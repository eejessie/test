1 0 0 2 0
2 4 1 0
2 5 1 0
1 1 0 2 0
2 6 1 1
2 15 1 1
1 2 0 2 0
2 26 1 2
2 28 1 2
1 3 0 2 0
2 29 1 3
2 30 1 3
2 31 1 11
2 32 1 11
2 33 1 12
2 34 1 12
2 35 1 17
2 36 1 17
2 37 1 20
2 38 1 20
2 39 1 23
2 40 1 23
0 7 5 1 1 4
0 8 5 1 1 6
0 9 5 1 1 26
0 10 5 1 1 29
0 11 7 2 2 5 28
0 12 5 2 1 31
0 13 7 1 2 7 9
0 14 5 1 1 13
3 77 7 0 2 33 14
0 16 7 1 2 15 30
0 17 5 2 1 16
0 18 7 1 2 8 10
0 19 5 1 1 18
0 20 7 2 2 35 19
0 21 5 1 1 37
0 22 7 1 2 32 38
0 23 5 2 1 22
0 24 7 1 2 34 21
0 25 5 1 1 24
3 78 7 0 2 39 25
0 27 7 1 2 36 40
3 79 5 0 1 27
