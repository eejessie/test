1 0 0 165 0
2 25 1 0
2 26 1 0
2 59236 1 0
2 59237 1 0
2 59238 1 0
2 59239 1 0
2 59240 1 0
2 59241 1 0
2 59242 1 0
2 59243 1 0
2 59244 1 0
2 59245 1 0
2 59246 1 0
2 59247 1 0
2 59248 1 0
2 59249 1 0
2 59250 1 0
2 59251 1 0
2 59252 1 0
2 59253 1 0
2 59254 1 0
2 59255 1 0
2 59256 1 0
2 59257 1 0
2 59258 1 0
2 59259 1 0
2 59260 1 0
2 59261 1 0
2 59262 1 0
2 59263 1 0
2 59264 1 0
2 59265 1 0
2 59266 1 0
2 59267 1 0
2 59268 1 0
2 59269 1 0
2 59270 1 0
2 59271 1 0
2 59272 1 0
2 59273 1 0
2 59274 1 0
2 59275 1 0
2 59276 1 0
2 59277 1 0
2 59278 1 0
2 59279 1 0
2 59280 1 0
2 59281 1 0
2 59282 1 0
2 59283 1 0
2 59284 1 0
2 59285 1 0
2 59286 1 0
2 59287 1 0
2 59288 1 0
2 59289 1 0
2 59290 1 0
2 59291 1 0
2 59292 1 0
2 59293 1 0
2 59294 1 0
2 59295 1 0
2 59296 1 0
2 59297 1 0
2 59298 1 0
2 59299 1 0
2 59300 1 0
2 59301 1 0
2 59302 1 0
2 59303 1 0
2 59304 1 0
2 59305 1 0
2 59306 1 0
2 59307 1 0
2 59308 1 0
2 59309 1 0
2 59310 1 0
2 59311 1 0
2 59312 1 0
2 59313 1 0
2 59314 1 0
2 59315 1 0
2 59316 1 0
2 59317 1 0
2 59318 1 0
2 59319 1 0
2 59320 1 0
2 59321 1 0
2 59322 1 0
2 59323 1 0
2 59324 1 0
2 59325 1 0
2 59326 1 0
2 59327 1 0
2 59328 1 0
2 59329 1 0
2 59330 1 0
2 59331 1 0
2 59332 1 0
2 59333 1 0
2 59334 1 0
2 59335 1 0
2 59336 1 0
2 59337 1 0
2 59338 1 0
2 59339 1 0
2 59340 1 0
2 59341 1 0
2 59342 1 0
2 59343 1 0
2 59344 1 0
2 59345 1 0
2 59346 1 0
2 59347 1 0
2 59348 1 0
2 59349 1 0
2 59350 1 0
2 59351 1 0
2 59352 1 0
2 59353 1 0
2 59354 1 0
2 59355 1 0
2 59356 1 0
2 59357 1 0
2 59358 1 0
2 59359 1 0
2 59360 1 0
2 59361 1 0
2 59362 1 0
2 59363 1 0
2 59364 1 0
2 59365 1 0
2 59366 1 0
2 59367 1 0
2 59368 1 0
2 59369 1 0
2 59370 1 0
2 59371 1 0
2 59372 1 0
2 59373 1 0
2 59374 1 0
2 59375 1 0
2 59376 1 0
2 59377 1 0
2 59378 1 0
2 59379 1 0
2 59380 1 0
2 59381 1 0
2 59382 1 0
2 59383 1 0
2 59384 1 0
2 59385 1 0
2 59386 1 0
2 59387 1 0
2 59388 1 0
2 59389 1 0
2 59390 1 0
2 59391 1 0
2 59392 1 0
2 59393 1 0
2 59394 1 0
2 59395 1 0
2 59396 1 0
2 59397 1 0
2 59398 1 0
1 1 0 325 0
2 59399 1 1
2 59400 1 1
2 59401 1 1
2 59402 1 1
2 59403 1 1
2 59404 1 1
2 59405 1 1
2 59406 1 1
2 59407 1 1
2 59408 1 1
2 59409 1 1
2 59410 1 1
2 59411 1 1
2 59412 1 1
2 59413 1 1
2 59414 1 1
2 59415 1 1
2 59416 1 1
2 59417 1 1
2 59418 1 1
2 59419 1 1
2 59420 1 1
2 59421 1 1
2 59422 1 1
2 59423 1 1
2 59424 1 1
2 59425 1 1
2 59426 1 1
2 59427 1 1
2 59428 1 1
2 59429 1 1
2 59430 1 1
2 59431 1 1
2 59432 1 1
2 59433 1 1
2 59434 1 1
2 59435 1 1
2 59436 1 1
2 59437 1 1
2 59438 1 1
2 59439 1 1
2 59440 1 1
2 59441 1 1
2 59442 1 1
2 59443 1 1
2 59444 1 1
2 59445 1 1
2 59446 1 1
2 59447 1 1
2 59448 1 1
2 59449 1 1
2 59450 1 1
2 59451 1 1
2 59452 1 1
2 59453 1 1
2 59454 1 1
2 59455 1 1
2 59456 1 1
2 59457 1 1
2 59458 1 1
2 59459 1 1
2 59460 1 1
2 59461 1 1
2 59462 1 1
2 59463 1 1
2 59464 1 1
2 59465 1 1
2 59466 1 1
2 59467 1 1
2 59468 1 1
2 59469 1 1
2 59470 1 1
2 59471 1 1
2 59472 1 1
2 59473 1 1
2 59474 1 1
2 59475 1 1
2 59476 1 1
2 59477 1 1
2 59478 1 1
2 59479 1 1
2 59480 1 1
2 59481 1 1
2 59482 1 1
2 59483 1 1
2 59484 1 1
2 59485 1 1
2 59486 1 1
2 59487 1 1
2 59488 1 1
2 59489 1 1
2 59490 1 1
2 59491 1 1
2 59492 1 1
2 59493 1 1
2 59494 1 1
2 59495 1 1
2 59496 1 1
2 59497 1 1
2 59498 1 1
2 59499 1 1
2 59500 1 1
2 59501 1 1
2 59502 1 1
2 59503 1 1
2 59504 1 1
2 59505 1 1
2 59506 1 1
2 59507 1 1
2 59508 1 1
2 59509 1 1
2 59510 1 1
2 59511 1 1
2 59512 1 1
2 59513 1 1
2 59514 1 1
2 59515 1 1
2 59516 1 1
2 59517 1 1
2 59518 1 1
2 59519 1 1
2 59520 1 1
2 59521 1 1
2 59522 1 1
2 59523 1 1
2 59524 1 1
2 59525 1 1
2 59526 1 1
2 59527 1 1
2 59528 1 1
2 59529 1 1
2 59530 1 1
2 59531 1 1
2 59532 1 1
2 59533 1 1
2 59534 1 1
2 59535 1 1
2 59536 1 1
2 59537 1 1
2 59538 1 1
2 59539 1 1
2 59540 1 1
2 59541 1 1
2 59542 1 1
2 59543 1 1
2 59544 1 1
2 59545 1 1
2 59546 1 1
2 59547 1 1
2 59548 1 1
2 59549 1 1
2 59550 1 1
2 59551 1 1
2 59552 1 1
2 59553 1 1
2 59554 1 1
2 59555 1 1
2 59556 1 1
2 59557 1 1
2 59558 1 1
2 59559 1 1
2 59560 1 1
2 59561 1 1
2 59562 1 1
2 59563 1 1
2 59564 1 1
2 59565 1 1
2 59566 1 1
2 59567 1 1
2 59568 1 1
2 59569 1 1
2 59570 1 1
2 59571 1 1
2 59572 1 1
2 59573 1 1
2 59574 1 1
2 59575 1 1
2 59576 1 1
2 59577 1 1
2 59578 1 1
2 59579 1 1
2 59580 1 1
2 59581 1 1
2 59582 1 1
2 59583 1 1
2 59584 1 1
2 59585 1 1
2 59586 1 1
2 59587 1 1
2 59588 1 1
2 59589 1 1
2 59590 1 1
2 59591 1 1
2 59592 1 1
2 59593 1 1
2 59594 1 1
2 59595 1 1
2 59596 1 1
2 59597 1 1
2 59598 1 1
2 59599 1 1
2 59600 1 1
2 59601 1 1
2 59602 1 1
2 59603 1 1
2 59604 1 1
2 59605 1 1
2 59606 1 1
2 59607 1 1
2 59608 1 1
2 59609 1 1
2 59610 1 1
2 59611 1 1
2 59612 1 1
2 59613 1 1
2 59614 1 1
2 59615 1 1
2 59616 1 1
2 59617 1 1
2 59618 1 1
2 59619 1 1
2 59620 1 1
2 59621 1 1
2 59622 1 1
2 59623 1 1
2 59624 1 1
2 59625 1 1
2 59626 1 1
2 59627 1 1
2 59628 1 1
2 59629 1 1
2 59630 1 1
2 59631 1 1
2 59632 1 1
2 59633 1 1
2 59634 1 1
2 59635 1 1
2 59636 1 1
2 59637 1 1
2 59638 1 1
2 59639 1 1
2 59640 1 1
2 59641 1 1
2 59642 1 1
2 59643 1 1
2 59644 1 1
2 59645 1 1
2 59646 1 1
2 59647 1 1
2 59648 1 1
2 59649 1 1
2 59650 1 1
2 59651 1 1
2 59652 1 1
2 59653 1 1
2 59654 1 1
2 59655 1 1
2 59656 1 1
2 59657 1 1
2 59658 1 1
2 59659 1 1
2 59660 1 1
2 59661 1 1
2 59662 1 1
2 59663 1 1
2 59664 1 1
2 59665 1 1
2 59666 1 1
2 59667 1 1
2 59668 1 1
2 59669 1 1
2 59670 1 1
2 59671 1 1
2 59672 1 1
2 59673 1 1
2 59674 1 1
2 59675 1 1
2 59676 1 1
2 59677 1 1
2 59678 1 1
2 59679 1 1
2 59680 1 1
2 59681 1 1
2 59682 1 1
2 59683 1 1
2 59684 1 1
2 59685 1 1
2 59686 1 1
2 59687 1 1
2 59688 1 1
2 59689 1 1
2 59690 1 1
2 59691 1 1
2 59692 1 1
2 59693 1 1
2 59694 1 1
2 59695 1 1
2 59696 1 1
2 59697 1 1
2 59698 1 1
2 59699 1 1
2 59700 1 1
2 59701 1 1
2 59702 1 1
2 59703 1 1
2 59704 1 1
2 59705 1 1
2 59706 1 1
2 59707 1 1
2 59708 1 1
2 59709 1 1
2 59710 1 1
2 59711 1 1
2 59712 1 1
2 59713 1 1
2 59714 1 1
2 59715 1 1
2 59716 1 1
2 59717 1 1
2 59718 1 1
2 59719 1 1
2 59720 1 1
2 59721 1 1
2 59722 1 1
2 59723 1 1
1 2 0 289 0
2 59724 1 2
2 59725 1 2
2 59726 1 2
2 59727 1 2
2 59728 1 2
2 59729 1 2
2 59730 1 2
2 59731 1 2
2 59732 1 2
2 59733 1 2
2 59734 1 2
2 59735 1 2
2 59736 1 2
2 59737 1 2
2 59738 1 2
2 59739 1 2
2 59740 1 2
2 59741 1 2
2 59742 1 2
2 59743 1 2
2 59744 1 2
2 59745 1 2
2 59746 1 2
2 59747 1 2
2 59748 1 2
2 59749 1 2
2 59750 1 2
2 59751 1 2
2 59752 1 2
2 59753 1 2
2 59754 1 2
2 59755 1 2
2 59756 1 2
2 59757 1 2
2 59758 1 2
2 59759 1 2
2 59760 1 2
2 59761 1 2
2 59762 1 2
2 59763 1 2
2 59764 1 2
2 59765 1 2
2 59766 1 2
2 59767 1 2
2 59768 1 2
2 59769 1 2
2 59770 1 2
2 59771 1 2
2 59772 1 2
2 59773 1 2
2 59774 1 2
2 59775 1 2
2 59776 1 2
2 59777 1 2
2 59778 1 2
2 59779 1 2
2 59780 1 2
2 59781 1 2
2 59782 1 2
2 59783 1 2
2 59784 1 2
2 59785 1 2
2 59786 1 2
2 59787 1 2
2 59788 1 2
2 59789 1 2
2 59790 1 2
2 59791 1 2
2 59792 1 2
2 59793 1 2
2 59794 1 2
2 59795 1 2
2 59796 1 2
2 59797 1 2
2 59798 1 2
2 59799 1 2
2 59800 1 2
2 59801 1 2
2 59802 1 2
2 59803 1 2
2 59804 1 2
2 59805 1 2
2 59806 1 2
2 59807 1 2
2 59808 1 2
2 59809 1 2
2 59810 1 2
2 59811 1 2
2 59812 1 2
2 59813 1 2
2 59814 1 2
2 59815 1 2
2 59816 1 2
2 59817 1 2
2 59818 1 2
2 59819 1 2
2 59820 1 2
2 59821 1 2
2 59822 1 2
2 59823 1 2
2 59824 1 2
2 59825 1 2
2 59826 1 2
2 59827 1 2
2 59828 1 2
2 59829 1 2
2 59830 1 2
2 59831 1 2
2 59832 1 2
2 59833 1 2
2 59834 1 2
2 59835 1 2
2 59836 1 2
2 59837 1 2
2 59838 1 2
2 59839 1 2
2 59840 1 2
2 59841 1 2
2 59842 1 2
2 59843 1 2
2 59844 1 2
2 59845 1 2
2 59846 1 2
2 59847 1 2
2 59848 1 2
2 59849 1 2
2 59850 1 2
2 59851 1 2
2 59852 1 2
2 59853 1 2
2 59854 1 2
2 59855 1 2
2 59856 1 2
2 59857 1 2
2 59858 1 2
2 59859 1 2
2 59860 1 2
2 59861 1 2
2 59862 1 2
2 59863 1 2
2 59864 1 2
2 59865 1 2
2 59866 1 2
2 59867 1 2
2 59868 1 2
2 59869 1 2
2 59870 1 2
2 59871 1 2
2 59872 1 2
2 59873 1 2
2 59874 1 2
2 59875 1 2
2 59876 1 2
2 59877 1 2
2 59878 1 2
2 59879 1 2
2 59880 1 2
2 59881 1 2
2 59882 1 2
2 59883 1 2
2 59884 1 2
2 59885 1 2
2 59886 1 2
2 59887 1 2
2 59888 1 2
2 59889 1 2
2 59890 1 2
2 59891 1 2
2 59892 1 2
2 59893 1 2
2 59894 1 2
2 59895 1 2
2 59896 1 2
2 59897 1 2
2 59898 1 2
2 59899 1 2
2 59900 1 2
2 59901 1 2
2 59902 1 2
2 59903 1 2
2 59904 1 2
2 59905 1 2
2 59906 1 2
2 59907 1 2
2 59908 1 2
2 59909 1 2
2 59910 1 2
2 59911 1 2
2 59912 1 2
2 59913 1 2
2 59914 1 2
2 59915 1 2
2 59916 1 2
2 59917 1 2
2 59918 1 2
2 59919 1 2
2 59920 1 2
2 59921 1 2
2 59922 1 2
2 59923 1 2
2 59924 1 2
2 59925 1 2
2 59926 1 2
2 59927 1 2
2 59928 1 2
2 59929 1 2
2 59930 1 2
2 59931 1 2
2 59932 1 2
2 59933 1 2
2 59934 1 2
2 59935 1 2
2 59936 1 2
2 59937 1 2
2 59938 1 2
2 59939 1 2
2 59940 1 2
2 59941 1 2
2 59942 1 2
2 59943 1 2
2 59944 1 2
2 59945 1 2
2 59946 1 2
2 59947 1 2
2 59948 1 2
2 59949 1 2
2 59950 1 2
2 59951 1 2
2 59952 1 2
2 59953 1 2
2 59954 1 2
2 59955 1 2
2 59956 1 2
2 59957 1 2
2 59958 1 2
2 59959 1 2
2 59960 1 2
2 59961 1 2
2 59962 1 2
2 59963 1 2
2 59964 1 2
2 59965 1 2
2 59966 1 2
2 59967 1 2
2 59968 1 2
2 59969 1 2
2 59970 1 2
2 59971 1 2
2 59972 1 2
2 59973 1 2
2 59974 1 2
2 59975 1 2
2 59976 1 2
2 59977 1 2
2 59978 1 2
2 59979 1 2
2 59980 1 2
2 59981 1 2
2 59982 1 2
2 59983 1 2
2 59984 1 2
2 59985 1 2
2 59986 1 2
2 59987 1 2
2 59988 1 2
2 59989 1 2
2 59990 1 2
2 59991 1 2
2 59992 1 2
2 59993 1 2
2 59994 1 2
2 59995 1 2
2 59996 1 2
2 59997 1 2
2 59998 1 2
2 59999 1 2
2 60000 1 2
2 60001 1 2
2 60002 1 2
2 60003 1 2
2 60004 1 2
2 60005 1 2
2 60006 1 2
2 60007 1 2
2 60008 1 2
2 60009 1 2
2 60010 1 2
2 60011 1 2
2 60012 1 2
1 3 0 171 0
2 60013 1 3
2 60014 1 3
2 60015 1 3
2 60016 1 3
2 60017 1 3
2 60018 1 3
2 60019 1 3
2 60020 1 3
2 60021 1 3
2 60022 1 3
2 60023 1 3
2 60024 1 3
2 60025 1 3
2 60026 1 3
2 60027 1 3
2 60028 1 3
2 60029 1 3
2 60030 1 3
2 60031 1 3
2 60032 1 3
2 60033 1 3
2 60034 1 3
2 60035 1 3
2 60036 1 3
2 60037 1 3
2 60038 1 3
2 60039 1 3
2 60040 1 3
2 60041 1 3
2 60042 1 3
2 60043 1 3
2 60044 1 3
2 60045 1 3
2 60046 1 3
2 60047 1 3
2 60048 1 3
2 60049 1 3
2 60050 1 3
2 60051 1 3
2 60052 1 3
2 60053 1 3
2 60054 1 3
2 60055 1 3
2 60056 1 3
2 60057 1 3
2 60058 1 3
2 60059 1 3
2 60060 1 3
2 60061 1 3
2 60062 1 3
2 60063 1 3
2 60064 1 3
2 60065 1 3
2 60066 1 3
2 60067 1 3
2 60068 1 3
2 60069 1 3
2 60070 1 3
2 60071 1 3
2 60072 1 3
2 60073 1 3
2 60074 1 3
2 60075 1 3
2 60076 1 3
2 60077 1 3
2 60078 1 3
2 60079 1 3
2 60080 1 3
2 60081 1 3
2 60082 1 3
2 60083 1 3
2 60084 1 3
2 60085 1 3
2 60086 1 3
2 60087 1 3
2 60088 1 3
2 60089 1 3
2 60090 1 3
2 60091 1 3
2 60092 1 3
2 60093 1 3
2 60094 1 3
2 60095 1 3
2 60096 1 3
2 60097 1 3
2 60098 1 3
2 60099 1 3
2 60100 1 3
2 60101 1 3
2 60102 1 3
2 60103 1 3
2 60104 1 3
2 60105 1 3
2 60106 1 3
2 60107 1 3
2 60108 1 3
2 60109 1 3
2 60110 1 3
2 60111 1 3
2 60112 1 3
2 60113 1 3
2 60114 1 3
2 60115 1 3
2 60116 1 3
2 60117 1 3
2 60118 1 3
2 60119 1 3
2 60120 1 3
2 60121 1 3
2 60122 1 3
2 60123 1 3
2 60124 1 3
2 60125 1 3
2 60126 1 3
2 60127 1 3
2 60128 1 3
2 60129 1 3
2 60130 1 3
2 60131 1 3
2 60132 1 3
2 60133 1 3
2 60134 1 3
2 60135 1 3
2 60136 1 3
2 60137 1 3
2 60138 1 3
2 60139 1 3
2 60140 1 3
2 60141 1 3
2 60142 1 3
2 60143 1 3
2 60144 1 3
2 60145 1 3
2 60146 1 3
2 60147 1 3
2 60148 1 3
2 60149 1 3
2 60150 1 3
2 60151 1 3
2 60152 1 3
2 60153 1 3
2 60154 1 3
2 60155 1 3
2 60156 1 3
2 60157 1 3
2 60158 1 3
2 60159 1 3
2 60160 1 3
2 60161 1 3
2 60162 1 3
2 60163 1 3
2 60164 1 3
2 60165 1 3
2 60166 1 3
2 60167 1 3
2 60168 1 3
2 60169 1 3
2 60170 1 3
2 60171 1 3
2 60172 1 3
2 60173 1 3
2 60174 1 3
2 60175 1 3
2 60176 1 3
2 60177 1 3
2 60178 1 3
2 60179 1 3
2 60180 1 3
2 60181 1 3
2 60182 1 3
2 60183 1 3
1 4 0 247 0
2 60184 1 4
2 60185 1 4
2 60186 1 4
2 60187 1 4
2 60188 1 4
2 60189 1 4
2 60190 1 4
2 60191 1 4
2 60192 1 4
2 60193 1 4
2 60194 1 4
2 60195 1 4
2 60196 1 4
2 60197 1 4
2 60198 1 4
2 60199 1 4
2 60200 1 4
2 60201 1 4
2 60202 1 4
2 60203 1 4
2 60204 1 4
2 60205 1 4
2 60206 1 4
2 60207 1 4
2 60208 1 4
2 60209 1 4
2 60210 1 4
2 60211 1 4
2 60212 1 4
2 60213 1 4
2 60214 1 4
2 60215 1 4
2 60216 1 4
2 60217 1 4
2 60218 1 4
2 60219 1 4
2 60220 1 4
2 60221 1 4
2 60222 1 4
2 60223 1 4
2 60224 1 4
2 60225 1 4
2 60226 1 4
2 60227 1 4
2 60228 1 4
2 60229 1 4
2 60230 1 4
2 60231 1 4
2 60232 1 4
2 60233 1 4
2 60234 1 4
2 60235 1 4
2 60236 1 4
2 60237 1 4
2 60238 1 4
2 60239 1 4
2 60240 1 4
2 60241 1 4
2 60242 1 4
2 60243 1 4
2 60244 1 4
2 60245 1 4
2 60246 1 4
2 60247 1 4
2 60248 1 4
2 60249 1 4
2 60250 1 4
2 60251 1 4
2 60252 1 4
2 60253 1 4
2 60254 1 4
2 60255 1 4
2 60256 1 4
2 60257 1 4
2 60258 1 4
2 60259 1 4
2 60260 1 4
2 60261 1 4
2 60262 1 4
2 60263 1 4
2 60264 1 4
2 60265 1 4
2 60266 1 4
2 60267 1 4
2 60268 1 4
2 60269 1 4
2 60270 1 4
2 60271 1 4
2 60272 1 4
2 60273 1 4
2 60274 1 4
2 60275 1 4
2 60276 1 4
2 60277 1 4
2 60278 1 4
2 60279 1 4
2 60280 1 4
2 60281 1 4
2 60282 1 4
2 60283 1 4
2 60284 1 4
2 60285 1 4
2 60286 1 4
2 60287 1 4
2 60288 1 4
2 60289 1 4
2 60290 1 4
2 60291 1 4
2 60292 1 4
2 60293 1 4
2 60294 1 4
2 60295 1 4
2 60296 1 4
2 60297 1 4
2 60298 1 4
2 60299 1 4
2 60300 1 4
2 60301 1 4
2 60302 1 4
2 60303 1 4
2 60304 1 4
2 60305 1 4
2 60306 1 4
2 60307 1 4
2 60308 1 4
2 60309 1 4
2 60310 1 4
2 60311 1 4
2 60312 1 4
2 60313 1 4
2 60314 1 4
2 60315 1 4
2 60316 1 4
2 60317 1 4
2 60318 1 4
2 60319 1 4
2 60320 1 4
2 60321 1 4
2 60322 1 4
2 60323 1 4
2 60324 1 4
2 60325 1 4
2 60326 1 4
2 60327 1 4
2 60328 1 4
2 60329 1 4
2 60330 1 4
2 60331 1 4
2 60332 1 4
2 60333 1 4
2 60334 1 4
2 60335 1 4
2 60336 1 4
2 60337 1 4
2 60338 1 4
2 60339 1 4
2 60340 1 4
2 60341 1 4
2 60342 1 4
2 60343 1 4
2 60344 1 4
2 60345 1 4
2 60346 1 4
2 60347 1 4
2 60348 1 4
2 60349 1 4
2 60350 1 4
2 60351 1 4
2 60352 1 4
2 60353 1 4
2 60354 1 4
2 60355 1 4
2 60356 1 4
2 60357 1 4
2 60358 1 4
2 60359 1 4
2 60360 1 4
2 60361 1 4
2 60362 1 4
2 60363 1 4
2 60364 1 4
2 60365 1 4
2 60366 1 4
2 60367 1 4
2 60368 1 4
2 60369 1 4
2 60370 1 4
2 60371 1 4
2 60372 1 4
2 60373 1 4
2 60374 1 4
2 60375 1 4
2 60376 1 4
2 60377 1 4
2 60378 1 4
2 60379 1 4
2 60380 1 4
2 60381 1 4
2 60382 1 4
2 60383 1 4
2 60384 1 4
2 60385 1 4
2 60386 1 4
2 60387 1 4
2 60388 1 4
2 60389 1 4
2 60390 1 4
2 60391 1 4
2 60392 1 4
2 60393 1 4
2 60394 1 4
2 60395 1 4
2 60396 1 4
2 60397 1 4
2 60398 1 4
2 60399 1 4
2 60400 1 4
2 60401 1 4
2 60402 1 4
2 60403 1 4
2 60404 1 4
2 60405 1 4
2 60406 1 4
2 60407 1 4
2 60408 1 4
2 60409 1 4
2 60410 1 4
2 60411 1 4
2 60412 1 4
2 60413 1 4
2 60414 1 4
2 60415 1 4
2 60416 1 4
2 60417 1 4
2 60418 1 4
2 60419 1 4
2 60420 1 4
2 60421 1 4
2 60422 1 4
2 60423 1 4
2 60424 1 4
2 60425 1 4
2 60426 1 4
2 60427 1 4
2 60428 1 4
2 60429 1 4
2 60430 1 4
1 5 0 214 0
2 60431 1 5
2 60432 1 5
2 60433 1 5
2 60434 1 5
2 60435 1 5
2 60436 1 5
2 60437 1 5
2 60438 1 5
2 60439 1 5
2 60440 1 5
2 60441 1 5
2 60442 1 5
2 60443 1 5
2 60444 1 5
2 60445 1 5
2 60446 1 5
2 60447 1 5
2 60448 1 5
2 60449 1 5
2 60450 1 5
2 60451 1 5
2 60452 1 5
2 60453 1 5
2 60454 1 5
2 60455 1 5
2 60456 1 5
2 60457 1 5
2 60458 1 5
2 60459 1 5
2 60460 1 5
2 60461 1 5
2 60462 1 5
2 60463 1 5
2 60464 1 5
2 60465 1 5
2 60466 1 5
2 60467 1 5
2 60468 1 5
2 60469 1 5
2 60470 1 5
2 60471 1 5
2 60472 1 5
2 60473 1 5
2 60474 1 5
2 60475 1 5
2 60476 1 5
2 60477 1 5
2 60478 1 5
2 60479 1 5
2 60480 1 5
2 60481 1 5
2 60482 1 5
2 60483 1 5
2 60484 1 5
2 60485 1 5
2 60486 1 5
2 60487 1 5
2 60488 1 5
2 60489 1 5
2 60490 1 5
2 60491 1 5
2 60492 1 5
2 60493 1 5
2 60494 1 5
2 60495 1 5
2 60496 1 5
2 60497 1 5
2 60498 1 5
2 60499 1 5
2 60500 1 5
2 60501 1 5
2 60502 1 5
2 60503 1 5
2 60504 1 5
2 60505 1 5
2 60506 1 5
2 60507 1 5
2 60508 1 5
2 60509 1 5
2 60510 1 5
2 60511 1 5
2 60512 1 5
2 60513 1 5
2 60514 1 5
2 60515 1 5
2 60516 1 5
2 60517 1 5
2 60518 1 5
2 60519 1 5
2 60520 1 5
2 60521 1 5
2 60522 1 5
2 60523 1 5
2 60524 1 5
2 60525 1 5
2 60526 1 5
2 60527 1 5
2 60528 1 5
2 60529 1 5
2 60530 1 5
2 60531 1 5
2 60532 1 5
2 60533 1 5
2 60534 1 5
2 60535 1 5
2 60536 1 5
2 60537 1 5
2 60538 1 5
2 60539 1 5
2 60540 1 5
2 60541 1 5
2 60542 1 5
2 60543 1 5
2 60544 1 5
2 60545 1 5
2 60546 1 5
2 60547 1 5
2 60548 1 5
2 60549 1 5
2 60550 1 5
2 60551 1 5
2 60552 1 5
2 60553 1 5
2 60554 1 5
2 60555 1 5
2 60556 1 5
2 60557 1 5
2 60558 1 5
2 60559 1 5
2 60560 1 5
2 60561 1 5
2 60562 1 5
2 60563 1 5
2 60564 1 5
2 60565 1 5
2 60566 1 5
2 60567 1 5
2 60568 1 5
2 60569 1 5
2 60570 1 5
2 60571 1 5
2 60572 1 5
2 60573 1 5
2 60574 1 5
2 60575 1 5
2 60576 1 5
2 60577 1 5
2 60578 1 5
2 60579 1 5
2 60580 1 5
2 60581 1 5
2 60582 1 5
2 60583 1 5
2 60584 1 5
2 60585 1 5
2 60586 1 5
2 60587 1 5
2 60588 1 5
2 60589 1 5
2 60590 1 5
2 60591 1 5
2 60592 1 5
2 60593 1 5
2 60594 1 5
2 60595 1 5
2 60596 1 5
2 60597 1 5
2 60598 1 5
2 60599 1 5
2 60600 1 5
2 60601 1 5
2 60602 1 5
2 60603 1 5
2 60604 1 5
2 60605 1 5
2 60606 1 5
2 60607 1 5
2 60608 1 5
2 60609 1 5
2 60610 1 5
2 60611 1 5
2 60612 1 5
2 60613 1 5
2 60614 1 5
2 60615 1 5
2 60616 1 5
2 60617 1 5
2 60618 1 5
2 60619 1 5
2 60620 1 5
2 60621 1 5
2 60622 1 5
2 60623 1 5
2 60624 1 5
2 60625 1 5
2 60626 1 5
2 60627 1 5
2 60628 1 5
2 60629 1 5
2 60630 1 5
2 60631 1 5
2 60632 1 5
2 60633 1 5
2 60634 1 5
2 60635 1 5
2 60636 1 5
2 60637 1 5
2 60638 1 5
2 60639 1 5
2 60640 1 5
2 60641 1 5
2 60642 1 5
2 60643 1 5
2 60644 1 5
1 6 0 103 0
2 60645 1 6
2 60646 1 6
2 60647 1 6
2 60648 1 6
2 60649 1 6
2 60650 1 6
2 60651 1 6
2 60652 1 6
2 60653 1 6
2 60654 1 6
2 60655 1 6
2 60656 1 6
2 60657 1 6
2 60658 1 6
2 60659 1 6
2 60660 1 6
2 60661 1 6
2 60662 1 6
2 60663 1 6
2 60664 1 6
2 60665 1 6
2 60666 1 6
2 60667 1 6
2 60668 1 6
2 60669 1 6
2 60670 1 6
2 60671 1 6
2 60672 1 6
2 60673 1 6
2 60674 1 6
2 60675 1 6
2 60676 1 6
2 60677 1 6
2 60678 1 6
2 60679 1 6
2 60680 1 6
2 60681 1 6
2 60682 1 6
2 60683 1 6
2 60684 1 6
2 60685 1 6
2 60686 1 6
2 60687 1 6
2 60688 1 6
2 60689 1 6
2 60690 1 6
2 60691 1 6
2 60692 1 6
2 60693 1 6
2 60694 1 6
2 60695 1 6
2 60696 1 6
2 60697 1 6
2 60698 1 6
2 60699 1 6
2 60700 1 6
2 60701 1 6
2 60702 1 6
2 60703 1 6
2 60704 1 6
2 60705 1 6
2 60706 1 6
2 60707 1 6
2 60708 1 6
2 60709 1 6
2 60710 1 6
2 60711 1 6
2 60712 1 6
2 60713 1 6
2 60714 1 6
2 60715 1 6
2 60716 1 6
2 60717 1 6
2 60718 1 6
2 60719 1 6
2 60720 1 6
2 60721 1 6
2 60722 1 6
2 60723 1 6
2 60724 1 6
2 60725 1 6
2 60726 1 6
2 60727 1 6
2 60728 1 6
2 60729 1 6
2 60730 1 6
2 60731 1 6
2 60732 1 6
2 60733 1 6
2 60734 1 6
2 60735 1 6
2 60736 1 6
2 60737 1 6
2 60738 1 6
2 60739 1 6
2 60740 1 6
2 60741 1 6
2 60742 1 6
2 60743 1 6
2 60744 1 6
2 60745 1 6
2 60746 1 6
2 60747 1 6
1 7 0 4 0
2 60748 1 7
2 60749 1 7
2 60750 1 7
2 60751 1 7
1 8 0 69 0
2 60752 1 8
2 60753 1 8
2 60754 1 8
2 60755 1 8
2 60756 1 8
2 60757 1 8
2 60758 1 8
2 60759 1 8
2 60760 1 8
2 60761 1 8
2 60762 1 8
2 60763 1 8
2 60764 1 8
2 60765 1 8
2 60766 1 8
2 60767 1 8
2 60768 1 8
2 60769 1 8
2 60770 1 8
2 60771 1 8
2 60772 1 8
2 60773 1 8
2 60774 1 8
2 60775 1 8
2 60776 1 8
2 60777 1 8
2 60778 1 8
2 60779 1 8
2 60780 1 8
2 60781 1 8
2 60782 1 8
2 60783 1 8
2 60784 1 8
2 60785 1 8
2 60786 1 8
2 60787 1 8
2 60788 1 8
2 60789 1 8
2 60790 1 8
2 60791 1 8
2 60792 1 8
2 60793 1 8
2 60794 1 8
2 60795 1 8
2 60796 1 8
2 60797 1 8
2 60798 1 8
2 60799 1 8
2 60800 1 8
2 60801 1 8
2 60802 1 8
2 60803 1 8
2 60804 1 8
2 60805 1 8
2 60806 1 8
2 60807 1 8
2 60808 1 8
2 60809 1 8
2 60810 1 8
2 60811 1 8
2 60812 1 8
2 60813 1 8
2 60814 1 8
2 60815 1 8
2 60816 1 8
2 60817 1 8
2 60818 1 8
2 60819 1 8
2 60820 1 8
1 9 0 147 0
2 60821 1 9
2 60822 1 9
2 60823 1 9
2 60824 1 9
2 60825 1 9
2 60826 1 9
2 60827 1 9
2 60828 1 9
2 60829 1 9
2 60830 1 9
2 60831 1 9
2 60832 1 9
2 60833 1 9
2 60834 1 9
2 60835 1 9
2 60836 1 9
2 60837 1 9
2 60838 1 9
2 60839 1 9
2 60840 1 9
2 60841 1 9
2 60842 1 9
2 60843 1 9
2 60844 1 9
2 60845 1 9
2 60846 1 9
2 60847 1 9
2 60848 1 9
2 60849 1 9
2 60850 1 9
2 60851 1 9
2 60852 1 9
2 60853 1 9
2 60854 1 9
2 60855 1 9
2 60856 1 9
2 60857 1 9
2 60858 1 9
2 60859 1 9
2 60860 1 9
2 60861 1 9
2 60862 1 9
2 60863 1 9
2 60864 1 9
2 60865 1 9
2 60866 1 9
2 60867 1 9
2 60868 1 9
2 60869 1 9
2 60870 1 9
2 60871 1 9
2 60872 1 9
2 60873 1 9
2 60874 1 9
2 60875 1 9
2 60876 1 9
2 60877 1 9
2 60878 1 9
2 60879 1 9
2 60880 1 9
2 60881 1 9
2 60882 1 9
2 60883 1 9
2 60884 1 9
2 60885 1 9
2 60886 1 9
2 60887 1 9
2 60888 1 9
2 60889 1 9
2 60890 1 9
2 60891 1 9
2 60892 1 9
2 60893 1 9
2 60894 1 9
2 60895 1 9
2 60896 1 9
2 60897 1 9
2 60898 1 9
2 60899 1 9
2 60900 1 9
2 60901 1 9
2 60902 1 9
2 60903 1 9
2 60904 1 9
2 60905 1 9
2 60906 1 9
2 60907 1 9
2 60908 1 9
2 60909 1 9
2 60910 1 9
2 60911 1 9
2 60912 1 9
2 60913 1 9
2 60914 1 9
2 60915 1 9
2 60916 1 9
2 60917 1 9
2 60918 1 9
2 60919 1 9
2 60920 1 9
2 60921 1 9
2 60922 1 9
2 60923 1 9
2 60924 1 9
2 60925 1 9
2 60926 1 9
2 60927 1 9
2 60928 1 9
2 60929 1 9
2 60930 1 9
2 60931 1 9
2 60932 1 9
2 60933 1 9
2 60934 1 9
2 60935 1 9
2 60936 1 9
2 60937 1 9
2 60938 1 9
2 60939 1 9
2 60940 1 9
2 60941 1 9
2 60942 1 9
2 60943 1 9
2 60944 1 9
2 60945 1 9
2 60946 1 9
2 60947 1 9
2 60948 1 9
2 60949 1 9
2 60950 1 9
2 60951 1 9
2 60952 1 9
2 60953 1 9
2 60954 1 9
2 60955 1 9
2 60956 1 9
2 60957 1 9
2 60958 1 9
2 60959 1 9
2 60960 1 9
2 60961 1 9
2 60962 1 9
2 60963 1 9
2 60964 1 9
2 60965 1 9
2 60966 1 9
2 60967 1 9
1 10 0 181 0
2 60968 1 10
2 60969 1 10
2 60970 1 10
2 60971 1 10
2 60972 1 10
2 60973 1 10
2 60974 1 10
2 60975 1 10
2 60976 1 10
2 60977 1 10
2 60978 1 10
2 60979 1 10
2 60980 1 10
2 60981 1 10
2 60982 1 10
2 60983 1 10
2 60984 1 10
2 60985 1 10
2 60986 1 10
2 60987 1 10
2 60988 1 10
2 60989 1 10
2 60990 1 10
2 60991 1 10
2 60992 1 10
2 60993 1 10
2 60994 1 10
2 60995 1 10
2 60996 1 10
2 60997 1 10
2 60998 1 10
2 60999 1 10
2 61000 1 10
2 61001 1 10
2 61002 1 10
2 61003 1 10
2 61004 1 10
2 61005 1 10
2 61006 1 10
2 61007 1 10
2 61008 1 10
2 61009 1 10
2 61010 1 10
2 61011 1 10
2 61012 1 10
2 61013 1 10
2 61014 1 10
2 61015 1 10
2 61016 1 10
2 61017 1 10
2 61018 1 10
2 61019 1 10
2 61020 1 10
2 61021 1 10
2 61022 1 10
2 61023 1 10
2 61024 1 10
2 61025 1 10
2 61026 1 10
2 61027 1 10
2 61028 1 10
2 61029 1 10
2 61030 1 10
2 61031 1 10
2 61032 1 10
2 61033 1 10
2 61034 1 10
2 61035 1 10
2 61036 1 10
2 61037 1 10
2 61038 1 10
2 61039 1 10
2 61040 1 10
2 61041 1 10
2 61042 1 10
2 61043 1 10
2 61044 1 10
2 61045 1 10
2 61046 1 10
2 61047 1 10
2 61048 1 10
2 61049 1 10
2 61050 1 10
2 61051 1 10
2 61052 1 10
2 61053 1 10
2 61054 1 10
2 61055 1 10
2 61056 1 10
2 61057 1 10
2 61058 1 10
2 61059 1 10
2 61060 1 10
2 61061 1 10
2 61062 1 10
2 61063 1 10
2 61064 1 10
2 61065 1 10
2 61066 1 10
2 61067 1 10
2 61068 1 10
2 61069 1 10
2 61070 1 10
2 61071 1 10
2 61072 1 10
2 61073 1 10
2 61074 1 10
2 61075 1 10
2 61076 1 10
2 61077 1 10
2 61078 1 10
2 61079 1 10
2 61080 1 10
2 61081 1 10
2 61082 1 10
2 61083 1 10
2 61084 1 10
2 61085 1 10
2 61086 1 10
2 61087 1 10
2 61088 1 10
2 61089 1 10
2 61090 1 10
2 61091 1 10
2 61092 1 10
2 61093 1 10
2 61094 1 10
2 61095 1 10
2 61096 1 10
2 61097 1 10
2 61098 1 10
2 61099 1 10
2 61100 1 10
2 61101 1 10
2 61102 1 10
2 61103 1 10
2 61104 1 10
2 61105 1 10
2 61106 1 10
2 61107 1 10
2 61108 1 10
2 61109 1 10
2 61110 1 10
2 61111 1 10
2 61112 1 10
2 61113 1 10
2 61114 1 10
2 61115 1 10
2 61116 1 10
2 61117 1 10
2 61118 1 10
2 61119 1 10
2 61120 1 10
2 61121 1 10
2 61122 1 10
2 61123 1 10
2 61124 1 10
2 61125 1 10
2 61126 1 10
2 61127 1 10
2 61128 1 10
2 61129 1 10
2 61130 1 10
2 61131 1 10
2 61132 1 10
2 61133 1 10
2 61134 1 10
2 61135 1 10
2 61136 1 10
2 61137 1 10
2 61138 1 10
2 61139 1 10
2 61140 1 10
2 61141 1 10
2 61142 1 10
2 61143 1 10
2 61144 1 10
2 61145 1 10
2 61146 1 10
2 61147 1 10
2 61148 1 10
1 11 0 227 0
2 61149 1 11
2 61150 1 11
2 61151 1 11
2 61152 1 11
2 61153 1 11
2 61154 1 11
2 61155 1 11
2 61156 1 11
2 61157 1 11
2 61158 1 11
2 61159 1 11
2 61160 1 11
2 61161 1 11
2 61162 1 11
2 61163 1 11
2 61164 1 11
2 61165 1 11
2 61166 1 11
2 61167 1 11
2 61168 1 11
2 61169 1 11
2 61170 1 11
2 61171 1 11
2 61172 1 11
2 61173 1 11
2 61174 1 11
2 61175 1 11
2 61176 1 11
2 61177 1 11
2 61178 1 11
2 61179 1 11
2 61180 1 11
2 61181 1 11
2 61182 1 11
2 61183 1 11
2 61184 1 11
2 61185 1 11
2 61186 1 11
2 61187 1 11
2 61188 1 11
2 61189 1 11
2 61190 1 11
2 61191 1 11
2 61192 1 11
2 61193 1 11
2 61194 1 11
2 61195 1 11
2 61196 1 11
2 61197 1 11
2 61198 1 11
2 61199 1 11
2 61200 1 11
2 61201 1 11
2 61202 1 11
2 61203 1 11
2 61204 1 11
2 61205 1 11
2 61206 1 11
2 61207 1 11
2 61208 1 11
2 61209 1 11
2 61210 1 11
2 61211 1 11
2 61212 1 11
2 61213 1 11
2 61214 1 11
2 61215 1 11
2 61216 1 11
2 61217 1 11
2 61218 1 11
2 61219 1 11
2 61220 1 11
2 61221 1 11
2 61222 1 11
2 61223 1 11
2 61224 1 11
2 61225 1 11
2 61226 1 11
2 61227 1 11
2 61228 1 11
2 61229 1 11
2 61230 1 11
2 61231 1 11
2 61232 1 11
2 61233 1 11
2 61234 1 11
2 61235 1 11
2 61236 1 11
2 61237 1 11
2 61238 1 11
2 61239 1 11
2 61240 1 11
2 61241 1 11
2 61242 1 11
2 61243 1 11
2 61244 1 11
2 61245 1 11
2 61246 1 11
2 61247 1 11
2 61248 1 11
2 61249 1 11
2 61250 1 11
2 61251 1 11
2 61252 1 11
2 61253 1 11
2 61254 1 11
2 61255 1 11
2 61256 1 11
2 61257 1 11
2 61258 1 11
2 61259 1 11
2 61260 1 11
2 61261 1 11
2 61262 1 11
2 61263 1 11
2 61264 1 11
2 61265 1 11
2 61266 1 11
2 61267 1 11
2 61268 1 11
2 61269 1 11
2 61270 1 11
2 61271 1 11
2 61272 1 11
2 61273 1 11
2 61274 1 11
2 61275 1 11
2 61276 1 11
2 61277 1 11
2 61278 1 11
2 61279 1 11
2 61280 1 11
2 61281 1 11
2 61282 1 11
2 61283 1 11
2 61284 1 11
2 61285 1 11
2 61286 1 11
2 61287 1 11
2 61288 1 11
2 61289 1 11
2 61290 1 11
2 61291 1 11
2 61292 1 11
2 61293 1 11
2 61294 1 11
2 61295 1 11
2 61296 1 11
2 61297 1 11
2 61298 1 11
2 61299 1 11
2 61300 1 11
2 61301 1 11
2 61302 1 11
2 61303 1 11
2 61304 1 11
2 61305 1 11
2 61306 1 11
2 61307 1 11
2 61308 1 11
2 61309 1 11
2 61310 1 11
2 61311 1 11
2 61312 1 11
2 61313 1 11
2 61314 1 11
2 61315 1 11
2 61316 1 11
2 61317 1 11
2 61318 1 11
2 61319 1 11
2 61320 1 11
2 61321 1 11
2 61322 1 11
2 61323 1 11
2 61324 1 11
2 61325 1 11
2 61326 1 11
2 61327 1 11
2 61328 1 11
2 61329 1 11
2 61330 1 11
2 61331 1 11
2 61332 1 11
2 61333 1 11
2 61334 1 11
2 61335 1 11
2 61336 1 11
2 61337 1 11
2 61338 1 11
2 61339 1 11
2 61340 1 11
2 61341 1 11
2 61342 1 11
2 61343 1 11
2 61344 1 11
2 61345 1 11
2 61346 1 11
2 61347 1 11
2 61348 1 11
2 61349 1 11
2 61350 1 11
2 61351 1 11
2 61352 1 11
2 61353 1 11
2 61354 1 11
2 61355 1 11
2 61356 1 11
2 61357 1 11
2 61358 1 11
2 61359 1 11
2 61360 1 11
2 61361 1 11
2 61362 1 11
2 61363 1 11
2 61364 1 11
2 61365 1 11
2 61366 1 11
2 61367 1 11
2 61368 1 11
2 61369 1 11
2 61370 1 11
2 61371 1 11
2 61372 1 11
2 61373 1 11
2 61374 1 11
2 61375 1 11
1 12 0 246 0
2 61376 1 12
2 61377 1 12
2 61378 1 12
2 61379 1 12
2 61380 1 12
2 61381 1 12
2 61382 1 12
2 61383 1 12
2 61384 1 12
2 61385 1 12
2 61386 1 12
2 61387 1 12
2 61388 1 12
2 61389 1 12
2 61390 1 12
2 61391 1 12
2 61392 1 12
2 61393 1 12
2 61394 1 12
2 61395 1 12
2 61396 1 12
2 61397 1 12
2 61398 1 12
2 61399 1 12
2 61400 1 12
2 61401 1 12
2 61402 1 12
2 61403 1 12
2 61404 1 12
2 61405 1 12
2 61406 1 12
2 61407 1 12
2 61408 1 12
2 61409 1 12
2 61410 1 12
2 61411 1 12
2 61412 1 12
2 61413 1 12
2 61414 1 12
2 61415 1 12
2 61416 1 12
2 61417 1 12
2 61418 1 12
2 61419 1 12
2 61420 1 12
2 61421 1 12
2 61422 1 12
2 61423 1 12
2 61424 1 12
2 61425 1 12
2 61426 1 12
2 61427 1 12
2 61428 1 12
2 61429 1 12
2 61430 1 12
2 61431 1 12
2 61432 1 12
2 61433 1 12
2 61434 1 12
2 61435 1 12
2 61436 1 12
2 61437 1 12
2 61438 1 12
2 61439 1 12
2 61440 1 12
2 61441 1 12
2 61442 1 12
2 61443 1 12
2 61444 1 12
2 61445 1 12
2 61446 1 12
2 61447 1 12
2 61448 1 12
2 61449 1 12
2 61450 1 12
2 61451 1 12
2 61452 1 12
2 61453 1 12
2 61454 1 12
2 61455 1 12
2 61456 1 12
2 61457 1 12
2 61458 1 12
2 61459 1 12
2 61460 1 12
2 61461 1 12
2 61462 1 12
2 61463 1 12
2 61464 1 12
2 61465 1 12
2 61466 1 12
2 61467 1 12
2 61468 1 12
2 61469 1 12
2 61470 1 12
2 61471 1 12
2 61472 1 12
2 61473 1 12
2 61474 1 12
2 61475 1 12
2 61476 1 12
2 61477 1 12
2 61478 1 12
2 61479 1 12
2 61480 1 12
2 61481 1 12
2 61482 1 12
2 61483 1 12
2 61484 1 12
2 61485 1 12
2 61486 1 12
2 61487 1 12
2 61488 1 12
2 61489 1 12
2 61490 1 12
2 61491 1 12
2 61492 1 12
2 61493 1 12
2 61494 1 12
2 61495 1 12
2 61496 1 12
2 61497 1 12
2 61498 1 12
2 61499 1 12
2 61500 1 12
2 61501 1 12
2 61502 1 12
2 61503 1 12
2 61504 1 12
2 61505 1 12
2 61506 1 12
2 61507 1 12
2 61508 1 12
2 61509 1 12
2 61510 1 12
2 61511 1 12
2 61512 1 12
2 61513 1 12
2 61514 1 12
2 61515 1 12
2 61516 1 12
2 61517 1 12
2 61518 1 12
2 61519 1 12
2 61520 1 12
2 61521 1 12
2 61522 1 12
2 61523 1 12
2 61524 1 12
2 61525 1 12
2 61526 1 12
2 61527 1 12
2 61528 1 12
2 61529 1 12
2 61530 1 12
2 61531 1 12
2 61532 1 12
2 61533 1 12
2 61534 1 12
2 61535 1 12
2 61536 1 12
2 61537 1 12
2 61538 1 12
2 61539 1 12
2 61540 1 12
2 61541 1 12
2 61542 1 12
2 61543 1 12
2 61544 1 12
2 61545 1 12
2 61546 1 12
2 61547 1 12
2 61548 1 12
2 61549 1 12
2 61550 1 12
2 61551 1 12
2 61552 1 12
2 61553 1 12
2 61554 1 12
2 61555 1 12
2 61556 1 12
2 61557 1 12
2 61558 1 12
2 61559 1 12
2 61560 1 12
2 61561 1 12
2 61562 1 12
2 61563 1 12
2 61564 1 12
2 61565 1 12
2 61566 1 12
2 61567 1 12
2 61568 1 12
2 61569 1 12
2 61570 1 12
2 61571 1 12
2 61572 1 12
2 61573 1 12
2 61574 1 12
2 61575 1 12
2 61576 1 12
2 61577 1 12
2 61578 1 12
2 61579 1 12
2 61580 1 12
2 61581 1 12
2 61582 1 12
2 61583 1 12
2 61584 1 12
2 61585 1 12
2 61586 1 12
2 61587 1 12
2 61588 1 12
2 61589 1 12
2 61590 1 12
2 61591 1 12
2 61592 1 12
2 61593 1 12
2 61594 1 12
2 61595 1 12
2 61596 1 12
2 61597 1 12
2 61598 1 12
2 61599 1 12
2 61600 1 12
2 61601 1 12
2 61602 1 12
2 61603 1 12
2 61604 1 12
2 61605 1 12
2 61606 1 12
2 61607 1 12
2 61608 1 12
2 61609 1 12
2 61610 1 12
2 61611 1 12
2 61612 1 12
2 61613 1 12
2 61614 1 12
2 61615 1 12
2 61616 1 12
2 61617 1 12
2 61618 1 12
2 61619 1 12
2 61620 1 12
2 61621 1 12
1 13 0 213 0
2 61622 1 13
2 61623 1 13
2 61624 1 13
2 61625 1 13
2 61626 1 13
2 61627 1 13
2 61628 1 13
2 61629 1 13
2 61630 1 13
2 61631 1 13
2 61632 1 13
2 61633 1 13
2 61634 1 13
2 61635 1 13
2 61636 1 13
2 61637 1 13
2 61638 1 13
2 61639 1 13
2 61640 1 13
2 61641 1 13
2 61642 1 13
2 61643 1 13
2 61644 1 13
2 61645 1 13
2 61646 1 13
2 61647 1 13
2 61648 1 13
2 61649 1 13
2 61650 1 13
2 61651 1 13
2 61652 1 13
2 61653 1 13
2 61654 1 13
2 61655 1 13
2 61656 1 13
2 61657 1 13
2 61658 1 13
2 61659 1 13
2 61660 1 13
2 61661 1 13
2 61662 1 13
2 61663 1 13
2 61664 1 13
2 61665 1 13
2 61666 1 13
2 61667 1 13
2 61668 1 13
2 61669 1 13
2 61670 1 13
2 61671 1 13
2 61672 1 13
2 61673 1 13
2 61674 1 13
2 61675 1 13
2 61676 1 13
2 61677 1 13
2 61678 1 13
2 61679 1 13
2 61680 1 13
2 61681 1 13
2 61682 1 13
2 61683 1 13
2 61684 1 13
2 61685 1 13
2 61686 1 13
2 61687 1 13
2 61688 1 13
2 61689 1 13
2 61690 1 13
2 61691 1 13
2 61692 1 13
2 61693 1 13
2 61694 1 13
2 61695 1 13
2 61696 1 13
2 61697 1 13
2 61698 1 13
2 61699 1 13
2 61700 1 13
2 61701 1 13
2 61702 1 13
2 61703 1 13
2 61704 1 13
2 61705 1 13
2 61706 1 13
2 61707 1 13
2 61708 1 13
2 61709 1 13
2 61710 1 13
2 61711 1 13
2 61712 1 13
2 61713 1 13
2 61714 1 13
2 61715 1 13
2 61716 1 13
2 61717 1 13
2 61718 1 13
2 61719 1 13
2 61720 1 13
2 61721 1 13
2 61722 1 13
2 61723 1 13
2 61724 1 13
2 61725 1 13
2 61726 1 13
2 61727 1 13
2 61728 1 13
2 61729 1 13
2 61730 1 13
2 61731 1 13
2 61732 1 13
2 61733 1 13
2 61734 1 13
2 61735 1 13
2 61736 1 13
2 61737 1 13
2 61738 1 13
2 61739 1 13
2 61740 1 13
2 61741 1 13
2 61742 1 13
2 61743 1 13
2 61744 1 13
2 61745 1 13
2 61746 1 13
2 61747 1 13
2 61748 1 13
2 61749 1 13
2 61750 1 13
2 61751 1 13
2 61752 1 13
2 61753 1 13
2 61754 1 13
2 61755 1 13
2 61756 1 13
2 61757 1 13
2 61758 1 13
2 61759 1 13
2 61760 1 13
2 61761 1 13
2 61762 1 13
2 61763 1 13
2 61764 1 13
2 61765 1 13
2 61766 1 13
2 61767 1 13
2 61768 1 13
2 61769 1 13
2 61770 1 13
2 61771 1 13
2 61772 1 13
2 61773 1 13
2 61774 1 13
2 61775 1 13
2 61776 1 13
2 61777 1 13
2 61778 1 13
2 61779 1 13
2 61780 1 13
2 61781 1 13
2 61782 1 13
2 61783 1 13
2 61784 1 13
2 61785 1 13
2 61786 1 13
2 61787 1 13
2 61788 1 13
2 61789 1 13
2 61790 1 13
2 61791 1 13
2 61792 1 13
2 61793 1 13
2 61794 1 13
2 61795 1 13
2 61796 1 13
2 61797 1 13
2 61798 1 13
2 61799 1 13
2 61800 1 13
2 61801 1 13
2 61802 1 13
2 61803 1 13
2 61804 1 13
2 61805 1 13
2 61806 1 13
2 61807 1 13
2 61808 1 13
2 61809 1 13
2 61810 1 13
2 61811 1 13
2 61812 1 13
2 61813 1 13
2 61814 1 13
2 61815 1 13
2 61816 1 13
2 61817 1 13
2 61818 1 13
2 61819 1 13
2 61820 1 13
2 61821 1 13
2 61822 1 13
2 61823 1 13
2 61824 1 13
2 61825 1 13
2 61826 1 13
2 61827 1 13
2 61828 1 13
2 61829 1 13
2 61830 1 13
2 61831 1 13
2 61832 1 13
2 61833 1 13
2 61834 1 13
1 14 0 126 0
2 61835 1 14
2 61836 1 14
2 61837 1 14
2 61838 1 14
2 61839 1 14
2 61840 1 14
2 61841 1 14
2 61842 1 14
2 61843 1 14
2 61844 1 14
2 61845 1 14
2 61846 1 14
2 61847 1 14
2 61848 1 14
2 61849 1 14
2 61850 1 14
2 61851 1 14
2 61852 1 14
2 61853 1 14
2 61854 1 14
2 61855 1 14
2 61856 1 14
2 61857 1 14
2 61858 1 14
2 61859 1 14
2 61860 1 14
2 61861 1 14
2 61862 1 14
2 61863 1 14
2 61864 1 14
2 61865 1 14
2 61866 1 14
2 61867 1 14
2 61868 1 14
2 61869 1 14
2 61870 1 14
2 61871 1 14
2 61872 1 14
2 61873 1 14
2 61874 1 14
2 61875 1 14
2 61876 1 14
2 61877 1 14
2 61878 1 14
2 61879 1 14
2 61880 1 14
2 61881 1 14
2 61882 1 14
2 61883 1 14
2 61884 1 14
2 61885 1 14
2 61886 1 14
2 61887 1 14
2 61888 1 14
2 61889 1 14
2 61890 1 14
2 61891 1 14
2 61892 1 14
2 61893 1 14
2 61894 1 14
2 61895 1 14
2 61896 1 14
2 61897 1 14
2 61898 1 14
2 61899 1 14
2 61900 1 14
2 61901 1 14
2 61902 1 14
2 61903 1 14
2 61904 1 14
2 61905 1 14
2 61906 1 14
2 61907 1 14
2 61908 1 14
2 61909 1 14
2 61910 1 14
2 61911 1 14
2 61912 1 14
2 61913 1 14
2 61914 1 14
2 61915 1 14
2 61916 1 14
2 61917 1 14
2 61918 1 14
2 61919 1 14
2 61920 1 14
2 61921 1 14
2 61922 1 14
2 61923 1 14
2 61924 1 14
2 61925 1 14
2 61926 1 14
2 61927 1 14
2 61928 1 14
2 61929 1 14
2 61930 1 14
2 61931 1 14
2 61932 1 14
2 61933 1 14
2 61934 1 14
2 61935 1 14
2 61936 1 14
2 61937 1 14
2 61938 1 14
2 61939 1 14
2 61940 1 14
2 61941 1 14
2 61942 1 14
2 61943 1 14
2 61944 1 14
2 61945 1 14
2 61946 1 14
2 61947 1 14
2 61948 1 14
2 61949 1 14
2 61950 1 14
2 61951 1 14
2 61952 1 14
2 61953 1 14
2 61954 1 14
2 61955 1 14
2 61956 1 14
2 61957 1 14
2 61958 1 14
2 61959 1 14
2 61960 1 14
1 15 0 5 0
2 61961 1 15
2 61962 1 15
2 61963 1 15
2 61964 1 15
2 61965 1 15
1 16 0 201 0
2 61966 1 16
2 61967 1 16
2 61968 1 16
2 61969 1 16
2 61970 1 16
2 61971 1 16
2 61972 1 16
2 61973 1 16
2 61974 1 16
2 61975 1 16
2 61976 1 16
2 61977 1 16
2 61978 1 16
2 61979 1 16
2 61980 1 16
2 61981 1 16
2 61982 1 16
2 61983 1 16
2 61984 1 16
2 61985 1 16
2 61986 1 16
2 61987 1 16
2 61988 1 16
2 61989 1 16
2 61990 1 16
2 61991 1 16
2 61992 1 16
2 61993 1 16
2 61994 1 16
2 61995 1 16
2 61996 1 16
2 61997 1 16
2 61998 1 16
2 61999 1 16
2 62000 1 16
2 62001 1 16
2 62002 1 16
2 62003 1 16
2 62004 1 16
2 62005 1 16
2 62006 1 16
2 62007 1 16
2 62008 1 16
2 62009 1 16
2 62010 1 16
2 62011 1 16
2 62012 1 16
2 62013 1 16
2 62014 1 16
2 62015 1 16
2 62016 1 16
2 62017 1 16
2 62018 1 16
2 62019 1 16
2 62020 1 16
2 62021 1 16
2 62022 1 16
2 62023 1 16
2 62024 1 16
2 62025 1 16
2 62026 1 16
2 62027 1 16
2 62028 1 16
2 62029 1 16
2 62030 1 16
2 62031 1 16
2 62032 1 16
2 62033 1 16
2 62034 1 16
2 62035 1 16
2 62036 1 16
2 62037 1 16
2 62038 1 16
2 62039 1 16
2 62040 1 16
2 62041 1 16
2 62042 1 16
2 62043 1 16
2 62044 1 16
2 62045 1 16
2 62046 1 16
2 62047 1 16
2 62048 1 16
2 62049 1 16
2 62050 1 16
2 62051 1 16
2 62052 1 16
2 62053 1 16
2 62054 1 16
2 62055 1 16
2 62056 1 16
2 62057 1 16
2 62058 1 16
2 62059 1 16
2 62060 1 16
2 62061 1 16
2 62062 1 16
2 62063 1 16
2 62064 1 16
2 62065 1 16
2 62066 1 16
2 62067 1 16
2 62068 1 16
2 62069 1 16
2 62070 1 16
2 62071 1 16
2 62072 1 16
2 62073 1 16
2 62074 1 16
2 62075 1 16
2 62076 1 16
2 62077 1 16
2 62078 1 16
2 62079 1 16
2 62080 1 16
2 62081 1 16
2 62082 1 16
2 62083 1 16
2 62084 1 16
2 62085 1 16
2 62086 1 16
2 62087 1 16
2 62088 1 16
2 62089 1 16
2 62090 1 16
2 62091 1 16
2 62092 1 16
2 62093 1 16
2 62094 1 16
2 62095 1 16
2 62096 1 16
2 62097 1 16
2 62098 1 16
2 62099 1 16
2 62100 1 16
2 62101 1 16
2 62102 1 16
2 62103 1 16
2 62104 1 16
2 62105 1 16
2 62106 1 16
2 62107 1 16
2 62108 1 16
2 62109 1 16
2 62110 1 16
2 62111 1 16
2 62112 1 16
2 62113 1 16
2 62114 1 16
2 62115 1 16
2 62116 1 16
2 62117 1 16
2 62118 1 16
2 62119 1 16
2 62120 1 16
2 62121 1 16
2 62122 1 16
2 62123 1 16
2 62124 1 16
2 62125 1 16
2 62126 1 16
2 62127 1 16
2 62128 1 16
2 62129 1 16
2 62130 1 16
2 62131 1 16
2 62132 1 16
2 62133 1 16
2 62134 1 16
2 62135 1 16
2 62136 1 16
2 62137 1 16
2 62138 1 16
2 62139 1 16
2 62140 1 16
2 62141 1 16
2 62142 1 16
2 62143 1 16
2 62144 1 16
2 62145 1 16
2 62146 1 16
2 62147 1 16
2 62148 1 16
2 62149 1 16
2 62150 1 16
2 62151 1 16
2 62152 1 16
2 62153 1 16
2 62154 1 16
2 62155 1 16
2 62156 1 16
2 62157 1 16
2 62158 1 16
2 62159 1 16
2 62160 1 16
2 62161 1 16
2 62162 1 16
2 62163 1 16
2 62164 1 16
2 62165 1 16
2 62166 1 16
1 17 0 247 0
2 62167 1 17
2 62168 1 17
2 62169 1 17
2 62170 1 17
2 62171 1 17
2 62172 1 17
2 62173 1 17
2 62174 1 17
2 62175 1 17
2 62176 1 17
2 62177 1 17
2 62178 1 17
2 62179 1 17
2 62180 1 17
2 62181 1 17
2 62182 1 17
2 62183 1 17
2 62184 1 17
2 62185 1 17
2 62186 1 17
2 62187 1 17
2 62188 1 17
2 62189 1 17
2 62190 1 17
2 62191 1 17
2 62192 1 17
2 62193 1 17
2 62194 1 17
2 62195 1 17
2 62196 1 17
2 62197 1 17
2 62198 1 17
2 62199 1 17
2 62200 1 17
2 62201 1 17
2 62202 1 17
2 62203 1 17
2 62204 1 17
2 62205 1 17
2 62206 1 17
2 62207 1 17
2 62208 1 17
2 62209 1 17
2 62210 1 17
2 62211 1 17
2 62212 1 17
2 62213 1 17
2 62214 1 17
2 62215 1 17
2 62216 1 17
2 62217 1 17
2 62218 1 17
2 62219 1 17
2 62220 1 17
2 62221 1 17
2 62222 1 17
2 62223 1 17
2 62224 1 17
2 62225 1 17
2 62226 1 17
2 62227 1 17
2 62228 1 17
2 62229 1 17
2 62230 1 17
2 62231 1 17
2 62232 1 17
2 62233 1 17
2 62234 1 17
2 62235 1 17
2 62236 1 17
2 62237 1 17
2 62238 1 17
2 62239 1 17
2 62240 1 17
2 62241 1 17
2 62242 1 17
2 62243 1 17
2 62244 1 17
2 62245 1 17
2 62246 1 17
2 62247 1 17
2 62248 1 17
2 62249 1 17
2 62250 1 17
2 62251 1 17
2 62252 1 17
2 62253 1 17
2 62254 1 17
2 62255 1 17
2 62256 1 17
2 62257 1 17
2 62258 1 17
2 62259 1 17
2 62260 1 17
2 62261 1 17
2 62262 1 17
2 62263 1 17
2 62264 1 17
2 62265 1 17
2 62266 1 17
2 62267 1 17
2 62268 1 17
2 62269 1 17
2 62270 1 17
2 62271 1 17
2 62272 1 17
2 62273 1 17
2 62274 1 17
2 62275 1 17
2 62276 1 17
2 62277 1 17
2 62278 1 17
2 62279 1 17
2 62280 1 17
2 62281 1 17
2 62282 1 17
2 62283 1 17
2 62284 1 17
2 62285 1 17
2 62286 1 17
2 62287 1 17
2 62288 1 17
2 62289 1 17
2 62290 1 17
2 62291 1 17
2 62292 1 17
2 62293 1 17
2 62294 1 17
2 62295 1 17
2 62296 1 17
2 62297 1 17
2 62298 1 17
2 62299 1 17
2 62300 1 17
2 62301 1 17
2 62302 1 17
2 62303 1 17
2 62304 1 17
2 62305 1 17
2 62306 1 17
2 62307 1 17
2 62308 1 17
2 62309 1 17
2 62310 1 17
2 62311 1 17
2 62312 1 17
2 62313 1 17
2 62314 1 17
2 62315 1 17
2 62316 1 17
2 62317 1 17
2 62318 1 17
2 62319 1 17
2 62320 1 17
2 62321 1 17
2 62322 1 17
2 62323 1 17
2 62324 1 17
2 62325 1 17
2 62326 1 17
2 62327 1 17
2 62328 1 17
2 62329 1 17
2 62330 1 17
2 62331 1 17
2 62332 1 17
2 62333 1 17
2 62334 1 17
2 62335 1 17
2 62336 1 17
2 62337 1 17
2 62338 1 17
2 62339 1 17
2 62340 1 17
2 62341 1 17
2 62342 1 17
2 62343 1 17
2 62344 1 17
2 62345 1 17
2 62346 1 17
2 62347 1 17
2 62348 1 17
2 62349 1 17
2 62350 1 17
2 62351 1 17
2 62352 1 17
2 62353 1 17
2 62354 1 17
2 62355 1 17
2 62356 1 17
2 62357 1 17
2 62358 1 17
2 62359 1 17
2 62360 1 17
2 62361 1 17
2 62362 1 17
2 62363 1 17
2 62364 1 17
2 62365 1 17
2 62366 1 17
2 62367 1 17
2 62368 1 17
2 62369 1 17
2 62370 1 17
2 62371 1 17
2 62372 1 17
2 62373 1 17
2 62374 1 17
2 62375 1 17
2 62376 1 17
2 62377 1 17
2 62378 1 17
2 62379 1 17
2 62380 1 17
2 62381 1 17
2 62382 1 17
2 62383 1 17
2 62384 1 17
2 62385 1 17
2 62386 1 17
2 62387 1 17
2 62388 1 17
2 62389 1 17
2 62390 1 17
2 62391 1 17
2 62392 1 17
2 62393 1 17
2 62394 1 17
2 62395 1 17
2 62396 1 17
2 62397 1 17
2 62398 1 17
2 62399 1 17
2 62400 1 17
2 62401 1 17
2 62402 1 17
2 62403 1 17
2 62404 1 17
2 62405 1 17
2 62406 1 17
2 62407 1 17
2 62408 1 17
2 62409 1 17
2 62410 1 17
2 62411 1 17
2 62412 1 17
2 62413 1 17
1 18 0 384 0
2 62414 1 18
2 62415 1 18
2 62416 1 18
2 62417 1 18
2 62418 1 18
2 62419 1 18
2 62420 1 18
2 62421 1 18
2 62422 1 18
2 62423 1 18
2 62424 1 18
2 62425 1 18
2 62426 1 18
2 62427 1 18
2 62428 1 18
2 62429 1 18
2 62430 1 18
2 62431 1 18
2 62432 1 18
2 62433 1 18
2 62434 1 18
2 62435 1 18
2 62436 1 18
2 62437 1 18
2 62438 1 18
2 62439 1 18
2 62440 1 18
2 62441 1 18
2 62442 1 18
2 62443 1 18
2 62444 1 18
2 62445 1 18
2 62446 1 18
2 62447 1 18
2 62448 1 18
2 62449 1 18
2 62450 1 18
2 62451 1 18
2 62452 1 18
2 62453 1 18
2 62454 1 18
2 62455 1 18
2 62456 1 18
2 62457 1 18
2 62458 1 18
2 62459 1 18
2 62460 1 18
2 62461 1 18
2 62462 1 18
2 62463 1 18
2 62464 1 18
2 62465 1 18
2 62466 1 18
2 62467 1 18
2 62468 1 18
2 62469 1 18
2 62470 1 18
2 62471 1 18
2 62472 1 18
2 62473 1 18
2 62474 1 18
2 62475 1 18
2 62476 1 18
2 62477 1 18
2 62478 1 18
2 62479 1 18
2 62480 1 18
2 62481 1 18
2 62482 1 18
2 62483 1 18
2 62484 1 18
2 62485 1 18
2 62486 1 18
2 62487 1 18
2 62488 1 18
2 62489 1 18
2 62490 1 18
2 62491 1 18
2 62492 1 18
2 62493 1 18
2 62494 1 18
2 62495 1 18
2 62496 1 18
2 62497 1 18
2 62498 1 18
2 62499 1 18
2 62500 1 18
2 62501 1 18
2 62502 1 18
2 62503 1 18
2 62504 1 18
2 62505 1 18
2 62506 1 18
2 62507 1 18
2 62508 1 18
2 62509 1 18
2 62510 1 18
2 62511 1 18
2 62512 1 18
2 62513 1 18
2 62514 1 18
2 62515 1 18
2 62516 1 18
2 62517 1 18
2 62518 1 18
2 62519 1 18
2 62520 1 18
2 62521 1 18
2 62522 1 18
2 62523 1 18
2 62524 1 18
2 62525 1 18
2 62526 1 18
2 62527 1 18
2 62528 1 18
2 62529 1 18
2 62530 1 18
2 62531 1 18
2 62532 1 18
2 62533 1 18
2 62534 1 18
2 62535 1 18
2 62536 1 18
2 62537 1 18
2 62538 1 18
2 62539 1 18
2 62540 1 18
2 62541 1 18
2 62542 1 18
2 62543 1 18
2 62544 1 18
2 62545 1 18
2 62546 1 18
2 62547 1 18
2 62548 1 18
2 62549 1 18
2 62550 1 18
2 62551 1 18
2 62552 1 18
2 62553 1 18
2 62554 1 18
2 62555 1 18
2 62556 1 18
2 62557 1 18
2 62558 1 18
2 62559 1 18
2 62560 1 18
2 62561 1 18
2 62562 1 18
2 62563 1 18
2 62564 1 18
2 62565 1 18
2 62566 1 18
2 62567 1 18
2 62568 1 18
2 62569 1 18
2 62570 1 18
2 62571 1 18
2 62572 1 18
2 62573 1 18
2 62574 1 18
2 62575 1 18
2 62576 1 18
2 62577 1 18
2 62578 1 18
2 62579 1 18
2 62580 1 18
2 62581 1 18
2 62582 1 18
2 62583 1 18
2 62584 1 18
2 62585 1 18
2 62586 1 18
2 62587 1 18
2 62588 1 18
2 62589 1 18
2 62590 1 18
2 62591 1 18
2 62592 1 18
2 62593 1 18
2 62594 1 18
2 62595 1 18
2 62596 1 18
2 62597 1 18
2 62598 1 18
2 62599 1 18
2 62600 1 18
2 62601 1 18
2 62602 1 18
2 62603 1 18
2 62604 1 18
2 62605 1 18
2 62606 1 18
2 62607 1 18
2 62608 1 18
2 62609 1 18
2 62610 1 18
2 62611 1 18
2 62612 1 18
2 62613 1 18
2 62614 1 18
2 62615 1 18
2 62616 1 18
2 62617 1 18
2 62618 1 18
2 62619 1 18
2 62620 1 18
2 62621 1 18
2 62622 1 18
2 62623 1 18
2 62624 1 18
2 62625 1 18
2 62626 1 18
2 62627 1 18
2 62628 1 18
2 62629 1 18
2 62630 1 18
2 62631 1 18
2 62632 1 18
2 62633 1 18
2 62634 1 18
2 62635 1 18
2 62636 1 18
2 62637 1 18
2 62638 1 18
2 62639 1 18
2 62640 1 18
2 62641 1 18
2 62642 1 18
2 62643 1 18
2 62644 1 18
2 62645 1 18
2 62646 1 18
2 62647 1 18
2 62648 1 18
2 62649 1 18
2 62650 1 18
2 62651 1 18
2 62652 1 18
2 62653 1 18
2 62654 1 18
2 62655 1 18
2 62656 1 18
2 62657 1 18
2 62658 1 18
2 62659 1 18
2 62660 1 18
2 62661 1 18
2 62662 1 18
2 62663 1 18
2 62664 1 18
2 62665 1 18
2 62666 1 18
2 62667 1 18
2 62668 1 18
2 62669 1 18
2 62670 1 18
2 62671 1 18
2 62672 1 18
2 62673 1 18
2 62674 1 18
2 62675 1 18
2 62676 1 18
2 62677 1 18
2 62678 1 18
2 62679 1 18
2 62680 1 18
2 62681 1 18
2 62682 1 18
2 62683 1 18
2 62684 1 18
2 62685 1 18
2 62686 1 18
2 62687 1 18
2 62688 1 18
2 62689 1 18
2 62690 1 18
2 62691 1 18
2 62692 1 18
2 62693 1 18
2 62694 1 18
2 62695 1 18
2 62696 1 18
2 62697 1 18
2 62698 1 18
2 62699 1 18
2 62700 1 18
2 62701 1 18
2 62702 1 18
2 62703 1 18
2 62704 1 18
2 62705 1 18
2 62706 1 18
2 62707 1 18
2 62708 1 18
2 62709 1 18
2 62710 1 18
2 62711 1 18
2 62712 1 18
2 62713 1 18
2 62714 1 18
2 62715 1 18
2 62716 1 18
2 62717 1 18
2 62718 1 18
2 62719 1 18
2 62720 1 18
2 62721 1 18
2 62722 1 18
2 62723 1 18
2 62724 1 18
2 62725 1 18
2 62726 1 18
2 62727 1 18
2 62728 1 18
2 62729 1 18
2 62730 1 18
2 62731 1 18
2 62732 1 18
2 62733 1 18
2 62734 1 18
2 62735 1 18
2 62736 1 18
2 62737 1 18
2 62738 1 18
2 62739 1 18
2 62740 1 18
2 62741 1 18
2 62742 1 18
2 62743 1 18
2 62744 1 18
2 62745 1 18
2 62746 1 18
2 62747 1 18
2 62748 1 18
2 62749 1 18
2 62750 1 18
2 62751 1 18
2 62752 1 18
2 62753 1 18
2 62754 1 18
2 62755 1 18
2 62756 1 18
2 62757 1 18
2 62758 1 18
2 62759 1 18
2 62760 1 18
2 62761 1 18
2 62762 1 18
2 62763 1 18
2 62764 1 18
2 62765 1 18
2 62766 1 18
2 62767 1 18
2 62768 1 18
2 62769 1 18
2 62770 1 18
2 62771 1 18
2 62772 1 18
2 62773 1 18
2 62774 1 18
2 62775 1 18
2 62776 1 18
2 62777 1 18
2 62778 1 18
2 62779 1 18
2 62780 1 18
2 62781 1 18
2 62782 1 18
2 62783 1 18
2 62784 1 18
2 62785 1 18
2 62786 1 18
2 62787 1 18
2 62788 1 18
2 62789 1 18
2 62790 1 18
2 62791 1 18
2 62792 1 18
2 62793 1 18
2 62794 1 18
2 62795 1 18
2 62796 1 18
2 62797 1 18
1 19 0 454 0
2 62798 1 19
2 62799 1 19
2 62800 1 19
2 62801 1 19
2 62802 1 19
2 62803 1 19
2 62804 1 19
2 62805 1 19
2 62806 1 19
2 62807 1 19
2 62808 1 19
2 62809 1 19
2 62810 1 19
2 62811 1 19
2 62812 1 19
2 62813 1 19
2 62814 1 19
2 62815 1 19
2 62816 1 19
2 62817 1 19
2 62818 1 19
2 62819 1 19
2 62820 1 19
2 62821 1 19
2 62822 1 19
2 62823 1 19
2 62824 1 19
2 62825 1 19
2 62826 1 19
2 62827 1 19
2 62828 1 19
2 62829 1 19
2 62830 1 19
2 62831 1 19
2 62832 1 19
2 62833 1 19
2 62834 1 19
2 62835 1 19
2 62836 1 19
2 62837 1 19
2 62838 1 19
2 62839 1 19
2 62840 1 19
2 62841 1 19
2 62842 1 19
2 62843 1 19
2 62844 1 19
2 62845 1 19
2 62846 1 19
2 62847 1 19
2 62848 1 19
2 62849 1 19
2 62850 1 19
2 62851 1 19
2 62852 1 19
2 62853 1 19
2 62854 1 19
2 62855 1 19
2 62856 1 19
2 62857 1 19
2 62858 1 19
2 62859 1 19
2 62860 1 19
2 62861 1 19
2 62862 1 19
2 62863 1 19
2 62864 1 19
2 62865 1 19
2 62866 1 19
2 62867 1 19
2 62868 1 19
2 62869 1 19
2 62870 1 19
2 62871 1 19
2 62872 1 19
2 62873 1 19
2 62874 1 19
2 62875 1 19
2 62876 1 19
2 62877 1 19
2 62878 1 19
2 62879 1 19
2 62880 1 19
2 62881 1 19
2 62882 1 19
2 62883 1 19
2 62884 1 19
2 62885 1 19
2 62886 1 19
2 62887 1 19
2 62888 1 19
2 62889 1 19
2 62890 1 19
2 62891 1 19
2 62892 1 19
2 62893 1 19
2 62894 1 19
2 62895 1 19
2 62896 1 19
2 62897 1 19
2 62898 1 19
2 62899 1 19
2 62900 1 19
2 62901 1 19
2 62902 1 19
2 62903 1 19
2 62904 1 19
2 62905 1 19
2 62906 1 19
2 62907 1 19
2 62908 1 19
2 62909 1 19
2 62910 1 19
2 62911 1 19
2 62912 1 19
2 62913 1 19
2 62914 1 19
2 62915 1 19
2 62916 1 19
2 62917 1 19
2 62918 1 19
2 62919 1 19
2 62920 1 19
2 62921 1 19
2 62922 1 19
2 62923 1 19
2 62924 1 19
2 62925 1 19
2 62926 1 19
2 62927 1 19
2 62928 1 19
2 62929 1 19
2 62930 1 19
2 62931 1 19
2 62932 1 19
2 62933 1 19
2 62934 1 19
2 62935 1 19
2 62936 1 19
2 62937 1 19
2 62938 1 19
2 62939 1 19
2 62940 1 19
2 62941 1 19
2 62942 1 19
2 62943 1 19
2 62944 1 19
2 62945 1 19
2 62946 1 19
2 62947 1 19
2 62948 1 19
2 62949 1 19
2 62950 1 19
2 62951 1 19
2 62952 1 19
2 62953 1 19
2 62954 1 19
2 62955 1 19
2 62956 1 19
2 62957 1 19
2 62958 1 19
2 62959 1 19
2 62960 1 19
2 62961 1 19
2 62962 1 19
2 62963 1 19
2 62964 1 19
2 62965 1 19
2 62966 1 19
2 62967 1 19
2 62968 1 19
2 62969 1 19
2 62970 1 19
2 62971 1 19
2 62972 1 19
2 62973 1 19
2 62974 1 19
2 62975 1 19
2 62976 1 19
2 62977 1 19
2 62978 1 19
2 62979 1 19
2 62980 1 19
2 62981 1 19
2 62982 1 19
2 62983 1 19
2 62984 1 19
2 62985 1 19
2 62986 1 19
2 62987 1 19
2 62988 1 19
2 62989 1 19
2 62990 1 19
2 62991 1 19
2 62992 1 19
2 62993 1 19
2 62994 1 19
2 62995 1 19
2 62996 1 19
2 62997 1 19
2 62998 1 19
2 62999 1 19
2 63000 1 19
2 63001 1 19
2 63002 1 19
2 63003 1 19
2 63004 1 19
2 63005 1 19
2 63006 1 19
2 63007 1 19
2 63008 1 19
2 63009 1 19
2 63010 1 19
2 63011 1 19
2 63012 1 19
2 63013 1 19
2 63014 1 19
2 63015 1 19
2 63016 1 19
2 63017 1 19
2 63018 1 19
2 63019 1 19
2 63020 1 19
2 63021 1 19
2 63022 1 19
2 63023 1 19
2 63024 1 19
2 63025 1 19
2 63026 1 19
2 63027 1 19
2 63028 1 19
2 63029 1 19
2 63030 1 19
2 63031 1 19
2 63032 1 19
2 63033 1 19
2 63034 1 19
2 63035 1 19
2 63036 1 19
2 63037 1 19
2 63038 1 19
2 63039 1 19
2 63040 1 19
2 63041 1 19
2 63042 1 19
2 63043 1 19
2 63044 1 19
2 63045 1 19
2 63046 1 19
2 63047 1 19
2 63048 1 19
2 63049 1 19
2 63050 1 19
2 63051 1 19
2 63052 1 19
2 63053 1 19
2 63054 1 19
2 63055 1 19
2 63056 1 19
2 63057 1 19
2 63058 1 19
2 63059 1 19
2 63060 1 19
2 63061 1 19
2 63062 1 19
2 63063 1 19
2 63064 1 19
2 63065 1 19
2 63066 1 19
2 63067 1 19
2 63068 1 19
2 63069 1 19
2 63070 1 19
2 63071 1 19
2 63072 1 19
2 63073 1 19
2 63074 1 19
2 63075 1 19
2 63076 1 19
2 63077 1 19
2 63078 1 19
2 63079 1 19
2 63080 1 19
2 63081 1 19
2 63082 1 19
2 63083 1 19
2 63084 1 19
2 63085 1 19
2 63086 1 19
2 63087 1 19
2 63088 1 19
2 63089 1 19
2 63090 1 19
2 63091 1 19
2 63092 1 19
2 63093 1 19
2 63094 1 19
2 63095 1 19
2 63096 1 19
2 63097 1 19
2 63098 1 19
2 63099 1 19
2 63100 1 19
2 63101 1 19
2 63102 1 19
2 63103 1 19
2 63104 1 19
2 63105 1 19
2 63106 1 19
2 63107 1 19
2 63108 1 19
2 63109 1 19
2 63110 1 19
2 63111 1 19
2 63112 1 19
2 63113 1 19
2 63114 1 19
2 63115 1 19
2 63116 1 19
2 63117 1 19
2 63118 1 19
2 63119 1 19
2 63120 1 19
2 63121 1 19
2 63122 1 19
2 63123 1 19
2 63124 1 19
2 63125 1 19
2 63126 1 19
2 63127 1 19
2 63128 1 19
2 63129 1 19
2 63130 1 19
2 63131 1 19
2 63132 1 19
2 63133 1 19
2 63134 1 19
2 63135 1 19
2 63136 1 19
2 63137 1 19
2 63138 1 19
2 63139 1 19
2 63140 1 19
2 63141 1 19
2 63142 1 19
2 63143 1 19
2 63144 1 19
2 63145 1 19
2 63146 1 19
2 63147 1 19
2 63148 1 19
2 63149 1 19
2 63150 1 19
2 63151 1 19
2 63152 1 19
2 63153 1 19
2 63154 1 19
2 63155 1 19
2 63156 1 19
2 63157 1 19
2 63158 1 19
2 63159 1 19
2 63160 1 19
2 63161 1 19
2 63162 1 19
2 63163 1 19
2 63164 1 19
2 63165 1 19
2 63166 1 19
2 63167 1 19
2 63168 1 19
2 63169 1 19
2 63170 1 19
2 63171 1 19
2 63172 1 19
2 63173 1 19
2 63174 1 19
2 63175 1 19
2 63176 1 19
2 63177 1 19
2 63178 1 19
2 63179 1 19
2 63180 1 19
2 63181 1 19
2 63182 1 19
2 63183 1 19
2 63184 1 19
2 63185 1 19
2 63186 1 19
2 63187 1 19
2 63188 1 19
2 63189 1 19
2 63190 1 19
2 63191 1 19
2 63192 1 19
2 63193 1 19
2 63194 1 19
2 63195 1 19
2 63196 1 19
2 63197 1 19
2 63198 1 19
2 63199 1 19
2 63200 1 19
2 63201 1 19
2 63202 1 19
2 63203 1 19
2 63204 1 19
2 63205 1 19
2 63206 1 19
2 63207 1 19
2 63208 1 19
2 63209 1 19
2 63210 1 19
2 63211 1 19
2 63212 1 19
2 63213 1 19
2 63214 1 19
2 63215 1 19
2 63216 1 19
2 63217 1 19
2 63218 1 19
2 63219 1 19
2 63220 1 19
2 63221 1 19
2 63222 1 19
2 63223 1 19
2 63224 1 19
2 63225 1 19
2 63226 1 19
2 63227 1 19
2 63228 1 19
2 63229 1 19
2 63230 1 19
2 63231 1 19
2 63232 1 19
2 63233 1 19
2 63234 1 19
2 63235 1 19
2 63236 1 19
2 63237 1 19
2 63238 1 19
2 63239 1 19
2 63240 1 19
2 63241 1 19
2 63242 1 19
2 63243 1 19
2 63244 1 19
2 63245 1 19
2 63246 1 19
2 63247 1 19
2 63248 1 19
2 63249 1 19
2 63250 1 19
2 63251 1 19
1 20 0 368 0
2 63252 1 20
2 63253 1 20
2 63254 1 20
2 63255 1 20
2 63256 1 20
2 63257 1 20
2 63258 1 20
2 63259 1 20
2 63260 1 20
2 63261 1 20
2 63262 1 20
2 63263 1 20
2 63264 1 20
2 63265 1 20
2 63266 1 20
2 63267 1 20
2 63268 1 20
2 63269 1 20
2 63270 1 20
2 63271 1 20
2 63272 1 20
2 63273 1 20
2 63274 1 20
2 63275 1 20
2 63276 1 20
2 63277 1 20
2 63278 1 20
2 63279 1 20
2 63280 1 20
2 63281 1 20
2 63282 1 20
2 63283 1 20
2 63284 1 20
2 63285 1 20
2 63286 1 20
2 63287 1 20
2 63288 1 20
2 63289 1 20
2 63290 1 20
2 63291 1 20
2 63292 1 20
2 63293 1 20
2 63294 1 20
2 63295 1 20
2 63296 1 20
2 63297 1 20
2 63298 1 20
2 63299 1 20
2 63300 1 20
2 63301 1 20
2 63302 1 20
2 63303 1 20
2 63304 1 20
2 63305 1 20
2 63306 1 20
2 63307 1 20
2 63308 1 20
2 63309 1 20
2 63310 1 20
2 63311 1 20
2 63312 1 20
2 63313 1 20
2 63314 1 20
2 63315 1 20
2 63316 1 20
2 63317 1 20
2 63318 1 20
2 63319 1 20
2 63320 1 20
2 63321 1 20
2 63322 1 20
2 63323 1 20
2 63324 1 20
2 63325 1 20
2 63326 1 20
2 63327 1 20
2 63328 1 20
2 63329 1 20
2 63330 1 20
2 63331 1 20
2 63332 1 20
2 63333 1 20
2 63334 1 20
2 63335 1 20
2 63336 1 20
2 63337 1 20
2 63338 1 20
2 63339 1 20
2 63340 1 20
2 63341 1 20
2 63342 1 20
2 63343 1 20
2 63344 1 20
2 63345 1 20
2 63346 1 20
2 63347 1 20
2 63348 1 20
2 63349 1 20
2 63350 1 20
2 63351 1 20
2 63352 1 20
2 63353 1 20
2 63354 1 20
2 63355 1 20
2 63356 1 20
2 63357 1 20
2 63358 1 20
2 63359 1 20
2 63360 1 20
2 63361 1 20
2 63362 1 20
2 63363 1 20
2 63364 1 20
2 63365 1 20
2 63366 1 20
2 63367 1 20
2 63368 1 20
2 63369 1 20
2 63370 1 20
2 63371 1 20
2 63372 1 20
2 63373 1 20
2 63374 1 20
2 63375 1 20
2 63376 1 20
2 63377 1 20
2 63378 1 20
2 63379 1 20
2 63380 1 20
2 63381 1 20
2 63382 1 20
2 63383 1 20
2 63384 1 20
2 63385 1 20
2 63386 1 20
2 63387 1 20
2 63388 1 20
2 63389 1 20
2 63390 1 20
2 63391 1 20
2 63392 1 20
2 63393 1 20
2 63394 1 20
2 63395 1 20
2 63396 1 20
2 63397 1 20
2 63398 1 20
2 63399 1 20
2 63400 1 20
2 63401 1 20
2 63402 1 20
2 63403 1 20
2 63404 1 20
2 63405 1 20
2 63406 1 20
2 63407 1 20
2 63408 1 20
2 63409 1 20
2 63410 1 20
2 63411 1 20
2 63412 1 20
2 63413 1 20
2 63414 1 20
2 63415 1 20
2 63416 1 20
2 63417 1 20
2 63418 1 20
2 63419 1 20
2 63420 1 20
2 63421 1 20
2 63422 1 20
2 63423 1 20
2 63424 1 20
2 63425 1 20
2 63426 1 20
2 63427 1 20
2 63428 1 20
2 63429 1 20
2 63430 1 20
2 63431 1 20
2 63432 1 20
2 63433 1 20
2 63434 1 20
2 63435 1 20
2 63436 1 20
2 63437 1 20
2 63438 1 20
2 63439 1 20
2 63440 1 20
2 63441 1 20
2 63442 1 20
2 63443 1 20
2 63444 1 20
2 63445 1 20
2 63446 1 20
2 63447 1 20
2 63448 1 20
2 63449 1 20
2 63450 1 20
2 63451 1 20
2 63452 1 20
2 63453 1 20
2 63454 1 20
2 63455 1 20
2 63456 1 20
2 63457 1 20
2 63458 1 20
2 63459 1 20
2 63460 1 20
2 63461 1 20
2 63462 1 20
2 63463 1 20
2 63464 1 20
2 63465 1 20
2 63466 1 20
2 63467 1 20
2 63468 1 20
2 63469 1 20
2 63470 1 20
2 63471 1 20
2 63472 1 20
2 63473 1 20
2 63474 1 20
2 63475 1 20
2 63476 1 20
2 63477 1 20
2 63478 1 20
2 63479 1 20
2 63480 1 20
2 63481 1 20
2 63482 1 20
2 63483 1 20
2 63484 1 20
2 63485 1 20
2 63486 1 20
2 63487 1 20
2 63488 1 20
2 63489 1 20
2 63490 1 20
2 63491 1 20
2 63492 1 20
2 63493 1 20
2 63494 1 20
2 63495 1 20
2 63496 1 20
2 63497 1 20
2 63498 1 20
2 63499 1 20
2 63500 1 20
2 63501 1 20
2 63502 1 20
2 63503 1 20
2 63504 1 20
2 63505 1 20
2 63506 1 20
2 63507 1 20
2 63508 1 20
2 63509 1 20
2 63510 1 20
2 63511 1 20
2 63512 1 20
2 63513 1 20
2 63514 1 20
2 63515 1 20
2 63516 1 20
2 63517 1 20
2 63518 1 20
2 63519 1 20
2 63520 1 20
2 63521 1 20
2 63522 1 20
2 63523 1 20
2 63524 1 20
2 63525 1 20
2 63526 1 20
2 63527 1 20
2 63528 1 20
2 63529 1 20
2 63530 1 20
2 63531 1 20
2 63532 1 20
2 63533 1 20
2 63534 1 20
2 63535 1 20
2 63536 1 20
2 63537 1 20
2 63538 1 20
2 63539 1 20
2 63540 1 20
2 63541 1 20
2 63542 1 20
2 63543 1 20
2 63544 1 20
2 63545 1 20
2 63546 1 20
2 63547 1 20
2 63548 1 20
2 63549 1 20
2 63550 1 20
2 63551 1 20
2 63552 1 20
2 63553 1 20
2 63554 1 20
2 63555 1 20
2 63556 1 20
2 63557 1 20
2 63558 1 20
2 63559 1 20
2 63560 1 20
2 63561 1 20
2 63562 1 20
2 63563 1 20
2 63564 1 20
2 63565 1 20
2 63566 1 20
2 63567 1 20
2 63568 1 20
2 63569 1 20
2 63570 1 20
2 63571 1 20
2 63572 1 20
2 63573 1 20
2 63574 1 20
2 63575 1 20
2 63576 1 20
2 63577 1 20
2 63578 1 20
2 63579 1 20
2 63580 1 20
2 63581 1 20
2 63582 1 20
2 63583 1 20
2 63584 1 20
2 63585 1 20
2 63586 1 20
2 63587 1 20
2 63588 1 20
2 63589 1 20
2 63590 1 20
2 63591 1 20
2 63592 1 20
2 63593 1 20
2 63594 1 20
2 63595 1 20
2 63596 1 20
2 63597 1 20
2 63598 1 20
2 63599 1 20
2 63600 1 20
2 63601 1 20
2 63602 1 20
2 63603 1 20
2 63604 1 20
2 63605 1 20
2 63606 1 20
2 63607 1 20
2 63608 1 20
2 63609 1 20
2 63610 1 20
2 63611 1 20
2 63612 1 20
2 63613 1 20
2 63614 1 20
2 63615 1 20
2 63616 1 20
2 63617 1 20
2 63618 1 20
2 63619 1 20
1 21 0 264 0
2 63620 1 21
2 63621 1 21
2 63622 1 21
2 63623 1 21
2 63624 1 21
2 63625 1 21
2 63626 1 21
2 63627 1 21
2 63628 1 21
2 63629 1 21
2 63630 1 21
2 63631 1 21
2 63632 1 21
2 63633 1 21
2 63634 1 21
2 63635 1 21
2 63636 1 21
2 63637 1 21
2 63638 1 21
2 63639 1 21
2 63640 1 21
2 63641 1 21
2 63642 1 21
2 63643 1 21
2 63644 1 21
2 63645 1 21
2 63646 1 21
2 63647 1 21
2 63648 1 21
2 63649 1 21
2 63650 1 21
2 63651 1 21
2 63652 1 21
2 63653 1 21
2 63654 1 21
2 63655 1 21
2 63656 1 21
2 63657 1 21
2 63658 1 21
2 63659 1 21
2 63660 1 21
2 63661 1 21
2 63662 1 21
2 63663 1 21
2 63664 1 21
2 63665 1 21
2 63666 1 21
2 63667 1 21
2 63668 1 21
2 63669 1 21
2 63670 1 21
2 63671 1 21
2 63672 1 21
2 63673 1 21
2 63674 1 21
2 63675 1 21
2 63676 1 21
2 63677 1 21
2 63678 1 21
2 63679 1 21
2 63680 1 21
2 63681 1 21
2 63682 1 21
2 63683 1 21
2 63684 1 21
2 63685 1 21
2 63686 1 21
2 63687 1 21
2 63688 1 21
2 63689 1 21
2 63690 1 21
2 63691 1 21
2 63692 1 21
2 63693 1 21
2 63694 1 21
2 63695 1 21
2 63696 1 21
2 63697 1 21
2 63698 1 21
2 63699 1 21
2 63700 1 21
2 63701 1 21
2 63702 1 21
2 63703 1 21
2 63704 1 21
2 63705 1 21
2 63706 1 21
2 63707 1 21
2 63708 1 21
2 63709 1 21
2 63710 1 21
2 63711 1 21
2 63712 1 21
2 63713 1 21
2 63714 1 21
2 63715 1 21
2 63716 1 21
2 63717 1 21
2 63718 1 21
2 63719 1 21
2 63720 1 21
2 63721 1 21
2 63722 1 21
2 63723 1 21
2 63724 1 21
2 63725 1 21
2 63726 1 21
2 63727 1 21
2 63728 1 21
2 63729 1 21
2 63730 1 21
2 63731 1 21
2 63732 1 21
2 63733 1 21
2 63734 1 21
2 63735 1 21
2 63736 1 21
2 63737 1 21
2 63738 1 21
2 63739 1 21
2 63740 1 21
2 63741 1 21
2 63742 1 21
2 63743 1 21
2 63744 1 21
2 63745 1 21
2 63746 1 21
2 63747 1 21
2 63748 1 21
2 63749 1 21
2 63750 1 21
2 63751 1 21
2 63752 1 21
2 63753 1 21
2 63754 1 21
2 63755 1 21
2 63756 1 21
2 63757 1 21
2 63758 1 21
2 63759 1 21
2 63760 1 21
2 63761 1 21
2 63762 1 21
2 63763 1 21
2 63764 1 21
2 63765 1 21
2 63766 1 21
2 63767 1 21
2 63768 1 21
2 63769 1 21
2 63770 1 21
2 63771 1 21
2 63772 1 21
2 63773 1 21
2 63774 1 21
2 63775 1 21
2 63776 1 21
2 63777 1 21
2 63778 1 21
2 63779 1 21
2 63780 1 21
2 63781 1 21
2 63782 1 21
2 63783 1 21
2 63784 1 21
2 63785 1 21
2 63786 1 21
2 63787 1 21
2 63788 1 21
2 63789 1 21
2 63790 1 21
2 63791 1 21
2 63792 1 21
2 63793 1 21
2 63794 1 21
2 63795 1 21
2 63796 1 21
2 63797 1 21
2 63798 1 21
2 63799 1 21
2 63800 1 21
2 63801 1 21
2 63802 1 21
2 63803 1 21
2 63804 1 21
2 63805 1 21
2 63806 1 21
2 63807 1 21
2 63808 1 21
2 63809 1 21
2 63810 1 21
2 63811 1 21
2 63812 1 21
2 63813 1 21
2 63814 1 21
2 63815 1 21
2 63816 1 21
2 63817 1 21
2 63818 1 21
2 63819 1 21
2 63820 1 21
2 63821 1 21
2 63822 1 21
2 63823 1 21
2 63824 1 21
2 63825 1 21
2 63826 1 21
2 63827 1 21
2 63828 1 21
2 63829 1 21
2 63830 1 21
2 63831 1 21
2 63832 1 21
2 63833 1 21
2 63834 1 21
2 63835 1 21
2 63836 1 21
2 63837 1 21
2 63838 1 21
2 63839 1 21
2 63840 1 21
2 63841 1 21
2 63842 1 21
2 63843 1 21
2 63844 1 21
2 63845 1 21
2 63846 1 21
2 63847 1 21
2 63848 1 21
2 63849 1 21
2 63850 1 21
2 63851 1 21
2 63852 1 21
2 63853 1 21
2 63854 1 21
2 63855 1 21
2 63856 1 21
2 63857 1 21
2 63858 1 21
2 63859 1 21
2 63860 1 21
2 63861 1 21
2 63862 1 21
2 63863 1 21
2 63864 1 21
2 63865 1 21
2 63866 1 21
2 63867 1 21
2 63868 1 21
2 63869 1 21
2 63870 1 21
2 63871 1 21
2 63872 1 21
2 63873 1 21
2 63874 1 21
2 63875 1 21
2 63876 1 21
2 63877 1 21
2 63878 1 21
2 63879 1 21
2 63880 1 21
2 63881 1 21
2 63882 1 21
2 63883 1 21
1 22 0 204 0
2 63884 1 22
2 63885 1 22
2 63886 1 22
2 63887 1 22
2 63888 1 22
2 63889 1 22
2 63890 1 22
2 63891 1 22
2 63892 1 22
2 63893 1 22
2 63894 1 22
2 63895 1 22
2 63896 1 22
2 63897 1 22
2 63898 1 22
2 63899 1 22
2 63900 1 22
2 63901 1 22
2 63902 1 22
2 63903 1 22
2 63904 1 22
2 63905 1 22
2 63906 1 22
2 63907 1 22
2 63908 1 22
2 63909 1 22
2 63910 1 22
2 63911 1 22
2 63912 1 22
2 63913 1 22
2 63914 1 22
2 63915 1 22
2 63916 1 22
2 63917 1 22
2 63918 1 22
2 63919 1 22
2 63920 1 22
2 63921 1 22
2 63922 1 22
2 63923 1 22
2 63924 1 22
2 63925 1 22
2 63926 1 22
2 63927 1 22
2 63928 1 22
2 63929 1 22
2 63930 1 22
2 63931 1 22
2 63932 1 22
2 63933 1 22
2 63934 1 22
2 63935 1 22
2 63936 1 22
2 63937 1 22
2 63938 1 22
2 63939 1 22
2 63940 1 22
2 63941 1 22
2 63942 1 22
2 63943 1 22
2 63944 1 22
2 63945 1 22
2 63946 1 22
2 63947 1 22
2 63948 1 22
2 63949 1 22
2 63950 1 22
2 63951 1 22
2 63952 1 22
2 63953 1 22
2 63954 1 22
2 63955 1 22
2 63956 1 22
2 63957 1 22
2 63958 1 22
2 63959 1 22
2 63960 1 22
2 63961 1 22
2 63962 1 22
2 63963 1 22
2 63964 1 22
2 63965 1 22
2 63966 1 22
2 63967 1 22
2 63968 1 22
2 63969 1 22
2 63970 1 22
2 63971 1 22
2 63972 1 22
2 63973 1 22
2 63974 1 22
2 63975 1 22
2 63976 1 22
2 63977 1 22
2 63978 1 22
2 63979 1 22
2 63980 1 22
2 63981 1 22
2 63982 1 22
2 63983 1 22
2 63984 1 22
2 63985 1 22
2 63986 1 22
2 63987 1 22
2 63988 1 22
2 63989 1 22
2 63990 1 22
2 63991 1 22
2 63992 1 22
2 63993 1 22
2 63994 1 22
2 63995 1 22
2 63996 1 22
2 63997 1 22
2 63998 1 22
2 63999 1 22
2 64000 1 22
2 64001 1 22
2 64002 1 22
2 64003 1 22
2 64004 1 22
2 64005 1 22
2 64006 1 22
2 64007 1 22
2 64008 1 22
2 64009 1 22
2 64010 1 22
2 64011 1 22
2 64012 1 22
2 64013 1 22
2 64014 1 22
2 64015 1 22
2 64016 1 22
2 64017 1 22
2 64018 1 22
2 64019 1 22
2 64020 1 22
2 64021 1 22
2 64022 1 22
2 64023 1 22
2 64024 1 22
2 64025 1 22
2 64026 1 22
2 64027 1 22
2 64028 1 22
2 64029 1 22
2 64030 1 22
2 64031 1 22
2 64032 1 22
2 64033 1 22
2 64034 1 22
2 64035 1 22
2 64036 1 22
2 64037 1 22
2 64038 1 22
2 64039 1 22
2 64040 1 22
2 64041 1 22
2 64042 1 22
2 64043 1 22
2 64044 1 22
2 64045 1 22
2 64046 1 22
2 64047 1 22
2 64048 1 22
2 64049 1 22
2 64050 1 22
2 64051 1 22
2 64052 1 22
2 64053 1 22
2 64054 1 22
2 64055 1 22
2 64056 1 22
2 64057 1 22
2 64058 1 22
2 64059 1 22
2 64060 1 22
2 64061 1 22
2 64062 1 22
2 64063 1 22
2 64064 1 22
2 64065 1 22
2 64066 1 22
2 64067 1 22
2 64068 1 22
2 64069 1 22
2 64070 1 22
2 64071 1 22
2 64072 1 22
2 64073 1 22
2 64074 1 22
2 64075 1 22
2 64076 1 22
2 64077 1 22
2 64078 1 22
2 64079 1 22
2 64080 1 22
2 64081 1 22
2 64082 1 22
2 64083 1 22
2 64084 1 22
2 64085 1 22
2 64086 1 22
2 64087 1 22
1 23 0 106 0
2 64088 1 23
2 64089 1 23
2 64090 1 23
2 64091 1 23
2 64092 1 23
2 64093 1 23
2 64094 1 23
2 64095 1 23
2 64096 1 23
2 64097 1 23
2 64098 1 23
2 64099 1 23
2 64100 1 23
2 64101 1 23
2 64102 1 23
2 64103 1 23
2 64104 1 23
2 64105 1 23
2 64106 1 23
2 64107 1 23
2 64108 1 23
2 64109 1 23
2 64110 1 23
2 64111 1 23
2 64112 1 23
2 64113 1 23
2 64114 1 23
2 64115 1 23
2 64116 1 23
2 64117 1 23
2 64118 1 23
2 64119 1 23
2 64120 1 23
2 64121 1 23
2 64122 1 23
2 64123 1 23
2 64124 1 23
2 64125 1 23
2 64126 1 23
2 64127 1 23
2 64128 1 23
2 64129 1 23
2 64130 1 23
2 64131 1 23
2 64132 1 23
2 64133 1 23
2 64134 1 23
2 64135 1 23
2 64136 1 23
2 64137 1 23
2 64138 1 23
2 64139 1 23
2 64140 1 23
2 64141 1 23
2 64142 1 23
2 64143 1 23
2 64144 1 23
2 64145 1 23
2 64146 1 23
2 64147 1 23
2 64148 1 23
2 64149 1 23
2 64150 1 23
2 64151 1 23
2 64152 1 23
2 64153 1 23
2 64154 1 23
2 64155 1 23
2 64156 1 23
2 64157 1 23
2 64158 1 23
2 64159 1 23
2 64160 1 23
2 64161 1 23
2 64162 1 23
2 64163 1 23
2 64164 1 23
2 64165 1 23
2 64166 1 23
2 64167 1 23
2 64168 1 23
2 64169 1 23
2 64170 1 23
2 64171 1 23
2 64172 1 23
2 64173 1 23
2 64174 1 23
2 64175 1 23
2 64176 1 23
2 64177 1 23
2 64178 1 23
2 64179 1 23
2 64180 1 23
2 64181 1 23
2 64182 1 23
2 64183 1 23
2 64184 1 23
2 64185 1 23
2 64186 1 23
2 64187 1 23
2 64188 1 23
2 64189 1 23
2 64190 1 23
2 64191 1 23
2 64192 1 23
2 64193 1 23
1 24 0 3 0
2 64194 1 24
2 64195 1 24
2 64196 1 24
2 64197 1 27
2 64198 1 27
2 64199 1 27
2 64200 1 27
2 64201 1 27
2 64202 1 27
2 64203 1 27
2 64204 1 27
2 64205 1 27
2 64206 1 27
2 64207 1 27
2 64208 1 27
2 64209 1 27
2 64210 1 27
2 64211 1 27
2 64212 1 27
2 64213 1 27
2 64214 1 27
2 64215 1 27
2 64216 1 27
2 64217 1 27
2 64218 1 27
2 64219 1 27
2 64220 1 27
2 64221 1 27
2 64222 1 27
2 64223 1 27
2 64224 1 27
2 64225 1 27
2 64226 1 27
2 64227 1 27
2 64228 1 27
2 64229 1 27
2 64230 1 27
2 64231 1 27
2 64232 1 27
2 64233 1 27
2 64234 1 27
2 64235 1 27
2 64236 1 27
2 64237 1 27
2 64238 1 27
2 64239 1 27
2 64240 1 27
2 64241 1 27
2 64242 1 27
2 64243 1 27
2 64244 1 27
2 64245 1 27
2 64246 1 27
2 64247 1 27
2 64248 1 27
2 64249 1 27
2 64250 1 27
2 64251 1 27
2 64252 1 27
2 64253 1 27
2 64254 1 27
2 64255 1 27
2 64256 1 27
2 64257 1 27
2 64258 1 27
2 64259 1 27
2 64260 1 27
2 64261 1 27
2 64262 1 27
2 64263 1 27
2 64264 1 27
2 64265 1 27
2 64266 1 27
2 64267 1 27
2 64268 1 27
2 64269 1 27
2 64270 1 27
2 64271 1 27
2 64272 1 27
2 64273 1 27
2 64274 1 27
2 64275 1 27
2 64276 1 27
2 64277 1 27
2 64278 1 27
2 64279 1 27
2 64280 1 27
2 64281 1 27
2 64282 1 27
2 64283 1 27
2 64284 1 27
2 64285 1 27
2 64286 1 27
2 64287 1 27
2 64288 1 27
2 64289 1 27
2 64290 1 27
2 64291 1 27
2 64292 1 27
2 64293 1 27
2 64294 1 27
2 64295 1 27
2 64296 1 27
2 64297 1 27
2 64298 1 27
2 64299 1 27
2 64300 1 27
2 64301 1 27
2 64302 1 27
2 64303 1 27
2 64304 1 27
2 64305 1 27
2 64306 1 27
2 64307 1 27
2 64308 1 27
2 64309 1 27
2 64310 1 27
2 64311 1 27
2 64312 1 27
2 64313 1 27
2 64314 1 27
2 64315 1 27
2 64316 1 27
2 64317 1 27
2 64318 1 27
2 64319 1 27
2 64320 1 27
2 64321 1 27
2 64322 1 27
2 64323 1 27
2 64324 1 27
2 64325 1 27
2 64326 1 27
2 64327 1 27
2 64328 1 27
2 64329 1 27
2 64330 1 27
2 64331 1 27
2 64332 1 27
2 64333 1 27
2 64334 1 27
2 64335 1 27
2 64336 1 27
2 64337 1 27
2 64338 1 27
2 64339 1 27
2 64340 1 27
2 64341 1 27
2 64342 1 27
2 64343 1 27
2 64344 1 27
2 64345 1 27
2 64346 1 27
2 64347 1 27
2 64348 1 27
2 64349 1 27
2 64350 1 27
2 64351 1 27
2 64352 1 27
2 64353 1 27
2 64354 1 27
2 64355 1 27
2 64356 1 27
2 64357 1 27
2 64358 1 27
2 64359 1 27
2 64360 1 27
2 64361 1 27
2 64362 1 27
2 64363 1 27
2 64364 1 27
2 64365 1 27
2 64366 1 27
2 64367 1 27
2 64368 1 27
2 64369 1 27
2 64370 1 27
2 64371 1 27
2 64372 1 27
2 64373 1 27
2 64374 1 28
2 64375 1 28
2 64376 1 28
2 64377 1 28
2 64378 1 28
2 64379 1 28
2 64380 1 28
2 64381 1 28
2 64382 1 28
2 64383 1 28
2 64384 1 28
2 64385 1 28
2 64386 1 28
2 64387 1 28
2 64388 1 28
2 64389 1 28
2 64390 1 28
2 64391 1 28
2 64392 1 28
2 64393 1 28
2 64394 1 28
2 64395 1 28
2 64396 1 28
2 64397 1 28
2 64398 1 28
2 64399 1 28
2 64400 1 28
2 64401 1 28
2 64402 1 28
2 64403 1 28
2 64404 1 28
2 64405 1 28
2 64406 1 28
2 64407 1 28
2 64408 1 28
2 64409 1 28
2 64410 1 28
2 64411 1 28
2 64412 1 28
2 64413 1 28
2 64414 1 28
2 64415 1 28
2 64416 1 28
2 64417 1 28
2 64418 1 28
2 64419 1 28
2 64420 1 28
2 64421 1 28
2 64422 1 28
2 64423 1 28
2 64424 1 28
2 64425 1 28
2 64426 1 28
2 64427 1 28
2 64428 1 28
2 64429 1 28
2 64430 1 28
2 64431 1 28
2 64432 1 28
2 64433 1 28
2 64434 1 28
2 64435 1 28
2 64436 1 28
2 64437 1 28
2 64438 1 28
2 64439 1 28
2 64440 1 28
2 64441 1 28
2 64442 1 28
2 64443 1 28
2 64444 1 28
2 64445 1 28
2 64446 1 28
2 64447 1 28
2 64448 1 28
2 64449 1 28
2 64450 1 28
2 64451 1 28
2 64452 1 28
2 64453 1 28
2 64454 1 28
2 64455 1 28
2 64456 1 28
2 64457 1 28
2 64458 1 28
2 64459 1 28
2 64460 1 28
2 64461 1 28
2 64462 1 28
2 64463 1 28
2 64464 1 28
2 64465 1 28
2 64466 1 28
2 64467 1 28
2 64468 1 28
2 64469 1 28
2 64470 1 28
2 64471 1 28
2 64472 1 28
2 64473 1 28
2 64474 1 28
2 64475 1 28
2 64476 1 28
2 64477 1 28
2 64478 1 28
2 64479 1 28
2 64480 1 28
2 64481 1 28
2 64482 1 28
2 64483 1 28
2 64484 1 28
2 64485 1 28
2 64486 1 28
2 64487 1 28
2 64488 1 28
2 64489 1 28
2 64490 1 28
2 64491 1 28
2 64492 1 28
2 64493 1 28
2 64494 1 28
2 64495 1 28
2 64496 1 28
2 64497 1 28
2 64498 1 28
2 64499 1 28
2 64500 1 28
2 64501 1 28
2 64502 1 28
2 64503 1 28
2 64504 1 28
2 64505 1 28
2 64506 1 28
2 64507 1 28
2 64508 1 28
2 64509 1 28
2 64510 1 28
2 64511 1 28
2 64512 1 28
2 64513 1 28
2 64514 1 28
2 64515 1 28
2 64516 1 28
2 64517 1 28
2 64518 1 28
2 64519 1 28
2 64520 1 28
2 64521 1 28
2 64522 1 28
2 64523 1 28
2 64524 1 28
2 64525 1 28
2 64526 1 28
2 64527 1 28
2 64528 1 28
2 64529 1 28
2 64530 1 28
2 64531 1 28
2 64532 1 28
2 64533 1 28
2 64534 1 28
2 64535 1 28
2 64536 1 28
2 64537 1 28
2 64538 1 28
2 64539 1 28
2 64540 1 28
2 64541 1 28
2 64542 1 28
2 64543 1 28
2 64544 1 28
2 64545 1 28
2 64546 1 28
2 64547 1 28
2 64548 1 28
2 64549 1 28
2 64550 1 28
2 64551 1 28
2 64552 1 28
2 64553 1 28
2 64554 1 28
2 64555 1 28
2 64556 1 28
2 64557 1 28
2 64558 1 28
2 64559 1 28
2 64560 1 28
2 64561 1 28
2 64562 1 28
2 64563 1 28
2 64564 1 28
2 64565 1 28
2 64566 1 28
2 64567 1 28
2 64568 1 28
2 64569 1 28
2 64570 1 28
2 64571 1 28
2 64572 1 28
2 64573 1 28
2 64574 1 28
2 64575 1 28
2 64576 1 28
2 64577 1 28
2 64578 1 28
2 64579 1 28
2 64580 1 28
2 64581 1 28
2 64582 1 28
2 64583 1 28
2 64584 1 28
2 64585 1 28
2 64586 1 28
2 64587 1 28
2 64588 1 28
2 64589 1 28
2 64590 1 28
2 64591 1 28
2 64592 1 28
2 64593 1 28
2 64594 1 28
2 64595 1 28
2 64596 1 28
2 64597 1 28
2 64598 1 28
2 64599 1 28
2 64600 1 28
2 64601 1 28
2 64602 1 28
2 64603 1 29
2 64604 1 29
2 64605 1 29
2 64606 1 29
2 64607 1 29
2 64608 1 29
2 64609 1 29
2 64610 1 29
2 64611 1 29
2 64612 1 29
2 64613 1 29
2 64614 1 29
2 64615 1 29
2 64616 1 29
2 64617 1 29
2 64618 1 29
2 64619 1 29
2 64620 1 29
2 64621 1 29
2 64622 1 29
2 64623 1 29
2 64624 1 29
2 64625 1 29
2 64626 1 29
2 64627 1 29
2 64628 1 29
2 64629 1 29
2 64630 1 29
2 64631 1 29
2 64632 1 29
2 64633 1 29
2 64634 1 29
2 64635 1 29
2 64636 1 29
2 64637 1 29
2 64638 1 29
2 64639 1 29
2 64640 1 29
2 64641 1 29
2 64642 1 29
2 64643 1 29
2 64644 1 29
2 64645 1 29
2 64646 1 29
2 64647 1 29
2 64648 1 29
2 64649 1 29
2 64650 1 29
2 64651 1 29
2 64652 1 29
2 64653 1 29
2 64654 1 29
2 64655 1 29
2 64656 1 29
2 64657 1 29
2 64658 1 29
2 64659 1 29
2 64660 1 29
2 64661 1 29
2 64662 1 29
2 64663 1 29
2 64664 1 29
2 64665 1 29
2 64666 1 29
2 64667 1 29
2 64668 1 29
2 64669 1 29
2 64670 1 29
2 64671 1 29
2 64672 1 29
2 64673 1 29
2 64674 1 29
2 64675 1 29
2 64676 1 29
2 64677 1 29
2 64678 1 29
2 64679 1 29
2 64680 1 29
2 64681 1 29
2 64682 1 29
2 64683 1 29
2 64684 1 29
2 64685 1 29
2 64686 1 29
2 64687 1 29
2 64688 1 29
2 64689 1 29
2 64690 1 29
2 64691 1 29
2 64692 1 29
2 64693 1 29
2 64694 1 29
2 64695 1 29
2 64696 1 29
2 64697 1 29
2 64698 1 29
2 64699 1 29
2 64700 1 29
2 64701 1 29
2 64702 1 29
2 64703 1 29
2 64704 1 29
2 64705 1 29
2 64706 1 29
2 64707 1 29
2 64708 1 29
2 64709 1 29
2 64710 1 29
2 64711 1 29
2 64712 1 29
2 64713 1 29
2 64714 1 29
2 64715 1 29
2 64716 1 29
2 64717 1 29
2 64718 1 29
2 64719 1 29
2 64720 1 29
2 64721 1 29
2 64722 1 29
2 64723 1 29
2 64724 1 29
2 64725 1 29
2 64726 1 29
2 64727 1 29
2 64728 1 29
2 64729 1 29
2 64730 1 29
2 64731 1 29
2 64732 1 29
2 64733 1 29
2 64734 1 29
2 64735 1 29
2 64736 1 29
2 64737 1 29
2 64738 1 29
2 64739 1 29
2 64740 1 29
2 64741 1 29
2 64742 1 29
2 64743 1 29
2 64744 1 29
2 64745 1 29
2 64746 1 29
2 64747 1 29
2 64748 1 29
2 64749 1 29
2 64750 1 29
2 64751 1 29
2 64752 1 29
2 64753 1 29
2 64754 1 29
2 64755 1 29
2 64756 1 29
2 64757 1 29
2 64758 1 29
2 64759 1 29
2 64760 1 29
2 64761 1 29
2 64762 1 29
2 64763 1 29
2 64764 1 29
2 64765 1 29
2 64766 1 29
2 64767 1 29
2 64768 1 29
2 64769 1 29
2 64770 1 29
2 64771 1 29
2 64772 1 29
2 64773 1 29
2 64774 1 29
2 64775 1 29
2 64776 1 29
2 64777 1 29
2 64778 1 29
2 64779 1 29
2 64780 1 29
2 64781 1 29
2 64782 1 29
2 64783 1 29
2 64784 1 29
2 64785 1 29
2 64786 1 29
2 64787 1 29
2 64788 1 29
2 64789 1 29
2 64790 1 29
2 64791 1 29
2 64792 1 29
2 64793 1 29
2 64794 1 29
2 64795 1 29
2 64796 1 29
2 64797 1 29
2 64798 1 29
2 64799 1 29
2 64800 1 29
2 64801 1 29
2 64802 1 29
2 64803 1 29
2 64804 1 29
2 64805 1 29
2 64806 1 29
2 64807 1 29
2 64808 1 29
2 64809 1 29
2 64810 1 29
2 64811 1 29
2 64812 1 29
2 64813 1 29
2 64814 1 29
2 64815 1 29
2 64816 1 29
2 64817 1 29
2 64818 1 29
2 64819 1 29
2 64820 1 29
2 64821 1 29
2 64822 1 29
2 64823 1 29
2 64824 1 29
2 64825 1 29
2 64826 1 29
2 64827 1 29
2 64828 1 29
2 64829 1 29
2 64830 1 29
2 64831 1 30
2 64832 1 30
2 64833 1 30
2 64834 1 30
2 64835 1 30
2 64836 1 30
2 64837 1 30
2 64838 1 30
2 64839 1 30
2 64840 1 30
2 64841 1 30
2 64842 1 30
2 64843 1 30
2 64844 1 30
2 64845 1 30
2 64846 1 30
2 64847 1 30
2 64848 1 30
2 64849 1 30
2 64850 1 30
2 64851 1 30
2 64852 1 30
2 64853 1 30
2 64854 1 30
2 64855 1 30
2 64856 1 30
2 64857 1 30
2 64858 1 30
2 64859 1 30
2 64860 1 30
2 64861 1 30
2 64862 1 30
2 64863 1 30
2 64864 1 30
2 64865 1 30
2 64866 1 30
2 64867 1 30
2 64868 1 30
2 64869 1 30
2 64870 1 30
2 64871 1 30
2 64872 1 30
2 64873 1 30
2 64874 1 30
2 64875 1 30
2 64876 1 30
2 64877 1 30
2 64878 1 30
2 64879 1 30
2 64880 1 30
2 64881 1 30
2 64882 1 30
2 64883 1 30
2 64884 1 30
2 64885 1 30
2 64886 1 30
2 64887 1 30
2 64888 1 30
2 64889 1 30
2 64890 1 30
2 64891 1 30
2 64892 1 30
2 64893 1 30
2 64894 1 30
2 64895 1 30
2 64896 1 30
2 64897 1 30
2 64898 1 30
2 64899 1 30
2 64900 1 30
2 64901 1 30
2 64902 1 30
2 64903 1 30
2 64904 1 30
2 64905 1 30
2 64906 1 30
2 64907 1 30
2 64908 1 30
2 64909 1 30
2 64910 1 30
2 64911 1 30
2 64912 1 30
2 64913 1 30
2 64914 1 30
2 64915 1 30
2 64916 1 30
2 64917 1 30
2 64918 1 30
2 64919 1 30
2 64920 1 30
2 64921 1 30
2 64922 1 30
2 64923 1 30
2 64924 1 30
2 64925 1 30
2 64926 1 30
2 64927 1 30
2 64928 1 30
2 64929 1 30
2 64930 1 30
2 64931 1 30
2 64932 1 30
2 64933 1 30
2 64934 1 30
2 64935 1 30
2 64936 1 30
2 64937 1 30
2 64938 1 30
2 64939 1 30
2 64940 1 30
2 64941 1 30
2 64942 1 30
2 64943 1 30
2 64944 1 30
2 64945 1 30
2 64946 1 30
2 64947 1 30
2 64948 1 30
2 64949 1 30
2 64950 1 30
2 64951 1 30
2 64952 1 30
2 64953 1 30
2 64954 1 30
2 64955 1 30
2 64956 1 30
2 64957 1 30
2 64958 1 30
2 64959 1 30
2 64960 1 30
2 64961 1 30
2 64962 1 30
2 64963 1 30
2 64964 1 30
2 64965 1 30
2 64966 1 30
2 64967 1 30
2 64968 1 30
2 64969 1 30
2 64970 1 30
2 64971 1 30
2 64972 1 30
2 64973 1 30
2 64974 1 30
2 64975 1 30
2 64976 1 30
2 64977 1 30
2 64978 1 30
2 64979 1 30
2 64980 1 30
2 64981 1 30
2 64982 1 30
2 64983 1 30
2 64984 1 30
2 64985 1 30
2 64986 1 30
2 64987 1 30
2 64988 1 30
2 64989 1 30
2 64990 1 30
2 64991 1 30
2 64992 1 30
2 64993 1 30
2 64994 1 30
2 64995 1 30
2 64996 1 30
2 64997 1 30
2 64998 1 30
2 64999 1 30
2 65000 1 30
2 65001 1 30
2 65002 1 30
2 65003 1 30
2 65004 1 30
2 65005 1 30
2 65006 1 30
2 65007 1 30
2 65008 1 30
2 65009 1 30
2 65010 1 30
2 65011 1 30
2 65012 1 30
2 65013 1 30
2 65014 1 30
2 65015 1 30
2 65016 1 30
2 65017 1 30
2 65018 1 30
2 65019 1 30
2 65020 1 30
2 65021 1 30
2 65022 1 30
2 65023 1 30
2 65024 1 30
2 65025 1 30
2 65026 1 30
2 65027 1 30
2 65028 1 30
2 65029 1 30
2 65030 1 30
2 65031 1 30
2 65032 1 30
2 65033 1 30
2 65034 1 30
2 65035 1 30
2 65036 1 30
2 65037 1 30
2 65038 1 30
2 65039 1 30
2 65040 1 30
2 65041 1 30
2 65042 1 31
2 65043 1 31
2 65044 1 31
2 65045 1 31
2 65046 1 31
2 65047 1 31
2 65048 1 31
2 65049 1 31
2 65050 1 31
2 65051 1 31
2 65052 1 31
2 65053 1 31
2 65054 1 31
2 65055 1 31
2 65056 1 31
2 65057 1 31
2 65058 1 31
2 65059 1 31
2 65060 1 31
2 65061 1 31
2 65062 1 31
2 65063 1 31
2 65064 1 31
2 65065 1 31
2 65066 1 31
2 65067 1 31
2 65068 1 31
2 65069 1 31
2 65070 1 31
2 65071 1 31
2 65072 1 31
2 65073 1 31
2 65074 1 31
2 65075 1 31
2 65076 1 31
2 65077 1 31
2 65078 1 31
2 65079 1 31
2 65080 1 31
2 65081 1 31
2 65082 1 31
2 65083 1 31
2 65084 1 31
2 65085 1 31
2 65086 1 31
2 65087 1 31
2 65088 1 31
2 65089 1 31
2 65090 1 31
2 65091 1 31
2 65092 1 31
2 65093 1 31
2 65094 1 31
2 65095 1 31
2 65096 1 31
2 65097 1 31
2 65098 1 31
2 65099 1 31
2 65100 1 31
2 65101 1 31
2 65102 1 31
2 65103 1 31
2 65104 1 31
2 65105 1 31
2 65106 1 31
2 65107 1 31
2 65108 1 31
2 65109 1 31
2 65110 1 31
2 65111 1 31
2 65112 1 31
2 65113 1 31
2 65114 1 31
2 65115 1 31
2 65116 1 31
2 65117 1 31
2 65118 1 31
2 65119 1 31
2 65120 1 31
2 65121 1 31
2 65122 1 31
2 65123 1 31
2 65124 1 31
2 65125 1 31
2 65126 1 31
2 65127 1 31
2 65128 1 31
2 65129 1 31
2 65130 1 31
2 65131 1 31
2 65132 1 31
2 65133 1 31
2 65134 1 31
2 65135 1 31
2 65136 1 31
2 65137 1 31
2 65138 1 31
2 65139 1 31
2 65140 1 31
2 65141 1 31
2 65142 1 31
2 65143 1 31
2 65144 1 31
2 65145 1 31
2 65146 1 31
2 65147 1 31
2 65148 1 31
2 65149 1 31
2 65150 1 31
2 65151 1 31
2 65152 1 31
2 65153 1 31
2 65154 1 31
2 65155 1 31
2 65156 1 31
2 65157 1 31
2 65158 1 31
2 65159 1 31
2 65160 1 31
2 65161 1 31
2 65162 1 31
2 65163 1 31
2 65164 1 31
2 65165 1 31
2 65166 1 31
2 65167 1 31
2 65168 1 31
2 65169 1 31
2 65170 1 31
2 65171 1 31
2 65172 1 31
2 65173 1 31
2 65174 1 31
2 65175 1 31
2 65176 1 31
2 65177 1 31
2 65178 1 31
2 65179 1 31
2 65180 1 31
2 65181 1 31
2 65182 1 31
2 65183 1 31
2 65184 1 31
2 65185 1 31
2 65186 1 31
2 65187 1 31
2 65188 1 31
2 65189 1 31
2 65190 1 31
2 65191 1 31
2 65192 1 31
2 65193 1 31
2 65194 1 31
2 65195 1 31
2 65196 1 31
2 65197 1 31
2 65198 1 31
2 65199 1 31
2 65200 1 31
2 65201 1 31
2 65202 1 31
2 65203 1 31
2 65204 1 31
2 65205 1 31
2 65206 1 31
2 65207 1 31
2 65208 1 31
2 65209 1 31
2 65210 1 31
2 65211 1 31
2 65212 1 31
2 65213 1 31
2 65214 1 31
2 65215 1 31
2 65216 1 31
2 65217 1 31
2 65218 1 31
2 65219 1 31
2 65220 1 31
2 65221 1 31
2 65222 1 31
2 65223 1 31
2 65224 1 31
2 65225 1 31
2 65226 1 31
2 65227 1 31
2 65228 1 31
2 65229 1 31
2 65230 1 31
2 65231 1 31
2 65232 1 31
2 65233 1 31
2 65234 1 31
2 65235 1 31
2 65236 1 31
2 65237 1 31
2 65238 1 31
2 65239 1 31
2 65240 1 31
2 65241 1 31
2 65242 1 31
2 65243 1 31
2 65244 1 31
2 65245 1 31
2 65246 1 31
2 65247 1 31
2 65248 1 31
2 65249 1 31
2 65250 1 31
2 65251 1 31
2 65252 1 31
2 65253 1 31
2 65254 1 31
2 65255 1 31
2 65256 1 31
2 65257 1 31
2 65258 1 31
2 65259 1 31
2 65260 1 31
2 65261 1 31
2 65262 1 31
2 65263 1 31
2 65264 1 31
2 65265 1 31
2 65266 1 31
2 65267 1 31
2 65268 1 31
2 65269 1 31
2 65270 1 31
2 65271 1 31
2 65272 1 31
2 65273 1 31
2 65274 1 31
2 65275 1 31
2 65276 1 31
2 65277 1 31
2 65278 1 31
2 65279 1 31
2 65280 1 31
2 65281 1 31
2 65282 1 31
2 65283 1 31
2 65284 1 31
2 65285 1 31
2 65286 1 31
2 65287 1 31
2 65288 1 31
2 65289 1 31
2 65290 1 31
2 65291 1 31
2 65292 1 31
2 65293 1 31
2 65294 1 31
2 65295 1 31
2 65296 1 31
2 65297 1 31
2 65298 1 31
2 65299 1 31
2 65300 1 31
2 65301 1 31
2 65302 1 31
2 65303 1 31
2 65304 1 31
2 65305 1 31
2 65306 1 31
2 65307 1 31
2 65308 1 31
2 65309 1 31
2 65310 1 31
2 65311 1 31
2 65312 1 32
2 65313 1 32
2 65314 1 32
2 65315 1 32
2 65316 1 32
2 65317 1 32
2 65318 1 32
2 65319 1 32
2 65320 1 32
2 65321 1 32
2 65322 1 32
2 65323 1 32
2 65324 1 32
2 65325 1 32
2 65326 1 32
2 65327 1 32
2 65328 1 32
2 65329 1 32
2 65330 1 32
2 65331 1 32
2 65332 1 32
2 65333 1 32
2 65334 1 32
2 65335 1 32
2 65336 1 32
2 65337 1 32
2 65338 1 32
2 65339 1 32
2 65340 1 32
2 65341 1 32
2 65342 1 32
2 65343 1 32
2 65344 1 32
2 65345 1 32
2 65346 1 32
2 65347 1 32
2 65348 1 32
2 65349 1 32
2 65350 1 32
2 65351 1 32
2 65352 1 32
2 65353 1 32
2 65354 1 32
2 65355 1 32
2 65356 1 32
2 65357 1 32
2 65358 1 32
2 65359 1 32
2 65360 1 32
2 65361 1 32
2 65362 1 32
2 65363 1 32
2 65364 1 32
2 65365 1 32
2 65366 1 32
2 65367 1 32
2 65368 1 32
2 65369 1 32
2 65370 1 32
2 65371 1 32
2 65372 1 32
2 65373 1 32
2 65374 1 32
2 65375 1 32
2 65376 1 32
2 65377 1 32
2 65378 1 32
2 65379 1 32
2 65380 1 32
2 65381 1 32
2 65382 1 32
2 65383 1 32
2 65384 1 32
2 65385 1 32
2 65386 1 32
2 65387 1 32
2 65388 1 32
2 65389 1 32
2 65390 1 32
2 65391 1 32
2 65392 1 32
2 65393 1 32
2 65394 1 32
2 65395 1 32
2 65396 1 32
2 65397 1 32
2 65398 1 32
2 65399 1 32
2 65400 1 32
2 65401 1 32
2 65402 1 32
2 65403 1 32
2 65404 1 32
2 65405 1 32
2 65406 1 32
2 65407 1 32
2 65408 1 32
2 65409 1 32
2 65410 1 32
2 65411 1 32
2 65412 1 32
2 65413 1 32
2 65414 1 32
2 65415 1 32
2 65416 1 32
2 65417 1 32
2 65418 1 32
2 65419 1 32
2 65420 1 32
2 65421 1 32
2 65422 1 32
2 65423 1 32
2 65424 1 32
2 65425 1 32
2 65426 1 32
2 65427 1 32
2 65428 1 32
2 65429 1 32
2 65430 1 32
2 65431 1 32
2 65432 1 32
2 65433 1 32
2 65434 1 32
2 65435 1 32
2 65436 1 32
2 65437 1 32
2 65438 1 32
2 65439 1 32
2 65440 1 32
2 65441 1 32
2 65442 1 32
2 65443 1 32
2 65444 1 32
2 65445 1 32
2 65446 1 32
2 65447 1 32
2 65448 1 32
2 65449 1 32
2 65450 1 32
2 65451 1 32
2 65452 1 32
2 65453 1 32
2 65454 1 32
2 65455 1 32
2 65456 1 32
2 65457 1 32
2 65458 1 32
2 65459 1 32
2 65460 1 32
2 65461 1 32
2 65462 1 32
2 65463 1 32
2 65464 1 32
2 65465 1 32
2 65466 1 32
2 65467 1 32
2 65468 1 32
2 65469 1 32
2 65470 1 32
2 65471 1 32
2 65472 1 32
2 65473 1 32
2 65474 1 32
2 65475 1 32
2 65476 1 32
2 65477 1 32
2 65478 1 32
2 65479 1 32
2 65480 1 32
2 65481 1 32
2 65482 1 32
2 65483 1 32
2 65484 1 32
2 65485 1 32
2 65486 1 32
2 65487 1 32
2 65488 1 32
2 65489 1 32
2 65490 1 32
2 65491 1 32
2 65492 1 32
2 65493 1 32
2 65494 1 32
2 65495 1 32
2 65496 1 32
2 65497 1 32
2 65498 1 32
2 65499 1 32
2 65500 1 32
2 65501 1 32
2 65502 1 32
2 65503 1 32
2 65504 1 32
2 65505 1 32
2 65506 1 32
2 65507 1 32
2 65508 1 32
2 65509 1 32
2 65510 1 32
2 65511 1 32
2 65512 1 32
2 65513 1 32
2 65514 1 32
2 65515 1 32
2 65516 1 32
2 65517 1 32
2 65518 1 32
2 65519 1 32
2 65520 1 32
2 65521 1 32
2 65522 1 32
2 65523 1 32
2 65524 1 32
2 65525 1 32
2 65526 1 32
2 65527 1 32
2 65528 1 32
2 65529 1 32
2 65530 1 32
2 65531 1 32
2 65532 1 32
2 65533 1 32
2 65534 1 32
2 65535 1 32
2 65536 1 32
2 65537 1 33
2 65538 1 33
2 65539 1 33
2 65540 1 33
2 65541 1 33
2 65542 1 33
2 65543 1 33
2 65544 1 33
2 65545 1 33
2 65546 1 33
2 65547 1 33
2 65548 1 33
2 65549 1 33
2 65550 1 33
2 65551 1 33
2 65552 1 33
2 65553 1 33
2 65554 1 33
2 65555 1 33
2 65556 1 33
2 65557 1 33
2 65558 1 33
2 65559 1 33
2 65560 1 33
2 65561 1 33
2 65562 1 33
2 65563 1 33
2 65564 1 33
2 65565 1 33
2 65566 1 33
2 65567 1 33
2 65568 1 33
2 65569 1 33
2 65570 1 33
2 65571 1 33
2 65572 1 33
2 65573 1 33
2 65574 1 33
2 65575 1 33
2 65576 1 33
2 65577 1 33
2 65578 1 33
2 65579 1 33
2 65580 1 33
2 65581 1 33
2 65582 1 33
2 65583 1 33
2 65584 1 33
2 65585 1 33
2 65586 1 33
2 65587 1 33
2 65588 1 33
2 65589 1 33
2 65590 1 33
2 65591 1 33
2 65592 1 33
2 65593 1 33
2 65594 1 33
2 65595 1 33
2 65596 1 33
2 65597 1 33
2 65598 1 33
2 65599 1 33
2 65600 1 33
2 65601 1 33
2 65602 1 33
2 65603 1 33
2 65604 1 33
2 65605 1 33
2 65606 1 33
2 65607 1 33
2 65608 1 33
2 65609 1 33
2 65610 1 33
2 65611 1 33
2 65612 1 33
2 65613 1 33
2 65614 1 33
2 65615 1 33
2 65616 1 33
2 65617 1 33
2 65618 1 33
2 65619 1 33
2 65620 1 33
2 65621 1 33
2 65622 1 33
2 65623 1 33
2 65624 1 33
2 65625 1 33
2 65626 1 33
2 65627 1 33
2 65628 1 33
2 65629 1 33
2 65630 1 33
2 65631 1 33
2 65632 1 33
2 65633 1 33
2 65634 1 33
2 65635 1 33
2 65636 1 33
2 65637 1 33
2 65638 1 33
2 65639 1 33
2 65640 1 33
2 65641 1 33
2 65642 1 33
2 65643 1 33
2 65644 1 33
2 65645 1 33
2 65646 1 33
2 65647 1 33
2 65648 1 33
2 65649 1 33
2 65650 1 33
2 65651 1 33
2 65652 1 33
2 65653 1 33
2 65654 1 33
2 65655 1 33
2 65656 1 33
2 65657 1 33
2 65658 1 33
2 65659 1 33
2 65660 1 33
2 65661 1 33
2 65662 1 33
2 65663 1 33
2 65664 1 34
2 65665 1 34
2 65666 1 34
2 65667 1 34
2 65668 1 34
2 65669 1 34
2 65670 1 34
2 65671 1 34
2 65672 1 35
2 65673 1 35
2 65674 1 35
2 65675 1 35
2 65676 1 35
2 65677 1 35
2 65678 1 35
2 65679 1 35
2 65680 1 35
2 65681 1 35
2 65682 1 35
2 65683 1 35
2 65684 1 35
2 65685 1 35
2 65686 1 35
2 65687 1 35
2 65688 1 35
2 65689 1 35
2 65690 1 35
2 65691 1 35
2 65692 1 35
2 65693 1 35
2 65694 1 35
2 65695 1 35
2 65696 1 35
2 65697 1 35
2 65698 1 35
2 65699 1 35
2 65700 1 35
2 65701 1 35
2 65702 1 35
2 65703 1 35
2 65704 1 35
2 65705 1 35
2 65706 1 35
2 65707 1 35
2 65708 1 35
2 65709 1 35
2 65710 1 35
2 65711 1 35
2 65712 1 35
2 65713 1 35
2 65714 1 35
2 65715 1 35
2 65716 1 35
2 65717 1 35
2 65718 1 35
2 65719 1 35
2 65720 1 35
2 65721 1 35
2 65722 1 35
2 65723 1 35
2 65724 1 35
2 65725 1 35
2 65726 1 35
2 65727 1 35
2 65728 1 35
2 65729 1 35
2 65730 1 35
2 65731 1 35
2 65732 1 35
2 65733 1 35
2 65734 1 35
2 65735 1 35
2 65736 1 35
2 65737 1 35
2 65738 1 35
2 65739 1 35
2 65740 1 35
2 65741 1 35
2 65742 1 35
2 65743 1 35
2 65744 1 35
2 65745 1 35
2 65746 1 35
2 65747 1 35
2 65748 1 35
2 65749 1 35
2 65750 1 35
2 65751 1 36
2 65752 1 36
2 65753 1 36
2 65754 1 36
2 65755 1 36
2 65756 1 36
2 65757 1 36
2 65758 1 36
2 65759 1 36
2 65760 1 36
2 65761 1 36
2 65762 1 36
2 65763 1 36
2 65764 1 36
2 65765 1 36
2 65766 1 36
2 65767 1 36
2 65768 1 36
2 65769 1 36
2 65770 1 36
2 65771 1 36
2 65772 1 36
2 65773 1 36
2 65774 1 36
2 65775 1 36
2 65776 1 36
2 65777 1 36
2 65778 1 36
2 65779 1 36
2 65780 1 36
2 65781 1 36
2 65782 1 36
2 65783 1 36
2 65784 1 36
2 65785 1 36
2 65786 1 36
2 65787 1 36
2 65788 1 36
2 65789 1 36
2 65790 1 36
2 65791 1 36
2 65792 1 36
2 65793 1 36
2 65794 1 36
2 65795 1 36
2 65796 1 36
2 65797 1 36
2 65798 1 36
2 65799 1 36
2 65800 1 36
2 65801 1 36
2 65802 1 36
2 65803 1 36
2 65804 1 36
2 65805 1 36
2 65806 1 36
2 65807 1 36
2 65808 1 36
2 65809 1 36
2 65810 1 36
2 65811 1 36
2 65812 1 36
2 65813 1 36
2 65814 1 36
2 65815 1 36
2 65816 1 36
2 65817 1 36
2 65818 1 36
2 65819 1 36
2 65820 1 36
2 65821 1 36
2 65822 1 36
2 65823 1 36
2 65824 1 36
2 65825 1 36
2 65826 1 36
2 65827 1 36
2 65828 1 36
2 65829 1 36
2 65830 1 36
2 65831 1 36
2 65832 1 36
2 65833 1 36
2 65834 1 36
2 65835 1 36
2 65836 1 36
2 65837 1 36
2 65838 1 36
2 65839 1 36
2 65840 1 36
2 65841 1 36
2 65842 1 36
2 65843 1 36
2 65844 1 36
2 65845 1 36
2 65846 1 36
2 65847 1 36
2 65848 1 36
2 65849 1 36
2 65850 1 36
2 65851 1 36
2 65852 1 36
2 65853 1 36
2 65854 1 36
2 65855 1 36
2 65856 1 36
2 65857 1 36
2 65858 1 36
2 65859 1 36
2 65860 1 36
2 65861 1 36
2 65862 1 36
2 65863 1 36
2 65864 1 36
2 65865 1 36
2 65866 1 36
2 65867 1 36
2 65868 1 36
2 65869 1 36
2 65870 1 36
2 65871 1 36
2 65872 1 36
2 65873 1 36
2 65874 1 36
2 65875 1 36
2 65876 1 36
2 65877 1 36
2 65878 1 36
2 65879 1 36
2 65880 1 36
2 65881 1 36
2 65882 1 36
2 65883 1 36
2 65884 1 36
2 65885 1 36
2 65886 1 36
2 65887 1 36
2 65888 1 36
2 65889 1 36
2 65890 1 36
2 65891 1 36
2 65892 1 36
2 65893 1 36
2 65894 1 36
2 65895 1 36
2 65896 1 36
2 65897 1 36
2 65898 1 36
2 65899 1 36
2 65900 1 36
2 65901 1 36
2 65902 1 36
2 65903 1 36
2 65904 1 36
2 65905 1 36
2 65906 1 36
2 65907 1 36
2 65908 1 36
2 65909 1 36
2 65910 1 36
2 65911 1 36
2 65912 1 36
2 65913 1 37
2 65914 1 37
2 65915 1 37
2 65916 1 37
2 65917 1 37
2 65918 1 37
2 65919 1 37
2 65920 1 37
2 65921 1 37
2 65922 1 37
2 65923 1 37
2 65924 1 37
2 65925 1 37
2 65926 1 37
2 65927 1 37
2 65928 1 37
2 65929 1 37
2 65930 1 37
2 65931 1 37
2 65932 1 37
2 65933 1 37
2 65934 1 37
2 65935 1 37
2 65936 1 37
2 65937 1 37
2 65938 1 37
2 65939 1 37
2 65940 1 37
2 65941 1 37
2 65942 1 37
2 65943 1 37
2 65944 1 37
2 65945 1 37
2 65946 1 37
2 65947 1 37
2 65948 1 37
2 65949 1 37
2 65950 1 37
2 65951 1 37
2 65952 1 37
2 65953 1 37
2 65954 1 37
2 65955 1 37
2 65956 1 37
2 65957 1 37
2 65958 1 37
2 65959 1 37
2 65960 1 37
2 65961 1 37
2 65962 1 37
2 65963 1 37
2 65964 1 37
2 65965 1 37
2 65966 1 37
2 65967 1 37
2 65968 1 37
2 65969 1 37
2 65970 1 37
2 65971 1 37
2 65972 1 37
2 65973 1 37
2 65974 1 37
2 65975 1 37
2 65976 1 37
2 65977 1 37
2 65978 1 37
2 65979 1 37
2 65980 1 37
2 65981 1 37
2 65982 1 37
2 65983 1 37
2 65984 1 37
2 65985 1 37
2 65986 1 37
2 65987 1 37
2 65988 1 37
2 65989 1 37
2 65990 1 37
2 65991 1 37
2 65992 1 37
2 65993 1 37
2 65994 1 37
2 65995 1 37
2 65996 1 37
2 65997 1 37
2 65998 1 37
2 65999 1 37
2 66000 1 37
2 66001 1 37
2 66002 1 37
2 66003 1 37
2 66004 1 37
2 66005 1 37
2 66006 1 37
2 66007 1 37
2 66008 1 37
2 66009 1 37
2 66010 1 37
2 66011 1 37
2 66012 1 37
2 66013 1 37
2 66014 1 37
2 66015 1 37
2 66016 1 37
2 66017 1 37
2 66018 1 37
2 66019 1 37
2 66020 1 37
2 66021 1 37
2 66022 1 37
2 66023 1 37
2 66024 1 37
2 66025 1 37
2 66026 1 37
2 66027 1 37
2 66028 1 37
2 66029 1 37
2 66030 1 37
2 66031 1 37
2 66032 1 37
2 66033 1 37
2 66034 1 37
2 66035 1 37
2 66036 1 37
2 66037 1 37
2 66038 1 37
2 66039 1 37
2 66040 1 37
2 66041 1 37
2 66042 1 37
2 66043 1 37
2 66044 1 37
2 66045 1 37
2 66046 1 37
2 66047 1 37
2 66048 1 37
2 66049 1 37
2 66050 1 37
2 66051 1 37
2 66052 1 37
2 66053 1 37
2 66054 1 37
2 66055 1 37
2 66056 1 37
2 66057 1 37
2 66058 1 37
2 66059 1 37
2 66060 1 37
2 66061 1 37
2 66062 1 37
2 66063 1 37
2 66064 1 37
2 66065 1 37
2 66066 1 37
2 66067 1 37
2 66068 1 37
2 66069 1 37
2 66070 1 37
2 66071 1 37
2 66072 1 37
2 66073 1 37
2 66074 1 37
2 66075 1 37
2 66076 1 37
2 66077 1 37
2 66078 1 37
2 66079 1 37
2 66080 1 37
2 66081 1 37
2 66082 1 37
2 66083 1 37
2 66084 1 37
2 66085 1 37
2 66086 1 37
2 66087 1 37
2 66088 1 37
2 66089 1 37
2 66090 1 38
2 66091 1 38
2 66092 1 38
2 66093 1 38
2 66094 1 38
2 66095 1 38
2 66096 1 38
2 66097 1 38
2 66098 1 38
2 66099 1 38
2 66100 1 38
2 66101 1 38
2 66102 1 38
2 66103 1 38
2 66104 1 38
2 66105 1 38
2 66106 1 38
2 66107 1 38
2 66108 1 38
2 66109 1 38
2 66110 1 38
2 66111 1 38
2 66112 1 38
2 66113 1 38
2 66114 1 38
2 66115 1 38
2 66116 1 38
2 66117 1 38
2 66118 1 38
2 66119 1 38
2 66120 1 38
2 66121 1 38
2 66122 1 38
2 66123 1 38
2 66124 1 38
2 66125 1 38
2 66126 1 38
2 66127 1 38
2 66128 1 38
2 66129 1 38
2 66130 1 38
2 66131 1 38
2 66132 1 38
2 66133 1 38
2 66134 1 38
2 66135 1 38
2 66136 1 38
2 66137 1 38
2 66138 1 38
2 66139 1 38
2 66140 1 38
2 66141 1 38
2 66142 1 38
2 66143 1 38
2 66144 1 38
2 66145 1 38
2 66146 1 38
2 66147 1 38
2 66148 1 38
2 66149 1 38
2 66150 1 38
2 66151 1 38
2 66152 1 38
2 66153 1 38
2 66154 1 38
2 66155 1 38
2 66156 1 38
2 66157 1 38
2 66158 1 38
2 66159 1 38
2 66160 1 38
2 66161 1 38
2 66162 1 38
2 66163 1 38
2 66164 1 38
2 66165 1 38
2 66166 1 38
2 66167 1 38
2 66168 1 38
2 66169 1 38
2 66170 1 38
2 66171 1 38
2 66172 1 38
2 66173 1 38
2 66174 1 38
2 66175 1 38
2 66176 1 38
2 66177 1 38
2 66178 1 38
2 66179 1 38
2 66180 1 38
2 66181 1 38
2 66182 1 38
2 66183 1 38
2 66184 1 38
2 66185 1 38
2 66186 1 38
2 66187 1 38
2 66188 1 38
2 66189 1 38
2 66190 1 38
2 66191 1 38
2 66192 1 38
2 66193 1 38
2 66194 1 38
2 66195 1 38
2 66196 1 38
2 66197 1 38
2 66198 1 38
2 66199 1 38
2 66200 1 38
2 66201 1 38
2 66202 1 38
2 66203 1 38
2 66204 1 38
2 66205 1 38
2 66206 1 38
2 66207 1 38
2 66208 1 38
2 66209 1 38
2 66210 1 38
2 66211 1 38
2 66212 1 38
2 66213 1 38
2 66214 1 38
2 66215 1 38
2 66216 1 38
2 66217 1 38
2 66218 1 38
2 66219 1 38
2 66220 1 38
2 66221 1 38
2 66222 1 38
2 66223 1 38
2 66224 1 38
2 66225 1 38
2 66226 1 38
2 66227 1 38
2 66228 1 38
2 66229 1 38
2 66230 1 38
2 66231 1 38
2 66232 1 38
2 66233 1 38
2 66234 1 38
2 66235 1 38
2 66236 1 38
2 66237 1 38
2 66238 1 38
2 66239 1 38
2 66240 1 38
2 66241 1 38
2 66242 1 38
2 66243 1 38
2 66244 1 38
2 66245 1 38
2 66246 1 38
2 66247 1 38
2 66248 1 38
2 66249 1 38
2 66250 1 38
2 66251 1 38
2 66252 1 38
2 66253 1 38
2 66254 1 38
2 66255 1 38
2 66256 1 38
2 66257 1 38
2 66258 1 38
2 66259 1 38
2 66260 1 38
2 66261 1 38
2 66262 1 38
2 66263 1 38
2 66264 1 38
2 66265 1 38
2 66266 1 38
2 66267 1 38
2 66268 1 38
2 66269 1 38
2 66270 1 38
2 66271 1 38
2 66272 1 38
2 66273 1 38
2 66274 1 38
2 66275 1 38
2 66276 1 38
2 66277 1 38
2 66278 1 38
2 66279 1 38
2 66280 1 38
2 66281 1 38
2 66282 1 38
2 66283 1 38
2 66284 1 38
2 66285 1 38
2 66286 1 38
2 66287 1 38
2 66288 1 38
2 66289 1 38
2 66290 1 38
2 66291 1 38
2 66292 1 38
2 66293 1 38
2 66294 1 38
2 66295 1 38
2 66296 1 38
2 66297 1 38
2 66298 1 38
2 66299 1 38
2 66300 1 38
2 66301 1 38
2 66302 1 38
2 66303 1 38
2 66304 1 38
2 66305 1 38
2 66306 1 38
2 66307 1 38
2 66308 1 38
2 66309 1 38
2 66310 1 38
2 66311 1 38
2 66312 1 38
2 66313 1 38
2 66314 1 38
2 66315 1 38
2 66316 1 38
2 66317 1 38
2 66318 1 38
2 66319 1 38
2 66320 1 38
2 66321 1 38
2 66322 1 38
2 66323 1 38
2 66324 1 38
2 66325 1 38
2 66326 1 38
2 66327 1 38
2 66328 1 38
2 66329 1 38
2 66330 1 38
2 66331 1 38
2 66332 1 38
2 66333 1 38
2 66334 1 38
2 66335 1 38
2 66336 1 38
2 66337 1 38
2 66338 1 38
2 66339 1 38
2 66340 1 38
2 66341 1 38
2 66342 1 38
2 66343 1 38
2 66344 1 38
2 66345 1 38
2 66346 1 38
2 66347 1 39
2 66348 1 39
2 66349 1 39
2 66350 1 39
2 66351 1 39
2 66352 1 39
2 66353 1 39
2 66354 1 39
2 66355 1 39
2 66356 1 39
2 66357 1 39
2 66358 1 39
2 66359 1 39
2 66360 1 39
2 66361 1 39
2 66362 1 39
2 66363 1 39
2 66364 1 39
2 66365 1 39
2 66366 1 39
2 66367 1 39
2 66368 1 39
2 66369 1 39
2 66370 1 39
2 66371 1 39
2 66372 1 39
2 66373 1 39
2 66374 1 39
2 66375 1 39
2 66376 1 39
2 66377 1 39
2 66378 1 39
2 66379 1 39
2 66380 1 39
2 66381 1 39
2 66382 1 39
2 66383 1 39
2 66384 1 39
2 66385 1 39
2 66386 1 39
2 66387 1 39
2 66388 1 39
2 66389 1 39
2 66390 1 39
2 66391 1 39
2 66392 1 39
2 66393 1 39
2 66394 1 39
2 66395 1 39
2 66396 1 39
2 66397 1 39
2 66398 1 39
2 66399 1 39
2 66400 1 39
2 66401 1 39
2 66402 1 39
2 66403 1 39
2 66404 1 39
2 66405 1 39
2 66406 1 39
2 66407 1 39
2 66408 1 39
2 66409 1 39
2 66410 1 39
2 66411 1 39
2 66412 1 39
2 66413 1 39
2 66414 1 39
2 66415 1 39
2 66416 1 39
2 66417 1 39
2 66418 1 39
2 66419 1 39
2 66420 1 39
2 66421 1 39
2 66422 1 39
2 66423 1 39
2 66424 1 39
2 66425 1 39
2 66426 1 39
2 66427 1 39
2 66428 1 39
2 66429 1 39
2 66430 1 39
2 66431 1 39
2 66432 1 39
2 66433 1 39
2 66434 1 39
2 66435 1 39
2 66436 1 39
2 66437 1 39
2 66438 1 39
2 66439 1 39
2 66440 1 39
2 66441 1 39
2 66442 1 39
2 66443 1 39
2 66444 1 39
2 66445 1 39
2 66446 1 39
2 66447 1 39
2 66448 1 39
2 66449 1 39
2 66450 1 39
2 66451 1 39
2 66452 1 39
2 66453 1 39
2 66454 1 39
2 66455 1 39
2 66456 1 39
2 66457 1 39
2 66458 1 39
2 66459 1 39
2 66460 1 39
2 66461 1 39
2 66462 1 39
2 66463 1 39
2 66464 1 39
2 66465 1 39
2 66466 1 39
2 66467 1 39
2 66468 1 39
2 66469 1 39
2 66470 1 39
2 66471 1 39
2 66472 1 39
2 66473 1 39
2 66474 1 39
2 66475 1 39
2 66476 1 39
2 66477 1 39
2 66478 1 39
2 66479 1 39
2 66480 1 39
2 66481 1 39
2 66482 1 39
2 66483 1 39
2 66484 1 39
2 66485 1 39
2 66486 1 39
2 66487 1 39
2 66488 1 39
2 66489 1 39
2 66490 1 39
2 66491 1 39
2 66492 1 39
2 66493 1 39
2 66494 1 39
2 66495 1 39
2 66496 1 39
2 66497 1 39
2 66498 1 39
2 66499 1 39
2 66500 1 39
2 66501 1 39
2 66502 1 39
2 66503 1 39
2 66504 1 39
2 66505 1 39
2 66506 1 39
2 66507 1 39
2 66508 1 39
2 66509 1 39
2 66510 1 39
2 66511 1 39
2 66512 1 39
2 66513 1 39
2 66514 1 39
2 66515 1 39
2 66516 1 39
2 66517 1 39
2 66518 1 39
2 66519 1 39
2 66520 1 39
2 66521 1 39
2 66522 1 39
2 66523 1 39
2 66524 1 39
2 66525 1 39
2 66526 1 39
2 66527 1 39
2 66528 1 39
2 66529 1 39
2 66530 1 39
2 66531 1 39
2 66532 1 39
2 66533 1 39
2 66534 1 39
2 66535 1 39
2 66536 1 39
2 66537 1 39
2 66538 1 39
2 66539 1 39
2 66540 1 39
2 66541 1 39
2 66542 1 39
2 66543 1 39
2 66544 1 39
2 66545 1 39
2 66546 1 39
2 66547 1 39
2 66548 1 39
2 66549 1 39
2 66550 1 39
2 66551 1 39
2 66552 1 39
2 66553 1 39
2 66554 1 39
2 66555 1 39
2 66556 1 39
2 66557 1 39
2 66558 1 39
2 66559 1 39
2 66560 1 39
2 66561 1 39
2 66562 1 39
2 66563 1 39
2 66564 1 39
2 66565 1 39
2 66566 1 39
2 66567 1 39
2 66568 1 39
2 66569 1 39
2 66570 1 39
2 66571 1 39
2 66572 1 39
2 66573 1 39
2 66574 1 39
2 66575 1 39
2 66576 1 39
2 66577 1 39
2 66578 1 39
2 66579 1 39
2 66580 1 39
2 66581 1 39
2 66582 1 39
2 66583 1 39
2 66584 1 39
2 66585 1 39
2 66586 1 39
2 66587 1 39
2 66588 1 39
2 66589 1 39
2 66590 1 39
2 66591 1 39
2 66592 1 39
2 66593 1 39
2 66594 1 39
2 66595 1 39
2 66596 1 39
2 66597 1 39
2 66598 1 39
2 66599 1 39
2 66600 1 39
2 66601 1 39
2 66602 1 39
2 66603 1 39
2 66604 1 39
2 66605 1 39
2 66606 1 39
2 66607 1 40
2 66608 1 40
2 66609 1 40
2 66610 1 40
2 66611 1 40
2 66612 1 40
2 66613 1 40
2 66614 1 40
2 66615 1 40
2 66616 1 40
2 66617 1 40
2 66618 1 40
2 66619 1 40
2 66620 1 40
2 66621 1 40
2 66622 1 40
2 66623 1 40
2 66624 1 40
2 66625 1 40
2 66626 1 40
2 66627 1 40
2 66628 1 40
2 66629 1 40
2 66630 1 40
2 66631 1 40
2 66632 1 40
2 66633 1 40
2 66634 1 40
2 66635 1 40
2 66636 1 40
2 66637 1 40
2 66638 1 40
2 66639 1 40
2 66640 1 40
2 66641 1 40
2 66642 1 40
2 66643 1 40
2 66644 1 40
2 66645 1 40
2 66646 1 40
2 66647 1 40
2 66648 1 40
2 66649 1 40
2 66650 1 40
2 66651 1 40
2 66652 1 40
2 66653 1 40
2 66654 1 40
2 66655 1 40
2 66656 1 40
2 66657 1 40
2 66658 1 40
2 66659 1 40
2 66660 1 40
2 66661 1 40
2 66662 1 40
2 66663 1 40
2 66664 1 40
2 66665 1 40
2 66666 1 40
2 66667 1 40
2 66668 1 40
2 66669 1 40
2 66670 1 40
2 66671 1 40
2 66672 1 40
2 66673 1 40
2 66674 1 40
2 66675 1 40
2 66676 1 40
2 66677 1 40
2 66678 1 40
2 66679 1 40
2 66680 1 40
2 66681 1 40
2 66682 1 40
2 66683 1 40
2 66684 1 40
2 66685 1 40
2 66686 1 40
2 66687 1 40
2 66688 1 40
2 66689 1 40
2 66690 1 40
2 66691 1 40
2 66692 1 40
2 66693 1 40
2 66694 1 40
2 66695 1 40
2 66696 1 40
2 66697 1 40
2 66698 1 40
2 66699 1 40
2 66700 1 40
2 66701 1 40
2 66702 1 40
2 66703 1 40
2 66704 1 40
2 66705 1 40
2 66706 1 40
2 66707 1 40
2 66708 1 40
2 66709 1 40
2 66710 1 40
2 66711 1 40
2 66712 1 40
2 66713 1 40
2 66714 1 40
2 66715 1 40
2 66716 1 40
2 66717 1 40
2 66718 1 40
2 66719 1 40
2 66720 1 40
2 66721 1 40
2 66722 1 40
2 66723 1 40
2 66724 1 40
2 66725 1 40
2 66726 1 40
2 66727 1 40
2 66728 1 40
2 66729 1 40
2 66730 1 40
2 66731 1 40
2 66732 1 40
2 66733 1 40
2 66734 1 40
2 66735 1 40
2 66736 1 40
2 66737 1 40
2 66738 1 40
2 66739 1 40
2 66740 1 40
2 66741 1 40
2 66742 1 40
2 66743 1 40
2 66744 1 40
2 66745 1 40
2 66746 1 40
2 66747 1 40
2 66748 1 40
2 66749 1 40
2 66750 1 40
2 66751 1 40
2 66752 1 40
2 66753 1 40
2 66754 1 40
2 66755 1 40
2 66756 1 40
2 66757 1 40
2 66758 1 40
2 66759 1 40
2 66760 1 40
2 66761 1 40
2 66762 1 40
2 66763 1 40
2 66764 1 40
2 66765 1 40
2 66766 1 40
2 66767 1 40
2 66768 1 40
2 66769 1 40
2 66770 1 40
2 66771 1 40
2 66772 1 40
2 66773 1 40
2 66774 1 40
2 66775 1 40
2 66776 1 40
2 66777 1 40
2 66778 1 40
2 66779 1 40
2 66780 1 40
2 66781 1 40
2 66782 1 40
2 66783 1 40
2 66784 1 40
2 66785 1 40
2 66786 1 40
2 66787 1 40
2 66788 1 40
2 66789 1 41
2 66790 1 41
2 66791 1 41
2 66792 1 41
2 66793 1 41
2 66794 1 41
2 66795 1 41
2 66796 1 41
2 66797 1 41
2 66798 1 41
2 66799 1 41
2 66800 1 41
2 66801 1 41
2 66802 1 41
2 66803 1 41
2 66804 1 41
2 66805 1 41
2 66806 1 41
2 66807 1 41
2 66808 1 41
2 66809 1 41
2 66810 1 41
2 66811 1 41
2 66812 1 41
2 66813 1 41
2 66814 1 41
2 66815 1 41
2 66816 1 41
2 66817 1 41
2 66818 1 41
2 66819 1 41
2 66820 1 41
2 66821 1 41
2 66822 1 41
2 66823 1 41
2 66824 1 41
2 66825 1 41
2 66826 1 41
2 66827 1 41
2 66828 1 41
2 66829 1 41
2 66830 1 41
2 66831 1 41
2 66832 1 41
2 66833 1 41
2 66834 1 41
2 66835 1 41
2 66836 1 41
2 66837 1 41
2 66838 1 41
2 66839 1 41
2 66840 1 41
2 66841 1 41
2 66842 1 41
2 66843 1 41
2 66844 1 41
2 66845 1 41
2 66846 1 41
2 66847 1 41
2 66848 1 41
2 66849 1 41
2 66850 1 41
2 66851 1 41
2 66852 1 41
2 66853 1 41
2 66854 1 41
2 66855 1 41
2 66856 1 41
2 66857 1 41
2 66858 1 41
2 66859 1 41
2 66860 1 41
2 66861 1 41
2 66862 1 41
2 66863 1 41
2 66864 1 41
2 66865 1 41
2 66866 1 41
2 66867 1 41
2 66868 1 41
2 66869 1 41
2 66870 1 41
2 66871 1 41
2 66872 1 41
2 66873 1 41
2 66874 1 41
2 66875 1 41
2 66876 1 41
2 66877 1 41
2 66878 1 41
2 66879 1 41
2 66880 1 41
2 66881 1 41
2 66882 1 41
2 66883 1 41
2 66884 1 41
2 66885 1 41
2 66886 1 41
2 66887 1 41
2 66888 1 41
2 66889 1 41
2 66890 1 41
2 66891 1 41
2 66892 1 41
2 66893 1 41
2 66894 1 41
2 66895 1 41
2 66896 1 41
2 66897 1 41
2 66898 1 41
2 66899 1 41
2 66900 1 41
2 66901 1 41
2 66902 1 41
2 66903 1 41
2 66904 1 41
2 66905 1 41
2 66906 1 41
2 66907 1 41
2 66908 1 41
2 66909 1 41
2 66910 1 41
2 66911 1 41
2 66912 1 41
2 66913 1 41
2 66914 1 41
2 66915 1 41
2 66916 1 41
2 66917 1 41
2 66918 1 41
2 66919 1 41
2 66920 1 41
2 66921 1 41
2 66922 1 41
2 66923 1 41
2 66924 1 41
2 66925 1 41
2 66926 1 41
2 66927 1 41
2 66928 1 41
2 66929 1 41
2 66930 1 41
2 66931 1 41
2 66932 1 41
2 66933 1 41
2 66934 1 41
2 66935 1 41
2 66936 1 41
2 66937 1 41
2 66938 1 41
2 66939 1 41
2 66940 1 41
2 66941 1 41
2 66942 1 42
2 66943 1 42
2 66944 1 42
2 66945 1 42
2 66946 1 42
2 66947 1 42
2 66948 1 42
2 66949 1 42
2 66950 1 42
2 66951 1 42
2 66952 1 42
2 66953 1 42
2 66954 1 42
2 66955 1 42
2 66956 1 43
2 66957 1 43
2 66958 1 43
2 66959 1 43
2 66960 1 43
2 66961 1 43
2 66962 1 43
2 66963 1 43
2 66964 1 43
2 66965 1 43
2 66966 1 43
2 66967 1 43
2 66968 1 43
2 66969 1 43
2 66970 1 43
2 66971 1 43
2 66972 1 43
2 66973 1 43
2 66974 1 43
2 66975 1 43
2 66976 1 43
2 66977 1 43
2 66978 1 43
2 66979 1 43
2 66980 1 43
2 66981 1 43
2 66982 1 43
2 66983 1 43
2 66984 1 43
2 66985 1 43
2 66986 1 43
2 66987 1 43
2 66988 1 43
2 66989 1 43
2 66990 1 43
2 66991 1 43
2 66992 1 43
2 66993 1 43
2 66994 1 43
2 66995 1 43
2 66996 1 43
2 66997 1 43
2 66998 1 43
2 66999 1 43
2 67000 1 43
2 67001 1 43
2 67002 1 43
2 67003 1 43
2 67004 1 43
2 67005 1 43
2 67006 1 43
2 67007 1 43
2 67008 1 43
2 67009 1 43
2 67010 1 43
2 67011 1 43
2 67012 1 43
2 67013 1 43
2 67014 1 43
2 67015 1 43
2 67016 1 43
2 67017 1 43
2 67018 1 43
2 67019 1 43
2 67020 1 43
2 67021 1 43
2 67022 1 43
2 67023 1 43
2 67024 1 43
2 67025 1 43
2 67026 1 43
2 67027 1 43
2 67028 1 43
2 67029 1 43
2 67030 1 43
2 67031 1 43
2 67032 1 43
2 67033 1 43
2 67034 1 43
2 67035 1 43
2 67036 1 43
2 67037 1 43
2 67038 1 43
2 67039 1 43
2 67040 1 43
2 67041 1 43
2 67042 1 43
2 67043 1 43
2 67044 1 43
2 67045 1 43
2 67046 1 43
2 67047 1 43
2 67048 1 43
2 67049 1 43
2 67050 1 43
2 67051 1 43
2 67052 1 43
2 67053 1 43
2 67054 1 43
2 67055 1 43
2 67056 1 43
2 67057 1 43
2 67058 1 43
2 67059 1 43
2 67060 1 43
2 67061 1 43
2 67062 1 43
2 67063 1 43
2 67064 1 43
2 67065 1 43
2 67066 1 43
2 67067 1 43
2 67068 1 43
2 67069 1 43
2 67070 1 43
2 67071 1 43
2 67072 1 43
2 67073 1 43
2 67074 1 43
2 67075 1 43
2 67076 1 43
2 67077 1 43
2 67078 1 43
2 67079 1 43
2 67080 1 43
2 67081 1 43
2 67082 1 43
2 67083 1 43
2 67084 1 43
2 67085 1 43
2 67086 1 43
2 67087 1 43
2 67088 1 43
2 67089 1 43
2 67090 1 43
2 67091 1 43
2 67092 1 43
2 67093 1 43
2 67094 1 43
2 67095 1 43
2 67096 1 43
2 67097 1 43
2 67098 1 43
2 67099 1 43
2 67100 1 43
2 67101 1 43
2 67102 1 43
2 67103 1 43
2 67104 1 43
2 67105 1 43
2 67106 1 43
2 67107 1 43
2 67108 1 43
2 67109 1 43
2 67110 1 43
2 67111 1 43
2 67112 1 43
2 67113 1 43
2 67114 1 43
2 67115 1 43
2 67116 1 43
2 67117 1 43
2 67118 1 43
2 67119 1 43
2 67120 1 43
2 67121 1 43
2 67122 1 43
2 67123 1 43
2 67124 1 43
2 67125 1 43
2 67126 1 43
2 67127 1 43
2 67128 1 43
2 67129 1 43
2 67130 1 43
2 67131 1 43
2 67132 1 43
2 67133 1 43
2 67134 1 43
2 67135 1 43
2 67136 1 43
2 67137 1 43
2 67138 1 43
2 67139 1 43
2 67140 1 43
2 67141 1 43
2 67142 1 43
2 67143 1 43
2 67144 1 43
2 67145 1 43
2 67146 1 43
2 67147 1 43
2 67148 1 43
2 67149 1 43
2 67150 1 43
2 67151 1 43
2 67152 1 43
2 67153 1 43
2 67154 1 43
2 67155 1 43
2 67156 1 43
2 67157 1 43
2 67158 1 43
2 67159 1 43
2 67160 1 44
2 67161 1 44
2 67162 1 44
2 67163 1 44
2 67164 1 44
2 67165 1 44
2 67166 1 44
2 67167 1 44
2 67168 1 44
2 67169 1 44
2 67170 1 44
2 67171 1 44
2 67172 1 44
2 67173 1 44
2 67174 1 44
2 67175 1 44
2 67176 1 44
2 67177 1 44
2 67178 1 44
2 67179 1 44
2 67180 1 44
2 67181 1 44
2 67182 1 44
2 67183 1 44
2 67184 1 44
2 67185 1 44
2 67186 1 44
2 67187 1 44
2 67188 1 44
2 67189 1 44
2 67190 1 44
2 67191 1 44
2 67192 1 44
2 67193 1 44
2 67194 1 44
2 67195 1 44
2 67196 1 44
2 67197 1 44
2 67198 1 44
2 67199 1 44
2 67200 1 44
2 67201 1 44
2 67202 1 44
2 67203 1 44
2 67204 1 44
2 67205 1 44
2 67206 1 44
2 67207 1 44
2 67208 1 44
2 67209 1 44
2 67210 1 44
2 67211 1 44
2 67212 1 44
2 67213 1 44
2 67214 1 44
2 67215 1 44
2 67216 1 44
2 67217 1 44
2 67218 1 44
2 67219 1 44
2 67220 1 44
2 67221 1 44
2 67222 1 44
2 67223 1 44
2 67224 1 44
2 67225 1 44
2 67226 1 44
2 67227 1 44
2 67228 1 44
2 67229 1 44
2 67230 1 44
2 67231 1 44
2 67232 1 44
2 67233 1 44
2 67234 1 44
2 67235 1 44
2 67236 1 44
2 67237 1 44
2 67238 1 44
2 67239 1 44
2 67240 1 44
2 67241 1 44
2 67242 1 44
2 67243 1 44
2 67244 1 44
2 67245 1 44
2 67246 1 44
2 67247 1 44
2 67248 1 44
2 67249 1 44
2 67250 1 44
2 67251 1 44
2 67252 1 44
2 67253 1 44
2 67254 1 44
2 67255 1 44
2 67256 1 44
2 67257 1 44
2 67258 1 44
2 67259 1 44
2 67260 1 44
2 67261 1 44
2 67262 1 44
2 67263 1 44
2 67264 1 44
2 67265 1 44
2 67266 1 44
2 67267 1 44
2 67268 1 44
2 67269 1 44
2 67270 1 44
2 67271 1 44
2 67272 1 44
2 67273 1 44
2 67274 1 44
2 67275 1 44
2 67276 1 44
2 67277 1 44
2 67278 1 44
2 67279 1 44
2 67280 1 44
2 67281 1 44
2 67282 1 44
2 67283 1 44
2 67284 1 44
2 67285 1 44
2 67286 1 44
2 67287 1 44
2 67288 1 44
2 67289 1 44
2 67290 1 44
2 67291 1 44
2 67292 1 44
2 67293 1 44
2 67294 1 44
2 67295 1 44
2 67296 1 44
2 67297 1 44
2 67298 1 44
2 67299 1 44
2 67300 1 44
2 67301 1 44
2 67302 1 44
2 67303 1 44
2 67304 1 44
2 67305 1 44
2 67306 1 44
2 67307 1 44
2 67308 1 44
2 67309 1 44
2 67310 1 44
2 67311 1 44
2 67312 1 44
2 67313 1 44
2 67314 1 44
2 67315 1 44
2 67316 1 44
2 67317 1 44
2 67318 1 44
2 67319 1 44
2 67320 1 44
2 67321 1 44
2 67322 1 44
2 67323 1 44
2 67324 1 44
2 67325 1 44
2 67326 1 44
2 67327 1 44
2 67328 1 44
2 67329 1 44
2 67330 1 44
2 67331 1 44
2 67332 1 44
2 67333 1 44
2 67334 1 44
2 67335 1 44
2 67336 1 44
2 67337 1 44
2 67338 1 44
2 67339 1 44
2 67340 1 44
2 67341 1 44
2 67342 1 44
2 67343 1 44
2 67344 1 44
2 67345 1 44
2 67346 1 44
2 67347 1 44
2 67348 1 44
2 67349 1 44
2 67350 1 44
2 67351 1 44
2 67352 1 44
2 67353 1 44
2 67354 1 44
2 67355 1 44
2 67356 1 44
2 67357 1 44
2 67358 1 44
2 67359 1 44
2 67360 1 44
2 67361 1 44
2 67362 1 44
2 67363 1 44
2 67364 1 44
2 67365 1 44
2 67366 1 44
2 67367 1 44
2 67368 1 44
2 67369 1 44
2 67370 1 44
2 67371 1 44
2 67372 1 44
2 67373 1 44
2 67374 1 44
2 67375 1 44
2 67376 1 44
2 67377 1 44
2 67378 1 44
2 67379 1 44
2 67380 1 44
2 67381 1 44
2 67382 1 44
2 67383 1 44
2 67384 1 44
2 67385 1 44
2 67386 1 44
2 67387 1 44
2 67388 1 44
2 67389 1 44
2 67390 1 44
2 67391 1 44
2 67392 1 44
2 67393 1 44
2 67394 1 44
2 67395 1 44
2 67396 1 44
2 67397 1 44
2 67398 1 44
2 67399 1 44
2 67400 1 45
2 67401 1 45
2 67402 1 45
2 67403 1 45
2 67404 1 45
2 67405 1 45
2 67406 1 45
2 67407 1 45
2 67408 1 45
2 67409 1 45
2 67410 1 45
2 67411 1 45
2 67412 1 45
2 67413 1 45
2 67414 1 45
2 67415 1 45
2 67416 1 45
2 67417 1 45
2 67418 1 45
2 67419 1 45
2 67420 1 45
2 67421 1 45
2 67422 1 45
2 67423 1 45
2 67424 1 45
2 67425 1 45
2 67426 1 45
2 67427 1 45
2 67428 1 45
2 67429 1 45
2 67430 1 45
2 67431 1 45
2 67432 1 45
2 67433 1 45
2 67434 1 45
2 67435 1 45
2 67436 1 45
2 67437 1 45
2 67438 1 45
2 67439 1 45
2 67440 1 45
2 67441 1 45
2 67442 1 45
2 67443 1 45
2 67444 1 45
2 67445 1 45
2 67446 1 45
2 67447 1 45
2 67448 1 45
2 67449 1 45
2 67450 1 45
2 67451 1 45
2 67452 1 45
2 67453 1 45
2 67454 1 45
2 67455 1 45
2 67456 1 45
2 67457 1 45
2 67458 1 45
2 67459 1 45
2 67460 1 45
2 67461 1 45
2 67462 1 45
2 67463 1 45
2 67464 1 45
2 67465 1 45
2 67466 1 45
2 67467 1 45
2 67468 1 45
2 67469 1 45
2 67470 1 45
2 67471 1 45
2 67472 1 45
2 67473 1 45
2 67474 1 45
2 67475 1 45
2 67476 1 45
2 67477 1 45
2 67478 1 45
2 67479 1 45
2 67480 1 45
2 67481 1 45
2 67482 1 45
2 67483 1 45
2 67484 1 45
2 67485 1 45
2 67486 1 45
2 67487 1 45
2 67488 1 45
2 67489 1 45
2 67490 1 45
2 67491 1 45
2 67492 1 45
2 67493 1 45
2 67494 1 45
2 67495 1 45
2 67496 1 45
2 67497 1 45
2 67498 1 45
2 67499 1 45
2 67500 1 45
2 67501 1 45
2 67502 1 45
2 67503 1 45
2 67504 1 45
2 67505 1 45
2 67506 1 45
2 67507 1 45
2 67508 1 45
2 67509 1 45
2 67510 1 45
2 67511 1 45
2 67512 1 45
2 67513 1 45
2 67514 1 45
2 67515 1 45
2 67516 1 45
2 67517 1 45
2 67518 1 45
2 67519 1 45
2 67520 1 45
2 67521 1 45
2 67522 1 45
2 67523 1 45
2 67524 1 45
2 67525 1 45
2 67526 1 45
2 67527 1 45
2 67528 1 45
2 67529 1 45
2 67530 1 45
2 67531 1 45
2 67532 1 45
2 67533 1 45
2 67534 1 45
2 67535 1 45
2 67536 1 45
2 67537 1 45
2 67538 1 45
2 67539 1 45
2 67540 1 45
2 67541 1 45
2 67542 1 45
2 67543 1 45
2 67544 1 45
2 67545 1 45
2 67546 1 45
2 67547 1 45
2 67548 1 45
2 67549 1 45
2 67550 1 45
2 67551 1 45
2 67552 1 45
2 67553 1 45
2 67554 1 45
2 67555 1 45
2 67556 1 45
2 67557 1 45
2 67558 1 45
2 67559 1 45
2 67560 1 45
2 67561 1 45
2 67562 1 45
2 67563 1 45
2 67564 1 45
2 67565 1 45
2 67566 1 45
2 67567 1 45
2 67568 1 45
2 67569 1 45
2 67570 1 45
2 67571 1 45
2 67572 1 45
2 67573 1 45
2 67574 1 45
2 67575 1 45
2 67576 1 45
2 67577 1 45
2 67578 1 45
2 67579 1 45
2 67580 1 45
2 67581 1 45
2 67582 1 45
2 67583 1 45
2 67584 1 45
2 67585 1 45
2 67586 1 45
2 67587 1 45
2 67588 1 45
2 67589 1 45
2 67590 1 45
2 67591 1 45
2 67592 1 45
2 67593 1 45
2 67594 1 45
2 67595 1 45
2 67596 1 45
2 67597 1 45
2 67598 1 45
2 67599 1 45
2 67600 1 45
2 67601 1 45
2 67602 1 45
2 67603 1 45
2 67604 1 45
2 67605 1 45
2 67606 1 45
2 67607 1 45
2 67608 1 45
2 67609 1 45
2 67610 1 45
2 67611 1 45
2 67612 1 45
2 67613 1 45
2 67614 1 45
2 67615 1 45
2 67616 1 45
2 67617 1 45
2 67618 1 45
2 67619 1 45
2 67620 1 45
2 67621 1 45
2 67622 1 45
2 67623 1 45
2 67624 1 45
2 67625 1 45
2 67626 1 45
2 67627 1 45
2 67628 1 45
2 67629 1 45
2 67630 1 45
2 67631 1 45
2 67632 1 45
2 67633 1 45
2 67634 1 45
2 67635 1 45
2 67636 1 45
2 67637 1 45
2 67638 1 45
2 67639 1 45
2 67640 1 45
2 67641 1 45
2 67642 1 45
2 67643 1 45
2 67644 1 45
2 67645 1 45
2 67646 1 45
2 67647 1 45
2 67648 1 45
2 67649 1 45
2 67650 1 45
2 67651 1 45
2 67652 1 45
2 67653 1 45
2 67654 1 45
2 67655 1 45
2 67656 1 45
2 67657 1 45
2 67658 1 45
2 67659 1 45
2 67660 1 45
2 67661 1 45
2 67662 1 45
2 67663 1 45
2 67664 1 45
2 67665 1 45
2 67666 1 45
2 67667 1 45
2 67668 1 45
2 67669 1 45
2 67670 1 45
2 67671 1 45
2 67672 1 45
2 67673 1 45
2 67674 1 45
2 67675 1 45
2 67676 1 45
2 67677 1 45
2 67678 1 45
2 67679 1 45
2 67680 1 45
2 67681 1 45
2 67682 1 45
2 67683 1 45
2 67684 1 45
2 67685 1 45
2 67686 1 45
2 67687 1 45
2 67688 1 45
2 67689 1 45
2 67690 1 45
2 67691 1 45
2 67692 1 45
2 67693 1 45
2 67694 1 45
2 67695 1 45
2 67696 1 45
2 67697 1 45
2 67698 1 45
2 67699 1 45
2 67700 1 45
2 67701 1 45
2 67702 1 45
2 67703 1 45
2 67704 1 45
2 67705 1 45
2 67706 1 45
2 67707 1 45
2 67708 1 45
2 67709 1 45
2 67710 1 45
2 67711 1 45
2 67712 1 45
2 67713 1 45
2 67714 1 45
2 67715 1 45
2 67716 1 45
2 67717 1 45
2 67718 1 45
2 67719 1 45
2 67720 1 45
2 67721 1 45
2 67722 1 45
2 67723 1 45
2 67724 1 45
2 67725 1 45
2 67726 1 45
2 67727 1 45
2 67728 1 45
2 67729 1 45
2 67730 1 45
2 67731 1 45
2 67732 1 45
2 67733 1 45
2 67734 1 45
2 67735 1 45
2 67736 1 45
2 67737 1 45
2 67738 1 45
2 67739 1 45
2 67740 1 45
2 67741 1 45
2 67742 1 45
2 67743 1 45
2 67744 1 45
2 67745 1 45
2 67746 1 45
2 67747 1 45
2 67748 1 45
2 67749 1 45
2 67750 1 45
2 67751 1 45
2 67752 1 45
2 67753 1 45
2 67754 1 45
2 67755 1 45
2 67756 1 45
2 67757 1 45
2 67758 1 45
2 67759 1 45
2 67760 1 45
2 67761 1 45
2 67762 1 45
2 67763 1 45
2 67764 1 45
2 67765 1 45
2 67766 1 45
2 67767 1 45
2 67768 1 45
2 67769 1 45
2 67770 1 45
2 67771 1 45
2 67772 1 45
2 67773 1 45
2 67774 1 45
2 67775 1 45
2 67776 1 45
2 67777 1 45
2 67778 1 45
2 67779 1 45
2 67780 1 45
2 67781 1 45
2 67782 1 45
2 67783 1 45
2 67784 1 45
2 67785 1 45
2 67786 1 45
2 67787 1 45
2 67788 1 45
2 67789 1 45
2 67790 1 45
2 67791 1 45
2 67792 1 45
2 67793 1 45
2 67794 1 45
2 67795 1 45
2 67796 1 45
2 67797 1 46
2 67798 1 46
2 67799 1 46
2 67800 1 46
2 67801 1 46
2 67802 1 46
2 67803 1 46
2 67804 1 46
2 67805 1 46
2 67806 1 46
2 67807 1 46
2 67808 1 46
2 67809 1 46
2 67810 1 46
2 67811 1 46
2 67812 1 46
2 67813 1 46
2 67814 1 46
2 67815 1 46
2 67816 1 46
2 67817 1 46
2 67818 1 46
2 67819 1 46
2 67820 1 46
2 67821 1 46
2 67822 1 46
2 67823 1 46
2 67824 1 46
2 67825 1 46
2 67826 1 46
2 67827 1 46
2 67828 1 46
2 67829 1 46
2 67830 1 46
2 67831 1 46
2 67832 1 46
2 67833 1 46
2 67834 1 46
2 67835 1 46
2 67836 1 46
2 67837 1 46
2 67838 1 46
2 67839 1 46
2 67840 1 46
2 67841 1 46
2 67842 1 46
2 67843 1 46
2 67844 1 46
2 67845 1 46
2 67846 1 46
2 67847 1 46
2 67848 1 46
2 67849 1 46
2 67850 1 46
2 67851 1 46
2 67852 1 46
2 67853 1 46
2 67854 1 46
2 67855 1 46
2 67856 1 46
2 67857 1 46
2 67858 1 46
2 67859 1 46
2 67860 1 46
2 67861 1 46
2 67862 1 46
2 67863 1 46
2 67864 1 46
2 67865 1 46
2 67866 1 46
2 67867 1 46
2 67868 1 46
2 67869 1 46
2 67870 1 46
2 67871 1 46
2 67872 1 46
2 67873 1 46
2 67874 1 46
2 67875 1 46
2 67876 1 46
2 67877 1 46
2 67878 1 46
2 67879 1 46
2 67880 1 46
2 67881 1 46
2 67882 1 46
2 67883 1 46
2 67884 1 46
2 67885 1 46
2 67886 1 46
2 67887 1 46
2 67888 1 46
2 67889 1 46
2 67890 1 46
2 67891 1 46
2 67892 1 46
2 67893 1 46
2 67894 1 46
2 67895 1 46
2 67896 1 46
2 67897 1 46
2 67898 1 46
2 67899 1 46
2 67900 1 46
2 67901 1 46
2 67902 1 46
2 67903 1 46
2 67904 1 46
2 67905 1 46
2 67906 1 46
2 67907 1 46
2 67908 1 46
2 67909 1 46
2 67910 1 46
2 67911 1 46
2 67912 1 46
2 67913 1 46
2 67914 1 46
2 67915 1 46
2 67916 1 46
2 67917 1 46
2 67918 1 46
2 67919 1 46
2 67920 1 46
2 67921 1 46
2 67922 1 46
2 67923 1 46
2 67924 1 46
2 67925 1 46
2 67926 1 46
2 67927 1 46
2 67928 1 46
2 67929 1 46
2 67930 1 46
2 67931 1 46
2 67932 1 46
2 67933 1 46
2 67934 1 46
2 67935 1 46
2 67936 1 46
2 67937 1 46
2 67938 1 46
2 67939 1 46
2 67940 1 46
2 67941 1 46
2 67942 1 46
2 67943 1 46
2 67944 1 46
2 67945 1 46
2 67946 1 46
2 67947 1 46
2 67948 1 46
2 67949 1 46
2 67950 1 46
2 67951 1 46
2 67952 1 46
2 67953 1 46
2 67954 1 46
2 67955 1 46
2 67956 1 46
2 67957 1 46
2 67958 1 46
2 67959 1 46
2 67960 1 46
2 67961 1 46
2 67962 1 46
2 67963 1 46
2 67964 1 46
2 67965 1 46
2 67966 1 46
2 67967 1 46
2 67968 1 46
2 67969 1 46
2 67970 1 46
2 67971 1 46
2 67972 1 46
2 67973 1 46
2 67974 1 46
2 67975 1 46
2 67976 1 46
2 67977 1 46
2 67978 1 46
2 67979 1 46
2 67980 1 46
2 67981 1 46
2 67982 1 46
2 67983 1 46
2 67984 1 46
2 67985 1 46
2 67986 1 46
2 67987 1 46
2 67988 1 46
2 67989 1 46
2 67990 1 46
2 67991 1 46
2 67992 1 46
2 67993 1 46
2 67994 1 46
2 67995 1 46
2 67996 1 46
2 67997 1 46
2 67998 1 46
2 67999 1 46
2 68000 1 46
2 68001 1 46
2 68002 1 46
2 68003 1 46
2 68004 1 46
2 68005 1 46
2 68006 1 46
2 68007 1 46
2 68008 1 46
2 68009 1 46
2 68010 1 46
2 68011 1 46
2 68012 1 46
2 68013 1 46
2 68014 1 46
2 68015 1 46
2 68016 1 46
2 68017 1 46
2 68018 1 46
2 68019 1 46
2 68020 1 46
2 68021 1 46
2 68022 1 46
2 68023 1 46
2 68024 1 46
2 68025 1 46
2 68026 1 46
2 68027 1 46
2 68028 1 46
2 68029 1 46
2 68030 1 46
2 68031 1 46
2 68032 1 46
2 68033 1 46
2 68034 1 46
2 68035 1 46
2 68036 1 46
2 68037 1 46
2 68038 1 46
2 68039 1 46
2 68040 1 46
2 68041 1 46
2 68042 1 46
2 68043 1 46
2 68044 1 46
2 68045 1 46
2 68046 1 46
2 68047 1 46
2 68048 1 46
2 68049 1 46
2 68050 1 46
2 68051 1 46
2 68052 1 46
2 68053 1 46
2 68054 1 46
2 68055 1 46
2 68056 1 46
2 68057 1 46
2 68058 1 46
2 68059 1 46
2 68060 1 46
2 68061 1 46
2 68062 1 46
2 68063 1 46
2 68064 1 46
2 68065 1 46
2 68066 1 46
2 68067 1 46
2 68068 1 46
2 68069 1 46
2 68070 1 46
2 68071 1 46
2 68072 1 46
2 68073 1 46
2 68074 1 46
2 68075 1 46
2 68076 1 46
2 68077 1 46
2 68078 1 46
2 68079 1 46
2 68080 1 46
2 68081 1 46
2 68082 1 46
2 68083 1 46
2 68084 1 46
2 68085 1 46
2 68086 1 46
2 68087 1 46
2 68088 1 46
2 68089 1 46
2 68090 1 46
2 68091 1 46
2 68092 1 46
2 68093 1 46
2 68094 1 46
2 68095 1 46
2 68096 1 46
2 68097 1 46
2 68098 1 46
2 68099 1 46
2 68100 1 46
2 68101 1 46
2 68102 1 46
2 68103 1 46
2 68104 1 46
2 68105 1 46
2 68106 1 46
2 68107 1 46
2 68108 1 46
2 68109 1 46
2 68110 1 46
2 68111 1 46
2 68112 1 46
2 68113 1 46
2 68114 1 46
2 68115 1 46
2 68116 1 46
2 68117 1 46
2 68118 1 46
2 68119 1 46
2 68120 1 46
2 68121 1 46
2 68122 1 46
2 68123 1 46
2 68124 1 46
2 68125 1 46
2 68126 1 46
2 68127 1 46
2 68128 1 46
2 68129 1 46
2 68130 1 46
2 68131 1 46
2 68132 1 46
2 68133 1 46
2 68134 1 46
2 68135 1 46
2 68136 1 46
2 68137 1 46
2 68138 1 46
2 68139 1 46
2 68140 1 46
2 68141 1 46
2 68142 1 46
2 68143 1 46
2 68144 1 46
2 68145 1 46
2 68146 1 46
2 68147 1 46
2 68148 1 46
2 68149 1 46
2 68150 1 46
2 68151 1 46
2 68152 1 46
2 68153 1 46
2 68154 1 46
2 68155 1 46
2 68156 1 46
2 68157 1 46
2 68158 1 46
2 68159 1 46
2 68160 1 46
2 68161 1 46
2 68162 1 46
2 68163 1 46
2 68164 1 46
2 68165 1 46
2 68166 1 46
2 68167 1 46
2 68168 1 46
2 68169 1 46
2 68170 1 46
2 68171 1 46
2 68172 1 46
2 68173 1 46
2 68174 1 46
2 68175 1 46
2 68176 1 46
2 68177 1 46
2 68178 1 46
2 68179 1 46
2 68180 1 46
2 68181 1 46
2 68182 1 46
2 68183 1 46
2 68184 1 46
2 68185 1 46
2 68186 1 46
2 68187 1 46
2 68188 1 47
2 68189 1 47
2 68190 1 47
2 68191 1 47
2 68192 1 47
2 68193 1 47
2 68194 1 47
2 68195 1 47
2 68196 1 47
2 68197 1 47
2 68198 1 47
2 68199 1 47
2 68200 1 47
2 68201 1 47
2 68202 1 47
2 68203 1 47
2 68204 1 47
2 68205 1 47
2 68206 1 47
2 68207 1 47
2 68208 1 47
2 68209 1 47
2 68210 1 47
2 68211 1 47
2 68212 1 47
2 68213 1 47
2 68214 1 47
2 68215 1 47
2 68216 1 47
2 68217 1 47
2 68218 1 47
2 68219 1 47
2 68220 1 47
2 68221 1 47
2 68222 1 47
2 68223 1 47
2 68224 1 47
2 68225 1 47
2 68226 1 47
2 68227 1 47
2 68228 1 47
2 68229 1 47
2 68230 1 47
2 68231 1 47
2 68232 1 47
2 68233 1 47
2 68234 1 47
2 68235 1 47
2 68236 1 47
2 68237 1 47
2 68238 1 47
2 68239 1 47
2 68240 1 47
2 68241 1 47
2 68242 1 47
2 68243 1 47
2 68244 1 47
2 68245 1 47
2 68246 1 47
2 68247 1 47
2 68248 1 47
2 68249 1 47
2 68250 1 47
2 68251 1 47
2 68252 1 47
2 68253 1 47
2 68254 1 47
2 68255 1 47
2 68256 1 47
2 68257 1 47
2 68258 1 47
2 68259 1 47
2 68260 1 47
2 68261 1 47
2 68262 1 47
2 68263 1 47
2 68264 1 47
2 68265 1 47
2 68266 1 47
2 68267 1 47
2 68268 1 47
2 68269 1 47
2 68270 1 47
2 68271 1 47
2 68272 1 47
2 68273 1 47
2 68274 1 47
2 68275 1 47
2 68276 1 47
2 68277 1 47
2 68278 1 47
2 68279 1 47
2 68280 1 47
2 68281 1 47
2 68282 1 47
2 68283 1 47
2 68284 1 47
2 68285 1 47
2 68286 1 47
2 68287 1 47
2 68288 1 47
2 68289 1 47
2 68290 1 47
2 68291 1 47
2 68292 1 47
2 68293 1 47
2 68294 1 47
2 68295 1 47
2 68296 1 47
2 68297 1 47
2 68298 1 47
2 68299 1 47
2 68300 1 47
2 68301 1 47
2 68302 1 47
2 68303 1 47
2 68304 1 47
2 68305 1 47
2 68306 1 47
2 68307 1 47
2 68308 1 47
2 68309 1 47
2 68310 1 47
2 68311 1 47
2 68312 1 47
2 68313 1 47
2 68314 1 47
2 68315 1 47
2 68316 1 47
2 68317 1 47
2 68318 1 47
2 68319 1 47
2 68320 1 47
2 68321 1 47
2 68322 1 47
2 68323 1 47
2 68324 1 47
2 68325 1 47
2 68326 1 47
2 68327 1 47
2 68328 1 47
2 68329 1 47
2 68330 1 47
2 68331 1 47
2 68332 1 47
2 68333 1 47
2 68334 1 47
2 68335 1 47
2 68336 1 47
2 68337 1 47
2 68338 1 47
2 68339 1 47
2 68340 1 47
2 68341 1 47
2 68342 1 47
2 68343 1 47
2 68344 1 47
2 68345 1 47
2 68346 1 47
2 68347 1 47
2 68348 1 47
2 68349 1 47
2 68350 1 47
2 68351 1 47
2 68352 1 47
2 68353 1 47
2 68354 1 47
2 68355 1 47
2 68356 1 47
2 68357 1 47
2 68358 1 47
2 68359 1 47
2 68360 1 47
2 68361 1 47
2 68362 1 47
2 68363 1 47
2 68364 1 47
2 68365 1 47
2 68366 1 47
2 68367 1 47
2 68368 1 47
2 68369 1 47
2 68370 1 47
2 68371 1 47
2 68372 1 47
2 68373 1 47
2 68374 1 47
2 68375 1 47
2 68376 1 47
2 68377 1 47
2 68378 1 47
2 68379 1 47
2 68380 1 47
2 68381 1 47
2 68382 1 47
2 68383 1 47
2 68384 1 47
2 68385 1 47
2 68386 1 47
2 68387 1 47
2 68388 1 47
2 68389 1 47
2 68390 1 47
2 68391 1 47
2 68392 1 47
2 68393 1 47
2 68394 1 47
2 68395 1 47
2 68396 1 47
2 68397 1 47
2 68398 1 47
2 68399 1 47
2 68400 1 47
2 68401 1 47
2 68402 1 47
2 68403 1 47
2 68404 1 47
2 68405 1 47
2 68406 1 47
2 68407 1 47
2 68408 1 47
2 68409 1 47
2 68410 1 47
2 68411 1 47
2 68412 1 47
2 68413 1 47
2 68414 1 47
2 68415 1 47
2 68416 1 47
2 68417 1 47
2 68418 1 47
2 68419 1 47
2 68420 1 47
2 68421 1 47
2 68422 1 47
2 68423 1 47
2 68424 1 47
2 68425 1 47
2 68426 1 47
2 68427 1 47
2 68428 1 47
2 68429 1 47
2 68430 1 47
2 68431 1 47
2 68432 1 47
2 68433 1 47
2 68434 1 47
2 68435 1 47
2 68436 1 47
2 68437 1 47
2 68438 1 47
2 68439 1 47
2 68440 1 47
2 68441 1 47
2 68442 1 47
2 68443 1 47
2 68444 1 47
2 68445 1 47
2 68446 1 47
2 68447 1 47
2 68448 1 47
2 68449 1 47
2 68450 1 47
2 68451 1 47
2 68452 1 47
2 68453 1 47
2 68454 1 47
2 68455 1 47
2 68456 1 47
2 68457 1 47
2 68458 1 47
2 68459 1 47
2 68460 1 47
2 68461 1 47
2 68462 1 47
2 68463 1 47
2 68464 1 47
2 68465 1 47
2 68466 1 47
2 68467 1 47
2 68468 1 47
2 68469 1 47
2 68470 1 47
2 68471 1 47
2 68472 1 47
2 68473 1 47
2 68474 1 47
2 68475 1 47
2 68476 1 47
2 68477 1 47
2 68478 1 47
2 68479 1 47
2 68480 1 47
2 68481 1 47
2 68482 1 47
2 68483 1 47
2 68484 1 47
2 68485 1 47
2 68486 1 47
2 68487 1 47
2 68488 1 47
2 68489 1 47
2 68490 1 47
2 68491 1 47
2 68492 1 47
2 68493 1 47
2 68494 1 47
2 68495 1 47
2 68496 1 47
2 68497 1 47
2 68498 1 47
2 68499 1 47
2 68500 1 47
2 68501 1 47
2 68502 1 47
2 68503 1 47
2 68504 1 47
2 68505 1 47
2 68506 1 47
2 68507 1 47
2 68508 1 47
2 68509 1 47
2 68510 1 47
2 68511 1 47
2 68512 1 47
2 68513 1 47
2 68514 1 47
2 68515 1 47
2 68516 1 47
2 68517 1 47
2 68518 1 47
2 68519 1 47
2 68520 1 47
2 68521 1 47
2 68522 1 47
2 68523 1 47
2 68524 1 47
2 68525 1 47
2 68526 1 47
2 68527 1 47
2 68528 1 47
2 68529 1 47
2 68530 1 47
2 68531 1 47
2 68532 1 47
2 68533 1 47
2 68534 1 47
2 68535 1 47
2 68536 1 47
2 68537 1 47
2 68538 1 47
2 68539 1 47
2 68540 1 47
2 68541 1 47
2 68542 1 47
2 68543 1 47
2 68544 1 47
2 68545 1 47
2 68546 1 47
2 68547 1 47
2 68548 1 47
2 68549 1 47
2 68550 1 47
2 68551 1 47
2 68552 1 47
2 68553 1 47
2 68554 1 47
2 68555 1 47
2 68556 1 47
2 68557 1 47
2 68558 1 47
2 68559 1 47
2 68560 1 47
2 68561 1 47
2 68562 1 47
2 68563 1 47
2 68564 1 47
2 68565 1 47
2 68566 1 47
2 68567 1 47
2 68568 1 47
2 68569 1 47
2 68570 1 47
2 68571 1 47
2 68572 1 47
2 68573 1 47
2 68574 1 47
2 68575 1 47
2 68576 1 47
2 68577 1 47
2 68578 1 47
2 68579 1 47
2 68580 1 47
2 68581 1 48
2 68582 1 48
2 68583 1 48
2 68584 1 48
2 68585 1 48
2 68586 1 48
2 68587 1 48
2 68588 1 48
2 68589 1 48
2 68590 1 48
2 68591 1 48
2 68592 1 48
2 68593 1 48
2 68594 1 48
2 68595 1 48
2 68596 1 48
2 68597 1 48
2 68598 1 48
2 68599 1 48
2 68600 1 48
2 68601 1 48
2 68602 1 48
2 68603 1 48
2 68604 1 48
2 68605 1 48
2 68606 1 48
2 68607 1 48
2 68608 1 48
2 68609 1 48
2 68610 1 48
2 68611 1 48
2 68612 1 48
2 68613 1 48
2 68614 1 48
2 68615 1 48
2 68616 1 48
2 68617 1 48
2 68618 1 48
2 68619 1 48
2 68620 1 48
2 68621 1 48
2 68622 1 48
2 68623 1 48
2 68624 1 48
2 68625 1 48
2 68626 1 48
2 68627 1 48
2 68628 1 48
2 68629 1 48
2 68630 1 48
2 68631 1 48
2 68632 1 48
2 68633 1 48
2 68634 1 48
2 68635 1 48
2 68636 1 48
2 68637 1 48
2 68638 1 48
2 68639 1 48
2 68640 1 48
2 68641 1 48
2 68642 1 48
2 68643 1 48
2 68644 1 48
2 68645 1 48
2 68646 1 48
2 68647 1 48
2 68648 1 48
2 68649 1 48
2 68650 1 48
2 68651 1 48
2 68652 1 48
2 68653 1 48
2 68654 1 48
2 68655 1 48
2 68656 1 48
2 68657 1 48
2 68658 1 48
2 68659 1 48
2 68660 1 48
2 68661 1 48
2 68662 1 48
2 68663 1 48
2 68664 1 48
2 68665 1 48
2 68666 1 48
2 68667 1 48
2 68668 1 48
2 68669 1 48
2 68670 1 48
2 68671 1 48
2 68672 1 48
2 68673 1 48
2 68674 1 48
2 68675 1 48
2 68676 1 48
2 68677 1 48
2 68678 1 48
2 68679 1 48
2 68680 1 48
2 68681 1 48
2 68682 1 48
2 68683 1 48
2 68684 1 48
2 68685 1 48
2 68686 1 48
2 68687 1 48
2 68688 1 48
2 68689 1 48
2 68690 1 48
2 68691 1 48
2 68692 1 48
2 68693 1 48
2 68694 1 48
2 68695 1 48
2 68696 1 48
2 68697 1 48
2 68698 1 48
2 68699 1 48
2 68700 1 48
2 68701 1 48
2 68702 1 48
2 68703 1 48
2 68704 1 48
2 68705 1 48
2 68706 1 48
2 68707 1 48
2 68708 1 48
2 68709 1 48
2 68710 1 48
2 68711 1 48
2 68712 1 48
2 68713 1 48
2 68714 1 48
2 68715 1 48
2 68716 1 48
2 68717 1 48
2 68718 1 48
2 68719 1 48
2 68720 1 48
2 68721 1 48
2 68722 1 48
2 68723 1 48
2 68724 1 48
2 68725 1 48
2 68726 1 48
2 68727 1 48
2 68728 1 48
2 68729 1 48
2 68730 1 48
2 68731 1 48
2 68732 1 48
2 68733 1 48
2 68734 1 48
2 68735 1 48
2 68736 1 48
2 68737 1 48
2 68738 1 48
2 68739 1 48
2 68740 1 48
2 68741 1 48
2 68742 1 48
2 68743 1 48
2 68744 1 48
2 68745 1 48
2 68746 1 48
2 68747 1 48
2 68748 1 48
2 68749 1 48
2 68750 1 48
2 68751 1 48
2 68752 1 48
2 68753 1 48
2 68754 1 48
2 68755 1 48
2 68756 1 48
2 68757 1 48
2 68758 1 48
2 68759 1 48
2 68760 1 48
2 68761 1 48
2 68762 1 48
2 68763 1 48
2 68764 1 48
2 68765 1 48
2 68766 1 48
2 68767 1 48
2 68768 1 48
2 68769 1 48
2 68770 1 48
2 68771 1 48
2 68772 1 48
2 68773 1 48
2 68774 1 48
2 68775 1 48
2 68776 1 48
2 68777 1 48
2 68778 1 48
2 68779 1 48
2 68780 1 48
2 68781 1 48
2 68782 1 48
2 68783 1 48
2 68784 1 48
2 68785 1 48
2 68786 1 48
2 68787 1 48
2 68788 1 48
2 68789 1 48
2 68790 1 48
2 68791 1 48
2 68792 1 48
2 68793 1 48
2 68794 1 48
2 68795 1 48
2 68796 1 48
2 68797 1 48
2 68798 1 48
2 68799 1 48
2 68800 1 48
2 68801 1 48
2 68802 1 48
2 68803 1 48
2 68804 1 48
2 68805 1 48
2 68806 1 48
2 68807 1 48
2 68808 1 48
2 68809 1 48
2 68810 1 48
2 68811 1 48
2 68812 1 48
2 68813 1 48
2 68814 1 48
2 68815 1 48
2 68816 1 48
2 68817 1 49
2 68818 1 49
2 68819 1 49
2 68820 1 49
2 68821 1 49
2 68822 1 49
2 68823 1 49
2 68824 1 49
2 68825 1 49
2 68826 1 49
2 68827 1 49
2 68828 1 49
2 68829 1 49
2 68830 1 49
2 68831 1 49
2 68832 1 49
2 68833 1 49
2 68834 1 49
2 68835 1 49
2 68836 1 49
2 68837 1 49
2 68838 1 49
2 68839 1 49
2 68840 1 49
2 68841 1 49
2 68842 1 49
2 68843 1 49
2 68844 1 49
2 68845 1 49
2 68846 1 49
2 68847 1 49
2 68848 1 49
2 68849 1 49
2 68850 1 49
2 68851 1 49
2 68852 1 49
2 68853 1 49
2 68854 1 49
2 68855 1 49
2 68856 1 49
2 68857 1 49
2 68858 1 49
2 68859 1 49
2 68860 1 49
2 68861 1 49
2 68862 1 49
2 68863 1 49
2 68864 1 49
2 68865 1 49
2 68866 1 49
2 68867 1 49
2 68868 1 49
2 68869 1 49
2 68870 1 49
2 68871 1 49
2 68872 1 49
2 68873 1 49
2 68874 1 49
2 68875 1 49
2 68876 1 49
2 68877 1 49
2 68878 1 49
2 68879 1 49
2 68880 1 49
2 68881 1 49
2 68882 1 49
2 68883 1 49
2 68884 1 49
2 68885 1 49
2 68886 1 49
2 68887 1 49
2 68888 1 49
2 68889 1 49
2 68890 1 49
2 68891 1 49
2 68892 1 49
2 68893 1 49
2 68894 1 49
2 68895 1 49
2 68896 1 49
2 68897 1 49
2 68898 1 49
2 68899 1 49
2 68900 1 49
2 68901 1 49
2 68902 1 49
2 68903 1 49
2 68904 1 49
2 68905 1 49
2 68906 1 49
2 68907 1 49
2 68908 1 49
2 68909 1 49
2 68910 1 49
2 68911 1 49
2 68912 1 49
2 68913 1 49
2 68914 1 49
2 68915 1 49
2 68916 1 49
2 68917 1 49
2 68918 1 49
2 68919 1 49
2 68920 1 49
2 68921 1 49
2 68922 1 49
2 68923 1 49
2 68924 1 49
2 68925 1 49
2 68926 1 49
2 68927 1 49
2 68928 1 49
2 68929 1 49
2 68930 1 49
2 68931 1 49
2 68932 1 49
2 68933 1 49
2 68934 1 49
2 68935 1 49
2 68936 1 49
2 68937 1 49
2 68938 1 49
2 68939 1 49
2 68940 1 49
2 68941 1 49
2 68942 1 49
2 68943 1 49
2 68944 1 49
2 68945 1 49
2 68946 1 49
2 68947 1 49
2 68948 1 49
2 68949 1 49
2 68950 1 49
2 68951 1 49
2 68952 1 49
2 68953 1 49
2 68954 1 49
2 68955 1 49
2 68956 1 49
2 68957 1 49
2 68958 1 49
2 68959 1 49
2 68960 1 49
2 68961 1 49
2 68962 1 49
2 68963 1 49
2 68964 1 49
2 68965 1 49
2 68966 1 49
2 68967 1 49
2 68968 1 49
2 68969 1 49
2 68970 1 49
2 68971 1 49
2 68972 1 49
2 68973 1 49
2 68974 1 49
2 68975 1 50
2 68976 1 50
2 68977 1 50
2 68978 1 50
2 68979 1 50
2 68980 1 50
2 68981 1 50
2 68982 1 50
2 68983 1 50
2 68984 1 50
2 68985 1 50
2 68986 1 50
2 68987 1 50
2 68988 1 50
2 68989 1 50
2 68990 1 50
2 68991 1 50
2 68992 1 50
2 68993 1 50
2 68994 1 50
2 68995 1 50
2 68996 1 50
2 68997 1 50
2 68998 1 50
2 68999 1 50
2 69000 1 50
2 69001 1 50
2 69002 1 50
2 69003 1 50
2 69004 1 50
2 69005 1 50
2 69006 1 50
2 69007 1 50
2 69008 1 50
2 69009 1 50
2 69010 1 50
2 69011 1 50
2 69012 1 50
2 69013 1 50
2 69014 1 50
2 69015 1 50
2 69016 1 50
2 69017 1 50
2 69018 1 50
2 69019 1 50
2 69020 1 50
2 69021 1 50
2 69022 1 50
2 69023 1 50
2 69024 1 50
2 69025 1 50
2 69026 1 50
2 69027 1 50
2 69028 1 50
2 69029 1 50
2 69030 1 50
2 69031 1 50
2 69032 1 50
2 69033 1 50
2 69034 1 50
2 69035 1 50
2 69036 1 50
2 69037 1 50
2 69038 1 50
2 69039 1 51
2 69040 1 51
2 69041 1 52
2 69042 1 52
2 69043 1 52
2 69044 1 52
2 69045 1 52
2 69046 1 52
2 69047 1 53
2 69048 1 53
2 69049 1 53
2 69050 1 53
2 69051 1 53
2 69052 1 53
2 69053 1 53
2 69054 1 53
2 69055 1 53
2 69056 1 53
2 69057 1 53
2 69058 1 53
2 69059 1 53
2 69060 1 53
2 69061 1 53
2 69062 1 53
2 69063 1 53
2 69064 1 53
2 69065 1 53
2 69066 1 53
2 69067 1 53
2 69068 1 53
2 69069 1 53
2 69070 1 53
2 69071 1 53
2 69072 1 53
2 69073 1 53
2 69074 1 53
2 69075 1 53
2 69076 1 53
2 69077 1 53
2 69078 1 54
2 69079 1 54
2 69080 1 54
2 69081 1 54
2 69082 1 54
2 69083 1 54
2 69084 1 54
2 69085 1 54
2 69086 1 54
2 69087 1 54
2 69088 1 54
2 69089 1 54
2 69090 1 54
2 69091 1 54
2 69092 1 54
2 69093 1 54
2 69094 1 54
2 69095 1 54
2 69096 1 54
2 69097 1 54
2 69098 1 54
2 69099 1 54
2 69100 1 54
2 69101 1 54
2 69102 1 54
2 69103 1 54
2 69104 1 54
2 69105 1 54
2 69106 1 54
2 69107 1 54
2 69108 1 54
2 69109 1 54
2 69110 1 54
2 69111 1 54
2 69112 1 54
2 69113 1 54
2 69114 1 54
2 69115 1 54
2 69116 1 54
2 69117 1 54
2 69118 1 54
2 69119 1 54
2 69120 1 54
2 69121 1 54
2 69122 1 54
2 69123 1 54
2 69124 1 54
2 69125 1 54
2 69126 1 54
2 69127 1 54
2 69128 1 54
2 69129 1 54
2 69130 1 54
2 69131 1 54
2 69132 1 54
2 69133 1 54
2 69134 1 54
2 69135 1 54
2 69136 1 54
2 69137 1 54
2 69138 1 54
2 69139 1 54
2 69140 1 54
2 69141 1 54
2 69142 1 54
2 69143 1 55
2 69144 1 55
2 69145 1 55
2 69146 1 55
2 69147 1 55
2 69148 1 56
2 69149 1 56
2 69150 1 56
2 69151 1 56
2 69152 1 56
2 69153 1 56
2 69154 1 56
2 69155 1 56
2 69156 1 56
2 69157 1 56
2 69158 1 56
2 69159 1 56
2 69160 1 56
2 69161 1 56
2 69162 1 56
2 69163 1 57
2 69164 1 57
2 69165 1 57
2 69166 1 57
2 69167 1 57
2 69168 1 57
2 69169 1 57
2 69170 1 57
2 69171 1 57
2 69172 1 57
2 69173 1 57
2 69174 1 57
2 69175 1 57
2 69176 1 57
2 69177 1 57
2 69178 1 57
2 69179 1 57
2 69180 1 57
2 69181 1 57
2 69182 1 57
2 69183 1 57
2 69184 1 57
2 69185 1 57
2 69186 1 57
2 69187 1 57
2 69188 1 57
2 69189 1 57
2 69190 1 57
2 69191 1 57
2 69192 1 57
2 69193 1 57
2 69194 1 57
2 69195 1 57
2 69196 1 57
2 69197 1 57
2 69198 1 57
2 69199 1 57
2 69200 1 57
2 69201 1 57
2 69202 1 57
2 69203 1 57
2 69204 1 57
2 69205 1 57
2 69206 1 57
2 69207 1 57
2 69208 1 57
2 69209 1 57
2 69210 1 57
2 69211 1 57
2 69212 1 57
2 69213 1 57
2 69214 1 57
2 69215 1 57
2 69216 1 57
2 69217 1 57
2 69218 1 57
2 69219 1 57
2 69220 1 58
2 69221 1 58
2 69222 1 58
2 69223 1 58
2 69224 1 58
2 69225 1 58
2 69226 1 58
2 69227 1 58
2 69228 1 58
2 69229 1 58
2 69230 1 58
2 69231 1 58
2 69232 1 58
2 69233 1 58
2 69234 1 58
2 69235 1 58
2 69236 1 58
2 69237 1 58
2 69238 1 58
2 69239 1 58
2 69240 1 58
2 69241 1 58
2 69242 1 58
2 69243 1 58
2 69244 1 58
2 69245 1 58
2 69246 1 58
2 69247 1 58
2 69248 1 58
2 69249 1 58
2 69250 1 58
2 69251 1 58
2 69252 1 58
2 69253 1 58
2 69254 1 58
2 69255 1 58
2 69256 1 58
2 69257 1 58
2 69258 1 58
2 69259 1 58
2 69260 1 58
2 69261 1 58
2 69262 1 58
2 69263 1 58
2 69264 1 58
2 69265 1 58
2 69266 1 58
2 69267 1 58
2 69268 1 58
2 69269 1 58
2 69270 1 58
2 69271 1 58
2 69272 1 58
2 69273 1 58
2 69274 1 58
2 69275 1 58
2 69276 1 58
2 69277 1 58
2 69278 1 58
2 69279 1 58
2 69280 1 58
2 69281 1 58
2 69282 1 58
2 69283 1 58
2 69284 1 58
2 69285 1 58
2 69286 1 59
2 69287 1 59
2 69288 1 59
2 69289 1 59
2 69290 1 59
2 69291 1 60
2 69292 1 60
2 69293 1 60
2 69294 1 60
2 69295 1 60
2 69296 1 60
2 69297 1 60
2 69298 1 60
2 69299 1 60
2 69300 1 60
2 69301 1 60
2 69302 1 60
2 69303 1 60
2 69304 1 60
2 69305 1 60
2 69306 1 60
2 69307 1 60
2 69308 1 60
2 69309 1 60
2 69310 1 60
2 69311 1 60
2 69312 1 60
2 69313 1 60
2 69314 1 60
2 69315 1 60
2 69316 1 60
2 69317 1 60
2 69318 1 60
2 69319 1 60
2 69320 1 60
2 69321 1 60
2 69322 1 60
2 69323 1 60
2 69324 1 60
2 69325 1 60
2 69326 1 60
2 69327 1 61
2 69328 1 61
2 69329 1 61
2 69330 1 61
2 69331 1 62
2 69332 1 62
2 69333 1 64
2 69334 1 64
2 69335 1 68
2 69336 1 68
2 69337 1 69
2 69338 1 69
2 69339 1 69
2 69340 1 69
2 69341 1 69
2 69342 1 69
2 69343 1 69
2 69344 1 69
2 69345 1 69
2 69346 1 69
2 69347 1 70
2 69348 1 70
2 69349 1 70
2 69350 1 70
2 69351 1 70
2 69352 1 70
2 69353 1 72
2 69354 1 72
2 69355 1 72
2 69356 1 73
2 69357 1 73
2 69358 1 73
2 69359 1 73
2 69360 1 73
2 69361 1 73
2 69362 1 73
2 69363 1 73
2 69364 1 73
2 69365 1 73
2 69366 1 73
2 69367 1 73
2 69368 1 73
2 69369 1 73
2 69370 1 73
2 69371 1 73
2 69372 1 73
2 69373 1 73
2 69374 1 73
2 69375 1 73
2 69376 1 73
2 69377 1 73
2 69378 1 73
2 69379 1 73
2 69380 1 73
2 69381 1 73
2 69382 1 74
2 69383 1 74
2 69384 1 74
2 69385 1 74
2 69386 1 74
2 69387 1 74
2 69388 1 74
2 69389 1 74
2 69390 1 74
2 69391 1 74
2 69392 1 74
2 69393 1 74
2 69394 1 74
2 69395 1 74
2 69396 1 74
2 69397 1 74
2 69398 1 74
2 69399 1 74
2 69400 1 74
2 69401 1 74
2 69402 1 74
2 69403 1 74
2 69404 1 74
2 69405 1 74
2 69406 1 74
2 69407 1 74
2 69408 1 74
2 69409 1 74
2 69410 1 74
2 69411 1 74
2 69412 1 74
2 69413 1 74
2 69414 1 74
2 69415 1 74
2 69416 1 74
2 69417 1 74
2 69418 1 74
2 69419 1 74
2 69420 1 74
2 69421 1 74
2 69422 1 74
2 69423 1 74
2 69424 1 74
2 69425 1 74
2 69426 1 74
2 69427 1 74
2 69428 1 74
2 69429 1 74
2 69430 1 74
2 69431 1 74
2 69432 1 74
2 69433 1 74
2 69434 1 74
2 69435 1 74
2 69436 1 74
2 69437 1 74
2 69438 1 74
2 69439 1 76
2 69440 1 76
2 69441 1 76
2 69442 1 76
2 69443 1 76
2 69444 1 76
2 69445 1 76
2 69446 1 76
2 69447 1 76
2 69448 1 77
2 69449 1 77
2 69450 1 78
2 69451 1 78
2 69452 1 78
2 69453 1 78
2 69454 1 78
2 69455 1 78
2 69456 1 78
2 69457 1 85
2 69458 1 85
2 69459 1 85
2 69460 1 85
2 69461 1 85
2 69462 1 85
2 69463 1 85
2 69464 1 85
2 69465 1 85
2 69466 1 85
2 69467 1 85
2 69468 1 86
2 69469 1 86
2 69470 1 86
2 69471 1 86
2 69472 1 86
2 69473 1 86
2 69474 1 87
2 69475 1 87
2 69476 1 87
2 69477 1 87
2 69478 1 87
2 69479 1 87
2 69480 1 87
2 69481 1 87
2 69482 1 87
2 69483 1 87
2 69484 1 87
2 69485 1 87
2 69486 1 87
2 69487 1 87
2 69488 1 87
2 69489 1 87
2 69490 1 87
2 69491 1 87
2 69492 1 87
2 69493 1 87
2 69494 1 87
2 69495 1 87
2 69496 1 87
2 69497 1 87
2 69498 1 87
2 69499 1 87
2 69500 1 87
2 69501 1 87
2 69502 1 87
2 69503 1 87
2 69504 1 87
2 69505 1 87
2 69506 1 87
2 69507 1 87
2 69508 1 87
2 69509 1 87
2 69510 1 87
2 69511 1 87
2 69512 1 87
2 69513 1 87
2 69514 1 87
2 69515 1 87
2 69516 1 87
2 69517 1 87
2 69518 1 87
2 69519 1 87
2 69520 1 87
2 69521 1 87
2 69522 1 87
2 69523 1 87
2 69524 1 87
2 69525 1 87
2 69526 1 87
2 69527 1 87
2 69528 1 87
2 69529 1 87
2 69530 1 87
2 69531 1 87
2 69532 1 87
2 69533 1 87
2 69534 1 87
2 69535 1 87
2 69536 1 87
2 69537 1 87
2 69538 1 87
2 69539 1 87
2 69540 1 87
2 69541 1 87
2 69542 1 87
2 69543 1 87
2 69544 1 87
2 69545 1 87
2 69546 1 87
2 69547 1 87
2 69548 1 87
2 69549 1 87
2 69550 1 87
2 69551 1 87
2 69552 1 87
2 69553 1 87
2 69554 1 87
2 69555 1 87
2 69556 1 87
2 69557 1 87
2 69558 1 87
2 69559 1 87
2 69560 1 87
2 69561 1 87
2 69562 1 87
2 69563 1 87
2 69564 1 87
2 69565 1 87
2 69566 1 87
2 69567 1 87
2 69568 1 87
2 69569 1 87
2 69570 1 87
2 69571 1 87
2 69572 1 87
2 69573 1 87
2 69574 1 87
2 69575 1 87
2 69576 1 87
2 69577 1 87
2 69578 1 87
2 69579 1 87
2 69580 1 87
2 69581 1 87
2 69582 1 87
2 69583 1 87
2 69584 1 87
2 69585 1 87
2 69586 1 87
2 69587 1 87
2 69588 1 87
2 69589 1 87
2 69590 1 87
2 69591 1 87
2 69592 1 87
2 69593 1 87
2 69594 1 87
2 69595 1 87
2 69596 1 87
2 69597 1 87
2 69598 1 87
2 69599 1 87
2 69600 1 87
2 69601 1 87
2 69602 1 87
2 69603 1 87
2 69604 1 87
2 69605 1 87
2 69606 1 87
2 69607 1 87
2 69608 1 87
2 69609 1 87
2 69610 1 87
2 69611 1 87
2 69612 1 87
2 69613 1 87
2 69614 1 87
2 69615 1 87
2 69616 1 87
2 69617 1 87
2 69618 1 87
2 69619 1 87
2 69620 1 87
2 69621 1 88
2 69622 1 88
2 69623 1 88
2 69624 1 88
2 69625 1 88
2 69626 1 88
2 69627 1 88
2 69628 1 88
2 69629 1 88
2 69630 1 88
2 69631 1 88
2 69632 1 88
2 69633 1 88
2 69634 1 88
2 69635 1 88
2 69636 1 88
2 69637 1 88
2 69638 1 88
2 69639 1 88
2 69640 1 88
2 69641 1 88
2 69642 1 88
2 69643 1 88
2 69644 1 88
2 69645 1 88
2 69646 1 88
2 69647 1 88
2 69648 1 88
2 69649 1 88
2 69650 1 88
2 69651 1 88
2 69652 1 88
2 69653 1 88
2 69654 1 88
2 69655 1 88
2 69656 1 88
2 69657 1 88
2 69658 1 88
2 69659 1 88
2 69660 1 88
2 69661 1 88
2 69662 1 88
2 69663 1 88
2 69664 1 88
2 69665 1 88
2 69666 1 88
2 69667 1 88
2 69668 1 88
2 69669 1 88
2 69670 1 88
2 69671 1 88
2 69672 1 88
2 69673 1 88
2 69674 1 88
2 69675 1 88
2 69676 1 88
2 69677 1 88
2 69678 1 88
2 69679 1 88
2 69680 1 88
2 69681 1 88
2 69682 1 88
2 69683 1 88
2 69684 1 88
2 69685 1 88
2 69686 1 88
2 69687 1 88
2 69688 1 88
2 69689 1 88
2 69690 1 88
2 69691 1 88
2 69692 1 88
2 69693 1 88
2 69694 1 88
2 69695 1 88
2 69696 1 88
2 69697 1 88
2 69698 1 88
2 69699 1 88
2 69700 1 88
2 69701 1 88
2 69702 1 88
2 69703 1 88
2 69704 1 88
2 69705 1 88
2 69706 1 88
2 69707 1 88
2 69708 1 88
2 69709 1 88
2 69710 1 88
2 69711 1 88
2 69712 1 88
2 69713 1 88
2 69714 1 88
2 69715 1 88
2 69716 1 89
2 69717 1 89
2 69718 1 89
2 69719 1 89
2 69720 1 89
2 69721 1 89
2 69722 1 89
2 69723 1 89
2 69724 1 89
2 69725 1 89
2 69726 1 89
2 69727 1 89
2 69728 1 89
2 69729 1 89
2 69730 1 89
2 69731 1 90
2 69732 1 90
2 69733 1 90
2 69734 1 90
2 69735 1 90
2 69736 1 90
2 69737 1 90
2 69738 1 90
2 69739 1 90
2 69740 1 90
2 69741 1 91
2 69742 1 91
2 69743 1 91
2 69744 1 91
2 69745 1 91
2 69746 1 91
2 69747 1 91
2 69748 1 91
2 69749 1 91
2 69750 1 91
2 69751 1 91
2 69752 1 91
2 69753 1 91
2 69754 1 91
2 69755 1 91
2 69756 1 91
2 69757 1 91
2 69758 1 91
2 69759 1 91
2 69760 1 91
2 69761 1 91
2 69762 1 91
2 69763 1 91
2 69764 1 91
2 69765 1 91
2 69766 1 91
2 69767 1 91
2 69768 1 91
2 69769 1 91
2 69770 1 91
2 69771 1 91
2 69772 1 91
2 69773 1 91
2 69774 1 91
2 69775 1 91
2 69776 1 91
2 69777 1 91
2 69778 1 91
2 69779 1 91
2 69780 1 91
2 69781 1 91
2 69782 1 91
2 69783 1 91
2 69784 1 91
2 69785 1 91
2 69786 1 91
2 69787 1 91
2 69788 1 91
2 69789 1 91
2 69790 1 91
2 69791 1 91
2 69792 1 91
2 69793 1 91
2 69794 1 91
2 69795 1 91
2 69796 1 91
2 69797 1 91
2 69798 1 91
2 69799 1 91
2 69800 1 91
2 69801 1 91
2 69802 1 91
2 69803 1 91
2 69804 1 91
2 69805 1 91
2 69806 1 91
2 69807 1 91
2 69808 1 91
2 69809 1 91
2 69810 1 91
2 69811 1 91
2 69812 1 91
2 69813 1 91
2 69814 1 91
2 69815 1 91
2 69816 1 91
2 69817 1 91
2 69818 1 91
2 69819 1 91
2 69820 1 91
2 69821 1 91
2 69822 1 91
2 69823 1 91
2 69824 1 91
2 69825 1 91
2 69826 1 91
2 69827 1 91
2 69828 1 91
2 69829 1 91
2 69830 1 91
2 69831 1 91
2 69832 1 91
2 69833 1 91
2 69834 1 91
2 69835 1 91
2 69836 1 91
2 69837 1 91
2 69838 1 91
2 69839 1 91
2 69840 1 91
2 69841 1 91
2 69842 1 91
2 69843 1 91
2 69844 1 91
2 69845 1 91
2 69846 1 91
2 69847 1 91
2 69848 1 91
2 69849 1 91
2 69850 1 91
2 69851 1 91
2 69852 1 91
2 69853 1 91
2 69854 1 91
2 69855 1 91
2 69856 1 91
2 69857 1 91
2 69858 1 91
2 69859 1 91
2 69860 1 91
2 69861 1 91
2 69862 1 91
2 69863 1 91
2 69864 1 92
2 69865 1 92
2 69866 1 92
2 69867 1 92
2 69868 1 92
2 69869 1 92
2 69870 1 92
2 69871 1 92
2 69872 1 92
2 69873 1 92
2 69874 1 92
2 69875 1 92
2 69876 1 92
2 69877 1 92
2 69878 1 92
2 69879 1 92
2 69880 1 92
2 69881 1 92
2 69882 1 92
2 69883 1 92
2 69884 1 92
2 69885 1 92
2 69886 1 92
2 69887 1 92
2 69888 1 92
2 69889 1 92
2 69890 1 92
2 69891 1 92
2 69892 1 92
2 69893 1 92
2 69894 1 92
2 69895 1 92
2 69896 1 92
2 69897 1 92
2 69898 1 92
2 69899 1 92
2 69900 1 92
2 69901 1 92
2 69902 1 92
2 69903 1 92
2 69904 1 92
2 69905 1 92
2 69906 1 92
2 69907 1 92
2 69908 1 92
2 69909 1 92
2 69910 1 92
2 69911 1 92
2 69912 1 92
2 69913 1 92
2 69914 1 92
2 69915 1 92
2 69916 1 92
2 69917 1 92
2 69918 1 92
2 69919 1 92
2 69920 1 92
2 69921 1 92
2 69922 1 92
2 69923 1 92
2 69924 1 92
2 69925 1 92
2 69926 1 92
2 69927 1 92
2 69928 1 92
2 69929 1 92
2 69930 1 92
2 69931 1 92
2 69932 1 92
2 69933 1 92
2 69934 1 92
2 69935 1 92
2 69936 1 92
2 69937 1 92
2 69938 1 92
2 69939 1 92
2 69940 1 92
2 69941 1 92
2 69942 1 92
2 69943 1 92
2 69944 1 92
2 69945 1 92
2 69946 1 92
2 69947 1 92
2 69948 1 92
2 69949 1 92
2 69950 1 92
2 69951 1 92
2 69952 1 92
2 69953 1 92
2 69954 1 92
2 69955 1 92
2 69956 1 92
2 69957 1 92
2 69958 1 92
2 69959 1 92
2 69960 1 92
2 69961 1 92
2 69962 1 92
2 69963 1 92
2 69964 1 92
2 69965 1 92
2 69966 1 92
2 69967 1 93
2 69968 1 93
2 69969 1 93
2 69970 1 93
2 69971 1 93
2 69972 1 93
2 69973 1 93
2 69974 1 94
2 69975 1 94
2 69976 1 94
2 69977 1 94
2 69978 1 94
2 69979 1 94
2 69980 1 94
2 69981 1 94
2 69982 1 94
2 69983 1 94
2 69984 1 94
2 69985 1 94
2 69986 1 94
2 69987 1 94
2 69988 1 94
2 69989 1 94
2 69990 1 94
2 69991 1 94
2 69992 1 94
2 69993 1 94
2 69994 1 94
2 69995 1 94
2 69996 1 94
2 69997 1 94
2 69998 1 94
2 69999 1 94
2 70000 1 95
2 70001 1 95
2 70002 1 95
2 70003 1 95
2 70004 1 96
2 70005 1 96
2 70006 1 101
2 70007 1 101
2 70008 1 101
2 70009 1 101
2 70010 1 101
2 70011 1 101
2 70012 1 101
2 70013 1 101
2 70014 1 101
2 70015 1 101
2 70016 1 101
2 70017 1 101
2 70018 1 101
2 70019 1 101
2 70020 1 101
2 70021 1 101
2 70022 1 101
2 70023 1 101
2 70024 1 101
2 70025 1 101
2 70026 1 101
2 70027 1 101
2 70028 1 101
2 70029 1 101
2 70030 1 101
2 70031 1 101
2 70032 1 101
2 70033 1 101
2 70034 1 101
2 70035 1 101
2 70036 1 101
2 70037 1 101
2 70038 1 101
2 70039 1 101
2 70040 1 101
2 70041 1 101
2 70042 1 101
2 70043 1 101
2 70044 1 101
2 70045 1 101
2 70046 1 101
2 70047 1 101
2 70048 1 101
2 70049 1 101
2 70050 1 101
2 70051 1 101
2 70052 1 101
2 70053 1 101
2 70054 1 101
2 70055 1 101
2 70056 1 101
2 70057 1 101
2 70058 1 101
2 70059 1 101
2 70060 1 101
2 70061 1 101
2 70062 1 101
2 70063 1 101
2 70064 1 101
2 70065 1 101
2 70066 1 101
2 70067 1 101
2 70068 1 101
2 70069 1 101
2 70070 1 101
2 70071 1 101
2 70072 1 101
2 70073 1 101
2 70074 1 101
2 70075 1 101
2 70076 1 101
2 70077 1 101
2 70078 1 101
2 70079 1 101
2 70080 1 101
2 70081 1 101
2 70082 1 101
2 70083 1 101
2 70084 1 101
2 70085 1 101
2 70086 1 101
2 70087 1 101
2 70088 1 101
2 70089 1 101
2 70090 1 101
2 70091 1 101
2 70092 1 101
2 70093 1 101
2 70094 1 101
2 70095 1 101
2 70096 1 101
2 70097 1 101
2 70098 1 102
2 70099 1 102
2 70100 1 102
2 70101 1 102
2 70102 1 102
2 70103 1 102
2 70104 1 102
2 70105 1 102
2 70106 1 102
2 70107 1 102
2 70108 1 102
2 70109 1 102
2 70110 1 102
2 70111 1 102
2 70112 1 102
2 70113 1 102
2 70114 1 102
2 70115 1 102
2 70116 1 102
2 70117 1 102
2 70118 1 102
2 70119 1 102
2 70120 1 102
2 70121 1 102
2 70122 1 102
2 70123 1 102
2 70124 1 102
2 70125 1 102
2 70126 1 102
2 70127 1 102
2 70128 1 102
2 70129 1 102
2 70130 1 102
2 70131 1 102
2 70132 1 102
2 70133 1 102
2 70134 1 102
2 70135 1 102
2 70136 1 102
2 70137 1 102
2 70138 1 102
2 70139 1 102
2 70140 1 102
2 70141 1 102
2 70142 1 102
2 70143 1 102
2 70144 1 102
2 70145 1 102
2 70146 1 102
2 70147 1 102
2 70148 1 102
2 70149 1 102
2 70150 1 102
2 70151 1 102
2 70152 1 102
2 70153 1 102
2 70154 1 102
2 70155 1 102
2 70156 1 102
2 70157 1 102
2 70158 1 102
2 70159 1 102
2 70160 1 102
2 70161 1 102
2 70162 1 102
2 70163 1 102
2 70164 1 102
2 70165 1 102
2 70166 1 102
2 70167 1 102
2 70168 1 102
2 70169 1 102
2 70170 1 102
2 70171 1 102
2 70172 1 102
2 70173 1 102
2 70174 1 102
2 70175 1 102
2 70176 1 102
2 70177 1 102
2 70178 1 102
2 70179 1 102
2 70180 1 102
2 70181 1 102
2 70182 1 102
2 70183 1 102
2 70184 1 102
2 70185 1 102
2 70186 1 102
2 70187 1 102
2 70188 1 102
2 70189 1 102
2 70190 1 102
2 70191 1 102
2 70192 1 102
2 70193 1 102
2 70194 1 102
2 70195 1 102
2 70196 1 102
2 70197 1 102
2 70198 1 102
2 70199 1 102
2 70200 1 102
2 70201 1 102
2 70202 1 102
2 70203 1 102
2 70204 1 102
2 70205 1 102
2 70206 1 102
2 70207 1 102
2 70208 1 102
2 70209 1 102
2 70210 1 102
2 70211 1 102
2 70212 1 102
2 70213 1 102
2 70214 1 102
2 70215 1 102
2 70216 1 102
2 70217 1 102
2 70218 1 102
2 70219 1 102
2 70220 1 102
2 70221 1 103
2 70222 1 103
2 70223 1 103
2 70224 1 103
2 70225 1 103
2 70226 1 103
2 70227 1 103
2 70228 1 103
2 70229 1 103
2 70230 1 103
2 70231 1 103
2 70232 1 103
2 70233 1 103
2 70234 1 103
2 70235 1 103
2 70236 1 103
2 70237 1 103
2 70238 1 104
2 70239 1 104
2 70240 1 104
2 70241 1 104
2 70242 1 105
2 70243 1 105
2 70244 1 105
2 70245 1 105
2 70246 1 105
2 70247 1 105
2 70248 1 106
2 70249 1 106
2 70250 1 107
2 70251 1 107
2 70252 1 107
2 70253 1 107
2 70254 1 107
2 70255 1 107
2 70256 1 107
2 70257 1 107
2 70258 1 108
2 70259 1 108
2 70260 1 108
2 70261 1 108
2 70262 1 108
2 70263 1 108
2 70264 1 108
2 70265 1 108
2 70266 1 111
2 70267 1 111
2 70268 1 111
2 70269 1 111
2 70270 1 111
2 70271 1 111
2 70272 1 111
2 70273 1 111
2 70274 1 111
2 70275 1 111
2 70276 1 111
2 70277 1 111
2 70278 1 111
2 70279 1 111
2 70280 1 111
2 70281 1 111
2 70282 1 111
2 70283 1 111
2 70284 1 111
2 70285 1 111
2 70286 1 111
2 70287 1 111
2 70288 1 111
2 70289 1 111
2 70290 1 111
2 70291 1 111
2 70292 1 111
2 70293 1 111
2 70294 1 111
2 70295 1 111
2 70296 1 112
2 70297 1 112
2 70298 1 112
2 70299 1 112
2 70300 1 112
2 70301 1 112
2 70302 1 112
2 70303 1 112
2 70304 1 112
2 70305 1 112
2 70306 1 112
2 70307 1 112
2 70308 1 112
2 70309 1 112
2 70310 1 112
2 70311 1 112
2 70312 1 112
2 70313 1 112
2 70314 1 112
2 70315 1 112
2 70316 1 112
2 70317 1 112
2 70318 1 112
2 70319 1 112
2 70320 1 112
2 70321 1 112
2 70322 1 112
2 70323 1 112
2 70324 1 112
2 70325 1 112
2 70326 1 112
2 70327 1 112
2 70328 1 112
2 70329 1 112
2 70330 1 112
2 70331 1 112
2 70332 1 112
2 70333 1 112
2 70334 1 112
2 70335 1 112
2 70336 1 112
2 70337 1 112
2 70338 1 112
2 70339 1 112
2 70340 1 112
2 70341 1 112
2 70342 1 112
2 70343 1 112
2 70344 1 112
2 70345 1 112
2 70346 1 112
2 70347 1 112
2 70348 1 112
2 70349 1 112
2 70350 1 112
2 70351 1 112
2 70352 1 112
2 70353 1 115
2 70354 1 115
2 70355 1 115
2 70356 1 116
2 70357 1 116
2 70358 1 116
2 70359 1 118
2 70360 1 118
2 70361 1 119
2 70362 1 119
2 70363 1 119
2 70364 1 120
2 70365 1 120
2 70366 1 120
2 70367 1 120
2 70368 1 120
2 70369 1 120
2 70370 1 120
2 70371 1 120
2 70372 1 120
2 70373 1 120
2 70374 1 120
2 70375 1 120
2 70376 1 120
2 70377 1 120
2 70378 1 120
2 70379 1 120
2 70380 1 120
2 70381 1 120
2 70382 1 120
2 70383 1 120
2 70384 1 122
2 70385 1 122
2 70386 1 123
2 70387 1 123
2 70388 1 124
2 70389 1 124
2 70390 1 124
2 70391 1 124
2 70392 1 125
2 70393 1 125
2 70394 1 125
2 70395 1 125
2 70396 1 125
2 70397 1 125
2 70398 1 125
2 70399 1 125
2 70400 1 125
2 70401 1 126
2 70402 1 126
2 70403 1 126
2 70404 1 126
2 70405 1 126
2 70406 1 126
2 70407 1 126
2 70408 1 126
2 70409 1 126
2 70410 1 126
2 70411 1 126
2 70412 1 129
2 70413 1 129
2 70414 1 129
2 70415 1 129
2 70416 1 129
2 70417 1 132
2 70418 1 132
2 70419 1 132
2 70420 1 132
2 70421 1 132
2 70422 1 134
2 70423 1 134
2 70424 1 135
2 70425 1 135
2 70426 1 135
2 70427 1 136
2 70428 1 136
2 70429 1 136
2 70430 1 138
2 70431 1 138
2 70432 1 139
2 70433 1 139
2 70434 1 139
2 70435 1 139
2 70436 1 140
2 70437 1 140
2 70438 1 141
2 70439 1 141
2 70440 1 141
2 70441 1 141
2 70442 1 141
2 70443 1 141
2 70444 1 141
2 70445 1 141
2 70446 1 141
2 70447 1 141
2 70448 1 141
2 70449 1 141
2 70450 1 141
2 70451 1 141
2 70452 1 141
2 70453 1 141
2 70454 1 141
2 70455 1 141
2 70456 1 141
2 70457 1 141
2 70458 1 141
2 70459 1 142
2 70460 1 142
2 70461 1 142
2 70462 1 142
2 70463 1 142
2 70464 1 142
2 70465 1 142
2 70466 1 142
2 70467 1 143
2 70468 1 143
2 70469 1 143
2 70470 1 143
2 70471 1 143
2 70472 1 143
2 70473 1 143
2 70474 1 143
2 70475 1 143
2 70476 1 143
2 70477 1 143
2 70478 1 143
2 70479 1 143
2 70480 1 143
2 70481 1 143
2 70482 1 143
2 70483 1 143
2 70484 1 143
2 70485 1 143
2 70486 1 143
2 70487 1 143
2 70488 1 143
2 70489 1 143
2 70490 1 143
2 70491 1 143
2 70492 1 143
2 70493 1 143
2 70494 1 143
2 70495 1 143
2 70496 1 143
2 70497 1 143
2 70498 1 143
2 70499 1 143
2 70500 1 143
2 70501 1 143
2 70502 1 143
2 70503 1 143
2 70504 1 143
2 70505 1 144
2 70506 1 144
2 70507 1 144
2 70508 1 144
2 70509 1 144
2 70510 1 144
2 70511 1 144
2 70512 1 144
2 70513 1 144
2 70514 1 144
2 70515 1 144
2 70516 1 144
2 70517 1 144
2 70518 1 144
2 70519 1 144
2 70520 1 144
2 70521 1 144
2 70522 1 144
2 70523 1 144
2 70524 1 144
2 70525 1 144
2 70526 1 144
2 70527 1 144
2 70528 1 144
2 70529 1 144
2 70530 1 144
2 70531 1 144
2 70532 1 144
2 70533 1 144
2 70534 1 144
2 70535 1 144
2 70536 1 144
2 70537 1 144
2 70538 1 144
2 70539 1 144
2 70540 1 144
2 70541 1 144
2 70542 1 144
2 70543 1 144
2 70544 1 144
2 70545 1 144
2 70546 1 145
2 70547 1 145
2 70548 1 145
2 70549 1 145
2 70550 1 147
2 70551 1 147
2 70552 1 150
2 70553 1 150
2 70554 1 150
2 70555 1 150
2 70556 1 150
2 70557 1 155
2 70558 1 155
2 70559 1 155
2 70560 1 155
2 70561 1 155
2 70562 1 155
2 70563 1 155
2 70564 1 155
2 70565 1 155
2 70566 1 155
2 70567 1 155
2 70568 1 155
2 70569 1 155
2 70570 1 155
2 70571 1 155
2 70572 1 155
2 70573 1 155
2 70574 1 155
2 70575 1 155
2 70576 1 155
2 70577 1 155
2 70578 1 155
2 70579 1 155
2 70580 1 155
2 70581 1 155
2 70582 1 155
2 70583 1 155
2 70584 1 155
2 70585 1 155
2 70586 1 155
2 70587 1 155
2 70588 1 155
2 70589 1 155
2 70590 1 155
2 70591 1 155
2 70592 1 155
2 70593 1 155
2 70594 1 155
2 70595 1 155
2 70596 1 155
2 70597 1 155
2 70598 1 155
2 70599 1 155
2 70600 1 155
2 70601 1 155
2 70602 1 155
2 70603 1 155
2 70604 1 155
2 70605 1 155
2 70606 1 155
2 70607 1 155
2 70608 1 155
2 70609 1 155
2 70610 1 155
2 70611 1 155
2 70612 1 155
2 70613 1 155
2 70614 1 155
2 70615 1 155
2 70616 1 155
2 70617 1 155
2 70618 1 155
2 70619 1 155
2 70620 1 155
2 70621 1 155
2 70622 1 155
2 70623 1 155
2 70624 1 155
2 70625 1 155
2 70626 1 155
2 70627 1 155
2 70628 1 155
2 70629 1 155
2 70630 1 155
2 70631 1 155
2 70632 1 155
2 70633 1 155
2 70634 1 155
2 70635 1 155
2 70636 1 155
2 70637 1 155
2 70638 1 155
2 70639 1 155
2 70640 1 155
2 70641 1 155
2 70642 1 155
2 70643 1 155
2 70644 1 155
2 70645 1 155
2 70646 1 155
2 70647 1 155
2 70648 1 155
2 70649 1 155
2 70650 1 155
2 70651 1 155
2 70652 1 155
2 70653 1 155
2 70654 1 155
2 70655 1 155
2 70656 1 155
2 70657 1 155
2 70658 1 155
2 70659 1 155
2 70660 1 155
2 70661 1 155
2 70662 1 155
2 70663 1 155
2 70664 1 155
2 70665 1 155
2 70666 1 155
2 70667 1 155
2 70668 1 155
2 70669 1 155
2 70670 1 155
2 70671 1 155
2 70672 1 155
2 70673 1 155
2 70674 1 155
2 70675 1 155
2 70676 1 155
2 70677 1 155
2 70678 1 155
2 70679 1 155
2 70680 1 155
2 70681 1 155
2 70682 1 155
2 70683 1 155
2 70684 1 155
2 70685 1 155
2 70686 1 155
2 70687 1 155
2 70688 1 155
2 70689 1 155
2 70690 1 155
2 70691 1 155
2 70692 1 155
2 70693 1 155
2 70694 1 155
2 70695 1 155
2 70696 1 155
2 70697 1 155
2 70698 1 155
2 70699 1 155
2 70700 1 155
2 70701 1 155
2 70702 1 155
2 70703 1 155
2 70704 1 155
2 70705 1 155
2 70706 1 155
2 70707 1 155
2 70708 1 155
2 70709 1 155
2 70710 1 155
2 70711 1 155
2 70712 1 155
2 70713 1 155
2 70714 1 155
2 70715 1 156
2 70716 1 156
2 70717 1 156
2 70718 1 156
2 70719 1 156
2 70720 1 156
2 70721 1 156
2 70722 1 156
2 70723 1 156
2 70724 1 156
2 70725 1 156
2 70726 1 156
2 70727 1 156
2 70728 1 156
2 70729 1 156
2 70730 1 156
2 70731 1 156
2 70732 1 156
2 70733 1 156
2 70734 1 156
2 70735 1 156
2 70736 1 156
2 70737 1 156
2 70738 1 156
2 70739 1 156
2 70740 1 156
2 70741 1 156
2 70742 1 156
2 70743 1 156
2 70744 1 156
2 70745 1 156
2 70746 1 156
2 70747 1 156
2 70748 1 156
2 70749 1 156
2 70750 1 156
2 70751 1 156
2 70752 1 156
2 70753 1 156
2 70754 1 156
2 70755 1 156
2 70756 1 156
2 70757 1 156
2 70758 1 156
2 70759 1 156
2 70760 1 156
2 70761 1 156
2 70762 1 156
2 70763 1 156
2 70764 1 156
2 70765 1 156
2 70766 1 156
2 70767 1 156
2 70768 1 156
2 70769 1 156
2 70770 1 156
2 70771 1 156
2 70772 1 156
2 70773 1 156
2 70774 1 156
2 70775 1 156
2 70776 1 156
2 70777 1 156
2 70778 1 156
2 70779 1 156
2 70780 1 156
2 70781 1 156
2 70782 1 156
2 70783 1 156
2 70784 1 156
2 70785 1 156
2 70786 1 156
2 70787 1 156
2 70788 1 156
2 70789 1 156
2 70790 1 156
2 70791 1 156
2 70792 1 156
2 70793 1 156
2 70794 1 156
2 70795 1 156
2 70796 1 156
2 70797 1 156
2 70798 1 156
2 70799 1 156
2 70800 1 156
2 70801 1 156
2 70802 1 156
2 70803 1 156
2 70804 1 156
2 70805 1 156
2 70806 1 156
2 70807 1 156
2 70808 1 156
2 70809 1 156
2 70810 1 156
2 70811 1 156
2 70812 1 156
2 70813 1 156
2 70814 1 156
2 70815 1 156
2 70816 1 156
2 70817 1 156
2 70818 1 156
2 70819 1 156
2 70820 1 156
2 70821 1 156
2 70822 1 156
2 70823 1 156
2 70824 1 156
2 70825 1 156
2 70826 1 156
2 70827 1 156
2 70828 1 156
2 70829 1 156
2 70830 1 156
2 70831 1 156
2 70832 1 156
2 70833 1 156
2 70834 1 156
2 70835 1 156
2 70836 1 156
2 70837 1 156
2 70838 1 156
2 70839 1 156
2 70840 1 156
2 70841 1 156
2 70842 1 156
2 70843 1 156
2 70844 1 156
2 70845 1 156
2 70846 1 156
2 70847 1 156
2 70848 1 156
2 70849 1 156
2 70850 1 156
2 70851 1 156
2 70852 1 156
2 70853 1 156
2 70854 1 156
2 70855 1 156
2 70856 1 156
2 70857 1 156
2 70858 1 156
2 70859 1 156
2 70860 1 156
2 70861 1 156
2 70862 1 156
2 70863 1 156
2 70864 1 156
2 70865 1 156
2 70866 1 156
2 70867 1 156
2 70868 1 156
2 70869 1 156
2 70870 1 156
2 70871 1 156
2 70872 1 156
2 70873 1 156
2 70874 1 156
2 70875 1 156
2 70876 1 156
2 70877 1 156
2 70878 1 156
2 70879 1 156
2 70880 1 156
2 70881 1 157
2 70882 1 157
2 70883 1 157
2 70884 1 157
2 70885 1 157
2 70886 1 158
2 70887 1 158
2 70888 1 159
2 70889 1 159
2 70890 1 159
2 70891 1 160
2 70892 1 160
2 70893 1 161
2 70894 1 161
2 70895 1 161
2 70896 1 161
2 70897 1 161
2 70898 1 161
2 70899 1 162
2 70900 1 162
2 70901 1 162
2 70902 1 162
2 70903 1 162
2 70904 1 162
2 70905 1 162
2 70906 1 162
2 70907 1 163
2 70908 1 163
2 70909 1 163
2 70910 1 163
2 70911 1 163
2 70912 1 163
2 70913 1 163
2 70914 1 163
2 70915 1 163
2 70916 1 164
2 70917 1 164
2 70918 1 164
2 70919 1 167
2 70920 1 167
2 70921 1 167
2 70922 1 167
2 70923 1 167
2 70924 1 167
2 70925 1 167
2 70926 1 167
2 70927 1 167
2 70928 1 167
2 70929 1 168
2 70930 1 168
2 70931 1 168
2 70932 1 168
2 70933 1 169
2 70934 1 169
2 70935 1 169
2 70936 1 169
2 70937 1 169
2 70938 1 171
2 70939 1 171
2 70940 1 171
2 70941 1 171
2 70942 1 171
2 70943 1 171
2 70944 1 171
2 70945 1 171
2 70946 1 171
2 70947 1 171
2 70948 1 171
2 70949 1 171
2 70950 1 171
2 70951 1 171
2 70952 1 172
2 70953 1 172
2 70954 1 172
2 70955 1 173
2 70956 1 173
2 70957 1 173
2 70958 1 173
2 70959 1 173
2 70960 1 174
2 70961 1 174
2 70962 1 176
2 70963 1 176
2 70964 1 178
2 70965 1 178
2 70966 1 179
2 70967 1 179
2 70968 1 179
2 70969 1 179
2 70970 1 179
2 70971 1 179
2 70972 1 179
2 70973 1 179
2 70974 1 179
2 70975 1 179
2 70976 1 179
2 70977 1 179
2 70978 1 179
2 70979 1 179
2 70980 1 180
2 70981 1 180
2 70982 1 180
2 70983 1 180
2 70984 1 180
2 70985 1 180
2 70986 1 180
2 70987 1 180
2 70988 1 180
2 70989 1 180
2 70990 1 182
2 70991 1 182
2 70992 1 192
2 70993 1 192
2 70994 1 196
2 70995 1 196
2 70996 1 196
2 70997 1 199
2 70998 1 199
2 70999 1 200
2 71000 1 200
2 71001 1 200
2 71002 1 200
2 71003 1 200
2 71004 1 200
2 71005 1 200
2 71006 1 200
2 71007 1 200
2 71008 1 200
2 71009 1 200
2 71010 1 200
2 71011 1 200
2 71012 1 200
2 71013 1 200
2 71014 1 200
2 71015 1 201
2 71016 1 201
2 71017 1 201
2 71018 1 201
2 71019 1 201
2 71020 1 201
2 71021 1 201
2 71022 1 201
2 71023 1 201
2 71024 1 201
2 71025 1 201
2 71026 1 201
2 71027 1 201
2 71028 1 201
2 71029 1 201
2 71030 1 201
2 71031 1 201
2 71032 1 201
2 71033 1 201
2 71034 1 202
2 71035 1 202
2 71036 1 202
2 71037 1 203
2 71038 1 203
2 71039 1 203
2 71040 1 203
2 71041 1 203
2 71042 1 203
2 71043 1 203
2 71044 1 203
2 71045 1 203
2 71046 1 203
2 71047 1 203
2 71048 1 203
2 71049 1 203
2 71050 1 203
2 71051 1 203
2 71052 1 203
2 71053 1 203
2 71054 1 203
2 71055 1 203
2 71056 1 203
2 71057 1 203
2 71058 1 203
2 71059 1 203
2 71060 1 203
2 71061 1 203
2 71062 1 203
2 71063 1 203
2 71064 1 203
2 71065 1 203
2 71066 1 203
2 71067 1 203
2 71068 1 203
2 71069 1 203
2 71070 1 203
2 71071 1 203
2 71072 1 203
2 71073 1 203
2 71074 1 203
2 71075 1 203
2 71076 1 203
2 71077 1 203
2 71078 1 203
2 71079 1 203
2 71080 1 203
2 71081 1 203
2 71082 1 203
2 71083 1 203
2 71084 1 203
2 71085 1 203
2 71086 1 203
2 71087 1 203
2 71088 1 203
2 71089 1 203
2 71090 1 203
2 71091 1 203
2 71092 1 203
2 71093 1 203
2 71094 1 203
2 71095 1 203
2 71096 1 203
2 71097 1 203
2 71098 1 203
2 71099 1 203
2 71100 1 203
2 71101 1 203
2 71102 1 203
2 71103 1 203
2 71104 1 203
2 71105 1 203
2 71106 1 203
2 71107 1 203
2 71108 1 203
2 71109 1 203
2 71110 1 203
2 71111 1 203
2 71112 1 203
2 71113 1 203
2 71114 1 203
2 71115 1 203
2 71116 1 203
2 71117 1 203
2 71118 1 203
2 71119 1 203
2 71120 1 203
2 71121 1 203
2 71122 1 203
2 71123 1 203
2 71124 1 203
2 71125 1 203
2 71126 1 203
2 71127 1 203
2 71128 1 203
2 71129 1 203
2 71130 1 203
2 71131 1 203
2 71132 1 203
2 71133 1 203
2 71134 1 203
2 71135 1 203
2 71136 1 203
2 71137 1 203
2 71138 1 203
2 71139 1 203
2 71140 1 203
2 71141 1 204
2 71142 1 204
2 71143 1 204
2 71144 1 204
2 71145 1 204
2 71146 1 204
2 71147 1 204
2 71148 1 204
2 71149 1 204
2 71150 1 204
2 71151 1 204
2 71152 1 204
2 71153 1 204
2 71154 1 204
2 71155 1 204
2 71156 1 204
2 71157 1 204
2 71158 1 204
2 71159 1 204
2 71160 1 204
2 71161 1 204
2 71162 1 204
2 71163 1 204
2 71164 1 204
2 71165 1 204
2 71166 1 204
2 71167 1 204
2 71168 1 204
2 71169 1 204
2 71170 1 204
2 71171 1 204
2 71172 1 204
2 71173 1 204
2 71174 1 204
2 71175 1 204
2 71176 1 204
2 71177 1 204
2 71178 1 204
2 71179 1 204
2 71180 1 204
2 71181 1 204
2 71182 1 204
2 71183 1 204
2 71184 1 204
2 71185 1 204
2 71186 1 204
2 71187 1 204
2 71188 1 204
2 71189 1 204
2 71190 1 204
2 71191 1 204
2 71192 1 204
2 71193 1 204
2 71194 1 204
2 71195 1 204
2 71196 1 204
2 71197 1 204
2 71198 1 204
2 71199 1 204
2 71200 1 204
2 71201 1 204
2 71202 1 204
2 71203 1 204
2 71204 1 204
2 71205 1 204
2 71206 1 204
2 71207 1 204
2 71208 1 204
2 71209 1 204
2 71210 1 204
2 71211 1 204
2 71212 1 204
2 71213 1 204
2 71214 1 204
2 71215 1 204
2 71216 1 204
2 71217 1 204
2 71218 1 204
2 71219 1 204
2 71220 1 204
2 71221 1 204
2 71222 1 204
2 71223 1 204
2 71224 1 204
2 71225 1 204
2 71226 1 204
2 71227 1 204
2 71228 1 204
2 71229 1 204
2 71230 1 204
2 71231 1 204
2 71232 1 204
2 71233 1 204
2 71234 1 204
2 71235 1 204
2 71236 1 204
2 71237 1 204
2 71238 1 204
2 71239 1 204
2 71240 1 204
2 71241 1 204
2 71242 1 204
2 71243 1 204
2 71244 1 204
2 71245 1 204
2 71246 1 204
2 71247 1 204
2 71248 1 204
2 71249 1 204
2 71250 1 204
2 71251 1 204
2 71252 1 204
2 71253 1 204
2 71254 1 204
2 71255 1 204
2 71256 1 204
2 71257 1 204
2 71258 1 204
2 71259 1 204
2 71260 1 204
2 71261 1 204
2 71262 1 204
2 71263 1 204
2 71264 1 204
2 71265 1 204
2 71266 1 204
2 71267 1 204
2 71268 1 204
2 71269 1 204
2 71270 1 205
2 71271 1 205
2 71272 1 205
2 71273 1 205
2 71274 1 205
2 71275 1 205
2 71276 1 206
2 71277 1 206
2 71278 1 206
2 71279 1 206
2 71280 1 206
2 71281 1 214
2 71282 1 214
2 71283 1 214
2 71284 1 214
2 71285 1 214
2 71286 1 214
2 71287 1 214
2 71288 1 214
2 71289 1 214
2 71290 1 214
2 71291 1 214
2 71292 1 214
2 71293 1 214
2 71294 1 214
2 71295 1 214
2 71296 1 214
2 71297 1 214
2 71298 1 215
2 71299 1 215
2 71300 1 215
2 71301 1 215
2 71302 1 215
2 71303 1 215
2 71304 1 215
2 71305 1 215
2 71306 1 215
2 71307 1 215
2 71308 1 215
2 71309 1 215
2 71310 1 215
2 71311 1 215
2 71312 1 215
2 71313 1 215
2 71314 1 215
2 71315 1 215
2 71316 1 215
2 71317 1 216
2 71318 1 216
2 71319 1 216
2 71320 1 216
2 71321 1 216
2 71322 1 216
2 71323 1 216
2 71324 1 216
2 71325 1 216
2 71326 1 216
2 71327 1 216
2 71328 1 216
2 71329 1 217
2 71330 1 217
2 71331 1 217
2 71332 1 217
2 71333 1 217
2 71334 1 217
2 71335 1 217
2 71336 1 217
2 71337 1 217
2 71338 1 217
2 71339 1 218
2 71340 1 218
2 71341 1 218
2 71342 1 219
2 71343 1 219
2 71344 1 219
2 71345 1 219
2 71346 1 219
2 71347 1 219
2 71348 1 219
2 71349 1 219
2 71350 1 219
2 71351 1 219
2 71352 1 219
2 71353 1 219
2 71354 1 219
2 71355 1 219
2 71356 1 219
2 71357 1 219
2 71358 1 219
2 71359 1 219
2 71360 1 219
2 71361 1 219
2 71362 1 219
2 71363 1 220
2 71364 1 220
2 71365 1 220
2 71366 1 220
2 71367 1 220
2 71368 1 220
2 71369 1 220
2 71370 1 220
2 71371 1 220
2 71372 1 220
2 71373 1 220
2 71374 1 220
2 71375 1 220
2 71376 1 220
2 71377 1 220
2 71378 1 221
2 71379 1 221
2 71380 1 221
2 71381 1 221
2 71382 1 222
2 71383 1 222
2 71384 1 223
2 71385 1 223
2 71386 1 223
2 71387 1 223
2 71388 1 223
2 71389 1 223
2 71390 1 223
2 71391 1 223
2 71392 1 223
2 71393 1 223
2 71394 1 223
2 71395 1 223
2 71396 1 223
2 71397 1 223
2 71398 1 223
2 71399 1 223
2 71400 1 224
2 71401 1 224
2 71402 1 225
2 71403 1 225
2 71404 1 225
2 71405 1 225
2 71406 1 225
2 71407 1 225
2 71408 1 226
2 71409 1 226
2 71410 1 226
2 71411 1 226
2 71412 1 226
2 71413 1 226
2 71414 1 226
2 71415 1 226
2 71416 1 226
2 71417 1 226
2 71418 1 226
2 71419 1 226
2 71420 1 226
2 71421 1 226
2 71422 1 226
2 71423 1 226
2 71424 1 226
2 71425 1 226
2 71426 1 226
2 71427 1 226
2 71428 1 226
2 71429 1 227
2 71430 1 227
2 71431 1 227
2 71432 1 227
2 71433 1 227
2 71434 1 227
2 71435 1 227
2 71436 1 227
2 71437 1 228
2 71438 1 228
2 71439 1 228
2 71440 1 228
2 71441 1 228
2 71442 1 228
2 71443 1 228
2 71444 1 230
2 71445 1 230
2 71446 1 230
2 71447 1 230
2 71448 1 233
2 71449 1 233
2 71450 1 233
2 71451 1 233
2 71452 1 233
2 71453 1 233
2 71454 1 233
2 71455 1 233
2 71456 1 233
2 71457 1 233
2 71458 1 233
2 71459 1 233
2 71460 1 233
2 71461 1 233
2 71462 1 233
2 71463 1 233
2 71464 1 234
2 71465 1 234
2 71466 1 234
2 71467 1 234
2 71468 1 234
2 71469 1 234
2 71470 1 234
2 71471 1 234
2 71472 1 234
2 71473 1 235
2 71474 1 235
2 71475 1 235
2 71476 1 235
2 71477 1 235
2 71478 1 235
2 71479 1 235
2 71480 1 235
2 71481 1 235
2 71482 1 235
2 71483 1 235
2 71484 1 235
2 71485 1 235
2 71486 1 235
2 71487 1 235
2 71488 1 235
2 71489 1 235
2 71490 1 235
2 71491 1 235
2 71492 1 235
2 71493 1 235
2 71494 1 235
2 71495 1 235
2 71496 1 235
2 71497 1 235
2 71498 1 235
2 71499 1 235
2 71500 1 235
2 71501 1 235
2 71502 1 235
2 71503 1 235
2 71504 1 235
2 71505 1 235
2 71506 1 235
2 71507 1 235
2 71508 1 235
2 71509 1 235
2 71510 1 235
2 71511 1 235
2 71512 1 236
2 71513 1 236
2 71514 1 236
2 71515 1 236
2 71516 1 236
2 71517 1 236
2 71518 1 236
2 71519 1 236
2 71520 1 236
2 71521 1 236
2 71522 1 236
2 71523 1 236
2 71524 1 236
2 71525 1 236
2 71526 1 236
2 71527 1 237
2 71528 1 237
2 71529 1 237
2 71530 1 237
2 71531 1 237
2 71532 1 237
2 71533 1 237
2 71534 1 237
2 71535 1 237
2 71536 1 237
2 71537 1 237
2 71538 1 237
2 71539 1 237
2 71540 1 237
2 71541 1 237
2 71542 1 237
2 71543 1 237
2 71544 1 237
2 71545 1 237
2 71546 1 237
2 71547 1 237
2 71548 1 237
2 71549 1 237
2 71550 1 237
2 71551 1 237
2 71552 1 237
2 71553 1 237
2 71554 1 237
2 71555 1 237
2 71556 1 237
2 71557 1 237
2 71558 1 237
2 71559 1 237
2 71560 1 237
2 71561 1 237
2 71562 1 237
2 71563 1 237
2 71564 1 237
2 71565 1 237
2 71566 1 237
2 71567 1 237
2 71568 1 237
2 71569 1 237
2 71570 1 237
2 71571 1 237
2 71572 1 237
2 71573 1 237
2 71574 1 237
2 71575 1 237
2 71576 1 237
2 71577 1 237
2 71578 1 237
2 71579 1 237
2 71580 1 237
2 71581 1 237
2 71582 1 237
2 71583 1 237
2 71584 1 237
2 71585 1 237
2 71586 1 237
2 71587 1 237
2 71588 1 238
2 71589 1 238
2 71590 1 239
2 71591 1 239
2 71592 1 239
2 71593 1 239
2 71594 1 239
2 71595 1 239
2 71596 1 239
2 71597 1 239
2 71598 1 239
2 71599 1 239
2 71600 1 239
2 71601 1 239
2 71602 1 239
2 71603 1 239
2 71604 1 239
2 71605 1 239
2 71606 1 239
2 71607 1 242
2 71608 1 242
2 71609 1 242
2 71610 1 242
2 71611 1 242
2 71612 1 242
2 71613 1 242
2 71614 1 242
2 71615 1 242
2 71616 1 242
2 71617 1 242
2 71618 1 242
2 71619 1 242
2 71620 1 242
2 71621 1 242
2 71622 1 242
2 71623 1 243
2 71624 1 243
2 71625 1 243
2 71626 1 243
2 71627 1 243
2 71628 1 243
2 71629 1 243
2 71630 1 243
2 71631 1 243
2 71632 1 245
2 71633 1 245
2 71634 1 245
2 71635 1 245
2 71636 1 245
2 71637 1 245
2 71638 1 245
2 71639 1 246
2 71640 1 246
2 71641 1 252
2 71642 1 252
2 71643 1 252
2 71644 1 252
2 71645 1 252
2 71646 1 252
2 71647 1 252
2 71648 1 252
2 71649 1 252
2 71650 1 252
2 71651 1 252
2 71652 1 252
2 71653 1 254
2 71654 1 254
2 71655 1 254
2 71656 1 266
2 71657 1 266
2 71658 1 266
2 71659 1 267
2 71660 1 267
2 71661 1 274
2 71662 1 274
2 71663 1 274
2 71664 1 274
2 71665 1 274
2 71666 1 274
2 71667 1 274
2 71668 1 274
2 71669 1 274
2 71670 1 274
2 71671 1 275
2 71672 1 275
2 71673 1 275
2 71674 1 275
2 71675 1 275
2 71676 1 275
2 71677 1 275
2 71678 1 275
2 71679 1 275
2 71680 1 275
2 71681 1 275
2 71682 1 275
2 71683 1 275
2 71684 1 275
2 71685 1 275
2 71686 1 275
2 71687 1 275
2 71688 1 275
2 71689 1 275
2 71690 1 275
2 71691 1 275
2 71692 1 275
2 71693 1 275
2 71694 1 275
2 71695 1 275
2 71696 1 275
2 71697 1 275
2 71698 1 275
2 71699 1 275
2 71700 1 275
2 71701 1 275
2 71702 1 275
2 71703 1 275
2 71704 1 275
2 71705 1 275
2 71706 1 275
2 71707 1 275
2 71708 1 275
2 71709 1 275
2 71710 1 275
2 71711 1 275
2 71712 1 275
2 71713 1 275
2 71714 1 275
2 71715 1 275
2 71716 1 275
2 71717 1 275
2 71718 1 275
2 71719 1 275
2 71720 1 275
2 71721 1 275
2 71722 1 275
2 71723 1 275
2 71724 1 275
2 71725 1 275
2 71726 1 275
2 71727 1 275
2 71728 1 275
2 71729 1 275
2 71730 1 275
2 71731 1 276
2 71732 1 276
2 71733 1 276
2 71734 1 276
2 71735 1 276
2 71736 1 276
2 71737 1 276
2 71738 1 276
2 71739 1 276
2 71740 1 276
2 71741 1 276
2 71742 1 276
2 71743 1 276
2 71744 1 276
2 71745 1 276
2 71746 1 276
2 71747 1 276
2 71748 1 276
2 71749 1 276
2 71750 1 276
2 71751 1 276
2 71752 1 276
2 71753 1 276
2 71754 1 276
2 71755 1 276
2 71756 1 276
2 71757 1 276
2 71758 1 276
2 71759 1 276
2 71760 1 276
2 71761 1 276
2 71762 1 276
2 71763 1 276
2 71764 1 276
2 71765 1 276
2 71766 1 276
2 71767 1 276
2 71768 1 276
2 71769 1 276
2 71770 1 276
2 71771 1 276
2 71772 1 276
2 71773 1 276
2 71774 1 276
2 71775 1 276
2 71776 1 276
2 71777 1 276
2 71778 1 276
2 71779 1 276
2 71780 1 276
2 71781 1 276
2 71782 1 276
2 71783 1 276
2 71784 1 276
2 71785 1 276
2 71786 1 276
2 71787 1 276
2 71788 1 276
2 71789 1 276
2 71790 1 276
2 71791 1 276
2 71792 1 276
2 71793 1 276
2 71794 1 276
2 71795 1 276
2 71796 1 276
2 71797 1 276
2 71798 1 276
2 71799 1 276
2 71800 1 276
2 71801 1 276
2 71802 1 276
2 71803 1 276
2 71804 1 276
2 71805 1 276
2 71806 1 276
2 71807 1 276
2 71808 1 276
2 71809 1 276
2 71810 1 276
2 71811 1 276
2 71812 1 276
2 71813 1 276
2 71814 1 276
2 71815 1 276
2 71816 1 276
2 71817 1 276
2 71818 1 276
2 71819 1 276
2 71820 1 276
2 71821 1 276
2 71822 1 276
2 71823 1 276
2 71824 1 276
2 71825 1 276
2 71826 1 276
2 71827 1 276
2 71828 1 276
2 71829 1 276
2 71830 1 276
2 71831 1 276
2 71832 1 276
2 71833 1 276
2 71834 1 276
2 71835 1 276
2 71836 1 276
2 71837 1 276
2 71838 1 276
2 71839 1 276
2 71840 1 276
2 71841 1 276
2 71842 1 276
2 71843 1 276
2 71844 1 277
2 71845 1 277
2 71846 1 277
2 71847 1 278
2 71848 1 278
2 71849 1 279
2 71850 1 279
2 71851 1 281
2 71852 1 281
2 71853 1 282
2 71854 1 282
2 71855 1 284
2 71856 1 284
2 71857 1 289
2 71858 1 289
2 71859 1 289
2 71860 1 289
2 71861 1 289
2 71862 1 289
2 71863 1 289
2 71864 1 289
2 71865 1 289
2 71866 1 289
2 71867 1 289
2 71868 1 289
2 71869 1 289
2 71870 1 289
2 71871 1 289
2 71872 1 289
2 71873 1 289
2 71874 1 289
2 71875 1 289
2 71876 1 289
2 71877 1 289
2 71878 1 289
2 71879 1 289
2 71880 1 289
2 71881 1 289
2 71882 1 289
2 71883 1 289
2 71884 1 289
2 71885 1 289
2 71886 1 289
2 71887 1 289
2 71888 1 289
2 71889 1 289
2 71890 1 289
2 71891 1 289
2 71892 1 289
2 71893 1 289
2 71894 1 289
2 71895 1 289
2 71896 1 289
2 71897 1 289
2 71898 1 289
2 71899 1 289
2 71900 1 289
2 71901 1 289
2 71902 1 289
2 71903 1 290
2 71904 1 290
2 71905 1 290
2 71906 1 290
2 71907 1 290
2 71908 1 290
2 71909 1 290
2 71910 1 290
2 71911 1 290
2 71912 1 290
2 71913 1 290
2 71914 1 290
2 71915 1 290
2 71916 1 290
2 71917 1 290
2 71918 1 290
2 71919 1 290
2 71920 1 290
2 71921 1 290
2 71922 1 290
2 71923 1 290
2 71924 1 290
2 71925 1 290
2 71926 1 290
2 71927 1 290
2 71928 1 290
2 71929 1 290
2 71930 1 290
2 71931 1 290
2 71932 1 290
2 71933 1 290
2 71934 1 290
2 71935 1 290
2 71936 1 290
2 71937 1 290
2 71938 1 290
2 71939 1 290
2 71940 1 290
2 71941 1 290
2 71942 1 291
2 71943 1 291
2 71944 1 291
2 71945 1 291
2 71946 1 291
2 71947 1 291
2 71948 1 291
2 71949 1 291
2 71950 1 291
2 71951 1 291
2 71952 1 291
2 71953 1 291
2 71954 1 291
2 71955 1 291
2 71956 1 291
2 71957 1 291
2 71958 1 291
2 71959 1 291
2 71960 1 291
2 71961 1 291
2 71962 1 291
2 71963 1 291
2 71964 1 291
2 71965 1 291
2 71966 1 291
2 71967 1 291
2 71968 1 291
2 71969 1 291
2 71970 1 291
2 71971 1 291
2 71972 1 291
2 71973 1 291
2 71974 1 291
2 71975 1 291
2 71976 1 291
2 71977 1 291
2 71978 1 291
2 71979 1 291
2 71980 1 291
2 71981 1 291
2 71982 1 291
2 71983 1 291
2 71984 1 291
2 71985 1 291
2 71986 1 291
2 71987 1 291
2 71988 1 291
2 71989 1 291
2 71990 1 291
2 71991 1 291
2 71992 1 291
2 71993 1 291
2 71994 1 291
2 71995 1 291
2 71996 1 291
2 71997 1 291
2 71998 1 291
2 71999 1 291
2 72000 1 291
2 72001 1 291
2 72002 1 291
2 72003 1 291
2 72004 1 291
2 72005 1 291
2 72006 1 291
2 72007 1 291
2 72008 1 291
2 72009 1 291
2 72010 1 291
2 72011 1 291
2 72012 1 291
2 72013 1 291
2 72014 1 291
2 72015 1 291
2 72016 1 291
2 72017 1 291
2 72018 1 291
2 72019 1 291
2 72020 1 291
2 72021 1 291
2 72022 1 291
2 72023 1 291
2 72024 1 291
2 72025 1 291
2 72026 1 291
2 72027 1 291
2 72028 1 291
2 72029 1 291
2 72030 1 291
2 72031 1 291
2 72032 1 291
2 72033 1 292
2 72034 1 292
2 72035 1 292
2 72036 1 292
2 72037 1 292
2 72038 1 292
2 72039 1 292
2 72040 1 292
2 72041 1 292
2 72042 1 292
2 72043 1 292
2 72044 1 292
2 72045 1 292
2 72046 1 292
2 72047 1 292
2 72048 1 292
2 72049 1 292
2 72050 1 292
2 72051 1 292
2 72052 1 292
2 72053 1 292
2 72054 1 292
2 72055 1 292
2 72056 1 292
2 72057 1 292
2 72058 1 292
2 72059 1 292
2 72060 1 292
2 72061 1 292
2 72062 1 292
2 72063 1 292
2 72064 1 292
2 72065 1 292
2 72066 1 292
2 72067 1 292
2 72068 1 292
2 72069 1 292
2 72070 1 292
2 72071 1 292
2 72072 1 292
2 72073 1 292
2 72074 1 292
2 72075 1 292
2 72076 1 292
2 72077 1 292
2 72078 1 292
2 72079 1 292
2 72080 1 292
2 72081 1 292
2 72082 1 292
2 72083 1 292
2 72084 1 292
2 72085 1 292
2 72086 1 292
2 72087 1 292
2 72088 1 292
2 72089 1 292
2 72090 1 292
2 72091 1 292
2 72092 1 292
2 72093 1 292
2 72094 1 292
2 72095 1 292
2 72096 1 292
2 72097 1 292
2 72098 1 292
2 72099 1 292
2 72100 1 292
2 72101 1 292
2 72102 1 292
2 72103 1 292
2 72104 1 292
2 72105 1 292
2 72106 1 292
2 72107 1 292
2 72108 1 292
2 72109 1 292
2 72110 1 292
2 72111 1 292
2 72112 1 292
2 72113 1 292
2 72114 1 292
2 72115 1 292
2 72116 1 292
2 72117 1 292
2 72118 1 292
2 72119 1 292
2 72120 1 292
2 72121 1 292
2 72122 1 292
2 72123 1 292
2 72124 1 292
2 72125 1 292
2 72126 1 292
2 72127 1 292
2 72128 1 292
2 72129 1 292
2 72130 1 292
2 72131 1 292
2 72132 1 292
2 72133 1 292
2 72134 1 292
2 72135 1 292
2 72136 1 292
2 72137 1 292
2 72138 1 292
2 72139 1 292
2 72140 1 292
2 72141 1 293
2 72142 1 293
2 72143 1 293
2 72144 1 294
2 72145 1 294
2 72146 1 294
2 72147 1 294
2 72148 1 294
2 72149 1 294
2 72150 1 301
2 72151 1 301
2 72152 1 301
2 72153 1 301
2 72154 1 301
2 72155 1 301
2 72156 1 302
2 72157 1 302
2 72158 1 302
2 72159 1 302
2 72160 1 302
2 72161 1 302
2 72162 1 302
2 72163 1 302
2 72164 1 303
2 72165 1 303
2 72166 1 303
2 72167 1 303
2 72168 1 303
2 72169 1 303
2 72170 1 303
2 72171 1 303
2 72172 1 303
2 72173 1 304
2 72174 1 304
2 72175 1 304
2 72176 1 304
2 72177 1 304
2 72178 1 304
2 72179 1 304
2 72180 1 304
2 72181 1 304
2 72182 1 304
2 72183 1 304
2 72184 1 304
2 72185 1 304
2 72186 1 304
2 72187 1 304
2 72188 1 304
2 72189 1 304
2 72190 1 304
2 72191 1 304
2 72192 1 304
2 72193 1 304
2 72194 1 304
2 72195 1 305
2 72196 1 305
2 72197 1 305
2 72198 1 305
2 72199 1 305
2 72200 1 305
2 72201 1 305
2 72202 1 305
2 72203 1 305
2 72204 1 305
2 72205 1 305
2 72206 1 305
2 72207 1 305
2 72208 1 305
2 72209 1 305
2 72210 1 305
2 72211 1 305
2 72212 1 305
2 72213 1 305
2 72214 1 305
2 72215 1 305
2 72216 1 305
2 72217 1 305
2 72218 1 305
2 72219 1 305
2 72220 1 305
2 72221 1 305
2 72222 1 305
2 72223 1 305
2 72224 1 305
2 72225 1 305
2 72226 1 305
2 72227 1 305
2 72228 1 305
2 72229 1 305
2 72230 1 305
2 72231 1 305
2 72232 1 305
2 72233 1 305
2 72234 1 305
2 72235 1 305
2 72236 1 305
2 72237 1 305
2 72238 1 305
2 72239 1 305
2 72240 1 305
2 72241 1 305
2 72242 1 305
2 72243 1 305
2 72244 1 305
2 72245 1 305
2 72246 1 305
2 72247 1 305
2 72248 1 305
2 72249 1 305
2 72250 1 305
2 72251 1 305
2 72252 1 305
2 72253 1 305
2 72254 1 305
2 72255 1 305
2 72256 1 305
2 72257 1 305
2 72258 1 305
2 72259 1 305
2 72260 1 305
2 72261 1 305
2 72262 1 305
2 72263 1 305
2 72264 1 305
2 72265 1 305
2 72266 1 305
2 72267 1 305
2 72268 1 305
2 72269 1 305
2 72270 1 305
2 72271 1 305
2 72272 1 305
2 72273 1 305
2 72274 1 305
2 72275 1 305
2 72276 1 305
2 72277 1 305
2 72278 1 305
2 72279 1 306
2 72280 1 306
2 72281 1 306
2 72282 1 306
2 72283 1 306
2 72284 1 306
2 72285 1 306
2 72286 1 306
2 72287 1 306
2 72288 1 306
2 72289 1 306
2 72290 1 306
2 72291 1 306
2 72292 1 306
2 72293 1 306
2 72294 1 306
2 72295 1 306
2 72296 1 306
2 72297 1 306
2 72298 1 306
2 72299 1 306
2 72300 1 306
2 72301 1 306
2 72302 1 306
2 72303 1 306
2 72304 1 306
2 72305 1 306
2 72306 1 306
2 72307 1 306
2 72308 1 306
2 72309 1 306
2 72310 1 306
2 72311 1 306
2 72312 1 306
2 72313 1 306
2 72314 1 306
2 72315 1 306
2 72316 1 306
2 72317 1 306
2 72318 1 306
2 72319 1 306
2 72320 1 306
2 72321 1 306
2 72322 1 306
2 72323 1 306
2 72324 1 306
2 72325 1 306
2 72326 1 306
2 72327 1 306
2 72328 1 306
2 72329 1 306
2 72330 1 306
2 72331 1 306
2 72332 1 306
2 72333 1 306
2 72334 1 306
2 72335 1 306
2 72336 1 306
2 72337 1 306
2 72338 1 306
2 72339 1 306
2 72340 1 306
2 72341 1 306
2 72342 1 306
2 72343 1 306
2 72344 1 306
2 72345 1 306
2 72346 1 306
2 72347 1 306
2 72348 1 306
2 72349 1 306
2 72350 1 306
2 72351 1 306
2 72352 1 306
2 72353 1 306
2 72354 1 306
2 72355 1 306
2 72356 1 306
2 72357 1 306
2 72358 1 306
2 72359 1 306
2 72360 1 306
2 72361 1 306
2 72362 1 306
2 72363 1 306
2 72364 1 306
2 72365 1 306
2 72366 1 306
2 72367 1 306
2 72368 1 306
2 72369 1 306
2 72370 1 306
2 72371 1 306
2 72372 1 306
2 72373 1 306
2 72374 1 306
2 72375 1 306
2 72376 1 306
2 72377 1 306
2 72378 1 306
2 72379 1 306
2 72380 1 306
2 72381 1 306
2 72382 1 306
2 72383 1 306
2 72384 1 306
2 72385 1 306
2 72386 1 306
2 72387 1 306
2 72388 1 306
2 72389 1 306
2 72390 1 306
2 72391 1 306
2 72392 1 306
2 72393 1 306
2 72394 1 306
2 72395 1 306
2 72396 1 306
2 72397 1 306
2 72398 1 306
2 72399 1 306
2 72400 1 306
2 72401 1 306
2 72402 1 306
2 72403 1 306
2 72404 1 306
2 72405 1 306
2 72406 1 307
2 72407 1 307
2 72408 1 307
2 72409 1 307
2 72410 1 307
2 72411 1 307
2 72412 1 307
2 72413 1 307
2 72414 1 307
2 72415 1 307
2 72416 1 307
2 72417 1 308
2 72418 1 308
2 72419 1 308
2 72420 1 308
2 72421 1 308
2 72422 1 308
2 72423 1 308
2 72424 1 309
2 72425 1 309
2 72426 1 310
2 72427 1 310
2 72428 1 310
2 72429 1 314
2 72430 1 314
2 72431 1 317
2 72432 1 317
2 72433 1 317
2 72434 1 317
2 72435 1 317
2 72436 1 317
2 72437 1 317
2 72438 1 317
2 72439 1 317
2 72440 1 318
2 72441 1 318
2 72442 1 318
2 72443 1 319
2 72444 1 319
2 72445 1 319
2 72446 1 319
2 72447 1 319
2 72448 1 319
2 72449 1 319
2 72450 1 320
2 72451 1 320
2 72452 1 320
2 72453 1 320
2 72454 1 320
2 72455 1 320
2 72456 1 320
2 72457 1 320
2 72458 1 321
2 72459 1 321
2 72460 1 322
2 72461 1 322
2 72462 1 322
2 72463 1 322
2 72464 1 323
2 72465 1 323
2 72466 1 323
2 72467 1 323
2 72468 1 323
2 72469 1 323
2 72470 1 324
2 72471 1 324
2 72472 1 324
2 72473 1 324
2 72474 1 324
2 72475 1 324
2 72476 1 324
2 72477 1 324
2 72478 1 325
2 72479 1 325
2 72480 1 338
2 72481 1 338
2 72482 1 338
2 72483 1 339
2 72484 1 339
2 72485 1 339
2 72486 1 339
2 72487 1 339
2 72488 1 339
2 72489 1 339
2 72490 1 339
2 72491 1 339
2 72492 1 339
2 72493 1 339
2 72494 1 339
2 72495 1 339
2 72496 1 339
2 72497 1 339
2 72498 1 339
2 72499 1 339
2 72500 1 339
2 72501 1 339
2 72502 1 339
2 72503 1 339
2 72504 1 339
2 72505 1 339
2 72506 1 339
2 72507 1 339
2 72508 1 339
2 72509 1 339
2 72510 1 339
2 72511 1 339
2 72512 1 339
2 72513 1 340
2 72514 1 340
2 72515 1 340
2 72516 1 340
2 72517 1 340
2 72518 1 340
2 72519 1 340
2 72520 1 340
2 72521 1 340
2 72522 1 340
2 72523 1 340
2 72524 1 340
2 72525 1 341
2 72526 1 341
2 72527 1 341
2 72528 1 341
2 72529 1 341
2 72530 1 341
2 72531 1 341
2 72532 1 341
2 72533 1 341
2 72534 1 341
2 72535 1 341
2 72536 1 341
2 72537 1 341
2 72538 1 341
2 72539 1 341
2 72540 1 341
2 72541 1 341
2 72542 1 341
2 72543 1 341
2 72544 1 341
2 72545 1 341
2 72546 1 341
2 72547 1 341
2 72548 1 341
2 72549 1 341
2 72550 1 341
2 72551 1 341
2 72552 1 341
2 72553 1 341
2 72554 1 341
2 72555 1 341
2 72556 1 341
2 72557 1 341
2 72558 1 341
2 72559 1 341
2 72560 1 341
2 72561 1 341
2 72562 1 341
2 72563 1 341
2 72564 1 342
2 72565 1 342
2 72566 1 342
2 72567 1 342
2 72568 1 342
2 72569 1 342
2 72570 1 342
2 72571 1 342
2 72572 1 342
2 72573 1 342
2 72574 1 342
2 72575 1 342
2 72576 1 343
2 72577 1 343
2 72578 1 343
2 72579 1 343
2 72580 1 343
2 72581 1 343
2 72582 1 343
2 72583 1 343
2 72584 1 343
2 72585 1 343
2 72586 1 343
2 72587 1 343
2 72588 1 343
2 72589 1 343
2 72590 1 343
2 72591 1 343
2 72592 1 343
2 72593 1 343
2 72594 1 343
2 72595 1 343
2 72596 1 343
2 72597 1 343
2 72598 1 343
2 72599 1 343
2 72600 1 343
2 72601 1 343
2 72602 1 343
2 72603 1 343
2 72604 1 343
2 72605 1 343
2 72606 1 343
2 72607 1 343
2 72608 1 343
2 72609 1 343
2 72610 1 344
2 72611 1 344
2 72612 1 344
2 72613 1 346
2 72614 1 346
2 72615 1 346
2 72616 1 346
2 72617 1 346
2 72618 1 346
2 72619 1 347
2 72620 1 347
2 72621 1 347
2 72622 1 348
2 72623 1 348
2 72624 1 349
2 72625 1 349
2 72626 1 350
2 72627 1 350
2 72628 1 350
2 72629 1 350
2 72630 1 351
2 72631 1 351
2 72632 1 351
2 72633 1 351
2 72634 1 351
2 72635 1 351
2 72636 1 352
2 72637 1 352
2 72638 1 352
2 72639 1 355
2 72640 1 355
2 72641 1 358
2 72642 1 358
2 72643 1 366
2 72644 1 366
2 72645 1 367
2 72646 1 367
2 72647 1 368
2 72648 1 368
2 72649 1 368
2 72650 1 370
2 72651 1 370
2 72652 1 370
2 72653 1 370
2 72654 1 370
2 72655 1 371
2 72656 1 371
2 72657 1 371
2 72658 1 371
2 72659 1 373
2 72660 1 373
2 72661 1 373
2 72662 1 373
2 72663 1 373
2 72664 1 374
2 72665 1 374
2 72666 1 374
2 72667 1 374
2 72668 1 374
2 72669 1 374
2 72670 1 374
2 72671 1 374
2 72672 1 374
2 72673 1 374
2 72674 1 374
2 72675 1 374
2 72676 1 374
2 72677 1 374
2 72678 1 375
2 72679 1 375
2 72680 1 375
2 72681 1 375
2 72682 1 375
2 72683 1 375
2 72684 1 375
2 72685 1 375
2 72686 1 375
2 72687 1 375
2 72688 1 375
2 72689 1 375
2 72690 1 375
2 72691 1 375
2 72692 1 375
2 72693 1 375
2 72694 1 375
2 72695 1 375
2 72696 1 375
2 72697 1 375
2 72698 1 375
2 72699 1 375
2 72700 1 375
2 72701 1 375
2 72702 1 375
2 72703 1 375
2 72704 1 375
2 72705 1 375
2 72706 1 375
2 72707 1 375
2 72708 1 375
2 72709 1 375
2 72710 1 375
2 72711 1 375
2 72712 1 375
2 72713 1 375
2 72714 1 375
2 72715 1 375
2 72716 1 375
2 72717 1 375
2 72718 1 375
2 72719 1 375
2 72720 1 375
2 72721 1 375
2 72722 1 375
2 72723 1 375
2 72724 1 375
2 72725 1 375
2 72726 1 375
2 72727 1 375
2 72728 1 377
2 72729 1 377
2 72730 1 379
2 72731 1 379
2 72732 1 379
2 72733 1 380
2 72734 1 380
2 72735 1 382
2 72736 1 382
2 72737 1 382
2 72738 1 382
2 72739 1 382
2 72740 1 382
2 72741 1 382
2 72742 1 382
2 72743 1 382
2 72744 1 385
2 72745 1 385
2 72746 1 395
2 72747 1 395
2 72748 1 395
2 72749 1 395
2 72750 1 395
2 72751 1 396
2 72752 1 396
2 72753 1 396
2 72754 1 396
2 72755 1 396
2 72756 1 397
2 72757 1 397
2 72758 1 398
2 72759 1 398
2 72760 1 398
2 72761 1 398
2 72762 1 398
2 72763 1 398
2 72764 1 398
2 72765 1 398
2 72766 1 398
2 72767 1 398
2 72768 1 398
2 72769 1 398
2 72770 1 398
2 72771 1 398
2 72772 1 398
2 72773 1 398
2 72774 1 399
2 72775 1 399
2 72776 1 399
2 72777 1 399
2 72778 1 399
2 72779 1 399
2 72780 1 399
2 72781 1 399
2 72782 1 399
2 72783 1 400
2 72784 1 400
2 72785 1 400
2 72786 1 400
2 72787 1 400
2 72788 1 400
2 72789 1 401
2 72790 1 401
2 72791 1 401
2 72792 1 401
2 72793 1 401
2 72794 1 402
2 72795 1 402
2 72796 1 402
2 72797 1 403
2 72798 1 403
2 72799 1 403
2 72800 1 403
2 72801 1 406
2 72802 1 406
2 72803 1 406
2 72804 1 406
2 72805 1 406
2 72806 1 406
2 72807 1 408
2 72808 1 408
2 72809 1 410
2 72810 1 410
2 72811 1 410
2 72812 1 410
2 72813 1 410
2 72814 1 410
2 72815 1 410
2 72816 1 410
2 72817 1 410
2 72818 1 410
2 72819 1 410
2 72820 1 410
2 72821 1 411
2 72822 1 411
2 72823 1 411
2 72824 1 414
2 72825 1 414
2 72826 1 414
2 72827 1 415
2 72828 1 415
2 72829 1 415
2 72830 1 415
2 72831 1 415
2 72832 1 415
2 72833 1 415
2 72834 1 415
2 72835 1 415
2 72836 1 415
2 72837 1 415
2 72838 1 415
2 72839 1 416
2 72840 1 416
2 72841 1 417
2 72842 1 417
2 72843 1 418
2 72844 1 418
2 72845 1 418
2 72846 1 418
2 72847 1 418
2 72848 1 418
2 72849 1 418
2 72850 1 418
2 72851 1 419
2 72852 1 419
2 72853 1 419
2 72854 1 419
2 72855 1 419
2 72856 1 419
2 72857 1 419
2 72858 1 420
2 72859 1 420
2 72860 1 420
2 72861 1 420
2 72862 1 420
2 72863 1 420
2 72864 1 420
2 72865 1 420
2 72866 1 420
2 72867 1 421
2 72868 1 421
2 72869 1 421
2 72870 1 422
2 72871 1 422
2 72872 1 422
2 72873 1 423
2 72874 1 423
2 72875 1 423
2 72876 1 423
2 72877 1 423
2 72878 1 423
2 72879 1 423
2 72880 1 423
2 72881 1 425
2 72882 1 425
2 72883 1 426
2 72884 1 426
2 72885 1 426
2 72886 1 442
2 72887 1 442
2 72888 1 442
2 72889 1 442
2 72890 1 442
2 72891 1 442
2 72892 1 443
2 72893 1 443
2 72894 1 443
2 72895 1 443
2 72896 1 443
2 72897 1 443
2 72898 1 443
2 72899 1 443
2 72900 1 443
2 72901 1 443
2 72902 1 443
2 72903 1 443
2 72904 1 443
2 72905 1 443
2 72906 1 443
2 72907 1 443
2 72908 1 443
2 72909 1 443
2 72910 1 443
2 72911 1 443
2 72912 1 443
2 72913 1 443
2 72914 1 443
2 72915 1 443
2 72916 1 443
2 72917 1 443
2 72918 1 443
2 72919 1 443
2 72920 1 443
2 72921 1 443
2 72922 1 443
2 72923 1 443
2 72924 1 443
2 72925 1 443
2 72926 1 443
2 72927 1 443
2 72928 1 443
2 72929 1 443
2 72930 1 443
2 72931 1 443
2 72932 1 443
2 72933 1 443
2 72934 1 443
2 72935 1 443
2 72936 1 443
2 72937 1 446
2 72938 1 446
2 72939 1 446
2 72940 1 446
2 72941 1 446
2 72942 1 446
2 72943 1 446
2 72944 1 446
2 72945 1 446
2 72946 1 446
2 72947 1 446
2 72948 1 446
2 72949 1 446
2 72950 1 446
2 72951 1 446
2 72952 1 446
2 72953 1 446
2 72954 1 446
2 72955 1 446
2 72956 1 446
2 72957 1 447
2 72958 1 447
2 72959 1 447
2 72960 1 447
2 72961 1 447
2 72962 1 448
2 72963 1 448
2 72964 1 448
2 72965 1 448
2 72966 1 448
2 72967 1 448
2 72968 1 448
2 72969 1 448
2 72970 1 449
2 72971 1 449
2 72972 1 449
2 72973 1 450
2 72974 1 450
2 72975 1 450
2 72976 1 450
2 72977 1 450
2 72978 1 450
2 72979 1 450
2 72980 1 450
2 72981 1 450
2 72982 1 450
2 72983 1 450
2 72984 1 450
2 72985 1 450
2 72986 1 450
2 72987 1 450
2 72988 1 450
2 72989 1 450
2 72990 1 453
2 72991 1 453
2 72992 1 453
2 72993 1 453
2 72994 1 453
2 72995 1 453
2 72996 1 453
2 72997 1 453
2 72998 1 453
2 72999 1 453
2 73000 1 453
2 73001 1 453
2 73002 1 453
2 73003 1 453
2 73004 1 453
2 73005 1 453
2 73006 1 453
2 73007 1 453
2 73008 1 453
2 73009 1 453
2 73010 1 453
2 73011 1 453
2 73012 1 453
2 73013 1 453
2 73014 1 453
2 73015 1 453
2 73016 1 453
2 73017 1 453
2 73018 1 453
2 73019 1 453
2 73020 1 453
2 73021 1 453
2 73022 1 453
2 73023 1 453
2 73024 1 453
2 73025 1 453
2 73026 1 454
2 73027 1 454
2 73028 1 454
2 73029 1 454
2 73030 1 454
2 73031 1 454
2 73032 1 454
2 73033 1 454
2 73034 1 454
2 73035 1 454
2 73036 1 454
2 73037 1 454
2 73038 1 454
2 73039 1 454
2 73040 1 454
2 73041 1 454
2 73042 1 454
2 73043 1 454
2 73044 1 454
2 73045 1 454
2 73046 1 454
2 73047 1 454
2 73048 1 454
2 73049 1 454
2 73050 1 454
2 73051 1 454
2 73052 1 454
2 73053 1 454
2 73054 1 454
2 73055 1 455
2 73056 1 455
2 73057 1 455
2 73058 1 457
2 73059 1 457
2 73060 1 457
2 73061 1 457
2 73062 1 457
2 73063 1 458
2 73064 1 458
2 73065 1 458
2 73066 1 459
2 73067 1 459
2 73068 1 459
2 73069 1 460
2 73070 1 460
2 73071 1 462
2 73072 1 462
2 73073 1 462
2 73074 1 470
2 73075 1 470
2 73076 1 470
2 73077 1 470
2 73078 1 472
2 73079 1 472
2 73080 1 472
2 73081 1 472
2 73082 1 472
2 73083 1 472
2 73084 1 472
2 73085 1 472
2 73086 1 472
2 73087 1 472
2 73088 1 472
2 73089 1 472
2 73090 1 472
2 73091 1 472
2 73092 1 472
2 73093 1 472
2 73094 1 472
2 73095 1 472
2 73096 1 472
2 73097 1 472
2 73098 1 472
2 73099 1 472
2 73100 1 472
2 73101 1 472
2 73102 1 472
2 73103 1 472
2 73104 1 472
2 73105 1 472
2 73106 1 472
2 73107 1 472
2 73108 1 472
2 73109 1 472
2 73110 1 472
2 73111 1 472
2 73112 1 472
2 73113 1 472
2 73114 1 472
2 73115 1 472
2 73116 1 472
2 73117 1 472
2 73118 1 472
2 73119 1 472
2 73120 1 472
2 73121 1 473
2 73122 1 473
2 73123 1 473
2 73124 1 473
2 73125 1 473
2 73126 1 473
2 73127 1 473
2 73128 1 473
2 73129 1 473
2 73130 1 473
2 73131 1 473
2 73132 1 473
2 73133 1 473
2 73134 1 473
2 73135 1 473
2 73136 1 473
2 73137 1 473
2 73138 1 473
2 73139 1 473
2 73140 1 474
2 73141 1 474
2 73142 1 474
2 73143 1 474
2 73144 1 475
2 73145 1 475
2 73146 1 476
2 73147 1 476
2 73148 1 480
2 73149 1 480
2 73150 1 487
2 73151 1 487
2 73152 1 487
2 73153 1 487
2 73154 1 487
2 73155 1 487
2 73156 1 487
2 73157 1 487
2 73158 1 487
2 73159 1 487
2 73160 1 487
2 73161 1 487
2 73162 1 487
2 73163 1 487
2 73164 1 487
2 73165 1 487
2 73166 1 487
2 73167 1 487
2 73168 1 487
2 73169 1 487
2 73170 1 487
2 73171 1 487
2 73172 1 488
2 73173 1 488
2 73174 1 488
2 73175 1 488
2 73176 1 488
2 73177 1 488
2 73178 1 488
2 73179 1 488
2 73180 1 488
2 73181 1 488
2 73182 1 488
2 73183 1 489
2 73184 1 489
2 73185 1 489
2 73186 1 489
2 73187 1 489
2 73188 1 489
2 73189 1 489
2 73190 1 489
2 73191 1 489
2 73192 1 489
2 73193 1 489
2 73194 1 489
2 73195 1 489
2 73196 1 489
2 73197 1 489
2 73198 1 489
2 73199 1 490
2 73200 1 490
2 73201 1 490
2 73202 1 490
2 73203 1 490
2 73204 1 490
2 73205 1 490
2 73206 1 490
2 73207 1 490
2 73208 1 490
2 73209 1 490
2 73210 1 490
2 73211 1 490
2 73212 1 490
2 73213 1 490
2 73214 1 490
2 73215 1 490
2 73216 1 490
2 73217 1 490
2 73218 1 490
2 73219 1 490
2 73220 1 490
2 73221 1 491
2 73222 1 491
2 73223 1 491
2 73224 1 491
2 73225 1 491
2 73226 1 491
2 73227 1 491
2 73228 1 491
2 73229 1 491
2 73230 1 491
2 73231 1 491
2 73232 1 492
2 73233 1 492
2 73234 1 492
2 73235 1 492
2 73236 1 492
2 73237 1 493
2 73238 1 493
2 73239 1 493
2 73240 1 493
2 73241 1 494
2 73242 1 494
2 73243 1 494
2 73244 1 494
2 73245 1 495
2 73246 1 495
2 73247 1 495
2 73248 1 495
2 73249 1 495
2 73250 1 495
2 73251 1 495
2 73252 1 495
2 73253 1 495
2 73254 1 496
2 73255 1 496
2 73256 1 496
2 73257 1 496
2 73258 1 496
2 73259 1 496
2 73260 1 496
2 73261 1 496
2 73262 1 497
2 73263 1 497
2 73264 1 497
2 73265 1 498
2 73266 1 498
2 73267 1 504
2 73268 1 504
2 73269 1 505
2 73270 1 505
2 73271 1 506
2 73272 1 506
2 73273 1 506
2 73274 1 506
2 73275 1 506
2 73276 1 507
2 73277 1 507
2 73278 1 507
2 73279 1 507
2 73280 1 507
2 73281 1 507
2 73282 1 507
2 73283 1 508
2 73284 1 508
2 73285 1 508
2 73286 1 508
2 73287 1 508
2 73288 1 508
2 73289 1 508
2 73290 1 509
2 73291 1 509
2 73292 1 509
2 73293 1 509
2 73294 1 510
2 73295 1 510
2 73296 1 510
2 73297 1 510
2 73298 1 511
2 73299 1 511
2 73300 1 511
2 73301 1 511
2 73302 1 511
2 73303 1 511
2 73304 1 511
2 73305 1 513
2 73306 1 513
2 73307 1 513
2 73308 1 513
2 73309 1 514
2 73310 1 514
2 73311 1 514
2 73312 1 515
2 73313 1 515
2 73314 1 515
2 73315 1 516
2 73316 1 516
2 73317 1 516
2 73318 1 516
2 73319 1 516
2 73320 1 516
2 73321 1 516
2 73322 1 516
2 73323 1 516
2 73324 1 516
2 73325 1 516
2 73326 1 516
2 73327 1 517
2 73328 1 517
2 73329 1 517
2 73330 1 517
2 73331 1 517
2 73332 1 517
2 73333 1 517
2 73334 1 517
2 73335 1 517
2 73336 1 517
2 73337 1 517
2 73338 1 517
2 73339 1 521
2 73340 1 521
2 73341 1 524
2 73342 1 524
2 73343 1 524
2 73344 1 524
2 73345 1 524
2 73346 1 524
2 73347 1 524
2 73348 1 524
2 73349 1 524
2 73350 1 524
2 73351 1 524
2 73352 1 524
2 73353 1 524
2 73354 1 525
2 73355 1 525
2 73356 1 525
2 73357 1 525
2 73358 1 525
2 73359 1 525
2 73360 1 525
2 73361 1 525
2 73362 1 525
2 73363 1 525
2 73364 1 525
2 73365 1 525
2 73366 1 525
2 73367 1 525
2 73368 1 525
2 73369 1 525
2 73370 1 525
2 73371 1 525
2 73372 1 525
2 73373 1 526
2 73374 1 526
2 73375 1 526
2 73376 1 526
2 73377 1 526
2 73378 1 527
2 73379 1 527
2 73380 1 527
2 73381 1 527
2 73382 1 527
2 73383 1 527
2 73384 1 527
2 73385 1 527
2 73386 1 527
2 73387 1 527
2 73388 1 528
2 73389 1 528
2 73390 1 529
2 73391 1 529
2 73392 1 530
2 73393 1 530
2 73394 1 530
2 73395 1 530
2 73396 1 530
2 73397 1 530
2 73398 1 530
2 73399 1 530
2 73400 1 530
2 73401 1 530
2 73402 1 530
2 73403 1 530
2 73404 1 530
2 73405 1 530
2 73406 1 530
2 73407 1 530
2 73408 1 530
2 73409 1 530
2 73410 1 530
2 73411 1 530
2 73412 1 530
2 73413 1 530
2 73414 1 530
2 73415 1 530
2 73416 1 530
2 73417 1 530
2 73418 1 530
2 73419 1 530
2 73420 1 530
2 73421 1 530
2 73422 1 530
2 73423 1 531
2 73424 1 531
2 73425 1 531
2 73426 1 531
2 73427 1 531
2 73428 1 532
2 73429 1 532
2 73430 1 532
2 73431 1 532
2 73432 1 532
2 73433 1 532
2 73434 1 532
2 73435 1 532
2 73436 1 532
2 73437 1 532
2 73438 1 532
2 73439 1 532
2 73440 1 533
2 73441 1 533
2 73442 1 534
2 73443 1 534
2 73444 1 534
2 73445 1 534
2 73446 1 534
2 73447 1 534
2 73448 1 534
2 73449 1 534
2 73450 1 534
2 73451 1 534
2 73452 1 534
2 73453 1 535
2 73454 1 535
2 73455 1 536
2 73456 1 536
2 73457 1 536
2 73458 1 536
2 73459 1 537
2 73460 1 537
2 73461 1 537
2 73462 1 537
2 73463 1 537
2 73464 1 544
2 73465 1 544
2 73466 1 544
2 73467 1 544
2 73468 1 544
2 73469 1 544
2 73470 1 544
2 73471 1 568
2 73472 1 568
2 73473 1 568
2 73474 1 568
2 73475 1 568
2 73476 1 568
2 73477 1 568
2 73478 1 568
2 73479 1 568
2 73480 1 568
2 73481 1 568
2 73482 1 568
2 73483 1 568
2 73484 1 568
2 73485 1 568
2 73486 1 568
2 73487 1 568
2 73488 1 568
2 73489 1 568
2 73490 1 568
2 73491 1 568
2 73492 1 569
2 73493 1 569
2 73494 1 569
2 73495 1 569
2 73496 1 570
2 73497 1 570
2 73498 1 570
2 73499 1 570
2 73500 1 570
2 73501 1 570
2 73502 1 570
2 73503 1 570
2 73504 1 570
2 73505 1 570
2 73506 1 570
2 73507 1 570
2 73508 1 570
2 73509 1 570
2 73510 1 570
2 73511 1 570
2 73512 1 570
2 73513 1 571
2 73514 1 571
2 73515 1 571
2 73516 1 571
2 73517 1 571
2 73518 1 571
2 73519 1 571
2 73520 1 571
2 73521 1 571
2 73522 1 571
2 73523 1 571
2 73524 1 571
2 73525 1 571
2 73526 1 571
2 73527 1 571
2 73528 1 571
2 73529 1 571
2 73530 1 571
2 73531 1 571
2 73532 1 572
2 73533 1 572
2 73534 1 572
2 73535 1 572
2 73536 1 572
2 73537 1 572
2 73538 1 573
2 73539 1 573
2 73540 1 577
2 73541 1 577
2 73542 1 578
2 73543 1 578
2 73544 1 578
2 73545 1 578
2 73546 1 579
2 73547 1 579
2 73548 1 579
2 73549 1 579
2 73550 1 579
2 73551 1 579
2 73552 1 579
2 73553 1 580
2 73554 1 580
2 73555 1 580
2 73556 1 580
2 73557 1 580
2 73558 1 580
2 73559 1 580
2 73560 1 580
2 73561 1 580
2 73562 1 580
2 73563 1 580
2 73564 1 580
2 73565 1 580
2 73566 1 580
2 73567 1 580
2 73568 1 580
2 73569 1 580
2 73570 1 580
2 73571 1 580
2 73572 1 580
2 73573 1 580
2 73574 1 580
2 73575 1 580
2 73576 1 580
2 73577 1 580
2 73578 1 580
2 73579 1 580
2 73580 1 580
2 73581 1 580
2 73582 1 581
2 73583 1 581
2 73584 1 581
2 73585 1 582
2 73586 1 582
2 73587 1 582
2 73588 1 590
2 73589 1 590
2 73590 1 590
2 73591 1 590
2 73592 1 590
2 73593 1 592
2 73594 1 592
2 73595 1 592
2 73596 1 593
2 73597 1 593
2 73598 1 593
2 73599 1 593
2 73600 1 593
2 73601 1 593
2 73602 1 593
2 73603 1 593
2 73604 1 593
2 73605 1 593
2 73606 1 593
2 73607 1 593
2 73608 1 593
2 73609 1 593
2 73610 1 593
2 73611 1 593
2 73612 1 593
2 73613 1 593
2 73614 1 593
2 73615 1 593
2 73616 1 593
2 73617 1 593
2 73618 1 593
2 73619 1 593
2 73620 1 594
2 73621 1 594
2 73622 1 594
2 73623 1 594
2 73624 1 594
2 73625 1 594
2 73626 1 594
2 73627 1 595
2 73628 1 595
2 73629 1 595
2 73630 1 595
2 73631 1 598
2 73632 1 598
2 73633 1 608
2 73634 1 608
2 73635 1 609
2 73636 1 609
2 73637 1 609
2 73638 1 609
2 73639 1 610
2 73640 1 610
2 73641 1 610
2 73642 1 610
2 73643 1 610
2 73644 1 610
2 73645 1 611
2 73646 1 611
2 73647 1 611
2 73648 1 613
2 73649 1 613
2 73650 1 613
2 73651 1 613
2 73652 1 613
2 73653 1 614
2 73654 1 614
2 73655 1 614
2 73656 1 614
2 73657 1 614
2 73658 1 614
2 73659 1 614
2 73660 1 614
2 73661 1 614
2 73662 1 614
2 73663 1 614
2 73664 1 614
2 73665 1 614
2 73666 1 614
2 73667 1 614
2 73668 1 614
2 73669 1 614
2 73670 1 614
2 73671 1 614
2 73672 1 614
2 73673 1 615
2 73674 1 615
2 73675 1 615
2 73676 1 615
2 73677 1 615
2 73678 1 616
2 73679 1 616
2 73680 1 617
2 73681 1 617
2 73682 1 617
2 73683 1 617
2 73684 1 617
2 73685 1 617
2 73686 1 617
2 73687 1 617
2 73688 1 617
2 73689 1 617
2 73690 1 617
2 73691 1 617
2 73692 1 618
2 73693 1 618
2 73694 1 618
2 73695 1 625
2 73696 1 625
2 73697 1 625
2 73698 1 625
2 73699 1 625
2 73700 1 626
2 73701 1 626
2 73702 1 626
2 73703 1 626
2 73704 1 626
2 73705 1 626
2 73706 1 626
2 73707 1 626
2 73708 1 626
2 73709 1 626
2 73710 1 626
2 73711 1 626
2 73712 1 626
2 73713 1 626
2 73714 1 626
2 73715 1 626
2 73716 1 626
2 73717 1 626
2 73718 1 626
2 73719 1 630
2 73720 1 630
2 73721 1 630
2 73722 1 631
2 73723 1 631
2 73724 1 631
2 73725 1 631
2 73726 1 632
2 73727 1 632
2 73728 1 632
2 73729 1 632
2 73730 1 632
2 73731 1 632
2 73732 1 632
2 73733 1 633
2 73734 1 633
2 73735 1 639
2 73736 1 639
2 73737 1 639
2 73738 1 639
2 73739 1 639
2 73740 1 639
2 73741 1 639
2 73742 1 639
2 73743 1 639
2 73744 1 639
2 73745 1 639
2 73746 1 640
2 73747 1 640
2 73748 1 640
2 73749 1 640
2 73750 1 640
2 73751 1 640
2 73752 1 641
2 73753 1 641
2 73754 1 647
2 73755 1 647
2 73756 1 647
2 73757 1 647
2 73758 1 647
2 73759 1 647
2 73760 1 647
2 73761 1 647
2 73762 1 647
2 73763 1 647
2 73764 1 648
2 73765 1 648
2 73766 1 649
2 73767 1 649
2 73768 1 649
2 73769 1 649
2 73770 1 649
2 73771 1 650
2 73772 1 650
2 73773 1 650
2 73774 1 653
2 73775 1 653
2 73776 1 653
2 73777 1 653
2 73778 1 653
2 73779 1 653
2 73780 1 653
2 73781 1 653
2 73782 1 653
2 73783 1 653
2 73784 1 653
2 73785 1 653
2 73786 1 653
2 73787 1 653
2 73788 1 653
2 73789 1 653
2 73790 1 653
2 73791 1 653
2 73792 1 653
2 73793 1 653
2 73794 1 653
2 73795 1 653
2 73796 1 653
2 73797 1 653
2 73798 1 653
2 73799 1 653
2 73800 1 653
2 73801 1 653
2 73802 1 654
2 73803 1 654
2 73804 1 654
2 73805 1 654
2 73806 1 654
2 73807 1 654
2 73808 1 654
2 73809 1 654
2 73810 1 654
2 73811 1 654
2 73812 1 654
2 73813 1 654
2 73814 1 654
2 73815 1 654
2 73816 1 654
2 73817 1 654
2 73818 1 654
2 73819 1 654
2 73820 1 654
2 73821 1 654
2 73822 1 654
2 73823 1 654
2 73824 1 654
2 73825 1 654
2 73826 1 654
2 73827 1 654
2 73828 1 654
2 73829 1 654
2 73830 1 654
2 73831 1 654
2 73832 1 654
2 73833 1 654
2 73834 1 656
2 73835 1 656
2 73836 1 656
2 73837 1 656
2 73838 1 656
2 73839 1 656
2 73840 1 656
2 73841 1 656
2 73842 1 656
2 73843 1 656
2 73844 1 657
2 73845 1 657
2 73846 1 658
2 73847 1 658
2 73848 1 658
2 73849 1 658
2 73850 1 658
2 73851 1 658
2 73852 1 658
2 73853 1 658
2 73854 1 658
2 73855 1 659
2 73856 1 659
2 73857 1 661
2 73858 1 661
2 73859 1 661
2 73860 1 661
2 73861 1 661
2 73862 1 661
2 73863 1 661
2 73864 1 661
2 73865 1 661
2 73866 1 661
2 73867 1 661
2 73868 1 661
2 73869 1 661
2 73870 1 661
2 73871 1 661
2 73872 1 661
2 73873 1 661
2 73874 1 661
2 73875 1 661
2 73876 1 661
2 73877 1 661
2 73878 1 661
2 73879 1 661
2 73880 1 661
2 73881 1 661
2 73882 1 661
2 73883 1 661
2 73884 1 662
2 73885 1 662
2 73886 1 663
2 73887 1 663
2 73888 1 663
2 73889 1 663
2 73890 1 663
2 73891 1 663
2 73892 1 663
2 73893 1 663
2 73894 1 663
2 73895 1 663
2 73896 1 663
2 73897 1 663
2 73898 1 665
2 73899 1 665
2 73900 1 665
2 73901 1 665
2 73902 1 665
2 73903 1 665
2 73904 1 665
2 73905 1 665
2 73906 1 665
2 73907 1 665
2 73908 1 665
2 73909 1 665
2 73910 1 665
2 73911 1 665
2 73912 1 665
2 73913 1 665
2 73914 1 665
2 73915 1 665
2 73916 1 665
2 73917 1 665
2 73918 1 665
2 73919 1 666
2 73920 1 666
2 73921 1 667
2 73922 1 667
2 73923 1 667
2 73924 1 667
2 73925 1 667
2 73926 1 668
2 73927 1 668
2 73928 1 668
2 73929 1 668
2 73930 1 680
2 73931 1 680
2 73932 1 681
2 73933 1 681
2 73934 1 681
2 73935 1 681
2 73936 1 685
2 73937 1 685
2 73938 1 686
2 73939 1 686
2 73940 1 687
2 73941 1 687
2 73942 1 695
2 73943 1 695
2 73944 1 695
2 73945 1 695
2 73946 1 695
2 73947 1 695
2 73948 1 695
2 73949 1 695
2 73950 1 695
2 73951 1 695
2 73952 1 695
2 73953 1 695
2 73954 1 695
2 73955 1 695
2 73956 1 695
2 73957 1 696
2 73958 1 696
2 73959 1 696
2 73960 1 696
2 73961 1 696
2 73962 1 696
2 73963 1 696
2 73964 1 697
2 73965 1 697
2 73966 1 705
2 73967 1 705
2 73968 1 705
2 73969 1 705
2 73970 1 705
2 73971 1 705
2 73972 1 705
2 73973 1 705
2 73974 1 706
2 73975 1 706
2 73976 1 706
2 73977 1 706
2 73978 1 707
2 73979 1 707
2 73980 1 707
2 73981 1 707
2 73982 1 707
2 73983 1 707
2 73984 1 709
2 73985 1 709
2 73986 1 710
2 73987 1 710
2 73988 1 710
2 73989 1 710
2 73990 1 710
2 73991 1 711
2 73992 1 711
2 73993 1 711
2 73994 1 711
2 73995 1 714
2 73996 1 714
2 73997 1 714
2 73998 1 714
2 73999 1 714
2 74000 1 714
2 74001 1 714
2 74002 1 714
2 74003 1 715
2 74004 1 715
2 74005 1 715
2 74006 1 715
2 74007 1 715
2 74008 1 715
2 74009 1 715
2 74010 1 715
2 74011 1 715
2 74012 1 715
2 74013 1 715
2 74014 1 715
2 74015 1 715
2 74016 1 715
2 74017 1 715
2 74018 1 715
2 74019 1 715
2 74020 1 715
2 74021 1 715
2 74022 1 715
2 74023 1 715
2 74024 1 715
2 74025 1 715
2 74026 1 715
2 74027 1 715
2 74028 1 715
2 74029 1 715
2 74030 1 715
2 74031 1 715
2 74032 1 715
2 74033 1 715
2 74034 1 715
2 74035 1 715
2 74036 1 715
2 74037 1 715
2 74038 1 715
2 74039 1 716
2 74040 1 716
2 74041 1 716
2 74042 1 716
2 74043 1 716
2 74044 1 716
2 74045 1 716
2 74046 1 716
2 74047 1 716
2 74048 1 717
2 74049 1 717
2 74050 1 717
2 74051 1 717
2 74052 1 717
2 74053 1 717
2 74054 1 717
2 74055 1 717
2 74056 1 717
2 74057 1 717
2 74058 1 717
2 74059 1 717
2 74060 1 717
2 74061 1 717
2 74062 1 717
2 74063 1 717
2 74064 1 717
2 74065 1 717
2 74066 1 717
2 74067 1 717
2 74068 1 717
2 74069 1 717
2 74070 1 717
2 74071 1 717
2 74072 1 717
2 74073 1 717
2 74074 1 717
2 74075 1 717
2 74076 1 717
2 74077 1 717
2 74078 1 717
2 74079 1 717
2 74080 1 718
2 74081 1 718
2 74082 1 718
2 74083 1 722
2 74084 1 722
2 74085 1 722
2 74086 1 722
2 74087 1 722
2 74088 1 722
2 74089 1 722
2 74090 1 722
2 74091 1 722
2 74092 1 722
2 74093 1 722
2 74094 1 722
2 74095 1 722
2 74096 1 722
2 74097 1 722
2 74098 1 722
2 74099 1 722
2 74100 1 722
2 74101 1 722
2 74102 1 722
2 74103 1 722
2 74104 1 722
2 74105 1 722
2 74106 1 722
2 74107 1 723
2 74108 1 723
2 74109 1 723
2 74110 1 723
2 74111 1 723
2 74112 1 723
2 74113 1 723
2 74114 1 723
2 74115 1 723
2 74116 1 723
2 74117 1 723
2 74118 1 723
2 74119 1 723
2 74120 1 723
2 74121 1 723
2 74122 1 723
2 74123 1 723
2 74124 1 723
2 74125 1 723
2 74126 1 723
2 74127 1 724
2 74128 1 724
2 74129 1 724
2 74130 1 724
2 74131 1 724
2 74132 1 724
2 74133 1 724
2 74134 1 725
2 74135 1 725
2 74136 1 725
2 74137 1 725
2 74138 1 725
2 74139 1 725
2 74140 1 725
2 74141 1 725
2 74142 1 729
2 74143 1 729
2 74144 1 729
2 74145 1 729
2 74146 1 729
2 74147 1 729
2 74148 1 729
2 74149 1 729
2 74150 1 729
2 74151 1 729
2 74152 1 729
2 74153 1 729
2 74154 1 729
2 74155 1 729
2 74156 1 730
2 74157 1 730
2 74158 1 731
2 74159 1 731
2 74160 1 732
2 74161 1 732
2 74162 1 732
2 74163 1 732
2 74164 1 732
2 74165 1 733
2 74166 1 733
2 74167 1 734
2 74168 1 734
2 74169 1 737
2 74170 1 737
2 74171 1 738
2 74172 1 738
2 74173 1 738
2 74174 1 738
2 74175 1 739
2 74176 1 739
2 74177 1 739
2 74178 1 740
2 74179 1 740
2 74180 1 740
2 74181 1 740
2 74182 1 740
2 74183 1 740
2 74184 1 740
2 74185 1 740
2 74186 1 740
2 74187 1 740
2 74188 1 740
2 74189 1 740
2 74190 1 741
2 74191 1 741
2 74192 1 742
2 74193 1 742
2 74194 1 751
2 74195 1 751
2 74196 1 751
2 74197 1 751
2 74198 1 751
2 74199 1 751
2 74200 1 751
2 74201 1 751
2 74202 1 751
2 74203 1 751
2 74204 1 751
2 74205 1 751
2 74206 1 751
2 74207 1 751
2 74208 1 752
2 74209 1 752
2 74210 1 752
2 74211 1 752
2 74212 1 760
2 74213 1 760
2 74214 1 760
2 74215 1 760
2 74216 1 760
2 74217 1 760
2 74218 1 760
2 74219 1 760
2 74220 1 760
2 74221 1 760
2 74222 1 760
2 74223 1 760
2 74224 1 760
2 74225 1 760
2 74226 1 760
2 74227 1 760
2 74228 1 761
2 74229 1 761
2 74230 1 761
2 74231 1 761
2 74232 1 761
2 74233 1 762
2 74234 1 762
2 74235 1 763
2 74236 1 763
2 74237 1 766
2 74238 1 766
2 74239 1 766
2 74240 1 767
2 74241 1 767
2 74242 1 771
2 74243 1 771
2 74244 1 773
2 74245 1 773
2 74246 1 773
2 74247 1 773
2 74248 1 773
2 74249 1 773
2 74250 1 773
2 74251 1 774
2 74252 1 774
2 74253 1 775
2 74254 1 775
2 74255 1 781
2 74256 1 781
2 74257 1 781
2 74258 1 782
2 74259 1 782
2 74260 1 782
2 74261 1 782
2 74262 1 782
2 74263 1 782
2 74264 1 782
2 74265 1 782
2 74266 1 783
2 74267 1 783
2 74268 1 796
2 74269 1 796
2 74270 1 797
2 74271 1 797
2 74272 1 797
2 74273 1 797
2 74274 1 797
2 74275 1 797
2 74276 1 797
2 74277 1 797
2 74278 1 797
2 74279 1 797
2 74280 1 797
2 74281 1 797
2 74282 1 797
2 74283 1 797
2 74284 1 797
2 74285 1 798
2 74286 1 798
2 74287 1 798
2 74288 1 799
2 74289 1 799
2 74290 1 800
2 74291 1 800
2 74292 1 800
2 74293 1 800
2 74294 1 801
2 74295 1 801
2 74296 1 803
2 74297 1 803
2 74298 1 803
2 74299 1 803
2 74300 1 803
2 74301 1 806
2 74302 1 806
2 74303 1 808
2 74304 1 808
2 74305 1 808
2 74306 1 808
2 74307 1 808
2 74308 1 808
2 74309 1 808
2 74310 1 809
2 74311 1 809
2 74312 1 811
2 74313 1 811
2 74314 1 811
2 74315 1 811
2 74316 1 815
2 74317 1 815
2 74318 1 816
2 74319 1 816
2 74320 1 816
2 74321 1 817
2 74322 1 817
2 74323 1 817
2 74324 1 817
2 74325 1 817
2 74326 1 817
2 74327 1 817
2 74328 1 820
2 74329 1 820
2 74330 1 820
2 74331 1 820
2 74332 1 820
2 74333 1 820
2 74334 1 820
2 74335 1 820
2 74336 1 820
2 74337 1 820
2 74338 1 820
2 74339 1 820
2 74340 1 820
2 74341 1 820
2 74342 1 820
2 74343 1 820
2 74344 1 820
2 74345 1 820
2 74346 1 820
2 74347 1 822
2 74348 1 822
2 74349 1 822
2 74350 1 822
2 74351 1 823
2 74352 1 823
2 74353 1 823
2 74354 1 823
2 74355 1 824
2 74356 1 824
2 74357 1 824
2 74358 1 824
2 74359 1 824
2 74360 1 824
2 74361 1 824
2 74362 1 824
2 74363 1 824
2 74364 1 824
2 74365 1 824
2 74366 1 824
2 74367 1 824
2 74368 1 824
2 74369 1 824
2 74370 1 824
2 74371 1 824
2 74372 1 824
2 74373 1 825
2 74374 1 825
2 74375 1 827
2 74376 1 827
2 74377 1 828
2 74378 1 828
2 74379 1 835
2 74380 1 835
2 74381 1 835
2 74382 1 835
2 74383 1 835
2 74384 1 836
2 74385 1 836
2 74386 1 836
2 74387 1 837
2 74388 1 837
2 74389 1 837
2 74390 1 837
2 74391 1 837
2 74392 1 837
2 74393 1 837
2 74394 1 837
2 74395 1 837
2 74396 1 837
2 74397 1 837
2 74398 1 837
2 74399 1 837
2 74400 1 837
2 74401 1 837
2 74402 1 837
2 74403 1 837
2 74404 1 837
2 74405 1 837
2 74406 1 838
2 74407 1 838
2 74408 1 838
2 74409 1 839
2 74410 1 839
2 74411 1 839
2 74412 1 839
2 74413 1 840
2 74414 1 840
2 74415 1 840
2 74416 1 840
2 74417 1 841
2 74418 1 841
2 74419 1 841
2 74420 1 841
2 74421 1 841
2 74422 1 842
2 74423 1 842
2 74424 1 842
2 74425 1 844
2 74426 1 844
2 74427 1 844
2 74428 1 849
2 74429 1 849
2 74430 1 849
2 74431 1 849
2 74432 1 849
2 74433 1 850
2 74434 1 850
2 74435 1 850
2 74436 1 850
2 74437 1 850
2 74438 1 851
2 74439 1 851
2 74440 1 853
2 74441 1 853
2 74442 1 854
2 74443 1 854
2 74444 1 855
2 74445 1 855
2 74446 1 855
2 74447 1 864
2 74448 1 864
2 74449 1 864
2 74450 1 864
2 74451 1 864
2 74452 1 864
2 74453 1 864
2 74454 1 864
2 74455 1 864
2 74456 1 864
2 74457 1 865
2 74458 1 865
2 74459 1 865
2 74460 1 865
2 74461 1 866
2 74462 1 866
2 74463 1 866
2 74464 1 866
2 74465 1 866
2 74466 1 866
2 74467 1 866
2 74468 1 867
2 74469 1 867
2 74470 1 867
2 74471 1 867
2 74472 1 867
2 74473 1 867
2 74474 1 868
2 74475 1 868
2 74476 1 868
2 74477 1 868
2 74478 1 868
2 74479 1 868
2 74480 1 868
2 74481 1 868
2 74482 1 868
2 74483 1 868
2 74484 1 868
2 74485 1 868
2 74486 1 868
2 74487 1 872
2 74488 1 872
2 74489 1 873
2 74490 1 873
2 74491 1 873
2 74492 1 873
2 74493 1 873
2 74494 1 873
2 74495 1 874
2 74496 1 874
2 74497 1 874
2 74498 1 874
2 74499 1 874
2 74500 1 874
2 74501 1 874
2 74502 1 874
2 74503 1 874
2 74504 1 876
2 74505 1 876
2 74506 1 876
2 74507 1 876
2 74508 1 876
2 74509 1 876
2 74510 1 876
2 74511 1 876
2 74512 1 876
2 74513 1 877
2 74514 1 877
2 74515 1 877
2 74516 1 877
2 74517 1 877
2 74518 1 877
2 74519 1 877
2 74520 1 877
2 74521 1 877
2 74522 1 877
2 74523 1 877
2 74524 1 880
2 74525 1 880
2 74526 1 881
2 74527 1 881
2 74528 1 894
2 74529 1 894
2 74530 1 894
2 74531 1 895
2 74532 1 895
2 74533 1 895
2 74534 1 895
2 74535 1 895
2 74536 1 901
2 74537 1 901
2 74538 1 901
2 74539 1 902
2 74540 1 902
2 74541 1 902
2 74542 1 902
2 74543 1 910
2 74544 1 910
2 74545 1 910
2 74546 1 910
2 74547 1 910
2 74548 1 910
2 74549 1 911
2 74550 1 911
2 74551 1 912
2 74552 1 912
2 74553 1 912
2 74554 1 913
2 74555 1 913
2 74556 1 921
2 74557 1 921
2 74558 1 921
2 74559 1 921
2 74560 1 921
2 74561 1 921
2 74562 1 921
2 74563 1 921
2 74564 1 921
2 74565 1 921
2 74566 1 921
2 74567 1 921
2 74568 1 921
2 74569 1 921
2 74570 1 921
2 74571 1 922
2 74572 1 922
2 74573 1 922
2 74574 1 922
2 74575 1 922
2 74576 1 922
2 74577 1 922
2 74578 1 922
2 74579 1 922
2 74580 1 922
2 74581 1 922
2 74582 1 922
2 74583 1 922
2 74584 1 922
2 74585 1 922
2 74586 1 922
2 74587 1 922
2 74588 1 922
2 74589 1 922
2 74590 1 922
2 74591 1 922
2 74592 1 922
2 74593 1 922
2 74594 1 922
2 74595 1 922
2 74596 1 922
2 74597 1 922
2 74598 1 922
2 74599 1 922
2 74600 1 922
2 74601 1 922
2 74602 1 922
2 74603 1 922
2 74604 1 922
2 74605 1 922
2 74606 1 922
2 74607 1 922
2 74608 1 922
2 74609 1 922
2 74610 1 923
2 74611 1 923
2 74612 1 923
2 74613 1 923
2 74614 1 924
2 74615 1 924
2 74616 1 924
2 74617 1 924
2 74618 1 924
2 74619 1 924
2 74620 1 924
2 74621 1 924
2 74622 1 924
2 74623 1 924
2 74624 1 924
2 74625 1 924
2 74626 1 924
2 74627 1 924
2 74628 1 924
2 74629 1 925
2 74630 1 925
2 74631 1 925
2 74632 1 925
2 74633 1 925
2 74634 1 925
2 74635 1 925
2 74636 1 926
2 74637 1 926
2 74638 1 926
2 74639 1 926
2 74640 1 926
2 74641 1 926
2 74642 1 926
2 74643 1 927
2 74644 1 927
2 74645 1 928
2 74646 1 928
2 74647 1 931
2 74648 1 931
2 74649 1 931
2 74650 1 931
2 74651 1 931
2 74652 1 931
2 74653 1 931
2 74654 1 931
2 74655 1 932
2 74656 1 932
2 74657 1 932
2 74658 1 932
2 74659 1 932
2 74660 1 932
2 74661 1 932
2 74662 1 939
2 74663 1 939
2 74664 1 939
2 74665 1 939
2 74666 1 940
2 74667 1 940
2 74668 1 940
2 74669 1 941
2 74670 1 941
2 74671 1 941
2 74672 1 941
2 74673 1 941
2 74674 1 941
2 74675 1 941
2 74676 1 941
2 74677 1 941
2 74678 1 941
2 74679 1 941
2 74680 1 941
2 74681 1 941
2 74682 1 941
2 74683 1 941
2 74684 1 941
2 74685 1 941
2 74686 1 942
2 74687 1 942
2 74688 1 942
2 74689 1 944
2 74690 1 944
2 74691 1 963
2 74692 1 963
2 74693 1 963
2 74694 1 963
2 74695 1 963
2 74696 1 972
2 74697 1 972
2 74698 1 983
2 74699 1 983
2 74700 1 983
2 74701 1 983
2 74702 1 983
2 74703 1 983
2 74704 1 983
2 74705 1 985
2 74706 1 985
2 74707 1 986
2 74708 1 986
2 74709 1 986
2 74710 1 986
2 74711 1 986
2 74712 1 986
2 74713 1 986
2 74714 1 986
2 74715 1 987
2 74716 1 987
2 74717 1 987
2 74718 1 987
2 74719 1 1000
2 74720 1 1000
2 74721 1 1000
2 74722 1 1000
2 74723 1 1000
2 74724 1 1000
2 74725 1 1000
2 74726 1 1000
2 74727 1 1000
2 74728 1 1000
2 74729 1 1000
2 74730 1 1000
2 74731 1 1000
2 74732 1 1000
2 74733 1 1000
2 74734 1 1000
2 74735 1 1000
2 74736 1 1000
2 74737 1 1000
2 74738 1 1000
2 74739 1 1000
2 74740 1 1000
2 74741 1 1001
2 74742 1 1001
2 74743 1 1001
2 74744 1 1001
2 74745 1 1001
2 74746 1 1002
2 74747 1 1002
2 74748 1 1002
2 74749 1 1003
2 74750 1 1003
2 74751 1 1008
2 74752 1 1008
2 74753 1 1008
2 74754 1 1008
2 74755 1 1009
2 74756 1 1009
2 74757 1 1009
2 74758 1 1009
2 74759 1 1009
2 74760 1 1009
2 74761 1 1010
2 74762 1 1010
2 74763 1 1010
2 74764 1 1010
2 74765 1 1011
2 74766 1 1011
2 74767 1 1011
2 74768 1 1011
2 74769 1 1011
2 74770 1 1011
2 74771 1 1011
2 74772 1 1012
2 74773 1 1012
2 74774 1 1016
2 74775 1 1016
2 74776 1 1016
2 74777 1 1016
2 74778 1 1016
2 74779 1 1025
2 74780 1 1025
2 74781 1 1025
2 74782 1 1025
2 74783 1 1025
2 74784 1 1025
2 74785 1 1025
2 74786 1 1025
2 74787 1 1025
2 74788 1 1025
2 74789 1 1026
2 74790 1 1026
2 74791 1 1026
2 74792 1 1026
2 74793 1 1026
2 74794 1 1026
2 74795 1 1026
2 74796 1 1026
2 74797 1 1026
2 74798 1 1026
2 74799 1 1026
2 74800 1 1026
2 74801 1 1026
2 74802 1 1026
2 74803 1 1026
2 74804 1 1026
2 74805 1 1026
2 74806 1 1026
2 74807 1 1026
2 74808 1 1028
2 74809 1 1028
2 74810 1 1028
2 74811 1 1028
2 74812 1 1036
2 74813 1 1036
2 74814 1 1036
2 74815 1 1036
2 74816 1 1036
2 74817 1 1036
2 74818 1 1036
2 74819 1 1036
2 74820 1 1037
2 74821 1 1037
2 74822 1 1037
2 74823 1 1040
2 74824 1 1040
2 74825 1 1040
2 74826 1 1040
2 74827 1 1040
2 74828 1 1040
2 74829 1 1040
2 74830 1 1040
2 74831 1 1041
2 74832 1 1041
2 74833 1 1050
2 74834 1 1050
2 74835 1 1050
2 74836 1 1050
2 74837 1 1050
2 74838 1 1050
2 74839 1 1050
2 74840 1 1051
2 74841 1 1051
2 74842 1 1051
2 74843 1 1052
2 74844 1 1052
2 74845 1 1052
2 74846 1 1052
2 74847 1 1052
2 74848 1 1052
2 74849 1 1052
2 74850 1 1052
2 74851 1 1053
2 74852 1 1053
2 74853 1 1059
2 74854 1 1059
2 74855 1 1059
2 74856 1 1061
2 74857 1 1061
2 74858 1 1062
2 74859 1 1062
2 74860 1 1062
2 74861 1 1062
2 74862 1 1062
2 74863 1 1062
2 74864 1 1062
2 74865 1 1062
2 74866 1 1062
2 74867 1 1062
2 74868 1 1062
2 74869 1 1062
2 74870 1 1063
2 74871 1 1063
2 74872 1 1064
2 74873 1 1064
2 74874 1 1078
2 74875 1 1078
2 74876 1 1083
2 74877 1 1083
2 74878 1 1083
2 74879 1 1083
2 74880 1 1083
2 74881 1 1083
2 74882 1 1083
2 74883 1 1083
2 74884 1 1083
2 74885 1 1083
2 74886 1 1083
2 74887 1 1084
2 74888 1 1084
2 74889 1 1084
2 74890 1 1084
2 74891 1 1084
2 74892 1 1084
2 74893 1 1084
2 74894 1 1084
2 74895 1 1084
2 74896 1 1084
2 74897 1 1084
2 74898 1 1084
2 74899 1 1084
2 74900 1 1084
2 74901 1 1084
2 74902 1 1085
2 74903 1 1085
2 74904 1 1085
2 74905 1 1093
2 74906 1 1093
2 74907 1 1093
2 74908 1 1093
2 74909 1 1093
2 74910 1 1094
2 74911 1 1094
2 74912 1 1094
2 74913 1 1095
2 74914 1 1095
2 74915 1 1095
2 74916 1 1095
2 74917 1 1095
2 74918 1 1095
2 74919 1 1095
2 74920 1 1096
2 74921 1 1096
2 74922 1 1104
2 74923 1 1104
2 74924 1 1104
2 74925 1 1104
2 74926 1 1104
2 74927 1 1104
2 74928 1 1104
2 74929 1 1104
2 74930 1 1104
2 74931 1 1104
2 74932 1 1104
2 74933 1 1104
2 74934 1 1104
2 74935 1 1104
2 74936 1 1104
2 74937 1 1104
2 74938 1 1104
2 74939 1 1106
2 74940 1 1106
2 74941 1 1113
2 74942 1 1113
2 74943 1 1113
2 74944 1 1113
2 74945 1 1113
2 74946 1 1113
2 74947 1 1113
2 74948 1 1113
2 74949 1 1113
2 74950 1 1113
2 74951 1 1113
2 74952 1 1114
2 74953 1 1114
2 74954 1 1115
2 74955 1 1115
2 74956 1 1115
2 74957 1 1116
2 74958 1 1116
2 74959 1 1116
2 74960 1 1116
2 74961 1 1116
2 74962 1 1117
2 74963 1 1117
2 74964 1 1117
2 74965 1 1117
2 74966 1 1117
2 74967 1 1117
2 74968 1 1117
2 74969 1 1117
2 74970 1 1118
2 74971 1 1118
2 74972 1 1118
2 74973 1 1118
2 74974 1 1118
2 74975 1 1118
2 74976 1 1118
2 74977 1 1118
2 74978 1 1118
2 74979 1 1119
2 74980 1 1119
2 74981 1 1127
2 74982 1 1127
2 74983 1 1127
2 74984 1 1127
2 74985 1 1127
2 74986 1 1127
2 74987 1 1127
2 74988 1 1127
2 74989 1 1127
2 74990 1 1127
2 74991 1 1127
2 74992 1 1127
2 74993 1 1127
2 74994 1 1127
2 74995 1 1127
2 74996 1 1127
2 74997 1 1128
2 74998 1 1128
2 74999 1 1128
2 75000 1 1128
2 75001 1 1128
2 75002 1 1128
2 75003 1 1129
2 75004 1 1129
2 75005 1 1129
2 75006 1 1130
2 75007 1 1130
2 75008 1 1130
2 75009 1 1130
2 75010 1 1130
2 75011 1 1130
2 75012 1 1130
2 75013 1 1130
2 75014 1 1130
2 75015 1 1130
2 75016 1 1130
2 75017 1 1130
2 75018 1 1130
2 75019 1 1130
2 75020 1 1130
2 75021 1 1130
2 75022 1 1130
2 75023 1 1130
2 75024 1 1130
2 75025 1 1130
2 75026 1 1130
2 75027 1 1130
2 75028 1 1130
2 75029 1 1130
2 75030 1 1130
2 75031 1 1130
2 75032 1 1130
2 75033 1 1131
2 75034 1 1131
2 75035 1 1131
2 75036 1 1131
2 75037 1 1131
2 75038 1 1131
2 75039 1 1131
2 75040 1 1131
2 75041 1 1131
2 75042 1 1131
2 75043 1 1133
2 75044 1 1133
2 75045 1 1133
2 75046 1 1133
2 75047 1 1133
2 75048 1 1133
2 75049 1 1133
2 75050 1 1133
2 75051 1 1133
2 75052 1 1133
2 75053 1 1133
2 75054 1 1133
2 75055 1 1133
2 75056 1 1133
2 75057 1 1134
2 75058 1 1134
2 75059 1 1138
2 75060 1 1138
2 75061 1 1138
2 75062 1 1138
2 75063 1 1138
2 75064 1 1138
2 75065 1 1138
2 75066 1 1138
2 75067 1 1138
2 75068 1 1138
2 75069 1 1138
2 75070 1 1138
2 75071 1 1138
2 75072 1 1138
2 75073 1 1138
2 75074 1 1138
2 75075 1 1138
2 75076 1 1138
2 75077 1 1138
2 75078 1 1138
2 75079 1 1139
2 75080 1 1139
2 75081 1 1139
2 75082 1 1139
2 75083 1 1146
2 75084 1 1146
2 75085 1 1146
2 75086 1 1147
2 75087 1 1147
2 75088 1 1147
2 75089 1 1148
2 75090 1 1148
2 75091 1 1148
2 75092 1 1148
2 75093 1 1148
2 75094 1 1148
2 75095 1 1148
2 75096 1 1148
2 75097 1 1148
2 75098 1 1148
2 75099 1 1148
2 75100 1 1148
2 75101 1 1148
2 75102 1 1156
2 75103 1 1156
2 75104 1 1156
2 75105 1 1156
2 75106 1 1156
2 75107 1 1156
2 75108 1 1156
2 75109 1 1156
2 75110 1 1156
2 75111 1 1156
2 75112 1 1156
2 75113 1 1156
2 75114 1 1156
2 75115 1 1156
2 75116 1 1156
2 75117 1 1156
2 75118 1 1156
2 75119 1 1156
2 75120 1 1156
2 75121 1 1156
2 75122 1 1156
2 75123 1 1156
2 75124 1 1157
2 75125 1 1157
2 75126 1 1157
2 75127 1 1157
2 75128 1 1157
2 75129 1 1157
2 75130 1 1158
2 75131 1 1158
2 75132 1 1167
2 75133 1 1167
2 75134 1 1167
2 75135 1 1167
2 75136 1 1167
2 75137 1 1167
2 75138 1 1167
2 75139 1 1167
2 75140 1 1167
2 75141 1 1167
2 75142 1 1167
2 75143 1 1167
2 75144 1 1167
2 75145 1 1167
2 75146 1 1168
2 75147 1 1168
2 75148 1 1168
2 75149 1 1168
2 75150 1 1168
2 75151 1 1168
2 75152 1 1168
2 75153 1 1168
2 75154 1 1169
2 75155 1 1169
2 75156 1 1172
2 75157 1 1172
2 75158 1 1172
2 75159 1 1172
2 75160 1 1172
2 75161 1 1172
2 75162 1 1172
2 75163 1 1172
2 75164 1 1172
2 75165 1 1172
2 75166 1 1172
2 75167 1 1172
2 75168 1 1172
2 75169 1 1172
2 75170 1 1172
2 75171 1 1172
2 75172 1 1172
2 75173 1 1172
2 75174 1 1172
2 75175 1 1172
2 75176 1 1172
2 75177 1 1172
2 75178 1 1172
2 75179 1 1172
2 75180 1 1172
2 75181 1 1172
2 75182 1 1172
2 75183 1 1172
2 75184 1 1172
2 75185 1 1172
2 75186 1 1172
2 75187 1 1172
2 75188 1 1172
2 75189 1 1172
2 75190 1 1172
2 75191 1 1172
2 75192 1 1172
2 75193 1 1172
2 75194 1 1172
2 75195 1 1172
2 75196 1 1172
2 75197 1 1172
2 75198 1 1172
2 75199 1 1172
2 75200 1 1172
2 75201 1 1172
2 75202 1 1172
2 75203 1 1172
2 75204 1 1172
2 75205 1 1172
2 75206 1 1172
2 75207 1 1172
2 75208 1 1172
2 75209 1 1172
2 75210 1 1172
2 75211 1 1172
2 75212 1 1172
2 75213 1 1172
2 75214 1 1172
2 75215 1 1172
2 75216 1 1172
2 75217 1 1172
2 75218 1 1172
2 75219 1 1172
2 75220 1 1172
2 75221 1 1172
2 75222 1 1172
2 75223 1 1172
2 75224 1 1172
2 75225 1 1172
2 75226 1 1172
2 75227 1 1172
2 75228 1 1172
2 75229 1 1172
2 75230 1 1172
2 75231 1 1172
2 75232 1 1172
2 75233 1 1172
2 75234 1 1172
2 75235 1 1172
2 75236 1 1172
2 75237 1 1172
2 75238 1 1172
2 75239 1 1172
2 75240 1 1172
2 75241 1 1172
2 75242 1 1172
2 75243 1 1172
2 75244 1 1173
2 75245 1 1173
2 75246 1 1173
2 75247 1 1173
2 75248 1 1173
2 75249 1 1173
2 75250 1 1173
2 75251 1 1173
2 75252 1 1173
2 75253 1 1173
2 75254 1 1173
2 75255 1 1173
2 75256 1 1173
2 75257 1 1173
2 75258 1 1173
2 75259 1 1173
2 75260 1 1173
2 75261 1 1173
2 75262 1 1173
2 75263 1 1173
2 75264 1 1173
2 75265 1 1173
2 75266 1 1173
2 75267 1 1173
2 75268 1 1173
2 75269 1 1173
2 75270 1 1173
2 75271 1 1173
2 75272 1 1173
2 75273 1 1173
2 75274 1 1173
2 75275 1 1173
2 75276 1 1173
2 75277 1 1173
2 75278 1 1173
2 75279 1 1173
2 75280 1 1173
2 75281 1 1173
2 75282 1 1173
2 75283 1 1173
2 75284 1 1173
2 75285 1 1173
2 75286 1 1173
2 75287 1 1173
2 75288 1 1173
2 75289 1 1173
2 75290 1 1173
2 75291 1 1173
2 75292 1 1173
2 75293 1 1173
2 75294 1 1173
2 75295 1 1173
2 75296 1 1173
2 75297 1 1173
2 75298 1 1173
2 75299 1 1173
2 75300 1 1173
2 75301 1 1173
2 75302 1 1173
2 75303 1 1173
2 75304 1 1173
2 75305 1 1173
2 75306 1 1173
2 75307 1 1173
2 75308 1 1173
2 75309 1 1173
2 75310 1 1173
2 75311 1 1173
2 75312 1 1173
2 75313 1 1173
2 75314 1 1173
2 75315 1 1173
2 75316 1 1173
2 75317 1 1173
2 75318 1 1173
2 75319 1 1173
2 75320 1 1173
2 75321 1 1173
2 75322 1 1173
2 75323 1 1173
2 75324 1 1173
2 75325 1 1173
2 75326 1 1173
2 75327 1 1173
2 75328 1 1173
2 75329 1 1173
2 75330 1 1173
2 75331 1 1173
2 75332 1 1173
2 75333 1 1173
2 75334 1 1173
2 75335 1 1173
2 75336 1 1173
2 75337 1 1173
2 75338 1 1173
2 75339 1 1173
2 75340 1 1173
2 75341 1 1173
2 75342 1 1173
2 75343 1 1173
2 75344 1 1173
2 75345 1 1173
2 75346 1 1173
2 75347 1 1173
2 75348 1 1173
2 75349 1 1173
2 75350 1 1173
2 75351 1 1173
2 75352 1 1173
2 75353 1 1173
2 75354 1 1173
2 75355 1 1173
2 75356 1 1173
2 75357 1 1173
2 75358 1 1173
2 75359 1 1173
2 75360 1 1173
2 75361 1 1173
2 75362 1 1173
2 75363 1 1173
2 75364 1 1173
2 75365 1 1173
2 75366 1 1173
2 75367 1 1173
2 75368 1 1173
2 75369 1 1173
2 75370 1 1173
2 75371 1 1173
2 75372 1 1173
2 75373 1 1173
2 75374 1 1173
2 75375 1 1173
2 75376 1 1173
2 75377 1 1173
2 75378 1 1173
2 75379 1 1173
2 75380 1 1173
2 75381 1 1173
2 75382 1 1173
2 75383 1 1174
2 75384 1 1174
2 75385 1 1174
2 75386 1 1174
2 75387 1 1174
2 75388 1 1174
2 75389 1 1174
2 75390 1 1174
2 75391 1 1174
2 75392 1 1174
2 75393 1 1174
2 75394 1 1174
2 75395 1 1174
2 75396 1 1174
2 75397 1 1174
2 75398 1 1174
2 75399 1 1174
2 75400 1 1174
2 75401 1 1174
2 75402 1 1174
2 75403 1 1175
2 75404 1 1175
2 75405 1 1175
2 75406 1 1175
2 75407 1 1176
2 75408 1 1176
2 75409 1 1176
2 75410 1 1176
2 75411 1 1176
2 75412 1 1176
2 75413 1 1176
2 75414 1 1176
2 75415 1 1176
2 75416 1 1176
2 75417 1 1176
2 75418 1 1176
2 75419 1 1176
2 75420 1 1176
2 75421 1 1176
2 75422 1 1176
2 75423 1 1176
2 75424 1 1177
2 75425 1 1177
2 75426 1 1177
2 75427 1 1177
2 75428 1 1177
2 75429 1 1178
2 75430 1 1178
2 75431 1 1178
2 75432 1 1178
2 75433 1 1178
2 75434 1 1178
2 75435 1 1178
2 75436 1 1178
2 75437 1 1178
2 75438 1 1178
2 75439 1 1178
2 75440 1 1178
2 75441 1 1178
2 75442 1 1178
2 75443 1 1178
2 75444 1 1178
2 75445 1 1178
2 75446 1 1178
2 75447 1 1178
2 75448 1 1180
2 75449 1 1180
2 75450 1 1180
2 75451 1 1180
2 75452 1 1189
2 75453 1 1189
2 75454 1 1191
2 75455 1 1191
2 75456 1 1191
2 75457 1 1192
2 75458 1 1192
2 75459 1 1192
2 75460 1 1192
2 75461 1 1192
2 75462 1 1195
2 75463 1 1195
2 75464 1 1195
2 75465 1 1195
2 75466 1 1195
2 75467 1 1195
2 75468 1 1195
2 75469 1 1195
2 75470 1 1195
2 75471 1 1195
2 75472 1 1195
2 75473 1 1195
2 75474 1 1195
2 75475 1 1195
2 75476 1 1195
2 75477 1 1195
2 75478 1 1195
2 75479 1 1195
2 75480 1 1195
2 75481 1 1195
2 75482 1 1195
2 75483 1 1195
2 75484 1 1195
2 75485 1 1195
2 75486 1 1195
2 75487 1 1195
2 75488 1 1195
2 75489 1 1195
2 75490 1 1195
2 75491 1 1195
2 75492 1 1195
2 75493 1 1195
2 75494 1 1195
2 75495 1 1195
2 75496 1 1195
2 75497 1 1195
2 75498 1 1195
2 75499 1 1195
2 75500 1 1195
2 75501 1 1195
2 75502 1 1195
2 75503 1 1195
2 75504 1 1195
2 75505 1 1195
2 75506 1 1195
2 75507 1 1195
2 75508 1 1195
2 75509 1 1195
2 75510 1 1195
2 75511 1 1195
2 75512 1 1195
2 75513 1 1195
2 75514 1 1195
2 75515 1 1195
2 75516 1 1195
2 75517 1 1195
2 75518 1 1195
2 75519 1 1195
2 75520 1 1195
2 75521 1 1195
2 75522 1 1195
2 75523 1 1195
2 75524 1 1195
2 75525 1 1195
2 75526 1 1195
2 75527 1 1195
2 75528 1 1195
2 75529 1 1195
2 75530 1 1195
2 75531 1 1195
2 75532 1 1195
2 75533 1 1195
2 75534 1 1195
2 75535 1 1195
2 75536 1 1195
2 75537 1 1195
2 75538 1 1196
2 75539 1 1196
2 75540 1 1196
2 75541 1 1196
2 75542 1 1196
2 75543 1 1196
2 75544 1 1196
2 75545 1 1196
2 75546 1 1196
2 75547 1 1196
2 75548 1 1196
2 75549 1 1196
2 75550 1 1196
2 75551 1 1196
2 75552 1 1196
2 75553 1 1196
2 75554 1 1196
2 75555 1 1196
2 75556 1 1196
2 75557 1 1196
2 75558 1 1196
2 75559 1 1196
2 75560 1 1196
2 75561 1 1196
2 75562 1 1196
2 75563 1 1196
2 75564 1 1196
2 75565 1 1196
2 75566 1 1196
2 75567 1 1196
2 75568 1 1196
2 75569 1 1196
2 75570 1 1196
2 75571 1 1196
2 75572 1 1196
2 75573 1 1196
2 75574 1 1196
2 75575 1 1196
2 75576 1 1196
2 75577 1 1196
2 75578 1 1196
2 75579 1 1196
2 75580 1 1196
2 75581 1 1196
2 75582 1 1196
2 75583 1 1196
2 75584 1 1196
2 75585 1 1196
2 75586 1 1196
2 75587 1 1196
2 75588 1 1196
2 75589 1 1196
2 75590 1 1196
2 75591 1 1196
2 75592 1 1196
2 75593 1 1196
2 75594 1 1196
2 75595 1 1196
2 75596 1 1196
2 75597 1 1196
2 75598 1 1196
2 75599 1 1196
2 75600 1 1196
2 75601 1 1196
2 75602 1 1196
2 75603 1 1196
2 75604 1 1196
2 75605 1 1196
2 75606 1 1196
2 75607 1 1196
2 75608 1 1196
2 75609 1 1196
2 75610 1 1196
2 75611 1 1196
2 75612 1 1196
2 75613 1 1196
2 75614 1 1196
2 75615 1 1196
2 75616 1 1196
2 75617 1 1196
2 75618 1 1196
2 75619 1 1196
2 75620 1 1196
2 75621 1 1196
2 75622 1 1196
2 75623 1 1196
2 75624 1 1196
2 75625 1 1196
2 75626 1 1196
2 75627 1 1196
2 75628 1 1196
2 75629 1 1196
2 75630 1 1196
2 75631 1 1196
2 75632 1 1196
2 75633 1 1196
2 75634 1 1196
2 75635 1 1196
2 75636 1 1196
2 75637 1 1196
2 75638 1 1196
2 75639 1 1196
2 75640 1 1196
2 75641 1 1196
2 75642 1 1196
2 75643 1 1196
2 75644 1 1196
2 75645 1 1196
2 75646 1 1196
2 75647 1 1196
2 75648 1 1196
2 75649 1 1196
2 75650 1 1196
2 75651 1 1196
2 75652 1 1196
2 75653 1 1196
2 75654 1 1196
2 75655 1 1196
2 75656 1 1196
2 75657 1 1196
2 75658 1 1196
2 75659 1 1196
2 75660 1 1196
2 75661 1 1196
2 75662 1 1196
2 75663 1 1197
2 75664 1 1197
2 75665 1 1197
2 75666 1 1197
2 75667 1 1197
2 75668 1 1197
2 75669 1 1197
2 75670 1 1197
2 75671 1 1197
2 75672 1 1205
2 75673 1 1205
2 75674 1 1205
2 75675 1 1205
2 75676 1 1205
2 75677 1 1205
2 75678 1 1205
2 75679 1 1205
2 75680 1 1205
2 75681 1 1205
2 75682 1 1205
2 75683 1 1205
2 75684 1 1205
2 75685 1 1205
2 75686 1 1205
2 75687 1 1205
2 75688 1 1205
2 75689 1 1205
2 75690 1 1205
2 75691 1 1205
2 75692 1 1205
2 75693 1 1205
2 75694 1 1205
2 75695 1 1205
2 75696 1 1205
2 75697 1 1206
2 75698 1 1206
2 75699 1 1206
2 75700 1 1206
2 75701 1 1207
2 75702 1 1207
2 75703 1 1207
2 75704 1 1207
2 75705 1 1207
2 75706 1 1207
2 75707 1 1207
2 75708 1 1207
2 75709 1 1207
2 75710 1 1207
2 75711 1 1207
2 75712 1 1207
2 75713 1 1207
2 75714 1 1207
2 75715 1 1207
2 75716 1 1207
2 75717 1 1207
2 75718 1 1207
2 75719 1 1208
2 75720 1 1208
2 75721 1 1208
2 75722 1 1209
2 75723 1 1209
2 75724 1 1209
2 75725 1 1209
2 75726 1 1209
2 75727 1 1210
2 75728 1 1210
2 75729 1 1212
2 75730 1 1212
2 75731 1 1219
2 75732 1 1219
2 75733 1 1219
2 75734 1 1220
2 75735 1 1220
2 75736 1 1220
2 75737 1 1220
2 75738 1 1220
2 75739 1 1220
2 75740 1 1220
2 75741 1 1220
2 75742 1 1220
2 75743 1 1221
2 75744 1 1221
2 75745 1 1221
2 75746 1 1221
2 75747 1 1222
2 75748 1 1222
2 75749 1 1222
2 75750 1 1222
2 75751 1 1222
2 75752 1 1222
2 75753 1 1222
2 75754 1 1222
2 75755 1 1222
2 75756 1 1223
2 75757 1 1223
2 75758 1 1223
2 75759 1 1223
2 75760 1 1223
2 75761 1 1234
2 75762 1 1234
2 75763 1 1235
2 75764 1 1235
2 75765 1 1235
2 75766 1 1235
2 75767 1 1236
2 75768 1 1236
2 75769 1 1236
2 75770 1 1239
2 75771 1 1239
2 75772 1 1239
2 75773 1 1241
2 75774 1 1241
2 75775 1 1241
2 75776 1 1241
2 75777 1 1241
2 75778 1 1241
2 75779 1 1241
2 75780 1 1244
2 75781 1 1244
2 75782 1 1244
2 75783 1 1244
2 75784 1 1244
2 75785 1 1244
2 75786 1 1244
2 75787 1 1244
2 75788 1 1244
2 75789 1 1245
2 75790 1 1245
2 75791 1 1245
2 75792 1 1245
2 75793 1 1255
2 75794 1 1255
2 75795 1 1256
2 75796 1 1256
2 75797 1 1256
2 75798 1 1256
2 75799 1 1256
2 75800 1 1256
2 75801 1 1257
2 75802 1 1257
2 75803 1 1257
2 75804 1 1257
2 75805 1 1257
2 75806 1 1257
2 75807 1 1257
2 75808 1 1258
2 75809 1 1258
2 75810 1 1258
2 75811 1 1259
2 75812 1 1259
2 75813 1 1259
2 75814 1 1260
2 75815 1 1260
2 75816 1 1260
2 75817 1 1260
2 75818 1 1260
2 75819 1 1266
2 75820 1 1266
2 75821 1 1266
2 75822 1 1266
2 75823 1 1266
2 75824 1 1266
2 75825 1 1266
2 75826 1 1266
2 75827 1 1266
2 75828 1 1266
2 75829 1 1266
2 75830 1 1266
2 75831 1 1266
2 75832 1 1266
2 75833 1 1266
2 75834 1 1266
2 75835 1 1266
2 75836 1 1266
2 75837 1 1266
2 75838 1 1266
2 75839 1 1266
2 75840 1 1266
2 75841 1 1266
2 75842 1 1266
2 75843 1 1266
2 75844 1 1266
2 75845 1 1266
2 75846 1 1266
2 75847 1 1266
2 75848 1 1266
2 75849 1 1266
2 75850 1 1266
2 75851 1 1266
2 75852 1 1266
2 75853 1 1266
2 75854 1 1266
2 75855 1 1266
2 75856 1 1266
2 75857 1 1267
2 75858 1 1267
2 75859 1 1268
2 75860 1 1268
2 75861 1 1268
2 75862 1 1269
2 75863 1 1269
2 75864 1 1269
2 75865 1 1269
2 75866 1 1273
2 75867 1 1273
2 75868 1 1274
2 75869 1 1274
2 75870 1 1274
2 75871 1 1274
2 75872 1 1274
2 75873 1 1274
2 75874 1 1274
2 75875 1 1274
2 75876 1 1274
2 75877 1 1274
2 75878 1 1274
2 75879 1 1274
2 75880 1 1274
2 75881 1 1274
2 75882 1 1274
2 75883 1 1274
2 75884 1 1274
2 75885 1 1275
2 75886 1 1275
2 75887 1 1275
2 75888 1 1275
2 75889 1 1275
2 75890 1 1290
2 75891 1 1290
2 75892 1 1291
2 75893 1 1291
2 75894 1 1296
2 75895 1 1296
2 75896 1 1296
2 75897 1 1296
2 75898 1 1296
2 75899 1 1296
2 75900 1 1296
2 75901 1 1296
2 75902 1 1296
2 75903 1 1296
2 75904 1 1296
2 75905 1 1296
2 75906 1 1296
2 75907 1 1296
2 75908 1 1296
2 75909 1 1296
2 75910 1 1296
2 75911 1 1296
2 75912 1 1297
2 75913 1 1297
2 75914 1 1298
2 75915 1 1298
2 75916 1 1298
2 75917 1 1298
2 75918 1 1298
2 75919 1 1298
2 75920 1 1298
2 75921 1 1298
2 75922 1 1298
2 75923 1 1298
2 75924 1 1298
2 75925 1 1298
2 75926 1 1299
2 75927 1 1299
2 75928 1 1299
2 75929 1 1299
2 75930 1 1299
2 75931 1 1299
2 75932 1 1301
2 75933 1 1301
2 75934 1 1301
2 75935 1 1306
2 75936 1 1306
2 75937 1 1306
2 75938 1 1306
2 75939 1 1306
2 75940 1 1306
2 75941 1 1306
2 75942 1 1306
2 75943 1 1306
2 75944 1 1307
2 75945 1 1307
2 75946 1 1317
2 75947 1 1317
2 75948 1 1317
2 75949 1 1318
2 75950 1 1318
2 75951 1 1319
2 75952 1 1319
2 75953 1 1319
2 75954 1 1319
2 75955 1 1319
2 75956 1 1319
2 75957 1 1320
2 75958 1 1320
2 75959 1 1320
2 75960 1 1320
2 75961 1 1320
2 75962 1 1320
2 75963 1 1320
2 75964 1 1320
2 75965 1 1320
2 75966 1 1320
2 75967 1 1320
2 75968 1 1320
2 75969 1 1320
2 75970 1 1320
2 75971 1 1322
2 75972 1 1322
2 75973 1 1322
2 75974 1 1322
2 75975 1 1332
2 75976 1 1332
2 75977 1 1336
2 75978 1 1336
2 75979 1 1336
2 75980 1 1336
2 75981 1 1336
2 75982 1 1337
2 75983 1 1337
2 75984 1 1337
2 75985 1 1338
2 75986 1 1338
2 75987 1 1338
2 75988 1 1340
2 75989 1 1340
2 75990 1 1343
2 75991 1 1343
2 75992 1 1350
2 75993 1 1350
2 75994 1 1350
2 75995 1 1350
2 75996 1 1350
2 75997 1 1350
2 75998 1 1350
2 75999 1 1350
2 76000 1 1350
2 76001 1 1351
2 76002 1 1351
2 76003 1 1351
2 76004 1 1351
2 76005 1 1351
2 76006 1 1351
2 76007 1 1351
2 76008 1 1351
2 76009 1 1351
2 76010 1 1351
2 76011 1 1351
2 76012 1 1351
2 76013 1 1351
2 76014 1 1364
2 76015 1 1364
2 76016 1 1364
2 76017 1 1364
2 76018 1 1364
2 76019 1 1365
2 76020 1 1365
2 76021 1 1365
2 76022 1 1365
2 76023 1 1372
2 76024 1 1372
2 76025 1 1372
2 76026 1 1373
2 76027 1 1373
2 76028 1 1373
2 76029 1 1376
2 76030 1 1376
2 76031 1 1376
2 76032 1 1377
2 76033 1 1377
2 76034 1 1377
2 76035 1 1383
2 76036 1 1383
2 76037 1 1386
2 76038 1 1386
2 76039 1 1386
2 76040 1 1386
2 76041 1 1387
2 76042 1 1387
2 76043 1 1387
2 76044 1 1387
2 76045 1 1387
2 76046 1 1387
2 76047 1 1387
2 76048 1 1387
2 76049 1 1387
2 76050 1 1387
2 76051 1 1387
2 76052 1 1387
2 76053 1 1387
2 76054 1 1387
2 76055 1 1387
2 76056 1 1387
2 76057 1 1387
2 76058 1 1387
2 76059 1 1387
2 76060 1 1387
2 76061 1 1387
2 76062 1 1387
2 76063 1 1387
2 76064 1 1388
2 76065 1 1388
2 76066 1 1389
2 76067 1 1389
2 76068 1 1389
2 76069 1 1389
2 76070 1 1389
2 76071 1 1389
2 76072 1 1389
2 76073 1 1389
2 76074 1 1389
2 76075 1 1390
2 76076 1 1390
2 76077 1 1390
2 76078 1 1390
2 76079 1 1390
2 76080 1 1390
2 76081 1 1390
2 76082 1 1390
2 76083 1 1390
2 76084 1 1391
2 76085 1 1391
2 76086 1 1391
2 76087 1 1398
2 76088 1 1398
2 76089 1 1398
2 76090 1 1398
2 76091 1 1398
2 76092 1 1398
2 76093 1 1398
2 76094 1 1398
2 76095 1 1399
2 76096 1 1399
2 76097 1 1399
2 76098 1 1399
2 76099 1 1399
2 76100 1 1399
2 76101 1 1400
2 76102 1 1400
2 76103 1 1404
2 76104 1 1404
2 76105 1 1404
2 76106 1 1404
2 76107 1 1404
2 76108 1 1404
2 76109 1 1405
2 76110 1 1405
2 76111 1 1405
2 76112 1 1405
2 76113 1 1405
2 76114 1 1407
2 76115 1 1407
2 76116 1 1407
2 76117 1 1407
2 76118 1 1407
2 76119 1 1407
2 76120 1 1407
2 76121 1 1407
2 76122 1 1419
2 76123 1 1419
2 76124 1 1419
2 76125 1 1419
2 76126 1 1419
2 76127 1 1419
2 76128 1 1419
2 76129 1 1419
2 76130 1 1420
2 76131 1 1420
2 76132 1 1420
2 76133 1 1422
2 76134 1 1422
2 76135 1 1427
2 76136 1 1427
2 76137 1 1428
2 76138 1 1428
2 76139 1 1428
2 76140 1 1428
2 76141 1 1428
2 76142 1 1428
2 76143 1 1428
2 76144 1 1428
2 76145 1 1428
2 76146 1 1428
2 76147 1 1428
2 76148 1 1428
2 76149 1 1428
2 76150 1 1428
2 76151 1 1428
2 76152 1 1428
2 76153 1 1429
2 76154 1 1429
2 76155 1 1429
2 76156 1 1435
2 76157 1 1435
2 76158 1 1435
2 76159 1 1435
2 76160 1 1435
2 76161 1 1435
2 76162 1 1435
2 76163 1 1435
2 76164 1 1435
2 76165 1 1435
2 76166 1 1435
2 76167 1 1435
2 76168 1 1435
2 76169 1 1435
2 76170 1 1435
2 76171 1 1435
2 76172 1 1435
2 76173 1 1435
2 76174 1 1435
2 76175 1 1435
2 76176 1 1435
2 76177 1 1435
2 76178 1 1435
2 76179 1 1435
2 76180 1 1435
2 76181 1 1435
2 76182 1 1435
2 76183 1 1435
2 76184 1 1435
2 76185 1 1435
2 76186 1 1435
2 76187 1 1435
2 76188 1 1435
2 76189 1 1435
2 76190 1 1435
2 76191 1 1435
2 76192 1 1435
2 76193 1 1435
2 76194 1 1436
2 76195 1 1436
2 76196 1 1436
2 76197 1 1436
2 76198 1 1436
2 76199 1 1436
2 76200 1 1436
2 76201 1 1436
2 76202 1 1436
2 76203 1 1436
2 76204 1 1436
2 76205 1 1436
2 76206 1 1436
2 76207 1 1436
2 76208 1 1436
2 76209 1 1436
2 76210 1 1436
2 76211 1 1436
2 76212 1 1436
2 76213 1 1436
2 76214 1 1436
2 76215 1 1436
2 76216 1 1436
2 76217 1 1437
2 76218 1 1437
2 76219 1 1437
2 76220 1 1437
2 76221 1 1438
2 76222 1 1438
2 76223 1 1438
2 76224 1 1438
2 76225 1 1439
2 76226 1 1439
2 76227 1 1440
2 76228 1 1440
2 76229 1 1443
2 76230 1 1443
2 76231 1 1443
2 76232 1 1443
2 76233 1 1443
2 76234 1 1443
2 76235 1 1444
2 76236 1 1444
2 76237 1 1455
2 76238 1 1455
2 76239 1 1455
2 76240 1 1455
2 76241 1 1455
2 76242 1 1455
2 76243 1 1456
2 76244 1 1456
2 76245 1 1456
2 76246 1 1456
2 76247 1 1456
2 76248 1 1456
2 76249 1 1456
2 76250 1 1456
2 76251 1 1456
2 76252 1 1456
2 76253 1 1456
2 76254 1 1456
2 76255 1 1456
2 76256 1 1456
2 76257 1 1456
2 76258 1 1456
2 76259 1 1456
2 76260 1 1456
2 76261 1 1456
2 76262 1 1456
2 76263 1 1456
2 76264 1 1456
2 76265 1 1456
2 76266 1 1456
2 76267 1 1456
2 76268 1 1456
2 76269 1 1456
2 76270 1 1456
2 76271 1 1456
2 76272 1 1456
2 76273 1 1456
2 76274 1 1456
2 76275 1 1456
2 76276 1 1456
2 76277 1 1456
2 76278 1 1456
2 76279 1 1456
2 76280 1 1456
2 76281 1 1456
2 76282 1 1456
2 76283 1 1456
2 76284 1 1456
2 76285 1 1456
2 76286 1 1456
2 76287 1 1456
2 76288 1 1456
2 76289 1 1456
2 76290 1 1456
2 76291 1 1456
2 76292 1 1456
2 76293 1 1456
2 76294 1 1456
2 76295 1 1456
2 76296 1 1456
2 76297 1 1456
2 76298 1 1456
2 76299 1 1456
2 76300 1 1456
2 76301 1 1456
2 76302 1 1456
2 76303 1 1456
2 76304 1 1456
2 76305 1 1457
2 76306 1 1457
2 76307 1 1458
2 76308 1 1458
2 76309 1 1458
2 76310 1 1460
2 76311 1 1460
2 76312 1 1460
2 76313 1 1463
2 76314 1 1463
2 76315 1 1463
2 76316 1 1463
2 76317 1 1463
2 76318 1 1463
2 76319 1 1463
2 76320 1 1463
2 76321 1 1464
2 76322 1 1464
2 76323 1 1464
2 76324 1 1464
2 76325 1 1464
2 76326 1 1464
2 76327 1 1464
2 76328 1 1464
2 76329 1 1464
2 76330 1 1464
2 76331 1 1471
2 76332 1 1471
2 76333 1 1471
2 76334 1 1471
2 76335 1 1471
2 76336 1 1471
2 76337 1 1471
2 76338 1 1471
2 76339 1 1471
2 76340 1 1471
2 76341 1 1471
2 76342 1 1471
2 76343 1 1471
2 76344 1 1471
2 76345 1 1471
2 76346 1 1471
2 76347 1 1471
2 76348 1 1471
2 76349 1 1471
2 76350 1 1471
2 76351 1 1471
2 76352 1 1471
2 76353 1 1472
2 76354 1 1472
2 76355 1 1472
2 76356 1 1472
2 76357 1 1472
2 76358 1 1472
2 76359 1 1472
2 76360 1 1472
2 76361 1 1472
2 76362 1 1472
2 76363 1 1472
2 76364 1 1472
2 76365 1 1472
2 76366 1 1472
2 76367 1 1472
2 76368 1 1472
2 76369 1 1472
2 76370 1 1472
2 76371 1 1472
2 76372 1 1472
2 76373 1 1472
2 76374 1 1472
2 76375 1 1472
2 76376 1 1473
2 76377 1 1473
2 76378 1 1480
2 76379 1 1480
2 76380 1 1481
2 76381 1 1481
2 76382 1 1481
2 76383 1 1481
2 76384 1 1481
2 76385 1 1481
2 76386 1 1481
2 76387 1 1481
2 76388 1 1481
2 76389 1 1491
2 76390 1 1491
2 76391 1 1494
2 76392 1 1494
2 76393 1 1495
2 76394 1 1495
2 76395 1 1499
2 76396 1 1499
2 76397 1 1513
2 76398 1 1513
2 76399 1 1514
2 76400 1 1514
2 76401 1 1514
2 76402 1 1514
2 76403 1 1514
2 76404 1 1514
2 76405 1 1514
2 76406 1 1514
2 76407 1 1514
2 76408 1 1514
2 76409 1 1514
2 76410 1 1514
2 76411 1 1514
2 76412 1 1514
2 76413 1 1514
2 76414 1 1514
2 76415 1 1514
2 76416 1 1514
2 76417 1 1514
2 76418 1 1514
2 76419 1 1514
2 76420 1 1515
2 76421 1 1515
2 76422 1 1515
2 76423 1 1515
2 76424 1 1515
2 76425 1 1515
2 76426 1 1515
2 76427 1 1515
2 76428 1 1515
2 76429 1 1515
2 76430 1 1515
2 76431 1 1515
2 76432 1 1516
2 76433 1 1516
2 76434 1 1516
2 76435 1 1516
2 76436 1 1516
2 76437 1 1517
2 76438 1 1517
2 76439 1 1517
2 76440 1 1517
2 76441 1 1517
2 76442 1 1517
2 76443 1 1517
2 76444 1 1517
2 76445 1 1517
2 76446 1 1517
2 76447 1 1517
2 76448 1 1517
2 76449 1 1517
2 76450 1 1517
2 76451 1 1517
2 76452 1 1517
2 76453 1 1517
2 76454 1 1517
2 76455 1 1518
2 76456 1 1518
2 76457 1 1518
2 76458 1 1530
2 76459 1 1530
2 76460 1 1531
2 76461 1 1531
2 76462 1 1541
2 76463 1 1541
2 76464 1 1546
2 76465 1 1546
2 76466 1 1552
2 76467 1 1552
2 76468 1 1553
2 76469 1 1553
2 76470 1 1559
2 76471 1 1559
2 76472 1 1561
2 76473 1 1561
2 76474 1 1561
2 76475 1 1563
2 76476 1 1563
2 76477 1 1564
2 76478 1 1564
2 76479 1 1564
2 76480 1 1564
2 76481 1 1564
2 76482 1 1564
2 76483 1 1567
2 76484 1 1567
2 76485 1 1568
2 76486 1 1568
2 76487 1 1568
2 76488 1 1568
2 76489 1 1568
2 76490 1 1568
2 76491 1 1568
2 76492 1 1568
2 76493 1 1568
2 76494 1 1568
2 76495 1 1568
2 76496 1 1568
2 76497 1 1568
2 76498 1 1568
2 76499 1 1568
2 76500 1 1568
2 76501 1 1568
2 76502 1 1568
2 76503 1 1568
2 76504 1 1568
2 76505 1 1568
2 76506 1 1569
2 76507 1 1569
2 76508 1 1569
2 76509 1 1569
2 76510 1 1569
2 76511 1 1569
2 76512 1 1569
2 76513 1 1570
2 76514 1 1570
2 76515 1 1571
2 76516 1 1571
2 76517 1 1571
2 76518 1 1587
2 76519 1 1587
2 76520 1 1595
2 76521 1 1595
2 76522 1 1595
2 76523 1 1595
2 76524 1 1596
2 76525 1 1596
2 76526 1 1596
2 76527 1 1597
2 76528 1 1597
2 76529 1 1597
2 76530 1 1598
2 76531 1 1598
2 76532 1 1600
2 76533 1 1600
2 76534 1 1603
2 76535 1 1603
2 76536 1 1604
2 76537 1 1604
2 76538 1 1604
2 76539 1 1604
2 76540 1 1604
2 76541 1 1604
2 76542 1 1605
2 76543 1 1605
2 76544 1 1608
2 76545 1 1608
2 76546 1 1609
2 76547 1 1609
2 76548 1 1609
2 76549 1 1609
2 76550 1 1609
2 76551 1 1609
2 76552 1 1609
2 76553 1 1609
2 76554 1 1609
2 76555 1 1609
2 76556 1 1609
2 76557 1 1609
2 76558 1 1609
2 76559 1 1609
2 76560 1 1609
2 76561 1 1609
2 76562 1 1609
2 76563 1 1609
2 76564 1 1609
2 76565 1 1609
2 76566 1 1609
2 76567 1 1609
2 76568 1 1609
2 76569 1 1609
2 76570 1 1610
2 76571 1 1610
2 76572 1 1610
2 76573 1 1610
2 76574 1 1610
2 76575 1 1610
2 76576 1 1611
2 76577 1 1611
2 76578 1 1611
2 76579 1 1611
2 76580 1 1611
2 76581 1 1611
2 76582 1 1612
2 76583 1 1612
2 76584 1 1617
2 76585 1 1617
2 76586 1 1617
2 76587 1 1617
2 76588 1 1617
2 76589 1 1617
2 76590 1 1617
2 76591 1 1617
2 76592 1 1619
2 76593 1 1619
2 76594 1 1619
2 76595 1 1619
2 76596 1 1620
2 76597 1 1620
2 76598 1 1620
2 76599 1 1620
2 76600 1 1636
2 76601 1 1636
2 76602 1 1643
2 76603 1 1643
2 76604 1 1644
2 76605 1 1644
2 76606 1 1646
2 76607 1 1646
2 76608 1 1651
2 76609 1 1651
2 76610 1 1651
2 76611 1 1651
2 76612 1 1651
2 76613 1 1651
2 76614 1 1651
2 76615 1 1651
2 76616 1 1651
2 76617 1 1651
2 76618 1 1651
2 76619 1 1651
2 76620 1 1651
2 76621 1 1651
2 76622 1 1651
2 76623 1 1651
2 76624 1 1651
2 76625 1 1651
2 76626 1 1651
2 76627 1 1651
2 76628 1 1651
2 76629 1 1651
2 76630 1 1651
2 76631 1 1651
2 76632 1 1651
2 76633 1 1651
2 76634 1 1651
2 76635 1 1651
2 76636 1 1651
2 76637 1 1651
2 76638 1 1651
2 76639 1 1651
2 76640 1 1651
2 76641 1 1651
2 76642 1 1651
2 76643 1 1651
2 76644 1 1651
2 76645 1 1651
2 76646 1 1651
2 76647 1 1651
2 76648 1 1651
2 76649 1 1651
2 76650 1 1651
2 76651 1 1651
2 76652 1 1651
2 76653 1 1651
2 76654 1 1651
2 76655 1 1651
2 76656 1 1652
2 76657 1 1652
2 76658 1 1652
2 76659 1 1652
2 76660 1 1652
2 76661 1 1652
2 76662 1 1652
2 76663 1 1652
2 76664 1 1652
2 76665 1 1652
2 76666 1 1652
2 76667 1 1652
2 76668 1 1652
2 76669 1 1652
2 76670 1 1652
2 76671 1 1652
2 76672 1 1652
2 76673 1 1652
2 76674 1 1652
2 76675 1 1652
2 76676 1 1652
2 76677 1 1652
2 76678 1 1652
2 76679 1 1652
2 76680 1 1653
2 76681 1 1653
2 76682 1 1653
2 76683 1 1653
2 76684 1 1657
2 76685 1 1657
2 76686 1 1665
2 76687 1 1665
2 76688 1 1666
2 76689 1 1666
2 76690 1 1667
2 76691 1 1667
2 76692 1 1667
2 76693 1 1667
2 76694 1 1667
2 76695 1 1667
2 76696 1 1667
2 76697 1 1667
2 76698 1 1667
2 76699 1 1667
2 76700 1 1667
2 76701 1 1667
2 76702 1 1667
2 76703 1 1667
2 76704 1 1667
2 76705 1 1667
2 76706 1 1667
2 76707 1 1667
2 76708 1 1668
2 76709 1 1668
2 76710 1 1669
2 76711 1 1669
2 76712 1 1677
2 76713 1 1677
2 76714 1 1677
2 76715 1 1677
2 76716 1 1677
2 76717 1 1677
2 76718 1 1677
2 76719 1 1677
2 76720 1 1677
2 76721 1 1678
2 76722 1 1678
2 76723 1 1679
2 76724 1 1679
2 76725 1 1679
2 76726 1 1679
2 76727 1 1680
2 76728 1 1680
2 76729 1 1680
2 76730 1 1680
2 76731 1 1680
2 76732 1 1680
2 76733 1 1680
2 76734 1 1681
2 76735 1 1681
2 76736 1 1685
2 76737 1 1685
2 76738 1 1685
2 76739 1 1685
2 76740 1 1685
2 76741 1 1685
2 76742 1 1685
2 76743 1 1685
2 76744 1 1685
2 76745 1 1685
2 76746 1 1685
2 76747 1 1685
2 76748 1 1685
2 76749 1 1685
2 76750 1 1685
2 76751 1 1685
2 76752 1 1685
2 76753 1 1685
2 76754 1 1685
2 76755 1 1686
2 76756 1 1686
2 76757 1 1686
2 76758 1 1686
2 76759 1 1686
2 76760 1 1686
2 76761 1 1686
2 76762 1 1686
2 76763 1 1686
2 76764 1 1686
2 76765 1 1686
2 76766 1 1686
2 76767 1 1686
2 76768 1 1686
2 76769 1 1686
2 76770 1 1686
2 76771 1 1686
2 76772 1 1686
2 76773 1 1686
2 76774 1 1686
2 76775 1 1686
2 76776 1 1686
2 76777 1 1686
2 76778 1 1686
2 76779 1 1686
2 76780 1 1686
2 76781 1 1686
2 76782 1 1686
2 76783 1 1686
2 76784 1 1686
2 76785 1 1686
2 76786 1 1686
2 76787 1 1686
2 76788 1 1686
2 76789 1 1686
2 76790 1 1686
2 76791 1 1686
2 76792 1 1686
2 76793 1 1686
2 76794 1 1686
2 76795 1 1686
2 76796 1 1686
2 76797 1 1686
2 76798 1 1686
2 76799 1 1686
2 76800 1 1686
2 76801 1 1686
2 76802 1 1686
2 76803 1 1686
2 76804 1 1686
2 76805 1 1686
2 76806 1 1686
2 76807 1 1686
2 76808 1 1686
2 76809 1 1686
2 76810 1 1686
2 76811 1 1686
2 76812 1 1686
2 76813 1 1695
2 76814 1 1695
2 76815 1 1695
2 76816 1 1695
2 76817 1 1695
2 76818 1 1695
2 76819 1 1695
2 76820 1 1695
2 76821 1 1695
2 76822 1 1695
2 76823 1 1695
2 76824 1 1695
2 76825 1 1695
2 76826 1 1695
2 76827 1 1695
2 76828 1 1695
2 76829 1 1695
2 76830 1 1695
2 76831 1 1695
2 76832 1 1696
2 76833 1 1696
2 76834 1 1696
2 76835 1 1696
2 76836 1 1696
2 76837 1 1696
2 76838 1 1696
2 76839 1 1696
2 76840 1 1696
2 76841 1 1696
2 76842 1 1696
2 76843 1 1696
2 76844 1 1696
2 76845 1 1696
2 76846 1 1696
2 76847 1 1696
2 76848 1 1696
2 76849 1 1696
2 76850 1 1696
2 76851 1 1696
2 76852 1 1696
2 76853 1 1696
2 76854 1 1697
2 76855 1 1697
2 76856 1 1697
2 76857 1 1698
2 76858 1 1698
2 76859 1 1698
2 76860 1 1698
2 76861 1 1699
2 76862 1 1699
2 76863 1 1700
2 76864 1 1700
2 76865 1 1700
2 76866 1 1700
2 76867 1 1700
2 76868 1 1700
2 76869 1 1700
2 76870 1 1700
2 76871 1 1700
2 76872 1 1700
2 76873 1 1700
2 76874 1 1701
2 76875 1 1701
2 76876 1 1701
2 76877 1 1701
2 76878 1 1701
2 76879 1 1701
2 76880 1 1702
2 76881 1 1702
2 76882 1 1702
2 76883 1 1702
2 76884 1 1702
2 76885 1 1702
2 76886 1 1702
2 76887 1 1702
2 76888 1 1703
2 76889 1 1703
2 76890 1 1705
2 76891 1 1705
2 76892 1 1710
2 76893 1 1710
2 76894 1 1724
2 76895 1 1724
2 76896 1 1724
2 76897 1 1725
2 76898 1 1725
2 76899 1 1725
2 76900 1 1725
2 76901 1 1725
2 76902 1 1725
2 76903 1 1725
2 76904 1 1726
2 76905 1 1726
2 76906 1 1726
2 76907 1 1726
2 76908 1 1726
2 76909 1 1726
2 76910 1 1726
2 76911 1 1726
2 76912 1 1726
2 76913 1 1727
2 76914 1 1727
2 76915 1 1728
2 76916 1 1728
2 76917 1 1728
2 76918 1 1728
2 76919 1 1728
2 76920 1 1728
2 76921 1 1728
2 76922 1 1729
2 76923 1 1729
2 76924 1 1729
2 76925 1 1729
2 76926 1 1729
2 76927 1 1729
2 76928 1 1729
2 76929 1 1729
2 76930 1 1729
2 76931 1 1729
2 76932 1 1729
2 76933 1 1729
2 76934 1 1729
2 76935 1 1729
2 76936 1 1729
2 76937 1 1730
2 76938 1 1730
2 76939 1 1735
2 76940 1 1735
2 76941 1 1742
2 76942 1 1742
2 76943 1 1742
2 76944 1 1742
2 76945 1 1742
2 76946 1 1743
2 76947 1 1743
2 76948 1 1746
2 76949 1 1746
2 76950 1 1750
2 76951 1 1750
2 76952 1 1755
2 76953 1 1755
2 76954 1 1755
2 76955 1 1755
2 76956 1 1755
2 76957 1 1755
2 76958 1 1755
2 76959 1 1755
2 76960 1 1755
2 76961 1 1755
2 76962 1 1755
2 76963 1 1756
2 76964 1 1756
2 76965 1 1757
2 76966 1 1757
2 76967 1 1757
2 76968 1 1763
2 76969 1 1763
2 76970 1 1763
2 76971 1 1763
2 76972 1 1763
2 76973 1 1767
2 76974 1 1767
2 76975 1 1767
2 76976 1 1768
2 76977 1 1768
2 76978 1 1768
2 76979 1 1768
2 76980 1 1768
2 76981 1 1768
2 76982 1 1779
2 76983 1 1779
2 76984 1 1779
2 76985 1 1779
2 76986 1 1779
2 76987 1 1780
2 76988 1 1780
2 76989 1 1780
2 76990 1 1780
2 76991 1 1780
2 76992 1 1780
2 76993 1 1780
2 76994 1 1780
2 76995 1 1780
2 76996 1 1780
2 76997 1 1780
2 76998 1 1780
2 76999 1 1780
2 77000 1 1780
2 77001 1 1780
2 77002 1 1780
2 77003 1 1780
2 77004 1 1780
2 77005 1 1780
2 77006 1 1780
2 77007 1 1780
2 77008 1 1780
2 77009 1 1780
2 77010 1 1780
2 77011 1 1780
2 77012 1 1780
2 77013 1 1780
2 77014 1 1780
2 77015 1 1780
2 77016 1 1781
2 77017 1 1781
2 77018 1 1781
2 77019 1 1781
2 77020 1 1781
2 77021 1 1781
2 77022 1 1781
2 77023 1 1781
2 77024 1 1782
2 77025 1 1782
2 77026 1 1782
2 77027 1 1782
2 77028 1 1783
2 77029 1 1783
2 77030 1 1783
2 77031 1 1783
2 77032 1 1783
2 77033 1 1783
2 77034 1 1783
2 77035 1 1783
2 77036 1 1783
2 77037 1 1783
2 77038 1 1783
2 77039 1 1783
2 77040 1 1783
2 77041 1 1783
2 77042 1 1783
2 77043 1 1783
2 77044 1 1783
2 77045 1 1783
2 77046 1 1784
2 77047 1 1784
2 77048 1 1784
2 77049 1 1784
2 77050 1 1784
2 77051 1 1784
2 77052 1 1784
2 77053 1 1784
2 77054 1 1784
2 77055 1 1784
2 77056 1 1785
2 77057 1 1785
2 77058 1 1797
2 77059 1 1797
2 77060 1 1797
2 77061 1 1797
2 77062 1 1797
2 77063 1 1797
2 77064 1 1797
2 77065 1 1797
2 77066 1 1797
2 77067 1 1797
2 77068 1 1797
2 77069 1 1797
2 77070 1 1797
2 77071 1 1797
2 77072 1 1797
2 77073 1 1797
2 77074 1 1797
2 77075 1 1797
2 77076 1 1797
2 77077 1 1797
2 77078 1 1797
2 77079 1 1797
2 77080 1 1797
2 77081 1 1797
2 77082 1 1799
2 77083 1 1799
2 77084 1 1800
2 77085 1 1800
2 77086 1 1801
2 77087 1 1801
2 77088 1 1801
2 77089 1 1801
2 77090 1 1801
2 77091 1 1801
2 77092 1 1801
2 77093 1 1801
2 77094 1 1801
2 77095 1 1801
2 77096 1 1801
2 77097 1 1801
2 77098 1 1801
2 77099 1 1801
2 77100 1 1801
2 77101 1 1801
2 77102 1 1802
2 77103 1 1802
2 77104 1 1802
2 77105 1 1802
2 77106 1 1804
2 77107 1 1804
2 77108 1 1805
2 77109 1 1805
2 77110 1 1810
2 77111 1 1810
2 77112 1 1810
2 77113 1 1810
2 77114 1 1810
2 77115 1 1810
2 77116 1 1810
2 77117 1 1810
2 77118 1 1810
2 77119 1 1810
2 77120 1 1810
2 77121 1 1811
2 77122 1 1811
2 77123 1 1811
2 77124 1 1811
2 77125 1 1811
2 77126 1 1811
2 77127 1 1812
2 77128 1 1812
2 77129 1 1815
2 77130 1 1815
2 77131 1 1821
2 77132 1 1821
2 77133 1 1821
2 77134 1 1821
2 77135 1 1821
2 77136 1 1821
2 77137 1 1826
2 77138 1 1826
2 77139 1 1828
2 77140 1 1828
2 77141 1 1842
2 77142 1 1842
2 77143 1 1842
2 77144 1 1842
2 77145 1 1842
2 77146 1 1842
2 77147 1 1842
2 77148 1 1844
2 77149 1 1844
2 77150 1 1844
2 77151 1 1845
2 77152 1 1845
2 77153 1 1846
2 77154 1 1846
2 77155 1 1846
2 77156 1 1846
2 77157 1 1846
2 77158 1 1846
2 77159 1 1846
2 77160 1 1846
2 77161 1 1846
2 77162 1 1846
2 77163 1 1846
2 77164 1 1846
2 77165 1 1846
2 77166 1 1847
2 77167 1 1847
2 77168 1 1847
2 77169 1 1847
2 77170 1 1847
2 77171 1 1847
2 77172 1 1847
2 77173 1 1847
2 77174 1 1848
2 77175 1 1848
2 77176 1 1848
2 77177 1 1849
2 77178 1 1849
2 77179 1 1849
2 77180 1 1849
2 77181 1 1849
2 77182 1 1849
2 77183 1 1849
2 77184 1 1849
2 77185 1 1849
2 77186 1 1849
2 77187 1 1849
2 77188 1 1849
2 77189 1 1849
2 77190 1 1849
2 77191 1 1849
2 77192 1 1849
2 77193 1 1849
2 77194 1 1849
2 77195 1 1849
2 77196 1 1849
2 77197 1 1849
2 77198 1 1850
2 77199 1 1850
2 77200 1 1850
2 77201 1 1850
2 77202 1 1851
2 77203 1 1851
2 77204 1 1851
2 77205 1 1862
2 77206 1 1862
2 77207 1 1864
2 77208 1 1864
2 77209 1 1864
2 77210 1 1864
2 77211 1 1865
2 77212 1 1865
2 77213 1 1865
2 77214 1 1865
2 77215 1 1865
2 77216 1 1865
2 77217 1 1865
2 77218 1 1865
2 77219 1 1865
2 77220 1 1865
2 77221 1 1866
2 77222 1 1866
2 77223 1 1866
2 77224 1 1876
2 77225 1 1876
2 77226 1 1876
2 77227 1 1876
2 77228 1 1876
2 77229 1 1876
2 77230 1 1876
2 77231 1 1876
2 77232 1 1876
2 77233 1 1876
2 77234 1 1876
2 77235 1 1876
2 77236 1 1876
2 77237 1 1876
2 77238 1 1876
2 77239 1 1876
2 77240 1 1876
2 77241 1 1877
2 77242 1 1877
2 77243 1 1877
2 77244 1 1877
2 77245 1 1877
2 77246 1 1878
2 77247 1 1878
2 77248 1 1878
2 77249 1 1878
2 77250 1 1878
2 77251 1 1878
2 77252 1 1879
2 77253 1 1879
2 77254 1 1880
2 77255 1 1880
2 77256 1 1880
2 77257 1 1880
2 77258 1 1880
2 77259 1 1880
2 77260 1 1881
2 77261 1 1881
2 77262 1 1881
2 77263 1 1881
2 77264 1 1882
2 77265 1 1882
2 77266 1 1883
2 77267 1 1883
2 77268 1 1886
2 77269 1 1886
2 77270 1 1889
2 77271 1 1889
2 77272 1 1890
2 77273 1 1890
2 77274 1 1891
2 77275 1 1891
2 77276 1 1891
2 77277 1 1892
2 77278 1 1892
2 77279 1 1896
2 77280 1 1896
2 77281 1 1896
2 77282 1 1909
2 77283 1 1909
2 77284 1 1909
2 77285 1 1909
2 77286 1 1909
2 77287 1 1909
2 77288 1 1909
2 77289 1 1909
2 77290 1 1909
2 77291 1 1909
2 77292 1 1909
2 77293 1 1909
2 77294 1 1909
2 77295 1 1909
2 77296 1 1909
2 77297 1 1909
2 77298 1 1909
2 77299 1 1909
2 77300 1 1909
2 77301 1 1909
2 77302 1 1909
2 77303 1 1910
2 77304 1 1910
2 77305 1 1910
2 77306 1 1910
2 77307 1 1910
2 77308 1 1910
2 77309 1 1910
2 77310 1 1910
2 77311 1 1910
2 77312 1 1919
2 77313 1 1919
2 77314 1 1919
2 77315 1 1919
2 77316 1 1919
2 77317 1 1919
2 77318 1 1919
2 77319 1 1919
2 77320 1 1919
2 77321 1 1919
2 77322 1 1920
2 77323 1 1920
2 77324 1 1920
2 77325 1 1920
2 77326 1 1920
2 77327 1 1920
2 77328 1 1920
2 77329 1 1921
2 77330 1 1921
2 77331 1 1921
2 77332 1 1921
2 77333 1 1922
2 77334 1 1922
2 77335 1 1923
2 77336 1 1923
2 77337 1 1923
2 77338 1 1923
2 77339 1 1923
2 77340 1 1923
2 77341 1 1923
2 77342 1 1924
2 77343 1 1924
2 77344 1 1926
2 77345 1 1926
2 77346 1 1926
2 77347 1 1926
2 77348 1 1926
2 77349 1 1926
2 77350 1 1926
2 77351 1 1926
2 77352 1 1926
2 77353 1 1926
2 77354 1 1926
2 77355 1 1926
2 77356 1 1927
2 77357 1 1927
2 77358 1 1927
2 77359 1 1927
2 77360 1 1934
2 77361 1 1934
2 77362 1 1934
2 77363 1 1935
2 77364 1 1935
2 77365 1 1936
2 77366 1 1936
2 77367 1 1936
2 77368 1 1936
2 77369 1 1936
2 77370 1 1936
2 77371 1 1936
2 77372 1 1936
2 77373 1 1936
2 77374 1 1936
2 77375 1 1936
2 77376 1 1936
2 77377 1 1936
2 77378 1 1936
2 77379 1 1936
2 77380 1 1937
2 77381 1 1937
2 77382 1 1937
2 77383 1 1937
2 77384 1 1937
2 77385 1 1937
2 77386 1 1937
2 77387 1 1937
2 77388 1 1938
2 77389 1 1938
2 77390 1 1938
2 77391 1 1938
2 77392 1 1938
2 77393 1 1938
2 77394 1 1938
2 77395 1 1938
2 77396 1 1938
2 77397 1 1938
2 77398 1 1938
2 77399 1 1938
2 77400 1 1938
2 77401 1 1938
2 77402 1 1938
2 77403 1 1938
2 77404 1 1938
2 77405 1 1941
2 77406 1 1941
2 77407 1 1943
2 77408 1 1943
2 77409 1 1946
2 77410 1 1946
2 77411 1 1946
2 77412 1 1946
2 77413 1 1946
2 77414 1 1946
2 77415 1 1946
2 77416 1 1946
2 77417 1 1946
2 77418 1 1946
2 77419 1 1946
2 77420 1 1946
2 77421 1 1946
2 77422 1 1946
2 77423 1 1946
2 77424 1 1946
2 77425 1 1946
2 77426 1 1946
2 77427 1 1946
2 77428 1 1946
2 77429 1 1946
2 77430 1 1946
2 77431 1 1946
2 77432 1 1946
2 77433 1 1946
2 77434 1 1946
2 77435 1 1946
2 77436 1 1946
2 77437 1 1946
2 77438 1 1946
2 77439 1 1946
2 77440 1 1946
2 77441 1 1946
2 77442 1 1946
2 77443 1 1947
2 77444 1 1947
2 77445 1 1947
2 77446 1 1947
2 77447 1 1947
2 77448 1 1947
2 77449 1 1948
2 77450 1 1948
2 77451 1 1954
2 77452 1 1954
2 77453 1 1954
2 77454 1 1954
2 77455 1 1954
2 77456 1 1954
2 77457 1 1954
2 77458 1 1954
2 77459 1 1954
2 77460 1 1954
2 77461 1 1954
2 77462 1 1954
2 77463 1 1954
2 77464 1 1954
2 77465 1 1954
2 77466 1 1954
2 77467 1 1954
2 77468 1 1954
2 77469 1 1954
2 77470 1 1954
2 77471 1 1954
2 77472 1 1954
2 77473 1 1954
2 77474 1 1954
2 77475 1 1954
2 77476 1 1954
2 77477 1 1954
2 77478 1 1954
2 77479 1 1954
2 77480 1 1954
2 77481 1 1954
2 77482 1 1954
2 77483 1 1954
2 77484 1 1954
2 77485 1 1954
2 77486 1 1954
2 77487 1 1954
2 77488 1 1954
2 77489 1 1954
2 77490 1 1954
2 77491 1 1954
2 77492 1 1954
2 77493 1 1954
2 77494 1 1955
2 77495 1 1955
2 77496 1 1955
2 77497 1 1955
2 77498 1 1955
2 77499 1 1955
2 77500 1 1955
2 77501 1 1955
2 77502 1 1955
2 77503 1 1955
2 77504 1 1955
2 77505 1 1955
2 77506 1 1955
2 77507 1 1955
2 77508 1 1955
2 77509 1 1955
2 77510 1 1955
2 77511 1 1956
2 77512 1 1956
2 77513 1 1956
2 77514 1 1956
2 77515 1 1956
2 77516 1 1956
2 77517 1 1956
2 77518 1 1956
2 77519 1 1957
2 77520 1 1957
2 77521 1 1958
2 77522 1 1958
2 77523 1 1959
2 77524 1 1959
2 77525 1 1966
2 77526 1 1966
2 77527 1 1966
2 77528 1 1966
2 77529 1 1966
2 77530 1 1966
2 77531 1 1968
2 77532 1 1968
2 77533 1 1968
2 77534 1 1968
2 77535 1 1968
2 77536 1 1968
2 77537 1 1968
2 77538 1 1985
2 77539 1 1985
2 77540 1 1985
2 77541 1 1985
2 77542 1 1985
2 77543 1 1985
2 77544 1 1985
2 77545 1 1985
2 77546 1 1985
2 77547 1 1985
2 77548 1 1985
2 77549 1 1985
2 77550 1 1985
2 77551 1 1985
2 77552 1 1985
2 77553 1 1985
2 77554 1 1985
2 77555 1 1985
2 77556 1 1985
2 77557 1 1985
2 77558 1 1985
2 77559 1 1985
2 77560 1 1985
2 77561 1 1985
2 77562 1 1985
2 77563 1 1985
2 77564 1 1985
2 77565 1 1985
2 77566 1 1985
2 77567 1 1985
2 77568 1 1985
2 77569 1 1985
2 77570 1 1985
2 77571 1 1985
2 77572 1 1985
2 77573 1 1985
2 77574 1 1985
2 77575 1 1985
2 77576 1 1985
2 77577 1 1985
2 77578 1 1985
2 77579 1 1985
2 77580 1 1985
2 77581 1 1985
2 77582 1 1985
2 77583 1 1985
2 77584 1 1985
2 77585 1 1985
2 77586 1 1985
2 77587 1 1985
2 77588 1 1986
2 77589 1 1986
2 77590 1 1986
2 77591 1 1986
2 77592 1 1986
2 77593 1 1986
2 77594 1 1986
2 77595 1 1986
2 77596 1 1986
2 77597 1 1986
2 77598 1 1986
2 77599 1 1986
2 77600 1 1986
2 77601 1 1986
2 77602 1 1986
2 77603 1 1986
2 77604 1 1986
2 77605 1 1986
2 77606 1 1986
2 77607 1 1986
2 77608 1 1986
2 77609 1 1986
2 77610 1 1986
2 77611 1 1987
2 77612 1 1987
2 77613 1 1987
2 77614 1 1987
2 77615 1 1987
2 77616 1 1987
2 77617 1 1987
2 77618 1 1989
2 77619 1 1989
2 77620 1 1990
2 77621 1 1990
2 77622 1 1991
2 77623 1 1991
2 77624 1 1991
2 77625 1 1991
2 77626 1 1991
2 77627 1 1999
2 77628 1 1999
2 77629 1 1999
2 77630 1 2006
2 77631 1 2006
2 77632 1 2006
2 77633 1 2006
2 77634 1 2007
2 77635 1 2007
2 77636 1 2007
2 77637 1 2007
2 77638 1 2009
2 77639 1 2009
2 77640 1 2009
2 77641 1 2009
2 77642 1 2009
2 77643 1 2009
2 77644 1 2010
2 77645 1 2010
2 77646 1 2010
2 77647 1 2011
2 77648 1 2011
2 77649 1 2020
2 77650 1 2020
2 77651 1 2040
2 77652 1 2040
2 77653 1 2043
2 77654 1 2043
2 77655 1 2045
2 77656 1 2045
2 77657 1 2045
2 77658 1 2045
2 77659 1 2045
2 77660 1 2045
2 77661 1 2046
2 77662 1 2046
2 77663 1 2059
2 77664 1 2059
2 77665 1 2059
2 77666 1 2059
2 77667 1 2059
2 77668 1 2059
2 77669 1 2060
2 77670 1 2060
2 77671 1 2060
2 77672 1 2060
2 77673 1 2062
2 77674 1 2062
2 77675 1 2063
2 77676 1 2063
2 77677 1 2063
2 77678 1 2064
2 77679 1 2064
2 77680 1 2067
2 77681 1 2067
2 77682 1 2077
2 77683 1 2077
2 77684 1 2078
2 77685 1 2078
2 77686 1 2078
2 77687 1 2078
2 77688 1 2078
2 77689 1 2078
2 77690 1 2078
2 77691 1 2078
2 77692 1 2078
2 77693 1 2078
2 77694 1 2078
2 77695 1 2079
2 77696 1 2079
2 77697 1 2079
2 77698 1 2079
2 77699 1 2079
2 77700 1 2079
2 77701 1 2079
2 77702 1 2079
2 77703 1 2079
2 77704 1 2079
2 77705 1 2079
2 77706 1 2079
2 77707 1 2079
2 77708 1 2079
2 77709 1 2080
2 77710 1 2080
2 77711 1 2081
2 77712 1 2081
2 77713 1 2081
2 77714 1 2081
2 77715 1 2081
2 77716 1 2082
2 77717 1 2082
2 77718 1 2082
2 77719 1 2082
2 77720 1 2084
2 77721 1 2084
2 77722 1 2084
2 77723 1 2084
2 77724 1 2085
2 77725 1 2085
2 77726 1 2085
2 77727 1 2085
2 77728 1 2085
2 77729 1 2085
2 77730 1 2085
2 77731 1 2085
2 77732 1 2085
2 77733 1 2085
2 77734 1 2085
2 77735 1 2085
2 77736 1 2085
2 77737 1 2085
2 77738 1 2085
2 77739 1 2085
2 77740 1 2085
2 77741 1 2085
2 77742 1 2085
2 77743 1 2085
2 77744 1 2085
2 77745 1 2085
2 77746 1 2085
2 77747 1 2086
2 77748 1 2086
2 77749 1 2086
2 77750 1 2086
2 77751 1 2086
2 77752 1 2087
2 77753 1 2087
2 77754 1 2087
2 77755 1 2098
2 77756 1 2098
2 77757 1 2098
2 77758 1 2098
2 77759 1 2098
2 77760 1 2098
2 77761 1 2098
2 77762 1 2098
2 77763 1 2098
2 77764 1 2098
2 77765 1 2098
2 77766 1 2098
2 77767 1 2098
2 77768 1 2098
2 77769 1 2098
2 77770 1 2098
2 77771 1 2098
2 77772 1 2098
2 77773 1 2098
2 77774 1 2098
2 77775 1 2098
2 77776 1 2098
2 77777 1 2098
2 77778 1 2098
2 77779 1 2098
2 77780 1 2098
2 77781 1 2098
2 77782 1 2098
2 77783 1 2098
2 77784 1 2098
2 77785 1 2098
2 77786 1 2098
2 77787 1 2098
2 77788 1 2098
2 77789 1 2098
2 77790 1 2098
2 77791 1 2098
2 77792 1 2098
2 77793 1 2098
2 77794 1 2098
2 77795 1 2098
2 77796 1 2098
2 77797 1 2098
2 77798 1 2098
2 77799 1 2098
2 77800 1 2098
2 77801 1 2098
2 77802 1 2098
2 77803 1 2098
2 77804 1 2099
2 77805 1 2099
2 77806 1 2099
2 77807 1 2099
2 77808 1 2100
2 77809 1 2100
2 77810 1 2100
2 77811 1 2100
2 77812 1 2101
2 77813 1 2101
2 77814 1 2103
2 77815 1 2103
2 77816 1 2103
2 77817 1 2103
2 77818 1 2104
2 77819 1 2104
2 77820 1 2107
2 77821 1 2107
2 77822 1 2116
2 77823 1 2116
2 77824 1 2116
2 77825 1 2116
2 77826 1 2116
2 77827 1 2116
2 77828 1 2116
2 77829 1 2116
2 77830 1 2116
2 77831 1 2116
2 77832 1 2116
2 77833 1 2116
2 77834 1 2116
2 77835 1 2116
2 77836 1 2116
2 77837 1 2116
2 77838 1 2117
2 77839 1 2117
2 77840 1 2117
2 77841 1 2117
2 77842 1 2117
2 77843 1 2118
2 77844 1 2118
2 77845 1 2118
2 77846 1 2118
2 77847 1 2119
2 77848 1 2119
2 77849 1 2128
2 77850 1 2128
2 77851 1 2128
2 77852 1 2128
2 77853 1 2128
2 77854 1 2128
2 77855 1 2128
2 77856 1 2128
2 77857 1 2128
2 77858 1 2128
2 77859 1 2128
2 77860 1 2128
2 77861 1 2128
2 77862 1 2128
2 77863 1 2128
2 77864 1 2128
2 77865 1 2128
2 77866 1 2128
2 77867 1 2128
2 77868 1 2128
2 77869 1 2128
2 77870 1 2128
2 77871 1 2128
2 77872 1 2129
2 77873 1 2129
2 77874 1 2130
2 77875 1 2130
2 77876 1 2130
2 77877 1 2131
2 77878 1 2131
2 77879 1 2131
2 77880 1 2131
2 77881 1 2131
2 77882 1 2131
2 77883 1 2131
2 77884 1 2131
2 77885 1 2131
2 77886 1 2131
2 77887 1 2131
2 77888 1 2131
2 77889 1 2131
2 77890 1 2131
2 77891 1 2131
2 77892 1 2131
2 77893 1 2131
2 77894 1 2131
2 77895 1 2131
2 77896 1 2131
2 77897 1 2131
2 77898 1 2131
2 77899 1 2131
2 77900 1 2131
2 77901 1 2131
2 77902 1 2131
2 77903 1 2131
2 77904 1 2131
2 77905 1 2131
2 77906 1 2131
2 77907 1 2131
2 77908 1 2131
2 77909 1 2131
2 77910 1 2131
2 77911 1 2131
2 77912 1 2131
2 77913 1 2131
2 77914 1 2131
2 77915 1 2131
2 77916 1 2131
2 77917 1 2131
2 77918 1 2131
2 77919 1 2131
2 77920 1 2131
2 77921 1 2131
2 77922 1 2131
2 77923 1 2131
2 77924 1 2131
2 77925 1 2131
2 77926 1 2131
2 77927 1 2131
2 77928 1 2131
2 77929 1 2131
2 77930 1 2131
2 77931 1 2131
2 77932 1 2131
2 77933 1 2131
2 77934 1 2131
2 77935 1 2131
2 77936 1 2131
2 77937 1 2131
2 77938 1 2132
2 77939 1 2132
2 77940 1 2132
2 77941 1 2132
2 77942 1 2132
2 77943 1 2132
2 77944 1 2132
2 77945 1 2132
2 77946 1 2132
2 77947 1 2132
2 77948 1 2132
2 77949 1 2133
2 77950 1 2133
2 77951 1 2135
2 77952 1 2135
2 77953 1 2141
2 77954 1 2141
2 77955 1 2141
2 77956 1 2141
2 77957 1 2144
2 77958 1 2144
2 77959 1 2144
2 77960 1 2144
2 77961 1 2144
2 77962 1 2144
2 77963 1 2144
2 77964 1 2144
2 77965 1 2144
2 77966 1 2144
2 77967 1 2144
2 77968 1 2144
2 77969 1 2144
2 77970 1 2144
2 77971 1 2144
2 77972 1 2144
2 77973 1 2144
2 77974 1 2144
2 77975 1 2144
2 77976 1 2145
2 77977 1 2145
2 77978 1 2145
2 77979 1 2145
2 77980 1 2145
2 77981 1 2145
2 77982 1 2153
2 77983 1 2153
2 77984 1 2153
2 77985 1 2153
2 77986 1 2153
2 77987 1 2153
2 77988 1 2153
2 77989 1 2153
2 77990 1 2153
2 77991 1 2153
2 77992 1 2153
2 77993 1 2153
2 77994 1 2153
2 77995 1 2154
2 77996 1 2154
2 77997 1 2154
2 77998 1 2154
2 77999 1 2154
2 78000 1 2155
2 78001 1 2155
2 78002 1 2155
2 78003 1 2155
2 78004 1 2155
2 78005 1 2155
2 78006 1 2155
2 78007 1 2155
2 78008 1 2155
2 78009 1 2155
2 78010 1 2156
2 78011 1 2156
2 78012 1 2156
2 78013 1 2156
2 78014 1 2157
2 78015 1 2157
2 78016 1 2157
2 78017 1 2157
2 78018 1 2157
2 78019 1 2167
2 78020 1 2167
2 78021 1 2167
2 78022 1 2168
2 78023 1 2168
2 78024 1 2168
2 78025 1 2169
2 78026 1 2169
2 78027 1 2169
2 78028 1 2169
2 78029 1 2169
2 78030 1 2169
2 78031 1 2169
2 78032 1 2169
2 78033 1 2169
2 78034 1 2169
2 78035 1 2169
2 78036 1 2170
2 78037 1 2170
2 78038 1 2170
2 78039 1 2170
2 78040 1 2170
2 78041 1 2170
2 78042 1 2171
2 78043 1 2171
2 78044 1 2171
2 78045 1 2172
2 78046 1 2172
2 78047 1 2191
2 78048 1 2191
2 78049 1 2191
2 78050 1 2191
2 78051 1 2191
2 78052 1 2191
2 78053 1 2191
2 78054 1 2191
2 78055 1 2191
2 78056 1 2191
2 78057 1 2191
2 78058 1 2191
2 78059 1 2191
2 78060 1 2191
2 78061 1 2191
2 78062 1 2191
2 78063 1 2191
2 78064 1 2191
2 78065 1 2191
2 78066 1 2191
2 78067 1 2191
2 78068 1 2192
2 78069 1 2192
2 78070 1 2192
2 78071 1 2192
2 78072 1 2192
2 78073 1 2193
2 78074 1 2193
2 78075 1 2193
2 78076 1 2194
2 78077 1 2194
2 78078 1 2194
2 78079 1 2194
2 78080 1 2194
2 78081 1 2196
2 78082 1 2196
2 78083 1 2199
2 78084 1 2199
2 78085 1 2205
2 78086 1 2205
2 78087 1 2205
2 78088 1 2205
2 78089 1 2206
2 78090 1 2206
2 78091 1 2213
2 78092 1 2213
2 78093 1 2214
2 78094 1 2214
2 78095 1 2214
2 78096 1 2221
2 78097 1 2221
2 78098 1 2222
2 78099 1 2222
2 78100 1 2222
2 78101 1 2223
2 78102 1 2223
2 78103 1 2225
2 78104 1 2225
2 78105 1 2229
2 78106 1 2229
2 78107 1 2229
2 78108 1 2229
2 78109 1 2229
2 78110 1 2229
2 78111 1 2229
2 78112 1 2229
2 78113 1 2230
2 78114 1 2230
2 78115 1 2230
2 78116 1 2230
2 78117 1 2230
2 78118 1 2231
2 78119 1 2231
2 78120 1 2231
2 78121 1 2231
2 78122 1 2231
2 78123 1 2231
2 78124 1 2231
2 78125 1 2231
2 78126 1 2231
2 78127 1 2231
2 78128 1 2231
2 78129 1 2231
2 78130 1 2231
2 78131 1 2231
2 78132 1 2231
2 78133 1 2231
2 78134 1 2231
2 78135 1 2231
2 78136 1 2231
2 78137 1 2231
2 78138 1 2231
2 78139 1 2231
2 78140 1 2231
2 78141 1 2231
2 78142 1 2232
2 78143 1 2232
2 78144 1 2232
2 78145 1 2232
2 78146 1 2232
2 78147 1 2232
2 78148 1 2232
2 78149 1 2232
2 78150 1 2232
2 78151 1 2233
2 78152 1 2233
2 78153 1 2233
2 78154 1 2233
2 78155 1 2233
2 78156 1 2233
2 78157 1 2233
2 78158 1 2233
2 78159 1 2233
2 78160 1 2233
2 78161 1 2233
2 78162 1 2233
2 78163 1 2233
2 78164 1 2233
2 78165 1 2233
2 78166 1 2234
2 78167 1 2234
2 78168 1 2238
2 78169 1 2238
2 78170 1 2243
2 78171 1 2243
2 78172 1 2243
2 78173 1 2243
2 78174 1 2243
2 78175 1 2243
2 78176 1 2243
2 78177 1 2243
2 78178 1 2243
2 78179 1 2243
2 78180 1 2243
2 78181 1 2243
2 78182 1 2243
2 78183 1 2243
2 78184 1 2243
2 78185 1 2243
2 78186 1 2243
2 78187 1 2243
2 78188 1 2243
2 78189 1 2243
2 78190 1 2243
2 78191 1 2243
2 78192 1 2243
2 78193 1 2243
2 78194 1 2243
2 78195 1 2243
2 78196 1 2243
2 78197 1 2243
2 78198 1 2243
2 78199 1 2243
2 78200 1 2243
2 78201 1 2243
2 78202 1 2243
2 78203 1 2244
2 78204 1 2244
2 78205 1 2244
2 78206 1 2244
2 78207 1 2245
2 78208 1 2245
2 78209 1 2245
2 78210 1 2245
2 78211 1 2245
2 78212 1 2246
2 78213 1 2246
2 78214 1 2246
2 78215 1 2249
2 78216 1 2249
2 78217 1 2249
2 78218 1 2249
2 78219 1 2249
2 78220 1 2249
2 78221 1 2250
2 78222 1 2250
2 78223 1 2250
2 78224 1 2250
2 78225 1 2250
2 78226 1 2250
2 78227 1 2250
2 78228 1 2250
2 78229 1 2253
2 78230 1 2253
2 78231 1 2270
2 78232 1 2270
2 78233 1 2273
2 78234 1 2273
2 78235 1 2273
2 78236 1 2274
2 78237 1 2274
2 78238 1 2274
2 78239 1 2274
2 78240 1 2281
2 78241 1 2281
2 78242 1 2281
2 78243 1 2281
2 78244 1 2281
2 78245 1 2281
2 78246 1 2281
2 78247 1 2281
2 78248 1 2281
2 78249 1 2281
2 78250 1 2281
2 78251 1 2281
2 78252 1 2281
2 78253 1 2281
2 78254 1 2281
2 78255 1 2281
2 78256 1 2281
2 78257 1 2281
2 78258 1 2281
2 78259 1 2281
2 78260 1 2281
2 78261 1 2281
2 78262 1 2281
2 78263 1 2281
2 78264 1 2281
2 78265 1 2281
2 78266 1 2281
2 78267 1 2281
2 78268 1 2282
2 78269 1 2282
2 78270 1 2282
2 78271 1 2282
2 78272 1 2282
2 78273 1 2282
2 78274 1 2282
2 78275 1 2282
2 78276 1 2282
2 78277 1 2282
2 78278 1 2282
2 78279 1 2283
2 78280 1 2283
2 78281 1 2283
2 78282 1 2283
2 78283 1 2283
2 78284 1 2292
2 78285 1 2292
2 78286 1 2292
2 78287 1 2292
2 78288 1 2292
2 78289 1 2292
2 78290 1 2292
2 78291 1 2292
2 78292 1 2292
2 78293 1 2292
2 78294 1 2293
2 78295 1 2293
2 78296 1 2293
2 78297 1 2293
2 78298 1 2293
2 78299 1 2293
2 78300 1 2294
2 78301 1 2294
2 78302 1 2294
2 78303 1 2294
2 78304 1 2302
2 78305 1 2302
2 78306 1 2303
2 78307 1 2303
2 78308 1 2304
2 78309 1 2304
2 78310 1 2304
2 78311 1 2304
2 78312 1 2305
2 78313 1 2305
2 78314 1 2305
2 78315 1 2305
2 78316 1 2305
2 78317 1 2305
2 78318 1 2307
2 78319 1 2307
2 78320 1 2307
2 78321 1 2307
2 78322 1 2307
2 78323 1 2321
2 78324 1 2321
2 78325 1 2324
2 78326 1 2324
2 78327 1 2326
2 78328 1 2326
2 78329 1 2326
2 78330 1 2326
2 78331 1 2326
2 78332 1 2327
2 78333 1 2327
2 78334 1 2327
2 78335 1 2327
2 78336 1 2328
2 78337 1 2328
2 78338 1 2332
2 78339 1 2332
2 78340 1 2332
2 78341 1 2332
2 78342 1 2333
2 78343 1 2333
2 78344 1 2333
2 78345 1 2333
2 78346 1 2333
2 78347 1 2333
2 78348 1 2333
2 78349 1 2333
2 78350 1 2333
2 78351 1 2333
2 78352 1 2338
2 78353 1 2338
2 78354 1 2338
2 78355 1 2338
2 78356 1 2339
2 78357 1 2339
2 78358 1 2339
2 78359 1 2339
2 78360 1 2339
2 78361 1 2339
2 78362 1 2339
2 78363 1 2354
2 78364 1 2354
2 78365 1 2354
2 78366 1 2354
2 78367 1 2354
2 78368 1 2354
2 78369 1 2354
2 78370 1 2354
2 78371 1 2354
2 78372 1 2354
2 78373 1 2354
2 78374 1 2354
2 78375 1 2354
2 78376 1 2354
2 78377 1 2354
2 78378 1 2354
2 78379 1 2354
2 78380 1 2354
2 78381 1 2354
2 78382 1 2354
2 78383 1 2354
2 78384 1 2354
2 78385 1 2355
2 78386 1 2355
2 78387 1 2355
2 78388 1 2355
2 78389 1 2355
2 78390 1 2355
2 78391 1 2357
2 78392 1 2357
2 78393 1 2357
2 78394 1 2357
2 78395 1 2361
2 78396 1 2361
2 78397 1 2361
2 78398 1 2361
2 78399 1 2361
2 78400 1 2361
2 78401 1 2361
2 78402 1 2361
2 78403 1 2370
2 78404 1 2370
2 78405 1 2370
2 78406 1 2370
2 78407 1 2370
2 78408 1 2370
2 78409 1 2370
2 78410 1 2371
2 78411 1 2371
2 78412 1 2371
2 78413 1 2371
2 78414 1 2371
2 78415 1 2371
2 78416 1 2371
2 78417 1 2372
2 78418 1 2372
2 78419 1 2372
2 78420 1 2373
2 78421 1 2373
2 78422 1 2373
2 78423 1 2373
2 78424 1 2373
2 78425 1 2373
2 78426 1 2373
2 78427 1 2376
2 78428 1 2376
2 78429 1 2380
2 78430 1 2380
2 78431 1 2390
2 78432 1 2390
2 78433 1 2390
2 78434 1 2390
2 78435 1 2390
2 78436 1 2390
2 78437 1 2390
2 78438 1 2390
2 78439 1 2390
2 78440 1 2391
2 78441 1 2391
2 78442 1 2391
2 78443 1 2391
2 78444 1 2391
2 78445 1 2392
2 78446 1 2392
2 78447 1 2401
2 78448 1 2401
2 78449 1 2406
2 78450 1 2406
2 78451 1 2407
2 78452 1 2407
2 78453 1 2409
2 78454 1 2409
2 78455 1 2420
2 78456 1 2420
2 78457 1 2421
2 78458 1 2421
2 78459 1 2421
2 78460 1 2421
2 78461 1 2421
2 78462 1 2421
2 78463 1 2421
2 78464 1 2421
2 78465 1 2421
2 78466 1 2423
2 78467 1 2423
2 78468 1 2424
2 78469 1 2424
2 78470 1 2424
2 78471 1 2425
2 78472 1 2425
2 78473 1 2425
2 78474 1 2425
2 78475 1 2425
2 78476 1 2425
2 78477 1 2425
2 78478 1 2425
2 78479 1 2425
2 78480 1 2425
2 78481 1 2425
2 78482 1 2425
2 78483 1 2425
2 78484 1 2426
2 78485 1 2426
2 78486 1 2426
2 78487 1 2426
2 78488 1 2427
2 78489 1 2427
2 78490 1 2427
2 78491 1 2428
2 78492 1 2428
2 78493 1 2430
2 78494 1 2430
2 78495 1 2434
2 78496 1 2434
2 78497 1 2437
2 78498 1 2437
2 78499 1 2441
2 78500 1 2441
2 78501 1 2441
2 78502 1 2441
2 78503 1 2442
2 78504 1 2442
2 78505 1 2443
2 78506 1 2443
2 78507 1 2443
2 78508 1 2443
2 78509 1 2443
2 78510 1 2443
2 78511 1 2443
2 78512 1 2443
2 78513 1 2443
2 78514 1 2443
2 78515 1 2443
2 78516 1 2445
2 78517 1 2445
2 78518 1 2445
2 78519 1 2453
2 78520 1 2453
2 78521 1 2453
2 78522 1 2453
2 78523 1 2453
2 78524 1 2453
2 78525 1 2453
2 78526 1 2453
2 78527 1 2453
2 78528 1 2453
2 78529 1 2453
2 78530 1 2453
2 78531 1 2453
2 78532 1 2453
2 78533 1 2453
2 78534 1 2453
2 78535 1 2453
2 78536 1 2455
2 78537 1 2455
2 78538 1 2455
2 78539 1 2456
2 78540 1 2456
2 78541 1 2456
2 78542 1 2467
2 78543 1 2467
2 78544 1 2467
2 78545 1 2467
2 78546 1 2467
2 78547 1 2467
2 78548 1 2467
2 78549 1 2467
2 78550 1 2467
2 78551 1 2467
2 78552 1 2467
2 78553 1 2467
2 78554 1 2467
2 78555 1 2467
2 78556 1 2467
2 78557 1 2467
2 78558 1 2467
2 78559 1 2467
2 78560 1 2467
2 78561 1 2467
2 78562 1 2467
2 78563 1 2467
2 78564 1 2467
2 78565 1 2467
2 78566 1 2467
2 78567 1 2467
2 78568 1 2467
2 78569 1 2467
2 78570 1 2467
2 78571 1 2467
2 78572 1 2467
2 78573 1 2467
2 78574 1 2467
2 78575 1 2467
2 78576 1 2467
2 78577 1 2467
2 78578 1 2467
2 78579 1 2467
2 78580 1 2467
2 78581 1 2467
2 78582 1 2468
2 78583 1 2468
2 78584 1 2468
2 78585 1 2468
2 78586 1 2468
2 78587 1 2468
2 78588 1 2468
2 78589 1 2468
2 78590 1 2468
2 78591 1 2468
2 78592 1 2468
2 78593 1 2468
2 78594 1 2468
2 78595 1 2468
2 78596 1 2468
2 78597 1 2468
2 78598 1 2468
2 78599 1 2468
2 78600 1 2468
2 78601 1 2468
2 78602 1 2468
2 78603 1 2468
2 78604 1 2468
2 78605 1 2469
2 78606 1 2469
2 78607 1 2471
2 78608 1 2471
2 78609 1 2471
2 78610 1 2471
2 78611 1 2471
2 78612 1 2472
2 78613 1 2472
2 78614 1 2472
2 78615 1 2472
2 78616 1 2473
2 78617 1 2473
2 78618 1 2473
2 78619 1 2473
2 78620 1 2473
2 78621 1 2473
2 78622 1 2473
2 78623 1 2473
2 78624 1 2473
2 78625 1 2473
2 78626 1 2473
2 78627 1 2473
2 78628 1 2474
2 78629 1 2474
2 78630 1 2474
2 78631 1 2474
2 78632 1 2474
2 78633 1 2475
2 78634 1 2475
2 78635 1 2475
2 78636 1 2475
2 78637 1 2475
2 78638 1 2476
2 78639 1 2476
2 78640 1 2476
2 78641 1 2476
2 78642 1 2477
2 78643 1 2477
2 78644 1 2478
2 78645 1 2478
2 78646 1 2478
2 78647 1 2478
2 78648 1 2480
2 78649 1 2480
2 78650 1 2483
2 78651 1 2483
2 78652 1 2484
2 78653 1 2484
2 78654 1 2484
2 78655 1 2484
2 78656 1 2484
2 78657 1 2484
2 78658 1 2484
2 78659 1 2484
2 78660 1 2484
2 78661 1 2484
2 78662 1 2484
2 78663 1 2484
2 78664 1 2484
2 78665 1 2484
2 78666 1 2484
2 78667 1 2484
2 78668 1 2484
2 78669 1 2484
2 78670 1 2484
2 78671 1 2484
2 78672 1 2484
2 78673 1 2484
2 78674 1 2485
2 78675 1 2485
2 78676 1 2490
2 78677 1 2490
2 78678 1 2494
2 78679 1 2494
2 78680 1 2494
2 78681 1 2494
2 78682 1 2494
2 78683 1 2494
2 78684 1 2495
2 78685 1 2495
2 78686 1 2495
2 78687 1 2495
2 78688 1 2496
2 78689 1 2496
2 78690 1 2500
2 78691 1 2500
2 78692 1 2500
2 78693 1 2500
2 78694 1 2500
2 78695 1 2500
2 78696 1 2500
2 78697 1 2500
2 78698 1 2500
2 78699 1 2500
2 78700 1 2500
2 78701 1 2500
2 78702 1 2500
2 78703 1 2500
2 78704 1 2500
2 78705 1 2500
2 78706 1 2500
2 78707 1 2500
2 78708 1 2500
2 78709 1 2500
2 78710 1 2500
2 78711 1 2500
2 78712 1 2500
2 78713 1 2500
2 78714 1 2501
2 78715 1 2501
2 78716 1 2501
2 78717 1 2501
2 78718 1 2502
2 78719 1 2502
2 78720 1 2511
2 78721 1 2511
2 78722 1 2512
2 78723 1 2512
2 78724 1 2513
2 78725 1 2513
2 78726 1 2514
2 78727 1 2514
2 78728 1 2514
2 78729 1 2525
2 78730 1 2525
2 78731 1 2546
2 78732 1 2546
2 78733 1 2546
2 78734 1 2546
2 78735 1 2546
2 78736 1 2546
2 78737 1 2546
2 78738 1 2546
2 78739 1 2546
2 78740 1 2546
2 78741 1 2546
2 78742 1 2546
2 78743 1 2546
2 78744 1 2546
2 78745 1 2546
2 78746 1 2546
2 78747 1 2546
2 78748 1 2546
2 78749 1 2546
2 78750 1 2546
2 78751 1 2546
2 78752 1 2546
2 78753 1 2546
2 78754 1 2546
2 78755 1 2546
2 78756 1 2546
2 78757 1 2546
2 78758 1 2546
2 78759 1 2546
2 78760 1 2546
2 78761 1 2546
2 78762 1 2546
2 78763 1 2546
2 78764 1 2546
2 78765 1 2546
2 78766 1 2546
2 78767 1 2546
2 78768 1 2546
2 78769 1 2546
2 78770 1 2546
2 78771 1 2546
2 78772 1 2546
2 78773 1 2546
2 78774 1 2546
2 78775 1 2546
2 78776 1 2546
2 78777 1 2546
2 78778 1 2546
2 78779 1 2546
2 78780 1 2546
2 78781 1 2546
2 78782 1 2546
2 78783 1 2546
2 78784 1 2546
2 78785 1 2546
2 78786 1 2546
2 78787 1 2546
2 78788 1 2546
2 78789 1 2547
2 78790 1 2547
2 78791 1 2547
2 78792 1 2547
2 78793 1 2548
2 78794 1 2548
2 78795 1 2548
2 78796 1 2548
2 78797 1 2548
2 78798 1 2548
2 78799 1 2548
2 78800 1 2548
2 78801 1 2548
2 78802 1 2548
2 78803 1 2548
2 78804 1 2548
2 78805 1 2548
2 78806 1 2548
2 78807 1 2548
2 78808 1 2549
2 78809 1 2549
2 78810 1 2549
2 78811 1 2550
2 78812 1 2550
2 78813 1 2551
2 78814 1 2551
2 78815 1 2552
2 78816 1 2552
2 78817 1 2553
2 78818 1 2553
2 78819 1 2558
2 78820 1 2558
2 78821 1 2558
2 78822 1 2561
2 78823 1 2561
2 78824 1 2566
2 78825 1 2566
2 78826 1 2576
2 78827 1 2576
2 78828 1 2576
2 78829 1 2576
2 78830 1 2576
2 78831 1 2577
2 78832 1 2577
2 78833 1 2577
2 78834 1 2577
2 78835 1 2577
2 78836 1 2586
2 78837 1 2586
2 78838 1 2586
2 78839 1 2586
2 78840 1 2586
2 78841 1 2587
2 78842 1 2587
2 78843 1 2587
2 78844 1 2593
2 78845 1 2593
2 78846 1 2601
2 78847 1 2601
2 78848 1 2601
2 78849 1 2601
2 78850 1 2602
2 78851 1 2602
2 78852 1 2603
2 78853 1 2603
2 78854 1 2603
2 78855 1 2603
2 78856 1 2604
2 78857 1 2604
2 78858 1 2604
2 78859 1 2604
2 78860 1 2604
2 78861 1 2605
2 78862 1 2605
2 78863 1 2605
2 78864 1 2605
2 78865 1 2605
2 78866 1 2605
2 78867 1 2605
2 78868 1 2605
2 78869 1 2605
2 78870 1 2605
2 78871 1 2605
2 78872 1 2605
2 78873 1 2605
2 78874 1 2605
2 78875 1 2606
2 78876 1 2606
2 78877 1 2606
2 78878 1 2607
2 78879 1 2607
2 78880 1 2607
2 78881 1 2607
2 78882 1 2607
2 78883 1 2614
2 78884 1 2614
2 78885 1 2614
2 78886 1 2614
2 78887 1 2614
2 78888 1 2614
2 78889 1 2614
2 78890 1 2616
2 78891 1 2616
2 78892 1 2616
2 78893 1 2616
2 78894 1 2617
2 78895 1 2617
2 78896 1 2617
2 78897 1 2617
2 78898 1 2617
2 78899 1 2625
2 78900 1 2625
2 78901 1 2628
2 78902 1 2628
2 78903 1 2628
2 78904 1 2628
2 78905 1 2628
2 78906 1 2629
2 78907 1 2629
2 78908 1 2629
2 78909 1 2629
2 78910 1 2629
2 78911 1 2629
2 78912 1 2629
2 78913 1 2629
2 78914 1 2629
2 78915 1 2630
2 78916 1 2630
2 78917 1 2630
2 78918 1 2631
2 78919 1 2631
2 78920 1 2643
2 78921 1 2643
2 78922 1 2643
2 78923 1 2643
2 78924 1 2644
2 78925 1 2644
2 78926 1 2647
2 78927 1 2647
2 78928 1 2647
2 78929 1 2647
2 78930 1 2647
2 78931 1 2647
2 78932 1 2647
2 78933 1 2647
2 78934 1 2647
2 78935 1 2647
2 78936 1 2648
2 78937 1 2648
2 78938 1 2648
2 78939 1 2648
2 78940 1 2648
2 78941 1 2648
2 78942 1 2649
2 78943 1 2649
2 78944 1 2649
2 78945 1 2649
2 78946 1 2651
2 78947 1 2651
2 78948 1 2668
2 78949 1 2668
2 78950 1 2668
2 78951 1 2668
2 78952 1 2668
2 78953 1 2668
2 78954 1 2669
2 78955 1 2669
2 78956 1 2669
2 78957 1 2669
2 78958 1 2671
2 78959 1 2671
2 78960 1 2671
2 78961 1 2671
2 78962 1 2671
2 78963 1 2671
2 78964 1 2671
2 78965 1 2671
2 78966 1 2671
2 78967 1 2671
2 78968 1 2671
2 78969 1 2671
2 78970 1 2671
2 78971 1 2671
2 78972 1 2671
2 78973 1 2671
2 78974 1 2671
2 78975 1 2672
2 78976 1 2672
2 78977 1 2682
2 78978 1 2682
2 78979 1 2683
2 78980 1 2683
2 78981 1 2683
2 78982 1 2686
2 78983 1 2686
2 78984 1 2686
2 78985 1 2688
2 78986 1 2688
2 78987 1 2700
2 78988 1 2700
2 78989 1 2700
2 78990 1 2700
2 78991 1 2700
2 78992 1 2700
2 78993 1 2700
2 78994 1 2700
2 78995 1 2700
2 78996 1 2702
2 78997 1 2702
2 78998 1 2702
2 78999 1 2703
2 79000 1 2703
2 79001 1 2703
2 79002 1 2703
2 79003 1 2703
2 79004 1 2703
2 79005 1 2703
2 79006 1 2703
2 79007 1 2703
2 79008 1 2703
2 79009 1 2703
2 79010 1 2703
2 79011 1 2703
2 79012 1 2703
2 79013 1 2703
2 79014 1 2703
2 79015 1 2703
2 79016 1 2703
2 79017 1 2703
2 79018 1 2703
2 79019 1 2703
2 79020 1 2703
2 79021 1 2703
2 79022 1 2703
2 79023 1 2703
2 79024 1 2703
2 79025 1 2703
2 79026 1 2705
2 79027 1 2705
2 79028 1 2713
2 79029 1 2713
2 79030 1 2713
2 79031 1 2713
2 79032 1 2713
2 79033 1 2713
2 79034 1 2713
2 79035 1 2713
2 79036 1 2713
2 79037 1 2713
2 79038 1 2713
2 79039 1 2713
2 79040 1 2713
2 79041 1 2713
2 79042 1 2713
2 79043 1 2713
2 79044 1 2713
2 79045 1 2713
2 79046 1 2713
2 79047 1 2713
2 79048 1 2713
2 79049 1 2714
2 79050 1 2714
2 79051 1 2714
2 79052 1 2714
2 79053 1 2714
2 79054 1 2714
2 79055 1 2714
2 79056 1 2714
2 79057 1 2714
2 79058 1 2714
2 79059 1 2719
2 79060 1 2719
2 79061 1 2719
2 79062 1 2719
2 79063 1 2719
2 79064 1 2719
2 79065 1 2719
2 79066 1 2719
2 79067 1 2719
2 79068 1 2719
2 79069 1 2719
2 79070 1 2721
2 79071 1 2721
2 79072 1 2721
2 79073 1 2729
2 79074 1 2729
2 79075 1 2729
2 79076 1 2729
2 79077 1 2729
2 79078 1 2730
2 79079 1 2730
2 79080 1 2739
2 79081 1 2739
2 79082 1 2742
2 79083 1 2742
2 79084 1 2742
2 79085 1 2742
2 79086 1 2742
2 79087 1 2742
2 79088 1 2743
2 79089 1 2743
2 79090 1 2743
2 79091 1 2747
2 79092 1 2747
2 79093 1 2761
2 79094 1 2761
2 79095 1 2769
2 79096 1 2769
2 79097 1 2769
2 79098 1 2769
2 79099 1 2769
2 79100 1 2769
2 79101 1 2769
2 79102 1 2769
2 79103 1 2769
2 79104 1 2769
2 79105 1 2769
2 79106 1 2771
2 79107 1 2771
2 79108 1 2773
2 79109 1 2773
2 79110 1 2775
2 79111 1 2775
2 79112 1 2775
2 79113 1 2776
2 79114 1 2776
2 79115 1 2777
2 79116 1 2777
2 79117 1 2777
2 79118 1 2790
2 79119 1 2790
2 79120 1 2790
2 79121 1 2790
2 79122 1 2790
2 79123 1 2790
2 79124 1 2790
2 79125 1 2790
2 79126 1 2791
2 79127 1 2791
2 79128 1 2815
2 79129 1 2815
2 79130 1 2815
2 79131 1 2815
2 79132 1 2815
2 79133 1 2815
2 79134 1 2815
2 79135 1 2815
2 79136 1 2815
2 79137 1 2815
2 79138 1 2815
2 79139 1 2815
2 79140 1 2815
2 79141 1 2815
2 79142 1 2815
2 79143 1 2815
2 79144 1 2815
2 79145 1 2816
2 79146 1 2816
2 79147 1 2816
2 79148 1 2816
2 79149 1 2816
2 79150 1 2817
2 79151 1 2817
2 79152 1 2824
2 79153 1 2824
2 79154 1 2841
2 79155 1 2841
2 79156 1 2841
2 79157 1 2842
2 79158 1 2842
2 79159 1 2842
2 79160 1 2849
2 79161 1 2849
2 79162 1 2850
2 79163 1 2850
2 79164 1 2862
2 79165 1 2862
2 79166 1 2862
2 79167 1 2871
2 79168 1 2871
2 79169 1 2897
2 79170 1 2897
2 79171 1 2897
2 79172 1 2897
2 79173 1 2898
2 79174 1 2898
2 79175 1 2918
2 79176 1 2918
2 79177 1 2921
2 79178 1 2921
2 79179 1 2921
2 79180 1 2922
2 79181 1 2922
2 79182 1 2922
2 79183 1 2922
2 79184 1 2922
2 79185 1 2922
2 79186 1 2935
2 79187 1 2935
2 79188 1 2935
2 79189 1 2935
2 79190 1 2935
2 79191 1 2935
2 79192 1 2935
2 79193 1 2937
2 79194 1 2937
2 79195 1 2951
2 79196 1 2951
2 79197 1 2951
2 79198 1 2951
2 79199 1 2951
2 79200 1 2951
2 79201 1 2951
2 79202 1 2951
2 79203 1 2951
2 79204 1 2951
2 79205 1 2951
2 79206 1 2951
2 79207 1 2951
2 79208 1 2951
2 79209 1 2951
2 79210 1 2951
2 79211 1 2951
2 79212 1 2951
2 79213 1 2952
2 79214 1 2952
2 79215 1 2952
2 79216 1 2957
2 79217 1 2957
2 79218 1 2958
2 79219 1 2958
2 79220 1 2959
2 79221 1 2959
2 79222 1 2959
2 79223 1 2966
2 79224 1 2966
2 79225 1 2966
2 79226 1 2967
2 79227 1 2967
2 79228 1 2987
2 79229 1 2987
2 79230 1 2987
2 79231 1 2987
2 79232 1 2987
2 79233 1 2987
2 79234 1 2987
2 79235 1 2987
2 79236 1 2988
2 79237 1 2988
2 79238 1 2991
2 79239 1 2991
2 79240 1 2992
2 79241 1 2992
2 79242 1 2992
2 79243 1 2992
2 79244 1 2992
2 79245 1 2993
2 79246 1 2993
2 79247 1 2994
2 79248 1 2994
2 79249 1 2994
2 79250 1 2994
2 79251 1 2994
2 79252 1 2994
2 79253 1 2994
2 79254 1 2994
2 79255 1 2994
2 79256 1 2994
2 79257 1 2994
2 79258 1 2994
2 79259 1 2994
2 79260 1 2994
2 79261 1 2994
2 79262 1 2994
2 79263 1 2994
2 79264 1 2994
2 79265 1 2994
2 79266 1 2994
2 79267 1 2994
2 79268 1 2994
2 79269 1 2994
2 79270 1 2994
2 79271 1 2994
2 79272 1 2994
2 79273 1 2995
2 79274 1 2995
2 79275 1 2995
2 79276 1 2997
2 79277 1 2997
2 79278 1 2997
2 79279 1 2997
2 79280 1 2997
2 79281 1 2997
2 79282 1 2998
2 79283 1 2998
2 79284 1 2998
2 79285 1 2998
2 79286 1 2998
2 79287 1 2998
2 79288 1 2998
2 79289 1 2998
2 79290 1 2998
2 79291 1 2998
2 79292 1 2998
2 79293 1 2998
2 79294 1 2998
2 79295 1 2998
2 79296 1 2998
2 79297 1 2999
2 79298 1 2999
2 79299 1 3000
2 79300 1 3000
2 79301 1 3000
2 79302 1 3001
2 79303 1 3001
2 79304 1 3001
2 79305 1 3006
2 79306 1 3006
2 79307 1 3006
2 79308 1 3006
2 79309 1 3006
2 79310 1 3006
2 79311 1 3007
2 79312 1 3007
2 79313 1 3007
2 79314 1 3007
2 79315 1 3007
2 79316 1 3007
2 79317 1 3007
2 79318 1 3007
2 79319 1 3007
2 79320 1 3007
2 79321 1 3007
2 79322 1 3007
2 79323 1 3007
2 79324 1 3007
2 79325 1 3007
2 79326 1 3007
2 79327 1 3007
2 79328 1 3007
2 79329 1 3007
2 79330 1 3007
2 79331 1 3007
2 79332 1 3007
2 79333 1 3007
2 79334 1 3007
2 79335 1 3007
2 79336 1 3008
2 79337 1 3008
2 79338 1 3014
2 79339 1 3014
2 79340 1 3014
2 79341 1 3014
2 79342 1 3014
2 79343 1 3014
2 79344 1 3014
2 79345 1 3015
2 79346 1 3015
2 79347 1 3015
2 79348 1 3015
2 79349 1 3015
2 79350 1 3015
2 79351 1 3016
2 79352 1 3016
2 79353 1 3021
2 79354 1 3021
2 79355 1 3021
2 79356 1 3021
2 79357 1 3029
2 79358 1 3029
2 79359 1 3029
2 79360 1 3029
2 79361 1 3029
2 79362 1 3029
2 79363 1 3029
2 79364 1 3029
2 79365 1 3029
2 79366 1 3030
2 79367 1 3030
2 79368 1 3030
2 79369 1 3030
2 79370 1 3030
2 79371 1 3030
2 79372 1 3030
2 79373 1 3030
2 79374 1 3030
2 79375 1 3030
2 79376 1 3030
2 79377 1 3030
2 79378 1 3030
2 79379 1 3030
2 79380 1 3030
2 79381 1 3030
2 79382 1 3030
2 79383 1 3030
2 79384 1 3031
2 79385 1 3031
2 79386 1 3031
2 79387 1 3031
2 79388 1 3031
2 79389 1 3032
2 79390 1 3032
2 79391 1 3034
2 79392 1 3034
2 79393 1 3034
2 79394 1 3034
2 79395 1 3034
2 79396 1 3035
2 79397 1 3035
2 79398 1 3035
2 79399 1 3035
2 79400 1 3035
2 79401 1 3035
2 79402 1 3035
2 79403 1 3035
2 79404 1 3035
2 79405 1 3035
2 79406 1 3035
2 79407 1 3037
2 79408 1 3037
2 79409 1 3037
2 79410 1 3048
2 79411 1 3048
2 79412 1 3048
2 79413 1 3050
2 79414 1 3050
2 79415 1 3050
2 79416 1 3051
2 79417 1 3051
2 79418 1 3051
2 79419 1 3051
2 79420 1 3051
2 79421 1 3051
2 79422 1 3054
2 79423 1 3054
2 79424 1 3055
2 79425 1 3055
2 79426 1 3055
2 79427 1 3064
2 79428 1 3064
2 79429 1 3064
2 79430 1 3064
2 79431 1 3064
2 79432 1 3064
2 79433 1 3064
2 79434 1 3064
2 79435 1 3064
2 79436 1 3064
2 79437 1 3064
2 79438 1 3064
2 79439 1 3064
2 79440 1 3064
2 79441 1 3064
2 79442 1 3064
2 79443 1 3064
2 79444 1 3064
2 79445 1 3064
2 79446 1 3064
2 79447 1 3064
2 79448 1 3064
2 79449 1 3064
2 79450 1 3064
2 79451 1 3064
2 79452 1 3064
2 79453 1 3064
2 79454 1 3064
2 79455 1 3064
2 79456 1 3065
2 79457 1 3065
2 79458 1 3065
2 79459 1 3065
2 79460 1 3066
2 79461 1 3066
2 79462 1 3066
2 79463 1 3069
2 79464 1 3069
2 79465 1 3069
2 79466 1 3069
2 79467 1 3069
2 79468 1 3069
2 79469 1 3069
2 79470 1 3069
2 79471 1 3069
2 79472 1 3070
2 79473 1 3070
2 79474 1 3070
2 79475 1 3071
2 79476 1 3071
2 79477 1 3071
2 79478 1 3071
2 79479 1 3071
2 79480 1 3071
2 79481 1 3071
2 79482 1 3071
2 79483 1 3071
2 79484 1 3071
2 79485 1 3071
2 79486 1 3071
2 79487 1 3071
2 79488 1 3071
2 79489 1 3071
2 79490 1 3071
2 79491 1 3071
2 79492 1 3071
2 79493 1 3071
2 79494 1 3071
2 79495 1 3072
2 79496 1 3072
2 79497 1 3072
2 79498 1 3072
2 79499 1 3082
2 79500 1 3082
2 79501 1 3082
2 79502 1 3082
2 79503 1 3082
2 79504 1 3082
2 79505 1 3082
2 79506 1 3082
2 79507 1 3082
2 79508 1 3082
2 79509 1 3082
2 79510 1 3082
2 79511 1 3082
2 79512 1 3082
2 79513 1 3082
2 79514 1 3082
2 79515 1 3082
2 79516 1 3082
2 79517 1 3082
2 79518 1 3082
2 79519 1 3082
2 79520 1 3082
2 79521 1 3082
2 79522 1 3082
2 79523 1 3082
2 79524 1 3082
2 79525 1 3082
2 79526 1 3082
2 79527 1 3090
2 79528 1 3090
2 79529 1 3090
2 79530 1 3090
2 79531 1 3090
2 79532 1 3090
2 79533 1 3090
2 79534 1 3090
2 79535 1 3090
2 79536 1 3090
2 79537 1 3090
2 79538 1 3090
2 79539 1 3090
2 79540 1 3090
2 79541 1 3090
2 79542 1 3090
2 79543 1 3092
2 79544 1 3092
2 79545 1 3092
2 79546 1 3092
2 79547 1 3092
2 79548 1 3103
2 79549 1 3103
2 79550 1 3103
2 79551 1 3103
2 79552 1 3103
2 79553 1 3103
2 79554 1 3103
2 79555 1 3103
2 79556 1 3103
2 79557 1 3103
2 79558 1 3103
2 79559 1 3103
2 79560 1 3103
2 79561 1 3103
2 79562 1 3103
2 79563 1 3103
2 79564 1 3103
2 79565 1 3104
2 79566 1 3104
2 79567 1 3105
2 79568 1 3105
2 79569 1 3105
2 79570 1 3105
2 79571 1 3105
2 79572 1 3105
2 79573 1 3129
2 79574 1 3129
2 79575 1 3129
2 79576 1 3135
2 79577 1 3135
2 79578 1 3135
2 79579 1 3135
2 79580 1 3150
2 79581 1 3150
2 79582 1 3155
2 79583 1 3155
2 79584 1 3155
2 79585 1 3155
2 79586 1 3155
2 79587 1 3155
2 79588 1 3155
2 79589 1 3155
2 79590 1 3155
2 79591 1 3155
2 79592 1 3155
2 79593 1 3157
2 79594 1 3157
2 79595 1 3157
2 79596 1 3158
2 79597 1 3158
2 79598 1 3158
2 79599 1 3162
2 79600 1 3162
2 79601 1 3162
2 79602 1 3165
2 79603 1 3165
2 79604 1 3171
2 79605 1 3171
2 79606 1 3171
2 79607 1 3171
2 79608 1 3171
2 79609 1 3171
2 79610 1 3171
2 79611 1 3171
2 79612 1 3171
2 79613 1 3171
2 79614 1 3171
2 79615 1 3171
2 79616 1 3171
2 79617 1 3171
2 79618 1 3171
2 79619 1 3171
2 79620 1 3171
2 79621 1 3171
2 79622 1 3171
2 79623 1 3171
2 79624 1 3171
2 79625 1 3171
2 79626 1 3171
2 79627 1 3171
2 79628 1 3171
2 79629 1 3171
2 79630 1 3171
2 79631 1 3171
2 79632 1 3171
2 79633 1 3171
2 79634 1 3171
2 79635 1 3171
2 79636 1 3171
2 79637 1 3171
2 79638 1 3171
2 79639 1 3171
2 79640 1 3171
2 79641 1 3171
2 79642 1 3172
2 79643 1 3172
2 79644 1 3172
2 79645 1 3172
2 79646 1 3172
2 79647 1 3172
2 79648 1 3172
2 79649 1 3172
2 79650 1 3172
2 79651 1 3172
2 79652 1 3172
2 79653 1 3172
2 79654 1 3172
2 79655 1 3172
2 79656 1 3172
2 79657 1 3172
2 79658 1 3172
2 79659 1 3172
2 79660 1 3172
2 79661 1 3172
2 79662 1 3172
2 79663 1 3172
2 79664 1 3172
2 79665 1 3172
2 79666 1 3172
2 79667 1 3172
2 79668 1 3172
2 79669 1 3172
2 79670 1 3172
2 79671 1 3172
2 79672 1 3172
2 79673 1 3172
2 79674 1 3172
2 79675 1 3172
2 79676 1 3172
2 79677 1 3172
2 79678 1 3172
2 79679 1 3172
2 79680 1 3172
2 79681 1 3172
2 79682 1 3172
2 79683 1 3172
2 79684 1 3172
2 79685 1 3172
2 79686 1 3172
2 79687 1 3172
2 79688 1 3172
2 79689 1 3172
2 79690 1 3172
2 79691 1 3172
2 79692 1 3172
2 79693 1 3172
2 79694 1 3172
2 79695 1 3172
2 79696 1 3173
2 79697 1 3173
2 79698 1 3173
2 79699 1 3173
2 79700 1 3173
2 79701 1 3173
2 79702 1 3173
2 79703 1 3173
2 79704 1 3174
2 79705 1 3174
2 79706 1 3174
2 79707 1 3174
2 79708 1 3174
2 79709 1 3174
2 79710 1 3174
2 79711 1 3174
2 79712 1 3174
2 79713 1 3174
2 79714 1 3174
2 79715 1 3174
2 79716 1 3174
2 79717 1 3174
2 79718 1 3174
2 79719 1 3174
2 79720 1 3174
2 79721 1 3174
2 79722 1 3174
2 79723 1 3174
2 79724 1 3174
2 79725 1 3174
2 79726 1 3176
2 79727 1 3176
2 79728 1 3176
2 79729 1 3176
2 79730 1 3176
2 79731 1 3176
2 79732 1 3176
2 79733 1 3177
2 79734 1 3177
2 79735 1 3177
2 79736 1 3187
2 79737 1 3187
2 79738 1 3187
2 79739 1 3187
2 79740 1 3187
2 79741 1 3187
2 79742 1 3187
2 79743 1 3187
2 79744 1 3187
2 79745 1 3187
2 79746 1 3187
2 79747 1 3187
2 79748 1 3187
2 79749 1 3187
2 79750 1 3187
2 79751 1 3187
2 79752 1 3187
2 79753 1 3187
2 79754 1 3187
2 79755 1 3189
2 79756 1 3189
2 79757 1 3189
2 79758 1 3190
2 79759 1 3190
2 79760 1 3193
2 79761 1 3193
2 79762 1 3193
2 79763 1 3193
2 79764 1 3193
2 79765 1 3193
2 79766 1 3193
2 79767 1 3193
2 79768 1 3193
2 79769 1 3193
2 79770 1 3193
2 79771 1 3193
2 79772 1 3193
2 79773 1 3193
2 79774 1 3193
2 79775 1 3193
2 79776 1 3193
2 79777 1 3193
2 79778 1 3193
2 79779 1 3193
2 79780 1 3193
2 79781 1 3193
2 79782 1 3193
2 79783 1 3193
2 79784 1 3193
2 79785 1 3193
2 79786 1 3193
2 79787 1 3193
2 79788 1 3193
2 79789 1 3193
2 79790 1 3193
2 79791 1 3193
2 79792 1 3193
2 79793 1 3193
2 79794 1 3193
2 79795 1 3193
2 79796 1 3193
2 79797 1 3193
2 79798 1 3193
2 79799 1 3194
2 79800 1 3194
2 79801 1 3194
2 79802 1 3194
2 79803 1 3194
2 79804 1 3194
2 79805 1 3194
2 79806 1 3194
2 79807 1 3194
2 79808 1 3194
2 79809 1 3194
2 79810 1 3194
2 79811 1 3194
2 79812 1 3194
2 79813 1 3194
2 79814 1 3194
2 79815 1 3194
2 79816 1 3194
2 79817 1 3194
2 79818 1 3194
2 79819 1 3194
2 79820 1 3194
2 79821 1 3194
2 79822 1 3194
2 79823 1 3201
2 79824 1 3201
2 79825 1 3201
2 79826 1 3201
2 79827 1 3201
2 79828 1 3201
2 79829 1 3202
2 79830 1 3202
2 79831 1 3210
2 79832 1 3210
2 79833 1 3210
2 79834 1 3210
2 79835 1 3210
2 79836 1 3211
2 79837 1 3211
2 79838 1 3211
2 79839 1 3211
2 79840 1 3211
2 79841 1 3215
2 79842 1 3215
2 79843 1 3215
2 79844 1 3215
2 79845 1 3215
2 79846 1 3215
2 79847 1 3216
2 79848 1 3216
2 79849 1 3216
2 79850 1 3216
2 79851 1 3216
2 79852 1 3216
2 79853 1 3241
2 79854 1 3241
2 79855 1 3241
2 79856 1 3241
2 79857 1 3241
2 79858 1 3241
2 79859 1 3241
2 79860 1 3241
2 79861 1 3241
2 79862 1 3241
2 79863 1 3242
2 79864 1 3242
2 79865 1 3243
2 79866 1 3243
2 79867 1 3245
2 79868 1 3245
2 79869 1 3245
2 79870 1 3245
2 79871 1 3246
2 79872 1 3246
2 79873 1 3253
2 79874 1 3253
2 79875 1 3253
2 79876 1 3253
2 79877 1 3253
2 79878 1 3253
2 79879 1 3253
2 79880 1 3253
2 79881 1 3253
2 79882 1 3253
2 79883 1 3253
2 79884 1 3253
2 79885 1 3253
2 79886 1 3253
2 79887 1 3253
2 79888 1 3253
2 79889 1 3253
2 79890 1 3253
2 79891 1 3253
2 79892 1 3253
2 79893 1 3253
2 79894 1 3253
2 79895 1 3253
2 79896 1 3253
2 79897 1 3253
2 79898 1 3254
2 79899 1 3254
2 79900 1 3254
2 79901 1 3254
2 79902 1 3254
2 79903 1 3254
2 79904 1 3255
2 79905 1 3255
2 79906 1 3255
2 79907 1 3255
2 79908 1 3255
2 79909 1 3255
2 79910 1 3255
2 79911 1 3255
2 79912 1 3255
2 79913 1 3262
2 79914 1 3262
2 79915 1 3262
2 79916 1 3262
2 79917 1 3262
2 79918 1 3262
2 79919 1 3263
2 79920 1 3263
2 79921 1 3263
2 79922 1 3263
2 79923 1 3263
2 79924 1 3263
2 79925 1 3263
2 79926 1 3263
2 79927 1 3268
2 79928 1 3268
2 79929 1 3269
2 79930 1 3269
2 79931 1 3269
2 79932 1 3269
2 79933 1 3270
2 79934 1 3270
2 79935 1 3272
2 79936 1 3272
2 79937 1 3280
2 79938 1 3280
2 79939 1 3280
2 79940 1 3280
2 79941 1 3281
2 79942 1 3281
2 79943 1 3281
2 79944 1 3281
2 79945 1 3282
2 79946 1 3282
2 79947 1 3282
2 79948 1 3283
2 79949 1 3283
2 79950 1 3288
2 79951 1 3288
2 79952 1 3288
2 79953 1 3289
2 79954 1 3289
2 79955 1 3289
2 79956 1 3297
2 79957 1 3297
2 79958 1 3297
2 79959 1 3298
2 79960 1 3298
2 79961 1 3299
2 79962 1 3299
2 79963 1 3303
2 79964 1 3303
2 79965 1 3303
2 79966 1 3303
2 79967 1 3306
2 79968 1 3306
2 79969 1 3326
2 79970 1 3326
2 79971 1 3327
2 79972 1 3327
2 79973 1 3327
2 79974 1 3327
2 79975 1 3327
2 79976 1 3333
2 79977 1 3333
2 79978 1 3333
2 79979 1 3333
2 79980 1 3333
2 79981 1 3333
2 79982 1 3334
2 79983 1 3334
2 79984 1 3334
2 79985 1 3334
2 79986 1 3334
2 79987 1 3334
2 79988 1 3334
2 79989 1 3334
2 79990 1 3334
2 79991 1 3338
2 79992 1 3338
2 79993 1 3339
2 79994 1 3339
2 79995 1 3339
2 79996 1 3340
2 79997 1 3340
2 79998 1 3340
2 79999 1 3340
2 80000 1 3340
2 80001 1 3344
2 80002 1 3344
2 80003 1 3344
2 80004 1 3344
2 80005 1 3344
2 80006 1 3344
2 80007 1 3344
2 80008 1 3344
2 80009 1 3345
2 80010 1 3345
2 80011 1 3345
2 80012 1 3359
2 80013 1 3359
2 80014 1 3359
2 80015 1 3359
2 80016 1 3359
2 80017 1 3359
2 80018 1 3359
2 80019 1 3359
2 80020 1 3359
2 80021 1 3359
2 80022 1 3359
2 80023 1 3359
2 80024 1 3359
2 80025 1 3359
2 80026 1 3359
2 80027 1 3359
2 80028 1 3359
2 80029 1 3359
2 80030 1 3359
2 80031 1 3359
2 80032 1 3359
2 80033 1 3359
2 80034 1 3359
2 80035 1 3359
2 80036 1 3359
2 80037 1 3359
2 80038 1 3359
2 80039 1 3359
2 80040 1 3359
2 80041 1 3359
2 80042 1 3359
2 80043 1 3359
2 80044 1 3359
2 80045 1 3359
2 80046 1 3359
2 80047 1 3360
2 80048 1 3360
2 80049 1 3360
2 80050 1 3360
2 80051 1 3360
2 80052 1 3360
2 80053 1 3360
2 80054 1 3361
2 80055 1 3361
2 80056 1 3361
2 80057 1 3362
2 80058 1 3362
2 80059 1 3370
2 80060 1 3370
2 80061 1 3370
2 80062 1 3371
2 80063 1 3371
2 80064 1 3373
2 80065 1 3373
2 80066 1 3375
2 80067 1 3375
2 80068 1 3375
2 80069 1 3375
2 80070 1 3375
2 80071 1 3376
2 80072 1 3376
2 80073 1 3376
2 80074 1 3376
2 80075 1 3376
2 80076 1 3377
2 80077 1 3377
2 80078 1 3377
2 80079 1 3377
2 80080 1 3377
2 80081 1 3377
2 80082 1 3378
2 80083 1 3378
2 80084 1 3379
2 80085 1 3379
2 80086 1 3379
2 80087 1 3379
2 80088 1 3381
2 80089 1 3381
2 80090 1 3382
2 80091 1 3382
2 80092 1 3382
2 80093 1 3386
2 80094 1 3386
2 80095 1 3386
2 80096 1 3386
2 80097 1 3399
2 80098 1 3399
2 80099 1 3400
2 80100 1 3400
2 80101 1 3400
2 80102 1 3400
2 80103 1 3401
2 80104 1 3401
2 80105 1 3401
2 80106 1 3401
2 80107 1 3401
2 80108 1 3401
2 80109 1 3401
2 80110 1 3401
2 80111 1 3401
2 80112 1 3401
2 80113 1 3401
2 80114 1 3401
2 80115 1 3401
2 80116 1 3401
2 80117 1 3401
2 80118 1 3401
2 80119 1 3401
2 80120 1 3402
2 80121 1 3402
2 80122 1 3415
2 80123 1 3415
2 80124 1 3415
2 80125 1 3415
2 80126 1 3415
2 80127 1 3415
2 80128 1 3415
2 80129 1 3415
2 80130 1 3416
2 80131 1 3416
2 80132 1 3417
2 80133 1 3417
2 80134 1 3420
2 80135 1 3420
2 80136 1 3421
2 80137 1 3421
2 80138 1 3421
2 80139 1 3423
2 80140 1 3423
2 80141 1 3427
2 80142 1 3427
2 80143 1 3440
2 80144 1 3440
2 80145 1 3440
2 80146 1 3440
2 80147 1 3440
2 80148 1 3440
2 80149 1 3452
2 80150 1 3452
2 80151 1 3452
2 80152 1 3452
2 80153 1 3452
2 80154 1 3452
2 80155 1 3452
2 80156 1 3454
2 80157 1 3454
2 80158 1 3454
2 80159 1 3459
2 80160 1 3459
2 80161 1 3459
2 80162 1 3459
2 80163 1 3459
2 80164 1 3459
2 80165 1 3459
2 80166 1 3459
2 80167 1 3459
2 80168 1 3459
2 80169 1 3459
2 80170 1 3459
2 80171 1 3459
2 80172 1 3459
2 80173 1 3459
2 80174 1 3459
2 80175 1 3459
2 80176 1 3459
2 80177 1 3461
2 80178 1 3461
2 80179 1 3461
2 80180 1 3461
2 80181 1 3461
2 80182 1 3462
2 80183 1 3462
2 80184 1 3462
2 80185 1 3462
2 80186 1 3464
2 80187 1 3464
2 80188 1 3464
2 80189 1 3464
2 80190 1 3464
2 80191 1 3464
2 80192 1 3464
2 80193 1 3464
2 80194 1 3464
2 80195 1 3465
2 80196 1 3465
2 80197 1 3465
2 80198 1 3465
2 80199 1 3465
2 80200 1 3486
2 80201 1 3486
2 80202 1 3498
2 80203 1 3498
2 80204 1 3498
2 80205 1 3498
2 80206 1 3499
2 80207 1 3499
2 80208 1 3499
2 80209 1 3499
2 80210 1 3500
2 80211 1 3500
2 80212 1 3501
2 80213 1 3501
2 80214 1 3519
2 80215 1 3519
2 80216 1 3519
2 80217 1 3520
2 80218 1 3520
2 80219 1 3520
2 80220 1 3520
2 80221 1 3521
2 80222 1 3521
2 80223 1 3521
2 80224 1 3521
2 80225 1 3522
2 80226 1 3522
2 80227 1 3522
2 80228 1 3522
2 80229 1 3529
2 80230 1 3529
2 80231 1 3530
2 80232 1 3530
2 80233 1 3531
2 80234 1 3531
2 80235 1 3534
2 80236 1 3534
2 80237 1 3535
2 80238 1 3535
2 80239 1 3536
2 80240 1 3536
2 80241 1 3536
2 80242 1 3543
2 80243 1 3543
2 80244 1 3543
2 80245 1 3543
2 80246 1 3543
2 80247 1 3543
2 80248 1 3547
2 80249 1 3547
2 80250 1 3548
2 80251 1 3548
2 80252 1 3548
2 80253 1 3550
2 80254 1 3550
2 80255 1 3551
2 80256 1 3551
2 80257 1 3551
2 80258 1 3551
2 80259 1 3551
2 80260 1 3551
2 80261 1 3551
2 80262 1 3551
2 80263 1 3551
2 80264 1 3552
2 80265 1 3552
2 80266 1 3552
2 80267 1 3567
2 80268 1 3567
2 80269 1 3567
2 80270 1 3568
2 80271 1 3568
2 80272 1 3568
2 80273 1 3568
2 80274 1 3568
2 80275 1 3568
2 80276 1 3568
2 80277 1 3568
2 80278 1 3568
2 80279 1 3568
2 80280 1 3568
2 80281 1 3568
2 80282 1 3568
2 80283 1 3568
2 80284 1 3568
2 80285 1 3568
2 80286 1 3568
2 80287 1 3568
2 80288 1 3568
2 80289 1 3568
2 80290 1 3568
2 80291 1 3568
2 80292 1 3569
2 80293 1 3569
2 80294 1 3570
2 80295 1 3570
2 80296 1 3570
2 80297 1 3570
2 80298 1 3570
2 80299 1 3570
2 80300 1 3571
2 80301 1 3571
2 80302 1 3571
2 80303 1 3571
2 80304 1 3571
2 80305 1 3571
2 80306 1 3573
2 80307 1 3573
2 80308 1 3573
2 80309 1 3573
2 80310 1 3573
2 80311 1 3575
2 80312 1 3575
2 80313 1 3575
2 80314 1 3575
2 80315 1 3575
2 80316 1 3575
2 80317 1 3583
2 80318 1 3583
2 80319 1 3583
2 80320 1 3583
2 80321 1 3583
2 80322 1 3583
2 80323 1 3584
2 80324 1 3584
2 80325 1 3585
2 80326 1 3585
2 80327 1 3597
2 80328 1 3597
2 80329 1 3618
2 80330 1 3618
2 80331 1 3618
2 80332 1 3618
2 80333 1 3618
2 80334 1 3618
2 80335 1 3618
2 80336 1 3618
2 80337 1 3618
2 80338 1 3618
2 80339 1 3618
2 80340 1 3618
2 80341 1 3618
2 80342 1 3618
2 80343 1 3619
2 80344 1 3619
2 80345 1 3619
2 80346 1 3619
2 80347 1 3619
2 80348 1 3620
2 80349 1 3620
2 80350 1 3620
2 80351 1 3620
2 80352 1 3620
2 80353 1 3620
2 80354 1 3620
2 80355 1 3620
2 80356 1 3620
2 80357 1 3620
2 80358 1 3620
2 80359 1 3620
2 80360 1 3620
2 80361 1 3620
2 80362 1 3620
2 80363 1 3620
2 80364 1 3620
2 80365 1 3620
2 80366 1 3621
2 80367 1 3621
2 80368 1 3621
2 80369 1 3621
2 80370 1 3621
2 80371 1 3621
2 80372 1 3621
2 80373 1 3622
2 80374 1 3622
2 80375 1 3622
2 80376 1 3622
2 80377 1 3622
2 80378 1 3622
2 80379 1 3623
2 80380 1 3623
2 80381 1 3623
2 80382 1 3623
2 80383 1 3623
2 80384 1 3623
2 80385 1 3623
2 80386 1 3623
2 80387 1 3623
2 80388 1 3623
2 80389 1 3623
2 80390 1 3623
2 80391 1 3623
2 80392 1 3623
2 80393 1 3623
2 80394 1 3623
2 80395 1 3623
2 80396 1 3623
2 80397 1 3623
2 80398 1 3623
2 80399 1 3623
2 80400 1 3623
2 80401 1 3623
2 80402 1 3623
2 80403 1 3623
2 80404 1 3623
2 80405 1 3623
2 80406 1 3623
2 80407 1 3623
2 80408 1 3623
2 80409 1 3623
2 80410 1 3623
2 80411 1 3623
2 80412 1 3623
2 80413 1 3623
2 80414 1 3623
2 80415 1 3623
2 80416 1 3623
2 80417 1 3623
2 80418 1 3623
2 80419 1 3623
2 80420 1 3623
2 80421 1 3623
2 80422 1 3623
2 80423 1 3623
2 80424 1 3623
2 80425 1 3623
2 80426 1 3623
2 80427 1 3624
2 80428 1 3624
2 80429 1 3624
2 80430 1 3625
2 80431 1 3625
2 80432 1 3625
2 80433 1 3626
2 80434 1 3626
2 80435 1 3626
2 80436 1 3628
2 80437 1 3628
2 80438 1 3633
2 80439 1 3633
2 80440 1 3634
2 80441 1 3634
2 80442 1 3634
2 80443 1 3640
2 80444 1 3640
2 80445 1 3640
2 80446 1 3640
2 80447 1 3642
2 80448 1 3642
2 80449 1 3642
2 80450 1 3647
2 80451 1 3647
2 80452 1 3652
2 80453 1 3652
2 80454 1 3652
2 80455 1 3652
2 80456 1 3652
2 80457 1 3652
2 80458 1 3652
2 80459 1 3652
2 80460 1 3652
2 80461 1 3652
2 80462 1 3653
2 80463 1 3653
2 80464 1 3654
2 80465 1 3654
2 80466 1 3654
2 80467 1 3654
2 80468 1 3654
2 80469 1 3654
2 80470 1 3654
2 80471 1 3658
2 80472 1 3658
2 80473 1 3664
2 80474 1 3664
2 80475 1 3672
2 80476 1 3672
2 80477 1 3672
2 80478 1 3672
2 80479 1 3672
2 80480 1 3672
2 80481 1 3673
2 80482 1 3673
2 80483 1 3673
2 80484 1 3673
2 80485 1 3673
2 80486 1 3682
2 80487 1 3682
2 80488 1 3682
2 80489 1 3682
2 80490 1 3682
2 80491 1 3682
2 80492 1 3682
2 80493 1 3682
2 80494 1 3682
2 80495 1 3682
2 80496 1 3683
2 80497 1 3683
2 80498 1 3683
2 80499 1 3691
2 80500 1 3691
2 80501 1 3692
2 80502 1 3692
2 80503 1 3695
2 80504 1 3695
2 80505 1 3695
2 80506 1 3695
2 80507 1 3705
2 80508 1 3705
2 80509 1 3705
2 80510 1 3705
2 80511 1 3705
2 80512 1 3705
2 80513 1 3705
2 80514 1 3705
2 80515 1 3705
2 80516 1 3705
2 80517 1 3705
2 80518 1 3705
2 80519 1 3705
2 80520 1 3706
2 80521 1 3706
2 80522 1 3706
2 80523 1 3706
2 80524 1 3706
2 80525 1 3707
2 80526 1 3707
2 80527 1 3707
2 80528 1 3707
2 80529 1 3707
2 80530 1 3707
2 80531 1 3707
2 80532 1 3707
2 80533 1 3707
2 80534 1 3707
2 80535 1 3707
2 80536 1 3707
2 80537 1 3707
2 80538 1 3707
2 80539 1 3707
2 80540 1 3707
2 80541 1 3707
2 80542 1 3707
2 80543 1 3707
2 80544 1 3707
2 80545 1 3707
2 80546 1 3708
2 80547 1 3708
2 80548 1 3708
2 80549 1 3708
2 80550 1 3708
2 80551 1 3708
2 80552 1 3708
2 80553 1 3708
2 80554 1 3717
2 80555 1 3717
2 80556 1 3717
2 80557 1 3717
2 80558 1 3717
2 80559 1 3717
2 80560 1 3717
2 80561 1 3717
2 80562 1 3717
2 80563 1 3717
2 80564 1 3717
2 80565 1 3717
2 80566 1 3717
2 80567 1 3718
2 80568 1 3718
2 80569 1 3718
2 80570 1 3718
2 80571 1 3721
2 80572 1 3721
2 80573 1 3721
2 80574 1 3723
2 80575 1 3723
2 80576 1 3723
2 80577 1 3723
2 80578 1 3723
2 80579 1 3724
2 80580 1 3724
2 80581 1 3724
2 80582 1 3725
2 80583 1 3725
2 80584 1 3725
2 80585 1 3725
2 80586 1 3725
2 80587 1 3725
2 80588 1 3725
2 80589 1 3726
2 80590 1 3726
2 80591 1 3726
2 80592 1 3726
2 80593 1 3727
2 80594 1 3727
2 80595 1 3727
2 80596 1 3732
2 80597 1 3732
2 80598 1 3732
2 80599 1 3732
2 80600 1 3733
2 80601 1 3733
2 80602 1 3733
2 80603 1 3733
2 80604 1 3733
2 80605 1 3733
2 80606 1 3733
2 80607 1 3733
2 80608 1 3733
2 80609 1 3733
2 80610 1 3733
2 80611 1 3734
2 80612 1 3734
2 80613 1 3734
2 80614 1 3734
2 80615 1 3734
2 80616 1 3741
2 80617 1 3741
2 80618 1 3741
2 80619 1 3741
2 80620 1 3741
2 80621 1 3741
2 80622 1 3741
2 80623 1 3741
2 80624 1 3741
2 80625 1 3741
2 80626 1 3741
2 80627 1 3741
2 80628 1 3742
2 80629 1 3742
2 80630 1 3744
2 80631 1 3744
2 80632 1 3744
2 80633 1 3745
2 80634 1 3745
2 80635 1 3745
2 80636 1 3745
2 80637 1 3745
2 80638 1 3745
2 80639 1 3746
2 80640 1 3746
2 80641 1 3746
2 80642 1 3746
2 80643 1 3746
2 80644 1 3759
2 80645 1 3759
2 80646 1 3759
2 80647 1 3771
2 80648 1 3771
2 80649 1 3771
2 80650 1 3771
2 80651 1 3771
2 80652 1 3771
2 80653 1 3771
2 80654 1 3771
2 80655 1 3772
2 80656 1 3772
2 80657 1 3773
2 80658 1 3773
2 80659 1 3773
2 80660 1 3773
2 80661 1 3773
2 80662 1 3773
2 80663 1 3780
2 80664 1 3780
2 80665 1 3780
2 80666 1 3780
2 80667 1 3780
2 80668 1 3780
2 80669 1 3780
2 80670 1 3781
2 80671 1 3781
2 80672 1 3782
2 80673 1 3782
2 80674 1 3782
2 80675 1 3790
2 80676 1 3790
2 80677 1 3805
2 80678 1 3805
2 80679 1 3805
2 80680 1 3805
2 80681 1 3805
2 80682 1 3805
2 80683 1 3805
2 80684 1 3805
2 80685 1 3805
2 80686 1 3805
2 80687 1 3805
2 80688 1 3805
2 80689 1 3805
2 80690 1 3805
2 80691 1 3805
2 80692 1 3805
2 80693 1 3805
2 80694 1 3806
2 80695 1 3806
2 80696 1 3806
2 80697 1 3815
2 80698 1 3815
2 80699 1 3815
2 80700 1 3815
2 80701 1 3820
2 80702 1 3820
2 80703 1 3820
2 80704 1 3820
2 80705 1 3820
2 80706 1 3822
2 80707 1 3822
2 80708 1 3822
2 80709 1 3825
2 80710 1 3825
2 80711 1 3825
2 80712 1 3825
2 80713 1 3825
2 80714 1 3825
2 80715 1 3825
2 80716 1 3825
2 80717 1 3825
2 80718 1 3833
2 80719 1 3833
2 80720 1 3833
2 80721 1 3833
2 80722 1 3833
2 80723 1 3833
2 80724 1 3833
2 80725 1 3833
2 80726 1 3833
2 80727 1 3833
2 80728 1 3833
2 80729 1 3833
2 80730 1 3833
2 80731 1 3833
2 80732 1 3833
2 80733 1 3833
2 80734 1 3833
2 80735 1 3833
2 80736 1 3833
2 80737 1 3833
2 80738 1 3833
2 80739 1 3833
2 80740 1 3833
2 80741 1 3834
2 80742 1 3834
2 80743 1 3834
2 80744 1 3834
2 80745 1 3834
2 80746 1 3835
2 80747 1 3835
2 80748 1 3835
2 80749 1 3835
2 80750 1 3835
2 80751 1 3835
2 80752 1 3835
2 80753 1 3835
2 80754 1 3835
2 80755 1 3835
2 80756 1 3835
2 80757 1 3835
2 80758 1 3844
2 80759 1 3844
2 80760 1 3844
2 80761 1 3844
2 80762 1 3844
2 80763 1 3844
2 80764 1 3845
2 80765 1 3845
2 80766 1 3846
2 80767 1 3846
2 80768 1 3847
2 80769 1 3847
2 80770 1 3848
2 80771 1 3848
2 80772 1 3848
2 80773 1 3850
2 80774 1 3850
2 80775 1 3850
2 80776 1 3850
2 80777 1 3850
2 80778 1 3850
2 80779 1 3850
2 80780 1 3851
2 80781 1 3851
2 80782 1 3851
2 80783 1 3851
2 80784 1 3851
2 80785 1 3851
2 80786 1 3851
2 80787 1 3852
2 80788 1 3852
2 80789 1 3852
2 80790 1 3852
2 80791 1 3858
2 80792 1 3858
2 80793 1 3858
2 80794 1 3858
2 80795 1 3860
2 80796 1 3860
2 80797 1 3860
2 80798 1 3860
2 80799 1 3863
2 80800 1 3863
2 80801 1 3863
2 80802 1 3864
2 80803 1 3864
2 80804 1 3864
2 80805 1 3864
2 80806 1 3864
2 80807 1 3864
2 80808 1 3864
2 80809 1 3864
2 80810 1 3864
2 80811 1 3864
2 80812 1 3864
2 80813 1 3864
2 80814 1 3864
2 80815 1 3864
2 80816 1 3864
2 80817 1 3864
2 80818 1 3864
2 80819 1 3864
2 80820 1 3864
2 80821 1 3864
2 80822 1 3866
2 80823 1 3866
2 80824 1 3866
2 80825 1 3881
2 80826 1 3881
2 80827 1 3881
2 80828 1 3881
2 80829 1 3881
2 80830 1 3882
2 80831 1 3882
2 80832 1 3882
2 80833 1 3882
2 80834 1 3882
2 80835 1 3882
2 80836 1 3882
2 80837 1 3882
2 80838 1 3882
2 80839 1 3882
2 80840 1 3882
2 80841 1 3882
2 80842 1 3882
2 80843 1 3882
2 80844 1 3882
2 80845 1 3882
2 80846 1 3882
2 80847 1 3882
2 80848 1 3882
2 80849 1 3882
2 80850 1 3882
2 80851 1 3882
2 80852 1 3882
2 80853 1 3882
2 80854 1 3882
2 80855 1 3882
2 80856 1 3882
2 80857 1 3882
2 80858 1 3882
2 80859 1 3882
2 80860 1 3882
2 80861 1 3882
2 80862 1 3882
2 80863 1 3882
2 80864 1 3882
2 80865 1 3882
2 80866 1 3882
2 80867 1 3882
2 80868 1 3882
2 80869 1 3882
2 80870 1 3882
2 80871 1 3882
2 80872 1 3882
2 80873 1 3882
2 80874 1 3882
2 80875 1 3882
2 80876 1 3882
2 80877 1 3882
2 80878 1 3882
2 80879 1 3882
2 80880 1 3882
2 80881 1 3882
2 80882 1 3882
2 80883 1 3882
2 80884 1 3882
2 80885 1 3882
2 80886 1 3882
2 80887 1 3882
2 80888 1 3882
2 80889 1 3882
2 80890 1 3882
2 80891 1 3882
2 80892 1 3882
2 80893 1 3882
2 80894 1 3882
2 80895 1 3882
2 80896 1 3883
2 80897 1 3883
2 80898 1 3883
2 80899 1 3883
2 80900 1 3883
2 80901 1 3883
2 80902 1 3883
2 80903 1 3883
2 80904 1 3883
2 80905 1 3883
2 80906 1 3883
2 80907 1 3883
2 80908 1 3883
2 80909 1 3883
2 80910 1 3883
2 80911 1 3883
2 80912 1 3883
2 80913 1 3884
2 80914 1 3884
2 80915 1 3884
2 80916 1 3884
2 80917 1 3884
2 80918 1 3884
2 80919 1 3884
2 80920 1 3884
2 80921 1 3886
2 80922 1 3886
2 80923 1 3894
2 80924 1 3894
2 80925 1 3894
2 80926 1 3894
2 80927 1 3894
2 80928 1 3894
2 80929 1 3894
2 80930 1 3894
2 80931 1 3894
2 80932 1 3894
2 80933 1 3903
2 80934 1 3903
2 80935 1 3903
2 80936 1 3919
2 80937 1 3919
2 80938 1 3919
2 80939 1 3921
2 80940 1 3921
2 80941 1 3921
2 80942 1 3921
2 80943 1 3921
2 80944 1 3921
2 80945 1 3921
2 80946 1 3921
2 80947 1 3921
2 80948 1 3921
2 80949 1 3921
2 80950 1 3921
2 80951 1 3921
2 80952 1 3921
2 80953 1 3921
2 80954 1 3921
2 80955 1 3921
2 80956 1 3921
2 80957 1 3921
2 80958 1 3921
2 80959 1 3921
2 80960 1 3921
2 80961 1 3921
2 80962 1 3921
2 80963 1 3921
2 80964 1 3921
2 80965 1 3921
2 80966 1 3921
2 80967 1 3921
2 80968 1 3922
2 80969 1 3922
2 80970 1 3922
2 80971 1 3923
2 80972 1 3923
2 80973 1 3933
2 80974 1 3933
2 80975 1 3933
2 80976 1 3933
2 80977 1 3935
2 80978 1 3935
2 80979 1 3935
2 80980 1 3935
2 80981 1 3935
2 80982 1 3935
2 80983 1 3935
2 80984 1 3935
2 80985 1 3935
2 80986 1 3935
2 80987 1 3937
2 80988 1 3937
2 80989 1 3937
2 80990 1 3937
2 80991 1 3937
2 80992 1 3937
2 80993 1 3937
2 80994 1 3937
2 80995 1 3937
2 80996 1 3937
2 80997 1 3937
2 80998 1 3937
2 80999 1 3937
2 81000 1 3937
2 81001 1 3937
2 81002 1 3937
2 81003 1 3937
2 81004 1 3937
2 81005 1 3947
2 81006 1 3947
2 81007 1 3947
2 81008 1 3947
2 81009 1 3947
2 81010 1 3947
2 81011 1 3947
2 81012 1 3947
2 81013 1 3947
2 81014 1 3947
2 81015 1 3947
2 81016 1 3947
2 81017 1 3947
2 81018 1 3947
2 81019 1 3947
2 81020 1 3947
2 81021 1 3947
2 81022 1 3947
2 81023 1 3947
2 81024 1 3947
2 81025 1 3947
2 81026 1 3947
2 81027 1 3947
2 81028 1 3947
2 81029 1 3947
2 81030 1 3947
2 81031 1 3947
2 81032 1 3948
2 81033 1 3948
2 81034 1 3948
2 81035 1 3952
2 81036 1 3952
2 81037 1 3952
2 81038 1 3952
2 81039 1 3955
2 81040 1 3955
2 81041 1 3964
2 81042 1 3964
2 81043 1 3964
2 81044 1 3964
2 81045 1 3964
2 81046 1 3964
2 81047 1 3964
2 81048 1 3964
2 81049 1 3964
2 81050 1 3964
2 81051 1 3964
2 81052 1 3964
2 81053 1 3964
2 81054 1 3965
2 81055 1 3965
2 81056 1 3965
2 81057 1 3965
2 81058 1 3965
2 81059 1 3965
2 81060 1 3966
2 81061 1 3966
2 81062 1 3966
2 81063 1 3966
2 81064 1 3967
2 81065 1 3967
2 81066 1 3967
2 81067 1 3967
2 81068 1 3967
2 81069 1 3972
2 81070 1 3972
2 81071 1 3973
2 81072 1 3973
2 81073 1 3974
2 81074 1 3974
2 81075 1 3974
2 81076 1 3974
2 81077 1 3974
2 81078 1 3974
2 81079 1 3974
2 81080 1 3974
2 81081 1 3974
2 81082 1 3974
2 81083 1 3974
2 81084 1 3975
2 81085 1 3975
2 81086 1 3975
2 81087 1 3991
2 81088 1 3991
2 81089 1 3991
2 81090 1 3991
2 81091 1 3991
2 81092 1 3991
2 81093 1 3991
2 81094 1 3991
2 81095 1 3991
2 81096 1 3992
2 81097 1 3992
2 81098 1 3992
2 81099 1 3992
2 81100 1 3992
2 81101 1 3992
2 81102 1 3992
2 81103 1 3992
2 81104 1 3992
2 81105 1 3992
2 81106 1 3992
2 81107 1 3992
2 81108 1 3992
2 81109 1 3992
2 81110 1 3992
2 81111 1 3992
2 81112 1 3992
2 81113 1 3992
2 81114 1 3993
2 81115 1 3993
2 81116 1 3994
2 81117 1 3994
2 81118 1 3994
2 81119 1 3994
2 81120 1 3994
2 81121 1 3994
2 81122 1 3995
2 81123 1 3995
2 81124 1 3995
2 81125 1 3995
2 81126 1 3995
2 81127 1 3995
2 81128 1 3995
2 81129 1 3995
2 81130 1 3996
2 81131 1 3996
2 81132 1 4000
2 81133 1 4000
2 81134 1 4000
2 81135 1 4006
2 81136 1 4006
2 81137 1 4006
2 81138 1 4013
2 81139 1 4013
2 81140 1 4013
2 81141 1 4022
2 81142 1 4022
2 81143 1 4022
2 81144 1 4022
2 81145 1 4022
2 81146 1 4022
2 81147 1 4022
2 81148 1 4022
2 81149 1 4022
2 81150 1 4022
2 81151 1 4022
2 81152 1 4022
2 81153 1 4022
2 81154 1 4022
2 81155 1 4022
2 81156 1 4022
2 81157 1 4022
2 81158 1 4022
2 81159 1 4022
2 81160 1 4022
2 81161 1 4022
2 81162 1 4022
2 81163 1 4022
2 81164 1 4022
2 81165 1 4022
2 81166 1 4022
2 81167 1 4022
2 81168 1 4022
2 81169 1 4022
2 81170 1 4022
2 81171 1 4022
2 81172 1 4022
2 81173 1 4022
2 81174 1 4022
2 81175 1 4022
2 81176 1 4022
2 81177 1 4022
2 81178 1 4022
2 81179 1 4022
2 81180 1 4022
2 81181 1 4022
2 81182 1 4022
2 81183 1 4022
2 81184 1 4022
2 81185 1 4022
2 81186 1 4022
2 81187 1 4022
2 81188 1 4022
2 81189 1 4022
2 81190 1 4022
2 81191 1 4022
2 81192 1 4022
2 81193 1 4022
2 81194 1 4022
2 81195 1 4023
2 81196 1 4023
2 81197 1 4023
2 81198 1 4037
2 81199 1 4037
2 81200 1 4037
2 81201 1 4037
2 81202 1 4037
2 81203 1 4037
2 81204 1 4037
2 81205 1 4037
2 81206 1 4038
2 81207 1 4038
2 81208 1 4038
2 81209 1 4039
2 81210 1 4039
2 81211 1 4043
2 81212 1 4043
2 81213 1 4044
2 81214 1 4044
2 81215 1 4044
2 81216 1 4044
2 81217 1 4044
2 81218 1 4044
2 81219 1 4044
2 81220 1 4052
2 81221 1 4052
2 81222 1 4052
2 81223 1 4052
2 81224 1 4052
2 81225 1 4053
2 81226 1 4053
2 81227 1 4060
2 81228 1 4060
2 81229 1 4062
2 81230 1 4062
2 81231 1 4062
2 81232 1 4062
2 81233 1 4070
2 81234 1 4070
2 81235 1 4072
2 81236 1 4072
2 81237 1 4077
2 81238 1 4077
2 81239 1 4079
2 81240 1 4079
2 81241 1 4079
2 81242 1 4079
2 81243 1 4079
2 81244 1 4087
2 81245 1 4087
2 81246 1 4087
2 81247 1 4088
2 81248 1 4088
2 81249 1 4100
2 81250 1 4100
2 81251 1 4100
2 81252 1 4100
2 81253 1 4100
2 81254 1 4100
2 81255 1 4100
2 81256 1 4101
2 81257 1 4101
2 81258 1 4110
2 81259 1 4110
2 81260 1 4110
2 81261 1 4110
2 81262 1 4110
2 81263 1 4117
2 81264 1 4117
2 81265 1 4138
2 81266 1 4138
2 81267 1 4138
2 81268 1 4138
2 81269 1 4138
2 81270 1 4138
2 81271 1 4138
2 81272 1 4138
2 81273 1 4138
2 81274 1 4138
2 81275 1 4139
2 81276 1 4139
2 81277 1 4139
2 81278 1 4140
2 81279 1 4140
2 81280 1 4140
2 81281 1 4140
2 81282 1 4140
2 81283 1 4140
2 81284 1 4140
2 81285 1 4140
2 81286 1 4140
2 81287 1 4140
2 81288 1 4140
2 81289 1 4141
2 81290 1 4141
2 81291 1 4141
2 81292 1 4141
2 81293 1 4141
2 81294 1 4149
2 81295 1 4149
2 81296 1 4149
2 81297 1 4149
2 81298 1 4149
2 81299 1 4149
2 81300 1 4149
2 81301 1 4149
2 81302 1 4150
2 81303 1 4150
2 81304 1 4150
2 81305 1 4151
2 81306 1 4151
2 81307 1 4151
2 81308 1 4151
2 81309 1 4151
2 81310 1 4151
2 81311 1 4151
2 81312 1 4152
2 81313 1 4152
2 81314 1 4152
2 81315 1 4152
2 81316 1 4152
2 81317 1 4152
2 81318 1 4152
2 81319 1 4160
2 81320 1 4160
2 81321 1 4160
2 81322 1 4160
2 81323 1 4160
2 81324 1 4160
2 81325 1 4160
2 81326 1 4160
2 81327 1 4160
2 81328 1 4160
2 81329 1 4160
2 81330 1 4161
2 81331 1 4161
2 81332 1 4162
2 81333 1 4162
2 81334 1 4162
2 81335 1 4162
2 81336 1 4163
2 81337 1 4163
2 81338 1 4163
2 81339 1 4163
2 81340 1 4164
2 81341 1 4164
2 81342 1 4166
2 81343 1 4166
2 81344 1 4168
2 81345 1 4168
2 81346 1 4168
2 81347 1 4168
2 81348 1 4168
2 81349 1 4168
2 81350 1 4168
2 81351 1 4168
2 81352 1 4168
2 81353 1 4170
2 81354 1 4170
2 81355 1 4172
2 81356 1 4172
2 81357 1 4172
2 81358 1 4172
2 81359 1 4187
2 81360 1 4187
2 81361 1 4188
2 81362 1 4188
2 81363 1 4188
2 81364 1 4191
2 81365 1 4191
2 81366 1 4192
2 81367 1 4192
2 81368 1 4194
2 81369 1 4194
2 81370 1 4194
2 81371 1 4197
2 81372 1 4197
2 81373 1 4197
2 81374 1 4210
2 81375 1 4210
2 81376 1 4211
2 81377 1 4211
2 81378 1 4211
2 81379 1 4211
2 81380 1 4212
2 81381 1 4212
2 81382 1 4212
2 81383 1 4219
2 81384 1 4219
2 81385 1 4219
2 81386 1 4219
2 81387 1 4219
2 81388 1 4219
2 81389 1 4219
2 81390 1 4219
2 81391 1 4219
2 81392 1 4219
2 81393 1 4219
2 81394 1 4219
2 81395 1 4220
2 81396 1 4220
2 81397 1 4220
2 81398 1 4220
2 81399 1 4221
2 81400 1 4221
2 81401 1 4221
2 81402 1 4223
2 81403 1 4223
2 81404 1 4237
2 81405 1 4237
2 81406 1 4237
2 81407 1 4237
2 81408 1 4237
2 81409 1 4243
2 81410 1 4243
2 81411 1 4243
2 81412 1 4243
2 81413 1 4244
2 81414 1 4244
2 81415 1 4247
2 81416 1 4247
2 81417 1 4247
2 81418 1 4247
2 81419 1 4248
2 81420 1 4248
2 81421 1 4248
2 81422 1 4248
2 81423 1 4248
2 81424 1 4248
2 81425 1 4249
2 81426 1 4249
2 81427 1 4249
2 81428 1 4249
2 81429 1 4249
2 81430 1 4250
2 81431 1 4250
2 81432 1 4250
2 81433 1 4250
2 81434 1 4250
2 81435 1 4250
2 81436 1 4251
2 81437 1 4251
2 81438 1 4251
2 81439 1 4253
2 81440 1 4253
2 81441 1 4255
2 81442 1 4255
2 81443 1 4255
2 81444 1 4255
2 81445 1 4256
2 81446 1 4256
2 81447 1 4257
2 81448 1 4257
2 81449 1 4258
2 81450 1 4258
2 81451 1 4258
2 81452 1 4258
2 81453 1 4259
2 81454 1 4259
2 81455 1 4263
2 81456 1 4263
2 81457 1 4263
2 81458 1 4263
2 81459 1 4263
2 81460 1 4264
2 81461 1 4264
2 81462 1 4264
2 81463 1 4266
2 81464 1 4266
2 81465 1 4266
2 81466 1 4266
2 81467 1 4266
2 81468 1 4266
2 81469 1 4266
2 81470 1 4266
2 81471 1 4276
2 81472 1 4276
2 81473 1 4276
2 81474 1 4276
2 81475 1 4276
2 81476 1 4276
2 81477 1 4277
2 81478 1 4277
2 81479 1 4277
2 81480 1 4277
2 81481 1 4277
2 81482 1 4277
2 81483 1 4280
2 81484 1 4280
2 81485 1 4281
2 81486 1 4281
2 81487 1 4291
2 81488 1 4291
2 81489 1 4291
2 81490 1 4291
2 81491 1 4291
2 81492 1 4291
2 81493 1 4291
2 81494 1 4291
2 81495 1 4291
2 81496 1 4291
2 81497 1 4291
2 81498 1 4291
2 81499 1 4291
2 81500 1 4291
2 81501 1 4293
2 81502 1 4293
2 81503 1 4293
2 81504 1 4294
2 81505 1 4294
2 81506 1 4295
2 81507 1 4295
2 81508 1 4295
2 81509 1 4295
2 81510 1 4298
2 81511 1 4298
2 81512 1 4298
2 81513 1 4300
2 81514 1 4300
2 81515 1 4307
2 81516 1 4307
2 81517 1 4323
2 81518 1 4323
2 81519 1 4341
2 81520 1 4341
2 81521 1 4341
2 81522 1 4341
2 81523 1 4341
2 81524 1 4341
2 81525 1 4341
2 81526 1 4341
2 81527 1 4341
2 81528 1 4341
2 81529 1 4341
2 81530 1 4341
2 81531 1 4341
2 81532 1 4341
2 81533 1 4341
2 81534 1 4341
2 81535 1 4341
2 81536 1 4341
2 81537 1 4341
2 81538 1 4341
2 81539 1 4341
2 81540 1 4341
2 81541 1 4341
2 81542 1 4341
2 81543 1 4341
2 81544 1 4341
2 81545 1 4341
2 81546 1 4342
2 81547 1 4342
2 81548 1 4342
2 81549 1 4342
2 81550 1 4342
2 81551 1 4342
2 81552 1 4342
2 81553 1 4342
2 81554 1 4342
2 81555 1 4342
2 81556 1 4342
2 81557 1 4342
2 81558 1 4344
2 81559 1 4344
2 81560 1 4344
2 81561 1 4344
2 81562 1 4345
2 81563 1 4345
2 81564 1 4345
2 81565 1 4345
2 81566 1 4345
2 81567 1 4345
2 81568 1 4345
2 81569 1 4345
2 81570 1 4345
2 81571 1 4345
2 81572 1 4345
2 81573 1 4345
2 81574 1 4345
2 81575 1 4345
2 81576 1 4345
2 81577 1 4354
2 81578 1 4354
2 81579 1 4354
2 81580 1 4354
2 81581 1 4355
2 81582 1 4355
2 81583 1 4367
2 81584 1 4367
2 81585 1 4375
2 81586 1 4375
2 81587 1 4375
2 81588 1 4375
2 81589 1 4377
2 81590 1 4377
2 81591 1 4377
2 81592 1 4395
2 81593 1 4395
2 81594 1 4395
2 81595 1 4395
2 81596 1 4395
2 81597 1 4395
2 81598 1 4402
2 81599 1 4402
2 81600 1 4402
2 81601 1 4402
2 81602 1 4402
2 81603 1 4402
2 81604 1 4402
2 81605 1 4403
2 81606 1 4403
2 81607 1 4403
2 81608 1 4403
2 81609 1 4411
2 81610 1 4411
2 81611 1 4412
2 81612 1 4412
2 81613 1 4412
2 81614 1 4412
2 81615 1 4412
2 81616 1 4412
2 81617 1 4412
2 81618 1 4412
2 81619 1 4413
2 81620 1 4413
2 81621 1 4413
2 81622 1 4414
2 81623 1 4414
2 81624 1 4414
2 81625 1 4414
2 81626 1 4414
2 81627 1 4415
2 81628 1 4415
2 81629 1 4425
2 81630 1 4425
2 81631 1 4425
2 81632 1 4425
2 81633 1 4425
2 81634 1 4425
2 81635 1 4425
2 81636 1 4425
2 81637 1 4426
2 81638 1 4426
2 81639 1 4427
2 81640 1 4427
2 81641 1 4427
2 81642 1 4427
2 81643 1 4427
2 81644 1 4427
2 81645 1 4427
2 81646 1 4427
2 81647 1 4428
2 81648 1 4428
2 81649 1 4428
2 81650 1 4428
2 81651 1 4429
2 81652 1 4429
2 81653 1 4429
2 81654 1 4429
2 81655 1 4430
2 81656 1 4430
2 81657 1 4430
2 81658 1 4430
2 81659 1 4431
2 81660 1 4431
2 81661 1 4433
2 81662 1 4433
2 81663 1 4433
2 81664 1 4442
2 81665 1 4442
2 81666 1 4442
2 81667 1 4446
2 81668 1 4446
2 81669 1 4449
2 81670 1 4449
2 81671 1 4451
2 81672 1 4451
2 81673 1 4451
2 81674 1 4459
2 81675 1 4459
2 81676 1 4459
2 81677 1 4459
2 81678 1 4459
2 81679 1 4461
2 81680 1 4461
2 81681 1 4467
2 81682 1 4467
2 81683 1 4479
2 81684 1 4479
2 81685 1 4488
2 81686 1 4488
2 81687 1 4488
2 81688 1 4488
2 81689 1 4488
2 81690 1 4488
2 81691 1 4489
2 81692 1 4489
2 81693 1 4489
2 81694 1 4489
2 81695 1 4489
2 81696 1 4489
2 81697 1 4489
2 81698 1 4489
2 81699 1 4489
2 81700 1 4489
2 81701 1 4489
2 81702 1 4489
2 81703 1 4489
2 81704 1 4489
2 81705 1 4489
2 81706 1 4489
2 81707 1 4501
2 81708 1 4501
2 81709 1 4503
2 81710 1 4503
2 81711 1 4503
2 81712 1 4504
2 81713 1 4504
2 81714 1 4509
2 81715 1 4509
2 81716 1 4511
2 81717 1 4511
2 81718 1 4518
2 81719 1 4518
2 81720 1 4535
2 81721 1 4535
2 81722 1 4535
2 81723 1 4538
2 81724 1 4538
2 81725 1 4538
2 81726 1 4538
2 81727 1 4538
2 81728 1 4538
2 81729 1 4538
2 81730 1 4539
2 81731 1 4539
2 81732 1 4539
2 81733 1 4539
2 81734 1 4539
2 81735 1 4540
2 81736 1 4540
2 81737 1 4540
2 81738 1 4540
2 81739 1 4540
2 81740 1 4540
2 81741 1 4540
2 81742 1 4540
2 81743 1 4540
2 81744 1 4542
2 81745 1 4542
2 81746 1 4557
2 81747 1 4557
2 81748 1 4557
2 81749 1 4557
2 81750 1 4557
2 81751 1 4557
2 81752 1 4557
2 81753 1 4557
2 81754 1 4557
2 81755 1 4557
2 81756 1 4557
2 81757 1 4557
2 81758 1 4557
2 81759 1 4557
2 81760 1 4557
2 81761 1 4557
2 81762 1 4557
2 81763 1 4563
2 81764 1 4563
2 81765 1 4563
2 81766 1 4563
2 81767 1 4563
2 81768 1 4563
2 81769 1 4563
2 81770 1 4563
2 81771 1 4563
2 81772 1 4563
2 81773 1 4563
2 81774 1 4563
2 81775 1 4563
2 81776 1 4563
2 81777 1 4563
2 81778 1 4563
2 81779 1 4563
2 81780 1 4563
2 81781 1 4565
2 81782 1 4565
2 81783 1 4565
2 81784 1 4566
2 81785 1 4566
2 81786 1 4566
2 81787 1 4566
2 81788 1 4571
2 81789 1 4571
2 81790 1 4571
2 81791 1 4571
2 81792 1 4571
2 81793 1 4571
2 81794 1 4571
2 81795 1 4571
2 81796 1 4571
2 81797 1 4571
2 81798 1 4572
2 81799 1 4572
2 81800 1 4572
2 81801 1 4581
2 81802 1 4581
2 81803 1 4581
2 81804 1 4600
2 81805 1 4600
2 81806 1 4600
2 81807 1 4600
2 81808 1 4600
2 81809 1 4600
2 81810 1 4600
2 81811 1 4600
2 81812 1 4600
2 81813 1 4600
2 81814 1 4600
2 81815 1 4601
2 81816 1 4601
2 81817 1 4602
2 81818 1 4602
2 81819 1 4602
2 81820 1 4602
2 81821 1 4602
2 81822 1 4603
2 81823 1 4603
2 81824 1 4603
2 81825 1 4603
2 81826 1 4625
2 81827 1 4625
2 81828 1 4625
2 81829 1 4625
2 81830 1 4626
2 81831 1 4626
2 81832 1 4626
2 81833 1 4626
2 81834 1 4626
2 81835 1 4626
2 81836 1 4626
2 81837 1 4626
2 81838 1 4626
2 81839 1 4637
2 81840 1 4637
2 81841 1 4637
2 81842 1 4637
2 81843 1 4638
2 81844 1 4638
2 81845 1 4638
2 81846 1 4638
2 81847 1 4638
2 81848 1 4640
2 81849 1 4640
2 81850 1 4650
2 81851 1 4650
2 81852 1 4650
2 81853 1 4650
2 81854 1 4658
2 81855 1 4658
2 81856 1 4659
2 81857 1 4659
2 81858 1 4659
2 81859 1 4675
2 81860 1 4675
2 81861 1 4675
2 81862 1 4676
2 81863 1 4676
2 81864 1 4676
2 81865 1 4676
2 81866 1 4676
2 81867 1 4676
2 81868 1 4676
2 81869 1 4676
2 81870 1 4676
2 81871 1 4689
2 81872 1 4689
2 81873 1 4690
2 81874 1 4690
2 81875 1 4690
2 81876 1 4690
2 81877 1 4691
2 81878 1 4691
2 81879 1 4699
2 81880 1 4699
2 81881 1 4699
2 81882 1 4700
2 81883 1 4700
2 81884 1 4700
2 81885 1 4700
2 81886 1 4701
2 81887 1 4701
2 81888 1 4701
2 81889 1 4701
2 81890 1 4701
2 81891 1 4701
2 81892 1 4701
2 81893 1 4701
2 81894 1 4701
2 81895 1 4705
2 81896 1 4705
2 81897 1 4708
2 81898 1 4708
2 81899 1 4708
2 81900 1 4708
2 81901 1 4709
2 81902 1 4709
2 81903 1 4709
2 81904 1 4709
2 81905 1 4717
2 81906 1 4717
2 81907 1 4717
2 81908 1 4717
2 81909 1 4717
2 81910 1 4717
2 81911 1 4717
2 81912 1 4729
2 81913 1 4729
2 81914 1 4729
2 81915 1 4729
2 81916 1 4729
2 81917 1 4729
2 81918 1 4758
2 81919 1 4758
2 81920 1 4758
2 81921 1 4758
2 81922 1 4759
2 81923 1 4759
2 81924 1 4767
2 81925 1 4767
2 81926 1 4769
2 81927 1 4769
2 81928 1 4769
2 81929 1 4776
2 81930 1 4776
2 81931 1 4776
2 81932 1 4777
2 81933 1 4777
2 81934 1 4777
2 81935 1 4777
2 81936 1 4777
2 81937 1 4782
2 81938 1 4782
2 81939 1 4783
2 81940 1 4783
2 81941 1 4794
2 81942 1 4794
2 81943 1 4805
2 81944 1 4805
2 81945 1 4805
2 81946 1 4813
2 81947 1 4813
2 81948 1 4813
2 81949 1 4813
2 81950 1 4813
2 81951 1 4813
2 81952 1 4813
2 81953 1 4814
2 81954 1 4814
2 81955 1 4822
2 81956 1 4822
2 81957 1 4823
2 81958 1 4823
2 81959 1 4836
2 81960 1 4836
2 81961 1 4836
2 81962 1 4836
2 81963 1 4836
2 81964 1 4839
2 81965 1 4839
2 81966 1 4839
2 81967 1 4839
2 81968 1 4839
2 81969 1 4839
2 81970 1 4839
2 81971 1 4839
2 81972 1 4841
2 81973 1 4841
2 81974 1 4841
2 81975 1 4842
2 81976 1 4842
2 81977 1 4842
2 81978 1 4842
2 81979 1 4842
2 81980 1 4842
2 81981 1 4842
2 81982 1 4842
2 81983 1 4856
2 81984 1 4856
2 81985 1 4856
2 81986 1 4856
2 81987 1 4856
2 81988 1 4856
2 81989 1 4856
2 81990 1 4856
2 81991 1 4856
2 81992 1 4856
2 81993 1 4856
2 81994 1 4856
2 81995 1 4856
2 81996 1 4856
2 81997 1 4856
2 81998 1 4856
2 81999 1 4856
2 82000 1 4856
2 82001 1 4856
2 82002 1 4856
2 82003 1 4856
2 82004 1 4856
2 82005 1 4856
2 82006 1 4856
2 82007 1 4860
2 82008 1 4860
2 82009 1 4860
2 82010 1 4860
2 82011 1 4860
2 82012 1 4860
2 82013 1 4864
2 82014 1 4864
2 82015 1 4864
2 82016 1 4865
2 82017 1 4865
2 82018 1 4865
2 82019 1 4866
2 82020 1 4866
2 82021 1 4866
2 82022 1 4866
2 82023 1 4866
2 82024 1 4867
2 82025 1 4867
2 82026 1 4869
2 82027 1 4869
2 82028 1 4869
2 82029 1 4869
2 82030 1 4869
2 82031 1 4870
2 82032 1 4870
2 82033 1 4870
2 82034 1 4870
2 82035 1 4874
2 82036 1 4874
2 82037 1 4874
2 82038 1 4876
2 82039 1 4876
2 82040 1 4876
2 82041 1 4876
2 82042 1 4877
2 82043 1 4877
2 82044 1 4897
2 82045 1 4897
2 82046 1 4897
2 82047 1 4897
2 82048 1 4908
2 82049 1 4908
2 82050 1 4908
2 82051 1 4908
2 82052 1 4909
2 82053 1 4909
2 82054 1 4914
2 82055 1 4914
2 82056 1 4914
2 82057 1 4914
2 82058 1 4918
2 82059 1 4918
2 82060 1 4918
2 82061 1 4918
2 82062 1 4918
2 82063 1 4918
2 82064 1 4918
2 82065 1 4930
2 82066 1 4930
2 82067 1 4930
2 82068 1 4930
2 82069 1 4931
2 82070 1 4931
2 82071 1 4933
2 82072 1 4933
2 82073 1 4938
2 82074 1 4938
2 82075 1 4938
2 82076 1 4939
2 82077 1 4939
2 82078 1 4939
2 82079 1 4939
2 82080 1 4939
2 82081 1 4940
2 82082 1 4940
2 82083 1 4941
2 82084 1 4941
2 82085 1 4941
2 82086 1 4944
2 82087 1 4944
2 82088 1 4944
2 82089 1 4964
2 82090 1 4964
2 82091 1 4964
2 82092 1 4975
2 82093 1 4975
2 82094 1 4979
2 82095 1 4979
2 82096 1 4980
2 82097 1 4980
2 82098 1 4980
2 82099 1 4980
2 82100 1 5013
2 82101 1 5013
2 82102 1 5028
2 82103 1 5028
2 82104 1 5028
2 82105 1 5028
2 82106 1 5028
2 82107 1 5028
2 82108 1 5028
2 82109 1 5028
2 82110 1 5028
2 82111 1 5028
2 82112 1 5028
2 82113 1 5028
2 82114 1 5030
2 82115 1 5030
2 82116 1 5030
2 82117 1 5030
2 82118 1 5030
2 82119 1 5030
2 82120 1 5030
2 82121 1 5030
2 82122 1 5031
2 82123 1 5031
2 82124 1 5042
2 82125 1 5042
2 82126 1 5060
2 82127 1 5060
2 82128 1 5069
2 82129 1 5069
2 82130 1 5069
2 82131 1 5069
2 82132 1 5069
2 82133 1 5069
2 82134 1 5069
2 82135 1 5071
2 82136 1 5071
2 82137 1 5071
2 82138 1 5071
2 82139 1 5071
2 82140 1 5071
2 82141 1 5072
2 82142 1 5072
2 82143 1 5072
2 82144 1 5072
2 82145 1 5072
2 82146 1 5075
2 82147 1 5075
2 82148 1 5075
2 82149 1 5075
2 82150 1 5075
2 82151 1 5075
2 82152 1 5075
2 82153 1 5081
2 82154 1 5081
2 82155 1 5092
2 82156 1 5092
2 82157 1 5092
2 82158 1 5095
2 82159 1 5095
2 82160 1 5095
2 82161 1 5096
2 82162 1 5096
2 82163 1 5096
2 82164 1 5105
2 82165 1 5105
2 82166 1 5105
2 82167 1 5105
2 82168 1 5105
2 82169 1 5105
2 82170 1 5105
2 82171 1 5105
2 82172 1 5105
2 82173 1 5105
2 82174 1 5105
2 82175 1 5105
2 82176 1 5105
2 82177 1 5105
2 82178 1 5105
2 82179 1 5105
2 82180 1 5105
2 82181 1 5105
2 82182 1 5105
2 82183 1 5105
2 82184 1 5105
2 82185 1 5105
2 82186 1 5105
2 82187 1 5105
2 82188 1 5105
2 82189 1 5106
2 82190 1 5106
2 82191 1 5106
2 82192 1 5107
2 82193 1 5107
2 82194 1 5107
2 82195 1 5107
2 82196 1 5107
2 82197 1 5107
2 82198 1 5107
2 82199 1 5118
2 82200 1 5118
2 82201 1 5118
2 82202 1 5119
2 82203 1 5119
2 82204 1 5123
2 82205 1 5123
2 82206 1 5123
2 82207 1 5124
2 82208 1 5124
2 82209 1 5125
2 82210 1 5125
2 82211 1 5125
2 82212 1 5125
2 82213 1 5136
2 82214 1 5136
2 82215 1 5140
2 82216 1 5140
2 82217 1 5140
2 82218 1 5154
2 82219 1 5154
2 82220 1 5156
2 82221 1 5156
2 82222 1 5168
2 82223 1 5168
2 82224 1 5168
2 82225 1 5168
2 82226 1 5168
2 82227 1 5169
2 82228 1 5169
2 82229 1 5182
2 82230 1 5182
2 82231 1 5182
2 82232 1 5182
2 82233 1 5182
2 82234 1 5182
2 82235 1 5182
2 82236 1 5182
2 82237 1 5182
2 82238 1 5183
2 82239 1 5183
2 82240 1 5190
2 82241 1 5190
2 82242 1 5199
2 82243 1 5199
2 82244 1 5201
2 82245 1 5201
2 82246 1 5201
2 82247 1 5201
2 82248 1 5208
2 82249 1 5208
2 82250 1 5216
2 82251 1 5216
2 82252 1 5216
2 82253 1 5217
2 82254 1 5217
2 82255 1 5217
2 82256 1 5217
2 82257 1 5217
2 82258 1 5224
2 82259 1 5224
2 82260 1 5224
2 82261 1 5224
2 82262 1 5224
2 82263 1 5224
2 82264 1 5224
2 82265 1 5224
2 82266 1 5224
2 82267 1 5224
2 82268 1 5224
2 82269 1 5224
2 82270 1 5224
2 82271 1 5224
2 82272 1 5224
2 82273 1 5224
2 82274 1 5224
2 82275 1 5224
2 82276 1 5224
2 82277 1 5224
2 82278 1 5224
2 82279 1 5225
2 82280 1 5225
2 82281 1 5225
2 82282 1 5225
2 82283 1 5225
2 82284 1 5225
2 82285 1 5225
2 82286 1 5225
2 82287 1 5225
2 82288 1 5225
2 82289 1 5225
2 82290 1 5225
2 82291 1 5227
2 82292 1 5227
2 82293 1 5231
2 82294 1 5231
2 82295 1 5231
2 82296 1 5231
2 82297 1 5232
2 82298 1 5232
2 82299 1 5232
2 82300 1 5235
2 82301 1 5235
2 82302 1 5235
2 82303 1 5235
2 82304 1 5235
2 82305 1 5235
2 82306 1 5235
2 82307 1 5235
2 82308 1 5235
2 82309 1 5235
2 82310 1 5235
2 82311 1 5235
2 82312 1 5236
2 82313 1 5236
2 82314 1 5237
2 82315 1 5237
2 82316 1 5238
2 82317 1 5238
2 82318 1 5238
2 82319 1 5238
2 82320 1 5238
2 82321 1 5238
2 82322 1 5238
2 82323 1 5238
2 82324 1 5238
2 82325 1 5238
2 82326 1 5238
2 82327 1 5238
2 82328 1 5238
2 82329 1 5238
2 82330 1 5240
2 82331 1 5240
2 82332 1 5240
2 82333 1 5250
2 82334 1 5250
2 82335 1 5260
2 82336 1 5260
2 82337 1 5260
2 82338 1 5260
2 82339 1 5260
2 82340 1 5260
2 82341 1 5260
2 82342 1 5260
2 82343 1 5260
2 82344 1 5260
2 82345 1 5260
2 82346 1 5260
2 82347 1 5260
2 82348 1 5260
2 82349 1 5260
2 82350 1 5261
2 82351 1 5261
2 82352 1 5261
2 82353 1 5261
2 82354 1 5261
2 82355 1 5261
2 82356 1 5262
2 82357 1 5262
2 82358 1 5262
2 82359 1 5275
2 82360 1 5275
2 82361 1 5277
2 82362 1 5277
2 82363 1 5277
2 82364 1 5277
2 82365 1 5277
2 82366 1 5277
2 82367 1 5277
2 82368 1 5277
2 82369 1 5277
2 82370 1 5277
2 82371 1 5277
2 82372 1 5277
2 82373 1 5277
2 82374 1 5277
2 82375 1 5277
2 82376 1 5277
2 82377 1 5277
2 82378 1 5278
2 82379 1 5278
2 82380 1 5278
2 82381 1 5278
2 82382 1 5278
2 82383 1 5278
2 82384 1 5278
2 82385 1 5278
2 82386 1 5278
2 82387 1 5278
2 82388 1 5279
2 82389 1 5279
2 82390 1 5280
2 82391 1 5280
2 82392 1 5284
2 82393 1 5284
2 82394 1 5284
2 82395 1 5284
2 82396 1 5284
2 82397 1 5284
2 82398 1 5284
2 82399 1 5284
2 82400 1 5284
2 82401 1 5284
2 82402 1 5284
2 82403 1 5284
2 82404 1 5284
2 82405 1 5284
2 82406 1 5284
2 82407 1 5284
2 82408 1 5284
2 82409 1 5284
2 82410 1 5284
2 82411 1 5284
2 82412 1 5284
2 82413 1 5284
2 82414 1 5284
2 82415 1 5284
2 82416 1 5284
2 82417 1 5284
2 82418 1 5284
2 82419 1 5284
2 82420 1 5284
2 82421 1 5284
2 82422 1 5284
2 82423 1 5285
2 82424 1 5285
2 82425 1 5285
2 82426 1 5286
2 82427 1 5286
2 82428 1 5287
2 82429 1 5287
2 82430 1 5295
2 82431 1 5295
2 82432 1 5295
2 82433 1 5296
2 82434 1 5296
2 82435 1 5298
2 82436 1 5298
2 82437 1 5299
2 82438 1 5299
2 82439 1 5300
2 82440 1 5300
2 82441 1 5305
2 82442 1 5305
2 82443 1 5317
2 82444 1 5317
2 82445 1 5318
2 82446 1 5318
2 82447 1 5320
2 82448 1 5320
2 82449 1 5320
2 82450 1 5322
2 82451 1 5322
2 82452 1 5323
2 82453 1 5323
2 82454 1 5324
2 82455 1 5324
2 82456 1 5325
2 82457 1 5325
2 82458 1 5325
2 82459 1 5325
2 82460 1 5325
2 82461 1 5325
2 82462 1 5325
2 82463 1 5325
2 82464 1 5326
2 82465 1 5326
2 82466 1 5326
2 82467 1 5330
2 82468 1 5330
2 82469 1 5330
2 82470 1 5330
2 82471 1 5330
2 82472 1 5331
2 82473 1 5331
2 82474 1 5331
2 82475 1 5339
2 82476 1 5339
2 82477 1 5347
2 82478 1 5347
2 82479 1 5348
2 82480 1 5348
2 82481 1 5348
2 82482 1 5348
2 82483 1 5359
2 82484 1 5359
2 82485 1 5359
2 82486 1 5362
2 82487 1 5362
2 82488 1 5364
2 82489 1 5364
2 82490 1 5365
2 82491 1 5365
2 82492 1 5365
2 82493 1 5365
2 82494 1 5366
2 82495 1 5366
2 82496 1 5366
2 82497 1 5366
2 82498 1 5366
2 82499 1 5366
2 82500 1 5366
2 82501 1 5366
2 82502 1 5366
2 82503 1 5366
2 82504 1 5366
2 82505 1 5367
2 82506 1 5367
2 82507 1 5377
2 82508 1 5377
2 82509 1 5377
2 82510 1 5387
2 82511 1 5387
2 82512 1 5387
2 82513 1 5387
2 82514 1 5387
2 82515 1 5387
2 82516 1 5387
2 82517 1 5388
2 82518 1 5388
2 82519 1 5388
2 82520 1 5388
2 82521 1 5389
2 82522 1 5389
2 82523 1 5389
2 82524 1 5389
2 82525 1 5389
2 82526 1 5390
2 82527 1 5390
2 82528 1 5390
2 82529 1 5394
2 82530 1 5394
2 82531 1 5394
2 82532 1 5395
2 82533 1 5395
2 82534 1 5395
2 82535 1 5403
2 82536 1 5403
2 82537 1 5404
2 82538 1 5404
2 82539 1 5411
2 82540 1 5411
2 82541 1 5411
2 82542 1 5411
2 82543 1 5425
2 82544 1 5425
2 82545 1 5425
2 82546 1 5427
2 82547 1 5427
2 82548 1 5436
2 82549 1 5436
2 82550 1 5448
2 82551 1 5448
2 82552 1 5448
2 82553 1 5448
2 82554 1 5448
2 82555 1 5448
2 82556 1 5448
2 82557 1 5448
2 82558 1 5450
2 82559 1 5450
2 82560 1 5450
2 82561 1 5450
2 82562 1 5450
2 82563 1 5450
2 82564 1 5450
2 82565 1 5451
2 82566 1 5451
2 82567 1 5451
2 82568 1 5451
2 82569 1 5451
2 82570 1 5451
2 82571 1 5451
2 82572 1 5451
2 82573 1 5451
2 82574 1 5451
2 82575 1 5451
2 82576 1 5451
2 82577 1 5451
2 82578 1 5451
2 82579 1 5451
2 82580 1 5451
2 82581 1 5463
2 82582 1 5463
2 82583 1 5463
2 82584 1 5463
2 82585 1 5482
2 82586 1 5482
2 82587 1 5482
2 82588 1 5482
2 82589 1 5482
2 82590 1 5482
2 82591 1 5482
2 82592 1 5483
2 82593 1 5483
2 82594 1 5483
2 82595 1 5484
2 82596 1 5484
2 82597 1 5485
2 82598 1 5485
2 82599 1 5485
2 82600 1 5485
2 82601 1 5485
2 82602 1 5485
2 82603 1 5485
2 82604 1 5485
2 82605 1 5485
2 82606 1 5485
2 82607 1 5485
2 82608 1 5485
2 82609 1 5485
2 82610 1 5485
2 82611 1 5485
2 82612 1 5485
2 82613 1 5485
2 82614 1 5485
2 82615 1 5485
2 82616 1 5485
2 82617 1 5485
2 82618 1 5485
2 82619 1 5486
2 82620 1 5486
2 82621 1 5487
2 82622 1 5487
2 82623 1 5489
2 82624 1 5489
2 82625 1 5489
2 82626 1 5489
2 82627 1 5489
2 82628 1 5497
2 82629 1 5497
2 82630 1 5497
2 82631 1 5498
2 82632 1 5498
2 82633 1 5498
2 82634 1 5503
2 82635 1 5503
2 82636 1 5506
2 82637 1 5506
2 82638 1 5508
2 82639 1 5508
2 82640 1 5508
2 82641 1 5509
2 82642 1 5509
2 82643 1 5509
2 82644 1 5509
2 82645 1 5509
2 82646 1 5509
2 82647 1 5509
2 82648 1 5509
2 82649 1 5509
2 82650 1 5509
2 82651 1 5509
2 82652 1 5509
2 82653 1 5509
2 82654 1 5509
2 82655 1 5509
2 82656 1 5509
2 82657 1 5509
2 82658 1 5509
2 82659 1 5509
2 82660 1 5509
2 82661 1 5510
2 82662 1 5510
2 82663 1 5510
2 82664 1 5510
2 82665 1 5517
2 82666 1 5517
2 82667 1 5518
2 82668 1 5518
2 82669 1 5518
2 82670 1 5522
2 82671 1 5522
2 82672 1 5523
2 82673 1 5523
2 82674 1 5523
2 82675 1 5523
2 82676 1 5523
2 82677 1 5523
2 82678 1 5523
2 82679 1 5523
2 82680 1 5523
2 82681 1 5523
2 82682 1 5524
2 82683 1 5524
2 82684 1 5524
2 82685 1 5524
2 82686 1 5533
2 82687 1 5533
2 82688 1 5535
2 82689 1 5535
2 82690 1 5588
2 82691 1 5588
2 82692 1 5595
2 82693 1 5595
2 82694 1 5595
2 82695 1 5608
2 82696 1 5608
2 82697 1 5608
2 82698 1 5608
2 82699 1 5608
2 82700 1 5609
2 82701 1 5609
2 82702 1 5610
2 82703 1 5610
2 82704 1 5611
2 82705 1 5611
2 82706 1 5620
2 82707 1 5620
2 82708 1 5628
2 82709 1 5628
2 82710 1 5628
2 82711 1 5628
2 82712 1 5629
2 82713 1 5629
2 82714 1 5642
2 82715 1 5642
2 82716 1 5642
2 82717 1 5644
2 82718 1 5644
2 82719 1 5644
2 82720 1 5644
2 82721 1 5644
2 82722 1 5644
2 82723 1 5644
2 82724 1 5655
2 82725 1 5655
2 82726 1 5655
2 82727 1 5657
2 82728 1 5657
2 82729 1 5657
2 82730 1 5668
2 82731 1 5668
2 82732 1 5668
2 82733 1 5668
2 82734 1 5668
2 82735 1 5669
2 82736 1 5669
2 82737 1 5669
2 82738 1 5669
2 82739 1 5670
2 82740 1 5670
2 82741 1 5678
2 82742 1 5678
2 82743 1 5678
2 82744 1 5678
2 82745 1 5679
2 82746 1 5679
2 82747 1 5679
2 82748 1 5701
2 82749 1 5701
2 82750 1 5701
2 82751 1 5739
2 82752 1 5739
2 82753 1 5739
2 82754 1 5739
2 82755 1 5739
2 82756 1 5748
2 82757 1 5748
2 82758 1 5748
2 82759 1 5749
2 82760 1 5749
2 82761 1 5749
2 82762 1 5757
2 82763 1 5757
2 82764 1 5757
2 82765 1 5757
2 82766 1 5760
2 82767 1 5760
2 82768 1 5760
2 82769 1 5769
2 82770 1 5769
2 82771 1 5769
2 82772 1 5769
2 82773 1 5770
2 82774 1 5770
2 82775 1 5770
2 82776 1 5770
2 82777 1 5770
2 82778 1 5778
2 82779 1 5778
2 82780 1 5778
2 82781 1 5778
2 82782 1 5778
2 82783 1 5778
2 82784 1 5778
2 82785 1 5779
2 82786 1 5779
2 82787 1 5779
2 82788 1 5779
2 82789 1 5779
2 82790 1 5779
2 82791 1 5779
2 82792 1 5779
2 82793 1 5779
2 82794 1 5779
2 82795 1 5780
2 82796 1 5780
2 82797 1 5781
2 82798 1 5781
2 82799 1 5781
2 82800 1 5781
2 82801 1 5781
2 82802 1 5781
2 82803 1 5781
2 82804 1 5781
2 82805 1 5781
2 82806 1 5781
2 82807 1 5781
2 82808 1 5781
2 82809 1 5781
2 82810 1 5781
2 82811 1 5781
2 82812 1 5793
2 82813 1 5793
2 82814 1 5793
2 82815 1 5793
2 82816 1 5793
2 82817 1 5795
2 82818 1 5795
2 82819 1 5795
2 82820 1 5795
2 82821 1 5795
2 82822 1 5795
2 82823 1 5808
2 82824 1 5808
2 82825 1 5809
2 82826 1 5809
2 82827 1 5870
2 82828 1 5870
2 82829 1 5870
2 82830 1 5870
2 82831 1 5870
2 82832 1 5870
2 82833 1 5870
2 82834 1 5870
2 82835 1 5870
2 82836 1 5871
2 82837 1 5871
2 82838 1 5874
2 82839 1 5874
2 82840 1 5874
2 82841 1 5874
2 82842 1 5886
2 82843 1 5886
2 82844 1 5886
2 82845 1 5886
2 82846 1 5886
2 82847 1 5886
2 82848 1 5888
2 82849 1 5888
2 82850 1 5889
2 82851 1 5889
2 82852 1 5908
2 82853 1 5908
2 82854 1 5908
2 82855 1 5908
2 82856 1 5912
2 82857 1 5912
2 82858 1 5923
2 82859 1 5923
2 82860 1 5923
2 82861 1 5923
2 82862 1 5923
2 82863 1 5923
2 82864 1 5923
2 82865 1 5923
2 82866 1 5923
2 82867 1 5925
2 82868 1 5925
2 82869 1 5925
2 82870 1 5926
2 82871 1 5926
2 82872 1 5938
2 82873 1 5938
2 82874 1 5938
2 82875 1 5938
2 82876 1 5965
2 82877 1 5965
2 82878 1 5968
2 82879 1 5968
2 82880 1 5969
2 82881 1 5969
2 82882 1 5977
2 82883 1 5977
2 82884 1 5978
2 82885 1 5978
2 82886 1 5978
2 82887 1 5978
2 82888 1 5979
2 82889 1 5979
2 82890 1 5979
2 82891 1 5987
2 82892 1 5987
2 82893 1 5987
2 82894 1 5988
2 82895 1 5988
2 82896 1 6001
2 82897 1 6001
2 82898 1 6001
2 82899 1 6001
2 82900 1 6001
2 82901 1 6002
2 82902 1 6002
2 82903 1 6002
2 82904 1 6003
2 82905 1 6003
2 82906 1 6003
2 82907 1 6003
2 82908 1 6003
2 82909 1 6003
2 82910 1 6003
2 82911 1 6003
2 82912 1 6007
2 82913 1 6007
2 82914 1 6007
2 82915 1 6007
2 82916 1 6007
2 82917 1 6007
2 82918 1 6007
2 82919 1 6007
2 82920 1 6007
2 82921 1 6007
2 82922 1 6007
2 82923 1 6007
2 82924 1 6007
2 82925 1 6007
2 82926 1 6007
2 82927 1 6007
2 82928 1 6007
2 82929 1 6007
2 82930 1 6007
2 82931 1 6007
2 82932 1 6007
2 82933 1 6007
2 82934 1 6007
2 82935 1 6007
2 82936 1 6007
2 82937 1 6008
2 82938 1 6008
2 82939 1 6008
2 82940 1 6008
2 82941 1 6008
2 82942 1 6008
2 82943 1 6008
2 82944 1 6008
2 82945 1 6008
2 82946 1 6008
2 82947 1 6008
2 82948 1 6008
2 82949 1 6008
2 82950 1 6008
2 82951 1 6008
2 82952 1 6008
2 82953 1 6010
2 82954 1 6010
2 82955 1 6010
2 82956 1 6010
2 82957 1 6010
2 82958 1 6010
2 82959 1 6010
2 82960 1 6010
2 82961 1 6010
2 82962 1 6010
2 82963 1 6010
2 82964 1 6010
2 82965 1 6011
2 82966 1 6011
2 82967 1 6011
2 82968 1 6021
2 82969 1 6021
2 82970 1 6021
2 82971 1 6021
2 82972 1 6021
2 82973 1 6021
2 82974 1 6021
2 82975 1 6021
2 82976 1 6021
2 82977 1 6021
2 82978 1 6021
2 82979 1 6021
2 82980 1 6021
2 82981 1 6021
2 82982 1 6021
2 82983 1 6021
2 82984 1 6021
2 82985 1 6022
2 82986 1 6022
2 82987 1 6022
2 82988 1 6022
2 82989 1 6025
2 82990 1 6025
2 82991 1 6025
2 82992 1 6025
2 82993 1 6025
2 82994 1 6025
2 82995 1 6025
2 82996 1 6028
2 82997 1 6028
2 82998 1 6033
2 82999 1 6033
2 83000 1 6033
2 83001 1 6033
2 83002 1 6033
2 83003 1 6033
2 83004 1 6034
2 83005 1 6034
2 83006 1 6046
2 83007 1 6046
2 83008 1 6046
2 83009 1 6046
2 83010 1 6046
2 83011 1 6046
2 83012 1 6046
2 83013 1 6049
2 83014 1 6049
2 83015 1 6050
2 83016 1 6050
2 83017 1 6050
2 83018 1 6050
2 83019 1 6050
2 83020 1 6050
2 83021 1 6050
2 83022 1 6051
2 83023 1 6051
2 83024 1 6051
2 83025 1 6051
2 83026 1 6051
2 83027 1 6051
2 83028 1 6051
2 83029 1 6051
2 83030 1 6052
2 83031 1 6052
2 83032 1 6052
2 83033 1 6061
2 83034 1 6061
2 83035 1 6061
2 83036 1 6061
2 83037 1 6061
2 83038 1 6061
2 83039 1 6061
2 83040 1 6062
2 83041 1 6062
2 83042 1 6062
2 83043 1 6062
2 83044 1 6062
2 83045 1 6063
2 83046 1 6063
2 83047 1 6063
2 83048 1 6070
2 83049 1 6070
2 83050 1 6070
2 83051 1 6070
2 83052 1 6070
2 83053 1 6070
2 83054 1 6070
2 83055 1 6070
2 83056 1 6070
2 83057 1 6070
2 83058 1 6070
2 83059 1 6070
2 83060 1 6070
2 83061 1 6070
2 83062 1 6070
2 83063 1 6070
2 83064 1 6070
2 83065 1 6070
2 83066 1 6070
2 83067 1 6071
2 83068 1 6071
2 83069 1 6072
2 83070 1 6072
2 83071 1 6072
2 83072 1 6073
2 83073 1 6073
2 83074 1 6084
2 83075 1 6084
2 83076 1 6101
2 83077 1 6101
2 83078 1 6142
2 83079 1 6142
2 83080 1 6148
2 83081 1 6148
2 83082 1 6164
2 83083 1 6164
2 83084 1 6171
2 83085 1 6171
2 83086 1 6171
2 83087 1 6171
2 83088 1 6171
2 83089 1 6171
2 83090 1 6171
2 83091 1 6171
2 83092 1 6171
2 83093 1 6171
2 83094 1 6171
2 83095 1 6171
2 83096 1 6171
2 83097 1 6171
2 83098 1 6171
2 83099 1 6171
2 83100 1 6171
2 83101 1 6171
2 83102 1 6171
2 83103 1 6171
2 83104 1 6171
2 83105 1 6171
2 83106 1 6171
2 83107 1 6171
2 83108 1 6171
2 83109 1 6171
2 83110 1 6171
2 83111 1 6171
2 83112 1 6171
2 83113 1 6171
2 83114 1 6171
2 83115 1 6171
2 83116 1 6171
2 83117 1 6172
2 83118 1 6172
2 83119 1 6172
2 83120 1 6172
2 83121 1 6172
2 83122 1 6188
2 83123 1 6188
2 83124 1 6189
2 83125 1 6189
2 83126 1 6189
2 83127 1 6193
2 83128 1 6193
2 83129 1 6195
2 83130 1 6195
2 83131 1 6209
2 83132 1 6209
2 83133 1 6213
2 83134 1 6213
2 83135 1 6213
2 83136 1 6213
2 83137 1 6214
2 83138 1 6214
2 83139 1 6214
2 83140 1 6226
2 83141 1 6226
2 83142 1 6232
2 83143 1 6232
2 83144 1 6232
2 83145 1 6233
2 83146 1 6233
2 83147 1 6272
2 83148 1 6272
2 83149 1 6272
2 83150 1 6272
2 83151 1 6272
2 83152 1 6272
2 83153 1 6272
2 83154 1 6272
2 83155 1 6272
2 83156 1 6280
2 83157 1 6280
2 83158 1 6280
2 83159 1 6280
2 83160 1 6281
2 83161 1 6281
2 83162 1 6282
2 83163 1 6282
2 83164 1 6285
2 83165 1 6285
2 83166 1 6285
2 83167 1 6285
2 83168 1 6285
2 83169 1 6286
2 83170 1 6286
2 83171 1 6293
2 83172 1 6293
2 83173 1 6302
2 83174 1 6302
2 83175 1 6302
2 83176 1 6321
2 83177 1 6321
2 83178 1 6336
2 83179 1 6336
2 83180 1 6337
2 83181 1 6337
2 83182 1 6337
2 83183 1 6337
2 83184 1 6337
2 83185 1 6337
2 83186 1 6337
2 83187 1 6337
2 83188 1 6337
2 83189 1 6337
2 83190 1 6337
2 83191 1 6337
2 83192 1 6337
2 83193 1 6337
2 83194 1 6337
2 83195 1 6337
2 83196 1 6337
2 83197 1 6337
2 83198 1 6337
2 83199 1 6337
2 83200 1 6337
2 83201 1 6338
2 83202 1 6338
2 83203 1 6338
2 83204 1 6338
2 83205 1 6338
2 83206 1 6338
2 83207 1 6338
2 83208 1 6338
2 83209 1 6347
2 83210 1 6347
2 83211 1 6348
2 83212 1 6348
2 83213 1 6348
2 83214 1 6359
2 83215 1 6359
2 83216 1 6359
2 83217 1 6359
2 83218 1 6359
2 83219 1 6359
2 83220 1 6360
2 83221 1 6360
2 83222 1 6360
2 83223 1 6361
2 83224 1 6361
2 83225 1 6365
2 83226 1 6365
2 83227 1 6365
2 83228 1 6374
2 83229 1 6374
2 83230 1 6380
2 83231 1 6380
2 83232 1 6380
2 83233 1 6381
2 83234 1 6381
2 83235 1 6384
2 83236 1 6384
2 83237 1 6402
2 83238 1 6402
2 83239 1 6408
2 83240 1 6408
2 83241 1 6410
2 83242 1 6410
2 83243 1 6413
2 83244 1 6413
2 83245 1 6413
2 83246 1 6413
2 83247 1 6413
2 83248 1 6413
2 83249 1 6413
2 83250 1 6413
2 83251 1 6413
2 83252 1 6413
2 83253 1 6413
2 83254 1 6414
2 83255 1 6414
2 83256 1 6418
2 83257 1 6418
2 83258 1 6427
2 83259 1 6427
2 83260 1 6428
2 83261 1 6428
2 83262 1 6428
2 83263 1 6431
2 83264 1 6431
2 83265 1 6432
2 83266 1 6432
2 83267 1 6433
2 83268 1 6433
2 83269 1 6434
2 83270 1 6434
2 83271 1 6434
2 83272 1 6449
2 83273 1 6449
2 83274 1 6451
2 83275 1 6451
2 83276 1 6462
2 83277 1 6462
2 83278 1 6464
2 83279 1 6464
2 83280 1 6466
2 83281 1 6466
2 83282 1 6472
2 83283 1 6472
2 83284 1 6488
2 83285 1 6488
2 83286 1 6488
2 83287 1 6488
2 83288 1 6489
2 83289 1 6489
2 83290 1 6489
2 83291 1 6489
2 83292 1 6489
2 83293 1 6498
2 83294 1 6498
2 83295 1 6511
2 83296 1 6511
2 83297 1 6515
2 83298 1 6515
2 83299 1 6515
2 83300 1 6515
2 83301 1 6515
2 83302 1 6515
2 83303 1 6515
2 83304 1 6515
2 83305 1 6515
2 83306 1 6515
2 83307 1 6516
2 83308 1 6516
2 83309 1 6516
2 83310 1 6516
2 83311 1 6516
2 83312 1 6516
2 83313 1 6517
2 83314 1 6517
2 83315 1 6561
2 83316 1 6561
2 83317 1 6562
2 83318 1 6562
2 83319 1 6573
2 83320 1 6573
2 83321 1 6573
2 83322 1 6574
2 83323 1 6574
2 83324 1 6574
2 83325 1 6582
2 83326 1 6582
2 83327 1 6582
2 83328 1 6582
2 83329 1 6582
2 83330 1 6582
2 83331 1 6583
2 83332 1 6583
2 83333 1 6583
2 83334 1 6583
2 83335 1 6583
2 83336 1 6583
2 83337 1 6583
2 83338 1 6583
2 83339 1 6590
2 83340 1 6590
2 83341 1 6590
2 83342 1 6590
2 83343 1 6590
2 83344 1 6590
2 83345 1 6590
2 83346 1 6590
2 83347 1 6591
2 83348 1 6591
2 83349 1 6591
2 83350 1 6591
2 83351 1 6591
2 83352 1 6591
2 83353 1 6591
2 83354 1 6591
2 83355 1 6599
2 83356 1 6599
2 83357 1 6599
2 83358 1 6599
2 83359 1 6599
2 83360 1 6599
2 83361 1 6613
2 83362 1 6613
2 83363 1 6619
2 83364 1 6619
2 83365 1 6619
2 83366 1 6619
2 83367 1 6620
2 83368 1 6620
2 83369 1 6639
2 83370 1 6639
2 83371 1 6640
2 83372 1 6640
2 83373 1 6650
2 83374 1 6650
2 83375 1 6650
2 83376 1 6650
2 83377 1 6651
2 83378 1 6651
2 83379 1 6651
2 83380 1 6654
2 83381 1 6654
2 83382 1 6654
2 83383 1 6654
2 83384 1 6654
2 83385 1 6666
2 83386 1 6666
2 83387 1 6676
2 83388 1 6676
2 83389 1 6688
2 83390 1 6688
2 83391 1 6689
2 83392 1 6689
2 83393 1 6691
2 83394 1 6691
2 83395 1 6704
2 83396 1 6704
2 83397 1 6704
2 83398 1 6704
2 83399 1 6704
2 83400 1 6704
2 83401 1 6704
2 83402 1 6704
2 83403 1 6704
2 83404 1 6704
2 83405 1 6704
2 83406 1 6704
2 83407 1 6704
2 83408 1 6704
2 83409 1 6704
2 83410 1 6704
2 83411 1 6705
2 83412 1 6705
2 83413 1 6705
2 83414 1 6705
2 83415 1 6705
2 83416 1 6705
2 83417 1 6705
2 83418 1 6705
2 83419 1 6706
2 83420 1 6706
2 83421 1 6712
2 83422 1 6712
2 83423 1 6713
2 83424 1 6713
2 83425 1 6713
2 83426 1 6713
2 83427 1 6713
2 83428 1 6726
2 83429 1 6726
2 83430 1 6726
2 83431 1 6726
2 83432 1 6726
2 83433 1 6726
2 83434 1 6734
2 83435 1 6734
2 83436 1 6734
2 83437 1 6752
2 83438 1 6752
2 83439 1 6752
2 83440 1 6752
2 83441 1 6752
2 83442 1 6763
2 83443 1 6763
2 83444 1 6763
2 83445 1 6763
2 83446 1 6763
2 83447 1 6763
2 83448 1 6763
2 83449 1 6763
2 83450 1 6763
2 83451 1 6774
2 83452 1 6774
2 83453 1 6774
2 83454 1 6775
2 83455 1 6775
2 83456 1 6775
2 83457 1 6776
2 83458 1 6776
2 83459 1 6776
2 83460 1 6776
2 83461 1 6776
2 83462 1 6777
2 83463 1 6777
2 83464 1 6778
2 83465 1 6778
2 83466 1 6778
2 83467 1 6778
2 83468 1 6778
2 83469 1 6779
2 83470 1 6779
2 83471 1 6779
2 83472 1 6779
2 83473 1 6780
2 83474 1 6780
2 83475 1 6780
2 83476 1 6780
2 83477 1 6780
2 83478 1 6780
2 83479 1 6780
2 83480 1 6780
2 83481 1 6781
2 83482 1 6781
2 83483 1 6781
2 83484 1 6781
2 83485 1 6781
2 83486 1 6781
2 83487 1 6782
2 83488 1 6782
2 83489 1 6782
2 83490 1 6782
2 83491 1 6782
2 83492 1 6782
2 83493 1 6782
2 83494 1 6782
2 83495 1 6782
2 83496 1 6782
2 83497 1 6782
2 83498 1 6783
2 83499 1 6783
2 83500 1 6783
2 83501 1 6783
2 83502 1 6801
2 83503 1 6801
2 83504 1 6801
2 83505 1 6809
2 83506 1 6809
2 83507 1 6811
2 83508 1 6811
2 83509 1 6811
2 83510 1 6811
2 83511 1 6811
2 83512 1 6812
2 83513 1 6812
2 83514 1 6820
2 83515 1 6820
2 83516 1 6820
2 83517 1 6820
2 83518 1 6820
2 83519 1 6820
2 83520 1 6820
2 83521 1 6820
2 83522 1 6820
2 83523 1 6820
2 83524 1 6820
2 83525 1 6820
2 83526 1 6820
2 83527 1 6820
2 83528 1 6820
2 83529 1 6820
2 83530 1 6820
2 83531 1 6820
2 83532 1 6820
2 83533 1 6820
2 83534 1 6820
2 83535 1 6820
2 83536 1 6820
2 83537 1 6820
2 83538 1 6820
2 83539 1 6820
2 83540 1 6820
2 83541 1 6820
2 83542 1 6820
2 83543 1 6820
2 83544 1 6820
2 83545 1 6820
2 83546 1 6820
2 83547 1 6820
2 83548 1 6820
2 83549 1 6820
2 83550 1 6820
2 83551 1 6820
2 83552 1 6820
2 83553 1 6820
2 83554 1 6820
2 83555 1 6820
2 83556 1 6820
2 83557 1 6820
2 83558 1 6820
2 83559 1 6820
2 83560 1 6820
2 83561 1 6820
2 83562 1 6820
2 83563 1 6820
2 83564 1 6820
2 83565 1 6820
2 83566 1 6820
2 83567 1 6820
2 83568 1 6820
2 83569 1 6820
2 83570 1 6820
2 83571 1 6820
2 83572 1 6820
2 83573 1 6820
2 83574 1 6820
2 83575 1 6821
2 83576 1 6821
2 83577 1 6821
2 83578 1 6829
2 83579 1 6829
2 83580 1 6829
2 83581 1 6829
2 83582 1 6829
2 83583 1 6829
2 83584 1 6829
2 83585 1 6829
2 83586 1 6829
2 83587 1 6829
2 83588 1 6829
2 83589 1 6829
2 83590 1 6829
2 83591 1 6829
2 83592 1 6830
2 83593 1 6830
2 83594 1 6830
2 83595 1 6830
2 83596 1 6831
2 83597 1 6831
2 83598 1 6832
2 83599 1 6832
2 83600 1 6832
2 83601 1 6832
2 83602 1 6832
2 83603 1 6832
2 83604 1 6833
2 83605 1 6833
2 83606 1 6833
2 83607 1 6833
2 83608 1 6834
2 83609 1 6834
2 83610 1 6834
2 83611 1 6841
2 83612 1 6841
2 83613 1 6847
2 83614 1 6847
2 83615 1 6847
2 83616 1 6847
2 83617 1 6854
2 83618 1 6854
2 83619 1 6854
2 83620 1 6854
2 83621 1 6854
2 83622 1 6854
2 83623 1 6854
2 83624 1 6854
2 83625 1 6854
2 83626 1 6854
2 83627 1 6854
2 83628 1 6854
2 83629 1 6854
2 83630 1 6854
2 83631 1 6854
2 83632 1 6867
2 83633 1 6867
2 83634 1 6867
2 83635 1 6867
2 83636 1 6867
2 83637 1 6867
2 83638 1 6867
2 83639 1 6867
2 83640 1 6867
2 83641 1 6869
2 83642 1 6869
2 83643 1 6870
2 83644 1 6870
2 83645 1 6876
2 83646 1 6876
2 83647 1 6876
2 83648 1 6876
2 83649 1 6876
2 83650 1 6876
2 83651 1 6876
2 83652 1 6876
2 83653 1 6889
2 83654 1 6889
2 83655 1 6890
2 83656 1 6890
2 83657 1 6890
2 83658 1 6897
2 83659 1 6897
2 83660 1 6897
2 83661 1 6897
2 83662 1 6897
2 83663 1 6897
2 83664 1 6897
2 83665 1 6897
2 83666 1 6897
2 83667 1 6897
2 83668 1 6911
2 83669 1 6911
2 83670 1 6911
2 83671 1 6911
2 83672 1 6911
2 83673 1 6911
2 83674 1 6911
2 83675 1 6911
2 83676 1 6911
2 83677 1 6912
2 83678 1 6912
2 83679 1 6912
2 83680 1 6915
2 83681 1 6915
2 83682 1 6915
2 83683 1 6915
2 83684 1 6915
2 83685 1 6916
2 83686 1 6916
2 83687 1 6916
2 83688 1 6916
2 83689 1 6942
2 83690 1 6942
2 83691 1 6942
2 83692 1 6945
2 83693 1 6945
2 83694 1 6948
2 83695 1 6948
2 83696 1 6948
2 83697 1 6948
2 83698 1 6948
2 83699 1 6948
2 83700 1 6948
2 83701 1 6948
2 83702 1 6948
2 83703 1 6948
2 83704 1 6948
2 83705 1 6948
2 83706 1 6948
2 83707 1 6948
2 83708 1 6948
2 83709 1 6949
2 83710 1 6949
2 83711 1 6949
2 83712 1 6949
2 83713 1 6949
2 83714 1 6949
2 83715 1 6949
2 83716 1 6949
2 83717 1 6949
2 83718 1 6949
2 83719 1 6949
2 83720 1 6949
2 83721 1 6949
2 83722 1 6949
2 83723 1 6950
2 83724 1 6950
2 83725 1 6950
2 83726 1 6950
2 83727 1 6950
2 83728 1 6950
2 83729 1 6951
2 83730 1 6951
2 83731 1 6951
2 83732 1 6951
2 83733 1 6951
2 83734 1 6951
2 83735 1 6951
2 83736 1 6951
2 83737 1 6951
2 83738 1 6951
2 83739 1 6951
2 83740 1 6951
2 83741 1 6951
2 83742 1 6951
2 83743 1 6951
2 83744 1 6951
2 83745 1 6951
2 83746 1 6951
2 83747 1 6951
2 83748 1 6951
2 83749 1 6951
2 83750 1 6951
2 83751 1 6951
2 83752 1 6951
2 83753 1 6951
2 83754 1 6951
2 83755 1 6951
2 83756 1 6951
2 83757 1 6952
2 83758 1 6952
2 83759 1 6952
2 83760 1 6952
2 83761 1 6952
2 83762 1 6952
2 83763 1 6952
2 83764 1 6953
2 83765 1 6953
2 83766 1 6953
2 83767 1 6953
2 83768 1 6953
2 83769 1 6963
2 83770 1 6963
2 83771 1 6964
2 83772 1 6964
2 83773 1 6965
2 83774 1 6965
2 83775 1 6965
2 83776 1 6966
2 83777 1 6966
2 83778 1 6988
2 83779 1 6988
2 83780 1 6988
2 83781 1 6988
2 83782 1 6988
2 83783 1 6988
2 83784 1 6988
2 83785 1 6988
2 83786 1 6988
2 83787 1 6989
2 83788 1 6989
2 83789 1 6990
2 83790 1 6990
2 83791 1 6997
2 83792 1 6997
2 83793 1 6997
2 83794 1 6997
2 83795 1 6997
2 83796 1 6998
2 83797 1 6998
2 83798 1 6999
2 83799 1 6999
2 83800 1 7001
2 83801 1 7001
2 83802 1 7002
2 83803 1 7002
2 83804 1 7002
2 83805 1 7002
2 83806 1 7002
2 83807 1 7002
2 83808 1 7002
2 83809 1 7002
2 83810 1 7002
2 83811 1 7003
2 83812 1 7003
2 83813 1 7003
2 83814 1 7004
2 83815 1 7004
2 83816 1 7004
2 83817 1 7004
2 83818 1 7004
2 83819 1 7006
2 83820 1 7006
2 83821 1 7006
2 83822 1 7006
2 83823 1 7007
2 83824 1 7007
2 83825 1 7012
2 83826 1 7012
2 83827 1 7012
2 83828 1 7012
2 83829 1 7012
2 83830 1 7012
2 83831 1 7012
2 83832 1 7012
2 83833 1 7032
2 83834 1 7032
2 83835 1 7032
2 83836 1 7044
2 83837 1 7044
2 83838 1 7044
2 83839 1 7044
2 83840 1 7044
2 83841 1 7044
2 83842 1 7044
2 83843 1 7044
2 83844 1 7044
2 83845 1 7044
2 83846 1 7044
2 83847 1 7044
2 83848 1 7044
2 83849 1 7044
2 83850 1 7044
2 83851 1 7044
2 83852 1 7044
2 83853 1 7047
2 83854 1 7047
2 83855 1 7050
2 83856 1 7050
2 83857 1 7066
2 83858 1 7066
2 83859 1 7067
2 83860 1 7067
2 83861 1 7077
2 83862 1 7077
2 83863 1 7077
2 83864 1 7084
2 83865 1 7084
2 83866 1 7084
2 83867 1 7084
2 83868 1 7084
2 83869 1 7084
2 83870 1 7084
2 83871 1 7084
2 83872 1 7085
2 83873 1 7085
2 83874 1 7085
2 83875 1 7085
2 83876 1 7085
2 83877 1 7085
2 83878 1 7085
2 83879 1 7085
2 83880 1 7085
2 83881 1 7092
2 83882 1 7092
2 83883 1 7092
2 83884 1 7092
2 83885 1 7093
2 83886 1 7093
2 83887 1 7093
2 83888 1 7093
2 83889 1 7093
2 83890 1 7093
2 83891 1 7093
2 83892 1 7093
2 83893 1 7096
2 83894 1 7096
2 83895 1 7096
2 83896 1 7096
2 83897 1 7096
2 83898 1 7096
2 83899 1 7096
2 83900 1 7096
2 83901 1 7096
2 83902 1 7096
2 83903 1 7096
2 83904 1 7096
2 83905 1 7096
2 83906 1 7096
2 83907 1 7096
2 83908 1 7096
2 83909 1 7096
2 83910 1 7096
2 83911 1 7096
2 83912 1 7096
2 83913 1 7096
2 83914 1 7096
2 83915 1 7097
2 83916 1 7097
2 83917 1 7097
2 83918 1 7097
2 83919 1 7097
2 83920 1 7097
2 83921 1 7097
2 83922 1 7097
2 83923 1 7105
2 83924 1 7105
2 83925 1 7105
2 83926 1 7113
2 83927 1 7113
2 83928 1 7114
2 83929 1 7114
2 83930 1 7114
2 83931 1 7115
2 83932 1 7115
2 83933 1 7126
2 83934 1 7126
2 83935 1 7126
2 83936 1 7126
2 83937 1 7126
2 83938 1 7126
2 83939 1 7126
2 83940 1 7126
2 83941 1 7126
2 83942 1 7127
2 83943 1 7127
2 83944 1 7127
2 83945 1 7145
2 83946 1 7145
2 83947 1 7145
2 83948 1 7145
2 83949 1 7145
2 83950 1 7145
2 83951 1 7156
2 83952 1 7156
2 83953 1 7156
2 83954 1 7156
2 83955 1 7159
2 83956 1 7159
2 83957 1 7162
2 83958 1 7162
2 83959 1 7191
2 83960 1 7191
2 83961 1 7192
2 83962 1 7192
2 83963 1 7193
2 83964 1 7193
2 83965 1 7193
2 83966 1 7211
2 83967 1 7211
2 83968 1 7225
2 83969 1 7225
2 83970 1 7260
2 83971 1 7260
2 83972 1 7263
2 83973 1 7263
2 83974 1 7289
2 83975 1 7289
2 83976 1 7299
2 83977 1 7299
2 83978 1 7299
2 83979 1 7299
2 83980 1 7299
2 83981 1 7299
2 83982 1 7299
2 83983 1 7301
2 83984 1 7301
2 83985 1 7302
2 83986 1 7302
2 83987 1 7304
2 83988 1 7304
2 83989 1 7309
2 83990 1 7309
2 83991 1 7312
2 83992 1 7312
2 83993 1 7320
2 83994 1 7320
2 83995 1 7320
2 83996 1 7320
2 83997 1 7322
2 83998 1 7322
2 83999 1 7322
2 84000 1 7333
2 84001 1 7333
2 84002 1 7333
2 84003 1 7333
2 84004 1 7335
2 84005 1 7335
2 84006 1 7336
2 84007 1 7336
2 84008 1 7336
2 84009 1 7339
2 84010 1 7339
2 84011 1 7339
2 84012 1 7339
2 84013 1 7343
2 84014 1 7343
2 84015 1 7343
2 84016 1 7343
2 84017 1 7343
2 84018 1 7344
2 84019 1 7344
2 84020 1 7344
2 84021 1 7344
2 84022 1 7363
2 84023 1 7363
2 84024 1 7373
2 84025 1 7373
2 84026 1 7373
2 84027 1 7373
2 84028 1 7373
2 84029 1 7400
2 84030 1 7400
2 84031 1 7400
2 84032 1 7400
2 84033 1 7401
2 84034 1 7401
2 84035 1 7405
2 84036 1 7405
2 84037 1 7405
2 84038 1 7405
2 84039 1 7414
2 84040 1 7414
2 84041 1 7417
2 84042 1 7417
2 84043 1 7432
2 84044 1 7432
2 84045 1 7432
2 84046 1 7439
2 84047 1 7439
2 84048 1 7439
2 84049 1 7441
2 84050 1 7441
2 84051 1 7442
2 84052 1 7442
2 84053 1 7442
2 84054 1 7442
2 84055 1 7457
2 84056 1 7457
2 84057 1 7462
2 84058 1 7462
2 84059 1 7463
2 84060 1 7463
2 84061 1 7467
2 84062 1 7467
2 84063 1 7491
2 84064 1 7491
2 84065 1 7494
2 84066 1 7494
2 84067 1 7497
2 84068 1 7497
2 84069 1 7497
2 84070 1 7514
2 84071 1 7514
2 84072 1 7514
2 84073 1 7514
2 84074 1 7514
2 84075 1 7516
2 84076 1 7516
2 84077 1 7516
2 84078 1 7516
2 84079 1 7516
2 84080 1 7516
2 84081 1 7516
2 84082 1 7516
2 84083 1 7516
2 84084 1 7516
2 84085 1 7516
2 84086 1 7516
2 84087 1 7517
2 84088 1 7517
2 84089 1 7517
2 84090 1 7517
2 84091 1 7518
2 84092 1 7518
2 84093 1 7524
2 84094 1 7524
2 84095 1 7524
2 84096 1 7525
2 84097 1 7525
2 84098 1 7525
2 84099 1 7525
2 84100 1 7525
2 84101 1 7526
2 84102 1 7526
2 84103 1 7526
2 84104 1 7526
2 84105 1 7526
2 84106 1 7527
2 84107 1 7527
2 84108 1 7530
2 84109 1 7530
2 84110 1 7545
2 84111 1 7545
2 84112 1 7545
2 84113 1 7545
2 84114 1 7545
2 84115 1 7550
2 84116 1 7550
2 84117 1 7556
2 84118 1 7556
2 84119 1 7556
2 84120 1 7557
2 84121 1 7557
2 84122 1 7557
2 84123 1 7557
2 84124 1 7557
2 84125 1 7557
2 84126 1 7573
2 84127 1 7573
2 84128 1 7578
2 84129 1 7578
2 84130 1 7594
2 84131 1 7594
2 84132 1 7604
2 84133 1 7604
2 84134 1 7607
2 84135 1 7607
2 84136 1 7607
2 84137 1 7607
2 84138 1 7607
2 84139 1 7607
2 84140 1 7607
2 84141 1 7607
2 84142 1 7607
2 84143 1 7607
2 84144 1 7607
2 84145 1 7607
2 84146 1 7610
2 84147 1 7610
2 84148 1 7610
2 84149 1 7611
2 84150 1 7611
2 84151 1 7611
2 84152 1 7611
2 84153 1 7611
2 84154 1 7611
2 84155 1 7611
2 84156 1 7612
2 84157 1 7612
2 84158 1 7612
2 84159 1 7612
2 84160 1 7612
2 84161 1 7612
2 84162 1 7620
2 84163 1 7620
2 84164 1 7621
2 84165 1 7621
2 84166 1 7621
2 84167 1 7621
2 84168 1 7621
2 84169 1 7621
2 84170 1 7621
2 84171 1 7621
2 84172 1 7621
2 84173 1 7630
2 84174 1 7630
2 84175 1 7630
2 84176 1 7630
2 84177 1 7630
2 84178 1 7630
2 84179 1 7630
2 84180 1 7630
2 84181 1 7630
2 84182 1 7630
2 84183 1 7630
2 84184 1 7630
2 84185 1 7630
2 84186 1 7630
2 84187 1 7630
2 84188 1 7630
2 84189 1 7630
2 84190 1 7630
2 84191 1 7630
2 84192 1 7630
2 84193 1 7630
2 84194 1 7630
2 84195 1 7630
2 84196 1 7630
2 84197 1 7630
2 84198 1 7630
2 84199 1 7630
2 84200 1 7630
2 84201 1 7630
2 84202 1 7630
2 84203 1 7630
2 84204 1 7630
2 84205 1 7630
2 84206 1 7630
2 84207 1 7630
2 84208 1 7630
2 84209 1 7630
2 84210 1 7630
2 84211 1 7630
2 84212 1 7632
2 84213 1 7632
2 84214 1 7632
2 84215 1 7632
2 84216 1 7632
2 84217 1 7632
2 84218 1 7632
2 84219 1 7632
2 84220 1 7641
2 84221 1 7641
2 84222 1 7641
2 84223 1 7641
2 84224 1 7641
2 84225 1 7641
2 84226 1 7642
2 84227 1 7642
2 84228 1 7643
2 84229 1 7643
2 84230 1 7643
2 84231 1 7643
2 84232 1 7643
2 84233 1 7643
2 84234 1 7643
2 84235 1 7644
2 84236 1 7644
2 84237 1 7644
2 84238 1 7644
2 84239 1 7645
2 84240 1 7645
2 84241 1 7646
2 84242 1 7646
2 84243 1 7646
2 84244 1 7646
2 84245 1 7646
2 84246 1 7647
2 84247 1 7647
2 84248 1 7668
2 84249 1 7668
2 84250 1 7668
2 84251 1 7668
2 84252 1 7668
2 84253 1 7668
2 84254 1 7668
2 84255 1 7668
2 84256 1 7669
2 84257 1 7669
2 84258 1 7669
2 84259 1 7669
2 84260 1 7669
2 84261 1 7669
2 84262 1 7671
2 84263 1 7671
2 84264 1 7671
2 84265 1 7671
2 84266 1 7671
2 84267 1 7671
2 84268 1 7671
2 84269 1 7671
2 84270 1 7671
2 84271 1 7671
2 84272 1 7671
2 84273 1 7672
2 84274 1 7672
2 84275 1 7672
2 84276 1 7680
2 84277 1 7680
2 84278 1 7680
2 84279 1 7680
2 84280 1 7680
2 84281 1 7680
2 84282 1 7682
2 84283 1 7682
2 84284 1 7682
2 84285 1 7682
2 84286 1 7682
2 84287 1 7682
2 84288 1 7682
2 84289 1 7682
2 84290 1 7683
2 84291 1 7683
2 84292 1 7683
2 84293 1 7683
2 84294 1 7683
2 84295 1 7683
2 84296 1 7687
2 84297 1 7687
2 84298 1 7687
2 84299 1 7688
2 84300 1 7688
2 84301 1 7689
2 84302 1 7689
2 84303 1 7689
2 84304 1 7689
2 84305 1 7689
2 84306 1 7689
2 84307 1 7689
2 84308 1 7689
2 84309 1 7691
2 84310 1 7691
2 84311 1 7699
2 84312 1 7699
2 84313 1 7703
2 84314 1 7703
2 84315 1 7703
2 84316 1 7716
2 84317 1 7716
2 84318 1 7724
2 84319 1 7724
2 84320 1 7724
2 84321 1 7735
2 84322 1 7735
2 84323 1 7740
2 84324 1 7740
2 84325 1 7740
2 84326 1 7740
2 84327 1 7740
2 84328 1 7740
2 84329 1 7740
2 84330 1 7740
2 84331 1 7740
2 84332 1 7740
2 84333 1 7740
2 84334 1 7740
2 84335 1 7740
2 84336 1 7740
2 84337 1 7740
2 84338 1 7740
2 84339 1 7740
2 84340 1 7740
2 84341 1 7740
2 84342 1 7740
2 84343 1 7740
2 84344 1 7740
2 84345 1 7740
2 84346 1 7740
2 84347 1 7740
2 84348 1 7740
2 84349 1 7740
2 84350 1 7740
2 84351 1 7740
2 84352 1 7740
2 84353 1 7740
2 84354 1 7740
2 84355 1 7740
2 84356 1 7740
2 84357 1 7740
2 84358 1 7740
2 84359 1 7740
2 84360 1 7740
2 84361 1 7740
2 84362 1 7740
2 84363 1 7740
2 84364 1 7740
2 84365 1 7740
2 84366 1 7740
2 84367 1 7740
2 84368 1 7740
2 84369 1 7740
2 84370 1 7740
2 84371 1 7741
2 84372 1 7741
2 84373 1 7742
2 84374 1 7742
2 84375 1 7742
2 84376 1 7742
2 84377 1 7742
2 84378 1 7742
2 84379 1 7742
2 84380 1 7742
2 84381 1 7742
2 84382 1 7742
2 84383 1 7742
2 84384 1 7742
2 84385 1 7742
2 84386 1 7742
2 84387 1 7742
2 84388 1 7742
2 84389 1 7743
2 84390 1 7743
2 84391 1 7743
2 84392 1 7743
2 84393 1 7744
2 84394 1 7744
2 84395 1 7744
2 84396 1 7758
2 84397 1 7758
2 84398 1 7758
2 84399 1 7759
2 84400 1 7759
2 84401 1 7760
2 84402 1 7760
2 84403 1 7760
2 84404 1 7760
2 84405 1 7761
2 84406 1 7761
2 84407 1 7773
2 84408 1 7773
2 84409 1 7773
2 84410 1 7773
2 84411 1 7773
2 84412 1 7773
2 84413 1 7774
2 84414 1 7774
2 84415 1 7775
2 84416 1 7775
2 84417 1 7775
2 84418 1 7775
2 84419 1 7794
2 84420 1 7794
2 84421 1 7796
2 84422 1 7796
2 84423 1 7796
2 84424 1 7796
2 84425 1 7796
2 84426 1 7796
2 84427 1 7796
2 84428 1 7796
2 84429 1 7796
2 84430 1 7796
2 84431 1 7796
2 84432 1 7796
2 84433 1 7796
2 84434 1 7796
2 84435 1 7796
2 84436 1 7796
2 84437 1 7796
2 84438 1 7796
2 84439 1 7796
2 84440 1 7796
2 84441 1 7796
2 84442 1 7796
2 84443 1 7796
2 84444 1 7796
2 84445 1 7796
2 84446 1 7796
2 84447 1 7796
2 84448 1 7796
2 84449 1 7796
2 84450 1 7796
2 84451 1 7796
2 84452 1 7796
2 84453 1 7796
2 84454 1 7798
2 84455 1 7798
2 84456 1 7801
2 84457 1 7801
2 84458 1 7801
2 84459 1 7801
2 84460 1 7802
2 84461 1 7802
2 84462 1 7802
2 84463 1 7803
2 84464 1 7803
2 84465 1 7812
2 84466 1 7812
2 84467 1 7812
2 84468 1 7812
2 84469 1 7812
2 84470 1 7812
2 84471 1 7812
2 84472 1 7812
2 84473 1 7812
2 84474 1 7812
2 84475 1 7812
2 84476 1 7812
2 84477 1 7812
2 84478 1 7812
2 84479 1 7812
2 84480 1 7812
2 84481 1 7812
2 84482 1 7812
2 84483 1 7812
2 84484 1 7812
2 84485 1 7812
2 84486 1 7812
2 84487 1 7812
2 84488 1 7812
2 84489 1 7812
2 84490 1 7812
2 84491 1 7812
2 84492 1 7812
2 84493 1 7812
2 84494 1 7812
2 84495 1 7812
2 84496 1 7812
2 84497 1 7812
2 84498 1 7812
2 84499 1 7812
2 84500 1 7812
2 84501 1 7812
2 84502 1 7812
2 84503 1 7812
2 84504 1 7812
2 84505 1 7812
2 84506 1 7812
2 84507 1 7812
2 84508 1 7812
2 84509 1 7812
2 84510 1 7812
2 84511 1 7812
2 84512 1 7812
2 84513 1 7812
2 84514 1 7812
2 84515 1 7812
2 84516 1 7812
2 84517 1 7812
2 84518 1 7812
2 84519 1 7812
2 84520 1 7812
2 84521 1 7812
2 84522 1 7812
2 84523 1 7812
2 84524 1 7812
2 84525 1 7812
2 84526 1 7812
2 84527 1 7812
2 84528 1 7812
2 84529 1 7812
2 84530 1 7812
2 84531 1 7812
2 84532 1 7812
2 84533 1 7812
2 84534 1 7812
2 84535 1 7812
2 84536 1 7812
2 84537 1 7812
2 84538 1 7812
2 84539 1 7812
2 84540 1 7812
2 84541 1 7812
2 84542 1 7812
2 84543 1 7813
2 84544 1 7813
2 84545 1 7813
2 84546 1 7813
2 84547 1 7813
2 84548 1 7813
2 84549 1 7813
2 84550 1 7813
2 84551 1 7813
2 84552 1 7813
2 84553 1 7813
2 84554 1 7813
2 84555 1 7813
2 84556 1 7813
2 84557 1 7813
2 84558 1 7813
2 84559 1 7813
2 84560 1 7813
2 84561 1 7813
2 84562 1 7813
2 84563 1 7813
2 84564 1 7813
2 84565 1 7813
2 84566 1 7813
2 84567 1 7813
2 84568 1 7821
2 84569 1 7821
2 84570 1 7822
2 84571 1 7822
2 84572 1 7827
2 84573 1 7827
2 84574 1 7827
2 84575 1 7828
2 84576 1 7828
2 84577 1 7838
2 84578 1 7838
2 84579 1 7838
2 84580 1 7838
2 84581 1 7839
2 84582 1 7839
2 84583 1 7839
2 84584 1 7840
2 84585 1 7840
2 84586 1 7840
2 84587 1 7840
2 84588 1 7840
2 84589 1 7840
2 84590 1 7840
2 84591 1 7840
2 84592 1 7840
2 84593 1 7840
2 84594 1 7841
2 84595 1 7841
2 84596 1 7841
2 84597 1 7841
2 84598 1 7841
2 84599 1 7841
2 84600 1 7841
2 84601 1 7841
2 84602 1 7841
2 84603 1 7841
2 84604 1 7841
2 84605 1 7841
2 84606 1 7841
2 84607 1 7841
2 84608 1 7841
2 84609 1 7841
2 84610 1 7842
2 84611 1 7842
2 84612 1 7842
2 84613 1 7843
2 84614 1 7843
2 84615 1 7843
2 84616 1 7843
2 84617 1 7859
2 84618 1 7859
2 84619 1 7859
2 84620 1 7859
2 84621 1 7859
2 84622 1 7860
2 84623 1 7860
2 84624 1 7861
2 84625 1 7861
2 84626 1 7869
2 84627 1 7869
2 84628 1 7869
2 84629 1 7869
2 84630 1 7869
2 84631 1 7878
2 84632 1 7878
2 84633 1 7878
2 84634 1 7878
2 84635 1 7878
2 84636 1 7878
2 84637 1 7878
2 84638 1 7878
2 84639 1 7882
2 84640 1 7882
2 84641 1 7882
2 84642 1 7882
2 84643 1 7882
2 84644 1 7883
2 84645 1 7883
2 84646 1 7883
2 84647 1 7883
2 84648 1 7883
2 84649 1 7883
2 84650 1 7884
2 84651 1 7884
2 84652 1 7897
2 84653 1 7897
2 84654 1 7897
2 84655 1 7897
2 84656 1 7897
2 84657 1 7897
2 84658 1 7897
2 84659 1 7898
2 84660 1 7898
2 84661 1 7898
2 84662 1 7898
2 84663 1 7898
2 84664 1 7898
2 84665 1 7909
2 84666 1 7909
2 84667 1 7909
2 84668 1 7909
2 84669 1 7910
2 84670 1 7910
2 84671 1 7913
2 84672 1 7913
2 84673 1 7913
2 84674 1 7913
2 84675 1 7922
2 84676 1 7922
2 84677 1 7922
2 84678 1 7931
2 84679 1 7931
2 84680 1 7932
2 84681 1 7932
2 84682 1 7936
2 84683 1 7936
2 84684 1 7936
2 84685 1 7936
2 84686 1 7936
2 84687 1 7936
2 84688 1 7936
2 84689 1 7937
2 84690 1 7937
2 84691 1 7946
2 84692 1 7946
2 84693 1 7946
2 84694 1 7947
2 84695 1 7947
2 84696 1 7947
2 84697 1 7947
2 84698 1 7949
2 84699 1 7949
2 84700 1 7957
2 84701 1 7957
2 84702 1 7968
2 84703 1 7968
2 84704 1 7969
2 84705 1 7969
2 84706 1 7975
2 84707 1 7975
2 84708 1 7978
2 84709 1 7978
2 84710 1 7978
2 84711 1 7978
2 84712 1 7979
2 84713 1 7979
2 84714 1 7980
2 84715 1 7980
2 84716 1 7980
2 84717 1 7980
2 84718 1 7989
2 84719 1 7989
2 84720 1 7991
2 84721 1 7991
2 84722 1 8000
2 84723 1 8000
2 84724 1 8000
2 84725 1 8001
2 84726 1 8001
2 84727 1 8011
2 84728 1 8011
2 84729 1 8011
2 84730 1 8011
2 84731 1 8011
2 84732 1 8011
2 84733 1 8011
2 84734 1 8011
2 84735 1 8011
2 84736 1 8011
2 84737 1 8011
2 84738 1 8011
2 84739 1 8011
2 84740 1 8011
2 84741 1 8011
2 84742 1 8011
2 84743 1 8012
2 84744 1 8012
2 84745 1 8012
2 84746 1 8013
2 84747 1 8013
2 84748 1 8013
2 84749 1 8014
2 84750 1 8014
2 84751 1 8014
2 84752 1 8019
2 84753 1 8019
2 84754 1 8020
2 84755 1 8020
2 84756 1 8020
2 84757 1 8031
2 84758 1 8031
2 84759 1 8033
2 84760 1 8033
2 84761 1 8044
2 84762 1 8044
2 84763 1 8044
2 84764 1 8044
2 84765 1 8044
2 84766 1 8045
2 84767 1 8045
2 84768 1 8045
2 84769 1 8045
2 84770 1 8045
2 84771 1 8045
2 84772 1 8045
2 84773 1 8045
2 84774 1 8045
2 84775 1 8045
2 84776 1 8045
2 84777 1 8045
2 84778 1 8045
2 84779 1 8045
2 84780 1 8045
2 84781 1 8045
2 84782 1 8046
2 84783 1 8046
2 84784 1 8047
2 84785 1 8047
2 84786 1 8048
2 84787 1 8048
2 84788 1 8049
2 84789 1 8049
2 84790 1 8049
2 84791 1 8055
2 84792 1 8055
2 84793 1 8055
2 84794 1 8055
2 84795 1 8061
2 84796 1 8061
2 84797 1 8061
2 84798 1 8061
2 84799 1 8061
2 84800 1 8061
2 84801 1 8061
2 84802 1 8061
2 84803 1 8061
2 84804 1 8061
2 84805 1 8061
2 84806 1 8061
2 84807 1 8061
2 84808 1 8061
2 84809 1 8061
2 84810 1 8061
2 84811 1 8061
2 84812 1 8061
2 84813 1 8062
2 84814 1 8062
2 84815 1 8071
2 84816 1 8071
2 84817 1 8071
2 84818 1 8071
2 84819 1 8071
2 84820 1 8071
2 84821 1 8081
2 84822 1 8081
2 84823 1 8081
2 84824 1 8081
2 84825 1 8081
2 84826 1 8081
2 84827 1 8081
2 84828 1 8081
2 84829 1 8081
2 84830 1 8081
2 84831 1 8081
2 84832 1 8081
2 84833 1 8081
2 84834 1 8081
2 84835 1 8081
2 84836 1 8081
2 84837 1 8081
2 84838 1 8082
2 84839 1 8082
2 84840 1 8082
2 84841 1 8082
2 84842 1 8082
2 84843 1 8083
2 84844 1 8083
2 84845 1 8083
2 84846 1 8083
2 84847 1 8083
2 84848 1 8087
2 84849 1 8087
2 84850 1 8088
2 84851 1 8088
2 84852 1 8089
2 84853 1 8089
2 84854 1 8089
2 84855 1 8089
2 84856 1 8089
2 84857 1 8089
2 84858 1 8089
2 84859 1 8100
2 84860 1 8100
2 84861 1 8104
2 84862 1 8104
2 84863 1 8104
2 84864 1 8104
2 84865 1 8104
2 84866 1 8104
2 84867 1 8104
2 84868 1 8104
2 84869 1 8104
2 84870 1 8104
2 84871 1 8104
2 84872 1 8104
2 84873 1 8104
2 84874 1 8104
2 84875 1 8112
2 84876 1 8112
2 84877 1 8113
2 84878 1 8113
2 84879 1 8113
2 84880 1 8113
2 84881 1 8113
2 84882 1 8113
2 84883 1 8113
2 84884 1 8113
2 84885 1 8113
2 84886 1 8114
2 84887 1 8114
2 84888 1 8114
2 84889 1 8133
2 84890 1 8133
2 84891 1 8133
2 84892 1 8141
2 84893 1 8141
2 84894 1 8141
2 84895 1 8156
2 84896 1 8156
2 84897 1 8160
2 84898 1 8160
2 84899 1 8169
2 84900 1 8169
2 84901 1 8169
2 84902 1 8169
2 84903 1 8169
2 84904 1 8169
2 84905 1 8169
2 84906 1 8169
2 84907 1 8169
2 84908 1 8169
2 84909 1 8170
2 84910 1 8170
2 84911 1 8170
2 84912 1 8170
2 84913 1 8170
2 84914 1 8170
2 84915 1 8170
2 84916 1 8170
2 84917 1 8189
2 84918 1 8189
2 84919 1 8189
2 84920 1 8189
2 84921 1 8191
2 84922 1 8191
2 84923 1 8204
2 84924 1 8204
2 84925 1 8205
2 84926 1 8205
2 84927 1 8205
2 84928 1 8206
2 84929 1 8206
2 84930 1 8206
2 84931 1 8216
2 84932 1 8216
2 84933 1 8216
2 84934 1 8216
2 84935 1 8217
2 84936 1 8217
2 84937 1 8217
2 84938 1 8218
2 84939 1 8218
2 84940 1 8218
2 84941 1 8219
2 84942 1 8219
2 84943 1 8227
2 84944 1 8227
2 84945 1 8227
2 84946 1 8227
2 84947 1 8227
2 84948 1 8227
2 84949 1 8227
2 84950 1 8227
2 84951 1 8227
2 84952 1 8229
2 84953 1 8229
2 84954 1 8229
2 84955 1 8238
2 84956 1 8238
2 84957 1 8247
2 84958 1 8247
2 84959 1 8247
2 84960 1 8247
2 84961 1 8251
2 84962 1 8251
2 84963 1 8251
2 84964 1 8254
2 84965 1 8254
2 84966 1 8258
2 84967 1 8258
2 84968 1 8279
2 84969 1 8279
2 84970 1 8279
2 84971 1 8285
2 84972 1 8285
2 84973 1 8289
2 84974 1 8289
2 84975 1 8290
2 84976 1 8290
2 84977 1 8290
2 84978 1 8290
2 84979 1 8294
2 84980 1 8294
2 84981 1 8295
2 84982 1 8295
2 84983 1 8295
2 84984 1 8295
2 84985 1 8313
2 84986 1 8313
2 84987 1 8313
2 84988 1 8313
2 84989 1 8313
2 84990 1 8314
2 84991 1 8314
2 84992 1 8314
2 84993 1 8316
2 84994 1 8316
2 84995 1 8322
2 84996 1 8322
2 84997 1 8326
2 84998 1 8326
2 84999 1 8327
2 85000 1 8327
2 85001 1 8327
2 85002 1 8327
2 85003 1 8328
2 85004 1 8328
2 85005 1 8328
2 85006 1 8328
2 85007 1 8335
2 85008 1 8335
2 85009 1 8335
2 85010 1 8335
2 85011 1 8335
2 85012 1 8335
2 85013 1 8336
2 85014 1 8336
2 85015 1 8336
2 85016 1 8336
2 85017 1 8336
2 85018 1 8337
2 85019 1 8337
2 85020 1 8340
2 85021 1 8340
2 85022 1 8346
2 85023 1 8346
2 85024 1 8348
2 85025 1 8348
2 85026 1 8365
2 85027 1 8365
2 85028 1 8365
2 85029 1 8368
2 85030 1 8368
2 85031 1 8378
2 85032 1 8378
2 85033 1 8380
2 85034 1 8380
2 85035 1 8380
2 85036 1 8380
2 85037 1 8380
2 85038 1 8380
2 85039 1 8380
2 85040 1 8380
2 85041 1 8380
2 85042 1 8380
2 85043 1 8380
2 85044 1 8380
2 85045 1 8380
2 85046 1 8380
2 85047 1 8380
2 85048 1 8380
2 85049 1 8380
2 85050 1 8381
2 85051 1 8381
2 85052 1 8381
2 85053 1 8381
2 85054 1 8381
2 85055 1 8381
2 85056 1 8382
2 85057 1 8382
2 85058 1 8394
2 85059 1 8394
2 85060 1 8394
2 85061 1 8394
2 85062 1 8394
2 85063 1 8394
2 85064 1 8395
2 85065 1 8395
2 85066 1 8395
2 85067 1 8395
2 85068 1 8401
2 85069 1 8401
2 85070 1 8404
2 85071 1 8404
2 85072 1 8404
2 85073 1 8404
2 85074 1 8405
2 85075 1 8405
2 85076 1 8414
2 85077 1 8414
2 85078 1 8414
2 85079 1 8415
2 85080 1 8415
2 85081 1 8416
2 85082 1 8416
2 85083 1 8416
2 85084 1 8416
2 85085 1 8417
2 85086 1 8417
2 85087 1 8417
2 85088 1 8421
2 85089 1 8421
2 85090 1 8429
2 85091 1 8429
2 85092 1 8429
2 85093 1 8430
2 85094 1 8430
2 85095 1 8430
2 85096 1 8431
2 85097 1 8431
2 85098 1 8431
2 85099 1 8432
2 85100 1 8432
2 85101 1 8442
2 85102 1 8442
2 85103 1 8442
2 85104 1 8458
2 85105 1 8458
2 85106 1 8458
2 85107 1 8458
2 85108 1 8458
2 85109 1 8459
2 85110 1 8459
2 85111 1 8459
2 85112 1 8459
2 85113 1 8459
2 85114 1 8459
2 85115 1 8459
2 85116 1 8475
2 85117 1 8475
2 85118 1 8475
2 85119 1 8490
2 85120 1 8490
2 85121 1 8497
2 85122 1 8497
2 85123 1 8499
2 85124 1 8499
2 85125 1 8500
2 85126 1 8500
2 85127 1 8511
2 85128 1 8511
2 85129 1 8511
2 85130 1 8511
2 85131 1 8511
2 85132 1 8511
2 85133 1 8511
2 85134 1 8511
2 85135 1 8511
2 85136 1 8511
2 85137 1 8511
2 85138 1 8511
2 85139 1 8511
2 85140 1 8511
2 85141 1 8511
2 85142 1 8511
2 85143 1 8511
2 85144 1 8511
2 85145 1 8512
2 85146 1 8512
2 85147 1 8512
2 85148 1 8512
2 85149 1 8512
2 85150 1 8513
2 85151 1 8513
2 85152 1 8513
2 85153 1 8514
2 85154 1 8514
2 85155 1 8514
2 85156 1 8515
2 85157 1 8515
2 85158 1 8517
2 85159 1 8517
2 85160 1 8517
2 85161 1 8520
2 85162 1 8520
2 85163 1 8520
2 85164 1 8545
2 85165 1 8545
2 85166 1 8576
2 85167 1 8576
2 85168 1 8576
2 85169 1 8576
2 85170 1 8577
2 85171 1 8577
2 85172 1 8578
2 85173 1 8578
2 85174 1 8580
2 85175 1 8580
2 85176 1 8580
2 85177 1 8587
2 85178 1 8587
2 85179 1 8587
2 85180 1 8587
2 85181 1 8587
2 85182 1 8587
2 85183 1 8587
2 85184 1 8587
2 85185 1 8587
2 85186 1 8587
2 85187 1 8587
2 85188 1 8587
2 85189 1 8587
2 85190 1 8587
2 85191 1 8587
2 85192 1 8587
2 85193 1 8588
2 85194 1 8588
2 85195 1 8588
2 85196 1 8588
2 85197 1 8588
2 85198 1 8588
2 85199 1 8588
2 85200 1 8588
2 85201 1 8589
2 85202 1 8589
2 85203 1 8590
2 85204 1 8590
2 85205 1 8590
2 85206 1 8590
2 85207 1 8591
2 85208 1 8591
2 85209 1 8595
2 85210 1 8595
2 85211 1 8603
2 85212 1 8603
2 85213 1 8605
2 85214 1 8605
2 85215 1 8605
2 85216 1 8605
2 85217 1 8606
2 85218 1 8606
2 85219 1 8617
2 85220 1 8617
2 85221 1 8617
2 85222 1 8618
2 85223 1 8618
2 85224 1 8620
2 85225 1 8620
2 85226 1 8622
2 85227 1 8622
2 85228 1 8622
2 85229 1 8628
2 85230 1 8628
2 85231 1 8636
2 85232 1 8636
2 85233 1 8636
2 85234 1 8637
2 85235 1 8637
2 85236 1 8641
2 85237 1 8641
2 85238 1 8642
2 85239 1 8642
2 85240 1 8644
2 85241 1 8644
2 85242 1 8644
2 85243 1 8644
2 85244 1 8645
2 85245 1 8645
2 85246 1 8646
2 85247 1 8646
2 85248 1 8646
2 85249 1 8646
2 85250 1 8655
2 85251 1 8655
2 85252 1 8655
2 85253 1 8656
2 85254 1 8656
2 85255 1 8659
2 85256 1 8659
2 85257 1 8664
2 85258 1 8664
2 85259 1 8664
2 85260 1 8664
2 85261 1 8676
2 85262 1 8676
2 85263 1 8680
2 85264 1 8680
2 85265 1 8680
2 85266 1 8681
2 85267 1 8681
2 85268 1 8681
2 85269 1 8700
2 85270 1 8700
2 85271 1 8700
2 85272 1 8700
2 85273 1 8700
2 85274 1 8700
2 85275 1 8713
2 85276 1 8713
2 85277 1 8713
2 85278 1 8714
2 85279 1 8714
2 85280 1 8722
2 85281 1 8722
2 85282 1 8722
2 85283 1 8723
2 85284 1 8723
2 85285 1 8726
2 85286 1 8726
2 85287 1 8742
2 85288 1 8742
2 85289 1 8742
2 85290 1 8743
2 85291 1 8743
2 85292 1 8743
2 85293 1 8743
2 85294 1 8743
2 85295 1 8743
2 85296 1 8743
2 85297 1 8747
2 85298 1 8747
2 85299 1 8747
2 85300 1 8747
2 85301 1 8747
2 85302 1 8747
2 85303 1 8747
2 85304 1 8747
2 85305 1 8747
2 85306 1 8747
2 85307 1 8748
2 85308 1 8748
2 85309 1 8748
2 85310 1 8751
2 85311 1 8751
2 85312 1 8751
2 85313 1 8752
2 85314 1 8752
2 85315 1 8752
2 85316 1 8770
2 85317 1 8770
2 85318 1 8773
2 85319 1 8773
2 85320 1 8773
2 85321 1 8773
2 85322 1 8773
2 85323 1 8773
2 85324 1 8773
2 85325 1 8773
2 85326 1 8773
2 85327 1 8773
2 85328 1 8773
2 85329 1 8774
2 85330 1 8774
2 85331 1 8789
2 85332 1 8789
2 85333 1 8789
2 85334 1 8789
2 85335 1 8794
2 85336 1 8794
2 85337 1 8794
2 85338 1 8795
2 85339 1 8795
2 85340 1 8795
2 85341 1 8795
2 85342 1 8795
2 85343 1 8795
2 85344 1 8795
2 85345 1 8795
2 85346 1 8795
2 85347 1 8795
2 85348 1 8795
2 85349 1 8795
2 85350 1 8795
2 85351 1 8796
2 85352 1 8796
2 85353 1 8796
2 85354 1 8796
2 85355 1 8796
2 85356 1 8798
2 85357 1 8798
2 85358 1 8799
2 85359 1 8799
2 85360 1 8799
2 85361 1 8813
2 85362 1 8813
2 85363 1 8815
2 85364 1 8815
2 85365 1 8815
2 85366 1 8815
2 85367 1 8815
2 85368 1 8815
2 85369 1 8815
2 85370 1 8815
2 85371 1 8818
2 85372 1 8818
2 85373 1 8819
2 85374 1 8819
2 85375 1 8819
2 85376 1 8819
2 85377 1 8819
2 85378 1 8819
2 85379 1 8820
2 85380 1 8820
2 85381 1 8820
2 85382 1 8822
2 85383 1 8822
2 85384 1 8822
2 85385 1 8822
2 85386 1 8822
2 85387 1 8823
2 85388 1 8823
2 85389 1 8831
2 85390 1 8831
2 85391 1 8861
2 85392 1 8861
2 85393 1 8862
2 85394 1 8862
2 85395 1 8862
2 85396 1 8862
2 85397 1 8862
2 85398 1 8869
2 85399 1 8869
2 85400 1 8869
2 85401 1 8869
2 85402 1 8870
2 85403 1 8870
2 85404 1 8870
2 85405 1 8870
2 85406 1 8871
2 85407 1 8871
2 85408 1 8871
2 85409 1 8871
2 85410 1 8871
2 85411 1 8872
2 85412 1 8872
2 85413 1 8880
2 85414 1 8880
2 85415 1 8880
2 85416 1 8883
2 85417 1 8883
2 85418 1 8883
2 85419 1 8883
2 85420 1 8883
2 85421 1 8886
2 85422 1 8886
2 85423 1 8886
2 85424 1 8897
2 85425 1 8897
2 85426 1 8897
2 85427 1 8897
2 85428 1 8897
2 85429 1 8897
2 85430 1 8897
2 85431 1 8898
2 85432 1 8898
2 85433 1 8899
2 85434 1 8899
2 85435 1 8916
2 85436 1 8916
2 85437 1 8941
2 85438 1 8941
2 85439 1 8941
2 85440 1 8941
2 85441 1 8941
2 85442 1 8941
2 85443 1 8941
2 85444 1 8941
2 85445 1 8941
2 85446 1 8941
2 85447 1 8941
2 85448 1 8941
2 85449 1 8941
2 85450 1 8941
2 85451 1 8941
2 85452 1 8941
2 85453 1 8941
2 85454 1 8941
2 85455 1 8941
2 85456 1 8941
2 85457 1 8941
2 85458 1 8942
2 85459 1 8942
2 85460 1 8942
2 85461 1 8942
2 85462 1 8942
2 85463 1 8942
2 85464 1 8943
2 85465 1 8943
2 85466 1 8943
2 85467 1 8943
2 85468 1 8943
2 85469 1 8944
2 85470 1 8944
2 85471 1 8944
2 85472 1 8947
2 85473 1 8947
2 85474 1 8948
2 85475 1 8948
2 85476 1 8951
2 85477 1 8951
2 85478 1 8951
2 85479 1 8951
2 85480 1 8951
2 85481 1 8951
2 85482 1 8952
2 85483 1 8952
2 85484 1 8959
2 85485 1 8959
2 85486 1 8979
2 85487 1 8979
2 85488 1 8979
2 85489 1 8979
2 85490 1 8979
2 85491 1 8979
2 85492 1 8983
2 85493 1 8983
2 85494 1 8986
2 85495 1 8986
2 85496 1 8986
2 85497 1 8987
2 85498 1 8987
2 85499 1 8987
2 85500 1 8987
2 85501 1 8988
2 85502 1 8988
2 85503 1 8988
2 85504 1 8988
2 85505 1 8988
2 85506 1 8988
2 85507 1 8988
2 85508 1 8988
2 85509 1 8988
2 85510 1 8988
2 85511 1 8988
2 85512 1 8988
2 85513 1 8988
2 85514 1 8988
2 85515 1 8988
2 85516 1 8988
2 85517 1 8988
2 85518 1 8988
2 85519 1 8988
2 85520 1 8988
2 85521 1 8988
2 85522 1 8988
2 85523 1 8988
2 85524 1 8988
2 85525 1 8988
2 85526 1 8988
2 85527 1 8988
2 85528 1 8988
2 85529 1 8988
2 85530 1 8988
2 85531 1 8988
2 85532 1 8988
2 85533 1 8988
2 85534 1 8988
2 85535 1 8988
2 85536 1 8988
2 85537 1 8988
2 85538 1 8988
2 85539 1 8988
2 85540 1 8988
2 85541 1 8988
2 85542 1 8988
2 85543 1 8989
2 85544 1 8989
2 85545 1 8989
2 85546 1 8989
2 85547 1 8990
2 85548 1 8990
2 85549 1 8990
2 85550 1 8990
2 85551 1 8990
2 85552 1 8990
2 85553 1 8990
2 85554 1 8990
2 85555 1 8992
2 85556 1 8992
2 85557 1 9011
2 85558 1 9011
2 85559 1 9012
2 85560 1 9012
2 85561 1 9012
2 85562 1 9013
2 85563 1 9013
2 85564 1 9013
2 85565 1 9013
2 85566 1 9013
2 85567 1 9014
2 85568 1 9014
2 85569 1 9014
2 85570 1 9022
2 85571 1 9022
2 85572 1 9040
2 85573 1 9040
2 85574 1 9040
2 85575 1 9050
2 85576 1 9050
2 85577 1 9058
2 85578 1 9058
2 85579 1 9058
2 85580 1 9068
2 85581 1 9068
2 85582 1 9068
2 85583 1 9068
2 85584 1 9069
2 85585 1 9069
2 85586 1 9082
2 85587 1 9082
2 85588 1 9082
2 85589 1 9082
2 85590 1 9083
2 85591 1 9083
2 85592 1 9083
2 85593 1 9083
2 85594 1 9083
2 85595 1 9083
2 85596 1 9083
2 85597 1 9083
2 85598 1 9095
2 85599 1 9095
2 85600 1 9095
2 85601 1 9104
2 85602 1 9104
2 85603 1 9104
2 85604 1 9104
2 85605 1 9104
2 85606 1 9104
2 85607 1 9104
2 85608 1 9104
2 85609 1 9111
2 85610 1 9111
2 85611 1 9113
2 85612 1 9113
2 85613 1 9116
2 85614 1 9116
2 85615 1 9116
2 85616 1 9116
2 85617 1 9117
2 85618 1 9117
2 85619 1 9118
2 85620 1 9118
2 85621 1 9136
2 85622 1 9136
2 85623 1 9136
2 85624 1 9136
2 85625 1 9137
2 85626 1 9137
2 85627 1 9137
2 85628 1 9138
2 85629 1 9138
2 85630 1 9139
2 85631 1 9139
2 85632 1 9141
2 85633 1 9141
2 85634 1 9142
2 85635 1 9142
2 85636 1 9149
2 85637 1 9149
2 85638 1 9151
2 85639 1 9151
2 85640 1 9152
2 85641 1 9152
2 85642 1 9152
2 85643 1 9152
2 85644 1 9152
2 85645 1 9152
2 85646 1 9152
2 85647 1 9154
2 85648 1 9154
2 85649 1 9168
2 85650 1 9168
2 85651 1 9168
2 85652 1 9168
2 85653 1 9169
2 85654 1 9169
2 85655 1 9169
2 85656 1 9175
2 85657 1 9175
2 85658 1 9175
2 85659 1 9175
2 85660 1 9175
2 85661 1 9188
2 85662 1 9188
2 85663 1 9188
2 85664 1 9189
2 85665 1 9189
2 85666 1 9192
2 85667 1 9192
2 85668 1 9192
2 85669 1 9192
2 85670 1 9192
2 85671 1 9192
2 85672 1 9192
2 85673 1 9192
2 85674 1 9192
2 85675 1 9192
2 85676 1 9193
2 85677 1 9193
2 85678 1 9193
2 85679 1 9193
2 85680 1 9193
2 85681 1 9193
2 85682 1 9193
2 85683 1 9193
2 85684 1 9193
2 85685 1 9193
2 85686 1 9193
2 85687 1 9193
2 85688 1 9194
2 85689 1 9194
2 85690 1 9195
2 85691 1 9195
2 85692 1 9195
2 85693 1 9203
2 85694 1 9203
2 85695 1 9203
2 85696 1 9203
2 85697 1 9203
2 85698 1 9203
2 85699 1 9203
2 85700 1 9203
2 85701 1 9203
2 85702 1 9203
2 85703 1 9203
2 85704 1 9203
2 85705 1 9203
2 85706 1 9203
2 85707 1 9203
2 85708 1 9203
2 85709 1 9203
2 85710 1 9203
2 85711 1 9203
2 85712 1 9203
2 85713 1 9203
2 85714 1 9203
2 85715 1 9203
2 85716 1 9203
2 85717 1 9207
2 85718 1 9207
2 85719 1 9227
2 85720 1 9227
2 85721 1 9233
2 85722 1 9233
2 85723 1 9244
2 85724 1 9244
2 85725 1 9244
2 85726 1 9245
2 85727 1 9245
2 85728 1 9247
2 85729 1 9247
2 85730 1 9249
2 85731 1 9249
2 85732 1 9257
2 85733 1 9257
2 85734 1 9264
2 85735 1 9264
2 85736 1 9265
2 85737 1 9265
2 85738 1 9267
2 85739 1 9267
2 85740 1 9268
2 85741 1 9268
2 85742 1 9268
2 85743 1 9268
2 85744 1 9268
2 85745 1 9275
2 85746 1 9275
2 85747 1 9302
2 85748 1 9302
2 85749 1 9303
2 85750 1 9303
2 85751 1 9303
2 85752 1 9313
2 85753 1 9313
2 85754 1 9314
2 85755 1 9314
2 85756 1 9314
2 85757 1 9314
2 85758 1 9314
2 85759 1 9321
2 85760 1 9321
2 85761 1 9321
2 85762 1 9322
2 85763 1 9322
2 85764 1 9329
2 85765 1 9329
2 85766 1 9336
2 85767 1 9336
2 85768 1 9336
2 85769 1 9336
2 85770 1 9339
2 85771 1 9339
2 85772 1 9339
2 85773 1 9340
2 85774 1 9340
2 85775 1 9340
2 85776 1 9340
2 85777 1 9340
2 85778 1 9340
2 85779 1 9340
2 85780 1 9340
2 85781 1 9356
2 85782 1 9356
2 85783 1 9356
2 85784 1 9356
2 85785 1 9356
2 85786 1 9356
2 85787 1 9369
2 85788 1 9369
2 85789 1 9378
2 85790 1 9378
2 85791 1 9378
2 85792 1 9378
2 85793 1 9378
2 85794 1 9378
2 85795 1 9384
2 85796 1 9384
2 85797 1 9384
2 85798 1 9384
2 85799 1 9389
2 85800 1 9389
2 85801 1 9389
2 85802 1 9402
2 85803 1 9402
2 85804 1 9402
2 85805 1 9403
2 85806 1 9403
2 85807 1 9403
2 85808 1 9403
2 85809 1 9404
2 85810 1 9404
2 85811 1 9404
2 85812 1 9405
2 85813 1 9405
2 85814 1 9405
2 85815 1 9405
2 85816 1 9405
2 85817 1 9405
2 85818 1 9405
2 85819 1 9405
2 85820 1 9406
2 85821 1 9406
2 85822 1 9406
2 85823 1 9407
2 85824 1 9407
2 85825 1 9408
2 85826 1 9408
2 85827 1 9408
2 85828 1 9408
2 85829 1 9424
2 85830 1 9424
2 85831 1 9424
2 85832 1 9424
2 85833 1 9426
2 85834 1 9426
2 85835 1 9426
2 85836 1 9427
2 85837 1 9427
2 85838 1 9427
2 85839 1 9427
2 85840 1 9427
2 85841 1 9427
2 85842 1 9427
2 85843 1 9427
2 85844 1 9427
2 85845 1 9427
2 85846 1 9427
2 85847 1 9427
2 85848 1 9427
2 85849 1 9427
2 85850 1 9427
2 85851 1 9427
2 85852 1 9427
2 85853 1 9427
2 85854 1 9427
2 85855 1 9427
2 85856 1 9427
2 85857 1 9428
2 85858 1 9428
2 85859 1 9428
2 85860 1 9429
2 85861 1 9429
2 85862 1 9429
2 85863 1 9430
2 85864 1 9430
2 85865 1 9439
2 85866 1 9439
2 85867 1 9439
2 85868 1 9439
2 85869 1 9440
2 85870 1 9440
2 85871 1 9440
2 85872 1 9440
2 85873 1 9440
2 85874 1 9441
2 85875 1 9441
2 85876 1 9441
2 85877 1 9455
2 85878 1 9455
2 85879 1 9455
2 85880 1 9455
2 85881 1 9455
2 85882 1 9455
2 85883 1 9455
2 85884 1 9455
2 85885 1 9456
2 85886 1 9456
2 85887 1 9456
2 85888 1 9458
2 85889 1 9458
2 85890 1 9458
2 85891 1 9462
2 85892 1 9462
2 85893 1 9463
2 85894 1 9463
2 85895 1 9463
2 85896 1 9463
2 85897 1 9463
2 85898 1 9463
2 85899 1 9463
2 85900 1 9463
2 85901 1 9463
2 85902 1 9463
2 85903 1 9463
2 85904 1 9463
2 85905 1 9463
2 85906 1 9463
2 85907 1 9463
2 85908 1 9463
2 85909 1 9463
2 85910 1 9463
2 85911 1 9463
2 85912 1 9463
2 85913 1 9463
2 85914 1 9463
2 85915 1 9463
2 85916 1 9463
2 85917 1 9463
2 85918 1 9463
2 85919 1 9463
2 85920 1 9463
2 85921 1 9463
2 85922 1 9463
2 85923 1 9463
2 85924 1 9463
2 85925 1 9464
2 85926 1 9464
2 85927 1 9464
2 85928 1 9464
2 85929 1 9464
2 85930 1 9464
2 85931 1 9464
2 85932 1 9464
2 85933 1 9464
2 85934 1 9464
2 85935 1 9477
2 85936 1 9477
2 85937 1 9478
2 85938 1 9478
2 85939 1 9490
2 85940 1 9490
2 85941 1 9490
2 85942 1 9490
2 85943 1 9490
2 85944 1 9490
2 85945 1 9490
2 85946 1 9490
2 85947 1 9490
2 85948 1 9490
2 85949 1 9490
2 85950 1 9491
2 85951 1 9491
2 85952 1 9491
2 85953 1 9491
2 85954 1 9491
2 85955 1 9491
2 85956 1 9491
2 85957 1 9495
2 85958 1 9495
2 85959 1 9496
2 85960 1 9496
2 85961 1 9496
2 85962 1 9498
2 85963 1 9498
2 85964 1 9507
2 85965 1 9507
2 85966 1 9507
2 85967 1 9507
2 85968 1 9508
2 85969 1 9508
2 85970 1 9508
2 85971 1 9508
2 85972 1 9509
2 85973 1 9509
2 85974 1 9510
2 85975 1 9510
2 85976 1 9510
2 85977 1 9510
2 85978 1 9510
2 85979 1 9513
2 85980 1 9513
2 85981 1 9531
2 85982 1 9531
2 85983 1 9531
2 85984 1 9531
2 85985 1 9532
2 85986 1 9532
2 85987 1 9534
2 85988 1 9534
2 85989 1 9535
2 85990 1 9535
2 85991 1 9535
2 85992 1 9536
2 85993 1 9536
2 85994 1 9536
2 85995 1 9537
2 85996 1 9537
2 85997 1 9538
2 85998 1 9538
2 85999 1 9539
2 86000 1 9539
2 86001 1 9539
2 86002 1 9539
2 86003 1 9540
2 86004 1 9540
2 86005 1 9548
2 86006 1 9548
2 86007 1 9549
2 86008 1 9549
2 86009 1 9549
2 86010 1 9549
2 86011 1 9549
2 86012 1 9549
2 86013 1 9550
2 86014 1 9550
2 86015 1 9550
2 86016 1 9550
2 86017 1 9550
2 86018 1 9550
2 86019 1 9554
2 86020 1 9554
2 86021 1 9562
2 86022 1 9562
2 86023 1 9562
2 86024 1 9562
2 86025 1 9563
2 86026 1 9563
2 86027 1 9563
2 86028 1 9564
2 86029 1 9564
2 86030 1 9565
2 86031 1 9565
2 86032 1 9565
2 86033 1 9565
2 86034 1 9585
2 86035 1 9585
2 86036 1 9585
2 86037 1 9585
2 86038 1 9585
2 86039 1 9592
2 86040 1 9592
2 86041 1 9592
2 86042 1 9597
2 86043 1 9597
2 86044 1 9597
2 86045 1 9611
2 86046 1 9611
2 86047 1 9613
2 86048 1 9613
2 86049 1 9613
2 86050 1 9613
2 86051 1 9617
2 86052 1 9617
2 86053 1 9636
2 86054 1 9636
2 86055 1 9636
2 86056 1 9636
2 86057 1 9636
2 86058 1 9636
2 86059 1 9636
2 86060 1 9637
2 86061 1 9637
2 86062 1 9637
2 86063 1 9637
2 86064 1 9637
2 86065 1 9638
2 86066 1 9638
2 86067 1 9638
2 86068 1 9639
2 86069 1 9639
2 86070 1 9646
2 86071 1 9646
2 86072 1 9646
2 86073 1 9646
2 86074 1 9646
2 86075 1 9646
2 86076 1 9646
2 86077 1 9646
2 86078 1 9646
2 86079 1 9646
2 86080 1 9646
2 86081 1 9646
2 86082 1 9646
2 86083 1 9646
2 86084 1 9646
2 86085 1 9646
2 86086 1 9646
2 86087 1 9646
2 86088 1 9646
2 86089 1 9646
2 86090 1 9646
2 86091 1 9646
2 86092 1 9646
2 86093 1 9646
2 86094 1 9646
2 86095 1 9646
2 86096 1 9646
2 86097 1 9646
2 86098 1 9646
2 86099 1 9646
2 86100 1 9646
2 86101 1 9646
2 86102 1 9646
2 86103 1 9646
2 86104 1 9646
2 86105 1 9646
2 86106 1 9646
2 86107 1 9646
2 86108 1 9646
2 86109 1 9646
2 86110 1 9646
2 86111 1 9646
2 86112 1 9646
2 86113 1 9646
2 86114 1 9646
2 86115 1 9646
2 86116 1 9646
2 86117 1 9646
2 86118 1 9647
2 86119 1 9647
2 86120 1 9647
2 86121 1 9647
2 86122 1 9647
2 86123 1 9647
2 86124 1 9647
2 86125 1 9647
2 86126 1 9649
2 86127 1 9649
2 86128 1 9650
2 86129 1 9650
2 86130 1 9650
2 86131 1 9650
2 86132 1 9650
2 86133 1 9651
2 86134 1 9651
2 86135 1 9651
2 86136 1 9651
2 86137 1 9660
2 86138 1 9660
2 86139 1 9660
2 86140 1 9672
2 86141 1 9672
2 86142 1 9672
2 86143 1 9672
2 86144 1 9672
2 86145 1 9672
2 86146 1 9672
2 86147 1 9673
2 86148 1 9673
2 86149 1 9673
2 86150 1 9694
2 86151 1 9694
2 86152 1 9694
2 86153 1 9694
2 86154 1 9694
2 86155 1 9694
2 86156 1 9694
2 86157 1 9694
2 86158 1 9694
2 86159 1 9694
2 86160 1 9694
2 86161 1 9694
2 86162 1 9694
2 86163 1 9694
2 86164 1 9694
2 86165 1 9694
2 86166 1 9694
2 86167 1 9694
2 86168 1 9694
2 86169 1 9694
2 86170 1 9694
2 86171 1 9694
2 86172 1 9694
2 86173 1 9694
2 86174 1 9694
2 86175 1 9694
2 86176 1 9694
2 86177 1 9694
2 86178 1 9694
2 86179 1 9694
2 86180 1 9694
2 86181 1 9694
2 86182 1 9694
2 86183 1 9694
2 86184 1 9694
2 86185 1 9694
2 86186 1 9694
2 86187 1 9694
2 86188 1 9694
2 86189 1 9694
2 86190 1 9694
2 86191 1 9694
2 86192 1 9694
2 86193 1 9694
2 86194 1 9707
2 86195 1 9707
2 86196 1 9707
2 86197 1 9709
2 86198 1 9709
2 86199 1 9709
2 86200 1 9709
2 86201 1 9713
2 86202 1 9713
2 86203 1 9713
2 86204 1 9713
2 86205 1 9713
2 86206 1 9716
2 86207 1 9716
2 86208 1 9716
2 86209 1 9716
2 86210 1 9716
2 86211 1 9716
2 86212 1 9716
2 86213 1 9716
2 86214 1 9716
2 86215 1 9716
2 86216 1 9717
2 86217 1 9717
2 86218 1 9717
2 86219 1 9724
2 86220 1 9724
2 86221 1 9724
2 86222 1 9724
2 86223 1 9724
2 86224 1 9725
2 86225 1 9725
2 86226 1 9725
2 86227 1 9738
2 86228 1 9738
2 86229 1 9740
2 86230 1 9740
2 86231 1 9740
2 86232 1 9740
2 86233 1 9740
2 86234 1 9740
2 86235 1 9740
2 86236 1 9740
2 86237 1 9741
2 86238 1 9741
2 86239 1 9741
2 86240 1 9741
2 86241 1 9741
2 86242 1 9741
2 86243 1 9741
2 86244 1 9741
2 86245 1 9743
2 86246 1 9743
2 86247 1 9743
2 86248 1 9745
2 86249 1 9745
2 86250 1 9745
2 86251 1 9746
2 86252 1 9746
2 86253 1 9753
2 86254 1 9753
2 86255 1 9753
2 86256 1 9753
2 86257 1 9753
2 86258 1 9753
2 86259 1 9753
2 86260 1 9753
2 86261 1 9753
2 86262 1 9753
2 86263 1 9753
2 86264 1 9753
2 86265 1 9754
2 86266 1 9754
2 86267 1 9754
2 86268 1 9767
2 86269 1 9767
2 86270 1 9767
2 86271 1 9769
2 86272 1 9769
2 86273 1 9778
2 86274 1 9778
2 86275 1 9794
2 86276 1 9794
2 86277 1 9794
2 86278 1 9794
2 86279 1 9794
2 86280 1 9794
2 86281 1 9794
2 86282 1 9794
2 86283 1 9794
2 86284 1 9794
2 86285 1 9794
2 86286 1 9794
2 86287 1 9802
2 86288 1 9802
2 86289 1 9802
2 86290 1 9802
2 86291 1 9802
2 86292 1 9802
2 86293 1 9803
2 86294 1 9803
2 86295 1 9804
2 86296 1 9804
2 86297 1 9804
2 86298 1 9807
2 86299 1 9807
2 86300 1 9807
2 86301 1 9807
2 86302 1 9807
2 86303 1 9807
2 86304 1 9807
2 86305 1 9807
2 86306 1 9807
2 86307 1 9807
2 86308 1 9807
2 86309 1 9812
2 86310 1 9812
2 86311 1 9812
2 86312 1 9812
2 86313 1 9812
2 86314 1 9812
2 86315 1 9812
2 86316 1 9812
2 86317 1 9812
2 86318 1 9813
2 86319 1 9813
2 86320 1 9813
2 86321 1 9822
2 86322 1 9822
2 86323 1 9822
2 86324 1 9822
2 86325 1 9822
2 86326 1 9822
2 86327 1 9822
2 86328 1 9822
2 86329 1 9823
2 86330 1 9823
2 86331 1 9823
2 86332 1 9823
2 86333 1 9824
2 86334 1 9824
2 86335 1 9825
2 86336 1 9825
2 86337 1 9832
2 86338 1 9832
2 86339 1 9832
2 86340 1 9832
2 86341 1 9832
2 86342 1 9835
2 86343 1 9835
2 86344 1 9836
2 86345 1 9836
2 86346 1 9836
2 86347 1 9857
2 86348 1 9857
2 86349 1 9857
2 86350 1 9858
2 86351 1 9858
2 86352 1 9858
2 86353 1 9858
2 86354 1 9858
2 86355 1 9858
2 86356 1 9858
2 86357 1 9858
2 86358 1 9858
2 86359 1 9858
2 86360 1 9869
2 86361 1 9869
2 86362 1 9869
2 86363 1 9869
2 86364 1 9869
2 86365 1 9869
2 86366 1 9870
2 86367 1 9870
2 86368 1 9877
2 86369 1 9877
2 86370 1 9877
2 86371 1 9877
2 86372 1 9877
2 86373 1 9877
2 86374 1 9877
2 86375 1 9878
2 86376 1 9878
2 86377 1 9878
2 86378 1 9878
2 86379 1 9887
2 86380 1 9887
2 86381 1 9887
2 86382 1 9887
2 86383 1 9887
2 86384 1 9887
2 86385 1 9887
2 86386 1 9887
2 86387 1 9887
2 86388 1 9887
2 86389 1 9891
2 86390 1 9891
2 86391 1 9891
2 86392 1 9891
2 86393 1 9891
2 86394 1 9926
2 86395 1 9926
2 86396 1 9927
2 86397 1 9927
2 86398 1 9927
2 86399 1 9927
2 86400 1 9927
2 86401 1 9927
2 86402 1 9927
2 86403 1 9927
2 86404 1 9935
2 86405 1 9935
2 86406 1 9935
2 86407 1 9935
2 86408 1 9936
2 86409 1 9936
2 86410 1 9944
2 86411 1 9944
2 86412 1 9944
2 86413 1 9944
2 86414 1 9944
2 86415 1 9944
2 86416 1 9948
2 86417 1 9948
2 86418 1 9951
2 86419 1 9951
2 86420 1 9951
2 86421 1 9951
2 86422 1 9951
2 86423 1 9951
2 86424 1 9951
2 86425 1 9951
2 86426 1 9955
2 86427 1 9955
2 86428 1 9971
2 86429 1 9971
2 86430 1 9971
2 86431 1 9971
2 86432 1 9971
2 86433 1 9971
2 86434 1 9971
2 86435 1 9971
2 86436 1 9971
2 86437 1 9971
2 86438 1 9973
2 86439 1 9973
2 86440 1 9996
2 86441 1 9996
2 86442 1 9996
2 86443 1 9997
2 86444 1 9997
2 86445 1 9997
2 86446 1 10009
2 86447 1 10009
2 86448 1 10012
2 86449 1 10012
2 86450 1 10012
2 86451 1 10013
2 86452 1 10013
2 86453 1 10013
2 86454 1 10013
2 86455 1 10013
2 86456 1 10013
2 86457 1 10013
2 86458 1 10014
2 86459 1 10014
2 86460 1 10021
2 86461 1 10021
2 86462 1 10021
2 86463 1 10021
2 86464 1 10035
2 86465 1 10035
2 86466 1 10035
2 86467 1 10035
2 86468 1 10035
2 86469 1 10035
2 86470 1 10035
2 86471 1 10035
2 86472 1 10035
2 86473 1 10035
2 86474 1 10035
2 86475 1 10035
2 86476 1 10035
2 86477 1 10035
2 86478 1 10035
2 86479 1 10035
2 86480 1 10036
2 86481 1 10036
2 86482 1 10037
2 86483 1 10037
2 86484 1 10037
2 86485 1 10037
2 86486 1 10060
2 86487 1 10060
2 86488 1 10071
2 86489 1 10071
2 86490 1 10071
2 86491 1 10072
2 86492 1 10072
2 86493 1 10072
2 86494 1 10072
2 86495 1 10072
2 86496 1 10072
2 86497 1 10086
2 86498 1 10086
2 86499 1 10087
2 86500 1 10087
2 86501 1 10087
2 86502 1 10087
2 86503 1 10087
2 86504 1 10087
2 86505 1 10087
2 86506 1 10087
2 86507 1 10112
2 86508 1 10112
2 86509 1 10112
2 86510 1 10113
2 86511 1 10113
2 86512 1 10113
2 86513 1 10113
2 86514 1 10113
2 86515 1 10113
2 86516 1 10113
2 86517 1 10114
2 86518 1 10114
2 86519 1 10114
2 86520 1 10114
2 86521 1 10118
2 86522 1 10118
2 86523 1 10134
2 86524 1 10134
2 86525 1 10134
2 86526 1 10135
2 86527 1 10135
2 86528 1 10136
2 86529 1 10136
2 86530 1 10136
2 86531 1 10136
2 86532 1 10136
2 86533 1 10136
2 86534 1 10145
2 86535 1 10145
2 86536 1 10145
2 86537 1 10145
2 86538 1 10145
2 86539 1 10155
2 86540 1 10155
2 86541 1 10155
2 86542 1 10155
2 86543 1 10155
2 86544 1 10165
2 86545 1 10165
2 86546 1 10165
2 86547 1 10165
2 86548 1 10165
2 86549 1 10166
2 86550 1 10166
2 86551 1 10166
2 86552 1 10166
2 86553 1 10166
2 86554 1 10186
2 86555 1 10186
2 86556 1 10186
2 86557 1 10186
2 86558 1 10196
2 86559 1 10196
2 86560 1 10197
2 86561 1 10197
2 86562 1 10197
2 86563 1 10197
2 86564 1 10197
2 86565 1 10198
2 86566 1 10198
2 86567 1 10203
2 86568 1 10203
2 86569 1 10204
2 86570 1 10204
2 86571 1 10204
2 86572 1 10204
2 86573 1 10204
2 86574 1 10204
2 86575 1 10205
2 86576 1 10205
2 86577 1 10205
2 86578 1 10213
2 86579 1 10213
2 86580 1 10213
2 86581 1 10213
2 86582 1 10213
2 86583 1 10213
2 86584 1 10214
2 86585 1 10214
2 86586 1 10214
2 86587 1 10218
2 86588 1 10218
2 86589 1 10228
2 86590 1 10228
2 86591 1 10228
2 86592 1 10228
2 86593 1 10228
2 86594 1 10228
2 86595 1 10228
2 86596 1 10228
2 86597 1 10234
2 86598 1 10234
2 86599 1 10234
2 86600 1 10234
2 86601 1 10234
2 86602 1 10234
2 86603 1 10234
2 86604 1 10234
2 86605 1 10235
2 86606 1 10235
2 86607 1 10243
2 86608 1 10243
2 86609 1 10243
2 86610 1 10243
2 86611 1 10243
2 86612 1 10243
2 86613 1 10244
2 86614 1 10244
2 86615 1 10244
2 86616 1 10244
2 86617 1 10252
2 86618 1 10252
2 86619 1 10252
2 86620 1 10263
2 86621 1 10263
2 86622 1 10263
2 86623 1 10263
2 86624 1 10263
2 86625 1 10263
2 86626 1 10264
2 86627 1 10264
2 86628 1 10265
2 86629 1 10265
2 86630 1 10272
2 86631 1 10272
2 86632 1 10274
2 86633 1 10274
2 86634 1 10277
2 86635 1 10277
2 86636 1 10277
2 86637 1 10285
2 86638 1 10285
2 86639 1 10285
2 86640 1 10286
2 86641 1 10286
2 86642 1 10286
2 86643 1 10286
2 86644 1 10286
2 86645 1 10289
2 86646 1 10289
2 86647 1 10289
2 86648 1 10289
2 86649 1 10332
2 86650 1 10332
2 86651 1 10332
2 86652 1 10332
2 86653 1 10332
2 86654 1 10332
2 86655 1 10332
2 86656 1 10332
2 86657 1 10332
2 86658 1 10332
2 86659 1 10332
2 86660 1 10333
2 86661 1 10333
2 86662 1 10333
2 86663 1 10333
2 86664 1 10333
2 86665 1 10333
2 86666 1 10333
2 86667 1 10335
2 86668 1 10335
2 86669 1 10335
2 86670 1 10336
2 86671 1 10336
2 86672 1 10342
2 86673 1 10342
2 86674 1 10342
2 86675 1 10342
2 86676 1 10342
2 86677 1 10342
2 86678 1 10342
2 86679 1 10342
2 86680 1 10343
2 86681 1 10343
2 86682 1 10346
2 86683 1 10346
2 86684 1 10347
2 86685 1 10347
2 86686 1 10347
2 86687 1 10347
2 86688 1 10347
2 86689 1 10356
2 86690 1 10356
2 86691 1 10356
2 86692 1 10356
2 86693 1 10356
2 86694 1 10357
2 86695 1 10357
2 86696 1 10357
2 86697 1 10382
2 86698 1 10382
2 86699 1 10382
2 86700 1 10382
2 86701 1 10382
2 86702 1 10382
2 86703 1 10382
2 86704 1 10382
2 86705 1 10382
2 86706 1 10382
2 86707 1 10382
2 86708 1 10382
2 86709 1 10382
2 86710 1 10382
2 86711 1 10382
2 86712 1 10382
2 86713 1 10382
2 86714 1 10382
2 86715 1 10382
2 86716 1 10382
2 86717 1 10382
2 86718 1 10382
2 86719 1 10382
2 86720 1 10382
2 86721 1 10382
2 86722 1 10382
2 86723 1 10382
2 86724 1 10382
2 86725 1 10382
2 86726 1 10382
2 86727 1 10382
2 86728 1 10382
2 86729 1 10382
2 86730 1 10382
2 86731 1 10382
2 86732 1 10382
2 86733 1 10382
2 86734 1 10383
2 86735 1 10383
2 86736 1 10383
2 86737 1 10383
2 86738 1 10383
2 86739 1 10383
2 86740 1 10383
2 86741 1 10383
2 86742 1 10383
2 86743 1 10384
2 86744 1 10384
2 86745 1 10384
2 86746 1 10384
2 86747 1 10384
2 86748 1 10384
2 86749 1 10384
2 86750 1 10384
2 86751 1 10384
2 86752 1 10384
2 86753 1 10384
2 86754 1 10384
2 86755 1 10384
2 86756 1 10384
2 86757 1 10384
2 86758 1 10384
2 86759 1 10384
2 86760 1 10384
2 86761 1 10384
2 86762 1 10384
2 86763 1 10384
2 86764 1 10384
2 86765 1 10384
2 86766 1 10384
2 86767 1 10384
2 86768 1 10384
2 86769 1 10385
2 86770 1 10385
2 86771 1 10385
2 86772 1 10385
2 86773 1 10385
2 86774 1 10386
2 86775 1 10386
2 86776 1 10386
2 86777 1 10386
2 86778 1 10386
2 86779 1 10386
2 86780 1 10386
2 86781 1 10386
2 86782 1 10386
2 86783 1 10386
2 86784 1 10386
2 86785 1 10386
2 86786 1 10386
2 86787 1 10386
2 86788 1 10386
2 86789 1 10386
2 86790 1 10386
2 86791 1 10386
2 86792 1 10386
2 86793 1 10386
2 86794 1 10386
2 86795 1 10386
2 86796 1 10386
2 86797 1 10386
2 86798 1 10386
2 86799 1 10386
2 86800 1 10386
2 86801 1 10386
2 86802 1 10386
2 86803 1 10386
2 86804 1 10386
2 86805 1 10386
2 86806 1 10386
2 86807 1 10386
2 86808 1 10386
2 86809 1 10386
2 86810 1 10386
2 86811 1 10386
2 86812 1 10386
2 86813 1 10386
2 86814 1 10386
2 86815 1 10386
2 86816 1 10386
2 86817 1 10386
2 86818 1 10386
2 86819 1 10386
2 86820 1 10386
2 86821 1 10386
2 86822 1 10386
2 86823 1 10387
2 86824 1 10387
2 86825 1 10387
2 86826 1 10388
2 86827 1 10388
2 86828 1 10388
2 86829 1 10388
2 86830 1 10388
2 86831 1 10388
2 86832 1 10388
2 86833 1 10388
2 86834 1 10388
2 86835 1 10388
2 86836 1 10388
2 86837 1 10388
2 86838 1 10388
2 86839 1 10388
2 86840 1 10388
2 86841 1 10389
2 86842 1 10389
2 86843 1 10389
2 86844 1 10389
2 86845 1 10390
2 86846 1 10390
2 86847 1 10393
2 86848 1 10393
2 86849 1 10393
2 86850 1 10393
2 86851 1 10393
2 86852 1 10393
2 86853 1 10401
2 86854 1 10401
2 86855 1 10402
2 86856 1 10402
2 86857 1 10402
2 86858 1 10402
2 86859 1 10402
2 86860 1 10402
2 86861 1 10402
2 86862 1 10410
2 86863 1 10410
2 86864 1 10410
2 86865 1 10410
2 86866 1 10411
2 86867 1 10411
2 86868 1 10411
2 86869 1 10411
2 86870 1 10411
2 86871 1 10420
2 86872 1 10420
2 86873 1 10421
2 86874 1 10421
2 86875 1 10421
2 86876 1 10421
2 86877 1 10421
2 86878 1 10421
2 86879 1 10430
2 86880 1 10430
2 86881 1 10430
2 86882 1 10431
2 86883 1 10431
2 86884 1 10431
2 86885 1 10432
2 86886 1 10432
2 86887 1 10440
2 86888 1 10440
2 86889 1 10440
2 86890 1 10440
2 86891 1 10441
2 86892 1 10441
2 86893 1 10452
2 86894 1 10452
2 86895 1 10452
2 86896 1 10464
2 86897 1 10464
2 86898 1 10464
2 86899 1 10464
2 86900 1 10464
2 86901 1 10465
2 86902 1 10465
2 86903 1 10465
2 86904 1 10465
2 86905 1 10477
2 86906 1 10477
2 86907 1 10477
2 86908 1 10477
2 86909 1 10477
2 86910 1 10477
2 86911 1 10477
2 86912 1 10477
2 86913 1 10477
2 86914 1 10477
2 86915 1 10478
2 86916 1 10478
2 86917 1 10478
2 86918 1 10479
2 86919 1 10479
2 86920 1 10492
2 86921 1 10492
2 86922 1 10492
2 86923 1 10492
2 86924 1 10513
2 86925 1 10513
2 86926 1 10522
2 86927 1 10522
2 86928 1 10522
2 86929 1 10523
2 86930 1 10523
2 86931 1 10539
2 86932 1 10539
2 86933 1 10539
2 86934 1 10539
2 86935 1 10539
2 86936 1 10539
2 86937 1 10539
2 86938 1 10539
2 86939 1 10540
2 86940 1 10540
2 86941 1 10548
2 86942 1 10548
2 86943 1 10554
2 86944 1 10554
2 86945 1 10570
2 86946 1 10570
2 86947 1 10570
2 86948 1 10570
2 86949 1 10570
2 86950 1 10571
2 86951 1 10571
2 86952 1 10572
2 86953 1 10572
2 86954 1 10582
2 86955 1 10582
2 86956 1 10583
2 86957 1 10583
2 86958 1 10583
2 86959 1 10584
2 86960 1 10584
2 86961 1 10605
2 86962 1 10605
2 86963 1 10605
2 86964 1 10605
2 86965 1 10605
2 86966 1 10605
2 86967 1 10605
2 86968 1 10611
2 86969 1 10611
2 86970 1 10611
2 86971 1 10611
2 86972 1 10611
2 86973 1 10611
2 86974 1 10611
2 86975 1 10611
2 86976 1 10611
2 86977 1 10611
2 86978 1 10611
2 86979 1 10611
2 86980 1 10611
2 86981 1 10612
2 86982 1 10612
2 86983 1 10612
2 86984 1 10612
2 86985 1 10612
2 86986 1 10612
2 86987 1 10613
2 86988 1 10613
2 86989 1 10613
2 86990 1 10613
2 86991 1 10613
2 86992 1 10614
2 86993 1 10614
2 86994 1 10614
2 86995 1 10614
2 86996 1 10614
2 86997 1 10614
2 86998 1 10614
2 86999 1 10614
2 87000 1 10614
2 87001 1 10615
2 87002 1 10615
2 87003 1 10615
2 87004 1 10615
2 87005 1 10621
2 87006 1 10621
2 87007 1 10622
2 87008 1 10622
2 87009 1 10622
2 87010 1 10624
2 87011 1 10624
2 87012 1 10637
2 87013 1 10637
2 87014 1 10643
2 87015 1 10643
2 87016 1 10643
2 87017 1 10643
2 87018 1 10643
2 87019 1 10643
2 87020 1 10643
2 87021 1 10643
2 87022 1 10643
2 87023 1 10653
2 87024 1 10653
2 87025 1 10653
2 87026 1 10653
2 87027 1 10653
2 87028 1 10653
2 87029 1 10653
2 87030 1 10653
2 87031 1 10653
2 87032 1 10653
2 87033 1 10654
2 87034 1 10654
2 87035 1 10654
2 87036 1 10654
2 87037 1 10654
2 87038 1 10657
2 87039 1 10657
2 87040 1 10658
2 87041 1 10658
2 87042 1 10666
2 87043 1 10666
2 87044 1 10666
2 87045 1 10666
2 87046 1 10666
2 87047 1 10668
2 87048 1 10668
2 87049 1 10668
2 87050 1 10669
2 87051 1 10669
2 87052 1 10669
2 87053 1 10670
2 87054 1 10670
2 87055 1 10671
2 87056 1 10671
2 87057 1 10671
2 87058 1 10686
2 87059 1 10686
2 87060 1 10689
2 87061 1 10689
2 87062 1 10706
2 87063 1 10706
2 87064 1 10720
2 87065 1 10720
2 87066 1 10720
2 87067 1 10720
2 87068 1 10720
2 87069 1 10720
2 87070 1 10720
2 87071 1 10720
2 87072 1 10720
2 87073 1 10720
2 87074 1 10720
2 87075 1 10720
2 87076 1 10720
2 87077 1 10720
2 87078 1 10720
2 87079 1 10720
2 87080 1 10720
2 87081 1 10720
2 87082 1 10721
2 87083 1 10721
2 87084 1 10730
2 87085 1 10730
2 87086 1 10730
2 87087 1 10734
2 87088 1 10734
2 87089 1 10734
2 87090 1 10735
2 87091 1 10735
2 87092 1 10735
2 87093 1 10736
2 87094 1 10736
2 87095 1 10736
2 87096 1 10736
2 87097 1 10736
2 87098 1 10736
2 87099 1 10736
2 87100 1 10737
2 87101 1 10737
2 87102 1 10739
2 87103 1 10739
2 87104 1 10739
2 87105 1 10739
2 87106 1 10739
2 87107 1 10739
2 87108 1 10739
2 87109 1 10740
2 87110 1 10740
2 87111 1 10754
2 87112 1 10754
2 87113 1 10754
2 87114 1 10754
2 87115 1 10754
2 87116 1 10754
2 87117 1 10754
2 87118 1 10754
2 87119 1 10754
2 87120 1 10754
2 87121 1 10754
2 87122 1 10754
2 87123 1 10754
2 87124 1 10754
2 87125 1 10754
2 87126 1 10754
2 87127 1 10754
2 87128 1 10754
2 87129 1 10754
2 87130 1 10754
2 87131 1 10754
2 87132 1 10755
2 87133 1 10755
2 87134 1 10755
2 87135 1 10755
2 87136 1 10756
2 87137 1 10756
2 87138 1 10756
2 87139 1 10756
2 87140 1 10756
2 87141 1 10756
2 87142 1 10756
2 87143 1 10756
2 87144 1 10756
2 87145 1 10767
2 87146 1 10767
2 87147 1 10767
2 87148 1 10767
2 87149 1 10767
2 87150 1 10767
2 87151 1 10767
2 87152 1 10767
2 87153 1 10769
2 87154 1 10769
2 87155 1 10769
2 87156 1 10769
2 87157 1 10770
2 87158 1 10770
2 87159 1 10770
2 87160 1 10770
2 87161 1 10770
2 87162 1 10770
2 87163 1 10770
2 87164 1 10770
2 87165 1 10770
2 87166 1 10770
2 87167 1 10770
2 87168 1 10770
2 87169 1 10770
2 87170 1 10770
2 87171 1 10770
2 87172 1 10770
2 87173 1 10770
2 87174 1 10770
2 87175 1 10770
2 87176 1 10770
2 87177 1 10770
2 87178 1 10770
2 87179 1 10770
2 87180 1 10770
2 87181 1 10770
2 87182 1 10770
2 87183 1 10770
2 87184 1 10770
2 87185 1 10770
2 87186 1 10770
2 87187 1 10770
2 87188 1 10770
2 87189 1 10770
2 87190 1 10770
2 87191 1 10770
2 87192 1 10770
2 87193 1 10770
2 87194 1 10770
2 87195 1 10770
2 87196 1 10770
2 87197 1 10770
2 87198 1 10770
2 87199 1 10770
2 87200 1 10770
2 87201 1 10771
2 87202 1 10771
2 87203 1 10779
2 87204 1 10779
2 87205 1 10779
2 87206 1 10779
2 87207 1 10779
2 87208 1 10779
2 87209 1 10779
2 87210 1 10779
2 87211 1 10779
2 87212 1 10779
2 87213 1 10779
2 87214 1 10779
2 87215 1 10779
2 87216 1 10779
2 87217 1 10779
2 87218 1 10780
2 87219 1 10780
2 87220 1 10781
2 87221 1 10781
2 87222 1 10782
2 87223 1 10782
2 87224 1 10782
2 87225 1 10782
2 87226 1 10782
2 87227 1 10783
2 87228 1 10783
2 87229 1 10784
2 87230 1 10784
2 87231 1 10784
2 87232 1 10784
2 87233 1 10784
2 87234 1 10785
2 87235 1 10785
2 87236 1 10785
2 87237 1 10785
2 87238 1 10785
2 87239 1 10785
2 87240 1 10785
2 87241 1 10785
2 87242 1 10785
2 87243 1 10785
2 87244 1 10785
2 87245 1 10785
2 87246 1 10785
2 87247 1 10786
2 87248 1 10786
2 87249 1 10786
2 87250 1 10786
2 87251 1 10788
2 87252 1 10788
2 87253 1 10795
2 87254 1 10795
2 87255 1 10796
2 87256 1 10796
2 87257 1 10806
2 87258 1 10806
2 87259 1 10806
2 87260 1 10806
2 87261 1 10806
2 87262 1 10806
2 87263 1 10806
2 87264 1 10806
2 87265 1 10806
2 87266 1 10806
2 87267 1 10807
2 87268 1 10807
2 87269 1 10807
2 87270 1 10807
2 87271 1 10807
2 87272 1 10807
2 87273 1 10810
2 87274 1 10810
2 87275 1 10810
2 87276 1 10810
2 87277 1 10810
2 87278 1 10810
2 87279 1 10810
2 87280 1 10810
2 87281 1 10830
2 87282 1 10830
2 87283 1 10835
2 87284 1 10835
2 87285 1 10836
2 87286 1 10836
2 87287 1 10843
2 87288 1 10843
2 87289 1 10843
2 87290 1 10843
2 87291 1 10843
2 87292 1 10843
2 87293 1 10843
2 87294 1 10843
2 87295 1 10843
2 87296 1 10843
2 87297 1 10843
2 87298 1 10844
2 87299 1 10844
2 87300 1 10844
2 87301 1 10844
2 87302 1 10844
2 87303 1 10844
2 87304 1 10844
2 87305 1 10844
2 87306 1 10845
2 87307 1 10845
2 87308 1 10845
2 87309 1 10852
2 87310 1 10852
2 87311 1 10852
2 87312 1 10852
2 87313 1 10852
2 87314 1 10852
2 87315 1 10852
2 87316 1 10852
2 87317 1 10852
2 87318 1 10852
2 87319 1 10852
2 87320 1 10852
2 87321 1 10853
2 87322 1 10853
2 87323 1 10853
2 87324 1 10855
2 87325 1 10855
2 87326 1 10855
2 87327 1 10855
2 87328 1 10857
2 87329 1 10857
2 87330 1 10857
2 87331 1 10859
2 87332 1 10859
2 87333 1 10859
2 87334 1 10859
2 87335 1 10859
2 87336 1 10859
2 87337 1 10859
2 87338 1 10859
2 87339 1 10859
2 87340 1 10860
2 87341 1 10860
2 87342 1 10860
2 87343 1 10860
2 87344 1 10860
2 87345 1 10860
2 87346 1 10861
2 87347 1 10861
2 87348 1 10861
2 87349 1 10877
2 87350 1 10877
2 87351 1 10898
2 87352 1 10898
2 87353 1 10898
2 87354 1 10899
2 87355 1 10899
2 87356 1 10899
2 87357 1 10899
2 87358 1 10899
2 87359 1 10899
2 87360 1 10900
2 87361 1 10900
2 87362 1 10908
2 87363 1 10908
2 87364 1 10913
2 87365 1 10913
2 87366 1 10913
2 87367 1 10913
2 87368 1 10913
2 87369 1 10913
2 87370 1 10913
2 87371 1 10917
2 87372 1 10917
2 87373 1 10917
2 87374 1 10917
2 87375 1 10917
2 87376 1 10919
2 87377 1 10919
2 87378 1 10920
2 87379 1 10920
2 87380 1 10920
2 87381 1 10920
2 87382 1 10932
2 87383 1 10932
2 87384 1 10932
2 87385 1 10932
2 87386 1 10932
2 87387 1 10932
2 87388 1 10932
2 87389 1 10932
2 87390 1 10932
2 87391 1 10932
2 87392 1 10932
2 87393 1 10932
2 87394 1 10932
2 87395 1 10932
2 87396 1 10932
2 87397 1 10932
2 87398 1 10932
2 87399 1 10932
2 87400 1 10932
2 87401 1 10932
2 87402 1 10932
2 87403 1 10932
2 87404 1 10939
2 87405 1 10939
2 87406 1 10939
2 87407 1 10939
2 87408 1 10941
2 87409 1 10941
2 87410 1 10941
2 87411 1 10947
2 87412 1 10947
2 87413 1 10963
2 87414 1 10963
2 87415 1 10963
2 87416 1 10963
2 87417 1 10966
2 87418 1 10966
2 87419 1 10966
2 87420 1 10966
2 87421 1 10966
2 87422 1 10967
2 87423 1 10967
2 87424 1 10967
2 87425 1 10967
2 87426 1 10967
2 87427 1 10967
2 87428 1 10967
2 87429 1 10967
2 87430 1 10967
2 87431 1 10967
2 87432 1 10967
2 87433 1 10967
2 87434 1 10967
2 87435 1 10967
2 87436 1 10967
2 87437 1 10967
2 87438 1 10967
2 87439 1 10967
2 87440 1 10982
2 87441 1 10982
2 87442 1 10983
2 87443 1 10983
2 87444 1 10983
2 87445 1 10983
2 87446 1 10983
2 87447 1 10983
2 87448 1 10993
2 87449 1 10993
2 87450 1 10993
2 87451 1 10994
2 87452 1 10994
2 87453 1 10997
2 87454 1 10997
2 87455 1 10997
2 87456 1 10997
2 87457 1 11012
2 87458 1 11012
2 87459 1 11012
2 87460 1 11012
2 87461 1 11012
2 87462 1 11012
2 87463 1 11012
2 87464 1 11012
2 87465 1 11015
2 87466 1 11015
2 87467 1 11015
2 87468 1 11015
2 87469 1 11016
2 87470 1 11016
2 87471 1 11016
2 87472 1 11025
2 87473 1 11025
2 87474 1 11025
2 87475 1 11025
2 87476 1 11025
2 87477 1 11033
2 87478 1 11033
2 87479 1 11034
2 87480 1 11034
2 87481 1 11034
2 87482 1 11034
2 87483 1 11034
2 87484 1 11042
2 87485 1 11042
2 87486 1 11042
2 87487 1 11042
2 87488 1 11046
2 87489 1 11046
2 87490 1 11055
2 87491 1 11055
2 87492 1 11063
2 87493 1 11063
2 87494 1 11063
2 87495 1 11063
2 87496 1 11066
2 87497 1 11066
2 87498 1 11067
2 87499 1 11067
2 87500 1 11067
2 87501 1 11067
2 87502 1 11067
2 87503 1 11067
2 87504 1 11067
2 87505 1 11067
2 87506 1 11067
2 87507 1 11067
2 87508 1 11067
2 87509 1 11067
2 87510 1 11068
2 87511 1 11068
2 87512 1 11068
2 87513 1 11068
2 87514 1 11068
2 87515 1 11068
2 87516 1 11068
2 87517 1 11068
2 87518 1 11068
2 87519 1 11070
2 87520 1 11070
2 87521 1 11072
2 87522 1 11072
2 87523 1 11073
2 87524 1 11073
2 87525 1 11073
2 87526 1 11073
2 87527 1 11073
2 87528 1 11073
2 87529 1 11073
2 87530 1 11073
2 87531 1 11073
2 87532 1 11077
2 87533 1 11077
2 87534 1 11078
2 87535 1 11078
2 87536 1 11083
2 87537 1 11083
2 87538 1 11083
2 87539 1 11100
2 87540 1 11100
2 87541 1 11100
2 87542 1 11100
2 87543 1 11103
2 87544 1 11103
2 87545 1 11114
2 87546 1 11114
2 87547 1 11123
2 87548 1 11123
2 87549 1 11123
2 87550 1 11123
2 87551 1 11123
2 87552 1 11124
2 87553 1 11124
2 87554 1 11124
2 87555 1 11135
2 87556 1 11135
2 87557 1 11135
2 87558 1 11135
2 87559 1 11136
2 87560 1 11136
2 87561 1 11137
2 87562 1 11137
2 87563 1 11141
2 87564 1 11141
2 87565 1 11141
2 87566 1 11142
2 87567 1 11142
2 87568 1 11156
2 87569 1 11156
2 87570 1 11157
2 87571 1 11157
2 87572 1 11165
2 87573 1 11165
2 87574 1 11165
2 87575 1 11165
2 87576 1 11165
2 87577 1 11165
2 87578 1 11165
2 87579 1 11165
2 87580 1 11166
2 87581 1 11166
2 87582 1 11174
2 87583 1 11174
2 87584 1 11176
2 87585 1 11176
2 87586 1 11176
2 87587 1 11176
2 87588 1 11176
2 87589 1 11177
2 87590 1 11177
2 87591 1 11177
2 87592 1 11177
2 87593 1 11177
2 87594 1 11177
2 87595 1 11181
2 87596 1 11181
2 87597 1 11181
2 87598 1 11181
2 87599 1 11182
2 87600 1 11182
2 87601 1 11182
2 87602 1 11183
2 87603 1 11183
2 87604 1 11183
2 87605 1 11183
2 87606 1 11183
2 87607 1 11192
2 87608 1 11192
2 87609 1 11192
2 87610 1 11192
2 87611 1 11192
2 87612 1 11192
2 87613 1 11192
2 87614 1 11193
2 87615 1 11193
2 87616 1 11193
2 87617 1 11194
2 87618 1 11194
2 87619 1 11205
2 87620 1 11205
2 87621 1 11205
2 87622 1 11205
2 87623 1 11205
2 87624 1 11205
2 87625 1 11205
2 87626 1 11219
2 87627 1 11219
2 87628 1 11219
2 87629 1 11219
2 87630 1 11219
2 87631 1 11219
2 87632 1 11219
2 87633 1 11220
2 87634 1 11220
2 87635 1 11221
2 87636 1 11221
2 87637 1 11221
2 87638 1 11221
2 87639 1 11221
2 87640 1 11221
2 87641 1 11221
2 87642 1 11221
2 87643 1 11221
2 87644 1 11221
2 87645 1 11222
2 87646 1 11222
2 87647 1 11241
2 87648 1 11241
2 87649 1 11241
2 87650 1 11241
2 87651 1 11242
2 87652 1 11242
2 87653 1 11252
2 87654 1 11252
2 87655 1 11253
2 87656 1 11253
2 87657 1 11253
2 87658 1 11253
2 87659 1 11253
2 87660 1 11253
2 87661 1 11265
2 87662 1 11265
2 87663 1 11265
2 87664 1 11265
2 87665 1 11265
2 87666 1 11265
2 87667 1 11265
2 87668 1 11265
2 87669 1 11265
2 87670 1 11265
2 87671 1 11271
2 87672 1 11271
2 87673 1 11273
2 87674 1 11273
2 87675 1 11273
2 87676 1 11274
2 87677 1 11274
2 87678 1 11279
2 87679 1 11279
2 87680 1 11282
2 87681 1 11282
2 87682 1 11282
2 87683 1 11282
2 87684 1 11283
2 87685 1 11283
2 87686 1 11288
2 87687 1 11288
2 87688 1 11309
2 87689 1 11309
2 87690 1 11309
2 87691 1 11329
2 87692 1 11329
2 87693 1 11343
2 87694 1 11343
2 87695 1 11351
2 87696 1 11351
2 87697 1 11351
2 87698 1 11359
2 87699 1 11359
2 87700 1 11360
2 87701 1 11360
2 87702 1 11360
2 87703 1 11360
2 87704 1 11368
2 87705 1 11368
2 87706 1 11378
2 87707 1 11378
2 87708 1 11378
2 87709 1 11379
2 87710 1 11379
2 87711 1 11379
2 87712 1 11379
2 87713 1 11380
2 87714 1 11380
2 87715 1 11380
2 87716 1 11380
2 87717 1 11380
2 87718 1 11381
2 87719 1 11381
2 87720 1 11381
2 87721 1 11381
2 87722 1 11382
2 87723 1 11382
2 87724 1 11383
2 87725 1 11383
2 87726 1 11383
2 87727 1 11383
2 87728 1 11388
2 87729 1 11388
2 87730 1 11388
2 87731 1 11388
2 87732 1 11388
2 87733 1 11388
2 87734 1 11388
2 87735 1 11388
2 87736 1 11405
2 87737 1 11405
2 87738 1 11405
2 87739 1 11417
2 87740 1 11417
2 87741 1 11427
2 87742 1 11427
2 87743 1 11428
2 87744 1 11428
2 87745 1 11434
2 87746 1 11434
2 87747 1 11451
2 87748 1 11451
2 87749 1 11451
2 87750 1 11452
2 87751 1 11452
2 87752 1 11453
2 87753 1 11453
2 87754 1 11461
2 87755 1 11461
2 87756 1 11461
2 87757 1 11461
2 87758 1 11461
2 87759 1 11461
2 87760 1 11461
2 87761 1 11461
2 87762 1 11461
2 87763 1 11461
2 87764 1 11462
2 87765 1 11462
2 87766 1 11462
2 87767 1 11462
2 87768 1 11463
2 87769 1 11463
2 87770 1 11463
2 87771 1 11468
2 87772 1 11468
2 87773 1 11472
2 87774 1 11472
2 87775 1 11472
2 87776 1 11482
2 87777 1 11482
2 87778 1 11483
2 87779 1 11483
2 87780 1 11492
2 87781 1 11492
2 87782 1 11493
2 87783 1 11493
2 87784 1 11493
2 87785 1 11493
2 87786 1 11496
2 87787 1 11496
2 87788 1 11497
2 87789 1 11497
2 87790 1 11497
2 87791 1 11497
2 87792 1 11497
2 87793 1 11497
2 87794 1 11506
2 87795 1 11506
2 87796 1 11507
2 87797 1 11507
2 87798 1 11515
2 87799 1 11515
2 87800 1 11515
2 87801 1 11515
2 87802 1 11515
2 87803 1 11515
2 87804 1 11517
2 87805 1 11517
2 87806 1 11517
2 87807 1 11518
2 87808 1 11518
2 87809 1 11521
2 87810 1 11521
2 87811 1 11521
2 87812 1 11521
2 87813 1 11522
2 87814 1 11522
2 87815 1 11530
2 87816 1 11530
2 87817 1 11554
2 87818 1 11554
2 87819 1 11554
2 87820 1 11556
2 87821 1 11556
2 87822 1 11556
2 87823 1 11556
2 87824 1 11556
2 87825 1 11556
2 87826 1 11556
2 87827 1 11557
2 87828 1 11557
2 87829 1 11557
2 87830 1 11557
2 87831 1 11557
2 87832 1 11557
2 87833 1 11558
2 87834 1 11558
2 87835 1 11567
2 87836 1 11567
2 87837 1 11567
2 87838 1 11571
2 87839 1 11571
2 87840 1 11582
2 87841 1 11582
2 87842 1 11582
2 87843 1 11582
2 87844 1 11582
2 87845 1 11582
2 87846 1 11582
2 87847 1 11583
2 87848 1 11583
2 87849 1 11583
2 87850 1 11584
2 87851 1 11584
2 87852 1 11585
2 87853 1 11585
2 87854 1 11585
2 87855 1 11585
2 87856 1 11585
2 87857 1 11585
2 87858 1 11585
2 87859 1 11585
2 87860 1 11585
2 87861 1 11585
2 87862 1 11585
2 87863 1 11585
2 87864 1 11585
2 87865 1 11585
2 87866 1 11585
2 87867 1 11585
2 87868 1 11585
2 87869 1 11585
2 87870 1 11585
2 87871 1 11585
2 87872 1 11585
2 87873 1 11586
2 87874 1 11586
2 87875 1 11588
2 87876 1 11588
2 87877 1 11595
2 87878 1 11595
2 87879 1 11595
2 87880 1 11595
2 87881 1 11595
2 87882 1 11595
2 87883 1 11596
2 87884 1 11596
2 87885 1 11599
2 87886 1 11599
2 87887 1 11600
2 87888 1 11600
2 87889 1 11605
2 87890 1 11605
2 87891 1 11605
2 87892 1 11605
2 87893 1 11605
2 87894 1 11605
2 87895 1 11612
2 87896 1 11612
2 87897 1 11612
2 87898 1 11620
2 87899 1 11620
2 87900 1 11640
2 87901 1 11640
2 87902 1 11640
2 87903 1 11644
2 87904 1 11644
2 87905 1 11644
2 87906 1 11653
2 87907 1 11653
2 87908 1 11653
2 87909 1 11653
2 87910 1 11667
2 87911 1 11667
2 87912 1 11667
2 87913 1 11667
2 87914 1 11667
2 87915 1 11667
2 87916 1 11667
2 87917 1 11667
2 87918 1 11668
2 87919 1 11668
2 87920 1 11668
2 87921 1 11673
2 87922 1 11673
2 87923 1 11674
2 87924 1 11674
2 87925 1 11674
2 87926 1 11674
2 87927 1 11674
2 87928 1 11675
2 87929 1 11675
2 87930 1 11675
2 87931 1 11679
2 87932 1 11679
2 87933 1 11679
2 87934 1 11679
2 87935 1 11687
2 87936 1 11687
2 87937 1 11696
2 87938 1 11696
2 87939 1 11699
2 87940 1 11699
2 87941 1 11699
2 87942 1 11699
2 87943 1 11699
2 87944 1 11699
2 87945 1 11700
2 87946 1 11700
2 87947 1 11710
2 87948 1 11710
2 87949 1 11713
2 87950 1 11713
2 87951 1 11713
2 87952 1 11713
2 87953 1 11713
2 87954 1 11713
2 87955 1 11713
2 87956 1 11732
2 87957 1 11732
2 87958 1 11733
2 87959 1 11733
2 87960 1 11733
2 87961 1 11745
2 87962 1 11745
2 87963 1 11760
2 87964 1 11760
2 87965 1 11760
2 87966 1 11761
2 87967 1 11761
2 87968 1 11774
2 87969 1 11774
2 87970 1 11774
2 87971 1 11774
2 87972 1 11774
2 87973 1 11775
2 87974 1 11775
2 87975 1 11801
2 87976 1 11801
2 87977 1 11802
2 87978 1 11802
2 87979 1 11820
2 87980 1 11820
2 87981 1 11827
2 87982 1 11827
2 87983 1 11829
2 87984 1 11829
2 87985 1 11830
2 87986 1 11830
2 87987 1 11830
2 87988 1 11862
2 87989 1 11862
2 87990 1 11890
2 87991 1 11890
2 87992 1 11890
2 87993 1 11890
2 87994 1 11890
2 87995 1 11890
2 87996 1 11891
2 87997 1 11891
2 87998 1 11891
2 87999 1 11891
2 88000 1 11891
2 88001 1 11891
2 88002 1 11892
2 88003 1 11892
2 88004 1 11892
2 88005 1 11893
2 88006 1 11893
2 88007 1 11893
2 88008 1 11893
2 88009 1 11901
2 88010 1 11901
2 88011 1 11901
2 88012 1 11901
2 88013 1 11901
2 88014 1 11901
2 88015 1 11901
2 88016 1 11901
2 88017 1 11902
2 88018 1 11902
2 88019 1 11902
2 88020 1 11902
2 88021 1 11902
2 88022 1 11902
2 88023 1 11902
2 88024 1 11902
2 88025 1 11903
2 88026 1 11903
2 88027 1 11920
2 88028 1 11920
2 88029 1 11920
2 88030 1 11920
2 88031 1 11921
2 88032 1 11921
2 88033 1 11921
2 88034 1 11921
2 88035 1 11926
2 88036 1 11926
2 88037 1 11926
2 88038 1 11926
2 88039 1 11926
2 88040 1 11926
2 88041 1 11928
2 88042 1 11928
2 88043 1 11930
2 88044 1 11930
2 88045 1 11930
2 88046 1 11930
2 88047 1 11931
2 88048 1 11931
2 88049 1 11932
2 88050 1 11932
2 88051 1 11932
2 88052 1 11933
2 88053 1 11933
2 88054 1 11940
2 88055 1 11940
2 88056 1 11940
2 88057 1 11940
2 88058 1 11941
2 88059 1 11941
2 88060 1 11941
2 88061 1 11953
2 88062 1 11953
2 88063 1 11967
2 88064 1 11967
2 88065 1 11978
2 88066 1 11978
2 88067 1 11978
2 88068 1 11978
2 88069 1 11978
2 88070 1 11978
2 88071 1 11978
2 88072 1 11978
2 88073 1 11978
2 88074 1 11978
2 88075 1 11978
2 88076 1 11978
2 88077 1 11986
2 88078 1 11986
2 88079 1 11990
2 88080 1 11990
2 88081 1 11990
2 88082 1 11990
2 88083 1 11990
2 88084 1 11990
2 88085 1 11990
2 88086 1 11990
2 88087 1 11990
2 88088 1 11990
2 88089 1 11990
2 88090 1 11990
2 88091 1 11990
2 88092 1 11990
2 88093 1 11991
2 88094 1 11991
2 88095 1 11991
2 88096 1 11992
2 88097 1 11992
2 88098 1 11992
2 88099 1 11992
2 88100 1 11992
2 88101 1 11992
2 88102 1 11992
2 88103 1 11992
2 88104 1 11992
2 88105 1 11992
2 88106 1 11992
2 88107 1 11992
2 88108 1 11992
2 88109 1 11992
2 88110 1 11992
2 88111 1 11992
2 88112 1 11993
2 88113 1 11993
2 88114 1 12000
2 88115 1 12000
2 88116 1 12000
2 88117 1 12000
2 88118 1 12000
2 88119 1 12000
2 88120 1 12000
2 88121 1 12000
2 88122 1 12000
2 88123 1 12000
2 88124 1 12000
2 88125 1 12000
2 88126 1 12017
2 88127 1 12017
2 88128 1 12017
2 88129 1 12017
2 88130 1 12017
2 88131 1 12017
2 88132 1 12025
2 88133 1 12025
2 88134 1 12025
2 88135 1 12025
2 88136 1 12025
2 88137 1 12025
2 88138 1 12025
2 88139 1 12025
2 88140 1 12026
2 88141 1 12026
2 88142 1 12039
2 88143 1 12039
2 88144 1 12043
2 88145 1 12043
2 88146 1 12074
2 88147 1 12074
2 88148 1 12074
2 88149 1 12075
2 88150 1 12075
2 88151 1 12075
2 88152 1 12075
2 88153 1 12075
2 88154 1 12075
2 88155 1 12084
2 88156 1 12084
2 88157 1 12097
2 88158 1 12097
2 88159 1 12097
2 88160 1 12097
2 88161 1 12114
2 88162 1 12114
2 88163 1 12114
2 88164 1 12114
2 88165 1 12115
2 88166 1 12115
2 88167 1 12115
2 88168 1 12115
2 88169 1 12115
2 88170 1 12125
2 88171 1 12125
2 88172 1 12126
2 88173 1 12126
2 88174 1 12126
2 88175 1 12128
2 88176 1 12128
2 88177 1 12128
2 88178 1 12133
2 88179 1 12133
2 88180 1 12133
2 88181 1 12146
2 88182 1 12146
2 88183 1 12161
2 88184 1 12161
2 88185 1 12161
2 88186 1 12161
2 88187 1 12161
2 88188 1 12161
2 88189 1 12161
2 88190 1 12161
2 88191 1 12163
2 88192 1 12163
2 88193 1 12163
2 88194 1 12163
2 88195 1 12163
2 88196 1 12163
2 88197 1 12163
2 88198 1 12163
2 88199 1 12163
2 88200 1 12163
2 88201 1 12165
2 88202 1 12165
2 88203 1 12167
2 88204 1 12167
2 88205 1 12169
2 88206 1 12169
2 88207 1 12187
2 88208 1 12187
2 88209 1 12216
2 88210 1 12216
2 88211 1 12216
2 88212 1 12216
2 88213 1 12216
2 88214 1 12228
2 88215 1 12228
2 88216 1 12245
2 88217 1 12245
2 88218 1 12245
2 88219 1 12255
2 88220 1 12255
2 88221 1 12262
2 88222 1 12262
2 88223 1 12262
2 88224 1 12262
2 88225 1 12273
2 88226 1 12273
2 88227 1 12273
2 88228 1 12273
2 88229 1 12273
2 88230 1 12274
2 88231 1 12274
2 88232 1 12274
2 88233 1 12274
2 88234 1 12274
2 88235 1 12274
2 88236 1 12274
2 88237 1 12274
2 88238 1 12274
2 88239 1 12275
2 88240 1 12275
2 88241 1 12276
2 88242 1 12276
2 88243 1 12284
2 88244 1 12284
2 88245 1 12285
2 88246 1 12285
2 88247 1 12285
2 88248 1 12285
2 88249 1 12285
2 88250 1 12286
2 88251 1 12286
2 88252 1 12287
2 88253 1 12287
2 88254 1 12287
2 88255 1 12297
2 88256 1 12297
2 88257 1 12305
2 88258 1 12305
2 88259 1 12313
2 88260 1 12313
2 88261 1 12313
2 88262 1 12313
2 88263 1 12313
2 88264 1 12313
2 88265 1 12348
2 88266 1 12348
2 88267 1 12349
2 88268 1 12349
2 88269 1 12349
2 88270 1 12350
2 88271 1 12350
2 88272 1 12350
2 88273 1 12350
2 88274 1 12364
2 88275 1 12364
2 88276 1 12370
2 88277 1 12370
2 88278 1 12380
2 88279 1 12380
2 88280 1 12380
2 88281 1 12381
2 88282 1 12381
2 88283 1 12409
2 88284 1 12409
2 88285 1 12409
2 88286 1 12409
2 88287 1 12428
2 88288 1 12428
2 88289 1 12428
2 88290 1 12429
2 88291 1 12429
2 88292 1 12429
2 88293 1 12436
2 88294 1 12436
2 88295 1 12437
2 88296 1 12437
2 88297 1 12438
2 88298 1 12438
2 88299 1 12438
2 88300 1 12438
2 88301 1 12460
2 88302 1 12460
2 88303 1 12469
2 88304 1 12469
2 88305 1 12470
2 88306 1 12470
2 88307 1 12471
2 88308 1 12471
2 88309 1 12481
2 88310 1 12481
2 88311 1 12481
2 88312 1 12490
2 88313 1 12490
2 88314 1 12497
2 88315 1 12497
2 88316 1 12519
2 88317 1 12519
2 88318 1 12519
2 88319 1 12519
2 88320 1 12519
2 88321 1 12545
2 88322 1 12545
2 88323 1 12545
2 88324 1 12545
2 88325 1 12553
2 88326 1 12553
2 88327 1 12564
2 88328 1 12564
2 88329 1 12564
2 88330 1 12564
2 88331 1 12566
2 88332 1 12566
2 88333 1 12566
2 88334 1 12566
2 88335 1 12567
2 88336 1 12567
2 88337 1 12567
2 88338 1 12584
2 88339 1 12584
2 88340 1 12584
2 88341 1 12584
2 88342 1 12584
2 88343 1 12584
2 88344 1 12584
2 88345 1 12591
2 88346 1 12591
2 88347 1 12600
2 88348 1 12600
2 88349 1 12619
2 88350 1 12619
2 88351 1 12621
2 88352 1 12621
2 88353 1 12621
2 88354 1 12621
2 88355 1 12625
2 88356 1 12625
2 88357 1 12625
2 88358 1 12625
2 88359 1 12625
2 88360 1 12625
2 88361 1 12625
2 88362 1 12625
2 88363 1 12625
2 88364 1 12626
2 88365 1 12626
2 88366 1 12626
2 88367 1 12626
2 88368 1 12626
2 88369 1 12629
2 88370 1 12629
2 88371 1 12630
2 88372 1 12630
2 88373 1 12649
2 88374 1 12649
2 88375 1 12652
2 88376 1 12652
2 88377 1 12655
2 88378 1 12655
2 88379 1 12656
2 88380 1 12656
2 88381 1 12656
2 88382 1 12657
2 88383 1 12657
2 88384 1 12658
2 88385 1 12658
2 88386 1 12662
2 88387 1 12662
2 88388 1 12670
2 88389 1 12670
2 88390 1 12670
2 88391 1 12670
2 88392 1 12670
2 88393 1 12670
2 88394 1 12670
2 88395 1 12670
2 88396 1 12670
2 88397 1 12673
2 88398 1 12673
2 88399 1 12687
2 88400 1 12687
2 88401 1 12687
2 88402 1 12688
2 88403 1 12688
2 88404 1 12688
2 88405 1 12689
2 88406 1 12689
2 88407 1 12690
2 88408 1 12690
2 88409 1 12694
2 88410 1 12694
2 88411 1 12695
2 88412 1 12695
2 88413 1 12695
2 88414 1 12695
2 88415 1 12695
2 88416 1 12695
2 88417 1 12695
2 88418 1 12695
2 88419 1 12695
2 88420 1 12696
2 88421 1 12696
2 88422 1 12696
2 88423 1 12696
2 88424 1 12696
2 88425 1 12696
2 88426 1 12696
2 88427 1 12696
2 88428 1 12705
2 88429 1 12705
2 88430 1 12705
2 88431 1 12706
2 88432 1 12706
2 88433 1 12709
2 88434 1 12709
2 88435 1 12730
2 88436 1 12730
2 88437 1 12731
2 88438 1 12731
2 88439 1 12731
2 88440 1 12731
2 88441 1 12732
2 88442 1 12732
2 88443 1 12745
2 88444 1 12745
2 88445 1 12745
2 88446 1 12747
2 88447 1 12747
2 88448 1 12747
2 88449 1 12747
2 88450 1 12747
2 88451 1 12747
2 88452 1 12748
2 88453 1 12748
2 88454 1 12748
2 88455 1 12748
2 88456 1 12749
2 88457 1 12749
2 88458 1 12749
2 88459 1 12749
2 88460 1 12749
2 88461 1 12749
2 88462 1 12749
2 88463 1 12749
2 88464 1 12749
2 88465 1 12749
2 88466 1 12749
2 88467 1 12749
2 88468 1 12749
2 88469 1 12749
2 88470 1 12749
2 88471 1 12749
2 88472 1 12749
2 88473 1 12749
2 88474 1 12749
2 88475 1 12749
2 88476 1 12749
2 88477 1 12749
2 88478 1 12749
2 88479 1 12749
2 88480 1 12749
2 88481 1 12749
2 88482 1 12749
2 88483 1 12750
2 88484 1 12750
2 88485 1 12752
2 88486 1 12752
2 88487 1 12752
2 88488 1 12753
2 88489 1 12753
2 88490 1 12753
2 88491 1 12755
2 88492 1 12755
2 88493 1 12755
2 88494 1 12755
2 88495 1 12755
2 88496 1 12759
2 88497 1 12759
2 88498 1 12761
2 88499 1 12761
2 88500 1 12767
2 88501 1 12767
2 88502 1 12773
2 88503 1 12773
2 88504 1 12773
2 88505 1 12774
2 88506 1 12774
2 88507 1 12774
2 88508 1 12774
2 88509 1 12774
2 88510 1 12774
2 88511 1 12774
2 88512 1 12775
2 88513 1 12775
2 88514 1 12777
2 88515 1 12777
2 88516 1 12777
2 88517 1 12778
2 88518 1 12778
2 88519 1 12778
2 88520 1 12778
2 88521 1 12778
2 88522 1 12779
2 88523 1 12779
2 88524 1 12781
2 88525 1 12781
2 88526 1 12795
2 88527 1 12795
2 88528 1 12795
2 88529 1 12796
2 88530 1 12796
2 88531 1 12796
2 88532 1 12796
2 88533 1 12802
2 88534 1 12802
2 88535 1 12805
2 88536 1 12805
2 88537 1 12805
2 88538 1 12809
2 88539 1 12809
2 88540 1 12809
2 88541 1 12809
2 88542 1 12809
2 88543 1 12809
2 88544 1 12809
2 88545 1 12816
2 88546 1 12816
2 88547 1 12816
2 88548 1 12816
2 88549 1 12823
2 88550 1 12823
2 88551 1 12824
2 88552 1 12824
2 88553 1 12831
2 88554 1 12831
2 88555 1 12832
2 88556 1 12832
2 88557 1 12832
2 88558 1 12842
2 88559 1 12842
2 88560 1 12843
2 88561 1 12843
2 88562 1 12843
2 88563 1 12844
2 88564 1 12844
2 88565 1 12848
2 88566 1 12848
2 88567 1 12848
2 88568 1 12848
2 88569 1 12849
2 88570 1 12849
2 88571 1 12849
2 88572 1 12849
2 88573 1 12849
2 88574 1 12851
2 88575 1 12851
2 88576 1 12859
2 88577 1 12859
2 88578 1 12860
2 88579 1 12860
2 88580 1 12860
2 88581 1 12860
2 88582 1 12860
2 88583 1 12860
2 88584 1 12860
2 88585 1 12867
2 88586 1 12867
2 88587 1 12867
2 88588 1 12868
2 88589 1 12868
2 88590 1 12869
2 88591 1 12869
2 88592 1 12869
2 88593 1 12870
2 88594 1 12870
2 88595 1 12883
2 88596 1 12883
2 88597 1 12883
2 88598 1 12883
2 88599 1 12894
2 88600 1 12894
2 88601 1 12895
2 88602 1 12895
2 88603 1 12896
2 88604 1 12896
2 88605 1 12896
2 88606 1 12896
2 88607 1 12896
2 88608 1 12896
2 88609 1 12896
2 88610 1 12896
2 88611 1 12896
2 88612 1 12896
2 88613 1 12896
2 88614 1 12896
2 88615 1 12896
2 88616 1 12896
2 88617 1 12896
2 88618 1 12896
2 88619 1 12896
2 88620 1 12896
2 88621 1 12920
2 88622 1 12920
2 88623 1 12937
2 88624 1 12937
2 88625 1 12937
2 88626 1 12937
2 88627 1 12937
2 88628 1 12937
2 88629 1 12937
2 88630 1 12938
2 88631 1 12938
2 88632 1 12938
2 88633 1 12938
2 88634 1 12939
2 88635 1 12939
2 88636 1 12939
2 88637 1 12941
2 88638 1 12941
2 88639 1 12943
2 88640 1 12943
2 88641 1 12943
2 88642 1 12943
2 88643 1 12951
2 88644 1 12951
2 88645 1 12951
2 88646 1 12951
2 88647 1 12951
2 88648 1 12951
2 88649 1 12951
2 88650 1 12964
2 88651 1 12964
2 88652 1 12964
2 88653 1 12964
2 88654 1 12964
2 88655 1 12964
2 88656 1 12964
2 88657 1 12966
2 88658 1 12966
2 88659 1 12976
2 88660 1 12976
2 88661 1 12996
2 88662 1 12996
2 88663 1 13000
2 88664 1 13000
2 88665 1 13008
2 88666 1 13008
2 88667 1 13009
2 88668 1 13009
2 88669 1 13018
2 88670 1 13018
2 88671 1 13018
2 88672 1 13021
2 88673 1 13021
2 88674 1 13022
2 88675 1 13022
2 88676 1 13028
2 88677 1 13028
2 88678 1 13039
2 88679 1 13039
2 88680 1 13054
2 88681 1 13054
2 88682 1 13061
2 88683 1 13061
2 88684 1 13061
2 88685 1 13062
2 88686 1 13062
2 88687 1 13062
2 88688 1 13062
2 88689 1 13069
2 88690 1 13069
2 88691 1 13069
2 88692 1 13069
2 88693 1 13070
2 88694 1 13070
2 88695 1 13073
2 88696 1 13073
2 88697 1 13074
2 88698 1 13074
2 88699 1 13074
2 88700 1 13076
2 88701 1 13076
2 88702 1 13081
2 88703 1 13081
2 88704 1 13081
2 88705 1 13093
2 88706 1 13093
2 88707 1 13093
2 88708 1 13094
2 88709 1 13094
2 88710 1 13095
2 88711 1 13095
2 88712 1 13095
2 88713 1 13095
2 88714 1 13096
2 88715 1 13096
2 88716 1 13096
2 88717 1 13096
2 88718 1 13096
2 88719 1 13096
2 88720 1 13113
2 88721 1 13113
2 88722 1 13113
2 88723 1 13113
2 88724 1 13124
2 88725 1 13124
2 88726 1 13132
2 88727 1 13132
2 88728 1 13133
2 88729 1 13133
2 88730 1 13133
2 88731 1 13134
2 88732 1 13134
2 88733 1 13134
2 88734 1 13140
2 88735 1 13140
2 88736 1 13140
2 88737 1 13140
2 88738 1 13140
2 88739 1 13140
2 88740 1 13141
2 88741 1 13141
2 88742 1 13141
2 88743 1 13148
2 88744 1 13148
2 88745 1 13148
2 88746 1 13148
2 88747 1 13148
2 88748 1 13150
2 88749 1 13150
2 88750 1 13151
2 88751 1 13151
2 88752 1 13151
2 88753 1 13151
2 88754 1 13151
2 88755 1 13151
2 88756 1 13151
2 88757 1 13152
2 88758 1 13152
2 88759 1 13152
2 88760 1 13152
2 88761 1 13162
2 88762 1 13162
2 88763 1 13162
2 88764 1 13163
2 88765 1 13163
2 88766 1 13163
2 88767 1 13163
2 88768 1 13163
2 88769 1 13163
2 88770 1 13163
2 88771 1 13163
2 88772 1 13163
2 88773 1 13191
2 88774 1 13191
2 88775 1 13191
2 88776 1 13198
2 88777 1 13198
2 88778 1 13200
2 88779 1 13200
2 88780 1 13200
2 88781 1 13201
2 88782 1 13201
2 88783 1 13205
2 88784 1 13205
2 88785 1 13211
2 88786 1 13211
2 88787 1 13214
2 88788 1 13214
2 88789 1 13215
2 88790 1 13215
2 88791 1 13217
2 88792 1 13217
2 88793 1 13234
2 88794 1 13234
2 88795 1 13238
2 88796 1 13238
2 88797 1 13241
2 88798 1 13241
2 88799 1 13244
2 88800 1 13244
2 88801 1 13272
2 88802 1 13272
2 88803 1 13272
2 88804 1 13272
2 88805 1 13274
2 88806 1 13274
2 88807 1 13274
2 88808 1 13277
2 88809 1 13277
2 88810 1 13277
2 88811 1 13277
2 88812 1 13277
2 88813 1 13277
2 88814 1 13277
2 88815 1 13278
2 88816 1 13278
2 88817 1 13278
2 88818 1 13278
2 88819 1 13278
2 88820 1 13281
2 88821 1 13281
2 88822 1 13282
2 88823 1 13282
2 88824 1 13282
2 88825 1 13282
2 88826 1 13283
2 88827 1 13283
2 88828 1 13283
2 88829 1 13284
2 88830 1 13284
2 88831 1 13284
2 88832 1 13284
2 88833 1 13284
2 88834 1 13285
2 88835 1 13285
2 88836 1 13291
2 88837 1 13291
2 88838 1 13293
2 88839 1 13293
2 88840 1 13294
2 88841 1 13294
2 88842 1 13295
2 88843 1 13295
2 88844 1 13296
2 88845 1 13296
2 88846 1 13297
2 88847 1 13297
2 88848 1 13297
2 88849 1 13297
2 88850 1 13299
2 88851 1 13299
2 88852 1 13302
2 88853 1 13302
2 88854 1 13313
2 88855 1 13313
2 88856 1 13313
2 88857 1 13313
2 88858 1 13313
2 88859 1 13313
2 88860 1 13313
2 88861 1 13313
2 88862 1 13313
2 88863 1 13314
2 88864 1 13314
2 88865 1 13314
2 88866 1 13316
2 88867 1 13316
2 88868 1 13316
2 88869 1 13316
2 88870 1 13317
2 88871 1 13317
2 88872 1 13331
2 88873 1 13331
2 88874 1 13333
2 88875 1 13333
2 88876 1 13333
2 88877 1 13334
2 88878 1 13334
2 88879 1 13334
2 88880 1 13334
2 88881 1 13334
2 88882 1 13334
2 88883 1 13334
2 88884 1 13335
2 88885 1 13335
2 88886 1 13336
2 88887 1 13336
2 88888 1 13336
2 88889 1 13336
2 88890 1 13336
2 88891 1 13352
2 88892 1 13352
2 88893 1 13352
2 88894 1 13352
2 88895 1 13383
2 88896 1 13383
2 88897 1 13383
2 88898 1 13389
2 88899 1 13389
2 88900 1 13411
2 88901 1 13411
2 88902 1 13411
2 88903 1 13411
2 88904 1 13412
2 88905 1 13412
2 88906 1 13412
2 88907 1 13412
2 88908 1 13412
2 88909 1 13417
2 88910 1 13417
2 88911 1 13426
2 88912 1 13426
2 88913 1 13426
2 88914 1 13426
2 88915 1 13427
2 88916 1 13427
2 88917 1 13427
2 88918 1 13427
2 88919 1 13427
2 88920 1 13432
2 88921 1 13432
2 88922 1 13433
2 88923 1 13433
2 88924 1 13438
2 88925 1 13438
2 88926 1 13438
2 88927 1 13438
2 88928 1 13438
2 88929 1 13438
2 88930 1 13439
2 88931 1 13439
2 88932 1 13439
2 88933 1 13439
2 88934 1 13439
2 88935 1 13439
2 88936 1 13439
2 88937 1 13439
2 88938 1 13439
2 88939 1 13447
2 88940 1 13447
2 88941 1 13448
2 88942 1 13448
2 88943 1 13448
2 88944 1 13449
2 88945 1 13449
2 88946 1 13449
2 88947 1 13449
2 88948 1 13449
2 88949 1 13449
2 88950 1 13449
2 88951 1 13449
2 88952 1 13449
2 88953 1 13449
2 88954 1 13449
2 88955 1 13449
2 88956 1 13449
2 88957 1 13449
2 88958 1 13449
2 88959 1 13449
2 88960 1 13449
2 88961 1 13452
2 88962 1 13452
2 88963 1 13452
2 88964 1 13453
2 88965 1 13453
2 88966 1 13461
2 88967 1 13461
2 88968 1 13463
2 88969 1 13463
2 88970 1 13480
2 88971 1 13480
2 88972 1 13480
2 88973 1 13480
2 88974 1 13481
2 88975 1 13481
2 88976 1 13486
2 88977 1 13486
2 88978 1 13486
2 88979 1 13486
2 88980 1 13486
2 88981 1 13486
2 88982 1 13486
2 88983 1 13486
2 88984 1 13486
2 88985 1 13500
2 88986 1 13500
2 88987 1 13500
2 88988 1 13507
2 88989 1 13507
2 88990 1 13507
2 88991 1 13507
2 88992 1 13507
2 88993 1 13507
2 88994 1 13507
2 88995 1 13507
2 88996 1 13507
2 88997 1 13507
2 88998 1 13507
2 88999 1 13507
2 89000 1 13508
2 89001 1 13508
2 89002 1 13509
2 89003 1 13509
2 89004 1 13510
2 89005 1 13510
2 89006 1 13510
2 89007 1 13520
2 89008 1 13520
2 89009 1 13520
2 89010 1 13536
2 89011 1 13536
2 89012 1 13538
2 89013 1 13538
2 89014 1 13549
2 89015 1 13549
2 89016 1 13549
2 89017 1 13550
2 89018 1 13550
2 89019 1 13553
2 89020 1 13553
2 89021 1 13577
2 89022 1 13577
2 89023 1 13577
2 89024 1 13577
2 89025 1 13577
2 89026 1 13578
2 89027 1 13578
2 89028 1 13578
2 89029 1 13580
2 89030 1 13580
2 89031 1 13580
2 89032 1 13580
2 89033 1 13587
2 89034 1 13587
2 89035 1 13587
2 89036 1 13602
2 89037 1 13602
2 89038 1 13603
2 89039 1 13603
2 89040 1 13603
2 89041 1 13603
2 89042 1 13609
2 89043 1 13609
2 89044 1 13609
2 89045 1 13609
2 89046 1 13609
2 89047 1 13609
2 89048 1 13610
2 89049 1 13610
2 89050 1 13610
2 89051 1 13610
2 89052 1 13610
2 89053 1 13610
2 89054 1 13610
2 89055 1 13613
2 89056 1 13613
2 89057 1 13613
2 89058 1 13613
2 89059 1 13613
2 89060 1 13613
2 89061 1 13613
2 89062 1 13613
2 89063 1 13614
2 89064 1 13614
2 89065 1 13614
2 89066 1 13614
2 89067 1 13644
2 89068 1 13644
2 89069 1 13644
2 89070 1 13644
2 89071 1 13644
2 89072 1 13645
2 89073 1 13645
2 89074 1 13656
2 89075 1 13656
2 89076 1 13660
2 89077 1 13660
2 89078 1 13661
2 89079 1 13661
2 89080 1 13661
2 89081 1 13670
2 89082 1 13670
2 89083 1 13676
2 89084 1 13676
2 89085 1 13679
2 89086 1 13679
2 89087 1 13679
2 89088 1 13679
2 89089 1 13700
2 89090 1 13700
2 89091 1 13704
2 89092 1 13704
2 89093 1 13714
2 89094 1 13714
2 89095 1 13714
2 89096 1 13714
2 89097 1 13714
2 89098 1 13715
2 89099 1 13715
2 89100 1 13715
2 89101 1 13715
2 89102 1 13715
2 89103 1 13715
2 89104 1 13715
2 89105 1 13715
2 89106 1 13715
2 89107 1 13715
2 89108 1 13717
2 89109 1 13717
2 89110 1 13717
2 89111 1 13719
2 89112 1 13719
2 89113 1 13727
2 89114 1 13727
2 89115 1 13738
2 89116 1 13738
2 89117 1 13740
2 89118 1 13740
2 89119 1 13754
2 89120 1 13754
2 89121 1 13755
2 89122 1 13755
2 89123 1 13762
2 89124 1 13762
2 89125 1 13762
2 89126 1 13762
2 89127 1 13762
2 89128 1 13764
2 89129 1 13764
2 89130 1 13764
2 89131 1 13764
2 89132 1 13773
2 89133 1 13773
2 89134 1 13774
2 89135 1 13774
2 89136 1 13774
2 89137 1 13794
2 89138 1 13794
2 89139 1 13799
2 89140 1 13799
2 89141 1 13802
2 89142 1 13802
2 89143 1 13802
2 89144 1 13802
2 89145 1 13802
2 89146 1 13802
2 89147 1 13802
2 89148 1 13803
2 89149 1 13803
2 89150 1 13806
2 89151 1 13806
2 89152 1 13810
2 89153 1 13810
2 89154 1 13810
2 89155 1 13820
2 89156 1 13820
2 89157 1 13820
2 89158 1 13821
2 89159 1 13821
2 89160 1 13821
2 89161 1 13821
2 89162 1 13822
2 89163 1 13822
2 89164 1 13822
2 89165 1 13822
2 89166 1 13824
2 89167 1 13824
2 89168 1 13825
2 89169 1 13825
2 89170 1 13826
2 89171 1 13826
2 89172 1 13827
2 89173 1 13827
2 89174 1 13837
2 89175 1 13837
2 89176 1 13853
2 89177 1 13853
2 89178 1 13866
2 89179 1 13866
2 89180 1 13866
2 89181 1 13866
2 89182 1 13866
2 89183 1 13866
2 89184 1 13866
2 89185 1 13867
2 89186 1 13867
2 89187 1 13867
2 89188 1 13868
2 89189 1 13868
2 89190 1 13868
2 89191 1 13869
2 89192 1 13869
2 89193 1 13869
2 89194 1 13869
2 89195 1 13870
2 89196 1 13870
2 89197 1 13873
2 89198 1 13873
2 89199 1 13873
2 89200 1 13877
2 89201 1 13877
2 89202 1 13877
2 89203 1 13877
2 89204 1 13878
2 89205 1 13878
2 89206 1 13882
2 89207 1 13882
2 89208 1 13882
2 89209 1 13882
2 89210 1 13883
2 89211 1 13883
2 89212 1 13883
2 89213 1 13883
2 89214 1 13883
2 89215 1 13895
2 89216 1 13895
2 89217 1 13895
2 89218 1 13895
2 89219 1 13896
2 89220 1 13896
2 89221 1 13929
2 89222 1 13929
2 89223 1 13929
2 89224 1 13929
2 89225 1 13930
2 89226 1 13930
2 89227 1 13931
2 89228 1 13931
2 89229 1 13939
2 89230 1 13939
2 89231 1 13940
2 89232 1 13940
2 89233 1 13940
2 89234 1 13942
2 89235 1 13942
2 89236 1 13943
2 89237 1 13943
2 89238 1 13943
2 89239 1 13947
2 89240 1 13947
2 89241 1 13967
2 89242 1 13967
2 89243 1 13967
2 89244 1 13974
2 89245 1 13974
2 89246 1 13978
2 89247 1 13978
2 89248 1 13978
2 89249 1 13978
2 89250 1 13978
2 89251 1 13981
2 89252 1 13981
2 89253 1 13981
2 89254 1 13981
2 89255 1 13981
2 89256 1 13981
2 89257 1 14003
2 89258 1 14003
2 89259 1 14016
2 89260 1 14016
2 89261 1 14016
2 89262 1 14027
2 89263 1 14027
2 89264 1 14027
2 89265 1 14027
2 89266 1 14027
2 89267 1 14028
2 89268 1 14028
2 89269 1 14028
2 89270 1 14063
2 89271 1 14063
2 89272 1 14076
2 89273 1 14076
2 89274 1 14077
2 89275 1 14077
2 89276 1 14077
2 89277 1 14092
2 89278 1 14092
2 89279 1 14113
2 89280 1 14113
2 89281 1 14113
2 89282 1 14123
2 89283 1 14123
2 89284 1 14142
2 89285 1 14142
2 89286 1 14142
2 89287 1 14142
2 89288 1 14145
2 89289 1 14145
2 89290 1 14160
2 89291 1 14160
2 89292 1 14161
2 89293 1 14161
2 89294 1 14162
2 89295 1 14162
2 89296 1 14162
2 89297 1 14162
2 89298 1 14171
2 89299 1 14171
2 89300 1 14172
2 89301 1 14172
2 89302 1 14172
2 89303 1 14172
2 89304 1 14172
2 89305 1 14175
2 89306 1 14175
2 89307 1 14176
2 89308 1 14176
2 89309 1 14177
2 89310 1 14177
2 89311 1 14177
2 89312 1 14177
2 89313 1 14177
2 89314 1 14177
2 89315 1 14177
2 89316 1 14177
2 89317 1 14177
2 89318 1 14177
2 89319 1 14177
2 89320 1 14177
2 89321 1 14177
2 89322 1 14177
2 89323 1 14177
2 89324 1 14177
2 89325 1 14177
2 89326 1 14177
2 89327 1 14177
2 89328 1 14177
2 89329 1 14177
2 89330 1 14177
2 89331 1 14177
2 89332 1 14177
2 89333 1 14178
2 89334 1 14178
2 89335 1 14178
2 89336 1 14178
2 89337 1 14178
2 89338 1 14178
2 89339 1 14178
2 89340 1 14178
2 89341 1 14179
2 89342 1 14179
2 89343 1 14180
2 89344 1 14180
2 89345 1 14180
2 89346 1 14180
2 89347 1 14182
2 89348 1 14182
2 89349 1 14182
2 89350 1 14192
2 89351 1 14192
2 89352 1 14192
2 89353 1 14192
2 89354 1 14192
2 89355 1 14192
2 89356 1 14192
2 89357 1 14192
2 89358 1 14194
2 89359 1 14194
2 89360 1 14195
2 89361 1 14195
2 89362 1 14196
2 89363 1 14196
2 89364 1 14196
2 89365 1 14196
2 89366 1 14196
2 89367 1 14196
2 89368 1 14198
2 89369 1 14198
2 89370 1 14205
2 89371 1 14205
2 89372 1 14205
2 89373 1 14206
2 89374 1 14206
2 89375 1 14209
2 89376 1 14209
2 89377 1 14214
2 89378 1 14214
2 89379 1 14216
2 89380 1 14216
2 89381 1 14216
2 89382 1 14216
2 89383 1 14217
2 89384 1 14217
2 89385 1 14217
2 89386 1 14217
2 89387 1 14219
2 89388 1 14219
2 89389 1 14219
2 89390 1 14225
2 89391 1 14225
2 89392 1 14253
2 89393 1 14253
2 89394 1 14253
2 89395 1 14254
2 89396 1 14254
2 89397 1 14257
2 89398 1 14257
2 89399 1 14257
2 89400 1 14257
2 89401 1 14257
2 89402 1 14257
2 89403 1 14257
2 89404 1 14257
2 89405 1 14257
2 89406 1 14257
2 89407 1 14257
2 89408 1 14258
2 89409 1 14258
2 89410 1 14258
2 89411 1 14258
2 89412 1 14258
2 89413 1 14258
2 89414 1 14260
2 89415 1 14260
2 89416 1 14261
2 89417 1 14261
2 89418 1 14261
2 89419 1 14264
2 89420 1 14264
2 89421 1 14267
2 89422 1 14267
2 89423 1 14267
2 89424 1 14269
2 89425 1 14269
2 89426 1 14276
2 89427 1 14276
2 89428 1 14276
2 89429 1 14276
2 89430 1 14289
2 89431 1 14289
2 89432 1 14291
2 89433 1 14291
2 89434 1 14301
2 89435 1 14301
2 89436 1 14301
2 89437 1 14301
2 89438 1 14301
2 89439 1 14303
2 89440 1 14303
2 89441 1 14303
2 89442 1 14304
2 89443 1 14304
2 89444 1 14304
2 89445 1 14305
2 89446 1 14305
2 89447 1 14307
2 89448 1 14307
2 89449 1 14316
2 89450 1 14316
2 89451 1 14316
2 89452 1 14316
2 89453 1 14316
2 89454 1 14316
2 89455 1 14317
2 89456 1 14317
2 89457 1 14317
2 89458 1 14318
2 89459 1 14318
2 89460 1 14318
2 89461 1 14318
2 89462 1 14321
2 89463 1 14321
2 89464 1 14329
2 89465 1 14329
2 89466 1 14329
2 89467 1 14331
2 89468 1 14331
2 89469 1 14342
2 89470 1 14342
2 89471 1 14342
2 89472 1 14342
2 89473 1 14342
2 89474 1 14342
2 89475 1 14343
2 89476 1 14343
2 89477 1 14343
2 89478 1 14343
2 89479 1 14344
2 89480 1 14344
2 89481 1 14344
2 89482 1 14344
2 89483 1 14344
2 89484 1 14344
2 89485 1 14344
2 89486 1 14344
2 89487 1 14344
2 89488 1 14344
2 89489 1 14344
2 89490 1 14344
2 89491 1 14344
2 89492 1 14344
2 89493 1 14345
2 89494 1 14345
2 89495 1 14347
2 89496 1 14347
2 89497 1 14347
2 89498 1 14360
2 89499 1 14360
2 89500 1 14371
2 89501 1 14371
2 89502 1 14371
2 89503 1 14371
2 89504 1 14371
2 89505 1 14371
2 89506 1 14371
2 89507 1 14372
2 89508 1 14372
2 89509 1 14372
2 89510 1 14372
2 89511 1 14372
2 89512 1 14372
2 89513 1 14373
2 89514 1 14373
2 89515 1 14373
2 89516 1 14382
2 89517 1 14382
2 89518 1 14382
2 89519 1 14382
2 89520 1 14382
2 89521 1 14382
2 89522 1 14382
2 89523 1 14382
2 89524 1 14382
2 89525 1 14383
2 89526 1 14383
2 89527 1 14383
2 89528 1 14383
2 89529 1 14383
2 89530 1 14383
2 89531 1 14421
2 89532 1 14421
2 89533 1 14421
2 89534 1 14422
2 89535 1 14422
2 89536 1 14422
2 89537 1 14422
2 89538 1 14422
2 89539 1 14422
2 89540 1 14444
2 89541 1 14444
2 89542 1 14444
2 89543 1 14445
2 89544 1 14445
2 89545 1 14445
2 89546 1 14445
2 89547 1 14445
2 89548 1 14458
2 89549 1 14458
2 89550 1 14458
2 89551 1 14458
2 89552 1 14458
2 89553 1 14459
2 89554 1 14459
2 89555 1 14459
2 89556 1 14459
2 89557 1 14459
2 89558 1 14460
2 89559 1 14460
2 89560 1 14460
2 89561 1 14460
2 89562 1 14460
2 89563 1 14461
2 89564 1 14461
2 89565 1 14461
2 89566 1 14461
2 89567 1 14463
2 89568 1 14463
2 89569 1 14465
2 89570 1 14465
2 89571 1 14467
2 89572 1 14467
2 89573 1 14473
2 89574 1 14473
2 89575 1 14474
2 89576 1 14474
2 89577 1 14476
2 89578 1 14476
2 89579 1 14476
2 89580 1 14476
2 89581 1 14493
2 89582 1 14493
2 89583 1 14493
2 89584 1 14494
2 89585 1 14494
2 89586 1 14494
2 89587 1 14494
2 89588 1 14494
2 89589 1 14494
2 89590 1 14494
2 89591 1 14495
2 89592 1 14495
2 89593 1 14495
2 89594 1 14502
2 89595 1 14502
2 89596 1 14508
2 89597 1 14508
2 89598 1 14511
2 89599 1 14511
2 89600 1 14512
2 89601 1 14512
2 89602 1 14512
2 89603 1 14513
2 89604 1 14513
2 89605 1 14513
2 89606 1 14528
2 89607 1 14528
2 89608 1 14529
2 89609 1 14529
2 89610 1 14530
2 89611 1 14530
2 89612 1 14530
2 89613 1 14530
2 89614 1 14552
2 89615 1 14552
2 89616 1 14561
2 89617 1 14561
2 89618 1 14562
2 89619 1 14562
2 89620 1 14563
2 89621 1 14563
2 89622 1 14568
2 89623 1 14568
2 89624 1 14569
2 89625 1 14569
2 89626 1 14569
2 89627 1 14569
2 89628 1 14569
2 89629 1 14571
2 89630 1 14571
2 89631 1 14578
2 89632 1 14578
2 89633 1 14600
2 89634 1 14600
2 89635 1 14618
2 89636 1 14618
2 89637 1 14618
2 89638 1 14618
2 89639 1 14618
2 89640 1 14627
2 89641 1 14627
2 89642 1 14627
2 89643 1 14627
2 89644 1 14627
2 89645 1 14628
2 89646 1 14628
2 89647 1 14628
2 89648 1 14628
2 89649 1 14628
2 89650 1 14628
2 89651 1 14629
2 89652 1 14629
2 89653 1 14635
2 89654 1 14635
2 89655 1 14652
2 89656 1 14652
2 89657 1 14652
2 89658 1 14652
2 89659 1 14670
2 89660 1 14670
2 89661 1 14670
2 89662 1 14671
2 89663 1 14671
2 89664 1 14684
2 89665 1 14684
2 89666 1 14685
2 89667 1 14685
2 89668 1 14686
2 89669 1 14686
2 89670 1 14690
2 89671 1 14690
2 89672 1 14711
2 89673 1 14711
2 89674 1 14712
2 89675 1 14712
2 89676 1 14712
2 89677 1 14726
2 89678 1 14726
2 89679 1 14727
2 89680 1 14727
2 89681 1 14728
2 89682 1 14728
2 89683 1 14728
2 89684 1 14728
2 89685 1 14728
2 89686 1 14728
2 89687 1 14728
2 89688 1 14728
2 89689 1 14728
2 89690 1 14728
2 89691 1 14728
2 89692 1 14728
2 89693 1 14728
2 89694 1 14728
2 89695 1 14728
2 89696 1 14728
2 89697 1 14728
2 89698 1 14729
2 89699 1 14729
2 89700 1 14732
2 89701 1 14732
2 89702 1 14732
2 89703 1 14732
2 89704 1 14732
2 89705 1 14732
2 89706 1 14732
2 89707 1 14732
2 89708 1 14732
2 89709 1 14732
2 89710 1 14732
2 89711 1 14732
2 89712 1 14732
2 89713 1 14732
2 89714 1 14732
2 89715 1 14732
2 89716 1 14732
2 89717 1 14743
2 89718 1 14743
2 89719 1 14743
2 89720 1 14743
2 89721 1 14743
2 89722 1 14743
2 89723 1 14743
2 89724 1 14744
2 89725 1 14744
2 89726 1 14747
2 89727 1 14747
2 89728 1 14747
2 89729 1 14756
2 89730 1 14756
2 89731 1 14759
2 89732 1 14759
2 89733 1 14770
2 89734 1 14770
2 89735 1 14770
2 89736 1 14777
2 89737 1 14777
2 89738 1 14778
2 89739 1 14778
2 89740 1 14778
2 89741 1 14778
2 89742 1 14778
2 89743 1 14778
2 89744 1 14780
2 89745 1 14780
2 89746 1 14780
2 89747 1 14792
2 89748 1 14792
2 89749 1 14792
2 89750 1 14792
2 89751 1 14792
2 89752 1 14792
2 89753 1 14792
2 89754 1 14792
2 89755 1 14793
2 89756 1 14793
2 89757 1 14801
2 89758 1 14801
2 89759 1 14817
2 89760 1 14817
2 89761 1 14817
2 89762 1 14834
2 89763 1 14834
2 89764 1 14834
2 89765 1 14834
2 89766 1 14834
2 89767 1 14834
2 89768 1 14834
2 89769 1 14834
2 89770 1 14834
2 89771 1 14834
2 89772 1 14834
2 89773 1 14834
2 89774 1 14834
2 89775 1 14834
2 89776 1 14834
2 89777 1 14834
2 89778 1 14834
2 89779 1 14834
2 89780 1 14834
2 89781 1 14848
2 89782 1 14848
2 89783 1 14848
2 89784 1 14856
2 89785 1 14856
2 89786 1 14856
2 89787 1 14864
2 89788 1 14864
2 89789 1 14866
2 89790 1 14866
2 89791 1 14866
2 89792 1 14866
2 89793 1 14866
2 89794 1 14866
2 89795 1 14867
2 89796 1 14867
2 89797 1 14867
2 89798 1 14868
2 89799 1 14868
2 89800 1 14868
2 89801 1 14878
2 89802 1 14878
2 89803 1 14880
2 89804 1 14880
2 89805 1 14890
2 89806 1 14890
2 89807 1 14905
2 89808 1 14905
2 89809 1 14905
2 89810 1 14905
2 89811 1 14905
2 89812 1 14905
2 89813 1 14905
2 89814 1 14905
2 89815 1 14905
2 89816 1 14905
2 89817 1 14905
2 89818 1 14905
2 89819 1 14905
2 89820 1 14905
2 89821 1 14905
2 89822 1 14905
2 89823 1 14905
2 89824 1 14913
2 89825 1 14913
2 89826 1 14913
2 89827 1 14928
2 89828 1 14928
2 89829 1 14929
2 89830 1 14929
2 89831 1 14929
2 89832 1 14930
2 89833 1 14930
2 89834 1 14930
2 89835 1 14930
2 89836 1 14930
2 89837 1 14930
2 89838 1 14931
2 89839 1 14931
2 89840 1 14932
2 89841 1 14932
2 89842 1 14945
2 89843 1 14945
2 89844 1 14946
2 89845 1 14946
2 89846 1 14948
2 89847 1 14948
2 89848 1 14948
2 89849 1 14956
2 89850 1 14956
2 89851 1 14966
2 89852 1 14966
2 89853 1 14966
2 89854 1 14967
2 89855 1 14967
2 89856 1 14975
2 89857 1 14975
2 89858 1 14975
2 89859 1 14975
2 89860 1 14975
2 89861 1 14975
2 89862 1 14976
2 89863 1 14976
2 89864 1 14976
2 89865 1 14998
2 89866 1 14998
2 89867 1 15007
2 89868 1 15007
2 89869 1 15016
2 89870 1 15016
2 89871 1 15017
2 89872 1 15017
2 89873 1 15017
2 89874 1 15017
2 89875 1 15017
2 89876 1 15017
2 89877 1 15017
2 89878 1 15017
2 89879 1 15017
2 89880 1 15018
2 89881 1 15018
2 89882 1 15022
2 89883 1 15022
2 89884 1 15022
2 89885 1 15023
2 89886 1 15023
2 89887 1 15030
2 89888 1 15030
2 89889 1 15030
2 89890 1 15045
2 89891 1 15045
2 89892 1 15075
2 89893 1 15075
2 89894 1 15080
2 89895 1 15080
2 89896 1 15080
2 89897 1 15080
2 89898 1 15080
2 89899 1 15080
2 89900 1 15080
2 89901 1 15081
2 89902 1 15081
2 89903 1 15083
2 89904 1 15083
2 89905 1 15083
2 89906 1 15101
2 89907 1 15101
2 89908 1 15102
2 89909 1 15102
2 89910 1 15102
2 89911 1 15104
2 89912 1 15104
2 89913 1 15111
2 89914 1 15111
2 89915 1 15119
2 89916 1 15119
2 89917 1 15119
2 89918 1 15128
2 89919 1 15128
2 89920 1 15137
2 89921 1 15137
2 89922 1 15137
2 89923 1 15137
2 89924 1 15137
2 89925 1 15137
2 89926 1 15137
2 89927 1 15137
2 89928 1 15137
2 89929 1 15137
2 89930 1 15137
2 89931 1 15137
2 89932 1 15137
2 89933 1 15137
2 89934 1 15137
2 89935 1 15137
2 89936 1 15137
2 89937 1 15137
2 89938 1 15137
2 89939 1 15137
2 89940 1 15137
2 89941 1 15137
2 89942 1 15137
2 89943 1 15137
2 89944 1 15137
2 89945 1 15137
2 89946 1 15138
2 89947 1 15138
2 89948 1 15138
2 89949 1 15138
2 89950 1 15138
2 89951 1 15138
2 89952 1 15138
2 89953 1 15138
2 89954 1 15139
2 89955 1 15139
2 89956 1 15139
2 89957 1 15139
2 89958 1 15139
2 89959 1 15139
2 89960 1 15148
2 89961 1 15148
2 89962 1 15156
2 89963 1 15156
2 89964 1 15156
2 89965 1 15156
2 89966 1 15156
2 89967 1 15156
2 89968 1 15157
2 89969 1 15157
2 89970 1 15165
2 89971 1 15165
2 89972 1 15165
2 89973 1 15165
2 89974 1 15165
2 89975 1 15165
2 89976 1 15165
2 89977 1 15166
2 89978 1 15166
2 89979 1 15166
2 89980 1 15167
2 89981 1 15167
2 89982 1 15184
2 89983 1 15184
2 89984 1 15184
2 89985 1 15187
2 89986 1 15187
2 89987 1 15190
2 89988 1 15190
2 89989 1 15190
2 89990 1 15202
2 89991 1 15202
2 89992 1 15206
2 89993 1 15206
2 89994 1 15214
2 89995 1 15214
2 89996 1 15223
2 89997 1 15223
2 89998 1 15223
2 89999 1 15223
2 90000 1 15242
2 90001 1 15242
2 90002 1 15275
2 90003 1 15275
2 90004 1 15275
2 90005 1 15290
2 90006 1 15290
2 90007 1 15290
2 90008 1 15290
2 90009 1 15290
2 90010 1 15292
2 90011 1 15292
2 90012 1 15301
2 90013 1 15301
2 90014 1 15301
2 90015 1 15301
2 90016 1 15302
2 90017 1 15302
2 90018 1 15302
2 90019 1 15316
2 90020 1 15316
2 90021 1 15316
2 90022 1 15316
2 90023 1 15316
2 90024 1 15319
2 90025 1 15319
2 90026 1 15334
2 90027 1 15334
2 90028 1 15343
2 90029 1 15343
2 90030 1 15343
2 90031 1 15344
2 90032 1 15344
2 90033 1 15345
2 90034 1 15345
2 90035 1 15345
2 90036 1 15345
2 90037 1 15345
2 90038 1 15345
2 90039 1 15346
2 90040 1 15346
2 90041 1 15346
2 90042 1 15346
2 90043 1 15346
2 90044 1 15346
2 90045 1 15346
2 90046 1 15349
2 90047 1 15349
2 90048 1 15377
2 90049 1 15377
2 90050 1 15378
2 90051 1 15378
2 90052 1 15386
2 90053 1 15386
2 90054 1 15390
2 90055 1 15390
2 90056 1 15394
2 90057 1 15394
2 90058 1 15394
2 90059 1 15394
2 90060 1 15394
2 90061 1 15394
2 90062 1 15394
2 90063 1 15412
2 90064 1 15412
2 90065 1 15412
2 90066 1 15412
2 90067 1 15412
2 90068 1 15412
2 90069 1 15412
2 90070 1 15412
2 90071 1 15412
2 90072 1 15412
2 90073 1 15413
2 90074 1 15413
2 90075 1 15413
2 90076 1 15414
2 90077 1 15414
2 90078 1 15415
2 90079 1 15415
2 90080 1 15419
2 90081 1 15419
2 90082 1 15419
2 90083 1 15423
2 90084 1 15423
2 90085 1 15426
2 90086 1 15426
2 90087 1 15429
2 90088 1 15429
2 90089 1 15437
2 90090 1 15437
2 90091 1 15444
2 90092 1 15444
2 90093 1 15460
2 90094 1 15460
2 90095 1 15461
2 90096 1 15461
2 90097 1 15461
2 90098 1 15461
2 90099 1 15461
2 90100 1 15471
2 90101 1 15471
2 90102 1 15471
2 90103 1 15473
2 90104 1 15473
2 90105 1 15473
2 90106 1 15477
2 90107 1 15477
2 90108 1 15477
2 90109 1 15477
2 90110 1 15477
2 90111 1 15477
2 90112 1 15477
2 90113 1 15477
2 90114 1 15477
2 90115 1 15477
2 90116 1 15477
2 90117 1 15477
2 90118 1 15477
2 90119 1 15478
2 90120 1 15478
2 90121 1 15478
2 90122 1 15478
2 90123 1 15478
2 90124 1 15478
2 90125 1 15478
2 90126 1 15478
2 90127 1 15478
2 90128 1 15478
2 90129 1 15478
2 90130 1 15478
2 90131 1 15479
2 90132 1 15479
2 90133 1 15479
2 90134 1 15480
2 90135 1 15480
2 90136 1 15480
2 90137 1 15485
2 90138 1 15485
2 90139 1 15485
2 90140 1 15485
2 90141 1 15485
2 90142 1 15485
2 90143 1 15485
2 90144 1 15485
2 90145 1 15485
2 90146 1 15485
2 90147 1 15485
2 90148 1 15486
2 90149 1 15486
2 90150 1 15496
2 90151 1 15496
2 90152 1 15498
2 90153 1 15498
2 90154 1 15498
2 90155 1 15498
2 90156 1 15498
2 90157 1 15498
2 90158 1 15498
2 90159 1 15498
2 90160 1 15498
2 90161 1 15498
2 90162 1 15498
2 90163 1 15498
2 90164 1 15500
2 90165 1 15500
2 90166 1 15500
2 90167 1 15510
2 90168 1 15510
2 90169 1 15516
2 90170 1 15516
2 90171 1 15516
2 90172 1 15516
2 90173 1 15516
2 90174 1 15516
2 90175 1 15516
2 90176 1 15516
2 90177 1 15516
2 90178 1 15516
2 90179 1 15516
2 90180 1 15516
2 90181 1 15516
2 90182 1 15516
2 90183 1 15516
2 90184 1 15516
2 90185 1 15516
2 90186 1 15516
2 90187 1 15517
2 90188 1 15517
2 90189 1 15518
2 90190 1 15518
2 90191 1 15519
2 90192 1 15519
2 90193 1 15519
2 90194 1 15519
2 90195 1 15519
2 90196 1 15519
2 90197 1 15519
2 90198 1 15519
2 90199 1 15519
2 90200 1 15519
2 90201 1 15519
2 90202 1 15519
2 90203 1 15519
2 90204 1 15519
2 90205 1 15519
2 90206 1 15519
2 90207 1 15519
2 90208 1 15519
2 90209 1 15519
2 90210 1 15519
2 90211 1 15519
2 90212 1 15521
2 90213 1 15521
2 90214 1 15521
2 90215 1 15521
2 90216 1 15521
2 90217 1 15521
2 90218 1 15545
2 90219 1 15545
2 90220 1 15553
2 90221 1 15553
2 90222 1 15556
2 90223 1 15556
2 90224 1 15556
2 90225 1 15557
2 90226 1 15557
2 90227 1 15563
2 90228 1 15563
2 90229 1 15568
2 90230 1 15568
2 90231 1 15569
2 90232 1 15569
2 90233 1 15571
2 90234 1 15571
2 90235 1 15576
2 90236 1 15576
2 90237 1 15578
2 90238 1 15578
2 90239 1 15583
2 90240 1 15583
2 90241 1 15584
2 90242 1 15584
2 90243 1 15584
2 90244 1 15591
2 90245 1 15591
2 90246 1 15591
2 90247 1 15591
2 90248 1 15591
2 90249 1 15604
2 90250 1 15604
2 90251 1 15618
2 90252 1 15618
2 90253 1 15619
2 90254 1 15619
2 90255 1 15625
2 90256 1 15625
2 90257 1 15635
2 90258 1 15635
2 90259 1 15642
2 90260 1 15642
2 90261 1 15645
2 90262 1 15645
2 90263 1 15645
2 90264 1 15645
2 90265 1 15645
2 90266 1 15646
2 90267 1 15646
2 90268 1 15646
2 90269 1 15646
2 90270 1 15646
2 90271 1 15646
2 90272 1 15648
2 90273 1 15648
2 90274 1 15648
2 90275 1 15649
2 90276 1 15649
2 90277 1 15650
2 90278 1 15650
2 90279 1 15652
2 90280 1 15652
2 90281 1 15667
2 90282 1 15667
2 90283 1 15667
2 90284 1 15667
2 90285 1 15670
2 90286 1 15670
2 90287 1 15670
2 90288 1 15671
2 90289 1 15671
2 90290 1 15678
2 90291 1 15678
2 90292 1 15687
2 90293 1 15687
2 90294 1 15687
2 90295 1 15688
2 90296 1 15688
2 90297 1 15720
2 90298 1 15720
2 90299 1 15733
2 90300 1 15733
2 90301 1 15733
2 90302 1 15734
2 90303 1 15734
2 90304 1 15735
2 90305 1 15735
2 90306 1 15738
2 90307 1 15738
2 90308 1 15738
2 90309 1 15753
2 90310 1 15753
2 90311 1 15753
2 90312 1 15767
2 90313 1 15767
2 90314 1 15767
2 90315 1 15771
2 90316 1 15771
2 90317 1 15771
2 90318 1 15771
2 90319 1 15774
2 90320 1 15774
2 90321 1 15786
2 90322 1 15786
2 90323 1 15786
2 90324 1 15787
2 90325 1 15787
2 90326 1 15798
2 90327 1 15798
2 90328 1 15798
2 90329 1 15798
2 90330 1 15798
2 90331 1 15798
2 90332 1 15798
2 90333 1 15799
2 90334 1 15799
2 90335 1 15802
2 90336 1 15802
2 90337 1 15802
2 90338 1 15822
2 90339 1 15822
2 90340 1 15822
2 90341 1 15838
2 90342 1 15838
2 90343 1 15838
2 90344 1 15838
2 90345 1 15838
2 90346 1 15839
2 90347 1 15839
2 90348 1 15839
2 90349 1 15856
2 90350 1 15856
2 90351 1 15860
2 90352 1 15860
2 90353 1 15867
2 90354 1 15867
2 90355 1 15886
2 90356 1 15886
2 90357 1 15887
2 90358 1 15887
2 90359 1 15888
2 90360 1 15888
2 90361 1 15888
2 90362 1 15888
2 90363 1 15888
2 90364 1 15889
2 90365 1 15889
2 90366 1 15897
2 90367 1 15897
2 90368 1 15907
2 90369 1 15907
2 90370 1 15908
2 90371 1 15908
2 90372 1 15908
2 90373 1 15930
2 90374 1 15930
2 90375 1 15930
2 90376 1 15930
2 90377 1 15931
2 90378 1 15931
2 90379 1 15931
2 90380 1 15943
2 90381 1 15943
2 90382 1 15943
2 90383 1 15943
2 90384 1 15943
2 90385 1 15943
2 90386 1 15943
2 90387 1 15943
2 90388 1 15944
2 90389 1 15944
2 90390 1 15944
2 90391 1 15945
2 90392 1 15945
2 90393 1 15947
2 90394 1 15947
2 90395 1 15950
2 90396 1 15950
2 90397 1 15950
2 90398 1 15950
2 90399 1 15962
2 90400 1 15962
2 90401 1 15969
2 90402 1 15969
2 90403 1 15969
2 90404 1 15970
2 90405 1 15970
2 90406 1 15971
2 90407 1 15971
2 90408 1 15972
2 90409 1 15972
2 90410 1 15972
2 90411 1 15974
2 90412 1 15974
2 90413 1 15974
2 90414 1 15990
2 90415 1 15990
2 90416 1 15993
2 90417 1 15993
2 90418 1 16002
2 90419 1 16002
2 90420 1 16003
2 90421 1 16003
2 90422 1 16012
2 90423 1 16012
2 90424 1 16021
2 90425 1 16021
2 90426 1 16034
2 90427 1 16034
2 90428 1 16036
2 90429 1 16036
2 90430 1 16038
2 90431 1 16038
2 90432 1 16038
2 90433 1 16038
2 90434 1 16038
2 90435 1 16038
2 90436 1 16039
2 90437 1 16039
2 90438 1 16039
2 90439 1 16039
2 90440 1 16040
2 90441 1 16040
2 90442 1 16040
2 90443 1 16041
2 90444 1 16041
2 90445 1 16041
2 90446 1 16060
2 90447 1 16060
2 90448 1 16060
2 90449 1 16061
2 90450 1 16061
2 90451 1 16061
2 90452 1 16074
2 90453 1 16074
2 90454 1 16075
2 90455 1 16075
2 90456 1 16076
2 90457 1 16076
2 90458 1 16079
2 90459 1 16079
2 90460 1 16079
2 90461 1 16113
2 90462 1 16113
2 90463 1 16113
2 90464 1 16113
2 90465 1 16113
2 90466 1 16116
2 90467 1 16116
2 90468 1 16116
2 90469 1 16132
2 90470 1 16132
2 90471 1 16133
2 90472 1 16133
2 90473 1 16133
2 90474 1 16149
2 90475 1 16149
2 90476 1 16153
2 90477 1 16153
2 90478 1 16153
2 90479 1 16153
2 90480 1 16179
2 90481 1 16179
2 90482 1 16195
2 90483 1 16195
2 90484 1 16206
2 90485 1 16206
2 90486 1 16206
2 90487 1 16211
2 90488 1 16211
2 90489 1 16228
2 90490 1 16228
2 90491 1 16228
2 90492 1 16228
2 90493 1 16228
2 90494 1 16229
2 90495 1 16229
2 90496 1 16229
2 90497 1 16229
2 90498 1 16229
2 90499 1 16229
2 90500 1 16229
2 90501 1 16229
2 90502 1 16229
2 90503 1 16229
2 90504 1 16229
2 90505 1 16229
2 90506 1 16229
2 90507 1 16229
2 90508 1 16229
2 90509 1 16237
2 90510 1 16237
2 90511 1 16242
2 90512 1 16242
2 90513 1 16242
2 90514 1 16243
2 90515 1 16243
2 90516 1 16243
2 90517 1 16248
2 90518 1 16248
2 90519 1 16249
2 90520 1 16249
2 90521 1 16250
2 90522 1 16250
2 90523 1 16262
2 90524 1 16262
2 90525 1 16264
2 90526 1 16264
2 90527 1 16265
2 90528 1 16265
2 90529 1 16266
2 90530 1 16266
2 90531 1 16269
2 90532 1 16269
2 90533 1 16279
2 90534 1 16279
2 90535 1 16280
2 90536 1 16280
2 90537 1 16280
2 90538 1 16281
2 90539 1 16281
2 90540 1 16282
2 90541 1 16282
2 90542 1 16282
2 90543 1 16287
2 90544 1 16287
2 90545 1 16294
2 90546 1 16294
2 90547 1 16295
2 90548 1 16295
2 90549 1 16300
2 90550 1 16300
2 90551 1 16300
2 90552 1 16311
2 90553 1 16311
2 90554 1 16315
2 90555 1 16315
2 90556 1 16330
2 90557 1 16330
2 90558 1 16330
2 90559 1 16336
2 90560 1 16336
2 90561 1 16344
2 90562 1 16344
2 90563 1 16350
2 90564 1 16350
2 90565 1 16363
2 90566 1 16363
2 90567 1 16364
2 90568 1 16364
2 90569 1 16365
2 90570 1 16365
2 90571 1 16365
2 90572 1 16365
2 90573 1 16369
2 90574 1 16369
2 90575 1 16372
2 90576 1 16372
2 90577 1 16372
2 90578 1 16372
2 90579 1 16372
2 90580 1 16373
2 90581 1 16373
2 90582 1 16375
2 90583 1 16375
2 90584 1 16384
2 90585 1 16384
2 90586 1 16387
2 90587 1 16387
2 90588 1 16396
2 90589 1 16396
2 90590 1 16396
2 90591 1 16396
2 90592 1 16396
2 90593 1 16408
2 90594 1 16408
2 90595 1 16419
2 90596 1 16419
2 90597 1 16419
2 90598 1 16419
2 90599 1 16419
2 90600 1 16419
2 90601 1 16419
2 90602 1 16419
2 90603 1 16419
2 90604 1 16419
2 90605 1 16419
2 90606 1 16419
2 90607 1 16419
2 90608 1 16419
2 90609 1 16419
2 90610 1 16419
2 90611 1 16419
2 90612 1 16419
2 90613 1 16419
2 90614 1 16419
2 90615 1 16419
2 90616 1 16420
2 90617 1 16420
2 90618 1 16420
2 90619 1 16420
2 90620 1 16420
2 90621 1 16420
2 90622 1 16420
2 90623 1 16421
2 90624 1 16421
2 90625 1 16456
2 90626 1 16456
2 90627 1 16475
2 90628 1 16475
2 90629 1 16475
2 90630 1 16475
2 90631 1 16475
2 90632 1 16479
2 90633 1 16479
2 90634 1 16479
2 90635 1 16479
2 90636 1 16479
2 90637 1 16479
2 90638 1 16479
2 90639 1 16479
2 90640 1 16479
2 90641 1 16479
2 90642 1 16479
2 90643 1 16479
2 90644 1 16479
2 90645 1 16479
2 90646 1 16491
2 90647 1 16491
2 90648 1 16491
2 90649 1 16519
2 90650 1 16519
2 90651 1 16519
2 90652 1 16520
2 90653 1 16520
2 90654 1 16520
2 90655 1 16521
2 90656 1 16521
2 90657 1 16522
2 90658 1 16522
2 90659 1 16524
2 90660 1 16524
2 90661 1 16524
2 90662 1 16524
2 90663 1 16538
2 90664 1 16538
2 90665 1 16546
2 90666 1 16546
2 90667 1 16553
2 90668 1 16553
2 90669 1 16558
2 90670 1 16558
2 90671 1 16565
2 90672 1 16565
2 90673 1 16582
2 90674 1 16582
2 90675 1 16585
2 90676 1 16585
2 90677 1 16585
2 90678 1 16585
2 90679 1 16588
2 90680 1 16588
2 90681 1 16589
2 90682 1 16589
2 90683 1 16589
2 90684 1 16590
2 90685 1 16590
2 90686 1 16592
2 90687 1 16592
2 90688 1 16592
2 90689 1 16605
2 90690 1 16605
2 90691 1 16637
2 90692 1 16637
2 90693 1 16637
2 90694 1 16637
2 90695 1 16637
2 90696 1 16646
2 90697 1 16646
2 90698 1 16646
2 90699 1 16651
2 90700 1 16651
2 90701 1 16652
2 90702 1 16652
2 90703 1 16663
2 90704 1 16663
2 90705 1 16663
2 90706 1 16664
2 90707 1 16664
2 90708 1 16665
2 90709 1 16665
2 90710 1 16675
2 90711 1 16675
2 90712 1 16684
2 90713 1 16684
2 90714 1 16684
2 90715 1 16684
2 90716 1 16684
2 90717 1 16685
2 90718 1 16685
2 90719 1 16710
2 90720 1 16710
2 90721 1 16710
2 90722 1 16710
2 90723 1 16710
2 90724 1 16711
2 90725 1 16711
2 90726 1 16715
2 90727 1 16715
2 90728 1 16715
2 90729 1 16718
2 90730 1 16718
2 90731 1 16718
2 90732 1 16719
2 90733 1 16719
2 90734 1 16719
2 90735 1 16733
2 90736 1 16733
2 90737 1 16734
2 90738 1 16734
2 90739 1 16734
2 90740 1 16734
2 90741 1 16785
2 90742 1 16785
2 90743 1 16799
2 90744 1 16799
2 90745 1 16814
2 90746 1 16814
2 90747 1 16814
2 90748 1 16815
2 90749 1 16815
2 90750 1 16817
2 90751 1 16817
2 90752 1 16822
2 90753 1 16822
2 90754 1 16835
2 90755 1 16835
2 90756 1 16851
2 90757 1 16851
2 90758 1 16865
2 90759 1 16865
2 90760 1 16866
2 90761 1 16866
2 90762 1 16866
2 90763 1 16867
2 90764 1 16867
2 90765 1 16867
2 90766 1 16867
2 90767 1 16867
2 90768 1 16867
2 90769 1 16867
2 90770 1 16867
2 90771 1 16867
2 90772 1 16867
2 90773 1 16867
2 90774 1 16867
2 90775 1 16867
2 90776 1 16867
2 90777 1 16867
2 90778 1 16867
2 90779 1 16867
2 90780 1 16867
2 90781 1 16867
2 90782 1 16867
2 90783 1 16868
2 90784 1 16868
2 90785 1 16868
2 90786 1 16869
2 90787 1 16869
2 90788 1 16877
2 90789 1 16877
2 90790 1 16877
2 90791 1 16877
2 90792 1 16877
2 90793 1 16878
2 90794 1 16878
2 90795 1 16880
2 90796 1 16880
2 90797 1 16880
2 90798 1 16880
2 90799 1 16892
2 90800 1 16892
2 90801 1 16892
2 90802 1 16897
2 90803 1 16897
2 90804 1 16917
2 90805 1 16917
2 90806 1 16917
2 90807 1 16917
2 90808 1 16917
2 90809 1 16930
2 90810 1 16930
2 90811 1 16930
2 90812 1 16930
2 90813 1 16931
2 90814 1 16931
2 90815 1 16960
2 90816 1 16960
2 90817 1 16973
2 90818 1 16973
2 90819 1 16982
2 90820 1 16982
2 90821 1 16983
2 90822 1 16983
2 90823 1 16992
2 90824 1 16992
2 90825 1 17002
2 90826 1 17002
2 90827 1 17058
2 90828 1 17058
2 90829 1 17058
2 90830 1 17060
2 90831 1 17060
2 90832 1 17107
2 90833 1 17107
2 90834 1 17115
2 90835 1 17115
2 90836 1 17115
2 90837 1 17162
2 90838 1 17162
2 90839 1 17163
2 90840 1 17163
2 90841 1 17172
2 90842 1 17172
2 90843 1 17173
2 90844 1 17173
2 90845 1 17178
2 90846 1 17178
2 90847 1 17182
2 90848 1 17182
2 90849 1 17191
2 90850 1 17191
2 90851 1 17209
2 90852 1 17209
2 90853 1 17221
2 90854 1 17221
2 90855 1 17228
2 90856 1 17228
2 90857 1 17229
2 90858 1 17229
2 90859 1 17229
2 90860 1 17229
2 90861 1 17229
2 90862 1 17230
2 90863 1 17230
2 90864 1 17230
2 90865 1 17230
2 90866 1 17258
2 90867 1 17258
2 90868 1 17259
2 90869 1 17259
2 90870 1 17260
2 90871 1 17260
2 90872 1 17260
2 90873 1 17260
2 90874 1 17261
2 90875 1 17261
2 90876 1 17261
2 90877 1 17261
2 90878 1 17261
2 90879 1 17261
2 90880 1 17264
2 90881 1 17264
2 90882 1 17265
2 90883 1 17265
2 90884 1 17279
2 90885 1 17279
2 90886 1 17283
2 90887 1 17283
2 90888 1 17289
2 90889 1 17289
2 90890 1 17305
2 90891 1 17305
2 90892 1 17311
2 90893 1 17311
2 90894 1 17311
2 90895 1 17322
2 90896 1 17322
2 90897 1 17331
2 90898 1 17331
2 90899 1 17331
2 90900 1 17331
2 90901 1 17331
2 90902 1 17331
2 90903 1 17332
2 90904 1 17332
2 90905 1 17340
2 90906 1 17340
2 90907 1 17353
2 90908 1 17353
2 90909 1 17353
2 90910 1 17354
2 90911 1 17354
2 90912 1 17354
2 90913 1 17378
2 90914 1 17378
2 90915 1 17393
2 90916 1 17393
2 90917 1 17404
2 90918 1 17404
2 90919 1 17407
2 90920 1 17407
2 90921 1 17420
2 90922 1 17420
2 90923 1 17421
2 90924 1 17421
2 90925 1 17421
2 90926 1 17421
2 90927 1 17421
2 90928 1 17421
2 90929 1 17421
2 90930 1 17421
2 90931 1 17450
2 90932 1 17450
2 90933 1 17454
2 90934 1 17454
2 90935 1 17454
2 90936 1 17463
2 90937 1 17463
2 90938 1 17463
2 90939 1 17463
2 90940 1 17463
2 90941 1 17464
2 90942 1 17464
2 90943 1 17477
2 90944 1 17477
2 90945 1 17481
2 90946 1 17481
2 90947 1 17485
2 90948 1 17485
2 90949 1 17486
2 90950 1 17486
2 90951 1 17486
2 90952 1 17486
2 90953 1 17487
2 90954 1 17487
2 90955 1 17487
2 90956 1 17488
2 90957 1 17488
2 90958 1 17489
2 90959 1 17489
2 90960 1 17489
2 90961 1 17494
2 90962 1 17494
2 90963 1 17494
2 90964 1 17494
2 90965 1 17495
2 90966 1 17495
2 90967 1 17495
2 90968 1 17497
2 90969 1 17497
2 90970 1 17497
2 90971 1 17497
2 90972 1 17503
2 90973 1 17503
2 90974 1 17503
2 90975 1 17509
2 90976 1 17509
2 90977 1 17509
2 90978 1 17509
2 90979 1 17509
2 90980 1 17509
2 90981 1 17509
2 90982 1 17510
2 90983 1 17510
2 90984 1 17510
2 90985 1 17510
2 90986 1 17514
2 90987 1 17514
2 90988 1 17564
2 90989 1 17564
2 90990 1 17604
2 90991 1 17604
2 90992 1 17604
2 90993 1 17611
2 90994 1 17611
2 90995 1 17611
2 90996 1 17616
2 90997 1 17616
2 90998 1 17642
2 90999 1 17642
2 91000 1 17642
2 91001 1 17642
2 91002 1 17644
2 91003 1 17644
2 91004 1 17644
2 91005 1 17645
2 91006 1 17645
2 91007 1 17645
2 91008 1 17669
2 91009 1 17669
2 91010 1 17669
2 91011 1 17669
2 91012 1 17669
2 91013 1 17669
2 91014 1 17669
2 91015 1 17669
2 91016 1 17678
2 91017 1 17678
2 91018 1 17689
2 91019 1 17689
2 91020 1 17689
2 91021 1 17738
2 91022 1 17738
2 91023 1 17746
2 91024 1 17746
2 91025 1 17748
2 91026 1 17748
2 91027 1 17748
2 91028 1 17785
2 91029 1 17785
2 91030 1 17785
2 91031 1 17788
2 91032 1 17788
2 91033 1 17792
2 91034 1 17792
2 91035 1 17793
2 91036 1 17793
2 91037 1 17811
2 91038 1 17811
2 91039 1 17811
2 91040 1 17819
2 91041 1 17819
2 91042 1 17819
2 91043 1 17833
2 91044 1 17833
2 91045 1 17834
2 91046 1 17834
2 91047 1 17834
2 91048 1 17835
2 91049 1 17835
2 91050 1 17861
2 91051 1 17861
2 91052 1 17861
2 91053 1 17861
2 91054 1 17861
2 91055 1 17861
2 91056 1 17865
2 91057 1 17865
2 91058 1 17865
2 91059 1 17872
2 91060 1 17872
2 91061 1 17880
2 91062 1 17880
2 91063 1 17880
2 91064 1 17880
2 91065 1 17896
2 91066 1 17896
2 91067 1 17909
2 91068 1 17909
2 91069 1 17909
2 91070 1 17909
2 91071 1 17909
2 91072 1 17909
2 91073 1 17909
2 91074 1 17909
2 91075 1 17909
2 91076 1 17910
2 91077 1 17910
2 91078 1 17912
2 91079 1 17912
2 91080 1 17912
2 91081 1 17931
2 91082 1 17931
2 91083 1 17931
2 91084 1 17932
2 91085 1 17932
2 91086 1 17935
2 91087 1 17935
2 91088 1 17935
2 91089 1 17935
2 91090 1 17957
2 91091 1 17957
2 91092 1 17957
2 91093 1 17957
2 91094 1 17984
2 91095 1 17984
2 91096 1 17997
2 91097 1 17997
2 91098 1 18005
2 91099 1 18005
2 91100 1 18005
2 91101 1 18005
2 91102 1 18005
2 91103 1 18005
2 91104 1 18014
2 91105 1 18014
2 91106 1 18032
2 91107 1 18032
2 91108 1 18033
2 91109 1 18033
2 91110 1 18033
2 91111 1 18033
2 91112 1 18033
2 91113 1 18034
2 91114 1 18034
2 91115 1 18034
2 91116 1 18035
2 91117 1 18035
2 91118 1 18049
2 91119 1 18049
2 91120 1 18061
2 91121 1 18061
2 91122 1 18061
2 91123 1 18061
2 91124 1 18061
2 91125 1 18061
2 91126 1 18061
2 91127 1 18061
2 91128 1 18061
2 91129 1 18061
2 91130 1 18061
2 91131 1 18062
2 91132 1 18062
2 91133 1 18062
2 91134 1 18062
2 91135 1 18062
2 91136 1 18062
2 91137 1 18063
2 91138 1 18063
2 91139 1 18063
2 91140 1 18081
2 91141 1 18081
2 91142 1 18090
2 91143 1 18090
2 91144 1 18090
2 91145 1 18090
2 91146 1 18092
2 91147 1 18092
2 91148 1 18095
2 91149 1 18095
2 91150 1 18095
2 91151 1 18095
2 91152 1 18105
2 91153 1 18105
2 91154 1 18105
2 91155 1 18120
2 91156 1 18120
2 91157 1 18120
2 91158 1 18120
2 91159 1 18120
2 91160 1 18120
2 91161 1 18120
2 91162 1 18120
2 91163 1 18120
2 91164 1 18120
2 91165 1 18120
2 91166 1 18121
2 91167 1 18121
2 91168 1 18129
2 91169 1 18129
2 91170 1 18129
2 91171 1 18130
2 91172 1 18130
2 91173 1 18130
2 91174 1 18130
2 91175 1 18148
2 91176 1 18148
2 91177 1 18148
2 91178 1 18148
2 91179 1 18148
2 91180 1 18155
2 91181 1 18155
2 91182 1 18155
2 91183 1 18155
2 91184 1 18155
2 91185 1 18164
2 91186 1 18164
2 91187 1 18165
2 91188 1 18165
2 91189 1 18166
2 91190 1 18166
2 91191 1 18178
2 91192 1 18178
2 91193 1 18178
2 91194 1 18178
2 91195 1 18178
2 91196 1 18178
2 91197 1 18191
2 91198 1 18191
2 91199 1 18191
2 91200 1 18192
2 91201 1 18192
2 91202 1 18192
2 91203 1 18194
2 91204 1 18194
2 91205 1 18196
2 91206 1 18196
2 91207 1 18196
2 91208 1 18196
2 91209 1 18212
2 91210 1 18212
2 91211 1 18212
2 91212 1 18212
2 91213 1 18212
2 91214 1 18212
2 91215 1 18212
2 91216 1 18213
2 91217 1 18213
2 91218 1 18213
2 91219 1 18259
2 91220 1 18259
2 91221 1 18259
2 91222 1 18260
2 91223 1 18260
2 91224 1 18261
2 91225 1 18261
2 91226 1 18279
2 91227 1 18279
2 91228 1 18279
2 91229 1 18279
2 91230 1 18289
2 91231 1 18289
2 91232 1 18289
2 91233 1 18292
2 91234 1 18292
2 91235 1 18293
2 91236 1 18293
2 91237 1 18315
2 91238 1 18315
2 91239 1 18315
2 91240 1 18316
2 91241 1 18316
2 91242 1 18316
2 91243 1 18319
2 91244 1 18319
2 91245 1 18319
2 91246 1 18319
2 91247 1 18338
2 91248 1 18338
2 91249 1 18344
2 91250 1 18344
2 91251 1 18344
2 91252 1 18345
2 91253 1 18345
2 91254 1 18368
2 91255 1 18368
2 91256 1 18369
2 91257 1 18369
2 91258 1 18435
2 91259 1 18435
2 91260 1 18435
2 91261 1 18435
2 91262 1 18436
2 91263 1 18436
2 91264 1 18457
2 91265 1 18457
2 91266 1 18459
2 91267 1 18459
2 91268 1 18465
2 91269 1 18465
2 91270 1 18477
2 91271 1 18477
2 91272 1 18477
2 91273 1 18478
2 91274 1 18478
2 91275 1 18503
2 91276 1 18503
2 91277 1 18504
2 91278 1 18504
2 91279 1 18523
2 91280 1 18523
2 91281 1 18523
2 91282 1 18524
2 91283 1 18524
2 91284 1 18525
2 91285 1 18525
2 91286 1 18532
2 91287 1 18532
2 91288 1 18532
2 91289 1 18532
2 91290 1 18533
2 91291 1 18533
2 91292 1 18556
2 91293 1 18556
2 91294 1 18556
2 91295 1 18567
2 91296 1 18567
2 91297 1 18567
2 91298 1 18567
2 91299 1 18568
2 91300 1 18568
2 91301 1 18568
2 91302 1 18571
2 91303 1 18571
2 91304 1 18572
2 91305 1 18572
2 91306 1 18572
2 91307 1 18572
2 91308 1 18577
2 91309 1 18577
2 91310 1 18577
2 91311 1 18577
2 91312 1 18577
2 91313 1 18591
2 91314 1 18591
2 91315 1 18592
2 91316 1 18592
2 91317 1 18611
2 91318 1 18611
2 91319 1 18611
2 91320 1 18623
2 91321 1 18623
2 91322 1 18623
2 91323 1 18623
2 91324 1 18623
2 91325 1 18623
2 91326 1 18623
2 91327 1 18624
2 91328 1 18624
2 91329 1 18625
2 91330 1 18625
2 91331 1 18625
2 91332 1 18631
2 91333 1 18631
2 91334 1 18631
2 91335 1 18632
2 91336 1 18632
2 91337 1 18658
2 91338 1 18658
2 91339 1 18691
2 91340 1 18691
2 91341 1 18691
2 91342 1 18691
2 91343 1 18722
2 91344 1 18722
2 91345 1 18722
2 91346 1 18722
2 91347 1 18722
2 91348 1 18722
2 91349 1 18724
2 91350 1 18724
2 91351 1 18737
2 91352 1 18737
2 91353 1 18741
2 91354 1 18741
2 91355 1 18753
2 91356 1 18753
2 91357 1 18753
2 91358 1 18757
2 91359 1 18757
2 91360 1 18757
2 91361 1 18757
2 91362 1 18757
2 91363 1 18757
2 91364 1 18757
2 91365 1 18757
2 91366 1 18757
2 91367 1 18757
2 91368 1 18757
2 91369 1 18767
2 91370 1 18767
2 91371 1 18770
2 91372 1 18770
2 91373 1 18773
2 91374 1 18773
2 91375 1 18773
2 91376 1 18773
2 91377 1 18773
2 91378 1 18774
2 91379 1 18774
2 91380 1 18777
2 91381 1 18777
2 91382 1 18793
2 91383 1 18793
2 91384 1 18793
2 91385 1 18793
2 91386 1 18794
2 91387 1 18794
2 91388 1 18794
2 91389 1 18795
2 91390 1 18795
2 91391 1 18811
2 91392 1 18811
2 91393 1 18812
2 91394 1 18812
2 91395 1 18812
2 91396 1 18812
2 91397 1 18824
2 91398 1 18824
2 91399 1 18825
2 91400 1 18825
2 91401 1 18825
2 91402 1 18845
2 91403 1 18845
2 91404 1 18845
2 91405 1 18845
2 91406 1 18846
2 91407 1 18846
2 91408 1 18846
2 91409 1 18848
2 91410 1 18848
2 91411 1 18848
2 91412 1 18848
2 91413 1 18848
2 91414 1 18848
2 91415 1 18849
2 91416 1 18849
2 91417 1 18851
2 91418 1 18851
2 91419 1 18851
2 91420 1 18851
2 91421 1 18873
2 91422 1 18873
2 91423 1 18873
2 91424 1 18873
2 91425 1 18873
2 91426 1 18875
2 91427 1 18875
2 91428 1 18876
2 91429 1 18876
2 91430 1 18876
2 91431 1 18876
2 91432 1 18876
2 91433 1 18876
2 91434 1 18885
2 91435 1 18885
2 91436 1 18889
2 91437 1 18889
2 91438 1 18889
2 91439 1 18904
2 91440 1 18904
2 91441 1 18904
2 91442 1 18904
2 91443 1 18904
2 91444 1 18904
2 91445 1 18908
2 91446 1 18908
2 91447 1 18928
2 91448 1 18928
2 91449 1 18928
2 91450 1 18930
2 91451 1 18930
2 91452 1 18956
2 91453 1 18956
2 91454 1 18957
2 91455 1 18957
2 91456 1 18957
2 91457 1 18957
2 91458 1 18960
2 91459 1 18960
2 91460 1 18965
2 91461 1 18965
2 91462 1 18965
2 91463 1 18965
2 91464 1 18968
2 91465 1 18968
2 91466 1 18977
2 91467 1 18977
2 91468 1 18977
2 91469 1 18996
2 91470 1 18996
2 91471 1 18996
2 91472 1 18996
2 91473 1 19022
2 91474 1 19022
2 91475 1 19022
2 91476 1 19022
2 91477 1 19037
2 91478 1 19037
2 91479 1 19044
2 91480 1 19044
2 91481 1 19045
2 91482 1 19045
2 91483 1 19045
2 91484 1 19045
2 91485 1 19047
2 91486 1 19047
2 91487 1 19047
2 91488 1 19051
2 91489 1 19051
2 91490 1 19058
2 91491 1 19058
2 91492 1 19060
2 91493 1 19060
2 91494 1 19061
2 91495 1 19061
2 91496 1 19106
2 91497 1 19106
2 91498 1 19106
2 91499 1 19115
2 91500 1 19115
2 91501 1 19115
2 91502 1 19130
2 91503 1 19130
2 91504 1 19130
2 91505 1 19137
2 91506 1 19137
2 91507 1 19137
2 91508 1 19137
2 91509 1 19137
2 91510 1 19179
2 91511 1 19179
2 91512 1 19179
2 91513 1 19179
2 91514 1 19194
2 91515 1 19194
2 91516 1 19194
2 91517 1 19194
2 91518 1 19196
2 91519 1 19196
2 91520 1 19212
2 91521 1 19212
2 91522 1 19237
2 91523 1 19237
2 91524 1 19245
2 91525 1 19245
2 91526 1 19245
2 91527 1 19245
2 91528 1 19245
2 91529 1 19245
2 91530 1 19245
2 91531 1 19245
2 91532 1 19245
2 91533 1 19246
2 91534 1 19246
2 91535 1 19246
2 91536 1 19246
2 91537 1 19246
2 91538 1 19246
2 91539 1 19246
2 91540 1 19246
2 91541 1 19247
2 91542 1 19247
2 91543 1 19247
2 91544 1 19247
2 91545 1 19247
2 91546 1 19247
2 91547 1 19250
2 91548 1 19250
2 91549 1 19252
2 91550 1 19252
2 91551 1 19253
2 91552 1 19253
2 91553 1 19253
2 91554 1 19254
2 91555 1 19254
2 91556 1 19254
2 91557 1 19254
2 91558 1 19254
2 91559 1 19255
2 91560 1 19255
2 91561 1 19270
2 91562 1 19270
2 91563 1 19278
2 91564 1 19278
2 91565 1 19278
2 91566 1 19279
2 91567 1 19279
2 91568 1 19316
2 91569 1 19316
2 91570 1 19328
2 91571 1 19328
2 91572 1 19328
2 91573 1 19328
2 91574 1 19329
2 91575 1 19329
2 91576 1 19329
2 91577 1 19340
2 91578 1 19340
2 91579 1 19340
2 91580 1 19340
2 91581 1 19340
2 91582 1 19344
2 91583 1 19344
2 91584 1 19354
2 91585 1 19354
2 91586 1 19364
2 91587 1 19364
2 91588 1 19365
2 91589 1 19365
2 91590 1 19366
2 91591 1 19366
2 91592 1 19366
2 91593 1 19366
2 91594 1 19366
2 91595 1 19366
2 91596 1 19366
2 91597 1 19366
2 91598 1 19366
2 91599 1 19367
2 91600 1 19367
2 91601 1 19367
2 91602 1 19370
2 91603 1 19370
2 91604 1 19370
2 91605 1 19397
2 91606 1 19397
2 91607 1 19397
2 91608 1 19410
2 91609 1 19410
2 91610 1 19412
2 91611 1 19412
2 91612 1 19421
2 91613 1 19421
2 91614 1 19424
2 91615 1 19424
2 91616 1 19431
2 91617 1 19431
2 91618 1 19431
2 91619 1 19461
2 91620 1 19461
2 91621 1 19477
2 91622 1 19477
2 91623 1 19498
2 91624 1 19498
2 91625 1 19498
2 91626 1 19498
2 91627 1 19498
2 91628 1 19499
2 91629 1 19499
2 91630 1 19500
2 91631 1 19500
2 91632 1 19524
2 91633 1 19524
2 91634 1 19542
2 91635 1 19542
2 91636 1 19543
2 91637 1 19543
2 91638 1 19570
2 91639 1 19570
2 91640 1 19588
2 91641 1 19588
2 91642 1 19588
2 91643 1 19589
2 91644 1 19589
2 91645 1 19590
2 91646 1 19590
2 91647 1 19601
2 91648 1 19601
2 91649 1 19601
2 91650 1 19601
2 91651 1 19602
2 91652 1 19602
2 91653 1 19620
2 91654 1 19620
2 91655 1 19620
2 91656 1 19620
2 91657 1 19620
2 91658 1 19620
2 91659 1 19620
2 91660 1 19620
2 91661 1 19620
2 91662 1 19620
2 91663 1 19620
2 91664 1 19621
2 91665 1 19621
2 91666 1 19621
2 91667 1 19621
2 91668 1 19621
2 91669 1 19621
2 91670 1 19621
2 91671 1 19621
2 91672 1 19621
2 91673 1 19621
2 91674 1 19621
2 91675 1 19621
2 91676 1 19621
2 91677 1 19621
2 91678 1 19621
2 91679 1 19621
2 91680 1 19621
2 91681 1 19621
2 91682 1 19621
2 91683 1 19621
2 91684 1 19621
2 91685 1 19621
2 91686 1 19621
2 91687 1 19621
2 91688 1 19621
2 91689 1 19621
2 91690 1 19621
2 91691 1 19621
2 91692 1 19621
2 91693 1 19621
2 91694 1 19621
2 91695 1 19621
2 91696 1 19621
2 91697 1 19621
2 91698 1 19621
2 91699 1 19621
2 91700 1 19621
2 91701 1 19621
2 91702 1 19621
2 91703 1 19621
2 91704 1 19621
2 91705 1 19621
2 91706 1 19621
2 91707 1 19621
2 91708 1 19621
2 91709 1 19621
2 91710 1 19621
2 91711 1 19621
2 91712 1 19621
2 91713 1 19621
2 91714 1 19621
2 91715 1 19621
2 91716 1 19621
2 91717 1 19621
2 91718 1 19621
2 91719 1 19621
2 91720 1 19621
2 91721 1 19621
2 91722 1 19621
2 91723 1 19621
2 91724 1 19621
2 91725 1 19621
2 91726 1 19621
2 91727 1 19621
2 91728 1 19621
2 91729 1 19621
2 91730 1 19621
2 91731 1 19621
2 91732 1 19621
2 91733 1 19621
2 91734 1 19621
2 91735 1 19621
2 91736 1 19621
2 91737 1 19621
2 91738 1 19621
2 91739 1 19622
2 91740 1 19622
2 91741 1 19622
2 91742 1 19622
2 91743 1 19628
2 91744 1 19628
2 91745 1 19642
2 91746 1 19642
2 91747 1 19650
2 91748 1 19650
2 91749 1 19650
2 91750 1 19650
2 91751 1 19655
2 91752 1 19655
2 91753 1 19672
2 91754 1 19672
2 91755 1 19672
2 91756 1 19672
2 91757 1 19672
2 91758 1 19672
2 91759 1 19672
2 91760 1 19672
2 91761 1 19672
2 91762 1 19672
2 91763 1 19672
2 91764 1 19672
2 91765 1 19672
2 91766 1 19673
2 91767 1 19673
2 91768 1 19674
2 91769 1 19674
2 91770 1 19675
2 91771 1 19675
2 91772 1 19675
2 91773 1 19685
2 91774 1 19685
2 91775 1 19685
2 91776 1 19685
2 91777 1 19685
2 91778 1 19686
2 91779 1 19686
2 91780 1 19695
2 91781 1 19695
2 91782 1 19695
2 91783 1 19706
2 91784 1 19706
2 91785 1 19706
2 91786 1 19717
2 91787 1 19717
2 91788 1 19718
2 91789 1 19718
2 91790 1 19727
2 91791 1 19727
2 91792 1 19728
2 91793 1 19728
2 91794 1 19730
2 91795 1 19730
2 91796 1 19730
2 91797 1 19730
2 91798 1 19739
2 91799 1 19739
2 91800 1 19747
2 91801 1 19747
2 91802 1 19750
2 91803 1 19750
2 91804 1 19752
2 91805 1 19752
2 91806 1 19783
2 91807 1 19783
2 91808 1 19783
2 91809 1 19783
2 91810 1 19783
2 91811 1 19783
2 91812 1 19783
2 91813 1 19783
2 91814 1 19783
2 91815 1 19783
2 91816 1 19783
2 91817 1 19783
2 91818 1 19795
2 91819 1 19795
2 91820 1 19795
2 91821 1 19795
2 91822 1 19795
2 91823 1 19795
2 91824 1 19795
2 91825 1 19795
2 91826 1 19795
2 91827 1 19795
2 91828 1 19795
2 91829 1 19795
2 91830 1 19795
2 91831 1 19795
2 91832 1 19795
2 91833 1 19795
2 91834 1 19795
2 91835 1 19796
2 91836 1 19796
2 91837 1 19796
2 91838 1 19798
2 91839 1 19798
2 91840 1 19815
2 91841 1 19815
2 91842 1 19817
2 91843 1 19817
2 91844 1 19817
2 91845 1 19817
2 91846 1 19817
2 91847 1 19817
2 91848 1 19817
2 91849 1 19817
2 91850 1 19817
2 91851 1 19817
2 91852 1 19818
2 91853 1 19818
2 91854 1 19818
2 91855 1 19818
2 91856 1 19818
2 91857 1 19818
2 91858 1 19818
2 91859 1 19818
2 91860 1 19818
2 91861 1 19818
2 91862 1 19818
2 91863 1 19818
2 91864 1 19818
2 91865 1 19818
2 91866 1 19818
2 91867 1 19818
2 91868 1 19818
2 91869 1 19818
2 91870 1 19818
2 91871 1 19818
2 91872 1 19818
2 91873 1 19818
2 91874 1 19818
2 91875 1 19818
2 91876 1 19818
2 91877 1 19818
2 91878 1 19818
2 91879 1 19818
2 91880 1 19818
2 91881 1 19818
2 91882 1 19818
2 91883 1 19818
2 91884 1 19829
2 91885 1 19829
2 91886 1 19829
2 91887 1 19829
2 91888 1 19829
2 91889 1 19829
2 91890 1 19829
2 91891 1 19830
2 91892 1 19830
2 91893 1 19830
2 91894 1 19830
2 91895 1 19830
2 91896 1 19830
2 91897 1 19830
2 91898 1 19832
2 91899 1 19832
2 91900 1 19874
2 91901 1 19874
2 91902 1 19874
2 91903 1 19875
2 91904 1 19875
2 91905 1 19875
2 91906 1 19896
2 91907 1 19896
2 91908 1 19896
2 91909 1 19905
2 91910 1 19905
2 91911 1 19905
2 91912 1 19914
2 91913 1 19914
2 91914 1 19932
2 91915 1 19932
2 91916 1 19934
2 91917 1 19934
2 91918 1 19934
2 91919 1 19934
2 91920 1 19934
2 91921 1 19952
2 91922 1 19952
2 91923 1 19952
2 91924 1 19967
2 91925 1 19967
2 91926 1 19977
2 91927 1 19977
2 91928 1 19977
2 91929 1 19977
2 91930 1 19988
2 91931 1 19988
2 91932 1 19996
2 91933 1 19996
2 91934 1 19997
2 91935 1 19997
2 91936 1 20021
2 91937 1 20021
2 91938 1 20022
2 91939 1 20022
2 91940 1 20023
2 91941 1 20023
2 91942 1 20031
2 91943 1 20031
2 91944 1 20031
2 91945 1 20031
2 91946 1 20031
2 91947 1 20031
2 91948 1 20037
2 91949 1 20037
2 91950 1 20037
2 91951 1 20037
2 91952 1 20046
2 91953 1 20046
2 91954 1 20071
2 91955 1 20071
2 91956 1 20071
2 91957 1 20072
2 91958 1 20072
2 91959 1 20077
2 91960 1 20077
2 91961 1 20077
2 91962 1 20080
2 91963 1 20080
2 91964 1 20109
2 91965 1 20109
2 91966 1 20127
2 91967 1 20127
2 91968 1 20151
2 91969 1 20151
2 91970 1 20153
2 91971 1 20153
2 91972 1 20189
2 91973 1 20189
2 91974 1 20202
2 91975 1 20202
2 91976 1 20202
2 91977 1 20203
2 91978 1 20203
2 91979 1 20211
2 91980 1 20211
2 91981 1 20219
2 91982 1 20219
2 91983 1 20219
2 91984 1 20219
2 91985 1 20219
2 91986 1 20222
2 91987 1 20222
2 91988 1 20222
2 91989 1 20222
2 91990 1 20223
2 91991 1 20223
2 91992 1 20239
2 91993 1 20239
2 91994 1 20239
2 91995 1 20239
2 91996 1 20239
2 91997 1 20239
2 91998 1 20239
2 91999 1 20239
2 92000 1 20239
2 92001 1 20240
2 92002 1 20240
2 92003 1 20247
2 92004 1 20247
2 92005 1 20247
2 92006 1 20247
2 92007 1 20247
2 92008 1 20247
2 92009 1 20247
2 92010 1 20256
2 92011 1 20256
2 92012 1 20256
2 92013 1 20256
2 92014 1 20256
2 92015 1 20256
2 92016 1 20265
2 92017 1 20265
2 92018 1 20278
2 92019 1 20278
2 92020 1 20278
2 92021 1 20278
2 92022 1 20278
2 92023 1 20282
2 92024 1 20282
2 92025 1 20282
2 92026 1 20282
2 92027 1 20282
2 92028 1 20282
2 92029 1 20282
2 92030 1 20290
2 92031 1 20290
2 92032 1 20290
2 92033 1 20290
2 92034 1 20291
2 92035 1 20291
2 92036 1 20291
2 92037 1 20291
2 92038 1 20291
2 92039 1 20292
2 92040 1 20292
2 92041 1 20300
2 92042 1 20300
2 92043 1 20300
2 92044 1 20300
2 92045 1 20300
2 92046 1 20300
2 92047 1 20302
2 92048 1 20302
2 92049 1 20302
2 92050 1 20303
2 92051 1 20303
2 92052 1 20306
2 92053 1 20306
2 92054 1 20306
2 92055 1 20306
2 92056 1 20306
2 92057 1 20307
2 92058 1 20307
2 92059 1 20326
2 92060 1 20326
2 92061 1 20326
2 92062 1 20326
2 92063 1 20326
2 92064 1 20336
2 92065 1 20336
2 92066 1 20337
2 92067 1 20337
2 92068 1 20346
2 92069 1 20346
2 92070 1 20358
2 92071 1 20358
2 92072 1 20370
2 92073 1 20370
2 92074 1 20371
2 92075 1 20371
2 92076 1 20379
2 92077 1 20379
2 92078 1 20380
2 92079 1 20380
2 92080 1 20380
2 92081 1 20380
2 92082 1 20380
2 92083 1 20385
2 92084 1 20385
2 92085 1 20396
2 92086 1 20396
2 92087 1 20399
2 92088 1 20399
2 92089 1 20399
2 92090 1 20401
2 92091 1 20401
2 92092 1 20413
2 92093 1 20413
2 92094 1 20413
2 92095 1 20413
2 92096 1 20413
2 92097 1 20413
2 92098 1 20413
2 92099 1 20431
2 92100 1 20431
2 92101 1 20437
2 92102 1 20437
2 92103 1 20437
2 92104 1 20437
2 92105 1 20437
2 92106 1 20439
2 92107 1 20439
2 92108 1 20455
2 92109 1 20455
2 92110 1 20455
2 92111 1 20456
2 92112 1 20456
2 92113 1 20457
2 92114 1 20457
2 92115 1 20472
2 92116 1 20472
2 92117 1 20472
2 92118 1 20472
2 92119 1 20472
2 92120 1 20472
2 92121 1 20472
2 92122 1 20472
2 92123 1 20472
2 92124 1 20472
2 92125 1 20472
2 92126 1 20472
2 92127 1 20472
2 92128 1 20472
2 92129 1 20472
2 92130 1 20473
2 92131 1 20473
2 92132 1 20473
2 92133 1 20492
2 92134 1 20492
2 92135 1 20492
2 92136 1 20497
2 92137 1 20497
2 92138 1 20497
2 92139 1 20497
2 92140 1 20508
2 92141 1 20508
2 92142 1 20508
2 92143 1 20508
2 92144 1 20518
2 92145 1 20518
2 92146 1 20518
2 92147 1 20521
2 92148 1 20521
2 92149 1 20521
2 92150 1 20521
2 92151 1 20521
2 92152 1 20521
2 92153 1 20525
2 92154 1 20525
2 92155 1 20525
2 92156 1 20525
2 92157 1 20525
2 92158 1 20546
2 92159 1 20546
2 92160 1 20546
2 92161 1 20546
2 92162 1 20546
2 92163 1 20546
2 92164 1 20548
2 92165 1 20548
2 92166 1 20553
2 92167 1 20553
2 92168 1 20553
2 92169 1 20553
2 92170 1 20561
2 92171 1 20561
2 92172 1 20562
2 92173 1 20562
2 92174 1 20562
2 92175 1 20562
2 92176 1 20562
2 92177 1 20562
2 92178 1 20562
2 92179 1 20563
2 92180 1 20563
2 92181 1 20580
2 92182 1 20580
2 92183 1 20580
2 92184 1 20580
2 92185 1 20585
2 92186 1 20585
2 92187 1 20585
2 92188 1 20616
2 92189 1 20616
2 92190 1 20620
2 92191 1 20620
2 92192 1 20621
2 92193 1 20621
2 92194 1 20621
2 92195 1 20621
2 92196 1 20622
2 92197 1 20622
2 92198 1 20640
2 92199 1 20640
2 92200 1 20642
2 92201 1 20642
2 92202 1 20652
2 92203 1 20652
2 92204 1 20652
2 92205 1 20656
2 92206 1 20656
2 92207 1 20664
2 92208 1 20664
2 92209 1 20665
2 92210 1 20665
2 92211 1 20666
2 92212 1 20666
2 92213 1 20666
2 92214 1 20666
2 92215 1 20666
2 92216 1 20674
2 92217 1 20674
2 92218 1 20690
2 92219 1 20690
2 92220 1 20691
2 92221 1 20691
2 92222 1 20694
2 92223 1 20694
2 92224 1 20708
2 92225 1 20708
2 92226 1 20708
2 92227 1 20708
2 92228 1 20708
2 92229 1 20708
2 92230 1 20719
2 92231 1 20719
2 92232 1 20719
2 92233 1 20719
2 92234 1 20719
2 92235 1 20728
2 92236 1 20728
2 92237 1 20739
2 92238 1 20739
2 92239 1 20780
2 92240 1 20780
2 92241 1 20780
2 92242 1 20781
2 92243 1 20781
2 92244 1 20781
2 92245 1 20783
2 92246 1 20783
2 92247 1 20783
2 92248 1 20795
2 92249 1 20795
2 92250 1 20798
2 92251 1 20798
2 92252 1 20800
2 92253 1 20800
2 92254 1 20810
2 92255 1 20810
2 92256 1 20810
2 92257 1 20810
2 92258 1 20836
2 92259 1 20836
2 92260 1 20850
2 92261 1 20850
2 92262 1 20872
2 92263 1 20872
2 92264 1 20874
2 92265 1 20874
2 92266 1 20874
2 92267 1 20874
2 92268 1 20874
2 92269 1 20874
2 92270 1 20874
2 92271 1 20874
2 92272 1 20874
2 92273 1 20874
2 92274 1 20874
2 92275 1 20875
2 92276 1 20875
2 92277 1 20875
2 92278 1 20883
2 92279 1 20883
2 92280 1 20883
2 92281 1 20883
2 92282 1 20883
2 92283 1 20883
2 92284 1 20883
2 92285 1 20883
2 92286 1 20883
2 92287 1 20883
2 92288 1 20884
2 92289 1 20884
2 92290 1 20885
2 92291 1 20885
2 92292 1 20886
2 92293 1 20886
2 92294 1 20886
2 92295 1 20887
2 92296 1 20887
2 92297 1 20891
2 92298 1 20891
2 92299 1 20891
2 92300 1 20896
2 92301 1 20896
2 92302 1 20896
2 92303 1 20896
2 92304 1 20897
2 92305 1 20897
2 92306 1 20900
2 92307 1 20900
2 92308 1 20900
2 92309 1 20900
2 92310 1 20900
2 92311 1 20900
2 92312 1 20900
2 92313 1 20900
2 92314 1 20900
2 92315 1 20900
2 92316 1 20900
2 92317 1 20900
2 92318 1 20900
2 92319 1 20902
2 92320 1 20902
2 92321 1 20902
2 92322 1 20902
2 92323 1 20903
2 92324 1 20903
2 92325 1 20905
2 92326 1 20905
2 92327 1 20905
2 92328 1 20905
2 92329 1 20905
2 92330 1 20907
2 92331 1 20907
2 92332 1 20907
2 92333 1 20907
2 92334 1 20907
2 92335 1 20907
2 92336 1 20907
2 92337 1 20908
2 92338 1 20908
2 92339 1 20909
2 92340 1 20909
2 92341 1 20909
2 92342 1 20922
2 92343 1 20922
2 92344 1 20923
2 92345 1 20923
2 92346 1 20923
2 92347 1 20923
2 92348 1 20924
2 92349 1 20924
2 92350 1 20924
2 92351 1 20924
2 92352 1 20924
2 92353 1 20932
2 92354 1 20932
2 92355 1 20932
2 92356 1 20932
2 92357 1 20932
2 92358 1 20932
2 92359 1 20934
2 92360 1 20934
2 92361 1 20934
2 92362 1 20934
2 92363 1 20949
2 92364 1 20949
2 92365 1 20950
2 92366 1 20950
2 92367 1 20951
2 92368 1 20951
2 92369 1 20966
2 92370 1 20966
2 92371 1 20966
2 92372 1 20966
2 92373 1 20966
2 92374 1 20966
2 92375 1 20966
2 92376 1 20966
2 92377 1 20967
2 92378 1 20967
2 92379 1 20970
2 92380 1 20970
2 92381 1 20987
2 92382 1 20987
2 92383 1 20988
2 92384 1 20988
2 92385 1 21004
2 92386 1 21004
2 92387 1 21004
2 92388 1 21004
2 92389 1 21005
2 92390 1 21005
2 92391 1 21012
2 92392 1 21012
2 92393 1 21026
2 92394 1 21026
2 92395 1 21029
2 92396 1 21029
2 92397 1 21047
2 92398 1 21047
2 92399 1 21047
2 92400 1 21048
2 92401 1 21048
2 92402 1 21049
2 92403 1 21049
2 92404 1 21054
2 92405 1 21054
2 92406 1 21055
2 92407 1 21055
2 92408 1 21056
2 92409 1 21056
2 92410 1 21056
2 92411 1 21056
2 92412 1 21056
2 92413 1 21069
2 92414 1 21069
2 92415 1 21070
2 92416 1 21070
2 92417 1 21070
2 92418 1 21070
2 92419 1 21070
2 92420 1 21070
2 92421 1 21080
2 92422 1 21080
2 92423 1 21101
2 92424 1 21101
2 92425 1 21101
2 92426 1 21101
2 92427 1 21121
2 92428 1 21121
2 92429 1 21125
2 92430 1 21125
2 92431 1 21128
2 92432 1 21128
2 92433 1 21128
2 92434 1 21129
2 92435 1 21129
2 92436 1 21142
2 92437 1 21142
2 92438 1 21143
2 92439 1 21143
2 92440 1 21146
2 92441 1 21146
2 92442 1 21160
2 92443 1 21160
2 92444 1 21175
2 92445 1 21175
2 92446 1 21184
2 92447 1 21184
2 92448 1 21197
2 92449 1 21197
2 92450 1 21197
2 92451 1 21197
2 92452 1 21197
2 92453 1 21197
2 92454 1 21197
2 92455 1 21198
2 92456 1 21198
2 92457 1 21198
2 92458 1 21198
2 92459 1 21198
2 92460 1 21199
2 92461 1 21199
2 92462 1 21199
2 92463 1 21217
2 92464 1 21217
2 92465 1 21247
2 92466 1 21247
2 92467 1 21248
2 92468 1 21248
2 92469 1 21257
2 92470 1 21257
2 92471 1 21271
2 92472 1 21271
2 92473 1 21286
2 92474 1 21286
2 92475 1 21293
2 92476 1 21293
2 92477 1 21293
2 92478 1 21293
2 92479 1 21293
2 92480 1 21293
2 92481 1 21293
2 92482 1 21293
2 92483 1 21293
2 92484 1 21294
2 92485 1 21294
2 92486 1 21325
2 92487 1 21325
2 92488 1 21325
2 92489 1 21325
2 92490 1 21325
2 92491 1 21371
2 92492 1 21371
2 92493 1 21372
2 92494 1 21372
2 92495 1 21393
2 92496 1 21393
2 92497 1 21415
2 92498 1 21415
2 92499 1 21415
2 92500 1 21422
2 92501 1 21422
2 92502 1 21422
2 92503 1 21423
2 92504 1 21423
2 92505 1 21439
2 92506 1 21439
2 92507 1 21439
2 92508 1 21439
2 92509 1 21468
2 92510 1 21468
2 92511 1 21476
2 92512 1 21476
2 92513 1 21476
2 92514 1 21476
2 92515 1 21476
2 92516 1 21477
2 92517 1 21477
2 92518 1 21477
2 92519 1 21478
2 92520 1 21478
2 92521 1 21487
2 92522 1 21487
2 92523 1 21487
2 92524 1 21487
2 92525 1 21487
2 92526 1 21487
2 92527 1 21514
2 92528 1 21514
2 92529 1 21514
2 92530 1 21514
2 92531 1 21514
2 92532 1 21516
2 92533 1 21516
2 92534 1 21516
2 92535 1 21516
2 92536 1 21520
2 92537 1 21520
2 92538 1 21524
2 92539 1 21524
2 92540 1 21524
2 92541 1 21524
2 92542 1 21524
2 92543 1 21524
2 92544 1 21540
2 92545 1 21540
2 92546 1 21540
2 92547 1 21540
2 92548 1 21540
2 92549 1 21546
2 92550 1 21546
2 92551 1 21554
2 92552 1 21554
2 92553 1 21559
2 92554 1 21559
2 92555 1 21559
2 92556 1 21559
2 92557 1 21559
2 92558 1 21560
2 92559 1 21560
2 92560 1 21560
2 92561 1 21560
2 92562 1 21560
2 92563 1 21560
2 92564 1 21565
2 92565 1 21565
2 92566 1 21566
2 92567 1 21566
2 92568 1 21569
2 92569 1 21569
2 92570 1 21569
2 92571 1 21569
2 92572 1 21569
2 92573 1 21570
2 92574 1 21570
2 92575 1 21585
2 92576 1 21585
2 92577 1 21617
2 92578 1 21617
2 92579 1 21618
2 92580 1 21618
2 92581 1 21627
2 92582 1 21627
2 92583 1 21627
2 92584 1 21628
2 92585 1 21628
2 92586 1 21630
2 92587 1 21630
2 92588 1 21639
2 92589 1 21639
2 92590 1 21642
2 92591 1 21642
2 92592 1 21642
2 92593 1 21642
2 92594 1 21642
2 92595 1 21642
2 92596 1 21642
2 92597 1 21654
2 92598 1 21654
2 92599 1 21654
2 92600 1 21654
2 92601 1 21655
2 92602 1 21655
2 92603 1 21667
2 92604 1 21667
2 92605 1 21667
2 92606 1 21678
2 92607 1 21678
2 92608 1 21689
2 92609 1 21689
2 92610 1 21694
2 92611 1 21694
2 92612 1 21698
2 92613 1 21698
2 92614 1 21733
2 92615 1 21733
2 92616 1 21741
2 92617 1 21741
2 92618 1 21741
2 92619 1 21742
2 92620 1 21742
2 92621 1 21742
2 92622 1 21742
2 92623 1 21757
2 92624 1 21757
2 92625 1 21761
2 92626 1 21761
2 92627 1 21761
2 92628 1 21761
2 92629 1 21761
2 92630 1 21761
2 92631 1 21773
2 92632 1 21773
2 92633 1 21774
2 92634 1 21774
2 92635 1 21774
2 92636 1 21799
2 92637 1 21799
2 92638 1 21799
2 92639 1 21799
2 92640 1 21799
2 92641 1 21799
2 92642 1 21799
2 92643 1 21799
2 92644 1 21799
2 92645 1 21801
2 92646 1 21801
2 92647 1 21801
2 92648 1 21811
2 92649 1 21811
2 92650 1 21818
2 92651 1 21818
2 92652 1 21819
2 92653 1 21819
2 92654 1 21848
2 92655 1 21848
2 92656 1 21848
2 92657 1 21849
2 92658 1 21849
2 92659 1 21849
2 92660 1 21849
2 92661 1 21850
2 92662 1 21850
2 92663 1 21851
2 92664 1 21851
2 92665 1 21852
2 92666 1 21852
2 92667 1 21852
2 92668 1 21852
2 92669 1 21852
2 92670 1 21852
2 92671 1 21852
2 92672 1 21852
2 92673 1 21852
2 92674 1 21852
2 92675 1 21852
2 92676 1 21852
2 92677 1 21874
2 92678 1 21874
2 92679 1 21874
2 92680 1 21875
2 92681 1 21875
2 92682 1 21876
2 92683 1 21876
2 92684 1 21882
2 92685 1 21882
2 92686 1 21883
2 92687 1 21883
2 92688 1 21923
2 92689 1 21923
2 92690 1 21925
2 92691 1 21925
2 92692 1 21942
2 92693 1 21942
2 92694 1 21942
2 92695 1 21986
2 92696 1 21986
2 92697 1 21986
2 92698 1 21986
2 92699 1 22024
2 92700 1 22024
2 92701 1 22024
2 92702 1 22051
2 92703 1 22051
2 92704 1 22051
2 92705 1 22051
2 92706 1 22051
2 92707 1 22085
2 92708 1 22085
2 92709 1 22086
2 92710 1 22086
2 92711 1 22087
2 92712 1 22087
2 92713 1 22090
2 92714 1 22090
2 92715 1 22101
2 92716 1 22101
2 92717 1 22153
2 92718 1 22153
2 92719 1 22153
2 92720 1 22153
2 92721 1 22153
2 92722 1 22192
2 92723 1 22192
2 92724 1 22194
2 92725 1 22194
2 92726 1 22194
2 92727 1 22196
2 92728 1 22196
2 92729 1 22209
2 92730 1 22209
2 92731 1 22210
2 92732 1 22210
2 92733 1 22210
2 92734 1 22240
2 92735 1 22240
2 92736 1 22240
2 92737 1 22240
2 92738 1 22241
2 92739 1 22241
2 92740 1 22241
2 92741 1 22241
2 92742 1 22241
2 92743 1 22241
2 92744 1 22241
2 92745 1 22241
2 92746 1 22241
2 92747 1 22244
2 92748 1 22244
2 92749 1 22268
2 92750 1 22268
2 92751 1 22268
2 92752 1 22268
2 92753 1 22268
2 92754 1 22268
2 92755 1 22275
2 92756 1 22275
2 92757 1 22278
2 92758 1 22278
2 92759 1 22297
2 92760 1 22297
2 92761 1 22309
2 92762 1 22309
2 92763 1 22309
2 92764 1 22309
2 92765 1 22309
2 92766 1 22322
2 92767 1 22322
2 92768 1 22322
2 92769 1 22322
2 92770 1 22322
2 92771 1 22322
2 92772 1 22322
2 92773 1 22322
2 92774 1 22322
2 92775 1 22322
2 92776 1 22322
2 92777 1 22322
2 92778 1 22323
2 92779 1 22323
2 92780 1 22323
2 92781 1 22323
2 92782 1 22323
2 92783 1 22323
2 92784 1 22323
2 92785 1 22324
2 92786 1 22324
2 92787 1 22324
2 92788 1 22324
2 92789 1 22370
2 92790 1 22370
2 92791 1 22370
2 92792 1 22370
2 92793 1 22370
2 92794 1 22370
2 92795 1 22371
2 92796 1 22371
2 92797 1 22374
2 92798 1 22374
2 92799 1 22374
2 92800 1 22374
2 92801 1 22374
2 92802 1 22375
2 92803 1 22375
2 92804 1 22378
2 92805 1 22378
2 92806 1 22378
2 92807 1 22390
2 92808 1 22390
2 92809 1 22399
2 92810 1 22399
2 92811 1 22399
2 92812 1 22399
2 92813 1 22400
2 92814 1 22400
2 92815 1 22400
2 92816 1 22401
2 92817 1 22401
2 92818 1 22401
2 92819 1 22401
2 92820 1 22401
2 92821 1 22402
2 92822 1 22402
2 92823 1 22403
2 92824 1 22403
2 92825 1 22403
2 92826 1 22403
2 92827 1 22408
2 92828 1 22408
2 92829 1 22408
2 92830 1 22408
2 92831 1 22408
2 92832 1 22424
2 92833 1 22424
2 92834 1 22424
2 92835 1 22425
2 92836 1 22425
2 92837 1 22425
2 92838 1 22425
2 92839 1 22425
2 92840 1 22453
2 92841 1 22453
2 92842 1 22453
2 92843 1 22453
2 92844 1 22453
2 92845 1 22453
2 92846 1 22461
2 92847 1 22461
2 92848 1 22476
2 92849 1 22476
2 92850 1 22484
2 92851 1 22484
2 92852 1 22484
2 92853 1 22502
2 92854 1 22502
2 92855 1 22502
2 92856 1 22502
2 92857 1 22502
2 92858 1 22502
2 92859 1 22502
2 92860 1 22502
2 92861 1 22503
2 92862 1 22503
2 92863 1 22503
2 92864 1 22531
2 92865 1 22531
2 92866 1 22531
2 92867 1 22531
2 92868 1 22531
2 92869 1 22531
2 92870 1 22531
2 92871 1 22531
2 92872 1 22547
2 92873 1 22547
2 92874 1 22547
2 92875 1 22556
2 92876 1 22556
2 92877 1 22565
2 92878 1 22565
2 92879 1 22645
2 92880 1 22645
2 92881 1 22660
2 92882 1 22660
2 92883 1 22660
2 92884 1 22660
2 92885 1 22660
2 92886 1 22661
2 92887 1 22661
2 92888 1 22661
2 92889 1 22680
2 92890 1 22680
2 92891 1 22680
2 92892 1 22686
2 92893 1 22686
2 92894 1 22697
2 92895 1 22697
2 92896 1 22724
2 92897 1 22724
2 92898 1 22725
2 92899 1 22725
2 92900 1 22725
2 92901 1 22725
2 92902 1 22778
2 92903 1 22778
2 92904 1 22806
2 92905 1 22806
2 92906 1 22806
2 92907 1 22806
2 92908 1 22807
2 92909 1 22807
2 92910 1 22811
2 92911 1 22811
2 92912 1 22826
2 92913 1 22826
2 92914 1 22827
2 92915 1 22827
2 92916 1 22828
2 92917 1 22828
2 92918 1 22842
2 92919 1 22842
2 92920 1 22843
2 92921 1 22843
2 92922 1 22850
2 92923 1 22850
2 92924 1 22850
2 92925 1 22851
2 92926 1 22851
2 92927 1 22898
2 92928 1 22898
2 92929 1 22927
2 92930 1 22927
2 92931 1 22943
2 92932 1 22943
2 92933 1 23001
2 92934 1 23001
2 92935 1 23001
2 92936 1 23017
2 92937 1 23017
2 92938 1 23017
2 92939 1 23049
2 92940 1 23049
2 92941 1 23049
2 92942 1 23096
2 92943 1 23096
2 92944 1 23097
2 92945 1 23097
2 92946 1 23097
2 92947 1 23110
2 92948 1 23110
2 92949 1 23117
2 92950 1 23117
2 92951 1 23120
2 92952 1 23120
2 92953 1 23128
2 92954 1 23128
2 92955 1 23128
2 92956 1 23128
2 92957 1 23128
2 92958 1 23128
2 92959 1 23128
2 92960 1 23138
2 92961 1 23138
2 92962 1 23150
2 92963 1 23150
2 92964 1 23150
2 92965 1 23150
2 92966 1 23159
2 92967 1 23159
2 92968 1 23216
2 92969 1 23216
2 92970 1 23230
2 92971 1 23230
2 92972 1 23231
2 92973 1 23231
2 92974 1 23276
2 92975 1 23276
2 92976 1 23276
2 92977 1 23294
2 92978 1 23294
2 92979 1 23316
2 92980 1 23316
2 92981 1 23316
2 92982 1 23316
2 92983 1 23316
2 92984 1 23316
2 92985 1 23316
2 92986 1 23316
2 92987 1 23372
2 92988 1 23372
2 92989 1 23412
2 92990 1 23412
2 92991 1 23438
2 92992 1 23438
2 92993 1 23438
2 92994 1 23451
2 92995 1 23451
2 92996 1 23455
2 92997 1 23455
2 92998 1 23528
2 92999 1 23528
2 93000 1 23534
2 93001 1 23534
2 93002 1 23539
2 93003 1 23539
2 93004 1 23541
2 93005 1 23541
2 93006 1 23564
2 93007 1 23564
2 93008 1 23569
2 93009 1 23569
2 93010 1 23575
2 93011 1 23575
2 93012 1 23575
2 93013 1 23575
2 93014 1 23587
2 93015 1 23587
2 93016 1 23588
2 93017 1 23588
2 93018 1 23588
2 93019 1 23602
2 93020 1 23602
2 93021 1 23605
2 93022 1 23605
2 93023 1 23606
2 93024 1 23606
2 93025 1 23606
2 93026 1 23613
2 93027 1 23613
2 93028 1 23613
2 93029 1 23613
2 93030 1 23646
2 93031 1 23646
2 93032 1 23660
2 93033 1 23660
2 93034 1 23683
2 93035 1 23683
2 93036 1 23696
2 93037 1 23696
2 93038 1 23696
2 93039 1 23696
2 93040 1 23696
2 93041 1 23696
2 93042 1 23699
2 93043 1 23699
2 93044 1 23712
2 93045 1 23712
2 93046 1 23715
2 93047 1 23715
2 93048 1 23756
2 93049 1 23756
2 93050 1 23760
2 93051 1 23760
2 93052 1 23762
2 93053 1 23762
2 93054 1 23766
2 93055 1 23766
2 93056 1 23767
2 93057 1 23767
2 93058 1 23767
2 93059 1 23788
2 93060 1 23788
2 93061 1 23806
2 93062 1 23806
2 93063 1 23812
2 93064 1 23812
2 93065 1 23851
2 93066 1 23851
2 93067 1 23853
2 93068 1 23853
2 93069 1 23856
2 93070 1 23856
2 93071 1 23857
2 93072 1 23857
2 93073 1 23884
2 93074 1 23884
2 93075 1 23884
2 93076 1 23890
2 93077 1 23890
2 93078 1 23890
2 93079 1 23900
2 93080 1 23900
2 93081 1 23900
2 93082 1 23912
2 93083 1 23912
2 93084 1 23913
2 93085 1 23913
2 93086 1 23913
2 93087 1 23917
2 93088 1 23917
2 93089 1 23958
2 93090 1 23958
2 93091 1 23959
2 93092 1 23959
2 93093 1 23960
2 93094 1 23960
2 93095 1 23960
2 93096 1 23996
2 93097 1 23996
2 93098 1 24005
2 93099 1 24005
2 93100 1 24015
2 93101 1 24015
2 93102 1 24015
2 93103 1 24016
2 93104 1 24016
2 93105 1 24027
2 93106 1 24027
2 93107 1 24028
2 93108 1 24028
2 93109 1 24040
2 93110 1 24040
2 93111 1 24040
2 93112 1 24051
2 93113 1 24051
2 93114 1 24052
2 93115 1 24052
2 93116 1 24066
2 93117 1 24066
2 93118 1 24082
2 93119 1 24082
2 93120 1 24115
2 93121 1 24115
2 93122 1 24115
2 93123 1 24122
2 93124 1 24122
2 93125 1 24126
2 93126 1 24126
2 93127 1 24145
2 93128 1 24145
2 93129 1 24146
2 93130 1 24146
2 93131 1 24176
2 93132 1 24176
2 93133 1 24189
2 93134 1 24189
2 93135 1 24205
2 93136 1 24205
2 93137 1 24212
2 93138 1 24212
2 93139 1 24236
2 93140 1 24236
2 93141 1 24273
2 93142 1 24273
2 93143 1 24282
2 93144 1 24282
2 93145 1 24283
2 93146 1 24283
2 93147 1 24288
2 93148 1 24288
2 93149 1 24297
2 93150 1 24297
2 93151 1 24315
2 93152 1 24315
2 93153 1 24321
2 93154 1 24321
2 93155 1 24321
2 93156 1 24334
2 93157 1 24334
2 93158 1 24334
2 93159 1 24340
2 93160 1 24340
2 93161 1 24340
2 93162 1 24343
2 93163 1 24343
2 93164 1 24357
2 93165 1 24357
2 93166 1 24357
2 93167 1 24370
2 93168 1 24370
2 93169 1 24384
2 93170 1 24384
2 93171 1 24406
2 93172 1 24406
2 93173 1 24407
2 93174 1 24407
2 93175 1 24437
2 93176 1 24437
2 93177 1 24437
2 93178 1 24437
2 93179 1 24437
2 93180 1 24437
2 93181 1 24437
2 93182 1 24448
2 93183 1 24448
2 93184 1 24450
2 93185 1 24450
2 93186 1 24454
2 93187 1 24454
2 93188 1 24454
2 93189 1 24454
2 93190 1 24465
2 93191 1 24465
2 93192 1 24472
2 93193 1 24472
2 93194 1 24472
2 93195 1 24474
2 93196 1 24474
2 93197 1 24474
2 93198 1 24474
2 93199 1 24474
2 93200 1 24474
2 93201 1 24474
2 93202 1 24474
2 93203 1 24474
2 93204 1 24475
2 93205 1 24475
2 93206 1 24475
2 93207 1 24475
2 93208 1 24475
2 93209 1 24475
2 93210 1 24475
2 93211 1 24475
2 93212 1 24475
2 93213 1 24475
2 93214 1 24475
2 93215 1 24476
2 93216 1 24476
2 93217 1 24476
2 93218 1 24476
2 93219 1 24480
2 93220 1 24480
2 93221 1 24506
2 93222 1 24506
2 93223 1 24506
2 93224 1 24508
2 93225 1 24508
2 93226 1 24520
2 93227 1 24520
2 93228 1 24528
2 93229 1 24528
2 93230 1 24528
2 93231 1 24528
2 93232 1 24534
2 93233 1 24534
2 93234 1 24551
2 93235 1 24551
2 93236 1 24601
2 93237 1 24601
2 93238 1 24601
2 93239 1 24601
2 93240 1 24603
2 93241 1 24603
2 93242 1 24610
2 93243 1 24610
2 93244 1 24610
2 93245 1 24621
2 93246 1 24621
2 93247 1 24633
2 93248 1 24633
2 93249 1 24643
2 93250 1 24643
2 93251 1 24643
2 93252 1 24644
2 93253 1 24644
2 93254 1 24644
2 93255 1 24644
2 93256 1 24671
2 93257 1 24671
2 93258 1 24671
2 93259 1 24671
2 93260 1 24674
2 93261 1 24674
2 93262 1 24674
2 93263 1 24687
2 93264 1 24687
2 93265 1 24701
2 93266 1 24701
2 93267 1 24701
2 93268 1 24701
2 93269 1 24701
2 93270 1 24701
2 93271 1 24701
2 93272 1 24702
2 93273 1 24702
2 93274 1 24702
2 93275 1 24717
2 93276 1 24717
2 93277 1 24718
2 93278 1 24718
2 93279 1 24732
2 93280 1 24732
2 93281 1 24732
2 93282 1 24761
2 93283 1 24761
2 93284 1 24782
2 93285 1 24782
2 93286 1 24800
2 93287 1 24800
2 93288 1 24824
2 93289 1 24824
2 93290 1 24824
2 93291 1 24838
2 93292 1 24838
2 93293 1 24847
2 93294 1 24847
2 93295 1 24847
2 93296 1 24868
2 93297 1 24868
2 93298 1 24868
2 93299 1 24889
2 93300 1 24889
2 93301 1 24903
2 93302 1 24903
2 93303 1 24904
2 93304 1 24904
2 93305 1 24912
2 93306 1 24912
2 93307 1 24916
2 93308 1 24916
2 93309 1 24916
2 93310 1 24916
2 93311 1 24916
2 93312 1 24916
2 93313 1 24918
2 93314 1 24918
2 93315 1 24919
2 93316 1 24919
2 93317 1 24945
2 93318 1 24945
2 93319 1 24946
2 93320 1 24946
2 93321 1 24947
2 93322 1 24947
2 93323 1 24966
2 93324 1 24966
2 93325 1 24995
2 93326 1 24995
2 93327 1 24995
2 93328 1 24995
2 93329 1 24995
2 93330 1 24995
2 93331 1 25003
2 93332 1 25003
2 93333 1 25003
2 93334 1 25039
2 93335 1 25039
2 93336 1 25039
2 93337 1 25039
2 93338 1 25040
2 93339 1 25040
2 93340 1 25069
2 93341 1 25069
2 93342 1 25075
2 93343 1 25075
2 93344 1 25088
2 93345 1 25088
2 93346 1 25127
2 93347 1 25127
2 93348 1 25139
2 93349 1 25139
2 93350 1 25139
2 93351 1 25143
2 93352 1 25143
2 93353 1 25158
2 93354 1 25158
2 93355 1 25184
2 93356 1 25184
2 93357 1 25184
2 93358 1 25184
2 93359 1 25194
2 93360 1 25194
2 93361 1 25195
2 93362 1 25195
2 93363 1 25200
2 93364 1 25200
2 93365 1 25200
2 93366 1 25200
2 93367 1 25200
2 93368 1 25200
2 93369 1 25200
2 93370 1 25200
2 93371 1 25201
2 93372 1 25201
2 93373 1 25201
2 93374 1 25201
2 93375 1 25201
2 93376 1 25201
2 93377 1 25201
2 93378 1 25223
2 93379 1 25223
2 93380 1 25241
2 93381 1 25241
2 93382 1 25241
2 93383 1 25241
2 93384 1 25241
2 93385 1 25241
2 93386 1 25241
2 93387 1 25246
2 93388 1 25246
2 93389 1 25246
2 93390 1 25246
2 93391 1 25263
2 93392 1 25263
2 93393 1 25346
2 93394 1 25346
2 93395 1 25346
2 93396 1 25399
2 93397 1 25399
2 93398 1 25399
2 93399 1 25399
2 93400 1 25405
2 93401 1 25405
2 93402 1 25406
2 93403 1 25406
2 93404 1 25412
2 93405 1 25412
2 93406 1 25412
2 93407 1 25412
2 93408 1 25412
2 93409 1 25426
2 93410 1 25426
2 93411 1 25463
2 93412 1 25463
2 93413 1 25483
2 93414 1 25483
2 93415 1 25485
2 93416 1 25485
2 93417 1 25496
2 93418 1 25496
2 93419 1 25496
2 93420 1 25517
2 93421 1 25517
2 93422 1 25517
2 93423 1 25517
2 93424 1 25517
2 93425 1 25532
2 93426 1 25532
2 93427 1 25532
2 93428 1 25532
2 93429 1 25532
2 93430 1 25553
2 93431 1 25553
2 93432 1 25556
2 93433 1 25556
2 93434 1 25565
2 93435 1 25565
2 93436 1 25578
2 93437 1 25578
2 93438 1 25579
2 93439 1 25579
2 93440 1 25579
2 93441 1 25579
2 93442 1 25579
2 93443 1 25606
2 93444 1 25606
2 93445 1 25636
2 93446 1 25636
2 93447 1 25663
2 93448 1 25663
2 93449 1 25666
2 93450 1 25666
2 93451 1 25700
2 93452 1 25700
2 93453 1 25711
2 93454 1 25711
2 93455 1 25712
2 93456 1 25712
2 93457 1 25728
2 93458 1 25728
2 93459 1 25728
2 93460 1 25728
2 93461 1 25737
2 93462 1 25737
2 93463 1 25776
2 93464 1 25776
2 93465 1 25794
2 93466 1 25794
2 93467 1 25794
2 93468 1 25797
2 93469 1 25797
2 93470 1 25812
2 93471 1 25812
2 93472 1 25924
2 93473 1 25924
2 93474 1 25924
2 93475 1 25927
2 93476 1 25927
2 93477 1 25986
2 93478 1 25986
2 93479 1 25986
2 93480 1 26001
2 93481 1 26001
2 93482 1 26034
2 93483 1 26034
2 93484 1 26040
2 93485 1 26040
2 93486 1 26048
2 93487 1 26048
2 93488 1 26048
2 93489 1 26048
2 93490 1 26048
2 93491 1 26090
2 93492 1 26090
2 93493 1 26098
2 93494 1 26098
2 93495 1 26107
2 93496 1 26107
2 93497 1 26107
2 93498 1 26116
2 93499 1 26116
2 93500 1 26118
2 93501 1 26118
2 93502 1 26119
2 93503 1 26119
2 93504 1 26120
2 93505 1 26120
2 93506 1 26120
2 93507 1 26120
2 93508 1 26120
2 93509 1 26123
2 93510 1 26123
2 93511 1 26123
2 93512 1 26143
2 93513 1 26143
2 93514 1 26143
2 93515 1 26158
2 93516 1 26158
2 93517 1 26172
2 93518 1 26172
2 93519 1 26193
2 93520 1 26193
2 93521 1 26193
2 93522 1 26202
2 93523 1 26202
2 93524 1 26202
2 93525 1 26214
2 93526 1 26214
2 93527 1 26225
2 93528 1 26225
2 93529 1 26226
2 93530 1 26226
2 93531 1 26233
2 93532 1 26233
2 93533 1 26233
2 93534 1 26233
2 93535 1 26233
2 93536 1 26233
2 93537 1 26234
2 93538 1 26234
2 93539 1 26234
2 93540 1 26234
2 93541 1 26235
2 93542 1 26235
2 93543 1 26242
2 93544 1 26242
2 93545 1 26242
2 93546 1 26242
2 93547 1 26242
2 93548 1 26242
2 93549 1 26299
2 93550 1 26299
2 93551 1 26304
2 93552 1 26304
2 93553 1 26318
2 93554 1 26318
2 93555 1 26330
2 93556 1 26330
2 93557 1 26338
2 93558 1 26338
2 93559 1 26372
2 93560 1 26372
2 93561 1 26372
2 93562 1 26381
2 93563 1 26381
2 93564 1 26382
2 93565 1 26382
2 93566 1 26399
2 93567 1 26399
2 93568 1 26399
2 93569 1 26412
2 93570 1 26412
2 93571 1 26421
2 93572 1 26421
2 93573 1 26423
2 93574 1 26423
2 93575 1 26441
2 93576 1 26441
2 93577 1 26441
2 93578 1 26441
2 93579 1 26442
2 93580 1 26442
2 93581 1 26445
2 93582 1 26445
2 93583 1 26445
2 93584 1 26445
2 93585 1 26446
2 93586 1 26446
2 93587 1 26446
2 93588 1 26446
2 93589 1 26448
2 93590 1 26448
2 93591 1 26455
2 93592 1 26455
2 93593 1 26455
2 93594 1 26455
2 93595 1 26456
2 93596 1 26456
2 93597 1 26456
2 93598 1 26479
2 93599 1 26479
2 93600 1 26480
2 93601 1 26480
2 93602 1 26495
2 93603 1 26495
2 93604 1 26523
2 93605 1 26523
2 93606 1 26540
2 93607 1 26540
2 93608 1 26549
2 93609 1 26549
2 93610 1 26549
2 93611 1 26567
2 93612 1 26567
2 93613 1 26585
2 93614 1 26585
2 93615 1 26597
2 93616 1 26597
2 93617 1 26626
2 93618 1 26626
2 93619 1 26626
2 93620 1 26637
2 93621 1 26637
2 93622 1 26649
2 93623 1 26649
2 93624 1 26649
2 93625 1 26671
2 93626 1 26671
2 93627 1 26671
2 93628 1 26671
2 93629 1 26671
2 93630 1 26671
2 93631 1 26671
2 93632 1 26671
2 93633 1 26671
2 93634 1 26682
2 93635 1 26682
2 93636 1 26698
2 93637 1 26698
2 93638 1 26699
2 93639 1 26699
2 93640 1 26699
2 93641 1 26699
2 93642 1 26699
2 93643 1 26701
2 93644 1 26701
2 93645 1 26717
2 93646 1 26717
2 93647 1 26718
2 93648 1 26718
2 93649 1 26742
2 93650 1 26742
2 93651 1 26742
2 93652 1 26760
2 93653 1 26760
2 93654 1 26760
2 93655 1 26760
2 93656 1 26769
2 93657 1 26769
2 93658 1 26777
2 93659 1 26777
2 93660 1 26777
2 93661 1 26777
2 93662 1 26779
2 93663 1 26779
2 93664 1 26779
2 93665 1 26795
2 93666 1 26795
2 93667 1 26798
2 93668 1 26798
2 93669 1 26799
2 93670 1 26799
2 93671 1 26799
2 93672 1 26808
2 93673 1 26808
2 93674 1 26808
2 93675 1 26808
2 93676 1 26816
2 93677 1 26816
2 93678 1 26835
2 93679 1 26835
2 93680 1 26843
2 93681 1 26843
2 93682 1 26852
2 93683 1 26852
2 93684 1 26861
2 93685 1 26861
2 93686 1 26876
2 93687 1 26876
2 93688 1 26876
2 93689 1 26893
2 93690 1 26893
2 93691 1 26893
2 93692 1 26905
2 93693 1 26905
2 93694 1 26906
2 93695 1 26906
2 93696 1 26907
2 93697 1 26907
2 93698 1 26907
2 93699 1 26907
2 93700 1 26908
2 93701 1 26908
2 93702 1 26915
2 93703 1 26915
2 93704 1 26925
2 93705 1 26925
2 93706 1 26925
2 93707 1 26926
2 93708 1 26926
2 93709 1 26927
2 93710 1 26927
2 93711 1 26939
2 93712 1 26939
2 93713 1 26958
2 93714 1 26958
2 93715 1 26958
2 93716 1 26958
2 93717 1 26959
2 93718 1 26959
2 93719 1 26959
2 93720 1 26989
2 93721 1 26989
2 93722 1 26989
2 93723 1 27005
2 93724 1 27005
2 93725 1 27065
2 93726 1 27065
2 93727 1 27065
2 93728 1 27065
2 93729 1 27065
2 93730 1 27082
2 93731 1 27082
2 93732 1 27082
2 93733 1 27083
2 93734 1 27083
2 93735 1 27086
2 93736 1 27086
2 93737 1 27086
2 93738 1 27086
2 93739 1 27093
2 93740 1 27093
2 93741 1 27093
2 93742 1 27093
2 93743 1 27093
2 93744 1 27107
2 93745 1 27107
2 93746 1 27123
2 93747 1 27123
2 93748 1 27136
2 93749 1 27136
2 93750 1 27167
2 93751 1 27167
2 93752 1 27168
2 93753 1 27168
2 93754 1 27168
2 93755 1 27168
2 93756 1 27168
2 93757 1 27184
2 93758 1 27184
2 93759 1 27185
2 93760 1 27185
2 93761 1 27185
2 93762 1 27185
2 93763 1 27211
2 93764 1 27211
2 93765 1 27212
2 93766 1 27212
2 93767 1 27212
2 93768 1 27212
2 93769 1 27212
2 93770 1 27226
2 93771 1 27226
2 93772 1 27226
2 93773 1 27226
2 93774 1 27226
2 93775 1 27226
2 93776 1 27226
2 93777 1 27240
2 93778 1 27240
2 93779 1 27240
2 93780 1 27283
2 93781 1 27283
2 93782 1 27300
2 93783 1 27300
2 93784 1 27300
2 93785 1 27310
2 93786 1 27310
2 93787 1 27317
2 93788 1 27317
2 93789 1 27335
2 93790 1 27335
2 93791 1 27341
2 93792 1 27341
2 93793 1 27341
2 93794 1 27341
2 93795 1 27341
2 93796 1 27403
2 93797 1 27403
2 93798 1 27406
2 93799 1 27406
2 93800 1 27406
2 93801 1 27406
2 93802 1 27406
2 93803 1 27407
2 93804 1 27407
2 93805 1 27407
2 93806 1 27440
2 93807 1 27440
2 93808 1 27463
2 93809 1 27463
2 93810 1 27486
2 93811 1 27486
2 93812 1 27504
2 93813 1 27504
2 93814 1 27524
2 93815 1 27524
2 93816 1 27537
2 93817 1 27537
2 93818 1 27542
2 93819 1 27542
2 93820 1 27570
2 93821 1 27570
2 93822 1 27570
2 93823 1 27570
2 93824 1 27571
2 93825 1 27571
2 93826 1 27647
2 93827 1 27647
2 93828 1 27651
2 93829 1 27651
2 93830 1 27667
2 93831 1 27667
2 93832 1 27668
2 93833 1 27668
2 93834 1 27702
2 93835 1 27702
2 93836 1 27702
2 93837 1 27703
2 93838 1 27703
2 93839 1 27703
2 93840 1 27703
2 93841 1 27713
2 93842 1 27713
2 93843 1 27713
2 93844 1 27713
2 93845 1 27730
2 93846 1 27730
2 93847 1 27767
2 93848 1 27767
2 93849 1 27780
2 93850 1 27780
2 93851 1 27780
2 93852 1 27781
2 93853 1 27781
2 93854 1 27785
2 93855 1 27785
2 93856 1 27787
2 93857 1 27787
2 93858 1 27814
2 93859 1 27814
2 93860 1 27827
2 93861 1 27827
2 93862 1 27835
2 93863 1 27835
2 93864 1 27840
2 93865 1 27840
2 93866 1 27840
2 93867 1 27864
2 93868 1 27864
2 93869 1 27864
2 93870 1 27864
2 93871 1 27865
2 93872 1 27865
2 93873 1 27865
2 93874 1 27865
2 93875 1 27891
2 93876 1 27891
2 93877 1 27891
2 93878 1 27905
2 93879 1 27905
2 93880 1 27905
2 93881 1 27913
2 93882 1 27913
2 93883 1 27930
2 93884 1 27930
2 93885 1 27931
2 93886 1 27931
2 93887 1 27936
2 93888 1 27936
2 93889 1 27936
2 93890 1 27936
2 93891 1 27937
2 93892 1 27937
2 93893 1 27937
2 93894 1 27937
2 93895 1 27945
2 93896 1 27945
2 93897 1 27953
2 93898 1 27953
2 93899 1 27955
2 93900 1 27955
2 93901 1 27960
2 93902 1 27960
2 93903 1 27981
2 93904 1 27981
2 93905 1 27981
2 93906 1 27983
2 93907 1 27983
2 93908 1 28021
2 93909 1 28021
2 93910 1 28059
2 93911 1 28059
2 93912 1 28061
2 93913 1 28061
2 93914 1 28076
2 93915 1 28076
2 93916 1 28076
2 93917 1 28076
2 93918 1 28086
2 93919 1 28086
2 93920 1 28090
2 93921 1 28090
2 93922 1 28090
2 93923 1 28114
2 93924 1 28114
2 93925 1 28115
2 93926 1 28115
2 93927 1 28131
2 93928 1 28131
2 93929 1 28131
2 93930 1 28131
2 93931 1 28131
2 93932 1 28131
2 93933 1 28131
2 93934 1 28153
2 93935 1 28153
2 93936 1 28156
2 93937 1 28156
2 93938 1 28156
2 93939 1 28156
2 93940 1 28156
2 93941 1 28161
2 93942 1 28161
2 93943 1 28162
2 93944 1 28162
2 93945 1 28170
2 93946 1 28170
2 93947 1 28204
2 93948 1 28204
2 93949 1 28204
2 93950 1 28207
2 93951 1 28207
2 93952 1 28215
2 93953 1 28215
2 93954 1 28229
2 93955 1 28229
2 93956 1 28243
2 93957 1 28243
2 93958 1 28277
2 93959 1 28277
2 93960 1 28327
2 93961 1 28327
2 93962 1 28330
2 93963 1 28330
2 93964 1 28347
2 93965 1 28347
2 93966 1 28365
2 93967 1 28365
2 93968 1 28365
2 93969 1 28365
2 93970 1 28368
2 93971 1 28368
2 93972 1 28368
2 93973 1 28372
2 93974 1 28372
2 93975 1 28372
2 93976 1 28372
2 93977 1 28372
2 93978 1 28373
2 93979 1 28373
2 93980 1 28398
2 93981 1 28398
2 93982 1 28398
2 93983 1 28398
2 93984 1 28398
2 93985 1 28399
2 93986 1 28399
2 93987 1 28399
2 93988 1 28401
2 93989 1 28401
2 93990 1 28417
2 93991 1 28417
2 93992 1 28417
2 93993 1 28453
2 93994 1 28453
2 93995 1 28494
2 93996 1 28494
2 93997 1 28498
2 93998 1 28498
2 93999 1 28516
2 94000 1 28516
2 94001 1 28516
2 94002 1 28524
2 94003 1 28524
2 94004 1 28524
2 94005 1 28559
2 94006 1 28559
2 94007 1 28584
2 94008 1 28584
2 94009 1 28594
2 94010 1 28594
2 94011 1 28637
2 94012 1 28637
2 94013 1 28657
2 94014 1 28657
2 94015 1 28702
2 94016 1 28702
2 94017 1 28702
2 94018 1 28718
2 94019 1 28718
2 94020 1 28718
2 94021 1 28718
2 94022 1 28719
2 94023 1 28719
2 94024 1 28737
2 94025 1 28737
2 94026 1 28752
2 94027 1 28752
2 94028 1 28813
2 94029 1 28813
2 94030 1 28827
2 94031 1 28827
2 94032 1 28839
2 94033 1 28839
2 94034 1 28843
2 94035 1 28843
2 94036 1 28844
2 94037 1 28844
2 94038 1 28889
2 94039 1 28889
2 94040 1 28925
2 94041 1 28925
2 94042 1 28925
2 94043 1 28960
2 94044 1 28960
2 94045 1 28960
2 94046 1 29050
2 94047 1 29050
2 94048 1 29056
2 94049 1 29056
2 94050 1 29156
2 94051 1 29156
2 94052 1 29201
2 94053 1 29201
2 94054 1 29201
2 94055 1 29228
2 94056 1 29228
2 94057 1 29228
2 94058 1 29235
2 94059 1 29235
2 94060 1 29250
2 94061 1 29250
2 94062 1 29277
2 94063 1 29277
2 94064 1 29285
2 94065 1 29285
2 94066 1 29290
2 94067 1 29290
2 94068 1 29293
2 94069 1 29293
2 94070 1 29293
2 94071 1 29340
2 94072 1 29340
2 94073 1 29361
2 94074 1 29361
2 94075 1 29362
2 94076 1 29362
2 94077 1 29364
2 94078 1 29364
2 94079 1 29365
2 94080 1 29365
2 94081 1 29365
2 94082 1 29365
2 94083 1 29365
2 94084 1 29365
2 94085 1 29365
2 94086 1 29384
2 94087 1 29384
2 94088 1 29385
2 94089 1 29385
2 94090 1 29397
2 94091 1 29397
2 94092 1 29397
2 94093 1 29432
2 94094 1 29432
2 94095 1 29432
2 94096 1 29440
2 94097 1 29440
2 94098 1 29459
2 94099 1 29459
2 94100 1 29469
2 94101 1 29469
2 94102 1 29469
2 94103 1 29469
2 94104 1 29469
2 94105 1 29470
2 94106 1 29470
2 94107 1 29491
2 94108 1 29491
2 94109 1 29491
2 94110 1 29491
2 94111 1 29497
2 94112 1 29497
2 94113 1 29546
2 94114 1 29546
2 94115 1 29547
2 94116 1 29547
2 94117 1 29563
2 94118 1 29563
2 94119 1 29563
2 94120 1 29571
2 94121 1 29571
2 94122 1 29571
2 94123 1 29650
2 94124 1 29650
2 94125 1 29690
2 94126 1 29690
2 94127 1 29694
2 94128 1 29694
2 94129 1 29694
2 94130 1 29694
2 94131 1 29695
2 94132 1 29695
2 94133 1 29717
2 94134 1 29717
2 94135 1 29722
2 94136 1 29722
2 94137 1 29722
2 94138 1 29722
2 94139 1 29722
2 94140 1 29722
2 94141 1 29722
2 94142 1 29722
2 94143 1 29722
2 94144 1 29722
2 94145 1 29738
2 94146 1 29738
2 94147 1 29746
2 94148 1 29746
2 94149 1 29746
2 94150 1 29746
2 94151 1 29746
2 94152 1 29746
2 94153 1 29766
2 94154 1 29766
2 94155 1 29768
2 94156 1 29768
2 94157 1 29768
2 94158 1 29769
2 94159 1 29769
2 94160 1 29769
2 94161 1 29769
2 94162 1 29769
2 94163 1 29769
2 94164 1 29769
2 94165 1 29770
2 94166 1 29770
2 94167 1 29770
2 94168 1 29770
2 94169 1 29770
2 94170 1 29773
2 94171 1 29773
2 94172 1 29773
2 94173 1 29774
2 94174 1 29774
2 94175 1 29774
2 94176 1 29774
2 94177 1 29774
2 94178 1 29774
2 94179 1 29774
2 94180 1 29774
2 94181 1 29774
2 94182 1 29774
2 94183 1 29774
2 94184 1 29774
2 94185 1 29774
2 94186 1 29774
2 94187 1 29774
2 94188 1 29774
2 94189 1 29774
2 94190 1 29776
2 94191 1 29776
2 94192 1 29787
2 94193 1 29787
2 94194 1 29787
2 94195 1 29795
2 94196 1 29795
2 94197 1 29795
2 94198 1 29797
2 94199 1 29797
2 94200 1 29797
2 94201 1 29797
2 94202 1 29807
2 94203 1 29807
2 94204 1 29807
2 94205 1 29816
2 94206 1 29816
2 94207 1 29816
2 94208 1 29816
2 94209 1 29816
2 94210 1 29816
2 94211 1 29816
2 94212 1 29816
2 94213 1 29816
2 94214 1 29816
2 94215 1 29816
2 94216 1 29816
2 94217 1 29816
2 94218 1 29816
2 94219 1 29816
2 94220 1 29816
2 94221 1 29816
2 94222 1 29816
2 94223 1 29816
2 94224 1 29816
2 94225 1 29817
2 94226 1 29817
2 94227 1 29817
2 94228 1 29817
2 94229 1 29817
2 94230 1 29817
2 94231 1 29817
2 94232 1 29818
2 94233 1 29818
2 94234 1 29818
2 94235 1 29818
2 94236 1 29819
2 94237 1 29819
2 94238 1 29819
2 94239 1 29820
2 94240 1 29820
2 94241 1 29821
2 94242 1 29821
2 94243 1 29821
2 94244 1 29822
2 94245 1 29822
2 94246 1 29822
2 94247 1 29838
2 94248 1 29838
2 94249 1 29846
2 94250 1 29846
2 94251 1 29846
2 94252 1 29846
2 94253 1 29846
2 94254 1 29846
2 94255 1 29846
2 94256 1 29846
2 94257 1 29846
2 94258 1 29846
2 94259 1 29848
2 94260 1 29848
2 94261 1 29848
2 94262 1 29857
2 94263 1 29857
2 94264 1 29865
2 94265 1 29865
2 94266 1 29891
2 94267 1 29891
2 94268 1 29892
2 94269 1 29892
2 94270 1 29894
2 94271 1 29894
2 94272 1 29896
2 94273 1 29896
2 94274 1 29896
2 94275 1 29896
2 94276 1 29896
2 94277 1 29896
2 94278 1 29897
2 94279 1 29897
2 94280 1 29897
2 94281 1 29903
2 94282 1 29903
2 94283 1 29903
2 94284 1 29905
2 94285 1 29905
2 94286 1 29905
2 94287 1 29905
2 94288 1 29905
2 94289 1 29910
2 94290 1 29910
2 94291 1 29924
2 94292 1 29924
2 94293 1 29931
2 94294 1 29931
2 94295 1 29940
2 94296 1 29940
2 94297 1 29940
2 94298 1 29941
2 94299 1 29941
2 94300 1 29943
2 94301 1 29943
2 94302 1 29965
2 94303 1 29965
2 94304 1 29978
2 94305 1 29978
2 94306 1 30034
2 94307 1 30034
2 94308 1 30047
2 94309 1 30047
2 94310 1 30052
2 94311 1 30052
2 94312 1 30052
2 94313 1 30052
2 94314 1 30079
2 94315 1 30079
2 94316 1 30082
2 94317 1 30082
2 94318 1 30087
2 94319 1 30087
2 94320 1 30087
2 94321 1 30087
2 94322 1 30087
2 94323 1 30109
2 94324 1 30109
2 94325 1 30147
2 94326 1 30147
2 94327 1 30147
2 94328 1 30159
2 94329 1 30159
2 94330 1 30175
2 94331 1 30175
2 94332 1 30184
2 94333 1 30184
2 94334 1 30184
2 94335 1 30184
2 94336 1 30184
2 94337 1 30217
2 94338 1 30217
2 94339 1 30231
2 94340 1 30231
2 94341 1 30234
2 94342 1 30234
2 94343 1 30258
2 94344 1 30258
2 94345 1 30258
2 94346 1 30258
2 94347 1 30258
2 94348 1 30258
2 94349 1 30258
2 94350 1 30258
2 94351 1 30258
2 94352 1 30258
2 94353 1 30258
2 94354 1 30258
2 94355 1 30259
2 94356 1 30259
2 94357 1 30260
2 94358 1 30260
2 94359 1 30268
2 94360 1 30268
2 94361 1 30268
2 94362 1 30270
2 94363 1 30270
2 94364 1 30298
2 94365 1 30298
2 94366 1 30336
2 94367 1 30336
2 94368 1 30359
2 94369 1 30359
2 94370 1 30372
2 94371 1 30372
2 94372 1 30377
2 94373 1 30377
2 94374 1 30378
2 94375 1 30378
2 94376 1 30392
2 94377 1 30392
2 94378 1 30393
2 94379 1 30393
2 94380 1 30415
2 94381 1 30415
2 94382 1 30426
2 94383 1 30426
2 94384 1 30436
2 94385 1 30436
2 94386 1 30444
2 94387 1 30444
2 94388 1 30445
2 94389 1 30445
2 94390 1 30462
2 94391 1 30462
2 94392 1 30462
2 94393 1 30463
2 94394 1 30463
2 94395 1 30463
2 94396 1 30503
2 94397 1 30503
2 94398 1 30554
2 94399 1 30554
2 94400 1 30554
2 94401 1 30572
2 94402 1 30572
2 94403 1 30580
2 94404 1 30580
2 94405 1 30580
2 94406 1 30580
2 94407 1 30580
2 94408 1 30580
2 94409 1 30580
2 94410 1 30580
2 94411 1 30581
2 94412 1 30581
2 94413 1 30582
2 94414 1 30582
2 94415 1 30590
2 94416 1 30590
2 94417 1 30617
2 94418 1 30617
2 94419 1 30617
2 94420 1 30618
2 94421 1 30618
2 94422 1 30618
2 94423 1 30619
2 94424 1 30619
2 94425 1 30651
2 94426 1 30651
2 94427 1 30655
2 94428 1 30655
2 94429 1 30686
2 94430 1 30686
2 94431 1 30695
2 94432 1 30695
2 94433 1 30695
2 94434 1 30709
2 94435 1 30709
2 94436 1 30709
2 94437 1 30709
2 94438 1 30710
2 94439 1 30710
2 94440 1 30710
2 94441 1 30710
2 94442 1 30710
2 94443 1 30710
2 94444 1 30710
2 94445 1 30745
2 94446 1 30745
2 94447 1 30775
2 94448 1 30775
2 94449 1 30775
2 94450 1 30775
2 94451 1 30776
2 94452 1 30776
2 94453 1 30783
2 94454 1 30783
2 94455 1 30806
2 94456 1 30806
2 94457 1 30808
2 94458 1 30808
2 94459 1 30814
2 94460 1 30814
2 94461 1 30814
2 94462 1 30814
2 94463 1 30827
2 94464 1 30827
2 94465 1 30836
2 94466 1 30836
2 94467 1 30844
2 94468 1 30844
2 94469 1 30867
2 94470 1 30867
2 94471 1 30867
2 94472 1 30867
2 94473 1 30867
2 94474 1 30867
2 94475 1 30897
2 94476 1 30897
2 94477 1 30917
2 94478 1 30917
2 94479 1 30917
2 94480 1 30940
2 94481 1 30940
2 94482 1 30948
2 94483 1 30948
2 94484 1 30951
2 94485 1 30951
2 94486 1 30951
2 94487 1 30951
2 94488 1 30951
2 94489 1 30968
2 94490 1 30968
2 94491 1 31030
2 94492 1 31030
2 94493 1 31031
2 94494 1 31031
2 94495 1 31033
2 94496 1 31033
2 94497 1 31041
2 94498 1 31041
2 94499 1 31041
2 94500 1 31085
2 94501 1 31085
2 94502 1 31085
2 94503 1 31085
2 94504 1 31104
2 94505 1 31104
2 94506 1 31106
2 94507 1 31106
2 94508 1 31107
2 94509 1 31107
2 94510 1 31108
2 94511 1 31108
2 94512 1 31125
2 94513 1 31125
2 94514 1 31130
2 94515 1 31130
2 94516 1 31130
2 94517 1 31130
2 94518 1 31130
2 94519 1 31148
2 94520 1 31148
2 94521 1 31164
2 94522 1 31164
2 94523 1 31199
2 94524 1 31199
2 94525 1 31223
2 94526 1 31223
2 94527 1 31231
2 94528 1 31231
2 94529 1 31234
2 94530 1 31234
2 94531 1 31270
2 94532 1 31270
2 94533 1 31270
2 94534 1 31270
2 94535 1 31271
2 94536 1 31271
2 94537 1 31272
2 94538 1 31272
2 94539 1 31333
2 94540 1 31333
2 94541 1 31353
2 94542 1 31353
2 94543 1 31353
2 94544 1 31379
2 94545 1 31379
2 94546 1 31417
2 94547 1 31417
2 94548 1 31422
2 94549 1 31422
2 94550 1 31422
2 94551 1 31458
2 94552 1 31458
2 94553 1 31479
2 94554 1 31479
2 94555 1 31479
2 94556 1 31512
2 94557 1 31512
2 94558 1 31512
2 94559 1 31519
2 94560 1 31519
2 94561 1 31545
2 94562 1 31545
2 94563 1 31546
2 94564 1 31546
2 94565 1 31547
2 94566 1 31547
2 94567 1 31548
2 94568 1 31548
2 94569 1 31548
2 94570 1 31580
2 94571 1 31580
2 94572 1 31619
2 94573 1 31619
2 94574 1 31628
2 94575 1 31628
2 94576 1 31628
2 94577 1 31629
2 94578 1 31629
2 94579 1 31631
2 94580 1 31631
2 94581 1 31631
2 94582 1 31632
2 94583 1 31632
2 94584 1 31632
2 94585 1 31632
2 94586 1 31633
2 94587 1 31633
2 94588 1 31759
2 94589 1 31759
2 94590 1 31779
2 94591 1 31779
2 94592 1 31808
2 94593 1 31808
2 94594 1 31809
2 94595 1 31809
2 94596 1 31820
2 94597 1 31820
2 94598 1 31823
2 94599 1 31823
2 94600 1 31832
2 94601 1 31832
2 94602 1 31833
2 94603 1 31833
2 94604 1 31884
2 94605 1 31884
2 94606 1 31884
2 94607 1 31884
2 94608 1 31884
2 94609 1 31884
2 94610 1 31884
2 94611 1 31885
2 94612 1 31885
2 94613 1 31885
2 94614 1 31913
2 94615 1 31913
2 94616 1 31914
2 94617 1 31914
2 94618 1 31918
2 94619 1 31918
2 94620 1 31918
2 94621 1 31920
2 94622 1 31920
2 94623 1 31924
2 94624 1 31924
2 94625 1 31940
2 94626 1 31940
2 94627 1 31940
2 94628 1 31962
2 94629 1 31962
2 94630 1 31973
2 94631 1 31973
2 94632 1 31985
2 94633 1 31985
2 94634 1 31985
2 94635 1 31985
2 94636 1 31985
2 94637 1 31985
2 94638 1 31985
2 94639 1 31986
2 94640 1 31986
2 94641 1 31987
2 94642 1 31987
2 94643 1 32002
2 94644 1 32002
2 94645 1 32002
2 94646 1 32002
2 94647 1 32002
2 94648 1 32002
2 94649 1 32003
2 94650 1 32003
2 94651 1 32003
2 94652 1 32003
2 94653 1 32003
2 94654 1 32003
2 94655 1 32003
2 94656 1 32014
2 94657 1 32014
2 94658 1 32024
2 94659 1 32024
2 94660 1 32025
2 94661 1 32025
2 94662 1 32025
2 94663 1 32027
2 94664 1 32027
2 94665 1 32028
2 94666 1 32028
2 94667 1 32028
2 94668 1 32039
2 94669 1 32039
2 94670 1 32048
2 94671 1 32048
2 94672 1 32058
2 94673 1 32058
2 94674 1 32060
2 94675 1 32060
2 94676 1 32061
2 94677 1 32061
2 94678 1 32086
2 94679 1 32086
2 94680 1 32107
2 94681 1 32107
2 94682 1 32136
2 94683 1 32136
2 94684 1 32144
2 94685 1 32144
2 94686 1 32151
2 94687 1 32151
2 94688 1 32152
2 94689 1 32152
2 94690 1 32166
2 94691 1 32166
2 94692 1 32178
2 94693 1 32178
2 94694 1 32186
2 94695 1 32186
2 94696 1 32186
2 94697 1 32186
2 94698 1 32189
2 94699 1 32189
2 94700 1 32190
2 94701 1 32190
2 94702 1 32190
2 94703 1 32306
2 94704 1 32306
2 94705 1 32344
2 94706 1 32344
2 94707 1 32378
2 94708 1 32378
2 94709 1 32383
2 94710 1 32383
2 94711 1 32406
2 94712 1 32406
2 94713 1 32414
2 94714 1 32414
2 94715 1 32414
2 94716 1 32414
2 94717 1 32414
2 94718 1 32414
2 94719 1 32414
2 94720 1 32414
2 94721 1 32414
2 94722 1 32414
2 94723 1 32414
2 94724 1 32414
2 94725 1 32414
2 94726 1 32414
2 94727 1 32414
2 94728 1 32437
2 94729 1 32437
2 94730 1 32437
2 94731 1 32437
2 94732 1 32437
2 94733 1 32437
2 94734 1 32437
2 94735 1 32437
2 94736 1 32437
2 94737 1 32438
2 94738 1 32438
2 94739 1 32440
2 94740 1 32440
2 94741 1 32440
2 94742 1 32466
2 94743 1 32466
2 94744 1 32466
2 94745 1 32484
2 94746 1 32484
2 94747 1 32492
2 94748 1 32492
2 94749 1 32492
2 94750 1 32492
2 94751 1 32492
2 94752 1 32492
2 94753 1 32492
2 94754 1 32492
2 94755 1 32492
2 94756 1 32492
2 94757 1 32492
2 94758 1 32492
2 94759 1 32492
2 94760 1 32492
2 94761 1 32492
2 94762 1 32492
2 94763 1 32492
2 94764 1 32492
2 94765 1 32492
2 94766 1 32492
2 94767 1 32492
2 94768 1 32492
2 94769 1 32492
2 94770 1 32492
2 94771 1 32492
2 94772 1 32492
2 94773 1 32492
2 94774 1 32492
2 94775 1 32492
2 94776 1 32524
2 94777 1 32524
2 94778 1 32533
2 94779 1 32533
2 94780 1 32600
2 94781 1 32600
2 94782 1 32600
2 94783 1 32600
2 94784 1 32601
2 94785 1 32601
2 94786 1 32617
2 94787 1 32617
2 94788 1 32627
2 94789 1 32627
2 94790 1 32628
2 94791 1 32628
2 94792 1 32628
2 94793 1 32641
2 94794 1 32641
2 94795 1 32656
2 94796 1 32656
2 94797 1 32656
2 94798 1 32663
2 94799 1 32663
2 94800 1 32663
2 94801 1 32696
2 94802 1 32696
2 94803 1 32700
2 94804 1 32700
2 94805 1 32700
2 94806 1 32701
2 94807 1 32701
2 94808 1 32704
2 94809 1 32704
2 94810 1 32717
2 94811 1 32717
2 94812 1 32720
2 94813 1 32720
2 94814 1 32766
2 94815 1 32766
2 94816 1 32769
2 94817 1 32769
2 94818 1 32775
2 94819 1 32775
2 94820 1 32812
2 94821 1 32812
2 94822 1 32832
2 94823 1 32832
2 94824 1 32863
2 94825 1 32863
2 94826 1 32863
2 94827 1 32863
2 94828 1 32863
2 94829 1 32866
2 94830 1 32866
2 94831 1 32896
2 94832 1 32896
2 94833 1 32897
2 94834 1 32897
2 94835 1 32899
2 94836 1 32899
2 94837 1 32910
2 94838 1 32910
2 94839 1 32923
2 94840 1 32923
2 94841 1 32930
2 94842 1 32930
2 94843 1 32933
2 94844 1 32933
2 94845 1 32996
2 94846 1 32996
2 94847 1 33006
2 94848 1 33006
2 94849 1 33046
2 94850 1 33046
2 94851 1 33046
2 94852 1 33046
2 94853 1 33053
2 94854 1 33053
2 94855 1 33070
2 94856 1 33070
2 94857 1 33070
2 94858 1 33070
2 94859 1 33071
2 94860 1 33071
2 94861 1 33131
2 94862 1 33131
2 94863 1 33316
2 94864 1 33316
2 94865 1 33316
2 94866 1 33317
2 94867 1 33317
2 94868 1 33317
2 94869 1 33338
2 94870 1 33338
2 94871 1 33344
2 94872 1 33344
2 94873 1 33344
2 94874 1 33344
2 94875 1 33344
2 94876 1 33371
2 94877 1 33371
2 94878 1 33371
2 94879 1 33371
2 94880 1 33371
2 94881 1 33371
2 94882 1 33371
2 94883 1 33391
2 94884 1 33391
2 94885 1 33432
2 94886 1 33432
2 94887 1 33457
2 94888 1 33457
2 94889 1 33475
2 94890 1 33475
2 94891 1 33482
2 94892 1 33482
2 94893 1 33485
2 94894 1 33485
2 94895 1 33491
2 94896 1 33491
2 94897 1 33495
2 94898 1 33495
2 94899 1 33495
2 94900 1 33498
2 94901 1 33498
2 94902 1 33498
2 94903 1 33505
2 94904 1 33505
2 94905 1 33512
2 94906 1 33512
2 94907 1 33512
2 94908 1 33528
2 94909 1 33528
2 94910 1 33530
2 94911 1 33530
2 94912 1 33530
2 94913 1 33530
2 94914 1 33530
2 94915 1 33530
2 94916 1 33542
2 94917 1 33542
2 94918 1 33543
2 94919 1 33543
2 94920 1 33543
2 94921 1 33543
2 94922 1 33552
2 94923 1 33552
2 94924 1 33561
2 94925 1 33561
2 94926 1 33568
2 94927 1 33568
2 94928 1 33568
2 94929 1 33584
2 94930 1 33584
2 94931 1 33593
2 94932 1 33593
2 94933 1 33593
2 94934 1 33593
2 94935 1 33593
2 94936 1 33594
2 94937 1 33594
2 94938 1 33594
2 94939 1 33594
2 94940 1 33596
2 94941 1 33596
2 94942 1 33598
2 94943 1 33598
2 94944 1 33607
2 94945 1 33607
2 94946 1 33607
2 94947 1 33622
2 94948 1 33622
2 94949 1 33632
2 94950 1 33632
2 94951 1 33640
2 94952 1 33640
2 94953 1 33641
2 94954 1 33641
2 94955 1 33641
2 94956 1 33644
2 94957 1 33644
2 94958 1 33672
2 94959 1 33672
2 94960 1 33677
2 94961 1 33677
2 94962 1 33679
2 94963 1 33679
2 94964 1 33679
2 94965 1 33683
2 94966 1 33683
2 94967 1 33684
2 94968 1 33684
2 94969 1 33707
2 94970 1 33707
2 94971 1 33724
2 94972 1 33724
2 94973 1 33724
2 94974 1 33757
2 94975 1 33757
2 94976 1 33757
2 94977 1 33758
2 94978 1 33758
2 94979 1 33761
2 94980 1 33761
2 94981 1 33762
2 94982 1 33762
2 94983 1 33767
2 94984 1 33767
2 94985 1 33803
2 94986 1 33803
2 94987 1 33803
2 94988 1 33804
2 94989 1 33804
2 94990 1 33806
2 94991 1 33806
2 94992 1 33806
2 94993 1 33835
2 94994 1 33835
2 94995 1 33839
2 94996 1 33839
2 94997 1 33839
2 94998 1 33839
2 94999 1 33866
2 95000 1 33866
2 95001 1 33869
2 95002 1 33869
2 95003 1 33869
2 95004 1 33870
2 95005 1 33870
2 95006 1 33897
2 95007 1 33897
2 95008 1 33905
2 95009 1 33905
2 95010 1 33921
2 95011 1 33921
2 95012 1 33960
2 95013 1 33960
2 95014 1 33961
2 95015 1 33961
2 95016 1 33987
2 95017 1 33987
2 95018 1 33987
2 95019 1 33987
2 95020 1 33992
2 95021 1 33992
2 95022 1 33992
2 95023 1 34003
2 95024 1 34003
2 95025 1 34011
2 95026 1 34011
2 95027 1 34011
2 95028 1 34011
2 95029 1 34032
2 95030 1 34032
2 95031 1 34036
2 95032 1 34036
2 95033 1 34042
2 95034 1 34042
2 95035 1 34048
2 95036 1 34048
2 95037 1 34049
2 95038 1 34049
2 95039 1 34058
2 95040 1 34058
2 95041 1 34071
2 95042 1 34071
2 95043 1 34197
2 95044 1 34197
2 95045 1 34199
2 95046 1 34199
2 95047 1 34202
2 95048 1 34202
2 95049 1 34207
2 95050 1 34207
2 95051 1 34211
2 95052 1 34211
2 95053 1 34263
2 95054 1 34263
2 95055 1 34263
2 95056 1 34292
2 95057 1 34292
2 95058 1 34296
2 95059 1 34296
2 95060 1 34300
2 95061 1 34300
2 95062 1 34317
2 95063 1 34317
2 95064 1 34318
2 95065 1 34318
2 95066 1 34318
2 95067 1 34377
2 95068 1 34377
2 95069 1 34391
2 95070 1 34391
2 95071 1 34414
2 95072 1 34414
2 95073 1 34415
2 95074 1 34415
2 95075 1 34449
2 95076 1 34449
2 95077 1 34466
2 95078 1 34466
2 95079 1 34469
2 95080 1 34469
2 95081 1 34475
2 95082 1 34475
2 95083 1 34510
2 95084 1 34510
2 95085 1 34521
2 95086 1 34521
2 95087 1 34546
2 95088 1 34546
2 95089 1 34546
2 95090 1 34546
2 95091 1 34546
2 95092 1 34546
2 95093 1 34546
2 95094 1 34547
2 95095 1 34547
2 95096 1 34547
2 95097 1 34567
2 95098 1 34567
2 95099 1 34581
2 95100 1 34581
2 95101 1 34618
2 95102 1 34618
2 95103 1 34618
2 95104 1 34618
2 95105 1 34646
2 95106 1 34646
2 95107 1 34646
2 95108 1 34648
2 95109 1 34648
2 95110 1 34650
2 95111 1 34650
2 95112 1 34680
2 95113 1 34680
2 95114 1 34680
2 95115 1 34693
2 95116 1 34693
2 95117 1 34704
2 95118 1 34704
2 95119 1 34704
2 95120 1 34720
2 95121 1 34720
2 95122 1 34722
2 95123 1 34722
2 95124 1 34778
2 95125 1 34778
2 95126 1 34793
2 95127 1 34793
2 95128 1 34795
2 95129 1 34795
2 95130 1 34795
2 95131 1 34795
2 95132 1 34831
2 95133 1 34831
2 95134 1 34831
2 95135 1 34841
2 95136 1 34841
2 95137 1 34879
2 95138 1 34879
2 95139 1 34896
2 95140 1 34896
2 95141 1 34934
2 95142 1 34934
2 95143 1 34934
2 95144 1 34934
2 95145 1 34934
2 95146 1 34972
2 95147 1 34972
2 95148 1 34972
2 95149 1 35001
2 95150 1 35001
2 95151 1 35003
2 95152 1 35003
2 95153 1 35029
2 95154 1 35029
2 95155 1 35030
2 95156 1 35030
2 95157 1 35030
2 95158 1 35030
2 95159 1 35030
2 95160 1 35068
2 95161 1 35068
2 95162 1 35068
2 95163 1 35073
2 95164 1 35073
2 95165 1 35076
2 95166 1 35076
2 95167 1 35084
2 95168 1 35084
2 95169 1 35098
2 95170 1 35098
2 95171 1 35110
2 95172 1 35110
2 95173 1 35112
2 95174 1 35112
2 95175 1 35116
2 95176 1 35116
2 95177 1 35123
2 95178 1 35123
2 95179 1 35126
2 95180 1 35126
2 95181 1 35126
2 95182 1 35126
2 95183 1 35131
2 95184 1 35131
2 95185 1 35131
2 95186 1 35132
2 95187 1 35132
2 95188 1 35187
2 95189 1 35187
2 95190 1 35193
2 95191 1 35193
2 95192 1 35242
2 95193 1 35242
2 95194 1 35242
2 95195 1 35242
2 95196 1 35242
2 95197 1 35253
2 95198 1 35253
2 95199 1 35263
2 95200 1 35263
2 95201 1 35290
2 95202 1 35290
2 95203 1 35294
2 95204 1 35294
2 95205 1 35327
2 95206 1 35327
2 95207 1 35327
2 95208 1 35334
2 95209 1 35334
2 95210 1 35374
2 95211 1 35374
2 95212 1 35468
2 95213 1 35468
2 95214 1 35468
2 95215 1 35493
2 95216 1 35493
2 95217 1 35500
2 95218 1 35500
2 95219 1 35529
2 95220 1 35529
2 95221 1 35540
2 95222 1 35540
2 95223 1 35575
2 95224 1 35575
2 95225 1 35575
2 95226 1 35575
2 95227 1 35577
2 95228 1 35577
2 95229 1 35577
2 95230 1 35577
2 95231 1 35577
2 95232 1 35577
2 95233 1 35585
2 95234 1 35585
2 95235 1 35606
2 95236 1 35606
2 95237 1 35606
2 95238 1 35609
2 95239 1 35609
2 95240 1 35616
2 95241 1 35616
2 95242 1 35622
2 95243 1 35622
2 95244 1 35622
2 95245 1 35622
2 95246 1 35623
2 95247 1 35623
2 95248 1 35623
2 95249 1 35643
2 95250 1 35643
2 95251 1 35643
2 95252 1 35643
2 95253 1 35643
2 95254 1 35643
2 95255 1 35643
2 95256 1 35644
2 95257 1 35644
2 95258 1 35645
2 95259 1 35645
2 95260 1 35645
2 95261 1 35645
2 95262 1 35645
2 95263 1 35645
2 95264 1 35645
2 95265 1 35662
2 95266 1 35662
2 95267 1 35664
2 95268 1 35664
2 95269 1 35665
2 95270 1 35665
2 95271 1 35730
2 95272 1 35730
2 95273 1 35738
2 95274 1 35738
2 95275 1 35738
2 95276 1 35775
2 95277 1 35775
2 95278 1 35809
2 95279 1 35809
2 95280 1 35818
2 95281 1 35818
2 95282 1 35819
2 95283 1 35819
2 95284 1 35834
2 95285 1 35834
2 95286 1 35883
2 95287 1 35883
2 95288 1 35883
2 95289 1 35883
2 95290 1 35883
2 95291 1 35883
2 95292 1 35883
2 95293 1 35883
2 95294 1 35883
2 95295 1 35883
2 95296 1 35883
2 95297 1 35883
2 95298 1 35883
2 95299 1 35883
2 95300 1 35883
2 95301 1 35883
2 95302 1 35883
2 95303 1 35883
2 95304 1 35883
2 95305 1 35883
2 95306 1 35883
2 95307 1 35883
2 95308 1 35883
2 95309 1 35883
2 95310 1 35883
2 95311 1 35883
2 95312 1 35883
2 95313 1 35883
2 95314 1 35883
2 95315 1 35883
2 95316 1 35883
2 95317 1 35883
2 95318 1 35883
2 95319 1 35883
2 95320 1 35883
2 95321 1 35883
2 95322 1 35883
2 95323 1 35883
2 95324 1 35883
2 95325 1 35883
2 95326 1 35883
2 95327 1 35883
2 95328 1 35885
2 95329 1 35885
2 95330 1 35888
2 95331 1 35888
2 95332 1 35888
2 95333 1 35888
2 95334 1 35889
2 95335 1 35889
2 95336 1 35889
2 95337 1 35892
2 95338 1 35892
2 95339 1 35892
2 95340 1 35910
2 95341 1 35910
2 95342 1 35911
2 95343 1 35911
2 95344 1 35912
2 95345 1 35912
2 95346 1 35918
2 95347 1 35918
2 95348 1 35918
2 95349 1 35921
2 95350 1 35921
2 95351 1 35934
2 95352 1 35934
2 95353 1 35962
2 95354 1 35962
2 95355 1 35966
2 95356 1 35966
2 95357 1 35970
2 95358 1 35970
2 95359 1 35986
2 95360 1 35986
2 95361 1 35999
2 95362 1 35999
2 95363 1 36026
2 95364 1 36026
2 95365 1 36035
2 95366 1 36035
2 95367 1 36064
2 95368 1 36064
2 95369 1 36067
2 95370 1 36067
2 95371 1 36116
2 95372 1 36116
2 95373 1 36149
2 95374 1 36149
2 95375 1 36162
2 95376 1 36162
2 95377 1 36172
2 95378 1 36172
2 95379 1 36176
2 95380 1 36176
2 95381 1 36222
2 95382 1 36222
2 95383 1 36224
2 95384 1 36224
2 95385 1 36253
2 95386 1 36253
2 95387 1 36258
2 95388 1 36258
2 95389 1 36281
2 95390 1 36281
2 95391 1 36334
2 95392 1 36334
2 95393 1 36334
2 95394 1 36342
2 95395 1 36342
2 95396 1 36348
2 95397 1 36348
2 95398 1 36351
2 95399 1 36351
2 95400 1 36367
2 95401 1 36367
2 95402 1 36369
2 95403 1 36369
2 95404 1 36377
2 95405 1 36377
2 95406 1 36380
2 95407 1 36380
2 95408 1 36382
2 95409 1 36382
2 95410 1 36382
2 95411 1 36407
2 95412 1 36407
2 95413 1 36420
2 95414 1 36420
2 95415 1 36423
2 95416 1 36423
2 95417 1 36423
2 95418 1 36465
2 95419 1 36465
2 95420 1 36465
2 95421 1 36467
2 95422 1 36467
2 95423 1 36469
2 95424 1 36469
2 95425 1 36485
2 95426 1 36485
2 95427 1 36501
2 95428 1 36501
2 95429 1 36501
2 95430 1 36520
2 95431 1 36520
2 95432 1 36522
2 95433 1 36522
2 95434 1 36522
2 95435 1 36525
2 95436 1 36525
2 95437 1 36526
2 95438 1 36526
2 95439 1 36544
2 95440 1 36544
2 95441 1 36547
2 95442 1 36547
2 95443 1 36547
2 95444 1 36547
2 95445 1 36548
2 95446 1 36548
2 95447 1 36551
2 95448 1 36551
2 95449 1 36627
2 95450 1 36627
2 95451 1 36649
2 95452 1 36649
2 95453 1 36650
2 95454 1 36650
2 95455 1 36656
2 95456 1 36656
2 95457 1 36657
2 95458 1 36657
2 95459 1 36658
2 95460 1 36658
2 95461 1 36670
2 95462 1 36670
2 95463 1 36672
2 95464 1 36672
2 95465 1 36681
2 95466 1 36681
2 95467 1 36739
2 95468 1 36739
2 95469 1 36739
2 95470 1 36739
2 95471 1 36739
2 95472 1 36739
2 95473 1 36739
2 95474 1 36739
2 95475 1 36739
2 95476 1 36739
2 95477 1 36739
2 95478 1 36739
2 95479 1 36739
2 95480 1 36739
2 95481 1 36740
2 95482 1 36740
2 95483 1 36741
2 95484 1 36741
2 95485 1 36742
2 95486 1 36742
2 95487 1 36771
2 95488 1 36771
2 95489 1 36771
2 95490 1 36771
2 95491 1 36771
2 95492 1 36800
2 95493 1 36800
2 95494 1 36800
2 95495 1 36800
2 95496 1 36841
2 95497 1 36841
2 95498 1 36841
2 95499 1 36842
2 95500 1 36842
2 95501 1 36844
2 95502 1 36844
2 95503 1 36845
2 95504 1 36845
2 95505 1 36846
2 95506 1 36846
2 95507 1 36846
2 95508 1 36867
2 95509 1 36867
2 95510 1 36878
2 95511 1 36878
2 95512 1 36878
2 95513 1 36878
2 95514 1 36883
2 95515 1 36883
2 95516 1 36900
2 95517 1 36900
2 95518 1 36910
2 95519 1 36910
2 95520 1 36911
2 95521 1 36911
2 95522 1 36966
2 95523 1 36966
2 95524 1 36967
2 95525 1 36967
2 95526 1 36968
2 95527 1 36968
2 95528 1 36970
2 95529 1 36970
2 95530 1 36978
2 95531 1 36978
2 95532 1 36981
2 95533 1 36981
2 95534 1 36986
2 95535 1 36986
2 95536 1 36993
2 95537 1 36993
2 95538 1 36993
2 95539 1 36994
2 95540 1 36994
2 95541 1 36994
2 95542 1 36994
2 95543 1 37033
2 95544 1 37033
2 95545 1 37034
2 95546 1 37034
2 95547 1 37065
2 95548 1 37065
2 95549 1 37072
2 95550 1 37072
2 95551 1 37105
2 95552 1 37105
2 95553 1 37105
2 95554 1 37106
2 95555 1 37106
2 95556 1 37107
2 95557 1 37107
2 95558 1 37116
2 95559 1 37116
2 95560 1 37117
2 95561 1 37117
2 95562 1 37119
2 95563 1 37119
2 95564 1 37149
2 95565 1 37149
2 95566 1 37172
2 95567 1 37172
2 95568 1 37172
2 95569 1 37186
2 95570 1 37186
2 95571 1 37189
2 95572 1 37189
2 95573 1 37196
2 95574 1 37196
2 95575 1 37212
2 95576 1 37212
2 95577 1 37229
2 95578 1 37229
2 95579 1 37232
2 95580 1 37232
2 95581 1 37240
2 95582 1 37240
2 95583 1 37241
2 95584 1 37241
2 95585 1 37285
2 95586 1 37285
2 95587 1 37290
2 95588 1 37290
2 95589 1 37293
2 95590 1 37293
2 95591 1 37299
2 95592 1 37299
2 95593 1 37310
2 95594 1 37310
2 95595 1 37324
2 95596 1 37324
2 95597 1 37324
2 95598 1 37324
2 95599 1 37325
2 95600 1 37325
2 95601 1 37325
2 95602 1 37325
2 95603 1 37362
2 95604 1 37362
2 95605 1 37385
2 95606 1 37385
2 95607 1 37448
2 95608 1 37448
2 95609 1 37453
2 95610 1 37453
2 95611 1 37506
2 95612 1 37506
2 95613 1 37511
2 95614 1 37511
2 95615 1 37522
2 95616 1 37522
2 95617 1 37526
2 95618 1 37526
2 95619 1 37534
2 95620 1 37534
2 95621 1 37534
2 95622 1 37556
2 95623 1 37556
2 95624 1 37556
2 95625 1 37579
2 95626 1 37579
2 95627 1 37590
2 95628 1 37590
2 95629 1 37641
2 95630 1 37641
2 95631 1 37697
2 95632 1 37697
2 95633 1 37697
2 95634 1 37697
2 95635 1 37697
2 95636 1 37697
2 95637 1 37697
2 95638 1 37697
2 95639 1 37697
2 95640 1 37697
2 95641 1 37697
2 95642 1 37697
2 95643 1 37704
2 95644 1 37704
2 95645 1 37705
2 95646 1 37705
2 95647 1 37705
2 95648 1 37705
2 95649 1 37735
2 95650 1 37735
2 95651 1 37735
2 95652 1 37761
2 95653 1 37761
2 95654 1 37764
2 95655 1 37764
2 95656 1 37768
2 95657 1 37768
2 95658 1 37772
2 95659 1 37772
2 95660 1 37786
2 95661 1 37786
2 95662 1 37786
2 95663 1 37786
2 95664 1 37786
2 95665 1 37820
2 95666 1 37820
2 95667 1 37840
2 95668 1 37840
2 95669 1 37841
2 95670 1 37841
2 95671 1 37852
2 95672 1 37852
2 95673 1 37874
2 95674 1 37874
2 95675 1 37898
2 95676 1 37898
2 95677 1 37902
2 95678 1 37902
2 95679 1 37912
2 95680 1 37912
2 95681 1 37944
2 95682 1 37944
2 95683 1 37987
2 95684 1 37987
2 95685 1 38012
2 95686 1 38012
2 95687 1 38024
2 95688 1 38024
2 95689 1 38069
2 95690 1 38069
2 95691 1 38139
2 95692 1 38139
2 95693 1 38146
2 95694 1 38146
2 95695 1 38179
2 95696 1 38179
2 95697 1 38179
2 95698 1 38184
2 95699 1 38184
2 95700 1 38184
2 95701 1 38185
2 95702 1 38185
2 95703 1 38185
2 95704 1 38194
2 95705 1 38194
2 95706 1 38194
2 95707 1 38194
2 95708 1 38194
2 95709 1 38194
2 95710 1 38194
2 95711 1 38195
2 95712 1 38195
2 95713 1 38196
2 95714 1 38196
2 95715 1 38196
2 95716 1 38196
2 95717 1 38196
2 95718 1 38196
2 95719 1 38196
2 95720 1 38196
2 95721 1 38196
2 95722 1 38196
2 95723 1 38198
2 95724 1 38198
2 95725 1 38268
2 95726 1 38268
2 95727 1 38268
2 95728 1 38268
2 95729 1 38298
2 95730 1 38298
2 95731 1 38299
2 95732 1 38299
2 95733 1 38299
2 95734 1 38319
2 95735 1 38319
2 95736 1 38319
2 95737 1 38323
2 95738 1 38323
2 95739 1 38325
2 95740 1 38325
2 95741 1 38332
2 95742 1 38332
2 95743 1 38332
2 95744 1 38332
2 95745 1 38332
2 95746 1 38332
2 95747 1 38335
2 95748 1 38335
2 95749 1 38335
2 95750 1 38336
2 95751 1 38336
2 95752 1 38358
2 95753 1 38358
2 95754 1 38361
2 95755 1 38361
2 95756 1 38412
2 95757 1 38412
2 95758 1 38459
2 95759 1 38459
2 95760 1 38485
2 95761 1 38485
2 95762 1 38543
2 95763 1 38543
2 95764 1 38545
2 95765 1 38545
2 95766 1 38561
2 95767 1 38561
2 95768 1 38572
2 95769 1 38572
2 95770 1 38577
2 95771 1 38577
2 95772 1 38614
2 95773 1 38614
2 95774 1 38615
2 95775 1 38615
2 95776 1 38632
2 95777 1 38632
2 95778 1 38640
2 95779 1 38640
2 95780 1 38640
2 95781 1 38688
2 95782 1 38688
2 95783 1 38689
2 95784 1 38689
2 95785 1 38707
2 95786 1 38707
2 95787 1 38734
2 95788 1 38734
2 95789 1 38738
2 95790 1 38738
2 95791 1 38740
2 95792 1 38740
2 95793 1 38740
2 95794 1 38762
2 95795 1 38762
2 95796 1 38780
2 95797 1 38780
2 95798 1 38780
2 95799 1 38804
2 95800 1 38804
2 95801 1 38820
2 95802 1 38820
2 95803 1 38828
2 95804 1 38828
2 95805 1 38828
2 95806 1 38828
2 95807 1 38828
2 95808 1 38845
2 95809 1 38845
2 95810 1 38853
2 95811 1 38853
2 95812 1 38853
2 95813 1 38853
2 95814 1 38853
2 95815 1 38853
2 95816 1 38868
2 95817 1 38868
2 95818 1 38893
2 95819 1 38893
2 95820 1 38893
2 95821 1 38895
2 95822 1 38895
2 95823 1 38961
2 95824 1 38961
2 95825 1 38967
2 95826 1 38967
2 95827 1 38967
2 95828 1 38967
2 95829 1 38986
2 95830 1 38986
2 95831 1 39002
2 95832 1 39002
2 95833 1 39003
2 95834 1 39003
2 95835 1 39003
2 95836 1 39003
2 95837 1 39003
2 95838 1 39018
2 95839 1 39018
2 95840 1 39018
2 95841 1 39020
2 95842 1 39020
2 95843 1 39048
2 95844 1 39048
2 95845 1 39051
2 95846 1 39051
2 95847 1 39089
2 95848 1 39089
2 95849 1 39097
2 95850 1 39097
2 95851 1 39135
2 95852 1 39135
2 95853 1 39135
2 95854 1 39135
2 95855 1 39152
2 95856 1 39152
2 95857 1 39172
2 95858 1 39172
2 95859 1 39189
2 95860 1 39189
2 95861 1 39189
2 95862 1 39194
2 95863 1 39194
2 95864 1 39202
2 95865 1 39202
2 95866 1 39214
2 95867 1 39214
2 95868 1 39228
2 95869 1 39228
2 95870 1 39228
2 95871 1 39228
2 95872 1 39228
2 95873 1 39235
2 95874 1 39235
2 95875 1 39235
2 95876 1 39236
2 95877 1 39236
2 95878 1 39243
2 95879 1 39243
2 95880 1 39244
2 95881 1 39244
2 95882 1 39244
2 95883 1 39246
2 95884 1 39246
2 95885 1 39259
2 95886 1 39259
2 95887 1 39260
2 95888 1 39260
2 95889 1 39303
2 95890 1 39303
2 95891 1 39331
2 95892 1 39331
2 95893 1 39336
2 95894 1 39336
2 95895 1 39355
2 95896 1 39355
2 95897 1 39364
2 95898 1 39364
2 95899 1 39373
2 95900 1 39373
2 95901 1 39380
2 95902 1 39380
2 95903 1 39399
2 95904 1 39399
2 95905 1 39409
2 95906 1 39409
2 95907 1 39409
2 95908 1 39411
2 95909 1 39411
2 95910 1 39411
2 95911 1 39415
2 95912 1 39415
2 95913 1 39459
2 95914 1 39459
2 95915 1 39459
2 95916 1 39459
2 95917 1 39459
2 95918 1 39459
2 95919 1 39460
2 95920 1 39460
2 95921 1 39480
2 95922 1 39480
2 95923 1 39480
2 95924 1 39481
2 95925 1 39481
2 95926 1 39481
2 95927 1 39484
2 95928 1 39484
2 95929 1 39511
2 95930 1 39511
2 95931 1 39512
2 95932 1 39512
2 95933 1 39512
2 95934 1 39512
2 95935 1 39532
2 95936 1 39532
2 95937 1 39540
2 95938 1 39540
2 95939 1 39540
2 95940 1 39546
2 95941 1 39546
2 95942 1 39546
2 95943 1 39553
2 95944 1 39553
2 95945 1 39557
2 95946 1 39557
2 95947 1 39557
2 95948 1 39567
2 95949 1 39567
2 95950 1 39570
2 95951 1 39570
2 95952 1 39570
2 95953 1 39570
2 95954 1 39572
2 95955 1 39572
2 95956 1 39576
2 95957 1 39576
2 95958 1 39576
2 95959 1 39590
2 95960 1 39590
2 95961 1 39590
2 95962 1 39590
2 95963 1 39601
2 95964 1 39601
2 95965 1 39609
2 95966 1 39609
2 95967 1 39610
2 95968 1 39610
2 95969 1 39610
2 95970 1 39610
2 95971 1 39612
2 95972 1 39612
2 95973 1 39617
2 95974 1 39617
2 95975 1 39617
2 95976 1 39617
2 95977 1 39617
2 95978 1 39617
2 95979 1 39620
2 95980 1 39620
2 95981 1 39620
2 95982 1 39641
2 95983 1 39641
2 95984 1 39642
2 95985 1 39642
2 95986 1 39642
2 95987 1 39644
2 95988 1 39644
2 95989 1 39644
2 95990 1 39644
2 95991 1 39645
2 95992 1 39645
2 95993 1 39659
2 95994 1 39659
2 95995 1 39685
2 95996 1 39685
2 95997 1 39685
2 95998 1 39686
2 95999 1 39686
2 96000 1 39690
2 96001 1 39690
2 96002 1 39697
2 96003 1 39697
2 96004 1 39708
2 96005 1 39708
2 96006 1 39712
2 96007 1 39712
2 96008 1 39712
2 96009 1 39715
2 96010 1 39715
2 96011 1 39715
2 96012 1 39715
2 96013 1 39723
2 96014 1 39723
2 96015 1 39727
2 96016 1 39727
2 96017 1 39727
2 96018 1 39727
2 96019 1 39727
2 96020 1 39727
2 96021 1 39727
2 96022 1 39727
2 96023 1 39727
2 96024 1 39728
2 96025 1 39728
2 96026 1 39728
2 96027 1 39729
2 96028 1 39729
2 96029 1 39739
2 96030 1 39739
2 96031 1 39756
2 96032 1 39756
2 96033 1 39756
2 96034 1 39759
2 96035 1 39759
2 96036 1 39760
2 96037 1 39760
2 96038 1 39786
2 96039 1 39786
2 96040 1 39806
2 96041 1 39806
2 96042 1 39814
2 96043 1 39814
2 96044 1 39822
2 96045 1 39822
2 96046 1 39822
2 96047 1 39835
2 96048 1 39835
2 96049 1 39845
2 96050 1 39845
2 96051 1 39846
2 96052 1 39846
2 96053 1 39846
2 96054 1 39846
2 96055 1 39848
2 96056 1 39848
2 96057 1 39855
2 96058 1 39855
2 96059 1 39864
2 96060 1 39864
2 96061 1 39873
2 96062 1 39873
2 96063 1 39875
2 96064 1 39875
2 96065 1 39875
2 96066 1 39875
2 96067 1 39875
2 96068 1 39875
2 96069 1 39875
2 96070 1 39876
2 96071 1 39876
2 96072 1 39876
2 96073 1 39878
2 96074 1 39878
2 96075 1 39886
2 96076 1 39886
2 96077 1 39888
2 96078 1 39888
2 96079 1 39893
2 96080 1 39893
2 96081 1 39893
2 96082 1 39893
2 96083 1 39893
2 96084 1 39902
2 96085 1 39902
2 96086 1 39921
2 96087 1 39921
2 96088 1 39921
2 96089 1 39921
2 96090 1 39933
2 96091 1 39933
2 96092 1 39933
2 96093 1 39933
2 96094 1 39942
2 96095 1 39942
2 96096 1 39942
2 96097 1 39956
2 96098 1 39956
2 96099 1 39986
2 96100 1 39986
2 96101 1 39997
2 96102 1 39997
2 96103 1 39998
2 96104 1 39998
2 96105 1 40014
2 96106 1 40014
2 96107 1 40021
2 96108 1 40021
2 96109 1 40021
2 96110 1 40034
2 96111 1 40034
2 96112 1 40064
2 96113 1 40064
2 96114 1 40072
2 96115 1 40072
2 96116 1 40072
2 96117 1 40073
2 96118 1 40073
2 96119 1 40103
2 96120 1 40103
2 96121 1 40103
2 96122 1 40103
2 96123 1 40103
2 96124 1 40104
2 96125 1 40104
2 96126 1 40104
2 96127 1 40104
2 96128 1 40108
2 96129 1 40108
2 96130 1 40124
2 96131 1 40124
2 96132 1 40124
2 96133 1 40125
2 96134 1 40125
2 96135 1 40133
2 96136 1 40133
2 96137 1 40148
2 96138 1 40148
2 96139 1 40148
2 96140 1 40149
2 96141 1 40149
2 96142 1 40160
2 96143 1 40160
2 96144 1 40161
2 96145 1 40161
2 96146 1 40161
2 96147 1 40198
2 96148 1 40198
2 96149 1 40223
2 96150 1 40223
2 96151 1 40243
2 96152 1 40243
2 96153 1 40243
2 96154 1 40246
2 96155 1 40246
2 96156 1 40246
2 96157 1 40254
2 96158 1 40254
2 96159 1 40261
2 96160 1 40261
2 96161 1 40261
2 96162 1 40263
2 96163 1 40263
2 96164 1 40272
2 96165 1 40272
2 96166 1 40274
2 96167 1 40274
2 96168 1 40274
2 96169 1 40283
2 96170 1 40283
2 96171 1 40283
2 96172 1 40286
2 96173 1 40286
2 96174 1 40286
2 96175 1 40286
2 96176 1 40286
2 96177 1 40286
2 96178 1 40286
2 96179 1 40296
2 96180 1 40296
2 96181 1 40296
2 96182 1 40296
2 96183 1 40303
2 96184 1 40303
2 96185 1 40312
2 96186 1 40312
2 96187 1 40312
2 96188 1 40312
2 96189 1 40312
2 96190 1 40312
2 96191 1 40312
2 96192 1 40338
2 96193 1 40338
2 96194 1 40339
2 96195 1 40339
2 96196 1 40339
2 96197 1 40339
2 96198 1 40357
2 96199 1 40357
2 96200 1 40357
2 96201 1 40379
2 96202 1 40379
2 96203 1 40379
2 96204 1 40379
2 96205 1 40397
2 96206 1 40397
2 96207 1 40397
2 96208 1 40416
2 96209 1 40416
2 96210 1 40419
2 96211 1 40419
2 96212 1 40423
2 96213 1 40423
2 96214 1 40423
2 96215 1 40441
2 96216 1 40441
2 96217 1 40445
2 96218 1 40445
2 96219 1 40445
2 96220 1 40445
2 96221 1 40464
2 96222 1 40464
2 96223 1 40465
2 96224 1 40465
2 96225 1 40510
2 96226 1 40510
2 96227 1 40544
2 96228 1 40544
2 96229 1 40556
2 96230 1 40556
2 96231 1 40556
2 96232 1 40556
2 96233 1 40564
2 96234 1 40564
2 96235 1 40572
2 96236 1 40572
2 96237 1 40572
2 96238 1 40572
2 96239 1 40572
2 96240 1 40596
2 96241 1 40596
2 96242 1 40596
2 96243 1 40596
2 96244 1 40596
2 96245 1 40596
2 96246 1 40596
2 96247 1 40596
2 96248 1 40598
2 96249 1 40598
2 96250 1 40598
2 96251 1 40607
2 96252 1 40607
2 96253 1 40608
2 96254 1 40608
2 96255 1 40608
2 96256 1 40614
2 96257 1 40614
2 96258 1 40628
2 96259 1 40628
2 96260 1 40630
2 96261 1 40630
2 96262 1 40666
2 96263 1 40666
2 96264 1 40666
2 96265 1 40666
2 96266 1 40667
2 96267 1 40667
2 96268 1 40667
2 96269 1 40667
2 96270 1 40667
2 96271 1 40667
2 96272 1 40677
2 96273 1 40677
2 96274 1 40702
2 96275 1 40702
2 96276 1 40707
2 96277 1 40707
2 96278 1 40754
2 96279 1 40754
2 96280 1 40754
2 96281 1 40756
2 96282 1 40756
2 96283 1 40756
2 96284 1 40756
2 96285 1 40766
2 96286 1 40766
2 96287 1 40793
2 96288 1 40793
2 96289 1 40794
2 96290 1 40794
2 96291 1 40816
2 96292 1 40816
2 96293 1 40816
2 96294 1 40816
2 96295 1 40816
2 96296 1 40817
2 96297 1 40817
2 96298 1 40831
2 96299 1 40831
2 96300 1 40831
2 96301 1 40835
2 96302 1 40835
2 96303 1 40849
2 96304 1 40849
2 96305 1 40850
2 96306 1 40850
2 96307 1 40859
2 96308 1 40859
2 96309 1 40877
2 96310 1 40877
2 96311 1 40877
2 96312 1 40877
2 96313 1 40877
2 96314 1 40877
2 96315 1 40877
2 96316 1 40887
2 96317 1 40887
2 96318 1 40901
2 96319 1 40901
2 96320 1 40902
2 96321 1 40902
2 96322 1 40923
2 96323 1 40923
2 96324 1 40923
2 96325 1 40923
2 96326 1 40923
2 96327 1 40923
2 96328 1 40923
2 96329 1 40923
2 96330 1 40923
2 96331 1 40923
2 96332 1 40923
2 96333 1 40923
2 96334 1 40923
2 96335 1 40923
2 96336 1 40923
2 96337 1 40923
2 96338 1 40925
2 96339 1 40925
2 96340 1 40943
2 96341 1 40943
2 96342 1 40953
2 96343 1 40953
2 96344 1 40977
2 96345 1 40977
2 96346 1 40982
2 96347 1 40982
2 96348 1 40982
2 96349 1 41032
2 96350 1 41032
2 96351 1 41042
2 96352 1 41042
2 96353 1 41072
2 96354 1 41072
2 96355 1 41073
2 96356 1 41073
2 96357 1 41112
2 96358 1 41112
2 96359 1 41118
2 96360 1 41118
2 96361 1 41119
2 96362 1 41119
2 96363 1 41121
2 96364 1 41121
2 96365 1 41134
2 96366 1 41134
2 96367 1 41153
2 96368 1 41153
2 96369 1 41156
2 96370 1 41156
2 96371 1 41157
2 96372 1 41157
2 96373 1 41158
2 96374 1 41158
2 96375 1 41160
2 96376 1 41160
2 96377 1 41175
2 96378 1 41175
2 96379 1 41187
2 96380 1 41187
2 96381 1 41192
2 96382 1 41192
2 96383 1 41192
2 96384 1 41204
2 96385 1 41204
2 96386 1 41204
2 96387 1 41205
2 96388 1 41205
2 96389 1 41205
2 96390 1 41206
2 96391 1 41206
2 96392 1 41207
2 96393 1 41207
2 96394 1 41207
2 96395 1 41220
2 96396 1 41220
2 96397 1 41223
2 96398 1 41223
2 96399 1 41227
2 96400 1 41227
2 96401 1 41244
2 96402 1 41244
2 96403 1 41248
2 96404 1 41248
2 96405 1 41261
2 96406 1 41261
2 96407 1 41268
2 96408 1 41268
2 96409 1 41272
2 96410 1 41272
2 96411 1 41292
2 96412 1 41292
2 96413 1 41303
2 96414 1 41303
2 96415 1 41303
2 96416 1 41303
2 96417 1 41318
2 96418 1 41318
2 96419 1 41321
2 96420 1 41321
2 96421 1 41321
2 96422 1 41321
2 96423 1 41321
2 96424 1 41354
2 96425 1 41354
2 96426 1 41363
2 96427 1 41363
2 96428 1 41380
2 96429 1 41380
2 96430 1 41387
2 96431 1 41387
2 96432 1 41391
2 96433 1 41391
2 96434 1 41434
2 96435 1 41434
2 96436 1 41434
2 96437 1 41434
2 96438 1 41434
2 96439 1 41435
2 96440 1 41435
2 96441 1 41435
2 96442 1 41439
2 96443 1 41439
2 96444 1 41439
2 96445 1 41439
2 96446 1 41439
2 96447 1 41460
2 96448 1 41460
2 96449 1 41475
2 96450 1 41475
2 96451 1 41480
2 96452 1 41480
2 96453 1 41487
2 96454 1 41487
2 96455 1 41489
2 96456 1 41489
2 96457 1 41496
2 96458 1 41496
2 96459 1 41497
2 96460 1 41497
2 96461 1 41506
2 96462 1 41506
2 96463 1 41507
2 96464 1 41507
2 96465 1 41512
2 96466 1 41512
2 96467 1 41513
2 96468 1 41513
2 96469 1 41513
2 96470 1 41513
2 96471 1 41513
2 96472 1 41531
2 96473 1 41531
2 96474 1 41539
2 96475 1 41539
2 96476 1 41597
2 96477 1 41597
2 96478 1 41612
2 96479 1 41612
2 96480 1 41635
2 96481 1 41635
2 96482 1 41675
2 96483 1 41675
2 96484 1 41675
2 96485 1 41675
2 96486 1 41686
2 96487 1 41686
2 96488 1 41686
2 96489 1 41686
2 96490 1 41686
2 96491 1 41686
2 96492 1 41686
2 96493 1 41686
2 96494 1 41686
2 96495 1 41687
2 96496 1 41687
2 96497 1 41687
2 96498 1 41734
2 96499 1 41734
2 96500 1 41734
2 96501 1 41734
2 96502 1 41735
2 96503 1 41735
2 96504 1 41735
2 96505 1 41736
2 96506 1 41736
2 96507 1 41784
2 96508 1 41784
2 96509 1 41784
2 96510 1 41784
2 96511 1 41784
2 96512 1 41806
2 96513 1 41806
2 96514 1 41807
2 96515 1 41807
2 96516 1 41807
2 96517 1 41826
2 96518 1 41826
2 96519 1 41826
2 96520 1 41826
2 96521 1 41826
2 96522 1 41844
2 96523 1 41844
2 96524 1 41844
2 96525 1 41852
2 96526 1 41852
2 96527 1 41852
2 96528 1 41853
2 96529 1 41853
2 96530 1 41856
2 96531 1 41856
2 96532 1 41856
2 96533 1 41856
2 96534 1 41856
2 96535 1 41856
2 96536 1 41856
2 96537 1 41860
2 96538 1 41860
2 96539 1 41873
2 96540 1 41873
2 96541 1 41873
2 96542 1 41880
2 96543 1 41880
2 96544 1 41913
2 96545 1 41913
2 96546 1 41919
2 96547 1 41919
2 96548 1 41920
2 96549 1 41920
2 96550 1 41929
2 96551 1 41929
2 96552 1 41934
2 96553 1 41934
2 96554 1 41934
2 96555 1 41934
2 96556 1 41934
2 96557 1 41934
2 96558 1 41947
2 96559 1 41947
2 96560 1 41957
2 96561 1 41957
2 96562 1 41960
2 96563 1 41960
2 96564 1 41981
2 96565 1 41981
2 96566 1 41981
2 96567 1 41982
2 96568 1 41982
2 96569 1 41982
2 96570 1 41989
2 96571 1 41989
2 96572 1 41989
2 96573 1 41989
2 96574 1 41989
2 96575 1 41989
2 96576 1 41990
2 96577 1 41990
2 96578 1 41990
2 96579 1 41997
2 96580 1 41997
2 96581 1 41997
2 96582 1 42018
2 96583 1 42018
2 96584 1 42018
2 96585 1 42018
2 96586 1 42028
2 96587 1 42028
2 96588 1 42028
2 96589 1 42028
2 96590 1 42035
2 96591 1 42035
2 96592 1 42050
2 96593 1 42050
2 96594 1 42058
2 96595 1 42058
2 96596 1 42078
2 96597 1 42078
2 96598 1 42090
2 96599 1 42090
2 96600 1 42090
2 96601 1 42090
2 96602 1 42090
2 96603 1 42091
2 96604 1 42091
2 96605 1 42108
2 96606 1 42108
2 96607 1 42109
2 96608 1 42109
2 96609 1 42109
2 96610 1 42109
2 96611 1 42118
2 96612 1 42118
2 96613 1 42121
2 96614 1 42121
2 96615 1 42124
2 96616 1 42124
2 96617 1 42124
2 96618 1 42163
2 96619 1 42163
2 96620 1 42163
2 96621 1 42163
2 96622 1 42179
2 96623 1 42179
2 96624 1 42188
2 96625 1 42188
2 96626 1 42232
2 96627 1 42232
2 96628 1 42232
2 96629 1 42241
2 96630 1 42241
2 96631 1 42243
2 96632 1 42243
2 96633 1 42252
2 96634 1 42252
2 96635 1 42258
2 96636 1 42258
2 96637 1 42261
2 96638 1 42261
2 96639 1 42261
2 96640 1 42261
2 96641 1 42268
2 96642 1 42268
2 96643 1 42275
2 96644 1 42275
2 96645 1 42283
2 96646 1 42283
2 96647 1 42287
2 96648 1 42287
2 96649 1 42295
2 96650 1 42295
2 96651 1 42295
2 96652 1 42312
2 96653 1 42312
2 96654 1 42325
2 96655 1 42325
2 96656 1 42329
2 96657 1 42329
2 96658 1 42333
2 96659 1 42333
2 96660 1 42338
2 96661 1 42338
2 96662 1 42376
2 96663 1 42376
2 96664 1 42389
2 96665 1 42389
2 96666 1 42389
2 96667 1 42389
2 96668 1 42398
2 96669 1 42398
2 96670 1 42398
2 96671 1 42398
2 96672 1 42398
2 96673 1 42398
2 96674 1 42399
2 96675 1 42399
2 96676 1 42410
2 96677 1 42410
2 96678 1 42410
2 96679 1 42410
2 96680 1 42410
2 96681 1 42410
2 96682 1 42411
2 96683 1 42411
2 96684 1 42430
2 96685 1 42430
2 96686 1 42431
2 96687 1 42431
2 96688 1 42431
2 96689 1 42431
2 96690 1 42431
2 96691 1 42433
2 96692 1 42433
2 96693 1 42434
2 96694 1 42434
2 96695 1 42480
2 96696 1 42480
2 96697 1 42493
2 96698 1 42493
2 96699 1 42529
2 96700 1 42529
2 96701 1 42529
2 96702 1 42545
2 96703 1 42545
2 96704 1 42545
2 96705 1 42545
2 96706 1 42545
2 96707 1 42545
2 96708 1 42545
2 96709 1 42545
2 96710 1 42545
2 96711 1 42546
2 96712 1 42546
2 96713 1 42546
2 96714 1 42546
2 96715 1 42550
2 96716 1 42550
2 96717 1 42567
2 96718 1 42567
2 96719 1 42578
2 96720 1 42578
2 96721 1 42586
2 96722 1 42586
2 96723 1 42595
2 96724 1 42595
2 96725 1 42595
2 96726 1 42595
2 96727 1 42595
2 96728 1 42616
2 96729 1 42616
2 96730 1 42616
2 96731 1 42616
2 96732 1 42616
2 96733 1 42616
2 96734 1 42616
2 96735 1 42616
2 96736 1 42616
2 96737 1 42617
2 96738 1 42617
2 96739 1 42633
2 96740 1 42633
2 96741 1 42641
2 96742 1 42641
2 96743 1 42659
2 96744 1 42659
2 96745 1 42683
2 96746 1 42683
2 96747 1 42726
2 96748 1 42726
2 96749 1 42754
2 96750 1 42754
2 96751 1 42785
2 96752 1 42785
2 96753 1 42786
2 96754 1 42786
2 96755 1 42803
2 96756 1 42803
2 96757 1 42806
2 96758 1 42806
2 96759 1 42819
2 96760 1 42819
2 96761 1 42825
2 96762 1 42825
2 96763 1 42825
2 96764 1 42890
2 96765 1 42890
2 96766 1 42897
2 96767 1 42897
2 96768 1 42897
2 96769 1 42899
2 96770 1 42899
2 96771 1 42901
2 96772 1 42901
2 96773 1 42916
2 96774 1 42916
2 96775 1 42926
2 96776 1 42926
2 96777 1 42954
2 96778 1 42954
2 96779 1 42954
2 96780 1 42954
2 96781 1 42954
2 96782 1 42954
2 96783 1 42954
2 96784 1 42963
2 96785 1 42963
2 96786 1 43019
2 96787 1 43019
2 96788 1 43019
2 96789 1 43019
2 96790 1 43021
2 96791 1 43021
2 96792 1 43053
2 96793 1 43053
2 96794 1 43053
2 96795 1 43053
2 96796 1 43053
2 96797 1 43053
2 96798 1 43060
2 96799 1 43060
2 96800 1 43112
2 96801 1 43112
2 96802 1 43112
2 96803 1 43122
2 96804 1 43122
2 96805 1 43124
2 96806 1 43124
2 96807 1 43124
2 96808 1 43124
2 96809 1 43171
2 96810 1 43171
2 96811 1 43232
2 96812 1 43232
2 96813 1 43251
2 96814 1 43251
2 96815 1 43277
2 96816 1 43277
2 96817 1 43292
2 96818 1 43292
2 96819 1 43340
2 96820 1 43340
2 96821 1 43341
2 96822 1 43341
2 96823 1 43353
2 96824 1 43353
2 96825 1 43353
2 96826 1 43355
2 96827 1 43355
2 96828 1 43410
2 96829 1 43410
2 96830 1 43410
2 96831 1 43410
2 96832 1 43410
2 96833 1 43413
2 96834 1 43413
2 96835 1 43422
2 96836 1 43422
2 96837 1 43423
2 96838 1 43423
2 96839 1 43449
2 96840 1 43449
2 96841 1 43451
2 96842 1 43451
2 96843 1 43452
2 96844 1 43452
2 96845 1 43452
2 96846 1 43452
2 96847 1 43452
2 96848 1 43452
2 96849 1 43452
2 96850 1 43452
2 96851 1 43452
2 96852 1 43475
2 96853 1 43475
2 96854 1 43480
2 96855 1 43480
2 96856 1 43480
2 96857 1 43480
2 96858 1 43481
2 96859 1 43481
2 96860 1 43482
2 96861 1 43482
2 96862 1 43494
2 96863 1 43494
2 96864 1 43503
2 96865 1 43503
2 96866 1 43509
2 96867 1 43509
2 96868 1 43509
2 96869 1 43510
2 96870 1 43510
2 96871 1 43548
2 96872 1 43548
2 96873 1 43549
2 96874 1 43549
2 96875 1 43557
2 96876 1 43557
2 96877 1 43557
2 96878 1 43557
2 96879 1 43557
2 96880 1 43557
2 96881 1 43557
2 96882 1 43557
2 96883 1 43557
2 96884 1 43557
2 96885 1 43574
2 96886 1 43574
2 96887 1 43636
2 96888 1 43636
2 96889 1 43639
2 96890 1 43639
2 96891 1 43655
2 96892 1 43655
2 96893 1 43726
2 96894 1 43726
2 96895 1 43741
2 96896 1 43741
2 96897 1 43741
2 96898 1 43741
2 96899 1 43741
2 96900 1 43742
2 96901 1 43742
2 96902 1 43742
2 96903 1 43745
2 96904 1 43745
2 96905 1 43745
2 96906 1 43745
2 96907 1 43746
2 96908 1 43746
2 96909 1 43746
2 96910 1 43749
2 96911 1 43749
2 96912 1 43749
2 96913 1 43749
2 96914 1 43749
2 96915 1 43760
2 96916 1 43760
2 96917 1 43760
2 96918 1 43760
2 96919 1 43760
2 96920 1 43760
2 96921 1 43760
2 96922 1 43760
2 96923 1 43760
2 96924 1 43760
2 96925 1 43760
2 96926 1 43760
2 96927 1 43760
2 96928 1 43760
2 96929 1 43760
2 96930 1 43760
2 96931 1 43760
2 96932 1 43760
2 96933 1 43760
2 96934 1 43760
2 96935 1 43782
2 96936 1 43782
2 96937 1 43802
2 96938 1 43802
2 96939 1 43821
2 96940 1 43821
2 96941 1 43821
2 96942 1 43821
2 96943 1 43821
2 96944 1 43821
2 96945 1 43833
2 96946 1 43833
2 96947 1 43902
2 96948 1 43902
2 96949 1 43902
2 96950 1 43902
2 96951 1 43902
2 96952 1 43902
2 96953 1 43903
2 96954 1 43903
2 96955 1 43903
2 96956 1 43903
2 96957 1 43907
2 96958 1 43907
2 96959 1 43907
2 96960 1 43908
2 96961 1 43908
2 96962 1 43954
2 96963 1 43954
2 96964 1 43964
2 96965 1 43964
2 96966 1 43969
2 96967 1 43969
2 96968 1 44003
2 96969 1 44003
2 96970 1 44006
2 96971 1 44006
2 96972 1 44009
2 96973 1 44009
2 96974 1 44012
2 96975 1 44012
2 96976 1 44053
2 96977 1 44053
2 96978 1 44065
2 96979 1 44065
2 96980 1 44065
2 96981 1 44065
2 96982 1 44065
2 96983 1 44065
2 96984 1 44065
2 96985 1 44065
2 96986 1 44091
2 96987 1 44091
2 96988 1 44091
2 96989 1 44091
2 96990 1 44091
2 96991 1 44091
2 96992 1 44091
2 96993 1 44091
2 96994 1 44094
2 96995 1 44094
2 96996 1 44096
2 96997 1 44096
2 96998 1 44098
2 96999 1 44098
2 97000 1 44099
2 97001 1 44099
2 97002 1 44099
2 97003 1 44103
2 97004 1 44103
2 97005 1 44107
2 97006 1 44107
2 97007 1 44107
2 97008 1 44107
2 97009 1 44107
2 97010 1 44108
2 97011 1 44108
2 97012 1 44108
2 97013 1 44108
2 97014 1 44108
2 97015 1 44108
2 97016 1 44108
2 97017 1 44110
2 97018 1 44110
2 97019 1 44111
2 97020 1 44111
2 97021 1 44112
2 97022 1 44112
2 97023 1 44112
2 97024 1 44113
2 97025 1 44113
2 97026 1 44114
2 97027 1 44114
2 97028 1 44114
2 97029 1 44118
2 97030 1 44118
2 97031 1 44118
2 97032 1 44118
2 97033 1 44120
2 97034 1 44120
2 97035 1 44128
2 97036 1 44128
2 97037 1 44130
2 97038 1 44130
2 97039 1 44132
2 97040 1 44132
2 97041 1 44133
2 97042 1 44133
2 97043 1 44198
2 97044 1 44198
2 97045 1 44216
2 97046 1 44216
2 97047 1 44219
2 97048 1 44219
2 97049 1 44280
2 97050 1 44280
2 97051 1 44301
2 97052 1 44301
2 97053 1 44349
2 97054 1 44349
2 97055 1 44375
2 97056 1 44375
2 97057 1 44415
2 97058 1 44415
2 97059 1 44429
2 97060 1 44429
2 97061 1 44436
2 97062 1 44436
2 97063 1 44437
2 97064 1 44437
2 97065 1 44457
2 97066 1 44457
2 97067 1 44484
2 97068 1 44484
2 97069 1 44487
2 97070 1 44487
2 97071 1 44498
2 97072 1 44498
2 97073 1 44500
2 97074 1 44500
2 97075 1 44510
2 97076 1 44510
2 97077 1 44511
2 97078 1 44511
2 97079 1 44578
2 97080 1 44578
2 97081 1 44578
2 97082 1 44606
2 97083 1 44606
2 97084 1 44629
2 97085 1 44629
2 97086 1 44629
2 97087 1 44646
2 97088 1 44646
2 97089 1 44666
2 97090 1 44666
2 97091 1 44666
2 97092 1 44685
2 97093 1 44685
2 97094 1 44693
2 97095 1 44693
2 97096 1 44705
2 97097 1 44705
2 97098 1 44716
2 97099 1 44716
2 97100 1 44716
2 97101 1 44716
2 97102 1 44716
2 97103 1 44729
2 97104 1 44729
2 97105 1 44790
2 97106 1 44790
2 97107 1 44790
2 97108 1 44817
2 97109 1 44817
2 97110 1 44837
2 97111 1 44837
2 97112 1 44839
2 97113 1 44839
2 97114 1 44841
2 97115 1 44841
2 97116 1 44841
2 97117 1 44863
2 97118 1 44863
2 97119 1 44878
2 97120 1 44878
2 97121 1 44878
2 97122 1 44915
2 97123 1 44915
2 97124 1 45060
2 97125 1 45060
2 97126 1 45095
2 97127 1 45095
2 97128 1 45128
2 97129 1 45128
2 97130 1 45163
2 97131 1 45163
2 97132 1 45175
2 97133 1 45175
2 97134 1 45175
2 97135 1 45176
2 97136 1 45176
2 97137 1 45190
2 97138 1 45190
2 97139 1 45212
2 97140 1 45212
2 97141 1 45256
2 97142 1 45256
2 97143 1 45353
2 97144 1 45353
2 97145 1 45353
2 97146 1 45353
2 97147 1 45372
2 97148 1 45372
2 97149 1 45377
2 97150 1 45377
2 97151 1 45390
2 97152 1 45390
2 97153 1 45390
2 97154 1 45390
2 97155 1 45394
2 97156 1 45394
2 97157 1 45408
2 97158 1 45408
2 97159 1 45413
2 97160 1 45413
2 97161 1 45417
2 97162 1 45417
2 97163 1 45471
2 97164 1 45471
2 97165 1 45521
2 97166 1 45521
2 97167 1 45555
2 97168 1 45555
2 97169 1 45555
2 97170 1 45558
2 97171 1 45558
2 97172 1 45558
2 97173 1 45566
2 97174 1 45566
2 97175 1 45566
2 97176 1 45566
2 97177 1 45567
2 97178 1 45567
2 97179 1 45567
2 97180 1 45599
2 97181 1 45599
2 97182 1 45637
2 97183 1 45637
2 97184 1 45637
2 97185 1 45654
2 97186 1 45654
2 97187 1 45700
2 97188 1 45700
2 97189 1 45708
2 97190 1 45708
2 97191 1 45742
2 97192 1 45742
2 97193 1 45761
2 97194 1 45761
2 97195 1 45778
2 97196 1 45778
2 97197 1 45800
2 97198 1 45800
2 97199 1 45800
2 97200 1 45808
2 97201 1 45808
2 97202 1 45811
2 97203 1 45811
2 97204 1 45813
2 97205 1 45813
2 97206 1 45825
2 97207 1 45825
2 97208 1 45832
2 97209 1 45832
2 97210 1 45832
2 97211 1 45832
2 97212 1 45832
2 97213 1 45832
2 97214 1 45833
2 97215 1 45833
2 97216 1 45910
2 97217 1 45910
2 97218 1 45924
2 97219 1 45924
2 97220 1 45956
2 97221 1 45956
2 97222 1 46063
2 97223 1 46063
2 97224 1 46077
2 97225 1 46077
2 97226 1 46181
2 97227 1 46181
2 97228 1 46182
2 97229 1 46182
2 97230 1 46262
2 97231 1 46262
2 97232 1 46294
2 97233 1 46294
2 97234 1 46302
2 97235 1 46302
2 97236 1 46303
2 97237 1 46303
2 97238 1 46303
2 97239 1 46326
2 97240 1 46326
2 97241 1 46350
2 97242 1 46350
2 97243 1 46483
2 97244 1 46483
2 97245 1 46485
2 97246 1 46485
2 97247 1 46491
2 97248 1 46491
2 97249 1 46502
2 97250 1 46502
2 97251 1 46531
2 97252 1 46531
2 97253 1 46537
2 97254 1 46537
2 97255 1 46537
2 97256 1 46537
2 97257 1 46537
2 97258 1 46537
2 97259 1 46537
2 97260 1 46538
2 97261 1 46538
2 97262 1 46541
2 97263 1 46541
2 97264 1 46555
2 97265 1 46555
2 97266 1 46556
2 97267 1 46556
2 97268 1 46558
2 97269 1 46558
2 97270 1 46567
2 97271 1 46567
2 97272 1 46570
2 97273 1 46570
2 97274 1 46572
2 97275 1 46572
2 97276 1 46574
2 97277 1 46574
2 97278 1 46577
2 97279 1 46577
2 97280 1 46607
2 97281 1 46607
2 97282 1 46632
2 97283 1 46632
2 97284 1 46633
2 97285 1 46633
2 97286 1 46633
2 97287 1 46633
2 97288 1 46633
2 97289 1 46633
2 97290 1 46637
2 97291 1 46637
2 97292 1 46721
2 97293 1 46721
2 97294 1 46748
2 97295 1 46748
2 97296 1 46778
2 97297 1 46778
2 97298 1 46851
2 97299 1 46851
2 97300 1 46852
2 97301 1 46852
2 97302 1 46884
2 97303 1 46884
2 97304 1 46885
2 97305 1 46885
2 97306 1 46898
2 97307 1 46898
2 97308 1 46898
2 97309 1 46899
2 97310 1 46899
2 97311 1 46899
2 97312 1 46899
2 97313 1 46933
2 97314 1 46933
2 97315 1 47017
2 97316 1 47017
2 97317 1 47218
2 97318 1 47218
2 97319 1 47335
2 97320 1 47335
2 97321 1 47372
2 97322 1 47372
2 97323 1 47373
2 97324 1 47373
2 97325 1 47375
2 97326 1 47375
2 97327 1 47401
2 97328 1 47401
2 97329 1 47401
2 97330 1 47401
2 97331 1 47444
2 97332 1 47444
2 97333 1 47444
2 97334 1 47444
2 97335 1 47445
2 97336 1 47445
2 97337 1 47446
2 97338 1 47446
2 97339 1 47483
2 97340 1 47483
2 97341 1 47553
2 97342 1 47553
2 97343 1 47565
2 97344 1 47565
2 97345 1 47565
2 97346 1 47565
2 97347 1 47566
2 97348 1 47566
2 97349 1 47567
2 97350 1 47567
2 97351 1 47567
2 97352 1 47571
2 97353 1 47571
2 97354 1 47592
2 97355 1 47592
2 97356 1 47599
2 97357 1 47599
2 97358 1 47599
2 97359 1 47599
2 97360 1 47599
2 97361 1 47639
2 97362 1 47639
2 97363 1 47644
2 97364 1 47644
2 97365 1 47657
2 97366 1 47657
2 97367 1 47664
2 97368 1 47664
2 97369 1 47674
2 97370 1 47674
2 97371 1 47674
2 97372 1 47674
2 97373 1 47674
2 97374 1 47674
2 97375 1 47676
2 97376 1 47676
2 97377 1 47676
2 97378 1 47677
2 97379 1 47677
2 97380 1 47687
2 97381 1 47687
2 97382 1 47688
2 97383 1 47688
2 97384 1 47697
2 97385 1 47697
2 97386 1 47698
2 97387 1 47698
2 97388 1 47698
2 97389 1 47698
2 97390 1 47731
2 97391 1 47731
2 97392 1 47731
2 97393 1 47740
2 97394 1 47740
2 97395 1 47779
2 97396 1 47779
2 97397 1 47779
2 97398 1 47779
2 97399 1 47779
2 97400 1 47779
2 97401 1 47779
2 97402 1 47779
2 97403 1 47779
2 97404 1 47779
2 97405 1 47779
2 97406 1 47779
2 97407 1 47779
2 97408 1 47779
2 97409 1 47779
2 97410 1 47779
2 97411 1 47779
2 97412 1 47779
2 97413 1 47779
2 97414 1 47781
2 97415 1 47781
2 97416 1 47782
2 97417 1 47782
2 97418 1 47790
2 97419 1 47790
2 97420 1 47796
2 97421 1 47796
2 97422 1 47804
2 97423 1 47804
2 97424 1 47804
2 97425 1 47804
2 97426 1 47804
2 97427 1 47804
2 97428 1 47804
2 97429 1 47805
2 97430 1 47805
2 97431 1 47805
2 97432 1 47805
2 97433 1 47805
2 97434 1 47805
2 97435 1 47805
2 97436 1 47805
2 97437 1 47805
2 97438 1 47805
2 97439 1 47805
2 97440 1 47805
2 97441 1 47805
2 97442 1 47805
2 97443 1 47825
2 97444 1 47825
2 97445 1 47832
2 97446 1 47832
2 97447 1 47832
2 97448 1 47832
2 97449 1 47842
2 97450 1 47842
2 97451 1 47842
2 97452 1 47843
2 97453 1 47843
2 97454 1 47843
2 97455 1 47844
2 97456 1 47844
2 97457 1 47845
2 97458 1 47845
2 97459 1 47846
2 97460 1 47846
2 97461 1 47846
2 97462 1 47856
2 97463 1 47856
2 97464 1 47862
2 97465 1 47862
2 97466 1 47876
2 97467 1 47876
2 97468 1 47876
2 97469 1 47876
2 97470 1 47876
2 97471 1 47876
2 97472 1 47877
2 97473 1 47877
2 97474 1 47885
2 97475 1 47885
2 97476 1 47885
2 97477 1 47885
2 97478 1 47886
2 97479 1 47886
2 97480 1 47886
2 97481 1 47887
2 97482 1 47887
2 97483 1 47896
2 97484 1 47896
2 97485 1 47897
2 97486 1 47897
2 97487 1 47899
2 97488 1 47899
2 97489 1 47899
2 97490 1 47907
2 97491 1 47907
2 97492 1 47907
2 97493 1 47915
2 97494 1 47915
2 97495 1 47915
2 97496 1 47928
2 97497 1 47928
2 97498 1 47928
2 97499 1 47939
2 97500 1 47939
2 97501 1 47942
2 97502 1 47942
2 97503 1 47945
2 97504 1 47945
2 97505 1 47960
2 97506 1 47960
2 97507 1 47960
2 97508 1 47966
2 97509 1 47966
2 97510 1 47975
2 97511 1 47975
2 97512 1 47985
2 97513 1 47985
2 97514 1 48003
2 97515 1 48003
2 97516 1 48003
2 97517 1 48003
2 97518 1 48011
2 97519 1 48011
2 97520 1 48011
2 97521 1 48012
2 97522 1 48012
2 97523 1 48019
2 97524 1 48019
2 97525 1 48032
2 97526 1 48032
2 97527 1 48032
2 97528 1 48032
2 97529 1 48039
2 97530 1 48039
2 97531 1 48048
2 97532 1 48048
2 97533 1 48056
2 97534 1 48056
2 97535 1 48056
2 97536 1 48056
2 97537 1 48057
2 97538 1 48057
2 97539 1 48069
2 97540 1 48069
2 97541 1 48084
2 97542 1 48084
2 97543 1 48110
2 97544 1 48110
2 97545 1 48110
2 97546 1 48123
2 97547 1 48123
2 97548 1 48124
2 97549 1 48124
2 97550 1 48124
2 97551 1 48128
2 97552 1 48128
2 97553 1 48140
2 97554 1 48140
2 97555 1 48160
2 97556 1 48160
2 97557 1 48162
2 97558 1 48162
2 97559 1 48163
2 97560 1 48163
2 97561 1 48192
2 97562 1 48192
2 97563 1 48201
2 97564 1 48201
2 97565 1 48201
2 97566 1 48202
2 97567 1 48202
2 97568 1 48210
2 97569 1 48210
2 97570 1 48210
2 97571 1 48211
2 97572 1 48211
2 97573 1 48212
2 97574 1 48212
2 97575 1 48212
2 97576 1 48233
2 97577 1 48233
2 97578 1 48233
2 97579 1 48233
2 97580 1 48233
2 97581 1 48245
2 97582 1 48245
2 97583 1 48254
2 97584 1 48254
2 97585 1 48254
2 97586 1 48254
2 97587 1 48254
2 97588 1 48254
2 97589 1 48255
2 97590 1 48255
2 97591 1 48270
2 97592 1 48270
2 97593 1 48271
2 97594 1 48271
2 97595 1 48274
2 97596 1 48274
2 97597 1 48274
2 97598 1 48275
2 97599 1 48275
2 97600 1 48277
2 97601 1 48277
2 97602 1 48277
2 97603 1 48277
2 97604 1 48294
2 97605 1 48294
2 97606 1 48295
2 97607 1 48295
2 97608 1 48297
2 97609 1 48297
2 97610 1 48301
2 97611 1 48301
2 97612 1 48301
2 97613 1 48302
2 97614 1 48302
2 97615 1 48303
2 97616 1 48303
2 97617 1 48304
2 97618 1 48304
2 97619 1 48306
2 97620 1 48306
2 97621 1 48308
2 97622 1 48308
2 97623 1 48323
2 97624 1 48323
2 97625 1 48324
2 97626 1 48324
2 97627 1 48326
2 97628 1 48326
2 97629 1 48326
2 97630 1 48335
2 97631 1 48335
2 97632 1 48335
2 97633 1 48337
2 97634 1 48337
2 97635 1 48337
2 97636 1 48338
2 97637 1 48338
2 97638 1 48347
2 97639 1 48347
2 97640 1 48347
2 97641 1 48350
2 97642 1 48350
2 97643 1 48350
2 97644 1 48351
2 97645 1 48351
2 97646 1 48351
2 97647 1 48351
2 97648 1 48351
2 97649 1 48359
2 97650 1 48359
2 97651 1 48362
2 97652 1 48362
2 97653 1 48362
2 97654 1 48362
2 97655 1 48362
2 97656 1 48362
2 97657 1 48363
2 97658 1 48363
2 97659 1 48369
2 97660 1 48369
2 97661 1 48369
2 97662 1 48369
2 97663 1 48369
2 97664 1 48369
2 97665 1 48370
2 97666 1 48370
2 97667 1 48370
2 97668 1 48378
2 97669 1 48378
2 97670 1 48378
2 97671 1 48378
2 97672 1 48378
2 97673 1 48379
2 97674 1 48379
2 97675 1 48379
2 97676 1 48380
2 97677 1 48380
2 97678 1 48381
2 97679 1 48381
2 97680 1 48381
2 97681 1 48381
2 97682 1 48383
2 97683 1 48383
2 97684 1 48383
2 97685 1 48392
2 97686 1 48392
2 97687 1 48410
2 97688 1 48410
2 97689 1 48410
2 97690 1 48411
2 97691 1 48411
2 97692 1 48426
2 97693 1 48426
2 97694 1 48426
2 97695 1 48429
2 97696 1 48429
2 97697 1 48429
2 97698 1 48430
2 97699 1 48430
2 97700 1 48430
2 97701 1 48431
2 97702 1 48431
2 97703 1 48431
2 97704 1 48432
2 97705 1 48432
2 97706 1 48444
2 97707 1 48444
2 97708 1 48448
2 97709 1 48448
2 97710 1 48471
2 97711 1 48471
2 97712 1 48474
2 97713 1 48474
2 97714 1 48474
2 97715 1 48474
2 97716 1 48484
2 97717 1 48484
2 97718 1 48495
2 97719 1 48495
2 97720 1 48497
2 97721 1 48497
2 97722 1 48521
2 97723 1 48521
2 97724 1 48521
2 97725 1 48522
2 97726 1 48522
2 97727 1 48522
2 97728 1 48522
2 97729 1 48551
2 97730 1 48551
2 97731 1 48560
2 97732 1 48560
2 97733 1 48560
2 97734 1 48560
2 97735 1 48560
2 97736 1 48560
2 97737 1 48569
2 97738 1 48569
2 97739 1 48569
2 97740 1 48569
2 97741 1 48569
2 97742 1 48569
2 97743 1 48569
2 97744 1 48569
2 97745 1 48570
2 97746 1 48570
2 97747 1 48570
2 97748 1 48575
2 97749 1 48575
2 97750 1 48575
2 97751 1 48576
2 97752 1 48576
2 97753 1 48585
2 97754 1 48585
2 97755 1 48585
2 97756 1 48591
2 97757 1 48591
2 97758 1 48591
2 97759 1 48591
2 97760 1 48592
2 97761 1 48592
2 97762 1 48637
2 97763 1 48637
2 97764 1 48637
2 97765 1 48637
2 97766 1 48637
2 97767 1 48637
2 97768 1 48637
2 97769 1 48637
2 97770 1 48637
2 97771 1 48637
2 97772 1 48650
2 97773 1 48650
2 97774 1 48650
2 97775 1 48650
2 97776 1 48650
2 97777 1 48650
2 97778 1 48662
2 97779 1 48662
2 97780 1 48674
2 97781 1 48674
2 97782 1 48703
2 97783 1 48703
2 97784 1 48707
2 97785 1 48707
2 97786 1 48707
2 97787 1 48732
2 97788 1 48732
2 97789 1 48732
2 97790 1 48732
2 97791 1 48732
2 97792 1 48747
2 97793 1 48747
2 97794 1 48747
2 97795 1 48755
2 97796 1 48755
2 97797 1 48755
2 97798 1 48755
2 97799 1 48755
2 97800 1 48755
2 97801 1 48755
2 97802 1 48755
2 97803 1 48755
2 97804 1 48755
2 97805 1 48755
2 97806 1 48755
2 97807 1 48758
2 97808 1 48758
2 97809 1 48759
2 97810 1 48759
2 97811 1 48766
2 97812 1 48766
2 97813 1 48770
2 97814 1 48770
2 97815 1 48770
2 97816 1 48770
2 97817 1 48772
2 97818 1 48772
2 97819 1 48774
2 97820 1 48774
2 97821 1 48775
2 97822 1 48775
2 97823 1 48803
2 97824 1 48803
2 97825 1 48803
2 97826 1 48836
2 97827 1 48836
2 97828 1 48837
2 97829 1 48837
2 97830 1 48840
2 97831 1 48840
2 97832 1 48840
2 97833 1 48849
2 97834 1 48849
2 97835 1 48850
2 97836 1 48850
2 97837 1 48882
2 97838 1 48882
2 97839 1 48903
2 97840 1 48903
2 97841 1 48904
2 97842 1 48904
2 97843 1 48914
2 97844 1 48914
2 97845 1 48914
2 97846 1 48914
2 97847 1 48914
2 97848 1 48923
2 97849 1 48923
2 97850 1 48924
2 97851 1 48924
2 97852 1 48954
2 97853 1 48954
2 97854 1 48954
2 97855 1 48962
2 97856 1 48962
2 97857 1 48962
2 97858 1 48962
2 97859 1 48962
2 97860 1 48963
2 97861 1 48963
2 97862 1 48965
2 97863 1 48965
2 97864 1 49017
2 97865 1 49017
2 97866 1 49035
2 97867 1 49035
2 97868 1 49041
2 97869 1 49041
2 97870 1 49048
2 97871 1 49048
2 97872 1 49048
2 97873 1 49083
2 97874 1 49083
2 97875 1 49083
2 97876 1 49083
2 97877 1 49088
2 97878 1 49088
2 97879 1 49092
2 97880 1 49092
2 97881 1 49126
2 97882 1 49126
2 97883 1 49141
2 97884 1 49141
2 97885 1 49142
2 97886 1 49142
2 97887 1 49142
2 97888 1 49150
2 97889 1 49150
2 97890 1 49150
2 97891 1 49150
2 97892 1 49157
2 97893 1 49157
2 97894 1 49179
2 97895 1 49179
2 97896 1 49198
2 97897 1 49198
2 97898 1 49199
2 97899 1 49199
2 97900 1 49199
2 97901 1 49214
2 97902 1 49214
2 97903 1 49230
2 97904 1 49230
2 97905 1 49261
2 97906 1 49261
2 97907 1 49298
2 97908 1 49298
2 97909 1 49331
2 97910 1 49331
2 97911 1 49388
2 97912 1 49388
2 97913 1 49393
2 97914 1 49393
2 97915 1 49397
2 97916 1 49397
2 97917 1 49397
2 97918 1 49397
2 97919 1 49401
2 97920 1 49401
2 97921 1 49401
2 97922 1 49401
2 97923 1 49416
2 97924 1 49416
2 97925 1 49418
2 97926 1 49418
2 97927 1 49419
2 97928 1 49419
2 97929 1 49419
2 97930 1 49432
2 97931 1 49432
2 97932 1 49432
2 97933 1 49433
2 97934 1 49433
2 97935 1 49467
2 97936 1 49467
2 97937 1 49467
2 97938 1 49468
2 97939 1 49468
2 97940 1 49468
2 97941 1 49470
2 97942 1 49470
2 97943 1 49487
2 97944 1 49487
2 97945 1 49496
2 97946 1 49496
2 97947 1 49496
2 97948 1 49496
2 97949 1 49523
2 97950 1 49523
2 97951 1 49524
2 97952 1 49524
2 97953 1 49526
2 97954 1 49526
2 97955 1 49532
2 97956 1 49532
2 97957 1 49532
2 97958 1 49539
2 97959 1 49539
2 97960 1 49583
2 97961 1 49583
2 97962 1 49583
2 97963 1 49601
2 97964 1 49601
2 97965 1 49618
2 97966 1 49618
2 97967 1 49619
2 97968 1 49619
2 97969 1 49628
2 97970 1 49628
2 97971 1 49630
2 97972 1 49630
2 97973 1 49630
2 97974 1 49630
2 97975 1 49643
2 97976 1 49643
2 97977 1 49662
2 97978 1 49662
2 97979 1 49663
2 97980 1 49663
2 97981 1 49666
2 97982 1 49666
2 97983 1 49678
2 97984 1 49678
2 97985 1 49678
2 97986 1 49725
2 97987 1 49725
2 97988 1 49733
2 97989 1 49733
2 97990 1 49743
2 97991 1 49743
2 97992 1 49743
2 97993 1 49743
2 97994 1 49776
2 97995 1 49776
2 97996 1 49778
2 97997 1 49778
2 97998 1 49785
2 97999 1 49785
2 98000 1 49793
2 98001 1 49793
2 98002 1 49793
2 98003 1 49793
2 98004 1 49809
2 98005 1 49809
2 98006 1 49810
2 98007 1 49810
2 98008 1 49817
2 98009 1 49817
2 98010 1 49818
2 98011 1 49818
2 98012 1 49861
2 98013 1 49861
2 98014 1 49869
2 98015 1 49869
2 98016 1 49870
2 98017 1 49870
2 98018 1 49870
2 98019 1 49870
2 98020 1 49870
2 98021 1 49870
2 98022 1 49870
2 98023 1 49870
2 98024 1 49870
2 98025 1 49870
2 98026 1 49870
2 98027 1 49870
2 98028 1 49870
2 98029 1 49870
2 98030 1 49870
2 98031 1 49871
2 98032 1 49871
2 98033 1 49871
2 98034 1 49894
2 98035 1 49894
2 98036 1 49903
2 98037 1 49903
2 98038 1 49903
2 98039 1 49903
2 98040 1 49903
2 98041 1 49903
2 98042 1 49915
2 98043 1 49915
2 98044 1 49942
2 98045 1 49942
2 98046 1 49949
2 98047 1 49949
2 98048 1 49965
2 98049 1 49965
2 98050 1 49965
2 98051 1 49998
2 98052 1 49998
2 98053 1 49998
2 98054 1 50001
2 98055 1 50001
2 98056 1 50001
2 98057 1 50006
2 98058 1 50006
2 98059 1 50013
2 98060 1 50013
2 98061 1 50013
2 98062 1 50015
2 98063 1 50015
2 98064 1 50026
2 98065 1 50026
2 98066 1 50040
2 98067 1 50040
2 98068 1 50041
2 98069 1 50041
2 98070 1 50044
2 98071 1 50044
2 98072 1 50047
2 98073 1 50047
2 98074 1 50047
2 98075 1 50050
2 98076 1 50050
2 98077 1 50054
2 98078 1 50054
2 98079 1 50054
2 98080 1 50054
2 98081 1 50054
2 98082 1 50072
2 98083 1 50072
2 98084 1 50072
2 98085 1 50073
2 98086 1 50073
2 98087 1 50073
2 98088 1 50073
2 98089 1 50084
2 98090 1 50084
2 98091 1 50088
2 98092 1 50088
2 98093 1 50091
2 98094 1 50091
2 98095 1 50091
2 98096 1 50115
2 98097 1 50115
2 98098 1 50115
2 98099 1 50123
2 98100 1 50123
2 98101 1 50125
2 98102 1 50125
2 98103 1 50126
2 98104 1 50126
2 98105 1 50149
2 98106 1 50149
2 98107 1 50168
2 98108 1 50168
2 98109 1 50182
2 98110 1 50182
2 98111 1 50194
2 98112 1 50194
2 98113 1 50196
2 98114 1 50196
2 98115 1 50222
2 98116 1 50222
2 98117 1 50231
2 98118 1 50231
2 98119 1 50232
2 98120 1 50232
2 98121 1 50232
2 98122 1 50251
2 98123 1 50251
2 98124 1 50251
2 98125 1 50277
2 98126 1 50277
2 98127 1 50280
2 98128 1 50280
2 98129 1 50281
2 98130 1 50281
2 98131 1 50314
2 98132 1 50314
2 98133 1 50317
2 98134 1 50317
2 98135 1 50338
2 98136 1 50338
2 98137 1 50346
2 98138 1 50346
2 98139 1 50371
2 98140 1 50371
2 98141 1 50371
2 98142 1 50379
2 98143 1 50379
2 98144 1 50379
2 98145 1 50379
2 98146 1 50426
2 98147 1 50426
2 98148 1 50456
2 98149 1 50456
2 98150 1 50495
2 98151 1 50495
2 98152 1 50535
2 98153 1 50535
2 98154 1 50544
2 98155 1 50544
2 98156 1 50545
2 98157 1 50545
2 98158 1 50585
2 98159 1 50585
2 98160 1 50620
2 98161 1 50620
2 98162 1 50635
2 98163 1 50635
2 98164 1 50644
2 98165 1 50644
2 98166 1 50644
2 98167 1 50665
2 98168 1 50665
2 98169 1 50665
2 98170 1 50665
2 98171 1 50666
2 98172 1 50666
2 98173 1 50673
2 98174 1 50673
2 98175 1 50673
2 98176 1 50674
2 98177 1 50674
2 98178 1 50684
2 98179 1 50684
2 98180 1 50684
2 98181 1 50684
2 98182 1 50732
2 98183 1 50732
2 98184 1 50751
2 98185 1 50751
2 98186 1 50758
2 98187 1 50758
2 98188 1 50763
2 98189 1 50763
2 98190 1 50772
2 98191 1 50772
2 98192 1 50772
2 98193 1 50772
2 98194 1 50785
2 98195 1 50785
2 98196 1 50785
2 98197 1 50785
2 98198 1 50785
2 98199 1 50799
2 98200 1 50799
2 98201 1 50800
2 98202 1 50800
2 98203 1 50811
2 98204 1 50811
2 98205 1 50811
2 98206 1 50818
2 98207 1 50818
2 98208 1 50818
2 98209 1 50818
2 98210 1 50826
2 98211 1 50826
2 98212 1 50826
2 98213 1 50827
2 98214 1 50827
2 98215 1 50845
2 98216 1 50845
2 98217 1 50846
2 98218 1 50846
2 98219 1 50867
2 98220 1 50867
2 98221 1 50867
2 98222 1 50867
2 98223 1 50896
2 98224 1 50896
2 98225 1 50902
2 98226 1 50902
2 98227 1 50916
2 98228 1 50916
2 98229 1 50930
2 98230 1 50930
2 98231 1 50967
2 98232 1 50967
2 98233 1 50980
2 98234 1 50980
2 98235 1 50980
2 98236 1 51001
2 98237 1 51001
2 98238 1 51005
2 98239 1 51005
2 98240 1 51014
2 98241 1 51014
2 98242 1 51037
2 98243 1 51037
2 98244 1 51040
2 98245 1 51040
2 98246 1 51040
2 98247 1 51040
2 98248 1 51040
2 98249 1 51084
2 98250 1 51084
2 98251 1 51115
2 98252 1 51115
2 98253 1 51124
2 98254 1 51124
2 98255 1 51156
2 98256 1 51156
2 98257 1 51157
2 98258 1 51157
2 98259 1 51159
2 98260 1 51159
2 98261 1 51161
2 98262 1 51161
2 98263 1 51171
2 98264 1 51171
2 98265 1 51173
2 98266 1 51173
2 98267 1 51173
2 98268 1 51175
2 98269 1 51175
2 98270 1 51184
2 98271 1 51184
2 98272 1 51184
2 98273 1 51235
2 98274 1 51235
2 98275 1 51270
2 98276 1 51270
2 98277 1 51271
2 98278 1 51271
2 98279 1 51272
2 98280 1 51272
2 98281 1 51280
2 98282 1 51280
2 98283 1 51280
2 98284 1 51281
2 98285 1 51281
2 98286 1 51283
2 98287 1 51283
2 98288 1 51288
2 98289 1 51288
2 98290 1 51289
2 98291 1 51289
2 98292 1 51293
2 98293 1 51293
2 98294 1 51293
2 98295 1 51293
2 98296 1 51308
2 98297 1 51308
2 98298 1 51308
2 98299 1 51319
2 98300 1 51319
2 98301 1 51322
2 98302 1 51322
2 98303 1 51322
2 98304 1 51322
2 98305 1 51323
2 98306 1 51323
2 98307 1 51328
2 98308 1 51328
2 98309 1 51339
2 98310 1 51339
2 98311 1 51352
2 98312 1 51352
2 98313 1 51385
2 98314 1 51385
2 98315 1 51387
2 98316 1 51387
2 98317 1 51401
2 98318 1 51401
2 98319 1 51403
2 98320 1 51403
2 98321 1 51403
2 98322 1 51437
2 98323 1 51437
2 98324 1 51437
2 98325 1 51437
2 98326 1 51437
2 98327 1 51447
2 98328 1 51447
2 98329 1 51461
2 98330 1 51461
2 98331 1 51461
2 98332 1 51461
2 98333 1 51461
2 98334 1 51461
2 98335 1 51489
2 98336 1 51489
2 98337 1 51516
2 98338 1 51516
2 98339 1 51540
2 98340 1 51540
2 98341 1 51562
2 98342 1 51562
2 98343 1 51566
2 98344 1 51566
2 98345 1 51567
2 98346 1 51567
2 98347 1 51571
2 98348 1 51571
2 98349 1 51588
2 98350 1 51588
2 98351 1 51606
2 98352 1 51606
2 98353 1 51606
2 98354 1 51611
2 98355 1 51611
2 98356 1 51620
2 98357 1 51620
2 98358 1 51620
2 98359 1 51623
2 98360 1 51623
2 98361 1 51626
2 98362 1 51626
2 98363 1 51626
2 98364 1 51626
2 98365 1 51628
2 98366 1 51628
2 98367 1 51628
2 98368 1 51659
2 98369 1 51659
2 98370 1 51661
2 98371 1 51661
2 98372 1 51663
2 98373 1 51663
2 98374 1 51688
2 98375 1 51688
2 98376 1 51707
2 98377 1 51707
2 98378 1 51716
2 98379 1 51716
2 98380 1 51757
2 98381 1 51757
2 98382 1 51760
2 98383 1 51760
2 98384 1 51762
2 98385 1 51762
2 98386 1 51790
2 98387 1 51790
2 98388 1 51827
2 98389 1 51827
2 98390 1 51838
2 98391 1 51838
2 98392 1 51843
2 98393 1 51843
2 98394 1 51893
2 98395 1 51893
2 98396 1 51893
2 98397 1 51940
2 98398 1 51940
2 98399 1 51948
2 98400 1 51948
2 98401 1 51962
2 98402 1 51962
2 98403 1 51963
2 98404 1 51963
2 98405 1 51971
2 98406 1 51971
2 98407 1 52021
2 98408 1 52021
2 98409 1 52043
2 98410 1 52043
2 98411 1 52067
2 98412 1 52067
2 98413 1 52067
2 98414 1 52068
2 98415 1 52068
2 98416 1 52101
2 98417 1 52101
2 98418 1 52111
2 98419 1 52111
2 98420 1 52135
2 98421 1 52135
2 98422 1 52163
2 98423 1 52163
2 98424 1 52176
2 98425 1 52176
2 98426 1 52218
2 98427 1 52218
2 98428 1 52233
2 98429 1 52233
2 98430 1 52245
2 98431 1 52245
2 98432 1 52248
2 98433 1 52248
2 98434 1 52249
2 98435 1 52249
2 98436 1 52310
2 98437 1 52310
2 98438 1 52504
2 98439 1 52504
2 98440 1 52525
2 98441 1 52525
2 98442 1 52525
2 98443 1 52525
2 98444 1 52525
2 98445 1 52543
2 98446 1 52543
2 98447 1 52567
2 98448 1 52567
2 98449 1 52591
2 98450 1 52591
2 98451 1 52619
2 98452 1 52619
2 98453 1 52630
2 98454 1 52630
2 98455 1 52705
2 98456 1 52705
2 98457 1 52720
2 98458 1 52720
2 98459 1 52779
2 98460 1 52779
2 98461 1 52788
2 98462 1 52788
2 98463 1 52788
2 98464 1 52789
2 98465 1 52789
2 98466 1 52800
2 98467 1 52800
2 98468 1 52829
2 98469 1 52829
2 98470 1 52829
2 98471 1 52857
2 98472 1 52857
2 98473 1 52866
2 98474 1 52866
2 98475 1 52892
2 98476 1 52892
2 98477 1 52895
2 98478 1 52895
2 98479 1 52908
2 98480 1 52908
2 98481 1 52920
2 98482 1 52920
2 98483 1 52931
2 98484 1 52931
2 98485 1 53041
2 98486 1 53041
2 98487 1 53042
2 98488 1 53042
2 98489 1 53047
2 98490 1 53047
2 98491 1 53134
2 98492 1 53134
2 98493 1 53137
2 98494 1 53137
2 98495 1 53191
2 98496 1 53191
2 98497 1 53212
2 98498 1 53212
2 98499 1 53214
2 98500 1 53214
2 98501 1 53230
2 98502 1 53230
2 98503 1 53253
2 98504 1 53253
2 98505 1 53261
2 98506 1 53261
2 98507 1 53263
2 98508 1 53263
2 98509 1 53292
2 98510 1 53292
2 98511 1 53338
2 98512 1 53338
2 98513 1 53338
2 98514 1 53409
2 98515 1 53409
2 98516 1 53457
2 98517 1 53457
2 98518 1 53457
2 98519 1 53470
2 98520 1 53470
2 98521 1 53482
2 98522 1 53482
2 98523 1 53502
2 98524 1 53502
2 98525 1 53510
2 98526 1 53510
2 98527 1 53581
2 98528 1 53581
2 98529 1 53582
2 98530 1 53582
2 98531 1 53600
2 98532 1 53600
2 98533 1 53600
2 98534 1 53600
2 98535 1 53600
2 98536 1 53601
2 98537 1 53601
2 98538 1 53605
2 98539 1 53605
2 98540 1 53653
2 98541 1 53653
2 98542 1 53712
2 98543 1 53712
2 98544 1 53762
2 98545 1 53762
2 98546 1 53763
2 98547 1 53763
2 98548 1 53820
2 98549 1 53820
2 98550 1 53820
2 98551 1 53835
2 98552 1 53835
2 98553 1 53835
2 98554 1 53868
2 98555 1 53868
2 98556 1 53890
2 98557 1 53890
2 98558 1 53896
2 98559 1 53896
2 98560 1 53956
2 98561 1 53956
2 98562 1 53987
2 98563 1 53987
2 98564 1 53988
2 98565 1 53988
2 98566 1 54058
2 98567 1 54058
2 98568 1 54065
2 98569 1 54065
2 98570 1 54067
2 98571 1 54067
2 98572 1 54096
2 98573 1 54096
2 98574 1 54377
2 98575 1 54377
2 98576 1 54715
2 98577 1 54715
2 98578 1 54927
2 98579 1 54927
2 98580 1 54960
2 98581 1 54960
2 98582 1 54962
2 98583 1 54962
2 98584 1 54973
2 98585 1 54973
2 98586 1 54978
2 98587 1 54978
2 98588 1 54981
2 98589 1 54981
2 98590 1 55031
2 98591 1 55031
2 98592 1 55056
2 98593 1 55056
2 98594 1 55057
2 98595 1 55057
2 98596 1 55064
2 98597 1 55064
2 98598 1 55330
2 98599 1 55330
2 98600 1 55536
2 98601 1 55536
2 98602 1 55539
2 98603 1 55539
2 98604 1 55547
2 98605 1 55547
2 98606 1 55588
2 98607 1 55588
2 98608 1 55590
2 98609 1 55590
2 98610 1 55590
2 98611 1 55596
2 98612 1 55596
2 98613 1 55614
2 98614 1 55614
2 98615 1 55653
2 98616 1 55653
2 98617 1 55682
2 98618 1 55682
2 98619 1 55697
2 98620 1 55697
2 98621 1 55733
2 98622 1 55733
2 98623 1 55776
2 98624 1 55776
2 98625 1 55782
2 98626 1 55782
2 98627 1 55782
2 98628 1 55782
2 98629 1 55782
2 98630 1 55846
2 98631 1 55846
2 98632 1 55857
2 98633 1 55857
2 98634 1 55917
2 98635 1 55917
2 98636 1 55917
2 98637 1 55917
2 98638 1 55921
2 98639 1 55921
2 98640 1 56019
2 98641 1 56019
2 98642 1 56046
2 98643 1 56046
2 98644 1 56061
2 98645 1 56061
2 98646 1 56061
2 98647 1 56082
2 98648 1 56082
2 98649 1 56284
2 98650 1 56284
2 98651 1 56287
2 98652 1 56287
2 98653 1 56287
2 98654 1 56334
2 98655 1 56334
2 98656 1 56334
2 98657 1 56358
2 98658 1 56358
2 98659 1 56384
2 98660 1 56384
2 98661 1 56384
2 98662 1 56476
2 98663 1 56476
2 98664 1 56477
2 98665 1 56477
2 98666 1 56590
2 98667 1 56590
2 98668 1 56672
2 98669 1 56672
2 98670 1 56711
2 98671 1 56711
2 98672 1 56714
2 98673 1 56714
2 98674 1 56747
2 98675 1 56747
2 98676 1 56756
2 98677 1 56756
2 98678 1 56818
2 98679 1 56818
2 98680 1 56885
2 98681 1 56885
2 98682 1 56937
2 98683 1 56937
2 98684 1 56938
2 98685 1 56938
2 98686 1 56952
2 98687 1 56952
2 98688 1 56953
2 98689 1 56953
2 98690 1 56971
2 98691 1 56971
2 98692 1 56976
2 98693 1 56976
2 98694 1 57008
2 98695 1 57008
2 98696 1 57044
2 98697 1 57044
2 98698 1 57051
2 98699 1 57051
2 98700 1 57054
2 98701 1 57054
2 98702 1 57073
2 98703 1 57073
2 98704 1 57073
2 98705 1 57094
2 98706 1 57094
2 98707 1 57101
2 98708 1 57101
2 98709 1 57174
2 98710 1 57174
2 98711 1 57257
2 98712 1 57257
2 98713 1 57262
2 98714 1 57262
2 98715 1 57262
2 98716 1 57294
2 98717 1 57294
2 98718 1 57410
2 98719 1 57410
2 98720 1 57435
2 98721 1 57435
2 98722 1 57474
2 98723 1 57474
2 98724 1 57493
2 98725 1 57493
2 98726 1 57546
2 98727 1 57546
2 98728 1 57593
2 98729 1 57593
2 98730 1 57633
2 98731 1 57633
2 98732 1 57638
2 98733 1 57638
2 98734 1 57639
2 98735 1 57639
2 98736 1 57723
2 98737 1 57723
2 98738 1 57724
2 98739 1 57724
2 98740 1 57728
2 98741 1 57728
2 98742 1 57728
2 98743 1 57870
2 98744 1 57870
2 98745 1 57946
2 98746 1 57946
2 98747 1 57970
2 98748 1 57970
2 98749 1 58009
2 98750 1 58009
2 98751 1 58010
2 98752 1 58010
2 98753 1 58074
2 98754 1 58074
2 98755 1 58074
2 98756 1 58074
2 98757 1 58093
2 98758 1 58093
2 98759 1 58187
2 98760 1 58187
2 98761 1 58420
2 98762 1 58420
2 98763 1 58464
2 98764 1 58464
2 98765 1 58554
2 98766 1 58554
2 98767 1 58568
2 98768 1 58568
2 98769 1 58662
2 98770 1 58662
2 98771 1 58814
2 98772 1 58814
2 98773 1 58815
2 98774 1 58815
2 98775 1 58837
2 98776 1 58837
2 98777 1 58978
2 98778 1 58978
2 98779 1 59014
2 98780 1 59014
2 98781 1 59028
2 98782 1 59028
2 98783 1 59039
2 98784 1 59039
2 98785 1 59042
2 98786 1 59042
2 98787 1 59099
2 98788 1 59099
2 98789 1 59099
2 98790 1 59123
2 98791 1 59123
0 27 5 177 1 25
0 28 5 229 1 59399
0 29 5 228 1 59724
0 30 5 211 1 60013
0 31 5 270 1 60184
0 32 5 225 1 60431
0 33 5 127 1 60645
0 34 5 8 1 60748
0 35 5 79 1 60752
0 36 5 162 1 60821
0 37 5 177 1 60968
0 38 5 257 1 61149
0 39 5 260 1 61376
0 40 5 182 1 61622
0 41 5 153 1 61835
0 42 5 14 1 61961
0 43 5 204 1 61966
0 44 5 240 1 62167
0 45 5 397 1 62414
0 46 5 391 1 62798
0 47 5 393 1 63252
0 48 5 236 1 63620
0 49 5 158 1 63884
0 50 5 64 1 64088
0 51 5 2 1 64194
0 52 7 6 2 60185 68188
0 53 7 31 2 65751 62168
0 54 5 65 1 69047
0 55 7 5 2 67400 69078
0 56 5 15 1 69143
0 57 7 57 2 60822 67160
0 58 5 66 1 69163
0 59 7 5 2 62415 69220
0 60 5 36 1 69286
0 61 7 4 2 66956 69291
0 62 5 2 1 69327
0 63 7 1 2 60753 69328
0 64 5 2 1 63
0 65 7 1 2 69148 69333
0 66 5 1 1 65
0 67 7 1 2 26 66
0 68 5 2 1 67
0 69 7 10 2 60754 67161
0 70 5 6 1 69337
0 71 7 1 2 65752 69347
0 72 5 3 1 71
0 73 7 26 2 65672 61967
0 74 5 57 1 69356
0 75 7 1 2 62169 69357
0 76 5 9 1 75
0 77 7 2 2 67401 69439
0 78 5 7 1 69448
0 79 7 1 2 69353 69449
0 80 5 1 1 79
0 81 7 1 2 69335 80
0 82 5 1 1 81
0 83 7 1 2 59400 82
0 84 5 1 1 83
0 85 7 11 2 60823 67402
0 86 5 6 1 69457
0 87 7 147 2 59236 60755
0 88 5 95 1 69474
0 89 7 15 2 66957 69475
0 90 5 10 1 69716
0 91 7 123 2 64197 65673
0 92 5 103 1 69741
0 93 7 7 2 67162 69864
0 94 5 26 1 69967
0 95 7 4 2 69731 69974
0 96 5 2 1 70000
0 97 7 1 2 69458 70004
0 98 5 1 1 97
0 99 7 1 2 84 98
0 100 5 1 1 99
0 101 7 92 2 64831 66090
0 102 5 123 1 70006
0 103 7 17 2 59725 70098
0 104 5 4 1 70221
0 105 7 6 2 60969 70099
0 106 5 2 1 70242
0 107 7 8 2 70238 70248
0 108 5 8 1 70250
0 109 7 1 2 100 70258
0 110 5 1 1 109
0 111 7 30 2 60756 66958
0 112 5 57 1 70266
0 113 7 1 2 70296 69221
0 114 5 1 1 113
0 115 7 3 2 69079 114
0 116 5 3 1 70353
0 117 7 1 2 59237 70354
0 118 5 2 1 117
0 119 7 3 2 60824 69382
0 120 5 20 1 70361
0 121 7 1 2 67163 70362
0 122 5 2 1 121
0 123 7 2 2 70359 70384
0 124 5 4 1 70386
0 125 7 9 2 67164 69383
0 126 5 11 1 70392
0 127 7 1 2 60825 69440
0 128 5 1 1 127
0 129 7 5 2 70401 128
0 130 5 1 1 70412
0 131 7 1 2 70297 69048
0 132 5 5 1 131
0 133 7 1 2 59238 70417
0 134 5 2 1 133
0 135 7 3 2 70413 70422
0 136 5 3 1 70424
0 137 7 1 2 59401 70427
0 138 5 2 1 137
0 139 7 4 2 70387 70430
0 140 5 2 1 70432
0 141 7 21 2 64198 64374
0 142 5 8 1 70438
0 143 7 38 2 61968 62170
0 144 5 41 1 70467
0 145 7 4 2 65674 70468
0 146 5 1 1 70546
0 147 7 2 2 70439 70547
0 148 5 1 1 70550
0 149 7 1 2 65753 70551
0 150 5 5 1 149
0 151 7 1 2 67403 70552
0 152 5 1 1 151
0 153 7 1 2 70433 152
0 154 5 1 1 153
0 155 7 158 2 60014 61150
0 156 5 166 1 70557
0 157 7 5 2 64603 70715
0 158 5 2 1 70881
0 159 7 3 2 65913 70716
0 160 5 2 1 70888
0 161 7 6 2 70886 70891
0 162 5 8 1 70893
0 163 7 9 2 70100 70894
0 164 5 3 1 70907
0 165 7 1 2 154 70908
0 166 5 1 1 165
0 167 7 10 2 64375 65914
0 168 5 4 1 70919
0 169 7 5 2 69742 70920
0 170 5 1 1 70933
0 171 7 14 2 65754 62416
0 172 5 3 1 70938
0 173 7 5 2 70469 70939
0 174 5 2 1 70955
0 175 7 1 2 70934 70956
0 176 5 2 1 175
0 177 7 1 2 59726 70962
0 178 5 2 1 177
0 179 7 14 2 64376 69743
0 180 5 10 1 70966
0 181 7 1 2 70967 70957
0 182 5 2 1 181
0 183 7 1 2 60970 70990
0 184 5 1 1 183
0 185 7 1 2 70964 184
0 186 5 1 1 185
0 187 7 1 2 70558 186
0 188 5 1 1 187
0 189 7 1 2 166 188
0 190 7 1 2 110 189
0 191 5 1 1 190
0 192 7 2 2 63885 191
0 193 7 1 2 69041 70992
0 194 5 1 1 193
0 195 7 1 2 69744 69149
0 196 5 3 1 195
0 197 7 1 2 70952 70994
0 198 5 1 1 197
0 199 7 2 2 68817 198
0 200 7 16 2 61969 63253
0 201 7 19 2 64832 65042
0 202 5 3 1 71015
0 203 7 104 2 64604 65915
0 204 5 129 1 71037
0 205 7 6 2 66091 71038
0 206 7 5 2 71016 71270
0 207 7 1 2 70999 71276
0 208 7 1 2 70997 207
0 209 5 1 1 208
0 210 7 1 2 194 209
0 211 5 1 1 210
0 212 7 1 2 66347 211
0 213 5 1 1 212
0 214 7 17 2 66959 69865
0 215 5 19 1 71281
0 216 7 12 2 69621 71298
0 217 5 10 1 71317
0 218 7 3 2 63254 71329
0 219 7 21 2 67165 67404
0 220 5 15 1 71342
0 221 7 4 2 61151 71343
0 222 7 2 2 71339 71378
0 223 7 16 2 60015 60186
0 224 5 2 1 71384
0 225 7 6 2 59402 71385
0 226 7 21 2 59727 60826
0 227 5 8 1 71408
0 228 7 7 2 60971 71409
0 229 5 1 1 71437
0 230 7 4 2 71402 71438
0 231 7 1 2 71382 71444
0 232 5 1 1 231
0 233 7 16 2 61970 69622
0 234 5 9 1 71448
0 235 7 39 2 69866 71464
0 236 7 15 2 60187 70101
0 237 5 61 1 71512
0 238 7 2 2 65916 69222
0 239 5 17 1 71588
0 240 7 1 2 71513 71590
0 241 5 1 1 240
0 242 7 16 2 60972 67166
0 243 5 9 1 71607
0 244 7 1 2 60827 71608
0 245 5 7 1 244
0 246 7 2 2 66092 71632
0 247 5 1 1 71639
0 248 7 1 2 64833 71640
0 249 5 1 1 248
0 250 7 1 2 60188 249
0 251 5 1 1 250
0 252 7 12 2 60828 61152
0 253 5 1 1 71641
0 254 7 3 2 71642 71609
0 255 5 1 1 71653
0 256 7 1 2 60016 71654
0 257 5 1 1 256
0 258 7 1 2 251 257
0 259 5 1 1 258
0 260 7 1 2 59728 259
0 261 5 1 1 260
0 262 7 1 2 241 261
0 263 5 1 1 262
0 264 7 1 2 59403 263
0 265 5 1 1 264
0 266 7 3 2 71514 71141
0 267 5 2 1 71656
0 268 7 1 2 69080 71657
0 269 5 1 1 268
0 270 7 1 2 265 269
0 271 5 1 1 270
0 272 7 1 2 67405 271
0 273 5 1 1 272
0 274 7 10 2 60189 67167
0 275 7 60 2 59404 60829
0 276 5 113 1 71671
0 277 7 3 2 71672 71142
0 278 5 2 1 71844
0 279 7 2 2 70102 71845
0 280 5 1 1 71849
0 281 7 2 2 70916 280
0 282 5 2 1 71851
0 283 7 1 2 71661 71853
0 284 5 2 1 283
0 285 7 1 2 273 71855
0 286 5 1 1 285
0 287 7 1 2 71473 286
0 288 5 1 1 287
0 289 7 46 2 60973 67406
0 290 5 39 1 71857
0 291 7 91 2 64377 65755
0 292 5 108 1 71942
0 293 7 3 2 60974 69867
0 294 5 6 1 72141
0 295 7 1 2 72033 72142
0 296 5 1 1 295
0 297 7 1 2 71903 296
0 298 5 1 1 297
0 299 7 1 2 59729 298
0 300 5 1 1 299
0 301 7 6 2 67168 72034
0 302 5 8 1 72150
0 303 7 9 2 71731 72156
0 304 5 22 1 72164
0 305 7 84 2 59730 60975
0 306 5 127 1 72195
0 307 7 11 2 67407 71143
0 308 5 7 1 72406
0 309 7 2 2 72279 72417
0 310 5 3 1 72424
0 311 7 1 2 72173 72426
0 312 5 1 1 311
0 313 7 1 2 300 312
0 314 5 2 1 313
0 315 7 1 2 70103 72429
0 316 5 1 1 315
0 317 7 9 2 65675 62171
0 318 5 3 1 72431
0 319 7 7 2 64199 72432
0 320 5 8 1 72443
0 321 7 2 2 72035 72450
0 322 5 4 1 72458
0 323 7 6 2 62417 71732
0 324 5 8 1 72464
0 325 7 2 2 72460 72465
0 326 5 1 1 72478
0 327 7 1 2 71039 72479
0 328 5 1 1 327
0 329 7 1 2 70559 328
0 330 5 1 1 329
0 331 7 1 2 316 330
0 332 5 1 1 331
0 333 7 1 2 60190 332
0 334 5 1 1 333
0 335 7 1 2 63255 334
0 336 7 1 2 288 335
0 337 5 1 1 336
0 338 7 3 2 70560 71144
0 339 5 30 1 72480
0 340 7 12 2 60830 69868
0 341 5 39 1 72513
0 342 7 12 2 59405 69869
0 343 5 34 1 72564
0 344 7 3 2 72525 72576
0 345 5 1 1 72610
0 346 7 6 2 64378 72280
0 347 5 3 1 72613
0 348 7 2 2 65756 72281
0 349 5 2 1 72622
0 350 7 4 2 72619 72624
0 351 5 6 1 72626
0 352 7 3 2 72611 72630
0 353 5 1 1 72636
0 354 7 1 2 71145 353
0 355 5 2 1 354
0 356 7 1 2 70717 72639
0 357 5 1 1 356
0 358 7 2 2 70104 357
0 359 5 1 1 72641
0 360 7 1 2 67169 72642
0 361 5 1 1 360
0 362 7 1 2 72483 361
0 363 5 1 1 362
0 364 7 1 2 65043 363
0 365 5 1 1 364
0 366 7 2 2 67170 71733
0 367 5 2 1 72643
0 368 7 3 2 65676 66960
0 369 5 1 1 72647
0 370 7 5 2 64200 72648
0 371 5 4 1 72650
0 372 7 1 2 72645 72655
0 373 5 5 1 372
0 374 7 14 2 60017 71146
0 375 5 50 1 72664
0 376 7 1 2 72659 72678
0 377 5 2 1 376
0 378 7 1 2 70968 71040
0 379 5 3 1 378
0 380 7 2 2 62172 72730
0 381 5 1 1 72733
0 382 7 9 2 59406 60018
0 383 5 1 1 72735
0 384 7 1 2 67171 383
0 385 5 2 1 384
0 386 7 1 2 72656 72744
0 387 7 1 2 381 386
0 388 5 1 1 387
0 389 7 1 2 66093 388
0 390 5 1 1 389
0 391 7 1 2 72728 390
0 392 5 1 1 391
0 393 7 1 2 60191 392
0 394 5 1 1 393
0 395 7 5 2 60019 65044
0 396 7 5 2 61153 72746
0 397 5 2 1 72751
0 398 7 16 2 65757 61971
0 399 5 9 1 72758
0 400 7 6 2 65677 72759
0 401 5 5 1 72783
0 402 7 3 2 72784 70440
0 403 5 4 1 72794
0 404 7 1 2 72752 72797
0 405 5 1 1 404
0 406 7 6 2 60020 66094
0 407 5 1 1 72801
0 408 7 2 2 62173 72802
0 409 5 1 1 72807
0 410 7 12 2 65045 61154
0 411 5 3 1 72809
0 412 7 1 2 409 72821
0 413 5 1 1 412
0 414 7 3 2 65758 70298
0 415 5 12 1 72824
0 416 7 2 2 59239 72827
0 417 5 2 1 72839
0 418 7 8 2 72841 70364
0 419 5 7 1 72843
0 420 7 9 2 59240 60831
0 421 5 3 1 72858
0 422 7 3 2 70267 72859
0 423 5 8 1 72870
0 424 7 1 2 64379 72873
0 425 5 2 1 424
0 426 7 3 2 72851 72881
0 427 5 1 1 72883
0 428 7 1 2 72884 71147
0 429 5 1 1 428
0 430 7 1 2 72196 72798
0 431 5 1 1 430
0 432 7 1 2 429 431
0 433 5 1 1 432
0 434 7 1 2 413 433
0 435 5 1 1 434
0 436 7 1 2 405 435
0 437 7 1 2 394 436
0 438 7 1 2 365 437
0 439 5 1 1 438
0 440 7 1 2 67408 439
0 441 5 1 1 440
0 442 7 6 2 64834 72282
0 443 5 45 1 72886
0 444 7 1 2 70436 72892
0 445 5 1 1 444
0 446 7 20 2 60021 60976
0 447 7 5 2 59731 72937
0 448 5 8 1 72957
0 449 7 3 2 65046 72962
0 450 5 17 1 72970
0 451 7 1 2 60022 70553
0 452 5 1 1 451
0 453 7 36 2 66961 67172
0 454 5 29 1 72990
0 455 7 3 2 59241 72991
0 456 5 1 1 73055
0 457 7 5 2 60757 60832
0 458 5 3 1 73058
0 459 7 3 2 59407 73059
0 460 5 2 1 73066
0 461 7 1 2 73056 73067
0 462 5 3 1 461
0 463 7 1 2 452 73071
0 464 5 1 1 463
0 465 7 1 2 71148 464
0 466 5 1 1 465
0 467 7 1 2 72971 466
0 468 7 1 2 445 467
0 469 5 1 1 468
0 470 7 4 2 62174 71041
0 471 5 1 1 73074
0 472 7 43 2 64380 62175
0 473 5 19 1 73078
0 474 7 4 2 72526 73079
0 475 5 2 1 73140
0 476 7 2 2 71149 73144
0 477 5 1 1 73146
0 478 7 1 2 62418 477
0 479 5 1 1 478
0 480 7 2 2 471 479
0 481 5 1 1 73148
0 482 7 1 2 60192 73149
0 483 5 1 1 482
0 484 7 1 2 61155 483
0 485 7 1 2 469 484
0 486 5 1 1 485
0 487 7 22 2 66095 62419
0 488 5 11 1 73150
0 489 7 16 2 59242 70268
0 490 5 22 1 73183
0 491 7 11 2 61972 69745
0 492 5 5 1 73221
0 493 7 4 2 59408 73232
0 494 5 4 1 73237
0 495 7 9 2 73199 73241
0 496 5 8 1 73245
0 497 7 3 2 60193 71150
0 498 5 2 1 73262
0 499 7 1 2 73246 73265
0 500 5 1 1 499
0 501 7 1 2 69081 72973
0 502 7 1 2 500 501
0 503 5 1 1 502
0 504 7 2 2 64381 69358
0 505 5 2 1 73267
0 506 7 5 2 59732 73269
0 507 5 7 1 73271
0 508 7 7 2 59409 70269
0 509 5 4 1 73283
0 510 7 4 2 64605 73290
0 511 5 7 1 73294
0 512 7 1 2 59243 73298
0 513 5 4 1 512
0 514 7 3 2 73276 73305
0 515 5 3 1 73309
0 516 7 12 2 60833 60977
0 517 7 12 2 67173 73315
0 518 7 1 2 60023 73327
0 519 5 1 1 518
0 520 7 1 2 65047 519
0 521 5 2 1 520
0 522 7 1 2 73312 73339
0 523 5 1 1 522
0 524 7 13 2 64382 61973
0 525 5 19 1 73341
0 526 7 5 2 69746 73342
0 527 5 10 1 73373
0 528 7 2 2 60194 73378
0 529 5 2 1 73388
0 530 7 31 2 59733 60024
0 531 5 5 1 73392
0 532 7 12 2 59410 60758
0 533 5 2 1 73428
0 534 7 11 2 59244 66962
0 535 5 2 1 73442
0 536 7 4 2 73429 73443
0 537 5 5 1 73455
0 538 7 1 2 73393 73456
0 539 5 1 1 538
0 540 7 1 2 73390 539
0 541 5 1 1 540
0 542 7 1 2 71591 541
0 543 5 1 1 542
0 544 7 7 2 60195 60978
0 545 7 1 2 59734 73464
0 546 5 1 1 545
0 547 7 1 2 543 546
0 548 7 1 2 523 547
0 549 7 1 2 503 548
0 550 5 1 1 549
0 551 7 1 2 73151 550
0 552 5 1 1 551
0 553 7 1 2 68189 552
0 554 7 1 2 486 553
0 555 7 1 2 441 554
0 556 5 1 1 555
0 557 7 1 2 61377 556
0 558 7 1 2 337 557
0 559 5 1 1 558
0 560 7 1 2 232 559
0 561 5 1 1 560
0 562 7 1 2 63886 561
0 563 5 1 1 562
0 564 7 1 2 213 563
0 565 5 1 1 564
0 566 7 1 2 62799 565
0 567 5 1 1 566
0 568 7 21 2 67797 63887
0 569 7 4 2 70007 72283
0 570 5 17 1 73492
0 571 7 19 2 62176 71734
0 572 5 6 1 73513
0 573 7 2 2 59735 73532
0 574 5 1 1 73538
0 575 7 1 2 71858 574
0 576 5 1 1 575
0 577 7 2 2 60025 65917
0 578 5 4 1 73540
0 579 7 7 2 59736 72036
0 580 5 29 1 73546
0 581 7 3 2 64835 73553
0 582 5 3 1 73582
0 583 7 1 2 62420 73585
0 584 5 1 1 583
0 585 7 1 2 73542 584
0 586 7 1 2 576 585
0 587 5 1 1 586
0 588 7 1 2 61156 587
0 589 5 1 1 588
0 590 7 5 2 59411 62421
0 591 7 1 2 69164 73588
0 592 5 3 1 591
0 593 7 24 2 62177 67409
0 594 5 7 1 73596
0 595 7 4 2 61974 73597
0 596 5 1 1 73627
0 597 7 1 2 62422 72174
0 598 5 2 1 597
0 599 7 1 2 596 73631
0 600 5 1 1 599
0 601 7 1 2 69476 600
0 602 5 1 1 601
0 603 7 1 2 73593 602
0 604 7 1 2 589 603
0 605 5 1 1 604
0 606 7 1 2 73496 605
0 607 5 1 1 606
0 608 7 2 2 62423 70105
0 609 5 4 1 73633
0 610 7 6 2 59245 69338
0 611 5 3 1 73639
0 612 7 1 2 71735 73645
0 613 5 5 1 612
0 614 7 20 2 61157 67174
0 615 5 5 1 73653
0 616 7 2 2 72037 73673
0 617 7 12 2 66963 62178
0 618 5 3 1 73680
0 619 7 1 2 67410 73692
0 620 7 1 2 73678 619
0 621 7 1 2 73648 620
0 622 5 1 1 621
0 623 7 1 2 73635 622
0 624 5 1 1 623
0 625 7 5 2 62179 69623
0 626 5 19 1 73695
0 627 7 1 2 71151 73700
0 628 7 1 2 624 627
0 629 5 1 1 628
0 630 7 3 2 60026 62424
0 631 5 4 1 73719
0 632 7 7 2 60979 66096
0 633 7 2 2 67411 73726
0 634 5 1 1 73733
0 635 7 1 2 73722 634
0 636 5 1 1 635
0 637 7 1 2 72038 636
0 638 5 1 1 637
0 639 7 11 2 66097 67412
0 640 5 6 1 73735
0 641 7 2 2 71610 73736
0 642 5 1 1 73752
0 643 7 1 2 638 642
0 644 5 1 1 643
0 645 7 1 2 59737 644
0 646 5 1 1 645
0 647 7 10 2 60027 67413
0 648 5 2 1 73754
0 649 7 5 2 66098 67175
0 650 5 3 1 73766
0 651 7 1 2 73755 73767
0 652 5 1 1 651
0 653 7 28 2 65918 62425
0 654 5 32 1 73774
0 655 7 1 2 60028 73802
0 656 5 10 1 655
0 657 7 2 2 61158 73803
0 658 5 9 1 73844
0 659 7 2 2 73834 73846
0 660 5 1 1 73855
0 661 7 27 2 64383 64606
0 662 5 2 1 73857
0 663 7 12 2 65759 73858
0 664 5 1 1 73886
0 665 7 21 2 61159 67414
0 666 5 2 1 73898
0 667 7 5 2 60980 73899
0 668 5 4 1 73921
0 669 7 1 2 664 73926
0 670 7 1 2 660 669
0 671 5 1 1 670
0 672 7 1 2 652 671
0 673 7 1 2 646 672
0 674 7 1 2 629 673
0 675 7 1 2 607 674
0 676 5 1 1 675
0 677 7 1 2 68190 676
0 678 5 1 1 677
0 679 7 1 2 71736 72679
0 680 5 2 1 679
0 681 7 4 2 72893 73930
0 682 5 1 1 73932
0 683 7 1 2 69477 73933
0 684 5 1 1 683
0 685 7 2 2 60029 72039
0 686 5 2 1 73936
0 687 7 2 2 73937 71152
0 688 5 1 1 73940
0 689 7 1 2 684 688
0 690 5 1 1 689
0 691 7 1 2 67176 690
0 692 5 1 1 691
0 693 7 1 2 72963 692
0 694 5 1 1 693
0 695 7 15 2 67415 63256
0 696 7 7 2 66964 73942
0 697 5 2 1 73957
0 698 7 1 2 61160 73958
0 699 7 1 2 694 698
0 700 5 1 1 699
0 701 7 1 2 678 700
0 702 5 1 1 701
0 703 7 1 2 65048 702
0 704 5 1 1 703
0 705 7 8 2 60030 63257
0 706 7 4 2 60981 69082
0 707 5 6 1 73974
0 708 7 1 2 59412 71592
0 709 5 2 1 708
0 710 7 5 2 73978 73984
0 711 5 4 1 73986
0 712 7 1 2 59738 73991
0 713 5 1 1 712
0 714 7 8 2 59413 67177
0 715 5 36 1 73995
0 716 7 9 2 60834 73996
0 717 5 32 1 74039
0 718 7 3 2 60982 74040
0 719 5 1 1 74080
0 720 7 1 2 713 719
0 721 5 1 1 720
0 722 7 24 2 66965 67416
0 723 5 20 1 74083
0 724 7 7 2 62426 69624
0 725 5 8 1 74127
0 726 7 1 2 74107 74134
0 727 7 1 2 721 726
0 728 5 1 1 727
0 729 7 14 2 59739 62427
0 730 5 2 1 74142
0 731 7 2 2 64384 69223
0 732 5 5 1 74158
0 733 7 2 2 74160 73975
0 734 5 2 1 74165
0 735 7 1 2 74143 74166
0 736 5 1 1 735
0 737 7 2 2 72040 69478
0 738 5 4 1 74169
0 739 7 3 2 71737 74171
0 740 5 12 1 74175
0 741 7 2 2 66966 71153
0 742 7 2 2 74178 74190
0 743 5 1 1 74192
0 744 7 1 2 73598 74193
0 745 5 1 1 744
0 746 7 1 2 736 745
0 747 7 1 2 728 746
0 748 5 1 1 747
0 749 7 1 2 61161 748
0 750 5 1 1 749
0 751 7 14 2 59740 71673
0 752 5 4 1 74194
0 753 7 1 2 74195 69717
0 754 7 1 2 73753 753
0 755 5 1 1 754
0 756 7 1 2 750 755
0 757 5 1 1 756
0 758 7 1 2 73966 757
0 759 5 1 1 758
0 760 7 16 2 61975 68191
0 761 7 5 2 62428 72484
0 762 7 2 2 73080 74228
0 763 5 2 1 74233
0 764 7 1 2 60196 74234
0 765 5 1 1 764
0 766 7 3 2 71042 73900
0 767 7 2 2 64836 74237
0 768 5 1 1 74240
0 769 7 1 2 67178 74241
0 770 5 1 1 769
0 771 7 2 2 765 770
0 772 5 1 1 74242
0 773 7 7 2 65049 67417
0 774 5 2 1 74244
0 775 7 2 2 73654 74245
0 776 5 1 1 74253
0 777 7 1 2 74243 776
0 778 5 1 1 777
0 779 7 1 2 74212 778
0 780 5 1 1 779
0 781 7 3 2 61162 73943
0 782 7 8 2 60197 66967
0 783 5 2 1 74258
0 784 7 1 2 74255 74259
0 785 5 1 1 784
0 786 7 1 2 780 785
0 787 5 1 1 786
0 788 7 1 2 72527 787
0 789 5 1 1 788
0 790 7 1 2 759 789
0 791 7 1 2 704 790
0 792 5 1 1 791
0 793 7 1 2 61378 792
0 794 5 1 1 793
0 795 7 1 2 66968 69625
0 796 5 2 1 795
0 797 7 15 2 61976 67179
0 798 5 3 1 74270
0 799 7 2 2 73693 74285
0 800 5 4 1 74288
0 801 7 2 2 69870 74290
0 802 5 1 1 74294
0 803 7 5 2 74268 74295
0 804 7 1 2 72041 74296
0 805 5 1 1 804
0 806 7 2 2 61977 69871
0 807 5 1 1 74301
0 808 7 7 2 70505 73026
0 809 5 2 1 74303
0 810 7 1 2 807 74310
0 811 5 4 1 810
0 812 7 1 2 71674 74312
0 813 5 1 1 812
0 814 7 1 2 805 813
0 815 5 2 1 814
0 816 7 3 2 66348 70718
0 817 5 7 1 74318
0 818 7 1 2 74316 74321
0 819 5 1 1 818
0 820 7 19 2 61163 66349
0 821 5 1 1 74328
0 822 7 4 2 60031 74329
0 823 5 4 1 74347
0 824 7 18 2 66099 61379
0 825 5 2 1 74355
0 826 7 1 2 74351 74373
0 827 5 2 1 826
0 828 7 2 2 66969 74375
0 829 7 1 2 72151 74377
0 830 5 1 1 829
0 831 7 1 2 819 830
0 832 5 1 1 831
0 833 7 1 2 67418 832
0 834 5 1 1 833
0 835 7 5 2 61978 70106
0 836 5 3 1 74379
0 837 7 19 2 67180 62429
0 838 5 3 1 74387
0 839 7 4 2 59414 71465
0 840 5 4 1 74409
0 841 7 5 2 74410 72514
0 842 5 3 1 74417
0 843 7 1 2 74388 74418
0 844 5 3 1 843
0 845 7 1 2 74384 74425
0 846 5 1 1 845
0 847 7 1 2 61380 846
0 848 5 1 1 847
0 849 7 5 2 64201 70299
0 850 5 5 1 74428
0 851 7 2 2 67181 74433
0 852 5 1 1 74438
0 853 7 2 2 69384 70561
0 854 5 2 1 74440
0 855 7 3 2 62430 71675
0 856 7 1 2 74441 74444
0 857 7 1 2 74439 856
0 858 5 1 1 857
0 859 7 1 2 848 858
0 860 7 1 2 834 859
0 861 5 1 1 860
0 862 7 1 2 71154 861
0 863 5 1 1 862
0 864 7 10 2 64385 69049
0 865 5 4 1 74447
0 866 7 7 2 69747 74448
0 867 5 6 1 74461
0 868 7 13 2 61979 67419
0 869 5 1 1 74474
0 870 7 1 2 74468 74475
0 871 5 1 1 870
0 872 7 2 2 59415 69083
0 873 5 6 1 74487
0 874 7 9 2 69224 74489
0 875 5 1 1 74495
0 876 7 9 2 62180 71943
0 877 5 11 1 74504
0 878 7 1 2 74513 71474
0 879 5 1 1 878
0 880 7 2 2 74496 879
0 881 5 2 1 74524
0 882 7 1 2 62431 74526
0 883 5 1 1 882
0 884 7 1 2 871 883
0 885 5 1 1 884
0 886 7 1 2 74322 885
0 887 5 1 1 886
0 888 7 1 2 67420 74378
0 889 5 1 1 888
0 890 7 1 2 887 889
0 891 5 1 1 890
0 892 7 1 2 72197 891
0 893 5 1 1 892
0 894 7 3 2 71299 74128
0 895 5 5 1 74528
0 896 7 1 2 74108 74514
0 897 7 1 2 74531 896
0 898 5 1 1 897
0 899 7 1 2 72042 74389
0 900 5 1 1 899
0 901 7 3 2 67421 69872
0 902 5 4 1 74536
0 903 7 1 2 61980 74537
0 904 5 1 1 903
0 905 7 1 2 900 904
0 906 7 1 2 898 905
0 907 5 1 1 906
0 908 7 1 2 61381 907
0 909 5 1 1 908
0 910 7 6 2 69479 74196
0 911 5 2 1 74543
0 912 7 3 2 66350 72992
0 913 5 2 1 74551
0 914 7 1 2 71859 74552
0 915 7 1 2 74544 914
0 916 5 1 1 915
0 917 7 1 2 909 916
0 918 5 1 1 917
0 919 7 1 2 70107 918
0 920 5 1 1 919
0 921 7 15 2 64607 71738
0 922 5 39 1 74556
0 923 7 4 2 65919 74557
0 924 5 15 1 74610
0 925 7 7 2 69339 73444
0 926 5 7 1 74629
0 927 7 2 2 67422 74630
0 928 5 2 1 74643
0 929 7 1 2 74376 74644
0 930 5 1 1 929
0 931 7 8 2 61382 70108
0 932 5 7 1 74647
0 933 7 1 2 62432 74648
0 934 5 1 1 933
0 935 7 1 2 930 934
0 936 5 1 1 935
0 937 7 1 2 74614 936
0 938 5 1 1 937
0 939 7 4 2 59416 74084
0 940 5 3 1 74662
0 941 7 17 2 61164 61383
0 942 5 3 1 74669
0 943 7 1 2 64837 74109
0 944 5 2 1 943
0 945 7 1 2 74670 74689
0 946 7 1 2 74666 945
0 947 5 1 1 946
0 948 7 1 2 63258 947
0 949 7 1 2 938 948
0 950 7 1 2 920 949
0 951 7 1 2 893 950
0 952 7 1 2 863 951
0 953 5 1 1 952
0 954 7 1 2 73640 73497
0 955 5 1 1 954
0 956 7 1 2 70239 955
0 957 5 1 1 956
0 958 7 1 2 72043 957
0 959 5 1 1 958
0 960 7 1 2 71676 73498
0 961 5 1 1 960
0 962 7 1 2 70251 961
0 963 5 5 1 962
0 964 7 1 2 73701 74691
0 965 5 1 1 964
0 966 7 1 2 70719 965
0 967 7 1 2 959 966
0 968 5 1 1 967
0 969 7 1 2 62433 968
0 970 5 1 1 969
0 971 7 1 2 65920 73901
0 972 5 2 1 971
0 973 7 1 2 72175 73499
0 974 5 1 1 973
0 975 7 1 2 70252 974
0 976 5 1 1 975
0 977 7 1 2 62434 976
0 978 5 1 1 977
0 979 7 1 2 74696 978
0 980 5 1 1 979
0 981 7 1 2 71282 980
0 982 5 1 1 981
0 983 7 7 2 65921 61165
0 984 7 1 2 60032 74698
0 985 5 2 1 984
0 986 7 8 2 64608 71944
0 987 5 4 1 74707
0 988 7 1 2 62435 70243
0 989 5 1 1 988
0 990 7 1 2 74697 989
0 991 5 1 1 990
0 992 7 1 2 74715 991
0 993 5 1 1 992
0 994 7 1 2 74705 993
0 995 7 1 2 982 994
0 996 7 1 2 970 995
0 997 5 1 1 996
0 998 7 1 2 66351 997
0 999 5 1 1 998
0 1000 7 22 2 66352 67423
0 1001 5 5 1 74719
0 1002 7 3 2 71155 74179
0 1003 5 2 1 74746
0 1004 7 1 2 72887 74749
0 1005 5 1 1 1004
0 1006 7 1 2 67182 1005
0 1007 5 1 1 1006
0 1008 7 4 2 60983 72044
0 1009 5 6 1 74751
0 1010 7 4 2 73554 74755
0 1011 5 7 1 74761
0 1012 7 2 2 73533 74765
0 1013 7 1 2 71283 74772
0 1014 5 1 1 1013
0 1015 7 1 2 71945 71300
0 1016 5 5 1 1015
0 1017 7 1 2 72894 74774
0 1018 5 1 1 1017
0 1019 7 1 2 73423 1018
0 1020 7 1 2 1014 1019
0 1021 7 1 2 1007 1020
0 1022 5 1 1 1021
0 1023 7 1 2 74720 1022
0 1024 5 1 1 1023
0 1025 7 10 2 64202 69359
0 1026 5 19 1 74779
0 1027 7 1 2 74789 73121
0 1028 5 4 1 1027
0 1029 7 1 2 61384 72680
0 1030 7 1 2 74808 1029
0 1031 5 1 1 1030
0 1032 7 1 2 1024 1031
0 1033 5 1 1 1032
0 1034 7 1 2 66100 1033
0 1035 5 1 1 1034
0 1036 7 8 2 60984 61166
0 1037 5 3 1 74812
0 1038 7 1 2 71739 74813
0 1039 5 1 1 1038
0 1040 7 8 2 61981 69480
0 1041 5 2 1 74823
0 1042 7 1 2 71847 73493
0 1043 5 1 1 1042
0 1044 7 1 2 74824 1043
0 1045 5 1 1 1044
0 1046 7 1 2 1039 1045
0 1047 5 1 1 1046
0 1048 7 1 2 74721 1047
0 1049 5 1 1 1048
0 1050 7 7 2 64838 73859
0 1051 5 3 1 74833
0 1052 7 8 2 65922 61385
0 1053 7 2 2 74834 74843
0 1054 5 1 1 74851
0 1055 7 1 2 1049 1054
0 1056 5 1 1 1055
0 1057 7 1 2 62181 1056
0 1058 5 1 1 1057
0 1059 7 3 2 64839 61386
0 1060 7 1 2 74853 73775
0 1061 5 2 1 1060
0 1062 7 12 2 60985 66353
0 1063 7 2 2 73902 74858
0 1064 5 2 1 74870
0 1065 7 1 2 74856 74872
0 1066 5 1 1 1065
0 1067 7 1 2 64609 1066
0 1068 5 1 1 1067
0 1069 7 1 2 68192 1068
0 1070 7 1 2 1058 1069
0 1071 7 1 2 1035 1070
0 1072 7 1 2 999 1071
0 1073 5 1 1 1072
0 1074 7 1 2 60198 1073
0 1075 7 1 2 953 1074
0 1076 5 1 1 1075
0 1077 7 1 2 74156 73746
0 1078 5 2 1 1077
0 1079 7 1 2 64840 71633
0 1080 5 1 1 1079
0 1081 7 1 2 74874 1080
0 1082 5 1 1 1081
0 1083 7 11 2 64610 62436
0 1084 5 15 1 74876
0 1085 7 3 2 61167 74887
0 1086 5 1 1 74902
0 1087 7 1 2 71904 74903
0 1088 5 1 1 1087
0 1089 7 1 2 1082 1088
0 1090 5 1 1 1089
0 1091 7 1 2 61387 1090
0 1092 5 1 1 1091
0 1093 7 5 2 60033 73655
0 1094 5 3 1 74905
0 1095 7 7 2 60835 66354
0 1096 5 2 1 74913
0 1097 7 1 2 71860 74914
0 1098 7 1 2 74906 1097
0 1099 5 1 1 1098
0 1100 7 1 2 1092 1099
0 1101 5 1 1 1100
0 1102 7 1 2 65050 1101
0 1103 5 1 1 1102
0 1104 7 17 2 66355 62437
0 1105 5 1 1 74922
0 1106 7 2 2 74907 71439
0 1107 7 1 2 74923 74939
0 1108 5 1 1 1107
0 1109 7 1 2 1103 1108
0 1110 5 1 1 1109
0 1111 7 1 2 68193 1110
0 1112 5 1 1 1111
0 1113 7 11 2 60986 61388
0 1114 5 2 1 74941
0 1115 7 3 2 60836 74942
0 1116 7 5 2 63259 74390
0 1117 7 8 2 59417 61168
0 1118 7 9 2 60034 74962
0 1119 5 2 1 74970
0 1120 7 1 2 74957 74971
0 1121 7 1 2 74954 1120
0 1122 5 1 1 1121
0 1123 7 1 2 1112 1122
0 1124 5 1 1 1123
0 1125 7 1 2 66970 1124
0 1126 5 1 1 1125
0 1127 7 16 2 61169 63260
0 1128 7 6 2 60035 74981
0 1129 5 3 1 74997
0 1130 7 27 2 59418 66971
0 1131 5 10 1 75006
0 1132 7 1 2 62438 75033
0 1133 5 14 1 1132
0 1134 7 2 2 74998 75043
0 1135 5 1 1 75057
0 1136 7 1 2 74110 75058
0 1137 5 1 1 1136
0 1138 7 20 2 65051 68194
0 1139 7 4 2 66101 74085
0 1140 7 1 2 75059 75079
0 1141 5 1 1 1140
0 1142 7 1 2 1137 1141
0 1143 5 1 1 1142
0 1144 7 1 2 59741 1143
0 1145 5 1 1 1144
0 1146 7 3 2 68195 70109
0 1147 5 3 1 75083
0 1148 7 13 2 66972 62439
0 1149 7 1 2 65052 75089
0 1150 7 1 2 75084 1149
0 1151 5 1 1 1150
0 1152 7 1 2 1145 1151
0 1153 5 1 1 1152
0 1154 7 1 2 61389 1153
0 1155 5 1 1 1154
0 1156 7 22 2 66973 68196
0 1157 5 6 1 75102
0 1158 7 2 2 75103 74722
0 1159 5 1 1 75130
0 1160 7 1 2 59742 72753
0 1161 7 1 2 75131 1160
0 1162 5 1 1 1161
0 1163 7 1 2 1155 1162
0 1164 5 1 1 1163
0 1165 7 1 2 71593 1164
0 1166 5 1 1 1165
0 1167 7 14 2 65053 61390
0 1168 5 8 1 75132
0 1169 7 2 2 66102 75104
0 1170 7 1 2 75133 75154
0 1171 5 1 1 1170
0 1172 7 88 2 65054 66356
0 1173 5 139 1 75156
0 1174 7 20 2 68197 75244
0 1175 5 4 1 75383
0 1176 7 17 2 66357 61982
0 1177 5 5 1 75407
0 1178 7 19 2 66974 63261
0 1179 5 1 1 75429
0 1180 7 4 2 75424 1179
0 1181 5 1 1 75448
0 1182 7 1 2 75449 70562
0 1183 7 1 2 75403 1182
0 1184 5 1 1 1183
0 1185 7 1 2 1171 1184
0 1186 5 1 1 1185
0 1187 7 1 2 72407 1186
0 1188 5 1 1 1187
0 1189 7 2 2 61391 73500
0 1190 5 1 1 75452
0 1191 7 3 2 70563 72198
0 1192 5 5 1 75454
0 1193 7 1 2 1190 75457
0 1194 5 1 1 1193
0 1195 7 76 2 60199 61392
0 1196 5 125 1 75462
0 1197 7 9 2 68198 75538
0 1198 7 1 2 75090 75663
0 1199 7 1 2 1194 1198
0 1200 5 1 1 1199
0 1201 7 1 2 1188 1200
0 1202 5 1 1 1201
0 1203 7 1 2 59419 1202
0 1204 5 1 1 1203
0 1205 7 25 2 62440 63262
0 1206 5 4 1 75672
0 1207 7 18 2 61170 66975
0 1208 5 3 1 75701
0 1209 7 5 2 59743 61393
0 1210 7 2 2 75722 72938
0 1211 5 1 1 75727
0 1212 7 2 2 75702 75728
0 1213 7 1 2 75673 75729
0 1214 5 1 1 1213
0 1215 7 1 2 1204 1214
0 1216 5 1 1 1215
0 1217 7 1 2 69084 1216
0 1218 5 1 1 1217
0 1219 7 3 2 61394 73944
0 1220 7 9 2 61171 61983
0 1221 7 4 2 60036 75734
0 1222 7 9 2 60987 69165
0 1223 5 5 1 75747
0 1224 7 1 2 75743 75748
0 1225 7 1 2 75731 1224
0 1226 5 1 1 1225
0 1227 7 1 2 1218 1226
0 1228 7 1 2 1166 1227
0 1229 7 1 2 1126 1228
0 1230 5 1 1 1229
0 1231 7 1 2 69873 1230
0 1232 5 1 1 1231
0 1233 7 1 2 69481 70470
0 1234 5 2 1 1233
0 1235 7 4 2 65055 67183
0 1236 5 3 1 75763
0 1237 7 1 2 75761 75767
0 1238 5 1 1 1237
0 1239 7 3 2 71156 72620
0 1240 5 1 1 75770
0 1241 7 7 2 72625 75771
0 1242 7 1 2 1238 75773
0 1243 5 1 1 1242
0 1244 7 9 2 67184 69482
0 1245 5 4 1 75780
0 1246 7 1 2 75789 72284
0 1247 5 1 1 1246
0 1248 7 1 2 65056 74766
0 1249 7 1 2 1247 1248
0 1250 5 1 1 1249
0 1251 7 1 2 1243 1250
0 1252 5 1 1 1251
0 1253 7 1 2 67424 1252
0 1254 5 1 1 1253
0 1255 7 2 2 62441 72199
0 1256 7 6 2 59420 69166
0 1257 5 7 1 75795
0 1258 7 3 2 69626 75801
0 1259 5 3 1 75808
0 1260 7 5 2 72176 75811
0 1261 5 1 1 75814
0 1262 7 1 2 75793 75815
0 1263 5 1 1 1262
0 1264 7 1 2 1254 1263
0 1265 5 1 1 1264
0 1266 7 38 2 66358 68199
0 1267 5 2 1 75819
0 1268 7 3 2 60037 75820
0 1269 5 4 1 75859
0 1270 7 1 2 61172 75860
0 1271 7 1 2 1265 1270
0 1272 5 1 1 1271
0 1273 7 2 2 72528 74213
0 1274 7 17 2 60200 66359
0 1275 5 5 1 75868
0 1276 7 1 2 75869 71379
0 1277 7 1 2 75866 1276
0 1278 5 1 1 1277
0 1279 7 1 2 1272 1278
0 1280 7 1 2 1232 1279
0 1281 7 1 2 1076 1280
0 1282 7 1 2 794 1281
0 1283 5 1 1 1282
0 1284 7 1 2 73471 1283
0 1285 5 1 1 1284
0 1286 7 1 2 567 1285
0 1287 5 1 1 1286
0 1288 7 1 2 63621 1287
0 1289 5 1 1 1288
0 1290 7 2 2 60759 69167
0 1291 5 2 1 75890
0 1292 7 1 2 70360 75892
0 1293 5 1 1 1292
0 1294 7 1 2 71157 1293
0 1295 5 1 1 1294
0 1296 7 18 2 65678 65760
0 1297 5 2 1 75894
0 1298 7 12 2 64203 75895
0 1299 5 6 1 75914
0 1300 7 1 2 75926 72200
0 1301 5 3 1 1300
0 1302 7 1 2 1295 75932
0 1303 5 1 1 1302
0 1304 7 1 2 59421 1303
0 1305 5 1 1 1304
0 1306 7 9 2 66976 73702
0 1307 5 2 1 75935
0 1308 7 1 2 72529 69975
0 1309 7 1 2 75944 1308
0 1310 5 1 1 1309
0 1311 7 1 2 72201 1310
0 1312 5 1 1 1311
0 1313 7 1 2 1305 1312
0 1314 5 1 1 1313
0 1315 7 1 2 70110 1314
0 1316 5 1 1 1315
0 1317 7 3 2 71740 75945
0 1318 5 2 1 75946
0 1319 7 6 2 65761 73081
0 1320 5 14 1 75951
0 1321 7 1 2 69874 75957
0 1322 5 4 1 1321
0 1323 7 1 2 71043 75971
0 1324 7 1 2 75947 1323
0 1325 5 1 1 1324
0 1326 7 1 2 70564 1325
0 1327 5 1 1 1326
0 1328 7 1 2 1316 1327
0 1329 5 1 1 1328
0 1330 7 1 2 67425 1329
0 1331 5 1 1 1330
0 1332 7 2 2 65057 75458
0 1333 5 1 1 75975
0 1334 7 1 2 1331 75976
0 1335 5 1 1 1334
0 1336 7 5 2 69748 71741
0 1337 5 3 1 75977
0 1338 7 3 2 67426 75978
0 1339 5 1 1 75985
0 1340 7 2 2 65923 74172
0 1341 5 1 1 75988
0 1342 7 1 2 74558 75989
0 1343 5 2 1 1342
0 1344 7 1 2 62442 75990
0 1345 5 1 1 1344
0 1346 7 1 2 1339 1345
0 1347 5 1 1 1346
0 1348 7 1 2 66977 1347
0 1349 5 1 1 1348
0 1350 7 9 2 67427 72045
0 1351 5 13 1 75992
0 1352 7 1 2 65924 75993
0 1353 5 1 1 1352
0 1354 7 1 2 71044 72466
0 1355 5 1 1 1354
0 1356 7 1 2 69875 71905
0 1357 7 1 2 1355 1356
0 1358 5 1 1 1357
0 1359 7 1 2 1353 1358
0 1360 7 1 2 1349 1359
0 1361 5 1 1 1360
0 1362 7 1 2 66103 1361
0 1363 5 1 1 1362
0 1364 7 5 2 64841 66978
0 1365 5 4 1 76014
0 1366 7 1 2 76015 75986
0 1367 5 1 1 1366
0 1368 7 1 2 1363 1367
0 1369 5 1 1 1368
0 1370 7 1 2 67185 1369
0 1371 5 1 1 1370
0 1372 7 3 2 62443 71158
0 1373 5 3 1 76023
0 1374 7 1 2 59246 76024
0 1375 5 1 1 1374
0 1376 7 3 2 59422 72860
0 1377 5 3 1 76029
0 1378 7 1 2 76001 76032
0 1379 5 1 1 1378
0 1380 7 1 2 71906 1379
0 1381 5 1 1 1380
0 1382 7 1 2 1375 1381
0 1383 5 2 1 1382
0 1384 7 1 2 69385 76035
0 1385 5 1 1 1384
0 1386 7 4 2 64386 70300
0 1387 5 23 1 76037
0 1388 7 2 2 65762 76038
0 1389 5 9 1 76064
0 1390 7 9 2 65925 67428
0 1391 5 3 1 76075
0 1392 7 1 2 59247 76076
0 1393 5 1 1 1392
0 1394 7 1 2 76026 1393
0 1395 5 1 1 1394
0 1396 7 1 2 76066 1395
0 1397 5 1 1 1396
0 1398 7 8 2 62444 70301
0 1399 5 6 1 76087
0 1400 7 2 2 71677 76095
0 1401 5 1 1 76101
0 1402 7 1 2 71907 76102
0 1403 5 1 1 1402
0 1404 7 6 2 60988 62445
0 1405 5 5 1 76103
0 1406 7 1 2 76084 76109
0 1407 5 8 1 1406
0 1408 7 1 2 59744 76114
0 1409 5 1 1 1408
0 1410 7 1 2 64842 71861
0 1411 5 1 1 1410
0 1412 7 1 2 1409 1411
0 1413 7 1 2 1403 1412
0 1414 7 1 2 1397 1413
0 1415 7 1 2 1385 1414
0 1416 5 1 1 1415
0 1417 7 1 2 66104 1416
0 1418 5 1 1 1417
0 1419 7 8 2 61173 62446
0 1420 5 3 1 76122
0 1421 7 1 2 72993 75987
0 1422 5 2 1 1421
0 1423 7 1 2 76130 76133
0 1424 5 1 1 1423
0 1425 7 1 2 65926 1424
0 1426 5 1 1 1425
0 1427 7 2 2 66105 71908
0 1428 5 16 1 76135
0 1429 7 3 2 70720 76137
0 1430 5 1 1 76153
0 1431 7 1 2 1426 1430
0 1432 5 1 1 1431
0 1433 7 1 2 64611 1432
0 1434 5 1 1 1433
0 1435 7 38 2 61984 62447
0 1436 5 23 1 76156
0 1437 7 4 2 65763 76157
0 1438 5 4 1 76217
0 1439 7 2 2 72665 76221
0 1440 5 2 1 76225
0 1441 7 1 2 61174 76226
0 1442 5 1 1 1441
0 1443 7 6 2 62182 72577
0 1444 5 2 1 76229
0 1445 7 1 2 76230 76138
0 1446 7 1 2 1442 1445
0 1447 5 1 1 1446
0 1448 7 1 2 60201 1447
0 1449 7 1 2 1434 1448
0 1450 7 1 2 1418 1449
0 1451 7 1 2 1371 1450
0 1452 5 1 1 1451
0 1453 7 1 2 1335 1452
0 1454 5 1 1 1453
0 1455 7 6 2 64387 69627
0 1456 5 62 1 76237
0 1457 7 2 2 69168 74086
0 1458 5 3 1 76305
0 1459 7 1 2 66106 76307
0 1460 5 3 1 1459
0 1461 7 1 2 60038 76310
0 1462 5 1 1 1461
0 1463 7 8 2 60837 71344
0 1464 5 10 1 76313
0 1465 7 1 2 75703 76314
0 1466 5 1 1 1465
0 1467 7 1 2 1462 1466
0 1468 5 1 1 1467
0 1469 7 1 2 71159 1468
0 1470 5 1 1 1469
0 1471 7 22 2 60838 66979
0 1472 5 23 1 76331
0 1473 7 2 2 76332 73656
0 1474 7 1 2 76376 72895
0 1475 5 1 1 1474
0 1476 7 1 2 1470 1475
0 1477 5 1 1 1476
0 1478 7 1 2 65058 1477
0 1479 5 1 1 1478
0 1480 7 2 2 71410 72939
0 1481 7 9 2 66107 66980
0 1482 5 1 1 76380
0 1483 7 1 2 76381 74391
0 1484 7 1 2 76378 1483
0 1485 5 1 1 1484
0 1486 7 1 2 1479 1485
0 1487 5 1 1 1486
0 1488 7 1 2 76243 1487
0 1489 5 1 1 1488
0 1490 7 1 2 72666 72810
0 1491 5 2 1 1490
0 1492 7 1 2 72811 72896
0 1493 5 1 1 1492
0 1494 7 2 2 73394 73727
0 1495 5 2 1 76391
0 1496 7 1 2 62448 76392
0 1497 5 1 1 1496
0 1498 7 1 2 1493 1497
0 1499 5 2 1 1498
0 1500 7 1 2 71678 76395
0 1501 5 1 1 1500
0 1502 7 1 2 76389 1501
0 1503 5 1 1 1502
0 1504 7 1 2 69876 1503
0 1505 5 1 1 1504
0 1506 7 1 2 72046 74246
0 1507 7 1 2 70909 1506
0 1508 5 1 1 1507
0 1509 7 1 2 1505 1508
0 1510 5 1 1 1509
0 1511 7 1 2 70506 1510
0 1512 5 1 1 1511
0 1513 7 2 2 65764 73027
0 1514 5 21 1 76397
0 1515 7 12 2 59248 59423
0 1516 5 5 1 76420
0 1517 7 18 2 60760 76421
0 1518 5 3 1 76437
0 1519 7 1 2 76438 76396
0 1520 5 1 1 1519
0 1521 7 1 2 76390 1520
0 1522 5 1 1 1521
0 1523 7 1 2 76399 1522
0 1524 5 1 1 1523
0 1525 7 1 2 62800 1524
0 1526 7 1 2 1512 1525
0 1527 7 1 2 1489 1526
0 1528 7 1 2 1454 1527
0 1529 5 1 1 1528
0 1530 7 2 2 61985 71679
0 1531 5 2 1 76458
0 1532 7 1 2 72047 74313
0 1533 5 1 1 1532
0 1534 7 1 2 76460 1533
0 1535 5 1 1 1534
0 1536 7 1 2 59745 1535
0 1537 5 1 1 1536
0 1538 7 1 2 74571 74297
0 1539 5 1 1 1538
0 1540 7 1 2 1537 1539
0 1541 5 2 1 1540
0 1542 7 1 2 70111 76462
0 1543 5 1 1 1542
0 1544 7 1 2 70565 73028
0 1545 5 1 1 1544
0 1546 7 2 2 1543 1545
0 1547 5 1 1 76464
0 1548 7 1 2 74559 72461
0 1549 5 1 1 1548
0 1550 7 1 2 61986 1549
0 1551 5 1 1 1550
0 1552 7 2 2 64612 75034
0 1553 5 2 1 76466
0 1554 7 1 2 62183 76468
0 1555 5 1 1 1554
0 1556 7 1 2 1551 1555
0 1557 5 1 1 1556
0 1558 7 1 2 70112 1557
0 1559 5 2 1 1558
0 1560 7 1 2 70008 74208
0 1561 5 3 1 1560
0 1562 7 1 2 74298 76472
0 1563 5 2 1 1562
0 1564 7 6 2 60839 62184
0 1565 5 1 1 76477
0 1566 7 1 2 60039 76478
0 1567 5 2 1 1566
0 1568 7 21 2 59424 59746
0 1569 5 7 1 76485
0 1570 7 2 2 67186 76506
0 1571 5 3 1 76513
0 1572 7 1 2 61175 76514
0 1573 5 1 1 1572
0 1574 7 1 2 76483 1573
0 1575 5 1 1 1574
0 1576 7 1 2 66981 1575
0 1577 5 1 1 1576
0 1578 7 1 2 76475 1577
0 1579 7 1 2 76470 1578
0 1580 5 1 1 1579
0 1581 7 1 2 60989 1580
0 1582 5 1 1 1581
0 1583 7 1 2 76465 1582
0 1584 5 1 1 1583
0 1585 7 1 2 62449 1584
0 1586 5 1 1 1585
0 1587 7 2 2 72202 74775
0 1588 5 1 1 76518
0 1589 7 1 2 71475 71846
0 1590 5 1 1 1589
0 1591 7 1 2 1588 1590
0 1592 5 1 1 1591
0 1593 7 1 2 71345 1592
0 1594 5 1 1 1593
0 1595 7 4 2 67187 71284
0 1596 5 3 1 76520
0 1597 7 3 2 74539 76524
0 1598 5 2 1 76527
0 1599 7 1 2 74173 76002
0 1600 5 2 1 1599
0 1601 7 1 2 76530 76532
0 1602 5 1 1 1601
0 1603 7 2 2 62450 73029
0 1604 5 6 1 76534
0 1605 7 2 2 59425 76536
0 1606 5 1 1 76542
0 1607 7 1 2 60840 76543
0 1608 5 2 1 1607
0 1609 7 24 2 59747 66982
0 1610 5 6 1 76546
0 1611 7 6 2 67188 76547
0 1612 5 2 1 76576
0 1613 7 1 2 76582 71909
0 1614 5 1 1 1613
0 1615 7 1 2 60040 1614
0 1616 5 1 1 1615
0 1617 7 8 2 59249 67429
0 1618 5 1 1 76584
0 1619 7 4 2 69340 76585
0 1620 5 4 1 76592
0 1621 7 1 2 1616 76596
0 1622 7 1 2 76544 1621
0 1623 7 1 2 1602 1622
0 1624 5 1 1 1623
0 1625 7 1 2 72897 1624
0 1626 5 1 1 1625
0 1627 7 1 2 1594 1626
0 1628 5 1 1 1627
0 1629 7 1 2 66108 1628
0 1630 5 1 1 1629
0 1631 7 1 2 1586 1630
0 1632 5 1 1 1631
0 1633 7 1 2 65059 1632
0 1634 5 1 1 1633
0 1635 7 1 2 75781 75091
0 1636 5 2 1 1635
0 1637 7 1 2 69877 73599
0 1638 5 1 1 1637
0 1639 7 1 2 76600 1638
0 1640 5 1 1 1639
0 1641 7 1 2 72048 1640
0 1642 5 1 1 1641
0 1643 7 2 2 59748 75092
0 1644 5 2 1 76602
0 1645 7 1 2 69483 74476
0 1646 5 2 1 1645
0 1647 7 1 2 76604 76606
0 1648 5 1 1 1647
0 1649 7 1 2 67189 1648
0 1650 5 1 1 1649
0 1651 7 48 2 62185 62451
0 1652 5 24 1 76608
0 1653 7 4 2 71363 76656
0 1654 7 1 2 71680 74286
0 1655 7 1 2 76680 1654
0 1656 5 1 1 1655
0 1657 7 2 2 60041 65765
0 1658 5 1 1 76684
0 1659 7 1 2 1656 1658
0 1660 7 1 2 1650 1659
0 1661 7 1 2 1642 1660
0 1662 5 1 1 1661
0 1663 7 1 2 72812 1662
0 1664 5 1 1 1663
0 1665 7 2 2 60202 76609
0 1666 5 2 1 76686
0 1667 7 18 2 64613 65766
0 1668 5 2 1 76690
0 1669 7 2 2 69749 76691
0 1670 5 1 1 76710
0 1671 7 1 2 76687 76711
0 1672 5 1 1 1671
0 1673 7 1 2 72756 1672
0 1674 5 1 1 1673
0 1675 7 1 2 64388 1674
0 1676 5 1 1 1675
0 1677 7 9 2 64204 65767
0 1678 5 2 1 76712
0 1679 7 4 2 69360 76713
0 1680 5 7 1 76723
0 1681 7 2 2 70721 76724
0 1682 5 1 1 76734
0 1683 7 1 2 71515 1682
0 1684 5 1 1 1683
0 1685 7 19 2 65060 70722
0 1686 5 58 1 76736
0 1687 7 1 2 64614 76755
0 1688 7 1 2 1684 1687
0 1689 5 1 1 1688
0 1690 7 1 2 1676 1689
0 1691 7 1 2 1664 1690
0 1692 5 1 1 1691
0 1693 7 1 2 65927 1692
0 1694 5 1 1 1693
0 1695 7 19 2 65768 69750
0 1696 7 22 2 66109 61987
0 1697 5 3 1 76832
0 1698 7 4 2 64843 76833
0 1699 5 2 1 76857
0 1700 7 11 2 64389 62452
0 1701 5 6 1 76863
0 1702 7 8 2 62186 70723
0 1703 5 2 1 76880
0 1704 7 1 2 76864 76881
0 1705 5 2 1 1704
0 1706 7 1 2 76861 76890
0 1707 5 1 1 1706
0 1708 7 1 2 60203 1707
0 1709 5 1 1 1708
0 1710 7 2 2 60990 74477
0 1711 7 1 2 72813 76892
0 1712 5 1 1 1711
0 1713 7 1 2 1709 1712
0 1714 5 1 1 1713
0 1715 7 1 2 76813 1714
0 1716 5 1 1 1715
0 1717 7 1 2 67798 1716
0 1718 7 1 2 1694 1717
0 1719 7 1 2 1634 1718
0 1720 5 1 1 1719
0 1721 7 1 2 63263 1720
0 1722 7 1 2 1529 1721
0 1723 5 1 1 1722
0 1724 7 3 2 59250 69386
0 1725 5 7 1 76894
0 1726 7 9 2 70302 76897
0 1727 5 2 1 76904
0 1728 7 7 2 64390 76905
0 1729 5 15 1 76915
0 1730 7 2 2 76922 71346
0 1731 5 1 1 76937
0 1732 7 1 2 67190 74776
0 1733 5 1 1 1732
0 1734 7 1 2 64615 1733
0 1735 5 2 1 1734
0 1736 7 1 2 60991 76939
0 1737 5 1 1 1736
0 1738 7 1 2 1731 1737
0 1739 5 1 1 1738
0 1740 7 1 2 64844 1739
0 1741 5 1 1 1740
0 1742 7 5 2 62187 72049
0 1743 7 2 2 72828 76041
0 1744 5 1 1 76946
0 1745 7 1 2 76941 76947
0 1746 5 2 1 1745
0 1747 7 1 2 76895 73030
0 1748 7 1 2 74457 1747
0 1749 5 1 1 1748
0 1750 7 2 2 76948 1749
0 1751 5 1 1 76950
0 1752 7 1 2 62453 76951
0 1753 5 1 1 1752
0 1754 7 1 2 59749 73122
0 1755 5 11 1 1754
0 1756 7 2 2 72530 76952
0 1757 5 3 1 76963
0 1758 7 1 2 67430 76965
0 1759 5 1 1 1758
0 1760 7 1 2 60992 1759
0 1761 7 1 2 1753 1760
0 1762 5 1 1 1761
0 1763 7 5 2 60761 61988
0 1764 5 1 1 76968
0 1765 7 1 2 69085 76969
0 1766 5 1 1 1765
0 1767 7 3 2 66983 72050
0 1768 5 6 1 76973
0 1769 7 1 2 62188 76974
0 1770 5 1 1 1769
0 1771 7 1 2 1766 1770
0 1772 5 1 1 1771
0 1773 7 1 2 59251 1772
0 1774 5 1 1 1773
0 1775 7 1 2 76949 1774
0 1776 5 1 1 1775
0 1777 7 1 2 74144 1776
0 1778 5 1 1 1777
0 1779 7 5 2 64616 69225
0 1780 5 29 1 76982
0 1781 7 8 2 64845 67431
0 1782 5 4 1 77016
0 1783 7 18 2 59426 69484
0 1784 5 10 1 77028
0 1785 7 2 2 76158 77029
0 1786 5 1 1 77056
0 1787 7 1 2 77024 1786
0 1788 5 1 1 1787
0 1789 7 1 2 76987 1788
0 1790 5 1 1 1789
0 1791 7 1 2 1778 1790
0 1792 7 1 2 1762 1791
0 1793 7 1 2 1741 1792
0 1794 5 1 1 1793
0 1795 7 1 2 65061 1794
0 1796 5 1 1 1795
0 1797 7 24 2 64617 64846
0 1798 5 1 1 77058
0 1799 7 2 2 60204 77059
0 1800 7 2 2 67432 73123
0 1801 5 16 1 77084
0 1802 7 4 2 64205 77086
0 1803 5 1 1 77102
0 1804 7 2 2 65679 77103
0 1805 5 2 1 77106
0 1806 7 1 2 74515 77108
0 1807 5 1 1 1806
0 1808 7 1 2 77082 1807
0 1809 5 1 1 1808
0 1810 7 11 2 59750 67191
0 1811 5 6 1 77110
0 1812 7 2 2 62454 77111
0 1813 5 1 1 77127
0 1814 7 1 2 72051 72646
0 1815 7 2 2 76681 1814
0 1816 5 1 1 77129
0 1817 7 1 2 1813 1816
0 1818 5 1 1 1817
0 1819 7 1 2 71285 1818
0 1820 5 1 1 1819
0 1821 7 6 2 67433 69485
0 1822 5 1 1 77131
0 1823 7 1 2 76942 77132
0 1824 5 1 1 1823
0 1825 7 1 2 73547 74392
0 1826 5 2 1 1825
0 1827 7 1 2 71681 73600
0 1828 5 2 1 1827
0 1829 7 1 2 77137 77139
0 1830 7 1 2 1824 1829
0 1831 7 1 2 1820 1830
0 1832 5 1 1 1831
0 1833 7 1 2 65062 1832
0 1834 5 1 1 1833
0 1835 7 1 2 1809 1834
0 1836 5 1 1 1835
0 1837 7 1 2 65928 1836
0 1838 5 1 1 1837
0 1839 7 1 2 66110 1838
0 1840 7 1 2 1796 1839
0 1841 5 1 1 1840
0 1842 7 7 2 65063 65929
0 1843 5 1 1 77141
0 1844 7 3 2 64618 77142
0 1845 5 2 1 77148
0 1846 7 13 2 64847 71045
0 1847 5 8 1 77153
0 1848 7 3 2 60205 77166
0 1849 5 21 1 77174
0 1850 7 4 2 69050 73343
0 1851 5 3 1 77198
0 1852 7 1 2 77177 77199
0 1853 5 1 1 1852
0 1854 7 1 2 77151 1853
0 1855 5 1 1 1854
0 1856 7 1 2 69751 1855
0 1857 5 1 1 1856
0 1858 7 1 2 71623 71017
0 1859 5 1 1 1858
0 1860 7 1 2 1857 1859
0 1861 5 1 1 1860
0 1862 7 2 2 62455 1861
0 1863 5 1 1 77205
0 1864 7 4 2 69878 71682
0 1865 5 10 1 77207
0 1866 7 3 2 65064 77060
0 1867 5 1 1 77221
0 1868 7 1 2 77211 77222
0 1869 5 1 1 1868
0 1870 7 1 2 61176 1869
0 1871 7 1 2 1863 1870
0 1872 5 1 1 1871
0 1873 7 1 2 62801 1872
0 1874 7 1 2 1841 1873
0 1875 5 1 1 1874
0 1876 7 17 2 64391 65680
0 1877 5 5 1 77224
0 1878 7 6 2 64206 64619
0 1879 5 2 1 77246
0 1880 7 6 2 77225 77247
0 1881 5 4 1 77254
0 1882 7 2 2 62189 77260
0 1883 5 2 1 77264
0 1884 7 1 2 77265 73152
0 1885 5 1 1 1884
0 1886 7 2 2 74111 76194
0 1887 7 1 2 77268 77107
0 1888 5 1 1 1887
0 1889 7 2 2 67434 72774
0 1890 5 2 1 77270
0 1891 7 3 2 64392 77272
0 1892 5 2 1 77274
0 1893 7 1 2 76682 77275
0 1894 5 1 1 1893
0 1895 7 1 2 65769 74393
0 1896 5 3 1 1895
0 1897 7 1 2 73747 77279
0 1898 7 1 2 1894 1897
0 1899 7 1 2 1888 1898
0 1900 5 1 1 1899
0 1901 7 1 2 71046 1900
0 1902 5 1 1 1901
0 1903 7 1 2 1885 1902
0 1904 5 1 1 1903
0 1905 7 1 2 64848 1904
0 1906 5 1 1 1905
0 1907 7 1 2 60993 73124
0 1908 5 1 1 1907
0 1909 7 21 2 65930 62190
0 1910 5 9 1 77282
0 1911 7 1 2 77303 73153
0 1912 7 1 2 76692 1911
0 1913 7 1 2 1908 1912
0 1914 5 1 1 1913
0 1915 7 1 2 1906 1914
0 1916 5 1 1 1915
0 1917 7 1 2 67799 1916
0 1918 5 1 1 1917
0 1919 7 10 2 64620 62191
0 1920 5 7 1 77312
0 1921 7 4 2 64393 77313
0 1922 5 2 1 77329
0 1923 7 7 2 65770 61177
0 1924 7 2 2 77330 77335
0 1925 5 1 1 77342
0 1926 7 12 2 64849 62456
0 1927 5 4 1 77344
0 1928 7 1 2 77343 77345
0 1929 5 1 1 1928
0 1930 7 1 2 1918 1929
0 1931 5 1 1 1930
0 1932 7 1 2 65065 1931
0 1933 5 1 1 1932
0 1934 7 3 2 62192 72531
0 1935 5 2 1 77360
0 1936 7 15 2 61178 62802
0 1937 5 8 1 77365
0 1938 7 17 2 66111 67800
0 1939 5 1 1 77388
0 1940 7 1 2 77389 74478
0 1941 5 2 1 1940
0 1942 7 1 2 77380 77405
0 1943 5 2 1 1942
0 1944 7 1 2 77361 77407
0 1945 5 1 1 1944
0 1946 7 34 2 62457 67801
0 1947 5 6 1 77409
0 1948 7 2 2 77410 73768
0 1949 5 1 1 77449
0 1950 7 1 2 1945 1949
0 1951 5 1 1 1950
0 1952 7 1 2 65066 1951
0 1953 5 1 1 1952
0 1954 7 43 2 62458 62803
0 1955 5 17 1 77451
0 1956 7 8 2 62193 77452
0 1957 5 2 1 77511
0 1958 7 2 2 76834 77512
0 1959 7 2 2 60206 75915
0 1960 7 1 2 77521 77523
0 1961 5 1 1 1960
0 1962 7 1 2 1953 1961
0 1963 5 1 1 1962
0 1964 7 1 2 64394 1963
0 1965 5 1 1 1964
0 1966 7 6 2 65067 65681
0 1967 5 1 1 77525
0 1968 7 7 2 64207 77526
0 1969 5 1 1 77531
0 1970 7 1 2 76382 77411
0 1971 7 1 2 77532 1970
0 1972 5 1 1 1971
0 1973 7 1 2 1965 1972
0 1974 5 1 1 1973
0 1975 7 1 2 72681 1974
0 1976 5 1 1 1975
0 1977 7 1 2 1933 1976
0 1978 7 1 2 1875 1977
0 1979 5 1 1 1978
0 1980 7 1 2 68200 1979
0 1981 5 1 1 1980
0 1982 7 1 2 66360 1981
0 1983 7 1 2 1723 1982
0 1984 5 1 1 1983
0 1985 7 50 2 68581 63888
0 1986 7 23 2 66112 68201
0 1987 7 7 2 64850 77588
0 1988 5 1 1 77611
0 1989 7 2 2 71047 77612
0 1990 5 2 1 77618
0 1991 7 5 2 61179 76159
0 1992 5 1 1 77622
0 1993 7 1 2 63264 77623
0 1994 5 1 1 1993
0 1995 7 1 2 77620 1994
0 1996 5 1 1 1995
0 1997 7 1 2 65771 1996
0 1998 5 1 1 1997
0 1999 7 3 2 72485 76139
0 2000 7 1 2 63265 77627
0 2001 5 1 1 2000
0 2002 7 1 2 1998 2001
0 2003 5 1 1 2002
0 2004 7 1 2 73082 2003
0 2005 5 1 1 2004
0 2006 7 4 2 60762 72994
0 2007 5 4 1 77630
0 2008 7 1 2 62459 77634
0 2009 5 6 1 2008
0 2010 7 3 2 59252 77638
0 2011 5 2 1 77644
0 2012 7 1 2 65931 77645
0 2013 5 1 1 2012
0 2014 7 1 2 76027 2013
0 2015 5 1 1 2014
0 2016 7 1 2 72052 2015
0 2017 5 1 1 2016
0 2018 7 1 2 60763 70507
0 2019 5 1 1 2018
0 2020 7 2 2 73031 2019
0 2021 5 1 1 77649
0 2022 7 1 2 2021 74615
0 2023 5 1 1 2022
0 2024 7 1 2 72285 2023
0 2025 5 1 1 2024
0 2026 7 1 2 62460 2025
0 2027 5 1 1 2026
0 2028 7 1 2 69441 76036
0 2029 5 1 1 2028
0 2030 7 1 2 74560 70001
0 2031 5 1 1 2030
0 2032 7 1 2 76077 2031
0 2033 5 1 1 2032
0 2034 7 1 2 2029 2033
0 2035 7 1 2 2027 2034
0 2036 7 1 2 2017 2035
0 2037 5 1 1 2036
0 2038 7 1 2 66113 2037
0 2039 5 1 1 2038
0 2040 7 2 2 64621 74820
0 2041 5 1 1 77651
0 2042 7 1 2 76085 73172
0 2043 7 2 2 77652 2042
0 2044 5 1 1 77653
0 2045 7 6 2 59751 61180
0 2046 5 2 1 77655
0 2047 7 1 2 64851 77661
0 2048 7 1 2 76140 2047
0 2049 5 1 1 2048
0 2050 7 1 2 2044 2049
0 2051 7 1 2 2039 2050
0 2052 5 1 1 2051
0 2053 7 1 2 63266 2052
0 2054 5 1 1 2053
0 2055 7 1 2 2005 2054
0 2056 5 1 1 2055
0 2057 7 1 2 62804 2056
0 2058 5 1 1 2057
0 2059 7 6 2 61181 62194
0 2060 5 4 1 77663
0 2061 7 1 2 77664 76227
0 2062 5 2 1 2061
0 2063 7 3 2 71742 72486
0 2064 5 2 1 77675
0 2065 7 1 2 72995 77676
0 2066 5 1 1 2065
0 2067 7 2 2 62195 73728
0 2068 5 1 1 77680
0 2069 7 1 2 2066 2068
0 2070 5 1 1 2069
0 2071 7 1 2 67435 2070
0 2072 5 1 1 2071
0 2073 7 1 2 77673 2072
0 2074 5 1 1 2073
0 2075 7 1 2 62805 2074
0 2076 5 1 1 2075
0 2077 7 2 2 61182 71160
0 2078 5 11 1 77682
0 2079 7 14 2 65932 66114
0 2080 5 2 1 77695
0 2081 7 5 2 64622 77696
0 2082 5 4 1 77711
0 2083 7 1 2 60042 77716
0 2084 5 4 1 2083
0 2085 7 23 2 77684 77720
0 2086 5 5 1 77724
0 2087 7 3 2 61989 77725
0 2088 5 1 1 77752
0 2089 7 1 2 2088 74235
0 2090 5 1 1 2089
0 2091 7 1 2 65772 67802
0 2092 7 1 2 2090 2091
0 2093 5 1 1 2092
0 2094 7 1 2 2076 2093
0 2095 5 1 1 2094
0 2096 7 1 2 63267 2095
0 2097 5 1 1 2096
0 2098 7 49 2 62806 68202
0 2099 5 4 1 77755
0 2100 7 4 2 76835 70940
0 2101 5 2 1 77808
0 2102 7 1 2 61183 76222
0 2103 5 4 1 2102
0 2104 7 2 2 64852 77814
0 2105 5 1 1 77818
0 2106 7 1 2 77812 2105
0 2107 5 2 1 2106
0 2108 7 1 2 71048 77820
0 2109 5 1 1 2108
0 2110 7 1 2 64853 77809
0 2111 5 1 1 2110
0 2112 7 1 2 2109 2111
0 2113 5 1 1 2112
0 2114 7 1 2 73083 2113
0 2115 5 1 1 2114
0 2116 7 16 2 65933 77061
0 2117 5 5 1 77822
0 2118 7 4 2 77823 73154
0 2119 5 2 1 77843
0 2120 7 1 2 2115 77847
0 2121 5 1 1 2120
0 2122 7 1 2 77756 2121
0 2123 5 1 1 2122
0 2124 7 1 2 2097 2123
0 2125 5 1 1 2124
0 2126 7 1 2 69752 2125
0 2127 5 1 1 2126
0 2128 7 23 2 64854 65934
0 2129 5 2 1 77849
0 2130 7 3 2 64623 77850
0 2131 7 61 2 67803 63268
0 2132 5 11 1 77877
0 2133 7 2 2 66115 77878
0 2134 7 1 2 77874 77949
0 2135 5 2 1 2134
0 2136 7 1 2 2127 77951
0 2137 7 1 2 2058 2136
0 2138 5 1 1 2137
0 2139 7 1 2 65068 2138
0 2140 5 1 1 2139
0 2141 7 4 2 60207 72682
0 2142 7 1 2 77953 77810
0 2143 5 1 1 2142
0 2144 7 19 2 65069 66116
0 2145 5 6 1 77957
0 2146 7 1 2 71049 77976
0 2147 7 1 2 77819 2146
0 2148 5 1 1 2147
0 2149 7 1 2 2143 2148
0 2150 5 1 1 2149
0 2151 7 1 2 76231 2150
0 2152 5 1 1 2151
0 2153 7 13 2 64624 66117
0 2154 5 5 1 77982
0 2155 7 10 2 77983 77851
0 2156 5 4 1 78000
0 2157 7 5 2 60208 62461
0 2158 5 1 1 78014
0 2159 7 1 2 2158 76134
0 2160 5 1 1 2159
0 2161 7 1 2 78001 2160
0 2162 5 1 1 2161
0 2163 7 1 2 2152 2162
0 2164 5 1 1 2163
0 2165 7 1 2 62807 2164
0 2166 5 1 1 2165
0 2167 7 3 2 69753 73887
0 2168 5 3 1 78019
0 2169 7 11 2 66118 62196
0 2170 5 6 1 78025
0 2171 7 3 2 65935 78026
0 2172 5 2 1 78042
0 2173 7 1 2 67804 77346
0 2174 7 1 2 78043 2173
0 2175 7 1 2 78020 2174
0 2176 5 1 1 2175
0 2177 7 1 2 2166 2176
0 2178 5 1 1 2177
0 2179 7 1 2 63269 2178
0 2180 5 1 1 2179
0 2181 7 1 2 61395 2180
0 2182 7 1 2 2140 2181
0 2183 5 1 1 2182
0 2184 7 1 2 77538 2183
0 2185 7 1 2 1984 2184
0 2186 5 1 1 2185
0 2187 7 1 2 1289 2186
0 2188 5 1 1 2187
0 2189 7 1 2 66607 2188
0 2190 5 1 1 2189
0 2191 7 21 2 61623 63889
0 2192 7 5 2 64855 68582
0 2193 7 3 2 61990 76610
0 2194 5 5 1 78073
0 2195 7 1 2 71161 78076
0 2196 5 2 1 2195
0 2197 7 1 2 69754 78081
0 2198 5 1 1 2197
0 2199 7 2 2 73344 76611
0 2200 5 1 1 78083
0 2201 7 1 2 2198 2200
0 2202 5 1 1 2201
0 2203 7 1 2 65773 2202
0 2204 5 1 1 2203
0 2205 7 4 2 64625 77087
0 2206 5 2 1 78085
0 2207 7 1 2 65936 78086
0 2208 5 1 1 2207
0 2209 7 1 2 2204 2208
0 2210 5 1 1 2209
0 2211 7 1 2 62808 2210
0 2212 5 1 1 2211
0 2213 7 2 2 69051 73776
0 2214 5 3 1 78091
0 2215 7 1 2 77255 78092
0 2216 5 1 1 2215
0 2217 7 1 2 2212 2216
0 2218 5 1 1 2217
0 2219 7 1 2 78068 2218
0 2220 5 1 1 2219
0 2221 7 2 2 59253 74616
0 2222 5 3 1 78096
0 2223 7 2 2 60764 78097
0 2224 5 1 1 78101
0 2225 7 2 2 74762 2224
0 2226 5 1 1 78103
0 2227 7 1 2 72286 78104
0 2228 5 1 1 2227
0 2229 7 8 2 62197 72287
0 2230 5 5 1 78105
0 2231 7 24 2 66984 67805
0 2232 5 9 1 78118
0 2233 7 15 2 67436 63622
0 2234 5 2 1 78151
0 2235 7 1 2 78119 78152
0 2236 7 1 2 78113 2235
0 2237 7 1 2 2228 2236
0 2238 5 2 1 2237
0 2239 7 1 2 2220 78168
0 2240 5 1 1 2239
0 2241 7 1 2 66119 2240
0 2242 5 1 1 2241
0 2243 7 33 2 67437 62809
0 2244 5 4 1 78170
0 2245 7 5 2 67192 78171
0 2246 5 3 1 78207
0 2247 7 1 2 78208 74419
0 2248 5 1 1 2247
0 2249 7 6 2 59427 69459
0 2250 5 8 1 78215
0 2251 7 1 2 71286 78216
0 2252 5 1 1 2251
0 2253 7 2 2 74690 2252
0 2254 5 1 1 78229
0 2255 7 1 2 62462 73649
0 2256 5 1 1 2255
0 2257 7 1 2 76528 2256
0 2258 5 1 1 2257
0 2259 7 1 2 74112 2258
0 2260 5 1 1 2259
0 2261 7 1 2 2254 2260
0 2262 5 1 1 2261
0 2263 7 1 2 67806 2262
0 2264 5 1 1 2263
0 2265 7 1 2 2248 2264
0 2266 5 1 1 2265
0 2267 7 1 2 61184 2266
0 2268 5 1 1 2267
0 2269 7 1 2 77443 77381
0 2270 5 2 1 2269
0 2271 7 1 2 71683 78231
0 2272 5 1 1 2271
0 2273 7 3 2 67438 70113
0 2274 5 4 1 78233
0 2275 7 1 2 62810 78234
0 2276 5 1 1 2275
0 2277 7 1 2 2272 2276
0 2278 5 1 1 2277
0 2279 7 1 2 72996 2278
0 2280 5 1 1 2279
0 2281 7 28 2 67439 67807
0 2282 5 11 1 78240
0 2283 7 5 2 61991 78241
0 2284 7 1 2 71684 78279
0 2285 5 1 1 2284
0 2286 7 1 2 2280 2285
0 2287 5 1 1 2286
0 2288 7 1 2 69879 2287
0 2289 5 1 1 2288
0 2290 7 1 2 77366 73650
0 2291 5 1 1 2290
0 2292 7 10 2 60841 67808
0 2293 5 6 1 78284
0 2294 7 4 2 59428 78285
0 2295 5 1 1 78300
0 2296 7 1 2 74304 78301
0 2297 5 1 1 2296
0 2298 7 1 2 2291 2297
0 2299 5 1 1 2298
0 2300 7 1 2 67440 2299
0 2301 5 1 1 2300
0 2302 7 2 2 59254 69169
0 2303 5 2 1 78304
0 2304 7 4 2 73430 78305
0 2305 5 6 1 78308
0 2306 7 1 2 64856 78312
0 2307 5 5 1 2306
0 2308 7 1 2 78232 78318
0 2309 5 1 1 2308
0 2310 7 1 2 74385 76131
0 2311 5 1 1 2310
0 2312 7 1 2 67809 2311
0 2313 5 1 1 2312
0 2314 7 1 2 2309 2313
0 2315 7 1 2 2301 2314
0 2316 7 1 2 2289 2315
0 2317 5 1 1 2316
0 2318 7 1 2 71162 2317
0 2319 5 1 1 2318
0 2320 7 1 2 67193 74135
0 2321 5 2 1 2320
0 2322 7 1 2 76529 78323
0 2323 5 1 1 2322
0 2324 7 2 2 74113 2323
0 2325 5 1 1 78325
0 2326 7 5 2 60842 62463
0 2327 7 4 2 59429 78327
0 2328 5 2 1 78332
0 2329 7 1 2 67810 78336
0 2330 7 1 2 2325 2329
0 2331 5 1 1 2330
0 2332 7 4 2 70393 74434
0 2333 5 10 1 78338
0 2334 7 1 2 78342 72467
0 2335 5 1 1 2334
0 2336 7 1 2 61185 2335
0 2337 5 1 1 2336
0 2338 7 4 2 76333 73997
0 2339 5 7 1 78352
0 2340 7 1 2 74538 78353
0 2341 5 1 1 2340
0 2342 7 1 2 62811 2341
0 2343 7 1 2 2337 2342
0 2344 5 1 1 2343
0 2345 7 1 2 72898 2344
0 2346 7 1 2 2331 2345
0 2347 5 1 1 2346
0 2348 7 1 2 62198 78120
0 2349 5 1 1 2348
0 2350 7 1 2 77382 2349
0 2351 5 1 1 2350
0 2352 7 1 2 69486 2351
0 2353 5 1 1 2352
0 2354 7 22 2 67194 67811
0 2355 5 6 1 78363
0 2356 7 1 2 75719 78385
0 2357 5 4 1 2356
0 2358 7 1 2 69880 78142
0 2359 7 1 2 78391 2358
0 2360 5 1 1 2359
0 2361 7 8 2 67195 70114
0 2362 5 1 1 78395
0 2363 7 1 2 62812 78396
0 2364 5 1 1 2363
0 2365 7 1 2 2360 2364
0 2366 7 1 2 2353 2365
0 2367 5 1 1 2366
0 2368 7 1 2 72408 2367
0 2369 5 1 1 2368
0 2370 7 7 2 62199 70303
0 2371 5 7 1 78403
0 2372 7 3 2 76898 78404
0 2373 5 7 1 78417
0 2374 7 1 2 62464 78418
0 2375 5 1 1 2374
0 2376 7 2 2 67812 74114
0 2377 7 1 2 73501 78427
0 2378 7 1 2 2375 2377
0 2379 5 1 1 2378
0 2380 7 2 2 61186 72451
0 2381 5 1 1 78429
0 2382 7 1 2 62813 72899
0 2383 7 1 2 78430 2382
0 2384 5 1 1 2383
0 2385 7 1 2 2379 2384
0 2386 7 1 2 2369 2385
0 2387 5 1 1 2386
0 2388 7 1 2 72053 2387
0 2389 5 1 1 2388
0 2390 7 9 2 60994 62814
0 2391 7 5 2 59752 78431
0 2392 5 2 1 78440
0 2393 7 1 2 73756 78441
0 2394 5 1 1 2393
0 2395 7 1 2 2389 2394
0 2396 7 1 2 2347 2395
0 2397 7 1 2 2319 2396
0 2398 7 1 2 2268 2397
0 2399 5 1 1 2398
0 2400 7 1 2 63623 2399
0 2401 5 2 1 2400
0 2402 7 1 2 2242 78447
0 2403 5 1 1 2402
0 2404 7 1 2 65070 2403
0 2405 5 1 1 2404
0 2406 7 2 2 61187 76657
0 2407 5 2 1 78449
0 2408 7 1 2 64395 78451
0 2409 5 2 1 2408
0 2410 7 1 2 61188 77109
0 2411 5 1 1 2410
0 2412 7 1 2 65774 2411
0 2413 5 1 1 2412
0 2414 7 1 2 78453 2413
0 2415 5 1 1 2414
0 2416 7 1 2 73173 2415
0 2417 5 1 1 2416
0 2418 7 1 2 69755 74490
0 2419 5 1 1 2418
0 2420 7 2 2 71946 73032
0 2421 5 9 1 78455
0 2422 7 1 2 2419 78457
0 2423 5 2 1 2422
0 2424 7 3 2 65775 69628
0 2425 5 13 1 78468
0 2426 7 4 2 67196 78471
0 2427 5 3 1 78484
0 2428 7 2 2 71050 78488
0 2429 5 1 1 78491
0 2430 7 2 2 78466 78492
0 2431 5 1 1 78493
0 2432 7 1 2 62465 78494
0 2433 5 1 1 2432
0 2434 7 2 2 73764 2433
0 2435 7 1 2 66120 78495
0 2436 5 1 1 2435
0 2437 7 2 2 2417 2436
0 2438 5 1 1 78497
0 2439 7 1 2 62815 78498
0 2440 5 1 1 2439
0 2441 7 4 2 66121 72683
0 2442 5 2 1 78499
0 2443 7 11 2 65776 65937
0 2444 5 1 1 78505
0 2445 7 3 2 61992 78506
0 2446 5 1 1 78516
0 2447 7 1 2 78087 78517
0 2448 5 1 1 2447
0 2449 7 1 2 78503 2448
0 2450 5 1 1 2449
0 2451 7 1 2 69756 2450
0 2452 5 1 1 2451
0 2453 7 17 2 65938 61993
0 2454 5 1 1 78519
0 2455 7 3 2 64626 78520
0 2456 5 3 1 78536
0 2457 7 1 2 73174 78539
0 2458 5 1 1 2457
0 2459 7 1 2 64857 2458
0 2460 5 1 1 2459
0 2461 7 1 2 67813 2460
0 2462 7 1 2 2452 2461
0 2463 5 1 1 2462
0 2464 7 1 2 60209 2463
0 2465 7 1 2 2440 2464
0 2466 5 1 1 2465
0 2467 7 40 2 66122 62816
0 2468 5 23 1 78542
0 2469 7 2 2 60043 78543
0 2470 5 1 1 78605
0 2471 7 5 2 65777 72578
0 2472 5 4 1 78607
0 2473 7 12 2 65682 70441
0 2474 5 5 1 78616
0 2475 7 5 2 59753 78628
0 2476 5 4 1 78633
0 2477 7 2 2 60995 78634
0 2478 5 4 1 78642
0 2479 7 1 2 78612 78643
0 2480 5 2 1 2479
0 2481 7 1 2 62200 78648
0 2482 5 1 1 2481
0 2483 7 2 2 60996 73548
0 2484 5 22 1 78650
0 2485 7 2 2 71476 75774
0 2486 5 1 1 78674
0 2487 7 1 2 78652 2486
0 2488 5 1 1 2487
0 2489 7 1 2 62466 2488
0 2490 7 2 2 2482 2489
0 2491 5 1 1 78676
0 2492 7 1 2 78606 78677
0 2493 5 1 1 2492
0 2494 7 6 2 67814 71051
0 2495 7 4 2 64858 61189
0 2496 5 2 1 78684
0 2497 7 1 2 72532 78685
0 2498 7 1 2 78678 2497
0 2499 5 1 1 2498
0 2500 7 24 2 62201 62817
0 2501 5 4 1 78690
0 2502 7 2 2 66123 78691
0 2503 5 1 1 78718
0 2504 7 1 2 69881 78719
0 2505 7 1 2 73941 2504
0 2506 5 1 1 2505
0 2507 7 1 2 2499 2506
0 2508 5 1 1 2507
0 2509 7 1 2 66985 2508
0 2510 5 1 1 2509
0 2511 7 2 2 61994 78309
0 2512 5 2 1 78720
0 2513 7 2 2 59430 76479
0 2514 5 3 1 78724
0 2515 7 1 2 74825 75958
0 2516 5 1 1 2515
0 2517 7 1 2 78726 2516
0 2518 5 1 1 2517
0 2519 7 1 2 71163 2518
0 2520 5 1 1 2519
0 2521 7 1 2 78722 2520
0 2522 5 1 1 2521
0 2523 7 1 2 60044 2522
0 2524 5 1 1 2523
0 2525 7 2 2 74041 72203
0 2526 5 1 1 78729
0 2527 7 1 2 74826 78730
0 2528 5 1 1 2527
0 2529 7 1 2 2524 2528
0 2530 5 1 1 2529
0 2531 7 1 2 78544 2530
0 2532 5 1 1 2531
0 2533 7 1 2 2510 2532
0 2534 5 1 1 2533
0 2535 7 1 2 67441 2534
0 2536 5 1 1 2535
0 2537 7 1 2 2493 2536
0 2538 7 1 2 2466 2537
0 2539 5 1 1 2538
0 2540 7 1 2 63624 2539
0 2541 5 1 1 2540
0 2542 7 1 2 2405 2541
0 2543 5 1 1 2542
0 2544 7 1 2 63270 2543
0 2545 5 1 1 2544
0 2546 7 58 2 68203 63625
0 2547 5 4 1 78731
0 2548 7 15 2 60210 66124
0 2549 5 3 1 78793
0 2550 7 2 2 64859 78794
0 2551 5 2 1 78811
0 2552 7 2 2 72822 78813
0 2553 5 2 1 78815
0 2554 7 1 2 73141 78817
0 2555 5 1 1 2554
0 2556 7 1 2 60997 70554
0 2557 5 1 1 2556
0 2558 7 3 2 76814 78521
0 2559 5 1 1 78819
0 2560 7 1 2 73084 78820
0 2561 5 2 1 2560
0 2562 7 1 2 59754 78822
0 2563 5 1 1 2562
0 2564 7 1 2 2557 2563
0 2565 7 1 2 70434 2564
0 2566 5 2 1 2565
0 2567 7 1 2 77958 78824
0 2568 5 1 1 2567
0 2569 7 1 2 2555 2568
0 2570 5 1 1 2569
0 2571 7 1 2 62467 2570
0 2572 5 1 1 2571
0 2573 7 1 2 71364 78818
0 2574 5 1 1 2573
0 2575 7 1 2 78808 78688
0 2576 5 5 1 2575
0 2577 7 5 2 62202 78826
0 2578 5 1 1 78831
0 2579 7 1 2 72533 76865
0 2580 7 1 2 78832 2579
0 2581 5 1 1 2580
0 2582 7 1 2 2574 2581
0 2583 5 1 1 2582
0 2584 7 1 2 71052 2583
0 2585 5 1 1 2584
0 2586 7 5 2 64860 67197
0 2587 5 3 1 78836
0 2588 7 1 2 253 78837
0 2589 5 1 1 2588
0 2590 7 1 2 66125 72734
0 2591 5 1 1 2590
0 2592 7 1 2 2589 2591
0 2593 5 2 1 2592
0 2594 7 1 2 74247 78844
0 2595 5 1 1 2594
0 2596 7 1 2 2585 2595
0 2597 7 1 2 2572 2596
0 2598 5 1 1 2597
0 2599 7 1 2 62818 2598
0 2600 5 1 1 2599
0 2601 7 4 2 71527 71053
0 2602 5 2 1 78846
0 2603 7 4 2 66986 78172
0 2604 5 5 1 78852
0 2605 7 14 2 62203 67815
0 2606 7 3 2 64396 76160
0 2607 5 5 1 78875
0 2608 7 1 2 78861 78876
0 2609 5 1 1 2608
0 2610 7 1 2 78856 2609
0 2611 5 1 1 2610
0 2612 7 1 2 69757 2611
0 2613 5 1 1 2612
0 2614 7 7 2 67816 76612
0 2615 5 1 1 78883
0 2616 7 4 2 64397 72760
0 2617 5 5 1 78890
0 2618 7 1 2 78884 78891
0 2619 5 1 1 2618
0 2620 7 1 2 78212 2619
0 2621 5 1 1 2620
0 2622 7 1 2 71743 2621
0 2623 5 1 1 2622
0 2624 7 1 2 2613 2623
0 2625 5 2 1 2624
0 2626 7 1 2 78847 78899
0 2627 5 1 1 2626
0 2628 7 5 2 65071 67817
0 2629 5 9 1 78901
0 2630 7 3 2 70009 78902
0 2631 5 2 1 78915
0 2632 7 1 2 74809 78916
0 2633 5 1 1 2632
0 2634 7 1 2 2627 2633
0 2635 7 1 2 2600 2634
0 2636 5 1 1 2635
0 2637 7 1 2 78732 2636
0 2638 5 1 1 2637
0 2639 7 1 2 2545 2638
0 2640 5 1 1 2639
0 2641 7 1 2 66361 2640
0 2642 5 1 1 2641
0 2643 7 4 2 62468 72534
0 2644 5 2 1 78920
0 2645 7 1 2 67818 75408
0 2646 5 1 1 2645
0 2647 7 10 2 65939 62819
0 2648 5 6 1 78926
0 2649 7 4 2 64627 61396
0 2650 7 1 2 78927 78942
0 2651 5 2 1 2650
0 2652 7 1 2 2646 78946
0 2653 5 1 1 2652
0 2654 7 1 2 78921 2653
0 2655 5 1 1 2654
0 2656 7 1 2 66362 78679
0 2657 5 1 1 2656
0 2658 7 1 2 2655 2657
0 2659 5 1 1 2658
0 2660 7 1 2 62204 2659
0 2661 5 1 1 2660
0 2662 7 1 2 66363 78209
0 2663 5 1 1 2662
0 2664 7 1 2 2661 2663
0 2665 5 1 1 2664
0 2666 7 1 2 64398 2665
0 2667 5 1 1 2666
0 2668 7 6 2 65683 66364
0 2669 7 4 2 64208 78948
0 2670 5 1 1 78954
0 2671 7 17 2 61995 67819
0 2672 7 2 2 71054 78958
0 2673 5 1 1 78975
0 2674 7 1 2 78857 2673
0 2675 5 1 1 2674
0 2676 7 1 2 78955 2675
0 2677 5 1 1 2676
0 2678 7 1 2 2667 2677
0 2679 5 1 1 2678
0 2680 7 1 2 68204 2679
0 2681 5 1 1 2680
0 2682 7 2 2 61397 77879
0 2683 5 3 1 78977
0 2684 7 1 2 71055 74540
0 2685 5 1 1 2684
0 2686 7 3 2 61996 77088
0 2687 5 1 1 78982
0 2688 7 2 2 75896 78983
0 2689 5 1 1 78985
0 2690 7 1 2 64209 78986
0 2691 5 1 1 2690
0 2692 7 1 2 2685 2691
0 2693 5 1 1 2692
0 2694 7 1 2 78978 2693
0 2695 5 1 1 2694
0 2696 7 1 2 2681 2695
0 2697 5 1 1 2696
0 2698 7 1 2 63626 2697
0 2699 5 1 1 2698
0 2700 7 9 2 65940 66365
0 2701 7 1 2 72579 78987
0 2702 7 3 2 72761 77314
0 2703 7 27 2 62820 68583
0 2704 5 1 1 78999
0 2705 7 2 2 75674 79000
0 2706 7 1 2 78996 79026
0 2707 7 1 2 2701 2706
0 2708 5 1 1 2707
0 2709 7 1 2 2699 2708
0 2710 5 1 1 2709
0 2711 7 1 2 65072 2710
0 2712 5 1 1 2711
0 2713 7 21 2 63271 63627
0 2714 7 10 2 60211 67820
0 2715 5 1 1 79049
0 2716 7 1 2 66366 79050
0 2717 7 1 2 78984 2716
0 2718 5 1 1 2717
0 2719 7 11 2 62821 71056
0 2720 5 1 1 79059
0 2721 7 3 2 64399 61398
0 2722 7 1 2 73601 79070
0 2723 7 1 2 79060 2722
0 2724 5 1 1 2723
0 2725 7 1 2 2718 2724
0 2726 5 1 1 2725
0 2727 7 1 2 76815 2726
0 2728 5 1 1 2727
0 2729 7 5 2 64628 66367
0 2730 7 2 2 60212 79073
0 2731 7 1 2 67821 73777
0 2732 7 1 2 79078 2731
0 2733 5 1 1 2732
0 2734 7 1 2 2728 2733
0 2735 5 1 1 2734
0 2736 7 1 2 79028 2735
0 2737 5 1 1 2736
0 2738 7 1 2 2712 2737
0 2739 5 2 1 2738
0 2740 7 1 2 70724 79080
0 2741 5 1 1 2740
0 2742 7 6 2 70725 71057
0 2743 5 3 1 79082
0 2744 7 1 2 60213 79083
0 2745 5 1 1 2744
0 2746 7 1 2 78816 2745
0 2747 5 2 1 2746
0 2748 7 1 2 73085 79091
0 2749 5 1 1 2748
0 2750 7 1 2 77959 2431
0 2751 5 1 1 2750
0 2752 7 1 2 2749 2751
0 2753 5 1 1 2752
0 2754 7 1 2 62822 2753
0 2755 5 1 1 2754
0 2756 7 1 2 62823 79092
0 2757 5 1 1 2756
0 2758 7 1 2 71528 78976
0 2759 5 1 1 2758
0 2760 7 1 2 2757 2759
0 2761 5 2 1 2760
0 2762 7 1 2 76816 79093
0 2763 5 1 1 2762
0 2764 7 1 2 78918 2763
0 2765 7 1 2 2755 2764
0 2766 5 1 1 2765
0 2767 7 1 2 62469 2766
0 2768 5 1 1 2767
0 2769 7 11 2 65073 62824
0 2770 5 1 1 79095
0 2771 7 2 2 70010 79096
0 2772 7 1 2 67442 79106
0 2773 5 2 1 2772
0 2774 7 1 2 67822 78540
0 2775 5 3 1 2774
0 2776 7 2 2 71529 74505
0 2777 5 3 1 79113
0 2778 7 1 2 77494 79114
0 2779 7 1 2 79110 2778
0 2780 5 1 1 2779
0 2781 7 1 2 78919 2780
0 2782 5 1 1 2781
0 2783 7 1 2 69758 2782
0 2784 5 1 1 2783
0 2785 7 1 2 79108 2784
0 2786 7 1 2 2768 2785
0 2787 5 1 1 2786
0 2788 7 1 2 63272 2787
0 2789 5 1 1 2788
0 2790 7 8 2 66126 71018
0 2791 5 2 1 79118
0 2792 7 1 2 77757 79119
0 2793 7 1 2 481 2792
0 2794 5 1 1 2793
0 2795 7 1 2 2789 2794
0 2796 5 1 1 2795
0 2797 7 1 2 61399 2796
0 2798 5 1 1 2797
0 2799 7 1 2 77149 77613
0 2800 7 1 2 78900 2799
0 2801 5 1 1 2800
0 2802 7 1 2 2798 2801
0 2803 5 1 1 2802
0 2804 7 1 2 63628 2803
0 2805 5 1 1 2804
0 2806 7 1 2 2741 2805
0 2807 7 1 2 2642 2806
0 2808 5 1 1 2807
0 2809 7 1 2 78047 2808
0 2810 5 1 1 2809
0 2811 7 1 2 2190 2810
0 2812 5 1 1 2811
0 2813 7 1 2 65312 2812
0 2814 5 1 1 2813
0 2815 7 17 2 60432 63890
0 2816 7 5 2 61997 72580
0 2817 5 2 1 79145
0 2818 7 1 2 62825 79146
0 2819 5 1 1 2818
0 2820 7 1 2 72731 2819
0 2821 5 1 1 2820
0 2822 7 1 2 76613 2821
0 2823 5 1 1 2822
0 2824 7 2 2 62826 69759
0 2825 5 1 1 79152
0 2826 7 1 2 71058 79153
0 2827 5 1 1 2826
0 2828 7 1 2 2823 2827
0 2829 5 1 1 2828
0 2830 7 1 2 65778 78069
0 2831 7 1 2 2829 2830
0 2832 5 1 1 2831
0 2833 7 1 2 78169 2832
0 2834 5 1 1 2833
0 2835 7 1 2 66127 2834
0 2836 5 1 1 2835
0 2837 7 1 2 78448 2836
0 2838 5 1 1 2837
0 2839 7 1 2 65074 2838
0 2840 5 1 1 2839
0 2841 7 3 2 67443 69387
0 2842 5 3 1 79154
0 2843 7 1 2 73033 79155
0 2844 5 1 1 2843
0 2845 7 1 2 76110 2844
0 2846 5 1 1 2845
0 2847 7 1 2 72054 2846
0 2848 5 1 1 2847
0 2849 7 2 2 869 78337
0 2850 5 2 1 79160
0 2851 7 1 2 76111 79161
0 2852 5 1 1 2851
0 2853 7 1 2 70394 2852
0 2854 5 1 1 2853
0 2855 7 1 2 2848 2854
0 2856 5 1 1 2855
0 2857 7 1 2 59255 2856
0 2858 5 1 1 2857
0 2859 7 1 2 62470 74756
0 2860 7 1 2 78356 2859
0 2861 5 1 1 2860
0 2862 7 3 2 67444 76353
0 2863 5 1 1 79164
0 2864 7 1 2 60765 71365
0 2865 7 1 2 2863 2864
0 2866 7 1 2 2861 2865
0 2867 5 1 1 2866
0 2868 7 1 2 73589 73976
0 2869 5 1 1 2868
0 2870 7 1 2 59431 73602
0 2871 5 2 1 2870
0 2872 7 1 2 62471 71611
0 2873 5 1 1 2872
0 2874 7 1 2 79167 2873
0 2875 5 1 1 2874
0 2876 7 1 2 72829 2875
0 2877 5 1 1 2876
0 2878 7 1 2 2869 2877
0 2879 7 1 2 2867 2878
0 2880 7 1 2 2858 2879
0 2881 5 1 1 2880
0 2882 7 1 2 59755 2881
0 2883 5 1 1 2882
0 2884 7 1 2 67445 1751
0 2885 5 1 1 2884
0 2886 7 1 2 74426 2885
0 2887 5 1 1 2886
0 2888 7 1 2 60998 2887
0 2889 5 1 1 2888
0 2890 7 1 2 67446 78721
0 2891 5 1 1 2890
0 2892 7 1 2 2889 2891
0 2893 7 1 2 2883 2892
0 2894 5 1 1 2893
0 2895 7 1 2 60045 2894
0 2896 5 1 1 2895
0 2897 7 4 2 59756 71612
0 2898 5 2 1 79169
0 2899 7 1 2 61998 76586
0 2900 7 1 2 73068 2899
0 2901 7 1 2 79170 2900
0 2902 5 1 1 2901
0 2903 7 1 2 2896 2902
0 2904 5 1 1 2903
0 2905 7 1 2 66128 2904
0 2906 5 1 1 2905
0 2907 7 1 2 60214 2438
0 2908 5 1 1 2907
0 2909 7 1 2 62827 2908
0 2910 7 1 2 2906 2909
0 2911 5 1 1 2910
0 2912 7 1 2 66987 74238
0 2913 5 1 1 2912
0 2914 7 1 2 78809 2913
0 2915 5 1 1 2914
0 2916 7 1 2 69760 2915
0 2917 5 1 1 2916
0 2918 7 2 2 60215 73155
0 2919 5 1 1 79175
0 2920 7 1 2 60216 61999
0 2921 5 3 1 2920
0 2922 7 6 2 65779 66988
0 2923 5 1 1 79180
0 2924 7 1 2 79181 73903
0 2925 5 1 1 2924
0 2926 7 1 2 79177 2925
0 2927 5 1 1 2926
0 2928 7 1 2 71059 2927
0 2929 5 1 1 2928
0 2930 7 1 2 2919 2929
0 2931 7 1 2 2917 2930
0 2932 5 1 1 2931
0 2933 7 1 2 64861 2932
0 2934 5 1 1 2933
0 2935 7 7 2 65684 77248
0 2936 5 1 1 79186
0 2937 7 2 2 60217 77697
0 2938 5 1 1 79193
0 2939 7 1 2 79187 79194
0 2940 5 1 1 2939
0 2941 7 1 2 67823 2940
0 2942 7 1 2 2934 2941
0 2943 5 1 1 2942
0 2944 7 1 2 63629 2943
0 2945 7 1 2 2911 2944
0 2946 5 1 1 2945
0 2947 7 1 2 2840 2946
0 2948 5 1 1 2947
0 2949 7 1 2 66368 2948
0 2950 5 1 1 2949
0 2951 7 18 2 61400 63630
0 2952 5 3 1 79195
0 2953 7 1 2 74541 78917
0 2954 5 1 1 2953
0 2955 7 1 2 65075 78496
0 2956 5 1 1 2955
0 2957 7 2 2 75927 73125
0 2958 5 2 1 79216
0 2959 7 3 2 62472 77954
0 2960 7 1 2 79218 79220
0 2961 5 1 1 2960
0 2962 7 1 2 2956 2961
0 2963 5 1 1 2962
0 2964 7 1 2 66129 2963
0 2965 5 1 1 2964
0 2966 7 3 2 71947 71530
0 2967 5 2 1 79223
0 2968 7 1 2 69761 73603
0 2969 7 1 2 79224 2968
0 2970 5 1 1 2969
0 2971 7 1 2 77178 76123
0 2972 7 1 2 79219 2971
0 2973 5 1 1 2972
0 2974 7 1 2 2970 2973
0 2975 7 1 2 2965 2974
0 2976 5 1 1 2975
0 2977 7 1 2 62828 2976
0 2978 5 1 1 2977
0 2979 7 1 2 2954 2978
0 2980 5 1 1 2979
0 2981 7 1 2 79196 2980
0 2982 5 1 1 2981
0 2983 7 1 2 2950 2982
0 2984 5 1 1 2983
0 2985 7 1 2 66608 2984
0 2986 5 1 1 2985
0 2987 7 8 2 66369 79001
0 2988 7 2 2 71277 79228
0 2989 5 1 1 79236
0 2990 7 1 2 66609 79237
0 2991 5 2 1 2990
0 2992 7 5 2 62000 71060
0 2993 5 2 1 79240
0 2994 7 26 2 66370 61624
0 2995 5 3 1 79247
0 2996 7 1 2 65076 79248
0 2997 5 6 1 2996
0 2998 7 15 2 66610 67824
0 2999 5 2 1 79282
0 3000 7 3 2 61401 79283
0 3001 5 3 1 79299
0 3002 7 1 2 79276 79302
0 3003 5 1 1 3002
0 3004 7 1 2 70011 3003
0 3005 5 1 1 3004
0 3006 7 6 2 75146 75885
0 3007 5 25 1 79305
0 3008 7 2 2 79311 79284
0 3009 5 1 1 79336
0 3010 7 1 2 3005 3009
0 3011 5 1 1 3010
0 3012 7 1 2 79241 3011
0 3013 5 1 1 3012
0 3014 7 7 2 61625 75157
0 3015 7 6 2 62829 70012
0 3016 5 2 1 79345
0 3017 7 1 2 79338 79346
0 3018 5 1 1 3017
0 3019 7 1 2 3013 3018
0 3020 5 1 1 3019
0 3021 7 4 2 64210 63631
0 3022 7 1 2 75897 79353
0 3023 7 1 2 3020 3022
0 3024 5 1 1 3023
0 3025 7 1 2 79238 3024
0 3026 5 1 1 3025
0 3027 7 1 2 77089 3026
0 3028 5 1 1 3027
0 3029 7 9 2 61626 62205
0 3030 7 18 2 62830 63632
0 3031 7 5 2 62473 79366
0 3032 7 2 2 79357 79384
0 3033 5 1 1 79389
0 3034 7 5 2 64862 66371
0 3035 7 11 2 64400 65077
0 3036 5 1 1 79396
0 3037 7 3 2 66130 79397
0 3038 7 1 2 79391 79407
0 3039 7 1 2 79390 3038
0 3040 5 1 1 3039
0 3041 7 1 2 3028 3040
0 3042 7 1 2 2986 3041
0 3043 5 1 1 3042
0 3044 7 1 2 63273 3043
0 3045 5 1 1 3044
0 3046 7 1 2 66611 79081
0 3047 5 1 1 3046
0 3048 7 3 2 75898 77104
0 3049 5 1 1 79410
0 3050 7 3 2 64401 76614
0 3051 5 6 1 79413
0 3052 7 1 2 3049 79416
0 3053 5 1 1 3052
0 3054 7 2 2 79029 78988
0 3055 7 3 2 64629 61627
0 3056 7 1 2 79097 79424
0 3057 7 1 2 79422 3056
0 3058 7 1 2 3053 3057
0 3059 5 1 1 3058
0 3060 7 1 2 3047 3059
0 3061 5 1 1 3060
0 3062 7 1 2 70726 3061
0 3063 5 1 1 3062
0 3064 7 29 2 66612 68205
0 3065 5 4 1 79427
0 3066 7 3 2 63633 79428
0 3067 7 1 2 66372 79094
0 3068 5 1 1 3067
0 3069 7 9 2 65078 70013
0 3070 5 3 1 79463
0 3071 7 20 2 66373 62831
0 3072 5 4 1 79475
0 3073 7 1 2 79464 79495
0 3074 7 1 2 79111 3073
0 3075 5 1 1 3074
0 3076 7 1 2 3068 3075
0 3077 5 1 1 3076
0 3078 7 1 2 73142 3077
0 3079 5 1 1 3078
0 3080 7 1 2 75158 78825
0 3081 5 1 1 3080
0 3082 7 28 2 75539 75245
0 3083 5 1 1 79499
0 3084 7 1 2 79500 77824
0 3085 5 1 1 3084
0 3086 7 1 2 3081 3085
0 3087 5 1 1 3086
0 3088 7 1 2 66131 3087
0 3089 5 1 1 3088
0 3090 7 16 2 64630 65079
0 3091 5 1 1 79527
0 3092 7 5 2 66374 79528
0 3093 7 1 2 74699 79543
0 3094 5 1 1 3093
0 3095 7 1 2 3089 3094
0 3096 5 1 1 3095
0 3097 7 1 2 62832 3096
0 3098 5 1 1 3097
0 3099 7 1 2 3079 3098
0 3100 5 1 1 3099
0 3101 7 1 2 62474 3100
0 3102 5 1 1 3101
0 3103 7 17 2 66132 66375
0 3104 5 2 1 79548
0 3105 7 6 2 64863 67825
0 3106 5 1 1 79567
0 3107 7 1 2 79549 79568
0 3108 7 1 2 74810 3107
0 3109 5 1 1 3108
0 3110 7 1 2 79565 73075
0 3111 5 1 1 3110
0 3112 7 1 2 66376 78845
0 3113 5 1 1 3112
0 3114 7 1 2 72660 71061
0 3115 5 1 1 3114
0 3116 7 1 2 3113 3115
0 3117 5 1 1 3116
0 3118 7 1 2 67447 3117
0 3119 5 1 1 3118
0 3120 7 1 2 3111 3119
0 3121 5 1 1 3120
0 3122 7 1 2 62833 74655
0 3123 7 1 2 3121 3122
0 3124 5 1 1 3123
0 3125 7 1 2 3109 3124
0 3126 5 1 1 3125
0 3127 7 1 2 65080 3126
0 3128 5 1 1 3127
0 3129 7 3 2 60218 62206
0 3130 5 1 1 79573
0 3131 7 1 2 67448 72661
0 3132 5 1 1 3131
0 3133 7 1 2 3130 3132
0 3134 5 1 1 3133
0 3135 7 4 2 66133 79476
0 3136 5 1 1 79576
0 3137 7 1 2 77825 79577
0 3138 7 1 2 3134 3137
0 3139 5 1 1 3138
0 3140 7 1 2 3128 3139
0 3141 7 1 2 3102 3140
0 3142 5 1 1 3141
0 3143 7 1 2 79460 3142
0 3144 5 1 1 3143
0 3145 7 1 2 3063 3144
0 3146 7 1 2 3045 3145
0 3147 5 1 1 3146
0 3148 7 1 2 79128 3147
0 3149 5 1 1 3148
0 3150 7 2 2 2814 3149
0 3151 5 1 1 79580
0 3152 7 1 2 66789 3151
0 3153 5 1 1 3152
0 3154 7 1 2 67826 76854
0 3155 5 11 1 3154
0 3156 7 1 2 60046 78582
0 3157 5 3 1 3156
0 3158 7 3 2 79582 79593
0 3159 7 1 2 71062 79596
0 3160 5 1 1 3159
0 3161 7 1 2 79351 3160
0 3162 5 3 1 3161
0 3163 7 1 2 79411 79599
0 3164 5 1 1 3163
0 3165 7 2 2 77726 73086
0 3166 5 1 1 79602
0 3167 7 1 2 79603 77453
0 3168 5 1 1 3167
0 3169 7 1 2 3164 3168
0 3170 5 1 1 3169
0 3171 7 38 2 65313 66613
0 3172 5 54 1 79604
0 3173 7 8 2 75159 79605
0 3174 7 22 2 61836 63634
0 3175 5 1 1 79704
0 3176 7 7 2 63274 63891
0 3177 7 3 2 79705 79726
0 3178 7 1 2 79696 79733
0 3179 7 1 2 3170 3178
0 3180 5 1 1 3179
0 3181 7 1 2 3153 3180
0 3182 5 1 1 3181
0 3183 7 1 2 60646 3182
0 3184 5 1 1 3183
0 3185 7 1 2 61837 79581
0 3186 5 1 1 3185
0 3187 7 19 2 66614 68818
0 3188 5 1 1 79736
0 3189 7 3 2 60766 75105
0 3190 5 2 1 79755
0 3191 7 1 2 79074 79756
0 3192 5 1 1 3191
0 3193 7 39 2 61402 63275
0 3194 5 24 1 79760
0 3195 7 1 2 79761 69361
0 3196 5 1 1 3195
0 3197 7 1 2 3192 3196
0 3198 5 1 1 3197
0 3199 7 1 2 59256 3198
0 3200 5 1 1 3199
0 3201 7 6 2 60767 61403
0 3202 7 2 2 64211 71000
0 3203 7 1 2 79823 79829
0 3204 5 1 1 3203
0 3205 7 1 2 3200 3204
0 3206 5 1 1 3205
0 3207 7 1 2 72055 71744
0 3208 7 1 2 3206 3207
0 3209 5 1 1 3208
0 3210 7 5 2 64212 62001
0 3211 5 5 1 79831
0 3212 7 1 2 64631 72056
0 3213 7 1 2 79836 3212
0 3214 5 1 1 3213
0 3215 7 6 2 62002 71745
0 3216 5 6 1 79841
0 3217 7 1 2 60843 77226
0 3218 5 1 1 3217
0 3219 7 1 2 79847 3218
0 3220 5 1 1 3219
0 3221 7 1 2 64213 59757
0 3222 7 1 2 3220 3221
0 3223 5 1 1 3222
0 3224 7 1 2 3214 3223
0 3225 5 1 1 3224
0 3226 7 1 2 79762 3225
0 3227 5 1 1 3226
0 3228 7 1 2 75821 71301
0 3229 7 1 2 74790 3228
0 3230 5 1 1 3229
0 3231 7 1 2 79799 3230
0 3232 5 1 1 3231
0 3233 7 1 2 73555 74572
0 3234 7 1 2 3232 3233
0 3235 5 1 1 3234
0 3236 7 1 2 3227 3235
0 3237 7 1 2 3209 3236
0 3238 5 1 1 3237
0 3239 7 1 2 67198 3238
0 3240 5 1 1 3239
0 3241 7 10 2 59758 68206
0 3242 5 2 1 79853
0 3243 7 2 2 75409 79854
0 3244 5 1 1 79865
0 3245 7 4 2 61404 75430
0 3246 5 2 1 79867
0 3247 7 1 2 59432 79868
0 3248 5 1 1 3247
0 3249 7 1 2 3244 3248
0 3250 5 1 1 3249
0 3251 7 1 2 69487 3250
0 3252 5 1 1 3251
0 3253 7 25 2 61405 66989
0 3254 5 6 1 79873
0 3255 7 9 2 59759 63276
0 3256 7 1 2 79874 79904
0 3257 5 1 1 3256
0 3258 7 1 2 3252 3257
0 3259 5 1 1 3258
0 3260 7 1 2 65780 3259
0 3261 5 1 1 3260
0 3262 7 6 2 63277 72057
0 3263 7 8 2 61406 62003
0 3264 5 1 1 79919
0 3265 7 1 2 79913 79920
0 3266 5 1 1 3265
0 3267 7 1 2 68207 75425
0 3268 5 2 1 3267
0 3269 7 4 2 60844 68208
0 3270 5 2 1 79929
0 3271 7 1 2 79898 79933
0 3272 5 2 1 3271
0 3273 7 1 2 64402 79935
0 3274 7 1 2 79927 3273
0 3275 5 1 1 3274
0 3276 7 1 2 3266 3275
0 3277 5 1 1 3276
0 3278 7 1 2 59760 3277
0 3279 5 1 1 3278
0 3280 7 4 2 61407 71001
0 3281 5 4 1 79937
0 3282 7 3 2 66377 75106
0 3283 5 2 1 79945
0 3284 7 1 2 73556 79946
0 3285 5 1 1 3284
0 3286 7 1 2 79941 3285
0 3287 5 1 1 3286
0 3288 7 3 2 69882 74573
0 3289 5 3 1 79950
0 3290 7 1 2 3287 79951
0 3291 5 1 1 3290
0 3292 7 1 2 3279 3291
0 3293 7 1 2 3261 3292
0 3294 5 1 1 3293
0 3295 7 1 2 62207 3294
0 3296 5 1 1 3295
0 3297 7 3 2 59761 62004
0 3298 5 2 1 79956
0 3299 7 2 2 75822 76817
0 3300 5 1 1 79961
0 3301 7 1 2 79957 79962
0 3302 5 1 1 3301
0 3303 7 4 2 68209 69488
0 3304 5 1 1 79963
0 3305 7 1 2 66378 3304
0 3306 5 2 1 3305
0 3307 7 1 2 64632 60845
0 3308 7 1 2 1181 3307
0 3309 7 1 2 79967 3308
0 3310 5 1 1 3309
0 3311 7 1 2 3302 3310
0 3312 5 1 1 3311
0 3313 7 1 2 59433 3312
0 3314 5 1 1 3313
0 3315 7 1 2 3296 3314
0 3316 7 1 2 3240 3315
0 3317 5 1 1 3316
0 3318 7 1 2 3317 79465
0 3319 5 1 1 3318
0 3320 7 1 2 60846 76923
0 3321 5 1 1 3320
0 3322 7 1 2 74413 3321
0 3323 5 1 1 3322
0 3324 7 1 2 59762 3323
0 3325 5 1 1 3324
0 3326 7 2 2 72058 74791
0 3327 5 5 1 79969
0 3328 7 1 2 74561 79971
0 3329 5 1 1 3328
0 3330 7 1 2 67199 3329
0 3331 7 1 2 3325 3330
0 3332 5 1 1 3331
0 3333 7 6 2 59434 76334
0 3334 5 9 1 79976
0 3335 7 1 2 64633 79977
0 3336 5 1 1 3335
0 3337 7 1 2 73557 69762
0 3338 5 2 1 3337
0 3339 7 3 2 74574 79991
0 3340 5 5 1 79993
0 3341 7 1 2 62005 79994
0 3342 5 1 1 3341
0 3343 7 1 2 64634 76455
0 3344 5 8 1 3343
0 3345 7 3 2 64403 59763
0 3346 5 1 1 80009
0 3347 7 1 2 60847 3346
0 3348 5 1 1 3347
0 3349 7 1 2 66990 3348
0 3350 7 1 2 80001 3349
0 3351 5 1 1 3350
0 3352 7 1 2 3342 3351
0 3353 5 1 1 3352
0 3354 7 1 2 62208 3353
0 3355 5 1 1 3354
0 3356 7 1 2 3336 3355
0 3357 7 1 2 3332 3356
0 3358 5 1 1 3357
0 3359 7 35 2 66379 63278
0 3360 5 7 1 80012
0 3361 7 3 2 80013 76756
0 3362 5 2 1 80054
0 3363 7 1 2 71531 80055
0 3364 7 1 2 3358 3363
0 3365 5 1 1 3364
0 3366 7 1 2 3319 3365
0 3367 5 1 1 3366
0 3368 7 1 2 79737 3367
0 3369 5 1 1 3368
0 3370 7 3 2 59764 72852
0 3371 5 2 1 80059
0 3372 7 1 2 64404 80062
0 3373 5 2 1 3372
0 3374 7 1 2 59765 72789
0 3375 5 5 1 3374
0 3376 7 5 2 60848 70270
0 3377 5 6 1 80071
0 3378 7 2 2 64635 80076
0 3379 5 4 1 80082
0 3380 7 1 2 59257 80084
0 3381 5 2 1 3380
0 3382 7 3 2 80066 80088
0 3383 5 1 1 80090
0 3384 7 1 2 80063 80091
0 3385 5 1 1 3384
0 3386 7 4 2 80064 3385
0 3387 5 1 1 80093
0 3388 7 1 2 79312 73657
0 3389 7 1 2 80094 3388
0 3390 5 1 1 3389
0 3391 7 1 2 75463 70882
0 3392 7 1 2 72662 3391
0 3393 5 1 1 3392
0 3394 7 1 2 3390 3393
0 3395 5 1 1 3394
0 3396 7 1 2 68210 3395
0 3397 5 1 1 3396
0 3398 7 1 2 74562 74174
0 3399 5 2 1 3398
0 3400 7 4 2 60219 61190
0 3401 7 17 2 67200 63279
0 3402 7 2 2 79875 80103
0 3403 5 1 1 80120
0 3404 7 1 2 80099 80121
0 3405 7 1 2 80097 3404
0 3406 5 1 1 3405
0 3407 7 1 2 3397 3406
0 3408 5 1 1 3407
0 3409 7 1 2 78048 3408
0 3410 5 1 1 3409
0 3411 7 1 2 3369 3410
0 3412 5 1 1 3411
0 3413 7 1 2 65941 3412
0 3414 5 1 1 3413
0 3415 7 8 2 64405 67201
0 3416 5 2 1 80122
0 3417 7 2 2 72657 80130
0 3418 5 1 1 80132
0 3419 7 1 2 77266 80133
0 3420 5 2 1 3419
0 3421 7 3 2 78795 74854
0 3422 7 1 2 80134 80136
0 3423 5 2 1 3422
0 3424 7 1 2 62209 70222
0 3425 7 1 2 72885 3424
0 3426 5 1 1 3425
0 3427 7 2 2 72658 77267
0 3428 7 1 2 80141 76515
0 3429 5 1 1 3428
0 3430 7 1 2 70566 3429
0 3431 5 1 1 3430
0 3432 7 1 2 3426 3431
0 3433 5 1 1 3432
0 3434 7 1 2 79501 3433
0 3435 5 1 1 3434
0 3436 7 1 2 80139 3435
0 3437 5 1 1 3436
0 3438 7 1 2 68211 3437
0 3439 5 1 1 3438
0 3440 7 6 2 63280 75464
0 3441 5 1 1 80143
0 3442 7 1 2 1547 80144
0 3443 5 1 1 3442
0 3444 7 1 2 3439 3443
0 3445 5 1 1 3444
0 3446 7 1 2 78049 3445
0 3447 5 1 1 3446
0 3448 7 1 2 3414 3447
0 3449 5 1 1 3448
0 3450 7 1 2 65314 3449
0 3451 5 1 1 3450
0 3452 7 7 2 63281 79313
0 3453 5 1 1 80149
0 3454 7 3 2 64406 80150
0 3455 5 1 1 80156
0 3456 7 1 2 76818 79358
0 3457 7 1 2 80157 3456
0 3458 5 1 1 3457
0 3459 7 18 2 61408 66615
0 3460 5 1 1 80159
0 3461 7 5 2 60220 80160
0 3462 5 4 1 80177
0 3463 7 1 2 79277 80182
0 3464 5 9 1 3463
0 3465 7 5 2 65942 68212
0 3466 7 1 2 64636 80195
0 3467 7 1 2 72663 3466
0 3468 7 1 2 80186 3467
0 3469 5 1 1 3468
0 3470 7 1 2 3458 3469
0 3471 5 1 1 3470
0 3472 7 1 2 70727 3471
0 3473 5 1 1 3472
0 3474 7 1 2 65943 80095
0 3475 5 1 1 3474
0 3476 7 1 2 60047 76507
0 3477 5 1 1 3476
0 3478 7 1 2 67202 3477
0 3479 7 1 2 3475 3478
0 3480 5 1 1 3479
0 3481 7 1 2 64864 427
0 3482 5 1 1 3481
0 3483 7 1 2 59766 3482
0 3484 5 1 1 3483
0 3485 7 1 2 60048 70980
0 3486 5 2 1 3485
0 3487 7 1 2 62210 80200
0 3488 7 1 2 3484 3487
0 3489 5 1 1 3488
0 3490 7 1 2 3480 3489
0 3491 5 1 1 3490
0 3492 7 1 2 60049 72651
0 3493 5 1 1 3492
0 3494 7 1 2 3491 3493
0 3495 5 1 1 3494
0 3496 7 1 2 61191 3495
0 3497 5 1 1 3496
0 3498 7 4 2 60050 62211
0 3499 5 4 1 80202
0 3500 7 2 2 80060 72882
0 3501 5 2 1 80210
0 3502 7 1 2 80203 80211
0 3503 5 1 1 3502
0 3504 7 1 2 3497 3503
0 3505 5 1 1 3504
0 3506 7 1 2 79502 3505
0 3507 5 1 1 3506
0 3508 7 1 2 80140 3507
0 3509 5 1 1 3508
0 3510 7 1 2 66616 3509
0 3511 5 1 1 3510
0 3512 7 1 2 79466 79249
0 3513 7 1 2 80135 3512
0 3514 5 1 1 3513
0 3515 7 1 2 68213 3514
0 3516 7 1 2 3511 3515
0 3517 5 1 1 3516
0 3518 7 1 2 69489 74575
0 3519 5 3 1 3518
0 3520 7 4 2 73558 80214
0 3521 5 4 1 80217
0 3522 7 4 2 66991 70115
0 3523 7 1 2 80221 80225
0 3524 5 1 1 3523
0 3525 7 1 2 70728 3524
0 3526 5 1 1 3525
0 3527 7 1 2 62212 3526
0 3528 5 1 1 3527
0 3529 7 2 2 65944 67203
0 3530 5 2 1 80229
0 3531 7 2 2 80230 75704
0 3532 5 1 1 80233
0 3533 7 1 2 69490 80234
0 3534 5 2 1 3533
0 3535 7 2 2 59767 72452
0 3536 5 3 1 80237
0 3537 7 1 2 74380 80238
0 3538 5 1 1 3537
0 3539 7 1 2 80235 3538
0 3540 5 1 1 3539
0 3541 7 1 2 72059 3540
0 3542 5 1 1 3541
0 3543 7 6 2 59435 71411
0 3544 5 1 1 80242
0 3545 7 1 2 70116 80243
0 3546 5 1 1 3545
0 3547 7 2 2 70729 3546
0 3548 5 3 1 80248
0 3549 7 1 2 62006 80250
0 3550 5 2 1 3549
0 3551 7 9 2 67204 74576
0 3552 5 3 1 80255
0 3553 7 1 2 66992 74700
0 3554 5 1 1 3553
0 3555 7 1 2 69883 74381
0 3556 5 1 1 3555
0 3557 7 1 2 3554 3556
0 3558 5 1 1 3557
0 3559 7 1 2 80256 3558
0 3560 5 1 1 3559
0 3561 7 1 2 80253 3560
0 3562 7 1 2 3542 3561
0 3563 7 1 2 3528 3562
0 3564 5 1 1 3563
0 3565 7 1 2 75160 3564
0 3566 5 1 1 3565
0 3567 7 3 2 61409 71516
0 3568 5 22 1 80267
0 3569 7 2 2 62213 80270
0 3570 7 6 2 64637 65685
0 3571 7 6 2 64214 80294
0 3572 5 1 1 80300
0 3573 7 5 2 65945 71948
0 3574 5 1 1 80306
0 3575 7 6 2 80301 80307
0 3576 7 1 2 75246 80311
0 3577 7 1 2 80292 3576
0 3578 5 1 1 3577
0 3579 7 1 2 3566 3578
0 3580 5 1 1 3579
0 3581 7 1 2 61628 3580
0 3582 5 1 1 3581
0 3583 7 6 2 66617 75465
0 3584 5 2 1 80317
0 3585 7 2 2 70117 74299
0 3586 5 1 1 80325
0 3587 7 1 2 3586 3532
0 3588 5 1 1 3587
0 3589 7 1 2 74577 3588
0 3590 5 1 1 3589
0 3591 7 1 2 70223 74314
0 3592 5 1 1 3591
0 3593 7 1 2 80236 3592
0 3594 5 1 1 3593
0 3595 7 1 2 72060 3594
0 3596 5 1 1 3595
0 3597 7 2 2 61192 80204
0 3598 5 1 1 80327
0 3599 7 1 2 3598 80254
0 3600 7 1 2 3596 3599
0 3601 7 1 2 3590 3600
0 3602 5 1 1 3601
0 3603 7 1 2 80318 3602
0 3604 5 1 1 3603
0 3605 7 1 2 63282 3604
0 3606 7 1 2 3582 3605
0 3607 5 1 1 3606
0 3608 7 1 2 3517 3607
0 3609 5 1 1 3608
0 3610 7 1 2 3473 3609
0 3611 5 1 1 3610
0 3612 7 1 2 79129 3611
0 3613 5 1 1 3612
0 3614 7 1 2 3451 3613
0 3615 5 1 1 3614
0 3616 7 1 2 62475 3615
0 3617 5 1 1 3616
0 3618 7 14 2 65315 61629
0 3619 5 5 1 80329
0 3620 7 18 2 60433 66618
0 3621 5 7 1 80348
0 3622 7 6 2 80343 80366
0 3623 5 48 1 80373
0 3624 7 3 2 63892 80379
0 3625 7 3 2 62007 71949
0 3626 5 3 1 80430
0 3627 7 1 2 69763 79842
0 3628 5 2 1 3627
0 3629 7 1 2 80433 80436
0 3630 5 1 1 3629
0 3631 7 1 2 62214 3630
0 3632 5 1 1 3631
0 3633 7 2 2 62008 72535
0 3634 5 3 1 80438
0 3635 7 1 2 73534 80440
0 3636 5 1 1 3635
0 3637 7 1 2 65946 3636
0 3638 5 1 1 3637
0 3639 7 1 2 60999 70508
0 3640 5 4 1 3639
0 3641 7 1 2 64638 80443
0 3642 5 3 1 3641
0 3643 7 1 2 61193 80447
0 3644 7 1 2 3638 3643
0 3645 7 1 2 3632 3644
0 3646 5 1 1 3645
0 3647 7 2 2 66134 79996
0 3648 5 1 1 80450
0 3649 7 1 2 60051 3648
0 3650 7 1 2 3646 3649
0 3651 5 1 1 3650
0 3652 7 10 2 59768 60768
0 3653 5 2 1 80452
0 3654 7 7 2 66135 72997
0 3655 5 1 1 80464
0 3656 7 1 2 80453 80465
0 3657 5 1 1 3656
0 3658 7 2 2 77283 75735
0 3659 5 1 1 80471
0 3660 7 1 2 3657 3659
0 3661 5 1 1 3660
0 3662 7 1 2 59258 3661
0 3663 5 1 1 3662
0 3664 7 2 2 60769 70471
0 3665 5 1 1 80473
0 3666 7 1 2 74701 80474
0 3667 5 1 1 3666
0 3668 7 1 2 3663 3667
0 3669 5 1 1 3668
0 3670 7 1 2 71685 3669
0 3671 5 1 1 3670
0 3672 7 6 2 77227 76714
0 3673 5 5 1 80475
0 3674 7 1 2 59769 80472
0 3675 7 1 2 80481 3674
0 3676 5 1 1 3675
0 3677 7 1 2 3671 3676
0 3678 7 1 2 3651 3677
0 3679 5 1 1 3678
0 3680 7 1 2 68214 3679
0 3681 5 1 1 3680
0 3682 7 10 2 60849 76486
0 3683 5 3 1 80486
0 3684 7 1 2 80487 74908
0 3685 7 1 2 71340 3684
0 3686 5 1 1 3685
0 3687 7 1 2 3681 3686
0 3688 5 1 1 3687
0 3689 7 1 2 80427 3688
0 3690 5 1 1 3689
0 3691 7 2 2 64407 71449
0 3692 5 2 1 80499
0 3693 7 1 2 59770 80501
0 3694 5 1 1 3693
0 3695 7 4 2 69362 77249
0 3696 7 1 2 64408 80503
0 3697 5 1 1 3696
0 3698 7 1 2 62215 3697
0 3699 7 1 2 3694 3698
0 3700 5 1 1 3699
0 3701 7 1 2 64639 72652
0 3702 5 1 1 3701
0 3703 7 1 2 3700 3702
0 3704 5 1 1 3703
0 3705 7 13 2 65316 66136
0 3706 7 5 2 64865 80507
0 3707 7 21 2 63283 68819
0 3708 7 8 2 66619 80525
0 3709 7 1 2 80546 78507
0 3710 7 1 2 80520 3709
0 3711 7 1 2 3704 3710
0 3712 5 1 1 3711
0 3713 7 1 2 3690 3712
0 3714 5 1 1 3713
0 3715 7 1 2 79503 3714
0 3716 5 1 1 3715
0 3717 7 13 2 65081 60434
0 3718 7 4 2 79250 80554
0 3719 5 1 1 80567
0 3720 7 1 2 75466 80380
0 3721 5 3 1 3720
0 3722 7 1 2 3719 80571
0 3723 5 5 1 3722
0 3724 7 3 2 63893 80574
0 3725 7 7 2 64409 70730
0 3726 5 4 1 80582
0 3727 7 3 2 64640 80583
0 3728 5 1 1 80593
0 3729 7 1 2 75867 80594
0 3730 5 1 1 3729
0 3731 7 1 2 60850 70981
0 3732 5 4 1 3731
0 3733 7 11 2 72581 80596
0 3734 5 5 1 80600
0 3735 7 1 2 74982 80611
0 3736 5 1 1 3735
0 3737 7 1 2 3730 3736
0 3738 5 1 1 3737
0 3739 7 1 2 62216 3738
0 3740 5 1 1 3739
0 3741 7 12 2 68215 70014
0 3742 7 2 2 64641 80616
0 3743 5 1 1 80628
0 3744 7 3 2 62009 80104
0 3745 7 6 2 60770 61194
0 3746 7 5 2 59259 80633
0 3747 7 1 2 80630 80639
0 3748 5 1 1 3747
0 3749 7 1 2 3743 3748
0 3750 7 1 2 3740 3749
0 3751 5 1 1 3750
0 3752 7 1 2 80579 3751
0 3753 5 1 1 3752
0 3754 7 1 2 64215 80010
0 3755 7 1 2 74999 3754
0 3756 5 1 1 3755
0 3757 7 1 2 59436 80629
0 3758 5 1 1 3757
0 3759 7 3 2 64410 70567
0 3760 7 1 2 63284 80644
0 3761 5 1 1 3760
0 3762 7 1 2 3758 3761
0 3763 5 1 1 3762
0 3764 7 1 2 69629 69884
0 3765 7 1 2 3763 3764
0 3766 5 1 1 3765
0 3767 7 1 2 3756 3766
0 3768 5 1 1 3767
0 3769 7 1 2 62010 3768
0 3770 5 1 1 3769
0 3771 7 8 2 64216 64866
0 3772 5 2 1 80647
0 3773 7 6 2 65686 80648
0 3774 7 1 2 75155 80657
0 3775 5 1 1 3774
0 3776 7 1 2 75003 3775
0 3777 5 1 1 3776
0 3778 7 1 2 59437 3777
0 3779 5 1 1 3778
0 3780 7 7 2 63285 70568
0 3781 5 2 1 80663
0 3782 7 3 2 64411 70015
0 3783 5 1 1 80672
0 3784 7 1 2 79757 80673
0 3785 5 1 1 3784
0 3786 7 1 2 80670 3785
0 3787 5 1 1 3786
0 3788 7 1 2 59260 3787
0 3789 5 1 1 3788
0 3790 7 2 2 75705 73967
0 3791 5 1 1 80675
0 3792 7 1 2 3789 3791
0 3793 7 1 2 3779 3792
0 3794 5 1 1 3793
0 3795 7 1 2 64642 3794
0 3796 5 1 1 3795
0 3797 7 1 2 3770 3796
0 3798 5 1 1 3797
0 3799 7 1 2 62217 3798
0 3800 5 1 1 3799
0 3801 7 1 2 80676 79188
0 3802 5 1 1 3801
0 3803 7 1 2 3800 3802
0 3804 5 1 1 3803
0 3805 7 17 2 68820 79606
0 3806 7 3 2 75161 80677
0 3807 7 1 2 65781 80694
0 3808 7 1 2 3804 3807
0 3809 5 1 1 3808
0 3810 7 1 2 3753 3809
0 3811 5 1 1 3810
0 3812 7 1 2 65947 3811
0 3813 5 1 1 3812
0 3814 7 1 2 76548 74042
0 3815 5 4 1 3814
0 3816 7 1 2 73938 80697
0 3817 5 1 1 3816
0 3818 7 1 2 69885 3817
0 3819 5 1 1 3818
0 3820 7 5 2 60052 60851
0 3821 5 1 1 80701
0 3822 7 3 2 59438 80702
0 3823 5 1 1 80706
0 3824 7 1 2 64867 80496
0 3825 5 9 1 3824
0 3826 7 1 2 75782 80709
0 3827 5 1 1 3826
0 3828 7 1 2 3823 3827
0 3829 7 1 2 3819 3828
0 3830 5 1 1 3829
0 3831 7 1 2 63286 3830
0 3832 5 1 1 3831
0 3833 7 23 2 62218 68216
0 3834 7 5 2 62011 80718
0 3835 7 12 2 64412 64868
0 3836 7 1 2 72536 80746
0 3837 7 1 2 80741 3836
0 3838 5 1 1 3837
0 3839 7 1 2 3832 3838
0 3840 5 1 1 3839
0 3841 7 1 2 66137 80575
0 3842 7 1 2 3840 3841
0 3843 5 1 1 3842
0 3844 7 6 2 60852 61410
0 3845 5 2 1 80758
0 3846 7 2 2 74963 80759
0 3847 5 2 1 80766
0 3848 7 3 2 59771 80767
0 3849 5 1 1 80770
0 3850 7 7 2 66620 69491
0 3851 7 7 2 60053 68217
0 3852 7 4 2 65317 66993
0 3853 7 1 2 80780 80787
0 3854 7 1 2 71662 3853
0 3855 7 1 2 80773 3854
0 3856 7 1 2 80771 3855
0 3857 5 1 1 3856
0 3858 7 4 2 59772 65082
0 3859 5 1 1 80791
0 3860 7 4 2 60771 66380
0 3861 7 1 2 80792 80795
0 3862 7 1 2 71643 3861
0 3863 7 3 2 59261 72736
0 3864 7 20 2 67205 68218
0 3865 5 1 1 80802
0 3866 7 3 2 66994 80803
0 3867 7 1 2 80381 80822
0 3868 7 1 2 80799 3867
0 3869 7 1 2 3862 3868
0 3870 5 1 1 3869
0 3871 7 1 2 3857 3870
0 3872 7 1 2 3843 3871
0 3873 5 1 1 3872
0 3874 7 1 2 63894 3873
0 3875 5 1 1 3874
0 3876 7 1 2 3813 3875
0 3877 7 1 2 3716 3876
0 3878 5 1 1 3877
0 3879 7 1 2 67449 3878
0 3880 5 1 1 3879
0 3881 7 5 2 63895 79314
0 3882 7 66 2 60435 61630
0 3883 5 17 1 80830
0 3884 7 8 2 63287 80831
0 3885 5 1 1 80913
0 3886 7 2 2 69764 77753
0 3887 5 1 1 80921
0 3888 7 1 2 65782 80922
0 3889 5 1 1 3888
0 3890 7 1 2 78010 3889
0 3891 5 1 1 3890
0 3892 7 1 2 80914 3891
0 3893 5 1 1 3892
0 3894 7 10 2 60054 67206
0 3895 7 1 2 77589 80923
0 3896 7 1 2 80382 3895
0 3897 7 1 2 80096 3896
0 3898 5 1 1 3897
0 3899 7 1 2 3893 3898
0 3900 5 1 1 3899
0 3901 7 1 2 80825 3900
0 3902 5 1 1 3901
0 3903 7 3 2 67207 80098
0 3904 7 1 2 80933 76383
0 3905 5 1 1 3904
0 3906 7 1 2 74702 74209
0 3907 5 1 1 3906
0 3908 7 1 2 3905 3907
0 3909 5 1 1 3908
0 3910 7 1 2 80580 73968
0 3911 7 1 2 3909 3910
0 3912 5 1 1 3911
0 3913 7 1 2 3902 3912
0 3914 7 1 2 3880 3913
0 3915 7 1 2 3617 3914
0 3916 5 1 1 3915
0 3917 7 1 2 67827 3916
0 3918 5 1 1 3917
0 3919 7 3 2 59439 61411
0 3920 5 1 1 80936
0 3921 7 29 2 67450 68219
0 3922 5 3 1 80939
0 3923 7 2 2 70118 80428
0 3924 7 1 2 80940 80971
0 3925 5 1 1 3924
0 3926 7 1 2 62476 80547
0 3927 7 1 2 80521 3926
0 3928 5 1 1 3927
0 3929 7 1 2 3925 3928
0 3930 5 1 1 3929
0 3931 7 1 2 80937 3930
0 3932 5 1 1 3931
0 3933 7 4 2 65318 77698
0 3934 7 1 2 67451 80747
0 3935 7 10 2 68220 68821
0 3936 5 1 1 80977
0 3937 7 18 2 66381 66621
0 3938 5 1 1 80987
0 3939 7 1 2 80978 80988
0 3940 7 1 2 3934 3939
0 3941 7 1 2 80973 3940
0 3942 5 1 1 3941
0 3943 7 1 2 3932 3942
0 3944 5 1 1 3943
0 3945 7 1 2 67208 3944
0 3946 5 1 1 3945
0 3947 7 27 2 68221 63896
0 3948 7 3 2 60436 79550
0 3949 7 1 2 61631 76615
0 3950 7 1 2 81032 3949
0 3951 5 1 1 3950
0 3952 7 4 2 61412 70569
0 3953 5 1 1 81035
0 3954 7 1 2 80383 81036
0 3955 5 2 1 3954
0 3956 7 1 2 3951 81039
0 3957 5 1 1 3956
0 3958 7 1 2 81005 3957
0 3959 5 1 1 3958
0 3960 7 1 2 3946 3959
0 3961 5 1 1 3960
0 3962 7 1 2 60853 3961
0 3963 5 1 1 3962
0 3964 7 13 2 61413 62477
0 3965 5 6 1 81041
0 3966 7 4 2 66138 81042
0 3967 5 5 1 81060
0 3968 7 1 2 74352 81064
0 3969 5 1 1 3968
0 3970 7 1 2 80915 3969
0 3971 5 1 1 3970
0 3972 7 2 2 62478 71624
0 3973 5 2 1 81069
0 3974 7 11 2 60437 66139
0 3975 7 3 2 79251 81073
0 3976 7 1 2 81070 81084
0 3977 5 1 1 3976
0 3978 7 1 2 81040 3977
0 3979 5 1 1 3978
0 3980 7 1 2 68222 73126
0 3981 7 1 2 3979 3980
0 3982 5 1 1 3981
0 3983 7 1 2 3971 3982
0 3984 5 1 1 3983
0 3985 7 1 2 63897 3984
0 3986 5 1 1 3985
0 3987 7 1 2 3963 3986
0 3988 5 1 1 3987
0 3989 7 1 2 65083 3988
0 3990 5 1 1 3989
0 3991 7 9 2 60221 63898
0 3992 7 18 2 61632 63288
0 3993 5 2 1 81096
0 3994 7 6 2 66382 81097
0 3995 5 8 1 81116
0 3996 7 2 2 73156 81117
0 3997 5 1 1 81130
0 3998 7 1 2 60438 81131
0 3999 5 1 1 3998
0 4000 7 3 2 66383 70119
0 4001 5 1 1 81132
0 4002 7 1 2 70731 78221
0 4003 5 1 1 4002
0 4004 7 1 2 81133 4003
0 4005 5 1 1 4004
0 4006 7 3 2 62479 74356
0 4007 7 1 2 65948 81135
0 4008 5 1 1 4007
0 4009 7 1 2 4005 4008
0 4010 5 1 1 4009
0 4011 7 1 2 67209 4010
0 4012 5 1 1 4011
0 4013 7 3 2 76616 74357
0 4014 5 1 1 81138
0 4015 7 1 2 74353 4014
0 4016 5 1 1 4015
0 4017 7 1 2 72061 4016
0 4018 5 1 1 4017
0 4019 7 1 2 68223 4018
0 4020 7 1 2 4012 4019
0 4021 5 1 1 4020
0 4022 7 54 2 79642 80896
0 4023 5 3 1 81141
0 4024 7 1 2 63289 3953
0 4025 5 1 1 4024
0 4026 7 1 2 81142 4025
0 4027 7 1 2 4021 4026
0 4028 5 1 1 4027
0 4029 7 1 2 3999 4028
0 4030 5 1 1 4029
0 4031 7 1 2 81087 4030
0 4032 5 1 1 4031
0 4033 7 1 2 3990 4032
0 4034 5 1 1 4033
0 4035 7 1 2 59773 4034
0 4036 5 1 1 4035
0 4037 7 8 2 68224 74723
0 4038 5 3 1 81198
0 4039 7 2 2 77284 81199
0 4040 5 1 1 81209
0 4041 7 1 2 66384 80231
0 4042 5 1 1 4041
0 4043 7 2 2 75857 79800
0 4044 5 7 1 81211
0 4045 7 1 2 78328 81213
0 4046 7 1 2 4042 4045
0 4047 5 1 1 4046
0 4048 7 1 2 4040 4047
0 4049 5 1 1 4048
0 4050 7 1 2 66140 4049
0 4051 5 1 1 4050
0 4052 7 5 2 60055 71644
0 4053 5 2 1 81220
0 4054 7 1 2 80014 81221
0 4055 5 1 1 4054
0 4056 7 1 2 4051 4055
0 4057 5 1 1 4056
0 4058 7 1 2 65084 4057
0 4059 5 1 1 4058
0 4060 7 2 2 62480 75870
0 4061 5 1 1 81227
0 4062 7 4 2 60854 66141
0 4063 7 1 2 63290 81229
0 4064 7 1 2 81228 4063
0 4065 5 1 1 4064
0 4066 7 1 2 4059 4065
0 4067 5 1 1 4066
0 4068 7 1 2 80832 4067
0 4069 5 1 1 4068
0 4070 7 2 2 61195 69292
0 4071 5 1 1 81233
0 4072 7 2 2 60056 81234
0 4073 5 1 1 81235
0 4074 7 1 2 79315 81236
0 4075 5 1 1 4074
0 4076 7 1 2 60855 74394
0 4077 5 2 1 4076
0 4078 7 1 2 73620 81237
0 4079 5 5 1 4078
0 4080 7 1 2 75467 77699
0 4081 7 1 2 81239 4080
0 4082 5 1 1 4081
0 4083 7 1 2 4075 4082
0 4084 5 1 1 4083
0 4085 7 1 2 68225 4084
0 4086 5 1 1 4085
0 4087 7 3 2 60222 60856
0 4088 7 2 2 63291 81244
0 4089 5 1 1 81247
0 4090 7 1 2 81037 81248
0 4091 5 1 1 4090
0 4092 7 1 2 4086 4091
0 4093 5 1 1 4092
0 4094 7 1 2 81143 4093
0 4095 5 1 1 4094
0 4096 7 1 2 4069 4095
0 4097 5 1 1 4096
0 4098 7 1 2 59440 4097
0 4099 5 1 1 4098
0 4100 7 7 2 61414 62219
0 4101 7 2 2 65949 81249
0 4102 7 1 2 78796 81256
0 4103 5 1 1 4102
0 4104 7 1 2 70570 79504
0 4105 5 1 1 4104
0 4106 7 1 2 4103 4105
0 4107 5 1 1 4106
0 4108 7 1 2 60857 4107
0 4109 5 1 1 4108
0 4110 7 5 2 67210 70571
0 4111 7 1 2 75871 81258
0 4112 5 1 1 4111
0 4113 7 1 2 4109 4112
0 4114 5 1 1 4113
0 4115 7 1 2 80384 4114
0 4116 5 1 1 4115
0 4117 7 2 2 60858 77285
0 4118 5 1 1 81263
0 4119 7 1 2 78841 4118
0 4120 5 1 1 4119
0 4121 7 1 2 66142 80568
0 4122 7 1 2 4120 4121
0 4123 5 1 1 4122
0 4124 7 1 2 4116 4123
0 4125 5 1 1 4124
0 4126 7 1 2 80941 4125
0 4127 5 1 1 4126
0 4128 7 1 2 4099 4127
0 4129 5 1 1 4128
0 4130 7 1 2 63899 4129
0 4131 5 1 1 4130
0 4132 7 1 2 4036 4131
0 4133 5 1 1 4132
0 4134 7 1 2 66995 4133
0 4135 5 1 1 4134
0 4136 7 1 2 71663 80972
0 4137 5 1 1 4136
0 4138 7 10 2 64869 65319
0 4139 7 3 2 81265 77960
0 4140 7 11 2 66622 62012
0 4141 7 5 2 62220 68822
0 4142 7 1 2 81278 81289
0 4143 7 1 2 81275 4142
0 4144 5 1 1 4143
0 4145 7 1 2 4137 4144
0 4146 5 1 1 4145
0 4147 7 1 2 60859 4146
0 4148 5 1 1 4147
0 4149 7 8 2 65085 66623
0 4150 7 3 2 70016 81294
0 4151 7 7 2 67211 68823
0 4152 7 7 2 65320 65950
0 4153 7 1 2 81305 81312
0 4154 7 1 2 81302 4153
0 4155 5 1 1 4154
0 4156 7 1 2 4148 4155
0 4157 5 1 1 4156
0 4158 7 1 2 76487 4157
0 4159 5 1 1 4158
0 4160 7 11 2 65951 70017
0 4161 7 2 2 59774 81319
0 4162 7 4 2 66624 81306
0 4163 7 4 2 65321 60860
0 4164 7 2 2 65086 81336
0 4165 7 1 2 81332 81340
0 4166 7 2 2 81330 4165
0 4167 5 1 1 81342
0 4168 7 9 2 61196 71386
0 4169 5 1 1 81344
0 4170 7 2 2 80385 81345
0 4171 5 1 1 81353
0 4172 7 4 2 61633 77143
0 4173 7 1 2 81074 81355
0 4174 5 1 1 4173
0 4175 7 1 2 4171 4174
0 4176 5 1 1 4175
0 4177 7 1 2 63900 75959
0 4178 7 1 2 4176 4177
0 4179 5 1 1 4178
0 4180 7 1 2 4167 4179
0 4181 7 1 2 4159 4180
0 4182 5 1 1 4181
0 4183 7 1 2 61415 4182
0 4184 5 1 1 4183
0 4185 7 1 2 71412 78397
0 4186 5 1 1 4185
0 4187 7 2 2 70732 4186
0 4188 5 3 1 81359
0 4189 7 1 2 59441 81361
0 4190 5 1 1 4189
0 4191 7 2 2 70572 69086
0 4192 5 2 1 81364
0 4193 7 1 2 4190 81366
0 4194 5 3 1 4193
0 4195 7 1 2 65087 81368
0 4196 5 1 1 4195
0 4197 7 3 2 60223 75960
0 4198 7 1 2 77700 81371
0 4199 5 1 1 4198
0 4200 7 1 2 4196 4199
0 4201 5 1 1 4200
0 4202 7 1 2 79130 79252
0 4203 7 1 2 4201 4202
0 4204 5 1 1 4203
0 4205 7 1 2 4184 4204
0 4206 5 1 1 4205
0 4207 7 1 2 67452 4206
0 4208 5 1 1 4207
0 4209 7 1 2 70573 80187
0 4210 5 2 1 4209
0 4211 7 4 2 61634 79316
0 4212 5 3 1 81376
0 4213 7 1 2 73157 81377
0 4214 5 1 1 4213
0 4215 7 1 2 81374 4214
0 4216 5 1 1 4215
0 4217 7 1 2 60439 4216
0 4218 5 1 1 4217
0 4219 7 12 2 60224 65322
0 4220 7 4 2 60057 81383
0 4221 7 3 2 61635 74671
0 4222 7 1 2 81395 81399
0 4223 5 2 1 4222
0 4224 7 1 2 4218 81402
0 4225 5 1 1 4224
0 4226 7 1 2 63901 80257
0 4227 7 1 2 4225 4226
0 4228 5 1 1 4227
0 4229 7 1 2 4208 4228
0 4230 5 1 1 4229
0 4231 7 1 2 63292 4230
0 4232 5 1 1 4231
0 4233 7 1 2 4135 4232
0 4234 5 1 1 4233
0 4235 7 1 2 69886 4234
0 4236 5 1 1 4235
0 4237 7 5 2 63293 72537
0 4238 5 1 1 81404
0 4239 7 1 2 79921 81405
0 4240 5 1 1 4239
0 4241 7 1 2 3300 4240
0 4242 5 1 1 4241
0 4243 7 4 2 73087 74877
0 4244 5 2 1 81409
0 4245 7 1 2 4242 81410
0 4246 5 1 1 4245
0 4247 7 4 2 67212 73233
0 4248 5 6 1 81415
0 4249 7 5 2 69732 81419
0 4250 5 6 1 81425
0 4251 7 3 2 72062 81430
0 4252 5 1 1 81436
0 4253 7 2 2 4252 74636
0 4254 5 1 1 81439
0 4255 7 4 2 59442 70509
0 4256 5 2 1 81441
0 4257 7 2 2 60861 81442
0 4258 5 4 1 81447
0 4259 7 2 2 81440 81449
0 4260 5 1 1 81453
0 4261 7 1 2 59775 4260
0 4262 5 1 1 4261
0 4263 7 5 2 60862 72998
0 4264 5 3 1 81455
0 4265 7 1 2 77030 81456
0 4266 5 8 1 4265
0 4267 7 1 2 4262 81463
0 4268 5 1 1 4267
0 4269 7 1 2 63294 74724
0 4270 7 1 2 4268 4269
0 4271 5 1 1 4270
0 4272 7 1 2 4246 4271
0 4273 5 1 1 4272
0 4274 7 1 2 65952 4273
0 4275 5 1 1 4274
0 4276 7 6 2 67453 70510
0 4277 5 6 1 81471
0 4278 7 1 2 76531 81477
0 4279 5 1 1 4278
0 4280 7 2 2 69492 74395
0 4281 5 2 1 81483
0 4282 7 1 2 4279 81485
0 4283 5 1 1 4282
0 4284 7 1 2 80015 80488
0 4285 7 1 2 4283 4284
0 4286 5 1 1 4285
0 4287 7 1 2 4275 4286
0 4288 5 1 1 4287
0 4289 7 1 2 79738 4288
0 4290 5 1 1 4289
0 4291 7 14 2 61416 61636
0 4292 5 1 1 81487
0 4293 7 3 2 63902 80942
0 4294 7 2 2 71950 76906
0 4295 5 4 1 81504
0 4296 7 1 2 67213 81506
0 4297 5 1 1 4296
0 4298 7 3 2 64643 4297
0 4299 5 1 1 81510
0 4300 7 2 2 81501 4299
0 4301 7 1 2 81488 81513
0 4302 5 1 1 4301
0 4303 7 1 2 4290 4302
0 4304 5 1 1 4303
0 4305 7 1 2 65323 4304
0 4306 5 1 1 4305
0 4307 7 2 2 61417 80349
0 4308 7 1 2 81514 81515
0 4309 5 1 1 4308
0 4310 7 1 2 4306 4309
0 4311 5 1 1 4310
0 4312 7 1 2 71532 76757
0 4313 7 1 2 4311 4312
0 4314 5 1 1 4313
0 4315 7 1 2 64870 76988
0 4316 5 1 1 4315
0 4317 7 1 2 76439 77286
0 4318 5 1 1 4317
0 4319 7 1 2 4316 4318
0 4320 5 1 1 4319
0 4321 7 1 2 77590 4320
0 4322 5 1 1 4321
0 4323 7 2 2 80719 77701
0 4324 5 1 1 81517
0 4325 7 1 2 73969 76577
0 4326 5 1 1 4325
0 4327 7 1 2 4324 4326
0 4328 5 1 1 4327
0 4329 7 1 2 60863 4328
0 4330 5 1 1 4329
0 4331 7 1 2 67214 80617
0 4332 5 1 1 4331
0 4333 7 1 2 4330 4332
0 4334 5 1 1 4333
0 4335 7 1 2 76244 4334
0 4336 5 1 1 4335
0 4337 7 1 2 4322 4336
0 4338 5 1 1 4337
0 4339 7 1 2 67454 4338
0 4340 5 1 1 4339
0 4341 7 27 2 62481 68226
0 4342 7 12 2 66143 81519
0 4343 5 1 1 81546
0 4344 7 4 2 59776 69087
0 4345 5 15 1 81558
0 4346 7 1 2 71625 81559
0 4347 5 1 1 4346
0 4348 7 1 2 76989 74827
0 4349 5 1 1 4348
0 4350 7 1 2 4347 4349
0 4351 5 1 1 4350
0 4352 7 1 2 59443 4351
0 4353 5 1 1 4352
0 4354 7 4 2 60864 65953
0 4355 7 2 2 59777 81577
0 4356 7 1 2 67215 81581
0 4357 5 1 1 4356
0 4358 7 1 2 4353 4357
0 4359 5 1 1 4358
0 4360 7 1 2 81547 4359
0 4361 5 1 1 4360
0 4362 7 1 2 64644 69331
0 4363 5 1 1 4362
0 4364 7 1 2 76245 4363
0 4365 5 1 1 4364
0 4366 7 1 2 80002 76400
0 4367 5 2 1 4366
0 4368 7 1 2 67455 76990
0 4369 5 1 1 4368
0 4370 7 1 2 81583 4369
0 4371 7 1 2 4365 4370
0 4372 5 1 1 4371
0 4373 7 1 2 60058 4372
0 4374 5 1 1 4373
0 4375 7 4 2 60865 76246
0 4376 5 1 1 81585
0 4377 7 3 2 67456 77112
0 4378 5 1 1 81589
0 4379 7 1 2 66996 81590
0 4380 7 1 2 81586 4379
0 4381 5 1 1 4380
0 4382 7 1 2 63295 4381
0 4383 7 1 2 4374 4382
0 4384 5 1 1 4383
0 4385 7 1 2 68227 74840
0 4386 5 1 1 4385
0 4387 7 1 2 61197 4386
0 4388 7 1 2 4384 4387
0 4389 5 1 1 4388
0 4390 7 1 2 4361 4389
0 4391 7 1 2 4340 4390
0 4392 5 1 1 4391
0 4393 7 1 2 65088 4392
0 4394 5 1 1 4393
0 4395 7 6 2 61198 68228
0 4396 7 1 2 77206 81592
0 4397 5 1 1 4396
0 4398 7 1 2 4394 4397
0 4399 5 1 1 4398
0 4400 7 1 2 80833 4399
0 4401 5 1 1 4400
0 4402 7 7 2 67216 76335
0 4403 5 4 1 81598
0 4404 7 1 2 64645 81605
0 4405 5 1 1 4404
0 4406 7 1 2 76247 4405
0 4407 5 1 1 4406
0 4408 7 1 2 81584 4407
0 4409 5 1 1 4408
0 4410 7 1 2 62482 4409
0 4411 5 2 1 4410
0 4412 7 8 2 66997 76248
0 4413 5 3 1 81611
0 4414 7 5 2 60866 70511
0 4415 5 2 1 81622
0 4416 7 1 2 64646 81627
0 4417 7 1 2 81619 4416
0 4418 5 1 1 4417
0 4419 7 1 2 76078 4418
0 4420 5 1 1 4419
0 4421 7 1 2 81609 4420
0 4422 5 1 1 4421
0 4423 7 1 2 66144 4422
0 4424 5 1 1 4423
0 4425 7 8 2 65687 66145
0 4426 5 2 1 81629
0 4427 7 8 2 64217 81630
0 4428 5 4 1 81639
0 4429 7 4 2 66998 71347
0 4430 5 4 1 81651
0 4431 7 2 2 81640 81652
0 4432 5 1 1 81659
0 4433 7 3 2 65783 75736
0 4434 5 1 1 81661
0 4435 7 1 2 76617 81662
0 4436 5 1 1 4435
0 4437 7 1 2 4432 4436
0 4438 5 1 1 4437
0 4439 7 1 2 64413 4438
0 4440 5 1 1 4439
0 4441 7 1 2 77665 76161
0 4442 5 3 1 4441
0 4443 7 1 2 67457 80466
0 4444 5 1 1 4443
0 4445 7 1 2 81664 4444
0 4446 5 2 1 4445
0 4447 7 1 2 75916 81667
0 4448 5 1 1 4447
0 4449 7 2 2 4440 4448
0 4450 5 1 1 81669
0 4451 7 3 2 64647 61199
0 4452 7 1 2 73835 81671
0 4453 5 1 1 4452
0 4454 7 1 2 81670 4453
0 4455 7 1 2 4424 4454
0 4456 5 1 1 4455
0 4457 7 1 2 63296 4456
0 4458 5 1 1 4457
0 4459 7 5 2 67217 69765
0 4460 5 1 1 81674
0 4461 7 2 2 74087 81675
0 4462 5 1 1 81679
0 4463 7 1 2 77669 4462
0 4464 5 1 1 4463
0 4465 7 1 2 64414 4464
0 4466 5 1 1 4465
0 4467 7 2 2 65784 72999
0 4468 5 1 1 81681
0 4469 7 1 2 67458 81682
0 4470 5 1 1 4469
0 4471 7 1 2 77670 4470
0 4472 5 1 1 4471
0 4473 7 1 2 69766 4472
0 4474 5 1 1 4473
0 4475 7 1 2 4466 4474
0 4476 5 1 1 4475
0 4477 7 1 2 63297 4476
0 4478 5 1 1 4477
0 4479 7 2 2 70472 81548
0 4480 5 1 1 81683
0 4481 7 1 2 65785 70969
0 4482 7 1 2 81684 4481
0 4483 5 1 1 4482
0 4484 7 1 2 4478 4483
0 4485 5 1 1 4484
0 4486 7 1 2 72684 4485
0 4487 5 1 1 4486
0 4488 7 6 2 64648 73778
0 4489 5 16 1 81685
0 4490 7 1 2 69767 80618
0 4491 7 1 2 81686 4490
0 4492 5 1 1 4491
0 4493 7 1 2 4487 4492
0 4494 7 1 2 4458 4493
0 4495 5 1 1 4494
0 4496 7 1 2 60440 4495
0 4497 5 1 1 4496
0 4498 7 1 2 80374 4497
0 4499 5 1 1 4498
0 4500 7 1 2 59778 69293
0 4501 5 2 1 4500
0 4502 7 1 2 81707 76321
0 4503 5 3 1 4502
0 4504 7 2 2 61200 81709
0 4505 5 1 1 81712
0 4506 7 1 2 66146 76322
0 4507 5 1 1 4506
0 4508 7 1 2 59779 4507
0 4509 5 2 1 4508
0 4510 7 1 2 81714 4071
0 4511 5 2 1 4510
0 4512 7 1 2 76440 81716
0 4513 5 1 1 4512
0 4514 7 1 2 4505 4513
0 4515 5 1 1 4514
0 4516 7 1 2 60059 4515
0 4517 5 1 1 4516
0 4518 7 2 2 71645 81591
0 4519 5 1 1 81718
0 4520 7 1 2 76441 81719
0 4521 5 1 1 4520
0 4522 7 1 2 4517 4521
0 4523 5 1 1 4522
0 4524 7 1 2 68229 4523
0 4525 5 1 1 4524
0 4526 7 1 2 80897 4525
0 4527 5 1 1 4526
0 4528 7 1 2 60225 4527
0 4529 7 1 2 4499 4528
0 4530 5 1 1 4529
0 4531 7 1 2 4401 4530
0 4532 5 1 1 4531
0 4533 7 1 2 63903 4532
0 4534 5 1 1 4533
0 4535 7 3 2 63904 79855
0 4536 7 1 2 76249 81354
0 4537 5 1 1 4536
0 4538 7 7 2 66147 61637
0 4539 7 5 2 60441 81723
0 4540 7 9 2 65089 62483
0 4541 5 1 1 81735
0 4542 7 2 2 81730 81736
0 4543 7 1 2 74828 81744
0 4544 5 1 1 4543
0 4545 7 1 2 4537 4544
0 4546 5 1 1 4545
0 4547 7 1 2 81720 4546
0 4548 5 1 1 4547
0 4549 7 1 2 70224 69718
0 4550 5 1 1 4549
0 4551 7 1 2 70733 4550
0 4552 5 1 1 4551
0 4553 7 1 2 65090 4552
0 4554 5 1 1 4553
0 4555 7 1 2 2938 4554
0 4556 5 1 1 4555
0 4557 7 17 2 63905 80834
0 4558 5 1 1 81746
0 4559 7 1 2 4556 81747
0 4560 5 1 1 4559
0 4561 7 1 2 63298 4560
0 4562 5 1 1 4561
0 4563 7 18 2 65091 65324
0 4564 5 1 1 81763
0 4565 7 3 2 66625 81764
0 4566 7 4 2 62013 68824
0 4567 7 1 2 69493 81784
0 4568 7 1 2 81781 4567
0 4569 7 1 2 81331 4568
0 4570 5 1 1 4569
0 4571 7 10 2 60226 70574
0 4572 5 3 1 81788
0 4573 7 1 2 80429 81789
0 4574 5 1 1 4573
0 4575 7 1 2 68230 4574
0 4576 7 1 2 4570 4575
0 4577 5 1 1 4576
0 4578 7 1 2 59444 4577
0 4579 7 1 2 4562 4578
0 4580 5 1 1 4579
0 4581 7 3 2 61638 75431
0 4582 7 1 2 80555 81801
0 4583 5 1 1 4582
0 4584 7 1 2 60227 79964
0 4585 7 1 2 80386 4584
0 4586 5 1 1 4585
0 4587 7 1 2 4583 4586
0 4588 5 1 1 4587
0 4589 7 1 2 63906 70575
0 4590 7 1 2 4588 4589
0 4591 5 1 1 4590
0 4592 7 1 2 4580 4591
0 4593 5 1 1 4592
0 4594 7 1 2 67459 4593
0 4595 5 1 1 4594
0 4596 7 1 2 4548 4595
0 4597 5 1 1 4596
0 4598 7 1 2 69088 4597
0 4599 5 1 1 4598
0 4600 7 11 2 60772 67460
0 4601 5 2 1 81804
0 4602 7 5 2 59262 81805
0 4603 5 4 1 81817
0 4604 7 1 2 74214 81818
0 4605 7 1 2 81343 4604
0 4606 5 1 1 4605
0 4607 7 1 2 66385 4606
0 4608 7 1 2 4599 4607
0 4609 7 1 2 4534 4608
0 4610 5 1 1 4609
0 4611 7 1 2 60060 81717
0 4612 5 1 1 4611
0 4613 7 1 2 4519 4612
0 4614 5 1 1 4613
0 4615 7 1 2 59445 4614
0 4616 5 1 1 4615
0 4617 7 1 2 81562 69468
0 4618 5 1 1 4617
0 4619 7 1 2 70576 4618
0 4620 5 1 1 4619
0 4621 7 1 2 4616 4620
0 4622 5 1 1 4621
0 4623 7 1 2 69494 4622
0 4624 5 1 1 4623
0 4625 7 4 2 81560 74161
0 4626 5 9 1 81826
0 4627 7 1 2 78222 81830
0 4628 5 1 1 4627
0 4629 7 1 2 70577 4628
0 4630 5 1 1 4629
0 4631 7 1 2 4624 4630
0 4632 5 1 1 4631
0 4633 7 1 2 68231 4632
0 4634 5 1 1 4633
0 4635 7 1 2 80898 4634
0 4636 5 1 1 4635
0 4637 7 4 2 63907 79643
0 4638 7 5 2 81628 81445
0 4639 5 1 1 81843
0 4640 7 2 2 74563 73200
0 4641 5 1 1 81848
0 4642 7 1 2 81844 81849
0 4643 5 1 1 4642
0 4644 7 1 2 76079 4643
0 4645 5 1 1 4644
0 4646 7 1 2 81610 4645
0 4647 5 1 1 4646
0 4648 7 1 2 66148 4647
0 4649 5 1 1 4648
0 4650 7 4 2 67461 73000
0 4651 5 1 1 81850
0 4652 7 1 2 81851 77677
0 4653 5 1 1 4652
0 4654 7 1 2 77674 4653
0 4655 5 1 1 4654
0 4656 7 1 2 69768 4655
0 4657 5 1 1 4656
0 4658 7 2 2 60061 73127
0 4659 5 3 1 81854
0 4660 7 1 2 76953 81856
0 4661 7 1 2 76228 4660
0 4662 5 1 1 4661
0 4663 7 1 2 81691 4662
0 4664 5 1 1 4663
0 4665 7 1 2 61201 4664
0 4666 5 1 1 4665
0 4667 7 1 2 4657 4666
0 4668 7 1 2 4649 4667
0 4669 5 1 1 4668
0 4670 7 1 2 63299 4669
0 4671 5 1 1 4670
0 4672 7 1 2 77754 74449
0 4673 5 1 1 4672
0 4674 7 1 2 78011 4673
0 4675 5 3 1 4674
0 4676 7 9 2 68232 69769
0 4677 5 1 1 81862
0 4678 7 1 2 62484 81863
0 4679 7 1 2 81859 4678
0 4680 5 1 1 4679
0 4681 7 1 2 80835 4680
0 4682 7 1 2 4671 4681
0 4683 5 1 1 4682
0 4684 7 1 2 81839 4683
0 4685 7 1 2 4636 4684
0 4686 5 1 1 4685
0 4687 7 1 2 80312 80720
0 4688 5 1 1 4687
0 4689 7 2 2 63300 76488
0 4690 7 4 2 72861 69341
0 4691 5 2 1 81873
0 4692 7 1 2 81871 81874
0 4693 5 1 1 4692
0 4694 7 1 2 4688 4693
0 4695 5 1 1 4694
0 4696 7 1 2 62485 4695
0 4697 5 1 1 4696
0 4698 7 1 2 59780 74516
0 4699 5 3 1 4698
0 4700 7 4 2 74048 81879
0 4701 5 9 1 81882
0 4702 7 1 2 69495 81886
0 4703 5 1 1 4702
0 4704 7 1 2 81831 4703
0 4705 5 2 1 4704
0 4706 7 1 2 66999 81895
0 4707 5 1 1 4706
0 4708 7 4 2 71413 73998
0 4709 5 4 1 81897
0 4710 7 1 2 4707 81901
0 4711 5 1 1 4710
0 4712 7 1 2 63301 76080
0 4713 7 1 2 4711 4712
0 4714 5 1 1 4713
0 4715 7 1 2 4697 4714
0 4716 5 1 1 4715
0 4717 7 7 2 66149 66626
0 4718 5 1 1 81905
0 4719 7 1 2 68825 81906
0 4720 7 1 2 81266 4719
0 4721 7 1 2 4716 4720
0 4722 5 1 1 4721
0 4723 7 1 2 4686 4722
0 4724 5 1 1 4723
0 4725 7 1 2 65092 4724
0 4726 5 1 1 4725
0 4727 7 1 2 76250 81362
0 4728 5 1 1 4727
0 4729 7 6 2 69496 76489
0 4730 5 1 1 81912
0 4731 7 1 2 70734 4730
0 4732 5 1 1 4731
0 4733 7 1 2 70120 69089
0 4734 7 1 2 4732 4733
0 4735 5 1 1 4734
0 4736 7 1 2 4728 4735
0 4737 5 1 1 4736
0 4738 7 1 2 67462 4737
0 4739 5 1 1 4738
0 4740 7 1 2 70578 80934
0 4741 5 1 1 4740
0 4742 7 1 2 4739 4741
0 4743 5 1 1 4742
0 4744 7 1 2 67000 4743
0 4745 5 1 1 4744
0 4746 7 1 2 74578 74136
0 4747 5 1 1 4746
0 4748 7 1 2 72063 71348
0 4749 5 1 1 4748
0 4750 7 1 2 73559 4749
0 4751 7 1 2 4747 4750
0 4752 5 1 1 4751
0 4753 7 1 2 70579 4752
0 4754 5 1 1 4753
0 4755 7 1 2 63302 4754
0 4756 7 1 2 4745 4755
0 4757 5 1 1 4756
0 4758 7 4 2 64415 61202
0 4759 5 2 1 81918
0 4760 7 1 2 64649 81919
0 4761 5 1 1 4760
0 4762 7 1 2 81071 4761
0 4763 5 1 1 4762
0 4764 7 1 2 64871 4763
0 4765 5 1 1 4764
0 4766 7 1 2 71164 77202
0 4767 5 2 1 4766
0 4768 7 1 2 69770 81924
0 4769 5 3 1 4768
0 4770 7 1 2 61203 81926
0 4771 5 1 1 4770
0 4772 7 1 2 62486 4771
0 4773 5 1 1 4772
0 4774 7 1 2 4765 4773
0 4775 5 1 1 4774
0 4776 7 3 2 59263 76970
0 4777 5 5 1 81929
0 4778 7 1 2 80232 81932
0 4779 5 1 1 4778
0 4780 7 1 2 72064 4779
0 4781 5 1 1 4780
0 4782 7 2 2 69497 74271
0 4783 5 2 1 81937
0 4784 7 1 2 78727 81939
0 4785 7 1 2 4781 4784
0 4786 5 1 1 4785
0 4787 7 1 2 59781 4786
0 4788 5 1 1 4787
0 4789 7 1 2 66150 78723
0 4790 7 1 2 4788 4789
0 4791 5 1 1 4790
0 4792 7 1 2 4775 4791
0 4793 5 1 1 4792
0 4794 7 2 2 73604 74180
0 4795 5 1 1 81941
0 4796 7 1 2 77702 81942
0 4797 5 1 1 4796
0 4798 7 1 2 68233 4797
0 4799 7 1 2 4793 4798
0 4800 5 1 1 4799
0 4801 7 1 2 80387 4800
0 4802 7 1 2 4757 4801
0 4803 5 1 1 4802
0 4804 7 1 2 73779 77062
0 4805 5 3 1 4804
0 4806 7 1 2 77838 76223
0 4807 5 1 1 4806
0 4808 7 1 2 72685 76232
0 4809 7 1 2 4807 4808
0 4810 5 1 1 4809
0 4811 7 1 2 81943 4810
0 4812 5 1 1 4811
0 4813 7 7 2 66151 63303
0 4814 5 2 1 81946
0 4815 7 1 2 80836 81947
0 4816 7 1 2 4812 4815
0 4817 5 1 1 4816
0 4818 7 1 2 4803 4817
0 4819 5 1 1 4818
0 4820 7 1 2 60228 4819
0 4821 5 1 1 4820
0 4822 7 2 2 60442 65954
0 4823 7 2 2 77063 81955
0 4824 7 1 2 81098 81957
0 4825 7 1 2 4450 4824
0 4826 5 1 1 4825
0 4827 7 1 2 4821 4826
0 4828 5 1 1 4827
0 4829 7 1 2 63908 4828
0 4830 5 1 1 4829
0 4831 7 1 2 61418 4830
0 4832 7 1 2 4726 4831
0 4833 5 1 1 4832
0 4834 7 1 2 4610 4833
0 4835 5 1 1 4834
0 4836 7 5 2 81006 74672
0 4837 7 1 2 77955 81959
0 4838 5 1 1 4837
0 4839 7 8 2 64872 62014
0 4840 5 1 1 81964
0 4841 7 3 2 81737 81965
0 4842 7 8 2 66386 80526
0 4843 7 1 2 77712 81975
0 4844 7 1 2 81972 4843
0 4845 5 1 1 4844
0 4846 7 1 2 4838 4845
0 4847 5 1 1 4846
0 4848 7 1 2 73088 4847
0 4849 5 1 1 4848
0 4850 7 1 2 81960 77083
0 4851 5 1 1 4850
0 4852 7 1 2 4849 4851
0 4853 5 1 1 4852
0 4854 7 1 2 81144 4853
0 4855 5 1 1 4854
0 4856 7 24 2 61639 68234
0 4857 5 1 1 81983
0 4858 7 1 2 63909 74330
0 4859 7 1 2 81984 4858
0 4860 7 6 2 64873 80556
0 4861 7 1 2 76954 82007
0 4862 7 1 2 4859 4861
0 4863 5 1 1 4862
0 4864 7 3 2 70018 79317
0 4865 5 3 1 82013
0 4866 7 5 2 65093 74331
0 4867 5 2 1 82019
0 4868 7 1 2 82016 82024
0 4869 5 5 1 4868
0 4870 7 4 2 79131 81985
0 4871 5 1 1 82031
0 4872 7 1 2 82026 82032
0 4873 5 1 1 4872
0 4874 7 3 2 71387 74332
0 4875 5 1 1 82035
0 4876 7 4 2 68826 75675
0 4877 7 2 2 65325 81279
0 4878 7 1 2 82038 82042
0 4879 7 1 2 82036 4878
0 4880 5 1 1 4879
0 4881 7 1 2 4873 4880
0 4882 5 1 1 4881
0 4883 7 1 2 71063 73089
0 4884 7 1 2 4882 4883
0 4885 5 1 1 4884
0 4886 7 1 2 4863 4885
0 4887 7 1 2 4855 4886
0 4888 5 1 1 4887
0 4889 7 1 2 72538 4888
0 4890 5 1 1 4889
0 4891 7 1 2 4835 4890
0 4892 7 1 2 4314 4891
0 4893 7 1 2 4236 4892
0 4894 5 1 1 4893
0 4895 7 1 2 62834 4894
0 4896 5 1 1 4895
0 4897 7 4 2 80748 76693
0 4898 5 1 1 82044
0 4899 7 1 2 80721 76124
0 4900 7 1 2 82045 4899
0 4901 7 1 2 80581 4900
0 4902 5 1 1 4901
0 4903 7 1 2 4896 4902
0 4904 7 1 2 3918 4903
0 4905 5 1 1 4904
0 4906 7 1 2 68584 4905
0 4907 5 1 1 4906
0 4908 7 4 2 64650 68235
0 4909 7 2 2 78522 82048
0 4910 5 1 1 82052
0 4911 7 1 2 79412 82053
0 4912 5 1 1 4911
0 4913 7 1 2 64651 73646
0 4914 5 4 1 4913
0 4915 7 1 2 72065 82054
0 4916 5 1 1 4915
0 4917 7 1 2 76983 74491
0 4918 5 7 1 4917
0 4919 7 1 2 71287 82058
0 4920 5 1 1 4919
0 4921 7 1 2 80264 4920
0 4922 7 1 2 4916 4921
0 4923 5 1 1 4922
0 4924 7 1 2 73945 4923
0 4925 5 1 1 4924
0 4926 7 1 2 4912 4925
0 4927 5 1 1 4926
0 4928 7 1 2 64874 4927
0 4929 5 1 1 4928
0 4930 7 4 2 65688 71746
0 4931 5 2 1 82065
0 4932 7 1 2 72152 82069
0 4933 5 2 1 4932
0 4934 7 1 2 79982 82071
0 4935 5 1 1 4934
0 4936 7 1 2 74145 4935
0 4937 5 1 1 4936
0 4938 7 3 2 62487 76354
0 4939 5 5 1 82073
0 4940 7 2 2 59782 82076
0 4941 5 3 1 82081
0 4942 7 1 2 81478 82082
0 4943 5 1 1 4942
0 4944 7 3 2 60867 70473
0 4945 5 1 1 82086
0 4946 7 1 2 67463 82087
0 4947 5 1 1 4946
0 4948 7 1 2 76605 4947
0 4949 5 1 1 4948
0 4950 7 1 2 59446 4949
0 4951 5 1 1 4950
0 4952 7 1 2 4943 4951
0 4953 5 1 1 4952
0 4954 7 1 2 60773 4953
0 4955 5 1 1 4954
0 4956 7 1 2 4955 77138
0 4957 5 1 1 4956
0 4958 7 1 2 59264 4957
0 4959 5 1 1 4958
0 4960 7 1 2 4937 4959
0 4961 5 1 1 4960
0 4962 7 1 2 65955 4961
0 4963 5 1 1 4962
0 4964 7 3 2 69887 80244
0 4965 7 1 2 78074 82089
0 4966 5 1 1 4965
0 4967 7 1 2 4963 4966
0 4968 5 1 1 4967
0 4969 7 1 2 63304 4968
0 4970 5 1 1 4969
0 4971 7 1 2 4929 4970
0 4972 5 1 1 4971
0 4973 7 1 2 66152 4972
0 4974 5 1 1 4973
0 4975 7 2 2 67464 72582
0 4976 5 1 1 82092
0 4977 7 1 2 82093 78997
0 4978 5 1 1 4977
0 4979 7 2 2 59783 75928
0 4980 5 4 1 82094
0 4981 7 1 2 62221 82096
0 4982 5 1 1 4981
0 4983 7 1 2 76966 4982
0 4984 5 1 1 4983
0 4985 7 1 2 62015 4984
0 4986 5 1 1 4985
0 4987 7 1 2 73034 73860
0 4988 5 1 1 4987
0 4989 7 1 2 4986 4988
0 4990 5 1 1 4989
0 4991 7 1 2 60062 4990
0 4992 5 1 1 4991
0 4993 7 1 2 78842 76019
0 4994 7 1 2 4992 4993
0 4995 5 1 1 4994
0 4996 7 1 2 62488 4995
0 4997 5 1 1 4996
0 4998 7 1 2 4978 4997
0 4999 5 1 1 4998
0 5000 7 1 2 65956 4999
0 5001 5 1 1 5000
0 5002 7 1 2 67465 77064
0 5003 7 1 2 80601 5002
0 5004 5 1 1 5003
0 5005 7 1 2 5001 5004
0 5006 5 1 1 5005
0 5007 7 1 2 74983 5006
0 5008 5 1 1 5007
0 5009 7 1 2 4974 5008
0 5010 5 1 1 5009
0 5011 7 1 2 62835 5010
0 5012 5 1 1 5011
0 5013 7 2 2 67218 80602
0 5014 7 1 2 70883 82100
0 5015 5 1 1 5014
0 5016 7 1 2 64652 81505
0 5017 5 1 1 5016
0 5018 7 1 2 70019 5017
0 5019 5 1 1 5018
0 5020 7 1 2 5015 5019
0 5021 5 1 1 5020
0 5022 7 1 2 65957 5021
0 5023 5 1 1 5022
0 5024 7 1 2 73771 1925
0 5025 5 1 1 5024
0 5026 7 1 2 75979 5025
0 5027 5 1 1 5026
0 5028 7 12 2 65786 66153
0 5029 5 1 1 82102
0 5030 7 8 2 64416 82103
0 5031 5 2 1 82114
0 5032 7 1 2 67219 82115
0 5033 5 1 1 5032
0 5034 7 1 2 5027 5033
0 5035 5 1 1 5034
0 5036 7 1 2 64875 5035
0 5037 5 1 1 5036
0 5038 7 1 2 5023 5037
0 5039 5 1 1 5038
0 5040 7 1 2 62489 5039
0 5041 5 1 1 5040
0 5042 7 2 2 67466 77727
0 5043 5 1 1 82124
0 5044 7 1 2 74462 82125
0 5045 5 1 1 5044
0 5046 7 1 2 5041 5045
0 5047 5 1 1 5046
0 5048 7 1 2 77880 5047
0 5049 5 1 1 5048
0 5050 7 1 2 5012 5049
0 5051 5 1 1 5050
0 5052 7 1 2 80388 5051
0 5053 5 1 1 5052
0 5054 7 1 2 80497 78485
0 5055 5 1 1 5054
0 5056 7 1 2 59784 69226
0 5057 5 1 1 5056
0 5058 7 1 2 69888 76943
0 5059 5 1 1 5058
0 5060 7 2 2 5057 5059
0 5061 5 1 1 82126
0 5062 7 1 2 69968 79182
0 5063 5 1 1 5062
0 5064 7 1 2 82127 5063
0 5065 7 1 2 5055 5064
0 5066 5 1 1 5065
0 5067 7 1 2 62490 5066
0 5068 5 1 1 5067
0 5069 7 7 2 65689 62491
0 5070 5 1 1 82128
0 5071 7 6 2 64218 82129
0 5072 5 5 1 82135
0 5073 7 1 2 69170 82136
0 5074 5 1 1 5073
0 5075 7 7 2 64653 67467
0 5076 7 1 2 72539 82146
0 5077 5 1 1 5076
0 5078 7 1 2 5074 5077
0 5079 7 1 2 5068 5078
0 5080 5 1 1 5079
0 5081 7 2 2 67828 5080
0 5082 5 1 1 82153
0 5083 7 1 2 80935 78853
0 5084 5 1 1 5083
0 5085 7 1 2 5082 5084
0 5086 5 1 1 5085
0 5087 7 1 2 65958 5086
0 5088 5 1 1 5087
0 5089 7 1 2 67468 76463
0 5090 5 1 1 5089
0 5091 7 1 2 72862 77631
0 5092 5 3 1 5091
0 5093 7 1 2 59447 70388
0 5094 5 1 1 5093
0 5095 7 3 2 82155 5094
0 5096 5 3 1 82158
0 5097 7 1 2 74146 82161
0 5098 5 1 1 5097
0 5099 7 1 2 5090 5098
0 5100 5 1 1 5099
0 5101 7 1 2 62836 5100
0 5102 5 1 1 5101
0 5103 7 1 2 5088 5102
0 5104 5 1 1 5103
0 5105 7 25 2 65326 68236
0 5106 5 3 1 82164
0 5107 7 7 2 66627 70580
0 5108 7 1 2 82165 82192
0 5109 7 1 2 5104 5108
0 5110 5 1 1 5109
0 5111 7 1 2 5053 5110
0 5112 5 1 1 5111
0 5113 7 1 2 68827 5112
0 5114 5 1 1 5113
0 5115 7 1 2 59785 76067
0 5116 5 1 1 5115
0 5117 7 1 2 71686 70271
0 5118 5 3 1 5117
0 5119 7 2 2 5116 82199
0 5120 5 1 1 82202
0 5121 7 1 2 62492 82203
0 5122 5 1 1 5121
0 5123 7 3 2 70304 73861
0 5124 5 2 1 82204
0 5125 7 4 2 65787 67469
0 5126 7 1 2 82205 82209
0 5127 5 1 1 5126
0 5128 7 1 2 5122 5127
0 5129 5 1 1 5128
0 5130 7 1 2 64876 5129
0 5131 5 1 1 5130
0 5132 7 1 2 71910 5131
0 5133 5 1 1 5132
0 5134 7 1 2 59448 72830
0 5135 5 1 1 5134
0 5136 7 2 2 62493 5135
0 5137 7 1 2 80083 82213
0 5138 5 1 1 5137
0 5139 7 1 2 67470 80441
0 5140 5 3 1 5139
0 5141 7 1 2 67220 82215
0 5142 7 1 2 5138 5141
0 5143 5 1 1 5142
0 5144 7 1 2 5133 5143
0 5145 5 1 1 5144
0 5146 7 1 2 61204 5145
0 5147 5 1 1 5146
0 5148 7 1 2 62494 74564
0 5149 5 1 1 5148
0 5150 7 1 2 70121 81479
0 5151 7 1 2 5149 5150
0 5152 5 1 1 5151
0 5153 7 1 2 59786 73737
0 5154 5 2 1 5153
0 5155 7 1 2 82218 73636
0 5156 5 2 1 5155
0 5157 7 1 2 72153 82220
0 5158 5 1 1 5157
0 5159 7 1 2 74197 73628
0 5160 5 1 1 5159
0 5161 7 1 2 5158 5160
0 5162 7 1 2 5152 5161
0 5163 5 1 1 5162
0 5164 7 1 2 60774 5163
0 5165 5 1 1 5164
0 5166 7 1 2 72177 82221
0 5167 5 1 1 5166
0 5168 7 5 2 67471 74814
0 5169 5 2 1 82222
0 5170 7 1 2 70240 78236
0 5171 5 1 1 5170
0 5172 7 1 2 82227 5171
0 5173 5 1 1 5172
0 5174 7 1 2 5167 5173
0 5175 5 1 1 5174
0 5176 7 1 2 67001 5175
0 5177 5 1 1 5176
0 5178 7 1 2 5165 5177
0 5179 5 1 1 5178
0 5180 7 1 2 59265 5179
0 5181 5 1 1 5180
0 5182 7 9 2 67472 69171
0 5183 5 2 1 82229
0 5184 7 1 2 66154 82230
0 5185 5 1 1 5184
0 5186 7 1 2 73723 5185
0 5187 5 1 1 5186
0 5188 7 1 2 59787 5187
0 5189 5 1 1 5188
0 5190 7 2 2 60063 73919
0 5191 7 1 2 69294 82240
0 5192 5 1 1 5191
0 5193 7 1 2 5189 5192
0 5194 5 1 1 5193
0 5195 7 1 2 76042 5194
0 5196 5 1 1 5195
0 5197 7 1 2 74888 82241
0 5198 5 1 1 5197
0 5199 7 2 2 73724 82219
0 5200 5 1 1 82242
0 5201 7 4 2 67002 73431
0 5202 7 1 2 5200 82244
0 5203 5 1 1 5202
0 5204 7 1 2 5198 5203
0 5205 5 1 1 5204
0 5206 7 1 2 69090 5205
0 5207 5 1 1 5206
0 5208 7 2 2 73395 73738
0 5209 5 1 1 82248
0 5210 7 1 2 67829 5209
0 5211 7 1 2 5207 5210
0 5212 7 1 2 5196 5211
0 5213 7 1 2 5181 5212
0 5214 7 1 2 5147 5213
0 5215 5 1 1 5214
0 5216 7 3 2 64654 73035
0 5217 5 5 1 82250
0 5218 7 1 2 62495 82251
0 5219 5 1 1 5218
0 5220 7 1 2 60064 5219
0 5221 5 1 1 5220
0 5222 7 1 2 70002 5221
0 5223 5 1 1 5222
0 5224 7 21 2 59788 67473
0 5225 5 12 1 82258
0 5226 7 1 2 64877 82279
0 5227 5 2 1 5226
0 5228 7 1 2 72066 82291
0 5229 7 1 2 5223 5228
0 5230 5 1 1 5229
0 5231 7 4 2 77647 69450
0 5232 5 3 1 82293
0 5233 7 1 2 80710 82297
0 5234 5 1 1 5233
0 5235 7 12 2 64219 62222
0 5236 5 2 1 82300
0 5237 7 2 2 69363 82301
0 5238 5 14 1 82314
0 5239 7 1 2 74579 82316
0 5240 5 3 1 5239
0 5241 7 1 2 82330 82280
0 5242 5 1 1 5241
0 5243 7 1 2 60065 5242
0 5244 5 1 1 5243
0 5245 7 1 2 5234 5244
0 5246 7 1 2 5230 5245
0 5247 5 1 1 5246
0 5248 7 1 2 61205 5247
0 5249 5 1 1 5248
0 5250 7 2 2 80612 82259
0 5251 5 1 1 82333
0 5252 7 1 2 80924 82334
0 5253 5 1 1 5252
0 5254 7 1 2 62837 5253
0 5255 7 1 2 5249 5254
0 5256 5 1 1 5255
0 5257 7 1 2 68237 5256
0 5258 7 1 2 5215 5257
0 5259 5 1 1 5258
0 5260 7 15 2 67474 77881
0 5261 5 6 1 82335
0 5262 7 3 2 70581 73001
0 5263 5 1 1 82356
0 5264 7 1 2 82336 82357
0 5265 7 1 2 80222 5264
0 5266 5 1 1 5265
0 5267 7 1 2 5259 5266
0 5268 5 1 1 5267
0 5269 7 1 2 81748 5268
0 5270 5 1 1 5269
0 5271 7 1 2 5114 5270
0 5272 5 1 1 5271
0 5273 7 1 2 79505 5272
0 5274 5 1 1 5273
0 5275 7 2 2 64878 60229
0 5276 5 1 1 82359
0 5277 7 17 2 62016 62838
0 5278 5 10 1 82361
0 5279 7 2 2 74358 82362
0 5280 7 2 2 82360 82388
0 5281 5 1 1 82390
0 5282 7 1 2 71064 82391
0 5283 5 1 1 5282
0 5284 7 31 2 66387 67830
0 5285 5 3 1 82392
0 5286 7 2 2 73658 82393
0 5287 5 2 1 82426
0 5288 7 1 2 64417 72747
0 5289 7 1 2 82427 5288
0 5290 5 1 1 5289
0 5291 7 1 2 5283 5290
0 5292 5 1 1 5291
0 5293 7 1 2 65788 5292
0 5294 5 1 1 5293
0 5295 7 3 2 65094 82394
0 5296 7 2 2 70225 74821
0 5297 7 1 2 71477 72178
0 5298 5 2 1 5297
0 5299 7 2 2 75802 82435
0 5300 5 2 1 82437
0 5301 7 1 2 82438 74706
0 5302 5 1 1 5301
0 5303 7 1 2 82433 5302
0 5304 5 1 1 5303
0 5305 7 2 2 61206 81507
0 5306 5 1 1 82441
0 5307 7 1 2 73541 82442
0 5308 5 1 1 5307
0 5309 7 1 2 5304 5308
0 5310 5 1 1 5309
0 5311 7 1 2 82430 5310
0 5312 5 1 1 5311
0 5313 7 1 2 5294 5312
0 5314 5 1 1 5313
0 5315 7 1 2 62496 5314
0 5316 5 1 1 5315
0 5317 7 2 2 65789 73605
0 5318 5 2 1 82443
0 5319 7 1 2 74406 82445
0 5320 5 3 1 5319
0 5321 7 1 2 64418 82447
0 5322 5 2 1 5321
0 5323 7 2 2 77280 82450
0 5324 5 2 1 82452
0 5325 7 8 2 60066 67831
0 5326 5 3 1 82456
0 5327 7 1 2 82020 82457
0 5328 7 1 2 82454 5327
0 5329 5 1 1 5328
0 5330 7 5 2 62017 69150
0 5331 5 3 1 82467
0 5332 7 1 2 80137 79061
0 5333 7 1 2 82468 5332
0 5334 5 1 1 5333
0 5335 7 1 2 5329 5334
0 5336 5 1 1 5335
0 5337 7 1 2 69771 5336
0 5338 5 1 1 5337
0 5339 7 2 2 59789 78410
0 5340 5 1 1 82475
0 5341 7 1 2 67475 70395
0 5342 5 1 1 5341
0 5343 7 1 2 5340 5342
0 5344 5 1 1 5343
0 5345 7 1 2 59266 5344
0 5346 5 1 1 5345
0 5347 7 2 2 64655 74115
0 5348 5 4 1 82477
0 5349 7 1 2 69342 82479
0 5350 5 1 1 5349
0 5351 7 1 2 82281 5350
0 5352 7 1 2 5346 5351
0 5353 5 1 1 5352
0 5354 7 1 2 72067 5353
0 5355 5 1 1 5354
0 5356 7 1 2 78420 82260
0 5357 5 1 1 5356
0 5358 7 1 2 64656 1618
0 5359 5 3 1 5358
0 5360 7 1 2 69388 82483
0 5361 5 1 1 5360
0 5362 7 2 2 67221 74889
0 5363 5 1 1 82486
0 5364 7 2 2 60775 74088
0 5365 5 4 1 82488
0 5366 7 11 2 59267 59790
0 5367 5 2 1 82494
0 5368 7 1 2 82490 82505
0 5369 7 1 2 5363 5368
0 5370 7 1 2 5361 5369
0 5371 5 1 1 5370
0 5372 7 1 2 71687 5371
0 5373 5 1 1 5372
0 5374 7 1 2 5357 5373
0 5375 7 1 2 5355 5374
0 5376 5 1 1 5375
0 5377 7 3 2 62839 75162
0 5378 5 1 1 82507
0 5379 7 1 2 70582 82508
0 5380 7 1 2 5376 5379
0 5381 5 1 1 5380
0 5382 7 1 2 5338 5381
0 5383 7 1 2 5316 5382
0 5384 5 1 1 5383
0 5385 7 1 2 63305 5384
0 5386 5 1 1 5385
0 5387 7 7 2 68238 75163
0 5388 7 4 2 67222 72565
0 5389 5 5 1 82517
0 5390 7 3 2 59791 82518
0 5391 5 1 1 82526
0 5392 7 1 2 81230 82527
0 5393 5 1 1 5392
0 5394 7 3 2 64220 61207
0 5395 7 3 2 60067 82529
0 5396 7 1 2 75899 76955
0 5397 7 1 2 82532 5396
0 5398 5 1 1 5397
0 5399 7 1 2 5393 5398
0 5400 5 1 1 5399
0 5401 7 1 2 62497 5400
0 5402 5 1 1 5401
0 5403 7 2 2 64419 77336
0 5404 7 2 2 79189 82535
0 5405 7 1 2 73606 82537
0 5406 5 1 1 5405
0 5407 7 1 2 5402 5406
0 5408 5 1 1 5407
0 5409 7 1 2 65959 5408
0 5410 5 1 1 5409
0 5411 7 4 2 67476 70020
0 5412 5 1 1 82539
0 5413 7 1 2 69889 81887
0 5414 5 1 1 5413
0 5415 7 1 2 81832 5414
0 5416 5 1 1 5415
0 5417 7 1 2 82540 5416
0 5418 5 1 1 5417
0 5419 7 1 2 5410 5418
0 5420 5 1 1 5419
0 5421 7 1 2 62018 5420
0 5422 5 1 1 5421
0 5423 7 1 2 67477 78838
0 5424 5 1 1 5423
0 5425 7 3 2 59449 76618
0 5426 5 1 1 82543
0 5427 7 2 2 69498 82544
0 5428 5 1 1 82546
0 5429 7 1 2 60868 82547
0 5430 5 1 1 5429
0 5431 7 1 2 5424 5430
0 5432 5 1 1 5431
0 5433 7 1 2 65960 5432
0 5434 5 1 1 5433
0 5435 7 1 2 76683 76533
0 5436 5 2 1 5435
0 5437 7 1 2 69499 73607
0 5438 5 1 1 5437
0 5439 7 1 2 73594 5438
0 5440 7 1 2 82548 5439
0 5441 5 1 1 5440
0 5442 7 1 2 64879 5441
0 5443 5 1 1 5442
0 5444 7 1 2 5434 5443
0 5445 5 1 1 5444
0 5446 7 1 2 59792 5445
0 5447 5 1 1 5446
0 5448 7 8 2 67223 71688
0 5449 5 1 1 82550
0 5450 7 7 2 69091 74162
0 5451 5 16 1 82558
0 5452 7 1 2 69500 82559
0 5453 5 1 1 5452
0 5454 7 1 2 5449 5453
0 5455 5 1 1 5454
0 5456 7 1 2 71626 77017
0 5457 7 1 2 5455 5456
0 5458 5 1 1 5457
0 5459 7 1 2 5447 5458
0 5460 5 1 1 5459
0 5461 7 1 2 76384 5460
0 5462 5 1 1 5461
0 5463 7 4 2 80295 80649
0 5464 7 1 2 71951 73904
0 5465 7 1 2 82581 5464
0 5466 5 1 1 5465
0 5467 7 1 2 5462 5466
0 5468 7 1 2 5422 5467
0 5469 5 1 1 5468
0 5470 7 1 2 62840 5469
0 5471 5 1 1 5470
0 5472 7 1 2 81320 82154
0 5473 5 1 1 5472
0 5474 7 1 2 5471 5473
0 5475 5 1 1 5474
0 5476 7 1 2 82510 5475
0 5477 5 1 1 5476
0 5478 7 1 2 5386 5477
0 5479 5 1 1 5478
0 5480 7 1 2 68828 5479
0 5481 5 1 1 5480
0 5482 7 7 2 59793 70583
0 5483 5 3 1 82585
0 5484 7 2 2 82586 82439
0 5485 7 22 2 61419 67478
0 5486 5 2 1 82597
0 5487 7 2 2 60230 82598
0 5488 5 1 1 82621
0 5489 7 5 2 67832 81007
0 5490 7 1 2 82622 82623
0 5491 7 1 2 82595 5490
0 5492 5 1 1 5491
0 5493 7 1 2 5481 5492
0 5494 5 1 1 5493
0 5495 7 1 2 81145 5494
0 5496 5 1 1 5495
0 5497 7 3 2 62019 77287
0 5498 5 3 1 82628
0 5499 7 1 2 60068 82631
0 5500 5 1 1 5499
0 5501 7 1 2 5500 82538
0 5502 5 1 1 5501
0 5503 7 2 2 60776 73681
0 5504 5 1 1 82634
0 5505 7 1 2 74287 5504
0 5506 5 2 1 5505
0 5507 7 1 2 59268 82636
0 5508 5 3 1 5507
0 5509 7 20 2 61000 67003
0 5510 5 4 1 82641
0 5511 7 1 2 70396 82661
0 5512 5 1 1 5511
0 5513 7 1 2 82638 5512
0 5514 5 1 1 5513
0 5515 7 1 2 74580 5514
0 5516 5 1 1 5515
0 5517 7 2 2 59794 73036
0 5518 5 3 1 82665
0 5519 7 1 2 82666 69442
0 5520 5 1 1 5519
0 5521 7 1 2 67004 69348
0 5522 5 2 1 5521
0 5523 7 10 2 64657 62020
0 5524 5 4 1 82672
0 5525 7 1 2 59269 82682
0 5526 7 1 2 82662 5525
0 5527 7 1 2 82670 5526
0 5528 5 1 1 5527
0 5529 7 1 2 5520 5528
0 5530 5 1 1 5529
0 5531 7 1 2 72068 5530
0 5532 5 1 1 5531
0 5533 7 2 2 59450 62021
0 5534 5 1 1 82686
0 5535 7 2 2 71414 82687
0 5536 5 1 1 82688
0 5537 7 1 2 5532 5536
0 5538 7 1 2 5516 5537
0 5539 5 1 1 5538
0 5540 7 1 2 70021 5539
0 5541 5 1 1 5540
0 5542 7 1 2 5502 5541
0 5543 5 1 1 5542
0 5544 7 1 2 68239 5543
0 5545 5 1 1 5544
0 5546 7 1 2 71478 82059
0 5547 5 1 1 5546
0 5548 7 1 2 81883 5547
0 5549 5 1 1 5548
0 5550 7 1 2 80664 5549
0 5551 5 1 1 5550
0 5552 7 1 2 5545 5551
0 5553 5 1 1 5552
0 5554 7 1 2 67479 5553
0 5555 5 1 1 5554
0 5556 7 1 2 60869 78523
0 5557 5 1 1 5556
0 5558 7 1 2 64880 70272
0 5559 5 1 1 5558
0 5560 7 1 2 5557 5559
0 5561 5 1 1 5560
0 5562 7 1 2 59270 5561
0 5563 5 1 1 5562
0 5564 7 1 2 65961 76971
0 5565 5 1 1 5564
0 5566 7 1 2 76020 5565
0 5567 5 1 1 5566
0 5568 7 1 2 60870 5567
0 5569 5 1 1 5568
0 5570 7 1 2 5563 5569
0 5571 5 1 1 5570
0 5572 7 1 2 67224 5571
0 5573 5 1 1 5572
0 5574 7 1 2 73184 81264
0 5575 5 1 1 5574
0 5576 7 1 2 5573 5575
0 5577 5 1 1 5576
0 5578 7 1 2 59451 5577
0 5579 5 1 1 5578
0 5580 7 1 2 81875 76016
0 5581 5 1 1 5580
0 5582 7 1 2 5579 5581
0 5583 5 1 1 5582
0 5584 7 1 2 77591 74147
0 5585 7 1 2 5583 5584
0 5586 5 1 1 5585
0 5587 7 1 2 72069 70005
0 5588 5 2 1 5587
0 5589 7 1 2 71689 82317
0 5590 5 1 1 5589
0 5591 7 1 2 82690 5590
0 5592 5 1 1 5591
0 5593 7 1 2 79905 5592
0 5594 5 1 1 5593
0 5595 7 3 2 72762 73780
0 5596 5 1 1 82692
0 5597 7 1 2 76956 81864
0 5598 7 1 2 82693 5597
0 5599 5 1 1 5598
0 5600 7 1 2 5594 5599
0 5601 5 1 1 5600
0 5602 7 1 2 70584 5601
0 5603 5 1 1 5602
0 5604 7 1 2 62841 5603
0 5605 7 1 2 5586 5604
0 5606 7 1 2 5555 5605
0 5607 5 1 1 5606
0 5608 7 5 2 61420 81384
0 5609 5 2 1 82695
0 5610 7 2 2 79739 82696
0 5611 5 2 1 82702
0 5612 7 1 2 79914 82434
0 5613 5 1 1 5612
0 5614 7 1 2 78508 77614
0 5615 5 1 1 5614
0 5616 7 1 2 5613 5615
0 5617 5 1 1 5616
0 5618 7 1 2 71479 5617
0 5619 5 1 1 5618
0 5620 7 2 2 80619 81578
0 5621 5 1 1 82706
0 5622 7 1 2 65790 75000
0 5623 5 1 1 5622
0 5624 7 1 2 5621 5623
0 5625 5 1 1 5624
0 5626 7 1 2 69772 5625
0 5627 5 1 1 5626
0 5628 7 4 2 59452 70122
0 5629 5 2 1 82708
0 5630 7 1 2 79906 74822
0 5631 7 1 2 82709 5630
0 5632 5 1 1 5631
0 5633 7 1 2 77621 5632
0 5634 5 1 1 5633
0 5635 7 1 2 60871 5634
0 5636 5 1 1 5635
0 5637 7 1 2 5627 5636
0 5638 7 1 2 5619 5637
0 5639 5 1 1 5638
0 5640 7 1 2 67225 5639
0 5641 5 1 1 5640
0 5642 7 3 2 74984 80711
0 5643 7 1 2 60069 74716
0 5644 5 7 1 5643
0 5645 7 1 2 71318 82717
0 5646 5 1 1 5645
0 5647 7 1 2 82714 5646
0 5648 5 1 1 5647
0 5649 7 1 2 80620 5061
0 5650 5 1 1 5649
0 5651 7 1 2 5648 5650
0 5652 5 1 1 5651
0 5653 7 1 2 65962 5652
0 5654 5 1 1 5653
0 5655 7 3 2 59453 66155
0 5656 5 1 1 82724
0 5657 7 3 2 59795 80703
0 5658 7 1 2 82725 82727
0 5659 7 1 2 71341 5658
0 5660 5 1 1 5659
0 5661 7 1 2 5654 5660
0 5662 7 1 2 5641 5661
0 5663 5 1 1 5662
0 5664 7 1 2 62498 5663
0 5665 5 1 1 5664
0 5666 7 1 2 74396 82707
0 5667 5 1 1 5666
0 5668 7 5 2 69773 69052
0 5669 5 4 1 82730
0 5670 7 2 2 73970 73905
0 5671 5 1 1 82739
0 5672 7 1 2 82731 82740
0 5673 5 1 1 5672
0 5674 7 1 2 5667 5673
0 5675 5 1 1 5674
0 5676 7 1 2 64420 5675
0 5677 5 1 1 5676
0 5678 7 4 2 64658 76081
0 5679 5 3 1 82741
0 5680 7 1 2 77615 82742
0 5681 5 1 1 5680
0 5682 7 1 2 80645 74958
0 5683 5 1 1 5682
0 5684 7 1 2 5681 5683
0 5685 5 1 1 5684
0 5686 7 1 2 72540 5685
0 5687 5 1 1 5686
0 5688 7 1 2 67833 5687
0 5689 7 1 2 5677 5688
0 5690 7 1 2 5665 5689
0 5691 5 1 1 5690
0 5692 7 1 2 82703 5691
0 5693 7 1 2 5607 5692
0 5694 5 1 1 5693
0 5695 7 1 2 66156 70397
0 5696 5 1 1 5695
0 5697 7 1 2 82639 5696
0 5698 5 1 1 5697
0 5699 7 1 2 82261 5698
0 5700 5 1 1 5699
0 5701 7 3 2 62223 76899
0 5702 5 1 1 82748
0 5703 7 1 2 76088 82749
0 5704 5 1 1 5703
0 5705 7 1 2 70123 74116
0 5706 7 1 2 5704 5705
0 5707 5 1 1 5706
0 5708 7 1 2 5700 5707
0 5709 5 1 1 5708
0 5710 7 1 2 72070 5709
0 5711 5 1 1 5710
0 5712 7 1 2 76473 78326
0 5713 5 1 1 5712
0 5714 7 1 2 80467 77133
0 5715 5 1 1 5714
0 5716 7 1 2 73637 5715
0 5717 5 1 1 5716
0 5718 7 1 2 74581 5717
0 5719 5 1 1 5718
0 5720 7 1 2 61208 78230
0 5721 5 1 1 5720
0 5722 7 1 2 73682 78217
0 5723 5 1 1 5722
0 5724 7 1 2 74386 5723
0 5725 5 1 1 5724
0 5726 7 1 2 59796 5725
0 5727 5 1 1 5726
0 5728 7 1 2 5721 5727
0 5729 7 1 2 5719 5728
0 5730 7 1 2 5713 5729
0 5731 7 1 2 5711 5730
0 5732 5 1 1 5731
0 5733 7 1 2 75468 5732
0 5734 5 1 1 5733
0 5735 7 1 2 67480 74317
0 5736 5 1 1 5735
0 5737 7 1 2 74427 5736
0 5738 5 1 1 5737
0 5739 7 5 2 61209 75247
0 5740 5 1 1 82751
0 5741 7 1 2 73396 82752
0 5742 7 1 2 5738 5741
0 5743 5 1 1 5742
0 5744 7 1 2 5734 5743
0 5745 5 1 1 5744
0 5746 7 1 2 73472 5745
0 5747 5 1 1 5746
0 5748 7 3 2 63910 75469
0 5749 7 3 2 67481 76924
0 5750 7 1 2 70226 82759
0 5751 5 1 1 5750
0 5752 7 1 2 74979 5751
0 5753 5 1 1 5752
0 5754 7 1 2 69092 5753
0 5755 5 1 1 5754
0 5756 7 1 2 66157 78223
0 5757 5 4 1 5756
0 5758 7 1 2 78339 82762
0 5759 5 1 1 5758
0 5760 7 3 2 61210 72071
0 5761 5 1 1 82766
0 5762 7 1 2 69890 82767
0 5763 5 1 1 5762
0 5764 7 1 2 81715 5763
0 5765 7 1 2 5759 5764
0 5766 5 1 1 5765
0 5767 7 1 2 60070 5766
0 5768 5 1 1 5767
0 5769 7 4 2 59797 69891
0 5770 5 5 1 82769
0 5771 7 1 2 71466 82710
0 5772 7 1 2 82770 5771
0 5773 5 1 1 5772
0 5774 7 1 2 70735 5773
0 5775 5 1 1 5774
0 5776 7 1 2 69295 5775
0 5777 5 1 1 5776
0 5778 7 7 2 59454 69389
0 5779 5 10 1 82778
0 5780 7 2 2 74435 82779
0 5781 5 15 1 82795
0 5782 7 1 2 64659 82797
0 5783 5 1 1 5782
0 5784 7 1 2 73659 69460
0 5785 7 1 2 5783 5784
0 5786 5 1 1 5785
0 5787 7 1 2 5777 5786
0 5788 7 1 2 5768 5787
0 5789 7 1 2 5755 5788
0 5790 5 1 1 5789
0 5791 7 1 2 82756 5790
0 5792 5 1 1 5791
0 5793 7 5 2 64660 75164
0 5794 5 1 1 82812
0 5795 7 6 2 81321 82813
0 5796 7 1 2 62022 82817
0 5797 7 1 2 70998 5796
0 5798 5 1 1 5797
0 5799 7 1 2 5792 5798
0 5800 5 1 1 5799
0 5801 7 1 2 62842 5800
0 5802 5 1 1 5801
0 5803 7 1 2 5747 5802
0 5804 5 1 1 5803
0 5805 7 1 2 63306 5804
0 5806 5 1 1 5805
0 5807 7 1 2 59798 70555
0 5808 5 2 1 5807
0 5809 7 2 2 70435 82823
0 5810 5 1 1 82825
0 5811 7 1 2 66158 82826
0 5812 5 1 1 5811
0 5813 7 1 2 61211 73147
0 5814 5 1 1 5813
0 5815 7 1 2 62499 5814
0 5816 7 1 2 5812 5815
0 5817 5 1 1 5816
0 5818 7 1 2 77288 81672
0 5819 5 1 1 5818
0 5820 7 1 2 80142 72745
0 5821 5 1 1 5820
0 5822 7 1 2 66159 5821
0 5823 5 1 1 5822
0 5824 7 1 2 72729 5823
0 5825 5 1 1 5824
0 5826 7 1 2 67482 5825
0 5827 5 1 1 5826
0 5828 7 1 2 5819 5827
0 5829 7 1 2 5817 5828
0 5830 5 1 1 5829
0 5831 7 1 2 60231 5830
0 5832 5 1 1 5831
0 5833 7 1 2 72871 73608
0 5834 5 1 1 5833
0 5835 7 1 2 70363 73609
0 5836 5 1 1 5835
0 5837 7 1 2 72840 76096
0 5838 7 1 2 81240 5837
0 5839 5 1 1 5838
0 5840 7 1 2 5836 5839
0 5841 5 1 1 5840
0 5842 7 1 2 59455 5841
0 5843 5 1 1 5842
0 5844 7 1 2 5834 5843
0 5845 5 1 1 5844
0 5846 7 1 2 59799 72803
0 5847 7 1 2 5845 5846
0 5848 5 1 1 5847
0 5849 7 1 2 62843 5848
0 5850 7 1 2 5832 5849
0 5851 5 1 1 5850
0 5852 7 1 2 72541 772
0 5853 5 1 1 5852
0 5854 7 1 2 81641 77956
0 5855 5 1 1 5854
0 5856 7 1 2 5853 5855
0 5857 5 1 1 5856
0 5858 7 1 2 62023 5857
0 5859 5 1 1 5858
0 5860 7 1 2 81944 3166
0 5861 5 1 1 5860
0 5862 7 1 2 60232 5861
0 5863 5 1 1 5862
0 5864 7 1 2 67834 5863
0 5865 7 1 2 5859 5864
0 5866 5 1 1 5865
0 5867 7 1 2 61421 5866
0 5868 7 1 2 5851 5867
0 5869 5 1 1 5868
0 5870 7 9 2 60233 62844
0 5871 5 2 1 82827
0 5872 7 1 2 69329 82828
0 5873 5 1 1 5872
0 5874 7 4 2 61212 78242
0 5875 5 1 1 82838
0 5876 7 1 2 4945 75768
0 5877 5 1 1 5876
0 5878 7 1 2 82839 5877
0 5879 5 1 1 5878
0 5880 7 1 2 5873 5879
0 5881 5 1 1 5880
0 5882 7 1 2 60777 5881
0 5883 5 1 1 5882
0 5884 7 1 2 62845 81245
0 5885 5 1 1 5884
0 5886 7 6 2 67835 72814
0 5887 5 1 1 82842
0 5888 7 2 2 67005 69093
0 5889 5 2 1 82848
0 5890 7 1 2 82843 82849
0 5891 5 1 1 5890
0 5892 7 1 2 5885 5891
0 5893 5 1 1 5892
0 5894 7 1 2 67483 5893
0 5895 5 1 1 5894
0 5896 7 1 2 5883 5895
0 5897 5 1 1 5896
0 5898 7 1 2 59271 5897
0 5899 5 1 1 5898
0 5900 7 1 2 69390 82829
0 5901 5 1 1 5900
0 5902 7 1 2 78411 82844
0 5903 5 1 1 5902
0 5904 7 1 2 5901 5903
0 5905 5 1 1 5904
0 5906 7 1 2 60872 5905
0 5907 5 1 1 5906
0 5908 7 4 2 67006 78364
0 5909 5 1 1 82852
0 5910 7 1 2 65095 80634
0 5911 7 1 2 82853 5910
0 5912 5 2 1 5911
0 5913 7 1 2 5907 82856
0 5914 5 1 1 5913
0 5915 7 1 2 67484 5914
0 5916 5 1 1 5915
0 5917 7 1 2 5899 5916
0 5918 5 1 1 5917
0 5919 7 1 2 59456 5918
0 5920 5 1 1 5919
0 5921 7 1 2 70398 82845
0 5922 5 1 1 5921
0 5923 7 9 2 67007 62846
0 5924 5 1 1 82858
0 5925 7 3 2 60234 60778
0 5926 7 2 2 82859 82867
0 5927 5 1 1 82870
0 5928 7 1 2 5922 5927
0 5929 5 1 1 5928
0 5930 7 1 2 59272 5929
0 5931 5 1 1 5930
0 5932 7 1 2 82857 5931
0 5933 5 1 1 5932
0 5934 7 1 2 69461 5933
0 5935 5 1 1 5934
0 5936 7 1 2 5920 5935
0 5937 5 1 1 5936
0 5938 7 4 2 59800 66388
0 5939 7 1 2 60071 82872
0 5940 7 1 2 5937 5939
0 5941 5 1 1 5940
0 5942 7 1 2 5869 5941
0 5943 5 1 1 5942
0 5944 7 1 2 81008 5943
0 5945 5 1 1 5944
0 5946 7 1 2 5806 5945
0 5947 5 1 1 5946
0 5948 7 1 2 80837 5947
0 5949 5 1 1 5948
0 5950 7 1 2 5694 5949
0 5951 7 1 2 5496 5950
0 5952 7 1 2 5274 5951
0 5953 5 1 1 5952
0 5954 7 1 2 63635 5953
0 5955 5 1 1 5954
0 5956 7 1 2 64881 3387
0 5957 5 1 1 5956
0 5958 7 1 2 66160 5957
0 5959 5 1 1 5958
0 5960 7 1 2 79997 75737
0 5961 5 1 1 5960
0 5962 7 1 2 67836 5961
0 5963 7 1 2 5959 5962
0 5964 5 1 1 5963
0 5965 7 2 2 70124 71480
0 5966 7 1 2 74582 82876
0 5967 5 1 1 5966
0 5968 7 2 2 72072 70227
0 5969 5 2 1 82878
0 5970 7 1 2 62847 82880
0 5971 7 1 2 5967 5970
0 5972 5 1 1 5971
0 5973 7 1 2 67226 5972
0 5974 7 1 2 5964 5973
0 5975 5 1 1 5974
0 5976 7 1 2 64421 80077
0 5977 5 2 1 5976
0 5978 7 4 2 72831 82882
0 5979 7 3 2 62848 70125
0 5980 5 1 1 82888
0 5981 7 1 2 59273 77390
0 5982 5 1 1 5981
0 5983 7 1 2 5980 5982
0 5984 5 1 1 5983
0 5985 7 1 2 82884 5984
0 5986 5 1 1 5985
0 5987 7 3 2 59274 72073
0 5988 5 2 1 82891
0 5989 7 1 2 82889 82892
0 5990 5 1 1 5989
0 5991 7 1 2 66161 78302
0 5992 5 1 1 5991
0 5993 7 1 2 5990 5992
0 5994 5 1 1 5993
0 5995 7 1 2 69391 5994
0 5996 5 1 1 5995
0 5997 7 1 2 5986 5996
0 5998 5 1 1 5997
0 5999 7 1 2 59801 5998
0 6000 5 1 1 5999
0 6001 7 5 2 61213 78121
0 6002 5 3 1 82896
0 6003 7 8 2 62224 73862
0 6004 5 1 1 82904
0 6005 7 1 2 82897 82905
0 6006 5 1 1 6005
0 6007 7 25 2 61214 67837
0 6008 5 16 1 82912
0 6009 7 1 2 66162 78143
0 6010 5 12 1 6009
0 6011 7 3 2 60072 82953
0 6012 5 1 1 82965
0 6013 7 1 2 82937 82966
0 6014 5 1 1 6013
0 6015 7 1 2 6006 6014
0 6016 7 1 2 6000 6015
0 6017 7 1 2 5975 6016
0 6018 5 1 1 6017
0 6019 7 1 2 67485 6018
0 6020 5 1 1 6019
0 6021 7 17 2 67227 62849
0 6022 7 4 2 67008 82968
0 6023 7 1 2 80454 82985
0 6024 5 1 1 6023
0 6025 7 7 2 59275 67838
0 6026 5 1 1 82989
0 6027 7 1 2 76619 82990
0 6028 5 2 1 6027
0 6029 7 1 2 6024 82996
0 6030 5 1 1 6029
0 6031 7 1 2 70126 6030
0 6032 5 1 1 6031
0 6033 7 6 2 60073 62850
0 6034 5 2 1 82998
0 6035 7 1 2 60779 77391
0 6036 5 1 1 6035
0 6037 7 1 2 83004 6036
0 6038 5 1 1 6037
0 6039 7 1 2 59276 76578
0 6040 7 1 2 6038 6039
0 6041 5 1 1 6040
0 6042 7 1 2 6032 6041
0 6043 5 1 1 6042
0 6044 7 1 2 60873 6043
0 6045 5 1 1 6044
0 6046 7 7 2 62851 70585
0 6047 7 1 2 83006 70418
0 6048 5 1 1 6047
0 6049 7 2 2 64661 69733
0 6050 5 7 1 83013
0 6051 7 8 2 67839 70127
0 6052 5 3 1 83022
0 6053 7 1 2 76620 83023
0 6054 7 1 2 83015 6053
0 6055 5 1 1 6054
0 6056 7 1 2 6048 6055
0 6057 7 1 2 6045 6056
0 6058 5 1 1 6057
0 6059 7 1 2 59457 6058
0 6060 5 1 1 6059
0 6061 7 7 2 62225 77412
0 6062 5 5 1 83033
0 6063 7 3 2 59277 71690
0 6064 7 1 2 82969 83045
0 6065 5 1 1 6064
0 6066 7 1 2 83040 6065
0 6067 5 1 1 6066
0 6068 7 1 2 59802 6067
0 6069 5 1 1 6068
0 6070 7 19 2 59458 67840
0 6071 5 2 1 83048
0 6072 7 3 2 60874 76621
0 6073 5 2 1 83069
0 6074 7 1 2 83049 83070
0 6075 5 1 1 6074
0 6076 7 1 2 59278 82999
0 6077 7 1 2 74458 6076
0 6078 5 1 1 6077
0 6079 7 1 2 6075 6078
0 6080 7 1 2 6069 6079
0 6081 5 1 1 6080
0 6082 7 1 2 61215 6081
0 6083 5 1 1 6082
0 6084 7 2 2 73720 78862
0 6085 7 1 2 74583 83074
0 6086 5 1 1 6085
0 6087 7 1 2 6083 6086
0 6088 5 1 1 6087
0 6089 7 1 2 69392 6088
0 6090 5 1 1 6089
0 6091 7 1 2 60780 82986
0 6092 5 1 1 6091
0 6093 7 1 2 2615 6092
0 6094 5 1 1 6093
0 6095 7 1 2 61216 6094
0 6096 5 1 1 6095
0 6097 7 1 2 77383 82997
0 6098 5 1 1 6097
0 6099 7 1 2 80085 6098
0 6100 5 1 1 6099
0 6101 7 2 2 61217 82970
0 6102 5 1 1 83076
0 6103 7 1 2 59803 78885
0 6104 5 1 1 6103
0 6105 7 1 2 6102 6104
0 6106 5 1 1 6105
0 6107 7 1 2 60875 6106
0 6108 5 1 1 6107
0 6109 7 1 2 6100 6108
0 6110 7 1 2 6096 6109
0 6111 5 1 1 6110
0 6112 7 1 2 60074 6111
0 6113 5 1 1 6112
0 6114 7 1 2 80089 71429
0 6115 5 1 1 6114
0 6116 7 1 2 61218 83034
0 6117 7 1 2 6115 6116
0 6118 5 1 1 6117
0 6119 7 1 2 6113 6118
0 6120 7 1 2 6090 6119
0 6121 7 1 2 6060 6120
0 6122 7 1 2 6020 6121
0 6123 5 1 1 6122
0 6124 7 1 2 68240 6123
0 6125 5 1 1 6124
0 6126 7 1 2 76570 69469
0 6127 5 1 1 6126
0 6128 7 1 2 59459 6127
0 6129 5 1 1 6128
0 6130 7 1 2 82083 6129
0 6131 5 1 1 6130
0 6132 7 1 2 60781 6131
0 6133 5 1 1 6132
0 6134 7 1 2 74584 74089
0 6135 5 1 1 6134
0 6136 7 1 2 6133 6135
0 6137 5 1 1 6136
0 6138 7 1 2 59279 6137
0 6139 5 1 1 6138
0 6140 7 1 2 67486 5120
0 6141 5 1 1 6140
0 6142 7 2 2 71415 75007
0 6143 5 1 1 83078
0 6144 7 1 2 6141 6143
0 6145 7 1 2 6139 6144
0 6146 5 1 1 6145
0 6147 7 1 2 67228 6146
0 6148 5 2 1 6147
0 6149 7 1 2 83080 5251
0 6150 5 1 1 6149
0 6151 7 1 2 73971 82913
0 6152 7 1 2 6150 6151
0 6153 5 1 1 6152
0 6154 7 1 2 6125 6153
0 6155 5 1 1 6154
0 6156 7 1 2 80389 6155
0 6157 5 1 1 6156
0 6158 7 1 2 76235 73397
0 6159 5 1 1 6158
0 6160 7 1 2 67487 6159
0 6161 5 1 1 6160
0 6162 7 1 2 59280 69443
0 6163 5 1 1 6162
0 6164 7 2 2 77650 6163
0 6165 7 1 2 74708 83082
0 6166 5 1 1 6165
0 6167 7 1 2 62500 6166
0 6168 5 1 1 6167
0 6169 7 1 2 6161 6168
0 6170 5 1 1 6169
0 6171 7 33 2 62852 63307
0 6172 5 5 1 83084
0 6173 7 1 2 81731 83085
0 6174 7 1 2 6170 6173
0 6175 5 1 1 6174
0 6176 7 1 2 6157 6175
0 6177 5 1 1 6176
0 6178 7 1 2 68585 6177
0 6179 5 1 1 6178
0 6180 7 1 2 69501 80712
0 6181 5 1 1 6180
0 6182 7 1 2 73939 6181
0 6183 5 1 1 6182
0 6184 7 1 2 67229 6183
0 6185 5 1 1 6184
0 6186 7 1 2 73424 6185
0 6187 5 1 1 6186
0 6188 7 2 2 78122 73906
0 6189 7 3 2 63308 83122
0 6190 5 1 1 83124
0 6191 7 1 2 6187 83125
0 6192 5 1 1 6191
0 6193 7 2 2 62501 82718
0 6194 5 1 1 83127
0 6195 7 2 2 73560 82691
0 6196 7 1 2 64882 83129
0 6197 5 1 1 6196
0 6198 7 1 2 6194 6197
0 6199 5 1 1 6198
0 6200 7 1 2 59804 81437
0 6201 5 1 1 6200
0 6202 7 1 2 80713 82318
0 6203 5 1 1 6202
0 6204 7 1 2 6201 6203
0 6205 7 1 2 6199 6204
0 6206 5 1 1 6205
0 6207 7 1 2 62853 6206
0 6208 5 1 1 6207
0 6209 7 2 2 76900 72825
0 6210 5 1 1 83131
0 6211 7 1 2 81411 83132
0 6212 5 1 1 6211
0 6213 7 4 2 67488 73535
0 6214 5 3 1 83133
0 6215 7 1 2 59805 83134
0 6216 5 1 1 6215
0 6217 7 1 2 67841 6216
0 6218 7 1 2 6212 6217
0 6219 5 1 1 6218
0 6220 7 1 2 6208 6219
0 6221 5 1 1 6220
0 6222 7 1 2 61219 6221
0 6223 5 1 1 6222
0 6224 7 1 2 80640 82987
0 6225 5 1 1 6224
0 6226 7 2 2 61220 74792
0 6227 5 1 1 83140
0 6228 7 1 2 2362 6227
0 6229 5 1 1 6228
0 6230 7 1 2 62854 6229
0 6231 5 1 1 6230
0 6232 7 3 2 61221 70512
0 6233 5 2 1 83142
0 6234 7 1 2 67842 83145
0 6235 7 1 2 78421 6234
0 6236 5 1 1 6235
0 6237 7 1 2 6231 6236
0 6238 5 1 1 6237
0 6239 7 1 2 67489 6238
0 6240 5 1 1 6239
0 6241 7 1 2 6225 6240
0 6242 5 1 1 6241
0 6243 7 1 2 74585 6242
0 6244 5 1 1 6243
0 6245 7 1 2 78340 74875
0 6246 5 1 1 6245
0 6247 7 1 2 82243 6246
0 6248 5 1 1 6247
0 6249 7 1 2 67843 6248
0 6250 5 1 1 6249
0 6251 7 1 2 69892 82971
0 6252 7 1 2 73757 6251
0 6253 5 1 1 6252
0 6254 7 1 2 6250 6253
0 6255 5 1 1 6254
0 6256 7 1 2 72074 6255
0 6257 5 1 1 6256
0 6258 7 1 2 80714 78422
0 6259 5 1 1 6258
0 6260 7 1 2 73425 6259
0 6261 5 1 1 6260
0 6262 7 1 2 77413 6261
0 6263 5 1 1 6262
0 6264 7 1 2 6257 6263
0 6265 7 1 2 6244 6264
0 6266 7 1 2 6223 6265
0 6267 5 1 1 6266
0 6268 7 1 2 68241 6267
0 6269 5 1 1 6268
0 6270 7 1 2 6192 6269
0 6271 5 1 1 6270
0 6272 7 9 2 63636 80838
0 6273 5 1 1 83147
0 6274 7 1 2 6271 83148
0 6275 5 1 1 6274
0 6276 7 1 2 6179 6275
0 6277 5 1 1 6276
0 6278 7 1 2 79506 6277
0 6279 5 1 1 6278
0 6280 7 4 2 60075 68586
0 6281 7 2 2 61422 75676
0 6282 5 2 1 83160
0 6283 7 1 2 82637 83161
0 6284 5 1 1 6283
0 6285 7 5 2 65096 75823
0 6286 5 2 1 83164
0 6287 7 1 2 77639 83165
0 6288 5 1 1 6287
0 6289 7 1 2 6284 6288
0 6290 5 1 1 6289
0 6291 7 1 2 82914 6290
0 6292 5 1 1 6291
0 6293 7 2 2 74397 77758
0 6294 5 1 1 83171
0 6295 7 1 2 76972 74359
0 6296 7 1 2 83172 6295
0 6297 5 1 1 6296
0 6298 7 1 2 6292 6297
0 6299 5 1 1 6298
0 6300 7 1 2 59281 6299
0 6301 5 1 1 6300
0 6302 7 3 2 71002 81043
0 6303 7 1 2 67230 83173
0 6304 5 1 1 6303
0 6305 7 1 2 65097 81200
0 6306 5 1 1 6305
0 6307 7 1 2 6304 6306
0 6308 5 1 1 6307
0 6309 7 1 2 60782 6308
0 6310 5 1 1 6309
0 6311 7 1 2 81472 82511
0 6312 5 1 1 6311
0 6313 7 1 2 6310 6312
0 6314 5 1 1 6313
0 6315 7 1 2 82915 6314
0 6316 5 1 1 6315
0 6317 7 1 2 6301 6316
0 6318 5 1 1 6317
0 6319 7 1 2 60876 6318
0 6320 5 1 1 6319
0 6321 7 2 2 68242 81431
0 6322 7 1 2 74725 82846
0 6323 7 1 2 83176 6322
0 6324 5 1 1 6323
0 6325 7 1 2 6320 6324
0 6326 5 1 1 6325
0 6327 7 1 2 59460 6326
0 6328 5 1 1 6327
0 6329 7 1 2 82512 82840
0 6330 7 1 2 70389 6329
0 6331 5 1 1 6330
0 6332 7 1 2 6328 6331
0 6333 5 1 1 6332
0 6334 7 1 2 59806 6333
0 6335 5 1 1 6334
0 6336 7 2 2 69502 75165
0 6337 7 21 2 59461 68243
0 6338 5 8 1 83180
0 6339 7 1 2 78243 83181
0 6340 7 1 2 83178 6339
0 6341 7 1 2 76377 6340
0 6342 5 1 1 6341
0 6343 7 1 2 6335 6342
0 6344 5 1 1 6343
0 6345 7 1 2 83156 6344
0 6346 5 1 1 6345
0 6347 7 2 2 59462 74890
0 6348 5 3 1 83209
0 6349 7 1 2 71481 83210
0 6350 5 1 1 6349
0 6351 7 1 2 82282 6350
0 6352 5 1 1 6351
0 6353 7 1 2 69094 6352
0 6354 5 1 1 6353
0 6355 7 1 2 76925 81710
0 6356 5 1 1 6355
0 6357 7 1 2 6354 6356
0 6358 5 1 1 6357
0 6359 7 6 2 70586 78733
0 6360 5 3 1 83214
0 6361 7 2 2 67844 83215
0 6362 7 1 2 6358 83223
0 6363 5 1 1 6362
0 6364 7 1 2 78635 78613
0 6365 5 3 1 6364
0 6366 7 1 2 64883 83225
0 6367 5 1 1 6366
0 6368 7 1 2 67490 6367
0 6369 5 1 1 6368
0 6370 7 1 2 66163 6369
0 6371 7 1 2 83081 6370
0 6372 5 1 1 6371
0 6373 7 1 2 73222 82210
0 6374 5 2 1 6373
0 6375 7 1 2 61222 83228
0 6376 5 1 1 6375
0 6377 7 1 2 63309 6376
0 6378 7 1 2 6372 6377
0 6379 5 1 1 6378
0 6380 7 3 2 76694 78027
0 6381 5 2 1 83230
0 6382 7 1 2 68244 83231
0 6383 5 1 1 6382
0 6384 7 2 2 80105 75706
0 6385 5 1 1 83235
0 6386 7 1 2 6383 6385
0 6387 5 1 1 6386
0 6388 7 1 2 64422 6387
0 6389 5 1 1 6388
0 6390 7 1 2 64662 73660
0 6391 5 1 1 6390
0 6392 7 1 2 76484 6391
0 6393 5 1 1 6392
0 6394 7 1 2 67009 6393
0 6395 5 1 1 6394
0 6396 7 1 2 76476 6395
0 6397 7 1 2 76471 6396
0 6398 5 1 1 6397
0 6399 7 1 2 63310 6398
0 6400 5 1 1 6399
0 6401 7 1 2 6389 6400
0 6402 5 2 1 6401
0 6403 7 1 2 62502 83237
0 6404 5 1 1 6403
0 6405 7 1 2 67845 6404
0 6406 7 1 2 6379 6405
0 6407 5 1 1 6406
0 6408 7 2 2 77592 76964
0 6409 5 1 1 83239
0 6410 7 2 2 63311 70128
0 6411 7 1 2 69095 73313
0 6412 5 1 1 6411
0 6413 7 11 2 67231 71416
0 6414 5 2 1 83243
0 6415 7 1 2 76991 73254
0 6416 5 1 1 6415
0 6417 7 1 2 83254 6416
0 6418 7 2 2 6412 6417
0 6419 5 1 1 83256
0 6420 7 1 2 70736 83257
0 6421 5 1 1 6420
0 6422 7 1 2 83241 6421
0 6423 5 1 1 6422
0 6424 7 1 2 6409 6423
0 6425 5 1 1 6424
0 6426 7 1 2 67491 6425
0 6427 5 2 1 6426
0 6428 7 3 2 67010 76622
0 6429 5 1 1 83260
0 6430 7 1 2 77593 83261
0 6431 5 2 1 6430
0 6432 7 2 2 81520 76836
0 6433 5 2 1 83265
0 6434 7 3 2 67011 80106
0 6435 7 1 2 70228 83269
0 6436 5 1 1 6435
0 6437 7 1 2 83267 6436
0 6438 5 1 1 6437
0 6439 7 1 2 60783 6438
0 6440 5 1 1 6439
0 6441 7 1 2 83263 6440
0 6442 5 1 1 6441
0 6443 7 1 2 72075 6442
0 6444 5 1 1 6443
0 6445 7 1 2 60784 76162
0 6446 5 1 1 6445
0 6447 7 1 2 76021 6446
0 6448 5 1 1 6447
0 6449 7 2 2 66164 80804
0 6450 7 1 2 6448 83272
0 6451 5 2 1 6450
0 6452 7 1 2 63312 80251
0 6453 5 1 1 6452
0 6454 7 1 2 83274 6453
0 6455 5 1 1 6454
0 6456 7 1 2 69444 6455
0 6457 5 1 1 6456
0 6458 7 1 2 6444 6457
0 6459 5 1 1 6458
0 6460 7 1 2 59282 6459
0 6461 5 1 1 6460
0 6462 7 2 2 60877 78412
0 6463 5 1 1 83276
0 6464 7 2 2 69393 83277
0 6465 5 1 1 83278
0 6466 7 2 2 76490 83279
0 6467 5 1 1 83280
0 6468 7 1 2 70129 83281
0 6469 5 1 1 6468
0 6470 7 1 2 73863 70402
0 6471 5 1 1 6470
0 6472 7 2 2 60076 6471
0 6473 5 1 1 83282
0 6474 7 1 2 61223 83283
0 6475 5 1 1 6474
0 6476 7 1 2 6469 6475
0 6477 5 1 1 6476
0 6478 7 1 2 63313 6477
0 6479 5 1 1 6478
0 6480 7 1 2 78843 5426
0 6481 5 1 1 6480
0 6482 7 1 2 77594 6481
0 6483 5 1 1 6482
0 6484 7 1 2 75004 6483
0 6485 5 1 1 6484
0 6486 7 1 2 72832 6485
0 6487 5 1 1 6486
0 6488 7 4 2 64663 74003
0 6489 5 5 1 83284
0 6490 7 1 2 64884 83288
0 6491 5 1 1 6490
0 6492 7 1 2 80072 76623
0 6493 5 1 1 6492
0 6494 7 1 2 6491 6493
0 6495 5 1 1 6494
0 6496 7 1 2 77595 6495
0 6497 5 1 1 6496
0 6498 7 2 2 6487 6497
0 6499 7 1 2 62855 83293
0 6500 7 1 2 6479 6499
0 6501 7 1 2 6461 6500
0 6502 7 1 2 83258 6501
0 6503 5 1 1 6502
0 6504 7 1 2 68587 6503
0 6505 7 1 2 6407 6504
0 6506 5 1 1 6505
0 6507 7 1 2 6363 6506
0 6508 5 1 1 6507
0 6509 7 1 2 61423 6508
0 6510 5 1 1 6509
0 6511 7 2 2 74985 77414
0 6512 5 1 1 83295
0 6513 7 1 2 74300 83296
0 6514 5 1 1 6513
0 6515 7 10 2 66389 67232
0 6516 5 6 1 83297
0 6517 7 2 2 69503 83298
0 6518 5 1 1 83313
0 6519 7 1 2 77759 83314
0 6520 5 1 1 6519
0 6521 7 1 2 6514 6520
0 6522 5 1 1 6521
0 6523 7 1 2 74198 83157
0 6524 7 1 2 6522 6523
0 6525 5 1 1 6524
0 6526 7 1 2 6510 6525
0 6527 5 1 1 6526
0 6528 7 1 2 60235 6527
0 6529 5 1 1 6528
0 6530 7 1 2 6346 6529
0 6531 5 1 1 6530
0 6532 7 1 2 81146 6531
0 6533 5 1 1 6532
0 6534 7 1 2 83270 77656
0 6535 5 1 1 6534
0 6536 7 1 2 83268 6535
0 6537 5 1 1 6536
0 6538 7 1 2 60785 6537
0 6539 5 1 1 6538
0 6540 7 1 2 6539 83264
0 6541 5 1 1 6540
0 6542 7 1 2 72076 6541
0 6543 5 1 1 6542
0 6544 7 1 2 146 82715
0 6545 5 1 1 6544
0 6546 7 1 2 83275 6545
0 6547 7 1 2 6543 6546
0 6548 5 1 1 6547
0 6549 7 1 2 59283 6548
0 6550 5 1 1 6549
0 6551 7 1 2 6467 6473
0 6552 5 1 1 6551
0 6553 7 1 2 74986 6552
0 6554 5 1 1 6553
0 6555 7 1 2 83294 6554
0 6556 7 1 2 6550 6555
0 6557 7 1 2 83259 6556
0 6558 5 1 1 6557
0 6559 7 1 2 65098 6558
0 6560 5 1 1 6559
0 6561 7 2 2 60878 72440
0 6562 5 2 1 83315
0 6563 7 1 2 62024 83317
0 6564 5 1 1 6563
0 6565 7 1 2 59284 69354
0 6566 7 1 2 6564 6565
0 6567 5 1 1 6566
0 6568 7 1 2 6465 6567
0 6569 5 1 1 6568
0 6570 7 1 2 59463 6569
0 6571 5 1 1 6570
0 6572 7 1 2 6571 82156
0 6573 5 3 1 6572
0 6574 7 3 2 63314 73398
0 6575 7 1 2 73158 83322
0 6576 7 1 2 83319 6575
0 6577 5 1 1 6576
0 6578 7 1 2 6560 6577
0 6579 5 1 1 6578
0 6580 7 1 2 68588 6579
0 6581 5 1 1 6580
0 6582 7 6 2 62503 74004
0 6583 5 8 1 83325
0 6584 7 1 2 3383 83331
0 6585 5 1 1 6584
0 6586 7 1 2 77121 83211
0 6587 5 1 1 6586
0 6588 7 1 2 72853 6587
0 6589 5 1 1 6588
0 6590 7 8 2 59464 67492
0 6591 5 8 1 83339
0 6592 7 1 2 72874 83347
0 6593 5 1 1 6592
0 6594 7 1 2 59807 6593
0 6595 5 1 1 6594
0 6596 7 1 2 6589 6595
0 6597 7 1 2 6585 6596
0 6598 5 1 1 6597
0 6599 7 6 2 60236 63637
0 6600 7 1 2 80781 83355
0 6601 7 1 2 6598 6600
0 6602 5 1 1 6601
0 6603 7 1 2 6581 6602
0 6604 5 1 1 6603
0 6605 7 1 2 66390 6604
0 6606 5 1 1 6605
0 6607 7 1 2 67233 82489
0 6608 5 1 1 6607
0 6609 7 1 2 64885 6608
0 6610 5 1 1 6609
0 6611 7 1 2 71417 6610
0 6612 5 1 1 6611
0 6613 7 2 2 67234 73758
0 6614 5 1 1 83361
0 6615 7 1 2 6612 6614
0 6616 5 1 1 6615
0 6617 7 1 2 59465 6616
0 6618 5 1 1 6617
0 6619 7 4 2 59285 71349
0 6620 5 2 1 83363
0 6621 7 1 2 69394 83364
0 6622 5 1 1 6621
0 6623 7 1 2 66165 6622
0 6624 5 1 1 6623
0 6625 7 1 2 80715 6624
0 6626 5 1 1 6625
0 6627 7 1 2 6618 6626
0 6628 5 1 1 6627
0 6629 7 1 2 63315 6628
0 6630 5 1 1 6629
0 6631 7 1 2 77596 71366
0 6632 7 1 2 74891 6631
0 6633 5 1 1 6632
0 6634 7 1 2 6630 6633
0 6635 5 1 1 6634
0 6636 7 1 2 60237 6635
0 6637 5 1 1 6636
0 6638 7 1 2 80943 72808
0 6639 5 2 1 6638
0 6640 7 2 2 69893 71517
0 6641 5 1 1 83371
0 6642 7 1 2 63316 83372
0 6643 5 1 1 6642
0 6644 7 1 2 83369 6643
0 6645 5 1 1 6644
0 6646 7 1 2 59808 6645
0 6647 5 1 1 6646
0 6648 7 1 2 68245 79176
0 6649 5 1 1 6648
0 6650 7 4 2 59286 60238
0 6651 7 3 2 67493 83242
0 6652 7 1 2 83373 83377
0 6653 5 1 1 6652
0 6654 7 5 2 67235 73399
0 6655 7 1 2 81549 83380
0 6656 5 1 1 6655
0 6657 7 1 2 6653 6656
0 6658 5 1 1 6657
0 6659 7 1 2 69395 6658
0 6660 5 1 1 6659
0 6661 7 1 2 6649 6660
0 6662 7 1 2 6647 6661
0 6663 5 1 1 6662
0 6664 7 1 2 72077 6663
0 6665 5 1 1 6664
0 6666 7 2 2 59287 81550
0 6667 5 1 1 83385
0 6668 7 1 2 73400 83386
0 6669 5 1 1 6668
0 6670 7 1 2 60239 83378
0 6671 5 1 1 6670
0 6672 7 1 2 6669 6671
0 6673 5 1 1 6672
0 6674 7 1 2 73128 6673
0 6675 5 1 1 6674
0 6676 7 2 2 60240 70229
0 6677 5 1 1 83387
0 6678 7 1 2 80107 83388
0 6679 5 1 1 6678
0 6680 7 1 2 77597 73610
0 6681 7 1 2 80800 6680
0 6682 5 1 1 6681
0 6683 7 1 2 6679 6682
0 6684 7 1 2 6675 6683
0 6685 5 1 1 6684
0 6686 7 1 2 72833 6685
0 6687 5 1 1 6686
0 6688 7 2 2 71418 72737
0 6689 5 2 1 83389
0 6690 7 1 2 65099 83391
0 6691 5 2 1 6690
0 6692 7 1 2 74987 83365
0 6693 5 1 1 6692
0 6694 7 1 2 4343 6693
0 6695 5 1 1 6694
0 6696 7 1 2 69396 6695
0 6697 5 1 1 6696
0 6698 7 1 2 67236 81551
0 6699 5 1 1 6698
0 6700 7 1 2 6697 6699
0 6701 5 1 1 6700
0 6702 7 1 2 83393 6701
0 6703 5 1 1 6702
0 6704 7 16 2 60241 63317
0 6705 5 8 1 83395
0 6706 7 2 2 83332 83396
0 6707 7 1 2 70130 83419
0 6708 5 1 1 6707
0 6709 7 1 2 59466 74398
0 6710 5 1 1 6709
0 6711 7 1 2 73621 6710
0 6712 5 2 1 6711
0 6713 7 5 2 59288 68246
0 6714 5 1 1 83423
0 6715 7 1 2 72804 83424
0 6716 7 1 2 83421 6715
0 6717 5 1 1 6716
0 6718 7 1 2 6708 6717
0 6719 5 1 1 6718
0 6720 7 1 2 80086 6719
0 6721 5 1 1 6720
0 6722 7 1 2 73999 74256
0 6723 5 1 1 6722
0 6724 7 1 2 6667 6723
0 6725 5 1 1 6724
0 6726 7 6 2 60879 73401
0 6727 5 1 1 83428
0 6728 7 1 2 70273 83429
0 6729 5 1 1 6728
0 6730 7 1 2 65100 6729
0 6731 5 1 1 6730
0 6732 7 1 2 6725 6731
0 6733 5 1 1 6732
0 6734 7 3 2 59289 83397
0 6735 5 1 1 83434
0 6736 7 1 2 78398 83435
0 6737 5 1 1 6736
0 6738 7 1 2 83370 6737
0 6739 5 1 1 6738
0 6740 7 1 2 74586 69397
0 6741 7 1 2 6739 6740
0 6742 5 1 1 6741
0 6743 7 1 2 6733 6742
0 6744 7 1 2 6721 6743
0 6745 7 1 2 6703 6744
0 6746 7 1 2 6687 6745
0 6747 7 1 2 6665 6746
0 6748 7 1 2 6637 6747
0 6749 5 1 1 6748
0 6750 7 1 2 61424 6749
0 6751 5 1 1 6750
0 6752 7 5 2 59467 81246
0 6753 7 1 2 73402 83437
0 6754 7 1 2 71383 6753
0 6755 5 1 1 6754
0 6756 7 1 2 6751 6755
0 6757 5 1 1 6756
0 6758 7 1 2 63638 6757
0 6759 5 1 1 6758
0 6760 7 1 2 62856 6759
0 6761 7 1 2 6606 6760
0 6762 5 1 1 6761
0 6763 7 9 2 65101 68589
0 6764 7 1 2 83442 83238
0 6765 5 1 1 6764
0 6766 7 1 2 78734 82596
0 6767 5 1 1 6766
0 6768 7 1 2 6765 6767
0 6769 5 1 1 6768
0 6770 7 1 2 66391 6769
0 6771 5 1 1 6770
0 6772 7 1 2 81888 71482
0 6773 5 1 1 6772
0 6774 7 3 2 81833 6773
0 6775 5 3 1 83451
0 6776 7 5 2 64886 75540
0 6777 5 2 1 83457
0 6778 7 5 2 66166 75541
0 6779 5 4 1 83464
0 6780 7 8 2 83462 83469
0 6781 5 6 1 83473
0 6782 7 11 2 75248 83474
0 6783 5 4 1 83487
0 6784 7 1 2 83454 83488
0 6785 5 1 1 6784
0 6786 7 1 2 80271 6785
0 6787 5 1 1 6786
0 6788 7 1 2 79030 6787
0 6789 5 1 1 6788
0 6790 7 1 2 62504 6789
0 6791 7 1 2 6771 6790
0 6792 5 1 1 6791
0 6793 7 1 2 64664 69349
0 6794 5 1 1 6793
0 6795 7 1 2 62025 6794
0 6796 5 1 1 6795
0 6797 7 1 2 82640 6796
0 6798 5 1 1 6797
0 6799 7 1 2 83489 6798
0 6800 5 1 1 6799
0 6801 7 3 2 61425 73002
0 6802 5 1 1 83502
0 6803 7 1 2 78797 83503
0 6804 5 1 1 6803
0 6805 7 1 2 6800 6804
0 6806 5 1 1 6805
0 6807 7 1 2 63318 6806
0 6808 5 1 1 6807
0 6809 7 2 2 64665 78343
0 6810 5 1 1 83505
0 6811 7 5 2 60077 81593
0 6812 5 2 1 83507
0 6813 7 1 2 75166 83508
0 6814 7 1 2 6810 6813
0 6815 5 1 1 6814
0 6816 7 1 2 6808 6815
0 6817 5 1 1 6816
0 6818 7 1 2 63639 6817
0 6819 5 1 1 6818
0 6820 7 61 2 63319 68590
0 6821 7 3 2 79551 83514
0 6822 7 1 2 72453 80793
0 6823 7 1 2 83575 6822
0 6824 5 1 1 6823
0 6825 7 1 2 6819 6824
0 6826 5 1 1 6825
0 6827 7 1 2 72078 6826
0 6828 5 1 1 6827
0 6829 7 14 2 67012 63640
0 6830 7 4 2 60078 75249
0 6831 5 2 1 83592
0 6832 7 6 2 59290 67237
0 6833 5 4 1 83598
0 6834 7 3 2 80455 83599
0 6835 7 1 2 74686 83608
0 6836 5 1 1 6835
0 6837 7 1 2 77671 6836
0 6838 5 1 1 6837
0 6839 7 1 2 83593 6838
0 6840 5 1 1 6839
0 6841 7 2 2 62226 75470
0 6842 5 1 1 83611
0 6843 7 1 2 6840 6842
0 6844 5 1 1 6843
0 6845 7 1 2 71691 6844
0 6846 5 1 1 6845
0 6847 7 4 2 61426 78798
0 6848 7 1 2 83613 82055
0 6849 5 1 1 6848
0 6850 7 1 2 6846 6849
0 6851 5 1 1 6850
0 6852 7 1 2 83578 6851
0 6853 5 1 1 6852
0 6854 7 15 2 68591 75167
0 6855 7 1 2 66167 80716
0 6856 5 1 1 6855
0 6857 7 1 2 69774 81663
0 6858 5 1 1 6857
0 6859 7 1 2 6856 6858
0 6860 5 1 1 6859
0 6861 7 1 2 83617 6860
0 6862 5 1 1 6861
0 6863 7 1 2 6853 6862
0 6864 5 1 1 6863
0 6865 7 1 2 63320 6864
0 6866 5 1 1 6865
0 6867 7 9 2 62026 63641
0 6868 7 1 2 83490 83632
0 6869 5 2 1 6868
0 6870 7 2 2 80468 83618
0 6871 5 1 1 83643
0 6872 7 1 2 83641 6871
0 6873 5 1 1 6872
0 6874 7 1 2 69894 6873
0 6875 5 1 1 6874
0 6876 7 8 2 66168 68592
0 6877 7 1 2 83645 83179
0 6878 5 1 1 6877
0 6879 7 1 2 83642 6878
0 6880 5 1 1 6879
0 6881 7 1 2 67238 6880
0 6882 5 1 1 6881
0 6883 7 1 2 6875 6882
0 6884 5 1 1 6883
0 6885 7 1 2 63321 6884
0 6886 5 1 1 6885
0 6887 7 1 2 65102 78413
0 6888 5 1 1 6887
0 6889 7 2 2 65103 67013
0 6890 5 3 1 83653
0 6891 7 1 2 3665 83655
0 6892 5 1 1 6891
0 6893 7 1 2 59291 6892
0 6894 5 1 1 6893
0 6895 7 1 2 6888 6894
0 6896 5 1 1 6895
0 6897 7 10 2 61224 63642
0 6898 7 1 2 83658 75861
0 6899 7 1 2 6896 6898
0 6900 5 1 1 6899
0 6901 7 1 2 6886 6900
0 6902 5 1 1 6901
0 6903 7 1 2 74587 6902
0 6904 5 1 1 6903
0 6905 7 1 2 67494 6904
0 6906 7 1 2 6866 6905
0 6907 7 1 2 6828 6906
0 6908 5 1 1 6907
0 6909 7 1 2 6792 6908
0 6910 5 1 1 6909
0 6911 7 9 2 60242 79197
0 6912 5 3 1 83668
0 6913 7 1 2 74382 83669
0 6914 5 1 1 6913
0 6915 7 5 2 76251 78472
0 6916 5 4 1 83680
0 6917 7 1 2 73549 83644
0 6918 7 1 2 83681 6917
0 6919 5 1 1 6918
0 6920 7 1 2 6914 6919
0 6921 5 1 1 6920
0 6922 7 1 2 63322 6921
0 6923 5 1 1 6922
0 6924 7 1 2 67846 6923
0 6925 7 1 2 6910 6924
0 6926 5 1 1 6925
0 6927 7 1 2 80839 6926
0 6928 7 1 2 6762 6927
0 6929 5 1 1 6928
0 6930 7 1 2 67495 130
0 6931 5 1 1 6930
0 6932 7 1 2 69336 6931
0 6933 5 1 1 6932
0 6934 7 1 2 59468 6933
0 6935 5 1 1 6934
0 6936 7 1 2 67496 70390
0 6937 5 1 1 6936
0 6938 7 1 2 6935 6937
0 6939 5 1 1 6938
0 6940 7 1 2 59809 6939
0 6941 5 1 1 6940
0 6942 7 3 2 69504 83340
0 6943 5 1 1 83689
0 6944 7 1 2 81457 83690
0 6945 5 2 1 6944
0 6946 7 1 2 6941 83692
0 6947 5 1 1 6946
0 6948 7 15 2 65327 61427
0 6949 5 14 1 83694
0 6950 7 6 2 66628 83695
0 6951 7 28 2 67847 68247
0 6952 5 7 1 83729
0 6953 7 5 2 68593 83730
0 6954 7 1 2 81790 83764
0 6955 7 1 2 83723 6954
0 6956 7 1 2 6947 6955
0 6957 5 1 1 6956
0 6958 7 1 2 63911 6957
0 6959 7 1 2 6929 6958
0 6960 7 1 2 6533 6959
0 6961 7 1 2 6279 6960
0 6962 5 1 1 6961
0 6963 7 2 2 64666 69976
0 6964 5 2 1 83769
0 6965 7 3 2 72433 70442
0 6966 5 2 1 83773
0 6967 7 1 2 83771 83776
0 6968 5 1 1 6967
0 6969 7 1 2 65791 6968
0 6970 5 1 1 6969
0 6971 7 1 2 77333 6970
0 6972 5 1 1 6971
0 6973 7 1 2 67848 6972
0 6974 5 1 1 6973
0 6975 7 1 2 79952 82972
0 6976 5 1 1 6975
0 6977 7 1 2 6974 6976
0 6978 5 1 1 6977
0 6979 7 1 2 67014 6978
0 6980 5 1 1 6979
0 6981 7 1 2 62857 80215
0 6982 5 1 1 6981
0 6983 7 1 2 67849 74717
0 6984 5 1 1 6983
0 6985 7 1 2 67239 6984
0 6986 7 1 2 6982 6985
0 6987 5 1 1 6986
0 6988 7 9 2 59810 62858
0 6989 5 2 1 83778
0 6990 7 2 2 71692 83779
0 6991 5 1 1 83789
0 6992 7 1 2 6987 6991
0 6993 7 1 2 6980 6992
0 6994 5 1 1 6993
0 6995 7 1 2 62505 6994
0 6996 5 1 1 6995
0 6997 7 5 2 64221 77228
0 6998 5 2 1 83791
0 6999 7 2 2 72583 83796
0 7000 5 1 1 83798
0 7001 7 2 2 62859 76323
0 7002 5 9 1 83800
0 7003 7 3 2 65792 76624
0 7004 5 5 1 83811
0 7005 7 1 2 67850 83814
0 7006 5 4 1 7005
0 7007 7 2 2 83802 83819
0 7008 7 1 2 83799 83823
0 7009 5 1 1 7008
0 7010 7 1 2 78173 78636
0 7011 5 1 1 7010
0 7012 7 8 2 62506 69775
0 7013 7 1 2 64423 78286
0 7014 7 1 2 83825 7013
0 7015 5 1 1 7014
0 7016 7 1 2 7011 7015
0 7017 5 1 1 7016
0 7018 7 1 2 62227 7017
0 7019 5 1 1 7018
0 7020 7 1 2 7009 7019
0 7021 5 1 1 7020
0 7022 7 1 2 62027 7021
0 7023 5 1 1 7022
0 7024 7 1 2 64667 81623
0 7025 5 1 1 7024
0 7026 7 1 2 69053 73185
0 7027 5 1 1 7026
0 7028 7 1 2 7025 7027
0 7029 5 1 1 7028
0 7030 7 1 2 59469 7029
0 7031 5 1 1 7030
0 7032 7 3 2 64424 73683
0 7033 7 1 2 59811 83833
0 7034 5 1 1 7033
0 7035 7 1 2 7031 7034
0 7036 5 1 1 7035
0 7037 7 1 2 78174 7036
0 7038 5 1 1 7037
0 7039 7 1 2 7023 7038
0 7040 7 1 2 6996 7039
0 7041 5 1 1 7040
0 7042 7 1 2 83619 7041
0 7043 5 1 1 7042
0 7044 7 17 2 63643 75471
0 7045 5 1 1 83836
0 7046 7 1 2 59812 76236
0 7047 5 2 1 7046
0 7048 7 1 2 77415 83853
0 7049 5 1 1 7048
0 7050 7 2 2 64668 76907
0 7051 5 1 1 83855
0 7052 7 1 2 67497 7051
0 7053 5 1 1 7052
0 7054 7 1 2 82331 7053
0 7055 5 1 1 7054
0 7056 7 1 2 62860 7055
0 7057 5 1 1 7056
0 7058 7 1 2 7049 7057
0 7059 5 1 1 7058
0 7060 7 1 2 83837 7059
0 7061 5 1 1 7060
0 7062 7 1 2 7043 7061
0 7063 5 1 1 7062
0 7064 7 1 2 61225 7063
0 7065 5 1 1 7064
0 7066 7 2 2 67498 78423
0 7067 5 2 1 83857
0 7068 7 1 2 83790 83838
0 7069 7 1 2 83858 7068
0 7070 5 1 1 7069
0 7071 7 1 2 7065 7070
0 7072 5 1 1 7071
0 7073 7 1 2 60079 7072
0 7074 5 1 1 7073
0 7075 7 1 2 83780 78424
0 7076 5 1 1 7075
0 7077 7 3 2 67851 82673
0 7078 7 1 2 62228 83861
0 7079 5 1 1 7078
0 7080 7 1 2 7076 7079
0 7081 5 1 1 7080
0 7082 7 1 2 62507 7081
0 7083 5 1 1 7082
0 7084 7 8 2 64669 62861
0 7085 5 9 1 83864
0 7086 7 1 2 81852 83865
0 7087 5 1 1 7086
0 7088 7 1 2 7083 7087
0 7089 5 1 1 7088
0 7090 7 1 2 83620 7089
0 7091 5 1 1 7090
0 7092 7 4 2 62508 73201
0 7093 5 8 1 83881
0 7094 7 1 2 83770 83882
0 7095 5 1 1 7094
0 7096 7 22 2 61428 62862
0 7097 5 8 1 83893
0 7098 7 1 2 83894 83356
0 7099 7 1 2 7095 7098
0 7100 5 1 1 7099
0 7101 7 1 2 7091 7100
0 7102 5 1 1 7101
0 7103 7 1 2 61226 7102
0 7104 5 1 1 7103
0 7105 7 3 2 83357 75723
0 7106 7 1 2 78210 83923
0 7107 7 1 2 71483 7106
0 7108 5 1 1 7107
0 7109 7 1 2 7104 7108
0 7110 5 1 1 7109
0 7111 7 1 2 60080 7110
0 7112 5 1 1 7111
0 7113 7 2 2 61227 82860
0 7114 5 3 1 83926
0 7115 7 2 2 82954 83030
0 7116 7 1 2 60786 83931
0 7117 5 1 1 7116
0 7118 7 1 2 83928 7117
0 7119 5 1 1 7118
0 7120 7 1 2 59292 7119
0 7121 5 1 1 7120
0 7122 7 1 2 70274 77367
0 7123 5 1 1 7122
0 7124 7 1 2 7121 7123
0 7125 5 1 1 7124
0 7126 7 9 2 59813 63644
0 7127 7 3 2 71664 82599
0 7128 5 1 1 83942
0 7129 7 1 2 83933 83943
0 7130 7 1 2 7125 7129
0 7131 5 1 1 7130
0 7132 7 1 2 7112 7131
0 7133 5 1 1 7132
0 7134 7 1 2 72079 7133
0 7135 5 1 1 7134
0 7136 7 1 2 74305 77392
0 7137 5 1 1 7136
0 7138 7 1 2 83929 7137
0 7139 5 1 1 7138
0 7140 7 1 2 69895 7139
0 7141 5 1 1 7140
0 7142 7 1 2 66169 78959
0 7143 5 1 1 7142
0 7144 7 1 2 77384 7143
0 7145 5 6 1 7144
0 7146 7 1 2 69505 83945
0 7147 5 1 1 7146
0 7148 7 1 2 67240 83932
0 7149 5 1 1 7148
0 7150 7 1 2 7147 7149
0 7151 7 1 2 7141 7150
0 7152 5 1 1 7151
0 7153 7 1 2 78218 83924
0 7154 7 1 2 7152 7153
0 7155 5 1 1 7154
0 7156 7 4 2 68594 70022
0 7157 7 1 2 62863 83452
0 7158 5 1 1 7157
0 7159 7 2 2 65690 76355
0 7160 5 1 1 83955
0 7161 7 1 2 64222 83956
0 7162 5 2 1 7161
0 7163 7 1 2 59814 83957
0 7164 5 1 1 7163
0 7165 7 1 2 59470 82683
0 7166 5 1 1 7165
0 7167 7 1 2 62229 80434
0 7168 7 1 2 7166 7167
0 7169 7 1 2 7164 7168
0 7170 5 1 1 7169
0 7171 7 1 2 3418 76695
0 7172 5 1 1 7171
0 7173 7 1 2 67852 7172
0 7174 7 1 2 7170 7173
0 7175 5 1 1 7174
0 7176 7 1 2 62509 7175
0 7177 7 1 2 7158 7176
0 7178 5 1 1 7177
0 7179 7 1 2 73432 79183
0 7180 5 1 1 7179
0 7181 7 1 2 79959 7180
0 7182 5 1 1 7181
0 7183 7 1 2 59293 7182
0 7184 5 1 1 7183
0 7185 7 1 2 75035 73272
0 7186 5 1 1 7185
0 7187 7 1 2 7184 7186
0 7188 5 1 1 7187
0 7189 7 1 2 62230 7188
0 7190 5 1 1 7189
0 7191 7 2 2 62231 76356
0 7192 5 2 1 83959
0 7193 7 3 2 59471 64670
0 7194 7 1 2 72775 83963
0 7195 7 1 2 83961 7194
0 7196 5 1 1 7195
0 7197 7 1 2 7190 7196
0 7198 5 1 1 7197
0 7199 7 1 2 78175 7198
0 7200 5 1 1 7199
0 7201 7 1 2 62028 7000
0 7202 5 1 1 7201
0 7203 7 1 2 76571 83824
0 7204 7 1 2 7202 7203
0 7205 5 1 1 7204
0 7206 7 1 2 7200 7205
0 7207 7 1 2 7178 7206
0 7208 5 1 1 7207
0 7209 7 1 2 83951 7208
0 7210 5 1 1 7209
0 7211 7 2 2 82458 83659
0 7212 7 1 2 82262 83966
0 7213 7 1 2 83320 7212
0 7214 5 1 1 7213
0 7215 7 1 2 7210 7214
0 7216 5 1 1 7215
0 7217 7 1 2 79507 7216
0 7218 5 1 1 7217
0 7219 7 1 2 7155 7218
0 7220 7 1 2 7135 7219
0 7221 7 1 2 7074 7220
0 7222 5 1 1 7221
0 7223 7 1 2 63323 7222
0 7224 5 1 1 7223
0 7225 7 2 2 71484 78365
0 7226 7 1 2 70023 83968
0 7227 5 1 1 7226
0 7228 7 1 2 62864 80326
0 7229 5 1 1 7228
0 7230 7 1 2 7227 7229
0 7231 5 1 1 7230
0 7232 7 1 2 59815 7231
0 7233 5 1 1 7232
0 7234 7 1 2 62865 75744
0 7235 5 1 1 7234
0 7236 7 1 2 7233 7235
0 7237 5 1 1 7236
0 7238 7 1 2 60880 7237
0 7239 5 1 1 7238
0 7240 7 1 2 74315 83007
0 7241 5 1 1 7240
0 7242 7 1 2 7239 7241
0 7243 5 1 1 7242
0 7244 7 1 2 59472 7243
0 7245 5 1 1 7244
0 7246 7 1 2 75936 5391
0 7247 5 1 1 7246
0 7248 7 1 2 62029 75929
0 7249 7 1 2 77363 7248
0 7250 5 1 1 7249
0 7251 7 1 2 82667 7250
0 7252 7 1 2 7247 7251
0 7253 5 1 1 7252
0 7254 7 1 2 83008 7253
0 7255 5 1 1 7254
0 7256 7 1 2 7245 7255
0 7257 5 1 1 7256
0 7258 7 1 2 79508 7257
0 7259 5 1 1 7258
0 7260 7 2 2 69896 76491
0 7261 5 1 1 83970
0 7262 7 1 2 64887 7261
0 7263 5 2 1 7262
0 7264 7 1 2 83972 78022
0 7265 5 1 1 7264
0 7266 7 1 2 67015 7265
0 7267 5 1 1 7266
0 7268 7 1 2 80482 81966
0 7269 5 1 1 7268
0 7270 7 1 2 7267 7269
0 7271 5 1 1 7270
0 7272 7 1 2 67241 7271
0 7273 5 1 1 7272
0 7274 7 1 2 62232 81612
0 7275 5 1 1 7274
0 7276 7 1 2 62030 72080
0 7277 7 1 2 75982 7276
0 7278 5 1 1 7277
0 7279 7 1 2 7278 82668
0 7280 7 1 2 7275 7279
0 7281 5 1 1 7280
0 7282 7 1 2 64888 7281
0 7283 5 1 1 7282
0 7284 7 1 2 7273 7283
0 7285 5 1 1 7284
0 7286 7 1 2 62866 83614
0 7287 7 1 2 7285 7286
0 7288 5 1 1 7287
0 7289 7 2 2 74199 74333
0 7290 5 1 1 83974
0 7291 7 1 2 72748 83975
0 7292 7 1 2 83969 7291
0 7293 5 1 1 7292
0 7294 7 1 2 7288 7293
0 7295 7 1 2 7259 7294
0 7296 5 1 1 7295
0 7297 7 1 2 63645 7296
0 7298 5 1 1 7297
0 7299 7 7 2 68595 79477
0 7300 5 1 1 83976
0 7301 7 2 2 79467 83977
0 7302 7 2 2 76336 80123
0 7303 5 1 1 83985
0 7304 7 2 2 62031 72179
0 7305 5 1 1 83987
0 7306 7 1 2 60787 83988
0 7307 5 1 1 7306
0 7308 7 1 2 7303 7307
0 7309 5 2 1 7308
0 7310 7 1 2 64671 83989
0 7311 5 1 1 7310
0 7312 7 2 2 59816 69398
0 7313 7 1 2 69054 75036
0 7314 7 1 2 83991 7313
0 7315 5 1 1 7314
0 7316 7 1 2 7311 7315
0 7317 5 1 1 7316
0 7318 7 1 2 59294 7317
0 7319 5 1 1 7318
0 7320 7 4 2 67016 76992
0 7321 5 1 1 83993
0 7322 7 3 2 64425 60788
0 7323 7 1 2 81563 83997
0 7324 7 1 2 83994 7323
0 7325 5 1 1 7324
0 7326 7 1 2 7319 7325
0 7327 5 1 1 7326
0 7328 7 1 2 83983 7327
0 7329 5 1 1 7328
0 7330 7 1 2 67499 7329
0 7331 7 1 2 7298 7330
0 7332 5 1 1 7331
0 7333 7 4 2 63646 72542
0 7334 7 1 2 70131 79306
0 7335 5 2 1 7334
0 7336 7 3 2 83475 84004
0 7337 7 1 2 84000 84006
0 7338 5 1 1 7337
0 7339 7 4 2 60881 62032
0 7340 5 1 1 84009
0 7341 7 1 2 73090 84010
0 7342 5 1 1 7341
0 7343 7 5 2 64426 71302
0 7344 5 4 1 84013
0 7345 7 1 2 81416 84014
0 7346 5 1 1 7345
0 7347 7 1 2 84018 74811
0 7348 5 1 1 7347
0 7349 7 1 2 7348 75762
0 7350 7 1 2 7346 7349
0 7351 5 1 1 7350
0 7352 7 1 2 65793 7351
0 7353 5 1 1 7352
0 7354 7 1 2 7342 7353
0 7355 5 1 1 7354
0 7356 7 1 2 75168 83952
0 7357 7 1 2 7355 7356
0 7358 5 1 1 7357
0 7359 7 1 2 7338 7358
0 7360 5 1 1 7359
0 7361 7 1 2 67853 7360
0 7362 5 1 1 7361
0 7363 7 2 2 75472 75738
0 7364 7 1 2 84022 79367
0 7365 7 1 2 74463 7364
0 7366 5 1 1 7365
0 7367 7 1 2 7362 7366
0 7368 5 1 1 7367
0 7369 7 1 2 64672 7368
0 7370 5 1 1 7369
0 7371 7 1 2 62867 6419
0 7372 5 1 1 7371
0 7373 7 5 2 64427 67854
0 7374 7 1 2 77362 84024
0 7375 5 1 1 7374
0 7376 7 1 2 7372 7375
0 7377 5 1 1 7376
0 7378 7 1 2 63647 84007
0 7379 7 1 2 7377 7378
0 7380 5 1 1 7379
0 7381 7 1 2 59295 83990
0 7382 5 1 1 7381
0 7383 7 1 2 81599 83998
0 7384 5 1 1 7383
0 7385 7 1 2 7382 7384
0 7386 5 1 1 7385
0 7387 7 1 2 59817 83984
0 7388 7 1 2 7386 7387
0 7389 5 1 1 7388
0 7390 7 1 2 62510 7389
0 7391 7 1 2 7380 7390
0 7392 7 1 2 7370 7391
0 7393 5 1 1 7392
0 7394 7 1 2 68248 7393
0 7395 7 1 2 7332 7394
0 7396 5 1 1 7395
0 7397 7 1 2 66629 7396
0 7398 7 1 2 7224 7397
0 7399 5 1 1 7398
0 7400 7 4 2 67500 75169
0 7401 7 2 2 802 74831
0 7402 5 1 1 84033
0 7403 7 1 2 74200 7402
0 7404 5 1 1 7403
0 7405 7 4 2 76549 74181
0 7406 5 1 1 84035
0 7407 7 1 2 78839 84036
0 7408 5 1 1 7407
0 7409 7 1 2 7404 7408
0 7410 5 1 1 7409
0 7411 7 1 2 84029 7410
0 7412 5 1 1 7411
0 7413 7 1 2 62233 77212
0 7414 5 2 1 7413
0 7415 7 1 2 59818 84039
0 7416 5 1 1 7415
0 7417 7 2 2 62511 79318
0 7418 7 1 2 64889 84041
0 7419 7 1 2 7416 7418
0 7420 5 1 1 7419
0 7421 7 1 2 7412 7420
0 7422 5 1 1 7421
0 7423 7 1 2 66170 7422
0 7424 5 1 1 7423
0 7425 7 1 2 72754 74924
0 7426 7 1 2 83854 7425
0 7427 5 1 1 7426
0 7428 7 1 2 7424 7427
0 7429 5 1 1 7428
0 7430 7 1 2 63324 7429
0 7431 5 1 1 7430
0 7432 7 3 2 71019 74925
0 7433 7 1 2 83240 84043
0 7434 5 1 1 7433
0 7435 7 1 2 7431 7434
0 7436 5 1 1 7435
0 7437 7 1 2 67855 7436
0 7438 5 1 1 7437
0 7439 7 3 2 59819 62234
0 7440 5 1 1 84046
0 7441 7 2 2 69630 73091
0 7442 5 4 1 84049
0 7443 7 1 2 76508 84051
0 7444 5 1 1 7443
0 7445 7 1 2 74090 7444
0 7446 5 1 1 7445
0 7447 7 1 2 79150 7446
0 7448 5 1 1 7447
0 7449 7 1 2 7440 7448
0 7450 5 1 1 7449
0 7451 7 1 2 80003 69096
0 7452 5 1 1 7451
0 7453 7 1 2 76993 76252
0 7454 5 1 1 7453
0 7455 7 1 2 62512 7454
0 7456 7 1 2 7452 7455
0 7457 5 2 1 7456
0 7458 7 1 2 76195 84055
0 7459 7 1 2 7450 7458
0 7460 5 1 1 7459
0 7461 7 1 2 69172 74148
0 7462 5 2 1 7461
0 7463 7 2 2 62513 72584
0 7464 5 1 1 84059
0 7465 7 1 2 76994 7464
0 7466 5 1 1 7465
0 7467 7 2 2 69097 78629
0 7468 5 1 1 84061
0 7469 7 1 2 74892 84062
0 7470 5 1 1 7469
0 7471 7 1 2 7466 7470
0 7472 5 1 1 7471
0 7473 7 1 2 74117 7472
0 7474 5 1 1 7473
0 7475 7 1 2 84057 7474
0 7476 7 1 2 7460 7475
0 7477 5 1 1 7476
0 7478 7 1 2 70024 7477
0 7479 5 1 1 7478
0 7480 7 1 2 81668 74709
0 7481 5 1 1 7480
0 7482 7 1 2 73003 82541
0 7483 5 1 1 7482
0 7484 7 1 2 7481 7483
0 7485 5 1 1 7484
0 7486 7 1 2 69776 7485
0 7487 5 1 1 7486
0 7488 7 1 2 68249 7487
0 7489 7 1 2 7479 7488
0 7490 5 1 1 7489
0 7491 7 2 2 60882 70132
0 7492 7 1 2 84063 76938
0 7493 5 1 1 7492
0 7494 7 2 2 69098 83341
0 7495 7 1 2 82877 84065
0 7496 5 1 1 7495
0 7497 7 3 2 76163 74450
0 7498 5 1 1 84067
0 7499 7 1 2 69777 84068
0 7500 5 1 1 7499
0 7501 7 1 2 70587 7500
0 7502 5 1 1 7501
0 7503 7 1 2 7496 7502
0 7504 7 1 2 7493 7503
0 7505 5 1 1 7504
0 7506 7 1 2 59820 7505
0 7507 5 1 1 7506
0 7508 7 1 2 62514 73063
0 7509 5 1 1 7508
0 7510 7 1 2 73445 7509
0 7511 5 1 1 7510
0 7512 7 1 2 64428 7511
0 7513 5 1 1 7512
0 7514 7 5 2 62515 69977
0 7515 5 1 1 84070
0 7516 7 12 2 62235 69778
0 7517 5 4 1 84075
0 7518 7 2 2 60883 84087
0 7519 5 1 1 84091
0 7520 7 1 2 84071 7519
0 7521 5 1 1 7520
0 7522 7 1 2 7513 7521
0 7523 5 1 1 7522
0 7524 7 3 2 62033 69227
0 7525 5 5 1 84093
0 7526 7 5 2 69296 84096
0 7527 7 2 2 60789 84101
0 7528 5 1 1 84106
0 7529 7 1 2 78473 75044
0 7530 5 2 1 7529
0 7531 7 1 2 78306 84108
0 7532 7 1 2 7528 7531
0 7533 7 1 2 7523 7532
0 7534 5 1 1 7533
0 7535 7 1 2 70588 7534
0 7536 5 1 1 7535
0 7537 7 1 2 63325 7536
0 7538 7 1 2 7507 7537
0 7539 5 1 1 7538
0 7540 7 1 2 65104 7539
0 7541 7 1 2 7490 7540
0 7542 5 1 1 7541
0 7543 7 1 2 79307 7542
0 7544 5 1 1 7543
0 7545 7 5 2 62516 70474
0 7546 7 1 2 79953 73583
0 7547 5 1 1 7546
0 7548 7 1 2 84110 7547
0 7549 5 1 1 7548
0 7550 7 2 2 74005 74118
0 7551 5 1 1 84115
0 7552 7 1 2 6463 84116
0 7553 5 1 1 7552
0 7554 7 1 2 59296 7553
0 7555 5 1 1 7554
0 7556 7 3 2 59821 70513
0 7557 5 6 1 84117
0 7558 7 1 2 62517 84120
0 7559 5 1 1 7558
0 7560 7 1 2 7559 82207
0 7561 5 1 1 7560
0 7562 7 1 2 82072 84109
0 7563 7 1 2 7561 7562
0 7564 7 1 2 7555 7563
0 7565 5 1 1 7564
0 7566 7 1 2 64890 7565
0 7567 5 1 1 7566
0 7568 7 1 2 7549 7567
0 7569 5 1 1 7568
0 7570 7 1 2 66171 7569
0 7571 5 1 1 7570
0 7572 7 1 2 66172 71350
0 7573 5 2 1 7572
0 7574 7 1 2 81665 84126
0 7575 5 1 1 7574
0 7576 7 1 2 78608 7575
0 7577 5 1 1 7576
0 7578 7 2 2 77666 78617
0 7579 7 1 2 76164 84128
0 7580 5 1 1 7579
0 7581 7 1 2 7577 7580
0 7582 5 1 1 7581
0 7583 7 1 2 64673 7582
0 7584 5 1 1 7583
0 7585 7 1 2 75250 7584
0 7586 7 1 2 7571 7585
0 7587 5 1 1 7586
0 7588 7 1 2 62868 75404
0 7589 7 1 2 7587 7588
0 7590 7 1 2 7544 7589
0 7591 5 1 1 7590
0 7592 7 1 2 7438 7591
0 7593 5 1 1 7592
0 7594 7 2 2 63648 7593
0 7595 5 1 1 84130
0 7596 7 1 2 61640 7595
0 7597 5 1 1 7596
0 7598 7 1 2 65328 7597
0 7599 7 1 2 7399 7598
0 7600 5 1 1 7599
0 7601 7 1 2 80350 84131
0 7602 5 1 1 7601
0 7603 7 1 2 69055 77416
0 7604 5 2 1 7603
0 7605 7 1 2 78213 84132
0 7606 5 1 1 7605
0 7607 7 12 2 63649 80390
0 7608 7 1 2 79190 84134
0 7609 5 1 1 7608
0 7610 7 3 2 59822 65329
0 7611 7 7 2 62034 68596
0 7612 7 6 2 64891 66630
0 7613 7 1 2 84149 84156
0 7614 7 1 2 84146 7613
0 7615 5 1 1 7614
0 7616 7 1 2 7609 7615
0 7617 5 1 1 7616
0 7618 7 1 2 80151 7617
0 7619 5 1 1 7618
0 7620 7 2 2 81267 83443
0 7621 7 9 2 59823 66631
0 7622 7 1 2 75824 84164
0 7623 7 1 2 74780 7622
0 7624 7 1 2 84162 7623
0 7625 5 1 1 7624
0 7626 7 1 2 7619 7625
0 7627 5 1 1 7626
0 7628 7 1 2 66173 7627
0 7629 5 1 1 7628
0 7630 7 39 2 65330 68597
0 7631 5 1 1 84173
0 7632 7 8 2 63326 84174
0 7633 7 1 2 75170 81280
0 7634 7 1 2 84212 7633
0 7635 7 1 2 82587 7634
0 7636 5 1 1 7635
0 7637 7 1 2 7629 7636
0 7638 5 1 1 7637
0 7639 7 1 2 64429 7638
0 7640 5 1 1 7639
0 7641 7 6 2 75171 80391
0 7642 5 2 1 84220
0 7643 7 7 2 80161 81385
0 7644 5 4 1 84228
0 7645 7 2 2 84226 84235
0 7646 5 5 1 84239
0 7647 7 2 2 63650 84241
0 7648 7 1 2 80665 84246
0 7649 5 1 1 7648
0 7650 7 1 2 7640 7649
0 7651 5 1 1 7650
0 7652 7 1 2 7606 7651
0 7653 5 1 1 7652
0 7654 7 1 2 68829 7653
0 7655 7 1 2 7602 7654
0 7656 7 1 2 7600 7655
0 7657 5 1 1 7656
0 7658 7 1 2 61001 7657
0 7659 7 1 2 6962 7658
0 7660 5 1 1 7659
0 7661 7 1 2 66790 7660
0 7662 7 1 2 5955 7661
0 7663 7 1 2 4907 7662
0 7664 5 1 1 7663
0 7665 7 1 2 65537 7664
0 7666 7 1 2 3186 7665
0 7667 5 1 1 7666
0 7668 7 8 2 65963 61641
0 7669 7 6 2 63651 84248
0 7670 5 1 1 84256
0 7671 7 11 2 61002 66632
0 7672 7 3 2 68598 84262
0 7673 5 1 1 84273
0 7674 7 1 2 64892 84274
0 7675 5 1 1 7674
0 7676 7 1 2 7670 7675
0 7677 5 1 1 7676
0 7678 7 1 2 82448 7677
0 7679 5 1 1 7678
0 7680 7 6 2 62518 69056
0 7681 5 1 1 84276
0 7682 7 8 2 61003 61642
0 7683 7 6 2 63652 84282
0 7684 5 1 1 84290
0 7685 7 1 2 84277 84291
0 7686 5 1 1 7685
0 7687 7 3 2 65964 66633
0 7688 7 2 2 64893 84296
0 7689 7 8 2 67501 68599
0 7690 5 1 1 84301
0 7691 7 2 2 67242 84302
0 7692 7 1 2 84299 84309
0 7693 5 1 1 7692
0 7694 7 1 2 7686 7693
0 7695 7 1 2 7679 7694
0 7696 5 1 1 7695
0 7697 7 1 2 77882 7696
0 7698 5 1 1 7697
0 7699 7 2 2 67502 79031
0 7700 7 1 2 61643 71613
0 7701 7 1 2 84311 7700
0 7702 5 1 1 7701
0 7703 7 3 2 68600 84157
0 7704 5 1 1 84313
0 7705 7 1 2 80196 84278
0 7706 7 1 2 84314 7705
0 7707 5 1 1 7706
0 7708 7 1 2 7702 7707
0 7709 5 1 1 7708
0 7710 7 1 2 62869 7709
0 7711 5 1 1 7710
0 7712 7 1 2 7698 7711
0 7713 5 1 1 7712
0 7714 7 1 2 65331 7713
0 7715 5 1 1 7714
0 7716 7 2 2 65965 74399
0 7717 5 1 1 84316
0 7718 7 1 2 69057 76115
0 7719 5 1 1 7718
0 7720 7 1 2 7717 7719
0 7721 5 1 1 7720
0 7722 7 1 2 67856 7721
0 7723 5 1 1 7722
0 7724 7 3 2 71614 78176
0 7725 5 1 1 84318
0 7726 7 1 2 7723 7725
0 7727 5 1 1 7726
0 7728 7 1 2 80351 79032
0 7729 7 1 2 7727 7728
0 7730 5 1 1 7729
0 7731 7 1 2 7715 7730
0 7732 5 1 1 7731
0 7733 7 1 2 64430 7732
0 7734 5 1 1 7733
0 7735 7 2 2 84135 78268
0 7736 5 1 1 84321
0 7737 7 1 2 76112 78936
0 7738 7 1 2 84322 7737
0 7739 5 1 1 7738
0 7740 7 48 2 66634 68601
0 7741 5 2 1 84323
0 7742 7 16 2 65332 67857
0 7743 5 4 1 84373
0 7744 7 3 2 84324 84374
0 7745 5 1 1 84393
0 7746 7 1 2 64894 76104
0 7747 7 1 2 84394 7746
0 7748 5 1 1 7747
0 7749 7 1 2 7739 7748
0 7750 5 1 1 7749
0 7751 7 1 2 65794 80108
0 7752 7 1 2 7750 7751
0 7753 5 1 1 7752
0 7754 7 1 2 7734 7753
0 7755 5 1 1 7754
0 7756 7 1 2 62035 7755
0 7757 5 1 1 7756
0 7758 7 3 2 62870 69228
0 7759 5 2 1 84396
0 7760 7 4 2 74492 84397
0 7761 5 2 1 84401
0 7762 7 1 2 81521 84402
0 7763 5 1 1 7762
0 7764 7 1 2 82350 7763
0 7765 5 1 1 7764
0 7766 7 1 2 77852 84136
0 7767 7 1 2 7765 7766
0 7768 5 1 1 7767
0 7769 7 1 2 7757 7768
0 7770 5 1 1 7769
0 7771 7 1 2 64674 7770
0 7772 5 1 1 7771
0 7773 7 6 2 64895 63327
0 7774 7 2 2 67503 79002
0 7775 7 4 2 65333 84263
0 7776 7 1 2 83986 84415
0 7777 7 1 2 84413 7776
0 7778 5 1 1 7777
0 7779 7 1 2 77304 69287
0 7780 5 1 1 7779
0 7781 7 1 2 82451 7780
0 7782 5 1 1 7781
0 7783 7 1 2 78960 84137
0 7784 7 1 2 7782 7783
0 7785 5 1 1 7784
0 7786 7 1 2 7778 7785
0 7787 5 1 1 7786
0 7788 7 1 2 84407 7787
0 7789 5 1 1 7788
0 7790 7 1 2 7772 7789
0 7791 5 1 1 7790
0 7792 7 1 2 79509 7791
0 7793 5 1 1 7792
0 7794 7 2 2 80352 76165
0 7795 5 1 1 84419
0 7796 7 33 2 67858 63653
0 7797 7 1 2 71594 84421
0 7798 7 2 2 74167 7797
0 7799 7 1 2 84420 84454
0 7800 5 1 1 7799
0 7801 7 4 2 71165 72288
0 7802 7 3 2 73092 77417
0 7803 5 2 1 84460
0 7804 7 1 2 84456 84461
0 7805 5 1 1 7804
0 7806 7 1 2 83964 84319
0 7807 5 1 1 7806
0 7808 7 1 2 7805 7807
0 7809 5 1 1 7808
0 7810 7 1 2 84325 7809
0 7811 5 1 1 7810
0 7812 7 78 2 61644 63654
0 7813 5 25 1 84465
0 7814 7 1 2 78961 84466
0 7815 7 1 2 84317 7814
0 7816 5 1 1 7815
0 7817 7 1 2 7811 7816
0 7818 5 1 1 7817
0 7819 7 1 2 60884 7818
0 7820 5 1 1 7819
0 7821 7 2 2 61645 76166
0 7822 5 2 1 84568
0 7823 7 1 2 84422 84569
0 7824 7 1 2 82565 7823
0 7825 5 1 1 7824
0 7826 7 1 2 83787 77444
0 7827 5 3 1 7826
0 7828 7 2 2 59473 84326
0 7829 5 1 1 84575
0 7830 7 1 2 69058 74157
0 7831 7 1 2 84576 7830
0 7832 7 1 2 84572 7831
0 7833 5 1 1 7832
0 7834 7 1 2 7825 7833
0 7835 5 1 1 7834
0 7836 7 1 2 61004 7835
0 7837 5 1 1 7836
0 7838 7 4 2 65795 73781
0 7839 5 3 1 84577
0 7840 7 10 2 62236 68602
0 7841 7 16 2 59824 67859
0 7842 5 3 1 84594
0 7843 7 4 2 59474 66635
0 7844 7 1 2 84595 84613
0 7845 7 1 2 84584 7844
0 7846 7 1 2 84578 7845
0 7847 5 1 1 7846
0 7848 7 1 2 7837 7847
0 7849 7 1 2 7820 7848
0 7850 5 1 1 7849
0 7851 7 1 2 65334 7850
0 7852 5 1 1 7851
0 7853 7 1 2 7800 7852
0 7854 5 1 1 7853
0 7855 7 1 2 75172 7854
0 7856 5 1 1 7855
0 7857 7 1 2 83862 84247
0 7858 5 1 1 7857
0 7859 7 5 2 59475 66392
0 7860 7 2 2 84165 84617
0 7861 7 2 2 67243 79003
0 7862 7 1 2 81341 84624
0 7863 7 1 2 84622 7862
0 7864 5 1 1 7863
0 7865 7 1 2 7858 7864
0 7866 5 1 1 7865
0 7867 7 1 2 76116 7866
0 7868 5 1 1 7867
0 7869 7 5 2 66636 76167
0 7870 7 1 2 82697 84626
0 7871 7 1 2 84455 7870
0 7872 5 1 1 7871
0 7873 7 1 2 7868 7872
0 7874 7 1 2 7856 7873
0 7875 5 1 1 7874
0 7876 7 1 2 68250 7875
0 7877 5 1 1 7876
0 7878 7 8 2 65335 65796
0 7879 7 1 2 84585 84631
0 7880 7 1 2 80178 7879
0 7881 5 1 1 7880
0 7882 7 5 2 66393 84586
0 7883 7 6 2 65105 65797
0 7884 5 2 1 84644
0 7885 7 1 2 80392 84645
0 7886 7 1 2 84639 7885
0 7887 5 1 1 7886
0 7888 7 1 2 7881 7887
0 7889 5 1 1 7888
0 7890 7 1 2 64431 7889
0 7891 5 1 1 7890
0 7892 7 1 2 63655 75803
0 7893 7 1 2 80576 7892
0 7894 5 1 1 7893
0 7895 7 1 2 7891 7894
0 7896 5 1 1 7895
0 7897 7 7 2 64675 78928
0 7898 5 6 1 84652
0 7899 7 1 2 75677 84653
0 7900 7 1 2 7896 7899
0 7901 5 1 1 7900
0 7902 7 1 2 7877 7901
0 7903 5 1 1 7902
0 7904 7 1 2 64896 7903
0 7905 5 1 1 7904
0 7906 7 1 2 66174 7905
0 7907 7 1 2 7793 7906
0 7908 5 1 1 7907
0 7909 7 4 2 64676 63656
0 7910 7 2 2 81967 78863
0 7911 7 1 2 80152 84669
0 7912 5 1 1 7911
0 7913 7 4 2 65966 67017
0 7914 5 1 1 84671
0 7915 7 1 2 82973 84672
0 7916 7 1 2 83166 7915
0 7917 5 1 1 7916
0 7918 7 1 2 7912 7917
0 7919 5 1 1 7918
0 7920 7 1 2 62519 7919
0 7921 5 1 1 7920
0 7922 7 3 2 71351 77883
0 7923 7 1 2 75173 82642
0 7924 7 1 2 84675 7923
0 7925 5 1 1 7924
0 7926 7 1 2 7921 7925
0 7927 5 1 1 7926
0 7928 7 1 2 61646 7927
0 7929 5 1 1 7928
0 7930 7 1 2 77884 71862
0 7931 5 2 1 7930
0 7932 7 2 2 73782 77760
0 7933 5 1 1 84680
0 7934 7 1 2 84678 7933
0 7935 5 1 1 7934
0 7936 7 7 2 66637 67244
0 7937 7 2 2 61429 84682
0 7938 7 1 2 74260 84689
0 7939 7 1 2 7935 7938
0 7940 5 1 1 7939
0 7941 7 1 2 7929 7940
0 7942 5 1 1 7941
0 7943 7 1 2 65798 7942
0 7944 5 1 1 7943
0 7945 7 1 2 73765 82663
0 7946 7 3 2 77269 7945
0 7947 7 4 2 61647 83086
0 7948 5 1 1 84694
0 7949 7 2 2 79319 84695
0 7950 7 1 2 84691 84698
0 7951 5 1 1 7950
0 7952 7 1 2 7944 7951
0 7953 5 1 1 7952
0 7954 7 1 2 64432 7953
0 7955 5 1 1 7954
0 7956 7 1 2 73684 73783
0 7957 5 2 1 7956
0 7958 7 1 2 65799 84692
0 7959 5 1 1 7958
0 7960 7 1 2 84700 7959
0 7961 5 1 1 7960
0 7962 7 1 2 84699 7961
0 7963 5 1 1 7962
0 7964 7 1 2 7955 7963
0 7965 5 1 1 7964
0 7966 7 1 2 84665 7965
0 7967 5 1 1 7966
0 7968 7 2 2 75174 84467
0 7969 5 2 1 84702
0 7970 7 1 2 80722 79062
0 7971 5 1 1 7970
0 7972 7 1 2 67860 80631
0 7973 5 1 1 7972
0 7974 7 1 2 7971 7973
0 7975 5 2 1 7974
0 7976 7 1 2 71747 84706
0 7977 5 1 1 7976
0 7978 7 4 2 61005 62036
0 7979 5 2 1 84708
0 7980 7 4 2 62237 77885
0 7981 5 1 1 84714
0 7982 7 1 2 84709 84715
0 7983 5 1 1 7982
0 7984 7 1 2 7977 7983
0 7985 5 1 1 7984
0 7986 7 1 2 62520 7985
0 7987 5 1 1 7986
0 7988 7 1 2 71952 80444
0 7989 5 2 1 7988
0 7990 7 1 2 71166 84718
0 7991 5 2 1 7990
0 7992 7 1 2 82337 84720
0 7993 5 1 1 7992
0 7994 7 1 2 7987 7993
0 7995 5 1 1 7994
0 7996 7 1 2 84703 7995
0 7997 5 1 1 7996
0 7998 7 1 2 61430 84707
0 7999 5 1 1 7998
0 8000 7 3 2 61006 62238
0 8001 5 2 1 84722
0 8002 7 1 2 75825 78962
0 8003 7 1 2 84723 8002
0 8004 5 1 1 8003
0 8005 7 1 2 7999 8004
0 8006 5 1 1 8005
0 8007 7 1 2 71748 8006
0 8008 5 1 1 8007
0 8009 7 1 2 73561 75826
0 8010 5 1 1 8009
0 8011 7 16 2 62239 63328
0 8012 5 3 1 84727
0 8013 7 3 2 61431 84728
0 8014 5 3 1 84746
0 8015 7 1 2 8010 84749
0 8016 5 1 1 8015
0 8017 7 1 2 61007 8016
0 8018 5 1 1 8017
0 8019 7 2 2 66394 80805
0 8020 5 3 1 84752
0 8021 7 1 2 81579 84753
0 8022 5 1 1 8021
0 8023 7 1 2 8018 8022
0 8024 5 1 1 8023
0 8025 7 1 2 78963 8024
0 8026 5 1 1 8025
0 8027 7 1 2 8008 8026
0 8028 5 1 1 8027
0 8029 7 1 2 62521 8028
0 8030 5 1 1 8029
0 8031 7 2 2 67504 84721
0 8032 5 1 1 84757
0 8033 7 2 2 67861 81214
0 8034 5 1 1 84759
0 8035 7 1 2 66395 79245
0 8036 5 1 1 8035
0 8037 7 1 2 84760 8036
0 8038 7 1 2 84758 8037
0 8039 5 1 1 8038
0 8040 7 1 2 8030 8039
0 8041 5 1 1 8040
0 8042 7 1 2 63657 8041
0 8043 5 1 1 8042
0 8044 7 5 2 66396 71953
0 8045 7 16 2 62522 68603
0 8046 7 2 2 78692 84766
0 8047 7 2 2 84761 84782
0 8048 5 2 1 84784
0 8049 7 3 2 63329 71065
0 8050 7 1 2 84785 84788
0 8051 5 1 1 8050
0 8052 7 1 2 60243 8051
0 8053 7 1 2 8043 8052
0 8054 5 1 1 8053
0 8055 7 4 2 82600 84423
0 8056 5 1 1 84791
0 8057 7 1 2 84786 8056
0 8058 5 1 1 8057
0 8059 7 1 2 71066 8058
0 8060 5 1 1 8059
0 8061 7 18 2 61008 67862
0 8062 5 2 1 84795
0 8063 7 1 2 63658 81044
0 8064 7 1 2 84796 8063
0 8065 7 1 2 81834 8064
0 8066 5 1 1 8065
0 8067 7 1 2 8060 8066
0 8068 5 1 1 8067
0 8069 7 1 2 68251 8068
0 8070 5 1 1 8069
0 8071 7 6 2 68604 77886
0 8072 5 1 1 84815
0 8073 7 1 2 73864 74859
0 8074 7 1 2 82444 8073
0 8075 7 1 2 84816 8074
0 8076 5 1 1 8075
0 8077 7 1 2 8070 8076
0 8078 5 1 1 8077
0 8079 7 1 2 62037 8078
0 8080 5 1 1 8079
0 8081 7 17 2 61432 67863
0 8082 5 5 1 84821
0 8083 7 5 2 63659 84822
0 8084 7 1 2 74215 73784
0 8085 7 1 2 84843 8084
0 8086 5 1 1 8085
0 8087 7 2 2 78177 83515
0 8088 5 2 1 84848
0 8089 7 7 2 64433 66397
0 8090 5 1 1 84852
0 8091 7 1 2 82643 84853
0 8092 7 1 2 84849 8091
0 8093 5 1 1 8092
0 8094 7 1 2 8086 8093
0 8095 5 1 1 8094
0 8096 7 1 2 60885 8095
0 8097 5 1 1 8096
0 8098 7 1 2 64434 76117
0 8099 5 1 1 8098
0 8100 7 2 2 61009 70941
0 8101 5 1 1 84859
0 8102 7 1 2 8099 8101
0 8103 5 1 1 8102
0 8104 7 14 2 68605 80016
0 8105 7 1 2 83863 84861
0 8106 7 1 2 8103 8105
0 8107 5 1 1 8106
0 8108 7 1 2 8097 8107
0 8109 5 1 1 8108
0 8110 7 1 2 67245 8109
0 8111 5 1 1 8110
0 8112 7 2 2 73888 74844
0 8113 7 9 2 62523 83087
0 8114 7 3 2 84587 84877
0 8115 5 1 1 84886
0 8116 7 1 2 84875 84887
0 8117 5 1 1 8116
0 8118 7 1 2 65106 8117
0 8119 7 1 2 8111 8118
0 8120 7 1 2 8080 8119
0 8121 5 1 1 8120
0 8122 7 1 2 66638 8121
0 8123 7 1 2 8054 8122
0 8124 5 1 1 8123
0 8125 7 1 2 7997 8124
0 8126 5 1 1 8125
0 8127 7 1 2 60081 8126
0 8128 5 1 1 8127
0 8129 7 1 2 7967 8128
0 8130 5 1 1 8129
0 8131 7 1 2 65336 8130
0 8132 5 1 1 8131
0 8133 7 3 2 63660 80353
0 8134 7 1 2 77305 76168
0 8135 7 1 2 74049 8134
0 8136 5 1 1 8135
0 8137 7 1 2 8032 8136
0 8138 5 1 1 8137
0 8139 7 1 2 60082 8138
0 8140 5 1 1 8139
0 8141 7 3 2 73004 71863
0 8142 5 1 1 84892
0 8143 7 1 2 74710 84893
0 8144 5 1 1 8143
0 8145 7 1 2 8140 8144
0 8146 5 1 1 8145
0 8147 7 1 2 66398 8146
0 8148 5 1 1 8147
0 8149 7 1 2 76169 81250
0 8150 7 1 2 82046 8149
0 8151 5 1 1 8150
0 8152 7 1 2 8148 8151
0 8153 5 1 1 8152
0 8154 7 1 2 67864 8153
0 8155 5 1 1 8154
0 8156 7 2 2 62871 78943
0 8157 7 1 2 71749 84693
0 8158 5 1 1 8157
0 8159 7 1 2 8158 84701
0 8160 5 2 1 8159
0 8161 7 1 2 84895 84897
0 8162 5 1 1 8161
0 8163 7 1 2 8155 8162
0 8164 5 1 1 8163
0 8165 7 1 2 65107 8164
0 8166 5 1 1 8165
0 8167 7 1 2 62872 84898
0 8168 5 1 1 8167
0 8169 7 10 2 65800 76866
0 8170 5 8 1 84899
0 8171 7 1 2 84900 84670
0 8172 5 1 1 8171
0 8173 7 1 2 8168 8172
0 8174 5 1 1 8173
0 8175 7 1 2 79079 8174
0 8176 5 1 1 8175
0 8177 7 1 2 8166 8176
0 8178 5 1 1 8177
0 8179 7 1 2 63330 8178
0 8180 5 1 1 8179
0 8181 7 1 2 80206 4468
0 8182 5 1 1 8181
0 8183 7 1 2 64435 8182
0 8184 5 1 1 8183
0 8185 7 1 2 60083 69059
0 8186 5 1 1 8185
0 8187 7 1 2 8184 8186
0 8188 5 1 1 8187
0 8189 7 4 2 68252 77454
0 8190 5 1 1 84917
0 8191 7 2 2 75175 71067
0 8192 7 1 2 84918 84921
0 8193 7 1 2 8188 8192
0 8194 5 1 1 8193
0 8195 7 1 2 8180 8194
0 8196 5 1 1 8195
0 8197 7 1 2 84889 8196
0 8198 5 1 1 8197
0 8199 7 1 2 61228 8198
0 8200 7 1 2 8132 8199
0 8201 5 1 1 8200
0 8202 7 1 2 7908 8201
0 8203 5 1 1 8202
0 8204 7 2 2 79320 80393
0 8205 7 3 2 77065 78524
0 8206 7 3 2 67865 79033
0 8207 7 1 2 84925 84928
0 8208 7 1 2 84923 8207
0 8209 7 1 2 82455 8208
0 8210 5 1 1 8209
0 8211 7 1 2 68830 8210
0 8212 7 1 2 8203 8211
0 8213 5 1 1 8212
0 8214 7 1 2 65967 74348
0 8215 5 1 1 8214
0 8216 7 4 2 64897 74360
0 8217 5 3 1 84931
0 8218 7 3 2 61010 73005
0 8219 5 2 1 84938
0 8220 7 1 2 74334 84939
0 8221 5 1 1 8220
0 8222 7 1 2 84935 8221
0 8223 5 1 1 8222
0 8224 7 1 2 62524 8223
0 8225 5 1 1 8224
0 8226 7 1 2 8215 8225
0 8227 7 9 2 61433 70475
0 8228 5 1 1 84943
0 8229 7 3 2 70942 70921
0 8230 5 1 1 84952
0 8231 7 1 2 84944 84953
0 8232 5 1 1 8231
0 8233 7 1 2 74873 8232
0 8234 5 1 1 8233
0 8235 7 1 2 64677 8234
0 8236 5 1 1 8235
0 8237 7 1 2 66399 73927
0 8238 5 2 1 8237
0 8239 7 1 2 82566 74656
0 8240 7 1 2 84955 8239
0 8241 5 1 1 8240
0 8242 7 1 2 8236 8241
0 8243 7 1 2 8226 8242
0 8244 5 1 1 8243
0 8245 7 1 2 65108 8244
0 8246 5 1 1 8245
0 8247 7 4 2 78799 79392
0 8248 5 1 1 84957
0 8249 7 1 2 69151 84958
0 8250 5 1 1 8249
0 8251 7 3 2 64898 79552
0 8252 7 1 2 79574 84961
0 8253 5 1 1 8252
0 8254 7 2 2 76625 79242
0 8255 5 1 1 84964
0 8256 7 1 2 8248 8255
0 8257 5 1 1 8256
0 8258 7 2 2 75251 74657
0 8259 7 1 2 65801 84966
0 8260 7 1 2 8257 8259
0 8261 5 1 1 8260
0 8262 7 1 2 8253 8261
0 8263 5 1 1 8262
0 8264 7 1 2 64436 8263
0 8265 5 1 1 8264
0 8266 7 1 2 8250 8265
0 8267 7 1 2 8246 8266
0 8268 5 1 1 8267
0 8269 7 1 2 63331 8268
0 8270 5 1 1 8269
0 8271 7 1 2 74878 84710
0 8272 5 1 1 8271
0 8273 7 1 2 71954 77018
0 8274 5 1 1 8273
0 8275 7 1 2 8272 8274
0 8276 5 1 1 8275
0 8277 7 1 2 73514 8276
0 8278 5 1 1 8277
0 8279 7 3 2 62038 74400
0 8280 5 1 1 84968
0 8281 7 1 2 64899 84969
0 8282 5 1 1 8281
0 8283 7 1 2 8278 8282
0 8284 5 1 1 8283
0 8285 7 2 2 77598 8284
0 8286 5 1 1 84971
0 8287 7 1 2 75176 84972
0 8288 5 1 1 8287
0 8289 7 2 2 72081 83135
0 8290 5 4 1 84973
0 8291 7 1 2 80153 84975
0 8292 5 1 1 8291
0 8293 7 1 2 76196 75961
0 8294 5 2 1 8293
0 8295 7 4 2 76658 84979
0 8296 7 1 2 83167 84981
0 8297 5 1 1 8296
0 8298 7 1 2 8292 8297
0 8299 5 1 1 8298
0 8300 7 1 2 71068 8299
0 8301 5 1 1 8300
0 8302 7 1 2 80158 70958
0 8303 5 1 1 8302
0 8304 7 1 2 8301 8303
0 8305 5 1 1 8304
0 8306 7 1 2 70737 8305
0 8307 5 1 1 8306
0 8308 7 1 2 8288 8307
0 8309 7 1 2 8270 8308
0 8310 5 1 1 8309
0 8311 7 1 2 67866 8310
0 8312 5 1 1 8311
0 8313 7 5 2 66400 80723
0 8314 5 3 1 84985
0 8315 7 1 2 79801 84990
0 8316 5 2 1 8315
0 8317 7 1 2 76737 76141
0 8318 5 1 1 8317
0 8319 7 1 2 77977 78848
0 8320 5 1 1 8319
0 8321 7 1 2 8318 8320
0 8322 5 2 1 8321
0 8323 7 1 2 84993 84995
0 8324 5 1 1 8323
0 8325 7 1 2 74335 83398
0 8326 5 2 1 8325
0 8327 7 4 2 70025 75060
0 8328 5 4 1 84999
0 8329 7 1 2 81251 85000
0 8330 5 1 1 8329
0 8331 7 1 2 84997 8330
0 8332 5 1 1 8331
0 8333 7 1 2 71069 8332
0 8334 5 1 1 8333
0 8335 7 6 2 63332 70738
0 8336 5 5 1 85007
0 8337 7 2 2 76142 85008
0 8338 5 1 1 85018
0 8339 7 1 2 75872 85019
0 8340 5 2 1 8339
0 8341 7 1 2 8334 85020
0 8342 7 1 2 8324 8341
0 8343 5 1 1 8342
0 8344 7 1 2 71750 8343
0 8345 5 1 1 8344
0 8346 7 2 2 61229 84729
0 8347 5 1 1 85022
0 8348 7 2 2 71955 80621
0 8349 5 1 1 85024
0 8350 7 1 2 8347 8349
0 8351 5 1 1 8350
0 8352 7 1 2 71070 8351
0 8353 5 1 1 8352
0 8354 7 1 2 76154 84730
0 8355 5 1 1 8354
0 8356 7 1 2 8353 8355
0 8357 5 1 1 8356
0 8358 7 1 2 79510 8357
0 8359 5 1 1 8358
0 8360 7 1 2 73562 76155
0 8361 5 1 1 8360
0 8362 7 1 2 74703 73889
0 8363 5 1 1 8362
0 8364 7 1 2 8361 8363
0 8365 5 3 1 8364
0 8366 7 1 2 82513 85026
0 8367 5 1 1 8366
0 8368 7 2 2 71071 81948
0 8369 7 1 2 64900 83612
0 8370 7 1 2 85029 8369
0 8371 5 1 1 8370
0 8372 7 1 2 8367 8371
0 8373 7 1 2 8359 8372
0 8374 7 1 2 8345 8373
0 8375 5 1 1 8374
0 8376 7 1 2 62873 8375
0 8377 5 1 1 8376
0 8378 7 2 2 64901 74565
0 8379 5 1 1 85031
0 8380 7 17 2 66401 62240
0 8381 5 6 1 85033
0 8382 7 2 2 81522 85034
0 8383 7 1 2 72815 85056
0 8384 7 1 2 85032 8383
0 8385 5 1 1 8384
0 8386 7 1 2 8377 8385
0 8387 5 1 1 8386
0 8388 7 1 2 62039 8387
0 8389 5 1 1 8388
0 8390 7 1 2 8312 8389
0 8391 5 1 1 8390
0 8392 7 1 2 80840 8391
0 8393 5 1 1 8392
0 8394 7 6 2 64902 62874
0 8395 5 4 1 85058
0 8396 7 1 2 77356 78937
0 8397 5 1 1 8396
0 8398 7 1 2 64678 8397
0 8399 5 1 1 8398
0 8400 7 1 2 85064 8399
0 8401 5 2 1 8400
0 8402 7 1 2 84945 85068
0 8403 5 1 1 8402
0 8404 7 4 2 66402 78244
0 8405 5 2 1 85070
0 8406 7 1 2 77872 72289
0 8407 7 1 2 84712 8406
0 8408 7 1 2 85071 8407
0 8409 5 1 1 8408
0 8410 7 1 2 8403 8409
0 8411 5 1 1 8410
0 8412 7 1 2 71751 8411
0 8413 5 1 1 8412
0 8414 7 3 2 62241 73563
0 8415 5 2 1 85076
0 8416 7 4 2 67505 82644
0 8417 5 3 1 85081
0 8418 7 1 2 85077 85082
0 8419 5 1 1 8418
0 8420 7 1 2 77306 76197
0 8421 5 2 1 8420
0 8422 7 1 2 60084 76659
0 8423 7 1 2 85088 8422
0 8424 5 1 1 8423
0 8425 7 1 2 8419 8424
0 8426 5 1 1 8425
0 8427 7 1 2 82395 8426
0 8428 5 1 1 8427
0 8429 7 3 2 61434 82363
0 8430 5 3 1 85090
0 8431 7 3 2 71956 71072
0 8432 5 2 1 85096
0 8433 7 1 2 73586 85099
0 8434 5 1 1 8433
0 8435 7 1 2 85091 8434
0 8436 5 1 1 8435
0 8437 7 1 2 8428 8436
0 8438 7 1 2 8413 8437
0 8439 5 1 1 8438
0 8440 7 1 2 61230 8439
0 8441 5 1 1 8440
0 8442 7 3 2 62525 79843
0 8443 5 1 1 85101
0 8444 7 1 2 77681 85102
0 8445 5 1 1 8444
0 8446 7 1 2 70889 84982
0 8447 5 1 1 8446
0 8448 7 1 2 8445 8447
0 8449 5 1 1 8448
0 8450 7 1 2 64679 8449
0 8451 5 1 1 8450
0 8452 7 1 2 70026 84983
0 8453 5 1 1 8452
0 8454 7 1 2 8451 8453
0 8455 5 1 1 8454
0 8456 7 1 2 67867 8455
0 8457 5 1 1 8456
0 8458 7 5 2 62040 78545
0 8459 5 7 1 85104
0 8460 7 1 2 71864 85105
0 8461 7 1 2 81835 8460
0 8462 5 1 1 8461
0 8463 7 1 2 8457 8462
0 8464 5 1 1 8463
0 8465 7 1 2 61435 8464
0 8466 5 1 1 8465
0 8467 7 1 2 8441 8466
0 8468 5 1 1 8467
0 8469 7 1 2 60244 8468
0 8470 5 1 1 8469
0 8471 7 1 2 81880 82645
0 8472 5 1 1 8471
0 8473 7 1 2 73543 8472
0 8474 5 1 1 8473
0 8475 7 3 2 67506 74050
0 8476 5 1 1 85116
0 8477 7 1 2 8474 85117
0 8478 5 1 1 8477
0 8479 7 1 2 80925 76170
0 8480 5 1 1 8479
0 8481 7 1 2 8478 8480
0 8482 5 1 1 8481
0 8483 7 1 2 61436 82847
0 8484 7 1 2 8482 8483
0 8485 5 1 1 8484
0 8486 7 1 2 8470 8485
0 8487 5 1 1 8486
0 8488 7 1 2 68253 8487
0 8489 5 1 1 8488
0 8490 7 2 2 61011 76537
0 8491 7 1 2 75994 73539
0 8492 5 1 1 8491
0 8493 7 1 2 85119 8492
0 8494 5 1 1 8493
0 8495 7 1 2 73544 8494
0 8496 5 1 1 8495
0 8497 7 2 2 74988 8496
0 8498 5 1 1 85121
0 8499 7 2 2 60245 84823
0 8500 5 2 1 85123
0 8501 7 1 2 85122 85124
0 8502 5 1 1 8501
0 8503 7 1 2 8489 8502
0 8504 5 1 1 8503
0 8505 7 1 2 81147 8504
0 8506 5 1 1 8505
0 8507 7 1 2 8393 8506
0 8508 5 1 1 8507
0 8509 7 1 2 68606 8508
0 8510 5 1 1 8509
0 8511 7 18 2 60443 63661
0 8512 5 5 1 85127
0 8513 7 3 2 81986 85128
0 8514 7 3 2 77066 74845
0 8515 5 2 1 85153
0 8516 7 1 2 3083 85156
0 8517 5 3 1 8516
0 8518 7 1 2 72644 85158
0 8519 5 1 1 8518
0 8520 7 3 2 62242 79321
0 8521 5 1 1 85161
0 8522 7 1 2 61012 85162
0 8523 5 1 1 8522
0 8524 7 1 2 8519 8523
0 8525 5 1 1 8524
0 8526 7 1 2 73907 8525
0 8527 5 1 1 8526
0 8528 7 1 2 71957 74229
0 8529 5 1 1 8528
0 8530 7 1 2 77747 8529
0 8531 5 1 1 8530
0 8532 7 1 2 62243 8531
0 8533 5 1 1 8532
0 8534 7 1 2 71752 78500
0 8535 5 1 1 8534
0 8536 7 1 2 8533 8535
0 8537 5 1 1 8536
0 8538 7 1 2 75473 8537
0 8539 5 1 1 8538
0 8540 7 1 2 8527 8539
0 8541 5 1 1 8540
0 8542 7 1 2 67868 8541
0 8543 5 1 1 8542
0 8544 7 1 2 71352 72487
0 8545 5 2 1 8544
0 8546 7 1 2 76125 74497
0 8547 5 1 1 8546
0 8548 7 1 2 85164 8547
0 8549 5 1 1 8548
0 8550 7 1 2 79922 82830
0 8551 7 1 2 8549 8550
0 8552 5 1 1 8551
0 8553 7 1 2 8543 8552
0 8554 5 1 1 8553
0 8555 7 1 2 85150 8554
0 8556 5 1 1 8555
0 8557 7 1 2 63912 8556
0 8558 7 1 2 8510 8557
0 8559 5 1 1 8558
0 8560 7 1 2 8213 8559
0 8561 5 1 1 8560
0 8562 7 1 2 66791 8561
0 8563 5 1 1 8562
0 8564 7 1 2 84327 85027
0 8565 5 1 1 8564
0 8566 7 1 2 61231 84901
0 8567 5 1 1 8566
0 8568 7 1 2 85165 8567
0 8569 5 1 1 8568
0 8570 7 1 2 84468 8569
0 8571 5 1 1 8570
0 8572 7 1 2 8565 8571
0 8573 5 1 1 8572
0 8574 7 1 2 62875 8573
0 8575 5 1 1 8574
0 8576 7 4 2 68607 77685
0 8577 7 2 2 77721 85166
0 8578 7 2 2 67246 77418
0 8579 5 1 1 85172
0 8580 7 3 2 66639 85173
0 8581 7 1 2 85170 85174
0 8582 5 1 1 8581
0 8583 7 1 2 8575 8582
0 8584 5 1 1 8583
0 8585 7 1 2 62041 8584
0 8586 5 1 1 8585
0 8587 7 16 2 62526 63662
0 8588 7 8 2 61648 85177
0 8589 5 2 1 85193
0 8590 7 4 2 64680 68608
0 8591 7 2 2 84297 85203
0 8592 5 1 1 85207
0 8593 7 1 2 85201 8592
0 8594 5 1 1 8593
0 8595 7 2 2 70739 8594
0 8596 5 1 1 85209
0 8597 7 1 2 62527 84543
0 8598 5 1 1 8597
0 8599 7 1 2 85210 8598
0 8600 5 1 1 8599
0 8601 7 1 2 73739 84315
0 8602 5 1 1 8601
0 8603 7 2 2 84249 85178
0 8604 5 1 1 85211
0 8605 7 4 2 64681 85212
0 8606 5 2 1 85213
0 8607 7 1 2 8602 85217
0 8608 7 1 2 8600 8607
0 8609 5 1 1 8608
0 8610 7 1 2 71958 78864
0 8611 7 1 2 8609 8610
0 8612 5 1 1 8611
0 8613 7 1 2 8586 8612
0 8614 5 1 1 8613
0 8615 7 1 2 66403 8614
0 8616 5 1 1 8615
0 8617 7 3 2 66175 78178
0 8618 5 2 1 85219
0 8619 7 1 2 74272 85220
0 8620 5 2 1 8619
0 8621 7 1 2 66176 78865
0 8622 5 3 1 8621
0 8623 7 1 2 85093 85226
0 8624 5 1 1 8623
0 8625 7 1 2 84902 8624
0 8626 5 1 1 8625
0 8627 7 1 2 85224 8626
0 8628 5 2 1 8627
0 8629 7 1 2 77826 84469
0 8630 7 1 2 85229 8629
0 8631 5 1 1 8630
0 8632 7 1 2 8616 8631
0 8633 5 1 1 8632
0 8634 7 1 2 65109 8633
0 8635 5 1 1 8634
0 8636 7 3 2 74273 78179
0 8637 5 2 1 85231
0 8638 7 1 2 65802 84462
0 8639 5 1 1 8638
0 8640 7 1 2 85234 8639
0 8641 5 2 1 8640
0 8642 7 2 2 72686 85236
0 8643 5 1 1 85238
0 8644 7 4 2 64903 62244
0 8645 5 2 1 85240
0 8646 7 4 2 71073 85241
0 8647 5 1 1 85246
0 8648 7 1 2 67869 85247
0 8649 5 1 1 8648
0 8650 7 1 2 8643 8649
0 8651 5 1 1 8650
0 8652 7 1 2 80319 8651
0 8653 5 1 1 8652
0 8654 7 1 2 78036 82378
0 8655 5 3 1 8654
0 8656 7 2 2 78583 85250
0 8657 7 1 2 84903 85253
0 8658 5 1 1 8657
0 8659 7 2 2 85225 8658
0 8660 5 1 1 85255
0 8661 7 1 2 80183 77839
0 8662 5 1 1 8661
0 8663 7 1 2 79273 80184
0 8664 5 4 1 8663
0 8665 7 1 2 8662 85257
0 8666 7 1 2 8660 8665
0 8667 5 1 1 8666
0 8668 7 1 2 8653 8667
0 8669 5 1 1 8668
0 8670 7 1 2 63663 8669
0 8671 5 1 1 8670
0 8672 7 1 2 8635 8671
0 8673 5 1 1 8672
0 8674 7 1 2 65337 8673
0 8675 5 1 1 8674
0 8676 7 2 2 80989 84175
0 8677 7 1 2 77628 85261
0 8678 5 1 1 8677
0 8679 7 1 2 61437 77167
0 8680 5 3 1 8679
0 8681 7 3 2 80394 85179
0 8682 5 1 1 85266
0 8683 7 1 2 79566 85267
0 8684 7 1 2 85263 8683
0 8685 5 1 1 8684
0 8686 7 1 2 8678 8685
0 8687 5 1 1 8686
0 8688 7 1 2 62876 8687
0 8689 5 1 1 8688
0 8690 7 1 2 66177 84813
0 8691 5 1 1 8690
0 8692 7 1 2 70740 74879
0 8693 7 1 2 85262 8692
0 8694 7 1 2 8691 8693
0 8695 5 1 1 8694
0 8696 7 1 2 8689 8695
0 8697 5 1 1 8696
0 8698 7 1 2 65110 8697
0 8699 5 1 1 8698
0 8700 7 6 2 71074 79393
0 8701 5 1 1 85269
0 8702 7 1 2 81148 85270
0 8703 5 1 1 8702
0 8704 7 1 2 84236 8703
0 8705 5 1 1 8704
0 8706 7 1 2 61232 79385
0 8707 7 1 2 8705 8706
0 8708 5 1 1 8707
0 8709 7 1 2 8699 8708
0 8710 5 1 1 8709
0 8711 7 1 2 70476 8710
0 8712 5 1 1 8711
0 8713 7 3 2 74704 77067
0 8714 7 2 2 65338 85275
0 8715 7 1 2 84683 84792
0 8716 7 1 2 85278 8715
0 8717 5 1 1 8716
0 8718 7 1 2 8712 8717
0 8719 5 1 1 8718
0 8720 7 1 2 71753 8719
0 8721 5 1 1 8720
0 8722 7 3 2 77853 79529
0 8723 5 2 1 85280
0 8724 7 1 2 85230 85281
0 8725 5 1 1 8724
0 8726 7 2 2 66404 77179
0 8727 7 1 2 65111 85239
0 8728 5 1 1 8727
0 8729 7 1 2 85256 8728
0 8730 5 1 1 8729
0 8731 7 1 2 85285 8730
0 8732 5 1 1 8731
0 8733 7 1 2 8725 8732
0 8734 5 1 1 8733
0 8735 7 1 2 84890 8734
0 8736 5 1 1 8735
0 8737 7 1 2 8721 8736
0 8738 7 1 2 8675 8737
0 8739 5 1 1 8738
0 8740 7 1 2 68254 8739
0 8741 5 1 1 8740
0 8742 7 3 2 60444 84470
0 8743 5 7 1 85287
0 8744 7 1 2 62877 85288
0 8745 7 1 2 81860 8744
0 8746 5 1 1 8745
0 8747 7 10 2 61233 66640
0 8748 7 3 2 84375 85297
0 8749 7 1 2 71865 85307
0 8750 5 1 1 8749
0 8751 7 3 2 62528 80395
0 8752 7 3 2 71959 70027
0 8753 7 1 2 82629 85313
0 8754 7 1 2 85310 8753
0 8755 5 1 1 8754
0 8756 7 1 2 8750 8755
0 8757 5 1 1 8756
0 8758 7 1 2 64682 8757
0 8759 5 1 1 8758
0 8760 7 1 2 74401 82646
0 8761 5 1 1 8760
0 8762 7 1 2 73545 8761
0 8763 5 1 1 8762
0 8764 7 1 2 85308 8763
0 8765 5 1 1 8764
0 8766 7 1 2 8759 8765
0 8767 5 1 1 8766
0 8768 7 1 2 68609 8767
0 8769 5 1 1 8768
0 8770 7 2 2 81724 85180
0 8771 7 1 2 81958 85316
0 8772 5 1 1 8771
0 8773 7 11 2 65339 84328
0 8774 7 2 2 82916 71866
0 8775 7 1 2 85318 85329
0 8776 5 1 1 8775
0 8777 7 1 2 8772 8776
0 8778 5 1 1 8777
0 8779 7 1 2 82567 8778
0 8780 5 1 1 8779
0 8781 7 1 2 8769 8780
0 8782 7 1 2 8746 8781
0 8783 5 1 1 8782
0 8784 7 1 2 75177 8783
0 8785 5 1 1 8784
0 8786 7 1 2 78180 84138
0 8787 7 1 2 81861 8786
0 8788 5 1 1 8787
0 8789 7 4 2 67870 71754
0 8790 7 1 2 72157 85331
0 8791 7 1 2 84139 8790
0 8792 7 1 2 77844 8791
0 8793 5 1 1 8792
0 8794 7 3 2 66178 81281
0 8795 7 13 2 67871 68610
0 8796 7 5 2 65340 85338
0 8797 5 1 1 85351
0 8798 7 2 2 85335 85352
0 8799 7 3 2 62529 71960
0 8800 5 1 1 85358
0 8801 7 1 2 85248 85359
0 8802 7 1 2 85356 8801
0 8803 5 1 1 8802
0 8804 7 1 2 8793 8803
0 8805 7 1 2 8788 8804
0 8806 5 1 1 8805
0 8807 7 1 2 61438 8806
0 8808 5 1 1 8807
0 8809 7 1 2 8785 8808
0 8810 5 1 1 8809
0 8811 7 1 2 63333 8810
0 8812 5 1 1 8811
0 8813 7 2 2 82166 71867
0 8814 5 1 1 85361
0 8815 7 8 2 66641 62245
0 8816 7 1 2 82917 85363
0 8817 7 1 2 85362 8816
0 8818 5 2 1 8817
0 8819 7 6 2 67507 83088
0 8820 5 3 1 85373
0 8821 7 1 2 68255 85109
0 8822 5 5 1 8821
0 8823 7 2 2 83117 85382
0 8824 7 1 2 84904 85387
0 8825 5 1 1 8824
0 8826 7 1 2 85379 8825
0 8827 5 1 1 8826
0 8828 7 1 2 72687 8827
0 8829 5 1 1 8828
0 8830 7 1 2 73611 82364
0 8831 5 2 1 8830
0 8832 7 1 2 67872 73159
0 8833 5 1 1 8832
0 8834 7 1 2 85389 8833
0 8835 5 1 1 8834
0 8836 7 1 2 71961 8835
0 8837 5 1 1 8836
0 8838 7 1 2 85222 8837
0 8839 5 1 1 8838
0 8840 7 1 2 63334 8839
0 8841 5 1 1 8840
0 8842 7 1 2 8829 8841
0 8843 5 1 1 8842
0 8844 7 1 2 81149 8843
0 8845 5 1 1 8844
0 8846 7 1 2 85371 8845
0 8847 5 1 1 8846
0 8848 7 1 2 63664 8847
0 8849 5 1 1 8848
0 8850 7 1 2 72688 85268
0 8851 5 1 1 8850
0 8852 7 1 2 77154 85319
0 8853 5 1 1 8852
0 8854 7 1 2 8851 8853
0 8855 5 1 1 8854
0 8856 7 1 2 85388 8855
0 8857 5 1 1 8856
0 8858 7 1 2 72689 85320
0 8859 5 1 1 8858
0 8860 7 1 2 8682 8859
0 8861 5 2 1 8860
0 8862 7 5 2 63335 77393
0 8863 7 1 2 85391 85393
0 8864 5 1 1 8863
0 8865 7 1 2 8857 8864
0 8866 5 1 1 8865
0 8867 7 1 2 62246 8866
0 8868 5 1 1 8867
0 8869 7 4 2 78735 78245
0 8870 5 4 1 85398
0 8871 7 5 2 65341 67247
0 8872 5 2 1 85406
0 8873 7 1 2 85298 85407
0 8874 7 1 2 85399 8873
0 8875 5 1 1 8874
0 8876 7 1 2 8868 8875
0 8877 5 1 1 8876
0 8878 7 1 2 71755 8877
0 8879 5 1 1 8878
0 8880 7 3 2 62530 77728
0 8881 5 1 1 85413
0 8882 7 1 2 61234 78077
0 8883 5 5 1 8882
0 8884 7 1 2 72690 85416
0 8885 5 1 1 8884
0 8886 7 3 2 70477 73160
0 8887 5 1 1 85421
0 8888 7 1 2 77840 8887
0 8889 7 1 2 8885 8888
0 8890 5 1 1 8889
0 8891 7 1 2 71962 8890
0 8892 5 1 1 8891
0 8893 7 1 2 8881 8892
0 8894 5 1 1 8893
0 8895 7 1 2 77887 8894
0 8896 5 1 1 8895
0 8897 7 7 2 62042 77761
0 8898 5 2 1 85424
0 8899 7 2 2 71963 78002
0 8900 7 1 2 85425 85433
0 8901 5 1 1 8900
0 8902 7 1 2 8896 8901
0 8903 5 1 1 8902
0 8904 7 1 2 85321 8903
0 8905 5 1 1 8904
0 8906 7 1 2 8879 8905
0 8907 7 1 2 8849 8906
0 8908 5 1 1 8907
0 8909 7 1 2 79511 8908
0 8910 5 1 1 8909
0 8911 7 1 2 8812 8910
0 8912 7 1 2 8741 8911
0 8913 5 1 1 8912
0 8914 7 1 2 63913 8913
0 8915 5 1 1 8914
0 8916 7 2 2 63336 82365
0 8917 7 1 2 79198 79221
0 8918 5 1 1 8917
0 8919 7 1 2 78070 84922
0 8920 5 1 1 8919
0 8921 7 1 2 8918 8920
0 8922 5 1 1 8921
0 8923 7 1 2 66179 8922
0 8924 5 1 1 8923
0 8925 7 1 2 76126 79199
0 8926 7 1 2 77875 8925
0 8927 5 1 1 8926
0 8928 7 1 2 8924 8927
0 8929 5 1 1 8928
0 8930 7 1 2 80396 8929
0 8931 5 1 1 8930
0 8932 7 1 2 61235 85392
0 8933 5 1 1 8932
0 8934 7 1 2 66180 84303
0 8935 7 1 2 84416 8934
0 8936 5 1 1 8935
0 8937 7 1 2 8933 8936
0 8938 5 1 1 8937
0 8939 7 1 2 79512 8938
0 8940 5 1 1 8939
0 8941 7 21 2 60445 66405
0 8942 5 6 1 85437
0 8943 7 5 2 61649 85438
0 8944 7 3 2 79120 85464
0 8945 7 1 2 85181 85469
0 8946 5 1 1 8945
0 8947 7 2 2 65342 83646
0 8948 5 2 1 85472
0 8949 7 1 2 80320 85473
0 8950 5 1 1 8949
0 8951 7 6 2 65112 85439
0 8952 5 2 1 85476
0 8953 7 1 2 85477 85194
0 8954 5 1 1 8953
0 8955 7 1 2 8950 8954
0 8956 5 1 1 8955
0 8957 7 1 2 64904 8956
0 8958 5 1 1 8957
0 8959 7 2 2 81075 85195
0 8960 5 1 1 85484
0 8961 7 1 2 75178 85485
0 8962 5 1 1 8961
0 8963 7 1 2 8958 8962
0 8964 5 1 1 8963
0 8965 7 1 2 71075 8964
0 8966 5 1 1 8965
0 8967 7 1 2 8946 8966
0 8968 7 1 2 8940 8967
0 8969 7 1 2 8931 8968
0 8970 5 1 1 8969
0 8971 7 1 2 85435 8970
0 8972 5 1 1 8971
0 8973 7 1 2 84242 78501
0 8974 5 1 1 8973
0 8975 7 1 2 77827 84221
0 8976 5 1 1 8975
0 8977 7 1 2 8974 8976
0 8978 5 1 1 8977
0 8979 7 6 2 63665 83731
0 8980 7 1 2 8978 85486
0 8981 5 1 1 8980
0 8982 7 1 2 8972 8981
0 8983 5 2 1 8982
0 8984 7 1 2 63914 85492
0 8985 5 1 1 8984
0 8986 7 3 2 80974 77223
0 8987 7 4 2 62878 74926
0 8988 7 42 2 63666 68831
0 8989 5 4 1 85501
0 8990 7 8 2 63337 85502
0 8991 5 1 1 85547
0 8992 7 2 2 85497 85548
0 8993 7 1 2 66642 85555
0 8994 7 1 2 85494 8993
0 8995 5 1 1 8994
0 8996 7 1 2 8985 8995
0 8997 5 1 1 8996
0 8998 7 1 2 74051 8997
0 8999 5 1 1 8998
0 9000 7 1 2 61838 8999
0 9001 7 1 2 8915 9000
0 9002 5 1 1 9001
0 9003 7 1 2 8563 9002
0 9004 5 1 1 9003
0 9005 7 1 2 65538 9004
0 9006 5 1 1 9005
0 9007 7 1 2 78849 85232
0 9008 5 1 1 9007
0 9009 7 1 2 64905 85254
0 9010 5 1 1 9009
0 9011 7 2 2 65113 78866
0 9012 5 3 1 85557
0 9013 7 5 2 66181 82366
0 9014 5 3 1 85562
0 9015 7 1 2 60246 85563
0 9016 5 1 1 9015
0 9017 7 1 2 85559 9016
0 9018 7 1 2 9010 9017
0 9019 5 1 1 9018
0 9020 7 1 2 71076 9019
0 9021 5 1 1 9020
0 9022 7 2 2 62879 75739
0 9023 5 1 1 85570
0 9024 7 1 2 65114 85571
0 9025 5 1 1 9024
0 9026 7 1 2 9021 9025
0 9027 5 1 1 9026
0 9028 7 1 2 84905 9027
0 9029 5 1 1 9028
0 9030 7 1 2 9008 9029
0 9031 5 1 1 9030
0 9032 7 1 2 66406 9031
0 9033 5 1 1 9032
0 9034 7 1 2 71278 85237
0 9035 5 1 1 9034
0 9036 7 1 2 9033 9035
0 9037 5 1 1 9036
0 9038 7 1 2 68256 9037
0 9039 5 1 1 9038
0 9040 7 3 2 71077 77419
0 9041 5 1 1 85572
0 9042 7 1 2 85390 9041
0 9043 5 1 1 9042
0 9044 7 1 2 71964 9043
0 9045 5 1 1 9044
0 9046 7 1 2 67508 79063
0 9047 5 1 1 9046
0 9048 7 1 2 9045 9047
0 9049 5 1 1 9048
0 9050 7 2 2 63338 9049
0 9051 5 1 1 85575
0 9052 7 1 2 84932 85576
0 9053 5 1 1 9052
0 9054 7 1 2 9039 9053
0 9055 5 1 1 9054
0 9056 7 1 2 81150 9055
0 9057 5 1 1 9056
0 9058 7 3 2 62880 74336
0 9059 5 1 1 85577
0 9060 7 1 2 74216 85578
0 9061 5 1 1 9060
0 9062 7 1 2 61439 77950
0 9063 5 1 1 9062
0 9064 7 1 2 9061 9063
0 9065 5 1 1 9064
0 9066 7 1 2 64906 9065
0 9067 5 1 1 9066
0 9068 7 4 2 60247 79553
0 9069 5 2 1 85580
0 9070 7 1 2 85426 85581
0 9071 5 1 1 9070
0 9072 7 1 2 9067 9071
0 9073 5 1 1 9072
0 9074 7 1 2 71078 9073
0 9075 5 1 1 9074
0 9076 7 1 2 82021 85427
0 9077 5 1 1 9076
0 9078 7 1 2 9075 9077
0 9079 5 1 1 9078
0 9080 7 1 2 81151 9079
0 9081 5 1 1 9080
0 9082 7 4 2 65343 74673
0 9083 7 8 2 60248 66643
0 9084 7 1 2 85428 85590
0 9085 7 1 2 85586 9084
0 9086 5 1 1 9085
0 9087 7 1 2 60446 81118
0 9088 7 1 2 71279 9087
0 9089 5 1 1 9088
0 9090 7 1 2 9086 9089
0 9091 7 1 2 9081 9090
0 9092 5 1 1 9091
0 9093 7 1 2 76626 9092
0 9094 5 1 1 9093
0 9095 7 3 2 82601 79429
0 9096 5 1 1 85598
0 9097 7 1 2 78366 85599
0 9098 7 1 2 85279 9097
0 9099 5 1 1 9098
0 9100 7 1 2 9094 9099
0 9101 5 1 1 9100
0 9102 7 1 2 71756 9101
0 9103 5 1 1 9102
0 9104 7 8 2 62043 77455
0 9105 7 1 2 85025 85601
0 9106 5 1 1 9105
0 9107 7 1 2 9051 9106
0 9108 5 1 1 9107
0 9109 7 1 2 81152 9108
0 9110 5 1 1 9109
0 9111 7 2 2 65344 78246
0 9112 5 1 1 85609
0 9113 7 2 2 73661 79430
0 9114 7 1 2 85610 85611
0 9115 5 1 1 9114
0 9116 7 4 2 76837 77762
0 9117 5 2 1 85613
0 9118 7 2 2 64907 85614
0 9119 5 1 1 85619
0 9120 7 1 2 71079 77888
0 9121 5 1 1 9120
0 9122 7 1 2 9119 9121
0 9123 5 1 1 9122
0 9124 7 1 2 62247 85311
0 9125 7 1 2 9123 9124
0 9126 5 1 1 9125
0 9127 7 1 2 9115 9126
0 9128 5 1 1 9127
0 9129 7 1 2 71757 9128
0 9130 5 1 1 9129
0 9131 7 1 2 85372 9130
0 9132 7 1 2 9110 9131
0 9133 5 1 1 9132
0 9134 7 1 2 79513 9133
0 9135 5 1 1 9134
0 9136 7 4 2 65345 83732
0 9137 5 3 1 85621
0 9138 7 2 2 80179 85622
0 9139 5 2 1 85628
0 9140 7 1 2 62248 85629
0 9141 5 2 1 9140
0 9142 7 2 2 80017 81725
0 9143 7 1 2 82008 85634
0 9144 5 1 1 9143
0 9145 7 1 2 85632 9144
0 9146 5 1 1 9145
0 9147 7 1 2 84906 9146
0 9148 5 1 1 9147
0 9149 7 2 2 68257 85233
0 9150 7 1 2 84229 85636
0 9151 5 2 1 9150
0 9152 7 7 2 66407 80557
0 9153 5 1 1 85640
0 9154 7 2 2 84696 85641
0 9155 7 1 2 66182 85647
0 9156 5 1 1 9155
0 9157 7 1 2 85633 9156
0 9158 5 1 1 9157
0 9159 7 1 2 64908 9158
0 9160 5 1 1 9159
0 9161 7 1 2 85638 9160
0 9162 7 1 2 9148 9161
0 9163 5 1 1 9162
0 9164 7 1 2 71080 9163
0 9165 5 1 1 9164
0 9166 7 1 2 84731 85470
0 9167 5 1 1 9166
0 9168 7 4 2 65346 61236
0 9169 7 3 2 60249 85649
0 9170 7 1 2 80162 81523
0 9171 7 1 2 85653 9170
0 9172 5 1 1 9171
0 9173 7 1 2 9167 9172
0 9174 5 1 1 9173
0 9175 7 5 2 64437 62881
0 9176 7 1 2 72763 85656
0 9177 7 1 2 9174 9176
0 9178 5 1 1 9177
0 9179 7 1 2 9165 9178
0 9180 7 1 2 9135 9179
0 9181 7 1 2 9103 9180
0 9182 7 1 2 9057 9181
0 9183 5 1 1 9182
0 9184 7 1 2 66792 9183
0 9185 5 1 1 9184
0 9186 7 1 2 62882 81925
0 9187 5 1 1 9186
0 9188 7 3 2 81687 74498
0 9189 5 2 1 85661
0 9190 7 1 2 9187 85664
0 9191 5 1 1 9190
0 9192 7 10 2 66408 61839
0 9193 7 12 2 66644 63339
0 9194 7 2 2 85666 85676
0 9195 5 3 1 85688
0 9196 7 1 2 81276 85689
0 9197 7 1 2 9191 9196
0 9198 5 1 1 9197
0 9199 7 1 2 9185 9198
0 9200 5 1 1 9199
0 9201 7 1 2 63667 9200
0 9202 5 1 1 9201
0 9203 7 24 2 66793 68611
0 9204 7 1 2 61237 85069
0 9205 5 1 1 9204
0 9206 7 1 2 78181 73729
0 9207 5 2 1 9206
0 9208 7 1 2 9205 85717
0 9209 5 1 1 9208
0 9210 7 1 2 73515 9209
0 9211 5 1 1 9210
0 9212 7 1 2 62883 85028
0 9213 5 1 1 9212
0 9214 7 1 2 9211 9213
0 9215 5 1 1 9214
0 9216 7 1 2 74217 9215
0 9217 5 1 1 9216
0 9218 7 1 2 8286 8498
0 9219 5 1 1 9218
0 9220 7 1 2 67873 9219
0 9221 5 1 1 9220
0 9222 7 1 2 66409 9221
0 9223 7 1 2 9217 9222
0 9224 5 1 1 9223
0 9225 7 1 2 70028 84976
0 9226 5 1 1 9225
0 9227 7 2 2 71965 84965
0 9228 5 1 1 85719
0 9229 7 1 2 9226 9228
0 9230 5 1 1 9229
0 9231 7 1 2 77889 9230
0 9232 5 1 1 9231
0 9233 7 2 2 81322 82674
0 9234 5 1 1 85721
0 9235 7 1 2 77763 74499
0 9236 7 1 2 85722 9235
0 9237 5 1 1 9236
0 9238 7 1 2 61440 9237
0 9239 7 1 2 9232 9238
0 9240 5 1 1 9239
0 9241 7 1 2 65115 9240
0 9242 7 1 2 9224 9241
0 9243 5 1 1 9242
0 9244 7 3 2 62531 77890
0 9245 5 2 1 85723
0 9246 7 1 2 74218 84654
0 9247 5 2 1 9246
0 9248 7 1 2 77938 85728
0 9249 5 2 1 9248
0 9250 7 1 2 69060 85730
0 9251 5 1 1 9250
0 9252 7 1 2 85726 9251
0 9253 5 1 1 9252
0 9254 7 1 2 84959 9253
0 9255 5 1 1 9254
0 9256 7 1 2 69229 77891
0 9257 5 2 1 9256
0 9258 7 1 2 80742 79064
0 9259 5 1 1 9258
0 9260 7 1 2 85732 9259
0 9261 5 1 1 9260
0 9262 7 1 2 84960 9261
0 9263 5 1 1 9262
0 9264 7 2 2 81045 84732
0 9265 5 2 1 85734
0 9266 7 1 2 67874 85735
0 9267 5 2 1 9266
0 9268 7 5 2 68258 79478
0 9269 7 1 2 60250 85740
0 9270 5 1 1 9269
0 9271 7 1 2 85738 9270
0 9272 5 1 1 9271
0 9273 7 1 2 70029 9272
0 9274 5 1 1 9273
0 9275 7 2 2 77892 85035
0 9276 5 1 1 85745
0 9277 7 1 2 78015 85746
0 9278 5 1 1 9277
0 9279 7 1 2 9274 9278
0 9280 5 1 1 9279
0 9281 7 1 2 76696 78525
0 9282 7 1 2 9280 9281
0 9283 5 1 1 9282
0 9284 7 1 2 9263 9283
0 9285 5 1 1 9284
0 9286 7 1 2 64438 9285
0 9287 5 1 1 9286
0 9288 7 1 2 9255 9287
0 9289 7 1 2 9243 9288
0 9290 5 1 1 9289
0 9291 7 1 2 66645 9290
0 9292 5 1 1 9291
0 9293 7 1 2 79468 81119
0 9294 7 1 2 85720 9293
0 9295 5 1 1 9294
0 9296 7 1 2 9292 9295
0 9297 5 1 1 9296
0 9298 7 1 2 65347 9297
0 9299 5 1 1 9298
0 9300 7 1 2 80558 77068
0 9301 7 1 2 84954 9300
0 9302 7 2 2 66183 80990
0 9303 7 3 2 62044 84733
0 9304 7 1 2 85747 85749
0 9305 7 1 2 9301 9304
0 9306 5 1 1 9305
0 9307 7 1 2 9299 9306
0 9308 5 1 1 9307
0 9309 7 1 2 85693 9308
0 9310 5 1 1 9309
0 9311 7 1 2 75134 85731
0 9312 5 1 1 9311
0 9313 7 2 2 60251 80018
0 9314 5 5 1 85752
0 9315 7 1 2 67875 85753
0 9316 5 1 1 9315
0 9317 7 1 2 9312 9316
0 9318 5 1 1 9317
0 9319 7 1 2 82568 9318
0 9320 5 1 1 9319
0 9321 7 3 2 67876 80724
0 9322 7 2 2 84646 84854
0 9323 7 1 2 85759 85762
0 9324 5 1 1 9323
0 9325 7 1 2 9320 9324
0 9326 5 1 1 9325
0 9327 7 1 2 62532 9326
0 9328 5 1 1 9327
0 9329 7 2 2 83089 73629
0 9330 7 1 2 84876 85764
0 9331 5 1 1 9330
0 9332 7 1 2 9328 9331
0 9333 5 1 1 9332
0 9334 7 1 2 80397 9333
0 9335 5 1 1 9334
0 9336 7 4 2 62533 83733
0 9337 7 1 2 84230 85766
0 9338 5 1 1 9337
0 9339 7 3 2 64683 83090
0 9340 7 8 2 61650 62045
0 9341 7 1 2 65968 85773
0 9342 7 1 2 85478 9341
0 9343 7 1 2 85770 9342
0 9344 5 1 1 9343
0 9345 7 1 2 9338 9344
0 9346 5 1 1 9345
0 9347 7 1 2 75952 9346
0 9348 5 1 1 9347
0 9349 7 1 2 85639 9348
0 9350 7 1 2 9335 9349
0 9351 5 1 1 9350
0 9352 7 1 2 63668 9351
0 9353 5 1 1 9352
0 9354 7 1 2 77420 85208
0 9355 5 1 1 9354
0 9356 7 6 2 61651 79368
0 9357 5 1 1 85781
0 9358 7 1 2 67509 85782
0 9359 5 1 1 9358
0 9360 7 1 2 9355 9359
0 9361 5 1 1 9360
0 9362 7 1 2 65348 9361
0 9363 5 1 1 9362
0 9364 7 1 2 78182 84891
0 9365 5 1 1 9364
0 9366 7 1 2 9363 9365
0 9367 5 1 1 9366
0 9368 7 1 2 66410 3865
0 9369 5 2 1 9368
0 9370 7 1 2 65116 79928
0 9371 7 1 2 85787 9370
0 9372 5 1 1 9371
0 9373 7 1 2 85754 9372
0 9374 5 1 1 9373
0 9375 7 1 2 9367 9374
0 9376 5 1 1 9375
0 9377 7 1 2 65969 76984
0 9378 5 6 1 9377
0 9379 7 1 2 70960 85789
0 9380 5 1 1 9379
0 9381 7 1 2 64439 9380
0 9382 5 1 1 9381
0 9383 7 1 2 77289 76697
0 9384 5 4 1 9383
0 9385 7 1 2 9382 85795
0 9386 5 1 1 9385
0 9387 7 1 2 80154 9386
0 9388 5 1 1 9387
0 9389 7 3 2 71966 79530
0 9390 5 1 1 85799
0 9391 7 1 2 81210 85800
0 9392 5 1 1 9391
0 9393 7 1 2 9388 9392
0 9394 5 1 1 9393
0 9395 7 1 2 84395 9394
0 9396 5 1 1 9395
0 9397 7 1 2 9376 9396
0 9398 7 1 2 9353 9397
0 9399 5 1 1 9398
0 9400 7 1 2 66794 9399
0 9401 5 1 1 9400
0 9402 7 3 2 61840 62046
0 9403 7 4 2 66646 85802
0 9404 7 3 2 79398 85805
0 9405 7 8 2 65803 62884
0 9406 5 3 1 85812
0 9407 7 2 2 64684 85813
0 9408 7 4 2 65349 62249
0 9409 7 1 2 79423 85825
0 9410 7 1 2 85823 9409
0 9411 7 1 2 85809 9410
0 9412 5 1 1 9411
0 9413 7 1 2 9401 9412
0 9414 5 1 1 9413
0 9415 7 1 2 70741 9414
0 9416 5 1 1 9415
0 9417 7 1 2 9310 9416
0 9418 7 1 2 9202 9417
0 9419 5 1 1 9418
0 9420 7 1 2 63915 9419
0 9421 5 1 1 9420
0 9422 7 1 2 66795 85493
0 9423 5 1 1 9422
0 9424 7 4 2 65117 77729
0 9425 5 1 1 85829
0 9426 7 3 2 75678 79369
0 9427 7 21 2 66647 61841
0 9428 5 3 1 85836
0 9429 7 3 2 65350 85837
0 9430 5 2 1 85860
0 9431 7 1 2 75410 85861
0 9432 7 1 2 85833 9431
0 9433 7 1 2 85830 9432
0 9434 5 1 1 9433
0 9435 7 1 2 9423 9434
0 9436 5 1 1 9435
0 9437 7 1 2 63916 9436
0 9438 5 1 1 9437
0 9439 7 4 2 80527 79370
0 9440 7 5 2 66796 62534
0 9441 7 3 2 80991 85869
0 9442 7 1 2 85865 85874
0 9443 7 1 2 85495 9442
0 9444 5 1 1 9443
0 9445 7 1 2 9438 9444
0 9446 5 1 1 9445
0 9447 7 1 2 74052 9446
0 9448 5 1 1 9447
0 9449 7 1 2 60647 9448
0 9450 7 1 2 9421 9449
0 9451 5 1 1 9450
0 9452 7 1 2 69631 9451
0 9453 7 1 2 9006 9452
0 9454 5 1 1 9453
0 9455 7 8 2 60648 63917
0 9456 7 3 2 68259 69897
0 9457 5 1 1 85885
0 9458 7 3 2 81215 9457
0 9459 5 1 1 85888
0 9460 7 1 2 84996 85889
0 9461 5 1 1 9460
0 9462 7 2 2 64223 71020
0 9463 7 32 2 61441 68260
0 9464 5 10 1 85893
0 9465 7 1 2 81631 85894
0 9466 7 1 2 85891 9465
0 9467 5 1 1 9466
0 9468 7 1 2 84998 9467
0 9469 5 1 1 9468
0 9470 7 1 2 71081 9469
0 9471 5 1 1 9470
0 9472 7 1 2 85021 9471
0 9473 7 1 2 9461 9472
0 9474 5 1 1 9473
0 9475 7 1 2 62885 9474
0 9476 5 1 1 9475
0 9477 7 2 2 61013 74989
0 9478 5 2 1 85935
0 9479 7 1 2 77730 81865
0 9480 5 1 1 9479
0 9481 7 1 2 85937 9480
0 9482 5 1 1 9481
0 9483 7 1 2 75179 78280
0 9484 7 1 2 9482 9483
0 9485 5 1 1 9484
0 9486 7 1 2 9476 9485
0 9487 5 1 1 9486
0 9488 7 1 2 65804 9487
0 9489 5 1 1 9488
0 9490 7 11 2 62535 77764
0 9491 5 7 1 85939
0 9492 7 1 2 82022 85940
0 9493 5 1 1 9492
0 9494 7 1 2 81552 85059
0 9495 5 2 1 9494
0 9496 7 3 2 73223 77893
0 9497 7 1 2 70742 85959
0 9498 5 2 1 9497
0 9499 7 1 2 85957 85962
0 9500 5 1 1 9499
0 9501 7 1 2 79514 9500
0 9502 5 1 1 9501
0 9503 7 1 2 9493 9502
0 9504 5 1 1 9503
0 9505 7 1 2 65970 9504
0 9506 5 1 1 9505
0 9507 7 4 2 66184 77765
0 9508 5 4 1 85964
0 9509 7 2 2 61238 77894
0 9510 5 5 1 85972
0 9511 7 1 2 85968 85974
0 9512 5 1 1 9511
0 9513 7 2 2 61014 9512
0 9514 7 1 2 84030 85979
0 9515 5 1 1 9514
0 9516 7 1 2 9506 9515
0 9517 5 1 1 9516
0 9518 7 1 2 64685 9517
0 9519 5 1 1 9518
0 9520 7 1 2 75180 73922
0 9521 5 1 1 9520
0 9522 7 1 2 82017 9521
0 9523 5 1 1 9522
0 9524 7 1 2 85960 9523
0 9525 5 1 1 9524
0 9526 7 1 2 9519 9525
0 9527 7 1 2 9489 9526
0 9528 5 1 1 9527
0 9529 7 1 2 68612 9528
0 9530 5 1 1 9529
0 9531 7 4 2 62047 72488
0 9532 5 2 1 85981
0 9533 7 1 2 67877 85985
0 9534 5 2 1 9533
0 9535 7 3 2 60252 78584
0 9536 5 3 1 85989
0 9537 7 2 2 61442 85990
0 9538 5 2 1 85995
0 9539 7 4 2 62536 78736
0 9540 7 2 2 76819 85999
0 9541 7 1 2 85996 86003
0 9542 7 1 2 85987 9541
0 9543 5 1 1 9542
0 9544 7 1 2 9530 9543
0 9545 5 1 1 9544
0 9546 7 1 2 79607 9545
0 9547 5 1 1 9546
0 9548 7 2 2 65971 78546
0 9549 7 6 2 77069 86005
0 9550 5 6 1 86007
0 9551 7 1 2 78924 86013
0 9552 5 1 1 9551
0 9553 7 1 2 79034 9552
0 9554 7 2 2 79600 9553
0 9555 7 1 2 80569 86019
0 9556 5 1 1 9555
0 9557 7 1 2 83946 85159
0 9558 5 1 1 9557
0 9559 7 1 2 75135 78964
0 9560 5 1 1 9559
0 9561 7 1 2 61443 78585
0 9562 5 4 1 9561
0 9563 7 3 2 67018 78586
0 9564 5 2 1 86025
0 9565 7 4 2 86021 86028
0 9566 7 1 2 60253 79496
0 9567 7 1 2 86030 9566
0 9568 5 1 1 9567
0 9569 7 1 2 9560 9568
0 9570 5 1 1 9569
0 9571 7 1 2 72691 9570
0 9572 5 1 1 9571
0 9573 7 1 2 9558 9572
0 9574 5 1 1 9573
0 9575 7 1 2 85182 9574
0 9576 5 1 1 9575
0 9577 7 1 2 2989 9576
0 9578 5 1 1 9577
0 9579 7 1 2 72543 9578
0 9580 5 1 1 9579
0 9581 7 1 2 78906 85223
0 9582 5 1 1 9581
0 9583 7 1 2 77828 9582
0 9584 5 1 1 9583
0 9585 7 5 2 62886 77961
0 9586 7 1 2 67510 86034
0 9587 5 1 1 9586
0 9588 7 1 2 9584 9587
0 9589 5 1 1 9588
0 9590 7 1 2 61444 9589
0 9591 5 1 1 9590
0 9592 7 3 2 74726 78123
0 9593 5 1 1 86039
0 9594 7 1 2 85276 86040
0 9595 5 1 1 9594
0 9596 7 1 2 78203 1939
0 9597 5 3 1 9596
0 9598 7 1 2 79322 72692
0 9599 7 1 2 86042 9598
0 9600 5 1 1 9599
0 9601 7 1 2 9595 9600
0 9602 7 1 2 9591 9601
0 9603 5 1 1 9602
0 9604 7 1 2 63669 9603
0 9605 5 1 1 9604
0 9606 7 1 2 9580 9605
0 9607 5 1 1 9606
0 9608 7 1 2 63340 9607
0 9609 5 1 1 9608
0 9610 7 1 2 65118 86031
0 9611 5 2 1 9610
0 9612 7 1 2 3136 86045
0 9613 5 4 1 9612
0 9614 7 1 2 72693 5378
0 9615 7 1 2 86047 9614
0 9616 5 1 1 9615
0 9617 7 2 2 79497 79583
0 9618 7 1 2 85282 86051
0 9619 5 1 1 9618
0 9620 7 1 2 83947 85286
0 9621 5 1 1 9620
0 9622 7 1 2 9619 9621
0 9623 7 1 2 9616 9622
0 9624 5 1 1 9623
0 9625 7 1 2 86004 9624
0 9626 5 1 1 9625
0 9627 7 1 2 9609 9626
0 9628 5 1 1 9627
0 9629 7 1 2 81153 9628
0 9630 5 1 1 9629
0 9631 7 1 2 9556 9630
0 9632 7 1 2 9547 9631
0 9633 5 1 1 9632
0 9634 7 1 2 66797 9633
0 9635 5 1 1 9634
0 9636 7 7 2 65119 80992
0 9637 7 5 2 65351 61842
0 9638 7 3 2 86053 86060
0 9639 5 2 1 86065
0 9640 7 1 2 86020 86066
0 9641 5 1 1 9640
0 9642 7 1 2 9635 9641
0 9643 5 1 1 9642
0 9644 7 1 2 85877 9643
0 9645 5 1 1 9644
0 9646 7 48 2 61843 63918
0 9647 5 8 1 86070
0 9648 7 1 2 72694 86071
0 9649 5 2 1 9648
0 9650 7 5 2 62537 68832
0 9651 7 4 2 66798 86128
0 9652 7 1 2 60085 69779
0 9653 7 1 2 79243 9652
0 9654 7 1 2 86133 9653
0 9655 5 1 1 9654
0 9656 7 1 2 86126 9655
0 9657 5 1 1 9656
0 9658 7 1 2 61239 9657
0 9659 5 1 1 9658
0 9660 7 3 2 59825 66799
0 9661 7 1 2 68833 76017
0 9662 7 1 2 86137 9661
0 9663 5 1 1 9662
0 9664 7 1 2 86118 9663
0 9665 5 1 1 9664
0 9666 7 1 2 73734 9665
0 9667 5 1 1 9666
0 9668 7 1 2 9659 9667
0 9669 5 1 1 9668
0 9670 7 1 2 84329 9669
0 9671 5 1 1 9670
0 9672 7 7 2 67019 68834
0 9673 7 3 2 66800 86140
0 9674 7 1 2 71082 86147
0 9675 5 1 1 9674
0 9676 7 1 2 86119 9675
0 9677 5 1 1 9676
0 9678 7 1 2 76127 84471
0 9679 7 1 2 9677 9678
0 9680 5 1 1 9679
0 9681 7 1 2 9671 9680
0 9682 5 1 1 9681
0 9683 7 1 2 63341 9682
0 9684 5 1 1 9683
0 9685 7 1 2 72695 85196
0 9686 5 1 1 9685
0 9687 7 1 2 77155 84330
0 9688 5 1 1 9687
0 9689 7 1 2 9686 9688
0 9690 5 1 1 9689
0 9691 7 1 2 69780 86072
0 9692 7 1 2 9690 9691
0 9693 5 1 1 9692
0 9694 7 44 2 66801 68835
0 9695 5 1 1 86150
0 9696 7 1 2 81968 86151
0 9697 7 1 2 85214 9696
0 9698 5 1 1 9697
0 9699 7 1 2 9693 9698
0 9700 5 1 1 9699
0 9701 7 1 2 77599 9700
0 9702 5 1 1 9701
0 9703 7 1 2 9684 9702
0 9704 5 1 1 9703
0 9705 7 1 2 65805 9704
0 9706 5 1 1 9705
0 9707 7 3 2 77539 85838
0 9708 5 1 1 86194
0 9709 7 4 2 68261 86195
0 9710 5 1 1 86197
0 9711 7 1 2 77845 86198
0 9712 5 1 1 9711
0 9713 7 5 2 66802 81785
0 9714 7 1 2 77619 86201
0 9715 5 1 1 9714
0 9716 7 10 2 61844 63342
0 9717 7 3 2 63919 86206
0 9718 7 1 2 61240 86216
0 9719 5 1 1 9718
0 9720 7 1 2 9715 9719
0 9721 5 1 1 9720
0 9722 7 1 2 83826 9721
0 9723 5 1 1 9722
0 9724 7 5 2 67511 63920
0 9725 7 3 2 61845 86219
0 9726 7 1 2 63343 72696
0 9727 7 1 2 86224 9726
0 9728 5 1 1 9727
0 9729 7 1 2 9723 9728
0 9730 5 1 1 9729
0 9731 7 1 2 84472 9730
0 9732 5 1 1 9731
0 9733 7 1 2 9712 9732
0 9734 7 1 2 9706 9733
0 9735 5 1 1 9734
0 9736 7 1 2 79515 9735
0 9737 5 1 1 9736
0 9738 7 2 2 75181 85839
0 9739 5 1 1 86227
0 9740 7 8 2 60254 61652
0 9741 7 8 2 61445 66803
0 9742 7 1 2 86229 86237
0 9743 5 3 1 9742
0 9744 7 1 2 9739 86245
0 9745 5 3 1 9744
0 9746 7 2 2 68613 86248
0 9747 7 1 2 77654 86251
0 9748 5 1 1 9747
0 9749 7 1 2 77629 86252
0 9750 5 1 1 9749
0 9751 7 1 2 75147 821
0 9752 5 1 1 9751
0 9753 7 12 2 61846 62538
0 9754 7 3 2 63670 86253
0 9755 7 1 2 77070 84250
0 9756 7 1 2 86265 9755
0 9757 7 1 2 9752 9756
0 9758 5 1 1 9757
0 9759 7 1 2 9750 9758
0 9760 5 1 1 9759
0 9761 7 1 2 76820 9760
0 9762 5 1 1 9761
0 9763 7 1 2 9748 9762
0 9764 5 1 1 9763
0 9765 7 1 2 68262 9764
0 9766 5 1 1 9765
0 9767 7 3 2 61446 78153
0 9768 5 1 1 86268
0 9769 7 2 2 80650 85204
0 9770 7 1 2 65972 78949
0 9771 7 1 2 86271 9770
0 9772 5 1 1 9771
0 9773 7 1 2 9768 9772
0 9774 5 1 1 9773
0 9775 7 1 2 65120 9774
0 9776 5 1 1 9775
0 9777 7 1 2 71083 77019
0 9778 5 2 1 9777
0 9779 7 1 2 72544 79222
0 9780 5 1 1 9779
0 9781 7 1 2 86273 9780
0 9782 5 1 1 9781
0 9783 7 1 2 79200 9782
0 9784 5 1 1 9783
0 9785 7 1 2 9776 9784
0 9786 5 1 1 9785
0 9787 7 1 2 66185 9786
0 9788 5 1 1 9787
0 9789 7 1 2 79201 85277
0 9790 7 1 2 78922 9789
0 9791 5 1 1 9790
0 9792 7 1 2 9788 9791
0 9793 5 1 1 9792
0 9794 7 12 2 61653 61847
0 9795 7 1 2 63344 86275
0 9796 7 1 2 9793 9795
0 9797 5 1 1 9796
0 9798 7 1 2 9766 9797
0 9799 5 1 1 9798
0 9800 7 1 2 63921 9799
0 9801 5 1 1 9800
0 9802 7 6 2 64909 82104
0 9803 5 2 1 86287
0 9804 7 3 2 83516 86288
0 9805 7 1 2 69781 86295
0 9806 5 1 1 9805
0 9807 7 11 2 68263 70589
0 9808 7 1 2 84001 86298
0 9809 5 1 1 9808
0 9810 7 1 2 9806 9809
0 9811 5 1 1 9810
0 9812 7 9 2 66804 62048
0 9813 7 3 2 86129 86309
0 9814 7 1 2 9811 86318
0 9815 5 1 1 9814
0 9816 7 1 2 86296 86073
0 9817 5 1 1 9816
0 9818 7 1 2 9815 9817
0 9819 5 1 1 9818
0 9820 7 1 2 71084 9819
0 9821 5 1 1 9820
0 9822 7 8 2 61848 68264
0 9823 7 4 2 63922 86321
0 9824 7 2 2 85183 86329
0 9825 7 2 2 69782 77337
0 9826 7 1 2 86333 86335
0 9827 5 1 1 9826
0 9828 7 1 2 9821 9827
0 9829 5 1 1 9828
0 9830 7 1 2 80188 9829
0 9831 5 1 1 9830
0 9832 7 5 2 65806 66648
0 9833 7 1 2 72204 86337
0 9834 7 1 2 73959 9833
0 9835 7 2 2 68836 85694
0 9836 7 3 2 74337 72749
0 9837 5 1 1 86344
0 9838 7 1 2 86342 86345
0 9839 7 1 2 9834 9838
0 9840 5 1 1 9839
0 9841 7 1 2 62887 9840
0 9842 7 1 2 9831 9841
0 9843 7 1 2 9801 9842
0 9844 7 1 2 9737 9843
0 9845 5 1 1 9844
0 9846 7 1 2 78509 86225
0 9847 5 1 1 9846
0 9848 7 1 2 66186 73316
0 9849 7 1 2 86134 9848
0 9850 5 1 1 9849
0 9851 7 1 2 9847 9850
0 9852 5 1 1 9851
0 9853 7 1 2 64686 9852
0 9854 5 1 1 9853
0 9855 7 1 2 81582 86135
0 9856 5 1 1 9855
0 9857 7 3 2 65807 63923
0 9858 7 10 2 61849 67512
0 9859 7 1 2 86347 86350
0 9860 5 1 1 9859
0 9861 7 1 2 9856 9860
0 9862 5 1 1 9861
0 9863 7 1 2 66187 9862
0 9864 5 1 1 9863
0 9865 7 1 2 9854 9864
0 9866 5 1 1 9865
0 9867 7 1 2 84331 9866
0 9868 5 1 1 9867
0 9869 7 6 2 65808 61654
0 9870 7 2 2 85184 86074
0 9871 7 1 2 86360 86366
0 9872 5 1 1 9871
0 9873 7 1 2 9868 9872
0 9874 5 1 1 9873
0 9875 7 1 2 66411 9874
0 9876 5 1 1 9875
0 9877 7 7 2 63924 79706
0 9878 7 4 2 66188 78510
0 9879 7 1 2 62539 79425
0 9880 7 1 2 86375 9879
0 9881 7 1 2 86368 9880
0 9882 5 1 1 9881
0 9883 7 1 2 9876 9882
0 9884 5 1 1 9883
0 9885 7 1 2 65121 9884
0 9886 5 1 1 9885
0 9887 7 10 2 66412 63671
0 9888 7 1 2 86254 86379
0 9889 7 1 2 77713 9888
0 9890 5 1 1 9889
0 9891 7 5 2 66805 67513
0 9892 7 1 2 75474 86389
0 9893 7 1 2 85167 9892
0 9894 5 1 1 9893
0 9895 7 1 2 9890 9894
0 9896 5 1 1 9895
0 9897 7 1 2 61655 9896
0 9898 5 1 1 9897
0 9899 7 1 2 80321 86266
0 9900 5 1 1 9899
0 9901 7 1 2 9898 9900
0 9902 5 1 1 9901
0 9903 7 1 2 86348 9902
0 9904 5 1 1 9903
0 9905 7 1 2 9886 9904
0 9906 5 1 1 9905
0 9907 7 1 2 68265 9906
0 9908 5 1 1 9907
0 9909 7 1 2 66649 85168
0 9910 5 1 1 9909
0 9911 7 1 2 85202 9910
0 9912 5 1 1 9911
0 9913 7 1 2 79323 9912
0 9914 5 1 1 9913
0 9915 7 1 2 78800 71085
0 9916 7 1 2 85197 9915
0 9917 5 1 1 9916
0 9918 7 1 2 9914 9917
0 9919 5 1 1 9918
0 9920 7 1 2 86217 9919
0 9921 5 1 1 9920
0 9922 7 1 2 9908 9921
0 9923 5 1 1 9922
0 9924 7 1 2 64910 9923
0 9925 5 1 1 9924
0 9926 7 2 2 67514 86249
0 9927 7 8 2 65973 76698
0 9928 5 1 1 86396
0 9929 7 1 2 77600 86397
0 9930 5 1 1 9929
0 9931 7 1 2 85938 9930
0 9932 5 1 1 9931
0 9933 7 1 2 86394 9932
0 9934 5 1 1 9933
0 9935 7 4 2 66650 86207
0 9936 5 2 1 86404
0 9937 7 1 2 79324 77714
0 9938 7 1 2 86405 9937
0 9939 5 1 1 9938
0 9940 7 1 2 9934 9939
0 9941 5 1 1 9940
0 9942 7 1 2 68614 9941
0 9943 5 1 1 9942
0 9944 7 6 2 65809 61447
0 9945 7 1 2 79431 86410
0 9946 5 1 1 9945
0 9947 7 1 2 81122 9946
0 9948 5 2 1 9947
0 9949 7 1 2 60255 86416
0 9950 5 1 1 9949
0 9951 7 8 2 65122 61656
0 9952 7 1 2 65810 75827
0 9953 5 1 1 9952
0 9954 7 1 2 79802 9953
0 9955 5 2 1 9954
0 9956 7 1 2 86418 86426
0 9957 5 1 1 9956
0 9958 7 1 2 9950 9957
0 9959 5 1 1 9958
0 9960 7 1 2 77686 86267
0 9961 7 1 2 9959 9960
0 9962 5 1 1 9961
0 9963 7 1 2 9943 9962
0 9964 5 1 1 9963
0 9965 7 1 2 63925 9964
0 9966 5 1 1 9965
0 9967 7 1 2 9925 9966
0 9968 5 1 1 9967
0 9969 7 1 2 62049 9968
0 9970 5 1 1 9969
0 9971 7 10 2 67020 68615
0 9972 7 1 2 63345 86428
0 9973 7 2 2 76118 9972
0 9974 7 1 2 66189 77071
0 9975 7 1 2 86438 9974
0 9976 5 1 1 9975
0 9977 7 1 2 61015 81594
0 9978 7 1 2 76685 85185
0 9979 7 1 2 9977 9978
0 9980 5 1 1 9979
0 9981 7 1 2 9976 9980
0 9982 5 1 1 9981
0 9983 7 1 2 79516 9982
0 9984 5 1 1 9983
0 9985 7 1 2 74349 79531
0 9986 7 1 2 86439 9985
0 9987 5 1 1 9986
0 9988 7 1 2 80622 83839
0 9989 7 1 2 84860 9988
0 9990 5 1 1 9989
0 9991 7 1 2 9987 9990
0 9992 7 1 2 9984 9991
0 9993 5 1 1 9992
0 9994 7 1 2 66651 9993
0 9995 5 1 1 9994
0 9996 7 3 2 71021 73730
0 9997 7 3 2 65811 79253
0 9998 7 1 2 86000 86443
0 9999 7 1 2 86440 9998
0 10000 5 1 1 9999
0 10001 7 1 2 9995 10000
0 10002 5 1 1 10001
0 10003 7 1 2 86152 10002
0 10004 5 1 1 10003
0 10005 7 1 2 9970 10004
0 10006 5 1 1 10005
0 10007 7 1 2 69783 10006
0 10008 5 1 1 10007
0 10009 7 2 2 68266 76119
0 10010 7 1 2 82193 86446
0 10011 5 1 1 10010
0 10012 7 3 2 64911 77703
0 10013 7 7 2 61657 67515
0 10014 7 2 2 63346 86451
0 10015 7 1 2 86448 86458
0 10016 5 1 1 10015
0 10017 7 1 2 10011 10016
0 10018 5 1 1 10017
0 10019 7 1 2 86153 10018
0 10020 5 1 1 10019
0 10021 7 4 2 81099 86075
0 10022 7 1 2 65974 86460
0 10023 7 1 2 77815 10022
0 10024 5 1 1 10023
0 10025 7 1 2 10020 10024
0 10026 5 1 1 10025
0 10027 7 1 2 64687 10026
0 10028 5 1 1 10027
0 10029 7 1 2 77821 86461
0 10030 5 1 1 10029
0 10031 7 1 2 10028 10030
0 10032 5 1 1 10031
0 10033 7 1 2 63672 10032
0 10034 5 1 1 10033
0 10035 7 16 2 68267 77540
0 10036 7 2 2 84283 86464
0 10037 7 4 2 61241 66806
0 10038 7 1 2 74091 76699
0 10039 7 1 2 86482 10038
0 10040 7 1 2 86480 10039
0 10041 5 1 1 10040
0 10042 7 1 2 10034 10041
0 10043 5 1 1 10042
0 10044 7 1 2 79517 10043
0 10045 5 1 1 10044
0 10046 7 1 2 80666 76082
0 10047 5 1 1 10046
0 10048 7 1 2 70030 86447
0 10049 5 1 1 10048
0 10050 7 1 2 10047 10049
0 10051 5 1 1 10050
0 10052 7 1 2 80189 86154
0 10053 7 1 2 10051 10052
0 10054 5 1 1 10053
0 10055 7 1 2 60256 77813
0 10056 5 1 1 10055
0 10057 7 1 2 61448 10056
0 10058 5 1 1 10057
0 10059 7 1 2 75707 74727
0 10060 5 2 1 10059
0 10061 7 1 2 10058 86486
0 10062 5 1 1 10061
0 10063 7 1 2 77854 86462
0 10064 7 1 2 10062 10063
0 10065 5 1 1 10064
0 10066 7 1 2 10054 10065
0 10067 5 1 1 10066
0 10068 7 1 2 84666 10067
0 10069 5 1 1 10068
0 10070 7 1 2 59826 72776
0 10071 5 3 1 10070
0 10072 7 6 2 63347 77541
0 10073 7 1 2 74815 86491
0 10074 7 1 2 86488 10073
0 10075 7 1 2 86395 10074
0 10076 5 1 1 10075
0 10077 7 1 2 67878 10076
0 10078 7 1 2 10069 10077
0 10079 7 1 2 10045 10078
0 10080 7 1 2 10008 10079
0 10081 5 1 1 10080
0 10082 7 1 2 9845 10081
0 10083 5 1 1 10082
0 10084 7 1 2 65352 10083
0 10085 5 1 1 10084
0 10086 7 2 2 63673 77456
0 10087 7 8 2 66190 61850
0 10088 7 1 2 72697 86499
0 10089 7 1 2 86497 10088
0 10090 5 1 1 10089
0 10091 7 1 2 82918 85695
0 10092 7 1 2 76893 10091
0 10093 5 1 1 10092
0 10094 7 1 2 10090 10093
0 10095 5 1 1 10094
0 10096 7 1 2 80190 10095
0 10097 5 1 1 10096
0 10098 7 1 2 80163 83948
0 10099 5 1 1 10098
0 10100 7 1 2 79339 79584
0 10101 5 1 1 10100
0 10102 7 1 2 10099 10101
0 10103 5 1 1 10102
0 10104 7 1 2 64912 10103
0 10105 5 1 1 10104
0 10106 7 1 2 62050 79337
0 10107 5 1 1 10106
0 10108 7 1 2 10105 10107
0 10109 5 1 1 10108
0 10110 7 1 2 71086 10109
0 10111 5 1 1 10110
0 10112 7 3 2 66652 79325
0 10113 7 7 2 62051 70743
0 10114 5 4 1 86510
0 10115 7 1 2 67879 86511
0 10116 5 1 1 10115
0 10117 7 1 2 77385 10116
0 10118 5 2 1 10117
0 10119 7 1 2 86507 86521
0 10120 5 1 1 10119
0 10121 7 1 2 10111 10120
0 10122 5 1 1 10121
0 10123 7 1 2 85186 10122
0 10124 5 1 1 10123
0 10125 7 1 2 79239 10124
0 10126 5 1 1 10125
0 10127 7 1 2 61851 10126
0 10128 5 1 1 10127
0 10129 7 1 2 10097 10128
0 10130 5 1 1 10129
0 10131 7 1 2 79727 10130
0 10132 5 1 1 10131
0 10133 7 1 2 82018 9837
0 10134 5 3 1 10133
0 10135 7 2 2 81282 85870
0 10136 7 6 2 68837 78737
0 10137 7 1 2 84655 86528
0 10138 7 1 2 86526 10137
0 10139 7 1 2 86523 10138
0 10140 5 1 1 10139
0 10141 7 1 2 10132 10140
0 10142 5 1 1 10141
0 10143 7 1 2 72545 10142
0 10144 5 1 1 10143
0 10145 7 5 2 61658 62888
0 10146 7 1 2 66191 4677
0 10147 5 1 1 10146
0 10148 7 1 2 71087 75086
0 10149 7 1 2 10147 10148
0 10150 5 1 1 10149
0 10151 7 1 2 8338 10150
0 10152 5 1 1 10151
0 10153 7 1 2 86534 10152
0 10154 5 1 1 10153
0 10155 7 5 2 80944 78124
0 10156 7 1 2 81673 84264
0 10157 7 1 2 86539 10156
0 10158 5 1 1 10157
0 10159 7 1 2 10154 10158
0 10160 5 1 1 10159
0 10161 7 1 2 65812 10160
0 10162 5 1 1 10161
0 10163 7 1 2 77731 85961
0 10164 5 1 1 10163
0 10165 7 5 2 64913 78547
0 10166 5 5 1 86544
0 10167 7 1 2 71088 81524
0 10168 7 1 2 86545 10167
0 10169 5 1 1 10168
0 10170 7 1 2 10164 10169
0 10171 5 1 1 10170
0 10172 7 1 2 61659 10171
0 10173 5 1 1 10172
0 10174 7 1 2 10162 10173
0 10175 5 1 1 10174
0 10176 7 1 2 85696 10175
0 10177 5 1 1 10176
0 10178 7 1 2 75917 85941
0 10179 5 1 1 10178
0 10180 7 1 2 77939 10179
0 10181 5 1 1 10180
0 10182 7 1 2 66192 10181
0 10183 5 1 1 10182
0 10184 7 1 2 85380 10183
0 10185 5 1 1 10184
0 10186 7 4 2 63674 85840
0 10187 5 1 1 86554
0 10188 7 1 2 72698 86555
0 10189 7 1 2 10185 10188
0 10190 5 1 1 10189
0 10191 7 1 2 10177 10190
0 10192 5 1 1 10191
0 10193 7 1 2 63926 10192
0 10194 5 1 1 10193
0 10195 7 1 2 77394 77020
0 10196 5 2 1 10195
0 10197 7 5 2 67021 77457
0 10198 5 2 1 86560
0 10199 7 1 2 77338 86561
0 10200 5 1 1 10199
0 10201 7 1 2 86558 10200
0 10202 5 1 1 10201
0 10203 7 2 2 64688 84298
0 10204 7 6 2 66807 63675
0 10205 7 3 2 80528 86569
0 10206 7 1 2 86567 86575
0 10207 7 1 2 10202 10206
0 10208 5 1 1 10207
0 10209 7 1 2 10194 10208
0 10210 5 1 1 10209
0 10211 7 1 2 79518 10210
0 10212 5 1 1 10211
0 10213 7 6 2 62052 63927
0 10214 7 3 2 61660 86578
0 10215 7 1 2 74846 86584
0 10216 7 1 2 77524 10215
0 10217 5 1 1 10216
0 10218 7 2 2 65123 61016
0 10219 7 1 2 79740 86587
0 10220 7 1 2 84962 10219
0 10221 5 1 1 10220
0 10222 7 1 2 10217 10221
0 10223 5 1 1 10222
0 10224 7 1 2 64689 10223
0 10225 5 1 1 10224
0 10226 7 1 2 75475 86585
0 10227 5 1 1 10226
0 10228 7 8 2 61017 68838
0 10229 7 1 2 70031 86589
0 10230 7 1 2 86054 10229
0 10231 5 1 1 10230
0 10232 7 1 2 10227 10231
0 10233 5 1 1 10232
0 10234 7 8 2 64224 70744
0 10235 5 2 1 86597
0 10236 7 1 2 75900 86598
0 10237 7 1 2 10233 10236
0 10238 5 1 1 10237
0 10239 7 1 2 10225 10238
0 10240 5 1 1 10239
0 10241 7 1 2 62540 10240
0 10242 5 1 1 10241
0 10243 7 6 2 67516 68839
0 10244 7 4 2 66653 86607
0 10245 5 1 1 86613
0 10246 7 1 2 82818 86614
0 10247 5 1 1 10246
0 10248 7 1 2 10242 10247
0 10249 5 1 1 10248
0 10250 7 1 2 68268 10249
0 10251 5 1 1 10250
0 10252 7 3 2 79741 80019
0 10253 7 1 2 71089 73759
0 10254 7 1 2 72816 10253
0 10255 7 1 2 86617 10254
0 10256 5 1 1 10255
0 10257 7 1 2 10251 10256
0 10258 5 1 1 10257
0 10259 7 1 2 67880 10258
0 10260 5 1 1 10259
0 10261 7 1 2 65691 81009
0 10262 7 1 2 77339 10261
0 10263 7 6 2 61661 75476
0 10264 5 2 1 86620
0 10265 7 2 2 64225 77458
0 10266 7 1 2 86621 86628
0 10267 7 1 2 10262 10266
0 10268 5 1 1 10267
0 10269 7 1 2 63676 10268
0 10270 7 1 2 10260 10269
0 10271 5 1 1 10270
0 10272 7 2 2 80191 81010
0 10273 7 1 2 67517 75930
0 10274 5 2 1 10273
0 10275 7 1 2 77368 86632
0 10276 5 1 1 10275
0 10277 7 3 2 75918 78281
0 10278 5 1 1 86634
0 10279 7 1 2 70745 86635
0 10280 5 1 1 10279
0 10281 7 1 2 10276 10280
0 10282 5 1 1 10281
0 10283 7 1 2 86630 10282
0 10284 5 1 1 10283
0 10285 7 3 2 63348 85814
0 10286 7 5 2 61449 78050
0 10287 7 1 2 78812 86640
0 10288 5 1 1 10287
0 10289 7 4 2 64226 75182
0 10290 5 1 1 86645
0 10291 7 1 2 79742 82130
0 10292 7 1 2 76858 10291
0 10293 7 1 2 86646 10292
0 10294 5 1 1 10293
0 10295 7 1 2 10288 10294
0 10296 5 1 1 10295
0 10297 7 1 2 86637 10296
0 10298 5 1 1 10297
0 10299 7 1 2 10284 10298
0 10300 5 1 1 10299
0 10301 7 1 2 65975 10300
0 10302 5 1 1 10301
0 10303 7 1 2 80192 86220
0 10304 7 1 2 85980 10303
0 10305 5 1 1 10304
0 10306 7 1 2 10302 10305
0 10307 5 1 1 10306
0 10308 7 1 2 64690 10307
0 10309 5 1 1 10308
0 10310 7 1 2 64914 77408
0 10311 5 1 1 10310
0 10312 7 1 2 85718 10311
0 10313 5 1 1 10312
0 10314 7 1 2 75919 86631
0 10315 7 1 2 10313 10314
0 10316 5 1 1 10315
0 10317 7 1 2 68616 10316
0 10318 7 1 2 10309 10317
0 10319 5 1 1 10318
0 10320 7 1 2 66808 10319
0 10321 7 1 2 10271 10320
0 10322 5 1 1 10321
0 10323 7 1 2 82819 84697
0 10324 5 1 1 10323
0 10325 7 1 2 81866 70943
0 10326 7 1 2 86052 10325
0 10327 5 1 1 10326
0 10328 7 1 2 78979 10327
0 10329 5 1 1 10328
0 10330 7 1 2 65124 10329
0 10331 5 1 1 10330
0 10332 7 11 2 63349 78247
0 10333 7 7 2 66413 67022
0 10334 5 1 1 86660
0 10335 7 3 2 61242 86661
0 10336 7 2 2 86649 86667
0 10337 5 1 1 86670
0 10338 7 1 2 10331 10337
0 10339 5 1 1 10338
0 10340 7 1 2 77156 10339
0 10341 5 1 1 10340
0 10342 7 8 2 61450 83091
0 10343 5 2 1 86672
0 10344 7 1 2 73740 86673
0 10345 5 1 1 10344
0 10346 7 2 2 68269 83949
0 10347 7 5 2 65813 66414
0 10348 7 1 2 82137 86684
0 10349 7 1 2 86682 10348
0 10350 5 1 1 10349
0 10351 7 1 2 10345 10350
0 10352 5 1 1 10351
0 10353 7 1 2 77180 10352
0 10354 5 1 1 10353
0 10355 7 1 2 72699 76218
0 10356 7 5 2 66415 83734
0 10357 5 3 1 86689
0 10358 7 1 2 77533 86690
0 10359 7 1 2 10355 10358
0 10360 5 1 1 10359
0 10361 7 1 2 10354 10360
0 10362 7 1 2 10341 10361
0 10363 5 1 1 10362
0 10364 7 1 2 66654 10363
0 10365 5 1 1 10364
0 10366 7 1 2 10324 10365
0 10367 5 1 1 10366
0 10368 7 1 2 86369 10367
0 10369 5 1 1 10368
0 10370 7 1 2 60447 10369
0 10371 7 1 2 10322 10370
0 10372 7 1 2 10212 10371
0 10373 7 1 2 10144 10372
0 10374 5 1 1 10373
0 10375 7 1 2 65539 10374
0 10376 7 1 2 10085 10375
0 10377 5 1 1 10376
0 10378 7 1 2 9645 10377
0 10379 5 1 1 10378
0 10380 7 1 2 74006 10379
0 10381 5 1 1 10380
0 10382 7 37 2 65540 66809
0 10383 5 9 1 86697
0 10384 7 26 2 60649 61852
0 10385 5 5 1 86743
0 10386 7 49 2 86734 86769
0 10387 5 3 1 86774
0 10388 7 15 2 62889 75542
0 10389 5 4 1 86826
0 10390 7 2 2 68270 86827
0 10391 7 1 2 75080 86845
0 10392 5 1 1 10391
0 10393 7 6 2 65814 63350
0 10394 7 1 2 81046 86847
0 10395 7 1 2 83950 10394
0 10396 5 1 1 10395
0 10397 7 1 2 10392 10396
0 10398 5 1 1 10397
0 10399 7 1 2 80398 10398
0 10400 5 1 1 10399
0 10401 7 2 2 65125 82105
0 10402 7 7 2 62053 75679
0 10403 7 1 2 85465 86855
0 10404 7 1 2 86853 10403
0 10405 5 1 1 10404
0 10406 7 1 2 10400 10405
0 10407 5 1 1 10406
0 10408 7 1 2 62250 10407
0 10409 5 1 1 10408
0 10410 7 4 2 67518 83735
0 10411 7 5 2 66655 74674
0 10412 7 1 2 74274 84632
0 10413 7 1 2 86866 10412
0 10414 7 1 2 86862 10413
0 10415 5 1 1 10414
0 10416 7 1 2 10409 10415
0 10417 5 1 1 10416
0 10418 7 1 2 64440 10417
0 10419 5 1 1 10418
0 10420 7 2 2 63351 80399
0 10421 7 6 2 67881 71353
0 10422 7 1 2 72764 74338
0 10423 7 1 2 86873 10422
0 10424 7 1 2 86871 10423
0 10425 5 1 1 10424
0 10426 7 1 2 10419 10425
0 10427 5 1 1 10426
0 10428 7 1 2 64227 10427
0 10429 5 1 1 10428
0 10430 7 3 2 65126 81076
0 10431 7 3 2 62890 79254
0 10432 5 2 1 86882
0 10433 7 1 2 62054 86883
0 10434 7 1 2 86879 10433
0 10435 5 1 1 10434
0 10436 7 1 2 75148 86487
0 10437 5 1 1 10436
0 10438 7 1 2 84025 10437
0 10439 5 1 1 10438
0 10440 7 4 2 62055 78183
0 10441 5 2 1 86887
0 10442 7 1 2 74361 86888
0 10443 5 1 1 10442
0 10444 7 1 2 10439 10443
0 10445 5 1 1 10444
0 10446 7 1 2 81154 10445
0 10447 5 1 1 10446
0 10448 7 1 2 10435 10447
0 10449 5 1 1 10448
0 10450 7 1 2 63352 10449
0 10451 5 1 1 10450
0 10452 7 3 2 79432 84824
0 10453 7 1 2 71967 81386
0 10454 7 1 2 86893 10453
0 10455 5 1 1 10454
0 10456 7 1 2 10451 10455
0 10457 5 1 1 10456
0 10458 7 1 2 62251 10457
0 10459 5 1 1 10458
0 10460 7 1 2 10429 10459
0 10461 5 1 1 10460
0 10462 7 1 2 65692 10461
0 10463 5 1 1 10462
0 10464 7 5 2 64228 71968
0 10465 5 4 1 86896
0 10466 7 1 2 67519 86901
0 10467 5 1 1 10466
0 10468 7 1 2 85648 10467
0 10469 5 1 1 10468
0 10470 7 1 2 85630 10469
0 10471 5 1 1 10470
0 10472 7 1 2 66193 10471
0 10473 5 1 1 10472
0 10474 7 1 2 73908 82396
0 10475 7 1 2 83834 10474
0 10476 5 1 1 10475
0 10477 7 10 2 64441 66194
0 10478 5 3 1 86905
0 10479 7 2 2 78184 86906
0 10480 5 1 1 86918
0 10481 7 1 2 64229 86919
0 10482 5 1 1 10481
0 10483 7 1 2 85560 10482
0 10484 5 1 1 10483
0 10485 7 1 2 61451 76432
0 10486 7 1 2 10484 10485
0 10487 5 1 1 10486
0 10488 7 1 2 10476 10487
0 10489 5 1 1 10488
0 10490 7 1 2 65815 10489
0 10491 5 1 1 10490
0 10492 7 4 2 61452 77459
0 10493 5 1 1 86920
0 10494 7 1 2 78801 86921
0 10495 5 1 1 10494
0 10496 7 1 2 10491 10495
0 10497 5 1 1 10496
0 10498 7 1 2 63353 10497
0 10499 5 1 1 10498
0 10500 7 1 2 77601 82431
0 10501 5 1 1 10500
0 10502 7 1 2 10499 10501
0 10503 5 1 1 10502
0 10504 7 1 2 81155 10503
0 10505 5 1 1 10504
0 10506 7 1 2 10473 10505
0 10507 7 1 2 10463 10506
0 10508 5 1 1 10507
0 10509 7 1 2 64915 10508
0 10510 5 1 1 10509
0 10511 7 1 2 65127 86671
0 10512 5 1 1 10511
0 10513 7 2 2 79763 78016
0 10514 7 1 2 82106 86924
0 10515 5 1 1 10514
0 10516 7 1 2 74092 83168
0 10517 5 1 1 10516
0 10518 7 1 2 10515 10517
0 10519 5 1 1 10518
0 10520 7 1 2 77229 10519
0 10521 5 1 1 10520
0 10522 7 3 2 75183 74219
0 10523 5 2 1 86926
0 10524 7 1 2 77340 86927
0 10525 5 1 1 10524
0 10526 7 1 2 10521 10525
0 10527 5 1 1 10526
0 10528 7 1 2 62891 82302
0 10529 7 1 2 10527 10528
0 10530 5 1 1 10529
0 10531 7 1 2 10512 10530
0 10532 5 1 1 10531
0 10533 7 1 2 81156 10532
0 10534 5 1 1 10533
0 10535 7 1 2 77230 74093
0 10536 5 1 1 10535
0 10537 7 1 2 4434 10536
0 10538 5 1 1 10537
0 10539 7 8 2 64230 62892
0 10540 5 2 1 86931
0 10541 7 1 2 80725 86932
0 10542 7 1 2 10538 10541
0 10543 5 1 1 10542
0 10544 7 1 2 6190 10543
0 10545 5 1 1 10544
0 10546 7 1 2 84231 10545
0 10547 5 1 1 10546
0 10548 7 2 2 84878 85036
0 10549 7 1 2 80559 86361
0 10550 7 1 2 70970 10549
0 10551 7 1 2 86941 10550
0 10552 5 1 1 10551
0 10553 7 1 2 78214 84463
0 10554 5 2 1 10553
0 10555 7 1 2 68271 86943
0 10556 7 1 2 84243 10555
0 10557 5 1 1 10556
0 10558 7 1 2 10552 10557
0 10559 5 1 1 10558
0 10560 7 1 2 70746 10559
0 10561 5 1 1 10560
0 10562 7 1 2 10547 10561
0 10563 7 1 2 10534 10562
0 10564 7 1 2 10510 10563
0 10565 5 1 1 10564
0 10566 7 1 2 86775 10565
0 10567 5 1 1 10566
0 10568 7 1 2 70747 86944
0 10569 5 1 1 10568
0 10570 7 5 2 65816 77231
0 10571 5 2 1 86945
0 10572 7 2 2 62252 86946
0 10573 5 1 1 86952
0 10574 7 1 2 61243 10573
0 10575 5 1 1 10574
0 10576 7 1 2 79569 10575
0 10577 5 1 1 10576
0 10578 7 1 2 10569 10577
0 10579 5 1 1 10578
0 10580 7 1 2 60257 10579
0 10581 5 1 1 10580
0 10582 7 2 2 60258 77667
0 10583 7 3 2 62056 85815
0 10584 5 2 1 86956
0 10585 7 1 2 86954 86957
0 10586 5 1 1 10585
0 10587 7 1 2 74261 78693
0 10588 5 1 1 10587
0 10589 7 1 2 73662 72765
0 10590 7 1 2 79570 10589
0 10591 5 1 1 10590
0 10592 7 1 2 10588 10591
0 10593 5 1 1 10592
0 10594 7 1 2 67520 77232
0 10595 7 1 2 10593 10594
0 10596 5 1 1 10595
0 10597 7 1 2 10586 10596
0 10598 5 1 1 10597
0 10599 7 1 2 64231 10598
0 10600 5 1 1 10599
0 10601 7 1 2 10581 10600
0 10602 5 1 1 10601
0 10603 7 1 2 68272 10602
0 10604 5 1 1 10603
0 10605 7 7 2 60259 67521
0 10606 7 1 2 75432 82919
0 10607 7 1 2 86961 10606
0 10608 5 1 1 10607
0 10609 7 1 2 10604 10608
0 10610 5 1 1 10609
0 10611 7 13 2 61662 66810
0 10612 7 6 2 60448 86968
0 10613 5 5 1 86981
0 10614 7 9 2 65541 61453
0 10615 7 4 2 86982 86992
0 10616 5 1 1 87001
0 10617 7 1 2 10610 87002
0 10618 5 1 1 10617
0 10619 7 1 2 62893 69451
0 10620 5 1 1 10619
0 10621 7 2 2 70478 82131
0 10622 5 3 1 87005
0 10623 7 1 2 67882 87007
0 10624 5 2 1 10623
0 10625 7 1 2 87010 86897
0 10626 5 1 1 10625
0 10627 7 1 2 10620 10626
0 10628 5 1 1 10627
0 10629 7 1 2 66195 10628
0 10630 5 1 1 10629
0 10631 7 1 2 74464 77460
0 10632 5 1 1 10631
0 10633 7 1 2 10630 10632
0 10634 5 1 1 10633
0 10635 7 1 2 64916 10634
0 10636 5 1 1 10635
0 10637 7 2 2 76627 78548
0 10638 5 1 1 87012
0 10639 7 1 2 80476 87013
0 10640 5 1 1 10639
0 10641 7 1 2 10636 10640
0 10642 5 1 1 10641
0 10643 7 9 2 60650 66416
0 10644 7 1 2 81765 87014
0 10645 7 1 2 86406 10644
0 10646 7 1 2 10642 10645
0 10647 5 1 1 10646
0 10648 7 1 2 10618 10647
0 10649 7 1 2 10567 10648
0 10650 5 1 1 10649
0 10651 7 1 2 63928 10650
0 10652 5 1 1 10651
0 10653 7 10 2 62541 70748
0 10654 7 5 2 61454 61853
0 10655 7 1 2 81088 87033
0 10656 7 1 2 87023 10655
0 10657 5 2 1 10656
0 10658 7 2 2 84008 86608
0 10659 7 1 2 66811 76715
0 10660 7 1 2 87040 10659
0 10661 5 1 1 10660
0 10662 7 1 2 87038 10661
0 10663 5 1 1 10662
0 10664 7 1 2 66656 10663
0 10665 5 1 1 10664
0 10666 7 5 2 62542 63929
0 10667 7 1 2 86500 87042
0 10668 5 3 1 10667
0 10669 7 3 2 61854 87043
0 10670 5 2 1 87050
0 10671 7 3 2 66812 86609
0 10672 7 1 2 66196 76716
0 10673 7 1 2 87055 10672
0 10674 5 1 1 10673
0 10675 7 1 2 87053 10674
0 10676 5 1 1 10675
0 10677 7 1 2 64917 10676
0 10678 5 1 1 10677
0 10679 7 1 2 87047 10678
0 10680 5 1 1 10679
0 10681 7 1 2 79340 10680
0 10682 5 1 1 10681
0 10683 7 1 2 65353 10682
0 10684 7 1 2 10665 10683
0 10685 5 1 1 10684
0 10686 7 2 2 70749 87044
0 10687 7 1 2 86250 87058
0 10688 5 1 1 10687
0 10689 7 2 2 60449 10688
0 10690 7 1 2 80651 80993
0 10691 7 1 2 86854 10690
0 10692 7 1 2 87056 10691
0 10693 5 1 1 10692
0 10694 7 1 2 87060 10693
0 10695 5 1 1 10694
0 10696 7 1 2 70305 10695
0 10697 7 1 2 10685 10696
0 10698 5 1 1 10697
0 10699 7 1 2 65693 86310
0 10700 7 1 2 87041 10699
0 10701 5 1 1 10700
0 10702 7 1 2 87039 10701
0 10703 5 1 1 10702
0 10704 7 1 2 66657 10703
0 10705 5 1 1 10704
0 10706 7 2 2 81632 86610
0 10707 7 1 2 86311 87062
0 10708 5 1 1 10707
0 10709 7 1 2 87054 10708
0 10710 5 1 1 10709
0 10711 7 1 2 64918 10710
0 10712 5 1 1 10711
0 10713 7 1 2 10712 87048
0 10714 5 1 1 10713
0 10715 7 1 2 79341 10714
0 10716 5 1 1 10715
0 10717 7 1 2 65354 10716
0 10718 7 1 2 10705 10717
0 10719 5 1 1 10718
0 10720 7 18 2 66658 66813
0 10721 7 2 2 71022 87064
0 10722 7 1 2 75411 87063
0 10723 7 1 2 87082 10722
0 10724 5 1 1 10723
0 10725 7 1 2 87061 10724
0 10726 5 1 1 10725
0 10727 7 1 2 65817 10726
0 10728 7 1 2 10719 10727
0 10729 5 1 1 10728
0 10730 7 3 2 65128 80400
0 10731 5 1 1 87084
0 10732 7 1 2 85667 87085
0 10733 5 1 1 10732
0 10734 7 3 2 61855 79608
0 10735 5 3 1 87087
0 10736 7 7 2 66814 80841
0 10737 5 2 1 87093
0 10738 7 1 2 87090 87100
0 10739 5 7 1 10738
0 10740 7 2 2 61455 87102
0 10741 5 1 1 87109
0 10742 7 1 2 60260 87110
0 10743 5 1 1 10742
0 10744 7 1 2 10733 10743
0 10745 5 1 1 10744
0 10746 7 1 2 64232 87059
0 10747 7 1 2 10745 10746
0 10748 5 1 1 10747
0 10749 7 1 2 10729 10748
0 10750 7 1 2 10698 10749
0 10751 5 1 1 10750
0 10752 7 1 2 65542 10751
0 10753 5 1 1 10752
0 10754 7 21 2 60651 66815
0 10755 5 4 1 87111
0 10756 7 9 2 63930 87112
0 10757 5 1 1 87136
0 10758 7 1 2 72875 87024
0 10759 7 1 2 87137 10758
0 10760 7 1 2 84244 10759
0 10761 5 1 1 10760
0 10762 7 1 2 10753 10761
0 10763 5 1 1 10762
0 10764 7 1 2 68273 10763
0 10765 5 1 1 10764
0 10766 7 1 2 70750 80826
0 10767 7 8 2 65543 61856
0 10768 5 1 1 87145
0 10769 7 4 2 87132 10768
0 10770 5 44 1 87153
0 10771 7 2 2 62543 87157
0 10772 7 1 2 86872 87201
0 10773 7 1 2 10766 10772
0 10774 5 1 1 10773
0 10775 7 1 2 10765 10774
0 10776 5 1 1 10775
0 10777 7 1 2 67883 10776
0 10778 5 1 1 10777
0 10779 7 15 2 60450 66816
0 10780 7 2 2 65544 87203
0 10781 7 2 2 86622 87218
0 10782 5 5 1 87220
0 10783 7 2 2 61456 79126
0 10784 5 5 1 87227
0 10785 7 13 2 71533 87229
0 10786 5 4 1 87234
0 10787 7 1 2 80401 87235
0 10788 5 2 1 10787
0 10789 7 1 2 84237 87251
0 10790 5 1 1 10789
0 10791 7 1 2 86776 10790
0 10792 5 1 1 10791
0 10793 7 1 2 87222 10792
0 10794 5 1 1 10793
0 10795 7 2 2 81011 78185
0 10796 7 2 2 65818 72649
0 10797 5 1 1 87255
0 10798 7 1 2 64233 87256
0 10799 7 1 2 87253 10798
0 10800 7 1 2 10794 10799
0 10801 5 1 1 10800
0 10802 7 1 2 10778 10801
0 10803 5 1 1 10802
0 10804 7 1 2 74007 10803
0 10805 5 1 1 10804
0 10806 7 10 2 62894 68840
0 10807 7 6 2 66817 87257
0 10808 7 1 2 73663 87267
0 10809 5 1 1 10808
0 10810 7 8 2 67884 86076
0 10811 7 1 2 62253 87273
0 10812 5 1 1 10811
0 10813 7 1 2 10809 10812
0 10814 5 1 1 10813
0 10815 7 1 2 73374 10814
0 10816 5 1 1 10815
0 10817 7 1 2 70751 87274
0 10818 5 1 1 10817
0 10819 7 1 2 10816 10818
0 10820 5 1 1 10819
0 10821 7 1 2 65819 10820
0 10822 5 1 1 10821
0 10823 7 1 2 86077 86522
0 10824 5 1 1 10823
0 10825 7 1 2 10822 10824
0 10826 5 1 1 10825
0 10827 7 1 2 62544 10826
0 10828 5 1 1 10827
0 10829 7 1 2 65820 79832
0 10830 5 2 1 10829
0 10831 7 1 2 73129 87281
0 10832 5 1 1 10831
0 10833 7 1 2 65694 10832
0 10834 5 1 1 10833
0 10835 7 2 2 76357 73093
0 10836 5 2 1 87283
0 10837 7 1 2 10834 87285
0 10838 5 1 1 10837
0 10839 7 1 2 66197 10838
0 10840 5 1 1 10839
0 10841 7 1 2 60086 10840
0 10842 5 1 1 10841
0 10843 7 11 2 61857 67885
0 10844 7 8 2 63931 87287
0 10845 7 3 2 64442 70479
0 10846 5 1 1 87306
0 10847 7 1 2 61244 10846
0 10848 5 1 1 10847
0 10849 7 1 2 87298 10848
0 10850 7 1 2 10842 10849
0 10851 5 1 1 10850
0 10852 7 12 2 62895 63932
0 10853 7 3 2 61858 87309
0 10854 5 1 1 87321
0 10855 7 4 2 65821 70443
0 10856 5 1 1 87324
0 10857 7 3 2 69445 10856
0 10858 5 1 1 87328
0 10859 7 9 2 67886 68841
0 10860 7 6 2 66818 87331
0 10861 5 3 1 87340
0 10862 7 1 2 70032 87341
0 10863 7 1 2 10858 10862
0 10864 5 1 1 10863
0 10865 7 1 2 10854 10864
0 10866 5 1 1 10865
0 10867 7 1 2 70590 87329
0 10868 5 1 1 10867
0 10869 7 1 2 67522 10868
0 10870 7 1 2 10866 10869
0 10871 5 1 1 10870
0 10872 7 1 2 10851 10871
0 10873 7 1 2 10828 10872
0 10874 5 1 1 10873
0 10875 7 1 2 65545 10874
0 10876 5 1 1 10875
0 10877 7 2 2 76628 78965
0 10878 7 1 2 65695 87349
0 10879 5 1 1 10878
0 10880 7 1 2 78204 10879
0 10881 5 1 1 10880
0 10882 7 1 2 64234 10881
0 10883 5 1 1 10882
0 10884 7 1 2 85227 10883
0 10885 5 1 1 10884
0 10886 7 1 2 65822 10885
0 10887 5 1 1 10886
0 10888 7 1 2 61245 4840
0 10889 5 1 1 10888
0 10890 7 1 2 70306 78867
0 10891 7 1 2 10889 10890
0 10892 5 1 1 10891
0 10893 7 1 2 10887 10892
0 10894 5 1 1 10893
0 10895 7 1 2 64443 10894
0 10896 5 1 1 10895
0 10897 7 1 2 62254 78186
0 10898 5 3 1 10897
0 10899 7 6 2 64235 67887
0 10900 7 2 2 66198 87354
0 10901 7 1 2 65823 87360
0 10902 5 1 1 10901
0 10903 7 1 2 87351 10902
0 10904 5 1 1 10903
0 10905 7 1 2 65696 10904
0 10906 5 1 1 10905
0 10907 7 1 2 67888 87025
0 10908 5 2 1 10907
0 10909 7 1 2 10906 87362
0 10910 5 1 1 10909
0 10911 7 1 2 62057 10910
0 10912 5 1 1 10911
0 10913 7 7 2 78269 77495
0 10914 7 1 2 70752 78294
0 10915 7 1 2 87364 10914
0 10916 5 1 1 10915
0 10917 7 5 2 62896 76128
0 10918 5 1 1 87371
0 10919 7 2 2 64919 77395
0 10920 5 4 1 87376
0 10921 7 1 2 10918 87378
0 10922 7 1 2 10916 10921
0 10923 7 1 2 10912 10922
0 10924 7 1 2 10896 10923
0 10925 5 1 1 10924
0 10926 7 1 2 87138 10925
0 10927 5 1 1 10926
0 10928 7 1 2 10876 10927
0 10929 5 1 1 10928
0 10930 7 1 2 63354 10929
0 10931 5 1 1 10930
0 10932 7 22 2 63933 87158
0 10933 7 1 2 64236 82469
0 10934 5 1 1 10933
0 10935 7 1 2 76660 10934
0 10936 5 1 1 10935
0 10937 7 1 2 87382 10936
0 10938 5 1 1 10937
0 10939 7 4 2 62255 70444
0 10940 5 1 1 87404
0 10941 7 3 2 65546 75901
0 10942 7 1 2 86319 87408
0 10943 7 1 2 87405 10942
0 10944 5 1 1 10943
0 10945 7 1 2 10938 10944
0 10946 5 1 1 10945
0 10947 7 2 2 70033 77766
0 10948 5 1 1 87411
0 10949 7 1 2 10946 87412
0 10950 5 1 1 10949
0 10951 7 1 2 85965 87307
0 10952 5 1 1 10951
0 10953 7 1 2 85727 10952
0 10954 5 1 1 10953
0 10955 7 1 2 64920 10954
0 10956 5 1 1 10955
0 10957 7 1 2 69152 85394
0 10958 5 1 1 10957
0 10959 7 1 2 10956 10958
0 10960 5 1 1 10959
0 10961 7 1 2 87383 10960
0 10962 5 1 1 10961
0 10963 7 4 2 64444 65547
0 10964 7 1 2 67023 77341
0 10965 7 1 2 87413 10964
0 10966 7 5 2 66819 80529
0 10967 7 18 2 62897 76629
0 10968 5 1 1 87422
0 10969 7 1 2 87417 87423
0 10970 7 1 2 10965 10969
0 10971 5 1 1 10970
0 10972 7 1 2 10962 10971
0 10973 5 1 1 10972
0 10974 7 1 2 69632 10973
0 10975 5 1 1 10974
0 10976 7 1 2 10950 10975
0 10977 7 1 2 10931 10976
0 10978 5 1 1 10977
0 10979 7 1 2 80402 10978
0 10980 5 1 1 10979
0 10981 7 1 2 74220 78868
0 10982 7 2 2 87057 10981
0 10983 7 6 2 64445 65355
0 10984 7 1 2 65548 69633
0 10985 7 1 2 87442 10984
0 10986 7 1 2 82194 10985
0 10987 7 1 2 87440 10986
0 10988 5 1 1 10987
0 10989 7 1 2 10980 10988
0 10990 5 1 1 10989
0 10991 7 1 2 79519 10990
0 10992 5 1 1 10991
0 10993 7 3 2 75680 87258
0 10994 7 2 2 78802 86238
0 10995 7 1 2 87448 87451
0 10996 5 1 1 10995
0 10997 7 4 2 65129 86078
0 10998 7 1 2 86691 87453
0 10999 5 1 1 10998
0 11000 7 1 2 10996 10999
0 11001 5 1 1 11000
0 11002 7 1 2 64237 11001
0 11003 5 1 1 11002
0 11004 7 1 2 78549 86322
0 11005 7 1 2 80827 11004
0 11006 5 1 1 11005
0 11007 7 1 2 11003 11006
0 11008 5 1 1 11007
0 11009 7 1 2 64921 11008
0 11010 5 1 1 11009
0 11011 7 1 2 68274 87454
0 11012 7 8 2 64238 66199
0 11013 5 1 1 87457
0 11014 7 1 2 67889 11013
0 11015 5 4 1 11014
0 11016 7 3 2 66417 78587
0 11017 5 1 1 87469
0 11018 7 1 2 87465 87470
0 11019 7 1 2 11011 11018
0 11020 5 1 1 11019
0 11021 7 1 2 11010 11020
0 11022 5 1 1 11021
0 11023 7 1 2 65824 11022
0 11024 5 1 1 11023
0 11025 7 5 2 67890 80530
0 11026 7 1 2 86346 86390
0 11027 7 1 2 87472 11026
0 11028 5 1 1 11027
0 11029 7 1 2 11024 11028
0 11030 5 1 1 11029
0 11031 7 1 2 65549 11030
0 11032 5 1 1 11031
0 11033 7 2 2 67891 86605
0 11034 5 5 1 87477
0 11035 7 1 2 87471 87479
0 11036 5 1 1 11035
0 11037 7 1 2 74362 85060
0 11038 5 1 1 11037
0 11039 7 1 2 65130 11038
0 11040 7 1 2 11036 11039
0 11041 5 1 1 11040
0 11042 7 4 2 70034 79479
0 11043 5 1 1 87484
0 11044 7 1 2 60261 11043
0 11045 5 1 1 11044
0 11046 7 2 2 86349 87113
0 11047 7 1 2 68275 87488
0 11048 7 1 2 11045 11047
0 11049 7 1 2 11041 11048
0 11050 5 1 1 11049
0 11051 7 1 2 11032 11050
0 11052 5 1 1 11051
0 11053 7 1 2 62256 11052
0 11054 5 1 1 11053
0 11055 7 2 2 82027 84919
0 11056 5 1 1 87490
0 11057 7 1 2 87384 87491
0 11058 5 1 1 11057
0 11059 7 1 2 11054 11058
0 11060 5 1 1 11059
0 11061 7 1 2 81157 11060
0 11062 5 1 1 11061
0 11063 7 4 2 79644 87159
0 11064 5 1 1 87492
0 11065 7 1 2 86987 86823
0 11066 5 2 1 11065
0 11067 7 12 2 11064 87496
0 11068 7 9 2 60262 74675
0 11069 5 1 1 87510
0 11070 7 2 2 81525 87511
0 11071 7 1 2 87310 87519
0 11072 5 2 1 11071
0 11073 7 9 2 65131 79554
0 11074 5 1 1 87523
0 11075 7 1 2 87524 87449
0 11076 5 1 1 11075
0 11077 7 2 2 75477 82624
0 11078 5 2 1 87532
0 11079 7 1 2 11076 87534
0 11080 5 1 1 11079
0 11081 7 1 2 64922 11080
0 11082 5 1 1 11081
0 11083 7 3 2 63934 83736
0 11084 7 1 2 83615 87536
0 11085 5 1 1 11084
0 11086 7 1 2 11082 11085
0 11087 5 1 1 11086
0 11088 7 1 2 64239 11087
0 11089 5 1 1 11088
0 11090 7 1 2 81961 82831
0 11091 5 1 1 11090
0 11092 7 1 2 11089 11091
0 11093 5 1 1 11092
0 11094 7 1 2 69061 11093
0 11095 5 1 1 11094
0 11096 7 1 2 87521 11095
0 11097 5 1 1 11096
0 11098 7 1 2 87498 11097
0 11099 5 1 1 11098
0 11100 7 4 2 65356 66820
0 11101 7 1 2 86993 87539
0 11102 7 1 2 81346 11101
0 11103 7 2 2 67523 85364
0 11104 7 1 2 87473 87543
0 11105 7 1 2 11102 11104
0 11106 5 1 1 11105
0 11107 7 1 2 11099 11106
0 11108 7 1 2 11062 11107
0 11109 5 1 1 11108
0 11110 7 1 2 82785 11109
0 11111 5 1 1 11110
0 11112 7 1 2 75184 77421
0 11113 5 1 1 11112
0 11114 7 2 2 67524 85657
0 11115 5 1 1 87545
0 11116 7 1 2 74275 83465
0 11117 7 1 2 87546 11116
0 11118 5 1 1 11117
0 11119 7 1 2 11113 11118
0 11120 5 1 1 11119
0 11121 7 1 2 68276 11120
0 11122 5 1 1 11121
0 11123 7 5 2 62545 73345
0 11124 5 3 1 87547
0 11125 7 1 2 83895 87548
0 11126 5 1 1 11125
0 11127 7 1 2 9593 11126
0 11128 5 1 1 11127
0 11129 7 1 2 85023 11128
0 11130 5 1 1 11129
0 11131 7 1 2 11122 11130
0 11132 5 1 1 11131
0 11133 7 1 2 64923 11132
0 11134 5 1 1 11133
0 11135 7 4 2 64446 82367
0 11136 5 2 1 87555
0 11137 7 2 2 81136 84734
0 11138 5 1 1 87561
0 11139 7 1 2 60263 87562
0 11140 5 1 1 11139
0 11141 7 3 2 66418 71354
0 11142 5 2 1 87563
0 11143 7 1 2 75061 87564
0 11144 5 1 1 11143
0 11145 7 1 2 11140 11144
0 11146 5 1 1 11145
0 11147 7 1 2 87556 11146
0 11148 5 1 1 11147
0 11149 7 1 2 85767 87525
0 11150 5 1 1 11149
0 11151 7 1 2 11148 11150
0 11152 7 1 2 11134 11151
0 11153 5 1 1 11152
0 11154 7 1 2 65825 11153
0 11155 5 1 1 11154
0 11156 7 2 2 80726 82368
0 11157 5 2 1 87568
0 11158 7 1 2 64447 82023
0 11159 7 1 2 87569 11158
0 11160 5 1 1 11159
0 11161 7 1 2 11155 11160
0 11162 5 1 1 11161
0 11163 7 1 2 87385 11162
0 11164 5 1 1 11163
0 11165 7 8 2 70035 75185
0 11166 5 2 1 87572
0 11167 7 1 2 87414 87573
0 11168 7 1 2 87441 11167
0 11169 5 1 1 11168
0 11170 7 1 2 11164 11169
0 11171 5 1 1 11170
0 11172 7 1 2 81158 11171
0 11173 5 1 1 11172
0 11174 7 2 2 65550 81489
0 11175 5 1 1 87582
0 11176 7 5 2 64448 60451
0 11177 7 6 2 60264 66821
0 11178 7 1 2 87584 87589
0 11179 7 1 2 87583 11178
0 11180 5 1 1 11179
0 11181 7 4 2 65357 80164
0 11182 5 3 1 87595
0 11183 7 5 2 64449 60265
0 11184 5 1 1 87602
0 11185 7 1 2 87160 87603
0 11186 7 1 2 87596 11185
0 11187 5 1 1 11186
0 11188 7 1 2 11180 11187
0 11189 5 1 1 11188
0 11190 7 1 2 85637 11189
0 11191 5 1 1 11190
0 11192 7 7 2 62058 78694
0 11193 5 3 1 87607
0 11194 7 2 2 79399 85440
0 11195 5 1 1 87617
0 11196 7 1 2 81100 87618
0 11197 7 1 2 87608 11196
0 11198 5 1 1 11197
0 11199 7 1 2 85631 11198
0 11200 5 1 1 11199
0 11201 7 1 2 87161 11200
0 11202 5 1 1 11201
0 11203 7 1 2 83737 87221
0 11204 5 1 1 11203
0 11205 7 7 2 60652 63355
0 11206 7 1 2 79480 85826
0 11207 7 1 2 87619 11206
0 11208 7 1 2 85810 11207
0 11209 5 1 1 11208
0 11210 7 1 2 11204 11209
0 11211 7 1 2 11202 11210
0 11212 5 1 1 11211
0 11213 7 1 2 87026 11212
0 11214 5 1 1 11213
0 11215 7 1 2 11191 11214
0 11216 5 1 1 11215
0 11217 7 1 2 65826 11216
0 11218 5 1 1 11217
0 11219 7 7 2 65551 61663
0 11220 5 2 1 87626
0 11221 7 10 2 87204 87627
0 11222 5 2 1 87635
0 11223 7 1 2 73346 87512
0 11224 7 1 2 87636 11223
0 11225 5 1 1 11224
0 11226 7 1 2 81283 87604
0 11227 7 1 2 85587 11226
0 11228 7 1 2 87162 11227
0 11229 5 1 1 11228
0 11230 7 1 2 11225 11229
0 11231 5 1 1 11230
0 11232 7 1 2 62257 77767
0 11233 7 1 2 11231 11232
0 11234 5 1 1 11233
0 11235 7 1 2 11218 11234
0 11236 5 1 1 11235
0 11237 7 1 2 63935 11236
0 11238 5 1 1 11237
0 11239 7 1 2 78803 80749
0 11240 7 1 2 84946 11239
0 11241 7 4 2 79609 86698
0 11242 7 2 2 80945 87332
0 11243 7 1 2 87647 87651
0 11244 7 1 2 11240 11243
0 11245 5 1 1 11244
0 11246 7 1 2 11238 11245
0 11247 7 1 2 11173 11246
0 11248 5 1 1 11247
0 11249 7 1 2 69634 11248
0 11250 5 1 1 11249
0 11251 7 1 2 67248 79837
0 11252 5 2 1 11251
0 11253 7 6 2 66419 71023
0 11254 7 1 2 87450 87655
0 11255 5 1 1 11254
0 11256 7 1 2 87535 11255
0 11257 5 1 1 11256
0 11258 7 1 2 75902 86907
0 11259 7 1 2 11257 11258
0 11260 5 1 1 11259
0 11261 7 1 2 87522 11260
0 11262 5 1 1 11261
0 11263 7 1 2 87499 11262
0 11264 5 1 1 11263
0 11265 7 10 2 66822 62898
0 11266 7 1 2 87605 87661
0 11267 7 1 2 82039 11266
0 11268 7 1 2 84933 87409
0 11269 7 1 2 11267 11268
0 11270 5 1 1 11269
0 11271 7 2 2 64924 79764
0 11272 5 1 1 87671
0 11273 7 3 2 64450 75828
0 11274 5 2 1 87673
0 11275 7 1 2 70753 87674
0 11276 5 1 1 11275
0 11277 7 1 2 11272 11276
0 11278 5 1 1 11277
0 11279 7 2 2 67892 75903
0 11280 7 1 2 11278 87678
0 11281 5 1 1 11280
0 11282 7 4 2 66420 81526
0 11283 5 2 1 87680
0 11284 7 1 2 77369 87681
0 11285 5 1 1 11284
0 11286 7 1 2 11281 11285
0 11287 5 1 1 11286
0 11288 7 2 2 65132 87163
0 11289 7 1 2 63936 87686
0 11290 7 1 2 11287 11289
0 11291 5 1 1 11290
0 11292 7 1 2 11270 11291
0 11293 5 1 1 11292
0 11294 7 1 2 81159 11293
0 11295 5 1 1 11294
0 11296 7 1 2 11264 11295
0 11297 5 1 1 11296
0 11298 7 1 2 87653 11297
0 11299 5 1 1 11298
0 11300 7 1 2 11250 11299
0 11301 7 1 2 11111 11300
0 11302 7 1 2 10992 11301
0 11303 7 1 2 10805 11302
0 11304 7 1 2 10652 11303
0 11305 5 1 1 11304
0 11306 7 1 2 63677 11305
0 11307 5 1 1 11306
0 11308 7 1 2 67249 75912
0 11309 5 3 1 11308
0 11310 7 1 2 64451 78903
0 11311 5 1 1 11310
0 11312 7 1 2 62059 85221
0 11313 5 1 1 11312
0 11314 7 1 2 11311 11313
0 11315 5 1 1 11314
0 11316 7 1 2 64240 11315
0 11317 5 1 1 11316
0 11318 7 1 2 10480 11317
0 11319 5 1 1 11318
0 11320 7 1 2 61457 11319
0 11321 5 1 1 11320
0 11322 7 1 2 64241 81920
0 11323 7 1 2 86041 11322
0 11324 5 1 1 11323
0 11325 7 1 2 11321 11324
0 11326 5 1 1 11325
0 11327 7 1 2 64925 11326
0 11328 5 1 1 11327
0 11329 7 2 2 67893 86908
0 11330 5 1 1 87691
0 11331 7 1 2 86891 11330
0 11332 5 1 1 11331
0 11333 7 1 2 64242 11332
0 11334 5 1 1 11333
0 11335 7 1 2 11115 11334
0 11336 5 1 1 11335
0 11337 7 1 2 79520 11336
0 11338 5 1 1 11337
0 11339 7 1 2 11328 11338
0 11340 5 1 1 11339
0 11341 7 1 2 63678 11340
0 11342 5 1 1 11341
0 11343 7 2 2 79555 79004
0 11344 7 1 2 81973 87693
0 11345 5 1 1 11344
0 11346 7 1 2 11342 11345
0 11347 5 1 1 11346
0 11348 7 1 2 87386 11347
0 11349 5 1 1 11348
0 11350 7 1 2 59476 79838
0 11351 5 3 1 11350
0 11352 7 1 2 82014 87695
0 11353 5 1 1 11352
0 11354 7 1 2 62060 75186
0 11355 7 1 2 82533 11354
0 11356 5 1 1 11355
0 11357 7 1 2 11353 11356
0 11358 5 1 1 11357
0 11359 7 2 2 67894 86699
0 11360 7 4 2 68842 78154
0 11361 7 1 2 87698 87700
0 11362 7 1 2 11358 11361
0 11363 5 1 1 11362
0 11364 7 1 2 11349 11363
0 11365 5 1 1 11364
0 11366 7 1 2 63356 11365
0 11367 5 1 1 11366
0 11368 7 2 2 86700 86922
0 11369 7 1 2 82530 87606
0 11370 7 1 2 86465 11369
0 11371 7 1 2 87704 11370
0 11372 5 1 1 11371
0 11373 7 1 2 11367 11372
0 11374 5 1 1 11373
0 11375 7 1 2 81160 11374
0 11376 5 1 1 11375
0 11377 7 1 2 80842 87164
0 11378 5 3 1 11377
0 11379 7 4 2 65358 60653
0 11380 7 5 2 85841 87709
0 11381 5 4 1 87713
0 11382 7 2 2 87706 87718
0 11383 5 4 1 87722
0 11384 7 1 2 79371 87574
0 11385 7 1 2 87696 11384
0 11386 7 1 2 87724 11385
0 11387 5 1 1 11386
0 11388 7 8 2 67895 70754
0 11389 5 1 1 87728
0 11390 7 1 2 87697 87729
0 11391 5 1 1 11390
0 11392 7 1 2 9023 11391
0 11393 5 1 1 11392
0 11394 7 1 2 79521 11393
0 11395 5 1 1 11394
0 11396 7 1 2 5281 11395
0 11397 5 1 1 11396
0 11398 7 1 2 84767 87500
0 11399 7 1 2 11397 11398
0 11400 5 1 1 11399
0 11401 7 1 2 11387 11400
0 11402 5 1 1 11401
0 11403 7 1 2 63357 11402
0 11404 5 1 1 11403
0 11405 7 3 2 81527 79005
0 11406 5 1 1 87736
0 11407 7 1 2 70445 87737
0 11408 7 1 2 82028 11407
0 11409 7 1 2 87501 11408
0 11410 5 1 1 11409
0 11411 7 1 2 11404 11410
0 11412 5 1 1 11411
0 11413 7 1 2 63937 11412
0 11414 5 1 1 11413
0 11415 7 1 2 79923 86962
0 11416 7 1 2 82534 11415
0 11417 7 2 2 77895 85503
0 11418 7 1 2 87648 87739
0 11419 7 1 2 11416 11418
0 11420 5 1 1 11419
0 11421 7 1 2 11414 11420
0 11422 7 1 2 11376 11421
0 11423 5 1 1 11422
0 11424 7 1 2 87688 11423
0 11425 5 1 1 11424
0 11426 7 1 2 67896 76882
0 11427 5 2 1 11426
0 11428 7 2 2 64452 86043
0 11429 5 1 1 87743
0 11430 7 1 2 87352 11429
0 11431 7 1 2 87741 11430
0 11432 5 1 1 11431
0 11433 7 1 2 67024 87353
0 11434 5 2 1 11433
0 11435 7 1 2 63358 87745
0 11436 7 1 2 11432 11435
0 11437 5 1 1 11436
0 11438 7 1 2 85958 11437
0 11439 5 1 1 11438
0 11440 7 1 2 60266 11439
0 11441 5 1 1 11440
0 11442 7 1 2 81528 79098
0 11443 5 1 1 11442
0 11444 7 1 2 64453 81969
0 11445 7 1 2 84676 11444
0 11446 5 1 1 11445
0 11447 7 1 2 11443 11446
0 11448 5 1 1 11447
0 11449 7 1 2 61246 11448
0 11450 5 1 1 11449
0 11451 7 3 2 70755 77090
0 11452 7 2 2 65133 74221
0 11453 5 2 1 87750
0 11454 7 1 2 67897 87751
0 11455 7 1 2 87747 11454
0 11456 5 1 1 11455
0 11457 7 1 2 66421 11456
0 11458 7 1 2 11450 11457
0 11459 7 1 2 11441 11458
0 11460 5 1 1 11459
0 11461 7 10 2 67898 70591
0 11462 5 4 1 87754
0 11463 7 3 2 63359 87764
0 11464 5 1 1 87768
0 11465 7 1 2 74008 77496
0 11466 7 1 2 87769 11465
0 11467 7 1 2 60267 86549
0 11468 5 2 1 11467
0 11469 7 1 2 87771 87746
0 11470 7 1 2 11466 11469
0 11471 5 1 1 11470
0 11472 7 3 2 65134 81529
0 11473 5 1 1 87773
0 11474 7 1 2 79347 87774
0 11475 5 1 1 11474
0 11476 7 1 2 61458 11475
0 11477 7 1 2 11471 11476
0 11478 5 1 1 11477
0 11479 7 1 2 63679 11478
0 11480 7 1 2 11460 11479
0 11481 5 1 1 11480
0 11482 7 2 2 74009 83517
0 11483 7 2 2 74927 85061
0 11484 5 1 1 87778
0 11485 7 1 2 77962 87779
0 11486 7 1 2 87776 11485
0 11487 5 1 1 11486
0 11488 7 1 2 11481 11487
0 11489 5 1 1 11488
0 11490 7 1 2 81161 11489
0 11491 5 1 1 11490
0 11492 7 2 2 67250 73354
0 11493 5 4 1 87780
0 11494 7 1 2 79372 85471
0 11495 5 1 1 11494
0 11496 7 2 2 70756 79326
0 11497 7 6 2 66659 84768
0 11498 5 1 1 87788
0 11499 7 1 2 84376 87789
0 11500 7 1 2 87786 11499
0 11501 5 1 1 11500
0 11502 7 1 2 11495 11501
0 11503 5 1 1 11502
0 11504 7 1 2 87782 11503
0 11505 5 1 1 11504
0 11506 7 2 2 83470 84005
0 11507 7 2 2 79006 87794
0 11508 7 1 2 79610 83326
0 11509 7 1 2 87796 11508
0 11510 5 1 1 11509
0 11511 7 1 2 11505 11510
0 11512 5 1 1 11511
0 11513 7 1 2 63360 11512
0 11514 5 1 1 11513
0 11515 7 6 2 68277 79611
0 11516 5 1 1 87798
0 11517 7 3 2 67899 75478
0 11518 7 2 2 63680 70757
0 11519 7 1 2 87804 87807
0 11520 5 1 1 11519
0 11521 7 4 2 62899 74010
0 11522 5 2 1 87809
0 11523 7 1 2 68617 87810
0 11524 7 1 2 82029 11523
0 11525 5 1 1 11524
0 11526 7 1 2 11520 11525
0 11527 5 1 1 11526
0 11528 7 1 2 62546 11527
0 11529 5 1 1 11528
0 11530 7 2 2 75479 73094
0 11531 7 1 2 87815 87808
0 11532 5 1 1 11531
0 11533 7 1 2 83621 82542
0 11534 5 1 1 11533
0 11535 7 1 2 11532 11534
0 11536 5 1 1 11535
0 11537 7 1 2 67900 11536
0 11538 5 1 1 11537
0 11539 7 1 2 11529 11538
0 11540 5 1 1 11539
0 11541 7 1 2 62061 11540
0 11542 5 1 1 11541
0 11543 7 1 2 79386 87513
0 11544 5 1 1 11543
0 11545 7 1 2 11542 11544
0 11546 5 1 1 11545
0 11547 7 1 2 87799 11546
0 11548 5 1 1 11547
0 11549 7 1 2 11514 11548
0 11550 7 1 2 11491 11549
0 11551 5 1 1 11550
0 11552 7 1 2 63938 11551
0 11553 5 1 1 11552
0 11554 7 3 2 82040 79373
0 11555 5 1 1 87817
0 11556 7 7 2 65359 66422
0 11557 5 6 1 87820
0 11558 7 2 2 81907 87821
0 11559 7 1 2 71024 87308
0 11560 7 1 2 87833 11559
0 11561 7 1 2 87818 11560
0 11562 5 1 1 11561
0 11563 7 1 2 11553 11562
0 11564 5 1 1 11563
0 11565 7 1 2 86777 11564
0 11566 5 1 1 11565
0 11567 7 3 2 81749 84769
0 11568 7 1 2 87787 87835
0 11569 5 1 1 11568
0 11570 7 1 2 81396 86867
0 11571 5 2 1 11570
0 11572 7 1 2 81162 86524
0 11573 5 1 1 11572
0 11574 7 1 2 87838 11573
0 11575 5 1 1 11574
0 11576 7 1 2 87701 11575
0 11577 5 1 1 11576
0 11578 7 1 2 11569 11577
0 11579 5 1 1 11578
0 11580 7 1 2 87699 11579
0 11581 5 1 1 11580
0 11582 7 7 2 65360 71025
0 11583 7 3 2 60654 66200
0 11584 7 2 2 87840 87847
0 11585 7 21 2 63681 63939
0 11586 7 2 2 79481 85842
0 11587 5 1 1 87873
0 11588 7 2 2 87852 87874
0 11589 7 1 2 87850 87875
0 11590 5 1 1 11589
0 11591 7 1 2 11581 11590
0 11592 5 1 1 11591
0 11593 7 1 2 87783 11592
0 11594 5 1 1 11593
0 11595 7 6 2 65135 62258
0 11596 7 2 2 75412 85504
0 11597 7 1 2 87877 87883
0 11598 5 1 1 11597
0 11599 7 2 2 75480 77542
0 11600 5 2 1 87885
0 11601 7 1 2 11598 87887
0 11602 5 1 1 11601
0 11603 7 1 2 70036 11602
0 11604 5 1 1 11603
0 11605 7 6 2 61247 68618
0 11606 7 1 2 80828 87889
0 11607 5 1 1 11606
0 11608 7 1 2 11604 11607
0 11609 5 1 1 11608
0 11610 7 1 2 61664 11609
0 11611 5 1 1 11610
0 11612 7 3 2 62259 81284
0 11613 7 1 2 80138 85505
0 11614 7 1 2 87895 11613
0 11615 5 1 1 11614
0 11616 7 1 2 11611 11615
0 11617 5 1 1 11616
0 11618 7 1 2 64454 11617
0 11619 5 1 1 11618
0 11620 7 2 2 79359 77543
0 11621 7 1 2 87795 87898
0 11622 5 1 1 11621
0 11623 7 1 2 11619 11622
0 11624 5 1 1 11623
0 11625 7 1 2 60452 11624
0 11626 5 1 1 11625
0 11627 7 1 2 85506 85774
0 11628 7 1 2 80522 11627
0 11629 7 1 2 87816 11628
0 11630 5 1 1 11629
0 11631 7 1 2 11626 11630
0 11632 5 1 1 11631
0 11633 7 1 2 77461 86701
0 11634 7 1 2 11632 11633
0 11635 5 1 1 11634
0 11636 7 1 2 11594 11635
0 11637 5 1 1 11636
0 11638 7 1 2 63361 11637
0 11639 5 1 1 11638
0 11640 7 3 2 68278 86702
0 11641 7 1 2 62062 81750
0 11642 7 1 2 87748 11641
0 11643 5 1 1 11642
0 11644 7 3 2 62260 86909
0 11645 5 1 1 87903
0 11646 7 1 2 80678 77021
0 11647 7 1 2 87904 11646
0 11648 5 1 1 11647
0 11649 7 1 2 11643 11648
0 11650 5 1 1 11649
0 11651 7 1 2 83840 11650
0 11652 5 1 1 11651
0 11653 7 4 2 67525 77544
0 11654 7 1 2 71026 85775
0 11655 7 1 2 81033 11654
0 11656 7 1 2 87906 11655
0 11657 5 1 1 11656
0 11658 7 1 2 11652 11657
0 11659 5 1 1 11658
0 11660 7 1 2 67901 11659
0 11661 5 1 1 11660
0 11662 7 1 2 75413 74011
0 11663 7 1 2 83444 11662
0 11664 5 1 1 11663
0 11665 7 1 2 83677 11664
0 11666 5 1 1 11665
0 11667 7 8 2 60453 78051
0 11668 5 3 1 87910
0 11669 7 1 2 87372 87911
0 11670 7 1 2 11666 11669
0 11671 5 1 1 11670
0 11672 7 1 2 11661 11671
0 11673 7 2 2 79007 86579
0 11674 7 5 2 61665 62547
0 11675 7 3 2 60454 87923
0 11676 7 1 2 70037 87928
0 11677 7 1 2 87921 11676
0 11678 5 1 1 11677
0 11679 7 4 2 79612 85507
0 11680 7 1 2 73612 87755
0 11681 7 1 2 87931 11680
0 11682 5 1 1 11681
0 11683 7 1 2 11678 11682
0 11684 5 1 1 11683
0 11685 7 1 2 64455 11684
0 11686 5 1 1 11685
0 11687 7 2 2 70480 78550
0 11688 5 1 1 87935
0 11689 7 1 2 64926 87936
0 11690 7 1 2 87836 11689
0 11691 5 1 1 11690
0 11692 7 1 2 11686 11691
0 11693 5 1 1 11692
0 11694 7 1 2 79327 11693
0 11695 5 1 1 11694
0 11696 7 2 2 79008 87045
0 11697 7 1 2 84023 87937
0 11698 5 1 1 11697
0 11699 7 6 2 68843 86380
0 11700 7 2 2 70038 73613
0 11701 5 1 1 87945
0 11702 7 1 2 78904 87946
0 11703 7 1 2 87939 11702
0 11704 5 1 1 11703
0 11705 7 1 2 11698 11704
0 11706 5 1 1 11705
0 11707 7 1 2 64456 11706
0 11708 5 1 1 11707
0 11709 7 1 2 76129 78695
0 11710 5 2 1 11709
0 11711 7 1 2 86559 87947
0 11712 5 1 1 11711
0 11713 7 7 2 68619 75481
0 11714 7 1 2 86580 87949
0 11715 7 1 2 11712 11714
0 11716 5 1 1 11715
0 11717 7 1 2 11708 11716
0 11718 5 1 1 11717
0 11719 7 1 2 81163 11718
0 11720 5 1 1 11719
0 11721 7 1 2 11695 11720
0 11722 7 1 2 11672 11721
0 11723 5 1 1 11722
0 11724 7 1 2 87900 11723
0 11725 5 1 1 11724
0 11726 7 1 2 11639 11725
0 11727 7 1 2 11566 11726
0 11728 5 1 1 11727
0 11729 7 1 2 72546 11728
0 11730 5 1 1 11729
0 11731 7 1 2 70039 74053
0 11732 5 2 1 11731
0 11733 7 3 2 70481 86947
0 11734 5 1 1 87958
0 11735 7 1 2 70133 11734
0 11736 5 1 1 11735
0 11737 7 1 2 86599 11736
0 11738 5 1 1 11737
0 11739 7 1 2 87956 11738
0 11740 5 1 1 11739
0 11741 7 1 2 67902 11740
0 11742 5 1 1 11741
0 11743 7 1 2 77370 87959
0 11744 5 1 1 11743
0 11745 7 2 2 61248 78696
0 11746 5 1 1 87961
0 11747 7 1 2 86898 87962
0 11748 5 1 1 11747
0 11749 7 1 2 87379 11748
0 11750 5 1 1 11749
0 11751 7 1 2 70307 11750
0 11752 5 1 1 11751
0 11753 7 1 2 11744 11752
0 11754 7 1 2 11742 11753
0 11755 5 1 1 11754
0 11756 7 1 2 63362 11755
0 11757 5 1 1 11756
0 11758 7 1 2 70134 87330
0 11759 5 1 1 11758
0 11760 7 3 2 67903 85009
0 11761 5 2 1 87963
0 11762 7 1 2 11759 87964
0 11763 5 1 1 11762
0 11764 7 1 2 72434 80623
0 11765 5 1 1 11764
0 11766 7 1 2 61249 79830
0 11767 5 1 1 11766
0 11768 7 1 2 11765 11767
0 11769 5 1 1 11768
0 11770 7 1 2 71758 11769
0 11771 5 1 1 11770
0 11772 7 1 2 80624 76717
0 11773 5 1 1 11772
0 11774 7 5 2 64457 63363
0 11775 5 2 1 87968
0 11776 7 1 2 61250 87969
0 11777 5 1 1 11776
0 11778 7 1 2 11773 11777
0 11779 5 1 1 11778
0 11780 7 1 2 70403 11779
0 11781 5 1 1 11780
0 11782 7 1 2 63364 86336
0 11783 5 1 1 11782
0 11784 7 1 2 80625 87284
0 11785 5 1 1 11784
0 11786 7 1 2 11783 11785
0 11787 7 1 2 11781 11786
0 11788 7 1 2 11771 11787
0 11789 5 1 1 11788
0 11790 7 1 2 62900 11789
0 11791 5 1 1 11790
0 11792 7 1 2 11763 11791
0 11793 5 1 1 11792
0 11794 7 1 2 62548 11793
0 11795 5 1 1 11794
0 11796 7 1 2 11757 11795
0 11797 5 1 1 11796
0 11798 7 1 2 79522 87502
0 11799 7 1 2 11797 11798
0 11800 5 1 1 11799
0 11801 7 2 2 65827 81420
0 11802 5 2 1 87975
0 11803 7 1 2 77046 87976
0 11804 5 1 1 11803
0 11805 7 1 2 62261 76039
0 11806 5 1 1 11805
0 11807 7 1 2 11804 11806
0 11808 5 1 1 11807
0 11809 7 1 2 62549 11808
0 11810 5 1 1 11809
0 11811 7 1 2 85244 11810
0 11812 5 1 1 11811
0 11813 7 1 2 77371 11812
0 11814 5 1 1 11813
0 11815 7 1 2 72454 6210
0 11816 5 1 1 11815
0 11817 7 1 2 64458 70514
0 11818 7 1 2 11816 11817
0 11819 5 1 1 11818
0 11820 7 2 2 65828 73685
0 11821 7 1 2 69784 87979
0 11822 5 1 1 11821
0 11823 7 1 2 11819 11822
0 11824 5 1 1 11823
0 11825 7 1 2 87027 11824
0 11826 5 1 1 11825
0 11827 7 2 2 64459 73614
0 11828 5 1 1 87981
0 11829 7 2 2 74407 11828
0 11830 5 3 1 87983
0 11831 7 1 2 72876 74012
0 11832 5 1 1 11831
0 11833 7 1 2 78474 11832
0 11834 5 1 1 11833
0 11835 7 1 2 67526 11834
0 11836 5 1 1 11835
0 11837 7 1 2 87984 11836
0 11838 5 1 1 11837
0 11839 7 1 2 70040 11838
0 11840 5 1 1 11839
0 11841 7 1 2 11826 11840
0 11842 5 1 1 11841
0 11843 7 1 2 67904 11842
0 11844 5 1 1 11843
0 11845 7 1 2 11814 11844
0 11846 5 1 1 11845
0 11847 7 1 2 66823 80577
0 11848 5 1 1 11847
0 11849 7 1 2 86068 11848
0 11850 5 1 1 11849
0 11851 7 1 2 65552 11850
0 11852 5 1 1 11851
0 11853 7 1 2 75187 87065
0 11854 7 1 2 87710 11853
0 11855 5 1 1 11854
0 11856 7 1 2 11852 11855
0 11857 5 1 1 11856
0 11858 7 1 2 68279 11857
0 11859 7 1 2 11846 11858
0 11860 5 1 1 11859
0 11861 7 1 2 65697 82470
0 11862 5 2 1 11861
0 11863 7 1 2 76661 87988
0 11864 5 1 1 11863
0 11865 7 1 2 64460 11864
0 11866 5 1 1 11865
0 11867 7 1 2 72826 77091
0 11868 5 1 1 11867
0 11869 7 1 2 78878 11868
0 11870 5 1 1 11869
0 11871 7 1 2 64243 11870
0 11872 5 1 1 11871
0 11873 7 1 2 11866 11872
0 11874 5 1 1 11873
0 11875 7 1 2 84245 86778
0 11876 5 1 1 11875
0 11877 7 1 2 87223 11876
0 11878 5 1 1 11877
0 11879 7 1 2 78551 84408
0 11880 7 1 2 11878 11879
0 11881 7 1 2 11874 11880
0 11882 5 1 1 11881
0 11883 7 1 2 11860 11882
0 11884 7 1 2 11800 11883
0 11885 5 1 1 11884
0 11886 7 1 2 63940 11885
0 11887 5 1 1 11886
0 11888 7 1 2 80531 72755
0 11889 7 1 2 87679 87406
0 11890 7 6 2 66423 66824
0 11891 7 6 2 65553 66660
0 11892 7 3 2 87990 87996
0 11893 7 4 2 65361 74094
0 11894 5 1 1 88005
0 11895 7 1 2 88002 88006
0 11896 7 1 2 11889 11895
0 11897 7 1 2 11888 11896
0 11898 5 1 1 11897
0 11899 7 1 2 80532 87066
0 11900 7 1 2 79523 11899
0 11901 7 8 2 67025 78248
0 11902 7 8 2 65362 65554
0 11903 7 2 2 70041 88017
0 11904 7 1 2 88009 88025
0 11905 7 1 2 11900 11904
0 11906 7 1 2 74465 11905
0 11907 5 1 1 11906
0 11908 7 1 2 11898 11907
0 11909 7 1 2 11887 11908
0 11910 5 1 1 11909
0 11911 7 1 2 68620 11910
0 11912 5 1 1 11911
0 11913 7 1 2 11730 11912
0 11914 7 1 2 11425 11913
0 11915 7 1 2 11307 11914
0 11916 5 1 1 11915
0 11917 7 1 2 72290 11916
0 11918 5 1 1 11917
0 11919 7 1 2 67905 79417
0 11920 5 4 1 11919
0 11921 7 4 2 85878 87088
0 11922 5 1 1 88031
0 11923 7 1 2 88027 88032
0 11924 5 1 1 11923
0 11925 7 1 2 67527 84088
0 11926 5 6 1 11925
0 11927 7 1 2 64461 88035
0 11928 5 2 1 11927
0 11929 7 1 2 76662 88041
0 11930 5 4 1 11929
0 11931 7 2 2 68844 88043
0 11932 7 3 2 65555 87662
0 11933 7 2 2 80843 88049
0 11934 7 1 2 88047 88052
0 11935 5 1 1 11934
0 11936 7 1 2 11924 11935
0 11937 5 1 1 11936
0 11938 7 1 2 66424 11937
0 11939 5 1 1 11938
0 11940 7 4 2 68845 80403
0 11941 7 3 2 67906 86391
0 11942 7 1 2 86994 88058
0 11943 7 1 2 88054 11942
0 11944 5 1 1 11943
0 11945 7 1 2 11939 11944
0 11946 5 1 1 11945
0 11947 7 1 2 65136 11946
0 11948 5 1 1 11947
0 11949 7 1 2 83896 88044
0 11950 5 1 1 11949
0 11951 7 1 2 85074 11950
0 11952 5 1 1 11951
0 11953 7 2 2 68846 87590
0 11954 5 1 1 88061
0 11955 7 1 2 65556 80404
0 11956 7 1 2 88062 11955
0 11957 7 1 2 11952 11956
0 11958 5 1 1 11957
0 11959 7 1 2 11948 11958
0 11960 5 1 1 11959
0 11961 7 1 2 70042 11960
0 11962 5 1 1 11961
0 11963 7 1 2 81397 79300
0 11964 5 1 1 11963
0 11965 7 1 2 72750 82397
0 11966 5 1 1 11965
0 11967 7 2 2 62901 70446
0 11968 5 1 1 88063
0 11969 7 1 2 65698 88064
0 11970 7 1 2 85163 11969
0 11971 5 1 1 11970
0 11972 7 1 2 11966 11971
0 11973 5 1 1 11972
0 11974 7 1 2 81164 11973
0 11975 5 1 1 11974
0 11976 7 1 2 11964 11975
0 11977 5 1 1 11976
0 11978 7 12 2 68847 86703
0 11979 7 1 2 73909 88065
0 11980 7 1 2 11977 11979
0 11981 5 1 1 11980
0 11982 7 1 2 11962 11981
0 11983 5 1 1 11982
0 11984 7 1 2 63365 11983
0 11985 5 1 1 11984
0 11986 7 2 2 62902 86130
0 11987 7 1 2 80205 86055
0 11988 7 1 2 88077 11987
0 11989 5 1 1 11988
0 11990 7 14 2 61666 67907
0 11991 7 3 2 63941 88079
0 11992 7 16 2 61459 67251
0 11993 5 2 1 88096
0 11994 7 1 2 77022 88097
0 11995 7 1 2 88093 11994
0 11996 5 1 1 11995
0 11997 7 1 2 61251 11996
0 11998 7 1 2 11989 11997
0 11999 5 1 1 11998
0 12000 7 12 2 66661 62903
0 12001 7 1 2 81290 77347
0 12002 7 1 2 88114 12001
0 12003 7 1 2 79328 12002
0 12004 5 1 1 12003
0 12005 7 1 2 79051 86641
0 12006 5 1 1 12005
0 12007 7 1 2 66201 12006
0 12008 7 1 2 12004 12007
0 12009 5 1 1 12008
0 12010 7 1 2 60455 12009
0 12011 7 1 2 11999 12010
0 12012 5 1 1 12011
0 12013 7 1 2 70043 81378
0 12014 5 1 1 12013
0 12015 7 1 2 81375 12014
0 12016 5 1 1 12015
0 12017 7 6 2 65363 68848
0 12018 7 1 2 87424 88126
0 12019 7 1 2 12016 12018
0 12020 5 1 1 12019
0 12021 7 1 2 12012 12020
0 12022 5 1 1 12021
0 12023 7 1 2 64462 12022
0 12024 5 1 1 12023
0 12025 7 8 2 60456 81490
0 12026 5 2 1 88132
0 12027 7 1 2 62262 81089
0 12028 7 1 2 87730 12027
0 12029 7 1 2 88133 12028
0 12030 5 1 1 12029
0 12031 7 1 2 12024 12030
0 12032 5 1 1 12031
0 12033 7 1 2 87901 12032
0 12034 5 1 1 12033
0 12035 7 1 2 11985 12034
0 12036 5 1 1 12035
0 12037 7 1 2 63682 12036
0 12038 5 1 1 12037
0 12039 7 2 2 77545 86704
0 12040 7 1 2 79329 77092
0 12041 7 1 2 87731 12040
0 12042 5 1 1 12041
0 12043 7 2 2 69785 81047
0 12044 5 1 1 88144
0 12045 7 1 2 85658 88145
0 12046 7 1 2 78833 12045
0 12047 5 1 1 12046
0 12048 7 1 2 12042 12047
0 12049 5 1 1 12048
0 12050 7 1 2 63366 12049
0 12051 5 1 1 12050
0 12052 7 1 2 11056 12051
0 12053 5 1 1 12052
0 12054 7 1 2 61667 12053
0 12055 5 1 1 12054
0 12056 7 1 2 87520 88115
0 12057 5 1 1 12056
0 12058 7 1 2 12055 12057
0 12059 5 1 1 12058
0 12060 7 1 2 60457 12059
0 12061 5 1 1 12060
0 12062 7 1 2 81530 74676
0 12063 7 1 2 81387 86535
0 12064 7 1 2 12062 12063
0 12065 5 1 1 12064
0 12066 7 1 2 12061 12065
0 12067 5 1 1 12066
0 12068 7 1 2 88142 12067
0 12069 5 1 1 12068
0 12070 7 1 2 12038 12069
0 12071 5 1 1 12070
0 12072 7 1 2 64691 12071
0 12073 5 1 1 12072
0 12074 7 3 2 80946 73473
0 12075 7 6 2 68621 86705
0 12076 7 1 2 80646 88149
0 12077 7 1 2 88146 12076
0 12078 7 1 2 84924 12077
0 12079 5 1 1 12078
0 12080 7 1 2 12073 12079
0 12081 5 1 1 12080
0 12082 7 1 2 65976 12081
0 12083 5 1 1 12082
0 12084 7 2 2 63942 86706
0 12085 7 1 2 76957 82223
0 12086 7 1 2 80578 12085
0 12087 5 1 1 12086
0 12088 7 1 2 80844 77093
0 12089 7 1 2 82015 12088
0 12090 5 1 1 12089
0 12091 7 1 2 12087 12090
0 12092 5 1 1 12091
0 12093 7 1 2 83518 12092
0 12094 5 1 1 12093
0 12095 7 1 2 74254 79071
0 12096 5 1 1 12095
0 12097 7 4 2 61252 74728
0 12098 5 1 1 88157
0 12099 7 1 2 67252 88158
0 12100 5 1 1 12099
0 12101 7 1 2 84936 12100
0 12102 5 1 1 12101
0 12103 7 1 2 60268 74013
0 12104 7 1 2 12102 12103
0 12105 5 1 1 12104
0 12106 7 1 2 12096 12105
0 12107 5 1 1 12106
0 12108 7 1 2 85151 12107
0 12109 5 1 1 12108
0 12110 7 1 2 12094 12109
0 12111 5 1 1 12110
0 12112 7 1 2 67908 12111
0 12113 5 1 1 12112
0 12114 7 4 2 60458 62550
0 12115 5 5 1 88161
0 12116 7 1 2 81101 88162
0 12117 7 1 2 83774 12116
0 12118 7 1 2 87797 12117
0 12119 5 1 1 12118
0 12120 7 1 2 12113 12119
0 12121 5 1 1 12120
0 12122 7 1 2 88155 12121
0 12123 5 1 1 12122
0 12124 7 1 2 80589 76888
0 12125 5 2 1 12124
0 12126 7 3 2 70253 88170
0 12127 5 1 1 88172
0 12128 7 3 2 81295 85441
0 12129 7 1 2 88173 88175
0 12130 5 1 1 12129
0 12131 7 1 2 71380 86508
0 12132 5 1 1 12131
0 12133 7 3 2 66662 71355
0 12134 5 1 1 88178
0 12135 7 1 2 74677 88179
0 12136 5 1 1 12135
0 12137 7 1 2 79278 12136
0 12138 5 1 1 12137
0 12139 7 1 2 77829 12138
0 12140 5 1 1 12139
0 12141 7 1 2 12132 12140
0 12142 5 1 1 12141
0 12143 7 1 2 64463 12142
0 12144 5 1 1 12143
0 12145 7 1 2 62263 77732
0 12146 5 2 1 12145
0 12147 7 1 2 64464 78502
0 12148 5 1 1 12147
0 12149 7 1 2 88181 12148
0 12150 5 1 1 12149
0 12151 7 1 2 80193 12150
0 12152 5 1 1 12151
0 12153 7 1 2 12144 12152
0 12154 5 1 1 12153
0 12155 7 1 2 65364 12154
0 12156 5 1 1 12155
0 12157 7 1 2 12130 12156
0 12158 5 1 1 12157
0 12159 7 1 2 84424 12158
0 12160 5 1 1 12159
0 12161 7 8 2 65365 62904
0 12162 5 1 1 88183
0 12163 7 10 2 66663 62551
0 12164 5 1 1 88191
0 12165 7 2 2 65977 68622
0 12166 5 1 1 88201
0 12167 7 2 2 88192 88202
0 12168 5 1 1 88203
0 12169 7 2 2 64692 88204
0 12170 5 1 1 88205
0 12171 7 1 2 88184 88206
0 12172 7 1 2 82030 12171
0 12173 5 1 1 12172
0 12174 7 1 2 12160 12173
0 12175 5 1 1 12174
0 12176 7 1 2 68280 12175
0 12177 5 1 1 12176
0 12178 7 1 2 61668 79578
0 12179 5 1 1 12178
0 12180 7 1 2 79303 12179
0 12181 5 1 1 12180
0 12182 7 1 2 64927 12181
0 12183 5 1 1 12182
0 12184 7 1 2 80165 86044
0 12185 5 1 1 12184
0 12186 7 1 2 70044 79255
0 12187 5 2 1 12186
0 12188 7 1 2 79304 88207
0 12189 5 1 1 12188
0 12190 7 1 2 79414 12189
0 12191 5 1 1 12190
0 12192 7 1 2 12185 12191
0 12193 7 1 2 12183 12192
0 12194 5 1 1 12193
0 12195 7 1 2 65137 12194
0 12196 5 1 1 12195
0 12197 7 1 2 67909 85582
0 12198 5 1 1 12197
0 12199 7 1 2 78205 84464
0 12200 7 1 2 12198 12199
0 12201 5 1 1 12200
0 12202 7 1 2 66664 84967
0 12203 7 1 2 12201 12202
0 12204 5 1 1 12203
0 12205 7 1 2 12196 12204
0 12206 5 1 1 12205
0 12207 7 1 2 71090 12206
0 12208 5 1 1 12207
0 12209 7 1 2 83024 76891
0 12210 5 1 1 12209
0 12211 7 1 2 62905 77025
0 12212 5 1 1 12211
0 12213 7 1 2 79330 12212
0 12214 7 1 2 12210 12213
0 12215 5 1 1 12214
0 12216 7 5 2 66202 82602
0 12217 5 1 1 88209
0 12218 7 1 2 79099 88210
0 12219 5 1 1 12218
0 12220 7 1 2 12215 12219
0 12221 5 1 1 12220
0 12222 7 1 2 66665 12221
0 12223 5 1 1 12222
0 12224 7 1 2 12208 12223
0 12225 5 1 1 12224
0 12226 7 1 2 63683 12225
0 12227 5 1 1 12226
0 12228 7 2 2 78618 77513
0 12229 5 1 1 88214
0 12230 7 1 2 86056 88215
0 12231 7 1 2 85171 12230
0 12232 5 1 1 12231
0 12233 7 1 2 60459 12232
0 12234 7 1 2 12227 12233
0 12235 5 1 1 12234
0 12236 7 1 2 76958 74871
0 12237 5 1 1 12236
0 12238 7 1 2 61460 70254
0 12239 7 1 2 87749 12238
0 12240 5 1 1 12239
0 12241 7 1 2 12237 12240
0 12242 5 1 1 12241
0 12243 7 1 2 84332 12242
0 12244 5 1 1 12243
0 12245 7 3 2 63684 81491
0 12246 5 1 1 88216
0 12247 7 1 2 77748 74236
0 12248 5 1 1 12247
0 12249 7 1 2 88217 12248
0 12250 5 1 1 12249
0 12251 7 1 2 12244 12250
0 12252 5 1 1 12251
0 12253 7 1 2 65138 12252
0 12254 5 1 1 12253
0 12255 7 2 2 84158 83647
0 12256 5 1 1 88219
0 12257 7 1 2 85218 12256
0 12258 7 1 2 8596 12257
0 12259 5 1 1 12258
0 12260 7 1 2 73095 12259
0 12261 5 1 1 12260
0 12262 7 4 2 66203 84473
0 12263 5 1 1 88221
0 12264 7 1 2 72700 88222
0 12265 5 1 1 12264
0 12266 7 1 2 77733 87790
0 12267 5 1 1 12266
0 12268 7 1 2 12265 12267
0 12269 7 1 2 12261 12268
0 12270 5 1 1 12269
0 12271 7 1 2 75873 12270
0 12272 5 1 1 12271
0 12273 7 5 2 64465 61669
0 12274 7 9 2 62264 63685
0 12275 7 2 2 88225 88230
0 12276 5 2 1 88239
0 12277 7 1 2 77830 81061
0 12278 7 1 2 88240 12277
0 12279 5 1 1 12278
0 12280 7 1 2 67910 12279
0 12281 7 1 2 12272 12280
0 12282 7 1 2 12254 12281
0 12283 5 1 1 12282
0 12284 7 2 2 78028 84770
0 12285 7 5 2 64244 65139
0 12286 5 2 1 88245
0 12287 7 3 2 77233 88246
0 12288 5 1 1 88252
0 12289 7 1 2 88243 88253
0 12290 5 1 1 12289
0 12291 7 1 2 60269 78155
0 12292 5 1 1 12291
0 12293 7 1 2 12290 12292
0 12294 5 1 1 12293
0 12295 7 1 2 72701 12294
0 12296 5 1 1 12295
0 12297 7 2 2 71027 84771
0 12298 7 1 2 77315 70935
0 12299 7 1 2 88255 12298
0 12300 5 1 1 12299
0 12301 7 1 2 12296 12300
0 12302 5 1 1 12301
0 12303 7 1 2 61670 12302
0 12304 5 1 1 12303
0 12305 7 2 2 84129 87791
0 12306 5 1 1 88257
0 12307 7 1 2 60270 88258
0 12308 5 1 1 12307
0 12309 7 1 2 12304 12308
0 12310 5 1 1 12309
0 12311 7 1 2 66425 12310
0 12312 5 1 1 12311
0 12313 7 6 2 61671 78156
0 12314 5 1 1 88259
0 12315 7 1 2 66204 88260
0 12316 5 1 1 12315
0 12317 7 1 2 12306 12316
0 12318 5 1 1 12317
0 12319 7 1 2 77181 12318
0 12320 5 1 1 12319
0 12321 7 1 2 78157 86419
0 12322 5 1 1 12321
0 12323 7 1 2 78619 85591
0 12324 7 1 2 88244 12323
0 12325 5 1 1 12324
0 12326 7 1 2 12322 12325
0 12327 5 1 1 12326
0 12328 7 1 2 72702 12327
0 12329 5 1 1 12328
0 12330 7 1 2 12320 12329
0 12331 5 1 1 12330
0 12332 7 1 2 61461 12331
0 12333 5 1 1 12332
0 12334 7 1 2 62906 12333
0 12335 7 1 2 12312 12334
0 12336 5 1 1 12335
0 12337 7 1 2 12283 12336
0 12338 5 1 1 12337
0 12339 7 1 2 65366 12338
0 12340 5 1 1 12339
0 12341 7 1 2 63367 12340
0 12342 7 1 2 12235 12341
0 12343 5 1 1 12342
0 12344 7 1 2 12177 12343
0 12345 5 1 1 12344
0 12346 7 1 2 63943 12345
0 12347 5 1 1 12346
0 12348 7 2 2 81908 78989
0 12349 7 3 2 81268 79532
0 12350 7 4 2 63686 83092
0 12351 7 1 2 88267 88270
0 12352 7 1 2 88265 12351
0 12353 7 1 2 88048 12352
0 12354 5 1 1 12353
0 12355 7 1 2 12347 12354
0 12356 5 1 1 12355
0 12357 7 1 2 86779 12356
0 12358 5 1 1 12357
0 12359 7 1 2 12123 12358
0 12360 7 1 2 12083 12359
0 12361 5 1 1 12360
0 12362 7 1 2 76358 12361
0 12363 5 1 1 12362
0 12364 7 2 2 66426 85831
0 12365 5 1 1 88274
0 12366 7 1 2 87165 87537
0 12367 7 1 2 88275 12366
0 12368 5 1 1 12367
0 12369 7 1 2 84735 87259
0 12370 7 2 2 77157 12369
0 12371 7 1 2 87452 87415
0 12372 7 1 2 88276 12371
0 12373 5 1 1 12372
0 12374 7 1 2 12368 12373
0 12375 5 1 1 12374
0 12376 7 1 2 80405 12375
0 12377 5 1 1 12376
0 12378 7 1 2 72703 87533
0 12379 5 1 1 12378
0 12380 7 3 2 64466 75188
0 12381 5 2 1 88278
0 12382 7 1 2 88277 88279
0 12383 5 1 1 12382
0 12384 7 1 2 12379 12383
0 12385 5 1 1 12384
0 12386 7 1 2 66205 87503
0 12387 7 1 2 12385 12386
0 12388 5 1 1 12387
0 12389 7 1 2 12377 12388
0 12390 5 1 1 12389
0 12391 7 1 2 63687 12390
0 12392 5 1 1 12391
0 12393 7 1 2 80829 84817
0 12394 7 1 2 87504 12393
0 12395 7 1 2 88174 12394
0 12396 5 1 1 12395
0 12397 7 1 2 12392 12396
0 12398 5 1 1 12397
0 12399 7 1 2 77273 12398
0 12400 5 1 1 12399
0 12401 7 1 2 68975 12400
0 12402 7 1 2 12363 12401
0 12403 7 1 2 11918 12402
0 12404 7 1 2 10381 12403
0 12405 7 1 2 9454 12404
0 12406 7 1 2 7667 12405
0 12407 7 1 2 3184 12406
0 12408 5 1 1 12407
0 12409 7 4 2 64467 85816
0 12410 5 1 1 88283
0 12411 7 1 2 70515 69734
0 12412 7 1 2 88284 12411
0 12413 5 1 1 12412
0 12414 7 1 2 78907 12413
0 12415 5 1 1 12414
0 12416 7 1 2 62552 12415
0 12417 5 1 1 12416
0 12418 7 1 2 81676 85602
0 12419 5 1 1 12418
0 12420 7 1 2 78908 12419
0 12421 5 1 1 12420
0 12422 7 1 2 71759 12421
0 12423 5 1 1 12422
0 12424 7 1 2 12417 12423
0 12425 5 1 1 12424
0 12426 7 1 2 70758 12425
0 12427 5 1 1 12426
0 12428 7 3 2 65829 76525
0 12429 5 3 1 88287
0 12430 7 1 2 84026 88288
0 12431 5 1 1 12430
0 12432 7 1 2 5924 12431
0 12433 5 1 1 12432
0 12434 7 1 2 71534 12433
0 12435 5 1 1 12434
0 12436 7 2 2 62907 78827
0 12437 5 2 1 88293
0 12438 7 4 2 67911 71535
0 12439 5 1 1 88297
0 12440 7 1 2 73202 88298
0 12441 5 1 1 12440
0 12442 7 1 2 88295 12441
0 12443 5 1 1 12442
0 12444 7 1 2 62265 12443
0 12445 5 1 1 12444
0 12446 7 1 2 74781 88299
0 12447 5 1 1 12446
0 12448 7 1 2 12445 12447
0 12449 5 1 1 12448
0 12450 7 1 2 71760 12449
0 12451 5 1 1 12450
0 12452 7 1 2 12435 12451
0 12453 5 1 1 12452
0 12454 7 1 2 62553 12453
0 12455 5 1 1 12454
0 12456 7 1 2 12427 12455
0 12457 5 1 1 12456
0 12458 7 1 2 72291 12457
0 12459 5 1 1 12458
0 12460 7 2 2 72435 87458
0 12461 5 1 1 88301
0 12462 7 1 2 65830 88302
0 12463 5 1 1 12462
0 12464 7 1 2 60271 12463
0 12465 5 1 1 12464
0 12466 7 1 2 64928 12465
0 12467 5 1 1 12466
0 12468 7 1 2 70045 72444
0 12469 5 2 1 12468
0 12470 7 2 2 65831 71536
0 12471 7 2 2 69978 88305
0 12472 5 1 1 88307
0 12473 7 1 2 88303 12472
0 12474 5 1 1 12473
0 12475 7 1 2 64468 12474
0 12476 5 1 1 12475
0 12477 7 1 2 12467 12476
0 12478 5 1 1 12477
0 12479 7 1 2 71091 12478
0 12480 5 1 1 12479
0 12481 7 3 2 66206 73516
0 12482 5 1 1 88309
0 12483 7 1 2 77534 88310
0 12484 5 1 1 12483
0 12485 7 1 2 12480 12484
0 12486 5 1 1 12485
0 12487 7 1 2 67912 12486
0 12488 5 1 1 12487
0 12489 7 1 2 67913 76738
0 12490 5 2 1 12489
0 12491 7 1 2 77514 78828
0 12492 5 1 1 12491
0 12493 7 1 2 88312 12492
0 12494 5 1 1 12493
0 12495 7 1 2 69635 12494
0 12496 5 1 1 12495
0 12497 7 2 2 71537 87355
0 12498 5 1 1 88314
0 12499 7 1 2 62266 82132
0 12500 7 1 2 88315 12499
0 12501 5 1 1 12500
0 12502 7 1 2 12496 12501
0 12503 5 1 1 12502
0 12504 7 1 2 62063 12503
0 12505 5 1 1 12504
0 12506 7 1 2 62908 6429
0 12507 5 1 1 12506
0 12508 7 1 2 69786 2715
0 12509 7 1 2 12507 12508
0 12510 5 1 1 12509
0 12511 7 1 2 85561 12510
0 12512 5 1 1 12511
0 12513 7 1 2 70759 12512
0 12514 5 1 1 12513
0 12515 7 1 2 12505 12514
0 12516 5 1 1 12515
0 12517 7 1 2 78653 12516
0 12518 5 1 1 12517
0 12519 7 5 2 62267 76838
0 12520 7 1 2 85332 88316
0 12521 5 1 1 12520
0 12522 7 1 2 86565 12521
0 12523 5 1 1 12522
0 12524 7 1 2 77182 12523
0 12525 5 1 1 12524
0 12526 7 1 2 87948 12439
0 12527 5 1 1 12526
0 12528 7 1 2 73890 78526
0 12529 7 1 2 12527 12528
0 12530 5 1 1 12529
0 12531 7 1 2 12525 12530
0 12532 5 1 1 12531
0 12533 7 1 2 69636 12532
0 12534 5 1 1 12533
0 12535 7 1 2 80313 87350
0 12536 5 1 1 12535
0 12537 7 1 2 62909 83654
0 12538 5 1 1 12537
0 12539 7 1 2 12536 12538
0 12540 5 1 1 12539
0 12541 7 1 2 70760 12540
0 12542 5 1 1 12541
0 12543 7 1 2 12534 12542
0 12544 7 1 2 12518 12543
0 12545 7 4 2 64469 79184
0 12546 5 1 1 88321
0 12547 7 1 2 78697 88322
0 12548 5 1 1 12547
0 12549 7 1 2 87380 12548
0 12550 5 1 1 12549
0 12551 7 1 2 69787 12550
0 12552 5 1 1 12551
0 12553 7 2 2 64929 82938
0 12554 7 1 2 78357 85567
0 12555 7 1 2 88325 12554
0 12556 5 1 1 12555
0 12557 7 1 2 12552 12556
0 12558 5 1 1 12557
0 12559 7 1 2 71092 12558
0 12560 5 1 1 12559
0 12561 7 1 2 82939 82379
0 12562 7 1 2 75804 12561
0 12563 5 1 1 12562
0 12564 7 4 2 64930 65832
0 12565 5 1 1 88327
0 12566 7 4 2 64470 88328
0 12567 5 3 1 88331
0 12568 7 1 2 82369 88335
0 12569 5 1 1 12568
0 12570 7 1 2 71303 77396
0 12571 5 1 1 12570
0 12572 7 1 2 12569 12571
0 12573 7 1 2 12563 12572
0 12574 5 1 1 12573
0 12575 7 1 2 65140 12574
0 12576 5 1 1 12575
0 12577 7 1 2 12560 12576
0 12578 5 1 1 12577
0 12579 7 1 2 62554 12578
0 12580 5 1 1 12579
0 12581 7 1 2 83859 78905
0 12582 7 1 2 76545 12581
0 12583 5 1 1 12582
0 12584 7 7 2 62910 75093
0 12585 7 1 2 71761 88338
0 12586 5 1 1 12585
0 12587 7 1 2 78909 12586
0 12588 5 1 1 12587
0 12589 7 1 2 66207 12588
0 12590 5 1 1 12589
0 12591 7 2 2 66208 82861
0 12592 5 1 1 88345
0 12593 7 1 2 67914 77527
0 12594 5 1 1 12593
0 12595 7 1 2 12592 12594
0 12596 5 1 1 12595
0 12597 7 1 2 64245 12596
0 12598 5 1 1 12597
0 12599 7 1 2 82671 79178
0 12600 5 2 1 12599
0 12601 7 1 2 78552 88347
0 12602 5 1 1 12601
0 12603 7 1 2 12598 12602
0 12604 5 1 1 12603
0 12605 7 1 2 62555 12604
0 12606 5 1 1 12605
0 12607 7 1 2 12590 12606
0 12608 7 1 2 12583 12607
0 12609 5 1 1 12608
0 12610 7 1 2 72704 12609
0 12611 5 1 1 12610
0 12612 7 1 2 12580 12611
0 12613 7 1 2 12544 12612
0 12614 7 1 2 12488 12613
0 12615 7 1 2 12459 12614
0 12616 5 1 1 12615
0 12617 7 1 2 63368 12616
0 12618 5 1 1 12617
0 12619 7 2 2 75062 87425
0 12620 5 1 1 88349
0 12621 7 4 2 76908 70761
0 12622 5 1 1 88351
0 12623 7 1 2 72631 88352
0 12624 5 1 1 12623
0 12625 7 9 2 72292 74763
0 12626 5 5 1 88355
0 12627 7 1 2 70135 88364
0 12628 5 1 1 12627
0 12629 7 2 2 70762 12628
0 12630 5 2 1 88369
0 12631 7 1 2 12624 88371
0 12632 5 1 1 12631
0 12633 7 1 2 88350 12632
0 12634 5 1 1 12633
0 12635 7 1 2 61462 12634
0 12636 7 1 2 12618 12635
0 12637 5 1 1 12636
0 12638 7 1 2 65141 86026
0 12639 5 1 1 12638
0 12640 7 1 2 77422 76839
0 12641 7 1 2 74459 12640
0 12642 5 1 1 12641
0 12643 7 1 2 12639 12642
0 12644 5 1 1 12643
0 12645 7 1 2 72900 12644
0 12646 5 1 1 12645
0 12647 7 1 2 65142 88336
0 12648 5 1 1 12647
0 12649 7 2 2 74276 72637
0 12650 5 1 1 88373
0 12651 7 1 2 82528 73317
0 12652 5 2 1 12651
0 12653 7 1 2 64931 88375
0 12654 5 1 1 12653
0 12655 7 2 2 69637 69062
0 12656 5 3 1 88377
0 12657 7 2 2 64471 87689
0 12658 5 2 1 88382
0 12659 7 1 2 62268 73064
0 12660 5 1 1 12659
0 12661 7 1 2 59297 12660
0 12662 5 2 1 12661
0 12663 7 1 2 88383 88386
0 12664 5 1 1 12663
0 12665 7 1 2 88379 12664
0 12666 5 1 1 12665
0 12667 7 1 2 72293 12666
0 12668 5 1 1 12667
0 12669 7 1 2 72566 69173
0 12670 5 9 1 12669
0 12671 7 1 2 71093 88388
0 12672 5 1 1 12671
0 12673 7 2 2 12668 12672
0 12674 5 1 1 88397
0 12675 7 1 2 12654 88398
0 12676 5 1 1 12675
0 12677 7 1 2 67026 12676
0 12678 5 1 1 12677
0 12679 7 1 2 12650 12678
0 12680 5 1 1 12679
0 12681 7 1 2 62556 12680
0 12682 5 1 1 12681
0 12683 7 1 2 12648 12682
0 12684 5 1 1 12683
0 12685 7 1 2 61253 12684
0 12686 5 1 1 12685
0 12687 7 3 2 61018 81561
0 12688 5 3 1 88399
0 12689 7 2 2 74163 88400
0 12690 5 2 1 88405
0 12691 7 1 2 71450 88407
0 12692 5 1 1 12691
0 12693 7 1 2 71762 88036
0 12694 5 2 1 12693
0 12695 7 9 2 62557 72294
0 12696 5 8 1 88411
0 12697 7 1 2 74517 78114
0 12698 7 1 2 88420 12697
0 12699 7 1 2 7515 12698
0 12700 7 1 2 88409 12699
0 12701 7 1 2 12692 12700
0 12702 5 1 1 12701
0 12703 7 1 2 66209 12702
0 12704 5 1 1 12703
0 12705 7 3 2 61254 76198
0 12706 5 2 1 88428
0 12707 7 1 2 72705 88431
0 12708 5 1 1 12707
0 12709 7 2 2 65699 78654
0 12710 5 1 1 88433
0 12711 7 1 2 64246 88434
0 12712 5 1 1 12711
0 12713 7 1 2 72627 12712
0 12714 5 1 1 12713
0 12715 7 1 2 85417 12714
0 12716 5 1 1 12715
0 12717 7 1 2 12708 12716
0 12718 7 1 2 12704 12717
0 12719 5 1 1 12718
0 12720 7 1 2 60272 12719
0 12721 5 1 1 12720
0 12722 7 1 2 12686 12721
0 12723 5 1 1 12722
0 12724 7 1 2 67915 12723
0 12725 5 1 1 12724
0 12726 7 1 2 12646 12725
0 12727 5 1 1 12726
0 12728 7 1 2 63369 12727
0 12729 5 1 1 12728
0 12730 7 2 2 67528 76727
0 12731 5 4 1 88435
0 12732 7 2 2 69638 88437
0 12733 5 1 1 88441
0 12734 7 1 2 77277 12733
0 12735 5 1 1 12734
0 12736 7 1 2 62269 12735
0 12737 5 1 1 12736
0 12738 7 1 2 76359 88045
0 12739 5 1 1 12738
0 12740 7 1 2 80442 83682
0 12741 5 1 1 12740
0 12742 7 1 2 62558 12741
0 12743 5 1 1 12742
0 12744 7 1 2 12739 12743
0 12745 7 3 2 12737 12744
0 12746 5 1 1 88443
0 12747 7 6 2 71167 88421
0 12748 7 4 2 69399 74436
0 12749 5 27 1 88452
0 12750 7 2 2 71763 88456
0 12751 5 1 1 88483
0 12752 7 3 2 72082 12751
0 12753 5 3 1 88485
0 12754 7 1 2 69898 79978
0 12755 5 5 1 12754
0 12756 7 1 2 62270 88491
0 12757 5 1 1 12756
0 12758 7 1 2 88486 12757
0 12759 5 2 1 12758
0 12760 7 1 2 72295 88496
0 12761 5 2 1 12760
0 12762 7 1 2 88446 88498
0 12763 7 1 2 88444 12762
0 12764 5 1 1 12763
0 12765 7 1 2 70763 12764
0 12766 5 1 1 12765
0 12767 7 2 2 70136 12766
0 12768 5 1 1 88500
0 12769 7 1 2 65143 12768
0 12770 5 1 1 12769
0 12771 7 1 2 75980 76976
0 12772 5 1 1 12771
0 12773 7 3 2 78894 12772
0 12774 5 7 1 88502
0 12775 7 2 2 73076 88505
0 12776 5 1 1 88512
0 12777 7 3 2 65700 73347
0 12778 5 5 1 88514
0 12779 7 2 2 61019 88517
0 12780 5 1 1 88522
0 12781 7 2 2 64247 12780
0 12782 5 1 1 88524
0 12783 7 1 2 77234 78527
0 12784 5 1 1 12783
0 12785 7 1 2 59827 12784
0 12786 5 1 1 12785
0 12787 7 1 2 88525 12786
0 12788 5 1 1 12787
0 12789 7 1 2 65978 73295
0 12790 5 1 1 12789
0 12791 7 1 2 12788 12790
0 12792 5 1 1 12791
0 12793 7 1 2 69230 12792
0 12794 5 1 1 12793
0 12795 7 3 2 81564 73979
0 12796 7 4 2 72296 88526
0 12797 5 1 1 88529
0 12798 7 1 2 73247 88530
0 12799 5 1 1 12798
0 12800 7 1 2 85796 12799
0 12801 7 1 2 12794 12800
0 12802 5 2 1 12801
0 12803 7 1 2 62559 88533
0 12804 5 1 1 12803
0 12805 7 3 2 12776 12804
0 12806 5 1 1 88535
0 12807 7 1 2 12770 88536
0 12808 5 1 1 12807
0 12809 7 7 2 68281 71538
0 12810 5 1 1 88538
0 12811 7 1 2 67916 88539
0 12812 7 1 2 12808 12811
0 12813 5 1 1 12812
0 12814 7 1 2 72640 78829
0 12815 5 1 1 12814
0 12816 7 4 2 64472 71028
0 12817 5 1 1 88545
0 12818 7 1 2 71539 12817
0 12819 5 1 1 12818
0 12820 7 1 2 62271 12819
0 12821 7 1 2 12815 12820
0 12822 5 1 1 12821
0 12823 7 2 2 69788 72297
0 12824 5 2 1 88549
0 12825 7 1 2 74764 88550
0 12826 5 1 1 12825
0 12827 7 1 2 74617 12826
0 12828 5 1 1 12827
0 12829 7 1 2 70764 12828
0 12830 5 1 1 12829
0 12831 7 2 2 72567 72205
0 12832 5 3 1 88553
0 12833 7 1 2 71540 88555
0 12834 5 1 1 12833
0 12835 7 1 2 67253 86293
0 12836 7 1 2 12834 12835
0 12837 7 1 2 12830 12836
0 12838 5 1 1 12837
0 12839 7 1 2 68282 12838
0 12840 7 1 2 12822 12839
0 12841 5 1 1 12840
0 12842 7 2 2 77031 71440
0 12843 5 3 1 88558
0 12844 7 2 2 60273 75433
0 12845 5 1 1 88563
0 12846 7 1 2 88560 88564
0 12847 5 1 1 12846
0 12848 7 4 2 68283 69639
0 12849 7 5 2 65833 70765
0 12850 5 1 1 88569
0 12851 7 2 2 80124 88570
0 12852 5 1 1 88574
0 12853 7 1 2 73517 78830
0 12854 5 1 1 12853
0 12855 7 1 2 12852 12854
0 12856 5 1 1 12855
0 12857 7 1 2 72298 12856
0 12858 5 1 1 12857
0 12859 7 2 2 77175 78504
0 12860 5 7 1 88576
0 12861 7 1 2 67254 88578
0 12862 5 1 1 12861
0 12863 7 1 2 12858 12862
0 12864 5 1 1 12863
0 12865 7 1 2 88565 12864
0 12866 5 1 1 12865
0 12867 7 3 2 61020 70230
0 12868 5 2 1 88585
0 12869 7 3 2 76739 88588
0 12870 5 2 1 88590
0 12871 7 1 2 63370 79115
0 12872 7 1 2 88593 12871
0 12873 5 1 1 12872
0 12874 7 1 2 12866 12873
0 12875 5 1 1 12874
0 12876 7 1 2 62064 12875
0 12877 5 1 1 12876
0 12878 7 1 2 12847 12877
0 12879 7 1 2 12841 12878
0 12880 5 1 1 12879
0 12881 7 1 2 62560 12880
0 12882 5 1 1 12881
0 12883 7 4 2 71693 72206
0 12884 5 1 1 88595
0 12885 7 1 2 75434 73769
0 12886 7 1 2 88596 12885
0 12887 5 1 1 12886
0 12888 7 1 2 62272 87775
0 12889 5 1 1 12888
0 12890 7 1 2 12887 12889
0 12891 5 1 1 12890
0 12892 7 1 2 69506 12891
0 12893 5 1 1 12892
0 12894 7 2 2 65144 80806
0 12895 5 2 1 88599
0 12896 7 18 2 61021 73403
0 12897 7 1 2 75435 88603
0 12898 5 1 1 12897
0 12899 7 1 2 88601 12898
0 12900 5 1 1 12899
0 12901 7 1 2 66210 12900
0 12902 5 1 1 12901
0 12903 7 1 2 88602 12845
0 12904 5 1 1 12903
0 12905 7 1 2 64932 12904
0 12906 5 1 1 12905
0 12907 7 1 2 12902 12906
0 12908 7 1 2 12893 12907
0 12909 7 1 2 12882 12908
0 12910 5 1 1 12909
0 12911 7 1 2 62911 12910
0 12912 5 1 1 12911
0 12913 7 1 2 66427 12912
0 12914 7 1 2 12813 12913
0 12915 7 1 2 12729 12914
0 12916 5 1 1 12915
0 12917 7 1 2 12637 12916
0 12918 5 1 1 12917
0 12919 7 1 2 64248 82974
0 12920 5 2 1 12919
0 12921 7 1 2 85228 88621
0 12922 5 1 1 12921
0 12923 7 1 2 88356 12922
0 12924 5 1 1 12923
0 12925 7 1 2 71094 85333
0 12926 5 1 1 12925
0 12927 7 1 2 88622 12926
0 12928 5 1 1 12927
0 12929 7 1 2 66211 12928
0 12930 5 1 1 12929
0 12931 7 1 2 12924 12930
0 12932 5 1 1 12931
0 12933 7 1 2 70308 12932
0 12934 5 1 1 12933
0 12935 7 1 2 77687 82975
0 12936 5 1 1 12935
0 12937 7 7 2 59477 71168
0 12938 5 4 1 88623
0 12939 7 3 2 67255 71169
0 12940 5 1 1 88634
0 12941 7 2 2 88630 12940
0 12942 5 1 1 88637
0 12943 7 4 2 72299 88638
0 12944 5 1 1 88639
0 12945 7 1 2 87361 88640
0 12946 5 1 1 12945
0 12947 7 1 2 12936 12946
0 12948 5 1 1 12947
0 12949 7 1 2 70365 12948
0 12950 5 1 1 12949
0 12951 7 7 2 61022 76492
0 12952 5 1 1 88643
0 12953 7 1 2 82976 12952
0 12954 5 1 1 12953
0 12955 7 1 2 82569 78680
0 12956 5 1 1 12955
0 12957 7 1 2 12954 12956
0 12958 5 1 1 12957
0 12959 7 1 2 66212 12958
0 12960 5 1 1 12959
0 12961 7 1 2 78714 87466
0 12962 7 1 2 80067 12961
0 12963 7 1 2 61023 72790
0 12964 5 7 1 12963
0 12965 7 1 2 72621 78115
0 12966 5 2 1 12965
0 12967 7 1 2 88650 88657
0 12968 7 1 2 12962 12967
0 12969 5 1 1 12968
0 12970 7 1 2 12960 12969
0 12971 7 1 2 12950 12970
0 12972 7 1 2 12934 12971
0 12973 5 1 1 12972
0 12974 7 1 2 62561 12973
0 12975 5 1 1 12974
0 12976 7 2 2 71095 78029
0 12977 5 1 1 88659
0 12978 7 1 2 67917 88660
0 12979 7 1 2 88506 12978
0 12980 5 1 1 12979
0 12981 7 1 2 12975 12980
0 12982 5 1 1 12981
0 12983 7 1 2 64933 12982
0 12984 5 1 1 12983
0 12985 7 1 2 71319 88357
0 12986 5 1 1 12985
0 12987 7 1 2 74618 12986
0 12988 5 1 1 12987
0 12989 7 1 2 74402 78553
0 12990 7 1 2 12988 12989
0 12991 5 1 1 12990
0 12992 7 1 2 12984 12991
0 12993 5 1 1 12992
0 12994 7 1 2 75063 12993
0 12995 5 1 1 12994
0 12996 7 2 2 64934 74054
0 12997 5 1 1 88661
0 12998 7 1 2 62065 12997
0 12999 5 1 1 12998
0 13000 7 2 2 72083 82635
0 13001 5 1 1 88663
0 13002 7 1 2 59298 88664
0 13003 5 1 1 13002
0 13004 7 1 2 12999 13003
0 13005 5 1 1 13004
0 13006 7 1 2 73161 13005
0 13007 5 1 1 13006
0 13008 7 2 2 66213 79983
0 13009 5 2 1 88665
0 13010 7 1 2 65145 88667
0 13011 5 1 1 13010
0 13012 7 1 2 13007 13011
0 13013 5 1 1 13012
0 13014 7 1 2 67918 13013
0 13015 5 1 1 13014
0 13016 7 1 2 62066 76758
0 13017 5 1 1 13016
0 13018 7 3 2 72084 83683
0 13019 5 1 1 88669
0 13020 7 1 2 67027 88670
0 13021 5 2 1 13020
0 13022 7 2 2 74055 88672
0 13023 5 1 1 88674
0 13024 7 1 2 70137 73037
0 13025 7 1 2 13023 13024
0 13026 5 1 1 13025
0 13027 7 1 2 13017 13026
0 13028 5 2 1 13027
0 13029 7 1 2 77462 88676
0 13030 5 1 1 13029
0 13031 7 1 2 13015 13030
0 13032 5 1 1 13031
0 13033 7 1 2 63371 13032
0 13034 5 1 1 13033
0 13035 7 1 2 13034 12620
0 13036 5 1 1 13035
0 13037 7 1 2 66428 13036
0 13038 5 1 1 13037
0 13039 7 2 2 71003 83897
0 13040 5 1 1 88678
0 13041 7 1 2 81738 88679
0 13042 5 1 1 13041
0 13043 7 1 2 13038 13042
0 13044 5 1 1 13043
0 13045 7 1 2 71170 13044
0 13046 5 1 1 13045
0 13047 7 1 2 12995 13046
0 13048 7 1 2 12918 13047
0 13049 5 1 1 13048
0 13050 7 1 2 80845 13049
0 13051 5 1 1 13050
0 13052 7 1 2 78486 86027
0 13053 5 1 1 13052
0 13054 7 2 2 60886 82955
0 13055 7 1 2 69507 88680
0 13056 5 1 1 13055
0 13057 7 1 2 13053 13056
0 13058 5 1 1 13057
0 13059 7 1 2 67529 13058
0 13060 5 1 1 13059
0 13061 7 3 2 65834 70482
0 13062 5 4 1 88682
0 13063 7 1 2 82920 88685
0 13064 5 1 1 13063
0 13065 7 1 2 13060 13064
0 13066 5 1 1 13065
0 13067 7 1 2 59478 13066
0 13068 5 1 1 13067
0 13069 7 4 2 69462 78367
0 13070 5 2 1 88689
0 13071 7 1 2 73186 88690
0 13072 5 1 1 13071
0 13073 7 2 2 67919 69099
0 13074 5 3 1 88695
0 13075 7 1 2 69508 83803
0 13076 5 2 1 13075
0 13077 7 1 2 88697 88700
0 13078 5 1 1 13077
0 13079 7 1 2 67028 13078
0 13080 5 1 1 13079
0 13081 7 3 2 67920 69297
0 13082 5 1 1 88702
0 13083 7 1 2 13080 13082
0 13084 5 1 1 13083
0 13085 7 1 2 61255 13084
0 13086 5 1 1 13085
0 13087 7 1 2 13072 13086
0 13088 7 1 2 13068 13087
0 13089 5 1 1 13088
0 13090 7 1 2 61024 13089
0 13091 5 1 1 13090
0 13092 7 1 2 62067 83348
0 13093 5 3 1 13092
0 13094 7 2 2 62562 77047
0 13095 5 4 1 88708
0 13096 7 6 2 88705 88710
0 13097 7 1 2 69100 88714
0 13098 5 1 1 13097
0 13099 7 1 2 69298 81613
0 13100 5 1 1 13099
0 13101 7 1 2 76324 13100
0 13102 7 1 2 13098 13101
0 13103 5 1 1 13102
0 13104 7 1 2 82921 13103
0 13105 5 1 1 13104
0 13106 7 1 2 13091 13105
0 13107 5 1 1 13106
0 13108 7 1 2 59828 13107
0 13109 5 1 1 13108
0 13110 7 1 2 73804 75816
0 13111 5 1 1 13110
0 13112 7 1 2 69640 74506
0 13113 5 4 1 13112
0 13114 7 1 2 71868 88720
0 13115 5 1 1 13114
0 13116 7 1 2 13111 13115
0 13117 5 1 1 13116
0 13118 7 1 2 67029 13117
0 13119 5 1 1 13118
0 13120 7 1 2 82560 71869
0 13121 5 1 1 13120
0 13122 7 1 2 13119 13121
0 13123 5 1 1 13122
0 13124 7 2 2 67921 13123
0 13125 5 1 1 88724
0 13126 7 1 2 61256 88725
0 13127 5 1 1 13126
0 13128 7 1 2 13109 13127
0 13129 5 1 1 13128
0 13130 7 1 2 60087 13129
0 13131 5 1 1 13130
0 13132 7 2 2 67030 75817
0 13133 7 3 2 59829 84797
0 13134 5 3 1 88728
0 13135 7 1 2 73910 88729
0 13136 7 1 2 88726 13135
0 13137 5 1 1 13136
0 13138 7 1 2 13131 13137
0 13139 5 1 1 13138
0 13140 7 6 2 60274 83696
0 13141 5 3 1 88734
0 13142 7 1 2 79433 88735
0 13143 7 1 2 13139 13142
0 13144 5 1 1 13143
0 13145 7 1 2 64473 72844
0 13146 5 1 1 13145
0 13147 7 1 2 76728 13146
0 13148 5 5 1 13147
0 13149 7 1 2 72300 88743
0 13150 5 2 1 13149
0 13151 7 7 2 69509 71694
0 13152 5 4 1 88750
0 13153 7 1 2 72489 88757
0 13154 5 1 1 13153
0 13155 7 1 2 62068 72706
0 13156 5 1 1 13155
0 13157 7 1 2 13154 13156
0 13158 7 1 2 88748 13157
0 13159 5 1 1 13158
0 13160 7 1 2 79052 13159
0 13161 5 1 1 13160
0 13162 7 3 2 65835 76238
0 13163 5 9 1 88761
0 13164 7 1 2 77372 88764
0 13165 5 1 1 13164
0 13166 7 1 2 76459 77397
0 13167 5 1 1 13166
0 13168 7 1 2 13165 13167
0 13169 5 1 1 13168
0 13170 7 1 2 72901 13169
0 13171 5 1 1 13170
0 13172 7 1 2 69510 71850
0 13173 5 1 1 13172
0 13174 7 1 2 72490 13173
0 13175 7 1 2 88604 88765
0 13176 5 1 1 13175
0 13177 7 1 2 78003 76239
0 13178 5 1 1 13177
0 13179 7 1 2 60275 13178
0 13180 5 1 1 13179
0 13181 7 1 2 13176 13180
0 13182 7 1 2 13174 13181
0 13183 5 1 1 13182
0 13184 7 1 2 62912 13183
0 13185 5 1 1 13184
0 13186 7 1 2 13171 13185
0 13187 7 1 2 13161 13186
0 13188 5 1 1 13187
0 13189 7 1 2 62563 13188
0 13190 5 1 1 13189
0 13191 7 3 2 67530 82832
0 13192 5 1 1 88773
0 13193 7 1 2 61025 80061
0 13194 5 1 1 13193
0 13195 7 1 2 64474 13194
0 13196 5 1 1 13195
0 13197 7 1 2 72791 72207
0 13198 5 2 1 13197
0 13199 7 1 2 65979 80078
0 13200 5 3 1 13199
0 13201 7 2 2 59299 88778
0 13202 5 1 1 88781
0 13203 7 1 2 80087 88782
0 13204 5 1 1 13203
0 13205 7 2 2 88776 13204
0 13206 5 1 1 88783
0 13207 7 1 2 13196 13206
0 13208 5 1 1 13207
0 13209 7 1 2 88774 13208
0 13210 5 1 1 13209
0 13211 7 2 2 72301 88492
0 13212 5 1 1 88785
0 13213 7 1 2 88503 13212
0 13214 5 2 1 13213
0 13215 7 2 2 61257 77026
0 13216 5 1 1 88789
0 13217 7 2 2 77978 13216
0 13218 7 1 2 88787 88791
0 13219 5 1 1 13218
0 13220 7 1 2 74239 88507
0 13221 5 1 1 13220
0 13222 7 1 2 13219 13221
0 13223 5 1 1 13222
0 13224 7 1 2 67922 13223
0 13225 5 1 1 13224
0 13226 7 1 2 13210 13225
0 13227 7 1 2 13190 13226
0 13228 5 1 1 13227
0 13229 7 1 2 62273 13228
0 13230 5 1 1 13229
0 13231 7 1 2 76442 72902
0 13232 5 1 1 13231
0 13233 7 1 2 72707 13232
0 13234 5 2 1 13233
0 13235 7 1 2 76401 88793
0 13236 5 1 1 13235
0 13237 7 1 2 71096 81606
0 13238 5 2 1 13237
0 13239 7 1 2 60088 88795
0 13240 5 1 1 13239
0 13241 7 2 2 60887 76550
0 13242 5 1 1 88797
0 13243 7 1 2 71615 88798
0 13244 5 2 1 13243
0 13245 7 1 2 13240 88799
0 13246 5 1 1 13245
0 13247 7 1 2 76253 13246
0 13248 5 1 1 13247
0 13249 7 1 2 13236 13248
0 13250 5 1 1 13249
0 13251 7 1 2 67531 13250
0 13252 5 1 1 13251
0 13253 7 1 2 80926 74747
0 13254 5 1 1 13253
0 13255 7 1 2 13252 13254
0 13256 5 1 1 13255
0 13257 7 1 2 66214 13256
0 13258 5 1 1 13257
0 13259 7 1 2 64475 88438
0 13260 5 1 1 13259
0 13261 7 1 2 74532 13260
0 13262 5 1 1 13261
0 13263 7 1 2 76663 13262
0 13264 5 1 1 13263
0 13265 7 1 2 82745 13264
0 13266 5 1 1 13265
0 13267 7 1 2 60276 13266
0 13268 5 1 1 13267
0 13269 7 1 2 62913 13268
0 13270 7 1 2 13258 13269
0 13271 5 1 1 13270
0 13272 7 4 2 80125 70944
0 13273 5 1 1 88801
0 13274 7 3 2 61258 72708
0 13275 7 1 2 88802 88805
0 13276 5 1 1 13275
0 13277 7 7 2 62564 71097
0 13278 5 5 1 88808
0 13279 7 1 2 74182 88815
0 13280 5 1 1 13279
0 13281 7 2 2 59830 73805
0 13282 5 4 1 88820
0 13283 7 3 2 64935 71911
0 13284 5 5 1 88826
0 13285 7 2 2 88822 88827
0 13286 5 1 1 88834
0 13287 7 1 2 13280 88835
0 13288 5 1 1 13287
0 13289 7 1 2 67256 13288
0 13290 5 1 1 13289
0 13291 7 2 2 59479 88816
0 13292 7 1 2 60888 88836
0 13293 5 2 1 13292
0 13294 7 2 2 66215 88828
0 13295 5 2 1 88840
0 13296 7 2 2 88823 88841
0 13297 5 4 1 88844
0 13298 7 1 2 88838 88845
0 13299 5 2 1 13298
0 13300 7 1 2 69511 88850
0 13301 5 1 1 13300
0 13302 7 2 2 72085 88846
0 13303 5 1 1 88852
0 13304 7 1 2 13301 13303
0 13305 7 1 2 13290 13304
0 13306 5 1 1 13305
0 13307 7 1 2 65146 13306
0 13308 5 1 1 13307
0 13309 7 1 2 13276 13308
0 13310 5 1 1 13309
0 13311 7 1 2 67031 13310
0 13312 5 1 1 13311
0 13313 7 9 2 64249 62565
0 13314 5 3 1 88854
0 13315 7 1 2 69364 88855
0 13316 5 4 1 13315
0 13317 7 2 2 61259 88866
0 13318 5 1 1 88870
0 13319 7 1 2 72709 13318
0 13320 5 1 1 13319
0 13321 7 1 2 79972 73162
0 13322 5 1 1 13321
0 13323 7 1 2 60277 13322
0 13324 7 1 2 13320 13323
0 13325 5 1 1 13324
0 13326 7 1 2 67257 88853
0 13327 5 1 1 13326
0 13328 7 1 2 71171 82763
0 13329 5 1 1 13328
0 13330 7 1 2 77984 73785
0 13331 5 2 1 13330
0 13332 7 1 2 60089 88872
0 13333 5 3 1 13332
0 13334 7 7 2 67532 72208
0 13335 5 2 1 88877
0 13336 7 5 2 61260 71695
0 13337 5 1 1 88886
0 13338 7 1 2 65147 13337
0 13339 7 1 2 88884 13338
0 13340 7 1 2 88874 13339
0 13341 7 1 2 13329 13340
0 13342 7 1 2 13327 13341
0 13343 5 1 1 13342
0 13344 7 1 2 13325 13343
0 13345 5 1 1 13344
0 13346 7 1 2 67923 768
0 13347 7 1 2 13345 13346
0 13348 7 1 2 13312 13347
0 13349 5 1 1 13348
0 13350 7 1 2 13271 13349
0 13351 5 1 1 13350
0 13352 7 4 2 67258 75708
0 13353 5 1 1 88891
0 13354 7 1 2 69641 88892
0 13355 5 1 1 13354
0 13356 7 1 2 79179 13355
0 13357 5 1 1 13356
0 13358 7 1 2 72710 13357
0 13359 5 1 1 13358
0 13360 7 1 2 78804 73203
0 13361 5 1 1 13360
0 13362 7 1 2 13359 13361
0 13363 5 1 1 13362
0 13364 7 1 2 62566 13363
0 13365 5 1 1 13364
0 13366 7 1 2 71320 72302
0 13367 7 1 2 88792 13366
0 13368 5 1 1 13367
0 13369 7 1 2 13365 13368
0 13370 5 1 1 13369
0 13371 7 1 2 67924 13370
0 13372 5 1 1 13371
0 13373 7 1 2 69735 72303
0 13374 7 1 2 88775 13373
0 13375 5 1 1 13374
0 13376 7 1 2 13372 13375
0 13377 5 1 1 13376
0 13378 7 1 2 71764 13377
0 13379 5 1 1 13378
0 13380 7 1 2 82841 88332
0 13381 5 1 1 13380
0 13382 7 1 2 67925 84909
0 13383 5 3 1 13382
0 13384 7 1 2 74782 77497
0 13385 7 1 2 88895 13384
0 13386 5 1 1 13385
0 13387 7 1 2 65836 87744
0 13388 5 1 1 13387
0 13389 7 2 2 62567 87765
0 13390 5 1 1 88898
0 13391 7 1 2 78715 88899
0 13392 5 1 1 13391
0 13393 7 1 2 13388 13392
0 13394 7 1 2 13386 13393
0 13395 5 1 1 13394
0 13396 7 1 2 60278 13395
0 13397 5 1 1 13396
0 13398 7 1 2 13381 13397
0 13399 5 1 1 13398
0 13400 7 1 2 72304 13399
0 13401 5 1 1 13400
0 13402 7 1 2 71172 73641
0 13403 5 1 1 13402
0 13404 7 1 2 72418 74645
0 13405 7 1 2 13403 13404
0 13406 5 1 1 13405
0 13407 7 1 2 72086 13406
0 13408 5 1 1 13407
0 13409 7 1 2 71173 75796
0 13410 5 1 1 13409
0 13411 7 4 2 71467 73703
0 13412 7 5 2 67533 74619
0 13413 7 1 2 88900 88904
0 13414 5 1 1 13413
0 13415 7 1 2 13410 13414
0 13416 7 1 2 13408 13415
0 13417 5 2 1 13416
0 13418 7 1 2 72817 88909
0 13419 5 1 1 13418
0 13420 7 1 2 68284 13419
0 13421 7 1 2 13401 13420
0 13422 7 1 2 13379 13421
0 13423 7 1 2 13351 13422
0 13424 7 1 2 13230 13423
0 13425 5 1 1 13424
0 13426 7 4 2 59831 82647
0 13427 5 5 1 88911
0 13428 7 1 2 78386 88915
0 13429 5 1 1 13428
0 13430 7 1 2 69512 13429
0 13431 5 1 1 13430
0 13432 7 2 2 76551 71616
0 13433 5 2 1 88920
0 13434 7 1 2 13431 88922
0 13435 5 1 1 13434
0 13436 7 1 2 67534 13435
0 13437 5 1 1 13436
0 13438 7 6 2 67926 71174
0 13439 5 9 1 88924
0 13440 7 1 2 69736 88412
0 13441 5 1 1 13440
0 13442 7 1 2 88925 13441
0 13443 5 1 1 13442
0 13444 7 1 2 13437 13443
0 13445 5 1 1 13444
0 13446 7 1 2 72087 13445
0 13447 5 2 1 13446
0 13448 7 3 2 62914 71912
0 13449 5 17 1 88941
0 13450 7 1 2 70516 88944
0 13451 5 1 1 13450
0 13452 7 3 2 67259 73806
0 13453 5 2 1 88961
0 13454 7 1 2 69719 88962
0 13455 5 1 1 13454
0 13456 7 1 2 13451 13455
0 13457 5 1 1 13456
0 13458 7 1 2 59832 13457
0 13459 5 1 1 13458
0 13460 7 1 2 62915 76597
0 13461 5 2 1 13460
0 13462 7 1 2 62069 78387
0 13463 5 2 1 13462
0 13464 7 1 2 61026 88968
0 13465 7 1 2 88966 13464
0 13466 5 1 1 13465
0 13467 7 1 2 13459 13466
0 13468 5 1 1 13467
0 13469 7 1 2 71696 13468
0 13470 5 1 1 13469
0 13471 7 1 2 88912 88967
0 13472 5 1 1 13471
0 13473 7 1 2 13470 13472
0 13474 7 1 2 88939 13473
0 13475 5 1 1 13474
0 13476 7 1 2 76759 13475
0 13477 5 1 1 13476
0 13478 7 1 2 81692 75937
0 13479 5 1 1 13478
0 13480 7 4 2 71913 88824
0 13481 7 2 2 62916 88970
0 13482 7 1 2 13479 88974
0 13483 5 1 1 13482
0 13484 7 1 2 60279 13483
0 13485 5 1 1 13484
0 13486 7 9 2 60790 82495
0 13487 5 1 1 88976
0 13488 7 1 2 71356 84798
0 13489 7 1 2 88977 13488
0 13490 5 1 1 13489
0 13491 7 1 2 13485 13490
0 13492 5 1 1 13491
0 13493 7 1 2 70138 13492
0 13494 5 1 1 13493
0 13495 7 1 2 81798 13494
0 13496 5 1 1 13495
0 13497 7 1 2 72088 13496
0 13498 5 1 1 13497
0 13499 7 1 2 60280 73006
0 13500 5 3 1 13499
0 13501 7 1 2 83050 71441
0 13502 5 1 1 13501
0 13503 7 1 2 88985 13502
0 13504 5 1 1 13503
0 13505 7 1 2 69513 13504
0 13506 5 1 1 13505
0 13507 7 12 2 59480 61027
0 13508 5 2 1 88988
0 13509 7 2 2 77113 78287
0 13510 5 3 1 89002
0 13511 7 1 2 88989 89003
0 13512 5 1 1 13511
0 13513 7 1 2 13506 13512
0 13514 5 1 1 13513
0 13515 7 1 2 67535 13514
0 13516 5 1 1 13515
0 13517 7 1 2 81624 88624
0 13518 5 1 1 13517
0 13519 7 1 2 62917 76572
0 13520 5 3 1 13519
0 13521 7 1 2 78938 79246
0 13522 7 1 2 89007 13521
0 13523 5 1 1 13522
0 13524 7 1 2 13518 13523
0 13525 5 1 1 13524
0 13526 7 1 2 60281 13525
0 13527 5 1 1 13526
0 13528 7 1 2 13516 13527
0 13529 5 1 1 13528
0 13530 7 1 2 70139 13529
0 13531 5 1 1 13530
0 13532 7 1 2 5875 88986
0 13533 5 1 1 13532
0 13534 7 1 2 69514 13533
0 13535 5 1 1 13534
0 13536 7 2 2 60282 70517
0 13537 5 1 1 89010
0 13538 7 2 2 61261 78368
0 13539 5 1 1 89012
0 13540 7 1 2 13537 13539
0 13541 5 1 1 13540
0 13542 7 1 2 67536 13541
0 13543 5 1 1 13542
0 13544 7 1 2 13535 13543
0 13545 5 1 1 13544
0 13546 7 1 2 60090 13545
0 13547 5 1 1 13546
0 13548 7 1 2 78388 83146
0 13549 5 3 1 13548
0 13550 7 2 2 67537 89014
0 13551 5 1 1 89017
0 13552 7 1 2 78270 13353
0 13553 5 2 1 13552
0 13554 7 1 2 69515 89019
0 13555 5 1 1 13554
0 13556 7 1 2 13551 13555
0 13557 5 1 1 13556
0 13558 7 1 2 60283 13557
0 13559 5 1 1 13558
0 13560 7 1 2 13547 13559
0 13561 5 1 1 13560
0 13562 7 1 2 74620 13561
0 13563 5 1 1 13562
0 13564 7 1 2 62918 78537
0 13565 5 1 1 13564
0 13566 7 1 2 81791 13565
0 13567 5 1 1 13566
0 13568 7 1 2 63372 13567
0 13569 7 1 2 13563 13568
0 13570 7 1 2 13531 13569
0 13571 7 1 2 13498 13570
0 13572 7 1 2 13477 13571
0 13573 5 1 1 13572
0 13574 7 1 2 61463 13573
0 13575 7 1 2 13425 13574
0 13576 5 1 1 13575
0 13577 7 5 2 66429 76760
0 13578 5 3 1 89021
0 13579 7 1 2 78144 71914
0 13580 5 4 1 13579
0 13581 7 1 2 69516 89029
0 13582 5 1 1 13581
0 13583 7 1 2 8142 13582
0 13584 5 1 1 13583
0 13585 7 1 2 60889 13584
0 13586 5 1 1 13585
0 13587 7 3 2 67260 88945
0 13588 5 1 1 89033
0 13589 7 1 2 69720 89034
0 13590 5 1 1 13589
0 13591 7 1 2 13586 13590
0 13592 5 1 1 13591
0 13593 7 1 2 59481 13592
0 13594 5 1 1 13593
0 13595 7 1 2 73807 88686
0 13596 5 1 1 13595
0 13597 7 1 2 81607 13596
0 13598 5 1 1 13597
0 13599 7 1 2 59482 13598
0 13600 5 1 1 13599
0 13601 7 1 2 62568 75756
0 13602 5 2 1 13601
0 13603 7 4 2 71595 89036
0 13604 5 1 1 89038
0 13605 7 1 2 13600 13604
0 13606 5 1 1 13605
0 13607 7 1 2 67927 13606
0 13608 5 1 1 13607
0 13609 7 6 2 67928 73808
0 13610 5 7 1 89042
0 13611 7 1 2 88380 89043
0 13612 5 1 1 13611
0 13613 7 8 2 60890 69517
0 13614 5 4 1 89055
0 13615 7 1 2 89056 89035
0 13616 5 1 1 13615
0 13617 7 1 2 13612 13616
0 13618 5 1 1 13617
0 13619 7 1 2 67032 13618
0 13620 5 1 1 13619
0 13621 7 1 2 13608 13620
0 13622 7 1 2 13594 13621
0 13623 5 1 1 13622
0 13624 7 1 2 59833 13623
0 13625 5 1 1 13624
0 13626 7 1 2 13125 13625
0 13627 5 1 1 13626
0 13628 7 1 2 89022 13627
0 13629 5 1 1 13628
0 13630 7 1 2 69642 85097
0 13631 5 1 1 13630
0 13632 7 1 2 87426 13631
0 13633 5 1 1 13632
0 13634 7 1 2 82423 13633
0 13635 5 1 1 13634
0 13636 7 1 2 81792 13635
0 13637 5 1 1 13636
0 13638 7 1 2 13629 13637
0 13639 5 1 1 13638
0 13640 7 1 2 68285 13639
0 13641 5 1 1 13640
0 13642 7 1 2 66430 88910
0 13643 5 1 1 13642
0 13644 7 5 2 72089 76630
0 13645 5 2 1 89067
0 13646 7 1 2 78442 89068
0 13647 5 1 1 13646
0 13648 7 1 2 69518 87427
0 13649 7 1 2 75775 13648
0 13650 5 1 1 13649
0 13651 7 1 2 13647 13650
0 13652 7 1 2 13643 13651
0 13653 5 1 1 13652
0 13654 7 1 2 69042 13653
0 13655 5 1 1 13654
0 13656 7 2 2 68286 75874
0 13657 5 1 1 89074
0 13658 7 1 2 79948 83411
0 13659 5 1 1 13658
0 13660 7 2 2 67538 13659
0 13661 7 3 2 69519 72209
0 13662 5 1 1 89078
0 13663 7 1 2 89076 89079
0 13664 5 1 1 13663
0 13665 7 1 2 13657 13664
0 13666 5 1 1 13665
0 13667 7 1 2 59483 13666
0 13668 5 1 1 13667
0 13669 7 1 2 75829 74262
0 13670 5 2 1 13669
0 13671 7 1 2 13668 89081
0 13672 5 1 1 13671
0 13673 7 1 2 69101 13672
0 13674 5 1 1 13673
0 13675 7 1 2 69231 88809
0 13676 5 2 1 13675
0 13677 7 1 2 89075 89083
0 13678 5 1 1 13677
0 13679 7 4 2 69174 72210
0 13680 5 1 1 89085
0 13681 7 1 2 89077 89086
0 13682 5 1 1 13681
0 13683 7 1 2 89082 13682
0 13684 5 1 1 13683
0 13685 7 1 2 76254 13684
0 13686 5 1 1 13685
0 13687 7 1 2 13678 13686
0 13688 7 1 2 13674 13687
0 13689 5 1 1 13688
0 13690 7 1 2 67929 13689
0 13691 5 1 1 13690
0 13692 7 1 2 13655 13691
0 13693 5 1 1 13692
0 13694 7 1 2 70140 13693
0 13695 5 1 1 13694
0 13696 7 1 2 5276 76393
0 13697 5 1 1 13696
0 13698 7 1 2 77768 13697
0 13699 5 1 1 13698
0 13700 7 2 2 65148 82940
0 13701 5 1 1 89089
0 13702 7 1 2 88605 13701
0 13703 5 1 1 13702
0 13704 7 2 2 61262 79053
0 13705 5 1 1 89091
0 13706 7 1 2 13703 13705
0 13707 5 1 1 13706
0 13708 7 1 2 63373 13707
0 13709 5 1 1 13708
0 13710 7 1 2 13699 13709
0 13711 5 1 1 13710
0 13712 7 1 2 61464 13711
0 13713 5 1 1 13712
0 13714 7 5 2 59834 60284
0 13715 7 10 2 72940 89093
0 13716 5 1 1 89098
0 13717 7 3 2 63374 82941
0 13718 5 1 1 89108
0 13719 7 2 2 85925 13718
0 13720 7 1 2 89099 89111
0 13721 5 1 1 13720
0 13722 7 1 2 61263 81216
0 13723 5 1 1 13722
0 13724 7 1 2 60285 78980
0 13725 7 1 2 13723 13724
0 13726 5 1 1 13725
0 13727 7 2 2 65149 85926
0 13728 5 1 1 89113
0 13729 7 1 2 77979 72903
0 13730 7 1 2 13728 13729
0 13731 7 1 2 13726 13730
0 13732 5 1 1 13731
0 13733 7 1 2 13721 13732
0 13734 7 1 2 13713 13733
0 13735 5 1 1 13734
0 13736 7 1 2 76664 13735
0 13737 5 1 1 13736
0 13738 7 2 2 70592 83399
0 13739 5 1 1 89115
0 13740 7 2 2 67930 73704
0 13741 5 1 1 89117
0 13742 7 1 2 81464 13741
0 13743 5 1 1 13742
0 13744 7 1 2 71175 13743
0 13745 5 1 1 13744
0 13746 7 1 2 2295 88923
0 13747 5 1 1 13746
0 13748 7 1 2 69520 13747
0 13749 5 1 1 13748
0 13750 7 1 2 13745 13749
0 13751 5 1 1 13750
0 13752 7 1 2 67539 13751
0 13753 5 1 1 13752
0 13754 7 2 2 70518 72211
0 13755 5 2 1 89119
0 13756 7 1 2 78389 89121
0 13757 5 1 1 13756
0 13758 7 1 2 67540 13757
0 13759 5 1 1 13758
0 13760 7 1 2 70519 88926
0 13761 5 1 1 13760
0 13762 7 5 2 60791 61028
0 13763 5 1 1 89123
0 13764 7 4 2 59300 89124
0 13765 5 1 1 89128
0 13766 7 1 2 76579 89129
0 13767 5 1 1 13766
0 13768 7 1 2 13761 13767
0 13769 7 1 2 13759 13768
0 13770 5 1 1 13769
0 13771 7 1 2 71697 13770
0 13772 5 1 1 13771
0 13773 7 2 2 76552 84799
0 13774 5 3 1 89132
0 13775 7 1 2 13772 89134
0 13776 7 1 2 13753 13775
0 13777 7 1 2 88940 13776
0 13778 5 1 1 13777
0 13779 7 1 2 89116 13778
0 13780 5 1 1 13779
0 13781 7 1 2 13737 13780
0 13782 7 1 2 13695 13781
0 13783 7 1 2 13641 13782
0 13784 7 1 2 13576 13783
0 13785 5 1 1 13784
0 13786 7 1 2 81165 13785
0 13787 5 1 1 13786
0 13788 7 1 2 13144 13787
0 13789 7 1 2 13051 13788
0 13790 5 1 1 13789
0 13791 7 1 2 68849 13790
0 13792 5 1 1 13791
0 13793 7 1 2 64250 70385
0 13794 5 2 1 13793
0 13795 7 1 2 70355 89137
0 13796 7 1 2 70428 13795
0 13797 5 1 1 13796
0 13798 7 1 2 70431 13797
0 13799 5 2 1 13798
0 13800 7 1 2 65980 81465
0 13801 5 1 1 13800
0 13802 7 7 2 59301 73433
0 13803 7 2 2 76337 71617
0 13804 5 1 1 89148
0 13805 7 1 2 89141 89149
0 13806 5 2 1 13805
0 13807 7 1 2 64693 89150
0 13808 5 1 1 13807
0 13809 7 1 2 13801 13808
0 13810 7 3 2 89139 13809
0 13811 5 1 1 89152
0 13812 7 1 2 60091 89153
0 13813 5 1 1 13812
0 13814 7 1 2 60286 13813
0 13815 5 1 1 13814
0 13816 7 1 2 76394 13815
0 13817 5 1 1 13816
0 13818 7 1 2 62919 13817
0 13819 5 1 1 13818
0 13820 7 3 2 64936 69643
0 13821 5 4 1 89155
0 13822 7 4 2 64694 69644
0 13823 5 1 1 89162
0 13824 7 2 2 65981 89163
0 13825 5 2 1 89166
0 13826 7 2 2 89158 89168
0 13827 5 2 1 89170
0 13828 7 1 2 84015 89172
0 13829 5 1 1 13828
0 13830 7 1 2 72904 13829
0 13831 5 1 1 13830
0 13832 7 1 2 69232 13831
0 13833 5 1 1 13832
0 13834 7 1 2 64937 88402
0 13835 5 1 1 13834
0 13836 7 1 2 85797 13835
0 13837 5 2 1 13836
0 13838 7 1 2 82798 89174
0 13839 5 1 1 13838
0 13840 7 1 2 77168 13839
0 13841 7 1 2 13833 13840
0 13842 5 1 1 13841
0 13843 7 1 2 67931 13842
0 13844 5 1 1 13843
0 13845 7 1 2 79848 75764
0 13846 7 1 2 88766 13845
0 13847 5 1 1 13846
0 13848 7 1 2 13844 13847
0 13849 5 1 1 13848
0 13850 7 1 2 61264 13849
0 13851 5 1 1 13850
0 13852 7 1 2 76402 81443
0 13853 5 2 1 13852
0 13854 7 1 2 81460 78554
0 13855 7 1 2 89176 13854
0 13856 5 1 1 13855
0 13857 7 1 2 72905 85992
0 13858 7 1 2 13856 13857
0 13859 5 1 1 13858
0 13860 7 1 2 13851 13859
0 13861 7 1 2 13819 13860
0 13862 5 1 1 13861
0 13863 7 1 2 63375 13862
0 13864 5 1 1 13863
0 13865 7 1 2 69233 69737
0 13866 5 7 1 13865
0 13867 7 3 2 73255 89178
0 13868 7 3 2 72180 89185
0 13869 5 4 1 89188
0 13870 7 2 2 72305 89191
0 13871 5 1 1 89195
0 13872 7 1 2 71176 13871
0 13873 5 3 1 13872
0 13874 7 1 2 71541 89197
0 13875 5 1 1 13874
0 13876 7 1 2 69789 88683
0 13877 5 4 1 13876
0 13878 7 2 2 64476 70414
0 13879 5 1 1 89204
0 13880 7 1 2 70423 89205
0 13881 5 1 1 13880
0 13882 7 4 2 89200 13881
0 13883 5 5 1 89206
0 13884 7 1 2 89210 88579
0 13885 5 1 1 13884
0 13886 7 1 2 76761 13885
0 13887 7 1 2 13875 13886
0 13888 5 1 1 13887
0 13889 7 1 2 77769 13888
0 13890 5 1 1 13889
0 13891 7 1 2 13864 13890
0 13892 5 1 1 13891
0 13893 7 1 2 66431 13892
0 13894 5 1 1 13893
0 13895 7 4 2 65150 77770
0 13896 5 2 1 89215
0 13897 7 1 2 77734 89211
0 13898 5 1 1 13897
0 13899 7 1 2 70046 89198
0 13900 5 1 1 13899
0 13901 7 1 2 13898 13900
0 13902 5 1 1 13901
0 13903 7 1 2 89216 13902
0 13904 5 1 1 13903
0 13905 7 1 2 13894 13904
0 13906 5 1 1 13905
0 13907 7 1 2 68850 13906
0 13908 5 1 1 13907
0 13909 7 1 2 83738 78895
0 13910 5 1 1 13909
0 13911 7 1 2 75124 82942
0 13912 5 1 1 13911
0 13913 7 1 2 71698 75783
0 13914 7 1 2 13912 13913
0 13915 5 1 1 13914
0 13916 7 1 2 13910 13915
0 13917 5 1 1 13916
0 13918 7 1 2 60092 13917
0 13919 5 1 1 13918
0 13920 7 1 2 62920 78313
0 13921 5 1 1 13920
0 13922 7 1 2 61265 75107
0 13923 7 1 2 13921 13922
0 13924 5 1 1 13923
0 13925 7 1 2 13919 13924
0 13926 5 1 1 13925
0 13927 7 1 2 72212 13926
0 13928 5 1 1 13927
0 13929 7 4 2 75108 70593
0 13930 5 2 1 89221
0 13931 7 2 2 67932 89222
0 13932 5 1 1 89227
0 13933 7 1 2 13928 13932
0 13934 5 1 1 13933
0 13935 7 1 2 81090 13934
0 13936 5 1 1 13935
0 13937 7 1 2 71542 13811
0 13938 5 1 1 13937
0 13939 7 2 2 65982 70425
0 13940 5 3 1 89229
0 13941 7 1 2 61029 69446
0 13942 5 2 1 13941
0 13943 7 3 2 65983 70404
0 13944 5 1 1 89236
0 13945 7 1 2 60891 13944
0 13946 5 1 1 13945
0 13947 7 2 2 89234 13946
0 13948 7 1 2 64251 89239
0 13949 5 1 1 13948
0 13950 7 1 2 65984 70356
0 13951 5 1 1 13950
0 13952 7 1 2 13949 13951
0 13953 5 1 1 13952
0 13954 7 1 2 64477 13953
0 13955 5 1 1 13954
0 13956 7 1 2 89231 13955
0 13957 5 1 1 13956
0 13958 7 1 2 64695 13957
0 13959 5 1 1 13958
0 13960 7 1 2 60287 78823
0 13961 7 1 2 13959 13960
0 13962 5 1 1 13961
0 13963 7 1 2 70766 13962
0 13964 5 1 1 13963
0 13965 7 1 2 13938 13964
0 13966 5 1 1 13965
0 13967 7 3 2 68851 83093
0 13968 7 1 2 13966 89241
0 13969 5 1 1 13968
0 13970 7 1 2 13936 13969
0 13971 5 1 1 13970
0 13972 7 1 2 61465 13971
0 13973 5 1 1 13972
0 13974 7 2 2 81976 78555
0 13975 5 1 1 89244
0 13976 7 1 2 78319 89245
0 13977 5 1 1 13976
0 13978 7 5 2 81091 85895
0 13979 7 1 2 74183 83025
0 13980 5 1 1 13979
0 13981 7 6 2 60093 60792
0 13982 7 1 2 59302 89251
0 13983 7 1 2 82768 13982
0 13984 5 1 1 13983
0 13985 7 1 2 13980 13984
0 13986 5 1 1 13985
0 13987 7 1 2 89246 13986
0 13988 5 1 1 13987
0 13989 7 1 2 13977 13988
0 13990 5 1 1 13989
0 13991 7 1 2 67033 13990
0 13992 5 1 1 13991
0 13993 7 1 2 74056 82464
0 13994 5 1 1 13993
0 13995 7 1 2 60288 85065
0 13996 7 1 2 81962 13995
0 13997 7 1 2 13994 13996
0 13998 5 1 1 13997
0 13999 7 1 2 13992 13998
0 14000 5 1 1 13999
0 14001 7 1 2 71177 14000
0 14002 5 1 1 14001
0 14003 7 2 2 72667 72628
0 14004 5 1 1 89257
0 14005 7 1 2 89247 89258
0 14006 5 1 1 14005
0 14007 7 1 2 75189 80533
0 14008 7 1 2 75991 14007
0 14009 5 1 1 14008
0 14010 7 1 2 14006 14009
0 14011 5 1 1 14010
0 14012 7 1 2 78392 14011
0 14013 5 1 1 14012
0 14014 7 1 2 82625 87514
0 14015 5 1 1 14014
0 14016 7 3 2 59303 80796
0 14017 7 1 2 80534 89259
0 14018 7 1 2 88346 14017
0 14019 5 1 1 14018
0 14020 7 1 2 14015 14019
0 14021 5 1 1 14020
0 14022 7 1 2 72906 14021
0 14023 5 1 1 14022
0 14024 7 1 2 81963 89100
0 14025 5 1 1 14024
0 14026 7 1 2 72823 2470
0 14027 5 5 1 14026
0 14028 7 3 2 66432 71178
0 14029 7 1 2 80535 89267
0 14030 7 1 2 89262 14029
0 14031 5 1 1 14030
0 14032 7 1 2 14025 14031
0 14033 7 1 2 14023 14032
0 14034 5 1 1 14033
0 14035 7 1 2 75962 14034
0 14036 5 1 1 14035
0 14037 7 1 2 14013 14036
0 14038 7 1 2 14002 14037
0 14039 7 1 2 13973 14038
0 14040 7 1 2 13908 14039
0 14041 5 1 1 14040
0 14042 7 1 2 67541 14041
0 14043 5 1 1 14042
0 14044 7 1 2 81502 87515
0 14045 5 1 1 14044
0 14046 7 1 2 14045 13975
0 14047 5 1 1 14046
0 14048 7 1 2 60094 14047
0 14049 5 1 1 14048
0 14050 7 1 2 81977 72818
0 14051 5 1 1 14050
0 14052 7 1 2 14049 14051
0 14053 5 1 1 14052
0 14054 7 1 2 73007 14053
0 14055 5 1 1 14054
0 14056 7 1 2 84031 87474
0 14057 5 1 1 14056
0 14058 7 1 2 14055 14057
0 14059 5 1 1 14058
0 14060 7 1 2 2226 14059
0 14061 5 1 1 14060
0 14062 7 1 2 82901 6012
0 14063 5 2 1 14062
0 14064 7 1 2 69521 73992
0 14065 5 1 1 14064
0 14066 7 1 2 74168 14065
0 14067 5 1 1 14066
0 14068 7 1 2 59835 14067
0 14069 5 1 1 14068
0 14070 7 1 2 77032 73328
0 14071 5 1 1 14070
0 14072 7 1 2 14069 14071
0 14073 5 1 1 14072
0 14074 7 1 2 89270 14073
0 14075 5 1 1 14074
0 14076 7 2 2 71098 73204
0 14077 5 3 1 89272
0 14078 7 1 2 75963 89274
0 14079 5 1 1 14078
0 14080 7 1 2 67034 85790
0 14081 5 1 1 14080
0 14082 7 1 2 72306 89177
0 14083 7 1 2 14081 14082
0 14084 7 1 2 14079 14083
0 14085 5 1 1 14084
0 14086 7 1 2 61266 14085
0 14087 5 1 1 14086
0 14088 7 1 2 2526 14087
0 14089 5 1 1 14088
0 14090 7 1 2 60095 14089
0 14091 5 1 1 14090
0 14092 7 2 2 74964 71442
0 14093 5 1 1 89277
0 14094 7 1 2 67261 89278
0 14095 5 1 1 14094
0 14096 7 1 2 14091 14095
0 14097 5 1 1 14096
0 14098 7 1 2 67933 14097
0 14099 5 1 1 14098
0 14100 7 1 2 14075 14099
0 14101 5 1 1 14100
0 14102 7 1 2 89248 14101
0 14103 5 1 1 14102
0 14104 7 1 2 14061 14103
0 14105 7 1 2 14043 14104
0 14106 5 1 1 14105
0 14107 7 1 2 80846 14106
0 14108 5 1 1 14107
0 14109 7 1 2 13792 14108
0 14110 5 1 1 14109
0 14111 7 1 2 68623 14110
0 14112 5 1 1 14111
0 14113 7 3 2 71699 75938
0 14114 5 1 1 89279
0 14115 7 1 2 72307 14114
0 14116 5 1 1 14115
0 14117 7 1 2 61267 14116
0 14118 5 1 1 14117
0 14119 7 1 2 72964 14118
0 14120 5 1 1 14119
0 14121 7 1 2 62569 14120
0 14122 5 1 1 14121
0 14123 7 2 2 72181 72958
0 14124 7 1 2 89186 89282
0 14125 5 1 1 14124
0 14126 7 1 2 61466 14125
0 14127 5 1 1 14126
0 14128 7 1 2 14122 14127
0 14129 5 1 1 14128
0 14130 7 1 2 62921 14129
0 14131 5 1 1 14130
0 14132 7 1 2 71304 75809
0 14133 5 1 1 14132
0 14134 7 1 2 89283 14133
0 14135 5 1 1 14134
0 14136 7 1 2 74363 14135
0 14137 5 1 1 14136
0 14138 7 1 2 14131 14137
0 14139 5 1 1 14138
0 14140 7 1 2 60289 14139
0 14141 5 1 1 14140
0 14142 7 4 2 61467 72213
0 14143 5 1 1 89284
0 14144 7 1 2 66433 72965
0 14145 5 2 1 14144
0 14146 7 1 2 89280 89288
0 14147 5 1 1 14146
0 14148 7 1 2 14143 14147
0 14149 5 1 1 14148
0 14150 7 1 2 61268 14149
0 14151 5 1 1 14150
0 14152 7 1 2 1211 14151
0 14153 5 1 1 14152
0 14154 7 1 2 77463 14153
0 14155 5 1 1 14154
0 14156 7 1 2 14141 14155
0 14157 5 1 1 14156
0 14158 7 1 2 61672 14157
0 14159 5 1 1 14158
0 14160 7 2 2 75939 77464
0 14161 7 2 2 71646 74943
0 14162 7 4 2 72738 89094
0 14163 7 1 2 89292 89294
0 14164 7 1 2 89290 14163
0 14165 5 1 1 14164
0 14166 7 1 2 14159 14165
0 14167 5 1 1 14166
0 14168 7 1 2 60460 14167
0 14169 5 1 1 14168
0 14170 7 1 2 66216 78314
0 14171 5 2 1 14170
0 14172 7 5 2 61468 79645
0 14173 5 1 1 89300
0 14174 7 1 2 60290 89301
0 14175 5 2 1 14174
0 14176 7 2 2 80899 89305
0 14177 5 24 1 89307
0 14178 7 8 2 60461 61469
0 14179 5 2 1 89333
0 14180 7 4 2 61673 89334
0 14181 5 1 1 89343
0 14182 7 3 2 89309 14181
0 14183 7 1 2 88606 89347
0 14184 5 1 1 14183
0 14185 7 1 2 60291 85466
0 14186 5 1 1 14185
0 14187 7 1 2 14184 14186
0 14188 5 1 1 14187
0 14189 7 1 2 89298 14188
0 14190 5 1 1 14189
0 14191 7 1 2 75886 81065
0 14192 5 8 1 14191
0 14193 7 1 2 72214 89350
0 14194 5 2 1 14193
0 14195 7 2 2 59836 74793
0 14196 5 6 1 89360
0 14197 7 1 2 61030 89361
0 14198 5 2 1 14197
0 14199 7 1 2 72419 89368
0 14200 5 1 1 14199
0 14201 7 1 2 60096 14200
0 14202 5 1 1 14201
0 14203 7 1 2 71765 14202
0 14204 5 1 1 14203
0 14205 7 3 2 62570 71305
0 14206 5 2 1 89370
0 14207 7 1 2 78655 89371
0 14208 5 1 1 14207
0 14209 7 2 2 14204 14208
0 14210 5 1 1 89375
0 14211 7 1 2 62274 14210
0 14212 5 1 1 14211
0 14213 7 1 2 74057 72711
0 14214 5 2 1 14213
0 14215 7 1 2 67542 75964
0 14216 5 4 1 14215
0 14217 7 4 2 71766 89379
0 14218 7 1 2 72308 89383
0 14219 5 3 1 14218
0 14220 7 1 2 89377 89387
0 14221 5 1 1 14220
0 14222 7 1 2 88457 14221
0 14223 5 1 1 14222
0 14224 7 1 2 82719 71915
0 14225 5 2 1 14224
0 14226 7 1 2 73564 73836
0 14227 5 1 1 14226
0 14228 7 1 2 61269 14227
0 14229 7 1 2 89390 14228
0 14230 7 1 2 14223 14229
0 14231 7 1 2 14212 14230
0 14232 5 1 1 14231
0 14233 7 1 2 61470 73748
0 14234 7 1 2 89299 14233
0 14235 7 1 2 14232 14234
0 14236 5 1 1 14235
0 14237 7 1 2 89358 14236
0 14238 5 1 1 14237
0 14239 7 1 2 80847 14238
0 14240 5 1 1 14239
0 14241 7 1 2 14190 14240
0 14242 5 1 1 14241
0 14243 7 1 2 67934 14242
0 14244 5 1 1 14243
0 14245 7 1 2 81400 71445
0 14246 7 1 2 89291 14245
0 14247 5 1 1 14246
0 14248 7 1 2 14244 14247
0 14249 7 1 2 14169 14248
0 14250 5 1 1 14249
0 14251 7 1 2 68287 14250
0 14252 5 1 1 14251
0 14253 7 3 2 67935 70520
0 14254 5 2 1 89392
0 14255 7 1 2 66217 89395
0 14256 5 1 1 14255
0 14257 7 11 2 63376 75252
0 14258 7 6 2 67543 89397
0 14259 7 1 2 75543 72966
0 14260 5 2 1 14259
0 14261 7 3 2 89408 89414
0 14262 7 1 2 14256 89416
0 14263 5 1 1 14262
0 14264 7 2 2 79876 77896
0 14265 5 1 1 89419
0 14266 7 1 2 77771 75094
0 14267 5 3 1 14266
0 14268 7 1 2 79803 89421
0 14269 5 2 1 14268
0 14270 7 1 2 61270 89424
0 14271 5 1 1 14270
0 14272 7 1 2 14265 14271
0 14273 5 1 1 14272
0 14274 7 1 2 72974 14273
0 14275 5 1 1 14274
0 14276 7 4 2 68288 79877
0 14277 7 1 2 87373 89426
0 14278 5 1 1 14277
0 14279 7 1 2 79907 73465
0 14280 7 1 2 82967 14279
0 14281 5 1 1 14280
0 14282 7 1 2 14278 14281
0 14283 7 1 2 14275 14282
0 14284 5 1 1 14283
0 14285 7 1 2 67262 14284
0 14286 5 1 1 14285
0 14287 7 1 2 75136 86863
0 14288 5 1 1 14287
0 14289 7 2 2 80947 82398
0 14290 7 1 2 72975 89430
0 14291 5 2 1 14290
0 14292 7 1 2 14288 89432
0 14293 7 1 2 14286 14292
0 14294 5 1 1 14293
0 14295 7 1 2 69522 14294
0 14296 5 1 1 14295
0 14297 7 1 2 14263 14296
0 14298 5 1 1 14297
0 14299 7 1 2 61674 14298
0 14300 5 1 1 14299
0 14301 7 5 2 61031 71388
0 14302 7 1 2 85896 89434
0 14303 7 3 2 88978 14302
0 14304 7 3 2 66666 78249
0 14305 5 2 1 89442
0 14306 7 1 2 74403 83927
0 14307 5 2 1 14306
0 14308 7 1 2 89445 89447
0 14309 5 1 1 14308
0 14310 7 1 2 89439 14309
0 14311 5 1 1 14310
0 14312 7 1 2 14300 14311
0 14313 5 1 1 14312
0 14314 7 1 2 60462 14313
0 14315 5 1 1 14314
0 14316 7 6 2 75253 80848
0 14317 5 3 1 89449
0 14318 7 4 2 63377 70521
0 14319 7 1 2 89450 89458
0 14320 5 1 1 14319
0 14321 7 2 2 68289 73705
0 14322 7 1 2 89462 89348
0 14323 5 1 1 14322
0 14324 7 1 2 14320 14323
0 14325 5 1 1 14324
0 14326 7 1 2 82922 14325
0 14327 5 1 1 14326
0 14328 7 1 2 79804 84754
0 14329 5 3 1 14328
0 14330 7 1 2 60292 89464
0 14331 5 2 1 14330
0 14332 7 1 2 85966 88098
0 14333 5 1 1 14332
0 14334 7 1 2 89467 14333
0 14335 5 1 1 14334
0 14336 7 1 2 80849 14335
0 14337 5 1 1 14336
0 14338 7 1 2 14327 14337
0 14339 5 1 1 14338
0 14340 7 1 2 67544 14339
0 14341 5 1 1 14340
0 14342 7 6 2 60293 79765
0 14343 5 4 1 89469
0 14344 7 14 2 67035 75254
0 14345 5 2 1 89479
0 14346 7 1 2 85950 85975
0 14347 5 3 1 14346
0 14348 7 1 2 89480 89495
0 14349 5 1 1 14348
0 14350 7 1 2 89475 14349
0 14351 5 1 1 14350
0 14352 7 1 2 80850 73642
0 14353 7 1 2 14351 14352
0 14354 5 1 1 14353
0 14355 7 1 2 14341 14354
0 14356 5 1 1 14355
0 14357 7 1 2 72907 14356
0 14358 5 1 1 14357
0 14359 7 1 2 70594 85258
0 14360 5 2 1 14359
0 14361 7 1 2 61675 89351
0 14362 5 1 1 14361
0 14363 7 1 2 89498 14362
0 14364 5 1 1 14363
0 14365 7 1 2 60463 14364
0 14366 5 1 1 14365
0 14367 7 1 2 81403 14366
0 14368 5 1 1 14367
0 14369 7 1 2 89118 14368
0 14370 5 1 1 14369
0 14371 7 7 2 83596 5740
0 14372 5 6 1 89500
0 14373 7 3 2 62571 70522
0 14374 7 1 2 62922 80851
0 14375 7 1 2 89513 14374
0 14376 7 1 2 89507 14375
0 14377 5 1 1 14376
0 14378 7 1 2 14370 14377
0 14379 5 1 1 14378
0 14380 7 1 2 68290 14379
0 14381 5 1 1 14380
0 14382 7 9 2 60097 82923
0 14383 5 6 1 89516
0 14384 7 1 2 76593 89271
0 14385 5 1 1 14384
0 14386 7 1 2 89525 14385
0 14387 5 1 1 14386
0 14388 7 1 2 75255 14387
0 14389 5 1 1 14388
0 14390 7 1 2 64938 76598
0 14391 5 1 1 14390
0 14392 7 1 2 75482 14391
0 14393 5 1 1 14392
0 14394 7 1 2 14389 14393
0 14395 5 1 1 14394
0 14396 7 1 2 80916 14395
0 14397 5 1 1 14396
0 14398 7 1 2 14381 14397
0 14399 5 1 1 14398
0 14400 7 1 2 71179 14399
0 14401 5 1 1 14400
0 14402 7 1 2 9112 89448
0 14403 5 1 1 14402
0 14404 7 1 2 61676 89440
0 14405 7 1 2 14403 14404
0 14406 5 1 1 14405
0 14407 7 1 2 14401 14406
0 14408 7 1 2 14358 14407
0 14409 7 1 2 14315 14408
0 14410 5 1 1 14409
0 14411 7 1 2 72090 14410
0 14412 5 1 1 14411
0 14413 7 1 2 75949 85942
0 14414 5 1 1 14413
0 14415 7 1 2 82338 89281
0 14416 5 1 1 14415
0 14417 7 1 2 14414 14416
0 14418 5 1 1 14417
0 14419 7 1 2 75256 14418
0 14420 5 1 1 14419
0 14421 7 3 2 66218 83898
0 14422 5 6 1 89531
0 14423 7 1 2 81212 89534
0 14424 5 1 1 14423
0 14425 7 1 2 65151 81217
0 14426 5 1 1 14425
0 14427 7 1 2 67545 14426
0 14428 7 1 2 14424 14427
0 14429 5 1 1 14428
0 14430 7 1 2 14420 14429
0 14431 5 1 1 14430
0 14432 7 1 2 80852 14431
0 14433 5 1 1 14432
0 14434 7 1 2 68291 72470
0 14435 7 1 2 89349 14434
0 14436 5 1 1 14435
0 14437 7 1 2 80853 74137
0 14438 7 1 2 89398 14437
0 14439 5 1 1 14438
0 14440 7 1 2 14436 14439
0 14441 5 1 1 14440
0 14442 7 1 2 67936 14441
0 14443 5 1 1 14442
0 14444 7 3 2 71700 73706
0 14445 7 5 2 67546 75257
0 14446 7 1 2 80917 89543
0 14447 7 1 2 89540 14446
0 14448 5 1 1 14447
0 14449 7 1 2 14443 14448
0 14450 5 1 1 14449
0 14451 7 1 2 61271 14450
0 14452 5 1 1 14451
0 14453 7 1 2 14433 14452
0 14454 5 1 1 14453
0 14455 7 1 2 60098 14454
0 14456 5 1 1 14455
0 14457 7 1 2 64939 78224
0 14458 5 5 1 14457
0 14459 7 5 2 65367 81492
0 14460 5 5 1 89553
0 14461 7 4 2 67263 83739
0 14462 7 1 2 60294 80641
0 14463 7 2 2 89563 14462
0 14464 7 1 2 89554 89567
0 14465 5 2 1 14464
0 14466 7 1 2 80166 89568
0 14467 5 2 1 14466
0 14468 7 1 2 73664 86692
0 14469 5 1 1 14468
0 14470 7 1 2 89476 14469
0 14471 5 1 1 14470
0 14472 7 1 2 69523 14471
0 14473 5 2 1 14472
0 14474 7 2 2 75544 82902
0 14475 5 1 1 89575
0 14476 7 4 2 75258 14475
0 14477 5 1 1 89577
0 14478 7 1 2 80109 89578
0 14479 5 1 1 14478
0 14480 7 1 2 89573 14479
0 14481 5 1 1 14480
0 14482 7 1 2 61677 14481
0 14483 5 1 1 14482
0 14484 7 1 2 89571 14483
0 14485 5 1 1 14484
0 14486 7 1 2 60464 14485
0 14487 5 1 1 14486
0 14488 7 1 2 89569 14487
0 14489 5 1 1 14488
0 14490 7 1 2 89548 14489
0 14491 5 1 1 14490
0 14492 7 1 2 67937 89352
0 14493 5 3 1 14492
0 14494 7 7 2 67547 71701
0 14495 7 3 2 75259 86022
0 14496 7 1 2 89584 89591
0 14497 5 1 1 14496
0 14498 7 1 2 89581 14497
0 14499 5 1 1 14498
0 14500 7 1 2 67264 14499
0 14501 5 1 1 14500
0 14502 7 2 2 87374 89481
0 14503 5 1 1 89594
0 14504 7 1 2 14501 14503
0 14505 5 1 1 14504
0 14506 7 1 2 69524 14505
0 14507 5 1 1 14506
0 14508 7 2 2 59484 81231
0 14509 7 1 2 84825 89596
0 14510 5 1 1 14509
0 14511 7 2 2 64478 73038
0 14512 5 3 1 89598
0 14513 7 3 2 76403 89600
0 14514 5 1 1 89603
0 14515 7 1 2 62923 82753
0 14516 7 1 2 89604 14515
0 14517 5 1 1 14516
0 14518 7 1 2 14510 14517
0 14519 5 1 1 14518
0 14520 7 1 2 62572 14519
0 14521 5 1 1 14520
0 14522 7 1 2 83438 82399
0 14523 5 1 1 14522
0 14524 7 1 2 68292 14523
0 14525 7 1 2 14521 14524
0 14526 7 1 2 14507 14525
0 14527 5 1 1 14526
0 14528 7 2 2 60295 88099
0 14529 5 2 1 89606
0 14530 7 4 2 59485 75260
0 14531 5 1 1 89610
0 14532 7 1 2 88010 89057
0 14533 7 1 2 89611 14532
0 14534 5 1 1 14533
0 14535 7 1 2 89608 14534
0 14536 5 1 1 14535
0 14537 7 1 2 61272 14536
0 14538 5 1 1 14537
0 14539 7 1 2 83504 79054
0 14540 5 1 1 14539
0 14541 7 1 2 63378 14540
0 14542 7 1 2 14538 14541
0 14543 5 1 1 14542
0 14544 7 1 2 80854 14543
0 14545 7 1 2 14527 14544
0 14546 5 1 1 14545
0 14547 7 1 2 14491 14546
0 14548 7 1 2 14456 14547
0 14549 5 1 1 14548
0 14550 7 1 2 71180 14549
0 14551 5 1 1 14550
0 14552 7 2 2 75261 82924
0 14553 7 1 2 75950 89614
0 14554 5 1 1 14553
0 14555 7 1 2 75483 73707
0 14556 5 1 1 14555
0 14557 7 1 2 14554 14556
0 14558 5 1 1 14557
0 14559 7 1 2 80918 14558
0 14560 5 1 1 14559
0 14561 7 2 2 68293 73651
0 14562 7 2 2 84826 85299
0 14563 5 2 1 89618
0 14564 7 1 2 79274 89620
0 14565 5 1 1 14564
0 14566 7 1 2 60296 14565
0 14567 5 1 1 14566
0 14568 7 2 2 61273 82400
0 14569 5 5 1 89622
0 14570 7 1 2 89535 89624
0 14571 5 2 1 14570
0 14572 7 1 2 61678 89629
0 14573 5 1 1 14572
0 14574 7 1 2 14567 14573
0 14575 5 1 1 14574
0 14576 7 1 2 60465 14575
0 14577 5 1 1 14576
0 14578 7 2 2 61471 88080
0 14579 7 1 2 85654 89631
0 14580 5 1 1 14579
0 14581 7 1 2 14577 14580
0 14582 5 1 1 14581
0 14583 7 1 2 89616 14582
0 14584 5 1 1 14583
0 14585 7 1 2 14560 14584
0 14586 5 1 1 14585
0 14587 7 1 2 67548 14586
0 14588 5 1 1 14587
0 14589 7 1 2 85976 89422
0 14590 5 1 1 14589
0 14591 7 1 2 69525 14590
0 14592 5 1 1 14591
0 14593 7 1 2 73008 89496
0 14594 5 1 1 14593
0 14595 7 1 2 14592 14594
0 14596 5 1 1 14595
0 14597 7 1 2 75262 14596
0 14598 5 1 1 14597
0 14599 7 1 2 83400 88100
0 14600 5 2 1 14599
0 14601 7 1 2 89574 89633
0 14602 7 1 2 14598 14601
0 14603 5 1 1 14602
0 14604 7 1 2 61679 14603
0 14605 5 1 1 14604
0 14606 7 1 2 89572 14605
0 14607 5 1 1 14606
0 14608 7 1 2 60466 14607
0 14609 5 1 1 14608
0 14610 7 1 2 89570 14609
0 14611 5 1 1 14610
0 14612 7 1 2 71702 14611
0 14613 5 1 1 14612
0 14614 7 1 2 14588 14613
0 14615 5 1 1 14614
0 14616 7 1 2 72908 14615
0 14617 5 1 1 14616
0 14618 7 5 2 60099 60467
0 14619 7 1 2 81379 89635
0 14620 5 1 1 14619
0 14621 7 1 2 85259 88607
0 14622 5 1 1 14621
0 14623 7 1 2 81380 14622
0 14624 5 1 1 14623
0 14625 7 1 2 60468 14624
0 14626 5 1 1 14625
0 14627 7 5 2 61032 81493
0 14628 7 6 2 60100 65368
0 14629 7 2 2 89645 89095
0 14630 7 1 2 89640 89651
0 14631 5 1 1 14630
0 14632 7 1 2 14626 14631
0 14633 5 1 1 14632
0 14634 7 1 2 72165 73647
0 14635 5 2 1 14634
0 14636 7 1 2 67549 89653
0 14637 7 1 2 14633 14636
0 14638 5 1 1 14637
0 14639 7 1 2 14620 14638
0 14640 5 1 1 14639
0 14641 7 1 2 68294 14640
0 14642 5 1 1 14641
0 14643 7 1 2 80707 75784
0 14644 7 1 2 85260 14643
0 14645 5 1 1 14644
0 14646 7 1 2 81381 14645
0 14647 5 1 1 14646
0 14648 7 1 2 80948 14647
0 14649 5 1 1 14648
0 14650 7 1 2 69645 85360
0 14651 5 1 1 14650
0 14652 7 4 2 60297 81494
0 14653 7 1 2 63379 89655
0 14654 7 1 2 14651 14653
0 14655 5 1 1 14654
0 14656 7 1 2 14649 14655
0 14657 5 1 1 14656
0 14658 7 1 2 60469 14657
0 14659 5 1 1 14658
0 14660 7 1 2 79930 71403
0 14661 7 1 2 76594 89555
0 14662 7 1 2 14660 14661
0 14663 5 1 1 14662
0 14664 7 1 2 14659 14663
0 14665 5 1 1 14664
0 14666 7 1 2 71181 14665
0 14667 5 1 1 14666
0 14668 7 1 2 75484 72909
0 14669 5 1 1 14668
0 14670 7 3 2 75263 89415
0 14671 7 2 2 71703 89659
0 14672 5 1 1 89662
0 14673 7 1 2 69526 89663
0 14674 5 1 1 14673
0 14675 7 1 2 14669 14674
0 14676 5 1 1 14675
0 14677 7 1 2 80919 14676
0 14678 5 1 1 14677
0 14679 7 1 2 14667 14678
0 14680 7 1 2 14642 14679
0 14681 5 1 1 14680
0 14682 7 1 2 78588 14681
0 14683 5 1 1 14682
0 14684 7 2 2 62573 74058
0 14685 5 2 1 89664
0 14686 7 2 2 73708 89666
0 14687 5 1 1 89668
0 14688 7 1 2 82956 89669
0 14689 5 1 1 14688
0 14690 7 2 2 67938 82764
0 14691 5 1 1 89670
0 14692 7 1 2 14689 14691
0 14693 5 1 1 14692
0 14694 7 1 2 89660 14693
0 14695 5 1 1 14694
0 14696 7 1 2 75485 88608
0 14697 5 1 1 14696
0 14698 7 1 2 14695 14697
0 14699 5 1 1 14698
0 14700 7 1 2 80920 14699
0 14701 5 1 1 14700
0 14702 7 1 2 14683 14701
0 14703 7 1 2 14617 14702
0 14704 7 1 2 14551 14703
0 14705 7 1 2 14412 14704
0 14706 7 1 2 14252 14705
0 14707 5 1 1 14706
0 14708 7 1 2 85508 14707
0 14709 5 1 1 14708
0 14710 7 1 2 83182 77465
0 14711 5 2 1 14710
0 14712 7 3 2 74000 78288
0 14713 5 1 1 89674
0 14714 7 1 2 73946 89675
0 14715 5 1 1 14714
0 14716 7 1 2 89672 14715
0 14717 5 1 1 14716
0 14718 7 1 2 75264 14717
0 14719 5 1 1 14718
0 14720 7 1 2 67036 89470
0 14721 5 1 1 14720
0 14722 7 1 2 14719 14721
0 14723 5 1 1 14722
0 14724 7 1 2 63688 14723
0 14725 5 1 1 14724
0 14726 7 2 2 60892 83299
0 14727 5 2 1 89677
0 14728 7 17 2 62924 83519
0 14729 5 2 1 89681
0 14730 7 1 2 76171 89682
0 14731 5 1 1 14730
0 14732 7 17 2 67939 78738
0 14733 7 1 2 74663 89700
0 14734 5 1 1 14733
0 14735 7 1 2 14731 14734
0 14736 5 1 1 14735
0 14737 7 1 2 89678 14736
0 14738 5 1 1 14737
0 14739 7 1 2 14725 14738
0 14740 5 1 1 14739
0 14741 7 1 2 80855 14740
0 14742 5 1 1 14741
0 14743 7 7 2 60893 62925
0 14744 7 2 2 76631 89717
0 14745 5 1 1 89724
0 14746 7 1 2 83307 14745
0 14747 5 3 1 14746
0 14748 7 1 2 60298 89726
0 14749 5 1 1 14748
0 14750 7 1 2 80760 77515
0 14751 5 1 1 14750
0 14752 7 1 2 14749 14751
0 14753 5 1 1 14752
0 14754 7 1 2 59486 14753
0 14755 5 1 1 14754
0 14756 7 2 2 66434 69299
0 14757 5 1 1 89729
0 14758 7 1 2 60299 89730
0 14759 5 2 1 14758
0 14760 7 1 2 14755 89731
0 14761 5 1 1 14760
0 14762 7 1 2 67037 14761
0 14763 5 1 1 14762
0 14764 7 1 2 71665 74729
0 14765 5 1 1 14764
0 14766 7 1 2 14763 14765
0 14767 5 1 1 14766
0 14768 7 1 2 68295 14767
0 14769 5 1 1 14768
0 14770 7 3 2 63380 69300
0 14771 7 1 2 75486 89733
0 14772 5 1 1 14771
0 14773 7 1 2 14769 14772
0 14774 5 1 1 14773
0 14775 7 1 2 68624 14774
0 14776 5 1 1 14775
0 14777 7 2 2 74095 88101
0 14778 7 6 2 59487 60300
0 14779 5 1 1 89738
0 14780 7 3 2 60894 89739
0 14781 7 1 2 89701 89744
0 14782 7 1 2 89736 14781
0 14783 5 1 1 14782
0 14784 7 1 2 14776 14783
0 14785 5 1 1 14784
0 14786 7 1 2 81166 14785
0 14787 5 1 1 14786
0 14788 7 1 2 14742 14787
0 14789 5 1 1 14788
0 14790 7 1 2 70141 14789
0 14791 5 1 1 14790
0 14792 7 8 2 68625 79434
0 14793 7 2 2 89263 89747
0 14794 7 1 2 82603 89755
0 14795 5 1 1 14794
0 14796 7 1 2 72091 89756
0 14797 5 1 1 14796
0 14798 7 1 2 61680 78556
0 14799 5 1 1 14798
0 14800 7 1 2 71389 85300
0 14801 5 2 1 14800
0 14802 7 1 2 14799 89757
0 14803 5 1 1 14802
0 14804 7 1 2 83183 14803
0 14805 5 1 1 14804
0 14806 7 1 2 76762 81102
0 14807 5 1 1 14806
0 14808 7 1 2 14805 14807
0 14809 5 1 1 14808
0 14810 7 1 2 60895 78158
0 14811 7 1 2 14809 14810
0 14812 5 1 1 14811
0 14813 7 1 2 14797 14812
0 14814 5 1 1 14813
0 14815 7 1 2 61472 14814
0 14816 5 1 1 14815
0 14817 7 3 2 59488 89023
0 14818 5 1 1 89759
0 14819 7 1 2 68296 89760
0 14820 5 1 1 14819
0 14821 7 1 2 13739 14820
0 14822 5 1 1 14821
0 14823 7 1 2 60896 88261
0 14824 7 1 2 14822 14823
0 14825 5 1 1 14824
0 14826 7 1 2 14816 14825
0 14827 5 1 1 14826
0 14828 7 1 2 67265 14827
0 14829 5 1 1 14828
0 14830 7 1 2 14795 14829
0 14831 5 1 1 14830
0 14832 7 1 2 67038 14831
0 14833 5 1 1 14832
0 14834 7 19 2 66435 68626
0 14835 5 1 1 89762
0 14836 7 1 2 76172 81232
0 14837 5 1 1 14836
0 14838 7 1 2 75769 14837
0 14839 5 1 1 14838
0 14840 7 1 2 59489 14839
0 14841 5 1 1 14840
0 14842 7 1 2 65152 84102
0 14843 5 1 1 14842
0 14844 7 1 2 14841 14843
0 14845 5 1 1 14844
0 14846 7 1 2 89763 14845
0 14847 5 1 1 14846
0 14848 7 3 2 63689 70523
0 14849 7 1 2 83491 89781
0 14850 5 1 1 14849
0 14851 7 1 2 14847 14850
0 14852 5 1 1 14851
0 14853 7 1 2 63381 14852
0 14854 5 1 1 14853
0 14855 7 1 2 81066 89026
0 14856 5 3 1 14855
0 14857 7 1 2 75008 78739
0 14858 7 1 2 89784 14857
0 14859 5 1 1 14858
0 14860 7 1 2 61681 14859
0 14861 7 1 2 14854 14860
0 14862 5 1 1 14861
0 14863 7 1 2 84097 89734
0 14864 7 2 2 83492 14863
0 14865 5 1 1 89787
0 14866 7 6 2 59490 69301
0 14867 5 3 1 89789
0 14868 7 3 2 68297 89790
0 14869 5 1 1 89798
0 14870 7 1 2 79308 72757
0 14871 5 1 1 14870
0 14872 7 1 2 89799 14871
0 14873 5 1 1 14872
0 14874 7 1 2 14865 14873
0 14875 5 1 1 14874
0 14876 7 1 2 68627 14875
0 14877 5 1 1 14876
0 14878 7 2 2 71390 80938
0 14879 5 1 1 89801
0 14880 7 2 2 75709 89802
0 14881 7 1 2 78740 89803
0 14882 5 1 1 14881
0 14883 7 1 2 66667 14882
0 14884 7 1 2 14877 14883
0 14885 5 1 1 14884
0 14886 7 1 2 67940 14885
0 14887 7 1 2 14862 14886
0 14888 5 1 1 14887
0 14889 7 1 2 79435 88102
0 14890 5 2 1 14889
0 14891 7 1 2 81123 89805
0 14892 5 1 1 14891
0 14893 7 1 2 84304 89264
0 14894 7 1 2 14892 14893
0 14895 5 1 1 14894
0 14896 7 1 2 14888 14895
0 14897 7 1 2 14833 14896
0 14898 5 1 1 14897
0 14899 7 1 2 60470 14898
0 14900 5 1 1 14899
0 14901 7 1 2 81382 89499
0 14902 5 1 1 14901
0 14903 7 1 2 83051 14902
0 14904 5 1 1 14903
0 14905 7 17 2 61682 67039
0 14906 7 1 2 61473 89807
0 14907 7 1 2 89265 14906
0 14908 5 1 1 14907
0 14909 7 1 2 14904 14908
0 14910 5 1 1 14909
0 14911 7 1 2 69302 14910
0 14912 5 1 1 14911
0 14913 7 3 2 61683 75045
0 14914 5 1 1 89824
0 14915 7 1 2 88103 89266
0 14916 7 1 2 89825 14915
0 14917 5 1 1 14916
0 14918 7 1 2 14912 14917
0 14919 5 1 1 14918
0 14920 7 1 2 68298 14919
0 14921 5 1 1 14920
0 14922 7 1 2 88081 89788
0 14923 5 1 1 14922
0 14924 7 1 2 14921 14923
0 14925 5 1 1 14924
0 14926 7 1 2 68628 14925
0 14927 5 1 1 14926
0 14928 7 2 2 59491 83804
0 14929 5 3 1 89827
0 14930 7 6 2 60301 79878
0 14931 5 2 1 89832
0 14932 7 2 2 61684 89833
0 14933 7 1 2 83216 89840
0 14934 7 1 2 89828 14933
0 14935 5 1 1 14934
0 14936 7 1 2 14927 14935
0 14937 5 1 1 14936
0 14938 7 1 2 65369 14937
0 14939 5 1 1 14938
0 14940 7 1 2 14900 14939
0 14941 7 1 2 14791 14940
0 14942 5 1 1 14941
0 14943 7 1 2 71182 14942
0 14944 5 1 1 14943
0 14945 7 2 2 74730 83445
0 14946 7 2 2 82957 89842
0 14947 5 1 1 89844
0 14948 7 3 2 83358 88609
0 14949 7 1 2 78589 88969
0 14950 7 1 2 89846 14949
0 14951 5 1 1 14950
0 14952 7 1 2 14947 14951
0 14953 5 1 1 14952
0 14954 7 1 2 63382 14953
0 14955 5 1 1 14954
0 14956 7 2 2 67266 81531
0 14957 7 1 2 79202 82943
0 14958 7 1 2 82958 14957
0 14959 7 1 2 89849 14958
0 14960 5 1 1 14959
0 14961 7 1 2 14955 14960
0 14962 5 1 1 14961
0 14963 7 1 2 61685 14962
0 14964 5 1 1 14963
0 14965 7 1 2 81048 83381
0 14966 7 3 2 60302 74816
0 14967 7 2 2 62926 78741
0 14968 7 1 2 89851 89854
0 14969 7 1 2 14965 14968
0 14970 5 1 1 14969
0 14971 7 1 2 14964 14970
0 14972 5 1 1 14971
0 14973 7 1 2 60471 14972
0 14974 5 1 1 14973
0 14975 7 6 2 61686 67267
0 14976 7 3 2 63690 89856
0 14977 7 1 2 87375 89862
0 14978 5 1 1 14977
0 14979 7 1 2 85322 89018
0 14980 5 1 1 14979
0 14981 7 1 2 14978 14980
0 14982 5 1 1 14981
0 14983 7 1 2 85897 89101
0 14984 7 1 2 14982 14983
0 14985 5 1 1 14984
0 14986 7 1 2 14974 14985
0 14987 5 1 1 14986
0 14988 7 1 2 60897 14987
0 14989 5 1 1 14988
0 14990 7 1 2 89847 89020
0 14991 5 1 1 14990
0 14992 7 1 2 67268 89845
0 14993 5 1 1 14992
0 14994 7 1 2 14991 14993
0 14995 5 1 1 14994
0 14996 7 1 2 63383 14995
0 14997 5 1 1 14996
0 14998 7 2 2 67550 75137
0 14999 5 1 1 89865
0 15000 7 1 2 82959 78742
0 15001 7 1 2 89866 15000
0 15002 5 1 1 15001
0 15003 7 1 2 14997 15002
0 15004 5 1 1 15003
0 15005 7 1 2 80856 15004
0 15006 5 1 1 15005
0 15007 7 2 2 81388 88610
0 15008 7 1 2 83765 86868
0 15009 7 1 2 89867 15008
0 15010 5 1 1 15009
0 15011 7 1 2 15006 15010
0 15012 7 1 2 14989 15011
0 15013 5 1 1 15012
0 15014 7 1 2 59492 15013
0 15015 5 1 1 15014
0 15016 7 2 2 66436 85776
0 15017 7 9 2 60472 62927
0 15018 7 2 2 75681 89871
0 15019 5 1 1 89880
0 15020 7 1 2 89869 89881
0 15021 5 1 1 15020
0 15022 7 3 2 61474 80110
0 15023 5 2 1 89882
0 15024 7 1 2 67551 89883
0 15025 5 1 1 15024
0 15026 7 1 2 86694 15025
0 15027 5 1 1 15026
0 15028 7 1 2 61274 15027
0 15029 5 1 1 15028
0 15030 7 3 2 67269 79879
0 15031 7 1 2 86650 89887
0 15032 5 1 1 15031
0 15033 7 1 2 15029 15032
0 15034 5 1 1 15033
0 15035 7 1 2 72092 15034
0 15036 5 1 1 15035
0 15037 7 1 2 75830 89015
0 15038 5 1 1 15037
0 15039 7 1 2 79766 82960
0 15040 5 1 1 15039
0 15041 7 1 2 15038 15040
0 15042 5 1 1 15041
0 15043 7 1 2 89585 15042
0 15044 5 1 1 15043
0 15045 7 2 2 68299 81252
0 15046 7 1 2 88339 89890
0 15047 5 1 1 15046
0 15048 7 1 2 82925 89465
0 15049 5 1 1 15048
0 15050 7 1 2 15047 15049
0 15051 7 1 2 15044 15050
0 15052 7 1 2 15036 15051
0 15053 5 1 1 15052
0 15054 7 1 2 81167 15053
0 15055 5 1 1 15054
0 15056 7 1 2 15021 15055
0 15057 5 1 1 15056
0 15058 7 1 2 68629 15057
0 15059 5 1 1 15058
0 15060 7 1 2 79871 6294
0 15061 5 1 1 15060
0 15062 7 1 2 60898 15061
0 15063 5 1 1 15062
0 15064 7 1 2 3403 81206
0 15065 7 1 2 15063 15064
0 15066 5 1 1 15065
0 15067 7 1 2 59493 15066
0 15068 5 1 1 15067
0 15069 7 1 2 76404 81201
0 15070 5 1 1 15069
0 15071 7 1 2 15068 15070
0 15072 5 1 1 15071
0 15073 7 1 2 61275 15072
0 15074 5 1 1 15073
0 15075 7 2 2 61276 79880
0 15076 7 1 2 89735 89892
0 15077 5 1 1 15076
0 15078 7 1 2 79869 71704
0 15079 5 1 1 15078
0 15080 7 7 2 74059 89380
0 15081 5 2 1 89894
0 15082 7 1 2 66437 75125
0 15083 5 3 1 15082
0 15084 7 1 2 85927 89903
0 15085 7 1 2 89901 15084
0 15086 5 1 1 15085
0 15087 7 1 2 15079 15086
0 15088 5 1 1 15087
0 15089 7 1 2 67941 15088
0 15090 5 1 1 15089
0 15091 7 1 2 15077 15090
0 15092 7 1 2 15074 15091
0 15093 5 1 1 15092
0 15094 7 1 2 83149 15093
0 15095 5 1 1 15094
0 15096 7 1 2 15059 15095
0 15097 5 1 1 15096
0 15098 7 1 2 72976 15097
0 15099 5 1 1 15098
0 15100 7 1 2 82604 88600
0 15101 5 2 1 15100
0 15102 7 3 2 63384 71391
0 15103 5 1 1 89908
0 15104 7 2 2 69303 72215
0 15105 7 1 2 89909 89911
0 15106 5 1 1 15105
0 15107 7 1 2 89906 15106
0 15108 5 1 1 15107
0 15109 7 1 2 67040 15108
0 15110 5 1 1 15109
0 15111 7 2 2 82605 75064
0 15112 5 1 1 89913
0 15113 7 1 2 60899 89914
0 15114 5 1 1 15113
0 15115 7 1 2 15110 15114
0 15116 5 1 1 15115
0 15117 7 1 2 63691 15116
0 15118 5 1 1 15117
0 15119 7 3 2 69175 84862
0 15120 5 1 1 89915
0 15121 7 1 2 74248 89916
0 15122 5 1 1 15121
0 15123 7 1 2 15118 15122
0 15124 5 1 1 15123
0 15125 7 1 2 61277 15124
0 15126 5 1 1 15125
0 15127 7 1 2 68300 85050
0 15128 5 2 1 15127
0 15129 7 1 2 81739 79009
0 15130 7 1 2 75450 15129
0 15131 7 1 2 89918 15130
0 15132 5 1 1 15131
0 15133 7 1 2 15126 15132
0 15134 5 1 1 15133
0 15135 7 1 2 80857 15134
0 15136 5 1 1 15135
0 15137 7 26 2 68301 68630
0 15138 7 8 2 66668 89920
0 15139 5 6 1 89946
0 15140 7 1 2 85588 89947
0 15141 5 1 1 15140
0 15142 7 1 2 73947 85289
0 15143 5 1 1 15142
0 15144 7 1 2 15141 15143
0 15145 5 1 1 15144
0 15146 7 1 2 89102 15145
0 15147 5 1 1 15146
0 15148 7 2 2 74096 78743
0 15149 7 1 2 80560 81495
0 15150 7 1 2 89960 15149
0 15151 5 1 1 15150
0 15152 7 1 2 15147 15151
0 15153 5 1 1 15152
0 15154 7 1 2 69102 15153
0 15155 5 1 1 15154
0 15156 7 6 2 65153 83520
0 15157 5 2 1 89962
0 15158 7 1 2 85467 89963
0 15159 7 1 2 76311 15158
0 15160 5 1 1 15159
0 15161 7 1 2 15155 15160
0 15162 5 1 1 15161
0 15163 7 1 2 67942 15162
0 15164 5 1 1 15163
0 15165 7 7 2 61475 78744
0 15166 5 3 1 89970
0 15167 7 2 2 68631 69103
0 15168 5 1 1 89980
0 15169 7 1 2 63385 89981
0 15170 5 1 1 15169
0 15171 7 1 2 89977 15170
0 15172 5 1 1 15171
0 15173 7 1 2 82961 89103
0 15174 7 1 2 15172 15173
0 15175 5 1 1 15174
0 15176 7 1 2 68632 79931
0 15177 7 1 2 75138 15176
0 15178 7 1 2 89016 15177
0 15179 5 1 1 15178
0 15180 7 1 2 15175 15179
0 15181 5 1 1 15180
0 15182 7 1 2 59494 15181
0 15183 5 1 1 15182
0 15184 7 3 2 67270 83521
0 15185 5 1 1 89982
0 15186 7 1 2 89978 15185
0 15187 5 2 1 15186
0 15188 7 1 2 88681 89985
0 15189 5 1 1 15188
0 15190 7 3 2 63692 80807
0 15191 7 1 2 79881 78590
0 15192 7 1 2 89987 15191
0 15193 5 1 1 15192
0 15194 7 1 2 15189 15193
0 15195 5 1 1 15194
0 15196 7 1 2 89104 15195
0 15197 5 1 1 15196
0 15198 7 1 2 15183 15197
0 15199 5 1 1 15198
0 15200 7 1 2 67552 15199
0 15201 5 1 1 15200
0 15202 7 2 2 61278 74518
0 15203 5 1 1 89990
0 15204 7 1 2 83446 89991
0 15205 5 1 1 15204
0 15206 7 2 2 71705 89435
0 15207 7 1 2 77114 83579
0 15208 7 1 2 89992 15207
0 15209 5 1 1 15208
0 15210 7 1 2 15205 15209
0 15211 5 1 1 15210
0 15212 7 1 2 83740 15211
0 15213 5 1 1 15212
0 15214 7 2 2 83522 72216
0 15215 7 1 2 71392 89994
0 15216 5 1 1 15215
0 15217 7 1 2 15213 15216
0 15218 5 1 1 15217
0 15219 7 1 2 61476 15218
0 15220 5 1 1 15219
0 15221 7 1 2 73694 85977
0 15222 5 1 1 15221
0 15223 7 4 2 59837 68633
0 15224 7 1 2 89436 89996
0 15225 7 1 2 89497 15224
0 15226 7 1 2 15222 15225
0 15227 5 1 1 15226
0 15228 7 1 2 15220 15227
0 15229 7 1 2 15201 15228
0 15230 5 1 1 15229
0 15231 7 1 2 81168 15230
0 15232 5 1 1 15231
0 15233 7 1 2 15164 15232
0 15234 7 1 2 15136 15233
0 15235 7 1 2 15099 15234
0 15236 7 1 2 15015 15235
0 15237 7 1 2 14944 15236
0 15238 5 1 1 15237
0 15239 7 1 2 68852 15238
0 15240 5 1 1 15239
0 15241 7 1 2 67553 83236
0 15242 5 2 1 15241
0 15243 7 1 2 75858 90000
0 15244 5 1 1 15243
0 15245 7 1 2 60303 15244
0 15246 5 1 1 15245
0 15247 7 1 2 4480 90001
0 15248 5 1 1 15247
0 15249 7 1 2 61477 15248
0 15250 5 1 1 15249
0 15251 7 1 2 15246 15250
0 15252 5 1 1 15251
0 15253 7 1 2 68634 15252
0 15254 5 1 1 15253
0 15255 7 1 2 87516 89961
0 15256 5 1 1 15255
0 15257 7 1 2 15254 15256
0 15258 5 1 1 15257
0 15259 7 1 2 67943 15258
0 15260 5 1 1 15259
0 15261 7 1 2 83944 83523
0 15262 5 1 1 15261
0 15263 7 1 2 15260 15262
0 15264 5 1 1 15263
0 15265 7 1 2 72093 15264
0 15266 5 1 1 15265
0 15267 7 1 2 70524 89592
0 15268 5 1 1 15267
0 15269 7 1 2 82428 15268
0 15270 5 1 1 15269
0 15271 7 1 2 89586 15270
0 15272 5 1 1 15271
0 15273 7 1 2 62275 89595
0 15274 5 1 1 15273
0 15275 7 3 2 75265 78369
0 15276 7 1 2 75545 90002
0 15277 5 1 1 15276
0 15278 7 1 2 68302 15277
0 15279 7 1 2 15274 15278
0 15280 7 1 2 15272 15279
0 15281 5 1 1 15280
0 15282 7 1 2 89579 89587
0 15283 5 1 1 15282
0 15284 7 1 2 63386 85997
0 15285 7 1 2 15283 15284
0 15286 5 1 1 15285
0 15287 7 1 2 68635 15286
0 15288 7 1 2 15281 15287
0 15289 5 1 1 15288
0 15290 7 5 2 67271 72471
0 15291 5 1 1 90005
0 15292 7 2 2 75487 75710
0 15293 7 1 2 85487 90010
0 15294 7 1 2 90006 15293
0 15295 5 1 1 15294
0 15296 7 1 2 15289 15295
0 15297 7 1 2 15266 15296
0 15298 5 1 1 15297
0 15299 7 1 2 81169 15298
0 15300 5 1 1 15299
0 15301 7 4 2 62070 77423
0 15302 5 3 1 90012
0 15303 7 1 2 78187 72182
0 15304 5 1 1 15303
0 15305 7 1 2 90016 15304
0 15306 5 1 1 15305
0 15307 7 1 2 66219 15306
0 15308 5 1 1 15307
0 15309 7 1 2 62928 77624
0 15310 5 1 1 15309
0 15311 7 1 2 15308 15310
0 15312 5 1 1 15311
0 15313 7 1 2 89764 15312
0 15314 5 1 1 15313
0 15315 7 1 2 69288 74493
0 15316 5 5 1 15315
0 15317 7 1 2 90019 89834
0 15318 5 1 1 15317
0 15319 7 2 2 79984 76003
0 15320 7 1 2 15291 90024
0 15321 5 1 1 15320
0 15322 7 1 2 89615 15321
0 15323 5 1 1 15322
0 15324 7 1 2 15318 15323
0 15325 5 1 1 15324
0 15326 7 1 2 63693 15325
0 15327 5 1 1 15326
0 15328 7 1 2 15314 15327
0 15329 5 1 1 15328
0 15330 7 1 2 63387 15329
0 15331 5 1 1 15330
0 15332 7 1 2 76405 89593
0 15333 5 1 1 15332
0 15334 7 2 2 66438 78125
0 15335 5 1 1 90026
0 15336 7 1 2 61279 69104
0 15337 7 1 2 90027 15336
0 15338 5 1 1 15337
0 15339 7 1 2 15333 15338
0 15340 5 1 1 15339
0 15341 7 1 2 67554 15340
0 15342 5 1 1 15341
0 15343 7 3 2 75711 82401
0 15344 5 2 1 90028
0 15345 7 6 2 62929 75266
0 15346 5 7 1 90033
0 15347 7 1 2 62574 90039
0 15348 5 1 1 15347
0 15349 7 2 2 75887 81054
0 15350 5 1 1 90046
0 15351 7 1 2 89536 90047
0 15352 5 1 1 15351
0 15353 7 1 2 15348 15352
0 15354 5 1 1 15353
0 15355 7 1 2 90031 15354
0 15356 5 1 1 15355
0 15357 7 1 2 89791 15356
0 15358 5 1 1 15357
0 15359 7 1 2 15342 15358
0 15360 5 1 1 15359
0 15361 7 1 2 78745 15360
0 15362 5 1 1 15361
0 15363 7 1 2 15331 15362
0 15364 5 1 1 15363
0 15365 7 1 2 80858 15364
0 15366 5 1 1 15365
0 15367 7 1 2 67944 89921
0 15368 7 1 2 82698 15367
0 15369 7 1 2 88180 88887
0 15370 7 1 2 15368 15369
0 15371 5 1 1 15370
0 15372 7 1 2 15366 15371
0 15373 7 1 2 15300 15372
0 15374 5 1 1 15373
0 15375 7 1 2 68853 15374
0 15376 5 1 1 15375
0 15377 7 2 2 78052 83766
0 15378 7 2 2 80100 89335
0 15379 7 1 2 90020 90050
0 15380 7 1 2 90048 15379
0 15381 5 1 1 15380
0 15382 7 1 2 15376 15381
0 15383 5 1 1 15382
0 15384 7 1 2 72910 15383
0 15385 5 1 1 15384
0 15386 7 2 2 63388 89740
0 15387 7 1 2 74649 90052
0 15388 5 1 1 15387
0 15389 7 1 2 3920 80968
0 15390 5 2 1 15389
0 15391 7 1 2 76763 85928
0 15392 7 1 2 90054 15391
0 15393 5 1 1 15392
0 15394 7 7 2 61280 72739
0 15395 7 1 2 83401 90056
0 15396 5 1 1 15395
0 15397 7 1 2 15112 15396
0 15398 7 1 2 15393 15397
0 15399 5 1 1 15398
0 15400 7 1 2 67945 15399
0 15401 5 1 1 15400
0 15402 7 1 2 15388 15401
0 15403 5 1 1 15402
0 15404 7 1 2 68636 15403
0 15405 5 1 1 15404
0 15406 7 1 2 83670 89228
0 15407 5 1 1 15406
0 15408 7 1 2 15405 15407
0 15409 5 1 1 15408
0 15410 7 1 2 81170 15409
0 15411 5 1 1 15410
0 15412 7 10 2 70595 75488
0 15413 5 3 1 90063
0 15414 7 2 2 84333 90064
0 15415 7 2 2 80949 84377
0 15416 5 1 1 90078
0 15417 7 1 2 90076 90079
0 15418 5 1 1 15417
0 15419 7 3 2 59495 83524
0 15420 5 1 1 90080
0 15421 7 1 2 75414 90081
0 15422 5 1 1 15421
0 15423 7 2 2 75267 78746
0 15424 5 1 1 90083
0 15425 7 1 2 15422 15424
0 15426 5 2 1 15425
0 15427 7 1 2 82890 90085
0 15428 5 1 1 15427
0 15429 7 2 2 76385 89702
0 15430 5 1 1 90087
0 15431 7 1 2 61478 90088
0 15432 5 1 1 15431
0 15433 7 1 2 15428 15432
0 15434 5 1 1 15433
0 15435 7 1 2 62575 15434
0 15436 5 1 1 15435
0 15437 7 2 2 59496 79767
0 15438 5 1 1 90089
0 15439 7 1 2 67555 90090
0 15440 5 1 1 15439
0 15441 7 1 2 86695 15440
0 15442 5 1 1 15441
0 15443 7 1 2 76764 15442
0 15444 5 2 1 15443
0 15445 7 1 2 74257 71404
0 15446 5 1 1 15445
0 15447 7 1 2 90091 15446
0 15448 5 1 1 15447
0 15449 7 1 2 83580 15448
0 15450 5 1 1 15449
0 15451 7 1 2 15436 15450
0 15452 5 1 1 15451
0 15453 7 1 2 80859 15452
0 15454 5 1 1 15453
0 15455 7 1 2 15418 15454
0 15456 7 1 2 15411 15455
0 15457 5 1 1 15456
0 15458 7 1 2 68854 15457
0 15459 5 1 1 15458
0 15460 7 2 2 70767 83031
0 15461 5 5 1 90093
0 15462 7 1 2 84305 85898
0 15463 7 1 2 89741 15462
0 15464 7 1 2 87912 15463
0 15465 7 1 2 90095 15464
0 15466 5 1 1 15465
0 15467 7 1 2 15459 15466
0 15468 5 1 1 15467
0 15469 7 1 2 69105 15468
0 15470 5 1 1 15469
0 15471 7 3 2 60900 75046
0 15472 5 1 1 90100
0 15473 7 3 2 67272 90101
0 15474 5 1 1 90103
0 15475 7 1 2 62930 15474
0 15476 5 1 1 15475
0 15477 7 13 2 63944 89922
0 15478 7 12 2 60304 60473
0 15479 7 3 2 60101 90119
0 15480 7 3 2 81401 90131
0 15481 7 1 2 90106 90134
0 15482 7 1 2 15476 15481
0 15483 5 1 1 15482
0 15484 7 1 2 74650 86230
0 15485 7 11 2 60474 68303
0 15486 7 2 2 77546 90137
0 15487 5 1 1 90148
0 15488 7 1 2 88691 90149
0 15489 7 1 2 15484 15488
0 15490 5 1 1 15489
0 15491 7 1 2 15483 15490
0 15492 7 1 2 15470 15491
0 15493 5 1 1 15492
0 15494 7 1 2 71183 15493
0 15495 5 1 1 15494
0 15496 7 2 2 68304 74519
0 15497 5 1 1 90150
0 15498 7 12 2 67946 69176
0 15499 5 1 1 90152
0 15500 7 3 2 83342 90153
0 15501 5 1 1 90164
0 15502 7 1 2 15497 15501
0 15503 5 1 1 15502
0 15504 7 1 2 67041 15503
0 15505 5 1 1 15504
0 15506 7 1 2 80969 15505
0 15507 5 1 1 15506
0 15508 7 1 2 61281 15507
0 15509 5 1 1 15508
0 15510 7 2 2 67947 90021
0 15511 5 1 1 90167
0 15512 7 1 2 68305 90168
0 15513 5 1 1 15512
0 15514 7 1 2 15509 15513
0 15515 5 1 1 15514
0 15516 7 18 2 61479 90120
0 15517 5 2 1 90169
0 15518 7 2 2 72959 90170
0 15519 7 21 2 61687 68637
0 15520 5 1 1 90191
0 15521 7 6 2 63945 90192
0 15522 5 1 1 90212
0 15523 7 1 2 90189 90213
0 15524 7 1 2 15515 15523
0 15525 5 1 1 15524
0 15526 7 1 2 15495 15525
0 15527 7 1 2 15385 15526
0 15528 7 1 2 15240 15527
0 15529 5 1 1 15528
0 15530 7 1 2 69899 15529
0 15531 5 1 1 15530
0 15532 7 1 2 14709 15531
0 15533 7 1 2 14112 15532
0 15534 5 1 1 15533
0 15535 7 1 2 86780 15534
0 15536 5 1 1 15535
0 15537 7 1 2 81876 74664
0 15538 5 1 1 15537
0 15539 7 1 2 66220 15538
0 15540 5 1 1 15539
0 15541 7 1 2 62071 89384
0 15542 5 1 1 15541
0 15543 7 1 2 76665 15542
0 15544 5 1 1 15543
0 15545 7 2 2 65701 15544
0 15546 5 1 1 90218
0 15547 7 1 2 62576 81845
0 15548 5 1 1 15547
0 15549 7 1 2 15546 15548
0 15550 5 1 1 15549
0 15551 7 1 2 64252 15550
0 15552 5 1 1 15551
0 15553 7 2 2 65702 81846
0 15554 5 1 1 90220
0 15555 7 1 2 67273 72777
0 15556 5 3 1 15555
0 15557 7 2 2 74494 90222
0 15558 5 1 1 90225
0 15559 7 1 2 15554 15558
0 15560 5 1 1 15559
0 15561 7 1 2 62577 15560
0 15562 5 1 1 15561
0 15563 7 2 2 15552 15562
0 15564 7 1 2 15540 90227
0 15565 5 1 1 15564
0 15566 7 1 2 64696 15565
0 15567 5 1 1 15566
0 15568 7 2 2 66221 73459
0 15569 5 2 1 90229
0 15570 7 1 2 78620 78528
0 15571 5 2 1 15570
0 15572 7 1 2 90231 90233
0 15573 5 1 1 15572
0 15574 7 1 2 69153 15573
0 15575 5 1 1 15574
0 15576 7 2 2 69304 71596
0 15577 7 1 2 65985 83349
0 15578 5 2 1 15577
0 15579 7 1 2 90235 90237
0 15580 5 1 1 15579
0 15581 7 1 2 66222 15580
0 15582 5 1 1 15581
0 15583 7 2 2 61033 70982
0 15584 5 3 1 90239
0 15585 7 1 2 83815 76855
0 15586 5 1 1 15585
0 15587 7 1 2 90241 15586
0 15588 5 1 1 15587
0 15589 7 1 2 15582 15588
0 15590 7 1 2 15575 15589
0 15591 7 5 2 65986 76632
0 15592 5 1 1 90244
0 15593 7 1 2 61282 84581
0 15594 5 1 1 15593
0 15595 7 1 2 84094 15594
0 15596 5 1 1 15595
0 15597 7 1 2 15592 15596
0 15598 5 1 1 15597
0 15599 7 1 2 72585 15598
0 15600 5 1 1 15599
0 15601 7 1 2 74757 85418
0 15602 5 1 1 15601
0 15603 7 1 2 78037 84582
0 15604 5 2 1 15603
0 15605 7 1 2 64479 90249
0 15606 5 1 1 15605
0 15607 7 1 2 15602 15606
0 15608 5 1 1 15607
0 15609 7 1 2 69646 15608
0 15610 5 1 1 15609
0 15611 7 1 2 15600 15610
0 15612 7 1 2 15590 15611
0 15613 7 1 2 15567 15612
0 15614 5 1 1 15613
0 15615 7 1 2 64940 15614
0 15616 5 1 1 15615
0 15617 7 1 2 60793 82648
0 15618 5 2 1 15617
0 15619 7 2 2 65703 78529
0 15620 5 1 1 90253
0 15621 7 1 2 62276 90254
0 15622 5 1 1 15621
0 15623 7 1 2 81072 15622
0 15624 5 1 1 15623
0 15625 7 2 2 90251 15624
0 15626 5 1 1 90255
0 15627 7 1 2 64253 90256
0 15628 5 1 1 15627
0 15629 7 1 2 76089 89235
0 15630 5 1 1 15629
0 15631 7 1 2 15628 15630
0 15632 5 1 1 15631
0 15633 7 1 2 65837 15632
0 15634 5 1 1 15633
0 15635 7 2 2 73786 81421
0 15636 5 1 1 90257
0 15637 7 1 2 15634 15636
0 15638 5 1 1 15637
0 15639 7 1 2 64480 15638
0 15640 5 1 1 15639
0 15641 7 1 2 78425 87977
0 15642 5 2 1 15641
0 15643 7 1 2 73787 90259
0 15644 5 1 1 15643
0 15645 7 5 2 67556 74794
0 15646 5 6 1 90261
0 15647 7 1 2 69234 90266
0 15648 5 3 1 15647
0 15649 7 2 2 74138 88381
0 15650 5 2 1 90275
0 15651 7 1 2 82472 90276
0 15652 7 2 2 90272 15651
0 15653 5 1 1 90279
0 15654 7 1 2 65987 15653
0 15655 5 1 1 15654
0 15656 7 1 2 62578 90260
0 15657 5 1 1 15656
0 15658 7 1 2 15655 15657
0 15659 5 1 1 15658
0 15660 7 1 2 64697 15659
0 15661 5 1 1 15660
0 15662 7 1 2 15644 15661
0 15663 7 1 2 15640 15662
0 15664 5 1 1 15663
0 15665 7 1 2 66223 15664
0 15666 5 1 1 15665
0 15667 7 4 2 64254 65988
0 15668 5 1 1 90281
0 15669 7 1 2 67557 15668
0 15670 5 3 1 15669
0 15671 7 2 2 65838 73205
0 15672 5 1 1 90288
0 15673 7 1 2 90285 90289
0 15674 5 1 1 15673
0 15675 7 1 2 65989 73206
0 15676 5 1 1 15675
0 15677 7 1 2 67558 15676
0 15678 5 2 1 15677
0 15679 7 1 2 73809 81417
0 15680 5 1 1 15679
0 15681 7 1 2 90290 15680
0 15682 5 1 1 15681
0 15683 7 1 2 15674 15682
0 15684 5 1 1 15683
0 15685 7 1 2 66224 15684
0 15686 5 1 1 15685
0 15687 7 3 2 65990 76173
0 15688 5 2 1 90292
0 15689 7 1 2 73810 76856
0 15690 5 1 1 15689
0 15691 7 1 2 65704 15690
0 15692 5 1 1 15691
0 15693 7 1 2 90295 15692
0 15694 5 1 1 15693
0 15695 7 1 2 82303 15694
0 15696 5 1 1 15695
0 15697 7 1 2 66225 73039
0 15698 5 1 1 15697
0 15699 7 1 2 60794 15698
0 15700 5 1 1 15699
0 15701 7 1 2 65991 85419
0 15702 7 1 2 15700 15701
0 15703 5 1 1 15702
0 15704 7 1 2 15696 15703
0 15705 5 1 1 15704
0 15706 7 1 2 65839 15705
0 15707 5 1 1 15706
0 15708 7 1 2 15686 15707
0 15709 5 1 1 15708
0 15710 7 1 2 73865 15709
0 15711 5 1 1 15710
0 15712 7 1 2 15666 15711
0 15713 7 1 2 15616 15712
0 15714 5 1 1 15713
0 15715 7 1 2 85642 15714
0 15716 5 1 1 15715
0 15717 7 1 2 79882 76633
0 15718 7 1 2 81642 15717
0 15719 5 1 1 15718
0 15720 7 2 2 69647 76174
0 15721 5 1 1 90297
0 15722 7 1 2 78030 90298
0 15723 5 1 1 15722
0 15724 7 1 2 61480 15723
0 15725 5 1 1 15724
0 15726 7 1 2 60475 74637
0 15727 7 1 2 15725 15726
0 15728 5 1 1 15727
0 15729 7 1 2 15719 15728
0 15730 5 1 1 15729
0 15731 7 1 2 65840 15730
0 15732 5 1 1 15731
0 15733 7 3 2 64255 70405
0 15734 5 2 1 90299
0 15735 7 2 2 67559 78414
0 15736 5 1 1 90304
0 15737 7 1 2 90302 90305
0 15738 5 3 1 15737
0 15739 7 1 2 85442 90306
0 15740 5 1 1 15739
0 15741 7 1 2 15732 15740
0 15742 5 1 1 15741
0 15743 7 1 2 64481 15742
0 15744 5 1 1 15743
0 15745 7 1 2 61283 90280
0 15746 5 1 1 15745
0 15747 7 1 2 85443 15746
0 15748 5 1 1 15747
0 15749 7 1 2 15744 15748
0 15750 5 1 1 15749
0 15751 7 1 2 65154 15750
0 15752 5 1 1 15751
0 15753 7 3 2 60476 85037
0 15754 5 1 1 90309
0 15755 7 1 2 82116 90310
0 15756 7 1 2 74529 15755
0 15757 5 1 1 15756
0 15758 7 1 2 15752 15757
0 15759 5 1 1 15758
0 15760 7 1 2 77158 15759
0 15761 5 1 1 15760
0 15762 7 1 2 15716 15761
0 15763 5 1 1 15762
0 15764 7 1 2 63389 15763
0 15765 5 1 1 15764
0 15766 7 1 2 67560 81432
0 15767 5 3 1 15766
0 15768 7 1 2 71767 76199
0 15769 7 1 2 90312 15768
0 15770 5 1 1 15769
0 15771 7 4 2 64256 69452
0 15772 5 1 1 90315
0 15773 7 1 2 76200 90316
0 15774 5 2 1 15773
0 15775 7 1 2 62579 88348
0 15776 5 1 1 15775
0 15777 7 1 2 90319 15776
0 15778 7 1 2 15770 15777
0 15779 5 1 1 15778
0 15780 7 1 2 66226 15779
0 15781 5 1 1 15780
0 15782 7 1 2 74251 15781
0 15783 5 1 1 15782
0 15784 7 1 2 72712 15783
0 15785 5 1 1 15784
0 15786 7 3 2 67561 71543
0 15787 5 2 1 90321
0 15788 7 1 2 81677 86512
0 15789 5 1 1 15788
0 15790 7 1 2 2578 15789
0 15791 5 1 1 15790
0 15792 7 1 2 62580 15791
0 15793 5 1 1 15792
0 15794 7 1 2 90324 15793
0 15795 5 1 1 15794
0 15796 7 1 2 71768 15795
0 15797 5 1 1 15796
0 15798 7 7 2 62581 71544
0 15799 5 2 1 90326
0 15800 7 1 2 67042 90327
0 15801 5 1 1 15800
0 15802 7 3 2 65841 80584
0 15803 7 1 2 70525 76090
0 15804 5 1 1 15803
0 15805 7 1 2 90320 15804
0 15806 5 1 1 15805
0 15807 7 1 2 90335 15806
0 15808 5 1 1 15807
0 15809 7 1 2 15801 15808
0 15810 7 1 2 15797 15809
0 15811 5 1 1 15810
0 15812 7 1 2 72309 15811
0 15813 5 1 1 15812
0 15814 7 1 2 76175 78834
0 15815 5 1 1 15814
0 15816 7 1 2 90325 15815
0 15817 5 1 1 15816
0 15818 7 1 2 69648 15817
0 15819 5 1 1 15818
0 15820 7 1 2 73040 90322
0 15821 5 1 1 15820
0 15822 7 3 2 62582 76883
0 15823 7 1 2 72653 90338
0 15824 5 1 1 15823
0 15825 7 1 2 15821 15824
0 15826 7 1 2 15819 15825
0 15827 5 1 1 15826
0 15828 7 1 2 78656 15827
0 15829 5 1 1 15828
0 15830 7 1 2 76821 83835
0 15831 5 1 1 15830
0 15832 7 1 2 61284 81970
0 15833 5 1 1 15832
0 15834 7 1 2 15831 15833
0 15835 5 1 1 15834
0 15836 7 1 2 71099 15835
0 15837 5 1 1 15836
0 15838 7 5 2 65155 62072
0 15839 5 3 1 90341
0 15840 7 1 2 90342 88337
0 15841 5 1 1 15840
0 15842 7 1 2 15837 15841
0 15843 5 1 1 15842
0 15844 7 1 2 62583 15843
0 15845 5 1 1 15844
0 15846 7 1 2 82743 78456
0 15847 5 1 1 15846
0 15848 7 1 2 83656 15847
0 15849 5 1 1 15848
0 15850 7 1 2 70768 15849
0 15851 5 1 1 15850
0 15852 7 1 2 61481 15851
0 15853 7 1 2 15845 15852
0 15854 7 1 2 62277 79844
0 15855 5 1 1 15854
0 15856 7 2 2 61285 15855
0 15857 5 1 1 90349
0 15858 7 1 2 67562 15857
0 15859 5 1 1 15858
0 15860 7 2 2 76201 90267
0 15861 7 1 2 74060 90351
0 15862 5 1 1 15861
0 15863 7 1 2 15859 15862
0 15864 5 1 1 15863
0 15865 7 1 2 77183 15864
0 15866 5 1 1 15865
0 15867 7 2 2 67563 70769
0 15868 5 1 1 90353
0 15869 7 1 2 81666 15868
0 15870 5 1 1 15869
0 15871 7 1 2 85098 15870
0 15872 5 1 1 15871
0 15873 7 1 2 77184 76202
0 15874 7 1 2 83137 15873
0 15875 5 1 1 15874
0 15876 7 1 2 15872 15875
0 15877 5 1 1 15876
0 15878 7 1 2 69649 15877
0 15879 5 1 1 15878
0 15880 7 1 2 15866 15879
0 15881 7 1 2 15853 15880
0 15882 7 1 2 15829 15881
0 15883 7 1 2 15813 15882
0 15884 7 1 2 15785 15883
0 15885 5 1 1 15884
0 15886 7 2 2 60305 76203
0 15887 7 2 2 76995 71597
0 15888 7 5 2 71184 90357
0 15889 7 2 2 69235 76240
0 15890 5 1 1 90364
0 15891 7 1 2 88401 15890
0 15892 5 1 1 15891
0 15893 7 1 2 77048 15892
0 15894 5 1 1 15893
0 15895 7 1 2 90359 15894
0 15896 5 1 1 15895
0 15897 7 2 2 67564 15896
0 15898 5 1 1 90366
0 15899 7 1 2 62584 88561
0 15900 5 1 1 15899
0 15901 7 1 2 60102 15900
0 15902 7 1 2 15898 15901
0 15903 5 1 1 15902
0 15904 7 1 2 90355 15903
0 15905 5 1 1 15904
0 15906 7 1 2 69790 74061
0 15907 5 2 1 15906
0 15908 7 3 2 81827 90368
0 15909 5 1 1 90370
0 15910 7 1 2 61034 90371
0 15911 5 1 1 15910
0 15912 7 1 2 86963 15911
0 15913 5 1 1 15912
0 15914 7 1 2 62585 72977
0 15915 7 1 2 79116 15914
0 15916 5 1 1 15915
0 15917 7 1 2 15913 15916
0 15918 5 1 1 15917
0 15919 7 1 2 62073 15918
0 15920 5 1 1 15919
0 15921 7 1 2 74520 77625
0 15922 5 1 1 15921
0 15923 7 1 2 66227 76338
0 15924 7 1 2 77134 15923
0 15925 5 1 1 15924
0 15926 7 1 2 15922 15925
0 15927 5 1 1 15926
0 15928 7 1 2 72911 15927
0 15929 5 1 1 15928
0 15930 7 4 2 65842 77290
0 15931 5 3 1 90373
0 15932 7 1 2 82249 90377
0 15933 5 1 1 15932
0 15934 7 1 2 66439 15933
0 15935 7 1 2 15929 15934
0 15936 7 1 2 15920 15935
0 15937 7 1 2 15905 15936
0 15938 5 1 1 15937
0 15939 7 1 2 15885 15938
0 15940 5 1 1 15939
0 15941 7 1 2 63390 15940
0 15942 5 1 1 15941
0 15943 7 8 2 62586 75546
0 15944 5 3 1 90380
0 15945 7 2 2 76884 90381
0 15946 5 1 1 90391
0 15947 7 2 2 11074 90392
0 15948 7 1 2 64257 90393
0 15949 5 1 1 15948
0 15950 7 4 2 87230 90323
0 15951 5 1 1 90395
0 15952 7 1 2 15949 15951
0 15953 5 1 1 15952
0 15954 7 1 2 71769 15953
0 15955 5 1 1 15954
0 15956 7 1 2 86600 88803
0 15957 5 1 1 15956
0 15958 7 1 2 11701 15957
0 15959 5 1 1 15958
0 15960 7 1 2 75547 15959
0 15961 5 1 1 15960
0 15962 7 2 2 74249 85038
0 15963 5 1 1 90399
0 15964 7 1 2 15961 15963
0 15965 7 1 2 15955 15964
0 15966 5 1 1 15965
0 15967 7 1 2 72310 15966
0 15968 5 1 1 15967
0 15969 7 3 2 75548 77735
0 15970 5 2 1 90401
0 15971 7 2 2 75268 90404
0 15972 5 3 1 90406
0 15973 7 1 2 75965 88863
0 15974 5 3 1 15973
0 15975 7 1 2 76666 90411
0 15976 7 1 2 90408 15975
0 15977 5 1 1 15976
0 15978 7 1 2 15968 15977
0 15979 5 1 1 15978
0 15980 7 1 2 70309 15979
0 15981 5 1 1 15980
0 15982 7 1 2 64482 90394
0 15983 5 1 1 15982
0 15984 7 1 2 64258 90396
0 15985 5 1 1 15984
0 15986 7 1 2 15983 15985
0 15987 5 1 1 15986
0 15988 7 1 2 72311 15987
0 15989 5 1 1 15988
0 15990 7 2 2 70447 90400
0 15991 5 1 1 90414
0 15992 7 1 2 67565 10940
0 15993 5 2 1 15992
0 15994 7 1 2 76667 90416
0 15995 7 1 2 90402 15994
0 15996 5 1 1 15995
0 15997 7 1 2 15991 15996
0 15998 7 1 2 15989 15997
0 15999 5 1 1 15998
0 16000 7 1 2 70366 15999
0 16001 5 1 1 16000
0 16002 7 2 2 66440 77980
0 16003 7 2 2 76885 90418
0 16004 5 1 1 90420
0 16005 7 1 2 74014 85051
0 16006 7 1 2 83481 16005
0 16007 5 1 1 16006
0 16008 7 1 2 16004 16007
0 16009 5 1 1 16008
0 16010 7 1 2 74880 16009
0 16011 5 1 1 16010
0 16012 7 2 2 64259 74015
0 16013 7 1 2 90397 90422
0 16014 5 1 1 16013
0 16015 7 1 2 16011 16014
0 16016 5 1 1 16015
0 16017 7 1 2 88651 16016
0 16018 5 1 1 16017
0 16019 7 1 2 76004 72312
0 16020 5 1 1 16019
0 16021 7 2 2 62587 69365
0 16022 5 1 1 90424
0 16023 7 1 2 60103 16022
0 16024 7 1 2 16020 16023
0 16025 5 1 1 16024
0 16026 7 1 2 76668 16025
0 16027 5 1 1 16026
0 16028 7 1 2 82746 16027
0 16029 5 1 1 16028
0 16030 7 1 2 75190 16029
0 16031 5 1 1 16030
0 16032 7 1 2 82147 90423
0 16033 5 1 1 16032
0 16034 7 2 2 62588 80126
0 16035 5 1 1 90426
0 16036 7 2 2 16033 16035
0 16037 5 1 1 90428
0 16038 7 6 2 62074 75549
0 16039 7 4 2 65705 65992
0 16040 5 3 1 90436
0 16041 7 3 2 88329 90437
0 16042 7 1 2 90430 90443
0 16043 5 1 1 16042
0 16044 7 1 2 75269 16043
0 16045 5 1 1 16044
0 16046 7 1 2 16037 16045
0 16047 5 1 1 16046
0 16048 7 1 2 68306 16047
0 16049 7 1 2 16031 16048
0 16050 7 1 2 16018 16049
0 16051 7 1 2 16001 16050
0 16052 7 1 2 72183 72409
0 16053 5 1 1 16052
0 16054 7 1 2 72888 16053
0 16055 5 1 1 16054
0 16056 7 1 2 75270 16055
0 16057 5 1 1 16056
0 16058 7 1 2 76669 16057
0 16059 5 1 1 16058
0 16060 7 3 2 75904 78530
0 16061 5 3 1 90446
0 16062 7 1 2 60104 90449
0 16063 5 1 1 16062
0 16064 7 1 2 75271 76634
0 16065 5 1 1 16064
0 16066 7 1 2 90429 16065
0 16067 5 1 1 16066
0 16068 7 1 2 16063 16067
0 16069 5 1 1 16068
0 16070 7 1 2 16059 16069
0 16071 5 1 1 16070
0 16072 7 1 2 83466 16071
0 16073 5 1 1 16072
0 16074 7 2 2 64941 74847
0 16075 7 2 2 69366 70945
0 16076 5 2 1 90454
0 16077 7 1 2 90452 90455
0 16078 5 1 1 16077
0 16079 7 3 2 67566 72313
0 16080 5 1 1 90458
0 16081 7 1 2 71770 90459
0 16082 5 1 1 16081
0 16083 7 1 2 69650 80750
0 16084 5 1 1 16083
0 16085 7 1 2 62589 16084
0 16086 5 1 1 16085
0 16087 7 1 2 16082 16086
0 16088 5 1 1 16087
0 16089 7 1 2 66441 16088
0 16090 5 1 1 16089
0 16091 7 1 2 16078 16090
0 16092 5 1 1 16091
0 16093 7 1 2 65156 16092
0 16094 5 1 1 16093
0 16095 7 1 2 76176 74339
0 16096 7 1 2 90444 16095
0 16097 5 1 1 16096
0 16098 7 1 2 16094 16097
0 16099 5 1 1 16098
0 16100 7 1 2 62278 16099
0 16101 5 1 1 16100
0 16102 7 1 2 16073 16101
0 16103 7 1 2 16051 16102
0 16104 7 1 2 15981 16103
0 16105 5 1 1 16104
0 16106 7 1 2 65370 16105
0 16107 7 1 2 15942 16106
0 16108 5 1 1 16107
0 16109 7 1 2 68638 16108
0 16110 7 1 2 15765 16109
0 16111 5 1 1 16110
0 16112 7 1 2 75191 72967
0 16113 5 5 1 16112
0 16114 7 1 2 89541 90461
0 16115 5 1 1 16114
0 16116 7 3 2 67274 75272
0 16117 7 1 2 59838 90466
0 16118 5 1 1 16117
0 16119 7 1 2 16115 16118
0 16120 5 1 1 16119
0 16121 7 1 2 61286 16120
0 16122 5 1 1 16121
0 16123 7 1 2 73404 90467
0 16124 5 1 1 16123
0 16125 7 1 2 16122 16124
0 16126 5 1 1 16125
0 16127 7 1 2 80788 16126
0 16128 5 1 1 16127
0 16129 7 1 2 64698 73460
0 16130 5 1 1 16129
0 16131 7 1 2 65993 73291
0 16132 5 2 1 16131
0 16133 7 3 2 12782 90469
0 16134 7 1 2 16130 90471
0 16135 5 1 1 16134
0 16136 7 1 2 76740 16135
0 16137 5 1 1 16136
0 16138 7 1 2 71545 78531
0 16139 7 1 2 77256 16138
0 16140 5 1 1 16139
0 16141 7 1 2 16137 16140
0 16142 5 1 1 16141
0 16143 7 1 2 69236 16142
0 16144 5 1 1 16143
0 16145 7 1 2 70770 73980
0 16146 5 1 1 16145
0 16147 7 1 2 59839 16146
0 16148 5 1 1 16147
0 16149 7 2 2 61287 90378
0 16150 5 1 1 90474
0 16151 7 1 2 60105 90475
0 16152 5 1 1 16151
0 16153 7 4 2 16148 16152
0 16154 5 1 1 90476
0 16155 7 1 2 65157 90477
0 16156 5 1 1 16155
0 16157 7 1 2 73077 86289
0 16158 5 1 1 16157
0 16159 7 1 2 16156 16158
0 16160 5 1 1 16159
0 16161 7 1 2 73248 16160
0 16162 5 1 1 16161
0 16163 7 1 2 70142 12797
0 16164 5 1 1 16163
0 16165 7 1 2 76741 16164
0 16166 5 1 1 16165
0 16167 7 1 2 16162 16166
0 16168 7 1 2 16144 16167
0 16169 5 1 1 16168
0 16170 7 1 2 60477 16169
0 16171 5 1 1 16170
0 16172 7 1 2 16128 16171
0 16173 5 1 1 16172
0 16174 7 1 2 62590 16173
0 16175 5 1 1 16174
0 16176 7 1 2 70143 89207
0 16177 5 1 1 16176
0 16178 7 1 2 70899 16177
0 16179 5 2 1 16178
0 16180 7 1 2 77736 89192
0 16181 5 1 1 16180
0 16182 7 1 2 90480 16181
0 16183 5 1 1 16182
0 16184 7 1 2 80561 16183
0 16185 5 1 1 16184
0 16186 7 1 2 88611 89189
0 16187 5 1 1 16186
0 16188 7 1 2 88736 16187
0 16189 5 1 1 16188
0 16190 7 1 2 16185 16189
0 16191 7 1 2 16175 16190
0 16192 5 1 1 16191
0 16193 7 1 2 68307 16192
0 16194 5 1 1 16193
0 16195 7 2 2 73709 79162
0 16196 5 1 1 90482
0 16197 7 1 2 82519 72217
0 16198 5 1 1 16197
0 16199 7 1 2 67567 6004
0 16200 7 1 2 16198 16199
0 16201 5 1 1 16200
0 16202 7 1 2 16196 16201
0 16203 5 1 1 16202
0 16204 7 1 2 61288 16203
0 16205 5 1 1 16204
0 16206 7 3 2 60306 71367
0 16207 5 1 1 90484
0 16208 7 1 2 84127 73725
0 16209 5 1 1 16208
0 16210 7 1 2 72218 16209
0 16211 5 2 1 16210
0 16212 7 1 2 16207 90487
0 16213 7 1 2 16205 16212
0 16214 5 1 1 16213
0 16215 7 1 2 60478 16214
0 16216 5 1 1 16215
0 16217 7 1 2 69527 79163
0 16218 5 1 1 16217
0 16219 7 1 2 73595 16218
0 16220 5 1 1 16219
0 16221 7 1 2 73405 89852
0 16222 7 1 2 16220 16221
0 16223 5 1 1 16222
0 16224 7 1 2 16216 16223
0 16225 5 1 1 16224
0 16226 7 1 2 63391 16225
0 16227 5 1 1 16226
0 16228 7 5 2 59840 71870
0 16229 5 15 1 90489
0 16230 7 1 2 70771 90494
0 16231 5 1 1 16230
0 16232 7 1 2 81693 16231
0 16233 5 1 1 16232
0 16234 7 1 2 89212 16233
0 16235 5 1 1 16234
0 16236 7 1 2 70772 88971
0 16237 5 2 1 16236
0 16238 7 1 2 71518 90509
0 16239 5 1 1 16238
0 16240 7 1 2 89193 16239
0 16241 5 1 1 16240
0 16242 7 3 2 61035 70596
0 16243 7 3 2 82263 90511
0 16244 5 1 1 90514
0 16245 7 1 2 65158 16244
0 16246 5 1 1 16245
0 16247 7 1 2 59841 76143
0 16248 5 2 1 16247
0 16249 7 2 2 73847 90517
0 16250 7 2 2 88875 90519
0 16251 5 1 1 90521
0 16252 7 1 2 16246 16251
0 16253 7 1 2 16241 16252
0 16254 7 1 2 16235 16253
0 16255 5 1 1 16254
0 16256 7 1 2 90138 16255
0 16257 5 1 1 16256
0 16258 7 1 2 16227 16257
0 16259 5 1 1 16258
0 16260 7 1 2 66442 16259
0 16261 5 1 1 16260
0 16262 7 2 2 63392 89336
0 16263 7 1 2 71185 69969
0 16264 5 2 1 16263
0 16265 7 2 2 1240 90525
0 16266 5 2 1 90527
0 16267 7 1 2 79418 88422
0 16268 7 1 2 90529 16267
0 16269 5 2 1 16268
0 16270 7 1 2 70773 90531
0 16271 5 1 1 16270
0 16272 7 1 2 65994 81412
0 16273 5 1 1 16272
0 16274 7 1 2 70144 16273
0 16275 7 1 2 16271 16274
0 16276 5 1 1 16275
0 16277 7 1 2 76360 16276
0 16278 5 1 1 16277
0 16279 7 2 2 64942 81633
0 16280 5 3 1 90533
0 16281 7 2 2 76700 90245
0 16282 5 3 1 90538
0 16283 7 1 2 90535 90540
0 16284 5 1 1 16283
0 16285 7 1 2 64260 16284
0 16286 5 1 1 16285
0 16287 7 2 2 72568 82728
0 16288 7 1 2 73009 73923
0 16289 7 1 2 90543 16288
0 16290 5 1 1 16289
0 16291 7 1 2 65159 16290
0 16292 5 1 1 16291
0 16293 7 1 2 16286 16292
0 16294 7 2 2 76701 90293
0 16295 5 2 1 90545
0 16296 7 1 2 70145 90547
0 16297 5 1 1 16296
0 16298 7 1 2 74016 16297
0 16299 5 1 1 16298
0 16300 7 3 2 64699 90438
0 16301 5 1 1 90549
0 16302 7 1 2 69063 90550
0 16303 5 1 1 16302
0 16304 7 1 2 70146 16303
0 16305 5 1 1 16304
0 16306 7 1 2 62591 16305
0 16307 5 1 1 16306
0 16308 7 1 2 16299 16307
0 16309 7 1 2 16293 16308
0 16310 7 1 2 84052 77271
0 16311 5 2 1 16310
0 16312 7 1 2 88171 90552
0 16313 5 1 1 16312
0 16314 7 1 2 83812 73375
0 16315 5 2 1 16314
0 16316 7 1 2 70147 90554
0 16317 7 1 2 16313 16316
0 16318 5 1 1 16317
0 16319 7 1 2 72314 16318
0 16320 5 1 1 16319
0 16321 7 1 2 70971 85982
0 16322 5 1 1 16321
0 16323 7 1 2 70895 16322
0 16324 5 1 1 16323
0 16325 7 1 2 90277 16324
0 16326 5 1 1 16325
0 16327 7 1 2 16320 16326
0 16328 7 1 2 16309 16327
0 16329 7 1 2 65843 72436
0 16330 5 3 1 16329
0 16331 7 1 2 71186 90556
0 16332 5 1 1 16331
0 16333 7 1 2 62592 16332
0 16334 5 1 1 16333
0 16335 7 1 2 71187 76224
0 16336 5 2 1 16335
0 16337 7 1 2 74017 90559
0 16338 5 1 1 16337
0 16339 7 1 2 83816 16301
0 16340 5 1 1 16339
0 16341 7 1 2 64261 16340
0 16342 5 1 1 16341
0 16343 7 1 2 16338 16342
0 16344 7 2 2 16334 16343
0 16345 5 1 1 90561
0 16346 7 1 2 70774 16345
0 16347 5 1 1 16346
0 16348 7 1 2 73224 70900
0 16349 5 1 1 16348
0 16350 7 2 2 69651 73242
0 16351 7 1 2 74230 90563
0 16352 5 1 1 16351
0 16353 7 1 2 16349 16352
0 16354 5 1 1 16353
0 16355 7 1 2 69237 16354
0 16356 5 1 1 16355
0 16357 7 1 2 16347 16356
0 16358 7 1 2 16328 16357
0 16359 7 1 2 16278 16358
0 16360 5 1 1 16359
0 16361 7 1 2 90523 16360
0 16362 5 1 1 16361
0 16363 7 2 2 65371 80808
0 16364 5 2 1 90565
0 16365 7 4 2 62593 75273
0 16366 7 1 2 69721 90569
0 16367 5 1 1 16366
0 16368 7 1 2 12217 16367
0 16369 5 2 1 16368
0 16370 7 1 2 90566 90573
0 16371 5 1 1 16370
0 16372 7 5 2 60479 80020
0 16373 5 2 1 90575
0 16374 7 1 2 73622 81486
0 16375 5 2 1 16374
0 16376 7 1 2 90576 90582
0 16377 5 1 1 16376
0 16378 7 1 2 16371 16377
0 16379 5 1 1 16378
0 16380 7 1 2 72912 16379
0 16381 5 1 1 16380
0 16382 7 1 2 82167 89482
0 16383 5 1 1 16382
0 16384 7 2 2 90580 16383
0 16385 5 1 1 90584
0 16386 7 1 2 65372 75109
0 16387 5 2 1 16386
0 16388 7 1 2 85755 90586
0 16389 5 1 1 16388
0 16390 7 1 2 88612 16389
0 16391 5 1 1 16390
0 16392 7 1 2 90585 16391
0 16393 5 1 1 16392
0 16394 7 1 2 81484 16393
0 16395 5 1 1 16394
0 16396 7 5 2 59842 74860
0 16397 7 1 2 73615 90588
0 16398 7 1 2 89910 16397
0 16399 5 1 1 16398
0 16400 7 1 2 16395 16399
0 16401 5 1 1 16400
0 16402 7 1 2 61289 16401
0 16403 5 1 1 16402
0 16404 7 1 2 16381 16403
0 16405 5 1 1 16404
0 16406 7 1 2 72094 16405
0 16407 5 1 1 16406
0 16408 7 2 2 67568 83697
0 16409 5 1 1 90593
0 16410 7 1 2 77602 90594
0 16411 5 1 1 16410
0 16412 7 1 2 62594 73710
0 16413 7 1 2 16385 16412
0 16414 5 1 1 16413
0 16415 7 1 2 16411 16414
0 16416 5 1 1 16415
0 16417 7 1 2 71706 16416
0 16418 5 1 1 16417
0 16419 7 21 2 60480 63393
0 16420 5 7 1 90595
0 16421 7 2 2 62595 74340
0 16422 5 1 1 90623
0 16423 7 1 2 90596 90624
0 16424 5 1 1 16423
0 16425 7 1 2 71004 85444
0 16426 5 1 1 16425
0 16427 7 1 2 83273 83698
0 16428 5 1 1 16427
0 16429 7 1 2 16426 16428
0 16430 5 1 1 16429
0 16431 7 1 2 77135 16430
0 16432 5 1 1 16431
0 16433 7 1 2 16424 16432
0 16434 7 1 2 16418 16433
0 16435 5 1 1 16434
0 16436 7 1 2 72913 16435
0 16437 5 1 1 16436
0 16438 7 1 2 63694 16437
0 16439 7 1 2 16407 16438
0 16440 7 1 2 16362 16439
0 16441 7 1 2 16261 16440
0 16442 7 1 2 16194 16441
0 16443 5 1 1 16442
0 16444 7 1 2 16111 16443
0 16445 5 1 1 16444
0 16446 7 1 2 79942 84991
0 16447 5 1 1 16446
0 16448 7 1 2 65160 16447
0 16449 5 1 1 16448
0 16450 7 1 2 80021 88677
0 16451 5 1 1 16450
0 16452 7 1 2 16449 16451
0 16453 5 1 1 16452
0 16454 7 1 2 84176 16453
0 16455 5 1 1 16454
0 16456 7 2 2 63695 70148
0 16457 7 1 2 90577 90625
0 16458 7 1 2 88721 16457
0 16459 5 1 1 16458
0 16460 7 1 2 62596 16459
0 16461 7 1 2 16455 16460
0 16462 5 1 1 16461
0 16463 7 1 2 85899 89646
0 16464 5 1 1 16463
0 16465 7 1 2 79965 83699
0 16466 5 1 1 16465
0 16467 7 1 2 90581 16466
0 16468 5 1 1 16467
0 16469 7 1 2 82551 16468
0 16470 5 1 1 16469
0 16471 7 1 2 16464 16470
0 16472 5 1 1 16471
0 16473 7 1 2 66228 16472
0 16474 5 1 1 16473
0 16475 7 5 2 60481 62279
0 16476 7 1 2 60106 90627
0 16477 5 1 1 16476
0 16478 7 1 2 65373 81799
0 16479 5 14 1 16478
0 16480 7 1 2 81930 72184
0 16481 7 1 2 90632 16480
0 16482 5 1 1 16481
0 16483 7 1 2 16477 16482
0 16484 5 1 1 16483
0 16485 7 1 2 80022 16484
0 16486 5 1 1 16485
0 16487 7 1 2 16474 16486
0 16488 5 1 1 16487
0 16489 7 1 2 63696 16488
0 16490 5 1 1 16489
0 16491 7 3 2 59497 89647
0 16492 7 1 2 83576 90646
0 16493 5 1 1 16492
0 16494 7 1 2 67569 16493
0 16495 7 1 2 16490 16494
0 16496 5 1 1 16495
0 16497 7 1 2 71188 16496
0 16498 7 1 2 16462 16497
0 16499 5 1 1 16498
0 16500 7 1 2 16445 16499
0 16501 5 1 1 16500
0 16502 7 1 2 62931 16501
0 16503 5 1 1 16502
0 16504 7 1 2 67043 90583
0 16505 5 1 1 16504
0 16506 7 1 2 76028 16505
0 16507 5 1 1 16506
0 16508 7 1 2 66229 16507
0 16509 5 1 1 16508
0 16510 7 1 2 67570 75765
0 16511 5 1 1 16510
0 16512 7 1 2 16509 16511
0 16513 5 1 1 16512
0 16514 7 1 2 72095 16513
0 16515 5 1 1 16514
0 16516 7 1 2 69528 78031
0 16517 5 1 1 16516
0 16518 7 1 2 65995 73565
0 16519 5 3 1 16518
0 16520 7 3 2 61290 74718
0 16521 5 2 1 90652
0 16522 7 2 2 90649 90653
0 16523 7 1 2 60107 90657
0 16524 5 4 1 16523
0 16525 7 1 2 81678 90659
0 16526 5 1 1 16525
0 16527 7 1 2 16517 16526
0 16528 5 1 1 16527
0 16529 7 1 2 67044 16528
0 16530 5 1 1 16529
0 16531 7 1 2 66230 78725
0 16532 5 1 1 16531
0 16533 7 1 2 3859 16532
0 16534 7 1 2 16530 16533
0 16535 5 1 1 16534
0 16536 7 1 2 67571 16535
0 16537 5 1 1 16536
0 16538 7 2 2 16515 16537
0 16539 7 1 2 74588 88901
0 16540 5 1 1 16539
0 16541 7 1 2 13765 16540
0 16542 5 1 1 16541
0 16543 7 1 2 62597 16542
0 16544 5 1 1 16543
0 16545 7 1 2 66231 16544
0 16546 5 2 1 16545
0 16547 7 1 2 64483 88403
0 16548 5 1 1 16547
0 16549 7 1 2 71485 16548
0 16550 5 1 1 16549
0 16551 7 1 2 88408 16550
0 16552 5 1 1 16551
0 16553 7 2 2 90360 16552
0 16554 7 1 2 70597 90667
0 16555 5 1 1 16554
0 16556 7 1 2 62598 16555
0 16557 5 1 1 16556
0 16558 7 2 2 82570 72315
0 16559 5 1 1 90669
0 16560 7 1 2 72668 16559
0 16561 5 1 1 16560
0 16562 7 1 2 71451 16561
0 16563 5 1 1 16562
0 16564 7 1 2 80603 78106
0 16565 5 2 1 16564
0 16566 7 1 2 72914 89378
0 16567 7 1 2 90671 16566
0 16568 7 1 2 16563 16567
0 16569 7 1 2 16557 16568
0 16570 5 1 1 16569
0 16571 7 1 2 90665 16570
0 16572 5 1 1 16571
0 16573 7 1 2 90663 16572
0 16574 5 1 1 16573
0 16575 7 1 2 66443 16574
0 16576 5 1 1 16575
0 16577 7 1 2 71546 88358
0 16578 5 1 1 16577
0 16579 7 1 2 76765 16578
0 16580 5 1 1 16579
0 16581 7 1 2 81680 16580
0 16582 5 2 1 16581
0 16583 7 1 2 16576 90673
0 16584 5 1 1 16583
0 16585 7 4 2 63697 90597
0 16586 7 1 2 16584 90675
0 16587 5 1 1 16586
0 16588 7 2 2 65161 79768
0 16589 5 3 1 90679
0 16590 7 2 2 62599 76840
0 16591 7 1 2 65162 80727
0 16592 5 3 1 16591
0 16593 7 1 2 79805 90686
0 16594 5 1 1 16593
0 16595 7 1 2 69791 16594
0 16596 5 1 1 16595
0 16597 7 1 2 84750 16596
0 16598 5 1 1 16597
0 16599 7 1 2 90684 16598
0 16600 5 1 1 16599
0 16601 7 1 2 90681 16600
0 16602 5 1 1 16601
0 16603 7 1 2 64943 16602
0 16604 5 1 1 16603
0 16605 7 2 2 84076 76841
0 16606 7 1 2 77348 90689
0 16607 5 1 1 16606
0 16608 7 1 2 60108 78038
0 16609 5 1 1 16608
0 16610 7 1 2 65163 69979
0 16611 7 1 2 16609 16610
0 16612 5 1 1 16611
0 16613 7 1 2 16607 16612
0 16614 5 1 1 16613
0 16615 7 1 2 68308 16614
0 16616 5 1 1 16615
0 16617 7 1 2 74277 83827
0 16618 5 1 1 16617
0 16619 7 1 2 77027 16618
0 16620 5 1 1 16619
0 16621 7 1 2 74990 16620
0 16622 5 1 1 16621
0 16623 7 1 2 16616 16622
0 16624 5 1 1 16623
0 16625 7 1 2 66444 16624
0 16626 5 1 1 16625
0 16627 7 1 2 86929 11138
0 16628 5 1 1 16627
0 16629 7 1 2 64944 16628
0 16630 5 1 1 16629
0 16631 7 1 2 75415 77603
0 16632 5 1 1 16631
0 16633 7 1 2 85736 16632
0 16634 5 1 1 16633
0 16635 7 1 2 65164 16634
0 16636 5 1 1 16635
0 16637 7 5 2 62280 75682
0 16638 5 1 1 90691
0 16639 7 1 2 86668 90692
0 16640 5 1 1 16639
0 16641 7 1 2 16636 16640
0 16642 7 1 2 16630 16641
0 16643 5 1 1 16642
0 16644 7 1 2 69652 16643
0 16645 5 1 1 16644
0 16646 7 3 2 65706 88247
0 16647 7 1 2 83174 90696
0 16648 5 1 1 16647
0 16649 7 1 2 65165 9459
0 16650 5 1 1 16649
0 16651 7 2 2 60307 80047
0 16652 5 2 1 90699
0 16653 7 1 2 85420 90701
0 16654 7 1 2 16650 16653
0 16655 5 1 1 16654
0 16656 7 1 2 16648 16655
0 16657 7 1 2 16645 16656
0 16658 7 1 2 16626 16657
0 16659 7 1 2 16604 16658
0 16660 5 1 1 16659
0 16661 7 1 2 68639 16660
0 16662 5 1 1 16661
0 16663 7 3 2 83660 85900
0 16664 7 2 2 62600 78344
0 16665 5 2 1 90706
0 16666 7 1 2 90703 90707
0 16667 5 1 1 16666
0 16668 7 1 2 16662 16667
0 16669 5 1 1 16668
0 16670 7 1 2 72316 16669
0 16671 5 1 1 16670
0 16672 7 1 2 64262 75831
0 16673 5 1 1 16672
0 16674 7 1 2 79806 16673
0 16675 5 2 1 16674
0 16676 7 1 2 65166 90710
0 16677 5 1 1 16676
0 16678 7 1 2 80023 88429
0 16679 5 1 1 16678
0 16680 7 1 2 16677 16679
0 16681 5 1 1 16680
0 16682 7 1 2 69453 16681
0 16683 5 1 1 16682
0 16684 7 5 2 65167 85039
0 16685 5 2 1 90712
0 16686 7 1 2 81532 90713
0 16687 5 1 1 16686
0 16688 7 1 2 75149 12098
0 16689 5 1 1 16688
0 16690 7 1 2 63394 82304
0 16691 7 1 2 16689 16690
0 16692 5 1 1 16691
0 16693 7 1 2 62601 82514
0 16694 5 1 1 16693
0 16695 7 1 2 16692 16694
0 16696 5 1 1 16695
0 16697 7 1 2 70310 16696
0 16698 5 1 1 16697
0 16699 7 1 2 16687 16698
0 16700 7 1 2 16683 16699
0 16701 5 1 1 16700
0 16702 7 1 2 68640 16701
0 16703 5 1 1 16702
0 16704 7 1 2 78345 90704
0 16705 5 1 1 16704
0 16706 7 1 2 16703 16705
0 16707 5 1 1 16706
0 16708 7 1 2 72713 16707
0 16709 5 1 1 16708
0 16710 7 5 2 65996 81533
0 16711 7 2 2 77072 90719
0 16712 5 1 1 90724
0 16713 7 1 2 65168 90725
0 16714 5 1 1 16713
0 16715 7 3 2 63395 75875
0 16716 7 1 2 82305 90726
0 16717 5 1 1 16716
0 16718 7 3 2 64263 63396
0 16719 5 3 1 90729
0 16720 7 1 2 81253 90730
0 16721 5 1 1 16720
0 16722 7 1 2 87684 16721
0 16723 5 1 1 16722
0 16724 7 1 2 77185 16723
0 16725 5 1 1 16724
0 16726 7 1 2 16717 16725
0 16727 7 1 2 16714 16726
0 16728 5 1 1 16727
0 16729 7 1 2 70311 16728
0 16730 5 1 1 16729
0 16731 7 1 2 77186 90711
0 16732 5 1 1 16731
0 16733 7 2 2 64264 77073
0 16734 7 4 2 68309 77144
0 16735 7 1 2 90735 90737
0 16736 5 1 1 16735
0 16737 7 1 2 85756 16736
0 16738 7 1 2 16732 16737
0 16739 5 1 1 16738
0 16740 7 1 2 69454 16739
0 16741 5 1 1 16740
0 16742 7 1 2 75274 77841
0 16743 5 1 1 16742
0 16744 7 1 2 80728 90382
0 16745 7 1 2 16743 16744
0 16746 5 1 1 16745
0 16747 7 1 2 16741 16746
0 16748 7 1 2 16730 16747
0 16749 5 1 1 16748
0 16750 7 1 2 83648 16749
0 16751 5 1 1 16750
0 16752 7 1 2 74678 82315
0 16753 7 1 2 86001 16752
0 16754 5 1 1 16753
0 16755 7 1 2 16751 16754
0 16756 7 1 2 16709 16755
0 16757 7 1 2 16671 16756
0 16758 5 1 1 16757
0 16759 7 1 2 71771 16758
0 16760 5 1 1 16759
0 16761 7 1 2 72714 79173
0 16762 5 1 1 16761
0 16763 7 1 2 66232 16762
0 16764 5 1 1 16763
0 16765 7 1 2 72669 74469
0 16766 5 1 1 16765
0 16767 7 1 2 60308 16766
0 16768 5 1 1 16767
0 16769 7 1 2 16764 16768
0 16770 5 1 1 16769
0 16771 7 1 2 62075 16770
0 16772 5 1 1 16771
0 16773 7 1 2 67045 88806
0 16774 5 1 1 16773
0 16775 7 1 2 78810 16774
0 16776 5 1 1 16775
0 16777 7 1 2 69980 16776
0 16778 5 1 1 16777
0 16779 7 1 2 62602 16778
0 16780 7 1 2 16772 16779
0 16781 5 1 1 16780
0 16782 7 1 2 65169 78102
0 16783 5 1 1 16782
0 16784 7 1 2 71969 78346
0 16785 5 2 1 16784
0 16786 7 1 2 77169 90741
0 16787 5 1 1 16786
0 16788 7 1 2 88807 16787
0 16789 5 1 1 16788
0 16790 7 1 2 67572 16789
0 16791 7 1 2 16783 16790
0 16792 5 1 1 16791
0 16793 7 1 2 16781 16792
0 16794 5 1 1 16793
0 16795 7 1 2 72670 90742
0 16796 5 1 1 16795
0 16797 7 1 2 78805 16796
0 16798 5 1 1 16797
0 16799 7 2 2 64945 71848
0 16800 5 1 1 90743
0 16801 7 1 2 66233 84970
0 16802 5 1 1 16801
0 16803 7 1 2 83657 16802
0 16804 5 1 1 16803
0 16805 7 1 2 16800 16804
0 16806 5 1 1 16805
0 16807 7 1 2 77170 72819
0 16808 5 1 1 16807
0 16809 7 1 2 66445 16808
0 16810 7 1 2 16806 16809
0 16811 7 1 2 16798 16810
0 16812 7 1 2 16794 16811
0 16813 5 1 1 16812
0 16814 7 3 2 70483 82138
0 16815 5 2 1 90745
0 16816 7 1 2 65997 83506
0 16817 5 2 1 16816
0 16818 7 1 2 90748 90750
0 16819 5 1 1 16818
0 16820 7 1 2 71970 16819
0 16821 5 1 1 16820
0 16822 7 2 2 62603 76526
0 16823 5 1 1 90752
0 16824 7 1 2 71100 90753
0 16825 5 1 1 16824
0 16826 7 1 2 16821 16825
0 16827 5 1 1 16826
0 16828 7 1 2 71547 16827
0 16829 5 1 1 16828
0 16830 7 1 2 60309 70991
0 16831 5 1 1 16830
0 16832 7 1 2 71101 16831
0 16833 5 1 1 16832
0 16834 7 1 2 62076 81822
0 16835 5 2 1 16834
0 16836 7 1 2 69970 90754
0 16837 5 1 1 16836
0 16838 7 1 2 65170 76005
0 16839 7 1 2 16837 16838
0 16840 5 1 1 16839
0 16841 7 1 2 16833 16840
0 16842 5 1 1 16841
0 16843 7 1 2 70775 16842
0 16844 5 1 1 16843
0 16845 7 1 2 87228 16844
0 16846 7 1 2 16829 16845
0 16847 5 1 1 16846
0 16848 7 1 2 63397 16847
0 16849 7 1 2 16813 16848
0 16850 5 1 1 16849
0 16851 7 2 2 65707 84980
0 16852 5 1 1 90756
0 16853 7 1 2 76670 16852
0 16854 5 1 1 16853
0 16855 7 1 2 64265 16854
0 16856 5 1 1 16855
0 16857 7 1 2 76097 78896
0 16858 5 1 1 16857
0 16859 7 1 2 62281 16858
0 16860 5 1 1 16859
0 16861 7 1 2 8800 16860
0 16862 7 1 2 12365 16861
0 16863 7 1 2 16856 16862
0 16864 5 1 1 16863
0 16865 7 2 2 87231 88540
0 16866 7 3 2 70776 75192
0 16867 5 20 1 90760
0 16868 7 3 2 71189 90763
0 16869 5 2 1 90783
0 16870 7 1 2 90758 90786
0 16871 7 1 2 16864 16870
0 16872 5 1 1 16871
0 16873 7 1 2 16850 16872
0 16874 5 1 1 16873
0 16875 7 1 2 68641 16874
0 16876 5 1 1 16875
0 16877 7 5 2 67573 72941
0 16878 5 2 1 90788
0 16879 7 1 2 65171 90793
0 16880 5 4 1 16879
0 16881 7 1 2 81218 90795
0 16882 5 1 1 16881
0 16883 7 1 2 66446 83412
0 16884 5 1 1 16883
0 16885 7 1 2 79979 72410
0 16886 5 1 1 16885
0 16887 7 1 2 682 16886
0 16888 5 1 1 16887
0 16889 7 1 2 69529 16888
0 16890 5 1 1 16889
0 16891 7 1 2 72942 86964
0 16892 5 3 1 16891
0 16893 7 1 2 16890 90799
0 16894 5 1 1 16893
0 16895 7 1 2 63398 16894
0 16896 5 1 1 16895
0 16897 7 2 2 62282 71306
0 16898 5 1 1 90802
0 16899 7 1 2 84910 89171
0 16900 5 1 1 16899
0 16901 7 1 2 90803 16900
0 16902 5 1 1 16901
0 16903 7 1 2 72715 76006
0 16904 5 1 1 16903
0 16905 7 1 2 16902 16904
0 16906 5 1 1 16905
0 16907 7 1 2 68310 16906
0 16908 5 1 1 16907
0 16909 7 1 2 16896 16908
0 16910 5 1 1 16909
0 16911 7 1 2 16884 16910
0 16912 5 1 1 16911
0 16913 7 1 2 16882 16912
0 16914 5 1 1 16913
0 16915 7 1 2 61291 16914
0 16916 5 1 1 16915
0 16917 7 5 2 76493 89130
0 16918 7 1 2 80927 74915
0 16919 7 1 2 90804 16918
0 16920 5 1 1 16919
0 16921 7 1 2 78310 89353
0 16922 5 1 1 16921
0 16923 7 1 2 16922 89359
0 16924 7 1 2 16920 16923
0 16925 5 1 1 16924
0 16926 7 1 2 68311 16925
0 16927 5 1 1 16926
0 16928 7 1 2 89354 89617
0 16929 5 1 1 16928
0 16930 7 4 2 59304 60109
0 16931 7 2 2 89742 90809
0 16932 7 1 2 73060 73960
0 16933 7 1 2 90813 16932
0 16934 5 1 1 16933
0 16935 7 1 2 16929 16934
0 16936 5 1 1 16935
0 16937 7 1 2 71190 16936
0 16938 5 1 1 16937
0 16939 7 1 2 88902 89105
0 16940 5 1 1 16939
0 16941 7 1 2 82606 72978
0 16942 5 1 1 16941
0 16943 7 1 2 16940 16942
0 16944 5 1 1 16943
0 16945 7 1 2 63399 71707
0 16946 7 1 2 16944 16945
0 16947 5 1 1 16946
0 16948 7 1 2 16938 16947
0 16949 7 1 2 16927 16948
0 16950 7 1 2 16916 16949
0 16951 5 1 1 16950
0 16952 7 1 2 63698 16951
0 16953 5 1 1 16952
0 16954 7 1 2 16876 16953
0 16955 7 1 2 16760 16954
0 16956 7 1 2 81508 89373
0 16957 5 1 1 16956
0 16958 7 1 2 62283 16957
0 16959 5 1 1 16958
0 16960 7 2 2 84911 16959
0 16961 5 1 1 90815
0 16962 7 1 2 60110 90816
0 16963 5 1 1 16962
0 16964 7 1 2 90705 16963
0 16965 5 1 1 16964
0 16966 7 1 2 71971 90328
0 16967 5 1 1 16966
0 16968 7 1 2 76766 16967
0 16969 5 1 1 16968
0 16970 7 1 2 61482 16969
0 16971 5 1 1 16970
0 16972 7 1 2 71972 75095
0 16973 5 2 1 16972
0 16974 7 1 2 88790 90817
0 16975 5 1 1 16974
0 16976 7 1 2 90419 16975
0 16977 5 1 1 16976
0 16978 7 1 2 16971 16977
0 16979 5 1 1 16978
0 16980 7 1 2 63400 16979
0 16981 5 1 1 16980
0 16982 7 2 2 73348 70946
0 16983 5 2 1 90819
0 16984 7 1 2 90759 90820
0 16985 5 1 1 16984
0 16986 7 1 2 16981 16985
0 16987 5 1 1 16986
0 16988 7 1 2 69981 16987
0 16989 5 1 1 16988
0 16990 7 1 2 79924 85010
0 16991 5 1 1 16990
0 16992 7 2 2 68312 76635
0 16993 7 1 2 71973 74658
0 16994 7 1 2 90823 16993
0 16995 5 1 1 16994
0 16996 7 1 2 16991 16995
0 16997 5 1 1 16996
0 16998 7 1 2 65172 16997
0 16999 5 1 1 16998
0 17000 7 1 2 82117 90824
0 17001 5 1 1 17000
0 17002 7 2 2 62077 73911
0 17003 5 1 1 90825
0 17004 7 1 2 63401 90826
0 17005 5 1 1 17004
0 17006 7 1 2 17001 17005
0 17007 5 1 1 17006
0 17008 7 1 2 64946 17007
0 17009 5 1 1 17008
0 17010 7 1 2 71005 78806
0 17011 5 1 1 17010
0 17012 7 1 2 17009 17011
0 17013 5 1 1 17012
0 17014 7 1 2 66447 17013
0 17015 5 1 1 17014
0 17016 7 1 2 16999 17015
0 17017 5 1 1 17016
0 17018 7 1 2 69653 17017
0 17019 5 1 1 17018
0 17020 7 1 2 79226 88304
0 17021 5 1 1 17020
0 17022 7 1 2 62078 17021
0 17023 5 1 1 17022
0 17024 7 1 2 71034 17023
0 17025 5 1 1 17024
0 17026 7 1 2 61483 17025
0 17027 5 1 1 17026
0 17028 7 1 2 67275 80431
0 17029 5 1 1 17028
0 17030 7 1 2 76022 17029
0 17031 5 1 1 17030
0 17032 7 1 2 74341 17031
0 17033 5 1 1 17032
0 17034 7 1 2 61292 82319
0 17035 5 1 1 17034
0 17036 7 1 2 79524 17035
0 17037 5 1 1 17036
0 17038 7 1 2 17033 17037
0 17039 7 1 2 17027 17038
0 17040 5 1 1 17039
0 17041 7 1 2 75683 17040
0 17042 5 1 1 17041
0 17043 7 1 2 75995 16898
0 17044 5 1 1 17043
0 17045 7 1 2 75832 76742
0 17046 7 1 2 17044 17045
0 17047 5 1 1 17046
0 17048 7 1 2 17042 17047
0 17049 7 1 2 17019 17048
0 17050 7 1 2 16989 17049
0 17051 5 1 1 17050
0 17052 7 1 2 68642 17051
0 17053 5 1 1 17052
0 17054 7 1 2 16965 17053
0 17055 5 1 1 17054
0 17056 7 1 2 72317 17055
0 17057 5 1 1 17056
0 17058 7 3 2 62079 72915
0 17059 5 1 1 90827
0 17060 7 2 2 71191 69722
0 17061 5 1 1 90830
0 17062 7 1 2 62284 90831
0 17063 5 1 1 17062
0 17064 7 1 2 17059 17063
0 17065 5 1 1 17064
0 17066 7 1 2 73163 17065
0 17067 5 1 1 17066
0 17068 7 1 2 66234 76599
0 17069 5 1 1 17068
0 17070 7 1 2 65173 17069
0 17071 5 1 1 17070
0 17072 7 1 2 17067 17071
0 17073 5 1 1 17072
0 17074 7 1 2 89765 17073
0 17075 5 1 1 17074
0 17076 7 1 2 66235 74646
0 17077 5 1 1 17076
0 17078 7 1 2 60310 17077
0 17079 5 1 1 17078
0 17080 7 1 2 66236 4378
0 17081 5 1 1 17080
0 17082 7 1 2 61484 17081
0 17083 5 1 1 17082
0 17084 7 1 2 17079 17083
0 17085 5 1 1 17084
0 17086 7 1 2 61036 17085
0 17087 5 1 1 17086
0 17088 7 1 2 59843 82754
0 17089 5 1 1 17088
0 17090 7 1 2 17087 17089
0 17091 5 1 1 17090
0 17092 7 1 2 60111 17091
0 17093 5 1 1 17092
0 17094 7 1 2 7128 17093
0 17095 5 1 1 17094
0 17096 7 1 2 63699 17095
0 17097 5 1 1 17096
0 17098 7 1 2 17075 17097
0 17099 5 1 1 17098
0 17100 7 1 2 63402 17099
0 17101 5 1 1 17100
0 17102 7 1 2 59844 89355
0 17103 5 1 1 17102
0 17104 7 1 2 74731 73406
0 17105 5 1 1 17104
0 17106 7 1 2 81067 17105
0 17107 5 2 1 17106
0 17108 7 1 2 61037 90832
0 17109 5 1 1 17108
0 17110 7 1 2 17109 14999
0 17111 7 1 2 17103 17110
0 17112 5 1 1 17111
0 17113 7 1 2 69530 17112
0 17114 5 1 1 17113
0 17115 7 3 2 71192 89356
0 17116 5 1 1 90834
0 17117 7 1 2 67276 90835
0 17118 5 1 1 17117
0 17119 7 1 2 17114 17118
0 17120 5 1 1 17119
0 17121 7 1 2 78747 17120
0 17122 5 1 1 17121
0 17123 7 1 2 17101 17122
0 17124 5 1 1 17123
0 17125 7 1 2 72096 17124
0 17126 5 1 1 17125
0 17127 7 1 2 17057 17126
0 17128 7 1 2 16955 17127
0 17129 5 1 1 17128
0 17130 7 1 2 65374 17129
0 17131 5 1 1 17130
0 17132 7 1 2 16587 17131
0 17133 5 1 1 17132
0 17134 7 1 2 67948 17133
0 17135 5 1 1 17134
0 17136 7 1 2 62285 72638
0 17137 5 1 1 17136
0 17138 7 1 2 74621 17137
0 17139 5 1 1 17138
0 17140 7 1 2 64947 17139
0 17141 5 1 1 17140
0 17142 7 1 2 70972 72716
0 17143 5 1 1 17142
0 17144 7 1 2 72916 17143
0 17145 5 1 1 17144
0 17146 7 1 2 69238 17145
0 17147 5 1 1 17146
0 17148 7 1 2 72586 89175
0 17149 5 1 1 17148
0 17150 7 1 2 17147 17149
0 17151 5 1 1 17150
0 17152 7 1 2 62604 17151
0 17153 5 1 1 17152
0 17154 7 1 2 77176 17153
0 17155 5 1 1 17154
0 17156 7 1 2 71368 17155
0 17157 5 1 1 17156
0 17158 7 1 2 17141 17157
0 17159 5 1 1 17158
0 17160 7 1 2 61485 17159
0 17161 5 1 1 17160
0 17162 7 2 2 74201 72943
0 17163 5 2 1 90837
0 17164 7 1 2 79525 90839
0 17165 5 1 1 17164
0 17166 7 1 2 17161 17165
0 17167 5 1 1 17166
0 17168 7 1 2 66237 17167
0 17169 5 1 1 17168
0 17170 7 1 2 71548 90495
0 17171 5 1 1 17170
0 17172 7 2 2 70777 88810
0 17173 5 2 1 90841
0 17174 7 1 2 17171 90843
0 17175 5 1 1 17174
0 17176 7 1 2 82571 17175
0 17177 5 1 1 17176
0 17178 7 2 2 71549 72425
0 17179 5 1 1 90845
0 17180 7 1 2 76767 17179
0 17181 7 1 2 17177 17180
0 17182 5 2 1 17181
0 17183 7 1 2 61486 90847
0 17184 5 1 1 17183
0 17185 7 1 2 85584 17184
0 17186 5 1 1 17185
0 17187 7 1 2 71452 17186
0 17188 5 1 1 17187
0 17189 7 1 2 77831 84279
0 17190 5 1 1 17189
0 17191 7 2 2 7681 88447
0 17192 7 1 2 72547 78107
0 17193 5 1 1 17192
0 17194 7 1 2 60112 17193
0 17195 7 1 2 90849 17194
0 17196 5 1 1 17195
0 17197 7 1 2 65174 17196
0 17198 5 1 1 17197
0 17199 7 1 2 17190 17198
0 17200 5 1 1 17199
0 17201 7 1 2 64484 17200
0 17202 5 1 1 17201
0 17203 7 1 2 60113 70995
0 17204 5 1 1 17203
0 17205 7 1 2 64700 17204
0 17206 5 1 1 17205
0 17207 7 1 2 82732 71916
0 17208 5 1 1 17207
0 17209 7 2 2 73788 82773
0 17210 5 1 1 90851
0 17211 7 1 2 17210 88829
0 17212 7 1 2 17208 17211
0 17213 7 1 2 17206 17212
0 17214 5 1 1 17213
0 17215 7 1 2 65175 17214
0 17216 5 1 1 17215
0 17217 7 1 2 72671 88423
0 17218 5 1 1 17217
0 17219 7 1 2 65176 17218
0 17220 5 1 1 17219
0 17221 7 2 2 62605 77187
0 17222 7 1 2 78621 90853
0 17223 5 1 1 17222
0 17224 7 1 2 17220 17223
0 17225 5 1 1 17224
0 17226 7 1 2 69239 17225
0 17227 5 1 1 17226
0 17228 7 2 2 69792 77349
0 17229 7 5 2 64701 69064
0 17230 5 4 1 90857
0 17231 7 1 2 65998 90858
0 17232 7 1 2 90855 17231
0 17233 5 1 1 17232
0 17234 7 1 2 17227 17233
0 17235 7 1 2 17216 17234
0 17236 7 1 2 17202 17235
0 17237 5 1 1 17236
0 17238 7 1 2 61487 17237
0 17239 5 1 1 17238
0 17240 7 1 2 17188 17239
0 17241 7 1 2 17169 17240
0 17242 5 1 1 17241
0 17243 7 1 2 60482 17242
0 17244 5 1 1 17243
0 17245 7 1 2 73665 85479
0 17246 5 1 1 17245
0 17247 7 1 2 72944 88737
0 17248 5 1 1 17247
0 17249 7 1 2 17246 17248
0 17250 5 1 1 17249
0 17251 7 1 2 67574 17250
0 17252 5 1 1 17251
0 17253 7 1 2 63403 17252
0 17254 7 1 2 17244 17253
0 17255 5 1 1 17254
0 17256 7 1 2 72318 16961
0 17257 5 1 1 17256
0 17258 7 2 2 64702 71917
0 17259 5 2 1 90866
0 17260 7 4 2 73811 90868
0 17261 5 6 1 90870
0 17262 7 1 2 78347 90874
0 17263 5 1 1 17262
0 17264 7 2 2 76177 84077
0 17265 5 2 1 90880
0 17266 7 1 2 17263 90882
0 17267 5 1 1 17266
0 17268 7 1 2 71772 17267
0 17269 5 1 1 17268
0 17270 7 1 2 74507 89372
0 17271 5 1 1 17270
0 17272 7 1 2 78426 75996
0 17273 5 1 1 17272
0 17274 7 1 2 71102 17273
0 17275 5 1 1 17274
0 17276 7 1 2 17271 17275
0 17277 7 1 2 17269 17276
0 17278 7 1 2 17257 17277
0 17279 5 2 1 17278
0 17280 7 1 2 71550 90884
0 17281 5 1 1 17280
0 17282 7 1 2 73866 84579
0 17283 5 2 1 17282
0 17284 7 1 2 60311 90886
0 17285 5 1 1 17284
0 17286 7 1 2 62286 17285
0 17287 5 1 1 17286
0 17288 7 1 2 65177 71773
0 17289 5 2 1 17288
0 17290 7 1 2 78075 74611
0 17291 5 1 1 17290
0 17292 7 1 2 90888 17291
0 17293 7 1 2 17287 17292
0 17294 5 1 1 17293
0 17295 7 1 2 65708 17294
0 17296 5 1 1 17295
0 17297 7 1 2 74062 90343
0 17298 5 1 1 17297
0 17299 7 1 2 17296 17298
0 17300 5 1 1 17299
0 17301 7 1 2 64266 17300
0 17302 5 1 1 17301
0 17303 7 1 2 69240 82786
0 17304 5 1 1 17303
0 17305 7 2 2 73270 17304
0 17306 7 1 2 69144 72219
0 17307 7 1 2 90890 17306
0 17308 5 1 1 17307
0 17309 7 1 2 65178 17308
0 17310 5 1 1 17309
0 17311 7 3 2 62606 70922
0 17312 5 1 1 90892
0 17313 7 1 2 78998 90893
0 17314 5 1 1 17313
0 17315 7 1 2 79472 17314
0 17316 7 1 2 17310 17315
0 17317 7 1 2 17302 17316
0 17318 5 1 1 17317
0 17319 7 1 2 70778 17318
0 17320 5 1 1 17319
0 17321 7 1 2 17281 17320
0 17322 5 2 1 17321
0 17323 7 1 2 60483 90895
0 17324 5 1 1 17323
0 17325 7 1 2 71193 78320
0 17326 5 1 1 17325
0 17327 7 1 2 72917 89654
0 17328 5 1 1 17327
0 17329 7 1 2 17326 17328
0 17330 5 1 1 17329
0 17331 7 6 2 65375 67575
0 17332 5 2 1 90897
0 17333 7 1 2 60312 90898
0 17334 7 1 2 17330 17333
0 17335 5 1 1 17334
0 17336 7 1 2 17324 17335
0 17337 5 1 1 17336
0 17338 7 1 2 66448 17337
0 17339 5 1 1 17338
0 17340 7 2 2 62607 80562
0 17341 7 1 2 72717 88508
0 17342 5 1 1 17341
0 17343 7 1 2 71307 72889
0 17344 5 1 1 17343
0 17345 7 1 2 17342 17344
0 17346 5 1 1 17345
0 17347 7 1 2 62287 17346
0 17348 5 1 1 17347
0 17349 7 1 2 77171 17348
0 17350 5 1 1 17349
0 17351 7 1 2 90905 17350
0 17352 5 1 1 17351
0 17353 7 3 2 74063 71103
0 17354 5 3 1 90907
0 17355 7 1 2 89388 90910
0 17356 5 1 1 17355
0 17357 7 1 2 82009 17356
0 17358 5 1 1 17357
0 17359 7 1 2 75805 82699
0 17360 5 1 1 17359
0 17361 7 1 2 17358 17360
0 17362 5 1 1 17361
0 17363 7 1 2 88458 17362
0 17364 5 1 1 17363
0 17365 7 1 2 72185 88613
0 17366 5 1 1 17365
0 17367 7 1 2 88738 17366
0 17368 5 1 1 17367
0 17369 7 1 2 82010 72166
0 17370 7 1 2 90875 17369
0 17371 5 1 1 17370
0 17372 7 1 2 17368 17371
0 17373 7 1 2 17364 17372
0 17374 7 1 2 17352 17373
0 17375 5 1 1 17374
0 17376 7 1 2 66238 17375
0 17377 5 1 1 17376
0 17378 7 2 2 62608 88513
0 17379 5 1 1 90913
0 17380 7 1 2 82011 90914
0 17381 5 1 1 17380
0 17382 7 1 2 68313 17381
0 17383 7 1 2 17377 17382
0 17384 7 1 2 17339 17383
0 17385 5 1 1 17384
0 17386 7 1 2 63700 17385
0 17387 7 1 2 17255 17386
0 17388 5 1 1 17387
0 17389 7 1 2 61293 77203
0 17390 5 1 1 17389
0 17391 7 1 2 65999 17390
0 17392 5 1 1 17391
0 17393 7 2 2 66239 74064
0 17394 7 1 2 76977 90915
0 17395 5 1 1 17394
0 17396 7 1 2 17392 17395
0 17397 5 1 1 17396
0 17398 7 1 2 65709 17397
0 17399 5 1 1 17398
0 17400 7 1 2 17399 12482
0 17401 5 1 1 17400
0 17402 7 1 2 64267 17401
0 17403 5 1 1 17402
0 17404 7 2 2 61038 78458
0 17405 5 1 1 90917
0 17406 7 1 2 78358 17405
0 17407 5 2 1 17406
0 17408 7 1 2 71774 78405
0 17409 5 1 1 17408
0 17410 7 1 2 90919 17409
0 17411 5 1 1 17410
0 17412 7 1 2 66240 17411
0 17413 5 1 1 17412
0 17414 7 1 2 17403 17413
0 17415 5 1 1 17414
0 17416 7 1 2 62609 17415
0 17417 5 1 1 17416
0 17418 7 1 2 72167 88459
0 17419 5 1 1 17418
0 17420 7 2 2 75966 17419
0 17421 5 8 1 90921
0 17422 7 1 2 77704 90923
0 17423 5 1 1 17422
0 17424 7 1 2 17417 17423
0 17425 5 1 1 17424
0 17426 7 1 2 64703 17425
0 17427 5 1 1 17426
0 17428 7 1 2 81433 88290
0 17429 5 1 1 17428
0 17430 7 1 2 66000 17429
0 17431 5 1 1 17430
0 17432 7 1 2 89201 17431
0 17433 5 1 1 17432
0 17434 7 1 2 64485 17433
0 17435 5 1 1 17434
0 17436 7 1 2 89232 17435
0 17437 5 1 1 17436
0 17438 7 1 2 73164 17437
0 17439 5 1 1 17438
0 17440 7 1 2 17427 17439
0 17441 5 1 1 17440
0 17442 7 1 2 64948 17441
0 17443 5 1 1 17442
0 17444 7 1 2 80314 85422
0 17445 5 1 1 17444
0 17446 7 1 2 17443 17445
0 17447 5 1 1 17446
0 17448 7 1 2 60484 17447
0 17449 5 1 1 17448
0 17450 7 2 2 61294 80789
0 17451 7 1 2 80004 69305
0 17452 5 1 1 17451
0 17453 7 1 2 77122 69470
0 17454 5 3 1 17453
0 17455 7 1 2 76255 90933
0 17456 5 1 1 17455
0 17457 7 1 2 17452 17456
0 17458 5 1 1 17457
0 17459 7 1 2 90931 17458
0 17460 5 1 1 17459
0 17461 7 1 2 17449 17460
0 17462 5 1 1 17461
0 17463 7 5 2 75193 83525
0 17464 5 2 1 90936
0 17465 7 1 2 17462 90937
0 17466 5 1 1 17465
0 17467 7 1 2 66669 17466
0 17468 7 1 2 17388 17467
0 17469 7 1 2 17135 17468
0 17470 7 1 2 16503 17469
0 17471 5 1 1 17470
0 17472 7 1 2 62610 90226
0 17473 5 1 1 17472
0 17474 7 1 2 64268 90219
0 17475 5 1 1 17474
0 17476 7 1 2 17473 17475
0 17477 5 2 1 17476
0 17478 7 1 2 66001 90943
0 17479 5 1 1 17478
0 17480 7 1 2 74451 83828
0 17481 5 2 1 17480
0 17482 7 1 2 17479 90945
0 17483 5 1 1 17482
0 17484 7 1 2 62932 17483
0 17485 5 2 1 17484
0 17486 7 4 2 62080 72319
0 17487 5 3 1 90949
0 17488 7 2 2 69793 90950
0 17489 5 3 1 90956
0 17490 7 1 2 88927 90958
0 17491 5 1 1 17490
0 17492 7 1 2 62611 17491
0 17493 5 1 1 17492
0 17494 7 4 2 65710 62933
0 17495 5 3 1 90961
0 17496 7 1 2 79833 90962
0 17497 5 4 1 17496
0 17498 7 1 2 17493 90968
0 17499 5 1 1 17498
0 17500 7 1 2 69241 17499
0 17501 5 1 1 17500
0 17502 7 1 2 67949 78078
0 17503 5 3 1 17502
0 17504 7 1 2 60901 82380
0 17505 5 1 1 17504
0 17506 7 1 2 72320 17505
0 17507 7 1 2 90972 17506
0 17508 5 1 1 17507
0 17509 7 7 2 67950 76204
0 17510 5 4 1 90975
0 17511 7 1 2 71104 90982
0 17512 5 1 1 17511
0 17513 7 1 2 80296 90282
0 17514 5 2 1 17513
0 17515 7 1 2 82381 90986
0 17516 5 1 1 17515
0 17517 7 1 2 69154 17516
0 17518 5 1 1 17517
0 17519 7 1 2 17512 17518
0 17520 7 1 2 17508 17519
0 17521 7 1 2 17501 17520
0 17522 5 1 1 17521
0 17523 7 1 2 64949 17522
0 17524 5 1 1 17523
0 17525 7 1 2 90947 17524
0 17526 5 1 1 17525
0 17527 7 1 2 66449 17526
0 17528 5 1 1 17527
0 17529 7 1 2 75426 90541
0 17530 5 1 1 17529
0 17531 7 1 2 69794 17530
0 17532 5 1 1 17531
0 17533 7 1 2 84098 72220
0 17534 5 1 1 17533
0 17535 7 1 2 66450 17534
0 17536 5 1 1 17535
0 17537 7 1 2 17532 17536
0 17538 5 1 1 17537
0 17539 7 1 2 62934 17538
0 17540 5 1 1 17539
0 17541 7 1 2 62288 90560
0 17542 5 1 1 17541
0 17543 7 1 2 9928 17542
0 17544 5 1 1 17543
0 17545 7 1 2 69795 17544
0 17546 5 1 1 17545
0 17547 7 1 2 69155 88930
0 17548 5 1 1 17547
0 17549 7 1 2 69289 82850
0 17550 5 1 1 17549
0 17551 7 1 2 69796 82074
0 17552 5 1 1 17551
0 17553 7 1 2 17550 17552
0 17554 5 1 1 17553
0 17555 7 1 2 72321 17554
0 17556 5 1 1 17555
0 17557 7 1 2 17548 17556
0 17558 7 1 2 17546 17557
0 17559 5 1 1 17558
0 17560 7 1 2 66451 17559
0 17561 5 1 1 17560
0 17562 7 1 2 17540 17561
0 17563 5 1 1 17562
0 17564 7 2 2 64486 17563
0 17565 5 1 1 90988
0 17566 7 1 2 64950 90989
0 17567 5 1 1 17566
0 17568 7 1 2 17528 17567
0 17569 5 1 1 17568
0 17570 7 1 2 66241 17569
0 17571 5 1 1 17570
0 17572 7 1 2 66002 89895
0 17573 5 1 1 17572
0 17574 7 1 2 76636 77213
0 17575 5 1 1 17574
0 17576 7 1 2 17573 17575
0 17577 5 1 1 17576
0 17578 7 1 2 62935 17577
0 17579 5 1 1 17578
0 17580 7 1 2 84405 90946
0 17581 5 1 1 17580
0 17582 7 1 2 66003 17581
0 17583 5 1 1 17582
0 17584 7 1 2 74758 88037
0 17585 5 1 1 17584
0 17586 7 1 2 75981 71918
0 17587 5 1 1 17586
0 17588 7 1 2 17585 17587
0 17589 5 1 1 17588
0 17590 7 1 2 62936 17589
0 17591 5 1 1 17590
0 17592 7 1 2 17583 17591
0 17593 5 1 1 17592
0 17594 7 1 2 62081 17593
0 17595 5 1 1 17594
0 17596 7 1 2 17579 17595
0 17597 5 1 1 17596
0 17598 7 1 2 64704 17597
0 17599 5 1 1 17598
0 17600 7 1 2 90948 17599
0 17601 5 1 1 17600
0 17602 7 1 2 64951 17601
0 17603 5 1 1 17602
0 17604 7 3 2 62612 79585
0 17605 7 1 2 84078 90990
0 17606 5 1 1 17605
0 17607 7 1 2 85110 17606
0 17608 5 1 1 17607
0 17609 7 1 2 71974 17608
0 17610 5 1 1 17609
0 17611 7 3 2 62082 69982
0 17612 5 1 1 90993
0 17613 7 1 2 64487 90994
0 17614 5 1 1 17613
0 17615 7 1 2 64488 69156
0 17616 5 2 1 17615
0 17617 7 1 2 82473 90996
0 17618 7 1 2 90273 17617
0 17619 7 1 2 17614 17618
0 17620 5 1 1 17619
0 17621 7 1 2 78557 17620
0 17622 5 1 1 17621
0 17623 7 1 2 17610 17622
0 17624 5 1 1 17623
0 17625 7 1 2 66004 17624
0 17626 5 1 1 17625
0 17627 7 1 2 78558 90944
0 17628 5 1 1 17627
0 17629 7 1 2 17626 17628
0 17630 5 1 1 17629
0 17631 7 1 2 64705 17630
0 17632 5 1 1 17631
0 17633 7 1 2 17603 17632
0 17634 5 1 1 17633
0 17635 7 1 2 66452 17634
0 17636 5 1 1 17635
0 17637 7 1 2 17571 17636
0 17638 5 1 1 17637
0 17639 7 1 2 65179 17638
0 17640 5 1 1 17639
0 17641 7 1 2 79556 82139
0 17642 7 4 2 62937 77074
0 17643 5 1 1 90998
0 17644 7 3 2 71975 77291
0 17645 5 3 1 91002
0 17646 7 1 2 90999 91003
0 17647 7 1 2 17641 17646
0 17648 5 1 1 17647
0 17649 7 1 2 17640 17648
0 17650 5 1 1 17649
0 17651 7 1 2 84177 17650
0 17652 5 1 1 17651
0 17653 7 1 2 65376 89630
0 17654 5 1 1 17653
0 17655 7 1 2 83709 85458
0 17656 5 1 1 17655
0 17657 7 1 2 65180 11017
0 17658 7 1 2 17656 17657
0 17659 5 1 1 17658
0 17660 7 1 2 17654 17659
0 17661 5 1 1 17660
0 17662 7 1 2 72718 17661
0 17663 5 1 1 17662
0 17664 7 1 2 75876 88185
0 17665 5 1 1 17664
0 17666 7 1 2 4564 77842
0 17667 5 1 1 17666
0 17668 7 1 2 83710 85482
0 17669 5 8 1 17668
0 17670 7 1 2 82944 91008
0 17671 7 1 2 17667 17670
0 17672 5 1 1 17671
0 17673 7 1 2 17665 17672
0 17674 7 1 2 17663 17673
0 17675 5 1 1 17674
0 17676 7 1 2 63701 17675
0 17677 5 1 1 17676
0 17678 7 2 2 75194 78559
0 17679 5 1 1 91016
0 17680 7 1 2 84178 72890
0 17681 7 1 2 91017 17680
0 17682 5 1 1 17681
0 17683 7 1 2 17677 17682
0 17684 5 1 1 17683
0 17685 7 1 2 71369 17684
0 17686 5 1 1 17685
0 17687 7 1 2 72322 88389
0 17688 5 1 1 17687
0 17689 7 3 2 82572 75972
0 17690 5 1 1 91018
0 17691 7 1 2 61295 17690
0 17692 7 1 2 17688 17691
0 17693 5 1 1 17692
0 17694 7 1 2 62613 17693
0 17695 5 1 1 17694
0 17696 7 1 2 73934 90672
0 17697 7 1 2 17695 17696
0 17698 5 1 1 17697
0 17699 7 1 2 90666 17698
0 17700 5 1 1 17699
0 17701 7 1 2 90664 17700
0 17702 5 1 1 17701
0 17703 7 1 2 66453 17702
0 17704 5 1 1 17703
0 17705 7 1 2 90674 17704
0 17706 5 1 1 17705
0 17707 7 1 2 67951 17706
0 17708 5 1 1 17707
0 17709 7 1 2 70526 88291
0 17710 5 1 1 17709
0 17711 7 1 2 64489 17710
0 17712 5 1 1 17711
0 17713 7 1 2 82474 17712
0 17714 5 1 1 17713
0 17715 7 1 2 70779 17714
0 17716 5 1 1 17715
0 17717 7 1 2 71976 90881
0 17718 5 1 1 17717
0 17719 7 1 2 70149 17718
0 17720 7 1 2 17716 17719
0 17721 5 1 1 17720
0 17722 7 1 2 72323 17721
0 17723 5 1 1 17722
0 17724 7 1 2 82320 76538
0 17725 5 1 1 17724
0 17726 7 1 2 65844 17725
0 17727 5 1 1 17726
0 17728 7 1 2 78079 17727
0 17729 5 1 1 17728
0 17730 7 1 2 64490 17729
0 17731 5 1 1 17730
0 17732 7 1 2 70961 17731
0 17733 5 1 1 17732
0 17734 7 1 2 72491 17733
0 17735 5 1 1 17734
0 17736 7 1 2 83829 85983
0 17737 5 1 1 17736
0 17738 7 2 2 70780 90268
0 17739 5 1 1 91021
0 17740 7 1 2 72324 91022
0 17741 5 1 1 17740
0 17742 7 1 2 17737 17741
0 17743 5 1 1 17742
0 17744 7 1 2 74065 17743
0 17745 5 1 1 17744
0 17746 7 2 2 77737 88493
0 17747 5 1 1 91023
0 17748 7 3 2 61296 69900
0 17749 7 1 2 67046 91025
0 17750 5 1 1 17749
0 17751 7 1 2 65181 17750
0 17752 5 1 1 17751
0 17753 7 1 2 61488 17752
0 17754 7 1 2 17747 17753
0 17755 7 1 2 17745 17754
0 17756 7 1 2 17735 17755
0 17757 7 1 2 17723 17756
0 17758 5 1 1 17757
0 17759 7 1 2 81933 5656
0 17760 5 1 1 17759
0 17761 7 1 2 69177 17760
0 17762 5 1 1 17761
0 17763 7 1 2 80207 17762
0 17764 5 1 1 17763
0 17765 7 1 2 67576 17764
0 17766 5 1 1 17765
0 17767 7 1 2 74829 84066
0 17768 5 1 1 17767
0 17769 7 1 2 73638 17768
0 17770 5 1 1 17769
0 17771 7 1 2 88722 17770
0 17772 5 1 1 17771
0 17773 7 1 2 17766 17772
0 17774 5 1 1 17773
0 17775 7 1 2 71194 17774
0 17776 5 1 1 17775
0 17777 7 1 2 76132 76607
0 17778 7 1 2 82549 17777
0 17779 7 1 2 90488 17778
0 17780 5 1 1 17779
0 17781 7 1 2 72918 17780
0 17782 5 1 1 17781
0 17783 7 1 2 67577 88556
0 17784 5 1 1 17783
0 17785 7 3 2 62614 72097
0 17786 5 1 1 91028
0 17787 7 1 2 69531 91029
0 17788 5 2 1 17787
0 17789 7 1 2 67277 91031
0 17790 7 1 2 17784 17789
0 17791 5 1 1 17790
0 17792 7 2 2 61297 77334
0 17793 5 2 1 91033
0 17794 7 1 2 76671 91034
0 17795 7 1 2 17791 17794
0 17796 5 1 1 17795
0 17797 7 1 2 72919 74445
0 17798 5 1 1 17797
0 17799 7 1 2 66242 17798
0 17800 5 1 1 17799
0 17801 7 1 2 90483 17800
0 17802 5 1 1 17801
0 17803 7 1 2 66454 17802
0 17804 7 1 2 17796 17803
0 17805 7 1 2 17782 17804
0 17806 7 1 2 17776 17805
0 17807 5 1 1 17806
0 17808 7 1 2 62938 17807
0 17809 7 1 2 17758 17808
0 17810 5 1 1 17809
0 17811 7 3 2 62289 90496
0 17812 5 1 1 91037
0 17813 7 1 2 69797 91038
0 17814 5 1 1 17813
0 17815 7 1 2 90871 17814
0 17816 5 1 1 17815
0 17817 7 1 2 71551 17816
0 17818 5 1 1 17817
0 17819 7 3 2 70781 84079
0 17820 5 1 1 91040
0 17821 7 1 2 88811 91041
0 17822 5 1 1 17821
0 17823 7 1 2 71035 17822
0 17824 7 1 2 17818 17823
0 17825 5 1 1 17824
0 17826 7 1 2 71775 17825
0 17827 5 1 1 17826
0 17828 7 1 2 71036 79117
0 17829 5 1 1 17828
0 17830 7 1 2 72325 17829
0 17831 5 1 1 17830
0 17832 7 1 2 71105 90336
0 17833 5 2 1 17832
0 17834 7 3 2 71552 72326
0 17835 5 2 1 91045
0 17836 7 1 2 79227 91048
0 17837 7 1 2 91043 17836
0 17838 5 1 1 17837
0 17839 7 1 2 84072 17838
0 17840 5 1 1 17839
0 17841 7 1 2 17831 17840
0 17842 7 1 2 17827 17841
0 17843 5 1 1 17842
0 17844 7 1 2 61489 17843
0 17845 5 1 1 17844
0 17846 7 1 2 73666 84032
0 17847 5 1 1 17846
0 17848 7 1 2 75139 82945
0 17849 5 1 1 17848
0 17850 7 1 2 85585 17849
0 17851 5 1 1 17850
0 17852 7 1 2 90840 17851
0 17853 5 1 1 17852
0 17854 7 1 2 17847 17853
0 17855 7 1 2 17845 17854
0 17856 7 1 2 17810 17855
0 17857 7 1 2 17708 17856
0 17858 5 1 1 17857
0 17859 7 1 2 65377 17858
0 17860 5 1 1 17859
0 17861 7 6 2 60485 65845
0 17862 7 1 2 76637 91050
0 17863 7 1 2 84963 17862
0 17864 5 1 1 17863
0 17865 7 3 2 61490 76638
0 17866 5 1 1 91056
0 17867 7 1 2 86290 91057
0 17868 5 1 1 17867
0 17869 7 1 2 85459 17868
0 17870 5 1 1 17869
0 17871 7 1 2 70598 83817
0 17872 5 2 1 17871
0 17873 7 1 2 65182 91059
0 17874 7 1 2 17870 17873
0 17875 5 1 1 17874
0 17876 7 1 2 17864 17875
0 17877 5 1 1 17876
0 17878 7 1 2 64491 17877
0 17879 5 1 1 17878
0 17880 7 4 2 80563 74319
0 17881 5 1 1 91061
0 17882 7 1 2 69242 91062
0 17883 5 1 1 17882
0 17884 7 1 2 17879 17883
0 17885 5 1 1 17884
0 17886 7 1 2 69798 17885
0 17887 5 1 1 17886
0 17888 7 1 2 84977 91063
0 17889 5 1 1 17888
0 17890 7 1 2 17887 17889
0 17891 5 1 1 17890
0 17892 7 1 2 62083 17891
0 17893 5 1 1 17892
0 17894 7 1 2 86633 89795
0 17895 5 1 1 17894
0 17896 7 2 2 70150 75967
0 17897 7 1 2 17895 91065
0 17898 5 1 1 17897
0 17899 7 1 2 91064 17898
0 17900 5 1 1 17899
0 17901 7 1 2 17893 17900
0 17902 5 1 1 17901
0 17903 7 1 2 62939 17902
0 17904 5 1 1 17903
0 17905 7 1 2 60486 89896
0 17906 5 1 1 17905
0 17907 7 1 2 60487 83138
0 17908 5 1 1 17907
0 17909 7 9 2 67278 78250
0 17910 5 2 1 91067
0 17911 7 1 2 88323 91068
0 17912 5 3 1 17911
0 17913 7 1 2 17908 91078
0 17914 5 1 1 17913
0 17915 7 1 2 69799 17914
0 17916 5 1 1 17915
0 17917 7 1 2 17906 17916
0 17918 5 1 1 17917
0 17919 7 1 2 87575 17918
0 17920 5 1 1 17919
0 17921 7 1 2 17904 17920
0 17922 5 1 1 17921
0 17923 7 1 2 72327 17922
0 17924 5 1 1 17923
0 17925 7 1 2 69800 89897
0 17926 5 1 1 17925
0 17927 7 1 2 90022 17926
0 17928 5 1 1 17927
0 17929 7 1 2 62084 17928
0 17930 5 1 1 17929
0 17931 7 3 2 73096 70947
0 17932 5 2 1 91081
0 17933 7 1 2 17930 91084
0 17934 5 1 1 17933
0 17935 7 4 2 87236 87827
0 17936 5 1 1 91086
0 17937 7 1 2 71106 91087
0 17938 5 1 1 17937
0 17939 7 1 2 17881 17938
0 17940 5 1 1 17939
0 17941 7 1 2 17934 17940
0 17942 5 1 1 17941
0 17943 7 1 2 85643 91024
0 17944 5 1 1 17943
0 17945 7 1 2 17942 17944
0 17946 5 1 1 17945
0 17947 7 1 2 62940 17946
0 17948 5 1 1 17947
0 17949 7 1 2 85414 91019
0 17950 5 1 1 17949
0 17951 7 1 2 74566 81323
0 17952 5 1 1 17951
0 17953 7 1 2 17950 17952
0 17954 5 1 1 17953
0 17955 7 1 2 60488 17954
0 17956 5 1 1 17955
0 17957 7 4 2 69801 77159
0 17958 7 1 2 76386 86874
0 17959 7 1 2 91090 17958
0 17960 5 1 1 17959
0 17961 7 1 2 17956 17960
0 17962 5 1 1 17961
0 17963 7 1 2 75195 17962
0 17964 5 1 1 17963
0 17965 7 1 2 17948 17964
0 17966 7 1 2 17924 17965
0 17967 7 1 2 17860 17966
0 17968 5 1 1 17967
0 17969 7 1 2 63702 17968
0 17970 5 1 1 17969
0 17971 7 1 2 17686 17970
0 17972 7 1 2 17652 17971
0 17973 5 1 1 17972
0 17974 7 1 2 63404 17973
0 17975 5 1 1 17974
0 17976 7 1 2 70782 89122
0 17977 5 1 1 17976
0 17978 7 1 2 62290 78538
0 17979 5 1 1 17978
0 17980 7 1 2 17977 17979
0 17981 5 1 1 17980
0 17982 7 1 2 66455 17981
0 17983 5 1 1 17982
0 17984 7 2 2 66243 70484
0 17985 7 1 2 77832 91094
0 17986 5 1 1 17985
0 17987 7 1 2 17983 17986
0 17988 5 1 1 17987
0 17989 7 1 2 65183 17988
0 17990 5 1 1 17989
0 17991 7 1 2 85271 88317
0 17992 5 1 1 17991
0 17993 7 1 2 17990 17992
0 17994 5 1 1 17993
0 17995 7 1 2 71977 17994
0 17996 5 1 1 17995
0 17997 7 2 2 80448 82632
0 17998 5 1 1 91096
0 17999 7 1 2 90761 17998
0 18000 5 1 1 17999
0 18001 7 1 2 17996 18000
0 18002 5 1 1 18001
0 18003 7 1 2 62941 18002
0 18004 5 1 1 18003
0 18005 7 6 2 64952 78032
0 18006 5 1 1 91098
0 18007 7 1 2 75196 91099
0 18008 7 1 2 72632 18007
0 18009 5 1 1 18008
0 18010 7 1 2 18004 18009
0 18011 5 1 1 18010
0 18012 7 1 2 62615 18011
0 18013 5 1 1 18012
0 18014 7 2 2 64953 79586
0 18015 5 1 1 91104
0 18016 7 1 2 78591 90379
0 18017 5 1 1 18016
0 18018 7 1 2 91105 18017
0 18019 5 1 1 18018
0 18020 7 1 2 78698 86376
0 18021 5 1 1 18020
0 18022 7 1 2 18019 18021
0 18023 5 1 1 18022
0 18024 7 1 2 79544 18023
0 18025 5 1 1 18024
0 18026 7 1 2 18013 18025
0 18027 5 1 1 18026
0 18028 7 1 2 84213 18027
0 18029 5 1 1 18028
0 18030 7 1 2 90842 91009
0 18031 5 1 1 18030
0 18032 7 2 2 66456 82946
0 18033 5 5 1 91106
0 18034 7 3 2 75550 91108
0 18035 7 2 2 65378 91113
0 18036 5 1 1 91116
0 18037 7 1 2 70047 91010
0 18038 5 1 1 18037
0 18039 7 1 2 18036 18038
0 18040 5 1 1 18039
0 18041 7 1 2 90497 18040
0 18042 5 1 1 18041
0 18043 7 1 2 18031 18042
0 18044 5 1 1 18043
0 18045 7 1 2 62085 18044
0 18046 5 1 1 18045
0 18047 7 1 2 72492 91011
0 18048 5 1 1 18047
0 18049 7 2 2 83458 71271
0 18050 5 1 1 91118
0 18051 7 1 2 87828 91119
0 18052 5 1 1 18051
0 18053 7 1 2 18048 18052
0 18054 5 1 1 18053
0 18055 7 1 2 77466 18054
0 18056 5 1 1 18055
0 18057 7 1 2 18046 18056
0 18058 5 1 1 18057
0 18059 7 1 2 87970 18058
0 18060 5 1 1 18059
0 18061 7 11 2 62942 70783
0 18062 5 6 1 91120
0 18063 7 3 2 70151 72427
0 18064 5 1 1 91137
0 18065 7 1 2 91121 18064
0 18066 5 1 1 18065
0 18067 7 1 2 9234 18066
0 18068 5 1 1 18067
0 18069 7 1 2 75551 18068
0 18070 5 1 1 18069
0 18071 7 1 2 75197 85988
0 18072 5 1 1 18071
0 18073 7 1 2 18070 18072
0 18074 5 1 1 18073
0 18075 7 1 2 82168 18074
0 18076 5 1 1 18075
0 18077 7 1 2 18060 18076
0 18078 5 1 1 18077
0 18079 7 1 2 63703 18078
0 18080 5 1 1 18079
0 18081 7 2 2 83526 87822
0 18082 7 1 2 79400 91140
0 18083 7 1 2 79601 18082
0 18084 5 1 1 18083
0 18085 7 1 2 18080 18084
0 18086 5 1 1 18085
0 18087 7 1 2 69243 18086
0 18088 5 1 1 18087
0 18089 7 1 2 67578 73977
0 18090 5 4 1 18089
0 18091 7 1 2 79807 87676
0 18092 5 2 1 18091
0 18093 7 1 2 71553 91146
0 18094 5 1 1 18093
0 18095 7 4 2 66457 77897
0 18096 7 1 2 61298 91148
0 18097 5 1 1 18096
0 18098 7 1 2 77616 79401
0 18099 5 1 1 18098
0 18100 7 1 2 18097 18099
0 18101 7 1 2 18094 18100
0 18102 5 1 1 18101
0 18103 7 1 2 62086 18102
0 18104 5 1 1 18103
0 18105 7 3 2 80585 86828
0 18106 5 1 1 91152
0 18107 7 1 2 68314 91153
0 18108 5 1 1 18107
0 18109 7 1 2 18104 18108
0 18110 5 1 1 18109
0 18111 7 1 2 65379 18110
0 18112 5 1 1 18111
0 18113 7 1 2 80024 76842
0 18114 7 1 2 82012 18113
0 18115 5 1 1 18114
0 18116 7 1 2 18112 18115
0 18117 5 1 1 18116
0 18118 7 1 2 84667 18117
0 18119 5 1 1 18118
0 18120 7 11 2 68643 83094
0 18121 7 2 2 87526 91155
0 18122 5 1 1 91166
0 18123 7 1 2 81269 91167
0 18124 5 1 1 18123
0 18125 7 1 2 18119 18124
0 18126 5 1 1 18125
0 18127 7 1 2 91142 18126
0 18128 5 1 1 18127
0 18129 7 3 2 62943 74881
0 18130 5 4 1 91168
0 18131 7 1 2 75427 91171
0 18132 5 1 1 18131
0 18133 7 1 2 73097 18132
0 18134 5 1 1 18133
0 18135 7 1 2 62616 75416
0 18136 5 1 1 18135
0 18137 7 1 2 18134 18136
0 18138 5 1 1 18137
0 18139 7 1 2 66005 18138
0 18140 5 1 1 18139
0 18141 7 1 2 82675 74928
0 18142 5 1 1 18141
0 18143 7 1 2 18140 18142
0 18144 5 1 1 18143
0 18145 7 1 2 65846 18144
0 18146 5 1 1 18145
0 18147 7 1 2 67952 90296
0 18148 5 5 1 18147
0 18149 7 1 2 84855 91175
0 18150 5 1 1 18149
0 18151 7 1 2 18146 18150
0 18152 5 1 1 18151
0 18153 7 1 2 82169 18152
0 18154 5 1 1 18153
0 18155 7 5 2 63405 77467
0 18156 5 1 1 91180
0 18157 7 1 2 86398 90311
0 18158 7 1 2 91181 18157
0 18159 5 1 1 18158
0 18160 7 1 2 18154 18159
0 18161 5 1 1 18160
0 18162 7 1 2 71554 18161
0 18163 5 1 1 18162
0 18164 7 2 2 62944 71776
0 18165 5 2 1 91185
0 18166 7 2 2 59845 70929
0 18167 5 1 1 91189
0 18168 7 1 2 91186 18167
0 18169 5 1 1 18168
0 18170 7 1 2 90548 18169
0 18171 5 1 1 18170
0 18172 7 1 2 62291 18171
0 18173 5 1 1 18172
0 18174 7 1 2 91172 18173
0 18175 5 1 1 18174
0 18176 7 1 2 91012 18175
0 18177 5 1 1 18176
0 18178 7 6 2 65380 62087
0 18179 7 1 2 75140 91191
0 18180 5 1 1 18179
0 18181 7 1 2 18177 18180
0 18182 5 1 1 18181
0 18183 7 1 2 63406 18182
0 18184 5 1 1 18183
0 18185 7 1 2 86928 87443
0 18186 5 1 1 18185
0 18187 7 1 2 18184 18186
0 18188 5 1 1 18187
0 18189 7 1 2 70784 18188
0 18190 5 1 1 18189
0 18191 7 3 2 62292 71919
0 18192 5 3 1 91197
0 18193 7 1 2 65847 91198
0 18194 5 2 1 18193
0 18195 7 1 2 73812 91203
0 18196 5 4 1 18195
0 18197 7 1 2 79597 91013
0 18198 5 1 1 18197
0 18199 7 1 2 62088 91117
0 18200 5 1 1 18199
0 18201 7 1 2 18198 18200
0 18202 5 1 1 18201
0 18203 7 1 2 63407 18202
0 18204 5 1 1 18203
0 18205 7 1 2 82170 91154
0 18206 5 1 1 18205
0 18207 7 1 2 18204 18206
0 18208 5 1 1 18207
0 18209 7 1 2 91205 18208
0 18210 5 1 1 18209
0 18211 7 1 2 60489 79473
0 18212 5 7 1 18211
0 18213 7 3 2 62945 91209
0 18214 5 1 1 91216
0 18215 7 1 2 74882 91147
0 18216 7 1 2 91217 18215
0 18217 5 1 1 18216
0 18218 7 1 2 74222 80508
0 18219 7 1 2 88546 18218
0 18220 5 1 1 18219
0 18221 7 1 2 18217 18220
0 18222 5 1 1 18221
0 18223 7 1 2 77292 18222
0 18224 5 1 1 18223
0 18225 7 1 2 83266 87841
0 18226 5 1 1 18225
0 18227 7 1 2 18224 18226
0 18228 5 1 1 18227
0 18229 7 1 2 72623 18228
0 18230 5 1 1 18229
0 18231 7 1 2 75740 91149
0 18232 5 1 1 18231
0 18233 7 1 2 77604 79402
0 18234 7 1 2 91176 18233
0 18235 5 1 1 18234
0 18236 7 1 2 18232 18235
0 18237 5 1 1 18236
0 18238 7 1 2 64954 18237
0 18239 5 1 1 18238
0 18240 7 1 2 71006 85583
0 18241 5 1 1 18240
0 18242 7 1 2 18239 18241
0 18243 5 1 1 18242
0 18244 7 1 2 65381 18243
0 18245 5 1 1 18244
0 18246 7 1 2 18230 18245
0 18247 7 1 2 18210 18246
0 18248 7 1 2 18190 18247
0 18249 7 1 2 18163 18248
0 18250 5 1 1 18249
0 18251 7 1 2 63704 18250
0 18252 5 1 1 18251
0 18253 7 1 2 18128 18252
0 18254 7 1 2 18088 18253
0 18255 7 1 2 18029 18254
0 18256 5 1 1 18255
0 18257 7 1 2 69654 18256
0 18258 5 1 1 18257
0 18259 7 3 2 75552 71107
0 18260 5 2 1 91219
0 18261 7 2 2 86841 91222
0 18262 5 1 1 91224
0 18263 7 1 2 70152 91225
0 18264 5 1 1 18263
0 18265 7 1 2 83476 84659
0 18266 5 1 1 18265
0 18267 7 1 2 18264 18266
0 18268 5 1 1 18267
0 18269 7 1 2 75275 18268
0 18270 5 1 1 18269
0 18271 7 1 2 62617 18270
0 18272 5 1 1 18271
0 18273 7 1 2 83482 78929
0 18274 5 1 1 18273
0 18275 7 1 2 18272 18274
0 18276 5 1 1 18275
0 18277 7 1 2 69065 18276
0 18278 5 1 1 18277
0 18279 7 4 2 70785 73856
0 18280 5 1 1 91226
0 18281 7 1 2 75276 18280
0 18282 5 1 1 18281
0 18283 7 1 2 86829 18282
0 18284 5 1 1 18283
0 18285 7 1 2 18278 18284
0 18286 5 1 1 18285
0 18287 7 1 2 72587 18286
0 18288 5 1 1 18287
0 18289 7 3 2 75553 83792
0 18290 7 1 2 77738 91230
0 18291 5 1 1 18290
0 18292 7 2 2 87232 91046
0 18293 5 2 1 91233
0 18294 7 1 2 77235 86647
0 18295 5 1 1 18294
0 18296 7 1 2 91235 18295
0 18297 7 1 2 18291 18296
0 18298 5 1 1 18297
0 18299 7 1 2 76639 18298
0 18300 5 1 1 18299
0 18301 7 1 2 18288 18300
0 18302 5 1 1 18301
0 18303 7 1 2 62089 18302
0 18304 5 1 1 18303
0 18305 7 1 2 72420 91234
0 18306 5 1 1 18305
0 18307 7 1 2 90764 18306
0 18308 5 1 1 18307
0 18309 7 1 2 72588 18308
0 18310 5 1 1 18309
0 18311 7 1 2 90510 89508
0 18312 5 1 1 18311
0 18313 7 1 2 75554 18312
0 18314 5 1 1 18313
0 18315 7 3 2 70599 73813
0 18316 5 3 1 91237
0 18317 7 1 2 64706 91240
0 18318 5 1 1 18317
0 18319 7 4 2 76144 88830
0 18320 5 1 1 91243
0 18321 7 1 2 18318 91244
0 18322 5 1 1 18321
0 18323 7 1 2 75555 18322
0 18324 5 1 1 18323
0 18325 7 1 2 77848 18324
0 18326 5 1 1 18325
0 18327 7 1 2 73376 18326
0 18328 5 1 1 18327
0 18329 7 1 2 18314 18328
0 18330 5 1 1 18329
0 18331 7 1 2 62946 75037
0 18332 7 1 2 18330 18331
0 18333 5 1 1 18332
0 18334 7 1 2 18310 18333
0 18335 5 1 1 18334
0 18336 7 1 2 69244 18335
0 18337 5 1 1 18336
0 18338 7 2 2 70973 73789
0 18339 5 1 1 91247
0 18340 7 1 2 88946 18339
0 18341 5 1 1 18340
0 18342 7 1 2 69066 18341
0 18343 5 1 1 18342
0 18344 7 3 2 62947 73790
0 18345 5 2 1 91249
0 18346 7 1 2 18343 91252
0 18347 5 1 1 18346
0 18348 7 1 2 64707 18347
0 18349 5 1 1 18348
0 18350 7 1 2 83813 78930
0 18351 5 1 1 18350
0 18352 7 1 2 18349 18351
0 18353 5 1 1 18352
0 18354 7 1 2 70786 18353
0 18355 5 1 1 18354
0 18356 7 1 2 78638 91206
0 18357 5 1 1 18356
0 18358 7 1 2 83872 78093
0 18359 7 1 2 18357 18358
0 18360 5 1 1 18359
0 18361 7 1 2 70048 18360
0 18362 5 1 1 18361
0 18363 7 1 2 18355 18362
0 18364 5 1 1 18363
0 18365 7 1 2 75556 18364
0 18366 5 1 1 18365
0 18367 7 1 2 82382 86915
0 18368 5 2 1 18367
0 18369 7 2 2 69802 91254
0 18370 5 1 1 91256
0 18371 7 1 2 60114 85111
0 18372 5 1 1 18371
0 18373 7 1 2 91257 18372
0 18374 5 1 1 18373
0 18375 7 1 2 85659 86513
0 18376 5 1 1 18375
0 18377 7 1 2 18374 18376
0 18378 5 1 1 18377
0 18379 7 1 2 64708 18378
0 18380 5 1 1 18379
0 18381 7 1 2 86550 18380
0 18382 5 1 1 18381
0 18383 7 1 2 75557 18382
0 18384 5 1 1 18383
0 18385 7 1 2 77261 89517
0 18386 5 1 1 18385
0 18387 7 1 2 75198 18386
0 18388 5 1 1 18387
0 18389 7 1 2 18384 18388
0 18390 5 1 1 18389
0 18391 7 1 2 91143 18390
0 18392 5 1 1 18391
0 18393 7 1 2 70231 70983
0 18394 5 1 1 18393
0 18395 7 1 2 91204 91238
0 18396 5 1 1 18395
0 18397 7 1 2 18394 18396
0 18398 5 1 1 18397
0 18399 7 1 2 62948 82592
0 18400 5 1 1 18399
0 18401 7 1 2 78094 18400
0 18402 7 1 2 18398 18401
0 18403 5 1 1 18402
0 18404 7 1 2 75199 18403
0 18405 5 1 1 18404
0 18406 7 1 2 18392 18405
0 18407 7 1 2 18366 18406
0 18408 7 1 2 18337 18407
0 18409 7 1 2 18304 18408
0 18410 5 1 1 18409
0 18411 7 1 2 65382 18410
0 18412 5 1 1 18411
0 18413 7 1 2 76178 82820
0 18414 7 1 2 75973 84403
0 18415 7 1 2 18413 18414
0 18416 5 1 1 18415
0 18417 7 1 2 18412 18416
0 18418 5 1 1 18417
0 18419 7 1 2 78748 18418
0 18420 5 1 1 18419
0 18421 7 1 2 61688 18420
0 18422 7 1 2 18258 18421
0 18423 7 1 2 17975 18422
0 18424 5 1 1 18423
0 18425 7 1 2 17471 18424
0 18426 5 1 1 18425
0 18427 7 1 2 68855 18426
0 18428 5 1 1 18427
0 18429 7 1 2 74414 82283
0 18430 5 1 1 18429
0 18431 7 1 2 82141 18430
0 18432 5 1 1 18431
0 18433 7 1 2 70049 18432
0 18434 5 1 1 18433
0 18435 7 4 2 69655 72328
0 18436 5 2 1 91258
0 18437 7 1 2 62618 91259
0 18438 5 1 1 18437
0 18439 7 1 2 90987 18438
0 18440 5 1 1 18439
0 18441 7 1 2 65848 18440
0 18442 5 1 1 18441
0 18443 7 1 2 88817 18442
0 18444 5 1 1 18443
0 18445 7 1 2 64492 18444
0 18446 5 1 1 18445
0 18447 7 1 2 72877 81688
0 18448 5 1 1 18447
0 18449 7 1 2 18446 18448
0 18450 5 1 1 18449
0 18451 7 1 2 62949 18450
0 18452 5 1 1 18451
0 18453 7 1 2 18434 18452
0 18454 5 1 1 18453
0 18455 7 1 2 62293 18454
0 18456 5 1 1 18455
0 18457 7 2 2 65849 73310
0 18458 5 1 1 91264
0 18459 7 2 2 64709 76241
0 18460 5 1 1 91266
0 18461 7 1 2 18458 18460
0 18462 5 1 1 18461
0 18463 7 1 2 77468 18462
0 18464 5 1 1 18463
0 18465 7 2 2 77075 76843
0 18466 5 1 1 91268
0 18467 7 1 2 18464 18466
0 18468 5 1 1 18467
0 18469 7 1 2 66006 18468
0 18470 5 1 1 18469
0 18471 7 1 2 62294 90963
0 18472 5 1 1 18471
0 18473 7 1 2 5596 18472
0 18474 5 1 1 18473
0 18475 7 1 2 64710 18474
0 18476 5 1 1 18475
0 18477 7 3 2 60902 82649
0 18478 5 2 1 91270
0 18479 7 1 2 72437 91273
0 18480 5 1 1 18479
0 18481 7 1 2 67579 18480
0 18482 5 1 1 18481
0 18483 7 1 2 59498 90236
0 18484 5 1 1 18483
0 18485 7 1 2 62950 18484
0 18486 7 1 2 18482 18485
0 18487 5 1 1 18486
0 18488 7 1 2 18476 18487
0 18489 5 1 1 18488
0 18490 7 1 2 64269 18489
0 18491 5 1 1 18490
0 18492 7 1 2 71777 82133
0 18493 5 1 1 18492
0 18494 7 1 2 67580 76469
0 18495 5 1 1 18494
0 18496 7 1 2 62295 82200
0 18497 7 1 2 18495 18496
0 18498 5 1 1 18497
0 18499 7 1 2 18493 18498
0 18500 5 1 1 18499
0 18501 7 1 2 62951 18500
0 18502 5 1 1 18501
0 18503 7 2 2 65711 90546
0 18504 5 2 1 91275
0 18505 7 1 2 64711 90246
0 18506 5 1 1 18505
0 18507 7 1 2 85820 18506
0 18508 5 1 1 18507
0 18509 7 1 2 82799 72329
0 18510 7 1 2 18508 18509
0 18511 5 1 1 18510
0 18512 7 1 2 91277 18511
0 18513 7 1 2 18502 18512
0 18514 7 1 2 18491 18513
0 18515 5 1 1 18514
0 18516 7 1 2 70787 18515
0 18517 5 1 1 18516
0 18518 7 1 2 18470 18517
0 18519 7 1 2 18456 18518
0 18520 5 1 1 18519
0 18521 7 1 2 75558 18520
0 18522 5 1 1 18521
0 18523 7 3 2 62952 72493
0 18524 5 2 1 91279
0 18525 7 2 2 90536 91282
0 18526 7 1 2 70788 90551
0 18527 5 1 1 18526
0 18528 7 1 2 91284 18527
0 18529 5 1 1 18528
0 18530 7 1 2 64493 18529
0 18531 5 1 1 18530
0 18532 7 4 2 64494 71108
0 18533 5 2 1 91286
0 18534 7 1 2 90965 91290
0 18535 5 1 1 18534
0 18536 7 1 2 70789 18535
0 18537 5 1 1 18536
0 18538 7 1 2 65712 79065
0 18539 5 1 1 18538
0 18540 7 1 2 3783 18539
0 18541 7 1 2 18537 18540
0 18542 5 1 1 18541
0 18543 7 1 2 64270 18542
0 18544 5 1 1 18543
0 18545 7 1 2 18531 18544
0 18546 5 1 1 18545
0 18547 7 1 2 75559 18546
0 18548 5 1 1 18547
0 18549 7 1 2 80297 77855
0 18550 7 1 2 78560 18549
0 18551 5 1 1 18550
0 18552 7 1 2 88281 18551
0 18553 5 1 1 18552
0 18554 7 1 2 64271 18553
0 18555 5 1 1 18554
0 18556 7 3 2 66458 77528
0 18557 5 1 1 91292
0 18558 7 1 2 86014 18557
0 18559 5 1 1 18558
0 18560 7 1 2 64495 18559
0 18561 5 1 1 18560
0 18562 7 1 2 18555 18561
0 18563 7 1 2 18548 18562
0 18564 5 1 1 18563
0 18565 7 1 2 62090 18564
0 18566 5 1 1 18565
0 18567 7 4 2 66459 71555
0 18568 5 3 1 91295
0 18569 7 1 2 78644 91296
0 18570 5 1 1 18569
0 18571 7 2 2 66244 72330
0 18572 5 4 1 91302
0 18573 7 1 2 71029 91303
0 18574 5 1 1 18573
0 18575 7 1 2 77257 78990
0 18576 5 1 1 18575
0 18577 7 5 2 75560 72331
0 18578 5 1 1 91308
0 18579 7 1 2 62953 91309
0 18580 5 1 1 18579
0 18581 7 1 2 18576 18580
0 18582 5 1 1 18581
0 18583 7 1 2 70790 18582
0 18584 5 1 1 18583
0 18585 7 1 2 18574 18584
0 18586 7 1 2 18570 18585
0 18587 7 1 2 18566 18586
0 18588 5 1 1 18587
0 18589 7 1 2 69157 18588
0 18590 5 1 1 18589
0 18591 7 2 2 61491 77519
0 18592 5 2 1 91313
0 18593 7 1 2 91260 91315
0 18594 5 1 1 18593
0 18595 7 1 2 84080 79066
0 18596 5 1 1 18595
0 18597 7 1 2 18594 18596
0 18598 5 1 1 18597
0 18599 7 1 2 65850 18598
0 18600 5 1 1 18599
0 18601 7 1 2 62954 74129
0 18602 5 1 1 18601
0 18603 7 1 2 61492 18602
0 18604 5 1 1 18603
0 18605 7 1 2 71109 18604
0 18606 5 1 1 18605
0 18607 7 1 2 18600 18606
0 18608 5 1 1 18607
0 18609 7 1 2 66245 18608
0 18610 5 1 1 18609
0 18611 7 3 2 66007 74929
0 18612 7 1 2 76702 91317
0 18613 5 1 1 18612
0 18614 7 1 2 61493 78045
0 18615 5 1 1 18614
0 18616 7 1 2 65184 18615
0 18617 5 1 1 18616
0 18618 7 1 2 18613 18617
0 18619 7 1 2 18610 18618
0 18620 5 1 1 18619
0 18621 7 1 2 64496 18620
0 18622 5 1 1 18621
0 18623 7 7 2 64272 66460
0 18624 5 2 1 91320
0 18625 7 3 2 82134 91321
0 18626 5 1 1 91329
0 18627 7 1 2 10638 18626
0 18628 5 1 1 18627
0 18629 7 1 2 65851 18628
0 18630 5 1 1 18629
0 18631 7 3 2 66246 69656
0 18632 5 2 1 91332
0 18633 7 1 2 66461 91333
0 18634 5 1 1 18633
0 18635 7 1 2 18630 18634
0 18636 5 1 1 18635
0 18637 7 1 2 66008 18636
0 18638 5 1 1 18637
0 18639 7 1 2 60313 12461
0 18640 5 1 1 18639
0 18641 7 1 2 66462 18640
0 18642 5 1 1 18641
0 18643 7 1 2 18638 18642
0 18644 5 1 1 18643
0 18645 7 1 2 64712 18644
0 18646 5 1 1 18645
0 18647 7 1 2 60314 77717
0 18648 5 1 1 18647
0 18649 7 1 2 66463 18648
0 18650 5 1 1 18649
0 18651 7 1 2 62619 79067
0 18652 7 1 2 90230 18651
0 18653 5 1 1 18652
0 18654 7 1 2 18650 18653
0 18655 5 1 1 18654
0 18656 7 1 2 69245 18655
0 18657 5 1 1 18656
0 18658 7 2 2 72766 78561
0 18659 5 1 1 91337
0 18660 7 1 2 91248 91338
0 18661 5 1 1 18660
0 18662 7 1 2 73187 82224
0 18663 5 1 1 18662
0 18664 7 1 2 75200 18663
0 18665 5 1 1 18664
0 18666 7 1 2 18661 18665
0 18667 7 1 2 18657 18666
0 18668 7 1 2 18646 18667
0 18669 7 1 2 18622 18668
0 18670 5 1 1 18669
0 18671 7 1 2 64955 18670
0 18672 5 1 1 18671
0 18673 7 1 2 62296 82800
0 18674 5 1 1 18673
0 18675 7 1 2 61299 18674
0 18676 5 1 1 18675
0 18677 7 1 2 82284 18676
0 18678 5 1 1 18677
0 18679 7 1 2 73188 75797
0 18680 5 1 1 18679
0 18681 7 1 2 77688 18680
0 18682 5 1 1 18681
0 18683 7 1 2 72332 88762
0 18684 5 1 1 18683
0 18685 7 1 2 77709 18684
0 18686 7 1 2 18682 18685
0 18687 7 1 2 18678 18686
0 18688 5 1 1 18687
0 18689 7 1 2 65185 18688
0 18690 5 1 1 18689
0 18691 7 4 2 62620 77705
0 18692 5 1 1 91339
0 18693 7 1 2 72589 76703
0 18694 7 1 2 91340 18693
0 18695 5 1 1 18694
0 18696 7 1 2 18690 18695
0 18697 5 1 1 18696
0 18698 7 1 2 66464 18697
0 18699 5 1 1 18698
0 18700 7 1 2 77307 70953
0 18701 5 1 1 18700
0 18702 7 1 2 77258 80272
0 18703 5 1 1 18702
0 18704 7 1 2 83477 18703
0 18705 5 1 1 18704
0 18706 7 1 2 62955 18705
0 18707 5 1 1 18706
0 18708 7 1 2 69657 87237
0 18709 5 1 1 18708
0 18710 7 1 2 18707 18709
0 18711 5 1 1 18710
0 18712 7 1 2 62091 18711
0 18713 5 1 1 18712
0 18714 7 1 2 18106 91299
0 18715 5 1 1 18714
0 18716 7 1 2 72590 18715
0 18717 5 1 1 18716
0 18718 7 1 2 18713 18717
0 18719 5 1 1 18718
0 18720 7 1 2 18701 18719
0 18721 5 1 1 18720
0 18722 7 6 2 62956 70485
0 18723 5 1 1 91343
0 18724 7 2 2 80273 72333
0 18725 7 1 2 91344 91349
0 18726 5 1 1 18725
0 18727 7 1 2 9425 18726
0 18728 5 1 1 18727
0 18729 7 1 2 62621 18728
0 18730 5 1 1 18729
0 18731 7 1 2 90951 91297
0 18732 5 1 1 18731
0 18733 7 1 2 18730 18732
0 18734 5 1 1 18733
0 18735 7 1 2 80604 18734
0 18736 5 1 1 18735
0 18737 7 2 2 70791 91310
0 18738 7 1 2 76916 91351
0 18739 5 1 1 18738
0 18740 7 1 2 90407 18739
0 18741 5 2 1 18740
0 18742 7 1 2 83820 91353
0 18743 5 1 1 18742
0 18744 7 1 2 18736 18743
0 18745 7 1 2 18721 18744
0 18746 7 1 2 18699 18745
0 18747 7 1 2 18672 18746
0 18748 7 1 2 18590 18747
0 18749 7 1 2 18522 18748
0 18750 5 1 1 18749
0 18751 7 1 2 80860 18750
0 18752 5 1 1 18751
0 18753 7 3 2 66670 71393
0 18754 7 1 2 76494 83077
0 18755 5 1 1 18754
0 18756 7 1 2 72863 83873
0 18757 7 11 2 60490 67953
0 18758 5 1 1 91358
0 18759 7 1 2 89125 18758
0 18760 7 1 2 18756 18759
0 18761 7 1 2 87813 18760
0 18762 5 1 1 18761
0 18763 7 1 2 18755 18762
0 18764 5 1 1 18763
0 18765 7 1 2 91355 18764
0 18766 5 1 1 18765
0 18767 7 2 2 67954 86420
0 18768 7 1 2 72441 3574
0 18769 5 1 1 18768
0 18770 7 2 2 64273 74759
0 18771 7 1 2 18769 91371
0 18772 5 1 1 18771
0 18773 7 5 2 64497 75905
0 18774 5 2 1 91373
0 18775 7 1 2 66009 91374
0 18776 5 1 1 18775
0 18777 7 2 2 18772 18776
0 18778 7 1 2 66010 78315
0 18779 5 1 1 18778
0 18780 7 1 2 72098 72442
0 18781 5 1 1 18780
0 18782 7 1 2 64274 18781
0 18783 5 1 1 18782
0 18784 7 1 2 86950 18783
0 18785 7 1 2 18779 18784
0 18786 5 1 1 18785
0 18787 7 1 2 64713 18786
0 18788 5 1 1 18787
0 18789 7 1 2 91380 18788
0 18790 5 1 1 18789
0 18791 7 1 2 70050 18790
0 18792 5 1 1 18791
0 18793 7 4 2 64275 69067
0 18794 5 3 1 91382
0 18795 7 2 2 70792 91383
0 18796 7 1 2 80298 70923
0 18797 7 1 2 91389 18796
0 18798 5 1 1 18797
0 18799 7 1 2 18792 18798
0 18800 5 1 1 18799
0 18801 7 1 2 91369 18800
0 18802 5 1 1 18801
0 18803 7 1 2 18766 18802
0 18804 5 1 1 18803
0 18805 7 1 2 67047 18804
0 18806 5 1 1 18805
0 18807 7 1 2 71030 81726
0 18808 7 1 2 88374 18807
0 18809 5 1 1 18808
0 18810 7 1 2 66247 76509
0 18811 5 2 1 18810
0 18812 7 4 2 65383 61039
0 18813 7 1 2 91356 91393
0 18814 7 1 2 91391 18813
0 18815 5 1 1 18814
0 18816 7 1 2 18809 18815
0 18817 5 1 1 18816
0 18818 7 1 2 67955 18817
0 18819 5 1 1 18818
0 18820 7 1 2 18806 18819
0 18821 5 1 1 18820
0 18822 7 1 2 67581 18821
0 18823 5 1 1 18822
0 18824 7 2 2 65384 78126
0 18825 5 3 1 91397
0 18826 7 1 2 77386 91399
0 18827 5 1 1 18826
0 18828 7 1 2 75785 18827
0 18829 5 1 1 18828
0 18830 7 1 2 74965 89718
0 18831 5 1 1 18830
0 18832 7 1 2 18829 18831
0 18833 5 1 1 18832
0 18834 7 1 2 85592 88614
0 18835 7 1 2 18833 18834
0 18836 5 1 1 18835
0 18837 7 1 2 18823 18836
0 18838 5 1 1 18837
0 18839 7 1 2 61494 18838
0 18840 5 1 1 18839
0 18841 7 1 2 18752 18840
0 18842 5 1 1 18841
0 18843 7 1 2 68315 18842
0 18844 5 1 1 18843
0 18845 7 4 2 60491 61300
0 18846 7 3 2 66671 91402
0 18847 5 1 1 91406
0 18848 7 6 2 66465 86536
0 18849 5 2 1 91409
0 18850 7 1 2 80367 91415
0 18851 5 4 1 18850
0 18852 7 1 2 80489 91417
0 18853 5 1 1 18852
0 18854 7 1 2 18847 18853
0 18855 5 1 1 18854
0 18856 7 1 2 75940 18855
0 18857 5 1 1 18856
0 18858 7 1 2 85301 88104
0 18859 7 1 2 88751 18858
0 18860 5 1 1 18859
0 18861 7 1 2 80344 18860
0 18862 5 1 1 18861
0 18863 7 1 2 84596 18862
0 18864 5 1 1 18863
0 18865 7 1 2 18857 18864
0 18866 5 1 1 18865
0 18867 7 1 2 89437 18866
0 18868 5 1 1 18867
0 18869 7 1 2 80274 89199
0 18870 5 1 1 18869
0 18871 7 1 2 89208 18870
0 18872 5 1 1 18871
0 18873 7 5 2 60492 88082
0 18874 5 1 1 91421
0 18875 7 2 2 80268 79088
0 18876 5 6 1 91426
0 18877 7 1 2 91422 91428
0 18878 7 1 2 18872 18877
0 18879 5 1 1 18878
0 18880 7 1 2 18868 18879
0 18881 5 1 1 18880
0 18882 7 1 2 67582 18881
0 18883 5 1 1 18882
0 18884 7 1 2 67279 7160
0 18885 5 2 1 18884
0 18886 7 1 2 64276 91434
0 18887 5 1 1 18886
0 18888 7 1 2 76406 18887
0 18889 5 3 1 18888
0 18890 7 1 2 72334 91436
0 18891 5 1 1 18890
0 18892 7 1 2 89202 18891
0 18893 5 1 1 18892
0 18894 7 1 2 64498 18893
0 18895 5 1 1 18894
0 18896 7 1 2 76339 82520
0 18897 5 1 1 18896
0 18898 7 1 2 71110 18897
0 18899 5 1 1 18898
0 18900 7 1 2 18895 18899
0 18901 5 1 1 18900
0 18902 7 1 2 62622 18901
0 18903 5 1 1 18902
0 18904 7 6 2 64277 72335
0 18905 7 1 2 62623 91439
0 18906 5 1 1 18905
0 18907 7 1 2 91291 18906
0 18908 5 2 1 18907
0 18909 7 1 2 70415 91445
0 18910 5 1 1 18909
0 18911 7 1 2 70548 86399
0 18912 5 1 1 18911
0 18913 7 1 2 71519 18912
0 18914 7 1 2 18910 18913
0 18915 7 1 2 18903 18914
0 18916 5 1 1 18915
0 18917 7 1 2 62957 18916
0 18918 5 1 1 18917
0 18919 7 1 2 72633 87428
0 18920 5 1 1 18919
0 18921 7 1 2 70793 88413
0 18922 5 1 1 18921
0 18923 7 1 2 91283 18922
0 18924 5 1 1 18923
0 18925 7 1 2 82573 18924
0 18926 5 1 1 18925
0 18927 7 1 2 64714 89048
0 18928 5 3 1 18927
0 18929 7 1 2 78939 91447
0 18930 5 2 1 18929
0 18931 7 1 2 70794 91450
0 18932 5 1 1 18931
0 18933 7 1 2 90333 18932
0 18934 7 1 2 18926 18933
0 18935 5 1 1 18934
0 18936 7 1 2 64278 18935
0 18937 5 1 1 18936
0 18938 7 1 2 18920 18937
0 18939 5 1 1 18938
0 18940 7 1 2 70312 18939
0 18941 5 1 1 18940
0 18942 7 1 2 77236 90952
0 18943 5 1 1 18942
0 18944 7 1 2 88928 18943
0 18945 5 1 1 18944
0 18946 7 1 2 62624 18945
0 18947 5 1 1 18946
0 18948 7 1 2 59846 88523
0 18949 5 1 1 18948
0 18950 7 1 2 62958 18949
0 18951 5 1 1 18950
0 18952 7 1 2 18947 18951
0 18953 5 1 1 18952
0 18954 7 1 2 69246 18953
0 18955 5 1 1 18954
0 18956 7 2 2 67956 74893
0 18957 5 4 1 91452
0 18958 7 1 2 73981 91454
0 18959 5 1 1 18958
0 18960 7 2 2 78095 18959
0 18961 7 1 2 83874 91458
0 18962 5 1 1 18961
0 18963 7 1 2 82787 18962
0 18964 5 1 1 18963
0 18965 7 4 2 67048 76495
0 18966 7 1 2 72143 91460
0 18967 5 1 1 18966
0 18968 7 2 2 72421 18967
0 18969 7 1 2 62959 91464
0 18970 5 1 1 18969
0 18971 7 1 2 60315 18970
0 18972 7 1 2 18964 18971
0 18973 7 1 2 18955 18972
0 18974 5 1 1 18973
0 18975 7 1 2 70795 18974
0 18976 5 1 1 18975
0 18977 7 3 2 61040 69400
0 18978 7 1 2 81898 91466
0 18979 5 1 1 18978
0 18980 7 1 2 90329 18979
0 18981 5 1 1 18980
0 18982 7 1 2 61495 18981
0 18983 7 1 2 18976 18982
0 18984 7 1 2 18941 18983
0 18985 7 1 2 18918 18984
0 18986 5 1 1 18985
0 18987 7 1 2 74420 72221
0 18988 5 1 1 18987
0 18989 7 1 2 77424 18988
0 18990 5 1 1 18989
0 18991 7 1 2 83005 78910
0 18992 7 1 2 18990 18991
0 18993 5 1 1 18992
0 18994 7 1 2 61301 18993
0 18995 5 1 1 18994
0 18996 7 4 2 59847 75009
0 18997 5 1 1 91469
0 18998 7 1 2 89719 91470
0 18999 5 1 1 18998
0 19000 7 1 2 67280 77398
0 19001 5 1 1 19000
0 19002 7 1 2 18999 19001
0 19003 5 1 1 19002
0 19004 7 1 2 69532 19003
0 19005 5 1 1 19004
0 19006 7 1 2 76553 82977
0 19007 5 1 1 19006
0 19008 7 1 2 83041 19007
0 19009 5 1 1 19008
0 19010 7 1 2 71708 19009
0 19011 5 1 1 19010
0 19012 7 1 2 60316 82947
0 19013 5 1 1 19012
0 19014 7 1 2 66466 19013
0 19015 7 1 2 19011 19014
0 19016 7 1 2 19005 19015
0 19017 7 1 2 18995 19016
0 19018 5 1 1 19017
0 19019 7 1 2 60493 19018
0 19020 7 1 2 18986 19019
0 19021 5 1 1 19020
0 19022 7 4 2 71709 73466
0 19023 7 1 2 83075 82873
0 19024 7 1 2 91473 19023
0 19025 5 1 1 19024
0 19026 7 1 2 19021 19025
0 19027 5 1 1 19026
0 19028 7 1 2 61689 19027
0 19029 5 1 1 19028
0 19030 7 1 2 18883 19029
0 19031 5 1 1 19030
0 19032 7 1 2 63408 19031
0 19033 5 1 1 19032
0 19034 7 1 2 68644 19033
0 19035 7 1 2 18844 19034
0 19036 5 1 1 19035
0 19037 7 2 2 73667 82607
0 19038 7 1 2 76340 77898
0 19039 7 1 2 89142 19038
0 19040 5 1 1 19039
0 19041 7 1 2 77804 19040
0 19042 5 1 1 19041
0 19043 7 1 2 91477 19042
0 19044 5 2 1 19043
0 19045 7 4 2 62625 69533
0 19046 7 1 2 78966 91481
0 19047 5 3 1 19046
0 19048 7 1 2 83930 91485
0 19049 5 1 1 19048
0 19050 7 1 2 85901 19049
0 19051 5 2 1 19050
0 19052 7 1 2 67281 77899
0 19053 7 1 2 73189 19052
0 19054 5 1 1 19053
0 19055 7 1 2 77805 19054
0 19056 5 1 1 19055
0 19057 7 1 2 74679 19056
0 19058 5 2 1 19057
0 19059 7 1 2 80642 89420
0 19060 5 2 1 19059
0 19061 7 2 2 67957 71468
0 19062 7 1 2 85302 91494
0 19063 5 1 1 19062
0 19064 7 1 2 83915 19063
0 19065 5 1 1 19064
0 19066 7 1 2 59499 89463
0 19067 7 1 2 19065 19066
0 19068 5 1 1 19067
0 19069 7 1 2 91492 19068
0 19070 5 1 1 19069
0 19071 7 1 2 60903 19070
0 19072 5 1 1 19071
0 19073 7 1 2 91490 19072
0 19074 5 1 1 19073
0 19075 7 1 2 67583 19074
0 19076 5 1 1 19075
0 19077 7 1 2 91488 19076
0 19078 5 1 1 19077
0 19079 7 1 2 59848 19078
0 19080 5 1 1 19079
0 19081 7 1 2 91479 19080
0 19082 5 1 1 19081
0 19083 7 1 2 89438 19082
0 19084 5 1 1 19083
0 19085 7 1 2 61496 89154
0 19086 5 1 1 19085
0 19087 7 1 2 71469 89542
0 19088 5 1 1 19087
0 19089 7 1 2 64956 19088
0 19090 5 1 1 19089
0 19091 7 1 2 61302 19090
0 19092 5 1 1 19091
0 19093 7 1 2 70153 76580
0 19094 5 1 1 19093
0 19095 7 1 2 66467 19094
0 19096 7 1 2 19092 19095
0 19097 5 1 1 19096
0 19098 7 1 2 67584 19097
0 19099 7 1 2 19086 19098
0 19100 5 1 1 19099
0 19101 7 1 2 80208 77672
0 19102 7 1 2 81934 19101
0 19103 5 1 1 19102
0 19104 7 1 2 75277 19103
0 19105 5 1 1 19104
0 19106 7 3 2 76443 79171
0 19107 5 1 1 91496
0 19108 7 1 2 61497 73130
0 19109 7 1 2 19107 19108
0 19110 5 1 1 19109
0 19111 7 1 2 19105 19110
0 19112 5 1 1 19111
0 19113 7 1 2 62626 19112
0 19114 5 1 1 19113
0 19115 7 3 2 69534 76179
0 19116 5 1 1 91499
0 19117 7 1 2 83308 19116
0 19118 5 1 1 19117
0 19119 7 1 2 88615 19118
0 19120 5 1 1 19119
0 19121 7 1 2 75278 76672
0 19122 7 1 2 90073 19121
0 19123 5 1 1 19122
0 19124 7 1 2 67958 19123
0 19125 7 1 2 19120 19124
0 19126 7 1 2 19114 19125
0 19127 7 1 2 19100 19126
0 19128 5 1 1 19127
0 19129 7 1 2 59849 76205
0 19130 5 3 1 19129
0 19131 7 1 2 71370 91502
0 19132 5 1 1 19131
0 19133 7 1 2 70600 19132
0 19134 5 1 1 19133
0 19135 7 1 2 78475 89483
0 19136 5 1 1 19135
0 19137 7 5 2 67585 73407
0 19138 7 1 2 60904 73711
0 19139 7 1 2 91505 19138
0 19140 5 1 1 19139
0 19141 7 1 2 19136 19140
0 19142 5 1 1 19141
0 19143 7 1 2 59500 19142
0 19144 5 1 1 19143
0 19145 7 1 2 19134 19144
0 19146 5 1 1 19145
0 19147 7 1 2 61041 19146
0 19148 5 1 1 19147
0 19149 7 1 2 61303 74841
0 19150 5 1 1 19149
0 19151 7 1 2 81806 83046
0 19152 5 1 1 19151
0 19153 7 1 2 19150 19152
0 19154 5 1 1 19153
0 19155 7 1 2 75279 19154
0 19156 5 1 1 19155
0 19157 7 1 2 86830 19156
0 19158 7 1 2 19148 19157
0 19159 5 1 1 19158
0 19160 7 1 2 19128 19159
0 19161 5 1 1 19160
0 19162 7 1 2 81049 79575
0 19163 5 1 1 19162
0 19164 7 1 2 68316 19163
0 19165 7 1 2 19161 19164
0 19166 5 1 1 19165
0 19167 7 1 2 74066 81565
0 19168 5 1 1 19167
0 19169 7 1 2 82898 19168
0 19170 5 1 1 19169
0 19171 7 1 2 80258 90789
0 19172 5 1 1 19171
0 19173 7 1 2 19170 19172
0 19174 5 1 1 19173
0 19175 7 1 2 75280 19174
0 19176 5 1 1 19175
0 19177 7 1 2 83123 76379
0 19178 5 1 1 19177
0 19179 7 4 2 61304 72945
0 19180 7 1 2 88011 91510
0 19181 5 1 1 19180
0 19182 7 1 2 75561 19181
0 19183 5 1 1 19182
0 19184 7 1 2 80259 19183
0 19185 5 1 1 19184
0 19186 7 1 2 19178 19185
0 19187 7 1 2 19176 19186
0 19188 5 1 1 19187
0 19189 7 1 2 69535 19188
0 19190 5 1 1 19189
0 19191 7 1 2 72946 89544
0 19192 5 1 1 19191
0 19193 7 1 2 75562 19192
0 19194 5 4 1 19193
0 19195 7 1 2 67959 77322
0 19196 5 2 1 19195
0 19197 7 1 2 74210 91518
0 19198 5 1 1 19197
0 19199 7 1 2 91514 19198
0 19200 5 1 1 19199
0 19201 7 1 2 63409 19200
0 19202 7 1 2 19190 19201
0 19203 5 1 1 19202
0 19204 7 1 2 61690 19203
0 19205 7 1 2 19166 19204
0 19206 5 1 1 19205
0 19207 7 1 2 19084 19206
0 19208 5 1 1 19207
0 19209 7 1 2 60494 19208
0 19210 5 1 1 19209
0 19211 7 1 2 83916 89625
0 19212 5 2 1 19211
0 19213 7 1 2 69536 91520
0 19214 5 1 1 19213
0 19215 7 1 2 83917 90032
0 19216 5 1 1 19215
0 19217 7 1 2 67282 19216
0 19218 5 1 1 19217
0 19219 7 1 2 19214 19218
0 19220 5 1 1 19219
0 19221 7 1 2 83184 19220
0 19222 5 1 1 19221
0 19223 7 1 2 91493 19222
0 19224 5 1 1 19223
0 19225 7 1 2 60905 19224
0 19226 5 1 1 19225
0 19227 7 1 2 91491 19226
0 19228 5 1 1 19227
0 19229 7 1 2 67586 19228
0 19230 5 1 1 19229
0 19231 7 1 2 91489 19230
0 19232 5 1 1 19231
0 19233 7 1 2 59850 19232
0 19234 5 1 1 19233
0 19235 7 1 2 91480 19234
0 19236 5 1 1 19235
0 19237 7 2 2 72947 86231
0 19238 7 1 2 19236 91522
0 19239 5 1 1 19238
0 19240 7 1 2 63705 19239
0 19241 7 1 2 19210 19240
0 19242 5 1 1 19241
0 19243 7 1 2 19036 19242
0 19244 5 1 1 19243
0 19245 7 9 2 59851 69178
0 19246 5 8 1 91524
0 19247 7 6 2 69537 88990
0 19248 5 1 1 91541
0 19249 7 1 2 91525 91542
0 19250 5 2 1 19249
0 19251 7 1 2 62297 72144
0 19252 5 2 1 19251
0 19253 7 3 2 66011 71778
0 19254 5 5 1 91551
0 19255 7 2 2 69538 91554
0 19256 5 1 1 91559
0 19257 7 1 2 74760 19256
0 19258 5 1 1 19257
0 19259 7 1 2 91549 19258
0 19260 5 1 1 19259
0 19261 7 1 2 64715 19260
0 19262 5 1 1 19261
0 19263 7 1 2 60115 91381
0 19264 7 1 2 19262 19263
0 19265 5 1 1 19264
0 19266 7 1 2 91547 19265
0 19267 5 1 1 19266
0 19268 7 1 2 83362 88559
0 19269 5 1 1 19268
0 19270 7 2 2 66248 19269
0 19271 5 1 1 91561
0 19272 7 1 2 60317 19271
0 19273 7 1 2 19267 19272
0 19274 5 1 1 19273
0 19275 7 1 2 67587 19274
0 19276 5 1 1 19275
0 19277 7 1 2 62298 89063
0 19278 5 3 1 19277
0 19279 7 2 2 78476 91563
0 19280 5 1 1 91566
0 19281 7 1 2 91562 91567
0 19282 5 1 1 19281
0 19283 7 1 2 19276 19282
0 19284 5 1 1 19283
0 19285 7 1 2 67049 19284
0 19286 5 1 1 19285
0 19287 7 1 2 78116 90708
0 19288 5 1 1 19287
0 19289 7 1 2 61305 19288
0 19290 5 1 1 19289
0 19291 7 1 2 71357 90957
0 19292 5 1 1 19291
0 19293 7 1 2 19290 19292
0 19294 5 1 1 19293
0 19295 7 1 2 71779 19294
0 19296 5 1 1 19295
0 19297 7 1 2 73696 76007
0 19298 5 1 1 19297
0 19299 7 1 2 71195 19298
0 19300 5 1 1 19299
0 19301 7 1 2 62092 19300
0 19302 5 1 1 19301
0 19303 7 1 2 62627 72462
0 19304 5 1 1 19303
0 19305 7 1 2 60318 19304
0 19306 7 1 2 19302 19305
0 19307 5 1 1 19306
0 19308 7 1 2 61306 19307
0 19309 5 1 1 19308
0 19310 7 1 2 62299 71453
0 19311 5 1 1 19310
0 19312 7 1 2 67588 19311
0 19313 5 1 1 19312
0 19314 7 1 2 61307 19313
0 19315 5 1 1 19314
0 19316 7 2 2 62093 71358
0 19317 5 1 1 91568
0 19318 7 1 2 71978 91569
0 19319 5 1 1 19318
0 19320 7 1 2 19315 19319
0 19321 5 1 1 19320
0 19322 7 1 2 72336 19321
0 19323 5 1 1 19322
0 19324 7 1 2 2444 74479
0 19325 5 1 1 19324
0 19326 7 1 2 73867 19325
0 19327 5 1 1 19326
0 19328 7 4 2 66249 74119
0 19329 5 3 1 91570
0 19330 7 1 2 73814 91571
0 19331 7 1 2 19327 19330
0 19332 5 1 1 19331
0 19333 7 1 2 67960 19332
0 19334 7 1 2 19323 19333
0 19335 7 1 2 19309 19334
0 19336 7 1 2 19296 19335
0 19337 7 1 2 19286 19336
0 19338 5 1 1 19337
0 19339 7 1 2 66012 77049
0 19340 5 5 1 19339
0 19341 7 1 2 59852 91577
0 19342 5 1 1 19341
0 19343 7 1 2 71196 74097
0 19344 5 2 1 19343
0 19345 7 1 2 19342 91582
0 19346 5 1 1 19345
0 19347 7 1 2 60906 19346
0 19348 5 1 1 19347
0 19349 7 1 2 70051 19348
0 19350 5 1 1 19349
0 19351 7 1 2 78487 19350
0 19352 5 1 1 19351
0 19353 7 1 2 60795 90953
0 19354 7 2 2 88448 19353
0 19355 5 1 1 91584
0 19356 7 1 2 59305 91585
0 19357 5 1 1 19356
0 19358 7 1 2 82712 19357
0 19359 7 1 2 19352 19358
0 19360 5 1 1 19359
0 19361 7 1 2 69106 19360
0 19362 5 1 1 19361
0 19363 7 1 2 64716 89064
0 19364 5 2 1 19363
0 19365 7 2 2 66013 74120
0 19366 5 9 1 91588
0 19367 7 3 2 67283 91590
0 19368 7 1 2 91586 91599
0 19369 5 1 1 19368
0 19370 7 3 2 78477 72222
0 19371 5 1 1 91602
0 19372 7 1 2 70154 74139
0 19373 5 1 1 19372
0 19374 7 1 2 19371 19373
0 19375 7 1 2 19369 19374
0 19376 5 1 1 19375
0 19377 7 1 2 59501 19376
0 19378 5 1 1 19377
0 19379 7 1 2 70155 91587
0 19380 5 1 1 19379
0 19381 7 1 2 65186 70249
0 19382 7 1 2 91122 19381
0 19383 7 1 2 19380 19382
0 19384 7 1 2 19378 19383
0 19385 7 1 2 19362 19384
0 19386 5 1 1 19385
0 19387 7 1 2 19338 19386
0 19388 5 1 1 19387
0 19389 7 1 2 60319 91572
0 19390 5 1 1 19389
0 19391 7 1 2 19388 19390
0 19392 5 1 1 19391
0 19393 7 1 2 61498 19392
0 19394 5 1 1 19393
0 19395 7 1 2 67284 80223
0 19396 5 1 1 19395
0 19397 7 3 2 72864 81807
0 19398 5 1 1 91605
0 19399 7 1 2 19396 19398
0 19400 5 1 1 19399
0 19401 7 1 2 67050 19400
0 19402 5 1 1 19401
0 19403 7 1 2 67589 91392
0 19404 5 1 1 19403
0 19405 7 1 2 19402 19404
0 19406 5 1 1 19405
0 19407 7 1 2 61042 19406
0 19408 5 1 1 19407
0 19409 7 1 2 66250 74211
0 19410 5 2 1 19409
0 19411 7 1 2 69539 91608
0 19412 5 2 1 19411
0 19413 7 1 2 5761 91610
0 19414 5 1 1 19413
0 19415 7 1 2 73010 19414
0 19416 5 1 1 19415
0 19417 7 1 2 19408 19416
0 19418 5 1 1 19417
0 19419 7 1 2 82402 19418
0 19420 5 1 1 19419
0 19421 7 2 2 61308 91591
0 19422 5 1 1 91612
0 19423 7 1 2 66251 85085
0 19424 5 2 1 19423
0 19425 7 1 2 59853 91614
0 19426 5 1 1 19425
0 19427 7 1 2 19422 19426
0 19428 5 1 1 19427
0 19429 7 1 2 71710 19428
0 19430 5 1 1 19429
0 19431 7 3 2 61043 75712
0 19432 7 1 2 67590 91616
0 19433 5 1 1 19432
0 19434 7 1 2 19430 19433
0 19435 5 1 1 19434
0 19436 7 1 2 69540 19435
0 19437 5 1 1 19436
0 19438 7 1 2 71647 85083
0 19439 5 1 1 19438
0 19440 7 1 2 59854 91613
0 19441 5 1 1 19440
0 19442 7 1 2 65187 19441
0 19443 5 1 1 19442
0 19444 7 1 2 88767 19443
0 19445 5 1 1 19444
0 19446 7 1 2 19439 19445
0 19447 7 1 2 19437 19446
0 19448 5 1 1 19447
0 19449 7 1 2 67285 19448
0 19450 5 1 1 19449
0 19451 7 1 2 83350 71272
0 19452 5 1 1 19451
0 19453 7 1 2 60320 19452
0 19454 5 1 1 19453
0 19455 7 1 2 67051 77683
0 19456 7 1 2 91606 19455
0 19457 5 1 1 19456
0 19458 7 1 2 61309 72223
0 19459 5 1 1 19458
0 19460 7 1 2 65188 19459
0 19461 5 2 1 19460
0 19462 7 1 2 74184 91619
0 19463 5 1 1 19462
0 19464 7 1 2 19457 19463
0 19465 7 1 2 19454 19464
0 19466 7 1 2 19450 19465
0 19467 5 1 1 19466
0 19468 7 1 2 62960 19467
0 19469 5 1 1 19468
0 19470 7 1 2 19420 19469
0 19471 5 1 1 19470
0 19472 7 1 2 60116 19471
0 19473 5 1 1 19472
0 19474 7 1 2 60907 7551
0 19475 5 1 1 19474
0 19476 7 1 2 81655 19475
0 19477 5 2 1 19476
0 19478 7 1 2 82833 91621
0 19479 5 1 1 19478
0 19480 7 1 2 74043 90029
0 19481 5 1 1 19480
0 19482 7 1 2 19479 19481
0 19483 5 1 1 19482
0 19484 7 1 2 69541 19483
0 19485 5 1 1 19484
0 19486 7 1 2 82834 76312
0 19487 5 1 1 19486
0 19488 7 1 2 19485 19487
0 19489 5 1 1 19488
0 19490 7 1 2 71197 19489
0 19491 5 1 1 19490
0 19492 7 1 2 82926 74861
0 19493 5 1 1 19492
0 19494 7 1 2 13192 19493
0 19495 5 1 1 19494
0 19496 7 1 2 76496 19495
0 19497 5 1 1 19496
0 19498 7 5 2 59502 62961
0 19499 7 2 2 69463 91623
0 19500 5 2 1 91628
0 19501 7 1 2 69542 91629
0 19502 5 1 1 19501
0 19503 7 1 2 78478 82403
0 19504 5 1 1 19503
0 19505 7 1 2 19502 19504
0 19506 5 1 1 19505
0 19507 7 1 2 91620 19506
0 19508 5 1 1 19507
0 19509 7 1 2 19497 19508
0 19510 5 1 1 19509
0 19511 7 1 2 67052 19510
0 19512 5 1 1 19511
0 19513 7 1 2 82835 91304
0 19514 7 1 2 88768 19513
0 19515 5 1 1 19514
0 19516 7 1 2 19512 19515
0 19517 5 1 1 19516
0 19518 7 1 2 67286 19517
0 19519 5 1 1 19518
0 19520 7 1 2 66252 72878
0 19521 5 1 1 19520
0 19522 7 1 2 82404 19521
0 19523 5 1 1 19522
0 19524 7 2 2 59503 73912
0 19525 5 1 1 91632
0 19526 7 1 2 74185 91305
0 19527 5 1 1 19526
0 19528 7 1 2 19525 19527
0 19529 5 1 1 19528
0 19530 7 1 2 62962 19529
0 19531 5 1 1 19530
0 19532 7 1 2 19523 19531
0 19533 5 1 1 19532
0 19534 7 1 2 60321 19533
0 19535 5 1 1 19534
0 19536 7 1 2 68317 19535
0 19537 7 1 2 19519 19536
0 19538 7 1 2 19491 19537
0 19539 7 1 2 19473 19538
0 19540 7 1 2 19394 19539
0 19541 5 1 1 19540
0 19542 7 2 2 83244 83052
0 19543 5 2 1 91634
0 19544 7 1 2 79899 91636
0 19545 5 1 1 19544
0 19546 7 1 2 61310 19545
0 19547 5 1 1 19546
0 19548 7 1 2 76554 72186
0 19549 5 1 1 19548
0 19550 7 1 2 78390 19549
0 19551 5 1 1 19550
0 19552 7 1 2 61499 19551
0 19553 5 1 1 19552
0 19554 7 1 2 19547 19553
0 19555 5 1 1 19554
0 19556 7 1 2 69543 19555
0 19557 5 1 1 19556
0 19558 7 1 2 81902 15203
0 19559 5 1 1 19558
0 19560 7 1 2 79883 19559
0 19561 5 1 1 19560
0 19562 7 1 2 19557 19561
0 19563 5 1 1 19562
0 19564 7 1 2 90796 19563
0 19565 5 1 1 19564
0 19566 7 1 2 3849 90800
0 19567 5 1 1 19566
0 19568 7 1 2 67287 19567
0 19569 5 1 1 19568
0 19570 7 2 2 70156 89545
0 19571 5 1 1 91638
0 19572 7 1 2 74767 91639
0 19573 5 1 1 19572
0 19574 7 1 2 19569 19573
0 19575 5 1 1 19574
0 19576 7 1 2 69544 19575
0 19577 5 1 1 19576
0 19578 7 1 2 11069 19577
0 19579 5 1 1 19578
0 19580 7 1 2 67961 19579
0 19581 5 1 1 19580
0 19582 7 1 2 63410 19581
0 19583 7 1 2 19565 19582
0 19584 5 1 1 19583
0 19585 7 1 2 68645 19584
0 19586 7 1 2 19541 19585
0 19587 5 1 1 19586
0 19588 7 3 2 76768 91049
0 19589 7 2 2 71711 91640
0 19590 5 2 1 91643
0 19591 7 1 2 6677 91645
0 19592 5 1 1 19591
0 19593 7 1 2 88903 19592
0 19594 5 1 1 19593
0 19595 7 1 2 74631 91641
0 19596 5 1 1 19595
0 19597 7 1 2 71659 19596
0 19598 5 1 1 19597
0 19599 7 1 2 72099 19598
0 19600 5 1 1 19599
0 19601 7 4 2 89159 91335
0 19602 5 2 1 91647
0 19603 7 1 2 71520 70892
0 19604 7 1 2 91648 19603
0 19605 5 1 1 19604
0 19606 7 1 2 19600 19605
0 19607 7 1 2 19594 19606
0 19608 5 1 1 19607
0 19609 7 1 2 67591 19608
0 19610 5 1 1 19609
0 19611 7 1 2 71856 19610
0 19612 5 1 1 19611
0 19613 7 1 2 61500 89703
0 19614 7 1 2 19612 19613
0 19615 5 1 1 19614
0 19616 7 1 2 19587 19615
0 19617 5 1 1 19616
0 19618 7 1 2 81171 19617
0 19619 5 1 1 19618
0 19620 7 11 2 65385 75563
0 19621 5 75 1 91653
0 19622 7 4 2 61044 91664
0 19623 7 1 2 83009 91739
0 19624 5 1 1 19623
0 19625 7 1 2 76769 89872
0 19626 5 1 1 19625
0 19627 7 1 2 66468 88731
0 19628 5 2 1 19627
0 19629 7 1 2 75428 84838
0 19630 7 1 2 90633 19629
0 19631 7 1 2 91743 19630
0 19632 5 1 1 19631
0 19633 7 1 2 19626 19632
0 19634 5 1 1 19633
0 19635 7 1 2 75786 19634
0 19636 5 1 1 19635
0 19637 7 1 2 19624 19636
0 19638 5 1 1 19637
0 19639 7 1 2 67592 19638
0 19640 5 1 1 19639
0 19641 7 1 2 65386 90074
0 19642 5 2 1 19641
0 19643 7 1 2 76770 83035
0 19644 7 1 2 91745 19643
0 19645 5 1 1 19644
0 19646 7 1 2 19640 19645
0 19647 5 1 1 19646
0 19648 7 1 2 61691 19647
0 19649 5 1 1 19648
0 19650 7 4 2 80101 89636
0 19651 7 1 2 66014 75790
0 19652 5 1 1 19651
0 19653 7 1 2 83899 19652
0 19654 5 1 1 19653
0 19655 7 2 2 82650 79285
0 19656 7 1 2 83609 91751
0 19657 5 1 1 19656
0 19658 7 1 2 19654 19657
0 19659 5 1 1 19658
0 19660 7 1 2 67593 19659
0 19661 5 1 1 19660
0 19662 7 1 2 61501 78886
0 19663 5 1 1 19662
0 19664 7 1 2 19661 19663
0 19665 5 1 1 19664
0 19666 7 1 2 91747 19665
0 19667 5 1 1 19666
0 19668 7 1 2 19649 19667
0 19669 5 1 1 19668
0 19670 7 1 2 63706 19669
0 19671 5 1 1 19670
0 19672 7 13 2 60495 67594
0 19673 5 2 1 91753
0 19674 7 2 2 84474 91754
0 19675 5 3 1 91768
0 19676 7 1 2 89260 91769
0 19677 5 1 1 19676
0 19678 7 1 2 81389 84334
0 19679 7 1 2 89285 19678
0 19680 5 1 1 19679
0 19681 7 1 2 19677 19680
0 19682 5 1 1 19681
0 19683 7 1 2 78127 19682
0 19684 5 1 1 19683
0 19685 7 5 2 59306 71871
0 19686 5 2 1 91773
0 19687 7 1 2 80456 79374
0 19688 7 1 2 91774 19687
0 19689 7 1 2 89310 19688
0 19690 5 1 1 19689
0 19691 7 1 2 19684 19690
0 19692 5 1 1 19691
0 19693 7 1 2 67288 19692
0 19694 5 1 1 19693
0 19695 7 3 2 84047 76105
0 19696 5 1 1 91780
0 19697 7 1 2 84425 91781
0 19698 7 1 2 89311 19697
0 19699 5 1 1 19698
0 19700 7 1 2 19694 19699
0 19701 5 1 1 19700
0 19702 7 1 2 70157 19701
0 19703 5 1 1 19702
0 19704 7 1 2 73712 78443
0 19705 5 1 1 19704
0 19706 7 3 2 65387 73011
0 19707 7 1 2 67962 91783
0 19708 5 1 1 19707
0 19709 7 1 2 19705 19708
0 19710 5 1 1 19709
0 19711 7 1 2 90077 19710
0 19712 5 1 1 19711
0 19713 7 1 2 68318 19712
0 19714 7 1 2 19703 19713
0 19715 7 1 2 19671 19714
0 19716 5 1 1 19715
0 19717 7 2 2 66469 82903
0 19718 5 2 1 91786
0 19719 7 1 2 65189 91787
0 19720 5 1 1 19719
0 19721 7 1 2 90790 19720
0 19722 5 1 1 19721
0 19723 7 1 2 14477 19722
0 19724 5 1 1 19723
0 19725 7 1 2 83934 19724
0 19726 5 1 1 19725
0 19727 7 2 2 69545 76555
0 19728 5 2 1 91790
0 19729 7 1 2 62963 91792
0 19730 5 4 1 19729
0 19731 7 1 2 68646 91107
0 19732 7 1 2 91794 19731
0 19733 5 1 1 19732
0 19734 7 1 2 19726 19733
0 19735 5 1 1 19734
0 19736 7 1 2 67289 19735
0 19737 5 1 1 19736
0 19738 7 1 2 62964 13487
0 19739 5 2 1 19738
0 19740 7 1 2 63707 91798
0 19741 7 1 2 91515 19740
0 19742 5 1 1 19741
0 19743 7 1 2 19737 19742
0 19744 5 1 1 19743
0 19745 7 1 2 61692 19744
0 19746 5 1 1 19745
0 19747 7 2 2 66672 87890
0 19748 5 1 1 91800
0 19749 7 1 2 83661 84827
0 19750 5 2 1 19749
0 19751 7 1 2 69546 84335
0 19752 5 2 1 19751
0 19753 7 1 2 91802 91804
0 19754 5 1 1 19753
0 19755 7 1 2 77115 19754
0 19756 5 1 1 19755
0 19757 7 1 2 19748 19756
0 19758 5 1 1 19757
0 19759 7 1 2 71394 85084
0 19760 7 1 2 19758 19759
0 19761 5 1 1 19760
0 19762 7 1 2 19746 19761
0 19763 5 1 1 19762
0 19764 7 1 2 60496 19763
0 19765 5 1 1 19764
0 19766 7 1 2 69547 83978
0 19767 5 1 1 19766
0 19768 7 1 2 91803 19767
0 19769 5 1 1 19768
0 19770 7 1 2 76556 19769
0 19771 5 1 1 19770
0 19772 7 1 2 8797 19771
0 19773 5 1 1 19772
0 19774 7 1 2 71359 91523
0 19775 7 1 2 19773 19774
0 19776 5 1 1 19775
0 19777 7 1 2 63411 19776
0 19778 7 1 2 19765 19777
0 19779 5 1 1 19778
0 19780 7 1 2 72100 19779
0 19781 7 1 2 19716 19780
0 19782 5 1 1 19781
0 19783 7 12 2 63708 89312
0 19784 5 1 1 91806
0 19785 7 1 2 59504 91807
0 19786 5 1 1 19785
0 19787 7 1 2 80180 84310
0 19788 5 1 1 19787
0 19789 7 1 2 19786 19788
0 19790 5 1 1 19789
0 19791 7 1 2 76341 19790
0 19792 5 1 1 19791
0 19793 7 1 2 84336 91622
0 19794 5 1 1 19793
0 19795 7 17 2 63709 79646
0 19796 5 3 1 91818
0 19797 7 1 2 62628 76978
0 19798 5 2 1 19797
0 19799 7 1 2 91819 91838
0 19800 5 1 1 19799
0 19801 7 1 2 19794 19800
0 19802 5 1 1 19801
0 19803 7 1 2 75489 19802
0 19804 5 1 1 19803
0 19805 7 1 2 83150 91839
0 19806 5 1 1 19805
0 19807 7 1 2 19804 19806
0 19808 5 1 1 19807
0 19809 7 1 2 69548 19808
0 19810 5 1 1 19809
0 19811 7 1 2 19792 19810
0 19812 5 1 1 19811
0 19813 7 1 2 70601 19812
0 19814 5 1 1 19813
0 19815 7 2 2 69549 82077
0 19816 5 1 1 91840
0 19817 7 10 2 60497 75281
0 19818 5 32 1 91842
0 19819 7 1 2 84475 91843
0 19820 7 1 2 91841 19819
0 19821 5 1 1 19820
0 19822 7 1 2 19814 19821
0 19823 5 1 1 19822
0 19824 7 1 2 77772 19823
0 19825 5 1 1 19824
0 19826 7 1 2 61693 69464
0 19827 7 1 2 84214 19826
0 19828 5 1 1 19827
0 19829 7 7 2 66673 67053
0 19830 7 7 2 67290 68647
0 19831 5 1 1 91891
0 19832 7 2 2 81337 91892
0 19833 7 1 2 91884 91898
0 19834 5 1 1 19833
0 19835 7 1 2 69107 76180
0 19836 7 1 2 91820 19835
0 19837 5 1 1 19836
0 19838 7 1 2 19834 19837
0 19839 5 1 1 19838
0 19840 7 1 2 79824 83425
0 19841 7 1 2 19839 19840
0 19842 5 1 1 19841
0 19843 7 1 2 19828 19842
0 19844 5 1 1 19843
0 19845 7 1 2 60322 19844
0 19846 5 1 1 19845
0 19847 7 1 2 69108 91500
0 19848 5 1 1 19847
0 19849 7 1 2 14757 19848
0 19850 5 1 1 19849
0 19851 7 1 2 85152 19850
0 19852 5 1 1 19851
0 19853 7 1 2 19846 19852
0 19854 5 1 1 19853
0 19855 7 1 2 59505 19854
0 19856 5 1 1 19855
0 19857 7 1 2 79256 91755
0 19858 7 1 2 78479 19857
0 19859 5 1 1 19858
0 19860 7 1 2 81938 78329
0 19861 7 1 2 89313 19860
0 19862 5 1 1 19861
0 19863 7 1 2 19859 19862
0 19864 5 1 1 19863
0 19865 7 1 2 78749 19864
0 19866 5 1 1 19865
0 19867 7 1 2 19856 19866
0 19868 5 1 1 19867
0 19869 7 1 2 70158 19868
0 19870 5 1 1 19869
0 19871 7 1 2 70602 89314
0 19872 5 1 1 19871
0 19873 7 1 2 19872 89455
0 19874 5 3 1 19873
0 19875 7 3 2 63710 80729
0 19876 7 1 2 62629 91903
0 19877 7 1 2 91900 19876
0 19878 5 1 1 19877
0 19879 7 1 2 80861 83577
0 19880 5 1 1 19879
0 19881 7 1 2 19878 19880
0 19882 7 1 2 19870 19881
0 19883 5 1 1 19882
0 19884 7 1 2 67963 19883
0 19885 5 1 1 19884
0 19886 7 1 2 19825 19885
0 19887 5 1 1 19886
0 19888 7 1 2 71198 19887
0 19889 5 1 1 19888
0 19890 7 1 2 90017 91630
0 19891 5 1 1 19890
0 19892 7 1 2 91808 19891
0 19893 5 1 1 19892
0 19894 7 1 2 84389 91631
0 19895 5 1 1 19894
0 19896 7 3 2 66674 73012
0 19897 5 1 1 91906
0 19898 7 1 2 87950 91907
0 19899 7 1 2 19895 19898
0 19900 5 1 1 19899
0 19901 7 1 2 19893 19900
0 19902 5 1 1 19901
0 19903 7 1 2 61311 19902
0 19904 5 1 1 19903
0 19905 7 3 2 84426 86452
0 19906 5 1 1 91909
0 19907 7 1 2 71712 85445
0 19908 7 1 2 91910 19907
0 19909 5 1 1 19908
0 19910 7 1 2 19904 19909
0 19911 5 1 1 19910
0 19912 7 1 2 69550 19911
0 19913 5 1 1 19912
0 19914 7 2 2 66470 78370
0 19915 5 1 1 91912
0 19916 7 1 2 67595 79980
0 19917 5 1 1 19916
0 19918 7 1 2 66253 19917
0 19919 5 1 1 19918
0 19920 7 1 2 91913 19919
0 19921 5 1 1 19920
0 19922 7 1 2 62965 89484
0 19923 5 1 1 19922
0 19924 7 1 2 19921 19923
0 19925 5 1 1 19924
0 19926 7 1 2 83151 19925
0 19927 5 1 1 19926
0 19928 7 1 2 19913 19927
0 19929 5 1 1 19928
0 19930 7 1 2 68319 19929
0 19931 5 1 1 19930
0 19932 7 2 2 66471 79360
0 19933 7 1 2 78017 91914
0 19934 7 5 2 67964 83527
0 19935 5 1 1 91916
0 19936 7 1 2 91917 88888
0 19937 7 1 2 19933 19936
0 19938 5 1 1 19937
0 19939 7 1 2 19931 19938
0 19940 5 1 1 19939
0 19941 7 1 2 72920 19940
0 19942 5 1 1 19941
0 19943 7 1 2 63946 19942
0 19944 7 1 2 19889 19943
0 19945 7 1 2 19782 19944
0 19946 7 1 2 19619 19945
0 19947 7 1 2 19244 19946
0 19948 5 1 1 19947
0 19949 7 1 2 86744 19948
0 19950 7 1 2 18428 19949
0 19951 5 1 1 19950
0 19952 7 3 2 68320 70527
0 19953 7 1 2 85129 91921
0 19954 5 1 1 19953
0 19955 7 1 2 79884 89983
0 19956 5 1 1 19955
0 19957 7 1 2 19954 19956
0 19958 5 1 1 19957
0 19959 7 1 2 88889 19958
0 19960 5 1 1 19959
0 19961 7 1 2 84179 85902
0 19962 5 1 1 19961
0 19963 7 1 2 19960 19962
0 19964 5 1 1 19963
0 19965 7 1 2 59855 19964
0 19966 5 1 1 19965
0 19967 7 2 2 67291 89923
0 19968 7 1 2 65388 80761
0 19969 7 1 2 91924 19968
0 19970 5 1 1 19969
0 19971 7 1 2 19966 19970
0 19972 5 1 1 19971
0 19973 7 1 2 67965 19972
0 19974 5 1 1 19973
0 19975 7 1 2 82552 90598
0 19976 5 1 1 19975
0 19977 7 4 2 68321 83900
0 19978 7 1 2 61312 91926
0 19979 5 1 1 19978
0 19980 7 1 2 19976 19979
0 19981 5 1 1 19980
0 19982 7 1 2 89997 19981
0 19983 5 1 1 19982
0 19984 7 1 2 19974 19983
0 19985 5 1 1 19984
0 19986 7 1 2 67596 19985
0 19987 5 1 1 19986
0 19988 7 2 2 74966 76557
0 19989 7 1 2 79010 85903
0 19990 7 1 2 91930 19989
0 19991 5 1 1 19990
0 19992 7 1 2 19987 19991
0 19993 5 1 1 19992
0 19994 7 1 2 72948 19993
0 19995 5 1 1 19994
0 19996 7 2 2 72101 72921
0 19997 5 2 1 91932
0 19998 7 1 2 84818 91403
0 19999 7 1 2 91933 19998
0 20000 5 1 1 19999
0 20001 7 1 2 19995 20000
0 20002 5 1 1 20001
0 20003 7 1 2 81092 20002
0 20004 5 1 1 20003
0 20005 7 1 2 71007 88594
0 20006 5 1 1 20005
0 20007 7 1 2 73686 75065
0 20008 5 1 1 20007
0 20009 7 1 2 20006 20008
0 20010 5 1 1 20009
0 20011 7 1 2 66472 20010
0 20012 5 1 1 20011
0 20013 7 1 2 62094 90680
0 20014 5 1 1 20013
0 20015 7 1 2 20012 20014
0 20016 5 1 1 20015
0 20017 7 1 2 68648 20016
0 20018 5 1 1 20017
0 20019 7 1 2 75282 73502
0 20020 5 1 1 20019
0 20021 7 2 2 75459 20020
0 20022 5 2 1 91936
0 20023 7 2 2 71713 91938
0 20024 5 1 1 91940
0 20025 7 1 2 89988 91941
0 20026 5 1 1 20025
0 20027 7 1 2 20018 20026
0 20028 5 1 1 20027
0 20029 7 1 2 62630 20028
0 20030 5 1 1 20029
0 20031 7 6 2 63711 85904
0 20032 5 1 1 91942
0 20033 7 1 2 78459 91943
0 20034 5 1 1 20033
0 20035 7 1 2 15120 20034
0 20036 5 1 1 20035
0 20037 7 4 2 67597 72922
0 20038 7 1 2 66254 91948
0 20039 7 1 2 20036 20038
0 20040 5 1 1 20039
0 20041 7 1 2 20030 20040
0 20042 5 1 1 20041
0 20043 7 1 2 62966 20042
0 20044 5 1 1 20043
0 20045 7 1 2 60908 78251
0 20046 5 2 1 20045
0 20047 7 1 2 75720 78295
0 20048 5 1 1 20047
0 20049 7 1 2 59506 20048
0 20050 5 1 1 20049
0 20051 7 1 2 61313 76342
0 20052 5 1 1 20051
0 20053 7 1 2 84610 20052
0 20054 7 1 2 20050 20053
0 20055 5 1 1 20054
0 20056 7 1 2 67292 20055
0 20057 5 1 1 20056
0 20058 7 1 2 91952 20057
0 20059 5 1 1 20058
0 20060 7 1 2 61502 20059
0 20061 5 1 1 20060
0 20062 7 1 2 76325 82084
0 20063 5 1 1 20062
0 20064 7 1 2 83053 72949
0 20065 7 1 2 20063 20064
0 20066 5 1 1 20065
0 20067 7 1 2 20061 20066
0 20068 5 1 1 20067
0 20069 7 1 2 60323 20068
0 20070 5 1 1 20069
0 20071 7 3 2 60117 69179
0 20072 5 2 1 91954
0 20073 7 1 2 74967 84597
0 20074 5 1 1 20073
0 20075 7 1 2 91957 20074
0 20076 5 1 1 20075
0 20077 7 3 2 67598 74944
0 20078 5 1 1 91959
0 20079 7 1 2 75721 83067
0 20080 5 2 1 20079
0 20081 7 1 2 91960 91962
0 20082 7 1 2 20076 20081
0 20083 5 1 1 20082
0 20084 7 1 2 20070 20083
0 20085 5 1 1 20084
0 20086 7 1 2 63412 20085
0 20087 5 1 1 20086
0 20088 7 1 2 75047 77900
0 20089 7 1 2 82755 20088
0 20090 5 1 1 20089
0 20091 7 1 2 60324 81202
0 20092 5 1 1 20091
0 20093 7 1 2 20090 20092
0 20094 5 1 1 20093
0 20095 7 1 2 60909 20094
0 20096 5 1 1 20095
0 20097 7 1 2 59507 89112
0 20098 5 1 1 20097
0 20099 7 1 2 68322 74553
0 20100 5 1 1 20099
0 20101 7 1 2 20098 20100
0 20102 5 1 1 20101
0 20103 7 1 2 86965 20102
0 20104 5 1 1 20103
0 20105 7 1 2 20096 20104
0 20106 5 1 1 20105
0 20107 7 1 2 72923 20106
0 20108 5 1 1 20107
0 20109 7 2 2 74364 85768
0 20110 5 1 1 91964
0 20111 7 1 2 78354 91965
0 20112 5 1 1 20111
0 20113 7 1 2 75732 91963
0 20114 5 1 1 20113
0 20115 7 1 2 79947 89676
0 20116 5 1 1 20115
0 20117 7 1 2 20114 20116
0 20118 5 1 1 20117
0 20119 7 1 2 72979 20118
0 20120 5 1 1 20119
0 20121 7 1 2 20112 20120
0 20122 7 1 2 20108 20121
0 20123 7 1 2 20087 20122
0 20124 5 1 1 20123
0 20125 7 1 2 63712 20124
0 20126 5 1 1 20125
0 20127 7 2 2 62631 79557
0 20128 7 1 2 90828 91966
0 20129 5 1 1 20128
0 20130 7 1 2 82025 20129
0 20131 5 1 1 20130
0 20132 7 1 2 91918 20131
0 20133 5 1 1 20132
0 20134 7 1 2 20126 20133
0 20135 7 1 2 20044 20134
0 20136 5 1 1 20135
0 20137 7 1 2 65389 20136
0 20138 5 1 1 20137
0 20139 7 1 2 75436 85579
0 20140 7 1 2 81241 20139
0 20141 7 1 2 89848 20140
0 20142 5 1 1 20141
0 20143 7 1 2 20138 20142
0 20144 5 1 1 20143
0 20145 7 1 2 68856 20144
0 20146 5 1 1 20145
0 20147 7 1 2 20004 20146
0 20148 5 1 1 20147
0 20149 7 1 2 66675 20148
0 20150 5 1 1 20149
0 20151 7 2 2 74991 83594
0 20152 5 1 1 91968
0 20153 7 2 2 68323 89357
0 20154 5 1 1 91970
0 20155 7 1 2 59508 91971
0 20156 5 1 1 20155
0 20157 7 1 2 20152 20156
0 20158 5 1 1 20157
0 20159 7 1 2 66676 20158
0 20160 5 1 1 20159
0 20161 7 1 2 3997 20160
0 20162 5 1 1 20161
0 20163 7 1 2 67054 20162
0 20164 5 1 1 20163
0 20165 7 1 2 74404 85635
0 20166 5 1 1 20165
0 20167 7 1 2 20164 20166
0 20168 5 1 1 20167
0 20169 7 1 2 63713 20168
0 20170 5 1 1 20169
0 20171 7 1 2 78333 84863
0 20172 7 1 2 85336 20171
0 20173 5 1 1 20172
0 20174 7 1 2 20170 20173
0 20175 5 1 1 20174
0 20176 7 1 2 67966 20175
0 20177 5 1 1 20176
0 20178 7 1 2 67599 78750
0 20179 7 1 2 84618 85593
0 20180 7 1 2 20178 20179
0 20181 7 1 2 81600 20180
0 20182 5 1 1 20181
0 20183 7 1 2 20177 20182
0 20184 5 1 1 20183
0 20185 7 1 2 68857 20184
0 20186 5 1 1 20185
0 20187 7 1 2 71405 73961
0 20188 5 1 1 20187
0 20189 7 2 2 81534 74365
0 20190 5 1 1 91972
0 20191 7 1 2 20188 20190
0 20192 5 1 1 20191
0 20193 7 1 2 73474 90193
0 20194 7 1 2 20192 20193
0 20195 5 1 1 20194
0 20196 7 1 2 20186 20195
0 20197 5 1 1 20196
0 20198 7 1 2 65390 20197
0 20199 5 1 1 20198
0 20200 7 1 2 84180 72805
0 20201 5 1 1 20200
0 20202 7 3 2 60910 63714
0 20203 7 2 2 59509 73687
0 20204 7 1 2 91974 91977
0 20205 7 1 2 90634 20204
0 20206 5 1 1 20205
0 20207 7 1 2 20201 20206
0 20208 5 1 1 20207
0 20209 7 1 2 80025 20208
0 20210 5 1 1 20209
0 20211 7 2 2 81338 75010
0 20212 7 1 2 73770 89971
0 20213 7 1 2 91979 20212
0 20214 5 1 1 20213
0 20215 7 1 2 20210 20214
0 20216 5 1 1 20215
0 20217 7 1 2 68858 20216
0 20218 5 1 1 20217
0 20219 7 5 2 70603 91665
0 20220 5 1 1 91981
0 20221 7 1 2 91852 20220
0 20222 5 4 1 20221
0 20223 7 2 2 69180 81012
0 20224 7 1 2 68649 91990
0 20225 7 1 2 91986 20224
0 20226 5 1 1 20225
0 20227 7 1 2 20218 20226
0 20228 5 1 1 20227
0 20229 7 1 2 66677 20228
0 20230 5 1 1 20229
0 20231 7 1 2 83581 91987
0 20232 5 1 1 20231
0 20233 7 1 2 90765 91899
0 20234 5 1 1 20233
0 20235 7 1 2 20232 20234
0 20236 5 1 1 20235
0 20237 7 1 2 81013 20236
0 20238 5 1 1 20237
0 20239 7 9 2 66473 85509
0 20240 7 2 2 84736 91992
0 20241 7 1 2 91980 92001
0 20242 5 1 1 20241
0 20243 7 1 2 20238 20242
0 20244 5 1 1 20243
0 20245 7 1 2 61694 20244
0 20246 5 1 1 20245
0 20247 7 7 2 61314 89637
0 20248 7 1 2 83582 92003
0 20249 7 1 2 89249 20248
0 20250 5 1 1 20249
0 20251 7 1 2 20246 20250
0 20252 7 1 2 20230 20251
0 20253 5 1 1 20252
0 20254 7 1 2 67600 20253
0 20255 5 1 1 20254
0 20256 7 6 2 68650 80406
0 20257 5 1 1 92010
0 20258 7 1 2 75011 92011
0 20259 5 1 1 20258
0 20260 7 1 2 6273 20259
0 20261 5 1 1 20260
0 20262 7 1 2 90766 20261
0 20263 5 1 1 20262
0 20264 7 1 2 75012 84337
0 20265 5 2 1 20264
0 20266 7 1 2 91835 92016
0 20267 5 1 1 20266
0 20268 7 1 2 90065 20267
0 20269 5 1 1 20268
0 20270 7 1 2 20263 20269
0 20271 5 1 1 20270
0 20272 7 1 2 91991 20271
0 20273 5 1 1 20272
0 20274 7 1 2 20255 20273
0 20275 5 1 1 20274
0 20276 7 1 2 62967 20275
0 20277 5 1 1 20276
0 20278 7 5 2 75283 80679
0 20279 5 1 1 92018
0 20280 7 1 2 62968 92019
0 20281 5 1 1 20280
0 20282 7 7 2 63947 89315
0 20283 7 1 2 76343 78869
0 20284 7 1 2 92023 20283
0 20285 5 1 1 20284
0 20286 7 1 2 20281 20285
0 20287 5 1 1 20286
0 20288 7 1 2 73590 20287
0 20289 5 1 1 20288
0 20290 7 4 2 60498 79257
0 20291 7 5 2 67601 73475
0 20292 7 2 2 92030 92034
0 20293 5 1 1 92039
0 20294 7 1 2 70528 92040
0 20295 5 1 1 20294
0 20296 7 1 2 20289 20295
0 20297 5 1 1 20296
0 20298 7 1 2 68324 20297
0 20299 5 1 1 20298
0 20300 7 6 2 68325 78252
0 20301 5 1 1 92041
0 20302 7 3 2 61503 63948
0 20303 7 2 2 92047 89011
0 20304 7 1 2 92042 92050
0 20305 5 1 1 20304
0 20306 7 5 2 62969 80536
0 20307 7 2 2 62632 86662
0 20308 7 1 2 92052 92057
0 20309 5 1 1 20308
0 20310 7 1 2 20305 20309
0 20311 5 1 1 20310
0 20312 7 1 2 81172 20311
0 20313 5 1 1 20312
0 20314 7 1 2 20299 20313
0 20315 5 1 1 20314
0 20316 7 1 2 63715 20315
0 20317 5 1 1 20316
0 20318 7 1 2 86131 88116
0 20319 7 1 2 91192 20318
0 20320 7 1 2 89917 20319
0 20321 5 1 1 20320
0 20322 7 1 2 20317 20321
0 20323 5 1 1 20322
0 20324 7 1 2 70159 20323
0 20325 5 1 1 20324
0 20326 7 5 2 67293 63716
0 20327 7 1 2 82626 92031
0 20328 5 1 1 20327
0 20329 7 1 2 67602 80548
0 20330 7 1 2 85655 20329
0 20331 5 1 1 20330
0 20332 7 1 2 20328 20331
0 20333 5 1 1 20332
0 20334 7 1 2 60118 20333
0 20335 5 1 1 20334
0 20336 7 2 2 60499 74342
0 20337 7 2 2 81014 88083
0 20338 7 1 2 92064 92066
0 20339 5 1 1 20338
0 20340 7 1 2 20335 20339
0 20341 5 1 1 20340
0 20342 7 1 2 92059 20341
0 20343 5 1 1 20342
0 20344 7 1 2 78399 89972
0 20345 5 1 1 20344
0 20346 7 2 2 73948 87891
0 20347 5 1 1 92068
0 20348 7 1 2 20345 20347
0 20349 5 1 1 20348
0 20350 7 1 2 60325 20349
0 20351 5 1 1 20350
0 20352 7 1 2 61504 92069
0 20353 5 1 1 20352
0 20354 7 1 2 20351 20353
0 20355 5 1 1 20354
0 20356 7 1 2 73476 20355
0 20357 5 1 1 20356
0 20358 7 2 2 85866 87565
0 20359 5 1 1 92070
0 20360 7 1 2 66255 92071
0 20361 5 1 1 20360
0 20362 7 1 2 20357 20361
0 20363 5 1 1 20362
0 20364 7 1 2 81173 20363
0 20365 5 1 1 20364
0 20366 7 1 2 20343 20365
0 20367 5 1 1 20366
0 20368 7 1 2 67055 20367
0 20369 5 1 1 20368
0 20370 7 2 2 66474 79286
0 20371 7 2 2 81766 92072
0 20372 7 1 2 81307 83528
0 20373 7 1 2 92074 20372
0 20374 5 1 1 20373
0 20375 7 1 2 20369 20374
0 20376 5 1 1 20375
0 20377 7 1 2 72102 20376
0 20378 5 1 1 20377
0 20379 7 2 2 77547 85905
0 20380 5 5 1 92076
0 20381 7 1 2 91993 89459
0 20382 5 1 1 20381
0 20383 7 1 2 92078 20382
0 20384 5 1 1 20383
0 20385 7 2 2 66678 81077
0 20386 7 1 2 77425 92083
0 20387 7 1 2 20384 20386
0 20388 5 1 1 20387
0 20389 7 1 2 20378 20388
0 20390 7 1 2 20325 20389
0 20391 7 1 2 20277 20390
0 20392 7 1 2 20199 20391
0 20393 5 1 1 20392
0 20394 7 1 2 71199 20393
0 20395 5 1 1 20394
0 20396 7 2 2 77373 88616
0 20397 5 1 1 92085
0 20398 7 1 2 69181 78188
0 20399 5 3 1 20398
0 20400 7 1 2 83042 92087
0 20401 5 2 1 20400
0 20402 7 1 2 80226 70896
0 20403 7 1 2 92090 20402
0 20404 5 1 1 20403
0 20405 7 1 2 20397 20404
0 20406 5 1 1 20405
0 20407 7 1 2 68326 20406
0 20408 5 1 1 20407
0 20409 7 1 2 82339 74940
0 20410 5 1 1 20409
0 20411 7 1 2 20408 20410
0 20412 5 1 1 20411
0 20413 7 7 2 75490 85130
0 20414 5 1 1 92092
0 20415 7 1 2 20412 92093
0 20416 5 1 1 20415
0 20417 7 1 2 69465 89652
0 20418 5 1 1 20417
0 20419 7 1 2 81078 83300
0 20420 5 1 1 20419
0 20421 7 1 2 20418 20420
0 20422 5 1 1 20421
0 20423 7 1 2 83529 20422
0 20424 5 1 1 20423
0 20425 7 1 2 74732 88597
0 20426 5 1 1 20425
0 20427 7 1 2 17866 20426
0 20428 5 1 1 20427
0 20429 7 1 2 90635 20428
0 20430 5 1 1 20429
0 20431 7 2 2 62633 76771
0 20432 5 1 1 92099
0 20433 7 1 2 90628 92100
0 20434 5 1 1 20433
0 20435 7 1 2 91666 91782
0 20436 5 1 1 20435
0 20437 7 5 2 59510 60500
0 20438 5 1 1 92101
0 20439 7 2 2 60911 92102
0 20440 7 1 2 74733 92106
0 20441 5 1 1 20440
0 20442 7 1 2 20436 20441
0 20443 5 1 1 20442
0 20444 7 1 2 70160 20443
0 20445 5 1 1 20444
0 20446 7 1 2 20434 20445
0 20447 7 1 2 20430 20446
0 20448 5 1 1 20447
0 20449 7 1 2 78751 20448
0 20450 5 1 1 20449
0 20451 7 1 2 20424 20450
0 20452 5 1 1 20451
0 20453 7 1 2 67967 20452
0 20454 5 1 1 20453
0 20455 7 3 2 60912 77773
0 20456 5 2 1 92108
0 20457 7 2 2 63413 74589
0 20458 7 1 2 72950 92113
0 20459 5 1 1 20458
0 20460 7 1 2 92111 20459
0 20461 5 1 1 20460
0 20462 7 1 2 91844 20461
0 20463 5 1 1 20462
0 20464 7 1 2 68327 89720
0 20465 7 1 2 91667 20464
0 20466 7 1 2 70910 20465
0 20467 5 1 1 20466
0 20468 7 1 2 20463 20467
0 20469 5 1 1 20468
0 20470 7 1 2 67603 20469
0 20471 5 1 1 20470
0 20472 7 15 2 60501 75491
0 20473 5 3 1 92115
0 20474 7 1 2 92114 92116
0 20475 5 1 1 20474
0 20476 7 1 2 20471 20475
0 20477 5 1 1 20476
0 20478 7 1 2 67294 20477
0 20479 5 1 1 20478
0 20480 7 1 2 60502 81872
0 20481 7 1 2 91516 20480
0 20482 5 1 1 20481
0 20483 7 1 2 20479 20482
0 20484 5 1 1 20483
0 20485 7 1 2 63717 20484
0 20486 5 1 1 20485
0 20487 7 1 2 20454 20486
0 20488 5 1 1 20487
0 20489 7 1 2 67056 20488
0 20490 5 1 1 20489
0 20491 7 1 2 73949 90154
0 20492 5 3 1 20491
0 20493 7 1 2 77806 92133
0 20494 5 1 1 20493
0 20495 7 1 2 91668 20494
0 20496 5 1 1 20495
0 20497 7 4 2 80950 78371
0 20498 7 1 2 71714 75877
0 20499 7 1 2 92136 20498
0 20500 5 1 1 20499
0 20501 7 1 2 20496 20500
0 20502 5 1 1 20501
0 20503 7 1 2 83662 20502
0 20504 5 1 1 20503
0 20505 7 1 2 59511 92091
0 20506 5 1 1 20505
0 20507 7 1 2 78330 78870
0 20508 5 4 1 20507
0 20509 7 1 2 20506 92140
0 20510 5 1 1 20509
0 20511 7 1 2 83402 89766
0 20512 7 1 2 20510 20511
0 20513 5 1 1 20512
0 20514 7 1 2 20504 20513
0 20515 5 1 1 20514
0 20516 7 1 2 60119 20515
0 20517 5 1 1 20516
0 20518 7 3 2 63718 77774
0 20519 7 1 2 91845 92144
0 20520 5 1 1 20519
0 20521 7 6 2 62634 83530
0 20522 5 1 1 92147
0 20523 7 1 2 86955 92148
0 20524 5 1 1 20523
0 20525 7 5 2 60503 78752
0 20526 5 1 1 92153
0 20527 7 1 2 82231 92154
0 20528 5 1 1 20527
0 20529 7 1 2 20524 20528
0 20530 5 1 1 20529
0 20531 7 1 2 59512 20530
0 20532 5 1 1 20531
0 20533 7 1 2 60326 76480
0 20534 7 1 2 75684 87892
0 20535 7 1 2 20533 20534
0 20536 5 1 1 20535
0 20537 7 1 2 20532 20536
0 20538 5 1 1 20537
0 20539 7 1 2 82405 20538
0 20540 5 1 1 20539
0 20541 7 1 2 20520 20540
0 20542 7 1 2 20517 20541
0 20543 5 1 1 20542
0 20544 7 1 2 61045 20543
0 20545 5 1 1 20544
0 20546 7 6 2 67968 75284
0 20547 7 1 2 83663 92158
0 20548 5 2 1 20547
0 20549 7 1 2 59513 83979
0 20550 5 1 1 20549
0 20551 7 1 2 92164 20550
0 20552 5 1 1 20551
0 20553 7 4 2 60504 60913
0 20554 7 1 2 80111 92166
0 20555 7 1 2 20552 20554
0 20556 5 1 1 20555
0 20557 7 1 2 20545 20556
0 20558 5 1 1 20557
0 20559 7 1 2 59856 20558
0 20560 5 1 1 20559
0 20561 7 2 2 67969 76673
0 20562 5 7 1 92170
0 20563 7 2 2 59514 92172
0 20564 7 1 2 78592 92179
0 20565 5 1 1 20564
0 20566 7 1 2 92141 20565
0 20567 5 1 1 20566
0 20568 7 1 2 60505 20567
0 20569 5 1 1 20568
0 20570 7 1 2 88947 92180
0 20571 5 1 1 20570
0 20572 7 1 2 92142 20571
0 20573 5 1 1 20572
0 20574 7 1 2 81347 20573
0 20575 5 1 1 20574
0 20576 7 1 2 20569 20575
0 20577 5 1 1 20576
0 20578 7 1 2 84864 20577
0 20579 5 1 1 20578
0 20580 7 4 2 59515 74916
0 20581 7 1 2 91069 92181
0 20582 5 1 1 20581
0 20583 7 1 2 90040 20582
0 20584 5 1 1 20583
0 20585 7 3 2 60506 70161
0 20586 7 1 2 78753 92185
0 20587 7 1 2 20584 20586
0 20588 5 1 1 20587
0 20589 7 1 2 20579 20588
0 20590 7 1 2 20560 20589
0 20591 7 1 2 20490 20590
0 20592 5 1 1 20591
0 20593 7 1 2 61695 20592
0 20594 5 1 1 20593
0 20595 7 1 2 20416 20594
0 20596 5 1 1 20595
0 20597 7 1 2 63949 20596
0 20598 5 1 1 20597
0 20599 7 1 2 63719 81473
0 20600 7 1 2 91644 20599
0 20601 5 1 1 20600
0 20602 7 1 2 68651 69306
0 20603 7 1 2 91573 20602
0 20604 5 1 1 20603
0 20605 7 1 2 20601 20604
0 20606 5 1 1 20605
0 20607 7 1 2 61505 20606
0 20608 5 1 1 20607
0 20609 7 1 2 76996 89767
0 20610 7 1 2 90797 20609
0 20611 5 1 1 20610
0 20612 7 1 2 20608 20611
0 20613 5 1 1 20612
0 20614 7 1 2 81015 20613
0 20615 5 1 1 20614
0 20616 7 2 2 73165 87940
0 20617 7 1 2 70529 92188
0 20618 5 1 1 20617
0 20619 7 1 2 75201 90794
0 20620 5 2 1 20619
0 20621 7 4 2 67057 77548
0 20622 7 2 2 61315 77116
0 20623 7 1 2 92192 92196
0 20624 7 1 2 92190 20623
0 20625 5 1 1 20624
0 20626 7 1 2 20618 20625
0 20627 5 1 1 20626
0 20628 7 1 2 71715 20627
0 20629 5 1 1 20628
0 20630 7 1 2 62300 79558
0 20631 7 1 2 87702 20630
0 20632 5 1 1 20631
0 20633 7 1 2 74680 77549
0 20634 7 1 2 72924 20633
0 20635 5 1 1 20634
0 20636 7 1 2 20632 20635
0 20637 5 1 1 20636
0 20638 7 1 2 72103 20637
0 20639 5 1 1 20638
0 20640 7 2 2 65190 83301
0 20641 7 1 2 87703 92198
0 20642 5 2 1 20641
0 20643 7 1 2 20639 92200
0 20644 7 1 2 20629 20643
0 20645 5 1 1 20644
0 20646 7 1 2 63414 20645
0 20647 5 1 1 20646
0 20648 7 1 2 20615 20647
0 20649 5 1 1 20648
0 20650 7 1 2 67970 20649
0 20651 5 1 1 20650
0 20652 7 3 2 75285 90107
0 20653 5 1 1 92202
0 20654 7 1 2 75048 92203
0 20655 5 1 1 20654
0 20656 7 2 2 68859 79035
0 20657 7 1 2 86663 92205
0 20658 7 1 2 81242 20657
0 20659 5 1 1 20658
0 20660 7 1 2 20655 20659
0 20661 5 1 1 20660
0 20662 7 1 2 73503 20661
0 20663 5 1 1 20662
0 20664 7 2 2 61046 75049
0 20665 5 2 1 92207
0 20666 7 5 2 61316 73408
0 20667 7 1 2 86466 92211
0 20668 7 1 2 92208 20667
0 20669 5 1 1 20668
0 20670 7 1 2 20663 20669
0 20671 5 1 1 20670
0 20672 7 1 2 62970 20671
0 20673 5 1 1 20672
0 20674 7 2 2 71716 75724
0 20675 7 1 2 67295 86492
0 20676 7 1 2 92216 20675
0 20677 7 1 2 90798 20676
0 20678 5 1 1 20677
0 20679 7 1 2 20673 20678
0 20680 7 1 2 20651 20679
0 20681 5 1 1 20680
0 20682 7 1 2 81174 20681
0 20683 5 1 1 20682
0 20684 7 1 2 20598 20683
0 20685 7 1 2 20395 20684
0 20686 7 1 2 20150 20685
0 20687 5 1 1 20686
0 20688 7 1 2 86745 20687
0 20689 5 1 1 20688
0 20690 7 2 2 67604 88625
0 20691 5 2 1 92218
0 20692 7 1 2 88916 92220
0 20693 5 1 1 20692
0 20694 7 2 2 60120 20693
0 20695 5 1 1 92222
0 20696 7 1 2 89493 20695
0 20697 5 1 1 20696
0 20698 7 1 2 82171 20697
0 20699 5 1 1 20698
0 20700 7 1 2 65391 90801
0 20701 5 1 1 20700
0 20702 7 1 2 80026 20701
0 20703 5 1 1 20702
0 20704 7 1 2 20699 20703
0 20705 5 1 1 20704
0 20706 7 1 2 68652 20705
0 20707 5 1 1 20706
0 20708 7 6 2 63720 91669
0 20709 7 1 2 80782 88626
0 20710 7 1 2 92224 20709
0 20711 5 1 1 20710
0 20712 7 1 2 20707 20711
0 20713 5 1 1 20712
0 20714 7 1 2 61317 20713
0 20715 5 1 1 20714
0 20716 7 1 2 60121 82651
0 20717 7 1 2 92225 20716
0 20718 5 1 1 20717
0 20719 7 5 2 68653 75286
0 20720 5 1 1 92230
0 20721 7 1 2 65392 92231
0 20722 5 1 1 20721
0 20723 7 1 2 20718 20722
0 20724 5 1 1 20723
0 20725 7 1 2 59857 20724
0 20726 5 1 1 20725
0 20727 7 1 2 60507 83583
0 20728 5 2 1 20727
0 20729 7 1 2 68654 91394
0 20730 5 1 1 20729
0 20731 7 1 2 92235 20730
0 20732 5 1 1 20731
0 20733 7 1 2 75287 20732
0 20734 5 1 1 20733
0 20735 7 1 2 20726 20734
0 20736 5 1 1 20735
0 20737 7 1 2 67605 20736
0 20738 5 1 1 20737
0 20739 7 2 2 75288 85131
0 20740 7 1 2 71200 92237
0 20741 5 1 1 20740
0 20742 7 1 2 20738 20741
0 20743 5 1 1 20742
0 20744 7 1 2 83185 20743
0 20745 5 1 1 20744
0 20746 7 1 2 20715 20745
0 20747 5 1 1 20746
0 20748 7 1 2 61696 20747
0 20749 5 1 1 20748
0 20750 7 1 2 59516 2041
0 20751 7 1 2 89973 90132
0 20752 7 1 2 20750 20751
0 20753 7 1 2 91615 20752
0 20754 5 1 1 20753
0 20755 7 1 2 20749 20754
0 20756 5 1 1 20755
0 20757 7 1 2 63950 20756
0 20758 5 1 1 20757
0 20759 7 1 2 65393 70259
0 20760 7 1 2 90086 20759
0 20761 5 1 1 20760
0 20762 7 1 2 65394 13716
0 20763 5 1 1 20762
0 20764 7 1 2 74992 75013
0 20765 7 1 2 86381 20764
0 20766 7 1 2 20763 20765
0 20767 5 1 1 20766
0 20768 7 1 2 20761 20767
0 20769 5 1 1 20768
0 20770 7 1 2 86132 20769
0 20771 5 1 1 20770
0 20772 7 1 2 91670 92223
0 20773 5 1 1 20772
0 20774 7 1 2 60508 89485
0 20775 5 1 1 20774
0 20776 7 1 2 20773 20775
0 20777 5 1 1 20776
0 20778 7 1 2 61318 20777
0 20779 5 1 1 20778
0 20780 7 3 2 61506 71201
0 20781 5 3 1 92239
0 20782 7 1 2 73266 92242
0 20783 5 3 1 20782
0 20784 7 1 2 59517 91756
0 20785 7 1 2 92245 20784
0 20786 5 1 1 20785
0 20787 7 1 2 20779 20786
0 20788 5 1 1 20787
0 20789 7 1 2 90108 20788
0 20790 5 1 1 20789
0 20791 7 1 2 20771 20790
0 20792 5 1 1 20791
0 20793 7 1 2 66679 20792
0 20794 5 1 1 20793
0 20795 7 2 2 78754 92024
0 20796 7 1 2 91633 92248
0 20797 5 1 1 20796
0 20798 7 2 2 74930 85549
0 20799 5 1 1 92250
0 20800 7 2 2 59518 92251
0 20801 5 1 1 92252
0 20802 7 1 2 20801 20653
0 20803 5 1 1 20802
0 20804 7 1 2 81175 20803
0 20805 5 1 1 20804
0 20806 7 1 2 20797 20805
0 20807 5 1 1 20806
0 20808 7 1 2 67058 20807
0 20809 5 1 1 20808
0 20810 7 4 2 59519 68860
0 20811 7 1 2 83531 90899
0 20812 7 1 2 92254 20811
0 20813 7 1 2 85748 20812
0 20814 5 1 1 20813
0 20815 7 1 2 20809 20814
0 20816 5 1 1 20815
0 20817 7 1 2 72925 20816
0 20818 5 1 1 20817
0 20819 7 1 2 61697 90932
0 20820 7 1 2 92253 20819
0 20821 5 1 1 20820
0 20822 7 1 2 62971 20821
0 20823 7 1 2 20818 20822
0 20824 7 1 2 20794 20823
0 20825 7 1 2 20758 20824
0 20826 5 1 1 20825
0 20827 7 1 2 61507 73175
0 20828 5 1 1 20827
0 20829 7 1 2 80407 20828
0 20830 7 1 2 92191 20829
0 20831 5 1 1 20830
0 20832 7 1 2 82608 84265
0 20833 7 1 2 81398 20832
0 20834 5 1 1 20833
0 20835 7 1 2 20831 20834
0 20836 5 2 1 20835
0 20837 7 1 2 89924 92258
0 20838 5 1 1 20837
0 20839 7 1 2 90791 89316
0 20840 5 1 1 20839
0 20841 7 1 2 89456 20840
0 20842 5 1 1 20841
0 20843 7 1 2 74993 83935
0 20844 7 1 2 20842 20843
0 20845 5 1 1 20844
0 20846 7 1 2 20838 20845
0 20847 5 1 1 20846
0 20848 7 1 2 59520 20847
0 20849 5 1 1 20848
0 20850 7 2 2 73962 90194
0 20851 7 1 2 81390 72951
0 20852 7 1 2 92260 20851
0 20853 5 1 1 20852
0 20854 7 1 2 20849 20853
0 20855 5 1 1 20854
0 20856 7 1 2 63951 20855
0 20857 5 1 1 20856
0 20858 7 1 2 88617 89409
0 20859 5 1 1 20858
0 20860 7 1 2 75110 90836
0 20861 5 1 1 20860
0 20862 7 1 2 20859 20861
0 20863 5 1 1 20862
0 20864 7 1 2 87932 20863
0 20865 5 1 1 20864
0 20866 7 1 2 67971 20865
0 20867 7 1 2 20857 20866
0 20868 5 1 1 20867
0 20869 7 1 2 20826 20868
0 20870 5 1 1 20869
0 20871 7 1 2 61047 74098
0 20872 7 2 2 74681 20871
0 20873 5 1 1 92262
0 20874 7 11 2 66680 63721
0 20875 7 3 2 80537 92264
0 20876 7 1 2 90647 92275
0 20877 7 1 2 92263 20876
0 20878 5 1 1 20877
0 20879 7 1 2 20870 20878
0 20880 5 1 1 20879
0 20881 7 1 2 86746 20880
0 20882 5 1 1 20881
0 20883 7 10 2 65557 68328
0 20884 5 2 1 92278
0 20885 7 2 2 85339 92279
0 20886 7 3 2 68861 92290
0 20887 7 2 2 87591 91757
0 20888 7 1 2 70604 92295
0 20889 7 1 2 89641 20888
0 20890 7 1 2 92292 20889
0 20891 5 3 1 20890
0 20892 7 1 2 20882 92297
0 20893 5 1 1 20892
0 20894 7 1 2 69109 20893
0 20895 5 1 1 20894
0 20896 7 4 2 60655 61048
0 20897 7 2 2 80862 92300
0 20898 7 1 2 79734 92304
0 20899 5 1 1 20898
0 20900 7 13 2 60656 66681
0 20901 5 1 1 92306
0 20902 7 4 2 61859 92307
0 20903 7 2 2 79036 92319
0 20904 5 1 1 92323
0 20905 7 5 2 65395 92324
0 20906 5 1 1 92325
0 20907 7 7 2 68655 86969
0 20908 7 2 2 90139 92330
0 20909 7 3 2 60327 65558
0 20910 7 1 2 61049 92339
0 20911 7 1 2 92337 20910
0 20912 5 1 1 20911
0 20913 7 1 2 20906 20912
0 20914 5 1 1 20913
0 20915 7 1 2 68862 74968
0 20916 7 1 2 20914 20915
0 20917 5 1 1 20916
0 20918 7 1 2 20899 20917
0 20919 5 1 1 20918
0 20920 7 1 2 61508 20919
0 20921 5 1 1 20920
0 20922 7 2 2 63722 86463
0 20923 7 4 2 60328 60657
0 20924 7 5 2 60509 61050
0 20925 7 1 2 92344 92348
0 20926 7 1 2 92342 20925
0 20927 5 1 1 20926
0 20928 7 1 2 20921 20927
0 20929 5 1 1 20928
0 20930 7 1 2 73760 20929
0 20931 5 1 1 20930
0 20932 7 6 2 60510 60658
0 20933 5 1 1 92353
0 20934 7 4 2 75492 92354
0 20935 7 1 2 92343 92359
0 20936 5 1 1 20935
0 20937 7 1 2 20931 20936
0 20938 5 1 1 20937
0 20939 7 1 2 62972 13242
0 20940 5 1 1 20939
0 20941 7 1 2 20938 20940
0 20942 5 1 1 20941
0 20943 7 1 2 20895 20942
0 20944 7 1 2 20689 20943
0 20945 5 1 1 20944
0 20946 7 1 2 69901 20945
0 20947 5 1 1 20946
0 20948 7 1 2 75833 89518
0 20949 5 2 1 20948
0 20950 7 2 2 59307 79825
0 20951 7 2 2 59858 83403
0 20952 5 1 1 92367
0 20953 7 1 2 92365 92368
0 20954 5 1 1 20953
0 20955 7 1 2 92363 20954
0 20956 5 1 1 20955
0 20957 7 1 2 85510 20956
0 20958 5 1 1 20957
0 20959 7 1 2 73409 83767
0 20960 7 1 2 92051 20959
0 20961 5 1 1 20960
0 20962 7 1 2 20958 20961
0 20963 5 1 1 20962
0 20964 7 1 2 66682 20963
0 20965 5 1 1 20964
0 20966 7 8 2 61698 77550
0 20967 5 2 1 92369
0 20968 7 1 2 76772 75941
0 20969 5 1 1 20968
0 20970 7 2 2 61319 84598
0 20971 5 1 1 92379
0 20972 7 1 2 20969 20971
0 20973 5 1 1 20972
0 20974 7 1 2 79769 20973
0 20975 5 1 1 20974
0 20976 7 1 2 73410 82406
0 20977 7 1 2 91922 20976
0 20978 5 1 1 20977
0 20979 7 1 2 20975 20978
0 20980 5 1 1 20979
0 20981 7 1 2 92370 20980
0 20982 5 1 1 20981
0 20983 7 1 2 20965 20982
0 20984 5 1 1 20983
0 20985 7 1 2 65396 20984
0 20986 5 1 1 20985
0 20987 7 2 2 60511 80994
0 20988 5 2 1 92381
0 20989 7 1 2 91925 92382
0 20990 5 1 1 20989
0 20991 7 1 2 85446 89948
0 20992 5 1 1 20991
0 20993 7 1 2 74994 75787
0 20994 7 1 2 91809 20993
0 20995 5 1 1 20994
0 20996 7 1 2 20992 20995
0 20997 5 1 1 20996
0 20998 7 1 2 67059 20997
0 20999 5 1 1 20998
0 21000 7 1 2 20990 20999
0 21001 5 1 1 21000
0 21002 7 1 2 67972 21001
0 21003 5 1 1 21002
0 21004 7 4 2 81103 79011
0 21005 7 2 2 60329 74343
0 21006 7 1 2 92385 92389
0 21007 5 1 1 21006
0 21008 7 1 2 21003 21007
0 21009 5 1 1 21008
0 21010 7 1 2 59859 21009
0 21011 5 1 1 21010
0 21012 7 2 2 83532 89808
0 21013 7 1 2 75878 73713
0 21014 7 1 2 92391 21013
0 21015 5 1 1 21014
0 21016 7 1 2 80809 91810
0 21017 5 1 1 21016
0 21018 7 1 2 21015 21017
0 21019 5 1 1 21018
0 21020 7 1 2 77374 21019
0 21021 5 1 1 21020
0 21022 7 1 2 21011 21021
0 21023 5 1 1 21022
0 21024 7 1 2 60122 21023
0 21025 5 1 1 21024
0 21026 7 2 2 81496 83359
0 21027 5 1 1 92393
0 21028 7 1 2 80323 86885
0 21029 5 2 1 21028
0 21030 7 1 2 68656 75942
0 21031 7 1 2 92395 21030
0 21032 5 1 1 21031
0 21033 7 1 2 21027 21032
0 21034 5 1 1 21033
0 21035 7 1 2 90599 21034
0 21036 5 1 1 21035
0 21037 7 1 2 21025 21036
0 21038 5 1 1 21037
0 21039 7 1 2 63952 21038
0 21040 5 1 1 21039
0 21041 7 1 2 20986 21040
0 21042 5 1 1 21041
0 21043 7 1 2 71717 21042
0 21044 5 1 1 21043
0 21045 7 1 2 75564 80375
0 21046 5 1 1 21045
0 21047 7 3 2 14173 21046
0 21048 7 2 2 70162 92397
0 21049 7 2 2 67973 79856
0 21050 7 1 2 92400 92402
0 21051 5 1 1 21050
0 21052 7 1 2 81793 91418
0 21053 5 1 1 21052
0 21054 7 2 2 85447 86537
0 21055 5 2 1 92404
0 21056 7 5 2 61509 76773
0 21057 5 1 1 92408
0 21058 7 1 2 80408 92409
0 21059 5 1 1 21058
0 21060 7 1 2 92406 21059
0 21061 7 1 2 21053 21060
0 21062 5 1 1 21061
0 21063 7 1 2 80112 21062
0 21064 5 1 1 21063
0 21065 7 1 2 21051 21064
0 21066 5 1 1 21065
0 21067 7 1 2 68657 21066
0 21068 5 1 1 21067
0 21069 7 2 2 61699 75289
0 21070 5 6 1 92413
0 21071 7 1 2 85132 85973
0 21072 7 1 2 92414 21071
0 21073 5 1 1 21072
0 21074 7 1 2 21068 21073
0 21075 5 1 1 21074
0 21076 7 1 2 63953 21075
0 21077 5 1 1 21076
0 21078 7 1 2 71556 74687
0 21079 5 1 1 21078
0 21080 7 2 2 80113 84427
0 21081 7 1 2 84166 88127
0 21082 7 1 2 92421 21081
0 21083 7 1 2 21079 21082
0 21084 5 1 1 21083
0 21085 7 1 2 21077 21084
0 21086 5 1 1 21085
0 21087 7 1 2 67060 21086
0 21088 5 1 1 21087
0 21089 7 1 2 79908 88105
0 21090 5 1 1 21089
0 21091 7 1 2 86696 21090
0 21092 5 1 1 21091
0 21093 7 1 2 80680 21092
0 21094 5 1 1 21093
0 21095 7 1 2 79728 89344
0 21096 5 1 1 21095
0 21097 7 1 2 21094 21096
0 21098 5 1 1 21097
0 21099 7 1 2 60330 21098
0 21100 5 1 1 21099
0 21101 7 4 2 79743 82172
0 21102 7 1 2 66475 87756
0 21103 7 1 2 92423 21102
0 21104 5 1 1 21103
0 21105 7 1 2 21100 21104
0 21106 5 1 1 21105
0 21107 7 1 2 63723 21106
0 21108 5 1 1 21107
0 21109 7 1 2 21088 21108
0 21110 5 1 1 21109
0 21111 7 1 2 69551 21110
0 21112 5 1 1 21111
0 21113 7 1 2 85340 92398
0 21114 5 1 1 21113
0 21115 7 1 2 83781 91811
0 21116 5 1 1 21115
0 21117 7 1 2 21114 21116
0 21118 5 1 1 21117
0 21119 7 1 2 70605 21118
0 21120 5 1 1 21119
0 21121 7 2 2 84378 89768
0 21122 5 1 1 92427
0 21123 7 1 2 86232 92428
0 21124 5 1 1 21123
0 21125 7 2 2 75290 85783
0 21126 7 1 2 59860 92429
0 21127 5 1 1 21126
0 21128 7 3 2 82407 84338
0 21129 5 2 1 92431
0 21130 7 1 2 60331 92432
0 21131 5 1 1 21130
0 21132 7 1 2 21127 21131
0 21133 5 1 1 21132
0 21134 7 1 2 60512 21133
0 21135 5 1 1 21134
0 21136 7 1 2 21124 21135
0 21137 7 1 2 21120 21136
0 21138 5 1 1 21137
0 21139 7 1 2 68329 21138
0 21140 5 1 1 21139
0 21141 7 1 2 60513 79482
0 21142 5 2 1 21141
0 21143 7 2 2 74344 83000
0 21144 5 1 1 92438
0 21145 7 1 2 83711 21144
0 21146 5 2 1 21145
0 21147 7 1 2 60332 92440
0 21148 5 1 1 21147
0 21149 7 1 2 92436 21148
0 21150 5 1 1 21149
0 21151 7 1 2 91893 21150
0 21152 5 1 1 21151
0 21153 7 1 2 63724 91359
0 21154 7 1 2 89509 21153
0 21155 5 1 1 21154
0 21156 7 1 2 21152 21155
0 21157 5 1 1 21156
0 21158 7 1 2 61700 21157
0 21159 5 1 1 21158
0 21160 7 2 2 68658 84684
0 21161 7 1 2 92117 92442
0 21162 5 1 1 21161
0 21163 7 1 2 21159 21162
0 21164 5 1 1 21163
0 21165 7 1 2 79909 21164
0 21166 5 1 1 21165
0 21167 7 1 2 21140 21166
0 21168 5 1 1 21167
0 21169 7 1 2 63954 21168
0 21170 5 1 1 21169
0 21171 7 1 2 21112 21170
0 21172 5 1 1 21171
0 21173 7 1 2 72104 21172
0 21174 5 1 1 21173
0 21175 7 2 2 60123 84476
0 21176 5 1 1 92444
0 21177 7 1 2 80245 84339
0 21178 5 1 1 21177
0 21179 7 1 2 21176 21178
0 21180 5 1 1 21179
0 21181 7 1 2 61320 21180
0 21182 5 1 1 21181
0 21183 7 1 2 84544 91805
0 21184 5 2 1 21183
0 21185 7 1 2 80928 92446
0 21186 5 1 1 21185
0 21187 7 1 2 83143 84477
0 21188 5 1 1 21187
0 21189 7 1 2 21186 21188
0 21190 5 1 1 21189
0 21191 7 1 2 74590 21190
0 21192 5 1 1 21191
0 21193 7 1 2 21182 21192
0 21194 5 1 1 21193
0 21195 7 1 2 60514 21194
0 21196 5 1 1 21195
0 21197 7 7 2 59521 68659
0 21198 7 5 2 61701 69552
0 21199 7 3 2 92448 92455
0 21200 7 1 2 69182 89648
0 21201 7 1 2 92460 21200
0 21202 5 1 1 21201
0 21203 7 1 2 21196 21202
0 21204 5 1 1 21203
0 21205 7 1 2 63955 21204
0 21206 5 1 1 21205
0 21207 7 1 2 64957 80698
0 21208 5 1 1 21207
0 21209 7 1 2 80681 83664
0 21210 7 1 2 82253 21209
0 21211 7 1 2 21208 21210
0 21212 5 1 1 21211
0 21213 7 1 2 21206 21212
0 21214 5 1 1 21213
0 21215 7 1 2 67974 21214
0 21216 5 1 1 21215
0 21217 7 2 2 84340 88893
0 21218 7 1 2 74591 92463
0 21219 5 1 1 21218
0 21220 7 1 2 83936 89857
0 21221 5 1 1 21220
0 21222 7 1 2 67061 91801
0 21223 5 1 1 21222
0 21224 7 1 2 21221 21223
0 21225 5 1 1 21224
0 21226 7 1 2 88752 21225
0 21227 5 1 1 21226
0 21228 7 1 2 21219 21227
0 21229 5 1 1 21228
0 21230 7 1 2 60124 79132
0 21231 7 1 2 21229 21230
0 21232 5 1 1 21231
0 21233 7 1 2 21216 21232
0 21234 5 1 1 21233
0 21235 7 1 2 63415 21234
0 21236 5 1 1 21235
0 21237 7 1 2 70052 80265
0 21238 5 1 1 21237
0 21239 7 1 2 87913 89855
0 21240 7 1 2 21238 21239
0 21241 5 1 1 21240
0 21242 7 1 2 21236 21241
0 21243 5 1 1 21242
0 21244 7 1 2 75291 21243
0 21245 5 1 1 21244
0 21246 7 1 2 9059 91400
0 21247 5 2 1 21246
0 21248 7 2 2 60125 61702
0 21249 7 1 2 92465 92467
0 21250 5 1 1 21249
0 21251 7 1 2 81176 91788
0 21252 5 1 1 21251
0 21253 7 1 2 21250 21252
0 21254 5 1 1 21253
0 21255 7 1 2 60333 21254
0 21256 5 1 1 21255
0 21257 7 2 2 67975 89809
0 21258 7 1 2 85589 92469
0 21259 5 1 1 21258
0 21260 7 1 2 78128 86869
0 21261 5 1 1 21260
0 21262 7 1 2 86886 21261
0 21263 5 1 1 21262
0 21264 7 1 2 60515 21263
0 21265 5 1 1 21264
0 21266 7 1 2 21259 21265
0 21267 7 1 2 21256 21266
0 21268 5 1 1 21267
0 21269 7 1 2 80260 21268
0 21270 5 1 1 21269
0 21271 7 2 2 60516 92396
0 21272 5 1 1 92471
0 21273 7 1 2 86233 92441
0 21274 5 1 1 21273
0 21275 7 1 2 21272 21274
0 21276 5 1 1 21275
0 21277 7 1 2 73550 21276
0 21278 5 1 1 21277
0 21279 7 1 2 21270 21278
0 21280 5 1 1 21279
0 21281 7 1 2 68660 21280
0 21282 5 1 1 21281
0 21283 7 1 2 62973 78359
0 21284 5 1 1 21283
0 21285 7 1 2 59861 21284
0 21286 5 2 1 21285
0 21287 7 1 2 67976 82561
0 21288 5 1 1 21287
0 21289 7 1 2 92473 21288
0 21290 5 1 1 21289
0 21291 7 1 2 70163 21290
0 21292 5 1 1 21291
0 21293 7 9 2 60126 75713
0 21294 5 2 1 92475
0 21295 7 1 2 74521 92476
0 21296 5 1 1 21295
0 21297 7 1 2 21292 21296
0 21298 5 1 1 21297
0 21299 7 1 2 75292 21298
0 21300 5 1 1 21299
0 21301 7 1 2 79885 81372
0 21302 5 1 1 21301
0 21303 7 1 2 21300 21302
0 21304 5 1 1 21303
0 21305 7 1 2 83152 21304
0 21306 5 1 1 21305
0 21307 7 1 2 21282 21306
0 21308 5 1 1 21307
0 21309 7 1 2 63416 21308
0 21310 5 1 1 21309
0 21311 7 1 2 81828 92401
0 21312 5 1 1 21311
0 21313 7 1 2 80409 89024
0 21314 5 1 1 21313
0 21315 7 1 2 87839 21314
0 21316 7 1 2 21312 21315
0 21317 5 1 1 21316
0 21318 7 1 2 83768 21317
0 21319 5 1 1 21318
0 21320 7 1 2 21310 21319
0 21321 5 1 1 21320
0 21322 7 1 2 63956 21321
0 21323 5 1 1 21322
0 21324 7 1 2 64958 91533
0 21325 5 5 1 21324
0 21326 7 1 2 74969 86693
0 21327 5 1 1 21326
0 21328 7 1 2 89477 21327
0 21329 5 1 1 21328
0 21330 7 1 2 92486 21329
0 21331 5 1 1 21330
0 21332 7 1 2 76497 80145
0 21333 5 1 1 21332
0 21334 7 1 2 92364 21333
0 21335 5 1 1 21334
0 21336 7 1 2 69110 21335
0 21337 5 1 1 21336
0 21338 7 1 2 79915 74682
0 21339 7 1 2 83382 21338
0 21340 5 1 1 21339
0 21341 7 1 2 21337 21340
0 21342 7 1 2 21331 21341
0 21343 5 1 1 21342
0 21344 7 1 2 67062 21343
0 21345 5 1 1 21344
0 21346 7 1 2 75565 80249
0 21347 5 1 1 21346
0 21348 7 1 2 63417 90003
0 21349 7 1 2 21347 21348
0 21350 5 1 1 21349
0 21351 7 1 2 21345 21350
0 21352 5 1 1 21351
0 21353 7 1 2 87933 21352
0 21354 5 1 1 21353
0 21355 7 1 2 21323 21354
0 21356 5 1 1 21355
0 21357 7 1 2 69902 21356
0 21358 5 1 1 21357
0 21359 7 1 2 67296 85784
0 21360 5 1 1 21359
0 21361 7 1 2 92434 21360
0 21362 5 1 1 21361
0 21363 7 1 2 60517 21362
0 21364 5 1 1 21363
0 21365 7 1 2 79258 85353
0 21366 5 1 1 21365
0 21367 7 1 2 21364 21366
0 21368 5 1 1 21367
0 21369 7 1 2 68330 21368
0 21370 5 1 1 21369
0 21371 7 2 2 79770 90195
0 21372 7 2 2 65397 92491
0 21373 7 1 2 73013 92493
0 21374 5 1 1 21373
0 21375 7 1 2 21370 21374
0 21376 5 1 1 21375
0 21377 7 1 2 61321 21376
0 21378 5 1 1 21377
0 21379 7 1 2 73643 84819
0 21380 7 1 2 89556 21379
0 21381 5 1 1 21380
0 21382 7 1 2 21378 21381
0 21383 5 1 1 21382
0 21384 7 1 2 60127 21383
0 21385 5 1 1 21384
0 21386 7 1 2 82978 85448
0 21387 7 1 2 92392 21386
0 21388 5 1 1 21387
0 21389 7 1 2 21385 21388
0 21390 5 1 1 21389
0 21391 7 1 2 59862 21390
0 21392 5 1 1 21391
0 21393 7 2 2 73668 73972
0 21394 5 1 1 92495
0 21395 7 1 2 82862 92496
0 21396 5 1 1 21395
0 21397 7 1 2 85625 21396
0 21398 5 1 1 21397
0 21399 7 1 2 61703 21398
0 21400 5 1 1 21399
0 21401 7 1 2 79436 91360
0 21402 5 1 1 21401
0 21403 7 1 2 21400 21402
0 21404 5 1 1 21403
0 21405 7 1 2 89769 21404
0 21406 5 1 1 21405
0 21407 7 1 2 79437 87757
0 21408 5 1 1 21407
0 21409 7 1 2 67297 81802
0 21410 5 1 1 21409
0 21411 7 1 2 21408 21410
0 21412 5 1 1 21411
0 21413 7 1 2 65398 21412
0 21414 5 1 1 21413
0 21415 7 3 2 63418 80354
0 21416 5 1 1 92497
0 21417 7 1 2 73014 92498
0 21418 5 1 1 21417
0 21419 7 1 2 68661 21418
0 21420 7 1 2 21414 21419
0 21421 5 1 1 21420
0 21422 7 3 2 68331 79647
0 21423 7 2 2 73669 83001
0 21424 7 1 2 92500 92503
0 21425 5 1 1 21424
0 21426 7 1 2 63725 3885
0 21427 7 1 2 21425 21426
0 21428 5 1 1 21427
0 21429 7 1 2 61510 21428
0 21430 7 1 2 21421 21429
0 21431 5 1 1 21430
0 21432 7 1 2 21406 21431
0 21433 5 1 1 21432
0 21434 7 1 2 59863 21433
0 21435 5 1 1 21434
0 21436 7 1 2 80410 89770
0 21437 7 1 2 91923 21436
0 21438 5 1 1 21437
0 21439 7 4 2 61704 79037
0 21440 7 1 2 89337 92505
0 21441 5 1 1 21440
0 21442 7 1 2 21438 21441
0 21443 5 1 1 21442
0 21444 7 1 2 67977 21443
0 21445 5 1 1 21444
0 21446 7 1 2 21435 21445
0 21447 5 1 1 21446
0 21448 7 1 2 60334 21447
0 21449 5 1 1 21448
0 21450 7 1 2 92065 92386
0 21451 5 1 1 21450
0 21452 7 1 2 21449 21451
0 21453 7 1 2 21392 21452
0 21454 5 1 1 21453
0 21455 7 1 2 63957 21454
0 21456 5 1 1 21455
0 21457 7 1 2 80572 92407
0 21458 5 1 1 21457
0 21459 7 1 2 63419 21458
0 21460 5 1 1 21459
0 21461 7 1 2 83741 83144
0 21462 7 1 2 92399 21461
0 21463 5 1 1 21462
0 21464 7 1 2 21460 21463
0 21465 5 1 1 21464
0 21466 7 1 2 77551 21465
0 21467 5 1 1 21466
0 21468 7 2 2 80114 85511
0 21469 5 1 1 92509
0 21470 7 1 2 84232 92510
0 21471 5 1 1 21470
0 21472 7 1 2 21467 21471
0 21473 5 1 1 21472
0 21474 7 1 2 80717 21473
0 21475 5 1 1 21474
0 21476 7 5 2 61322 61705
0 21477 7 3 2 77901 77552
0 21478 7 2 2 75293 92516
0 21479 7 1 2 92511 92519
0 21480 5 1 1 21479
0 21481 7 1 2 76387 89683
0 21482 5 1 1 21481
0 21483 7 1 2 61323 89704
0 21484 5 1 1 21483
0 21485 7 1 2 21482 21484
0 21486 5 1 1 21485
0 21487 7 6 2 59864 68863
0 21488 7 1 2 80995 92521
0 21489 7 1 2 21486 21488
0 21490 5 1 1 21489
0 21491 7 1 2 21480 21490
0 21492 5 1 1 21491
0 21493 7 1 2 65399 21492
0 21494 5 1 1 21493
0 21495 7 1 2 91407 92520
0 21496 5 1 1 21495
0 21497 7 1 2 21494 21496
0 21498 5 1 1 21497
0 21499 7 1 2 78321 21498
0 21500 5 1 1 21499
0 21501 7 1 2 84233 73411
0 21502 7 1 2 85550 21501
0 21503 5 1 1 21502
0 21504 7 1 2 21500 21503
0 21505 7 1 2 21475 21504
0 21506 7 1 2 21456 21505
0 21507 7 1 2 21358 21506
0 21508 7 1 2 21245 21507
0 21509 7 1 2 21174 21508
0 21510 7 1 2 21044 21509
0 21511 5 1 1 21510
0 21512 7 1 2 86747 21511
0 21513 5 1 1 21512
0 21514 7 5 2 60659 86208
0 21515 5 1 1 92527
0 21516 7 4 2 66476 79744
0 21517 7 1 2 72806 82988
0 21518 7 1 2 92532 21517
0 21519 5 1 1 21518
0 21520 7 2 2 60128 78372
0 21521 5 1 1 92536
0 21522 7 1 2 79900 21521
0 21523 5 1 1 21522
0 21524 7 6 2 59865 61706
0 21525 5 1 1 92538
0 21526 7 1 2 81093 92539
0 21527 7 1 2 21523 21526
0 21528 5 1 1 21527
0 21529 7 1 2 21519 21528
0 21530 5 1 1 21529
0 21531 7 1 2 65400 21530
0 21532 5 1 1 21531
0 21533 7 1 2 63958 76558
0 21534 7 1 2 92472 21533
0 21535 5 1 1 21534
0 21536 7 1 2 21532 21535
0 21537 5 1 1 21536
0 21538 7 1 2 68662 21537
0 21539 5 1 1 21538
0 21540 7 5 2 67298 63959
0 21541 7 1 2 80863 92544
0 21542 5 1 1 21541
0 21543 7 1 2 60129 80682
0 21544 5 1 1 21543
0 21545 7 1 2 21542 21544
0 21546 5 2 1 21545
0 21547 7 1 2 83841 92549
0 21548 5 1 1 21547
0 21549 7 1 2 21539 21548
0 21550 5 1 1 21549
0 21551 7 1 2 92528 21550
0 21552 5 1 1 21551
0 21553 7 1 2 85133 89810
0 21554 5 2 1 21553
0 21555 7 1 2 59866 92012
0 21556 5 1 1 21555
0 21557 7 1 2 92551 21556
0 21558 5 1 1 21557
0 21559 7 5 2 63960 75294
0 21560 7 6 2 61860 67299
0 21561 7 1 2 87620 92558
0 21562 7 1 2 92553 21561
0 21563 7 1 2 21558 21562
0 21564 5 1 1 21563
0 21565 7 2 2 65401 87015
0 21566 7 2 2 92559 92564
0 21567 7 1 2 92265 92566
0 21568 5 1 1 21567
0 21569 7 5 2 66825 67063
0 21570 7 2 2 87628 92568
0 21571 7 1 2 89998 92118
0 21572 7 1 2 92573 21571
0 21573 5 1 1 21572
0 21574 7 1 2 21568 21573
0 21575 5 1 1 21574
0 21576 7 1 2 68864 80783
0 21577 7 1 2 21575 21576
0 21578 5 1 1 21577
0 21579 7 1 2 21564 21578
0 21580 5 1 1 21579
0 21581 7 1 2 67978 21580
0 21582 5 1 1 21581
0 21583 7 1 2 67300 80695
0 21584 5 1 1 21583
0 21585 7 2 2 61511 80411
0 21586 5 1 1 92575
0 21587 7 1 2 60335 91419
0 21588 5 1 1 21587
0 21589 7 1 2 21586 21588
0 21590 5 1 1 21589
0 21591 7 1 2 63961 73412
0 21592 7 1 2 21590 21591
0 21593 5 1 1 21592
0 21594 7 1 2 21584 21593
0 21595 5 1 1 21594
0 21596 7 1 2 86429 92529
0 21597 7 1 2 21595 21596
0 21598 5 1 1 21597
0 21599 7 1 2 21582 21598
0 21600 5 1 1 21599
0 21601 7 1 2 61324 21600
0 21602 5 1 1 21601
0 21603 7 1 2 21552 21602
0 21604 5 1 1 21603
0 21605 7 1 2 88769 21604
0 21606 5 1 1 21605
0 21607 7 1 2 59867 77241
0 21608 5 1 1 21607
0 21609 7 1 2 73306 21608
0 21610 5 1 1 21609
0 21611 7 1 2 69111 21610
0 21612 5 1 1 21611
0 21613 7 1 2 72879 86489
0 21614 5 1 1 21613
0 21615 7 1 2 67301 21614
0 21616 5 1 1 21615
0 21617 7 2 2 67302 72515
0 21618 5 2 1 92577
0 21619 7 1 2 81608 82774
0 21620 7 1 2 92579 21619
0 21621 5 1 1 21620
0 21622 7 1 2 59522 21621
0 21623 5 1 1 21622
0 21624 7 1 2 21616 21623
0 21625 7 1 2 21612 21624
0 21626 5 1 1 21625
0 21627 7 3 2 65559 89925
0 21628 7 2 2 87094 92581
0 21629 5 1 1 92584
0 21630 7 2 2 87333 92585
0 21631 7 1 2 90066 92586
0 21632 7 1 2 21626 21631
0 21633 5 1 1 21632
0 21634 7 1 2 21606 21633
0 21635 7 1 2 21513 21634
0 21636 5 1 1 21635
0 21637 7 1 2 73815 21636
0 21638 5 1 1 21637
0 21639 7 2 2 78755 72980
0 21640 7 1 2 66477 92588
0 21641 5 1 1 21640
0 21642 7 7 2 66478 83533
0 21643 5 1 1 92590
0 21644 7 1 2 67303 92591
0 21645 5 1 1 21644
0 21646 7 1 2 89979 21645
0 21647 5 1 1 21646
0 21648 7 1 2 65191 21647
0 21649 5 1 1 21648
0 21650 7 1 2 21641 21649
0 21651 5 1 1 21650
0 21652 7 1 2 88128 21651
0 21653 5 1 1 21652
0 21654 7 4 2 75295 83534
0 21655 7 2 2 79133 72672
0 21656 7 1 2 92597 92601
0 21657 5 1 1 21656
0 21658 7 1 2 21653 21657
0 21659 5 1 1 21658
0 21660 7 1 2 66683 21659
0 21661 5 1 1 21660
0 21662 7 1 2 63962 72673
0 21663 7 1 2 92494 21662
0 21664 5 1 1 21663
0 21665 7 1 2 21661 21664
0 21666 5 1 1 21665
0 21667 7 3 2 69903 75997
0 21668 5 1 1 92603
0 21669 7 1 2 21666 92604
0 21670 5 1 1 21669
0 21671 7 1 2 67606 73935
0 21672 5 1 1 21671
0 21673 7 1 2 14004 21672
0 21674 5 1 1 21673
0 21675 7 1 2 75296 80355
0 21676 5 1 1 21675
0 21677 7 1 2 89558 21676
0 21678 5 2 1 21677
0 21679 7 1 2 21674 92606
0 21680 5 1 1 21679
0 21681 7 1 2 80573 21680
0 21682 5 1 1 21681
0 21683 7 1 2 92545 21682
0 21684 5 1 1 21683
0 21685 7 1 2 80696 88905
0 21686 5 1 1 21685
0 21687 7 1 2 21684 21686
0 21688 5 1 1 21687
0 21689 7 2 2 68663 69904
0 21690 5 1 1 92608
0 21691 7 1 2 21688 92609
0 21692 5 1 1 21691
0 21693 7 1 2 78053 92349
0 21694 5 2 1 21693
0 21695 7 1 2 81308 84417
0 21696 5 1 1 21695
0 21697 7 1 2 87918 21696
0 21698 5 2 1 21697
0 21699 7 1 2 59868 92612
0 21700 5 1 1 21699
0 21701 7 1 2 92610 21700
0 21702 5 1 1 21701
0 21703 7 1 2 60130 21702
0 21704 5 1 1 21703
0 21705 7 1 2 81333 81391
0 21706 5 1 1 21705
0 21707 7 1 2 21704 21706
0 21708 5 1 1 21707
0 21709 7 1 2 61512 21708
0 21710 5 1 1 21709
0 21711 7 1 2 86234 92602
0 21712 5 1 1 21711
0 21713 7 1 2 21710 21712
0 21714 5 1 1 21713
0 21715 7 1 2 69553 21714
0 21716 5 1 1 21715
0 21717 7 1 2 81334 89649
0 21718 5 1 1 21717
0 21719 7 1 2 21718 92611
0 21720 5 1 1 21719
0 21721 7 1 2 59869 21720
0 21722 5 1 1 21721
0 21723 7 1 2 60131 92613
0 21724 5 1 1 21723
0 21725 7 1 2 21722 21724
0 21726 5 1 1 21725
0 21727 7 1 2 69554 21726
0 21728 5 1 1 21727
0 21729 7 1 2 72224 92550
0 21730 5 1 1 21729
0 21731 7 1 2 79745 81392
0 21732 5 1 1 21731
0 21733 7 2 2 80929 81751
0 21734 5 1 1 92614
0 21735 7 1 2 21732 21734
0 21736 7 1 2 21730 21735
0 21737 7 1 2 21728 21736
0 21738 5 1 1 21737
0 21739 7 1 2 61513 21738
0 21740 5 1 1 21739
0 21741 7 3 2 63963 72926
0 21742 7 4 2 61707 90121
0 21743 7 1 2 73714 92619
0 21744 7 1 2 92616 21743
0 21745 5 1 1 21744
0 21746 7 1 2 21740 21745
0 21747 5 1 1 21746
0 21748 7 1 2 67607 21747
0 21749 5 1 1 21748
0 21750 7 1 2 92246 92615
0 21751 5 1 1 21750
0 21752 7 1 2 21749 21751
0 21753 7 1 2 21716 21752
0 21754 5 1 1 21753
0 21755 7 1 2 72105 21754
0 21756 5 1 1 21755
0 21757 7 2 2 69555 81752
0 21758 5 1 1 92623
0 21759 7 1 2 89549 92624
0 21760 5 1 1 21759
0 21761 7 6 2 60914 66684
0 21762 7 1 2 86611 92625
0 21763 7 1 2 90648 21762
0 21764 5 1 1 21763
0 21765 7 1 2 21760 21764
0 21766 5 1 1 21765
0 21767 7 1 2 75297 21766
0 21768 5 1 1 21767
0 21769 7 1 2 82704 21768
0 21770 5 1 1 21769
0 21771 7 1 2 67304 21770
0 21772 5 1 1 21771
0 21773 7 2 2 71718 79826
0 21774 7 3 2 59308 65402
0 21775 7 1 2 86615 92633
0 21776 7 1 2 92631 21775
0 21777 5 1 1 21776
0 21778 7 1 2 78054 72472
0 21779 7 1 2 91846 21778
0 21780 5 1 1 21779
0 21781 7 1 2 21777 21780
0 21782 5 1 1 21781
0 21783 7 1 2 60132 21782
0 21784 5 1 1 21783
0 21785 7 1 2 21772 21784
0 21786 5 1 1 21785
0 21787 7 1 2 71202 21786
0 21788 5 1 1 21787
0 21789 7 1 2 69556 90007
0 21790 5 1 1 21789
0 21791 7 1 2 78225 21790
0 21792 5 1 1 21791
0 21793 7 1 2 72927 21792
0 21794 5 1 1 21793
0 21795 7 1 2 72968 21794
0 21796 5 1 1 21795
0 21797 7 1 2 81753 21796
0 21798 5 1 1 21797
0 21799 7 9 2 66685 67608
0 21800 5 1 1 92636
0 21801 7 3 2 61051 92637
0 21802 7 1 2 83383 88129
0 21803 7 1 2 92645 21802
0 21804 5 1 1 21803
0 21805 7 1 2 21798 21804
0 21806 5 1 1 21805
0 21807 7 1 2 60336 21806
0 21808 5 1 1 21807
0 21809 7 1 2 80683 72981
0 21810 5 1 1 21809
0 21811 7 2 2 60518 92456
0 21812 7 1 2 92617 92648
0 21813 5 1 1 21812
0 21814 7 1 2 21810 21813
0 21815 5 1 1 21814
0 21816 7 1 2 90008 21815
0 21817 5 1 1 21816
0 21818 7 2 2 65403 60796
0 21819 7 2 2 59309 92650
0 21820 7 1 2 86616 92652
0 21821 5 1 1 21820
0 21822 7 1 2 87919 21821
0 21823 5 1 1 21822
0 21824 7 1 2 72982 21823
0 21825 5 1 1 21824
0 21826 7 1 2 80864 78219
0 21827 7 1 2 92618 21826
0 21828 5 1 1 21827
0 21829 7 1 2 21825 21828
0 21830 7 1 2 21817 21829
0 21831 5 1 1 21830
0 21832 7 1 2 61514 21831
0 21833 5 1 1 21832
0 21834 7 1 2 21808 21833
0 21835 7 1 2 21788 21834
0 21836 7 1 2 21756 21835
0 21837 5 1 1 21836
0 21838 7 1 2 63726 21837
0 21839 5 1 1 21838
0 21840 7 1 2 21692 21839
0 21841 5 1 1 21840
0 21842 7 1 2 63420 21841
0 21843 5 1 1 21842
0 21844 7 1 2 21670 21843
0 21845 5 1 1 21844
0 21846 7 1 2 86748 21845
0 21847 5 1 1 21846
0 21848 7 3 2 59523 73413
0 21849 7 4 2 65560 69557
0 21850 7 2 2 92654 92657
0 21851 7 2 2 80762 84284
0 21852 7 12 2 68664 68865
0 21853 7 1 2 68332 92665
0 21854 7 1 2 92296 21853
0 21855 7 1 2 92663 21854
0 21856 7 1 2 92661 21855
0 21857 5 1 1 21856
0 21858 7 1 2 21847 21857
0 21859 5 1 1 21858
0 21860 7 1 2 82962 21859
0 21861 5 1 1 21860
0 21862 7 1 2 5306 74549
0 21863 5 1 1 21862
0 21864 7 1 2 67305 21863
0 21865 5 1 1 21864
0 21866 7 1 2 77662 21865
0 21867 5 1 1 21866
0 21868 7 1 2 75298 21867
0 21869 5 1 1 21868
0 21870 7 1 2 80768 21869
0 21871 5 1 1 21870
0 21872 7 1 2 67979 21871
0 21873 5 1 1 21872
0 21874 7 3 2 64717 72591
0 21875 5 2 1 92677
0 21876 7 2 2 69247 81620
0 21877 5 1 1 92682
0 21878 7 1 2 92678 92683
0 21879 5 1 1 21878
0 21880 7 1 2 60337 21879
0 21881 5 1 1 21880
0 21882 7 2 2 67306 71648
0 21883 7 2 2 76559 76256
0 21884 5 1 1 92686
0 21885 7 1 2 92684 92687
0 21886 5 1 1 21885
0 21887 7 1 2 80643 91461
0 21888 5 1 1 21887
0 21889 7 1 2 73391 21888
0 21890 5 1 1 21889
0 21891 7 1 2 69112 21890
0 21892 5 1 1 21891
0 21893 7 1 2 21886 21892
0 21894 7 1 2 21881 21893
0 21895 5 1 1 21894
0 21896 7 1 2 61515 21895
0 21897 5 1 1 21896
0 21898 7 1 2 21873 21897
0 21899 5 1 1 21898
0 21900 7 1 2 77553 21899
0 21901 5 1 1 21900
0 21902 7 1 2 78911 11746
0 21903 5 1 1 21902
0 21904 7 1 2 87941 21903
0 21905 5 1 1 21904
0 21906 7 1 2 21901 21905
0 21907 5 1 1 21906
0 21908 7 1 2 63421 21907
0 21909 5 1 1 21908
0 21910 7 1 2 82332 83130
0 21911 5 1 1 21910
0 21912 7 1 2 61325 21911
0 21913 5 1 1 21912
0 21914 7 1 2 65192 21913
0 21915 5 1 1 21914
0 21916 7 1 2 82408 90109
0 21917 7 1 2 21915 21916
0 21918 5 1 1 21917
0 21919 7 1 2 21909 21918
0 21920 5 1 1 21919
0 21921 7 1 2 81177 21920
0 21922 5 1 1 21921
0 21923 7 2 2 69905 75299
0 21924 7 1 2 79746 84379
0 21925 5 2 1 21924
0 21926 7 1 2 67064 87914
0 21927 5 1 1 21926
0 21928 7 1 2 92690 21927
0 21929 5 1 1 21928
0 21930 7 1 2 92688 21929
0 21931 5 1 1 21930
0 21932 7 1 2 78129 92020
0 21933 5 1 1 21932
0 21934 7 1 2 21931 21933
0 21935 5 1 1 21934
0 21936 7 1 2 61326 21935
0 21937 5 1 1 21936
0 21938 7 1 2 82705 21937
0 21939 5 1 1 21938
0 21940 7 1 2 67307 21939
0 21941 5 1 1 21940
0 21942 7 3 2 68866 71486
0 21943 7 1 2 84234 92692
0 21944 5 1 1 21943
0 21945 7 1 2 21941 21944
0 21946 5 1 1 21945
0 21947 7 1 2 63727 21946
0 21948 5 1 1 21947
0 21949 7 1 2 80509 81335
0 21950 7 1 2 69723 21949
0 21951 5 1 1 21950
0 21952 7 1 2 87920 21951
0 21953 5 1 1 21952
0 21954 7 1 2 83980 21953
0 21955 5 1 1 21954
0 21956 7 1 2 21948 21955
0 21957 5 1 1 21956
0 21958 7 1 2 63422 21957
0 21959 5 1 1 21958
0 21960 7 1 2 82321 87886
0 21961 5 1 1 21960
0 21962 7 1 2 83302 85512
0 21963 7 1 2 76913 21962
0 21964 5 1 1 21963
0 21965 7 1 2 21961 21964
0 21966 5 1 1 21965
0 21967 7 1 2 82927 87800
0 21968 7 1 2 21966 21967
0 21969 5 1 1 21968
0 21970 7 1 2 21959 21969
0 21971 5 1 1 21970
0 21972 7 1 2 74592 21971
0 21973 5 1 1 21972
0 21974 7 1 2 80469 79229
0 21975 5 1 1 21974
0 21976 7 1 2 7045 21975
0 21977 5 1 1 21976
0 21978 7 1 2 59870 21977
0 21979 5 1 1 21978
0 21980 7 1 2 60797 89580
0 21981 5 1 1 21980
0 21982 7 1 2 89838 21981
0 21983 5 1 1 21982
0 21984 7 1 2 59310 21983
0 21985 5 1 1 21984
0 21986 7 4 2 61516 70275
0 21987 5 1 1 92695
0 21988 7 1 2 60338 92696
0 21989 5 1 1 21988
0 21990 7 1 2 21985 21989
0 21991 5 1 1 21990
0 21992 7 1 2 92060 21991
0 21993 5 1 1 21992
0 21994 7 1 2 21979 21993
0 21995 5 1 1 21994
0 21996 7 1 2 80684 21995
0 21997 5 1 1 21996
0 21998 7 1 2 84089 79230
0 21999 5 1 1 21998
0 22000 7 1 2 80457 78393
0 22001 5 1 1 22000
0 22002 7 1 2 82948 22001
0 22003 5 1 1 22002
0 22004 7 1 2 63728 75300
0 22005 7 1 2 22003 22004
0 22006 5 1 1 22005
0 22007 7 1 2 21999 22006
0 22008 5 1 1 22007
0 22009 7 1 2 60519 22008
0 22010 5 1 1 22009
0 22011 7 1 2 78394 92238
0 22012 5 1 1 22011
0 22013 7 1 2 73670 89771
0 22014 7 1 2 82871 22013
0 22015 5 1 1 22014
0 22016 7 1 2 22012 22015
0 22017 5 1 1 22016
0 22018 7 1 2 82496 22017
0 22019 5 1 1 22018
0 22020 7 1 2 22010 22019
0 22021 5 1 1 22020
0 22022 7 1 2 61708 22021
0 22023 5 1 1 22022
0 22024 7 3 2 59871 90122
0 22025 7 1 2 69558 92699
0 22026 7 1 2 92464 22025
0 22027 5 1 1 22026
0 22028 7 1 2 22023 22027
0 22029 5 1 1 22028
0 22030 7 1 2 63964 22029
0 22031 5 1 1 22030
0 22032 7 1 2 63423 22031
0 22033 7 1 2 21997 22032
0 22034 5 1 1 22033
0 22035 7 1 2 80458 91994
0 22036 5 1 1 22035
0 22037 7 1 2 87951 92546
0 22038 5 1 1 22037
0 22039 7 1 2 22036 22038
0 22040 5 1 1 22039
0 22041 7 1 2 59311 22040
0 22042 5 1 1 22041
0 22043 7 1 2 70276 91995
0 22044 5 1 1 22043
0 22045 7 1 2 87888 22044
0 22046 5 1 1 22045
0 22047 7 1 2 59872 22046
0 22048 5 1 1 22047
0 22049 7 1 2 62301 73453
0 22050 5 1 1 22049
0 22051 7 5 2 61517 77554
0 22052 5 1 1 92702
0 22053 7 1 2 82868 92703
0 22054 5 1 1 22053
0 22055 7 1 2 59873 87942
0 22056 5 1 1 22055
0 22057 7 1 2 22054 22056
0 22058 5 1 1 22057
0 22059 7 1 2 22050 22058
0 22060 5 1 1 22059
0 22061 7 1 2 22048 22060
0 22062 7 1 2 22042 22061
0 22063 5 1 1 22062
0 22064 7 1 2 85309 22063
0 22065 5 1 1 22064
0 22066 7 1 2 78055 79375
0 22067 7 1 2 90123 22066
0 22068 5 1 1 22067
0 22069 7 1 2 68333 22068
0 22070 7 1 2 22065 22069
0 22071 5 1 1 22070
0 22072 7 1 2 72106 22071
0 22073 7 1 2 22034 22072
0 22074 5 1 1 22073
0 22075 7 1 2 81219 85991
0 22076 5 1 1 22075
0 22077 7 1 2 75150 7290
0 22078 5 1 1 22077
0 22079 7 1 2 83742 22078
0 22080 5 1 1 22079
0 22081 7 1 2 22076 22080
0 22082 5 1 1 22081
0 22083 7 1 2 80685 22082
0 22084 5 1 1 22083
0 22085 7 2 2 59874 77775
0 22086 5 2 1 92707
0 22087 7 2 2 74783 77316
0 22088 5 1 1 92711
0 22089 7 1 2 61327 22088
0 22090 5 2 1 22089
0 22091 7 1 2 76498 84092
0 22092 5 1 1 22091
0 22093 7 1 2 92713 22092
0 22094 5 1 1 22093
0 22095 7 1 2 77902 22094
0 22096 5 1 1 22095
0 22097 7 1 2 92709 22096
0 22098 5 1 1 22097
0 22099 7 1 2 75301 22098
0 22100 5 1 1 22099
0 22101 7 2 2 67308 77776
0 22102 5 1 1 92715
0 22103 7 1 2 79808 22102
0 22104 5 1 1 22103
0 22105 7 1 2 60339 22104
0 22106 5 1 1 22105
0 22107 7 1 2 73671 77777
0 22108 7 1 2 80246 22107
0 22109 5 1 1 22108
0 22110 7 1 2 22106 22109
0 22111 7 1 2 22100 22110
0 22112 5 1 1 22111
0 22113 7 1 2 61709 22112
0 22114 5 1 1 22113
0 22115 7 1 2 82979 69043
0 22116 7 1 2 80772 22115
0 22117 5 1 1 22116
0 22118 7 1 2 22114 22117
0 22119 5 1 1 22118
0 22120 7 1 2 79134 22119
0 22121 5 1 1 22120
0 22122 7 1 2 22084 22121
0 22123 5 1 1 22122
0 22124 7 1 2 63729 22123
0 22125 5 1 1 22124
0 22126 7 1 2 75437 89772
0 22127 5 1 1 22126
0 22128 7 1 2 20032 22127
0 22129 5 1 1 22128
0 22130 7 1 2 68867 81296
0 22131 7 1 2 85650 22130
0 22132 5 1 1 22131
0 22133 7 1 2 60520 75968
0 22134 5 1 1 22133
0 22135 7 1 2 92197 89745
0 22136 5 1 1 22135
0 22137 7 1 2 22134 22136
0 22138 5 1 1 22137
0 22139 7 1 2 61710 87311
0 22140 7 1 2 22138 22139
0 22141 5 1 1 22140
0 22142 7 1 2 22132 22141
0 22143 5 1 1 22142
0 22144 7 1 2 22129 22143
0 22145 5 1 1 22144
0 22146 7 1 2 60340 74202
0 22147 7 1 2 92466 22146
0 22148 5 1 1 22147
0 22149 7 1 2 92437 22148
0 22150 5 1 1 22149
0 22151 7 1 2 69971 22150
0 22152 5 1 1 22151
0 22153 7 5 2 59524 89096
0 22154 7 1 2 71649 92717
0 22155 5 1 1 22154
0 22156 7 1 2 65404 22155
0 22157 5 1 1 22156
0 22158 7 1 2 69724 79483
0 22159 7 1 2 22157 22158
0 22160 5 1 1 22159
0 22161 7 1 2 22152 22160
0 22162 5 1 1 22161
0 22163 7 1 2 61711 22162
0 22164 5 1 1 22163
0 22165 7 1 2 59875 75943
0 22166 5 1 1 22165
0 22167 7 1 2 62974 22166
0 22168 5 1 1 22167
0 22169 7 1 2 83439 91408
0 22170 7 1 2 22168 22169
0 22171 5 1 1 22170
0 22172 7 1 2 22164 22171
0 22173 5 1 1 22172
0 22174 7 1 2 86493 22173
0 22175 5 1 1 22174
0 22176 7 1 2 22145 22175
0 22177 7 1 2 22125 22176
0 22178 7 1 2 22074 22177
0 22179 7 1 2 21973 22178
0 22180 7 1 2 21922 22179
0 22181 5 1 1 22180
0 22182 7 1 2 86749 22181
0 22183 5 1 1 22182
0 22184 7 1 2 75493 77657
0 22185 7 1 2 92587 22184
0 22186 7 1 2 82162 22185
0 22187 5 1 1 22186
0 22188 7 1 2 22183 22187
0 22189 5 1 1 22188
0 22190 7 1 2 88831 22189
0 22191 5 1 1 22190
0 22192 7 2 2 60341 74862
0 22193 5 1 1 92722
0 22194 7 3 2 78056 79012
0 22195 5 1 1 92724
0 22196 7 2 2 92723 92725
0 22197 5 1 1 92727
0 22198 7 1 2 92025 88644
0 22199 5 1 1 22198
0 22200 7 1 2 20279 22199
0 22201 5 1 1 22200
0 22202 7 1 2 84428 22201
0 22203 5 1 1 22202
0 22204 7 1 2 22197 22203
0 22205 5 1 1 22204
0 22206 7 1 2 61328 22205
0 22207 5 1 1 22206
0 22208 7 1 2 82726 79231
0 22209 5 2 1 22208
0 22210 7 3 2 63730 84599
0 22211 7 1 2 73467 92731
0 22212 5 1 1 22211
0 22213 7 1 2 92729 22212
0 22214 5 1 1 22213
0 22215 7 1 2 80686 22214
0 22216 5 1 1 22215
0 22217 7 1 2 22207 22216
0 22218 5 1 1 22217
0 22219 7 1 2 60133 22218
0 22220 5 1 1 22219
0 22221 7 1 2 92165 92730
0 22222 5 1 1 22221
0 22223 7 1 2 84418 92522
0 22224 7 1 2 22222 22223
0 22225 5 1 1 22224
0 22226 7 1 2 22220 22225
0 22227 5 1 1 22226
0 22228 7 1 2 67609 22227
0 22229 5 1 1 22228
0 22230 7 1 2 92732 89612
0 22231 5 1 1 22230
0 22232 7 1 2 7300 22231
0 22233 5 1 1 22232
0 22234 7 1 2 79135 92512
0 22235 7 1 2 22233 22234
0 22236 5 1 1 22235
0 22237 7 1 2 63424 22236
0 22238 7 1 2 22229 22237
0 22239 5 1 1 22238
0 22240 7 4 2 59525 63965
0 22241 7 9 2 62975 90767
0 22242 7 1 2 71203 92738
0 22243 5 1 1 22242
0 22244 7 2 2 60134 74863
0 22245 7 1 2 67980 92747
0 22246 5 1 1 22245
0 22247 7 1 2 22243 22246
0 22248 5 1 1 22247
0 22249 7 1 2 67610 22248
0 22250 5 1 1 22249
0 22251 7 1 2 89582 22250
0 22252 5 1 1 22251
0 22253 7 1 2 80412 22252
0 22254 5 1 1 22253
0 22255 7 1 2 61052 84380
0 22256 5 1 1 22255
0 22257 7 1 2 71204 77375
0 22258 5 1 1 22257
0 22259 7 1 2 22256 22258
0 22260 5 1 1 22259
0 22261 7 1 2 80181 73761
0 22262 7 1 2 22260 22261
0 22263 5 1 1 22262
0 22264 7 1 2 22254 22263
0 22265 5 1 1 22264
0 22266 7 1 2 68665 22265
0 22267 5 1 1 22266
0 22268 7 6 2 59876 60521
0 22269 7 1 2 92430 92749
0 22270 5 1 1 22269
0 22271 7 1 2 22267 22270
0 22272 5 1 1 22271
0 22273 7 1 2 92734 22272
0 22274 5 1 1 22273
0 22275 7 2 2 75302 70260
0 22276 5 1 1 92755
0 22277 7 1 2 80687 86498
0 22278 7 2 2 92756 22277
0 22279 5 1 1 92757
0 22280 7 1 2 68334 22279
0 22281 7 1 2 22274 22280
0 22282 5 1 1 22281
0 22283 7 1 2 86750 22282
0 22284 7 1 2 22239 22283
0 22285 5 1 1 22284
0 22286 7 1 2 92298 22285
0 22287 5 1 1 22286
0 22288 7 1 2 70530 15672
0 22289 7 1 2 22287 22288
0 22290 5 1 1 22289
0 22291 7 1 2 63425 92697
0 22292 5 1 1 22291
0 22293 7 1 2 81207 22292
0 22294 5 1 1 22293
0 22295 7 1 2 72983 22294
0 22296 5 1 1 22295
0 22297 7 2 2 73015 89252
0 22298 5 1 1 92759
0 22299 7 1 2 89268 92760
0 22300 5 1 1 22299
0 22301 7 1 2 75151 22300
0 22302 5 1 1 22301
0 22303 7 1 2 80951 22302
0 22304 5 1 1 22303
0 22305 7 1 2 22296 22304
0 22306 5 1 1 22305
0 22307 7 1 2 63731 22306
0 22308 5 1 1 22307
0 22309 7 5 2 67611 83535
0 22310 7 1 2 92199 92761
0 22311 5 1 1 22310
0 22312 7 1 2 22308 22311
0 22313 5 1 1 22312
0 22314 7 1 2 59526 22313
0 22315 5 1 1 22314
0 22316 7 1 2 72411 90938
0 22317 5 1 1 22316
0 22318 7 1 2 22315 22317
0 22319 5 1 1 22318
0 22320 7 1 2 87714 22319
0 22321 5 1 1 22320
0 22322 7 12 2 60522 65561
0 22323 7 7 2 61712 85697
0 22324 7 4 2 92766 92778
0 22325 7 1 2 81853 92785
0 22326 7 1 2 89441 22325
0 22327 5 1 1 22326
0 22328 7 1 2 22321 22327
0 22329 5 1 1 22328
0 22330 7 1 2 60915 22329
0 22331 5 1 1 22330
0 22332 7 1 2 89989 88645
0 22333 5 1 1 22332
0 22334 7 1 2 89968 22333
0 22335 5 1 1 22334
0 22336 7 1 2 60135 22335
0 22337 5 1 1 22336
0 22338 7 1 2 12944 89964
0 22339 5 1 1 22338
0 22340 7 1 2 60342 78756
0 22341 7 1 2 83289 22340
0 22342 5 1 1 22341
0 22343 7 1 2 22339 22342
0 22344 7 1 2 22337 22343
0 22345 5 1 1 22344
0 22346 7 1 2 66479 22345
0 22347 5 1 1 22346
0 22348 7 1 2 83290 75066
0 22349 5 1 1 22348
0 22350 7 1 2 20952 22349
0 22351 5 1 1 22350
0 22352 7 1 2 79203 22351
0 22353 5 1 1 22352
0 22354 7 1 2 22347 22353
0 22355 5 1 1 22354
0 22356 7 1 2 67612 22355
0 22357 5 1 1 22356
0 22358 7 1 2 83622 88913
0 22359 5 1 1 22358
0 22360 7 1 2 83671 75772
0 22361 5 1 1 22360
0 22362 7 1 2 22359 22361
0 22363 5 1 1 22362
0 22364 7 1 2 63426 22363
0 22365 5 1 1 22364
0 22366 7 1 2 22357 22365
0 22367 5 1 1 22366
0 22368 7 1 2 87715 22367
0 22369 5 1 1 22368
0 22370 7 6 2 67309 80952
0 22371 7 2 2 63732 79331
0 22372 7 1 2 87716 92795
0 22373 5 1 1 22372
0 22374 7 5 2 66686 79707
0 22375 5 2 1 92797
0 22376 7 1 2 92565 92798
0 22377 5 1 1 22376
0 22378 7 3 2 83374 92103
0 22379 7 1 2 86995 92331
0 22380 7 1 2 92804 22379
0 22381 5 1 1 22380
0 22382 7 1 2 22377 22381
0 22383 5 1 1 22382
0 22384 7 1 2 88618 22383
0 22385 5 1 1 22384
0 22386 7 1 2 22373 22385
0 22387 5 1 1 22386
0 22388 7 1 2 92789 22387
0 22389 5 1 1 22388
0 22390 7 2 2 65405 86751
0 22391 7 1 2 80167 79038
0 22392 7 1 2 73263 22391
0 22393 7 1 2 92807 22392
0 22394 5 1 1 22393
0 22395 7 1 2 22389 22394
0 22396 5 1 1 22395
0 22397 7 1 2 72834 22396
0 22398 5 1 1 22397
0 22399 7 4 2 59527 65562
0 22400 7 3 2 61713 92809
0 22401 7 5 2 60916 80810
0 22402 5 2 1 92816
0 22403 7 4 2 66826 84306
0 22404 7 1 2 92817 92823
0 22405 7 1 2 92813 22404
0 22406 7 1 2 90190 22405
0 22407 5 1 1 22406
0 22408 7 5 2 61053 63427
0 22409 5 1 1 92827
0 22410 7 1 2 87566 22409
0 22411 5 1 1 22410
0 22412 7 1 2 80048 83394
0 22413 7 1 2 22411 22412
0 22414 5 1 1 22413
0 22415 7 1 2 92790 92748
0 22416 5 1 1 22415
0 22417 7 1 2 89478 22416
0 22418 5 1 1 22417
0 22419 7 1 2 74593 22418
0 22420 5 1 1 22419
0 22421 7 1 2 89907 22420
0 22422 7 1 2 22414 22421
0 22423 5 1 1 22422
0 22424 7 3 2 66687 92634
0 22425 7 5 2 63733 86752
0 22426 7 1 2 92832 92835
0 22427 7 1 2 22423 22426
0 22428 5 1 1 22427
0 22429 7 1 2 22407 22428
0 22430 5 1 1 22429
0 22431 7 1 2 69401 22430
0 22432 5 1 1 22431
0 22433 7 1 2 22398 22432
0 22434 7 1 2 22369 22433
0 22435 7 1 2 22331 22434
0 22436 5 1 1 22435
0 22437 7 1 2 68868 22436
0 22438 5 1 1 22437
0 22439 7 1 2 326 72984
0 22440 5 1 1 22439
0 22441 7 1 2 73762 74773
0 22442 5 1 1 22441
0 22443 7 1 2 77188 22442
0 22444 7 1 2 22440 22443
0 22445 5 1 1 22444
0 22446 7 1 2 92576 22445
0 22447 5 1 1 22446
0 22448 7 1 2 60523 91357
0 22449 7 1 2 72430 22448
0 22450 5 1 1 22449
0 22451 7 1 2 22447 22450
0 22452 5 1 1 22451
0 22453 7 6 2 61861 85879
0 22454 7 1 2 83536 92840
0 22455 7 1 2 22452 22454
0 22456 5 1 1 22455
0 22457 7 1 2 22438 22456
0 22458 5 1 1 22457
0 22459 7 1 2 78593 22458
0 22460 5 1 1 22459
0 22461 7 2 2 77555 92405
0 22462 5 1 1 92846
0 22463 7 1 2 60136 92728
0 22464 5 1 1 22463
0 22465 7 1 2 72928 84429
0 22466 7 1 2 92021 22465
0 22467 5 1 1 22466
0 22468 7 1 2 22464 22467
0 22469 5 1 1 22468
0 22470 7 1 2 67613 22469
0 22471 5 1 1 22470
0 22472 7 1 2 22462 22471
0 22473 5 1 1 22472
0 22474 7 1 2 61329 22473
0 22475 5 1 1 22474
0 22476 7 2 2 85513 92638
0 22477 7 1 2 67981 92848
0 22478 7 1 2 89868 22477
0 22479 5 1 1 22478
0 22480 7 1 2 22475 22479
0 22481 5 1 1 22480
0 22482 7 1 2 59528 22481
0 22483 5 1 1 22482
0 22484 7 3 2 62976 92666
0 22485 7 1 2 79559 89650
0 22486 7 1 2 92646 22485
0 22487 7 1 2 92850 22486
0 22488 5 1 1 22487
0 22489 7 1 2 63428 22488
0 22490 7 1 2 22483 22489
0 22491 5 1 1 22490
0 22492 7 1 2 80865 83665
0 22493 5 1 1 22492
0 22494 7 1 2 67614 73504
0 22495 7 1 2 92013 22494
0 22496 5 1 1 22495
0 22497 7 1 2 22493 22496
0 22498 5 1 1 22497
0 22499 7 1 2 75303 22498
0 22500 5 1 1 22499
0 22501 7 1 2 80324 81195
0 22502 5 8 1 22501
0 22503 7 3 2 68666 92853
0 22504 7 1 2 90515 92861
0 22505 5 1 1 22504
0 22506 7 1 2 22500 22505
0 22507 5 1 1 22506
0 22508 7 1 2 62977 22507
0 22509 5 1 1 22508
0 22510 7 1 2 59877 92259
0 22511 5 1 1 22510
0 22512 7 1 2 61518 73731
0 22513 7 1 2 85312 22512
0 22514 5 1 1 22513
0 22515 7 1 2 22511 22514
0 22516 5 1 1 22515
0 22517 7 1 2 85341 22516
0 22518 5 1 1 22517
0 22519 7 1 2 22509 22518
0 22520 5 1 1 22519
0 22521 7 1 2 63966 22520
0 22522 5 1 1 22521
0 22523 7 1 2 59529 92758
0 22524 5 1 1 22523
0 22525 7 1 2 68335 22524
0 22526 7 1 2 22522 22525
0 22527 5 1 1 22526
0 22528 7 1 2 86753 22527
0 22529 7 1 2 22491 22528
0 22530 5 1 1 22529
0 22531 7 8 2 61054 66827
0 22532 7 1 2 73913 92864
0 22533 7 1 2 71406 22532
0 22534 7 1 2 88134 22533
0 22535 7 1 2 92293 22534
0 22536 5 1 1 22535
0 22537 7 1 2 22530 22536
0 22538 5 1 1 22537
0 22539 7 1 2 88687 22538
0 22540 5 1 1 22539
0 22541 7 1 2 77469 92022
0 22542 5 1 1 22541
0 22543 7 1 2 20293 22542
0 22544 5 1 1 22543
0 22545 7 1 2 90626 22544
0 22546 5 1 1 22545
0 22547 7 3 2 62978 77556
0 22548 7 1 2 72740 92639
0 22549 7 1 2 87517 22548
0 22550 7 1 2 92872 22549
0 22551 5 1 1 22550
0 22552 7 1 2 22546 22551
0 22553 5 1 1 22552
0 22554 7 1 2 68336 22553
0 22555 5 1 1 22554
0 22556 7 2 2 78057 92592
0 22557 5 1 1 92875
0 22558 7 1 2 83010 86966
0 22559 7 1 2 92876 22558
0 22560 5 1 1 22559
0 22561 7 1 2 22555 22560
0 22562 5 1 1 22561
0 22563 7 1 2 61055 22562
0 22564 5 1 1 22563
0 22565 7 2 2 61056 78189
0 22566 7 1 2 90768 92877
0 22567 5 1 1 22566
0 22568 7 1 2 89583 22567
0 22569 5 1 1 22568
0 22570 7 1 2 92449 22569
0 22571 5 1 1 22570
0 22572 7 1 2 83666 87805
0 22573 5 1 1 22572
0 22574 7 1 2 82459 83672
0 22575 5 1 1 22574
0 22576 7 1 2 22573 22575
0 22577 5 1 1 22576
0 22578 7 1 2 71872 22577
0 22579 5 1 1 22578
0 22580 7 1 2 22571 22579
0 22581 5 1 1 22580
0 22582 7 1 2 81016 22581
0 22583 5 1 1 22582
0 22584 7 1 2 74931 73732
0 22585 7 1 2 87740 22584
0 22586 5 1 1 22585
0 22587 7 1 2 22583 22586
0 22588 5 1 1 22587
0 22589 7 1 2 81178 22588
0 22590 5 1 1 22589
0 22591 7 1 2 74995 92847
0 22592 5 1 1 22591
0 22593 7 1 2 22590 22592
0 22594 7 1 2 22564 22593
0 22595 5 1 1 22594
0 22596 7 1 2 86754 22595
0 22597 5 1 1 22596
0 22598 7 1 2 92299 22597
0 22599 5 1 1 22598
0 22600 7 1 2 82254 22599
0 22601 5 1 1 22600
0 22602 7 1 2 64089 22601
0 22603 7 1 2 22540 22602
0 22604 7 1 2 22460 22603
0 22605 7 1 2 22290 22604
0 22606 7 1 2 22191 22605
0 22607 7 1 2 21861 22606
0 22608 7 1 2 21638 22607
0 22609 7 1 2 20947 22608
0 22610 7 1 2 19951 22609
0 22611 7 1 2 15536 22610
0 22612 5 1 1 22611
0 22613 7 1 2 12408 22612
0 22614 5 1 1 22613
0 22615 7 1 2 66942 22614
0 22616 5 1 1 22615
0 22617 7 1 2 77632 74768
0 22618 5 1 1 22617
0 22619 7 1 2 72337 90744
0 22620 5 1 1 22619
0 22621 7 1 2 78415 22620
0 22622 5 1 1 22621
0 22623 7 1 2 22618 22622
0 22624 5 1 1 22623
0 22625 7 1 2 67615 22624
0 22626 5 1 1 22625
0 22627 7 1 2 91934 22626
0 22628 5 1 1 22627
0 22629 7 1 2 77646 22628
0 22630 5 1 1 22629
0 22631 7 1 2 59312 73931
0 22632 5 1 1 22631
0 22633 7 1 2 76008 22632
0 22634 5 1 1 22633
0 22635 7 1 2 69447 22634
0 22636 5 1 1 22635
0 22637 7 1 2 70399 72473
0 22638 5 1 1 22637
0 22639 7 1 2 1401 22638
0 22640 7 1 2 22636 22639
0 22641 5 1 1 22640
0 22642 7 1 2 72929 22641
0 22643 5 1 1 22642
0 22644 7 1 2 71979 76091
0 22645 5 2 1 22644
0 22646 7 1 2 60137 92879
0 22647 5 1 1 22646
0 22648 7 1 2 70400 89550
0 22649 5 1 1 22648
0 22650 7 1 2 22647 22649
0 22651 5 1 1 22650
0 22652 7 1 2 71205 22651
0 22653 5 1 1 22652
0 22654 7 1 2 72972 22653
0 22655 7 1 2 22643 22654
0 22656 7 1 2 22630 22655
0 22657 5 1 1 22656
0 22658 7 1 2 63429 22657
0 22659 5 1 1 22658
0 22660 7 5 2 68337 72592
0 22661 7 3 2 80597 92881
0 22662 7 1 2 84111 92886
0 22663 5 1 1 22662
0 22664 7 1 2 22659 22663
0 22665 5 1 1 22664
0 22666 7 1 2 61519 22665
0 22667 5 1 1 22666
0 22668 7 1 2 72930 89902
0 22669 5 1 1 22668
0 22670 7 1 2 89551 88635
0 22671 5 1 1 22670
0 22672 7 1 2 22669 22671
0 22673 5 1 1 22672
0 22674 7 1 2 59313 75834
0 22675 5 1 1 22674
0 22676 7 1 2 83413 22675
0 22677 5 1 1 22676
0 22678 7 1 2 22673 22677
0 22679 5 1 1 22678
0 22680 7 3 2 61057 75835
0 22681 5 1 1 92889
0 22682 7 1 2 4089 22681
0 22683 5 1 1 22682
0 22684 7 1 2 60138 22683
0 22685 5 1 1 22684
0 22686 7 2 2 60343 73318
0 22687 7 1 2 63430 92892
0 22688 5 1 1 22687
0 22689 7 1 2 75862 22688
0 22690 5 1 1 22689
0 22691 7 1 2 59878 22690
0 22692 5 1 1 22691
0 22693 7 1 2 22685 22692
0 22694 5 1 1 22693
0 22695 7 1 2 59530 22694
0 22696 5 1 1 22695
0 22697 7 2 2 60917 75836
0 22698 5 1 1 92894
0 22699 7 1 2 83414 22698
0 22700 5 1 1 22699
0 22701 7 1 2 72674 22700
0 22702 5 1 1 22701
0 22703 7 1 2 22696 22702
0 22704 5 1 1 22703
0 22705 7 1 2 59314 22704
0 22706 5 1 1 22705
0 22707 7 1 2 22679 22706
0 22708 5 1 1 22707
0 22709 7 1 2 69402 22708
0 22710 5 1 1 22709
0 22711 7 1 2 73131 83436
0 22712 5 1 1 22711
0 22713 7 1 2 83186 83303
0 22714 5 1 1 22713
0 22715 7 1 2 22712 22714
0 22716 5 1 1 22715
0 22717 7 1 2 67616 22716
0 22718 5 1 1 22717
0 22719 7 1 2 75863 22718
0 22720 5 1 1 22719
0 22721 7 1 2 59879 22720
0 22722 5 1 1 22721
0 22723 7 1 2 83415 84755
0 22724 5 2 1 22723
0 22725 7 4 2 59315 63431
0 22726 7 1 2 71666 92898
0 22727 5 1 1 22726
0 22728 7 1 2 64499 22727
0 22729 5 1 1 22728
0 22730 7 1 2 92896 22729
0 22731 5 1 1 22730
0 22732 7 1 2 81208 22731
0 22733 5 1 1 22732
0 22734 7 1 2 60139 22733
0 22735 5 1 1 22734
0 22736 7 1 2 22722 22735
0 22737 5 1 1 22736
0 22738 7 1 2 88779 22737
0 22739 5 1 1 22738
0 22740 7 1 2 73132 81203
0 22741 5 1 1 22740
0 22742 7 1 2 59316 83420
0 22743 5 1 1 22742
0 22744 7 1 2 22741 22743
0 22745 5 1 1 22744
0 22746 7 1 2 72931 22745
0 22747 5 1 1 22746
0 22748 7 1 2 60140 92897
0 22749 5 1 1 22748
0 22750 7 1 2 83404 83366
0 22751 5 1 1 22750
0 22752 7 1 2 75864 22751
0 22753 5 1 1 22752
0 22754 7 1 2 59531 22753
0 22755 5 1 1 22754
0 22756 7 1 2 22749 22755
0 22757 5 1 1 22756
0 22758 7 1 2 71206 22757
0 22759 5 1 1 22758
0 22760 7 1 2 22747 22759
0 22761 5 1 1 22760
0 22762 7 1 2 72835 22761
0 22763 5 1 1 22762
0 22764 7 1 2 72719 72168
0 22765 5 1 1 22764
0 22766 7 1 2 91949 22765
0 22767 5 1 1 22766
0 22768 7 1 2 72969 22767
0 22769 5 1 1 22768
0 22770 7 1 2 83405 22769
0 22771 5 1 1 22770
0 22772 7 1 2 91271 89253
0 22773 5 1 1 22772
0 22774 7 1 2 65193 22773
0 22775 5 1 1 22774
0 22776 7 1 2 75837 22775
0 22777 5 1 1 22776
0 22778 7 2 2 61058 80073
0 22779 5 1 1 92902
0 22780 7 1 2 64959 22779
0 22781 5 1 1 22780
0 22782 7 1 2 59532 75838
0 22783 5 1 1 22782
0 22784 7 1 2 6735 22783
0 22785 5 1 1 22784
0 22786 7 1 2 82487 22785
0 22787 5 1 1 22786
0 22788 7 1 2 82484 90053
0 22789 5 1 1 22788
0 22790 7 1 2 59880 81204
0 22791 5 1 1 22790
0 22792 7 1 2 22789 22791
0 22793 7 1 2 22787 22792
0 22794 5 1 1 22793
0 22795 7 1 2 22781 22794
0 22796 5 1 1 22795
0 22797 7 1 2 22777 22796
0 22798 7 1 2 22771 22797
0 22799 7 1 2 22763 22798
0 22800 7 1 2 22739 22799
0 22801 7 1 2 22710 22800
0 22802 7 1 2 22667 22801
0 22803 5 1 1 22802
0 22804 7 1 2 63734 22803
0 22805 5 1 1 22804
0 22806 7 4 2 64718 70448
0 22807 7 2 2 90445 92904
0 22808 5 1 1 92908
0 22809 7 1 2 90939 22808
0 22810 5 1 1 22809
0 22811 7 2 2 83537 78991
0 22812 5 1 1 92910
0 22813 7 1 2 77023 92911
0 22814 5 1 1 22813
0 22815 7 1 2 74466 91944
0 22816 5 1 1 22815
0 22817 7 1 2 22814 22816
0 22818 5 1 1 22817
0 22819 7 1 2 64719 22818
0 22820 5 1 1 22819
0 22821 7 1 2 22810 22820
0 22822 7 1 2 22805 22821
0 22823 5 1 1 22822
0 22824 7 1 2 61330 22823
0 22825 5 1 1 22824
0 22826 7 2 2 59317 76043
0 22827 5 2 1 92912
0 22828 7 2 2 89399 92913
0 22829 5 1 1 92916
0 22830 7 1 2 75839 73284
0 22831 5 1 1 22830
0 22832 7 1 2 22829 22831
0 22833 5 1 1 22832
0 22834 7 1 2 74894 22833
0 22835 5 1 1 22834
0 22836 7 1 2 59881 89410
0 22837 5 1 1 22836
0 22838 7 1 2 22835 22837
0 22839 5 1 1 22838
0 22840 7 1 2 67310 22839
0 22841 5 1 1 22840
0 22842 7 2 2 76560 73434
0 22843 5 2 1 92918
0 22844 7 1 2 89400 92919
0 22845 5 1 1 22844
0 22846 7 1 2 22841 22845
0 22847 5 1 1 22846
0 22848 7 1 2 61059 22847
0 22849 5 1 1 22848
0 22850 7 3 2 77117 73190
0 22851 5 2 1 92922
0 22852 7 1 2 89411 92923
0 22853 5 1 1 22852
0 22854 7 1 2 22849 22853
0 22855 5 1 1 22854
0 22856 7 1 2 60918 22855
0 22857 5 1 1 22856
0 22858 7 1 2 89486 91497
0 22859 5 1 1 22858
0 22860 7 1 2 75566 22859
0 22861 5 1 1 22860
0 22862 7 1 2 63432 22861
0 22863 5 1 1 22862
0 22864 7 1 2 22857 22863
0 22865 5 1 1 22864
0 22866 7 1 2 60141 22865
0 22867 5 1 1 22866
0 22868 7 1 2 59882 73340
0 22869 5 1 1 22868
0 22870 7 1 2 73763 75749
0 22871 5 1 1 22870
0 22872 7 1 2 22869 22871
0 22873 5 1 1 22872
0 22874 7 1 2 59533 22873
0 22875 5 1 1 22874
0 22876 7 1 2 81566 73987
0 22877 5 1 1 22876
0 22878 7 1 2 60344 22877
0 22879 5 1 1 22878
0 22880 7 1 2 73993 91506
0 22881 5 1 1 22880
0 22882 7 1 2 22879 22881
0 22883 7 1 2 22875 22882
0 22884 5 1 1 22883
0 22885 7 1 2 66480 22884
0 22886 5 1 1 22885
0 22887 7 1 2 81881 73988
0 22888 5 1 1 22887
0 22889 7 1 2 81062 22888
0 22890 5 1 1 22889
0 22891 7 1 2 22886 22890
0 22892 5 1 1 22891
0 22893 7 1 2 61520 73264
0 22894 5 1 1 22893
0 22895 7 1 2 63433 22894
0 22896 7 1 2 14672 22895
0 22897 5 1 1 22896
0 22898 7 2 2 59318 22897
0 22899 5 1 1 92927
0 22900 7 1 2 22892 92928
0 22901 5 1 1 22900
0 22902 7 1 2 74594 91517
0 22903 5 1 1 22902
0 22904 7 1 2 75567 83392
0 22905 5 1 1 22904
0 22906 7 1 2 75304 73816
0 22907 7 1 2 22905 22906
0 22908 5 1 1 22907
0 22909 7 1 2 22903 22908
0 22910 5 1 1 22909
0 22911 7 1 2 67311 22910
0 22912 5 1 1 22911
0 22913 7 1 2 75998 89661
0 22914 5 1 1 22913
0 22915 7 1 2 22899 22914
0 22916 7 1 2 22912 22915
0 22917 5 1 1 22916
0 22918 7 1 2 63434 22917
0 22919 5 1 1 22918
0 22920 7 1 2 22901 22919
0 22921 5 1 1 22920
0 22922 7 1 2 69403 22921
0 22923 5 1 1 22922
0 22924 7 1 2 80801 89412
0 22925 5 1 1 22924
0 22926 7 1 2 20154 22925
0 22927 5 2 1 22926
0 22928 7 1 2 71207 92929
0 22929 5 1 1 22928
0 22930 7 1 2 81205 72960
0 22931 5 1 1 22930
0 22932 7 1 2 22929 22931
0 22933 5 1 1 22932
0 22934 7 1 2 70277 22933
0 22935 5 1 1 22934
0 22936 7 1 2 59534 89417
0 22937 5 1 1 22936
0 22938 7 1 2 22935 22937
0 22939 5 1 1 22938
0 22940 7 1 2 69113 22939
0 22941 5 1 1 22940
0 22942 7 1 2 83604 76065
0 22943 5 2 1 22942
0 22944 7 1 2 76997 92931
0 22945 5 1 1 22944
0 22946 7 1 2 62635 22945
0 22947 5 1 1 22946
0 22948 7 1 2 59319 74164
0 22949 5 1 1 22948
0 22950 7 1 2 64720 22949
0 22951 5 1 1 22950
0 22952 7 1 2 22947 22951
0 22953 5 1 1 22952
0 22954 7 1 2 66015 22953
0 22955 5 1 1 22954
0 22956 7 1 2 80146 82208
0 22957 7 1 2 22955 22956
0 22958 5 1 1 22957
0 22959 7 1 2 59883 92930
0 22960 5 1 1 22959
0 22961 7 1 2 67617 89471
0 22962 5 1 1 22961
0 22963 7 1 2 22960 22962
0 22964 5 1 1 22963
0 22965 7 1 2 71598 22964
0 22966 5 1 1 22965
0 22967 7 1 2 74864 91507
0 22968 5 1 1 22967
0 22969 7 1 2 17116 22968
0 22970 5 1 1 22969
0 22971 7 1 2 83187 22970
0 22972 5 1 1 22971
0 22973 7 1 2 59320 89418
0 22974 5 1 1 22973
0 22975 7 1 2 22972 22974
0 22976 5 1 1 22975
0 22977 7 1 2 70419 22976
0 22978 5 1 1 22977
0 22979 7 1 2 80811 90833
0 22980 5 1 1 22979
0 22981 7 1 2 89468 22980
0 22982 5 1 1 22981
0 22983 7 1 2 60919 22982
0 22984 5 1 1 22983
0 22985 7 1 2 83375 89884
0 22986 5 1 1 22985
0 22987 7 1 2 22984 22986
0 22988 5 1 1 22987
0 22989 7 1 2 90470 22988
0 22990 5 1 1 22989
0 22991 7 1 2 22978 22990
0 22992 7 1 2 22966 22991
0 22993 7 1 2 22958 22992
0 22994 7 1 2 22941 22993
0 22995 7 1 2 22923 22994
0 22996 7 1 2 22867 22995
0 22997 5 1 1 22996
0 22998 7 1 2 63735 22997
0 22999 5 1 1 22998
0 23000 7 1 2 66016 82478
0 23001 5 3 1 23000
0 23002 7 1 2 72154 92933
0 23003 5 1 1 23002
0 23004 7 1 2 74099 74622
0 23005 5 1 1 23004
0 23006 7 1 2 23003 23005
0 23007 5 1 1 23006
0 23008 7 1 2 69906 23007
0 23009 5 1 1 23008
0 23010 7 1 2 67618 88723
0 23011 5 1 1 23010
0 23012 7 1 2 79985 23011
0 23013 5 1 1 23012
0 23014 7 1 2 71208 23013
0 23015 5 1 1 23014
0 23016 7 1 2 76206 72932
0 23017 5 3 1 23016
0 23018 7 1 2 67619 75818
0 23019 5 1 1 23018
0 23020 7 1 2 92936 23019
0 23021 7 1 2 23015 23020
0 23022 7 1 2 23009 23021
0 23023 5 1 1 23022
0 23024 7 1 2 66481 23023
0 23025 5 1 1 23024
0 23026 7 1 2 74857 23025
0 23027 5 1 1 23026
0 23028 7 1 2 65194 23027
0 23029 5 1 1 23028
0 23030 7 1 2 59535 83316
0 23031 5 1 1 23030
0 23032 7 1 2 64960 23031
0 23033 5 1 1 23032
0 23034 7 1 2 62095 23033
0 23035 5 1 1 23034
0 23036 7 1 2 76461 13001
0 23037 5 1 1 23036
0 23038 7 1 2 59321 23037
0 23039 5 1 1 23038
0 23040 7 1 2 23035 23039
0 23041 5 1 1 23040
0 23042 7 1 2 71209 23041
0 23043 5 1 1 23042
0 23044 7 1 2 74470 90829
0 23045 5 1 1 23044
0 23046 7 1 2 66482 23045
0 23047 7 1 2 23043 23046
0 23048 5 1 1 23047
0 23049 7 3 2 73566 69983
0 23050 7 1 2 77856 92939
0 23051 5 1 1 23050
0 23052 7 1 2 61521 90346
0 23053 7 1 2 23051 23052
0 23054 5 1 1 23053
0 23055 7 1 2 62636 23054
0 23056 7 1 2 23048 23055
0 23057 5 1 1 23056
0 23058 7 1 2 77293 86411
0 23059 7 1 2 82582 23058
0 23060 5 1 1 23059
0 23061 7 1 2 23057 23060
0 23062 5 1 1 23061
0 23063 7 1 2 66256 23062
0 23064 5 1 1 23063
0 23065 7 1 2 63435 23064
0 23066 7 1 2 23029 23065
0 23067 5 1 1 23066
0 23068 7 1 2 71980 80239
0 23069 5 1 1 23068
0 23070 7 1 2 74460 82142
0 23071 7 1 2 88410 23070
0 23072 5 1 1 23071
0 23073 7 1 2 62096 23072
0 23074 5 1 1 23073
0 23075 7 1 2 23069 23074
0 23076 5 1 1 23075
0 23077 7 1 2 75202 23076
0 23078 5 1 1 23077
0 23079 7 1 2 76967 82735
0 23080 5 1 1 23079
0 23081 7 1 2 76181 23080
0 23082 5 1 1 23081
0 23083 7 1 2 82078 82736
0 23084 5 1 1 23083
0 23085 7 1 2 73868 23084
0 23086 5 1 1 23085
0 23087 7 1 2 23082 23086
0 23088 5 1 1 23087
0 23089 7 1 2 66017 83459
0 23090 7 1 2 23088 23089
0 23091 5 1 1 23090
0 23092 7 1 2 23078 23091
0 23093 5 1 1 23092
0 23094 7 1 2 66257 23093
0 23095 5 1 1 23094
0 23096 7 2 2 62637 75203
0 23097 7 3 2 77857 92942
0 23098 5 1 1 92944
0 23099 7 1 2 68338 23098
0 23100 7 1 2 23095 23099
0 23101 5 1 1 23100
0 23102 7 1 2 68667 23101
0 23103 7 1 2 23067 23102
0 23104 5 1 1 23103
0 23105 7 1 2 22999 23104
0 23106 7 1 2 22825 23105
0 23107 5 1 1 23106
0 23108 7 1 2 68869 23107
0 23109 5 1 1 23108
0 23110 7 2 2 75494 89926
0 23111 7 1 2 70993 92947
0 23112 5 1 1 23111
0 23113 7 1 2 23109 23112
0 23114 5 1 1 23113
0 23115 7 1 2 65406 23114
0 23116 5 1 1 23115
0 23117 7 2 2 66258 87943
0 23118 7 1 2 80115 92949
0 23119 5 1 1 23118
0 23120 7 2 2 64500 86412
0 23121 7 1 2 80730 77557
0 23122 7 1 2 92951 23121
0 23123 5 1 1 23122
0 23124 7 1 2 23119 23123
0 23125 5 1 1 23124
0 23126 7 1 2 69803 23125
0 23127 5 1 1 23126
0 23128 7 7 2 61522 68668
0 23129 5 1 1 92953
0 23130 7 1 2 82107 92954
0 23131 5 1 1 23130
0 23132 7 1 2 64279 83318
0 23133 5 1 1 23132
0 23134 7 1 2 59536 69355
0 23135 7 1 2 23133 23134
0 23136 5 1 1 23135
0 23137 7 1 2 81877 23136
0 23138 5 2 1 23137
0 23139 7 1 2 83667 89106
0 23140 7 1 2 92960 23139
0 23141 5 1 1 23140
0 23142 7 1 2 23131 23141
0 23143 5 1 1 23142
0 23144 7 1 2 81017 23143
0 23145 5 1 1 23144
0 23146 7 1 2 23127 23145
0 23147 5 1 1 23146
0 23148 7 1 2 67065 23147
0 23149 5 1 1 23148
0 23150 7 4 2 68339 87853
0 23151 7 1 2 73715 91026
0 23152 7 1 2 92962 23151
0 23153 7 1 2 71446 23152
0 23154 5 1 1 23153
0 23155 7 1 2 23149 23154
0 23156 5 1 1 23155
0 23157 7 1 2 67620 23156
0 23158 5 1 1 23157
0 23159 7 2 2 68669 81094
0 23160 7 1 2 79916 75983
0 23161 7 1 2 92966 23160
0 23162 7 1 2 70911 23161
0 23163 5 1 1 23162
0 23164 7 1 2 23158 23163
0 23165 5 1 1 23164
0 23166 7 1 2 60524 23165
0 23167 5 1 1 23166
0 23168 7 1 2 86494 91478
0 23169 7 1 2 71330 23168
0 23170 7 1 2 71447 23169
0 23171 5 1 1 23170
0 23172 7 1 2 23167 23171
0 23173 7 1 2 23116 23172
0 23174 5 1 1 23173
0 23175 7 1 2 67982 23174
0 23176 5 1 1 23175
0 23177 7 1 2 88770 91950
0 23178 5 1 1 23177
0 23179 7 1 2 71210 76257
0 23180 7 1 2 89160 23179
0 23181 7 1 2 89552 23180
0 23182 5 1 1 23181
0 23183 7 1 2 23178 23182
0 23184 5 1 1 23183
0 23185 7 1 2 67312 23184
0 23186 5 1 1 23185
0 23187 7 1 2 69307 88794
0 23188 5 1 1 23187
0 23189 7 1 2 81587 91951
0 23190 5 1 1 23189
0 23191 7 1 2 23188 23190
0 23192 7 1 2 23186 23191
0 23193 5 1 1 23192
0 23194 7 1 2 67066 23193
0 23195 5 1 1 23194
0 23196 7 1 2 72569 72933
0 23197 5 1 1 23196
0 23198 7 1 2 72720 23197
0 23199 5 1 1 23198
0 23200 7 1 2 69114 23199
0 23201 5 1 1 23200
0 23202 7 1 2 60142 85791
0 23203 5 1 1 23202
0 23204 7 1 2 13680 23203
0 23205 5 1 1 23204
0 23206 7 1 2 78630 23205
0 23207 5 1 1 23206
0 23208 7 1 2 23201 23207
0 23209 5 1 1 23208
0 23210 7 1 2 67621 23209
0 23211 5 1 1 23210
0 23212 7 1 2 23195 23211
0 23213 5 1 1 23212
0 23214 7 1 2 66483 23213
0 23215 5 1 1 23214
0 23216 7 2 2 67622 74848
0 23217 5 1 1 92968
0 23218 7 1 2 77076 92969
0 23219 5 1 1 23218
0 23220 7 1 2 75568 76207
0 23221 7 1 2 89289 23220
0 23222 5 1 1 23221
0 23223 7 1 2 23219 23222
0 23224 7 1 2 23215 23223
0 23225 5 1 1 23224
0 23226 7 1 2 66259 23225
0 23227 5 1 1 23226
0 23228 7 1 2 72570 71211
0 23229 5 1 1 23228
0 23230 7 2 2 72338 23229
0 23231 5 2 1 92970
0 23232 7 1 2 69115 92972
0 23233 5 1 1 23232
0 23234 7 1 2 70984 90361
0 23235 5 1 1 23234
0 23236 7 1 2 81367 23235
0 23237 7 1 2 23233 23236
0 23238 5 1 1 23237
0 23239 7 1 2 70164 23238
0 23240 5 1 1 23239
0 23241 7 1 2 70606 72732
0 23242 5 1 1 23241
0 23243 7 1 2 60345 78039
0 23244 5 1 1 23243
0 23245 7 1 2 62097 23244
0 23246 7 1 2 23242 23245
0 23247 7 1 2 23240 23246
0 23248 5 1 1 23247
0 23249 7 1 2 67067 11184
0 23250 5 1 1 23249
0 23251 7 1 2 74932 23250
0 23252 7 1 2 23248 23251
0 23253 5 1 1 23252
0 23254 7 1 2 74852 79165
0 23255 5 1 1 23254
0 23256 7 1 2 70165 92058
0 23257 7 1 2 74748 23256
0 23258 5 1 1 23257
0 23259 7 1 2 23255 23258
0 23260 5 1 1 23259
0 23261 7 1 2 62302 23260
0 23262 5 1 1 23261
0 23263 7 1 2 65852 90352
0 23264 5 1 1 23263
0 23265 7 1 2 1992 23264
0 23266 5 1 1 23265
0 23267 7 1 2 85154 23266
0 23268 5 1 1 23267
0 23269 7 1 2 23262 23268
0 23270 7 1 2 23253 23269
0 23271 7 1 2 23227 23270
0 23272 5 1 1 23271
0 23273 7 1 2 83538 23272
0 23274 5 1 1 23273
0 23275 7 1 2 62303 76926
0 23276 5 3 1 23275
0 23277 7 1 2 76516 4460
0 23278 7 1 2 92974 23277
0 23279 5 1 1 23278
0 23280 7 1 2 62638 23279
0 23281 5 1 1 23280
0 23282 7 1 2 73143 74480
0 23283 5 1 1 23282
0 23284 7 1 2 78452 8647
0 23285 5 1 1 23284
0 23286 7 1 2 23283 23285
0 23287 7 1 2 23281 23286
0 23288 5 1 1 23287
0 23289 7 1 2 66484 23288
0 23290 5 1 1 23289
0 23291 7 1 2 72548 74121
0 23292 7 1 2 87985 23291
0 23293 5 1 1 23292
0 23294 7 2 2 73749 23293
0 23295 7 1 2 83327 85052
0 23296 5 1 1 23295
0 23297 7 1 2 92977 23296
0 23298 5 1 1 23297
0 23299 7 1 2 77160 23298
0 23300 5 1 1 23299
0 23301 7 1 2 23290 23300
0 23302 5 1 1 23301
0 23303 7 1 2 65195 23302
0 23304 5 1 1 23303
0 23305 7 1 2 83328 78040
0 23306 5 1 1 23305
0 23307 7 1 2 92978 23306
0 23308 5 1 1 23307
0 23309 7 1 2 85272 23308
0 23310 5 1 1 23309
0 23311 7 1 2 68670 23310
0 23312 7 1 2 23304 23311
0 23313 5 1 1 23312
0 23314 7 1 2 90462 88727
0 23315 5 1 1 23314
0 23316 7 8 2 61060 75305
0 23317 7 1 2 59884 92979
0 23318 5 1 1 23317
0 23319 7 1 2 23315 23318
0 23320 5 1 1 23319
0 23321 7 1 2 61331 23320
0 23322 5 1 1 23321
0 23323 7 1 2 73414 92980
0 23324 5 1 1 23323
0 23325 7 1 2 23322 23324
0 23326 5 1 1 23325
0 23327 7 1 2 62639 23326
0 23328 5 1 1 23327
0 23329 7 1 2 81847 75948
0 23330 5 1 1 23329
0 23331 7 1 2 75306 73634
0 23332 7 1 2 23330 23331
0 23333 5 1 1 23332
0 23334 7 1 2 78322 88211
0 23335 5 1 1 23334
0 23336 7 1 2 89597 89737
0 23337 5 1 1 23336
0 23338 7 1 2 90570 91066
0 23339 5 1 1 23338
0 23340 7 1 2 23337 23339
0 23341 5 1 1 23340
0 23342 7 1 2 69907 23341
0 23343 5 1 1 23342
0 23344 7 1 2 23335 23343
0 23345 7 1 2 23333 23344
0 23346 5 1 1 23345
0 23347 7 1 2 71212 23346
0 23348 5 1 1 23347
0 23349 7 1 2 78334 89487
0 23350 5 1 1 23349
0 23351 7 1 2 81819 74366
0 23352 5 1 1 23351
0 23353 7 1 2 23350 23352
0 23354 5 1 1 23353
0 23355 7 1 2 67313 23354
0 23356 5 1 1 23355
0 23357 7 1 2 72187 90574
0 23358 5 1 1 23357
0 23359 7 1 2 78460 88212
0 23360 5 1 1 23359
0 23361 7 1 2 74044 90571
0 23362 5 1 1 23361
0 23363 7 1 2 23360 23362
0 23364 5 1 1 23363
0 23365 7 1 2 69908 23364
0 23366 5 1 1 23365
0 23367 7 1 2 23358 23366
0 23368 7 1 2 23356 23367
0 23369 5 1 1 23368
0 23370 7 1 2 72934 23369
0 23371 5 1 1 23370
0 23372 7 2 2 62640 73672
0 23373 7 1 2 77208 92987
0 23374 7 1 2 90463 23373
0 23375 5 1 1 23374
0 23376 7 1 2 75495 81857
0 23377 5 1 1 23376
0 23378 7 1 2 63736 23377
0 23379 7 1 2 23375 23378
0 23380 7 1 2 23371 23379
0 23381 7 1 2 23348 23380
0 23382 7 1 2 23328 23381
0 23383 5 1 1 23382
0 23384 7 1 2 68340 23383
0 23385 7 1 2 23313 23384
0 23386 5 1 1 23385
0 23387 7 1 2 23274 23386
0 23388 5 1 1 23387
0 23389 7 1 2 62979 23388
0 23390 5 1 1 23389
0 23391 7 1 2 59537 89039
0 23392 5 1 1 23391
0 23393 7 1 2 91144 23392
0 23394 5 1 1 23393
0 23395 7 1 2 59885 23394
0 23396 5 1 1 23395
0 23397 7 1 2 72188 88847
0 23398 5 1 1 23397
0 23399 7 1 2 70053 90498
0 23400 5 1 1 23399
0 23401 7 1 2 81694 23400
0 23402 5 1 1 23401
0 23403 7 1 2 23398 23402
0 23404 5 1 1 23403
0 23405 7 1 2 71487 23404
0 23406 5 1 1 23405
0 23407 7 1 2 87957 91245
0 23408 5 1 1 23407
0 23409 7 1 2 59538 89084
0 23410 5 1 1 23409
0 23411 7 1 2 73817 90862
0 23412 5 2 1 23411
0 23413 7 1 2 81567 92989
0 23414 7 1 2 23410 23413
0 23415 5 1 1 23414
0 23416 7 1 2 70166 23415
0 23417 5 1 1 23416
0 23418 7 1 2 23408 23417
0 23419 7 1 2 23406 23418
0 23420 7 1 2 23396 23419
0 23421 5 1 1 23420
0 23422 7 1 2 63436 23421
0 23423 5 1 1 23422
0 23424 7 1 2 61061 81855
0 23425 5 1 1 23424
0 23426 7 1 2 77605 23425
0 23427 5 1 1 23426
0 23428 7 1 2 23423 23427
0 23429 5 1 1 23428
0 23430 7 1 2 61523 23429
0 23431 5 1 1 23430
0 23432 7 1 2 75840 71331
0 23433 5 1 1 23432
0 23434 7 1 2 80671 23433
0 23435 5 1 1 23434
0 23436 7 1 2 71719 23435
0 23437 5 1 1 23436
0 23438 7 3 2 60143 69909
0 23439 5 1 1 92991
0 23440 7 1 2 79917 75714
0 23441 7 1 2 92992 23440
0 23442 5 1 1 23441
0 23443 7 1 2 23437 23442
0 23444 5 1 1 23443
0 23445 7 1 2 67314 23444
0 23446 5 1 1 23445
0 23447 7 1 2 75865 23446
0 23448 5 1 1 23447
0 23449 7 1 2 71213 23448
0 23450 5 1 1 23449
0 23451 7 2 2 80930 77658
0 23452 5 1 1 92994
0 23453 7 1 2 92828 92995
0 23454 5 1 1 23453
0 23455 7 2 2 78489 78467
0 23456 5 1 1 92996
0 23457 7 1 2 75841 72935
0 23458 7 1 2 23456 23457
0 23459 5 1 1 23458
0 23460 7 1 2 23454 23459
0 23461 7 1 2 23450 23460
0 23462 5 1 1 23461
0 23463 7 1 2 67623 23462
0 23464 5 1 1 23463
0 23465 7 1 2 23431 23464
0 23466 5 1 1 23465
0 23467 7 1 2 60346 23466
0 23468 5 1 1 23467
0 23469 7 1 2 79771 72189
0 23470 5 1 1 23469
0 23471 7 1 2 75842 74045
0 23472 5 1 1 23471
0 23473 7 1 2 23470 23472
0 23474 5 1 1 23473
0 23475 7 1 2 71488 23474
0 23476 5 1 1 23475
0 23477 7 1 2 79772 75798
0 23478 5 1 1 23477
0 23479 7 1 2 23476 23478
0 23480 5 1 1 23479
0 23481 7 1 2 71214 23480
0 23482 5 1 1 23481
0 23483 7 1 2 75843 80613
0 23484 5 1 1 23483
0 23485 7 1 2 81509 89466
0 23486 5 1 1 23485
0 23487 7 1 2 89885 23486
0 23488 7 1 2 23484 23487
0 23489 5 1 1 23488
0 23490 7 1 2 72225 23489
0 23491 5 1 1 23490
0 23492 7 1 2 23482 23491
0 23493 5 1 1 23492
0 23494 7 1 2 67624 23493
0 23495 5 1 1 23494
0 23496 7 1 2 75725 92829
0 23497 7 1 2 82440 23496
0 23498 5 1 1 23497
0 23499 7 1 2 23495 23498
0 23500 5 1 1 23499
0 23501 7 1 2 70607 23500
0 23502 5 1 1 23501
0 23503 7 1 2 23468 23502
0 23504 5 1 1 23503
0 23505 7 1 2 63737 23504
0 23506 5 1 1 23505
0 23507 7 1 2 67625 4254
0 23508 5 1 1 23507
0 23509 7 1 2 82298 74623
0 23510 5 1 1 23509
0 23511 7 1 2 74769 76539
0 23512 5 1 1 23511
0 23513 7 1 2 92937 23512
0 23514 7 1 2 23510 23513
0 23515 7 1 2 23508 23514
0 23516 5 1 1 23515
0 23517 7 1 2 72820 84865
0 23518 7 1 2 23516 23517
0 23519 5 1 1 23518
0 23520 7 1 2 23506 23519
0 23521 7 1 2 23390 23520
0 23522 5 1 1 23521
0 23523 7 1 2 65407 23522
0 23524 5 1 1 23523
0 23525 7 1 2 71288 75776
0 23526 5 1 1 23525
0 23527 7 1 2 78657 23526
0 23528 5 2 1 23527
0 23529 7 1 2 62304 92998
0 23530 5 1 1 23529
0 23531 7 1 2 84711 88979
0 23532 5 1 1 23531
0 23533 7 1 2 23530 23532
0 23534 5 2 1 23533
0 23535 7 1 2 67626 93000
0 23536 5 1 1 23535
0 23537 7 1 2 74149 74081
0 23538 5 1 1 23537
0 23539 7 2 2 74150 82652
0 23540 5 1 1 93002
0 23541 7 2 2 60798 74122
0 23542 7 1 2 90872 93004
0 23543 5 1 1 23542
0 23544 7 1 2 23540 23543
0 23545 5 1 1 23544
0 23546 7 1 2 59322 23545
0 23547 5 1 1 23546
0 23548 7 1 2 76603 89126
0 23549 5 1 1 23548
0 23550 7 1 2 23547 23549
0 23551 5 1 1 23550
0 23552 7 1 2 72190 23551
0 23553 5 1 1 23552
0 23554 7 1 2 23538 23553
0 23555 7 1 2 23536 23554
0 23556 5 1 1 23555
0 23557 7 1 2 82037 88271
0 23558 7 1 2 23556 23557
0 23559 5 1 1 23558
0 23560 7 1 2 23524 23559
0 23561 5 1 1 23560
0 23562 7 1 2 68870 23561
0 23563 5 1 1 23562
0 23564 7 2 2 76344 88991
0 23565 5 1 1 93006
0 23566 7 1 2 76595 93007
0 23567 5 1 1 23566
0 23568 7 1 2 60920 82322
0 23569 5 2 1 23568
0 23570 7 1 2 89237 93008
0 23571 5 1 1 23570
0 23572 7 1 2 59539 23571
0 23573 5 1 1 23572
0 23574 7 1 2 66018 77635
0 23575 5 4 1 23574
0 23576 7 1 2 59323 93010
0 23577 5 1 1 23576
0 23578 7 1 2 89240 23577
0 23579 7 1 2 23573 23578
0 23580 5 1 1 23579
0 23581 7 1 2 67627 23580
0 23582 5 1 1 23581
0 23583 7 1 2 76896 73994
0 23584 5 1 1 23583
0 23585 7 1 2 71720 93011
0 23586 5 1 1 23585
0 23587 7 2 2 70278 71618
0 23588 5 3 1 93014
0 23589 7 1 2 23586 93016
0 23590 7 1 2 23584 23589
0 23591 7 1 2 23582 23590
0 23592 5 1 1 23591
0 23593 7 1 2 61332 23592
0 23594 5 1 1 23593
0 23595 7 1 2 23567 23594
0 23596 5 1 1 23595
0 23597 7 1 2 91927 23596
0 23598 5 1 1 23597
0 23599 7 1 2 71721 76145
0 23600 5 1 1 23599
0 23601 7 1 2 73848 23600
0 23602 5 2 1 23601
0 23603 7 1 2 90600 93019
0 23604 5 1 1 23603
0 23605 7 2 2 72107 77778
0 23606 7 3 2 61333 82609
0 23607 7 1 2 93021 93023
0 23608 5 1 1 23607
0 23609 7 1 2 23604 23608
0 23610 5 1 1 23609
0 23611 7 1 2 59324 23610
0 23612 5 1 1 23611
0 23613 7 4 2 61524 74817
0 23614 7 1 2 93022 93026
0 23615 5 1 1 23614
0 23616 7 1 2 23612 23615
0 23617 5 1 1 23616
0 23618 7 1 2 78416 23617
0 23619 5 1 1 23618
0 23620 7 1 2 69725 76146
0 23621 5 1 1 23620
0 23622 7 1 2 73849 23621
0 23623 5 1 1 23622
0 23624 7 1 2 72108 23623
0 23625 5 1 1 23624
0 23626 7 1 2 69404 93020
0 23627 5 1 1 23626
0 23628 7 1 2 23625 23627
0 23629 5 1 1 23628
0 23630 7 1 2 67315 23629
0 23631 5 1 1 23630
0 23632 7 1 2 71780 71920
0 23633 7 1 2 79973 23632
0 23634 5 1 1 23633
0 23635 7 1 2 73845 23634
0 23636 5 1 1 23635
0 23637 7 1 2 23631 23636
0 23638 5 1 1 23637
0 23639 7 1 2 90601 23638
0 23640 5 1 1 23639
0 23641 7 1 2 23619 23640
0 23642 7 1 2 23598 23641
0 23643 5 1 1 23642
0 23644 7 1 2 59886 23643
0 23645 5 1 1 23644
0 23646 7 2 2 61062 88453
0 23647 5 1 1 93030
0 23648 7 1 2 90291 23647
0 23649 5 1 1 23648
0 23650 7 1 2 67316 23649
0 23651 5 1 1 23650
0 23652 7 1 2 61063 90262
0 23653 5 1 1 23652
0 23654 7 1 2 23651 23653
0 23655 5 1 1 23654
0 23656 7 1 2 91928 23655
0 23657 5 1 1 23656
0 23658 7 1 2 81426 71921
0 23659 5 1 1 23658
0 23660 7 2 2 63437 73818
0 23661 7 1 2 60525 93032
0 23662 7 1 2 23659 23661
0 23663 5 1 1 23662
0 23664 7 1 2 23657 23663
0 23665 5 1 1 23664
0 23666 7 1 2 60921 23665
0 23667 5 1 1 23666
0 23668 7 1 2 82299 90602
0 23669 5 1 1 23668
0 23670 7 1 2 62980 82610
0 23671 7 1 2 83177 23670
0 23672 5 1 1 23671
0 23673 7 1 2 23669 23672
0 23674 5 1 1 23673
0 23675 7 1 2 61064 23674
0 23676 5 1 1 23675
0 23677 7 1 2 23667 23676
0 23678 5 1 1 23677
0 23679 7 1 2 59540 23678
0 23680 5 1 1 23679
0 23681 7 1 2 74795 90603
0 23682 5 1 1 23681
0 23683 7 2 2 69559 75111
0 23684 7 1 2 83901 93034
0 23685 5 1 1 23684
0 23686 7 1 2 23682 23685
0 23687 5 1 1 23686
0 23688 7 1 2 69116 23687
0 23689 5 1 1 23688
0 23690 7 1 2 69405 91929
0 23691 5 1 1 23690
0 23692 7 1 2 90616 23691
0 23693 5 1 1 23692
0 23694 7 1 2 69183 23693
0 23695 5 1 1 23694
0 23696 7 6 2 60526 60799
0 23697 7 1 2 75438 93036
0 23698 5 1 1 23697
0 23699 7 2 2 69184 85906
0 23700 5 1 1 93042
0 23701 7 1 2 62981 93043
0 23702 5 1 1 23701
0 23703 7 1 2 23698 23702
0 23704 5 1 1 23703
0 23705 7 1 2 59325 23704
0 23706 5 1 1 23705
0 23707 7 1 2 23695 23706
0 23708 7 1 2 23689 23707
0 23709 5 1 1 23708
0 23710 7 1 2 67628 23709
0 23711 5 1 1 23710
0 23712 7 2 2 59326 93037
0 23713 7 1 2 76345 80116
0 23714 7 1 2 93044 23713
0 23715 5 2 1 23714
0 23716 7 1 2 23711 93046
0 23717 5 1 1 23716
0 23718 7 1 2 61065 23717
0 23719 5 1 1 23718
0 23720 7 1 2 83271 75999
0 23721 7 1 2 93045 23720
0 23722 5 1 1 23721
0 23723 7 1 2 23719 23722
0 23724 7 1 2 23680 23723
0 23725 5 1 1 23724
0 23726 7 1 2 61334 23725
0 23727 5 1 1 23726
0 23728 7 1 2 23645 23727
0 23729 5 1 1 23728
0 23730 7 1 2 60144 23729
0 23731 5 1 1 23730
0 23732 7 1 2 70391 90604
0 23733 5 1 1 23732
0 23734 7 1 2 85907 89721
0 23735 7 1 2 74632 23734
0 23736 5 1 1 23735
0 23737 7 1 2 23733 23736
0 23738 5 1 1 23737
0 23739 7 1 2 59541 23738
0 23740 5 1 1 23739
0 23741 7 1 2 93047 23740
0 23742 5 1 1 23741
0 23743 7 1 2 59887 73924
0 23744 7 1 2 23742 23743
0 23745 5 1 1 23744
0 23746 7 1 2 23731 23745
0 23747 5 1 1 23746
0 23748 7 1 2 92967 23747
0 23749 5 1 1 23748
0 23750 7 1 2 23563 23749
0 23751 7 1 2 23176 23750
0 23752 5 1 1 23751
0 23753 7 1 2 66688 23752
0 23754 5 1 1 23753
0 23755 7 1 2 66260 82159
0 23756 5 2 1 23755
0 23757 7 1 2 71215 93048
0 23758 5 1 1 23757
0 23759 7 1 2 71981 78406
0 23760 5 2 1 23759
0 23761 7 1 2 59327 93050
0 23762 5 2 1 23761
0 23763 7 1 2 69406 75969
0 23764 5 1 1 23763
0 23765 7 1 2 74500 23764
0 23766 7 2 2 93052 23765
0 23767 5 3 1 93054
0 23768 7 1 2 73505 93056
0 23769 5 1 1 23768
0 23770 7 1 2 77722 23769
0 23771 7 1 2 23758 23770
0 23772 5 1 1 23771
0 23773 7 1 2 62982 23772
0 23774 5 1 1 23773
0 23775 7 1 2 5887 23774
0 23776 5 1 1 23775
0 23777 7 1 2 66485 23776
0 23778 5 1 1 23777
0 23779 7 1 2 66019 81511
0 23780 5 1 1 23779
0 23781 7 1 2 66486 23780
0 23782 5 1 1 23781
0 23783 7 1 2 86274 23782
0 23784 5 1 1 23783
0 23785 7 1 2 67983 23784
0 23786 5 1 1 23785
0 23787 7 1 2 76208 76708
0 23788 5 2 1 23787
0 23789 7 1 2 62983 93059
0 23790 5 1 1 23789
0 23791 7 1 2 66020 73098
0 23792 5 1 1 23791
0 23793 7 1 2 60145 23792
0 23794 5 1 1 23793
0 23795 7 1 2 83830 23794
0 23796 5 1 1 23795
0 23797 7 1 2 23790 23796
0 23798 5 1 1 23797
0 23799 7 1 2 61525 23798
0 23800 5 1 1 23799
0 23801 7 1 2 23786 23800
0 23802 5 1 1 23801
0 23803 7 1 2 66261 23802
0 23804 5 1 1 23803
0 23805 7 1 2 75984 76944
0 23806 5 2 1 23805
0 23807 7 1 2 81922 93061
0 23808 5 1 1 23807
0 23809 7 1 2 82409 23808
0 23810 5 1 1 23809
0 23811 7 1 2 64961 78931
0 23812 5 2 1 23811
0 23813 7 1 2 3091 93063
0 23814 5 1 1 23813
0 23815 7 1 2 61526 23814
0 23816 5 1 1 23815
0 23817 7 1 2 23810 23816
0 23818 5 1 1 23817
0 23819 7 1 2 62641 23818
0 23820 5 1 1 23819
0 23821 7 1 2 71216 93057
0 23822 5 1 1 23821
0 23823 7 1 2 73494 23822
0 23824 7 1 2 82160 23823
0 23825 5 1 1 23824
0 23826 7 1 2 66487 23825
0 23827 5 1 1 23826
0 23828 7 1 2 62984 23827
0 23829 5 1 1 23828
0 23830 7 1 2 67629 18262
0 23831 7 1 2 23829 23830
0 23832 5 1 1 23831
0 23833 7 1 2 23820 23832
0 23834 7 1 2 23804 23833
0 23835 7 1 2 23778 23834
0 23836 5 1 1 23835
0 23837 7 1 2 60527 23836
0 23838 5 1 1 23837
0 23839 7 1 2 78190 82163
0 23840 5 1 1 23839
0 23841 7 1 2 80614 78887
0 23842 5 1 1 23841
0 23843 7 1 2 23840 23842
0 23844 5 1 1 23843
0 23845 7 1 2 70912 23844
0 23846 5 1 1 23845
0 23847 7 1 2 62642 93055
0 23848 5 1 1 23847
0 23849 7 1 2 72226 23848
0 23850 5 1 1 23849
0 23851 7 2 2 62643 73292
0 23852 5 1 1 93065
0 23853 7 2 2 59328 23852
0 23854 5 1 1 93067
0 23855 7 1 2 67630 88518
0 23856 5 2 1 23855
0 23857 7 2 2 23854 93069
0 23858 5 1 1 93071
0 23859 7 1 2 69117 23858
0 23860 5 1 1 23859
0 23861 7 1 2 69308 73256
0 23862 5 1 1 23861
0 23863 7 1 2 76326 23862
0 23864 7 1 2 23860 23863
0 23865 5 1 1 23864
0 23866 7 1 2 71217 23865
0 23867 5 1 1 23866
0 23868 7 1 2 23850 23867
0 23869 5 1 1 23868
0 23870 7 1 2 83011 23869
0 23871 5 1 1 23870
0 23872 7 1 2 23846 23871
0 23873 5 1 1 23872
0 23874 7 1 2 75879 23873
0 23875 5 1 1 23874
0 23876 7 1 2 23838 23875
0 23877 5 1 1 23876
0 23878 7 1 2 63438 23877
0 23879 5 1 1 23878
0 23880 7 1 2 77873 87559
0 23881 5 1 1 23880
0 23882 7 1 2 69804 23881
0 23883 5 1 1 23882
0 23884 7 3 2 62985 78532
0 23885 5 1 1 93073
0 23886 7 1 2 23883 23885
0 23887 5 1 1 23886
0 23888 7 1 2 65853 23887
0 23889 5 1 1 23888
0 23890 7 3 2 80751 77294
0 23891 5 1 1 93076
0 23892 7 1 2 23889 23891
0 23893 5 1 1 23892
0 23894 7 1 2 64721 23893
0 23895 5 1 1 23894
0 23896 7 1 2 93064 23895
0 23897 5 1 1 23896
0 23898 7 1 2 75569 23897
0 23899 5 1 1 23898
0 23900 7 3 2 62986 73869
0 23901 5 1 1 93079
0 23902 7 1 2 66021 93080
0 23903 5 1 1 23902
0 23904 7 1 2 1969 23903
0 23905 5 1 1 23904
0 23906 7 1 2 86685 23905
0 23907 5 1 1 23906
0 23908 7 1 2 23899 23907
0 23909 5 1 1 23908
0 23910 7 1 2 62644 23909
0 23911 5 1 1 23910
0 23912 7 2 2 64501 75417
0 23913 5 3 1 93082
0 23914 7 1 2 73870 88038
0 23915 5 1 1 23914
0 23916 7 1 2 90883 23915
0 23917 5 2 1 23916
0 23918 7 1 2 62987 93087
0 23919 5 1 1 23918
0 23920 7 1 2 93084 23919
0 23921 5 1 1 23920
0 23922 7 1 2 65854 23921
0 23923 5 1 1 23922
0 23924 7 1 2 62988 78877
0 23925 5 1 1 23924
0 23926 7 1 2 85053 90347
0 23927 7 1 2 23925 23926
0 23928 5 1 1 23927
0 23929 7 1 2 64722 23928
0 23930 5 1 1 23929
0 23931 7 1 2 90388 23930
0 23932 7 1 2 23923 23931
0 23933 5 1 1 23932
0 23934 7 1 2 78622 90383
0 23935 5 1 1 23934
0 23936 7 1 2 61066 23935
0 23937 5 1 1 23936
0 23938 7 1 2 64962 23937
0 23939 7 1 2 23933 23938
0 23940 5 1 1 23939
0 23941 7 1 2 75204 6727
0 23942 5 1 1 23941
0 23943 7 1 2 72445 75038
0 23944 5 1 1 23943
0 23945 7 1 2 73884 23944
0 23946 5 1 1 23945
0 23947 7 1 2 65855 23946
0 23948 5 1 1 23947
0 23949 7 1 2 78879 23948
0 23950 5 1 1 23949
0 23951 7 1 2 86831 23950
0 23952 5 1 1 23951
0 23953 7 1 2 23942 23952
0 23954 7 1 2 23940 23953
0 23955 5 1 1 23954
0 23956 7 1 2 66262 23955
0 23957 5 1 1 23956
0 23958 7 2 2 64502 79533
0 23959 5 2 1 93089
0 23960 7 3 2 64503 84647
0 23961 5 1 1 93093
0 23962 7 1 2 17643 23961
0 23963 5 1 1 23962
0 23964 7 1 2 69805 23963
0 23965 5 1 1 23964
0 23966 7 1 2 93091 23965
0 23967 5 1 1 23966
0 23968 7 1 2 62305 23967
0 23969 5 1 1 23968
0 23970 7 1 2 1867 23969
0 23971 5 1 1 23970
0 23972 7 1 2 66488 23971
0 23973 5 1 1 23972
0 23974 7 1 2 23957 23973
0 23975 7 1 2 23911 23974
0 23976 5 1 1 23975
0 23977 7 1 2 90140 23976
0 23978 5 1 1 23977
0 23979 7 1 2 23879 23978
0 23980 5 1 1 23979
0 23981 7 1 2 63967 23980
0 23982 5 1 1 23981
0 23983 7 1 2 72446 73166
0 23984 7 1 2 80308 88268
0 23985 7 1 2 89242 23984
0 23986 7 1 2 23983 23985
0 23987 5 1 1 23986
0 23988 7 1 2 23982 23987
0 23989 5 1 1 23988
0 23990 7 1 2 68671 23989
0 23991 5 1 1 23990
0 23992 7 1 2 77426 93001
0 23993 5 1 1 23992
0 23994 7 1 2 80490 84320
0 23995 5 1 1 23994
0 23996 7 2 2 69910 72227
0 23997 7 1 2 78854 93096
0 23998 5 1 1 23997
0 23999 7 1 2 90499 88931
0 24000 5 1 1 23999
0 24001 7 1 2 69560 90983
0 24002 7 1 2 24000 24001
0 24003 5 1 1 24002
0 24004 7 1 2 23998 24003
0 24005 5 2 1 24004
0 24006 7 1 2 72191 93098
0 24007 5 1 1 24006
0 24008 7 1 2 23995 24007
0 24009 7 1 2 23993 24008
0 24010 5 1 1 24009
0 24011 7 1 2 74651 24010
0 24012 5 1 1 24011
0 24013 7 1 2 83902 7498
0 24014 5 1 1 24013
0 24015 7 3 2 67984 74734
0 24016 7 2 2 79849 72192
0 24017 7 1 2 69561 93103
0 24018 5 1 1 24017
0 24019 7 1 2 78360 24018
0 24020 5 1 1 24019
0 24021 7 1 2 93100 24020
0 24022 5 1 1 24021
0 24023 7 1 2 24014 24022
0 24024 5 1 1 24023
0 24025 7 1 2 61067 24024
0 24026 5 1 1 24025
0 24027 7 2 2 70279 82893
0 24028 5 2 1 93105
0 24029 7 1 2 62989 90025
0 24030 7 1 2 93107 24029
0 24031 7 1 2 14687 24030
0 24032 5 1 1 24031
0 24033 7 1 2 61527 92173
0 24034 7 1 2 24032 24033
0 24035 5 1 1 24034
0 24036 7 1 2 24026 24035
0 24037 5 1 1 24036
0 24038 7 1 2 59888 24037
0 24039 5 1 1 24038
0 24040 7 3 2 59889 73319
0 24041 7 1 2 74735 89393
0 24042 7 1 2 93109 24041
0 24043 5 1 1 24042
0 24044 7 1 2 69118 83903
0 24045 7 1 2 92934 24044
0 24046 5 1 1 24045
0 24047 7 1 2 24043 24046
0 24048 5 1 1 24047
0 24049 7 1 2 72571 24048
0 24050 5 1 1 24049
0 24051 7 2 2 73688 77427
0 24052 5 2 1 93112
0 24053 7 1 2 60922 91600
0 24054 5 1 1 24053
0 24055 7 1 2 59890 71599
0 24056 5 1 1 24055
0 24057 7 1 2 91583 24056
0 24058 7 1 2 24054 24057
0 24059 5 1 1 24058
0 24060 7 1 2 62990 24059
0 24061 5 1 1 24060
0 24062 7 1 2 93114 24061
0 24063 5 1 1 24062
0 24064 7 1 2 69911 24063
0 24065 5 1 1 24064
0 24066 7 2 2 67631 91555
0 24067 7 1 2 73716 93116
0 24068 5 1 1 24067
0 24069 7 1 2 81444 73320
0 24070 5 1 1 24069
0 24071 7 1 2 24068 24070
0 24072 5 1 1 24071
0 24073 7 1 2 62991 24072
0 24074 5 1 1 24073
0 24075 7 1 2 81935 84725
0 24076 5 1 1 24075
0 24077 7 1 2 77428 24076
0 24078 5 1 1 24077
0 24079 7 1 2 71371 82664
0 24080 5 1 1 24079
0 24081 7 1 2 69562 24080
0 24082 5 2 1 24081
0 24083 7 1 2 88942 93118
0 24084 5 1 1 24083
0 24085 7 1 2 72109 92174
0 24086 7 1 2 24084 24085
0 24087 5 1 1 24086
0 24088 7 1 2 24078 24087
0 24089 7 1 2 24074 24088
0 24090 7 1 2 24065 24089
0 24091 5 1 1 24090
0 24092 7 1 2 61528 24091
0 24093 5 1 1 24092
0 24094 7 1 2 24050 24093
0 24095 7 1 2 24039 24094
0 24096 5 1 1 24095
0 24097 7 1 2 70608 24096
0 24098 5 1 1 24097
0 24099 7 1 2 24012 24098
0 24100 5 1 1 24099
0 24101 7 1 2 60347 24100
0 24102 5 1 1 24101
0 24103 7 1 2 70167 88796
0 24104 5 1 1 24103
0 24105 7 1 2 88800 24104
0 24106 5 1 1 24105
0 24107 7 1 2 76258 24106
0 24108 5 1 1 24107
0 24109 7 1 2 76444 73506
0 24110 5 1 1 24109
0 24111 7 1 2 70255 24110
0 24112 5 1 1 24111
0 24113 7 1 2 76407 24112
0 24114 5 1 1 24113
0 24115 7 3 2 71308 69984
0 24116 5 1 1 93120
0 24117 7 1 2 74692 24116
0 24118 5 1 1 24117
0 24119 7 1 2 70917 24118
0 24120 7 1 2 24114 24119
0 24121 7 1 2 24108 24120
0 24122 5 2 1 24121
0 24123 7 1 2 66489 93123
0 24124 5 1 1 24123
0 24125 7 1 2 76729 87286
0 24126 5 2 1 24125
0 24127 7 1 2 61529 93125
0 24128 5 1 1 24127
0 24129 7 1 2 67985 74374
0 24130 7 1 2 24128 24129
0 24131 7 1 2 24124 24130
0 24132 5 1 1 24131
0 24133 7 1 2 59542 85792
0 24134 5 1 1 24133
0 24135 7 1 2 88531 24134
0 24136 5 1 1 24135
0 24137 7 1 2 90769 24136
0 24138 5 1 1 24137
0 24139 7 1 2 72169 90787
0 24140 5 1 1 24139
0 24141 7 1 2 71332 24140
0 24142 5 1 1 24141
0 24143 7 1 2 24138 24142
0 24144 5 1 1 24143
0 24145 7 2 2 66490 88591
0 24146 5 2 1 93127
0 24147 7 1 2 24144 93129
0 24148 5 1 1 24147
0 24149 7 1 2 74046 88586
0 24150 5 1 1 24149
0 24151 7 1 2 62992 89501
0 24152 7 1 2 24150 24151
0 24153 7 1 2 24148 24152
0 24154 5 1 1 24153
0 24155 7 1 2 67632 24154
0 24156 7 1 2 24132 24155
0 24157 5 1 1 24156
0 24158 7 1 2 62993 88673
0 24159 5 1 1 24158
0 24160 7 1 2 71218 92175
0 24161 7 1 2 24159 24160
0 24162 5 1 1 24161
0 24163 7 1 2 76561 78432
0 24164 5 1 1 24163
0 24165 7 1 2 74832 92975
0 24166 5 1 1 24165
0 24167 7 1 2 77429 24166
0 24168 5 1 1 24167
0 24169 7 1 2 24164 24168
0 24170 7 1 2 24162 24169
0 24171 5 1 1 24170
0 24172 7 1 2 90770 24171
0 24173 5 1 1 24172
0 24174 7 1 2 73225 91287
0 24175 5 1 1 24174
0 24176 7 2 2 62994 24175
0 24177 5 1 1 93131
0 24178 7 1 2 83043 24177
0 24179 5 1 1 24178
0 24180 7 1 2 75307 24179
0 24181 5 1 1 24180
0 24182 7 1 2 76521 89269
0 24183 5 1 1 24182
0 24184 7 1 2 19696 24183
0 24185 5 1 1 24184
0 24186 7 1 2 72110 24185
0 24187 5 1 1 24186
0 24188 7 1 2 71289 76640
0 24189 5 2 1 24188
0 24190 7 1 2 83309 93133
0 24191 5 1 1 24190
0 24192 7 1 2 75777 24191
0 24193 5 1 1 24192
0 24194 7 1 2 24187 24193
0 24195 5 1 1 24194
0 24196 7 1 2 67986 24195
0 24197 5 1 1 24196
0 24198 7 1 2 24181 24197
0 24199 5 1 1 24198
0 24200 7 1 2 70168 24199
0 24201 5 1 1 24200
0 24202 7 1 2 60800 90013
0 24203 5 1 1 24202
0 24204 7 1 2 77387 24203
0 24205 5 2 1 24204
0 24206 7 1 2 60146 93135
0 24207 5 1 1 24206
0 24208 7 1 2 80635 90014
0 24209 5 1 1 24208
0 24210 7 1 2 90041 24209
0 24211 7 1 2 24207 24210
0 24212 5 2 1 24211
0 24213 7 1 2 59329 93137
0 24214 5 1 1 24213
0 24215 7 1 2 77242 92739
0 24216 5 1 1 24215
0 24217 7 1 2 24214 24216
0 24218 5 1 1 24217
0 24219 7 1 2 90362 24218
0 24220 5 1 1 24219
0 24221 7 1 2 77057 88929
0 24222 5 1 1 24221
0 24223 7 1 2 90042 24222
0 24224 5 1 1 24223
0 24225 7 1 2 70169 24224
0 24226 5 1 1 24225
0 24227 7 1 2 92740 92973
0 24228 5 1 1 24227
0 24229 7 1 2 24226 24228
0 24230 5 1 1 24229
0 24231 7 1 2 69119 24230
0 24232 5 1 1 24231
0 24233 7 1 2 62645 76510
0 24234 5 1 1 24233
0 24235 7 1 2 61335 24234
0 24236 5 2 1 24235
0 24237 7 1 2 78373 93139
0 24238 5 1 1 24237
0 24239 7 1 2 76688 24238
0 24240 5 1 1 24239
0 24241 7 1 2 61530 24240
0 24242 5 1 1 24241
0 24243 7 1 2 82836 19915
0 24244 5 1 1 24243
0 24245 7 1 2 70609 24244
0 24246 5 1 1 24245
0 24247 7 1 2 83918 92143
0 24248 7 1 2 24246 24247
0 24249 5 1 1 24248
0 24250 7 1 2 76774 24249
0 24251 5 1 1 24250
0 24252 7 1 2 24242 24251
0 24253 7 1 2 24232 24252
0 24254 7 1 2 24220 24253
0 24255 7 1 2 24201 24254
0 24256 7 1 2 24173 24255
0 24257 7 1 2 24157 24256
0 24258 5 1 1 24257
0 24259 7 1 2 60528 24258
0 24260 5 1 1 24259
0 24261 7 1 2 24102 24260
0 24262 5 1 1 24261
0 24263 7 1 2 81018 24262
0 24264 5 1 1 24263
0 24265 7 1 2 83014 93009
0 24266 5 1 1 24265
0 24267 7 1 2 59543 24266
0 24268 5 1 1 24267
0 24269 7 1 2 74018 76985
0 24270 5 1 1 24269
0 24271 7 1 2 73234 24270
0 24272 5 1 1 24271
0 24273 7 2 2 69120 83016
0 24274 5 1 1 93141
0 24275 7 1 2 66263 24274
0 24276 7 1 2 24272 24275
0 24277 7 1 2 24268 24276
0 24278 5 1 1 24277
0 24279 7 1 2 60147 24278
0 24280 5 1 1 24279
0 24281 7 1 2 69185 73285
0 24282 5 2 1 24281
0 24283 7 2 2 66264 93143
0 24284 5 1 1 93145
0 24285 7 1 2 59891 24284
0 24286 5 1 1 24285
0 24287 7 1 2 64504 70357
0 24288 5 2 1 24287
0 24289 7 1 2 61336 70420
0 24290 7 1 2 93147 24289
0 24291 5 1 1 24290
0 24292 7 1 2 24286 24291
0 24293 5 1 1 24292
0 24294 7 1 2 59330 24293
0 24295 5 1 1 24294
0 24296 7 1 2 81568 88515
0 24297 5 2 1 24296
0 24298 7 1 2 76998 93149
0 24299 5 1 1 24298
0 24300 7 1 2 69407 74488
0 24301 5 1 1 24300
0 24302 7 1 2 24299 24301
0 24303 5 1 1 24302
0 24304 7 1 2 61337 24303
0 24305 5 1 1 24304
0 24306 7 1 2 75570 24305
0 24307 7 1 2 24295 24306
0 24308 7 1 2 24280 24307
0 24309 5 1 1 24308
0 24310 7 1 2 67987 24309
0 24311 5 1 1 24310
0 24312 7 1 2 83478 82060
0 24313 5 1 1 24312
0 24314 7 1 2 81369 71489
0 24315 5 2 1 24314
0 24316 7 1 2 24313 93151
0 24317 7 1 2 24311 24316
0 24318 5 1 1 24317
0 24319 7 1 2 75308 24318
0 24320 5 1 1 24319
0 24321 7 3 2 61531 71490
0 24322 7 1 2 81373 93153
0 24323 5 1 1 24322
0 24324 7 1 2 24320 24323
0 24325 5 1 1 24324
0 24326 7 1 2 73819 24325
0 24327 5 1 1 24326
0 24328 7 1 2 69912 91955
0 24329 5 1 1 24328
0 24330 7 1 2 65196 24329
0 24331 5 1 1 24330
0 24332 7 1 2 59892 24331
0 24333 5 1 1 24332
0 24334 7 3 2 72572 73415
0 24335 5 1 1 93156
0 24336 7 1 2 65197 24335
0 24337 5 1 1 24336
0 24338 7 1 2 69121 24337
0 24339 5 1 1 24338
0 24340 7 3 2 71419 80931
0 24341 5 1 1 93159
0 24342 7 1 2 65198 24341
0 24343 5 2 1 24342
0 24344 7 1 2 59544 93162
0 24345 5 1 1 24344
0 24346 7 1 2 74266 24345
0 24347 7 1 2 24339 24346
0 24348 7 1 2 24333 24347
0 24349 5 1 1 24348
0 24350 7 1 2 67988 24349
0 24351 5 1 1 24350
0 24352 7 1 2 71400 24351
0 24353 5 1 1 24352
0 24354 7 1 2 84956 24353
0 24355 5 1 1 24354
0 24356 7 1 2 73914 74945
0 24357 5 3 1 24356
0 24358 7 1 2 71395 92578
0 24359 5 1 1 24358
0 24360 7 1 2 93164 24359
0 24361 5 1 1 24360
0 24362 7 1 2 59893 24361
0 24363 5 1 1 24362
0 24364 7 1 2 71667 83430
0 24365 5 1 1 24364
0 24366 7 1 2 93165 24365
0 24367 5 1 1 24366
0 24368 7 1 2 59545 24367
0 24369 5 1 1 24368
0 24370 7 2 2 92718 92993
0 24371 5 1 1 93167
0 24372 7 1 2 93166 24371
0 24373 5 1 1 24372
0 24374 7 1 2 69122 24373
0 24375 5 1 1 24374
0 24376 7 1 2 20873 24375
0 24377 7 1 2 24369 24376
0 24378 7 1 2 24363 24377
0 24379 5 1 1 24378
0 24380 7 1 2 67989 24379
0 24381 5 1 1 24380
0 24382 7 1 2 69123 83973
0 24383 5 1 1 24382
0 24384 7 2 2 60148 73355
0 24385 5 1 1 93169
0 24386 7 1 2 64723 24385
0 24387 5 1 1 24386
0 24388 7 1 2 92580 88662
0 24389 5 1 1 24388
0 24390 7 1 2 24387 24389
0 24391 5 1 1 24390
0 24392 7 1 2 24383 24391
0 24393 5 1 1 24392
0 24394 7 1 2 92159 24393
0 24395 5 1 1 24394
0 24396 7 1 2 75571 24395
0 24397 5 1 1 24396
0 24398 7 1 2 76147 24397
0 24399 5 1 1 24398
0 24400 7 1 2 72952 93024
0 24401 5 1 1 24400
0 24402 7 1 2 67068 81889
0 24403 5 1 1 24402
0 24404 7 1 2 62995 24403
0 24405 5 1 1 24404
0 24406 7 2 2 70170 91246
0 24407 5 2 1 93171
0 24408 7 1 2 75572 93173
0 24409 5 1 1 24408
0 24410 7 1 2 92689 24409
0 24411 7 1 2 24405 24410
0 24412 5 1 1 24411
0 24413 7 1 2 24401 24412
0 24414 7 1 2 24399 24413
0 24415 7 1 2 24381 24414
0 24416 7 1 2 24355 24415
0 24417 7 1 2 24327 24416
0 24418 5 1 1 24417
0 24419 7 1 2 60529 24418
0 24420 5 1 1 24419
0 24421 7 1 2 82963 71873
0 24422 5 1 1 24421
0 24423 7 1 2 89576 24422
0 24424 5 1 1 24423
0 24425 7 1 2 91847 24424
0 24426 5 1 1 24425
0 24427 7 1 2 78145 76136
0 24428 5 1 1 24427
0 24429 7 1 2 75309 24428
0 24430 5 1 1 24429
0 24431 7 1 2 78130 73925
0 24432 5 1 1 24431
0 24433 7 1 2 24430 24432
0 24434 5 1 1 24433
0 24435 7 1 2 60530 24434
0 24436 5 1 1 24435
0 24437 7 7 2 67990 71874
0 24438 7 1 2 90011 93175
0 24439 5 1 1 24438
0 24440 7 1 2 24436 24439
0 24441 5 1 1 24440
0 24442 7 1 2 60149 24441
0 24443 5 1 1 24442
0 24444 7 1 2 24426 24443
0 24445 5 1 1 24444
0 24446 7 1 2 81896 24445
0 24447 5 1 1 24446
0 24448 7 2 2 84974 90369
0 24449 5 1 1 93182
0 24450 7 2 2 61532 82928
0 24451 7 1 2 89107 93184
0 24452 7 1 2 93183 24451
0 24453 5 1 1 24452
0 24454 7 4 2 67991 91671
0 24455 5 1 1 93186
0 24456 7 1 2 92477 88963
0 24457 7 1 2 74545 24456
0 24458 7 1 2 93187 24457
0 24459 5 1 1 24458
0 24460 7 1 2 63968 24459
0 24461 7 1 2 24453 24460
0 24462 7 1 2 24447 24461
0 24463 7 1 2 24420 24462
0 24464 5 1 1 24463
0 24465 7 2 2 65856 76959
0 24466 5 1 1 93190
0 24467 7 1 2 74784 93191
0 24468 5 1 1 24467
0 24469 7 1 2 76361 82906
0 24470 5 1 1 24469
0 24471 7 1 2 24468 24470
0 24472 5 3 1 24471
0 24473 7 1 2 75152 85460
0 24474 5 9 1 24473
0 24475 7 11 2 62646 77858
0 24476 5 4 1 93204
0 24477 7 1 2 93195 93205
0 24478 5 1 1 24477
0 24479 7 1 2 85483 24478
0 24480 5 2 1 24479
0 24481 7 1 2 66265 93219
0 24482 7 1 2 93192 24481
0 24483 5 1 1 24482
0 24484 7 1 2 71430 81956
0 24485 7 1 2 84044 24484
0 24486 5 1 1 24485
0 24487 7 1 2 24483 24486
0 24488 5 1 1 24487
0 24489 7 1 2 62996 24488
0 24490 5 1 1 24489
0 24491 7 1 2 61338 82737
0 24492 5 1 1 24491
0 24493 7 1 2 85273 90906
0 24494 7 1 2 24492 24493
0 24495 5 1 1 24494
0 24496 7 1 2 68871 24495
0 24497 7 1 2 24490 24496
0 24498 5 1 1 24497
0 24499 7 1 2 63439 24498
0 24500 7 1 2 24464 24499
0 24501 5 1 1 24500
0 24502 7 1 2 24264 24501
0 24503 5 1 1 24502
0 24504 7 1 2 63738 24503
0 24505 5 1 1 24504
0 24506 7 3 2 60531 73950
0 24507 5 1 1 93221
0 24508 7 2 2 73477 93222
0 24509 7 1 2 84150 93224
0 24510 5 1 1 24509
0 24511 7 1 2 85617 90617
0 24512 5 1 1 24511
0 24513 7 1 2 81740 91996
0 24514 7 1 2 24512 24513
0 24515 5 1 1 24514
0 24516 7 1 2 24510 24515
0 24517 5 1 1 24516
0 24518 7 1 2 64724 24517
0 24519 5 1 1 24518
0 24520 7 2 2 77779 77558
0 24521 7 1 2 76182 81079
0 24522 7 1 2 93226 24521
0 24523 5 1 1 24522
0 24524 7 1 2 24519 24523
0 24525 5 1 1 24524
0 24526 7 1 2 77859 24525
0 24527 5 1 1 24526
0 24528 7 4 2 68672 79136
0 24529 5 1 1 93228
0 24530 7 1 2 82351 85969
0 24531 5 1 1 24530
0 24532 7 1 2 90431 24531
0 24533 5 1 1 24532
0 24534 7 2 2 63440 89532
0 24535 5 1 1 93232
0 24536 7 1 2 24533 24535
0 24537 5 1 1 24536
0 24538 7 1 2 93229 24537
0 24539 5 1 1 24538
0 24540 7 1 2 24527 24539
0 24541 5 1 1 24540
0 24542 7 1 2 62306 24541
0 24543 5 1 1 24542
0 24544 7 1 2 81535 77559
0 24545 7 1 2 85644 24544
0 24546 5 1 1 24545
0 24547 7 1 2 24543 24546
0 24548 5 1 1 24547
0 24549 7 1 2 64505 24548
0 24550 5 1 1 24549
0 24551 7 2 2 80049 85383
0 24552 7 1 2 77189 93234
0 24553 5 1 1 24552
0 24554 7 1 2 85618 85978
0 24555 5 1 1 24554
0 24556 7 1 2 66491 24555
0 24557 5 1 1 24556
0 24558 7 1 2 24553 24557
0 24559 5 1 1 24558
0 24560 7 1 2 62647 24559
0 24561 5 1 1 24560
0 24562 7 1 2 79534 84986
0 24563 5 1 1 24562
0 24564 7 1 2 24561 24563
0 24565 5 1 1 24564
0 24566 7 1 2 93230 24565
0 24567 5 1 1 24566
0 24568 7 1 2 24550 24567
0 24569 5 1 1 24568
0 24570 7 1 2 72549 24569
0 24571 5 1 1 24570
0 24572 7 1 2 24505 24571
0 24573 7 1 2 23991 24572
0 24574 5 1 1 24573
0 24575 7 1 2 61714 24574
0 24576 5 1 1 24575
0 24577 7 1 2 59331 93136
0 24578 5 1 1 24577
0 24579 7 1 2 60801 77376
0 24580 5 1 1 24579
0 24581 7 1 2 24578 24580
0 24582 5 1 1 24581
0 24583 7 1 2 71219 24582
0 24584 5 1 1 24583
0 24585 7 1 2 78191 91306
0 24586 7 1 2 76914 24585
0 24587 5 1 1 24586
0 24588 7 1 2 24584 24587
0 24589 5 1 1 24588
0 24590 7 1 2 68341 24589
0 24591 5 1 1 24590
0 24592 7 1 2 82340 72228
0 24593 7 1 2 83141 24592
0 24594 5 1 1 24593
0 24595 7 1 2 24591 24594
0 24596 5 1 1 24595
0 24597 7 1 2 59546 24596
0 24598 5 1 1 24597
0 24599 7 1 2 73820 77780
0 24600 5 1 1 24599
0 24601 7 4 2 59332 61068
0 24602 5 1 1 93236
0 24603 7 2 2 70280 93237
0 24604 7 1 2 86651 93240
0 24605 5 1 1 24604
0 24606 7 1 2 24600 24605
0 24607 5 1 1 24606
0 24608 7 1 2 59894 24607
0 24609 5 1 1 24608
0 24610 7 3 2 68342 78192
0 24611 7 1 2 61069 93242
0 24612 5 1 1 24611
0 24613 7 1 2 24609 24612
0 24614 5 1 1 24613
0 24615 7 1 2 61339 24614
0 24616 5 1 1 24615
0 24617 7 1 2 24598 24616
0 24618 5 1 1 24617
0 24619 7 1 2 60150 24618
0 24620 5 1 1 24619
0 24621 7 2 2 59547 93099
0 24622 5 1 1 93245
0 24623 7 1 2 81595 93246
0 24624 5 1 1 24623
0 24625 7 1 2 24620 24624
0 24626 5 1 1 24625
0 24627 7 1 2 69124 24626
0 24628 5 1 1 24627
0 24629 7 1 2 81446 70003
0 24630 5 1 1 24629
0 24631 7 1 2 60923 24630
0 24632 5 1 1 24631
0 24633 7 2 2 73461 24632
0 24634 5 1 1 93247
0 24635 7 1 2 91503 93248
0 24636 5 1 1 24635
0 24637 7 1 2 61070 24636
0 24638 5 1 1 24637
0 24639 7 1 2 7406 24638
0 24640 5 1 1 24639
0 24641 7 1 2 62997 24640
0 24642 5 1 1 24641
0 24643 7 3 2 64725 78511
0 24644 5 4 1 93249
0 24645 7 1 2 84016 93250
0 24646 5 1 1 24645
0 24647 7 1 2 83036 24646
0 24648 5 1 1 24647
0 24649 7 1 2 24642 24648
0 24650 5 1 1 24649
0 24651 7 1 2 70610 24650
0 24652 5 1 1 24651
0 24653 7 1 2 83782 82760
0 24654 5 1 1 24653
0 24655 7 1 2 91486 24654
0 24656 5 1 1 24655
0 24657 7 1 2 70796 71634
0 24658 5 1 1 24657
0 24659 7 1 2 24656 24658
0 24660 5 1 1 24659
0 24661 7 1 2 83037 92999
0 24662 5 1 1 24661
0 24663 7 1 2 24660 24662
0 24664 5 1 1 24663
0 24665 7 1 2 70171 24664
0 24666 5 1 1 24665
0 24667 7 1 2 24652 24666
0 24668 5 1 1 24667
0 24669 7 1 2 68343 24668
0 24670 5 1 1 24669
0 24671 7 4 2 60151 77377
0 24672 7 1 2 69913 82480
0 24673 5 1 1 24672
0 24674 7 3 2 81823 24673
0 24675 5 1 1 93260
0 24676 7 1 2 83212 93261
0 24677 5 1 1 24676
0 24678 7 1 2 93256 24677
0 24679 5 1 1 24678
0 24680 7 1 2 74383 77430
0 24681 7 1 2 88980 24680
0 24682 5 1 1 24681
0 24683 7 1 2 24679 24682
0 24684 5 1 1 24683
0 24685 7 1 2 68344 24684
0 24686 5 1 1 24685
0 24687 7 2 2 77033 73416
0 24688 7 1 2 83126 93263
0 24689 5 1 1 24688
0 24690 7 1 2 24686 24689
0 24691 5 1 1 24690
0 24692 7 1 2 71600 24691
0 24693 5 1 1 24692
0 24694 7 1 2 82264 88519
0 24695 5 1 1 24694
0 24696 7 1 2 74895 73299
0 24697 7 1 2 93068 24696
0 24698 5 1 1 24697
0 24699 7 1 2 24695 24698
0 24700 5 1 1 24699
0 24701 7 7 2 69186 84800
0 24702 5 3 1 93265
0 24703 7 1 2 75001 93266
0 24704 7 1 2 24700 24703
0 24705 5 1 1 24704
0 24706 7 1 2 24693 24705
0 24707 7 1 2 24670 24706
0 24708 7 1 2 24628 24707
0 24709 5 1 1 24708
0 24710 7 1 2 87854 90171
0 24711 7 1 2 24709 24710
0 24712 5 1 1 24711
0 24713 7 1 2 66828 24712
0 24714 7 1 2 24576 24713
0 24715 7 1 2 23754 24714
0 24716 5 1 1 24715
0 24717 7 2 2 70172 76730
0 24718 5 2 1 93275
0 24719 7 1 2 59333 92903
0 24720 5 1 1 24719
0 24721 7 1 2 93277 24720
0 24722 5 1 1 24721
0 24723 7 1 2 60348 24722
0 24724 5 1 1 24723
0 24725 7 1 2 72865 89254
0 24726 7 1 2 91617 24725
0 24727 5 1 1 24726
0 24728 7 1 2 24724 24727
0 24729 5 1 1 24728
0 24730 7 1 2 59895 24729
0 24731 5 1 1 24730
0 24732 7 3 2 88652 13202
0 24733 5 1 1 93279
0 24734 7 1 2 71521 24733
0 24735 5 1 1 24734
0 24736 7 1 2 24731 24735
0 24737 5 1 1 24736
0 24738 7 1 2 59548 24737
0 24739 5 1 1 24738
0 24740 7 1 2 72854 70261
0 24741 5 1 1 24740
0 24742 7 1 2 70918 24741
0 24743 5 1 1 24742
0 24744 7 1 2 60349 24743
0 24745 5 1 1 24744
0 24746 7 1 2 66689 24745
0 24747 7 1 2 24739 24746
0 24748 5 1 1 24747
0 24749 7 1 2 77190 72795
0 24750 5 1 1 24749
0 24751 7 1 2 77152 24750
0 24752 5 1 1 24751
0 24753 7 1 2 66266 24752
0 24754 5 1 1 24753
0 24755 7 1 2 61715 85283
0 24756 7 1 2 24754 24755
0 24757 5 1 1 24756
0 24758 7 1 2 67317 24757
0 24759 7 1 2 24748 24758
0 24760 5 1 1 24759
0 24761 7 2 2 83793 93251
0 24762 5 1 1 93282
0 24763 7 1 2 62098 93283
0 24764 5 1 1 24763
0 24765 7 1 2 70611 24764
0 24766 5 1 1 24765
0 24767 7 1 2 72339 74750
0 24768 5 1 1 24767
0 24769 7 1 2 67069 24768
0 24770 5 1 1 24769
0 24771 7 1 2 69914 75778
0 24772 5 1 1 24771
0 24773 7 1 2 78658 24772
0 24774 7 1 2 24770 24773
0 24775 5 1 1 24774
0 24776 7 1 2 70173 24775
0 24777 5 1 1 24776
0 24778 7 1 2 24766 24777
0 24779 5 1 1 24778
0 24780 7 1 2 85594 24779
0 24781 5 1 1 24780
0 24782 7 2 2 67070 70797
0 24783 7 1 2 79535 84251
0 24784 7 1 2 93284 24783
0 24785 5 1 1 24784
0 24786 7 1 2 24781 24785
0 24787 7 1 2 24760 24786
0 24788 5 1 1 24787
0 24789 7 1 2 62648 24788
0 24790 5 1 1 24789
0 24791 7 1 2 71660 91646
0 24792 5 1 1 24791
0 24793 7 1 2 69915 24792
0 24794 5 1 1 24793
0 24795 7 1 2 71522 88365
0 24796 5 1 1 24795
0 24797 7 1 2 24794 24796
0 24798 5 1 1 24797
0 24799 7 1 2 70486 24798
0 24800 5 2 1 24799
0 24801 7 1 2 73041 87585
0 24802 5 1 1 24801
0 24803 7 1 2 93286 24802
0 24804 5 1 1 24803
0 24805 7 1 2 92640 24804
0 24806 5 1 1 24805
0 24807 7 1 2 24790 24806
0 24808 5 1 1 24807
0 24809 7 1 2 67992 24808
0 24810 5 1 1 24809
0 24811 7 1 2 70487 82097
0 24812 5 1 1 24811
0 24813 7 1 2 60152 24812
0 24814 5 1 1 24813
0 24815 7 1 2 81745 24814
0 24816 5 1 1 24815
0 24817 7 1 2 24810 24816
0 24818 5 1 1 24817
0 24819 7 1 2 66492 24818
0 24820 5 1 1 24819
0 24821 7 1 2 73674 85645
0 24822 5 1 1 24821
0 24823 7 1 2 61340 80483
0 24824 5 3 1 24823
0 24825 7 1 2 81689 93196
0 24826 7 1 2 93288 24825
0 24827 5 1 1 24826
0 24828 7 1 2 24822 24827
0 24829 5 1 1 24828
0 24830 7 1 2 64963 24829
0 24831 5 1 1 24830
0 24832 7 1 2 79075 86880
0 24833 5 1 1 24832
0 24834 7 1 2 24831 24833
0 24835 5 1 1 24834
0 24836 7 1 2 61716 24835
0 24837 5 1 1 24836
0 24838 7 2 2 60350 80996
0 24839 7 1 2 70612 82061
0 24840 5 1 1 24839
0 24841 7 1 2 93152 24840
0 24842 5 1 1 24841
0 24843 7 1 2 73821 24842
0 24844 5 1 1 24843
0 24845 7 1 2 83455 93172
0 24846 5 1 1 24845
0 24847 7 3 2 70613 71875
0 24848 5 1 1 93293
0 24849 7 1 2 24846 24848
0 24850 7 1 2 24844 24849
0 24851 5 1 1 24850
0 24852 7 1 2 93291 24851
0 24853 5 1 1 24852
0 24854 7 1 2 24837 24853
0 24855 5 1 1 24854
0 24856 7 1 2 62998 24855
0 24857 5 1 1 24856
0 24858 7 1 2 80356 77450
0 24859 7 1 2 72796 24858
0 24860 5 1 1 24859
0 24861 7 1 2 24857 24860
0 24862 7 1 2 24820 24861
0 24863 5 1 1 24862
0 24864 7 1 2 63441 24863
0 24865 5 1 1 24864
0 24866 7 1 2 90771 92935
0 24867 5 1 1 24866
0 24868 7 3 2 67071 70244
0 24869 7 1 2 82265 93296
0 24870 5 1 1 24869
0 24871 7 1 2 24867 24870
0 24872 5 1 1 24871
0 24873 7 1 2 69916 24872
0 24874 5 1 1 24873
0 24875 7 1 2 77136 93130
0 24876 5 1 1 24875
0 24877 7 1 2 24874 24876
0 24878 5 1 1 24877
0 24879 7 1 2 67318 24878
0 24880 5 1 1 24879
0 24881 7 1 2 83885 90784
0 24882 5 1 1 24881
0 24883 7 1 2 91937 24882
0 24884 7 1 2 24880 24883
0 24885 5 1 1 24884
0 24886 7 1 2 72111 24885
0 24887 5 1 1 24886
0 24888 7 1 2 66022 76909
0 24889 5 2 1 24888
0 24890 7 1 2 67633 93299
0 24891 5 1 1 24890
0 24892 7 1 2 74796 91556
0 24893 5 1 1 24892
0 24894 7 1 2 88964 24893
0 24895 7 1 2 24891 24894
0 24896 5 1 1 24895
0 24897 7 1 2 59896 24896
0 24898 5 1 1 24897
0 24899 7 1 2 71321 71627
0 24900 5 1 1 24899
0 24901 7 1 2 93117 24900
0 24902 5 1 1 24901
0 24903 7 2 2 61071 74797
0 24904 5 2 1 93301
0 24905 7 1 2 71722 93302
0 24906 5 1 1 24905
0 24907 7 1 2 24902 24906
0 24908 7 1 2 24898 24907
0 24909 5 1 1 24908
0 24910 7 1 2 90772 24909
0 24911 5 1 1 24910
0 24912 7 2 2 74203 71876
0 24913 5 1 1 93305
0 24914 7 1 2 5702 93306
0 24915 5 1 1 24914
0 24916 7 6 2 59549 73321
0 24917 5 1 1 93307
0 24918 7 2 2 76562 81808
0 24919 5 2 1 93313
0 24920 7 1 2 93308 93314
0 24921 5 1 1 24920
0 24922 7 1 2 75310 82323
0 24923 5 1 1 24922
0 24924 7 1 2 24921 24923
0 24925 7 1 2 24915 24924
0 24926 5 1 1 24925
0 24927 7 1 2 70174 24926
0 24928 5 1 1 24927
0 24929 7 1 2 82553 90773
0 24930 5 1 1 24929
0 24931 7 1 2 89502 24930
0 24932 5 1 1 24931
0 24933 7 1 2 81695 24932
0 24934 5 1 1 24933
0 24935 7 1 2 83498 24934
0 24936 7 1 2 24928 24935
0 24937 7 1 2 24911 24936
0 24938 7 1 2 24887 24937
0 24939 5 1 1 24938
0 24940 7 1 2 62999 24939
0 24941 5 1 1 24940
0 24942 7 1 2 67634 93124
0 24943 5 1 1 24942
0 24944 7 1 2 69917 76975
0 24945 5 2 1 24944
0 24946 7 2 2 71781 93317
0 24947 5 2 1 93319
0 24948 7 1 2 70901 93320
0 24949 5 1 1 24948
0 24950 7 1 2 67319 77749
0 24951 7 1 2 24949 24950
0 24952 5 1 1 24951
0 24953 7 1 2 66493 24952
0 24954 7 1 2 24943 24953
0 24955 5 1 1 24954
0 24956 7 1 2 61533 73772
0 24957 5 1 1 24956
0 24958 7 1 2 67993 24957
0 24959 7 1 2 24955 24958
0 24960 5 1 1 24959
0 24961 7 1 2 24941 24960
0 24962 5 1 1 24961
0 24963 7 1 2 66690 24962
0 24964 5 1 1 24963
0 24965 7 1 2 65199 71852
0 24966 5 2 1 24965
0 24967 7 1 2 71290 93323
0 24968 5 1 1 24967
0 24969 7 1 2 61072 82879
0 24970 5 1 1 24969
0 24971 7 1 2 66494 24970
0 24972 7 1 2 24968 24971
0 24973 5 1 1 24972
0 24974 7 1 2 70924 79536
0 24975 7 1 2 71309 24974
0 24976 5 1 1 24975
0 24977 7 1 2 24973 24976
0 24978 5 1 1 24977
0 24979 7 1 2 76775 85100
0 24980 5 1 1 24979
0 24981 7 1 2 89503 24980
0 24982 7 1 2 24978 24981
0 24983 5 1 1 24982
0 24984 7 1 2 85365 86842
0 24985 7 1 2 24983 24984
0 24986 5 1 1 24985
0 24987 7 1 2 79287 88106
0 24988 5 1 1 24987
0 24989 7 1 2 81356 78699
0 24990 5 1 1 24989
0 24991 7 1 2 24988 24990
0 24992 5 1 1 24991
0 24993 7 1 2 64506 24992
0 24994 5 1 1 24993
0 24995 7 6 2 64964 77145
0 24996 7 1 2 81727 93325
0 24997 5 1 1 24996
0 24998 7 1 2 24994 24997
0 24999 7 1 2 24986 24998
0 25000 5 1 1 24999
0 25001 7 1 2 62649 25000
0 25002 5 1 1 25001
0 25003 7 3 2 77295 86362
0 25004 7 1 2 88547 93331
0 25005 5 1 1 25004
0 25006 7 1 2 61534 85175
0 25007 5 1 1 25006
0 25008 7 1 2 25005 25007
0 25009 5 1 1 25008
0 25010 7 1 2 64726 25009
0 25011 5 1 1 25010
0 25012 7 1 2 77357 11645
0 25013 5 1 1 25012
0 25014 7 1 2 76822 25013
0 25015 5 1 1 25014
0 25016 7 1 2 70798 82907
0 25017 5 1 1 25016
0 25018 7 1 2 25015 25017
0 25019 5 1 1 25018
0 25020 7 1 2 81357 25019
0 25021 5 1 1 25020
0 25022 7 1 2 72193 70262
0 25023 5 1 1 25022
0 25024 7 1 2 93128 25023
0 25025 5 1 1 25024
0 25026 7 1 2 79288 91482
0 25027 7 1 2 25025 25026
0 25028 5 1 1 25027
0 25029 7 1 2 25021 25028
0 25030 5 1 1 25029
0 25031 7 1 2 62099 25030
0 25032 5 1 1 25031
0 25033 7 1 2 25011 25032
0 25034 7 1 2 25002 25033
0 25035 7 1 2 24964 25034
0 25036 5 1 1 25035
0 25037 7 1 2 68345 25036
0 25038 5 1 1 25037
0 25039 7 4 2 75799 88454
0 25040 5 2 1 93334
0 25041 7 1 2 90846 93338
0 25042 5 1 1 25041
0 25043 7 1 2 76776 25042
0 25044 5 1 1 25043
0 25045 7 1 2 91138 93335
0 25046 5 1 1 25045
0 25047 7 1 2 82266 70245
0 25048 5 1 1 25047
0 25049 7 1 2 76777 81696
0 25050 5 1 1 25049
0 25051 7 1 2 25048 25050
0 25052 5 1 1 25051
0 25053 7 1 2 74527 25052
0 25054 5 1 1 25053
0 25055 7 1 2 25046 25054
0 25056 7 1 2 25044 25055
0 25057 5 1 1 25056
0 25058 7 1 2 61535 25057
0 25059 5 1 1 25058
0 25060 7 1 2 67635 93015
0 25061 5 1 1 25060
0 25062 7 1 2 77640 88821
0 25063 7 1 2 93012 25062
0 25064 5 1 1 25063
0 25065 7 1 2 25061 25064
0 25066 5 1 1 25065
0 25067 7 1 2 71723 25066
0 25068 5 1 1 25067
0 25069 7 2 2 77633 90490
0 25070 5 1 1 93340
0 25071 7 1 2 25068 25070
0 25072 5 1 1 25071
0 25073 7 1 2 59334 25072
0 25074 5 1 1 25073
0 25075 7 2 2 73061 88992
0 25076 5 1 1 93342
0 25077 7 1 2 82267 93343
0 25078 5 1 1 25077
0 25079 7 1 2 25074 25078
0 25080 5 1 1 25079
0 25081 7 1 2 61536 25080
0 25082 5 1 1 25081
0 25083 7 1 2 79954 72145
0 25084 7 1 2 88359 25083
0 25085 5 1 1 25084
0 25086 7 1 2 61537 25085
0 25087 5 1 1 25086
0 25088 7 2 2 69563 89488
0 25089 5 1 1 93344
0 25090 7 1 2 67320 93345
0 25091 5 1 1 25090
0 25092 7 1 2 25087 25091
0 25093 5 1 1 25092
0 25094 7 1 2 67636 25093
0 25095 5 1 1 25094
0 25096 7 1 2 74595 93013
0 25097 5 1 1 25096
0 25098 7 1 2 80498 93017
0 25099 7 1 2 25097 25098
0 25100 5 1 1 25099
0 25101 7 1 2 59335 25100
0 25102 5 1 1 25101
0 25103 7 1 2 61073 86951
0 25104 5 1 1 25103
0 25105 7 1 2 73069 25104
0 25106 5 1 1 25105
0 25107 7 1 2 59897 25106
0 25108 5 1 1 25107
0 25109 7 1 2 25076 25108
0 25110 7 1 2 25102 25109
0 25111 5 1 1 25110
0 25112 7 1 2 61538 25111
0 25113 5 1 1 25112
0 25114 7 1 2 25095 25113
0 25115 5 1 1 25114
0 25116 7 1 2 70175 25115
0 25117 5 1 1 25116
0 25118 7 1 2 72629 92240
0 25119 5 1 1 25118
0 25120 7 1 2 75311 88906
0 25121 5 1 1 25120
0 25122 7 1 2 25119 25121
0 25123 5 1 1 25122
0 25124 7 1 2 70176 25123
0 25125 5 1 1 25124
0 25126 7 1 2 89286 89588
0 25127 5 2 1 25126
0 25128 7 1 2 25125 93346
0 25129 5 1 1 25128
0 25130 7 1 2 70531 25129
0 25131 5 1 1 25130
0 25132 7 1 2 81434 88878
0 25133 5 1 1 25132
0 25134 7 1 2 66495 25133
0 25135 5 1 1 25134
0 25136 7 1 2 72112 25135
0 25137 5 1 1 25136
0 25138 7 1 2 66496 83693
0 25139 5 3 1 25138
0 25140 7 1 2 71220 93348
0 25141 5 1 1 25140
0 25142 7 1 2 66497 24913
0 25143 5 2 1 25142
0 25144 7 1 2 70532 93351
0 25145 5 1 1 25144
0 25146 7 1 2 61539 82143
0 25147 5 1 1 25146
0 25148 7 1 2 59336 93341
0 25149 5 1 1 25148
0 25150 7 1 2 25147 25149
0 25151 7 1 2 25145 25150
0 25152 7 1 2 25141 25151
0 25153 7 1 2 25137 25152
0 25154 5 1 1 25153
0 25155 7 1 2 76778 25154
0 25156 5 1 1 25155
0 25157 7 1 2 70614 86967
0 25158 5 2 1 25157
0 25159 7 1 2 59898 91961
0 25160 5 1 1 25159
0 25161 7 1 2 70177 92241
0 25162 5 1 1 25161
0 25163 7 1 2 19571 25162
0 25164 7 1 2 25160 25163
0 25165 5 1 1 25164
0 25166 7 1 2 81438 25165
0 25167 5 1 1 25166
0 25168 7 1 2 93353 25167
0 25169 7 1 2 25156 25168
0 25170 7 1 2 25131 25169
0 25171 7 1 2 25117 25170
0 25172 7 1 2 25082 25171
0 25173 5 1 1 25172
0 25174 7 1 2 67994 25173
0 25175 5 1 1 25174
0 25176 7 1 2 25059 25175
0 25177 5 1 1 25176
0 25178 7 1 2 85677 25177
0 25179 5 1 1 25178
0 25180 7 1 2 25038 25179
0 25181 5 1 1 25180
0 25182 7 1 2 65408 25181
0 25183 5 1 1 25182
0 25184 7 4 2 64727 60532
0 25185 7 1 2 85366 93355
0 25186 7 1 2 80477 25185
0 25187 5 1 1 25186
0 25188 7 1 2 59899 79217
0 25189 5 1 1 25188
0 25190 7 1 2 66267 25189
0 25191 5 1 1 25190
0 25192 7 1 2 69918 73356
0 25193 5 1 1 25192
0 25194 7 2 2 75039 25193
0 25195 7 2 2 62307 93359
0 25196 7 1 2 76704 93361
0 25197 5 1 1 25196
0 25198 7 1 2 25191 25197
0 25199 5 1 1 25198
0 25200 7 8 2 64965 73791
0 25201 5 7 1 93363
0 25202 7 1 2 79259 93364
0 25203 7 1 2 25199 25202
0 25204 5 1 1 25203
0 25205 7 1 2 25187 25204
0 25206 5 1 1 25205
0 25207 7 1 2 89217 25206
0 25208 5 1 1 25207
0 25209 7 1 2 63739 25208
0 25210 7 1 2 25183 25209
0 25211 7 1 2 24865 25210
0 25212 5 1 1 25211
0 25213 7 1 2 66268 2429
0 25214 5 1 1 25213
0 25215 7 1 2 83072 73773
0 25216 5 1 1 25215
0 25217 7 1 2 59550 25216
0 25218 5 1 1 25217
0 25219 7 1 2 3655 89072
0 25220 5 1 1 25219
0 25221 7 1 2 69919 25220
0 25222 5 1 1 25221
0 25223 7 2 2 60351 76874
0 25224 5 1 1 93378
0 25225 7 1 2 61341 25224
0 25226 5 1 1 25225
0 25227 7 1 2 82747 25226
0 25228 7 1 2 25222 25227
0 25229 7 1 2 25218 25228
0 25230 7 1 2 25214 25229
0 25231 5 1 1 25230
0 25232 7 1 2 77903 25231
0 25233 5 1 1 25232
0 25234 7 1 2 76823 90854
0 25235 5 1 1 25234
0 25236 7 1 2 77981 25235
0 25237 5 1 1 25236
0 25238 7 1 2 71431 25237
0 25239 5 1 1 25238
0 25240 7 1 2 60352 93371
0 25241 5 7 1 25240
0 25242 7 1 2 77317 93380
0 25243 5 1 1 25242
0 25244 7 1 2 72767 81324
0 25245 5 1 1 25244
0 25246 7 4 2 62650 70054
0 25247 5 1 1 93387
0 25248 7 1 2 65857 87878
0 25249 5 1 1 25248
0 25250 7 1 2 25247 25249
0 25251 5 1 1 25250
0 25252 7 1 2 69806 25251
0 25253 5 1 1 25252
0 25254 7 1 2 25245 25253
0 25255 7 1 2 25243 25254
0 25256 5 1 1 25255
0 25257 7 1 2 64507 25256
0 25258 5 1 1 25257
0 25259 7 1 2 60353 78046
0 25260 5 1 1 25259
0 25261 7 1 2 64728 25260
0 25262 5 1 1 25261
0 25263 7 2 2 60354 73822
0 25264 5 1 1 93391
0 25265 7 1 2 66269 25264
0 25266 5 1 1 25265
0 25267 7 1 2 25262 25266
0 25268 5 1 1 25267
0 25269 7 1 2 64966 25268
0 25270 5 1 1 25269
0 25271 7 1 2 25258 25270
0 25272 7 1 2 25239 25271
0 25273 5 1 1 25272
0 25274 7 1 2 68346 25273
0 25275 5 1 1 25274
0 25276 7 1 2 25233 25275
0 25277 5 1 1 25276
0 25278 7 1 2 66498 25277
0 25279 5 1 1 25278
0 25280 7 1 2 81139 70936
0 25281 5 1 1 25280
0 25282 7 1 2 67995 76083
0 25283 5 1 1 25282
0 25284 7 1 2 81055 25283
0 25285 5 1 1 25284
0 25286 7 1 2 79537 25285
0 25287 5 1 1 25286
0 25288 7 1 2 25281 25287
0 25289 5 1 1 25288
0 25290 7 1 2 63442 25289
0 25291 5 1 1 25290
0 25292 7 1 2 86916 93252
0 25293 5 1 1 25292
0 25294 7 1 2 69807 25293
0 25295 5 1 1 25294
0 25296 7 1 2 66023 91035
0 25297 5 1 1 25296
0 25298 7 1 2 25295 25297
0 25299 5 1 1 25298
0 25300 7 1 2 62651 25299
0 25301 5 1 1 25300
0 25302 7 1 2 77323 78897
0 25303 5 1 1 25302
0 25304 7 1 2 77706 25303
0 25305 5 1 1 25304
0 25306 7 1 2 25301 25305
0 25307 5 1 1 25306
0 25308 7 1 2 75067 25307
0 25309 5 1 1 25308
0 25310 7 1 2 67637 78681
0 25311 5 1 1 25310
0 25312 7 1 2 12044 25311
0 25313 5 1 1 25312
0 25314 7 1 2 81949 25313
0 25315 5 1 1 25314
0 25316 7 1 2 25309 25315
0 25317 5 1 1 25316
0 25318 7 1 2 64967 25317
0 25319 5 1 1 25318
0 25320 7 1 2 25291 25319
0 25321 7 1 2 25279 25320
0 25322 5 1 1 25321
0 25323 7 1 2 66691 25322
0 25324 5 1 1 25323
0 25325 7 1 2 82821 82341
0 25326 5 1 1 25325
0 25327 7 1 2 25324 25326
0 25328 5 1 1 25327
0 25329 7 1 2 65409 25328
0 25330 5 1 1 25329
0 25331 7 1 2 75573 88193
0 25332 5 1 1 25331
0 25333 7 1 2 65858 93088
0 25334 5 1 1 25333
0 25335 7 1 2 64729 87549
0 25336 5 1 1 25335
0 25337 7 1 2 25334 25336
0 25338 5 1 1 25337
0 25339 7 1 2 66270 92415
0 25340 7 1 2 25338 25339
0 25341 5 1 1 25340
0 25342 7 1 2 25332 25341
0 25343 5 1 1 25342
0 25344 7 1 2 64968 25343
0 25345 5 1 1 25344
0 25346 7 3 2 65859 75574
0 25347 7 1 2 76467 88194
0 25348 7 1 2 93393 25347
0 25349 5 1 1 25348
0 25350 7 1 2 25345 25349
0 25351 5 1 1 25350
0 25352 7 1 2 66024 25351
0 25353 5 1 1 25352
0 25354 7 1 2 85245 90821
0 25355 5 1 1 25354
0 25356 7 1 2 69808 25355
0 25357 5 1 1 25356
0 25358 7 1 2 82122 25357
0 25359 5 1 1 25358
0 25360 7 1 2 64730 25359
0 25361 5 1 1 25360
0 25362 7 1 2 75920 88318
0 25363 5 1 1 25362
0 25364 7 1 2 25361 25363
0 25365 5 1 1 25364
0 25366 7 1 2 75575 25365
0 25367 5 1 1 25366
0 25368 7 1 2 76209 82738
0 25369 5 1 1 25368
0 25370 7 1 2 79408 25369
0 25371 5 1 1 25370
0 25372 7 1 2 25367 25371
0 25373 5 1 1 25372
0 25374 7 1 2 66692 25373
0 25375 5 1 1 25374
0 25376 7 1 2 25353 25375
0 25377 5 1 1 25376
0 25378 7 1 2 65410 25377
0 25379 5 1 1 25378
0 25380 7 1 2 73885 82324
0 25381 5 1 1 25380
0 25382 7 1 2 66693 84580
0 25383 7 1 2 87576 25382
0 25384 7 1 2 25381 25383
0 25385 5 1 1 25384
0 25386 7 1 2 68347 25385
0 25387 7 1 2 25379 25386
0 25388 5 1 1 25387
0 25389 7 1 2 81697 93049
0 25390 5 1 1 25389
0 25391 7 1 2 88848 93058
0 25392 5 1 1 25391
0 25393 7 1 2 66499 90500
0 25394 7 1 2 88876 25393
0 25395 7 1 2 25392 25394
0 25396 7 1 2 25390 25395
0 25397 5 1 1 25396
0 25398 7 1 2 61540 93372
0 25399 5 4 1 25398
0 25400 7 1 2 79613 93396
0 25401 7 1 2 25397 25400
0 25402 5 1 1 25401
0 25403 7 1 2 83724 93060
0 25404 5 1 1 25403
0 25405 7 2 2 76824 77318
0 25406 5 2 1 93400
0 25407 7 1 2 73567 84073
0 25408 5 1 1 25407
0 25409 7 1 2 93402 25408
0 25410 5 1 1 25409
0 25411 7 1 2 3460 80345
0 25412 5 5 1 25411
0 25413 7 1 2 93326 93404
0 25414 7 1 2 25410 25413
0 25415 5 1 1 25414
0 25416 7 1 2 25404 25415
0 25417 5 1 1 25416
0 25418 7 1 2 66271 25417
0 25419 5 1 1 25418
0 25420 7 1 2 63443 25419
0 25421 7 1 2 25402 25420
0 25422 5 1 1 25421
0 25423 7 1 2 63000 25422
0 25424 7 1 2 25388 25423
0 25425 5 1 1 25424
0 25426 7 2 2 64731 82342
0 25427 5 1 1 93409
0 25428 7 1 2 81325 86057
0 25429 7 1 2 93410 25428
0 25430 5 1 1 25429
0 25431 7 1 2 68673 25430
0 25432 7 1 2 25425 25431
0 25433 7 1 2 25330 25432
0 25434 5 1 1 25433
0 25435 7 1 2 63969 25434
0 25436 7 1 2 25212 25435
0 25437 5 1 1 25436
0 25438 7 1 2 77833 78282
0 25439 5 1 1 25438
0 25440 7 1 2 89537 25439
0 25441 5 1 1 25440
0 25442 7 1 2 73099 25441
0 25443 5 1 1 25442
0 25444 7 1 2 85157 89626
0 25445 5 1 1 25444
0 25446 7 1 2 62652 25445
0 25447 5 1 1 25446
0 25448 7 1 2 25443 25447
0 25449 5 1 1 25448
0 25450 7 1 2 63444 25449
0 25451 5 1 1 25450
0 25452 7 1 2 73100 93397
0 25453 5 1 1 25452
0 25454 7 1 2 81945 25453
0 25455 5 1 1 25454
0 25456 7 1 2 85615 25455
0 25457 5 1 1 25456
0 25458 7 1 2 25451 25457
0 25459 5 1 1 25458
0 25460 7 1 2 84341 25459
0 25461 5 1 1 25460
0 25462 7 1 2 73167 77781
0 25463 5 2 1 25462
0 25464 7 1 2 73101 82343
0 25465 5 1 1 25464
0 25466 7 1 2 93411 25465
0 25467 5 1 1 25466
0 25468 7 1 2 61717 8701
0 25469 5 1 1 25468
0 25470 7 1 2 25467 25469
0 25471 5 1 1 25470
0 25472 7 1 2 64969 91318
0 25473 5 1 1 25472
0 25474 7 1 2 61718 25473
0 25475 5 1 1 25474
0 25476 7 1 2 73102 85967
0 25477 7 1 2 25475 25476
0 25478 5 1 1 25477
0 25479 7 1 2 25471 25478
0 25480 5 1 1 25479
0 25481 7 1 2 68674 25480
0 25482 5 1 1 25481
0 25483 7 2 2 64732 76886
0 25484 5 1 1 93413
0 25485 7 2 2 64970 76867
0 25486 5 1 1 93415
0 25487 7 1 2 25484 25486
0 25488 5 1 1 25487
0 25489 7 1 2 80197 84478
0 25490 7 1 2 25488 25489
0 25491 5 1 1 25490
0 25492 7 1 2 25482 25491
0 25493 5 1 1 25492
0 25494 7 1 2 62100 25493
0 25495 5 1 1 25494
0 25496 7 3 2 81536 78700
0 25497 5 1 1 93417
0 25498 7 1 2 84257 93418
0 25499 5 1 1 25498
0 25500 7 1 2 77324 76875
0 25501 5 1 1 25500
0 25502 7 1 2 75844 25501
0 25503 5 1 1 25502
0 25504 7 1 2 83162 25503
0 25505 5 1 1 25504
0 25506 7 1 2 84342 25505
0 25507 5 1 1 25506
0 25508 7 1 2 25499 25507
0 25509 7 1 2 25495 25508
0 25510 5 1 1 25509
0 25511 7 1 2 65200 25510
0 25512 5 1 1 25511
0 25513 7 1 2 25461 25512
0 25514 5 1 1 25513
0 25515 7 1 2 65411 25514
0 25516 5 1 1 25515
0 25517 7 5 2 63001 89927
0 25518 7 1 2 84300 93420
0 25519 5 1 1 25518
0 25520 7 1 2 61719 90676
0 25521 5 1 1 25520
0 25522 7 1 2 25519 25521
0 25523 5 1 1 25522
0 25524 7 1 2 78084 25523
0 25525 5 1 1 25524
0 25526 7 1 2 80866 88272
0 25527 5 1 1 25526
0 25528 7 1 2 25525 25527
0 25529 5 1 1 25528
0 25530 7 1 2 65201 25529
0 25531 5 1 1 25530
0 25532 7 5 2 64971 60533
0 25533 7 1 2 84252 93425
0 25534 7 1 2 85834 25533
0 25535 5 1 1 25534
0 25536 7 1 2 25531 25535
0 25537 5 1 1 25536
0 25538 7 1 2 66272 25537
0 25539 5 1 1 25538
0 25540 7 1 2 74481 79289
0 25541 5 1 1 25540
0 25542 7 1 2 78701 79538
0 25543 7 1 2 88226 25542
0 25544 5 1 1 25543
0 25545 7 1 2 25541 25544
0 25546 5 1 1 25545
0 25547 7 1 2 90677 25546
0 25548 5 1 1 25547
0 25549 7 1 2 25539 25548
0 25550 5 1 1 25549
0 25551 7 1 2 66500 25550
0 25552 5 1 1 25551
0 25553 7 2 2 74367 84409
0 25554 5 1 1 93430
0 25555 7 1 2 78932 85198
0 25556 7 2 2 93431 25555
0 25557 5 1 1 93432
0 25558 7 1 2 65202 93433
0 25559 5 1 1 25558
0 25560 7 1 2 25552 25559
0 25561 7 1 2 25516 25560
0 25562 5 1 1 25561
0 25563 7 1 2 63970 25562
0 25564 5 1 1 25563
0 25565 7 2 2 81782 91997
0 25566 7 1 2 82908 93365
0 25567 7 1 2 85384 25566
0 25568 7 1 2 93434 25567
0 25569 5 1 1 25568
0 25570 7 1 2 25564 25569
0 25571 5 1 1 25570
0 25572 7 1 2 72550 25571
0 25573 5 1 1 25572
0 25574 7 1 2 87656 90852
0 25575 5 1 1 25574
0 25576 7 1 2 75576 93206
0 25577 5 1 1 25576
0 25578 7 2 2 75312 25577
0 25579 5 5 1 93436
0 25580 7 1 2 63002 93438
0 25581 7 1 2 93193 25580
0 25582 5 1 1 25581
0 25583 7 1 2 25575 25582
0 25584 5 1 1 25583
0 25585 7 1 2 66273 25584
0 25586 5 1 1 25585
0 25587 7 1 2 63003 71432
0 25588 5 1 1 25587
0 25589 7 1 2 93403 25588
0 25590 5 1 1 25589
0 25591 7 1 2 92945 25590
0 25592 5 1 1 25591
0 25593 7 1 2 25586 25592
0 25594 5 1 1 25593
0 25595 7 1 2 80688 79039
0 25596 7 1 2 25594 25595
0 25597 5 1 1 25596
0 25598 7 1 2 61862 25597
0 25599 7 1 2 25573 25598
0 25600 7 1 2 25437 25599
0 25601 5 1 1 25600
0 25602 7 1 2 65563 25601
0 25603 7 1 2 24716 25602
0 25604 5 1 1 25603
0 25605 7 1 2 73235 89601
0 25606 5 2 1 25605
0 25607 7 1 2 60534 93443
0 25608 5 1 1 25607
0 25609 7 1 2 93287 25608
0 25610 5 1 1 25609
0 25611 7 1 2 66501 25610
0 25612 5 1 1 25611
0 25613 7 1 2 76362 73249
0 25614 5 1 1 25613
0 25615 7 1 2 91939 25614
0 25616 5 1 1 25615
0 25617 7 1 2 80462 73307
0 25618 5 1 1 25617
0 25619 7 1 2 61074 90774
0 25620 7 1 2 25618 25619
0 25621 5 1 1 25620
0 25622 7 1 2 6641 25621
0 25623 5 1 1 25622
0 25624 7 1 2 60924 25623
0 25625 5 1 1 25624
0 25626 7 1 2 25616 25625
0 25627 5 1 1 25626
0 25628 7 1 2 67321 25627
0 25629 5 1 1 25628
0 25630 7 1 2 80636 91462
0 25631 5 1 1 25630
0 25632 7 1 2 66502 25631
0 25633 5 1 1 25632
0 25634 7 1 2 60153 25633
0 25635 5 1 1 25634
0 25636 7 2 2 60802 76499
0 25637 7 1 2 89489 93445
0 25638 5 1 1 25637
0 25639 7 1 2 74688 25638
0 25640 7 1 2 25635 25639
0 25641 5 1 1 25640
0 25642 7 1 2 59337 25641
0 25643 5 1 1 25642
0 25644 7 1 2 60803 74652
0 25645 5 1 1 25644
0 25646 7 1 2 25643 25645
0 25647 5 1 1 25646
0 25648 7 1 2 71601 25647
0 25649 5 1 1 25648
0 25650 7 1 2 92243 25089
0 25651 5 1 1 25650
0 25652 7 1 2 72113 25651
0 25653 5 1 1 25652
0 25654 7 1 2 79955 72340
0 25655 5 1 1 25654
0 25656 7 1 2 61541 25655
0 25657 5 1 1 25656
0 25658 7 1 2 25653 25657
0 25659 5 1 1 25658
0 25660 7 1 2 70178 25659
0 25661 5 1 1 25660
0 25662 7 1 2 20024 22276
0 25663 5 2 1 25662
0 25664 7 1 2 70533 93447
0 25665 5 1 1 25664
0 25666 7 2 2 61542 72573
0 25667 5 1 1 93449
0 25668 7 1 2 73207 25667
0 25669 5 1 1 25668
0 25670 7 1 2 71443 90775
0 25671 7 1 2 25669 25670
0 25672 5 1 1 25671
0 25673 7 1 2 83499 25672
0 25674 7 1 2 25665 25673
0 25675 7 1 2 25661 25674
0 25676 7 1 2 25649 25675
0 25677 7 1 2 25629 25676
0 25678 5 1 1 25677
0 25679 7 1 2 65412 25678
0 25680 5 1 1 25679
0 25681 7 1 2 25612 25680
0 25682 5 1 1 25681
0 25683 7 1 2 67638 25682
0 25684 5 1 1 25683
0 25685 7 1 2 61075 5810
0 25686 5 1 1 25685
0 25687 7 1 2 59900 70437
0 25688 5 1 1 25687
0 25689 7 1 2 73072 25688
0 25690 7 1 2 25686 25689
0 25691 5 1 1 25690
0 25692 7 1 2 4061 83712
0 25693 5 1 1 25692
0 25694 7 1 2 70179 25693
0 25695 7 1 2 25691 25694
0 25696 5 1 1 25695
0 25697 7 1 2 79827 91784
0 25698 7 1 2 88598 25697
0 25699 5 1 1 25698
0 25700 7 2 2 70281 69187
0 25701 5 1 1 93451
0 25702 7 1 2 75794 93452
0 25703 7 1 2 89761 25702
0 25704 5 1 1 25703
0 25705 7 1 2 25699 25704
0 25706 5 1 1 25705
0 25707 7 1 2 59338 25706
0 25708 5 1 1 25707
0 25709 7 1 2 73721 92390
0 25710 5 1 1 25709
0 25711 7 2 2 65413 92410
0 25712 5 2 1 93453
0 25713 7 1 2 25710 93455
0 25714 5 1 1 25713
0 25715 7 1 2 80309 92712
0 25716 5 1 1 25715
0 25717 7 1 2 25714 25716
0 25718 5 1 1 25717
0 25719 7 1 2 25708 25718
0 25720 7 1 2 25696 25719
0 25721 7 1 2 25684 25720
0 25722 5 1 1 25721
0 25723 7 1 2 67996 25722
0 25724 5 1 1 25723
0 25725 7 1 2 60355 79484
0 25726 5 1 1 25725
0 25727 7 1 2 83713 25726
0 25728 5 4 1 25727
0 25729 7 1 2 70615 93457
0 25730 5 1 1 25729
0 25731 7 1 2 82700 25730
0 25732 5 1 1 25731
0 25733 7 1 2 82062 25732
0 25734 5 1 1 25733
0 25735 7 1 2 81370 93458
0 25736 5 1 1 25735
0 25737 7 2 2 61543 75970
0 25738 7 1 2 81393 93461
0 25739 5 1 1 25738
0 25740 7 1 2 25736 25739
0 25741 5 1 1 25740
0 25742 7 1 2 71491 25741
0 25743 5 1 1 25742
0 25744 7 1 2 25734 25743
0 25745 5 1 1 25744
0 25746 7 1 2 73823 25745
0 25747 5 1 1 25746
0 25748 7 1 2 60154 93459
0 25749 7 1 2 83456 25748
0 25750 5 1 1 25749
0 25751 7 1 2 88740 25750
0 25752 5 1 1 25751
0 25753 7 1 2 76148 25752
0 25754 5 1 1 25753
0 25755 7 1 2 64972 83453
0 25756 5 1 1 25755
0 25757 7 1 2 82228 88741
0 25758 5 1 1 25757
0 25759 7 1 2 93460 25758
0 25760 7 1 2 25756 25759
0 25761 5 1 1 25760
0 25762 7 1 2 25754 25761
0 25763 7 1 2 25747 25762
0 25764 7 1 2 25724 25763
0 25765 5 1 1 25764
0 25766 7 1 2 63445 25765
0 25767 5 1 1 25766
0 25768 7 1 2 78331 91978
0 25769 5 1 1 25768
0 25770 7 1 2 66503 81474
0 25771 5 1 1 25770
0 25772 7 1 2 25769 25771
0 25773 5 1 1 25772
0 25774 7 1 2 69920 25773
0 25775 5 1 1 25774
0 25776 7 2 2 79850 72474
0 25777 5 1 1 93463
0 25778 7 1 2 67322 93464
0 25779 5 1 1 25778
0 25780 7 1 2 81824 25779
0 25781 5 1 1 25780
0 25782 7 1 2 66504 25781
0 25783 5 1 1 25782
0 25784 7 1 2 25775 25783
0 25785 5 1 1 25784
0 25786 7 1 2 70180 25785
0 25787 5 1 1 25786
0 25788 7 1 2 62653 80328
0 25789 5 1 1 25788
0 25790 7 1 2 25787 25789
0 25791 5 1 1 25790
0 25792 7 1 2 67997 25791
0 25793 5 1 1 25792
0 25794 7 3 2 60925 82863
0 25795 7 1 2 74972 93465
0 25796 5 1 1 25795
0 25797 7 2 2 70181 82410
0 25798 5 1 1 93468
0 25799 7 1 2 16823 93469
0 25800 5 1 1 25799
0 25801 7 1 2 73191 93257
0 25802 5 1 1 25801
0 25803 7 1 2 25800 25802
0 25804 5 1 1 25803
0 25805 7 1 2 72114 25804
0 25806 5 1 1 25805
0 25807 7 1 2 25796 25806
0 25808 7 1 2 25793 25807
0 25809 5 1 1 25808
0 25810 7 1 2 71221 25809
0 25811 5 1 1 25810
0 25812 7 2 2 77689 743
0 25813 5 1 1 93470
0 25814 7 1 2 65203 88432
0 25815 7 1 2 77723 25814
0 25816 7 1 2 92938 25815
0 25817 7 1 2 93471 25816
0 25818 5 1 1 25817
0 25819 7 1 2 63004 25818
0 25820 5 1 1 25819
0 25821 7 1 2 67323 93140
0 25822 5 1 1 25821
0 25823 7 1 2 78004 84017
0 25824 5 1 1 25823
0 25825 7 1 2 76641 25824
0 25826 5 1 1 25825
0 25827 7 1 2 25822 25826
0 25828 5 1 1 25827
0 25829 7 1 2 67998 25828
0 25830 5 1 1 25829
0 25831 7 1 2 76689 25830
0 25832 7 1 2 25820 25831
0 25833 5 1 1 25832
0 25834 7 1 2 61544 25833
0 25835 5 1 1 25834
0 25836 7 1 2 83321 93101
0 25837 5 1 1 25836
0 25838 7 1 2 63005 90356
0 25839 5 1 1 25838
0 25840 7 1 2 25837 25839
0 25841 5 1 1 25840
0 25842 7 1 2 73507 25841
0 25843 5 1 1 25842
0 25844 7 1 2 90043 24622
0 25845 5 1 1 25844
0 25846 7 1 2 70182 25845
0 25847 5 1 1 25846
0 25848 7 1 2 72146 93262
0 25849 5 1 1 25848
0 25850 7 1 2 59551 25849
0 25851 5 1 1 25850
0 25852 7 1 2 88972 25851
0 25853 5 1 1 25852
0 25854 7 1 2 92741 25853
0 25855 5 1 1 25854
0 25856 7 1 2 25847 25855
0 25857 5 1 1 25856
0 25858 7 1 2 69125 25857
0 25859 5 1 1 25858
0 25860 7 1 2 25843 25859
0 25861 7 1 2 25835 25860
0 25862 7 1 2 59901 93138
0 25863 5 1 1 25862
0 25864 7 1 2 79156 92742
0 25865 5 1 1 25864
0 25866 7 1 2 25863 25865
0 25867 5 1 1 25866
0 25868 7 1 2 59339 25867
0 25869 5 1 1 25868
0 25870 7 1 2 60804 82481
0 25871 5 1 1 25870
0 25872 7 1 2 83213 25871
0 25873 5 1 1 25872
0 25874 7 1 2 92743 25873
0 25875 5 1 1 25874
0 25876 7 1 2 25869 25875
0 25877 5 1 1 25876
0 25878 7 1 2 71602 25877
0 25879 5 1 1 25878
0 25880 7 1 2 75313 70985
0 25881 5 1 1 25880
0 25882 7 1 2 76927 91508
0 25883 5 1 1 25882
0 25884 7 1 2 25881 25883
0 25885 5 1 1 25884
0 25886 7 1 2 63006 25885
0 25887 5 1 1 25886
0 25888 7 1 2 82460 91501
0 25889 5 1 1 25888
0 25890 7 1 2 25887 25889
0 25891 5 1 1 25890
0 25892 7 1 2 247 25891
0 25893 5 1 1 25892
0 25894 7 1 2 63007 25813
0 25895 5 1 1 25894
0 25896 7 1 2 77718 85066
0 25897 7 1 2 92176 25896
0 25898 5 1 1 25897
0 25899 7 1 2 71310 88333
0 25900 5 1 1 25899
0 25901 7 1 2 78888 25900
0 25902 5 1 1 25901
0 25903 7 1 2 25898 25902
0 25904 7 1 2 25895 25903
0 25905 5 1 1 25904
0 25906 7 1 2 60356 25905
0 25907 5 1 1 25906
0 25908 7 1 2 75205 255
0 25909 5 1 1 25908
0 25910 7 1 2 62101 89156
0 25911 5 1 1 25910
0 25912 7 1 2 69921 25911
0 25913 5 1 1 25912
0 25914 7 1 2 64508 25913
0 25915 5 1 1 25914
0 25916 7 1 2 63008 82292
0 25917 7 1 2 25915 25916
0 25918 5 1 1 25917
0 25919 7 1 2 91487 25918
0 25920 5 1 1 25919
0 25921 7 1 2 25909 25920
0 25922 5 1 1 25921
0 25923 7 1 2 66505 76674
0 25924 5 3 1 25923
0 25925 7 1 2 89073 93472
0 25926 7 1 2 93134 25925
0 25927 5 2 1 25926
0 25928 7 1 2 87758 93475
0 25929 5 1 1 25928
0 25930 7 1 2 83026 93476
0 25931 5 1 1 25930
0 25932 7 1 2 83002 88430
0 25933 5 1 1 25932
0 25934 7 1 2 25931 25933
0 25935 5 1 1 25934
0 25936 7 1 2 72229 25935
0 25937 5 1 1 25936
0 25938 7 1 2 25929 25937
0 25939 7 1 2 25922 25938
0 25940 7 1 2 25907 25939
0 25941 7 1 2 25893 25940
0 25942 7 1 2 25879 25941
0 25943 7 1 2 25861 25942
0 25944 7 1 2 25811 25943
0 25945 5 1 1 25944
0 25946 7 1 2 82173 25945
0 25947 5 1 1 25946
0 25948 7 1 2 63740 25947
0 25949 7 1 2 25767 25948
0 25950 5 1 1 25949
0 25951 7 1 2 82325 88849
0 25952 5 1 1 25951
0 25953 7 1 2 81698 74633
0 25954 5 1 1 25953
0 25955 7 1 2 25952 25954
0 25956 5 1 1 25955
0 25957 7 1 2 72115 25956
0 25958 5 1 1 25957
0 25959 7 1 2 81435 88851
0 25960 5 1 1 25959
0 25961 7 1 2 73824 76474
0 25962 5 1 1 25961
0 25963 7 1 2 74596 88842
0 25964 5 1 1 25963
0 25965 7 1 2 91123 25964
0 25966 7 1 2 25962 25965
0 25967 7 1 2 25960 25966
0 25968 7 1 2 25958 25967
0 25969 5 1 1 25968
0 25970 7 1 2 66274 90751
0 25971 5 1 1 25970
0 25972 7 1 2 81923 78728
0 25973 5 1 1 25972
0 25974 7 1 2 62654 25973
0 25975 5 1 1 25974
0 25976 7 1 2 72455 73623
0 25977 7 1 2 73679 25976
0 25978 5 1 1 25977
0 25979 7 1 2 67999 25978
0 25980 7 1 2 25975 25979
0 25981 7 1 2 25971 25980
0 25982 5 1 1 25981
0 25983 7 1 2 66506 25982
0 25984 7 1 2 25969 25983
0 25985 5 1 1 25984
0 25986 7 3 2 62308 89049
0 25987 5 1 1 93477
0 25988 7 1 2 64509 93478
0 25989 5 1 1 25988
0 25990 7 1 2 77358 25989
0 25991 5 1 1 25990
0 25992 7 1 2 74368 25991
0 25993 5 1 1 25992
0 25994 7 1 2 78967 87982
0 25995 5 1 1 25994
0 25996 7 1 2 81056 25995
0 25997 5 1 1 25996
0 25998 7 1 2 77191 25997
0 25999 5 1 1 25998
0 26000 7 1 2 74345 77431
0 26001 5 2 1 26000
0 26002 7 1 2 25999 93480
0 26003 7 1 2 25993 26002
0 26004 5 1 1 26003
0 26005 7 1 2 69809 26004
0 26006 5 1 1 26005
0 26007 7 1 2 77985 78253
0 26008 5 1 1 26007
0 26009 7 1 2 10493 26008
0 26010 5 1 1 26009
0 26011 7 1 2 64973 26010
0 26012 5 1 1 26011
0 26013 7 1 2 68000 75577
0 26014 7 1 2 82148 26013
0 26015 5 1 1 26014
0 26016 7 1 2 26012 26015
0 26017 5 1 1 26016
0 26018 7 1 2 66025 26017
0 26019 5 1 1 26018
0 26020 7 1 2 61545 74883
0 26021 5 1 1 26020
0 26022 7 1 2 89627 26021
0 26023 5 1 1 26022
0 26024 7 1 2 65204 26023
0 26025 5 1 1 26024
0 26026 7 1 2 81050 85564
0 26027 5 1 1 26026
0 26028 7 1 2 63446 26027
0 26029 7 1 2 26025 26028
0 26030 7 1 2 26019 26029
0 26031 7 1 2 26006 26030
0 26032 7 1 2 25985 26031
0 26033 5 1 1 26032
0 26034 7 2 2 81326 85603
0 26035 5 1 1 93482
0 26036 7 1 2 90717 26035
0 26037 5 1 1 26036
0 26038 7 1 2 64733 26037
0 26039 5 1 1 26038
0 26040 7 2 2 62655 77963
0 26041 5 1 1 93484
0 26042 7 1 2 82370 93485
0 26043 5 1 1 26042
0 26044 7 1 2 26039 26043
0 26045 5 1 1 26044
0 26046 7 1 2 72593 26045
0 26047 5 1 1 26046
0 26048 7 5 2 76183 78702
0 26049 7 1 2 78623 93486
0 26050 5 1 1 26049
0 26051 7 1 2 75578 77319
0 26052 5 1 1 26051
0 26053 7 1 2 90389 26052
0 26054 7 1 2 26050 26053
0 26055 5 1 1 26054
0 26056 7 1 2 77860 26055
0 26057 5 1 1 26056
0 26058 7 1 2 75206 73426
0 26059 5 1 1 26058
0 26060 7 1 2 77359 87614
0 26061 5 1 1 26060
0 26062 7 1 2 75579 78624
0 26063 7 1 2 26061 26062
0 26064 5 1 1 26063
0 26065 7 1 2 26059 26064
0 26066 7 1 2 26057 26065
0 26067 5 1 1 26066
0 26068 7 1 2 66275 26067
0 26069 5 1 1 26068
0 26070 7 1 2 2825 17312
0 26071 5 1 1 26070
0 26072 7 1 2 77320 26071
0 26073 5 1 1 26072
0 26074 7 1 2 5794 91253
0 26075 7 1 2 26073 26074
0 26076 5 1 1 26075
0 26077 7 1 2 83460 26076
0 26078 5 1 1 26077
0 26079 7 1 2 79403 91330
0 26080 5 1 1 26079
0 26081 7 1 2 68348 26080
0 26082 7 1 2 26078 26081
0 26083 7 1 2 26069 26082
0 26084 7 1 2 26047 26083
0 26085 5 1 1 26084
0 26086 7 1 2 65414 26085
0 26087 7 1 2 26033 26086
0 26088 5 1 1 26087
0 26089 7 1 2 64734 79773
0 26090 5 2 1 26089
0 26091 7 1 2 80743 84856
0 26092 5 1 1 26091
0 26093 7 1 2 93491 26092
0 26094 5 1 1 26093
0 26095 7 1 2 69810 26094
0 26096 5 1 1 26095
0 26097 7 1 2 78944 84737
0 26098 5 2 1 26097
0 26099 7 1 2 26096 93493
0 26100 5 1 1 26099
0 26101 7 1 2 77470 26100
0 26102 5 1 1 26101
0 26103 7 1 2 79076 86652
0 26104 5 1 1 26103
0 26105 7 1 2 26102 26104
0 26106 5 1 1 26105
0 26107 7 3 2 77861 77964
0 26108 7 1 2 26106 93495
0 26109 5 1 1 26108
0 26110 7 1 2 68675 26109
0 26111 7 1 2 26088 26110
0 26112 5 1 1 26111
0 26113 7 1 2 66829 26112
0 26114 7 1 2 25950 26113
0 26115 5 1 1 26114
0 26116 7 2 2 75207 83095
0 26117 5 1 1 93498
0 26118 7 2 2 66276 93499
0 26119 5 2 1 93500
0 26120 7 5 2 63009 79560
0 26121 7 1 2 76960 93504
0 26122 5 1 1 26121
0 26123 7 3 2 65713 86032
0 26124 5 1 1 93509
0 26125 7 1 2 64280 93510
0 26126 5 1 1 26125
0 26127 7 1 2 64735 86023
0 26128 5 1 1 26127
0 26129 7 1 2 93085 26128
0 26130 7 1 2 26126 26129
0 26131 5 1 1 26130
0 26132 7 1 2 63447 26131
0 26133 5 1 1 26132
0 26134 7 1 2 26122 26133
0 26135 5 1 1 26134
0 26136 7 1 2 62656 77146
0 26137 7 1 2 26135 26136
0 26138 5 1 1 26137
0 26139 7 1 2 93502 26138
0 26140 5 1 1 26139
0 26141 7 1 2 64974 26140
0 26142 5 1 1 26141
0 26143 7 3 2 80027 78562
0 26144 5 1 1 93512
0 26145 7 1 2 82775 93513
0 26146 7 1 2 93381 26145
0 26147 5 1 1 26146
0 26148 7 1 2 26142 26147
0 26149 5 1 1 26148
0 26150 7 1 2 63741 86061
0 26151 7 1 2 26149 26150
0 26152 5 1 1 26151
0 26153 7 1 2 26115 26152
0 26154 5 1 1 26153
0 26155 7 1 2 66694 26154
0 26156 5 1 1 26155
0 26157 7 1 2 84772 91193
0 26158 5 2 1 26157
0 26159 7 1 2 62309 85134
0 26160 5 1 1 26159
0 26161 7 1 2 93515 26160
0 26162 5 1 1 26161
0 26163 7 1 2 82049 26162
0 26164 5 1 1 26163
0 26165 7 1 2 84410 92955
0 26166 7 1 2 91341 26165
0 26167 5 1 1 26166
0 26168 7 1 2 26164 26167
0 26169 5 1 1 26168
0 26170 7 1 2 79100 26169
0 26171 5 1 1 26170
0 26172 7 2 2 74278 75685
0 26173 7 1 2 77399 85135
0 26174 7 1 2 93517 26173
0 26175 5 1 1 26174
0 26176 7 1 2 26171 26175
0 26177 5 1 1 26176
0 26178 7 1 2 69811 26177
0 26179 5 1 1 26178
0 26180 7 1 2 68349 84121
0 26181 7 1 2 93382 26180
0 26182 5 1 1 26181
0 26183 7 1 2 84751 26182
0 26184 5 1 1 26183
0 26185 7 1 2 63010 26184
0 26186 5 1 1 26185
0 26187 7 1 2 74223 93327
0 26188 5 1 1 26187
0 26189 7 1 2 26186 26188
0 26190 5 1 1 26189
0 26191 7 1 2 65415 26190
0 26192 5 1 1 26191
0 26193 7 3 2 75686 78703
0 26194 5 1 1 93519
0 26195 7 1 2 71031 74849
0 26196 7 1 2 93520 26195
0 26197 5 1 1 26196
0 26198 7 1 2 26192 26197
0 26199 5 1 1 26198
0 26200 7 1 2 66277 26199
0 26201 5 1 1 26200
0 26202 7 3 2 64736 81767
0 26203 7 1 2 84681 93522
0 26204 5 1 1 26203
0 26205 7 1 2 26201 26204
0 26206 5 1 1 26205
0 26207 7 1 2 68676 26206
0 26208 5 1 1 26207
0 26209 7 1 2 26179 26208
0 26210 5 1 1 26209
0 26211 7 1 2 66695 26210
0 26212 5 1 1 26211
0 26213 7 1 2 64737 79204
0 26214 5 2 1 26213
0 26215 7 1 2 85474 93525
0 26216 5 1 1 26215
0 26217 7 1 2 69812 26216
0 26218 5 1 1 26217
0 26219 7 1 2 80510 84588
0 26220 5 1 1 26219
0 26221 7 1 2 26218 26220
0 26222 5 1 1 26221
0 26223 7 1 2 83096 26222
0 26224 5 1 1 26223
0 26225 7 2 2 65416 78757
0 26226 5 2 1 93527
0 26227 7 1 2 62102 93528
0 26228 5 1 1 26227
0 26229 7 1 2 26224 26228
0 26230 5 1 1 26229
0 26231 7 1 2 62657 26230
0 26232 5 1 1 26231
0 26233 7 6 2 64738 65417
0 26234 7 4 2 62310 78758
0 26235 5 2 1 93537
0 26236 7 1 2 93531 93538
0 26237 5 1 1 26236
0 26238 7 1 2 26232 26237
0 26239 5 1 1 26238
0 26240 7 1 2 64975 26239
0 26241 5 1 1 26240
0 26242 7 6 2 65418 69367
0 26243 5 1 1 93543
0 26244 7 1 2 87459 93539
0 26245 7 1 2 93544 26244
0 26246 5 1 1 26245
0 26247 7 1 2 26241 26246
0 26248 5 1 1 26247
0 26249 7 1 2 81358 26248
0 26250 5 1 1 26249
0 26251 7 1 2 26212 26250
0 26252 5 1 1 26251
0 26253 7 1 2 64510 26252
0 26254 5 1 1 26253
0 26255 7 1 2 80564 84738
0 26256 5 1 1 26255
0 26257 7 1 2 90618 90687
0 26258 5 1 1 26257
0 26259 7 1 2 69813 93366
0 26260 7 1 2 26258 26259
0 26261 5 1 1 26260
0 26262 7 1 2 26256 26261
0 26263 5 1 1 26262
0 26264 7 1 2 84479 26263
0 26265 5 1 1 26264
0 26266 7 1 2 79121 88039
0 26267 5 1 1 26266
0 26268 7 1 2 12164 26267
0 26269 5 1 1 26268
0 26270 7 1 2 66026 26269
0 26271 5 1 1 26270
0 26272 7 1 2 4718 26271
0 26273 5 1 1 26272
0 26274 7 1 2 65419 26273
0 26275 5 1 1 26274
0 26276 7 1 2 88195 93496
0 26277 5 1 1 26276
0 26278 7 1 2 26275 26277
0 26279 5 1 1 26278
0 26280 7 1 2 89928 26279
0 26281 5 1 1 26280
0 26282 7 1 2 26265 26281
0 26283 5 1 1 26282
0 26284 7 1 2 73871 26283
0 26285 5 1 1 26284
0 26286 7 1 2 80900 77862
0 26287 7 1 2 81741 26286
0 26288 5 1 1 26287
0 26289 7 1 2 79648 26288
0 26290 5 1 1 26289
0 26291 7 1 2 83649 26290
0 26292 5 1 1 26291
0 26293 7 1 2 71032 85215
0 26294 5 1 1 26293
0 26295 7 1 2 26292 26294
0 26296 5 1 1 26295
0 26297 7 1 2 76233 26296
0 26298 5 1 1 26297
0 26299 7 2 2 66696 70974
0 26300 5 1 1 93549
0 26301 7 1 2 61076 26300
0 26302 5 1 1 26301
0 26303 7 1 2 61720 79474
0 26304 5 2 1 26303
0 26305 7 1 2 84773 93532
0 26306 7 1 2 93551 26305
0 26307 7 1 2 26302 26306
0 26308 5 1 1 26307
0 26309 7 1 2 26298 26308
0 26310 5 1 1 26309
0 26311 7 1 2 84181 79571
0 26312 7 1 2 82744 26311
0 26313 5 1 1 26312
0 26314 7 1 2 8960 26313
0 26315 5 1 1 26314
0 26316 7 1 2 64511 26315
0 26317 5 1 1 26316
0 26318 7 2 2 60535 69814
0 26319 7 1 2 85317 93553
0 26320 5 1 1 26319
0 26321 7 1 2 26317 26320
0 26322 5 1 1 26321
0 26323 7 1 2 87879 26322
0 26324 5 1 1 26323
0 26325 7 1 2 85136 89443
0 26326 5 1 1 26325
0 26327 7 1 2 63448 26326
0 26328 7 1 2 26324 26327
0 26329 5 1 1 26328
0 26330 7 2 2 62103 26329
0 26331 7 1 2 26310 93555
0 26332 5 1 1 26331
0 26333 7 1 2 69815 75068
0 26334 5 1 1 26333
0 26335 7 1 2 90619 26334
0 26336 5 1 1 26335
0 26337 7 1 2 65205 90605
0 26338 5 2 1 26337
0 26339 7 1 2 93215 93557
0 26340 5 1 1 26339
0 26341 7 1 2 88223 26340
0 26342 7 1 2 26336 26341
0 26343 5 1 1 26342
0 26344 7 1 2 26332 26343
0 26345 7 1 2 26285 26344
0 26346 5 1 1 26345
0 26347 7 1 2 63011 26346
0 26348 5 1 1 26347
0 26349 7 1 2 64512 81313
0 26350 7 1 2 88220 26349
0 26351 5 1 1 26350
0 26352 7 1 2 68350 26351
0 26353 5 1 1 26352
0 26354 7 1 2 93556 26353
0 26355 5 1 1 26354
0 26356 7 1 2 61342 77325
0 26357 7 1 2 88042 26356
0 26358 5 1 1 26357
0 26359 7 1 2 75069 26358
0 26360 5 1 1 26359
0 26361 7 1 2 6512 26360
0 26362 5 1 1 26361
0 26363 7 1 2 85323 26362
0 26364 5 1 1 26363
0 26365 7 1 2 26355 26364
0 26366 7 1 2 26348 26365
0 26367 5 1 1 26366
0 26368 7 1 2 66507 26367
0 26369 5 1 1 26368
0 26370 7 1 2 76184 87801
0 26371 5 1 1 26370
0 26372 7 3 2 64976 81950
0 26373 5 1 1 93559
0 26374 7 1 2 84081 93405
0 26375 7 1 2 93560 26374
0 26376 5 1 1 26375
0 26377 7 1 2 26371 26376
0 26378 5 1 1 26377
0 26379 7 1 2 85205 26378
0 26380 5 1 1 26379
0 26381 7 2 2 65420 80731
0 26382 5 2 1 93562
0 26383 7 1 2 25554 93564
0 26384 5 1 1 26383
0 26385 7 1 2 85199 26384
0 26386 5 1 1 26385
0 26387 7 1 2 26380 26386
0 26388 5 1 1 26387
0 26389 7 1 2 66027 26388
0 26390 5 1 1 26389
0 26391 7 1 2 69816 70488
0 26392 7 1 2 80511 26391
0 26393 7 1 2 89748 26392
0 26394 5 1 1 26393
0 26395 7 1 2 26390 26394
0 26396 5 1 1 26395
0 26397 7 1 2 65206 26396
0 26398 5 1 1 26397
0 26399 7 3 2 80658 90720
0 26400 5 1 1 93566
0 26401 7 1 2 70489 93567
0 26402 5 1 1 26401
0 26403 7 1 2 93492 26402
0 26404 5 1 1 26403
0 26405 7 1 2 79614 83650
0 26406 7 1 2 26404 26405
0 26407 5 1 1 26406
0 26408 7 1 2 26398 26407
0 26409 5 1 1 26408
0 26410 7 1 2 63012 26409
0 26411 5 1 1 26410
0 26412 7 2 2 82174 84343
0 26413 5 1 1 93569
0 26414 7 1 2 76844 88227
0 26415 7 1 2 92422 26414
0 26416 5 1 1 26415
0 26417 7 1 2 26413 26416
0 26418 5 1 1 26417
0 26419 7 1 2 91331 26418
0 26420 5 1 1 26419
0 26421 7 2 2 77904 74482
0 26422 5 1 1 93571
0 26423 7 2 2 69817 78563
0 26424 5 1 1 93573
0 26425 7 1 2 68351 93574
0 26426 5 1 1 26425
0 26427 7 1 2 26422 26426
0 26428 5 1 1 26427
0 26429 7 1 2 73103 26428
0 26430 5 1 1 26429
0 26431 7 1 2 62658 93235
0 26432 5 1 1 26431
0 26433 7 1 2 26430 26432
0 26434 5 1 1 26433
0 26435 7 1 2 85324 26434
0 26436 5 1 1 26435
0 26437 7 1 2 26420 26436
0 26438 5 1 1 26437
0 26439 7 1 2 77192 26438
0 26440 5 1 1 26439
0 26441 7 4 2 61721 88231
0 26442 5 2 1 93575
0 26443 7 1 2 82676 93576
0 26444 5 1 1 26443
0 26445 7 4 2 61722 83633
0 26446 5 4 1 93581
0 26447 7 1 2 64739 84344
0 26448 5 2 1 26447
0 26449 7 1 2 93585 93589
0 26450 5 1 1 26449
0 26451 7 1 2 90856 26450
0 26452 5 1 1 26451
0 26453 7 1 2 26444 26452
0 26454 5 1 1 26453
0 26455 7 4 2 65421 70799
0 26456 5 3 1 93591
0 26457 7 1 2 90738 93592
0 26458 7 1 2 26454 26457
0 26459 5 1 1 26458
0 26460 7 1 2 26440 26459
0 26461 7 1 2 26411 26460
0 26462 7 1 2 26369 26461
0 26463 7 1 2 26254 26462
0 26464 5 1 1 26463
0 26465 7 1 2 65860 26464
0 26466 5 1 1 26465
0 26467 7 1 2 82776 93220
0 26468 5 1 1 26467
0 26469 7 1 2 60536 87657
0 26470 5 1 1 26469
0 26471 7 1 2 26468 26470
0 26472 5 1 1 26471
0 26473 7 1 2 63013 26472
0 26474 5 1 1 26473
0 26475 7 1 2 60155 148
0 26476 5 1 1 26475
0 26477 7 1 2 60537 26476
0 26478 5 1 1 26477
0 26479 7 2 2 66028 89394
0 26480 5 2 1 93598
0 26481 7 1 2 62104 90629
0 26482 5 1 1 26481
0 26483 7 1 2 93600 26482
0 26484 5 1 1 26483
0 26485 7 1 2 64740 26484
0 26486 5 1 1 26485
0 26487 7 1 2 26478 26486
0 26488 5 1 1 26487
0 26489 7 1 2 92943 26488
0 26490 5 1 1 26489
0 26491 7 1 2 26474 26490
0 26492 5 1 1 26491
0 26493 7 1 2 63449 26492
0 26494 5 1 1 26493
0 26495 7 2 2 66508 83866
0 26496 5 1 1 93602
0 26497 7 1 2 60538 26496
0 26498 5 1 1 26497
0 26499 7 1 2 77350 26498
0 26500 5 1 1 26499
0 26501 7 1 2 62105 93533
0 26502 5 1 1 26501
0 26503 7 1 2 11484 26502
0 26504 5 1 1 26503
0 26505 7 1 2 64513 26504
0 26506 5 1 1 26505
0 26507 7 1 2 77250 93545
0 26508 5 1 1 26507
0 26509 7 1 2 26506 26508
0 26510 5 1 1 26509
0 26511 7 1 2 62311 26510
0 26512 5 1 1 26511
0 26513 7 1 2 26500 26512
0 26514 5 1 1 26513
0 26515 7 1 2 90739 26514
0 26516 5 1 1 26515
0 26517 7 1 2 26494 26516
0 26518 5 1 1 26517
0 26519 7 1 2 66278 26518
0 26520 5 1 1 26519
0 26521 7 1 2 73872 90578
0 26522 5 1 1 26521
0 26523 7 2 2 65422 81537
0 26524 5 1 1 93604
0 26525 7 1 2 66029 93605
0 26526 5 1 1 26525
0 26527 7 1 2 26522 26526
0 26528 5 1 1 26527
0 26529 7 1 2 69818 26528
0 26530 5 1 1 26529
0 26531 7 1 2 64977 90579
0 26532 5 1 1 26531
0 26533 7 1 2 82175 90894
0 26534 5 1 1 26533
0 26535 7 1 2 26532 26534
0 26536 7 1 2 26530 26535
0 26537 5 1 1 26536
0 26538 7 1 2 63014 26537
0 26539 5 1 1 26538
0 26540 7 2 2 64741 79147
0 26541 5 1 1 93606
0 26542 7 1 2 77863 82176
0 26543 7 1 2 93607 26542
0 26544 5 1 1 26543
0 26545 7 1 2 26539 26544
0 26546 5 1 1 26545
0 26547 7 1 2 62312 26546
0 26548 5 1 1 26547
0 26549 7 3 2 68352 87444
0 26550 7 1 2 73226 93608
0 26551 5 1 1 26550
0 26552 7 1 2 79077 70534
0 26553 7 1 2 77905 26552
0 26554 5 1 1 26553
0 26555 7 1 2 26551 26554
0 26556 5 1 1 26555
0 26557 7 1 2 93207 26556
0 26558 5 1 1 26557
0 26559 7 1 2 26548 26558
0 26560 5 1 1 26559
0 26561 7 1 2 65207 26560
0 26562 5 1 1 26561
0 26563 7 1 2 26520 26562
0 26564 5 1 1 26563
0 26565 7 1 2 63742 26564
0 26566 5 1 1 26565
0 26567 7 2 2 71273 87842
0 26568 7 1 2 84074 89684
0 26569 7 1 2 93611 26568
0 26570 5 1 1 26569
0 26571 7 1 2 26566 26570
0 26572 5 1 1 26571
0 26573 7 1 2 61723 26572
0 26574 5 1 1 26573
0 26575 7 1 2 25427 93412
0 26576 5 1 1 26575
0 26577 7 1 2 73104 26576
0 26578 5 1 1 26577
0 26579 7 1 2 77606 91169
0 26580 5 1 1 26579
0 26581 7 1 2 26578 26580
0 26582 5 1 1 26581
0 26583 7 1 2 69819 26582
0 26584 5 1 1 26583
0 26585 7 2 2 64514 77986
0 26586 5 1 1 93613
0 26587 7 1 2 85943 93614
0 26588 5 1 1 26587
0 26589 7 1 2 26584 26588
0 26590 5 1 1 26589
0 26591 7 1 2 62106 26590
0 26592 5 1 1 26591
0 26593 7 1 2 82149 85395
0 26594 5 1 1 26593
0 26595 7 1 2 26592 26594
0 26596 5 1 1 26595
0 26597 7 2 2 64978 81314
0 26598 7 1 2 83623 93615
0 26599 7 1 2 26596 26598
0 26600 5 1 1 26599
0 26601 7 1 2 26574 26600
0 26602 7 1 2 26466 26601
0 26603 5 1 1 26602
0 26604 7 1 2 66830 26603
0 26605 5 1 1 26604
0 26606 7 1 2 64742 93362
0 26607 5 1 1 26606
0 26608 7 1 2 81647 26607
0 26609 5 1 1 26608
0 26610 7 1 2 66509 26609
0 26611 5 1 1 26610
0 26612 7 1 2 81953 26611
0 26613 5 1 1 26612
0 26614 7 1 2 63015 26613
0 26615 5 1 1 26614
0 26616 7 1 2 80028 75040
0 26617 5 1 1 26616
0 26618 7 1 2 26615 26617
0 26619 5 1 1 26618
0 26620 7 1 2 65208 26619
0 26621 5 1 1 26620
0 26622 7 1 2 26144 26621
0 26623 5 1 1 26622
0 26624 7 1 2 93216 93503
0 26625 5 1 1 26624
0 26626 7 3 2 79615 79708
0 26627 7 1 2 65861 93617
0 26628 7 1 2 26625 26627
0 26629 7 1 2 26623 26628
0 26630 5 1 1 26629
0 26631 7 1 2 26605 26630
0 26632 7 1 2 26156 26631
0 26633 5 1 1 26632
0 26634 7 1 2 63971 26633
0 26635 5 1 1 26634
0 26636 7 1 2 66510 89090
0 26637 5 2 1 26636
0 26638 7 1 2 66279 86832
0 26639 7 1 2 93126 26638
0 26640 5 1 1 26639
0 26641 7 1 2 93620 26640
0 26642 5 1 1 26641
0 26643 7 1 2 64743 26642
0 26644 5 1 1 26643
0 26645 7 1 2 81648 85821
0 26646 5 1 1 26645
0 26647 7 1 2 75208 26646
0 26648 5 1 1 26647
0 26649 7 3 2 75906 76845
0 26650 7 1 2 86833 87407
0 26651 7 1 2 93622 26650
0 26652 5 1 1 26651
0 26653 7 1 2 26648 26652
0 26654 7 1 2 26644 26653
0 26655 5 1 1 26654
0 26656 7 1 2 63450 26655
0 26657 5 1 1 26656
0 26658 7 1 2 83201 82814
0 26659 7 1 2 80598 26658
0 26660 7 1 2 76234 85385
0 26661 7 1 2 26659 26660
0 26662 5 1 1 26661
0 26663 7 1 2 26657 26662
0 26664 5 1 1 26663
0 26665 7 1 2 93208 26664
0 26666 5 1 1 26665
0 26667 7 1 2 93194 93501
0 26668 5 1 1 26667
0 26669 7 1 2 26666 26668
0 26670 5 1 1 26669
0 26671 7 9 2 66831 85514
0 26672 7 1 2 79616 93625
0 26673 7 1 2 26670 26672
0 26674 5 1 1 26673
0 26675 7 1 2 26635 26674
0 26676 5 1 1 26675
0 26677 7 1 2 60660 26676
0 26678 5 1 1 26677
0 26679 7 1 2 68353 77965
0 26680 7 1 2 88012 26679
0 26681 5 1 1 26680
0 26682 7 2 2 62659 90606
0 26683 5 1 1 93634
0 26684 7 1 2 26681 26683
0 26685 5 1 1 26684
0 26686 7 1 2 78058 26685
0 26687 5 1 1 26686
0 26688 7 1 2 76210 83097
0 26689 7 1 2 80689 26688
0 26690 7 1 2 82216 26689
0 26691 5 1 1 26690
0 26692 7 1 2 26687 26691
0 26693 5 1 1 26692
0 26694 7 1 2 61546 26693
0 26695 5 1 1 26694
0 26696 7 1 2 81754 78923
0 26697 5 1 1 26696
0 26698 7 2 2 74483 87260
0 26699 7 5 2 64281 65423
0 26700 5 1 1 93638
0 26701 7 2 2 65714 93639
0 26702 7 1 2 86338 93643
0 26703 7 1 2 93636 26702
0 26704 5 1 1 26703
0 26705 7 1 2 26697 26704
0 26706 5 1 1 26705
0 26707 7 1 2 75664 26706
0 26708 5 1 1 26707
0 26709 7 1 2 63451 87915
0 26710 7 1 2 86636 26709
0 26711 5 1 1 26710
0 26712 7 1 2 26708 26711
0 26713 7 1 2 26695 26712
0 26714 5 1 1 26713
0 26715 7 1 2 66832 26714
0 26716 5 1 1 26715
0 26717 7 2 2 72768 82344
0 26718 5 2 1 93645
0 26719 7 1 2 87685 93647
0 26720 5 1 1 26719
0 26721 7 1 2 66697 26720
0 26722 5 1 1 26721
0 26723 7 1 2 66511 93646
0 26724 5 1 1 26723
0 26725 7 1 2 62660 79438
0 26726 5 1 1 26725
0 26727 7 1 2 26724 26726
0 26728 5 1 1 26727
0 26729 7 1 2 65209 26728
0 26730 5 1 1 26729
0 26731 7 1 2 26722 26730
0 26732 5 1 1 26731
0 26733 7 1 2 65424 26732
0 26734 5 1 1 26733
0 26735 7 1 2 75209 86339
0 26736 7 1 2 93572 26735
0 26737 5 1 1 26736
0 26738 7 1 2 26734 26737
0 26739 5 1 1 26738
0 26740 7 1 2 69820 26739
0 26741 5 1 1 26740
0 26742 7 3 2 65862 75665
0 26743 5 1 1 93649
0 26744 7 1 2 79809 26743
0 26745 5 1 1 26744
0 26746 7 1 2 62661 79617
0 26747 7 1 2 26745 26746
0 26748 5 1 1 26747
0 26749 7 1 2 26741 26748
0 26750 5 1 1 26749
0 26751 7 1 2 86079 26750
0 26752 5 1 1 26751
0 26753 7 1 2 26716 26752
0 26754 5 1 1 26753
0 26755 7 1 2 68677 26754
0 26756 5 1 1 26755
0 26757 7 1 2 75141 85843
0 26758 7 1 2 88147 26757
0 26759 5 1 1 26758
0 26760 7 4 2 61547 86970
0 26761 5 1 1 93652
0 26762 7 1 2 85863 26761
0 26763 5 1 1 26762
0 26764 7 1 2 65210 26763
0 26765 5 1 1 26764
0 26766 7 1 2 66512 87103
0 26767 5 1 1 26766
0 26768 7 1 2 26765 26767
0 26769 5 2 1 26768
0 26770 7 1 2 73168 89243
0 26771 7 1 2 93656 26770
0 26772 5 1 1 26771
0 26773 7 1 2 26759 26772
0 26774 5 1 1 26773
0 26775 7 1 2 72551 26774
0 26776 5 1 1 26775
0 26777 7 4 2 66513 90697
0 26778 5 1 1 93658
0 26779 7 3 2 66833 81987
0 26780 5 1 1 93662
0 26781 7 1 2 87091 26780
0 26782 5 1 1 26781
0 26783 7 1 2 82108 88078
0 26784 7 1 2 26782 26783
0 26785 7 1 2 93659 26784
0 26786 5 1 1 26785
0 26787 7 1 2 26776 26786
0 26788 5 1 1 26787
0 26789 7 1 2 83634 26788
0 26790 5 1 1 26789
0 26791 7 1 2 26756 26790
0 26792 5 1 1 26791
0 26793 7 1 2 64744 26792
0 26794 5 1 1 26793
0 26795 7 2 2 68872 87104
0 26796 7 1 2 89109 93665
0 26797 5 1 1 26796
0 26798 7 2 2 66280 72552
0 26799 7 3 2 61863 81019
0 26800 5 1 1 93669
0 26801 7 1 2 86538 93670
0 26802 7 1 2 93667 26801
0 26803 5 1 1 26802
0 26804 7 1 2 26797 26803
0 26805 5 1 1 26804
0 26806 7 1 2 66514 26805
0 26807 5 1 1 26806
0 26808 7 4 2 61724 86080
0 26809 5 1 1 93672
0 26810 7 1 2 93233 93673
0 26811 5 1 1 26810
0 26812 7 1 2 26807 26811
0 26813 5 1 1 26812
0 26814 7 1 2 65211 26813
0 26815 5 1 1 26814
0 26816 7 2 2 86209 87312
0 26817 7 1 2 81085 93676
0 26818 5 1 1 26817
0 26819 7 1 2 26815 26818
0 26820 5 1 1 26819
0 26821 7 1 2 85187 26820
0 26822 5 1 1 26821
0 26823 7 1 2 26794 26822
0 26824 5 1 1 26823
0 26825 7 1 2 66030 26824
0 26826 5 1 1 26825
0 26827 7 1 2 81063 86495
0 26828 7 1 2 87105 26827
0 26829 5 1 1 26828
0 26830 7 1 2 26826 26829
0 26831 5 1 1 26830
0 26832 7 1 2 64979 26831
0 26833 5 1 1 26832
0 26834 7 1 2 81057 10278
0 26835 5 2 1 26834
0 26836 7 1 2 65212 93678
0 26837 5 1 1 26836
0 26838 7 1 2 62107 93102
0 26839 5 1 1 26838
0 26840 7 1 2 89538 26839
0 26841 5 1 1 26840
0 26842 7 1 2 76825 26841
0 26843 5 2 1 26842
0 26844 7 1 2 26837 93680
0 26845 5 1 1 26844
0 26846 7 1 2 63972 87106
0 26847 7 1 2 26845 26846
0 26848 5 1 1 26847
0 26849 7 1 2 75142 86562
0 26850 5 1 1 26849
0 26851 7 1 2 65863 77400
0 26852 5 2 1 26851
0 26853 7 1 2 86892 93682
0 26854 5 1 1 26853
0 26855 7 1 2 69821 26854
0 26856 5 1 1 26855
0 26857 7 1 2 64745 77401
0 26858 5 1 1 26857
0 26859 7 1 2 65864 86889
0 26860 5 1 1 26859
0 26861 7 2 2 26858 26860
0 26862 5 1 1 93684
0 26863 7 1 2 26856 93685
0 26864 5 1 1 26863
0 26865 7 1 2 79526 26864
0 26866 5 1 1 26865
0 26867 7 1 2 26850 26866
0 26868 5 1 1 26867
0 26869 7 1 2 79747 87540
0 26870 7 1 2 26868 26869
0 26871 5 1 1 26870
0 26872 7 1 2 26848 26871
0 26873 5 1 1 26872
0 26874 7 1 2 68678 26873
0 26875 5 1 1 26874
0 26876 7 3 2 75921 86081
0 26877 5 1 1 93686
0 26878 7 1 2 80867 93687
0 26879 5 1 1 26878
0 26880 7 1 2 72553 76846
0 26881 7 1 2 93666 26880
0 26882 5 1 1 26881
0 26883 7 1 2 26879 26882
0 26884 5 1 1 26883
0 26885 7 1 2 64746 26884
0 26886 5 1 1 26885
0 26887 7 1 2 81755 86501
0 26888 5 1 1 26887
0 26889 7 1 2 26886 26888
0 26890 5 1 1 26889
0 26891 7 1 2 79101 26890
0 26892 5 1 1 26891
0 26893 7 3 2 60539 73478
0 26894 7 1 2 86340 86351
0 26895 7 1 2 93689 26894
0 26896 5 1 1 26895
0 26897 7 1 2 26892 26896
0 26898 5 1 1 26897
0 26899 7 1 2 86382 26898
0 26900 5 1 1 26899
0 26901 7 1 2 26875 26900
0 26902 5 1 1 26901
0 26903 7 1 2 63452 26902
0 26904 5 1 1 26903
0 26905 7 2 2 74484 87275
0 26906 5 2 1 93692
0 26907 7 4 2 66281 86155
0 26908 5 2 1 93696
0 26909 7 1 2 60357 93697
0 26910 5 1 1 26909
0 26911 7 1 2 93694 26910
0 26912 5 1 1 26911
0 26913 7 1 2 69822 26912
0 26914 5 1 1 26913
0 26915 7 2 2 87261 87592
0 26916 5 1 1 93702
0 26917 7 1 2 93695 26916
0 26918 5 1 1 26917
0 26919 7 1 2 65865 26918
0 26920 5 1 1 26919
0 26921 7 1 2 26914 26920
0 26922 5 1 1 26921
0 26923 7 1 2 79205 26922
0 26924 5 1 1 26923
0 26925 7 3 2 66282 86082
0 26926 5 2 1 93704
0 26927 7 2 2 66834 76826
0 26928 7 1 2 93637 93709
0 26929 5 1 1 26928
0 26930 7 1 2 93707 26929
0 26931 5 1 1 26930
0 26932 7 1 2 83624 26931
0 26933 5 1 1 26932
0 26934 7 1 2 26924 26933
0 26935 5 1 1 26934
0 26936 7 1 2 79618 26935
0 26937 5 1 1 26936
0 26938 7 1 2 75210 83651
0 26939 5 2 1 26938
0 26940 7 1 2 82611 78968
0 26941 7 1 2 84002 26940
0 26942 5 1 1 26941
0 26943 7 1 2 93711 26942
0 26944 5 1 1 26943
0 26945 7 1 2 78059 87205
0 26946 7 1 2 26944 26945
0 26947 5 1 1 26946
0 26948 7 1 2 26937 26947
0 26949 5 1 1 26948
0 26950 7 1 2 68354 26949
0 26951 5 1 1 26950
0 26952 7 1 2 65564 26951
0 26953 7 1 2 26904 26952
0 26954 7 1 2 26833 26953
0 26955 5 1 1 26954
0 26956 7 1 2 89110 92946
0 26957 5 1 1 26956
0 26958 7 4 2 63453 75580
0 26959 5 3 1 93713
0 26960 7 1 2 72554 93714
0 26961 5 1 1 26960
0 26962 7 1 2 75211 75922
0 26963 5 1 1 26962
0 26964 7 1 2 26961 26963
0 26965 5 1 1 26964
0 26966 7 1 2 93209 26965
0 26967 5 1 1 26966
0 26968 7 1 2 75212 81406
0 26969 5 1 1 26968
0 26970 7 1 2 26967 26969
0 26971 5 1 1 26970
0 26972 7 1 2 83867 76847
0 26973 7 1 2 26971 26972
0 26974 5 1 1 26973
0 26975 7 1 2 26957 26974
0 26976 5 1 1 26975
0 26977 7 1 2 87934 26976
0 26978 5 1 1 26977
0 26979 7 1 2 71111 93679
0 26980 5 1 1 26979
0 26981 7 1 2 81068 26980
0 26982 5 1 1 26981
0 26983 7 1 2 64980 26982
0 26984 5 1 1 26983
0 26985 7 1 2 93681 26984
0 26986 5 1 1 26985
0 26987 7 1 2 84182 26986
0 26988 5 1 1 26987
0 26989 7 3 2 84430 91758
0 26990 7 1 2 86686 93720
0 26991 5 1 1 26990
0 26992 7 1 2 26988 26991
0 26993 5 1 1 26992
0 26994 7 1 2 66698 26993
0 26995 5 1 1 26994
0 26996 7 1 2 79387 86449
0 26997 7 1 2 92032 26996
0 26998 5 1 1 26997
0 26999 7 1 2 26995 26998
0 27000 5 1 1 26999
0 27001 7 1 2 63454 27000
0 27002 5 1 1 27001
0 27003 7 1 2 79619 77607
0 27004 5 1 1 27003
0 27005 7 2 2 80901 86653
0 27006 7 1 2 72769 91091
0 27007 7 1 2 93723 27006
0 27008 5 1 1 27007
0 27009 7 1 2 27004 27008
0 27010 5 1 1 27009
0 27011 7 1 2 68679 27010
0 27012 5 1 1 27011
0 27013 7 1 2 86848 93356
0 27014 5 1 1 27013
0 27015 7 1 2 77608 93210
0 27016 5 1 1 27015
0 27017 7 1 2 27014 27016
0 27018 5 1 1 27017
0 27019 7 1 2 69823 27018
0 27020 5 1 1 27019
0 27021 7 1 2 88330 90721
0 27022 5 1 1 27021
0 27023 7 1 2 90620 27022
0 27024 5 1 1 27023
0 27025 7 1 2 66283 27024
0 27026 5 1 1 27025
0 27027 7 1 2 27020 27026
0 27028 5 1 1 27027
0 27029 7 1 2 85785 27028
0 27030 5 1 1 27029
0 27031 7 1 2 27012 27030
0 27032 5 1 1 27031
0 27033 7 1 2 66515 27032
0 27034 5 1 1 27033
0 27035 7 1 2 16712 93648
0 27036 5 1 1 27035
0 27037 7 1 2 69824 27036
0 27038 5 1 1 27037
0 27039 7 1 2 68355 78512
0 27040 7 1 2 77077 27039
0 27041 5 1 1 27040
0 27042 7 1 2 79810 27041
0 27043 5 1 1 27042
0 27044 7 1 2 62662 27043
0 27045 5 1 1 27044
0 27046 7 1 2 27038 27045
0 27047 5 1 1 27046
0 27048 7 1 2 84183 27047
0 27049 5 1 1 27048
0 27050 7 1 2 80953 78969
0 27051 7 1 2 85155 27050
0 27052 7 1 2 84003 27051
0 27053 5 1 1 27052
0 27054 7 1 2 27049 27053
0 27055 5 1 1 27054
0 27056 7 1 2 66699 27055
0 27057 5 1 1 27056
0 27058 7 1 2 25557 27057
0 27059 7 1 2 27034 27058
0 27060 5 1 1 27059
0 27061 7 1 2 65213 27060
0 27062 5 1 1 27061
0 27063 7 1 2 84774 85274
0 27064 5 1 1 27063
0 27065 7 5 2 68001 82612
0 27066 7 1 2 83635 93725
0 27067 5 1 1 27066
0 27068 7 1 2 27064 27067
0 27069 5 1 1 27068
0 27070 7 1 2 72555 87802
0 27071 7 1 2 27069 27070
0 27072 5 1 1 27071
0 27073 7 1 2 27062 27072
0 27074 7 1 2 27002 27073
0 27075 5 1 1 27074
0 27076 7 1 2 63973 27075
0 27077 5 1 1 27076
0 27078 7 1 2 26978 27077
0 27079 5 1 1 27078
0 27080 7 1 2 66835 27079
0 27081 5 1 1 27080
0 27082 7 3 2 63455 75213
0 27083 5 2 1 93730
0 27084 7 1 2 72516 93717
0 27085 5 1 1 27084
0 27086 7 4 2 75314 93718
0 27087 5 1 1 93735
0 27088 7 1 2 93211 27087
0 27089 7 1 2 27085 27088
0 27090 5 1 1 27089
0 27091 7 1 2 93733 27090
0 27092 5 1 1 27091
0 27093 7 5 2 63974 85844
0 27094 7 1 2 80512 79376
0 27095 7 1 2 93739 27094
0 27096 7 1 2 27092 27095
0 27097 5 1 1 27096
0 27098 7 1 2 60661 27097
0 27099 7 1 2 27081 27098
0 27100 5 1 1 27099
0 27101 7 1 2 26955 27100
0 27102 5 1 1 27101
0 27103 7 1 2 93526 93712
0 27104 5 1 1 27103
0 27105 7 1 2 76827 27104
0 27106 5 1 1 27105
0 27107 7 2 2 66284 79206
0 27108 5 1 1 93744
0 27109 7 1 2 27106 27108
0 27110 5 1 1 27109
0 27111 7 1 2 63016 27110
0 27112 5 1 1 27111
0 27113 7 1 2 84045 85169
0 27114 5 1 1 27113
0 27115 7 1 2 27112 27114
0 27116 5 1 1 27115
0 27117 7 1 2 63456 27116
0 27118 5 1 1 27117
0 27119 7 1 2 78564 93398
0 27120 5 1 1 27119
0 27121 7 1 2 86046 27120
0 27122 5 1 1 27121
0 27123 7 2 2 72556 27122
0 27124 7 1 2 78759 93746
0 27125 5 1 1 27124
0 27126 7 1 2 27118 27125
0 27127 5 1 1 27126
0 27128 7 1 2 87139 27127
0 27129 5 1 1 27128
0 27130 7 1 2 86202 93668
0 27131 5 1 1 27130
0 27132 7 1 2 26877 27131
0 27133 5 1 1 27132
0 27134 7 1 2 64747 27133
0 27135 5 1 1 27134
0 27136 7 2 2 86156 93383
0 27137 5 1 1 93748
0 27138 7 1 2 93708 27137
0 27139 7 1 2 27135 27138
0 27140 5 1 1 27139
0 27141 7 1 2 63017 27140
0 27142 5 1 1 27141
0 27143 7 1 2 66285 93749
0 27144 5 1 1 27143
0 27145 7 1 2 27142 27144
0 27146 5 1 1 27145
0 27147 7 1 2 79207 27146
0 27148 5 1 1 27147
0 27149 7 1 2 78565 93688
0 27150 5 1 1 27149
0 27151 7 1 2 77690 86083
0 27152 5 1 1 27151
0 27153 7 1 2 71112 87268
0 27154 5 1 1 27153
0 27155 7 1 2 27152 27154
0 27156 5 1 1 27155
0 27157 7 1 2 77351 27156
0 27158 5 1 1 27157
0 27159 7 1 2 27150 27158
0 27160 5 1 1 27159
0 27161 7 1 2 83625 27160
0 27162 5 1 1 27161
0 27163 7 1 2 63457 27162
0 27164 7 1 2 27148 27163
0 27165 5 1 1 27164
0 27166 7 1 2 75496 93217
0 27167 5 2 1 27166
0 27168 7 5 2 65715 76848
0 27169 7 1 2 77251 93752
0 27170 7 1 2 93750 27169
0 27171 5 1 1 27170
0 27172 7 1 2 93437 27171
0 27173 5 1 1 27172
0 27174 7 1 2 85817 27173
0 27175 5 1 1 27174
0 27176 7 1 2 69825 81327
0 27177 7 1 2 90384 27176
0 27178 5 1 1 27177
0 27179 7 1 2 27175 27178
0 27180 5 1 1 27179
0 27181 7 1 2 85515 27180
0 27182 5 1 1 27181
0 27183 7 1 2 61343 82144
0 27184 5 2 1 27183
0 27185 7 4 2 68002 77560
0 27186 7 1 2 61548 91574
0 27187 7 1 2 93759 27186
0 27188 7 1 2 93757 27187
0 27189 5 1 1 27188
0 27190 7 1 2 27182 27189
0 27191 5 1 1 27190
0 27192 7 1 2 66836 27191
0 27193 5 1 1 27192
0 27194 7 1 2 86370 93747
0 27195 5 1 1 27194
0 27196 7 1 2 68356 27195
0 27197 7 1 2 27193 27196
0 27198 5 1 1 27197
0 27199 7 1 2 65565 27198
0 27200 7 1 2 27165 27199
0 27201 5 1 1 27200
0 27202 7 1 2 27129 27201
0 27203 5 1 1 27202
0 27204 7 1 2 81179 27203
0 27205 5 1 1 27204
0 27206 7 1 2 27102 27205
0 27207 5 1 1 27206
0 27208 7 1 2 74019 27207
0 27209 5 1 1 27208
0 27210 7 1 2 60540 85284
0 27211 5 2 1 27210
0 27212 7 5 2 68357 80168
0 27213 7 1 2 82449 93765
0 27214 5 1 1 27213
0 27215 7 1 2 76388 84280
0 27216 5 1 1 27215
0 27217 7 1 2 74741 27216
0 27218 5 1 1 27217
0 27219 7 1 2 63458 88228
0 27220 7 1 2 27218 27219
0 27221 5 1 1 27220
0 27222 7 1 2 27214 27221
0 27223 5 1 1 27222
0 27224 7 1 2 63743 27223
0 27225 5 1 1 27224
0 27226 7 7 2 66700 83539
0 27227 7 1 2 74452 74736
0 27228 7 1 2 93770 27227
0 27229 5 1 1 27228
0 27230 7 1 2 27225 27229
0 27231 5 1 1 27230
0 27232 7 1 2 68003 27231
0 27233 5 1 1 27232
0 27234 7 1 2 85750 86413
0 27235 5 1 1 27234
0 27236 7 1 2 64515 87682
0 27237 5 1 1 27236
0 27238 7 1 2 27235 27237
0 27239 5 1 1 27238
0 27240 7 3 2 81909 79013
0 27241 7 1 2 27239 93777
0 27242 5 1 1 27241
0 27243 7 1 2 76849 89685
0 27244 5 1 1 27243
0 27245 7 1 2 85402 27244
0 27246 5 1 1 27245
0 27247 7 1 2 79072 27246
0 27248 5 1 1 27247
0 27249 7 1 2 81553 83981
0 27250 5 1 1 27249
0 27251 7 1 2 27248 27250
0 27252 5 1 1 27251
0 27253 7 1 2 66701 27252
0 27254 5 1 1 27253
0 27255 7 1 2 79260 73951
0 27256 7 1 2 84431 27255
0 27257 5 1 1 27256
0 27258 7 1 2 27254 27257
0 27259 5 1 1 27258
0 27260 7 1 2 69248 27259
0 27261 5 1 1 27260
0 27262 7 1 2 27242 27261
0 27263 7 1 2 27233 27262
0 27264 5 1 1 27263
0 27265 7 1 2 87166 27264
0 27266 5 1 1 27265
0 27267 7 1 2 75081 92291
0 27268 7 1 2 93653 27267
0 27269 5 1 1 27268
0 27270 7 1 2 27266 27269
0 27271 5 1 1 27270
0 27272 7 1 2 63975 27271
0 27273 5 1 1 27272
0 27274 7 1 2 86363 86910
0 27275 7 1 2 85551 27274
0 27276 7 1 2 87705 27275
0 27277 5 1 1 27276
0 27278 7 1 2 27273 27277
0 27279 5 1 1 27278
0 27280 7 1 2 93763 27279
0 27281 5 1 1 27280
0 27282 7 1 2 73518 78533
0 27283 5 2 1 27282
0 27284 7 1 2 68004 93780
0 27285 5 1 1 27284
0 27286 7 1 2 75687 27285
0 27287 5 1 1 27286
0 27288 7 1 2 71008 73850
0 27289 5 1 1 27288
0 27290 7 1 2 76642 86006
0 27291 5 1 1 27290
0 27292 7 1 2 27289 27291
0 27293 5 1 1 27292
0 27294 7 1 2 71982 27293
0 27295 5 1 1 27294
0 27296 7 1 2 27287 27295
0 27297 5 1 1 27296
0 27298 7 1 2 64981 27297
0 27299 5 1 1 27298
0 27300 7 3 2 63018 73519
0 27301 5 1 1 93782
0 27302 7 1 2 81951 93783
0 27303 5 1 1 27302
0 27304 7 1 2 27299 27303
0 27305 5 1 1 27304
0 27306 7 1 2 64748 27305
0 27307 5 1 1 27306
0 27308 7 1 2 76868 86849
0 27309 7 1 2 91124 27308
0 27310 5 2 1 27309
0 27311 7 1 2 27307 93785
0 27312 5 1 1 27311
0 27313 7 1 2 93435 27312
0 27314 5 1 1 27313
0 27315 7 1 2 84151 83725
0 27316 5 1 1 27315
0 27317 7 2 2 83584 88084
0 27318 5 1 1 93787
0 27319 7 1 2 79561 75953
0 27320 7 1 2 93788 27319
0 27321 5 1 1 27320
0 27322 7 1 2 27316 27321
0 27323 5 1 1 27322
0 27324 7 1 2 62663 27323
0 27325 5 1 1 27324
0 27326 7 1 2 65425 91911
0 27327 5 1 1 27326
0 27328 7 1 2 81285 87586
0 27329 7 1 2 87694 27328
0 27330 5 1 1 27329
0 27331 7 1 2 27327 27330
0 27332 5 1 1 27331
0 27333 7 1 2 69249 27332
0 27334 5 1 1 27333
0 27335 7 2 2 62313 93778
0 27336 5 1 1 93789
0 27337 7 1 2 72770 85449
0 27338 7 1 2 93790 27337
0 27339 5 1 1 27338
0 27340 7 1 2 84371 84545
0 27341 5 5 1 27340
0 27342 7 1 2 84027 90900
0 27343 7 1 2 15168 27342
0 27344 7 1 2 93791 27343
0 27345 5 1 1 27344
0 27346 7 1 2 27339 27345
0 27347 7 1 2 27334 27346
0 27348 7 1 2 27325 27347
0 27349 5 1 1 27348
0 27350 7 1 2 63459 27349
0 27351 5 1 1 27350
0 27352 7 1 2 63744 85450
0 27353 7 1 2 73520 27352
0 27354 5 1 1 27353
0 27355 7 1 2 84775 88186
0 27356 7 1 2 90916 27355
0 27357 5 1 1 27356
0 27358 7 1 2 27354 27357
0 27359 5 1 1 27358
0 27360 7 1 2 79439 27359
0 27361 5 1 1 27360
0 27362 7 1 2 27351 27361
0 27363 5 1 1 27362
0 27364 7 1 2 77193 27363
0 27365 5 1 1 27364
0 27366 7 1 2 74508 78254
0 27367 5 1 1 27366
0 27368 7 1 2 84570 27367
0 27369 5 1 1 27368
0 27370 7 1 2 65426 27369
0 27371 5 1 1 27370
0 27372 7 1 2 7795 27371
0 27373 5 1 1 27372
0 27374 7 1 2 89773 27373
0 27375 5 1 1 27374
0 27376 7 1 2 85604 88218
0 27377 7 1 2 74501 27376
0 27378 5 1 1 27377
0 27379 7 1 2 27375 27378
0 27380 5 1 1 27379
0 27381 7 1 2 65214 27380
0 27382 5 1 1 27381
0 27383 7 1 2 87550 91410
0 27384 5 1 1 27383
0 27385 7 1 2 89446 27384
0 27386 5 1 1 27385
0 27387 7 1 2 69250 27386
0 27388 5 1 1 27387
0 27389 7 1 2 64516 89444
0 27390 5 1 1 27389
0 27391 7 1 2 86444 93487
0 27392 5 1 1 27391
0 27393 7 1 2 27390 27392
0 27394 7 1 2 27388 27393
0 27395 5 1 1 27394
0 27396 7 1 2 85137 27395
0 27397 5 1 1 27396
0 27398 7 1 2 27382 27397
0 27399 5 1 1 27398
0 27400 7 1 2 77864 27399
0 27401 5 1 1 27400
0 27402 7 1 2 60541 3938
0 27403 7 2 2 92416 27402
0 27404 5 1 1 93796
0 27405 7 1 2 89559 27404
0 27406 5 5 1 27405
0 27407 7 3 2 83636 74502
0 27408 7 1 2 63019 93803
0 27409 7 1 2 93798 27408
0 27410 5 1 1 27409
0 27411 7 1 2 27401 27410
0 27412 5 1 1 27411
0 27413 7 1 2 64749 27412
0 27414 5 1 1 27413
0 27415 7 1 2 91319 93426
0 27416 5 1 1 27415
0 27417 7 1 2 83714 27416
0 27418 5 1 1 27417
0 27419 7 1 2 63745 27418
0 27420 5 1 1 27419
0 27421 7 1 2 84184 82574
0 27422 5 1 1 27421
0 27423 7 1 2 66516 85145
0 27424 7 1 2 27422 27423
0 27425 5 1 1 27424
0 27426 7 1 2 65215 23129
0 27427 7 1 2 93399 27426
0 27428 7 1 2 27425 27427
0 27429 5 1 1 27428
0 27430 7 1 2 27420 27429
0 27431 5 1 1 27430
0 27432 7 1 2 61725 27431
0 27433 5 1 1 27432
0 27434 7 1 2 63746 81516
0 27435 5 1 1 27434
0 27436 7 1 2 27433 27435
0 27437 5 1 1 27436
0 27438 7 1 2 82371 27437
0 27439 5 1 1 27438
0 27440 7 2 2 91051 92266
0 27441 7 1 2 64517 93113
0 27442 7 1 2 93806 27441
0 27443 5 1 1 27442
0 27444 7 1 2 27439 27443
0 27445 5 1 1 27444
0 27446 7 1 2 66286 27445
0 27447 5 1 1 27446
0 27448 7 1 2 65427 77626
0 27449 7 1 2 92433 27448
0 27450 5 1 1 27449
0 27451 7 1 2 63460 27450
0 27452 7 1 2 27447 27451
0 27453 7 1 2 27414 27452
0 27454 5 1 1 27453
0 27455 7 1 2 70490 93807
0 27456 5 1 1 27455
0 27457 7 1 2 84163 91342
0 27458 5 1 1 27457
0 27459 7 1 2 27456 27458
0 27460 5 1 1 27459
0 27461 7 1 2 64750 27460
0 27462 5 1 1 27461
0 27463 7 2 2 83637 87924
0 27464 5 1 1 93808
0 27465 7 1 2 93497 93809
0 27466 5 1 1 27465
0 27467 7 1 2 27462 27466
0 27468 5 1 1 27467
0 27469 7 1 2 63020 27468
0 27470 5 1 1 27469
0 27471 7 1 2 62108 87792
0 27472 5 1 1 27471
0 27473 7 1 2 93579 27472
0 27474 5 1 1 27473
0 27475 7 1 2 81768 27474
0 27476 5 1 1 27475
0 27477 7 1 2 64982 88232
0 27478 7 1 2 92084 27477
0 27479 5 1 1 27478
0 27480 7 1 2 27476 27479
0 27481 7 1 2 27470 27480
0 27482 5 1 1 27481
0 27483 7 1 2 64518 27482
0 27484 5 1 1 27483
0 27485 7 1 2 84589 91194
0 27486 5 2 1 27485
0 27487 7 1 2 85146 93810
0 27488 5 1 1 27487
0 27489 7 1 2 65216 27488
0 27490 5 1 1 27489
0 27491 7 1 2 66031 85188
0 27492 7 1 2 93427 27491
0 27493 5 1 1 27492
0 27494 7 1 2 27490 27493
0 27495 5 1 1 27494
0 27496 7 1 2 66702 27495
0 27497 5 1 1 27496
0 27498 7 1 2 81769 84480
0 27499 5 1 1 27498
0 27500 7 1 2 27497 27499
0 27501 5 1 1 27500
0 27502 7 1 2 73568 27501
0 27503 5 1 1 27502
0 27504 7 2 2 78566 93367
0 27505 7 1 2 76986 84185
0 27506 5 1 1 27505
0 27507 7 1 2 65866 93582
0 27508 5 1 1 27507
0 27509 7 1 2 27506 27508
0 27510 5 1 1 27509
0 27511 7 1 2 93812 27510
0 27512 5 1 1 27511
0 27513 7 1 2 84633 93577
0 27514 5 1 1 27513
0 27515 7 1 2 27512 27514
0 27516 5 1 1 27515
0 27517 7 1 2 65217 27516
0 27518 5 1 1 27517
0 27519 7 1 2 27503 27518
0 27520 7 1 2 27484 27519
0 27521 5 1 1 27520
0 27522 7 1 2 66517 27521
0 27523 5 1 1 27522
0 27524 7 2 2 71782 93483
0 27525 5 1 1 93814
0 27526 7 1 2 84140 93815
0 27527 5 1 1 27526
0 27528 7 1 2 68358 27527
0 27529 7 1 2 27523 27528
0 27530 5 1 1 27529
0 27531 7 1 2 27454 27530
0 27532 5 1 1 27531
0 27533 7 1 2 27365 27532
0 27534 5 1 1 27533
0 27535 7 1 2 63976 27534
0 27536 5 1 1 27535
0 27537 7 2 2 27314 27536
0 27538 5 1 1 93816
0 27539 7 1 2 61864 93817
0 27540 5 1 1 27539
0 27541 7 1 2 70491 73891
0 27542 5 2 1 27541
0 27543 7 1 2 73587 93818
0 27544 5 1 1 27543
0 27545 7 1 2 66032 27544
0 27546 5 1 1 27545
0 27547 7 1 2 71983 88319
0 27548 5 1 1 27547
0 27549 7 1 2 27546 27548
0 27550 5 1 1 27549
0 27551 7 1 2 84222 27550
0 27552 5 1 1 27551
0 27553 7 1 2 82118 84947
0 27554 5 1 1 27553
0 27555 7 1 2 10334 27554
0 27556 5 1 1 27555
0 27557 7 1 2 60358 27556
0 27558 5 1 1 27557
0 27559 7 1 2 79886 77194
0 27560 5 1 1 27559
0 27561 7 1 2 27558 27560
0 27562 5 1 1 27561
0 27563 7 1 2 79620 27562
0 27564 5 1 1 27563
0 27565 7 1 2 68680 27564
0 27566 7 1 2 27552 27565
0 27567 5 1 1 27566
0 27568 7 1 2 73569 93799
0 27569 5 1 1 27568
0 27570 7 4 2 71783 75581
0 27571 7 2 2 62314 87829
0 27572 5 1 1 93824
0 27573 7 1 2 93820 93825
0 27574 5 1 1 27573
0 27575 7 1 2 84857 91052
0 27576 5 1 1 27575
0 27577 7 1 2 27574 27576
0 27578 5 1 1 27577
0 27579 7 1 2 77987 84253
0 27580 7 1 2 27578 27579
0 27581 5 1 1 27580
0 27582 7 1 2 27569 27581
0 27583 5 1 1 27582
0 27584 7 1 2 64983 27583
0 27585 5 1 1 27584
0 27586 7 1 2 82119 93797
0 27587 5 1 1 27586
0 27588 7 1 2 63747 27587
0 27589 7 1 2 27585 27588
0 27590 5 1 1 27589
0 27591 7 1 2 63021 27590
0 27592 7 1 2 27567 27591
0 27593 5 1 1 27592
0 27594 7 1 2 78945 93804
0 27595 5 1 1 27594
0 27596 7 1 2 79409 84640
0 27597 5 1 1 27596
0 27598 7 1 2 27595 27597
0 27599 5 1 1 27598
0 27600 7 1 2 80413 27599
0 27601 5 1 1 27600
0 27602 7 1 2 80868 82815
0 27603 7 1 2 93805 27602
0 27604 5 1 1 27603
0 27605 7 1 2 27601 27604
0 27606 5 1 1 27605
0 27607 7 1 2 77865 27606
0 27608 5 1 1 27607
0 27609 7 1 2 63461 27608
0 27610 7 1 2 27593 27609
0 27611 5 1 1 27610
0 27612 7 1 2 63748 91000
0 27613 7 1 2 93332 27612
0 27614 5 1 1 27613
0 27615 7 1 2 7745 27614
0 27616 5 1 1 27615
0 27617 7 1 2 75214 27616
0 27618 5 1 1 27617
0 27619 7 1 2 85249 85818
0 27620 7 1 2 84141 27619
0 27621 5 1 1 27620
0 27622 7 1 2 27618 27621
0 27623 5 1 1 27622
0 27624 7 1 2 64519 27623
0 27625 5 1 1 27624
0 27626 7 1 2 68681 69251
0 27627 7 1 2 92075 27626
0 27628 5 1 1 27627
0 27629 7 1 2 27625 27628
0 27630 5 1 1 27629
0 27631 7 1 2 66287 27630
0 27632 5 1 1 27631
0 27633 7 1 2 74279 79014
0 27634 7 1 2 79697 27633
0 27635 5 1 1 27634
0 27636 7 1 2 68359 27635
0 27637 7 1 2 27632 27636
0 27638 5 1 1 27637
0 27639 7 1 2 27611 27638
0 27640 5 1 1 27639
0 27641 7 1 2 68873 27640
0 27642 5 1 1 27641
0 27643 7 1 2 65218 93083
0 27644 5 1 1 27643
0 27645 7 1 2 86015 27644
0 27646 5 1 1 27645
0 27647 7 2 2 68360 74067
0 27648 7 1 2 27646 93826
0 27649 5 1 1 27648
0 27650 7 1 2 75497 77172
0 27651 5 2 1 27650
0 27652 7 1 2 71009 91109
0 27653 7 1 2 93828 27652
0 27654 5 1 1 27653
0 27655 7 1 2 27649 27654
0 27656 5 1 1 27655
0 27657 7 1 2 80869 27656
0 27658 5 1 1 27657
0 27659 7 1 2 75741 85908
0 27660 7 1 2 80414 27659
0 27661 7 1 2 85334 27660
0 27662 5 1 1 27661
0 27663 7 1 2 27658 27662
0 27664 5 1 1 27663
0 27665 7 1 2 68682 27664
0 27666 5 1 1 27665
0 27667 7 2 2 78374 78760
0 27668 5 2 1 93830
0 27669 7 1 2 88135 93831
0 27670 5 1 1 27669
0 27671 7 1 2 63977 27670
0 27672 7 1 2 27666 27671
0 27673 5 1 1 27672
0 27674 7 1 2 62664 27673
0 27675 7 1 2 27642 27674
0 27676 5 1 1 27675
0 27677 7 1 2 77834 86654
0 27678 5 1 1 27677
0 27679 7 1 2 86930 27678
0 27680 5 1 1 27679
0 27681 7 1 2 73105 27680
0 27682 5 1 1 27681
0 27683 7 1 2 66518 77078
0 27684 7 1 2 85429 27683
0 27685 5 1 1 27684
0 27686 7 1 2 27682 27685
0 27687 5 1 1 27686
0 27688 7 1 2 65867 27687
0 27689 5 1 1 27688
0 27690 7 1 2 80744 79545
0 27691 5 1 1 27690
0 27692 7 1 2 27689 27691
0 27693 5 1 1 27692
0 27694 7 1 2 61726 27693
0 27695 5 1 1 27694
0 27696 7 1 2 75082 86894
0 27697 5 1 1 27696
0 27698 7 1 2 27695 27697
0 27699 5 1 1 27698
0 27700 7 1 2 79137 27699
0 27701 5 1 1 27700
0 27702 7 3 2 81770 84762
0 27703 7 4 2 63022 80979
0 27704 7 1 2 87544 93837
0 27705 7 1 2 93834 27704
0 27706 5 1 1 27705
0 27707 7 1 2 27701 27706
0 27708 5 1 1 27707
0 27709 7 1 2 68683 27708
0 27710 5 1 1 27709
0 27711 7 1 2 66288 92796
0 27712 5 1 1 27711
0 27713 7 4 2 63749 75582
0 27714 7 1 2 72158 91110
0 27715 7 1 2 93841 27714
0 27716 5 1 1 27715
0 27717 7 1 2 66519 12166
0 27718 5 1 1 27717
0 27719 7 1 2 85314 20720
0 27720 7 1 2 27718 27719
0 27721 5 1 1 27720
0 27722 7 1 2 27716 27721
0 27723 5 1 1 27722
0 27724 7 1 2 74567 27723
0 27725 5 1 1 27724
0 27726 7 1 2 27712 27725
0 27727 5 1 1 27726
0 27728 7 1 2 80538 27727
0 27729 5 1 1 27728
0 27730 7 2 2 82929 86467
0 27731 5 1 1 93845
0 27732 7 1 2 61549 85078
0 27733 7 1 2 93846 27732
0 27734 5 1 1 27733
0 27735 7 1 2 27729 27734
0 27736 5 1 1 27735
0 27737 7 1 2 62109 27736
0 27738 5 1 1 27737
0 27739 7 1 2 66289 81254
0 27740 7 1 2 74568 27739
0 27741 7 1 2 85867 27740
0 27742 5 1 1 27741
0 27743 7 1 2 27738 27742
0 27744 5 1 1 27743
0 27745 7 1 2 81180 27744
0 27746 5 1 1 27745
0 27747 7 1 2 81756 82389
0 27748 5 1 1 27747
0 27749 7 1 2 80690 77498
0 27750 7 1 2 79587 27749
0 27751 7 1 2 85160 27750
0 27752 5 1 1 27751
0 27753 7 1 2 27748 27752
0 27754 5 1 1 27753
0 27755 7 1 2 83540 27754
0 27756 5 1 1 27755
0 27757 7 1 2 82033 84793
0 27758 5 1 1 27757
0 27759 7 1 2 27756 27758
0 27760 5 1 1 27759
0 27761 7 1 2 82575 27760
0 27762 5 1 1 27761
0 27763 7 1 2 64984 78892
0 27764 5 1 1 27763
0 27765 7 1 2 27301 27764
0 27766 5 1 1 27765
0 27767 7 2 2 79040 79539
0 27768 7 1 2 68874 81086
0 27769 7 1 2 93847 27768
0 27770 7 1 2 27766 27769
0 27771 5 1 1 27770
0 27772 7 1 2 66837 27771
0 27773 7 1 2 27762 27772
0 27774 7 1 2 27746 27773
0 27775 7 1 2 27710 27774
0 27776 7 1 2 27676 27775
0 27777 5 1 1 27776
0 27778 7 1 2 27540 27777
0 27779 5 1 1 27778
0 27780 7 3 2 85516 88196
0 27781 5 2 1 93849
0 27782 7 1 2 68684 86586
0 27783 5 1 1 27782
0 27784 7 1 2 93852 27783
0 27785 5 2 1 27784
0 27786 7 1 2 66290 83098
0 27787 7 2 2 93854 27786
0 27788 5 1 1 93856
0 27789 7 1 2 61727 92963
0 27790 5 1 1 27789
0 27791 7 1 2 27788 27790
0 27792 5 1 1 27791
0 27793 7 1 2 71784 27792
0 27794 5 1 1 27793
0 27795 7 1 2 84627 86468
0 27796 5 1 1 27795
0 27797 7 1 2 27794 27796
0 27798 5 1 1 27797
0 27799 7 1 2 66033 27798
0 27800 5 1 1 27799
0 27801 7 1 2 85337 86469
0 27802 5 1 1 27801
0 27803 7 1 2 27800 27802
0 27804 5 1 1 27803
0 27805 7 1 2 64751 27804
0 27806 5 1 1 27805
0 27807 7 1 2 72771 84345
0 27808 7 1 2 73851 27807
0 27809 5 1 1 27808
0 27810 7 1 2 12263 27809
0 27811 5 1 1 27810
0 27812 7 1 2 64520 27811
0 27813 5 1 1 27812
0 27814 7 2 2 63023 88197
0 27815 7 1 2 68685 93858
0 27816 5 1 1 27815
0 27817 7 1 2 27813 27816
0 27818 5 1 1 27817
0 27819 7 1 2 81020 27818
0 27820 5 1 1 27819
0 27821 7 1 2 27806 27820
0 27822 5 1 1 27821
0 27823 7 1 2 64985 27822
0 27824 5 1 1 27823
0 27825 7 1 2 11498 93586
0 27826 5 1 1 27825
0 27827 7 2 2 63024 81021
0 27828 7 1 2 73892 93860
0 27829 7 1 2 27826 27828
0 27830 5 1 1 27829
0 27831 7 1 2 27824 27830
0 27832 5 1 1 27831
0 27833 7 1 2 65428 27832
0 27834 5 1 1 27833
0 27835 7 2 2 92267 93225
0 27836 5 1 1 93862
0 27837 7 1 2 61865 27836
0 27838 7 1 2 27834 27837
0 27839 5 1 1 27838
0 27840 7 3 2 63025 80415
0 27841 7 1 2 80539 77988
0 27842 7 1 2 93864 27841
0 27843 5 1 1 27842
0 27844 7 1 2 4871 27843
0 27845 5 1 1 27844
0 27846 7 1 2 76185 27845
0 27847 5 1 1 27846
0 27848 7 1 2 64752 78193
0 27849 7 1 2 92424 27848
0 27850 5 1 1 27849
0 27851 7 1 2 27847 27850
0 27852 5 1 1 27851
0 27853 7 1 2 66034 27852
0 27854 5 1 1 27853
0 27855 7 1 2 63978 74224
0 27856 7 1 2 81732 27855
0 27857 5 1 1 27856
0 27858 7 1 2 27854 27857
0 27859 5 1 1 27858
0 27860 7 1 2 64986 27859
0 27861 5 1 1 27860
0 27862 7 1 2 68361 91173
0 27863 5 1 1 27862
0 27864 7 4 2 63462 78271
0 27865 5 4 1 93867
0 27866 7 1 2 81757 93871
0 27867 7 1 2 27863 27866
0 27868 5 1 1 27867
0 27869 7 1 2 27861 27868
0 27870 5 1 1 27869
0 27871 7 1 2 68686 27870
0 27872 5 1 1 27871
0 27873 7 1 2 83868 73852
0 27874 5 1 1 27873
0 27875 7 1 2 62110 81328
0 27876 5 1 1 27875
0 27877 7 1 2 27874 27876
0 27878 5 1 1 27877
0 27879 7 1 2 78761 88055
0 27880 7 1 2 27878 27879
0 27881 5 1 1 27880
0 27882 7 1 2 27872 27881
0 27883 5 1 1 27882
0 27884 7 1 2 71984 27883
0 27885 5 1 1 27884
0 27886 7 1 2 82677 87837
0 27887 5 1 1 27886
0 27888 7 1 2 66291 82678
0 27889 5 1 1 27888
0 27890 7 1 2 77499 27889
0 27891 5 3 1 27890
0 27892 7 1 2 84142 93875
0 27893 5 1 1 27892
0 27894 7 1 2 81910 74884
0 27895 7 1 2 85354 27894
0 27896 5 1 1 27895
0 27897 7 1 2 27893 27896
0 27898 5 1 1 27897
0 27899 7 1 2 68875 27898
0 27900 5 1 1 27899
0 27901 7 1 2 27887 27900
0 27902 5 1 1 27901
0 27903 7 1 2 66035 27902
0 27904 5 1 1 27903
0 27905 7 3 2 80870 77561
0 27906 5 1 1 93878
0 27907 7 1 2 93876 93879
0 27908 5 1 1 27907
0 27909 7 1 2 27904 27908
0 27910 5 1 1 27909
0 27911 7 1 2 64987 27910
0 27912 5 1 1 27911
0 27913 7 2 2 62665 92726
0 27914 5 1 1 93881
0 27915 7 1 2 81080 93882
0 27916 5 1 1 27915
0 27917 7 1 2 27912 27916
0 27918 5 1 1 27917
0 27919 7 1 2 68362 27918
0 27920 5 1 1 27919
0 27921 7 1 2 66838 27920
0 27922 7 1 2 27885 27921
0 27923 5 1 1 27922
0 27924 7 1 2 62315 27923
0 27925 7 1 2 27839 27924
0 27926 5 1 1 27925
0 27927 7 1 2 83638 89873
0 27928 7 1 2 93705 27927
0 27929 5 1 1 27928
0 27930 7 2 2 61866 86581
0 27931 5 2 1 93883
0 27932 7 1 2 68005 93698
0 27933 5 1 1 27932
0 27934 7 1 2 93885 27933
0 27935 5 1 1 27934
0 27936 7 4 2 65429 84776
0 27937 5 4 1 93887
0 27938 7 1 2 77835 93888
0 27939 7 1 2 27935 27938
0 27940 5 1 1 27939
0 27941 7 1 2 27929 27940
0 27942 5 1 1 27941
0 27943 7 1 2 68363 27942
0 27944 5 1 1 27943
0 27945 7 2 2 73479 86352
0 27946 5 1 1 93895
0 27947 7 1 2 90678 93896
0 27948 5 1 1 27947
0 27949 7 1 2 27944 27948
0 27950 5 1 1 27949
0 27951 7 1 2 66703 27950
0 27952 5 1 1 27951
0 27953 7 2 2 61728 81022
0 27954 5 1 1 93897
0 27955 7 2 2 84777 87206
0 27956 5 1 1 93899
0 27957 7 1 2 83639 86062
0 27958 5 1 1 27957
0 27959 7 1 2 27956 27958
0 27960 5 2 1 27959
0 27961 7 1 2 78567 93901
0 27962 5 1 1 27961
0 27963 7 1 2 84926 93900
0 27964 5 1 1 27963
0 27965 7 1 2 27962 27964
0 27966 5 1 1 27965
0 27967 7 1 2 93898 27966
0 27968 5 1 1 27967
0 27969 7 1 2 27952 27968
0 27970 5 1 1 27969
0 27971 7 1 2 71785 27970
0 27972 5 1 1 27971
0 27973 7 1 2 71985 93857
0 27974 5 1 1 27973
0 27975 7 1 2 81023 85200
0 27976 5 1 1 27975
0 27977 7 1 2 27974 27976
0 27978 5 1 1 27977
0 27979 7 1 2 61867 27978
0 27980 5 1 1 27979
0 27981 7 3 2 84346 86157
0 27982 5 1 1 93903
0 27983 7 2 2 74280 77471
0 27984 7 1 2 68364 93906
0 27985 7 1 2 93904 27984
0 27986 5 1 1 27985
0 27987 7 1 2 27980 27986
0 27988 5 1 1 27987
0 27989 7 1 2 66036 27988
0 27990 5 1 1 27989
0 27991 7 1 2 65868 85806
0 27992 7 1 2 93227 27991
0 27993 5 1 1 27992
0 27994 7 1 2 27990 27993
0 27995 5 1 1 27994
0 27996 7 1 2 64753 27995
0 27997 5 1 1 27996
0 27998 7 1 2 71986 84254
0 27999 7 1 2 86334 27998
0 28000 5 1 1 27999
0 28001 7 1 2 27997 28000
0 28002 5 1 1 28001
0 28003 7 1 2 81270 28002
0 28004 5 1 1 28003
0 28005 7 1 2 27972 28004
0 28006 7 1 2 27926 28005
0 28007 5 1 1 28006
0 28008 7 1 2 75583 28007
0 28009 5 1 1 28008
0 28010 7 1 2 65566 28009
0 28011 7 1 2 27779 28010
0 28012 5 1 1 28011
0 28013 7 1 2 66839 27538
0 28014 5 1 1 28013
0 28015 7 1 2 73106 73853
0 28016 5 1 1 28015
0 28017 7 1 2 91448 28016
0 28018 5 1 1 28017
0 28019 7 1 2 65869 28018
0 28020 5 1 1 28019
0 28021 7 2 2 62316 77989
0 28022 5 1 1 93908
0 28023 7 1 2 28020 28022
0 28024 5 1 1 28023
0 28025 7 1 2 81971 28024
0 28026 5 1 1 28025
0 28027 7 1 2 83128 78704
0 28028 5 1 1 28027
0 28029 7 1 2 28026 28028
0 28030 5 1 1 28029
0 28031 7 1 2 85325 28030
0 28032 5 1 1 28031
0 28033 7 1 2 71987 87609
0 28034 5 1 1 28033
0 28035 7 1 2 93373 28034
0 28036 5 1 1 28035
0 28037 7 1 2 64754 28036
0 28038 5 1 1 28037
0 28039 7 1 2 80752 90250
0 28040 5 1 1 28039
0 28041 7 1 2 28038 28040
0 28042 5 1 1 28041
0 28043 7 1 2 80330 28042
0 28044 5 1 1 28043
0 28045 7 1 2 79361 77161
0 28046 5 1 1 28045
0 28047 7 1 2 85112 28046
0 28048 5 1 1 28047
0 28049 7 1 2 71786 80416
0 28050 7 1 2 28048 28049
0 28051 5 1 1 28050
0 28052 7 1 2 28044 28051
0 28053 5 1 1 28052
0 28054 7 1 2 63750 28053
0 28055 5 1 1 28054
0 28056 7 1 2 68365 28055
0 28057 7 1 2 28032 28056
0 28058 5 1 1 28057
0 28059 7 2 2 81315 79015
0 28060 5 1 1 93910
0 28061 7 2 2 64521 79362
0 28062 7 1 2 91269 93912
0 28063 7 1 2 93911 28062
0 28064 5 1 1 28063
0 28065 7 1 2 86341 93721
0 28066 5 1 1 28065
0 28067 7 1 2 63463 28066
0 28068 7 1 2 28064 28067
0 28069 5 1 1 28068
0 28070 7 1 2 63979 28069
0 28071 7 1 2 28058 28070
0 28072 5 1 1 28071
0 28073 7 1 2 74020 93863
0 28074 5 1 1 28073
0 28075 7 1 2 80549 74835
0 28076 7 4 2 78705 85189
0 28077 7 1 2 80975 93914
0 28078 7 1 2 28075 28077
0 28079 5 1 1 28078
0 28080 7 1 2 28074 28079
0 28081 7 1 2 28072 28080
0 28082 5 1 1 28081
0 28083 7 1 2 66840 28082
0 28084 5 1 1 28083
0 28085 7 1 2 66704 79735
0 28086 7 2 2 76850 77472
0 28087 7 1 2 93616 93918
0 28088 7 1 2 28085 28087
0 28089 5 1 1 28088
0 28090 7 3 2 66705 83640
0 28091 7 1 2 87051 93920
0 28092 5 1 1 28091
0 28093 7 1 2 66292 66841
0 28094 7 1 2 93855 28093
0 28095 5 1 1 28094
0 28096 7 1 2 28092 28095
0 28097 5 1 1 28096
0 28098 7 1 2 86638 28097
0 28099 5 1 1 28098
0 28100 7 1 2 81024 86312
0 28101 7 1 2 87793 28100
0 28102 5 1 1 28101
0 28103 7 1 2 28099 28102
0 28104 5 1 1 28103
0 28105 7 1 2 74021 77866
0 28106 7 1 2 93534 28105
0 28107 7 1 2 28104 28106
0 28108 5 1 1 28107
0 28109 7 1 2 28089 28108
0 28110 7 1 2 28084 28109
0 28111 5 1 1 28110
0 28112 7 1 2 75584 28111
0 28113 5 1 1 28112
0 28114 7 2 2 65870 82679
0 28115 5 2 1 93923
0 28116 7 1 2 63026 93924
0 28117 5 1 1 28116
0 28118 7 1 2 93374 28117
0 28119 5 1 1 28118
0 28120 7 1 2 74022 28119
0 28121 5 1 1 28120
0 28122 7 1 2 65871 93368
0 28123 5 1 1 28122
0 28124 7 1 2 85568 28123
0 28125 7 1 2 28121 28124
0 28126 5 1 1 28125
0 28127 7 1 2 63464 28126
0 28128 5 1 1 28127
0 28129 7 1 2 27525 28128
0 28130 5 1 1 28129
0 28131 7 7 2 61868 87855
0 28132 7 1 2 79698 93927
0 28133 7 1 2 28130 28132
0 28134 5 1 1 28133
0 28135 7 1 2 60662 28134
0 28136 7 1 2 28113 28135
0 28137 7 1 2 28014 28136
0 28138 5 1 1 28137
0 28139 7 1 2 28012 28138
0 28140 5 1 1 28139
0 28141 7 1 2 27281 28140
0 28142 5 1 1 28141
0 28143 7 1 2 69658 28142
0 28144 5 1 1 28143
0 28145 7 1 2 69350 75041
0 28146 5 1 1 28145
0 28147 7 1 2 59340 28146
0 28148 5 1 1 28147
0 28149 7 1 2 63027 28148
0 28150 7 1 2 82214 28149
0 28151 5 1 1 28150
0 28152 7 1 2 87856 93868
0 28153 7 2 2 28151 28152
0 28154 7 1 2 85668 93934
0 28155 5 1 1 28154
0 28156 7 5 2 80029 85517
0 28157 7 1 2 78706 93936
0 28158 5 1 1 28157
0 28159 7 1 2 73652 92598
0 28160 5 1 1 28159
0 28161 7 2 2 68687 69564
0 28162 7 2 2 86664 93941
0 28163 5 1 1 93943
0 28164 7 1 2 83678 28163
0 28165 5 1 1 28164
0 28166 7 1 2 72116 28165
0 28167 5 1 1 28166
0 28168 7 1 2 74917 92450
0 28169 5 1 1 28168
0 28170 7 2 2 67072 83673
0 28171 5 1 1 93945
0 28172 7 1 2 28169 28171
0 28173 5 1 1 28172
0 28174 7 1 2 67324 28173
0 28175 5 1 1 28174
0 28176 7 1 2 69565 83842
0 28177 5 1 1 28176
0 28178 7 1 2 86430 92182
0 28179 5 1 1 28178
0 28180 7 1 2 28177 28179
0 28181 7 1 2 28175 28180
0 28182 7 1 2 28167 28181
0 28183 5 1 1 28182
0 28184 7 1 2 68366 28183
0 28185 5 1 1 28184
0 28186 7 1 2 28160 28185
0 28187 5 1 1 28186
0 28188 7 1 2 73480 28187
0 28189 5 1 1 28188
0 28190 7 1 2 28158 28189
0 28191 5 1 1 28190
0 28192 7 1 2 67639 28191
0 28193 5 1 1 28192
0 28194 7 1 2 83757 77562
0 28195 7 1 2 93736 28194
0 28196 5 1 1 28195
0 28197 7 1 2 74777 85556
0 28198 5 1 1 28197
0 28199 7 1 2 28196 28198
0 28200 7 1 2 28193 28199
0 28201 5 1 1 28200
0 28202 7 1 2 70183 28201
0 28203 5 1 1 28202
0 28204 7 3 2 75315 77563
0 28205 7 1 2 83027 93947
0 28206 5 1 1 28205
0 28207 7 2 2 86383 87262
0 28208 7 1 2 73675 69126
0 28209 7 1 2 93950 28208
0 28210 5 1 1 28209
0 28211 7 1 2 28206 28210
0 28212 5 1 1 28211
0 28213 7 1 2 59552 28212
0 28214 5 1 1 28213
0 28215 7 2 2 60926 82980
0 28216 7 1 2 92950 93952
0 28217 5 1 1 28216
0 28218 7 1 2 28214 28217
0 28219 5 1 1 28218
0 28220 7 1 2 63465 28219
0 28221 5 1 1 28220
0 28222 7 1 2 81095 83028
0 28223 7 1 2 89974 28222
0 28224 5 1 1 28223
0 28225 7 1 2 28221 28224
0 28226 5 1 1 28225
0 28227 7 1 2 67073 28226
0 28228 5 1 1 28227
0 28229 7 2 2 69188 77782
0 28230 5 1 1 93954
0 28231 7 1 2 15438 28230
0 28232 5 1 1 28231
0 28233 7 1 2 76779 28232
0 28234 5 1 1 28233
0 28235 7 1 2 83919 25798
0 28236 5 1 1 28235
0 28237 7 1 2 92818 28236
0 28238 5 1 1 28237
0 28239 7 1 2 28234 28238
0 28240 5 1 1 28239
0 28241 7 1 2 68688 28240
0 28242 5 1 1 28241
0 28243 7 2 2 78400 83843
0 28244 7 1 2 83743 93956
0 28245 5 1 1 28244
0 28246 7 1 2 28242 28245
0 28247 5 1 1 28246
0 28248 7 1 2 63980 28247
0 28249 5 1 1 28248
0 28250 7 1 2 28228 28249
0 28251 5 1 1 28250
0 28252 7 1 2 69922 28251
0 28253 5 1 1 28252
0 28254 7 1 2 74047 78568
0 28255 5 1 1 28254
0 28256 7 1 2 78912 28255
0 28257 5 1 1 28256
0 28258 7 1 2 66520 28257
0 28259 5 1 1 28258
0 28260 7 1 2 82981 74918
0 28261 7 1 2 74830 28260
0 28262 5 1 1 28261
0 28263 7 1 2 28259 28262
0 28264 5 1 1 28263
0 28265 7 1 2 85518 28264
0 28266 5 1 1 28265
0 28267 7 1 2 72117 77564
0 28268 7 1 2 84099 28267
0 28269 7 1 2 92411 28268
0 28270 5 1 1 28269
0 28271 7 1 2 28266 28270
0 28272 5 1 1 28271
0 28273 7 1 2 63466 28272
0 28274 5 1 1 28273
0 28275 7 1 2 74369 78970
0 28276 5 1 1 28275
0 28277 7 2 2 63028 74638
0 28278 5 1 1 93958
0 28279 7 1 2 81450 93959
0 28280 5 1 1 28279
0 28281 7 1 2 84839 90776
0 28282 7 1 2 28280 28281
0 28283 5 1 1 28282
0 28284 7 1 2 28276 28283
0 28285 5 1 1 28284
0 28286 7 1 2 86470 28285
0 28287 5 1 1 28286
0 28288 7 1 2 28274 28287
0 28289 7 1 2 28253 28288
0 28290 5 1 1 28289
0 28291 7 1 2 67640 28290
0 28292 5 1 1 28291
0 28293 7 1 2 89510 93336
0 28294 5 1 1 28293
0 28295 7 1 2 83500 28294
0 28296 5 1 1 28295
0 28297 7 1 2 77565 28296
0 28298 5 1 1 28297
0 28299 7 1 2 71988 83083
0 28300 5 1 1 28299
0 28301 7 1 2 92189 28300
0 28302 5 1 1 28301
0 28303 7 1 2 28298 28302
0 28304 5 1 1 28303
0 28305 7 1 2 63467 28304
0 28306 5 1 1 28305
0 28307 7 1 2 93321 93957
0 28308 5 1 1 28307
0 28309 7 1 2 73379 89785
0 28310 5 1 1 28309
0 28311 7 1 2 70184 70282
0 28312 7 1 2 83600 28311
0 28313 7 1 2 92183 28312
0 28314 5 1 1 28313
0 28315 7 1 2 28310 28314
0 28316 5 1 1 28315
0 28317 7 1 2 68689 28316
0 28318 5 1 1 28317
0 28319 7 1 2 28308 28318
0 28320 5 1 1 28319
0 28321 7 1 2 81025 28320
0 28322 5 1 1 28321
0 28323 7 1 2 28306 28322
0 28324 5 1 1 28323
0 28325 7 1 2 68006 28324
0 28326 5 1 1 28325
0 28327 7 2 2 67074 77783
0 28328 5 1 1 93960
0 28329 7 1 2 79811 28328
0 28330 5 2 1 28329
0 28331 7 1 2 72517 93962
0 28332 5 1 1 28331
0 28333 7 1 2 79872 92112
0 28334 5 1 1 28333
0 28335 7 1 2 69566 28334
0 28336 5 1 1 28335
0 28337 7 1 2 28332 28336
0 28338 5 1 1 28337
0 28339 7 1 2 76780 28338
0 28340 5 1 1 28339
0 28341 7 1 2 92109 93154
0 28342 5 1 1 28341
0 28343 7 1 2 28340 28342
0 28344 5 1 1 28343
0 28345 7 1 2 59553 28344
0 28346 5 1 1 28345
0 28347 7 2 2 75439 89058
0 28348 7 1 2 92412 93964
0 28349 5 1 1 28348
0 28350 7 1 2 28346 28349
0 28351 5 1 1 28350
0 28352 7 1 2 63981 91894
0 28353 7 1 2 28351 28352
0 28354 5 1 1 28353
0 28355 7 1 2 28326 28354
0 28356 7 1 2 28292 28355
0 28357 7 1 2 28203 28356
0 28358 5 1 1 28357
0 28359 7 1 2 66842 28358
0 28360 5 1 1 28359
0 28361 7 1 2 28155 28360
0 28362 5 1 1 28361
0 28363 7 1 2 65567 28362
0 28364 5 1 1 28363
0 28365 7 4 2 60663 87991
0 28366 7 1 2 93935 93966
0 28367 5 1 1 28366
0 28368 7 3 2 70185 92232
0 28369 5 1 1 93970
0 28370 7 1 2 88059 93971
0 28371 5 1 1 28370
0 28372 7 5 2 61869 63029
0 28373 7 2 2 66521 93973
0 28374 5 1 1 93978
0 28375 7 1 2 63751 93979
0 28376 5 1 1 28375
0 28377 7 1 2 28371 28376
0 28378 5 1 1 28377
0 28379 7 1 2 65568 28378
0 28380 5 1 1 28379
0 28381 7 1 2 79377 93967
0 28382 5 1 1 28381
0 28383 7 1 2 28380 28382
0 28384 5 1 1 28383
0 28385 7 1 2 67075 28384
0 28386 5 1 1 28385
0 28387 7 1 2 76781 86996
0 28388 7 1 2 92824 28387
0 28389 5 1 1 28388
0 28390 7 1 2 28386 28389
0 28391 5 1 1 28390
0 28392 7 1 2 63468 28391
0 28393 5 1 1 28392
0 28394 7 1 2 81134 91131
0 28395 5 1 1 28394
0 28396 7 1 2 90044 28395
0 28397 5 1 1 28396
0 28398 7 5 2 59554 66843
0 28399 7 3 2 65569 67641
0 28400 5 1 1 93985
0 28401 7 2 2 93980 93986
0 28402 7 1 2 89929 93988
0 28403 7 1 2 28397 28402
0 28404 5 1 1 28403
0 28405 7 1 2 28393 28404
0 28406 5 1 1 28405
0 28407 7 1 2 69923 28406
0 28408 5 1 1 28407
0 28409 7 1 2 20110 90092
0 28410 5 1 1 28409
0 28411 7 1 2 88150 28410
0 28412 5 1 1 28411
0 28413 7 1 2 28408 28412
0 28414 5 1 1 28413
0 28415 7 1 2 63982 28414
0 28416 5 1 1 28415
0 28417 7 3 2 69567 92810
0 28418 7 1 2 78194 86313
0 28419 7 1 2 93937 28418
0 28420 7 1 2 93990 28419
0 28421 5 1 1 28420
0 28422 7 1 2 28416 28421
0 28423 5 1 1 28422
0 28424 7 1 2 69127 28423
0 28425 5 1 1 28424
0 28426 7 1 2 28367 28425
0 28427 7 1 2 28364 28426
0 28428 5 1 1 28427
0 28429 7 1 2 71222 28428
0 28430 5 1 1 28429
0 28431 7 1 2 89984 93155
0 28432 5 1 1 28431
0 28433 7 1 2 71492 89986
0 28434 5 1 1 28433
0 28435 7 1 2 78762 88107
0 28436 7 1 2 74798 28435
0 28437 5 1 1 28436
0 28438 7 1 2 28434 28437
0 28439 5 1 1 28438
0 28440 7 1 2 72985 28439
0 28441 5 1 1 28440
0 28442 7 1 2 28432 28441
0 28443 5 1 1 28442
0 28444 7 1 2 71724 28443
0 28445 5 1 1 28444
0 28446 7 1 2 74170 89888
0 28447 7 1 2 92589 28446
0 28448 5 1 1 28447
0 28449 7 1 2 28445 28448
0 28450 5 1 1 28449
0 28451 7 1 2 67642 28450
0 28452 5 1 1 28451
0 28453 7 2 2 73417 92890
0 28454 5 1 1 93993
0 28455 7 1 2 83416 4910
0 28456 5 1 1 28455
0 28457 7 1 2 61550 28456
0 28458 5 1 1 28457
0 28459 7 1 2 28454 28458
0 28460 5 1 1 28459
0 28461 7 1 2 68690 28460
0 28462 5 1 1 28461
0 28463 7 1 2 28452 28462
0 28464 5 1 1 28463
0 28465 7 1 2 63983 28464
0 28466 5 1 1 28465
0 28467 7 1 2 92704 92882
0 28468 5 1 1 28467
0 28469 7 1 2 69826 87971
0 28470 7 1 2 91998 28469
0 28471 5 1 1 28470
0 28472 7 1 2 28468 28471
0 28473 5 1 1 28472
0 28474 7 1 2 62666 28473
0 28475 5 1 1 28474
0 28476 7 1 2 73873 92002
0 28477 5 1 1 28476
0 28478 7 1 2 28475 28477
0 28479 5 1 1 28478
0 28480 7 1 2 65872 28479
0 28481 5 1 1 28480
0 28482 7 1 2 68007 28481
0 28483 7 1 2 28466 28482
0 28484 5 1 1 28483
0 28485 7 1 2 4976 91032
0 28486 5 1 1 28485
0 28487 7 1 2 67325 28486
0 28488 5 1 1 28487
0 28489 7 1 2 80209 79168
0 28490 7 1 2 28488 28489
0 28491 5 1 1 28490
0 28492 7 1 2 93938 28491
0 28493 5 1 1 28492
0 28494 7 2 2 78324 25777
0 28495 5 1 1 93995
0 28496 7 1 2 83597 93996
0 28497 5 1 1 28496
0 28498 7 2 2 86471 90464
0 28499 7 1 2 28497 93997
0 28500 5 1 1 28499
0 28501 7 1 2 63030 28500
0 28502 7 1 2 28493 28501
0 28503 5 1 1 28502
0 28504 7 1 2 28484 28503
0 28505 5 1 1 28504
0 28506 7 1 2 73624 73632
0 28507 5 1 1 28506
0 28508 7 1 2 93939 28507
0 28509 5 1 1 28508
0 28510 7 1 2 74522 93998
0 28511 5 1 1 28510
0 28512 7 1 2 28509 28511
0 28513 5 1 1 28512
0 28514 7 1 2 82864 28513
0 28515 5 1 1 28514
0 28516 7 3 2 63469 72986
0 28517 7 1 2 72118 92705
0 28518 7 1 2 93999 28517
0 28519 5 1 1 28518
0 28520 7 1 2 28515 28519
0 28521 5 1 1 28520
0 28522 7 1 2 69924 28521
0 28523 5 1 1 28522
0 28524 7 3 2 63984 92956
0 28525 7 1 2 72468 76979
0 28526 5 1 1 28525
0 28527 7 1 2 72987 28526
0 28528 5 1 1 28527
0 28529 7 1 2 71401 28528
0 28530 5 1 1 28529
0 28531 7 1 2 94002 28530
0 28532 5 1 1 28531
0 28533 7 1 2 92201 28532
0 28534 5 1 1 28533
0 28535 7 1 2 63470 28534
0 28536 5 1 1 28535
0 28537 7 1 2 28523 28536
0 28538 7 1 2 28505 28537
0 28539 5 1 1 28538
0 28540 7 1 2 61344 28539
0 28541 5 1 1 28540
0 28542 7 1 2 69925 83406
0 28543 5 1 1 28542
0 28544 7 1 2 81554 83601
0 28545 5 1 1 28544
0 28546 7 1 2 28543 28545
0 28547 5 1 1 28546
0 28548 7 1 2 72119 28547
0 28549 5 1 1 28548
0 28550 7 1 2 81555 82554
0 28551 5 1 1 28550
0 28552 7 1 2 15103 28551
0 28553 7 1 2 28549 28552
0 28554 7 1 2 60805 81556
0 28555 5 1 1 28554
0 28556 7 1 2 83417 28555
0 28557 5 1 1 28556
0 28558 7 1 2 71989 73454
0 28559 5 2 1 28558
0 28560 7 1 2 73536 94005
0 28561 7 1 2 28557 28560
0 28562 5 1 1 28561
0 28563 7 1 2 77609 78335
0 28564 5 1 1 28563
0 28565 7 1 2 69343 83407
0 28566 5 1 1 28565
0 28567 7 1 2 28564 28566
0 28568 5 1 1 28567
0 28569 7 1 2 79839 28568
0 28570 5 1 1 28569
0 28571 7 1 2 67076 77617
0 28572 5 1 1 28571
0 28573 7 1 2 83418 28572
0 28574 5 1 1 28573
0 28575 7 1 2 67643 28574
0 28576 5 1 1 28575
0 28577 7 1 2 28570 28576
0 28578 7 1 2 28562 28577
0 28579 7 1 2 28553 28578
0 28580 5 1 1 28579
0 28581 7 1 2 61551 28580
0 28582 5 1 1 28581
0 28583 7 1 2 73973 72230
0 28584 5 2 1 28583
0 28585 7 1 2 68367 80797
0 28586 5 1 1 28585
0 28587 7 1 2 94007 28586
0 28588 5 1 1 28587
0 28589 7 1 2 94006 28588
0 28590 5 1 1 28589
0 28591 7 1 2 79840 89127
0 28592 7 1 2 83323 28591
0 28593 5 1 1 28592
0 28594 7 2 2 71787 82894
0 28595 5 1 1 94009
0 28596 7 1 2 75845 28595
0 28597 5 1 1 28596
0 28598 7 1 2 28593 28597
0 28599 7 1 2 28590 28598
0 28600 5 1 1 28599
0 28601 7 1 2 67326 28600
0 28602 5 1 1 28601
0 28603 7 1 2 73238 92895
0 28604 5 1 1 28603
0 28605 7 1 2 84756 94008
0 28606 5 1 1 28605
0 28607 7 1 2 67644 28606
0 28608 5 1 1 28607
0 28609 7 1 2 28604 28608
0 28610 7 1 2 28602 28609
0 28611 5 1 1 28610
0 28612 7 1 2 60359 28611
0 28613 5 1 1 28612
0 28614 7 1 2 69926 72194
0 28615 5 1 1 28614
0 28616 7 1 2 74639 81480
0 28617 7 1 2 81451 28616
0 28618 7 1 2 28615 28617
0 28619 5 1 1 28618
0 28620 7 1 2 93994 28619
0 28621 5 1 1 28620
0 28622 7 1 2 28613 28621
0 28623 7 1 2 28582 28622
0 28624 5 1 1 28623
0 28625 7 1 2 68008 28624
0 28626 5 1 1 28625
0 28627 7 1 2 79774 72836
0 28628 7 1 2 72988 28627
0 28629 5 1 1 28628
0 28630 7 1 2 70283 92110
0 28631 7 1 2 90465 28630
0 28632 5 1 1 28631
0 28633 7 1 2 28629 28632
0 28634 5 1 1 28633
0 28635 7 1 2 59555 28634
0 28636 5 1 1 28635
0 28637 7 2 2 79828 76346
0 28638 7 1 2 94000 94011
0 28639 5 1 1 28638
0 28640 7 1 2 28636 28639
0 28641 5 1 1 28640
0 28642 7 1 2 59341 28641
0 28643 5 1 1 28642
0 28644 7 1 2 92632 94001
0 28645 5 1 1 28644
0 28646 7 1 2 28643 28645
0 28647 5 1 1 28646
0 28648 7 1 2 71360 28647
0 28649 5 1 1 28648
0 28650 7 1 2 81538 83616
0 28651 5 1 1 28650
0 28652 7 1 2 28649 28651
0 28653 7 1 2 28626 28652
0 28654 5 1 1 28653
0 28655 7 1 2 68691 28654
0 28656 5 1 1 28655
0 28657 7 2 2 63752 76675
0 28658 7 1 2 69044 94013
0 28659 5 1 1 28658
0 28660 7 1 2 62667 92997
0 28661 5 1 1 28660
0 28662 7 1 2 83541 28661
0 28663 5 1 1 28662
0 28664 7 1 2 28659 28663
0 28665 5 1 1 28664
0 28666 7 1 2 60156 28665
0 28667 5 1 1 28666
0 28668 7 1 2 68692 81557
0 28669 5 1 1 28668
0 28670 7 1 2 28667 28669
0 28671 5 1 1 28670
0 28672 7 1 2 61552 88730
0 28673 7 1 2 28671 28672
0 28674 5 1 1 28673
0 28675 7 1 2 28656 28674
0 28676 5 1 1 28675
0 28677 7 1 2 63985 28676
0 28678 5 1 1 28677
0 28679 7 1 2 59556 71372
0 28680 7 1 2 74533 28679
0 28681 5 1 1 28680
0 28682 7 1 2 76601 28681
0 28683 5 1 1 28682
0 28684 7 1 2 60927 28683
0 28685 5 1 1 28684
0 28686 7 1 2 72855 83422
0 28687 5 1 1 28686
0 28688 7 1 2 73616 73239
0 28689 5 1 1 28688
0 28690 7 1 2 28687 28689
0 28691 7 1 2 28685 28690
0 28692 5 1 1 28691
0 28693 7 1 2 68009 28692
0 28694 5 1 1 28693
0 28695 7 1 2 73625 72231
0 28696 7 1 2 87365 28695
0 28697 5 1 1 28696
0 28698 7 1 2 28694 28697
0 28699 5 1 1 28698
0 28700 7 1 2 66293 28699
0 28701 5 1 1 28700
0 28702 7 3 2 74151 78433
0 28703 5 1 1 94015
0 28704 7 1 2 78913 28703
0 28705 5 1 1 28704
0 28706 7 1 2 60157 28705
0 28707 5 1 1 28706
0 28708 7 1 2 63031 90485
0 28709 5 1 1 28708
0 28710 7 1 2 63471 28709
0 28711 7 1 2 28707 28710
0 28712 7 1 2 28701 28711
0 28713 5 1 1 28712
0 28714 7 1 2 61345 93925
0 28715 5 1 1 28714
0 28716 7 1 2 93212 28715
0 28717 5 1 1 28716
0 28718 7 4 2 64755 78569
0 28719 5 2 1 94018
0 28720 7 1 2 80439 94019
0 28721 5 1 1 28720
0 28722 7 1 2 68010 1670
0 28723 5 1 1 28722
0 28724 7 1 2 93384 28723
0 28725 5 1 1 28724
0 28726 7 1 2 28721 28725
0 28727 7 1 2 28717 28726
0 28728 5 1 1 28727
0 28729 7 1 2 64522 28728
0 28730 5 1 1 28729
0 28731 7 1 2 82694 82583
0 28732 5 1 1 28731
0 28733 7 1 2 28730 28732
0 28734 5 1 1 28733
0 28735 7 1 2 62317 28734
0 28736 5 1 1 28735
0 28737 7 2 2 59902 76782
0 28738 5 1 1 94024
0 28739 7 1 2 63032 93385
0 28740 7 1 2 28738 28739
0 28741 5 1 1 28740
0 28742 7 1 2 80201 77966
0 28743 5 1 1 28742
0 28744 7 1 2 68368 28743
0 28745 7 1 2 28741 28744
0 28746 7 1 2 28736 28745
0 28747 5 1 1 28746
0 28748 7 1 2 66522 28747
0 28749 7 1 2 28713 28748
0 28750 5 1 1 28749
0 28751 7 1 2 79812 87752
0 28752 5 2 1 28751
0 28753 7 1 2 78594 93375
0 28754 5 1 1 28753
0 28755 7 1 2 94026 28754
0 28756 5 1 1 28755
0 28757 7 1 2 73792 85620
0 28758 5 1 1 28757
0 28759 7 1 2 28756 28758
0 28760 5 1 1 28759
0 28761 7 1 2 65873 28760
0 28762 5 1 1 28761
0 28763 7 1 2 85616 90698
0 28764 5 1 1 28763
0 28765 7 1 2 79813 26400
0 28766 5 1 1 28765
0 28767 7 1 2 84650 85113
0 28768 5 1 1 28767
0 28769 7 1 2 28766 28768
0 28770 5 1 1 28769
0 28771 7 1 2 28764 28770
0 28772 7 1 2 28762 28771
0 28773 5 1 1 28772
0 28774 7 1 2 73107 28773
0 28775 5 1 1 28774
0 28776 7 1 2 82949 93386
0 28777 5 1 1 28776
0 28778 7 1 2 76828 85106
0 28779 5 1 1 28778
0 28780 7 1 2 28777 28779
0 28781 5 1 1 28780
0 28782 7 1 2 79775 28781
0 28783 5 1 1 28782
0 28784 7 1 2 85944 93328
0 28785 5 1 1 28784
0 28786 7 1 2 28783 28785
0 28787 7 1 2 28775 28786
0 28788 5 1 1 28787
0 28789 7 1 2 64756 28788
0 28790 5 1 1 28789
0 28791 7 1 2 81225 86674
0 28792 5 1 1 28791
0 28793 7 1 2 73108 90722
0 28794 7 1 2 88326 28793
0 28795 5 1 1 28794
0 28796 7 1 2 28792 28795
0 28797 5 1 1 28796
0 28798 7 1 2 65219 28797
0 28799 5 1 1 28798
0 28800 7 1 2 83794 91095
0 28801 5 1 1 28800
0 28802 7 1 2 93376 28801
0 28803 5 1 1 28802
0 28804 7 1 2 83099 86414
0 28805 7 1 2 28803 28804
0 28806 5 1 1 28805
0 28807 7 1 2 28799 28806
0 28808 7 1 2 28790 28807
0 28809 7 1 2 28750 28808
0 28810 5 1 1 28809
0 28811 7 1 2 63753 28810
0 28812 5 1 1 28811
0 28813 7 2 2 73176 83875
0 28814 5 1 1 94028
0 28815 7 1 2 73109 28814
0 28816 5 1 1 28815
0 28817 7 1 2 91174 28816
0 28818 5 1 1 28817
0 28819 7 1 2 65874 28818
0 28820 5 1 1 28819
0 28821 7 1 2 68011 82255
0 28822 5 1 1 28821
0 28823 7 1 2 73169 28822
0 28824 5 1 1 28823
0 28825 7 1 2 28820 28824
0 28826 5 1 1 28825
0 28827 7 2 2 84866 93329
0 28828 7 1 2 28826 94030
0 28829 5 1 1 28828
0 28830 7 1 2 28812 28829
0 28831 5 1 1 28830
0 28832 7 1 2 68876 28831
0 28833 5 1 1 28832
0 28834 7 1 2 28678 28833
0 28835 7 1 2 28541 28834
0 28836 5 1 1 28835
0 28837 7 1 2 86707 28836
0 28838 5 1 1 28837
0 28839 7 2 2 79709 87313
0 28840 7 1 2 80030 94032
0 28841 5 1 1 28840
0 28842 7 1 2 73617 93951
0 28843 5 2 1 28842
0 28844 7 2 2 77473 91999
0 28845 5 1 1 94036
0 28846 7 1 2 60928 94037
0 28847 5 1 1 28846
0 28848 7 1 2 89671 93948
0 28849 5 1 1 28848
0 28850 7 1 2 28847 28849
0 28851 5 1 1 28850
0 28852 7 1 2 67327 28851
0 28853 5 1 1 28852
0 28854 7 1 2 94034 28853
0 28855 5 1 1 28854
0 28856 7 1 2 67077 28855
0 28857 5 1 1 28856
0 28858 7 1 2 78296 89829
0 28859 5 1 1 28858
0 28860 7 1 2 61346 28859
0 28861 5 1 1 28860
0 28862 7 1 2 14779 28861
0 28863 5 1 1 28862
0 28864 7 1 2 94003 28863
0 28865 5 1 1 28864
0 28866 7 1 2 28857 28865
0 28867 5 1 1 28866
0 28868 7 1 2 63472 28867
0 28869 5 1 1 28868
0 28870 7 1 2 92206 88340
0 28871 5 1 1 28870
0 28872 7 1 2 27731 28871
0 28873 5 1 1 28872
0 28874 7 1 2 84619 28873
0 28875 5 1 1 28874
0 28876 7 1 2 60360 93963
0 28877 5 1 1 28876
0 28878 7 1 2 63033 89427
0 28879 5 1 1 28878
0 28880 7 1 2 28877 28879
0 28881 5 1 1 28880
0 28882 7 1 2 77566 28881
0 28883 5 1 1 28882
0 28884 7 1 2 28875 28883
0 28885 5 1 1 28884
0 28886 7 1 2 69128 28885
0 28887 5 1 1 28886
0 28888 7 1 2 75050 90034
0 28889 5 2 1 28888
0 28890 7 1 2 69309 89623
0 28891 5 1 1 28890
0 28892 7 1 2 94038 28891
0 28893 5 1 1 28892
0 28894 7 1 2 68693 28893
0 28895 5 1 1 28894
0 28896 7 1 2 83440 89782
0 28897 7 1 2 93726 28896
0 28898 5 1 1 28897
0 28899 7 1 2 28895 28898
0 28900 5 1 1 28899
0 28901 7 1 2 81026 28900
0 28902 5 1 1 28901
0 28903 7 1 2 28887 28902
0 28904 7 1 2 28869 28903
0 28905 5 1 1 28904
0 28906 7 1 2 69927 28905
0 28907 5 1 1 28906
0 28908 7 1 2 76676 83844
0 28909 5 1 1 28908
0 28910 7 1 2 70535 89774
0 28911 7 1 2 72475 28910
0 28912 5 1 1 28911
0 28913 7 1 2 28909 28912
0 28914 5 1 1 28913
0 28915 7 1 2 61347 28914
0 28916 5 1 1 28915
0 28917 7 1 2 86669 91895
0 28918 5 1 1 28917
0 28919 7 1 2 83441 86269
0 28920 5 1 1 28919
0 28921 7 1 2 28918 28920
0 28922 5 1 1 28921
0 28923 7 1 2 69568 28922
0 28924 5 1 1 28923
0 28925 7 3 2 59557 79887
0 28926 5 1 1 94040
0 28927 7 1 2 69466 92061
0 28928 7 1 2 94041 28927
0 28929 5 1 1 28928
0 28930 7 1 2 14835 28929
0 28931 5 1 1 28930
0 28932 7 1 2 60361 28931
0 28933 5 1 1 28932
0 28934 7 1 2 28924 28933
0 28935 7 1 2 28916 28934
0 28936 5 1 1 28935
0 28937 7 1 2 68369 28936
0 28938 5 1 1 28937
0 28939 7 1 2 75788 82765
0 28940 5 1 1 28939
0 28941 7 1 2 73920 28940
0 28942 5 1 1 28941
0 28943 7 1 2 75316 28942
0 28944 5 1 1 28943
0 28945 7 1 2 80769 28944
0 28946 5 1 1 28945
0 28947 7 1 2 83542 28946
0 28948 5 1 1 28947
0 28949 7 1 2 28938 28948
0 28950 5 1 1 28949
0 28951 7 1 2 68012 28950
0 28952 5 1 1 28951
0 28953 7 1 2 63473 72476
0 28954 7 1 2 87952 28953
0 28955 5 1 1 28954
0 28956 7 1 2 28952 28955
0 28957 5 1 1 28956
0 28958 7 1 2 63986 28957
0 28959 5 1 1 28958
0 28960 7 3 2 70284 83047
0 28961 5 1 1 94043
0 28962 7 1 2 71361 86472
0 28963 7 1 2 94044 28962
0 28964 5 1 1 28963
0 28965 7 1 2 20799 28964
0 28966 5 1 1 28965
0 28967 7 1 2 61348 28966
0 28968 5 1 1 28967
0 28969 7 1 2 92204 28495
0 28970 5 1 1 28969
0 28971 7 1 2 63474 81820
0 28972 7 1 2 87884 28971
0 28973 5 1 1 28972
0 28974 7 1 2 28970 28973
0 28975 7 1 2 28968 28974
0 28976 5 1 1 28975
0 28977 7 1 2 63034 28976
0 28978 5 1 1 28977
0 28979 7 1 2 68694 91521
0 28980 5 1 1 28979
0 28981 7 1 2 74634 84844
0 28982 5 1 1 28981
0 28983 7 1 2 2704 28982
0 28984 5 1 1 28983
0 28985 7 1 2 60362 28984
0 28986 5 1 1 28985
0 28987 7 1 2 28980 28986
0 28988 5 1 1 28987
0 28989 7 1 2 81503 28988
0 28990 5 1 1 28989
0 28991 7 1 2 87907 89893
0 28992 5 1 1 28991
0 28993 7 1 2 28992 28845
0 28994 5 1 1 28993
0 28995 7 1 2 69569 28994
0 28996 5 1 1 28995
0 28997 7 1 2 83471 86843
0 28998 7 1 2 93949 28997
0 28999 5 1 1 28998
0 29000 7 1 2 28996 28999
0 29001 5 1 1 29000
0 29002 7 1 2 67328 29001
0 29003 5 1 1 29002
0 29004 7 1 2 82757 86431
0 29005 5 1 1 29004
0 29006 7 1 2 94035 29005
0 29007 7 1 2 29003 29006
0 29008 5 1 1 29007
0 29009 7 1 2 63475 29008
0 29010 5 1 1 29009
0 29011 7 1 2 28990 29010
0 29012 5 1 1 29011
0 29013 7 1 2 72120 29012
0 29014 5 1 1 29013
0 29015 7 1 2 28978 29014
0 29016 7 1 2 28959 29015
0 29017 7 1 2 28907 29016
0 29018 5 1 1 29017
0 29019 7 1 2 66844 29018
0 29020 5 1 1 29019
0 29021 7 1 2 28841 29020
0 29022 5 1 1 29021
0 29023 7 1 2 65570 29022
0 29024 5 1 1 29023
0 29025 7 1 2 79041 87314
0 29026 7 1 2 93968 29025
0 29027 5 1 1 29026
0 29028 7 1 2 29024 29027
0 29029 5 1 1 29028
0 29030 7 1 2 72936 29029
0 29031 5 1 1 29030
0 29032 7 1 2 81649 1798
0 29033 5 1 1 29032
0 29034 7 1 2 75585 29033
0 29035 5 1 1 29034
0 29036 7 1 2 76705 93360
0 29037 5 1 1 29036
0 29038 7 1 2 86917 29037
0 29039 5 1 1 29038
0 29040 7 1 2 64988 29039
0 29041 5 1 1 29040
0 29042 7 1 2 2670 29041
0 29043 5 1 1 29042
0 29044 7 1 2 63035 29043
0 29045 5 1 1 29044
0 29046 7 1 2 29035 29045
0 29047 5 1 1 29046
0 29048 7 1 2 62668 29047
0 29049 5 1 1 29048
0 29050 7 2 2 69827 70800
0 29051 5 1 1 94046
0 29052 7 1 2 12565 29051
0 29053 5 1 1 29052
0 29054 7 1 2 64757 29053
0 29055 5 1 1 29054
0 29056 7 2 2 76829 86911
0 29057 5 1 1 94048
0 29058 7 1 2 29055 29057
0 29059 5 1 1 29058
0 29060 7 1 2 75418 29059
0 29061 5 1 1 29060
0 29062 7 1 2 29049 29061
0 29063 5 1 1 29062
0 29064 7 1 2 62318 29063
0 29065 5 1 1 29064
0 29066 7 1 2 93086 26424
0 29067 5 1 1 29066
0 29068 7 1 2 65875 29067
0 29069 5 1 1 29068
0 29070 7 1 2 94022 29069
0 29071 5 1 1 29070
0 29072 7 1 2 77352 29071
0 29073 5 1 1 29072
0 29074 7 1 2 29065 29073
0 29075 5 1 1 29074
0 29076 7 1 2 66037 29075
0 29077 5 1 1 29076
0 29078 7 1 2 76718 93511
0 29079 5 1 1 29078
0 29080 7 1 2 78595 85054
0 29081 5 1 1 29080
0 29082 7 1 2 64758 29081
0 29083 5 1 1 29082
0 29084 7 1 2 79352 91111
0 29085 7 1 2 29083 29084
0 29086 7 1 2 29079 29085
0 29087 5 1 1 29086
0 29088 7 1 2 65220 29087
0 29089 5 1 1 29088
0 29090 7 1 2 82098 93505
0 29091 5 1 1 29090
0 29092 7 1 2 68370 29091
0 29093 7 1 2 29089 29092
0 29094 7 1 2 29077 29093
0 29095 5 1 1 29094
0 29096 7 1 2 8228 93601
0 29097 5 1 1 29096
0 29098 7 1 2 64759 29097
0 29099 5 1 1 29098
0 29100 7 1 2 60158 77204
0 29101 5 1 1 29100
0 29102 7 1 2 61553 29101
0 29103 5 1 1 29102
0 29104 7 1 2 29099 29103
0 29105 5 1 1 29104
0 29106 7 1 2 66294 29105
0 29107 5 1 1 29106
0 29108 7 1 2 77079 93599
0 29109 5 1 1 29108
0 29110 7 1 2 4001 29109
0 29111 7 1 2 29107 29110
0 29112 5 1 1 29111
0 29113 7 1 2 62669 29112
0 29114 5 1 1 29113
0 29115 7 1 2 67645 93322
0 29116 5 1 1 29115
0 29117 7 1 2 71493 90009
0 29118 5 1 1 29117
0 29119 7 1 2 79562 29118
0 29120 7 1 2 29116 29119
0 29121 5 1 1 29120
0 29122 7 1 2 72557 91036
0 29123 5 1 1 29122
0 29124 7 1 2 60159 77995
0 29125 5 1 1 29124
0 29126 7 1 2 73676 29125
0 29127 5 1 1 29126
0 29128 7 1 2 61554 29127
0 29129 7 1 2 29123 29128
0 29130 5 1 1 29129
0 29131 7 1 2 63036 29130
0 29132 7 1 2 29121 29131
0 29133 5 1 1 29132
0 29134 7 1 2 83501 78255
0 29135 5 1 1 29134
0 29136 7 1 2 63476 29135
0 29137 7 1 2 29133 29136
0 29138 7 1 2 29114 29137
0 29139 5 1 1 29138
0 29140 7 1 2 63754 29139
0 29141 7 1 2 29095 29140
0 29142 5 1 1 29141
0 29143 7 1 2 66295 92940
0 29144 5 1 1 29143
0 29145 7 1 2 60363 29144
0 29146 5 1 1 29145
0 29147 7 1 2 63037 29146
0 29148 5 1 1 29147
0 29149 7 1 2 72558 79540
0 29150 5 1 1 29149
0 29151 7 1 2 29148 29150
0 29152 5 1 1 29151
0 29153 7 1 2 62670 29152
0 29154 5 1 1 29153
0 29155 7 1 2 82733 94020
0 29156 5 2 1 29155
0 29157 7 1 2 29154 94050
0 29158 5 1 1 29157
0 29159 7 1 2 66038 29158
0 29160 5 1 1 29159
0 29161 7 1 2 77967 83831
0 29162 5 1 1 29161
0 29163 7 1 2 29160 29162
0 29164 5 1 1 29163
0 29165 7 1 2 64989 29164
0 29166 5 1 1 29165
0 29167 7 1 2 76211 24466
0 29168 5 1 1 29167
0 29169 7 1 2 86035 29168
0 29170 5 1 1 29169
0 29171 7 1 2 29166 29170
0 29172 5 1 1 29171
0 29173 7 1 2 84867 29172
0 29174 5 1 1 29173
0 29175 7 1 2 29142 29174
0 29176 5 1 1 29175
0 29177 7 1 2 87387 29176
0 29178 5 1 1 29177
0 29179 7 1 2 78956 85552
0 29180 5 1 1 29179
0 29181 7 1 2 92079 29180
0 29182 5 1 1 29181
0 29183 7 1 2 82930 29182
0 29184 5 1 1 29183
0 29185 7 1 2 82372 94031
0 29186 5 1 1 29185
0 29187 7 1 2 90682 93218
0 29188 5 1 1 29187
0 29189 7 1 2 63755 69828
0 29190 7 1 2 94027 29189
0 29191 7 1 2 29188 29190
0 29192 5 1 1 29191
0 29193 7 1 2 29186 29192
0 29194 5 1 1 29193
0 29195 7 1 2 68877 29194
0 29196 5 1 1 29195
0 29197 7 1 2 29184 29196
0 29198 5 1 1 29197
0 29199 7 1 2 66845 29198
0 29200 5 1 1 29199
0 29201 7 3 2 66039 75846
0 29202 5 1 1 94052
0 29203 7 1 2 76851 86371
0 29204 7 1 2 94053 29203
0 29205 5 1 1 29204
0 29206 7 1 2 29200 29205
0 29207 5 1 1 29206
0 29208 7 1 2 64760 29207
0 29209 5 1 1 29208
0 29210 7 1 2 79938 81643
0 29211 5 1 1 29210
0 29212 7 1 2 77784 78992
0 29213 5 1 1 29212
0 29214 7 1 2 29211 29213
0 29215 5 1 1 29214
0 29216 7 1 2 86367 29215
0 29217 5 1 1 29216
0 29218 7 1 2 29209 29217
0 29219 5 1 1 29218
0 29220 7 1 2 65571 29219
0 29221 5 1 1 29220
0 29222 7 1 2 93877 94054
0 29223 5 1 1 29222
0 29224 7 1 2 81644 83175
0 29225 5 1 1 29224
0 29226 7 1 2 29223 29225
0 29227 5 1 1 29226
0 29228 7 3 2 87114 87857
0 29229 7 1 2 29227 94055
0 29230 5 1 1 29229
0 29231 7 1 2 29221 29230
0 29232 5 1 1 29231
0 29233 7 1 2 62319 29232
0 29234 5 1 1 29233
0 29235 7 2 2 66296 92340
0 29236 7 1 2 87418 94058
0 29237 5 1 1 29236
0 29238 7 1 2 86582 87167
0 29239 7 1 2 93568 29238
0 29240 5 1 1 29239
0 29241 7 1 2 29237 29240
0 29242 5 1 1 29241
0 29243 7 1 2 86384 29242
0 29244 5 1 1 29243
0 29245 7 1 2 29234 29244
0 29246 5 1 1 29245
0 29247 7 1 2 71788 29246
0 29248 5 1 1 29247
0 29249 7 1 2 67646 77785
0 29250 5 2 1 29249
0 29251 7 1 2 89886 94060
0 29252 5 1 1 29251
0 29253 7 1 2 61349 72989
0 29254 7 1 2 29252 29253
0 29255 5 1 1 29254
0 29256 7 1 2 82613 86683
0 29257 5 1 1 29256
0 29258 7 1 2 89433 29257
0 29259 7 1 2 29255 29258
0 29260 5 1 1 29259
0 29261 7 1 2 85698 29260
0 29262 5 1 1 29261
0 29263 7 1 2 66523 86255
0 29264 7 1 2 84929 29263
0 29265 5 1 1 29264
0 29266 7 1 2 29262 29265
0 29267 5 1 1 29266
0 29268 7 1 2 65572 29267
0 29269 5 1 1 29268
0 29270 7 1 2 77432 79042
0 29271 7 1 2 93969 29270
0 29272 5 1 1 29271
0 29273 7 1 2 29269 29272
0 29274 5 1 1 29273
0 29275 7 1 2 63987 29274
0 29276 5 1 1 29275
0 29277 7 2 2 85519 93731
0 29278 7 1 2 86708 86875
0 29279 7 1 2 94062 29278
0 29280 5 1 1 29279
0 29281 7 1 2 29276 29280
0 29282 5 1 1 29281
0 29283 7 1 2 80484 29282
0 29284 5 1 1 29283
0 29285 7 2 2 82482 91592
0 29286 7 1 2 90785 94064
0 29287 5 1 1 29286
0 29288 7 1 2 89504 29287
0 29289 5 1 1 29288
0 29290 7 2 2 86709 89930
0 29291 7 1 2 29289 94066
0 29292 5 1 1 29291
0 29293 7 3 2 79043 87168
0 29294 7 1 2 66524 81699
0 29295 7 1 2 94068 29294
0 29296 5 1 1 29295
0 29297 7 1 2 29292 29296
0 29298 5 1 1 29297
0 29299 7 1 2 63038 29298
0 29300 5 1 1 29299
0 29301 7 1 2 76563 92891
0 29302 5 1 1 29301
0 29303 7 1 2 71223 89413
0 29304 5 1 1 29303
0 29305 7 1 2 29302 29304
0 29306 5 1 1 29305
0 29307 7 1 2 70186 29306
0 29308 5 1 1 29307
0 29309 7 1 2 75112 89786
0 29310 5 1 1 29309
0 29311 7 1 2 29308 29310
0 29312 5 1 1 29311
0 29313 7 1 2 85342 86710
0 29314 7 1 2 29312 29313
0 29315 5 1 1 29314
0 29316 7 1 2 29300 29315
0 29317 5 1 1 29316
0 29318 7 1 2 72121 29317
0 29319 5 1 1 29318
0 29320 7 1 2 88973 88839
0 29321 5 1 1 29320
0 29322 7 1 2 76783 29321
0 29323 5 1 1 29322
0 29324 7 1 2 78220 88587
0 29325 5 1 1 29324
0 29326 7 1 2 71557 29325
0 29327 7 1 2 29323 29326
0 29328 5 1 1 29327
0 29329 7 1 2 79870 88151
0 29330 7 1 2 29328 29329
0 29331 5 1 1 29330
0 29332 7 1 2 29319 29331
0 29333 5 1 1 29332
0 29334 7 1 2 63988 29333
0 29335 5 1 1 29334
0 29336 7 1 2 62671 74693
0 29337 5 1 1 29336
0 29338 7 1 2 17003 29337
0 29339 5 1 1 29338
0 29340 7 2 2 65573 83100
0 29341 7 1 2 85520 87992
0 29342 7 1 2 94071 29341
0 29343 7 1 2 29339 29342
0 29344 5 1 1 29343
0 29345 7 1 2 29335 29344
0 29346 5 1 1 29345
0 29347 7 1 2 73717 29346
0 29348 5 1 1 29347
0 29349 7 1 2 81653 84432
0 29350 5 1 1 29349
0 29351 7 1 2 84787 29350
0 29352 5 1 1 29351
0 29353 7 1 2 93699 29352
0 29354 5 1 1 29353
0 29355 7 1 2 63756 93693
0 29356 5 1 1 29355
0 29357 7 1 2 29354 29356
0 29358 5 1 1 29357
0 29359 7 1 2 69829 29358
0 29360 5 1 1 29359
0 29361 7 2 2 64523 76363
0 29362 5 2 1 94073
0 29363 7 1 2 72778 94075
0 29364 5 2 1 29363
0 29365 7 7 2 63989 84433
0 29366 7 1 2 86353 94079
0 29367 7 1 2 94077 29366
0 29368 5 1 1 29367
0 29369 7 1 2 29360 29368
0 29370 5 1 1 29369
0 29371 7 1 2 65574 29370
0 29372 5 1 1 29371
0 29373 7 1 2 79851 79970
0 29374 5 1 1 29373
0 29375 7 1 2 78256 94056
0 29376 7 1 2 29374 29375
0 29377 5 1 1 29376
0 29378 7 1 2 29372 29377
0 29379 5 1 1 29378
0 29380 7 1 2 63477 29379
0 29381 5 1 1 29380
0 29382 7 1 2 76364 87388
0 29383 5 1 1 29382
0 29384 7 2 2 65575 65716
0 29385 7 2 2 64282 94086
0 29386 7 1 2 86320 94088
0 29387 5 1 1 29386
0 29388 7 1 2 29383 29387
0 29389 5 1 1 29388
0 29390 7 1 2 84858 91904
0 29391 7 1 2 29389 29390
0 29392 5 1 1 29391
0 29393 7 1 2 29381 29392
0 29394 5 1 1 29393
0 29395 7 1 2 77195 29394
0 29396 5 1 1 29395
0 29397 7 3 2 78763 87389
0 29398 7 1 2 81858 79563
0 29399 7 1 2 94090 29398
0 29400 5 1 1 29399
0 29401 7 1 2 81978 86314
0 29402 7 1 2 86272 87410
0 29403 7 1 2 29401 29402
0 29404 5 1 1 29403
0 29405 7 1 2 69830 84868
0 29406 5 1 1 29405
0 29407 7 1 2 78789 29406
0 29408 5 1 1 29407
0 29409 7 1 2 66297 87390
0 29410 7 1 2 29408 29409
0 29411 5 1 1 29410
0 29412 7 1 2 29404 29411
0 29413 5 1 1 29412
0 29414 7 1 2 65221 73110
0 29415 7 1 2 29413 29414
0 29416 5 1 1 29415
0 29417 7 1 2 29400 29416
0 29418 5 1 1 29417
0 29419 7 1 2 89050 29418
0 29420 5 1 1 29419
0 29421 7 1 2 29396 29420
0 29422 7 1 2 29348 29421
0 29423 7 1 2 29284 29422
0 29424 7 1 2 29248 29423
0 29425 7 1 2 29178 29424
0 29426 7 1 2 29031 29425
0 29427 7 1 2 28838 29426
0 29428 7 1 2 28430 29427
0 29429 5 1 1 29428
0 29430 7 1 2 81181 29429
0 29431 5 1 1 29430
0 29432 7 3 2 65717 85777
0 29433 7 1 2 74959 87325
0 29434 7 1 2 94093 29433
0 29435 5 1 1 29434
0 29436 7 1 2 9096 29435
0 29437 5 1 1 29436
0 29438 7 1 2 66298 29437
0 29439 5 1 1 29438
0 29440 7 2 2 80169 80732
0 29441 5 1 1 94096
0 29442 7 1 2 81124 29441
0 29443 5 1 1 29442
0 29444 7 1 2 94074 29443
0 29445 5 1 1 29444
0 29446 7 1 2 69831 86417
0 29447 5 1 1 29446
0 29448 7 1 2 63478 86445
0 29449 5 1 1 29448
0 29450 7 1 2 29447 29449
0 29451 5 1 1 29450
0 29452 7 1 2 62111 29451
0 29453 5 1 1 29452
0 29454 7 1 2 29445 29453
0 29455 5 1 1 29454
0 29456 7 1 2 67647 29455
0 29457 5 1 1 29456
0 29458 7 1 2 29439 29457
0 29459 5 2 1 29458
0 29460 7 1 2 86084 94098
0 29461 5 1 1 29460
0 29462 7 1 2 81979 86971
0 29463 7 1 2 81660 29462
0 29464 5 1 1 29463
0 29465 7 1 2 29461 29464
0 29466 5 1 1 29465
0 29467 7 1 2 63757 29466
0 29468 5 1 1 29467
0 29469 7 5 2 61870 80997
0 29470 7 2 2 71010 94100
0 29471 7 1 2 72559 94105
0 29472 5 1 1 29471
0 29473 7 1 2 79888 81988
0 29474 7 1 2 93710 29473
0 29475 5 1 1 29474
0 29476 7 1 2 29472 29475
0 29477 5 1 1 29476
0 29478 7 1 2 73111 29477
0 29479 5 1 1 29478
0 29480 7 1 2 79889 82109
0 29481 7 1 2 93663 29480
0 29482 5 1 1 29481
0 29483 7 1 2 29479 29482
0 29484 5 1 1 29483
0 29485 7 1 2 87908 29484
0 29486 5 1 1 29485
0 29487 7 1 2 29468 29486
0 29488 5 1 1 29487
0 29489 7 1 2 68013 29488
0 29490 5 1 1 29489
0 29491 7 4 2 86256 86583
0 29492 7 1 2 75847 94107
0 29493 5 1 1 29492
0 29494 7 1 2 61555 92569
0 29495 7 1 2 82041 29494
0 29496 5 1 1 29495
0 29497 7 2 2 81027 85669
0 29498 5 1 1 94111
0 29499 7 1 2 29496 29498
0 29500 5 1 1 29499
0 29501 7 1 2 74453 29500
0 29502 5 1 1 29501
0 29503 7 1 2 29493 29502
0 29504 5 1 1 29503
0 29505 7 1 2 69832 29504
0 29506 5 1 1 29505
0 29507 7 1 2 85103 94112
0 29508 5 1 1 29507
0 29509 7 1 2 29506 29508
0 29510 5 1 1 29509
0 29511 7 1 2 93779 29510
0 29512 5 1 1 29511
0 29513 7 1 2 29490 29512
0 29514 5 1 1 29513
0 29515 7 1 2 65576 29514
0 29516 5 1 1 29515
0 29517 7 1 2 63758 94099
0 29518 5 1 1 29517
0 29519 7 1 2 73349 92641
0 29520 7 1 2 84641 29519
0 29521 7 1 2 81407 29520
0 29522 5 1 1 29521
0 29523 7 1 2 29518 29522
0 29524 5 1 1 29523
0 29525 7 1 2 68014 29524
0 29526 5 1 1 29525
0 29527 7 1 2 64283 90757
0 29528 5 1 1 29527
0 29529 7 1 2 8443 29528
0 29530 5 1 1 29529
0 29531 7 1 2 89949 93506
0 29532 7 1 2 29530 29531
0 29533 5 1 1 29532
0 29534 7 1 2 29526 29533
0 29535 5 1 1 29534
0 29536 7 1 2 87140 29535
0 29537 5 1 1 29536
0 29538 7 1 2 29516 29537
0 29539 5 1 1 29538
0 29540 7 1 2 93764 29539
0 29541 5 1 1 29540
0 29542 7 1 2 69833 26862
0 29543 5 1 1 29542
0 29544 7 1 2 76186 92909
0 29545 5 1 1 29544
0 29546 7 2 2 63039 77094
0 29547 5 2 1 94113
0 29548 7 1 2 76365 94114
0 29549 7 1 2 29545 29548
0 29550 5 1 1 29549
0 29551 7 1 2 74454 77402
0 29552 5 1 1 29551
0 29553 7 1 2 86566 93683
0 29554 5 1 1 29553
0 29555 7 1 2 64761 29554
0 29556 5 1 1 29555
0 29557 7 1 2 29552 29556
0 29558 7 1 2 29550 29557
0 29559 7 1 2 29543 29558
0 29560 5 1 1 29559
0 29561 7 1 2 83543 29560
0 29562 5 1 1 29561
0 29563 7 3 2 67648 78596
0 29564 5 1 1 94117
0 29565 7 1 2 81512 91552
0 29566 5 1 1 29565
0 29567 7 1 2 94118 29566
0 29568 5 1 1 29567
0 29569 7 1 2 69928 82964
0 29570 5 1 1 29569
0 29571 7 3 2 60806 82991
0 29572 5 1 1 94120
0 29573 7 1 2 29570 29572
0 29574 5 1 1 29573
0 29575 7 1 2 76000 29574
0 29576 5 1 1 29575
0 29577 7 1 2 79594 29576
0 29578 7 1 2 29568 29577
0 29579 5 1 1 29578
0 29580 7 1 2 78764 29579
0 29581 5 1 1 29580
0 29582 7 1 2 29562 29581
0 29583 5 1 1 29582
0 29584 7 1 2 66706 29583
0 29585 5 1 1 29584
0 29586 7 1 2 70055 92506
0 29587 5 1 1 29586
0 29588 7 1 2 29585 29587
0 29589 5 1 1 29588
0 29590 7 1 2 68878 29589
0 29591 5 1 1 29590
0 29592 7 1 2 91575 90049
0 29593 5 1 1 29592
0 29594 7 1 2 65430 29593
0 29595 7 1 2 29591 29594
0 29596 5 1 1 29595
0 29597 7 1 2 84159 85521
0 29598 5 1 1 29597
0 29599 7 1 2 92377 29598
0 29600 5 1 1 29599
0 29601 7 1 2 66299 29600
0 29602 5 1 1 29601
0 29603 7 1 2 22195 29602
0 29604 5 1 1 29603
0 29605 7 1 2 63479 29604
0 29606 5 1 1 29605
0 29607 7 1 2 84347 91576
0 29608 5 1 1 29607
0 29609 7 1 2 61729 94014
0 29610 5 1 1 29609
0 29611 7 1 2 29608 29610
0 29612 5 1 1 29611
0 29613 7 1 2 87538 29612
0 29614 5 1 1 29613
0 29615 7 1 2 60542 29614
0 29616 7 1 2 29606 29615
0 29617 5 1 1 29616
0 29618 7 1 2 65577 29617
0 29619 7 1 2 29596 29618
0 29620 5 1 1 29619
0 29621 7 1 2 87154 29620
0 29622 5 1 1 29621
0 29623 7 1 2 82950 85326
0 29624 5 1 1 29623
0 29625 7 1 2 7736 29624
0 29626 5 1 1 29625
0 29627 7 1 2 63480 29626
0 29628 5 1 1 29627
0 29629 7 1 2 79621 76677
0 29630 7 1 2 89705 29629
0 29631 5 1 1 29630
0 29632 7 1 2 29628 29631
0 29633 5 1 1 29632
0 29634 7 1 2 63990 29633
0 29635 5 1 1 29634
0 29636 7 1 2 86735 29635
0 29637 5 1 1 29636
0 29638 7 1 2 79332 29637
0 29639 7 1 2 29622 29638
0 29640 5 1 1 29639
0 29641 7 1 2 29541 29640
0 29642 7 1 2 29431 29641
0 29643 7 1 2 28144 29642
0 29644 7 1 2 27209 29643
0 29645 7 1 2 26678 29644
0 29646 7 1 2 25604 29645
0 29647 5 1 1 29646
0 29648 7 1 2 64090 29647
0 29649 5 1 1 29648
0 29650 7 2 2 12498 88296
0 29651 5 1 1 94123
0 29652 7 1 2 63481 29651
0 29653 5 1 1 29652
0 29654 7 1 2 80586 89218
0 29655 5 1 1 29654
0 29656 7 1 2 29653 29655
0 29657 5 1 1 29656
0 29658 7 1 2 61556 29657
0 29659 5 1 1 29658
0 29660 7 1 2 87675 88294
0 29661 5 1 1 29660
0 29662 7 1 2 29659 29661
0 29663 5 1 1 29662
0 29664 7 1 2 86158 29663
0 29665 5 1 1 29664
0 29666 7 1 2 64524 86085
0 29667 7 1 2 87672 29666
0 29668 5 1 1 29667
0 29669 7 1 2 29665 29668
0 29670 5 1 1 29669
0 29671 7 1 2 66707 29670
0 29672 5 1 1 29671
0 29673 7 1 2 87527 87269
0 29674 5 1 1 29673
0 29675 7 1 2 86834 87460
0 29676 5 1 1 29675
0 29677 7 1 2 88282 29676
0 29678 5 1 1 29677
0 29679 7 1 2 64990 86086
0 29680 7 1 2 29678 29679
0 29681 5 1 1 29680
0 29682 7 1 2 29674 29681
0 29683 5 1 1 29682
0 29684 7 1 2 81104 29683
0 29685 5 1 1 29684
0 29686 7 1 2 29672 29685
0 29687 5 1 1 29686
0 29688 7 1 2 65431 29687
0 29689 5 1 1 29688
0 29690 7 2 2 87067 87263
0 29691 7 1 2 75215 81081
0 29692 7 1 2 94125 29691
0 29693 5 1 1 29692
0 29694 7 4 2 64284 78570
0 29695 5 2 1 94127
0 29696 7 1 2 93197 94128
0 29697 5 1 1 29696
0 29698 7 1 2 11195 29697
0 29699 5 1 1 29698
0 29700 7 1 2 85845 29699
0 29701 5 1 1 29700
0 29702 7 1 2 87587 93654
0 29703 5 1 1 29702
0 29704 7 1 2 29701 29703
0 29705 5 1 1 29704
0 29706 7 1 2 64991 63991
0 29707 7 1 2 29705 29706
0 29708 5 1 1 29707
0 29709 7 1 2 29693 29708
0 29710 5 1 1 29709
0 29711 7 1 2 63482 29710
0 29712 5 1 1 29711
0 29713 7 1 2 29689 29712
0 29714 5 1 1 29713
0 29715 7 1 2 65578 29714
0 29716 5 1 1 29715
0 29717 7 2 2 79102 93406
0 29718 7 1 2 87461 94133
0 29719 5 1 1 29718
0 29720 7 1 2 80170 87445
0 29721 5 1 1 29720
0 29722 7 10 2 66525 80417
0 29723 5 1 1 94135
0 29724 7 1 2 3036 94131
0 29725 5 1 1 29724
0 29726 7 1 2 94136 29725
0 29727 5 1 1 29726
0 29728 7 1 2 29721 29727
0 29729 7 1 2 29719 29728
0 29730 5 1 1 29729
0 29731 7 1 2 84411 87141
0 29732 7 1 2 29730 29731
0 29733 5 1 1 29732
0 29734 7 1 2 29716 29733
0 29735 5 1 1 29734
0 29736 7 1 2 68695 29735
0 29737 5 1 1 29736
0 29738 7 2 2 80418 83461
0 29739 7 1 2 94091 94145
0 29740 5 1 1 29739
0 29741 7 1 2 29737 29740
0 29742 5 1 1 29741
0 29743 7 1 2 62672 29742
0 29744 5 1 1 29743
0 29745 7 1 2 79279 81196
0 29746 5 6 1 29745
0 29747 7 1 2 70801 70449
0 29748 7 1 2 92035 29747
0 29749 7 1 2 94069 29748
0 29750 7 1 2 94147 29749
0 29751 5 1 1 29750
0 29752 7 1 2 29744 29751
0 29753 5 1 1 29752
0 29754 7 1 2 62320 29753
0 29755 5 1 1 29754
0 29756 7 1 2 82352 87677
0 29757 5 1 1 29756
0 29758 7 1 2 65222 29757
0 29759 5 1 1 29758
0 29760 7 1 2 74659 86655
0 29761 5 1 1 29760
0 29762 7 1 2 29759 29761
0 29763 5 1 1 29762
0 29764 7 1 2 87637 29763
0 29765 5 1 1 29764
0 29766 7 2 2 86058 93609
0 29767 5 1 1 94153
0 29768 7 3 2 91853 92417
0 29769 5 7 1 94155
0 29770 7 5 2 80902 94156
0 29771 7 1 2 70056 94165
0 29772 5 1 1 29771
0 29773 7 3 2 75586 79622
0 29774 5 17 1 94170
0 29775 7 1 2 29772 94173
0 29776 5 2 1 29775
0 29777 7 1 2 86656 94190
0 29778 5 1 1 29777
0 29779 7 1 2 29767 29778
0 29780 5 1 1 29779
0 29781 7 1 2 86781 29780
0 29782 5 1 1 29781
0 29783 7 1 2 29765 29782
0 29784 5 1 1 29783
0 29785 7 1 2 63992 29784
0 29786 5 1 1 29785
0 29787 7 3 2 68879 87238
0 29788 7 1 2 87649 93243
0 29789 7 1 2 94192 29788
0 29790 5 1 1 29789
0 29791 7 1 2 29786 29790
0 29792 5 1 1 29791
0 29793 7 1 2 68696 29792
0 29794 5 1 1 29793
0 29795 7 3 2 68371 87169
0 29796 7 1 2 76743 80171
0 29797 7 4 2 68015 87858
0 29798 7 1 2 90427 94198
0 29799 7 1 2 29796 29798
0 29800 7 1 2 94195 29799
0 29801 5 1 1 29800
0 29802 7 1 2 29794 29801
0 29803 5 1 1 29802
0 29804 7 1 2 64285 29803
0 29805 5 1 1 29804
0 29806 7 1 2 78686 86618
0 29807 7 3 2 68016 88018
0 29808 7 1 2 92825 94202
0 29809 7 1 2 29806 29808
0 29810 5 1 1 29809
0 29811 7 1 2 29805 29810
0 29812 7 1 2 29755 29811
0 29813 5 1 1 29812
0 29814 7 1 2 64091 29813
0 29815 5 1 1 29814
0 29816 7 20 2 63759 68976
0 29817 7 7 2 79729 94205
0 29818 7 4 2 87068 94225
0 29819 7 3 2 79485 94232
0 29820 7 2 2 64286 80753
0 29821 7 3 2 65223 65579
0 29822 7 3 2 80513 94241
0 29823 7 1 2 94239 94244
0 29824 7 1 2 94236 29823
0 29825 5 1 1 29824
0 29826 7 1 2 29815 29825
0 29827 5 1 1 29826
0 29828 7 1 2 70367 29827
0 29829 5 1 1 29828
0 29830 7 1 2 86675 93285
0 29831 5 1 1 29830
0 29832 7 1 2 85760 87239
0 29833 5 1 1 29832
0 29834 7 1 2 29831 29833
0 29835 5 1 1 29834
0 29836 7 1 2 86159 29835
0 29837 5 1 1 29836
0 29838 7 2 2 80733 86546
0 29839 5 1 1 94247
0 29840 7 1 2 86087 94248
0 29841 5 1 1 29840
0 29842 7 1 2 29837 29841
0 29843 5 1 1 29842
0 29844 7 1 2 65876 29843
0 29845 5 1 1 29844
0 29846 7 10 2 66846 68017
0 29847 5 1 1 94249
0 29848 7 3 2 86141 94250
0 29849 5 1 1 94259
0 29850 7 1 2 80031 77668
0 29851 7 1 2 94260 29850
0 29852 5 1 1 29851
0 29853 7 1 2 29845 29852
0 29854 5 1 1 29853
0 29855 7 1 2 64525 29854
0 29856 5 1 1 29855
0 29857 7 2 2 62321 86687
0 29858 7 1 2 82899 87419
0 29859 7 1 2 94262 29858
0 29860 5 1 1 29859
0 29861 7 1 2 29856 29860
0 29862 5 1 1 29861
0 29863 7 1 2 68697 29862
0 29864 5 1 1 29863
0 29865 7 2 2 77968 85670
0 29866 7 1 2 85868 94264
0 29867 5 1 1 29866
0 29868 7 1 2 29864 29867
0 29869 5 1 1 29868
0 29870 7 1 2 62673 29869
0 29871 5 1 1 29870
0 29872 7 1 2 82536 93540
0 29873 5 1 1 29872
0 29874 7 1 2 70802 89965
0 29875 5 1 1 29874
0 29876 7 1 2 29873 29875
0 29877 5 1 1 29876
0 29878 7 1 2 61557 29877
0 29879 5 1 1 29878
0 29880 7 1 2 78807 92593
0 29881 5 1 1 29880
0 29882 7 1 2 29879 29881
0 29883 5 1 1 29882
0 29884 7 1 2 81786 94251
0 29885 7 1 2 29883 29884
0 29886 5 1 1 29885
0 29887 7 1 2 29871 29886
0 29888 5 1 1 29887
0 29889 7 1 2 69659 29888
0 29890 5 1 1 29889
0 29891 7 2 2 62322 72867
0 29892 5 2 1 94266
0 29893 7 1 2 64526 78307
0 29894 5 2 1 29893
0 29895 7 1 2 94268 94270
0 29896 5 6 1 29895
0 29897 7 3 2 67649 75587
0 29898 5 1 1 94278
0 29899 7 1 2 94272 94279
0 29900 5 1 1 29899
0 29901 7 1 2 16422 29900
0 29902 5 1 1 29901
0 29903 7 3 2 68018 29902
0 29904 5 1 1 94281
0 29905 7 5 2 68019 73741
0 29906 7 1 2 94284 94273
0 29907 5 1 1 29906
0 29908 7 1 2 81051 93289
0 29909 5 1 1 29908
0 29910 7 2 2 65718 70948
0 29911 5 1 1 94289
0 29912 7 1 2 84948 94290
0 29913 5 1 1 29912
0 29914 7 1 2 29909 29913
0 29915 7 1 2 29907 29914
0 29916 5 1 1 29915
0 29917 7 1 2 64992 29916
0 29918 5 1 1 29917
0 29919 7 1 2 29904 29918
0 29920 5 1 1 29919
0 29921 7 1 2 63483 29920
0 29922 5 1 1 29921
0 29923 7 1 2 79852 82312
0 29924 5 2 1 29923
0 29925 7 1 2 75588 94291
0 29926 5 1 1 29925
0 29927 7 1 2 76219 94240
0 29928 5 1 1 29927
0 29929 7 1 2 29926 29928
0 29930 5 1 1 29929
0 29931 7 2 2 81634 77786
0 29932 7 1 2 29930 94293
0 29933 5 1 1 29932
0 29934 7 1 2 29922 29933
0 29935 5 1 1 29934
0 29936 7 1 2 86088 29935
0 29937 5 1 1 29936
0 29938 7 1 2 84763 93907
0 29939 5 1 1 29938
0 29940 7 3 2 81052 78707
0 29941 5 2 1 94295
0 29942 7 1 2 82424 94298
0 29943 5 2 1 29942
0 29944 7 1 2 65877 94300
0 29945 5 1 1 29944
0 29946 7 1 2 63040 77281
0 29947 5 1 1 29946
0 29948 7 1 2 64527 84840
0 29949 7 1 2 29947 29948
0 29950 5 1 1 29949
0 29951 7 1 2 29945 29950
0 29952 5 1 1 29951
0 29953 7 1 2 62112 29952
0 29954 5 1 1 29953
0 29955 7 1 2 78871 91322
0 29956 5 1 1 29955
0 29957 7 1 2 29954 29956
0 29958 5 1 1 29957
0 29959 7 1 2 65224 29958
0 29960 5 1 1 29959
0 29961 7 1 2 29939 29960
0 29962 5 1 1 29961
0 29963 7 1 2 70803 29962
0 29964 5 1 1 29963
0 29965 7 2 2 87233 88300
0 29966 7 1 2 70450 94302
0 29967 5 1 1 29966
0 29968 7 1 2 79486 78835
0 29969 5 1 1 29968
0 29970 7 1 2 29967 29969
0 29971 5 1 1 29970
0 29972 7 1 2 76220 29971
0 29973 5 1 1 29972
0 29974 7 1 2 29964 29973
0 29975 5 1 1 29974
0 29976 7 1 2 65719 29975
0 29977 5 1 1 29976
0 29978 7 2 2 67329 75589
0 29979 7 1 2 93388 94304
0 29980 5 1 1 29979
0 29981 7 1 2 90398 94274
0 29982 5 1 1 29981
0 29983 7 1 2 29980 29982
0 29984 5 1 1 29983
0 29985 7 1 2 63041 29984
0 29986 5 1 1 29985
0 29987 7 1 2 68372 29986
0 29988 7 1 2 29977 29987
0 29989 5 1 1 29988
0 29990 7 1 2 75923 90030
0 29991 5 1 1 29990
0 29992 7 1 2 61558 94124
0 29993 5 1 1 29992
0 29994 7 1 2 62323 74920
0 29995 7 1 2 91789 29994
0 29996 7 1 2 29993 29995
0 29997 5 1 1 29996
0 29998 7 1 2 29991 29997
0 29999 5 1 1 29998
0 30000 7 1 2 64528 29999
0 30001 5 1 1 30000
0 30002 7 1 2 78914 90096
0 30003 5 1 1 30002
0 30004 7 1 2 61559 78716
0 30005 7 1 2 30003 30004
0 30006 5 1 1 30005
0 30007 7 1 2 82429 30006
0 30008 5 1 1 30007
0 30009 7 1 2 80605 30008
0 30010 5 1 1 30009
0 30011 7 1 2 68020 78950
0 30012 5 1 1 30011
0 30013 7 1 2 89539 30012
0 30014 5 1 1 30013
0 30015 7 1 2 60364 30014
0 30016 5 1 1 30015
0 30017 7 1 2 83904 78687
0 30018 5 1 1 30017
0 30019 7 1 2 30016 30018
0 30020 5 1 1 30019
0 30021 7 1 2 82306 30020
0 30022 5 1 1 30021
0 30023 7 1 2 71789 79055
0 30024 7 1 2 85040 30023
0 30025 5 1 1 30024
0 30026 7 1 2 62113 30025
0 30027 7 1 2 30022 30026
0 30028 7 1 2 30010 30027
0 30029 5 1 1 30028
0 30030 7 1 2 70187 17820
0 30031 5 1 1 30030
0 30032 7 1 2 83905 30031
0 30033 5 1 1 30032
0 30034 7 2 2 74346 79572
0 30035 5 1 1 94306
0 30036 7 1 2 67078 30035
0 30037 7 1 2 30033 30036
0 30038 5 1 1 30037
0 30039 7 1 2 30029 30038
0 30040 5 1 1 30039
0 30041 7 1 2 30001 30040
0 30042 5 1 1 30041
0 30043 7 1 2 62674 30042
0 30044 5 1 1 30043
0 30045 7 1 2 74023 94307
0 30046 5 1 1 30045
0 30047 7 2 2 73268 91390
0 30048 5 1 1 94308
0 30049 7 1 2 61560 94309
0 30050 5 1 1 30049
0 30051 7 1 2 71725 83602
0 30052 5 4 1 30051
0 30053 7 1 2 79309 78814
0 30054 5 1 1 30053
0 30055 7 1 2 94310 30054
0 30056 5 1 1 30055
0 30057 7 1 2 30050 30056
0 30058 5 1 1 30057
0 30059 7 1 2 63042 30058
0 30060 5 1 1 30059
0 30061 7 1 2 30046 30060
0 30062 5 1 1 30061
0 30063 7 1 2 67650 30062
0 30064 5 1 1 30063
0 30065 7 1 2 63484 30064
0 30066 7 1 2 30044 30065
0 30067 5 1 1 30066
0 30068 7 1 2 86160 30067
0 30069 7 1 2 29989 30068
0 30070 5 1 1 30069
0 30071 7 1 2 29937 30070
0 30072 5 1 1 30071
0 30073 7 1 2 68698 30072
0 30074 5 1 1 30073
0 30075 7 1 2 75742 83038
0 30076 5 1 1 30075
0 30077 7 1 2 82837 30076
0 30078 5 1 1 30077
0 30079 7 2 2 80980 86239
0 30080 7 1 2 30078 94314
0 30081 5 1 1 30080
0 30082 7 2 2 82614 82627
0 30083 5 1 1 94316
0 30084 7 1 2 94311 94317
0 30085 5 1 1 30084
0 30086 7 1 2 83101 86899
0 30087 7 5 2 68880 70804
0 30088 7 1 2 91293 94318
0 30089 7 1 2 30086 30088
0 30090 5 1 1 30089
0 30091 7 1 2 30085 30090
0 30092 5 1 1 30091
0 30093 7 1 2 61871 30092
0 30094 5 1 1 30093
0 30095 7 1 2 30081 30094
0 30096 5 1 1 30095
0 30097 7 1 2 63760 30096
0 30098 5 1 1 30097
0 30099 7 1 2 65432 30098
0 30100 7 1 2 30074 30099
0 30101 7 1 2 29890 30100
0 30102 5 1 1 30101
0 30103 7 1 2 81058 91079
0 30104 5 1 1 30103
0 30105 7 1 2 71558 30104
0 30106 5 1 1 30105
0 30107 7 1 2 86665 91070
0 30108 5 1 1 30107
0 30109 7 2 2 70805 83906
0 30110 5 1 1 94323
0 30111 7 1 2 30108 30110
0 30112 5 1 1 30111
0 30113 7 1 2 71990 30112
0 30114 5 1 1 30113
0 30115 7 1 2 93481 30114
0 30116 7 1 2 30106 30115
0 30117 5 1 1 30116
0 30118 7 1 2 65720 30117
0 30119 5 1 1 30118
0 30120 7 1 2 63043 81137
0 30121 5 1 1 30120
0 30122 7 1 2 30119 30121
0 30123 5 1 1 30122
0 30124 7 1 2 64287 30123
0 30125 5 1 1 30124
0 30126 7 1 2 75888 90966
0 30127 5 1 1 30126
0 30128 7 1 2 66300 15350
0 30129 7 1 2 30127 30128
0 30130 5 1 1 30129
0 30131 7 1 2 79487 71381
0 30132 5 1 1 30131
0 30133 7 1 2 30130 30132
0 30134 7 1 2 30125 30133
0 30135 5 1 1 30134
0 30136 7 1 2 86161 30135
0 30137 5 1 1 30136
0 30138 7 1 2 75096 89065
0 30139 5 1 1 30138
0 30140 7 1 2 83229 30139
0 30141 5 1 1 30140
0 30142 7 1 2 74024 30141
0 30143 5 1 1 30142
0 30144 7 1 2 67330 69368
0 30145 5 1 1 30144
0 30146 7 1 2 2923 30145
0 30147 5 3 1 30146
0 30148 7 1 2 64288 94325
0 30149 5 1 1 30148
0 30150 7 1 2 72837 89602
0 30151 5 1 1 30150
0 30152 7 1 2 70536 30151
0 30153 5 1 1 30152
0 30154 7 1 2 30149 30153
0 30155 5 1 1 30154
0 30156 7 1 2 62675 30155
0 30157 5 1 1 30156
0 30158 7 1 2 30143 30157
0 30159 5 2 1 30158
0 30160 7 1 2 70806 94328
0 30161 5 1 1 30160
0 30162 7 1 2 67651 80275
0 30163 5 1 1 30162
0 30164 7 1 2 30161 30163
0 30165 5 1 1 30164
0 30166 7 1 2 68021 30165
0 30167 5 1 1 30166
0 30168 7 1 2 77353 84949
0 30169 5 1 1 30168
0 30170 7 1 2 30167 30169
0 30171 5 1 1 30170
0 30172 7 1 2 86089 30171
0 30173 5 1 1 30172
0 30174 7 1 2 30137 30173
0 30175 5 2 1 30174
0 30176 7 1 2 63485 94330
0 30177 5 1 1 30176
0 30178 7 1 2 86162 93094
0 30179 5 1 1 30178
0 30180 7 1 2 87049 30179
0 30181 5 1 1 30180
0 30182 7 1 2 66526 30181
0 30183 5 1 1 30182
0 30184 7 5 2 63044 71559
0 30185 7 1 2 71991 94332
0 30186 5 1 1 30185
0 30187 7 1 2 26041 30186
0 30188 5 1 1 30187
0 30189 7 1 2 86090 30188
0 30190 5 1 1 30189
0 30191 7 1 2 30183 30190
0 30192 5 1 1 30191
0 30193 7 1 2 69660 30192
0 30194 5 1 1 30193
0 30195 7 1 2 85062 93706
0 30196 5 1 1 30195
0 30197 7 1 2 66847 94193
0 30198 5 1 1 30197
0 30199 7 1 2 30196 30198
0 30200 5 1 1 30199
0 30201 7 1 2 62676 30200
0 30202 5 1 1 30201
0 30203 7 1 2 30194 30202
0 30204 5 1 1 30203
0 30205 7 1 2 62114 30204
0 30206 5 1 1 30205
0 30207 7 1 2 87052 88548
0 30208 5 1 1 30207
0 30209 7 1 2 30206 30208
0 30210 5 1 1 30209
0 30211 7 1 2 80734 30210
0 30212 5 1 1 30211
0 30213 7 1 2 30177 30212
0 30214 5 1 1 30213
0 30215 7 1 2 63761 30214
0 30216 5 1 1 30215
0 30217 7 2 2 85909 88013
0 30218 7 1 2 66848 94337
0 30219 5 1 1 30218
0 30220 7 1 2 70451 78571
0 30221 5 1 1 30220
0 30222 7 1 2 65225 72785
0 30223 5 1 1 30222
0 30224 7 1 2 30221 30223
0 30225 5 1 1 30224
0 30226 7 1 2 62324 30225
0 30227 5 1 1 30226
0 30228 7 1 2 80606 85565
0 30229 5 1 1 30228
0 30230 7 1 2 65226 93290
0 30231 5 2 1 30230
0 30232 7 1 2 30229 94339
0 30233 7 1 2 30227 30232
0 30234 5 2 1 30233
0 30235 7 1 2 75688 85671
0 30236 7 1 2 94341 30235
0 30237 5 1 1 30236
0 30238 7 1 2 30219 30237
0 30239 5 1 1 30238
0 30240 7 1 2 64993 30239
0 30241 5 1 1 30240
0 30242 7 1 2 64529 94326
0 30243 5 1 1 30242
0 30244 7 1 2 65721 69252
0 30245 7 1 2 74306 30244
0 30246 5 1 1 30245
0 30247 7 1 2 30243 30246
0 30248 5 1 1 30247
0 30249 7 1 2 64289 30248
0 30250 5 1 1 30249
0 30251 7 1 2 1482 76068
0 30252 5 1 1 30251
0 30253 7 1 2 70537 30252
0 30254 5 1 1 30253
0 30255 7 1 2 67652 30254
0 30256 7 1 2 30250 30255
0 30257 5 1 1 30256
0 30258 7 12 2 66849 68373
0 30259 5 2 1 94343
0 30260 7 2 2 84828 94344
0 30261 7 1 2 73177 94357
0 30262 7 1 2 30257 30261
0 30263 5 1 1 30262
0 30264 7 1 2 30241 30263
0 30265 5 1 1 30264
0 30266 7 1 2 63993 30265
0 30267 5 1 1 30266
0 30268 7 3 2 68881 72594
0 30269 7 1 2 66850 80599
0 30270 7 2 2 94359 30269
0 30271 7 1 2 86856 87577
0 30272 7 1 2 94362 30271
0 30273 5 1 1 30272
0 30274 7 1 2 30267 30273
0 30275 5 1 1 30274
0 30276 7 1 2 68699 30275
0 30277 5 1 1 30276
0 30278 7 1 2 60543 30277
0 30279 7 1 2 30216 30278
0 30280 5 1 1 30279
0 30281 7 1 2 30102 30280
0 30282 5 1 1 30281
0 30283 7 1 2 75907 86514
0 30284 7 1 2 87986 30283
0 30285 5 1 1 30284
0 30286 7 1 2 5412 30285
0 30287 5 1 1 30286
0 30288 7 1 2 64290 30287
0 30289 5 1 1 30288
0 30290 7 1 2 74408 8476
0 30291 5 1 1 30290
0 30292 7 1 2 70057 30291
0 30293 5 1 1 30292
0 30294 7 1 2 30289 30293
0 30295 5 1 1 30294
0 30296 7 1 2 91945 30295
0 30297 5 1 1 30296
0 30298 7 2 2 74737 83544
0 30299 7 1 2 70058 94364
0 30300 7 1 2 94275 30299
0 30301 5 1 1 30300
0 30302 7 1 2 30297 30301
0 30303 5 1 1 30302
0 30304 7 1 2 68022 30303
0 30305 5 1 1 30304
0 30306 7 1 2 86427 90300
0 30307 5 1 1 30306
0 30308 7 1 2 65722 84987
0 30309 5 1 1 30308
0 30310 7 1 2 79943 30309
0 30311 5 1 1 30310
0 30312 7 1 2 65878 30311
0 30313 5 1 1 30312
0 30314 7 1 2 30307 30313
0 30315 5 1 1 30314
0 30316 7 1 2 64530 30315
0 30317 5 1 1 30316
0 30318 7 1 2 79939 75924
0 30319 5 1 1 30318
0 30320 7 1 2 30317 30319
0 30321 5 1 1 30320
0 30322 7 1 2 84778 86547
0 30323 7 1 2 30321 30322
0 30324 5 1 1 30323
0 30325 7 1 2 30305 30324
0 30326 5 1 1 30325
0 30327 7 1 2 87455 30326
0 30328 5 1 1 30327
0 30329 7 1 2 66708 30328
0 30330 7 1 2 30282 30329
0 30331 5 1 1 30330
0 30332 7 1 2 65433 94331
0 30333 5 1 1 30332
0 30334 7 1 2 87276 94329
0 30335 5 1 1 30334
0 30336 7 2 2 68882 87207
0 30337 7 1 2 86948 86933
0 30338 7 1 2 94366 30337
0 30339 5 1 1 30338
0 30340 7 1 2 30335 30339
0 30341 5 1 1 30340
0 30342 7 1 2 70807 30341
0 30343 5 1 1 30342
0 30344 7 1 2 88165 91080
0 30345 5 1 1 30344
0 30346 7 1 2 69834 86163
0 30347 7 1 2 30345 30346
0 30348 5 1 1 30347
0 30349 7 1 2 27946 30348
0 30350 5 1 1 30349
0 30351 7 1 2 66301 30350
0 30352 5 1 1 30351
0 30353 7 1 2 90630 94108
0 30354 5 1 1 30353
0 30355 7 1 2 30352 30354
0 30356 5 1 1 30355
0 30357 7 1 2 64994 30356
0 30358 5 1 1 30357
0 30359 7 2 2 69661 86164
0 30360 7 1 2 81082 77474
0 30361 7 1 2 94368 30360
0 30362 5 1 1 30361
0 30363 7 1 2 30358 30362
0 30364 7 1 2 30343 30363
0 30365 5 1 1 30364
0 30366 7 1 2 75216 30365
0 30367 5 1 1 30366
0 30368 7 1 2 63762 30367
0 30369 7 1 2 30333 30368
0 30370 5 1 1 30369
0 30371 7 1 2 70538 70459
0 30372 5 2 1 30371
0 30373 7 1 2 75908 94370
0 30374 5 1 1 30373
0 30375 7 1 2 61350 30374
0 30376 5 1 1 30375
0 30377 7 2 2 81771 85672
0 30378 5 2 1 94372
0 30379 7 1 2 61561 87208
0 30380 5 1 1 30379
0 30381 7 1 2 94374 30380
0 30382 5 1 1 30381
0 30383 7 1 2 30376 30382
0 30384 5 1 1 30383
0 30385 7 1 2 64531 70406
0 30386 5 1 1 30385
0 30387 7 1 2 72792 30386
0 30388 5 1 1 30387
0 30389 7 1 2 64291 30388
0 30390 5 1 1 30389
0 30391 7 1 2 78898 30390
0 30392 5 2 1 30391
0 30393 7 2 2 65434 93974
0 30394 5 1 1 94378
0 30395 7 1 2 83467 94379
0 30396 7 1 2 94376 30395
0 30397 5 1 1 30396
0 30398 7 1 2 30384 30397
0 30399 5 1 1 30398
0 30400 7 1 2 62677 30399
0 30401 5 1 1 30400
0 30402 7 1 2 81083 88060
0 30403 7 1 2 94276 30402
0 30404 5 1 1 30403
0 30405 7 1 2 30401 30404
0 30406 5 1 1 30405
0 30407 7 1 2 64995 30406
0 30408 5 1 1 30407
0 30409 7 1 2 87209 94282
0 30410 5 1 1 30409
0 30411 7 1 2 30408 30410
0 30412 5 1 1 30411
0 30413 7 1 2 63994 30412
0 30414 5 1 1 30413
0 30415 7 2 2 66527 80514
0 30416 7 1 2 81974 94380
0 30417 7 1 2 94363 30416
0 30418 5 1 1 30417
0 30419 7 1 2 68700 30418
0 30420 7 1 2 30414 30419
0 30421 5 1 1 30420
0 30422 7 1 2 30370 30421
0 30423 5 1 1 30422
0 30424 7 1 2 63486 30423
0 30425 5 1 1 30424
0 30426 7 2 2 61872 88233
0 30427 7 1 2 91854 94382
0 30428 5 1 1 30427
0 30429 7 1 2 85699 87588
0 30430 7 1 2 76830 30429
0 30431 5 1 1 30430
0 30432 7 1 2 30428 30431
0 30433 5 1 1 30432
0 30434 7 1 2 77354 30433
0 30435 5 1 1 30434
0 30436 7 2 2 65723 68701
0 30437 7 1 2 87210 94384
0 30438 7 1 2 93821 30437
0 30439 5 1 1 30438
0 30440 7 1 2 30435 30439
0 30441 5 1 1 30440
0 30442 7 1 2 63045 30441
0 30443 5 1 1 30442
0 30444 7 2 2 84829 85700
0 30445 7 2 2 78840 74250
0 30446 7 1 2 94386 94388
0 30447 7 1 2 80607 30446
0 30448 5 1 1 30447
0 30449 7 1 2 30443 30448
0 30450 5 1 1 30449
0 30451 7 1 2 66302 30450
0 30452 5 1 1 30451
0 30453 7 1 2 79103 93428
0 30454 5 1 1 30453
0 30455 7 1 2 64292 83700
0 30456 7 1 2 91071 30455
0 30457 5 1 1 30456
0 30458 7 1 2 30454 30457
0 30459 5 1 1 30458
0 30460 7 1 2 82066 30459
0 30461 5 1 1 30460
0 30462 7 3 2 64532 84634
0 30463 7 3 2 82615 78375
0 30464 7 1 2 94390 94393
0 30465 5 1 1 30464
0 30466 7 1 2 30461 30465
0 30467 5 1 1 30466
0 30468 7 1 2 85701 30467
0 30469 5 1 1 30468
0 30470 7 1 2 30452 30469
0 30471 5 1 1 30470
0 30472 7 1 2 62115 30471
0 30473 5 1 1 30472
0 30474 7 1 2 84082 91210
0 30475 5 1 1 30474
0 30476 7 1 2 93595 30475
0 30477 5 1 1 30476
0 30478 7 1 2 86432 30477
0 30479 5 1 1 30478
0 30480 7 1 2 85138 94312
0 30481 5 1 1 30480
0 30482 7 1 2 30479 30481
0 30483 5 1 1 30482
0 30484 7 1 2 67653 30483
0 30485 5 1 1 30484
0 30486 7 1 2 61351 93889
0 30487 5 1 1 30486
0 30488 7 1 2 30485 30487
0 30489 5 1 1 30488
0 30490 7 1 2 84830 30489
0 30491 5 1 1 30490
0 30492 7 1 2 78033 79232
0 30493 7 1 2 93554 30492
0 30494 5 1 1 30493
0 30495 7 1 2 30491 30494
0 30496 5 1 1 30495
0 30497 7 1 2 66851 30496
0 30498 5 1 1 30497
0 30499 7 1 2 30473 30498
0 30500 5 1 1 30499
0 30501 7 1 2 63995 30500
0 30502 5 1 1 30501
0 30503 7 2 2 66852 92957
0 30504 7 1 2 88014 94396
0 30505 5 1 1 30504
0 30506 7 1 2 66528 79710
0 30507 7 1 2 87610 30506
0 30508 5 1 1 30507
0 30509 7 1 2 30505 30508
0 30510 5 1 1 30509
0 30511 7 1 2 65227 30510
0 30512 5 1 1 30511
0 30513 7 1 2 78708 93902
0 30514 5 1 1 30513
0 30515 7 1 2 30512 30514
0 30516 5 1 1 30515
0 30517 7 1 2 70059 30516
0 30518 5 1 1 30517
0 30519 7 1 2 88007 94387
0 30520 5 1 1 30519
0 30521 7 1 2 30518 30520
0 30522 5 1 1 30521
0 30523 7 1 2 71992 30522
0 30524 5 1 1 30523
0 30525 7 1 2 76187 86502
0 30526 7 1 2 88234 30525
0 30527 7 1 2 91654 30526
0 30528 5 1 1 30527
0 30529 7 1 2 30524 30528
0 30530 5 1 1 30529
0 30531 7 1 2 63996 30530
0 30532 5 1 1 30531
0 30533 7 1 2 70492 93626
0 30534 7 1 2 93835 30533
0 30535 5 1 1 30534
0 30536 7 1 2 30532 30535
0 30537 5 1 1 30536
0 30538 7 1 2 69662 30537
0 30539 5 1 1 30538
0 30540 7 1 2 65435 86570
0 30541 7 1 2 84112 30540
0 30542 7 1 2 94194 30541
0 30543 5 1 1 30542
0 30544 7 1 2 68374 30543
0 30545 7 1 2 30539 30544
0 30546 7 1 2 30502 30545
0 30547 5 1 1 30546
0 30548 7 1 2 30425 30547
0 30549 5 1 1 30548
0 30550 7 1 2 61730 30549
0 30551 5 1 1 30550
0 30552 7 1 2 30331 30551
0 30553 5 1 1 30552
0 30554 7 3 2 69663 81422
0 30555 5 1 1 94398
0 30556 7 1 2 84920 94399
0 30557 5 1 1 30556
0 30558 7 1 2 82353 30557
0 30559 5 1 1 30558
0 30560 7 1 2 65879 30559
0 30561 5 1 1 30560
0 30562 7 1 2 83605 86657
0 30563 5 1 1 30562
0 30564 7 1 2 30561 30563
0 30565 5 1 1 30564
0 30566 7 1 2 64533 30565
0 30567 5 1 1 30566
0 30568 7 1 2 82345 94267
0 30569 5 1 1 30568
0 30570 7 1 2 30567 30569
0 30571 5 1 1 30570
0 30572 7 2 2 81277 89775
0 30573 5 1 1 94401
0 30574 7 1 2 86091 94402
0 30575 7 1 2 30571 30574
0 30576 5 1 1 30575
0 30577 7 1 2 65580 30576
0 30578 7 1 2 30553 30577
0 30579 5 1 1 30578
0 30580 7 8 2 63487 79649
0 30581 7 2 2 89457 94403
0 30582 7 2 2 74025 94411
0 30583 5 1 1 94413
0 30584 7 1 2 79404 94097
0 30585 5 1 1 30584
0 30586 7 1 2 30583 30585
0 30587 5 1 1 30586
0 30588 7 1 2 67654 30587
0 30589 5 1 1 30588
0 30590 7 2 2 75143 89850
0 30591 5 1 1 94415
0 30592 7 1 2 66709 94416
0 30593 5 1 1 30592
0 30594 7 1 2 30589 30593
0 30595 5 1 1 30594
0 30596 7 1 2 69835 30595
0 30597 5 1 1 30596
0 30598 7 1 2 74960 94148
0 30599 5 1 1 30598
0 30600 7 1 2 30597 30599
0 30601 5 1 1 30600
0 30602 7 1 2 62116 30601
0 30603 5 1 1 30602
0 30604 7 1 2 75097 94414
0 30605 5 1 1 30604
0 30606 7 1 2 30603 30605
0 30607 5 1 1 30606
0 30608 7 1 2 65880 30607
0 30609 5 1 1 30608
0 30610 7 1 2 89514 93444
0 30611 7 1 2 94412 30610
0 30612 5 1 1 30611
0 30613 7 1 2 30609 30612
0 30614 5 1 1 30613
0 30615 7 1 2 73481 30614
0 30616 5 1 1 30615
0 30617 7 3 2 65436 65724
0 30618 7 3 2 65228 94417
0 30619 7 2 2 70452 94420
0 30620 7 1 2 86639 92533
0 30621 7 1 2 94423 30620
0 30622 5 1 1 30621
0 30623 7 1 2 30616 30622
0 30624 5 1 1 30623
0 30625 7 1 2 70808 30624
0 30626 5 1 1 30625
0 30627 7 1 2 93766 94313
0 30628 5 1 1 30627
0 30629 7 1 2 81125 30628
0 30630 5 1 1 30629
0 30631 7 1 2 91211 30630
0 30632 5 1 1 30631
0 30633 7 1 2 71560 81182
0 30634 5 1 1 30633
0 30635 7 1 2 92383 30634
0 30636 5 1 1 30635
0 30637 7 1 2 63488 30636
0 30638 5 1 1 30637
0 30639 7 1 2 30632 30638
0 30640 5 1 1 30639
0 30641 7 1 2 67655 30640
0 30642 5 1 1 30641
0 30643 7 1 2 84160 75766
0 30644 7 1 2 91973 30643
0 30645 5 1 1 30644
0 30646 7 1 2 30642 30645
0 30647 5 1 1 30646
0 30648 7 1 2 68023 30647
0 30649 5 1 1 30648
0 30650 7 1 2 85970 90621
0 30651 5 2 1 30650
0 30652 7 1 2 79342 94425
0 30653 5 1 1 30652
0 30654 7 1 2 79814 85971
0 30655 5 2 1 30654
0 30656 7 1 2 81183 94427
0 30657 5 1 1 30656
0 30658 7 1 2 30653 30657
0 30659 5 1 1 30658
0 30660 7 1 2 62117 30659
0 30661 5 1 1 30660
0 30662 7 1 2 68375 80357
0 30663 7 1 2 79405 30662
0 30664 5 1 1 30663
0 30665 7 1 2 30661 30664
0 30666 5 1 1 30665
0 30667 7 1 2 62678 85242
0 30668 7 1 2 30666 30667
0 30669 5 1 1 30668
0 30670 7 1 2 30649 30669
0 30671 5 1 1 30670
0 30672 7 1 2 63997 30671
0 30673 5 1 1 30672
0 30674 7 1 2 30626 30673
0 30675 5 1 1 30674
0 30676 7 1 2 63763 30675
0 30677 5 1 1 30676
0 30678 7 1 2 94134 94377
0 30679 5 1 1 30678
0 30680 7 1 2 87599 30679
0 30681 5 1 1 30680
0 30682 7 1 2 66303 30681
0 30683 5 1 1 30682
0 30684 7 1 2 94137 94342
0 30685 5 1 1 30684
0 30686 7 2 2 65725 86415
0 30687 7 1 2 79623 94371
0 30688 7 1 2 94429 30687
0 30689 5 1 1 30688
0 30690 7 1 2 30685 30689
0 30691 7 1 2 30683 30690
0 30692 5 1 1 30691
0 30693 7 1 2 62679 30692
0 30694 5 1 1 30693
0 30695 7 3 2 94166 94285
0 30696 5 1 1 94431
0 30697 7 1 2 94432 94277
0 30698 5 1 1 30697
0 30699 7 1 2 30694 30698
0 30700 5 1 1 30699
0 30701 7 1 2 64996 30700
0 30702 5 1 1 30701
0 30703 7 1 2 79624 94283
0 30704 5 1 1 30703
0 30705 7 1 2 30702 30704
0 30706 5 1 1 30705
0 30707 7 1 2 63489 30706
0 30708 5 1 1 30707
0 30709 7 4 2 66710 75590
0 30710 5 7 1 94434
0 30711 7 1 2 94292 94435
0 30712 5 1 1 30711
0 30713 7 1 2 79845 80652
0 30714 7 1 2 84907 92418
0 30715 7 1 2 30713 30714
0 30716 5 1 1 30715
0 30717 7 1 2 30712 30716
0 30718 5 1 1 30717
0 30719 7 1 2 65437 30718
0 30720 5 1 1 30719
0 30721 7 1 2 84628 86900
0 30722 7 1 2 87658 30721
0 30723 5 1 1 30722
0 30724 7 1 2 30720 30723
0 30725 5 1 1 30724
0 30726 7 1 2 94294 30725
0 30727 5 1 1 30726
0 30728 7 1 2 30708 30727
0 30729 5 1 1 30728
0 30730 7 1 2 77567 30729
0 30731 5 1 1 30730
0 30732 7 1 2 30677 30731
0 30733 5 1 1 30732
0 30734 7 1 2 66853 30733
0 30735 5 1 1 30734
0 30736 7 1 2 84143 90432
0 30737 5 1 1 30736
0 30738 7 1 2 78071 88285
0 30739 7 1 2 94167 30738
0 30740 5 1 1 30739
0 30741 7 1 2 30737 30740
0 30742 5 1 1 30741
0 30743 7 1 2 80735 30742
0 30744 5 1 1 30743
0 30745 7 2 2 74068 94149
0 30746 7 1 2 75440 84434
0 30747 7 1 2 94445 30746
0 30748 5 1 1 30747
0 30749 7 1 2 30744 30748
0 30750 5 1 1 30749
0 30751 7 1 2 66304 30750
0 30752 5 1 1 30751
0 30753 7 1 2 76018 84930
0 30754 7 1 2 94446 30753
0 30755 5 1 1 30754
0 30756 7 1 2 30752 30755
0 30757 5 1 1 30756
0 30758 7 1 2 62680 30757
0 30759 5 1 1 30758
0 30760 7 1 2 80368 88208
0 30761 5 1 1 30760
0 30762 7 1 2 65229 30761
0 30763 5 1 1 30762
0 30764 7 1 2 70060 81184
0 30765 5 1 1 30764
0 30766 7 1 2 30763 30765
0 30767 5 1 1 30766
0 30768 7 1 2 77200 92145
0 30769 7 1 2 30767 30768
0 30770 5 1 1 30769
0 30771 7 1 2 30759 30770
0 30772 5 1 1 30771
0 30773 7 1 2 63998 30772
0 30774 5 1 1 30773
0 30775 7 4 2 65438 80998
0 30776 7 2 2 77969 94447
0 30777 7 1 2 87819 94451
0 30778 5 1 1 30777
0 30779 7 1 2 30774 30778
0 30780 5 1 1 30779
0 30781 7 1 2 66854 30780
0 30782 5 1 1 30781
0 30783 7 2 2 78709 87859
0 30784 7 1 2 86291 87823
0 30785 7 1 2 94453 30784
0 30786 7 1 2 85811 30785
0 30787 5 1 1 30786
0 30788 7 1 2 30782 30787
0 30789 5 1 1 30788
0 30790 7 1 2 69664 30789
0 30791 5 1 1 30790
0 30792 7 1 2 79378 87046
0 30793 7 1 2 87843 30792
0 30794 7 1 2 88320 94101
0 30795 7 1 2 30793 30794
0 30796 5 1 1 30795
0 30797 7 1 2 60664 30796
0 30798 7 1 2 30791 30797
0 30799 7 1 2 30735 30798
0 30800 5 1 1 30799
0 30801 7 1 2 64092 30800
0 30802 7 1 2 30579 30801
0 30803 5 1 1 30802
0 30804 7 1 2 74405 93767
0 30805 5 1 1 30804
0 30806 7 2 2 62325 73952
0 30807 5 1 1 94455
0 30808 7 2 2 79261 94456
0 30809 5 1 1 94457
0 30810 7 1 2 30805 30809
0 30811 5 1 1 30810
0 30812 7 1 2 65230 30811
0 30813 5 1 1 30812
0 30814 7 4 2 62326 80419
0 30815 7 1 2 73953 94459
0 30816 5 1 1 30815
0 30817 7 1 2 30813 30816
0 30818 5 1 1 30817
0 30819 7 1 2 90337 30818
0 30820 5 1 1 30819
0 30821 7 1 2 85600 91212
0 30822 5 1 1 30821
0 30823 7 1 2 30820 30822
0 30824 5 1 1 30823
0 30825 7 1 2 68024 30824
0 30826 5 1 1 30825
0 30827 7 2 2 64997 75666
0 30828 5 1 1 94463
0 30829 7 1 2 88856 94460
0 30830 7 1 2 94464 30829
0 30831 5 1 1 30830
0 30832 7 1 2 30826 30831
0 30833 5 1 1 30832
0 30834 7 1 2 87170 30833
0 30835 5 1 1 30834
0 30836 7 2 2 80954 94252
0 30837 7 1 2 81497 92767
0 30838 7 1 2 94465 30837
0 30839 5 1 1 30838
0 30840 7 1 2 30835 30839
0 30841 5 1 1 30840
0 30842 7 1 2 87860 30841
0 30843 5 1 1 30842
0 30844 7 2 2 77787 87462
0 30845 5 1 1 94467
0 30846 7 1 2 82354 30845
0 30847 5 1 1 30846
0 30848 7 1 2 75591 30847
0 30849 5 1 1 30848
0 30850 7 1 2 85737 89219
0 30851 5 1 1 30850
0 30852 7 1 2 64293 30851
0 30853 5 1 1 30852
0 30854 7 1 2 67656 85396
0 30855 5 1 1 30854
0 30856 7 1 2 30853 30855
0 30857 5 1 1 30856
0 30858 7 1 2 64998 30857
0 30859 5 1 1 30858
0 30860 7 1 2 30849 30859
0 30861 5 1 1 30860
0 30862 7 1 2 87638 30861
0 30863 5 1 1 30862
0 30864 7 1 2 94171 94468
0 30865 5 1 1 30864
0 30866 7 1 2 84227 87600
0 30867 5 6 1 30866
0 30868 7 1 2 64294 94469
0 30869 5 1 1 30868
0 30870 7 1 2 80420 93507
0 30871 5 1 1 30870
0 30872 7 1 2 86036 93407
0 30873 5 1 1 30872
0 30874 7 1 2 30871 30873
0 30875 7 1 2 30869 30874
0 30876 5 1 1 30875
0 30877 7 1 2 76643 30876
0 30878 5 1 1 30877
0 30879 7 1 2 30696 30878
0 30880 5 1 1 30879
0 30881 7 1 2 64999 30880
0 30882 5 1 1 30881
0 30883 7 1 2 78257 94172
0 30884 5 1 1 30883
0 30885 7 1 2 30882 30884
0 30886 5 1 1 30885
0 30887 7 1 2 63490 30886
0 30888 5 1 1 30887
0 30889 7 1 2 30865 30888
0 30890 5 1 1 30889
0 30891 7 1 2 86782 30890
0 30892 5 1 1 30891
0 30893 7 1 2 30863 30892
0 30894 5 1 1 30893
0 30895 7 1 2 63999 30894
0 30896 5 1 1 30895
0 30897 7 2 2 74738 77788
0 30898 5 1 1 94475
0 30899 7 1 2 85739 30898
0 30900 5 1 1 30899
0 30901 7 1 2 71561 30900
0 30902 5 1 1 30901
0 30903 7 1 2 76744 94301
0 30904 5 1 1 30903
0 30905 7 1 2 77475 90421
0 30906 5 1 1 30905
0 30907 7 1 2 30904 30906
0 30908 5 1 1 30907
0 30909 7 1 2 64295 30908
0 30910 5 1 1 30909
0 30911 7 1 2 79109 30910
0 30912 5 1 1 30911
0 30913 7 1 2 68376 30912
0 30914 5 1 1 30913
0 30915 7 1 2 30902 30914
0 30916 5 1 1 30915
0 30917 7 3 2 80691 86711
0 30918 7 1 2 30916 94477
0 30919 5 1 1 30918
0 30920 7 1 2 30896 30919
0 30921 5 1 1 30920
0 30922 7 1 2 71790 30921
0 30923 5 1 1 30922
0 30924 7 1 2 84161 82531
0 30925 7 1 2 88066 30924
0 30926 5 1 1 30925
0 30927 7 1 2 62327 87391
0 30928 7 1 2 93552 30927
0 30929 5 1 1 30928
0 30930 7 1 2 30926 30929
0 30931 5 1 1 30930
0 30932 7 1 2 68025 30931
0 30933 5 1 1 30932
0 30934 7 1 2 87997 93703
0 30935 5 1 1 30934
0 30936 7 1 2 30933 30935
0 30937 5 1 1 30936
0 30938 7 1 2 80032 30937
0 30939 5 1 1 30938
0 30940 7 2 2 62328 86712
0 30941 7 1 2 81303 93838
0 30942 7 1 2 94480 30941
0 30943 5 1 1 30942
0 30944 7 1 2 30939 30943
0 30945 5 1 1 30944
0 30946 7 1 2 65439 30945
0 30947 5 1 1 30946
0 30948 7 2 2 78872 79730
0 30949 7 1 2 87171 94482
0 30950 5 1 1 30949
0 30951 7 5 2 86713 87264
0 30952 7 1 2 84994 94484
0 30953 5 1 1 30952
0 30954 7 1 2 30950 30953
0 30955 5 1 1 30954
0 30956 7 1 2 79625 30955
0 30957 5 1 1 30956
0 30958 7 1 2 87639 94483
0 30959 5 1 1 30958
0 30960 7 1 2 30957 30959
0 30961 5 1 1 30960
0 30962 7 1 2 71562 30961
0 30963 5 1 1 30962
0 30964 7 1 2 81304 86783
0 30965 5 1 1 30964
0 30966 7 1 2 87645 30965
0 30967 5 1 1 30966
0 30968 7 2 2 68026 79731
0 30969 7 1 2 85041 94489
0 30970 7 1 2 30967 30969
0 30971 5 1 1 30970
0 30972 7 1 2 30963 30971
0 30973 7 1 2 30947 30972
0 30974 5 1 1 30973
0 30975 7 1 2 67657 30974
0 30976 5 1 1 30975
0 30977 7 1 2 87489 94154
0 30978 5 1 1 30977
0 30979 7 1 2 79262 81028
0 30980 7 1 2 79406 91053
0 30981 7 1 2 30979 30980
0 30982 5 1 1 30981
0 30983 7 1 2 75592 79440
0 30984 7 1 2 88575 30983
0 30985 5 1 1 30984
0 30986 7 1 2 66305 81105
0 30987 7 1 2 90714 30986
0 30988 5 1 1 30987
0 30989 7 1 2 30985 30988
0 30990 5 1 1 30989
0 30991 7 1 2 65440 30990
0 30992 5 1 1 30991
0 30993 7 1 2 85042 85678
0 30994 7 1 2 86881 30993
0 30995 5 1 1 30994
0 30996 7 1 2 30992 30995
0 30997 5 1 1 30996
0 30998 7 1 2 87265 88857
0 30999 7 1 2 30997 30998
0 31000 5 1 1 30999
0 31001 7 1 2 30982 31000
0 31002 5 1 1 31001
0 31003 7 1 2 66855 31002
0 31004 5 1 1 31003
0 31005 7 1 2 86059 93671
0 31006 7 1 2 94391 31005
0 31007 5 1 1 31006
0 31008 7 1 2 31004 31007
0 31009 5 1 1 31008
0 31010 7 1 2 65581 31009
0 31011 5 1 1 31010
0 31012 7 1 2 30978 31011
0 31013 7 1 2 30976 31012
0 31014 7 1 2 30923 31013
0 31015 5 1 1 31014
0 31016 7 1 2 68702 31015
0 31017 5 1 1 31016
0 31018 7 1 2 30843 31017
0 31019 5 1 1 31018
0 31020 7 1 2 64093 31019
0 31021 5 1 1 31020
0 31022 7 1 2 84635 87416
0 31023 7 1 2 79122 31022
0 31024 7 1 2 94237 31023
0 31025 5 1 1 31024
0 31026 7 1 2 31021 31025
0 31027 5 1 1 31026
0 31028 7 1 2 70313 31027
0 31029 5 1 1 31028
0 31030 7 2 2 64534 94461
0 31031 7 2 2 65000 94092
0 31032 5 1 1 94493
0 31033 7 2 2 80540 79016
0 31034 7 1 2 77970 86714
0 31035 7 1 2 94495 31034
0 31036 5 1 1 31035
0 31037 7 1 2 31032 31036
0 31038 5 1 1 31037
0 31039 7 1 2 94491 31038
0 31040 5 1 1 31039
0 31041 7 3 2 77568 87505
0 31042 5 1 1 94497
0 31043 7 1 2 75070 94498
0 31044 5 1 1 31043
0 31045 7 1 2 31040 31044
0 31046 5 1 1 31045
0 31047 7 1 2 66529 31046
0 31048 5 1 1 31047
0 31049 7 1 2 81772 93913
0 31050 7 1 2 94494 31049
0 31051 5 1 1 31050
0 31052 7 1 2 31048 31051
0 31053 5 1 1 31052
0 31054 7 1 2 64094 31053
0 31055 5 1 1 31054
0 31056 7 1 2 82509 88026
0 31057 7 1 2 94233 31056
0 31058 5 1 1 31057
0 31059 7 1 2 31055 31058
0 31060 5 1 1 31059
0 31061 7 1 2 88439 31060
0 31062 5 1 1 31061
0 31063 7 1 2 31029 31062
0 31064 7 1 2 30803 31063
0 31065 7 1 2 29829 31064
0 31066 5 1 1 31065
0 31067 7 1 2 72341 31066
0 31068 5 1 1 31067
0 31069 7 1 2 81645 79104
0 31070 7 1 2 81980 31069
0 31071 5 1 1 31070
0 31072 7 1 2 30083 31071
0 31073 5 1 1 31072
0 31074 7 1 2 65441 31073
0 31075 5 1 1 31074
0 31076 7 1 2 68377 84764
0 31077 5 1 1 31076
0 31078 7 1 2 82355 31077
0 31079 5 1 1 31078
0 31080 7 1 2 88666 31079
0 31081 5 1 1 31080
0 31082 7 1 2 79940 80608
0 31083 5 1 1 31082
0 31084 7 1 2 70986 78614
0 31085 5 4 1 31084
0 31086 7 1 2 85107 94500
0 31087 5 1 1 31086
0 31088 7 1 2 70975 86688
0 31089 5 1 1 31088
0 31090 7 1 2 94340 31089
0 31091 7 1 2 31087 31090
0 31092 5 1 1 31091
0 31093 7 1 2 68378 31092
0 31094 5 1 1 31093
0 31095 7 1 2 31083 31094
0 31096 5 1 1 31095
0 31097 7 1 2 62681 31096
0 31098 5 1 1 31097
0 31099 7 1 2 31081 31098
0 31100 5 1 1 31099
0 31101 7 1 2 62329 31100
0 31102 5 1 1 31101
0 31103 7 1 2 73750 13273
0 31104 5 2 1 31103
0 31105 7 1 2 69836 94504
0 31106 5 2 1 31105
0 31107 7 2 2 66306 71791
0 31108 5 2 1 94508
0 31109 7 1 2 67658 94509
0 31110 5 1 1 31109
0 31111 7 1 2 94506 31110
0 31112 5 1 1 31111
0 31113 7 1 2 62118 31112
0 31114 5 1 1 31113
0 31115 7 1 2 82211 86912
0 31116 5 1 1 31115
0 31117 7 1 2 31114 31116
0 31118 5 1 1 31117
0 31119 7 1 2 77906 31118
0 31120 5 1 1 31119
0 31121 7 1 2 31102 31120
0 31122 5 1 1 31121
0 31123 7 1 2 60544 31122
0 31124 5 1 1 31123
0 31125 7 2 2 62119 76678
0 31126 7 1 2 24449 94512
0 31127 5 1 1 31126
0 31128 7 1 2 82453 31127
0 31129 5 1 1 31128
0 31130 7 5 2 61562 83744
0 31131 7 1 2 77971 94514
0 31132 7 1 2 31129 31131
0 31133 5 1 1 31132
0 31134 7 1 2 31124 31133
0 31135 5 1 1 31134
0 31136 7 1 2 64000 31135
0 31137 5 1 1 31136
0 31138 7 1 2 31075 31137
0 31139 5 1 1 31138
0 31140 7 1 2 61873 31139
0 31141 5 1 1 31140
0 31142 7 1 2 84831 85651
0 31143 5 1 1 31142
0 31144 7 1 2 9153 31143
0 31145 5 1 1 31144
0 31146 7 1 2 86203 31145
0 31147 5 1 1 31146
0 31148 7 2 2 76869 91054
0 31149 5 1 1 94519
0 31150 7 1 2 75419 94520
0 31151 5 1 1 31150
0 31152 7 1 2 77972 93727
0 31153 5 1 1 31152
0 31154 7 1 2 31151 31153
0 31155 5 1 1 31154
0 31156 7 1 2 71792 86092
0 31157 7 1 2 31155 31156
0 31158 5 1 1 31157
0 31159 7 1 2 31147 31158
0 31160 5 1 1 31159
0 31161 7 1 2 68379 31160
0 31162 5 1 1 31161
0 31163 7 1 2 73751 90818
0 31164 5 2 1 31163
0 31165 7 1 2 86218 91361
0 31166 7 1 2 94521 31165
0 31167 5 1 1 31166
0 31168 7 1 2 31162 31167
0 31169 5 1 1 31168
0 31170 7 1 2 62330 31169
0 31171 5 1 1 31170
0 31172 7 1 2 84648 85910
0 31173 5 1 1 31172
0 31174 7 1 2 90622 31173
0 31175 5 1 1 31174
0 31176 7 1 2 64535 31175
0 31177 5 1 1 31176
0 31178 7 1 2 60545 86850
0 31179 5 1 1 31178
0 31180 7 1 2 31177 31179
0 31181 5 1 1 31180
0 31182 7 1 2 67659 31181
0 31183 5 1 1 31182
0 31184 7 1 2 30591 31183
0 31185 5 1 1 31184
0 31186 7 1 2 77403 86093
0 31187 7 1 2 31185 31186
0 31188 5 1 1 31187
0 31189 7 1 2 31171 31188
0 31190 5 1 1 31189
0 31191 7 1 2 69665 31190
0 31192 5 1 1 31191
0 31193 7 1 2 72654 84677
0 31194 5 1 1 31193
0 31195 7 1 2 85423 92887
0 31196 5 1 1 31195
0 31197 7 1 2 31194 31196
0 31198 5 1 1 31197
0 31199 7 2 2 75593 31198
0 31200 5 1 1 94523
0 31201 7 1 2 94367 94524
0 31202 5 1 1 31201
0 31203 7 1 2 63764 31202
0 31204 7 1 2 31192 31203
0 31205 7 1 2 31141 31204
0 31206 5 1 1 31205
0 31207 7 1 2 73178 84406
0 31208 5 1 1 31207
0 31209 7 1 2 79925 31208
0 31210 5 1 1 31209
0 31211 7 1 2 74509 94286
0 31212 5 1 1 31211
0 31213 7 1 2 31210 31212
0 31214 5 1 1 31213
0 31215 7 1 2 63491 31214
0 31216 5 1 1 31215
0 31217 7 1 2 83169 31216
0 31218 5 1 1 31217
0 31219 7 1 2 69666 31218
0 31220 5 1 1 31219
0 31221 7 1 2 83920 77406
0 31222 5 1 1 31221
0 31223 7 2 2 69837 31222
0 31224 5 1 1 94525
0 31225 7 1 2 84739 94526
0 31226 5 1 1 31225
0 31227 7 1 2 83170 31226
0 31228 5 1 1 31227
0 31229 7 1 2 71793 31228
0 31230 5 1 1 31229
0 31231 7 2 2 68380 73042
0 31232 7 1 2 75217 94527
0 31233 5 1 1 31232
0 31234 7 2 2 76852 86658
0 31235 7 1 2 69985 94529
0 31236 5 1 1 31235
0 31237 7 1 2 84083 86846
0 31238 5 1 1 31237
0 31239 7 1 2 31236 31238
0 31240 5 1 1 31239
0 31241 7 1 2 71993 31240
0 31242 5 1 1 31241
0 31243 7 1 2 31233 31242
0 31244 7 1 2 31230 31243
0 31245 7 1 2 31220 31244
0 31246 5 1 1 31245
0 31247 7 1 2 86094 31246
0 31248 5 1 1 31247
0 31249 7 1 2 75667 84984
0 31250 5 1 1 31249
0 31251 7 1 2 67660 875
0 31252 5 1 1 31251
0 31253 7 1 2 79776 76212
0 31254 7 1 2 31252 31253
0 31255 5 1 1 31254
0 31256 7 1 2 31250 31255
0 31257 5 1 1 31256
0 31258 7 1 2 69667 31257
0 31259 5 1 1 31258
0 31260 7 1 2 79777 72595
0 31261 5 1 1 31260
0 31262 7 1 2 68381 91231
0 31263 5 1 1 31262
0 31264 7 1 2 31261 31263
0 31265 5 1 1 31264
0 31266 7 1 2 69253 31265
0 31267 5 1 1 31266
0 31268 7 1 2 79778 7468
0 31269 5 1 1 31268
0 31270 7 4 2 62331 75594
0 31271 5 2 1 94531
0 31272 7 2 2 68382 94532
0 31273 7 1 2 78609 94537
0 31274 5 1 1 31273
0 31275 7 1 2 31269 31274
0 31276 7 1 2 31267 31275
0 31277 5 1 1 31276
0 31278 7 1 2 62120 31277
0 31279 5 1 1 31278
0 31280 7 1 2 79779 75954
0 31281 5 1 1 31280
0 31282 7 1 2 67661 31281
0 31283 7 1 2 31279 31282
0 31284 5 1 1 31283
0 31285 7 1 2 77214 94305
0 31286 5 1 1 31285
0 31287 7 1 2 8521 31286
0 31288 5 1 1 31287
0 31289 7 1 2 68383 31288
0 31290 5 1 1 31289
0 31291 7 1 2 79780 90348
0 31292 7 1 2 78361 31291
0 31293 5 1 1 31292
0 31294 7 1 2 62682 31293
0 31295 7 1 2 31290 31294
0 31296 5 1 1 31295
0 31297 7 1 2 31284 31296
0 31298 5 1 1 31297
0 31299 7 1 2 31259 31298
0 31300 5 1 1 31299
0 31301 7 1 2 66307 31300
0 31302 5 1 1 31301
0 31303 7 1 2 63492 81921
0 31304 7 1 2 81255 70949
0 31305 7 1 2 31303 31304
0 31306 7 1 2 71454 31305
0 31307 5 1 1 31306
0 31308 7 1 2 63046 31307
0 31309 7 1 2 79890 80478
0 31310 7 1 2 90693 31309
0 31311 5 1 1 31310
0 31312 7 1 2 75405 93734
0 31313 7 1 2 94280 31312
0 31314 5 1 1 31313
0 31315 7 1 2 31311 31314
0 31316 7 1 2 31308 31315
0 31317 7 1 2 31302 31316
0 31318 5 1 1 31317
0 31319 7 1 2 75098 88390
0 31320 5 1 1 31319
0 31321 7 1 2 67662 90924
0 31322 5 1 1 31321
0 31323 7 1 2 31320 31322
0 31324 5 1 1 31323
0 31325 7 1 2 61352 31324
0 31326 5 1 1 31325
0 31327 7 1 2 62121 78018
0 31328 5 1 1 31327
0 31329 7 1 2 31326 31328
0 31330 5 1 1 31329
0 31331 7 1 2 63493 31330
0 31332 5 1 1 31331
0 31333 7 2 2 62122 77215
0 31334 5 1 1 94539
0 31335 7 1 2 75812 31334
0 31336 5 1 1 31335
0 31337 7 1 2 62683 31336
0 31338 5 1 1 31337
0 31339 7 1 2 74471 31338
0 31340 5 1 1 31339
0 31341 7 1 2 75071 31340
0 31342 5 1 1 31341
0 31343 7 1 2 31332 31342
0 31344 5 1 1 31343
0 31345 7 1 2 66530 31344
0 31346 5 1 1 31345
0 31347 7 1 2 82734 86913
0 31348 5 1 1 31347
0 31349 7 1 2 60365 31348
0 31350 5 1 1 31349
0 31351 7 1 2 62684 31350
0 31352 5 1 1 31351
0 31353 7 3 2 65231 69668
0 31354 5 1 1 94541
0 31355 7 1 2 82576 94542
0 31356 5 1 1 31355
0 31357 7 1 2 31352 31356
0 31358 5 1 1 31357
0 31359 7 1 2 62123 31358
0 31360 5 1 1 31359
0 31361 7 1 2 73521 77535
0 31362 5 1 1 31361
0 31363 7 1 2 31360 31362
0 31364 5 1 1 31363
0 31365 7 1 2 79781 31364
0 31366 5 1 1 31365
0 31367 7 1 2 68027 31366
0 31368 7 1 2 31346 31367
0 31369 5 1 1 31368
0 31370 7 1 2 86165 31369
0 31371 7 1 2 31318 31370
0 31372 5 1 1 31371
0 31373 7 1 2 31248 31372
0 31374 5 1 1 31373
0 31375 7 1 2 65442 31374
0 31376 5 1 1 31375
0 31377 7 1 2 94109 94430
0 31378 5 1 1 31377
0 31379 7 2 2 66531 86166
0 31380 7 1 2 60546 94544
0 31381 5 1 1 31380
0 31382 7 1 2 31378 31381
0 31383 5 1 1 31382
0 31384 7 1 2 65232 31383
0 31385 5 1 1 31384
0 31386 7 1 2 78951 91055
0 31387 7 1 2 94110 31386
0 31388 5 1 1 31387
0 31389 7 1 2 31385 31388
0 31390 5 1 1 31389
0 31391 7 1 2 70453 31390
0 31392 5 1 1 31391
0 31393 7 1 2 72856 82883
0 31394 5 1 1 31393
0 31395 7 1 2 85646 86167
0 31396 7 1 2 31394 31395
0 31397 5 1 1 31396
0 31398 7 1 2 31392 31397
0 31399 5 1 1 31398
0 31400 7 1 2 66308 31399
0 31401 5 1 1 31400
0 31402 7 1 2 85480 86095
0 31403 7 1 2 88484 31402
0 31404 5 1 1 31403
0 31405 7 1 2 31401 31404
0 31406 5 1 1 31405
0 31407 7 1 2 63047 31406
0 31408 5 1 1 31407
0 31409 7 1 2 75218 86096
0 31410 7 1 2 94287 31409
0 31411 7 1 2 88744 31410
0 31412 5 1 1 31411
0 31413 7 1 2 31408 31412
0 31414 5 1 1 31413
0 31415 7 1 2 62332 31414
0 31416 5 1 1 31415
0 31417 7 2 2 77404 82212
0 31418 5 1 1 94546
0 31419 7 1 2 70976 94547
0 31420 5 1 1 31419
0 31421 7 1 2 73179 12410
0 31422 5 3 1 31421
0 31423 7 1 2 60547 69669
0 31424 7 1 2 94548 31423
0 31425 5 1 1 31424
0 31426 7 1 2 31420 31425
0 31427 5 1 1 31426
0 31428 7 1 2 75420 87456
0 31429 7 1 2 31427 31428
0 31430 5 1 1 31429
0 31431 7 1 2 31416 31430
0 31432 5 1 1 31431
0 31433 7 1 2 63494 31432
0 31434 5 1 1 31433
0 31435 7 1 2 79891 87211
0 31436 7 1 2 88148 31435
0 31437 7 1 2 78316 31436
0 31438 5 1 1 31437
0 31439 7 1 2 68703 31438
0 31440 7 1 2 31434 31439
0 31441 7 1 2 31376 31440
0 31442 5 1 1 31441
0 31443 7 1 2 66711 31442
0 31444 7 1 2 31206 31443
0 31445 5 1 1 31444
0 31446 7 1 2 85094 31418
0 31447 5 1 1 31446
0 31448 7 1 2 65726 31447
0 31449 5 1 1 31448
0 31450 7 1 2 82110 78283
0 31451 5 1 1 31450
0 31452 7 1 2 31449 31451
0 31453 5 1 1 31452
0 31454 7 1 2 64536 31453
0 31455 5 1 1 31454
0 31456 7 1 2 85095 31224
0 31457 5 1 1 31456
0 31458 7 2 2 69670 31457
0 31459 7 1 2 65881 94551
0 31460 5 1 1 31459
0 31461 7 1 2 31455 31460
0 31462 5 1 1 31461
0 31463 7 1 2 62333 31462
0 31464 5 1 1 31463
0 31465 7 1 2 70416 94288
0 31466 5 1 1 31465
0 31467 7 1 2 78407 83907
0 31468 5 1 1 31467
0 31469 7 1 2 31466 31468
0 31470 5 1 1 31469
0 31471 7 1 2 70454 31470
0 31472 5 1 1 31471
0 31473 7 1 2 31464 31472
0 31474 5 1 1 31473
0 31475 7 1 2 63495 31474
0 31476 5 1 1 31475
0 31477 7 1 2 65233 73073
0 31478 5 1 1 31477
0 31479 7 3 2 63048 77237
0 31480 5 1 1 94553
0 31481 7 1 2 91384 94554
0 31482 5 1 1 31481
0 31483 7 1 2 31478 31482
0 31484 5 1 1 31483
0 31485 7 1 2 75848 31484
0 31486 5 1 1 31485
0 31487 7 1 2 79782 71455
0 31488 5 1 1 31487
0 31489 7 1 2 81867 87880
0 31490 5 1 1 31489
0 31491 7 1 2 31488 31490
0 31492 5 1 1 31491
0 31493 7 1 2 94549 31492
0 31494 5 1 1 31493
0 31495 7 1 2 31486 31494
0 31496 7 1 2 31476 31495
0 31497 5 1 1 31496
0 31498 7 1 2 60548 31497
0 31499 5 1 1 31498
0 31500 7 1 2 76719 77529
0 31501 7 1 2 87905 31500
0 31502 5 1 1 31501
0 31503 7 1 2 60549 31502
0 31504 5 1 1 31503
0 31505 7 1 2 78317 94338
0 31506 7 1 2 31504 31505
0 31507 5 1 1 31506
0 31508 7 1 2 31499 31507
0 31509 5 1 1 31508
0 31510 7 1 2 68704 31509
0 31511 5 1 1 31510
0 31512 7 3 2 61563 78258
0 31513 7 1 2 92155 94556
0 31514 5 1 1 31513
0 31515 7 1 2 66856 31514
0 31516 7 1 2 31511 31515
0 31517 5 1 1 31516
0 31518 7 1 2 74069 73742
0 31519 5 2 1 31518
0 31520 7 1 2 94507 94559
0 31521 5 1 1 31520
0 31522 7 1 2 62124 31521
0 31523 5 1 1 31522
0 31524 7 1 2 73743 74503
0 31525 5 1 1 31524
0 31526 7 1 2 73689 84908
0 31527 5 1 1 31526
0 31528 7 1 2 94560 31527
0 31529 5 1 1 31528
0 31530 7 1 2 69671 31529
0 31531 5 1 1 31530
0 31532 7 1 2 31525 31531
0 31533 7 1 2 31523 31532
0 31534 5 1 1 31533
0 31535 7 1 2 77907 31534
0 31536 5 1 1 31535
0 31537 7 1 2 77522 92888
0 31538 5 1 1 31537
0 31539 7 1 2 31536 31538
0 31540 5 1 1 31539
0 31541 7 1 2 91855 31540
0 31542 5 1 1 31541
0 31543 7 1 2 81408 91014
0 31544 5 1 1 31543
0 31545 7 2 2 66532 69672
0 31546 5 2 1 94561
0 31547 7 2 2 31354 94563
0 31548 5 3 1 94565
0 31549 7 1 2 65882 82177
0 31550 7 1 2 94567 31549
0 31551 5 1 1 31550
0 31552 7 1 2 31544 31551
0 31553 5 1 1 31552
0 31554 7 1 2 62125 31553
0 31555 5 1 1 31554
0 31556 7 1 2 93644 93650
0 31557 5 1 1 31556
0 31558 7 1 2 31555 31557
0 31559 5 1 1 31558
0 31560 7 1 2 62685 31559
0 31561 5 1 1 31560
0 31562 7 1 2 80515 93651
0 31563 5 1 1 31562
0 31564 7 1 2 31561 31563
0 31565 5 1 1 31564
0 31566 7 1 2 64537 31565
0 31567 5 1 1 31566
0 31568 7 1 2 75925 86857
0 31569 7 1 2 91015 31568
0 31570 5 1 1 31569
0 31571 7 1 2 31567 31570
0 31572 5 1 1 31571
0 31573 7 1 2 62334 31572
0 31574 5 1 1 31573
0 31575 7 1 2 31542 31574
0 31576 5 1 1 31575
0 31577 7 1 2 63765 31576
0 31578 5 1 1 31577
0 31579 7 1 2 72438 73170
0 31580 5 2 1 31579
0 31581 7 1 2 75317 94570
0 31582 5 1 1 31581
0 31583 7 1 2 93394 31582
0 31584 5 1 1 31583
0 31585 7 1 2 90718 31584
0 31586 5 1 1 31585
0 31587 7 1 2 64296 31586
0 31588 5 1 1 31587
0 31589 7 1 2 69254 91294
0 31590 5 1 1 31589
0 31591 7 1 2 31588 31590
0 31592 5 1 1 31591
0 31593 7 1 2 64538 31592
0 31594 5 1 1 31593
0 31595 7 1 2 75219 88378
0 31596 5 1 1 31595
0 31597 7 1 2 31594 31596
0 31598 5 1 1 31597
0 31599 7 1 2 63049 31598
0 31600 5 1 1 31599
0 31601 7 1 2 74130 87528
0 31602 5 1 1 31601
0 31603 7 1 2 31600 31602
0 31604 5 1 1 31603
0 31605 7 1 2 62126 31604
0 31606 5 1 1 31605
0 31607 7 1 2 93784 93660
0 31608 5 1 1 31607
0 31609 7 1 2 31606 31608
0 31610 5 1 1 31609
0 31611 7 1 2 84215 31610
0 31612 5 1 1 31611
0 31613 7 1 2 61874 31612
0 31614 7 1 2 31578 31613
0 31615 5 1 1 31614
0 31616 7 1 2 64001 31615
0 31617 7 1 2 31517 31616
0 31618 5 1 1 31617
0 31619 7 2 2 62335 75421
0 31620 7 1 2 69673 75072
0 31621 7 1 2 94572 31620
0 31622 5 1 1 31621
0 31623 7 1 2 31200 31622
0 31624 5 1 1 31623
0 31625 7 1 2 63766 31624
0 31626 5 1 1 31625
0 31627 7 1 2 71726 69408
0 31628 5 3 1 31627
0 31629 7 2 2 64297 94574
0 31630 5 1 1 94577
0 31631 7 3 2 82885 31630
0 31632 5 4 1 94579
0 31633 7 2 2 85043 89966
0 31634 7 1 2 78572 94586
0 31635 7 1 2 94582 31634
0 31636 5 1 1 31635
0 31637 7 1 2 31626 31636
0 31638 5 1 1 31637
0 31639 7 1 2 68883 87541
0 31640 7 1 2 31638 31639
0 31641 5 1 1 31640
0 31642 7 1 2 31618 31641
0 31643 5 1 1 31642
0 31644 7 1 2 61731 31643
0 31645 5 1 1 31644
0 31646 7 1 2 77973 86354
0 31647 7 1 2 87824 31646
0 31648 7 1 2 92517 31647
0 31649 7 1 2 89213 31648
0 31650 5 1 1 31649
0 31651 7 1 2 65582 31650
0 31652 7 1 2 31645 31651
0 31653 7 1 2 31445 31652
0 31654 5 1 1 31653
0 31655 7 1 2 92419 94530
0 31656 5 1 1 31655
0 31657 7 1 2 81106 90685
0 31658 5 1 1 31657
0 31659 7 1 2 79456 31658
0 31660 5 1 1 31659
0 31661 7 1 2 62336 86835
0 31662 7 1 2 31660 31661
0 31663 5 1 1 31662
0 31664 7 1 2 31656 31663
0 31665 5 1 1 31664
0 31666 7 1 2 65443 31665
0 31667 5 1 1 31666
0 31668 7 1 2 85075 94299
0 31669 5 1 1 31668
0 31670 7 1 2 65234 31669
0 31671 5 1 1 31670
0 31672 7 1 2 77516 85451
0 31673 5 1 1 31672
0 31674 7 1 2 31671 31673
0 31675 5 1 1 31674
0 31676 7 1 2 81952 81286
0 31677 7 1 2 31675 31676
0 31678 5 1 1 31677
0 31679 7 1 2 31667 31678
0 31680 5 1 1 31679
0 31681 7 1 2 69838 31680
0 31682 5 1 1 31681
0 31683 7 1 2 73630 85397
0 31684 7 1 2 94168 31683
0 31685 5 1 1 31684
0 31686 7 1 2 31682 31685
0 31687 5 1 1 31686
0 31688 7 1 2 71994 31687
0 31689 5 1 1 31688
0 31690 7 1 2 79699 94528
0 31691 5 1 1 31690
0 31692 7 1 2 68705 31691
0 31693 7 1 2 31689 31692
0 31694 5 1 1 31693
0 31695 7 1 2 76853 93728
0 31696 5 1 1 31695
0 31697 7 1 2 31149 31696
0 31698 5 1 1 31697
0 31699 7 1 2 69839 31698
0 31700 5 1 1 31699
0 31701 7 1 2 71995 94557
0 31702 5 1 1 31701
0 31703 7 1 2 88166 31702
0 31704 5 1 1 31703
0 31705 7 1 2 66309 31704
0 31706 5 1 1 31705
0 31707 7 1 2 31700 31706
0 31708 5 1 1 31707
0 31709 7 1 2 81297 31708
0 31710 5 1 1 31709
0 31711 7 1 2 65444 86421
0 31712 5 1 1 31711
0 31713 7 1 2 29723 31712
0 31714 5 1 1 31713
0 31715 7 1 2 71996 93758
0 31716 7 1 2 31714 31715
0 31717 5 1 1 31716
0 31718 7 1 2 31710 31717
0 31719 5 1 1 31718
0 31720 7 1 2 68384 31719
0 31721 5 1 1 31720
0 31722 7 1 2 71997 86858
0 31723 7 1 2 93800 31722
0 31724 5 1 1 31723
0 31725 7 1 2 31721 31724
0 31726 5 1 1 31725
0 31727 7 1 2 62337 31726
0 31728 5 1 1 31727
0 31729 7 1 2 82120 93419
0 31730 5 1 1 31729
0 31731 7 1 2 69986 77908
0 31732 7 1 2 94505 31731
0 31733 5 1 1 31732
0 31734 7 1 2 31730 31733
0 31735 5 1 1 31734
0 31736 7 1 2 62127 31735
0 31737 5 1 1 31736
0 31738 7 1 2 82121 82346
0 31739 5 1 1 31738
0 31740 7 1 2 31737 31739
0 31741 5 1 1 31740
0 31742 7 1 2 94150 31741
0 31743 5 1 1 31742
0 31744 7 1 2 77974 76009
0 31745 7 1 2 94513 31744
0 31746 5 1 1 31745
0 31747 7 1 2 90903 31746
0 31748 5 1 1 31747
0 31749 7 1 2 86895 31748
0 31750 5 1 1 31749
0 31751 7 1 2 63767 31750
0 31752 7 1 2 31743 31751
0 31753 7 1 2 31728 31752
0 31754 5 1 1 31753
0 31755 7 1 2 31694 31754
0 31756 5 1 1 31755
0 31757 7 1 2 81911 93729
0 31758 5 1 1 31757
0 31759 7 2 2 62128 80331
0 31760 7 1 2 76644 94588
0 31761 5 1 1 31760
0 31762 7 1 2 31758 31761
0 31763 5 1 1 31762
0 31764 7 1 2 65235 31763
0 31765 5 1 1 31764
0 31766 7 1 2 84113 94138
0 31767 5 1 1 31766
0 31768 7 1 2 31765 31767
0 31769 5 1 1 31768
0 31770 7 1 2 71998 31769
0 31771 5 1 1 31770
0 31772 7 1 2 65236 74370
0 31773 7 1 2 85176 31772
0 31774 5 1 1 31773
0 31775 7 1 2 31771 31774
0 31776 5 1 1 31775
0 31777 7 1 2 63768 31776
0 31778 5 1 1 31777
0 31779 7 2 2 68706 79626
0 31780 7 1 2 75220 94590
0 31781 5 1 1 31780
0 31782 7 1 2 68385 31781
0 31783 7 1 2 31778 31782
0 31784 5 1 1 31783
0 31785 7 1 2 75955 94433
0 31786 5 1 1 31785
0 31787 7 1 2 62129 94550
0 31788 7 1 2 94470 31787
0 31789 5 1 1 31788
0 31790 7 1 2 31786 31789
0 31791 5 1 1 31790
0 31792 7 1 2 68707 31791
0 31793 5 1 1 31792
0 31794 7 1 2 62338 84435
0 31795 7 1 2 94151 31794
0 31796 7 1 2 94522 31795
0 31797 5 1 1 31796
0 31798 7 1 2 63496 31797
0 31799 7 1 2 31793 31798
0 31800 5 1 1 31799
0 31801 7 1 2 69674 31800
0 31802 7 1 2 31784 31801
0 31803 5 1 1 31802
0 31804 7 1 2 31756 31803
0 31805 5 1 1 31804
0 31806 7 1 2 66857 31805
0 31807 5 1 1 31806
0 31808 7 2 2 80516 93661
0 31809 7 2 2 85807 93915
0 31810 7 1 2 94592 94594
0 31811 5 1 1 31810
0 31812 7 1 2 90690 93724
0 31813 5 1 1 31812
0 31814 7 1 2 11516 31813
0 31815 5 1 1 31814
0 31816 7 1 2 68708 31815
0 31817 5 1 1 31816
0 31818 7 1 2 90746 94426
0 31819 5 1 1 31818
0 31820 7 2 2 74640 77909
0 31821 5 1 1 94596
0 31822 7 1 2 73744 94597
0 31823 5 2 1 31822
0 31824 7 1 2 31819 94598
0 31825 5 1 1 31824
0 31826 7 1 2 84481 31825
0 31827 5 1 1 31826
0 31828 7 1 2 31817 31827
0 31829 5 1 1 31828
0 31830 7 1 2 66533 31829
0 31831 5 1 1 31830
0 31832 7 2 2 66310 78765
0 31833 5 2 1 94600
0 31834 7 1 2 80172 92171
0 31835 7 1 2 94601 31834
0 31836 7 1 2 90313 31835
0 31837 5 1 1 31836
0 31838 7 1 2 31831 31837
0 31839 5 1 1 31838
0 31840 7 1 2 65237 31839
0 31841 5 1 1 31840
0 31842 7 1 2 90747 94428
0 31843 5 1 1 31842
0 31844 7 1 2 94599 31843
0 31845 5 1 1 31844
0 31846 7 1 2 63769 31845
0 31847 5 1 1 31846
0 31848 7 1 2 90715 91156
0 31849 7 1 2 88460 31848
0 31850 5 1 1 31849
0 31851 7 1 2 31847 31850
0 31852 5 1 1 31851
0 31853 7 1 2 81185 31852
0 31854 5 1 1 31853
0 31855 7 1 2 84740 94591
0 31856 7 1 2 94552 31855
0 31857 5 1 1 31856
0 31858 7 1 2 31854 31857
0 31859 7 1 2 31841 31858
0 31860 5 1 1 31859
0 31861 7 1 2 66858 31860
0 31862 5 1 1 31861
0 31863 7 1 2 31811 31862
0 31864 5 1 1 31863
0 31865 7 1 2 71794 31864
0 31866 5 1 1 31865
0 31867 7 1 2 66311 93836
0 31868 7 1 2 94595 31867
0 31869 5 1 1 31868
0 31870 7 1 2 31866 31869
0 31871 7 1 2 31807 31870
0 31872 5 1 1 31871
0 31873 7 1 2 64002 31872
0 31874 5 1 1 31873
0 31875 7 1 2 87663 92276
0 31876 7 1 2 94593 31875
0 31877 5 1 1 31876
0 31878 7 1 2 60665 31877
0 31879 7 1 2 31874 31878
0 31880 5 1 1 31879
0 31881 7 1 2 64095 31880
0 31882 7 1 2 31654 31881
0 31883 5 1 1 31882
0 31884 7 7 2 68977 87861
0 31885 7 3 2 83102 94604
0 31886 7 1 2 85875 94245
0 31887 7 1 2 94611 31886
0 31888 7 1 2 88488 31887
0 31889 5 1 1 31888
0 31890 7 1 2 31883 31889
0 31891 5 1 1 31890
0 31892 7 1 2 72721 31891
0 31893 5 1 1 31892
0 31894 7 1 2 84704 27336
0 31895 5 1 1 31894
0 31896 7 1 2 91655 31895
0 31897 5 1 1 31896
0 31898 7 1 2 85481 92268
0 31899 5 1 1 31898
0 31900 7 1 2 31897 31899
0 31901 5 1 1 31900
0 31902 7 1 2 68386 31901
0 31903 5 1 1 31902
0 31904 7 1 2 80736 94169
0 31905 5 1 1 31904
0 31906 7 1 2 75144 85679
0 31907 5 1 1 31906
0 31908 7 1 2 31905 31907
0 31909 5 1 1 31908
0 31910 7 1 2 68709 78573
0 31911 7 1 2 31909 31910
0 31912 5 1 1 31911
0 31913 7 2 2 80812 84845
0 31914 5 2 1 94614
0 31915 7 1 2 81298 94615
0 31916 5 1 1 31915
0 31917 7 1 2 83545 78574
0 31918 5 3 1 31917
0 31919 7 1 2 78790 94618
0 31920 5 2 1 31919
0 31921 7 1 2 61732 91656
0 31922 5 1 1 31921
0 31923 7 1 2 92384 31922
0 31924 5 2 1 31923
0 31925 7 1 2 94621 94623
0 31926 5 1 1 31925
0 31927 7 1 2 31916 31926
0 31928 7 1 2 31912 31927
0 31929 5 1 1 31928
0 31930 7 1 2 62686 31929
0 31931 5 1 1 31930
0 31932 7 1 2 80517 89950
0 31933 5 1 1 31932
0 31934 7 1 2 84436 94458
0 31935 5 1 1 31934
0 31936 7 1 2 31933 31935
0 31937 5 1 1 31936
0 31938 7 1 2 65238 31937
0 31939 5 1 1 31938
0 31940 7 3 2 68028 73618
0 31941 7 1 2 92507 94625
0 31942 5 1 1 31941
0 31943 7 1 2 79564 89951
0 31944 5 1 1 31943
0 31945 7 1 2 31942 31944
0 31946 5 1 1 31945
0 31947 7 1 2 65445 31946
0 31948 5 1 1 31947
0 31949 7 1 2 84437 85367
0 31950 7 1 2 93223 31949
0 31951 5 1 1 31950
0 31952 7 1 2 31948 31951
0 31953 7 1 2 31939 31952
0 31954 7 1 2 31931 31953
0 31955 5 1 1 31954
0 31956 7 1 2 77867 31955
0 31957 5 1 1 31956
0 31958 7 1 2 31903 31957
0 31959 5 1 1 31958
0 31960 7 1 2 64762 31959
0 31961 5 1 1 31960
0 31962 7 2 2 66534 80332
0 31963 5 1 1 94628
0 31964 7 1 2 10731 31963
0 31965 5 1 1 31964
0 31966 7 1 2 79044 94626
0 31967 7 1 2 31965 31966
0 31968 5 1 1 31967
0 31969 7 1 2 31961 31968
0 31970 5 1 1 31969
0 31971 7 1 2 86784 31970
0 31972 5 1 1 31971
0 31973 7 2 2 75221 92326
0 31974 7 1 2 93213 94630
0 31975 5 1 1 31974
0 31976 7 1 2 83652 82050
0 31977 7 1 2 88053 31976
0 31978 7 1 2 93751 31977
0 31979 5 1 1 31978
0 31980 7 1 2 31975 31979
0 31981 5 1 1 31980
0 31982 7 1 2 62339 31981
0 31983 5 1 1 31982
0 31984 7 1 2 77990 85468
0 31985 7 7 2 66859 89931
0 31986 7 2 2 65583 66040
0 31987 7 2 2 65001 94639
0 31988 7 1 2 94632 94641
0 31989 7 1 2 31984 31988
0 31990 5 1 1 31989
0 31991 7 1 2 31983 31990
0 31992 7 1 2 31972 31991
0 31993 5 1 1 31992
0 31994 7 1 2 64003 31993
0 31995 5 1 1 31994
0 31996 7 1 2 80737 93439
0 31997 5 1 1 31996
0 31998 7 1 2 79783 93369
0 31999 5 1 1 31998
0 32000 7 1 2 31997 31999
0 32001 5 1 1 32000
0 32002 7 6 2 68884 87069
0 32003 7 7 2 65584 68029
0 32004 5 1 1 94649
0 32005 7 1 2 77991 84186
0 32006 7 1 2 94650 32005
0 32007 7 1 2 94643 32006
0 32008 7 1 2 32001 32007
0 32009 5 1 1 32008
0 32010 7 1 2 31995 32009
0 32011 5 1 1 32010
0 32012 7 1 2 64096 32011
0 32013 5 1 1 32012
0 32014 7 2 2 65585 85496
0 32015 7 1 2 94238 94656
0 32016 5 1 1 32015
0 32017 7 1 2 32013 32016
0 32018 5 1 1 32017
0 32019 7 1 2 79986 32018
0 32020 5 1 1 32019
0 32021 7 1 2 82383 5029
0 32022 5 1 1 32021
0 32023 7 1 2 78766 85044
0 32024 5 2 1 32023
0 32025 7 3 2 69840 74026
0 32026 5 1 1 94660
0 32027 7 2 2 73133 32026
0 32028 5 3 1 94663
0 32029 7 1 2 84869 94665
0 32030 5 1 1 32029
0 32031 7 1 2 93541 32030
0 32032 5 1 1 32031
0 32033 7 1 2 65239 32032
0 32034 5 1 1 32033
0 32035 7 1 2 94658 32034
0 32036 5 1 1 32035
0 32037 7 1 2 72342 32036
0 32038 5 1 1 32037
0 32039 7 2 2 77259 78767
0 32040 7 1 2 77296 94668
0 32041 5 1 1 32040
0 32042 7 1 2 90941 32041
0 32043 5 1 1 32042
0 32044 7 1 2 65002 32043
0 32045 5 1 1 32044
0 32046 7 1 2 77150 92594
0 32047 5 1 1 32046
0 32048 7 2 2 68387 93842
0 32049 7 1 2 83775 94670
0 32050 5 1 1 32049
0 32051 7 1 2 32047 32050
0 32052 7 1 2 32045 32051
0 32053 7 1 2 32038 32052
0 32054 5 1 1 32053
0 32055 7 1 2 86972 32054
0 32056 5 1 1 32055
0 32057 7 1 2 83463 91223
0 32058 5 2 1 32057
0 32059 7 1 2 68388 94672
0 32060 5 2 1 32059
0 32061 7 2 2 63497 72343
0 32062 7 1 2 61564 69987
0 32063 7 1 2 94676 32062
0 32064 5 1 1 32063
0 32065 7 1 2 94674 32064
0 32066 5 1 1 32065
0 32067 7 1 2 85702 32066
0 32068 5 1 1 32067
0 32069 7 1 2 69675 93715
0 32070 5 1 1 32069
0 32071 7 1 2 26778 32070
0 32072 5 1 1 32071
0 32073 7 1 2 77162 94383
0 32074 7 1 2 32072 32073
0 32075 5 1 1 32074
0 32076 7 1 2 32068 32075
0 32077 5 1 1 32076
0 32078 7 1 2 64539 32077
0 32079 5 1 1 32078
0 32080 7 1 2 75595 81868
0 32081 5 1 1 32080
0 32082 7 1 2 79815 32081
0 32083 5 1 1 32082
0 32084 7 1 2 72722 32083
0 32085 5 1 1 32084
0 32086 7 2 2 79784 78108
0 32087 5 1 1 94678
0 32088 7 1 2 69841 94679
0 32089 5 1 1 32088
0 32090 7 1 2 32085 32089
0 32091 5 1 1 32090
0 32092 7 1 2 85703 32091
0 32093 5 1 1 32092
0 32094 7 1 2 32079 32093
0 32095 5 1 1 32094
0 32096 7 1 2 66712 32095
0 32097 5 1 1 32096
0 32098 7 1 2 32056 32097
0 32099 5 1 1 32098
0 32100 7 1 2 62687 32099
0 32101 5 1 1 32100
0 32102 7 1 2 79045 82909
0 32103 7 1 2 86228 32102
0 32104 5 1 1 32103
0 32105 7 1 2 72723 93578
0 32106 5 1 1 32105
0 32107 7 2 2 68710 72344
0 32108 7 1 2 66713 80754
0 32109 7 1 2 94680 32108
0 32110 5 1 1 32109
0 32111 7 1 2 32106 32110
0 32112 5 1 1 32111
0 32113 7 1 2 66860 75668
0 32114 7 1 2 32112 32113
0 32115 5 1 1 32114
0 32116 7 1 2 32104 32115
0 32117 5 1 1 32116
0 32118 7 1 2 69676 32117
0 32119 5 1 1 32118
0 32120 7 1 2 32101 32119
0 32121 5 1 1 32120
0 32122 7 1 2 65446 32121
0 32123 5 1 1 32122
0 32124 7 1 2 79280 80369
0 32125 5 1 1 32124
0 32126 7 1 2 70977 77163
0 32127 7 1 2 32125 32126
0 32128 5 1 1 32127
0 32129 7 1 2 60550 94436
0 32130 7 1 2 78645 32129
0 32131 5 1 1 32130
0 32132 7 1 2 32128 32131
0 32133 5 1 1 32132
0 32134 7 1 2 78768 32133
0 32135 5 1 1 32134
0 32136 7 2 2 83546 72345
0 32137 7 1 2 72596 88176
0 32138 7 1 2 94682 32137
0 32139 5 1 1 32138
0 32140 7 1 2 32135 32139
0 32141 5 1 1 32140
0 32142 7 1 2 62688 32141
0 32143 5 1 1 32142
0 32144 7 2 2 79461 85452
0 32145 7 1 2 89173 94684
0 32146 5 1 1 32145
0 32147 7 1 2 32143 32146
0 32148 5 1 1 32147
0 32149 7 1 2 62340 32148
0 32150 5 1 1 32149
0 32151 7 2 2 77238 91440
0 32152 5 2 1 94686
0 32153 7 1 2 72675 94688
0 32154 5 1 1 32153
0 32155 7 1 2 88177 92149
0 32156 7 1 2 32154 32155
0 32157 5 1 1 32156
0 32158 7 1 2 32150 32157
0 32159 5 1 1 32158
0 32160 7 1 2 66861 32159
0 32161 5 1 1 32160
0 32162 7 1 2 32123 32161
0 32163 5 1 1 32162
0 32164 7 1 2 64004 32163
0 32165 5 1 1 32164
0 32166 7 2 2 78993 92277
0 32167 7 1 2 85871 87844
0 32168 7 1 2 94690 32167
0 32169 5 1 1 32168
0 32170 7 1 2 60666 32169
0 32171 7 1 2 32165 32170
0 32172 5 1 1 32171
0 32173 7 1 2 72724 91657
0 32174 5 1 1 32173
0 32175 7 1 2 77836 91856
0 32176 5 1 1 32175
0 32177 7 1 2 91672 32176
0 32178 5 2 1 32177
0 32179 7 1 2 62689 77239
0 32180 7 1 2 94692 32179
0 32181 5 1 1 32180
0 32182 7 1 2 32174 32181
0 32183 5 1 1 32182
0 32184 7 1 2 64298 32183
0 32185 5 1 1 32184
0 32186 7 4 2 65003 65727
0 32187 5 1 1 94694
0 32188 7 1 2 67663 90440
0 32189 5 2 1 32188
0 32190 7 3 2 88825 94698
0 32191 5 1 1 94700
0 32192 7 1 2 32187 32191
0 32193 5 1 1 32192
0 32194 7 1 2 91658 32193
0 32195 5 1 1 32194
0 32196 7 1 2 32185 32195
0 32197 5 1 1 32196
0 32198 7 1 2 61733 32197
0 32199 5 1 1 32198
0 32200 7 1 2 78625 93829
0 32201 5 1 1 32200
0 32202 7 1 2 18578 32201
0 32203 5 1 1 32202
0 32204 7 1 2 62690 32203
0 32205 5 1 1 32204
0 32206 7 1 2 72725 94562
0 32207 5 1 1 32206
0 32208 7 1 2 32205 32207
0 32209 5 1 1 32208
0 32210 7 1 2 80358 32209
0 32211 5 1 1 32210
0 32212 7 1 2 32199 32211
0 32213 5 1 1 32212
0 32214 7 1 2 62341 86097
0 32215 7 1 2 32213 32214
0 32216 5 1 1 32215
0 32217 7 1 2 81186 93440
0 32218 5 1 1 32217
0 32219 7 1 2 84238 32218
0 32220 5 1 1 32219
0 32221 7 1 2 82521 86168
0 32222 7 1 2 32220 32221
0 32223 5 1 1 32222
0 32224 7 1 2 32216 32223
0 32225 5 1 1 32224
0 32226 7 1 2 63770 32225
0 32227 5 1 1 32226
0 32228 7 1 2 84060 87107
0 32229 7 1 2 94673 32228
0 32230 5 1 1 32229
0 32231 7 1 2 75596 85862
0 32232 5 1 1 32231
0 32233 7 1 2 66862 92033
0 32234 5 1 1 32233
0 32235 7 1 2 32232 32234
0 32236 5 1 1 32235
0 32237 7 1 2 72614 89157
0 32238 7 1 2 32236 32237
0 32239 5 1 1 32238
0 32240 7 1 2 32230 32239
0 32241 5 1 1 32240
0 32242 7 1 2 77569 32241
0 32243 5 1 1 32242
0 32244 7 1 2 68389 32243
0 32245 7 1 2 32227 32244
0 32246 5 1 1 32245
0 32247 7 1 2 77147 92000
0 32248 5 1 1 32247
0 32249 7 1 2 22052 32248
0 32250 5 1 1 32249
0 32251 7 1 2 65004 32250
0 32252 5 1 1 32251
0 32253 7 1 2 71224 94664
0 32254 5 1 1 32253
0 32255 7 1 2 72346 94004
0 32256 7 1 2 32254 32255
0 32257 5 1 1 32256
0 32258 7 1 2 32252 32257
0 32259 5 1 1 32258
0 32260 7 1 2 87108 32259
0 32261 5 1 1 32260
0 32262 7 1 2 90453 93627
0 32263 5 1 1 32262
0 32264 7 1 2 86098 94666
0 32265 5 1 1 32264
0 32266 7 1 2 85243 94369
0 32267 5 1 1 32266
0 32268 7 1 2 32265 32267
0 32269 5 1 1 32268
0 32270 7 1 2 72347 32269
0 32271 5 1 1 32270
0 32272 7 1 2 77868 86169
0 32273 7 1 2 78639 32272
0 32274 5 1 1 32273
0 32275 7 1 2 86127 32274
0 32276 7 1 2 32271 32275
0 32277 5 1 1 32276
0 32278 7 1 2 83626 32277
0 32279 5 1 1 32278
0 32280 7 1 2 32263 32279
0 32281 5 1 1 32280
0 32282 7 1 2 81187 32281
0 32283 5 1 1 32282
0 32284 7 1 2 32261 32283
0 32285 5 1 1 32284
0 32286 7 1 2 62691 32285
0 32287 5 1 1 32286
0 32288 7 1 2 84642 91092
0 32289 5 1 1 32288
0 32290 7 1 2 79213 32289
0 32291 5 1 1 32290
0 32292 7 1 2 86170 87086
0 32293 7 1 2 32291 32292
0 32294 5 1 1 32293
0 32295 7 1 2 63498 32294
0 32296 7 1 2 32287 32295
0 32297 5 1 1 32296
0 32298 7 1 2 32246 32297
0 32299 5 1 1 32298
0 32300 7 1 2 65586 32299
0 32301 5 1 1 32300
0 32302 7 1 2 64097 32301
0 32303 7 1 2 32172 32302
0 32304 5 1 1 32303
0 32305 7 1 2 76259 73718
0 32306 5 2 1 32305
0 32307 7 1 2 85876 94640
0 32308 7 1 2 88269 94226
0 32309 7 1 2 32307 32308
0 32310 7 1 2 94703 32309
0 32311 5 1 1 32310
0 32312 7 1 2 32304 32311
0 32313 5 1 1 32312
0 32314 7 1 2 32022 32313
0 32315 5 1 1 32314
0 32316 7 1 2 94471 94683
0 32317 5 1 1 32316
0 32318 7 1 2 66714 80565
0 32319 7 1 2 91905 32318
0 32320 5 1 1 32319
0 32321 7 1 2 32317 32320
0 32322 5 1 1 32321
0 32323 7 1 2 91651 32322
0 32324 5 1 1 32323
0 32325 7 1 2 61734 94693
0 32326 5 1 1 32325
0 32327 7 1 2 80359 85264
0 32328 5 1 1 32327
0 32329 7 1 2 32326 32328
0 32330 5 1 1 32329
0 32331 7 1 2 66312 32330
0 32332 5 1 1 32331
0 32333 7 1 2 80566 86568
0 32334 5 1 1 32333
0 32335 7 1 2 32332 32334
0 32336 5 1 1 32335
0 32337 7 1 2 73697 78769
0 32338 7 1 2 32336 32337
0 32339 5 1 1 32338
0 32340 7 1 2 32324 32339
0 32341 5 1 1 32340
0 32342 7 1 2 62130 32341
0 32343 5 1 1 32342
0 32344 7 2 2 75669 85327
0 32345 5 1 1 94705
0 32346 7 1 2 80659 77297
0 32347 7 1 2 94706 32346
0 32348 5 1 1 32347
0 32349 7 1 2 32343 32348
0 32350 5 1 1 32349
0 32351 7 1 2 64005 32350
0 32352 5 1 1 32351
0 32353 7 1 2 90736 94421
0 32354 7 1 2 94691 32353
0 32355 5 1 1 32354
0 32356 7 1 2 32352 32355
0 32357 5 1 1 32356
0 32358 7 1 2 86785 32357
0 32359 5 1 1 32358
0 32360 7 1 2 83547 87003
0 32361 5 1 1 32360
0 32362 7 1 2 81271 87881
0 32363 7 1 2 88266 32362
0 32364 7 1 2 92836 32363
0 32365 5 1 1 32364
0 32366 7 1 2 32361 32365
0 32367 5 1 1 32366
0 32368 7 1 2 70884 32367
0 32369 5 1 1 32368
0 32370 7 1 2 79785 70890
0 32371 7 1 2 92786 32370
0 32372 5 1 1 32371
0 32373 7 1 2 32369 32372
0 32374 5 1 1 32373
0 32375 7 1 2 71456 32374
0 32376 5 1 1 32375
0 32377 7 1 2 76745 72348
0 32378 5 2 1 32377
0 32379 7 1 2 66041 79394
0 32380 5 1 1 32379
0 32381 7 1 2 94707 32380
0 32382 5 1 1 32381
0 32383 7 2 2 68711 80738
0 32384 7 1 2 69842 87640
0 32385 7 1 2 94709 32384
0 32386 7 1 2 32382 32385
0 32387 5 1 1 32386
0 32388 7 1 2 32376 32387
0 32389 5 1 1 32388
0 32390 7 1 2 64006 32389
0 32391 5 1 1 32390
0 32392 7 1 2 77739 93801
0 32393 5 1 1 32392
0 32394 7 1 2 75145 81188
0 32395 5 1 1 32394
0 32396 7 1 2 32393 32395
0 32397 5 1 1 32396
0 32398 7 1 2 86576 94089
0 32399 7 1 2 32397 32398
0 32400 5 1 1 32399
0 32401 7 1 2 32391 32400
0 32402 7 1 2 32359 32401
0 32403 5 1 1 32402
0 32404 7 1 2 64098 32403
0 32405 5 1 1 32404
0 32406 7 2 2 85368 94227
0 32407 7 1 2 87993 94711
0 32408 7 1 2 94657 32407
0 32409 5 1 1 32408
0 32410 7 1 2 32405 32409
0 32411 5 1 1 32410
0 32412 7 1 2 88896 32411
0 32413 5 1 1 32412
0 32414 7 15 2 68712 64099
0 32415 7 1 2 88566 94448
0 32416 5 1 1 32415
0 32417 7 1 2 82522 94139
0 32418 5 1 1 32417
0 32419 7 1 2 69843 93077
0 32420 7 1 2 93408 32419
0 32421 5 1 1 32420
0 32422 7 1 2 32418 32421
0 32423 5 1 1 32422
0 32424 7 1 2 85771 32423
0 32425 5 1 1 32424
0 32426 7 1 2 32416 32425
0 32427 5 1 1 32426
0 32428 7 1 2 87172 32427
0 32429 5 1 1 32428
0 32430 7 1 2 66535 87641
0 32431 7 1 2 88567 32430
0 32432 5 1 1 32431
0 32433 7 1 2 32429 32432
0 32434 5 1 1 32433
0 32435 7 1 2 94713 32434
0 32436 5 1 1 32435
0 32437 7 9 2 68978 87070
0 32438 7 2 2 88019 94728
0 32439 5 1 1 94737
0 32440 7 3 2 63771 94738
0 32441 5 1 1 94739
0 32442 7 1 2 80033 85063
0 32443 7 1 2 89167 32442
0 32444 7 1 2 94740 32443
0 32445 5 1 1 32444
0 32446 7 1 2 32436 32445
0 32447 5 1 1 32446
0 32448 7 1 2 65240 32447
0 32449 5 1 1 32448
0 32450 7 1 2 82523 87004
0 32451 5 1 1 32450
0 32452 7 1 2 93078 94140
0 32453 5 1 1 32452
0 32454 7 1 2 87601 32453
0 32455 5 1 1 32454
0 32456 7 1 2 69844 32455
0 32457 5 1 1 32456
0 32458 7 1 2 74027 83726
0 32459 5 1 1 32458
0 32460 7 1 2 32457 32459
0 32461 5 1 1 32460
0 32462 7 1 2 86786 32461
0 32463 5 1 1 32462
0 32464 7 1 2 32451 32463
0 32465 5 1 1 32464
0 32466 7 3 2 64100 83548
0 32467 7 1 2 83869 94742
0 32468 7 1 2 32465 32467
0 32469 5 1 1 32468
0 32470 7 1 2 32449 32469
0 32471 5 1 1 32470
0 32472 7 1 2 64007 32471
0 32473 5 1 1 32472
0 32474 7 1 2 83701 91919
0 32475 7 1 2 93550 32474
0 32476 5 1 1 32475
0 32477 7 1 2 80421 86385
0 32478 7 1 2 92883 32477
0 32479 5 1 1 32478
0 32480 7 1 2 32476 32479
0 32481 5 1 1 32480
0 32482 7 1 2 65241 32481
0 32483 5 1 1 32482
0 32484 7 2 2 70455 83549
0 32485 7 1 2 75318 79290
0 32486 7 1 2 94418 32485
0 32487 7 1 2 94745 32486
0 32488 7 1 2 85265 32487
0 32489 5 1 1 32488
0 32490 7 1 2 32483 32489
0 32491 5 1 1 32490
0 32492 7 29 2 68885 64101
0 32493 7 1 2 94481 94747
0 32494 7 1 2 32491 32493
0 32495 5 1 1 32494
0 32496 7 1 2 32473 32495
0 32497 5 1 1 32496
0 32498 7 1 2 77816 32497
0 32499 5 1 1 32498
0 32500 7 1 2 77996 86959
0 32501 5 1 1 32500
0 32502 7 1 2 60160 170
0 32503 5 1 1 32502
0 32504 7 1 2 75670 32503
0 32505 5 1 1 32504
0 32506 7 1 2 66042 82524
0 32507 5 1 1 32506
0 32508 7 1 2 83777 32507
0 32509 5 1 1 32508
0 32510 7 1 2 79786 32509
0 32511 5 1 1 32510
0 32512 7 1 2 32505 32511
0 32513 5 1 1 32512
0 32514 7 1 2 94499 32513
0 32515 5 1 1 32514
0 32516 7 1 2 22812 93542
0 32517 5 1 1 32516
0 32518 7 1 2 65242 32517
0 32519 5 1 1 32518
0 32520 7 1 2 32519 94659
0 32521 5 1 1 32520
0 32522 7 1 2 87392 32521
0 32523 5 1 1 32522
0 32524 7 2 2 86715 92667
0 32525 5 1 1 94776
0 32526 7 1 2 80034 93330
0 32527 7 1 2 94777 32526
0 32528 5 1 1 32527
0 32529 7 1 2 32523 32528
0 32530 5 1 1 32529
0 32531 7 1 2 72597 32530
0 32532 5 1 1 32531
0 32533 7 2 2 78770 86171
0 32534 7 1 2 94642 94778
0 32535 5 1 1 32534
0 32536 7 1 2 87393 90242
0 32537 7 1 2 94587 32536
0 32538 5 1 1 32537
0 32539 7 1 2 32535 32538
0 32540 5 1 1 32539
0 32541 7 1 2 75597 32540
0 32542 5 1 1 32541
0 32543 7 1 2 32532 32542
0 32544 5 1 1 32543
0 32545 7 1 2 81189 32544
0 32546 5 1 1 32545
0 32547 7 1 2 32515 32546
0 32548 5 1 1 32547
0 32549 7 1 2 62692 32548
0 32550 5 1 1 32549
0 32551 7 1 2 77298 94695
0 32552 7 1 2 94746 32551
0 32553 5 1 1 32552
0 32554 7 1 2 78791 32553
0 32555 5 1 1 32554
0 32556 7 1 2 84223 32555
0 32557 5 1 1 32556
0 32558 7 1 2 79462 88739
0 32559 5 1 1 32558
0 32560 7 1 2 32557 32559
0 32561 5 1 1 32560
0 32562 7 1 2 88067 32561
0 32563 5 1 1 32562
0 32564 7 1 2 87420 88256
0 32565 5 1 1 32564
0 32566 7 1 2 80198 86372
0 32567 5 1 1 32566
0 32568 7 1 2 32565 32567
0 32569 5 1 1 32568
0 32570 7 1 2 65587 32569
0 32571 5 1 1 32570
0 32572 7 1 2 80199 94057
0 32573 5 1 1 32572
0 32574 7 1 2 32571 32573
0 32575 5 1 1 32574
0 32576 7 1 2 94492 32575
0 32577 5 1 1 32576
0 32578 7 1 2 77869 90110
0 32579 7 1 2 87506 32578
0 32580 5 1 1 32579
0 32581 7 1 2 32577 32580
0 32582 5 1 1 32581
0 32583 7 1 2 66536 32582
0 32584 5 1 1 32583
0 32585 7 1 2 7704 88241
0 32586 5 1 1 32585
0 32587 7 1 2 65447 90740
0 32588 7 1 2 87394 32587
0 32589 7 1 2 32586 32588
0 32590 5 1 1 32589
0 32591 7 1 2 32584 32590
0 32592 5 1 1 32591
0 32593 7 1 2 69677 32592
0 32594 5 1 1 32593
0 32595 7 1 2 32563 32594
0 32596 7 1 2 32550 32595
0 32597 5 1 1 32596
0 32598 7 1 2 64102 32597
0 32599 5 1 1 32598
0 32600 7 4 2 65588 66537
0 32601 7 2 2 81316 94780
0 32602 7 1 2 80755 81742
0 32603 7 1 2 73698 32602
0 32604 7 1 2 94784 32603
0 32605 7 1 2 94234 32604
0 32606 5 1 1 32605
0 32607 7 1 2 32599 32606
0 32608 5 1 1 32607
0 32609 7 1 2 32501 32608
0 32610 5 1 1 32609
0 32611 7 1 2 32499 32610
0 32612 7 1 2 32413 32611
0 32613 7 1 2 32315 32612
0 32614 7 1 2 32020 32613
0 32615 7 1 2 31893 32614
0 32616 7 1 2 31068 32615
0 32617 7 2 2 29649 32616
0 32618 5 1 1 94786
0 32619 7 1 2 84187 78957
0 32620 5 1 1 32619
0 32621 7 1 2 77321 93745
0 32622 5 1 1 32621
0 32623 7 1 2 32620 32622
0 32624 5 1 1 32623
0 32625 7 1 2 64540 32624
0 32626 5 1 1 32625
0 32627 7 2 2 64763 70314
0 32628 7 3 2 82750 94788
0 32629 5 1 1 94790
0 32630 7 1 2 74371 94791
0 32631 5 1 1 32630
0 32632 7 1 2 85461 32631
0 32633 5 1 1 32632
0 32634 7 1 2 63772 32633
0 32635 5 1 1 32634
0 32636 7 1 2 32626 32635
0 32637 5 1 1 32636
0 32638 7 1 2 65883 32637
0 32639 5 1 1 32638
0 32640 7 1 2 7631 85147
0 32641 5 2 1 32640
0 32642 7 1 2 64764 21690
0 32643 7 1 2 94793 32642
0 32644 5 1 1 32643
0 32645 7 1 2 82801 85139
0 32646 5 1 1 32645
0 32647 7 1 2 85475 32646
0 32648 7 1 2 32644 32647
0 32649 5 1 1 32648
0 32650 7 1 2 66538 32649
0 32651 5 1 1 32650
0 32652 7 1 2 32639 32651
0 32653 5 1 1 32652
0 32654 7 1 2 65243 32653
0 32655 5 1 1 32654
0 32656 7 3 2 82111 85045
0 32657 7 1 2 93357 94795
0 32658 7 1 2 82802 32657
0 32659 5 1 1 32658
0 32660 7 1 2 83715 32659
0 32661 5 1 1 32660
0 32662 7 1 2 80491 71494
0 32663 5 3 1 32662
0 32664 7 1 2 63773 94798
0 32665 7 1 2 32661 32664
0 32666 5 1 1 32665
0 32667 7 1 2 32655 32666
0 32668 5 1 1 32667
0 32669 7 1 2 63499 32668
0 32670 5 1 1 32669
0 32671 7 1 2 75598 91195
0 32672 5 1 1 32671
0 32673 7 1 2 81635 90859
0 32674 7 1 2 91857 32673
0 32675 5 1 1 32674
0 32676 7 1 2 32672 32675
0 32677 5 1 1 32676
0 32678 7 1 2 64541 32677
0 32679 5 1 1 32678
0 32680 7 1 2 84636 90433
0 32681 5 1 1 32680
0 32682 7 1 2 32679 32681
0 32683 5 1 1 32682
0 32684 7 1 2 64299 32683
0 32685 5 1 1 32684
0 32686 7 1 2 93546 93822
0 32687 5 1 1 32686
0 32688 7 1 2 32685 32687
0 32689 5 1 1 32688
0 32690 7 1 2 78771 32689
0 32691 5 1 1 32690
0 32692 7 1 2 32670 32691
0 32693 5 1 1 32692
0 32694 7 1 2 78060 32693
0 32695 5 1 1 32694
0 32696 7 2 2 62131 73570
0 32697 5 1 1 94801
0 32698 7 1 2 71795 89362
0 32699 5 1 1 32698
0 32700 7 3 2 32697 32699
0 32701 5 2 1 94803
0 32702 7 1 2 94533 94806
0 32703 5 1 1 32702
0 32704 7 2 2 83472 32703
0 32705 5 1 1 94808
0 32706 7 1 2 68390 32705
0 32707 5 1 1 32706
0 32708 7 1 2 61353 79992
0 32709 5 1 1 32708
0 32710 7 1 2 79787 32709
0 32711 5 1 1 32710
0 32712 7 1 2 32707 32711
0 32713 5 1 1 32712
0 32714 7 1 2 77570 32713
0 32715 5 1 1 32714
0 32716 7 1 2 61354 90863
0 32717 5 2 1 32716
0 32718 7 1 2 77997 75014
0 32719 5 1 1 32718
0 32720 7 2 2 94810 32719
0 32721 7 1 2 94063 94812
0 32722 5 1 1 32721
0 32723 7 1 2 32715 32722
0 32724 5 1 1 32723
0 32725 7 1 2 65448 32724
0 32726 5 1 1 32725
0 32727 7 1 2 72122 79214
0 32728 5 1 1 32727
0 32729 7 1 2 74422 32728
0 32730 5 1 1 32729
0 32731 7 1 2 59903 32730
0 32732 5 1 1 32731
0 32733 7 1 2 77536 89776
0 32734 5 1 1 32733
0 32735 7 1 2 79215 32734
0 32736 5 1 1 32735
0 32737 7 1 2 63500 32736
0 32738 7 1 2 32732 32737
0 32739 5 1 1 32738
0 32740 7 1 2 83685 90434
0 32741 5 1 1 32740
0 32742 7 1 2 12288 32741
0 32743 5 1 1 32742
0 32744 7 1 2 78772 32743
0 32745 5 1 1 32744
0 32746 7 1 2 69068 94669
0 32747 5 1 1 32746
0 32748 7 1 2 90942 32747
0 32749 5 1 1 32748
0 32750 7 1 2 66313 32749
0 32751 5 1 1 32750
0 32752 7 1 2 32745 32751
0 32753 7 1 2 32739 32752
0 32754 5 1 1 32753
0 32755 7 1 2 79138 32754
0 32756 5 1 1 32755
0 32757 7 1 2 32726 32756
0 32758 5 1 1 32757
0 32759 7 1 2 66715 32758
0 32760 5 1 1 32759
0 32761 7 1 2 68886 79354
0 32762 7 1 2 93547 32761
0 32763 5 1 1 32762
0 32764 7 1 2 24529 32763
0 32765 5 1 1 32764
0 32766 7 2 2 64542 32765
0 32767 7 1 2 80035 94814
0 32768 5 1 1 32767
0 32769 7 2 2 60551 92964
0 32770 5 1 1 94816
0 32771 7 1 2 32768 32770
0 32772 5 1 1 32771
0 32773 7 1 2 66716 32772
0 32774 5 1 1 32773
0 32775 7 2 2 64543 77571
0 32776 7 1 2 65449 81120
0 32777 7 1 2 94818 32776
0 32778 5 1 1 32777
0 32779 7 1 2 32774 32778
0 32780 5 1 1 32779
0 32781 7 1 2 65244 32780
0 32782 5 1 1 32781
0 32783 7 1 2 83702 85680
0 32784 7 1 2 94819 32783
0 32785 5 1 1 32784
0 32786 7 1 2 32782 32785
0 32787 5 1 1 32786
0 32788 7 1 2 81569 32787
0 32789 5 1 1 32788
0 32790 7 1 2 32760 32789
0 32791 7 1 2 32695 32790
0 32792 5 1 1 32791
0 32793 7 1 2 63050 32792
0 32794 5 1 1 32793
0 32795 7 1 2 80550 88254
0 32796 5 1 1 32795
0 32797 7 1 2 27954 32796
0 32798 5 1 1 32797
0 32799 7 1 2 65450 32798
0 32800 5 1 1 32799
0 32801 7 1 2 83103 88229
0 32802 7 1 2 88461 32801
0 32803 5 1 1 32802
0 32804 7 1 2 79457 32803
0 32805 5 1 1 32804
0 32806 7 1 2 79139 32805
0 32807 5 1 1 32806
0 32808 7 1 2 32800 32807
0 32809 5 1 1 32808
0 32810 7 1 2 66539 32809
0 32811 5 1 1 32810
0 32812 7 2 2 79788 88462
0 32813 5 1 1 94820
0 32814 7 1 2 85660 94821
0 32815 5 1 1 32814
0 32816 7 1 2 82189 32815
0 32817 5 1 1 32816
0 32818 7 1 2 64008 86422
0 32819 7 1 2 32817 32818
0 32820 5 1 1 32819
0 32821 7 1 2 32811 32820
0 32822 5 1 1 32821
0 32823 7 1 2 66314 32822
0 32824 5 1 1 32823
0 32825 7 1 2 79700 85436
0 32826 7 1 2 94360 32825
0 32827 5 1 1 32826
0 32828 7 1 2 32824 32827
0 32829 5 1 1 32828
0 32830 7 1 2 63774 32829
0 32831 5 1 1 32830
0 32832 7 2 2 83550 87315
0 32833 7 1 2 94472 94822
0 32834 5 1 1 32833
0 32835 7 1 2 32831 32834
0 32836 5 1 1 32835
0 32837 7 1 2 64765 32836
0 32838 5 1 1 32837
0 32839 7 1 2 79140 92884
0 32840 5 1 1 32839
0 32841 7 1 2 80518 81981
0 32842 5 1 1 32841
0 32843 7 1 2 32840 32842
0 32844 5 1 1 32843
0 32845 7 1 2 81299 79379
0 32846 7 1 2 32844 32845
0 32847 5 1 1 32846
0 32848 7 1 2 32838 32847
0 32849 5 1 1 32848
0 32850 7 1 2 69255 32849
0 32851 5 1 1 32850
0 32852 7 1 2 89969 93832
0 32853 5 1 1 32852
0 32854 7 1 2 61565 32853
0 32855 5 1 1 32854
0 32856 7 1 2 89932 94534
0 32857 7 1 2 80451 32856
0 32858 5 1 1 32857
0 32859 7 1 2 32855 32858
0 32860 5 1 1 32859
0 32861 7 1 2 66717 32860
0 32862 5 1 1 32861
0 32863 7 5 2 63775 81989
0 32864 5 1 1 94824
0 32865 7 1 2 80005 88771
0 32866 5 2 1 32865
0 32867 7 1 2 83468 94829
0 32868 5 1 1 32867
0 32869 7 1 2 75319 32868
0 32870 5 1 1 32869
0 32871 7 1 2 94825 32870
0 32872 5 1 1 32871
0 32873 7 1 2 32862 32872
0 32874 5 1 1 32873
0 32875 7 1 2 65451 32874
0 32876 5 1 1 32875
0 32877 7 1 2 66315 94830
0 32878 5 1 1 32877
0 32879 7 1 2 60366 32878
0 32880 5 1 1 32879
0 32881 7 1 2 94685 32880
0 32882 5 1 1 32881
0 32883 7 1 2 32876 32882
0 32884 5 1 1 32883
0 32885 7 1 2 64009 32884
0 32886 5 1 1 32885
0 32887 7 1 2 79627 93848
0 32888 7 1 2 94796 32887
0 32889 7 1 2 94361 32888
0 32890 5 1 1 32889
0 32891 7 1 2 61875 32890
0 32892 7 1 2 32886 32891
0 32893 7 1 2 32851 32892
0 32894 7 1 2 32794 32893
0 32895 5 1 1 32894
0 32896 7 2 2 69069 73874
0 32897 5 2 1 94831
0 32898 7 1 2 82384 94833
0 32899 5 2 1 32898
0 32900 7 1 2 69845 94835
0 32901 5 1 1 32900
0 32902 7 1 2 84118 93104
0 32903 5 1 1 32902
0 32904 7 1 2 63051 32903
0 32905 5 1 1 32904
0 32906 7 1 2 32901 32905
0 32907 5 1 1 32906
0 32908 7 1 2 66316 32907
0 32909 5 1 1 32908
0 32910 7 2 2 82680 84404
0 32911 5 1 1 94837
0 32912 7 1 2 75974 94838
0 32913 5 1 1 32912
0 32914 7 1 2 32909 32913
0 32915 5 1 1 32914
0 32916 7 1 2 75599 32915
0 32917 5 1 1 32916
0 32918 7 1 2 75222 15909
0 32919 5 1 1 32918
0 32920 7 1 2 68391 32919
0 32921 7 1 2 32917 32920
0 32922 5 1 1 32921
0 32923 7 2 2 61355 74472
0 32924 5 1 1 94839
0 32925 7 1 2 82373 32924
0 32926 5 1 1 32925
0 32927 7 1 2 69846 85251
0 32928 5 1 1 32927
0 32929 7 1 2 87615 32928
0 32930 5 2 1 32929
0 32931 7 1 2 71796 94841
0 32932 5 1 1 32931
0 32933 7 2 2 82326 78461
0 32934 5 1 1 94843
0 32935 7 1 2 63052 32934
0 32936 5 1 1 32935
0 32937 7 1 2 66317 74510
0 32938 5 1 1 32937
0 32939 7 1 2 32936 32938
0 32940 7 1 2 32932 32939
0 32941 5 1 1 32940
0 32942 7 1 2 64766 32941
0 32943 5 1 1 32942
0 32944 7 1 2 32926 32943
0 32945 5 1 1 32944
0 32946 7 1 2 61566 32945
0 32947 5 1 1 32946
0 32948 7 1 2 81903 91112
0 32949 7 1 2 85998 32948
0 32950 5 1 1 32949
0 32951 7 1 2 63501 32950
0 32952 7 1 2 32947 32951
0 32953 5 1 1 32952
0 32954 7 1 2 32922 32953
0 32955 5 1 1 32954
0 32956 7 1 2 71797 86048
0 32957 5 1 1 32956
0 32958 7 1 2 78034 86836
0 32959 5 1 1 32958
0 32960 7 1 2 32957 32959
0 32961 5 1 1 32960
0 32962 7 1 2 68392 32961
0 32963 5 1 1 32962
0 32964 7 1 2 71011 91114
0 32965 5 1 1 32964
0 32966 7 1 2 32963 32965
0 32967 5 1 1 32966
0 32968 7 1 2 69678 32967
0 32969 5 1 1 32968
0 32970 7 1 2 32955 32969
0 32971 5 1 1 32970
0 32972 7 1 2 63776 32971
0 32973 5 1 1 32972
0 32974 7 1 2 82056 88772
0 32975 7 1 2 94804 32974
0 32976 5 1 1 32975
0 32977 7 1 2 86037 92595
0 32978 7 1 2 32976 32977
0 32979 5 1 1 32978
0 32980 7 1 2 32973 32979
0 32981 5 1 1 32980
0 32982 7 1 2 66718 32981
0 32983 5 1 1 32982
0 32984 7 1 2 64767 94842
0 32985 5 1 1 32984
0 32986 7 1 2 78597 32985
0 32987 5 1 1 32986
0 32988 7 1 2 71798 32987
0 32989 5 1 1 32988
0 32990 7 1 2 77331 82112
0 32991 5 1 1 32990
0 32992 7 1 2 73016 77998
0 32993 5 1 1 32992
0 32994 7 1 2 90655 32993
0 32995 5 1 1 32994
0 32996 7 2 2 73571 70493
0 32997 5 1 1 94845
0 32998 7 1 2 69847 94846
0 32999 5 1 1 32998
0 33000 7 1 2 32995 32999
0 33001 5 1 1 33000
0 33002 7 1 2 63053 33001
0 33003 5 1 1 33002
0 33004 7 1 2 32991 33003
0 33005 7 1 2 32989 33004
0 33006 5 2 1 33005
0 33007 7 1 2 79046 79343
0 33008 7 1 2 94847 33007
0 33009 5 1 1 33008
0 33010 7 1 2 60552 33009
0 33011 7 1 2 32983 33010
0 33012 5 1 1 33011
0 33013 7 1 2 79281 89621
0 33014 5 1 1 33013
0 33015 7 1 2 59904 72459
0 33016 5 1 1 33015
0 33017 7 1 2 33014 33016
0 33018 5 1 1 33017
0 33019 7 1 2 73893 85252
0 33020 5 1 1 33019
0 33021 7 1 2 85569 33020
0 33022 5 1 1 33021
0 33023 7 1 2 65728 33022
0 33024 5 1 1 33023
0 33025 7 1 2 2503 33024
0 33026 5 1 1 33025
0 33027 7 1 2 64300 33026
0 33028 5 1 1 33027
0 33029 7 1 2 72123 82476
0 33030 5 1 1 33029
0 33031 7 1 2 66318 33030
0 33032 5 1 1 33031
0 33033 7 1 2 93819 33032
0 33034 5 1 1 33033
0 33035 7 1 2 63054 33034
0 33036 5 1 1 33035
0 33037 7 1 2 33028 33036
0 33038 5 1 1 33037
0 33039 7 1 2 61735 75600
0 33040 7 1 2 33038 33039
0 33041 5 1 1 33040
0 33042 7 1 2 33018 33041
0 33043 5 1 1 33042
0 33044 7 1 2 63777 33043
0 33045 5 1 1 33044
0 33046 7 4 2 61736 84668
0 33047 7 1 2 63055 94849
0 33048 5 1 1 33047
0 33049 7 1 2 92435 33048
0 33050 5 1 1 33049
0 33051 7 1 2 73227 33050
0 33052 5 1 1 33051
0 33053 7 2 2 84546 93590
0 33054 5 1 1 94853
0 33055 7 1 2 78598 94854
0 33056 5 1 1 33055
0 33057 7 1 2 63056 84547
0 33058 5 1 1 33057
0 33059 7 1 2 86024 33058
0 33060 7 1 2 33056 33059
0 33061 5 1 1 33060
0 33062 7 1 2 33052 33061
0 33063 5 1 1 33062
0 33064 7 1 2 62342 33063
0 33065 5 1 1 33064
0 33066 7 1 2 78599 91327
0 33067 5 1 1 33066
0 33068 7 1 2 70315 33067
0 33069 5 1 1 33068
0 33070 7 4 2 65729 75422
0 33071 5 2 1 94855
0 33072 7 1 2 94132 94859
0 33073 7 1 2 33069 33072
0 33074 5 1 1 33073
0 33075 7 1 2 84482 33074
0 33076 5 1 1 33075
0 33077 7 1 2 33065 33076
0 33078 5 1 1 33077
0 33079 7 1 2 65245 33078
0 33080 5 1 1 33079
0 33081 7 1 2 78348 89619
0 33082 5 1 1 33081
0 33083 7 1 2 74641 91411
0 33084 7 1 2 92714 33083
0 33085 5 1 1 33084
0 33086 7 1 2 33082 33085
0 33087 5 1 1 33086
0 33088 7 1 2 63778 33087
0 33089 5 1 1 33088
0 33090 7 1 2 33080 33089
0 33091 5 1 1 33090
0 33092 7 1 2 71799 33091
0 33093 5 1 1 33092
0 33094 7 1 2 68030 90654
0 33095 7 1 2 32997 33094
0 33096 5 1 1 33095
0 33097 7 1 2 80999 83447
0 33098 7 1 2 78717 33097
0 33099 7 1 2 33096 33098
0 33100 5 1 1 33099
0 33101 7 1 2 33093 33100
0 33102 7 1 2 33045 33101
0 33103 5 1 1 33102
0 33104 7 1 2 68393 33103
0 33105 5 1 1 33104
0 33106 7 1 2 61567 94848
0 33107 5 1 1 33106
0 33108 7 1 2 74411 83245
0 33109 5 1 1 33108
0 33110 7 1 2 91115 33109
0 33111 5 1 1 33110
0 33112 7 1 2 33107 33111
0 33113 5 1 1 33112
0 33114 7 1 2 84483 33113
0 33115 5 1 1 33114
0 33116 7 1 2 82385 89628
0 33117 7 1 2 86509 33116
0 33118 5 1 1 33117
0 33119 7 1 2 64768 25701
0 33120 5 1 1 33119
0 33121 7 1 2 64301 80068
0 33122 5 1 1 33121
0 33123 7 1 2 33120 33122
0 33124 7 1 2 80065 33123
0 33125 5 1 1 33124
0 33126 7 1 2 79263 86038
0 33127 7 1 2 33125 33126
0 33128 5 1 1 33127
0 33129 7 1 2 33118 33128
0 33130 5 1 1 33129
0 33131 7 2 2 61356 85079
0 33132 5 1 1 94861
0 33133 7 1 2 68031 79995
0 33134 7 1 2 94862 33133
0 33135 5 1 1 33134
0 33136 7 1 2 68713 33135
0 33137 7 1 2 33130 33136
0 33138 5 1 1 33137
0 33139 7 1 2 33115 33138
0 33140 5 1 1 33139
0 33141 7 1 2 63502 33140
0 33142 5 1 1 33141
0 33143 7 1 2 65452 33142
0 33144 7 1 2 33105 33143
0 33145 5 1 1 33144
0 33146 7 1 2 68887 33145
0 33147 7 1 2 33012 33146
0 33148 5 1 1 33147
0 33149 7 1 2 9390 94809
0 33150 5 1 1 33149
0 33151 7 1 2 68394 33150
0 33152 5 1 1 33151
0 33153 7 1 2 79789 33132
0 33154 5 1 1 33153
0 33155 7 1 2 33152 33154
0 33156 5 1 1 33155
0 33157 7 1 2 63057 33156
0 33158 5 1 1 33157
0 33159 7 1 2 66319 84988
0 33160 5 1 1 33159
0 33161 7 1 2 86680 33160
0 33162 5 1 1 33161
0 33163 7 1 2 79998 33162
0 33164 5 1 1 33163
0 33165 7 1 2 82051 88311
0 33166 5 1 1 33165
0 33167 7 1 2 79816 33166
0 33168 5 1 1 33167
0 33169 7 1 2 65246 33168
0 33170 5 1 1 33169
0 33171 7 1 2 33164 33170
0 33172 7 1 2 33158 33171
0 33173 5 1 1 33172
0 33174 7 1 2 68714 33173
0 33175 5 1 1 33174
0 33176 7 1 2 94616 33175
0 33177 5 1 1 33176
0 33178 7 1 2 81758 33177
0 33179 5 1 1 33178
0 33180 7 1 2 66863 33179
0 33181 7 1 2 33148 33180
0 33182 5 1 1 33181
0 33183 7 1 2 32895 33182
0 33184 5 1 1 33183
0 33185 7 1 2 65589 33184
0 33186 5 1 1 33185
0 33187 7 1 2 72598 86033
0 33188 5 1 1 33187
0 33189 7 1 2 8090 85114
0 33190 5 1 1 33189
0 33191 7 1 2 69679 33190
0 33192 5 1 1 33191
0 33193 7 1 2 33188 33192
0 33194 5 1 1 33193
0 33195 7 1 2 63503 33194
0 33196 5 1 1 33195
0 33197 7 1 2 83795 79579
0 33198 5 1 1 33197
0 33199 7 1 2 33196 33198
0 33200 5 1 1 33199
0 33201 7 1 2 65247 33200
0 33202 5 1 1 33201
0 33203 7 1 2 82803 93514
0 33204 5 1 1 33203
0 33205 7 1 2 33202 33204
0 33206 5 1 1 33205
0 33207 7 1 2 69070 33206
0 33208 5 1 1 33207
0 33209 7 1 2 26117 33208
0 33210 5 1 1 33209
0 33211 7 1 2 64769 33210
0 33212 5 1 1 33211
0 33213 7 1 2 80036 91255
0 33214 7 1 2 94543 33213
0 33215 5 1 1 33214
0 33216 7 1 2 33212 33215
0 33217 5 1 1 33216
0 33218 7 1 2 79711 33217
0 33219 5 1 1 33218
0 33220 7 1 2 81650 82386
0 33221 5 1 1 33220
0 33222 7 1 2 94538 33221
0 33223 5 1 1 33222
0 33224 7 1 2 69848 86676
0 33225 5 1 1 33224
0 33226 7 1 2 33223 33225
0 33227 5 1 1 33226
0 33228 7 1 2 73572 33227
0 33229 5 1 1 33228
0 33230 7 1 2 79790 85993
0 33231 5 1 1 33230
0 33232 7 1 2 64770 82951
0 33233 5 1 1 33232
0 33234 7 1 2 90969 33233
0 33235 5 1 1 33234
0 33236 7 1 2 73522 33235
0 33237 5 1 1 33236
0 33238 7 1 2 78600 33237
0 33239 5 1 1 33238
0 33240 7 1 2 75671 33239
0 33241 5 1 1 33240
0 33242 7 1 2 33231 33241
0 33243 7 1 2 33229 33242
0 33244 5 1 1 33243
0 33245 7 1 2 68715 33244
0 33246 5 1 1 33245
0 33247 7 1 2 94617 33246
0 33248 5 1 1 33247
0 33249 7 1 2 66864 33248
0 33250 5 1 1 33249
0 33251 7 1 2 33219 33250
0 33252 5 1 1 33251
0 33253 7 1 2 64010 33252
0 33254 5 1 1 33253
0 33255 7 1 2 63058 94813
0 33256 5 1 1 33255
0 33257 7 1 2 78610 93909
0 33258 5 1 1 33257
0 33259 7 1 2 33256 33258
0 33260 5 1 1 33259
0 33261 7 1 2 93628 93732
0 33262 7 1 2 33260 33261
0 33263 5 1 1 33262
0 33264 7 1 2 33254 33263
0 33265 5 1 1 33264
0 33266 7 1 2 66719 33265
0 33267 5 1 1 33266
0 33268 7 1 2 86677 94799
0 33269 5 1 1 33268
0 33270 7 1 2 63059 71457
0 33271 5 1 1 33270
0 33272 7 1 2 77999 33271
0 33273 5 1 1 33272
0 33274 7 1 2 75601 33273
0 33275 5 1 1 33274
0 33276 7 1 2 94051 33275
0 33277 5 1 1 33276
0 33278 7 1 2 64544 33277
0 33279 5 1 1 33278
0 33280 7 1 2 86958 94568
0 33281 5 1 1 33280
0 33282 7 1 2 75320 33281
0 33283 7 1 2 33279 33282
0 33284 5 1 1 33283
0 33285 7 1 2 68395 33284
0 33286 5 1 1 33285
0 33287 7 1 2 33269 33286
0 33288 5 1 1 33287
0 33289 7 1 2 63779 33288
0 33290 5 1 1 33289
0 33291 7 1 2 90940 90964
0 33292 5 1 1 33291
0 33293 7 1 2 94602 33292
0 33294 5 1 1 33293
0 33295 7 1 2 64302 75602
0 33296 7 1 2 33294 33295
0 33297 5 1 1 33296
0 33298 7 1 2 81636 94671
0 33299 5 1 1 33298
0 33300 7 1 2 33297 33299
0 33301 5 1 1 33300
0 33302 7 1 2 73573 33301
0 33303 5 1 1 33302
0 33304 7 1 2 18122 33303
0 33305 7 1 2 33290 33304
0 33306 5 1 1 33305
0 33307 7 1 2 64011 86973
0 33308 7 1 2 33306 33307
0 33309 5 1 1 33308
0 33310 7 1 2 33267 33309
0 33311 5 1 1 33310
0 33312 7 1 2 65453 33311
0 33313 5 1 1 33312
0 33314 7 1 2 94345 94624
0 33315 5 1 1 33314
0 33316 7 3 2 63060 71322
0 33317 5 3 1 94863
0 33318 7 1 2 87972 94864
0 33319 7 1 2 93657 33318
0 33320 5 1 1 33319
0 33321 7 1 2 33315 33320
0 33322 5 1 1 33321
0 33323 7 1 2 66320 33322
0 33324 5 1 1 33323
0 33325 7 1 2 94106 94424
0 33326 5 1 1 33325
0 33327 7 1 2 33324 33326
0 33328 5 1 1 33327
0 33329 7 1 2 63780 33328
0 33330 5 1 1 33329
0 33331 7 1 2 83551 87664
0 33332 7 1 2 94473 33331
0 33333 5 1 1 33332
0 33334 7 1 2 33330 33333
0 33335 5 1 1 33334
0 33336 7 1 2 64771 33335
0 33337 5 1 1 33336
0 33338 7 2 2 86210 94381
0 33339 5 1 1 94869
0 33340 7 1 2 69680 94870
0 33341 5 1 1 33340
0 33342 7 1 2 72574 33341
0 33343 5 1 1 33342
0 33344 7 5 2 63061 90141
0 33345 5 1 1 94871
0 33346 7 1 2 66865 94872
0 33347 5 1 1 33346
0 33348 7 1 2 33339 33347
0 33349 5 1 1 33348
0 33350 7 1 2 63781 81300
0 33351 7 1 2 33349 33350
0 33352 7 1 2 33343 33351
0 33353 5 1 1 33352
0 33354 7 1 2 33337 33353
0 33355 5 1 1 33354
0 33356 7 1 2 64012 33355
0 33357 5 1 1 33356
0 33358 7 1 2 87560 18370
0 33359 5 1 1 33358
0 33360 7 1 2 64772 33359
0 33361 5 1 1 33360
0 33362 7 1 2 78601 33361
0 33363 5 1 1 33362
0 33364 7 1 2 79701 86577
0 33365 7 1 2 33363 33364
0 33366 5 1 1 33365
0 33367 7 1 2 33357 33366
0 33368 5 1 1 33367
0 33369 7 1 2 69256 33368
0 33370 5 1 1 33369
0 33371 7 7 2 66866 64013
0 33372 7 1 2 77610 74467
0 33373 5 1 1 33372
0 33374 7 1 2 79817 33373
0 33375 5 1 1 33374
0 33376 7 1 2 64773 33375
0 33377 5 1 1 33376
0 33378 7 1 2 71470 87973
0 33379 7 1 2 78631 33378
0 33380 7 1 2 4238 33379
0 33381 5 1 1 33380
0 33382 7 1 2 68396 90889
0 33383 5 1 1 33382
0 33384 7 1 2 80050 33383
0 33385 7 1 2 33381 33384
0 33386 5 1 1 33385
0 33387 7 1 2 33377 33386
0 33388 5 1 1 33387
0 33389 7 1 2 79380 33388
0 33390 5 1 1 33389
0 33391 7 2 2 69681 73574
0 33392 7 1 2 77537 89686
0 33393 5 1 1 33392
0 33394 7 1 2 94603 33393
0 33395 5 1 1 33394
0 33396 7 1 2 94883 33395
0 33397 5 1 1 33396
0 33398 7 1 2 83686 82374
0 33399 5 1 1 33398
0 33400 7 1 2 26586 33399
0 33401 5 1 1 33400
0 33402 7 1 2 78773 33401
0 33403 5 1 1 33402
0 33404 7 1 2 60367 33403
0 33405 5 1 1 33404
0 33406 7 1 2 94622 33405
0 33407 5 1 1 33406
0 33408 7 1 2 33397 33407
0 33409 5 1 1 33408
0 33410 7 1 2 66540 33409
0 33411 5 1 1 33410
0 33412 7 1 2 33390 33411
0 33413 5 1 1 33412
0 33414 7 1 2 66720 33413
0 33415 5 1 1 33414
0 33416 7 1 2 83232 82804
0 33417 5 1 1 33416
0 33418 7 1 2 60368 33417
0 33419 5 1 1 33418
0 33420 7 1 2 79488 92508
0 33421 7 1 2 94800 33420
0 33422 7 1 2 33419 33421
0 33423 5 1 1 33422
0 33424 7 1 2 33415 33423
0 33425 5 1 1 33424
0 33426 7 1 2 60553 33425
0 33427 5 1 1 33426
0 33428 7 1 2 64545 85890
0 33429 5 1 1 33428
0 33430 7 1 2 32813 33429
0 33431 5 1 1 33430
0 33432 7 2 2 65248 84484
0 33433 5 1 1 94885
0 33434 7 1 2 78035 85824
0 33435 7 1 2 94886 33434
0 33436 7 1 2 33431 33435
0 33437 5 1 1 33436
0 33438 7 1 2 33427 33437
0 33439 5 1 1 33438
0 33440 7 1 2 94876 33439
0 33441 5 1 1 33440
0 33442 7 1 2 87665 94815
0 33443 5 1 1 33442
0 33444 7 1 2 80519 93928
0 33445 5 1 1 33444
0 33446 7 1 2 33443 33445
0 33447 5 1 1 33446
0 33448 7 1 2 80037 33447
0 33449 5 1 1 33448
0 33450 7 1 2 87666 94817
0 33451 5 1 1 33450
0 33452 7 1 2 33449 33451
0 33453 5 1 1 33452
0 33454 7 1 2 66721 33453
0 33455 5 1 1 33454
0 33456 7 1 2 64546 94877
0 33457 7 2 2 91157 33456
0 33458 7 1 2 94629 94887
0 33459 5 1 1 33458
0 33460 7 1 2 33455 33459
0 33461 5 1 1 33460
0 33462 7 1 2 65249 33461
0 33463 5 1 1 33462
0 33464 7 1 2 87597 94888
0 33465 5 1 1 33464
0 33466 7 1 2 33463 33465
0 33467 5 1 1 33466
0 33468 7 1 2 81570 33467
0 33469 5 1 1 33468
0 33470 7 1 2 60667 33469
0 33471 7 1 2 33441 33470
0 33472 7 1 2 33370 33471
0 33473 7 1 2 33313 33472
0 33474 5 1 1 33473
0 33475 7 2 2 33186 33474
0 33476 7 1 2 64103 94889
0 33477 5 1 1 33476
0 33478 7 1 2 73575 71323
0 33479 5 1 1 33478
0 33480 7 1 2 74597 33479
0 33481 5 1 1 33480
0 33482 7 2 2 66541 78710
0 33483 7 1 2 94246 94891
0 33484 7 1 2 94235 33483
0 33485 7 2 2 33481 33484
0 33486 5 1 1 94893
0 33487 7 1 2 33477 33486
0 33488 5 1 1 33487
0 33489 7 1 2 73837 33488
0 33490 5 1 1 33489
0 33491 7 2 2 69988 87395
0 33492 5 1 1 94895
0 33493 7 1 2 71563 94896
0 33494 5 1 1 33493
0 33495 7 3 2 86172 94242
0 33496 5 1 1 94897
0 33497 7 1 2 86517 91649
0 33498 5 3 1 33497
0 33499 7 1 2 94898 94900
0 33500 5 1 1 33499
0 33501 7 1 2 33494 33500
0 33502 5 1 1 33501
0 33503 7 1 2 63062 33502
0 33504 5 1 1 33503
0 33505 7 2 2 79123 88068
0 33506 7 1 2 69989 94903
0 33507 5 1 1 33506
0 33508 7 1 2 33504 33507
0 33509 5 1 1 33508
0 33510 7 1 2 94141 33509
0 33511 5 1 1 33510
0 33512 7 3 2 71564 88069
0 33513 5 1 1 94905
0 33514 7 1 2 84381 94906
0 33515 5 1 1 33514
0 33516 7 1 2 87396 91218
0 33517 5 1 1 33516
0 33518 7 1 2 33515 33517
0 33519 5 1 1 33518
0 33520 7 1 2 66722 33519
0 33521 5 1 1 33520
0 33522 7 1 2 87316 87642
0 33523 5 1 1 33522
0 33524 7 1 2 33521 33523
0 33525 5 1 1 33524
0 33526 7 1 2 61568 33525
0 33527 5 1 1 33526
0 33528 7 2 2 63063 87397
0 33529 5 1 1 94908
0 33530 7 6 2 65005 81728
0 33531 7 1 2 81773 94910
0 33532 7 1 2 94909 33531
0 33533 5 1 1 33532
0 33534 7 1 2 33527 33533
0 33535 5 1 1 33534
0 33536 7 1 2 69990 33535
0 33537 5 1 1 33536
0 33538 7 1 2 33511 33537
0 33539 5 1 1 33538
0 33540 7 1 2 65884 33539
0 33541 5 1 1 33540
0 33542 7 2 2 66542 94243
0 33543 7 4 2 69849 86315
0 33544 7 1 2 91125 94918
0 33545 7 1 2 94916 33544
0 33546 7 1 2 88056 33545
0 33547 5 1 1 33546
0 33548 7 1 2 33541 33547
0 33549 5 1 1 33548
0 33550 7 1 2 64547 33549
0 33551 5 1 1 33550
0 33552 7 2 2 70809 93278
0 33553 7 1 2 84224 94485
0 33554 7 1 2 94922 33553
0 33555 5 1 1 33554
0 33556 7 1 2 33551 33555
0 33557 5 1 1 33556
0 33558 7 1 2 64774 33557
0 33559 5 1 1 33558
0 33560 7 1 2 82771 82555
0 33561 5 2 1 33560
0 33562 7 1 2 86787 94474
0 33563 5 1 1 33562
0 33564 7 1 2 10616 33563
0 33565 5 1 1 33564
0 33566 7 1 2 87317 33565
0 33567 5 1 1 33566
0 33568 7 3 2 79291 86173
0 33569 5 1 1 94926
0 33570 7 1 2 81774 86997
0 33571 7 1 2 94927 33570
0 33572 5 1 1 33571
0 33573 7 1 2 33567 33572
0 33574 5 1 1 33573
0 33575 7 1 2 70810 33574
0 33576 5 1 1 33575
0 33577 7 1 2 87342 94059
0 33578 7 1 2 94449 33577
0 33579 5 1 1 33578
0 33580 7 1 2 33576 33579
0 33581 5 1 1 33580
0 33582 7 1 2 94924 33581
0 33583 5 1 1 33582
0 33584 7 2 2 63064 81466
0 33585 5 1 1 94929
0 33586 7 1 2 94142 94904
0 33587 7 1 2 94930 33586
0 33588 5 1 1 33587
0 33589 7 1 2 68716 33588
0 33590 7 1 2 33583 33589
0 33591 7 1 2 33559 33590
0 33592 5 1 1 33591
0 33593 7 5 2 60554 87629
0 33594 5 4 1 94931
0 33595 7 1 2 65454 92308
0 33596 5 2 1 33595
0 33597 7 1 2 94936 94940
0 33598 5 2 1 33597
0 33599 7 1 2 94319 94942
0 33600 5 1 1 33599
0 33601 7 1 2 60668 81759
0 33602 5 1 1 33601
0 33603 7 1 2 33600 33602
0 33604 5 1 1 33603
0 33605 7 1 2 66543 33604
0 33606 5 1 1 33605
0 33607 7 3 2 65006 87848
0 33608 7 1 2 86642 94944
0 33609 5 1 1 33608
0 33610 7 1 2 33606 33609
0 33611 5 1 1 33610
0 33612 7 1 2 64548 33611
0 33613 5 1 1 33612
0 33614 7 1 2 85880 87830
0 33615 7 1 2 74660 33614
0 33616 7 1 2 94094 33615
0 33617 5 1 1 33616
0 33618 7 1 2 33613 33617
0 33619 5 1 1 33618
0 33620 7 1 2 65250 33619
0 33621 5 1 1 33620
0 33622 7 2 2 64014 79264
0 33623 7 1 2 87849 93429
0 33624 7 1 2 82788 33623
0 33625 7 1 2 94947 33624
0 33626 5 1 1 33625
0 33627 7 1 2 33621 33626
0 33628 5 1 1 33627
0 33629 7 1 2 66867 33628
0 33630 5 1 1 33629
0 33631 7 1 2 65590 94102
0 33632 7 2 2 64549 81775
0 33633 7 1 2 94320 94949
0 33634 7 1 2 33631 33633
0 33635 5 1 1 33634
0 33636 7 1 2 33630 33635
0 33637 5 1 1 33636
0 33638 7 1 2 81571 33637
0 33639 5 1 1 33638
0 33640 7 2 2 79702 87146
0 33641 7 3 2 89363 94321
0 33642 7 1 2 94951 94953
0 33643 5 1 1 33642
0 33644 7 2 2 79344 92768
0 33645 7 1 2 94954 94956
0 33646 5 1 1 33645
0 33647 7 1 2 81783 94955
0 33648 5 1 1 33647
0 33649 7 1 2 71565 87916
0 33650 7 1 2 73277 33649
0 33651 5 1 1 33650
0 33652 7 1 2 33648 33651
0 33653 5 1 1 33652
0 33654 7 1 2 66544 33653
0 33655 5 1 1 33654
0 33656 7 1 2 79469 86643
0 33657 7 1 2 73278 33656
0 33658 5 1 1 33657
0 33659 7 1 2 33655 33658
0 33660 5 1 1 33659
0 33661 7 1 2 60669 33660
0 33662 5 1 1 33661
0 33663 7 1 2 33646 33662
0 33664 5 1 1 33663
0 33665 7 1 2 66868 33664
0 33666 5 1 1 33665
0 33667 7 1 2 33643 33666
0 33668 5 1 1 33667
0 33669 7 1 2 69257 33668
0 33670 5 1 1 33669
0 33671 7 1 2 81287 86503
0 33672 7 2 2 65007 65591
0 33673 7 1 2 94419 94958
0 33674 7 1 2 33671 33673
0 33675 7 1 2 68888 69071
0 33676 7 1 2 92905 33675
0 33677 7 2 2 33674 33676
0 33678 5 1 1 94960
0 33679 7 3 2 87219 94911
0 33680 5 1 1 94962
0 33681 7 1 2 73377 90860
0 33682 5 1 1 33681
0 33683 7 2 2 70188 33682
0 33684 5 2 1 94965
0 33685 7 1 2 87147 94967
0 33686 5 1 1 33685
0 33687 7 1 2 66869 94945
0 33688 5 1 1 33687
0 33689 7 1 2 33686 33688
0 33690 5 1 1 33689
0 33691 7 1 2 79628 33690
0 33692 5 1 1 33691
0 33693 7 1 2 33680 33692
0 33694 5 1 1 33693
0 33695 7 1 2 68889 33694
0 33696 5 1 1 33695
0 33697 7 1 2 72779 90303
0 33698 5 1 1 33697
0 33699 7 1 2 64550 33698
0 33700 5 1 1 33699
0 33701 7 1 2 82684 91386
0 33702 7 1 2 33700 33701
0 33703 5 1 1 33702
0 33704 7 1 2 68890 87507
0 33705 7 1 2 33703 33704
0 33706 5 1 1 33705
0 33707 7 2 2 61737 86788
0 33708 5 1 1 94969
0 33709 7 1 2 79141 94970
0 33710 5 1 1 33709
0 33711 7 1 2 11922 33710
0 33712 7 1 2 33706 33711
0 33713 5 1 1 33712
0 33714 7 1 2 70811 33713
0 33715 5 1 1 33714
0 33716 7 1 2 33696 33715
0 33717 5 1 1 33716
0 33718 7 1 2 66545 33717
0 33719 5 1 1 33718
0 33720 7 1 2 33678 33719
0 33721 5 1 1 33720
0 33722 7 1 2 65251 33721
0 33723 5 1 1 33722
0 33724 7 3 2 73523 94322
0 33725 7 1 2 79703 94971
0 33726 5 1 1 33725
0 33727 7 1 2 64303 78061
0 33728 7 1 2 81836 33727
0 33729 7 1 2 91088 33728
0 33730 5 1 1 33729
0 33731 7 1 2 33726 33730
0 33732 5 1 1 33731
0 33733 7 1 2 60670 33732
0 33734 5 1 1 33733
0 33735 7 1 2 94957 94972
0 33736 5 1 1 33735
0 33737 7 1 2 33734 33736
0 33738 5 1 1 33737
0 33739 7 1 2 66870 33738
0 33740 5 1 1 33739
0 33741 7 1 2 94952 94973
0 33742 5 1 1 33741
0 33743 7 1 2 33740 33742
0 33744 5 1 1 33743
0 33745 7 1 2 70316 33744
0 33746 5 1 1 33745
0 33747 7 1 2 66546 94961
0 33748 5 1 1 33747
0 33749 7 1 2 91298 94943
0 33750 5 1 1 33749
0 33751 7 1 2 11175 94941
0 33752 5 1 1 33751
0 33753 7 1 2 79124 33752
0 33754 5 1 1 33753
0 33755 7 1 2 33750 33754
0 33756 5 1 1 33755
0 33757 7 3 2 59905 76928
0 33758 5 2 1 94974
0 33759 7 1 2 69258 94977
0 33760 5 1 1 33759
0 33761 7 2 2 81572 82805
0 33762 5 2 1 94979
0 33763 7 1 2 33760 94981
0 33764 5 1 1 33763
0 33765 7 1 2 86099 33764
0 33766 5 1 1 33765
0 33767 7 2 2 81291 94919
0 33768 5 1 1 94983
0 33769 7 1 2 73894 94984
0 33770 5 1 1 33769
0 33771 7 1 2 33766 33770
0 33772 5 1 1 33771
0 33773 7 1 2 33756 33772
0 33774 5 1 1 33773
0 33775 7 1 2 33748 33774
0 33776 7 1 2 33746 33775
0 33777 7 1 2 33723 33776
0 33778 7 1 2 33670 33777
0 33779 7 1 2 33639 33778
0 33780 5 1 1 33779
0 33781 7 1 2 63065 33780
0 33782 5 1 1 33781
0 33783 7 1 2 86120 33768
0 33784 5 1 1 33783
0 33785 7 1 2 65592 33784
0 33786 5 1 1 33785
0 33787 7 1 2 10757 33786
0 33788 5 1 1 33787
0 33789 7 1 2 63066 33788
0 33790 5 1 1 33789
0 33791 7 1 2 33790 33496
0 33792 5 1 1 33791
0 33793 7 1 2 70812 33792
0 33794 5 1 1 33793
0 33795 7 1 2 60369 94966
0 33796 5 1 1 33795
0 33797 7 1 2 94486 33796
0 33798 5 1 1 33797
0 33799 7 1 2 33794 33798
0 33800 5 1 1 33799
0 33801 7 1 2 61569 33800
0 33802 5 1 1 33801
0 33803 7 3 2 65593 61357
0 33804 7 2 2 82411 86174
0 33805 5 1 1 94988
0 33806 7 3 2 94985 94989
0 33807 5 1 1 94990
0 33808 7 1 2 65008 94991
0 33809 5 1 1 33808
0 33810 7 1 2 70813 73043
0 33811 7 1 2 88070 33810
0 33812 5 1 1 33811
0 33813 7 1 2 33492 33812
0 33814 5 1 1 33813
0 33815 7 1 2 63067 33814
0 33816 5 1 1 33815
0 33817 7 1 2 62343 94907
0 33818 5 1 1 33817
0 33819 7 1 2 33816 33818
0 33820 5 1 1 33819
0 33821 7 1 2 61570 33820
0 33822 5 1 1 33821
0 33823 7 1 2 62344 94992
0 33824 5 1 1 33823
0 33825 7 1 2 33822 33824
0 33826 5 1 1 33825
0 33827 7 1 2 73576 33826
0 33828 5 1 1 33827
0 33829 7 1 2 33809 33828
0 33830 7 1 2 33513 33529
0 33831 5 1 1 33830
0 33832 7 1 2 61571 33831
0 33833 5 1 1 33832
0 33834 7 1 2 33807 33833
0 33835 5 2 1 33834
0 33836 7 1 2 62132 81837
0 33837 7 1 2 94993 33836
0 33838 5 1 1 33837
0 33839 7 4 2 81292 91126
0 33840 7 1 2 66871 71800
0 33841 7 1 2 86998 33840
0 33842 7 1 2 94995 33841
0 33843 5 1 1 33842
0 33844 7 1 2 33838 33843
0 33845 5 1 1 33844
0 33846 7 1 2 69682 33845
0 33847 5 1 1 33846
0 33848 7 1 2 80240 94994
0 33849 5 1 1 33848
0 33850 7 1 2 59906 17612
0 33851 5 1 1 33850
0 33852 7 1 2 88071 94324
0 33853 7 1 2 33851 33852
0 33854 5 1 1 33853
0 33855 7 1 2 33849 33854
0 33856 5 1 1 33855
0 33857 7 1 2 71801 33856
0 33858 5 1 1 33857
0 33859 7 1 2 33847 33858
0 33860 7 1 2 33829 33859
0 33861 7 1 2 33802 33860
0 33862 5 1 1 33861
0 33863 7 1 2 81190 33862
0 33864 5 1 1 33863
0 33865 7 1 2 93886 93700
0 33866 5 2 1 33865
0 33867 7 1 2 60671 94999
0 33868 5 1 1 33867
0 33869 7 3 2 68891 87148
0 33870 7 2 2 66321 95001
0 33871 5 1 1 95004
0 33872 7 1 2 33868 33871
0 33873 5 1 1 33872
0 33874 7 1 2 79629 33873
0 33875 5 1 1 33874
0 33876 7 1 2 81733 88072
0 33877 5 1 1 33876
0 33878 7 1 2 33875 33877
0 33879 5 1 1 33878
0 33880 7 1 2 65009 33879
0 33881 5 1 1 33880
0 33882 7 1 2 85881 86504
0 33883 7 1 2 82043 33882
0 33884 5 1 1 33883
0 33885 7 1 2 33881 33884
0 33886 5 1 1 33885
0 33887 7 1 2 80241 33886
0 33888 5 1 1 33887
0 33889 7 1 2 88033 93414
0 33890 5 1 1 33889
0 33891 7 1 2 33888 33890
0 33892 5 1 1 33891
0 33893 7 1 2 71802 33892
0 33894 5 1 1 33893
0 33895 7 1 2 70885 92841
0 33896 5 1 1 33895
0 33897 7 2 2 68892 87173
0 33898 7 1 2 64551 76859
0 33899 7 1 2 95006 33898
0 33900 5 1 1 33899
0 33901 7 1 2 33896 33900
0 33902 5 1 1 33901
0 33903 7 1 2 79630 33902
0 33904 5 1 1 33903
0 33905 7 2 2 81729 92769
0 33906 7 1 2 80756 86204
0 33907 7 1 2 95008 33906
0 33908 5 1 1 33907
0 33909 7 1 2 33904 33908
0 33910 5 1 1 33909
0 33911 7 1 2 69259 33910
0 33912 5 1 1 33911
0 33913 7 1 2 70061 86205
0 33914 5 1 1 33913
0 33915 7 1 2 80587 86100
0 33916 5 1 1 33915
0 33917 7 1 2 33914 33916
0 33918 5 1 1 33917
0 33919 7 1 2 60672 33918
0 33920 5 1 1 33919
0 33921 7 2 2 65010 95005
0 33922 5 1 1 95010
0 33923 7 1 2 62133 95011
0 33924 5 1 1 33923
0 33925 7 1 2 33920 33924
0 33926 5 1 1 33925
0 33927 7 1 2 79631 33926
0 33928 5 1 1 33927
0 33929 7 1 2 81787 94963
0 33930 5 1 1 33929
0 33931 7 1 2 33928 33930
0 33932 5 1 1 33931
0 33933 7 1 2 81573 33932
0 33934 5 1 1 33933
0 33935 7 1 2 33912 33934
0 33936 5 1 1 33935
0 33937 7 1 2 69683 33936
0 33938 5 1 1 33937
0 33939 7 1 2 81293 94964
0 33940 5 1 1 33939
0 33941 7 1 2 65011 95000
0 33942 5 1 1 33941
0 33943 7 1 2 66322 93884
0 33944 5 1 1 33943
0 33945 7 1 2 33942 33944
0 33946 5 1 1 33945
0 33947 7 1 2 60673 33946
0 33948 5 1 1 33947
0 33949 7 1 2 33948 33922
0 33950 5 1 1 33949
0 33951 7 1 2 79632 69991
0 33952 7 1 2 33950 33951
0 33953 5 1 1 33952
0 33954 7 1 2 33940 33953
0 33955 5 1 1 33954
0 33956 7 1 2 73577 33955
0 33957 5 1 1 33956
0 33958 7 1 2 73875 88571
0 33959 5 1 1 33958
0 33960 7 2 2 70189 33959
0 33961 5 2 1 95012
0 33962 7 1 2 88034 95014
0 33963 5 1 1 33962
0 33964 7 1 2 33957 33963
0 33965 7 1 2 33938 33964
0 33966 7 1 2 33894 33965
0 33967 5 1 1 33966
0 33968 7 1 2 75223 33967
0 33969 5 1 1 33968
0 33970 7 1 2 63782 33969
0 33971 7 1 2 33864 33970
0 33972 7 1 2 33782 33971
0 33973 5 1 1 33972
0 33974 7 1 2 63504 33973
0 33975 7 1 2 33592 33974
0 33976 5 1 1 33975
0 33977 7 1 2 79301 85652
0 33978 5 1 1 33977
0 33979 7 1 2 87252 33978
0 33980 5 1 1 33979
0 33981 7 1 2 88073 33980
0 33982 5 1 1 33981
0 33983 7 1 2 60555 87578
0 33984 5 1 1 33983
0 33985 7 1 2 80376 33984
0 33986 5 1 1 33985
0 33987 7 4 2 63068 80276
0 33988 7 1 2 87398 95016
0 33989 7 1 2 33986 33988
0 33990 5 1 1 33989
0 33991 7 1 2 33982 33990
0 33992 5 3 1 33991
0 33993 7 1 2 62134 95020
0 33994 5 1 1 33993
0 33995 7 1 2 83483 88050
0 33996 7 1 2 88057 33995
0 33997 5 1 1 33996
0 33998 7 1 2 33994 33997
0 33999 5 1 1 33998
0 34000 7 1 2 68397 33999
0 34001 5 1 1 34000
0 34002 7 1 2 81000 87322
0 34003 7 2 2 87851 34002
0 34004 5 1 1 95023
0 34005 7 1 2 62135 95024
0 34006 5 1 1 34005
0 34007 7 1 2 34001 34006
0 34008 5 1 1 34007
0 34009 7 1 2 71803 34008
0 34010 5 1 1 34009
0 34011 7 4 2 68398 70814
0 34012 7 1 2 94462 94487
0 34013 5 1 1 34012
0 34014 7 1 2 86364 87446
0 34015 7 1 2 87399 34014
0 34016 5 1 1 34015
0 34017 7 1 2 34013 34016
0 34018 5 1 1 34017
0 34019 7 1 2 75603 34018
0 34020 5 1 1 34019
0 34021 7 1 2 80360 84765
0 34022 7 1 2 87400 34021
0 34023 5 1 1 34022
0 34024 7 1 2 34020 34023
0 34025 5 1 1 34024
0 34026 7 1 2 95025 34025
0 34027 5 1 1 34026
0 34028 7 1 2 34010 34027
0 34029 5 1 1 34028
0 34030 7 1 2 64775 34029
0 34031 5 1 1 34030
0 34032 7 2 2 66872 71999
0 34033 7 1 2 94996 95029
0 34034 5 1 1 34033
0 34035 7 1 2 71566 86101
0 34036 5 2 1 34035
0 34037 7 1 2 34034 95031
0 34038 5 1 1 34037
0 34039 7 1 2 65594 34038
0 34040 5 1 1 34039
0 34041 7 1 2 71567 87142
0 34042 5 2 1 34041
0 34043 7 1 2 34040 95033
0 34044 5 1 1 34043
0 34045 7 1 2 94143 34044
0 34046 5 1 1 34045
0 34047 7 1 2 80523 93674
0 34048 5 2 1 34047
0 34049 7 2 2 80422 94997
0 34050 7 1 2 95030 95037
0 34051 5 1 1 34050
0 34052 7 1 2 95035 34051
0 34053 5 1 1 34052
0 34054 7 1 2 65595 34053
0 34055 5 1 1 34054
0 34056 7 1 2 87711 94878
0 34057 7 1 2 94912 34056
0 34058 5 2 1 34057
0 34059 7 1 2 34055 95039
0 34060 5 1 1 34059
0 34061 7 1 2 65252 34060
0 34062 5 1 1 34061
0 34063 7 1 2 34046 34062
0 34064 5 1 1 34063
0 34065 7 1 2 68399 34064
0 34066 5 1 1 34065
0 34067 7 1 2 34031 34066
0 34068 5 1 1 34067
0 34069 7 1 2 63783 34068
0 34070 5 1 1 34069
0 34071 7 2 2 80423 93185
0 34072 5 1 1 95041
0 34073 7 1 2 86716 95042
0 34074 5 1 1 34073
0 34075 7 1 2 75321 95013
0 34076 5 1 1 34075
0 34077 7 1 2 75604 87508
0 34078 7 1 2 34076 34077
0 34079 5 1 1 34078
0 34080 7 1 2 34074 34079
0 34081 5 1 1 34080
0 34082 7 1 2 70494 90111
0 34083 7 1 2 34081 34082
0 34084 5 1 1 34083
0 34085 7 1 2 34070 34084
0 34086 5 1 1 34085
0 34087 7 1 2 69684 34086
0 34088 5 1 1 34087
0 34089 7 1 2 68400 95021
0 34090 5 1 1 34089
0 34091 7 1 2 34004 34090
0 34092 5 1 1 34091
0 34093 7 1 2 69992 34092
0 34094 5 1 1 34093
0 34095 7 1 2 81288 85453
0 34096 5 1 1 34095
0 34097 7 1 2 75605 94589
0 34098 5 1 1 34097
0 34099 7 1 2 34096 34098
0 34100 5 1 1 34099
0 34101 7 1 2 69850 87401
0 34102 7 1 2 34100 34101
0 34103 5 1 1 34102
0 34104 7 1 2 80333 94488
0 34105 5 1 1 34104
0 34106 7 1 2 92770 94126
0 34107 5 1 1 34106
0 34108 7 1 2 34105 34107
0 34109 5 1 1 34108
0 34110 7 1 2 75606 73044
0 34111 7 1 2 34109 34110
0 34112 5 1 1 34111
0 34113 7 1 2 34103 34112
0 34114 5 1 1 34113
0 34115 7 1 2 95026 34114
0 34116 5 1 1 34115
0 34117 7 1 2 34094 34116
0 34118 5 1 1 34117
0 34119 7 1 2 64776 34118
0 34120 5 1 1 34119
0 34121 7 1 2 94920 94998
0 34122 5 1 1 34121
0 34123 7 1 2 95032 34122
0 34124 5 1 1 34123
0 34125 7 1 2 65596 34124
0 34126 5 1 1 34125
0 34127 7 1 2 95034 34126
0 34128 5 1 1 34127
0 34129 7 1 2 94144 34128
0 34130 5 1 1 34129
0 34131 7 1 2 94921 95038
0 34132 5 1 1 34131
0 34133 7 1 2 95036 34132
0 34134 5 1 1 34133
0 34135 7 1 2 65597 34134
0 34136 5 1 1 34135
0 34137 7 1 2 95040 34136
0 34138 5 1 1 34137
0 34139 7 1 2 65253 34138
0 34140 5 1 1 34139
0 34141 7 1 2 34130 34140
0 34142 5 1 1 34141
0 34143 7 1 2 68401 34142
0 34144 5 1 1 34143
0 34145 7 1 2 34120 34144
0 34146 5 1 1 34145
0 34147 7 1 2 63784 34146
0 34148 5 1 1 34147
0 34149 7 1 2 80277 80504
0 34150 5 1 1 34149
0 34151 7 1 2 83479 34150
0 34152 5 1 1 34151
0 34153 7 1 2 63069 34152
0 34154 5 1 1 34153
0 34155 7 1 2 87247 34154
0 34156 5 1 1 34155
0 34157 7 1 2 80871 34156
0 34158 5 1 1 34157
0 34159 7 1 2 34072 34158
0 34160 5 1 1 34159
0 34161 7 1 2 66873 34160
0 34162 5 1 1 34161
0 34163 7 1 2 87155 34162
0 34164 5 1 1 34163
0 34165 7 1 2 80505 94191
0 34166 5 1 1 34165
0 34167 7 1 2 93593 94437
0 34168 5 1 1 34167
0 34169 7 1 2 34166 34168
0 34170 5 1 1 34169
0 34171 7 1 2 63070 34170
0 34172 5 1 1 34171
0 34173 7 1 2 79633 87240
0 34174 5 1 1 34173
0 34175 7 1 2 86736 34174
0 34176 7 1 2 34172 34175
0 34177 5 1 1 34176
0 34178 7 1 2 64015 34177
0 34179 7 1 2 34164 34178
0 34180 5 1 1 34179
0 34181 7 1 2 80506 87241
0 34182 5 1 1 34181
0 34183 7 1 2 90777 34182
0 34184 5 1 1 34183
0 34185 7 1 2 88020 94928
0 34186 7 1 2 34184 34185
0 34187 5 1 1 34186
0 34188 7 1 2 34180 34187
0 34189 5 1 1 34188
0 34190 7 1 2 94710 34189
0 34191 5 1 1 34190
0 34192 7 1 2 34148 34191
0 34193 5 1 1 34192
0 34194 7 1 2 71804 34193
0 34195 5 1 1 34194
0 34196 7 1 2 80361 79381
0 34197 5 2 1 34196
0 34198 7 1 2 84152 85369
0 34199 5 2 1 34198
0 34200 7 1 2 84548 95045
0 34201 5 1 1 34200
0 34202 7 2 2 63071 34201
0 34203 5 1 1 95047
0 34204 7 1 2 84084 84348
0 34205 5 1 1 34204
0 34206 7 1 2 93587 34205
0 34207 5 2 1 34206
0 34208 7 1 2 66323 95049
0 34209 5 1 1 34208
0 34210 7 1 2 34203 34209
0 34211 5 2 1 34210
0 34212 7 1 2 65455 95051
0 34213 5 1 1 34212
0 34214 7 1 2 95043 34213
0 34215 5 1 1 34214
0 34216 7 1 2 75607 34215
0 34217 5 1 1 34216
0 34218 7 1 2 81034 93921
0 34219 5 1 1 34218
0 34220 7 1 2 34217 34219
0 34221 5 1 1 34220
0 34222 7 1 2 87143 34221
0 34223 5 1 1 34222
0 34224 7 1 2 72447 90214
0 34225 5 1 1 34224
0 34226 7 1 2 85522 88117
0 34227 5 1 1 34226
0 34228 7 1 2 34225 34227
0 34229 5 1 1 34228
0 34230 7 1 2 66324 34229
0 34231 5 1 1 34230
0 34232 7 1 2 87611 92371
0 34233 5 1 1 34232
0 34234 7 1 2 81301 85523
0 34235 5 1 1 34234
0 34236 7 1 2 34233 34235
0 34237 7 1 2 34231 34236
0 34238 5 1 1 34237
0 34239 7 1 2 66874 34238
0 34240 5 1 1 34239
0 34241 7 1 2 63785 79588
0 34242 7 1 2 93740 34241
0 34243 5 1 1 34242
0 34244 7 1 2 34240 34243
0 34245 5 1 1 34244
0 34246 7 1 2 66547 34245
0 34247 5 1 1 34246
0 34248 7 1 2 86121 93701
0 34249 5 1 1 34248
0 34250 7 1 2 92269 34249
0 34251 5 1 1 34250
0 34252 7 1 2 86316 87899
0 34253 5 1 1 34252
0 34254 7 1 2 34251 34253
0 34255 5 1 1 34254
0 34256 7 1 2 79105 34255
0 34257 5 1 1 34256
0 34258 7 1 2 60556 34257
0 34259 7 1 2 34247 34258
0 34260 5 1 1 34259
0 34261 7 1 2 86102 95052
0 34262 5 1 1 34261
0 34263 7 3 2 84485 86175
0 34264 7 1 2 78575 95053
0 34265 5 1 1 34264
0 34266 7 1 2 34262 34265
0 34267 5 1 1 34266
0 34268 7 1 2 75608 34267
0 34269 5 1 1 34268
0 34270 7 1 2 85343 87896
0 34271 5 1 1 34270
0 34272 7 1 2 84549 34271
0 34273 5 1 1 34272
0 34274 7 1 2 75224 34273
0 34275 5 1 1 34274
0 34276 7 1 2 84438 86870
0 34277 5 1 1 34276
0 34278 7 1 2 34275 34277
0 34279 5 1 1 34278
0 34280 7 1 2 86176 34279
0 34281 5 1 1 34280
0 34282 7 1 2 65456 34281
0 34283 7 1 2 34269 34282
0 34284 5 1 1 34283
0 34285 7 1 2 65598 34284
0 34286 7 1 2 34260 34285
0 34287 5 1 1 34286
0 34288 7 1 2 34223 34287
0 34289 5 1 1 34288
0 34290 7 1 2 82720 34289
0 34291 5 1 1 34290
0 34292 7 2 2 74711 79348
0 34293 5 1 1 95056
0 34294 7 1 2 60557 34293
0 34295 5 1 1 34294
0 34296 7 2 2 76583 84486
0 34297 5 1 1 95058
0 34298 7 1 2 34295 95059
0 34299 5 1 1 34298
0 34300 7 2 2 72000 77992
0 34301 7 1 2 80903 91345
0 34302 7 1 2 95060 34301
0 34303 5 1 1 34302
0 34304 7 1 2 79650 34303
0 34305 5 1 1 34304
0 34306 7 1 2 79634 2381
0 34307 5 1 1 34306
0 34308 7 1 2 60161 34307
0 34309 5 1 1 34308
0 34310 7 1 2 68717 34309
0 34311 7 1 2 34305 34310
0 34312 5 1 1 34311
0 34313 7 1 2 34299 34312
0 34314 5 1 1 34313
0 34315 7 1 2 87687 34314
0 34316 5 1 1 34315
0 34317 7 2 2 60370 4898
0 34318 5 3 1 95062
0 34319 7 1 2 93922 95064
0 34320 5 1 1 34319
0 34321 7 1 2 77123 92270
0 34322 7 1 2 71568 34321
0 34323 5 1 1 34322
0 34324 7 1 2 34320 34323
0 34325 5 1 1 34324
0 34326 7 1 2 86789 34325
0 34327 5 1 1 34326
0 34328 7 1 2 70815 86423
0 34329 7 1 2 88152 34328
0 34330 5 1 1 34329
0 34331 7 1 2 65599 72448
0 34332 7 1 2 92779 34331
0 34333 7 1 2 95065 34332
0 34334 5 1 1 34333
0 34335 7 1 2 34330 34334
0 34336 7 1 2 34327 34335
0 34337 5 1 1 34336
0 34338 7 1 2 60558 34337
0 34339 5 1 1 34338
0 34340 7 1 2 34316 34339
0 34341 5 1 1 34340
0 34342 7 1 2 66548 34341
0 34343 5 1 1 34342
0 34344 7 1 2 70495 92787
0 34345 5 1 1 34344
0 34346 7 1 2 80377 95046
0 34347 5 1 1 34346
0 34348 7 1 2 87174 20257
0 34349 7 1 2 34347 34348
0 34350 5 1 1 34349
0 34351 7 1 2 34345 34350
0 34352 5 1 1 34351
0 34353 7 1 2 95057 34352
0 34354 5 1 1 34353
0 34355 7 1 2 34343 34354
0 34356 5 1 1 34355
0 34357 7 1 2 64016 34356
0 34358 5 1 1 34357
0 34359 7 1 2 65457 95048
0 34360 5 1 1 34359
0 34361 7 1 2 95044 34360
0 34362 5 1 1 34361
0 34363 7 1 2 66325 34362
0 34364 5 1 1 34363
0 34365 7 1 2 77124 88224
0 34366 5 1 1 34365
0 34367 7 1 2 74712 95050
0 34368 5 1 1 34367
0 34369 7 1 2 34366 34368
0 34370 5 1 1 34369
0 34371 7 1 2 81272 34370
0 34372 5 1 1 34371
0 34373 7 1 2 34364 34372
0 34374 5 1 1 34373
0 34375 7 1 2 87175 34374
0 34376 5 1 1 34375
0 34377 7 2 2 78711 86317
0 34378 7 1 2 68718 95009
0 34379 7 1 2 95067 34378
0 34380 5 1 1 34379
0 34381 7 1 2 34376 34380
0 34382 5 1 1 34381
0 34383 7 1 2 64017 34382
0 34384 5 1 1 34383
0 34385 7 1 2 84144 82952
0 34386 5 1 1 34385
0 34387 7 1 2 62345 85357
0 34388 5 1 1 34387
0 34389 7 1 2 34386 34388
0 34390 5 1 1 34389
0 34391 7 2 2 86177 34390
0 34392 7 1 2 73895 94959
0 34393 7 1 2 95069 34392
0 34394 5 1 1 34393
0 34395 7 1 2 34384 34394
0 34396 5 1 1 34395
0 34397 7 1 2 75609 34396
0 34398 5 1 1 34397
0 34399 7 1 2 94917 95070
0 34400 5 1 1 34399
0 34401 7 1 2 34398 34400
0 34402 7 1 2 34358 34401
0 34403 7 1 2 34291 34402
0 34404 5 1 1 34403
0 34405 7 1 2 68402 34404
0 34406 5 1 1 34405
0 34407 7 1 2 84145 88074
0 34408 7 1 2 90995 34407
0 34409 5 1 1 34408
0 34410 7 1 2 31042 34409
0 34411 5 1 1 34410
0 34412 7 1 2 86837 34411
0 34413 5 1 1 34412
0 34414 7 2 2 81776 87071
0 34415 7 2 2 94781 95071
0 34416 7 1 2 68893 85344
0 34417 7 1 2 95073 34416
0 34418 5 1 1 34417
0 34419 7 1 2 34413 34418
0 34420 5 1 1 34419
0 34421 7 1 2 70816 34420
0 34422 5 1 1 34421
0 34423 7 1 2 63786 84085
0 34424 7 1 2 95022 34423
0 34425 5 1 1 34424
0 34426 7 1 2 34422 34425
0 34427 5 1 1 34426
0 34428 7 1 2 68403 34427
0 34429 5 1 1 34428
0 34430 7 1 2 85846 91323
0 34431 7 1 2 94422 34430
0 34432 7 1 2 94454 94946
0 34433 7 1 2 34431 34432
0 34434 5 1 1 34433
0 34435 7 1 2 34429 34434
0 34436 5 1 1 34435
0 34437 7 1 2 73578 34436
0 34438 5 1 1 34437
0 34439 7 1 2 60674 65885
0 34440 7 1 2 74836 34439
0 34441 7 1 2 94033 34440
0 34442 7 1 2 94452 34441
0 34443 5 1 1 34442
0 34444 7 1 2 34438 34443
0 34445 7 1 2 34406 34444
0 34446 7 1 2 34195 34445
0 34447 7 1 2 34088 34446
0 34448 7 1 2 33976 34447
0 34449 5 2 1 34448
0 34450 7 1 2 64104 95075
0 34451 5 1 1 34450
0 34452 7 1 2 92906 93623
0 34453 5 1 1 34452
0 34454 7 1 2 71495 94510
0 34455 5 1 1 34454
0 34456 7 1 2 63072 90656
0 34457 7 1 2 34455 34456
0 34458 5 1 1 34457
0 34459 7 1 2 34453 34458
0 34460 5 1 1 34459
0 34461 7 1 2 65012 34460
0 34462 5 1 1 34461
0 34463 7 1 2 94865 95061
0 34464 5 1 1 34463
0 34465 7 1 2 34462 34464
0 34466 5 2 1 34465
0 34467 7 1 2 84741 94605
0 34468 7 1 2 95074 34467
0 34469 7 2 2 95077 34468
0 34470 5 1 1 95079
0 34471 7 1 2 34451 34470
0 34472 5 1 1 34471
0 34473 7 1 2 71922 34472
0 34474 5 1 1 34473
0 34475 7 2 2 87016 95072
0 34476 5 1 1 95081
0 34477 7 1 2 66875 93802
0 34478 5 1 1 34477
0 34479 7 1 2 86069 34478
0 34480 5 1 1 34479
0 34481 7 1 2 65600 34480
0 34482 5 1 1 34481
0 34483 7 1 2 34476 34482
0 34484 5 1 1 34483
0 34485 7 1 2 73524 73838
0 34486 5 1 1 34485
0 34487 7 1 2 8230 34486
0 34488 5 1 1 34487
0 34489 7 1 2 64777 34488
0 34490 5 1 1 34489
0 34491 7 1 2 93377 34490
0 34492 5 1 1 34491
0 34493 7 1 2 63505 34492
0 34494 7 1 2 34484 34493
0 34495 5 1 1 34494
0 34496 7 1 2 59558 84583
0 34497 5 1 1 34496
0 34498 7 1 2 92990 94146
0 34499 7 1 2 34497 34498
0 34500 5 1 1 34499
0 34501 7 1 2 84240 34500
0 34502 5 1 1 34501
0 34503 7 1 2 86717 93827
0 34504 7 1 2 34502 34503
0 34505 5 1 1 34504
0 34506 7 1 2 34495 34505
0 34507 5 1 1 34506
0 34508 7 1 2 63787 34507
0 34509 5 1 1 34508
0 34510 7 2 2 66876 63506
0 34511 7 1 2 65601 78072
0 34512 7 1 2 95083 34511
0 34513 7 1 2 80424 90716
0 34514 7 1 2 34512 34513
0 34515 7 1 2 74612 34514
0 34516 5 1 1 34515
0 34517 7 1 2 34509 34516
0 34518 5 1 1 34517
0 34519 7 1 2 69685 34518
0 34520 5 1 1 34519
0 34521 7 2 2 72726 91935
0 34522 7 1 2 69851 95085
0 34523 5 1 1 34522
0 34524 7 1 2 71805 72891
0 34525 5 1 1 34524
0 34526 7 1 2 34523 34525
0 34527 5 1 1 34526
0 34528 7 1 2 88153 90694
0 34529 7 1 2 84225 34528
0 34530 7 1 2 34527 34529
0 34531 5 1 1 34530
0 34532 7 1 2 34520 34531
0 34533 5 1 1 34532
0 34534 7 1 2 94748 34533
0 34535 5 1 1 34534
0 34536 7 1 2 81107 88235
0 34537 7 1 2 94696 34536
0 34538 7 1 2 93198 34537
0 34539 5 1 1 34538
0 34540 7 1 2 32345 34539
0 34541 5 1 1 34540
0 34542 7 1 2 64778 34541
0 34543 5 1 1 34542
0 34544 7 1 2 84349 84747
0 34545 5 1 1 34544
0 34546 7 7 2 61738 78774
0 34547 5 3 1 95087
0 34548 7 1 2 77530 95088
0 34549 5 1 1 34548
0 34550 7 1 2 34545 34549
0 34551 5 1 1 34550
0 34552 7 1 2 65458 34551
0 34553 5 1 1 34552
0 34554 7 1 2 34543 34553
0 34555 5 1 1 34554
0 34556 7 1 2 66043 34555
0 34557 5 1 1 34556
0 34558 7 1 2 93494 30828
0 34559 5 1 1 34558
0 34560 7 1 2 85328 34559
0 34561 5 1 1 34560
0 34562 7 1 2 34557 34561
0 34563 5 1 1 34562
0 34564 7 1 2 64304 34563
0 34565 5 1 1 34564
0 34566 7 1 2 94675 32087
0 34567 5 2 1 34566
0 34568 7 1 2 79635 94385
0 34569 7 1 2 95097 34568
0 34570 5 1 1 34569
0 34571 7 1 2 34565 34570
0 34572 5 1 1 34571
0 34573 7 1 2 62693 34572
0 34574 5 1 1 34573
0 34575 7 1 2 84350 91311
0 34576 5 1 1 34575
0 34577 7 1 2 33433 34576
0 34578 5 1 1 34577
0 34579 7 1 2 69852 34578
0 34580 5 1 1 34579
0 34581 7 2 2 86424 88236
0 34582 5 1 1 95099
0 34583 7 1 2 34580 34582
0 34584 5 1 1 34583
0 34585 7 1 2 65013 82178
0 34586 7 1 2 34584 34585
0 34587 5 1 1 34586
0 34588 7 1 2 34574 34587
0 34589 5 1 1 34588
0 34590 7 1 2 71806 34589
0 34591 5 1 1 34590
0 34592 7 1 2 80302 84487
0 34593 5 1 1 34592
0 34594 7 1 2 12168 34593
0 34595 5 1 1 34594
0 34596 7 1 2 72001 34595
0 34597 5 1 1 34596
0 34598 7 1 2 80660 84488
0 34599 5 1 1 34598
0 34600 7 1 2 12170 34599
0 34601 7 1 2 34597 34600
0 34602 5 1 1 34601
0 34603 7 1 2 73699 34602
0 34604 5 1 1 34603
0 34605 7 1 2 73839 94850
0 34606 5 1 1 34605
0 34607 7 1 2 65014 33054
0 34608 5 1 1 34607
0 34609 7 1 2 8604 34608
0 34610 5 1 1 34609
0 34611 7 1 2 72002 34610
0 34612 5 1 1 34611
0 34613 7 1 2 34606 34612
0 34614 7 1 2 34604 34613
0 34615 5 1 1 34614
0 34616 7 1 2 82179 34615
0 34617 5 1 1 34616
0 34618 7 4 2 62694 79047
0 34619 7 1 2 74855 73876
0 34620 7 1 2 93333 34619
0 34621 7 1 2 95101 34620
0 34622 5 1 1 34621
0 34623 7 1 2 34617 34622
0 34624 5 1 1 34623
0 34625 7 1 2 65254 34624
0 34626 5 1 1 34625
0 34627 7 1 2 90247 94884
0 34628 5 1 1 34627
0 34629 7 1 2 95063 34628
0 34630 5 1 1 34629
0 34631 7 1 2 93570 34630
0 34632 5 1 1 34631
0 34633 7 1 2 77299 80872
0 34634 7 1 2 95102 34633
0 34635 7 1 2 95066 34634
0 34636 5 1 1 34635
0 34637 7 1 2 34632 34636
0 34638 5 1 1 34637
0 34639 7 1 2 66549 34638
0 34640 5 1 1 34639
0 34641 7 1 2 34626 34640
0 34642 7 1 2 34591 34641
0 34643 5 1 1 34642
0 34644 7 1 2 86790 34643
0 34645 5 1 1 34644
0 34646 7 3 2 92280 92332
0 34647 5 1 1 95105
0 34648 7 2 2 90631 95106
0 34649 5 1 1 95108
0 34650 7 2 2 77080 92327
0 34651 5 1 1 95110
0 34652 7 1 2 65730 95111
0 34653 5 1 1 34652
0 34654 7 1 2 34649 34653
0 34655 5 1 1 34654
0 34656 7 1 2 64305 34655
0 34657 5 1 1 34656
0 34658 7 1 2 92338 94087
0 34659 5 1 1 34658
0 34660 7 1 2 34651 34659
0 34661 5 1 1 34660
0 34662 7 1 2 62346 34661
0 34663 5 1 1 34662
0 34664 7 1 2 34657 34663
0 34665 5 1 1 34664
0 34666 7 1 2 72003 34665
0 34667 5 1 1 34666
0 34668 7 1 2 89164 95109
0 34669 5 1 1 34668
0 34670 7 1 2 34667 34669
0 34671 5 1 1 34670
0 34672 7 1 2 75610 34671
0 34673 5 1 1 34672
0 34674 7 1 2 69993 94631
0 34675 5 1 1 34674
0 34676 7 1 2 34673 34675
0 34677 5 1 1 34676
0 34678 7 1 2 73793 34677
0 34679 5 1 1 34678
0 34680 7 3 2 66550 87176
0 34681 7 1 2 73840 83226
0 34682 5 1 1 34681
0 34683 7 1 2 65015 77216
0 34684 5 1 1 34683
0 34685 7 1 2 78023 34684
0 34686 5 1 1 34685
0 34687 7 1 2 62347 34686
0 34688 5 1 1 34687
0 34689 7 1 2 34682 34688
0 34690 5 1 1 34689
0 34691 7 1 2 78775 34690
0 34692 5 1 1 34691
0 34693 7 2 2 62695 78109
0 34694 5 1 1 95115
0 34695 7 1 2 83687 89967
0 34696 7 1 2 95116 34695
0 34697 5 1 1 34696
0 34698 7 1 2 34692 34697
0 34699 5 1 1 34698
0 34700 7 1 2 95112 34699
0 34701 5 1 1 34700
0 34702 7 1 2 87593 89933
0 34703 5 1 1 34702
0 34704 7 3 2 61876 62348
0 34705 7 1 2 66044 95117
0 34706 7 1 2 95103 34705
0 34707 5 1 1 34706
0 34708 7 1 2 34703 34707
0 34709 5 1 1 34708
0 34710 7 1 2 86999 34709
0 34711 5 1 1 34710
0 34712 7 1 2 81257 87115
0 34713 7 1 2 95104 34712
0 34714 5 1 1 34713
0 34715 7 1 2 34711 34714
0 34716 7 1 2 34701 34715
0 34717 5 1 1 34716
0 34718 7 1 2 81191 34717
0 34719 5 1 1 34718
0 34720 7 2 2 75225 73841
0 34721 5 1 1 95120
0 34722 7 2 2 64779 93441
0 34723 7 1 2 72449 95122
0 34724 5 1 1 34723
0 34725 7 1 2 34721 34724
0 34726 5 1 1 34725
0 34727 7 1 2 92328 34726
0 34728 5 1 1 34727
0 34729 7 1 2 74131 95098
0 34730 5 1 1 34729
0 34731 7 1 2 72349 79395
0 34732 7 1 2 81869 34731
0 34733 5 1 1 34732
0 34734 7 1 2 34730 34733
0 34735 5 1 1 34734
0 34736 7 1 2 92788 34735
0 34737 5 1 1 34736
0 34738 7 1 2 34728 34737
0 34739 5 1 1 34738
0 34740 7 1 2 71807 34739
0 34741 5 1 1 34740
0 34742 7 1 2 69994 82721
0 34743 7 1 2 92329 34742
0 34744 5 1 1 34743
0 34745 7 1 2 21629 34744
0 34746 5 1 1 34745
0 34747 7 1 2 65255 34746
0 34748 5 1 1 34747
0 34749 7 1 2 86365 92771
0 34750 7 1 2 74837 34749
0 34751 7 1 2 94633 34750
0 34752 5 1 1 34751
0 34753 7 1 2 34748 34752
0 34754 5 1 1 34753
0 34755 7 1 2 66551 34754
0 34756 5 1 1 34755
0 34757 7 1 2 34741 34756
0 34758 7 1 2 34719 34757
0 34759 7 1 2 34679 34758
0 34760 7 1 2 34645 34759
0 34761 5 1 1 34760
0 34762 7 1 2 64105 34761
0 34763 5 1 1 34762
0 34764 7 1 2 69853 81884
0 34765 5 1 1 34764
0 34766 7 1 2 82063 34765
0 34767 5 1 1 34766
0 34768 7 1 2 75689 94206
0 34769 7 1 2 87083 34768
0 34770 7 1 2 94785 34769
0 34771 7 1 2 34767 34770
0 34772 5 1 1 34771
0 34773 7 1 2 34763 34772
0 34774 5 1 1 34773
0 34775 7 1 2 64018 34774
0 34776 5 1 1 34775
0 34777 7 1 2 34535 34776
0 34778 5 2 1 34777
0 34779 7 1 2 79589 95124
0 34780 5 1 1 34779
0 34781 7 1 2 61962 34780
0 34782 7 1 2 34474 34781
0 34783 7 1 2 33490 34782
0 34784 7 1 2 94787 34783
0 34785 5 1 1 34784
0 34786 7 1 2 65664 34785
0 34787 7 1 2 22616 34786
0 34788 5 1 1 34787
0 34789 7 1 2 66943 32618
0 34790 5 1 1 34789
0 34791 7 1 2 66944 94890
0 34792 5 1 1 34791
0 34793 7 2 2 61963 79636
0 34794 7 1 2 86718 87862
0 34795 7 4 2 95126 34794
0 34796 7 1 2 85115 26124
0 34797 5 1 1 34796
0 34798 7 1 2 65256 34797
0 34799 5 1 1 34798
0 34800 7 1 2 70317 93508
0 34801 5 1 1 34800
0 34802 7 1 2 34799 34801
0 34803 5 1 1 34802
0 34804 7 1 2 64306 34803
0 34805 5 1 1 34804
0 34806 7 1 2 86838 93753
0 34807 5 1 1 34806
0 34808 7 1 2 34805 34807
0 34809 5 1 1 34808
0 34810 7 1 2 74159 34809
0 34811 5 1 1 34810
0 34812 7 1 2 62349 78611
0 34813 7 1 2 86049 34812
0 34814 5 1 1 34813
0 34815 7 1 2 93621 34814
0 34816 7 1 2 34811 34815
0 34817 5 1 1 34816
0 34818 7 1 2 64780 34817
0 34819 5 1 1 34818
0 34820 7 1 2 75322 83233
0 34821 5 1 1 34820
0 34822 7 1 2 82375 34821
0 34823 5 1 1 34822
0 34824 7 1 2 88280 94811
0 34825 5 1 1 34824
0 34826 7 1 2 34823 34825
0 34827 5 1 1 34826
0 34828 7 1 2 94569 34827
0 34829 5 1 1 34828
0 34830 7 1 2 69260 77050
0 34831 5 3 1 34830
0 34832 7 1 2 69129 95132
0 34833 5 1 1 34832
0 34834 7 1 2 87529 34833
0 34835 5 1 1 34834
0 34836 7 1 2 34829 34835
0 34837 7 1 2 34819 34836
0 34838 5 1 1 34837
0 34839 7 1 2 63507 34838
0 34840 5 1 1 34839
0 34841 7 2 2 70978 79541
0 34842 7 1 2 78576 94263
0 34843 7 1 2 95135 34842
0 34844 5 1 1 34843
0 34845 7 1 2 34840 34844
0 34846 5 1 1 34845
0 34847 7 1 2 95128 34846
0 34848 5 1 1 34847
0 34849 7 1 2 34792 34848
0 34850 5 1 1 34849
0 34851 7 1 2 64106 34850
0 34852 5 1 1 34851
0 34853 7 1 2 66945 94894
0 34854 5 1 1 34853
0 34855 7 1 2 34852 34854
0 34856 5 1 1 34855
0 34857 7 1 2 73842 34856
0 34858 5 1 1 34857
0 34859 7 1 2 66946 95076
0 34860 5 1 1 34859
0 34861 7 1 2 70887 11968
0 34862 5 1 1 34861
0 34863 7 1 2 69261 34862
0 34864 5 1 1 34863
0 34865 7 1 2 80590 86939
0 34866 5 1 1 34865
0 34867 7 1 2 81574 34866
0 34868 5 1 1 34867
0 34869 7 1 2 34864 34868
0 34870 5 1 1 34869
0 34871 7 1 2 70318 34870
0 34872 5 1 1 34871
0 34873 7 1 2 3728 87478
0 34874 5 1 1 34873
0 34875 7 1 2 69262 73279
0 34876 7 1 2 34874 34875
0 34877 5 1 1 34876
0 34878 7 1 2 68032 90864
0 34879 5 2 1 34878
0 34880 7 1 2 70817 95137
0 34881 5 1 1 34880
0 34882 7 1 2 81575 82789
0 34883 7 1 2 87480 34882
0 34884 5 1 1 34883
0 34885 7 1 2 70190 34884
0 34886 7 1 2 34881 34885
0 34887 7 1 2 34877 34886
0 34888 7 1 2 34872 34887
0 34889 5 1 1 34888
0 34890 7 1 2 75226 34889
0 34891 5 1 1 34890
0 34892 7 1 2 81838 88463
0 34893 5 1 1 34892
0 34894 7 1 2 81890 34893
0 34895 5 1 1 34894
0 34896 7 2 2 70062 34895
0 34897 7 1 2 86839 95139
0 34898 5 1 1 34897
0 34899 7 1 2 34891 34898
0 34900 5 1 1 34899
0 34901 7 1 2 63508 34900
0 34902 5 1 1 34901
0 34903 7 1 2 84040 88487
0 34904 5 1 1 34903
0 34905 7 1 2 64781 34904
0 34906 5 1 1 34905
0 34907 7 1 2 74473 34906
0 34908 5 1 1 34907
0 34909 7 1 2 78577 87659
0 34910 7 1 2 34908 34909
0 34911 5 1 1 34910
0 34912 7 1 2 34902 34911
0 34913 5 1 1 34912
0 34914 7 1 2 95129 34913
0 34915 5 1 1 34914
0 34916 7 1 2 34860 34915
0 34917 5 1 1 34916
0 34918 7 1 2 64107 34917
0 34919 5 1 1 34918
0 34920 7 1 2 66947 95080
0 34921 5 1 1 34920
0 34922 7 1 2 34919 34921
0 34923 5 1 1 34922
0 34924 7 1 2 71923 34923
0 34925 5 1 1 34924
0 34926 7 1 2 66948 95125
0 34927 5 1 1 34926
0 34928 7 1 2 91020 95123
0 34929 5 1 1 34928
0 34930 7 1 2 88391 95121
0 34931 5 1 1 34930
0 34932 7 1 2 34929 34931
0 34933 5 1 1 34932
0 34934 7 5 2 63509 64108
0 34935 7 1 2 95130 95141
0 34936 7 1 2 34933 34935
0 34937 5 1 1 34936
0 34938 7 1 2 34927 34937
0 34939 5 1 1 34938
0 34940 7 1 2 79590 34939
0 34941 5 1 1 34940
0 34942 7 1 2 86050 93214
0 34943 5 1 1 34942
0 34944 7 1 2 17679 34943
0 34945 5 1 1 34944
0 34946 7 1 2 88392 34945
0 34947 5 1 1 34946
0 34948 7 1 2 66326 94836
0 34949 5 1 1 34948
0 34950 7 1 2 32911 34949
0 34951 5 1 1 34950
0 34952 7 1 2 69686 34951
0 34953 5 1 1 34952
0 34954 7 1 2 94023 34953
0 34955 5 1 1 34954
0 34956 7 1 2 93442 34955
0 34957 5 1 1 34956
0 34958 7 1 2 81829 75813
0 34959 5 1 1 34958
0 34960 7 1 2 73794 34959
0 34961 5 1 1 34960
0 34962 7 1 2 78602 34961
0 34963 5 1 1 34962
0 34964 7 1 2 87660 34963
0 34965 5 1 1 34964
0 34966 7 1 2 34957 34965
0 34967 7 1 2 34947 34966
0 34968 5 1 1 34967
0 34969 7 1 2 63510 34968
0 34970 5 1 1 34969
0 34971 7 1 2 69687 79846
0 34972 5 3 1 34971
0 34973 7 1 2 90372 95146
0 34974 5 1 1 34973
0 34975 7 1 2 73795 34974
0 34976 5 1 1 34975
0 34977 7 1 2 76709 82145
0 34978 5 1 1 34977
0 34979 7 1 2 64552 34978
0 34980 5 1 1 34979
0 34981 7 1 2 90650 34980
0 34982 5 1 1 34981
0 34983 7 1 2 69688 34982
0 34984 5 1 1 34983
0 34985 7 1 2 82095 74752
0 34986 5 1 1 34985
0 34987 7 1 2 62696 34986
0 34988 5 1 1 34987
0 34989 7 1 2 34984 34988
0 34990 5 1 1 34989
0 34991 7 1 2 70496 34990
0 34992 5 1 1 34991
0 34993 7 1 2 34976 34992
0 34994 5 1 1 34993
0 34995 7 1 2 66327 34994
0 34996 5 1 1 34995
0 34997 7 1 2 17379 34996
0 34998 5 1 1 34997
0 34999 7 1 2 63073 34998
0 35000 5 1 1 34999
0 35001 7 2 2 77300 82113
0 35002 5 1 1 95149
0 35003 7 2 2 74530 95150
0 35004 7 1 2 73877 95151
0 35005 5 1 1 35004
0 35006 7 1 2 35000 35005
0 35007 5 1 1 35006
0 35008 7 1 2 65016 35007
0 35009 5 1 1 35008
0 35010 7 1 2 77715 93488
0 35011 7 1 2 80609 35010
0 35012 5 1 1 35011
0 35013 7 1 2 35009 35012
0 35014 5 1 1 35013
0 35015 7 1 2 75227 35014
0 35016 5 1 1 35015
0 35017 7 1 2 34970 35016
0 35018 5 1 1 35017
0 35019 7 1 2 64109 95131
0 35020 7 1 2 35018 35019
0 35021 5 1 1 35020
0 35022 7 1 2 34941 35021
0 35023 7 1 2 34925 35022
0 35024 7 1 2 34858 35023
0 35025 7 1 2 34790 35024
0 35026 5 1 1 35025
0 35027 7 1 2 60749 35026
0 35028 5 1 1 35027
0 35029 7 2 2 407 78689
0 35030 5 5 1 95153
0 35031 7 1 2 62136 83227
0 35032 5 1 1 35031
0 35033 7 1 2 80224 35032
0 35034 5 1 1 35033
0 35035 7 1 2 62697 35034
0 35036 5 1 1 35035
0 35037 7 1 2 82681 94501
0 35038 5 1 1 35037
0 35039 7 1 2 61077 35038
0 35040 7 1 2 35036 35039
0 35041 5 1 1 35040
0 35042 7 1 2 67079 80218
0 35043 5 1 1 35042
0 35044 7 1 2 72004 74302
0 35045 5 1 1 35044
0 35046 7 1 2 35043 35045
0 35047 5 1 1 35046
0 35048 7 1 2 67664 35047
0 35049 5 1 1 35048
0 35050 7 1 2 82099 74485
0 35051 5 1 1 35050
0 35052 7 1 2 71496 82075
0 35053 5 1 1 35052
0 35054 7 1 2 35051 35053
0 35055 5 1 1 35054
0 35056 7 1 2 59559 35055
0 35057 5 1 1 35056
0 35058 7 1 2 70954 77278
0 35059 5 1 1 35058
0 35060 7 1 2 59907 35059
0 35061 5 1 1 35060
0 35062 7 1 2 66045 35061
0 35063 7 1 2 35057 35062
0 35064 7 1 2 35049 35063
0 35065 5 1 1 35064
0 35066 7 1 2 35041 35065
0 35067 5 1 1 35066
0 35068 7 3 2 69689 74100
0 35069 5 1 1 95160
0 35070 7 1 2 74713 95161
0 35071 5 1 1 35070
0 35072 7 1 2 35067 35071
0 35073 5 2 1 35072
0 35074 7 1 2 63074 95163
0 35075 5 1 1 35074
0 35076 7 2 2 85573 88509
0 35077 5 1 1 95165
0 35078 7 1 2 35075 35077
0 35079 5 1 1 35078
0 35080 7 1 2 61572 35079
0 35081 5 1 1 35080
0 35082 7 1 2 73446 83999
0 35083 5 1 1 35082
0 35084 7 2 2 369 1764
0 35085 5 1 1 95167
0 35086 7 1 2 64307 59560
0 35087 7 1 2 35085 35086
0 35088 5 1 1 35087
0 35089 7 1 2 35083 35088
0 35090 5 1 1 35089
0 35091 7 1 2 73322 85072
0 35092 7 1 2 35090 35091
0 35093 5 1 1 35092
0 35094 7 1 2 35081 35093
0 35095 5 1 1 35094
0 35096 7 1 2 62350 35095
0 35097 5 1 1 35096
0 35098 7 2 2 74281 75909
0 35099 5 1 1 95169
0 35100 7 1 2 7914 35099
0 35101 5 1 1 35100
0 35102 7 1 2 64553 35101
0 35103 5 1 1 35102
0 35104 7 1 2 66046 94327
0 35105 5 1 1 35104
0 35106 7 1 2 35103 35105
0 35107 5 1 1 35106
0 35108 7 1 2 64308 35107
0 35109 5 1 1 35108
0 35110 7 2 2 67331 73350
0 35111 5 1 1 95171
0 35112 7 2 2 65886 73440
0 35113 5 1 1 95173
0 35114 7 1 2 77243 35113
0 35115 5 1 1 35114
0 35116 7 2 2 67080 35115
0 35117 5 1 1 95175
0 35118 7 1 2 35111 35117
0 35119 5 1 1 35118
0 35120 7 1 2 66047 35119
0 35121 5 1 1 35120
0 35122 7 1 2 35109 35121
0 35123 5 2 1 35122
0 35124 7 1 2 84896 95177
0 35125 5 1 1 35124
0 35126 7 4 2 59342 72232
0 35127 5 1 1 95179
0 35128 7 1 2 69344 82865
0 35129 7 1 2 95180 35128
0 35130 5 1 1 35129
0 35131 7 3 2 64309 70497
0 35132 5 2 1 95183
0 35133 7 1 2 80463 95184
0 35134 5 1 1 35133
0 35135 7 1 2 68033 84457
0 35136 7 1 2 35134 35135
0 35137 5 1 1 35136
0 35138 7 1 2 35130 35137
0 35139 5 1 1 35138
0 35140 7 1 2 59561 35139
0 35141 5 1 1 35140
0 35142 7 1 2 59343 77240
0 35143 7 1 2 71619 78971
0 35144 7 1 2 35142 35143
0 35145 5 1 1 35144
0 35146 7 1 2 35141 35145
0 35147 5 1 1 35146
0 35148 7 1 2 60929 35147
0 35149 5 1 1 35148
0 35150 7 1 2 76044 10797
0 35151 5 1 1 35150
0 35152 7 1 2 87356 89120
0 35153 7 1 2 35151 35152
0 35154 5 1 1 35153
0 35155 7 1 2 35149 35154
0 35156 5 1 1 35155
0 35157 7 1 2 66552 35156
0 35158 5 1 1 35157
0 35159 7 1 2 35125 35158
0 35160 5 1 1 35159
0 35161 7 1 2 67665 35160
0 35162 5 1 1 35161
0 35163 7 1 2 59562 88780
0 35164 5 1 1 35163
0 35165 7 1 2 90252 35164
0 35166 5 1 1 35165
0 35167 7 1 2 67332 35166
0 35168 5 1 1 35167
0 35169 7 1 2 24917 35168
0 35170 5 1 1 35169
0 35171 7 1 2 59344 35170
0 35172 5 1 1 35171
0 35173 7 1 2 70368 69351
0 35174 5 1 1 35173
0 35175 7 1 2 88993 35174
0 35176 5 1 1 35175
0 35177 7 1 2 35172 35176
0 35178 5 1 1 35177
0 35179 7 1 2 82412 35178
0 35180 5 1 1 35179
0 35181 7 1 2 80310 83908
0 35182 5 1 1 35181
0 35183 7 1 2 35180 35182
0 35184 5 1 1 35183
0 35185 7 1 2 59908 35184
0 35186 5 1 1 35185
0 35187 7 2 2 73250 72350
0 35188 5 1 1 95188
0 35189 7 1 2 71603 95189
0 35190 5 1 1 35189
0 35191 7 1 2 81580 83965
0 35192 5 1 1 35191
0 35193 7 2 2 35190 35192
0 35194 7 1 2 61078 91265
0 35195 5 1 1 35194
0 35196 7 1 2 95190 35195
0 35197 5 1 1 35196
0 35198 7 1 2 83909 35197
0 35199 5 1 1 35198
0 35200 7 1 2 35186 35199
0 35201 5 1 1 35200
0 35202 7 1 2 62698 35201
0 35203 5 1 1 35202
0 35204 7 1 2 35162 35203
0 35205 7 1 2 35097 35204
0 35206 5 1 1 35205
0 35207 7 1 2 65257 35206
0 35208 5 1 1 35207
0 35209 7 1 2 62351 95164
0 35210 5 1 1 35209
0 35211 7 1 2 82150 95178
0 35212 5 1 1 35211
0 35213 7 1 2 61079 73311
0 35214 5 1 1 35213
0 35215 7 1 2 59909 70925
0 35216 5 1 1 35215
0 35217 7 1 2 35214 35216
0 35218 5 1 1 35217
0 35219 7 1 2 65887 35218
0 35220 5 1 1 35219
0 35221 7 1 2 95191 35220
0 35222 5 1 1 35221
0 35223 7 1 2 62699 35222
0 35224 5 1 1 35223
0 35225 7 1 2 35212 35224
0 35226 7 1 2 35210 35225
0 35227 5 1 1 35226
0 35228 7 1 2 63075 35227
0 35229 5 1 1 35228
0 35230 7 1 2 62352 95166
0 35231 5 1 1 35230
0 35232 7 1 2 35229 35231
0 35233 5 1 1 35232
0 35234 7 1 2 75880 35233
0 35235 5 1 1 35234
0 35236 7 1 2 35208 35235
0 35237 5 1 1 35236
0 35238 7 1 2 68719 35237
0 35239 5 1 1 35238
0 35240 7 1 2 84458 89843
0 35241 5 1 1 35240
0 35242 7 5 2 60371 74946
0 35243 5 1 1 95192
0 35244 7 1 2 67081 85190
0 35245 7 1 2 95193 35244
0 35246 5 1 1 35245
0 35247 7 1 2 35241 35246
0 35248 5 1 1 35247
0 35249 7 1 2 69929 35248
0 35250 5 1 1 35249
0 35251 7 1 2 83627 93003
0 35252 5 1 1 35251
0 35253 7 2 2 69570 91593
0 35254 5 1 1 95197
0 35255 7 1 2 83845 71924
0 35256 7 1 2 95198 35255
0 35257 5 1 1 35256
0 35258 7 1 2 35252 35257
0 35259 7 1 2 35250 35258
0 35260 5 1 1 35259
0 35261 7 1 2 67333 35260
0 35262 5 1 1 35261
0 35263 7 2 2 73045 83846
0 35264 5 1 1 95199
0 35265 7 1 2 71877 95200
0 35266 5 1 1 35265
0 35267 7 1 2 65258 76120
0 35268 7 1 2 93944 35267
0 35269 5 1 1 35268
0 35270 7 1 2 4651 79208
0 35271 7 1 2 93392 35270
0 35272 5 1 1 35271
0 35273 7 1 2 35269 35272
0 35274 5 1 1 35273
0 35275 7 1 2 59910 35274
0 35276 5 1 1 35275
0 35277 7 1 2 35266 35276
0 35278 7 1 2 35262 35277
0 35279 5 1 1 35278
0 35280 7 1 2 68034 35279
0 35281 5 1 1 35280
0 35282 7 1 2 79068 91896
0 35283 7 1 2 84042 35282
0 35284 5 1 1 35283
0 35285 7 1 2 35281 35284
0 35286 5 1 1 35285
0 35287 7 1 2 72124 35286
0 35288 5 1 1 35287
0 35289 7 1 2 73626 76113
0 35290 5 2 1 35289
0 35291 7 1 2 67082 95201
0 35292 5 1 1 35291
0 35293 7 1 2 19317 35292
0 35294 5 2 1 35293
0 35295 7 1 2 69930 95203
0 35296 5 1 1 35295
0 35297 7 1 2 71925 91601
0 35298 5 1 1 35297
0 35299 7 1 2 59345 73825
0 35300 7 1 2 93005 35299
0 35301 5 1 1 35300
0 35302 7 1 2 35298 35301
0 35303 7 1 2 35296 35302
0 35304 5 1 1 35303
0 35305 7 1 2 74598 35304
0 35306 5 1 1 35305
0 35307 7 1 2 73017 74550
0 35308 5 1 1 35307
0 35309 7 1 2 82669 84034
0 35310 7 1 2 35308 35309
0 35311 5 1 1 35310
0 35312 7 1 2 71878 35311
0 35313 5 1 1 35312
0 35314 7 1 2 35306 35313
0 35315 5 1 1 35314
0 35316 7 1 2 79209 79056
0 35317 7 1 2 35315 35316
0 35318 5 1 1 35317
0 35319 7 1 2 35288 35318
0 35320 7 1 2 35239 35319
0 35321 5 1 1 35320
0 35322 7 1 2 63511 35321
0 35323 5 1 1 35322
0 35324 7 1 2 81238 82446
0 35325 5 1 1 35324
0 35326 7 1 2 79910 84801
0 35327 5 3 1 35326
0 35328 7 1 2 91288 93961
0 35329 5 1 1 35328
0 35330 7 1 2 95205 35329
0 35331 5 1 1 35330
0 35332 7 1 2 69931 35331
0 35333 5 1 1 35332
0 35334 7 2 2 75441 83054
0 35335 7 1 2 61080 95208
0 35336 5 1 1 35335
0 35337 7 1 2 85729 35336
0 35338 5 1 1 35337
0 35339 7 1 2 69571 35338
0 35340 5 1 1 35339
0 35341 7 1 2 84656 88568
0 35342 5 1 1 35341
0 35343 7 1 2 35342 95206
0 35344 5 1 1 35343
0 35345 7 1 2 59563 35344
0 35346 5 1 1 35345
0 35347 7 1 2 35340 35346
0 35348 7 1 2 35333 35347
0 35349 5 1 1 35348
0 35350 7 1 2 83628 35349
0 35351 5 1 1 35350
0 35352 7 1 2 66048 83847
0 35353 7 1 2 85430 35352
0 35354 5 1 1 35353
0 35355 7 1 2 35351 35354
0 35356 5 1 1 35355
0 35357 7 1 2 35325 35356
0 35358 5 1 1 35357
0 35359 7 1 2 75750 86270
0 35360 5 1 1 35359
0 35361 7 1 2 78513 84779
0 35362 7 1 2 80303 35361
0 35363 7 1 2 94573 35362
0 35364 5 1 1 35363
0 35365 7 1 2 35360 35364
0 35366 5 1 1 35365
0 35367 7 1 2 64554 35366
0 35368 5 1 1 35367
0 35369 7 1 2 62353 94978
0 35370 5 1 1 35369
0 35371 7 1 2 71497 79172
0 35372 5 1 1 35371
0 35373 7 1 2 71113 82806
0 35374 5 2 1 35373
0 35375 7 1 2 60930 95210
0 35376 7 1 2 35372 35375
0 35377 7 1 2 35370 35376
0 35378 5 1 1 35377
0 35379 7 1 2 71333 71628
0 35380 7 1 2 12942 35379
0 35381 5 1 1 35380
0 35382 7 1 2 77308 75757
0 35383 7 1 2 91190 35382
0 35384 5 1 1 35383
0 35385 7 1 2 35381 35384
0 35386 7 1 2 35378 35385
0 35387 5 1 1 35386
0 35388 7 1 2 67666 35387
0 35389 5 1 1 35388
0 35390 7 1 2 2491 35389
0 35391 5 1 1 35390
0 35392 7 1 2 79210 35391
0 35393 5 1 1 35392
0 35394 7 1 2 35368 35393
0 35395 5 1 1 35394
0 35396 7 1 2 65259 35395
0 35397 5 1 1 35396
0 35398 7 1 2 71433 88631
0 35399 5 1 1 35398
0 35400 7 1 2 73619 35399
0 35401 5 1 1 35400
0 35402 7 1 2 3544 73796
0 35403 5 1 1 35402
0 35404 7 1 2 80261 71926
0 35405 7 1 2 35403 35404
0 35406 5 1 1 35405
0 35407 7 1 2 35401 35406
0 35408 5 1 1 35407
0 35409 7 1 2 71498 35408
0 35410 5 1 1 35409
0 35411 7 1 2 72125 76121
0 35412 7 1 2 91550 35411
0 35413 5 1 1 35412
0 35414 7 1 2 71727 95202
0 35415 5 1 1 35414
0 35416 7 1 2 69263 71879
0 35417 5 1 1 35416
0 35418 7 1 2 35415 35417
0 35419 7 1 2 35413 35418
0 35420 5 1 1 35419
0 35421 7 1 2 59911 35420
0 35422 5 1 1 35421
0 35423 7 1 2 82151 73329
0 35424 5 1 1 35423
0 35425 7 1 2 66553 35424
0 35426 7 1 2 35422 35425
0 35427 7 1 2 35410 35426
0 35428 5 1 1 35427
0 35429 7 1 2 85662 88464
0 35430 5 1 1 35429
0 35431 7 1 2 79415 86400
0 35432 5 1 1 35431
0 35433 7 1 2 61573 35432
0 35434 7 1 2 35430 35433
0 35435 5 1 1 35434
0 35436 7 1 2 35428 35435
0 35437 5 1 1 35436
0 35438 7 1 2 74739 75751
0 35439 7 1 2 82807 35438
0 35440 5 1 1 35439
0 35441 7 1 2 35437 35440
0 35442 5 1 1 35441
0 35443 7 1 2 83360 35442
0 35444 5 1 1 35443
0 35445 7 1 2 68035 35444
0 35446 7 1 2 35397 35445
0 35447 5 1 1 35446
0 35448 7 1 2 67334 73251
0 35449 5 1 1 35448
0 35450 7 1 2 92976 35449
0 35451 5 1 1 35450
0 35452 7 1 2 65888 35451
0 35453 5 1 1 35452
0 35454 7 1 2 69854 95172
0 35455 5 1 1 35454
0 35456 7 1 2 1565 35455
0 35457 5 1 1 35456
0 35458 7 1 2 82808 35457
0 35459 5 1 1 35458
0 35460 7 1 2 35453 35459
0 35461 5 1 1 35460
0 35462 7 1 2 83629 35461
0 35463 5 1 1 35462
0 35464 7 1 2 35264 35463
0 35465 5 1 1 35464
0 35466 7 1 2 62700 35465
0 35467 5 1 1 35466
0 35468 7 3 2 75910 84153
0 35469 7 1 2 90415 95212
0 35470 5 1 1 35469
0 35471 7 1 2 35467 35470
0 35472 5 1 1 35471
0 35473 7 1 2 84459 35472
0 35474 5 1 1 35473
0 35475 7 1 2 78632 83674
0 35476 5 1 1 35475
0 35477 7 1 2 64782 83630
0 35478 7 1 2 89143 35477
0 35479 5 1 1 35478
0 35480 7 1 2 35476 35479
0 35481 5 1 1 35480
0 35482 7 1 2 69130 35481
0 35483 5 1 1 35482
0 35484 7 1 2 72575 83848
0 35485 5 1 1 35484
0 35486 7 1 2 35483 35485
0 35487 5 1 1 35486
0 35488 7 1 2 62137 35487
0 35489 5 1 1 35488
0 35490 7 1 2 75791 76260
0 35491 5 1 1 35490
0 35492 7 1 2 76517 35491
0 35493 5 2 1 35492
0 35494 7 1 2 93946 95215
0 35495 5 1 1 35494
0 35496 7 1 2 66049 35495
0 35497 7 1 2 35489 35496
0 35498 5 1 1 35497
0 35499 7 1 2 72005 80794
0 35500 7 2 2 89777 35499
0 35501 5 1 1 95217
0 35502 7 1 2 64310 95218
0 35503 5 1 1 35502
0 35504 7 1 2 83679 35503
0 35505 5 1 1 35504
0 35506 7 1 2 1744 35505
0 35507 5 1 1 35506
0 35508 7 1 2 83849 94010
0 35509 5 1 1 35508
0 35510 7 1 2 64311 83850
0 35511 5 1 1 35510
0 35512 7 1 2 35501 35511
0 35513 5 1 1 35512
0 35514 7 1 2 69369 35513
0 35515 5 1 1 35514
0 35516 7 1 2 35509 35515
0 35517 7 1 2 35507 35516
0 35518 5 1 1 35517
0 35519 7 1 2 62354 35518
0 35520 5 1 1 35519
0 35521 7 1 2 62138 83675
0 35522 7 1 2 80610 35521
0 35523 5 1 1 35522
0 35524 7 1 2 61081 35523
0 35525 7 1 2 35520 35524
0 35526 5 1 1 35525
0 35527 7 1 2 35498 35526
0 35528 5 1 1 35527
0 35529 7 2 2 73018 80219
0 35530 5 1 1 95219
0 35531 7 1 2 83851 95220
0 35532 5 1 1 35531
0 35533 7 1 2 62701 35532
0 35534 7 1 2 35528 35533
0 35535 5 1 1 35534
0 35536 7 1 2 79999 80445
0 35537 5 1 1 35536
0 35538 7 1 2 72634 94400
0 35539 5 1 1 35538
0 35540 7 2 2 35537 35539
0 35541 7 1 2 73046 88360
0 35542 5 1 1 35541
0 35543 7 1 2 77301 79148
0 35544 5 1 1 35543
0 35545 7 1 2 35542 35544
0 35546 7 1 2 95221 35545
0 35547 5 1 1 35546
0 35548 7 1 2 75498 35547
0 35549 5 1 1 35548
0 35550 7 1 2 79333 88921
0 35551 7 1 2 88671 35550
0 35552 5 1 1 35551
0 35553 7 1 2 35549 35552
0 35554 5 1 1 35553
0 35555 7 1 2 63788 35554
0 35556 5 1 1 35555
0 35557 7 1 2 67335 84154
0 35558 7 1 2 78994 35557
0 35559 7 1 2 95136 35558
0 35560 5 1 1 35559
0 35561 7 1 2 67667 35560
0 35562 7 1 2 35556 35561
0 35563 5 1 1 35562
0 35564 7 1 2 35535 35563
0 35565 5 1 1 35564
0 35566 7 1 2 63076 35565
0 35567 7 1 2 35474 35566
0 35568 5 1 1 35567
0 35569 7 1 2 68404 35568
0 35570 7 1 2 35447 35569
0 35571 5 1 1 35570
0 35572 7 1 2 35358 35571
0 35573 7 1 2 35323 35572
0 35574 5 1 1 35573
0 35575 7 4 2 65665 66949
0 35576 5 1 1 95223
0 35577 7 6 2 68979 95224
0 35578 7 1 2 94478 95227
0 35579 7 1 2 35574 35578
0 35580 5 1 1 35579
0 35581 7 1 2 67668 76940
0 35582 5 1 1 35581
0 35583 7 1 2 84941 35582
0 35584 5 1 1 35583
0 35585 7 2 2 77910 35584
0 35586 5 1 1 95233
0 35587 7 1 2 73551 95147
0 35588 5 1 1 35587
0 35589 7 1 2 77302 81539
0 35590 7 1 2 35588 35589
0 35591 5 1 1 35590
0 35592 7 1 2 35586 35591
0 35593 5 1 1 35592
0 35594 7 1 2 75228 35593
0 35595 5 1 1 35594
0 35596 7 1 2 82090 90755
0 35597 5 1 1 35596
0 35598 7 1 2 82515 35597
0 35599 5 1 1 35598
0 35600 7 1 2 3453 35599
0 35601 5 1 1 35600
0 35602 7 1 2 88943 35601
0 35603 5 1 1 35602
0 35604 7 1 2 35595 35603
0 35605 5 1 1 35604
0 35606 7 3 2 66950 68980
0 35607 7 1 2 35605 95235
0 35608 5 1 1 35607
0 35609 7 2 2 82413 95142
0 35610 7 1 2 61964 95238
0 35611 5 1 1 35610
0 35612 7 1 2 35608 35611
0 35613 5 1 1 35612
0 35614 7 1 2 65666 35613
0 35615 5 1 1 35614
0 35616 7 2 2 60750 66951
0 35617 7 1 2 95240 95239
0 35618 5 1 1 35617
0 35619 7 1 2 68720 35618
0 35620 7 1 2 35615 35619
0 35621 5 1 1 35620
0 35622 7 4 2 61082 78259
0 35623 5 3 1 95242
0 35624 7 1 2 79334 95243
0 35625 5 1 1 35624
0 35626 7 1 2 83910 90486
0 35627 5 1 1 35626
0 35628 7 1 2 35625 35627
0 35629 5 1 1 35628
0 35630 7 1 2 68405 35629
0 35631 5 1 1 35630
0 35632 7 1 2 82347 89835
0 35633 5 1 1 35632
0 35634 7 1 2 35631 35633
0 35635 5 1 1 35634
0 35636 7 1 2 95228 35635
0 35637 5 1 1 35636
0 35638 7 1 2 63789 35637
0 35639 5 1 1 35638
0 35640 7 1 2 87509 35639
0 35641 7 1 2 35621 35640
0 35642 5 1 1 35641
0 35643 7 7 2 61877 66952
0 35644 7 2 2 88085 95249
0 35645 7 7 2 65667 92355
0 35646 7 1 2 89778 95143
0 35647 7 1 2 95258 35646
0 35648 7 1 2 95256 35647
0 35649 5 1 1 35648
0 35650 7 1 2 35642 35649
0 35651 5 1 1 35650
0 35652 7 1 2 64019 35651
0 35653 5 1 1 35652
0 35654 7 1 2 75499 95234
0 35655 5 1 1 35654
0 35656 7 1 2 81454 84122
0 35657 5 1 1 35656
0 35658 7 1 2 67669 35657
0 35659 5 1 1 35658
0 35660 7 1 2 67670 78024
0 35661 5 1 1 35660
0 35662 7 2 2 59346 76069
0 35663 5 1 1 95265
0 35664 7 2 2 70369 82790
0 35665 7 2 2 35663 95267
0 35666 7 1 2 74569 95269
0 35667 5 1 1 35666
0 35668 7 1 2 67336 35667
0 35669 5 1 1 35668
0 35670 7 1 2 35661 35669
0 35671 5 1 1 35670
0 35672 7 1 2 61083 35671
0 35673 5 1 1 35672
0 35674 7 1 2 75611 35673
0 35675 7 1 2 35659 35674
0 35676 5 1 1 35675
0 35677 7 1 2 59912 91187
0 35678 7 1 2 95148 35677
0 35679 5 1 1 35678
0 35680 7 1 2 92177 35679
0 35681 5 1 1 35680
0 35682 7 1 2 91085 94866
0 35683 7 1 2 35681 35682
0 35684 5 1 1 35683
0 35685 7 1 2 66050 35684
0 35686 5 1 1 35685
0 35687 7 1 2 72518 91471
0 35688 5 1 1 35687
0 35689 7 1 2 77476 35688
0 35690 5 1 1 35689
0 35691 7 1 2 75500 35690
0 35692 7 1 2 35686 35691
0 35693 5 1 1 35692
0 35694 7 1 2 75384 86844
0 35695 7 1 2 35693 35694
0 35696 7 1 2 35676 35695
0 35697 5 1 1 35696
0 35698 7 1 2 35655 35697
0 35699 5 1 1 35698
0 35700 7 1 2 88143 35699
0 35701 5 1 1 35700
0 35702 7 1 2 75849 71373
0 35703 5 1 1 35702
0 35704 7 1 2 83163 35703
0 35705 5 1 1 35704
0 35706 7 1 2 63077 35705
0 35707 5 1 1 35706
0 35708 7 1 2 75442 85073
0 35709 5 1 1 35708
0 35710 7 1 2 35707 35709
0 35711 5 1 1 35710
0 35712 7 1 2 65260 35711
0 35713 5 1 1 35712
0 35714 7 1 2 75881 84879
0 35715 5 1 1 35714
0 35716 7 1 2 35713 35715
0 35717 5 1 1 35716
0 35718 7 1 2 87402 35717
0 35719 5 1 1 35718
0 35720 7 1 2 74599 95204
0 35721 5 1 1 35720
0 35722 7 1 2 74289 17786
0 35723 5 1 1 35722
0 35724 7 1 2 85120 35723
0 35725 5 1 1 35724
0 35726 7 1 2 35721 35725
0 35727 5 1 1 35726
0 35728 7 1 2 77911 35727
0 35729 5 1 1 35728
0 35730 7 2 2 62702 93074
0 35731 7 1 2 90151 95271
0 35732 5 1 1 35731
0 35733 7 1 2 35729 35732
0 35734 5 1 1 35733
0 35735 7 1 2 69932 35734
0 35736 5 1 1 35735
0 35737 7 1 2 71808 81427
0 35738 5 3 1 35737
0 35739 7 1 2 61084 82327
0 35740 7 1 2 95273 35739
0 35741 5 1 1 35740
0 35742 7 1 2 67083 95216
0 35743 5 1 1 35742
0 35744 7 1 2 66051 7305
0 35745 7 1 2 35743 35744
0 35746 5 1 1 35745
0 35747 7 1 2 35741 35746
0 35748 5 1 1 35747
0 35749 7 1 2 62703 35530
0 35750 7 1 2 35748 35749
0 35751 5 1 1 35750
0 35752 7 1 2 77217 82630
0 35753 5 1 1 35752
0 35754 7 1 2 67671 35753
0 35755 7 1 2 95222 35754
0 35756 5 1 1 35755
0 35757 7 1 2 77789 35756
0 35758 7 1 2 35751 35757
0 35759 5 1 1 35758
0 35760 7 1 2 35736 35759
0 35761 7 1 2 77807 88361
0 35762 5 1 1 35761
0 35763 7 1 2 77940 88366
0 35764 5 1 1 35763
0 35765 7 1 2 67672 35764
0 35766 7 1 2 35762 35765
0 35767 5 1 1 35766
0 35768 7 1 2 71225 85945
0 35769 7 1 2 78659 35768
0 35770 5 1 1 35769
0 35771 7 1 2 35767 35770
0 35772 5 1 1 35771
0 35773 7 1 2 73047 35772
0 35774 5 1 1 35773
0 35775 7 2 2 64783 90925
0 35776 7 1 2 90723 95276
0 35777 5 1 1 35776
0 35778 7 1 2 73019 1341
0 35779 7 1 2 88562 35778
0 35780 5 1 1 35779
0 35781 7 1 2 67337 84673
0 35782 5 1 1 35781
0 35783 7 1 2 81936 35782
0 35784 5 1 1 35783
0 35785 7 1 2 74624 35784
0 35786 5 1 1 35785
0 35787 7 1 2 67673 35786
0 35788 7 1 2 35780 35787
0 35789 5 1 1 35788
0 35790 7 1 2 84056 93033
0 35791 7 1 2 35789 35790
0 35792 5 1 1 35791
0 35793 7 1 2 35777 35792
0 35794 5 1 1 35793
0 35795 7 1 2 68036 35794
0 35796 5 1 1 35795
0 35797 7 1 2 35774 35796
0 35798 7 1 2 35760 35797
0 35799 5 1 1 35798
0 35800 7 1 2 66554 35799
0 35801 5 1 1 35800
0 35802 7 1 2 79310 35801
0 35803 5 1 1 35802
0 35804 7 1 2 78640 79166
0 35805 5 1 1 35804
0 35806 7 1 2 62139 77262
0 35807 5 1 1 35806
0 35808 7 1 2 67084 88758
0 35809 5 2 1 35808
0 35810 7 1 2 35807 95278
0 35811 5 1 1 35810
0 35812 7 1 2 62704 35811
0 35813 5 1 1 35812
0 35814 7 1 2 35805 35813
0 35815 5 1 1 35814
0 35816 7 1 2 62355 35815
0 35817 5 1 1 35816
0 35818 7 2 2 67085 74176
0 35819 5 2 1 95280
0 35820 7 1 2 59913 95282
0 35821 5 1 1 35820
0 35822 7 1 2 89515 35821
0 35823 5 1 1 35822
0 35824 7 1 2 35817 35823
0 35825 5 1 1 35824
0 35826 7 1 2 63078 35825
0 35827 5 1 1 35826
0 35828 7 1 2 67674 78514
0 35829 5 1 1 35828
0 35830 7 1 2 8280 35829
0 35831 5 1 1 35830
0 35832 7 1 2 63079 35831
0 35833 5 1 1 35832
0 35834 7 2 2 61085 72780
0 35835 5 1 1 95284
0 35836 7 1 2 59914 95285
0 35837 5 1 1 35836
0 35838 7 1 2 62356 87366
0 35839 7 1 2 88932 35838
0 35840 7 1 2 35837 35839
0 35841 5 1 1 35840
0 35842 7 1 2 35833 35841
0 35843 5 1 1 35842
0 35844 7 1 2 72599 35843
0 35845 5 1 1 35844
0 35846 7 1 2 78206 84133
0 35847 5 1 1 35846
0 35848 7 1 2 80502 78637
0 35849 5 1 1 35848
0 35850 7 1 2 35847 35849
0 35851 5 1 1 35850
0 35852 7 1 2 78195 83960
0 35853 5 1 1 35852
0 35854 7 1 2 71458 69471
0 35855 7 1 2 87367 91519
0 35856 7 1 2 35854 35855
0 35857 5 1 1 35856
0 35858 7 1 2 35853 35857
0 35859 7 1 2 35851 35858
0 35860 5 1 1 35859
0 35861 7 1 2 66052 35860
0 35862 5 1 1 35861
0 35863 7 1 2 75323 35862
0 35864 7 1 2 35845 35863
0 35865 7 1 2 35827 35864
0 35866 5 1 1 35865
0 35867 7 1 2 75406 88075
0 35868 7 1 2 35866 35867
0 35869 7 1 2 35803 35868
0 35870 5 1 1 35869
0 35871 7 1 2 35719 35870
0 35872 5 1 1 35871
0 35873 7 1 2 63790 35872
0 35874 5 1 1 35873
0 35875 7 1 2 35701 35874
0 35876 5 1 1 35875
0 35877 7 1 2 95229 35876
0 35878 5 1 1 35877
0 35879 7 1 2 78428 92077
0 35880 5 1 1 35879
0 35881 7 1 2 20359 35880
0 35882 5 1 1 35881
0 35883 7 42 2 60751 61965
0 35884 5 1 1 95286
0 35885 7 2 2 35576 35884
0 35886 7 1 2 86719 95328
0 35887 5 1 1 35886
0 35888 7 4 2 60675 65668
0 35889 7 3 2 95250 95330
0 35890 5 1 1 95334
0 35891 7 1 2 35887 35890
0 35892 5 3 1 35891
0 35893 7 1 2 64110 95337
0 35894 7 1 2 35882 35893
0 35895 5 1 1 35894
0 35896 7 1 2 35878 35895
0 35897 5 1 1 35896
0 35898 7 1 2 81192 35897
0 35899 5 1 1 35898
0 35900 7 1 2 35653 35899
0 35901 7 1 2 35580 35900
0 35902 5 1 1 35901
0 35903 7 1 2 95155 35902
0 35904 5 1 1 35903
0 35905 7 1 2 35028 35904
0 35906 7 1 2 34788 35905
0 35907 5 1 1 35906
0 35908 7 1 2 69039 35907
0 35909 5 1 1 35908
0 35910 7 2 2 71311 77912
0 35911 5 2 1 95340
0 35912 7 2 2 85994 86029
0 35913 5 1 1 95344
0 35914 7 1 2 18015 35913
0 35915 5 1 1 35914
0 35916 7 1 2 65731 35915
0 35917 5 1 1 35916
0 35918 7 3 2 63080 86515
0 35919 5 1 1 95346
0 35920 7 1 2 35917 35919
0 35921 5 2 1 35920
0 35922 7 1 2 64312 95349
0 35923 5 1 1 35922
0 35924 7 1 2 65732 95347
0 35925 5 1 1 35924
0 35926 7 1 2 35923 35925
0 35927 5 1 1 35926
0 35928 7 1 2 68406 35927
0 35929 5 1 1 35928
0 35930 7 1 2 95342 35929
0 35931 5 1 1 35930
0 35932 7 1 2 72006 35931
0 35933 5 1 1 35932
0 35934 7 2 2 87772 89526
0 35935 7 1 2 68407 95351
0 35936 5 1 1 35935
0 35937 7 1 2 35933 35936
0 35938 5 1 1 35937
0 35939 7 1 2 66053 35938
0 35940 5 1 1 35939
0 35941 7 1 2 93095 95027
0 35942 5 1 1 35941
0 35943 7 1 2 35940 35942
0 35944 5 1 1 35943
0 35945 7 1 2 64784 35944
0 35946 5 1 1 35945
0 35947 7 1 2 64555 93280
0 35948 5 1 1 35947
0 35949 7 1 2 66054 72845
0 35950 5 1 1 35949
0 35951 7 1 2 35948 35950
0 35952 5 1 1 35951
0 35953 7 1 2 64785 35952
0 35954 5 1 1 35953
0 35955 7 1 2 64556 78821
0 35956 5 1 1 35955
0 35957 7 1 2 35954 35956
0 35958 5 1 1 35957
0 35959 7 1 2 71569 35958
0 35960 5 1 1 35959
0 35961 7 1 2 72233 94580
0 35962 5 2 1 35961
0 35963 7 1 2 76746 95353
0 35964 5 1 1 35963
0 35965 7 1 2 35960 35964
0 35966 5 2 1 35965
0 35967 7 1 2 68408 95355
0 35968 5 1 1 35967
0 35969 7 1 2 60372 88372
0 35970 5 2 1 35969
0 35971 7 1 2 88465 95357
0 35972 5 1 1 35971
0 35973 7 1 2 71809 88580
0 35974 5 1 1 35973
0 35975 7 1 2 68409 35974
0 35976 7 1 2 35972 35975
0 35977 5 1 1 35976
0 35978 7 1 2 72126 89275
0 35979 5 1 1 35978
0 35980 7 1 2 78098 94677
0 35981 7 1 2 35979 35980
0 35982 5 1 1 35981
0 35983 7 1 2 63081 35982
0 35984 7 1 2 35977 35983
0 35985 5 1 1 35984
0 35986 7 2 2 73208 72494
0 35987 5 1 1 95359
0 35988 7 1 2 77678 35987
0 35989 7 1 2 88749 35988
0 35990 5 1 1 35989
0 35991 7 1 2 77913 35990
0 35992 5 1 1 35991
0 35993 7 1 2 35985 35992
0 35994 7 1 2 35968 35993
0 35995 5 1 1 35994
0 35996 7 1 2 62705 35995
0 35997 5 1 1 35996
0 35998 7 1 2 81870 90344
0 35999 5 2 1 35998
0 36000 7 1 2 95361 95343
0 36001 5 1 1 36000
0 36002 7 1 2 70818 36001
0 36003 5 1 1 36002
0 36004 7 1 2 71570 74225
0 36005 5 1 1 36004
0 36006 7 1 2 73964 36005
0 36007 5 1 1 36006
0 36008 7 1 2 69690 36007
0 36009 5 1 1 36008
0 36010 7 1 2 69855 88541
0 36011 5 1 1 36010
0 36012 7 1 2 79944 36011
0 36013 7 1 2 36009 36012
0 36014 5 1 1 36013
0 36015 7 1 2 63082 36014
0 36016 5 1 1 36015
0 36017 7 1 2 36003 36016
0 36018 5 1 1 36017
0 36019 7 1 2 78660 36018
0 36020 5 1 1 36019
0 36021 7 1 2 73209 75073
0 36022 5 1 1 36021
0 36023 7 1 2 77941 36022
0 36024 5 1 1 36023
0 36025 7 1 2 70819 36024
0 36026 5 2 1 36025
0 36027 7 1 2 73965 12810
0 36028 5 1 1 36027
0 36029 7 1 2 63083 36028
0 36030 5 1 1 36029
0 36031 7 1 2 95363 36030
0 36032 5 1 1 36031
0 36033 7 1 2 72351 36032
0 36034 5 1 1 36033
0 36035 7 2 2 72676 82931
0 36036 5 1 1 95365
0 36037 7 1 2 63512 79498
0 36038 7 1 2 73228 36037
0 36039 7 1 2 36036 36038
0 36040 5 1 1 36039
0 36041 7 1 2 36034 36040
0 36042 5 1 1 36041
0 36043 7 1 2 71810 36042
0 36044 5 1 1 36043
0 36045 7 1 2 70926 88572
0 36046 5 1 1 36045
0 36047 7 1 2 90097 36046
0 36048 5 1 1 36047
0 36049 7 1 2 75074 36048
0 36050 5 1 1 36049
0 36051 7 1 2 36044 36050
0 36052 7 1 2 36020 36051
0 36053 7 1 2 35997 36052
0 36054 7 1 2 35946 36053
0 36055 5 1 1 36054
0 36056 7 1 2 62357 36055
0 36057 5 1 1 36056
0 36058 7 1 2 62706 90564
0 36059 5 1 1 36058
0 36060 7 1 2 90959 36059
0 36061 5 1 1 36060
0 36062 7 1 2 69264 36061
0 36063 5 1 1 36062
0 36064 7 2 2 82653 82232
0 36065 5 1 1 95367
0 36066 7 1 2 81913 95368
0 36067 5 2 1 36066
0 36068 7 1 2 63084 95369
0 36069 5 1 1 36068
0 36070 7 1 2 73020 95244
0 36071 7 1 2 82091 36070
0 36072 5 1 1 36071
0 36073 7 1 2 66328 36072
0 36074 5 1 1 36073
0 36075 7 1 2 90553 88658
0 36076 5 1 1 36075
0 36077 7 1 2 73380 91262
0 36078 5 1 1 36077
0 36079 7 1 2 69158 36078
0 36080 5 1 1 36079
0 36081 7 1 2 36076 36080
0 36082 7 1 2 36074 36081
0 36083 7 1 2 36069 36082
0 36084 7 1 2 76366 90532
0 36085 5 1 1 36084
0 36086 7 1 2 90562 36085
0 36087 7 1 2 36083 36086
0 36088 7 1 2 36063 36087
0 36089 5 1 1 36088
0 36090 7 1 2 65017 36089
0 36091 5 1 1 36090
0 36092 7 1 2 2936 83333
0 36093 7 1 2 83291 36092
0 36094 5 1 1 36093
0 36095 7 1 2 66329 36094
0 36096 5 1 1 36095
0 36097 7 1 2 23901 36096
0 36098 5 1 1 36097
0 36099 7 1 2 35835 36098
0 36100 5 1 1 36099
0 36101 7 1 2 73112 1086
0 36102 5 1 1 36101
0 36103 7 1 2 94029 36102
0 36104 5 1 1 36103
0 36105 7 1 2 64313 36104
0 36106 5 1 1 36105
0 36107 7 1 2 94115 36106
0 36108 5 1 1 36107
0 36109 7 1 2 88653 36108
0 36110 5 1 1 36109
0 36111 7 1 2 76876 17812
0 36112 5 1 1 36111
0 36113 7 1 2 87467 36112
0 36114 5 1 1 36113
0 36115 7 1 2 74028 88812
0 36116 5 2 1 36115
0 36117 7 1 2 63085 72615
0 36118 5 1 1 36117
0 36119 7 1 2 95371 36118
0 36120 5 1 1 36119
0 36121 7 1 2 64314 36120
0 36122 5 1 1 36121
0 36123 7 1 2 36114 36122
0 36124 5 1 1 36123
0 36125 7 1 2 70370 36124
0 36126 5 1 1 36125
0 36127 7 1 2 36110 36126
0 36128 7 1 2 36100 36127
0 36129 7 1 2 66055 82285
0 36130 5 1 1 36129
0 36131 7 1 2 77309 88551
0 36132 5 1 1 36131
0 36133 7 1 2 64557 36132
0 36134 5 1 1 36133
0 36135 7 1 2 36130 36134
0 36136 5 1 1 36135
0 36137 7 1 2 66330 36136
0 36138 5 1 1 36137
0 36139 7 1 2 71114 88028
0 36140 5 1 1 36139
0 36141 7 1 2 36138 36140
0 36142 5 1 1 36141
0 36143 7 1 2 76367 36142
0 36144 5 1 1 36143
0 36145 7 1 2 86940 93253
0 36146 5 1 1 36145
0 36147 7 1 2 76092 36146
0 36148 5 1 1 36147
0 36149 7 2 2 59915 75913
0 36150 5 1 1 95373
0 36151 7 1 2 62707 36150
0 36152 5 1 1 36151
0 36153 7 1 2 68037 2446
0 36154 7 1 2 36152 36153
0 36155 5 1 1 36154
0 36156 7 1 2 66331 36155
0 36157 5 1 1 36156
0 36158 7 1 2 36148 36157
0 36159 5 1 1 36158
0 36160 7 1 2 74029 36159
0 36161 5 1 1 36160
0 36162 7 2 2 88894 93176
0 36163 7 1 2 90544 95375
0 36164 5 1 1 36163
0 36165 7 1 2 65261 36164
0 36166 5 1 1 36165
0 36167 7 1 2 66332 80079
0 36168 5 1 1 36167
0 36169 7 1 2 59347 36168
0 36170 5 1 1 36169
0 36171 7 1 2 73113 82286
0 36172 5 2 1 36171
0 36173 7 1 2 91453 95377
0 36174 5 1 1 36173
0 36175 7 1 2 61358 90450
0 36176 5 2 1 36175
0 36177 7 1 2 36174 95379
0 36178 7 1 2 36170 36177
0 36179 5 1 1 36178
0 36180 7 1 2 88873 36179
0 36181 7 1 2 36166 36180
0 36182 7 1 2 36161 36181
0 36183 7 1 2 36144 36182
0 36184 7 1 2 36128 36183
0 36185 7 1 2 83136 87282
0 36186 5 1 1 36185
0 36187 7 1 2 66333 36186
0 36188 5 1 1 36187
0 36189 7 1 2 81413 36188
0 36190 5 1 1 36189
0 36191 7 1 2 66056 36190
0 36192 5 1 1 36191
0 36193 7 1 2 83234 36192
0 36194 5 1 1 36193
0 36195 7 1 2 65733 36194
0 36196 5 1 1 36195
0 36197 7 1 2 1803 70930
0 36198 5 1 1 36197
0 36199 7 1 2 65889 36198
0 36200 5 1 1 36199
0 36201 7 1 2 62358 91441
0 36202 5 1 1 36201
0 36203 7 1 2 36200 36202
0 36204 5 1 1 36203
0 36205 7 1 2 70319 36204
0 36206 5 1 1 36205
0 36207 7 1 2 66057 69352
0 36208 5 1 1 36207
0 36209 7 1 2 73915 36208
0 36210 7 1 2 88384 36209
0 36211 5 1 1 36210
0 36212 7 1 2 90518 36211
0 36213 5 1 1 36212
0 36214 7 1 2 79419 36213
0 36215 7 1 2 36206 36214
0 36216 5 1 1 36215
0 36217 7 1 2 63086 36216
0 36218 5 1 1 36217
0 36219 7 1 2 36196 36218
0 36220 7 1 2 36184 36219
0 36221 7 1 2 36091 36220
0 36222 5 2 1 36221
0 36223 7 1 2 68410 95381
0 36224 5 2 1 36223
0 36225 7 1 2 69933 76098
0 36226 5 1 1 36225
0 36227 7 1 2 72007 36226
0 36228 5 1 1 36227
0 36229 7 1 2 88864 36228
0 36230 5 1 1 36229
0 36231 7 1 2 71115 36230
0 36232 5 1 1 36231
0 36233 7 1 2 76679 36232
0 36234 5 1 1 36233
0 36235 7 1 2 74070 79125
0 36236 7 1 2 36234 36235
0 36237 5 1 1 36236
0 36238 7 1 2 63513 36237
0 36239 5 1 1 36238
0 36240 7 1 2 95383 36239
0 36241 5 1 1 36240
0 36242 7 1 2 66555 36241
0 36243 5 1 1 36242
0 36244 7 1 2 71571 28961
0 36245 5 1 1 36244
0 36246 7 1 2 87028 88489
0 36247 5 1 1 36246
0 36248 7 1 2 36245 36247
0 36249 5 1 1 36248
0 36250 7 1 2 68411 36249
0 36251 5 1 1 36250
0 36252 7 1 2 67675 89460
0 36253 5 2 1 36252
0 36254 7 1 2 36251 95385
0 36255 5 1 1 36254
0 36256 7 1 2 71116 36255
0 36257 5 1 1 36256
0 36258 7 2 2 71811 71572
0 36259 7 1 2 88858 95387
0 36260 5 1 1 36259
0 36261 7 1 2 76784 36260
0 36262 5 1 1 36261
0 36263 7 1 2 68412 36262
0 36264 5 1 1 36263
0 36265 7 1 2 79791 88859
0 36266 5 1 1 36265
0 36267 7 1 2 36264 36266
0 36268 5 1 1 36267
0 36269 7 1 2 70320 36268
0 36270 5 1 1 36269
0 36271 7 1 2 59348 89589
0 36272 5 1 1 36271
0 36273 7 1 2 75075 36272
0 36274 5 1 1 36273
0 36275 7 1 2 79818 36274
0 36276 5 1 1 36275
0 36277 7 1 2 70820 36276
0 36278 5 1 1 36277
0 36279 7 1 2 79792 94575
0 36280 5 1 1 36279
0 36281 7 2 2 71812 69370
0 36282 7 1 2 88542 95389
0 36283 5 1 1 36282
0 36284 7 1 2 36280 36283
0 36285 5 1 1 36284
0 36286 7 1 2 62708 36285
0 36287 5 1 1 36286
0 36288 7 1 2 85003 36287
0 36289 7 1 2 36278 36288
0 36290 7 1 2 36270 36289
0 36291 7 1 2 36257 36290
0 36292 5 1 1 36291
0 36293 7 1 2 63087 36292
0 36294 5 1 1 36293
0 36295 7 1 2 79974 77914
0 36296 5 1 1 36295
0 36297 7 1 2 73210 79225
0 36298 5 1 1 36297
0 36299 7 1 2 76785 36298
0 36300 5 1 1 36299
0 36301 7 1 2 68413 36300
0 36302 5 1 1 36301
0 36303 7 1 2 36296 36302
0 36304 5 1 1 36303
0 36305 7 1 2 71117 36304
0 36306 5 1 1 36305
0 36307 7 1 2 77942 95362
0 36308 5 1 1 36307
0 36309 7 1 2 36308 95360
0 36310 5 1 1 36309
0 36311 7 1 2 74226 77707
0 36312 7 1 2 82584 36311
0 36313 5 1 1 36312
0 36314 7 1 2 36310 36313
0 36315 5 1 1 36314
0 36316 7 1 2 71813 36315
0 36317 5 1 1 36316
0 36318 7 1 2 85004 85963
0 36319 7 1 2 36317 36318
0 36320 7 1 2 36306 36319
0 36321 5 1 1 36320
0 36322 7 1 2 62709 36321
0 36323 5 1 1 36322
0 36324 7 1 2 90970 17739
0 36325 5 1 1 36324
0 36326 7 1 2 65262 36325
0 36327 5 1 1 36326
0 36328 7 1 2 80661 85108
0 36329 5 1 1 36328
0 36330 7 1 2 36327 36329
0 36331 5 1 1 36330
0 36332 7 1 2 71814 36331
0 36333 5 1 1 36332
0 36334 7 3 2 63088 69691
0 36335 5 1 1 95391
0 36336 7 1 2 71291 36335
0 36337 5 1 1 36336
0 36338 7 1 2 72008 36337
0 36339 7 1 2 95352 36338
0 36340 5 1 1 36339
0 36341 7 1 2 76747 83032
0 36342 5 2 1 36341
0 36343 7 1 2 68414 95394
0 36344 7 1 2 36340 36343
0 36345 7 1 2 36333 36344
0 36346 5 1 1 36345
0 36347 7 1 2 63089 95162
0 36348 5 2 1 36347
0 36349 7 1 2 68038 94047
0 36350 5 1 1 36349
0 36351 7 2 2 95396 36350
0 36352 5 1 1 95398
0 36353 7 1 2 71459 87732
0 36354 5 1 1 36353
0 36355 7 1 2 85235 36354
0 36356 7 1 2 95399 36355
0 36357 5 1 1 36356
0 36358 7 1 2 71815 36357
0 36359 5 1 1 36358
0 36360 7 1 2 80479 78972
0 36361 5 1 1 36360
0 36362 7 1 2 83921 36361
0 36363 5 1 1 36362
0 36364 7 1 2 62710 36363
0 36365 5 1 1 36364
0 36366 7 1 2 78858 11389
0 36367 5 2 1 36366
0 36368 7 1 2 72009 95400
0 36369 5 2 1 36368
0 36370 7 1 2 63514 95402
0 36371 7 1 2 36365 36370
0 36372 7 1 2 36359 36371
0 36373 5 1 1 36372
0 36374 7 1 2 72352 36373
0 36375 7 1 2 36346 36374
0 36376 5 1 1 36375
0 36377 7 2 2 73229 78211
0 36378 5 1 1 95404
0 36379 7 1 2 63515 95405
0 36380 5 2 1 36379
0 36381 7 1 2 68415 94333
0 36382 5 3 1 36381
0 36383 7 1 2 95364 95408
0 36384 5 1 1 36383
0 36385 7 1 2 62711 36384
0 36386 5 1 1 36385
0 36387 7 1 2 95406 36386
0 36388 5 1 1 36387
0 36389 7 1 2 78661 36388
0 36390 5 1 1 36389
0 36391 7 1 2 75076 88494
0 36392 5 1 1 36391
0 36393 7 1 2 77943 36392
0 36394 5 1 1 36393
0 36395 7 1 2 77740 36394
0 36396 5 1 1 36395
0 36397 7 1 2 90683 36396
0 36398 7 1 2 36390 36397
0 36399 7 1 2 36376 36398
0 36400 7 1 2 36323 36399
0 36401 7 1 2 36294 36400
0 36402 7 1 2 36243 36401
0 36403 7 1 2 36057 36402
0 36404 5 1 1 36403
0 36405 7 1 2 65459 36404
0 36406 5 1 1 36405
0 36407 7 2 2 74311 74269
0 36408 5 1 1 95411
0 36409 7 1 2 78196 36408
0 36410 5 1 1 36409
0 36411 7 1 2 60162 88871
0 36412 5 1 1 36411
0 36413 7 1 2 62359 36412
0 36414 5 1 1 36413
0 36415 7 1 2 12622 36414
0 36416 5 1 1 36415
0 36417 7 1 2 68039 36416
0 36418 5 1 1 36417
0 36419 7 1 2 36410 36418
0 36420 5 2 1 36419
0 36421 7 1 2 75229 95413
0 36422 5 1 1 36421
0 36423 7 3 2 63090 93199
0 36424 7 1 2 76910 90339
0 36425 7 1 2 95415 36424
0 36426 5 1 1 36425
0 36427 7 1 2 36422 36426
0 36428 5 1 1 36427
0 36429 7 1 2 71816 36428
0 36430 5 1 1 36429
0 36431 7 1 2 77477 91089
0 36432 5 1 1 36431
0 36433 7 1 2 91127 93200
0 36434 5 1 1 36433
0 36435 7 1 2 68040 86648
0 36436 5 1 1 36435
0 36437 7 1 2 36434 36436
0 36438 5 1 1 36437
0 36439 7 1 2 70407 36438
0 36440 5 1 1 36439
0 36441 7 1 2 86601 95416
0 36442 5 1 1 36441
0 36443 7 1 2 66556 85558
0 36444 5 1 1 36443
0 36445 7 1 2 36442 36444
0 36446 5 1 1 36445
0 36447 7 1 2 70321 36446
0 36448 5 1 1 36447
0 36449 7 1 2 36440 36448
0 36450 5 1 1 36449
0 36451 7 1 2 62712 36450
0 36452 5 1 1 36451
0 36453 7 1 2 75230 95401
0 36454 5 1 1 36453
0 36455 7 1 2 36452 36454
0 36456 5 1 1 36455
0 36457 7 1 2 72010 36456
0 36458 5 1 1 36457
0 36459 7 1 2 36432 36458
0 36460 7 1 2 36430 36459
0 36461 5 1 1 36460
0 36462 7 1 2 72353 36461
0 36463 5 1 1 36462
0 36464 7 1 2 67676 82328
0 36465 5 3 1 36464
0 36466 7 1 2 71817 95418
0 36467 5 2 1 36466
0 36468 7 1 2 90709 95421
0 36469 5 2 1 36468
0 36470 7 1 2 70063 95423
0 36471 5 1 1 36470
0 36472 7 1 2 74542 90278
0 36473 5 1 1 36472
0 36474 7 1 2 73145 36473
0 36475 5 1 1 36474
0 36476 7 1 2 62140 36475
0 36477 5 1 1 36476
0 36478 7 1 2 83334 78925
0 36479 7 1 2 36477 36478
0 36480 5 1 1 36479
0 36481 7 1 2 79084 36480
0 36482 5 1 1 36481
0 36483 7 1 2 36471 36482
0 36484 5 1 1 36483
0 36485 7 2 2 63091 36484
0 36486 5 1 1 95425
0 36487 7 1 2 85454 95426
0 36488 5 1 1 36487
0 36489 7 1 2 65263 36352
0 36490 5 1 1 36489
0 36491 7 1 2 71573 89874
0 36492 5 1 1 36491
0 36493 7 1 2 88313 36492
0 36494 5 1 1 36493
0 36495 7 1 2 62141 36494
0 36496 5 1 1 36495
0 36497 7 1 2 36490 36496
0 36498 5 1 1 36497
0 36499 7 1 2 62360 36498
0 36500 5 1 1 36499
0 36501 7 3 2 87363 36378
0 36502 5 1 1 95427
0 36503 7 1 2 65264 36502
0 36504 5 1 1 36503
0 36505 7 1 2 36500 36504
0 36506 5 1 1 36505
0 36507 7 1 2 66557 36506
0 36508 5 1 1 36507
0 36509 7 1 2 79107 84950
0 36510 5 1 1 36509
0 36511 7 1 2 36508 36510
0 36512 5 1 1 36511
0 36513 7 1 2 78662 36512
0 36514 5 1 1 36513
0 36515 7 1 2 36488 36514
0 36516 7 1 2 36463 36515
0 36517 7 1 2 72011 77741
0 36518 5 1 1 36517
0 36519 7 1 2 73508 36518
0 36520 5 2 1 36519
0 36521 7 1 2 69692 74291
0 36522 7 3 2 69995 36521
0 36523 7 1 2 95430 95432
0 36524 5 1 1 36523
0 36525 7 2 2 70539 71118
0 36526 5 2 1 95435
0 36527 7 1 2 12546 95412
0 36528 5 1 1 36527
0 36529 7 1 2 72635 36528
0 36530 5 1 1 36529
0 36531 7 1 2 95437 36530
0 36532 5 1 1 36531
0 36533 7 1 2 70064 36532
0 36534 5 1 1 36533
0 36535 7 1 2 36524 36534
0 36536 5 1 1 36535
0 36537 7 1 2 78197 36536
0 36538 5 1 1 36537
0 36539 7 1 2 87377 12806
0 36540 5 1 1 36539
0 36541 7 1 2 36538 36540
0 36542 5 1 1 36541
0 36543 7 1 2 75612 36542
0 36544 5 2 1 36543
0 36545 7 1 2 87759 88445
0 36546 5 1 1 36545
0 36547 7 4 2 63092 81481
0 36548 5 2 1 95441
0 36549 7 1 2 71119 95445
0 36550 7 1 2 36546 36549
0 36551 5 2 1 36550
0 36552 7 1 2 89875 95419
0 36553 5 1 1 36552
0 36554 7 1 2 82294 87733
0 36555 5 1 1 36554
0 36556 7 1 2 36553 36555
0 36557 5 1 1 36556
0 36558 7 1 2 71818 36557
0 36559 5 1 1 36558
0 36560 7 1 2 62713 70408
0 36561 7 1 2 87481 36560
0 36562 5 1 1 36561
0 36563 7 1 2 90098 36562
0 36564 5 1 1 36563
0 36565 7 1 2 12162 36564
0 36566 5 1 1 36565
0 36567 7 1 2 64315 89876
0 36568 5 1 1 36567
0 36569 7 1 2 87742 36568
0 36570 5 1 1 36569
0 36571 7 1 2 76093 36570
0 36572 5 1 1 36571
0 36573 7 1 2 66558 36572
0 36574 7 1 2 36566 36573
0 36575 7 1 2 36559 36574
0 36576 7 1 2 95447 36575
0 36577 5 1 1 36576
0 36578 7 1 2 61574 36486
0 36579 5 1 1 36578
0 36580 7 1 2 65265 36579
0 36581 7 1 2 36577 36580
0 36582 5 1 1 36581
0 36583 7 1 2 95439 36582
0 36584 7 1 2 36516 36583
0 36585 5 1 1 36584
0 36586 7 1 2 63516 36585
0 36587 5 1 1 36586
0 36588 7 1 2 71927 95078
0 36589 5 1 1 36588
0 36590 7 1 2 69693 94802
0 36591 7 1 2 91227 36590
0 36592 5 1 1 36591
0 36593 7 1 2 78012 36592
0 36594 5 1 1 36593
0 36595 7 1 2 63093 36594
0 36596 5 1 1 36595
0 36597 7 1 2 74177 77846
0 36598 5 1 1 36597
0 36599 7 1 2 73843 78578
0 36600 5 1 1 36599
0 36601 7 1 2 77870 90991
0 36602 5 1 1 36601
0 36603 7 1 2 36600 36602
0 36604 5 1 1 36603
0 36605 7 1 2 80000 36604
0 36606 5 1 1 36605
0 36607 7 1 2 36598 36606
0 36608 7 1 2 36596 36607
0 36609 7 1 2 36589 36608
0 36610 5 1 1 36609
0 36611 7 1 2 62361 36610
0 36612 5 1 1 36611
0 36613 7 1 2 71819 88860
0 36614 5 1 1 36613
0 36615 7 1 2 88367 36614
0 36616 5 1 1 36615
0 36617 7 1 2 63094 36616
0 36618 5 1 1 36617
0 36619 7 1 2 90887 36618
0 36620 5 1 1 36619
0 36621 7 1 2 70322 36620
0 36622 5 1 1 36621
0 36623 7 1 2 64316 91451
0 36624 5 1 1 36623
0 36625 7 1 2 77500 36624
0 36626 5 1 1 36625
0 36627 7 2 2 71820 95268
0 36628 7 1 2 36626 95449
0 36629 5 1 1 36628
0 36630 7 1 2 76030 88424
0 36631 5 1 1 36630
0 36632 7 1 2 88975 36631
0 36633 5 1 1 36632
0 36634 7 1 2 36629 36633
0 36635 7 1 2 36622 36634
0 36636 5 1 1 36635
0 36637 7 1 2 70065 36636
0 36638 5 1 1 36637
0 36639 7 1 2 74885 78933
0 36640 7 1 2 88490 36639
0 36641 5 1 1 36640
0 36642 7 1 2 36638 36641
0 36643 5 1 1 36642
0 36644 7 1 2 70821 36643
0 36645 5 1 1 36644
0 36646 7 1 2 36612 36645
0 36647 5 1 1 36646
0 36648 7 1 2 82516 36647
0 36649 5 2 1 36648
0 36650 7 2 2 36587 95451
0 36651 7 1 2 36406 95453
0 36652 5 1 1 36651
0 36653 7 1 2 66723 36652
0 36654 5 1 1 36653
0 36655 7 1 2 71821 95414
0 36656 5 2 1 36655
0 36657 7 2 2 62714 81428
0 36658 5 2 1 95457
0 36659 7 1 2 70616 95459
0 36660 5 1 1 36659
0 36661 7 1 2 68041 36660
0 36662 5 1 1 36661
0 36663 7 1 2 78859 36662
0 36664 5 1 1 36663
0 36665 7 1 2 72012 36664
0 36666 5 1 1 36665
0 36667 7 1 2 95455 36666
0 36668 5 1 1 36667
0 36669 7 1 2 72354 36668
0 36670 5 2 1 36669
0 36671 7 1 2 71312 87734
0 36672 5 2 1 36671
0 36673 7 1 2 95463 95397
0 36674 5 1 1 36673
0 36675 7 1 2 62362 36674
0 36676 5 1 1 36675
0 36677 7 1 2 95428 36676
0 36678 5 1 1 36677
0 36679 7 1 2 78663 36678
0 36680 5 1 1 36679
0 36681 7 2 2 71822 82295
0 36682 5 1 1 95465
0 36683 7 1 2 70191 95460
0 36684 7 1 2 36682 36683
0 36685 5 1 1 36684
0 36686 7 1 2 87735 36685
0 36687 5 1 1 36686
0 36688 7 1 2 36680 36687
0 36689 7 1 2 95448 36688
0 36690 7 1 2 95461 36689
0 36691 5 1 1 36690
0 36692 7 1 2 75231 36691
0 36693 5 1 1 36692
0 36694 7 1 2 95440 36693
0 36695 5 1 1 36694
0 36696 7 1 2 63517 36695
0 36697 5 1 1 36696
0 36698 7 1 2 95452 36697
0 36699 5 1 1 36698
0 36700 7 1 2 65460 36699
0 36701 5 1 1 36700
0 36702 7 1 2 36654 36701
0 36703 5 1 1 36702
0 36704 7 1 2 60676 36703
0 36705 5 1 1 36704
0 36706 7 1 2 87156 36705
0 36707 5 1 1 36706
0 36708 7 1 2 81222 85769
0 36709 5 1 1 36708
0 36710 7 1 2 63518 92186
0 36711 5 1 1 36710
0 36712 7 1 2 36709 36711
0 36713 5 1 1 36712
0 36714 7 1 2 67086 36713
0 36715 5 1 1 36714
0 36716 7 1 2 75745 86864
0 36717 5 1 1 36716
0 36718 7 1 2 36715 36717
0 36719 5 1 1 36718
0 36720 7 1 2 60807 36719
0 36721 5 1 1 36720
0 36722 7 1 2 81540 82932
0 36723 7 1 2 80708 36722
0 36724 5 1 1 36723
0 36725 7 1 2 36721 36724
0 36726 5 1 1 36725
0 36727 7 1 2 61086 36726
0 36728 5 1 1 36727
0 36729 7 1 2 33345 36728
0 36730 5 1 1 36729
0 36731 7 1 2 67338 36730
0 36732 5 1 1 36731
0 36733 7 1 2 83379 92107
0 36734 5 1 1 36733
0 36735 7 1 2 36732 36734
0 36736 5 1 1 36735
0 36737 7 1 2 59916 36736
0 36738 5 1 1 36737
0 36739 7 14 2 61087 68416
0 36740 5 2 1 95467
0 36741 7 2 2 78260 95468
0 36742 7 2 2 84048 95483
0 36743 5 1 1 95485
0 36744 7 1 2 60559 80117
0 36745 5 1 1 36744
0 36746 7 1 2 36743 36745
0 36747 5 1 1 36746
0 36748 7 1 2 70617 36747
0 36749 5 1 1 36748
0 36750 7 1 2 77641 94873
0 36751 5 1 1 36750
0 36752 7 1 2 36749 36751
0 36753 5 1 1 36752
0 36754 7 1 2 72127 36753
0 36755 5 1 1 36754
0 36756 7 1 2 74071 82491
0 36757 5 1 1 36756
0 36758 7 1 2 77790 36757
0 36759 5 1 1 36758
0 36760 7 1 2 80667 77642
0 36761 5 1 1 36760
0 36762 7 1 2 36759 36761
0 36763 5 1 1 36762
0 36764 7 1 2 60560 36763
0 36765 5 1 1 36764
0 36766 7 1 2 36755 36765
0 36767 7 1 2 36738 36766
0 36768 5 1 1 36767
0 36769 7 1 2 66724 36768
0 36770 5 1 1 36769
0 36771 7 5 2 78712 93635
0 36772 5 1 1 95487
0 36773 7 1 2 82886 95488
0 36774 7 1 2 70913 36773
0 36775 5 1 1 36774
0 36776 7 1 2 36770 36775
0 36777 5 1 1 36776
0 36778 7 1 2 59349 36777
0 36779 5 1 1 36778
0 36780 7 1 2 75455 95489
0 36781 5 1 1 36780
0 36782 7 1 2 69310 93297
0 36783 5 1 1 36782
0 36784 7 1 2 74910 36783
0 36785 5 1 1 36784
0 36786 7 1 2 59917 36785
0 36787 5 1 1 36786
0 36788 7 1 2 3821 84814
0 36789 5 1 1 36788
0 36790 7 1 2 73916 36789
0 36791 5 1 1 36790
0 36792 7 1 2 36787 36791
0 36793 5 1 1 36792
0 36794 7 1 2 63519 36793
0 36795 5 1 1 36794
0 36796 7 1 2 65018 76327
0 36797 5 1 1 36796
0 36798 7 1 2 77791 36797
0 36799 5 1 1 36798
0 36800 7 4 2 83758 83118
0 36801 7 1 2 76149 3106
0 36802 7 1 2 95492 36801
0 36803 5 1 1 36802
0 36804 7 1 2 36799 36803
0 36805 7 1 2 36795 36804
0 36806 5 1 1 36805
0 36807 7 1 2 60561 36806
0 36808 5 1 1 36807
0 36809 7 1 2 93038 93466
0 36810 5 1 1 36809
0 36811 7 1 2 90512 94627
0 36812 7 1 2 95374 36811
0 36813 5 1 1 36812
0 36814 7 1 2 36810 36813
0 36815 5 1 1 36814
0 36816 7 1 2 68417 36815
0 36817 5 1 1 36816
0 36818 7 1 2 90934 93298
0 36819 5 1 1 36818
0 36820 7 1 2 4073 36819
0 36821 5 1 1 36820
0 36822 7 1 2 90607 36821
0 36823 5 1 1 36822
0 36824 7 1 2 36817 36823
0 36825 5 1 1 36824
0 36826 7 1 2 59564 36825
0 36827 5 1 1 36826
0 36828 7 1 2 80637 80704
0 36829 7 1 2 95486 36828
0 36830 5 1 1 36829
0 36831 7 1 2 36827 36830
0 36832 7 1 2 36808 36831
0 36833 5 1 1 36832
0 36834 7 1 2 66725 36833
0 36835 5 1 1 36834
0 36836 7 1 2 36781 36835
0 36837 7 1 2 36779 36836
0 36838 5 1 1 36837
0 36839 7 1 2 75324 36838
0 36840 5 1 1 36839
0 36841 7 3 2 61359 83595
0 36842 5 2 1 95496
0 36843 7 1 2 89341 95497
0 36844 5 2 1 36843
0 36845 7 2 2 85462 88742
0 36846 5 3 1 95503
0 36847 7 1 2 95501 95504
0 36848 5 1 1 36847
0 36849 7 1 2 76519 36848
0 36850 5 1 1 36849
0 36851 7 1 2 70192 84019
0 36852 7 1 2 95505 36851
0 36853 5 1 1 36852
0 36854 7 1 2 36850 36853
0 36855 5 1 1 36854
0 36856 7 1 2 67339 36855
0 36857 5 1 1 36856
0 36858 7 1 2 70246 95506
0 36859 5 1 1 36858
0 36860 7 1 2 36857 36859
0 36861 5 1 1 36860
0 36862 7 1 2 67677 36861
0 36863 5 1 1 36862
0 36864 7 1 2 70618 95507
0 36865 5 1 1 36864
0 36866 7 1 2 72519 91618
0 36867 7 2 2 89295 36866
0 36868 5 1 1 95508
0 36869 7 1 2 61575 95509
0 36870 5 1 1 36869
0 36871 7 1 2 91848 36870
0 36872 5 1 1 36871
0 36873 7 1 2 36865 36872
0 36874 7 1 2 36863 36873
0 36875 5 1 1 36874
0 36876 7 1 2 68042 36875
0 36877 5 1 1 36876
0 36878 7 4 2 60373 89338
0 36879 5 1 1 95510
0 36880 7 1 2 63095 95511
0 36881 5 1 1 36880
0 36882 7 1 2 71629 73462
0 36883 5 2 1 36882
0 36884 7 1 2 70232 95514
0 36885 5 1 1 36884
0 36886 7 1 2 70619 82313
0 36887 5 1 1 36886
0 36888 7 1 2 36885 36887
0 36889 5 1 1 36888
0 36890 7 1 2 60931 36889
0 36891 5 1 1 36890
0 36892 7 1 2 66058 92914
0 36893 5 1 1 36892
0 36894 7 1 2 70620 36893
0 36895 5 1 1 36894
0 36896 7 1 2 36891 36895
0 36897 5 1 1 36896
0 36898 7 1 2 63096 36897
0 36899 5 1 1 36898
0 36900 7 2 2 81940 93062
0 36901 5 1 1 95516
0 36902 7 1 2 68043 73509
0 36903 7 1 2 36901 36902
0 36904 5 1 1 36903
0 36905 7 1 2 36899 36904
0 36906 5 1 1 36905
0 36907 7 1 2 67678 36906
0 36908 5 1 1 36907
0 36909 7 1 2 70066 91534
0 36910 5 2 1 36909
0 36911 7 2 2 77433 95518
0 36912 7 1 2 61088 95520
0 36913 5 1 1 36912
0 36914 7 1 2 77378 91956
0 36915 5 1 1 36914
0 36916 7 1 2 36913 36915
0 36917 5 1 1 36916
0 36918 7 1 2 76045 36917
0 36919 5 1 1 36918
0 36920 7 1 2 73300 92504
0 36921 5 1 1 36920
0 36922 7 1 2 36919 36921
0 36923 5 1 1 36922
0 36924 7 1 2 59350 36923
0 36925 5 1 1 36924
0 36926 7 1 2 82245 78434
0 36927 5 1 1 36926
0 36928 7 1 2 8579 36927
0 36929 5 1 1 36928
0 36930 7 1 2 70233 36929
0 36931 5 1 1 36930
0 36932 7 1 2 77379 75015
0 36933 7 1 2 89255 36932
0 36934 5 1 1 36933
0 36935 7 1 2 36931 36934
0 36936 5 1 1 36935
0 36937 7 1 2 60932 36936
0 36938 5 1 1 36937
0 36939 7 1 2 36925 36938
0 36940 7 1 2 36908 36939
0 36941 5 1 1 36940
0 36942 7 1 2 91673 36941
0 36943 5 1 1 36942
0 36944 7 1 2 36881 36943
0 36945 7 1 2 36877 36944
0 36946 5 1 1 36945
0 36947 7 1 2 68418 36946
0 36948 5 1 1 36947
0 36949 7 1 2 64786 72842
0 36950 5 1 1 36949
0 36951 7 1 2 67340 36950
0 36952 5 1 1 36951
0 36953 7 1 2 76721 83335
0 36954 5 1 1 36953
0 36955 7 1 2 83351 86548
0 36956 7 1 2 36954 36955
0 36957 7 1 2 36952 36956
0 36958 5 1 1 36957
0 36959 7 1 2 75501 90608
0 36960 7 1 2 36958 36959
0 36961 5 1 1 36960
0 36962 7 1 2 36948 36961
0 36963 5 1 1 36962
0 36964 7 1 2 66726 36963
0 36965 5 1 1 36964
0 36966 7 2 2 74072 76010
0 36967 5 2 1 95522
0 36968 7 2 2 69572 95524
0 36969 5 1 1 95526
0 36970 7 2 2 80227 95527
0 36971 5 1 1 95528
0 36972 7 1 2 75325 95529
0 36973 5 1 1 36972
0 36974 7 1 2 93354 36973
0 36975 5 1 1 36974
0 36976 7 1 2 90609 36975
0 36977 5 1 1 36976
0 36978 7 2 2 79901 69409
0 36979 7 1 2 74437 95530
0 36980 7 1 2 90165 36979
0 36981 5 2 1 36980
0 36982 7 1 2 83911 76070
0 36983 5 1 1 36982
0 36984 7 1 2 95532 36983
0 36985 5 1 1 36984
0 36986 7 2 2 68419 90636
0 36987 7 1 2 36985 95534
0 36988 5 1 1 36987
0 36989 7 1 2 36977 36988
0 36990 5 1 1 36989
0 36991 7 1 2 66727 36990
0 36992 5 1 1 36991
0 36993 7 3 2 69189 79441
0 36994 7 4 2 60562 67087
0 36995 5 1 1 95539
0 36996 7 1 2 78261 36995
0 36997 7 1 2 95536 36996
0 36998 7 1 2 71334 36997
0 36999 5 1 1 36998
0 37000 7 1 2 36772 36999
0 37001 5 1 1 37000
0 37002 7 1 2 59565 37001
0 37003 5 1 1 37002
0 37004 7 1 2 76722 87429
0 37005 5 1 1 37004
0 37006 7 1 2 21800 37005
0 37007 5 1 1 37006
0 37008 7 1 2 90610 37007
0 37009 5 1 1 37008
0 37010 7 1 2 37003 37009
0 37011 5 1 1 37010
0 37012 7 1 2 61576 37011
0 37013 5 1 1 37012
0 37014 7 1 2 80362 77792
0 37015 7 1 2 76071 37014
0 37016 5 1 1 37015
0 37017 7 1 2 37013 37016
0 37018 5 1 1 37017
0 37019 7 1 2 76786 37018
0 37020 5 1 1 37019
0 37021 7 1 2 81794 86902
0 37022 7 1 2 95490 37021
0 37023 5 1 1 37022
0 37024 7 1 2 37020 37023
0 37025 7 1 2 36992 37024
0 37026 5 1 1 37025
0 37027 7 1 2 71226 37026
0 37028 5 1 1 37027
0 37029 7 1 2 59351 82887
0 37030 5 1 1 37029
0 37031 7 1 2 72355 37030
0 37032 5 1 1 37031
0 37033 7 2 2 83104 37032
0 37034 7 2 2 91058 95543
0 37035 5 1 1 95545
0 37036 7 1 2 90124 95546
0 37037 5 1 1 37036
0 37038 7 1 2 86770 37037
0 37039 7 1 2 37028 37038
0 37040 7 1 2 36965 37039
0 37041 7 1 2 36840 37040
0 37042 5 1 1 37041
0 37043 7 1 2 68981 37042
0 37044 7 1 2 36707 37043
0 37045 5 1 1 37044
0 37046 7 1 2 67679 95515
0 37047 5 1 1 37046
0 37048 7 1 2 59566 93031
0 37049 5 1 1 37048
0 37050 7 1 2 37047 37049
0 37051 5 1 1 37050
0 37052 7 1 2 77659 37051
0 37053 5 1 1 37052
0 37054 7 1 2 61360 77643
0 37055 5 1 1 37054
0 37056 7 1 2 73677 93315
0 37057 5 1 1 37056
0 37058 7 1 2 59567 37057
0 37059 5 1 1 37058
0 37060 7 1 2 37055 37059
0 37061 5 1 1 37060
0 37062 7 1 2 59352 37061
0 37063 5 1 1 37062
0 37064 7 1 2 61361 95372
0 37065 5 2 1 37064
0 37066 7 1 2 76433 95547
0 37067 5 1 1 37066
0 37068 7 1 2 69371 77691
0 37069 5 1 1 37068
0 37070 7 1 2 37067 37069
0 37071 5 1 1 37070
0 37072 7 2 2 71374 73293
0 37073 5 1 1 95549
0 37074 7 1 2 37071 95550
0 37075 5 1 1 37074
0 37076 7 1 2 91307 37075
0 37077 5 1 1 37076
0 37078 7 1 2 37063 37077
0 37079 5 1 1 37078
0 37080 7 1 2 60163 37079
0 37081 5 1 1 37080
0 37082 7 1 2 37053 37081
0 37083 5 1 1 37082
0 37084 7 1 2 60933 37083
0 37085 5 1 1 37084
0 37086 7 1 2 76917 71928
0 37087 5 1 1 37086
0 37088 7 1 2 71227 37087
0 37089 5 1 1 37088
0 37090 7 1 2 73192 83336
0 37091 5 1 1 37090
0 37092 7 1 2 77125 83352
0 37093 5 1 1 37092
0 37094 7 1 2 73236 37093
0 37095 5 1 1 37094
0 37096 7 1 2 37091 37095
0 37097 7 1 2 37089 37096
0 37098 5 1 1 37097
0 37099 7 1 2 70621 37098
0 37100 5 1 1 37099
0 37101 7 1 2 37085 37100
0 37102 5 1 1 37101
0 37103 7 1 2 61577 37102
0 37104 5 1 1 37103
0 37105 7 3 2 83883 73243
0 37106 5 2 1 95551
0 37107 7 2 2 67341 95554
0 37108 7 1 2 67680 78675
0 37109 5 1 1 37108
0 37110 7 1 2 229 37109
0 37111 5 1 1 37110
0 37112 7 1 2 95556 37111
0 37113 5 1 1 37112
0 37114 7 1 2 72234 92605
0 37115 5 1 1 37114
0 37116 7 2 2 37113 37115
0 37117 5 2 1 95558
0 37118 7 1 2 69934 91594
0 37119 5 2 1 37118
0 37120 7 1 2 71434 95562
0 37121 5 1 1 37120
0 37122 7 1 2 67342 37121
0 37123 5 1 1 37122
0 37124 7 1 2 70822 92209
0 37125 7 1 2 93119 37124
0 37126 7 1 2 37123 37125
0 37127 5 1 1 37126
0 37128 7 1 2 74653 37127
0 37129 5 1 1 37128
0 37130 7 1 2 95559 37129
0 37131 5 1 1 37130
0 37132 7 1 2 68044 74323
0 37133 7 1 2 37131 37132
0 37134 5 1 1 37133
0 37135 7 1 2 37104 37134
0 37136 5 1 1 37135
0 37137 7 1 2 60374 37136
0 37138 5 1 1 37137
0 37139 7 1 2 61578 87760
0 37140 7 1 2 95560 37139
0 37141 5 1 1 37140
0 37142 7 1 2 37138 37141
0 37143 5 1 1 37142
0 37144 7 1 2 87902 37143
0 37145 5 1 1 37144
0 37146 7 1 2 80615 91564
0 37147 5 1 1 37146
0 37148 7 1 2 67088 72520
0 37149 5 2 1 37148
0 37150 7 1 2 37147 95564
0 37151 5 1 1 37150
0 37152 7 1 2 61089 37151
0 37153 5 1 1 37152
0 37154 7 1 2 82252 37153
0 37155 5 1 1 37154
0 37156 7 1 2 77085 37155
0 37157 5 1 1 37156
0 37158 7 1 2 75933 37157
0 37159 5 1 1 37158
0 37160 7 1 2 90997 91200
0 37161 5 1 1 37160
0 37162 7 1 2 69694 37161
0 37163 5 1 1 37162
0 37164 7 1 2 76720 94699
0 37165 5 1 1 37164
0 37166 7 1 2 29911 37165
0 37167 7 1 2 37163 37166
0 37168 5 1 1 37167
0 37169 7 1 2 62142 37168
0 37170 5 1 1 37169
0 37171 7 1 2 67681 2454
0 37172 5 3 1 37171
0 37173 7 1 2 64558 95566
0 37174 5 1 1 37173
0 37175 7 1 2 91201 37174
0 37176 5 1 1 37175
0 37177 7 1 2 72560 37176
0 37178 5 1 1 37177
0 37179 7 1 2 79420 37178
0 37180 7 1 2 37170 37179
0 37181 7 1 2 37159 37180
0 37182 5 1 1 37181
0 37183 7 1 2 71574 37182
0 37184 5 1 1 37183
0 37185 7 1 2 69265 73797
0 37186 5 2 1 37185
0 37187 7 1 2 59568 95569
0 37188 5 1 1 37187
0 37189 7 2 2 91207 37188
0 37190 5 1 1 95571
0 37191 7 1 2 64787 95572
0 37192 5 1 1 37191
0 37193 7 1 2 72013 90248
0 37194 5 1 1 37193
0 37195 7 1 2 37192 37194
0 37196 5 2 1 37195
0 37197 7 1 2 88353 95573
0 37198 5 1 1 37197
0 37199 7 1 2 70823 85663
0 37200 5 1 1 37199
0 37201 7 1 2 37198 37200
0 37202 7 1 2 37184 37201
0 37203 5 1 1 37202
0 37204 7 1 2 63097 37203
0 37205 5 1 1 37204
0 37206 7 1 2 83684 94076
0 37207 5 1 1 37206
0 37208 7 1 2 66334 37207
0 37209 5 1 1 37208
0 37210 7 1 2 63098 74415
0 37211 5 1 1 37210
0 37212 7 2 2 61362 72799
0 37213 5 1 1 95575
0 37214 7 1 2 62715 37213
0 37215 5 1 1 37214
0 37216 7 1 2 37211 37215
0 37217 7 1 2 37209 37216
0 37218 5 1 1 37217
0 37219 7 1 2 62363 37218
0 37220 5 1 1 37219
0 37221 7 1 2 68045 90232
0 37222 5 1 1 37221
0 37223 7 1 2 29564 37222
0 37224 5 1 1 37223
0 37225 7 1 2 37220 37224
0 37226 5 1 1 37225
0 37227 7 1 2 72356 37226
0 37228 5 1 1 37227
0 37229 7 2 2 64317 82791
0 37230 5 1 1 95577
0 37231 7 1 2 68046 81637
0 37232 5 2 1 37231
0 37233 7 1 2 95578 95579
0 37234 5 1 1 37233
0 37235 7 1 2 73180 31480
0 37236 7 1 2 37234 37235
0 37237 5 1 1 37236
0 37238 7 1 2 72357 37237
0 37239 5 1 1 37238
0 37240 7 2 2 67343 76261
0 37241 5 2 1 95581
0 37242 7 1 2 88709 95583
0 37243 5 1 1 37242
0 37244 7 1 2 68047 37243
0 37245 5 1 1 37244
0 37246 7 1 2 77692 37245
0 37247 5 1 1 37246
0 37248 7 1 2 74785 77693
0 37249 5 1 1 37248
0 37250 7 1 2 94867 37249
0 37251 5 1 1 37250
0 37252 7 1 2 77095 37251
0 37253 5 1 1 37252
0 37254 7 1 2 37247 37253
0 37255 7 1 2 37239 37254
0 37256 5 1 1 37255
0 37257 7 1 2 65890 37256
0 37258 5 1 1 37257
0 37259 7 1 2 78082 86914
0 37260 5 1 1 37259
0 37261 7 1 2 71228 15721
0 37262 7 1 2 78454 37261
0 37263 5 1 1 37262
0 37264 7 1 2 87811 37263
0 37265 5 1 1 37264
0 37266 7 1 2 37260 37265
0 37267 7 1 2 91336 89276
0 37268 5 1 1 37267
0 37269 7 1 2 88029 37268
0 37270 5 1 1 37269
0 37271 7 1 2 71650 84802
0 37272 7 1 2 93157 37271
0 37273 5 1 1 37272
0 37274 7 1 2 65266 37273
0 37275 5 1 1 37274
0 37276 7 1 2 37270 37275
0 37277 7 1 2 37266 37276
0 37278 7 1 2 37258 37277
0 37279 7 1 2 62143 91199
0 37280 5 1 1 37279
0 37281 7 1 2 80449 37280
0 37282 5 1 1 37281
0 37283 7 1 2 77218 37282
0 37284 5 1 1 37283
0 37285 7 2 2 74818 74546
0 37286 5 1 1 95585
0 37287 7 1 2 63099 37286
0 37288 5 1 1 37287
0 37289 7 1 2 72521 88646
0 37290 5 2 1 37289
0 37291 7 1 2 66335 95587
0 37292 5 1 1 37291
0 37293 7 2 2 76398 72616
0 37294 5 1 1 95589
0 37295 7 1 2 37292 37294
0 37296 7 1 2 37288 37295
0 37297 7 1 2 37284 37296
0 37298 7 1 2 67682 91378
0 37299 5 2 1 37298
0 37300 7 1 2 72358 95591
0 37301 5 1 1 37300
0 37302 7 1 2 72014 69455
0 37303 5 1 1 37302
0 37304 7 1 2 37301 37303
0 37305 5 1 1 37304
0 37306 7 1 2 77648 37305
0 37307 5 1 1 37306
0 37308 7 1 2 88425 30555
0 37309 5 1 1 37308
0 37310 7 2 2 71823 90501
0 37311 7 1 2 37309 95593
0 37312 5 1 1 37311
0 37313 7 1 2 37307 37312
0 37314 7 1 2 37297 37313
0 37315 5 1 1 37314
0 37316 7 1 2 65019 37315
0 37317 5 1 1 37316
0 37318 7 1 2 62144 90520
0 37319 5 1 1 37318
0 37320 7 1 2 77501 37319
0 37321 5 1 1 37320
0 37322 7 1 2 74030 37321
0 37323 5 1 1 37322
0 37324 7 4 2 63100 72359
0 37325 5 4 1 95595
0 37326 7 1 2 87784 95596
0 37327 5 1 1 37326
0 37328 7 1 2 77719 37327
0 37329 7 1 2 37323 37328
0 37330 5 1 1 37329
0 37331 7 1 2 72561 37330
0 37332 5 1 1 37331
0 37333 7 1 2 37317 37332
0 37334 7 1 2 37278 37333
0 37335 7 1 2 37228 37334
0 37336 5 1 1 37335
0 37337 7 1 2 66559 37336
0 37338 5 1 1 37337
0 37339 7 1 2 61579 2770
0 37340 5 1 1 37339
0 37341 7 1 2 70824 88933
0 37342 7 1 2 37340 37341
0 37343 5 1 1 37342
0 37344 7 1 2 91300 37343
0 37345 5 1 1 37344
0 37346 7 1 2 81656 37345
0 37347 5 1 1 37346
0 37348 7 1 2 68420 37347
0 37349 7 1 2 37338 37348
0 37350 7 1 2 37205 37349
0 37351 5 1 1 37350
0 37352 7 1 2 70622 74534
0 37353 7 1 2 95422 37352
0 37354 5 1 1 37353
0 37355 7 1 2 61580 37354
0 37356 5 1 1 37355
0 37357 7 1 2 72880 72360
0 37358 5 1 1 37357
0 37359 7 1 2 76645 37358
0 37360 5 1 1 37359
0 37361 7 1 2 67683 95436
0 37362 5 2 1 37361
0 37363 7 1 2 63101 95603
0 37364 7 1 2 37360 37363
0 37365 7 1 2 37356 37364
0 37366 5 1 1 37365
0 37367 7 1 2 59353 76099
0 37368 5 1 1 37367
0 37369 7 1 2 95592 37368
0 37370 5 1 1 37369
0 37371 7 1 2 80435 37370
0 37372 5 1 1 37371
0 37373 7 1 2 71120 37372
0 37374 5 1 1 37373
0 37375 7 1 2 62716 94901
0 37376 5 1 1 37375
0 37377 7 1 2 37374 37376
0 37378 5 1 1 37377
0 37379 7 1 2 62364 37378
0 37380 5 1 1 37379
0 37381 7 1 2 72495 95466
0 37382 5 1 1 37381
0 37383 7 1 2 79975 71121
0 37384 5 1 1 37383
0 37385 7 2 2 69856 86516
0 37386 5 1 1 95605
0 37387 7 1 2 37384 37386
0 37388 5 1 1 37387
0 37389 7 1 2 62717 37388
0 37390 5 1 1 37389
0 37391 7 1 2 68048 77750
0 37392 7 1 2 37390 37391
0 37393 7 1 2 37382 37392
0 37394 7 1 2 37380 37393
0 37395 5 1 1 37394
0 37396 7 1 2 37366 37395
0 37397 5 1 1 37396
0 37398 7 1 2 3264 35069
0 37399 5 1 1 37398
0 37400 7 1 2 63102 37399
0 37401 5 1 1 37400
0 37402 7 1 2 95464 37401
0 37403 5 1 1 37402
0 37404 7 1 2 62365 37403
0 37405 5 1 1 37404
0 37406 7 1 2 95429 37405
0 37407 5 1 1 37406
0 37408 7 1 2 78664 37407
0 37409 5 1 1 37408
0 37410 7 1 2 75931 83337
0 37411 5 1 1 37410
0 37412 7 1 2 1606 87579
0 37413 7 1 2 37411 37412
0 37414 5 1 1 37413
0 37415 7 1 2 75613 37414
0 37416 5 1 1 37415
0 37417 7 1 2 72800 87430
0 37418 5 1 1 37417
0 37419 7 1 2 93473 37418
0 37420 5 1 1 37419
0 37421 7 1 2 71229 37420
0 37422 5 1 1 37421
0 37423 7 1 2 63103 82545
0 37424 5 1 1 37423
0 37425 7 1 2 83310 37424
0 37426 5 1 1 37425
0 37427 7 1 2 72857 37426
0 37428 5 1 1 37427
0 37429 7 1 2 83912 88414
0 37430 5 1 1 37429
0 37431 7 1 2 63520 37430
0 37432 7 1 2 37428 37431
0 37433 7 1 2 37422 37432
0 37434 7 1 2 37416 37433
0 37435 7 1 2 37409 37434
0 37436 7 1 2 37397 37435
0 37437 7 1 2 95462 37436
0 37438 5 1 1 37437
0 37439 7 1 2 87177 37438
0 37440 7 1 2 37351 37439
0 37441 5 1 1 37440
0 37442 7 1 2 37145 37441
0 37443 5 1 1 37442
0 37444 7 1 2 68982 37443
0 37445 5 1 1 37444
0 37446 7 1 2 64788 93318
0 37447 5 1 1 37446
0 37448 7 2 2 70193 88108
0 37449 7 1 2 37447 95607
0 37450 5 1 1 37449
0 37451 7 1 2 69695 93121
0 37452 5 1 1 37451
0 37453 7 2 2 61363 37452
0 37454 7 1 2 83390 95609
0 37455 5 1 1 37454
0 37456 7 1 2 70194 87978
0 37457 5 1 1 37456
0 37458 7 1 2 71313 73878
0 37459 5 1 1 37458
0 37460 7 1 2 61364 37459
0 37461 5 1 1 37460
0 37462 7 1 2 77209 84119
0 37463 5 1 1 37462
0 37464 7 1 2 91611 37463
0 37465 7 1 2 37461 37464
0 37466 7 1 2 37457 37465
0 37467 5 1 1 37466
0 37468 7 1 2 61581 37467
0 37469 5 1 1 37468
0 37470 7 1 2 37455 37469
0 37471 5 1 1 37470
0 37472 7 1 2 67684 37471
0 37473 5 1 1 37472
0 37474 7 1 2 37450 37473
0 37475 5 1 1 37474
0 37476 7 1 2 61090 37475
0 37477 5 1 1 37476
0 37478 7 1 2 78226 82085
0 37479 5 1 1 37478
0 37480 7 1 2 69935 37479
0 37481 5 1 1 37480
0 37482 7 1 2 4376 74123
0 37483 5 1 1 37482
0 37484 7 1 2 59918 37483
0 37485 5 1 1 37484
0 37486 7 1 2 37481 37485
0 37487 5 1 1 37486
0 37488 7 1 2 95608 37487
0 37489 5 1 1 37488
0 37490 7 1 2 37477 37489
0 37491 5 1 1 37490
0 37492 7 1 2 68049 37491
0 37493 5 1 1 37492
0 37494 7 1 2 71499 93160
0 37495 5 1 1 37494
0 37496 7 1 2 76918 73427
0 37497 5 1 1 37496
0 37498 7 1 2 61365 92487
0 37499 7 1 2 37497 37498
0 37500 5 1 1 37499
0 37501 7 1 2 37495 37500
0 37502 5 1 1 37501
0 37503 7 1 2 67685 37502
0 37504 5 1 1 37503
0 37505 7 1 2 75715 73418
0 37506 5 2 1 37505
0 37507 7 1 2 37504 95611
0 37508 5 1 1 37507
0 37509 7 1 2 61091 37508
0 37510 5 1 1 37509
0 37511 7 2 2 70623 91526
0 37512 7 1 2 69936 95613
0 37513 5 1 1 37512
0 37514 7 1 2 37510 37513
0 37515 5 1 1 37514
0 37516 7 1 2 61582 37515
0 37517 5 1 1 37516
0 37518 7 1 2 37493 37517
0 37519 5 1 1 37518
0 37520 7 1 2 60375 37519
0 37521 5 1 1 37520
0 37522 7 2 2 76046 92488
0 37523 5 1 1 95615
0 37524 7 1 2 67686 95616
0 37525 5 1 1 37524
0 37526 7 2 2 68050 72128
0 37527 5 1 1 95617
0 37528 7 1 2 59919 95618
0 37529 5 1 1 37528
0 37530 7 1 2 37525 37529
0 37531 5 1 1 37530
0 37532 7 1 2 59354 37531
0 37533 5 1 1 37532
0 37534 7 3 2 60808 68051
0 37535 7 1 2 73579 74667
0 37536 5 1 1 37535
0 37537 7 1 2 95619 37536
0 37538 5 1 1 37537
0 37539 7 1 2 37533 37538
0 37540 5 1 1 37539
0 37541 7 1 2 61092 37540
0 37542 5 1 1 37541
0 37543 7 1 2 23439 93316
0 37544 5 1 1 37543
0 37545 7 1 2 72129 37544
0 37546 5 1 1 37545
0 37547 7 1 2 22298 37546
0 37548 5 1 1 37547
0 37549 7 1 2 68052 37548
0 37550 5 1 1 37549
0 37551 7 1 2 37542 37550
0 37552 5 1 1 37551
0 37553 7 1 2 61366 37552
0 37554 5 1 1 37553
0 37555 7 1 2 82492 72147
0 37556 5 3 1 37555
0 37557 7 1 2 72130 95622
0 37558 5 1 1 37557
0 37559 7 1 2 93144 37558
0 37560 5 1 1 37559
0 37561 7 1 2 59920 37560
0 37562 5 1 1 37561
0 37563 7 1 2 73286 71880
0 37564 5 1 1 37563
0 37565 7 1 2 37562 37564
0 37566 5 1 1 37565
0 37567 7 1 2 82461 37566
0 37568 5 1 1 37567
0 37569 7 1 2 37554 37568
0 37570 5 1 1 37569
0 37571 7 1 2 75326 37570
0 37572 5 1 1 37571
0 37573 7 1 2 71881 89511
0 37574 5 1 1 37573
0 37575 7 1 2 78237 91958
0 37576 5 1 1 37575
0 37577 7 1 2 75327 37576
0 37578 5 1 1 37577
0 37579 7 2 2 76315 91511
0 37580 5 1 1 95625
0 37581 7 1 2 37578 37580
0 37582 5 1 1 37581
0 37583 7 1 2 59921 37582
0 37584 5 1 1 37583
0 37585 7 1 2 37574 37584
0 37586 5 1 1 37585
0 37587 7 1 2 59569 37586
0 37588 5 1 1 37587
0 37589 7 1 2 82268 84064
0 37590 5 2 1 37589
0 37591 7 1 2 74911 95627
0 37592 5 1 1 37591
0 37593 7 1 2 75328 37592
0 37594 5 1 1 37593
0 37595 7 1 2 89609 37594
0 37596 7 1 2 37588 37595
0 37597 5 1 1 37596
0 37598 7 1 2 82992 37597
0 37599 5 1 1 37598
0 37600 7 1 2 75614 73928
0 37601 5 1 1 37600
0 37602 7 1 2 92489 89613
0 37603 7 1 2 37601 37602
0 37604 5 1 1 37603
0 37605 7 1 2 37599 37604
0 37606 5 1 1 37605
0 37607 7 1 2 69410 37606
0 37608 5 1 1 37607
0 37609 7 1 2 37523 37527
0 37610 5 1 1 37609
0 37611 7 1 2 59355 37610
0 37612 5 1 1 37611
0 37613 7 1 2 78462 95620
0 37614 5 1 1 37613
0 37615 7 1 2 90094 37614
0 37616 7 1 2 37612 37615
0 37617 5 1 1 37616
0 37618 7 1 2 75502 37617
0 37619 5 1 1 37618
0 37620 7 1 2 73435 83431
0 37621 7 1 2 95376 37620
0 37622 5 1 1 37621
0 37623 7 1 2 37619 37622
0 37624 7 1 2 37608 37623
0 37625 7 1 2 37572 37624
0 37626 5 1 1 37625
0 37627 7 1 2 68421 37626
0 37628 5 1 1 37627
0 37629 7 1 2 78376 88879
0 37630 5 1 1 37629
0 37631 7 1 2 92244 37630
0 37632 5 1 1 37631
0 37633 7 1 2 70624 37632
0 37634 5 1 1 37633
0 37635 7 1 2 75453 91072
0 37636 5 1 1 37635
0 37637 7 1 2 37634 37636
0 37638 5 1 1 37637
0 37639 7 1 2 67089 37638
0 37640 5 1 1 37639
0 37641 7 2 2 61093 88109
0 37642 7 1 2 83029 95629
0 37643 5 1 1 37642
0 37644 7 1 2 37640 37643
0 37645 5 1 1 37644
0 37646 7 1 2 60376 37645
0 37647 5 1 1 37646
0 37648 7 1 2 75730 91073
0 37649 5 1 1 37648
0 37650 7 1 2 37647 37649
0 37651 5 1 1 37650
0 37652 7 1 2 74186 37651
0 37653 5 1 1 37652
0 37654 7 1 2 83426 76047
0 37655 5 1 1 37654
0 37656 7 1 2 82465 37655
0 37657 5 1 1 37656
0 37658 7 1 2 76901 82206
0 37659 5 1 1 37658
0 37660 7 1 2 37657 37659
0 37661 5 1 1 37660
0 37662 7 1 2 68422 82780
0 37663 5 1 1 37662
0 37664 7 1 2 37661 37663
0 37665 5 1 1 37664
0 37666 7 1 2 75503 37665
0 37667 5 1 1 37666
0 37668 7 1 2 76048 90810
0 37669 5 1 1 37668
0 37670 7 1 2 68053 73287
0 37671 5 1 1 37670
0 37672 7 1 2 65020 6026
0 37673 5 1 1 37672
0 37674 7 1 2 82781 37673
0 37675 5 1 1 37674
0 37676 7 1 2 37671 37675
0 37677 7 1 2 37669 37676
0 37678 5 1 1 37677
0 37679 7 1 2 75385 37678
0 37680 5 1 1 37679
0 37681 7 1 2 14879 37680
0 37682 5 1 1 37681
0 37683 7 1 2 91527 37682
0 37684 5 1 1 37683
0 37685 7 1 2 37667 37684
0 37686 5 1 1 37685
0 37687 7 1 2 76150 37686
0 37688 5 1 1 37687
0 37689 7 1 2 90838 94558
0 37690 7 1 2 95610 37689
0 37691 5 1 1 37690
0 37692 7 1 2 37688 37691
0 37693 7 1 2 37653 37692
0 37694 7 1 2 37628 37693
0 37695 7 1 2 37521 37694
0 37696 5 1 1 37695
0 37697 7 12 2 64111 86755
0 37698 7 1 2 37696 95631
0 37699 5 1 1 37698
0 37700 7 1 2 37445 37699
0 37701 5 1 1 37700
0 37702 7 1 2 60563 37701
0 37703 5 1 1 37702
0 37704 7 2 2 76787 78850
0 37705 5 4 1 95643
0 37706 7 1 2 88745 95645
0 37707 5 1 1 37706
0 37708 7 1 2 70263 94045
0 37709 5 1 1 37708
0 37710 7 1 2 88592 37709
0 37711 5 1 1 37710
0 37712 7 1 2 37707 37711
0 37713 5 1 1 37712
0 37714 7 1 2 94515 37713
0 37715 5 1 1 37714
0 37716 7 1 2 81348 95544
0 37717 5 1 1 37716
0 37718 7 1 2 94516 95356
0 37719 5 1 1 37718
0 37720 7 1 2 37717 37719
0 37721 5 1 1 37720
0 37722 7 1 2 62366 37721
0 37723 5 1 1 37722
0 37724 7 1 2 37715 37723
0 37725 5 1 1 37724
0 37726 7 1 2 62718 37725
0 37727 5 1 1 37726
0 37728 7 1 2 76748 80080
0 37729 5 1 1 37728
0 37730 7 1 2 78518 90534
0 37731 5 1 1 37730
0 37732 7 1 2 60377 37731
0 37733 5 1 1 37732
0 37734 7 1 2 70625 90451
0 37735 5 3 1 37734
0 37736 7 1 2 64318 95649
0 37737 7 1 2 37733 37736
0 37738 5 1 1 37737
0 37739 7 1 2 37729 37738
0 37740 5 1 1 37739
0 37741 7 1 2 64789 37740
0 37742 5 1 1 37741
0 37743 7 1 2 76749 93281
0 37744 5 1 1 37743
0 37745 7 1 2 37742 37744
0 37746 5 1 1 37745
0 37747 7 1 2 64559 37746
0 37748 5 1 1 37747
0 37749 7 1 2 72846 70902
0 37750 5 1 1 37749
0 37751 7 1 2 77751 37750
0 37752 5 1 1 37751
0 37753 7 1 2 65267 37752
0 37754 5 1 1 37753
0 37755 7 1 2 37748 37754
0 37756 5 1 1 37755
0 37757 7 1 2 62367 37756
0 37758 5 1 1 37757
0 37759 7 1 2 70067 88557
0 37760 5 1 1 37759
0 37761 7 2 2 72600 86490
0 37762 7 1 2 61094 93926
0 37763 5 1 1 37762
0 37764 7 2 2 95652 37763
0 37765 5 1 1 95654
0 37766 7 1 2 70825 95655
0 37767 5 1 1 37766
0 37768 7 2 2 37760 37767
0 37769 7 1 2 70264 94689
0 37770 5 1 1 37769
0 37771 7 1 2 86518 12850
0 37772 5 2 1 37771
0 37773 7 1 2 37770 95658
0 37774 5 1 1 37773
0 37775 7 1 2 95656 37774
0 37776 5 1 1 37775
0 37777 7 1 2 65268 37776
0 37778 5 1 1 37777
0 37779 7 1 2 65461 36868
0 37780 5 1 1 37779
0 37781 7 1 2 37778 37780
0 37782 7 1 2 37758 37781
0 37783 5 1 1 37782
0 37784 7 1 2 68054 37783
0 37785 5 1 1 37784
0 37786 7 5 2 59570 65462
0 37787 7 1 2 60809 95660
0 37788 7 1 2 93467 37787
0 37789 5 1 1 37788
0 37790 7 1 2 37785 37789
0 37791 5 1 1 37790
0 37792 7 1 2 85911 37791
0 37793 5 1 1 37792
0 37794 7 1 2 76072 92744
0 37795 5 1 1 37794
0 37796 7 1 2 37795 95533
0 37797 5 1 1 37796
0 37798 7 1 2 68423 37797
0 37799 5 1 1 37798
0 37800 7 1 2 67687 76788
0 37801 5 1 1 37800
0 37802 7 1 2 36971 37801
0 37803 5 1 1 37802
0 37804 7 1 2 79793 37803
0 37805 5 1 1 37804
0 37806 7 1 2 37799 37805
0 37807 5 1 1 37806
0 37808 7 1 2 65463 37807
0 37809 5 1 1 37808
0 37810 7 1 2 74324 87431
0 37811 5 1 1 37810
0 37812 7 1 2 80228 80798
0 37813 7 1 2 95525 37812
0 37814 5 1 1 37813
0 37815 7 1 2 37811 37814
0 37816 5 1 1 37815
0 37817 7 1 2 59356 37816
0 37818 5 1 1 37817
0 37819 7 1 2 78713 91030
0 37820 5 2 1 37819
0 37821 7 1 2 74742 95665
0 37822 5 1 1 37821
0 37823 7 1 2 74325 37822
0 37824 5 1 1 37823
0 37825 7 1 2 37818 37824
0 37826 5 1 1 37825
0 37827 7 1 2 60378 37826
0 37828 5 1 1 37827
0 37829 7 1 2 70626 86903
0 37830 7 1 2 94296 37829
0 37831 5 1 1 37830
0 37832 7 1 2 37828 37831
0 37833 5 1 1 37832
0 37834 7 1 2 63521 37833
0 37835 5 1 1 37834
0 37836 7 1 2 37809 37835
0 37837 5 1 1 37836
0 37838 7 1 2 71230 37837
0 37839 5 1 1 37838
0 37840 7 2 2 59357 77793
0 37841 5 2 1 95667
0 37842 7 1 2 79819 95669
0 37843 5 1 1 37842
0 37844 7 1 2 74600 37843
0 37845 5 1 1 37844
0 37846 7 1 2 77794 93106
0 37847 5 1 1 37846
0 37848 7 1 2 37845 37847
0 37849 5 1 1 37848
0 37850 7 1 2 67344 37849
0 37851 5 1 1 37850
0 37852 7 2 2 75113 73436
0 37853 5 1 1 95671
0 37854 7 1 2 89722 95672
0 37855 5 1 1 37854
0 37856 7 1 2 8034 37855
0 37857 7 1 2 37851 37856
0 37858 5 1 1 37857
0 37859 7 1 2 65464 37858
0 37860 5 1 1 37859
0 37861 7 1 2 80668 82414
0 37862 5 1 1 37861
0 37863 7 1 2 83703 77795
0 37864 5 1 1 37863
0 37865 7 1 2 37862 37864
0 37866 5 1 1 37865
0 37867 7 1 2 60379 37866
0 37868 5 1 1 37867
0 37869 7 1 2 37035 37868
0 37870 7 1 2 37860 37869
0 37871 5 1 1 37870
0 37872 7 1 2 76789 37871
0 37873 5 1 1 37872
0 37874 7 2 2 74152 84803
0 37875 5 1 1 95673
0 37876 7 1 2 60934 95674
0 37877 5 1 1 37876
0 37878 7 1 2 63104 92698
0 37879 5 1 1 37878
0 37880 7 1 2 37877 37879
0 37881 5 1 1 37880
0 37882 7 1 2 59571 37881
0 37883 5 1 1 37882
0 37884 7 1 2 83922 37875
0 37885 5 1 1 37884
0 37886 7 1 2 80074 37885
0 37887 5 1 1 37886
0 37888 7 1 2 37883 37887
0 37889 5 1 1 37888
0 37890 7 1 2 59358 37889
0 37891 5 1 1 37890
0 37892 7 1 2 79892 78435
0 37893 5 1 1 37892
0 37894 7 1 2 37891 37893
0 37895 5 1 1 37894
0 37896 7 1 2 82180 37895
0 37897 5 1 1 37896
0 37898 7 2 2 59922 91395
0 37899 7 1 2 89431 95675
0 37900 5 1 1 37899
0 37901 7 1 2 82701 95502
0 37902 5 2 1 37901
0 37903 7 1 2 92899 95677
0 37904 5 1 1 37903
0 37905 7 1 2 37900 37904
0 37906 5 1 1 37905
0 37907 7 1 2 76073 37906
0 37908 5 1 1 37907
0 37909 7 1 2 83704 95668
0 37910 5 1 1 37909
0 37911 7 1 2 74350 83408
0 37912 5 2 1 37911
0 37913 7 1 2 37910 95679
0 37914 5 1 1 37913
0 37915 7 1 2 74601 37914
0 37916 5 1 1 37915
0 37917 7 1 2 37908 37916
0 37918 7 1 2 37897 37917
0 37919 5 1 1 37918
0 37920 7 1 2 67345 37919
0 37921 5 1 1 37920
0 37922 7 1 2 65465 80955
0 37923 7 1 2 92745 37922
0 37924 7 1 2 95266 37923
0 37925 5 1 1 37924
0 37926 7 1 2 37921 37925
0 37927 7 1 2 37873 37926
0 37928 7 1 2 37839 37927
0 37929 7 1 2 37793 37928
0 37930 7 1 2 69696 88362
0 37931 5 1 1 37930
0 37932 7 1 2 74625 37931
0 37933 5 1 1 37932
0 37934 7 1 2 71575 37933
0 37935 5 1 1 37934
0 37936 7 1 2 70247 74547
0 37937 5 1 1 37936
0 37938 7 1 2 76750 37937
0 37939 5 1 1 37938
0 37940 7 1 2 37935 37939
0 37941 5 1 1 37940
0 37942 7 1 2 89889 37941
0 37943 5 1 1 37942
0 37944 7 2 2 65466 71604
0 37945 7 1 2 90778 95681
0 37946 5 1 1 37945
0 37947 7 1 2 37943 37946
0 37948 5 1 1 37947
0 37949 7 1 2 63105 37948
0 37950 5 1 1 37949
0 37951 7 1 2 84147 78873
0 37952 7 1 2 93309 37951
0 37953 5 1 1 37952
0 37954 7 1 2 37950 37953
0 37955 5 1 1 37954
0 37956 7 1 2 68424 37955
0 37957 5 1 1 37956
0 37958 7 1 2 82772 74753
0 37959 7 1 2 85761 37958
0 37960 5 1 1 37959
0 37961 7 1 2 89564 95181
0 37962 7 1 2 95531 37961
0 37963 5 1 1 37962
0 37964 7 1 2 37960 37963
0 37965 5 1 1 37964
0 37966 7 1 2 65467 37965
0 37967 5 1 1 37966
0 37968 7 1 2 63522 93454
0 37969 5 1 1 37968
0 37970 7 1 2 95680 37969
0 37971 5 1 1 37970
0 37972 7 1 2 86904 37971
0 37973 5 1 1 37972
0 37974 7 1 2 37967 37973
0 37975 7 1 2 37957 37974
0 37976 5 1 1 37975
0 37977 7 1 2 67688 37976
0 37978 5 1 1 37977
0 37979 7 1 2 82181 37073
0 37980 5 1 1 37979
0 37981 7 1 2 76646 92917
0 37982 5 1 1 37981
0 37983 7 1 2 37980 37982
0 37984 5 1 1 37983
0 37985 7 1 2 61095 37984
0 37986 5 1 1 37985
0 37987 7 2 2 59359 95661
0 37988 7 1 2 75114 81809
0 37989 7 1 2 95683 37988
0 37990 5 1 1 37989
0 37991 7 1 2 37986 37990
0 37992 5 1 1 37991
0 37993 7 1 2 60935 37992
0 37994 5 1 1 37993
0 37995 7 1 2 83262 91543
0 37996 7 1 2 89401 37995
0 37997 5 1 1 37996
0 37998 7 1 2 37994 37997
0 37999 5 1 1 37998
0 38000 7 1 2 59923 37999
0 38001 5 1 1 38000
0 38002 7 1 2 75329 82182
0 38003 5 1 1 38002
0 38004 7 1 2 38001 38003
0 38005 5 1 1 38004
0 38006 7 1 2 63106 38005
0 38007 5 1 1 38006
0 38008 7 1 2 78227 93018
0 38009 5 1 1 38008
0 38010 7 1 2 59360 38009
0 38011 5 1 1 38010
0 38012 7 2 2 62719 72159
0 38013 5 1 1 95685
0 38014 7 1 2 82654 38013
0 38015 5 1 1 38014
0 38016 7 1 2 38011 38015
0 38017 5 1 1 38016
0 38018 7 1 2 59924 38017
0 38019 5 1 1 38018
0 38020 7 1 2 63107 79987
0 38021 5 1 1 38020
0 38022 7 1 2 71882 38021
0 38023 5 1 1 38022
0 38024 7 2 2 38019 38023
0 38025 5 1 1 95687
0 38026 7 1 2 65269 95688
0 38027 5 1 1 38026
0 38028 7 1 2 79794 38027
0 38029 5 1 1 38028
0 38030 7 1 2 66059 456
0 38031 5 1 1 38030
0 38032 7 1 2 66560 38031
0 38033 5 1 1 38032
0 38034 7 1 2 95517 38033
0 38035 5 1 1 38034
0 38036 7 1 2 67689 38035
0 38037 5 1 1 38036
0 38038 7 1 2 59361 76106
0 38039 5 1 1 38038
0 38040 7 1 2 87567 38039
0 38041 5 1 1 38040
0 38042 7 1 2 76049 38041
0 38043 5 1 1 38042
0 38044 7 1 2 84058 38043
0 38045 7 1 2 38037 38044
0 38046 5 1 1 38045
0 38047 7 1 2 83745 38046
0 38048 5 1 1 38047
0 38049 7 1 2 38029 38048
0 38050 5 1 1 38049
0 38051 7 1 2 65468 38050
0 38052 5 1 1 38051
0 38053 7 1 2 90727 38025
0 38054 5 1 1 38053
0 38055 7 1 2 38052 38054
0 38056 7 1 2 38007 38055
0 38057 5 1 1 38056
0 38058 7 1 2 70195 38057
0 38059 5 1 1 38058
0 38060 7 1 2 37978 38059
0 38061 7 1 2 37929 38060
0 38062 7 1 2 37727 38061
0 38063 5 1 1 38062
0 38064 7 1 2 87178 38063
0 38065 5 1 1 38064
0 38066 7 1 2 69266 91354
0 38067 5 1 1 38066
0 38068 7 1 2 74412 93097
0 38069 5 2 1 38068
0 38070 7 1 2 87242 95689
0 38071 5 1 1 38070
0 38072 7 1 2 83484 82809
0 38073 7 1 2 88532 38072
0 38074 5 1 1 38073
0 38075 7 1 2 38071 38074
0 38076 7 1 2 38067 38075
0 38077 5 1 1 38076
0 38078 7 1 2 62720 38077
0 38079 5 1 1 38078
0 38080 7 1 2 75232 78649
0 38081 5 1 1 38080
0 38082 7 1 2 77742 94502
0 38083 5 1 1 38082
0 38084 7 1 2 73510 38083
0 38085 5 1 1 38084
0 38086 7 1 2 75615 38085
0 38087 5 1 1 38086
0 38088 7 1 2 38081 38087
0 38089 5 1 1 38088
0 38090 7 1 2 70498 38089
0 38091 5 1 1 38090
0 38092 7 1 2 90779 38091
0 38093 7 1 2 38079 38092
0 38094 5 1 1 38093
0 38095 7 1 2 88187 92530
0 38096 7 1 2 38094 38095
0 38097 5 1 1 38096
0 38098 7 1 2 38065 38097
0 38099 5 1 1 38098
0 38100 7 1 2 68983 38099
0 38101 5 1 1 38100
0 38102 7 1 2 82497 89723
0 38103 5 1 1 38102
0 38104 7 1 2 77445 38103
0 38105 5 1 1 38104
0 38106 7 1 2 70196 38105
0 38107 5 1 1 38106
0 38108 7 1 2 77434 83246
0 38109 5 1 1 38108
0 38110 7 1 2 38107 38109
0 38111 5 1 1 38110
0 38112 7 1 2 88994 38111
0 38113 5 1 1 38112
0 38114 7 1 2 77126 95523
0 38115 7 1 2 78099 38114
0 38116 5 1 1 38115
0 38117 7 1 2 92746 38116
0 38118 5 1 1 38117
0 38119 7 1 2 38113 38118
0 38120 5 1 1 38119
0 38121 7 1 2 68425 38120
0 38122 5 1 1 38121
0 38123 7 1 2 67346 76790
0 38124 5 1 1 38123
0 38125 7 1 2 95628 38124
0 38126 5 1 1 38125
0 38127 7 1 2 59572 38126
0 38128 5 1 1 38127
0 38129 7 1 2 76791 69311
0 38130 5 1 1 38129
0 38131 7 1 2 38128 38130
0 38132 5 1 1 38131
0 38133 7 1 2 79795 38132
0 38134 5 1 1 38133
0 38135 7 1 2 38122 38134
0 38136 5 1 1 38135
0 38137 7 1 2 65469 38136
0 38138 5 1 1 38137
0 38139 7 2 2 77679 70914
0 38140 7 1 2 94297 95691
0 38141 5 1 1 38140
0 38142 7 1 2 59573 89727
0 38143 5 1 1 38142
0 38144 7 1 2 59925 87432
0 38145 5 1 1 38144
0 38146 7 2 2 38143 38145
0 38147 5 1 1 95693
0 38148 7 1 2 89679 95694
0 38149 5 1 1 38148
0 38150 7 1 2 61367 38149
0 38151 5 1 1 38150
0 38152 7 1 2 61096 87433
0 38153 5 1 1 38152
0 38154 7 1 2 74743 38153
0 38155 7 1 2 38151 38154
0 38156 5 1 1 38155
0 38157 7 1 2 60164 91609
0 38158 7 1 2 38156 38157
0 38159 5 1 1 38158
0 38160 7 1 2 61583 74626
0 38161 5 1 1 38160
0 38162 7 1 2 14093 38161
0 38163 5 1 1 38162
0 38164 7 1 2 87434 38163
0 38165 5 1 1 38164
0 38166 7 1 2 74204 88159
0 38167 5 1 1 38166
0 38168 7 1 2 38165 38167
0 38169 7 1 2 38159 38168
0 38170 5 1 1 38169
0 38171 7 1 2 60380 38170
0 38172 5 1 1 38171
0 38173 7 1 2 38141 38172
0 38174 5 1 1 38173
0 38175 7 1 2 63523 38174
0 38176 5 1 1 38175
0 38177 7 1 2 38138 38176
0 38178 5 1 1 38177
0 38179 7 3 2 68984 87179
0 38180 7 1 2 38178 95695
0 38181 5 1 1 38180
0 38182 7 1 2 64112 80813
0 38183 7 1 2 74955 38182
0 38184 7 3 2 60677 86355
0 38185 7 3 2 72741 82498
0 38186 7 1 2 89092 95701
0 38187 7 1 2 95698 38186
0 38188 7 1 2 38183 38187
0 38189 5 1 1 38188
0 38190 7 1 2 38181 38189
0 38191 5 1 1 38190
0 38192 7 1 2 69411 38191
0 38193 5 1 1 38192
0 38194 7 7 2 68426 64113
0 38195 7 2 2 91074 95704
0 38196 7 10 2 61878 67090
0 38197 7 1 2 74683 95713
0 38198 7 2 2 95711 38197
0 38199 7 1 2 73062 92301
0 38200 7 1 2 89296 38199
0 38201 7 1 2 95723 38200
0 38202 5 1 1 38201
0 38203 7 1 2 38193 38202
0 38204 7 1 2 38101 38203
0 38205 7 1 2 37703 38204
0 38206 5 1 1 38205
0 38207 7 1 2 61739 38206
0 38208 5 1 1 38207
0 38209 7 1 2 80262 91988
0 38210 5 1 1 38209
0 38211 7 1 2 70234 76031
0 38212 7 1 2 91740 38211
0 38213 5 1 1 38212
0 38214 7 1 2 38210 38213
0 38215 5 1 1 38214
0 38216 7 1 2 94196 38215
0 38217 5 1 1 38216
0 38218 7 1 2 90695 92808
0 38219 5 1 1 38218
0 38220 7 1 2 59362 94197
0 38221 7 1 2 91989 38220
0 38222 5 1 1 38221
0 38223 7 1 2 38219 38222
0 38224 5 1 1 38223
0 38225 7 1 2 74627 38224
0 38226 5 1 1 38225
0 38227 7 1 2 38217 38226
0 38228 5 1 1 38227
0 38229 7 1 2 63108 38228
0 38230 5 1 1 38229
0 38231 7 1 2 63524 92567
0 38232 5 1 1 38231
0 38233 7 1 2 21394 94061
0 38234 5 1 1 38233
0 38235 7 1 2 75330 38234
0 38236 5 1 1 38235
0 38237 7 1 2 78198 86299
0 38238 5 1 1 38237
0 38239 7 1 2 89634 38238
0 38240 7 1 2 38236 38239
0 38241 5 1 1 38240
0 38242 7 1 2 60564 38241
0 38243 5 1 1 38242
0 38244 7 1 2 90067 93244
0 38245 5 1 1 38244
0 38246 7 1 2 38243 38245
0 38247 5 1 1 38246
0 38248 7 1 2 86791 38247
0 38249 5 1 1 38248
0 38250 7 1 2 38232 38249
0 38251 5 1 1 38250
0 38252 7 1 2 72131 38251
0 38253 5 1 1 38252
0 38254 7 1 2 38230 38253
0 38255 5 1 1 38254
0 38256 7 1 2 66728 38255
0 38257 5 1 1 38256
0 38258 7 1 2 75331 95692
0 38259 5 1 1 38258
0 38260 7 1 2 75504 74628
0 38261 5 1 1 38260
0 38262 7 1 2 38259 38261
0 38263 5 1 1 38262
0 38264 7 1 2 95491 38263
0 38265 5 1 1 38264
0 38266 7 1 2 82716 91759
0 38267 5 1 1 38266
0 38268 7 4 2 61097 83746
0 38269 7 1 2 92988 95725
0 38270 5 1 1 38269
0 38271 7 1 2 24507 38270
0 38272 5 1 1 38271
0 38273 7 1 2 60165 74205
0 38274 7 1 2 38272 38273
0 38275 5 1 1 38274
0 38276 7 1 2 38267 38275
0 38277 5 1 1 38276
0 38278 7 1 2 75332 38277
0 38279 5 1 1 38278
0 38280 7 1 2 80147 91760
0 38281 5 1 1 38280
0 38282 7 1 2 83188 91741
0 38283 7 1 2 95521 38282
0 38284 5 1 1 38283
0 38285 7 1 2 38281 38284
0 38286 7 1 2 38279 38285
0 38287 5 1 1 38286
0 38288 7 1 2 66729 38287
0 38289 5 1 1 38288
0 38290 7 1 2 38265 38289
0 38291 5 1 1 38290
0 38292 7 1 2 86792 38291
0 38293 5 1 1 38292
0 38294 7 1 2 38257 38293
0 38295 5 1 1 38294
0 38296 7 1 2 68985 38295
0 38297 5 1 1 38296
0 38298 7 2 2 73468 91404
0 38299 7 3 2 60678 60936
0 38300 7 1 2 87034 95731
0 38301 7 1 2 95702 38300
0 38302 7 1 2 95729 38301
0 38303 7 1 2 95712 38302
0 38304 5 1 1 38303
0 38305 7 1 2 38297 38304
0 38306 5 1 1 38305
0 38307 7 1 2 69412 38306
0 38308 5 1 1 38307
0 38309 7 1 2 80459 92356
0 38310 7 1 2 89993 38309
0 38311 7 1 2 95724 38310
0 38312 5 1 1 38311
0 38313 7 1 2 38308 38312
0 38314 7 1 2 38208 38313
0 38315 7 1 2 37045 38314
0 38316 5 1 1 38315
0 38317 7 1 2 68721 38316
0 38318 5 1 1 38317
0 38319 7 3 2 87180 89317
0 38320 5 1 1 95734
0 38321 7 1 2 87719 38320
0 38322 5 1 1 38321
0 38323 7 2 2 95519 38322
0 38324 5 1 1 95737
0 38325 7 2 2 75333 87493
0 38326 7 1 2 95614 95739
0 38327 5 1 1 38326
0 38328 7 1 2 38324 38327
0 38329 5 1 1 38328
0 38330 7 1 2 94207 38329
0 38331 5 1 1 38330
0 38332 7 6 2 60679 64114
0 38333 7 1 2 69190 95741
0 38334 7 1 2 93027 38333
0 38335 7 3 2 59926 71396
0 38336 7 2 2 60565 86276
0 38337 7 1 2 95747 95750
0 38338 7 1 2 38334 38337
0 38339 5 1 1 38338
0 38340 7 1 2 38331 38339
0 38341 5 1 1 38340
0 38342 7 1 2 73381 38341
0 38343 5 1 1 38342
0 38344 7 1 2 75616 81360
0 38345 5 1 1 38344
0 38346 7 1 2 95740 38345
0 38347 5 1 1 38346
0 38348 7 1 2 87723 38347
0 38349 5 1 1 38348
0 38350 7 1 2 68986 83585
0 38351 7 1 2 91544 38350
0 38352 7 1 2 38349 38351
0 38353 5 1 1 38352
0 38354 7 1 2 38343 38353
0 38355 5 1 1 38354
0 38356 7 1 2 78262 38355
0 38357 5 1 1 38356
0 38358 7 2 2 86623 87212
0 38359 5 1 1 95752
0 38360 7 1 2 77478 85046
0 38361 5 2 1 38360
0 38362 7 1 2 74570 76980
0 38363 5 1 1 38362
0 38364 7 1 2 70627 90651
0 38365 7 1 2 38363 38364
0 38366 5 1 1 38365
0 38367 7 1 2 65734 38366
0 38368 5 1 1 38367
0 38369 7 1 2 68055 38368
0 38370 5 1 1 38369
0 38371 7 1 2 64319 38370
0 38372 5 1 1 38371
0 38373 7 1 2 62145 82722
0 38374 5 1 1 38373
0 38375 7 1 2 74206 78940
0 38376 5 1 1 38375
0 38377 7 1 2 82466 38376
0 38378 5 1 1 38377
0 38379 7 1 2 38374 38378
0 38380 7 1 2 38372 38379
0 38381 5 1 1 38380
0 38382 7 1 2 62721 38381
0 38383 5 1 1 38382
0 38384 7 1 2 80069 70456
0 38385 5 1 1 38384
0 38386 7 1 2 60166 38385
0 38387 5 1 1 38386
0 38388 7 1 2 62722 38387
0 38389 5 1 1 38388
0 38390 7 1 2 70931 88865
0 38391 5 1 1 38390
0 38392 7 1 2 64790 38391
0 38393 5 1 1 38392
0 38394 7 1 2 80591 38393
0 38395 5 1 1 38394
0 38396 7 1 2 70371 38395
0 38397 5 1 1 38396
0 38398 7 1 2 76877 15620
0 38399 5 1 1 38398
0 38400 7 1 2 76706 38399
0 38401 5 1 1 38400
0 38402 7 1 2 70826 88777
0 38403 5 1 1 38402
0 38404 7 1 2 38401 38403
0 38405 7 1 2 38397 38404
0 38406 7 1 2 38389 38405
0 38407 5 1 1 38406
0 38408 7 1 2 62368 38407
0 38409 5 1 1 38408
0 38410 7 1 2 78665 95392
0 38411 5 1 1 38410
0 38412 7 2 2 64791 90286
0 38413 5 1 1 95756
0 38414 7 1 2 86606 38413
0 38415 5 1 1 38414
0 38416 7 1 2 73525 38415
0 38417 5 1 1 38416
0 38418 7 1 2 77502 38417
0 38419 5 1 1 38418
0 38420 7 1 2 70323 38419
0 38421 5 1 1 38420
0 38422 7 1 2 38411 38421
0 38423 7 1 2 38409 38422
0 38424 7 1 2 38383 38423
0 38425 5 1 1 38424
0 38426 7 1 2 75617 38425
0 38427 5 1 1 38426
0 38428 7 1 2 95754 38427
0 38429 5 1 1 38428
0 38430 7 1 2 65470 38429
0 38431 5 1 1 38430
0 38432 7 1 2 66060 90317
0 38433 5 1 1 38432
0 38434 7 1 2 89161 38433
0 38435 5 1 1 38434
0 38436 7 1 2 66336 38435
0 38437 5 1 1 38436
0 38438 7 1 2 64320 93370
0 38439 5 1 1 38438
0 38440 7 1 2 38437 38439
0 38441 5 1 1 38440
0 38442 7 1 2 73580 38441
0 38443 5 1 1 38442
0 38444 7 1 2 64792 90301
0 38445 5 1 1 38444
0 38446 7 1 2 60167 38445
0 38447 5 1 1 38446
0 38448 7 1 2 77708 38447
0 38449 5 1 1 38448
0 38450 7 1 2 70265 90960
0 38451 5 1 1 38450
0 38452 7 1 2 87029 38451
0 38453 5 1 1 38452
0 38454 7 1 2 38449 38453
0 38455 5 1 1 38454
0 38456 7 1 2 71824 38455
0 38457 5 1 1 38456
0 38458 7 1 2 64321 71929
0 38459 5 2 1 38458
0 38460 7 1 2 90441 95758
0 38461 5 1 1 38460
0 38462 7 1 2 82047 38461
0 38463 5 1 1 38462
0 38464 7 1 2 77310 95759
0 38465 5 1 1 38464
0 38466 7 1 2 82723 38465
0 38467 5 1 1 38466
0 38468 7 1 2 13286 38467
0 38469 5 1 1 38468
0 38470 7 1 2 66337 38469
0 38471 5 1 1 38470
0 38472 7 1 2 38463 38471
0 38473 7 1 2 38457 38472
0 38474 7 1 2 38443 38473
0 38475 5 1 1 38474
0 38476 7 1 2 63109 38475
0 38477 5 1 1 38476
0 38478 7 1 2 60168 84912
0 38479 5 1 1 38478
0 38480 7 1 2 63110 38479
0 38481 5 1 1 38480
0 38482 7 1 2 63111 76011
0 38483 5 1 1 38482
0 38484 7 1 2 68056 80655
0 38485 5 2 1 38484
0 38486 7 1 2 73526 95760
0 38487 5 1 1 38486
0 38488 7 1 2 38483 38487
0 38489 5 1 1 38488
0 38490 7 1 2 64793 38489
0 38491 5 1 1 38490
0 38492 7 1 2 38481 38491
0 38493 5 1 1 38492
0 38494 7 1 2 66338 38493
0 38495 5 1 1 38494
0 38496 7 1 2 73584 77479
0 38497 5 1 1 38496
0 38498 7 1 2 38495 38497
0 38499 5 1 1 38498
0 38500 7 1 2 66061 38499
0 38501 5 1 1 38500
0 38502 7 1 2 77480 95015
0 38503 5 1 1 38502
0 38504 7 1 2 38501 38503
0 38505 5 1 1 38504
0 38506 7 1 2 70324 38505
0 38507 5 1 1 38506
0 38508 7 1 2 62723 91372
0 38509 5 1 1 38508
0 38510 7 1 2 93781 38509
0 38511 5 1 1 38510
0 38512 7 1 2 65735 38511
0 38513 5 1 1 38512
0 38514 7 1 2 91005 38513
0 38515 5 1 1 38514
0 38516 7 1 2 64794 38515
0 38517 5 1 1 38516
0 38518 7 1 2 70950 70937
0 38519 5 1 1 38518
0 38520 7 1 2 38517 38519
0 38521 5 1 1 38520
0 38522 7 1 2 70068 38521
0 38523 5 1 1 38522
0 38524 7 1 2 38507 38523
0 38525 7 1 2 38477 38524
0 38526 5 1 1 38525
0 38527 7 1 2 91858 38526
0 38528 5 1 1 38527
0 38529 7 1 2 70069 94807
0 38530 5 1 1 38529
0 38531 7 1 2 70070 80212
0 38532 5 1 1 38531
0 38533 7 1 2 80595 76725
0 38534 5 1 1 38533
0 38535 7 1 2 38532 38534
0 38536 5 1 1 38535
0 38537 7 1 2 62369 38536
0 38538 5 1 1 38537
0 38539 7 1 2 38530 38538
0 38540 5 1 1 38539
0 38541 7 1 2 91859 38540
0 38542 5 1 1 38541
0 38543 7 2 2 94844 95274
0 38544 7 1 2 64795 78362
0 38545 5 2 1 38544
0 38546 7 1 2 70628 95764
0 38547 7 1 2 95762 38546
0 38548 5 1 1 38547
0 38549 7 1 2 91659 38548
0 38550 5 1 1 38549
0 38551 7 1 2 38542 38550
0 38552 5 1 1 38551
0 38553 7 1 2 89051 38552
0 38554 5 1 1 38553
0 38555 7 1 2 73181 78941
0 38556 5 1 1 38555
0 38557 7 1 2 80699 91660
0 38558 5 1 1 38557
0 38559 7 1 2 70556 95763
0 38560 5 1 1 38559
0 38561 7 2 2 82824 38560
0 38562 7 1 2 65021 91860
0 38563 7 1 2 95766 38562
0 38564 5 1 1 38563
0 38565 7 1 2 38558 38564
0 38566 5 1 1 38565
0 38567 7 1 2 38556 38566
0 38568 5 1 1 38567
0 38569 7 1 2 72015 72496
0 38570 5 1 1 38569
0 38571 7 1 2 70897 38570
0 38572 5 2 1 38571
0 38573 7 1 2 88466 95768
0 38574 5 1 1 38573
0 38575 7 1 2 60381 71854
0 38576 7 1 2 38574 38575
0 38577 5 2 1 38576
0 38578 7 1 2 65471 95770
0 38579 5 1 1 38578
0 38580 7 1 2 72016 71280
0 38581 7 1 2 88467 38580
0 38582 5 1 1 38581
0 38583 7 1 2 38579 38582
0 38584 5 1 1 38583
0 38585 7 1 2 91316 38584
0 38586 5 1 1 38585
0 38587 7 1 2 60566 95755
0 38588 5 1 1 38587
0 38589 7 1 2 72017 95646
0 38590 5 1 1 38589
0 38591 7 1 2 94708 38590
0 38592 5 1 1 38591
0 38593 7 1 2 88468 38592
0 38594 5 1 1 38593
0 38595 7 1 2 93324 38594
0 38596 5 1 1 38595
0 38597 7 1 2 38588 38596
0 38598 5 1 1 38597
0 38599 7 1 2 61740 38598
0 38600 7 1 2 38586 38599
0 38601 7 1 2 38568 38600
0 38602 7 1 2 38554 38601
0 38603 7 1 2 38528 38602
0 38604 7 1 2 38431 38603
0 38605 5 1 1 38604
0 38606 7 1 2 60567 95771
0 38607 5 1 1 38606
0 38608 7 1 2 76792 92184
0 38609 5 1 1 38608
0 38610 7 1 2 38607 38609
0 38611 5 1 1 38610
0 38612 7 1 2 62724 38611
0 38613 5 1 1 38612
0 38614 7 2 2 81059 87831
0 38615 7 2 2 80278 95772
0 38616 7 1 2 95354 95774
0 38617 5 1 1 38616
0 38618 7 1 2 79085 94583
0 38619 5 1 1 38618
0 38620 7 1 2 72617 76735
0 38621 5 1 1 38620
0 38622 7 1 2 38619 38621
0 38623 5 1 1 38622
0 38624 7 1 2 82616 38623
0 38625 5 1 1 38624
0 38626 7 1 2 38617 38625
0 38627 7 1 2 38613 38626
0 38628 5 1 1 38627
0 38629 7 1 2 62370 38628
0 38630 5 1 1 38629
0 38631 7 1 2 73798 93358
0 38632 5 2 1 38631
0 38633 7 1 2 88167 23217
0 38634 5 1 1 38633
0 38635 7 1 2 64796 38634
0 38636 5 1 1 38635
0 38637 7 1 2 60568 73799
0 38638 5 1 1 38637
0 38639 7 1 2 38636 38638
0 38640 5 3 1 38639
0 38641 7 1 2 72018 95778
0 38642 5 1 1 38641
0 38643 7 1 2 95776 38642
0 38644 5 1 1 38643
0 38645 7 1 2 70827 38644
0 38646 5 1 1 38645
0 38647 7 1 2 71576 88163
0 38648 5 1 1 38647
0 38649 7 1 2 78666 95775
0 38650 5 1 1 38649
0 38651 7 1 2 38648 38650
0 38652 7 1 2 38646 38651
0 38653 5 1 1 38652
0 38654 7 1 2 73211 38653
0 38655 5 1 1 38654
0 38656 7 1 2 73230 95779
0 38657 5 1 1 38656
0 38658 7 1 2 95777 38657
0 38659 5 1 1 38658
0 38660 7 1 2 70828 38659
0 38661 5 1 1 38660
0 38662 7 1 2 89369 95773
0 38663 5 1 1 38662
0 38664 7 1 2 88168 38663
0 38665 5 1 1 38664
0 38666 7 1 2 80279 38665
0 38667 5 1 1 38666
0 38668 7 1 2 38661 38667
0 38669 5 1 1 38668
0 38670 7 1 2 71825 38669
0 38671 5 1 1 38670
0 38672 7 1 2 71577 95780
0 38673 5 1 1 38672
0 38674 7 1 2 72422 13662
0 38675 5 1 1 38674
0 38676 7 1 2 70629 38675
0 38677 5 1 1 38676
0 38678 7 1 2 60569 21057
0 38679 7 1 2 38677 38678
0 38680 5 1 1 38679
0 38681 7 1 2 38673 38680
0 38682 7 1 2 38671 38681
0 38683 7 1 2 38655 38682
0 38684 7 1 2 38630 38683
0 38685 5 1 1 38684
0 38686 7 1 2 63112 38685
0 38687 5 1 1 38686
0 38688 7 2 2 65736 76647
0 38689 5 2 1 95781
0 38690 7 1 2 71231 95783
0 38691 5 1 1 38690
0 38692 7 1 2 62146 38691
0 38693 5 1 1 38692
0 38694 7 1 2 65737 90876
0 38695 5 1 1 38694
0 38696 7 1 2 38693 38695
0 38697 5 1 1 38696
0 38698 7 1 2 65891 38697
0 38699 5 1 1 38698
0 38700 7 1 2 62725 89238
0 38701 5 1 1 38700
0 38702 7 1 2 65738 85089
0 38703 5 1 1 38702
0 38704 7 1 2 62371 95567
0 38705 5 1 1 38704
0 38706 7 1 2 38703 38705
0 38707 5 2 1 38706
0 38708 7 1 2 64797 95785
0 38709 5 1 1 38708
0 38710 7 1 2 38701 38709
0 38711 7 1 2 38699 38710
0 38712 5 1 1 38711
0 38713 7 1 2 64322 38712
0 38714 5 1 1 38713
0 38715 7 1 2 73065 88415
0 38716 5 1 1 38715
0 38717 7 1 2 93254 38716
0 38718 5 1 1 38717
0 38719 7 1 2 62372 38718
0 38720 5 1 1 38719
0 38721 7 1 2 84095 94701
0 38722 5 1 1 38721
0 38723 7 1 2 88818 38722
0 38724 7 1 2 38720 38723
0 38725 7 1 2 38714 38724
0 38726 5 1 1 38725
0 38727 7 1 2 64560 38726
0 38728 5 1 1 38727
0 38729 7 1 2 81601 88554
0 38730 5 1 1 38729
0 38731 7 1 2 62726 38730
0 38732 5 1 1 38731
0 38733 7 1 2 90668 38732
0 38734 5 2 1 38733
0 38735 7 1 2 70829 95787
0 38736 5 1 1 38735
0 38737 7 1 2 64798 70426
0 38738 5 2 1 38737
0 38739 7 1 2 73021 72522
0 38740 5 3 1 38739
0 38741 7 1 2 71122 95791
0 38742 5 1 1 38741
0 38743 7 1 2 89233 38742
0 38744 7 1 2 95789 38743
0 38745 5 1 1 38744
0 38746 7 1 2 62727 38745
0 38747 5 1 1 38746
0 38748 7 1 2 78515 94792
0 38749 5 1 1 38748
0 38750 7 1 2 71523 38749
0 38751 7 1 2 38747 38750
0 38752 7 1 2 38736 38751
0 38753 7 1 2 38728 38752
0 38754 5 1 1 38753
0 38755 7 1 2 85455 38754
0 38756 5 1 1 38755
0 38757 7 1 2 1843 83705
0 38758 5 1 1 38757
0 38759 7 1 2 72612 38758
0 38760 5 1 1 38759
0 38761 7 1 2 83716 89027
0 38762 5 2 1 38761
0 38763 7 1 2 83717 77520
0 38764 5 1 1 38763
0 38765 7 1 2 95794 38764
0 38766 7 1 2 38760 38765
0 38767 5 1 1 38766
0 38768 7 1 2 66730 38767
0 38769 7 1 2 38756 38768
0 38770 7 1 2 38687 38769
0 38771 5 1 1 38770
0 38772 7 1 2 61879 38771
0 38773 7 1 2 38605 38772
0 38774 5 1 1 38773
0 38775 7 1 2 38359 38774
0 38776 5 1 1 38775
0 38777 7 1 2 60680 38776
0 38778 5 1 1 38777
0 38779 7 1 2 74865 77517
0 38780 5 3 1 38779
0 38781 7 1 2 65472 81602
0 38782 5 1 1 38781
0 38783 7 1 2 95796 38782
0 38784 5 1 1 38783
0 38785 7 1 2 69937 38784
0 38786 5 1 1 38785
0 38787 7 1 2 90904 95797
0 38788 5 1 1 38787
0 38789 7 1 2 60937 38788
0 38790 5 1 1 38789
0 38791 7 1 2 38786 38790
0 38792 5 1 1 38791
0 38793 7 1 2 59927 38792
0 38794 5 1 1 38793
0 38795 7 1 2 91775 92651
0 38796 5 1 1 38795
0 38797 7 1 2 38794 38796
0 38798 5 1 1 38797
0 38799 7 1 2 85847 38798
0 38800 5 1 1 38799
0 38801 7 1 2 81878 72148
0 38802 7 1 2 95792 38801
0 38803 5 1 1 38802
0 38804 7 2 2 89318 38803
0 38805 7 1 2 86138 95799
0 38806 5 1 1 38805
0 38807 7 1 2 38800 38806
0 38808 5 1 1 38807
0 38809 7 1 2 60681 38808
0 38810 5 1 1 38809
0 38811 7 1 2 71335 95735
0 38812 5 1 1 38811
0 38813 7 1 2 71292 87717
0 38814 5 1 1 38813
0 38815 7 1 2 38812 38814
0 38816 5 1 1 38815
0 38817 7 1 2 67690 38816
0 38818 5 1 1 38817
0 38819 7 1 2 67347 77481
0 38820 7 2 2 85808 38819
0 38821 7 1 2 87017 89059
0 38822 7 1 2 95801 38821
0 38823 5 1 1 38822
0 38824 7 1 2 38818 38823
0 38825 5 1 1 38824
0 38826 7 1 2 71232 38825
0 38827 5 1 1 38826
0 38828 7 5 2 59928 65602
0 38829 7 1 2 61880 95803
0 38830 7 1 2 95800 38829
0 38831 5 1 1 38830
0 38832 7 1 2 38827 38831
0 38833 7 1 2 38810 38832
0 38834 5 1 1 38833
0 38835 7 1 2 59574 38834
0 38836 5 1 1 38835
0 38837 7 1 2 75334 87725
0 38838 5 1 1 38837
0 38839 7 1 2 1822 95563
0 38840 5 1 1 38839
0 38841 7 1 2 95736 38840
0 38842 5 1 1 38841
0 38843 7 1 2 11894 95798
0 38844 5 1 1 38843
0 38845 7 2 2 69938 92309
0 38846 7 1 2 61881 95808
0 38847 7 1 2 38844 38846
0 38848 5 1 1 38847
0 38849 7 1 2 38842 38848
0 38850 5 1 1 38849
0 38851 7 1 2 60938 38850
0 38852 5 1 1 38851
0 38853 7 6 2 60682 69573
0 38854 7 1 2 74866 95810
0 38855 7 1 2 95802 38854
0 38856 5 1 1 38855
0 38857 7 1 2 38852 38856
0 38858 5 1 1 38857
0 38859 7 1 2 59929 38858
0 38860 5 1 1 38859
0 38861 7 1 2 38838 38860
0 38862 7 1 2 38836 38861
0 38863 5 1 1 38862
0 38864 7 1 2 70197 38863
0 38865 5 1 1 38864
0 38866 7 1 2 72019 94702
0 38867 5 1 1 38866
0 38868 7 2 2 81700 38867
0 38869 5 1 1 95816
0 38870 7 1 2 69697 73527
0 38871 5 1 1 38870
0 38872 7 1 2 67691 38871
0 38873 7 1 2 12710 38872
0 38874 5 1 1 38873
0 38875 7 1 2 70830 38874
0 38876 5 1 1 38875
0 38877 7 1 2 95817 38876
0 38878 5 1 1 38877
0 38879 7 1 2 62147 38878
0 38880 5 1 1 38879
0 38881 7 1 2 69857 73528
0 38882 5 1 1 38881
0 38883 7 1 2 73826 38882
0 38884 5 1 1 38883
0 38885 7 1 2 70831 38884
0 38886 5 1 1 38885
0 38887 7 1 2 70198 38886
0 38888 7 1 2 38880 38887
0 38889 5 1 1 38888
0 38890 7 1 2 65270 38889
0 38891 5 1 1 38890
0 38892 7 1 2 69738 90258
0 38893 5 3 1 38892
0 38894 7 1 2 64323 95786
0 38895 5 2 1 38894
0 38896 7 1 2 66062 69456
0 38897 5 1 1 38896
0 38898 7 1 2 78080 38897
0 38899 7 1 2 95821 38898
0 38900 5 1 1 38899
0 38901 7 1 2 64799 38900
0 38902 5 1 1 38901
0 38903 7 1 2 95818 38902
0 38904 5 1 1 38903
0 38905 7 1 2 95388 38904
0 38906 5 1 1 38905
0 38907 7 1 2 61368 95784
0 38908 5 1 1 38907
0 38909 7 1 2 65271 72361
0 38910 5 1 1 38909
0 38911 7 1 2 72020 77196
0 38912 5 1 1 38911
0 38913 7 1 2 38910 38912
0 38914 5 1 1 38913
0 38915 7 1 2 79834 38914
0 38916 5 1 1 38915
0 38917 7 1 2 71826 79542
0 38918 5 1 1 38917
0 38919 7 1 2 38916 38918
0 38920 5 1 1 38919
0 38921 7 1 2 38908 38920
0 38922 5 1 1 38921
0 38923 7 1 2 76751 94925
0 38924 5 1 1 38923
0 38925 7 1 2 73879 88308
0 38926 5 1 1 38925
0 38927 7 1 2 38924 38926
0 38928 5 1 1 38927
0 38929 7 1 2 71930 38928
0 38930 5 1 1 38929
0 38931 7 1 2 60382 94571
0 38932 5 1 1 38931
0 38933 7 1 2 79835 95086
0 38934 5 1 1 38933
0 38935 7 1 2 8379 38934
0 38936 5 1 1 38935
0 38937 7 1 2 38932 38936
0 38938 5 1 1 38937
0 38939 7 1 2 76860 38869
0 38940 5 1 1 38939
0 38941 7 1 2 65272 73854
0 38942 5 1 1 38941
0 38943 7 1 2 60169 38942
0 38944 5 1 1 38943
0 38945 7 1 2 60383 18692
0 38946 5 1 1 38945
0 38947 7 1 2 92941 38946
0 38948 7 1 2 38944 38947
0 38949 5 1 1 38948
0 38950 7 1 2 38940 38949
0 38951 7 1 2 38938 38950
0 38952 7 1 2 38930 38951
0 38953 7 1 2 38922 38952
0 38954 7 1 2 38906 38953
0 38955 7 1 2 38891 38954
0 38956 5 1 1 38955
0 38957 7 1 2 87035 92310
0 38958 7 1 2 38956 38957
0 38959 5 1 1 38958
0 38960 7 1 2 66063 82810
0 38961 5 2 1 38960
0 38962 7 1 2 71420 90468
0 38963 7 1 2 95823 38962
0 38964 5 1 1 38963
0 38965 7 1 2 75618 38964
0 38966 5 1 1 38965
0 38967 7 4 2 70630 79651
0 38968 7 1 2 38966 95825
0 38969 5 1 1 38968
0 38970 7 1 2 88140 38969
0 38971 5 1 1 38970
0 38972 7 1 2 87181 38971
0 38973 5 1 1 38972
0 38974 7 1 2 76793 87726
0 38975 5 1 1 38974
0 38976 7 1 2 95738 95824
0 38977 5 1 1 38976
0 38978 7 1 2 38975 38977
0 38979 7 1 2 38973 38978
0 38980 7 1 2 38959 38979
0 38981 5 1 1 38980
0 38982 7 1 2 68057 38981
0 38983 5 1 1 38982
0 38984 7 1 2 65473 84020
0 38985 5 1 1 38984
0 38986 7 2 2 85605 89261
0 38987 5 1 1 95829
0 38988 7 1 2 38985 38987
0 38989 5 1 1 38988
0 38990 7 1 2 92320 38989
0 38991 5 1 1 38990
0 38992 7 1 2 80904 93347
0 38993 5 1 1 38992
0 38994 7 1 2 71500 87494
0 38995 7 1 2 38993 38994
0 38996 5 1 1 38995
0 38997 7 1 2 38991 38996
0 38998 5 1 1 38997
0 38999 7 1 2 76794 38998
0 39000 5 1 1 38999
0 39001 7 1 2 80905 4169
0 39002 5 2 1 39001
0 39003 7 5 2 79652 95831
0 39004 7 1 2 87182 95833
0 39005 5 1 1 39004
0 39006 7 1 2 87720 39005
0 39007 5 1 1 39006
0 39008 7 1 2 71501 93352
0 39009 7 1 2 39007 39008
0 39010 5 1 1 39009
0 39011 7 1 2 39000 39010
0 39012 5 1 1 39011
0 39013 7 1 2 67348 39012
0 39014 5 1 1 39013
0 39015 7 1 2 345 87183
0 39016 7 1 2 91901 39015
0 39017 5 1 1 39016
0 39018 7 3 2 86277 92119
0 39019 7 1 2 65603 95838
0 39020 5 2 1 39019
0 39021 7 1 2 39017 95841
0 39022 7 1 2 39014 39021
0 39023 7 1 2 38983 39022
0 39024 7 1 2 38865 39023
0 39025 7 1 2 38778 39024
0 39026 5 1 1 39025
0 39027 7 1 2 94208 39026
0 39028 5 1 1 39027
0 39029 7 1 2 38357 39028
0 39030 5 1 1 39029
0 39031 7 1 2 68427 39030
0 39032 5 1 1 39031
0 39033 7 1 2 75619 359
0 39034 5 1 1 39033
0 39035 7 1 2 91849 39034
0 39036 5 1 1 39035
0 39037 7 1 2 61741 39036
0 39038 5 1 1 39037
0 39039 7 1 2 80774 93448
0 39040 5 1 1 39039
0 39041 7 1 2 39038 39040
0 39042 5 1 1 39041
0 39043 7 1 2 62148 39042
0 39044 5 1 1 39043
0 39045 7 1 2 61742 90409
0 39046 5 1 1 39045
0 39047 7 1 2 81197 39046
0 39048 5 2 1 39047
0 39049 7 1 2 88759 95843
0 39050 5 1 1 39049
0 39051 7 2 2 61743 91312
0 39052 7 1 2 80588 78469
0 39053 7 1 2 95845 39052
0 39054 5 1 1 39053
0 39055 7 1 2 39050 39054
0 39056 7 1 2 39044 39055
0 39057 5 1 1 39056
0 39058 7 1 2 62373 39057
0 39059 5 1 1 39058
0 39060 7 1 2 94584 95844
0 39061 5 1 1 39060
0 39062 7 1 2 82713 95846
0 39063 7 1 2 94923 39062
0 39064 5 1 1 39063
0 39065 7 1 2 75460 94152
0 39066 5 1 1 39065
0 39067 7 1 2 67692 39066
0 39068 7 1 2 39064 39067
0 39069 7 1 2 39061 39068
0 39070 7 1 2 39059 39069
0 39071 5 1 1 39070
0 39072 7 1 2 61584 95647
0 39073 5 1 1 39072
0 39074 7 1 2 72497 85456
0 39075 5 1 1 39074
0 39076 7 1 2 39073 39075
0 39077 5 1 1 39076
0 39078 7 1 2 73114 39077
0 39079 5 1 1 39078
0 39080 7 1 2 67349 91352
0 39081 5 1 1 39080
0 39082 7 1 2 39079 39081
0 39083 5 1 1 39082
0 39084 7 1 2 72847 39083
0 39085 5 1 1 39084
0 39086 7 1 2 88641 93201
0 39087 5 1 1 39086
0 39088 7 1 2 80131 27572
0 39089 5 2 1 39088
0 39090 7 1 2 75620 95847
0 39091 7 1 2 88784 39090
0 39092 5 1 1 39091
0 39093 7 1 2 39087 39092
0 39094 5 1 1 39093
0 39095 7 1 2 70832 39094
0 39096 5 1 1 39095
0 39097 7 2 2 76919 78005
0 39098 7 1 2 84649 95849
0 39099 5 1 1 39098
0 39100 7 1 2 65474 39099
0 39101 5 1 1 39100
0 39102 7 1 2 76831 79244
0 39103 7 1 2 80280 39102
0 39104 7 1 2 95848 39103
0 39105 5 1 1 39104
0 39106 7 1 2 17936 39105
0 39107 7 1 2 39101 39106
0 39108 7 1 2 39096 39107
0 39109 7 1 2 39085 39108
0 39110 5 1 1 39109
0 39111 7 1 2 61744 39110
0 39112 5 1 1 39111
0 39113 7 1 2 91861 95850
0 39114 5 1 1 39113
0 39115 7 1 2 91674 39114
0 39116 5 1 1 39115
0 39117 7 1 2 76920 72498
0 39118 5 1 1 39117
0 39119 7 1 2 75335 81363
0 39120 7 1 2 39118 39119
0 39121 5 1 1 39120
0 39122 7 1 2 39116 39121
0 39123 5 1 1 39122
0 39124 7 1 2 66731 39123
0 39125 5 1 1 39124
0 39126 7 1 2 62728 39125
0 39127 7 1 2 39112 39126
0 39128 5 1 1 39127
0 39129 7 1 2 63113 39128
0 39130 7 1 2 39071 39129
0 39131 5 1 1 39130
0 39132 7 1 2 88086 90896
0 39133 5 1 1 39132
0 39134 7 1 2 80346 89758
0 39135 5 4 1 39134
0 39136 7 1 2 77503 95851
0 39137 5 1 1 39136
0 39138 7 1 2 67091 92961
0 39139 5 1 1 39138
0 39140 7 1 2 88393 39139
0 39141 5 1 1 39140
0 39142 7 1 2 91642 39141
0 39143 5 1 1 39142
0 39144 7 1 2 93122 95590
0 39145 5 1 1 39144
0 39146 7 1 2 71658 39145
0 39147 5 1 1 39146
0 39148 7 1 2 39143 39147
0 39149 5 1 1 39148
0 39150 7 1 2 67693 39149
0 39151 5 1 1 39150
0 39152 7 2 2 68058 73257
0 39153 7 1 2 76151 93163
0 39154 5 1 1 39153
0 39155 7 1 2 65273 73929
0 39156 5 1 1 39155
0 39157 7 1 2 92490 39156
0 39158 5 1 1 39157
0 39159 7 1 2 39154 39158
0 39160 5 1 1 39159
0 39161 7 1 2 95855 39160
0 39162 5 1 1 39161
0 39163 7 1 2 39151 39162
0 39164 5 1 1 39163
0 39165 7 1 2 66732 39164
0 39166 5 1 1 39165
0 39167 7 1 2 39137 39166
0 39168 7 1 2 39133 39167
0 39169 5 1 1 39168
0 39170 7 1 2 66561 39169
0 39171 5 1 1 39170
0 39172 7 2 2 71233 88499
0 39173 5 1 1 95857
0 39174 7 1 2 62729 39173
0 39175 5 1 1 39174
0 39176 7 1 2 64800 73989
0 39177 5 1 1 39176
0 39178 7 1 2 91006 39177
0 39179 5 1 1 39178
0 39180 7 1 2 88469 39179
0 39181 5 1 1 39180
0 39182 7 1 2 72160 74613
0 39183 5 1 1 39182
0 39184 7 1 2 39181 39183
0 39185 7 1 2 39175 39184
0 39186 5 1 1 39185
0 39187 7 1 2 70071 39186
0 39188 5 1 1 39187
0 39189 7 3 2 62374 88510
0 39190 5 1 1 95859
0 39191 7 1 2 85415 95860
0 39192 5 1 1 39191
0 39193 7 1 2 39188 39192
0 39194 5 2 1 39193
0 39195 7 1 2 91370 95862
0 39196 5 1 1 39195
0 39197 7 1 2 89376 94511
0 39198 5 1 1 39197
0 39199 7 1 2 62375 39198
0 39200 5 1 1 39199
0 39201 7 1 2 74073 72499
0 39202 5 2 1 39201
0 39203 7 1 2 89389 95864
0 39204 5 1 1 39203
0 39205 7 1 2 88470 39204
0 39206 5 1 1 39205
0 39207 7 1 2 82881 91241
0 39208 5 1 1 39207
0 39209 7 1 2 60384 76152
0 39210 7 1 2 89391 39209
0 39211 7 1 2 39208 39210
0 39212 7 1 2 39206 39211
0 39213 7 1 2 39200 39212
0 39214 5 2 1 39213
0 39215 7 1 2 63114 74252
0 39216 5 1 1 39215
0 39217 7 1 2 80425 39216
0 39218 7 1 2 95866 39217
0 39219 5 1 1 39218
0 39220 7 1 2 39196 39219
0 39221 7 1 2 39171 39220
0 39222 7 1 2 39131 39221
0 39223 5 1 1 39222
0 39224 7 1 2 63525 39223
0 39225 5 1 1 39224
0 39226 7 1 2 67694 74694
0 39227 5 1 1 39226
0 39228 7 5 2 68059 71421
0 39229 7 1 2 59575 95868
0 39230 5 1 1 39229
0 39231 7 1 2 39227 39230
0 39232 5 1 1 39231
0 39233 7 1 2 67350 39232
0 39234 5 1 1 39233
0 39235 7 3 2 68060 88843
0 39236 5 2 1 95873
0 39237 7 1 2 59576 95874
0 39238 5 1 1 39237
0 39239 7 1 2 39234 39238
0 39240 5 1 1 39239
0 39241 7 1 2 69413 39240
0 39242 5 1 1 39241
0 39243 7 2 2 59930 88948
0 39244 5 3 1 95878
0 39245 7 1 2 78238 95880
0 39246 5 2 1 39245
0 39247 7 1 2 69191 95883
0 39248 5 1 1 39247
0 39249 7 1 2 95876 39248
0 39250 5 1 1 39249
0 39251 7 1 2 59363 39250
0 39252 5 1 1 39251
0 39253 7 1 2 71234 78235
0 39254 5 1 1 39253
0 39255 7 1 2 39252 39254
0 39256 5 1 1 39255
0 39257 7 1 2 76050 39256
0 39258 5 1 1 39257
0 39259 7 2 2 65892 83606
0 39260 5 2 1 95885
0 39261 7 1 2 82246 73511
0 39262 5 1 1 39261
0 39263 7 1 2 70256 39262
0 39264 5 1 1 39263
0 39265 7 1 2 95887 39264
0 39266 5 1 1 39265
0 39267 7 1 2 73447 74695
0 39268 5 1 1 39267
0 39269 7 1 2 88589 39268
0 39270 7 1 2 39266 39269
0 39271 5 1 1 39270
0 39272 7 1 2 67695 39271
0 39273 5 1 1 39272
0 39274 7 1 2 76795 77504
0 39275 5 1 1 39274
0 39276 7 1 2 39273 39275
0 39277 7 1 2 39258 39276
0 39278 7 1 2 39242 39277
0 39279 5 1 1 39278
0 39280 7 1 2 83727 39279
0 39281 5 1 1 39280
0 39282 7 1 2 60683 39281
0 39283 7 1 2 39225 39282
0 39284 5 1 1 39283
0 39285 7 1 2 80757 78579
0 39286 7 1 2 83856 39285
0 39287 5 1 1 39286
0 39288 7 1 2 75505 39287
0 39289 5 1 1 39288
0 39290 7 1 2 91778 13588
0 39291 5 1 1 39290
0 39292 7 1 2 71422 39291
0 39293 5 1 1 39292
0 39294 7 1 2 69472 24602
0 39295 5 1 1 39294
0 39296 7 1 2 78401 39295
0 39297 5 1 1 39296
0 39298 7 1 2 95877 39297
0 39299 7 1 2 39293 39298
0 39300 5 1 1 39299
0 39301 7 1 2 59577 39300
0 39302 5 1 1 39301
0 39303 7 2 2 59364 70631
0 39304 5 1 1 95889
0 39305 7 1 2 62730 72868
0 39306 5 1 1 39305
0 39307 7 1 2 88636 39306
0 39308 5 1 1 39307
0 39309 7 1 2 91779 39308
0 39310 5 1 1 39309
0 39311 7 1 2 70199 39310
0 39312 5 1 1 39311
0 39313 7 1 2 39304 39312
0 39314 7 1 2 39302 39313
0 39315 5 1 1 39314
0 39316 7 1 2 69414 39315
0 39317 5 1 1 39316
0 39318 7 1 2 59365 95884
0 39319 5 1 1 39318
0 39320 7 1 2 70257 39319
0 39321 5 1 1 39320
0 39322 7 1 2 69192 39321
0 39323 5 1 1 39322
0 39324 7 1 2 59366 95875
0 39325 5 1 1 39324
0 39326 7 1 2 93174 39325
0 39327 7 1 2 39323 39326
0 39328 5 1 1 39327
0 39329 7 1 2 76051 39328
0 39330 5 1 1 39329
0 39331 7 2 2 78402 73301
0 39332 5 1 1 95891
0 39333 7 1 2 70241 95886
0 39334 5 1 1 39333
0 39335 7 1 2 70072 92920
0 39336 5 2 1 39335
0 39337 7 1 2 67696 95893
0 39338 7 1 2 39334 39337
0 39339 5 1 1 39338
0 39340 7 1 2 39332 39339
0 39341 5 1 1 39340
0 39342 7 1 2 61098 39341
0 39343 5 1 1 39342
0 39344 7 1 2 70632 83876
0 39345 5 1 1 39344
0 39346 7 1 2 76587 95892
0 39347 5 1 1 39346
0 39348 7 1 2 39345 39347
0 39349 7 1 2 39343 39348
0 39350 7 1 2 39330 39349
0 39351 7 1 2 39317 39350
0 39352 5 1 1 39351
0 39353 7 1 2 75336 39352
0 39354 5 1 1 39353
0 39355 7 2 2 39289 39354
0 39356 5 1 1 95895
0 39357 7 1 2 71651 71883
0 39358 7 1 2 93264 39357
0 39359 5 1 1 39358
0 39360 7 1 2 95896 39359
0 39361 5 1 1 39360
0 39362 7 1 2 60570 39361
0 39363 5 1 1 39362
0 39364 7 2 2 69574 73419
0 39365 7 1 2 91474 93025
0 39366 7 1 2 95897 39365
0 39367 5 1 1 39366
0 39368 7 1 2 39363 39367
0 39369 5 1 1 39368
0 39370 7 1 2 61745 39369
0 39371 5 1 1 39370
0 39372 7 1 2 93294 95856
0 39373 5 2 1 39372
0 39374 7 1 2 82933 88832
0 39375 5 1 1 39374
0 39376 7 1 2 72953 94119
0 39377 5 1 1 39376
0 39378 7 1 2 39375 39377
0 39379 5 1 1 39378
0 39380 7 2 2 67351 39379
0 39381 7 1 2 71423 73258
0 39382 7 1 2 95901 39381
0 39383 5 1 1 39382
0 39384 7 1 2 72562 75792
0 39385 5 1 1 39384
0 39386 7 1 2 90792 91931
0 39387 7 1 2 39385 39386
0 39388 5 1 1 39387
0 39389 7 1 2 39383 39388
0 39390 7 1 2 95899 39389
0 39391 5 1 1 39390
0 39392 7 1 2 89319 39391
0 39393 5 1 1 39392
0 39394 7 1 2 65604 39393
0 39395 7 1 2 39371 39394
0 39396 5 1 1 39395
0 39397 7 1 2 39284 39396
0 39398 5 1 1 39397
0 39399 7 2 2 82869 92167
0 39400 7 1 2 74947 85303
0 39401 7 1 2 95703 39400
0 39402 7 1 2 95903 39401
0 39403 7 1 2 85765 39402
0 39404 5 1 1 39403
0 39405 7 1 2 39398 39404
0 39406 5 1 1 39405
0 39407 7 1 2 61882 39406
0 39408 5 1 1 39407
0 39409 7 3 2 66877 89320
0 39410 5 1 1 95905
0 39411 7 3 2 60684 95906
0 39412 5 1 1 95908
0 39413 7 1 2 80873 39356
0 39414 5 1 1 39413
0 39415 7 2 2 68061 74799
0 39416 5 1 1 95911
0 39417 7 1 2 88833 92685
0 39418 7 1 2 95912 39417
0 39419 5 1 1 39418
0 39420 7 1 2 81418 78603
0 39421 5 1 1 39420
0 39422 7 1 2 61369 71502
0 39423 5 1 1 39422
0 39424 7 1 2 39421 39423
0 39425 5 1 1 39424
0 39426 7 1 2 60939 39425
0 39427 5 1 1 39426
0 39428 7 1 2 75716 73644
0 39429 5 1 1 39428
0 39430 7 1 2 39427 39429
0 39431 5 1 1 39430
0 39432 7 1 2 60170 71884
0 39433 7 1 2 39431 39432
0 39434 5 1 1 39433
0 39435 7 1 2 39419 39434
0 39436 5 1 1 39435
0 39437 7 1 2 59578 39436
0 39438 5 1 1 39437
0 39439 7 1 2 72872 95902
0 39440 5 1 1 39439
0 39441 7 1 2 39438 39440
0 39442 5 1 1 39441
0 39443 7 1 2 59931 39442
0 39444 5 1 1 39443
0 39445 7 1 2 95900 39444
0 39446 7 1 2 39414 39445
0 39447 5 1 1 39446
0 39448 7 1 2 95909 39447
0 39449 5 1 1 39448
0 39450 7 1 2 39408 39449
0 39451 5 1 1 39450
0 39452 7 1 2 94209 39451
0 39453 5 1 1 39452
0 39454 7 1 2 39032 39453
0 39455 7 1 2 38318 39454
0 39456 5 1 1 39455
0 39457 7 1 2 68894 39456
0 39458 5 1 1 39457
0 39459 7 6 2 60685 94749
0 39460 7 2 2 95751 95913
0 39461 7 1 2 59367 93972
0 39462 5 1 1 39461
0 39463 7 1 2 87518 92655
0 39464 5 1 1 39463
0 39465 7 1 2 39462 39464
0 39466 5 1 1 39465
0 39467 7 1 2 69415 39466
0 39468 5 1 1 39467
0 39469 7 1 2 59368 75506
0 39470 7 1 2 92212 39469
0 39471 5 1 1 39470
0 39472 7 1 2 28369 39471
0 39473 5 1 1 39472
0 39474 7 1 2 76052 39473
0 39475 5 1 1 39474
0 39476 7 1 2 39468 39475
0 39477 5 1 1 39476
0 39478 7 1 2 68062 39477
0 39479 5 1 1 39478
0 39480 7 3 2 75621 95499
0 39481 5 3 1 95921
0 39482 7 1 2 73382 95924
0 39483 5 1 1 39482
0 39484 7 2 2 75337 70235
0 39485 7 1 2 73457 95927
0 39486 5 1 1 39485
0 39487 7 1 2 39483 39486
0 39488 5 1 1 39487
0 39489 7 1 2 68722 39488
0 39490 5 1 1 39489
0 39491 7 1 2 39479 39490
0 39492 5 1 1 39491
0 39493 7 1 2 71885 39492
0 39494 5 1 1 39493
0 39495 7 1 2 73389 74654
0 39496 5 1 1 39495
0 39497 7 1 2 59579 91795
0 39498 7 1 2 83493 39497
0 39499 5 1 1 39498
0 39500 7 1 2 39496 39499
0 39501 5 1 1 39500
0 39502 7 1 2 68723 39501
0 39503 5 1 1 39502
0 39504 7 1 2 39494 39503
0 39505 5 1 1 39504
0 39506 7 1 2 68428 39505
0 39507 5 1 1 39506
0 39508 7 1 2 70633 88949
0 39509 5 1 1 39508
0 39510 7 1 2 72677 91027
0 39511 5 2 1 39510
0 39512 7 4 2 60171 73917
0 39513 5 1 1 95931
0 39514 7 1 2 70236 88950
0 39515 5 1 1 39514
0 39516 7 1 2 39513 39515
0 39517 5 1 1 39516
0 39518 7 1 2 71503 39517
0 39519 5 1 1 39518
0 39520 7 1 2 95929 39519
0 39521 5 1 1 39520
0 39522 7 1 2 59580 39521
0 39523 5 1 1 39522
0 39524 7 1 2 39509 39523
0 39525 5 1 1 39524
0 39526 7 1 2 87953 39525
0 39527 5 1 1 39526
0 39528 7 1 2 39507 39527
0 39529 5 1 1 39528
0 39530 7 1 2 95919 39529
0 39531 5 1 1 39530
0 39532 7 2 2 92372 90172
0 39533 7 1 2 59581 95623
0 39534 5 1 1 39533
0 39535 7 1 2 18320 39534
0 39536 5 1 1 39535
0 39537 7 1 2 68429 91132
0 39538 7 1 2 39536 39537
0 39539 5 1 1 39538
0 39540 7 3 2 82269 88995
0 39541 7 1 2 68430 95937
0 39542 5 1 1 39541
0 39543 7 1 2 59582 80956
0 39544 5 1 1 39543
0 39545 7 1 2 82593 39544
0 39546 5 3 1 39545
0 39547 7 1 2 82993 95940
0 39548 5 1 1 39547
0 39549 7 1 2 39542 39548
0 39550 5 1 1 39549
0 39551 7 1 2 69416 39550
0 39552 5 1 1 39551
0 39553 7 2 2 76588 95469
0 39554 7 1 2 76053 95943
0 39555 5 1 1 39554
0 39556 7 1 2 76054 89519
0 39557 5 3 1 39556
0 39558 7 1 2 83055 85886
0 39559 5 1 1 39558
0 39560 7 1 2 95945 39559
0 39561 7 1 2 39555 39560
0 39562 5 1 1 39561
0 39563 7 1 2 59932 39562
0 39564 5 1 1 39563
0 39565 7 1 2 39552 39564
0 39566 7 1 2 39539 39565
0 39567 5 2 1 39566
0 39568 7 1 2 95935 95948
0 39569 5 1 1 39568
0 39570 7 4 2 59583 91675
0 39571 5 1 1 95950
0 39572 7 2 2 77796 84351
0 39573 5 1 1 95954
0 39574 7 1 2 95951 95955
0 39575 5 1 1 39574
0 39576 7 3 2 81990 79017
0 39577 7 1 2 95662 95956
0 39578 5 1 1 39577
0 39579 7 1 2 39575 39578
0 39580 5 1 1 39579
0 39581 7 1 2 70634 39580
0 39582 5 1 1 39581
0 39583 7 1 2 93771 95890
0 39584 5 1 1 39583
0 39585 7 1 2 95094 39584
0 39586 5 1 1 39585
0 39587 7 1 2 59584 39586
0 39588 5 1 1 39587
0 39589 7 1 2 70635 84489
0 39590 5 4 1 39589
0 39591 7 1 2 39588 95959
0 39592 5 1 1 39591
0 39593 7 1 2 61099 39592
0 39594 5 1 1 39593
0 39595 7 1 2 76500 95089
0 39596 5 1 1 39595
0 39597 7 1 2 39594 39596
0 39598 5 1 1 39597
0 39599 7 1 2 69417 39598
0 39600 5 1 1 39599
0 39601 7 2 2 76055 82499
0 39602 7 1 2 95090 95963
0 39603 5 1 1 39602
0 39604 7 1 2 39600 39603
0 39605 5 1 1 39604
0 39606 7 1 2 91676 39605
0 39607 5 1 1 39606
0 39608 7 1 2 64324 74980
0 39609 5 2 1 39608
0 39610 7 4 2 80592 85013
0 39611 5 1 1 95967
0 39612 7 2 2 84490 95968
0 39613 7 1 2 95965 95971
0 39614 5 1 1 39613
0 39615 7 1 2 82588 93772
0 39616 5 1 1 39615
0 39617 7 6 2 68724 85681
0 39618 7 1 2 90057 95973
0 39619 5 1 1 39618
0 39620 7 3 2 59369 84491
0 39621 5 1 1 95979
0 39622 7 1 2 68431 95980
0 39623 5 1 1 39622
0 39624 7 1 2 39619 39623
0 39625 5 1 1 39624
0 39626 7 1 2 70285 39625
0 39627 5 1 1 39626
0 39628 7 1 2 39616 39627
0 39629 7 1 2 39614 39628
0 39630 5 1 1 39629
0 39631 7 1 2 91677 39630
0 39632 5 1 1 39631
0 39633 7 1 2 79758 39611
0 39634 5 1 1 39633
0 39635 7 1 2 39634 95966
0 39636 5 1 1 39635
0 39637 7 1 2 74442 39636
0 39638 5 1 1 39637
0 39639 7 1 2 92094 39638
0 39640 5 1 1 39639
0 39641 7 2 2 75507 92156
0 39642 5 3 1 95982
0 39643 7 1 2 75889 83718
0 39644 5 4 1 39643
0 39645 7 2 2 90196 92900
0 39646 7 1 2 95987 95991
0 39647 5 1 1 39646
0 39648 7 1 2 95984 39647
0 39649 5 1 1 39648
0 39650 7 1 2 59585 39649
0 39651 5 1 1 39650
0 39652 7 1 2 70636 84620
0 39653 7 1 2 95992 39652
0 39654 5 1 1 39653
0 39655 7 1 2 39651 39654
0 39656 5 1 1 39655
0 39657 7 1 2 69418 39656
0 39658 5 1 1 39657
0 39659 7 2 2 61746 83552
0 39660 7 1 2 73302 95993
0 39661 7 1 2 95795 39660
0 39662 5 1 1 39661
0 39663 7 1 2 39658 39662
0 39664 7 1 2 39640 39663
0 39665 7 1 2 39632 39664
0 39666 5 1 1 39665
0 39667 7 1 2 61100 39666
0 39668 5 1 1 39667
0 39669 7 1 2 95964 95983
0 39670 5 1 1 39669
0 39671 7 1 2 60571 69419
0 39672 7 1 2 91946 39671
0 39673 7 1 2 92719 39672
0 39674 5 1 1 39673
0 39675 7 1 2 39670 39674
0 39676 7 1 2 39668 39675
0 39677 7 1 2 39607 39676
0 39678 5 1 1 39677
0 39679 7 1 2 68063 39678
0 39680 5 1 1 39679
0 39681 7 1 2 39582 39680
0 39682 5 1 1 39681
0 39683 7 1 2 67697 39682
0 39684 5 1 1 39683
0 39685 7 3 2 59586 70637
0 39686 7 2 2 60810 78131
0 39687 7 1 2 82500 95998
0 39688 5 1 1 39687
0 39689 7 1 2 63526 39688
0 39690 5 2 1 39689
0 39691 7 1 2 95995 96000
0 39692 5 1 1 39691
0 39693 7 1 2 66733 39692
0 39694 5 1 1 39693
0 39695 7 1 2 92095 39694
0 39696 5 1 1 39695
0 39697 7 2 2 59587 96001
0 39698 5 1 1 96002
0 39699 7 1 2 84492 91982
0 39700 7 1 2 96003 39699
0 39701 5 1 1 39700
0 39702 7 1 2 39696 39701
0 39703 7 1 2 39684 39702
0 39704 5 1 1 39703
0 39705 7 1 2 68895 39704
0 39706 5 1 1 39705
0 39707 7 1 2 39569 39706
0 39708 5 2 1 39707
0 39709 7 1 2 61883 96004
0 39710 5 1 1 39709
0 39711 7 1 2 70833 88732
0 39712 5 3 1 39711
0 39713 7 1 2 68432 96006
0 39714 5 1 1 39713
0 39715 7 4 2 69939 91495
0 39716 5 1 1 96009
0 39717 7 1 2 91512 96010
0 39718 5 1 1 39717
0 39719 7 1 2 39714 39718
0 39720 5 1 1 39719
0 39721 7 1 2 59588 39720
0 39722 5 1 1 39721
0 39723 7 2 2 72954 92380
0 39724 5 1 1 96013
0 39725 7 1 2 39722 39724
0 39726 5 1 1 39725
0 39727 7 9 2 86235 89339
0 39728 5 3 1 96015
0 39729 7 2 2 86343 96016
0 39730 7 1 2 67698 96027
0 39731 7 1 2 39726 39730
0 39732 5 1 1 39731
0 39733 7 1 2 65605 39732
0 39734 7 1 2 39710 39733
0 39735 5 1 1 39734
0 39736 7 1 2 66878 96005
0 39737 5 1 1 39736
0 39738 7 1 2 59933 85014
0 39739 5 2 1 39738
0 39740 7 1 2 79759 74443
0 39741 5 1 1 39740
0 39742 7 1 2 59589 39741
0 39743 5 1 1 39742
0 39744 7 1 2 96029 39743
0 39745 5 1 1 39744
0 39746 7 1 2 61101 39745
0 39747 5 1 1 39746
0 39748 7 1 2 70638 83992
0 39749 5 1 1 39748
0 39750 7 1 2 83759 39749
0 39751 5 1 1 39750
0 39752 7 1 2 59590 39751
0 39753 5 1 1 39752
0 39754 7 1 2 39747 39753
0 39755 5 1 1 39754
0 39756 7 3 2 64020 89302
0 39757 7 1 2 39755 96031
0 39758 5 1 1 39757
0 39759 7 2 2 84266 91150
0 39760 7 2 2 68896 88520
0 39761 7 1 2 96034 96036
0 39762 5 1 1 39761
0 39763 7 1 2 39758 39762
0 39764 5 1 1 39763
0 39765 7 1 2 67699 39764
0 39766 5 1 1 39765
0 39767 7 1 2 70639 76056
0 39768 7 1 2 72412 39767
0 39769 5 1 1 39768
0 39770 7 1 2 91467 95941
0 39771 5 1 1 39770
0 39772 7 1 2 95946 39771
0 39773 7 1 2 39769 39772
0 39774 5 1 1 39773
0 39775 7 1 2 96032 39774
0 39776 5 1 1 39775
0 39777 7 1 2 71931 92921
0 39778 5 1 1 39777
0 39779 7 1 2 81001 87475
0 39780 7 1 2 39778 39779
0 39781 5 1 1 39780
0 39782 7 1 2 39776 39781
0 39783 5 1 1 39782
0 39784 7 1 2 59370 39783
0 39785 5 1 1 39784
0 39786 7 2 2 90954 95599
0 39787 7 1 2 59591 96038
0 39788 5 1 1 39787
0 39789 7 1 2 83068 88917
0 39790 5 1 1 39789
0 39791 7 1 2 60811 39790
0 39792 5 1 1 39791
0 39793 7 1 2 84611 39792
0 39794 7 1 2 39788 39793
0 39795 5 1 1 39794
0 39796 7 1 2 70640 96033
0 39797 7 1 2 39795 39796
0 39798 5 1 1 39797
0 39799 7 1 2 39785 39798
0 39800 7 1 2 39766 39799
0 39801 5 1 1 39800
0 39802 7 1 2 63791 39801
0 39803 5 1 1 39802
0 39804 7 1 2 80173 95949
0 39805 5 1 1 39804
0 39806 7 2 2 79265 77915
0 39807 5 1 1 96040
0 39808 7 1 2 94975 96041
0 39809 5 1 1 39808
0 39810 7 1 2 39805 39809
0 39811 5 1 1 39810
0 39812 7 1 2 77572 39811
0 39813 5 1 1 39812
0 39814 7 2 2 83886 77573
0 39815 7 1 2 74973 72235
0 39816 7 1 2 96042 39815
0 39817 5 1 1 39816
0 39818 7 1 2 93853 39817
0 39819 5 1 1 39818
0 39820 7 1 2 79796 39819
0 39821 5 1 1 39820
0 39822 7 3 2 66562 87925
0 39823 5 1 1 96044
0 39824 7 1 2 86473 96045
0 39825 5 1 1 39824
0 39826 7 1 2 39821 39825
0 39827 5 1 1 39826
0 39828 7 1 2 63115 39827
0 39829 5 1 1 39828
0 39830 7 1 2 39813 39829
0 39831 7 1 2 39803 39830
0 39832 5 1 1 39831
0 39833 7 1 2 60385 39832
0 39834 5 1 1 39833
0 39835 7 2 2 82777 72149
0 39836 5 1 1 96047
0 39837 7 1 2 82493 96048
0 39838 5 1 1 39837
0 39839 7 1 2 92014 39838
0 39840 5 1 1 39839
0 39841 7 1 2 91770 39840
0 39842 5 1 1 39841
0 39843 7 1 2 68433 39842
0 39844 5 1 1 39843
0 39845 7 2 2 59934 84352
0 39846 5 4 1 96049
0 39847 7 1 2 39621 96051
0 39848 5 2 1 39847
0 39849 7 1 2 92004 96055
0 39850 5 1 1 39849
0 39851 7 1 2 39844 39850
0 39852 5 1 1 39851
0 39853 7 1 2 64021 39852
0 39854 5 1 1 39853
0 39855 7 2 2 72413 86529
0 39856 7 1 2 92833 96057
0 39857 5 1 1 39856
0 39858 7 1 2 39854 39857
0 39859 5 1 1 39858
0 39860 7 1 2 59592 39859
0 39861 5 1 1 39860
0 39862 7 1 2 95663 96058
0 39863 5 1 1 39862
0 39864 7 2 2 59371 95942
0 39865 5 1 1 96059
0 39866 7 1 2 93231 96060
0 39867 5 1 1 39866
0 39868 7 1 2 39863 39867
0 39869 5 1 1 39868
0 39870 7 1 2 66734 39869
0 39871 5 1 1 39870
0 39872 7 1 2 80038 70641
0 39873 5 2 1 39872
0 39874 7 1 2 83719 96061
0 39875 5 7 1 39874
0 39876 7 3 2 86590 92271
0 39877 5 1 1 96070
0 39878 7 2 2 67700 96071
0 39879 5 1 1 96073
0 39880 7 1 2 82501 92373
0 39881 5 1 1 39880
0 39882 7 1 2 39879 39881
0 39883 5 1 1 39882
0 39884 7 1 2 96063 39883
0 39885 5 1 1 39884
0 39886 7 2 2 70642 85140
0 39887 5 1 1 96075
0 39888 7 2 2 67701 89934
0 39889 7 1 2 92635 96077
0 39890 5 1 1 39889
0 39891 7 1 2 39887 39890
0 39892 5 1 1 39891
0 39893 7 5 2 59593 61747
0 39894 7 1 2 64022 96079
0 39895 7 1 2 39892 39894
0 39896 5 1 1 39895
0 39897 7 1 2 39885 39896
0 39898 7 1 2 39871 39897
0 39899 5 1 1 39898
0 39900 7 1 2 69420 39899
0 39901 5 1 1 39900
0 39902 7 2 2 59935 89638
0 39903 7 1 2 77574 85304
0 39904 7 1 2 96084 39903
0 39905 5 1 1 39904
0 39906 7 1 2 82270 92425
0 39907 5 1 1 39906
0 39908 7 1 2 70643 87917
0 39909 5 1 1 39908
0 39910 7 1 2 39907 39909
0 39911 5 1 1 39910
0 39912 7 1 2 59372 63792
0 39913 7 1 2 39911 39912
0 39914 5 1 1 39913
0 39915 7 1 2 39905 39914
0 39916 5 1 1 39915
0 39917 7 1 2 70286 39916
0 39918 5 1 1 39917
0 39919 7 1 2 70460 96074
0 39920 5 1 1 39919
0 39921 7 4 2 60812 61748
0 39922 7 1 2 59936 96086
0 39923 7 1 2 92193 39922
0 39924 5 1 1 39923
0 39925 7 1 2 39920 39924
0 39926 5 1 1 39925
0 39927 7 1 2 96064 39926
0 39928 5 1 1 39927
0 39929 7 1 2 76501 96065
0 39930 5 1 1 39929
0 39931 7 1 2 8814 39930
0 39932 5 1 1 39931
0 39933 7 4 2 67092 85524
0 39934 7 1 2 80775 96090
0 39935 5 1 1 39934
0 39936 7 1 2 92378 39935
0 39937 5 1 1 39936
0 39938 7 1 2 39932 39937
0 39939 5 1 1 39938
0 39940 7 1 2 71886 89749
0 39941 5 1 1 39940
0 39942 7 3 2 61370 84493
0 39943 7 1 2 73420 96094
0 39944 5 1 1 39943
0 39945 7 1 2 39941 39944
0 39946 5 1 1 39945
0 39947 7 1 2 79142 39946
0 39948 5 1 1 39947
0 39949 7 1 2 68064 39948
0 39950 7 1 2 39939 39949
0 39951 7 1 2 39928 39950
0 39952 7 1 2 39918 39951
0 39953 7 1 2 39901 39952
0 39954 7 1 2 39861 39953
0 39955 5 1 1 39954
0 39956 7 2 2 81991 74933
0 39957 5 1 1 96097
0 39958 7 1 2 88647 94404
0 39959 7 1 2 83887 39958
0 39960 5 1 1 39959
0 39961 7 1 2 39957 39960
0 39962 5 1 1 39961
0 39963 7 1 2 70644 77575
0 39964 7 1 2 39962 39963
0 39965 5 1 1 39964
0 39966 7 1 2 90611 93850
0 39967 5 1 1 39966
0 39968 7 1 2 63116 39967
0 39969 7 1 2 39965 39968
0 39970 5 1 1 39969
0 39971 7 1 2 39955 39970
0 39972 5 1 1 39971
0 39973 7 1 2 67702 95996
0 39974 5 1 1 39973
0 39975 7 1 2 39865 39974
0 39976 5 1 1 39975
0 39977 7 1 2 84494 39976
0 39978 5 1 1 39977
0 39979 7 1 2 59937 84614
0 39980 7 1 2 96078 39979
0 39981 5 1 1 39980
0 39982 7 1 2 39978 39981
0 39983 5 1 1 39982
0 39984 7 1 2 61102 39983
0 39985 5 1 1 39984
0 39986 7 2 2 83343 84495
0 39987 5 1 1 96099
0 39988 7 1 2 92213 96100
0 39989 5 1 1 39988
0 39990 7 1 2 39985 39989
0 39991 5 1 1 39990
0 39992 7 1 2 69421 39991
0 39993 5 1 1 39992
0 39994 7 1 2 82485 72955
0 39995 7 1 2 96095 39994
0 39996 5 1 1 39995
0 39997 7 2 2 84267 89935
0 39998 5 2 1 96101
0 39999 7 1 2 96103 95960
0 40000 5 1 1 39999
0 40001 7 1 2 59373 82271
0 40002 7 1 2 40000 40001
0 40003 5 1 1 40002
0 40004 7 1 2 39996 40003
0 40005 5 1 1 40004
0 40006 7 1 2 76057 40005
0 40007 5 1 1 40006
0 40008 7 1 2 37853 96030
0 40009 5 1 1 40008
0 40010 7 1 2 71887 84496
0 40011 7 1 2 40009 40010
0 40012 5 1 1 40011
0 40013 7 1 2 84353 86300
0 40014 5 2 1 40013
0 40015 7 1 2 40012 96105
0 40016 7 1 2 40007 40015
0 40017 7 1 2 39993 40016
0 40018 5 1 1 40017
0 40019 7 1 2 79143 40018
0 40020 5 1 1 40019
0 40021 7 3 2 59594 85525
0 40022 5 1 1 96107
0 40023 7 1 2 65475 93768
0 40024 7 1 2 96108 40023
0 40025 5 1 1 40024
0 40026 7 1 2 40020 40025
0 40027 7 1 2 39972 40026
0 40028 7 1 2 39834 40027
0 40029 5 1 1 40028
0 40030 7 1 2 61884 40029
0 40031 5 1 1 40030
0 40032 7 1 2 83105 88648
0 40033 7 1 2 90135 40032
0 40034 7 2 2 96043 40033
0 40035 5 1 1 96110
0 40036 7 1 2 60686 40035
0 40037 7 1 2 40031 40036
0 40038 7 1 2 39737 40037
0 40039 5 1 1 40038
0 40040 7 1 2 39735 40039
0 40041 5 1 1 40040
0 40042 7 1 2 73193 95054
0 40043 5 1 1 40042
0 40044 7 1 2 9708 40043
0 40045 5 1 1 40044
0 40046 7 1 2 59595 40045
0 40047 5 1 1 40046
0 40048 7 1 2 68725 71324
0 40049 5 1 1 40048
0 40050 7 1 2 86103 93792
0 40051 7 1 2 40049 40050
0 40052 5 1 1 40051
0 40053 7 1 2 40047 40052
0 40054 5 1 1 40053
0 40055 7 1 2 68065 40054
0 40056 5 1 1 40055
0 40057 7 1 2 87667 89750
0 40058 7 1 2 96037 40057
0 40059 5 1 1 40058
0 40060 7 1 2 40056 40059
0 40061 5 1 1 40060
0 40062 7 1 2 59938 40061
0 40063 5 1 1 40062
0 40064 7 2 2 86142 94346
0 40065 5 1 1 96112
0 40066 7 1 2 59596 87277
0 40067 5 1 1 40066
0 40068 7 1 2 40065 40067
0 40069 5 1 1 40068
0 40070 7 1 2 69940 40069
0 40071 5 1 1 40070
0 40072 7 3 2 66879 80981
0 40073 5 2 1 96114
0 40074 7 1 2 76262 96115
0 40075 5 1 1 40074
0 40076 7 1 2 40071 40075
0 40077 5 1 1 40076
0 40078 7 1 2 84497 40077
0 40079 5 1 1 40078
0 40080 7 1 2 9710 40079
0 40081 7 1 2 40063 40080
0 40082 5 1 1 40081
0 40083 7 1 2 71888 40082
0 40084 5 1 1 40083
0 40085 7 1 2 69422 96056
0 40086 5 1 1 40085
0 40087 7 1 2 82502 84354
0 40088 5 1 1 40087
0 40089 7 1 2 40086 40088
0 40090 5 1 1 40089
0 40091 7 1 2 59597 40090
0 40092 5 1 1 40091
0 40093 7 1 2 84355 91796
0 40094 5 1 1 40093
0 40095 7 1 2 40092 40094
0 40096 5 1 1 40095
0 40097 7 1 2 86330 40096
0 40098 5 1 1 40097
0 40099 7 1 2 40084 40098
0 40100 5 1 1 40099
0 40101 7 1 2 91678 40100
0 40102 5 1 1 40101
0 40103 7 5 2 75508 87213
0 40104 5 4 1 96119
0 40105 7 1 2 69575 96120
0 40106 5 1 1 40105
0 40107 7 1 2 85864 96124
0 40108 5 2 1 40107
0 40109 7 1 2 84021 96128
0 40110 5 1 1 40109
0 40111 7 1 2 40106 40110
0 40112 5 1 1 40111
0 40113 7 1 2 68434 40112
0 40114 5 1 1 40113
0 40115 7 1 2 85690 96125
0 40116 5 1 1 40115
0 40117 7 1 2 91463 94121
0 40118 7 1 2 40116 40117
0 40119 5 1 1 40118
0 40120 7 1 2 40114 40119
0 40121 5 1 1 40120
0 40122 7 1 2 63793 40121
0 40123 5 1 1 40122
0 40124 7 3 2 63527 95988
0 40125 7 2 2 92680 96130
0 40126 5 1 1 96133
0 40127 7 1 2 92333 96134
0 40128 5 1 1 40127
0 40129 7 1 2 40123 40128
0 40130 5 1 1 40129
0 40131 7 1 2 71889 40130
0 40132 5 1 1 40131
0 40133 7 2 2 82782 95989
0 40134 7 1 2 92780 96135
0 40135 5 1 1 40134
0 40136 7 1 2 75882 92799
0 40137 5 1 1 40136
0 40138 7 1 2 40135 40137
0 40139 5 1 1 40138
0 40140 7 1 2 63528 40139
0 40141 5 1 1 40140
0 40142 7 1 2 83706 92800
0 40143 5 1 1 40142
0 40144 7 1 2 40141 40143
0 40145 5 1 1 40144
0 40146 7 1 2 82994 40145
0 40147 5 1 1 40146
0 40148 7 3 2 81992 85704
0 40149 7 2 2 83783 71890
0 40150 5 1 1 96140
0 40151 7 1 2 96137 96141
0 40152 5 1 1 40151
0 40153 7 1 2 61885 80174
0 40154 7 1 2 84439 40153
0 40155 5 1 1 40154
0 40156 7 1 2 40152 40155
0 40157 5 1 1 40156
0 40158 7 1 2 65476 40157
0 40159 5 1 1 40158
0 40160 7 2 2 82415 92272
0 40161 7 3 2 61886 96142
0 40162 5 1 1 96144
0 40163 7 1 2 83409 96145
0 40164 5 1 1 40163
0 40165 7 1 2 40159 40164
0 40166 5 1 1 40165
0 40167 7 1 2 88521 40166
0 40168 5 1 1 40167
0 40169 7 1 2 40147 40168
0 40170 7 1 2 40132 40169
0 40171 5 1 1 40170
0 40172 7 1 2 68897 40171
0 40173 5 1 1 40172
0 40174 7 1 2 92120 93929
0 40175 5 1 1 40174
0 40176 7 1 2 63117 91679
0 40177 7 1 2 91776 93905
0 40178 7 1 2 40176 40177
0 40179 5 1 1 40178
0 40180 7 1 2 40175 40179
0 40181 5 1 1 40180
0 40182 7 1 2 68435 40181
0 40183 5 1 1 40182
0 40184 7 1 2 77797 91777
0 40185 5 1 1 40184
0 40186 7 1 2 78981 40185
0 40187 5 1 1 40186
0 40188 7 1 2 85705 88130
0 40189 7 1 2 40187 40188
0 40190 5 1 1 40189
0 40191 7 1 2 84870 87343
0 40192 5 1 1 40191
0 40193 7 1 2 86104 89975
0 40194 5 1 1 40193
0 40195 7 1 2 40192 40194
0 40196 5 1 1 40195
0 40197 7 1 2 60386 40196
0 40198 5 2 1 40197
0 40199 7 1 2 86373 90142
0 40200 5 1 1 40199
0 40201 7 1 2 96147 40200
0 40202 7 1 2 40190 40201
0 40203 5 1 1 40202
0 40204 7 1 2 61749 40203
0 40205 5 1 1 40204
0 40206 7 1 2 40183 40205
0 40207 5 1 1 40206
0 40208 7 1 2 73303 40207
0 40209 5 1 1 40208
0 40210 7 1 2 60687 40209
0 40211 7 1 2 40173 40210
0 40212 7 1 2 6714 95246
0 40213 5 1 1 40212
0 40214 7 1 2 96121 40213
0 40215 5 1 1 40214
0 40216 7 1 2 61887 74867
0 40217 7 1 2 86659 40216
0 40218 5 1 1 40217
0 40219 7 1 2 40215 40218
0 40220 5 1 1 40219
0 40221 7 1 2 76058 40220
0 40222 5 1 1 40221
0 40223 7 2 2 81541 78436
0 40224 5 1 1 96149
0 40225 7 1 2 85673 96150
0 40226 5 1 1 40225
0 40227 7 1 2 40222 40226
0 40228 5 1 1 40227
0 40229 7 1 2 59939 40228
0 40230 5 1 1 40229
0 40231 7 1 2 88951 96122
0 40232 5 1 1 40231
0 40233 7 1 2 68066 86063
0 40234 5 1 1 40233
0 40235 7 1 2 40232 40234
0 40236 5 1 1 40235
0 40237 7 1 2 68436 40236
0 40238 5 1 1 40237
0 40239 7 1 2 40230 40238
0 40240 5 1 1 40239
0 40241 7 1 2 90197 40240
0 40242 5 1 1 40241
0 40243 7 3 2 59598 61888
0 40244 7 1 2 78776 96151
0 40245 5 1 1 40244
0 40246 7 3 2 59940 84285
0 40247 7 1 2 78263 85706
0 40248 7 1 2 96154 40247
0 40249 5 1 1 40248
0 40250 7 1 2 40245 40249
0 40251 5 1 1 40250
0 40252 7 1 2 59374 40251
0 40253 5 1 1 40252
0 40254 7 2 2 89999 94347
0 40255 7 1 2 96080 96157
0 40256 5 1 1 40255
0 40257 7 1 2 40253 40256
0 40258 5 1 1 40257
0 40259 7 1 2 90173 40258
0 40260 5 1 1 40259
0 40261 7 3 2 77916 90198
0 40262 5 1 1 96159
0 40263 7 2 2 66563 96160
0 40264 5 1 1 96162
0 40265 7 1 2 86356 95182
0 40266 7 1 2 96163 40265
0 40267 5 1 1 40266
0 40268 7 1 2 40260 40267
0 40269 5 1 1 40268
0 40270 7 1 2 69423 40269
0 40271 5 1 1 40270
0 40272 7 2 2 84804 85141
0 40273 5 1 1 96164
0 40274 7 3 2 75509 96165
0 40275 7 1 2 86357 92681
0 40276 7 1 2 96166 40275
0 40277 5 1 1 40276
0 40278 7 1 2 40271 40277
0 40279 7 1 2 40242 40278
0 40280 5 1 1 40279
0 40281 7 1 2 64023 40280
0 40282 5 1 1 40281
0 40283 7 3 2 79653 79712
0 40284 5 1 1 96169
0 40285 7 1 2 85857 86988
0 40286 5 7 1 40285
0 40287 7 1 2 68726 76422
0 40288 7 1 2 96172 40287
0 40289 5 1 1 40288
0 40290 7 1 2 40284 40289
0 40291 5 1 1 40290
0 40292 7 1 2 69424 40291
0 40293 5 1 1 40292
0 40294 7 1 2 70461 91821
0 40295 5 1 1 40294
0 40296 7 4 2 66735 86433
0 40297 7 1 2 73437 96179
0 40298 5 1 1 40297
0 40299 7 1 2 40295 40298
0 40300 5 1 1 40299
0 40301 7 1 2 61889 40300
0 40302 5 1 1 40301
0 40303 7 2 2 85707 89811
0 40304 7 1 2 59599 93039
0 40305 7 1 2 96183 40304
0 40306 5 1 1 40305
0 40307 7 1 2 40302 40306
0 40308 7 1 2 40293 40307
0 40309 5 1 1 40308
0 40310 7 1 2 95484 40309
0 40311 5 1 1 40310
0 40312 7 7 2 61890 79654
0 40313 5 1 1 96185
0 40314 7 1 2 70987 89687
0 40315 7 1 2 96186 40314
0 40316 5 1 1 40315
0 40317 7 1 2 40311 40316
0 40318 5 1 1 40317
0 40319 7 1 2 59941 40318
0 40320 5 1 1 40319
0 40321 7 1 2 86540 91545
0 40322 7 1 2 96170 40321
0 40323 5 1 1 40322
0 40324 7 1 2 64024 40323
0 40325 7 1 2 40320 40324
0 40326 5 1 1 40325
0 40327 7 1 2 63118 18997
0 40328 5 1 1 40327
0 40329 7 1 2 84498 40328
0 40330 5 1 1 40329
0 40331 7 1 2 59600 89030
0 40332 7 1 2 93773 40331
0 40333 5 1 1 40332
0 40334 7 1 2 40330 40333
0 40335 5 1 1 40334
0 40336 7 1 2 69941 40335
0 40337 5 1 1 40336
0 40338 7 2 2 61750 84440
0 40339 5 4 1 96192
0 40340 7 1 2 19935 21525
0 40341 5 1 1 40340
0 40342 7 1 2 69576 15520
0 40343 7 1 2 40341 40342
0 40344 5 1 1 40343
0 40345 7 1 2 96194 40344
0 40346 5 1 1 40345
0 40347 7 1 2 59601 40346
0 40348 5 1 1 40347
0 40349 7 1 2 93774 95879
0 40350 5 1 1 40349
0 40351 7 1 2 27318 40350
0 40352 7 1 2 40348 40351
0 40353 7 1 2 40337 40352
0 40354 5 1 1 40353
0 40355 7 1 2 87214 40354
0 40356 5 1 1 40355
0 40357 7 3 2 79048 85848
0 40358 7 1 2 94016 96198
0 40359 5 1 1 40358
0 40360 7 1 2 68898 40359
0 40361 7 1 2 40356 40360
0 40362 5 1 1 40361
0 40363 7 1 2 75338 40362
0 40364 7 1 2 40326 40363
0 40365 5 1 1 40364
0 40366 7 1 2 40282 40365
0 40367 7 1 2 40211 40366
0 40368 7 1 2 40102 40367
0 40369 5 1 1 40368
0 40370 7 1 2 86211 96136
0 40371 5 1 1 40370
0 40372 7 1 2 69045 86240
0 40373 7 1 2 92750 40372
0 40374 5 1 1 40373
0 40375 7 1 2 40371 40374
0 40376 5 1 1 40375
0 40377 7 1 2 59375 40376
0 40378 5 1 1 40377
0 40379 7 4 2 75510 92751
0 40380 7 1 2 77244 94348
0 40381 7 1 2 96201 40380
0 40382 5 1 1 40381
0 40383 7 1 2 40378 40382
0 40384 5 1 1 40383
0 40385 7 1 2 68067 40384
0 40386 5 1 1 40385
0 40387 7 1 2 30394 96126
0 40388 5 1 1 40387
0 40389 7 1 2 95944 40388
0 40390 5 1 1 40389
0 40391 7 1 2 87288 96131
0 40392 5 1 1 40391
0 40393 7 1 2 40390 40392
0 40394 5 1 1 40393
0 40395 7 1 2 73304 40394
0 40396 5 1 1 40395
0 40397 7 3 2 68437 88188
0 40398 7 1 2 73273 96205
0 40399 5 1 1 40398
0 40400 7 1 2 40126 40399
0 40401 5 1 1 40400
0 40402 7 1 2 61891 40401
0 40403 5 1 1 40402
0 40404 7 1 2 68438 96123
0 40405 7 1 2 73274 40404
0 40406 5 1 1 40405
0 40407 7 1 2 40403 40406
0 40408 5 1 1 40407
0 40409 7 1 2 71891 40408
0 40410 5 1 1 40409
0 40411 7 1 2 40396 40410
0 40412 7 1 2 40386 40411
0 40413 5 1 1 40412
0 40414 7 1 2 68899 40413
0 40415 5 1 1 40414
0 40416 7 2 2 68439 88952
0 40417 5 1 1 96208
0 40418 7 1 2 75126 95247
0 40419 5 2 1 40418
0 40420 7 1 2 76263 96210
0 40421 5 1 1 40420
0 40422 7 1 2 78132 71892
0 40423 5 3 1 40422
0 40424 7 1 2 83202 96212
0 40425 5 1 1 40424
0 40426 7 1 2 69942 40425
0 40427 5 1 1 40426
0 40428 7 1 2 40421 40427
0 40429 5 1 1 40428
0 40430 7 1 2 59942 40429
0 40431 5 1 1 40430
0 40432 7 1 2 40417 40431
0 40433 5 1 1 40432
0 40434 7 1 2 86105 92121
0 40435 7 1 2 40433 40434
0 40436 5 1 1 40435
0 40437 7 1 2 40415 40436
0 40438 5 1 1 40437
0 40439 7 1 2 68727 40438
0 40440 5 1 1 40439
0 40441 7 2 2 68440 71504
0 40442 5 1 1 96215
0 40443 7 1 2 40442 39698
0 40444 5 1 1 40443
0 40445 7 4 2 61892 68900
0 40446 7 1 2 78159 96217
0 40447 7 1 2 91742 40446
0 40448 7 1 2 40444 40447
0 40449 5 1 1 40448
0 40450 7 1 2 40440 40449
0 40451 5 1 1 40450
0 40452 7 1 2 61751 40451
0 40453 5 1 1 40452
0 40454 7 1 2 60572 92733
0 40455 5 1 1 40454
0 40456 7 1 2 39573 40455
0 40457 5 1 1 40456
0 40458 7 1 2 75016 40457
0 40459 5 1 1 40458
0 40460 7 1 2 20526 40459
0 40461 5 1 1 40460
0 40462 7 1 2 60813 40461
0 40463 5 1 1 40462
0 40464 7 2 2 84167 79018
0 40465 5 2 1 96221
0 40466 7 1 2 92236 96223
0 40467 5 1 1 40466
0 40468 7 1 2 68441 40467
0 40469 5 1 1 40468
0 40470 7 1 2 40463 40469
0 40471 5 1 1 40470
0 40472 7 1 2 59376 40471
0 40473 5 1 1 40472
0 40474 7 1 2 69425 96222
0 40475 5 1 1 40474
0 40476 7 1 2 76040 40475
0 40477 5 1 1 40476
0 40478 7 1 2 85148 96224
0 40479 5 1 1 40478
0 40480 7 1 2 68442 40479
0 40481 7 1 2 40477 40480
0 40482 5 1 1 40481
0 40483 7 1 2 40473 40482
0 40484 5 1 1 40483
0 40485 7 1 2 75511 40484
0 40486 5 1 1 40485
0 40487 7 1 2 84356 94874
0 40488 7 1 2 73314 40487
0 40489 5 1 1 40488
0 40490 7 1 2 40486 40489
0 40491 5 1 1 40490
0 40492 7 1 2 71893 96218
0 40493 7 1 2 40491 40492
0 40494 5 1 1 40493
0 40495 7 1 2 65606 40494
0 40496 7 1 2 40453 40495
0 40497 5 1 1 40496
0 40498 7 1 2 40369 40497
0 40499 5 1 1 40498
0 40500 7 1 2 92653 92849
0 40501 5 1 1 40500
0 40502 7 1 2 74124 79019
0 40503 7 1 2 94948 40502
0 40504 7 1 2 95555 40503
0 40505 5 1 1 40504
0 40506 7 1 2 40501 40505
0 40507 5 1 1 40506
0 40508 7 1 2 61893 40507
0 40509 5 1 1 40508
0 40510 7 2 2 73383 92854
0 40511 7 1 2 85345 86136
0 40512 7 1 2 96225 40511
0 40513 5 1 1 40512
0 40514 7 1 2 40509 40513
0 40515 5 1 1 40514
0 40516 7 1 2 68443 40515
0 40517 5 1 1 40516
0 40518 7 1 2 79655 92194
0 40519 5 1 1 40518
0 40520 7 1 2 84615 85191
0 40521 7 1 2 92693 40520
0 40522 5 1 1 40521
0 40523 7 1 2 40519 40522
0 40524 5 1 1 40523
0 40525 7 1 2 86212 90035
0 40526 7 1 2 40524 40525
0 40527 5 1 1 40526
0 40528 7 1 2 40517 40527
0 40529 5 1 1 40528
0 40530 7 1 2 60688 40529
0 40531 5 1 1 40530
0 40532 7 1 2 86257 96226
0 40533 5 1 1 40532
0 40534 7 1 2 87215 89841
0 40535 5 1 1 40534
0 40536 7 1 2 40533 40535
0 40537 5 1 1 40536
0 40538 7 1 2 92294 40537
0 40539 5 1 1 40538
0 40540 7 1 2 40531 40539
0 40541 5 1 1 40540
0 40542 7 1 2 71235 40541
0 40543 5 1 1 40542
0 40544 7 2 2 84357 87476
0 40545 5 1 1 96227
0 40546 7 1 2 90112 93177
0 40547 5 1 1 40546
0 40548 7 1 2 85543 40547
0 40549 5 1 1 40548
0 40550 7 1 2 92540 40549
0 40551 5 1 1 40550
0 40552 7 1 2 40545 40551
0 40553 5 1 1 40552
0 40554 7 1 2 76423 40553
0 40555 5 1 1 40554
0 40556 7 4 2 68068 85526
0 40557 5 1 1 96229
0 40558 7 1 2 61752 96230
0 40559 5 1 1 40558
0 40560 7 1 2 40555 40559
0 40561 5 1 1 40560
0 40562 7 1 2 69426 40561
0 40563 5 1 1 40562
0 40564 7 2 2 71894 95974
0 40565 5 1 1 96233
0 40566 7 1 2 59602 96234
0 40567 5 1 1 40566
0 40568 7 1 2 96195 40567
0 40569 5 1 1 40568
0 40570 7 1 2 59377 40569
0 40571 5 1 1 40570
0 40572 7 5 2 59603 84499
0 40573 7 1 2 59943 70287
0 40574 5 1 1 40573
0 40575 7 1 2 63119 40574
0 40576 5 1 1 40575
0 40577 7 1 2 96235 40576
0 40578 5 1 1 40577
0 40579 7 1 2 73438 89031
0 40580 5 1 1 40579
0 40581 7 1 2 95881 40580
0 40582 5 1 1 40581
0 40583 7 1 2 95975 40582
0 40584 5 1 1 40583
0 40585 7 1 2 40578 40584
0 40586 7 1 2 40571 40585
0 40587 5 1 1 40586
0 40588 7 1 2 68901 40587
0 40589 5 1 1 40588
0 40590 7 1 2 88015 93446
0 40591 7 1 2 86481 40590
0 40592 5 1 1 40591
0 40593 7 1 2 40589 40592
0 40594 7 1 2 40563 40593
0 40595 5 1 1 40594
0 40596 7 8 2 60573 61894
0 40597 5 1 1 96240
0 40598 7 3 2 65607 75339
0 40599 7 1 2 96241 96248
0 40600 7 1 2 40595 40599
0 40601 5 1 1 40600
0 40602 7 1 2 40543 40601
0 40603 7 1 2 40499 40602
0 40604 5 1 1 40603
0 40605 7 1 2 70200 40604
0 40606 5 1 1 40605
0 40607 7 2 2 92005 92374
0 40608 7 3 2 59944 73259
0 40609 5 1 1 96253
0 40610 7 1 2 63120 40609
0 40611 5 1 1 40610
0 40612 7 1 2 61103 40611
0 40613 5 1 1 40612
0 40614 7 2 2 71505 83056
0 40615 5 1 1 96256
0 40616 7 1 2 40613 40615
0 40617 5 1 1 40616
0 40618 7 1 2 67703 40617
0 40619 5 1 1 40618
0 40620 7 1 2 83057 39836
0 40621 5 1 1 40620
0 40622 7 1 2 40619 40621
0 40623 5 1 1 40622
0 40624 7 1 2 96251 40623
0 40625 5 1 1 40624
0 40626 7 1 2 80426 78199
0 40627 5 1 1 40626
0 40628 7 2 2 67093 77435
0 40629 5 1 1 96258
0 40630 7 2 2 72956 85305
0 40631 7 1 2 88981 96260
0 40632 7 1 2 96259 40631
0 40633 5 1 1 40632
0 40634 7 1 2 40627 40633
0 40635 5 1 1 40634
0 40636 7 1 2 68728 40635
0 40637 5 1 1 40636
0 40638 7 1 2 85290 40637
0 40639 5 1 1 40638
0 40640 7 1 2 59604 40639
0 40641 5 1 1 40640
0 40642 7 1 2 19355 88918
0 40643 5 1 1 40642
0 40644 7 1 2 59378 40643
0 40645 5 1 1 40644
0 40646 7 1 2 90263 88627
0 40647 5 1 1 40646
0 40648 7 1 2 76094 88632
0 40649 5 1 1 40648
0 40650 7 1 2 72236 40649
0 40651 5 1 1 40650
0 40652 7 1 2 40647 40651
0 40653 7 1 2 40645 40652
0 40654 5 1 1 40653
0 40655 7 1 2 84441 95826
0 40656 7 1 2 40654 40655
0 40657 5 1 1 40656
0 40658 7 1 2 40641 40657
0 40659 5 1 1 40658
0 40660 7 1 2 68902 40659
0 40661 5 1 1 40660
0 40662 7 1 2 40625 40661
0 40663 5 1 1 40662
0 40664 7 1 2 68444 40663
0 40665 5 1 1 40664
0 40666 7 4 2 61753 83586
0 40667 5 6 1 96262
0 40668 7 1 2 77034 96263
0 40669 5 1 1 40668
0 40670 7 1 2 40565 40669
0 40671 5 1 1 40670
0 40672 7 1 2 59945 40671
0 40673 5 1 1 40672
0 40674 7 1 2 76424 93775
0 40675 5 1 1 40674
0 40676 7 1 2 84550 40675
0 40677 5 2 1 40676
0 40678 7 1 2 69427 96272
0 40679 5 1 1 40678
0 40680 7 1 2 73288 95976
0 40681 5 1 1 40680
0 40682 7 1 2 70462 84500
0 40683 5 1 1 40682
0 40684 7 1 2 40681 40683
0 40685 7 1 2 40679 40684
0 40686 5 1 1 40685
0 40687 7 1 2 71895 40686
0 40688 5 1 1 40687
0 40689 7 1 2 40673 40688
0 40690 5 1 1 40689
0 40691 7 1 2 68069 40690
0 40692 5 1 1 40691
0 40693 7 1 2 95961 40692
0 40694 5 1 1 40693
0 40695 7 1 2 60574 68903
0 40696 7 1 2 40694 40695
0 40697 5 1 1 40696
0 40698 7 1 2 40665 40697
0 40699 5 1 1 40698
0 40700 7 1 2 86793 40699
0 40701 5 1 1 40700
0 40702 7 2 2 74800 84501
0 40703 5 1 1 96274
0 40704 7 1 2 71236 96275
0 40705 5 1 1 40704
0 40706 7 1 2 72237 91158
0 40707 5 2 1 40706
0 40708 7 1 2 40705 96276
0 40709 5 1 1 40708
0 40710 7 1 2 60575 40709
0 40711 5 1 1 40710
0 40712 7 1 2 91159 96155
0 40713 5 1 1 40712
0 40714 7 1 2 40711 40713
0 40715 5 1 1 40714
0 40716 7 1 2 67704 40715
0 40717 5 1 1 40716
0 40718 7 1 2 96052 40703
0 40719 5 1 1 40718
0 40720 7 1 2 91362 40719
0 40721 5 1 1 40720
0 40722 7 1 2 40717 40721
0 40723 5 1 1 40722
0 40724 7 1 2 92842 40723
0 40725 5 1 1 40724
0 40726 7 1 2 86226 92311
0 40727 5 1 1 40726
0 40728 7 1 2 92772 96087
0 40729 7 1 2 94261 40728
0 40730 5 1 1 40729
0 40731 7 1 2 40727 40730
0 40732 5 1 1 40731
0 40733 7 1 2 59379 40732
0 40734 5 1 1 40733
0 40735 7 1 2 87344 94932
0 40736 5 1 1 40735
0 40737 7 1 2 60689 69428
0 40738 7 1 2 93741 40737
0 40739 5 1 1 40738
0 40740 7 1 2 40736 40739
0 40741 5 1 1 40740
0 40742 7 1 2 67705 40741
0 40743 5 1 1 40742
0 40744 7 1 2 40734 40743
0 40745 5 1 1 40744
0 40746 7 1 2 59946 40745
0 40747 5 1 1 40746
0 40748 7 1 2 87299 95809
0 40749 5 1 1 40748
0 40750 7 1 2 40747 40749
0 40751 5 1 1 40750
0 40752 7 1 2 68729 40751
0 40753 5 1 1 40752
0 40754 7 3 2 79656 93930
0 40755 5 1 1 96278
0 40756 7 4 2 60690 67706
0 40757 7 1 2 71506 96281
0 40758 7 1 2 96279 40757
0 40759 5 1 1 40758
0 40760 7 1 2 40753 40759
0 40761 5 1 1 40760
0 40762 7 1 2 61104 40761
0 40763 5 1 1 40762
0 40764 7 1 2 84358 24675
0 40765 5 1 1 40764
0 40766 7 2 2 67707 91822
0 40767 5 1 1 96285
0 40768 7 1 2 40765 40767
0 40769 5 1 1 40768
0 40770 7 1 2 60691 87300
0 40771 7 1 2 40769 40770
0 40772 5 1 1 40771
0 40773 7 1 2 40763 40772
0 40774 5 1 1 40773
0 40775 7 1 2 86301 40774
0 40776 5 1 1 40775
0 40777 7 1 2 40725 40776
0 40778 5 1 1 40777
0 40779 7 1 2 59605 40778
0 40780 5 1 1 40779
0 40781 7 1 2 91797 93295
0 40782 5 1 1 40781
0 40783 7 1 2 65477 40782
0 40784 5 1 1 40783
0 40785 7 1 2 68445 40784
0 40786 5 1 1 40785
0 40787 7 1 2 92752 96011
0 40788 5 1 1 40787
0 40789 7 1 2 40786 40788
0 40790 5 1 1 40789
0 40791 7 1 2 84359 40790
0 40792 5 1 1 40791
0 40793 7 2 2 60576 96088
0 40794 7 2 2 73448 96287
0 40795 5 1 1 96289
0 40796 7 1 2 95470 95827
0 40797 5 1 1 40796
0 40798 7 1 2 40795 40797
0 40799 5 1 1 40798
0 40800 7 1 2 67708 40799
0 40801 5 1 1 40800
0 40802 7 1 2 18874 40801
0 40803 5 1 1 40802
0 40804 7 1 2 59947 40803
0 40805 5 1 1 40804
0 40806 7 1 2 88953 96290
0 40807 5 1 1 40806
0 40808 7 1 2 40805 40807
0 40809 5 1 1 40808
0 40810 7 1 2 63794 40809
0 40811 5 1 1 40810
0 40812 7 1 2 40792 40811
0 40813 5 1 1 40812
0 40814 7 1 2 64025 40813
0 40815 5 1 1 40814
0 40816 7 5 2 74996 83003
0 40817 5 2 1 96291
0 40818 7 1 2 93851 96292
0 40819 5 1 1 40818
0 40820 7 1 2 40815 40819
0 40821 5 1 1 40820
0 40822 7 1 2 86756 40821
0 40823 5 1 1 40822
0 40824 7 1 2 40780 40823
0 40825 7 1 2 40701 40824
0 40826 5 1 1 40825
0 40827 7 1 2 75340 40826
0 40828 5 1 1 40827
0 40829 7 1 2 61895 96111
0 40830 5 1 1 40829
0 40831 7 3 2 68904 83747
0 40832 7 1 2 60577 94438
0 40833 5 1 1 40832
0 40834 7 1 2 86626 40833
0 40835 5 2 1 40834
0 40836 7 1 2 86794 96301
0 40837 5 1 1 40836
0 40838 7 1 2 87721 40837
0 40839 5 1 1 40838
0 40840 7 1 2 96298 40839
0 40841 5 1 1 40840
0 40842 7 1 2 64026 86757
0 40843 7 1 2 89451 40842
0 40844 5 1 1 40843
0 40845 7 1 2 40841 40844
0 40846 5 1 1 40845
0 40847 7 1 2 83587 40846
0 40848 5 1 1 40847
0 40849 7 2 2 66564 86278
0 40850 7 2 2 83189 77576
0 40851 7 1 2 82376 96282
0 40852 7 1 2 96305 40851
0 40853 7 1 2 96303 40852
0 40854 5 1 1 40853
0 40855 7 1 2 40848 40854
0 40856 5 1 1 40855
0 40857 7 1 2 69943 40856
0 40858 5 1 1 40857
0 40859 7 2 2 75512 94779
0 40860 7 1 2 68070 96307
0 40861 5 1 1 40860
0 40862 7 1 2 89490 92451
0 40863 7 1 2 93677 40862
0 40864 5 1 1 40863
0 40865 7 1 2 40861 40864
0 40866 5 1 1 40865
0 40867 7 1 2 69577 40866
0 40868 5 1 1 40867
0 40869 7 1 2 93379 93629
0 40870 7 1 2 94517 40869
0 40871 5 1 1 40870
0 40872 7 1 2 40868 40871
0 40873 5 1 1 40872
0 40874 7 1 2 60692 40873
0 40875 5 1 1 40874
0 40876 7 1 2 64561 74132
0 40877 5 7 1 40876
0 40878 7 1 2 68071 79211
0 40879 7 1 2 69046 40878
0 40880 7 1 2 95002 40879
0 40881 7 1 2 96309 40880
0 40882 5 1 1 40881
0 40883 7 1 2 40875 40882
0 40884 5 1 1 40883
0 40885 7 1 2 79657 40884
0 40886 5 1 1 40885
0 40887 7 2 2 63795 96310
0 40888 7 1 2 87727 96316
0 40889 5 1 1 40888
0 40890 7 1 2 87202 92855
0 40891 5 1 1 40890
0 40892 7 1 2 87224 40891
0 40893 5 1 1 40892
0 40894 7 1 2 69726 92452
0 40895 7 1 2 40893 40894
0 40896 5 1 1 40895
0 40897 7 1 2 40889 40896
0 40898 5 1 1 40897
0 40899 7 1 2 96299 40898
0 40900 5 1 1 40899
0 40901 7 2 2 92357 93675
0 40902 5 2 1 96318
0 40903 7 1 2 75341 96319
0 40904 7 1 2 96317 40903
0 40905 5 1 1 40904
0 40906 7 1 2 40900 40905
0 40907 7 1 2 40886 40906
0 40908 7 1 2 40858 40907
0 40909 5 1 1 40908
0 40910 7 1 2 73512 40909
0 40911 5 1 1 40910
0 40912 7 1 2 40830 40911
0 40913 7 1 2 40828 40912
0 40914 7 1 2 40606 40913
0 40915 7 1 2 40041 40914
0 40916 5 1 1 40915
0 40917 7 1 2 68987 40916
0 40918 5 1 1 40917
0 40919 7 1 2 39531 40918
0 40920 5 1 1 40919
0 40921 7 1 2 69131 40920
0 40922 5 1 1 40921
0 40923 7 16 2 64027 68988
0 40924 7 1 2 69267 70903
0 40925 5 2 1 40924
0 40926 7 1 2 64562 90478
0 40927 5 1 1 40926
0 40928 7 1 2 96338 40927
0 40929 5 1 1 40928
0 40930 7 1 2 69858 40929
0 40931 5 1 1 40930
0 40932 7 1 2 70834 90670
0 40933 5 1 1 40932
0 40934 7 1 2 88577 40933
0 40935 7 1 2 40931 40934
0 40936 5 1 1 40935
0 40937 7 1 2 62149 40936
0 40938 5 1 1 40937
0 40939 7 1 2 70835 12674
0 40940 5 1 1 40939
0 40941 7 1 2 70073 88376
0 40942 5 1 1 40941
0 40943 7 2 2 71655 93158
0 40944 5 1 1 96340
0 40945 7 1 2 65274 40944
0 40946 5 1 1 40945
0 40947 7 1 2 40942 40946
0 40948 7 1 2 40940 40947
0 40949 7 1 2 40938 40948
0 40950 5 1 1 40949
0 40951 7 1 2 61585 40950
0 40952 5 1 1 40951
0 40953 7 2 2 83797 83247
0 40954 5 1 1 96342
0 40955 7 1 2 62150 74868
0 40956 7 1 2 96343 40955
0 40957 5 1 1 40956
0 40958 7 1 2 40952 40957
0 40959 5 1 1 40958
0 40960 7 1 2 67709 40959
0 40961 5 1 1 40960
0 40962 7 1 2 69578 77130
0 40963 5 1 1 40962
0 40964 7 1 2 77140 40963
0 40965 5 1 1 40964
0 40966 7 1 2 90589 40965
0 40967 5 1 1 40966
0 40968 7 1 2 77051 90479
0 40969 5 1 1 40968
0 40970 7 1 2 72500 90365
0 40971 5 1 1 40970
0 40972 7 1 2 79089 96339
0 40973 7 1 2 40971 40972
0 40974 7 1 2 40969 40973
0 40975 5 1 1 40974
0 40976 7 1 2 81053 40975
0 40977 5 2 1 40976
0 40978 7 1 2 40967 96344
0 40979 5 1 1 40978
0 40980 7 1 2 67094 40979
0 40981 5 1 1 40980
0 40982 7 3 2 79926 82101
0 40983 5 1 1 96346
0 40984 7 1 2 74231 96347
0 40985 5 1 1 40984
0 40986 7 1 2 40981 40985
0 40987 7 1 2 40961 40986
0 40988 5 1 1 40987
0 40989 7 1 2 68446 40988
0 40990 5 1 1 40989
0 40991 7 1 2 67710 88455
0 40992 5 1 1 40991
0 40993 7 1 2 65893 40992
0 40994 5 1 1 40993
0 40995 7 1 2 95557 40994
0 40996 5 1 1 40995
0 40997 7 1 2 21668 40996
0 40998 5 1 1 40997
0 40999 7 1 2 89287 40998
0 41000 5 1 1 40999
0 41001 7 1 2 95500 41000
0 41002 5 1 1 41001
0 41003 7 1 2 63529 41002
0 41004 5 1 1 41003
0 41005 7 1 2 60172 94840
0 41006 5 1 1 41005
0 41007 7 1 2 76188 41006
0 41008 5 1 1 41007
0 41009 7 1 2 61586 41008
0 41010 5 1 1 41009
0 41011 7 1 2 72362 41010
0 41012 5 1 1 41011
0 41013 7 1 2 77210 74326
0 41014 5 1 1 41013
0 41015 7 1 2 76648 85984
0 41016 5 1 1 41015
0 41017 7 1 2 61587 41016
0 41018 5 1 1 41017
0 41019 7 1 2 41014 41018
0 41020 5 1 1 41019
0 41021 7 1 2 90334 41020
0 41022 7 1 2 41012 41021
0 41023 5 1 1 41022
0 41024 7 1 2 60578 41023
0 41025 5 1 1 41024
0 41026 7 1 2 41004 41025
0 41027 7 1 2 40990 41026
0 41028 5 1 1 41027
0 41029 7 1 2 63121 41028
0 41030 5 1 1 41029
0 41031 7 1 2 68447 91328
0 41032 5 2 1 41031
0 41033 7 1 2 90660 96349
0 41034 5 1 1 41033
0 41035 7 1 2 66565 91039
0 41036 5 1 1 41035
0 41037 7 1 2 75697 41036
0 41038 5 1 1 41037
0 41039 7 1 2 71827 41038
0 41040 5 1 1 41039
0 41041 7 1 2 1105 84743
0 41042 5 2 1 41041
0 41043 7 1 2 78667 96351
0 41044 5 1 1 41043
0 41045 7 1 2 16638 41044
0 41046 7 1 2 41040 41045
0 41047 5 1 1 41046
0 41048 7 1 2 64325 41047
0 41049 5 1 1 41048
0 41050 7 1 2 41034 41049
0 41051 5 1 1 41050
0 41052 7 1 2 70325 41051
0 41053 5 1 1 41052
0 41054 7 1 2 69132 90891
0 41055 5 1 1 41054
0 41056 7 1 2 63530 41055
0 41057 5 1 1 41056
0 41058 7 1 2 69372 72170
0 41059 5 1 1 41058
0 41060 7 1 2 71237 74523
0 41061 7 1 2 41059 41060
0 41062 5 1 1 41061
0 41063 7 1 2 66566 41062
0 41064 5 1 1 41063
0 41065 7 1 2 41057 41064
0 41066 5 1 1 41065
0 41067 7 1 2 62731 41066
0 41068 5 1 1 41067
0 41069 7 1 2 82272 74082
0 41070 5 1 1 41069
0 41071 7 1 2 70836 41070
0 41072 5 2 1 41071
0 41073 7 2 2 90911 96353
0 41074 7 1 2 71524 96355
0 41075 5 1 1 41074
0 41076 7 1 2 85929 41075
0 41077 5 1 1 41076
0 41078 7 1 2 90732 94860
0 41079 5 1 1 41078
0 41080 7 1 2 90661 41079
0 41081 5 1 1 41080
0 41082 7 1 2 85751 86949
0 41083 5 1 1 41082
0 41084 7 1 2 76012 85047
0 41085 5 1 1 41084
0 41086 7 1 2 75698 41085
0 41087 7 1 2 85055 90733
0 41088 5 1 1 41087
0 41089 7 1 2 95390 41088
0 41090 5 1 1 41089
0 41091 7 1 2 94576 96352
0 41092 5 1 1 41091
0 41093 7 1 2 41090 41092
0 41094 7 1 2 41086 41093
0 41095 5 1 1 41094
0 41096 7 1 2 72363 41095
0 41097 5 1 1 41096
0 41098 7 1 2 41083 41097
0 41099 7 1 2 41081 41098
0 41100 7 1 2 41077 41099
0 41101 7 1 2 41068 41100
0 41102 7 1 2 41053 41101
0 41103 5 1 1 41102
0 41104 7 1 2 60579 41103
0 41105 5 1 1 41104
0 41106 7 1 2 64563 91145
0 41107 5 1 1 41106
0 41108 7 1 2 89040 41107
0 41109 5 1 1 41108
0 41110 7 1 2 64801 41109
0 41111 5 1 1 41110
0 41112 7 2 2 37190 41111
0 41113 5 1 1 96357
0 41114 7 1 2 71578 41113
0 41115 5 1 1 41114
0 41116 7 1 2 88471 90848
0 41117 5 1 1 41116
0 41118 7 2 2 76316 72238
0 41119 5 2 1 96359
0 41120 7 1 2 65275 96361
0 41121 5 2 1 41120
0 41122 7 1 2 59606 96363
0 41123 5 1 1 41122
0 41124 7 1 2 60387 90542
0 41125 5 1 1 41124
0 41126 7 1 2 70837 41125
0 41127 7 1 2 41123 41126
0 41128 5 1 1 41127
0 41129 7 1 2 79127 41128
0 41130 7 1 2 41117 41129
0 41131 7 1 2 41115 41130
0 41132 5 1 1 41131
0 41133 7 1 2 84832 41132
0 41134 5 2 1 41133
0 41135 7 1 2 69859 85086
0 41136 5 1 1 41135
0 41137 7 1 2 78480 41136
0 41138 5 1 1 41137
0 41139 7 1 2 64564 41138
0 41140 5 1 1 41139
0 41141 7 1 2 78297 85087
0 41142 5 1 1 41141
0 41143 7 1 2 67352 41142
0 41144 7 1 2 41140 41143
0 41145 5 1 1 41144
0 41146 7 1 2 61105 90976
0 41147 5 1 1 41146
0 41148 7 1 2 41145 41147
0 41149 5 1 1 41148
0 41150 7 1 2 59948 41149
0 41151 5 1 1 41150
0 41152 7 1 2 66567 95248
0 41153 5 2 1 41152
0 41154 7 1 2 59607 96367
0 41155 5 1 1 41154
0 41156 7 2 2 69579 93178
0 41157 5 2 1 96369
0 41158 7 2 2 41155 96371
0 41159 7 1 2 66568 96213
0 41160 5 2 1 41159
0 41161 7 1 2 69944 96375
0 41162 5 1 1 41161
0 41163 7 1 2 80764 41162
0 41164 7 1 2 96373 41163
0 41165 7 1 2 41151 41164
0 41166 5 1 1 41165
0 41167 7 1 2 65478 41166
0 41168 5 1 1 41167
0 41169 7 1 2 96365 41168
0 41170 5 1 1 41169
0 41171 7 1 2 68448 41170
0 41172 5 1 1 41171
0 41173 7 1 2 71932 91535
0 41174 5 1 1 41173
0 41175 7 2 2 68072 41174
0 41176 5 1 1 96377
0 41177 7 1 2 65276 41176
0 41178 5 1 1 41177
0 41179 7 1 2 83707 41178
0 41180 5 1 1 41179
0 41181 7 1 2 41172 41180
0 41182 7 1 2 41105 41181
0 41183 7 1 2 41030 41182
0 41184 5 1 1 41183
0 41185 7 1 2 61754 41184
0 41186 5 1 1 41185
0 41187 7 2 2 67711 76408
0 41188 5 1 1 96379
0 41189 7 1 2 89796 41188
0 41190 5 1 1 41189
0 41191 7 1 2 86678 41190
0 41192 5 3 1 41191
0 41193 7 1 2 92626 92791
0 41194 5 1 1 41193
0 41195 7 1 2 96381 41194
0 41196 5 1 1 41195
0 41197 7 1 2 69945 41196
0 41198 5 1 1 41197
0 41199 7 1 2 79442 90977
0 41200 5 1 1 41199
0 41201 7 1 2 19816 15472
0 41202 5 1 1 41201
0 41203 7 1 2 86679 41202
0 41204 5 3 1 41203
0 41205 7 3 2 67712 73357
0 41206 5 2 1 96387
0 41207 7 3 2 68449 96388
0 41208 7 1 2 92627 96392
0 41209 5 1 1 41208
0 41210 7 1 2 96384 41209
0 41211 5 1 1 41210
0 41212 7 1 2 67353 41211
0 41213 5 1 1 41212
0 41214 7 1 2 41200 41213
0 41215 7 1 2 41198 41214
0 41216 5 1 1 41215
0 41217 7 1 2 61106 41216
0 41218 5 1 1 41217
0 41219 7 1 2 66569 83203
0 41220 5 2 1 41219
0 41221 7 1 2 85930 15499
0 41222 5 1 1 41221
0 41223 7 2 2 96395 41222
0 41224 5 1 1 96397
0 41225 7 1 2 66736 96398
0 41226 5 1 1 41225
0 41227 7 2 2 80814 79292
0 41228 7 1 2 72523 96399
0 41229 5 1 1 41228
0 41230 7 1 2 41226 41229
0 41231 7 1 2 41218 41230
0 41232 5 1 1 41231
0 41233 7 1 2 59949 41232
0 41234 5 1 1 41233
0 41235 7 1 2 89877 91969
0 41236 5 1 1 41235
0 41237 7 1 2 61588 82387
0 41238 5 1 1 41237
0 41239 7 1 2 96374 41238
0 41240 5 1 1 41239
0 41241 7 1 2 68450 41240
0 41242 5 1 1 41241
0 41243 7 1 2 71896 84833
0 41244 5 2 1 41243
0 41245 7 1 2 85887 96376
0 41246 5 1 1 41245
0 41247 7 1 2 96401 41246
0 41248 7 2 2 41242 41247
0 41249 7 1 2 90187 96403
0 41250 5 1 1 41249
0 41251 7 1 2 66737 41250
0 41252 5 1 1 41251
0 41253 7 1 2 41236 41252
0 41254 7 1 2 41234 41253
0 41255 5 1 1 41254
0 41256 7 1 2 90637 41255
0 41257 5 1 1 41256
0 41258 7 1 2 68730 41257
0 41259 7 1 2 41186 41258
0 41260 5 1 1 41259
0 41261 7 2 2 81821 75017
0 41262 5 1 1 96405
0 41263 7 1 2 91536 41262
0 41264 5 1 1 41263
0 41265 7 1 2 61107 41264
0 41266 5 1 1 41265
0 41267 7 1 2 64565 90269
0 41268 5 2 1 41267
0 41269 7 1 2 74535 91528
0 41270 7 1 2 96407 41269
0 41271 5 1 1 41270
0 41272 7 2 2 41266 41271
0 41273 7 1 2 63531 96409
0 41274 5 1 1 41273
0 41275 7 1 2 61589 41274
0 41276 5 1 1 41275
0 41277 7 1 2 71589 95270
0 41278 5 1 1 41277
0 41279 7 1 2 67713 41278
0 41280 5 1 1 41279
0 41281 7 1 2 74602 74801
0 41282 5 1 1 41281
0 41283 7 1 2 93108 41282
0 41284 5 1 1 41283
0 41285 7 1 2 67354 41284
0 41286 5 1 1 41285
0 41287 7 1 2 74423 41286
0 41288 7 1 2 41280 41287
0 41289 5 1 1 41288
0 41290 7 1 2 68451 41289
0 41291 5 1 1 41290
0 41292 7 2 2 79893 76445
0 41293 5 1 1 96411
0 41294 7 1 2 20078 41293
0 41295 7 1 2 41291 41294
0 41296 5 1 1 41295
0 41297 7 1 2 68073 41296
0 41298 5 1 1 41297
0 41299 7 1 2 41276 41298
0 41300 5 1 1 41299
0 41301 7 1 2 95834 41300
0 41302 5 1 1 41301
0 41303 7 4 2 80874 81795
0 41304 5 1 1 96413
0 41305 7 1 2 63796 41304
0 41306 7 1 2 41302 41305
0 41307 5 1 1 41306
0 41308 7 1 2 61896 41307
0 41309 7 1 2 41260 41308
0 41310 5 1 1 41309
0 41311 7 1 2 72524 89565
0 41312 5 1 1 41311
0 41313 7 1 2 41224 41312
0 41314 5 1 1 41313
0 41315 7 1 2 59950 41314
0 41316 5 1 1 41315
0 41317 7 1 2 96404 41316
0 41318 5 2 1 41317
0 41319 7 1 2 66880 96417
0 41320 5 1 1 41319
0 41321 7 5 2 60940 66881
0 41322 7 1 2 92792 96419
0 41323 5 1 1 41322
0 41324 7 1 2 96382 41323
0 41325 5 1 1 41324
0 41326 7 1 2 69946 41325
0 41327 5 1 1 41326
0 41328 7 1 2 96393 96420
0 41329 5 1 1 41328
0 41330 7 1 2 96385 41329
0 41331 5 1 1 41330
0 41332 7 1 2 67355 41331
0 41333 5 1 1 41332
0 41334 7 1 2 90978 94349
0 41335 5 1 1 41334
0 41336 7 1 2 41333 41335
0 41337 7 1 2 41327 41336
0 41338 5 1 1 41337
0 41339 7 1 2 72239 41338
0 41340 5 1 1 41339
0 41341 7 1 2 41320 41340
0 41342 5 1 1 41341
0 41343 7 1 2 68731 96414
0 41344 7 1 2 41342 41343
0 41345 5 1 1 41344
0 41346 7 1 2 41310 41345
0 41347 5 1 1 41346
0 41348 7 1 2 60693 41347
0 41349 5 1 1 41348
0 41350 7 1 2 79191 87557
0 41351 5 1 1 41350
0 41352 7 1 2 60580 41351
0 41353 5 1 1 41352
0 41354 7 2 2 67714 73384
0 41355 5 1 1 96424
0 41356 7 1 2 89087 96425
0 41357 5 1 1 41356
0 41358 7 1 2 59951 24634
0 41359 5 1 1 41358
0 41360 7 1 2 62732 73441
0 41361 5 1 1 41360
0 41362 7 1 2 59380 41361
0 41363 5 2 1 41362
0 41364 7 1 2 81815 96426
0 41365 5 1 1 41364
0 41366 7 1 2 67095 41365
0 41367 5 1 1 41366
0 41368 7 1 2 76264 82079
0 41369 5 1 1 41368
0 41370 7 1 2 91504 41369
0 41371 7 1 2 41367 41370
0 41372 5 1 1 41371
0 41373 7 1 2 61108 41372
0 41374 5 1 1 41373
0 41375 7 1 2 41359 41374
0 41376 5 1 1 41375
0 41377 7 1 2 68074 41376
0 41378 5 1 1 41377
0 41379 7 1 2 41357 41378
0 41380 5 2 1 41379
0 41381 7 1 2 61590 96428
0 41382 5 1 1 41381
0 41383 7 1 2 41353 41382
0 41384 5 1 1 41383
0 41385 7 1 2 84360 41384
0 41386 5 1 1 41385
0 41387 7 2 2 68732 77482
0 41388 5 1 1 96430
0 41389 7 1 2 94794 41388
0 41390 5 1 1 41389
0 41391 7 2 2 62733 89779
0 41392 5 1 1 96432
0 41393 7 1 2 93132 96433
0 41394 5 1 1 41393
0 41395 7 1 2 41390 41394
0 41396 5 1 1 41395
0 41397 7 1 2 61755 41396
0 41398 5 1 1 41397
0 41399 7 1 2 59381 69312
0 41400 5 1 1 41399
0 41401 7 1 2 70288 95888
0 41402 5 1 1 41401
0 41403 7 1 2 41400 41402
0 41404 5 1 1 41403
0 41405 7 1 2 59608 41404
0 41406 5 1 1 41405
0 41407 7 1 2 59952 92932
0 41408 5 1 1 41407
0 41409 7 1 2 61109 92880
0 41410 5 1 1 41409
0 41411 7 1 2 82238 41410
0 41412 7 1 2 41408 41411
0 41413 7 1 2 41406 41412
0 41414 7 1 2 80266 76013
0 41415 7 1 2 78100 41414
0 41416 5 1 1 41415
0 41417 7 1 2 69429 41416
0 41418 5 1 1 41417
0 41419 7 1 2 69473 69334
0 41420 5 1 1 41419
0 41421 7 1 2 59382 41420
0 41422 5 1 1 41421
0 41423 7 1 2 41418 41422
0 41424 7 1 2 41413 41423
0 41425 5 1 1 41424
0 41426 7 1 2 79658 84846
0 41427 7 1 2 41425 41426
0 41428 5 1 1 41427
0 41429 7 1 2 41398 41428
0 41430 7 1 2 41386 41429
0 41431 5 1 1 41430
0 41432 7 1 2 68452 41431
0 41433 5 1 1 41432
0 41434 7 5 2 63122 94405
0 41435 5 3 1 96434
0 41436 7 1 2 95561 96435
0 41437 5 1 1 41436
0 41438 7 1 2 80370 81126
0 41439 5 5 1 41438
0 41440 7 1 2 96378 96442
0 41441 5 1 1 41440
0 41442 7 1 2 41437 41441
0 41443 5 1 1 41442
0 41444 7 1 2 68733 41443
0 41445 5 1 1 41444
0 41446 7 1 2 71933 73463
0 41447 5 1 1 41446
0 41448 7 1 2 68075 41447
0 41449 5 1 1 41448
0 41450 7 1 2 66570 41449
0 41451 7 1 2 96410 41450
0 41452 5 1 1 41451
0 41453 7 1 2 83153 41452
0 41454 5 1 1 41453
0 41455 7 1 2 41445 41454
0 41456 7 1 2 41433 41455
0 41457 5 1 1 41456
0 41458 7 1 2 61897 41457
0 41459 5 1 1 41458
0 41460 7 2 2 89936 96429
0 41461 7 1 2 80875 86241
0 41462 7 1 2 96447 41461
0 41463 5 1 1 41462
0 41464 7 1 2 41459 41463
0 41465 5 1 1 41464
0 41466 7 1 2 60694 41465
0 41467 5 1 1 41466
0 41468 7 1 2 87149 88136
0 41469 7 1 2 96448 41468
0 41470 5 1 1 41469
0 41471 7 1 2 41467 41470
0 41472 5 1 1 41471
0 41473 7 1 2 76796 41472
0 41474 5 1 1 41473
0 41475 7 2 2 92893 94394
0 41476 5 1 1 96449
0 41477 7 1 2 59953 96450
0 41478 5 1 1 41477
0 41479 7 1 2 66571 71325
0 41480 5 2 1 41479
0 41481 7 1 2 74786 95882
0 41482 5 1 1 41481
0 41483 7 1 2 96451 41482
0 41484 5 1 1 41483
0 41485 7 1 2 64566 41484
0 41486 5 1 1 41485
0 41487 7 2 2 60388 96368
0 41488 5 1 1 96453
0 41489 7 2 2 61591 88954
0 41490 5 1 1 96455
0 41491 7 1 2 91537 41490
0 41492 5 1 1 41491
0 41493 7 1 2 96454 41492
0 41494 7 1 2 41486 41493
0 41495 5 1 1 41494
0 41496 7 2 2 76929 72240
0 41497 5 2 1 96457
0 41498 7 1 2 80763 86876
0 41499 7 1 2 96458 41498
0 41500 5 1 1 41499
0 41501 7 1 2 41495 41500
0 41502 5 1 1 41501
0 41503 7 1 2 68453 41502
0 41504 5 1 1 41503
0 41505 7 1 2 41478 41504
0 41506 5 2 1 41505
0 41507 7 2 2 80876 85708
0 41508 7 1 2 96461 96463
0 41509 5 1 1 41508
0 41510 7 1 2 72132 78264
0 41511 5 1 1 41510
0 41512 7 2 2 63123 82287
0 41513 5 5 1 96465
0 41514 7 1 2 91188 96467
0 41515 7 1 2 80263 41514
0 41516 5 1 1 41515
0 41517 7 1 2 41511 41516
0 41518 5 1 1 41517
0 41519 7 1 2 69580 41518
0 41520 5 1 1 41519
0 41521 7 1 2 59609 90935
0 41522 5 1 1 41521
0 41523 7 1 2 81708 41522
0 41524 5 1 1 41523
0 41525 7 1 2 68076 41524
0 41526 5 1 1 41525
0 41527 7 1 2 41520 41526
0 41528 5 1 1 41527
0 41529 7 1 2 61110 41528
0 41530 5 1 1 41529
0 41531 7 2 2 76502 94122
0 41532 5 1 1 96472
0 41533 7 1 2 69193 96473
0 41534 5 1 1 41533
0 41535 7 1 2 41530 41534
0 41536 5 1 1 41535
0 41537 7 1 2 91680 41536
0 41538 5 1 1 41537
0 41539 7 2 2 95471 95869
0 41540 5 1 1 96474
0 41541 7 1 2 65479 41540
0 41542 5 1 1 41541
0 41543 7 1 2 69947 41542
0 41544 5 1 1 41543
0 41545 7 1 2 72866 80460
0 41546 7 1 2 92043 41545
0 41547 5 1 1 41546
0 41548 7 1 2 41544 41547
0 41549 5 1 1 41548
0 41550 7 1 2 59610 41549
0 41551 5 1 1 41550
0 41552 7 1 2 91766 41551
0 41553 5 1 1 41552
0 41554 7 1 2 75342 41553
0 41555 5 1 1 41554
0 41556 7 1 2 63797 41555
0 41557 7 1 2 41538 41556
0 41558 5 1 1 41557
0 41559 7 1 2 91538 19248
0 41560 5 1 1 41559
0 41561 7 1 2 62734 41560
0 41562 5 1 1 41561
0 41563 7 1 2 4795 41562
0 41564 5 1 1 41563
0 41565 7 1 2 75850 41564
0 41566 5 1 1 41565
0 41567 7 1 2 71375 13763
0 41568 5 1 1 41567
0 41569 7 1 2 59383 41568
0 41570 5 1 1 41569
0 41571 7 1 2 67356 81810
0 41572 5 1 1 41571
0 41573 7 1 2 89000 41572
0 41574 7 1 2 41570 41573
0 41575 5 1 1 41574
0 41576 7 1 2 89402 41575
0 41577 5 1 1 41576
0 41578 7 1 2 41566 41577
0 41579 5 1 1 41578
0 41580 7 1 2 63124 41579
0 41581 5 1 1 41580
0 41582 7 1 2 66064 95584
0 41583 5 1 1 41582
0 41584 7 1 2 67715 41583
0 41585 5 1 1 41584
0 41586 7 1 2 63125 41585
0 41587 5 1 1 41586
0 41588 7 1 2 82183 41587
0 41589 5 1 1 41588
0 41590 7 1 2 68734 41589
0 41591 7 1 2 41581 41590
0 41592 5 1 1 41591
0 41593 7 1 2 61756 41592
0 41594 7 1 2 41558 41593
0 41595 5 1 1 41594
0 41596 7 1 2 80363 89937
0 41597 5 2 1 41596
0 41598 7 1 2 89954 40273
0 41599 5 1 1 41598
0 41600 7 1 2 75513 41599
0 41601 5 1 1 41600
0 41602 7 1 2 96476 41601
0 41603 5 1 1 41602
0 41604 7 1 2 60941 41603
0 41605 5 1 1 41604
0 41606 7 1 2 76265 96167
0 41607 5 1 1 41606
0 41608 7 1 2 41605 41607
0 41609 5 1 1 41608
0 41610 7 1 2 67357 41609
0 41611 5 1 1 41610
0 41612 7 2 2 60389 92350
0 41613 7 1 2 84794 96478
0 41614 5 1 1 41613
0 41615 7 1 2 41611 41614
0 41616 5 1 1 41615
0 41617 7 1 2 59954 41616
0 41618 5 1 1 41617
0 41619 7 1 2 68735 12134
0 41620 5 1 1 41619
0 41621 7 1 2 63798 20438
0 41622 5 1 1 41621
0 41623 7 1 2 96475 41622
0 41624 7 1 2 41620 41623
0 41625 5 1 1 41624
0 41626 7 1 2 67358 91761
0 41627 7 1 2 89688 41626
0 41628 5 1 1 41627
0 41629 7 1 2 41625 41628
0 41630 5 1 1 41629
0 41631 7 1 2 69948 41630
0 41632 5 1 1 41631
0 41633 7 1 2 74207 85400
0 41634 5 1 1 41633
0 41635 7 2 2 83553 78437
0 41636 5 1 1 96480
0 41637 7 1 2 41634 41636
0 41638 5 1 1 41637
0 41639 7 1 2 69581 41638
0 41640 5 1 1 41639
0 41641 7 1 2 88996 89689
0 41642 5 1 1 41641
0 41643 7 1 2 41640 41642
0 41644 5 1 1 41643
0 41645 7 1 2 60581 41644
0 41646 5 1 1 41645
0 41647 7 1 2 41632 41646
0 41648 5 1 1 41647
0 41649 7 1 2 75343 41648
0 41650 5 1 1 41649
0 41651 7 1 2 92062 92753
0 41652 7 1 2 88753 41651
0 41653 5 1 1 41652
0 41654 7 1 2 89955 41653
0 41655 5 1 1 41654
0 41656 7 1 2 75514 41655
0 41657 5 1 1 41656
0 41658 7 1 2 41657 96477
0 41659 5 1 1 41658
0 41660 7 1 2 88955 41659
0 41661 5 1 1 41660
0 41662 7 1 2 78228 36969
0 41663 5 1 1 41662
0 41664 7 1 2 41663 96168
0 41665 5 1 1 41664
0 41666 7 1 2 41661 41665
0 41667 7 1 2 41650 41666
0 41668 7 1 2 41618 41667
0 41669 7 1 2 41595 41668
0 41670 5 1 1 41669
0 41671 7 1 2 67096 41670
0 41672 5 1 1 41671
0 41673 7 1 2 70988 91681
0 41674 5 1 1 41673
0 41675 7 4 2 75344 76266
0 41676 7 1 2 93179 96482
0 41677 5 1 1 41676
0 41678 7 1 2 41674 41677
0 41679 5 1 1 41678
0 41680 7 1 2 83248 41679
0 41681 5 1 1 41680
0 41682 7 1 2 91862 41681
0 41683 5 1 1 41682
0 41684 7 1 2 66738 41683
0 41685 5 1 1 41684
0 41686 7 9 2 66739 91682
0 41687 5 3 1 96486
0 41688 7 1 2 88956 96487
0 41689 5 1 1 41688
0 41690 7 1 2 74869 86890
0 41691 5 1 1 41690
0 41692 7 1 2 84390 41691
0 41693 5 1 1 41692
0 41694 7 1 2 61757 41693
0 41695 5 1 1 41694
0 41696 7 1 2 41689 41695
0 41697 5 1 1 41696
0 41698 7 1 2 77263 41697
0 41699 5 1 1 41698
0 41700 7 1 2 65277 40954
0 41701 5 1 1 41700
0 41702 7 1 2 85498 41701
0 41703 5 1 1 41702
0 41704 7 1 2 83720 41703
0 41705 5 1 1 41704
0 41706 7 1 2 61758 41705
0 41707 5 1 1 41706
0 41708 7 1 2 41699 41707
0 41709 7 1 2 41685 41708
0 41710 5 1 1 41709
0 41711 7 1 2 68454 41710
0 41712 5 1 1 41711
0 41713 7 1 2 96364 96443
0 41714 5 1 1 41713
0 41715 7 1 2 81394 96360
0 41716 5 1 1 41715
0 41717 7 1 2 80378 41716
0 41718 5 1 1 41717
0 41719 7 1 2 61592 41718
0 41720 5 1 1 41719
0 41721 7 1 2 41714 41720
0 41722 5 1 1 41721
0 41723 7 1 2 68077 41722
0 41724 5 1 1 41723
0 41725 7 1 2 66065 81816
0 41726 5 1 1 41725
0 41727 7 1 2 59384 41726
0 41728 5 1 1 41727
0 41729 7 1 2 61111 5070
0 41730 5 1 1 41729
0 41731 7 1 2 71435 41730
0 41732 7 1 2 41728 41731
0 41733 5 1 1 41732
0 41734 7 4 2 63532 90036
0 41735 7 3 2 79659 96498
0 41736 5 2 1 96502
0 41737 7 1 2 91202 96503
0 41738 7 1 2 41733 41737
0 41739 5 1 1 41738
0 41740 7 1 2 41724 41739
0 41741 7 1 2 41712 41740
0 41742 5 1 1 41741
0 41743 7 1 2 68736 41742
0 41744 5 1 1 41743
0 41745 7 1 2 71376 77052
0 41746 5 1 1 41745
0 41747 7 1 2 71424 92160
0 41748 7 1 2 41746 41747
0 41749 5 1 1 41748
0 41750 7 1 2 5488 41749
0 41751 5 1 1 41750
0 41752 7 1 2 61112 41751
0 41753 5 1 1 41752
0 41754 7 1 2 85125 41753
0 41755 5 1 1 41754
0 41756 7 1 2 79660 41755
0 41757 5 1 1 41756
0 41758 7 1 2 80877 88957
0 41759 5 1 1 41758
0 41760 7 1 2 41757 41759
0 41761 5 1 1 41760
0 41762 7 1 2 68455 41761
0 41763 5 1 1 41762
0 41764 7 1 2 67716 77245
0 41765 5 1 1 41764
0 41766 7 1 2 78934 41765
0 41767 7 1 2 96427 41766
0 41768 5 1 1 41767
0 41769 7 1 2 89452 41768
0 41770 5 1 1 41769
0 41771 7 1 2 41763 41770
0 41772 5 1 1 41771
0 41773 7 1 2 63799 41772
0 41774 5 1 1 41773
0 41775 7 1 2 41744 41774
0 41776 7 1 2 41672 41775
0 41777 5 1 1 41776
0 41778 7 1 2 61898 41777
0 41779 5 1 1 41778
0 41780 7 1 2 41509 41779
0 41781 5 1 1 41780
0 41782 7 1 2 60695 41781
0 41783 5 1 1 41782
0 41784 7 5 2 68737 87630
0 41785 7 1 2 96242 96507
0 41786 7 1 2 96462 41785
0 41787 5 1 1 41786
0 41788 7 1 2 41783 41787
0 41789 5 1 1 41788
0 41790 7 1 2 70201 41789
0 41791 5 1 1 41790
0 41792 7 1 2 66740 73212
0 41793 5 1 1 41792
0 41794 7 1 2 72133 93793
0 41795 7 1 2 41793 41794
0 41796 5 1 1 41795
0 41797 7 1 2 71336 84502
0 41798 5 1 1 41797
0 41799 7 1 2 71728 96180
0 41800 5 1 1 41799
0 41801 7 1 2 41798 41800
0 41802 7 1 2 41796 41801
0 41803 5 1 1 41802
0 41804 7 1 2 90638 41803
0 41805 5 1 1 41804
0 41806 7 2 2 81796 85142
0 41807 5 3 1 96512
0 41808 7 1 2 65480 89144
0 41809 5 1 1 41808
0 41810 7 1 2 65894 41809
0 41811 5 1 1 41810
0 41812 7 1 2 80334 86434
0 41813 7 1 2 76267 41812
0 41814 7 1 2 41811 41813
0 41815 5 1 1 41814
0 41816 7 1 2 96514 41815
0 41817 5 1 1 41816
0 41818 7 1 2 72021 71326
0 41819 5 1 1 41818
0 41820 7 1 2 41817 41819
0 41821 5 1 1 41820
0 41822 7 1 2 41805 41821
0 41823 5 1 1 41822
0 41824 7 1 2 61899 41823
0 41825 5 1 1 41824
0 41826 7 5 2 60173 86483
0 41827 7 1 2 86435 92620
0 41828 7 1 2 96517 41827
0 41829 7 1 2 74187 41828
0 41830 5 1 1 41829
0 41831 7 1 2 41825 41830
0 41832 5 1 1 41831
0 41833 7 1 2 60696 41832
0 41834 5 1 1 41833
0 41835 7 1 2 80102 83158
0 41836 7 1 2 95714 41835
0 41837 7 1 2 94933 41836
0 41838 7 1 2 74188 41837
0 41839 5 1 1 41838
0 41840 7 1 2 41834 41839
0 41841 5 1 1 41840
0 41842 7 1 2 68078 41841
0 41843 5 1 1 41842
0 41844 7 3 2 68738 86279
0 41845 7 1 2 87712 96522
0 41846 7 1 2 93349 41845
0 41847 5 1 1 41846
0 41848 7 1 2 41843 41847
0 41849 5 1 1 41848
0 41850 7 1 2 68456 41849
0 41851 5 1 1 41850
0 41852 7 3 2 60582 86737
0 41853 7 2 2 61759 96525
0 41854 5 1 1 96528
0 41855 7 1 2 86771 41854
0 41856 5 7 1 41855
0 41857 7 1 2 81349 96530
0 41858 5 1 1 41857
0 41859 7 1 2 60697 96187
0 41860 5 2 1 41859
0 41861 7 1 2 41858 96537
0 41862 5 1 1 41861
0 41863 7 1 2 75733 84625
0 41864 7 1 2 74421 41863
0 41865 7 1 2 41862 41864
0 41866 5 1 1 41865
0 41867 7 1 2 41851 41866
0 41868 5 1 1 41867
0 41869 7 1 2 71238 41868
0 41870 5 1 1 41869
0 41871 7 1 2 65608 96418
0 41872 5 1 1 41871
0 41873 7 3 2 65609 69194
0 41874 7 1 2 80957 96539
0 41875 5 1 1 41874
0 41876 7 1 2 96383 41875
0 41877 5 1 1 41876
0 41878 7 1 2 69949 41877
0 41879 5 1 1 41878
0 41880 7 2 2 65610 60942
0 41881 7 1 2 96394 96542
0 41882 5 1 1 41881
0 41883 7 1 2 96386 41882
0 41884 5 1 1 41883
0 41885 7 1 2 67359 41884
0 41886 5 1 1 41885
0 41887 7 1 2 90979 92281
0 41888 5 1 1 41887
0 41889 7 1 2 41886 41888
0 41890 7 1 2 41879 41889
0 41891 5 1 1 41890
0 41892 7 1 2 72241 41891
0 41893 5 1 1 41892
0 41894 7 1 2 41872 41893
0 41895 5 1 1 41894
0 41896 7 1 2 91748 96523
0 41897 7 1 2 41895 41896
0 41898 5 1 1 41897
0 41899 7 1 2 41870 41898
0 41900 7 1 2 41791 41899
0 41901 7 1 2 41474 41900
0 41902 7 1 2 41349 41901
0 41903 5 1 1 41902
0 41904 7 1 2 96322 41903
0 41905 5 1 1 41904
0 41906 7 1 2 59611 96089
0 41907 7 1 2 92195 41906
0 41908 5 1 1 41907
0 41909 7 1 2 40557 41908
0 41910 5 1 1 41909
0 41911 7 1 2 59385 41910
0 41912 5 1 1 41911
0 41913 7 2 2 83058 85527
0 41914 5 1 1 96544
0 41915 7 1 2 41912 41914
0 41916 5 1 1 41915
0 41917 7 1 2 75386 41916
0 41918 5 1 1 41917
0 41919 7 2 2 85528 94439
0 41920 7 2 2 68079 96546
0 41921 5 1 1 96548
0 41922 7 1 2 41918 41921
0 41923 5 1 1 41922
0 41924 7 1 2 66882 41923
0 41925 5 1 1 41924
0 41926 7 1 2 75387 93931
0 41927 5 1 1 41926
0 41928 7 1 2 66883 96228
0 41929 5 2 1 41928
0 41930 7 1 2 41927 96550
0 41931 5 1 1 41930
0 41932 7 1 2 76059 41931
0 41933 5 1 1 41932
0 41934 7 6 2 79713 94440
0 41935 5 1 1 96552
0 41936 7 1 2 64028 70463
0 41937 7 1 2 96553 41936
0 41938 5 1 1 41937
0 41939 7 1 2 41933 41938
0 41940 7 1 2 41925 41939
0 41941 5 1 1 41940
0 41942 7 1 2 61113 41941
0 41943 5 1 1 41942
0 41944 7 1 2 81029 92161
0 41945 7 1 2 92781 41944
0 41946 5 1 1 41945
0 41947 7 2 2 61593 86106
0 41948 5 1 1 96558
0 41949 7 1 2 87334 94350
0 41950 5 1 1 41949
0 41951 7 1 2 41948 41950
0 41952 5 1 1 41951
0 41953 7 1 2 60390 41952
0 41954 5 1 1 41953
0 41955 7 1 2 85912 87345
0 41956 5 1 1 41955
0 41957 7 2 2 26809 41956
0 41958 5 1 1 96560
0 41959 7 1 2 41954 96561
0 41960 5 2 1 41959
0 41961 7 1 2 63800 76425
0 41962 7 1 2 96562 41961
0 41963 5 1 1 41962
0 41964 7 1 2 41946 41963
0 41965 5 1 1 41964
0 41966 7 1 2 70289 41965
0 41967 5 1 1 41966
0 41968 7 1 2 41943 41967
0 41969 5 1 1 41968
0 41970 7 1 2 68989 41969
0 41971 5 1 1 41970
0 41972 7 1 2 61114 79714
0 41973 5 1 1 41972
0 41974 7 1 2 68080 92782
0 41975 5 1 1 41974
0 41976 7 1 2 41973 41975
0 41977 5 1 1 41976
0 41978 7 1 2 68457 92554
0 41979 7 1 2 41977 41978
0 41980 5 1 1 41979
0 41981 7 3 2 61115 87072
0 41982 7 3 2 83554 87335
0 41983 7 1 2 96564 96567
0 41984 5 1 1 41983
0 41985 7 1 2 41980 41984
0 41986 5 1 1 41985
0 41987 7 1 2 68990 41986
0 41988 5 1 1 41987
0 41989 7 6 2 61900 68739
0 41990 7 3 2 94750 96570
0 41991 7 1 2 89656 96576
0 41992 5 1 1 41991
0 41993 7 1 2 41988 41992
0 41994 5 1 1 41993
0 41995 7 1 2 59386 41994
0 41996 5 1 1 41995
0 41997 7 3 2 61116 94210
0 41998 7 1 2 96563 96579
0 41999 5 1 1 41998
0 42000 7 1 2 41996 41999
0 42001 5 1 1 42000
0 42002 7 1 2 69430 42001
0 42003 5 1 1 42002
0 42004 7 1 2 21987 95481
0 42005 5 1 1 42004
0 42006 7 1 2 68740 42005
0 42007 5 1 1 42006
0 42008 7 1 2 95726 96412
0 42009 5 1 1 42008
0 42010 7 1 2 42007 42009
0 42011 5 1 1 42010
0 42012 7 1 2 60391 42011
0 42013 5 1 1 42012
0 42014 7 1 2 92958 95472
0 42015 5 1 1 42014
0 42016 7 1 2 42013 42015
0 42017 5 1 1 42016
0 42018 7 4 2 86280 94751
0 42019 7 1 2 42017 96582
0 42020 5 1 1 42019
0 42021 7 1 2 42003 42020
0 42022 7 1 2 41971 42021
0 42023 5 1 1 42022
0 42024 7 1 2 70645 42023
0 42025 5 1 1 42024
0 42026 7 1 2 85858 86246
0 42027 5 1 1 42026
0 42028 7 4 2 68741 42027
0 42029 7 1 2 76446 82655
0 42030 5 1 1 42029
0 42031 7 1 2 39716 42030
0 42032 5 1 1 42031
0 42033 7 1 2 96586 42032
0 42034 5 1 1 42033
0 42035 7 2 2 61117 76930
0 42036 7 1 2 96554 96590
0 42037 5 1 1 42036
0 42038 7 1 2 42034 42037
0 42039 5 1 1 42038
0 42040 7 1 2 64029 42039
0 42041 5 1 1 42040
0 42042 7 1 2 66884 96549
0 42043 7 1 2 90472 42042
0 42044 5 1 1 42043
0 42045 7 1 2 42041 42044
0 42046 5 1 1 42045
0 42047 7 1 2 68458 42046
0 42048 5 1 1 42047
0 42049 7 1 2 84503 86107
0 42050 5 2 1 42049
0 42051 7 1 2 96551 96592
0 42052 5 1 1 42051
0 42053 7 1 2 59612 42052
0 42054 5 1 1 42053
0 42055 7 1 2 64326 87346
0 42056 5 1 1 42055
0 42057 7 1 2 86122 87347
0 42058 5 2 1 42057
0 42059 7 1 2 84504 96594
0 42060 7 1 2 42056 42059
0 42061 5 1 1 42060
0 42062 7 1 2 59387 87073
0 42063 7 1 2 96568 42062
0 42064 5 1 1 42063
0 42065 7 1 2 96593 42064
0 42066 5 1 1 42065
0 42067 7 1 2 69431 42066
0 42068 5 1 1 42067
0 42069 7 1 2 70290 87074
0 42070 7 1 2 96569 42069
0 42071 5 1 1 42070
0 42072 7 1 2 42068 42071
0 42073 7 1 2 42061 42072
0 42074 7 1 2 42054 42073
0 42075 5 1 1 42074
0 42076 7 1 2 61118 42075
0 42077 5 1 1 42076
0 42078 7 2 2 87863 95715
0 42079 7 1 2 59613 92457
0 42080 7 1 2 96596 42079
0 42081 5 1 1 42080
0 42082 7 1 2 42077 42081
0 42083 5 1 1 42082
0 42084 7 1 2 75345 42083
0 42085 5 1 1 42084
0 42086 7 1 2 42048 42085
0 42087 5 1 1 42086
0 42088 7 1 2 68991 42087
0 42089 5 1 1 42088
0 42090 7 5 2 90199 94752
0 42091 5 2 1 96598
0 42092 7 1 2 86323 95194
0 42093 7 1 2 96599 42092
0 42094 5 1 1 42093
0 42095 7 1 2 42089 42094
0 42096 7 1 2 42025 42095
0 42097 5 1 1 42096
0 42098 7 1 2 60583 42097
0 42099 5 1 1 42098
0 42100 7 1 2 84275 86108
0 42101 5 1 1 42100
0 42102 7 1 2 88087 93630
0 42103 5 1 1 42102
0 42104 7 1 2 42101 42103
0 42105 5 1 1 42104
0 42106 7 1 2 75018 42105
0 42107 5 1 1 42106
0 42108 7 2 2 66741 85346
0 42109 5 4 1 96605
0 42110 7 1 2 7684 96607
0 42111 5 1 1 42110
0 42112 7 1 2 86109 42111
0 42113 5 1 1 42112
0 42114 7 1 2 42107 42113
0 42115 5 1 1 42114
0 42116 7 1 2 60814 42115
0 42117 5 1 1 42116
0 42118 7 2 2 64030 95716
0 42119 5 1 1 96611
0 42120 7 1 2 87348 42119
0 42121 5 2 1 42120
0 42122 7 1 2 84292 96613
0 42123 5 1 1 42122
0 42124 7 3 2 66742 95717
0 42125 7 1 2 93760 96615
0 42126 5 1 1 42125
0 42127 7 1 2 42123 42126
0 42128 7 1 2 42117 42127
0 42129 5 1 1 42128
0 42130 7 1 2 59388 42129
0 42131 5 1 1 42130
0 42132 7 1 2 86196 95999
0 42133 5 1 1 42132
0 42134 7 1 2 59614 96595
0 42135 5 1 1 42134
0 42136 7 1 2 60815 96614
0 42137 5 1 1 42136
0 42138 7 1 2 29849 42137
0 42139 7 1 2 42135 42138
0 42140 5 1 1 42139
0 42141 7 1 2 84293 42140
0 42142 5 1 1 42141
0 42143 7 1 2 42133 42142
0 42144 7 1 2 42131 42143
0 42145 5 1 1 42144
0 42146 7 1 2 85913 42145
0 42147 5 1 1 42146
0 42148 7 1 2 76931 92334
0 42149 5 1 1 42148
0 42150 7 1 2 92802 42149
0 42151 5 1 1 42150
0 42152 7 1 2 81982 84805
0 42153 7 1 2 42151 42152
0 42154 5 1 1 42153
0 42155 7 1 2 42147 42154
0 42156 5 1 1 42155
0 42157 7 1 2 76797 42156
0 42158 5 1 1 42157
0 42159 7 1 2 68459 90473
0 42160 5 1 1 42159
0 42161 7 1 2 74952 42160
0 42162 5 1 1 42161
0 42163 7 4 2 70646 86974
0 42164 7 1 2 60392 96618
0 42165 5 1 1 42164
0 42166 7 1 2 87092 42165
0 42167 5 1 1 42166
0 42168 7 1 2 63801 42167
0 42169 7 1 2 42162 42168
0 42170 5 1 1 42169
0 42171 7 1 2 92830 94397
0 42172 7 1 2 95852 42171
0 42173 7 1 2 76932 42172
0 42174 5 1 1 42173
0 42175 7 1 2 42170 42174
0 42176 5 1 1 42175
0 42177 7 1 2 68905 42176
0 42178 5 1 1 42177
0 42179 7 2 2 64031 96571
0 42180 7 1 2 95853 96622
0 42181 7 1 2 96216 42180
0 42182 5 1 1 42181
0 42183 7 1 2 42178 42182
0 42184 5 1 1 42183
0 42185 7 1 2 68081 42184
0 42186 5 1 1 42185
0 42187 7 1 2 12246 96104
0 42188 5 2 1 42187
0 42189 7 1 2 75019 96624
0 42190 5 1 1 42189
0 42191 7 1 2 61119 95091
0 42192 5 1 1 42191
0 42193 7 1 2 42190 42192
0 42194 5 1 1 42193
0 42195 7 1 2 69582 42194
0 42196 5 1 1 42195
0 42197 7 1 2 69950 89904
0 42198 5 1 1 42197
0 42199 7 1 2 61594 73358
0 42200 5 1 1 42199
0 42201 7 1 2 83204 42200
0 42202 7 1 2 42198 42201
0 42203 5 1 1 42202
0 42204 7 1 2 84294 42203
0 42205 5 1 1 42204
0 42206 7 1 2 42196 42205
0 42207 5 1 1 42206
0 42208 7 1 2 81797 86110
0 42209 7 1 2 42207 42208
0 42210 5 1 1 42209
0 42211 7 1 2 42186 42210
0 42212 7 1 2 42158 42211
0 42213 5 1 1 42212
0 42214 7 1 2 68992 42213
0 42215 5 1 1 42214
0 42216 7 1 2 42099 42215
0 42217 5 1 1 42216
0 42218 7 1 2 67717 42217
0 42219 5 1 1 42218
0 42220 7 1 2 75020 96444
0 42221 5 1 1 42220
0 42222 7 1 2 61120 93769
0 42223 5 1 1 42222
0 42224 7 1 2 42221 42223
0 42225 5 1 1 42224
0 42226 7 1 2 68742 42225
0 42227 5 1 1 42226
0 42228 7 1 2 85291 42227
0 42229 5 1 1 42228
0 42230 7 1 2 61901 42229
0 42231 5 1 1 42230
0 42232 7 3 2 68743 92865
0 42233 5 1 1 96626
0 42234 7 1 2 80878 85914
0 42235 7 1 2 96627 42234
0 42236 5 1 1 42235
0 42237 7 1 2 42231 42236
0 42238 5 1 1 42237
0 42239 7 1 2 64032 42238
0 42240 5 1 1 42239
0 42241 7 2 2 75021 85529
0 42242 5 1 1 96629
0 42243 7 2 2 79661 96630
0 42244 5 1 1 96631
0 42245 7 1 2 86242 95473
0 42246 7 1 2 96632 42245
0 42247 5 1 1 42246
0 42248 7 1 2 42240 42247
0 42249 5 1 1 42248
0 42250 7 1 2 76798 42249
0 42251 5 1 1 42250
0 42252 7 2 2 79662 78777
0 42253 7 1 2 86591 96633
0 42254 5 1 1 42253
0 42255 7 1 2 89340 90215
0 42256 5 1 1 42255
0 42257 7 1 2 42254 42256
0 42258 5 2 1 42257
0 42259 7 1 2 75022 96635
0 42260 5 1 1 42259
0 42261 7 4 2 60584 84286
0 42262 7 1 2 90113 96637
0 42263 5 1 1 42262
0 42264 7 1 2 42260 42263
0 42265 5 1 1 42264
0 42266 7 1 2 81350 42265
0 42267 5 1 1 42266
0 42268 7 2 2 80879 88997
0 42269 7 1 2 67097 86530
0 42270 7 1 2 96641 42269
0 42271 5 1 1 42270
0 42272 7 1 2 66885 42271
0 42273 7 1 2 42267 42272
0 42274 5 1 1 42273
0 42275 7 2 2 90200 92048
0 42276 5 1 1 96643
0 42277 7 1 2 68460 96072
0 42278 5 1 1 42277
0 42279 7 1 2 42276 42278
0 42280 5 1 1 42279
0 42281 7 1 2 65481 42280
0 42282 5 1 1 42281
0 42283 7 2 2 66743 90639
0 42284 5 1 1 96645
0 42285 7 1 2 92706 96646
0 42286 5 1 1 42285
0 42287 7 2 2 42282 42286
0 42288 5 1 1 96647
0 42289 7 1 2 75023 42288
0 42290 5 1 1 42289
0 42291 7 1 2 90640 96625
0 42292 5 1 1 42291
0 42293 7 1 2 75515 96076
0 42294 5 1 1 42293
0 42295 7 3 2 68461 90201
0 42296 7 1 2 91396 96649
0 42297 5 1 1 42296
0 42298 7 1 2 42294 42297
0 42299 7 1 2 42292 42298
0 42300 5 1 1 42299
0 42301 7 1 2 64033 42300
0 42302 5 1 1 42301
0 42303 7 1 2 61902 42302
0 42304 7 1 2 42290 42303
0 42305 5 1 1 42304
0 42306 7 1 2 42274 42305
0 42307 5 1 1 42306
0 42308 7 1 2 42251 42307
0 42309 5 1 1 42308
0 42310 7 1 2 68082 42309
0 42311 5 1 1 42310
0 42312 7 2 2 67098 87036
0 42313 7 1 2 87864 88998
0 42314 7 1 2 96652 42313
0 42315 7 1 2 95835 42314
0 42316 5 1 1 42315
0 42317 7 1 2 76799 96597
0 42318 7 1 2 96642 42317
0 42319 5 1 1 42318
0 42320 7 1 2 42316 42319
0 42321 7 1 2 42311 42320
0 42322 5 1 1 42321
0 42323 7 1 2 69951 42322
0 42324 5 1 1 42323
0 42325 7 2 2 67099 73482
0 42326 7 1 2 61903 96654
0 42327 5 1 1 42326
0 42328 7 1 2 96117 42327
0 42329 5 2 1 42328
0 42330 7 1 2 95836 96656
0 42331 5 1 1 42330
0 42332 7 1 2 80982 87089
0 42333 5 2 1 42332
0 42334 7 1 2 42331 96658
0 42335 5 1 1 42334
0 42336 7 1 2 79212 42335
0 42337 5 1 1 42336
0 42338 7 2 2 95832 96280
0 42339 7 1 2 74948 96660
0 42340 5 1 1 42339
0 42341 7 1 2 61904 96648
0 42342 5 1 1 42341
0 42343 7 1 2 81351 96636
0 42344 5 1 1 42343
0 42345 7 1 2 86531 96638
0 42346 5 1 1 42345
0 42347 7 1 2 66886 42346
0 42348 7 1 2 42344 42347
0 42349 5 1 1 42348
0 42350 7 1 2 68083 42349
0 42351 7 1 2 42342 42350
0 42352 5 1 1 42351
0 42353 7 1 2 42340 42352
0 42354 5 1 1 42353
0 42355 7 1 2 69583 42354
0 42356 5 1 1 42355
0 42357 7 1 2 84834 96661
0 42358 5 1 1 42357
0 42359 7 1 2 42356 42358
0 42360 5 1 1 42359
0 42361 7 1 2 59615 42360
0 42362 5 1 1 42361
0 42363 7 1 2 42337 42362
0 42364 7 1 2 42324 42363
0 42365 5 1 1 42364
0 42366 7 1 2 68993 42365
0 42367 5 1 1 42366
0 42368 7 1 2 60585 41958
0 42369 5 1 1 42368
0 42370 7 1 2 93655 96300
0 42371 5 1 1 42370
0 42372 7 1 2 42369 42371
0 42373 5 1 1 42372
0 42374 7 1 2 89131 42373
0 42375 5 1 1 42374
0 42376 7 2 2 80880 87301
0 42377 5 1 1 96662
0 42378 7 1 2 42375 42377
0 42379 5 1 1 42378
0 42380 7 1 2 59616 42379
0 42381 5 1 1 42380
0 42382 7 1 2 80881 96657
0 42383 5 1 1 42382
0 42384 7 1 2 96659 42383
0 42385 7 1 2 42381 42384
0 42386 5 1 1 42385
0 42387 7 1 2 63802 42386
0 42388 5 1 1 42387
0 42389 7 4 2 69584 83059
0 42390 5 1 1 96664
0 42391 7 1 2 96623 96665
0 42392 7 1 2 96445 42391
0 42393 5 1 1 42392
0 42394 7 1 2 42388 42393
0 42395 5 1 1 42394
0 42396 7 1 2 68994 42395
0 42397 5 1 1 42396
0 42398 7 6 2 83748 94714
0 42399 7 2 2 96219 96668
0 42400 7 1 2 88137 96674
0 42401 5 1 1 42400
0 42402 7 1 2 42397 42401
0 42403 5 1 1 42402
0 42404 7 1 2 76800 42403
0 42405 5 1 1 42404
0 42406 7 1 2 96415 96675
0 42407 5 1 1 42406
0 42408 7 1 2 69952 73469
0 42409 7 1 2 92006 42408
0 42410 7 6 2 68744 94753
0 42411 7 2 2 61595 86281
0 42412 7 1 2 96676 96682
0 42413 7 1 2 42409 42412
0 42414 5 1 1 42413
0 42415 7 1 2 42407 42414
0 42416 7 1 2 42405 42415
0 42417 7 1 2 42367 42416
0 42418 7 1 2 42219 42417
0 42419 5 1 1 42418
0 42420 7 1 2 60698 42419
0 42421 5 1 1 42420
0 42422 7 1 2 89321 96209
0 42423 5 1 1 42422
0 42424 7 1 2 75346 91423
0 42425 5 1 1 42424
0 42426 7 1 2 42423 42425
0 42427 5 1 1 42426
0 42428 7 1 2 85530 42427
0 42429 5 1 1 42428
0 42430 7 2 2 88141 94158
0 42431 7 5 2 63533 96684
0 42432 5 1 1 96686
0 42433 7 2 2 68462 92856
0 42434 7 2 2 74802 96691
0 42435 7 1 2 62735 96693
0 42436 5 1 1 42435
0 42437 7 1 2 42432 42436
0 42438 5 1 1 42437
0 42439 7 1 2 68084 42438
0 42440 5 1 1 42439
0 42441 7 1 2 92878 96694
0 42442 5 1 1 42441
0 42443 7 1 2 42440 42442
0 42444 5 1 1 42443
0 42445 7 1 2 59617 42444
0 42446 5 1 1 42445
0 42447 7 1 2 96012 96687
0 42448 5 1 1 42447
0 42449 7 1 2 80322 91767
0 42450 5 1 1 42449
0 42451 7 1 2 81193 82619
0 42452 5 1 1 42451
0 42453 7 1 2 42450 42452
0 42454 5 1 1 42453
0 42455 7 1 2 89044 42454
0 42456 5 1 1 42455
0 42457 7 1 2 76086 73194
0 42458 7 1 2 87368 42457
0 42459 7 1 2 92857 42458
0 42460 5 1 1 42459
0 42461 7 1 2 42456 42460
0 42462 5 1 1 42461
0 42463 7 1 2 68463 42462
0 42464 5 1 1 42463
0 42465 7 1 2 42448 42464
0 42466 7 1 2 42446 42465
0 42467 5 1 1 42466
0 42468 7 1 2 68906 42467
0 42469 5 1 1 42468
0 42470 7 1 2 60816 96211
0 42471 5 1 1 42470
0 42472 7 1 2 96214 42471
0 42473 5 1 1 42472
0 42474 7 1 2 59389 42473
0 42475 5 1 1 42474
0 42476 7 1 2 70291 93180
0 42477 5 1 1 42476
0 42478 7 1 2 42475 42477
0 42479 5 1 1 42478
0 42480 7 2 2 59618 80882
0 42481 7 1 2 82758 96695
0 42482 7 1 2 42479 42481
0 42483 5 1 1 42482
0 42484 7 1 2 42469 42483
0 42485 5 1 1 42484
0 42486 7 1 2 68745 42485
0 42487 5 1 1 42486
0 42488 7 1 2 42429 42487
0 42489 5 1 1 42488
0 42490 7 1 2 86795 42489
0 42491 5 1 1 42490
0 42492 7 1 2 81127 96495
0 42493 5 2 1 42492
0 42494 7 1 2 71293 95245
0 42495 5 1 1 42494
0 42496 7 1 2 96372 42495
0 42497 5 1 1 42496
0 42498 7 1 2 96697 42497
0 42499 5 1 1 42498
0 42500 7 1 2 69953 96504
0 42501 5 1 1 42500
0 42502 7 1 2 93035 96488
0 42503 5 1 1 42502
0 42504 7 1 2 42501 42503
0 42505 7 1 2 42499 42504
0 42506 5 1 1 42505
0 42507 7 1 2 59619 42506
0 42508 5 1 1 42507
0 42509 7 1 2 94406 96483
0 42510 5 1 1 42509
0 42511 7 1 2 91578 96098
0 42512 5 1 1 42511
0 42513 7 1 2 42510 42512
0 42514 5 1 1 42513
0 42515 7 1 2 63126 42514
0 42516 5 1 1 42515
0 42517 7 1 2 82184 86453
0 42518 5 1 1 42517
0 42519 7 1 2 42516 42518
0 42520 5 1 1 42519
0 42521 7 1 2 67100 42520
0 42522 5 1 1 42521
0 42523 7 1 2 42508 42522
0 42524 5 1 1 42523
0 42525 7 1 2 77577 42524
0 42526 5 1 1 42525
0 42527 7 1 2 80692 91579
0 42528 5 1 1 42527
0 42529 7 3 2 75347 81840
0 42530 7 1 2 84806 96699
0 42531 7 1 2 73260 42530
0 42532 5 1 1 42531
0 42533 7 1 2 42528 42532
0 42534 5 1 1 42533
0 42535 7 1 2 67718 42534
0 42536 5 1 1 42535
0 42537 7 1 2 76933 92026
0 42538 5 1 1 42537
0 42539 7 1 2 92691 42538
0 42540 7 1 2 42536 42539
0 42541 5 1 1 42540
0 42542 7 1 2 68464 42541
0 42543 5 1 1 42542
0 42544 7 1 2 83721 85757
0 42545 5 9 1 42544
0 42546 7 4 2 68085 96702
0 42547 5 1 1 96711
0 42548 7 1 2 79748 96712
0 42549 5 1 1 42548
0 42550 7 2 2 88198 92053
0 42551 5 1 1 96715
0 42552 7 1 2 96591 96716
0 42553 5 1 1 42552
0 42554 7 1 2 4558 42553
0 42555 5 1 1 42554
0 42556 7 1 2 75348 42555
0 42557 5 1 1 42556
0 42558 7 1 2 42549 42557
0 42559 7 1 2 42543 42558
0 42560 5 1 1 42559
0 42561 7 1 2 63803 42560
0 42562 5 1 1 42561
0 42563 7 1 2 42526 42562
0 42564 5 1 1 42563
0 42565 7 1 2 86758 42564
0 42566 5 1 1 42565
0 42567 7 2 2 89322 92837
0 42568 5 1 1 96717
0 42569 7 1 2 73483 96718
0 42570 5 1 1 42569
0 42571 7 1 2 87184 92668
0 42572 7 1 2 96688 42571
0 42573 5 1 1 42572
0 42574 7 1 2 42570 42573
0 42575 5 1 1 42574
0 42576 7 1 2 67719 42575
0 42577 5 1 1 42576
0 42578 7 2 2 60699 86258
0 42579 7 1 2 91412 90114
0 42580 7 1 2 96719 42579
0 42581 5 1 1 42580
0 42582 7 1 2 42577 42581
0 42583 5 1 1 42582
0 42584 7 1 2 61121 42583
0 42585 5 1 1 42584
0 42586 7 2 2 78200 86474
0 42587 7 1 2 61760 85803
0 42588 7 1 2 87018 42587
0 42589 7 1 2 96721 42588
0 42590 5 1 1 42589
0 42591 7 1 2 42585 42590
0 42592 5 1 1 42591
0 42593 7 1 2 70989 42592
0 42594 5 1 1 42593
0 42595 7 5 2 68907 86975
0 42596 7 1 2 90125 92582
0 42597 7 1 2 96723 42596
0 42598 7 1 2 96456 42597
0 42599 7 1 2 73261 42598
0 42600 5 1 1 42599
0 42601 7 1 2 42594 42600
0 42602 7 1 2 42566 42601
0 42603 7 1 2 42491 42602
0 42604 5 1 1 42603
0 42605 7 1 2 68995 42604
0 42606 5 1 1 42605
0 42607 7 1 2 96402 41488
0 42608 5 1 1 42607
0 42609 7 1 2 89938 95920
0 42610 7 1 2 42608 42609
0 42611 5 1 1 42610
0 42612 7 1 2 42606 42611
0 42613 5 1 1 42612
0 42614 7 1 2 70202 42613
0 42615 5 1 1 42614
0 42616 7 9 2 65611 68996
0 42617 7 2 2 87909 91546
0 42618 7 1 2 92478 96737
0 42619 5 1 1 42618
0 42620 7 1 2 85544 42619
0 42621 5 1 1 42620
0 42622 7 1 2 75349 42621
0 42623 5 1 1 42622
0 42624 7 1 2 70647 85531
0 42625 5 1 1 42624
0 42626 7 1 2 89836 96738
0 42627 5 1 1 42626
0 42628 7 1 2 42625 42627
0 42629 7 1 2 42623 42628
0 42630 5 1 1 42629
0 42631 7 1 2 80883 42630
0 42632 5 1 1 42631
0 42633 7 2 2 68908 71397
0 42634 7 1 2 74684 91823
0 42635 7 1 2 96739 42634
0 42636 5 1 1 42635
0 42637 7 1 2 42632 42636
0 42638 5 1 1 42637
0 42639 7 1 2 86324 42638
0 42640 5 1 1 42639
0 42641 7 2 2 68465 83494
0 42642 7 1 2 70464 96741
0 42643 5 1 1 42642
0 42644 7 1 2 90075 42643
0 42645 5 1 1 42644
0 42646 7 1 2 79663 42645
0 42647 5 1 1 42646
0 42648 7 1 2 68466 70465
0 42649 5 1 1 42648
0 42650 7 1 2 90762 42649
0 42651 5 1 1 42650
0 42652 7 1 2 80884 42651
0 42653 5 1 1 42652
0 42654 7 1 2 42647 42653
0 42655 5 1 1 42654
0 42656 7 1 2 79715 42655
0 42657 5 1 1 42656
0 42658 7 1 2 79275 80371
0 42659 5 2 1 42658
0 42660 7 1 2 76801 96743
0 42661 5 1 1 42660
0 42662 7 1 2 80347 42284
0 42663 5 1 1 42662
0 42664 7 1 2 61596 42663
0 42665 5 1 1 42664
0 42666 7 1 2 42661 42665
0 42667 5 1 1 42666
0 42668 7 1 2 86213 42667
0 42669 5 1 1 42668
0 42670 7 1 2 86243 96416
0 42671 5 1 1 42670
0 42672 7 1 2 42669 42671
0 42673 5 1 1 42672
0 42674 7 1 2 68746 76060
0 42675 7 1 2 42673 42674
0 42676 5 1 1 42675
0 42677 7 1 2 42657 42676
0 42678 5 1 1 42677
0 42679 7 1 2 67720 42678
0 42680 5 1 1 42679
0 42681 7 1 2 80906 95922
0 42682 5 1 1 42681
0 42683 7 2 2 96634 42682
0 42684 7 1 2 61905 73289
0 42685 7 1 2 96745 42684
0 42686 5 1 1 42685
0 42687 7 1 2 42680 42686
0 42688 5 1 1 42687
0 42689 7 1 2 61122 42688
0 42690 5 1 1 42689
0 42691 7 1 2 61906 96406
0 42692 7 1 2 96746 42691
0 42693 5 1 1 42692
0 42694 7 1 2 42690 42693
0 42695 5 1 1 42694
0 42696 7 1 2 68909 42695
0 42697 5 1 1 42696
0 42698 7 1 2 82617 95977
0 42699 5 1 1 42698
0 42700 7 1 2 68467 96236
0 42701 5 1 1 42700
0 42702 7 1 2 42699 42701
0 42703 5 1 1 42702
0 42704 7 1 2 90641 42703
0 42705 5 1 1 42704
0 42706 7 1 2 89557 92762
0 42707 5 1 1 42706
0 42708 7 1 2 81596 85143
0 42709 7 1 2 71407 42708
0 42710 5 1 1 42709
0 42711 7 1 2 42707 42710
0 42712 7 1 2 42705 42711
0 42713 5 1 1 42712
0 42714 7 1 2 59390 42713
0 42715 5 1 1 42714
0 42716 7 1 2 88262 95535
0 42717 5 1 1 42716
0 42718 7 1 2 78778 73918
0 42719 7 1 2 90133 42718
0 42720 5 1 1 42719
0 42721 7 1 2 42717 42720
0 42722 7 1 2 42715 42721
0 42723 5 1 1 42722
0 42724 7 1 2 86592 42723
0 42725 5 1 1 42724
0 42726 7 2 2 83555 96744
0 42727 7 1 2 76589 96747
0 42728 5 1 1 42727
0 42729 7 1 2 62736 76434
0 42730 5 1 1 42729
0 42731 7 1 2 78779 89303
0 42732 7 1 2 42730 42731
0 42733 5 1 1 42732
0 42734 7 1 2 42728 42733
0 42735 5 1 1 42734
0 42736 7 1 2 86593 42735
0 42737 5 1 1 42736
0 42738 7 1 2 76590 90143
0 42739 7 1 2 96644 42738
0 42740 5 1 1 42739
0 42741 7 1 2 42737 42740
0 42742 5 1 1 42741
0 42743 7 1 2 76802 42742
0 42744 5 1 1 42743
0 42745 7 1 2 83376 90055
0 42746 7 1 2 96252 42745
0 42747 5 1 1 42746
0 42748 7 1 2 42744 42747
0 42749 7 1 2 42725 42748
0 42750 5 1 1 42749
0 42751 7 1 2 61907 42750
0 42752 5 1 1 42751
0 42753 7 1 2 68747 76591
0 42754 7 2 2 93028 42753
0 42755 7 1 2 86983 96740
0 42756 7 1 2 96749 42755
0 42757 5 1 1 42756
0 42758 7 1 2 42752 42757
0 42759 5 1 1 42758
0 42760 7 1 2 69432 42759
0 42761 5 1 1 42760
0 42762 7 1 2 60817 89804
0 42763 5 1 1 42762
0 42764 7 1 2 95624 96742
0 42765 5 1 1 42764
0 42766 7 1 2 42763 42765
0 42767 5 1 1 42766
0 42768 7 1 2 81760 96572
0 42769 7 1 2 42767 42768
0 42770 5 1 1 42769
0 42771 7 1 2 42761 42770
0 42772 7 1 2 42697 42771
0 42773 5 1 1 42772
0 42774 7 1 2 68086 42773
0 42775 5 1 1 42774
0 42776 7 1 2 42640 42775
0 42777 5 1 1 42776
0 42778 7 1 2 96728 42777
0 42779 5 1 1 42778
0 42780 7 1 2 42615 42779
0 42781 7 1 2 42421 42780
0 42782 5 1 1 42781
0 42783 7 1 2 76999 42782
0 42784 5 1 1 42783
0 42785 7 2 2 68087 77000
0 42786 5 2 1 96751
0 42787 7 1 2 74803 85532
0 42788 5 1 1 42787
0 42789 7 1 2 92080 42788
0 42790 5 1 1 42789
0 42791 7 1 2 96752 42790
0 42792 5 1 1 42791
0 42793 7 1 2 68748 83603
0 42794 7 1 2 81721 42793
0 42795 7 1 2 94012 42794
0 42796 5 1 1 42795
0 42797 7 1 2 42792 42796
0 42798 5 1 1 42797
0 42799 7 1 2 59620 42798
0 42800 5 1 1 42799
0 42801 7 1 2 69585 83995
0 42802 5 1 1 42801
0 42803 7 2 2 91539 42802
0 42804 5 1 1 96755
0 42805 7 1 2 68088 42804
0 42806 5 2 1 42805
0 42807 7 1 2 80039 96757
0 42808 5 1 1 42807
0 42809 7 1 2 85533 42808
0 42810 5 1 1 42809
0 42811 7 1 2 42800 42810
0 42812 5 1 1 42811
0 42813 7 1 2 60586 42812
0 42814 5 1 1 42813
0 42815 7 1 2 76061 95870
0 42816 5 1 1 42815
0 42817 7 1 2 66572 42816
0 42818 5 1 1 42817
0 42819 7 2 2 63534 42818
0 42820 5 1 1 96759
0 42821 7 1 2 89342 96760
0 42822 5 1 1 42821
0 42823 7 1 2 74804 96206
0 42824 5 1 1 42823
0 42825 7 3 2 59391 71425
0 42826 5 1 1 96761
0 42827 7 1 2 69433 91151
0 42828 7 1 2 96762 42827
0 42829 5 1 1 42828
0 42830 7 1 2 42824 42829
0 42831 7 1 2 42822 42830
0 42832 5 1 1 42831
0 42833 7 1 2 67360 42832
0 42834 5 1 1 42833
0 42835 7 1 2 59955 96207
0 42836 5 1 1 42835
0 42837 7 1 2 42834 42836
0 42838 5 1 1 42837
0 42839 7 1 2 92669 42838
0 42840 5 1 1 42839
0 42841 7 1 2 42814 42840
0 42842 5 1 1 42841
0 42843 7 1 2 61761 42842
0 42844 5 1 1 42843
0 42845 7 1 2 68089 42826
0 42846 5 1 1 42845
0 42847 7 1 2 69434 95493
0 42848 7 1 2 42846 42847
0 42849 5 1 1 42848
0 42850 7 1 2 95670 42849
0 42851 7 1 2 42820 42850
0 42852 5 1 1 42851
0 42853 7 1 2 67361 42852
0 42854 5 1 1 42853
0 42855 7 1 2 92710 42854
0 42856 5 1 1 42855
0 42857 7 1 2 80364 92670
0 42858 7 1 2 42856 42857
0 42859 5 1 1 42858
0 42860 7 1 2 42844 42859
0 42861 5 1 1 42860
0 42862 7 1 2 76803 42861
0 42863 5 1 1 42862
0 42864 7 1 2 76347 83610
0 42865 5 1 1 42864
0 42866 7 1 2 96753 42865
0 42867 5 1 1 42866
0 42868 7 1 2 42867 96306
0 42869 5 1 1 42868
0 42870 7 1 2 85545 42869
0 42871 5 1 1 42870
0 42872 7 1 2 61762 42871
0 42873 5 1 1 42872
0 42874 7 1 2 81309 93776
0 42875 5 1 1 42874
0 42876 7 1 2 42873 42875
0 42877 5 1 1 42876
0 42878 7 1 2 60587 42877
0 42879 5 1 1 42878
0 42880 7 1 2 80040 89858
0 42881 7 1 2 92671 42880
0 42882 5 1 1 42881
0 42883 7 1 2 42879 42882
0 42884 5 1 1 42883
0 42885 7 1 2 81352 42884
0 42886 5 1 1 42885
0 42887 7 1 2 42863 42886
0 42888 7 1 2 77001 95981
0 42889 5 1 1 42888
0 42890 7 2 2 69195 84168
0 42891 7 1 2 83556 96764
0 42892 5 1 1 42891
0 42893 7 1 2 42889 42892
0 42894 5 1 1 42893
0 42895 7 1 2 90642 42894
0 42896 5 1 1 42895
0 42897 7 3 2 59956 81339
0 42898 7 1 2 80118 90202
0 42899 7 2 2 96766 42898
0 42900 5 1 1 96769
0 42901 7 2 2 77002 96513
0 42902 7 1 2 59392 96771
0 42903 5 1 1 42902
0 42904 7 1 2 42900 42903
0 42905 7 1 2 42896 42904
0 42906 5 1 1 42905
0 42907 7 1 2 76062 42906
0 42908 5 1 1 42907
0 42909 7 1 2 63804 91529
0 42910 7 1 2 95837 42909
0 42911 5 1 1 42910
0 42912 7 1 2 42908 42911
0 42913 5 1 1 42912
0 42914 7 1 2 68910 42913
0 42915 5 1 1 42914
0 42916 7 2 2 91749 92375
0 42917 5 1 1 96773
0 42918 7 1 2 69268 73296
0 42919 5 1 1 42918
0 42920 7 1 2 96774 42919
0 42921 5 1 1 42920
0 42922 7 1 2 42915 42921
0 42923 5 1 1 42922
0 42924 7 1 2 68090 42923
0 42925 5 1 1 42924
0 42926 7 2 2 83557 84685
0 42927 5 1 1 96775
0 42928 7 1 2 96763 96776
0 42929 5 1 1 42928
0 42930 7 1 2 77003 96237
0 42931 5 1 1 42930
0 42932 7 1 2 42929 42931
0 42933 5 1 1 42932
0 42934 7 1 2 68091 42933
0 42935 5 1 1 42934
0 42936 7 1 2 82982 89952
0 42937 5 1 1 42936
0 42938 7 1 2 42935 42937
0 42939 5 1 1 42938
0 42940 7 1 2 90643 42939
0 42941 5 1 1 42940
0 42942 7 1 2 59393 96770
0 42943 5 1 1 42942
0 42944 7 1 2 59621 96772
0 42945 5 1 1 42944
0 42946 7 1 2 42943 42945
0 42947 5 1 1 42946
0 42948 7 1 2 68092 42947
0 42949 5 1 1 42948
0 42950 7 1 2 42941 42949
0 42951 5 1 1 42950
0 42952 7 1 2 68911 42951
0 42953 5 1 1 42952
0 42954 7 7 2 60174 92513
0 42955 7 1 2 92805 93761
0 42956 7 1 2 96777 42955
0 42957 5 1 1 42956
0 42958 7 1 2 42953 42957
0 42959 5 1 1 42958
0 42960 7 1 2 69435 42959
0 42961 5 1 1 42960
0 42962 7 1 2 64802 83607
0 42963 5 2 1 42962
0 42964 7 1 2 63127 84361
0 42965 7 1 2 96784 42964
0 42966 5 1 1 42965
0 42967 7 1 2 84551 42966
0 42968 5 1 1 42967
0 42969 7 1 2 90644 42968
0 42970 5 1 1 42969
0 42971 7 1 2 88189 90203
0 42972 7 1 2 83772 42971
0 42973 5 1 1 42972
0 42974 7 1 2 96515 42973
0 42975 7 1 2 42970 42974
0 42976 5 1 1 42975
0 42977 7 1 2 68912 42976
0 42978 5 1 1 42977
0 42979 7 1 2 42917 42978
0 42980 5 1 1 42979
0 42981 7 1 2 68468 42980
0 42982 5 1 1 42981
0 42983 7 1 2 42961 42982
0 42984 7 1 2 42925 42983
0 42985 5 1 1 42984
0 42986 7 1 2 61597 42985
0 42987 5 1 1 42986
0 42988 7 1 2 59957 72155
0 42989 5 1 1 42988
0 42990 7 1 2 78146 42989
0 42991 5 1 1 42990
0 42992 7 1 2 96689 42991
0 42993 5 1 1 42992
0 42994 7 1 2 76503 93955
0 42995 7 1 2 92858 42994
0 42996 5 1 1 42995
0 42997 7 1 2 42993 42996
0 42998 5 1 1 42997
0 42999 7 1 2 68749 42998
0 43000 5 1 1 42999
0 43001 7 1 2 80815 94441
0 43002 5 1 1 43001
0 43003 7 1 2 92420 43002
0 43004 5 1 1 43003
0 43005 7 1 2 60588 43004
0 43006 5 1 1 43005
0 43007 7 1 2 80816 86624
0 43008 5 1 1 43007
0 43009 7 1 2 43006 43008
0 43010 5 1 1 43009
0 43011 7 1 2 74603 83588
0 43012 7 1 2 43010 43011
0 43013 5 1 1 43012
0 43014 7 1 2 43000 43013
0 43015 5 1 1 43014
0 43016 7 1 2 69954 43015
0 43017 5 1 1 43016
0 43018 7 1 2 63128 83255
0 43019 5 4 1 43018
0 43020 7 1 2 59622 96786
0 43021 5 2 1 43020
0 43022 7 1 2 68093 13823
0 43023 5 1 1 43022
0 43024 7 1 2 96790 43023
0 43025 5 1 1 43024
0 43026 7 1 2 96690 43025
0 43027 5 1 1 43026
0 43028 7 1 2 82983 84037
0 43029 7 1 2 96692 43028
0 43030 5 1 1 43029
0 43031 7 1 2 43027 43030
0 43032 5 1 1 43031
0 43033 7 1 2 68750 43032
0 43034 5 1 1 43033
0 43035 7 1 2 63129 80220
0 43036 5 1 1 43035
0 43037 7 1 2 89453 43036
0 43038 5 1 1 43037
0 43039 7 1 2 71436 80216
0 43040 5 1 1 43039
0 43041 7 1 2 80817 43040
0 43042 7 1 2 96302 43041
0 43043 5 1 1 43042
0 43044 7 1 2 43038 43043
0 43045 5 1 1 43044
0 43046 7 1 2 63805 43045
0 43047 5 1 1 43046
0 43048 7 1 2 43034 43047
0 43049 7 1 2 43017 43048
0 43050 5 1 1 43049
0 43051 7 1 2 68913 43050
0 43052 5 1 1 43051
0 43053 7 6 2 59623 77004
0 43054 5 1 1 96792
0 43055 7 1 2 63130 7321
0 43056 7 1 2 43054 43055
0 43057 5 1 1 43056
0 43058 7 1 2 68469 43057
0 43059 5 1 1 43058
0 43060 7 2 2 75127 89004
0 43061 5 1 1 96798
0 43062 7 1 2 77035 43061
0 43063 5 1 1 43062
0 43064 7 1 2 68470 77005
0 43065 5 1 1 43064
0 43066 7 1 2 78355 84600
0 43067 5 1 1 43066
0 43068 7 1 2 43065 43067
0 43069 5 1 1 43068
0 43070 7 1 2 69955 43069
0 43071 5 1 1 43070
0 43072 7 1 2 43063 43071
0 43073 7 1 2 43059 43072
0 43074 5 1 1 43073
0 43075 7 1 2 95936 43074
0 43076 5 1 1 43075
0 43077 7 1 2 43052 43076
0 43078 5 1 1 43077
0 43079 7 1 2 70203 43078
0 43080 5 1 1 43079
0 43081 7 1 2 42987 43080
0 43082 7 1 2 42887 43081
0 43083 5 1 1 43082
0 43084 7 1 2 61908 43083
0 43085 5 1 1 43084
0 43086 7 1 2 76426 96748
0 43087 5 1 1 43086
0 43088 7 1 2 85292 43087
0 43089 5 1 1 43088
0 43090 7 1 2 76804 43089
0 43091 5 1 1 43090
0 43092 7 1 2 90645 96273
0 43093 5 1 1 43092
0 43094 7 1 2 95684 95994
0 43095 5 1 1 43094
0 43096 7 1 2 96516 43095
0 43097 7 1 2 43093 43096
0 43098 5 1 1 43097
0 43099 7 1 2 61598 43098
0 43100 5 1 1 43099
0 43101 7 1 2 43091 43100
0 43102 5 1 1 43101
0 43103 7 1 2 92523 43102
0 43104 5 1 1 43103
0 43105 7 1 2 90811 90051
0 43106 7 1 2 90216 43105
0 43107 5 1 1 43106
0 43108 7 1 2 43104 43107
0 43109 5 1 1 43108
0 43110 7 1 2 68094 43109
0 43111 5 1 1 43110
0 43112 7 3 2 75516 92104
0 43113 7 1 2 75085 92376
0 43114 7 1 2 96800 43113
0 43115 5 1 1 43114
0 43116 7 1 2 43111 43115
0 43117 5 1 1 43116
0 43118 7 1 2 69436 43117
0 43119 5 1 1 43118
0 43120 7 1 2 95894 96685
0 43121 5 1 1 43120
0 43122 7 2 2 80461 92479
0 43123 5 1 1 96803
0 43124 7 4 2 59624 94174
0 43125 7 1 2 4292 96805
0 43126 7 1 2 96804 43125
0 43127 5 1 1 43126
0 43128 7 1 2 43121 43127
0 43129 5 1 1 43128
0 43130 7 1 2 83558 43129
0 43131 5 1 1 43130
0 43132 7 1 2 76511 73308
0 43133 5 1 1 43132
0 43134 7 1 2 63806 43133
0 43135 7 1 2 91902 43134
0 43136 5 1 1 43135
0 43137 7 1 2 43131 43136
0 43138 5 1 1 43137
0 43139 7 1 2 68095 43138
0 43140 5 1 1 43139
0 43141 7 1 2 70237 83190
0 43142 7 1 2 91812 43141
0 43143 5 1 1 43142
0 43144 7 1 2 43140 43143
0 43145 5 1 1 43144
0 43146 7 1 2 68914 43145
0 43147 5 1 1 43146
0 43148 7 1 2 64803 92915
0 43149 5 1 1 43148
0 43150 7 1 2 70074 84612
0 43151 5 1 1 43150
0 43152 7 1 2 68471 43151
0 43153 7 1 2 43149 43152
0 43154 5 1 1 43153
0 43155 7 1 2 95947 43154
0 43156 5 1 1 43155
0 43157 7 1 2 75517 43156
0 43158 5 1 1 43157
0 43159 7 1 2 75350 83749
0 43160 7 1 2 92214 43159
0 43161 5 1 1 43160
0 43162 7 1 2 43158 43161
0 43163 5 1 1 43162
0 43164 7 1 2 93880 43163
0 43165 5 1 1 43164
0 43166 7 1 2 43147 43165
0 43167 7 1 2 43119 43166
0 43168 5 1 1 43167
0 43169 7 1 2 61909 43168
0 43170 5 1 1 43169
0 43171 7 2 2 85709 87336
0 43172 7 1 2 82783 82503
0 43173 7 1 2 96809 43172
0 43174 7 1 2 90136 43173
0 43175 5 1 1 43174
0 43176 7 1 2 75087 43123
0 43177 5 1 1 43176
0 43178 7 1 2 87337 92783
0 43179 7 1 2 96801 43178
0 43180 7 1 2 43177 43179
0 43181 5 1 1 43180
0 43182 7 1 2 43175 43181
0 43183 7 1 2 43170 43182
0 43184 5 1 1 43183
0 43185 7 1 2 69133 43184
0 43186 5 1 1 43185
0 43187 7 1 2 78298 96791
0 43188 5 1 1 43187
0 43189 7 1 2 69956 43188
0 43190 5 1 1 43189
0 43191 7 1 2 67362 84038
0 43192 5 1 1 43191
0 43193 7 1 2 96754 43192
0 43194 7 1 2 43190 43193
0 43195 5 1 1 43194
0 43196 7 1 2 70204 43195
0 43197 5 1 1 43196
0 43198 7 1 2 69957 74909
0 43199 5 1 1 43198
0 43200 7 1 2 70648 82256
0 43201 5 1 1 43200
0 43202 7 1 2 43199 43201
0 43203 7 1 2 43197 43202
0 43204 5 1 1 43203
0 43205 7 1 2 68472 43204
0 43206 5 1 1 43205
0 43207 7 1 2 71294 93161
0 43208 5 1 1 43207
0 43209 7 1 2 83432 95582
0 43210 5 1 1 43209
0 43211 7 1 2 43208 43210
0 43212 5 1 1 43211
0 43213 7 1 2 82934 43212
0 43214 5 1 1 43213
0 43215 7 1 2 43206 43214
0 43216 5 1 1 43215
0 43217 7 1 2 43216 96028
0 43218 5 1 1 43217
0 43219 7 1 2 43186 43218
0 43220 7 1 2 43085 43219
0 43221 5 1 1 43220
0 43222 7 1 2 96729 43221
0 43223 5 1 1 43222
0 43224 7 1 2 83017 86111
0 43225 5 1 1 43224
0 43226 7 1 2 87270 92924
0 43227 5 1 1 43226
0 43228 7 1 2 43225 43227
0 43229 5 1 1 43228
0 43230 7 1 2 87954 43229
0 43231 5 1 1 43230
0 43232 7 2 2 67363 85534
0 43233 5 1 1 96811
0 43234 7 1 2 61910 84148
0 43235 7 1 2 96812 43234
0 43236 5 1 1 43235
0 43237 7 1 2 43231 43236
0 43238 5 1 1 43237
0 43239 7 1 2 79443 43238
0 43240 5 1 1 43239
0 43241 7 1 2 92555 93975
0 43242 5 1 1 43241
0 43243 7 1 2 77118 86178
0 43244 7 1 2 95990 43243
0 43245 5 1 1 43244
0 43246 7 1 2 43242 43245
0 43247 5 1 1 43246
0 43248 7 1 2 69958 43247
0 43249 5 1 1 43248
0 43250 7 1 2 87318 92560
0 43251 5 2 1 43250
0 43252 7 1 2 33805 96813
0 43253 5 1 1 43252
0 43254 7 1 2 60393 43253
0 43255 5 1 1 43254
0 43256 7 1 2 84382 86179
0 43257 5 1 1 43256
0 43258 7 1 2 96814 43257
0 43259 5 1 1 43258
0 43260 7 1 2 61599 43259
0 43261 5 1 1 43260
0 43262 7 1 2 43255 43261
0 43263 7 1 2 43249 43262
0 43264 5 1 1 43263
0 43265 7 1 2 63535 43264
0 43266 5 1 1 43265
0 43267 7 1 2 66887 88982
0 43268 7 1 2 91785 93839
0 43269 7 1 2 43267 43268
0 43270 5 1 1 43269
0 43271 7 1 2 43266 43270
0 43272 5 1 1 43271
0 43273 7 1 2 68751 43272
0 43274 5 1 1 43273
0 43275 7 1 2 71668 94315
0 43276 5 1 1 43275
0 43277 7 2 2 69727 87302
0 43278 5 1 1 96815
0 43279 7 1 2 93737 94535
0 43280 7 1 2 96816 43279
0 43281 5 1 1 43280
0 43282 7 1 2 43276 43281
0 43283 5 1 1 43282
0 43284 7 1 2 59958 43283
0 43285 5 1 1 43284
0 43286 7 1 2 61911 89250
0 43287 5 1 1 43286
0 43288 7 1 2 43285 43287
0 43289 5 1 1 43288
0 43290 7 1 2 63807 43289
0 43291 5 1 1 43290
0 43292 7 2 2 87289 92547
0 43293 7 1 2 69959 83925
0 43294 7 1 2 96817 43293
0 43295 5 1 1 43294
0 43296 7 1 2 43291 43295
0 43297 7 1 2 43274 43296
0 43298 5 1 1 43297
0 43299 7 1 2 61763 43298
0 43300 5 1 1 43299
0 43301 7 1 2 43240 43300
0 43302 5 1 1 43301
0 43303 7 1 2 72134 43302
0 43304 5 1 1 43303
0 43305 7 1 2 68473 77326
0 43306 5 1 1 43305
0 43307 7 1 2 91637 43306
0 43308 5 1 1 43307
0 43309 7 1 2 84505 43308
0 43310 5 1 1 43309
0 43311 7 1 2 89751 28278
0 43312 5 1 1 43311
0 43313 7 1 2 43310 43312
0 43314 5 1 1 43313
0 43315 7 1 2 92049 43314
0 43316 5 1 1 43315
0 43317 7 1 2 85553 92073
0 43318 5 1 1 43317
0 43319 7 1 2 43316 43318
0 43320 5 1 1 43319
0 43321 7 1 2 60394 43320
0 43322 5 1 1 43321
0 43323 7 1 2 7948 89806
0 43324 5 1 1 43323
0 43325 7 1 2 60395 43324
0 43326 5 1 1 43325
0 43327 7 1 2 81108 83913
0 43328 5 1 1 43327
0 43329 7 1 2 43326 43328
0 43330 5 1 1 43329
0 43331 7 1 2 77578 43330
0 43332 5 1 1 43331
0 43333 7 1 2 79637 86532
0 43334 7 1 2 76522 43333
0 43335 5 1 1 43334
0 43336 7 1 2 43332 43335
0 43337 5 1 1 43336
0 43338 7 1 2 74604 43337
0 43339 5 1 1 43338
0 43340 7 2 2 81993 77579
0 43341 5 2 1 96819
0 43342 7 1 2 80175 85535
0 43343 5 1 1 43342
0 43344 7 1 2 96821 43343
0 43345 5 1 1 43344
0 43346 7 1 2 84383 43345
0 43347 5 1 1 43346
0 43348 7 1 2 43339 43347
0 43349 7 1 2 43322 43348
0 43350 5 1 1 43349
0 43351 7 1 2 61912 43350
0 43352 5 1 1 43351
0 43353 7 3 2 63131 74074
0 43354 5 1 1 96823
0 43355 7 2 2 68752 96132
0 43356 7 1 2 43354 96826
0 43357 5 1 1 43356
0 43358 7 1 2 91947 89746
0 43359 5 1 1 43358
0 43360 7 1 2 43357 43359
0 43361 5 1 1 43360
0 43362 7 1 2 59959 43361
0 43363 5 1 1 43362
0 43364 7 1 2 78377 96827
0 43365 5 1 1 43364
0 43366 7 1 2 43363 43365
0 43367 5 1 1 43366
0 43368 7 1 2 96724 43367
0 43369 5 1 1 43368
0 43370 7 1 2 74605 96308
0 43371 5 1 1 43370
0 43372 7 1 2 80492 85674
0 43373 7 1 2 92518 43372
0 43374 5 1 1 43373
0 43375 7 1 2 43371 43374
0 43376 5 1 1 43375
0 43377 7 1 2 67364 43376
0 43378 5 1 1 43377
0 43379 7 1 2 79797 86180
0 43380 7 1 2 85355 43379
0 43381 5 1 1 43380
0 43382 7 1 2 96148 43381
0 43383 7 1 2 43378 43382
0 43384 5 1 1 43383
0 43385 7 1 2 61764 43384
0 43386 5 1 1 43385
0 43387 7 1 2 85595 92561
0 43388 7 1 2 92217 43387
0 43389 7 1 2 93762 43388
0 43390 5 1 1 43389
0 43391 7 1 2 43386 43390
0 43392 5 1 1 43391
0 43393 7 1 2 71507 43392
0 43394 5 1 1 43393
0 43395 7 1 2 43369 43394
0 43396 7 1 2 43352 43395
0 43397 7 1 2 43304 43396
0 43398 5 1 1 43397
0 43399 7 1 2 70205 43398
0 43400 5 1 1 43399
0 43401 7 1 2 81891 87303
0 43402 5 1 1 43401
0 43403 7 1 2 82589 87271
0 43404 5 1 1 43403
0 43405 7 1 2 43402 43404
0 43406 5 1 1 43405
0 43407 7 1 2 80335 43406
0 43408 5 1 1 43407
0 43409 7 1 2 86123 9695
0 43410 5 5 1 43409
0 43411 7 1 2 68915 83788
0 43412 5 1 1 43411
0 43413 7 2 2 96828 43412
0 43414 7 1 2 70649 96833
0 43415 5 1 1 43414
0 43416 7 1 2 73552 87278
0 43417 5 1 1 43416
0 43418 7 1 2 43415 43417
0 43419 5 1 1 43418
0 43420 7 1 2 85596 43419
0 43421 5 1 1 43420
0 43422 7 2 2 80336 87272
0 43423 5 2 1 96835
0 43424 7 1 2 60818 92628
0 43425 7 1 2 92720 43424
0 43426 7 1 2 96612 43425
0 43427 5 1 1 43426
0 43428 7 1 2 96837 43427
0 43429 5 1 1 43428
0 43430 7 1 2 59394 43429
0 43431 5 1 1 43430
0 43432 7 1 2 60819 96836
0 43433 5 1 1 43432
0 43434 7 1 2 74606 85597
0 43435 7 1 2 87279 43434
0 43436 5 1 1 43435
0 43437 7 1 2 43433 43436
0 43438 7 1 2 43431 43437
0 43439 5 1 1 43438
0 43440 7 1 2 67365 43439
0 43441 5 1 1 43440
0 43442 7 1 2 43421 43441
0 43443 5 1 1 43442
0 43444 7 1 2 61600 43443
0 43445 5 1 1 43444
0 43446 7 1 2 63132 82157
0 43447 5 1 1 43446
0 43448 7 1 2 59625 43447
0 43449 5 2 1 43448
0 43450 7 1 2 88698 96839
0 43451 5 2 1 43450
0 43452 7 9 2 60175 85306
0 43453 7 1 2 86112 96843
0 43454 7 1 2 96841 43453
0 43455 5 1 1 43454
0 43456 7 1 2 96838 43455
0 43457 5 1 1 43456
0 43458 7 1 2 59960 43457
0 43459 5 1 1 43458
0 43460 7 1 2 88890 92537
0 43461 7 1 2 93742 43460
0 43462 5 1 1 43461
0 43463 7 1 2 43459 43462
0 43464 7 1 2 43445 43463
0 43465 5 1 1 43464
0 43466 7 1 2 75351 43465
0 43467 5 1 1 43466
0 43468 7 1 2 43408 43467
0 43469 5 1 1 43468
0 43470 7 1 2 68474 43469
0 43471 5 1 1 43470
0 43472 7 1 2 68916 76512
0 43473 5 1 1 43472
0 43474 7 1 2 96829 43473
0 43475 7 2 2 71337 43474
0 43476 7 1 2 69134 3936
0 43477 7 1 2 94355 43476
0 43478 7 1 2 96852 43477
0 43479 5 1 1 43478
0 43480 7 4 2 59626 86113
0 43481 5 2 1 96854
0 43482 7 2 2 87421 91530
0 43483 5 1 1 96860
0 43484 7 1 2 96858 43483
0 43485 5 1 1 43484
0 43486 7 1 2 71508 43485
0 43487 5 1 1 43486
0 43488 7 1 2 77006 86114
0 43489 5 1 1 43488
0 43490 7 1 2 59627 96861
0 43491 5 1 1 43490
0 43492 7 1 2 43489 43491
0 43493 7 1 2 43487 43492
0 43494 7 2 2 43479 43493
0 43495 5 1 1 96862
0 43496 7 1 2 61601 95854
0 43497 7 1 2 43495 43496
0 43498 5 1 1 43497
0 43499 7 1 2 80185 81128
0 43500 5 1 1 43499
0 43501 7 1 2 70650 43500
0 43502 5 1 1 43501
0 43503 7 2 2 61765 96703
0 43504 5 1 1 96864
0 43505 7 1 2 43502 43504
0 43506 5 1 1 43505
0 43507 7 1 2 96855 43506
0 43508 5 1 1 43507
0 43509 7 3 2 61766 76805
0 43510 7 2 2 80041 96866
0 43511 7 1 2 96853 96869
0 43512 5 1 1 43511
0 43513 7 1 2 43508 43512
0 43514 5 1 1 43513
0 43515 7 1 2 69135 43514
0 43516 5 1 1 43515
0 43517 7 1 2 86181 91531
0 43518 5 1 1 43517
0 43519 7 1 2 96859 43518
0 43520 5 1 1 43519
0 43521 7 1 2 71509 43520
0 43522 5 1 1 43521
0 43523 7 1 2 69196 86115
0 43524 5 1 1 43523
0 43525 7 1 2 68917 74075
0 43526 5 1 1 43525
0 43527 7 1 2 59961 96830
0 43528 7 1 2 43526 43527
0 43529 5 1 1 43528
0 43530 7 1 2 43524 43529
0 43531 7 1 2 43522 43530
0 43532 5 1 1 43531
0 43533 7 1 2 96870 43532
0 43534 5 1 1 43533
0 43535 7 1 2 43516 43534
0 43536 7 1 2 43498 43535
0 43537 5 1 1 43536
0 43538 7 1 2 68096 43537
0 43539 5 1 1 43538
0 43540 7 1 2 80119 96725
0 43541 7 1 2 95678 43540
0 43542 5 1 1 43541
0 43543 7 1 2 43539 43542
0 43544 7 1 2 43471 43543
0 43545 5 1 1 43544
0 43546 7 1 2 68753 43545
0 43547 5 1 1 43546
0 43548 7 2 2 60396 85915
0 43549 5 2 1 96871
0 43550 7 1 2 93719 95498
0 43551 5 1 1 43550
0 43552 7 1 2 96873 43551
0 43553 5 1 1 43552
0 43554 7 1 2 78062 43553
0 43555 5 1 1 43554
0 43556 7 1 2 80057 83722
0 43557 5 10 1 43556
0 43558 7 1 2 79749 89179
0 43559 7 1 2 96875 43558
0 43560 5 1 1 43559
0 43561 7 1 2 43555 43560
0 43562 5 1 1 43561
0 43563 7 1 2 59962 43562
0 43564 5 1 1 43563
0 43565 7 1 2 86644 89743
0 43566 5 1 1 43565
0 43567 7 1 2 67366 92534
0 43568 7 1 2 93965 43567
0 43569 5 1 1 43568
0 43570 7 1 2 43566 43569
0 43571 5 1 1 43570
0 43572 7 1 2 70651 43571
0 43573 5 1 1 43572
0 43574 7 2 2 68918 92629
0 43575 7 1 2 74635 96885
0 43576 7 1 2 96704 43575
0 43577 5 1 1 43576
0 43578 7 1 2 43573 43577
0 43579 7 1 2 43564 43578
0 43580 5 1 1 43579
0 43581 7 1 2 68097 43580
0 43582 5 1 1 43581
0 43583 7 1 2 76806 92426
0 43584 5 1 1 43583
0 43585 7 1 2 78063 92819
0 43586 7 1 2 83495 43585
0 43587 7 1 2 94976 43586
0 43588 5 1 1 43587
0 43589 7 1 2 43584 43588
0 43590 7 1 2 43582 43589
0 43591 5 1 1 43590
0 43592 7 1 2 61913 43591
0 43593 5 1 1 43592
0 43594 7 1 2 85691 86247
0 43595 5 1 1 43594
0 43596 7 1 2 70652 43595
0 43597 5 1 1 43596
0 43598 7 1 2 85849 96705
0 43599 5 1 1 43598
0 43600 7 1 2 43597 43599
0 43601 5 1 1 43600
0 43602 7 1 2 83018 87338
0 43603 7 1 2 43601 43602
0 43604 5 1 1 43603
0 43605 7 1 2 86331 92541
0 43606 7 1 2 71338 43605
0 43607 7 1 2 83496 43606
0 43608 5 1 1 43607
0 43609 7 1 2 43604 43608
0 43610 5 1 1 43609
0 43611 7 1 2 59628 43610
0 43612 5 1 1 43611
0 43613 7 1 2 78064 87290
0 43614 7 1 2 90068 43613
0 43615 5 1 1 43614
0 43616 7 1 2 43612 43615
0 43617 5 1 1 43616
0 43618 7 1 2 69136 43617
0 43619 5 1 1 43618
0 43620 7 1 2 63536 96758
0 43621 5 1 1 43620
0 43622 7 1 2 90069 96726
0 43623 7 1 2 43621 43622
0 43624 5 1 1 43623
0 43625 7 1 2 43619 43624
0 43626 7 1 2 43593 43625
0 43627 5 1 1 43626
0 43628 7 1 2 63808 43627
0 43629 5 1 1 43628
0 43630 7 1 2 43547 43629
0 43631 7 1 2 43400 43630
0 43632 5 1 1 43631
0 43633 7 1 2 68997 43632
0 43634 5 1 1 43633
0 43635 7 1 2 82436 96824
0 43636 5 2 1 43635
0 43637 7 1 2 81994 96887
0 43638 5 1 1 43637
0 43639 7 2 2 70653 79057
0 43640 7 1 2 61602 96889
0 43641 5 1 1 43640
0 43642 7 1 2 43638 43641
0 43643 5 1 1 43642
0 43644 7 1 2 59963 43643
0 43645 5 1 1 43644
0 43646 7 1 2 93462 96890
0 43647 5 1 1 43646
0 43648 7 1 2 43645 43647
0 43649 5 1 1 43648
0 43650 7 1 2 63809 43649
0 43651 5 1 1 43650
0 43652 7 1 2 59964 96842
0 43653 5 1 1 43652
0 43654 7 1 2 14713 43653
0 43655 5 2 1 43654
0 43656 7 1 2 89752 96891
0 43657 5 1 1 43656
0 43658 7 1 2 43651 43657
0 43659 5 1 1 43658
0 43660 7 1 2 61914 43659
0 43661 5 1 1 43660
0 43662 7 1 2 64804 74525
0 43663 5 1 1 43662
0 43664 7 1 2 68098 43663
0 43665 5 1 1 43664
0 43666 7 1 2 63537 43665
0 43667 5 1 1 43666
0 43668 7 1 2 87955 96619
0 43669 7 1 2 43667 43668
0 43670 5 1 1 43669
0 43671 7 1 2 43661 43670
0 43672 5 1 1 43671
0 43673 7 1 2 64034 43672
0 43674 5 1 1 43673
0 43675 7 1 2 84552 42927
0 43676 5 1 1 43675
0 43677 7 1 2 68919 43676
0 43678 5 1 1 43677
0 43679 7 1 2 96892 96820
0 43680 5 1 1 43679
0 43681 7 1 2 43678 43680
0 43682 5 1 1 43681
0 43683 7 1 2 66888 43682
0 43684 5 1 1 43683
0 43685 7 1 2 81722 79716
0 43686 7 1 2 96888 43685
0 43687 5 1 1 43686
0 43688 7 1 2 43684 43687
0 43689 5 1 1 43688
0 43690 7 1 2 95925 43689
0 43691 5 1 1 43690
0 43692 7 1 2 68475 96834
0 43693 5 1 1 43692
0 43694 7 1 2 69137 96856
0 43695 5 1 1 43694
0 43696 7 1 2 96863 43695
0 43697 5 1 1 43696
0 43698 7 1 2 68099 43697
0 43699 5 1 1 43698
0 43700 7 1 2 43693 43699
0 43701 5 1 1 43700
0 43702 7 1 2 84362 43701
0 43703 5 1 1 43702
0 43704 7 1 2 86116 94834
0 43705 5 1 1 43704
0 43706 7 1 2 59629 93142
0 43707 5 1 1 43706
0 43708 7 1 2 96756 43707
0 43709 5 1 1 43708
0 43710 7 1 2 86182 43709
0 43711 5 1 1 43710
0 43712 7 1 2 43705 43711
0 43713 5 1 1 43712
0 43714 7 1 2 68100 43713
0 43715 5 1 1 43714
0 43716 7 1 2 96118 43715
0 43717 5 1 1 43716
0 43718 7 1 2 84506 43717
0 43719 5 1 1 43718
0 43720 7 1 2 43703 43719
0 43721 5 1 1 43720
0 43722 7 1 2 90780 43721
0 43723 5 1 1 43722
0 43724 7 1 2 83019 82562
0 43725 5 1 1 43724
0 43726 7 2 2 91793 43725
0 43727 5 1 1 96893
0 43728 7 1 2 68101 43727
0 43729 5 1 1 43728
0 43730 7 1 2 63538 43729
0 43731 5 1 1 43730
0 43732 7 1 2 90070 93631
0 43733 7 1 2 43731 43732
0 43734 5 1 1 43733
0 43735 7 1 2 43723 43734
0 43736 7 1 2 43691 43735
0 43737 7 1 2 43674 43736
0 43738 5 1 1 43737
0 43739 7 1 2 68998 43738
0 43740 5 1 1 43739
0 43741 7 5 2 68754 68999
0 43742 7 3 2 83106 96895
0 43743 7 1 2 86117 96900
0 43744 5 1 1 43743
0 43745 7 4 2 68476 94715
0 43746 7 3 2 87291 96903
0 43747 7 1 2 67367 96907
0 43748 5 1 1 43747
0 43749 7 5 2 69000 86571
0 43750 5 1 1 96910
0 43751 7 1 2 43748 43750
0 43752 5 1 1 43751
0 43753 7 1 2 61767 92694
0 43754 7 1 2 43752 43753
0 43755 5 1 1 43754
0 43756 7 1 2 43744 43755
0 43757 5 1 1 43756
0 43758 7 1 2 74607 43757
0 43759 5 1 1 43758
0 43760 7 20 2 66889 69001
0 43761 7 1 2 68102 32629
0 43762 5 1 1 43761
0 43763 7 1 2 81904 43762
0 43764 5 1 1 43763
0 43765 7 1 2 95978 43764
0 43766 5 1 1 43765
0 43767 7 1 2 96196 43766
0 43768 5 1 1 43767
0 43769 7 1 2 96915 43768
0 43770 5 1 1 43769
0 43771 7 1 2 61768 80247
0 43772 7 1 2 96908 43771
0 43773 5 1 1 43772
0 43774 7 1 2 43770 43773
0 43775 5 1 1 43774
0 43776 7 1 2 68920 43775
0 43777 5 1 1 43776
0 43778 7 1 2 43759 43777
0 43779 5 1 1 43778
0 43780 7 1 2 75352 43779
0 43781 5 1 1 43780
0 43782 7 2 2 69345 87668
0 43783 7 1 2 68921 73449
0 43784 7 1 2 96935 43783
0 43785 5 1 1 43784
0 43786 7 1 2 86124 43785
0 43787 5 1 1 43786
0 43788 7 1 2 66744 43787
0 43789 5 1 1 43788
0 43790 7 1 2 86625 94879
0 43791 5 1 1 43790
0 43792 7 1 2 43789 43791
0 43793 5 1 1 43792
0 43794 7 1 2 68477 43793
0 43795 5 1 1 43794
0 43796 7 1 2 69972 89403
0 43797 7 1 2 94644 43796
0 43798 5 1 1 43797
0 43799 7 1 2 68755 43798
0 43800 7 1 2 43795 43799
0 43801 5 1 1 43800
0 43802 7 2 2 61603 80818
0 43803 5 1 1 96937
0 43804 7 1 2 66745 43803
0 43805 5 1 1 43804
0 43806 7 1 2 11954 43278
0 43807 5 1 1 43806
0 43808 7 1 2 43805 43807
0 43809 5 1 1 43808
0 43810 7 1 2 69973 87280
0 43811 7 1 2 94442 43810
0 43812 5 1 1 43811
0 43813 7 1 2 63810 43812
0 43814 7 1 2 43809 43813
0 43815 5 1 1 43814
0 43816 7 1 2 69002 43815
0 43817 7 1 2 43801 43816
0 43818 5 1 1 43817
0 43819 7 1 2 94211 96727
0 43820 5 1 1 43819
0 43821 7 6 2 63811 96323
0 43822 7 1 2 73195 96939
0 43823 5 1 1 43822
0 43824 7 1 2 96603 43823
0 43825 5 1 1 43824
0 43826 7 1 2 60397 87292
0 43827 7 1 2 43825 43826
0 43828 5 1 1 43827
0 43829 7 1 2 43820 43828
0 43830 5 1 1 43829
0 43831 7 1 2 85788 43830
0 43832 5 1 1 43831
0 43833 7 2 2 80819 88088
0 43834 7 1 2 87037 96677
0 43835 7 1 2 96945 43834
0 43836 5 1 1 43835
0 43837 7 1 2 43832 43836
0 43838 7 1 2 43818 43837
0 43839 5 1 1 43838
0 43840 7 1 2 59965 43839
0 43841 5 1 1 43840
0 43842 7 1 2 69728 96587
0 43843 5 1 1 43842
0 43844 7 1 2 41935 43843
0 43845 5 1 1 43844
0 43846 7 1 2 68478 43845
0 43847 5 1 1 43846
0 43848 7 1 2 72456 93976
0 43849 7 1 2 92599 43848
0 43850 5 1 1 43849
0 43851 7 1 2 43847 43850
0 43852 5 1 1 43851
0 43853 7 1 2 64035 43852
0 43854 5 1 1 43853
0 43855 7 1 2 68103 92600
0 43856 7 1 2 94645 43855
0 43857 5 1 1 43856
0 43858 7 1 2 43854 43857
0 43859 5 1 1 43858
0 43860 7 1 2 69003 43859
0 43861 5 1 1 43860
0 43862 7 1 2 43841 43861
0 43863 5 1 1 43862
0 43864 7 1 2 72135 43863
0 43865 5 1 1 43864
0 43866 7 1 2 67368 4641
0 43867 5 1 1 43866
0 43868 7 1 2 63133 43867
0 43869 5 1 1 43868
0 43870 7 1 2 96588 43869
0 43871 5 1 1 43870
0 43872 7 1 2 77327 96555
0 43873 5 1 1 43872
0 43874 7 1 2 43871 43873
0 43875 5 1 1 43874
0 43876 7 1 2 64036 43875
0 43877 5 1 1 43876
0 43878 7 1 2 71729 86139
0 43879 7 1 2 96547 43878
0 43880 5 1 1 43879
0 43881 7 1 2 43877 43880
0 43882 5 1 1 43881
0 43883 7 1 2 68479 43882
0 43884 5 1 1 43883
0 43885 7 1 2 81899 73484
0 43886 7 1 2 96556 43885
0 43887 5 1 1 43886
0 43888 7 1 2 43884 43887
0 43889 5 1 1 43888
0 43890 7 1 2 69004 43889
0 43891 5 1 1 43890
0 43892 7 1 2 92948 96583
0 43893 5 1 1 43892
0 43894 7 1 2 91635 96589
0 43895 5 1 1 43894
0 43896 7 1 2 68480 96557
0 43897 5 1 1 43896
0 43898 7 1 2 43895 43897
0 43899 5 1 1 43898
0 43900 7 1 2 96324 43899
0 43901 5 1 1 43900
0 43902 7 6 2 64115 85347
0 43903 7 4 2 86282 96947
0 43904 5 1 1 96953
0 43905 7 1 2 75518 96954
0 43906 5 1 1 43905
0 43907 7 3 2 68481 94212
0 43908 7 2 2 66890 67369
0 43909 7 1 2 94443 96960
0 43910 7 1 2 96957 43909
0 43911 5 1 1 43910
0 43912 7 1 2 43906 43911
0 43913 5 1 1 43912
0 43914 7 1 2 68922 74608
0 43915 7 1 2 43913 43914
0 43916 5 1 1 43915
0 43917 7 1 2 43901 43916
0 43918 5 1 1 43917
0 43919 7 1 2 71510 43918
0 43920 5 1 1 43919
0 43921 7 1 2 43893 43920
0 43922 7 1 2 43891 43921
0 43923 7 1 2 43865 43922
0 43924 7 1 2 43781 43923
0 43925 5 1 1 43924
0 43926 7 1 2 70206 43925
0 43927 5 1 1 43926
0 43928 7 1 2 68756 81892
0 43929 5 1 1 43928
0 43930 7 1 2 63134 43929
0 43931 5 1 1 43930
0 43932 7 1 2 75115 69197
0 43933 7 1 2 81914 43932
0 43934 5 1 1 43933
0 43935 7 1 2 63812 43934
0 43936 5 1 1 43935
0 43937 7 1 2 90071 43936
0 43938 7 1 2 43931 43937
0 43939 5 1 1 43938
0 43940 7 1 2 63135 96894
0 43941 5 1 1 43940
0 43942 7 1 2 89939 95926
0 43943 7 1 2 43941 43942
0 43944 5 1 1 43943
0 43945 7 1 2 43939 43944
0 43946 5 1 1 43945
0 43947 7 1 2 96584 43946
0 43948 5 1 1 43947
0 43949 7 1 2 43927 43948
0 43950 7 1 2 43740 43949
0 43951 5 1 1 43950
0 43952 7 1 2 60589 43951
0 43953 5 1 1 43952
0 43954 7 2 2 70207 82064
0 43955 7 1 2 84363 96962
0 43956 5 1 1 43955
0 43957 7 1 2 78378 91824
0 43958 5 1 1 43957
0 43959 7 1 2 43956 43958
0 43960 5 1 1 43959
0 43961 7 1 2 85916 43960
0 43962 5 1 1 43961
0 43963 7 1 2 85144 88089
0 43964 5 2 1 43963
0 43965 7 1 2 43962 96964
0 43966 5 1 1 43965
0 43967 7 1 2 64037 43966
0 43968 5 1 1 43967
0 43969 7 2 2 81893 84442
0 43970 7 1 2 86619 96966
0 43971 5 1 1 43970
0 43972 7 1 2 61915 43971
0 43973 7 1 2 43968 43972
0 43974 5 1 1 43973
0 43975 7 1 2 92015 92716
0 43976 5 1 1 43975
0 43977 7 1 2 70654 89304
0 43978 5 1 1 43977
0 43979 7 1 2 80907 43978
0 43980 5 1 1 43979
0 43981 7 1 2 96967 43980
0 43982 5 1 1 43981
0 43983 7 1 2 43976 43982
0 43984 5 1 1 43983
0 43985 7 1 2 68923 43984
0 43986 5 1 1 43985
0 43987 7 1 2 86475 89345
0 43988 7 1 2 96963 43987
0 43989 5 1 1 43988
0 43990 7 1 2 66891 43989
0 43991 7 1 2 43986 43990
0 43992 5 1 1 43991
0 43993 7 1 2 60398 43992
0 43994 7 1 2 43974 43993
0 43995 5 1 1 43994
0 43996 7 1 2 80820 94159
0 43997 5 1 1 43996
0 43998 7 1 2 92130 43997
0 43999 5 1 1 43998
0 44000 7 1 2 61916 94080
0 44001 7 1 2 43999 44000
0 44002 5 1 1 44001
0 44003 7 2 2 81310 93421
0 44004 7 1 2 87075 96968
0 44005 5 1 1 44004
0 44006 7 2 2 79717 88094
0 44007 5 1 1 96970
0 44008 7 1 2 44005 44007
0 44009 5 2 1 44008
0 44010 7 1 2 91683 96972
0 44011 5 1 1 44010
0 44012 7 2 2 65482 86976
0 44013 7 1 2 96969 96974
0 44014 5 1 1 44013
0 44015 7 1 2 44011 44014
0 44016 7 1 2 44002 44015
0 44017 5 1 1 44016
0 44018 7 1 2 80252 44017
0 44019 5 1 1 44018
0 44020 7 1 2 82711 86199
0 44021 5 1 1 44020
0 44022 7 1 2 85536 92542
0 44023 7 1 2 94253 44022
0 44024 7 1 2 74327 44023
0 44025 5 1 1 44024
0 44026 7 1 2 44021 44025
0 44027 5 1 1 44026
0 44028 7 1 2 69138 44027
0 44029 5 1 1 44028
0 44030 7 1 2 95092 96818
0 44031 5 1 1 44030
0 44032 7 1 2 61604 96973
0 44033 5 1 1 44032
0 44034 7 1 2 44031 44033
0 44035 7 1 2 44029 44034
0 44036 5 1 1 44035
0 44037 7 1 2 60590 44036
0 44038 5 1 1 44037
0 44039 7 1 2 85692 86989
0 44040 5 1 1 44039
0 44041 7 1 2 70655 44040
0 44042 5 1 1 44041
0 44043 7 1 2 10741 44042
0 44044 5 1 1 44043
0 44045 7 1 2 96545 44044
0 44046 5 1 1 44045
0 44047 7 1 2 86200 92187
0 44048 5 1 1 44047
0 44049 7 1 2 44046 44048
0 44050 5 1 1 44049
0 44051 7 1 2 77007 44050
0 44052 5 1 1 44051
0 44053 7 2 2 68924 79718
0 44054 7 1 2 84169 88696
0 44055 7 1 2 96976 44054
0 44056 7 1 2 96066 44055
0 44057 5 1 1 44056
0 44058 7 1 2 44052 44057
0 44059 7 1 2 44038 44058
0 44060 7 1 2 44019 44059
0 44061 7 1 2 43995 44060
0 44062 5 1 1 44061
0 44063 7 1 2 69005 44062
0 44064 5 1 1 44063
0 44065 7 8 2 64116 92672
0 44066 7 1 2 81995 96243
0 44067 7 1 2 96978 44066
0 44068 7 1 2 81894 44067
0 44069 7 1 2 83497 44068
0 44070 5 1 1 44069
0 44071 7 1 2 44064 44070
0 44072 5 1 1 44071
0 44073 7 1 2 74805 44072
0 44074 5 1 1 44073
0 44075 7 1 2 43953 44074
0 44076 7 1 2 43634 44075
0 44077 5 1 1 44076
0 44078 7 1 2 60700 44077
0 44079 5 1 1 44078
0 44080 7 1 2 43223 44079
0 44081 5 1 1 44080
0 44082 7 1 2 73827 44081
0 44083 5 1 1 44082
0 44084 7 1 2 42784 44083
0 44085 7 1 2 41905 44084
0 44086 7 1 2 40922 44085
0 44087 7 1 2 39458 44086
0 44088 5 1 1 44087
0 44089 7 1 2 95329 44088
0 44090 5 1 1 44089
0 44091 7 8 2 61769 91684
0 44092 5 1 1 96986
0 44093 7 1 2 87185 96987
0 44094 5 2 1 44093
0 44095 7 1 2 86214 92312
0 44096 5 2 1 44095
0 44097 7 1 2 86408 87133
0 44098 5 2 1 44097
0 44099 7 3 2 60591 96998
0 44100 5 1 1 97000
0 44101 7 1 2 75519 97001
0 44102 5 1 1 44101
0 44103 7 2 2 96996 44102
0 44104 5 1 1 97003
0 44105 7 1 2 96994 97004
0 44106 5 1 1 44105
0 44107 7 5 2 64117 44106
0 44108 7 7 2 63813 95287
0 44109 7 1 2 97005 97010
0 44110 5 2 1 44109
0 44111 7 2 2 68482 96896
0 44112 7 3 2 95251 97019
0 44113 7 2 2 61770 97021
0 44114 7 3 2 90174 95331
0 44115 7 1 2 97024 97026
0 44116 5 1 1 44115
0 44117 7 1 2 97017 44116
0 44118 5 4 1 44117
0 44119 7 1 2 70838 91076
0 44120 5 2 1 44119
0 44121 7 1 2 72242 91650
0 44122 7 1 2 97033 44121
0 44123 5 1 1 44122
0 44124 7 1 2 89527 44123
0 44125 5 1 1 44124
0 44126 7 1 2 97029 44125
0 44127 5 1 1 44126
0 44128 7 2 2 76911 87435
0 44129 5 1 1 97035
0 44130 7 2 2 85434 97036
0 44131 5 1 1 97037
0 44132 7 2 2 74031 90270
0 44133 5 2 1 97039
0 44134 7 1 2 89381 89066
0 44135 5 1 1 44134
0 44136 7 1 2 97041 44135
0 44137 5 1 1 44136
0 44138 7 1 2 64805 44137
0 44139 5 1 1 44138
0 44140 7 1 2 90822 44139
0 44141 5 1 1 44140
0 44142 7 1 2 65022 44141
0 44143 5 1 1 44142
0 44144 7 1 2 72848 74032
0 44145 5 1 1 44144
0 44146 7 1 2 83338 76731
0 44147 7 1 2 44145 44146
0 44148 5 1 1 44147
0 44149 7 1 2 64806 44148
0 44150 5 1 1 44149
0 44151 7 1 2 80092 77096
0 44152 5 1 1 44151
0 44153 7 1 2 76870 90223
0 44154 5 1 1 44153
0 44155 7 1 2 65023 82506
0 44156 5 1 1 44155
0 44157 7 1 2 44154 44156
0 44158 7 1 2 44152 44157
0 44159 7 1 2 44150 44158
0 44160 5 1 1 44159
0 44161 7 1 2 66339 44160
0 44162 5 1 1 44161
0 44163 7 1 2 44143 44162
0 44164 5 1 1 44163
0 44165 7 1 2 66066 44164
0 44166 5 1 1 44165
0 44167 7 1 2 60176 77364
0 44168 5 1 1 44167
0 44169 7 1 2 66340 44168
0 44170 5 1 1 44169
0 44171 7 1 2 4639 73385
0 44172 5 1 1 44171
0 44173 7 1 2 69698 44172
0 44174 5 1 1 44173
0 44175 7 1 2 44170 44174
0 44176 5 1 1 44175
0 44177 7 1 2 87030 44176
0 44178 5 1 1 44177
0 44179 7 1 2 65024 93146
0 44180 5 1 1 44179
0 44181 7 1 2 44178 44180
0 44182 5 1 1 44181
0 44183 7 1 2 72364 44182
0 44184 5 1 1 44183
0 44185 7 1 2 65025 72171
0 44186 5 1 1 44185
0 44187 7 1 2 67721 44186
0 44188 5 1 1 44187
0 44189 7 1 2 81638 78541
0 44190 5 1 1 44189
0 44191 7 1 2 62376 87326
0 44192 5 1 1 44191
0 44193 7 1 2 60177 44192
0 44194 5 1 1 44193
0 44195 7 1 2 44190 44194
0 44196 7 1 2 44188 44195
0 44197 5 1 1 44196
0 44198 7 2 2 65895 74033
0 44199 7 1 2 73134 73450
0 44200 5 1 1 44199
0 44201 7 1 2 97043 44200
0 44202 5 1 1 44201
0 44203 7 1 2 2687 44202
0 44204 7 1 2 90274 44203
0 44205 7 1 2 96408 44204
0 44206 5 1 1 44205
0 44207 7 1 2 70075 44206
0 44208 5 1 1 44207
0 44209 7 1 2 44197 44208
0 44210 7 1 2 44184 44209
0 44211 7 1 2 44166 44210
0 44212 5 1 1 44211
0 44213 7 1 2 63136 44212
0 44214 5 1 1 44213
0 44215 7 1 2 88426 89169
0 44216 5 2 1 44215
0 44217 7 1 2 71828 97045
0 44218 5 1 1 44217
0 44219 7 2 2 62737 78668
0 44220 7 1 2 69860 97047
0 44221 5 1 1 44220
0 44222 7 1 2 44218 44221
0 44223 5 1 1 44222
0 44224 7 1 2 65026 44223
0 44225 5 1 1 44224
0 44226 7 1 2 80480 81690
0 44227 5 1 1 44226
0 44228 7 1 2 44225 44227
0 44229 5 1 1 44228
0 44230 7 1 2 62377 44229
0 44231 5 1 1 44230
0 44232 7 1 2 77164 88763
0 44233 5 1 1 44232
0 44234 7 1 2 44231 44233
0 44235 5 1 1 44234
0 44236 7 1 2 79591 44235
0 44237 5 1 1 44236
0 44238 7 1 2 66067 81461
0 44239 5 1 1 44238
0 44240 7 1 2 65739 73115
0 44241 5 1 1 44240
0 44242 7 1 2 44239 44241
0 44243 5 1 1 44242
0 44244 7 1 2 64807 44243
0 44245 5 1 1 44244
0 44246 7 1 2 87785 95174
0 44247 5 1 1 44246
0 44248 7 1 2 82067 76981
0 44249 5 1 1 44248
0 44250 7 1 2 69139 44249
0 44251 5 1 1 44250
0 44252 7 1 2 64327 44251
0 44253 5 1 1 44252
0 44254 7 1 2 44247 44253
0 44255 7 1 2 44245 44254
0 44256 5 1 1 44255
0 44257 7 1 2 88416 44256
0 44258 5 1 1 44257
0 44259 7 1 2 86401 94667
0 44260 5 1 1 44259
0 44261 7 1 2 44258 44260
0 44262 5 1 1 44261
0 44263 7 1 2 70076 44262
0 44264 5 1 1 44263
0 44265 7 1 2 77710 86960
0 44266 5 1 1 44265
0 44267 7 1 2 65027 44266
0 44268 5 1 1 44267
0 44269 7 1 2 18659 44268
0 44270 5 1 1 44269
0 44271 7 1 2 62738 92679
0 44272 5 1 1 44271
0 44273 7 1 2 84053 44272
0 44274 5 1 1 44273
0 44275 7 1 2 67722 3572
0 44276 5 1 1 44275
0 44277 7 1 2 44274 44276
0 44278 7 1 2 44270 44277
0 44279 5 1 1 44278
0 44280 7 2 2 73880 87436
0 44281 5 1 1 97049
0 44282 7 1 2 80656 44281
0 44283 5 1 1 44282
0 44284 7 1 2 81414 83877
0 44285 7 1 2 94116 44284
0 44286 5 1 1 44285
0 44287 7 1 2 95380 44286
0 44288 7 1 2 44283 44287
0 44289 5 1 1 44288
0 44290 7 1 2 44279 44289
0 44291 7 1 2 44264 44290
0 44292 7 1 2 44237 44291
0 44293 7 1 2 44214 44292
0 44294 5 1 1 44293
0 44295 7 1 2 66573 44294
0 44296 5 1 1 44295
0 44297 7 1 2 44131 44296
0 44298 5 1 1 44297
0 44299 7 1 2 65278 44298
0 44300 5 1 1 44299
0 44301 7 2 2 70208 83818
0 44302 5 1 1 97051
0 44303 7 1 2 70839 44302
0 44304 5 1 1 44303
0 44305 7 1 2 71123 91060
0 44306 5 1 1 44305
0 44307 7 1 2 44304 44306
0 44308 5 1 1 44307
0 44309 7 1 2 69699 44308
0 44310 5 1 1 44309
0 44311 7 1 2 88182 44310
0 44312 5 1 1 44311
0 44313 7 1 2 63137 44312
0 44314 5 1 1 44313
0 44315 7 1 2 77165 81646
0 44316 5 1 1 44315
0 44317 7 1 2 84927 91334
0 44318 5 1 1 44317
0 44319 7 1 2 44316 44318
0 44320 7 1 2 44314 44319
0 44321 5 1 1 44320
0 44322 7 1 2 64567 44321
0 44323 5 1 1 44322
0 44324 7 1 2 88495 95686
0 44325 5 1 1 44324
0 44326 7 1 2 89385 88472
0 44327 5 1 1 44326
0 44328 7 1 2 44325 44327
0 44329 5 1 1 44328
0 44330 7 1 2 70077 44329
0 44331 5 1 1 44330
0 44332 7 1 2 69269 93072
0 44333 5 1 1 44332
0 44334 7 1 2 73252 69159
0 44335 5 1 1 44334
0 44336 7 1 2 44335 97052
0 44337 7 1 2 44333 44336
0 44338 5 1 1 44337
0 44339 7 1 2 91128 44338
0 44340 5 1 1 44339
0 44341 7 1 2 44331 44340
0 44342 5 1 1 44341
0 44343 7 1 2 72365 44342
0 44344 5 1 1 44343
0 44345 7 1 2 71460 78006
0 44346 5 1 1 44345
0 44347 7 1 2 69700 77743
0 44348 5 1 1 44347
0 44349 7 2 2 70979 76189
0 44350 7 1 2 72501 97053
0 44351 5 1 1 44350
0 44352 7 1 2 44348 44351
0 44353 5 1 1 44352
0 44354 7 1 2 63138 44353
0 44355 5 1 1 44354
0 44356 7 1 2 44346 44355
0 44357 5 1 1 44356
0 44358 7 1 2 69270 44357
0 44359 5 1 1 44358
0 44360 7 1 2 70457 95782
0 44361 5 1 1 44360
0 44362 7 1 2 87814 44361
0 44363 5 1 1 44362
0 44364 7 1 2 76368 44363
0 44365 5 1 1 44364
0 44366 7 1 2 63139 82217
0 44367 5 1 1 44366
0 44368 7 1 2 44365 44367
0 44369 5 1 1 44368
0 44370 7 1 2 77744 44369
0 44371 5 1 1 44370
0 44372 7 1 2 71124 89528
0 44373 5 1 1 44372
0 44374 7 1 2 90099 44373
0 44375 5 2 1 44374
0 44376 7 1 2 70959 97055
0 44377 5 1 1 44376
0 44378 7 1 2 71125 91100
0 44379 5 1 1 44378
0 44380 7 1 2 44377 44379
0 44381 5 1 1 44380
0 44382 7 1 2 72601 44381
0 44383 5 1 1 44382
0 44384 7 1 2 78615 69145
0 44385 5 1 1 44384
0 44386 7 1 2 78007 44385
0 44387 5 1 1 44386
0 44388 7 1 2 44383 44387
0 44389 7 1 2 44371 44388
0 44390 7 1 2 44359 44389
0 44391 7 1 2 44344 44390
0 44392 7 1 2 44323 44391
0 44393 5 1 1 44392
0 44394 7 1 2 75622 44393
0 44395 5 1 1 44394
0 44396 7 1 2 72457 91263
0 44397 5 1 1 44396
0 44398 7 1 2 62151 44397
0 44399 5 1 1 44398
0 44400 7 1 2 78117 44399
0 44401 5 1 1 44400
0 44402 7 1 2 65896 44401
0 44403 5 1 1 44402
0 44404 7 1 2 70656 91097
0 44405 7 1 2 44403 44404
0 44406 5 1 1 44405
0 44407 7 1 2 62739 44406
0 44408 5 1 1 44407
0 44409 7 1 2 69160 72366
0 44410 5 1 1 44409
0 44411 7 1 2 72481 44410
0 44412 5 1 1 44411
0 44413 7 1 2 88473 44412
0 44414 5 1 1 44413
0 44415 7 2 2 72781 83958
0 44416 5 1 1 97057
0 44417 7 1 2 76649 44416
0 44418 5 1 1 44417
0 44419 7 1 2 44414 44418
0 44420 5 1 1 44419
0 44421 7 1 2 64568 44420
0 44422 5 1 1 44421
0 44423 7 1 2 70209 16154
0 44424 7 1 2 44422 44423
0 44425 7 1 2 44408 44424
0 44426 5 1 1 44425
0 44427 7 1 2 75233 44426
0 44428 5 1 1 44427
0 44429 7 2 2 61123 96254
0 44430 5 1 1 97059
0 44431 7 1 2 67723 81365
0 44432 7 1 2 97060 44431
0 44433 5 1 1 44432
0 44434 7 1 2 75234 44433
0 44435 5 1 1 44434
0 44436 7 2 2 73244 89273
0 44437 5 2 1 97061
0 44438 7 1 2 70078 84281
0 44439 7 1 2 97062 44438
0 44440 5 1 1 44439
0 44441 7 1 2 44435 44440
0 44442 5 1 1 44441
0 44443 7 1 2 63140 44442
0 44444 5 1 1 44443
0 44445 7 1 2 91093 93919
0 44446 5 1 1 44445
0 44447 7 1 2 88449 89520
0 44448 5 1 1 44447
0 44449 7 1 2 75235 44448
0 44450 5 1 1 44449
0 44451 7 1 2 44446 44450
0 44452 5 1 1 44451
0 44453 7 1 2 64569 44452
0 44454 5 1 1 44453
0 44455 7 1 2 63141 73213
0 44456 5 1 1 44455
0 44457 7 2 2 90869 91239
0 44458 5 1 1 97065
0 44459 7 1 2 71327 95930
0 44460 7 1 2 44458 44459
0 44461 5 1 1 44460
0 44462 7 1 2 44456 44461
0 44463 5 1 1 44462
0 44464 7 1 2 75236 44463
0 44465 5 1 1 44464
0 44466 7 1 2 44454 44465
0 44467 5 1 1 44466
0 44468 7 1 2 69271 44467
0 44469 5 1 1 44468
0 44470 7 1 2 44444 44469
0 44471 7 1 2 44428 44470
0 44472 7 1 2 44395 44471
0 44473 5 1 1 44472
0 44474 7 1 2 63539 44473
0 44475 5 1 1 44474
0 44476 7 1 2 66574 97038
0 44477 5 1 1 44476
0 44478 7 1 2 44475 44477
0 44479 7 1 2 44300 44478
0 44480 5 1 1 44479
0 44481 7 1 2 65483 44480
0 44482 5 1 1 44481
0 44483 7 1 2 82822 91182
0 44484 7 2 2 89214 44483
0 44485 5 1 1 97067
0 44486 7 1 2 44482 44485
0 44487 5 2 1 44486
0 44488 7 1 2 66746 97069
0 44489 5 1 1 44488
0 44490 7 1 2 86942 93612
0 44491 7 1 2 88746 44490
0 44492 5 1 1 44491
0 44493 7 1 2 44489 44492
0 44494 5 1 1 44493
0 44495 7 1 2 60701 44494
0 44496 5 1 1 44495
0 44497 7 1 2 80653 84880
0 44498 7 2 2 79266 81777
0 44499 5 1 1 97071
0 44500 7 2 2 77993 70927
0 44501 5 1 1 97073
0 44502 7 1 2 95170 97074
0 44503 7 1 2 97072 44502
0 44504 7 1 2 44497 44503
0 44505 5 1 1 44504
0 44506 7 1 2 44496 44505
0 44507 5 1 1 44506
0 44508 7 1 2 86572 44507
0 44509 5 1 1 44508
0 44510 7 2 2 72161 82895
0 44511 7 2 2 70326 97075
0 44512 5 1 1 97077
0 44513 7 1 2 91170 97078
0 44514 5 1 1 44513
0 44515 7 1 2 91455 95185
0 44516 5 1 1 44515
0 44517 7 1 2 96468 44516
0 44518 5 1 1 44517
0 44519 7 1 2 65740 44518
0 44520 5 1 1 44519
0 44521 7 1 2 76213 82257
0 44522 5 1 1 44521
0 44523 7 1 2 63142 44522
0 44524 5 1 1 44523
0 44525 7 1 2 44520 44524
0 44526 5 1 1 44525
0 44527 7 1 2 64570 44526
0 44528 5 1 1 44527
0 44529 7 1 2 65741 87654
0 44530 5 1 1 44529
0 44531 7 1 2 81475 44530
0 44532 5 1 1 44531
0 44533 7 1 2 64808 44532
0 44534 5 1 1 44533
0 44535 7 1 2 88867 44534
0 44536 5 1 1 44535
0 44537 7 1 2 63143 44536
0 44538 5 1 1 44537
0 44539 7 1 2 44528 44538
0 44540 5 1 1 44539
0 44541 7 1 2 65897 44540
0 44542 5 1 1 44541
0 44543 7 1 2 62740 82307
0 44544 5 1 1 44543
0 44545 7 1 2 78089 44544
0 44546 5 1 1 44545
0 44547 7 1 2 70327 44546
0 44548 5 1 1 44547
0 44549 7 1 2 62741 83285
0 44550 5 1 1 44549
0 44551 7 1 2 44548 44550
0 44552 5 1 1 44551
0 44553 7 1 2 63144 44552
0 44554 5 1 1 44553
0 44555 7 1 2 44542 44554
0 44556 5 1 1 44555
0 44557 7 1 2 66068 44556
0 44558 5 1 1 44557
0 44559 7 1 2 44514 44558
0 44560 5 1 1 44559
0 44561 7 1 2 68483 44560
0 44562 5 1 1 44561
0 44563 7 1 2 85381 44562
0 44564 5 1 1 44563
0 44565 7 1 2 91863 44564
0 44566 5 1 1 44565
0 44567 7 1 2 82201 78110
0 44568 5 1 1 44567
0 44569 7 1 2 71239 44568
0 44570 5 1 1 44569
0 44571 7 1 2 84881 93202
0 44572 7 1 2 44570 44571
0 44573 5 1 1 44572
0 44574 7 1 2 44566 44573
0 44575 5 1 1 44574
0 44576 7 1 2 63814 44575
0 44577 5 1 1 44576
0 44578 7 3 2 65279 87825
0 44579 7 1 2 89690 97079
0 44580 5 1 1 44579
0 44581 7 1 2 44577 44580
0 44582 5 1 1 44581
0 44583 7 1 2 61771 44582
0 44584 5 1 1 44583
0 44585 7 1 2 74034 89364
0 44586 5 1 1 44585
0 44587 7 1 2 70328 76961
0 44588 5 1 1 44587
0 44589 7 1 2 44586 44588
0 44590 5 1 1 44589
0 44591 7 1 2 67724 44590
0 44592 5 1 1 44591
0 44593 7 1 2 67370 93066
0 44594 5 1 1 44593
0 44595 7 1 2 44592 44594
0 44596 5 1 1 44595
0 44597 7 1 2 84507 44596
0 44598 5 1 1 44597
0 44599 7 1 2 73690 82152
0 44600 5 1 1 44599
0 44601 7 1 2 84571 44600
0 44602 5 1 1 44601
0 44603 7 1 2 64571 44602
0 44604 5 1 1 44603
0 44605 7 1 2 79363 76190
0 44606 5 2 1 44605
0 44607 7 1 2 44604 97082
0 44608 5 1 1 44607
0 44609 7 1 2 69701 44608
0 44610 5 1 1 44609
0 44611 7 1 2 82910 85778
0 44612 5 1 1 44611
0 44613 7 1 2 66747 71377
0 44614 5 1 1 44613
0 44615 7 1 2 67725 82685
0 44616 5 1 1 44615
0 44617 7 1 2 94661 44616
0 44618 7 1 2 44614 44617
0 44619 5 1 1 44618
0 44620 7 1 2 44612 44619
0 44621 7 1 2 44610 44620
0 44622 5 1 1 44621
0 44623 7 1 2 84188 44622
0 44624 5 1 1 44623
0 44625 7 1 2 44598 44624
0 44626 5 1 1 44625
0 44627 7 1 2 65898 44626
0 44628 5 1 1 44627
0 44629 7 3 2 68757 93640
0 44630 5 1 1 97084
0 44631 7 1 2 76962 97085
0 44632 5 1 1 44631
0 44633 7 1 2 63815 80127
0 44634 5 1 1 44633
0 44635 7 1 2 44632 44634
0 44636 5 1 1 44635
0 44637 7 1 2 62742 44636
0 44638 5 1 1 44637
0 44639 7 1 2 83286 78160
0 44640 5 1 1 44639
0 44641 7 1 2 44638 44640
0 44642 5 1 1 44641
0 44643 7 1 2 70329 44642
0 44644 5 1 1 44643
0 44645 7 1 2 74787 84189
0 44646 5 2 1 44645
0 44647 7 1 2 78166 97087
0 44648 5 1 1 44647
0 44649 7 1 2 82911 44648
0 44650 5 1 1 44649
0 44651 7 1 2 44644 44650
0 44652 5 1 1 44651
0 44653 7 1 2 61772 44652
0 44654 5 1 1 44653
0 44655 7 1 2 44628 44654
0 44656 5 1 1 44655
0 44657 7 1 2 66069 44656
0 44658 5 1 1 44657
0 44659 7 1 2 63816 88804
0 44660 5 1 1 44659
0 44661 7 1 2 62378 44630
0 44662 5 1 1 44661
0 44663 7 1 2 71829 19831
0 44664 7 1 2 44662 44663
0 44665 5 1 1 44664
0 44666 7 3 2 68758 94392
0 44667 5 1 1 97089
0 44668 7 1 2 64328 97090
0 44669 5 1 1 44668
0 44670 7 1 2 62743 44669
0 44671 7 1 2 44665 44670
0 44672 5 1 1 44671
0 44673 7 1 2 70330 7690
0 44674 7 1 2 89382 44673
0 44675 7 1 2 44672 44674
0 44676 5 1 1 44675
0 44677 7 1 2 44660 44676
0 44678 5 1 1 44677
0 44679 7 1 2 79426 44678
0 44680 5 1 1 44679
0 44681 7 1 2 44658 44680
0 44682 5 1 1 44681
0 44683 7 1 2 63145 44682
0 44684 5 1 1 44683
0 44685 7 2 2 63817 88511
0 44686 7 1 2 79364 85574
0 44687 7 1 2 97092 44686
0 44688 5 1 1 44687
0 44689 7 1 2 44684 44688
0 44690 5 1 1 44689
0 44691 7 1 2 63540 44690
0 44692 5 1 1 44691
0 44693 7 2 2 70331 91442
0 44694 5 1 1 97094
0 44695 7 1 2 72428 44694
0 44696 5 1 1 44695
0 44697 7 1 2 82185 84508
0 44698 7 1 2 44696 44697
0 44699 5 1 1 44698
0 44700 7 1 2 44692 44699
0 44701 5 1 1 44700
0 44702 7 1 2 75623 44701
0 44703 5 1 1 44702
0 44704 7 1 2 74429 89898
0 44705 5 2 1 44704
0 44706 7 1 2 2689 97096
0 44707 5 1 1 44706
0 44708 7 1 2 64809 44707
0 44709 5 1 1 44708
0 44710 7 1 2 84114 91375
0 44711 5 1 1 44710
0 44712 7 1 2 44709 44711
0 44713 5 1 1 44712
0 44714 7 1 2 77798 44713
0 44715 5 1 1 44714
0 44716 7 5 2 62152 77917
0 44717 5 1 1 97098
0 44718 7 1 2 75911 97099
0 44719 5 1 1 44718
0 44720 7 1 2 44715 44719
0 44721 5 1 1 44720
0 44722 7 1 2 66070 44721
0 44723 5 1 1 44722
0 44724 7 1 2 69072 85946
0 44725 5 1 1 44724
0 44726 7 1 2 77944 44725
0 44727 5 1 1 44726
0 44728 7 1 2 64572 44727
0 44729 5 2 1 44728
0 44730 7 1 2 68104 86851
0 44731 5 1 1 44730
0 44732 7 1 2 97103 44731
0 44733 5 1 1 44732
0 44734 7 1 2 70332 44733
0 44735 5 1 1 44734
0 44736 7 1 2 72439 77918
0 44737 5 1 1 44736
0 44738 7 1 2 44735 44737
0 44739 5 1 1 44738
0 44740 7 1 2 64329 44739
0 44741 5 1 1 44740
0 44742 7 1 2 62379 79988
0 44743 5 1 1 44742
0 44744 7 1 2 67726 44743
0 44745 5 1 1 44744
0 44746 7 1 2 77919 44745
0 44747 5 1 1 44746
0 44748 7 1 2 44741 44747
0 44749 7 1 2 44723 44748
0 44750 5 1 1 44749
0 44751 7 1 2 94681 97080
0 44752 7 1 2 44750 44751
0 44753 5 1 1 44752
0 44754 7 1 2 44703 44753
0 44755 7 1 2 44584 44754
0 44756 5 1 1 44755
0 44757 7 1 2 70840 44756
0 44758 5 1 1 44757
0 44759 7 1 2 70409 77920
0 44760 5 1 1 44759
0 44761 7 1 2 80739 95350
0 44762 5 1 1 44761
0 44763 7 1 2 44760 44762
0 44764 5 1 1 44763
0 44765 7 1 2 62744 44764
0 44766 5 1 1 44765
0 44767 7 1 2 1967 78604
0 44768 5 1 1 44767
0 44769 7 1 2 65028 44768
0 44770 5 1 1 44769
0 44771 7 1 2 65280 95580
0 44772 5 1 1 44771
0 44773 7 1 2 44770 44772
0 44774 5 1 1 44773
0 44775 7 1 2 68484 44774
0 44776 5 1 1 44775
0 44777 7 1 2 44766 44776
0 44778 5 1 1 44777
0 44779 7 1 2 64330 44778
0 44780 5 1 1 44779
0 44781 7 1 2 65281 73048
0 44782 5 1 1 44781
0 44783 7 1 2 63146 87006
0 44784 5 1 1 44783
0 44785 7 1 2 44782 44784
0 44786 5 1 1 44785
0 44787 7 1 2 95028 44786
0 44788 5 1 1 44787
0 44789 7 1 2 77436 84742
0 44790 5 3 1 44789
0 44791 7 1 2 95409 97105
0 44792 5 1 1 44791
0 44793 7 1 2 70333 44792
0 44794 5 1 1 44793
0 44795 7 1 2 44788 44794
0 44796 7 1 2 44780 44795
0 44797 5 1 1 44796
0 44798 7 1 2 72022 44797
0 44799 5 1 1 44798
0 44800 7 1 2 95456 95403
0 44801 5 1 1 44800
0 44802 7 1 2 63541 44801
0 44803 5 1 1 44802
0 44804 7 1 2 76752 90307
0 44805 5 1 1 44804
0 44806 7 1 2 81423 94334
0 44807 5 1 1 44806
0 44808 7 1 2 44805 44807
0 44809 5 1 1 44808
0 44810 7 1 2 71830 44809
0 44811 5 1 1 44810
0 44812 7 1 2 95395 44811
0 44813 5 1 1 44812
0 44814 7 1 2 68485 44813
0 44815 5 1 1 44814
0 44816 7 1 2 75690 83914
0 44817 5 2 1 44816
0 44818 7 1 2 44815 97108
0 44819 7 1 2 44803 44818
0 44820 7 1 2 44799 44819
0 44821 5 1 1 44820
0 44822 7 1 2 72367 44821
0 44823 5 1 1 44822
0 44824 7 1 2 60943 76540
0 44825 5 1 1 44824
0 44826 7 1 2 65282 89797
0 44827 7 1 2 44825 44826
0 44828 5 1 1 44827
0 44829 7 1 2 63542 44828
0 44830 5 1 1 44829
0 44831 7 1 2 95384 44830
0 44832 5 1 1 44831
0 44833 7 1 2 66575 44832
0 44834 5 1 1 44833
0 44835 7 1 2 71579 81467
0 44836 5 1 1 44835
0 44837 7 2 2 70334 89899
0 44838 7 1 2 76902 97110
0 44839 5 2 1 44838
0 44840 7 1 2 90023 97112
0 44841 5 3 1 44840
0 44842 7 1 2 70841 97114
0 44843 5 1 1 44842
0 44844 7 1 2 44836 44843
0 44845 5 1 1 44844
0 44846 7 1 2 68486 44845
0 44847 5 1 1 44846
0 44848 7 1 2 95386 44847
0 44849 5 1 1 44848
0 44850 7 1 2 63147 44849
0 44851 5 1 1 44850
0 44852 7 1 2 72849 90330
0 44853 5 1 1 44852
0 44854 7 1 2 76807 44853
0 44855 5 1 1 44854
0 44856 7 1 2 68487 44855
0 44857 5 1 1 44856
0 44858 7 1 2 77921 77276
0 44859 5 1 1 44858
0 44860 7 1 2 64573 88543
0 44861 5 1 1 44860
0 44862 7 1 2 77945 44861
0 44863 5 2 1 44862
0 44864 7 1 2 88442 97117
0 44865 5 1 1 44864
0 44866 7 1 2 44859 44865
0 44867 7 1 2 44857 44866
0 44868 5 1 1 44867
0 44869 7 1 2 62380 44868
0 44870 5 1 1 44869
0 44871 7 1 2 72850 97118
0 44872 5 1 1 44871
0 44873 7 1 2 74788 88306
0 44874 5 1 1 44873
0 44875 7 1 2 68488 76808
0 44876 7 1 2 44874 44875
0 44877 5 1 1 44876
0 44878 7 3 2 63543 76268
0 44879 5 1 1 97119
0 44880 7 1 2 83119 44879
0 44881 7 1 2 44877 44880
0 44882 5 1 1 44881
0 44883 7 1 2 44872 44882
0 44884 5 1 1 44883
0 44885 7 1 2 62745 44884
0 44886 5 1 1 44885
0 44887 7 1 2 73116 90331
0 44888 5 1 1 44887
0 44889 7 1 2 76809 44888
0 44890 5 1 1 44889
0 44891 7 1 2 68489 44890
0 44892 5 1 1 44891
0 44893 7 1 2 77922 88046
0 44894 5 1 1 44893
0 44895 7 1 2 44892 44894
0 44896 5 1 1 44895
0 44897 7 1 2 76369 44896
0 44898 5 1 1 44897
0 44899 7 1 2 76753 92885
0 44900 5 1 1 44899
0 44901 7 1 2 87966 44900
0 44902 7 1 2 44898 44901
0 44903 7 1 2 44886 44902
0 44904 7 1 2 44870 44903
0 44905 7 1 2 44851 44904
0 44906 5 1 1 44905
0 44907 7 1 2 71126 44906
0 44908 5 1 1 44907
0 44909 7 1 2 81429 75077
0 44910 5 1 1 44909
0 44911 7 1 2 31821 44910
0 44912 5 1 1 44911
0 44913 7 1 2 62746 44912
0 44914 5 1 1 44913
0 44915 7 2 2 63544 87357
0 44916 5 1 1 97122
0 44917 7 1 2 70549 97123
0 44918 5 1 1 44917
0 44919 7 1 2 44914 44918
0 44920 5 1 1 44919
0 44921 7 1 2 70842 44920
0 44922 5 1 1 44921
0 44923 7 1 2 79798 95420
0 44924 5 1 1 44923
0 44925 7 1 2 78349 90332
0 44926 5 1 1 44925
0 44927 7 1 2 76810 44926
0 44928 5 1 1 44927
0 44929 7 1 2 68490 44928
0 44930 5 1 1 44929
0 44931 7 1 2 44924 44930
0 44932 5 1 1 44931
0 44933 7 1 2 63148 44932
0 44934 5 1 1 44933
0 44935 7 1 2 85005 44934
0 44936 7 1 2 44922 44935
0 44937 5 1 1 44936
0 44938 7 1 2 71831 44937
0 44939 5 1 1 44938
0 44940 7 1 2 73182 87616
0 44941 5 1 1 44940
0 44942 7 1 2 65283 44941
0 44943 5 1 1 44942
0 44944 7 1 2 4541 11688
0 44945 5 1 1 44944
0 44946 7 1 2 65029 44945
0 44947 5 1 1 44946
0 44948 7 1 2 44943 44947
0 44949 5 1 1 44948
0 44950 7 1 2 68491 44949
0 44951 5 1 1 44950
0 44952 7 1 2 73691 85374
0 44953 5 1 1 44952
0 44954 7 1 2 44951 44953
0 44955 5 1 1 44954
0 44956 7 1 2 69702 44955
0 44957 5 1 1 44956
0 44958 7 1 2 11473 44717
0 44959 5 1 1 44958
0 44960 7 1 2 70843 44959
0 44961 5 1 1 44960
0 44962 7 1 2 13040 44961
0 44963 5 1 1 44962
0 44964 7 1 2 62381 44963
0 44965 5 1 1 44964
0 44966 7 1 2 77946 87753
0 44967 5 1 1 44966
0 44968 7 1 2 70844 44967
0 44969 5 1 1 44968
0 44970 7 1 2 95410 44969
0 44971 5 1 1 44970
0 44972 7 1 2 88040 44971
0 44973 5 1 1 44972
0 44974 7 1 2 95407 44973
0 44975 7 1 2 44965 44974
0 44976 7 1 2 44957 44975
0 44977 5 1 1 44976
0 44978 7 1 2 78669 44977
0 44979 5 1 1 44978
0 44980 7 1 2 60399 87008
0 44981 5 1 1 44980
0 44982 7 1 2 70079 44981
0 44983 5 1 1 44982
0 44984 7 1 2 87882 90425
0 44985 5 1 1 44984
0 44986 7 1 2 44983 44985
0 44987 5 1 1 44986
0 44988 7 1 2 68492 44987
0 44989 5 1 1 44988
0 44990 7 1 2 83367 75078
0 44991 5 1 1 44990
0 44992 7 1 2 79820 44991
0 44993 5 1 1 44992
0 44994 7 1 2 70845 44993
0 44995 5 1 1 44994
0 44996 7 1 2 59966 84724
0 44997 5 1 1 44996
0 44998 7 1 2 61605 69373
0 44999 5 1 1 44998
0 45000 7 1 2 44997 44999
0 45001 5 1 1 45000
0 45002 7 1 2 75691 45001
0 45003 5 1 1 45002
0 45004 7 1 2 44995 45003
0 45005 7 1 2 44989 45004
0 45006 5 1 1 45005
0 45007 7 1 2 63149 45006
0 45008 5 1 1 45007
0 45009 7 1 2 81657 85001
0 45010 5 1 1 45009
0 45011 7 1 2 75153 87381
0 45012 5 1 1 45011
0 45013 7 1 2 63545 45012
0 45014 5 1 1 45013
0 45015 7 1 2 45010 45014
0 45016 7 1 2 45008 45015
0 45017 7 1 2 77947 90688
0 45018 5 1 1 45017
0 45019 7 1 2 62153 87031
0 45020 7 1 2 45018 45019
0 45021 5 1 1 45020
0 45022 7 1 2 85006 45021
0 45023 5 1 1 45022
0 45024 7 1 2 65742 45023
0 45025 5 1 1 45024
0 45026 7 1 2 76650 87965
0 45027 5 1 1 45026
0 45028 7 1 2 45025 45027
0 45029 5 1 1 45028
0 45030 7 1 2 64331 45029
0 45031 5 1 1 45030
0 45032 7 1 2 89220 97106
0 45033 5 1 1 45032
0 45034 7 1 2 70846 45033
0 45035 5 1 1 45034
0 45036 7 1 2 62382 88544
0 45037 5 1 1 45036
0 45038 7 1 2 79821 45037
0 45039 5 1 1 45038
0 45040 7 1 2 86629 45039
0 45041 5 1 1 45040
0 45042 7 1 2 45035 45041
0 45043 5 1 1 45042
0 45044 7 1 2 70335 45043
0 45045 5 1 1 45044
0 45046 7 1 2 45031 45045
0 45047 7 1 2 45016 45046
0 45048 7 1 2 44979 45047
0 45049 7 1 2 44939 45048
0 45050 7 1 2 44908 45049
0 45051 7 1 2 44834 45050
0 45052 7 1 2 44823 45051
0 45053 5 1 1 45052
0 45054 7 1 2 65484 45053
0 45055 5 1 1 45054
0 45056 7 1 2 68759 95454
0 45057 7 1 2 45055 45056
0 45058 5 1 1 45057
0 45059 7 1 2 76348 91498
0 45060 5 2 1 45059
0 45061 7 1 2 89878 97124
0 45062 5 1 1 45061
0 45063 7 1 2 65899 78646
0 45064 5 1 1 45063
0 45065 7 1 2 88552 45064
0 45066 5 1 1 45065
0 45067 7 1 2 62154 45066
0 45068 5 1 1 45067
0 45069 7 1 2 71832 91261
0 45070 5 1 1 45069
0 45071 7 1 2 71240 45070
0 45072 7 1 2 45068 45071
0 45073 5 1 1 45072
0 45074 7 1 2 62383 45073
0 45075 5 1 1 45074
0 45076 7 1 2 76370 90528
0 45077 5 1 1 45076
0 45078 7 1 2 37765 45077
0 45079 7 1 2 45075 45078
0 45080 5 1 1 45079
0 45081 7 1 2 84835 45080
0 45082 5 1 1 45081
0 45083 7 1 2 45062 45082
0 45084 5 1 1 45083
0 45085 7 1 2 62747 45084
0 45086 5 1 1 45085
0 45087 7 1 2 61606 78682
0 45088 7 1 2 90926 45087
0 45089 5 1 1 45088
0 45090 7 1 2 45086 45089
0 45091 5 1 1 45090
0 45092 7 1 2 71580 45091
0 45093 5 1 1 45092
0 45094 7 1 2 17565 91301
0 45095 7 2 2 85606 90861
0 45096 7 1 2 70928 97126
0 45097 5 1 1 45096
0 45098 7 1 2 69272 79112
0 45099 5 1 1 45098
0 45100 7 1 2 34694 45099
0 45101 5 1 1 45100
0 45102 7 1 2 64574 45101
0 45103 5 1 1 45102
0 45104 7 1 2 63150 90502
0 45105 5 1 1 45104
0 45106 7 1 2 64810 95568
0 45107 5 1 1 45106
0 45108 7 1 2 89045 45107
0 45109 5 1 1 45108
0 45110 7 1 2 69073 45109
0 45111 5 1 1 45110
0 45112 7 1 2 45105 45111
0 45113 7 1 2 45103 45112
0 45114 5 1 1 45113
0 45115 7 1 2 66576 45114
0 45116 5 1 1 45115
0 45117 7 1 2 45097 45116
0 45118 5 1 1 45117
0 45119 7 1 2 69703 45118
0 45120 5 1 1 45119
0 45121 7 1 2 62155 93479
0 45122 5 1 1 45121
0 45123 7 1 2 77505 45122
0 45124 5 1 1 45123
0 45125 7 1 2 65900 45124
0 45126 5 1 1 45125
0 45127 7 1 2 68105 88868
0 45128 5 2 1 45127
0 45129 7 1 2 72368 97128
0 45130 5 1 1 45129
0 45131 7 1 2 88819 90971
0 45132 7 1 2 45130 45131
0 45133 7 1 2 45126 45132
0 45134 5 1 1 45133
0 45135 7 1 2 69273 45134
0 45136 5 1 1 45135
0 45137 7 1 2 70996 90980
0 45138 5 1 1 45137
0 45139 7 1 2 66071 45138
0 45140 5 1 1 45139
0 45141 7 1 2 74125 90984
0 45142 7 1 2 88699 45141
0 45143 5 1 1 45142
0 45144 7 1 2 45140 45143
0 45145 5 1 1 45144
0 45146 7 1 2 64811 45145
0 45147 5 1 1 45146
0 45148 7 1 2 63151 91589
0 45149 5 1 1 45148
0 45150 7 1 2 45147 45149
0 45151 7 1 2 45136 45150
0 45152 5 1 1 45151
0 45153 7 1 2 66577 45152
0 45154 5 1 1 45153
0 45155 7 1 2 45120 45154
0 45156 7 1 2 45094 45155
0 45157 5 1 1 45156
0 45158 7 1 2 60592 45157
0 45159 5 1 1 45158
0 45160 7 1 2 82308 78670
0 45161 5 1 1 45160
0 45162 7 1 2 88368 45161
0 45163 5 2 1 45162
0 45164 7 1 2 70336 97130
0 45165 5 1 1 45164
0 45166 7 1 2 77252 73135
0 45167 5 1 1 45166
0 45168 7 1 2 88654 45167
0 45169 5 1 1 45168
0 45170 7 1 2 2559 45169
0 45171 7 1 2 64812 71630
0 45172 7 1 2 73985 45171
0 45173 5 1 1 45172
0 45174 7 1 2 67371 70466
0 45175 5 3 1 45174
0 45176 7 2 2 70372 97132
0 45177 5 1 1 97135
0 45178 7 1 2 72369 97136
0 45179 5 1 1 45178
0 45180 7 1 2 45173 45179
0 45181 7 1 2 45170 45180
0 45182 7 1 2 45165 45181
0 45183 5 1 1 45182
0 45184 7 1 2 62748 45183
0 45185 5 1 1 45184
0 45186 7 1 2 75520 45185
0 45187 5 1 1 45186
0 45188 7 1 2 89879 45187
0 45189 5 1 1 45188
0 45190 7 2 2 65284 84836
0 45191 5 1 1 97137
0 45192 7 1 2 85463 45191
0 45193 5 1 1 45192
0 45194 7 1 2 95788 45193
0 45195 5 1 1 45194
0 45196 7 1 2 77437 84951
0 45197 7 1 2 80315 45196
0 45198 5 1 1 45197
0 45199 7 1 2 45195 45198
0 45200 7 1 2 45189 45199
0 45201 5 1 1 45200
0 45202 7 1 2 70847 45201
0 45203 5 1 1 45202
0 45204 7 1 2 74919 87437
0 45205 5 1 1 45204
0 45206 7 1 2 85411 45205
0 45207 5 1 1 45206
0 45208 7 1 2 59630 45207
0 45209 5 1 1 45208
0 45210 7 1 2 67372 95830
0 45211 5 1 1 45210
0 45212 7 2 2 45209 45211
0 45213 5 1 1 97139
0 45214 7 1 2 84391 97140
0 45215 5 1 1 45214
0 45216 7 1 2 76811 45215
0 45217 5 1 1 45216
0 45218 7 1 2 79470 84837
0 45219 5 1 1 45218
0 45220 7 1 2 84601 88999
0 45221 5 1 1 45220
0 45222 7 1 2 75624 88112
0 45223 7 1 2 45221 45222
0 45224 5 1 1 45223
0 45225 7 1 2 65485 94566
0 45226 7 1 2 45224 45225
0 45227 5 1 1 45226
0 45228 7 1 2 45219 45227
0 45229 7 1 2 45217 45228
0 45230 7 1 2 45203 45229
0 45231 7 1 2 45159 45230
0 45232 7 1 2 45093 45231
0 45233 5 1 1 45232
0 45234 7 1 2 68493 45233
0 45235 5 1 1 45234
0 45236 7 1 2 60593 95867
0 45237 5 1 1 45236
0 45238 7 1 2 4875 45237
0 45239 5 1 1 45238
0 45240 7 1 2 63546 45239
0 45241 5 1 1 45240
0 45242 7 1 2 80042 73330
0 45243 7 1 2 94025 45242
0 45244 5 1 1 45243
0 45245 7 1 2 95630 96767
0 45246 5 1 1 45245
0 45247 7 1 2 93456 45246
0 45248 7 1 2 45244 45247
0 45249 7 1 2 45241 45248
0 45250 5 1 1 45249
0 45251 7 1 2 68106 45250
0 45252 5 1 1 45251
0 45253 7 1 2 63152 82088
0 45254 5 1 1 45253
0 45255 7 1 2 74554 45254
0 45256 5 2 1 45255
0 45257 7 1 2 70657 97141
0 45258 5 1 1 45257
0 45259 7 1 2 83304 74263
0 45260 5 1 1 45259
0 45261 7 1 2 45258 45260
0 45262 5 1 1 45261
0 45263 7 1 2 63547 45262
0 45264 5 1 1 45263
0 45265 7 1 2 79936 85408
0 45266 5 1 1 45265
0 45267 7 1 2 45264 45266
0 45268 5 1 1 45267
0 45269 7 1 2 69586 45268
0 45270 5 1 1 45269
0 45271 7 1 2 85626 45270
0 45272 5 1 1 45271
0 45273 7 1 2 59631 45272
0 45274 5 1 1 45273
0 45275 7 1 2 90587 96062
0 45276 5 1 1 45275
0 45277 7 1 2 68107 45276
0 45278 5 1 1 45277
0 45279 7 1 2 45274 45278
0 45280 5 1 1 45279
0 45281 7 1 2 72243 45280
0 45282 5 1 1 45281
0 45283 7 1 2 88581 88747
0 45284 5 1 1 45283
0 45285 7 1 2 71581 73049
0 45286 5 1 1 45285
0 45287 7 1 2 30048 45286
0 45288 5 1 1 45287
0 45289 7 1 2 72370 45288
0 45290 5 1 1 45289
0 45291 7 1 2 78851 45290
0 45292 7 1 2 45284 45291
0 45293 5 1 1 45292
0 45294 7 1 2 85917 45293
0 45295 5 1 1 45294
0 45296 7 1 2 75456 94581
0 45297 5 1 1 45296
0 45298 7 1 2 90612 45297
0 45299 5 1 1 45298
0 45300 7 1 2 85918 91047
0 45301 5 1 1 45300
0 45302 7 1 2 62384 90613
0 45303 5 1 1 45302
0 45304 7 1 2 45301 45303
0 45305 5 1 1 45304
0 45306 7 1 2 88760 45305
0 45307 5 1 1 45306
0 45308 7 1 2 88582 89891
0 45309 7 1 2 94585 45308
0 45310 5 1 1 45309
0 45311 7 1 2 45307 45310
0 45312 7 1 2 45299 45311
0 45313 7 1 2 45295 45312
0 45314 5 1 1 45313
0 45315 7 1 2 63153 45314
0 45316 5 1 1 45315
0 45317 7 1 2 83512 90702
0 45318 5 1 1 45317
0 45319 7 1 2 65486 45318
0 45320 5 1 1 45319
0 45321 7 1 2 93558 45320
0 45322 7 1 2 45316 45321
0 45323 7 1 2 45282 45322
0 45324 5 1 1 45323
0 45325 7 1 2 67727 45324
0 45326 5 1 1 45325
0 45327 7 1 2 63818 45326
0 45328 7 1 2 45252 45327
0 45329 7 1 2 45235 45328
0 45330 5 1 1 45329
0 45331 7 1 2 66748 45330
0 45332 7 1 2 45058 45331
0 45333 5 1 1 45332
0 45334 7 1 2 64813 96390
0 45335 5 1 1 45334
0 45336 7 1 2 88869 45335
0 45337 5 1 1 45336
0 45338 7 1 2 75625 45337
0 45339 5 1 1 45338
0 45340 7 1 2 79192 90345
0 45341 5 1 1 45340
0 45342 7 1 2 45339 45341
0 45343 5 1 1 45342
0 45344 7 1 2 65901 45343
0 45345 5 1 1 45344
0 45346 7 1 2 73881 90385
0 45347 5 1 1 45346
0 45348 7 1 2 45345 45347
0 45349 5 1 1 45348
0 45350 7 1 2 84190 45349
0 45351 5 1 1 45350
0 45352 7 1 2 67728 72793
0 45353 5 4 1 45352
0 45354 7 1 2 65285 97143
0 45355 5 1 1 45354
0 45356 7 1 2 65902 94856
0 45357 5 1 1 45356
0 45358 7 1 2 45355 45357
0 45359 5 1 1 45358
0 45360 7 1 2 64575 45359
0 45361 5 1 1 45360
0 45362 7 1 2 65286 82140
0 45363 5 1 1 45362
0 45364 7 1 2 45361 45363
0 45365 5 1 1 45364
0 45366 7 1 2 84509 45365
0 45367 5 1 1 45366
0 45368 7 1 2 45351 45367
0 45369 5 1 1 45368
0 45370 7 1 2 66072 45369
0 45371 5 1 1 45370
0 45372 7 2 2 85192 86425
0 45373 7 1 2 95653 97147
0 45374 5 1 1 45373
0 45375 7 1 2 78647 97148
0 45376 5 1 1 45375
0 45377 7 2 2 71127 84191
0 45378 5 1 1 97149
0 45379 7 1 2 91232 97150
0 45380 5 1 1 45379
0 45381 7 1 2 45376 45380
0 45382 5 1 1 45381
0 45383 7 1 2 76371 45382
0 45384 5 1 1 45383
0 45385 7 1 2 45374 45384
0 45386 7 1 2 45371 45385
0 45387 5 1 1 45386
0 45388 7 1 2 62385 45387
0 45389 5 1 1 45388
0 45390 7 4 2 65743 93583
0 45391 5 1 1 97151
0 45392 7 1 2 82288 97152
0 45393 5 1 1 45392
0 45394 7 2 2 84192 76871
0 45395 5 1 1 97155
0 45396 7 1 2 89365 97156
0 45397 5 1 1 45396
0 45398 7 1 2 45393 45397
0 45399 5 1 1 45398
0 45400 7 1 2 66073 93395
0 45401 7 1 2 45399 45400
0 45402 5 1 1 45401
0 45403 7 1 2 68108 84705
0 45404 7 1 2 45402 45403
0 45405 7 1 2 45389 45404
0 45406 5 1 1 45405
0 45407 7 1 2 84590 93548
0 45408 5 2 1 45407
0 45409 7 1 2 78167 97157
0 45410 5 1 1 45409
0 45411 7 1 2 64332 45410
0 45412 5 1 1 45411
0 45413 7 2 2 67729 69274
0 45414 5 1 1 97159
0 45415 7 1 2 63819 97160
0 45416 5 1 1 45415
0 45417 7 2 2 67730 88688
0 45418 5 1 1 97161
0 45419 7 1 2 84193 45418
0 45420 5 1 1 45419
0 45421 7 1 2 45416 45420
0 45422 7 1 2 45412 45421
0 45423 5 1 1 45422
0 45424 7 1 2 65287 45423
0 45425 5 1 1 45424
0 45426 7 1 2 64333 92063
0 45427 7 1 2 91276 45426
0 45428 5 1 1 45427
0 45429 7 1 2 45425 45428
0 45430 5 1 1 45429
0 45431 7 1 2 61773 45430
0 45432 5 1 1 45431
0 45433 7 1 2 69704 88404
0 45434 5 1 1 45433
0 45435 7 1 2 90358 45434
0 45436 5 1 1 45435
0 45437 7 1 2 67101 45436
0 45438 5 1 1 45437
0 45439 7 1 2 74282 75934
0 45440 5 1 1 45439
0 45441 7 1 2 45438 45440
0 45442 5 1 1 45441
0 45443 7 1 2 83448 90901
0 45444 7 1 2 45442 45443
0 45445 5 1 1 45444
0 45446 7 1 2 45432 45445
0 45447 5 1 1 45446
0 45448 7 1 2 64576 45447
0 45449 5 1 1 45448
0 45450 7 1 2 81482 72371
0 45451 5 1 1 45450
0 45452 7 1 2 62386 88440
0 45453 5 1 1 45452
0 45454 7 1 2 45451 45453
0 45455 5 1 1 45454
0 45456 7 1 2 61774 45455
0 45457 5 1 1 45456
0 45458 7 1 2 67102 19280
0 45459 5 1 1 45458
0 45460 7 1 2 74283 72563
0 45461 5 1 1 45460
0 45462 7 1 2 95438 45461
0 45463 7 1 2 45459 45462
0 45464 5 1 1 45463
0 45465 7 1 2 90460 45464
0 45466 5 1 1 45465
0 45467 7 1 2 45457 45466
0 45468 5 1 1 45467
0 45469 7 1 2 84194 45468
0 45470 5 1 1 45469
0 45471 7 2 2 63820 86454
0 45472 7 1 2 72244 94269
0 45473 5 1 1 45472
0 45474 7 1 2 97163 45473
0 45475 5 1 1 45474
0 45476 7 1 2 45470 45475
0 45477 5 1 1 45476
0 45478 7 1 2 65288 45477
0 45479 5 1 1 45478
0 45480 7 1 2 63154 45479
0 45481 7 1 2 45449 45480
0 45482 5 1 1 45481
0 45483 7 1 2 45406 45482
0 45484 5 1 1 45483
0 45485 7 1 2 84510 86923
0 45486 5 1 1 45485
0 45487 7 1 2 21122 45486
0 45488 5 1 1 45487
0 45489 7 1 2 78534 93401
0 45490 5 1 1 45489
0 45491 7 1 2 60400 45490
0 45492 5 1 1 45491
0 45493 7 1 2 45488 45492
0 45494 5 1 1 45493
0 45495 7 1 2 63548 45494
0 45496 7 1 2 45484 45495
0 45497 5 1 1 45496
0 45498 7 1 2 90447 97050
0 45499 5 1 1 45498
0 45500 7 1 2 60594 45499
0 45501 5 1 1 45500
0 45502 7 1 2 84511 45501
0 45503 5 1 1 45502
0 45504 7 1 2 68109 91007
0 45505 5 1 1 45504
0 45506 7 1 2 84195 45505
0 45507 5 1 1 45506
0 45508 7 1 2 80437 74754
0 45509 5 1 1 45508
0 45510 7 1 2 71314 45509
0 45511 5 1 1 45510
0 45512 7 1 2 68110 45511
0 45513 5 1 1 45512
0 45514 7 1 2 84512 45513
0 45515 5 1 1 45514
0 45516 7 1 2 45507 45515
0 45517 5 1 1 45516
0 45518 7 1 2 64814 45517
0 45519 5 1 1 45518
0 45520 7 1 2 74806 88292
0 45521 5 2 1 45520
0 45522 7 1 2 64577 97165
0 45523 5 1 1 45522
0 45524 7 1 2 76732 45523
0 45525 5 1 1 45524
0 45526 7 1 2 84258 45525
0 45527 5 1 1 45526
0 45528 7 1 2 45519 45527
0 45529 5 1 1 45528
0 45530 7 1 2 62749 45529
0 45531 5 1 1 45530
0 45532 7 1 2 81317 95213
0 45533 5 1 1 45532
0 45534 7 1 2 88242 45533
0 45535 5 1 1 45534
0 45536 7 1 2 64334 45535
0 45537 5 1 1 45536
0 45538 7 1 2 73990 84513
0 45539 5 1 1 45538
0 45540 7 1 2 45537 45539
0 45541 5 1 1 45540
0 45542 7 1 2 91456 45541
0 45543 5 1 1 45542
0 45544 7 1 2 84591 87447
0 45545 7 1 2 90448 45544
0 45546 5 1 1 45545
0 45547 7 1 2 9357 45546
0 45548 5 1 1 45547
0 45549 7 1 2 64335 45548
0 45550 5 1 1 45549
0 45551 7 1 2 71635 84514
0 45552 5 1 1 45551
0 45553 7 1 2 59632 45552
0 45554 5 1 1 45553
0 45555 7 3 2 68760 85827
0 45556 5 1 1 97167
0 45557 7 1 2 84553 45556
0 45558 5 3 1 45557
0 45559 7 1 2 63155 97170
0 45560 7 1 2 45554 45559
0 45561 5 1 1 45560
0 45562 7 1 2 45550 45561
0 45563 5 1 1 45562
0 45564 7 1 2 82289 45563
0 45565 5 1 1 45564
0 45566 7 4 2 65487 79020
0 45567 5 3 1 97173
0 45568 7 1 2 97044 97153
0 45569 5 1 1 45568
0 45570 7 1 2 97177 45569
0 45571 5 1 1 45570
0 45572 7 1 2 90908 45571
0 45573 5 1 1 45572
0 45574 7 1 2 45565 45573
0 45575 7 1 2 45543 45574
0 45576 7 1 2 45531 45575
0 45577 5 1 1 45576
0 45578 7 1 2 66578 45577
0 45579 5 1 1 45578
0 45580 7 1 2 45503 45579
0 45581 5 1 1 45580
0 45582 7 1 2 65289 45581
0 45583 5 1 1 45582
0 45584 7 1 2 74934 87960
0 45585 5 1 1 45584
0 45586 7 1 2 60595 45585
0 45587 5 1 1 45586
0 45588 7 1 2 63156 45587
0 45589 5 1 1 45588
0 45590 7 1 2 62750 95565
0 45591 5 1 1 45590
0 45592 7 1 2 74001 45591
0 45593 5 1 1 45592
0 45594 7 1 2 65488 97144
0 45595 7 1 2 45593 45594
0 45596 5 1 1 45595
0 45597 7 1 2 45589 45596
0 45598 5 1 1 45597
0 45599 7 2 2 71128 84515
0 45600 5 1 1 97180
0 45601 7 1 2 45598 97181
0 45602 5 1 1 45601
0 45603 7 1 2 68494 45602
0 45604 7 1 2 45583 45603
0 45605 5 1 1 45604
0 45606 7 1 2 70080 45605
0 45607 7 1 2 45497 45606
0 45608 5 1 1 45607
0 45609 7 1 2 84992 44916
0 45610 5 1 1 45609
0 45611 7 1 2 72469 45610
0 45612 5 1 1 45611
0 45613 7 1 2 84716 87327
0 45614 5 1 1 45613
0 45615 7 1 2 45612 45614
0 45616 5 1 1 45615
0 45617 7 1 2 72372 45616
0 45618 5 1 1 45617
0 45619 7 1 2 82563 88880
0 45620 5 1 1 45619
0 45621 7 1 2 75851 45620
0 45622 5 1 1 45621
0 45623 7 1 2 63549 85118
0 45624 5 1 1 45623
0 45625 7 1 2 45622 45624
0 45626 5 1 1 45625
0 45627 7 1 2 63157 45626
0 45628 5 1 1 45627
0 45629 7 1 2 45618 45628
0 45630 5 1 1 45629
0 45631 7 1 2 91213 45630
0 45632 5 1 1 45631
0 45633 7 1 2 85733 97104
0 45634 5 1 1 45633
0 45635 7 1 2 75626 45634
0 45636 5 1 1 45635
0 45637 7 3 2 68495 91864
0 45638 7 1 2 82577 97182
0 45639 5 1 1 45638
0 45640 7 1 2 45636 45639
0 45641 5 1 1 45640
0 45642 7 1 2 64336 45641
0 45643 5 1 1 45642
0 45644 7 1 2 92952 93521
0 45645 5 1 1 45644
0 45646 7 1 2 45643 45645
0 45647 5 1 1 45646
0 45648 7 1 2 78008 45647
0 45649 5 1 1 45648
0 45650 7 1 2 45632 45649
0 45651 5 1 1 45650
0 45652 7 1 2 63821 45651
0 45653 5 1 1 45652
0 45654 7 2 2 81273 87463
0 45655 7 1 2 81743 91160
0 45656 7 1 2 97185 45655
0 45657 5 1 1 45656
0 45658 7 1 2 45653 45657
0 45659 5 1 1 45658
0 45660 7 1 2 61775 45659
0 45661 5 1 1 45660
0 45662 7 1 2 7981 29202
0 45663 5 1 1 45662
0 45664 7 1 2 65903 45663
0 45665 5 1 1 45664
0 45666 7 1 2 80740 78995
0 45667 5 1 1 45666
0 45668 7 1 2 45665 45667
0 45669 5 1 1 45668
0 45670 7 1 2 64815 45669
0 45671 5 1 1 45670
0 45672 7 1 2 77923 90374
0 45673 5 1 1 45672
0 45674 7 1 2 45671 45673
0 45675 5 1 1 45674
0 45676 7 1 2 64578 45675
0 45677 5 1 1 45676
0 45678 7 1 2 84989 86402
0 45679 5 1 1 45678
0 45680 7 1 2 75806 88934
0 45681 7 1 2 95494 96350
0 45682 7 1 2 45680 45681
0 45683 5 1 1 45682
0 45684 7 1 2 45679 45683
0 45685 7 1 2 45677 45684
0 45686 5 1 1 45685
0 45687 7 1 2 62751 45686
0 45688 5 1 1 45687
0 45689 7 1 2 85741 97131
0 45690 5 1 1 45689
0 45691 7 1 2 45688 45690
0 45692 5 1 1 45691
0 45693 7 1 2 65290 45692
0 45694 5 1 1 45693
0 45695 7 1 2 82416 84789
0 45696 7 1 2 89665 45695
0 45697 5 1 1 45696
0 45698 7 1 2 45694 45697
0 45699 5 1 1 45698
0 45700 7 2 2 70081 84196
0 45701 5 1 1 97187
0 45702 7 1 2 45699 97188
0 45703 5 1 1 45702
0 45704 7 1 2 45661 45703
0 45705 5 1 1 45704
0 45706 7 1 2 70337 45705
0 45707 5 1 1 45706
0 45708 7 2 2 63550 84028
0 45709 5 1 1 97189
0 45710 7 1 2 91129 97133
0 45711 5 1 1 45710
0 45712 7 1 2 64337 91101
0 45713 5 1 1 45712
0 45714 7 1 2 45711 45713
0 45715 5 1 1 45714
0 45716 7 1 2 68496 45715
0 45717 5 1 1 45716
0 45718 7 1 2 45709 45717
0 45719 5 1 1 45718
0 45720 7 1 2 88417 45719
0 45721 5 1 1 45720
0 45722 7 1 2 68497 12127
0 45723 5 1 1 45722
0 45724 7 1 2 75699 86934
0 45725 7 1 2 45723 45724
0 45726 5 1 1 45725
0 45727 7 1 2 74838 81518
0 45728 5 1 1 45727
0 45729 7 1 2 45726 45728
0 45730 7 1 2 45721 45729
0 45731 5 1 1 45730
0 45732 7 1 2 91865 45731
0 45733 5 1 1 45732
0 45734 7 1 2 78935 84412
0 45735 7 1 2 81140 45734
0 45736 7 1 2 92907 45735
0 45737 5 1 1 45736
0 45738 7 1 2 45733 45737
0 45739 5 1 1 45738
0 45740 7 1 2 63822 45739
0 45741 5 1 1 45740
0 45742 7 2 2 81778 74935
0 45743 7 1 2 89691 97191
0 45744 5 1 1 45743
0 45745 7 1 2 45741 45744
0 45746 5 1 1 45745
0 45747 7 1 2 61776 45746
0 45748 5 1 1 45747
0 45749 7 1 2 79355 87987
0 45750 5 1 1 45749
0 45751 7 1 2 73117 93890
0 45752 5 1 1 45751
0 45753 7 1 2 45750 45752
0 45754 5 1 1 45753
0 45755 7 1 2 83107 45754
0 45756 5 1 1 45755
0 45757 7 1 2 64338 78161
0 45758 5 1 1 45757
0 45759 7 1 2 93891 45758
0 45760 5 1 1 45759
0 45761 7 2 2 85772 45760
0 45762 5 1 1 97193
0 45763 7 1 2 66074 97194
0 45764 5 1 1 45763
0 45765 7 1 2 93529 45764
0 45766 7 1 2 45756 45765
0 45767 5 1 1 45766
0 45768 7 1 2 70904 45767
0 45769 5 1 1 45768
0 45770 7 1 2 80524 79027
0 45771 5 1 1 45770
0 45772 7 1 2 77799 93641
0 45773 5 1 1 45772
0 45774 7 1 2 77952 45773
0 45775 5 1 1 45774
0 45776 7 1 2 74035 45775
0 45777 5 1 1 45776
0 45778 7 2 2 64339 70082
0 45779 5 1 1 97195
0 45780 7 1 2 85375 97196
0 45781 5 1 1 45780
0 45782 7 1 2 70083 97190
0 45783 5 1 1 45782
0 45784 7 1 2 64340 93563
0 45785 5 1 1 45784
0 45786 7 1 2 45783 45785
0 45787 5 1 1 45786
0 45788 7 1 2 88418 45787
0 45789 5 1 1 45788
0 45790 7 1 2 45781 45789
0 45791 7 1 2 45777 45790
0 45792 5 1 1 45791
0 45793 7 1 2 63823 45792
0 45794 5 1 1 45793
0 45795 7 1 2 45771 45794
0 45796 7 1 2 45769 45795
0 45797 5 1 1 45796
0 45798 7 1 2 61777 45797
0 45799 5 1 1 45798
0 45800 7 3 2 77438 83559
0 45801 7 1 2 97186 97197
0 45802 7 1 2 88642 45801
0 45803 5 1 1 45802
0 45804 7 1 2 45799 45803
0 45805 5 1 1 45804
0 45806 7 1 2 75627 45805
0 45807 5 1 1 45806
0 45808 7 2 2 77924 91866
0 45809 7 1 2 74036 97200
0 45810 5 1 1 45809
0 45811 7 2 2 90731 93203
0 45812 5 1 1 97202
0 45813 7 2 2 77483 97203
0 45814 5 1 1 97204
0 45815 7 1 2 75628 82186
0 45816 5 1 1 45815
0 45817 7 1 2 45814 45816
0 45818 5 1 1 45817
0 45819 7 1 2 73118 45818
0 45820 5 1 1 45819
0 45821 7 1 2 45810 45820
0 45822 5 1 1 45821
0 45823 7 1 2 84516 45822
0 45824 5 1 1 45823
0 45825 7 2 2 87358 97192
0 45826 7 1 2 83560 97206
0 45827 5 1 1 45826
0 45828 7 1 2 45824 45827
0 45829 5 1 1 45828
0 45830 7 1 2 72502 45829
0 45831 5 1 1 45830
0 45832 7 6 2 83449 87826
0 45833 5 2 1 97208
0 45834 7 1 2 10948 97107
0 45835 5 1 1 45834
0 45836 7 1 2 64341 45835
0 45837 5 1 1 45836
0 45838 7 1 2 87967 45837
0 45839 5 1 1 45838
0 45840 7 1 2 64579 45839
0 45841 5 1 1 45840
0 45842 7 1 2 29839 45841
0 45843 5 1 1 45842
0 45844 7 1 2 72373 45843
0 45845 5 1 1 45844
0 45846 7 1 2 71129 79595
0 45847 7 1 2 87468 45846
0 45848 5 1 1 45847
0 45849 7 1 2 86551 45848
0 45850 5 1 1 45849
0 45851 7 1 2 68498 83329
0 45852 7 1 2 45850 45851
0 45853 5 1 1 45852
0 45854 7 1 2 45845 45853
0 45855 5 1 1 45854
0 45856 7 1 2 97209 45855
0 45857 5 1 1 45856
0 45858 7 1 2 45831 45857
0 45859 7 1 2 45807 45858
0 45860 7 1 2 45748 45859
0 45861 5 1 1 45860
0 45862 7 1 2 70373 45861
0 45863 5 1 1 45862
0 45864 7 1 2 67731 95433
0 45865 5 1 1 45864
0 45866 7 1 2 62387 85779
0 45867 5 1 1 45866
0 45868 7 1 2 45865 45867
0 45869 5 1 1 45868
0 45870 7 1 2 84871 45869
0 45871 5 1 1 45870
0 45872 7 1 2 77636 94826
0 45873 5 1 1 45872
0 45874 7 1 2 45871 45873
0 45875 5 1 1 45874
0 45876 7 1 2 65489 45875
0 45877 5 1 1 45876
0 45878 7 1 2 80043 88263
0 45879 5 1 1 45878
0 45880 7 1 2 45877 45879
0 45881 5 1 1 45880
0 45882 7 1 2 63158 45881
0 45883 5 1 1 45882
0 45884 7 1 2 88237 96046
0 45885 7 1 2 95341 45884
0 45886 5 1 1 45885
0 45887 7 1 2 45883 45886
0 45888 5 1 1 45887
0 45889 7 1 2 78671 45888
0 45890 5 1 1 45889
0 45891 7 1 2 65490 83120
0 45892 7 1 2 85931 45891
0 45893 5 1 1 45892
0 45894 7 1 2 78952 97100
0 45895 5 1 1 45894
0 45896 7 1 2 64816 93610
0 45897 5 1 1 45896
0 45898 7 1 2 45895 45897
0 45899 5 1 1 45898
0 45900 7 1 2 73529 88861
0 45901 7 1 2 45899 45900
0 45902 5 1 1 45901
0 45903 7 1 2 45893 45902
0 45904 5 1 1 45903
0 45905 7 1 2 84517 45904
0 45906 5 1 1 45905
0 45907 7 1 2 45890 45906
0 45908 7 1 2 77097 97040
0 45909 5 1 1 45908
0 45910 7 2 2 70421 76100
0 45911 5 1 1 97216
0 45912 7 1 2 64342 79157
0 45913 7 1 2 45911 45912
0 45914 5 1 1 45913
0 45915 7 1 2 45909 45914
0 45916 5 1 1 45915
0 45917 7 1 2 61778 45916
0 45918 5 1 1 45917
0 45919 7 1 2 95604 45918
0 45920 5 1 1 45919
0 45921 7 1 2 84872 45920
0 45922 5 1 1 45921
0 45923 7 1 2 73136 82273
0 45924 5 2 1 45923
0 45925 7 1 2 64343 97218
0 45926 5 1 1 45925
0 45927 7 1 2 70292 89667
0 45928 5 1 1 45927
0 45929 7 1 2 83139 45928
0 45930 5 1 1 45929
0 45931 7 1 2 45926 45930
0 45932 5 1 1 45931
0 45933 7 1 2 94827 45932
0 45934 5 1 1 45933
0 45935 7 1 2 45922 45934
0 45936 5 1 1 45935
0 45937 7 1 2 65491 45936
0 45938 5 1 1 45937
0 45939 7 1 2 73537 73196
0 45940 5 1 1 45939
0 45941 7 1 2 74037 45940
0 45942 5 1 1 45941
0 45943 7 1 2 72838 45942
0 45944 5 1 1 45943
0 45945 7 1 2 67732 45944
0 45946 5 1 1 45945
0 45947 7 1 2 88169 45946
0 45948 5 1 1 45947
0 45949 7 1 2 81109 86386
0 45950 7 1 2 45948 45949
0 45951 5 1 1 45950
0 45952 7 1 2 45938 45951
0 45953 5 1 1 45952
0 45954 7 1 2 63159 45953
0 45955 5 1 1 45954
0 45956 7 2 2 78855 84873
0 45957 5 1 1 97220
0 45958 7 1 2 86002 94095
0 45959 5 1 1 45958
0 45960 7 1 2 45957 45959
0 45961 5 1 1 45960
0 45962 7 1 2 64344 45961
0 45963 5 1 1 45962
0 45964 7 1 2 74307 94365
0 45965 5 1 1 45964
0 45966 7 1 2 95095 45965
0 45967 5 1 1 45966
0 45968 7 1 2 63160 45967
0 45969 5 1 1 45968
0 45970 7 1 2 65744 97221
0 45971 5 1 1 45970
0 45972 7 1 2 62752 78408
0 45973 7 1 2 94828 45972
0 45974 5 1 1 45973
0 45975 7 1 2 45971 45974
0 45976 7 1 2 45969 45975
0 45977 7 1 2 45963 45976
0 45978 5 1 1 45977
0 45979 7 1 2 65492 45978
0 45980 5 1 1 45979
0 45981 7 1 2 66579 75692
0 45982 7 1 2 96193 45981
0 45983 7 1 2 852 45982
0 45984 5 1 1 45983
0 45985 7 1 2 45980 45984
0 45986 5 1 1 45985
0 45987 7 1 2 71833 45986
0 45988 5 1 1 45987
0 45989 7 1 2 9276 26524
0 45990 5 1 1 45989
0 45991 7 1 2 65745 45990
0 45992 5 1 1 45991
0 45993 7 1 2 75423 84717
0 45994 5 1 1 45993
0 45995 7 1 2 45992 45994
0 45996 5 1 1 45995
0 45997 7 1 2 64345 45996
0 45998 5 1 1 45997
0 45999 7 1 2 82187 76535
0 46000 5 1 1 45999
0 46001 7 1 2 45998 46000
0 46002 5 1 1 46001
0 46003 7 1 2 84518 46002
0 46004 5 1 1 46003
0 46005 7 1 2 70338 83039
0 46006 5 1 1 46005
0 46007 7 1 2 78860 46006
0 46008 5 1 1 46007
0 46009 7 1 2 91141 46008
0 46010 5 1 1 46009
0 46011 7 1 2 46004 46010
0 46012 5 1 1 46011
0 46013 7 1 2 72023 46012
0 46014 5 1 1 46013
0 46015 7 1 2 78792 21643
0 46016 5 1 1 46015
0 46017 7 1 2 87926 88190
0 46018 7 1 2 46016 46017
0 46019 5 1 1 46018
0 46020 7 1 2 46014 46019
0 46021 7 1 2 45988 46020
0 46022 5 1 1 46021
0 46023 7 1 2 72374 46022
0 46024 5 1 1 46023
0 46025 7 1 2 45955 46024
0 46026 7 1 2 45907 46025
0 46027 5 1 1 46026
0 46028 7 1 2 71582 46027
0 46029 5 1 1 46028
0 46030 7 1 2 93530 45762
0 46031 5 1 1 46030
0 46032 7 1 2 74038 46031
0 46033 5 1 1 46032
0 46034 7 1 2 64346 80128
0 46035 7 1 2 85835 46034
0 46036 5 1 1 46035
0 46037 7 1 2 46033 46036
0 46038 5 1 1 46037
0 46039 7 1 2 75629 46038
0 46040 5 1 1 46039
0 46041 7 1 2 62388 97205
0 46042 5 1 1 46041
0 46043 7 1 2 64817 77105
0 46044 5 1 1 46043
0 46045 7 1 2 68499 79421
0 46046 7 1 2 46044 46045
0 46047 5 1 1 46046
0 46048 7 1 2 91867 95495
0 46049 7 1 2 46047 46048
0 46050 5 1 1 46049
0 46051 7 1 2 46042 46050
0 46052 5 1 1 46051
0 46053 7 1 2 63824 46052
0 46054 5 1 1 46053
0 46055 7 1 2 46040 46054
0 46056 5 1 1 46055
0 46057 7 1 2 61779 46056
0 46058 5 1 1 46057
0 46059 7 1 2 73119 85947
0 46060 5 1 1 46059
0 46061 7 1 2 77948 46060
0 46062 5 1 1 46061
0 46063 7 2 2 84197 79546
0 46064 5 1 1 97222
0 46065 7 1 2 46062 97223
0 46066 5 1 1 46065
0 46067 7 1 2 46058 46066
0 46068 5 1 1 46067
0 46069 7 1 2 70848 46068
0 46070 5 1 1 46069
0 46071 7 1 2 80281 84519
0 46072 5 1 1 46071
0 46073 7 1 2 83953 79547
0 46074 5 1 1 46073
0 46075 7 1 2 46072 46074
0 46076 5 1 1 46075
0 46077 7 2 2 68500 88030
0 46078 7 1 2 46076 97224
0 46079 5 1 1 46078
0 46080 7 1 2 83287 92150
0 46081 7 1 2 94303 46080
0 46082 5 1 1 46081
0 46083 7 1 2 46079 46082
0 46084 5 1 1 46083
0 46085 7 1 2 64347 46084
0 46086 5 1 1 46085
0 46087 7 1 2 77925 94851
0 46088 5 1 1 46087
0 46089 7 1 2 83982 85002
0 46090 5 1 1 46089
0 46091 7 1 2 46088 46090
0 46092 5 1 1 46091
0 46093 7 1 2 77098 46092
0 46094 5 1 1 46093
0 46095 7 1 2 46086 46094
0 46096 5 1 1 46095
0 46097 7 1 2 65493 46096
0 46098 5 1 1 46097
0 46099 7 1 2 77926 78088
0 46100 7 1 2 87243 46099
0 46101 5 1 1 46100
0 46102 7 1 2 79471 91324
0 46103 7 1 2 97225 46102
0 46104 5 1 1 46103
0 46105 7 1 2 46101 46104
0 46106 5 1 1 46105
0 46107 7 1 2 84520 46106
0 46108 5 1 1 46107
0 46109 7 1 2 46098 46108
0 46110 7 1 2 46070 46109
0 46111 5 1 1 46110
0 46112 7 1 2 88655 46111
0 46113 5 1 1 46112
0 46114 7 1 2 97201 97219
0 46115 5 1 1 46114
0 46116 7 1 2 74961 86935
0 46117 5 1 1 46116
0 46118 7 1 2 82190 46117
0 46119 5 1 1 46118
0 46120 7 1 2 64580 46119
0 46121 5 1 1 46120
0 46122 7 1 2 93565 46121
0 46123 5 1 1 46122
0 46124 7 1 2 75630 46123
0 46125 5 1 1 46124
0 46126 7 1 2 64581 97183
0 46127 5 1 1 46126
0 46128 7 1 2 45812 46127
0 46129 5 1 1 46128
0 46130 7 1 2 87438 46129
0 46131 5 1 1 46130
0 46132 7 1 2 46125 46131
0 46133 5 1 1 46132
0 46134 7 1 2 64818 46133
0 46135 5 1 1 46134
0 46136 7 1 2 46115 46135
0 46137 5 1 1 46136
0 46138 7 1 2 84521 46137
0 46139 5 1 1 46138
0 46140 7 1 2 87777 97207
0 46141 5 1 1 46140
0 46142 7 1 2 46139 46141
0 46143 5 1 1 46142
0 46144 7 1 2 95650 46143
0 46145 5 1 1 46144
0 46146 7 1 2 87359 91868
0 46147 5 1 1 46146
0 46148 7 1 2 91082 95417
0 46149 5 1 1 46148
0 46150 7 1 2 46147 46149
0 46151 5 1 1 46150
0 46152 7 1 2 84522 46151
0 46153 5 1 1 46152
0 46154 7 1 2 74936 83450
0 46155 7 1 2 84384 46154
0 46156 5 1 1 46155
0 46157 7 1 2 46153 46156
0 46158 5 1 1 46157
0 46159 7 1 2 63551 74076
0 46160 7 1 2 46158 46159
0 46161 5 1 1 46160
0 46162 7 1 2 72162 93823
0 46163 5 1 1 46162
0 46164 7 1 2 76651 88286
0 46165 5 1 1 46164
0 46166 7 1 2 46163 46165
0 46167 5 1 1 46166
0 46168 7 1 2 65494 46167
0 46169 5 1 1 46168
0 46170 7 1 2 85763 87439
0 46171 5 1 1 46170
0 46172 7 1 2 46169 46171
0 46173 5 1 1 46172
0 46174 7 1 2 81996 79356
0 46175 7 1 2 46173 46174
0 46176 5 1 1 46175
0 46177 7 1 2 46161 46176
0 46178 5 1 1 46177
0 46179 7 1 2 70339 46178
0 46180 5 1 1 46179
0 46181 7 2 2 71730 76523
0 46182 5 2 1 97226
0 46183 7 1 2 62753 97228
0 46184 5 1 1 46183
0 46185 7 1 2 68111 46184
0 46186 5 1 1 46185
0 46187 7 1 2 81997 93843
0 46188 7 1 2 46186 46187
0 46189 5 1 1 46188
0 46190 7 1 2 74778 90264
0 46191 5 1 1 46190
0 46192 7 1 2 73530 46191
0 46193 5 1 1 46192
0 46194 7 1 2 84913 46193
0 46195 5 1 1 46194
0 46196 7 1 2 83631 77927
0 46197 7 1 2 46195 46196
0 46198 5 1 1 46197
0 46199 7 1 2 46189 46198
0 46200 5 1 1 46199
0 46201 7 1 2 65495 46200
0 46202 5 1 1 46201
0 46203 7 1 2 46180 46202
0 46204 5 1 1 46203
0 46205 7 1 2 72503 46204
0 46206 5 1 1 46205
0 46207 7 1 2 64819 91437
0 46208 5 1 1 46207
0 46209 7 1 2 66075 97166
0 46210 5 1 1 46209
0 46211 7 1 2 46208 46210
0 46212 5 1 1 46211
0 46213 7 1 2 64582 46212
0 46214 5 1 1 46213
0 46215 7 1 2 72786 91443
0 46216 5 1 1 46215
0 46217 7 1 2 46214 46216
0 46218 5 1 1 46217
0 46219 7 1 2 87683 46218
0 46220 5 1 1 46219
0 46221 7 1 2 63552 84651
0 46222 5 1 1 46221
0 46223 7 1 2 75852 79174
0 46224 5 1 1 46223
0 46225 7 1 2 46222 46224
0 46226 5 1 1 46225
0 46227 7 1 2 62754 46226
0 46228 5 1 1 46227
0 46229 7 1 2 64583 72869
0 46230 5 1 1 46229
0 46231 7 1 2 72245 46230
0 46232 5 1 1 46231
0 46233 7 1 2 75700 89919
0 46234 7 1 2 46232 46233
0 46235 5 1 1 46234
0 46236 7 1 2 75853 91553
0 46237 5 1 1 46236
0 46238 7 1 2 75854 82290
0 46239 5 1 1 46238
0 46240 7 1 2 30807 46239
0 46241 5 1 1 46240
0 46242 7 1 2 76033 46241
0 46243 5 1 1 46242
0 46244 7 1 2 46237 46243
0 46245 7 1 2 46235 46244
0 46246 7 1 2 46228 46245
0 46247 5 1 1 46246
0 46248 7 1 2 63161 46247
0 46249 5 1 1 46248
0 46250 7 1 2 78889 88788
0 46251 5 1 1 46250
0 46252 7 1 2 75631 82417
0 46253 5 1 1 46252
0 46254 7 1 2 29898 46253
0 46255 7 1 2 46251 46254
0 46256 5 1 1 46255
0 46257 7 1 2 63553 46256
0 46258 5 1 1 46257
0 46259 7 1 2 46249 46258
0 46260 7 1 2 46220 46259
0 46261 5 1 1 46260
0 46262 7 2 2 65496 84523
0 46263 5 1 1 97230
0 46264 7 1 2 46261 97231
0 46265 5 1 1 46264
0 46266 7 1 2 46206 46265
0 46267 7 1 2 46145 46266
0 46268 7 1 2 46113 46267
0 46269 7 1 2 46029 46268
0 46270 7 1 2 45863 46269
0 46271 7 1 2 45707 46270
0 46272 7 1 2 45608 46271
0 46273 7 1 2 45333 46272
0 46274 7 1 2 44758 46273
0 46275 5 1 1 46274
0 46276 7 1 2 66892 46275
0 46277 5 1 1 46276
0 46278 7 1 2 65497 97068
0 46279 5 1 1 46278
0 46280 7 1 2 61780 46279
0 46281 5 1 1 46280
0 46282 7 1 2 79719 46281
0 46283 7 1 2 97070 46282
0 46284 5 1 1 46283
0 46285 7 1 2 46277 46284
0 46286 5 1 1 46285
0 46287 7 1 2 65612 46286
0 46288 5 1 1 46287
0 46289 7 1 2 69006 46288
0 46290 7 1 2 44509 46289
0 46291 5 1 1 46290
0 46292 7 1 2 79720 87019
0 46293 5 1 1 46292
0 46294 7 2 2 73421 96961
0 46295 7 1 2 95904 97232
0 46296 7 1 2 96750 46295
0 46297 5 1 1 46296
0 46298 7 1 2 46293 46297
0 46299 5 1 1 46298
0 46300 7 1 2 83060 46299
0 46301 5 1 1 46300
0 46302 7 2 2 76328 72375
0 46303 5 3 1 97234
0 46304 7 1 2 75237 97235
0 46305 5 1 1 46304
0 46306 7 1 2 70340 90412
0 46307 5 1 1 46306
0 46308 7 1 2 70374 90417
0 46309 5 1 1 46308
0 46310 7 1 2 72772 94662
0 46311 5 1 1 46310
0 46312 7 1 2 76878 46311
0 46313 7 1 2 46309 46312
0 46314 7 1 2 46307 46313
0 46315 5 1 1 46314
0 46316 7 1 2 63162 46315
0 46317 5 1 1 46316
0 46318 7 1 2 63163 90308
0 46319 5 1 1 46318
0 46320 7 1 2 63164 77637
0 46321 5 1 1 46320
0 46322 7 1 2 59395 46321
0 46323 5 1 1 46322
0 46324 7 1 2 71834 87011
0 46325 7 1 2 46323 46324
0 46326 5 2 1 46325
0 46327 7 1 2 46319 97239
0 46328 5 1 1 46327
0 46329 7 1 2 72376 46328
0 46330 5 1 1 46329
0 46331 7 1 2 90662 90973
0 46332 5 1 1 46331
0 46333 7 1 2 90175 46332
0 46334 7 1 2 46330 46333
0 46335 7 1 2 46317 46334
0 46336 5 1 1 46335
0 46337 7 1 2 46305 46336
0 46338 5 1 1 46337
0 46339 7 1 2 67103 1261
0 46340 5 1 1 46339
0 46341 7 1 2 67373 94540
0 46342 5 1 1 46341
0 46343 7 1 2 46340 46342
0 46344 5 1 1 46343
0 46345 7 1 2 62755 46344
0 46346 5 1 1 46345
0 46347 7 1 2 67733 95861
0 46348 5 1 1 46347
0 46349 7 1 2 46346 46348
0 46350 5 2 1 46349
0 46351 7 1 2 72504 97241
0 46352 5 1 1 46351
0 46353 7 1 2 72024 95434
0 46354 5 1 1 46353
0 46355 7 1 2 70849 70540
0 46356 5 1 1 46355
0 46357 7 1 2 46354 46356
0 46358 5 1 1 46357
0 46359 7 1 2 62756 46358
0 46360 5 1 1 46359
0 46361 7 1 2 90354 88497
0 46362 5 1 1 46361
0 46363 7 1 2 46360 46362
0 46364 5 1 1 46363
0 46365 7 1 2 72377 46364
0 46366 5 1 1 46365
0 46367 7 1 2 70084 70541
0 46368 5 1 1 46367
0 46369 7 1 2 74921 46368
0 46370 7 1 2 5043 46369
0 46371 7 1 2 46366 46370
0 46372 7 1 2 46352 46371
0 46373 5 1 1 46372
0 46374 7 1 2 68112 46373
0 46375 5 1 1 46374
0 46376 7 1 2 46338 46375
0 46377 5 1 1 46376
0 46378 7 1 2 92838 46377
0 46379 5 1 1 46378
0 46380 7 1 2 46301 46379
0 46381 5 1 1 46380
0 46382 7 1 2 68501 46381
0 46383 5 1 1 46382
0 46384 7 1 2 66580 95382
0 46385 5 1 1 46384
0 46386 7 1 2 78470 93489
0 46387 5 1 1 46386
0 46388 7 1 2 67734 91565
0 46389 7 1 2 97058 46388
0 46390 5 1 1 46389
0 46391 7 1 2 65291 46390
0 46392 5 1 1 46391
0 46393 7 1 2 46387 46392
0 46394 5 1 1 46393
0 46395 7 1 2 64584 46394
0 46396 5 1 1 46395
0 46397 7 1 2 90557 97162
0 46398 5 1 1 46397
0 46399 7 1 2 65292 75893
0 46400 7 1 2 46398 46399
0 46401 5 1 1 46400
0 46402 7 1 2 46396 46401
0 46403 5 1 1 46402
0 46404 7 1 2 70850 46403
0 46405 5 1 1 46404
0 46406 7 1 2 76733 44512
0 46407 5 1 1 46406
0 46408 7 1 2 94335 46407
0 46409 5 1 1 46408
0 46410 7 1 2 65293 77099
0 46411 5 1 1 46410
0 46412 7 1 2 80662 91083
0 46413 5 1 1 46412
0 46414 7 1 2 46411 46413
0 46415 5 1 1 46414
0 46416 7 1 2 79592 46415
0 46417 5 1 1 46416
0 46418 7 1 2 75956 83832
0 46419 5 1 1 46418
0 46420 7 1 2 60178 46419
0 46421 5 1 1 46420
0 46422 7 1 2 77100 95345
0 46423 7 1 2 46421 46422
0 46424 5 1 1 46423
0 46425 7 1 2 46417 46424
0 46426 7 1 2 46409 46425
0 46427 7 1 2 46405 46426
0 46428 5 1 1 46427
0 46429 7 1 2 72378 46428
0 46430 5 1 1 46429
0 46431 7 1 2 88583 97111
0 46432 5 1 1 46431
0 46433 7 1 2 95644 46432
0 46434 5 1 1 46433
0 46435 7 1 2 64348 46434
0 46436 5 1 1 46435
0 46437 7 1 2 66076 94789
0 46438 5 1 1 46437
0 46439 7 1 2 90456 46438
0 46440 5 1 1 46439
0 46441 7 1 2 71583 46440
0 46442 5 1 1 46441
0 46443 7 1 2 60401 91278
0 46444 5 1 1 46443
0 46445 7 1 2 70341 70851
0 46446 7 1 2 46444 46445
0 46447 5 1 1 46446
0 46448 7 1 2 46442 46447
0 46449 7 1 2 46436 46448
0 46450 5 1 1 46449
0 46451 7 1 2 63165 46450
0 46452 5 1 1 46451
0 46453 7 1 2 77197 77811
0 46454 5 1 1 46453
0 46455 7 1 2 72727 77817
0 46456 5 1 1 46455
0 46457 7 1 2 77173 46456
0 46458 5 1 1 46457
0 46459 7 1 2 65294 46458
0 46460 5 1 1 46459
0 46461 7 1 2 46454 46460
0 46462 5 1 1 46461
0 46463 7 1 2 82525 46462
0 46464 5 1 1 46463
0 46465 7 1 2 76372 85832
0 46466 5 1 1 46465
0 46467 7 1 2 81603 93450
0 46468 5 1 1 46467
0 46469 7 1 2 65498 46468
0 46470 5 1 1 46469
0 46471 7 1 2 76754 91444
0 46472 7 1 2 97145 46471
0 46473 5 1 1 46472
0 46474 7 1 2 46470 46473
0 46475 7 1 2 46466 46474
0 46476 7 1 2 90558 88385
0 46477 5 1 1 46476
0 46478 7 1 2 62757 80081
0 46479 7 1 2 95648 46478
0 46480 7 1 2 46477 46479
0 46481 5 1 1 46480
0 46482 7 1 2 73120 97146
0 46483 5 2 1 46482
0 46484 7 1 2 70375 83330
0 46485 5 2 1 46484
0 46486 7 1 2 97243 97245
0 46487 5 1 1 46486
0 46488 7 1 2 64820 90283
0 46489 5 1 1 46488
0 46490 7 1 2 68113 46489
0 46491 5 2 1 46490
0 46492 7 1 2 71584 97247
0 46493 5 1 1 46492
0 46494 7 1 2 84660 88250
0 46495 5 1 1 46494
0 46496 7 1 2 70852 46495
0 46497 5 1 1 46496
0 46498 7 1 2 46493 46497
0 46499 5 1 1 46498
0 46500 7 1 2 46487 46499
0 46501 5 1 1 46500
0 46502 7 2 2 72379 97134
0 46503 7 1 2 94336 97249
0 46504 5 1 1 46503
0 46505 7 1 2 70853 88248
0 46506 7 1 2 78111 46505
0 46507 5 1 1 46506
0 46508 7 1 2 46504 46507
0 46509 5 1 1 46508
0 46510 7 1 2 70376 46509
0 46511 5 1 1 46510
0 46512 7 1 2 46501 46511
0 46513 7 1 2 46481 46512
0 46514 7 1 2 46475 46513
0 46515 7 1 2 46464 46514
0 46516 7 1 2 46452 46515
0 46517 7 1 2 46430 46516
0 46518 7 1 2 46385 46517
0 46519 5 1 1 46518
0 46520 7 1 2 63554 46519
0 46521 5 1 1 46520
0 46522 7 1 2 63166 88354
0 46523 5 1 1 46522
0 46524 7 1 2 80654 93754
0 46525 5 1 1 46524
0 46526 7 1 2 46523 46525
0 46527 5 1 1 46526
0 46528 7 1 2 75632 46527
0 46529 5 1 1 46528
0 46530 7 1 2 88249 94857
0 46531 5 2 1 46530
0 46532 7 1 2 46529 97251
0 46533 5 1 1 46532
0 46534 7 1 2 88813 46533
0 46535 5 1 1 46534
0 46536 7 1 2 60596 87248
0 46537 5 7 1 46536
0 46538 7 2 2 63167 97253
0 46539 7 1 2 76912 97260
0 46540 5 1 1 46539
0 46541 7 2 2 86602 91869
0 46542 5 1 1 97262
0 46543 7 1 2 69374 97263
0 46544 5 1 1 46543
0 46545 7 1 2 46540 46544
0 46546 5 1 1 46545
0 46547 7 1 2 90503 46546
0 46548 5 1 1 46547
0 46549 7 1 2 80304 90294
0 46550 5 1 1 46549
0 46551 7 1 2 80269 46550
0 46552 5 1 1 46551
0 46553 7 1 2 65499 46552
0 46554 5 1 1 46553
0 46555 7 2 2 90781 93596
0 46556 5 2 1 97264
0 46557 7 1 2 90877 97266
0 46558 5 2 1 46557
0 46559 7 1 2 87580 97268
0 46560 7 1 2 46554 46559
0 46561 7 1 2 46548 46560
0 46562 7 1 2 46535 46561
0 46563 5 1 1 46562
0 46564 7 1 2 82578 46563
0 46565 5 1 1 46564
0 46566 7 1 2 71897 84602
0 46567 5 2 1 46566
0 46568 7 1 2 65500 97270
0 46569 5 1 1 46568
0 46570 7 2 2 69074 91289
0 46571 7 1 2 83884 97272
0 46572 5 2 1 46571
0 46573 7 1 2 74511 90504
0 46574 5 2 1 46573
0 46575 7 1 2 72423 97095
0 46576 5 1 1 46575
0 46577 7 2 2 97276 46576
0 46578 7 1 2 71130 79158
0 46579 5 1 1 46578
0 46580 7 1 2 97278 46579
0 46581 5 1 1 46580
0 46582 7 1 2 63168 46581
0 46583 5 1 1 46582
0 46584 7 1 2 97274 46583
0 46585 5 1 1 46584
0 46586 7 1 2 66581 46585
0 46587 5 1 1 46586
0 46588 7 1 2 46569 46587
0 46589 5 1 1 46588
0 46590 7 1 2 71585 46589
0 46591 5 1 1 46590
0 46592 7 1 2 90386 91004
0 46593 5 1 1 46592
0 46594 7 1 2 60597 46593
0 46595 5 1 1 46594
0 46596 7 1 2 64821 46595
0 46597 5 1 1 46596
0 46598 7 1 2 65295 94858
0 46599 5 1 1 46598
0 46600 7 1 2 65501 71934
0 46601 5 1 1 46600
0 46602 7 1 2 46599 46601
0 46603 7 1 2 46597 46602
0 46604 5 1 1 46603
0 46605 7 1 2 63169 46604
0 46606 5 1 1 46605
0 46607 7 2 2 60402 81701
0 46608 5 1 1 97280
0 46609 7 1 2 65502 46608
0 46610 5 1 1 46609
0 46611 7 1 2 63170 74430
0 46612 5 1 1 46611
0 46613 7 1 2 97277 46612
0 46614 5 1 1 46613
0 46615 7 1 2 69739 91870
0 46616 7 1 2 46614 46615
0 46617 5 1 1 46616
0 46618 7 1 2 46610 46617
0 46619 7 1 2 46606 46618
0 46620 5 1 1 46619
0 46621 7 1 2 70854 46620
0 46622 5 1 1 46621
0 46623 7 1 2 81702 97279
0 46624 5 1 1 46623
0 46625 7 1 2 63171 46624
0 46626 5 1 1 46625
0 46627 7 1 2 97275 46626
0 46628 5 1 1 46627
0 46629 7 1 2 91214 46628
0 46630 5 1 1 46629
0 46631 7 1 2 60598 87581
0 46632 5 2 1 46631
0 46633 7 6 2 80282 97282
0 46634 5 1 1 97284
0 46635 7 1 2 97269 46634
0 46636 5 1 1 46635
0 46637 7 2 2 70342 74077
0 46638 5 1 1 97290
0 46639 7 1 2 46636 97291
0 46640 5 1 1 46639
0 46641 7 1 2 18214 46542
0 46642 5 1 1 46641
0 46643 7 1 2 90878 46642
0 46644 5 1 1 46643
0 46645 7 1 2 74937 95597
0 46646 5 1 1 46645
0 46647 7 1 2 26700 46646
0 46648 5 1 1 46647
0 46649 7 1 2 71586 46648
0 46650 5 1 1 46649
0 46651 7 1 2 63172 93594
0 46652 5 1 1 46651
0 46653 7 1 2 91215 91325
0 46654 5 1 1 46653
0 46655 7 1 2 46652 46654
0 46656 7 1 2 46650 46655
0 46657 7 1 2 46644 46656
0 46658 5 1 1 46657
0 46659 7 1 2 69198 82784
0 46660 5 1 1 46659
0 46661 7 1 2 46658 46660
0 46662 5 1 1 46661
0 46663 7 1 2 46640 46662
0 46664 7 1 2 46630 46663
0 46665 7 1 2 46622 46664
0 46666 7 1 2 46591 46665
0 46667 7 1 2 46565 46666
0 46668 7 1 2 46521 46667
0 46669 5 1 1 46668
0 46670 7 1 2 68761 46669
0 46671 5 1 1 46670
0 46672 7 1 2 70210 96356
0 46673 5 1 1 46672
0 46674 7 1 2 65296 46673
0 46675 5 1 1 46674
0 46676 7 1 2 70085 90909
0 46677 5 1 1 46676
0 46678 7 1 2 46675 46677
0 46679 5 1 1 46678
0 46680 7 1 2 63173 46679
0 46681 5 1 1 46680
0 46682 7 1 2 65297 90522
0 46683 5 1 1 46682
0 46684 7 1 2 79058 90516
0 46685 5 1 1 46684
0 46686 7 1 2 65503 46685
0 46687 5 1 1 46686
0 46688 7 1 2 46683 46687
0 46689 7 1 2 46681 46688
0 46690 5 1 1 46689
0 46691 7 1 2 68762 46690
0 46692 5 1 1 46691
0 46693 7 1 2 85149 46692
0 46694 5 1 1 46693
0 46695 7 1 2 85932 46694
0 46696 5 1 1 46695
0 46697 7 1 2 63825 89472
0 46698 5 1 1 46697
0 46699 7 1 2 46696 46698
0 46700 7 1 2 46671 46699
0 46701 5 1 1 46700
0 46702 7 1 2 86759 46701
0 46703 5 1 1 46702
0 46704 7 1 2 46383 46703
0 46705 5 1 1 46704
0 46706 7 1 2 66749 46705
0 46707 5 1 1 46706
0 46708 7 1 2 70855 89196
0 46709 5 1 1 46708
0 46710 7 1 2 89209 46709
0 46711 5 1 1 46710
0 46712 7 1 2 72505 46711
0 46713 5 1 1 46712
0 46714 7 1 2 91427 46713
0 46715 5 1 1 46714
0 46716 7 1 2 90572 46715
0 46717 5 1 1 46716
0 46718 7 1 2 82579 90505
0 46719 5 1 1 46718
0 46720 7 1 2 97066 46719
0 46721 5 2 1 46720
0 46722 7 1 2 88474 97292
0 46723 5 1 1 46722
0 46724 7 1 2 71525 96354
0 46725 7 1 2 46723 46724
0 46726 7 1 2 96358 46725
0 46727 5 1 1 46726
0 46728 7 1 2 61607 46727
0 46729 5 1 1 46728
0 46730 7 1 2 69313 90590
0 46731 5 1 1 46730
0 46732 7 1 2 63174 89028
0 46733 7 1 2 46731 46732
0 46734 7 1 2 46729 46733
0 46735 5 1 1 46734
0 46736 7 1 2 89194 88584
0 46737 5 1 1 46736
0 46738 7 1 2 60599 1333
0 46739 7 1 2 46737 46738
0 46740 7 1 2 90481 46739
0 46741 5 1 1 46740
0 46742 7 1 2 67735 46741
0 46743 5 1 1 46742
0 46744 7 1 2 89853 91509
0 46745 7 1 2 89190 46744
0 46746 5 1 1 46745
0 46747 7 1 2 62758 78490
0 46748 5 2 1 46747
0 46749 7 1 2 66582 97294
0 46750 7 1 2 46746 46749
0 46751 5 1 1 46750
0 46752 7 1 2 68114 46751
0 46753 7 1 2 46743 46752
0 46754 5 1 1 46753
0 46755 7 1 2 46735 46754
0 46756 5 1 1 46755
0 46757 7 1 2 46717 46756
0 46758 5 1 1 46757
0 46759 7 1 2 68502 46758
0 46760 5 1 1 46759
0 46761 7 1 2 85457 20301
0 46762 5 1 1 46761
0 46763 7 1 2 89293 93168
0 46764 5 1 1 46763
0 46765 7 1 2 90782 46764
0 46766 5 1 1 46765
0 46767 7 1 2 7340 74555
0 46768 5 1 1 46767
0 46769 7 1 2 90805 46768
0 46770 5 1 1 46769
0 46771 7 1 2 46766 46770
0 46772 5 1 1 46771
0 46773 7 1 2 67736 46772
0 46774 5 1 1 46773
0 46775 7 1 2 68115 46774
0 46776 5 1 1 46775
0 46777 7 1 2 63175 75461
0 46778 5 2 1 46777
0 46779 7 1 2 63555 87552
0 46780 7 1 2 97296 46779
0 46781 7 1 2 46776 46780
0 46782 5 1 1 46781
0 46783 7 1 2 46762 46782
0 46784 7 1 2 46760 46783
0 46785 5 1 1 46784
0 46786 7 1 2 61781 46785
0 46787 5 1 1 46786
0 46788 7 1 2 83012 87553
0 46789 5 1 1 46788
0 46790 7 1 2 83061 74486
0 46791 7 1 2 89060 46790
0 46792 5 1 1 46791
0 46793 7 1 2 46789 46792
0 46794 5 1 1 46793
0 46795 7 1 2 72246 46794
0 46796 5 1 1 46795
0 46797 7 1 2 61782 78272
0 46798 5 1 1 46797
0 46799 7 1 2 46796 46798
0 46800 5 1 1 46799
0 46801 7 1 2 63556 46800
0 46802 5 1 1 46801
0 46803 7 1 2 68503 78481
0 46804 5 1 1 46803
0 46805 7 1 2 73197 95938
0 46806 5 1 1 46805
0 46807 7 1 2 46804 46806
0 46808 5 1 1 46807
0 46809 7 1 2 68116 46808
0 46810 5 1 1 46809
0 46811 7 1 2 68504 93110
0 46812 5 1 1 46811
0 46813 7 1 2 46810 46812
0 46814 5 1 1 46813
0 46815 7 1 2 67374 46814
0 46816 5 1 1 46815
0 46817 7 1 2 80958 95600
0 46818 5 1 1 46817
0 46819 7 1 2 46816 46818
0 46820 5 1 1 46819
0 46821 7 1 2 66750 46820
0 46822 5 1 1 46821
0 46823 7 1 2 46802 46822
0 46824 5 1 1 46823
0 46825 7 1 2 91685 46824
0 46826 5 1 1 46825
0 46827 7 1 2 70658 96489
0 46828 5 1 1 46827
0 46829 7 1 2 89560 46828
0 46830 5 1 1 46829
0 46831 7 1 2 93872 46830
0 46832 5 1 1 46831
0 46833 7 1 2 92137 96261
0 46834 7 1 2 74548 46833
0 46835 5 1 1 46834
0 46836 7 1 2 90176 93869
0 46837 5 1 1 46836
0 46838 7 1 2 68763 46837
0 46839 7 1 2 46835 46838
0 46840 7 1 2 46832 46839
0 46841 7 1 2 46826 46840
0 46842 7 1 2 46787 46841
0 46843 5 1 1 46842
0 46844 7 1 2 78880 89323
0 46845 5 1 1 46844
0 46846 7 1 2 73214 82239
0 46847 5 1 1 46846
0 46848 7 1 2 89792 46847
0 46849 5 1 1 46848
0 46850 7 1 2 76308 46849
0 46851 5 2 1 46850
0 46852 7 2 2 72247 97298
0 46853 5 1 1 97300
0 46854 7 1 2 70659 94175
0 46855 7 1 2 97301 46854
0 46856 5 1 1 46855
0 46857 7 1 2 46845 46856
0 46858 5 1 1 46857
0 46859 7 1 2 68117 46858
0 46860 5 1 1 46859
0 46861 7 1 2 89324 97236
0 46862 5 1 1 46861
0 46863 7 1 2 46860 46862
0 46864 5 1 1 46863
0 46865 7 1 2 68505 46864
0 46866 5 1 1 46865
0 46867 7 1 2 63826 96024
0 46868 7 1 2 46866 46867
0 46869 5 1 1 46868
0 46870 7 1 2 87186 46869
0 46871 7 1 2 46843 46870
0 46872 5 1 1 46871
0 46873 7 1 2 63557 88935
0 46874 5 1 1 46873
0 46875 7 1 2 84657 90927
0 46876 5 1 1 46875
0 46877 7 1 2 46874 46876
0 46878 5 1 1 46877
0 46879 7 1 2 62759 46878
0 46880 5 1 1 46879
0 46881 7 1 2 73050 84790
0 46882 5 1 1 46881
0 46883 7 1 2 77484 90928
0 46884 5 2 1 46883
0 46885 7 2 2 74101 78379
0 46886 5 1 1 97304
0 46887 7 1 2 63558 46886
0 46888 5 1 1 46887
0 46889 7 1 2 97302 46888
0 46890 5 1 1 46889
0 46891 7 1 2 66341 46890
0 46892 5 1 1 46891
0 46893 7 1 2 46882 46892
0 46894 7 1 2 46880 46893
0 46895 5 1 1 46894
0 46896 7 1 2 84198 46895
0 46897 5 1 1 46896
0 46898 7 3 2 78133 78780
0 46899 5 4 1 97306
0 46900 7 1 2 97088 97309
0 46901 5 1 1 46900
0 46902 7 1 2 71835 46901
0 46903 5 1 1 46902
0 46904 7 1 2 69705 97307
0 46905 5 1 1 46904
0 46906 7 1 2 69740 97091
0 46907 5 1 1 46906
0 46908 7 1 2 46905 46907
0 46909 7 1 2 46903 46908
0 46910 5 1 1 46909
0 46911 7 1 2 62760 46910
0 46912 5 1 1 46911
0 46913 7 1 2 92044 97093
0 46914 5 1 1 46913
0 46915 7 1 2 97178 46914
0 46916 7 1 2 46912 46915
0 46917 5 1 1 46916
0 46918 7 1 2 62389 46917
0 46919 5 1 1 46918
0 46920 7 1 2 65504 95214
0 46921 5 1 1 46920
0 46922 7 1 2 97310 46921
0 46923 5 1 1 46922
0 46924 7 1 2 64585 46923
0 46925 5 1 1 46924
0 46926 7 1 2 79185 89706
0 46927 5 1 1 46926
0 46928 7 1 2 46925 46927
0 46929 5 1 1 46928
0 46930 7 1 2 62761 46929
0 46931 5 1 1 46930
0 46932 7 1 2 79021 91196
0 46933 5 2 1 46932
0 46934 7 1 2 46931 97313
0 46935 5 1 1 46934
0 46936 7 1 2 64349 46935
0 46937 5 1 1 46936
0 46938 7 1 2 79159 97174
0 46939 5 1 1 46938
0 46940 7 1 2 77439 78781
0 46941 7 1 2 95176 46940
0 46942 5 1 1 46941
0 46943 7 1 2 46939 46942
0 46944 7 1 2 46937 46943
0 46945 7 1 2 46919 46944
0 46946 5 1 1 46945
0 46947 7 1 2 71274 46946
0 46948 5 1 1 46947
0 46949 7 1 2 46897 46948
0 46950 5 1 1 46949
0 46951 7 1 2 65030 46950
0 46952 5 1 1 46951
0 46953 7 1 2 85828 91161
0 46954 5 1 1 46953
0 46955 7 1 2 74284 78009
0 46956 7 1 2 89707 46955
0 46957 5 1 1 46956
0 46958 7 1 2 46954 46957
0 46959 5 1 1 46958
0 46960 7 1 2 62762 46959
0 46961 5 1 1 46960
0 46962 7 1 2 68506 86552
0 46963 5 1 1 46962
0 46964 7 1 2 79086 46963
0 46965 5 1 1 46964
0 46966 7 1 2 26373 46965
0 46967 5 1 1 46966
0 46968 7 1 2 84199 46967
0 46969 5 1 1 46968
0 46970 7 1 2 46961 46969
0 46971 5 1 1 46970
0 46972 7 1 2 77219 46971
0 46973 5 1 1 46972
0 46974 7 1 2 68507 44501
0 46975 5 1 1 46974
0 46976 7 1 2 69275 46975
0 46977 5 1 1 46976
0 46978 7 1 2 76707 78044
0 46979 5 1 1 46978
0 46980 7 1 2 87974 46979
0 46981 7 1 2 46977 46980
0 46982 5 1 1 46981
0 46983 7 1 2 71461 46982
0 46984 5 1 1 46983
0 46985 7 1 2 68508 24762
0 46986 5 1 1 46985
0 46987 7 1 2 66342 46986
0 46988 5 1 1 46987
0 46989 7 1 2 68509 12977
0 46990 5 1 1 46989
0 46991 7 1 2 94503 46990
0 46992 5 1 1 46991
0 46993 7 1 2 46988 46992
0 46994 7 1 2 46984 46993
0 46995 5 1 1 46994
0 46996 7 1 2 62763 46995
0 46997 5 1 1 46996
0 46998 7 1 2 71315 86852
0 46999 7 1 2 84050 46998
0 47000 5 1 1 46999
0 47001 7 1 2 46997 47000
0 47002 5 1 1 47001
0 47003 7 1 2 63176 47002
0 47004 5 1 1 47003
0 47005 7 1 2 81658 85030
0 47006 5 1 1 47005
0 47007 7 1 2 47004 47006
0 47008 5 1 1 47007
0 47009 7 1 2 84200 47008
0 47010 5 1 1 47009
0 47011 7 1 2 46973 47010
0 47012 7 1 2 46952 47011
0 47013 5 1 1 47012
0 47014 7 1 2 75633 47013
0 47015 5 1 1 47014
0 47016 7 1 2 64586 91438
0 47017 5 2 1 47016
0 47018 7 1 2 68118 97315
0 47019 5 1 1 47018
0 47020 7 1 2 70660 73137
0 47021 5 1 1 47020
0 47022 7 1 2 47019 47021
0 47023 5 1 1 47022
0 47024 7 1 2 93276 47023
0 47025 5 1 1 47024
0 47026 7 1 2 87770 47025
0 47027 5 1 1 47026
0 47028 7 1 2 69276 94129
0 47029 5 1 1 47028
0 47030 7 1 2 84744 47029
0 47031 5 1 1 47030
0 47032 7 1 2 65031 47031
0 47033 5 1 1 47032
0 47034 7 1 2 78041 85822
0 47035 5 1 1 47034
0 47036 7 1 2 63559 47035
0 47037 5 1 1 47036
0 47038 7 1 2 47033 47037
0 47039 5 1 1 47038
0 47040 7 1 2 64587 47039
0 47041 5 1 1 47040
0 47042 7 1 2 68510 86294
0 47043 5 1 1 47042
0 47044 7 1 2 86936 47043
0 47045 5 1 1 47044
0 47046 7 1 2 63560 88573
0 47047 5 1 1 47046
0 47048 7 1 2 47045 47047
0 47049 5 1 1 47048
0 47050 7 1 2 62390 47049
0 47051 5 1 1 47050
0 47052 7 1 2 47041 47051
0 47053 5 1 1 47052
0 47054 7 1 2 70343 47053
0 47055 5 1 1 47054
0 47056 7 1 2 90734 18006
0 47057 5 1 1 47056
0 47058 7 1 2 64588 47057
0 47059 5 1 1 47058
0 47060 7 1 2 84745 47059
0 47061 5 1 1 47060
0 47062 7 1 2 63177 47061
0 47063 5 1 1 47062
0 47064 7 1 2 82309 85011
0 47065 5 1 1 47064
0 47066 7 1 2 47063 47065
0 47067 5 1 1 47066
0 47068 7 1 2 70377 47067
0 47069 5 1 1 47068
0 47070 7 1 2 69375 86292
0 47071 7 1 2 87812 47070
0 47072 5 1 1 47071
0 47073 7 1 2 47069 47072
0 47074 7 1 2 47055 47073
0 47075 7 1 2 47027 47074
0 47076 5 1 1 47075
0 47077 7 1 2 75634 47076
0 47078 5 1 1 47077
0 47079 7 1 2 70661 90922
0 47080 5 1 1 47079
0 47081 7 1 2 63178 47080
0 47082 5 1 1 47081
0 47083 7 1 2 68511 47082
0 47084 5 1 1 47083
0 47085 7 1 2 75238 47084
0 47086 5 1 1 47085
0 47087 7 1 2 47078 47086
0 47088 5 1 1 47087
0 47089 7 1 2 84201 47088
0 47090 5 1 1 47089
0 47091 7 1 2 88394 97175
0 47092 5 1 1 47091
0 47093 7 1 2 80129 76726
0 47094 7 1 2 89708 47093
0 47095 5 1 1 47094
0 47096 7 1 2 47092 47095
0 47097 5 1 1 47096
0 47098 7 1 2 66343 47097
0 47099 5 1 1 47098
0 47100 7 1 2 79989 84216
0 47101 5 1 1 47100
0 47102 7 1 2 47099 47101
0 47103 5 1 1 47102
0 47104 7 1 2 65032 47103
0 47105 5 1 1 47104
0 47106 7 1 2 60179 81954
0 47107 5 1 1 47106
0 47108 7 1 2 84202 47107
0 47109 7 1 2 85386 47108
0 47110 5 1 1 47109
0 47111 7 1 2 80674 85488
0 47112 7 1 2 87980 47111
0 47113 5 1 1 47112
0 47114 7 1 2 47110 47113
0 47115 5 1 1 47114
0 47116 7 1 2 69706 47115
0 47117 5 1 1 47116
0 47118 7 1 2 68119 88668
0 47119 5 1 1 47118
0 47120 7 1 2 84217 47119
0 47121 5 1 1 47120
0 47122 7 1 2 47117 47121
0 47123 7 1 2 47105 47122
0 47124 5 1 1 47123
0 47125 7 1 2 75635 47124
0 47126 5 1 1 47125
0 47127 7 1 2 83561 95348
0 47128 5 1 1 47127
0 47129 7 1 2 97311 47128
0 47130 5 1 1 47129
0 47131 7 1 2 69707 47130
0 47132 5 1 1 47131
0 47133 7 1 2 69861 83562
0 47134 7 1 2 79598 47133
0 47135 5 1 1 47134
0 47136 7 1 2 47132 47135
0 47137 5 1 1 47136
0 47138 7 1 2 74455 47137
0 47139 5 1 1 47138
0 47140 7 1 2 94619 97312
0 47141 5 1 1 47140
0 47142 7 1 2 65033 47141
0 47143 5 1 1 47142
0 47144 7 1 2 15430 47143
0 47145 7 1 2 47139 47144
0 47146 5 1 1 47145
0 47147 7 1 2 91871 47146
0 47148 5 1 1 47147
0 47149 7 1 2 63179 93339
0 47150 5 1 1 47149
0 47151 7 1 2 69140 94271
0 47152 7 1 2 46638 47151
0 47153 7 1 2 89138 47152
0 47154 5 1 1 47153
0 47155 7 1 2 70856 47154
0 47156 5 1 1 47155
0 47157 7 1 2 47150 47156
0 47158 5 1 1 47157
0 47159 7 1 2 97210 47158
0 47160 5 1 1 47159
0 47161 7 1 2 83305 89709
0 47162 5 1 1 47161
0 47163 7 1 2 63561 97168
0 47164 5 1 1 47163
0 47165 7 1 2 47162 47164
0 47166 5 1 1 47165
0 47167 7 1 2 65298 47166
0 47168 5 1 1 47167
0 47169 7 1 2 62391 92596
0 47170 5 1 1 47169
0 47171 7 1 2 93833 47170
0 47172 5 1 1 47171
0 47173 7 1 2 65505 47172
0 47174 5 1 1 47173
0 47175 7 1 2 47168 47174
0 47176 5 1 1 47175
0 47177 7 1 2 60180 95576
0 47178 5 1 1 47177
0 47179 7 1 2 47176 47178
0 47180 5 1 1 47179
0 47181 7 1 2 47160 47180
0 47182 7 1 2 47148 47181
0 47183 7 1 2 47126 47182
0 47184 5 1 1 47183
0 47185 7 1 2 62764 47184
0 47186 5 1 1 47185
0 47187 7 1 2 47090 47186
0 47188 5 1 1 47187
0 47189 7 1 2 72380 47188
0 47190 5 1 1 47189
0 47191 7 1 2 70542 85489
0 47192 5 1 1 47191
0 47193 7 1 2 70429 93148
0 47194 5 1 1 47193
0 47195 7 1 2 62765 47194
0 47196 5 1 1 47195
0 47197 7 1 2 69314 87989
0 47198 5 1 1 47197
0 47199 7 1 2 70458 47198
0 47200 5 1 1 47199
0 47201 7 1 2 33585 47200
0 47202 7 1 2 47196 47201
0 47203 5 1 1 47202
0 47204 7 1 2 71131 83563
0 47205 7 1 2 47203 47204
0 47206 5 1 1 47205
0 47207 7 1 2 47192 47206
0 47208 5 1 1 47207
0 47209 7 1 2 70086 47208
0 47210 5 1 1 47209
0 47211 7 1 2 87464 89692
0 47212 5 1 1 47211
0 47213 7 1 2 85403 47212
0 47214 5 1 1 47213
0 47215 7 1 2 65034 47214
0 47216 5 1 1 47215
0 47217 7 1 2 73745 89710
0 47218 5 2 1 47217
0 47219 7 1 2 47216 97317
0 47220 5 1 1 47219
0 47221 7 1 2 64589 47220
0 47222 5 1 1 47221
0 47223 7 1 2 91102 89693
0 47224 5 1 1 47223
0 47225 7 1 2 47222 47224
0 47226 5 1 1 47225
0 47227 7 1 2 70378 47226
0 47228 5 1 1 47227
0 47229 7 1 2 85404 94620
0 47230 5 1 1 47229
0 47231 7 1 2 65035 47230
0 47232 5 1 1 47231
0 47233 7 1 2 97318 47232
0 47234 5 1 1 47233
0 47235 7 1 2 62392 47234
0 47236 5 1 1 47235
0 47237 7 1 2 82377 86297
0 47238 5 1 1 47237
0 47239 7 1 2 47236 47238
0 47240 5 1 1 47239
0 47241 7 1 2 72602 47240
0 47242 5 1 1 47241
0 47243 7 1 2 71836 74431
0 47244 5 1 1 47243
0 47245 7 1 2 82851 87690
0 47246 5 1 1 47245
0 47247 7 1 2 47244 47246
0 47248 5 1 1 47247
0 47249 7 1 2 70857 85401
0 47250 7 1 2 47248 47249
0 47251 5 1 1 47250
0 47252 7 1 2 91379 95186
0 47253 5 1 1 47252
0 47254 7 1 2 79022 93561
0 47255 7 1 2 47253 47254
0 47256 5 1 1 47255
0 47257 7 1 2 47251 47256
0 47258 7 1 2 47242 47257
0 47259 7 1 2 47228 47258
0 47260 5 1 1 47259
0 47261 7 1 2 72381 47260
0 47262 5 1 1 47261
0 47263 7 1 2 91162 97115
0 47264 5 1 1 47263
0 47265 7 1 2 85405 47264
0 47266 5 1 1 47265
0 47267 7 1 2 77745 47266
0 47268 5 1 1 47267
0 47269 7 1 2 47262 47268
0 47270 7 1 2 47210 47269
0 47271 5 1 1 47270
0 47272 7 1 2 91872 47271
0 47273 5 1 1 47272
0 47274 7 1 2 73215 15511
0 47275 5 1 1 47274
0 47276 7 1 2 74456 90271
0 47277 5 1 1 47276
0 47278 7 1 2 74078 97129
0 47279 5 1 1 47278
0 47280 7 1 2 47277 47279
0 47281 7 1 2 47275 47280
0 47282 5 1 1 47281
0 47283 7 1 2 93716 47282
0 47284 5 1 1 47283
0 47285 7 1 2 78341 89590
0 47286 5 1 1 47285
0 47287 7 1 2 63180 47286
0 47288 5 1 1 47287
0 47289 7 1 2 62393 72787
0 47290 5 1 1 47289
0 47291 7 1 2 93051 47290
0 47292 7 1 2 13879 47291
0 47293 5 1 1 47292
0 47294 7 1 2 62766 93053
0 47295 7 1 2 47293 47294
0 47296 5 1 1 47295
0 47297 7 1 2 47288 47296
0 47298 5 1 1 47297
0 47299 7 1 2 75239 47298
0 47300 5 1 1 47299
0 47301 7 1 2 47284 47300
0 47302 5 1 1 47301
0 47303 7 1 2 84203 47302
0 47304 5 1 1 47303
0 47305 7 1 2 84443 97184
0 47306 7 1 2 97242 47305
0 47307 5 1 1 47306
0 47308 7 1 2 47304 47307
0 47309 5 1 1 47308
0 47310 7 1 2 72506 47309
0 47311 5 1 1 47310
0 47312 7 1 2 70662 97227
0 47313 5 1 1 47312
0 47314 7 1 2 63562 47313
0 47315 5 1 1 47314
0 47316 7 1 2 78273 75088
0 47317 5 1 1 47316
0 47318 7 1 2 90844 47317
0 47319 7 1 2 97303 47318
0 47320 7 1 2 47315 47319
0 47321 5 1 1 47320
0 47322 7 1 2 97211 47321
0 47323 5 1 1 47322
0 47324 7 1 2 47311 47323
0 47325 7 1 2 47273 47324
0 47326 7 1 2 47190 47325
0 47327 7 1 2 47015 47326
0 47328 5 1 1 47327
0 47329 7 1 2 86760 47328
0 47330 5 1 1 47329
0 47331 7 1 2 64350 90221
0 47332 5 1 1 47331
0 47333 7 1 2 78463 47332
0 47334 5 1 1 47333
0 47335 7 2 2 62767 47334
0 47336 5 1 1 97319
0 47337 7 1 2 63181 83368
0 47338 5 1 1 47337
0 47339 7 1 2 47336 47338
0 47340 5 1 1 47339
0 47341 7 1 2 80283 47340
0 47342 5 1 1 47341
0 47343 7 1 2 72025 90318
0 47344 5 1 1 47343
0 47345 7 1 2 87009 47344
0 47346 5 1 1 47345
0 47347 7 1 2 63182 47346
0 47348 5 1 1 47347
0 47349 7 1 2 90390 47348
0 47350 5 1 1 47349
0 47351 7 1 2 70858 47350
0 47352 5 1 1 47351
0 47353 7 1 2 47342 47352
0 47354 5 1 1 47353
0 47355 7 1 2 63563 47354
0 47356 5 1 1 47355
0 47357 7 1 2 68512 44129
0 47358 5 1 1 47357
0 47359 7 1 2 83485 47358
0 47360 5 1 1 47359
0 47361 7 1 2 69708 80284
0 47362 5 1 1 47361
0 47363 7 1 2 91133 47362
0 47364 5 1 1 47363
0 47365 7 1 2 75693 81424
0 47366 7 1 2 47364 47365
0 47367 5 1 1 47366
0 47368 7 1 2 47360 47367
0 47369 5 1 1 47368
0 47370 7 1 2 71837 47369
0 47371 5 1 1 47370
0 47372 7 2 2 76872 85819
0 47373 5 2 1 97321
0 47374 7 1 2 68513 97323
0 47375 5 2 1 47374
0 47376 7 1 2 70859 97325
0 47377 5 1 1 47376
0 47378 7 1 2 65036 94130
0 47379 5 1 1 47378
0 47380 7 1 2 47377 47379
0 47381 5 1 1 47380
0 47382 7 1 2 75636 47381
0 47383 5 1 1 47382
0 47384 7 1 2 86937 91873
0 47385 5 1 1 47384
0 47386 7 1 2 47383 47385
0 47387 5 1 1 47386
0 47388 7 1 2 70410 47387
0 47389 5 1 1 47388
0 47390 7 1 2 77506 97240
0 47391 5 1 1 47390
0 47392 7 1 2 97254 47391
0 47393 5 1 1 47392
0 47394 7 1 2 47389 47393
0 47395 7 1 2 47371 47394
0 47396 7 1 2 47356 47395
0 47397 5 1 1 47396
0 47398 7 1 2 72382 47397
0 47399 5 1 1 47398
0 47400 7 1 2 90405 91850
0 47401 5 4 1 47400
0 47402 7 1 2 90413 97327
0 47403 5 1 1 47402
0 47404 7 1 2 69277 91429
0 47405 5 1 1 47404
0 47406 7 1 2 74232 91385
0 47407 5 1 1 47406
0 47408 7 1 2 47405 47407
0 47409 5 1 1 47408
0 47410 7 1 2 64590 47409
0 47411 5 1 1 47410
0 47412 7 1 2 69161 91430
0 47413 5 1 1 47412
0 47414 7 1 2 47411 47413
0 47415 5 1 1 47414
0 47416 7 1 2 63564 47415
0 47417 5 1 1 47416
0 47418 7 1 2 47403 47417
0 47419 5 1 1 47418
0 47420 7 1 2 63183 47419
0 47421 5 1 1 47420
0 47422 7 1 2 63565 80285
0 47423 5 1 1 47422
0 47424 7 1 2 62394 97255
0 47425 5 1 1 47424
0 47426 7 1 2 47423 47425
0 47427 5 1 1 47426
0 47428 7 1 2 63184 47427
0 47429 5 1 1 47428
0 47430 7 1 2 75637 97326
0 47431 5 1 1 47430
0 47432 7 1 2 26194 47431
0 47433 5 1 1 47432
0 47434 7 1 2 86603 47433
0 47435 5 1 1 47434
0 47436 7 1 2 93786 47435
0 47437 7 1 2 47429 47436
0 47438 5 1 1 47437
0 47439 7 1 2 72383 47438
0 47440 5 1 1 47439
0 47441 7 1 2 80286 71132
0 47442 5 1 1 47441
0 47443 7 1 2 83480 47442
0 47444 5 4 1 47443
0 47445 7 2 2 64351 97331
0 47446 7 2 2 63566 71838
0 47447 7 1 2 72163 97337
0 47448 7 1 2 97335 47447
0 47449 5 1 1 47448
0 47450 7 1 2 47440 47449
0 47451 7 1 2 47421 47450
0 47452 5 1 1 47451
0 47453 7 1 2 70344 47452
0 47454 5 1 1 47453
0 47455 7 1 2 41355 97328
0 47456 5 1 1 47455
0 47457 7 1 2 67737 37230
0 47458 5 1 1 47457
0 47459 7 1 2 63567 91431
0 47460 7 1 2 47458 47459
0 47461 5 1 1 47460
0 47462 7 1 2 47456 47461
0 47463 5 1 1 47462
0 47464 7 1 2 63185 47463
0 47465 5 1 1 47464
0 47466 7 1 2 63568 93070
0 47467 7 1 2 97332 47466
0 47468 5 1 1 47467
0 47469 7 1 2 47465 47468
0 47470 5 1 1 47469
0 47471 7 1 2 69278 47470
0 47472 5 1 1 47471
0 47473 7 1 2 72026 97256
0 47474 5 1 1 47473
0 47475 7 1 2 80287 97338
0 47476 5 1 1 47475
0 47477 7 1 2 47474 47476
0 47478 5 1 1 47477
0 47479 7 1 2 72384 47478
0 47480 5 1 1 47479
0 47481 7 1 2 72507 91874
0 47482 5 1 1 47481
0 47483 7 2 2 18050 47482
0 47484 5 1 1 97339
0 47485 7 1 2 47480 97340
0 47486 5 1 1 47485
0 47487 7 1 2 90974 47486
0 47488 5 1 1 47487
0 47489 7 1 2 69960 75024
0 47490 5 1 1 47489
0 47491 7 1 2 62768 47490
0 47492 5 1 1 47491
0 47493 7 1 2 68120 47492
0 47494 5 1 1 47493
0 47495 7 1 2 75521 78013
0 47496 5 1 1 47495
0 47497 7 1 2 47494 47496
0 47498 5 1 1 47497
0 47499 7 1 2 91376 93490
0 47500 5 1 1 47499
0 47501 7 1 2 70860 91220
0 47502 5 1 1 47501
0 47503 7 1 2 47500 47502
0 47504 7 1 2 47498 47503
0 47505 5 1 1 47504
0 47506 7 1 2 72508 47505
0 47507 5 1 1 47506
0 47508 7 1 2 69146 73386
0 47509 5 1 1 47508
0 47510 7 1 2 63186 47509
0 47511 5 1 1 47510
0 47512 7 1 2 90555 47511
0 47513 5 1 1 47512
0 47514 7 1 2 76435 91432
0 47515 7 1 2 47513 47514
0 47516 5 1 1 47515
0 47517 7 1 2 87249 47516
0 47518 7 1 2 47507 47517
0 47519 5 1 1 47518
0 47520 7 1 2 63569 47519
0 47521 5 1 1 47520
0 47522 7 1 2 65506 96874
0 47523 5 1 1 47522
0 47524 7 1 2 67738 91387
0 47525 5 1 1 47524
0 47526 7 1 2 63187 47525
0 47527 7 1 2 97329 47526
0 47528 5 1 1 47527
0 47529 7 1 2 63570 69075
0 47530 7 1 2 97333 47529
0 47531 5 1 1 47530
0 47532 7 1 2 47528 47531
0 47533 5 1 1 47532
0 47534 7 1 2 82792 47533
0 47535 5 1 1 47534
0 47536 7 1 2 47523 47535
0 47537 7 1 2 47521 47536
0 47538 7 1 2 47488 47537
0 47539 7 1 2 47472 47538
0 47540 7 1 2 47454 47539
0 47541 7 1 2 47399 47540
0 47542 5 1 1 47541
0 47543 7 1 2 86761 47542
0 47544 5 1 1 47543
0 47545 7 1 2 73422 94358
0 47546 7 1 2 95730 47545
0 47547 7 1 2 97299 47546
0 47548 5 1 1 47547
0 47549 7 1 2 63827 47548
0 47550 7 1 2 47544 47549
0 47551 5 1 1 47550
0 47552 7 1 2 60944 71012
0 47553 5 2 1 47552
0 47554 7 1 2 65613 73022
0 47555 5 1 1 47554
0 47556 7 1 2 97341 47555
0 47557 5 1 1 47556
0 47558 7 1 2 96666 47557
0 47559 5 1 1 47558
0 47560 7 1 2 92288 96296
0 47561 7 1 2 47559 47560
0 47562 5 1 1 47561
0 47563 7 1 2 67739 47562
0 47564 5 1 1 47563
0 47565 7 4 2 65614 67375
0 47566 5 2 1 97343
0 47567 7 3 2 68514 97344
0 47568 5 1 1 97349
0 47569 7 1 2 60945 97350
0 47570 5 1 1 47569
0 47571 7 2 2 63188 73359
0 47572 5 1 1 97352
0 47573 7 1 2 75002 97353
0 47574 5 1 1 47573
0 47575 7 1 2 47570 47574
0 47576 7 1 2 47564 47575
0 47577 5 1 1 47576
0 47578 7 1 2 72248 47577
0 47579 5 1 1 47578
0 47580 7 1 2 70663 93873
0 47581 5 1 1 47580
0 47582 7 1 2 83750 97295
0 47583 5 1 1 47582
0 47584 7 1 2 47581 47583
0 47585 5 1 1 47584
0 47586 7 1 2 65615 47585
0 47587 5 1 1 47586
0 47588 7 1 2 47579 47587
0 47589 5 1 1 47588
0 47590 7 1 2 60600 47589
0 47591 5 1 1 47590
0 47592 7 2 2 85330 92820
0 47593 7 1 2 92662 97354
0 47594 5 1 1 47593
0 47595 7 1 2 47591 47594
0 47596 5 1 1 47595
0 47597 7 1 2 75522 47596
0 47598 5 1 1 47597
0 47599 7 5 2 59396 76504
0 47600 7 1 2 89256 92773
0 47601 7 1 2 97356 47600
0 47602 7 1 2 97355 47601
0 47603 5 1 1 47602
0 47604 7 1 2 47598 47603
0 47605 5 1 1 47604
0 47606 7 1 2 66893 47605
0 47607 5 1 1 47606
0 47608 7 1 2 70861 88534
0 47609 5 1 1 47608
0 47610 7 1 2 89187 88406
0 47611 5 1 1 47610
0 47612 7 1 2 70087 47611
0 47613 5 1 1 47612
0 47614 7 1 2 47609 47613
0 47615 5 1 1 47614
0 47616 7 1 2 92045 94373
0 47617 7 1 2 47615 47616
0 47618 5 1 1 47617
0 47619 7 1 2 68764 47618
0 47620 7 1 2 47607 47619
0 47621 5 1 1 47620
0 47622 7 1 2 61783 47621
0 47623 7 1 2 47551 47622
0 47624 5 1 1 47623
0 47625 7 1 2 64118 47624
0 47626 7 1 2 47330 47625
0 47627 7 1 2 46872 47626
0 47628 7 1 2 46707 47627
0 47629 5 1 1 47628
0 47630 7 1 2 95288 47629
0 47631 7 1 2 46291 47630
0 47632 5 1 1 47631
0 47633 7 1 2 44127 47632
0 47634 5 1 1 47633
0 47635 7 1 2 68925 47634
0 47636 5 1 1 47635
0 47637 7 1 2 92134 25497
0 47638 5 1 1 47637
0 47639 7 2 2 59633 47638
0 47640 5 1 1 97361
0 47641 7 1 2 76481 85948
0 47642 5 1 1 47641
0 47643 7 1 2 47640 47642
0 47644 5 2 1 47643
0 47645 7 1 2 66751 97363
0 47646 5 1 1 47645
0 47647 7 1 2 47568 47646
0 47648 5 1 1 47647
0 47649 7 1 2 68926 47648
0 47650 5 1 1 47649
0 47651 7 1 2 60702 92036
0 47652 5 1 1 47651
0 47653 7 1 2 47650 47652
0 47654 5 1 1 47653
0 47655 7 1 2 67104 47654
0 47656 5 1 1 47655
0 47657 7 2 2 67376 95732
0 47658 7 1 2 73485 97365
0 47659 5 1 1 47658
0 47660 7 1 2 47656 47659
0 47661 5 1 1 47660
0 47662 7 1 2 63828 47661
0 47663 5 1 1 47662
0 47664 7 2 2 77928 90104
0 47665 5 1 1 97367
0 47666 7 1 2 85951 47665
0 47667 5 1 1 47666
0 47668 7 1 2 90217 47667
0 47669 5 1 1 47668
0 47670 7 1 2 47663 47669
0 47671 5 1 1 47670
0 47672 7 1 2 61917 47671
0 47673 5 1 1 47672
0 47674 7 6 2 60703 63829
0 47675 7 1 2 63571 88693
0 47676 5 3 1 47675
0 47677 7 2 2 97369 97375
0 47678 7 1 2 67105 97378
0 47679 5 1 1 47678
0 47680 7 1 2 90204 92282
0 47681 7 1 2 69315 47680
0 47682 5 1 1 47681
0 47683 7 1 2 47679 47682
0 47684 5 1 1 47683
0 47685 7 1 2 86183 47684
0 47686 5 1 1 47685
0 47687 7 2 2 77580 89812
0 47688 5 2 1 97380
0 47689 7 1 2 87621 90155
0 47690 7 1 2 97381 47689
0 47691 5 1 1 47690
0 47692 7 1 2 47686 47691
0 47693 5 1 1 47692
0 47694 7 1 2 59634 47693
0 47695 5 1 1 47694
0 47696 7 1 2 85952 92135
0 47697 5 2 1 47696
0 47698 7 4 2 60704 68765
0 47699 7 1 2 78065 97386
0 47700 7 1 2 97384 47699
0 47701 5 1 1 47700
0 47702 7 1 2 47695 47701
0 47703 7 1 2 47673 47702
0 47704 5 1 1 47703
0 47705 7 1 2 60601 47704
0 47706 5 1 1 47705
0 47707 7 1 2 84103 84524
0 47708 5 1 1 47707
0 47709 7 1 2 83564 90105
0 47710 5 1 1 47709
0 47711 7 1 2 47708 47710
0 47712 5 1 1 47711
0 47713 7 1 2 68121 47712
0 47714 5 1 1 47713
0 47715 7 1 2 11406 47714
0 47716 5 1 1 47715
0 47717 7 1 2 92843 47716
0 47718 5 1 1 47717
0 47719 7 1 2 47706 47718
0 47720 5 1 1 47719
0 47721 7 1 2 64119 47720
0 47722 5 1 1 47721
0 47723 7 1 2 76309 89396
0 47724 5 1 1 47723
0 47725 7 1 2 91825 47724
0 47726 5 1 1 47725
0 47727 7 1 2 84104 96606
0 47728 5 1 1 47727
0 47729 7 1 2 47726 47728
0 47730 5 1 1 47729
0 47731 7 3 2 69007 81030
0 47732 7 1 2 86720 97390
0 47733 7 1 2 47730 47732
0 47734 5 1 1 47733
0 47735 7 1 2 47722 47734
0 47736 5 1 1 47735
0 47737 7 1 2 70664 47736
0 47738 5 1 1 47737
0 47739 7 1 2 78289 91762
0 47740 7 2 2 90115 47739
0 47741 7 1 2 61784 73023
0 47742 7 1 2 97393 47741
0 47743 5 1 1 47742
0 47744 7 1 2 84105 96436
0 47745 5 1 1 47744
0 47746 7 1 2 89800 96844
0 47747 5 1 1 47746
0 47748 7 1 2 47745 47747
0 47749 5 1 1 47748
0 47750 7 1 2 68766 47749
0 47751 5 1 1 47750
0 47752 7 1 2 70665 75025
0 47753 7 1 2 97376 47752
0 47754 5 1 1 47753
0 47755 7 1 2 65507 47754
0 47756 5 1 1 47755
0 47757 7 1 2 61785 89783
0 47758 7 1 2 47756 47757
0 47759 5 1 1 47758
0 47760 7 1 2 47751 47759
0 47761 5 1 1 47760
0 47762 7 1 2 68927 47761
0 47763 5 1 1 47762
0 47764 7 1 2 47743 47763
0 47765 5 1 1 47764
0 47766 7 1 2 64120 47765
0 47767 5 1 1 47766
0 47768 7 1 2 75051 93953
0 47769 5 1 1 47768
0 47770 7 1 2 90018 47769
0 47771 5 1 1 47770
0 47772 7 1 2 85682 94606
0 47773 7 1 2 47771 47772
0 47774 5 1 1 47773
0 47775 7 1 2 47767 47774
0 47776 5 1 1 47775
0 47777 7 1 2 87187 47776
0 47778 5 1 1 47777
0 47779 7 19 2 69008 86721
0 47780 7 1 2 96181 97395
0 47781 5 2 1 47780
0 47782 7 2 2 86325 97370
0 47783 7 1 2 64121 69316
0 47784 7 1 2 97416 47783
0 47785 5 1 1 47784
0 47786 7 1 2 97414 47785
0 47787 5 1 1 47786
0 47788 7 1 2 59635 47787
0 47789 5 1 1 47788
0 47790 7 2 2 87631 96911
0 47791 5 1 1 97418
0 47792 7 1 2 47789 47791
0 47793 5 1 1 47792
0 47794 7 1 2 60602 47793
0 47795 5 1 1 47794
0 47796 7 2 2 82233 84364
0 47797 5 1 1 97420
0 47798 7 1 2 67106 97421
0 47799 5 1 1 47798
0 47800 7 1 2 84525 89793
0 47801 5 1 1 47800
0 47802 7 1 2 47799 47801
0 47803 5 1 1 47802
0 47804 7 7 2 60705 68515
0 47805 7 14 2 61918 64122
0 47806 7 1 2 97422 97429
0 47807 7 1 2 47803 47806
0 47808 5 1 1 47807
0 47809 7 1 2 47795 47808
0 47810 5 1 1 47809
0 47811 7 1 2 68122 47810
0 47812 5 1 1 47811
0 47813 7 1 2 84554 84850
0 47814 5 1 1 47813
0 47815 7 1 2 60603 47814
0 47816 5 1 1 47815
0 47817 7 1 2 67740 92387
0 47818 5 1 1 47817
0 47819 7 1 2 47816 47818
0 47820 5 1 1 47819
0 47821 7 1 2 75026 47820
0 47822 5 1 1 47821
0 47823 7 1 2 91771 47822
0 47824 5 1 1 47823
0 47825 7 2 2 69199 97396
0 47826 7 1 2 47824 97443
0 47827 5 1 1 47826
0 47828 7 1 2 47812 47827
0 47829 5 1 1 47828
0 47830 7 1 2 64038 47829
0 47831 5 1 1 47830
0 47832 7 4 2 64123 85537
0 47833 7 1 2 92321 89461
0 47834 7 1 2 97445 47833
0 47835 5 1 1 47834
0 47836 7 1 2 47831 47835
0 47837 7 1 2 47778 47836
0 47838 7 1 2 47738 47837
0 47839 5 1 1 47838
0 47840 7 1 2 95289 47839
0 47841 5 1 1 47840
0 47842 7 3 2 69009 83751
0 47843 7 3 2 92673 97449
0 47844 7 2 2 81259 86283
0 47845 7 2 2 76349 95225
0 47846 7 3 2 59636 60706
0 47847 7 1 2 91763 97459
0 47848 7 1 2 97457 47847
0 47849 7 1 2 97455 47848
0 47850 7 1 2 97452 47849
0 47851 5 1 1 47850
0 47852 7 1 2 47841 47851
0 47853 5 1 1 47852
0 47854 7 1 2 71241 47853
0 47855 5 1 1 47854
0 47856 7 2 2 94823 96730
0 47857 5 1 1 97462
0 47858 7 1 2 83967 95914
0 47859 5 1 1 47858
0 47860 7 1 2 47857 47859
0 47861 5 1 1 47860
0 47862 7 2 2 72249 47861
0 47863 5 1 1 97464
0 47864 7 1 2 94651 96325
0 47865 5 1 1 47864
0 47866 7 1 2 67107 95915
0 47867 5 1 1 47866
0 47868 7 1 2 47865 47867
0 47869 5 1 1 47868
0 47870 7 1 2 83217 47869
0 47871 5 1 1 47870
0 47872 7 1 2 47863 47871
0 47873 5 1 1 47872
0 47874 7 1 2 66894 47873
0 47875 5 1 1 47874
0 47876 7 6 2 64124 70666
0 47877 7 2 2 85538 97466
0 47878 7 1 2 75116 87150
0 47879 7 1 2 97472 47878
0 47880 5 1 1 47879
0 47881 7 1 2 47875 47880
0 47882 5 1 1 47881
0 47883 7 1 2 59637 47882
0 47884 5 1 1 47883
0 47885 7 4 2 65616 61124
0 47886 7 3 2 92215 97474
0 47887 7 2 2 66895 75117
0 47888 7 1 2 96940 97481
0 47889 7 1 2 97478 47888
0 47890 5 1 1 47889
0 47891 7 1 2 47884 47890
0 47892 5 1 1 47891
0 47893 7 1 2 79664 47892
0 47894 5 1 1 47893
0 47895 7 1 2 60707 85683
0 47896 5 2 1 47895
0 47897 7 2 2 94937 97483
0 47898 7 1 2 87633 21416
0 47899 5 3 1 47898
0 47900 7 1 2 96014 97487
0 47901 5 1 1 47900
0 47902 7 1 2 97485 47901
0 47903 5 1 1 47902
0 47904 7 1 2 96109 47903
0 47905 5 1 1 47904
0 47906 7 1 2 20901 94938
0 47907 5 3 1 47906
0 47908 7 1 2 90116 89133
0 47909 7 1 2 97490 47908
0 47910 5 1 1 47909
0 47911 7 1 2 47905 47910
0 47912 5 1 1 47911
0 47913 7 1 2 61919 47912
0 47914 5 1 1 47913
0 47915 7 3 2 83752 77581
0 47916 7 1 2 88914 97493
0 47917 5 1 1 47916
0 47918 7 1 2 40022 47917
0 47919 5 1 1 47918
0 47920 7 1 2 60708 86984
0 47921 7 1 2 47919 47920
0 47922 5 1 1 47921
0 47923 7 1 2 47914 47922
0 47924 5 1 1 47923
0 47925 7 1 2 64125 47924
0 47926 5 1 1 47925
0 47927 7 1 2 84555 92017
0 47928 5 3 1 47927
0 47929 7 1 2 93690 97397
0 47930 7 1 2 97496 47929
0 47931 5 1 1 47930
0 47932 7 1 2 47926 47931
0 47933 7 1 2 47894 47932
0 47934 5 1 1 47933
0 47935 7 1 2 69317 47934
0 47936 5 1 1 47935
0 47937 7 1 2 70862 96362
0 47938 5 1 1 47937
0 47939 7 2 2 87188 87339
0 47940 7 1 2 47938 97499
0 47941 5 1 1 47940
0 47942 7 2 2 67108 70667
0 47943 5 1 1 97501
0 47944 7 1 2 68123 97237
0 47945 5 2 1 47944
0 47946 7 1 2 81625 88881
0 47947 5 1 1 47946
0 47948 7 1 2 97503 47947
0 47949 5 1 1 47948
0 47950 7 1 2 59638 47949
0 47951 5 1 1 47950
0 47952 7 1 2 47943 47951
0 47953 5 1 1 47952
0 47954 7 1 2 92844 47953
0 47955 5 1 1 47954
0 47956 7 1 2 47941 47955
0 47957 5 1 1 47956
0 47958 7 1 2 68516 47957
0 47959 5 1 1 47958
0 47960 7 3 2 83805 72250
0 47961 5 1 1 97505
0 47962 7 1 2 76350 91075
0 47963 5 1 1 47962
0 47964 7 1 2 47961 47963
0 47965 5 1 1 47964
0 47966 7 2 2 70668 47965
0 47967 5 1 1 97508
0 47968 7 1 2 92845 97509
0 47969 5 1 1 47968
0 47970 7 1 2 47959 47969
0 47971 5 1 1 47970
0 47972 7 1 2 79665 47971
0 47973 5 1 1 47972
0 47974 7 1 2 87707 96997
0 47975 5 2 1 47974
0 47976 7 1 2 76351 92255
0 47977 7 1 2 97510 47976
0 47978 5 1 1 47977
0 47979 7 1 2 63830 96320
0 47980 7 1 2 47978 47979
0 47981 7 1 2 47973 47980
0 47982 5 1 1 47981
0 47983 7 1 2 78290 73954
0 47984 7 1 2 74292 47983
0 47985 5 2 1 47984
0 47986 7 1 2 92289 97512
0 47987 5 1 1 47986
0 47988 7 1 2 87095 47987
0 47989 5 1 1 47988
0 47990 7 1 2 79458 97513
0 47991 5 1 1 47990
0 47992 7 1 2 86796 47991
0 47993 5 1 1 47992
0 47994 7 1 2 47989 47993
0 47995 5 1 1 47994
0 47996 7 1 2 72251 47995
0 47997 5 1 1 47996
0 47998 7 1 2 65617 96173
0 47999 5 1 1 47998
0 48000 7 1 2 60709 87076
0 48001 5 1 1 48000
0 48002 7 1 2 47999 48001
0 48003 5 4 1 48002
0 48004 7 1 2 68517 83806
0 48005 7 1 2 97514 48004
0 48006 5 1 1 48005
0 48007 7 1 2 47997 48006
0 48008 5 1 1 48007
0 48009 7 1 2 92256 48008
0 48010 5 1 1 48009
0 48011 7 3 2 63572 72252
0 48012 7 2 2 67109 83807
0 48013 7 1 2 59639 97521
0 48014 5 1 1 48013
0 48015 7 1 2 78274 48014
0 48016 5 1 1 48015
0 48017 7 1 2 97518 48016
0 48018 5 1 1 48017
0 48019 7 2 2 68518 95442
0 48020 7 1 2 69318 97523
0 48021 5 1 1 48020
0 48022 7 1 2 48018 48021
0 48023 5 1 1 48022
0 48024 7 1 2 64039 96531
0 48025 7 1 2 48023 48024
0 48026 5 1 1 48025
0 48027 7 1 2 48010 48026
0 48028 5 1 1 48027
0 48029 7 1 2 70669 48028
0 48030 5 1 1 48029
0 48031 7 1 2 77446 92088
0 48032 5 4 1 48031
0 48033 7 1 2 67110 97525
0 48034 5 1 1 48033
0 48035 7 1 2 78445 48034
0 48036 5 1 1 48035
0 48037 7 1 2 94407 48036
0 48038 5 1 1 48037
0 48039 7 2 2 73024 92046
0 48040 7 1 2 80493 84268
0 48041 7 1 2 97529 48040
0 48042 5 1 1 48041
0 48043 7 1 2 48038 48042
0 48044 5 1 1 48043
0 48045 7 1 2 87189 48044
0 48046 5 1 1 48045
0 48047 7 1 2 92138 92570
0 48048 7 2 2 71426 92351
0 48049 7 1 2 92814 97531
0 48050 7 1 2 48047 48049
0 48051 5 1 1 48050
0 48052 7 1 2 48046 48051
0 48053 5 1 1 48052
0 48054 7 1 2 68928 48053
0 48055 5 1 1 48054
0 48056 7 4 2 59640 79666
0 48057 7 2 2 85882 86215
0 48058 7 1 2 97533 97537
0 48059 5 1 1 48058
0 48060 7 1 2 68767 48059
0 48061 7 1 2 48055 48060
0 48062 7 1 2 48030 48061
0 48063 5 1 1 48062
0 48064 7 1 2 47982 48063
0 48065 5 1 1 48064
0 48066 7 1 2 64126 48065
0 48067 5 1 1 48066
0 48068 7 1 2 76191 90156
0 48069 5 2 1 48068
0 48070 7 1 2 75052 78444
0 48071 5 1 1 48070
0 48072 7 1 2 97539 48071
0 48073 5 1 1 48072
0 48074 7 1 2 94070 48073
0 48075 5 1 1 48074
0 48076 7 1 2 65508 47967
0 48077 5 1 1 48076
0 48078 7 1 2 94067 48077
0 48079 5 1 1 48078
0 48080 7 1 2 48075 48079
0 48081 5 1 1 48080
0 48082 7 1 2 66752 48081
0 48083 5 1 1 48082
0 48084 7 2 2 75118 83062
0 48085 5 1 1 97541
0 48086 7 1 2 81223 97542
0 48087 5 1 1 48086
0 48088 7 1 2 72253 89826
0 48089 5 1 1 48088
0 48090 7 1 2 48087 48089
0 48091 5 1 1 48090
0 48092 7 1 2 60604 48091
0 48093 5 1 1 48092
0 48094 7 1 2 61786 78303
0 48095 7 1 2 89223 48094
0 48096 5 1 1 48095
0 48097 7 1 2 48093 48096
0 48098 5 1 1 48097
0 48099 7 1 2 63831 86722
0 48100 7 1 2 48098 48099
0 48101 5 1 1 48100
0 48102 7 1 2 48083 48101
0 48103 5 1 1 48102
0 48104 7 1 2 64040 48103
0 48105 5 1 1 48104
0 48106 7 1 2 75694 93258
0 48107 5 1 1 48106
0 48108 7 1 2 90567 48107
0 48109 5 1 1 48108
0 48110 7 3 2 66896 87998
0 48111 7 1 2 96091 97543
0 48112 7 1 2 48109 48111
0 48113 5 1 1 48112
0 48114 7 1 2 69010 48113
0 48115 7 1 2 48105 48114
0 48116 5 1 1 48115
0 48117 7 1 2 48067 48116
0 48118 5 1 1 48117
0 48119 7 1 2 47936 48118
0 48120 5 1 1 48119
0 48121 7 1 2 95290 48120
0 48122 5 1 1 48121
0 48123 7 2 2 68929 97025
0 48124 7 3 2 60710 68124
0 48125 7 1 2 65669 74819
0 48126 7 1 2 97548 48125
0 48127 7 1 2 96085 48126
0 48128 7 2 2 97546 48127
0 48129 5 1 1 97551
0 48130 7 1 2 89794 97552
0 48131 5 1 1 48130
0 48132 7 1 2 86392 97465
0 48133 5 1 1 48132
0 48134 7 1 2 94716 97538
0 48135 5 1 1 48134
0 48136 7 1 2 48133 48135
0 48137 5 1 1 48136
0 48138 7 1 2 79667 48137
0 48139 5 1 1 48138
0 48140 7 2 2 63832 97488
0 48141 7 1 2 88882 97553
0 48142 5 1 1 48141
0 48143 7 1 2 66753 92583
0 48144 5 1 1 48143
0 48145 7 1 2 48142 48144
0 48146 5 1 1 48145
0 48147 7 1 2 61920 48146
0 48148 5 1 1 48147
0 48149 7 1 2 94634 97491
0 48150 5 1 1 48149
0 48151 7 1 2 48148 48150
0 48152 5 1 1 48151
0 48153 7 1 2 87761 94754
0 48154 7 1 2 48152 48153
0 48155 5 1 1 48154
0 48156 7 1 2 48139 48155
0 48157 5 1 1 48156
0 48158 7 1 2 95291 48157
0 48159 5 1 1 48158
0 48160 7 2 2 80983 96897
0 48161 7 1 2 95226 96283
0 48162 7 2 2 97555 48161
0 48163 7 2 2 77660 92468
0 48164 7 1 2 87293 92352
0 48165 7 1 2 97559 48164
0 48166 7 1 2 97557 48165
0 48167 5 1 1 48166
0 48168 7 1 2 48159 48167
0 48169 5 1 1 48168
0 48170 7 1 2 76409 48169
0 48171 5 1 1 48170
0 48172 7 1 2 48131 48171
0 48173 7 1 2 48122 48172
0 48174 7 1 2 47855 48173
0 48175 5 1 1 48174
0 48176 7 1 2 75353 48175
0 48177 5 1 1 48176
0 48178 7 1 2 91983 97351
0 48179 5 1 1 48178
0 48180 7 1 2 84748 90126
0 48181 5 1 1 48180
0 48182 7 1 2 48179 48181
0 48183 5 1 1 48182
0 48184 7 1 2 67111 48183
0 48185 5 1 1 48184
0 48186 7 1 2 80632 92122
0 48187 5 1 1 48186
0 48188 7 1 2 48185 48187
0 48189 5 1 1 48188
0 48190 7 1 2 61787 48189
0 48191 5 1 1 48190
0 48192 7 2 2 67112 79444
0 48193 5 1 1 97561
0 48194 7 1 2 81260 92123
0 48195 7 1 2 97562 48194
0 48196 5 1 1 48195
0 48197 7 1 2 48191 48196
0 48198 5 1 1 48197
0 48199 7 1 2 95871 48198
0 48200 5 1 1 48199
0 48201 7 3 2 75523 92774
0 48202 5 2 1 97563
0 48203 7 1 2 81998 97564
0 48204 5 1 1 48203
0 48205 7 1 2 48200 48204
0 48206 5 1 1 48205
0 48207 7 1 2 66897 48206
0 48208 5 1 1 48207
0 48209 7 1 2 91416 96496
0 48210 5 3 1 48209
0 48211 7 2 2 68519 97568
0 48212 5 3 1 97571
0 48213 7 1 2 80823 96845
0 48214 5 1 1 48213
0 48215 7 1 2 63573 74293
0 48216 7 1 2 94176 48215
0 48217 5 1 1 48216
0 48218 7 1 2 48214 48217
0 48219 5 1 1 48218
0 48220 7 1 2 95872 48219
0 48221 5 1 1 48220
0 48222 7 1 2 97573 48221
0 48223 5 1 1 48222
0 48224 7 1 2 86797 48223
0 48225 5 1 1 48224
0 48226 7 1 2 48208 48225
0 48227 5 1 1 48226
0 48228 7 1 2 68930 48227
0 48229 5 1 1 48228
0 48230 7 1 2 75524 96532
0 48231 5 1 1 48230
0 48232 7 1 2 96538 48231
0 48233 5 5 1 48232
0 48234 7 1 2 76564 69200
0 48235 7 1 2 79732 48234
0 48236 7 1 2 97576 48235
0 48237 5 1 1 48236
0 48238 7 1 2 48229 48237
0 48239 5 1 1 48238
0 48240 7 1 2 68768 48239
0 48241 5 1 1 48240
0 48242 7 1 2 59967 81626
0 48243 5 1 1 48242
0 48244 7 1 2 63189 48243
0 48245 5 2 1 48244
0 48246 7 1 2 86302 87865
0 48247 7 1 2 97581 48246
0 48248 7 1 2 97577 48247
0 48249 5 1 1 48248
0 48250 7 1 2 48241 48249
0 48251 5 1 1 48250
0 48252 7 1 2 64127 48251
0 48253 5 1 1 48252
0 48254 7 6 2 69011 87999
0 48255 7 2 2 93632 97583
0 48256 7 1 2 96876 97582
0 48257 5 1 1 48256
0 48258 7 1 2 80824 96768
0 48259 5 1 1 48258
0 48260 7 1 2 48257 48259
0 48261 5 1 1 48260
0 48262 7 1 2 97589 48261
0 48263 5 1 1 48262
0 48264 7 1 2 48253 48263
0 48265 5 1 1 48264
0 48266 7 1 2 59641 48265
0 48267 5 1 1 48266
0 48268 7 1 2 83249 89711
0 48269 5 1 1 48268
0 48270 7 2 2 75443 79023
0 48271 5 2 1 97591
0 48272 7 1 2 48269 97593
0 48273 5 1 1 48272
0 48274 7 3 2 70670 94755
0 48275 7 2 2 48273 97595
0 48276 7 1 2 86824 97566
0 48277 5 4 1 48276
0 48278 7 1 2 97598 97600
0 48279 5 1 1 48278
0 48280 7 1 2 77119 84011
0 48281 7 1 2 79489 48280
0 48282 5 1 1 48281
0 48283 7 1 2 91401 48282
0 48284 5 1 1 48283
0 48285 7 1 2 86476 97398
0 48286 7 1 2 48284 48285
0 48287 5 1 1 48286
0 48288 7 1 2 48279 48287
0 48289 5 1 1 48288
0 48290 7 1 2 61788 48289
0 48291 5 1 1 48290
0 48292 7 1 2 78147 91540
0 48293 5 1 1 48292
0 48294 7 2 2 64041 48293
0 48295 7 2 2 79721 92360
0 48296 5 1 1 97606
0 48297 7 2 2 64128 97607
0 48298 5 1 1 97608
0 48299 7 1 2 97604 97609
0 48300 5 1 1 48299
0 48301 7 3 2 61789 79722
0 48302 7 2 2 95742 97610
0 48303 5 2 1 97613
0 48304 7 2 2 89940 97399
0 48305 7 1 2 66754 97617
0 48306 5 2 1 48305
0 48307 7 1 2 97615 97619
0 48308 5 2 1 48307
0 48309 7 1 2 97605 97621
0 48310 5 1 1 48309
0 48311 7 1 2 86798 97599
0 48312 5 1 1 48311
0 48313 7 1 2 48310 48312
0 48314 5 1 1 48313
0 48315 7 1 2 91686 48314
0 48316 5 1 1 48315
0 48317 7 1 2 48300 48316
0 48318 7 1 2 48291 48317
0 48319 7 1 2 48267 48318
0 48320 5 1 1 48319
0 48321 7 1 2 95292 48320
0 48322 5 1 1 48321
0 48323 7 2 2 85623 97590
0 48324 5 2 1 97623
0 48325 7 1 2 85859 87134
0 48326 5 3 1 48325
0 48327 7 1 2 89224 97627
0 48328 5 1 1 48327
0 48329 7 1 2 81110 86738
0 48330 5 1 1 48329
0 48331 7 1 2 48328 48330
0 48332 5 1 1 48331
0 48333 7 1 2 96948 48332
0 48334 5 1 1 48333
0 48335 7 3 2 83108 96846
0 48336 5 1 1 97630
0 48337 7 3 2 65618 75119
0 48338 5 2 1 97633
0 48339 7 1 2 48336 97636
0 48340 5 1 1 48339
0 48341 7 1 2 96912 48340
0 48342 5 1 1 48341
0 48343 7 1 2 48334 48342
0 48344 5 1 1 48343
0 48345 7 1 2 60605 48344
0 48346 5 1 1 48345
0 48347 7 3 2 97430 97549
0 48348 5 1 1 97638
0 48349 7 1 2 83565 97639
0 48350 5 3 1 48349
0 48351 7 5 2 85015 86519
0 48352 7 1 2 97419 97644
0 48353 5 1 1 48352
0 48354 7 1 2 97641 48353
0 48355 7 1 2 48346 48354
0 48356 5 1 1 48355
0 48357 7 1 2 75525 48356
0 48358 5 1 1 48357
0 48359 7 2 2 91687 96904
0 48360 7 1 2 92470 97649
0 48361 5 1 1 48360
0 48362 7 6 2 69012 92273
0 48363 7 2 2 83109 97651
0 48364 5 1 1 97657
0 48365 7 1 2 48361 48364
0 48366 5 1 1 48365
0 48367 7 1 2 70671 48366
0 48368 5 1 1 48367
0 48369 7 6 2 66755 94213
0 48370 7 3 2 77800 86666
0 48371 5 1 1 97665
0 48372 7 1 2 97659 97666
0 48373 5 1 1 48372
0 48374 7 1 2 48368 48373
0 48375 5 1 1 48374
0 48376 7 1 2 86799 48375
0 48377 5 1 1 48376
0 48378 7 5 2 92775 96916
0 48379 7 3 2 84526 97668
0 48380 5 2 1 97673
0 48381 7 4 2 60711 85850
0 48382 5 1 1 97678
0 48383 7 3 2 96669 97679
0 48384 7 1 2 67113 97682
0 48385 5 1 1 48384
0 48386 7 1 2 97676 48385
0 48387 5 1 1 48386
0 48388 7 1 2 70672 48387
0 48389 5 1 1 48388
0 48390 7 1 2 87622 96955
0 48391 5 1 1 48390
0 48392 7 2 2 86977 94214
0 48393 7 1 2 97685 97634
0 48394 5 1 1 48393
0 48395 7 1 2 97642 48394
0 48396 5 1 1 48395
0 48397 7 1 2 60606 48396
0 48398 5 1 1 48397
0 48399 7 1 2 48391 48398
0 48400 7 1 2 48389 48399
0 48401 7 1 2 48377 48400
0 48402 7 1 2 48358 48401
0 48403 5 1 1 48402
0 48404 7 1 2 64042 48403
0 48405 5 1 1 48404
0 48406 7 1 2 97625 48405
0 48407 5 1 1 48406
0 48408 7 1 2 95293 48407
0 48409 5 1 1 48408
0 48410 7 3 2 90072 95259
0 48411 7 2 2 90205 97687
0 48412 7 1 2 86143 87294
0 48413 7 1 2 95236 48412
0 48414 7 1 2 97690 48413
0 48415 5 1 1 48414
0 48416 7 1 2 48409 48415
0 48417 5 1 1 48416
0 48418 7 1 2 77008 48417
0 48419 5 1 1 48418
0 48420 7 1 2 96231 97006
0 48421 5 1 1 48420
0 48422 7 1 2 94177 96518
0 48423 7 1 2 97463 48422
0 48424 5 1 1 48423
0 48425 7 1 2 48421 48424
0 48426 5 3 1 48425
0 48427 7 1 2 95294 97692
0 48428 5 1 1 48427
0 48429 7 3 2 95252 97556
0 48430 7 3 2 68125 97695
0 48431 7 3 2 89657 95260
0 48432 7 2 2 97698 97701
0 48433 5 1 1 97704
0 48434 7 1 2 48428 48433
0 48435 5 1 1 48434
0 48436 7 1 2 78464 95765
0 48437 7 1 2 48435 48436
0 48438 5 1 1 48437
0 48439 7 1 2 48419 48438
0 48440 7 1 2 48322 48439
0 48441 5 1 1 48440
0 48442 7 1 2 67741 48441
0 48443 5 1 1 48442
0 48444 7 2 2 60181 94986
0 48445 7 1 2 97706 97686
0 48446 5 1 1 48445
0 48447 7 1 2 48446 97643
0 48448 5 2 1 48447
0 48449 7 1 2 60607 97708
0 48450 5 1 1 48449
0 48451 7 1 2 60712 96956
0 48452 5 1 1 48451
0 48453 7 1 2 79382 96847
0 48454 7 1 2 95696 48453
0 48455 5 1 1 48454
0 48456 7 1 2 48452 48455
0 48457 5 1 1 48456
0 48458 7 1 2 63574 48457
0 48459 5 1 1 48458
0 48460 7 1 2 48450 48459
0 48461 5 1 1 48460
0 48462 7 1 2 64043 48461
0 48463 5 1 1 48462
0 48464 7 1 2 97626 48463
0 48465 5 1 1 48464
0 48466 7 1 2 77009 48465
0 48467 5 1 1 48466
0 48468 7 1 2 92157 96585
0 48469 5 1 1 48468
0 48470 7 1 2 70673 96446
0 48471 5 2 1 48470
0 48472 7 1 2 89561 97710
0 48473 5 1 1 48472
0 48474 7 4 2 68769 96326
0 48475 7 1 2 94254 97712
0 48476 7 1 2 48473 48475
0 48477 5 1 1 48476
0 48478 7 1 2 48469 48477
0 48479 5 1 1 48478
0 48480 7 1 2 65619 48479
0 48481 5 1 1 48480
0 48482 7 1 2 87101 10968
0 48483 5 1 1 48482
0 48484 7 2 2 97423 97446
0 48485 7 1 2 96174 97716
0 48486 7 1 2 48483 48485
0 48487 5 1 1 48486
0 48488 7 1 2 48481 48487
0 48489 7 1 2 48467 48488
0 48490 5 1 1 48489
0 48491 7 1 2 59642 48490
0 48492 5 1 1 48491
0 48493 7 1 2 97473 97511
0 48494 5 1 1 48493
0 48495 7 2 2 87994 92313
0 48496 7 1 2 69201 83784
0 48497 5 2 1 48496
0 48498 7 1 2 83044 97720
0 48499 5 1 1 48498
0 48500 7 1 2 97718 48499
0 48501 5 1 1 48500
0 48502 7 1 2 92178 94103
0 48503 5 1 1 48502
0 48504 7 1 2 86990 48503
0 48505 5 1 1 48504
0 48506 7 1 2 65620 96787
0 48507 7 1 2 48505 48506
0 48508 5 1 1 48507
0 48509 7 1 2 48501 48508
0 48510 5 1 1 48509
0 48511 7 1 2 96327 48510
0 48512 5 1 1 48511
0 48513 7 1 2 85851 95916
0 48514 7 1 2 89728 48513
0 48515 5 1 1 48514
0 48516 7 1 2 48512 48515
0 48517 5 1 1 48516
0 48518 7 1 2 63833 48517
0 48519 5 1 1 48518
0 48520 7 1 2 87708 48382
0 48521 5 3 1 48520
0 48522 7 4 2 64129 77582
0 48523 7 1 2 83433 89013
0 48524 7 1 2 97725 48523
0 48525 7 1 2 97722 48524
0 48526 5 1 1 48525
0 48527 7 1 2 48519 48526
0 48528 5 1 1 48527
0 48529 7 1 2 68520 48528
0 48530 5 1 1 48529
0 48531 7 1 2 48494 48530
0 48532 7 1 2 48492 48531
0 48533 5 1 1 48532
0 48534 7 1 2 95295 48533
0 48535 5 1 1 48534
0 48536 7 1 2 95917 95969
0 48537 5 1 1 48536
0 48538 7 1 2 96793 97631
0 48539 5 1 1 48538
0 48540 7 1 2 92283 96788
0 48541 5 1 1 48540
0 48542 7 1 2 48539 48541
0 48543 5 1 1 48542
0 48544 7 1 2 96328 48543
0 48545 5 1 1 48544
0 48546 7 1 2 48537 48545
0 48547 5 1 1 48546
0 48548 7 1 2 63834 48547
0 48549 5 1 1 48548
0 48550 7 1 2 83384 83753
0 48551 7 2 2 60713 71652
0 48552 7 1 2 97726 97729
0 48553 7 1 2 48550 48552
0 48554 5 1 1 48553
0 48555 7 1 2 48549 48554
0 48556 5 1 1 48555
0 48557 7 1 2 66898 48556
0 48558 5 1 1 48557
0 48559 7 1 2 63575 78066
0 48560 7 6 2 68126 64130
0 48561 7 1 2 97387 97731
0 48562 7 1 2 48559 48561
0 48563 7 1 2 96794 48562
0 48564 5 1 1 48563
0 48565 7 1 2 48558 48564
0 48566 5 1 1 48565
0 48567 7 1 2 60608 48566
0 48568 5 1 1 48567
0 48569 7 8 2 64131 87190
0 48570 7 3 2 68931 97737
0 48571 7 1 2 95972 97745
0 48572 5 1 1 48571
0 48573 7 1 2 77010 97709
0 48574 5 1 1 48573
0 48575 7 3 2 87077 96731
0 48576 7 2 2 82462 87893
0 48577 7 1 2 97748 97751
0 48578 5 1 1 48577
0 48579 7 1 2 48574 48578
0 48580 5 1 1 48579
0 48581 7 1 2 59643 48580
0 48582 5 1 1 48581
0 48583 7 1 2 97738 97752
0 48584 5 1 1 48583
0 48585 7 3 2 86573 96732
0 48586 5 1 1 97753
0 48587 7 1 2 48584 48586
0 48588 5 1 1 48587
0 48589 7 1 2 83250 48588
0 48590 5 1 1 48589
0 48591 7 4 2 69013 84444
0 48592 7 2 2 86723 97756
0 48593 5 1 1 97760
0 48594 7 1 2 48590 48593
0 48595 5 1 1 48594
0 48596 7 1 2 81999 48595
0 48597 5 1 1 48596
0 48598 7 1 2 48582 48597
0 48599 5 1 1 48598
0 48600 7 1 2 64044 48599
0 48601 5 1 1 48600
0 48602 7 1 2 48572 48601
0 48603 7 1 2 48568 48602
0 48604 5 1 1 48603
0 48605 7 1 2 95296 48604
0 48606 5 1 1 48605
0 48607 7 1 2 66756 95144
0 48608 7 1 2 97011 48607
0 48609 5 1 1 48608
0 48610 7 1 2 63576 89005
0 48611 5 1 1 48610
0 48612 7 1 2 61790 97388
0 48613 7 1 2 95230 48612
0 48614 7 1 2 48611 48613
0 48615 5 1 1 48614
0 48616 7 1 2 48609 48615
0 48617 5 1 1 48616
0 48618 7 1 2 70674 48617
0 48619 5 1 1 48618
0 48620 7 1 2 88118 89069
0 48621 5 1 1 48620
0 48622 7 1 2 97347 48621
0 48623 5 1 1 48622
0 48624 7 1 2 95705 97012
0 48625 7 1 2 48623 48624
0 48626 5 1 1 48625
0 48627 7 1 2 48619 48626
0 48628 5 1 1 48627
0 48629 7 1 2 68932 48628
0 48630 5 1 1 48629
0 48631 7 1 2 82729 85612
0 48632 5 1 1 48631
0 48633 7 1 2 81111 96795
0 48634 5 1 1 48633
0 48635 7 1 2 48632 48634
0 48636 5 1 1 48635
0 48637 7 10 2 64045 95297
0 48638 7 1 2 96949 97762
0 48639 7 1 2 48636 48638
0 48640 5 1 1 48639
0 48641 7 1 2 48630 48640
0 48642 5 1 1 48641
0 48643 7 1 2 96244 48642
0 48644 5 1 1 48643
0 48645 7 1 2 48606 48644
0 48646 5 1 1 48645
0 48647 7 1 2 61608 48646
0 48648 5 1 1 48647
0 48649 7 1 2 81121 83063
0 48650 7 6 2 86724 95298
0 48651 7 1 2 97713 97772
0 48652 7 1 2 48649 48651
0 48653 5 1 1 48652
0 48654 7 1 2 48648 48653
0 48655 5 1 1 48654
0 48656 7 1 2 60403 48655
0 48657 5 1 1 48656
0 48658 7 1 2 48535 48657
0 48659 5 1 1 48658
0 48660 7 1 2 67114 48659
0 48661 5 1 1 48660
0 48662 7 2 2 97547 97688
0 48663 5 1 1 97778
0 48664 7 1 2 67377 97779
0 48665 5 1 1 48664
0 48666 7 1 2 84888 86184
0 48667 5 1 1 48666
0 48668 7 1 2 89566 93932
0 48669 5 1 1 48668
0 48670 7 1 2 48667 48669
0 48671 5 1 1 48670
0 48672 7 1 2 65509 48671
0 48673 5 1 1 48672
0 48674 7 2 2 89521 93933
0 48675 5 1 1 97780
0 48676 7 1 2 86859 97781
0 48677 5 1 1 48676
0 48678 7 1 2 48673 48677
0 48679 5 1 1 48678
0 48680 7 1 2 66757 48679
0 48681 5 1 1 48680
0 48682 7 1 2 76889 85016
0 48683 7 1 2 96988 48682
0 48684 5 1 1 48683
0 48685 7 1 2 90127 96938
0 48686 5 1 1 48685
0 48687 7 1 2 48684 48686
0 48688 5 1 1 48687
0 48689 7 1 2 84445 94880
0 48690 7 1 2 48688 48689
0 48691 5 1 1 48690
0 48692 7 1 2 48681 48691
0 48693 5 1 1 48692
0 48694 7 1 2 69014 48693
0 48695 5 1 1 48694
0 48696 7 1 2 92226 94756
0 48697 7 1 2 97456 48696
0 48698 5 1 1 48697
0 48699 7 1 2 48695 48698
0 48700 5 1 1 48699
0 48701 7 1 2 65621 48700
0 48702 5 1 1 48701
0 48703 7 2 2 81261 93633
0 48704 5 1 1 97782
0 48705 7 1 2 61791 97783
0 48706 5 1 1 48705
0 48707 7 3 2 63190 86259
0 48708 7 1 2 86477 97784
0 48709 5 1 1 48708
0 48710 7 1 2 48706 48709
0 48711 5 1 1 48710
0 48712 7 1 2 91688 48711
0 48713 5 1 1 48712
0 48714 7 1 2 82000 87938
0 48715 5 1 1 48714
0 48716 7 1 2 48704 48715
0 48717 5 1 1 48716
0 48718 7 1 2 90177 48717
0 48719 5 1 1 48718
0 48720 7 1 2 48713 48719
0 48721 5 1 1 48720
0 48722 7 1 2 64132 48721
0 48723 5 1 1 48722
0 48724 7 1 2 67378 87078
0 48725 7 1 2 85624 48724
0 48726 7 1 2 94607 48725
0 48727 5 1 1 48726
0 48728 7 1 2 48723 48727
0 48729 5 1 1 48728
0 48730 7 1 2 60714 48729
0 48731 5 1 1 48730
0 48732 7 5 2 63835 70675
0 48733 7 1 2 92067 96796
0 48734 5 1 1 48733
0 48735 7 1 2 67379 80551
0 48736 5 1 1 48735
0 48737 7 1 2 48734 48736
0 48738 5 1 1 48737
0 48739 7 1 2 97787 48738
0 48740 5 1 1 48739
0 48741 7 1 2 78067 87738
0 48742 5 1 1 48741
0 48743 7 1 2 48740 48742
0 48744 5 1 1 48743
0 48745 7 1 2 97431 48744
0 48746 5 1 1 48745
0 48747 7 3 2 77929 96329
0 48748 7 1 2 86527 97788
0 48749 7 1 2 97792 48748
0 48750 5 1 1 48749
0 48751 7 1 2 48746 48750
0 48752 7 1 2 48731 48751
0 48753 5 1 1 48752
0 48754 7 1 2 65622 92131
0 48755 5 12 1 48754
0 48756 7 1 2 48753 97795
0 48757 5 1 1 48756
0 48758 7 2 2 96877 97757
0 48759 7 2 2 97544 97807
0 48760 5 1 1 97809
0 48761 7 1 2 68933 97810
0 48762 5 1 1 48761
0 48763 7 1 2 86800 97569
0 48764 5 1 1 48763
0 48765 7 1 2 87225 48764
0 48766 5 2 1 48765
0 48767 7 1 2 92674 97811
0 48768 5 1 1 48767
0 48769 7 1 2 66899 80908
0 48770 5 4 1 48769
0 48771 7 1 2 75526 97813
0 48772 5 2 1 48771
0 48773 7 1 2 40597 97817
0 48774 5 2 1 48773
0 48775 7 2 2 87866 97550
0 48776 7 1 2 70676 97821
0 48777 7 1 2 97819 48776
0 48778 5 1 1 48777
0 48779 7 1 2 48768 48778
0 48780 5 1 1 48779
0 48781 7 1 2 95706 48780
0 48782 5 1 1 48781
0 48783 7 1 2 48762 48782
0 48784 5 1 1 48783
0 48785 7 1 2 96797 48784
0 48786 5 1 1 48785
0 48787 7 1 2 48757 48786
0 48788 7 1 2 48702 48787
0 48789 5 1 1 48788
0 48790 7 1 2 95299 48789
0 48791 5 1 1 48790
0 48792 7 1 2 48665 48791
0 48793 7 1 2 48661 48792
0 48794 7 1 2 48443 48793
0 48795 5 1 1 48794
0 48796 7 1 2 61125 48795
0 48797 5 1 1 48796
0 48798 7 1 2 84218 38147
0 48799 5 1 1 48798
0 48800 7 1 2 92439 89070
0 48801 5 1 1 48800
0 48802 7 1 2 81458 84603
0 48803 5 3 1 48802
0 48804 7 1 2 66583 97823
0 48805 5 1 1 48804
0 48806 7 1 2 59644 48805
0 48807 5 1 1 48806
0 48808 7 1 2 82274 78380
0 48809 5 1 1 48808
0 48810 7 1 2 66584 48809
0 48811 5 1 1 48810
0 48812 7 1 2 60946 48811
0 48813 5 1 1 48812
0 48814 7 1 2 5263 48813
0 48815 7 1 2 48807 48814
0 48816 5 1 1 48815
0 48817 7 1 2 65510 48816
0 48818 5 1 1 48817
0 48819 7 1 2 48801 48818
0 48820 5 1 1 48819
0 48821 7 1 2 68521 48820
0 48822 5 1 1 48821
0 48823 7 1 2 90166 96067
0 48824 5 1 1 48823
0 48825 7 1 2 86563 90614
0 48826 5 1 1 48825
0 48827 7 1 2 48824 48826
0 48828 7 1 2 48822 48827
0 48829 5 1 1 48828
0 48830 7 1 2 63836 48829
0 48831 5 1 1 48830
0 48832 7 1 2 48799 48831
0 48833 5 1 1 48832
0 48834 7 1 2 96917 48833
0 48835 5 1 1 48834
0 48836 7 2 2 68127 76410
0 48837 5 2 1 97826
0 48838 7 1 2 89830 97828
0 48839 5 1 1 48838
0 48840 7 3 2 64133 96245
0 48841 7 1 2 89941 97830
0 48842 7 1 2 48839 48841
0 48843 5 1 1 48842
0 48844 7 1 2 48835 48843
0 48845 5 1 1 48844
0 48846 7 1 2 66758 48845
0 48847 5 1 1 48846
0 48848 7 1 2 40629 97721
0 48849 5 2 1 48848
0 48850 7 2 2 63577 97833
0 48851 7 1 2 95828 97835
0 48852 5 1 1 48851
0 48853 7 1 2 59645 45414
0 48854 5 1 1 48853
0 48855 7 1 2 97829 48854
0 48856 5 1 1 48855
0 48857 7 1 2 68522 79267
0 48858 7 1 2 87369 48857
0 48859 7 1 2 48856 48858
0 48860 5 1 1 48859
0 48861 7 1 2 48852 48860
0 48862 5 1 1 48861
0 48863 7 1 2 68770 48862
0 48864 5 1 1 48863
0 48865 7 1 2 79863 81226
0 48866 5 1 1 48865
0 48867 7 1 2 59646 48866
0 48868 5 1 1 48867
0 48869 7 1 2 82594 48868
0 48870 5 1 1 48869
0 48871 7 1 2 67115 48870
0 48872 5 1 1 48871
0 48873 7 1 2 83760 23452
0 48874 7 1 2 48872 48873
0 48875 5 1 1 48874
0 48876 7 1 2 83154 48875
0 48877 5 1 1 48876
0 48878 7 1 2 48864 48877
0 48879 5 1 1 48878
0 48880 7 1 2 97432 48879
0 48881 5 1 1 48880
0 48882 7 2 2 91183 94215
0 48883 7 1 2 80790 86978
0 48884 7 1 2 97837 48883
0 48885 5 1 1 48884
0 48886 7 1 2 48881 48885
0 48887 7 1 2 48847 48886
0 48888 5 1 1 48887
0 48889 7 1 2 65623 48888
0 48890 5 1 1 48889
0 48891 7 1 2 59647 81711
0 48892 5 1 1 48891
0 48893 7 1 2 5909 48892
0 48894 5 1 1 48893
0 48895 7 1 2 92335 48894
0 48896 5 1 1 48895
0 48897 7 1 2 76581 79723
0 48898 5 1 1 48897
0 48899 7 1 2 48896 48898
0 48900 5 1 1 48899
0 48901 7 1 2 65624 48900
0 48902 5 1 1 48901
0 48903 7 2 2 61921 76565
0 48904 7 2 2 93916 97839
0 48905 5 1 1 97841
0 48906 7 1 2 66759 97842
0 48907 5 1 1 48906
0 48908 7 1 2 94255 96508
0 48909 5 1 1 48908
0 48910 7 1 2 48907 48909
0 48911 5 1 1 48910
0 48912 7 1 2 72136 48911
0 48913 5 1 1 48912
0 48914 7 5 2 60715 67116
0 48915 7 1 2 83937 93981
0 48916 7 1 2 97843 48915
0 48917 5 1 1 48916
0 48918 7 1 2 48913 48917
0 48919 7 1 2 48902 48918
0 48920 5 1 1 48919
0 48921 7 1 2 60609 48920
0 48922 5 1 1 48921
0 48923 7 2 2 67117 91826
0 48924 5 2 1 97848
0 48925 7 1 2 96053 97850
0 48926 5 1 1 48925
0 48927 7 1 2 69319 48926
0 48928 5 1 1 48927
0 48929 7 1 2 83938 89813
0 48930 5 1 1 48929
0 48931 7 1 2 47797 48930
0 48932 7 1 2 48928 48931
0 48933 5 1 1 48932
0 48934 7 1 2 59648 48933
0 48935 5 1 1 48934
0 48936 7 1 2 68771 91908
0 48937 5 1 1 48936
0 48938 7 1 2 72137 84365
0 48939 5 1 1 48938
0 48940 7 1 2 91836 48939
0 48941 7 1 2 48937 48940
0 48942 5 1 1 48941
0 48943 7 1 2 68128 48942
0 48944 5 1 1 48943
0 48945 7 1 2 48935 48944
0 48946 5 1 1 48945
0 48947 7 1 2 86801 48946
0 48948 5 1 1 48947
0 48949 7 1 2 48922 48948
0 48950 5 1 1 48949
0 48951 7 1 2 61609 64134
0 48952 7 1 2 48950 48951
0 48953 5 1 1 48952
0 48954 7 3 2 63191 94216
0 48955 7 1 2 88003 89071
0 48956 7 1 2 97852 48955
0 48957 5 1 1 48956
0 48958 7 1 2 48953 48957
0 48959 5 1 1 48958
0 48960 7 1 2 68523 48959
0 48961 5 1 1 48960
0 48962 7 5 2 63578 69015
0 48963 7 2 2 77485 97855
0 48964 7 1 2 67118 97545
0 48965 7 2 2 97860 48964
0 48966 5 1 1 97862
0 48967 7 1 2 76373 69290
0 48968 5 1 1 48967
0 48969 7 1 2 59649 48968
0 48970 5 1 1 48969
0 48971 7 1 2 84123 48970
0 48972 5 1 1 48971
0 48973 7 1 2 33708 44100
0 48974 5 1 1 48973
0 48975 7 1 2 97467 48974
0 48976 7 1 2 48972 48975
0 48977 5 1 1 48976
0 48978 7 1 2 48966 48977
0 48979 5 1 1 48978
0 48980 7 1 2 61610 48979
0 48981 5 1 1 48980
0 48982 7 1 2 59968 88703
0 48983 5 1 1 48982
0 48984 7 1 2 88694 48983
0 48985 5 1 1 48984
0 48986 7 1 2 59650 97856
0 48987 7 1 2 88004 48986
0 48988 7 1 2 48985 48987
0 48989 5 1 1 48988
0 48990 7 1 2 48981 48989
0 48991 5 1 1 48990
0 48992 7 1 2 63837 48991
0 48993 5 1 1 48992
0 48994 7 1 2 81038 94743
0 48995 7 1 2 87497 48994
0 48996 7 1 2 97834 48995
0 48997 5 1 1 48996
0 48998 7 1 2 48993 48997
0 48999 7 1 2 48961 48998
0 49000 5 1 1 48999
0 49001 7 1 2 60404 49000
0 49002 5 1 1 49001
0 49003 7 1 2 79990 84124
0 49004 5 1 1 49003
0 49005 7 1 2 86409 86991
0 49006 5 1 1 49005
0 49007 7 1 2 63838 49006
0 49008 7 1 2 49004 49007
0 49009 5 1 1 49008
0 49010 7 1 2 79668 85710
0 49011 7 1 2 97836 49010
0 49012 5 1 1 49011
0 49013 7 1 2 49009 49012
0 49014 5 1 1 49013
0 49015 7 1 2 70677 49014
0 49016 5 1 1 49015
0 49017 7 2 2 87216 96081
0 49018 5 1 1 97864
0 49019 7 1 2 67380 94104
0 49020 5 1 1 49019
0 49021 7 1 2 49018 49020
0 49022 5 1 1 49021
0 49023 7 1 2 83939 49022
0 49024 5 1 1 49023
0 49025 7 1 2 80372 39823
0 49026 5 1 1 49025
0 49027 7 1 2 78381 85711
0 49028 7 1 2 49026 49027
0 49029 5 1 1 49028
0 49030 7 1 2 49024 49029
0 49031 5 1 1 49030
0 49032 7 1 2 67119 49031
0 49033 5 1 1 49032
0 49034 7 1 2 40162 49033
0 49035 7 2 2 85348 87217
0 49036 5 1 1 97866
0 49037 7 1 2 48905 49036
0 49038 5 1 1 49037
0 49039 7 1 2 66760 49038
0 49040 5 1 1 49039
0 49041 7 2 2 85872 90206
0 49042 7 1 2 82418 97868
0 49043 5 1 1 49042
0 49044 7 1 2 49040 49043
0 49045 5 1 1 49044
0 49046 7 1 2 72138 49045
0 49047 5 1 1 49046
0 49048 7 3 2 68772 91420
0 49049 7 1 2 74002 69467
0 49050 7 1 2 97870 49049
0 49051 5 1 1 49050
0 49052 7 1 2 96965 49051
0 49053 5 1 1 49052
0 49054 7 1 2 66900 49053
0 49055 5 1 1 49054
0 49056 7 1 2 49047 49055
0 49057 7 1 2 49034 49056
0 49058 5 1 1 49057
0 49059 7 1 2 68524 49058
0 49060 5 1 1 49059
0 49061 7 1 2 49016 49060
0 49062 5 1 1 49061
0 49063 7 1 2 95743 49062
0 49064 5 1 1 49063
0 49065 7 1 2 59969 97871
0 49066 5 1 1 49065
0 49067 7 1 2 92552 49066
0 49068 5 1 1 49067
0 49069 7 1 2 68525 49068
0 49070 5 1 1 49069
0 49071 7 1 2 89639 96096
0 49072 5 1 1 49071
0 49073 7 1 2 49070 49072
0 49074 5 1 1 49073
0 49075 7 1 2 66901 49074
0 49076 5 1 1 49075
0 49077 7 1 2 79949 75005
0 49078 5 1 1 49077
0 49079 7 1 2 86556 49078
0 49080 5 1 1 49079
0 49081 7 1 2 49076 49080
0 49082 5 1 1 49081
0 49083 7 4 2 59651 64135
0 49084 7 1 2 49082 97873
0 49085 5 1 1 49084
0 49086 7 1 2 60716 49085
0 49087 5 1 1 49086
0 49088 7 2 2 94729 96068
0 49089 5 1 1 97877
0 49090 7 1 2 84604 97878
0 49091 5 1 1 49090
0 49092 7 2 2 64136 80885
0 49093 7 1 2 61922 97879
0 49094 7 1 2 97645 49093
0 49095 5 1 1 49094
0 49096 7 1 2 49091 49095
0 49097 5 1 1 49096
0 49098 7 1 2 63839 49097
0 49099 5 1 1 49098
0 49100 7 1 2 79857 97433
0 49101 7 1 2 97872 49100
0 49102 5 1 1 49101
0 49103 7 1 2 65625 49102
0 49104 7 1 2 49099 49103
0 49105 5 1 1 49104
0 49106 7 1 2 59652 49105
0 49107 5 1 1 49106
0 49108 7 1 2 83566 96918
0 49109 7 1 2 94450 49108
0 49110 5 1 1 49109
0 49111 7 1 2 49107 49110
0 49112 5 1 1 49111
0 49113 7 1 2 69320 49112
0 49114 7 1 2 49087 49113
0 49115 5 1 1 49114
0 49116 7 1 2 49064 49115
0 49117 7 1 2 49002 49116
0 49118 7 1 2 48890 49117
0 49119 5 1 1 49118
0 49120 7 1 2 95300 49119
0 49121 5 1 1 49120
0 49122 7 1 2 83205 97824
0 49123 5 1 1 49122
0 49124 7 1 2 67742 49123
0 49125 5 1 1 49124
0 49126 7 2 2 68526 74609
0 49127 7 1 2 70543 97881
0 49128 5 1 1 49127
0 49129 7 1 2 49125 49128
0 49130 5 1 1 49129
0 49131 7 1 2 61923 95237
0 49132 7 1 2 97691 49131
0 49133 7 1 2 49130 49132
0 49134 5 1 1 49133
0 49135 7 1 2 49121 49134
0 49136 5 1 1 49135
0 49137 7 1 2 68934 49136
0 49138 5 1 1 49137
0 49139 7 1 2 96293 97746
0 49140 5 1 1 49139
0 49141 7 2 2 65626 87079
0 49142 7 3 2 97450 97883
0 49143 5 1 1 97885
0 49144 7 1 2 64046 97886
0 49145 5 1 1 49144
0 49146 7 1 2 49140 49145
0 49147 5 1 1 49146
0 49148 7 1 2 68773 49147
0 49149 5 1 1 49148
0 49150 7 4 2 64137 86284
0 49151 7 1 2 97822 97888
0 49152 5 1 1 49151
0 49153 7 1 2 49149 49152
0 49154 5 1 1 49153
0 49155 7 1 2 91689 49154
0 49156 5 1 1 49155
0 49157 7 2 2 94496 96519
0 49158 5 1 1 97892
0 49159 7 1 2 61792 97893
0 49160 5 1 1 49159
0 49161 7 1 2 86762 94081
0 49162 5 1 1 49161
0 49163 7 1 2 49160 49162
0 49164 5 1 1 49163
0 49165 7 1 2 90178 49164
0 49166 5 1 1 49165
0 49167 7 1 2 70678 92388
0 49168 7 1 2 95007 49167
0 49169 5 1 1 49168
0 49170 7 1 2 49166 49169
0 49171 5 1 1 49170
0 49172 7 1 2 64138 49171
0 49173 5 1 1 49172
0 49174 7 1 2 93664 94203
0 49175 7 1 2 97714 49174
0 49176 5 1 1 49175
0 49177 7 1 2 49173 49176
0 49178 7 1 2 49156 49177
0 49179 5 2 1 49178
0 49180 7 1 2 77011 97894
0 49181 5 1 1 49180
0 49182 7 1 2 81900 97693
0 49183 5 1 1 49182
0 49184 7 1 2 49181 49183
0 49185 5 1 1 49184
0 49186 7 1 2 95301 49185
0 49187 5 1 1 49186
0 49188 7 1 2 89859 95253
0 49189 7 1 2 80494 49188
0 49190 7 1 2 97027 49189
0 49191 7 1 2 97453 49190
0 49192 5 1 1 49191
0 49193 7 1 2 49187 49192
0 49194 5 1 1 49193
0 49195 7 1 2 91595 49194
0 49196 5 1 1 49195
0 49197 7 1 2 86772 90188
0 49198 5 2 1 49197
0 49199 7 3 2 86739 97896
0 49200 7 1 2 70863 97825
0 49201 5 1 1 49200
0 49202 7 1 2 59653 49201
0 49203 5 1 1 49202
0 49204 7 1 2 71427 86877
0 49205 5 1 1 49204
0 49206 7 1 2 70679 76411
0 49207 5 1 1 49206
0 49208 7 1 2 49205 49207
0 49209 7 1 2 49203 49208
0 49210 5 1 1 49209
0 49211 7 1 2 63579 49210
0 49212 5 1 1 49211
0 49213 7 1 2 69279 74886
0 49214 5 2 1 49213
0 49215 7 1 2 97524 97901
0 49216 5 1 1 49215
0 49217 7 1 2 49212 49216
0 49218 5 1 1 49217
0 49219 7 1 2 68774 49218
0 49220 5 1 1 49219
0 49221 7 1 2 72742 89712
0 49222 7 1 2 81713 49221
0 49223 5 1 1 49222
0 49224 7 1 2 49220 49223
0 49225 5 1 1 49224
0 49226 7 1 2 97898 49225
0 49227 5 1 1 49226
0 49228 7 1 2 70864 96799
0 49229 5 1 1 49228
0 49230 7 2 2 86763 49229
0 49231 7 1 2 92227 97903
0 49232 5 1 1 49231
0 49233 7 1 2 49227 49232
0 49234 5 1 1 49233
0 49235 7 1 2 64139 49234
0 49236 5 1 1 49235
0 49237 7 1 2 95209 97902
0 49238 5 1 1 49237
0 49239 7 1 2 85953 49238
0 49240 5 1 1 49239
0 49241 7 1 2 89025 49240
0 49242 5 1 1 49241
0 49243 7 1 2 92821 28926
0 49244 5 1 1 49243
0 49245 7 1 2 59970 49244
0 49246 5 1 1 49245
0 49247 7 1 2 69321 94042
0 49248 5 1 1 49247
0 49249 7 1 2 49246 49248
0 49250 5 1 1 49249
0 49251 7 1 2 68129 49250
0 49252 5 1 1 49251
0 49253 7 1 2 85933 49252
0 49254 5 1 1 49253
0 49255 7 1 2 65511 49254
0 49256 5 1 1 49255
0 49257 7 1 2 49242 49256
0 49258 5 1 1 49257
0 49259 7 1 2 68775 49258
0 49260 5 1 1 49259
0 49261 7 2 2 84125 83353
0 49262 5 1 1 97905
0 49263 7 1 2 68527 49262
0 49264 5 1 1 49263
0 49265 7 1 2 60182 74904
0 49266 5 1 1 49265
0 49267 7 1 2 49264 49266
0 49268 5 1 1 49267
0 49269 7 1 2 68130 49268
0 49270 5 1 1 49269
0 49271 7 1 2 83761 95612
0 49272 5 1 1 49271
0 49273 7 1 2 59654 49272
0 49274 5 1 1 49273
0 49275 7 1 2 82275 97646
0 49276 5 1 1 49275
0 49277 7 1 2 89529 49276
0 49278 7 1 2 49274 49277
0 49279 5 1 1 49278
0 49280 7 1 2 67381 49279
0 49281 5 1 1 49280
0 49282 7 1 2 48085 49281
0 49283 5 1 1 49282
0 49284 7 1 2 60947 49283
0 49285 5 1 1 49284
0 49286 7 1 2 49270 49285
0 49287 5 1 1 49286
0 49288 7 1 2 92228 49287
0 49289 5 1 1 49288
0 49290 7 1 2 49260 49289
0 49291 5 1 1 49290
0 49292 7 1 2 97400 49291
0 49293 5 1 1 49292
0 49294 7 1 2 49236 49293
0 49295 5 1 1 49294
0 49296 7 1 2 61793 49295
0 49297 5 1 1 49296
0 49298 7 2 2 77012 86860
0 49299 7 1 2 66761 97907
0 49300 5 1 1 49299
0 49301 7 1 2 28400 49300
0 49302 5 1 1 49301
0 49303 7 1 2 70680 49302
0 49304 5 1 1 49303
0 49305 7 1 2 81452 97906
0 49306 5 1 1 49305
0 49307 7 1 2 92284 49306
0 49308 5 1 1 49307
0 49309 7 1 2 49304 49308
0 49310 5 1 1 49309
0 49311 7 1 2 68131 49310
0 49312 5 1 1 49311
0 49313 7 1 2 75053 97632
0 49314 5 1 1 49313
0 49315 7 1 2 67743 97635
0 49316 5 1 1 49315
0 49317 7 1 2 49314 49316
0 49318 5 1 1 49317
0 49319 7 1 2 83251 49318
0 49320 5 1 1 49319
0 49321 7 1 2 49312 49320
0 49322 5 1 1 49321
0 49323 7 1 2 96919 49322
0 49324 5 1 1 49323
0 49325 7 1 2 64140 97904
0 49326 5 1 1 49325
0 49327 7 1 2 49324 49326
0 49328 5 1 1 49327
0 49329 7 1 2 63840 49328
0 49330 5 1 1 49329
0 49331 7 2 2 82590 76306
0 49332 7 1 2 96670 97628
0 49333 7 1 2 97909 49332
0 49334 5 1 1 49333
0 49335 7 1 2 49330 49334
0 49336 5 1 1 49335
0 49337 7 1 2 90179 49336
0 49338 5 1 1 49337
0 49339 7 1 2 80044 97652
0 49340 5 1 1 49339
0 49341 7 1 2 83252 89814
0 49342 7 1 2 97650 49341
0 49343 5 1 1 49342
0 49344 7 1 2 49340 49343
0 49345 5 1 1 49344
0 49346 7 1 2 70681 49345
0 49347 5 1 1 49346
0 49348 7 1 2 65512 96396
0 49349 5 1 1 49348
0 49350 7 1 2 85758 49349
0 49351 5 1 1 49350
0 49352 7 1 2 97653 49351
0 49353 5 1 1 49352
0 49354 7 1 2 49347 49353
0 49355 5 1 1 49354
0 49356 7 1 2 67744 49355
0 49357 5 1 1 49356
0 49358 7 1 2 75099 85048
0 49359 5 1 1 49358
0 49360 7 1 2 85412 49359
0 49361 5 1 1 49360
0 49362 7 1 2 97882 49361
0 49363 5 1 1 49362
0 49364 7 1 2 70682 97908
0 49365 5 1 1 49364
0 49366 7 1 2 49363 49365
0 49367 5 1 1 49366
0 49368 7 1 2 97654 49367
0 49369 5 1 1 49368
0 49370 7 1 2 49357 49369
0 49371 5 1 1 49370
0 49372 7 1 2 68132 49371
0 49373 5 1 1 49372
0 49374 7 1 2 1135 1159
0 49375 5 1 1 49374
0 49376 7 1 2 96765 97853
0 49377 7 1 2 49375 49376
0 49378 5 1 1 49377
0 49379 7 1 2 49373 49378
0 49380 5 1 1 49379
0 49381 7 1 2 86802 49380
0 49382 5 1 1 49381
0 49383 7 1 2 97683 97910
0 49384 5 1 1 49383
0 49385 7 1 2 59971 97368
0 49386 5 1 1 49385
0 49387 7 1 2 80959 87612
0 49388 5 2 1 49387
0 49389 7 1 2 49386 97911
0 49390 5 1 1 49389
0 49391 7 1 2 95632 49390
0 49392 5 1 1 49391
0 49393 7 2 2 78265 97749
0 49394 5 1 1 97913
0 49395 7 1 2 75027 97914
0 49396 5 1 1 49395
0 49397 7 4 2 87623 97434
0 49398 5 1 1 97915
0 49399 7 1 2 78465 97916
0 49400 5 1 1 49399
0 49401 7 4 2 92285 94730
0 49402 5 1 1 97919
0 49403 7 1 2 49400 49402
0 49404 7 1 2 49396 49403
0 49405 5 1 1 49404
0 49406 7 1 2 70683 49405
0 49407 5 1 1 49406
0 49408 7 1 2 91532 97887
0 49409 5 1 1 49408
0 49410 7 1 2 49407 49409
0 49411 7 1 2 49392 49410
0 49412 5 1 1 49411
0 49413 7 1 2 68776 49412
0 49414 5 1 1 49413
0 49415 7 1 2 77801 94717
0 49416 7 2 2 96720 49415
0 49417 5 1 1 97923
0 49418 7 2 2 63841 64141
0 49419 7 3 2 68528 97925
0 49420 7 1 2 95699 97927
0 49421 5 1 1 49420
0 49422 7 1 2 97415 49421
0 49423 5 1 1 49422
0 49424 7 1 2 59655 89522
0 49425 7 1 2 49423 49424
0 49426 5 1 1 49425
0 49427 7 1 2 49417 49426
0 49428 5 1 1 49427
0 49429 7 1 2 77013 49428
0 49430 5 1 1 49429
0 49431 7 1 2 80932 97730
0 49432 7 3 2 61924 76505
0 49433 7 2 2 78782 97732
0 49434 7 1 2 97930 97933
0 49435 7 1 2 49431 49434
0 49436 5 1 1 49435
0 49437 7 1 2 49430 49436
0 49438 7 1 2 49414 49437
0 49439 5 1 1 49438
0 49440 7 1 2 91690 49439
0 49441 5 1 1 49440
0 49442 7 1 2 49384 49441
0 49443 7 1 2 49382 49442
0 49444 7 1 2 49338 49443
0 49445 7 1 2 49297 49444
0 49446 5 1 1 49445
0 49447 7 1 2 97763 49446
0 49448 5 1 1 49447
0 49449 7 1 2 49196 49448
0 49450 7 1 2 49138 49449
0 49451 7 1 2 48797 49450
0 49452 7 1 2 48177 49451
0 49453 5 1 1 49452
0 49454 7 1 2 69961 49453
0 49455 5 1 1 49454
0 49456 7 1 2 88199 96941
0 49457 5 1 1 49456
0 49458 7 1 2 91607 90058
0 49459 7 1 2 96979 49458
0 49460 5 1 1 49459
0 49461 7 1 2 49457 49460
0 49462 5 1 1 49461
0 49463 7 1 2 71013 49462
0 49464 5 1 1 49463
0 49465 7 1 2 80886 90117
0 49466 5 1 1 49465
0 49467 7 3 2 66762 84307
0 49468 5 3 1 97935
0 49469 7 1 2 84556 97938
0 49470 5 2 1 49469
0 49471 7 1 2 70684 86144
0 49472 7 1 2 97941 49471
0 49473 5 1 1 49472
0 49474 7 1 2 49466 49473
0 49475 5 1 1 49474
0 49476 7 1 2 76269 49475
0 49477 5 1 1 49476
0 49478 7 1 2 91827 88715
0 49479 5 1 1 49478
0 49480 7 1 2 77036 97936
0 49481 5 1 1 49480
0 49482 7 1 2 49479 49481
0 49483 5 1 1 49482
0 49484 7 1 2 68529 49483
0 49485 5 1 1 49484
0 49486 7 1 2 86455 97789
0 49487 5 2 1 49486
0 49488 7 1 2 49485 97943
0 49489 5 1 1 49488
0 49490 7 1 2 68935 49489
0 49491 5 1 1 49490
0 49492 7 1 2 49477 49491
0 49493 5 1 1 49492
0 49494 7 1 2 60948 49493
0 49495 5 1 1 49494
0 49496 7 4 2 80638 90812
0 49497 7 1 2 86612 97945
0 49498 7 1 2 97497 49497
0 49499 5 1 1 49498
0 49500 7 1 2 49495 49499
0 49501 5 1 1 49500
0 49502 7 1 2 67382 49501
0 49503 5 1 1 49502
0 49504 7 1 2 27906 42244
0 49505 5 1 1 49504
0 49506 7 1 2 69587 49505
0 49507 5 1 1 49506
0 49508 7 1 2 81761 92453
0 49509 5 1 1 49508
0 49510 7 1 2 49507 49509
0 49511 5 1 1 49510
0 49512 7 1 2 80960 49511
0 49513 5 1 1 49512
0 49514 7 1 2 49503 49513
0 49515 5 1 1 49514
0 49516 7 1 2 64142 49515
0 49517 5 1 1 49516
0 49518 7 1 2 49464 49517
0 49519 5 1 1 49518
0 49520 7 1 2 68133 49519
0 49521 5 1 1 49520
0 49522 7 1 2 59656 94612
0 49523 5 2 1 49522
0 49524 7 2 2 89942 94757
0 49525 7 1 2 92480 97951
0 49526 5 2 1 49525
0 49527 7 1 2 97949 97953
0 49528 5 1 1 49527
0 49529 7 1 2 69588 49528
0 49530 5 1 1 49529
0 49531 7 1 2 86303 96980
0 49532 5 3 1 49531
0 49533 7 1 2 84100 94613
0 49534 5 1 1 49533
0 49535 7 1 2 97955 49534
0 49536 5 1 1 49535
0 49537 7 1 2 69322 49536
0 49538 5 1 1 49537
0 49539 7 2 2 69016 86221
0 49540 7 1 2 88273 97958
0 49541 5 1 1 49540
0 49542 7 1 2 97954 49541
0 49543 5 1 1 49542
0 49544 7 1 2 59657 49543
0 49545 5 1 1 49544
0 49546 7 1 2 49538 49545
0 49547 7 1 2 49530 49546
0 49548 5 1 1 49547
0 49549 7 1 2 66763 49548
0 49550 5 1 1 49549
0 49551 7 1 2 78881 91163
0 49552 5 1 1 49551
0 49553 7 1 2 83220 49552
0 49554 5 1 1 49553
0 49555 7 1 2 79669 49554
0 49556 5 1 1 49555
0 49557 7 1 2 85293 49556
0 49558 5 1 1 49557
0 49559 7 1 2 94758 49558
0 49560 5 1 1 49559
0 49561 7 1 2 49550 49560
0 49562 7 1 2 49521 49561
0 49563 5 1 1 49562
0 49564 7 1 2 61126 49563
0 49565 5 1 1 49564
0 49566 7 1 2 70685 84399
0 49567 5 1 1 49566
0 49568 7 1 2 88754 97305
0 49569 5 1 1 49568
0 49570 7 1 2 49567 49569
0 49571 5 1 1 49570
0 49572 7 1 2 78783 49571
0 49573 5 1 1 49572
0 49574 7 1 2 63192 88675
0 49575 5 1 1 49574
0 49576 7 1 2 68777 93870
0 49577 7 1 2 49575 49576
0 49578 5 1 1 49577
0 49579 7 1 2 49573 49578
0 49580 5 1 1 49579
0 49581 7 1 2 79670 49580
0 49582 5 1 1 49581
0 49583 7 3 2 79445 86436
0 49584 5 1 1 97960
0 49585 7 1 2 83064 97164
0 49586 5 1 1 49585
0 49587 7 1 2 49584 49586
0 49588 5 1 1 49587
0 49589 7 1 2 69589 49588
0 49590 5 1 1 49589
0 49591 7 1 2 75054 89753
0 49592 5 1 1 49591
0 49593 7 1 2 49590 49592
0 49594 5 1 1 49593
0 49595 7 1 2 81262 49594
0 49596 5 1 1 49595
0 49597 7 1 2 85294 49596
0 49598 5 1 1 49597
0 49599 7 1 2 60949 49598
0 49600 5 1 1 49599
0 49601 7 2 2 69709 89599
0 49602 5 1 1 97963
0 49603 7 1 2 83155 49602
0 49604 5 1 1 49603
0 49605 7 1 2 49600 49604
0 49606 7 1 2 49582 49605
0 49607 5 1 1 49606
0 49608 7 1 2 68936 49607
0 49609 5 1 1 49608
0 49610 7 1 2 76270 89860
0 49611 7 1 2 97394 49610
0 49612 5 1 1 49611
0 49613 7 1 2 49609 49612
0 49614 5 1 1 49613
0 49615 7 1 2 64143 49614
0 49616 5 1 1 49615
0 49617 7 1 2 76456 96391
0 49618 5 2 1 49617
0 49619 7 2 2 82984 92630
0 49620 7 1 2 94228 97967
0 49621 7 1 2 97965 49620
0 49622 5 1 1 49621
0 49623 7 1 2 49616 49622
0 49624 7 1 2 49565 49623
0 49625 5 1 1 49624
0 49626 7 1 2 59972 49625
0 49627 5 1 1 49626
0 49628 7 2 2 81811 93238
0 49629 5 1 1 97969
0 49630 7 4 2 68134 92501
0 49631 7 1 2 97970 97971
0 49632 5 1 1 49631
0 49633 7 1 2 80909 49632
0 49634 5 1 1 49633
0 49635 7 1 2 67120 49634
0 49636 5 1 1 49635
0 49637 7 1 2 96370 96778
0 49638 5 1 1 49637
0 49639 7 1 2 49636 49638
0 49640 5 1 1 49639
0 49641 7 1 2 94759 49640
0 49642 5 1 1 49641
0 49643 7 2 2 83110 96330
0 49644 7 1 2 74140 84269
0 49645 7 1 2 97975 49644
0 49646 5 1 1 49645
0 49647 7 1 2 49642 49646
0 49648 5 1 1 49647
0 49649 7 1 2 67383 49648
0 49650 5 1 1 49649
0 49651 7 1 2 92649 94760
0 49652 5 1 1 49651
0 49653 7 1 2 75100 85370
0 49654 7 1 2 97793 49653
0 49655 5 1 1 49654
0 49656 7 1 2 49652 49655
0 49657 7 1 2 49650 49656
0 49658 5 1 1 49657
0 49659 7 1 2 60950 49658
0 49660 5 1 1 49659
0 49661 7 1 2 63193 81825
0 49662 5 2 1 49661
0 49663 7 2 2 79671 86304
0 49664 7 1 2 97977 97979
0 49665 5 1 1 49664
0 49666 7 2 2 60610 89815
0 49667 5 1 1 97981
0 49668 7 1 2 67745 97982
0 49669 5 1 1 49668
0 49670 7 1 2 49665 49669
0 49671 5 1 1 49670
0 49672 7 1 2 94761 49671
0 49673 5 1 1 49672
0 49674 7 1 2 49660 49673
0 49675 5 1 1 49674
0 49676 7 1 2 59658 49675
0 49677 5 1 1 49676
0 49678 7 3 2 66764 97976
0 49679 5 1 1 97983
0 49680 7 1 2 70865 36065
0 49681 5 1 1 49680
0 49682 7 1 2 97984 49681
0 49683 5 1 1 49682
0 49684 7 1 2 75758 91177
0 49685 5 1 1 49684
0 49686 7 1 2 97980 49685
0 49687 5 1 1 49686
0 49688 7 1 2 83111 84942
0 49689 7 1 2 35254 49688
0 49690 5 1 1 49689
0 49691 7 1 2 80887 49690
0 49692 5 1 1 49691
0 49693 7 1 2 49687 49692
0 49694 5 1 1 49693
0 49695 7 1 2 94762 49694
0 49696 5 1 1 49695
0 49697 7 1 2 49683 49696
0 49698 7 1 2 49677 49697
0 49699 5 1 1 49698
0 49700 7 1 2 63842 49699
0 49701 5 1 1 49700
0 49702 7 1 2 96639 97447
0 49703 5 1 1 49702
0 49704 7 1 2 79672 96481
0 49705 5 1 1 49704
0 49706 7 1 2 60611 89863
0 49707 5 1 1 49706
0 49708 7 1 2 49705 49707
0 49709 5 1 1 49708
0 49710 7 1 2 94763 49709
0 49711 5 1 1 49710
0 49712 7 1 2 77440 94712
0 49713 5 1 1 49712
0 49714 7 1 2 49711 49713
0 49715 5 1 1 49714
0 49716 7 1 2 69729 49715
0 49717 5 1 1 49716
0 49718 7 1 2 49703 49717
0 49719 5 1 1 49718
0 49720 7 1 2 72139 49719
0 49721 5 1 1 49720
0 49722 7 1 2 63194 91274
0 49723 5 1 1 49722
0 49724 7 1 2 69590 49723
0 49725 5 2 1 49724
0 49726 7 1 2 61127 90102
0 49727 5 1 1 49726
0 49728 7 1 2 97986 49727
0 49729 5 1 1 49728
0 49730 7 1 2 67384 49729
0 49731 5 1 1 49730
0 49732 7 1 2 78275 49731
0 49733 5 2 1 49732
0 49734 7 1 2 79446 97988
0 49735 5 1 1 49734
0 49736 7 1 2 96439 49735
0 49737 5 1 1 49736
0 49738 7 1 2 70686 49737
0 49739 5 1 1 49738
0 49740 7 1 2 80365 93874
0 49741 5 1 1 49740
0 49742 7 1 2 66077 76242
0 49743 5 4 1 49742
0 49744 7 1 2 77441 97990
0 49745 5 1 1 49744
0 49746 7 1 2 81448 78438
0 49747 5 1 1 49746
0 49748 7 1 2 49745 49747
0 49749 5 1 1 49748
0 49750 7 1 2 94408 49749
0 49751 5 1 1 49750
0 49752 7 1 2 49741 49751
0 49753 7 1 2 49739 49752
0 49754 5 1 1 49753
0 49755 7 1 2 68937 49754
0 49756 5 1 1 49755
0 49757 7 1 2 70687 18723
0 49758 5 1 1 49757
0 49759 7 1 2 76271 93267
0 49760 5 1 1 49759
0 49761 7 1 2 49758 49760
0 49762 5 1 1 49761
0 49763 7 1 2 82034 13390
0 49764 7 1 2 49762 49763
0 49765 5 1 1 49764
0 49766 7 1 2 49756 49765
0 49767 5 1 1 49766
0 49768 7 1 2 94718 49767
0 49769 5 1 1 49768
0 49770 7 1 2 49721 49769
0 49771 7 1 2 49701 49770
0 49772 7 1 2 49627 49771
0 49773 5 1 1 49772
0 49774 7 1 2 86803 49773
0 49775 5 1 1 49774
0 49776 7 2 2 79447 96331
0 49777 5 1 1 97994
0 49778 7 2 2 91363 89861
0 49779 7 1 2 94764 97996
0 49780 5 1 1 49779
0 49781 7 1 2 49777 49780
0 49782 5 1 1 49781
0 49783 7 1 2 97502 49782
0 49784 5 1 1 49783
0 49785 7 2 2 82001 94765
0 49786 7 1 2 69202 91364
0 49787 7 1 2 97998 49786
0 49788 5 1 1 49787
0 49789 7 1 2 49784 49788
0 49790 5 1 1 49789
0 49791 7 1 2 68778 49790
0 49792 5 1 1 49791
0 49793 7 4 2 63580 94217
0 49794 7 1 2 91346 96886
0 49795 7 1 2 98000 49794
0 49796 5 1 1 49795
0 49797 7 1 2 49792 49796
0 49798 5 1 1 49797
0 49799 7 1 2 65627 49798
0 49800 5 1 1 49799
0 49801 7 1 2 92168 96678
0 49802 7 1 2 96779 97101
0 49803 7 1 2 49801 49802
0 49804 5 1 1 49803
0 49805 7 1 2 49800 49804
0 49806 5 1 1 49805
0 49807 7 1 2 66902 49806
0 49808 5 1 1 49807
0 49809 7 2 2 64047 64144
0 49810 7 2 2 69203 83567
0 49811 5 1 1 98006
0 49812 7 1 2 96266 49811
0 49813 5 1 1 49812
0 49814 7 1 2 61925 49813
0 49815 5 1 1 49814
0 49816 7 1 2 61926 83589
0 49817 5 2 1 49816
0 49818 7 2 2 61794 98007
0 49819 5 1 1 98010
0 49820 7 1 2 98008 49819
0 49821 5 1 1 49820
0 49822 7 1 2 60612 49821
0 49823 5 1 1 49822
0 49824 7 1 2 49815 49823
0 49825 5 1 1 49824
0 49826 7 1 2 60717 49825
0 49827 5 1 1 49826
0 49828 7 1 2 96246 98011
0 49829 5 1 1 49828
0 49830 7 1 2 49827 49829
0 49831 5 1 1 49830
0 49832 7 1 2 70688 49831
0 49833 5 1 1 49832
0 49834 7 1 2 79673 76412
0 49835 7 1 2 97417 49834
0 49836 5 1 1 49835
0 49837 7 1 2 49833 49836
0 49838 5 1 1 49837
0 49839 7 1 2 98004 49838
0 49840 5 1 1 49839
0 49841 7 1 2 49808 49840
0 49842 5 1 1 49841
0 49843 7 1 2 69591 49842
0 49844 5 1 1 49843
0 49845 7 1 2 91975 92562
0 49846 5 1 1 49845
0 49847 7 1 2 40262 49846
0 49848 5 1 1 49847
0 49849 7 1 2 60613 49848
0 49850 5 1 1 49849
0 49851 7 1 2 60951 89864
0 49852 5 1 1 49851
0 49853 7 1 2 8072 49852
0 49854 5 1 1 49853
0 49855 7 1 2 61927 49854
0 49856 5 1 1 49855
0 49857 7 1 2 49850 49856
0 49858 5 1 1 49857
0 49859 7 1 2 60718 49858
0 49860 5 1 1 49859
0 49861 7 2 2 81112 96573
0 49862 7 1 2 91365 98012
0 49863 5 1 1 49862
0 49864 7 1 2 49860 49863
0 49865 5 1 1 49864
0 49866 7 1 2 97468 49865
0 49867 5 1 1 49866
0 49868 7 1 2 96920 97707
0 49869 5 2 1 49868
0 49870 7 15 2 60719 97435
0 49871 5 3 1 98016
0 49872 7 1 2 81604 98017
0 49873 5 1 1 49872
0 49874 7 1 2 98014 49873
0 49875 5 1 1 49874
0 49876 7 1 2 91828 49875
0 49877 5 1 1 49876
0 49878 7 1 2 70689 97444
0 49879 5 1 1 49878
0 49880 7 1 2 48348 49879
0 49881 5 1 1 49880
0 49882 7 1 2 84366 49881
0 49883 5 1 1 49882
0 49884 7 1 2 49877 49883
0 49885 5 1 1 49884
0 49886 7 1 2 68530 49885
0 49887 5 1 1 49886
0 49888 7 1 2 97677 49887
0 49889 7 1 2 49867 49888
0 49890 5 1 1 49889
0 49891 7 1 2 64048 49890
0 49892 5 1 1 49891
0 49893 7 1 2 82358 91424
0 49894 7 2 2 65628 96421
0 49895 7 1 2 96981 98034
0 49896 7 1 2 49893 49895
0 49897 5 1 1 49896
0 49898 7 1 2 49892 49897
0 49899 7 1 2 49844 49898
0 49900 5 1 1 49899
0 49901 7 1 2 59659 49900
0 49902 5 1 1 49901
0 49903 7 6 2 92286 96921
0 49904 5 1 1 98036
0 49905 7 1 2 69592 98037
0 49906 5 1 1 49905
0 49907 7 1 2 63195 81462
0 49908 5 1 1 49907
0 49909 7 1 2 95633 49908
0 49910 5 1 1 49909
0 49911 7 1 2 49906 49910
0 49912 5 1 1 49911
0 49913 7 1 2 91829 49912
0 49914 5 1 1 49913
0 49915 7 2 2 79448 96922
0 49916 7 1 2 96540 98042
0 49917 5 1 1 49916
0 49918 7 1 2 68135 95145
0 49919 7 1 2 96533 49918
0 49920 5 1 1 49919
0 49921 7 1 2 49917 49920
0 49922 5 1 1 49921
0 49923 7 1 2 67121 49922
0 49924 5 1 1 49923
0 49925 7 1 2 49143 49924
0 49926 5 1 1 49925
0 49927 7 1 2 68779 49926
0 49928 5 1 1 49927
0 49929 7 1 2 49914 49928
0 49930 5 1 1 49929
0 49931 7 1 2 70690 49930
0 49932 5 1 1 49931
0 49933 7 1 2 91164 97401
0 49934 5 1 1 49933
0 49935 7 1 2 95718 95733
0 49936 7 1 2 97928 49935
0 49937 5 1 1 49936
0 49938 7 1 2 49934 49937
0 49939 5 1 1 49938
0 49940 7 1 2 69593 49939
0 49941 5 1 1 49940
0 49942 7 2 2 96901 98035
0 49943 5 1 1 98044
0 49944 7 1 2 49941 49943
0 49945 5 1 1 49944
0 49946 7 1 2 67385 49945
0 49947 5 1 1 49946
0 49948 7 1 2 89713 98018
0 49949 5 2 1 49948
0 49950 7 1 2 49947 98046
0 49951 5 1 1 49950
0 49952 7 1 2 79674 49951
0 49953 5 1 1 49952
0 49954 7 1 2 67122 97674
0 49955 5 1 1 49954
0 49956 7 1 2 69594 92314
0 49957 7 1 2 96909 49956
0 49958 5 1 1 49957
0 49959 7 1 2 49955 49958
0 49960 7 1 2 49953 49959
0 49961 7 1 2 49932 49960
0 49962 5 1 1 49961
0 49963 7 1 2 64049 49962
0 49964 5 1 1 49963
0 49965 7 3 2 63843 96999
0 49966 7 1 2 78482 98048
0 49967 5 1 1 49966
0 49968 7 1 2 65629 89061
0 49969 7 1 2 96184 49968
0 49970 5 1 1 49969
0 49971 7 1 2 49967 49970
0 49972 5 1 1 49971
0 49973 7 1 2 78382 49972
0 49974 5 1 1 49973
0 49975 7 1 2 34647 49974
0 49976 5 1 1 49975
0 49977 7 1 2 60614 97596
0 49978 7 1 2 49976 49977
0 49979 5 1 1 49978
0 49980 7 1 2 49964 49979
0 49981 7 1 2 49902 49980
0 49982 5 1 1 49981
0 49983 7 1 2 67746 49982
0 49984 5 1 1 49983
0 49985 7 1 2 21877 95107
0 49986 5 1 1 49985
0 49987 7 1 2 81614 90157
0 49988 7 1 2 98049 49987
0 49989 5 1 1 49988
0 49990 7 1 2 49986 49989
0 49991 5 1 1 49990
0 49992 7 1 2 92007 49991
0 49993 5 1 1 49992
0 49994 7 1 2 20904 49993
0 49995 5 1 1 49994
0 49996 7 1 2 94766 49995
0 49997 5 1 1 49996
0 49998 7 3 2 91830 98019
0 49999 5 1 1 98051
0 50000 7 1 2 97620 49999
0 50001 5 3 1 50000
0 50002 7 1 2 78148 96840
0 50003 5 1 1 50002
0 50004 7 1 2 98054 50003
0 50005 5 1 1 50004
0 50006 7 2 2 94719 96534
0 50007 7 1 2 77930 95133
0 50008 5 1 1 50007
0 50009 7 1 2 85954 50008
0 50010 5 1 1 50009
0 50011 7 1 2 98057 50010
0 50012 5 1 1 50011
0 50013 7 3 2 91831 98038
0 50014 5 1 1 98059
0 50015 7 2 2 67386 81588
0 50016 5 1 1 98062
0 50017 7 1 2 63196 50016
0 50018 5 1 1 50017
0 50019 7 1 2 98060 50018
0 50020 5 1 1 50019
0 50021 7 1 2 50012 50020
0 50022 7 1 2 50005 50021
0 50023 5 1 1 50022
0 50024 7 1 2 70691 50023
0 50025 5 1 1 50024
0 50026 7 2 2 89953 98020
0 50027 7 1 2 90158 98064
0 50028 5 1 1 50027
0 50029 7 1 2 67387 98045
0 50030 5 1 1 50029
0 50031 7 1 2 98047 50030
0 50032 5 1 1 50031
0 50033 7 1 2 67123 79675
0 50034 7 1 2 50032 50033
0 50035 5 1 1 50034
0 50036 7 1 2 50028 50035
0 50037 5 1 1 50036
0 50038 7 1 2 76272 50037
0 50039 5 1 1 50038
0 50040 7 2 2 60615 85712
0 50041 7 2 2 97584 98066
0 50042 5 1 1 98068
0 50043 7 1 2 68136 98069
0 50044 5 2 1 50043
0 50045 7 1 2 92502 97640
0 50046 5 1 1 50045
0 50047 7 3 2 94934 96923
0 50048 5 1 1 98072
0 50049 7 1 2 50046 50048
0 50050 5 2 1 50049
0 50051 7 1 2 69204 98075
0 50052 5 1 1 50051
0 50053 7 1 2 63197 77053
0 50054 5 5 1 50053
0 50055 7 1 2 98077 98073
0 50056 5 1 1 50055
0 50057 7 1 2 50052 50056
0 50058 5 1 1 50057
0 50059 7 1 2 63844 50058
0 50060 5 1 1 50059
0 50061 7 1 2 98070 50060
0 50062 7 1 2 50039 50061
0 50063 7 1 2 50025 50062
0 50064 5 1 1 50063
0 50065 7 1 2 64050 50064
0 50066 5 1 1 50065
0 50067 7 1 2 49997 50066
0 50068 7 1 2 49984 50067
0 50069 5 1 1 50068
0 50070 7 1 2 61128 50069
0 50071 5 1 1 50070
0 50072 7 3 2 60952 78383
0 50073 5 4 1 98082
0 50074 7 1 2 78299 88701
0 50075 5 1 1 50074
0 50076 7 1 2 67124 50075
0 50077 5 1 1 50076
0 50078 7 1 2 98085 50077
0 50079 5 1 1 50078
0 50080 7 1 2 59660 50079
0 50081 5 1 1 50080
0 50082 7 1 2 80075 82995
0 50083 5 1 1 50082
0 50084 7 2 2 50081 50083
0 50085 5 1 1 98089
0 50086 7 1 2 63581 98090
0 50087 5 1 1 50086
0 50088 7 2 2 96171 50087
0 50089 7 1 2 60720 98091
0 50090 5 1 1 50089
0 50091 7 3 2 69205 77931
0 50092 5 1 1 98093
0 50093 7 1 2 98094 97966
0 50094 5 1 1 50093
0 50095 7 1 2 97912 50094
0 50096 5 1 1 50095
0 50097 7 1 2 68780 96535
0 50098 7 1 2 50096 50097
0 50099 5 1 1 50098
0 50100 7 1 2 50090 50099
0 50101 5 1 1 50100
0 50102 7 1 2 64145 50101
0 50103 5 1 1 50102
0 50104 7 1 2 77037 96182
0 50105 5 1 1 50104
0 50106 7 1 2 65904 97964
0 50107 5 1 1 50106
0 50108 7 1 2 91832 50107
0 50109 5 1 1 50108
0 50110 7 1 2 50105 50109
0 50111 5 1 1 50110
0 50112 7 1 2 68137 50111
0 50113 5 1 1 50112
0 50114 7 1 2 79293 86437
0 50115 5 3 1 50114
0 50116 7 1 2 67388 96286
0 50117 5 1 1 50116
0 50118 7 1 2 98096 50117
0 50119 5 1 1 50118
0 50120 7 1 2 76273 50119
0 50121 5 1 1 50120
0 50122 7 1 2 81812 73451
0 50123 5 2 1 50122
0 50124 7 1 2 63198 98099
0 50125 5 2 1 50124
0 50126 7 2 2 59661 98101
0 50127 5 1 1 98103
0 50128 7 1 2 92443 98104
0 50129 5 1 1 50128
0 50130 7 1 2 50121 50129
0 50131 5 1 1 50130
0 50132 7 1 2 60953 50131
0 50133 5 1 1 50132
0 50134 7 1 2 50113 50133
0 50135 5 1 1 50134
0 50136 7 1 2 98039 50135
0 50137 5 1 1 50136
0 50138 7 1 2 50103 50137
0 50139 5 1 1 50138
0 50140 7 1 2 70692 50139
0 50141 5 1 1 50140
0 50142 7 1 2 19906 89956
0 50143 5 1 1 50142
0 50144 7 1 2 97402 50143
0 50145 5 1 1 50144
0 50146 7 1 2 97616 50145
0 50147 5 1 1 50146
0 50148 7 1 2 60616 50147
0 50149 5 2 1 50148
0 50150 7 1 2 59662 97684
0 50151 5 1 1 50150
0 50152 7 1 2 73360 97675
0 50153 5 1 1 50152
0 50154 7 1 2 50151 50153
0 50155 5 1 1 50154
0 50156 7 1 2 67747 50155
0 50157 5 1 1 50156
0 50158 7 1 2 96238 97669
0 50159 5 1 1 50158
0 50160 7 1 2 86358 92315
0 50161 7 1 2 96671 50160
0 50162 5 1 1 50161
0 50163 7 1 2 50159 50162
0 50164 5 1 1 50163
0 50165 7 1 2 69595 50164
0 50166 5 1 1 50165
0 50167 7 1 2 50166 98071
0 50168 7 2 2 50157 50167
0 50169 5 1 1 98107
0 50170 7 1 2 93989 96902
0 50171 5 1 1 50170
0 50172 7 1 2 97308 98021
0 50173 5 1 1 50172
0 50174 7 1 2 50171 50173
0 50175 5 1 1 50174
0 50176 7 1 2 69596 50175
0 50177 5 1 1 50176
0 50178 7 1 2 75055 89714
0 50179 7 1 2 98022 50178
0 50180 5 1 1 50179
0 50181 7 1 2 50177 50180
0 50182 5 2 1 50181
0 50183 7 1 2 79676 98109
0 50184 5 1 1 50183
0 50185 7 1 2 98108 50184
0 50186 5 1 1 50185
0 50187 7 1 2 69206 50186
0 50188 5 1 1 50187
0 50189 7 1 2 98105 50188
0 50190 7 1 2 50141 50189
0 50191 5 1 1 50190
0 50192 7 1 2 64051 50191
0 50193 5 1 1 50192
0 50194 7 2 2 86725 96848
0 50195 7 1 2 97838 98111
0 50196 5 2 1 50195
0 50197 7 1 2 83071 88119
0 50198 5 1 1 50197
0 50199 7 1 2 97348 50198
0 50200 5 1 1 50199
0 50201 7 1 2 80784 91405
0 50202 7 1 2 50200 50201
0 50203 5 1 1 50202
0 50204 7 1 2 97484 50203
0 50205 5 1 1 50204
0 50206 7 1 2 76274 50205
0 50207 5 1 1 50206
0 50208 7 1 2 76413 87624
0 50209 5 1 1 50208
0 50210 7 1 2 60617 97946
0 50211 7 1 2 97362 50210
0 50212 5 1 1 50211
0 50213 7 1 2 50209 50212
0 50214 5 1 1 50213
0 50215 7 1 2 66765 50214
0 50216 5 1 1 50215
0 50217 7 1 2 50207 50216
0 50218 5 1 1 50217
0 50219 7 1 2 61928 50218
0 50220 5 1 1 50219
0 50221 7 1 2 60183 92105
0 50222 7 2 2 95811 50221
0 50223 7 1 2 86484 88692
0 50224 7 1 2 98115 50223
0 50225 5 1 1 50224
0 50226 7 1 2 50220 50225
0 50227 5 1 1 50226
0 50228 7 1 2 63845 50227
0 50229 5 1 1 50228
0 50230 7 1 2 62769 81621
0 50231 5 2 1 50230
0 50232 7 3 2 70693 80888
0 50233 7 1 2 94635 96541
0 50234 7 1 2 98119 50233
0 50235 7 1 2 98117 50234
0 50236 5 1 1 50235
0 50237 7 1 2 50229 50236
0 50238 5 1 1 50237
0 50239 7 1 2 64146 50238
0 50240 5 1 1 50239
0 50241 7 1 2 98113 50240
0 50242 5 1 1 50241
0 50243 7 1 2 68938 50242
0 50244 5 1 1 50243
0 50245 7 1 2 50193 50244
0 50246 7 1 2 50071 50245
0 50247 5 1 1 50246
0 50248 7 1 2 59973 50247
0 50249 5 1 1 50248
0 50250 7 1 2 77932 73331
0 50251 5 3 1 50250
0 50252 7 1 2 89423 98122
0 50253 5 1 1 50252
0 50254 7 1 2 69597 50253
0 50255 5 1 1 50254
0 50256 7 1 2 87570 98123
0 50257 5 1 1 50256
0 50258 7 1 2 67748 50257
0 50259 5 1 1 50258
0 50260 7 1 2 50255 50259
0 50261 5 1 1 50260
0 50262 7 1 2 59663 50261
0 50263 5 1 1 50262
0 50264 7 1 2 82854 92831
0 50265 5 1 1 50264
0 50266 7 1 2 87571 50265
0 50267 5 1 1 50266
0 50268 7 1 2 60954 50267
0 50269 5 1 1 50268
0 50270 7 1 2 87613 95474
0 50271 5 1 1 50270
0 50272 7 1 2 50269 50271
0 50273 5 1 1 50272
0 50274 7 1 2 67749 50273
0 50275 5 1 1 50274
0 50276 7 1 2 50263 50275
0 50277 5 2 1 50276
0 50278 7 1 2 97814 98125
0 50279 5 1 1 50278
0 50280 7 2 2 68531 95446
0 50281 5 2 1 98127
0 50282 7 1 2 85852 98128
0 50283 5 1 1 50282
0 50284 7 1 2 50279 50283
0 50285 5 1 1 50284
0 50286 7 1 2 68781 50285
0 50287 5 1 1 50286
0 50288 7 1 2 76873 95393
0 50289 5 1 1 50288
0 50290 7 1 2 68532 50289
0 50291 5 1 1 50290
0 50292 7 1 2 66078 50291
0 50293 5 1 1 50292
0 50294 7 1 2 98092 50293
0 50295 5 1 1 50294
0 50296 7 1 2 50287 50295
0 50297 5 1 1 50296
0 50298 7 1 2 60721 50297
0 50299 5 1 1 50298
0 50300 7 1 2 80889 96574
0 50301 7 1 2 98126 50300
0 50302 5 1 1 50301
0 50303 7 1 2 50299 50302
0 50304 5 1 1 50303
0 50305 7 1 2 64147 50304
0 50306 5 1 1 50305
0 50307 7 1 2 96102 50085
0 50308 5 1 1 50307
0 50309 7 1 2 69207 89032
0 50310 5 1 1 50309
0 50311 7 1 2 68138 91596
0 50312 5 1 1 50311
0 50313 7 1 2 50310 50312
0 50314 5 2 1 50313
0 50315 7 1 2 76275 98131
0 50316 5 1 1 50315
0 50317 7 2 2 68139 91580
0 50318 7 1 2 76414 98133
0 50319 5 1 1 50318
0 50320 7 1 2 50316 50319
0 50321 5 1 1 50320
0 50322 7 1 2 78784 50321
0 50323 5 1 1 50322
0 50324 7 1 2 89698 50323
0 50325 5 1 1 50324
0 50326 7 1 2 79677 50325
0 50327 5 1 1 50326
0 50328 7 1 2 85295 50327
0 50329 7 1 2 50308 50328
0 50330 5 1 1 50329
0 50331 7 1 2 97403 50330
0 50332 5 1 1 50331
0 50333 7 1 2 50306 50332
0 50334 5 1 1 50333
0 50335 7 1 2 70694 50334
0 50336 5 1 1 50335
0 50337 7 1 2 96267 97939
0 50338 5 2 1 50337
0 50339 7 1 2 69598 98135
0 50340 5 1 1 50339
0 50341 7 1 2 12314 50340
0 50342 5 1 1 50341
0 50343 7 1 2 59664 50342
0 50344 5 1 1 50343
0 50345 7 1 2 78162 89816
0 50346 5 2 1 50345
0 50347 7 1 2 89957 98137
0 50348 7 1 2 50344 50347
0 50349 5 1 1 50348
0 50350 7 1 2 68140 50349
0 50351 5 1 1 50350
0 50352 7 1 2 68782 87551
0 50353 5 1 1 50352
0 50354 7 1 2 68533 93794
0 50355 7 1 2 50353 50354
0 50356 5 1 1 50355
0 50357 7 1 2 50351 50356
0 50358 5 1 1 50357
0 50359 7 1 2 97404 50358
0 50360 5 1 1 50359
0 50361 7 1 2 73351 84882
0 50362 5 1 1 50361
0 50363 7 1 2 97614 50362
0 50364 5 1 1 50363
0 50365 7 1 2 50360 50364
0 50366 5 1 1 50365
0 50367 7 1 2 60618 50366
0 50368 5 1 1 50367
0 50369 7 1 2 73323 98110
0 50370 5 1 1 50369
0 50371 7 3 2 86764 94744
0 50372 5 1 1 98139
0 50373 7 1 2 69599 98140
0 50374 5 1 1 50373
0 50375 7 1 2 50370 50374
0 50376 5 1 1 50375
0 50377 7 1 2 67389 50376
0 50378 5 1 1 50377
0 50379 7 4 2 64148 97389
0 50380 7 1 2 61929 18156
0 50381 7 1 2 98142 50380
0 50382 7 1 2 98129 50381
0 50383 5 1 1 50382
0 50384 7 1 2 50378 50383
0 50385 5 1 1 50384
0 50386 7 1 2 79678 50385
0 50387 5 1 1 50386
0 50388 7 1 2 69208 50169
0 50389 5 1 1 50388
0 50390 7 1 2 98106 50389
0 50391 5 1 1 50390
0 50392 7 1 2 61129 50391
0 50393 5 1 1 50392
0 50394 7 1 2 50387 50393
0 50395 7 1 2 50368 50394
0 50396 7 1 2 50336 50395
0 50397 5 1 1 50396
0 50398 7 1 2 64052 50397
0 50399 5 1 1 50398
0 50400 7 1 2 66079 69332
0 50401 5 1 1 50400
0 50402 7 1 2 76276 50401
0 50403 5 1 1 50402
0 50404 7 1 2 76415 91581
0 50405 5 1 1 50404
0 50406 7 1 2 63199 50405
0 50407 7 1 2 50403 50406
0 50408 5 1 1 50407
0 50409 7 1 2 76447 91366
0 50410 7 1 2 95626 50409
0 50411 5 1 1 50410
0 50412 7 1 2 65630 50411
0 50413 5 1 1 50412
0 50414 7 1 2 63582 50413
0 50415 7 1 2 50408 50414
0 50416 5 1 1 50415
0 50417 7 1 2 76652 90513
0 50418 7 1 2 94875 50417
0 50419 7 1 2 74189 50418
0 50420 5 1 1 50419
0 50421 7 1 2 50416 50420
0 50422 5 1 1 50421
0 50423 7 1 2 66766 50422
0 50424 5 1 1 50423
0 50425 7 1 2 80821 91557
0 50426 7 2 2 70695 92776
0 50427 7 1 2 69710 89001
0 50428 5 1 1 50427
0 50429 7 1 2 98146 50428
0 50430 7 1 2 50425 50429
0 50431 5 1 1 50430
0 50432 7 1 2 50424 50431
0 50433 5 1 1 50432
0 50434 7 1 2 61930 50433
0 50435 5 1 1 50434
0 50436 7 1 2 84807 86485
0 50437 7 1 2 76317 50436
0 50438 7 1 2 98116 50437
0 50439 5 1 1 50438
0 50440 7 1 2 50435 50439
0 50441 5 1 1 50440
0 50442 7 1 2 63846 50441
0 50443 5 1 1 50442
0 50444 7 1 2 96138 98147
0 50445 7 1 2 97989 50444
0 50446 5 1 1 50445
0 50447 7 1 2 50443 50446
0 50448 5 1 1 50447
0 50449 7 1 2 64149 50448
0 50450 5 1 1 50449
0 50451 7 1 2 70696 97991
0 50452 5 1 1 50451
0 50453 7 1 2 65513 50452
0 50454 5 1 1 50453
0 50455 7 1 2 84883 86726
0 50456 7 2 2 97655 50455
0 50457 5 1 1 98148
0 50458 7 1 2 50454 98149
0 50459 5 1 1 50458
0 50460 7 1 2 88021 97660
0 50461 5 1 1 50460
0 50462 7 1 2 74102 96509
0 50463 5 1 1 50462
0 50464 7 1 2 59665 97371
0 50465 5 1 1 50464
0 50466 7 1 2 50463 50465
0 50467 5 1 1 50466
0 50468 7 1 2 69600 50467
0 50469 5 1 1 50468
0 50470 7 1 2 63200 74668
0 50471 5 1 1 50470
0 50472 7 1 2 96510 50471
0 50473 5 1 1 50472
0 50474 7 1 2 50469 50473
0 50475 5 1 1 50474
0 50476 7 1 2 64150 92008
0 50477 7 1 2 50475 50476
0 50478 5 1 1 50477
0 50479 7 1 2 50461 50478
0 50480 5 1 1 50479
0 50481 7 1 2 94351 50480
0 50482 5 1 1 50481
0 50483 7 1 2 73955 97926
0 50484 7 1 2 97680 50483
0 50485 5 1 1 50484
0 50486 7 1 2 50482 50485
0 50487 5 1 1 50486
0 50488 7 1 2 85793 50487
0 50489 5 1 1 50488
0 50490 7 1 2 50459 50489
0 50491 7 1 2 50450 50490
0 50492 5 1 1 50491
0 50493 7 1 2 68939 50492
0 50494 5 1 1 50493
0 50495 7 2 2 59666 92447
0 50496 5 1 1 98150
0 50497 7 1 2 96268 50496
0 50498 5 1 1 50497
0 50499 7 1 2 97670 50498
0 50500 5 1 1 50499
0 50501 7 1 2 75444 76448
0 50502 7 1 2 98058 50501
0 50503 5 1 1 50502
0 50504 7 1 2 50014 50503
0 50505 5 1 1 50504
0 50506 7 1 2 70697 50505
0 50507 5 1 1 50506
0 50508 7 1 2 97647 98052
0 50509 5 1 1 50508
0 50510 7 1 2 97020 98112
0 50511 5 1 1 50510
0 50512 7 1 2 50509 50511
0 50513 5 1 1 50512
0 50514 7 1 2 76277 50513
0 50515 5 1 1 50514
0 50516 7 1 2 50042 50515
0 50517 7 1 2 50507 50516
0 50518 5 1 1 50517
0 50519 7 1 2 67750 50518
0 50520 5 1 1 50519
0 50521 7 1 2 50500 50520
0 50522 5 1 1 50521
0 50523 7 1 2 68141 50522
0 50524 5 1 1 50523
0 50525 7 1 2 81597 77486
0 50526 7 1 2 93170 50525
0 50527 7 1 2 97815 50526
0 50528 5 1 1 50527
0 50529 7 1 2 63583 96188
0 50530 5 1 1 50529
0 50531 7 1 2 50528 50530
0 50532 5 1 1 50531
0 50533 7 1 2 60722 50532
0 50534 5 1 1 50533
0 50535 7 2 2 68534 73361
0 50536 5 1 1 98152
0 50537 7 1 2 97785 98153
0 50538 7 1 2 98120 50537
0 50539 5 1 1 50538
0 50540 7 1 2 50534 50539
0 50541 5 1 1 50540
0 50542 7 1 2 94720 50541
0 50543 5 1 1 50542
0 50544 7 2 2 76427 93040
0 50545 7 2 2 67751 94218
0 50546 7 1 2 92574 98156
0 50547 7 1 2 98154 50546
0 50548 5 1 1 50547
0 50549 7 1 2 50543 50548
0 50550 7 1 2 50524 50549
0 50551 5 1 1 50550
0 50552 7 1 2 64053 50551
0 50553 5 1 1 50552
0 50554 7 1 2 97950 97956
0 50555 5 1 1 50554
0 50556 7 1 2 69601 50555
0 50557 5 1 1 50556
0 50558 7 1 2 74974 97952
0 50559 5 1 1 50558
0 50560 7 1 2 50557 50559
0 50561 5 1 1 50560
0 50562 7 1 2 74103 50561
0 50563 5 1 1 50562
0 50564 7 1 2 59667 76192
0 50565 7 1 2 94229 50564
0 50566 5 1 1 50565
0 50567 7 1 2 97957 50566
0 50568 5 1 1 50567
0 50569 7 1 2 68142 50568
0 50570 5 1 1 50569
0 50571 7 1 2 50563 50570
0 50572 5 1 1 50571
0 50573 7 1 2 66767 50572
0 50574 5 1 1 50573
0 50575 7 1 2 78785 74975
0 50576 5 1 1 50575
0 50577 7 1 2 84851 50576
0 50578 5 1 1 50577
0 50579 7 1 2 69602 50578
0 50580 5 1 1 50579
0 50581 7 1 2 65514 83513
0 50582 5 1 1 50581
0 50583 7 1 2 63847 50582
0 50584 5 1 1 50583
0 50585 7 2 2 83568 91624
0 50586 5 1 1 98158
0 50587 7 1 2 50584 50586
0 50588 5 1 1 50587
0 50589 7 1 2 67752 50588
0 50590 5 1 1 50589
0 50591 7 1 2 50580 50590
0 50592 5 1 1 50591
0 50593 7 1 2 61795 50592
0 50594 5 1 1 50593
0 50595 7 1 2 76278 91165
0 50596 5 1 1 50595
0 50597 7 1 2 83221 50596
0 50598 5 1 1 50597
0 50599 7 1 2 91764 50598
0 50600 5 1 1 50599
0 50601 7 1 2 50594 50600
0 50602 5 1 1 50601
0 50603 7 1 2 94767 50602
0 50604 5 1 1 50603
0 50605 7 1 2 50574 50604
0 50606 5 1 1 50605
0 50607 7 1 2 86804 50606
0 50608 5 1 1 50607
0 50609 7 1 2 50553 50608
0 50610 5 1 1 50609
0 50611 7 1 2 85794 50610
0 50612 5 1 1 50611
0 50613 7 1 2 50494 50612
0 50614 7 1 2 50399 50613
0 50615 7 1 2 50249 50614
0 50616 7 1 2 49775 50615
0 50617 5 1 1 50616
0 50618 7 1 2 95302 50617
0 50619 5 1 1 50618
0 50620 7 2 2 90238 88706
0 50621 7 1 2 69603 98160
0 50622 5 1 1 50621
0 50623 7 1 2 92210 50622
0 50624 5 1 1 50623
0 50625 7 1 2 60955 50624
0 50626 5 1 1 50625
0 50627 7 1 2 49629 50626
0 50628 5 1 1 50627
0 50629 7 1 2 59974 50628
0 50630 5 1 1 50629
0 50631 7 1 2 71898 88755
0 50632 5 1 1 50631
0 50633 7 1 2 50630 50632
0 50634 5 1 1 50633
0 50635 7 2 2 67390 97699
0 50636 7 1 2 95332 98121
0 50637 7 1 2 98162 50636
0 50638 7 1 2 50634 50637
0 50639 5 1 1 50638
0 50640 7 1 2 50619 50639
0 50641 5 1 1 50640
0 50642 7 1 2 75354 50641
0 50643 5 1 1 50642
0 50644 7 3 2 83569 94178
0 50645 7 1 2 59975 98164
0 50646 5 1 1 50645
0 50647 7 1 2 67125 91813
0 50648 5 1 1 50647
0 50649 7 1 2 50646 50648
0 50650 5 1 1 50649
0 50651 7 1 2 61931 50650
0 50652 5 1 1 50651
0 50653 7 1 2 92700 92492
0 50654 5 1 1 50653
0 50655 7 1 2 50652 50654
0 50656 5 1 1 50655
0 50657 7 1 2 60723 50656
0 50658 5 1 1 50657
0 50659 7 1 2 96202 98013
0 50660 5 1 1 50659
0 50661 7 1 2 50658 50660
0 50662 5 1 1 50661
0 50663 7 1 2 98005 50662
0 50664 5 1 1 50663
0 50665 7 4 2 64151 97578
0 50666 7 2 2 86496 98167
0 50667 7 1 2 61130 98171
0 50668 5 1 1 50667
0 50669 7 1 2 50664 50668
0 50670 5 1 1 50669
0 50671 7 1 2 59668 50670
0 50672 5 1 1 50671
0 50673 7 3 2 96706 97585
0 50674 5 2 1 98173
0 50675 7 1 2 85539 92866
0 50676 7 1 2 98174 50675
0 50677 5 1 1 50676
0 50678 7 1 2 50672 50677
0 50679 5 1 1 50678
0 50680 7 1 2 68143 50679
0 50681 5 1 1 50680
0 50682 7 1 2 82656 87876
0 50683 5 1 1 50682
0 50684 7 4 2 61131 79268
0 50685 7 1 2 87922 98178
0 50686 5 1 1 50685
0 50687 7 1 2 79638 96232
0 50688 5 1 1 50687
0 50689 7 1 2 50686 50688
0 50690 5 1 1 50689
0 50691 7 1 2 59976 50690
0 50692 5 1 1 50691
0 50693 7 1 2 39877 97382
0 50694 5 1 1 50693
0 50695 7 1 2 84385 50694
0 50696 5 1 1 50695
0 50697 7 1 2 79894 87867
0 50698 7 1 2 96479 50697
0 50699 5 1 1 50698
0 50700 7 1 2 50696 50699
0 50701 7 1 2 50692 50700
0 50702 5 1 1 50701
0 50703 7 1 2 66903 50702
0 50704 5 1 1 50703
0 50705 7 1 2 50683 50704
0 50706 5 1 1 50705
0 50707 7 1 2 59669 50706
0 50708 5 1 1 50707
0 50709 7 1 2 94082 96129
0 50710 5 1 1 50709
0 50711 7 1 2 50708 50710
0 50712 5 1 1 50711
0 50713 7 1 2 69017 50712
0 50714 5 1 1 50713
0 50715 7 1 2 61796 96628
0 50716 5 1 1 50715
0 50717 7 1 2 98009 50716
0 50718 5 1 1 50717
0 50719 7 1 2 90180 50718
0 50720 5 1 1 50719
0 50721 7 1 2 63201 96575
0 50722 7 1 2 98179 50721
0 50723 5 1 1 50722
0 50724 7 1 2 50720 50723
0 50725 5 1 1 50724
0 50726 7 1 2 94768 50725
0 50727 5 1 1 50726
0 50728 7 1 2 50714 50727
0 50729 5 1 1 50728
0 50730 7 1 2 65631 50729
0 50731 5 1 1 50730
0 50732 7 2 2 69018 94881
0 50733 7 1 2 96054 96269
0 50734 5 1 1 50733
0 50735 7 1 2 61132 50734
0 50736 5 1 1 50735
0 50737 7 1 2 98097 50736
0 50738 5 1 1 50737
0 50739 7 1 2 59670 50738
0 50740 5 1 1 50739
0 50741 7 1 2 96197 50740
0 50742 5 1 1 50741
0 50743 7 1 2 98182 50742
0 50744 5 1 1 50743
0 50745 7 1 2 84270 96577
0 50746 5 1 1 50745
0 50747 7 1 2 50744 50746
0 50748 5 1 1 50747
0 50749 7 1 2 65632 50748
0 50750 5 1 1 50749
0 50751 7 2 2 84271 85713
0 50752 7 1 2 95918 98184
0 50753 5 1 1 50752
0 50754 7 1 2 50750 50753
0 50755 5 1 1 50754
0 50756 7 1 2 91691 50755
0 50757 5 1 1 50756
0 50758 7 2 2 59671 91885
0 50759 7 1 2 96942 98186
0 50760 5 1 1 50759
0 50761 7 1 2 96604 50760
0 50762 5 1 1 50761
0 50763 7 2 2 63202 50762
0 50764 7 1 2 92867 98188
0 50765 5 1 1 50764
0 50766 7 1 2 96616 97448
0 50767 5 1 1 50766
0 50768 7 1 2 50765 50767
0 50769 5 1 1 50768
0 50770 7 1 2 66585 50769
0 50771 5 1 1 50770
0 50772 7 4 2 65515 94731
0 50773 5 1 1 98190
0 50774 7 1 2 94199 98191
0 50775 5 1 1 50774
0 50776 7 1 2 50771 50775
0 50777 5 1 1 50776
0 50778 7 1 2 60724 50777
0 50779 5 1 1 50778
0 50780 7 1 2 50757 50779
0 50781 7 1 2 50731 50780
0 50782 5 1 1 50781
0 50783 7 1 2 68535 50782
0 50784 5 1 1 50783
0 50785 7 5 2 64152 89325
0 50786 7 1 2 72254 97460
0 50787 7 1 2 86374 50786
0 50788 7 1 2 98194 50787
0 50789 5 1 1 50788
0 50790 7 1 2 50784 50789
0 50791 7 1 2 50681 50790
0 50792 5 1 1 50791
0 50793 7 1 2 67753 50792
0 50794 5 1 1 50793
0 50795 7 1 2 83206 92484
0 50796 5 1 1 50795
0 50797 7 1 2 96490 50796
0 50798 5 1 1 50797
0 50799 7 2 2 68536 95664
0 50800 5 2 1 98199
0 50801 7 1 2 67126 96878
0 50802 5 1 1 50801
0 50803 7 1 2 98201 50802
0 50804 5 1 1 50803
0 50805 7 1 2 61797 50804
0 50806 5 1 1 50805
0 50807 7 1 2 50798 50806
0 50808 5 1 1 50807
0 50809 7 1 2 97405 50808
0 50810 5 1 1 50809
0 50811 7 3 2 63584 98168
0 50812 7 1 2 82657 98203
0 50813 5 1 1 50812
0 50814 7 1 2 50810 50813
0 50815 5 1 1 50814
0 50816 7 1 2 68783 50815
0 50817 5 1 1 50816
0 50818 7 4 2 91814 98023
0 50819 7 1 2 59672 98206
0 50820 5 1 1 50819
0 50821 7 1 2 50817 50820
0 50822 5 1 1 50821
0 50823 7 1 2 59977 50822
0 50824 5 1 1 50823
0 50825 7 1 2 92302 97436
0 50826 5 3 1 50825
0 50827 7 2 2 82195 86861
0 50828 7 1 2 96924 98213
0 50829 5 1 1 50828
0 50830 7 1 2 98210 50829
0 50831 5 1 1 50830
0 50832 7 1 2 90181 50831
0 50833 5 1 1 50832
0 50834 7 1 2 95697 98214
0 50835 5 1 1 50834
0 50836 7 1 2 98015 98211
0 50837 5 1 1 50836
0 50838 7 1 2 96989 50837
0 50839 5 1 1 50838
0 50840 7 1 2 50835 50839
0 50841 7 1 2 50833 50840
0 50842 5 1 1 50841
0 50843 7 1 2 63848 50842
0 50844 5 1 1 50843
0 50845 7 2 2 92859 96733
0 50846 7 2 2 94636 98215
0 50847 5 1 1 98217
0 50848 7 1 2 61133 98218
0 50849 5 1 1 50848
0 50850 7 1 2 50844 50849
0 50851 5 1 1 50850
0 50852 7 1 2 59673 50851
0 50853 5 1 1 50852
0 50854 7 1 2 50824 50853
0 50855 5 1 1 50854
0 50856 7 1 2 68144 50855
0 50857 5 1 1 50856
0 50858 7 1 2 59674 97924
0 50859 5 1 1 50858
0 50860 7 1 2 89817 96913
0 50861 7 1 2 97479 50860
0 50862 5 1 1 50861
0 50863 7 1 2 50859 50862
0 50864 5 1 1 50863
0 50865 7 1 2 91692 50864
0 50866 5 1 1 50865
0 50867 7 4 2 64153 90207
0 50868 7 1 2 83191 86260
0 50869 7 1 2 98219 50868
0 50870 5 1 1 50869
0 50871 7 1 2 75717 87080
0 50872 7 1 2 83324 50871
0 50873 7 1 2 96580 50872
0 50874 5 1 1 50873
0 50875 7 1 2 50870 50874
0 50876 5 1 1 50875
0 50877 7 1 2 97796 50876
0 50878 5 1 1 50877
0 50879 7 1 2 75527 97461
0 50880 7 1 2 87929 50879
0 50881 7 1 2 96905 50880
0 50882 5 1 1 50881
0 50883 7 1 2 96617 98001
0 50884 7 1 2 97480 50883
0 50885 5 1 1 50884
0 50886 7 1 2 50882 50885
0 50887 7 1 2 50878 50886
0 50888 5 1 1 50887
0 50889 7 1 2 63203 50888
0 50890 5 1 1 50889
0 50891 7 1 2 50866 50890
0 50892 7 1 2 50857 50891
0 50893 5 1 1 50892
0 50894 7 1 2 64054 50893
0 50895 5 1 1 50894
0 50896 7 2 2 92274 92524
0 50897 5 1 1 98223
0 50898 7 1 2 97383 50897
0 50899 5 1 1 50898
0 50900 7 1 2 96879 50899
0 50901 5 1 1 50900
0 50902 7 2 2 64055 91693
0 50903 7 1 2 84367 92481
0 50904 7 1 2 98225 50903
0 50905 5 1 1 50904
0 50906 7 1 2 50901 50905
0 50907 5 1 1 50906
0 50908 7 1 2 68145 50907
0 50909 5 1 1 50908
0 50910 7 1 2 91472 92249
0 50911 5 1 1 50910
0 50912 7 1 2 50909 50911
0 50913 5 1 1 50912
0 50914 7 1 2 69019 50913
0 50915 5 1 1 50914
0 50916 7 2 2 82002 96679
0 50917 5 1 1 98227
0 50918 7 1 2 96203 98228
0 50919 5 1 1 50918
0 50920 7 1 2 50915 50919
0 50921 5 1 1 50920
0 50922 7 1 2 65633 50921
0 50923 5 1 1 50922
0 50924 7 1 2 73486 89818
0 50925 7 1 2 95997 50924
0 50926 5 1 1 50925
0 50927 7 1 2 3188 50926
0 50928 5 1 1 50927
0 50929 7 1 2 91694 50928
0 50930 5 2 1 50929
0 50931 7 1 2 92124 90059
0 50932 7 1 2 96655 50931
0 50933 5 1 1 50932
0 50934 7 1 2 98229 50933
0 50935 5 1 1 50934
0 50936 7 1 2 94721 50935
0 50937 5 1 1 50936
0 50938 7 1 2 66586 98189
0 50939 5 1 1 50938
0 50940 7 1 2 50937 50939
0 50941 5 1 1 50940
0 50942 7 1 2 59978 50941
0 50943 5 1 1 50942
0 50944 7 1 2 96092 98195
0 50945 5 1 1 50944
0 50946 7 1 2 50943 50945
0 50947 5 1 1 50946
0 50948 7 1 2 97424 50947
0 50949 5 1 1 50948
0 50950 7 1 2 50923 50949
0 50951 5 1 1 50950
0 50952 7 1 2 66904 50951
0 50953 5 1 1 50952
0 50954 7 1 2 68940 86884
0 50955 5 1 1 50954
0 50956 7 1 2 98230 50955
0 50957 5 1 1 50956
0 50958 7 1 2 94722 50957
0 50959 5 1 1 50958
0 50960 7 1 2 79490 94608
0 50961 7 1 2 98187 50960
0 50962 5 1 1 50961
0 50963 7 1 2 50959 50962
0 50964 5 1 1 50963
0 50965 7 1 2 65634 50964
0 50966 5 1 1 50965
0 50967 7 2 2 91695 97372
0 50968 5 1 1 98231
0 50969 7 1 2 97498 97797
0 50970 5 1 1 50969
0 50971 7 1 2 50968 50970
0 50972 5 1 1 50971
0 50973 7 1 2 73487 97469
0 50974 7 1 2 50972 50973
0 50975 5 1 1 50974
0 50976 7 1 2 50966 50975
0 50977 5 1 1 50976
0 50978 7 1 2 59979 50977
0 50979 5 1 1 50978
0 50980 7 3 2 91696 94769
0 50981 7 1 2 65635 96264
0 50982 7 1 2 98233 50981
0 50983 5 1 1 50982
0 50984 7 1 2 50979 50983
0 50985 5 1 1 50984
0 50986 7 1 2 61932 50985
0 50987 5 1 1 50986
0 50988 7 1 2 74685 87868
0 50989 7 1 2 95744 50988
0 50990 7 1 2 91425 95748
0 50991 7 1 2 50989 50990
0 50992 5 1 1 50991
0 50993 7 1 2 50987 50992
0 50994 5 1 1 50993
0 50995 7 1 2 68537 50994
0 50996 5 1 1 50995
0 50997 7 1 2 50953 50996
0 50998 5 1 1 50997
0 50999 7 1 2 73828 50998
0 51000 5 1 1 50999
0 51001 7 2 2 89694 97601
0 51002 7 1 2 88628 96780
0 51003 7 1 2 98236 51002
0 51004 5 1 1 51003
0 51005 7 2 2 87191 91697
0 51006 7 1 2 72482 98159
0 51007 5 1 1 51006
0 51008 7 1 2 76566 95093
0 51009 5 1 1 51008
0 51010 7 1 2 51007 51009
0 51011 5 1 1 51010
0 51012 7 1 2 98238 51011
0 51013 5 1 1 51012
0 51014 7 2 2 92345 92754
0 51015 7 1 2 89976 92571
0 51016 7 1 2 98240 51015
0 51017 5 1 1 51016
0 51018 7 1 2 51013 51017
0 51019 7 1 2 51004 51018
0 51020 5 1 1 51019
0 51021 7 1 2 64154 51020
0 51022 5 1 1 51021
0 51023 7 1 2 87542 95804
0 51024 7 1 2 91752 51023
0 51025 7 1 2 96958 51024
0 51026 5 1 1 51025
0 51027 7 1 2 51022 51026
0 51028 5 1 1 51027
0 51029 7 1 2 68941 51028
0 51030 5 1 1 51029
0 51031 7 1 2 51000 51030
0 51032 7 1 2 50895 51031
0 51033 7 1 2 50794 51032
0 51034 5 1 1 51033
0 51035 7 1 2 95303 51034
0 51036 5 1 1 51035
0 51037 7 2 2 68538 69020
0 51038 7 1 2 95335 98242
0 51039 5 1 1 51038
0 51040 7 5 2 64155 95304
0 51041 7 1 2 66905 83112
0 51042 7 1 2 98244 51041
0 51043 5 1 1 51042
0 51044 7 1 2 69021 84808
0 51045 7 1 2 95336 51044
0 51046 5 1 1 51045
0 51047 7 1 2 51043 51046
0 51048 5 1 1 51047
0 51049 7 1 2 75028 51048
0 51050 5 1 1 51049
0 51051 7 1 2 51039 51050
0 51052 5 1 1 51051
0 51053 7 1 2 68784 51052
0 51054 5 1 1 51053
0 51055 7 1 2 72255 93982
0 51056 7 1 2 95305 51055
0 51057 7 1 2 97934 51056
0 51058 5 1 1 51057
0 51059 7 1 2 51054 51058
0 51060 5 1 1 51059
0 51061 7 1 2 61798 51060
0 51062 5 1 1 51061
0 51063 7 1 2 98245 98050
0 51064 5 1 1 51063
0 51065 7 1 2 51062 51064
0 51066 5 1 1 51065
0 51067 7 1 2 60619 51066
0 51068 5 1 1 51067
0 51069 7 1 2 72256 89715
0 51070 5 1 1 51069
0 51071 7 1 2 97594 51070
0 51072 5 1 1 51071
0 51073 7 1 2 59675 51072
0 51074 5 1 1 51073
0 51075 7 1 2 84557 51074
0 51076 5 1 1 51075
0 51077 7 1 2 95306 97739
0 51078 7 1 2 51076 51077
0 51079 5 1 1 51078
0 51080 7 1 2 51068 51079
0 51081 5 1 1 51080
0 51082 7 1 2 75528 51081
0 51083 5 1 1 51082
0 51084 7 2 2 68146 69022
0 51085 7 1 2 92868 94782
0 51086 7 1 2 98249 51085
0 51087 5 1 1 51086
0 51088 7 1 2 98031 51087
0 51089 5 1 1 51088
0 51090 7 1 2 85684 51089
0 51091 5 1 1 51090
0 51092 7 1 2 88649 97972
0 51093 5 1 1 51092
0 51094 7 1 2 80910 51093
0 51095 5 1 1 51094
0 51096 7 1 2 97740 51095
0 51097 5 1 1 51096
0 51098 7 1 2 51091 51097
0 51099 5 1 1 51098
0 51100 7 1 2 63849 51099
0 51101 5 1 1 51100
0 51102 7 1 2 97592 97874
0 51103 7 1 2 87495 51102
0 51104 5 1 1 51103
0 51105 7 1 2 51101 51104
0 51106 5 1 1 51105
0 51107 7 1 2 95307 51106
0 51108 5 1 1 51107
0 51109 7 1 2 51083 51108
0 51110 5 1 1 51109
0 51111 7 1 2 68942 51110
0 51112 5 1 1 51111
0 51113 7 1 2 87625 88120
0 51114 5 1 1 51113
0 51115 7 2 2 94939 51114
0 51116 5 1 1 98251
0 51117 7 1 2 63204 92499
0 51118 5 1 1 51117
0 51119 7 1 2 87634 51118
0 51120 5 1 1 51119
0 51121 7 1 2 75529 51120
0 51122 5 1 1 51121
0 51123 7 1 2 98252 51122
0 51124 5 2 1 51123
0 51125 7 1 2 66906 98253
0 51126 5 1 1 51125
0 51127 7 1 2 85853 94072
0 51128 5 1 1 51127
0 51129 7 1 2 51126 51128
0 51130 5 1 1 51129
0 51131 7 1 2 71242 94219
0 51132 7 1 2 51130 51131
0 51133 5 1 1 51132
0 51134 7 1 2 97629 97897
0 51135 5 1 1 51134
0 51136 7 1 2 96995 51135
0 51137 5 1 1 51136
0 51138 7 1 2 82658 96672
0 51139 7 1 2 51137 51138
0 51140 5 1 1 51139
0 51141 7 1 2 51133 51140
0 51142 5 1 1 51141
0 51143 7 1 2 59676 51142
0 51144 5 1 1 51143
0 51145 7 1 2 78786 84809
0 51146 7 1 2 98169 51145
0 51147 5 1 1 51146
0 51148 7 1 2 51144 51147
0 51149 5 1 1 51148
0 51150 7 1 2 97764 51149
0 51151 5 1 1 51150
0 51152 7 1 2 51112 51151
0 51153 5 1 1 51152
0 51154 7 1 2 95932 51153
0 51155 5 1 1 51154
0 51156 7 2 2 68943 69023
0 51157 7 2 2 68785 98255
0 51158 7 1 2 81498 95254
0 51159 7 2 2 98257 51158
0 51160 7 1 2 61371 95261
0 51161 7 2 2 98259 51160
0 51162 7 1 2 73829 78134
0 51163 7 1 2 89297 51162
0 51164 7 1 2 98261 51163
0 51165 5 1 1 51164
0 51166 7 1 2 51155 51165
0 51167 7 1 2 51036 51166
0 51168 5 1 1 51167
0 51169 7 1 2 69962 51168
0 51170 5 1 1 51169
0 51171 7 2 2 90128 95333
0 51172 7 1 2 81499 98263
0 51173 7 3 2 97696 51172
0 51174 7 1 2 78149 50127
0 51175 5 2 1 51174
0 51176 7 1 2 98265 98268
0 51177 5 1 1 51176
0 51178 7 1 2 91483 98165
0 51179 5 1 1 51178
0 51180 7 1 2 19784 51179
0 51181 5 1 1 51180
0 51182 7 1 2 59677 51181
0 51183 5 1 1 51182
0 51184 7 3 2 75355 80961
0 51185 5 1 1 98270
0 51186 7 1 2 89839 51185
0 51187 5 1 1 51186
0 51188 7 1 2 79679 51187
0 51189 5 1 1 51188
0 51190 7 1 2 49667 51189
0 51191 5 1 1 51190
0 51192 7 1 2 63850 51191
0 51193 5 1 1 51192
0 51194 7 1 2 51183 51193
0 51195 5 1 1 51194
0 51196 7 1 2 60725 51195
0 51197 5 1 1 51196
0 51198 7 1 2 92151 89658
0 51199 7 1 2 98155 51198
0 51200 5 1 1 51199
0 51201 7 1 2 51197 51200
0 51202 5 1 1 51201
0 51203 7 1 2 66907 51202
0 51204 5 1 1 51203
0 51205 7 1 2 73362 96199
0 51206 7 1 2 97798 51205
0 51207 5 1 1 51206
0 51208 7 1 2 51204 51207
0 51209 5 1 1 51208
0 51210 7 1 2 68147 51209
0 51211 5 1 1 51210
0 51212 7 1 2 86407 97799
0 51213 5 1 1 51212
0 51214 7 1 2 39412 51213
0 51215 5 1 1 51214
0 51216 7 1 2 73458 78163
0 51217 7 1 2 51215 51216
0 51218 5 1 1 51217
0 51219 7 1 2 51211 51218
0 51220 5 1 1 51219
0 51221 7 1 2 68944 51220
0 51222 5 1 1 51221
0 51223 7 1 2 76449 91833
0 51224 5 1 1 51223
0 51225 7 1 2 96608 51224
0 51226 5 1 1 51225
0 51227 7 1 2 61933 51226
0 51228 5 1 1 51227
0 51229 7 1 2 61799 97867
0 51230 5 1 1 51229
0 51231 7 1 2 51228 51230
0 51232 5 1 1 51231
0 51233 7 1 2 75388 51232
0 51234 5 1 1 51233
0 51235 7 2 2 67754 91815
0 51236 5 1 1 98273
0 51237 7 1 2 61934 98274
0 51238 5 1 1 51237
0 51239 7 1 2 51234 51238
0 51240 5 1 1 51239
0 51241 7 1 2 85883 51240
0 51242 5 1 1 51241
0 51243 7 1 2 51222 51242
0 51244 5 1 1 51243
0 51245 7 1 2 64156 51244
0 51246 5 1 1 51245
0 51247 7 1 2 85780 92826
0 51248 5 1 1 51247
0 51249 7 1 2 92803 51248
0 51250 5 1 1 51249
0 51251 7 1 2 79491 51250
0 51252 5 1 1 51251
0 51253 7 1 2 91698 97942
0 51254 5 1 1 51253
0 51255 7 1 2 76450 88016
0 51256 7 1 2 94160 51255
0 51257 5 1 1 51256
0 51258 7 1 2 36879 51257
0 51259 5 1 1 51258
0 51260 7 1 2 63851 51259
0 51261 5 1 1 51260
0 51262 7 1 2 51254 51261
0 51263 5 1 1 51262
0 51264 7 1 2 66908 51263
0 51265 5 1 1 51264
0 51266 7 1 2 51252 51265
0 51267 5 1 1 51266
0 51268 7 1 2 68539 51267
0 51269 5 1 1 51268
0 51270 7 2 2 89494 14531
0 51271 5 2 1 98275
0 51272 7 2 2 66909 79024
0 51273 7 1 2 94409 98279
0 51274 7 1 2 98277 51273
0 51275 5 1 1 51274
0 51276 7 1 2 51269 51275
0 51277 5 1 1 51276
0 51278 7 1 2 69024 51277
0 51279 5 1 1 51278
0 51280 7 3 2 64157 89943
0 51281 7 2 2 89454 98281
0 51282 5 1 1 98284
0 51283 7 2 2 87295 98285
0 51284 5 1 1 98286
0 51285 7 1 2 64056 51284
0 51286 7 1 2 51279 51285
0 51287 5 1 1 51286
0 51288 7 2 2 66910 97857
0 51289 7 2 2 93859 98288
0 51290 5 1 1 98290
0 51291 7 1 2 76451 98291
0 51292 5 1 1 51291
0 51293 7 4 2 64158 79680
0 51294 7 1 2 80962 87296
0 51295 7 1 2 98292 51294
0 51296 5 1 1 51295
0 51297 7 1 2 51292 51296
0 51298 5 1 1 51297
0 51299 7 1 2 75356 51298
0 51300 5 1 1 51299
0 51301 7 1 2 91699 97889
0 51302 7 1 2 98269 51301
0 51303 5 1 1 51302
0 51304 7 1 2 51300 51303
0 51305 5 1 1 51304
0 51306 7 1 2 63852 51305
0 51307 5 1 1 51306
0 51308 7 3 2 61935 94179
0 51309 7 1 2 75695 94723
0 51310 7 1 2 96667 51309
0 51311 7 1 2 98296 51310
0 51312 5 1 1 51311
0 51313 7 1 2 68945 51312
0 51314 7 1 2 51307 51313
0 51315 5 1 1 51314
0 51316 7 1 2 65636 51315
0 51317 7 1 2 51287 51316
0 51318 5 1 1 51317
0 51319 7 2 2 77802 94609
0 51320 7 1 2 97719 98299
0 51321 5 1 1 51320
0 51322 7 4 2 64159 97899
0 51323 7 2 2 61800 98301
0 51324 5 1 1 98305
0 51325 7 1 2 91700 95634
0 51326 5 1 1 51325
0 51327 7 1 2 51324 51326
0 51328 5 2 1 51327
0 51329 7 1 2 92763 98307
0 51330 5 1 1 51329
0 51331 7 1 2 97406 97961
0 51332 5 1 1 51331
0 51333 7 1 2 95635 96265
0 51334 5 1 1 51333
0 51335 7 1 2 51332 51334
0 51336 5 1 1 51335
0 51337 7 1 2 91701 51336
0 51338 5 1 1 51337
0 51339 7 2 2 79492 87927
0 51340 5 1 1 98309
0 51341 7 1 2 97618 98310
0 51342 5 1 1 51341
0 51343 7 1 2 48298 51342
0 51344 5 1 1 51343
0 51345 7 1 2 67127 51344
0 51346 5 1 1 51345
0 51347 7 1 2 51338 51346
0 51348 7 1 2 51330 51347
0 51349 5 1 1 51348
0 51350 7 1 2 64057 51349
0 51351 5 1 1 51350
0 51352 7 2 2 75357 87192
0 51353 7 1 2 97851 97940
0 51354 5 1 1 51353
0 51355 7 1 2 98311 51354
0 51356 5 1 1 51355
0 51357 7 1 2 67755 87643
0 51358 7 1 2 92233 51357
0 51359 5 1 1 51358
0 51360 7 1 2 51356 51359
0 51361 5 1 1 51360
0 51362 7 1 2 97733 51361
0 51363 5 1 1 51362
0 51364 7 1 2 67756 94741
0 51365 5 1 1 51364
0 51366 7 1 2 51363 51365
0 51367 5 1 1 51366
0 51368 7 1 2 80984 51367
0 51369 5 1 1 51368
0 51370 7 1 2 51351 51369
0 51371 5 1 1 51370
0 51372 7 1 2 76279 51371
0 51373 5 1 1 51372
0 51374 7 1 2 51321 51373
0 51375 7 1 2 51318 51374
0 51376 7 1 2 51246 51375
0 51377 5 1 1 51376
0 51378 7 1 2 95308 51377
0 51379 5 1 1 51378
0 51380 7 1 2 51177 51379
0 51381 5 1 1 51380
0 51382 7 1 2 71243 51381
0 51383 5 1 1 51382
0 51384 7 1 2 59678 75389
0 51385 5 2 1 51384
0 51386 7 1 2 91661 98313
0 51387 5 2 1 51386
0 51388 7 1 2 77583 98315
0 51389 5 1 1 51388
0 51390 7 1 2 75029 93940
0 51391 5 1 1 51390
0 51392 7 1 2 51389 51391
0 51393 5 1 1 51392
0 51394 7 1 2 66768 51393
0 51395 5 1 1 51394
0 51396 7 1 2 22557 51395
0 51397 5 1 1 51396
0 51398 7 1 2 97407 51397
0 51399 5 1 1 51398
0 51400 7 1 2 75358 96189
0 51401 5 2 1 51400
0 51402 7 1 2 40313 97818
0 51403 5 3 1 51402
0 51404 7 1 2 75120 98319
0 51405 5 1 1 51404
0 51406 7 1 2 98317 51405
0 51407 5 1 1 51406
0 51408 7 1 2 60726 51407
0 51409 5 1 1 51408
0 51410 7 1 2 86326 89819
0 51411 7 1 2 95512 51410
0 51412 5 1 1 51411
0 51413 7 1 2 51409 51412
0 51414 5 1 1 51413
0 51415 7 1 2 87869 97875
0 51416 7 1 2 51414 51415
0 51417 5 1 1 51416
0 51418 7 1 2 51399 51417
0 51419 5 1 1 51418
0 51420 7 1 2 68148 51419
0 51421 5 1 1 51420
0 51422 7 1 2 86681 97637
0 51423 5 1 1 51422
0 51424 7 1 2 60405 51423
0 51425 5 1 1 51424
0 51426 7 1 2 65637 89428
0 51427 5 1 1 51426
0 51428 7 1 2 51425 51427
0 51429 5 1 1 51428
0 51430 7 1 2 96982 97865
0 51431 7 1 2 51429 51430
0 51432 5 1 1 51431
0 51433 7 1 2 51421 51432
0 51434 5 1 1 51433
0 51435 7 1 2 67757 51434
0 51436 5 1 1 51435
0 51437 7 5 2 64160 75359
0 51438 7 1 2 90118 88341
0 51439 7 1 2 98322 51438
0 51440 7 1 2 96536 51439
0 51441 5 1 1 51440
0 51442 7 1 2 51436 51441
0 51443 5 1 1 51442
0 51444 7 1 2 69604 51443
0 51445 5 1 1 51444
0 51446 7 1 2 96673 96696
0 51447 5 2 1 51446
0 51448 7 1 2 91184 97661
0 51449 5 1 1 51448
0 51450 7 1 2 98327 51449
0 51451 5 1 1 51450
0 51452 7 1 2 96249 51451
0 51453 5 1 1 51452
0 51454 7 1 2 64161 96017
0 51455 7 1 2 97198 51454
0 51456 5 1 1 51455
0 51457 7 1 2 51453 51456
0 51458 5 1 1 51457
0 51459 7 1 2 86185 51458
0 51460 5 1 1 51459
0 51461 7 6 2 94783 96925
0 51462 5 1 1 98329
0 51463 7 1 2 59679 82348
0 51464 5 1 1 51463
0 51465 7 1 2 8190 51464
0 51466 5 1 1 51465
0 51467 7 1 2 98330 51466
0 51468 5 1 1 51467
0 51469 7 1 2 60406 89425
0 51470 5 1 1 51469
0 51471 7 1 2 85919 88342
0 51472 5 1 1 51471
0 51473 7 1 2 51470 51472
0 51474 5 1 1 51473
0 51475 7 1 2 96526 51474
0 51476 5 1 1 51475
0 51477 7 1 2 21515 51476
0 51478 5 1 1 51477
0 51479 7 1 2 97876 51478
0 51480 5 1 1 51479
0 51481 7 1 2 51468 51480
0 51482 5 1 1 51481
0 51483 7 1 2 61801 51482
0 51484 5 1 1 51483
0 51485 7 1 2 49398 49394
0 51486 5 1 1 51485
0 51487 7 1 2 91702 51486
0 51488 5 1 1 51487
0 51489 7 2 2 75390 98024
0 51490 5 1 1 98335
0 51491 7 1 2 88343 98336
0 51492 5 1 1 51491
0 51493 7 1 2 51488 51492
0 51494 5 1 1 51493
0 51495 7 1 2 59680 51494
0 51496 5 1 1 51495
0 51497 7 1 2 91703 97920
0 51498 5 1 1 51497
0 51499 7 1 2 68786 51498
0 51500 7 1 2 51496 51499
0 51501 7 1 2 51484 51500
0 51502 5 1 1 51501
0 51503 7 1 2 78135 92811
0 51504 7 1 2 96926 51503
0 51505 5 1 1 51504
0 51506 7 1 2 98032 51505
0 51507 5 1 1 51506
0 51508 7 1 2 91704 51507
0 51509 5 1 1 51508
0 51510 7 1 2 51509 51490
0 51511 5 1 1 51510
0 51512 7 1 2 61802 51511
0 51513 5 1 1 51512
0 51514 7 1 2 93738 98025
0 51515 5 1 1 51514
0 51516 7 2 2 93987 96927
0 51517 7 1 2 87806 98337
0 51518 5 1 1 51517
0 51519 7 1 2 51515 51518
0 51520 5 1 1 51519
0 51521 7 1 2 60620 51520
0 51522 5 1 1 51521
0 51523 7 1 2 63853 51522
0 51524 7 1 2 51513 51523
0 51525 5 1 1 51524
0 51526 7 1 2 64058 51525
0 51527 7 1 2 51502 51526
0 51528 5 1 1 51527
0 51529 7 1 2 51460 51528
0 51530 7 1 2 51445 51529
0 51531 5 1 1 51530
0 51532 7 1 2 72257 51531
0 51533 5 1 1 51532
0 51534 7 1 2 84170 86594
0 51535 5 1 1 51534
0 51536 7 1 2 21758 51535
0 51537 5 1 1 51536
0 51538 7 1 2 92454 51537
0 51539 5 1 1 51538
0 51540 7 2 2 79681 83940
0 51541 5 1 1 98339
0 51542 7 1 2 86595 98340
0 51543 5 1 1 51542
0 51544 7 1 2 51539 51543
0 51545 5 1 1 51544
0 51546 7 1 2 83754 51545
0 51547 5 1 1 51546
0 51548 7 1 2 92675 96437
0 51549 5 1 1 51548
0 51550 7 1 2 51547 51549
0 51551 5 1 1 51550
0 51552 7 1 2 75360 51551
0 51553 5 1 1 51552
0 51554 7 1 2 76107 92525
0 51555 7 1 2 91920 51554
0 51556 7 1 2 94180 51555
0 51557 5 1 1 51556
0 51558 7 1 2 51553 51557
0 51559 5 1 1 51558
0 51560 7 1 2 64162 51559
0 51561 5 1 1 51560
0 51562 7 2 2 81002 77038
0 51563 7 1 2 98341 98300
0 51564 5 1 1 51563
0 51565 7 1 2 63585 88733
0 51566 5 2 1 51565
0 51567 7 2 2 83762 98343
0 51568 7 1 2 81003 96332
0 51569 7 1 2 98345 51568
0 51570 5 1 1 51569
0 51571 7 2 2 80985 98293
0 51572 7 1 2 96484 96039
0 51573 7 1 2 98347 51572
0 51574 5 1 1 51573
0 51575 7 1 2 51570 51574
0 51576 5 1 1 51575
0 51577 7 1 2 63854 51576
0 51578 5 1 1 51577
0 51579 7 1 2 79144 88090
0 51580 5 1 1 51579
0 51581 7 1 2 79750 82659
0 51582 7 1 2 81915 51581
0 51583 5 1 1 51582
0 51584 7 1 2 51580 51583
0 51585 5 1 1 51584
0 51586 7 1 2 75391 51585
0 51587 5 1 1 51586
0 51588 7 2 2 92054 94181
0 51589 7 1 2 90806 98349
0 51590 5 1 1 51589
0 51591 7 1 2 51587 51590
0 51592 5 1 1 51591
0 51593 7 1 2 94724 51592
0 51594 5 1 1 51593
0 51595 7 1 2 51578 51594
0 51596 5 1 1 51595
0 51597 7 1 2 67758 51596
0 51598 5 1 1 51597
0 51599 7 1 2 51564 51598
0 51600 7 1 2 51561 51599
0 51601 5 1 1 51600
0 51602 7 1 2 86805 51601
0 51603 5 1 1 51602
0 51604 7 1 2 96311 97624
0 51605 5 1 1 51604
0 51606 7 3 2 69025 75361
0 51607 7 1 2 83113 97515
0 51608 5 1 1 51607
0 51609 7 1 2 87646 51608
0 51610 5 1 1 51609
0 51611 7 2 2 98351 51610
0 51612 7 1 2 63855 98354
0 51613 5 1 1 51612
0 51614 7 1 2 85349 98204
0 51615 5 1 1 51614
0 51616 7 1 2 51613 51615
0 51617 5 1 1 51616
0 51618 7 1 2 96312 51617
0 51619 5 1 1 51618
0 51620 7 3 2 67759 81615
0 51621 5 1 1 98356
0 51622 7 1 2 63205 51621
0 51623 5 2 1 51622
0 51624 7 1 2 98359 98207
0 51625 5 1 1 51624
0 51626 7 4 2 89326 97754
0 51627 5 1 1 98361
0 51628 7 3 2 75362 96950
0 51629 7 1 2 92322 98365
0 51630 5 1 1 51629
0 51631 7 1 2 51627 51630
0 51632 5 1 1 51631
0 51633 7 1 2 88711 51632
0 51634 5 1 1 51633
0 51635 7 1 2 96491 98360
0 51636 5 1 1 51635
0 51637 7 1 2 68149 80337
0 51638 5 1 1 51637
0 51639 7 1 2 51636 51638
0 51640 5 1 1 51639
0 51641 7 1 2 86727 96898
0 51642 7 1 2 51640 51641
0 51643 5 1 1 51642
0 51644 7 1 2 51634 51643
0 51645 5 1 1 51644
0 51646 7 1 2 68540 51645
0 51647 5 1 1 51646
0 51648 7 1 2 51625 51647
0 51649 7 1 2 51619 51648
0 51650 5 1 1 51649
0 51651 7 1 2 64059 51650
0 51652 5 1 1 51651
0 51653 7 1 2 51605 51652
0 51654 7 1 2 51603 51653
0 51655 7 1 2 51533 51654
0 51656 5 1 1 51655
0 51657 7 1 2 95309 51656
0 51658 5 1 1 51657
0 51659 7 2 2 68946 97572
0 51660 5 1 1 98368
0 51661 7 2 2 80890 92735
0 51662 5 1 1 98370
0 51663 7 2 2 68947 71244
0 51664 7 1 2 92642 98372
0 51665 5 1 1 51664
0 51666 7 1 2 51662 51665
0 51667 5 1 1 51666
0 51668 7 1 2 75392 51667
0 51669 5 1 1 51668
0 51670 7 1 2 80541 76025
0 51671 7 1 2 96806 51670
0 51672 5 1 1 51671
0 51673 7 1 2 51669 51672
0 51674 5 1 1 51673
0 51675 7 1 2 68150 51674
0 51676 5 1 1 51675
0 51677 7 1 2 95939 98350
0 51678 5 1 1 51677
0 51679 7 1 2 51676 51678
0 51680 5 1 1 51679
0 51681 7 1 2 67128 51680
0 51682 5 1 1 51681
0 51683 7 1 2 51660 51682
0 51684 5 1 1 51683
0 51685 7 1 2 60727 51684
0 51686 5 1 1 51685
0 51687 7 1 2 87370 16080
0 51688 7 2 2 98373 51687
0 51689 7 1 2 74264 96082
0 51690 7 1 2 90524 51689
0 51691 7 1 2 98374 51690
0 51692 5 1 1 51691
0 51693 7 1 2 51686 51692
0 51694 5 1 1 51693
0 51695 7 1 2 66911 51694
0 51696 5 1 1 51695
0 51697 7 1 2 65638 80911
0 51698 5 1 1 51697
0 51699 7 1 2 94017 51698
0 51700 5 1 1 51699
0 51701 7 1 2 78136 97492
0 51702 5 1 1 51701
0 51703 7 1 2 51700 51702
0 51704 5 1 1 51703
0 51705 7 1 2 92736 51704
0 51706 5 1 1 51705
0 51707 7 2 2 71245 78266
0 51708 5 1 1 98376
0 51709 7 1 2 86145 88000
0 51710 7 1 2 98377 51709
0 51711 5 1 1 51710
0 51712 7 1 2 51706 51711
0 51713 5 1 1 51712
0 51714 7 1 2 61936 51713
0 51715 5 1 1 51714
0 51716 7 2 2 59681 74153
0 51717 7 1 2 87319 92305
0 51718 7 1 2 98378 51717
0 51719 5 1 1 51718
0 51720 7 1 2 51715 51719
0 51721 5 1 1 51720
0 51722 7 1 2 75363 51721
0 51723 5 1 1 51722
0 51724 7 1 2 95003 97570
0 51725 5 1 1 51724
0 51726 7 1 2 51723 51725
0 51727 5 1 1 51726
0 51728 7 1 2 68541 51727
0 51729 5 1 1 51728
0 51730 7 1 2 92812 98375
0 51731 5 1 1 51730
0 51732 7 1 2 59980 60728
0 51733 7 1 2 86222 51732
0 51734 5 1 1 51733
0 51735 7 1 2 51731 51734
0 51736 5 1 1 51735
0 51737 7 1 2 98297 51736
0 51738 5 1 1 51737
0 51739 7 1 2 75726 86223
0 51740 7 1 2 86740 51739
0 51741 7 1 2 92621 51740
0 51742 5 1 1 51741
0 51743 7 1 2 51738 51742
0 51744 5 1 1 51743
0 51745 7 1 2 75445 51744
0 51746 5 1 1 51745
0 51747 7 1 2 51729 51746
0 51748 7 1 2 51696 51747
0 51749 5 1 1 51748
0 51750 7 1 2 64163 51749
0 51751 5 1 1 51750
0 51752 7 1 2 96497 51340
0 51753 5 1 1 51752
0 51754 7 1 2 83192 51753
0 51755 5 1 1 51754
0 51756 7 1 2 96505 51755
0 51757 5 2 1 51756
0 51758 7 1 2 71246 98380
0 51759 5 1 1 51758
0 51760 7 2 2 75030 95475
0 51761 7 1 2 59981 92162
0 51762 7 2 2 98382 51761
0 51763 5 1 1 98384
0 51764 7 1 2 83207 89135
0 51765 5 1 1 51764
0 51766 7 1 2 91705 51765
0 51767 5 1 1 51766
0 51768 7 1 2 51763 51767
0 51769 5 1 1 51768
0 51770 7 1 2 66769 51769
0 51771 5 1 1 51770
0 51772 7 1 2 78137 97519
0 51773 5 1 1 51772
0 51774 7 1 2 74227 91625
0 51775 5 1 1 51774
0 51776 7 1 2 51773 51775
0 51777 5 1 1 51776
0 51778 7 1 2 79269 51777
0 51779 5 1 1 51778
0 51780 7 1 2 51771 51779
0 51781 5 1 1 51780
0 51782 7 1 2 67760 51781
0 51783 5 1 1 51782
0 51784 7 1 2 51759 51783
0 51785 5 1 1 51784
0 51786 7 1 2 96333 51785
0 51787 5 1 1 51786
0 51788 7 1 2 90182 97999
0 51789 5 1 1 51788
0 51790 7 2 2 68948 98323
0 51791 7 1 2 80891 71247
0 51792 7 1 2 86541 51791
0 51793 7 1 2 98386 51792
0 51794 5 1 1 51793
0 51795 7 1 2 51789 51794
0 51796 7 1 2 51787 51795
0 51797 5 1 1 51796
0 51798 7 1 2 86728 51797
0 51799 5 1 1 51798
0 51800 7 1 2 68787 51799
0 51801 7 1 2 51751 51800
0 51802 5 1 1 51801
0 51803 7 1 2 74949 97831
0 51804 5 1 1 51803
0 51805 7 1 2 51462 51804
0 51806 5 1 1 51805
0 51807 7 1 2 60407 51806
0 51808 5 1 1 51807
0 51809 7 1 2 51808 98212
0 51810 5 1 1 51809
0 51811 7 1 2 85685 51810
0 51812 5 1 1 51811
0 51813 7 1 2 96640 97741
0 51814 5 1 1 51813
0 51815 7 1 2 51812 51814
0 51816 5 1 1 51815
0 51817 7 1 2 68151 51816
0 51818 5 1 1 51817
0 51819 7 1 2 71248 97863
0 51820 5 1 1 51819
0 51821 7 1 2 97742 97973
0 51822 5 1 1 51821
0 51823 7 1 2 51820 51822
0 51824 5 1 1 51823
0 51825 7 1 2 88837 51824
0 51826 5 1 1 51825
0 51827 7 2 2 59982 97475
0 51828 7 1 2 86359 95707
0 51829 7 1 2 95540 51828
0 51830 7 1 2 98388 51829
0 51831 5 1 1 51830
0 51832 7 1 2 51826 51831
0 51833 5 1 1 51832
0 51834 7 1 2 75364 51833
0 51835 5 1 1 51834
0 51836 7 1 2 66770 20933
0 51837 5 1 1 51836
0 51838 7 2 2 97743 51837
0 51839 7 1 2 73470 98390
0 51840 5 1 1 51839
0 51841 7 1 2 32439 51840
0 51842 5 1 1 51841
0 51843 7 2 2 67129 79858
0 51844 5 1 1 98392
0 51845 7 1 2 67761 98393
0 51846 5 1 1 51845
0 51847 7 1 2 84841 51846
0 51848 5 1 1 51847
0 51849 7 1 2 51842 51848
0 51850 5 1 1 51849
0 51851 7 1 2 90491 89429
0 51852 7 1 2 98391 51851
0 51853 5 1 1 51852
0 51854 7 1 2 68949 51853
0 51855 7 1 2 51850 51854
0 51856 7 1 2 51835 51855
0 51857 7 1 2 51818 51856
0 51858 5 1 1 51857
0 51859 7 1 2 79958 76108
0 51860 5 1 1 51859
0 51861 7 1 2 71249 74740
0 51862 5 1 1 51861
0 51863 7 1 2 51860 51862
0 51864 5 1 1 51863
0 51865 7 1 2 77933 51864
0 51866 5 1 1 51865
0 51867 7 1 2 48371 51866
0 51868 5 1 1 51867
0 51869 7 1 2 87193 51868
0 51870 5 1 1 51869
0 51871 7 1 2 62156 92869
0 51872 7 1 2 85724 51871
0 51873 7 1 2 96204 51872
0 51874 5 1 1 51873
0 51875 7 1 2 51870 51874
0 51876 5 1 1 51875
0 51877 7 1 2 66771 51876
0 51878 5 1 1 51877
0 51879 7 1 2 75128 51708
0 51880 5 1 1 51879
0 51881 7 1 2 89327 51880
0 51882 5 1 1 51881
0 51883 7 1 2 93188 96156
0 51884 5 1 1 51883
0 51885 7 1 2 51882 51884
0 51886 5 1 1 51885
0 51887 7 1 2 86729 51886
0 51888 5 1 1 51887
0 51889 7 1 2 51878 51888
0 51890 5 1 1 51889
0 51891 7 1 2 69026 51890
0 51892 5 1 1 51891
0 51893 7 3 2 68542 71250
0 51894 5 1 1 98394
0 51895 7 1 2 97271 51894
0 51896 5 1 1 51895
0 51897 7 1 2 89491 51896
0 51898 5 1 1 51897
0 51899 7 1 2 61611 97281
0 51900 5 1 1 51899
0 51901 7 1 2 51898 51900
0 51902 5 1 1 51901
0 51903 7 1 2 79682 51902
0 51904 5 1 1 51903
0 51905 7 1 2 80892 81703
0 51906 5 1 1 51905
0 51907 7 1 2 51904 51906
0 51908 5 1 1 51907
0 51909 7 1 2 95636 51908
0 51910 5 1 1 51909
0 51911 7 1 2 51892 51910
0 51912 5 1 1 51911
0 51913 7 1 2 59682 51912
0 51914 5 1 1 51913
0 51915 7 1 2 67130 98355
0 51916 5 1 1 51915
0 51917 7 1 2 72258 98338
0 51918 5 1 1 51917
0 51919 7 1 2 98033 51918
0 51920 5 1 1 51919
0 51921 7 1 2 75365 97974
0 51922 7 1 2 51920 51921
0 51923 5 1 1 51922
0 51924 7 1 2 64060 51923
0 51925 7 1 2 51916 51924
0 51926 7 1 2 51914 51925
0 51927 5 1 1 51926
0 51928 7 1 2 51858 51927
0 51929 5 1 1 51928
0 51930 7 1 2 63856 51929
0 51931 5 1 1 51930
0 51932 7 1 2 95310 51931
0 51933 7 1 2 51802 51932
0 51934 5 1 1 51933
0 51935 7 1 2 61134 97705
0 51936 5 1 1 51935
0 51937 7 1 2 59983 97030
0 51938 5 1 1 51937
0 51939 7 1 2 87803 94220
0 51940 7 2 2 97773 51939
0 51941 5 1 1 98397
0 51942 7 1 2 67131 98398
0 51943 5 1 1 51942
0 51944 7 1 2 51938 51943
0 51945 5 1 1 51944
0 51946 7 1 2 68950 51945
0 51947 5 1 1 51946
0 51948 7 2 2 95311 98172
0 51949 5 1 1 98399
0 51950 7 1 2 67132 98400
0 51951 5 1 1 51950
0 51952 7 1 2 51947 51951
0 51953 5 1 1 51952
0 51954 7 1 2 88958 51953
0 51955 5 1 1 51954
0 51956 7 1 2 51936 51955
0 51957 7 1 2 51934 51956
0 51958 5 1 1 51957
0 51959 7 1 2 69963 51958
0 51960 5 1 1 51959
0 51961 7 1 2 79751 96707
0 51962 5 2 1 51961
0 51963 7 2 2 68543 96700
0 51964 5 1 1 98403
0 51965 7 1 2 88883 98404
0 51966 5 1 1 51965
0 51967 7 1 2 98401 51966
0 51968 5 1 1 51967
0 51969 7 1 2 97761 51968
0 51970 5 1 1 51969
0 51971 7 2 2 78164 44104
0 51972 7 1 2 72259 98405
0 51973 5 1 1 51972
0 51974 7 1 2 96139 97565
0 51975 5 1 1 51974
0 51976 7 1 2 82276 84295
0 51977 5 1 1 51976
0 51978 7 1 2 89958 51977
0 51979 5 1 1 51978
0 51980 7 1 2 91706 51979
0 51981 5 1 1 51980
0 51982 7 1 2 82003 79233
0 51983 5 1 1 51982
0 51984 7 1 2 51981 51983
0 51985 5 1 1 51984
0 51986 7 1 2 86806 51985
0 51987 5 1 1 51986
0 51988 7 1 2 51975 51987
0 51989 7 1 2 51973 51988
0 51990 5 1 1 51989
0 51991 7 1 2 68951 51990
0 51992 5 1 1 51991
0 51993 7 1 2 83755 92839
0 51994 7 1 2 96701 51993
0 51995 5 1 1 51994
0 51996 7 1 2 51992 51995
0 51997 5 1 1 51996
0 51998 7 1 2 64164 51997
0 51999 5 1 1 51998
0 52000 7 1 2 51970 51999
0 52001 5 1 1 52000
0 52002 7 1 2 95312 52001
0 52003 5 1 1 52002
0 52004 7 1 2 61937 89642
0 52005 7 1 2 92701 52004
0 52006 7 1 2 97558 52005
0 52007 5 1 1 52006
0 52008 7 1 2 52003 52007
0 52009 5 1 1 52008
0 52010 7 1 2 73363 52009
0 52011 5 1 1 52010
0 52012 7 1 2 92257 97007
0 52013 5 1 1 52012
0 52014 7 1 2 98389 98183
0 52015 7 1 2 96990 52014
0 52016 5 1 1 52015
0 52017 7 1 2 52013 52016
0 52018 5 1 1 52017
0 52019 7 1 2 84446 52018
0 52020 5 1 1 52019
0 52021 7 2 2 94161 96334
0 52022 7 1 2 88051 90082
0 52023 7 1 2 98407 52022
0 52024 5 1 1 52023
0 52025 7 1 2 52020 52024
0 52026 5 1 1 52025
0 52027 7 1 2 95313 52026
0 52028 5 1 1 52027
0 52029 7 1 2 96083 97028
0 52030 7 1 2 97700 52029
0 52031 5 1 1 52030
0 52032 7 1 2 52028 52031
0 52033 5 1 1 52032
0 52034 7 1 2 83888 52033
0 52035 5 1 1 52034
0 52036 7 1 2 52011 52035
0 52037 7 1 2 51960 52036
0 52038 7 1 2 51658 52037
0 52039 7 1 2 51383 52038
0 52040 5 1 1 52039
0 52041 7 1 2 70211 52040
0 52042 5 1 1 52041
0 52043 7 2 2 68952 91886
0 52044 5 1 1 98409
0 52045 7 1 2 92037 96781
0 52046 5 1 1 52045
0 52047 7 1 2 52044 52046
0 52048 5 1 1 52047
0 52049 7 1 2 69605 52048
0 52050 5 1 1 52049
0 52051 7 1 2 10245 52050
0 52052 5 1 1 52051
0 52053 7 1 2 59683 52052
0 52054 5 1 1 52053
0 52055 7 1 2 86146 92643
0 52056 5 1 1 52055
0 52057 7 1 2 52054 52056
0 52058 5 1 1 52057
0 52059 7 1 2 68544 52058
0 52060 5 1 1 52059
0 52061 7 1 2 92055 95933
0 52062 5 1 1 52061
0 52063 7 1 2 52060 52062
0 52064 5 1 1 52063
0 52065 7 1 2 68788 52064
0 52066 5 1 1 52065
0 52067 7 3 2 63857 76280
0 52068 7 2 2 68953 98411
0 52069 5 1 1 98414
0 52070 7 1 2 82004 98415
0 52071 5 1 1 52070
0 52072 7 1 2 52066 52071
0 52073 5 1 1 52072
0 52074 7 1 2 91707 52073
0 52075 5 1 1 52074
0 52076 7 1 2 75855 88716
0 52077 5 1 1 52076
0 52078 7 1 2 5671 52077
0 52079 5 1 1 52078
0 52080 7 1 2 87266 90208
0 52081 7 1 2 52079 52080
0 52082 5 1 1 52081
0 52083 7 1 2 52075 52082
0 52084 5 1 1 52083
0 52085 7 1 2 61938 52084
0 52086 5 1 1 52085
0 52087 7 1 2 68954 94637
0 52088 7 1 2 96018 52087
0 52089 7 1 2 88717 52088
0 52090 5 1 1 52089
0 52091 7 1 2 65639 52090
0 52092 7 1 2 52086 52091
0 52093 5 1 1 52092
0 52094 7 1 2 86261 92873
0 52095 5 1 1 52094
0 52096 7 1 2 74976 92038
0 52097 7 1 2 93942 52096
0 52098 5 1 1 52097
0 52099 7 1 2 52069 52098
0 52100 5 1 1 52099
0 52101 7 2 2 66912 52100
0 52102 5 1 1 98416
0 52103 7 1 2 61803 98417
0 52104 5 1 1 52103
0 52105 7 1 2 52095 52104
0 52106 5 1 1 52105
0 52107 7 1 2 91708 52106
0 52108 5 1 1 52107
0 52109 7 1 2 64061 84847
0 52110 7 1 2 91750 52109
0 52111 5 2 1 52110
0 52112 7 1 2 79234 86186
0 52113 5 1 1 52112
0 52114 7 1 2 98418 52113
0 52115 5 1 1 52114
0 52116 7 1 2 61804 52115
0 52117 5 1 1 52116
0 52118 7 1 2 27982 48675
0 52119 5 1 1 52118
0 52120 7 1 2 91709 52119
0 52121 5 1 1 52120
0 52122 7 1 2 52117 52121
0 52123 5 1 1 52122
0 52124 7 1 2 88718 52123
0 52125 5 1 1 52124
0 52126 7 1 2 27914 52102
0 52127 5 1 1 52126
0 52128 7 1 2 90183 52127
0 52129 5 1 1 52128
0 52130 7 1 2 52125 52129
0 52131 7 1 2 52108 52130
0 52132 5 1 1 52131
0 52133 7 1 2 68545 52132
0 52134 5 1 1 52133
0 52135 7 2 2 81616 83570
0 52136 5 1 1 98420
0 52137 7 1 2 84558 52136
0 52138 5 1 1 52137
0 52139 7 1 2 87304 52138
0 52140 5 1 1 52139
0 52141 7 1 2 49158 52140
0 52142 5 1 1 52141
0 52143 7 1 2 91710 52142
0 52144 5 1 1 52143
0 52145 7 1 2 61805 98421
0 52146 5 1 1 52145
0 52147 7 1 2 3175 52146
0 52148 5 1 1 52147
0 52149 7 1 2 73488 90184
0 52150 7 1 2 52148 52149
0 52151 5 1 1 52150
0 52152 7 1 2 52144 52151
0 52153 5 1 1 52152
0 52154 7 1 2 67762 52153
0 52155 5 1 1 52154
0 52156 7 1 2 60729 52155
0 52157 7 1 2 52134 52156
0 52158 5 1 1 52157
0 52159 7 1 2 64165 52158
0 52160 7 1 2 52093 52159
0 52161 5 1 1 52160
0 52162 7 1 2 96609 98138
0 52163 5 2 1 52162
0 52164 7 1 2 91711 98422
0 52165 5 1 1 52164
0 52166 7 1 2 40264 52165
0 52167 5 1 1 52166
0 52168 7 1 2 70698 52167
0 52169 5 1 1 52168
0 52170 7 1 2 90209 96713
0 52171 5 1 1 52170
0 52172 7 1 2 52169 52171
0 52173 5 1 1 52172
0 52174 7 1 2 66913 52173
0 52175 5 1 1 52174
0 52176 7 2 2 70699 74104
0 52177 7 1 2 83114 86557
0 52178 7 1 2 98424 52177
0 52179 5 1 1 52178
0 52180 7 1 2 52175 52179
0 52181 5 1 1 52180
0 52182 7 1 2 76281 52181
0 52183 5 1 1 52182
0 52184 7 1 2 92862 94466
0 52185 5 1 1 52184
0 52186 7 1 2 75746 85725
0 52187 5 1 1 52186
0 52188 7 1 2 77039 94476
0 52189 5 1 1 52188
0 52190 7 1 2 52187 52189
0 52191 5 1 1 52190
0 52192 7 1 2 85854 52191
0 52193 5 1 1 52192
0 52194 7 1 2 80963 77040
0 52195 5 1 1 52194
0 52196 7 1 2 87766 52195
0 52197 5 1 1 52196
0 52198 7 1 2 96991 52197
0 52199 5 1 1 52198
0 52200 7 1 2 81813 85920
0 52201 7 1 2 92806 52200
0 52202 5 1 1 52201
0 52203 7 1 2 52199 52202
0 52204 5 1 1 52203
0 52205 7 1 2 66914 52204
0 52206 5 1 1 52205
0 52207 7 1 2 52193 52206
0 52208 5 1 1 52207
0 52209 7 1 2 63858 52208
0 52210 5 1 1 52209
0 52211 7 1 2 52185 52210
0 52212 7 1 2 52183 52211
0 52213 5 1 1 52212
0 52214 7 1 2 64062 52213
0 52215 5 1 1 52214
0 52216 7 1 2 88719 96880
0 52217 5 1 1 52216
0 52218 7 2 2 68546 88008
0 52219 5 1 1 98426
0 52220 7 1 2 76282 98427
0 52221 5 1 1 52220
0 52222 7 1 2 52217 52221
0 52223 5 1 1 52222
0 52224 7 1 2 84447 94646
0 52225 7 1 2 52223 52224
0 52226 5 1 1 52225
0 52227 7 1 2 52215 52226
0 52228 5 1 1 52227
0 52229 7 1 2 65640 52228
0 52230 5 1 1 52229
0 52231 7 1 2 81004 78201
0 52232 7 1 2 87870 52231
0 52233 7 2 2 66915 83193
0 52234 7 1 2 95812 98428
0 52235 7 1 2 52232 52234
0 52236 5 1 1 52235
0 52237 7 1 2 52230 52236
0 52238 5 1 1 52237
0 52239 7 1 2 69027 52238
0 52240 5 1 1 52239
0 52241 7 1 2 87669 94221
0 52242 7 1 2 96849 52241
0 52243 5 1 1 52242
0 52244 7 1 2 43904 52243
0 52245 5 2 1 52244
0 52246 7 1 2 97120 98430
0 52247 5 1 1 52246
0 52248 7 2 2 61939 97734
0 52249 7 2 2 82005 97790
0 52250 7 1 2 98432 98434
0 52251 5 1 1 52250
0 52252 7 1 2 52247 52251
0 52253 5 1 1 52252
0 52254 7 1 2 67133 52253
0 52255 5 1 1 52254
0 52256 7 1 2 83509 98433
0 52257 7 1 2 98151 52256
0 52258 5 1 1 52257
0 52259 7 1 2 52255 52258
0 52260 5 1 1 52259
0 52261 7 1 2 67763 52260
0 52262 5 1 1 52261
0 52263 7 1 2 61806 93977
0 52264 7 1 2 98282 52263
0 52265 5 1 1 52264
0 52266 7 1 2 82196 96914
0 52267 7 1 2 97102 52266
0 52268 5 1 1 52267
0 52269 7 1 2 52265 52268
0 52270 5 1 1 52269
0 52271 7 1 2 62770 52270
0 52272 5 1 1 52271
0 52273 7 1 2 76428 95621
0 52274 7 1 2 95719 52273
0 52275 7 1 2 96782 97929
0 52276 7 1 2 52274 52275
0 52277 5 1 1 52276
0 52278 7 1 2 52272 52277
0 52279 7 1 2 52262 52278
0 52280 5 1 1 52279
0 52281 7 1 2 64063 52280
0 52282 5 1 1 52281
0 52283 7 1 2 86393 96600
0 52284 7 1 2 96294 52283
0 52285 5 1 1 52284
0 52286 7 1 2 52282 52285
0 52287 5 1 1 52286
0 52288 7 1 2 97800 52287
0 52289 5 1 1 52288
0 52290 7 1 2 52240 52289
0 52291 7 1 2 52161 52290
0 52292 5 1 1 52291
0 52293 7 1 2 95314 52292
0 52294 5 1 1 52293
0 52295 7 1 2 81814 82935
0 52296 7 1 2 90814 52295
0 52297 7 1 2 95262 52296
0 52298 7 1 2 98260 52297
0 52299 5 1 1 52298
0 52300 7 1 2 52294 52299
0 52301 5 1 1 52300
0 52302 7 1 2 71251 52301
0 52303 5 1 1 52302
0 52304 7 1 2 83115 92870
0 52305 7 1 2 95805 52304
0 52306 7 1 2 97715 52305
0 52307 5 1 1 52306
0 52308 7 1 2 71252 86332
0 52309 5 1 1 52308
0 52310 7 2 2 61135 86187
0 52311 7 1 2 82591 98436
0 52312 5 1 1 52311
0 52313 7 1 2 52309 52312
0 52314 5 1 1 52313
0 52315 7 1 2 97373 97735
0 52316 7 1 2 52314 52315
0 52317 5 1 1 52316
0 52318 7 1 2 52307 52317
0 52319 5 1 1 52318
0 52320 7 1 2 79683 52319
0 52321 5 1 1 52320
0 52322 7 1 2 68789 98395
0 52323 7 1 2 97516 52322
0 52324 5 1 1 52323
0 52325 7 1 2 72260 87297
0 52326 7 1 2 97554 52325
0 52327 5 1 1 52326
0 52328 7 1 2 52324 52327
0 52329 5 1 1 52328
0 52330 7 1 2 97597 52329
0 52331 5 1 1 52330
0 52332 7 1 2 52321 52331
0 52333 5 1 1 52332
0 52334 7 1 2 95315 52333
0 52335 5 1 1 52334
0 52336 7 1 2 48129 52335
0 52337 5 1 1 52336
0 52338 7 1 2 59684 52337
0 52339 5 1 1 52338
0 52340 7 1 2 84448 97765
0 52341 7 1 2 98074 52340
0 52342 5 1 1 52341
0 52343 7 1 2 52339 52342
0 52344 5 1 1 52343
0 52345 7 1 2 83889 52344
0 52346 5 1 1 52345
0 52347 7 1 2 96431 97063
0 52348 5 1 1 52347
0 52349 7 1 2 91837 52348
0 52350 5 1 1 52349
0 52351 7 1 2 68547 52350
0 52352 5 1 1 52351
0 52353 7 1 2 72414 35188
0 52354 5 1 1 52353
0 52355 7 1 2 96459 52354
0 52356 5 1 1 52355
0 52357 7 1 2 84820 52356
0 52358 5 1 1 52357
0 52359 7 1 2 52352 52358
0 52360 5 1 1 52359
0 52361 7 1 2 86765 52360
0 52362 5 1 1 52361
0 52363 7 1 2 92221 35127
0 52364 5 1 1 52363
0 52365 7 1 2 77934 52364
0 52366 5 1 1 52365
0 52367 7 1 2 89673 52366
0 52368 5 1 1 52367
0 52369 7 1 2 69437 52368
0 52370 5 1 1 52369
0 52371 7 1 2 71253 82349
0 52372 5 1 1 52371
0 52373 7 1 2 85955 52372
0 52374 5 1 1 52373
0 52375 7 1 2 59397 52374
0 52376 5 1 1 52375
0 52377 7 1 2 95207 52376
0 52378 5 1 1 52377
0 52379 7 1 2 76063 52378
0 52380 5 1 1 52379
0 52381 7 1 2 84679 85956
0 52382 5 1 1 52381
0 52383 7 1 2 59984 52382
0 52384 5 1 1 52383
0 52385 7 1 2 40224 52384
0 52386 7 1 2 52380 52385
0 52387 7 1 2 52370 52386
0 52388 5 1 1 52387
0 52389 7 1 2 68790 96529
0 52390 7 1 2 52388 52389
0 52391 5 1 1 52390
0 52392 7 1 2 52362 52391
0 52393 5 1 1 52392
0 52394 7 1 2 64166 52393
0 52395 5 1 1 52394
0 52396 7 1 2 64591 39416
0 52397 5 1 1 52396
0 52398 7 1 2 84661 94868
0 52399 7 1 2 52397 52398
0 52400 5 1 1 52399
0 52401 7 1 2 72385 52400
0 52402 5 1 1 52401
0 52403 7 1 2 67764 52402
0 52404 5 1 1 52403
0 52405 7 1 2 95690 52404
0 52406 5 1 1 52405
0 52407 7 1 2 98061 52406
0 52408 5 1 1 52407
0 52409 7 1 2 62771 92971
0 52410 5 1 1 52409
0 52411 7 1 2 68152 95211
0 52412 7 1 2 52410 52411
0 52413 5 1 1 52412
0 52414 7 1 2 71899 96255
0 52415 5 1 1 52414
0 52416 7 1 2 52413 52415
0 52417 5 1 1 52416
0 52418 7 1 2 98055 52417
0 52419 5 1 1 52418
0 52420 7 1 2 52408 52419
0 52421 7 1 2 52395 52420
0 52422 5 1 1 52421
0 52423 7 1 2 70700 52422
0 52424 5 1 1 52423
0 52425 7 1 2 72386 98100
0 52426 5 1 1 52425
0 52427 7 1 2 59685 52426
0 52428 5 1 1 52427
0 52429 7 1 2 74807 88450
0 52430 5 1 1 52429
0 52431 7 1 2 52428 52430
0 52432 5 1 1 52431
0 52433 7 1 2 85490 52432
0 52434 5 1 1 52433
0 52435 7 1 2 15420 52434
0 52436 5 1 1 52435
0 52437 7 1 2 79684 52436
0 52438 5 1 1 52437
0 52439 7 1 2 82796 88451
0 52440 5 1 1 52439
0 52441 7 1 2 90506 52440
0 52442 5 1 1 52441
0 52443 7 1 2 83756 84368
0 52444 7 1 2 52442 52443
0 52445 5 1 1 52444
0 52446 7 1 2 85296 52445
0 52447 7 1 2 52438 52446
0 52448 5 1 1 52447
0 52449 7 1 2 95637 52448
0 52450 5 1 1 52449
0 52451 7 1 2 76283 98423
0 52452 5 1 1 52451
0 52453 7 1 2 39987 98098
0 52454 5 1 1 52453
0 52455 7 1 2 69964 52454
0 52456 5 1 1 52455
0 52457 7 1 2 52452 52456
0 52458 5 1 1 52457
0 52459 7 1 2 71254 52458
0 52460 5 1 1 52459
0 52461 7 1 2 68153 73240
0 52462 5 1 1 52461
0 52463 7 1 2 88936 88885
0 52464 7 1 2 52462 52463
0 52465 5 1 1 52464
0 52466 7 1 2 84527 52465
0 52467 5 1 1 52466
0 52468 7 1 2 83941 84287
0 52469 5 1 1 52468
0 52470 7 1 2 68154 97937
0 52471 5 1 1 52470
0 52472 7 1 2 52469 52471
0 52473 5 1 1 52472
0 52474 7 1 2 76934 52473
0 52475 5 1 1 52474
0 52476 7 1 2 89959 52475
0 52477 7 1 2 52467 52476
0 52478 7 1 2 52460 52477
0 52479 5 1 1 52478
0 52480 7 1 2 97671 52479
0 52481 5 1 1 52480
0 52482 7 1 2 64064 52481
0 52483 7 1 2 52450 52482
0 52484 7 1 2 52424 52483
0 52485 5 1 1 52484
0 52486 7 1 2 84312 97681
0 52487 5 1 1 52486
0 52488 7 1 2 61136 92777
0 52489 7 1 2 94638 52488
0 52490 7 1 2 97560 52489
0 52491 5 1 1 52490
0 52492 7 1 2 52487 52491
0 52493 5 1 1 52492
0 52494 7 1 2 73387 52493
0 52495 5 1 1 52494
0 52496 7 1 2 76935 97374
0 52497 5 1 1 52496
0 52498 7 1 2 90265 96511
0 52499 5 1 1 52498
0 52500 7 1 2 52497 52499
0 52501 5 1 1 52500
0 52502 7 1 2 71255 52501
0 52503 5 1 1 52502
0 52504 7 2 2 68791 98102
0 52505 7 1 2 92815 98438
0 52506 5 1 1 52505
0 52507 7 1 2 52503 52506
0 52508 5 1 1 52507
0 52509 7 1 2 92009 94352
0 52510 7 1 2 52508 52509
0 52511 5 1 1 52510
0 52512 7 1 2 52495 52511
0 52513 5 1 1 52512
0 52514 7 1 2 64167 52513
0 52515 5 1 1 52514
0 52516 7 1 2 68955 98114
0 52517 7 1 2 52515 52516
0 52518 5 1 1 52517
0 52519 7 1 2 52485 52518
0 52520 5 1 1 52519
0 52521 7 1 2 89145 89695
0 52522 5 1 1 52521
0 52523 7 1 2 70866 89136
0 52524 5 1 1 52523
0 52525 7 5 2 68548 76284
0 52526 5 1 1 98440
0 52527 7 1 2 63859 98441
0 52528 7 1 2 52524 52527
0 52529 5 1 1 52528
0 52530 7 1 2 52522 52529
0 52531 5 1 1 52530
0 52532 7 1 2 67765 52531
0 52533 5 1 1 52532
0 52534 7 1 2 83222 20522
0 52535 5 1 1 52534
0 52536 7 1 2 68155 52535
0 52537 5 1 1 52536
0 52538 7 1 2 96277 52537
0 52539 7 1 2 52533 52538
0 52540 5 1 1 52539
0 52541 7 1 2 79685 52540
0 52542 5 1 1 52541
0 52543 7 2 2 79449 90060
0 52544 5 1 1 98445
0 52545 7 1 2 98439 98446
0 52546 5 1 1 52545
0 52547 7 1 2 79450 87894
0 52548 7 1 2 88619 52547
0 52549 5 1 1 52548
0 52550 7 1 2 91772 52549
0 52551 5 1 1 52550
0 52552 7 1 2 73364 52551
0 52553 5 1 1 52552
0 52554 7 1 2 52546 52553
0 52555 7 1 2 52542 52554
0 52556 5 1 1 52555
0 52557 7 1 2 68956 52556
0 52558 5 1 1 52557
0 52559 7 1 2 80893 72261
0 52560 7 1 2 97494 52559
0 52561 7 1 2 88712 52560
0 52562 5 1 1 52561
0 52563 7 1 2 52558 52562
0 52564 5 1 1 52563
0 52565 7 1 2 64168 52564
0 52566 5 1 1 52565
0 52567 7 2 2 67134 97658
0 52568 5 1 1 98447
0 52569 7 1 2 98328 52568
0 52570 5 1 1 52569
0 52571 7 1 2 69606 52570
0 52572 5 1 1 52571
0 52573 7 1 2 59686 98448
0 52574 5 1 1 52573
0 52575 7 1 2 52572 52574
0 52576 5 1 1 52575
0 52577 7 1 2 64065 52576
0 52578 5 1 1 52577
0 52579 7 1 2 86305 91887
0 52580 5 1 1 52579
0 52581 7 1 2 96440 52580
0 52582 5 1 1 52581
0 52583 7 1 2 96983 52582
0 52584 5 1 1 52583
0 52585 7 1 2 52578 52584
0 52586 5 1 1 52585
0 52587 7 1 2 67766 52586
0 52588 5 1 1 52587
0 52589 7 1 2 84629 97794
0 52590 5 1 1 52589
0 52591 7 2 2 61807 94770
0 52592 7 1 2 76285 86306
0 52593 7 1 2 98449 52592
0 52594 5 1 1 52593
0 52595 7 1 2 52590 52594
0 52596 5 1 1 52595
0 52597 7 1 2 63860 52596
0 52598 5 1 1 52597
0 52599 7 1 2 52588 52598
0 52600 5 1 1 52599
0 52601 7 1 2 71256 52600
0 52602 5 1 1 52601
0 52603 7 1 2 92647 96943
0 52604 5 1 1 52603
0 52605 7 1 2 79686 91597
0 52606 7 1 2 96984 52605
0 52607 5 1 1 52606
0 52608 7 1 2 52604 52607
0 52609 5 1 1 52608
0 52610 7 1 2 63206 52609
0 52611 5 1 1 52610
0 52612 7 1 2 84449 96335
0 52613 7 1 2 84630 52612
0 52614 5 1 1 52613
0 52615 7 1 2 52611 52614
0 52616 5 1 1 52615
0 52617 7 1 2 63586 52616
0 52618 5 1 1 52617
0 52619 7 2 2 61808 74105
0 52620 7 1 2 91367 95476
0 52621 7 1 2 97727 52620
0 52622 7 1 2 98451 52621
0 52623 5 1 1 52622
0 52624 7 1 2 52618 52623
0 52625 5 1 1 52624
0 52626 7 1 2 59687 52625
0 52627 5 1 1 52626
0 52628 7 1 2 97985 98161
0 52629 5 1 1 52628
0 52630 7 2 2 70701 89820
0 52631 5 1 1 98453
0 52632 7 1 2 93181 97534
0 52633 5 1 1 52632
0 52634 7 1 2 52631 52633
0 52635 5 1 1 52634
0 52636 7 1 2 64169 80986
0 52637 7 1 2 52635 52636
0 52638 5 1 1 52637
0 52639 7 1 2 52629 52638
0 52640 5 1 1 52639
0 52641 7 1 2 63861 52640
0 52642 5 1 1 52641
0 52643 7 1 2 92056 97535
0 52644 5 1 1 52643
0 52645 7 1 2 78138 98371
0 52646 5 1 1 52645
0 52647 7 1 2 68957 96850
0 52648 5 1 1 52647
0 52649 7 1 2 52646 52648
0 52650 5 1 1 52649
0 52651 7 1 2 68549 73830
0 52652 7 1 2 52650 52651
0 52653 5 1 1 52652
0 52654 7 1 2 52644 52653
0 52655 5 1 1 52654
0 52656 7 1 2 94725 52655
0 52657 5 1 1 52656
0 52658 7 1 2 52642 52657
0 52659 5 1 1 52658
0 52660 7 1 2 59985 52659
0 52661 5 1 1 52660
0 52662 7 1 2 80912 89225
0 52663 5 1 1 52662
0 52664 7 1 2 91834 52663
0 52665 5 1 1 52664
0 52666 7 1 2 91513 89754
0 52667 5 1 1 52666
0 52668 7 1 2 52665 52667
0 52669 5 1 1 52668
0 52670 7 1 2 67767 52669
0 52671 5 1 1 52670
0 52672 7 1 2 82660 98435
0 52673 5 1 1 52672
0 52674 7 1 2 52671 52673
0 52675 5 1 1 52674
0 52676 7 1 2 94771 52675
0 52677 5 1 1 52676
0 52678 7 1 2 52661 52677
0 52679 7 1 2 52627 52678
0 52680 5 1 1 52679
0 52681 7 1 2 69965 52680
0 52682 5 1 1 52681
0 52683 7 1 2 83785 84272
0 52684 7 1 2 94230 52683
0 52685 7 1 2 96313 52684
0 52686 5 1 1 52685
0 52687 7 1 2 52682 52686
0 52688 7 1 2 52602 52687
0 52689 7 1 2 52566 52688
0 52690 5 1 1 52689
0 52691 7 1 2 86807 52690
0 52692 5 1 1 52691
0 52693 7 1 2 52520 52692
0 52694 5 1 1 52693
0 52695 7 1 2 95316 52694
0 52696 5 1 1 52695
0 52697 7 1 2 52346 52696
0 52698 5 1 1 52697
0 52699 7 1 2 75366 52698
0 52700 5 1 1 52699
0 52701 7 1 2 80776 97774
0 52702 7 1 2 98226 52701
0 52703 5 1 1 52702
0 52704 7 1 2 66953 81500
0 52705 7 2 2 89097 52704
0 52706 7 1 2 61940 86596
0 52707 7 1 2 95263 52706
0 52708 7 1 2 98455 52707
0 52709 5 1 1 52708
0 52710 7 1 2 52703 52709
0 52711 5 1 1 52710
0 52712 7 1 2 95970 52711
0 52713 5 1 1 52712
0 52714 7 1 2 70702 80176
0 52715 5 1 1 52714
0 52716 7 1 2 81129 52715
0 52717 5 1 1 52716
0 52718 7 1 2 60408 52717
0 52719 5 1 1 52718
0 52720 7 2 2 97711 52719
0 52721 7 1 2 79968 80338
0 52722 5 1 1 52721
0 52723 7 1 2 98457 52722
0 52724 5 1 1 52723
0 52725 7 1 2 59688 52724
0 52726 5 1 1 52725
0 52727 7 1 2 92458 96881
0 52728 5 1 1 52727
0 52729 7 1 2 52726 52728
0 52730 5 1 1 52729
0 52731 7 1 2 64066 97775
0 52732 7 1 2 52730 52731
0 52733 5 1 1 52732
0 52734 7 1 2 52713 52733
0 52735 5 1 1 52734
0 52736 7 1 2 68792 52735
0 52737 5 1 1 52736
0 52738 7 1 2 77041 86148
0 52739 5 1 1 52738
0 52740 7 1 2 86125 52739
0 52741 5 1 1 52740
0 52742 7 1 2 80056 52741
0 52743 5 1 1 52742
0 52744 7 1 2 86149 92366
0 52745 5 1 1 52744
0 52746 7 1 2 26800 52745
0 52747 5 1 1 52746
0 52748 7 1 2 59689 52747
0 52749 5 1 1 52748
0 52750 7 1 2 72262 96116
0 52751 5 1 1 52750
0 52752 7 1 2 52749 52751
0 52753 5 1 1 52752
0 52754 7 1 2 65516 52753
0 52755 5 1 1 52754
0 52756 7 1 2 52743 52755
0 52757 5 1 1 52756
0 52758 7 1 2 66772 52757
0 52759 5 1 1 52758
0 52760 7 1 2 92027 98429
0 52761 5 1 1 52760
0 52762 7 1 2 52759 52761
0 52763 5 1 1 52762
0 52764 7 1 2 65641 52763
0 52765 5 1 1 52764
0 52766 7 1 2 80058 98202
0 52767 5 1 1 52766
0 52768 7 1 2 92316 94882
0 52769 7 1 2 52767 52768
0 52770 5 1 1 52769
0 52771 7 1 2 52765 52770
0 52772 5 1 1 52771
0 52773 7 1 2 97013 52772
0 52774 5 1 1 52773
0 52775 7 1 2 52737 52774
0 52776 5 1 1 52775
0 52777 7 1 2 67768 52776
0 52778 5 1 1 52777
0 52779 7 2 2 65670 60820
0 52780 7 1 2 92303 95255
0 52781 7 1 2 98459 52780
0 52782 7 1 2 68958 90210
0 52783 7 1 2 92125 52782
0 52784 7 1 2 97357 52783
0 52785 7 1 2 52781 52784
0 52786 5 1 1 52785
0 52787 7 1 2 92132 44092
0 52788 5 3 1 52787
0 52789 7 2 2 67769 87871
0 52790 7 1 2 97776 98464
0 52791 7 1 2 98461 52790
0 52792 5 1 1 52791
0 52793 7 1 2 52786 52792
0 52794 5 1 1 52793
0 52795 7 1 2 97648 52794
0 52796 5 1 1 52795
0 52797 7 1 2 98412 98454
0 52798 5 1 1 52797
0 52799 7 1 2 95477 96050
0 52800 5 2 1 52799
0 52801 7 1 2 52798 98466
0 52802 5 1 1 52801
0 52803 7 1 2 91712 52802
0 52804 5 1 1 52803
0 52805 7 1 2 95676 96650
0 52806 5 1 1 52805
0 52807 7 1 2 52804 52806
0 52808 5 1 1 52807
0 52809 7 1 2 64067 52808
0 52810 5 1 1 52809
0 52811 7 1 2 73365 96882
0 52812 5 1 1 52811
0 52813 7 1 2 65517 98442
0 52814 5 1 1 52813
0 52815 7 1 2 52812 52814
0 52816 5 1 1 52815
0 52817 7 1 2 61137 98224
0 52818 7 1 2 52816 52817
0 52819 5 1 1 52818
0 52820 7 1 2 52810 52819
0 52821 5 1 1 52820
0 52822 7 1 2 97777 52821
0 52823 5 1 1 52822
0 52824 7 1 2 52796 52823
0 52825 7 1 2 52778 52824
0 52826 5 1 1 52825
0 52827 7 1 2 69028 52826
0 52828 5 1 1 52827
0 52829 7 3 2 68959 83890
0 52830 7 1 2 96239 98468
0 52831 5 1 1 52830
0 52832 7 1 2 90211 92737
0 52833 5 1 1 52832
0 52834 7 1 2 67770 96093
0 52835 5 1 1 52834
0 52836 7 1 2 52833 52835
0 52837 5 1 1 52836
0 52838 7 1 2 69607 52837
0 52839 5 1 1 52838
0 52840 7 1 2 15522 42242
0 52841 5 1 1 52840
0 52842 7 1 2 67771 52841
0 52843 5 1 1 52842
0 52844 7 1 2 52839 52843
0 52845 5 1 1 52844
0 52846 7 1 2 86307 52845
0 52847 5 1 1 52846
0 52848 7 1 2 52831 52847
0 52849 5 1 1 52848
0 52850 7 1 2 72263 52849
0 52851 5 1 1 52850
0 52852 7 1 2 84559 7829
0 52853 5 1 1 52852
0 52854 7 1 2 68550 52853
0 52855 5 1 1 52854
0 52856 7 1 2 70703 92152
0 52857 5 2 1 52856
0 52858 7 1 2 52855 98471
0 52859 5 1 1 52858
0 52860 7 1 2 68960 52859
0 52861 5 1 1 52860
0 52862 7 1 2 52851 52861
0 52863 5 1 1 52862
0 52864 7 1 2 91713 52863
0 52865 5 1 1 52864
0 52866 7 2 2 75718 78165
0 52867 7 1 2 72961 98473
0 52868 5 1 1 52867
0 52869 7 1 2 41392 52868
0 52870 5 1 1 52869
0 52871 7 1 2 59690 52870
0 52872 5 1 1 52871
0 52873 7 1 2 83590 82225
0 52874 7 1 2 95898 52873
0 52875 5 1 1 52874
0 52876 7 1 2 52872 52875
0 52877 5 1 1 52876
0 52878 7 1 2 68551 52877
0 52879 5 1 1 52878
0 52880 7 1 2 98472 52879
0 52881 5 1 1 52880
0 52882 7 1 2 61809 52881
0 52883 5 1 1 52882
0 52884 7 1 2 95985 52883
0 52885 5 1 1 52884
0 52886 7 1 2 68961 52885
0 52887 5 1 1 52886
0 52888 7 1 2 52865 52887
0 52889 5 1 1 52888
0 52890 7 1 2 86808 52889
0 52891 5 1 1 52890
0 52892 7 2 2 64068 73366
0 52893 7 1 2 61810 83510
0 52894 7 1 2 98475 52893
0 52895 5 2 1 52894
0 52896 7 1 2 63587 84616
0 52897 7 1 2 98469 52896
0 52898 5 1 1 52897
0 52899 7 1 2 98477 52898
0 52900 5 1 1 52899
0 52901 7 1 2 63862 52900
0 52902 5 1 1 52901
0 52903 7 1 2 81114 52544
0 52904 5 1 1 52903
0 52905 7 1 2 69608 52904
0 52906 5 1 1 52905
0 52907 7 1 2 81113 76879
0 52908 5 2 1 52907
0 52909 7 1 2 80964 82197
0 52910 5 1 1 52909
0 52911 7 1 2 98479 52910
0 52912 7 1 2 52906 52911
0 52913 5 1 1 52912
0 52914 7 1 2 77584 52913
0 52915 5 1 1 52914
0 52916 7 1 2 52902 52915
0 52917 5 1 1 52916
0 52918 7 1 2 72264 52917
0 52919 5 1 1 52918
0 52920 7 2 2 59691 97947
0 52921 7 1 2 92965 98452
0 52922 7 1 2 98481 52921
0 52923 5 1 1 52922
0 52924 7 1 2 52919 52923
0 52925 5 1 1 52924
0 52926 7 1 2 97801 52925
0 52927 5 1 1 52926
0 52928 7 1 2 66773 89226
0 52929 5 1 1 52928
0 52930 7 1 2 6943 72387
0 52931 5 2 1 52930
0 52932 7 1 2 52929 98483
0 52933 5 1 1 52932
0 52934 7 1 2 61372 95478
0 52935 7 1 2 92656 52934
0 52936 5 1 1 52935
0 52937 7 1 2 52933 52936
0 52938 5 1 1 52937
0 52939 7 1 2 63863 52938
0 52940 5 1 1 52939
0 52941 7 1 2 89995 96314
0 52942 5 1 1 52941
0 52943 7 1 2 52940 52942
0 52944 5 1 1 52943
0 52945 7 1 2 91714 52944
0 52946 5 1 1 52945
0 52947 7 1 2 92096 98484
0 52948 5 1 1 52947
0 52949 7 1 2 52946 52948
0 52950 5 1 1 52949
0 52951 7 1 2 85884 52950
0 52952 5 1 1 52951
0 52953 7 1 2 52927 52952
0 52954 5 1 1 52953
0 52955 7 1 2 61941 52954
0 52956 5 1 1 52955
0 52957 7 1 2 93983 98470
0 52958 5 1 1 52957
0 52959 7 1 2 98478 52958
0 52960 5 1 1 52959
0 52961 7 1 2 63864 52960
0 52962 5 1 1 52961
0 52963 7 1 2 90061 94353
0 52964 5 1 1 52963
0 52965 7 1 2 81115 52964
0 52966 5 1 1 52965
0 52967 7 1 2 69609 52966
0 52968 5 1 1 52967
0 52969 7 1 2 80965 96520
0 52970 5 1 1 52969
0 52971 7 1 2 98480 52970
0 52972 7 1 2 52968 52971
0 52973 5 1 1 52972
0 52974 7 1 2 77585 52973
0 52975 5 1 1 52974
0 52976 7 1 2 52962 52975
0 52977 5 1 1 52976
0 52978 7 1 2 60730 52977
0 52979 5 1 1 52978
0 52980 7 1 2 95055 98425
0 52981 7 1 2 98443 52980
0 52982 5 1 1 52981
0 52983 7 1 2 52979 52982
0 52984 5 1 1 52983
0 52985 7 1 2 72265 52984
0 52986 5 1 1 52985
0 52987 7 1 2 92482 95813
0 52988 7 1 2 98465 52987
0 52989 5 1 1 52988
0 52990 7 1 2 32525 52989
0 52991 5 1 1 52990
0 52992 7 1 2 83194 52991
0 52993 5 1 1 52992
0 52994 7 1 2 80542 84780
0 52995 7 1 2 96521 52994
0 52996 5 1 1 52995
0 52997 7 1 2 52993 52996
0 52998 5 1 1 52997
0 52999 7 1 2 61811 52998
0 53000 5 1 1 52999
0 53001 7 1 2 52986 53000
0 53002 5 1 1 53001
0 53003 7 1 2 90185 53002
0 53004 5 1 1 53003
0 53005 7 1 2 52956 53004
0 53006 7 1 2 52891 53005
0 53007 5 1 1 53006
0 53008 7 1 2 98246 53007
0 53009 5 1 1 53008
0 53010 7 1 2 52828 53009
0 53011 5 1 1 53010
0 53012 7 1 2 68156 53011
0 53013 5 1 1 53012
0 53014 7 1 2 70704 98406
0 53015 5 1 1 53014
0 53016 7 1 2 96019 97476
0 53017 7 1 2 96158 53016
0 53018 5 1 1 53017
0 53019 7 1 2 97944 98467
0 53020 5 1 1 53019
0 53021 7 1 2 91715 53020
0 53022 5 1 1 53021
0 53023 7 1 2 90591 95957
0 53024 5 1 1 53023
0 53025 7 1 2 53022 53024
0 53026 5 1 1 53025
0 53027 7 1 2 87194 53026
0 53028 5 1 1 53027
0 53029 7 1 2 53018 53028
0 53030 7 1 2 53015 53029
0 53031 5 1 1 53030
0 53032 7 1 2 98247 53031
0 53033 5 1 1 53032
0 53034 7 1 2 86456 97022
0 53035 7 1 2 97689 53034
0 53036 5 1 1 53035
0 53037 7 1 2 53033 53036
0 53038 5 1 1 53037
0 53039 7 1 2 73367 53038
0 53040 5 1 1 53039
0 53041 7 2 2 69610 72743
0 53042 7 2 2 92514 98237
0 53043 7 1 2 98485 98487
0 53044 5 1 1 53043
0 53045 7 1 2 87195 92126
0 53046 5 1 1 53045
0 53047 7 2 2 66587 92317
0 53048 5 1 1 98489
0 53049 7 1 2 61942 98490
0 53050 5 1 1 53049
0 53051 7 1 2 53046 53050
0 53052 5 1 1 53051
0 53053 7 1 2 98413 53052
0 53054 5 1 1 53053
0 53055 7 1 2 28374 96127
0 53056 5 1 1 53055
0 53057 7 1 2 65642 53056
0 53058 5 1 1 53057
0 53059 7 1 2 87020 87670
0 53060 5 1 1 53059
0 53061 7 1 2 53058 53060
0 53062 5 1 1 53061
0 53063 7 1 2 67135 92461
0 53064 7 1 2 53062 53063
0 53065 5 1 1 53064
0 53066 7 1 2 53054 53065
0 53067 5 1 1 53066
0 53068 7 1 2 68552 53067
0 53069 5 1 1 53068
0 53070 7 1 2 53044 53069
0 53071 5 1 1 53070
0 53072 7 1 2 67772 53071
0 53073 5 1 1 53072
0 53074 7 1 2 88620 98488
0 53075 5 1 1 53074
0 53076 7 1 2 53073 53075
0 53077 5 1 1 53076
0 53078 7 1 2 64170 53077
0 53079 5 1 1 53078
0 53080 7 1 2 96297 48193
0 53081 5 1 1 53080
0 53082 7 1 2 83691 53081
0 53083 5 1 1 53082
0 53084 7 1 2 63588 92086
0 53085 5 1 1 53084
0 53086 7 1 2 53083 53085
0 53087 5 1 1 53086
0 53088 7 1 2 68793 53087
0 53089 5 1 1 53088
0 53090 7 1 2 88264 98444
0 53091 5 1 1 53090
0 53092 7 1 2 53089 53091
0 53093 5 1 1 53092
0 53094 7 1 2 97744 53093
0 53095 5 1 1 53094
0 53096 7 1 2 50457 53095
0 53097 5 1 1 53096
0 53098 7 1 2 91716 53097
0 53099 5 1 1 53098
0 53100 7 1 2 83728 83195
0 53101 7 1 2 97755 53100
0 53102 5 1 1 53101
0 53103 7 1 2 53099 53102
0 53104 7 1 2 53079 53103
0 53105 5 1 1 53104
0 53106 7 1 2 95317 53105
0 53107 5 1 1 53106
0 53108 7 1 2 53040 53107
0 53109 5 1 1 53108
0 53110 7 1 2 68962 53109
0 53111 5 1 1 53110
0 53112 7 1 2 81617 98308
0 53113 5 1 1 53112
0 53114 7 1 2 96867 98331
0 53115 5 1 1 53114
0 53116 7 1 2 53113 53115
0 53117 5 1 1 53116
0 53118 7 1 2 77487 53117
0 53119 5 1 1 53118
0 53120 7 1 2 91984 97750
0 53121 5 1 1 53120
0 53122 7 1 2 53119 53121
0 53123 5 1 1 53122
0 53124 7 1 2 68553 53123
0 53125 5 1 1 53124
0 53126 7 1 2 90062 98205
0 53127 5 1 1 53126
0 53128 7 1 2 53125 53127
0 53129 5 1 1 53128
0 53130 7 1 2 68794 53129
0 53131 5 1 1 53130
0 53132 7 1 2 85017 98208
0 53133 5 1 1 53132
0 53134 7 2 2 68554 88713
0 53135 7 1 2 95113 98491
0 53136 5 1 1 53135
0 53137 7 2 2 70705 96315
0 53138 7 1 2 63589 97602
0 53139 7 1 2 98493 53138
0 53140 5 1 1 53139
0 53141 7 1 2 53136 53140
0 53142 5 1 1 53141
0 53143 7 1 2 88121 53142
0 53144 5 1 1 53143
0 53145 7 1 2 98462 98492
0 53146 5 1 1 53145
0 53147 7 1 2 96992 98494
0 53148 5 1 1 53147
0 53149 7 1 2 53146 53148
0 53150 5 1 1 53149
0 53151 7 1 2 86730 53150
0 53152 5 1 1 53151
0 53153 7 1 2 53144 53152
0 53154 5 1 1 53153
0 53155 7 1 2 63865 53154
0 53156 5 1 1 53155
0 53157 7 1 2 79451 91717
0 53158 7 1 2 98357 53157
0 53159 5 1 1 53158
0 53160 7 1 2 83891 96295
0 53161 7 1 2 96807 53160
0 53162 5 1 1 53161
0 53163 7 1 2 53159 53162
0 53164 5 1 1 53163
0 53165 7 1 2 88154 53164
0 53166 5 1 1 53165
0 53167 7 1 2 53156 53166
0 53168 5 1 1 53167
0 53169 7 1 2 69029 53168
0 53170 5 1 1 53169
0 53171 7 1 2 98358 98209
0 53172 5 1 1 53171
0 53173 7 1 2 53170 53172
0 53174 5 1 1 53173
0 53175 7 1 2 72266 53174
0 53176 5 1 1 53175
0 53177 7 1 2 53133 53176
0 53178 7 1 2 53131 53177
0 53179 5 1 1 53178
0 53180 7 1 2 97766 53179
0 53181 5 1 1 53180
0 53182 7 1 2 53111 53181
0 53183 7 1 2 53013 53182
0 53184 7 1 2 52700 53183
0 53185 7 1 2 52303 53184
0 53186 7 1 2 52042 53185
0 53187 7 1 2 51170 53186
0 53188 5 1 1 53187
0 53189 7 1 2 69141 53188
0 53190 5 1 1 53189
0 53191 7 2 2 89146 90159
0 53192 5 1 1 98495
0 53193 7 1 2 70867 53192
0 53194 5 1 1 53193
0 53195 7 1 2 97023 97702
0 53196 5 1 1 53195
0 53197 7 1 2 97018 53196
0 53198 5 1 1 53197
0 53199 7 1 2 67773 53198
0 53200 5 1 1 53199
0 53201 7 1 2 79639 97014
0 53202 7 1 2 98040 53201
0 53203 5 1 1 53202
0 53204 7 1 2 53200 53203
0 53205 5 1 1 53204
0 53206 7 1 2 68963 53205
0 53207 5 1 1 53206
0 53208 7 1 2 51949 53207
0 53209 5 1 1 53208
0 53210 7 1 2 53194 53209
0 53211 5 1 1 53210
0 53212 7 2 2 64171 95958
0 53213 7 1 2 86262 98497
0 53214 5 2 1 53213
0 53215 7 1 2 84686 96422
0 53216 7 1 2 97854 53215
0 53217 7 1 2 97948 53216
0 53218 5 1 1 53217
0 53219 7 1 2 67774 89180
0 53220 7 1 2 98431 53219
0 53221 5 1 1 53220
0 53222 7 1 2 53218 53221
0 53223 5 1 1 53222
0 53224 7 1 2 63590 53223
0 53225 5 1 1 53224
0 53226 7 1 2 98499 53225
0 53227 5 1 1 53226
0 53228 7 1 2 59692 53227
0 53229 5 1 1 53228
0 53230 7 2 2 95118 98498
0 53231 5 1 1 98501
0 53232 7 1 2 67775 98502
0 53233 5 1 1 53232
0 53234 7 1 2 77442 87081
0 53235 7 1 2 74977 53234
0 53236 7 1 2 98002 53235
0 53237 5 1 1 53236
0 53238 7 1 2 53233 53237
0 53239 5 1 1 53238
0 53240 7 1 2 62157 53239
0 53241 5 1 1 53240
0 53242 7 1 2 60956 83218
0 53243 7 1 2 86878 97890
0 53244 7 1 2 53242 53243
0 53245 5 1 1 53244
0 53246 7 1 2 53241 53245
0 53247 7 1 2 53229 53246
0 53248 5 1 1 53247
0 53249 7 1 2 64069 53248
0 53250 5 1 1 53249
0 53251 7 1 2 89181 89696
0 53252 5 1 1 53251
0 53253 7 2 2 82234 85491
0 53254 5 1 1 98503
0 53255 7 1 2 69730 98504
0 53256 5 1 1 53255
0 53257 7 1 2 53252 53256
0 53258 5 1 1 53257
0 53259 7 1 2 96620 53258
0 53260 5 1 1 53259
0 53261 7 2 2 69611 76653
0 53262 5 1 1 98505
0 53263 7 2 2 85855 92146
0 53264 5 1 1 98507
0 53265 7 1 2 98506 98508
0 53266 5 1 1 53265
0 53267 7 1 2 53260 53266
0 53268 5 1 1 53267
0 53269 7 1 2 59693 53268
0 53270 5 1 1 53269
0 53271 7 1 2 96621 97199
0 53272 5 1 1 53271
0 53273 7 1 2 53270 53272
0 53274 5 1 1 53273
0 53275 7 1 2 94772 53274
0 53276 5 1 1 53275
0 53277 7 1 2 53250 53276
0 53278 5 1 1 53277
0 53279 7 1 2 97802 53278
0 53280 5 1 1 53279
0 53281 7 1 2 69209 85376
0 53282 5 1 1 53281
0 53283 7 1 2 79297 53282
0 53284 5 1 1 53283
0 53285 7 1 2 76452 53284
0 53286 5 1 1 53285
0 53287 7 1 2 79459 53286
0 53288 5 1 1 53287
0 53289 7 1 2 68795 53288
0 53290 5 1 1 53289
0 53291 7 1 2 59398 84107
0 53292 5 2 1 53291
0 53293 7 1 2 83801 98509
0 53294 5 1 1 53293
0 53295 7 1 2 59694 53294
0 53296 5 1 1 53295
0 53297 7 1 2 78276 53296
0 53298 5 1 1 53297
0 53299 7 1 2 84528 53298
0 53300 5 1 1 53299
0 53301 7 1 2 53290 53300
0 53302 5 1 1 53301
0 53303 7 1 2 91718 53302
0 53304 5 1 1 53303
0 53305 7 1 2 90981 92097
0 53306 5 1 1 53305
0 53307 7 1 2 82425 92089
0 53308 5 1 1 53307
0 53309 7 1 2 63591 92462
0 53310 7 1 2 53308 53309
0 53311 5 1 1 53310
0 53312 7 1 2 53306 53311
0 53313 7 1 2 53304 53312
0 53314 5 1 1 53313
0 53315 7 1 2 66916 53314
0 53316 5 1 1 53315
0 53317 7 1 2 76329 98510
0 53318 5 1 1 53317
0 53319 7 1 2 91626 53318
0 53320 5 1 1 53319
0 53321 7 1 2 76214 82419
0 53322 5 1 1 53321
0 53323 7 1 2 78973 73591
0 53324 5 1 1 53323
0 53325 7 1 2 53322 53324
0 53326 7 1 2 53320 53325
0 53327 5 1 1 53326
0 53328 7 1 2 96200 53327
0 53329 5 1 1 53328
0 53330 7 1 2 81542 85714
0 53331 7 1 2 91413 53330
0 53332 5 1 1 53331
0 53333 7 1 2 53329 53332
0 53334 7 1 2 53316 53333
0 53335 5 1 1 53334
0 53336 7 1 2 70706 53335
0 53337 5 1 1 53336
0 53338 7 3 2 59695 89182
0 53339 5 1 1 98511
0 53340 7 1 2 92863 98512
0 53341 5 1 1 53340
0 53342 7 1 2 53341 51236
0 53343 5 1 1 53342
0 53344 7 1 2 66917 53343
0 53345 5 1 1 53344
0 53346 7 1 2 84914 93618
0 53347 5 1 1 53346
0 53348 7 1 2 53345 53347
0 53349 5 1 1 53348
0 53350 7 1 2 68157 53349
0 53351 5 1 1 53350
0 53352 7 1 2 86236 98280
0 53353 5 1 1 53352
0 53354 7 1 2 78874 79724
0 53355 7 1 2 80777 53354
0 53356 5 1 1 53355
0 53357 7 1 2 53353 53356
0 53358 5 1 1 53357
0 53359 7 1 2 74938 53358
0 53360 5 1 1 53359
0 53361 7 1 2 80339 93350
0 53362 5 1 1 53361
0 53363 7 1 2 73452 92644
0 53364 7 1 2 75891 53363
0 53365 7 1 2 95952 53364
0 53366 5 1 1 53365
0 53367 7 1 2 53362 53366
0 53368 5 1 1 53367
0 53369 7 1 2 85715 53368
0 53370 5 1 1 53369
0 53371 7 1 2 53360 53370
0 53372 7 1 2 53351 53371
0 53373 5 1 1 53372
0 53374 7 1 2 68555 53373
0 53375 5 1 1 53374
0 53376 7 1 2 76215 92801
0 53377 5 1 1 53376
0 53378 7 1 2 89147 92784
0 53379 5 1 1 53378
0 53380 7 1 2 53377 53379
0 53381 5 1 1 53380
0 53382 7 1 2 96714 53381
0 53383 5 1 1 53382
0 53384 7 1 2 53375 53383
0 53385 7 1 2 53337 53384
0 53386 5 1 1 53385
0 53387 7 1 2 96734 53386
0 53388 5 1 1 53387
0 53389 7 1 2 69210 83219
0 53390 5 1 1 53389
0 53391 7 1 2 83571 98513
0 53392 5 1 1 53391
0 53393 7 1 2 53390 53392
0 53394 5 1 1 53393
0 53395 7 1 2 68158 53394
0 53396 5 1 1 53395
0 53397 7 1 2 70499 93422
0 53398 5 1 1 53397
0 53399 7 1 2 53396 53398
0 53400 5 1 1 53399
0 53401 7 1 2 67776 53400
0 53402 5 1 1 53401
0 53403 7 1 2 73592 93423
0 53404 5 1 1 53403
0 53405 7 1 2 53402 53404
0 53406 5 1 1 53405
0 53407 7 1 2 97820 53406
0 53408 5 1 1 53407
0 53409 7 2 2 79725 89328
0 53410 7 1 2 69612 97522
0 53411 5 1 1 53410
0 53412 7 1 2 98086 53411
0 53413 5 1 1 53412
0 53414 7 1 2 59696 53413
0 53415 5 1 1 53414
0 53416 7 1 2 85012 53415
0 53417 5 1 1 53416
0 53418 7 1 2 98514 53417
0 53419 5 1 1 53418
0 53420 7 1 2 53408 53419
0 53421 5 1 1 53420
0 53422 7 1 2 64172 53421
0 53423 5 1 1 53422
0 53424 7 1 2 76216 96883
0 53425 5 1 1 53424
0 53426 7 1 2 65518 84915
0 53427 5 1 1 53426
0 53428 7 1 2 85049 91484
0 53429 5 1 1 53428
0 53430 7 1 2 53427 53429
0 53431 5 1 1 53430
0 53432 7 1 2 68556 53431
0 53433 5 1 1 53432
0 53434 7 1 2 53425 53433
0 53435 5 1 1 53434
0 53436 7 1 2 84450 94732
0 53437 7 1 2 53435 53436
0 53438 5 1 1 53437
0 53439 7 1 2 53423 53438
0 53440 5 1 1 53439
0 53441 7 1 2 60731 53440
0 53442 5 1 1 53441
0 53443 7 1 2 64070 53442
0 53444 7 1 2 53388 53443
0 53445 5 1 1 53444
0 53446 7 1 2 86327 98196
0 53447 5 1 1 53446
0 53448 7 1 2 80045 94733
0 53449 5 1 1 53448
0 53450 7 1 2 95708 96653
0 53451 7 1 2 98482 53450
0 53452 5 1 1 53451
0 53453 7 1 2 53449 53452
0 53454 5 1 1 53453
0 53455 7 1 2 60409 53454
0 53456 5 1 1 53455
0 53457 7 3 2 79687 97437
0 53458 7 1 2 70707 73198
0 53459 7 1 2 98516 53458
0 53460 5 1 1 53459
0 53461 7 1 2 50773 53460
0 53462 5 1 1 53461
0 53463 7 1 2 83196 53462
0 53464 5 1 1 53463
0 53465 7 1 2 49089 53464
0 53466 7 1 2 53456 53465
0 53467 5 1 1 53466
0 53468 7 1 2 69211 53467
0 53469 5 1 1 53468
0 53470 7 2 2 66918 98243
0 53471 7 1 2 82247 92834
0 53472 7 1 2 98519 53471
0 53473 5 1 1 53472
0 53474 7 1 2 53469 53473
0 53475 5 1 1 53474
0 53476 7 1 2 67777 53475
0 53477 5 1 1 53476
0 53478 7 1 2 53447 53477
0 53479 5 1 1 53478
0 53480 7 1 2 68159 53479
0 53481 5 1 1 53480
0 53482 7 2 2 86285 95709
0 53483 7 1 2 77042 98521
0 53484 5 1 1 53483
0 53485 7 1 2 51290 53484
0 53486 5 1 1 53485
0 53487 7 1 2 91719 53486
0 53488 5 1 1 53487
0 53489 7 1 2 96975 97861
0 53490 5 1 1 53489
0 53491 7 1 2 63866 53490
0 53492 7 1 2 53488 53491
0 53493 7 1 2 53481 53492
0 53494 5 1 1 53493
0 53495 7 1 2 93474 95666
0 53496 5 1 1 53495
0 53497 7 1 2 98192 53496
0 53498 5 1 1 53497
0 53499 7 1 2 89183 91627
0 53500 5 1 1 53499
0 53501 7 1 2 77447 53500
0 53502 5 2 1 53501
0 53503 7 1 2 97470 98298
0 53504 7 1 2 98523 53503
0 53505 5 1 1 53504
0 53506 7 1 2 53498 53505
0 53507 5 1 1 53506
0 53508 7 1 2 63592 53507
0 53509 5 1 1 53508
0 53510 7 2 2 79270 97526
0 53511 5 1 1 98525
0 53512 7 1 2 83808 96492
0 53513 5 1 1 53512
0 53514 7 1 2 53511 53513
0 53515 5 1 1 53514
0 53516 7 1 2 61943 53515
0 53517 5 1 1 53516
0 53518 7 1 2 83809 95753
0 53519 5 1 1 53518
0 53520 7 1 2 53517 53519
0 53521 5 1 1 53520
0 53522 7 1 2 95710 53521
0 53523 5 1 1 53522
0 53524 7 1 2 68796 53523
0 53525 7 1 2 53509 53524
0 53526 5 1 1 53525
0 53527 7 1 2 65643 53526
0 53528 7 1 2 53494 53527
0 53529 5 1 1 53528
0 53530 7 1 2 61812 98078
0 53531 5 1 1 53530
0 53532 7 1 2 82900 82235
0 53533 7 1 2 98486 53532
0 53534 5 1 1 53533
0 53535 7 1 2 53531 53534
0 53536 5 1 1 53535
0 53537 7 1 2 63867 53536
0 53538 5 1 1 53537
0 53539 7 1 2 83810 84369
0 53540 5 1 1 53539
0 53541 7 1 2 53538 53540
0 53542 5 1 1 53541
0 53543 7 1 2 91720 53542
0 53544 5 1 1 53543
0 53545 7 1 2 92098 98079
0 53546 5 1 1 53545
0 53547 7 1 2 68797 98526
0 53548 5 1 1 53547
0 53549 7 1 2 53546 53548
0 53550 7 1 2 53544 53549
0 53551 5 1 1 53550
0 53552 7 1 2 68557 53551
0 53553 5 1 1 53552
0 53554 7 1 2 83572 91985
0 53555 7 1 2 98524 53554
0 53556 5 1 1 53555
0 53557 7 1 2 53553 53556
0 53558 5 1 1 53557
0 53559 7 1 2 66919 53558
0 53560 5 1 1 53559
0 53561 7 1 2 68558 96146
0 53562 5 1 1 53561
0 53563 7 1 2 53560 53562
0 53564 5 1 1 53563
0 53565 7 1 2 95745 53564
0 53566 5 1 1 53565
0 53567 7 1 2 68964 53566
0 53568 7 1 2 53529 53567
0 53569 5 1 1 53568
0 53570 7 1 2 53445 53569
0 53571 5 1 1 53570
0 53572 7 1 2 53280 53571
0 53573 5 1 1 53572
0 53574 7 1 2 95318 53573
0 53575 5 1 1 53574
0 53576 7 1 2 53211 53575
0 53577 5 1 1 53576
0 53578 7 1 2 71257 53577
0 53579 5 1 1 53578
0 53580 7 1 2 71133 77054
0 53581 5 2 1 53580
0 53582 7 2 2 68965 97008
0 53583 5 1 1 98529
0 53584 7 1 2 70708 98530
0 53585 5 1 1 53584
0 53586 7 1 2 88156 97451
0 53587 7 1 2 89329 53586
0 53588 5 1 1 53587
0 53589 7 1 2 53585 53588
0 53590 5 1 1 53589
0 53591 7 1 2 97015 53590
0 53592 5 1 1 53591
0 53593 7 1 2 48663 53592
0 53594 5 1 1 53593
0 53595 7 1 2 76416 53594
0 53596 5 1 1 53595
0 53597 7 1 2 60732 94182
0 53598 5 1 1 53597
0 53599 7 1 2 96025 53598
0 53600 5 5 1 53599
0 53601 7 2 2 77586 98531
0 53602 7 1 2 88344 98536
0 53603 5 1 1 53602
0 53604 7 1 2 65644 98463
0 53605 5 2 1 53604
0 53606 7 1 2 98538 53048
0 53607 5 1 1 53606
0 53608 7 1 2 69323 85540
0 53609 7 1 2 53607 53608
0 53610 5 1 1 53609
0 53611 7 1 2 53603 53610
0 53612 5 1 1 53611
0 53613 7 1 2 68559 53612
0 53614 5 1 1 53613
0 53615 7 1 2 73963 90160
0 53616 7 1 2 98537 53615
0 53617 5 1 1 53616
0 53618 7 1 2 53614 53617
0 53619 5 1 1 53618
0 53620 7 1 2 64173 53619
0 53621 5 1 1 53620
0 53622 7 1 2 81224 85377
0 53623 5 1 1 53622
0 53624 7 1 2 85627 53623
0 53625 5 1 1 53624
0 53626 7 1 2 91888 97345
0 53627 7 1 2 94610 53626
0 53628 7 1 2 53625 53627
0 53629 5 1 1 53628
0 53630 7 1 2 61944 53629
0 53631 7 1 2 53621 53630
0 53632 5 1 1 53631
0 53633 7 1 2 89562 98458
0 53634 5 1 1 53633
0 53635 7 1 2 68798 96543
0 53636 7 1 2 53634 53635
0 53637 5 1 1 53636
0 53638 7 1 2 79640 78787
0 53639 7 1 2 97844 53638
0 53640 5 1 1 53639
0 53641 7 1 2 53637 53640
0 53642 5 1 1 53641
0 53643 7 1 2 68160 53642
0 53644 5 1 1 53643
0 53645 7 1 2 80705 98474
0 53646 7 1 2 98254 53645
0 53647 5 1 1 53646
0 53648 7 1 2 53644 53647
0 53649 5 1 1 53648
0 53650 7 1 2 67391 53649
0 53651 5 1 1 53650
0 53652 7 1 2 91721 98136
0 53653 5 2 1 53652
0 53654 7 1 2 86459 89780
0 53655 5 1 1 53654
0 53656 7 1 2 98540 53655
0 53657 5 1 1 53656
0 53658 7 1 2 70709 53657
0 53659 5 1 1 53658
0 53660 7 1 2 84308 96865
0 53661 5 1 1 53660
0 53662 7 1 2 53659 53661
0 53663 5 1 1 53662
0 53664 7 1 2 94652 53663
0 53665 5 1 1 53664
0 53666 7 1 2 53651 53665
0 53667 5 1 1 53666
0 53668 7 1 2 64071 53667
0 53669 5 1 1 53668
0 53670 7 1 2 8115 53254
0 53671 5 1 1 53670
0 53672 7 1 2 88022 98410
0 53673 7 1 2 53671 53672
0 53674 5 1 1 53673
0 53675 7 1 2 53669 53674
0 53676 5 1 1 53675
0 53677 7 1 2 69030 53676
0 53678 5 1 1 53677
0 53679 7 1 2 69324 97717
0 53680 7 1 2 89330 53679
0 53681 5 1 1 53680
0 53682 7 1 2 66920 53681
0 53683 7 1 2 53678 53682
0 53684 5 1 1 53683
0 53685 7 1 2 53632 53684
0 53686 5 1 1 53685
0 53687 7 1 2 92361 89821
0 53688 7 1 2 97728 53687
0 53689 7 1 2 97385 53688
0 53690 5 1 1 53689
0 53691 7 1 2 53686 53690
0 53692 5 1 1 53691
0 53693 7 1 2 95319 53692
0 53694 5 1 1 53693
0 53695 7 1 2 53596 53694
0 53696 5 1 1 53695
0 53697 7 1 2 98527 53696
0 53698 5 1 1 53697
0 53699 7 1 2 66774 98239
0 53700 5 1 1 53699
0 53701 7 1 2 87226 53700
0 53702 5 1 1 53701
0 53703 7 1 2 98344 53702
0 53704 5 1 1 53703
0 53705 7 1 2 79271 86809
0 53706 7 1 2 98346 53705
0 53707 5 1 1 53706
0 53708 7 1 2 53704 53707
0 53709 5 1 1 53708
0 53710 7 1 2 96985 53709
0 53711 5 1 1 53710
0 53712 7 2 2 64072 98170
0 53713 7 1 2 86308 98542
0 53714 5 1 1 53713
0 53715 7 1 2 86188 97586
0 53716 7 1 2 96884 53715
0 53717 5 1 1 53716
0 53718 7 1 2 53714 53717
0 53719 5 1 1 53718
0 53720 7 1 2 63868 95601
0 53721 7 1 2 53719 53720
0 53722 5 1 1 53721
0 53723 7 1 2 53711 53722
0 53724 5 1 1 53723
0 53725 7 1 2 67778 53724
0 53726 5 1 1 53725
0 53727 7 1 2 72267 97694
0 53728 5 1 1 53727
0 53729 7 1 2 67392 53728
0 53730 7 1 2 53726 53729
0 53731 5 1 1 53730
0 53732 7 1 2 95806 98180
0 53733 7 1 2 96722 53732
0 53734 5 1 1 53733
0 53735 7 1 2 88023 92851
0 53736 5 1 1 53735
0 53737 7 1 2 87872 87762
0 53738 7 1 2 97803 53737
0 53739 5 1 1 53738
0 53740 7 1 2 53736 53739
0 53741 5 1 1 53740
0 53742 7 1 2 63593 88200
0 53743 7 1 2 53741 53742
0 53744 5 1 1 53743
0 53745 7 1 2 53734 53744
0 53746 5 1 1 53745
0 53747 7 1 2 66921 53746
0 53748 5 1 1 53747
0 53749 7 1 2 75696 87151
0 53750 7 1 2 94200 53749
0 53751 7 1 2 96851 53750
0 53752 5 1 1 53751
0 53753 7 1 2 53748 53752
0 53754 5 1 1 53753
0 53755 7 1 2 69031 53754
0 53756 5 1 1 53755
0 53757 7 1 2 62395 53756
0 53758 5 1 1 53757
0 53759 7 1 2 60957 53758
0 53760 7 1 2 53731 53759
0 53761 5 1 1 53760
0 53762 7 2 2 96143 97858
0 53763 5 2 1 98544
0 53764 7 1 2 88138 96906
0 53765 5 1 1 53764
0 53766 7 1 2 98546 53765
0 53767 5 1 1 53766
0 53768 7 1 2 60410 53767
0 53769 5 1 1 53768
0 53770 7 1 2 79294 94222
0 53771 7 1 2 96069 53770
0 53772 5 1 1 53771
0 53773 7 1 2 53769 53772
0 53774 5 1 1 53773
0 53775 7 1 2 68966 53774
0 53776 5 1 1 53775
0 53777 7 1 2 85409 96651
0 53778 7 1 2 97959 53777
0 53779 5 1 1 53778
0 53780 7 1 2 53776 53779
0 53781 5 1 1 53780
0 53782 7 1 2 86731 53781
0 53783 5 1 1 53782
0 53784 7 1 2 83224 98543
0 53785 5 1 1 53784
0 53786 7 1 2 53783 53785
0 53787 5 1 1 53786
0 53788 7 1 2 72268 53787
0 53789 5 1 1 53788
0 53790 7 1 2 84219 92535
0 53791 5 1 1 53790
0 53792 7 1 2 98419 53791
0 53793 5 1 1 53792
0 53794 7 1 2 96928 97346
0 53795 7 1 2 53793 53794
0 53796 5 1 1 53795
0 53797 7 1 2 92548 97808
0 53798 5 1 1 53797
0 53799 7 1 2 72269 89944
0 53800 7 1 2 98234 53799
0 53801 5 1 1 53800
0 53802 7 1 2 53798 53801
0 53803 5 1 1 53802
0 53804 7 1 2 66775 53803
0 53805 5 1 1 53804
0 53806 7 1 2 92708 96680
0 53807 7 1 2 98181 53806
0 53808 5 1 1 53807
0 53809 7 1 2 53805 53808
0 53810 5 1 1 53809
0 53811 7 1 2 86810 53810
0 53812 5 1 1 53811
0 53813 7 1 2 53796 53812
0 53814 7 1 2 53789 53813
0 53815 7 1 2 53761 53814
0 53816 5 1 1 53815
0 53817 7 1 2 67136 53816
0 53818 5 1 1 53817
0 53819 7 1 2 76318 97495
0 53820 5 3 1 53819
0 53821 7 1 2 11555 98548
0 53822 5 1 1 53821
0 53823 7 1 2 98216 53822
0 53824 5 1 1 53823
0 53825 7 1 2 80669 96681
0 53826 7 1 2 97527 53825
0 53827 7 1 2 98532 53826
0 53828 5 1 1 53827
0 53829 7 1 2 53824 53828
0 53830 5 1 1 53829
0 53831 7 1 2 66922 53830
0 53832 5 1 1 53831
0 53833 7 1 2 92028 97379
0 53834 5 1 1 53833
0 53835 7 3 2 80543 94183
0 53836 7 1 2 83159 94987
0 53837 7 1 2 97528 53836
0 53838 7 1 2 98551 53837
0 53839 5 1 1 53838
0 53840 7 1 2 53834 53839
0 53841 5 1 1 53840
0 53842 7 1 2 97438 53841
0 53843 5 1 1 53842
0 53844 7 1 2 53832 53843
0 53845 7 1 2 53818 53844
0 53846 5 1 1 53845
0 53847 7 1 2 95320 53846
0 53848 5 1 1 53847
0 53849 7 1 2 8991 98549
0 53850 5 1 1 53849
0 53851 7 1 2 70710 53850
0 53852 5 1 1 53851
0 53853 7 1 2 86533 89725
0 53854 5 1 1 53853
0 53855 7 1 2 53852 53854
0 53856 5 1 1 53855
0 53857 7 1 2 97804 53856
0 53858 5 1 1 53857
0 53859 7 1 2 67393 97425
0 53860 7 1 2 87944 53859
0 53861 5 1 1 53860
0 53862 7 1 2 53858 53861
0 53863 5 1 1 53862
0 53864 7 1 2 66776 53863
0 53865 5 1 1 53864
0 53866 7 1 2 85546 98550
0 53867 5 1 1 53866
0 53868 7 2 2 70711 53867
0 53869 7 1 2 96993 98554
0 53870 5 1 1 53869
0 53871 7 1 2 85541 90144
0 53872 7 1 2 89607 53871
0 53873 5 1 1 53872
0 53874 7 1 2 53870 53873
0 53875 5 1 1 53874
0 53876 7 1 2 65645 53875
0 53877 5 1 1 53876
0 53878 7 1 2 53865 53877
0 53879 5 1 1 53878
0 53880 7 1 2 61945 53879
0 53881 5 1 1 53880
0 53882 7 1 2 95910 98555
0 53883 5 1 1 53882
0 53884 7 1 2 53881 53883
0 53885 5 1 1 53884
0 53886 7 1 2 64174 53885
0 53887 5 1 1 53886
0 53888 7 1 2 82080 97895
0 53889 5 1 1 53888
0 53890 7 2 2 94653 95907
0 53891 5 1 1 98556
0 53892 7 1 2 11587 39410
0 53893 5 1 1 53892
0 53894 7 1 2 65646 53893
0 53895 5 1 1 53894
0 53896 7 2 2 66588 88122
0 53897 7 1 2 87116 98558
0 53898 5 1 1 53897
0 53899 7 1 2 53895 53898
0 53900 5 1 1 53899
0 53901 7 1 2 82236 53900
0 53902 5 1 1 53901
0 53903 7 1 2 53891 53902
0 53904 5 1 1 53903
0 53905 7 1 2 78788 96336
0 53906 7 1 2 53904 53905
0 53907 5 1 1 53906
0 53908 7 1 2 53889 53907
0 53909 7 1 2 53887 53908
0 53910 5 1 1 53909
0 53911 7 1 2 95321 53910
0 53912 5 1 1 53911
0 53913 7 1 2 71398 97377
0 53914 7 1 2 98262 53913
0 53915 5 1 1 53914
0 53916 7 1 2 53912 53915
0 53917 5 1 1 53916
0 53918 7 1 2 71258 53917
0 53919 5 1 1 53918
0 53920 7 1 2 97812 98283
0 53921 5 1 1 53920
0 53922 7 1 2 48760 53921
0 53923 5 1 1 53922
0 53924 7 1 2 71259 53923
0 53925 5 1 1 53924
0 53926 7 1 2 97009 97791
0 53927 5 1 1 53926
0 53928 7 1 2 53925 53927
0 53929 5 1 1 53928
0 53930 7 1 2 95322 53929
0 53931 5 1 1 53930
0 53932 7 1 2 90129 92515
0 53933 7 1 2 92959 53932
0 53934 7 1 2 80785 86766
0 53935 7 1 2 95231 53934
0 53936 7 1 2 53933 53935
0 53937 5 1 1 53936
0 53938 7 1 2 53931 53937
0 53939 5 1 1 53938
0 53940 7 1 2 67137 53939
0 53941 5 1 1 53940
0 53942 7 1 2 93029 96899
0 53943 7 1 2 95264 95257
0 53944 7 1 2 95749 53943
0 53945 7 1 2 53942 53944
0 53946 5 1 1 53945
0 53947 7 1 2 53941 53946
0 53948 5 1 1 53947
0 53949 7 1 2 68967 53948
0 53950 5 1 1 53949
0 53951 7 1 2 42233 96270
0 53952 5 1 1 53951
0 53953 7 1 2 59986 53952
0 53954 5 1 1 53953
0 53955 7 1 2 83591 84288
0 53956 5 2 1 53955
0 53957 7 1 2 53954 98560
0 53958 5 1 1 53957
0 53959 7 1 2 92362 53958
0 53960 5 1 1 53959
0 53961 7 1 2 7673 96271
0 53962 5 1 1 53961
0 53963 7 1 2 59987 53962
0 53964 5 1 1 53963
0 53965 7 1 2 98561 53964
0 53966 5 1 1 53965
0 53967 7 1 2 97805 53966
0 53968 5 1 1 53967
0 53969 7 1 2 74191 98232
0 53970 5 1 1 53969
0 53971 7 1 2 53968 53970
0 53972 5 1 1 53971
0 53973 7 1 2 61946 53972
0 53974 5 1 1 53973
0 53975 7 1 2 53960 53974
0 53976 5 1 1 53975
0 53977 7 1 2 97471 53976
0 53978 5 1 1 53977
0 53979 7 1 2 67138 98362
0 53980 5 1 1 53979
0 53981 7 1 2 53978 53980
0 53982 5 1 1 53981
0 53983 7 1 2 68161 53982
0 53984 5 1 1 53983
0 53985 7 1 2 72270 98363
0 53986 5 1 1 53985
0 53987 7 2 2 79493 97656
0 53988 5 2 1 98562
0 53989 7 1 2 87763 91722
0 53990 7 1 2 98220 53989
0 53991 5 1 1 53990
0 53992 7 1 2 98564 53991
0 53993 5 1 1 53992
0 53994 7 1 2 72271 53993
0 53995 5 1 1 53994
0 53996 7 1 2 91398 97662
0 53997 5 1 1 53996
0 53998 7 1 2 53995 53997
0 53999 5 1 1 53998
0 54000 7 1 2 86811 53999
0 54001 5 1 1 54000
0 54002 7 1 2 53986 54001
0 54003 7 1 2 53984 54002
0 54004 5 1 1 54003
0 54005 7 1 2 81031 95323
0 54006 7 1 2 54004 54005
0 54007 5 1 1 54006
0 54008 7 1 2 53950 54007
0 54009 5 1 1 54008
0 54010 7 1 2 69325 54009
0 54011 5 1 1 54010
0 54012 7 1 2 89643 92563
0 54013 7 1 2 97458 98241
0 54014 7 1 2 54012 54013
0 54015 7 1 2 97454 54014
0 54016 5 1 1 54015
0 54017 7 1 2 54011 54016
0 54018 7 1 2 53919 54017
0 54019 7 1 2 53848 54018
0 54020 5 1 1 54019
0 54021 7 1 2 76286 54020
0 54022 5 1 1 54021
0 54023 7 1 2 97366 98197
0 54024 5 1 1 54023
0 54025 7 1 2 98176 54024
0 54026 5 1 1 54025
0 54027 7 1 2 67779 54026
0 54028 5 1 1 54027
0 54029 7 1 2 65519 96735
0 54030 7 1 2 95537 54029
0 54031 5 1 1 54030
0 54032 7 1 2 54028 54031
0 54033 5 1 1 54032
0 54034 7 1 2 66923 54033
0 54035 5 1 1 54034
0 54036 7 1 2 75530 97489
0 54037 5 1 1 54036
0 54038 7 1 2 97486 54037
0 54039 5 1 1 54038
0 54040 7 1 2 82237 97439
0 54041 7 1 2 54039 54040
0 54042 5 1 1 54041
0 54043 7 1 2 54035 54042
0 54044 5 1 1 54043
0 54045 7 1 2 68968 54044
0 54046 5 1 1 54045
0 54047 7 1 2 87554 98026
0 54048 5 1 1 54047
0 54049 7 1 2 49904 54048
0 54050 5 1 1 54049
0 54051 7 1 2 92029 54050
0 54052 5 1 1 54051
0 54053 7 1 2 54046 54052
0 54054 5 1 1 54053
0 54055 7 1 2 63869 54054
0 54056 5 1 1 54055
0 54057 7 1 2 69212 97917
0 54058 5 2 1 54057
0 54059 7 1 2 78882 97921
0 54060 5 1 1 54059
0 54061 7 1 2 98566 54060
0 54062 5 1 1 54061
0 54063 7 1 2 91723 54062
0 54064 5 1 1 54063
0 54065 7 2 2 63594 98302
0 54066 7 1 2 69213 98568
0 54067 5 2 1 54066
0 54068 7 1 2 90902 98041
0 54069 5 1 1 54068
0 54070 7 1 2 98570 54069
0 54071 5 1 1 54070
0 54072 7 1 2 61813 54071
0 54073 5 1 1 54072
0 54074 7 1 2 54064 54073
0 54075 5 1 1 54074
0 54076 7 1 2 77587 54075
0 54077 5 1 1 54076
0 54078 7 1 2 54056 54077
0 54079 5 1 1 54078
0 54080 7 1 2 95324 54079
0 54081 5 1 1 54080
0 54082 7 1 2 76319 98266
0 54083 5 1 1 54082
0 54084 7 1 2 54081 54083
0 54085 5 1 1 54084
0 54086 7 1 2 96007 54085
0 54087 5 1 1 54086
0 54088 7 1 2 54022 54087
0 54089 7 1 2 53698 54088
0 54090 7 1 2 53579 54089
0 54091 7 1 2 53190 54090
0 54092 7 1 2 50643 54091
0 54093 7 1 2 49455 54092
0 54094 7 1 2 70379 70905
0 54095 5 1 1 54094
0 54096 7 2 2 70868 88656
0 54097 5 1 1 98572
0 54098 7 1 2 59988 54097
0 54099 5 1 1 54098
0 54100 7 1 2 64592 95651
0 54101 7 1 2 54099 54100
0 54102 5 1 1 54101
0 54103 7 1 2 54095 54102
0 54104 5 1 1 54103
0 54105 7 1 2 64352 54104
0 54106 5 1 1 54105
0 54107 7 1 2 72782 71260
0 54108 7 1 2 82070 54107
0 54109 5 1 1 54108
0 54110 7 1 2 70906 54109
0 54111 5 1 1 54110
0 54112 7 1 2 70212 54111
0 54113 7 1 2 54106 54112
0 54114 5 1 1 54113
0 54115 7 1 2 62396 54114
0 54116 5 1 1 54115
0 54117 7 1 2 67139 96341
0 54118 5 1 1 54117
0 54119 7 1 2 65299 54118
0 54120 5 1 1 54119
0 54121 7 1 2 70213 90530
0 54122 5 1 1 54121
0 54123 7 1 2 95659 54122
0 54124 5 1 1 54123
0 54125 7 1 2 95657 54124
0 54126 7 1 2 54120 54125
0 54127 7 1 2 54116 54126
0 54128 5 1 1 54127
0 54129 7 1 2 61612 54128
0 54130 5 1 1 54129
0 54131 7 1 2 66589 71620
0 54132 7 1 2 82689 54131
0 54133 5 1 1 54132
0 54134 7 1 2 54130 54133
0 54135 5 1 1 54134
0 54136 7 1 2 67780 54135
0 54137 5 1 1 54136
0 54138 7 1 2 81243 90807
0 54139 5 1 1 54138
0 54140 7 1 2 20432 54139
0 54141 5 1 1 54140
0 54142 7 1 2 66590 54141
0 54143 5 1 1 54142
0 54144 7 1 2 96345 54143
0 54145 5 1 1 54144
0 54146 7 1 2 67140 54145
0 54147 5 1 1 54146
0 54148 7 1 2 72509 96348
0 54149 5 1 1 54148
0 54150 7 1 2 14818 54149
0 54151 5 1 1 54150
0 54152 7 1 2 62772 54151
0 54153 5 1 1 54152
0 54154 7 1 2 54147 54153
0 54155 7 1 2 54137 54154
0 54156 5 1 1 54155
0 54157 7 1 2 63207 54156
0 54158 5 1 1 54157
0 54159 7 1 2 67141 97506
0 54160 5 1 1 54159
0 54161 7 1 2 59697 91744
0 54162 5 1 1 54161
0 54163 7 1 2 60411 77507
0 54164 5 1 1 54163
0 54165 7 1 2 80765 87767
0 54166 7 1 2 54164 54165
0 54167 7 1 2 54162 54166
0 54168 7 1 2 54160 54167
0 54169 5 1 1 54168
0 54170 7 1 2 65520 54169
0 54171 5 1 1 54170
0 54172 7 1 2 96366 54171
0 54173 7 1 2 54158 54172
0 54174 5 1 1 54173
0 54175 7 1 2 68560 54174
0 54176 5 1 1 54175
0 54177 7 1 2 65300 97504
0 54178 5 1 1 54177
0 54179 7 1 2 83708 54178
0 54180 5 1 1 54179
0 54181 7 1 2 71462 97293
0 54182 5 1 1 54181
0 54183 7 1 2 84090 88427
0 54184 5 1 1 54183
0 54185 7 1 2 95594 54184
0 54186 5 1 1 54185
0 54187 7 1 2 63208 95588
0 54188 5 1 1 54187
0 54189 7 1 2 97034 54188
0 54190 7 1 2 54186 54189
0 54191 7 1 2 90526 97048
0 54192 5 1 1 54191
0 54193 7 1 2 62397 88363
0 54194 5 1 1 54193
0 54195 7 1 2 54192 54194
0 54196 7 1 2 54190 54195
0 54197 7 1 2 54182 54196
0 54198 5 1 1 54197
0 54199 7 1 2 66591 54198
0 54200 5 1 1 54199
0 54201 7 1 2 72510 77220
0 54202 5 1 1 54201
0 54203 7 1 2 65905 94687
0 54204 5 1 1 54203
0 54205 7 1 2 54202 54204
0 54206 5 1 1 54205
0 54207 7 1 2 88113 54206
0 54208 5 1 1 54207
0 54209 7 1 2 70898 54208
0 54210 5 1 1 54209
0 54211 7 1 2 79902 54210
0 54212 5 1 1 54211
0 54213 7 1 2 71526 54212
0 54214 7 1 2 54200 54213
0 54215 5 1 1 54214
0 54216 7 1 2 61613 77508
0 54217 5 1 1 54216
0 54218 7 1 2 60621 54217
0 54219 7 1 2 54215 54218
0 54220 5 1 1 54219
0 54221 7 1 2 54180 54220
0 54222 7 1 2 54176 54221
0 54223 5 1 1 54222
0 54224 7 1 2 68799 54223
0 54225 5 1 1 54224
0 54226 7 1 2 20414 54225
0 54227 5 1 1 54226
0 54228 7 1 2 61814 54227
0 54229 5 1 1 54228
0 54230 7 1 2 68800 95538
0 54231 5 1 1 54230
0 54232 7 1 2 95962 54231
0 54233 5 1 1 54232
0 54234 7 1 2 96389 54233
0 54235 5 1 1 54234
0 54236 7 1 2 84529 95134
0 54237 5 1 1 54236
0 54238 7 1 2 63209 54237
0 54239 5 1 1 54238
0 54240 7 1 2 70712 93795
0 54241 7 1 2 54239 54240
0 54242 5 1 1 54241
0 54243 7 1 2 54235 54242
0 54244 5 1 1 54243
0 54245 7 1 2 72272 54244
0 54246 5 1 1 54245
0 54247 7 1 2 89080 97962
0 54248 5 1 1 54247
0 54249 7 1 2 82936 92445
0 54250 5 1 1 54249
0 54251 7 1 2 54248 54250
0 54252 5 1 1 54251
0 54253 7 1 2 59698 54252
0 54254 5 1 1 54253
0 54255 7 1 2 67142 84451
0 54256 7 1 2 96783 54255
0 54257 5 1 1 54256
0 54258 7 1 2 54254 54257
0 54259 5 1 1 54258
0 54260 7 1 2 69326 54259
0 54261 5 1 1 54260
0 54262 7 1 2 68801 82198
0 54263 5 1 1 54262
0 54264 7 1 2 32864 54263
0 54265 5 1 1 54264
0 54266 7 1 2 76320 54265
0 54267 5 1 1 54266
0 54268 7 1 2 96106 54267
0 54269 5 1 1 54268
0 54270 7 1 2 68162 54269
0 54271 5 1 1 54270
0 54272 7 1 2 54261 54271
0 54273 7 1 2 54246 54272
0 54274 5 1 1 54273
0 54275 7 1 2 91724 54274
0 54276 5 1 1 54275
0 54277 7 1 2 80970 92485
0 54278 5 1 1 54277
0 54279 7 1 2 69214 54278
0 54280 5 1 1 54279
0 54281 7 1 2 73368 95934
0 54282 5 1 1 54281
0 54283 7 1 2 54280 54282
0 54284 5 1 1 54283
0 54285 7 1 2 84452 54284
0 54286 5 1 1 54285
0 54287 7 1 2 84372 54286
0 54288 5 1 1 54287
0 54289 7 1 2 90186 54288
0 54290 5 1 1 54289
0 54291 7 1 2 66924 54290
0 54292 7 1 2 54276 54291
0 54293 7 1 2 54229 54292
0 54294 5 1 1 54293
0 54295 7 1 2 88395 97056
0 54296 5 1 1 54295
0 54297 7 1 2 63210 86953
0 54298 5 1 1 54297
0 54299 7 1 2 70214 54298
0 54300 5 1 1 54299
0 54301 7 1 2 64353 54300
0 54302 5 1 1 54301
0 54303 7 1 2 79090 54302
0 54304 5 1 1 54303
0 54305 7 1 2 69711 54304
0 54306 5 1 1 54305
0 54307 7 1 2 91285 54306
0 54308 5 1 1 54307
0 54309 7 1 2 62158 54308
0 54310 5 1 1 54309
0 54311 7 1 2 54296 54310
0 54312 5 1 1 54311
0 54313 7 1 2 62773 54312
0 54314 5 1 1 54313
0 54315 7 1 2 71328 91280
0 54316 5 1 1 54315
0 54317 7 1 2 3887 54316
0 54318 5 1 1 54317
0 54319 7 1 2 82580 54318
0 54320 5 1 1 54319
0 54321 7 1 2 71134 94902
0 54322 5 1 1 54321
0 54323 7 1 2 70088 73216
0 54324 5 1 1 54323
0 54325 7 1 2 84662 54324
0 54326 7 1 2 54322 54325
0 54327 5 1 1 54326
0 54328 7 1 2 74512 54327
0 54329 5 1 1 54328
0 54330 7 1 2 70089 88937
0 54331 5 1 1 54330
0 54332 7 1 2 91130 88633
0 54333 7 1 2 88527 54332
0 54334 5 1 1 54333
0 54335 7 1 2 54331 54334
0 54336 7 1 2 54329 54335
0 54337 7 1 2 54320 54336
0 54338 7 1 2 54314 54337
0 54339 5 1 1 54338
0 54340 7 1 2 61815 54339
0 54341 5 1 1 54340
0 54342 7 1 2 80470 86865
0 54343 5 1 1 54342
0 54344 7 1 2 97083 54343
0 54345 5 1 1 54344
0 54346 7 1 2 65037 54345
0 54347 5 1 1 54346
0 54348 7 1 2 79365 90992
0 54349 5 1 1 54348
0 54350 7 1 2 54347 54349
0 54351 5 1 1 54350
0 54352 7 1 2 69712 54351
0 54353 5 1 1 54352
0 54354 7 1 2 62774 91042
0 54355 5 1 1 54354
0 54356 7 1 2 69996 85607
0 54357 5 1 1 54356
0 54358 7 1 2 70090 73051
0 54359 5 1 1 54358
0 54360 7 1 2 91134 54359
0 54361 7 1 2 54357 54360
0 54362 7 1 2 54355 54361
0 54363 5 1 1 54362
0 54364 7 1 2 61816 54363
0 54365 5 1 1 54364
0 54366 7 1 2 54353 54365
0 54367 5 1 1 54366
0 54368 7 1 2 71839 54367
0 54369 5 1 1 54368
0 54370 7 1 2 78350 88897
0 54371 5 1 1 54370
0 54372 7 1 2 77509 54371
0 54373 5 1 1 54372
0 54374 7 1 2 70869 54373
0 54375 5 1 1 54374
0 54376 7 1 2 69376 77488
0 54377 5 2 1 54376
0 54378 7 1 2 70215 98574
0 54379 5 1 1 54378
0 54380 7 1 2 62398 54379
0 54381 5 1 1 54380
0 54382 7 1 2 76862 97324
0 54383 5 1 1 54382
0 54384 7 1 2 65746 54383
0 54385 5 1 1 54384
0 54386 7 1 2 54381 54385
0 54387 5 1 1 54386
0 54388 7 1 2 64354 54387
0 54389 5 1 1 54388
0 54390 7 1 2 73052 97322
0 54391 5 1 1 54390
0 54392 7 1 2 70091 15736
0 54393 5 1 1 54392
0 54394 7 1 2 54391 54393
0 54395 7 1 2 54389 54394
0 54396 7 1 2 54375 54395
0 54397 5 1 1 54396
0 54398 7 1 2 61817 54397
0 54399 5 1 1 54398
0 54400 7 1 2 85315 97530
0 54401 5 1 1 54400
0 54402 7 1 2 54399 54401
0 54403 7 1 2 54369 54402
0 54404 5 1 1 54403
0 54405 7 1 2 72388 54404
0 54406 5 1 1 54405
0 54407 7 1 2 54341 54406
0 54408 5 1 1 54407
0 54409 7 1 2 91875 54408
0 54410 5 1 1 54409
0 54411 7 1 2 70345 86008
0 54412 5 1 1 54411
0 54413 7 1 2 26243 54412
0 54414 5 1 1 54413
0 54415 7 1 2 64355 54414
0 54416 5 1 1 54415
0 54417 7 1 2 69377 86009
0 54418 5 1 1 54417
0 54419 7 1 2 54416 54418
0 54420 5 1 1 54419
0 54421 7 1 2 69280 54420
0 54422 5 1 1 54421
0 54423 7 1 2 65521 73217
0 54424 5 1 1 54423
0 54425 7 1 2 86016 54424
0 54426 5 1 1 54425
0 54427 7 1 2 69076 54426
0 54428 5 1 1 54427
0 54429 7 1 2 54422 54428
0 54430 5 1 1 54429
0 54431 7 1 2 64593 54430
0 54432 5 1 1 54431
0 54433 7 1 2 71511 75800
0 54434 5 1 1 54433
0 54435 7 1 2 65522 54434
0 54436 5 1 1 54435
0 54437 7 1 2 77876 78580
0 54438 7 1 2 95793 54437
0 54439 5 1 1 54438
0 54440 7 1 2 54436 54439
0 54441 5 1 1 54440
0 54442 7 1 2 62775 54441
0 54443 5 1 1 54442
0 54444 7 1 2 77081 86377
0 54445 7 1 2 78419 54444
0 54446 5 1 1 54445
0 54447 7 1 2 60622 54446
0 54448 5 1 1 54447
0 54449 7 1 2 63211 54448
0 54450 5 1 1 54449
0 54451 7 1 2 78021 76887
0 54452 7 1 2 95272 54451
0 54453 5 1 1 54452
0 54454 7 1 2 71261 89203
0 54455 5 1 1 54454
0 54456 7 1 2 78581 93416
0 54457 5 1 1 54456
0 54458 7 1 2 60623 54457
0 54459 5 1 1 54458
0 54460 7 1 2 54455 54459
0 54461 5 1 1 54460
0 54462 7 1 2 93597 54461
0 54463 7 1 2 54453 54462
0 54464 7 1 2 54450 54463
0 54465 7 1 2 54443 54464
0 54466 7 1 2 54432 54465
0 54467 5 1 1 54466
0 54468 7 1 2 61818 54467
0 54469 5 1 1 54468
0 54470 7 1 2 65523 90314
0 54471 5 1 1 54470
0 54472 7 1 2 79349 97320
0 54473 5 1 1 54472
0 54474 7 1 2 54471 54473
0 54475 5 1 1 54474
0 54476 7 1 2 61819 54475
0 54477 5 1 1 54476
0 54478 7 1 2 85410 86542
0 54479 5 1 1 54478
0 54480 7 1 2 77518 94913
0 54481 5 1 1 54480
0 54482 7 1 2 54479 54481
0 54483 5 1 1 54482
0 54484 7 1 2 69713 54483
0 54485 5 1 1 54484
0 54486 7 1 2 65524 73053
0 54487 5 1 1 54486
0 54488 7 1 2 69997 77355
0 54489 7 1 2 85566 54488
0 54490 5 1 1 54489
0 54491 7 1 2 54487 54490
0 54492 5 1 1 54491
0 54493 7 1 2 61820 54492
0 54494 5 1 1 54493
0 54495 7 1 2 54485 54494
0 54496 5 1 1 54495
0 54497 7 1 2 71840 54496
0 54498 5 1 1 54497
0 54499 7 1 2 84386 88324
0 54500 7 1 2 92793 54499
0 54501 5 1 1 54500
0 54502 7 1 2 54498 54501
0 54503 7 1 2 54477 54502
0 54504 5 1 1 54503
0 54505 7 1 2 72389 54504
0 54506 5 1 1 54505
0 54507 7 1 2 54469 54506
0 54508 5 1 1 54507
0 54509 7 1 2 75638 54508
0 54510 5 1 1 54509
0 54511 7 1 2 44499 54510
0 54512 7 1 2 54410 54511
0 54513 5 1 1 54512
0 54514 7 1 2 63870 54513
0 54515 5 1 1 54514
0 54516 7 1 2 62399 80213
0 54517 5 1 1 54516
0 54518 7 1 2 70216 94805
0 54519 7 1 2 54517 54518
0 54520 5 1 1 54519
0 54521 7 1 2 74320 54520
0 54522 5 1 1 54521
0 54523 7 1 2 80305 77201
0 54524 7 1 2 74661 54523
0 54525 5 1 1 54524
0 54526 7 1 2 54522 54525
0 54527 5 1 1 54526
0 54528 7 1 2 63212 54527
0 54529 5 1 1 54528
0 54530 7 1 2 66592 95140
0 54531 5 1 1 54530
0 54532 7 1 2 54529 54531
0 54533 5 1 1 54532
0 54534 7 1 2 71935 54533
0 54535 5 1 1 54534
0 54536 7 1 2 91242 95767
0 54537 5 1 1 54536
0 54538 7 1 2 69862 88370
0 54539 5 1 1 54538
0 54540 7 1 2 80700 91228
0 54541 5 1 1 54540
0 54542 7 1 2 74133 95769
0 54543 5 1 1 54542
0 54544 7 1 2 54541 54543
0 54545 7 1 2 54539 54544
0 54546 7 1 2 54537 54545
0 54547 5 1 1 54546
0 54548 7 1 2 63213 54547
0 54549 5 1 1 54548
0 54550 7 1 2 59989 93337
0 54551 5 1 1 54550
0 54552 7 1 2 77871 73171
0 54553 7 1 2 54551 54552
0 54554 5 1 1 54553
0 54555 7 1 2 91229 95277
0 54556 5 1 1 54555
0 54557 7 1 2 54554 54556
0 54558 7 1 2 54549 54557
0 54559 5 1 1 54558
0 54560 7 1 2 66593 54559
0 54561 5 1 1 54560
0 54562 7 1 2 69378 81576
0 54563 5 1 1 54562
0 54564 7 1 2 77014 54563
0 54565 5 1 1 54564
0 54566 7 1 2 64356 54565
0 54567 5 1 1 54566
0 54568 7 1 2 64822 70358
0 54569 5 1 1 54568
0 54570 7 1 2 54567 54569
0 54571 5 1 1 54570
0 54572 7 1 2 64594 54571
0 54573 5 1 1 54572
0 54574 7 1 2 95790 54573
0 54575 5 1 1 54574
0 54576 7 1 2 93813 54575
0 54577 5 1 1 54576
0 54578 7 1 2 54561 54577
0 54579 7 1 2 54535 54578
0 54580 5 1 1 54579
0 54581 7 1 2 65301 54580
0 54582 5 1 1 54581
0 54583 7 1 2 66080 82296
0 54584 5 1 1 54583
0 54585 7 1 2 90749 54584
0 54586 5 1 1 54585
0 54587 7 1 2 65906 54586
0 54588 5 1 1 54587
0 54589 7 1 2 95819 54588
0 54590 5 1 1 54589
0 54591 7 1 2 64595 54590
0 54592 5 1 1 54591
0 54593 7 1 2 62776 89230
0 54594 5 1 1 54593
0 54595 7 1 2 70963 54594
0 54596 7 1 2 54592 54595
0 54597 5 1 1 54596
0 54598 7 1 2 70965 87485
0 54599 7 1 2 54597 54598
0 54600 5 1 1 54599
0 54601 7 1 2 54582 54600
0 54602 5 1 1 54601
0 54603 7 1 2 84204 54602
0 54604 5 1 1 54603
0 54605 7 1 2 87482 88419
0 54606 5 1 1 54605
0 54607 7 1 2 72511 86938
0 54608 5 1 1 54607
0 54609 7 1 2 54606 54608
0 54610 5 1 1 54609
0 54611 7 1 2 71841 54610
0 54612 5 1 1 54611
0 54613 7 1 2 91044 54612
0 54614 5 1 1 54613
0 54615 7 1 2 62400 54614
0 54616 5 1 1 54615
0 54617 7 1 2 62777 95358
0 54618 5 1 1 54617
0 54619 7 1 2 72027 84658
0 54620 5 1 1 54619
0 54621 7 1 2 54618 54620
0 54622 5 1 1 54621
0 54623 7 1 2 64357 54622
0 54624 5 1 1 54623
0 54625 7 1 2 54616 54624
0 54626 5 1 1 54625
0 54627 7 1 2 85921 54626
0 54628 5 1 1 54627
0 54629 7 1 2 88164 91326
0 54630 5 1 1 54629
0 54631 7 1 2 62401 71587
0 54632 5 1 1 54631
0 54633 7 1 2 63214 86604
0 54634 5 1 1 54633
0 54635 7 1 2 54632 54634
0 54636 5 1 1 54635
0 54637 7 1 2 85922 54636
0 54638 5 1 1 54637
0 54639 7 1 2 15754 54638
0 54640 5 1 1 54639
0 54641 7 1 2 78672 54640
0 54642 5 1 1 54641
0 54643 7 1 2 54630 54642
0 54644 7 1 2 54628 54643
0 54645 5 1 1 54644
0 54646 7 1 2 70346 54645
0 54647 5 1 1 54646
0 54648 7 1 2 91388 97316
0 54649 5 1 1 54648
0 54650 7 1 2 72390 54649
0 54651 5 1 1 54650
0 54652 7 1 2 71135 75042
0 54653 5 1 1 54652
0 54654 7 1 2 81927 54653
0 54655 7 1 2 54651 54654
0 54656 5 1 1 54655
0 54657 7 1 2 62778 54656
0 54658 5 1 1 54657
0 54659 7 1 2 70870 91465
0 54660 5 1 1 54659
0 54661 7 1 2 70217 54660
0 54662 7 1 2 54658 54661
0 54663 5 1 1 54662
0 54664 7 1 2 63215 54663
0 54665 5 1 1 54664
0 54666 7 1 2 64358 90375
0 54667 5 1 1 54666
0 54668 7 1 2 68163 54667
0 54669 5 1 1 54668
0 54670 7 1 2 64823 54669
0 54671 5 1 1 54670
0 54672 7 1 2 91459 54671
0 54673 5 1 1 54672
0 54674 7 1 2 70871 54673
0 54675 5 1 1 54674
0 54676 7 1 2 83870 90376
0 54677 5 1 1 54676
0 54678 7 1 2 54675 54677
0 54679 5 1 1 54678
0 54680 7 1 2 82793 54679
0 54681 5 1 1 54680
0 54682 7 1 2 69379 91446
0 54683 5 1 1 54682
0 54684 7 1 2 81704 54683
0 54685 5 1 1 54684
0 54686 7 1 2 63216 54685
0 54687 5 1 1 54686
0 54688 7 1 2 73275 88959
0 54689 5 1 1 54688
0 54690 7 1 2 89052 54689
0 54691 5 1 1 54690
0 54692 7 1 2 88516 95757
0 54693 5 1 1 54692
0 54694 7 1 2 54691 54693
0 54695 5 1 1 54694
0 54696 7 1 2 70872 54695
0 54697 5 1 1 54696
0 54698 7 1 2 54687 54697
0 54699 5 1 1 54698
0 54700 7 1 2 69281 54699
0 54701 5 1 1 54700
0 54702 7 1 2 62779 91103
0 54703 5 1 1 54702
0 54704 7 1 2 82463 78450
0 54705 5 1 1 54704
0 54706 7 1 2 65302 54705
0 54707 5 1 1 54706
0 54708 7 1 2 54703 54707
0 54709 7 1 2 54701 54708
0 54710 7 1 2 54681 54709
0 54711 7 1 2 54665 54710
0 54712 5 1 1 54711
0 54713 7 1 2 85923 54712
0 54714 5 1 1 54713
0 54715 7 2 2 59990 95479
0 54716 5 1 1 98576
0 54717 7 1 2 61614 76541
0 54718 5 1 1 54717
0 54719 7 1 2 68561 81476
0 54720 5 1 1 54719
0 54721 7 1 2 54718 54720
0 54722 5 1 1 54721
0 54723 7 1 2 60958 54722
0 54724 5 1 1 54723
0 54725 7 1 2 54716 54724
0 54726 5 1 1 54725
0 54727 7 1 2 65525 54726
0 54728 5 1 1 54727
0 54729 7 1 2 85057 89062
0 54730 5 1 1 54729
0 54731 7 1 2 16409 54730
0 54732 5 1 1 54731
0 54733 7 1 2 59699 54732
0 54734 5 1 1 54733
0 54735 7 1 2 91350 92794
0 54736 7 1 2 95281 54735
0 54737 5 1 1 54736
0 54738 7 1 2 54734 54737
0 54739 7 1 2 54728 54738
0 54740 5 1 1 54739
0 54741 7 1 2 68164 54740
0 54742 5 1 1 54741
0 54743 7 1 2 70411 78673
0 54744 5 1 1 54743
0 54745 7 1 2 70500 82068
0 54746 5 1 1 54745
0 54747 7 1 2 54744 54746
0 54748 5 1 1 54747
0 54749 7 1 2 64359 54748
0 54750 5 1 1 54749
0 54751 7 1 2 80495 91468
0 54752 5 1 1 54751
0 54753 7 1 2 62780 54752
0 54754 5 1 1 54753
0 54755 7 1 2 72391 14514
0 54756 5 1 1 54755
0 54757 7 1 2 71262 54756
0 54758 7 1 2 54754 54757
0 54759 7 1 2 54750 54758
0 54760 5 1 1 54759
0 54761 7 1 2 79822 87832
0 54762 7 1 2 80288 54761
0 54763 7 1 2 54760 54762
0 54764 5 1 1 54763
0 54765 7 1 2 60624 81800
0 54766 5 1 1 54765
0 54767 7 1 2 68562 93259
0 54768 5 1 1 54767
0 54769 7 1 2 54766 54768
0 54770 5 1 1 54769
0 54771 7 1 2 66594 54770
0 54772 5 1 1 54771
0 54773 7 1 2 65526 90700
0 54774 5 1 1 54773
0 54775 7 1 2 63871 54774
0 54776 7 1 2 54772 54775
0 54777 7 1 2 54764 54776
0 54778 7 1 2 54742 54777
0 54779 7 1 2 54714 54778
0 54780 7 1 2 54647 54779
0 54781 5 1 1 54780
0 54782 7 1 2 82811 90539
0 54783 5 1 1 54782
0 54784 7 1 2 69863 82471
0 54785 5 1 1 54784
0 54786 7 1 2 72273 54785
0 54787 5 1 1 54786
0 54788 7 1 2 91435 88387
0 54789 7 1 2 54787 54788
0 54790 5 1 1 54789
0 54791 7 1 2 90850 54790
0 54792 5 1 1 54791
0 54793 7 1 2 64596 54792
0 54794 5 1 1 54793
0 54795 7 1 2 73218 91208
0 54796 5 1 1 54795
0 54797 7 1 2 69147 90442
0 54798 5 1 1 54797
0 54799 7 1 2 64360 54798
0 54800 5 1 1 54799
0 54801 7 1 2 91598 97217
0 54802 7 1 2 54800 54801
0 54803 5 1 1 54802
0 54804 7 1 2 64824 54803
0 54805 5 1 1 54804
0 54806 7 1 2 54796 54805
0 54807 7 1 2 54794 54806
0 54808 5 1 1 54807
0 54809 7 1 2 63217 54808
0 54810 5 1 1 54809
0 54811 7 1 2 54783 54810
0 54812 5 1 1 54811
0 54813 7 1 2 97267 54812
0 54814 5 1 1 54813
0 54815 7 1 2 72618 88475
0 54816 5 1 1 54815
0 54817 7 1 2 95366 54816
0 54818 5 1 1 54817
0 54819 7 1 2 65527 54818
0 54820 5 1 1 54819
0 54821 7 1 2 73253 86010
0 54822 5 1 1 54821
0 54823 7 1 2 60625 54822
0 54824 5 1 1 54823
0 54825 7 1 2 62781 96460
0 54826 7 1 2 54824 54825
0 54827 5 1 1 54826
0 54828 7 1 2 54820 54827
0 54829 5 1 1 54828
0 54830 7 1 2 75639 54829
0 54831 5 1 1 54830
0 54832 7 1 2 79151 72415
0 54833 5 1 1 54832
0 54834 7 1 2 95598 54833
0 54835 5 1 1 54834
0 54836 7 1 2 76921 88814
0 54837 5 1 1 54836
0 54838 7 1 2 54835 54837
0 54839 5 1 1 54838
0 54840 7 1 2 70873 54839
0 54841 5 1 1 54840
0 54842 7 1 2 91281 95552
0 54843 5 1 1 54842
0 54844 7 1 2 64597 90507
0 54845 7 1 2 88476 54844
0 54846 5 1 1 54845
0 54847 7 1 2 68165 90873
0 54848 7 1 2 54846 54847
0 54849 5 1 1 54848
0 54850 7 1 2 70092 54849
0 54851 5 1 1 54850
0 54852 7 1 2 54843 54851
0 54853 7 1 2 54841 54852
0 54854 5 1 1 54853
0 54855 7 1 2 91876 54854
0 54856 5 1 1 54855
0 54857 7 1 2 54831 54856
0 54858 5 1 1 54857
0 54859 7 1 2 69282 54858
0 54860 5 1 1 54859
0 54861 7 1 2 63218 94968
0 54862 5 1 1 54861
0 54863 7 1 2 70093 94980
0 54864 5 1 1 54863
0 54865 7 1 2 54862 54864
0 54866 5 1 1 54865
0 54867 7 1 2 91877 54866
0 54868 5 1 1 54867
0 54869 7 1 2 89523 94982
0 54870 5 1 1 54869
0 54871 7 1 2 65528 54870
0 54872 5 1 1 54871
0 54873 7 1 2 70501 91001
0 54874 7 1 2 94049 54873
0 54875 5 1 1 54874
0 54876 7 1 2 54872 54875
0 54877 5 1 1 54876
0 54878 7 1 2 75640 54877
0 54879 5 1 1 54878
0 54880 7 1 2 54868 54879
0 54881 5 1 1 54880
0 54882 7 1 2 71936 54881
0 54883 5 1 1 54882
0 54884 7 1 2 90865 93150
0 54885 5 1 1 54884
0 54886 7 1 2 64361 54885
0 54887 5 1 1 54886
0 54888 7 1 2 69077 73297
0 54889 5 1 1 54888
0 54890 7 1 2 54887 54889
0 54891 5 1 1 54890
0 54892 7 1 2 97261 54891
0 54893 5 1 1 54892
0 54894 7 1 2 71471 83971
0 54895 5 1 1 54894
0 54896 7 1 2 97285 54895
0 54897 5 1 1 54896
0 54898 7 1 2 54893 54897
0 54899 5 1 1 54898
0 54900 7 1 2 73800 54899
0 54901 5 1 1 54900
0 54902 7 1 2 95928 96257
0 54903 5 1 1 54902
0 54904 7 1 2 65529 95923
0 54905 7 1 2 54903 54904
0 54906 5 1 1 54905
0 54907 7 1 2 72603 95138
0 54908 5 1 1 54907
0 54909 7 1 2 88684 89165
0 54910 5 1 1 54909
0 54911 7 1 2 89008 54910
0 54912 7 1 2 54908 54911
0 54913 5 1 1 54912
0 54914 7 1 2 97286 54913
0 54915 5 1 1 54914
0 54916 7 1 2 68802 54915
0 54917 7 1 2 54906 54916
0 54918 7 1 2 54901 54917
0 54919 7 1 2 54883 54918
0 54920 7 1 2 54860 54919
0 54921 7 1 2 54814 54920
0 54922 5 1 1 54921
0 54923 7 1 2 66777 54922
0 54924 7 1 2 54781 54923
0 54925 5 1 1 54924
0 54926 7 1 2 54604 54925
0 54927 7 2 2 54515 54926
0 54928 5 1 1 98578
0 54929 7 1 2 61947 98579
0 54930 5 1 1 54929
0 54931 7 1 2 65647 54930
0 54932 7 1 2 54294 54931
0 54933 5 1 1 54932
0 54934 7 1 2 75367 88501
0 54935 5 1 1 54934
0 54936 7 1 2 91662 54935
0 54937 5 1 1 54936
0 54938 7 1 2 88537 54937
0 54939 5 1 1 54938
0 54940 7 1 2 61948 97287
0 54941 7 1 2 54939 54940
0 54942 5 1 1 54941
0 54943 7 1 2 78483 82226
0 54944 7 1 2 94184 97233
0 54945 7 1 2 54943 54944
0 54946 5 1 1 54945
0 54947 7 1 2 54942 54946
0 54948 5 1 1 54947
0 54949 7 1 2 63219 54948
0 54950 5 1 1 54949
0 54951 7 1 2 64362 89900
0 54952 5 1 1 54951
0 54953 7 1 2 72392 97076
0 54954 5 1 1 54953
0 54955 7 1 2 71263 54954
0 54956 7 1 2 54952 54955
0 54957 5 1 1 54956
0 54958 7 1 2 70347 54957
0 54959 5 1 1 54958
0 54960 7 2 2 67781 77253
0 54961 5 1 1 98580
0 54962 7 2 2 73138 98581
0 54963 5 1 1 98582
0 54964 7 1 2 60959 83292
0 54965 5 1 1 54964
0 54966 7 1 2 89366 54965
0 54967 5 1 1 54966
0 54968 7 1 2 98583 54967
0 54969 5 1 1 54968
0 54970 7 1 2 66081 54969
0 54971 5 1 1 54970
0 54972 7 1 2 81654 95586
0 54973 5 2 1 54972
0 54974 7 1 2 65038 98584
0 54975 5 1 1 54974
0 54976 7 1 2 70380 97250
0 54977 5 1 1 54976
0 54978 7 2 2 97246 54977
0 54979 5 1 1 98586
0 54980 7 1 2 72788 54963
0 54981 5 2 1 54980
0 54982 7 1 2 74896 95378
0 54983 7 1 2 98588 54982
0 54984 7 1 2 98587 54983
0 54985 7 1 2 54975 54984
0 54986 7 1 2 54971 54985
0 54987 7 1 2 54959 54986
0 54988 5 1 1 54987
0 54989 7 1 2 65303 54988
0 54990 5 1 1 54989
0 54991 7 1 2 88477 95574
0 54992 5 1 1 54991
0 54993 7 1 2 65304 95370
0 54994 5 1 1 54993
0 54995 7 1 2 85665 54994
0 54996 7 1 2 54992 54995
0 54997 5 1 1 54996
0 54998 7 1 2 66344 54997
0 54999 5 1 1 54998
0 55000 7 1 2 61373 84916
0 55001 5 1 1 55000
0 55002 7 1 2 82310 55001
0 55003 5 1 1 55002
0 55004 7 1 2 82123 55003
0 55005 5 1 1 55004
0 55006 7 1 2 70348 55005
0 55007 5 1 1 55006
0 55008 7 1 2 65747 84069
0 55009 5 1 1 55008
0 55010 7 1 2 73139 88436
0 55011 5 1 1 55010
0 55012 7 1 2 66345 55011
0 55013 5 1 1 55012
0 55014 7 1 2 55009 55013
0 55015 7 1 2 55007 55014
0 55016 5 1 1 55015
0 55017 7 1 2 72393 55016
0 55018 5 1 1 55017
0 55019 7 1 2 90457 97244
0 55020 7 1 2 97097 55019
0 55021 5 1 1 55020
0 55022 7 1 2 77694 55021
0 55023 5 1 1 55022
0 55024 7 1 2 81468 71275
0 55025 5 1 1 55024
0 55026 7 1 2 95548 54979
0 55027 5 1 1 55026
0 55028 7 1 2 55025 55027
0 55029 7 1 2 55023 55028
0 55030 7 1 2 55018 55029
0 55031 5 2 1 55030
0 55032 7 1 2 65039 98590
0 55033 5 1 1 55032
0 55034 7 1 2 54999 55033
0 55035 7 1 2 54990 55034
0 55036 5 1 1 55035
0 55037 7 1 2 86064 55036
0 55038 5 1 1 55037
0 55039 7 1 2 94256 96868
0 55040 7 1 2 97238 55039
0 55041 5 1 1 55040
0 55042 7 1 2 55038 55041
0 55043 5 1 1 55042
0 55044 7 1 2 66595 55043
0 55045 5 1 1 55044
0 55046 7 1 2 87096 98585
0 55047 5 1 1 55046
0 55048 7 1 2 61949 81779
0 55049 7 1 2 98591 55048
0 55050 5 1 1 55049
0 55051 7 1 2 55047 55050
0 55052 5 1 1 55051
0 55053 7 1 2 65040 55052
0 55054 5 1 1 55053
0 55055 7 1 2 64363 87097
0 55056 5 2 1 55055
0 55057 7 2 2 81780 86263
0 55058 7 1 2 77994 98594
0 55059 5 1 1 55058
0 55060 7 1 2 98592 55059
0 55061 5 1 1 55060
0 55062 7 1 2 64598 55061
0 55063 5 1 1 55062
0 55064 7 2 2 76654 86505
0 55065 7 1 2 93523 98596
0 55066 5 1 1 55065
0 55067 7 1 2 55063 55066
0 55068 5 1 1 55067
0 55069 7 1 2 70381 55068
0 55070 5 1 1 55069
0 55071 7 1 2 93624 98595
0 55072 5 1 1 55071
0 55073 7 1 2 75807 86985
0 55074 5 1 1 55073
0 55075 7 1 2 55072 55074
0 55076 5 1 1 55075
0 55077 7 1 2 64825 55076
0 55078 5 1 1 55077
0 55079 7 1 2 66925 87930
0 55080 5 1 1 55079
0 55081 7 1 2 94950 98597
0 55082 5 1 1 55081
0 55083 7 1 2 55082 98593
0 55084 5 1 1 55083
0 55085 7 1 2 80070 55084
0 55086 5 1 1 55085
0 55087 7 1 2 55080 55086
0 55088 7 1 2 55078 55087
0 55089 7 1 2 55070 55088
0 55090 5 1 1 55089
0 55091 7 1 2 66082 55090
0 55092 5 1 1 55091
0 55093 7 1 2 74424 87098
0 55094 5 1 1 55093
0 55095 7 1 2 84637 86506
0 55096 7 1 2 93090 55095
0 55097 7 1 2 88478 55096
0 55098 5 1 1 55097
0 55099 7 1 2 55094 55098
0 55100 5 1 1 55099
0 55101 7 1 2 62402 55100
0 55102 5 1 1 55101
0 55103 7 1 2 66926 81734
0 55104 5 1 1 55103
0 55105 7 1 2 55102 55104
0 55106 7 1 2 55092 55105
0 55107 5 1 1 55106
0 55108 7 1 2 71937 55107
0 55109 5 1 1 55108
0 55110 7 1 2 72477 85080
0 55111 5 1 1 55110
0 55112 7 1 2 64364 55111
0 55113 5 1 1 55112
0 55114 7 1 2 90658 55113
0 55115 5 1 1 55114
0 55116 7 1 2 70349 55115
0 55117 5 1 1 55116
0 55118 7 1 2 64599 54961
0 55119 5 1 1 55118
0 55120 7 1 2 77328 55119
0 55121 5 1 1 55120
0 55122 7 1 2 70382 55121
0 55123 5 1 1 55122
0 55124 7 1 2 82504 82556
0 55125 5 1 1 55124
0 55126 7 1 2 66346 55125
0 55127 5 1 1 55126
0 55128 7 1 2 60412 78090
0 55129 7 1 2 98589 55128
0 55130 7 1 2 55127 55129
0 55131 7 1 2 55123 55130
0 55132 7 1 2 55117 55131
0 55133 5 1 1 55132
0 55134 7 1 2 86986 55133
0 55135 5 1 1 55134
0 55136 7 1 2 77975 81318
0 55137 7 1 2 86264 55136
0 55138 7 1 2 74432 55137
0 55139 7 1 2 81885 55138
0 55140 5 1 1 55139
0 55141 7 1 2 55135 55140
0 55142 7 1 2 55109 55141
0 55143 7 1 2 55054 55142
0 55144 7 1 2 55045 55143
0 55145 7 1 2 54950 55144
0 55146 5 1 1 55145
0 55147 7 1 2 68803 55146
0 55148 5 1 1 55147
0 55149 7 1 2 74141 84054
0 55150 7 1 2 97042 55149
0 55151 5 1 1 55150
0 55152 7 1 2 66083 55151
0 55153 5 1 1 55152
0 55154 7 1 2 68166 55153
0 55155 7 1 2 90228 55154
0 55156 5 1 1 55155
0 55157 7 1 2 75641 55156
0 55158 5 1 1 55157
0 55159 7 1 2 60413 91314
0 55160 5 1 1 55159
0 55161 7 1 2 72604 55160
0 55162 5 1 1 55161
0 55163 7 1 2 94536 55162
0 55164 5 1 1 55163
0 55165 7 1 2 62159 55164
0 55166 5 1 1 55165
0 55167 7 1 2 75642 94704
0 55168 5 1 1 55167
0 55169 7 1 2 55166 55168
0 55170 5 1 1 55169
0 55171 7 1 2 65907 55170
0 55172 5 1 1 55171
0 55173 7 1 2 75643 77101
0 55174 5 1 1 55173
0 55175 7 1 2 12229 55174
0 55176 7 1 2 55172 55175
0 55177 5 1 1 55176
0 55178 7 1 2 66084 76374
0 55179 7 1 2 55177 55178
0 55180 5 1 1 55179
0 55181 7 1 2 55158 55180
0 55182 5 1 1 55181
0 55183 7 1 2 64826 55182
0 55184 5 1 1 55183
0 55185 7 1 2 82633 84719
0 55186 5 1 1 55185
0 55187 7 1 2 62782 55186
0 55188 5 1 1 55187
0 55189 7 1 2 62160 96825
0 55190 5 1 1 55189
0 55191 7 1 2 55188 55190
0 55192 5 1 1 55191
0 55193 7 1 2 69714 55192
0 55194 5 1 1 55193
0 55195 7 1 2 65908 91178
0 55196 5 1 1 55195
0 55197 7 1 2 25987 55196
0 55198 5 1 1 55197
0 55199 7 1 2 72605 55198
0 55200 5 1 1 55199
0 55201 7 1 2 68167 90234
0 55202 5 1 1 55201
0 55203 7 1 2 69162 55202
0 55204 5 1 1 55203
0 55205 7 1 2 83821 90243
0 55206 5 1 1 55205
0 55207 7 1 2 75368 55206
0 55208 7 1 2 55204 55207
0 55209 7 1 2 55200 55208
0 55210 7 1 2 55194 55209
0 55211 5 1 1 55210
0 55212 7 1 2 75644 55211
0 55213 5 1 1 55212
0 55214 7 1 2 55184 55213
0 55215 5 1 1 55214
0 55216 7 1 2 70874 55215
0 55217 5 1 1 55216
0 55218 7 1 2 90885 95017
0 55219 5 1 1 55218
0 55220 7 1 2 84894 88756
0 55221 5 1 1 55220
0 55222 7 1 2 64827 55221
0 55223 5 1 1 55222
0 55224 7 1 2 81469 71938
0 55225 5 1 1 55224
0 55226 7 1 2 89046 55225
0 55227 7 1 2 55223 55226
0 55228 7 1 2 89140 55227
0 55229 5 1 1 55228
0 55230 7 1 2 97257 55229
0 55231 5 1 1 55230
0 55232 7 1 2 62783 80289
0 55233 7 1 2 88479 97273
0 55234 7 1 2 55232 55233
0 55235 5 1 1 55234
0 55236 7 1 2 91746 55235
0 55237 7 1 2 55231 55236
0 55238 7 1 2 55219 55237
0 55239 7 1 2 55217 55238
0 55240 5 1 1 55239
0 55241 7 1 2 97611 55240
0 55242 5 1 1 55241
0 55243 7 1 2 55148 55242
0 55244 5 1 1 55243
0 55245 7 1 2 65648 55244
0 55246 5 1 1 55245
0 55247 7 1 2 63220 95863
0 55248 5 1 1 55247
0 55249 7 1 2 74839 95152
0 55250 5 1 1 55249
0 55251 7 1 2 55248 55250
0 55252 5 1 1 55251
0 55253 7 1 2 75240 55252
0 55254 5 1 1 55253
0 55255 7 1 2 69438 93310
0 55256 5 1 1 55255
0 55257 7 1 2 70875 55256
0 55258 5 1 1 55257
0 55259 7 1 2 78893 90439
0 55260 5 1 1 55259
0 55261 7 1 2 55258 55260
0 55262 5 1 1 55261
0 55263 7 1 2 75645 55262
0 55264 5 1 1 55263
0 55265 7 1 2 66085 88334
0 55266 7 1 2 93755 55265
0 55267 5 1 1 55266
0 55268 7 1 2 55264 55267
0 55269 5 1 1 55268
0 55270 7 1 2 64828 55269
0 55271 5 1 1 55270
0 55272 7 1 2 66086 70383
0 55273 5 1 1 55272
0 55274 7 1 2 59700 55273
0 55275 5 1 1 55274
0 55276 7 1 2 98573 55275
0 55277 5 1 1 55276
0 55278 7 1 2 89512 55277
0 55279 5 1 1 55278
0 55280 7 1 2 75646 55279
0 55281 5 1 1 55280
0 55282 7 1 2 80290 88786
0 55283 5 1 1 55282
0 55284 7 1 2 88504 55283
0 55285 5 1 1 55284
0 55286 7 1 2 63221 91433
0 55287 7 1 2 55285 55286
0 55288 5 1 1 55287
0 55289 7 1 2 55281 55288
0 55290 7 1 2 55271 55289
0 55291 5 1 1 55290
0 55292 7 1 2 62403 55291
0 55293 5 1 1 55292
0 55294 7 1 2 75647 87483
0 55295 5 1 1 55294
0 55296 7 1 2 86553 55295
0 55297 5 1 1 55296
0 55298 7 1 2 72394 95450
0 55299 7 1 2 55297 55298
0 55300 5 1 1 55299
0 55301 7 1 2 76034 79087
0 55302 5 1 1 55301
0 55303 7 1 2 91135 55302
0 55304 5 1 1 55303
0 55305 7 1 2 75648 55304
0 55306 5 1 1 55305
0 55307 7 1 2 76429 93111
0 55308 5 1 1 55307
0 55309 7 1 2 70218 84663
0 55310 5 1 1 55309
0 55311 7 1 2 75649 55310
0 55312 5 1 1 55311
0 55313 7 1 2 75369 86017
0 55314 7 1 2 55312 55313
0 55315 5 1 1 55314
0 55316 7 1 2 55308 55315
0 55317 5 1 1 55316
0 55318 7 1 2 55306 55317
0 55319 7 1 2 55300 55318
0 55320 7 1 2 55293 55319
0 55321 5 1 1 55320
0 55322 7 1 2 62784 55321
0 55323 5 1 1 55322
0 55324 7 1 2 89386 95018
0 55325 5 1 1 55324
0 55326 7 1 2 15946 55325
0 55327 5 1 1 55326
0 55328 7 1 2 64365 55327
0 55329 5 1 1 55328
0 55330 7 2 2 72028 75650
0 55331 7 1 2 87032 98598
0 55332 5 1 1 55331
0 55333 7 1 2 87250 55332
0 55334 7 1 2 55329 55333
0 55335 5 1 1 55334
0 55336 7 1 2 72395 55335
0 55337 5 1 1 55336
0 55338 7 1 2 84978 90410
0 55339 5 1 1 55338
0 55340 7 1 2 59701 84400
0 55341 5 1 1 55340
0 55342 7 1 2 83822 55341
0 55343 7 1 2 97336 55342
0 55344 5 1 1 55343
0 55345 7 1 2 55339 55344
0 55346 7 1 2 55337 55345
0 55347 5 1 1 55346
0 55348 7 1 2 70350 55347
0 55349 5 1 1 55348
0 55350 7 1 2 70876 97248
0 55351 5 1 1 55350
0 55352 7 1 2 84664 45779
0 55353 7 1 2 55351 55352
0 55354 5 1 1 55353
0 55355 7 1 2 75651 55354
0 55356 5 1 1 55355
0 55357 7 1 2 86018 10290
0 55358 7 1 2 55356 55357
0 55359 5 1 1 55358
0 55360 7 1 2 82794 55359
0 55361 5 1 1 55360
0 55362 7 1 2 91236 55361
0 55363 5 1 1 55362
0 55364 7 1 2 69283 55363
0 55365 5 1 1 55364
0 55366 7 1 2 73882 95606
0 55367 5 1 1 55366
0 55368 7 1 2 76436 89505
0 55369 5 1 1 55368
0 55370 7 1 2 80299 87558
0 55371 5 1 1 55370
0 55372 7 1 2 91136 55371
0 55373 7 1 2 55369 55372
0 55374 7 1 2 55367 55373
0 55375 5 1 1 55374
0 55376 7 1 2 73982 55375
0 55377 5 1 1 55376
0 55378 7 1 2 88938 89506
0 55379 5 1 1 55378
0 55380 7 1 2 73280 95761
0 55381 5 1 1 55380
0 55382 7 1 2 74842 55381
0 55383 5 1 1 55382
0 55384 7 1 2 16150 55383
0 55385 5 1 1 55384
0 55386 7 1 2 55379 55385
0 55387 7 1 2 55377 55386
0 55388 5 1 1 55387
0 55389 7 1 2 75652 55388
0 55390 5 1 1 55389
0 55391 7 1 2 85067 88251
0 55392 5 1 1 55391
0 55393 7 1 2 73281 55392
0 55394 5 1 1 55393
0 55395 7 1 2 93092 55394
0 55396 5 1 1 55395
0 55397 7 1 2 61615 35002
0 55398 5 1 1 55397
0 55399 7 1 2 55396 55398
0 55400 5 1 1 55399
0 55401 7 1 2 90284 94797
0 55402 5 1 1 55401
0 55403 7 1 2 63222 71033
0 55404 5 1 1 55403
0 55405 7 1 2 55402 55404
0 55406 5 1 1 55405
0 55407 7 1 2 73282 55406
0 55408 5 1 1 55407
0 55409 7 1 2 77332 86378
0 55410 5 1 1 55409
0 55411 7 1 2 76812 55410
0 55412 5 1 1 55411
0 55413 7 1 2 66596 55412
0 55414 5 1 1 55413
0 55415 7 1 2 73352 94697
0 55416 7 1 2 73983 55415
0 55417 7 1 2 94021 55416
0 55418 5 1 1 55417
0 55419 7 1 2 55414 55418
0 55420 7 1 2 55408 55419
0 55421 7 1 2 55400 55420
0 55422 7 1 2 55390 55421
0 55423 7 1 2 55365 55422
0 55424 7 1 2 55349 55423
0 55425 7 1 2 55323 55424
0 55426 5 1 1 55425
0 55427 7 1 2 65530 55426
0 55428 5 1 1 55427
0 55429 7 1 2 55254 55428
0 55430 5 1 1 55429
0 55431 7 1 2 86767 55430
0 55432 5 1 1 55431
0 55433 7 1 2 61616 90367
0 55434 5 1 1 55433
0 55435 7 1 2 89732 55434
0 55436 5 1 1 55435
0 55437 7 1 2 67143 55436
0 55438 5 1 1 55437
0 55439 7 1 2 59702 75883
0 55440 5 1 1 55439
0 55441 7 1 2 40983 55440
0 55442 5 1 1 55441
0 55443 7 1 2 67782 55442
0 55444 5 1 1 55443
0 55445 7 1 2 55438 55444
0 55446 5 1 1 55445
0 55447 7 1 2 68168 55446
0 55448 5 1 1 55447
0 55449 7 1 2 62785 73070
0 55450 5 1 1 55449
0 55451 7 1 2 71399 94065
0 55452 7 1 2 55450 55451
0 55453 7 1 2 15772 90350
0 55454 7 1 2 55452 55453
0 55455 5 1 1 55454
0 55456 7 1 2 60626 55455
0 55457 5 1 1 55456
0 55458 7 1 2 55448 55457
0 55459 5 1 1 55458
0 55460 7 1 2 86812 55459
0 55461 5 1 1 55460
0 55462 7 1 2 78446 93115
0 55463 5 1 1 55462
0 55464 7 1 2 69613 55463
0 55465 5 1 1 55464
0 55466 7 1 2 40150 97540
0 55467 7 1 2 55465 55466
0 55468 5 1 1 55467
0 55469 7 1 2 59703 55468
0 55470 5 1 1 55469
0 55471 7 1 2 74126 84398
0 55472 5 1 1 55471
0 55473 7 1 2 72274 90985
0 55474 7 1 2 55472 55473
0 55475 5 1 1 55474
0 55476 7 1 2 55470 55475
0 55477 5 1 1 55476
0 55478 7 1 2 97603 55477
0 55479 5 1 1 55478
0 55480 7 1 2 88704 88707
0 55481 7 1 2 95114 55480
0 55482 5 1 1 55481
0 55483 7 1 2 55479 55482
0 55484 5 1 1 55483
0 55485 7 1 2 70713 55484
0 55486 5 1 1 55485
0 55487 7 1 2 63872 55486
0 55488 7 1 2 55461 55487
0 55489 7 1 2 55432 55488
0 55490 5 1 1 55489
0 55491 7 1 2 90340 88480
0 55492 5 1 1 55491
0 55493 7 1 2 90537 55492
0 55494 5 1 1 55493
0 55495 7 1 2 55494 98599
0 55496 5 1 1 55495
0 55497 7 1 2 67783 95187
0 55498 7 1 2 45177 55497
0 55499 7 1 2 72606 90224
0 55500 5 1 1 55499
0 55501 7 1 2 91377 91878
0 55502 5 1 1 55501
0 55503 7 1 2 97265 55502
0 55504 7 1 2 55500 55503
0 55505 7 1 2 55498 55504
0 55506 5 1 1 55505
0 55507 7 1 2 97258 55506
0 55508 5 1 1 55507
0 55509 7 1 2 55496 55508
0 55510 5 1 1 55509
0 55511 7 1 2 72396 55510
0 55512 5 1 1 55511
0 55513 7 1 2 90403 97116
0 55514 5 1 1 55513
0 55515 7 1 2 70714 82564
0 55516 5 1 1 55515
0 55517 7 1 2 78239 55516
0 55518 5 1 1 55517
0 55519 7 1 2 97113 55518
0 55520 5 1 1 55519
0 55521 7 1 2 91879 55520
0 55522 5 1 1 55521
0 55523 7 1 2 81470 47484
0 55524 5 1 1 55523
0 55525 7 1 2 91725 55524
0 55526 7 1 2 55522 55525
0 55527 7 1 2 55514 55526
0 55528 7 1 2 55512 55527
0 55529 5 1 1 55528
0 55530 7 1 2 86813 55529
0 55531 5 1 1 55530
0 55532 7 1 2 87196 90435
0 55533 7 1 2 91652 55532
0 55534 5 1 1 55533
0 55535 7 1 2 60733 81274
0 55536 7 2 2 87530 55535
0 55537 5 1 1 98600
0 55538 7 1 2 86825 55537
0 55539 5 2 1 55538
0 55540 7 1 2 80293 95553
0 55541 7 1 2 98602 55540
0 55542 5 1 1 55541
0 55543 7 1 2 55534 55542
0 55544 5 1 1 55543
0 55545 7 1 2 65909 55544
0 55546 5 1 1 55545
0 55547 7 2 2 83486 87197
0 55548 7 1 2 72607 98604
0 55549 5 1 1 55548
0 55550 7 1 2 80291 97054
0 55551 7 1 2 98603 55550
0 55552 5 1 1 55551
0 55553 7 1 2 55549 55552
0 55554 5 1 1 55553
0 55555 7 1 2 69284 55554
0 55556 5 1 1 55555
0 55557 7 1 2 83962 82761
0 55558 5 1 1 55557
0 55559 7 1 2 98605 55558
0 55560 5 1 1 55559
0 55561 7 1 2 55556 55560
0 55562 7 1 2 55546 55561
0 55563 5 1 1 55562
0 55564 7 1 2 72397 55563
0 55565 5 1 1 55564
0 55566 7 1 2 86814 97330
0 55567 5 1 1 55566
0 55568 7 1 2 71136 98601
0 55569 5 1 1 55568
0 55570 7 1 2 86815 97334
0 55571 5 1 1 55570
0 55572 7 1 2 55569 55571
0 55573 5 1 1 55572
0 55574 7 1 2 12746 55573
0 55575 5 1 1 55574
0 55576 7 1 2 55567 55575
0 55577 7 1 2 55565 55576
0 55578 5 1 1 55577
0 55579 7 1 2 63223 55578
0 55580 5 1 1 55579
0 55581 7 1 2 68804 55580
0 55582 7 1 2 55531 55581
0 55583 5 1 1 55582
0 55584 7 1 2 66778 55583
0 55585 7 1 2 55490 55584
0 55586 5 1 1 55585
0 55587 7 1 2 84560 44667
0 55588 5 2 1 55587
0 55589 7 1 2 65910 84530
0 55590 5 3 1 55589
0 55591 7 1 2 71472 98608
0 55592 5 1 1 55591
0 55593 7 1 2 72398 55592
0 55594 7 1 2 98606 55593
0 55595 5 1 1 55594
0 55596 7 2 2 72029 84531
0 55597 5 1 1 98611
0 55598 7 1 2 45378 55597
0 55599 5 1 1 55598
0 55600 7 1 2 71463 55599
0 55601 5 1 1 55600
0 55602 7 1 2 80485 71264
0 55603 5 1 1 55602
0 55604 7 1 2 84532 55603
0 55605 5 1 1 55604
0 55606 7 1 2 55601 55605
0 55607 7 1 2 55595 55606
0 55608 5 1 1 55607
0 55609 7 1 2 62404 55608
0 55610 5 1 1 55609
0 55611 7 1 2 84155 84638
0 55612 5 1 1 55611
0 55613 7 1 2 84561 55612
0 55614 5 2 1 55613
0 55615 7 1 2 63224 98613
0 55616 5 1 1 55615
0 55617 7 1 2 80500 84205
0 55618 5 1 1 55617
0 55619 7 1 2 76457 84533
0 55620 5 1 1 55619
0 55621 7 1 2 55618 55620
0 55622 5 1 1 55621
0 55623 7 1 2 71137 55622
0 55624 5 1 1 55623
0 55625 7 1 2 55616 55624
0 55626 7 1 2 55610 55625
0 55627 5 1 1 55626
0 55628 7 1 2 62786 55627
0 55629 5 1 1 55628
0 55630 7 1 2 70293 84562
0 55631 5 1 1 55630
0 55632 7 1 2 94578 55631
0 55633 7 1 2 98607 55632
0 55634 5 1 1 55633
0 55635 7 1 2 59704 98609
0 55636 5 1 1 55635
0 55637 7 1 2 65748 98614
0 55638 7 1 2 55636 55637
0 55639 5 1 1 55638
0 55640 7 1 2 55634 55639
0 55641 5 1 1 55640
0 55642 7 1 2 71138 55641
0 55643 5 1 1 55642
0 55644 7 1 2 45395 98610
0 55645 5 1 1 55644
0 55646 7 1 2 63225 55645
0 55647 5 1 1 55646
0 55648 7 1 2 55643 55647
0 55649 5 1 1 55648
0 55650 7 1 2 62405 55649
0 55651 5 1 1 55650
0 55652 7 1 2 93588 93892
0 55653 5 2 1 55652
0 55654 7 1 2 88528 98615
0 55655 5 1 1 55654
0 55656 7 1 2 27464 97179
0 55657 7 1 2 55655 55656
0 55658 5 1 1 55657
0 55659 7 1 2 78626 55658
0 55660 5 1 1 55659
0 55661 7 1 2 62787 98612
0 55662 5 1 1 55661
0 55663 7 1 2 97314 55662
0 55664 5 1 1 55663
0 55665 7 1 2 83688 55664
0 55666 5 1 1 55665
0 55667 7 1 2 84563 93893
0 55668 5 1 1 55667
0 55669 7 1 2 63226 55668
0 55670 5 1 1 55669
0 55671 7 1 2 55666 55670
0 55672 7 1 2 55660 55671
0 55673 5 1 1 55672
0 55674 7 1 2 72399 55673
0 55675 5 1 1 55674
0 55676 7 1 2 63227 75810
0 55677 5 1 1 55676
0 55678 7 1 2 85798 55677
0 55679 5 1 1 55678
0 55680 7 1 2 98616 55679
0 55681 5 1 1 55680
0 55682 7 2 2 64600 84534
0 55683 5 1 1 98617
0 55684 7 1 2 93516 55683
0 55685 5 1 1 55684
0 55686 7 1 2 90967 93255
0 55687 5 1 1 55686
0 55688 7 1 2 64366 55687
0 55689 5 1 1 55688
0 55690 7 1 2 65749 86403
0 55691 5 1 1 55690
0 55692 7 1 2 55689 55691
0 55693 5 1 1 55692
0 55694 7 1 2 55685 55693
0 55695 5 1 1 55694
0 55696 7 1 2 84206 79069
0 55697 5 2 1 55696
0 55698 7 1 2 55695 98619
0 55699 7 1 2 55681 55698
0 55700 7 1 2 55675 55699
0 55701 7 1 2 55651 55700
0 55702 7 1 2 55629 55701
0 55703 5 1 1 55702
0 55704 7 1 2 75653 55703
0 55705 5 1 1 55704
0 55706 7 1 2 84535 91880
0 55707 5 1 1 55706
0 55708 7 1 2 69346 71900
0 55709 7 1 2 97358 55708
0 55710 5 1 1 55709
0 55711 7 1 2 97212 55710
0 55712 5 1 1 55711
0 55713 7 1 2 55707 55712
0 55714 7 1 2 55705 55713
0 55715 5 1 1 55714
0 55716 7 1 2 87117 55715
0 55717 5 1 1 55716
0 55718 7 1 2 63228 80446
0 55719 5 1 1 55718
0 55720 7 1 2 91449 55719
0 55721 5 1 1 55720
0 55722 7 1 2 84207 55721
0 55723 5 1 1 55722
0 55724 7 1 2 90867 93584
0 55725 5 1 1 55724
0 55726 7 1 2 84536 91179
0 55727 5 1 1 55726
0 55728 7 1 2 55725 55727
0 55729 7 1 2 55723 55728
0 55730 5 1 1 55729
0 55731 7 1 2 65911 55730
0 55732 5 1 1 55731
0 55733 7 2 2 65531 85206
0 55734 5 1 1 98621
0 55735 7 1 2 84564 55734
0 55736 5 1 1 55735
0 55737 7 1 2 89053 55736
0 55738 5 1 1 55737
0 55739 7 1 2 62788 94852
0 55740 5 1 1 55739
0 55741 7 1 2 28060 55740
0 55742 7 1 2 55738 55741
0 55743 5 1 1 55742
0 55744 7 1 2 62406 55743
0 55745 5 1 1 55744
0 55746 7 1 2 55732 55745
0 55747 5 1 1 55746
0 55748 7 1 2 75654 55747
0 55749 5 1 1 55748
0 55750 7 1 2 84259 97127
0 55751 5 1 1 55750
0 55752 7 1 2 55749 55751
0 55753 5 1 1 55752
0 55754 7 1 2 87118 55753
0 55755 5 1 1 55754
0 55756 7 1 2 70951 85675
0 55757 7 1 2 93535 55756
0 55758 7 1 2 93075 95100
0 55759 7 1 2 55757 55758
0 55760 5 1 1 55759
0 55761 7 1 2 55755 55760
0 55762 5 1 1 55761
0 55763 7 1 2 72608 55762
0 55764 5 1 1 55763
0 55765 7 1 2 64601 97176
0 55766 5 1 1 55765
0 55767 7 1 2 45600 55766
0 55768 5 1 1 55767
0 55769 7 1 2 90387 55768
0 55770 5 1 1 55769
0 55771 7 1 2 97214 55770
0 55772 5 1 1 55771
0 55773 7 1 2 87119 55772
0 55774 5 1 1 55773
0 55775 7 1 2 87135 94375
0 55776 5 2 1 55775
0 55777 7 1 2 78627 85216
0 55778 7 1 2 98623 55777
0 55779 5 1 1 55778
0 55780 7 1 2 82277 90240
0 55781 5 1 1 55780
0 55782 7 5 2 68805 87120
0 55783 7 1 2 91663 98625
0 55784 7 1 2 55781 55783
0 55785 5 1 1 55784
0 55786 7 1 2 55779 55785
0 55787 5 1 1 55786
0 55788 7 1 2 63229 55787
0 55789 5 1 1 55788
0 55790 7 1 2 87121 91221
0 55791 7 1 2 98618 55790
0 55792 5 1 1 55791
0 55793 7 1 2 55789 55792
0 55794 5 1 1 55793
0 55795 7 1 2 62407 55794
0 55796 5 1 1 55795
0 55797 7 1 2 55774 55796
0 55798 5 1 1 55797
0 55799 7 1 2 76375 55798
0 55800 5 1 1 55799
0 55801 7 1 2 55764 55800
0 55802 7 1 2 55717 55801
0 55803 5 1 1 55802
0 55804 7 1 2 70877 55803
0 55805 5 1 1 55804
0 55806 7 1 2 66087 84208
0 55807 5 1 1 55806
0 55808 7 1 2 84565 55807
0 55809 5 1 1 55808
0 55810 7 1 2 64367 55809
0 55811 5 1 1 55810
0 55812 7 1 2 93894 55811
0 55813 5 1 1 55812
0 55814 7 1 2 69380 55813
0 55815 5 1 1 55814
0 55816 7 1 2 82311 84537
0 55817 5 1 1 55816
0 55818 7 1 2 64829 97171
0 55819 5 1 1 55818
0 55820 7 1 2 55817 55819
0 55821 7 1 2 55815 55820
0 55822 5 1 1 55821
0 55823 7 1 2 70094 55822
0 55824 5 1 1 55823
0 55825 7 1 2 82329 96785
0 55826 5 1 1 55825
0 55827 7 1 2 84209 55826
0 55828 5 1 1 55827
0 55829 7 1 2 45391 55828
0 55830 5 1 1 55829
0 55831 7 1 2 91250 55830
0 55832 5 1 1 55831
0 55833 7 1 2 55824 55832
0 55834 5 1 1 55833
0 55835 7 1 2 75655 55834
0 55836 5 1 1 55835
0 55837 7 1 2 81329 84783
0 55838 5 1 1 55837
0 55839 7 1 2 84566 55838
0 55840 5 1 1 55839
0 55841 7 1 2 89367 55840
0 55842 5 1 1 55841
0 55843 7 1 2 84781 86011
0 55844 5 1 1 55843
0 55845 7 1 2 93580 55844
0 55846 5 2 1 55845
0 55847 7 1 2 64368 98630
0 55848 5 1 1 55847
0 55849 7 1 2 55842 55848
0 55850 5 1 1 55849
0 55851 7 1 2 91881 55850
0 55852 5 1 1 55851
0 55853 7 1 2 84643 93524
0 55854 5 1 1 55853
0 55855 7 1 2 90287 97213
0 55856 5 1 1 55855
0 55857 7 2 2 79383 84255
0 55858 5 1 1 98632
0 55859 7 1 2 93389 98633
0 55860 5 1 1 55859
0 55861 7 1 2 55856 55860
0 55862 5 1 1 55861
0 55863 7 1 2 69381 55862
0 55864 5 1 1 55863
0 55865 7 1 2 55854 55864
0 55866 7 1 2 55852 55865
0 55867 7 1 2 55836 55866
0 55868 5 1 1 55867
0 55869 7 1 2 87122 55868
0 55870 5 1 1 55869
0 55871 7 1 2 45701 55858
0 55872 5 1 1 55871
0 55873 7 1 2 64369 55872
0 55874 5 1 1 55873
0 55875 7 1 2 98620 55874
0 55876 5 1 1 55875
0 55877 7 1 2 62789 55876
0 55878 5 1 1 55877
0 55879 7 1 2 88238 94914
0 55880 5 1 1 55879
0 55881 7 1 2 55878 55880
0 55882 5 1 1 55881
0 55883 7 1 2 75656 55882
0 55884 5 1 1 55883
0 55885 7 1 2 91882 98631
0 55886 5 1 1 55885
0 55887 7 1 2 79350 84260
0 55888 5 1 1 55887
0 55889 7 1 2 97215 55888
0 55890 5 1 1 55889
0 55891 7 1 2 88862 55890
0 55892 5 1 1 55891
0 55893 7 1 2 55886 55892
0 55894 7 1 2 55884 55893
0 55895 5 1 1 55894
0 55896 7 1 2 87123 55895
0 55897 5 1 1 55896
0 55898 7 1 2 80976 79388
0 55899 7 1 2 85892 96304
0 55900 7 1 2 55898 55899
0 55901 5 1 1 55900
0 55902 7 1 2 55897 55901
0 55903 5 1 1 55902
0 55904 7 1 2 70351 55903
0 55905 5 1 1 55904
0 55906 7 1 2 87244 97172
0 55907 5 1 1 55906
0 55908 7 1 2 46263 55907
0 55909 5 1 1 55908
0 55910 7 1 2 87124 55909
0 55911 5 1 1 55910
0 55912 7 1 2 75657 87125
0 55913 5 1 1 55912
0 55914 7 1 2 70095 98624
0 55915 5 1 1 55914
0 55916 7 1 2 55913 55915
0 55917 5 4 1 55916
0 55918 7 1 2 78351 84538
0 55919 7 1 2 98634 55918
0 55920 5 1 1 55919
0 55921 7 2 2 84592 97288
0 55922 7 1 2 73231 87126
0 55923 7 1 2 98638 55922
0 55924 5 1 1 55923
0 55925 7 1 2 55920 55924
0 55926 5 1 1 55925
0 55927 7 1 2 83871 55926
0 55928 5 1 1 55927
0 55929 7 1 2 55911 55928
0 55930 5 1 1 55929
0 55931 7 1 2 71939 55930
0 55932 5 1 1 55931
0 55933 7 1 2 83954 93536
0 55934 5 1 1 55933
0 55935 7 1 2 3033 55934
0 55936 5 1 1 55935
0 55937 7 1 2 75658 55936
0 55938 5 1 1 55937
0 55939 7 1 2 93917 94915
0 55940 5 1 1 55939
0 55941 7 1 2 46064 55940
0 55942 7 1 2 55938 55941
0 55943 5 1 1 55942
0 55944 7 1 2 87127 55943
0 55945 5 1 1 55944
0 55946 7 1 2 85786 95119
0 55947 7 1 2 87845 91967
0 55948 7 1 2 55946 55947
0 55949 5 1 1 55948
0 55950 7 1 2 55945 55949
0 55951 5 1 1 55950
0 55952 7 1 2 93303 55951
0 55953 5 1 1 55952
0 55954 7 1 2 86286 86387
0 55955 7 1 2 87846 55954
0 55956 7 1 2 91251 93756
0 55957 7 1 2 55955 55956
0 55958 5 1 1 55957
0 55959 7 1 2 55953 55958
0 55960 7 1 2 55932 55959
0 55961 7 1 2 55905 55960
0 55962 7 1 2 55870 55961
0 55963 5 1 1 55962
0 55964 7 1 2 71842 55963
0 55965 5 1 1 55964
0 55966 7 1 2 72773 93081
0 55967 5 1 1 55966
0 55968 7 1 2 96452 55967
0 55969 5 1 1 55968
0 55970 7 1 2 65305 55969
0 55971 5 1 1 55970
0 55972 7 1 2 80432 93603
0 55973 5 1 1 55972
0 55974 7 1 2 55971 55973
0 55975 5 1 1 55974
0 55976 7 1 2 97169 55975
0 55977 5 1 1 55976
0 55978 7 1 2 84539 92925
0 55979 5 1 1 55978
0 55980 7 1 2 78409 97086
0 55981 5 1 1 55980
0 55982 7 1 2 97158 55981
0 55983 7 1 2 55979 55982
0 55984 5 1 1 55983
0 55985 7 1 2 65306 55984
0 55986 5 1 1 55985
0 55987 7 1 2 84567 93811
0 55988 5 1 1 55987
0 55989 7 1 2 63230 73896
0 55990 5 1 1 55989
0 55991 7 1 2 94564 55990
0 55992 5 1 1 55991
0 55993 7 1 2 55988 55992
0 55994 5 1 1 55993
0 55995 7 1 2 84086 84210
0 55996 5 1 1 55995
0 55997 7 1 2 34297 55996
0 55998 5 1 1 55997
0 55999 7 1 2 66597 55998
0 56000 5 1 1 55999
0 56001 7 1 2 55994 56000
0 56002 7 1 2 55986 56001
0 56003 5 1 1 56002
0 56004 7 1 2 70096 56003
0 56005 5 1 1 56004
0 56006 7 1 2 91883 92926
0 56007 5 1 1 56006
0 56008 7 1 2 73897 86840
0 56009 5 1 1 56008
0 56010 7 1 2 56007 56009
0 56011 5 1 1 56010
0 56012 7 1 2 84540 56011
0 56013 5 1 1 56012
0 56014 7 1 2 56005 56013
0 56015 7 1 2 55977 56014
0 56016 5 1 1 56015
0 56017 7 1 2 71940 56016
0 56018 5 1 1 56017
0 56019 7 2 2 62408 97154
0 56020 5 1 1 98640
0 56021 7 1 2 74714 84211
0 56022 5 1 1 56021
0 56023 7 1 2 56020 56022
0 56024 5 1 1 56023
0 56025 7 1 2 64370 56024
0 56026 5 1 1 56025
0 56027 7 1 2 77311 76074
0 56028 5 1 1 56027
0 56029 7 1 2 98622 56028
0 56030 5 1 1 56029
0 56031 7 1 2 56026 56030
0 56032 5 1 1 56031
0 56033 7 1 2 87245 56032
0 56034 5 1 1 56033
0 56035 7 1 2 93642 98641
0 56036 5 1 1 56035
0 56037 7 1 2 80340 93844
0 56038 5 1 1 56037
0 56039 7 1 2 30573 56038
0 56040 7 1 2 56036 56039
0 56041 7 1 2 56034 56040
0 56042 7 1 2 56018 56041
0 56043 5 1 1 56042
0 56044 7 1 2 87128 56043
0 56045 5 1 1 56044
0 56046 7 2 2 87129 97259
0 56047 5 1 1 98642
0 56048 7 1 2 74642 98643
0 56049 5 1 1 56048
0 56050 7 1 2 73831 89374
0 56051 7 1 2 93300 56050
0 56052 5 1 1 56051
0 56053 7 1 2 63231 88965
0 56054 7 1 2 98635 56053
0 56055 7 1 2 56052 56054
0 56056 5 1 1 56055
0 56057 7 1 2 56049 56056
0 56058 5 1 1 56057
0 56059 7 1 2 84541 56058
0 56060 5 1 1 56059
0 56061 7 3 2 65532 87246
0 56062 7 1 2 73219 98644
0 56063 5 1 1 56062
0 56064 7 1 2 95019 97283
0 56065 7 1 2 95458 56064
0 56066 5 1 1 56065
0 56067 7 1 2 56063 56066
0 56068 5 1 1 56067
0 56069 7 1 2 66088 56068
0 56070 5 1 1 56069
0 56071 7 1 2 83860 98645
0 56072 5 1 1 56071
0 56073 7 1 2 56070 56072
0 56074 5 1 1 56073
0 56075 7 1 2 98626 56074
0 56076 5 1 1 56075
0 56077 7 1 2 56060 56076
0 56078 5 1 1 56077
0 56079 7 1 2 73581 56078
0 56080 5 1 1 56079
0 56081 7 1 2 65912 98627
0 56082 7 2 2 97289 56081
0 56083 7 1 2 91267 98647
0 56084 5 1 1 56083
0 56085 7 1 2 71316 84261
0 56086 7 1 2 98636 56085
0 56087 5 1 1 56086
0 56088 7 1 2 56084 56087
0 56089 5 1 1 56088
0 56090 7 1 2 62409 56089
0 56091 5 1 1 56090
0 56092 7 1 2 73883 93304
0 56093 7 1 2 98648 56092
0 56094 5 1 1 56093
0 56095 7 1 2 56091 56094
0 56096 5 1 1 56095
0 56097 7 1 2 62790 56096
0 56098 5 1 1 56097
0 56099 7 1 2 80316 87130
0 56100 7 1 2 98639 56099
0 56101 5 1 1 56100
0 56102 7 1 2 56098 56101
0 56103 5 1 1 56102
0 56104 7 1 2 63232 56103
0 56105 5 1 1 56104
0 56106 7 1 2 88481 94832
0 56107 7 1 2 98637 56106
0 56108 5 1 1 56107
0 56109 7 1 2 56047 56108
0 56110 5 1 1 56109
0 56111 7 1 2 84542 56110
0 56112 5 1 1 56111
0 56113 7 1 2 98628 98646
0 56114 5 1 1 56113
0 56115 7 1 2 56112 56114
0 56116 5 1 1 56115
0 56117 7 1 2 89054 56116
0 56118 5 1 1 56117
0 56119 7 1 2 70502 98629
0 56120 5 1 1 56119
0 56121 7 1 2 65533 97612
0 56122 5 1 1 56121
0 56123 7 1 2 56120 56122
0 56124 5 1 1 56123
0 56125 7 1 2 71941 85801
0 56126 7 1 2 87486 56125
0 56127 7 1 2 56124 56126
0 56128 5 1 1 56127
0 56129 7 1 2 56118 56128
0 56130 7 1 2 56105 56129
0 56131 7 1 2 56080 56130
0 56132 7 1 2 56045 56131
0 56133 7 1 2 55965 56132
0 56134 7 1 2 55805 56133
0 56135 7 1 2 55586 56134
0 56136 7 1 2 55246 56135
0 56137 5 1 1 56136
0 56138 7 1 2 63595 56137
0 56139 5 1 1 56138
0 56140 7 1 2 66927 54928
0 56141 5 1 1 56140
0 56142 7 1 2 62791 73531
0 56143 5 1 1 56142
0 56144 7 1 2 86520 56143
0 56145 5 1 1 56144
0 56146 7 1 2 69715 56145
0 56147 5 1 1 56146
0 56148 7 1 2 69998 94078
0 56149 5 1 1 56148
0 56150 7 1 2 62161 72463
0 56151 5 1 1 56150
0 56152 7 1 2 56149 56151
0 56153 5 1 1 56152
0 56154 7 1 2 62792 56153
0 56155 5 1 1 56154
0 56156 7 1 2 56147 56155
0 56157 5 1 1 56156
0 56158 7 1 2 72400 56157
0 56159 5 1 1 56158
0 56160 7 1 2 90508 88396
0 56161 5 1 1 56160
0 56162 7 1 2 91139 56161
0 56163 5 1 1 56162
0 56164 7 1 2 70878 56163
0 56165 5 1 1 56164
0 56166 7 1 2 85986 90912
0 56167 7 1 2 81928 56166
0 56168 5 1 1 56167
0 56169 7 1 2 62793 56168
0 56170 5 1 1 56169
0 56171 7 1 2 56165 56170
0 56172 7 1 2 56159 56171
0 56173 5 1 1 56172
0 56174 7 1 2 63233 56173
0 56175 5 1 1 56174
0 56176 7 1 2 74897 89047
0 56177 5 1 1 56176
0 56178 7 1 2 70879 56177
0 56179 5 1 1 56178
0 56180 7 1 2 2720 56179
0 56181 5 1 1 56180
0 56182 7 1 2 90929 56181
0 56183 5 1 1 56182
0 56184 7 1 2 77746 95424
0 56185 5 1 1 56184
0 56186 7 1 2 72416 89605
0 56187 5 1 1 56186
0 56188 7 1 2 73495 56187
0 56189 5 1 1 56188
0 56190 7 1 2 56185 56189
0 56191 7 1 2 56183 56190
0 56192 7 1 2 56175 56191
0 56193 5 1 1 56192
0 56194 7 1 2 66598 56193
0 56195 5 1 1 56194
0 56196 7 1 2 86012 90930
0 56197 5 1 1 56196
0 56198 7 1 2 64602 88289
0 56199 5 1 1 56198
0 56200 7 1 2 95275 56199
0 56201 5 1 1 56200
0 56202 7 1 2 72401 56201
0 56203 5 1 1 56202
0 56204 7 1 2 71139 97229
0 56205 5 1 1 56204
0 56206 7 1 2 56203 56205
0 56207 5 1 1 56206
0 56208 7 1 2 63234 93390
0 56209 7 1 2 56207 56208
0 56210 5 1 1 56209
0 56211 7 1 2 56197 56210
0 56212 7 1 2 56195 56211
0 56213 5 1 1 56212
0 56214 7 1 2 65307 56213
0 56215 5 1 1 56214
0 56216 7 1 2 61617 98575
0 56217 5 1 1 56216
0 56218 7 1 2 65308 56217
0 56219 5 1 1 56218
0 56220 7 1 2 78953 85608
0 56221 5 1 1 56220
0 56222 7 1 2 56219 56221
0 56223 5 1 1 56222
0 56224 7 1 2 64371 56223
0 56225 5 1 1 56224
0 56226 7 1 2 70352 75241
0 56227 5 1 1 56226
0 56228 7 1 2 56225 56227
0 56229 5 1 1 56228
0 56230 7 1 2 62410 56229
0 56231 5 1 1 56230
0 56232 7 1 2 97252 56231
0 56233 5 1 1 56232
0 56234 7 1 2 95431 56233
0 56235 5 1 1 56234
0 56236 7 1 2 15626 95822
0 56237 5 1 1 56236
0 56238 7 1 2 64830 56237
0 56239 5 1 1 56238
0 56240 7 1 2 95820 56239
0 56241 5 1 1 56240
0 56242 7 1 2 71843 56241
0 56243 5 1 1 56242
0 56244 7 1 2 72030 90879
0 56245 5 1 1 56244
0 56246 7 1 2 81705 56245
0 56247 5 1 1 56246
0 56248 7 1 2 69999 56247
0 56249 5 1 1 56248
0 56250 7 1 2 72031 97046
0 56251 5 1 1 56250
0 56252 7 1 2 81706 56251
0 56253 5 1 1 56252
0 56254 7 1 2 62162 56253
0 56255 5 1 1 56254
0 56256 7 1 2 56249 56255
0 56257 7 1 2 56243 56256
0 56258 5 1 1 56257
0 56259 7 1 2 87487 56258
0 56260 5 1 1 56259
0 56261 7 1 2 56235 56260
0 56262 7 1 2 56215 56261
0 56263 5 1 1 56262
0 56264 7 1 2 93619 56263
0 56265 5 1 1 56264
0 56266 7 1 2 56141 56265
0 56267 5 1 1 56266
0 56268 7 1 2 60734 56267
0 56269 5 1 1 56268
0 56270 7 1 2 72402 95720
0 56271 7 1 2 87834 56270
0 56272 7 1 2 89716 94389
0 56273 7 1 2 56271 56272
0 56274 7 1 2 13019 56273
0 56275 5 1 1 56274
0 56276 7 1 2 56269 56275
0 56277 7 1 2 56139 56276
0 56278 7 1 2 54933 56277
0 56279 5 1 1 56278
0 56280 7 1 2 69032 56279
0 56281 5 1 1 56280
0 56282 7 1 2 69215 73369
0 56283 5 1 1 56282
0 56284 7 2 2 72403 56283
0 56285 5 1 1 98649
0 56286 7 1 2 77489 56285
0 56287 5 3 1 56286
0 56288 7 1 2 79298 98651
0 56289 5 1 1 56288
0 56290 7 1 2 91726 56289
0 56291 5 1 1 56290
0 56292 7 1 2 72032 78112
0 56293 5 1 1 56292
0 56294 7 1 2 95865 56293
0 56295 5 1 1 56294
0 56296 7 1 2 88482 56295
0 56297 5 1 1 56296
0 56298 7 1 2 72512 72172
0 56299 5 1 1 56298
0 56300 7 1 2 70915 92127
0 56301 7 1 2 56299 56300
0 56302 7 1 2 56297 56301
0 56303 5 1 1 56302
0 56304 7 1 2 68169 56303
0 56305 5 1 1 56304
0 56306 7 1 2 89524 39190
0 56307 7 1 2 95858 56306
0 56308 5 1 1 56307
0 56309 7 1 2 62794 56308
0 56310 5 1 1 56309
0 56311 7 1 2 56305 56310
0 56312 5 1 1 56311
0 56313 7 1 2 63235 98650
0 56314 5 1 1 56313
0 56315 7 1 2 61821 56314
0 56316 7 1 2 56312 56315
0 56317 5 1 1 56316
0 56318 7 1 2 56291 56317
0 56319 5 1 1 56318
0 56320 7 1 2 68563 56319
0 56321 5 1 1 56320
0 56322 7 1 2 59705 97507
0 56323 5 1 1 56322
0 56324 7 1 2 74912 56323
0 56325 5 1 1 56324
0 56326 7 1 2 69614 56325
0 56327 5 1 1 56326
0 56328 7 1 2 70880 73353
0 56329 5 1 1 56328
0 56330 7 1 2 67784 56329
0 56331 7 1 2 96008 56330
0 56332 5 1 1 56331
0 56333 7 1 2 89530 56332
0 56334 7 3 2 56327 56333
0 56335 5 1 1 98654
0 56336 7 1 2 86627 98655
0 56337 5 1 1 56336
0 56338 7 1 2 63596 56337
0 56339 5 1 1 56338
0 56340 7 1 2 60627 98130
0 56341 5 1 1 56340
0 56342 7 1 2 56339 56341
0 56343 5 1 1 56342
0 56344 7 1 2 75659 98656
0 56345 5 1 1 56344
0 56346 7 1 2 63597 91727
0 56347 7 1 2 56345 56346
0 56348 5 1 1 56347
0 56349 7 1 2 66779 56348
0 56350 5 1 1 56349
0 56351 7 1 2 56343 56350
0 56352 5 1 1 56351
0 56353 7 1 2 56321 56352
0 56354 5 1 1 56353
0 56355 7 1 2 61950 56354
0 56356 5 1 1 56355
0 56357 7 1 2 63598 96020
0 56358 7 2 2 56335 56357
0 56359 5 1 1 98657
0 56360 7 1 2 29847 98652
0 56361 5 1 1 56360
0 56362 7 1 2 82006 92128
0 56363 7 1 2 56361 56362
0 56364 5 1 1 56363
0 56365 7 1 2 56359 56364
0 56366 7 1 2 56356 56365
0 56367 5 1 1 56366
0 56368 7 1 2 60735 56367
0 56369 5 1 1 56368
0 56370 7 1 2 75531 96175
0 56371 5 1 1 56370
0 56372 7 1 2 96021 97297
0 56373 5 1 1 56372
0 56374 7 1 2 96190 56373
0 56375 5 1 1 56374
0 56376 7 1 2 56371 56375
0 56377 5 1 1 56376
0 56378 7 1 2 60736 56377
0 56379 5 1 1 56378
0 56380 7 1 2 95842 56379
0 56381 5 1 1 56380
0 56382 7 1 2 70544 56381
0 56383 5 1 1 56382
0 56384 7 3 2 62163 76945
0 56385 7 1 2 95839 98659
0 56386 5 1 1 56385
0 56387 7 1 2 91728 98660
0 56388 5 1 1 56387
0 56389 7 1 2 5534 95279
0 56390 5 1 1 56389
0 56391 7 1 2 62411 56390
0 56392 5 1 1 56391
0 56393 7 1 2 67394 79149
0 56394 5 1 1 56393
0 56395 7 1 2 95283 56394
0 56396 7 1 2 56392 56395
0 56397 5 1 1 56396
0 56398 7 1 2 61822 56397
0 56399 5 1 1 56398
0 56400 7 1 2 56388 56399
0 56401 5 1 1 56400
0 56402 7 1 2 61951 56401
0 56403 5 1 1 56402
0 56404 7 1 2 96022 98661
0 56405 5 1 1 56404
0 56406 7 1 2 56403 56405
0 56407 5 1 1 56406
0 56408 7 1 2 60737 56407
0 56409 5 1 1 56408
0 56410 7 1 2 56386 56409
0 56411 5 1 1 56410
0 56412 7 1 2 63236 56411
0 56413 5 1 1 56412
0 56414 7 1 2 56383 56413
0 56415 5 1 1 56414
0 56416 7 1 2 67785 56415
0 56417 5 1 1 56416
0 56418 7 1 2 32004 98653
0 56419 5 1 1 56418
0 56420 7 1 2 95840 56419
0 56421 5 1 1 56420
0 56422 7 1 2 56417 56421
0 56423 5 1 1 56422
0 56424 7 1 2 68564 56423
0 56425 5 1 1 56424
0 56426 7 1 2 61952 98658
0 56427 5 1 1 56426
0 56428 7 1 2 68806 56427
0 56429 7 1 2 56425 56428
0 56430 7 1 2 56369 56429
0 56431 5 1 1 56430
0 56432 7 1 2 77510 11464
0 56433 5 1 1 56432
0 56434 7 1 2 46853 56433
0 56435 5 1 1 56434
0 56436 7 1 2 89331 56435
0 56437 5 1 1 56436
0 56438 7 1 2 96026 56437
0 56439 5 1 1 56438
0 56440 7 1 2 86768 56439
0 56441 5 1 1 56440
0 56442 7 1 2 77043 96380
0 56443 5 1 1 56442
0 56444 7 1 2 63237 56443
0 56445 5 1 1 56444
0 56446 7 1 2 83511 89912
0 56447 7 1 2 56445 56446
0 56448 7 1 2 97579 56447
0 56449 5 1 1 56448
0 56450 7 1 2 63873 56449
0 56451 7 1 2 56441 56450
0 56452 5 1 1 56451
0 56453 7 1 2 64175 56452
0 56454 7 1 2 56431 56453
0 56455 5 1 1 56454
0 56456 7 1 2 56281 56455
0 56457 5 1 1 56456
0 56458 7 1 2 97767 56457
0 56459 5 1 1 56458
0 56460 7 1 2 80552 82874
0 56461 5 1 1 56460
0 56462 7 1 2 51964 56461
0 56463 5 1 1 56462
0 56464 7 1 2 84810 56463
0 56465 5 1 1 56464
0 56466 7 1 2 98402 56465
0 56467 5 1 1 56466
0 56468 7 1 2 91976 56467
0 56469 5 1 1 56468
0 56470 7 1 2 80341 86478
0 56471 5 1 1 56470
0 56472 7 1 2 56469 56471
0 56473 5 1 1 56472
0 56474 7 1 2 69033 56473
0 56475 5 1 1 56474
0 56476 7 2 2 75393 72275
0 56477 5 2 1 98662
0 56478 7 1 2 85126 98664
0 56479 5 1 1 56478
0 56480 7 1 2 92169 96601
0 56481 7 1 2 56479 56480
0 56482 5 1 1 56481
0 56483 7 1 2 56475 56482
0 56484 5 1 1 56483
0 56485 7 1 2 66928 56484
0 56486 5 1 1 56485
0 56487 7 1 2 24455 98665
0 56488 5 1 1 56487
0 56489 7 1 2 66780 56488
0 56490 5 1 1 56489
0 56491 7 1 2 39807 56490
0 56492 5 1 1 56491
0 56493 7 1 2 60960 96578
0 56494 7 1 2 56492 56493
0 56495 5 1 1 56494
0 56496 7 1 2 56486 56495
0 56497 5 1 1 56496
0 56498 7 1 2 65649 56497
0 56499 5 1 1 56498
0 56500 7 1 2 92526 98185
0 56501 5 1 1 56500
0 56502 7 1 2 40755 56501
0 56503 5 1 1 56502
0 56504 7 1 2 75370 56503
0 56505 5 1 1 56504
0 56506 7 1 2 72276 94083
0 56507 7 1 2 98320 56506
0 56508 5 1 1 56507
0 56509 7 1 2 56505 56508
0 56510 5 1 1 56509
0 56511 7 1 2 68565 56510
0 56512 5 1 1 56511
0 56513 7 1 2 96698 96810
0 56514 5 1 1 56513
0 56515 7 1 2 56512 56514
0 56516 5 1 1 56515
0 56517 7 1 2 60738 56516
0 56518 5 1 1 56517
0 56519 7 1 2 92129 98577
0 56520 7 1 2 96971 56519
0 56521 5 1 1 56520
0 56522 7 1 2 56518 56521
0 56523 5 1 1 56522
0 56524 7 1 2 60961 64176
0 56525 7 1 2 56523 56524
0 56526 5 1 1 56525
0 56527 7 1 2 56499 56526
0 56528 5 1 1 56527
0 56529 7 1 2 67395 56528
0 56530 5 1 1 56529
0 56531 7 1 2 75371 98065
0 56532 5 1 1 56531
0 56533 7 1 2 94223 98557
0 56534 5 1 1 56533
0 56535 7 1 2 56532 56534
0 56536 5 1 1 56535
0 56537 7 1 2 59991 56536
0 56538 5 1 1 56537
0 56539 7 1 2 91915 93424
0 56540 5 1 1 56539
0 56541 7 1 2 84811 91816
0 56542 5 1 1 56541
0 56543 7 1 2 56540 56542
0 56544 5 1 1 56543
0 56545 7 1 2 97408 56544
0 56546 5 1 1 56545
0 56547 7 1 2 94224 96035
0 56548 5 1 1 56547
0 56549 7 1 2 98547 51282
0 56550 5 1 1 56549
0 56551 7 1 2 59992 56550
0 56552 5 1 1 56551
0 56553 7 1 2 56548 56552
0 56554 5 1 1 56553
0 56555 7 1 2 86816 56554
0 56556 5 1 1 56555
0 56557 7 1 2 56546 56556
0 56558 7 1 2 56538 56557
0 56559 5 1 1 56558
0 56560 7 1 2 60962 64073
0 56561 7 1 2 56559 56560
0 56562 5 1 1 56561
0 56563 7 1 2 56530 56562
0 56564 5 1 1 56563
0 56565 7 1 2 67144 56564
0 56566 5 1 1 56565
0 56567 7 1 2 98396 98053
0 56568 5 1 1 56567
0 56569 7 1 2 75752 84605
0 56570 7 1 2 98056 56569
0 56571 5 1 1 56570
0 56572 7 1 2 56568 56571
0 56573 5 1 1 56572
0 56574 7 1 2 75372 56573
0 56575 5 1 1 56574
0 56576 7 1 2 68566 98364
0 56577 5 1 1 56576
0 56578 7 1 2 56575 56577
0 56579 5 1 1 56578
0 56580 7 1 2 64074 56579
0 56581 5 1 1 56580
0 56582 7 1 2 83786 75753
0 56583 5 1 1 56582
0 56584 7 1 2 71265 78974
0 56585 5 1 1 56584
0 56586 7 1 2 56583 56585
0 56587 5 1 1 56586
0 56588 7 1 2 97747 98166
0 56589 5 1 1 56588
0 56590 7 2 2 64177 80544
0 56591 7 1 2 92336 95513
0 56592 7 1 2 98666 56591
0 56593 5 1 1 56592
0 56594 7 1 2 56589 56593
0 56595 5 1 1 56594
0 56596 7 1 2 56587 56595
0 56597 5 1 1 56596
0 56598 7 1 2 96959 98559
0 56599 7 1 2 87403 56598
0 56600 5 1 1 56599
0 56601 7 1 2 56597 56600
0 56602 7 1 2 56581 56601
0 56603 7 1 2 56566 56602
0 56604 5 1 1 56603
0 56605 7 1 2 76287 56604
0 56606 5 1 1 56605
0 56607 7 1 2 69216 86773
0 56608 5 1 1 56607
0 56609 7 1 2 61138 91347
0 56610 5 1 1 56609
0 56611 7 1 2 56608 56610
0 56612 5 1 1 56611
0 56613 7 1 2 75394 56612
0 56614 5 1 1 56613
0 56615 7 1 2 94356 98124
0 56616 5 1 1 56615
0 56617 7 1 2 89492 56616
0 56618 5 1 1 56617
0 56619 7 1 2 3441 56618
0 56620 5 1 1 56619
0 56621 7 1 2 69615 56620
0 56622 5 1 1 56621
0 56623 7 1 2 56614 56622
0 56624 5 1 1 56623
0 56625 7 1 2 59993 56624
0 56626 5 1 1 56625
0 56627 7 1 2 68170 89473
0 56628 5 1 1 56627
0 56629 7 1 2 56626 56628
0 56630 5 1 1 56629
0 56631 7 1 2 86741 56630
0 56632 5 1 1 56631
0 56633 7 1 2 92981 95814
0 56634 7 1 2 97482 56633
0 56635 5 1 1 56634
0 56636 7 1 2 56632 56635
0 56637 5 1 1 56636
0 56638 7 1 2 60628 56637
0 56639 5 1 1 56638
0 56640 7 1 2 91799 92531
0 56641 5 1 1 56640
0 56642 7 1 2 56639 56641
0 56643 5 1 1 56642
0 56644 7 1 2 64178 56643
0 56645 5 1 1 56644
0 56646 7 1 2 92247 97832
0 56647 5 1 1 56646
0 56648 7 1 2 94892 96929
0 56649 5 1 1 56648
0 56650 7 1 2 56647 56649
0 56651 5 1 1 56650
0 56652 7 1 2 75121 56651
0 56653 5 1 1 56652
0 56654 7 1 2 87995 97859
0 56655 7 1 2 93268 56654
0 56656 5 1 1 56655
0 56657 7 1 2 56653 56656
0 56658 5 1 1 56657
0 56659 7 1 2 92658 56658
0 56660 5 1 1 56659
0 56661 7 1 2 63238 79866
0 56662 7 1 2 97409 56661
0 56663 5 1 1 56662
0 56664 7 1 2 56660 56663
0 56665 7 1 2 56645 56664
0 56666 5 1 1 56665
0 56667 7 1 2 59706 56666
0 56668 5 1 1 56667
0 56669 7 1 2 83116 97410
0 56670 5 1 1 56669
0 56671 7 1 2 63239 71631
0 56672 5 2 1 56671
0 56673 7 1 2 87198 98668
0 56674 5 1 1 56673
0 56675 7 1 2 73324 86742
0 56676 7 1 2 91348 56675
0 56677 5 1 1 56676
0 56678 7 1 2 56674 56677
0 56679 5 1 1 56678
0 56680 7 1 2 64179 90145
0 56681 7 1 2 56679 56680
0 56682 5 1 1 56681
0 56683 7 1 2 56670 56682
0 56684 5 1 1 56683
0 56685 7 1 2 59994 56684
0 56686 5 1 1 56685
0 56687 7 1 2 92901 96736
0 56688 7 1 2 96936 56687
0 56689 5 1 1 56688
0 56690 7 1 2 56686 56689
0 56691 5 1 1 56690
0 56692 7 1 2 75373 56691
0 56693 5 1 1 56692
0 56694 7 1 2 78139 98569
0 56695 5 1 1 56694
0 56696 7 1 2 85431 50092
0 56697 5 1 1 56696
0 56698 7 1 2 59995 98332
0 56699 7 1 2 56697 56698
0 56700 5 1 1 56699
0 56701 7 1 2 98571 56700
0 56702 5 1 1 56701
0 56703 7 1 2 61139 56702
0 56704 5 1 1 56703
0 56705 7 1 2 56695 56704
0 56706 7 1 2 56693 56705
0 56707 7 1 2 56668 56706
0 56708 5 1 1 56707
0 56709 7 1 2 61823 56708
0 56710 5 1 1 56709
0 56711 7 2 2 63599 97672
0 56712 7 1 2 82057 98670
0 56713 5 1 1 56712
0 56714 7 2 2 80745 98027
0 56715 7 1 2 78651 98672
0 56716 5 1 1 56715
0 56717 7 1 2 56713 56716
0 56718 5 1 1 56717
0 56719 7 1 2 63240 56718
0 56720 5 1 1 56719
0 56721 7 1 2 79452 98669
0 56722 5 1 1 56721
0 56723 7 1 2 79453 89184
0 56724 5 1 1 56723
0 56725 7 1 2 93241 98095
0 56726 5 1 1 56725
0 56727 7 1 2 56724 56726
0 56728 5 1 1 56727
0 56729 7 1 2 59707 56728
0 56730 5 1 1 56729
0 56731 7 1 2 56722 56730
0 56732 5 1 1 56731
0 56733 7 1 2 59996 56732
0 56734 5 1 1 56733
0 56735 7 1 2 80778 98383
0 56736 5 1 1 56735
0 56737 7 1 2 56734 56736
0 56738 5 1 1 56737
0 56739 7 1 2 95638 56738
0 56740 5 1 1 56739
0 56741 7 1 2 56720 56740
0 56742 5 1 1 56741
0 56743 7 1 2 75374 56742
0 56744 5 1 1 56743
0 56745 7 1 2 79911 98028
0 56746 5 1 1 56745
0 56747 7 2 2 96930 97477
0 56748 7 1 2 78291 84687
0 56749 7 1 2 98674 56748
0 56750 5 1 1 56749
0 56751 7 1 2 56746 56750
0 56752 5 1 1 56751
0 56753 7 1 2 69616 56752
0 56754 5 1 1 56753
0 56755 7 1 2 77935 98029
0 56756 5 2 1 56755
0 56757 7 1 2 65650 84171
0 56758 7 1 2 98520 56757
0 56759 5 1 1 56758
0 56760 7 1 2 98676 56759
0 56761 7 1 2 56754 56760
0 56762 5 1 1 56761
0 56763 7 1 2 59708 56762
0 56764 5 1 1 56763
0 56765 7 1 2 93991 98043
0 56766 5 1 1 56765
0 56767 7 1 2 56766 98677
0 56768 5 1 1 56767
0 56769 7 1 2 67145 56768
0 56770 5 1 1 56769
0 56771 7 1 2 63600 98087
0 56772 5 1 1 56771
0 56773 7 1 2 94734 95807
0 56774 7 1 2 56772 56773
0 56775 5 1 1 56774
0 56776 7 1 2 98567 56775
0 56777 5 1 1 56776
0 56778 7 1 2 61140 56777
0 56779 5 1 1 56778
0 56780 7 1 2 56770 56779
0 56781 7 1 2 56764 56780
0 56782 5 1 1 56781
0 56783 7 1 2 91729 56782
0 56784 5 1 1 56783
0 56785 7 1 2 56744 56784
0 56786 7 1 2 56710 56785
0 56787 5 1 1 56786
0 56788 7 1 2 68807 56787
0 56789 5 1 1 56788
0 56790 7 1 2 76573 53339
0 56791 5 1 1 56790
0 56792 7 1 2 91730 56791
0 56793 5 1 1 56792
0 56794 7 1 2 83253 75395
0 56795 5 1 1 56794
0 56796 7 1 2 56793 56795
0 56797 5 1 1 56796
0 56798 7 1 2 61824 56797
0 56799 5 1 1 56798
0 56800 7 1 2 79903 92822
0 56801 5 1 1 56800
0 56802 7 1 2 60414 56801
0 56803 5 1 1 56802
0 56804 7 1 2 23700 56803
0 56805 5 1 1 56804
0 56806 7 1 2 59997 56805
0 56807 5 1 1 56806
0 56808 7 1 2 75532 82557
0 56809 5 1 1 56808
0 56810 7 1 2 56807 56809
0 56811 5 1 1 56810
0 56812 7 1 2 60629 56811
0 56813 5 1 1 56812
0 56814 7 1 2 56799 56813
0 56815 5 1 1 56814
0 56816 7 1 2 65651 56815
0 56817 5 1 1 56816
0 56818 7 2 2 85686 87021
0 56819 5 1 1 98678
0 56820 7 1 2 76574 74079
0 56821 5 1 1 56820
0 56822 7 1 2 98679 56821
0 56823 5 1 1 56822
0 56824 7 1 2 56817 56823
0 56825 5 1 1 56824
0 56826 7 1 2 68171 56825
0 56827 5 1 1 56826
0 56828 7 1 2 75446 81916
0 56829 7 1 2 97968 56828
0 56830 7 1 2 97806 56829
0 56831 5 1 1 56830
0 56832 7 1 2 56827 56831
0 56833 5 1 1 56832
0 56834 7 1 2 61141 56833
0 56835 5 1 1 56834
0 56836 7 1 2 87022 88123
0 56837 5 1 1 56836
0 56838 7 1 2 98539 56837
0 56839 5 1 1 56838
0 56840 7 1 2 68567 56839
0 56841 5 1 1 56840
0 56842 7 1 2 97567 56819
0 56843 5 1 1 56842
0 56844 7 1 2 77044 78140
0 56845 7 1 2 56843 56844
0 56846 5 1 1 56845
0 56847 7 1 2 56841 56846
0 56848 5 1 1 56847
0 56849 7 1 2 71266 56848
0 56850 5 1 1 56849
0 56851 7 1 2 98278 51116
0 56852 5 1 1 56851
0 56853 7 1 2 66929 56852
0 56854 7 1 2 56850 56853
0 56855 7 1 2 56835 56854
0 56856 5 1 1 56855
0 56857 7 1 2 97125 98276
0 56858 5 1 1 56857
0 56859 7 1 2 63241 56858
0 56860 5 1 1 56859
0 56861 7 1 2 75759 17061
0 56862 5 1 1 56861
0 56863 7 1 2 59709 56862
0 56864 5 1 1 56863
0 56865 7 1 2 88919 56864
0 56866 5 1 1 56865
0 56867 7 1 2 82420 56866
0 56868 5 1 1 56867
0 56869 7 1 2 56860 56868
0 56870 5 1 1 56869
0 56871 7 1 2 63601 56870
0 56872 5 1 1 56871
0 56873 7 1 2 71267 85742
0 56874 5 1 1 56873
0 56875 7 1 2 56872 56874
0 56876 5 1 1 56875
0 56877 7 1 2 88001 56876
0 56878 5 1 1 56877
0 56879 7 1 2 61953 56878
0 56880 5 1 1 56879
0 56881 7 1 2 69034 56880
0 56882 7 1 2 56856 56881
0 56883 5 1 1 56882
0 56884 7 1 2 59710 83020
0 56885 5 2 1 56884
0 56886 7 1 2 72404 98680
0 56887 5 1 1 56886
0 56888 7 1 2 89332 56887
0 56889 5 1 1 56888
0 56890 7 1 2 79688 75396
0 56891 7 1 2 95602 56890
0 56892 5 1 1 56891
0 56893 7 1 2 56889 56892
0 56894 5 1 1 56893
0 56895 7 1 2 95639 56894
0 56896 5 1 1 56895
0 56897 7 1 2 56883 56896
0 56898 5 1 1 56897
0 56899 7 1 2 63874 56898
0 56900 5 1 1 56899
0 56901 7 1 2 89945 92982
0 56902 7 1 2 97723 56901
0 56903 5 1 1 56902
0 56904 7 1 2 42568 56903
0 56905 5 1 1 56904
0 56906 7 1 2 64180 56905
0 56907 5 1 1 56906
0 56908 7 1 2 56907 50847
0 56909 5 1 1 56908
0 56910 7 1 2 89009 56909
0 56911 5 1 1 56910
0 56912 7 1 2 64075 56911
0 56913 7 1 2 56900 56912
0 56914 7 1 2 56789 56913
0 56915 5 1 1 56914
0 56916 7 1 2 83763 74953
0 56917 5 1 1 56916
0 56918 7 1 2 65534 56917
0 56919 5 1 1 56918
0 56920 7 1 2 60415 97142
0 56921 5 1 1 56920
0 56922 7 1 2 76482 85092
0 56923 5 1 1 56922
0 56924 7 1 2 56921 56923
0 56925 5 1 1 56924
0 56926 7 1 2 69617 56925
0 56927 5 1 1 56926
0 56928 7 1 2 22193 56927
0 56929 5 1 1 56928
0 56930 7 1 2 63602 56929
0 56931 5 1 1 56930
0 56932 7 1 2 56919 56931
0 56933 5 1 1 56932
0 56934 7 1 2 97587 56933
0 56935 5 1 1 56934
0 56936 7 1 2 78150 71636
0 56937 5 2 1 56936
0 56938 7 2 2 94162 98682
0 56939 7 1 2 79966 95746
0 56940 7 1 2 98684 56939
0 56941 5 1 1 56940
0 56942 7 1 2 56935 56941
0 56943 5 1 1 56942
0 56944 7 1 2 63875 56943
0 56945 5 1 1 56944
0 56946 7 1 2 60963 81931
0 56947 5 1 1 56946
0 56948 7 1 2 84726 56947
0 56949 5 1 1 56948
0 56950 7 1 2 98533 56949
0 56951 5 1 1 56950
0 56952 7 2 2 83306 89822
0 56953 5 2 1 98686
0 56954 7 1 2 95815 98687
0 56955 5 1 1 56954
0 56956 7 1 2 56951 56955
0 56957 5 1 1 56956
0 56958 7 1 2 63603 56957
0 56959 5 1 1 56958
0 56960 7 1 2 92318 93041
0 56961 7 1 2 73057 56960
0 56962 5 1 1 56961
0 56963 7 1 2 56959 56962
0 56964 5 1 1 56963
0 56965 7 1 2 96951 56964
0 56966 5 1 1 56965
0 56967 7 1 2 56945 56966
0 56968 5 1 1 56967
0 56969 7 1 2 59711 56968
0 56970 5 1 1 56969
0 56971 7 2 2 69217 95727
0 56972 5 1 1 98690
0 56973 7 1 2 68172 84940
0 56974 5 1 1 56973
0 56975 7 1 2 63604 56974
0 56976 5 2 1 56975
0 56977 7 1 2 60416 98692
0 56978 5 1 1 56977
0 56979 7 1 2 56972 56978
0 56980 5 1 1 56979
0 56981 7 1 2 60630 87000
0 56982 7 1 2 56980 56981
0 56983 5 1 1 56982
0 56984 7 1 2 60739 85743
0 56985 5 1 1 56984
0 56986 7 1 2 56983 56985
0 56987 5 1 1 56986
0 56988 7 1 2 98221 56987
0 56989 5 1 1 56988
0 56990 7 1 2 79689 98143
0 56991 5 1 1 56990
0 56992 7 1 2 87897 92659
0 56993 7 1 2 96581 56992
0 56994 5 1 1 56993
0 56995 7 1 2 56991 56994
0 56996 5 1 1 56995
0 56997 7 1 2 90037 56996
0 56998 5 1 1 56997
0 56999 7 1 2 92341 97663
0 57000 5 1 1 56999
0 57001 7 1 2 71621 97845
0 57002 7 1 2 98222 57001
0 57003 5 1 1 57002
0 57004 7 1 2 57000 57003
0 57005 5 1 1 57004
0 57006 7 1 2 66599 57005
0 57007 5 1 1 57006
0 57008 7 2 2 60964 73054
0 57009 5 1 1 98694
0 57010 7 1 2 61142 94726
0 57011 7 1 2 98695 57010
0 57012 7 1 2 98534 57011
0 57013 5 1 1 57012
0 57014 7 1 2 57007 57013
0 57015 5 1 1 57014
0 57016 7 1 2 68173 57015
0 57017 5 1 1 57016
0 57018 7 1 2 56998 57017
0 57019 5 1 1 57018
0 57020 7 1 2 63605 57019
0 57021 5 1 1 57020
0 57022 7 1 2 91731 98693
0 57023 5 1 1 57022
0 57024 7 1 2 61618 98691
0 57025 5 1 1 57024
0 57026 7 1 2 57023 57025
0 57027 5 1 1 57026
0 57028 7 1 2 98144 57027
0 57029 5 1 1 57028
0 57030 7 1 2 88024 89905
0 57031 7 1 2 97758 57030
0 57032 5 1 1 57031
0 57033 7 1 2 57029 57032
0 57034 5 1 1 57033
0 57035 7 1 2 66781 57034
0 57036 5 1 1 57035
0 57037 7 1 2 57021 57036
0 57038 7 1 2 56989 57037
0 57039 7 1 2 56970 57038
0 57040 5 1 1 57039
0 57041 7 1 2 66930 57040
0 57042 5 1 1 57041
0 57043 7 1 2 84713 57009
0 57044 5 2 1 57043
0 57045 7 1 2 94185 98696
0 57046 5 1 1 57045
0 57047 7 1 2 98688 57046
0 57048 5 1 1 57047
0 57049 7 1 2 63606 57048
0 57050 5 1 1 57049
0 57051 7 2 2 73439 83427
0 57052 5 1 1 98698
0 57053 7 1 2 88987 57052
0 57054 5 2 1 57053
0 57055 7 1 2 61619 98700
0 57056 5 1 1 57055
0 57057 7 1 2 60631 73025
0 57058 5 1 1 57057
0 57059 7 1 2 57056 57058
0 57060 5 1 1 57059
0 57061 7 1 2 66782 57060
0 57062 5 1 1 57061
0 57063 7 1 2 57050 57062
0 57064 5 1 1 57063
0 57065 7 1 2 68808 57064
0 57066 5 1 1 57065
0 57067 7 1 2 75397 97849
0 57068 5 1 1 57067
0 57069 7 1 2 57066 57068
0 57070 5 1 1 57069
0 57071 7 1 2 68174 57070
0 57072 5 1 1 57071
0 57073 7 3 2 79690 90084
0 57074 5 1 1 98702
0 57075 7 1 2 73332 98703
0 57076 5 1 1 57075
0 57077 7 1 2 57072 57076
0 57078 5 1 1 57077
0 57079 7 1 2 87199 57078
0 57080 5 1 1 57079
0 57081 7 1 2 65652 98701
0 57082 5 1 1 57081
0 57083 7 1 2 83410 98697
0 57084 5 1 1 57083
0 57085 7 1 2 57082 57084
0 57086 5 1 1 57085
0 57087 7 1 2 89632 98067
0 57088 7 1 2 57086 57087
0 57089 5 1 1 57088
0 57090 7 1 2 57080 57089
0 57091 5 1 1 57090
0 57092 7 1 2 64181 57091
0 57093 5 1 1 57092
0 57094 7 2 2 97426 98294
0 57095 7 1 2 92163 98705
0 57096 5 1 1 57095
0 57097 7 1 2 98177 57096
0 57098 5 1 1 57097
0 57099 7 1 2 63876 57098
0 57100 5 1 1 57099
0 57101 7 2 2 62412 83573
0 57102 7 1 2 97736 98707
0 57103 7 1 2 98535 57102
0 57104 5 1 1 57103
0 57105 7 1 2 57100 57104
0 57106 5 1 1 57105
0 57107 7 1 2 66931 57106
0 57108 5 1 1 57107
0 57109 7 1 2 84593 89474
0 57110 5 1 1 57109
0 57111 7 1 2 79691 98708
0 57112 5 1 1 57111
0 57113 7 1 2 57074 57112
0 57114 7 1 2 57110 57113
0 57115 5 1 1 57114
0 57116 7 1 2 94654 97440
0 57117 7 1 2 57115 57116
0 57118 5 1 1 57117
0 57119 7 1 2 57108 57118
0 57120 5 1 1 57119
0 57121 7 1 2 70932 57120
0 57122 5 1 1 57121
0 57123 7 1 2 89404 92660
0 57124 7 1 2 95068 97664
0 57125 7 1 2 57123 57124
0 57126 5 1 1 57125
0 57127 7 1 2 57122 57126
0 57128 7 1 2 57093 57127
0 57129 5 1 1 57128
0 57130 7 1 2 59998 57129
0 57131 5 1 1 57130
0 57132 7 1 2 79934 74267
0 57133 5 1 1 57132
0 57134 7 1 2 84690 57133
0 57135 5 1 1 57134
0 57136 7 1 2 62413 79918
0 57137 7 1 2 94186 57136
0 57138 5 1 1 57137
0 57139 7 1 2 57135 57138
0 57140 5 1 1 57139
0 57141 7 1 2 61143 57140
0 57142 5 1 1 57141
0 57143 7 1 2 19897 97342
0 57144 5 1 1 57143
0 57145 7 1 2 60632 57144
0 57146 5 1 1 57145
0 57147 7 1 2 84012 94444
0 57148 5 1 1 57147
0 57149 7 1 2 98689 57148
0 57150 5 1 1 57149
0 57151 7 1 2 63607 57150
0 57152 5 1 1 57151
0 57153 7 1 2 57146 57152
0 57154 7 1 2 57142 57153
0 57155 5 1 1 57154
0 57156 7 1 2 98134 57155
0 57157 5 1 1 57156
0 57158 7 1 2 68809 96506
0 57159 7 1 2 97574 57158
0 57160 7 1 2 57157 57159
0 57161 5 1 1 57160
0 57162 7 1 2 98685 98699
0 57163 5 1 1 57162
0 57164 7 1 2 63877 57163
0 57165 5 1 1 57164
0 57166 7 1 2 64182 87152
0 57167 7 1 2 57165 57166
0 57168 7 1 2 57161 57167
0 57169 5 1 1 57168
0 57170 7 1 2 79864 6802
0 57171 5 1 1 57170
0 57172 7 1 2 76453 57171
0 57173 5 1 1 57172
0 57174 7 2 2 79932 71622
0 57175 5 1 1 98709
0 57176 7 1 2 57173 57175
0 57177 5 1 1 57176
0 57178 7 1 2 60417 96952
0 57179 7 1 2 97517 57178
0 57180 5 1 1 57179
0 57181 7 1 2 32441 57180
0 57182 5 1 1 57181
0 57183 7 1 2 57177 57182
0 57184 5 1 1 57183
0 57185 7 1 2 68969 57184
0 57186 7 1 2 57169 57185
0 57187 7 1 2 57131 57186
0 57188 7 1 2 57042 57187
0 57189 5 1 1 57188
0 57190 7 1 2 56915 57189
0 57191 5 1 1 57190
0 57192 7 1 2 56606 57191
0 57193 5 1 1 57192
0 57194 7 1 2 67786 57193
0 57195 5 1 1 57194
0 57196 7 1 2 85744 97992
0 57197 5 1 1 57196
0 57198 7 1 2 83311 53262
0 57199 5 1 1 57198
0 57200 7 1 2 72140 57199
0 57201 5 1 1 57200
0 57202 7 1 2 6518 57201
0 57203 5 1 1 57202
0 57204 7 1 2 67146 57203
0 57205 5 1 1 57204
0 57206 7 1 2 74308 74446
0 57207 5 1 1 57206
0 57208 7 1 2 57205 57207
0 57209 5 1 1 57208
0 57210 7 1 2 84812 57209
0 57211 5 1 1 57210
0 57212 7 1 2 90045 57211
0 57213 5 1 1 57212
0 57214 7 1 2 63608 57213
0 57215 5 1 1 57214
0 57216 7 1 2 57197 57215
0 57217 5 1 1 57216
0 57218 7 1 2 59999 57217
0 57219 5 1 1 57218
0 57220 7 1 2 84842 89405
0 57221 7 1 2 98080 57220
0 57222 5 1 1 57221
0 57223 7 1 2 80051 84387
0 57224 5 1 1 57223
0 57225 7 1 2 57222 57224
0 57226 7 1 2 57219 57225
0 57227 5 1 1 57226
0 57228 7 1 2 93743 57227
0 57229 5 1 1 57228
0 57230 7 1 2 95480 45213
0 57231 5 1 1 57230
0 57232 7 1 2 42547 57231
0 57233 5 1 1 57232
0 57234 7 1 2 79752 57233
0 57235 5 1 1 57234
0 57236 7 1 2 82855 95195
0 57237 5 1 1 57236
0 57238 7 1 2 4857 57237
0 57239 5 1 1 57238
0 57240 7 1 2 76288 57239
0 57241 5 1 1 57240
0 57242 7 1 2 78292 87781
0 57243 5 1 1 57242
0 57244 7 1 2 63609 57243
0 57245 5 1 1 57244
0 57246 7 1 2 61144 57245
0 57247 5 1 1 57246
0 57248 7 1 2 75242 57247
0 57249 5 1 1 57248
0 57250 7 1 2 61825 57249
0 57251 5 1 1 57250
0 57252 7 1 2 57241 57251
0 57253 5 1 1 57252
0 57254 7 1 2 60633 57253
0 57255 5 1 1 57254
0 57256 7 1 2 78384 91272
0 57257 5 2 1 57256
0 57258 7 1 2 66600 98711
0 57259 5 1 1 57258
0 57260 7 1 2 60418 57259
0 57261 5 1 1 57260
0 57262 7 3 2 74950 98083
0 57263 5 1 1 98713
0 57264 7 1 2 67147 98714
0 57265 5 1 1 57264
0 57266 7 1 2 57261 57265
0 57267 5 1 1 57266
0 57268 7 1 2 76289 57267
0 57269 5 1 1 57268
0 57270 7 1 2 35243 57269
0 57271 5 1 1 57270
0 57272 7 1 2 68568 57271
0 57273 5 1 1 57272
0 57274 7 1 2 89837 93269
0 57275 5 1 1 57274
0 57276 7 1 2 57273 57275
0 57277 7 1 2 57255 57276
0 57278 5 1 1 57277
0 57279 7 1 2 79692 57278
0 57280 5 1 1 57279
0 57281 7 1 2 88110 88091
0 57282 7 1 2 91475 57281
0 57283 5 1 1 57282
0 57284 7 1 2 57280 57283
0 57285 5 1 1 57284
0 57286 7 1 2 64076 57285
0 57287 5 1 1 57286
0 57288 7 1 2 57235 57287
0 57289 5 1 1 57288
0 57290 7 1 2 60000 57289
0 57291 5 1 1 57290
0 57292 7 1 2 80342 84884
0 57293 5 1 1 57292
0 57294 7 2 2 73333 77490
0 57295 5 1 1 98716
0 57296 7 1 2 15335 57295
0 57297 5 1 1 57296
0 57298 7 1 2 89406 57297
0 57299 5 1 1 57298
0 57300 7 1 2 79895 84388
0 57301 5 1 1 57300
0 57302 7 1 2 57299 57301
0 57303 5 1 1 57302
0 57304 7 1 2 76290 57303
0 57305 5 1 1 57304
0 57306 7 1 2 66601 42390
0 57307 5 1 1 57306
0 57308 7 1 2 82188 57307
0 57309 5 1 1 57308
0 57310 7 1 2 82191 97109
0 57311 5 1 1 57310
0 57312 7 1 2 60419 57311
0 57313 5 1 1 57312
0 57314 7 1 2 15019 57313
0 57315 7 1 2 57309 57314
0 57316 7 1 2 57305 57315
0 57317 5 1 1 57316
0 57318 7 1 2 66783 57317
0 57319 5 1 1 57318
0 57320 7 1 2 57293 57319
0 57321 5 1 1 57320
0 57322 7 1 2 68970 57321
0 57323 5 1 1 57322
0 57324 7 1 2 91851 98081
0 57325 5 1 1 57324
0 57326 7 1 2 63610 89151
0 57327 5 1 1 57326
0 57328 7 1 2 93189 57327
0 57329 5 1 1 57328
0 57330 7 1 2 57325 57329
0 57331 5 1 1 57330
0 57332 7 1 2 61826 57331
0 57333 5 1 1 57332
0 57334 7 1 2 90130 94518
0 57335 5 1 1 57334
0 57336 7 1 2 57333 57335
0 57337 5 1 1 57336
0 57338 7 1 2 64077 57337
0 57339 5 1 1 57338
0 57340 7 1 2 57323 57339
0 57341 7 1 2 57291 57340
0 57342 5 1 1 57341
0 57343 7 1 2 66932 57342
0 57344 5 1 1 57343
0 57345 7 1 2 57229 57344
0 57346 5 1 1 57345
0 57347 7 1 2 63878 57346
0 57348 5 1 1 57347
0 57349 7 1 2 73334 85499
0 57350 5 1 1 57349
0 57351 7 1 2 84392 57350
0 57352 5 1 1 57351
0 57353 7 1 2 73370 57352
0 57354 5 1 1 57353
0 57355 7 1 2 59712 91791
0 57356 5 1 1 57355
0 57357 7 1 2 65309 57356
0 57358 5 1 1 57357
0 57359 7 1 2 85500 57358
0 57360 5 1 1 57359
0 57361 7 1 2 68569 57360
0 57362 7 1 2 57354 57361
0 57363 5 1 1 57362
0 57364 7 1 2 65310 91548
0 57365 5 1 1 57364
0 57366 7 1 2 82421 57365
0 57367 5 1 1 57366
0 57368 7 1 2 75760 21884
0 57369 5 1 1 57368
0 57370 7 1 2 90038 57369
0 57371 5 1 1 57370
0 57372 7 1 2 63611 57371
0 57373 7 1 2 57367 57372
0 57374 5 1 1 57373
0 57375 7 1 2 61827 57374
0 57376 7 1 2 57363 57375
0 57377 5 1 1 57376
0 57378 7 1 2 76291 95541
0 57379 7 1 2 96499 57378
0 57380 5 1 1 57379
0 57381 7 1 2 75129 93272
0 57382 5 1 1 57381
0 57383 7 1 2 80779 95953
0 57384 7 1 2 57382 57383
0 57385 5 1 1 57384
0 57386 7 1 2 57380 57385
0 57387 5 1 1 57386
0 57388 7 1 2 60001 57387
0 57389 5 1 1 57388
0 57390 7 1 2 83121 92607
0 57391 5 1 1 57390
0 57392 7 1 2 60634 75754
0 57393 7 1 2 96500 57392
0 57394 5 1 1 57393
0 57395 7 1 2 57391 57394
0 57396 7 1 2 57389 57395
0 57397 7 1 2 57377 57396
0 57398 5 1 1 57397
0 57399 7 1 2 64078 57398
0 57400 5 1 1 57399
0 57401 7 1 2 80046 80693
0 57402 5 1 1 57401
0 57403 7 1 2 57400 57402
0 57404 5 1 1 57403
0 57405 7 1 2 85716 57404
0 57406 5 1 1 57405
0 57407 7 1 2 69035 57406
0 57408 7 1 2 57348 57407
0 57409 5 1 1 57408
0 57410 7 2 2 67148 98369
0 57411 5 1 1 98718
0 57412 7 1 2 90146 92543
0 57413 7 1 2 92556 57412
0 57414 5 1 1 57413
0 57415 7 1 2 62795 73335
0 57416 7 1 2 98552 57415
0 57417 5 1 1 57416
0 57418 7 1 2 57414 57417
0 57419 5 1 1 57418
0 57420 7 1 2 68175 57419
0 57421 5 1 1 57420
0 57422 7 1 2 57411 57421
0 57423 5 1 1 57422
0 57424 7 1 2 61954 57423
0 57425 5 1 1 57424
0 57426 7 1 2 96023 96113
0 57427 5 1 1 57426
0 57428 7 1 2 57425 57427
0 57429 5 1 1 57428
0 57430 7 1 2 76292 57429
0 57431 5 1 1 57430
0 57432 7 1 2 96663 98663
0 57433 5 1 1 57432
0 57434 7 1 2 77448 47572
0 57435 5 2 1 57434
0 57436 7 1 2 94410 98720
0 57437 5 1 1 57436
0 57438 7 1 2 91603 96400
0 57439 5 1 1 57438
0 57440 7 1 2 57437 57439
0 57441 5 1 1 57440
0 57442 7 1 2 75375 57441
0 57443 5 1 1 57442
0 57444 7 1 2 79272 84573
0 57445 5 1 1 57444
0 57446 7 1 2 83878 96493
0 57447 5 1 1 57446
0 57448 7 1 2 57445 57447
0 57449 5 1 1 57448
0 57450 7 1 2 68570 57449
0 57451 5 1 1 57450
0 57452 7 1 2 57443 57451
0 57453 5 1 1 57452
0 57454 7 1 2 61955 57453
0 57455 5 1 1 57454
0 57456 7 1 2 75533 83879
0 57457 5 1 1 57456
0 57458 7 1 2 91604 90004
0 57459 5 1 1 57458
0 57460 7 1 2 57457 57459
0 57461 5 1 1 57460
0 57462 7 1 2 86979 90147
0 57463 7 1 2 57461 57462
0 57464 5 1 1 57463
0 57465 7 1 2 57455 57464
0 57466 5 1 1 57465
0 57467 7 1 2 68971 57466
0 57468 5 1 1 57467
0 57469 7 1 2 57433 57468
0 57470 7 1 2 57431 57469
0 57471 5 1 1 57470
0 57472 7 1 2 68810 57471
0 57473 5 1 1 57472
0 57474 7 2 2 75243 93273
0 57475 5 1 1 98722
0 57476 7 1 2 60635 57475
0 57477 5 1 1 57476
0 57478 7 1 2 60420 98715
0 57479 5 1 1 57478
0 57480 7 1 2 57477 57479
0 57481 5 1 1 57480
0 57482 7 1 2 61828 57481
0 57483 5 1 1 57482
0 57484 7 1 2 88983 98683
0 57485 5 1 1 57484
0 57486 7 1 2 93274 57485
0 57487 5 1 1 57486
0 57488 7 1 2 59713 57487
0 57489 5 1 1 57488
0 57490 7 1 2 57489 98712
0 57491 5 1 1 57490
0 57492 7 1 2 94163 57491
0 57493 5 2 1 57492
0 57494 7 1 2 89308 98724
0 57495 5 1 1 57494
0 57496 7 1 2 68571 57495
0 57497 5 1 1 57496
0 57498 7 1 2 57483 57497
0 57499 5 1 1 57498
0 57500 7 1 2 96977 57499
0 57501 5 1 1 57500
0 57502 7 1 2 64183 57501
0 57503 7 1 2 57473 57502
0 57504 5 1 1 57503
0 57505 7 1 2 65653 57504
0 57506 7 1 2 57409 57505
0 57507 5 1 1 57506
0 57508 7 1 2 89306 98725
0 57509 5 1 1 57508
0 57510 7 1 2 68572 57509
0 57511 5 1 1 57510
0 57512 7 1 2 73325 97997
0 57513 5 1 1 57512
0 57514 7 1 2 66784 57263
0 57515 5 1 1 57514
0 57516 7 1 2 60636 57515
0 57517 5 1 1 57516
0 57518 7 1 2 89644 90161
0 57519 5 1 1 57518
0 57520 7 1 2 57517 57519
0 57521 5 1 1 57520
0 57522 7 1 2 60421 57521
0 57523 5 1 1 57522
0 57524 7 1 2 57513 57523
0 57525 7 1 2 57511 57524
0 57526 5 1 1 57525
0 57527 7 1 2 66933 57526
0 57528 5 1 1 57527
0 57529 7 1 2 63612 98723
0 57530 5 1 1 57529
0 57531 7 1 2 85856 85934
0 57532 7 1 2 57530 57531
0 57533 5 1 1 57532
0 57534 7 1 2 57528 57533
0 57535 5 1 1 57534
0 57536 7 1 2 94773 57535
0 57537 5 1 1 57536
0 57538 7 1 2 73489 98193
0 57539 5 1 1 57538
0 57540 7 1 2 96831 97880
0 57541 5 1 1 57540
0 57542 7 1 2 57539 57541
0 57543 5 1 1 57542
0 57544 7 1 2 80052 57543
0 57545 5 1 1 57544
0 57546 7 2 2 75398 98517
0 57547 5 1 1 98726
0 57548 7 1 2 76293 98727
0 57549 5 1 1 57548
0 57550 7 1 2 83312 83073
0 57551 5 1 1 57550
0 57552 7 1 2 76294 57551
0 57553 5 1 1 57552
0 57554 7 1 2 5428 89680
0 57555 7 1 2 57553 57554
0 57556 5 1 1 57555
0 57557 7 1 2 94735 97520
0 57558 7 1 2 57556 57557
0 57559 5 1 1 57558
0 57560 7 1 2 57549 57559
0 57561 5 1 1 57560
0 57562 7 1 2 67149 57561
0 57563 5 1 1 57562
0 57564 7 1 2 93292 98289
0 57565 5 1 1 57564
0 57566 7 1 2 93311 93518
0 57567 7 1 2 94736 57566
0 57568 5 1 1 57567
0 57569 7 1 2 57547 57568
0 57570 5 1 1 57569
0 57571 7 1 2 60002 57570
0 57572 5 1 1 57571
0 57573 7 1 2 57565 57572
0 57574 7 1 2 57563 57573
0 57575 5 1 1 57574
0 57576 7 1 2 68176 57575
0 57577 5 1 1 57576
0 57578 7 1 2 92983 98063
0 57579 5 1 1 57578
0 57580 7 1 2 75660 57579
0 57581 5 1 1 57580
0 57582 7 1 2 98518 57581
0 57583 5 1 1 57582
0 57584 7 1 2 82875 88124
0 57585 7 1 2 96931 57584
0 57586 7 1 2 97993 57585
0 57587 5 1 1 57586
0 57588 7 1 2 57583 57587
0 57589 5 1 1 57588
0 57590 7 1 2 68573 57589
0 57591 5 1 1 57590
0 57592 7 1 2 88125 95084
0 57593 7 2 2 98352 57592
0 57594 5 1 1 98728
0 57595 7 1 2 97840 98198
0 57596 5 1 1 57595
0 57597 7 1 2 57594 57596
0 57598 5 1 1 57597
0 57599 7 1 2 76454 57598
0 57600 5 1 1 57599
0 57601 7 1 2 92622 97441
0 57602 5 1 1 57601
0 57603 7 1 2 60003 98729
0 57604 5 1 1 57603
0 57605 7 1 2 57602 57604
0 57606 7 1 2 57600 57605
0 57607 7 1 2 57591 57606
0 57608 7 1 2 57577 57607
0 57609 5 1 1 57608
0 57610 7 1 2 64079 57609
0 57611 5 1 1 57610
0 57612 7 1 2 57545 57611
0 57613 7 1 2 57537 57612
0 57614 5 1 1 57613
0 57615 7 1 2 63879 57614
0 57616 5 1 1 57615
0 57617 7 1 2 79859 92557
0 57618 7 1 2 96176 57617
0 57619 5 1 1 57618
0 57620 7 1 2 73336 85873
0 57621 7 1 2 98553 57620
0 57622 5 1 1 57621
0 57623 7 1 2 57619 57622
0 57624 5 1 1 57623
0 57625 7 1 2 68177 57624
0 57626 5 1 1 57625
0 57627 7 1 2 66934 98719
0 57628 5 1 1 57627
0 57629 7 1 2 57626 57628
0 57630 5 1 1 57629
0 57631 7 1 2 76295 57630
0 57632 5 1 1 57631
0 57633 7 2 2 61956 95443
0 57634 5 1 1 98730
0 57635 7 1 2 66935 84606
0 57636 5 1 1 57635
0 57637 7 1 2 76575 98681
0 57638 5 2 1 57637
0 57639 7 2 2 69218 77491
0 57640 5 1 1 98734
0 57641 7 1 2 98732 98735
0 57642 5 1 1 57641
0 57643 7 1 2 57636 57642
0 57644 5 1 1 57643
0 57645 7 1 2 92984 57644
0 57646 5 1 1 57645
0 57647 7 1 2 75534 95444
0 57648 5 1 1 57647
0 57649 7 1 2 57646 57648
0 57650 5 1 1 57649
0 57651 7 1 2 60637 57650
0 57652 5 1 1 57651
0 57653 7 1 2 57634 57652
0 57654 5 1 1 57653
0 57655 7 1 2 64080 57654
0 57656 5 1 1 57655
0 57657 7 1 2 84574 94545
0 57658 5 1 1 57657
0 57659 7 1 2 57656 57658
0 57660 5 1 1 57659
0 57661 7 1 2 61829 57660
0 57662 5 1 1 57661
0 57663 7 1 2 84607 94647
0 57664 5 1 1 57663
0 57665 7 1 2 76352 77492
0 57666 7 1 2 96857 57665
0 57667 5 1 1 57666
0 57668 7 1 2 57664 57667
0 57669 5 1 1 57668
0 57670 7 1 2 69618 57669
0 57671 5 1 1 57670
0 57672 7 1 2 97786 98476
0 57673 5 1 1 57672
0 57674 7 1 2 33569 57673
0 57675 5 1 1 57674
0 57676 7 1 2 71428 57675
0 57677 5 1 1 57676
0 57678 7 1 2 57671 57677
0 57679 5 1 1 57678
0 57680 7 1 2 67396 57679
0 57681 5 1 1 57680
0 57682 7 1 2 84172 87305
0 57683 5 1 1 57682
0 57684 7 1 2 57681 57683
0 57685 5 1 1 57684
0 57686 7 1 2 92985 57685
0 57687 5 1 1 57686
0 57688 7 1 2 83880 94648
0 57689 5 1 1 57688
0 57690 7 1 2 64081 98731
0 57691 5 1 1 57690
0 57692 7 1 2 57689 57691
0 57693 5 1 1 57692
0 57694 7 1 2 91732 57693
0 57695 5 1 1 57694
0 57696 7 1 2 68574 57695
0 57697 7 1 2 57687 57696
0 57698 7 1 2 57662 57697
0 57699 5 1 1 57698
0 57700 7 1 2 77120 91560
0 57701 7 1 2 98321 57700
0 57702 5 1 1 57701
0 57703 7 1 2 98318 57702
0 57704 5 1 1 57703
0 57705 7 1 2 64082 57704
0 57706 5 1 1 57705
0 57707 7 1 2 86189 94164
0 57708 7 1 2 98721 57707
0 57709 5 1 1 57708
0 57710 7 1 2 63613 57709
0 57711 7 1 2 57706 57710
0 57712 5 1 1 57711
0 57713 7 1 2 57699 57712
0 57714 5 1 1 57713
0 57715 7 1 2 57632 57714
0 57716 5 1 1 57715
0 57717 7 1 2 94727 57716
0 57718 5 1 1 57717
0 57719 7 1 2 57616 57718
0 57720 5 1 1 57719
0 57721 7 1 2 60740 57720
0 57722 5 1 1 57721
0 57723 7 2 2 67397 64184
0 57724 7 2 2 96524 98736
0 57725 5 1 1 98738
0 57726 7 1 2 60965 98739
0 57727 5 1 1 57726
0 57728 7 3 2 76655 97759
0 57729 7 1 2 91889 92871
0 57730 7 1 2 98740 57729
0 57731 5 1 1 57730
0 57732 7 1 2 57727 57731
0 57733 5 1 1 57732
0 57734 7 1 2 59714 57733
0 57735 5 1 1 57734
0 57736 7 1 2 91890 96423
0 57737 7 1 2 98741 57736
0 57738 5 1 1 57737
0 57739 7 1 2 57725 57738
0 57740 5 1 1 57739
0 57741 7 1 2 61145 57740
0 57742 5 1 1 57741
0 57743 7 1 2 57735 57742
0 57744 5 1 1 57743
0 57745 7 1 2 69619 57744
0 57746 5 1 1 57745
0 57747 7 1 2 79981 96565
0 57748 7 1 2 98742 57747
0 57749 5 1 1 57748
0 57750 7 1 2 57746 57749
0 57751 5 1 1 57750
0 57752 7 1 2 79912 57751
0 57753 5 1 1 57752
0 57754 7 1 2 90162 96566
0 57755 7 1 2 98379 98003
0 57756 7 1 2 57754 57755
0 57757 5 1 1 57756
0 57758 7 1 2 53231 57757
0 57759 5 1 1 57758
0 57760 7 1 2 62164 57759
0 57761 5 1 1 57760
0 57762 7 1 2 98500 57761
0 57763 7 1 2 57753 57762
0 57764 5 1 1 57763
0 57765 7 1 2 64083 57764
0 57766 5 1 1 57765
0 57767 7 1 2 76296 97869
0 57768 5 1 1 57767
0 57769 7 1 2 10187 57768
0 57770 5 1 1 57769
0 57771 7 1 2 93270 98667
0 57772 7 1 2 57770 57771
0 57773 5 1 1 57772
0 57774 7 1 2 57766 57773
0 57775 5 1 1 57774
0 57776 7 1 2 75535 57775
0 57777 5 1 1 57776
0 57778 7 1 2 81543 69219
0 57779 7 1 2 92874 57778
0 57780 7 1 2 92986 97891
0 57781 7 1 2 57779 57780
0 57782 7 1 2 98733 57781
0 57783 5 1 1 57782
0 57784 7 1 2 57777 57783
0 57785 5 1 1 57784
0 57786 7 1 2 60638 57785
0 57787 5 1 1 57786
0 57788 7 1 2 85350 86328
0 57789 7 1 2 98387 57788
0 57790 5 1 1 57789
0 57791 7 1 2 94490 95721
0 57792 5 1 1 57791
0 57793 7 1 2 66936 76193
0 57794 7 1 2 93840 57793
0 57795 5 1 1 57794
0 57796 7 1 2 57792 57795
0 57797 5 1 1 57796
0 57798 7 1 2 69036 86388
0 57799 7 1 2 57797 57798
0 57800 5 1 1 57799
0 57801 7 1 2 57790 57800
0 57802 5 1 1 57801
0 57803 7 1 2 66785 57802
0 57804 5 1 1 57803
0 57805 7 1 2 79896 96944
0 57806 5 1 1 57805
0 57807 7 1 2 50917 57806
0 57808 5 1 1 57807
0 57809 7 1 2 60422 57808
0 57810 5 1 1 57809
0 57811 7 1 2 85924 96602
0 57812 5 1 1 57811
0 57813 7 1 2 57810 57812
0 57814 5 1 1 57813
0 57815 7 1 2 60639 94257
0 57816 7 1 2 57814 57815
0 57817 5 1 1 57816
0 57818 7 1 2 57804 57817
0 57819 5 1 1 57818
0 57820 7 1 2 78311 57819
0 57821 5 1 1 57820
0 57822 7 1 2 94258 97391
0 57823 7 1 2 92860 57822
0 57824 5 1 1 57823
0 57825 7 1 2 96220 98324
0 57826 7 1 2 96438 57825
0 57827 5 1 1 57826
0 57828 7 1 2 57824 57827
0 57829 5 1 1 57828
0 57830 7 1 2 68811 57829
0 57831 5 1 1 57830
0 57832 7 1 2 65654 57831
0 57833 7 1 2 57821 57832
0 57834 5 1 1 57833
0 57835 7 1 2 73490 98515
0 57836 5 1 1 57835
0 57837 7 1 2 79454 98496
0 57838 5 1 1 57837
0 57839 7 1 2 96441 57838
0 57840 5 1 1 57839
0 57841 7 1 2 86190 92234
0 57842 7 1 2 57840 57841
0 57843 5 1 1 57842
0 57844 7 1 2 57836 57843
0 57845 5 1 1 57844
0 57846 7 1 2 64185 57845
0 57847 5 1 1 57846
0 57848 7 1 2 92572 94231
0 57849 7 1 2 98084 57848
0 57850 7 1 2 98342 57849
0 57851 5 1 1 57850
0 57852 7 1 2 60741 57851
0 57853 7 1 2 57847 57852
0 57854 5 1 1 57853
0 57855 7 1 2 71268 57854
0 57856 7 1 2 57834 57855
0 57857 5 1 1 57856
0 57858 7 1 2 57787 57857
0 57859 7 1 2 57722 57858
0 57860 7 1 2 57507 57859
0 57861 7 1 2 57195 57860
0 57862 5 1 1 57861
0 57863 7 1 2 95325 57862
0 57864 5 1 1 57863
0 57865 7 1 2 75101 90363
0 57866 5 1 1 57865
0 57867 7 1 2 74309 88907
0 57868 5 1 1 57867
0 57869 7 1 2 57866 57868
0 57870 5 2 1 57869
0 57871 7 1 2 80148 98743
0 57872 5 1 1 57871
0 57873 7 1 2 60004 90918
0 57874 5 1 1 57873
0 57875 7 1 2 71140 76330
0 57876 5 1 1 57875
0 57877 7 1 2 59715 69330
0 57878 7 1 2 57876 57877
0 57879 5 1 1 57878
0 57880 7 1 2 57874 57879
0 57881 5 1 1 57880
0 57882 7 1 2 65655 75399
0 57883 7 1 2 57881 57882
0 57884 5 1 1 57883
0 57885 7 1 2 57872 57884
0 57886 5 1 1 57885
0 57887 7 1 2 68178 57886
0 57888 5 1 1 57887
0 57889 7 1 2 71669 76567
0 57890 7 1 2 74956 57889
0 57891 7 1 2 85378 57890
0 57892 5 1 1 57891
0 57893 7 1 2 89546 89088
0 57894 5 1 1 57893
0 57895 7 1 2 75661 57894
0 57896 5 1 1 57895
0 57897 7 1 2 59716 92287
0 57898 7 1 2 57896 57897
0 57899 5 1 1 57898
0 57900 7 1 2 57892 57899
0 57901 7 1 2 57888 57900
0 57902 5 1 1 57901
0 57903 7 1 2 96464 57902
0 57904 5 1 1 57903
0 57905 7 1 2 92474 98088
0 57906 5 1 1 57905
0 57907 7 1 2 73832 57906
0 57908 5 1 1 57907
0 57909 7 1 2 59717 83996
0 57910 5 1 1 57909
0 57911 7 1 2 63242 57910
0 57912 5 1 1 57911
0 57913 7 1 2 71901 57912
0 57914 5 1 1 57913
0 57915 7 1 2 89006 57914
0 57916 7 1 2 57908 57915
0 57917 5 1 1 57916
0 57918 7 1 2 98704 57917
0 57919 5 1 1 57918
0 57920 7 1 2 60005 98132
0 57921 5 1 1 57920
0 57922 7 1 2 78141 89041
0 57923 5 1 1 57922
0 57924 7 1 2 57921 57923
0 57925 5 1 1 57924
0 57926 7 1 2 59718 57925
0 57927 5 1 1 57926
0 57928 7 1 2 72277 97827
0 57929 5 1 1 57928
0 57930 7 1 2 57927 57929
0 57931 5 1 1 57930
0 57932 7 1 2 75376 57931
0 57933 5 1 1 57932
0 57934 7 1 2 39571 57933
0 57935 5 1 1 57934
0 57936 7 1 2 66786 57935
0 57937 5 1 1 57936
0 57938 7 1 2 59719 91414
0 57939 5 1 1 57938
0 57940 7 1 2 68575 57939
0 57941 7 1 2 57937 57940
0 57942 5 1 1 57941
0 57943 7 1 2 68179 94187
0 57944 7 1 2 98744 57943
0 57945 5 1 1 57944
0 57946 7 2 2 81459 90492
0 57947 5 1 1 98745
0 57948 7 1 2 94188 98746
0 57949 5 1 1 57948
0 57950 7 1 2 94157 57949
0 57951 5 1 1 57950
0 57952 7 1 2 63243 57951
0 57953 5 1 1 57952
0 57954 7 1 2 63614 57953
0 57955 7 1 2 57945 57954
0 57956 5 1 1 57955
0 57957 7 1 2 68812 57956
0 57958 7 1 2 57942 57957
0 57959 5 1 1 57958
0 57960 7 1 2 57919 57959
0 57961 5 1 1 57960
0 57962 7 1 2 86817 57961
0 57963 5 1 1 57962
0 57964 7 1 2 57904 57963
0 57965 5 1 1 57964
0 57966 7 1 2 64186 57965
0 57967 5 1 1 57966
0 57968 7 1 2 66602 97364
0 57969 5 1 1 57968
0 57970 7 2 2 75377 84885
0 57971 5 1 1 98747
0 57972 7 1 2 90568 57971
0 57973 5 1 1 57972
0 57974 7 1 2 67150 57973
0 57975 5 1 1 57974
0 57976 7 1 2 57969 57975
0 57977 5 1 1 57976
0 57978 7 1 2 61146 57977
0 57979 5 1 1 57978
0 57980 7 1 2 71362 96708
0 57981 5 1 1 57980
0 57982 7 1 2 82620 14869
0 57983 5 1 1 57982
0 57984 7 1 2 65535 57983
0 57985 5 1 1 57984
0 57986 7 1 2 74744 57640
0 57987 5 1 1 57986
0 57988 7 1 2 89407 57987
0 57989 5 1 1 57988
0 57990 7 1 2 57985 57989
0 57991 5 1 1 57990
0 57992 7 1 2 67151 57991
0 57993 5 1 1 57992
0 57994 7 1 2 57981 57993
0 57995 7 1 2 57979 57994
0 57996 5 1 1 57995
0 57997 7 1 2 60006 57996
0 57998 5 1 1 57997
0 57999 7 1 2 91558 96709
0 58000 5 1 1 57999
0 58001 7 1 2 83197 95682
0 58002 5 1 1 58001
0 58003 7 1 2 58000 58002
0 58004 5 1 1 58003
0 58005 7 1 2 67787 58004
0 58006 5 1 1 58005
0 58007 7 1 2 73337 98748
0 58008 5 1 1 58007
0 58009 7 2 2 63244 71637
0 58010 5 2 1 98749
0 58011 7 1 2 98200 98751
0 58012 5 1 1 58011
0 58013 7 1 2 58008 58012
0 58014 7 1 2 58006 58013
0 58015 5 1 1 58014
0 58016 7 1 2 67152 58015
0 58017 5 1 1 58016
0 58018 7 1 2 67398 71902
0 58019 5 1 1 58018
0 58020 7 1 2 89831 58019
0 58021 5 1 1 58020
0 58022 7 1 2 96710 58021
0 58023 5 1 1 58022
0 58024 7 1 2 15416 58023
0 58025 7 1 2 58017 58024
0 58026 7 1 2 57998 58025
0 58027 5 1 1 58026
0 58028 7 1 2 86574 97588
0 58029 7 1 2 58027 58028
0 58030 5 1 1 58029
0 58031 7 1 2 57967 58030
0 58032 5 1 1 58031
0 58033 7 1 2 95326 58032
0 58034 5 1 1 58033
0 58035 7 1 2 73833 96789
0 58036 5 1 1 58035
0 58037 7 1 2 77015 88960
0 58038 5 1 1 58037
0 58039 7 1 2 58036 58038
0 58040 5 1 1 58039
0 58041 7 1 2 59720 58040
0 58042 5 1 1 58041
0 58043 7 1 2 91077 12884
0 58044 5 1 1 58043
0 58045 7 1 2 67153 58044
0 58046 5 1 1 58045
0 58047 7 1 2 91953 58046
0 58048 7 1 2 58042 58047
0 58049 5 1 1 58048
0 58050 7 1 2 97031 58049
0 58051 5 1 1 58050
0 58052 7 1 2 58034 58051
0 58053 5 1 1 58052
0 58054 7 1 2 68972 58053
0 58055 5 1 1 58054
0 58056 7 1 2 83208 57947
0 58057 5 1 1 58056
0 58058 7 1 2 68180 58057
0 58059 5 1 1 58058
0 58060 7 1 2 70545 88908
0 58061 5 1 1 58060
0 58062 7 1 2 13804 58061
0 58063 5 1 1 58062
0 58064 7 1 2 68576 58063
0 58065 5 1 1 58064
0 58066 7 1 2 58059 58065
0 58067 5 1 1 58066
0 58068 7 1 2 75378 58067
0 58069 5 1 1 58068
0 58070 7 1 2 83344 75755
0 58071 7 1 2 92403 58070
0 58072 5 1 1 58071
0 58073 7 1 2 71638 96466
0 58074 5 4 1 58073
0 58075 7 1 2 75536 98753
0 58076 5 1 1 58075
0 58077 7 1 2 58072 58076
0 58078 7 1 2 58069 58077
0 58079 5 1 1 58078
0 58080 7 1 2 79693 58079
0 58081 5 1 1 58080
0 58082 7 1 2 79860 91476
0 58083 7 1 2 94395 58082
0 58084 5 1 1 58083
0 58085 7 1 2 80894 98754
0 58086 5 1 1 58085
0 58087 7 1 2 58084 58086
0 58088 7 1 2 58081 58087
0 58089 5 1 1 58088
0 58090 7 1 2 61957 58089
0 58091 5 1 1 58090
0 58092 7 1 2 60640 73326
0 58093 7 2 2 92721 58092
0 58094 7 1 2 82618 96946
0 58095 7 1 2 98757 58094
0 58096 5 1 1 58095
0 58097 7 1 2 58091 58096
0 58098 5 1 1 58097
0 58099 7 1 2 60742 58098
0 58100 5 1 1 58099
0 58101 7 1 2 92139 96683
0 58102 7 1 2 98758 58101
0 58103 5 1 1 58102
0 58104 7 1 2 64187 58103
0 58105 7 1 2 58100 58104
0 58106 5 1 1 58105
0 58107 7 1 2 83079 95728
0 58108 5 1 1 58107
0 58109 7 1 2 14914 58108
0 58110 5 1 1 58109
0 58111 7 1 2 75379 58110
0 58112 5 1 1 58111
0 58113 7 1 2 41476 58112
0 58114 5 1 1 58113
0 58115 7 1 2 60641 58114
0 58116 5 1 1 58115
0 58117 7 1 2 60966 61830
0 58118 7 1 2 98385 58117
0 58119 5 1 1 58118
0 58120 7 1 2 58116 58119
0 58121 5 1 1 58120
0 58122 7 1 2 86732 58121
0 58123 5 1 1 58122
0 58124 7 1 2 62165 74154
0 58125 5 1 1 58124
0 58126 7 1 2 74745 58125
0 58127 5 1 1 58126
0 58128 7 1 2 93271 58127
0 58129 5 1 1 58128
0 58130 7 1 2 94039 58129
0 58131 5 1 1 58130
0 58132 7 1 2 87200 58131
0 58133 5 1 1 58132
0 58134 7 1 2 71670 86244
0 58135 7 1 2 90015 58134
0 58136 7 1 2 97532 58135
0 58137 5 1 1 58136
0 58138 7 1 2 58133 58137
0 58139 5 1 1 58138
0 58140 7 1 2 85687 58139
0 58141 5 1 1 58140
0 58142 7 1 2 69037 58141
0 58143 7 1 2 58123 58142
0 58144 5 1 1 58143
0 58145 7 1 2 63880 58144
0 58146 7 1 2 58106 58145
0 58147 5 1 1 58146
0 58148 7 1 2 63881 98316
0 58149 5 1 1 58148
0 58150 7 1 2 75031 84874
0 58151 5 1 1 58150
0 58152 7 1 2 58149 58151
0 58153 5 1 1 58152
0 58154 7 1 2 78267 58153
0 58155 5 1 1 58154
0 58156 7 1 2 81544 79235
0 58157 5 1 1 58156
0 58158 7 1 2 58155 58157
0 58159 5 1 1 58158
0 58160 7 1 2 61831 58159
0 58161 5 1 1 58160
0 58162 7 1 2 75662 98314
0 58163 5 1 1 58162
0 58164 7 1 2 93722 58163
0 58165 5 1 1 58164
0 58166 7 1 2 68181 74665
0 58167 5 1 1 58166
0 58168 7 1 2 63615 58167
0 58169 5 1 1 58168
0 58170 7 1 2 84370 91733
0 58171 7 1 2 58169 58170
0 58172 5 1 1 58171
0 58173 7 1 2 58165 58172
0 58174 7 1 2 58161 58173
0 58175 5 1 1 58174
0 58176 7 1 2 60007 58175
0 58177 5 1 1 58176
0 58178 7 1 2 84414 89870
0 58179 5 1 1 58178
0 58180 7 1 2 83852 95542
0 58181 5 1 1 58180
0 58182 7 1 2 58179 58181
0 58183 7 1 2 98541 58182
0 58184 5 1 1 58183
0 58185 7 1 2 68577 58184
0 58186 5 1 1 58185
0 58187 7 2 2 75380 97536
0 58188 7 1 2 89697 98759
0 58189 5 1 1 58188
0 58190 7 1 2 58186 58189
0 58191 7 1 2 58177 58190
0 58192 5 1 1 58191
0 58193 7 1 2 97411 58192
0 58194 5 1 1 58193
0 58195 7 1 2 96610 51541
0 58196 5 1 1 58195
0 58197 7 1 2 75400 58196
0 58198 5 1 1 58197
0 58199 7 1 2 92764 96808
0 58200 5 1 1 58199
0 58201 7 1 2 58198 58200
0 58202 5 1 1 58201
0 58203 7 1 2 67154 58202
0 58204 5 1 1 58203
0 58205 7 1 2 74898 91817
0 58206 5 1 1 58205
0 58207 7 1 2 58204 58206
0 58208 5 1 1 58207
0 58209 7 1 2 61958 58208
0 58210 5 1 1 58209
0 58211 7 1 2 92261 96802
0 58212 5 1 1 58211
0 58213 7 1 2 58210 58212
0 58214 5 1 1 58213
0 58215 7 1 2 60743 58214
0 58216 5 1 1 58215
0 58217 7 1 2 74265 96152
0 58218 7 1 2 89346 58217
0 58219 7 1 2 92765 58218
0 58220 5 1 1 58219
0 58221 7 1 2 58216 58220
0 58222 5 1 1 58221
0 58223 7 1 2 64188 58222
0 58224 5 1 1 58223
0 58225 7 1 2 80895 98366
0 58226 5 1 1 58225
0 58227 7 1 2 98565 58226
0 58228 5 1 1 58227
0 58229 7 1 2 75122 58228
0 58230 5 1 1 58229
0 58231 7 1 2 82278 98545
0 58232 5 1 1 58231
0 58233 7 1 2 58230 58232
0 58234 5 1 1 58233
0 58235 7 1 2 86818 58234
0 58236 5 1 1 58235
0 58237 7 1 2 58224 58236
0 58238 7 1 2 58194 58237
0 58239 5 1 1 58238
0 58240 7 1 2 71605 58239
0 58241 5 1 1 58240
0 58242 7 1 2 67788 79960
0 58243 5 1 1 58242
0 58244 7 1 2 98333 58243
0 58245 7 1 2 89037 58244
0 58246 5 1 1 58245
0 58247 7 1 2 70503 92219
0 58248 5 1 1 58247
0 58249 7 1 2 61147 77128
0 58250 5 1 1 58249
0 58251 7 1 2 58248 58250
0 58252 5 1 1 58251
0 58253 7 1 2 60967 58252
0 58254 5 1 1 58253
0 58255 7 1 2 70504 90493
0 58256 5 1 1 58255
0 58257 7 1 2 58254 58256
0 58258 5 1 1 58257
0 58259 7 1 2 96527 98325
0 58260 7 1 2 58258 58259
0 58261 5 1 1 58260
0 58262 7 1 2 58246 58261
0 58263 5 1 1 58262
0 58264 7 1 2 63245 58263
0 58265 5 1 1 58264
0 58266 7 1 2 91765 98737
0 58267 7 1 2 74770 58266
0 58268 7 1 2 98312 58267
0 58269 5 1 1 58268
0 58270 7 1 2 94204 96932
0 58271 5 1 1 58270
0 58272 7 1 2 68578 58271
0 58273 7 1 2 58269 58272
0 58274 7 1 2 58265 58273
0 58275 5 1 1 58274
0 58276 7 1 2 72278 98303
0 58277 5 1 1 58276
0 58278 7 1 2 78202 86733
0 58279 7 1 2 98353 58278
0 58280 5 1 1 58279
0 58281 7 1 2 58277 58280
0 58282 5 1 1 58281
0 58283 7 1 2 76417 58282
0 58284 5 1 1 58283
0 58285 7 1 2 60008 95570
0 58286 5 1 1 58285
0 58287 7 1 2 98750 58286
0 58288 5 1 1 58287
0 58289 7 1 2 59721 90955
0 58290 7 1 2 58288 58289
0 58291 5 1 1 58290
0 58292 7 1 2 78277 58291
0 58293 5 1 1 58292
0 58294 7 1 2 98304 58293
0 58295 5 1 1 58294
0 58296 7 1 2 63616 58295
0 58297 7 1 2 58284 58296
0 58298 5 1 1 58297
0 58299 7 1 2 61832 58298
0 58300 7 1 2 58275 58299
0 58301 5 1 1 58300
0 58302 7 1 2 76418 98671
0 58303 5 1 1 58302
0 58304 7 1 2 75779 98673
0 58305 5 1 1 58304
0 58306 7 1 2 58303 58305
0 58307 5 1 1 58306
0 58308 7 1 2 63246 58307
0 58309 5 1 1 58308
0 58310 7 1 2 74771 95640
0 58311 5 1 1 58310
0 58312 7 1 2 76568 78293
0 58313 7 1 2 98675 58312
0 58314 5 1 1 58313
0 58315 7 1 2 58311 58314
0 58316 5 1 1 58315
0 58317 7 1 2 68579 84688
0 58318 7 1 2 58316 58317
0 58319 5 1 1 58318
0 58320 7 1 2 58309 58319
0 58321 5 1 1 58320
0 58322 7 1 2 67789 58321
0 58323 5 1 1 58322
0 58324 7 1 2 79861 98030
0 58325 7 1 2 98717 58324
0 58326 5 1 1 58325
0 58327 7 1 2 58323 58326
0 58328 5 1 1 58327
0 58329 7 1 2 75381 58328
0 58330 5 1 1 58329
0 58331 7 1 2 97922 98755
0 58332 5 1 1 58331
0 58333 7 1 2 60009 90920
0 58334 5 1 1 58333
0 58335 7 1 2 75032 98756
0 58336 5 1 1 58335
0 58337 7 1 2 78278 58336
0 58338 7 1 2 58334 58337
0 58339 5 1 1 58338
0 58340 7 1 2 97918 58339
0 58341 5 1 1 58340
0 58342 7 1 2 58332 58341
0 58343 5 1 1 58342
0 58344 7 1 2 91734 58343
0 58345 5 1 1 58344
0 58346 7 1 2 58330 58345
0 58347 7 1 2 58301 58346
0 58348 5 1 1 58347
0 58349 7 1 2 68813 58348
0 58350 5 1 1 58349
0 58351 7 1 2 73338 93984
0 58352 7 1 2 96161 58351
0 58353 5 1 1 58352
0 58354 7 1 2 53264 58353
0 58355 5 1 1 58354
0 58356 7 1 2 66603 58355
0 58357 5 1 1 58356
0 58358 7 1 2 79295 91897
0 58359 7 1 2 93312 58358
0 58360 5 1 1 58359
0 58361 7 1 2 95096 95986
0 58362 7 1 2 58360 58361
0 58363 5 1 1 58362
0 58364 7 1 2 66937 91735
0 58365 7 1 2 58363 58364
0 58366 5 1 1 58365
0 58367 7 1 2 58357 58366
0 58368 5 1 1 58367
0 58369 7 1 2 67155 58368
0 58370 5 1 1 58369
0 58371 7 1 2 84453 98710
0 58372 5 1 1 58371
0 58373 7 1 2 89699 58372
0 58374 5 1 1 58373
0 58375 7 1 2 98760 58374
0 58376 5 1 1 58375
0 58377 7 1 2 84289 90163
0 58378 7 1 2 92229 58377
0 58379 5 1 1 58378
0 58380 7 1 2 58376 58379
0 58381 5 1 1 58380
0 58382 7 1 2 66938 58381
0 58383 5 1 1 58382
0 58384 7 1 2 58370 58383
0 58385 5 1 1 58384
0 58386 7 1 2 69038 58385
0 58387 5 1 1 58386
0 58388 7 1 2 67156 98287
0 58389 5 1 1 58388
0 58390 7 1 2 58387 58389
0 58391 5 1 1 58390
0 58392 7 1 2 65656 58391
0 58393 5 1 1 58392
0 58394 7 1 2 66939 98563
0 58395 5 1 1 58394
0 58396 7 1 2 96177 98367
0 58397 5 1 1 58396
0 58398 7 1 2 58395 58397
0 58399 5 1 1 58398
0 58400 7 1 2 60744 75123
0 58401 7 1 2 58399 58400
0 58402 5 1 1 58401
0 58403 7 1 2 58393 58402
0 58404 5 1 1 58403
0 58405 7 1 2 74899 58404
0 58406 5 1 1 58405
0 58407 7 1 2 58350 58406
0 58408 7 1 2 58241 58407
0 58409 7 1 2 58147 58408
0 58410 5 1 1 58409
0 58411 7 1 2 97768 58410
0 58412 5 1 1 58411
0 58413 7 1 2 58055 58412
0 58414 5 1 1 58413
0 58415 7 1 2 69966 58414
0 58416 5 1 1 58415
0 58417 7 1 2 81618 96469
0 58418 5 1 1 58417
0 58419 7 1 2 91457 58418
0 58420 5 2 1 58419
0 58421 7 1 2 98761 98267
0 58422 5 1 1 58421
0 58423 7 1 2 68182 76297
0 58424 7 1 2 96178 58423
0 58425 5 1 1 58424
0 58426 7 1 2 81917 86564
0 58427 7 1 2 97816 58426
0 58428 5 1 1 58427
0 58429 7 1 2 58425 58428
0 58430 5 1 1 58429
0 58431 7 1 2 60745 58430
0 58432 5 1 1 58431
0 58433 7 1 2 77493 95722
0 58434 7 1 2 96288 58433
0 58435 7 1 2 97359 58434
0 58436 5 1 1 58435
0 58437 7 1 2 58432 58436
0 58438 5 1 1 58437
0 58439 7 1 2 75401 58438
0 58440 5 1 1 58439
0 58441 7 1 2 67790 80006
0 58442 5 1 1 58441
0 58443 7 1 2 63247 58442
0 58444 5 1 1 58443
0 58445 7 1 2 63617 58444
0 58446 7 1 2 97580 58445
0 58447 5 1 1 58446
0 58448 7 1 2 58440 58447
0 58449 5 1 1 58448
0 58450 7 1 2 64189 58449
0 58451 5 1 1 58450
0 58452 7 1 2 77936 88984
0 58453 5 1 1 58452
0 58454 7 1 2 85432 58453
0 58455 5 1 1 58454
0 58456 7 1 2 83345 58455
0 58457 5 1 1 58456
0 58458 7 1 2 76569 85949
0 58459 5 1 1 58458
0 58460 7 1 2 58457 58459
0 58461 5 1 1 58460
0 58462 7 1 2 66604 58461
0 58463 5 1 1 58462
0 58464 7 2 2 75056 96501
0 58465 5 1 1 98763
0 58466 7 1 2 58465 52219
0 58467 7 1 2 58463 58466
0 58468 5 1 1 58467
0 58469 7 1 2 61833 58468
0 58470 5 1 1 58469
0 58471 7 1 2 41532 50536
0 58472 5 1 1 58471
0 58473 7 1 2 67791 58472
0 58474 5 1 1 58473
0 58475 7 1 2 51844 58474
0 58476 5 1 1 58475
0 58477 7 1 2 96494 58476
0 58478 5 1 1 58477
0 58479 7 1 2 83021 98381
0 58480 5 1 1 58479
0 58481 7 1 2 60642 98764
0 58482 5 1 1 58481
0 58483 7 1 2 58480 58482
0 58484 7 1 2 58478 58483
0 58485 7 1 2 58470 58484
0 58486 5 1 1 58485
0 58487 7 1 2 96933 58486
0 58488 5 1 1 58487
0 58489 7 1 2 91368 98522
0 58490 7 1 2 96485 58489
0 58491 5 1 1 58490
0 58492 7 1 2 58488 58491
0 58493 5 1 1 58492
0 58494 7 1 2 65657 58493
0 58495 5 1 1 58494
0 58496 7 1 2 58451 58495
0 58497 5 1 1 58496
0 58498 7 1 2 64084 58497
0 58499 5 1 1 58498
0 58500 7 1 2 76298 86925
0 58501 5 1 1 58500
0 58502 7 1 2 80966 96250
0 58503 5 1 1 58502
0 58504 7 1 2 58501 58503
0 58505 5 1 1 58504
0 58506 7 1 2 60010 58505
0 58507 5 1 1 58506
0 58508 7 1 2 93992 98271
0 58509 5 1 1 58508
0 58510 7 1 2 58507 58509
0 58511 5 1 1 58510
0 58512 7 1 2 68183 58511
0 58513 5 1 1 58512
0 58514 7 1 2 65658 96872
0 58515 5 1 1 58514
0 58516 7 1 2 58513 58515
0 58517 5 1 1 58516
0 58518 7 1 2 87099 58517
0 58519 5 1 1 58518
0 58520 7 1 2 74155 94189
0 58521 7 1 2 97121 58520
0 58522 5 1 1 58521
0 58523 7 1 2 79455 89547
0 58524 7 1 2 80007 58523
0 58525 5 1 1 58524
0 58526 7 1 2 58522 58525
0 58527 5 1 1 58526
0 58528 7 1 2 68184 58527
0 58529 5 1 1 58528
0 58530 7 1 2 97575 58529
0 58531 5 1 1 58530
0 58532 7 1 2 86819 58531
0 58533 5 1 1 58532
0 58534 7 1 2 58519 58533
0 58535 5 1 1 58534
0 58536 7 1 2 94774 58535
0 58537 5 1 1 58536
0 58538 7 1 2 68814 58537
0 58539 7 1 2 58499 58538
0 58540 5 1 1 58539
0 58541 7 1 2 83346 84608
0 58542 5 1 1 58541
0 58543 7 1 2 52526 58542
0 58544 5 1 1 58543
0 58545 7 1 2 79694 58544
0 58546 5 1 1 58545
0 58547 7 1 2 70294 88092
0 58548 7 1 2 97360 58547
0 58549 5 1 1 58548
0 58550 7 1 2 58546 58549
0 58551 5 1 1 58550
0 58552 7 1 2 97412 58551
0 58553 5 1 1 58552
0 58554 7 2 2 73371 98295
0 58555 7 1 2 95700 98765
0 58556 5 1 1 58555
0 58557 7 1 2 58553 58556
0 58558 5 1 1 58557
0 58559 7 1 2 64085 58558
0 58560 5 1 1 58559
0 58561 7 1 2 94775 97002
0 58562 7 1 2 98762 58561
0 58563 5 1 1 58562
0 58564 7 1 2 58560 58563
0 58565 5 1 1 58564
0 58566 7 1 2 60423 58565
0 58567 5 1 1 58566
0 58568 7 2 2 64190 81841
0 58569 7 1 2 97427 97931
0 58570 7 1 2 98767 58569
0 58571 5 1 1 58570
0 58572 7 1 2 58567 58571
0 58573 5 1 1 58572
0 58574 7 1 2 61620 58573
0 58575 5 1 1 58574
0 58576 7 1 2 96153 97978
0 58577 7 1 2 98348 58576
0 58578 5 1 1 58577
0 58579 7 1 2 81842 86543
0 58580 5 1 1 58579
0 58581 7 1 2 42551 58580
0 58582 5 1 1 58581
0 58583 7 1 2 76299 96934
0 58584 7 1 2 58582 58583
0 58585 5 1 1 58584
0 58586 7 1 2 58578 58585
0 58587 5 1 1 58586
0 58588 7 1 2 65659 58587
0 58589 5 1 1 58588
0 58590 7 1 2 83065 86191
0 58591 5 1 1 58590
0 58592 7 1 2 68973 83354
0 58593 5 1 1 58592
0 58594 7 1 2 69620 96832
0 58595 7 1 2 58593 58594
0 58596 5 1 1 58595
0 58597 7 1 2 58591 58596
0 58598 5 1 1 58597
0 58599 7 1 2 98706 58598
0 58600 5 1 1 58599
0 58601 7 1 2 58589 58600
0 58602 5 1 1 58601
0 58603 7 1 2 60011 58602
0 58604 5 1 1 58603
0 58605 7 1 2 64086 98076
0 58606 5 1 1 58605
0 58607 7 1 2 87652 98766
0 58608 5 1 1 58607
0 58609 7 1 2 49679 58608
0 58610 5 1 1 58609
0 58611 7 1 2 86820 58610
0 58612 5 1 1 58611
0 58613 7 1 2 58606 58612
0 58614 7 1 2 58604 58613
0 58615 5 1 1 58614
0 58616 7 1 2 75382 58615
0 58617 5 1 1 58616
0 58618 7 1 2 80967 98256
0 58619 7 1 2 87650 58618
0 58620 5 1 1 58619
0 58621 7 1 2 92346 96559
0 58622 5 1 1 58621
0 58623 7 1 2 75402 97500
0 58624 5 1 1 58623
0 58625 7 1 2 58622 58624
0 58626 5 1 1 58625
0 58627 7 1 2 79695 58626
0 58628 5 1 1 58627
0 58629 7 1 2 96321 58628
0 58630 5 1 1 58629
0 58631 7 1 2 67157 64191
0 58632 7 1 2 58630 58631
0 58633 5 1 1 58632
0 58634 7 1 2 58620 58633
0 58635 5 1 1 58634
0 58636 7 1 2 80008 58635
0 58637 5 1 1 58636
0 58638 7 1 2 79494 97995
0 58639 5 1 1 58638
0 58640 7 1 2 89823 96470
0 58641 7 1 2 98235 58640
0 58642 5 1 1 58641
0 58643 7 1 2 58639 58642
0 58644 5 1 1 58643
0 58645 7 1 2 76300 58644
0 58646 5 1 1 58645
0 58647 7 1 2 74900 91736
0 58648 7 1 2 98450 58647
0 58649 5 1 1 58648
0 58650 7 1 2 73956 96337
0 58651 7 1 2 84623 58650
0 58652 5 1 1 58651
0 58653 7 1 2 58649 58652
0 58654 5 1 1 58653
0 58655 7 1 2 68185 58654
0 58656 5 1 1 58655
0 58657 7 1 2 58646 58656
0 58658 5 1 1 58657
0 58659 7 1 2 86821 58658
0 58660 5 1 1 58659
0 58661 7 1 2 74901 95641
0 58662 5 2 1 58661
0 58663 7 1 2 84609 97413
0 58664 7 1 2 83892 58663
0 58665 5 1 1 58664
0 58666 7 1 2 98769 58665
0 58667 5 1 1 58666
0 58668 7 1 2 59722 58667
0 58669 5 1 1 58668
0 58670 7 1 2 74106 95642
0 58671 5 1 1 58670
0 58672 7 1 2 58669 58671
0 58673 5 1 1 58672
0 58674 7 1 2 81762 58673
0 58675 5 1 1 58674
0 58676 7 1 2 87644 97392
0 58677 5 1 1 58676
0 58678 7 1 2 97442 97846
0 58679 7 1 2 80553 58678
0 58680 7 1 2 96471 58679
0 58681 5 1 1 58680
0 58682 7 1 2 58677 58681
0 58683 5 1 1 58682
0 58684 7 1 2 76301 58683
0 58685 5 1 1 58684
0 58686 7 1 2 92347 97932
0 58687 7 1 2 98768 58686
0 58688 5 1 1 58687
0 58689 7 1 2 88131 98250
0 58690 7 1 2 97884 58689
0 58691 5 1 1 58690
0 58692 7 1 2 58688 58691
0 58693 5 1 1 58692
0 58694 7 1 2 80053 58693
0 58695 5 1 1 58694
0 58696 7 1 2 60424 98334
0 58697 5 1 1 58696
0 58698 7 1 2 58697 98770
0 58699 5 1 1 58698
0 58700 7 1 2 80545 79296
0 58701 7 1 2 58699 58700
0 58702 5 1 1 58701
0 58703 7 1 2 63882 58702
0 58704 7 1 2 58695 58703
0 58705 7 1 2 58685 58704
0 58706 7 1 2 58675 58705
0 58707 7 1 2 58660 58706
0 58708 7 1 2 58637 58707
0 58709 7 1 2 58617 58708
0 58710 7 1 2 58575 58709
0 58711 5 1 1 58710
0 58712 7 1 2 95327 58711
0 58713 7 1 2 58540 58712
0 58714 5 1 1 58713
0 58715 7 1 2 58422 58714
0 58716 5 1 1 58715
0 58717 7 1 2 71606 58716
0 58718 5 1 1 58717
0 58719 7 1 2 97032 98118
0 58720 5 1 1 58719
0 58721 7 1 2 58720 51941
0 58722 5 1 1 58721
0 58723 7 1 2 68974 58722
0 58724 5 1 1 58723
0 58725 7 1 2 65660 76430
0 58726 7 1 2 70295 86980
0 58727 7 1 2 58725 58726
0 58728 7 1 2 98157 58727
0 58729 5 1 1 58728
0 58730 7 1 2 50372 58729
0 58731 5 1 1 58730
0 58732 7 1 2 91737 58731
0 58733 5 1 1 58732
0 58734 7 1 2 83574 98306
0 58735 5 1 1 58734
0 58736 7 1 2 58733 58735
0 58737 5 1 1 58736
0 58738 7 1 2 97769 58737
0 58739 5 1 1 58738
0 58740 7 1 2 58724 58739
0 58741 5 1 1 58740
0 58742 7 1 2 60012 58741
0 58743 5 1 1 58742
0 58744 7 1 2 73372 97622
0 58745 5 1 1 58744
0 58746 7 1 2 77045 98141
0 58747 5 1 1 58746
0 58748 7 1 2 58745 58747
0 58749 5 1 1 58748
0 58750 7 1 2 91738 58749
0 58751 5 1 1 58750
0 58752 7 1 2 97724 98272
0 58753 5 1 1 58752
0 58754 7 1 2 63618 92459
0 58755 7 1 2 97900 58754
0 58756 5 1 1 58755
0 58757 7 1 2 58753 58756
0 58758 5 1 1 58757
0 58759 7 1 2 68815 58758
0 58760 5 1 1 58759
0 58761 7 1 2 48296 58760
0 58762 5 1 1 58761
0 58763 7 1 2 59723 58762
0 58764 5 1 1 58763
0 58765 7 1 2 96247 97847
0 58766 7 1 2 83676 58765
0 58767 5 1 1 58766
0 58768 7 1 2 58764 58767
0 58769 5 1 1 58768
0 58770 7 1 2 64192 58769
0 58771 5 1 1 58770
0 58772 7 1 2 58751 58771
0 58773 5 1 1 58772
0 58774 7 1 2 97770 58773
0 58775 5 1 1 58774
0 58776 7 1 2 58743 58775
0 58777 5 1 1 58776
0 58778 7 1 2 98752 58777
0 58779 5 1 1 58778
0 58780 7 1 2 71269 86192
0 58781 7 1 2 98175 58780
0 58782 5 1 1 58781
0 58783 7 1 2 64087 97428
0 58784 7 1 2 96191 58783
0 58785 7 1 2 98326 58784
0 58786 7 1 2 98528 58785
0 58787 5 1 1 58786
0 58788 7 1 2 58782 58787
0 58789 5 1 1 58788
0 58790 7 1 2 67792 58789
0 58791 5 1 1 58790
0 58792 7 1 2 94354 94655
0 58793 7 1 2 98408 58792
0 58794 5 1 1 58793
0 58795 7 1 2 53583 58794
0 58796 5 1 1 58795
0 58797 7 1 2 90808 58796
0 58798 5 1 1 58797
0 58799 7 1 2 58791 58798
0 58800 5 1 1 58799
0 58801 7 1 2 97016 58800
0 58802 5 1 1 58801
0 58803 7 1 2 92358 93239
0 58804 7 1 2 98460 58803
0 58805 7 1 2 61959 83198
0 58806 7 1 2 98258 58805
0 58807 7 1 2 58804 58806
0 58808 7 1 2 98456 58807
0 58809 5 1 1 58808
0 58810 7 1 2 58802 58809
0 58811 5 1 1 58810
0 58812 7 1 2 76419 58811
0 58813 5 1 1 58812
0 58814 7 2 2 85542 88111
0 58815 5 2 1 98771
0 58816 7 1 2 90615 98772
0 58817 5 1 1 58816
0 58818 7 1 2 60746 86479
0 58819 5 1 1 58818
0 58820 7 1 2 58817 58819
0 58821 5 1 1 58820
0 58822 7 1 2 60425 58821
0 58823 5 1 1 58822
0 58824 7 1 2 92081 21469
0 58825 5 1 1 58824
0 58826 7 1 2 60747 58825
0 58827 5 1 1 58826
0 58828 7 1 2 58823 58827
0 58829 5 1 1 58828
0 58830 7 1 2 66787 58829
0 58831 5 1 1 58830
0 58832 7 1 2 15487 98773
0 58833 5 1 1 58832
0 58834 7 1 2 60426 58833
0 58835 5 1 1 58834
0 58836 7 1 2 92082 43233
0 58837 5 2 1 58836
0 58838 7 1 2 60643 98775
0 58839 5 1 1 58838
0 58840 7 1 2 58835 58839
0 58841 5 1 1 58840
0 58842 7 1 2 87632 58841
0 58843 5 1 1 58842
0 58844 7 1 2 58831 58843
0 58845 5 1 1 58844
0 58846 7 1 2 61960 58845
0 58847 5 1 1 58846
0 58848 7 1 2 96822 98774
0 58849 5 1 1 58848
0 58850 7 1 2 60427 58849
0 58851 5 1 1 58850
0 58852 7 1 2 61834 98776
0 58853 5 1 1 58852
0 58854 7 1 2 58851 58853
0 58855 5 1 1 58854
0 58856 7 1 2 60644 58855
0 58857 5 1 1 58856
0 58858 7 1 2 81311 92394
0 58859 5 1 1 58858
0 58860 7 1 2 58857 58859
0 58861 5 1 1 58860
0 58862 7 1 2 87131 58861
0 58863 5 1 1 58862
0 58864 7 1 2 58847 58863
0 58865 5 1 1 58864
0 58866 7 1 2 98248 58865
0 58867 5 1 1 58866
0 58868 7 1 2 67399 97697
0 58869 7 1 2 97703 58868
0 58870 5 1 1 58869
0 58871 7 1 2 58867 58870
0 58872 5 1 1 58871
0 58873 7 1 2 23565 97987
0 58874 5 1 1 58873
0 58875 7 1 2 67793 58874
0 58876 7 1 2 58872 58875
0 58877 5 1 1 58876
0 58878 7 1 2 92664 98264
0 58879 7 1 2 98163 58878
0 58880 5 1 1 58879
0 58881 7 1 2 58877 58880
0 58882 7 1 2 58813 58881
0 58883 7 1 2 58779 58882
0 58884 7 1 2 58718 58883
0 58885 7 1 2 58416 58884
0 58886 7 1 2 57864 58885
0 58887 5 1 1 58886
0 58888 7 1 2 70219 58887
0 58889 5 1 1 58888
0 58890 7 1 2 56459 58889
0 58891 7 1 2 54093 58890
0 58892 7 1 2 47636 58891
0 58893 7 1 2 44090 58892
0 58894 5 1 1 58893
0 58895 7 1 2 64195 58894
0 58896 5 1 1 58895
0 58897 7 1 2 88139 94201
0 58898 5 1 1 58897
0 58899 7 1 2 79753 79025
0 58900 7 1 2 97081 58899
0 58901 5 1 1 58900
0 58902 7 1 2 58898 58901
0 58903 5 1 1 58902
0 58904 7 1 2 95338 58903
0 58905 5 1 1 58904
0 58906 7 1 2 94084 95127
0 58907 5 1 1 58906
0 58908 7 1 2 60428 66954
0 58909 7 1 2 92676 58908
0 58910 7 1 2 93865 58909
0 58911 5 1 1 58910
0 58912 7 1 2 58907 58911
0 58913 5 1 1 58912
0 58914 7 1 2 61621 58913
0 58915 5 1 1 58914
0 58916 7 1 2 66955 80570
0 58917 7 1 2 92852 58916
0 58918 5 1 1 58917
0 58919 7 1 2 58915 58918
0 58920 5 1 1 58919
0 58921 7 1 2 65671 58920
0 58922 5 1 1 58921
0 58923 7 1 2 87598 95241
0 58924 7 1 2 94085 58923
0 58925 5 1 1 58924
0 58926 7 1 2 58922 58925
0 58927 5 1 1 58926
0 58928 7 1 2 86822 58927
0 58929 5 1 1 58928
0 58930 7 1 2 58905 58929
0 58931 5 1 1 58930
0 58932 7 1 2 81545 58931
0 58933 5 1 1 58932
0 58934 7 1 2 85554 88160
0 58935 7 1 2 93866 58934
0 58936 7 1 2 95339 58935
0 58937 5 1 1 58936
0 58938 7 1 2 58933 58937
0 58939 5 1 1 58938
0 58940 7 1 2 64193 58939
0 58941 5 1 1 58940
0 58942 7 1 2 83199 82816
0 58943 5 1 1 58942
0 58944 7 1 2 3455 58943
0 58945 5 1 1 58944
0 58946 7 1 2 71295 58945
0 58947 5 1 1 58946
0 58948 7 1 2 76302 73220
0 58949 7 1 2 80155 58948
0 58950 5 1 1 58949
0 58951 7 1 2 58947 58950
0 58952 5 1 1 58951
0 58953 7 1 2 66089 95156
0 58954 7 1 2 58952 58953
0 58955 5 1 1 58954
0 58956 7 1 2 79862 84621
0 58957 7 1 2 71296 58956
0 58958 7 1 2 86441 58957
0 58959 5 1 1 58958
0 58960 7 1 2 58955 58959
0 58961 5 1 1 58960
0 58962 7 1 2 63248 58961
0 58963 5 1 1 58962
0 58964 7 1 2 77937 84674
0 58965 7 1 2 72609 58964
0 58966 7 1 2 76303 58965
0 58967 7 1 2 86525 58966
0 58968 5 1 1 58967
0 58969 7 1 2 58963 58968
0 58970 5 1 1 58969
0 58971 7 1 2 79754 58970
0 58972 5 1 1 58971
0 58973 7 1 2 79335 80786
0 58974 5 1 1 58973
0 58975 7 1 2 75447 95196
0 58976 5 1 1 58975
0 58977 7 1 2 58974 58976
0 58978 5 2 1 58977
0 58979 7 1 2 61374 98777
0 58980 5 1 1 58979
0 58981 7 1 2 75537 80626
0 58982 5 1 1 58981
0 58983 7 1 2 58980 58982
0 58984 5 1 1 58983
0 58985 7 1 2 88095 58984
0 58986 5 1 1 58985
0 58987 7 1 2 58972 58986
0 58988 5 1 1 58987
0 58989 7 1 2 65536 58988
0 58990 5 1 1 58989
0 58991 7 1 2 66788 98778
0 58992 5 1 1 58991
0 58993 7 1 2 66605 86588
0 58994 7 1 2 81803 58993
0 58995 5 1 1 58994
0 58996 7 1 2 58992 58995
0 58997 5 1 1 58996
0 58998 7 1 2 61375 58997
0 58999 5 1 1 58998
0 59000 7 1 2 80194 80627
0 59001 5 1 1 59000
0 59002 7 1 2 58999 59001
0 59003 5 1 1 59002
0 59004 7 1 2 93691 59003
0 59005 5 1 1 59004
0 59006 7 1 2 58990 59005
0 59007 5 1 1 59006
0 59008 7 1 2 66940 59007
0 59009 5 1 1 59008
0 59010 7 1 2 67158 85936
0 59011 5 1 1 59010
0 59012 7 1 2 1988 59011
0 59013 5 1 1 59012
0 59014 7 2 2 73491 59013
0 59015 7 1 2 86067 98779
0 59016 5 1 1 59015
0 59017 7 1 2 59009 59016
0 59018 5 1 1 59017
0 59019 7 1 2 65661 59018
0 59020 5 1 1 59019
0 59021 7 1 2 95082 98780
0 59022 5 1 1 59021
0 59023 7 1 2 59020 59022
0 59024 5 1 1 59023
0 59025 7 1 2 62796 59024
0 59026 5 1 1 59025
0 59027 7 1 2 74354 84937
0 59028 5 2 1 59027
0 59029 7 1 2 74416 78683
0 59030 5 1 1 59029
0 59031 7 1 2 76304 77055
0 59032 5 1 1 59031
0 59033 7 1 2 67159 59032
0 59034 5 1 1 59033
0 59035 7 1 2 78439 26541
0 59036 7 1 2 59034 59035
0 59037 5 1 1 59036
0 59038 7 1 2 59030 59037
0 59039 5 2 1 59038
0 59040 7 1 2 98781 98783
0 59041 5 1 1 59040
0 59042 7 2 2 61148 82422
0 59043 7 1 2 80011 98785
0 59044 5 1 1 59043
0 59045 7 1 2 74850 94555
0 59046 5 1 1 59045
0 59047 7 1 2 68186 90592
0 59048 5 1 1 59047
0 59049 7 1 2 59046 59048
0 59050 5 1 1 59049
0 59051 7 1 2 64372 59050
0 59052 5 1 1 59051
0 59053 7 1 2 65750 76431
0 59054 7 1 2 98786 59053
0 59055 5 1 1 59054
0 59056 7 1 2 78947 59055
0 59057 7 1 2 59052 59056
0 59058 5 1 1 59057
0 59059 7 1 2 62166 59058
0 59060 5 1 1 59059
0 59061 7 1 2 59044 59060
0 59062 5 1 1 59061
0 59063 7 1 2 95157 59062
0 59064 5 1 1 59063
0 59065 7 1 2 59041 59064
0 59066 5 1 1 59065
0 59067 7 1 2 63619 59066
0 59068 5 1 1 59067
0 59069 7 1 2 71297 88629
0 59070 5 1 1 59069
0 59071 7 1 2 72405 59070
0 59072 5 1 1 59071
0 59073 7 1 2 65041 59072
0 59074 7 1 2 44430 59073
0 59075 5 1 1 59074
0 59076 7 1 2 95154 59075
0 59077 5 1 1 59076
0 59078 7 1 2 70220 97064
0 59079 5 1 1 59078
0 59080 7 1 2 63249 59079
0 59081 7 1 2 59077 59080
0 59082 5 1 1 59081
0 59083 7 1 2 64373 95168
0 59084 5 1 1 59083
0 59085 7 1 2 76903 77837
0 59086 7 1 2 87692 59085
0 59087 7 1 2 59084 59086
0 59088 5 1 1 59087
0 59089 7 1 2 59082 59088
0 59090 5 1 1 59089
0 59091 7 1 2 75856 59090
0 59092 5 1 1 59091
0 59093 7 1 2 59068 59092
0 59094 5 1 1 59093
0 59095 7 1 2 65311 59094
0 59096 5 1 1 59095
0 59097 7 1 2 70097 98784
0 59098 5 1 1 59097
0 59099 7 3 2 63250 95158
0 59100 7 1 2 78641 78535
0 59101 7 1 2 98787 59100
0 59102 5 1 1 59101
0 59103 7 1 2 59098 59102
0 59104 5 1 1 59103
0 59105 7 1 2 90728 59104
0 59106 5 1 1 59105
0 59107 7 1 2 59096 59106
0 59108 5 1 1 59107
0 59109 7 1 2 67794 94479
0 59110 7 1 2 59108 59109
0 59111 5 1 1 59110
0 59112 7 1 2 68816 59111
0 59113 7 1 2 59026 59112
0 59114 5 1 1 59113
0 59115 7 1 2 74372 87323
0 59116 5 1 1 59115
0 59117 7 1 2 68187 95159
0 59118 7 1 2 76936 59117
0 59119 5 1 1 59118
0 59120 7 1 2 63251 92483
0 59121 5 1 1 59120
0 59122 7 1 2 59119 59121
0 59123 5 2 1 59122
0 59124 7 1 2 66606 98790
0 59125 5 1 1 59124
0 59126 7 1 2 82866 84934
0 59127 5 1 1 59126
0 59128 7 1 2 59125 59127
0 59129 5 1 1 59128
0 59130 7 1 2 98437 59129
0 59131 5 1 1 59130
0 59132 7 1 2 59116 59131
0 59133 5 1 1 59132
0 59134 7 1 2 65662 59133
0 59135 5 1 1 59134
0 59136 7 1 2 87144 89533
0 59137 5 1 1 59136
0 59138 7 1 2 59135 59137
0 59139 5 1 1 59138
0 59140 7 1 2 60429 59139
0 59141 5 1 1 59140
0 59142 7 1 2 74951 94899
0 59143 7 1 2 98791 59142
0 59144 5 1 1 59143
0 59145 7 1 2 59141 59144
0 59146 5 1 1 59145
0 59147 7 1 2 67795 59146
0 59148 5 1 1 59147
0 59149 7 1 2 83066 98782
0 59150 5 1 1 59149
0 59151 7 1 2 79897 98788
0 59152 5 1 1 59151
0 59153 7 1 2 59150 59152
0 59154 5 1 1 59153
0 59155 7 1 2 60430 59154
0 59156 5 1 1 59155
0 59157 7 1 2 74978 97138
0 59158 5 1 1 59157
0 59159 7 1 2 59156 59158
0 59160 5 1 1 59159
0 59161 7 1 2 73801 88076
0 59162 7 1 2 59160 59161
0 59163 5 1 1 59162
0 59164 7 1 2 59148 59163
0 59165 5 1 1 59164
0 59166 7 1 2 79641 59165
0 59167 5 1 1 59166
0 59168 7 1 2 87320 87594
0 59169 7 1 2 88213 59168
0 59170 7 1 2 94935 59169
0 59171 5 1 1 59170
0 59172 7 1 2 59167 59171
0 59173 5 1 1 59172
0 59174 7 1 2 68580 59173
0 59175 5 1 1 59174
0 59176 7 1 2 71014 75884
0 59177 5 1 1 59176
0 59178 7 1 2 75451 95482
0 59179 7 1 2 89114 59178
0 59180 5 1 1 59179
0 59181 7 1 2 59177 59180
0 59182 5 1 1 59181
0 59183 7 1 2 98789 59182
0 59184 5 1 1 59183
0 59185 7 1 2 83200 82432
0 59186 7 1 2 86450 59185
0 59187 5 1 1 59186
0 59188 7 1 2 59184 59187
0 59189 5 1 1 59188
0 59190 7 1 2 62797 59189
0 59191 5 1 1 59190
0 59192 7 1 2 67796 86442
0 59193 7 1 2 97667 59192
0 59194 5 1 1 59193
0 59195 7 1 2 59191 59194
0 59196 5 1 1 59195
0 59197 7 1 2 86193 59196
0 59198 5 1 1 59197
0 59199 7 1 2 87254 94265
0 59200 5 1 1 59199
0 59201 7 1 2 59198 59200
0 59202 5 1 1 59201
0 59203 7 1 2 65663 59202
0 59204 5 1 1 59203
0 59205 7 1 2 66941 96284
0 59206 7 1 2 87531 59205
0 59207 7 1 2 93861 59206
0 59208 5 1 1 59207
0 59209 7 1 2 59204 59208
0 59210 5 1 1 59209
0 59211 7 1 2 81194 59210
0 59212 5 1 1 59211
0 59213 7 1 2 63883 59212
0 59214 7 1 2 59175 59213
0 59215 5 1 1 59214
0 59216 7 1 2 95232 59215
0 59217 7 1 2 59114 59216
0 59218 5 1 1 59217
0 59219 7 1 2 58941 59218
0 59220 5 1 1 59219
0 59221 7 1 2 69040 59220
0 59222 5 1 1 59221
0 59223 7 1 2 64196 77803
0 59224 7 1 2 85804 86457
0 59225 7 1 2 59223 59224
0 59226 7 1 2 97771 98145
0 59227 7 1 2 59225 59226
0 59228 5 1 1 59227
0 59229 7 1 2 59222 59228
0 59230 5 1 1 59229
0 59231 7 1 2 69142 69285
0 59232 7 1 2 59230 59231
0 59233 5 1 1 59232
0 59234 7 1 2 58896 59233
0 59235 7 1 2 35909 59234
3 129999 5 0 1 59235
