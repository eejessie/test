1 0 0 2 0
2 49 1 0
2 1482 1 0
1 1 0 2 0
2 1483 1 1
2 1484 1 1
1 2 0 2 0
2 1485 1 2
2 1486 1 2
1 3 0 2 0
2 1487 1 3
2 1488 1 3
1 4 0 2 0
2 1489 1 4
2 1490 1 4
1 5 0 2 0
2 1491 1 5
2 1492 1 5
1 6 0 2 0
2 1493 1 6
2 1494 1 6
1 7 0 2 0
2 1495 1 7
2 1496 1 7
1 8 0 2 0
2 1497 1 8
2 1498 1 8
1 9 0 2 0
2 1499 1 9
2 1500 1 9
1 10 0 2 0
2 1501 1 10
2 1502 1 10
1 11 0 2 0
2 1503 1 11
2 1504 1 11
1 12 0 2 0
2 1505 1 12
2 1506 1 12
1 13 0 2 0
2 1507 1 13
2 1508 1 13
1 14 0 2 0
2 1509 1 14
2 1510 1 14
1 15 0 2 0
2 1511 1 15
2 1512 1 15
1 16 0 2 0
2 1513 1 16
2 1514 1 16
1 17 0 2 0
2 1515 1 17
2 1516 1 17
1 18 0 2 0
2 1517 1 18
2 1518 1 18
1 19 0 2 0
2 1519 1 19
2 1520 1 19
1 20 0 2 0
2 1521 1 20
2 1522 1 20
1 21 0 2 0
2 1523 1 21
2 1524 1 21
1 22 0 2 0
2 1525 1 22
2 1526 1 22
1 23 0 2 0
2 1527 1 23
2 1528 1 23
1 24 0 2 0
2 1529 1 24
2 1530 1 24
1 25 0 2 0
2 1531 1 25
2 1532 1 25
1 26 0 2 0
2 1533 1 26
2 1534 1 26
1 27 0 2 0
2 1535 1 27
2 1536 1 27
1 28 0 2 0
2 1537 1 28
2 1538 1 28
1 29 0 2 0
2 1539 1 29
2 1540 1 29
1 30 0 2 0
2 1541 1 30
2 1542 1 30
1 31 0 2 0
2 1543 1 31
2 1544 1 31
1 32 0 3 0
2 1545 1 32
2 1546 1 32
2 1547 1 32
1 33 0 2 0
2 1548 1 33
2 1549 1 33
1 34 0 2 0
2 1550 1 34
2 1551 1 34
1 35 0 2 0
2 1552 1 35
2 1553 1 35
1 36 0 2 0
2 1554 1 36
2 1555 1 36
1 37 0 2 0
2 1556 1 37
2 1557 1 37
1 38 0 2 0
2 1558 1 38
2 1559 1 38
1 39 0 2 0
2 1560 1 39
2 1561 1 39
1 40 0 2 0
2 1562 1 40
2 1563 1 40
1 41 0 2 0
2 1564 1 41
2 1565 1 41
1 42 0 2 0
2 1566 1 42
2 1567 1 42
1 43 0 2 0
2 1568 1 43
2 1569 1 43
1 44 0 2 0
2 1570 1 44
2 1571 1 44
1 45 0 2 0
2 1572 1 45
2 1573 1 45
1 46 0 2 0
2 1574 1 46
2 1575 1 46
1 47 0 2 0
2 1576 1 47
2 1577 1 47
1 48 0 2 0
2 1578 1 48
2 1579 1 48
2 1580 1 69
2 1581 1 69
2 1582 1 70
2 1583 1 70
2 1584 1 71
2 1585 1 71
2 1586 1 72
2 1587 1 72
2 1588 1 73
2 1589 1 73
2 1590 1 74
2 1591 1 74
2 1592 1 75
2 1593 1 75
2 1594 1 76
2 1595 1 76
2 1596 1 77
2 1597 1 77
2 1598 1 78
2 1599 1 78
2 1600 1 79
2 1601 1 79
2 1602 1 80
2 1603 1 80
2 1604 1 81
2 1605 1 81
2 1606 1 98
2 1607 1 98
2 1608 1 100
2 1609 1 100
2 1610 1 102
2 1611 1 102
2 1612 1 104
2 1613 1 104
2 1614 1 106
2 1615 1 106
2 1616 1 107
2 1617 1 107
2 1618 1 108
2 1619 1 108
2 1620 1 108
2 1621 1 111
2 1622 1 111
2 1623 1 112
2 1624 1 112
2 1625 1 115
2 1626 1 115
2 1627 1 118
2 1628 1 118
2 1629 1 120
2 1630 1 120
2 1631 1 123
2 1632 1 123
2 1633 1 126
2 1634 1 126
2 1635 1 128
2 1636 1 128
2 1637 1 131
2 1638 1 131
2 1639 1 134
2 1640 1 134
2 1641 1 136
2 1642 1 136
2 1643 1 139
2 1644 1 139
2 1645 1 142
2 1646 1 142
2 1647 1 144
2 1648 1 144
2 1649 1 147
2 1650 1 147
2 1651 1 150
2 1652 1 150
2 1653 1 152
2 1654 1 152
2 1655 1 155
2 1656 1 155
2 1657 1 158
2 1658 1 158
2 1659 1 160
2 1660 1 160
2 1661 1 163
2 1662 1 163
2 1663 1 166
2 1664 1 166
2 1665 1 168
2 1666 1 168
2 1667 1 171
2 1668 1 171
2 1669 1 174
2 1670 1 174
2 1671 1 176
2 1672 1 176
2 1673 1 179
2 1674 1 179
2 1675 1 182
2 1676 1 182
2 1677 1 184
2 1678 1 184
2 1679 1 187
2 1680 1 187
2 1681 1 190
2 1682 1 190
2 1683 1 192
2 1684 1 192
2 1685 1 195
2 1686 1 195
2 1687 1 198
2 1688 1 198
2 1689 1 200
2 1690 1 200
2 1691 1 203
2 1692 1 203
2 1693 1 206
2 1694 1 206
2 1695 1 208
2 1696 1 208
2 1697 1 211
2 1698 1 211
2 1699 1 214
2 1700 1 214
2 1701 1 216
2 1702 1 216
2 1703 1 219
2 1704 1 219
2 1705 1 219
2 1706 1 219
2 1707 1 220
2 1708 1 220
2 1709 1 221
2 1710 1 221
2 1711 1 222
2 1712 1 222
2 1713 1 222
2 1714 1 222
2 1715 1 224
2 1716 1 224
2 1717 1 224
2 1718 1 224
2 1719 1 225
2 1720 1 225
2 1721 1 231
2 1722 1 231
2 1723 1 231
2 1724 1 231
2 1725 1 232
2 1726 1 232
2 1727 1 232
2 1728 1 234
2 1729 1 234
2 1730 1 234
2 1731 1 236
2 1732 1 236
2 1733 1 236
2 1734 1 237
2 1735 1 237
2 1736 1 243
2 1737 1 243
2 1738 1 243
2 1739 1 243
2 1740 1 244
2 1741 1 244
2 1742 1 244
2 1743 1 246
2 1744 1 246
2 1745 1 246
2 1746 1 248
2 1747 1 248
2 1748 1 248
2 1749 1 249
2 1750 1 249
2 1751 1 255
2 1752 1 255
2 1753 1 255
2 1754 1 255
2 1755 1 256
2 1756 1 256
2 1757 1 256
2 1758 1 258
2 1759 1 258
2 1760 1 258
2 1761 1 260
2 1762 1 260
2 1763 1 260
2 1764 1 261
2 1765 1 261
2 1766 1 267
2 1767 1 267
2 1768 1 267
2 1769 1 267
2 1770 1 268
2 1771 1 268
2 1772 1 270
2 1773 1 270
2 1774 1 270
2 1775 1 272
2 1776 1 272
2 1777 1 272
2 1778 1 273
2 1779 1 273
2 1780 1 279
2 1781 1 279
2 1782 1 279
2 1783 1 279
2 1784 1 280
2 1785 1 280
2 1786 1 280
2 1787 1 282
2 1788 1 282
2 1789 1 282
2 1790 1 284
2 1791 1 284
2 1792 1 284
2 1793 1 285
2 1794 1 285
2 1795 1 291
2 1796 1 291
2 1797 1 291
2 1798 1 292
2 1799 1 292
2 1800 1 292
2 1801 1 294
2 1802 1 294
2 1803 1 294
2 1804 1 296
2 1805 1 296
2 1806 1 296
2 1807 1 297
2 1808 1 297
2 1809 1 303
2 1810 1 303
2 1811 1 303
2 1812 1 303
2 1813 1 304
2 1814 1 304
2 1815 1 304
2 1816 1 306
2 1817 1 306
2 1818 1 306
2 1819 1 308
2 1820 1 308
2 1821 1 308
2 1822 1 309
2 1823 1 309
2 1824 1 315
2 1825 1 315
2 1826 1 315
2 1827 1 316
2 1828 1 316
2 1829 1 316
2 1830 1 318
2 1831 1 318
2 1832 1 318
2 1833 1 320
2 1834 1 320
2 1835 1 320
2 1836 1 321
2 1837 1 321
2 1838 1 327
2 1839 1 327
2 1840 1 327
2 1841 1 327
2 1842 1 328
2 1843 1 328
2 1844 1 328
2 1845 1 330
2 1846 1 330
2 1847 1 330
2 1848 1 332
2 1849 1 332
2 1850 1 332
2 1851 1 333
2 1852 1 333
2 1853 1 339
2 1854 1 339
2 1855 1 340
2 1856 1 340
2 1857 1 340
2 1858 1 342
2 1859 1 342
2 1860 1 342
2 1861 1 344
2 1862 1 344
2 1863 1 344
2 1864 1 345
2 1865 1 345
2 1866 1 351
2 1867 1 351
2 1868 1 351
2 1869 1 351
2 1870 1 352
2 1871 1 352
2 1872 1 352
2 1873 1 354
2 1874 1 354
2 1875 1 354
2 1876 1 356
2 1877 1 356
2 1878 1 356
2 1879 1 357
2 1880 1 357
2 1881 1 363
2 1882 1 363
2 1883 1 364
2 1884 1 364
2 1885 1 364
2 1886 1 366
2 1887 1 366
2 1888 1 366
2 1889 1 368
2 1890 1 368
2 1891 1 368
2 1892 1 369
2 1893 1 369
2 1894 1 375
2 1895 1 375
2 1896 1 375
2 1897 1 375
2 1898 1 376
2 1899 1 376
2 1900 1 376
2 1901 1 378
2 1902 1 378
2 1903 1 378
2 1904 1 380
2 1905 1 380
2 1906 1 380
2 1907 1 381
2 1908 1 381
2 1909 1 387
2 1910 1 387
2 1911 1 387
2 1912 1 387
2 1913 1 390
2 1914 1 390
2 1915 1 390
2 1916 1 392
2 1917 1 392
2 1918 1 392
2 1919 1 393
2 1920 1 393
2 1921 1 399
2 1922 1 399
2 1923 1 399
2 1924 1 399
2 1925 1 400
2 1926 1 400
2 1927 1 400
2 1928 1 402
2 1929 1 402
2 1930 1 402
2 1931 1 404
2 1932 1 404
2 1933 1 404
2 1934 1 407
2 1935 1 407
2 1936 1 407
2 1937 1 408
2 1938 1 408
2 1939 1 409
2 1940 1 409
2 1941 1 410
2 1942 1 410
2 1943 1 410
2 1944 1 413
2 1945 1 413
2 1946 1 414
2 1947 1 414
2 1948 1 417
2 1949 1 417
2 1950 1 418
2 1951 1 418
2 1952 1 421
2 1953 1 421
2 1954 1 422
2 1955 1 422
2 1956 1 425
2 1957 1 425
2 1958 1 426
2 1959 1 426
2 1960 1 429
2 1961 1 429
2 1962 1 430
2 1963 1 430
2 1964 1 433
2 1965 1 433
2 1966 1 434
2 1967 1 434
2 1968 1 437
2 1969 1 437
2 1970 1 438
2 1971 1 438
2 1972 1 441
2 1973 1 441
2 1974 1 442
2 1975 1 442
2 1976 1 445
2 1977 1 445
2 1978 1 446
2 1979 1 446
2 1980 1 449
2 1981 1 449
2 1982 1 450
2 1983 1 450
2 1984 1 453
2 1985 1 453
2 1986 1 454
2 1987 1 454
2 1988 1 457
2 1989 1 457
2 1990 1 458
2 1991 1 458
2 1992 1 461
2 1993 1 461
2 1994 1 462
2 1995 1 462
2 1996 1 465
2 1997 1 465
2 1998 1 466
2 1999 1 466
2 2000 1 469
2 2001 1 469
2 2002 1 469
2 2003 1 470
2 2004 1 470
2 2005 1 470
2 2006 1 473
2 2007 1 473
2 2008 1 474
2 2009 1 474
2 2010 1 475
2 2011 1 475
2 2012 1 475
2 2013 1 476
2 2014 1 476
2 2015 1 481
2 2016 1 481
2 2017 1 481
2 2018 1 482
2 2019 1 482
2 2020 1 484
2 2021 1 484
2 2022 1 485
2 2023 1 485
2 2024 1 485
2 2025 1 486
2 2026 1 486
2 2027 1 491
2 2028 1 491
2 2029 1 491
2 2030 1 492
2 2031 1 492
2 2032 1 493
2 2033 1 493
2 2034 1 493
2 2035 1 494
2 2036 1 494
2 2037 1 499
2 2038 1 499
2 2039 1 502
2 2040 1 502
2 2041 1 503
2 2042 1 503
2 2043 1 503
2 2044 1 504
2 2045 1 504
2 2046 1 509
2 2047 1 509
2 2048 1 509
2 2049 1 510
2 2050 1 510
2 2051 1 512
2 2052 1 512
2 2053 1 513
2 2054 1 513
2 2055 1 513
2 2056 1 514
2 2057 1 514
2 2058 1 519
2 2059 1 519
2 2060 1 519
2 2061 1 520
2 2062 1 520
2 2063 1 522
2 2064 1 522
2 2065 1 523
2 2066 1 523
2 2067 1 523
2 2068 1 524
2 2069 1 524
2 2070 1 529
2 2071 1 529
2 2072 1 529
2 2073 1 530
2 2074 1 530
2 2075 1 532
2 2076 1 532
2 2077 1 533
2 2078 1 533
2 2079 1 533
2 2080 1 534
2 2081 1 534
2 2082 1 539
2 2083 1 539
2 2084 1 539
2 2085 1 540
2 2086 1 540
2 2087 1 542
2 2088 1 542
2 2089 1 543
2 2090 1 543
2 2091 1 543
2 2092 1 544
2 2093 1 544
2 2094 1 549
2 2095 1 549
2 2096 1 549
2 2097 1 550
2 2098 1 550
2 2099 1 552
2 2100 1 552
2 2101 1 553
2 2102 1 553
2 2103 1 553
2 2104 1 554
2 2105 1 554
2 2106 1 559
2 2107 1 559
2 2108 1 559
2 2109 1 560
2 2110 1 560
2 2111 1 562
2 2112 1 562
2 2113 1 563
2 2114 1 563
2 2115 1 563
2 2116 1 564
2 2117 1 564
2 2118 1 569
2 2119 1 569
2 2120 1 569
2 2121 1 570
2 2122 1 570
2 2123 1 572
2 2124 1 572
2 2125 1 573
2 2126 1 573
2 2127 1 573
2 2128 1 574
2 2129 1 574
2 2130 1 579
2 2131 1 579
2 2132 1 579
2 2133 1 580
2 2134 1 580
2 2135 1 582
2 2136 1 582
2 2137 1 583
2 2138 1 583
2 2139 1 583
2 2140 1 584
2 2141 1 584
2 2142 1 589
2 2143 1 589
2 2144 1 589
2 2145 1 590
2 2146 1 590
2 2147 1 592
2 2148 1 592
2 2149 1 593
2 2150 1 593
2 2151 1 593
2 2152 1 594
2 2153 1 594
2 2154 1 599
2 2155 1 599
2 2156 1 599
2 2157 1 600
2 2158 1 600
2 2159 1 602
2 2160 1 602
2 2161 1 603
2 2162 1 603
2 2163 1 603
2 2164 1 604
2 2165 1 604
2 2166 1 609
2 2167 1 609
2 2168 1 609
2 2169 1 610
2 2170 1 610
2 2171 1 612
2 2172 1 612
2 2173 1 613
2 2174 1 613
2 2175 1 613
2 2176 1 614
2 2177 1 614
2 2178 1 619
2 2179 1 619
2 2180 1 619
2 2181 1 620
2 2182 1 620
2 2183 1 622
2 2184 1 622
2 2185 1 623
2 2186 1 623
2 2187 1 623
2 2188 1 624
2 2189 1 624
2 2190 1 629
2 2191 1 629
2 2192 1 632
2 2193 1 632
2 2194 1 633
2 2195 1 633
2 2196 1 634
2 2197 1 634
2 2198 1 634
2 2199 1 635
2 2200 1 635
2 2201 1 635
2 2202 1 636
2 2203 1 636
2 2204 1 637
2 2205 1 637
2 2206 1 638
2 2207 1 638
2 2208 1 641
2 2209 1 641
2 2210 1 644
2 2211 1 644
2 2212 1 645
2 2213 1 645
2 2214 1 649
2 2215 1 649
2 2216 1 652
2 2217 1 652
2 2218 1 653
2 2219 1 653
2 2220 1 657
2 2221 1 657
2 2222 1 660
2 2223 1 660
2 2224 1 661
2 2225 1 661
2 2226 1 665
2 2227 1 665
2 2228 1 668
2 2229 1 668
2 2230 1 669
2 2231 1 669
2 2232 1 673
2 2233 1 673
2 2234 1 676
2 2235 1 676
2 2236 1 677
2 2237 1 677
2 2238 1 681
2 2239 1 681
2 2240 1 684
2 2241 1 684
2 2242 1 685
2 2243 1 685
2 2244 1 689
2 2245 1 689
2 2246 1 692
2 2247 1 692
2 2248 1 693
2 2249 1 693
2 2250 1 697
2 2251 1 697
2 2252 1 700
2 2253 1 700
2 2254 1 701
2 2255 1 701
2 2256 1 705
2 2257 1 705
2 2258 1 708
2 2259 1 708
2 2260 1 709
2 2261 1 709
2 2262 1 713
2 2263 1 713
2 2264 1 716
2 2265 1 716
2 2266 1 717
2 2267 1 717
2 2268 1 721
2 2269 1 721
2 2270 1 724
2 2271 1 724
2 2272 1 725
2 2273 1 725
2 2274 1 729
2 2275 1 729
2 2276 1 732
2 2277 1 732
2 2278 1 733
2 2279 1 733
2 2280 1 737
2 2281 1 737
2 2282 1 740
2 2283 1 740
2 2284 1 741
2 2285 1 741
2 2286 1 745
2 2287 1 745
2 2288 1 748
2 2289 1 748
2 2290 1 749
2 2291 1 749
2 2292 1 753
2 2293 1 753
2 2294 1 756
2 2295 1 756
2 2296 1 757
2 2297 1 757
2 2298 1 763
2 2299 1 763
2 2300 1 766
2 2301 1 766
2 2302 1 768
2 2303 1 768
2 2304 1 775
2 2305 1 775
2 2306 1 781
2 2307 1 781
2 2308 1 793
2 2309 1 793
2 2310 1 801
2 2311 1 801
2 2312 1 809
2 2313 1 809
2 2314 1 815
2 2315 1 815
2 2316 1 823
2 2317 1 823
2 2318 1 827
2 2319 1 827
2 2320 1 835
2 2321 1 835
2 2322 1 839
2 2323 1 839
2 2324 1 847
2 2325 1 847
2 2326 1 849
2 2327 1 849
2 2328 1 850
2 2329 1 850
2 2330 1 851
2 2331 1 851
2 2332 1 856
2 2333 1 856
2 2334 1 867
2 2335 1 867
2 2336 1 875
2 2337 1 875
2 2338 1 887
2 2339 1 887
2 2340 1 899
2 2341 1 899
2 2342 1 920
2 2343 1 920
2 2344 1 931
2 2345 1 931
2 2346 1 939
2 2347 1 939
2 2348 1 947
2 2349 1 947
2 2350 1 976
2 2351 1 976
2 2352 1 977
2 2353 1 977
2 2354 1 980
2 2355 1 980
2 2356 1 980
2 2357 1 984
2 2358 1 984
2 2359 1 985
2 2360 1 985
2 2361 1 988
2 2362 1 988
2 2363 1 989
2 2364 1 989
2 2365 1 992
2 2366 1 992
2 2367 1 993
2 2368 1 993
2 2369 1 996
2 2370 1 996
2 2371 1 997
2 2372 1 997
2 2373 1 1000
2 2374 1 1000
2 2375 1 1001
2 2376 1 1001
2 2377 1 1004
2 2378 1 1004
2 2379 1 1005
2 2380 1 1005
2 2381 1 1008
2 2382 1 1008
2 2383 1 1009
2 2384 1 1009
2 2385 1 1012
2 2386 1 1012
2 2387 1 1013
2 2388 1 1013
2 2389 1 1016
2 2390 1 1016
2 2391 1 1017
2 2392 1 1017
2 2393 1 1020
2 2394 1 1020
2 2395 1 1021
2 2396 1 1021
2 2397 1 1024
2 2398 1 1024
2 2399 1 1025
2 2400 1 1025
2 2401 1 1028
2 2402 1 1028
2 2403 1 1029
2 2404 1 1029
2 2405 1 1032
2 2406 1 1032
2 2407 1 1032
2 2408 1 1033
2 2409 1 1033
2 2410 1 1033
2 2411 1 1036
2 2412 1 1036
2 2413 1 1036
2 2414 1 1037
2 2415 1 1037
2 2416 1 1044
2 2417 1 1044
2 2418 1 1044
2 2419 1 1045
2 2420 1 1045
2 2421 1 1050
2 2422 1 1050
2 2423 1 1053
2 2424 1 1053
2 2425 1 1058
2 2426 1 1058
2 2427 1 1058
2 2428 1 1059
2 2429 1 1059
2 2430 1 1064
2 2431 1 1064
2 2432 1 1064
2 2433 1 1065
2 2434 1 1065
2 2435 1 1067
2 2436 1 1067
2 2437 1 1072
2 2438 1 1072
2 2439 1 1072
2 2440 1 1073
2 2441 1 1073
2 2442 1 1075
2 2443 1 1075
2 2444 1 1080
2 2445 1 1080
2 2446 1 1080
2 2447 1 1081
2 2448 1 1081
2 2449 1 1083
2 2450 1 1083
2 2451 1 1088
2 2452 1 1088
2 2453 1 1088
2 2454 1 1089
2 2455 1 1089
2 2456 1 1091
2 2457 1 1091
2 2458 1 1096
2 2459 1 1096
2 2460 1 1096
2 2461 1 1097
2 2462 1 1097
2 2463 1 1099
2 2464 1 1099
2 2465 1 1104
2 2466 1 1104
2 2467 1 1104
2 2468 1 1105
2 2469 1 1105
2 2470 1 1107
2 2471 1 1107
2 2472 1 1112
2 2473 1 1112
2 2474 1 1112
2 2475 1 1113
2 2476 1 1113
2 2477 1 1115
2 2478 1 1115
2 2479 1 1120
2 2480 1 1120
2 2481 1 1120
2 2482 1 1121
2 2483 1 1121
2 2484 1 1123
2 2485 1 1123
2 2486 1 1128
2 2487 1 1128
2 2488 1 1128
2 2489 1 1129
2 2490 1 1129
2 2491 1 1131
2 2492 1 1131
2 2493 1 1136
2 2494 1 1136
2 2495 1 1136
2 2496 1 1137
2 2497 1 1137
2 2498 1 1139
2 2499 1 1139
2 2500 1 1144
2 2501 1 1144
2 2502 1 1144
2 2503 1 1145
2 2504 1 1145
2 2505 1 1147
2 2506 1 1147
2 2507 1 1152
2 2508 1 1152
2 2509 1 1152
2 2510 1 1152
2 2511 1 1155
2 2512 1 1155
2 2513 1 1158
2 2514 1 1158
2 2515 1 1161
2 2516 1 1161
2 2517 1 1162
2 2518 1 1162
2 2519 1 1163
2 2520 1 1163
2 2521 1 1166
2 2522 1 1166
2 2523 1 1169
2 2524 1 1169
2 2525 1 1170
2 2526 1 1170
2 2527 1 1174
2 2528 1 1174
2 2529 1 1177
2 2530 1 1177
2 2531 1 1178
2 2532 1 1178
2 2533 1 1182
2 2534 1 1182
2 2535 1 1185
2 2536 1 1185
2 2537 1 1186
2 2538 1 1186
2 2539 1 1190
2 2540 1 1190
2 2541 1 1193
2 2542 1 1193
2 2543 1 1194
2 2544 1 1194
2 2545 1 1198
2 2546 1 1198
2 2547 1 1201
2 2548 1 1201
2 2549 1 1202
2 2550 1 1202
2 2551 1 1206
2 2552 1 1206
2 2553 1 1209
2 2554 1 1209
2 2555 1 1210
2 2556 1 1210
2 2557 1 1214
2 2558 1 1214
2 2559 1 1217
2 2560 1 1217
2 2561 1 1218
2 2562 1 1218
2 2563 1 1222
2 2564 1 1222
2 2565 1 1225
2 2566 1 1225
2 2567 1 1226
2 2568 1 1226
2 2569 1 1230
2 2570 1 1230
2 2571 1 1233
2 2572 1 1233
2 2573 1 1234
2 2574 1 1234
2 2575 1 1238
2 2576 1 1238
2 2577 1 1241
2 2578 1 1241
2 2579 1 1242
2 2580 1 1242
2 2581 1 1246
2 2582 1 1246
2 2583 1 1249
2 2584 1 1249
2 2585 1 1250
2 2586 1 1250
2 2587 1 1254
2 2588 1 1254
2 2589 1 1257
2 2590 1 1257
2 2591 1 1258
2 2592 1 1258
2 2593 1 1262
2 2594 1 1262
2 2595 1 1265
2 2596 1 1265
2 2597 1 1266
2 2598 1 1266
2 2599 1 1270
2 2600 1 1270
2 2601 1 1273
2 2602 1 1273
2 2603 1 1274
2 2604 1 1274
2 2605 1 1280
2 2606 1 1280
2 2607 1 1286
2 2608 1 1286
2 2609 1 1288
2 2610 1 1288
2 2611 1 1291
2 2612 1 1291
2 2613 1 1300
2 2614 1 1300
2 2615 1 1306
2 2616 1 1306
2 2617 1 1314
2 2618 1 1314
2 2619 1 1322
2 2620 1 1322
2 2621 1 1326
2 2622 1 1326
2 2623 1 1334
2 2624 1 1334
2 2625 1 1338
2 2626 1 1338
2 2627 1 1346
2 2628 1 1346
2 2629 1 1350
2 2630 1 1350
2 2631 1 1358
2 2632 1 1358
2 2633 1 1362
2 2634 1 1362
2 2635 1 1370
2 2636 1 1370
2 2637 1 1374
2 2638 1 1374
2 2639 1 1389
2 2640 1 1389
2 2641 1 1401
2 2642 1 1401
2 2643 1 1413
2 2644 1 1413
2 2645 1 1425
2 2646 1 1425
2 2647 1 1437
2 2648 1 1437
2 2649 1 1452
2 2650 1 1452
0 50 5 1 1 49
0 51 5 1 1 1483
0 52 5 1 1 1485
0 53 5 1 1 1487
0 54 5 1 1 1489
0 55 5 1 1 1491
0 56 5 1 1 1493
0 57 5 1 1 1495
0 58 5 1 1 1497
0 59 5 1 1 1499
0 60 5 1 1 1501
0 61 5 1 1 1503
0 62 5 1 1 1505
0 63 5 1 1 1507
0 64 5 1 1 1509
0 65 5 1 1 1511
0 66 5 1 1 1513
0 67 5 1 1 1515
0 68 5 1 1 1517
0 69 5 2 1 1519
0 70 5 2 1 1521
0 71 5 2 1 1523
0 72 5 2 1 1525
0 73 5 2 1 1527
0 74 5 2 1 1529
0 75 5 2 1 1531
0 76 5 2 1 1533
0 77 5 2 1 1535
0 78 5 2 1 1537
0 79 5 2 1 1539
0 80 5 2 1 1541
0 81 5 2 1 1543
0 82 5 1 1 1545
0 83 5 1 1 1548
0 84 5 1 1 1550
0 85 5 1 1 1552
0 86 5 1 1 1554
0 87 5 1 1 1556
0 88 5 1 1 1558
0 89 5 1 1 1560
0 90 5 1 1 1562
0 91 5 1 1 1564
0 92 5 1 1 1566
0 93 5 1 1 1568
0 94 5 1 1 1570
0 95 5 1 1 1572
0 96 5 1 1 1574
0 97 5 1 1 1576
0 98 5 2 1 1578
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 1486 1518
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 1484 1516
0 106 5 2 1 105
0 107 7 2 2 1482 1514
0 108 5 3 1 1616
0 109 7 1 2 1614 1618
0 110 5 1 1 109
0 111 7 2 2 1612 110
0 112 5 2 1 1621
0 113 7 1 2 1610 1623
0 114 5 1 1 113
0 115 7 2 2 1608 114
0 116 5 1 1 1625
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 1488 1626
0 120 5 2 1 119
0 121 7 1 2 1580 1629
0 122 5 1 1 121
0 123 7 2 2 1627 122
0 124 5 1 1 1631
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 1490 1632
0 128 5 2 1 127
0 129 7 1 2 1582 1635
0 130 5 1 1 129
0 131 7 2 2 1633 130
0 132 5 1 1 1637
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 1492 1638
0 136 5 2 1 135
0 137 7 1 2 1584 1641
0 138 5 1 1 137
0 139 7 2 2 1639 138
0 140 5 1 1 1643
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 1494 1644
0 144 5 2 1 143
0 145 7 1 2 1586 1647
0 146 5 1 1 145
0 147 7 2 2 1645 146
0 148 5 1 1 1649
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 1496 1650
0 152 5 2 1 151
0 153 7 1 2 1588 1653
0 154 5 1 1 153
0 155 7 2 2 1651 154
0 156 5 1 1 1655
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 1498 1656
0 160 5 2 1 159
0 161 7 1 2 1590 1659
0 162 5 1 1 161
0 163 7 2 2 1657 162
0 164 5 1 1 1661
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 1500 1662
0 168 5 2 1 167
0 169 7 1 2 1592 1665
0 170 5 1 1 169
0 171 7 2 2 1663 170
0 172 5 1 1 1667
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 1502 1668
0 176 5 2 1 175
0 177 7 1 2 1594 1671
0 178 5 1 1 177
0 179 7 2 2 1669 178
0 180 5 1 1 1673
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 1504 1674
0 184 5 2 1 183
0 185 7 1 2 1596 1677
0 186 5 1 1 185
0 187 7 2 2 1675 186
0 188 5 1 1 1679
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 1506 1680
0 192 5 2 1 191
0 193 7 1 2 1598 1683
0 194 5 1 1 193
0 195 7 2 2 1681 194
0 196 5 1 1 1685
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 1508 1686
0 200 5 2 1 199
0 201 7 1 2 1600 1689
0 202 5 1 1 201
0 203 7 2 2 1687 202
0 204 5 1 1 1691
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 1510 1692
0 208 5 2 1 207
0 209 7 1 2 1602 1695
0 210 5 1 1 209
0 211 7 2 2 1693 210
0 212 5 1 1 1697
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 1512 1698
0 216 5 2 1 215
0 217 7 1 2 1604 1701
0 218 5 1 1 217
0 219 7 4 2 1699 218
0 220 5 2 1 1703
0 221 7 2 2 1579 1707
0 222 5 4 1 1709
0 223 7 1 2 1606 1704
0 224 5 4 1 223
0 225 7 2 2 1700 1702
0 226 5 1 1 1719
0 227 7 1 2 1544 226
0 228 5 1 1 227
0 229 7 1 2 1605 1720
0 230 5 1 1 229
0 231 7 4 2 228 230
0 232 5 3 1 1721
0 233 7 1 2 1577 1722
0 234 5 3 1 233
0 235 7 1 2 97 1725
0 236 5 3 1 235
0 237 7 2 2 1694 1696
0 238 5 1 1 1734
0 239 7 1 2 1542 1735
0 240 5 1 1 239
0 241 7 1 2 1603 238
0 242 5 1 1 241
0 243 7 4 2 240 242
0 244 5 3 1 1736
0 245 7 1 2 1575 1740
0 246 5 3 1 245
0 247 7 1 2 96 1737
0 248 5 3 1 247
0 249 7 2 2 1688 1690
0 250 5 1 1 1749
0 251 7 1 2 1540 1750
0 252 5 1 1 251
0 253 7 1 2 1601 250
0 254 5 1 1 253
0 255 7 4 2 252 254
0 256 5 3 1 1751
0 257 7 1 2 1573 1755
0 258 5 3 1 257
0 259 7 1 2 95 1752
0 260 5 3 1 259
0 261 7 2 2 1682 1684
0 262 5 1 1 1764
0 263 7 1 2 1538 1765
0 264 5 1 1 263
0 265 7 1 2 1599 262
0 266 5 1 1 265
0 267 7 4 2 264 266
0 268 5 2 1 1766
0 269 7 1 2 1571 1770
0 270 5 3 1 269
0 271 7 1 2 94 1767
0 272 5 3 1 271
0 273 7 2 2 1676 1678
0 274 5 1 1 1778
0 275 7 1 2 1536 1779
0 276 5 1 1 275
0 277 7 1 2 1597 274
0 278 5 1 1 277
0 279 7 4 2 276 278
0 280 5 3 1 1780
0 281 7 1 2 1569 1784
0 282 5 3 1 281
0 283 7 1 2 93 1781
0 284 5 3 1 283
0 285 7 2 2 1670 1672
0 286 5 1 1 1793
0 287 7 1 2 1534 1794
0 288 5 1 1 287
0 289 7 1 2 1595 286
0 290 5 1 1 289
0 291 7 3 2 288 290
0 292 5 3 1 1795
0 293 7 1 2 1567 1798
0 294 5 3 1 293
0 295 7 1 2 92 1796
0 296 5 3 1 295
0 297 7 2 2 1664 1666
0 298 5 1 1 1807
0 299 7 1 2 1532 1808
0 300 5 1 1 299
0 301 7 1 2 1593 298
0 302 5 1 1 301
0 303 7 4 2 300 302
0 304 5 3 1 1809
0 305 7 1 2 1565 1813
0 306 5 3 1 305
0 307 7 1 2 91 1810
0 308 5 3 1 307
0 309 7 2 2 1658 1660
0 310 5 1 1 1822
0 311 7 1 2 1530 1823
0 312 5 1 1 311
0 313 7 1 2 1591 310
0 314 5 1 1 313
0 315 7 3 2 312 314
0 316 5 3 1 1824
0 317 7 1 2 1563 1827
0 318 5 3 1 317
0 319 7 1 2 90 1825
0 320 5 3 1 319
0 321 7 2 2 1652 1654
0 322 5 1 1 1836
0 323 7 1 2 1528 1837
0 324 5 1 1 323
0 325 7 1 2 1589 322
0 326 5 1 1 325
0 327 7 4 2 324 326
0 328 5 3 1 1838
0 329 7 1 2 1561 1842
0 330 5 3 1 329
0 331 7 1 2 89 1839
0 332 5 3 1 331
0 333 7 2 2 1646 1648
0 334 5 1 1 1851
0 335 7 1 2 1526 1852
0 336 5 1 1 335
0 337 7 1 2 1587 334
0 338 5 1 1 337
0 339 7 2 2 336 338
0 340 5 3 1 1853
0 341 7 1 2 1559 1855
0 342 5 3 1 341
0 343 7 1 2 88 1854
0 344 5 3 1 343
0 345 7 2 2 1640 1642
0 346 5 1 1 1864
0 347 7 1 2 1524 1865
0 348 5 1 1 347
0 349 7 1 2 1585 346
0 350 5 1 1 349
0 351 7 4 2 348 350
0 352 5 3 1 1866
0 353 7 1 2 1557 1870
0 354 5 3 1 353
0 355 7 1 2 87 1867
0 356 5 3 1 355
0 357 7 2 2 1634 1636
0 358 5 1 1 1879
0 359 7 1 2 1522 1880
0 360 5 1 1 359
0 361 7 1 2 1583 358
0 362 5 1 1 361
0 363 7 2 2 360 362
0 364 5 3 1 1881
0 365 7 1 2 1555 1883
0 366 5 3 1 365
0 367 7 1 2 86 1882
0 368 5 3 1 367
0 369 7 2 2 1628 1630
0 370 5 1 1 1892
0 371 7 1 2 1520 1893
0 372 5 1 1 371
0 373 7 1 2 1581 370
0 374 5 1 1 373
0 375 7 4 2 372 374
0 376 5 3 1 1894
0 377 7 1 2 1553 1898
0 378 5 3 1 377
0 379 7 1 2 85 1895
0 380 5 3 1 379
0 381 7 2 2 1609 1611
0 382 5 1 1 1907
0 383 7 1 2 1622 382
0 384 5 1 1 383
0 385 7 1 2 1624 1908
0 386 5 1 1 385
0 387 7 4 2 384 386
0 388 5 1 1 1909
0 389 7 1 2 1551 1910
0 390 5 3 1 389
0 391 7 1 2 84 388
0 392 5 3 1 391
0 393 7 2 2 1613 1615
0 394 5 1 1 1919
0 395 7 1 2 1617 394
0 396 5 1 1 395
0 397 7 1 2 1619 1920
0 398 5 1 1 397
0 399 7 4 2 396 398
0 400 5 3 1 1921
0 401 7 1 2 1549 1922
0 402 5 3 1 401
0 403 7 1 2 83 1925
0 404 5 3 1 403
0 405 7 1 2 50 66
0 406 5 1 1 405
0 407 7 3 2 1620 406
0 408 5 2 1 1934
0 409 7 2 2 82 1935
0 410 5 3 1 1939
0 411 7 1 2 1931 1941
0 412 5 1 1 411
0 413 7 2 2 1928 412
0 414 5 2 1 1944
0 415 7 1 2 1916 1946
0 416 5 1 1 415
0 417 7 2 2 1913 416
0 418 5 2 1 1948
0 419 7 1 2 1904 1950
0 420 5 1 1 419
0 421 7 2 2 1901 420
0 422 5 2 1 1952
0 423 7 1 2 1889 1954
0 424 5 1 1 423
0 425 7 2 2 1886 424
0 426 5 2 1 1956
0 427 7 1 2 1876 1958
0 428 5 1 1 427
0 429 7 2 2 1873 428
0 430 5 2 1 1960
0 431 7 1 2 1861 1962
0 432 5 1 1 431
0 433 7 2 2 1858 432
0 434 5 2 1 1964
0 435 7 1 2 1848 1966
0 436 5 1 1 435
0 437 7 2 2 1845 436
0 438 5 2 1 1968
0 439 7 1 2 1833 1970
0 440 5 1 1 439
0 441 7 2 2 1830 440
0 442 5 2 1 1972
0 443 7 1 2 1819 1974
0 444 5 1 1 443
0 445 7 2 2 1816 444
0 446 5 2 1 1976
0 447 7 1 2 1804 1978
0 448 5 1 1 447
0 449 7 2 2 1801 448
0 450 5 2 1 1980
0 451 7 1 2 1790 1982
0 452 5 1 1 451
0 453 7 2 2 1787 452
0 454 5 2 1 1984
0 455 7 1 2 1775 1986
0 456 5 1 1 455
0 457 7 2 2 1772 456
0 458 5 2 1 1988
0 459 7 1 2 1761 1990
0 460 5 1 1 459
0 461 7 2 2 1758 460
0 462 5 2 1 1992
0 463 7 1 2 1746 1994
0 464 5 1 1 463
0 465 7 2 2 1743 464
0 466 5 2 1 1996
0 467 7 1 2 1731 1998
0 468 5 1 1 467
0 469 7 3 2 1728 468
0 470 5 3 1 2000
0 471 7 1 2 1715 2003
0 472 5 1 1 471
0 473 7 2 2 1711 472
0 474 5 2 1 2006
0 475 7 3 2 1729 1732
0 476 5 2 1 2010
0 477 7 1 2 1997 2013
0 478 5 1 1 477
0 479 7 1 2 1999 2011
0 480 5 1 1 479
0 481 7 3 2 478 480
0 482 5 2 1 2015
0 483 7 1 2 2007 2016
0 484 5 2 1 483
0 485 7 3 2 1744 1747
0 486 5 2 1 2022
0 487 7 1 2 1993 2025
0 488 5 1 1 487
0 489 7 1 2 1995 2023
0 490 5 1 1 489
0 491 7 3 2 488 490
0 492 5 2 1 2027
0 493 7 3 2 1712 1716
0 494 5 2 1 2032
0 495 7 1 2 2004 2033
0 496 5 1 1 495
0 497 7 1 2 2001 2035
0 498 5 1 1 497
0 499 7 2 2 496 498
0 500 5 1 1 2037
0 501 7 1 2 2028 2038
0 502 5 2 1 501
0 503 7 3 2 1759 1762
0 504 5 2 1 2041
0 505 7 1 2 1989 2044
0 506 5 1 1 505
0 507 7 1 2 1991 2042
0 508 5 1 1 507
0 509 7 3 2 506 508
0 510 5 2 1 2046
0 511 7 1 2 2017 2047
0 512 5 2 1 511
0 513 7 3 2 1773 1776
0 514 5 2 1 2053
0 515 7 1 2 1985 2056
0 516 5 1 1 515
0 517 7 1 2 1987 2054
0 518 5 1 1 517
0 519 7 3 2 516 518
0 520 5 2 1 2058
0 521 7 1 2 2029 2059
0 522 5 2 1 521
0 523 7 3 2 1788 1791
0 524 5 2 1 2065
0 525 7 1 2 1981 2068
0 526 5 1 1 525
0 527 7 1 2 1983 2066
0 528 5 1 1 527
0 529 7 3 2 526 528
0 530 5 2 1 2070
0 531 7 1 2 2048 2071
0 532 5 2 1 531
0 533 7 3 2 1802 1805
0 534 5 2 1 2077
0 535 7 1 2 1977 2080
0 536 5 1 1 535
0 537 7 1 2 1979 2078
0 538 5 1 1 537
0 539 7 3 2 536 538
0 540 5 2 1 2082
0 541 7 1 2 2060 2083
0 542 5 2 1 541
0 543 7 3 2 1817 1820
0 544 5 2 1 2089
0 545 7 1 2 1973 2092
0 546 5 1 1 545
0 547 7 1 2 1975 2090
0 548 5 1 1 547
0 549 7 3 2 546 548
0 550 5 2 1 2094
0 551 7 1 2 2072 2095
0 552 5 2 1 551
0 553 7 3 2 1831 1834
0 554 5 2 1 2101
0 555 7 1 2 1969 2104
0 556 5 1 1 555
0 557 7 1 2 1971 2102
0 558 5 1 1 557
0 559 7 3 2 556 558
0 560 5 2 1 2106
0 561 7 1 2 2084 2107
0 562 5 2 1 561
0 563 7 3 2 1846 1849
0 564 5 2 1 2113
0 565 7 1 2 1965 2116
0 566 5 1 1 565
0 567 7 1 2 1967 2114
0 568 5 1 1 567
0 569 7 3 2 566 568
0 570 5 2 1 2118
0 571 7 1 2 2096 2119
0 572 5 2 1 571
0 573 7 3 2 1859 1862
0 574 5 2 1 2125
0 575 7 1 2 1961 2128
0 576 5 1 1 575
0 577 7 1 2 1963 2126
0 578 5 1 1 577
0 579 7 3 2 576 578
0 580 5 2 1 2130
0 581 7 1 2 2108 2131
0 582 5 2 1 581
0 583 7 3 2 1874 1877
0 584 5 2 1 2137
0 585 7 1 2 1957 2140
0 586 5 1 1 585
0 587 7 1 2 1959 2138
0 588 5 1 1 587
0 589 7 3 2 586 588
0 590 5 2 1 2142
0 591 7 1 2 2120 2143
0 592 5 2 1 591
0 593 7 3 2 1887 1890
0 594 5 2 1 2149
0 595 7 1 2 1953 2152
0 596 5 1 1 595
0 597 7 1 2 1955 2150
0 598 5 1 1 597
0 599 7 3 2 596 598
0 600 5 2 1 2154
0 601 7 1 2 2132 2155
0 602 5 2 1 601
0 603 7 3 2 1902 1905
0 604 5 2 1 2161
0 605 7 1 2 1949 2164
0 606 5 1 1 605
0 607 7 1 2 1951 2162
0 608 5 1 1 607
0 609 7 3 2 606 608
0 610 5 2 1 2166
0 611 7 1 2 2144 2167
0 612 5 2 1 611
0 613 7 3 2 1914 1917
0 614 5 2 1 2173
0 615 7 1 2 1945 2176
0 616 5 1 1 615
0 617 7 1 2 1947 2174
0 618 5 1 1 617
0 619 7 3 2 616 618
0 620 5 2 1 2178
0 621 7 1 2 2156 2179
0 622 5 2 1 621
0 623 7 3 2 1929 1932
0 624 5 2 1 2185
0 625 7 1 2 1942 2186
0 626 5 1 1 625
0 627 7 1 2 1940 2188
0 628 5 1 1 627
0 629 7 2 2 626 628
0 630 5 1 1 2190
0 631 7 1 2 2168 2191
0 632 5 2 1 631
0 633 7 2 2 1546 1937
0 634 5 3 1 2194
0 635 7 3 2 1943 2196
0 636 5 2 1 2199
0 637 7 2 2 2180 2202
0 638 5 2 1 2204
0 639 7 1 2 2169 630
0 640 5 1 1 639
0 641 7 2 2 2192 640
0 642 5 1 1 2208
0 643 7 1 2 2205 2209
0 644 5 2 1 643
0 645 7 2 2 2193 2210
0 646 5 1 1 2212
0 647 7 1 2 2157 2181
0 648 5 1 1 647
0 649 7 2 2 2183 648
0 650 5 1 1 2214
0 651 7 1 2 646 2215
0 652 5 2 1 651
0 653 7 2 2 2184 2216
0 654 5 1 1 2218
0 655 7 1 2 2145 2170
0 656 5 1 1 655
0 657 7 2 2 2171 656
0 658 5 1 1 2220
0 659 7 1 2 654 2221
0 660 5 2 1 659
0 661 7 2 2 2172 2222
0 662 5 1 1 2224
0 663 7 1 2 2133 2158
0 664 5 1 1 663
0 665 7 2 2 2159 664
0 666 5 1 1 2226
0 667 7 1 2 662 2227
0 668 5 2 1 667
0 669 7 2 2 2160 2228
0 670 5 1 1 2230
0 671 7 1 2 2121 2146
0 672 5 1 1 671
0 673 7 2 2 2147 672
0 674 5 1 1 2232
0 675 7 1 2 670 2233
0 676 5 2 1 675
0 677 7 2 2 2148 2234
0 678 5 1 1 2236
0 679 7 1 2 2109 2134
0 680 5 1 1 679
0 681 7 2 2 2135 680
0 682 5 1 1 2238
0 683 7 1 2 678 2239
0 684 5 2 1 683
0 685 7 2 2 2136 2240
0 686 5 1 1 2242
0 687 7 1 2 2097 2122
0 688 5 1 1 687
0 689 7 2 2 2123 688
0 690 5 1 1 2244
0 691 7 1 2 686 2245
0 692 5 2 1 691
0 693 7 2 2 2124 2246
0 694 5 1 1 2248
0 695 7 1 2 2085 2110
0 696 5 1 1 695
0 697 7 2 2 2111 696
0 698 5 1 1 2250
0 699 7 1 2 694 2251
0 700 5 2 1 699
0 701 7 2 2 2112 2252
0 702 5 1 1 2254
0 703 7 1 2 2073 2098
0 704 5 1 1 703
0 705 7 2 2 2099 704
0 706 5 1 1 2256
0 707 7 1 2 702 2257
0 708 5 2 1 707
0 709 7 2 2 2100 2258
0 710 5 1 1 2260
0 711 7 1 2 2061 2086
0 712 5 1 1 711
0 713 7 2 2 2087 712
0 714 5 1 1 2262
0 715 7 1 2 710 2263
0 716 5 2 1 715
0 717 7 2 2 2088 2264
0 718 5 1 1 2266
0 719 7 1 2 2049 2074
0 720 5 1 1 719
0 721 7 2 2 2075 720
0 722 5 1 1 2268
0 723 7 1 2 718 2269
0 724 5 2 1 723
0 725 7 2 2 2076 2270
0 726 5 1 1 2272
0 727 7 1 2 2030 2062
0 728 5 1 1 727
0 729 7 2 2 2063 728
0 730 5 1 1 2274
0 731 7 1 2 726 2275
0 732 5 2 1 731
0 733 7 2 2 2064 2276
0 734 5 1 1 2278
0 735 7 1 2 2018 2050
0 736 5 1 1 735
0 737 7 2 2 2051 736
0 738 5 1 1 2280
0 739 7 1 2 734 2281
0 740 5 2 1 739
0 741 7 2 2 2052 2282
0 742 5 1 1 2284
0 743 7 1 2 2031 500
0 744 5 1 1 743
0 745 7 2 2 2039 744
0 746 5 1 1 2286
0 747 7 1 2 742 2287
0 748 5 2 1 747
0 749 7 2 2 2040 2288
0 750 5 1 1 2290
0 751 7 1 2 2008 2019
0 752 5 1 1 751
0 753 7 2 2 2020 752
0 754 5 1 1 2292
0 755 7 1 2 750 2293
0 756 5 2 1 755
0 757 7 2 2 2021 2294
0 758 5 1 1 2296
0 759 7 1 2 1717 2002
0 760 5 1 1 759
0 761 7 1 2 1713 2005
0 762 5 1 1 761
0 763 7 2 2 760 762
0 764 5 1 1 2298
0 765 7 1 2 758 2299
0 766 5 2 1 765
0 767 7 1 2 2297 764
0 768 5 2 1 767
0 769 7 1 2 2300 2302
0 770 5 1 1 769
0 771 7 1 2 1705 770
0 772 5 1 1 771
0 773 7 1 2 2291 754
0 774 5 1 1 773
0 775 7 2 2 2295 774
0 776 5 1 1 2304
0 777 7 1 2 1723 2305
0 778 5 1 1 777
0 779 7 1 2 2285 746
0 780 5 1 1 779
0 781 7 2 2 2289 780
0 782 5 1 1 2306
0 783 7 1 2 1738 782
0 784 5 1 1 783
0 785 7 1 2 1741 2307
0 786 5 1 1 785
0 787 7 1 2 2279 738
0 788 5 1 1 787
0 789 7 1 2 2283 788
0 790 5 1 1 789
0 791 7 1 2 2273 730
0 792 5 1 1 791
0 793 7 2 2 2277 792
0 794 5 1 1 2308
0 795 7 1 2 2267 722
0 796 5 1 1 795
0 797 7 1 2 2271 796
0 798 5 1 1 797
0 799 7 1 2 2255 706
0 800 5 1 1 799
0 801 7 2 2 2259 800
0 802 5 1 1 2310
0 803 7 1 2 1811 802
0 804 5 1 1 803
0 805 7 1 2 1814 2311
0 806 5 1 1 805
0 807 7 1 2 2249 698
0 808 5 1 1 807
0 809 7 2 2 2253 808
0 810 5 1 1 2312
0 811 7 1 2 1828 2313
0 812 5 1 1 811
0 813 7 1 2 2243 690
0 814 5 1 1 813
0 815 7 2 2 2247 814
0 816 5 1 1 2314
0 817 7 1 2 1843 2315
0 818 5 1 1 817
0 819 7 1 2 1840 816
0 820 5 1 1 819
0 821 7 1 2 2237 682
0 822 5 1 1 821
0 823 7 2 2 2241 822
0 824 5 1 1 2316
0 825 7 1 2 2231 674
0 826 5 1 1 825
0 827 7 2 2 2235 826
0 828 5 1 1 2318
0 829 7 1 2 1871 2319
0 830 5 1 1 829
0 831 7 1 2 1868 828
0 832 5 1 1 831
0 833 7 1 2 2225 666
0 834 5 1 1 833
0 835 7 2 2 2229 834
0 836 5 1 1 2320
0 837 7 1 2 2219 658
0 838 5 1 1 837
0 839 7 2 2 2223 838
0 840 5 1 1 2322
0 841 7 1 2 1899 2323
0 842 5 1 1 841
0 843 7 1 2 1896 840
0 844 5 1 1 843
0 845 7 1 2 2213 650
0 846 5 1 1 845
0 847 7 2 2 2217 846
0 848 5 1 1 2324
0 849 7 2 2 2187 2197
0 850 5 2 1 2326
0 851 7 2 2 1547 2327
0 852 5 1 1 2330
0 853 7 1 2 1936 2331
0 854 5 1 1 853
0 855 7 1 2 1938 2328
0 856 5 2 1 855
0 857 7 1 2 2182 2200
0 858 5 1 1 857
0 859 7 1 2 2206 858
0 860 5 1 1 859
0 861 7 1 2 2332 860
0 862 5 1 1 861
0 863 7 1 2 854 862
0 864 5 1 1 863
0 865 7 1 2 2207 642
0 866 5 1 1 865
0 867 7 2 2 2211 866
0 868 5 1 1 2334
0 869 7 1 2 1923 2335
0 870 5 1 1 869
0 871 7 1 2 864 870
0 872 5 1 1 871
0 873 7 1 2 1926 868
0 874 5 1 1 873
0 875 7 2 2 872 874
0 876 5 1 1 2336
0 877 7 1 2 848 876
0 878 5 1 1 877
0 879 7 1 2 1911 878
0 880 5 1 1 879
0 881 7 1 2 2325 2337
0 882 5 1 1 881
0 883 7 1 2 880 882
0 884 5 1 1 883
0 885 7 1 2 844 884
0 886 5 1 1 885
0 887 7 2 2 842 886
0 888 5 1 1 2338
0 889 7 1 2 2321 888
0 890 5 1 1 889
0 891 7 1 2 836 2339
0 892 5 1 1 891
0 893 7 1 2 1884 892
0 894 5 1 1 893
0 895 7 1 2 890 894
0 896 5 1 1 895
0 897 7 1 2 832 896
0 898 5 1 1 897
0 899 7 2 2 830 898
0 900 5 1 1 2340
0 901 7 1 2 2317 900
0 902 5 1 1 901
0 903 7 1 2 824 2341
0 904 5 1 1 903
0 905 7 1 2 1856 904
0 906 5 1 1 905
0 907 7 1 2 902 906
0 908 5 1 1 907
0 909 7 1 2 820 908
0 910 5 1 1 909
0 911 7 1 2 818 910
0 912 7 1 2 812 911
0 913 5 1 1 912
0 914 7 1 2 1826 810
0 915 5 1 1 914
0 916 7 1 2 913 915
0 917 5 1 1 916
0 918 7 1 2 806 917
0 919 5 1 1 918
0 920 7 2 2 804 919
0 921 5 1 1 2342
0 922 7 1 2 1799 2343
0 923 5 1 1 922
0 924 7 1 2 1797 921
0 925 5 1 1 924
0 926 7 1 2 2261 714
0 927 5 1 1 926
0 928 7 1 2 2265 927
0 929 7 1 2 925 928
0 930 5 1 1 929
0 931 7 2 2 923 930
0 932 5 1 1 2344
0 933 7 1 2 1785 932
0 934 5 1 1 933
0 935 7 1 2 798 934
0 936 5 1 1 935
0 937 7 1 2 1782 2345
0 938 5 1 1 937
0 939 7 2 2 936 938
0 940 5 1 1 2346
0 941 7 1 2 2309 2347
0 942 5 1 1 941
0 943 7 1 2 1768 942
0 944 5 1 1 943
0 945 7 1 2 794 940
0 946 5 1 1 945
0 947 7 2 2 944 946
0 948 5 1 1 2348
0 949 7 1 2 1756 2349
0 950 5 1 1 949
0 951 7 1 2 790 950
0 952 5 1 1 951
0 953 7 1 2 1753 948
0 954 5 1 1 953
0 955 7 1 2 952 954
0 956 5 1 1 955
0 957 7 1 2 786 956
0 958 5 1 1 957
0 959 7 1 2 784 958
0 960 5 1 1 959
0 961 7 1 2 778 960
0 962 5 1 1 961
0 963 7 1 2 1726 776
0 964 5 1 1 963
0 965 7 1 2 962 964
0 966 7 1 2 772 965
0 967 5 1 1 966
0 968 7 1 2 1708 2303
0 969 5 1 1 968
0 970 7 1 2 2009 2301
0 971 7 1 2 969 970
0 972 7 1 2 967 971
0 973 5 1 1 972
0 974 7 1 2 1930 2198
0 975 5 1 1 974
0 976 7 2 2 1933 975
0 977 5 2 1 2350
0 978 7 1 2 1915 2352
0 979 5 1 1 978
0 980 7 3 2 1918 979
0 981 5 1 1 2354
0 982 7 1 2 1906 2355
0 983 5 1 1 982
0 984 7 2 2 1903 983
0 985 5 2 1 2357
0 986 7 1 2 1891 2359
0 987 5 1 1 986
0 988 7 2 2 1888 987
0 989 5 2 1 2361
0 990 7 1 2 1878 2363
0 991 5 1 1 990
0 992 7 2 2 1875 991
0 993 5 2 1 2365
0 994 7 1 2 1863 2367
0 995 5 1 1 994
0 996 7 2 2 1860 995
0 997 5 2 1 2369
0 998 7 1 2 1850 2371
0 999 5 1 1 998
0 1000 7 2 2 1847 999
0 1001 5 2 1 2373
0 1002 7 1 2 1835 2375
0 1003 5 1 1 1002
0 1004 7 2 2 1832 1003
0 1005 5 2 1 2377
0 1006 7 1 2 1821 2379
0 1007 5 1 1 1006
0 1008 7 2 2 1818 1007
0 1009 5 2 1 2381
0 1010 7 1 2 1806 2383
0 1011 5 1 1 1010
0 1012 7 2 2 1803 1011
0 1013 5 2 1 2385
0 1014 7 1 2 1792 2387
0 1015 5 1 1 1014
0 1016 7 2 2 1789 1015
0 1017 5 2 1 2389
0 1018 7 1 2 1777 2391
0 1019 5 1 1 1018
0 1020 7 2 2 1774 1019
0 1021 5 2 1 2393
0 1022 7 1 2 1763 2395
0 1023 5 1 1 1022
0 1024 7 2 2 1760 1023
0 1025 5 2 1 2397
0 1026 7 1 2 1748 2399
0 1027 5 1 1 1026
0 1028 7 2 2 1745 1027
0 1029 5 2 1 2401
0 1030 7 1 2 1733 2403
0 1031 5 1 1 1030
0 1032 7 3 2 1730 1031
0 1033 5 3 1 2405
0 1034 7 1 2 1718 2408
0 1035 5 1 1 1034
0 1036 7 3 2 1714 1035
0 1037 5 2 1 2411
0 1038 7 1 2 973 2414
0 1039 5 1 1 1038
0 1040 7 1 2 2026 2398
0 1041 5 1 1 1040
0 1042 7 1 2 2024 2400
0 1043 5 1 1 1042
0 1044 7 3 2 1041 1043
0 1045 5 2 1 2416
0 1046 7 1 2 2036 2406
0 1047 5 1 1 1046
0 1048 7 1 2 2034 2409
0 1049 5 1 1 1048
0 1050 7 2 2 1047 1049
0 1051 5 1 1 2421
0 1052 7 1 2 2419 1051
0 1053 5 2 1 1052
0 1054 7 1 2 2045 2394
0 1055 5 1 1 1054
0 1056 7 1 2 2043 2396
0 1057 5 1 1 1056
0 1058 7 3 2 1055 1057
0 1059 5 2 1 2425
0 1060 7 1 2 2014 2402
0 1061 5 1 1 1060
0 1062 7 1 2 2012 2404
0 1063 5 1 1 1062
0 1064 7 3 2 1061 1063
0 1065 5 2 1 2430
0 1066 7 1 2 2428 2433
0 1067 5 2 1 1066
0 1068 7 1 2 2057 2390
0 1069 5 1 1 1068
0 1070 7 1 2 2055 2392
0 1071 5 1 1 1070
0 1072 7 3 2 1069 1071
0 1073 5 2 1 2437
0 1074 7 1 2 2420 2440
0 1075 5 2 1 1074
0 1076 7 1 2 2069 2386
0 1077 5 1 1 1076
0 1078 7 1 2 2067 2388
0 1079 5 1 1 1078
0 1080 7 3 2 1077 1079
0 1081 5 2 1 2444
0 1082 7 1 2 2429 2447
0 1083 5 2 1 1082
0 1084 7 1 2 2081 2382
0 1085 5 1 1 1084
0 1086 7 1 2 2079 2384
0 1087 5 1 1 1086
0 1088 7 3 2 1085 1087
0 1089 5 2 1 2451
0 1090 7 1 2 2441 2454
0 1091 5 2 1 1090
0 1092 7 1 2 2093 2378
0 1093 5 1 1 1092
0 1094 7 1 2 2091 2380
0 1095 5 1 1 1094
0 1096 7 3 2 1093 1095
0 1097 5 2 1 2458
0 1098 7 1 2 2448 2461
0 1099 5 2 1 1098
0 1100 7 1 2 2105 2374
0 1101 5 1 1 1100
0 1102 7 1 2 2103 2376
0 1103 5 1 1 1102
0 1104 7 3 2 1101 1103
0 1105 5 2 1 2465
0 1106 7 1 2 2455 2468
0 1107 5 2 1 1106
0 1108 7 1 2 2117 2370
0 1109 5 1 1 1108
0 1110 7 1 2 2115 2372
0 1111 5 1 1 1110
0 1112 7 3 2 1109 1111
0 1113 5 2 1 2472
0 1114 7 1 2 2462 2475
0 1115 5 2 1 1114
0 1116 7 1 2 2129 2366
0 1117 5 1 1 1116
0 1118 7 1 2 2127 2368
0 1119 5 1 1 1118
0 1120 7 3 2 1117 1119
0 1121 5 2 1 2479
0 1122 7 1 2 2469 2482
0 1123 5 2 1 1122
0 1124 7 1 2 2141 2362
0 1125 5 1 1 1124
0 1126 7 1 2 2139 2364
0 1127 5 1 1 1126
0 1128 7 3 2 1125 1127
0 1129 5 2 1 2486
0 1130 7 1 2 2476 2489
0 1131 5 2 1 1130
0 1132 7 1 2 2153 2358
0 1133 5 1 1 1132
0 1134 7 1 2 2151 2360
0 1135 5 1 1 1134
0 1136 7 3 2 1133 1135
0 1137 5 2 1 2493
0 1138 7 1 2 2483 2496
0 1139 5 2 1 1138
0 1140 7 1 2 2163 981
0 1141 5 1 1 1140
0 1142 7 1 2 2165 2356
0 1143 5 1 1 1142
0 1144 7 3 2 1141 1143
0 1145 5 2 1 2500
0 1146 7 1 2 2490 2501
0 1147 5 2 1 1146
0 1148 7 1 2 2175 2353
0 1149 5 1 1 1148
0 1150 7 1 2 2177 2351
0 1151 5 1 1 1150
0 1152 7 4 2 1149 1151
0 1153 5 1 1 2507
0 1154 7 1 2 2497 2508
0 1155 5 2 1 1154
0 1156 7 1 2 2189 2195
0 1157 5 1 1 1156
0 1158 7 2 2 2329 1157
0 1159 5 1 1 2513
0 1160 7 1 2 2502 2514
0 1161 5 2 1 1160
0 1162 7 2 2 2203 2509
0 1163 5 2 1 2517
0 1164 7 1 2 2503 1159
0 1165 5 1 1 1164
0 1166 7 2 2 2515 1165
0 1167 5 1 1 2521
0 1168 7 1 2 2518 2522
0 1169 5 2 1 1168
0 1170 7 2 2 2516 2523
0 1171 5 1 1 2525
0 1172 7 1 2 2494 1153
0 1173 5 1 1 1172
0 1174 7 2 2 2511 1173
0 1175 5 1 1 2527
0 1176 7 1 2 1171 2528
0 1177 5 2 1 1176
0 1178 7 2 2 2512 2529
0 1179 5 1 1 2531
0 1180 7 1 2 2487 2504
0 1181 5 1 1 1180
0 1182 7 2 2 2505 1181
0 1183 5 1 1 2533
0 1184 7 1 2 1179 2534
0 1185 5 2 1 1184
0 1186 7 2 2 2506 2535
0 1187 5 1 1 2537
0 1188 7 1 2 2480 2495
0 1189 5 1 1 1188
0 1190 7 2 2 2498 1189
0 1191 5 1 1 2539
0 1192 7 1 2 1187 2540
0 1193 5 2 1 1192
0 1194 7 2 2 2499 2541
0 1195 5 1 1 2543
0 1196 7 1 2 2473 2488
0 1197 5 1 1 1196
0 1198 7 2 2 2491 1197
0 1199 5 1 1 2545
0 1200 7 1 2 1195 2546
0 1201 5 2 1 1200
0 1202 7 2 2 2492 2547
0 1203 5 1 1 2549
0 1204 7 1 2 2466 2481
0 1205 5 1 1 1204
0 1206 7 2 2 2484 1205
0 1207 5 1 1 2551
0 1208 7 1 2 1203 2552
0 1209 5 2 1 1208
0 1210 7 2 2 2485 2553
0 1211 5 1 1 2555
0 1212 7 1 2 2459 2474
0 1213 5 1 1 1212
0 1214 7 2 2 2477 1213
0 1215 5 1 1 2557
0 1216 7 1 2 1211 2558
0 1217 5 2 1 1216
0 1218 7 2 2 2478 2559
0 1219 5 1 1 2561
0 1220 7 1 2 2452 2467
0 1221 5 1 1 1220
0 1222 7 2 2 2470 1221
0 1223 5 1 1 2563
0 1224 7 1 2 1219 2564
0 1225 5 2 1 1224
0 1226 7 2 2 2471 2565
0 1227 5 1 1 2567
0 1228 7 1 2 2445 2460
0 1229 5 1 1 1228
0 1230 7 2 2 2463 1229
0 1231 5 1 1 2569
0 1232 7 1 2 1227 2570
0 1233 5 2 1 1232
0 1234 7 2 2 2464 2571
0 1235 5 1 1 2573
0 1236 7 1 2 2438 2453
0 1237 5 1 1 1236
0 1238 7 2 2 2456 1237
0 1239 5 1 1 2575
0 1240 7 1 2 1235 2576
0 1241 5 2 1 1240
0 1242 7 2 2 2457 2577
0 1243 5 1 1 2579
0 1244 7 1 2 2426 2446
0 1245 5 1 1 1244
0 1246 7 2 2 2449 1245
0 1247 5 1 1 2581
0 1248 7 1 2 1243 2582
0 1249 5 2 1 1248
0 1250 7 2 2 2450 2583
0 1251 5 1 1 2585
0 1252 7 1 2 2417 2439
0 1253 5 1 1 1252
0 1254 7 2 2 2442 1253
0 1255 5 1 1 2587
0 1256 7 1 2 1251 2588
0 1257 5 2 1 1256
0 1258 7 2 2 2443 2589
0 1259 5 1 1 2591
0 1260 7 1 2 2427 2431
0 1261 5 1 1 1260
0 1262 7 2 2 2435 1261
0 1263 5 1 1 2593
0 1264 7 1 2 1259 2594
0 1265 5 2 1 1264
0 1266 7 2 2 2436 2595
0 1267 5 1 1 2597
0 1268 7 1 2 2418 2422
0 1269 5 1 1 1268
0 1270 7 2 2 2423 1269
0 1271 5 1 1 2599
0 1272 7 1 2 1267 2600
0 1273 5 2 1 1272
0 1274 7 2 2 2424 2601
0 1275 5 1 1 2603
0 1276 7 1 2 2415 2432
0 1277 5 1 1 1276
0 1278 7 1 2 2412 2434
0 1279 5 1 1 1278
0 1280 7 2 2 1277 1279
0 1281 5 1 1 2605
0 1282 7 1 2 2604 2606
0 1283 5 1 1 1282
0 1284 7 1 2 1607 2407
0 1285 5 1 1 1284
0 1286 7 2 2 1706 1285
0 1287 5 1 1 2607
0 1288 7 2 2 1283 1287
0 1289 5 1 1 2609
0 1290 7 1 2 1275 1281
0 1291 5 2 1 1290
0 1292 7 1 2 2608 2611
0 1293 5 1 1 1292
0 1294 7 1 2 1724 1293
0 1295 5 1 1 1294
0 1296 7 1 2 1289 1295
0 1297 5 1 1 1296
0 1298 7 1 2 2598 1271
0 1299 5 1 1 1298
0 1300 7 2 2 2602 1299
0 1301 5 1 1 2613
0 1302 7 1 2 1742 2614
0 1303 5 1 1 1302
0 1304 7 1 2 2586 1255
0 1305 5 1 1 1304
0 1306 7 2 2 2590 1305
0 1307 5 1 1 2615
0 1308 7 1 2 1769 1307
0 1309 5 1 1 1308
0 1310 7 1 2 1771 2616
0 1311 5 1 1 1310
0 1312 7 1 2 2580 1247
0 1313 5 1 1 1312
0 1314 7 2 2 2584 1313
0 1315 5 1 1 2617
0 1316 7 1 2 1783 1315
0 1317 5 1 1 1316
0 1318 7 1 2 1786 2618
0 1319 5 1 1 1318
0 1320 7 1 2 2574 1239
0 1321 5 1 1 1320
0 1322 7 2 2 2578 1321
0 1323 5 1 1 2619
0 1324 7 1 2 2568 1231
0 1325 5 1 1 1324
0 1326 7 2 2 2572 1325
0 1327 5 1 1 2621
0 1328 7 1 2 1815 2622
0 1329 5 1 1 1328
0 1330 7 1 2 1812 1327
0 1331 5 1 1 1330
0 1332 7 1 2 2562 1223
0 1333 5 1 1 1332
0 1334 7 2 2 2566 1333
0 1335 5 1 1 2623
0 1336 7 1 2 2556 1215
0 1337 5 1 1 1336
0 1338 7 2 2 2560 1337
0 1339 5 1 1 2625
0 1340 7 1 2 1844 2626
0 1341 5 1 1 1340
0 1342 7 1 2 1841 1339
0 1343 5 1 1 1342
0 1344 7 1 2 2550 1207
0 1345 5 1 1 1344
0 1346 7 2 2 2554 1345
0 1347 5 1 1 2627
0 1348 7 1 2 2544 1199
0 1349 5 1 1 1348
0 1350 7 2 2 2548 1349
0 1351 5 1 1 2629
0 1352 7 1 2 1872 2630
0 1353 5 1 1 1352
0 1354 7 1 2 1869 1351
0 1355 5 1 1 1354
0 1356 7 1 2 2538 1191
0 1357 5 1 1 1356
0 1358 7 2 2 2542 1357
0 1359 5 1 1 2631
0 1360 7 1 2 2532 1183
0 1361 5 1 1 1360
0 1362 7 2 2 2536 1361
0 1363 5 1 1 2633
0 1364 7 1 2 1900 2634
0 1365 5 1 1 1364
0 1366 7 1 2 1897 1363
0 1367 5 1 1 1366
0 1368 7 1 2 2526 1175
0 1369 5 1 1 1368
0 1370 7 2 2 2530 1369
0 1371 5 1 1 2635
0 1372 7 1 2 2519 1167
0 1373 5 1 1 1372
0 1374 7 2 2 2524 1373
0 1375 5 1 1 2637
0 1376 7 1 2 1924 2638
0 1377 5 1 1 1376
0 1378 7 1 2 852 2510
0 1379 5 1 1 1378
0 1380 7 1 2 2201 1379
0 1381 5 1 1 1380
0 1382 7 1 2 2520 1381
0 1383 5 1 1 1382
0 1384 7 1 2 2333 1383
0 1385 7 1 2 1377 1384
0 1386 5 1 1 1385
0 1387 7 1 2 1927 1375
0 1388 5 1 1 1387
0 1389 7 2 2 1386 1388
0 1390 5 1 1 2639
0 1391 7 1 2 1371 1390
0 1392 5 1 1 1391
0 1393 7 1 2 1912 1392
0 1394 5 1 1 1393
0 1395 7 1 2 2636 2640
0 1396 5 1 1 1395
0 1397 7 1 2 1394 1396
0 1398 5 1 1 1397
0 1399 7 1 2 1367 1398
0 1400 5 1 1 1399
0 1401 7 2 2 1365 1400
0 1402 5 1 1 2641
0 1403 7 1 2 2632 1402
0 1404 5 1 1 1403
0 1405 7 1 2 1359 2642
0 1406 5 1 1 1405
0 1407 7 1 2 1885 1406
0 1408 5 1 1 1407
0 1409 7 1 2 1404 1408
0 1410 5 1 1 1409
0 1411 7 1 2 1355 1410
0 1412 5 1 1 1411
0 1413 7 2 2 1353 1412
0 1414 5 1 1 2643
0 1415 7 1 2 2628 1414
0 1416 5 1 1 1415
0 1417 7 1 2 1347 2644
0 1418 5 1 1 1417
0 1419 7 1 2 1857 1418
0 1420 5 1 1 1419
0 1421 7 1 2 1416 1420
0 1422 5 1 1 1421
0 1423 7 1 2 1343 1422
0 1424 5 1 1 1423
0 1425 7 2 2 1341 1424
0 1426 5 1 1 2645
0 1427 7 1 2 2624 1426
0 1428 5 1 1 1427
0 1429 7 1 2 1335 2646
0 1430 5 1 1 1429
0 1431 7 1 2 1829 1430
0 1432 5 1 1 1431
0 1433 7 1 2 1428 1432
0 1434 5 1 1 1433
0 1435 7 1 2 1331 1434
0 1436 5 1 1 1435
0 1437 7 2 2 1329 1436
0 1438 5 1 1 2647
0 1439 7 1 2 2620 1438
0 1440 5 1 1 1439
0 1441 7 1 2 1323 2648
0 1442 5 1 1 1441
0 1443 7 1 2 1800 1442
0 1444 5 1 1 1443
0 1445 7 1 2 1440 1444
0 1446 7 1 2 1319 1445
0 1447 5 1 1 1446
0 1448 7 1 2 1317 1447
0 1449 5 1 1 1448
0 1450 7 1 2 1311 1449
0 1451 5 1 1 1450
0 1452 7 2 2 1309 1451
0 1453 5 1 1 2649
0 1454 7 1 2 1757 2650
0 1455 5 1 1 1454
0 1456 7 1 2 1754 1453
0 1457 5 1 1 1456
0 1458 7 1 2 2592 1263
0 1459 5 1 1 1458
0 1460 7 1 2 2596 1459
0 1461 7 1 2 1457 1460
0 1462 5 1 1 1461
0 1463 7 1 2 1455 1462
0 1464 7 1 2 1303 1463
0 1465 5 1 1 1464
0 1466 7 1 2 1739 1301
0 1467 5 1 1 1466
0 1468 7 1 2 1465 1467
0 1469 7 1 2 1297 1468
0 1470 5 1 1 1469
0 1471 7 1 2 1727 2612
0 1472 5 1 1 1471
0 1473 7 1 2 2610 1472
0 1474 5 1 1 1473
0 1475 7 1 2 1710 2410
0 1476 5 1 1 1475
0 1477 7 1 2 1474 1476
0 1478 7 1 2 1470 1477
0 1479 5 1 1 1478
0 1480 7 1 2 2413 1479
0 1481 5 1 1 1480
3 3499 7 0 2 1039 1481
