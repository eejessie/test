1 0 0 8 0
2 32 1 0
2 1937 1 0
2 1938 1 0
2 1939 1 0
2 1940 1 0
2 1941 1 0
2 1942 1 0
2 1943 1 0
1 1 0 9 0
2 1944 1 1
2 1945 1 1
2 1946 1 1
2 1947 1 1
2 1948 1 1
2 1949 1 1
2 1950 1 1
2 1951 1 1
2 1952 1 1
1 2 0 10 0
2 1953 1 2
2 1954 1 2
2 1955 1 2
2 1956 1 2
2 1957 1 2
2 1958 1 2
2 1959 1 2
2 1960 1 2
2 1961 1 2
2 1962 1 2
1 3 0 11 0
2 1963 1 3
2 1964 1 3
2 1965 1 3
2 1966 1 3
2 1967 1 3
2 1968 1 3
2 1969 1 3
2 1970 1 3
2 1971 1 3
2 1972 1 3
2 1973 1 3
1 4 0 10 0
2 1974 1 4
2 1975 1 4
2 1976 1 4
2 1977 1 4
2 1978 1 4
2 1979 1 4
2 1980 1 4
2 1981 1 4
2 1982 1 4
2 1983 1 4
1 5 0 11 0
2 1984 1 5
2 1985 1 5
2 1986 1 5
2 1987 1 5
2 1988 1 5
2 1989 1 5
2 1990 1 5
2 1991 1 5
2 1992 1 5
2 1993 1 5
2 1994 1 5
1 6 0 10 0
2 1995 1 6
2 1996 1 6
2 1997 1 6
2 1998 1 6
2 1999 1 6
2 2000 1 6
2 2001 1 6
2 2002 1 6
2 2003 1 6
2 2004 1 6
1 7 0 10 0
2 2005 1 7
2 2006 1 7
2 2007 1 7
2 2008 1 7
2 2009 1 7
2 2010 1 7
2 2011 1 7
2 2012 1 7
2 2013 1 7
2 2014 1 7
1 8 0 10 0
2 2015 1 8
2 2016 1 8
2 2017 1 8
2 2018 1 8
2 2019 1 8
2 2020 1 8
2 2021 1 8
2 2022 1 8
2 2023 1 8
2 2024 1 8
1 9 0 10 0
2 2025 1 9
2 2026 1 9
2 2027 1 9
2 2028 1 9
2 2029 1 9
2 2030 1 9
2 2031 1 9
2 2032 1 9
2 2033 1 9
2 2034 1 9
1 10 0 11 0
2 2035 1 10
2 2036 1 10
2 2037 1 10
2 2038 1 10
2 2039 1 10
2 2040 1 10
2 2041 1 10
2 2042 1 10
2 2043 1 10
2 2044 1 10
2 2045 1 10
1 11 0 10 0
2 2046 1 11
2 2047 1 11
2 2048 1 11
2 2049 1 11
2 2050 1 11
2 2051 1 11
2 2052 1 11
2 2053 1 11
2 2054 1 11
2 2055 1 11
1 12 0 10 0
2 2056 1 12
2 2057 1 12
2 2058 1 12
2 2059 1 12
2 2060 1 12
2 2061 1 12
2 2062 1 12
2 2063 1 12
2 2064 1 12
2 2065 1 12
1 13 0 10 0
2 2066 1 13
2 2067 1 13
2 2068 1 13
2 2069 1 13
2 2070 1 13
2 2071 1 13
2 2072 1 13
2 2073 1 13
2 2074 1 13
2 2075 1 13
1 14 0 10 0
2 2076 1 14
2 2077 1 14
2 2078 1 14
2 2079 1 14
2 2080 1 14
2 2081 1 14
2 2082 1 14
2 2083 1 14
2 2084 1 14
2 2085 1 14
1 15 0 10 0
2 2086 1 15
2 2087 1 15
2 2088 1 15
2 2089 1 15
2 2090 1 15
2 2091 1 15
2 2092 1 15
2 2093 1 15
2 2094 1 15
2 2095 1 15
1 16 0 3 0
2 2096 1 16
2 2097 1 16
2 2098 1 16
1 17 0 3 0
2 2099 1 17
2 2100 1 17
2 2101 1 17
1 18 0 3 0
2 2102 1 18
2 2103 1 18
2 2104 1 18
1 19 0 3 0
2 2105 1 19
2 2106 1 19
2 2107 1 19
1 20 0 3 0
2 2108 1 20
2 2109 1 20
2 2110 1 20
1 21 0 3 0
2 2111 1 21
2 2112 1 21
2 2113 1 21
1 22 0 3 0
2 2114 1 22
2 2115 1 22
2 2116 1 22
1 23 0 3 0
2 2117 1 23
2 2118 1 23
2 2119 1 23
1 24 0 3 0
2 2120 1 24
2 2121 1 24
2 2122 1 24
1 25 0 3 0
2 2123 1 25
2 2124 1 25
2 2125 1 25
1 26 0 3 0
2 2126 1 26
2 2127 1 26
2 2128 1 26
1 27 0 3 0
2 2129 1 27
2 2130 1 27
2 2131 1 27
1 28 0 4 0
2 2132 1 28
2 2133 1 28
2 2134 1 28
2 2135 1 28
1 29 0 3 0
2 2136 1 29
2 2137 1 29
2 2138 1 29
1 30 0 4 0
2 2139 1 30
2 2140 1 30
2 2141 1 30
2 2142 1 30
1 31 0 4 0
2 2143 1 31
2 2144 1 31
2 2145 1 31
2 2146 1 31
2 2147 1 34
2 2148 1 34
2 2149 1 35
2 2150 1 35
2 2151 1 36
2 2152 1 36
2 2153 1 37
2 2154 1 37
2 2155 1 38
2 2156 1 38
2 2157 1 39
2 2158 1 39
2 2159 1 40
2 2160 1 40
2 2161 1 41
2 2162 1 41
2 2163 1 42
2 2164 1 42
2 2165 1 43
2 2166 1 43
2 2167 1 44
2 2168 1 44
2 2169 1 45
2 2170 1 45
2 2171 1 46
2 2172 1 46
2 2173 1 47
2 2174 1 47
2 2175 1 48
2 2176 1 48
2 2177 1 48
2 2178 1 49
2 2179 1 49
2 2180 1 49
2 2181 1 50
2 2182 1 50
2 2183 1 50
2 2184 1 51
2 2185 1 51
2 2186 1 51
2 2187 1 52
2 2188 1 52
2 2189 1 52
2 2190 1 53
2 2191 1 53
2 2192 1 53
2 2193 1 54
2 2194 1 54
2 2195 1 54
2 2196 1 55
2 2197 1 55
2 2198 1 55
2 2199 1 56
2 2200 1 56
2 2201 1 56
2 2202 1 57
2 2203 1 57
2 2204 1 57
2 2205 1 58
2 2206 1 58
2 2207 1 58
2 2208 1 59
2 2209 1 59
2 2210 1 59
2 2211 1 60
2 2212 1 60
2 2213 1 60
2 2214 1 60
2 2215 1 61
2 2216 1 61
2 2217 1 61
2 2218 1 62
2 2219 1 62
2 2220 1 63
2 2221 1 63
2 2222 1 64
2 2223 1 64
2 2224 1 66
2 2225 1 66
2 2226 1 66
2 2227 1 68
2 2228 1 68
2 2229 1 74
2 2230 1 74
2 2231 1 76
2 2232 1 76
2 2233 1 81
2 2234 1 81
2 2235 1 84
2 2236 1 84
2 2237 1 87
2 2238 1 87
2 2239 1 89
2 2240 1 89
2 2241 1 90
2 2242 1 90
2 2243 1 95
2 2244 1 95
2 2245 1 98
2 2246 1 98
2 2247 1 103
2 2248 1 103
2 2249 1 104
2 2250 1 104
2 2251 1 105
2 2252 1 105
2 2253 1 108
2 2254 1 108
2 2255 1 111
2 2256 1 111
2 2257 1 113
2 2258 1 113
2 2259 1 114
2 2260 1 114
2 2261 1 119
2 2262 1 119
2 2263 1 122
2 2264 1 122
2 2265 1 127
2 2266 1 127
2 2267 1 127
2 2268 1 129
2 2269 1 129
2 2270 1 132
2 2271 1 132
2 2272 1 135
2 2273 1 135
2 2274 1 137
2 2275 1 137
2 2276 1 138
2 2277 1 138
2 2278 1 143
2 2279 1 143
2 2280 1 146
2 2281 1 146
2 2282 1 151
2 2283 1 151
2 2284 1 151
2 2285 1 153
2 2286 1 153
2 2287 1 156
2 2288 1 156
2 2289 1 159
2 2290 1 159
2 2291 1 161
2 2292 1 161
2 2293 1 162
2 2294 1 162
2 2295 1 167
2 2296 1 167
2 2297 1 170
2 2298 1 170
2 2299 1 175
2 2300 1 175
2 2301 1 175
2 2302 1 177
2 2303 1 177
2 2304 1 180
2 2305 1 180
2 2306 1 183
2 2307 1 183
2 2308 1 185
2 2309 1 185
2 2310 1 186
2 2311 1 186
2 2312 1 191
2 2313 1 191
2 2314 1 194
2 2315 1 194
2 2316 1 199
2 2317 1 199
2 2318 1 199
2 2319 1 201
2 2320 1 201
2 2321 1 204
2 2322 1 204
2 2323 1 207
2 2324 1 207
2 2325 1 209
2 2326 1 209
2 2327 1 210
2 2328 1 210
2 2329 1 215
2 2330 1 215
2 2331 1 218
2 2332 1 218
2 2333 1 223
2 2334 1 223
2 2335 1 223
2 2336 1 225
2 2337 1 225
2 2338 1 228
2 2339 1 228
2 2340 1 231
2 2341 1 231
2 2342 1 233
2 2343 1 233
2 2344 1 234
2 2345 1 234
2 2346 1 239
2 2347 1 239
2 2348 1 242
2 2349 1 242
2 2350 1 247
2 2351 1 247
2 2352 1 247
2 2353 1 249
2 2354 1 249
2 2355 1 252
2 2356 1 252
2 2357 1 255
2 2358 1 255
2 2359 1 257
2 2360 1 257
2 2361 1 258
2 2362 1 258
2 2363 1 263
2 2364 1 263
2 2365 1 266
2 2366 1 266
2 2367 1 271
2 2368 1 271
2 2369 1 271
2 2370 1 273
2 2371 1 273
2 2372 1 276
2 2373 1 276
2 2374 1 279
2 2375 1 279
2 2376 1 281
2 2377 1 281
2 2378 1 282
2 2379 1 282
2 2380 1 287
2 2381 1 287
2 2382 1 290
2 2383 1 290
2 2384 1 295
2 2385 1 295
2 2386 1 295
2 2387 1 297
2 2388 1 297
2 2389 1 300
2 2390 1 300
2 2391 1 303
2 2392 1 303
2 2393 1 305
2 2394 1 305
2 2395 1 306
2 2396 1 306
2 2397 1 311
2 2398 1 311
2 2399 1 314
2 2400 1 314
2 2401 1 319
2 2402 1 319
2 2403 1 319
2 2404 1 321
2 2405 1 321
2 2406 1 324
2 2407 1 324
2 2408 1 327
2 2409 1 327
2 2410 1 329
2 2411 1 329
2 2412 1 330
2 2413 1 330
2 2414 1 335
2 2415 1 335
2 2416 1 338
2 2417 1 338
2 2418 1 343
2 2419 1 343
2 2420 1 343
2 2421 1 345
2 2422 1 345
2 2423 1 348
2 2424 1 348
2 2425 1 351
2 2426 1 351
2 2427 1 353
2 2428 1 353
2 2429 1 354
2 2430 1 354
2 2431 1 359
2 2432 1 359
2 2433 1 362
2 2434 1 362
2 2435 1 367
2 2436 1 367
2 2437 1 367
2 2438 1 369
2 2439 1 369
2 2440 1 372
2 2441 1 372
2 2442 1 375
2 2443 1 375
2 2444 1 377
2 2445 1 377
2 2446 1 378
2 2447 1 378
2 2448 1 383
2 2449 1 383
2 2450 1 386
2 2451 1 386
2 2452 1 391
2 2453 1 391
2 2454 1 391
2 2455 1 393
2 2456 1 393
2 2457 1 396
2 2458 1 396
2 2459 1 399
2 2460 1 399
2 2461 1 401
2 2462 1 401
2 2463 1 402
2 2464 1 402
2 2465 1 407
2 2466 1 407
2 2467 1 410
2 2468 1 410
2 2469 1 415
2 2470 1 415
2 2471 1 415
2 2472 1 417
2 2473 1 417
2 2474 1 420
2 2475 1 420
2 2476 1 423
2 2477 1 423
2 2478 1 425
2 2479 1 425
2 2480 1 426
2 2481 1 426
2 2482 1 431
2 2483 1 431
2 2484 1 434
2 2485 1 434
2 2486 1 439
2 2487 1 439
2 2488 1 439
2 2489 1 441
2 2490 1 441
2 2491 1 444
2 2492 1 444
2 2493 1 447
2 2494 1 447
2 2495 1 449
2 2496 1 449
2 2497 1 450
2 2498 1 450
2 2499 1 455
2 2500 1 455
2 2501 1 458
2 2502 1 458
2 2503 1 463
2 2504 1 463
2 2505 1 463
2 2506 1 465
2 2507 1 465
2 2508 1 468
2 2509 1 468
2 2510 1 471
2 2511 1 471
2 2512 1 473
2 2513 1 473
2 2514 1 474
2 2515 1 474
2 2516 1 479
2 2517 1 479
2 2518 1 482
2 2519 1 482
2 2520 1 487
2 2521 1 487
2 2522 1 487
2 2523 1 489
2 2524 1 489
2 2525 1 492
2 2526 1 492
2 2527 1 495
2 2528 1 495
2 2529 1 497
2 2530 1 497
2 2531 1 498
2 2532 1 498
2 2533 1 503
2 2534 1 503
2 2535 1 506
2 2536 1 506
2 2537 1 511
2 2538 1 511
2 2539 1 511
2 2540 1 513
2 2541 1 513
2 2542 1 516
2 2543 1 516
2 2544 1 519
2 2545 1 519
2 2546 1 521
2 2547 1 521
2 2548 1 522
2 2549 1 522
2 2550 1 527
2 2551 1 527
2 2552 1 530
2 2553 1 530
2 2554 1 535
2 2555 1 535
2 2556 1 535
2 2557 1 537
2 2558 1 537
2 2559 1 540
2 2560 1 540
2 2561 1 543
2 2562 1 543
2 2563 1 545
2 2564 1 545
2 2565 1 546
2 2566 1 546
2 2567 1 551
2 2568 1 551
2 2569 1 554
2 2570 1 554
2 2571 1 559
2 2572 1 559
2 2573 1 559
2 2574 1 561
2 2575 1 561
2 2576 1 564
2 2577 1 564
2 2578 1 567
2 2579 1 567
2 2580 1 569
2 2581 1 569
2 2582 1 570
2 2583 1 570
2 2584 1 575
2 2585 1 575
2 2586 1 578
2 2587 1 578
2 2588 1 583
2 2589 1 583
2 2590 1 583
2 2591 1 585
2 2592 1 585
2 2593 1 588
2 2594 1 588
2 2595 1 591
2 2596 1 591
2 2597 1 593
2 2598 1 593
2 2599 1 594
2 2600 1 594
2 2601 1 599
2 2602 1 599
2 2603 1 602
2 2604 1 602
2 2605 1 607
2 2606 1 607
2 2607 1 607
2 2608 1 609
2 2609 1 609
2 2610 1 612
2 2611 1 612
2 2612 1 615
2 2613 1 615
2 2614 1 617
2 2615 1 617
2 2616 1 618
2 2617 1 618
2 2618 1 623
2 2619 1 623
2 2620 1 626
2 2621 1 626
2 2622 1 631
2 2623 1 631
2 2624 1 631
2 2625 1 633
2 2626 1 633
2 2627 1 636
2 2628 1 636
2 2629 1 639
2 2630 1 639
2 2631 1 641
2 2632 1 641
2 2633 1 642
2 2634 1 642
2 2635 1 647
2 2636 1 647
2 2637 1 650
2 2638 1 650
2 2639 1 655
2 2640 1 655
2 2641 1 655
2 2642 1 657
2 2643 1 657
2 2644 1 660
2 2645 1 660
2 2646 1 663
2 2647 1 663
2 2648 1 665
2 2649 1 665
2 2650 1 666
2 2651 1 666
2 2652 1 671
2 2653 1 671
2 2654 1 674
2 2655 1 674
2 2656 1 679
2 2657 1 679
2 2658 1 679
2 2659 1 681
2 2660 1 681
2 2661 1 686
2 2662 1 686
2 2663 1 687
2 2664 1 687
2 2665 1 687
2 2666 1 689
2 2667 1 689
2 2668 1 694
2 2669 1 694
2 2670 1 697
2 2671 1 697
2 2672 1 702
2 2673 1 702
2 2674 1 708
2 2675 1 708
2 2676 1 711
2 2677 1 711
2 2678 1 713
2 2679 1 713
2 2680 1 722
2 2681 1 722
2 2682 1 728
2 2683 1 728
2 2684 1 730
2 2685 1 730
2 2686 1 732
2 2687 1 732
2 2688 1 733
2 2689 1 733
2 2690 1 734
2 2691 1 734
2 2692 1 736
2 2693 1 736
2 2694 1 739
2 2695 1 739
2 2696 1 742
2 2697 1 742
2 2698 1 745
2 2699 1 745
2 2700 1 746
2 2701 1 746
2 2702 1 748
2 2703 1 748
2 2704 1 750
2 2705 1 750
2 2706 1 756
2 2707 1 756
2 2708 1 759
2 2709 1 759
2 2710 1 759
2 2711 1 763
2 2712 1 763
2 2713 1 764
2 2714 1 764
2 2715 1 766
2 2716 1 766
2 2717 1 769
2 2718 1 769
2 2719 1 770
2 2720 1 770
2 2721 1 774
2 2722 1 774
2 2723 1 777
2 2724 1 777
2 2725 1 778
2 2726 1 778
2 2727 1 782
2 2728 1 782
2 2729 1 785
2 2730 1 785
2 2731 1 786
2 2732 1 786
2 2733 1 790
2 2734 1 790
2 2735 1 793
2 2736 1 793
2 2737 1 794
2 2738 1 794
2 2739 1 796
2 2740 1 796
2 2741 1 799
2 2742 1 799
2 2743 1 800
2 2744 1 800
2 2745 1 804
2 2746 1 804
2 2747 1 807
2 2748 1 807
2 2749 1 808
2 2750 1 808
2 2751 1 812
2 2752 1 812
2 2753 1 815
2 2754 1 815
2 2755 1 816
2 2756 1 816
2 2757 1 820
2 2758 1 820
2 2759 1 823
2 2760 1 823
2 2761 1 824
2 2762 1 824
2 2763 1 828
2 2764 1 828
2 2765 1 831
2 2766 1 831
2 2767 1 832
2 2768 1 832
2 2769 1 836
2 2770 1 836
2 2771 1 839
2 2772 1 839
2 2773 1 840
2 2774 1 840
2 2775 1 844
2 2776 1 844
2 2777 1 847
2 2778 1 847
2 2779 1 848
2 2780 1 848
2 2781 1 852
2 2782 1 852
2 2783 1 855
2 2784 1 855
2 2785 1 856
2 2786 1 856
2 2787 1 858
2 2788 1 858
2 2789 1 860
2 2790 1 860
2 2791 1 861
2 2792 1 861
2 2793 1 862
2 2794 1 862
2 2795 1 863
2 2796 1 863
2 2797 1 864
2 2798 1 864
2 2799 1 867
2 2800 1 867
2 2801 1 868
2 2802 1 868
2 2803 1 872
2 2804 1 872
2 2805 1 875
2 2806 1 875
2 2807 1 876
2 2808 1 876
2 2809 1 880
2 2810 1 880
2 2811 1 883
2 2812 1 883
2 2813 1 884
2 2814 1 884
2 2815 1 888
2 2816 1 888
2 2817 1 891
2 2818 1 891
2 2819 1 892
2 2820 1 892
2 2821 1 896
2 2822 1 896
2 2823 1 899
2 2824 1 899
2 2825 1 900
2 2826 1 900
2 2827 1 904
2 2828 1 904
2 2829 1 907
2 2830 1 907
2 2831 1 908
2 2832 1 908
2 2833 1 912
2 2834 1 912
2 2835 1 915
2 2836 1 915
2 2837 1 916
2 2838 1 916
2 2839 1 920
2 2840 1 920
2 2841 1 923
2 2842 1 923
2 2843 1 924
2 2844 1 924
2 2845 1 926
2 2846 1 926
2 2847 1 929
2 2848 1 929
2 2849 1 932
2 2850 1 932
2 2851 1 936
2 2852 1 936
2 2853 1 939
2 2854 1 939
2 2855 1 940
2 2856 1 940
2 2857 1 944
2 2858 1 944
2 2859 1 947
2 2860 1 947
2 2861 1 948
2 2862 1 948
2 2863 1 950
2 2864 1 950
2 2865 1 953
2 2866 1 953
2 2867 1 954
2 2868 1 954
2 2869 1 956
2 2870 1 956
2 2871 1 962
2 2872 1 962
2 2873 1 965
2 2874 1 965
2 2875 1 968
2 2876 1 968
2 2877 1 971
2 2878 1 971
2 2879 1 974
2 2880 1 974
2 2881 1 978
2 2882 1 978
2 2883 1 981
2 2884 1 981
2 2885 1 982
2 2886 1 982
2 2887 1 986
2 2888 1 986
2 2889 1 989
2 2890 1 989
2 2891 1 990
2 2892 1 990
2 2893 1 992
2 2894 1 992
2 2895 1 995
2 2896 1 995
2 2897 1 998
2 2898 1 998
2 2899 1 1002
2 2900 1 1002
2 2901 1 1005
2 2902 1 1005
2 2903 1 1006
2 2904 1 1006
2 2905 1 1010
2 2906 1 1010
2 2907 1 1013
2 2908 1 1013
2 2909 1 1014
2 2910 1 1014
2 2911 1 1018
2 2912 1 1018
2 2913 1 1021
2 2914 1 1021
2 2915 1 1022
2 2916 1 1022
2 2917 1 1026
2 2918 1 1026
2 2919 1 1029
2 2920 1 1029
2 2921 1 1030
2 2922 1 1030
2 2923 1 1034
2 2924 1 1034
2 2925 1 1037
2 2926 1 1037
2 2927 1 1038
2 2928 1 1038
2 2929 1 1040
2 2930 1 1040
2 2931 1 1043
2 2932 1 1043
2 2933 1 1044
2 2934 1 1044
2 2935 1 1048
2 2936 1 1048
2 2937 1 1051
2 2938 1 1051
2 2939 1 1052
2 2940 1 1052
2 2941 1 1054
2 2942 1 1054
2 2943 1 1056
2 2944 1 1056
2 2945 1 1059
2 2946 1 1059
2 2947 1 1060
2 2948 1 1060
2 2949 1 1062
2 2950 1 1062
2 2951 1 1064
2 2952 1 1064
2 2953 1 1066
2 2954 1 1066
2 2955 1 1068
2 2956 1 1068
2 2957 1 1069
2 2958 1 1069
2 2959 1 1070
2 2960 1 1070
2 2961 1 1071
2 2962 1 1071
2 2963 1 1072
2 2964 1 1072
2 2965 1 1073
2 2966 1 1073
2 2967 1 1074
2 2968 1 1074
2 2969 1 1075
2 2970 1 1075
2 2971 1 1077
2 2972 1 1077
2 2973 1 1080
2 2974 1 1080
2 2975 1 1084
2 2976 1 1084
2 2977 1 1087
2 2978 1 1087
2 2979 1 1090
2 2980 1 1090
2 2981 1 1094
2 2982 1 1094
2 2983 1 1097
2 2984 1 1097
2 2985 1 1098
2 2986 1 1098
2 2987 1 1101
2 2988 1 1101
2 2989 1 1102
2 2990 1 1102
2 2991 1 1106
2 2992 1 1106
2 2993 1 1109
2 2994 1 1109
2 2995 1 1110
2 2996 1 1110
2 2997 1 1114
2 2998 1 1114
2 2999 1 1117
2 3000 1 1117
2 3001 1 1118
2 3002 1 1118
2 3003 1 1122
2 3004 1 1122
2 3005 1 1125
2 3006 1 1125
2 3007 1 1128
2 3008 1 1128
2 3009 1 1132
2 3010 1 1132
2 3011 1 1135
2 3012 1 1135
2 3013 1 1138
2 3014 1 1138
2 3015 1 1142
2 3016 1 1142
2 3017 1 1145
2 3018 1 1145
2 3019 1 1146
2 3020 1 1146
2 3021 1 1148
2 3022 1 1148
2 3023 1 1151
2 3024 1 1151
2 3025 1 1152
2 3026 1 1152
2 3027 1 1156
2 3028 1 1156
2 3029 1 1159
2 3030 1 1159
2 3031 1 1160
2 3032 1 1160
2 3033 1 1164
2 3034 1 1164
2 3035 1 1167
2 3036 1 1167
2 3037 1 1168
2 3038 1 1168
2 3039 1 1172
2 3040 1 1172
2 3041 1 1175
2 3042 1 1175
2 3043 1 1176
2 3044 1 1176
2 3045 1 1180
2 3046 1 1180
2 3047 1 1183
2 3048 1 1183
2 3049 1 1184
2 3050 1 1184
2 3051 1 1188
2 3052 1 1188
2 3053 1 1191
2 3054 1 1191
2 3055 1 1192
2 3056 1 1192
2 3057 1 1194
2 3058 1 1194
2 3059 1 1200
2 3060 1 1200
2 3061 1 1203
2 3062 1 1203
2 3063 1 1206
2 3064 1 1206
2 3065 1 1209
2 3066 1 1209
2 3067 1 1212
2 3068 1 1212
2 3069 1 1216
2 3070 1 1216
2 3071 1 1219
2 3072 1 1219
2 3073 1 1220
2 3074 1 1220
2 3075 1 1224
2 3076 1 1224
2 3077 1 1227
2 3078 1 1227
2 3079 1 1228
2 3080 1 1228
2 3081 1 1232
2 3082 1 1232
2 3083 1 1235
2 3084 1 1235
2 3085 1 1236
2 3086 1 1236
2 3087 1 1240
2 3088 1 1240
2 3089 1 1243
2 3090 1 1243
2 3091 1 1244
2 3092 1 1244
2 3093 1 1248
2 3094 1 1248
2 3095 1 1251
2 3096 1 1251
2 3097 1 1252
2 3098 1 1252
2 3099 1 1256
2 3100 1 1256
2 3101 1 1259
2 3102 1 1259
2 3103 1 1260
2 3104 1 1260
2 3105 1 1264
2 3106 1 1264
2 3107 1 1267
2 3108 1 1267
2 3109 1 1268
2 3110 1 1268
2 3111 1 1270
2 3112 1 1270
2 3113 1 1273
2 3114 1 1273
2 3115 1 1276
2 3116 1 1276
2 3117 1 1280
2 3118 1 1280
2 3119 1 1283
2 3120 1 1283
2 3121 1 1284
2 3122 1 1284
2 3123 1 1288
2 3124 1 1288
2 3125 1 1291
2 3126 1 1291
2 3127 1 1292
2 3128 1 1292
2 3129 1 1296
2 3130 1 1296
2 3131 1 1299
2 3132 1 1299
2 3133 1 1300
2 3134 1 1300
2 3135 1 1304
2 3136 1 1304
2 3137 1 1307
2 3138 1 1307
2 3139 1 1308
2 3140 1 1308
2 3141 1 1314
2 3142 1 1314
2 3143 1 1317
2 3144 1 1317
2 3145 1 1318
2 3146 1 1318
2 3147 1 1322
2 3148 1 1322
2 3149 1 1325
2 3150 1 1325
2 3151 1 1326
2 3152 1 1326
2 3153 1 1330
2 3154 1 1330
2 3155 1 1333
2 3156 1 1333
2 3157 1 1334
2 3158 1 1334
2 3159 1 1338
2 3160 1 1338
2 3161 1 1341
2 3162 1 1341
2 3163 1 1342
2 3164 1 1342
2 3165 1 1344
2 3166 1 1344
2 3167 1 1347
2 3168 1 1347
2 3169 1 1350
2 3170 1 1350
2 3171 1 1354
2 3172 1 1354
2 3173 1 1357
2 3174 1 1357
2 3175 1 1358
2 3176 1 1358
2 3177 1 1362
2 3178 1 1362
2 3179 1 1365
2 3180 1 1365
2 3181 1 1368
2 3182 1 1368
2 3183 1 1370
2 3184 1 1370
2 3185 1 1372
2 3186 1 1372
2 3187 1 1374
2 3188 1 1374
2 3189 1 1376
2 3190 1 1376
2 3191 1 1378
2 3192 1 1378
2 3193 1 1380
2 3194 1 1380
2 3195 1 1381
2 3196 1 1381
2 3197 1 1382
2 3198 1 1382
2 3199 1 1382
2 3200 1 1385
2 3201 1 1385
2 3202 1 1388
2 3203 1 1388
2 3204 1 1396
2 3205 1 1396
2 3206 1 1399
2 3207 1 1399
2 3208 1 1400
2 3209 1 1400
2 3210 1 1404
2 3211 1 1404
2 3212 1 1407
2 3213 1 1407
2 3214 1 1410
2 3215 1 1410
2 3216 1 1412
2 3217 1 1412
2 3218 1 1414
2 3219 1 1414
2 3220 1 1416
2 3221 1 1416
2 3222 1 1417
2 3223 1 1417
2 3224 1 1419
2 3225 1 1419
2 3226 1 1420
2 3227 1 1420
2 3228 1 1424
2 3229 1 1424
2 3230 1 1427
2 3231 1 1427
2 3232 1 1428
2 3233 1 1428
2 3234 1 1432
2 3235 1 1432
2 3236 1 1435
2 3237 1 1435
2 3238 1 1436
2 3239 1 1436
2 3240 1 1440
2 3241 1 1440
2 3242 1 1443
2 3243 1 1443
2 3244 1 1444
2 3245 1 1444
2 3246 1 1448
2 3247 1 1448
2 3248 1 1451
2 3249 1 1451
2 3250 1 1452
2 3251 1 1452
2 3252 1 1456
2 3253 1 1456
2 3254 1 1459
2 3255 1 1459
2 3256 1 1460
2 3257 1 1460
2 3258 1 1464
2 3259 1 1464
2 3260 1 1467
2 3261 1 1467
2 3262 1 1468
2 3263 1 1468
2 3264 1 1472
2 3265 1 1472
2 3266 1 1475
2 3267 1 1475
2 3268 1 1476
2 3269 1 1476
2 3270 1 1480
2 3271 1 1480
2 3272 1 1483
2 3273 1 1483
2 3274 1 1484
2 3275 1 1484
2 3276 1 1488
2 3277 1 1488
2 3278 1 1491
2 3279 1 1491
2 3280 1 1492
2 3281 1 1492
2 3282 1 1496
2 3283 1 1496
2 3284 1 1499
2 3285 1 1499
2 3286 1 1500
2 3287 1 1500
2 3288 1 1504
2 3289 1 1504
2 3290 1 1507
2 3291 1 1507
2 3292 1 1508
2 3293 1 1508
2 3294 1 1512
2 3295 1 1512
2 3296 1 1515
2 3297 1 1515
2 3298 1 1516
2 3299 1 1516
2 3300 1 1518
2 3301 1 1518
2 3302 1 1519
2 3303 1 1519
2 3304 1 1522
2 3305 1 1522
2 3306 1 1525
2 3307 1 1525
2 3308 1 1525
2 3309 1 1526
2 3310 1 1526
2 3311 1 1527
2 3312 1 1527
2 3313 1 1528
2 3314 1 1528
2 3315 1 1531
2 3316 1 1531
2 3317 1 1534
2 3318 1 1534
2 3319 1 1534
2 3320 1 1534
2 3321 1 1536
2 3322 1 1536
2 3323 1 1536
2 3324 1 1536
2 3325 1 1539
2 3326 1 1539
2 3327 1 1542
2 3328 1 1542
2 3329 1 1542
2 3330 1 1542
2 3331 1 1542
2 3332 1 1544
2 3333 1 1544
2 3334 1 1547
2 3335 1 1547
2 3336 1 1550
2 3337 1 1550
2 3338 1 1550
2 3339 1 1550
2 3340 1 1550
2 3341 1 1551
2 3342 1 1551
2 3343 1 1551
2 3344 1 1553
2 3345 1 1553
2 3346 1 1553
2 3347 1 1553
2 3348 1 1556
2 3349 1 1556
2 3350 1 1559
2 3351 1 1559
2 3352 1 1559
2 3353 1 1561
2 3354 1 1561
2 3355 1 1561
2 3356 1 1561
2 3357 1 1564
2 3358 1 1564
2 3359 1 1567
2 3360 1 1567
2 3361 1 1567
2 3362 1 1569
2 3363 1 1569
2 3364 1 1569
2 3365 1 1572
2 3366 1 1572
2 3367 1 1574
2 3368 1 1574
2 3369 1 1574
2 3370 1 1575
2 3371 1 1575
2 3372 1 1575
2 3373 1 1575
2 3374 1 1576
2 3375 1 1576
2 3376 1 1576
2 3377 1 1577
2 3378 1 1577
2 3379 1 1577
2 3380 1 1580
2 3381 1 1580
2 3382 1 1583
2 3383 1 1583
2 3384 1 1583
2 3385 1 1583
2 3386 1 1584
2 3387 1 1584
2 3388 1 1585
2 3389 1 1585
2 3390 1 1585
2 3391 1 1585
2 3392 1 1588
2 3393 1 1588
2 3394 1 1591
2 3395 1 1591
2 3396 1 1591
2 3397 1 1591
2 3398 1 1592
2 3399 1 1592
2 3400 1 1593
2 3401 1 1593
2 3402 1 1593
2 3403 1 1596
2 3404 1 1596
2 3405 1 1598
2 3406 1 1598
2 3407 1 1599
2 3408 1 1599
2 3409 1 1599
2 3410 1 1599
2 3411 1 1599
2 3412 1 1601
2 3413 1 1601
2 3414 1 1601
2 3415 1 1601
2 3416 1 1604
2 3417 1 1604
2 3418 1 1607
2 3419 1 1607
2 3420 1 1607
2 3421 1 1609
2 3422 1 1609
2 3423 1 1609
2 3424 1 1609
2 3425 1 1612
2 3426 1 1612
2 3427 1 1615
2 3428 1 1615
2 3429 1 1615
2 3430 1 1617
2 3431 1 1617
2 3432 1 1617
2 3433 1 1617
2 3434 1 1620
2 3435 1 1620
2 3436 1 1623
2 3437 1 1623
2 3438 1 1626
2 3439 1 1626
2 3440 1 1630
2 3441 1 1630
2 3442 1 1633
2 3443 1 1633
2 3444 1 1638
2 3445 1 1638
2 3446 1 1640
2 3447 1 1640
2 3448 1 1644
2 3449 1 1644
2 3450 1 1646
2 3451 1 1646
2 3452 1 1646
2 3453 1 1650
2 3454 1 1650
2 3455 1 1651
2 3456 1 1651
2 3457 1 1654
2 3458 1 1654
2 3459 1 1657
2 3460 1 1657
2 3461 1 1662
2 3462 1 1662
2 3463 1 1664
2 3464 1 1664
2 3465 1 1665
2 3466 1 1665
2 3467 1 1667
2 3468 1 1667
2 3469 1 1671
2 3470 1 1671
2 3471 1 1672
2 3472 1 1672
2 3473 1 1675
2 3474 1 1675
2 3475 1 1677
2 3476 1 1677
2 3477 1 1681
2 3478 1 1681
2 3479 1 1686
2 3480 1 1686
2 3481 1 1688
2 3482 1 1688
2 3483 1 1688
2 3484 1 1688
2 3485 1 1693
2 3486 1 1693
2 3487 1 1694
2 3488 1 1694
2 3489 1 1695
2 3490 1 1695
2 3491 1 1698
2 3492 1 1698
2 3493 1 1698
2 3494 1 1702
2 3495 1 1702
2 3496 1 1703
2 3497 1 1703
2 3498 1 1706
2 3499 1 1706
2 3500 1 1707
2 3501 1 1707
2 3502 1 1710
2 3503 1 1710
2 3504 1 1714
2 3505 1 1714
2 3506 1 1717
2 3507 1 1717
2 3508 1 1720
2 3509 1 1720
2 3510 1 1726
2 3511 1 1726
2 3512 1 1727
2 3513 1 1727
2 3514 1 1730
2 3515 1 1730
2 3516 1 1731
2 3517 1 1731
2 3518 1 1732
2 3519 1 1732
2 3520 1 1734
2 3521 1 1734
2 3522 1 1737
2 3523 1 1737
2 3524 1 1740
2 3525 1 1740
2 3526 1 1746
2 3527 1 1746
2 3528 1 1747
2 3529 1 1747
2 3530 1 1756
2 3531 1 1756
2 3532 1 1756
2 3533 1 1757
2 3534 1 1757
2 3535 1 1764
2 3536 1 1764
2 3537 1 1764
2 3538 1 1765
2 3539 1 1765
2 3540 1 1780
2 3541 1 1780
2 3542 1 1788
2 3543 1 1788
2 3544 1 1791
2 3545 1 1791
2 3546 1 1791
2 3547 1 1792
2 3548 1 1792
2 3549 1 1795
2 3550 1 1795
2 3551 1 1795
2 3552 1 1796
2 3553 1 1796
2 3554 1 1800
2 3555 1 1800
2 3556 1 1828
2 3557 1 1828
2 3558 1 1830
2 3559 1 1830
2 3560 1 1837
2 3561 1 1837
2 3562 1 1838
2 3563 1 1838
2 3564 1 1901
2 3565 1 1901
0 33 5 1 1 1944
0 34 5 2 1 1953
0 35 5 2 1 1963
0 36 5 2 1 1974
0 37 5 2 1 1984
0 38 5 2 1 1995
0 39 5 2 1 2005
0 40 5 2 1 2015
0 41 5 2 1 2025
0 42 5 2 1 2035
0 43 5 2 1 2046
0 44 5 2 1 2056
0 45 5 2 1 2066
0 46 5 2 1 2076
0 47 5 2 1 2086
0 48 5 3 1 2096
0 49 5 3 1 2099
0 50 5 3 1 2102
0 51 5 3 1 2105
0 52 5 3 1 2108
0 53 5 3 1 2111
0 54 5 3 1 2114
0 55 5 3 1 2117
0 56 5 3 1 2120
0 57 5 3 1 2123
0 58 5 3 1 2126
0 59 5 3 1 2129
0 60 5 4 1 2132
0 61 5 3 1 2136
0 62 5 2 1 2139
0 63 5 2 1 2143
0 64 7 2 2 2215 2218
0 65 5 1 1 2222
0 66 7 3 2 2144 2223
0 67 5 1 1 2224
0 68 7 2 2 2216 2145
0 69 5 1 1 2227
0 70 7 1 2 65 2228
0 71 5 1 1 70
0 72 7 1 2 2137 2220
0 73 5 1 1 72
0 74 7 2 2 71 73
0 75 5 1 1 2229
0 76 7 2 2 2211 2230
0 77 5 1 1 2231
0 78 7 1 2 2140 69
0 79 7 1 2 77 78
0 80 5 1 1 79
0 81 7 2 2 67 80
0 82 5 1 1 2233
0 83 7 1 2 2212 82
0 84 5 2 1 83
0 85 7 1 2 2133 2234
0 86 5 1 1 85
0 87 7 2 2 2235 86
0 88 5 1 1 2237
0 89 7 2 2 2208 2238
0 90 5 2 1 2239
0 91 7 1 2 75 2236
0 92 5 1 1 91
0 93 7 1 2 2213 2225
0 94 5 1 1 93
0 95 7 2 2 92 94
0 96 5 1 1 2243
0 97 7 1 2 2241 96
0 98 5 2 1 97
0 99 7 1 2 2141 2232
0 100 5 1 1 99
0 101 7 1 2 2134 2226
0 102 5 1 1 101
0 103 7 2 2 100 102
0 104 5 2 1 2247
0 105 7 2 2 2245 2248
0 106 5 1 1 2251
0 107 7 1 2 2209 106
0 108 5 2 1 107
0 109 7 1 2 2130 2252
0 110 5 1 1 109
0 111 7 2 2 2253 110
0 112 5 1 1 2255
0 113 7 2 2 2205 2256
0 114 5 2 1 2257
0 115 7 1 2 88 2254
0 116 5 1 1 115
0 117 7 1 2 2240 2249
0 118 5 1 1 117
0 119 7 2 2 116 118
0 120 5 1 1 2261
0 121 7 1 2 2259 120
0 122 5 2 1 121
0 123 7 1 2 2242 2250
0 124 5 1 1 123
0 125 7 1 2 2244 124
0 126 5 1 1 125
0 127 7 3 2 2246 126
0 128 5 1 1 2265
0 129 7 2 2 2263 128
0 130 5 1 1 2268
0 131 7 1 2 2206 130
0 132 5 2 1 131
0 133 7 1 2 2127 2269
0 134 5 1 1 133
0 135 7 2 2 2270 134
0 136 5 1 1 2272
0 137 7 2 2 2202 2273
0 138 5 2 1 2274
0 139 7 1 2 112 2271
0 140 5 1 1 139
0 141 7 1 2 2258 2266
0 142 5 1 1 141
0 143 7 2 2 140 142
0 144 5 1 1 2278
0 145 7 1 2 2276 144
0 146 5 2 1 145
0 147 7 1 2 2260 2267
0 148 5 1 1 147
0 149 7 1 2 2262 148
0 150 5 1 1 149
0 151 7 3 2 2264 150
0 152 5 1 1 2282
0 153 7 2 2 2280 152
0 154 5 1 1 2285
0 155 7 1 2 2203 154
0 156 5 2 1 155
0 157 7 1 2 2124 2286
0 158 5 1 1 157
0 159 7 2 2 2287 158
0 160 5 1 1 2289
0 161 7 2 2 2199 2290
0 162 5 2 1 2291
0 163 7 1 2 136 2288
0 164 5 1 1 163
0 165 7 1 2 2275 2283
0 166 5 1 1 165
0 167 7 2 2 164 166
0 168 5 1 1 2295
0 169 7 1 2 2293 168
0 170 5 2 1 169
0 171 7 1 2 2277 2284
0 172 5 1 1 171
0 173 7 1 2 2279 172
0 174 5 1 1 173
0 175 7 3 2 2281 174
0 176 5 1 1 2299
0 177 7 2 2 2297 176
0 178 5 1 1 2302
0 179 7 1 2 2200 178
0 180 5 2 1 179
0 181 7 1 2 2121 2303
0 182 5 1 1 181
0 183 7 2 2 2304 182
0 184 5 1 1 2306
0 185 7 2 2 2196 2307
0 186 5 2 1 2308
0 187 7 1 2 160 2305
0 188 5 1 1 187
0 189 7 1 2 2292 2300
0 190 5 1 1 189
0 191 7 2 2 188 190
0 192 5 1 1 2312
0 193 7 1 2 2310 192
0 194 5 2 1 193
0 195 7 1 2 2294 2301
0 196 5 1 1 195
0 197 7 1 2 2296 196
0 198 5 1 1 197
0 199 7 3 2 2298 198
0 200 5 1 1 2316
0 201 7 2 2 2314 200
0 202 5 1 1 2319
0 203 7 1 2 2197 202
0 204 5 2 1 203
0 205 7 1 2 2118 2320
0 206 5 1 1 205
0 207 7 2 2 2321 206
0 208 5 1 1 2323
0 209 7 2 2 2193 2324
0 210 5 2 1 2325
0 211 7 1 2 184 2322
0 212 5 1 1 211
0 213 7 1 2 2309 2317
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 1 1 2329
0 217 7 1 2 2327 216
0 218 5 2 1 217
0 219 7 1 2 2311 2318
0 220 5 1 1 219
0 221 7 1 2 2313 220
0 222 5 1 1 221
0 223 7 3 2 2315 222
0 224 5 1 1 2333
0 225 7 2 2 2331 224
0 226 5 1 1 2336
0 227 7 1 2 2194 226
0 228 5 2 1 227
0 229 7 1 2 2115 2337
0 230 5 1 1 229
0 231 7 2 2 2338 230
0 232 5 1 1 2340
0 233 7 2 2 2190 2341
0 234 5 2 1 2342
0 235 7 1 2 208 2339
0 236 5 1 1 235
0 237 7 1 2 2326 2334
0 238 5 1 1 237
0 239 7 2 2 236 238
0 240 5 1 1 2346
0 241 7 1 2 2344 240
0 242 5 2 1 241
0 243 7 1 2 2328 2335
0 244 5 1 1 243
0 245 7 1 2 2330 244
0 246 5 1 1 245
0 247 7 3 2 2332 246
0 248 5 1 1 2350
0 249 7 2 2 2348 248
0 250 5 1 1 2353
0 251 7 1 2 2191 250
0 252 5 2 1 251
0 253 7 1 2 2112 2354
0 254 5 1 1 253
0 255 7 2 2 2355 254
0 256 5 1 1 2357
0 257 7 2 2 2187 2358
0 258 5 2 1 2359
0 259 7 1 2 232 2356
0 260 5 1 1 259
0 261 7 1 2 2343 2351
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 2363
0 265 7 1 2 2361 264
0 266 5 2 1 265
0 267 7 1 2 2345 2352
0 268 5 1 1 267
0 269 7 1 2 2347 268
0 270 5 1 1 269
0 271 7 3 2 2349 270
0 272 5 1 1 2367
0 273 7 2 2 2365 272
0 274 5 1 1 2370
0 275 7 1 2 2188 274
0 276 5 2 1 275
0 277 7 1 2 2109 2371
0 278 5 1 1 277
0 279 7 2 2 2372 278
0 280 5 1 1 2374
0 281 7 2 2 2184 2375
0 282 5 2 1 2376
0 283 7 1 2 256 2373
0 284 5 1 1 283
0 285 7 1 2 2360 2368
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 2380
0 289 7 1 2 2378 288
0 290 5 2 1 289
0 291 7 1 2 2362 2369
0 292 5 1 1 291
0 293 7 1 2 2364 292
0 294 5 1 1 293
0 295 7 3 2 2366 294
0 296 5 1 1 2384
0 297 7 2 2 2382 296
0 298 5 1 1 2387
0 299 7 1 2 2185 298
0 300 5 2 1 299
0 301 7 1 2 2106 2388
0 302 5 1 1 301
0 303 7 2 2 2389 302
0 304 5 1 1 2391
0 305 7 2 2 2181 2392
0 306 5 2 1 2393
0 307 7 1 2 280 2390
0 308 5 1 1 307
0 309 7 1 2 2377 2385
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 2397
0 313 7 1 2 2395 312
0 314 5 2 1 313
0 315 7 1 2 2379 2386
0 316 5 1 1 315
0 317 7 1 2 2381 316
0 318 5 1 1 317
0 319 7 3 2 2383 318
0 320 5 1 1 2401
0 321 7 2 2 2399 320
0 322 5 1 1 2404
0 323 7 1 2 2182 322
0 324 5 2 1 323
0 325 7 1 2 2103 2405
0 326 5 1 1 325
0 327 7 2 2 2406 326
0 328 5 1 1 2408
0 329 7 2 2 2178 2409
0 330 5 2 1 2410
0 331 7 1 2 304 2407
0 332 5 1 1 331
0 333 7 1 2 2394 2402
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 2414
0 337 7 1 2 2412 336
0 338 5 2 1 337
0 339 7 1 2 2396 2403
0 340 5 1 1 339
0 341 7 1 2 2398 340
0 342 5 1 1 341
0 343 7 3 2 2400 342
0 344 5 1 1 2418
0 345 7 2 2 2416 344
0 346 5 1 1 2421
0 347 7 1 2 2179 346
0 348 5 2 1 347
0 349 7 1 2 2100 2422
0 350 5 1 1 349
0 351 7 2 2 2423 350
0 352 5 1 1 2425
0 353 7 2 2 2175 2426
0 354 5 2 1 2427
0 355 7 1 2 328 2424
0 356 5 1 1 355
0 357 7 1 2 2411 2419
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 2431
0 361 7 1 2 2429 360
0 362 5 2 1 361
0 363 7 1 2 2413 2420
0 364 5 1 1 363
0 365 7 1 2 2415 364
0 366 5 1 1 365
0 367 7 3 2 2417 366
0 368 5 1 1 2435
0 369 7 2 2 2433 368
0 370 5 1 1 2438
0 371 7 1 2 2176 370
0 372 5 2 1 371
0 373 7 1 2 2097 2439
0 374 5 1 1 373
0 375 7 2 2 2440 374
0 376 5 1 1 2442
0 377 7 2 2 2173 2443
0 378 5 2 1 2444
0 379 7 1 2 352 2441
0 380 5 1 1 379
0 381 7 1 2 2428 2436
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 2448
0 385 7 1 2 2446 384
0 386 5 2 1 385
0 387 7 1 2 2430 2437
0 388 5 1 1 387
0 389 7 1 2 2432 388
0 390 5 1 1 389
0 391 7 3 2 2434 390
0 392 5 1 1 2452
0 393 7 2 2 2450 392
0 394 5 1 1 2455
0 395 7 1 2 2174 394
0 396 5 2 1 395
0 397 7 1 2 2087 2456
0 398 5 1 1 397
0 399 7 2 2 2457 398
0 400 5 1 1 2459
0 401 7 2 2 2171 2460
0 402 5 2 1 2461
0 403 7 1 2 376 2458
0 404 5 1 1 403
0 405 7 1 2 2445 2453
0 406 5 1 1 405
0 407 7 2 2 404 406
0 408 5 1 1 2465
0 409 7 1 2 2463 408
0 410 5 2 1 409
0 411 7 1 2 2447 2454
0 412 5 1 1 411
0 413 7 1 2 2449 412
0 414 5 1 1 413
0 415 7 3 2 2451 414
0 416 5 1 1 2469
0 417 7 2 2 2467 416
0 418 5 1 1 2472
0 419 7 1 2 2172 418
0 420 5 2 1 419
0 421 7 1 2 2077 2473
0 422 5 1 1 421
0 423 7 2 2 2474 422
0 424 5 1 1 2476
0 425 7 2 2 2169 2477
0 426 5 2 1 2478
0 427 7 1 2 400 2475
0 428 5 1 1 427
0 429 7 1 2 2462 2470
0 430 5 1 1 429
0 431 7 2 2 428 430
0 432 5 1 1 2482
0 433 7 1 2 2480 432
0 434 5 2 1 433
0 435 7 1 2 2464 2471
0 436 5 1 1 435
0 437 7 1 2 2466 436
0 438 5 1 1 437
0 439 7 3 2 2468 438
0 440 5 1 1 2486
0 441 7 2 2 2484 440
0 442 5 1 1 2489
0 443 7 1 2 2170 442
0 444 5 2 1 443
0 445 7 1 2 2067 2490
0 446 5 1 1 445
0 447 7 2 2 2491 446
0 448 5 1 1 2493
0 449 7 2 2 2167 2494
0 450 5 2 1 2495
0 451 7 1 2 424 2492
0 452 5 1 1 451
0 453 7 1 2 2479 2487
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 2499
0 457 7 1 2 2497 456
0 458 5 2 1 457
0 459 7 1 2 2481 2488
0 460 5 1 1 459
0 461 7 1 2 2483 460
0 462 5 1 1 461
0 463 7 3 2 2485 462
0 464 5 1 1 2503
0 465 7 2 2 2501 464
0 466 5 1 1 2506
0 467 7 1 2 2168 466
0 468 5 2 1 467
0 469 7 1 2 2057 2507
0 470 5 1 1 469
0 471 7 2 2 2508 470
0 472 5 1 1 2510
0 473 7 2 2 2165 2511
0 474 5 2 1 2512
0 475 7 1 2 448 2509
0 476 5 1 1 475
0 477 7 1 2 2496 2504
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 2516
0 481 7 1 2 2514 480
0 482 5 2 1 481
0 483 7 1 2 2498 2505
0 484 5 1 1 483
0 485 7 1 2 2500 484
0 486 5 1 1 485
0 487 7 3 2 2502 486
0 488 5 1 1 2520
0 489 7 2 2 2518 488
0 490 5 1 1 2523
0 491 7 1 2 2166 490
0 492 5 2 1 491
0 493 7 1 2 2047 2524
0 494 5 1 1 493
0 495 7 2 2 2525 494
0 496 5 1 1 2527
0 497 7 2 2 2163 2528
0 498 5 2 1 2529
0 499 7 1 2 472 2526
0 500 5 1 1 499
0 501 7 1 2 2513 2521
0 502 5 1 1 501
0 503 7 2 2 500 502
0 504 5 1 1 2533
0 505 7 1 2 2531 504
0 506 5 2 1 505
0 507 7 1 2 2515 2522
0 508 5 1 1 507
0 509 7 1 2 2517 508
0 510 5 1 1 509
0 511 7 3 2 2519 510
0 512 5 1 1 2537
0 513 7 2 2 2535 512
0 514 5 1 1 2540
0 515 7 1 2 2164 514
0 516 5 2 1 515
0 517 7 1 2 2036 2541
0 518 5 1 1 517
0 519 7 2 2 2542 518
0 520 5 1 1 2544
0 521 7 2 2 2161 2545
0 522 5 2 1 2546
0 523 7 1 2 496 2543
0 524 5 1 1 523
0 525 7 1 2 2530 2538
0 526 5 1 1 525
0 527 7 2 2 524 526
0 528 5 1 1 2550
0 529 7 1 2 2548 528
0 530 5 2 1 529
0 531 7 1 2 2532 2539
0 532 5 1 1 531
0 533 7 1 2 2534 532
0 534 5 1 1 533
0 535 7 3 2 2536 534
0 536 5 1 1 2554
0 537 7 2 2 2552 536
0 538 5 1 1 2557
0 539 7 1 2 2162 538
0 540 5 2 1 539
0 541 7 1 2 2026 2558
0 542 5 1 1 541
0 543 7 2 2 2559 542
0 544 5 1 1 2561
0 545 7 2 2 2159 2562
0 546 5 2 1 2563
0 547 7 1 2 520 2560
0 548 5 1 1 547
0 549 7 1 2 2547 2555
0 550 5 1 1 549
0 551 7 2 2 548 550
0 552 5 1 1 2567
0 553 7 1 2 2565 552
0 554 5 2 1 553
0 555 7 1 2 2549 2556
0 556 5 1 1 555
0 557 7 1 2 2551 556
0 558 5 1 1 557
0 559 7 3 2 2553 558
0 560 5 1 1 2571
0 561 7 2 2 2569 560
0 562 5 1 1 2574
0 563 7 1 2 2160 562
0 564 5 2 1 563
0 565 7 1 2 2016 2575
0 566 5 1 1 565
0 567 7 2 2 2576 566
0 568 5 1 1 2578
0 569 7 2 2 2157 2579
0 570 5 2 1 2580
0 571 7 1 2 544 2577
0 572 5 1 1 571
0 573 7 1 2 2564 2572
0 574 5 1 1 573
0 575 7 2 2 572 574
0 576 5 1 1 2584
0 577 7 1 2 2582 576
0 578 5 2 1 577
0 579 7 1 2 2566 2573
0 580 5 1 1 579
0 581 7 1 2 2568 580
0 582 5 1 1 581
0 583 7 3 2 2570 582
0 584 5 1 1 2588
0 585 7 2 2 2586 584
0 586 5 1 1 2591
0 587 7 1 2 2158 586
0 588 5 2 1 587
0 589 7 1 2 2006 2592
0 590 5 1 1 589
0 591 7 2 2 2593 590
0 592 5 1 1 2595
0 593 7 2 2 2155 2596
0 594 5 2 1 2597
0 595 7 1 2 568 2594
0 596 5 1 1 595
0 597 7 1 2 2581 2589
0 598 5 1 1 597
0 599 7 2 2 596 598
0 600 5 1 1 2601
0 601 7 1 2 2599 600
0 602 5 2 1 601
0 603 7 1 2 2583 2590
0 604 5 1 1 603
0 605 7 1 2 2585 604
0 606 5 1 1 605
0 607 7 3 2 2587 606
0 608 5 1 1 2605
0 609 7 2 2 2603 608
0 610 5 1 1 2608
0 611 7 1 2 2156 610
0 612 5 2 1 611
0 613 7 1 2 1996 2609
0 614 5 1 1 613
0 615 7 2 2 2610 614
0 616 5 1 1 2612
0 617 7 2 2 2153 2613
0 618 5 2 1 2614
0 619 7 1 2 592 2611
0 620 5 1 1 619
0 621 7 1 2 2598 2606
0 622 5 1 1 621
0 623 7 2 2 620 622
0 624 5 1 1 2618
0 625 7 1 2 2616 624
0 626 5 2 1 625
0 627 7 1 2 2600 2607
0 628 5 1 1 627
0 629 7 1 2 2602 628
0 630 5 1 1 629
0 631 7 3 2 2604 630
0 632 5 1 1 2622
0 633 7 2 2 2620 632
0 634 5 1 1 2625
0 635 7 1 2 2154 634
0 636 5 2 1 635
0 637 7 1 2 1985 2626
0 638 5 1 1 637
0 639 7 2 2 2627 638
0 640 5 1 1 2629
0 641 7 2 2 2151 2630
0 642 5 2 1 2631
0 643 7 1 2 616 2628
0 644 5 1 1 643
0 645 7 1 2 2615 2623
0 646 5 1 1 645
0 647 7 2 2 644 646
0 648 5 1 1 2635
0 649 7 1 2 2633 648
0 650 5 2 1 649
0 651 7 1 2 2617 2624
0 652 5 1 1 651
0 653 7 1 2 2619 652
0 654 5 1 1 653
0 655 7 3 2 2621 654
0 656 5 1 1 2639
0 657 7 2 2 2637 656
0 658 5 1 1 2642
0 659 7 1 2 2152 658
0 660 5 2 1 659
0 661 7 1 2 1975 2643
0 662 5 1 1 661
0 663 7 2 2 2644 662
0 664 5 1 1 2646
0 665 7 2 2 2149 2647
0 666 5 2 1 2648
0 667 7 1 2 640 2645
0 668 5 1 1 667
0 669 7 1 2 2632 2640
0 670 5 1 1 669
0 671 7 2 2 668 670
0 672 5 1 1 2652
0 673 7 1 2 2650 672
0 674 5 2 1 673
0 675 7 1 2 2634 2641
0 676 5 1 1 675
0 677 7 1 2 2636 676
0 678 5 1 1 677
0 679 7 3 2 2638 678
0 680 5 1 1 2656
0 681 7 2 2 2654 680
0 682 5 1 1 2659
0 683 7 1 2 1964 2660
0 684 5 1 1 683
0 685 7 1 2 2150 682
0 686 5 2 1 685
0 687 7 3 2 684 2661
0 688 7 1 2 2147 2663
0 689 5 2 1 688
0 690 7 1 2 664 2662
0 691 5 1 1 690
0 692 7 1 2 2649 2657
0 693 5 1 1 692
0 694 7 2 2 691 693
0 695 5 1 1 2668
0 696 7 1 2 2666 695
0 697 5 2 1 696
0 698 7 1 2 2651 2658
0 699 5 1 1 698
0 700 7 1 2 2653 699
0 701 5 1 1 700
0 702 7 2 2 2655 701
0 703 5 1 1 2672
0 704 7 1 2 2667 2673
0 705 5 1 1 704
0 706 7 1 2 2669 705
0 707 5 1 1 706
0 708 7 2 2 2670 707
0 709 7 1 2 2664 2674
0 710 5 1 1 709
0 711 7 2 2 2671 703
0 712 5 1 1 2676
0 713 7 2 2 2148 712
0 714 5 1 1 2678
0 715 7 1 2 2675 2679
0 716 5 1 1 715
0 717 7 1 2 1954 2677
0 718 5 1 1 717
0 719 7 1 2 33 714
0 720 7 1 2 718 719
0 721 5 1 1 720
0 722 7 2 2 716 721
0 723 5 1 1 2680
0 724 7 1 2 710 2681
0 725 5 1 1 724
0 726 7 1 2 2665 723
0 727 5 1 1 726
0 728 7 2 2 725 727
0 729 5 1 1 2682
0 730 7 2 2 2007 2088
0 731 5 1 1 2684
0 732 7 2 2 1997 2078
0 733 5 2 1 2686
0 734 7 2 2 2008 2068
0 735 5 1 1 2690
0 736 7 2 2 1986 2089
0 737 5 1 1 2692
0 738 7 1 2 2691 2693
0 739 5 2 1 738
0 740 7 1 2 735 737
0 741 5 1 1 740
0 742 7 2 2 741 2694
0 743 5 1 1 2696
0 744 7 1 2 2687 2697
0 745 5 2 1 744
0 746 7 2 2 2695 2698
0 747 5 1 1 2700
0 748 7 2 2 1998 2090
0 749 5 1 1 2702
0 750 7 2 2 2009 2079
0 751 5 1 1 2704
0 752 7 1 2 749 2705
0 753 5 1 1 752
0 754 7 1 2 2703 751
0 755 5 1 1 754
0 756 7 2 2 753 755
0 757 5 1 1 2706
0 758 7 1 2 747 757
0 759 5 3 1 758
0 760 7 1 2 2688 2708
0 761 5 1 1 760
0 762 7 1 2 2685 761
0 763 5 2 1 762
0 764 7 2 2 1976 2091
0 765 5 1 1 2713
0 766 7 2 2 2010 2058
0 767 5 1 1 2715
0 768 7 1 2 2714 2716
0 769 5 2 1 768
0 770 7 2 2 1999 2069
0 771 5 1 1 2719
0 772 7 1 2 765 767
0 773 5 1 1 772
0 774 7 2 2 2717 773
0 775 5 1 1 2721
0 776 7 1 2 2720 2722
0 777 5 2 1 776
0 778 7 2 2 2718 2723
0 779 5 1 1 2725
0 780 7 1 2 2689 743
0 781 5 1 1 780
0 782 7 2 2 2699 781
0 783 5 1 1 2727
0 784 7 1 2 779 2728
0 785 5 2 1 784
0 786 7 2 2 1987 2080
0 787 5 1 1 2731
0 788 7 1 2 771 775
0 789 5 1 1 788
0 790 7 2 2 2724 789
0 791 5 1 1 2733
0 792 7 1 2 2732 2734
0 793 5 2 1 792
0 794 7 2 2 1965 2092
0 795 5 1 1 2737
0 796 7 2 2 2011 2048
0 797 5 1 1 2739
0 798 7 1 2 2738 2740
0 799 5 2 1 798
0 800 7 2 2 2000 2059
0 801 5 1 1 2743
0 802 7 1 2 795 797
0 803 5 1 1 802
0 804 7 2 2 2741 803
0 805 5 1 1 2745
0 806 7 1 2 2744 2746
0 807 5 2 1 806
0 808 7 2 2 2742 2747
0 809 5 1 1 2749
0 810 7 1 2 787 791
0 811 5 1 1 810
0 812 7 2 2 2735 811
0 813 5 1 1 2751
0 814 7 1 2 809 2752
0 815 5 2 1 814
0 816 7 2 2 2736 2753
0 817 5 1 1 2755
0 818 7 1 2 2726 783
0 819 5 1 1 818
0 820 7 2 2 2729 819
0 821 5 1 1 2757
0 822 7 1 2 817 2758
0 823 5 2 1 822
0 824 7 2 2 2730 2759
0 825 5 1 1 2761
0 826 7 1 2 2701 2707
0 827 5 1 1 826
0 828 7 2 2 2709 827
0 829 5 1 1 2763
0 830 7 1 2 825 2764
0 831 5 2 1 830
0 832 7 2 2 1977 2081
0 833 5 1 1 2767
0 834 7 1 2 801 805
0 835 5 1 1 834
0 836 7 2 2 2748 835
0 837 5 1 1 2769
0 838 7 1 2 2768 2770
0 839 5 2 1 838
0 840 7 2 2 1988 2070
0 841 5 1 1 2773
0 842 7 1 2 833 837
0 843 5 1 1 842
0 844 7 2 2 2771 843
0 845 5 1 1 2775
0 846 7 1 2 2774 2776
0 847 5 2 1 846
0 848 7 2 2 2772 2777
0 849 5 1 1 2779
0 850 7 1 2 2750 813
0 851 5 1 1 850
0 852 7 2 2 2754 851
0 853 5 1 1 2781
0 854 7 1 2 849 2782
0 855 5 2 1 854
0 856 7 2 2 2012 2017
0 857 5 1 1 2785
0 858 7 2 2 2001 2027
0 859 5 1 1 2787
0 860 7 2 2 2786 2788
0 861 5 2 1 2789
0 862 7 2 2 2037 2790
0 863 5 2 1 2793
0 864 7 2 2 1955 2093
0 865 5 1 1 2797
0 866 7 1 2 2794 2798
0 867 5 2 1 866
0 868 7 2 2 2013 2038
0 869 5 1 1 2801
0 870 7 1 2 2795 865
0 871 5 1 1 870
0 872 7 2 2 2799 871
0 873 5 1 1 2803
0 874 7 1 2 2802 2804
0 875 5 2 1 874
0 876 7 2 2 2800 2805
0 877 5 1 1 2807
0 878 7 1 2 841 845
0 879 5 1 1 878
0 880 7 2 2 2778 879
0 881 5 1 1 2809
0 882 7 1 2 877 2810
0 883 5 2 1 882
0 884 7 2 2 1989 2060
0 885 5 1 1 2813
0 886 7 1 2 869 873
0 887 5 1 1 886
0 888 7 2 2 2806 887
0 889 5 1 1 2815
0 890 7 1 2 2814 2816
0 891 5 2 1 890
0 892 7 2 2 2002 2049
0 893 5 1 1 2819
0 894 7 1 2 885 889
0 895 5 1 1 894
0 896 7 2 2 2817 895
0 897 5 1 1 2821
0 898 7 1 2 2820 2822
0 899 5 2 1 898
0 900 7 2 2 2818 2823
0 901 5 1 1 2825
0 902 7 1 2 2808 881
0 903 5 1 1 902
0 904 7 2 2 2811 903
0 905 5 1 1 2827
0 906 7 1 2 901 2828
0 907 5 2 1 906
0 908 7 2 2 2812 2829
0 909 5 1 1 2831
0 910 7 1 2 2780 853
0 911 5 1 1 910
0 912 7 2 2 2783 911
0 913 5 1 1 2833
0 914 7 1 2 909 2834
0 915 5 2 1 914
0 916 7 2 2 2784 2835
0 917 5 1 1 2837
0 918 7 1 2 2756 821
0 919 5 1 1 918
0 920 7 2 2 2760 919
0 921 5 1 1 2839
0 922 7 1 2 917 2840
0 923 5 2 1 922
0 924 7 2 2 1966 2082
0 925 5 1 1 2843
0 926 7 2 2 1978 2071
0 927 5 1 1 2845
0 928 7 1 2 2844 2846
0 929 5 2 1 928
0 930 7 1 2 893 897
0 931 5 1 1 930
0 932 7 2 2 2824 931
0 933 5 1 1 2849
0 934 7 1 2 925 927
0 935 5 1 1 934
0 936 7 2 2 2847 935
0 937 5 1 1 2851
0 938 7 1 2 2850 2852
0 939 5 2 1 938
0 940 7 2 2 2848 2853
0 941 5 1 1 2855
0 942 7 1 2 2826 905
0 943 5 1 1 942
0 944 7 2 2 2830 943
0 945 5 1 1 2857
0 946 7 1 2 941 2858
0 947 5 2 1 946
0 948 7 2 2 1990 2050
0 949 5 1 1 2861
0 950 7 2 2 1956 2083
0 951 5 1 1 2863
0 952 7 1 2 2862 2864
0 953 5 2 1 952
0 954 7 2 2 1945 2094
0 955 5 1 1 2867
0 956 7 2 2 1979 2061
0 957 5 1 1 2869
0 958 7 1 2 2003 2039
0 959 5 1 1 958
0 960 7 1 2 2791 959
0 961 5 1 1 960
0 962 7 2 2 2796 961
0 963 5 1 1 2871
0 964 7 1 2 2870 2872
0 965 5 2 1 964
0 966 7 1 2 957 963
0 967 5 1 1 966
0 968 7 2 2 2873 967
0 969 5 1 1 2875
0 970 7 1 2 2868 2876
0 971 5 2 1 970
0 972 7 1 2 955 969
0 973 5 1 1 972
0 974 7 2 2 2877 973
0 975 5 1 1 2879
0 976 7 1 2 949 951
0 977 5 1 1 976
0 978 7 2 2 2865 977
0 979 5 1 1 2881
0 980 7 1 2 2880 2882
0 981 5 2 1 980
0 982 7 2 2 2866 2883
0 983 5 1 1 2885
0 984 7 1 2 933 937
0 985 5 1 1 984
0 986 7 2 2 2854 985
0 987 5 1 1 2887
0 988 7 1 2 983 2888
0 989 5 2 1 988
0 990 7 2 2 2014 2028
0 991 5 1 1 2891
0 992 7 2 2 1967 2072
0 993 5 1 1 2893
0 994 7 1 2 2892 2894
0 995 5 2 1 994
0 996 7 1 2 975 979
0 997 5 1 1 996
0 998 7 2 2 2884 997
0 999 5 1 1 2897
0 1000 7 1 2 991 993
0 1001 5 1 1 1000
0 1002 7 2 2 2895 1001
0 1003 5 1 1 2899
0 1004 7 1 2 2898 2900
0 1005 5 2 1 1004
0 1006 7 2 2 2896 2901
0 1007 5 1 1 2903
0 1008 7 1 2 2886 987
0 1009 5 1 1 1008
0 1010 7 2 2 2889 1009
0 1011 5 1 1 2905
0 1012 7 1 2 1007 2906
0 1013 5 2 1 1012
0 1014 7 2 2 2890 2907
0 1015 5 1 1 2909
0 1016 7 1 2 2856 945
0 1017 5 1 1 1016
0 1018 7 2 2 2859 1017
0 1019 5 1 1 2911
0 1020 7 1 2 1015 2912
0 1021 5 2 1 1020
0 1022 7 2 2 2860 2913
0 1023 5 1 1 2915
0 1024 7 1 2 2832 913
0 1025 5 1 1 1024
0 1026 7 2 2 2836 1025
0 1027 5 1 1 2917
0 1028 7 1 2 1023 2918
0 1029 5 2 1 1028
0 1030 7 2 2 2874 2878
0 1031 5 1 1 2921
0 1032 7 1 2 2904 1011
0 1033 5 1 1 1032
0 1034 7 2 2 2908 1033
0 1035 5 1 1 2923
0 1036 7 1 2 1031 2924
0 1037 5 2 1 1036
0 1038 7 2 2 1991 2040
0 1039 5 1 1 2927
0 1040 7 2 2 1980 2051
0 1041 5 1 1 2929
0 1042 7 1 2 2928 2930
0 1043 5 2 1 1042
0 1044 7 2 2 1946 2084
0 1045 5 1 1 2933
0 1046 7 1 2 1039 1041
0 1047 5 1 1 1046
0 1048 7 2 2 2931 1047
0 1049 5 1 1 2935
0 1050 7 1 2 2934 2936
0 1051 5 2 1 1050
0 1052 7 2 2 2932 2937
0 1053 5 1 1 2939
0 1054 7 2 2 1957 2073
0 1055 5 1 1 2941
0 1056 7 2 2 32 2095
0 1057 5 1 1 2943
0 1058 7 1 2 2942 2944
0 1059 5 2 1 1058
0 1060 7 2 2 1968 2062
0 1061 5 1 1 2947
0 1062 7 2 2 1981 2029
0 1063 5 1 1 2949
0 1064 7 2 2 1937 2052
0 1065 5 1 1 2951
0 1066 7 2 2 1958 2030
0 1067 5 1 1 2953
0 1068 7 2 2 2952 2954
0 1069 5 2 1 2955
0 1070 7 2 2 1969 2956
0 1071 5 2 1 2959
0 1072 7 2 2 2950 2960
0 1073 5 2 1 2963
0 1074 7 2 2 1992 2964
0 1075 5 2 1 2967
0 1076 7 1 2 2948 2968
0 1077 5 2 1 1076
0 1078 7 1 2 1061 2969
0 1079 5 1 1 1078
0 1080 7 2 2 2971 1079
0 1081 5 1 1 2973
0 1082 7 1 2 857 859
0 1083 5 1 1 1082
0 1084 7 2 2 2792 1083
0 1085 5 1 1 2975
0 1086 7 1 2 2974 2976
0 1087 5 2 1 1086
0 1088 7 1 2 1081 1085
0 1089 5 1 1 1088
0 1090 7 2 2 2977 1089
0 1091 5 1 1 2979
0 1092 7 1 2 1055 1057
0 1093 5 1 1 1092
0 1094 7 2 2 2945 1093
0 1095 5 1 1 2981
0 1096 7 1 2 2980 2982
0 1097 5 2 1 1096
0 1098 7 2 2 2946 2983
0 1099 5 1 1 2985
0 1100 7 1 2 1053 1099
0 1101 5 2 1 1100
0 1102 7 2 2 2972 2978
0 1103 5 1 1 2989
0 1104 7 1 2 2940 2986
0 1105 5 1 1 1104
0 1106 7 2 2 2987 1105
0 1107 5 1 1 2991
0 1108 7 1 2 1103 2992
0 1109 5 2 1 1108
0 1110 7 2 2 2988 2993
0 1111 5 1 1 2995
0 1112 7 1 2 2922 1035
0 1113 5 1 1 1112
0 1114 7 2 2 2925 1113
0 1115 5 1 1 2997
0 1116 7 1 2 1111 2998
0 1117 5 2 1 1116
0 1118 7 2 2 2926 2999
0 1119 5 1 1 3001
0 1120 7 1 2 2910 1019
0 1121 5 1 1 1120
0 1122 7 2 2 2914 1121
0 1123 5 1 1 3003
0 1124 7 1 2 1119 3004
0 1125 5 2 1 1124
0 1126 7 1 2 999 1003
0 1127 5 1 1 1126
0 1128 7 2 2 2902 1127
0 1129 5 1 1 3007
0 1130 7 1 2 2990 1107
0 1131 5 1 1 1130
0 1132 7 2 2 2994 1131
0 1133 5 1 1 3009
0 1134 7 1 2 3008 3010
0 1135 5 2 1 1134
0 1136 7 1 2 1045 1049
0 1137 5 1 1 1136
0 1138 7 2 2 2938 1137
0 1139 5 1 1 3013
0 1140 7 1 2 1091 1095
0 1141 5 1 1 1140
0 1142 7 2 2 2984 1141
0 1143 5 1 1 3015
0 1144 7 1 2 3014 3016
0 1145 5 2 1 1144
0 1146 7 2 2 1970 2053
0 1147 5 1 1 3019
0 1148 7 2 2 1959 2063
0 1149 5 1 1 3021
0 1150 7 1 2 3020 3022
0 1151 5 2 1 1150
0 1152 7 2 2 1947 2074
0 1153 5 1 1 3025
0 1154 7 1 2 1147 1149
0 1155 5 1 1 1154
0 1156 7 2 2 3023 1155
0 1157 5 1 1 3027
0 1158 7 1 2 3026 3028
0 1159 5 2 1 1158
0 1160 7 2 2 3024 3029
0 1161 5 1 1 3031
0 1162 7 1 2 1139 1143
0 1163 5 1 1 1162
0 1164 7 2 2 3017 1163
0 1165 5 1 1 3033
0 1166 7 1 2 1161 3034
0 1167 5 2 1 1166
0 1168 7 2 2 3018 3035
0 1169 5 1 1 3037
0 1170 7 1 2 1129 1133
0 1171 5 1 1 1170
0 1172 7 2 2 3011 1171
0 1173 5 1 1 3039
0 1174 7 1 2 1169 3040
0 1175 5 2 1 1174
0 1176 7 2 2 3012 3041
0 1177 5 1 1 3043
0 1178 7 1 2 2996 1115
0 1179 5 1 1 1178
0 1180 7 2 2 3000 1179
0 1181 5 1 1 3045
0 1182 7 1 2 1177 3046
0 1183 5 2 1 1182
0 1184 7 2 2 1938 2085
0 1185 5 1 1 3049
0 1186 7 1 2 1153 1157
0 1187 5 1 1 1186
0 1188 7 2 2 3030 1187
0 1189 5 1 1 3051
0 1190 7 1 2 3050 3052
0 1191 5 2 1 1190
0 1192 7 2 2 2004 2018
0 1193 5 1 1 3055
0 1194 7 2 2 1982 2041
0 1195 5 1 1 3057
0 1196 7 1 2 1993 2031
0 1197 5 1 1 1196
0 1198 7 1 2 2965 1197
0 1199 5 1 1 1198
0 1200 7 2 2 2970 1199
0 1201 5 1 1 3059
0 1202 7 1 2 3058 3060
0 1203 5 2 1 1202
0 1204 7 1 2 1195 1201
0 1205 5 1 1 1204
0 1206 7 2 2 3061 1205
0 1207 5 1 1 3063
0 1208 7 1 2 3056 3064
0 1209 5 2 1 1208
0 1210 7 1 2 1193 1207
0 1211 5 1 1 1210
0 1212 7 2 2 3065 1211
0 1213 5 1 1 3067
0 1214 7 1 2 1185 1189
0 1215 5 1 1 1214
0 1216 7 2 2 3053 1215
0 1217 5 1 1 3069
0 1218 7 1 2 3068 3070
0 1219 5 2 1 1218
0 1220 7 2 2 3054 3071
0 1221 5 1 1 3073
0 1222 7 1 2 3032 1165
0 1223 5 1 1 1222
0 1224 7 2 2 3036 1223
0 1225 5 1 1 3075
0 1226 7 1 2 1221 3076
0 1227 5 2 1 1226
0 1228 7 2 2 3062 3066
0 1229 5 1 1 3079
0 1230 7 1 2 3074 1225
0 1231 5 1 1 1230
0 1232 7 2 2 3077 1231
0 1233 5 1 1 3081
0 1234 7 1 2 1229 3082
0 1235 5 2 1 1234
0 1236 7 2 2 3078 3083
0 1237 5 1 1 3085
0 1238 7 1 2 3038 1173
0 1239 5 1 1 1238
0 1240 7 2 2 3042 1239
0 1241 5 1 1 3087
0 1242 7 1 2 1237 3088
0 1243 5 2 1 1242
0 1244 7 2 2 1971 2042
0 1245 5 1 1 3091
0 1246 7 1 2 1063 2961
0 1247 5 1 1 1246
0 1248 7 2 2 2966 1247
0 1249 5 1 1 3093
0 1250 7 1 2 3092 3094
0 1251 5 2 1 1250
0 1252 7 2 2 1994 2019
0 1253 5 1 1 3097
0 1254 7 1 2 1245 1249
0 1255 5 1 1 1254
0 1256 7 2 2 3095 1255
0 1257 5 1 1 3099
0 1258 7 1 2 3098 3100
0 1259 5 2 1 1258
0 1260 7 2 2 3096 3101
0 1261 5 1 1 3103
0 1262 7 1 2 1213 1217
0 1263 5 1 1 1262
0 1264 7 2 2 3072 1263
0 1265 5 1 1 3105
0 1266 7 1 2 1261 3106
0 1267 5 2 1 1266
0 1268 7 2 2 1960 2054
0 1269 5 1 1 3109
0 1270 7 2 2 1939 2075
0 1271 5 1 1 3111
0 1272 7 1 2 3110 3112
0 1273 5 2 1 1272
0 1274 7 1 2 1253 1257
0 1275 5 1 1 1274
0 1276 7 2 2 3102 1275
0 1277 5 1 1 3115
0 1278 7 1 2 1269 1271
0 1279 5 1 1 1278
0 1280 7 2 2 3113 1279
0 1281 5 1 1 3117
0 1282 7 1 2 3116 3118
0 1283 5 2 1 1282
0 1284 7 2 2 3114 3119
0 1285 5 1 1 3121
0 1286 7 1 2 3104 1265
0 1287 5 1 1 1286
0 1288 7 2 2 3107 1287
0 1289 5 1 1 3123
0 1290 7 1 2 1285 3124
0 1291 5 2 1 1290
0 1292 7 2 2 3108 3125
0 1293 5 1 1 3127
0 1294 7 1 2 3080 1233
0 1295 5 1 1 1294
0 1296 7 2 2 3084 1295
0 1297 5 1 1 3129
0 1298 7 1 2 1293 3130
0 1299 5 2 1 1298
0 1300 7 2 2 1948 2064
0 1301 5 1 1 3133
0 1302 7 1 2 1277 1281
0 1303 5 1 1 1302
0 1304 7 2 2 3120 1303
0 1305 5 1 1 3135
0 1306 7 1 2 3134 3136
0 1307 5 2 1 1306
0 1308 7 2 2 1961 2043
0 1309 5 1 1 3139
0 1310 7 1 2 1972 2032
0 1311 5 1 1 1310
0 1312 7 1 2 2957 1311
0 1313 5 1 1 1312
0 1314 7 2 2 2962 1313
0 1315 5 1 1 3141
0 1316 7 1 2 3140 3142
0 1317 5 2 1 1316
0 1318 7 2 2 1983 2020
0 1319 5 1 1 3145
0 1320 7 1 2 1309 1315
0 1321 5 1 1 1320
0 1322 7 2 2 3143 1321
0 1323 5 1 1 3147
0 1324 7 1 2 3146 3148
0 1325 5 2 1 1324
0 1326 7 2 2 3144 3149
0 1327 5 1 1 3151
0 1328 7 1 2 1301 1305
0 1329 5 1 1 1328
0 1330 7 2 2 3137 1329
0 1331 5 1 1 3153
0 1332 7 1 2 1327 3154
0 1333 5 2 1 1332
0 1334 7 2 2 3138 3155
0 1335 5 1 1 3157
0 1336 7 1 2 3122 1289
0 1337 5 1 1 1336
0 1338 7 2 2 3126 1337
0 1339 5 1 1 3159
0 1340 7 1 2 1335 3160
0 1341 5 2 1 1340
0 1342 7 2 2 1940 2065
0 1343 5 1 1 3163
0 1344 7 2 2 1949 2055
0 1345 5 1 1 3165
0 1346 7 1 2 3164 3166
0 1347 5 2 1 1346
0 1348 7 1 2 1319 1323
0 1349 5 1 1 1348
0 1350 7 2 2 3150 1349
0 1351 5 1 1 3169
0 1352 7 1 2 1343 1345
0 1353 5 1 1 1352
0 1354 7 2 2 3167 1353
0 1355 5 1 1 3171
0 1356 7 1 2 3170 3172
0 1357 5 2 1 1356
0 1358 7 2 2 3168 3173
0 1359 5 1 1 3175
0 1360 7 1 2 3152 1331
0 1361 5 1 1 1360
0 1362 7 2 2 3156 1361
0 1363 5 1 1 3177
0 1364 7 1 2 1359 3178
0 1365 5 2 1 1364
0 1366 7 1 2 1351 1355
0 1367 5 1 1 1366
0 1368 7 2 2 3174 1367
0 1369 5 1 1 3181
0 1370 7 2 2 1950 2044
0 1371 5 1 1 3183
0 1372 7 2 2 1973 2021
0 1373 5 1 1 3185
0 1374 7 2 2 3184 3186
0 1375 5 1 1 3187
0 1376 7 2 2 1951 2033
0 1377 5 1 1 3189
0 1378 7 2 2 1941 2045
0 1379 5 1 1 3191
0 1380 7 2 2 3190 3192
0 1381 5 2 1 3193
0 1382 7 3 2 1375 3195
0 1383 5 1 1 3197
0 1384 7 1 2 3182 1383
0 1385 5 2 1 1384
0 1386 7 1 2 1065 1067
0 1387 5 1 1 1386
0 1388 7 2 2 2958 1387
0 1389 5 1 1 3202
0 1390 7 1 2 1371 1373
0 1391 5 1 1 1390
0 1392 7 1 2 3198 1391
0 1393 5 1 1 1392
0 1394 7 1 2 3188 3194
0 1395 5 1 1 1394
0 1396 7 2 2 1393 1395
0 1397 5 1 1 3204
0 1398 7 1 2 3203 1397
0 1399 5 2 1 1398
0 1400 7 2 2 1962 2022
0 1401 5 1 1 3208
0 1402 7 1 2 1377 1379
0 1403 5 1 1 1402
0 1404 7 2 2 3196 1403
0 1405 5 1 1 3210
0 1406 7 1 2 3209 3211
0 1407 5 2 1 1406
0 1408 7 1 2 1401 1405
0 1409 5 1 1 1408
0 1410 7 2 2 3212 1409
0 1411 5 1 1 3214
0 1412 7 2 2 1942 2034
0 1413 5 1 1 3216
0 1414 7 2 2 1952 2023
0 1415 5 1 1 3218
0 1416 7 2 2 3217 3219
0 1417 5 2 1 3220
0 1418 7 1 2 3215 3221
0 1419 5 2 1 1418
0 1420 7 2 2 3213 3224
0 1421 5 1 1 3226
0 1422 7 1 2 1389 3205
0 1423 5 1 1 1422
0 1424 7 2 2 3206 1423
0 1425 5 1 1 3228
0 1426 7 1 2 1421 3229
0 1427 5 2 1 1426
0 1428 7 2 2 3207 3230
0 1429 5 1 1 3232
0 1430 7 1 2 1369 3199
0 1431 5 1 1 1430
0 1432 7 2 2 3200 1431
0 1433 5 1 1 3234
0 1434 7 1 2 1429 3235
0 1435 5 2 1 1434
0 1436 7 2 2 3201 3236
0 1437 5 1 1 3238
0 1438 7 1 2 3176 1363
0 1439 5 1 1 1438
0 1440 7 2 2 3179 1439
0 1441 5 1 1 3240
0 1442 7 1 2 1437 3241
0 1443 5 2 1 1442
0 1444 7 2 2 3180 3242
0 1445 5 1 1 3244
0 1446 7 1 2 3158 1339
0 1447 5 1 1 1446
0 1448 7 2 2 3161 1447
0 1449 5 1 1 3246
0 1450 7 1 2 1445 3247
0 1451 5 2 1 1450
0 1452 7 2 2 3162 3248
0 1453 5 1 1 3250
0 1454 7 1 2 3128 1297
0 1455 5 1 1 1454
0 1456 7 2 2 3131 1455
0 1457 5 1 1 3252
0 1458 7 1 2 1453 3253
0 1459 5 2 1 1458
0 1460 7 2 2 3132 3254
0 1461 5 1 1 3256
0 1462 7 1 2 3086 1241
0 1463 5 1 1 1462
0 1464 7 2 2 3089 1463
0 1465 5 1 1 3258
0 1466 7 1 2 1461 3259
0 1467 5 2 1 1466
0 1468 7 2 2 3090 3260
0 1469 5 1 1 3262
0 1470 7 1 2 3044 1181
0 1471 5 1 1 1470
0 1472 7 2 2 3047 1471
0 1473 5 1 1 3264
0 1474 7 1 2 1469 3265
0 1475 5 2 1 1474
0 1476 7 2 2 3048 3266
0 1477 5 1 1 3268
0 1478 7 1 2 3002 1123
0 1479 5 1 1 1478
0 1480 7 2 2 3005 1479
0 1481 5 1 1 3270
0 1482 7 1 2 1477 3271
0 1483 5 2 1 1482
0 1484 7 2 2 3006 3272
0 1485 5 1 1 3274
0 1486 7 1 2 2916 1027
0 1487 5 1 1 1486
0 1488 7 2 2 2919 1487
0 1489 5 1 1 3276
0 1490 7 1 2 1485 3277
0 1491 5 2 1 1490
0 1492 7 2 2 2920 3278
0 1493 5 1 1 3280
0 1494 7 1 2 2838 921
0 1495 5 1 1 1494
0 1496 7 2 2 2841 1495
0 1497 5 1 1 3282
0 1498 7 1 2 1493 3283
0 1499 5 2 1 1498
0 1500 7 2 2 2842 3284
0 1501 5 1 1 3286
0 1502 7 1 2 2762 829
0 1503 5 1 1 1502
0 1504 7 2 2 2765 1503
0 1505 5 1 1 3288
0 1506 7 1 2 1501 3289
0 1507 5 2 1 1506
0 1508 7 2 2 2766 3290
0 1509 5 1 1 3292
0 1510 7 1 2 2710 731
0 1511 5 1 1 1510
0 1512 7 2 2 2711 1511
0 1513 5 1 1 3294
0 1514 7 1 2 1509 3295
0 1515 5 2 1 1514
0 1516 7 2 2 2712 3296
0 1517 5 1 1 3298
0 1518 7 2 2 2221 1517
0 1519 5 2 1 3300
0 1520 7 1 2 3293 1513
0 1521 5 1 1 1520
0 1522 7 2 2 3297 1521
0 1523 5 1 1 3304
0 1524 7 1 2 2142 1523
0 1525 5 3 1 1524
0 1526 7 2 2 2146 3299
0 1527 5 2 1 3309
0 1528 7 2 2 3306 3311
0 1529 7 1 2 3287 1505
0 1530 5 1 1 1529
0 1531 7 2 2 3291 1530
0 1532 5 1 1 3315
0 1533 7 1 2 2138 1532
0 1534 5 4 1 1533
0 1535 7 1 2 2217 3316
0 1536 5 4 1 1535
0 1537 7 1 2 3281 1497
0 1538 5 1 1 1537
0 1539 7 2 2 3285 1538
0 1540 5 1 1 3325
0 1541 7 1 2 2135 1540
0 1542 5 5 1 1541
0 1543 7 1 2 2214 3326
0 1544 5 2 1 1543
0 1545 7 1 2 3275 1489
0 1546 5 1 1 1545
0 1547 7 2 2 3279 1546
0 1548 5 1 1 3334
0 1549 7 1 2 2210 3335
0 1550 5 5 1 1549
0 1551 7 3 2 3332 3336
0 1552 7 1 2 2131 1548
0 1553 5 4 1 1552
0 1554 7 1 2 3269 1481
0 1555 5 1 1 1554
0 1556 7 2 2 3273 1555
0 1557 5 1 1 3348
0 1558 7 1 2 2128 1557
0 1559 5 3 1 1558
0 1560 7 1 2 2207 3349
0 1561 5 4 1 1560
0 1562 7 1 2 3263 1473
0 1563 5 1 1 1562
0 1564 7 2 2 3267 1563
0 1565 5 1 1 3357
0 1566 7 1 2 2125 1565
0 1567 5 3 1 1566
0 1568 7 1 2 2204 3358
0 1569 5 3 1 1568
0 1570 7 1 2 3257 1465
0 1571 5 1 1 1570
0 1572 7 2 2 3261 1571
0 1573 5 1 1 3365
0 1574 7 3 2 2201 3366
0 1575 5 4 1 3367
0 1576 7 3 2 2122 1573
0 1577 5 3 1 3374
0 1578 7 1 2 3251 1457
0 1579 5 1 1 1578
0 1580 7 2 2 3255 1579
0 1581 5 1 1 3380
0 1582 7 1 2 2198 3381
0 1583 5 4 1 1582
0 1584 7 2 2 2119 1581
0 1585 5 4 1 3386
0 1586 7 1 2 3245 1449
0 1587 5 1 1 1586
0 1588 7 2 2 3249 1587
0 1589 5 1 1 3392
0 1590 7 1 2 2116 1589
0 1591 5 4 1 1590
0 1592 7 2 2 2195 3393
0 1593 5 3 1 3398
0 1594 7 1 2 3239 1441
0 1595 5 1 1 1594
0 1596 7 2 2 3243 1595
0 1597 5 1 1 3403
0 1598 7 2 2 2192 3404
0 1599 5 5 1 3405
0 1600 7 1 2 2113 1597
0 1601 5 4 1 1600
0 1602 7 1 2 3233 1433
0 1603 5 1 1 1602
0 1604 7 2 2 3237 1603
0 1605 5 1 1 3416
0 1606 7 1 2 2110 1605
0 1607 5 3 1 1606
0 1608 7 1 2 2189 3417
0 1609 5 4 1 1608
0 1610 7 1 2 3227 1425
0 1611 5 1 1 1610
0 1612 7 2 2 3231 1611
0 1613 5 1 1 3425
0 1614 7 1 2 2107 1613
0 1615 5 3 1 1614
0 1616 7 1 2 2186 3426
0 1617 5 4 1 1616
0 1618 7 1 2 1411 3222
0 1619 5 1 1 1618
0 1620 7 2 2 3225 1619
0 1621 5 1 1 3434
0 1622 7 1 2 2183 3435
0 1623 5 2 1 1622
0 1624 7 1 2 1413 1415
0 1625 5 1 1 1624
0 1626 7 2 2 3223 1625
0 1627 5 1 1 3438
0 1628 7 1 2 2180 3439
0 1629 5 1 1 1628
0 1630 7 2 2 3436 1629
0 1631 5 1 1 3440
0 1632 7 1 2 2104 1621
0 1633 5 2 1 1632
0 1634 7 1 2 1631 3442
0 1635 5 1 1 1634
0 1636 7 1 2 2101 1627
0 1637 5 1 1 1636
0 1638 7 2 2 3443 1637
0 1639 5 1 1 3444
0 1640 7 2 2 1943 2024
0 1641 5 1 1 3446
0 1642 7 1 2 2098 1641
0 1643 5 1 1 1642
0 1644 7 2 2 3445 1643
0 1645 5 1 1 3448
0 1646 7 3 2 1635 1645
0 1647 5 1 1 3450
0 1648 7 1 2 3430 3451
0 1649 5 1 1 1648
0 1650 7 2 2 3427 1649
0 1651 5 2 1 3453
0 1652 7 1 2 3421 3455
0 1653 5 1 1 1652
0 1654 7 2 2 3418 1653
0 1655 5 1 1 3457
0 1656 7 1 2 3412 3458
0 1657 5 2 1 1656
0 1658 7 1 2 3407 3459
0 1659 7 1 2 3400 1658
0 1660 5 1 1 1659
0 1661 7 1 2 3394 1660
0 1662 7 2 2 3388 1661
0 1663 5 1 1 3461
0 1664 7 2 2 3382 1663
0 1665 5 2 1 3463
0 1666 7 1 2 3377 3465
0 1667 5 2 1 1666
0 1668 7 1 2 3370 3467
0 1669 7 1 2 3362 1668
0 1670 5 1 1 1669
0 1671 7 2 2 3359 1670
0 1672 5 2 1 3469
0 1673 7 1 2 3353 3471
0 1674 5 1 1 1673
0 1675 7 2 2 3350 1674
0 1676 5 1 1 3473
0 1677 7 2 2 3344 3474
0 1678 5 1 1 3475
0 1679 7 1 2 3341 1678
0 1680 5 1 1 1679
0 1681 7 2 2 3327 1680
0 1682 5 1 1 3477
0 1683 7 1 2 3321 1682
0 1684 5 1 1 1683
0 1685 7 1 2 3317 1684
0 1686 5 2 1 1685
0 1687 7 1 2 2219 3305
0 1688 5 4 1 1687
0 1689 7 1 2 3479 3481
0 1690 5 1 1 1689
0 1691 7 1 2 3313 1690
0 1692 5 1 1 1691
0 1693 7 2 2 3302 1692
0 1694 5 2 1 3485
0 1695 7 2 2 3371 3363
0 1696 7 1 2 2177 3447
0 1697 5 1 1 1696
0 1698 7 3 2 3441 1697
0 1699 5 1 1 3491
0 1700 7 1 2 3437 1639
0 1701 5 1 1 1700
0 1702 7 2 2 1699 1701
0 1703 5 2 1 3494
0 1704 7 1 2 3431 3496
0 1705 5 1 1 1704
0 1706 7 2 2 3428 1705
0 1707 5 2 1 3498
0 1708 7 1 2 3422 3500
0 1709 5 1 1 1708
0 1710 7 2 2 3419 1709
0 1711 5 1 1 3502
0 1712 7 1 2 3408 1711
0 1713 5 1 1 1712
0 1714 7 2 2 3395 1713
0 1715 7 1 2 3413 3504
0 1716 5 1 1 1715
0 1717 7 2 2 3383 3401
0 1718 7 1 2 1716 3506
0 1719 5 1 1 1718
0 1720 7 2 2 3389 1719
0 1721 5 1 1 3508
0 1722 7 1 2 3378 3509
0 1723 5 1 1 1722
0 1724 7 1 2 3489 1723
0 1725 5 1 1 1724
0 1726 7 2 2 3360 1725
0 1727 5 2 1 3510
0 1728 7 1 2 3354 3512
0 1729 5 1 1 1728
0 1730 7 2 2 3351 1729
0 1731 5 2 1 3514
0 1732 7 2 2 3345 3515
0 1733 5 1 1 3518
0 1734 7 2 2 3342 1733
0 1735 5 1 1 3520
0 1736 7 1 2 3328 1735
0 1737 5 2 1 1736
0 1738 7 1 2 3322 3522
0 1739 5 1 1 1738
0 1740 7 2 2 3318 1739
0 1741 5 1 1 3524
0 1742 7 1 2 3314 3525
0 1743 5 1 1 1742
0 1744 7 1 2 3310 3482
0 1745 5 1 1 1744
0 1746 7 2 2 3319 3323
0 1747 5 2 1 3526
0 1748 7 1 2 3523 3528
0 1749 5 1 1 1748
0 1750 7 1 2 3337 3519
0 1751 5 1 1 1750
0 1752 7 1 2 3338 3346
0 1753 5 1 1 1752
0 1754 7 1 2 3516 1753
0 1755 5 1 1 1754
0 1756 7 3 2 3352 3355
0 1757 5 2 1 3530
0 1758 7 1 2 3511 3533
0 1759 5 1 1 1758
0 1760 7 1 2 3513 3531
0 1761 5 1 1 1760
0 1762 7 1 2 1759 1761
0 1763 5 1 1 1762
0 1764 7 3 2 3361 3364
0 1765 5 2 1 3535
0 1766 7 1 2 3372 1721
0 1767 5 1 1 1766
0 1768 7 1 2 3368 3390
0 1769 5 1 1 1768
0 1770 7 1 2 3379 1769
0 1771 7 1 2 1767 1770
0 1772 7 1 2 3536 1771
0 1773 5 1 1 1772
0 1774 7 1 2 3375 3387
0 1775 7 1 2 3538 1774
0 1776 5 1 1 1775
0 1777 7 1 2 1773 1776
0 1778 5 1 1 1777
0 1779 7 1 2 3391 3384
0 1780 5 2 1 1779
0 1781 7 1 2 3396 3540
0 1782 5 1 1 1781
0 1783 7 1 2 3505 3402
0 1784 5 1 1 1783
0 1785 7 1 2 3414 1784
0 1786 5 1 1 1785
0 1787 7 1 2 3415 3409
0 1788 5 2 1 1787
0 1789 7 1 2 3503 3542
0 1790 5 1 1 1789
0 1791 7 3 2 3420 3423
0 1792 5 2 1 3544
0 1793 7 1 2 3499 3545
0 1794 5 1 1 1793
0 1795 7 3 2 3429 3432
0 1796 5 2 1 3549
0 1797 7 1 2 3497 3550
0 1798 5 1 1 1797
0 1799 7 1 2 3492 3449
0 1800 5 2 1 1799
0 1801 7 1 2 3495 3552
0 1802 5 1 1 1801
0 1803 7 1 2 3554 1802
0 1804 7 1 2 1798 1803
0 1805 5 1 1 1804
0 1806 7 1 2 3501 3547
0 1807 5 1 1 1806
0 1808 7 1 2 1805 1807
0 1809 7 1 2 1794 1808
0 1810 5 1 1 1809
0 1811 7 1 2 1790 1810
0 1812 7 1 2 1786 1811
0 1813 7 1 2 1782 1812
0 1814 7 1 2 1778 1813
0 1815 5 1 1 1814
0 1816 7 1 2 1763 1815
0 1817 7 1 2 1755 1816
0 1818 7 1 2 1751 1817
0 1819 7 1 2 1749 1818
0 1820 7 1 2 1745 1819
0 1821 7 1 2 1743 1820
0 1822 7 1 2 3329 3521
0 1823 5 1 1 1822
0 1824 7 1 2 3330 3527
0 1825 5 1 1 1824
0 1826 7 1 2 3339 3517
0 1827 5 1 1 1826
0 1828 7 2 2 3331 3333
0 1829 5 1 1 3556
0 1830 7 2 2 3347 1829
0 1831 5 1 1 3558
0 1832 7 1 2 1827 3559
0 1833 7 1 2 1825 1832
0 1834 5 1 1 1833
0 1835 7 1 2 1823 1834
0 1836 5 1 1 1835
0 1837 7 2 2 3307 3483
0 1838 5 2 1 3560
0 1839 7 1 2 1741 3562
0 1840 5 1 1 1839
0 1841 7 1 2 1836 1840
0 1842 7 1 2 1821 1841
0 1843 7 1 2 3486 1842
0 1844 5 1 1 1843
0 1845 7 1 2 3478 3529
0 1846 5 1 1 1845
0 1847 7 1 2 3468 3537
0 1848 5 1 1 1847
0 1849 7 1 2 3373 1848
0 1850 5 1 1 1849
0 1851 7 1 2 3466 3539
0 1852 5 1 1 1851
0 1853 7 1 2 3369 1852
0 1854 5 1 1 1853
0 1855 7 1 2 3376 3464
0 1856 5 1 1 1855
0 1857 7 1 2 3406 3399
0 1858 5 1 1 1857
0 1859 7 1 2 3541 1858
0 1860 5 1 1 1859
0 1861 7 1 2 3385 3462
0 1862 5 1 1 1861
0 1863 7 1 2 3397 3460
0 1864 5 1 1 1863
0 1865 7 1 2 3410 1864
0 1866 5 1 1 1865
0 1867 7 1 2 1655 3543
0 1868 5 1 1 1867
0 1869 7 1 2 3456 3546
0 1870 5 1 1 1869
0 1871 7 1 2 3452 3553
0 1872 5 1 1 1871
0 1873 7 1 2 1647 3551
0 1874 5 1 1 1873
0 1875 7 1 2 3555 1874
0 1876 7 1 2 1872 1875
0 1877 5 1 1 1876
0 1878 7 1 2 3454 3548
0 1879 5 1 1 1878
0 1880 7 1 2 1877 1879
0 1881 7 1 2 1870 1880
0 1882 5 1 1 1881
0 1883 7 1 2 1868 1882
0 1884 7 1 2 1866 1883
0 1885 7 1 2 1862 1884
0 1886 7 1 2 1860 1885
0 1887 7 1 2 1856 1886
0 1888 7 1 2 1854 1887
0 1889 7 1 2 1850 1888
0 1890 5 1 1 1889
0 1891 7 1 2 3472 3532
0 1892 5 1 1 1891
0 1893 7 1 2 3470 3534
0 1894 5 1 1 1893
0 1895 7 1 2 1892 1894
0 1896 7 1 2 1890 1895
0 1897 7 1 2 3312 1896
0 1898 7 1 2 1846 1897
0 1899 7 1 2 3308 3301
0 1900 5 1 1 1899
0 1901 7 2 2 3340 3557
0 1902 5 1 1 3564
0 1903 7 1 2 3476 3565
0 1904 5 1 1 1903
0 1905 7 1 2 1676 1831
0 1906 7 1 2 1902 1905
0 1907 5 1 1 1906
0 1908 7 1 2 1904 1907
0 1909 5 1 1 1908
0 1910 7 1 2 1900 1909
0 1911 7 1 2 1898 1910
0 1912 7 1 2 3480 3561
0 1913 5 1 1 1912
0 1914 7 1 2 3320 3563
0 1915 5 1 1 1914
0 1916 7 1 2 1913 1915
0 1917 7 1 2 1911 1916
0 1918 7 1 2 3487 1917
0 1919 5 1 1 1918
0 1920 7 1 2 1844 1919
0 1921 7 1 2 729 1920
0 1922 5 1 1 1921
0 1923 7 1 2 3433 3493
0 1924 7 1 2 3424 1923
0 1925 7 1 2 3411 1924
0 1926 7 1 2 3507 1925
0 1927 7 1 2 3490 1926
0 1928 7 1 2 3356 1927
0 1929 7 1 2 3343 1928
0 1930 7 1 2 3324 1929
0 1931 7 1 2 3303 1930
0 1932 7 1 2 3484 1931
0 1933 7 1 2 3488 1932
0 1934 5 1 1 1933
0 1935 7 1 2 2683 1934
0 1936 5 1 1 1935
3 4099 7 0 2 1922 1936
