1 0 0 2 0
2 32 1 0
2 33 1 0
1 1 0 2 0
2 34 1 1
2 35 1 1
1 2 0 2 0
2 36 1 2
2 37 1 2
1 3 0 2 0
2 38 1 3
2 39 1 3
1 4 0 2 0
2 40 1 4
2 41 1 4
1 5 0 2 0
2 42 1 5
2 43 1 5
1 6 0 2 0
2 44 1 6
2 45 1 6
1 7 0 2 0
2 46 1 7
2 47 1 7
1 8 0 2 0
2 48 1 8
2 85 1 8
1 9 0 2 0
2 96 1 9
2 109 1 9
1 10 0 2 0
2 122 1 10
2 135 1 10
1 11 0 2 0
2 148 1 11
2 161 1 11
1 12 0 2 0
2 174 1 12
2 187 1 12
1 13 0 2 0
2 206 1 13
2 223 1 13
1 14 0 2 0
2 240 1 14
2 259 1 14
1 15 0 2 0
2 278 1 15
2 297 1 15
1 16 0 2 0
2 319 1 16
2 325 1 16
1 17 0 2 0
2 326 1 17
2 327 1 17
1 18 0 2 0
2 328 1 18
2 329 1 18
1 19 0 2 0
2 330 1 19
2 331 1 19
1 20 0 2 0
2 332 1 20
2 333 1 20
1 21 0 2 0
2 334 1 21
2 335 1 21
1 22 0 2 0
2 336 1 22
2 337 1 22
1 23 0 2 0
2 338 1 23
2 339 1 23
1 24 0 2 0
2 340 1 24
2 341 1 24
1 25 0 2 0
2 342 1 25
2 343 1 25
1 26 0 2 0
2 344 1 26
2 345 1 26
1 27 0 2 0
2 346 1 27
2 347 1 27
1 28 0 2 0
2 348 1 28
2 349 1 28
1 29 0 2 0
2 350 1 29
2 351 1 29
1 30 0 2 0
2 352 1 30
2 353 1 30
1 31 0 2 0
2 354 1 31
2 355 1 31
2 356 1 81
2 357 1 81
2 358 1 82
2 359 1 82
2 360 1 87
2 361 1 87
2 362 1 90
2 363 1 90
2 364 1 93
2 365 1 93
2 366 1 97
2 367 1 97
2 368 1 100
2 369 1 100
2 370 1 103
2 371 1 103
2 372 1 106
2 373 1 106
2 374 1 110
2 375 1 110
2 376 1 113
2 377 1 113
2 378 1 116
2 379 1 116
2 380 1 119
2 381 1 119
2 382 1 126
2 383 1 126
2 384 1 127
2 385 1 127
2 386 1 129
2 387 1 129
2 388 1 132
2 389 1 132
2 390 1 139
2 391 1 139
2 392 1 140
2 393 1 140
2 394 1 142
2 395 1 142
2 396 1 145
2 397 1 145
2 398 1 150
2 399 1 150
2 400 1 153
2 401 1 153
2 402 1 155
2 403 1 155
2 404 1 158
2 405 1 158
2 406 1 162
2 407 1 162
2 408 1 163
2 409 1 163
2 410 1 164
2 411 1 164
2 412 1 165
2 413 1 165
2 414 1 168
2 415 1 168
2 416 1 168
2 417 1 171
2 418 1 171
2 419 1 176
2 420 1 176
2 421 1 176
2 422 1 178
2 423 1 178
2 424 1 179
2 425 1 179
2 426 1 179
2 427 1 181
2 428 1 181
2 429 1 186
2 430 1 186
2 431 1 189
2 432 1 189
2 433 1 189
2 434 1 191
2 435 1 191
2 436 1 192
2 437 1 192
2 438 1 200
2 439 1 200
2 440 1 203
2 441 1 203
2 442 1 207
2 443 1 207
2 444 1 208
2 445 1 208
2 446 1 210
2 447 1 210
2 448 1 211
2 449 1 211
2 450 1 211
2 451 1 216
2 452 1 216
2 453 1 216
2 454 1 225
2 455 1 225
2 456 1 225
2 457 1 227
2 458 1 227
2 459 1 228
2 460 1 228
2 461 1 228
2 462 1 234
2 463 1 234
2 464 1 236
2 465 1 236
2 466 1 236
2 467 1 241
2 468 1 241
2 469 1 242
2 470 1 242
2 471 1 244
2 472 1 244
2 473 1 244
2 474 1 245
2 475 1 245
2 476 1 245
2 477 1 253
2 478 1 253
2 479 1 254
2 480 1 254
2 481 1 261
2 482 1 261
2 483 1 261
2 484 1 263
2 485 1 263
2 486 1 263
2 487 1 264
2 488 1 264
2 489 1 264
2 490 1 268
2 491 1 268
2 492 1 272
2 493 1 272
2 494 1 280
2 495 1 280
2 496 1 282
2 497 1 282
2 498 1 282
2 499 1 283
2 500 1 283
2 501 1 285
2 502 1 285
2 503 1 291
2 504 1 291
2 505 1 294
2 506 1 294
2 507 1 299
2 508 1 299
2 509 1 301
2 510 1 301
2 511 1 302
2 512 1 302
2 513 1 313
2 514 1 313
0 49 5 1 1 32
0 50 5 1 1 34
0 51 5 1 1 36
0 52 5 1 1 38
0 53 5 1 1 40
0 54 5 1 1 42
0 55 5 1 1 44
0 56 5 1 1 46
0 57 5 1 1 48
0 58 5 1 1 96
0 59 5 1 1 122
0 60 5 1 1 148
0 61 5 1 1 174
0 62 5 1 1 206
0 63 5 1 1 240
0 64 5 1 1 278
0 65 5 1 1 319
0 66 5 1 1 326
0 67 5 1 1 328
0 68 5 1 1 330
0 69 5 1 1 332
0 70 5 1 1 334
0 71 5 1 1 336
0 72 5 1 1 338
0 73 5 1 1 340
0 74 5 1 1 342
0 75 5 1 1 344
0 76 5 1 1 346
0 77 5 1 1 348
0 78 5 1 1 350
0 79 5 1 1 352
0 80 5 1 1 354
0 81 7 2 2 33 325
0 82 5 2 1 356
0 83 7 1 2 49 65
0 84 5 1 1 83
3 683 7 0 2 358 84
0 86 7 1 2 35 327
0 87 5 2 1 86
0 88 7 1 2 50 66
0 89 5 1 1 88
0 90 7 2 2 360 89
0 91 5 1 1 362
0 92 7 1 2 357 363
0 93 5 2 1 92
0 94 7 1 2 359 91
0 95 5 1 1 94
3 684 7 0 2 364 95
0 97 7 2 2 361 365
0 98 5 1 1 366
0 99 7 1 2 37 329
0 100 5 2 1 99
0 101 7 1 2 51 67
0 102 5 1 1 101
0 103 7 2 2 368 102
0 104 5 1 1 370
0 105 7 1 2 98 371
0 106 5 2 1 105
0 107 7 1 2 367 104
0 108 5 1 1 107
3 685 7 0 2 372 108
0 110 7 2 2 369 373
0 111 5 1 1 374
0 112 7 1 2 39 331
0 113 5 2 1 112
0 114 7 1 2 52 68
0 115 5 1 1 114
0 116 7 2 2 376 115
0 117 5 1 1 378
0 118 7 1 2 111 379
0 119 5 2 1 118
0 120 7 1 2 375 117
0 121 5 1 1 120
3 686 7 0 2 380 121
0 123 7 1 2 53 69
0 124 5 1 1 123
0 125 7 1 2 41 333
0 126 5 2 1 125
0 127 7 2 2 124 382
0 128 5 1 1 384
0 129 7 2 2 377 381
0 130 5 1 1 386
0 131 7 1 2 385 130
0 132 5 2 1 131
0 133 7 1 2 128 387
0 134 5 1 1 133
3 687 7 0 2 388 134
0 136 7 1 2 54 70
0 137 5 1 1 136
0 138 7 1 2 43 335
0 139 5 2 1 138
0 140 7 2 2 137 390
0 141 5 1 1 392
0 142 7 2 2 383 389
0 143 5 1 1 394
0 144 7 1 2 393 143
0 145 5 2 1 144
0 146 7 1 2 141 395
0 147 5 1 1 146
3 688 7 0 2 396 147
0 149 7 1 2 45 337
0 150 5 2 1 149
0 151 7 1 2 55 71
0 152 5 1 1 151
0 153 7 2 2 398 152
0 154 5 1 1 400
0 155 7 2 2 391 397
0 156 5 1 1 402
0 157 7 1 2 401 156
0 158 5 2 1 157
0 159 7 1 2 154 403
0 160 5 1 1 159
3 689 7 0 2 404 160
0 162 7 2 2 399 405
0 163 5 2 1 406
0 164 7 2 2 47 339
0 165 5 2 1 410
0 166 7 1 2 56 72
0 167 5 1 1 166
0 168 7 3 2 412 167
0 169 5 1 1 414
0 170 7 1 2 408 415
0 171 5 2 1 170
0 172 7 1 2 407 169
0 173 5 1 1 172
3 690 7 0 2 417 173
0 175 7 1 2 85 341
0 176 5 3 1 175
0 177 7 1 2 57 73
0 178 5 2 1 177
0 179 7 3 2 419 422
0 180 5 1 1 424
0 181 7 2 2 413 418
0 182 5 1 1 427
0 183 7 1 2 180 428
0 184 5 1 1 183
0 185 7 1 2 425 182
0 186 5 2 1 185
3 691 7 0 2 184 429
0 188 7 1 2 109 343
0 189 5 3 1 188
0 190 7 1 2 58 74
0 191 5 2 1 190
0 192 7 2 2 431 434
0 193 5 1 1 436
0 194 7 1 2 416 426
0 195 7 1 2 409 194
0 196 5 1 1 195
0 197 7 1 2 411 423
0 198 5 1 1 197
0 199 7 1 2 420 198
0 200 7 2 2 196 199
0 201 5 1 1 438
0 202 7 1 2 437 201
0 203 5 2 1 202
0 204 7 1 2 193 439
0 205 5 1 1 204
3 692 7 0 2 440 205
0 207 7 2 2 135 345
0 208 5 2 1 442
0 209 7 1 2 59 75
0 210 5 2 1 209
0 211 7 3 2 444 446
0 212 5 1 1 448
0 213 7 1 2 421 432
0 214 7 1 2 430 213
0 215 5 1 1 214
0 216 7 3 2 435 215
0 217 5 1 1 451
0 218 7 1 2 449 217
0 219 5 1 1 218
0 220 7 1 2 212 452
0 221 5 1 1 220
0 222 7 1 2 219 221
3 693 5 0 1 222
0 224 7 1 2 161 347
0 225 5 3 1 224
0 226 7 1 2 60 76
0 227 5 2 1 226
0 228 7 3 2 454 457
0 229 5 1 1 459
0 230 7 1 2 433 441
0 231 5 1 1 230
0 232 7 1 2 447 231
0 233 5 1 1 232
0 234 7 2 2 445 233
0 235 5 1 1 462
0 236 7 3 2 460 235
0 237 5 1 1 464
0 238 7 1 2 229 463
0 239 5 1 1 238
3 694 7 0 2 237 239
0 241 7 2 2 187 349
0 242 5 2 1 467
0 243 7 1 2 61 77
0 244 5 3 1 243
0 245 7 3 2 469 471
0 246 5 1 1 474
0 247 7 1 2 450 461
0 248 7 1 2 453 247
0 249 5 1 1 248
0 250 7 1 2 443 458
0 251 5 1 1 250
0 252 7 1 2 455 251
0 253 7 2 2 249 252
0 254 5 2 1 477
0 255 7 1 2 475 479
0 256 5 1 1 255
0 257 7 1 2 246 478
0 258 5 1 1 257
3 695 7 0 2 256 258
0 260 7 1 2 223 351
0 261 5 3 1 260
0 262 7 1 2 62 78
0 263 5 3 1 262
0 264 7 3 2 481 484
0 265 5 1 1 487
0 266 7 1 2 456 470
0 267 5 1 1 266
0 268 7 2 2 472 267
0 269 5 1 1 490
0 270 7 1 2 465 473
0 271 5 1 1 270
0 272 7 2 2 269 271
0 273 5 1 1 492
0 274 7 1 2 488 273
0 275 5 1 1 274
0 276 7 1 2 265 493
0 277 5 1 1 276
3 696 7 0 2 275 277
0 279 7 1 2 63 79
0 280 5 2 1 279
0 281 7 1 2 259 353
0 282 5 3 1 281
0 283 7 2 2 494 496
0 284 5 1 1 499
0 285 7 2 2 476 489
0 286 7 1 2 480 501
0 287 5 1 1 286
0 288 7 1 2 468 485
0 289 5 1 1 288
0 290 7 1 2 482 289
0 291 7 2 2 287 290
0 292 5 1 1 503
0 293 7 1 2 500 292
0 294 5 2 1 293
0 295 7 1 2 284 504
0 296 5 1 1 295
3 697 7 0 2 505 296
0 298 7 1 2 64 80
0 299 5 2 1 298
0 300 7 1 2 297 355
0 301 5 2 1 300
0 302 7 2 2 507 509
0 303 5 1 1 511
0 304 7 1 2 466 502
0 305 5 1 1 304
0 306 7 1 2 486 491
0 307 5 1 1 306
0 308 7 1 2 483 307
0 309 7 1 2 305 308
0 310 5 1 1 309
0 311 7 1 2 495 310
0 312 5 1 1 311
0 313 7 2 2 497 312
0 314 5 1 1 513
0 315 7 1 2 512 314
0 316 5 1 1 315
0 317 7 1 2 303 514
0 318 5 1 1 317
3 698 7 0 2 316 318
0 320 7 1 2 498 506
0 321 5 1 1 320
0 322 7 1 2 508 321
0 323 5 1 1 322
0 324 7 1 2 510 323
3 699 5 0 1 324
