1 0 0 2 0
2 49 1 0
2 1708 1 0
1 1 0 2 0
2 1709 1 1
2 1710 1 1
1 2 0 2 0
2 1711 1 2
2 1712 1 2
1 3 0 2 0
2 1713 1 3
2 1714 1 3
1 4 0 2 0
2 1715 1 4
2 1716 1 4
1 5 0 2 0
2 1717 1 5
2 1718 1 5
1 6 0 2 0
2 1719 1 6
2 1720 1 6
1 7 0 2 0
2 1721 1 7
2 1722 1 7
1 8 0 2 0
2 1723 1 8
2 1724 1 8
1 9 0 2 0
2 1725 1 9
2 1726 1 9
1 10 0 2 0
2 1727 1 10
2 1728 1 10
1 11 0 2 0
2 1729 1 11
2 1730 1 11
1 12 0 2 0
2 1731 1 12
2 1732 1 12
1 13 0 2 0
2 1733 1 13
2 1734 1 13
1 14 0 2 0
2 1735 1 14
2 1736 1 14
1 15 0 2 0
2 1737 1 15
2 1738 1 15
1 16 0 2 0
2 1739 1 16
2 1740 1 16
1 17 0 2 0
2 1741 1 17
2 1742 1 17
1 18 0 2 0
2 1743 1 18
2 1744 1 18
1 19 0 2 0
2 1745 1 19
2 1746 1 19
1 20 0 2 0
2 1747 1 20
2 1748 1 20
1 21 0 2 0
2 1749 1 21
2 1750 1 21
1 22 0 2 0
2 1751 1 22
2 1752 1 22
1 23 0 2 0
2 1753 1 23
2 1754 1 23
1 24 0 2 0
2 1755 1 24
2 1756 1 24
1 25 0 2 0
2 1757 1 25
2 1758 1 25
1 26 0 2 0
2 1759 1 26
2 1760 1 26
1 27 0 2 0
2 1761 1 27
2 1762 1 27
1 28 0 2 0
2 1763 1 28
2 1764 1 28
1 29 0 2 0
2 1765 1 29
2 1766 1 29
1 30 0 2 0
2 1767 1 30
2 1768 1 30
1 31 0 2 0
2 1769 1 31
2 1770 1 31
1 32 0 2 0
2 1771 1 32
2 1772 1 32
1 33 0 2 0
2 1773 1 33
2 1774 1 33
1 34 0 2 0
2 1775 1 34
2 1776 1 34
1 35 0 2 0
2 1777 1 35
2 1778 1 35
1 36 0 2 0
2 1779 1 36
2 1780 1 36
1 37 0 2 0
2 1781 1 37
2 1782 1 37
1 38 0 2 0
2 1783 1 38
2 1784 1 38
1 39 0 2 0
2 1785 1 39
2 1786 1 39
1 40 0 2 0
2 1787 1 40
2 1788 1 40
1 41 0 2 0
2 1789 1 41
2 1790 1 41
1 42 0 2 0
2 1791 1 42
2 1792 1 42
1 43 0 2 0
2 1793 1 43
2 1794 1 43
1 44 0 2 0
2 1795 1 44
2 1796 1 44
1 45 0 2 0
2 1797 1 45
2 1798 1 45
1 46 0 2 0
2 1799 1 46
2 1800 1 46
1 47 0 2 0
2 1801 1 47
2 1802 1 47
1 48 0 2 0
2 1803 1 48
2 1804 1 48
2 1805 1 68
2 1806 1 68
2 1807 1 69
2 1808 1 69
2 1809 1 70
2 1810 1 70
2 1811 1 71
2 1812 1 71
2 1813 1 72
2 1814 1 72
2 1815 1 73
2 1816 1 73
2 1817 1 74
2 1818 1 74
2 1819 1 75
2 1820 1 75
2 1821 1 76
2 1822 1 76
2 1823 1 77
2 1824 1 77
2 1825 1 78
2 1826 1 78
2 1827 1 79
2 1828 1 79
2 1829 1 80
2 1830 1 80
2 1831 1 100
2 1832 1 100
2 1833 1 102
2 1834 1 102
2 1835 1 104
2 1836 1 104
2 1837 1 105
2 1838 1 105
2 1839 1 106
2 1840 1 106
2 1841 1 106
2 1842 1 109
2 1843 1 109
2 1844 1 112
2 1845 1 112
2 1846 1 114
2 1847 1 114
2 1848 1 117
2 1849 1 117
2 1850 1 120
2 1851 1 120
2 1852 1 122
2 1853 1 122
2 1854 1 125
2 1855 1 125
2 1856 1 128
2 1857 1 128
2 1858 1 130
2 1859 1 130
2 1860 1 133
2 1861 1 133
2 1862 1 136
2 1863 1 136
2 1864 1 138
2 1865 1 138
2 1866 1 141
2 1867 1 141
2 1868 1 144
2 1869 1 144
2 1870 1 146
2 1871 1 146
2 1872 1 149
2 1873 1 149
2 1874 1 152
2 1875 1 152
2 1876 1 154
2 1877 1 154
2 1878 1 157
2 1879 1 157
2 1880 1 160
2 1881 1 160
2 1882 1 162
2 1883 1 162
2 1884 1 165
2 1885 1 165
2 1886 1 168
2 1887 1 168
2 1888 1 170
2 1889 1 170
2 1890 1 173
2 1891 1 173
2 1892 1 176
2 1893 1 176
2 1894 1 178
2 1895 1 178
2 1896 1 181
2 1897 1 181
2 1898 1 184
2 1899 1 184
2 1900 1 186
2 1901 1 186
2 1902 1 189
2 1903 1 189
2 1904 1 192
2 1905 1 192
2 1906 1 194
2 1907 1 194
2 1908 1 197
2 1909 1 197
2 1910 1 200
2 1911 1 200
2 1912 1 202
2 1913 1 202
2 1914 1 205
2 1915 1 205
2 1916 1 208
2 1917 1 208
2 1918 1 210
2 1919 1 210
2 1920 1 213
2 1921 1 213
2 1922 1 214
2 1923 1 214
2 1924 1 216
2 1925 1 216
2 1926 1 219
2 1927 1 219
2 1928 1 219
2 1929 1 219
2 1930 1 220
2 1931 1 220
2 1932 1 220
2 1933 1 221
2 1934 1 221
2 1935 1 227
2 1936 1 227
2 1937 1 227
2 1938 1 227
2 1939 1 228
2 1940 1 228
2 1941 1 228
2 1942 1 230
2 1943 1 230
2 1944 1 230
2 1945 1 232
2 1946 1 232
2 1947 1 232
2 1948 1 233
2 1949 1 233
2 1950 1 239
2 1951 1 239
2 1952 1 239
2 1953 1 239
2 1954 1 240
2 1955 1 240
2 1956 1 240
2 1957 1 242
2 1958 1 242
2 1959 1 242
2 1960 1 244
2 1961 1 244
2 1962 1 244
2 1963 1 245
2 1964 1 245
2 1965 1 251
2 1966 1 251
2 1967 1 251
2 1968 1 251
2 1969 1 252
2 1970 1 252
2 1971 1 252
2 1972 1 254
2 1973 1 254
2 1974 1 254
2 1975 1 256
2 1976 1 256
2 1977 1 256
2 1978 1 257
2 1979 1 257
2 1980 1 263
2 1981 1 263
2 1982 1 263
2 1983 1 263
2 1984 1 264
2 1985 1 264
2 1986 1 264
2 1987 1 266
2 1988 1 266
2 1989 1 266
2 1990 1 268
2 1991 1 268
2 1992 1 268
2 1993 1 269
2 1994 1 269
2 1995 1 275
2 1996 1 275
2 1997 1 275
2 1998 1 276
2 1999 1 276
2 2000 1 278
2 2001 1 278
2 2002 1 278
2 2003 1 280
2 2004 1 280
2 2005 1 280
2 2006 1 281
2 2007 1 281
2 2008 1 287
2 2009 1 287
2 2010 1 288
2 2011 1 288
2 2012 1 290
2 2013 1 290
2 2014 1 290
2 2015 1 292
2 2016 1 292
2 2017 1 292
2 2018 1 293
2 2019 1 293
2 2020 1 299
2 2021 1 299
2 2022 1 302
2 2023 1 302
2 2024 1 302
2 2025 1 304
2 2026 1 304
2 2027 1 304
2 2028 1 307
2 2029 1 307
2 2030 1 309
2 2031 1 309
2 2032 1 310
2 2033 1 310
2 2034 1 310
2 2035 1 313
2 2036 1 313
2 2037 1 314
2 2038 1 314
2 2039 1 317
2 2040 1 317
2 2041 1 318
2 2042 1 318
2 2043 1 321
2 2044 1 321
2 2045 1 322
2 2046 1 322
2 2047 1 325
2 2048 1 325
2 2049 1 326
2 2050 1 326
2 2051 1 329
2 2052 1 329
2 2053 1 330
2 2054 1 330
2 2055 1 333
2 2056 1 333
2 2057 1 334
2 2058 1 334
2 2059 1 337
2 2060 1 337
2 2061 1 338
2 2062 1 338
2 2063 1 339
2 2064 1 339
2 2065 1 345
2 2066 1 345
2 2067 1 345
2 2068 1 345
2 2069 1 346
2 2070 1 346
2 2071 1 346
2 2072 1 348
2 2073 1 348
2 2074 1 348
2 2075 1 350
2 2076 1 350
2 2077 1 350
2 2078 1 351
2 2079 1 351
2 2080 1 351
2 2081 1 352
2 2082 1 352
2 2083 1 357
2 2084 1 357
2 2085 1 357
2 2086 1 357
2 2087 1 358
2 2088 1 358
2 2089 1 358
2 2090 1 359
2 2091 1 359
2 2092 1 365
2 2093 1 365
2 2094 1 365
2 2095 1 365
2 2096 1 366
2 2097 1 366
2 2098 1 366
2 2099 1 368
2 2100 1 368
2 2101 1 368
2 2102 1 370
2 2103 1 370
2 2104 1 370
2 2105 1 371
2 2106 1 371
2 2107 1 371
2 2108 1 372
2 2109 1 372
2 2110 1 373
2 2111 1 373
2 2112 1 379
2 2113 1 379
2 2114 1 380
2 2115 1 380
2 2116 1 380
2 2117 1 382
2 2118 1 382
2 2119 1 382
2 2120 1 384
2 2121 1 384
2 2122 1 384
2 2123 1 385
2 2124 1 385
2 2125 1 391
2 2126 1 391
2 2127 1 391
2 2128 1 391
2 2129 1 392
2 2130 1 392
2 2131 1 392
2 2132 1 394
2 2133 1 394
2 2134 1 394
2 2135 1 396
2 2136 1 396
2 2137 1 396
2 2138 1 397
2 2139 1 397
2 2140 1 403
2 2141 1 403
2 2142 1 404
2 2143 1 404
2 2144 1 404
2 2145 1 406
2 2146 1 406
2 2147 1 406
2 2148 1 408
2 2149 1 408
2 2150 1 408
2 2151 1 411
2 2152 1 411
2 2153 1 412
2 2154 1 412
2 2155 1 415
2 2156 1 415
2 2157 1 416
2 2158 1 416
2 2159 1 419
2 2160 1 419
2 2161 1 420
2 2162 1 420
2 2163 1 423
2 2164 1 423
2 2165 1 424
2 2166 1 424
2 2167 1 429
2 2168 1 429
2 2169 1 429
2 2170 1 429
2 2171 1 429
2 2172 1 430
2 2173 1 430
2 2174 1 430
2 2175 1 432
2 2176 1 432
2 2177 1 435
2 2178 1 435
2 2179 1 437
2 2180 1 437
2 2181 1 437
2 2182 1 438
2 2183 1 438
2 2184 1 443
2 2185 1 443
2 2186 1 443
2 2187 1 443
2 2188 1 444
2 2189 1 444
2 2190 1 444
2 2191 1 446
2 2192 1 446
2 2193 1 447
2 2194 1 447
2 2195 1 449
2 2196 1 449
2 2197 1 449
2 2198 1 450
2 2199 1 450
2 2200 1 455
2 2201 1 455
2 2202 1 455
2 2203 1 455
2 2204 1 456
2 2205 1 456
2 2206 1 456
2 2207 1 456
2 2208 1 457
2 2209 1 457
2 2210 1 463
2 2211 1 463
2 2212 1 464
2 2213 1 464
2 2214 1 464
2 2215 1 466
2 2216 1 466
2 2217 1 466
2 2218 1 468
2 2219 1 468
2 2220 1 468
2 2221 1 469
2 2222 1 469
2 2223 1 469
2 2224 1 470
2 2225 1 470
2 2226 1 473
2 2227 1 473
2 2228 1 474
2 2229 1 474
2 2230 1 479
2 2231 1 479
2 2232 1 479
2 2233 1 479
2 2234 1 480
2 2235 1 480
2 2236 1 482
2 2237 1 482
2 2238 1 485
2 2239 1 485
2 2240 1 488
2 2241 1 488
2 2242 1 491
2 2243 1 491
2 2244 1 494
2 2245 1 494
2 2246 1 495
2 2247 1 495
2 2248 1 495
2 2249 1 496
2 2250 1 496
2 2251 1 501
2 2252 1 501
2 2253 1 501
2 2254 1 501
2 2255 1 501
2 2256 1 502
2 2257 1 502
2 2258 1 502
2 2259 1 503
2 2260 1 503
2 2261 1 503
2 2262 1 504
2 2263 1 504
2 2264 1 509
2 2265 1 509
2 2266 1 509
2 2267 1 509
2 2268 1 510
2 2269 1 510
2 2270 1 510
2 2271 1 512
2 2272 1 512
2 2273 1 515
2 2274 1 515
2 2275 1 518
2 2276 1 518
2 2277 1 519
2 2278 1 519
2 2279 1 523
2 2280 1 523
2 2281 1 526
2 2282 1 526
2 2283 1 527
2 2284 1 527
2 2285 1 527
2 2286 1 528
2 2287 1 528
2 2288 1 533
2 2289 1 533
2 2290 1 533
2 2291 1 533
2 2292 1 534
2 2293 1 534
2 2294 1 534
2 2295 1 536
2 2296 1 536
2 2297 1 539
2 2298 1 539
2 2299 1 542
2 2300 1 542
2 2301 1 543
2 2302 1 543
2 2303 1 547
2 2304 1 547
2 2305 1 550
2 2306 1 550
2 2307 1 551
2 2308 1 551
2 2309 1 551
2 2310 1 552
2 2311 1 552
2 2312 1 557
2 2313 1 557
2 2314 1 557
2 2315 1 557
2 2316 1 558
2 2317 1 558
2 2318 1 558
2 2319 1 560
2 2320 1 560
2 2321 1 563
2 2322 1 563
2 2323 1 566
2 2324 1 566
2 2325 1 567
2 2326 1 567
2 2327 1 571
2 2328 1 571
2 2329 1 574
2 2330 1 574
2 2331 1 575
2 2332 1 575
2 2333 1 575
2 2334 1 576
2 2335 1 576
2 2336 1 581
2 2337 1 581
2 2338 1 581
2 2339 1 581
2 2340 1 582
2 2341 1 582
2 2342 1 582
2 2343 1 584
2 2344 1 584
2 2345 1 587
2 2346 1 587
2 2347 1 590
2 2348 1 590
2 2349 1 591
2 2350 1 591
2 2351 1 595
2 2352 1 595
2 2353 1 598
2 2354 1 598
2 2355 1 599
2 2356 1 599
2 2357 1 599
2 2358 1 600
2 2359 1 600
2 2360 1 605
2 2361 1 605
2 2362 1 605
2 2363 1 605
2 2364 1 606
2 2365 1 606
2 2366 1 606
2 2367 1 606
2 2368 1 608
2 2369 1 608
2 2370 1 611
2 2371 1 611
2 2372 1 614
2 2373 1 614
2 2374 1 615
2 2375 1 615
2 2376 1 619
2 2377 1 619
2 2378 1 622
2 2379 1 622
2 2380 1 623
2 2381 1 623
2 2382 1 623
2 2383 1 624
2 2384 1 624
2 2385 1 629
2 2386 1 629
2 2387 1 629
2 2388 1 629
2 2389 1 630
2 2390 1 630
2 2391 1 630
2 2392 1 632
2 2393 1 632
2 2394 1 635
2 2395 1 635
2 2396 1 638
2 2397 1 638
2 2398 1 639
2 2399 1 639
2 2400 1 643
2 2401 1 643
2 2402 1 646
2 2403 1 646
2 2404 1 647
2 2405 1 647
2 2406 1 647
2 2407 1 648
2 2408 1 648
2 2409 1 653
2 2410 1 653
2 2411 1 653
2 2412 1 653
2 2413 1 654
2 2414 1 654
2 2415 1 656
2 2416 1 656
2 2417 1 659
2 2418 1 659
2 2419 1 662
2 2420 1 662
2 2421 1 663
2 2422 1 663
2 2423 1 667
2 2424 1 667
2 2425 1 670
2 2426 1 670
2 2427 1 671
2 2428 1 671
2 2429 1 672
2 2430 1 672
2 2431 1 675
2 2432 1 675
2 2433 1 678
2 2434 1 678
2 2435 1 681
2 2436 1 681
2 2437 1 683
2 2438 1 683
2 2439 1 683
2 2440 1 684
2 2441 1 684
2 2442 1 685
2 2443 1 685
2 2444 1 685
2 2445 1 686
2 2446 1 686
2 2447 1 686
2 2448 1 686
2 2449 1 686
2 2450 1 689
2 2451 1 689
2 2452 1 690
2 2453 1 690
2 2454 1 693
2 2455 1 693
2 2456 1 696
2 2457 1 696
2 2458 1 697
2 2459 1 697
2 2460 1 701
2 2461 1 701
2 2462 1 704
2 2463 1 704
2 2464 1 705
2 2465 1 705
2 2466 1 709
2 2467 1 709
2 2468 1 712
2 2469 1 712
2 2470 1 713
2 2471 1 713
2 2472 1 717
2 2473 1 717
2 2474 1 720
2 2475 1 720
2 2476 1 721
2 2477 1 721
2 2478 1 725
2 2479 1 725
2 2480 1 728
2 2481 1 728
2 2482 1 729
2 2483 1 729
2 2484 1 733
2 2485 1 733
2 2486 1 736
2 2487 1 736
2 2488 1 737
2 2489 1 737
2 2490 1 741
2 2491 1 741
2 2492 1 744
2 2493 1 744
2 2494 1 745
2 2495 1 745
2 2496 1 749
2 2497 1 749
2 2498 1 752
2 2499 1 752
2 2500 1 753
2 2501 1 753
2 2502 1 757
2 2503 1 757
2 2504 1 760
2 2505 1 760
2 2506 1 761
2 2507 1 761
2 2508 1 761
2 2509 1 762
2 2510 1 762
2 2511 1 763
2 2512 1 763
2 2513 1 765
2 2514 1 765
2 2515 1 771
2 2516 1 771
2 2517 1 771
2 2518 1 771
2 2519 1 772
2 2520 1 772
2 2521 1 772
2 2522 1 774
2 2523 1 774
2 2524 1 774
2 2525 1 776
2 2526 1 776
2 2527 1 776
2 2528 1 777
2 2529 1 777
2 2530 1 777
2 2531 1 778
2 2532 1 778
2 2533 1 781
2 2534 1 781
2 2535 1 782
2 2536 1 782
2 2537 1 787
2 2538 1 787
2 2539 1 788
2 2540 1 788
2 2541 1 790
2 2542 1 790
2 2543 1 793
2 2544 1 793
2 2545 1 796
2 2546 1 796
2 2547 1 799
2 2548 1 799
2 2549 1 802
2 2550 1 802
2 2551 1 803
2 2552 1 803
2 2553 1 804
2 2554 1 804
2 2555 1 805
2 2556 1 805
2 2557 1 815
2 2558 1 815
2 2559 1 821
2 2560 1 821
2 2561 1 821
2 2562 1 821
2 2563 1 822
2 2564 1 822
2 2565 1 822
2 2566 1 825
2 2567 1 825
2 2568 1 831
2 2569 1 831
2 2570 1 839
2 2571 1 839
2 2572 1 843
2 2573 1 843
2 2574 1 851
2 2575 1 851
2 2576 1 855
2 2577 1 855
2 2578 1 863
2 2579 1 863
2 2580 1 867
2 2581 1 867
2 2582 1 875
2 2583 1 875
2 2584 1 881
2 2585 1 881
2 2586 1 882
2 2587 1 882
2 2588 1 887
2 2589 1 887
2 2590 1 895
2 2591 1 895
2 2592 1 903
2 2593 1 903
2 2594 1 906
2 2595 1 906
2 2596 1 908
2 2597 1 908
2 2598 1 932
2 2599 1 932
2 2600 1 944
2 2601 1 944
2 2602 1 956
2 2603 1 956
2 2604 1 977
2 2605 1 977
2 2606 1 977
2 2607 1 979
2 2608 1 979
2 2609 1 979
2 2610 1 980
2 2611 1 980
2 2612 1 980
2 2613 1 981
2 2614 1 981
2 2615 1 984
2 2616 1 984
2 2617 1 985
2 2618 1 985
2 2619 1 990
2 2620 1 990
2 2621 1 991
2 2622 1 991
2 2623 1 993
2 2624 1 993
2 2625 1 995
2 2626 1 995
2 2627 1 996
2 2628 1 996
2 2629 1 998
2 2630 1 998
2 2631 1 1004
2 2632 1 1004
2 2633 1 1018
2 2634 1 1018
2 2635 1 1019
2 2636 1 1019
2 2637 1 1019
2 2638 1 1023
2 2639 1 1023
2 2640 1 1025
2 2641 1 1025
2 2642 1 1025
2 2643 1 1028
2 2644 1 1028
2 2645 1 1046
2 2646 1 1046
2 2647 1 1061
2 2648 1 1061
2 2649 1 1062
2 2650 1 1062
2 2651 1 1065
2 2652 1 1065
2 2653 1 1066
2 2654 1 1066
2 2655 1 1069
2 2656 1 1069
2 2657 1 1070
2 2658 1 1070
2 2659 1 1073
2 2660 1 1073
2 2661 1 1074
2 2662 1 1074
2 2663 1 1077
2 2664 1 1077
2 2665 1 1078
2 2666 1 1078
2 2667 1 1081
2 2668 1 1081
2 2669 1 1082
2 2670 1 1082
2 2671 1 1085
2 2672 1 1085
2 2673 1 1086
2 2674 1 1086
2 2675 1 1089
2 2676 1 1089
2 2677 1 1090
2 2678 1 1090
2 2679 1 1093
2 2680 1 1093
2 2681 1 1094
2 2682 1 1094
2 2683 1 1097
2 2684 1 1097
2 2685 1 1098
2 2686 1 1098
2 2687 1 1101
2 2688 1 1101
2 2689 1 1102
2 2690 1 1102
2 2691 1 1107
2 2692 1 1107
2 2693 1 1107
2 2694 1 1107
2 2695 1 1108
2 2696 1 1108
2 2697 1 1108
2 2698 1 1113
2 2699 1 1113
2 2700 1 1113
2 2701 1 1113
2 2702 1 1114
2 2703 1 1114
2 2704 1 1114
2 2705 1 1116
2 2706 1 1116
2 2707 1 1119
2 2708 1 1119
2 2709 1 1125
2 2710 1 1125
2 2711 1 1125
2 2712 1 1125
2 2713 1 1126
2 2714 1 1126
2 2715 1 1126
2 2716 1 1128
2 2717 1 1128
2 2718 1 1129
2 2719 1 1129
2 2720 1 1133
2 2721 1 1133
2 2722 1 1134
2 2723 1 1134
2 2724 1 1139
2 2725 1 1139
2 2726 1 1139
2 2727 1 1140
2 2728 1 1140
2 2729 1 1140
2 2730 1 1142
2 2731 1 1142
2 2732 1 1145
2 2733 1 1145
2 2734 1 1151
2 2735 1 1151
2 2736 1 1151
2 2737 1 1151
2 2738 1 1152
2 2739 1 1152
2 2740 1 1152
2 2741 1 1154
2 2742 1 1154
2 2743 1 1157
2 2744 1 1157
2 2745 1 1160
2 2746 1 1160
2 2747 1 1165
2 2748 1 1165
2 2749 1 1165
2 2750 1 1165
2 2751 1 1166
2 2752 1 1166
2 2753 1 1166
2 2754 1 1171
2 2755 1 1171
2 2756 1 1171
2 2757 1 1171
2 2758 1 1172
2 2759 1 1172
2 2760 1 1172
2 2761 1 1174
2 2762 1 1174
2 2763 1 1177
2 2764 1 1177
2 2765 1 1180
2 2766 1 1180
2 2767 1 1181
2 2768 1 1181
2 2769 1 1185
2 2770 1 1185
2 2771 1 1188
2 2772 1 1188
2 2773 1 1193
2 2774 1 1193
2 2775 1 1193
2 2776 1 1193
2 2777 1 1194
2 2778 1 1194
2 2779 1 1194
2 2780 1 1196
2 2781 1 1196
2 2782 1 1199
2 2783 1 1199
2 2784 1 1202
2 2785 1 1202
2 2786 1 1203
2 2787 1 1203
2 2788 1 1207
2 2789 1 1207
2 2790 1 1210
2 2791 1 1210
2 2792 1 1215
2 2793 1 1215
2 2794 1 1215
2 2795 1 1215
2 2796 1 1216
2 2797 1 1216
2 2798 1 1216
2 2799 1 1218
2 2800 1 1218
2 2801 1 1221
2 2802 1 1221
2 2803 1 1224
2 2804 1 1224
2 2805 1 1225
2 2806 1 1225
2 2807 1 1229
2 2808 1 1229
2 2809 1 1232
2 2810 1 1232
2 2811 1 1237
2 2812 1 1237
2 2813 1 1237
2 2814 1 1237
2 2815 1 1238
2 2816 1 1238
2 2817 1 1238
2 2818 1 1240
2 2819 1 1240
2 2820 1 1243
2 2821 1 1243
2 2822 1 1246
2 2823 1 1246
2 2824 1 1247
2 2825 1 1247
2 2826 1 1251
2 2827 1 1251
2 2828 1 1254
2 2829 1 1254
2 2830 1 1259
2 2831 1 1259
2 2832 1 1259
2 2833 1 1259
2 2834 1 1259
2 2835 1 1260
2 2836 1 1260
2 2837 1 1260
2 2838 1 1262
2 2839 1 1262
2 2840 1 1265
2 2841 1 1265
2 2842 1 1268
2 2843 1 1268
2 2844 1 1269
2 2845 1 1269
2 2846 1 1273
2 2847 1 1273
2 2848 1 1276
2 2849 1 1276
2 2850 1 1281
2 2851 1 1281
2 2852 1 1281
2 2853 1 1281
2 2854 1 1282
2 2855 1 1282
2 2856 1 1282
2 2857 1 1284
2 2858 1 1284
2 2859 1 1287
2 2860 1 1287
2 2861 1 1290
2 2862 1 1290
2 2863 1 1291
2 2864 1 1291
2 2865 1 1295
2 2866 1 1295
2 2867 1 1298
2 2868 1 1298
2 2869 1 1303
2 2870 1 1303
2 2871 1 1303
2 2872 1 1304
2 2873 1 1304
2 2874 1 1304
2 2875 1 1306
2 2876 1 1306
2 2877 1 1309
2 2878 1 1309
2 2879 1 1312
2 2880 1 1312
2 2881 1 1313
2 2882 1 1313
2 2883 1 1317
2 2884 1 1317
2 2885 1 1320
2 2886 1 1320
2 2887 1 1321
2 2888 1 1321
2 2889 1 1322
2 2890 1 1322
2 2891 1 1325
2 2892 1 1325
2 2893 1 1328
2 2894 1 1328
2 2895 1 1331
2 2896 1 1331
2 2897 1 1335
2 2898 1 1335
2 2899 1 1336
2 2900 1 1336
2 2901 1 1339
2 2902 1 1339
2 2903 1 1342
2 2904 1 1342
2 2905 1 1343
2 2906 1 1343
2 2907 1 1347
2 2908 1 1347
2 2909 1 1350
2 2910 1 1350
2 2911 1 1351
2 2912 1 1351
2 2913 1 1355
2 2914 1 1355
2 2915 1 1358
2 2916 1 1358
2 2917 1 1359
2 2918 1 1359
2 2919 1 1363
2 2920 1 1363
2 2921 1 1366
2 2922 1 1366
2 2923 1 1367
2 2924 1 1367
2 2925 1 1371
2 2926 1 1371
2 2927 1 1374
2 2928 1 1374
2 2929 1 1375
2 2930 1 1375
2 2931 1 1379
2 2932 1 1379
2 2933 1 1382
2 2934 1 1382
2 2935 1 1383
2 2936 1 1383
2 2937 1 1387
2 2938 1 1387
2 2939 1 1390
2 2940 1 1390
2 2941 1 1391
2 2942 1 1391
2 2943 1 1395
2 2944 1 1395
2 2945 1 1398
2 2946 1 1398
2 2947 1 1399
2 2948 1 1399
2 2949 1 1403
2 2950 1 1403
2 2951 1 1406
2 2952 1 1406
2 2953 1 1407
2 2954 1 1407
2 2955 1 1409
2 2956 1 1409
2 2957 1 1413
2 2958 1 1413
2 2959 1 1414
2 2960 1 1414
2 2961 1 1419
2 2962 1 1419
2 2963 1 1419
2 2964 1 1419
2 2965 1 1420
2 2966 1 1420
2 2967 1 1420
2 2968 1 1422
2 2969 1 1422
2 2970 1 1425
2 2971 1 1425
2 2972 1 1428
2 2973 1 1428
2 2974 1 1431
2 2975 1 1431
2 2976 1 1434
2 2977 1 1434
2 2978 1 1437
2 2979 1 1437
2 2980 1 1440
2 2981 1 1440
2 2982 1 1443
2 2983 1 1443
2 2984 1 1449
2 2985 1 1449
2 2986 1 1450
2 2987 1 1450
2 2988 1 1453
2 2989 1 1453
2 2990 1 1454
2 2991 1 1454
2 2992 1 1457
2 2993 1 1457
2 2994 1 1457
2 2995 1 1457
2 2996 1 1458
2 2997 1 1458
2 2998 1 1463
2 2999 1 1463
2 3000 1 1463
2 3001 1 1464
2 3002 1 1464
2 3003 1 1466
2 3004 1 1466
2 3005 1 1469
2 3006 1 1469
2 3007 1 1469
2 3008 1 1470
2 3009 1 1470
2 3010 1 1472
2 3011 1 1472
2 3012 1 1473
2 3013 1 1473
2 3014 1 1475
2 3015 1 1475
2 3016 1 1481
2 3017 1 1481
2 3018 1 1481
2 3019 1 1482
2 3020 1 1482
2 3021 1 1487
2 3022 1 1487
2 3023 1 1491
2 3024 1 1491
2 3025 1 1494
2 3026 1 1494
2 3027 1 1497
2 3028 1 1497
2 3029 1 1498
2 3030 1 1498
2 3031 1 1500
2 3032 1 1500
2 3033 1 1503
2 3034 1 1503
2 3035 1 1506
2 3036 1 1506
2 3037 1 1512
2 3038 1 1512
2 3039 1 1515
2 3040 1 1515
2 3041 1 1522
2 3042 1 1522
2 3043 1 1524
2 3044 1 1524
2 3045 1 1528
2 3046 1 1528
2 3047 1 1542
2 3048 1 1542
2 3049 1 1550
2 3050 1 1550
2 3051 1 1554
2 3052 1 1554
2 3053 1 1562
2 3054 1 1562
2 3055 1 1566
2 3056 1 1566
2 3057 1 1574
2 3058 1 1574
2 3059 1 1578
2 3060 1 1578
2 3061 1 1586
2 3062 1 1586
2 3063 1 1592
2 3064 1 1592
2 3065 1 1593
2 3066 1 1593
2 3067 1 1598
2 3068 1 1598
2 3069 1 1606
2 3070 1 1606
2 3071 1 1637
2 3072 1 1637
2 3073 1 1649
2 3074 1 1649
2 3075 1 1661
2 3076 1 1661
2 3077 1 1677
2 3078 1 1677
0 50 5 1 1 49
0 51 5 1 1 1709
0 52 5 1 1 1711
0 53 5 1 1 1713
0 54 5 1 1 1715
0 55 5 1 1 1717
0 56 5 1 1 1719
0 57 5 1 1 1721
0 58 5 1 1 1723
0 59 5 1 1 1725
0 60 5 1 1 1727
0 61 5 1 1 1729
0 62 5 1 1 1731
0 63 5 1 1 1733
0 64 5 1 1 1735
0 65 5 1 1 1737
0 66 5 1 1 1739
0 67 5 1 1 1741
0 68 5 2 1 1743
0 69 5 2 1 1745
0 70 5 2 1 1747
0 71 5 2 1 1749
0 72 5 2 1 1751
0 73 5 2 1 1753
0 74 5 2 1 1755
0 75 5 2 1 1757
0 76 5 2 1 1759
0 77 5 2 1 1761
0 78 5 2 1 1763
0 79 5 2 1 1765
0 80 5 2 1 1767
0 81 5 1 1 1769
0 82 5 1 1 1771
0 83 5 1 1 1773
0 84 5 1 1 1775
0 85 5 1 1 1777
0 86 5 1 1 1779
0 87 5 1 1 1781
0 88 5 1 1 1783
0 89 5 1 1 1785
0 90 5 1 1 1787
0 91 5 1 1 1789
0 92 5 1 1 1791
0 93 5 1 1 1793
0 94 5 1 1 1795
0 95 5 1 1 1797
0 96 5 1 1 1799
0 97 5 1 1 1801
0 98 5 1 1 1803
0 99 7 1 2 65 81
0 100 5 2 1 99
0 101 7 1 2 51 67
0 102 5 2 1 101
0 103 7 1 2 1710 1742
0 104 5 2 1 103
0 105 7 2 2 1708 1740
0 106 5 3 1 1837
0 107 7 1 2 1835 1839
0 108 5 1 1 107
0 109 7 2 2 1833 108
0 110 5 1 1 1842
0 111 7 1 2 52 110
0 112 5 2 1 111
0 113 7 1 2 1712 1843
0 114 5 2 1 113
0 115 7 1 2 1805 1846
0 116 5 1 1 115
0 117 7 2 2 1844 116
0 118 5 1 1 1848
0 119 7 1 2 53 118
0 120 5 2 1 119
0 121 7 1 2 1714 1849
0 122 5 2 1 121
0 123 7 1 2 1807 1852
0 124 5 1 1 123
0 125 7 2 2 1850 124
0 126 5 1 1 1854
0 127 7 1 2 54 126
0 128 5 2 1 127
0 129 7 1 2 1716 1855
0 130 5 2 1 129
0 131 7 1 2 1809 1858
0 132 5 1 1 131
0 133 7 2 2 1856 132
0 134 5 1 1 1860
0 135 7 1 2 55 134
0 136 5 2 1 135
0 137 7 1 2 1718 1861
0 138 5 2 1 137
0 139 7 1 2 1811 1864
0 140 5 1 1 139
0 141 7 2 2 1862 140
0 142 5 1 1 1866
0 143 7 1 2 56 142
0 144 5 2 1 143
0 145 7 1 2 1720 1867
0 146 5 2 1 145
0 147 7 1 2 1813 1870
0 148 5 1 1 147
0 149 7 2 2 1868 148
0 150 5 1 1 1872
0 151 7 1 2 57 150
0 152 5 2 1 151
0 153 7 1 2 1722 1873
0 154 5 2 1 153
0 155 7 1 2 1815 1876
0 156 5 1 1 155
0 157 7 2 2 1874 156
0 158 5 1 1 1878
0 159 7 1 2 58 158
0 160 5 2 1 159
0 161 7 1 2 1724 1879
0 162 5 2 1 161
0 163 7 1 2 1817 1882
0 164 5 1 1 163
0 165 7 2 2 1880 164
0 166 5 1 1 1884
0 167 7 1 2 59 166
0 168 5 2 1 167
0 169 7 1 2 1726 1885
0 170 5 2 1 169
0 171 7 1 2 1819 1888
0 172 5 1 1 171
0 173 7 2 2 1886 172
0 174 5 1 1 1890
0 175 7 1 2 60 174
0 176 5 2 1 175
0 177 7 1 2 1728 1891
0 178 5 2 1 177
0 179 7 1 2 1821 1894
0 180 5 1 1 179
0 181 7 2 2 1892 180
0 182 5 1 1 1896
0 183 7 1 2 61 182
0 184 5 2 1 183
0 185 7 1 2 1730 1897
0 186 5 2 1 185
0 187 7 1 2 1823 1900
0 188 5 1 1 187
0 189 7 2 2 1898 188
0 190 5 1 1 1902
0 191 7 1 2 62 190
0 192 5 2 1 191
0 193 7 1 2 1732 1903
0 194 5 2 1 193
0 195 7 1 2 1825 1906
0 196 5 1 1 195
0 197 7 2 2 1904 196
0 198 5 1 1 1908
0 199 7 1 2 63 198
0 200 5 2 1 199
0 201 7 1 2 1734 1909
0 202 5 2 1 201
0 203 7 1 2 1827 1912
0 204 5 1 1 203
0 205 7 2 2 1910 204
0 206 5 1 1 1914
0 207 7 1 2 64 206
0 208 5 2 1 207
0 209 7 1 2 1736 1915
0 210 5 2 1 209
0 211 7 1 2 1829 1918
0 212 5 1 1 211
0 213 7 2 2 1916 212
0 214 5 2 1 1920
0 215 7 1 2 1738 1770
0 216 5 2 1 215
0 217 7 1 2 1922 1924
0 218 5 1 1 217
0 219 7 4 2 1831 218
0 220 5 3 1 1926
0 221 7 2 2 1875 1877
0 222 5 1 1 1933
0 223 7 1 2 1754 1934
0 224 5 1 1 223
0 225 7 1 2 1816 222
0 226 5 1 1 225
0 227 7 4 2 224 226
0 228 5 3 1 1935
0 229 7 1 2 89 1936
0 230 5 3 1 229
0 231 7 1 2 1786 1939
0 232 5 3 1 231
0 233 7 2 2 1869 1871
0 234 5 1 1 1948
0 235 7 1 2 1752 1949
0 236 5 1 1 235
0 237 7 1 2 1814 234
0 238 5 1 1 237
0 239 7 4 2 236 238
0 240 5 3 1 1950
0 241 7 1 2 88 1951
0 242 5 3 1 241
0 243 7 1 2 1784 1954
0 244 5 3 1 243
0 245 7 2 2 1863 1865
0 246 5 1 1 1963
0 247 7 1 2 1750 1964
0 248 5 1 1 247
0 249 7 1 2 1812 246
0 250 5 1 1 249
0 251 7 4 2 248 250
0 252 5 3 1 1965
0 253 7 1 2 87 1966
0 254 5 3 1 253
0 255 7 1 2 1782 1969
0 256 5 3 1 255
0 257 7 2 2 1857 1859
0 258 5 1 1 1978
0 259 7 1 2 1748 1979
0 260 5 1 1 259
0 261 7 1 2 1810 258
0 262 5 1 1 261
0 263 7 4 2 260 262
0 264 5 3 1 1980
0 265 7 1 2 86 1981
0 266 5 3 1 265
0 267 7 1 2 1780 1984
0 268 5 3 1 267
0 269 7 2 2 1851 1853
0 270 5 1 1 1993
0 271 7 1 2 1746 1994
0 272 5 1 1 271
0 273 7 1 2 1808 270
0 274 5 1 1 273
0 275 7 3 2 272 274
0 276 5 2 1 1995
0 277 7 1 2 85 1996
0 278 5 3 1 277
0 279 7 1 2 1778 1998
0 280 5 3 1 279
0 281 7 2 2 1845 1847
0 282 5 1 1 2006
0 283 7 1 2 1744 2007
0 284 5 1 1 283
0 285 7 1 2 1806 282
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 2 1 2008
0 289 7 1 2 84 2009
0 290 5 3 1 289
0 291 7 1 2 1776 2010
0 292 5 3 1 291
0 293 7 2 2 1834 1836
0 294 5 1 1 2018
0 295 7 1 2 1838 294
0 296 5 1 1 295
0 297 7 1 2 1840 2019
0 298 5 1 1 297
0 299 7 2 2 296 298
0 300 5 1 1 2020
0 301 7 1 2 83 300
0 302 5 3 1 301
0 303 7 1 2 1774 2021
0 304 5 3 1 303
0 305 7 1 2 50 66
0 306 5 1 1 305
0 307 7 2 2 1841 306
0 308 5 1 1 2028
0 309 7 2 2 1772 308
0 310 5 3 1 2030
0 311 7 1 2 2025 2032
0 312 5 1 1 311
0 313 7 2 2 2022 312
0 314 5 2 1 2035
0 315 7 1 2 2015 2037
0 316 5 1 1 315
0 317 7 2 2 2012 316
0 318 5 2 1 2039
0 319 7 1 2 2003 2041
0 320 5 1 1 319
0 321 7 2 2 2000 320
0 322 5 2 1 2043
0 323 7 1 2 1990 2045
0 324 5 1 1 323
0 325 7 2 2 1987 324
0 326 5 2 1 2047
0 327 7 1 2 1975 2049
0 328 5 1 1 327
0 329 7 2 2 1972 328
0 330 5 2 1 2051
0 331 7 1 2 1960 2053
0 332 5 1 1 331
0 333 7 2 2 1957 332
0 334 5 2 1 2055
0 335 7 1 2 1945 2057
0 336 5 1 1 335
0 337 7 2 2 1942 336
0 338 5 2 1 2059
0 339 7 2 2 1881 1883
0 340 5 1 1 2063
0 341 7 1 2 1756 2064
0 342 5 1 1 341
0 343 7 1 2 1818 340
0 344 5 1 1 343
0 345 7 4 2 342 344
0 346 5 3 1 2065
0 347 7 1 2 90 2066
0 348 5 3 1 347
0 349 7 1 2 1788 2069
0 350 5 3 1 349
0 351 7 3 2 2072 2075
0 352 5 2 1 2078
0 353 7 1 2 2060 2079
0 354 5 1 1 353
0 355 7 1 2 2061 2081
0 356 5 1 1 355
0 357 7 4 2 354 356
0 358 5 3 1 2083
0 359 7 2 2 1905 1907
0 360 5 1 1 2090
0 361 7 1 2 1764 2091
0 362 5 1 1 361
0 363 7 1 2 1826 360
0 364 5 1 1 363
0 365 7 4 2 362 364
0 366 5 3 1 2092
0 367 7 1 2 94 2093
0 368 5 3 1 367
0 369 7 1 2 1796 2096
0 370 5 3 1 369
0 371 7 3 2 2099 2102
0 372 5 2 1 2105
0 373 7 2 2 1899 1901
0 374 5 1 1 2110
0 375 7 1 2 1762 2111
0 376 5 1 1 375
0 377 7 1 2 1824 374
0 378 5 1 1 377
0 379 7 2 2 376 378
0 380 5 3 1 2112
0 381 7 1 2 93 2113
0 382 5 3 1 381
0 383 7 1 2 1794 2114
0 384 5 3 1 383
0 385 7 2 2 1893 1895
0 386 5 1 1 2123
0 387 7 1 2 1760 2124
0 388 5 1 1 387
0 389 7 1 2 1822 386
0 390 5 1 1 389
0 391 7 4 2 388 390
0 392 5 3 1 2125
0 393 7 1 2 92 2126
0 394 5 3 1 393
0 395 7 1 2 1792 2129
0 396 5 3 1 395
0 397 7 2 2 1887 1889
0 398 5 1 1 2138
0 399 7 1 2 1758 2139
0 400 5 1 1 399
0 401 7 1 2 1820 398
0 402 5 1 1 401
0 403 7 2 2 400 402
0 404 5 3 1 2140
0 405 7 1 2 91 2141
0 406 5 3 1 405
0 407 7 1 2 1790 2142
0 408 5 3 1 407
0 409 7 1 2 2076 2062
0 410 5 1 1 409
0 411 7 2 2 2073 410
0 412 5 2 1 2151
0 413 7 1 2 2148 2153
0 414 5 1 1 413
0 415 7 2 2 2145 414
0 416 5 2 1 2155
0 417 7 1 2 2135 2157
0 418 5 1 1 417
0 419 7 2 2 2132 418
0 420 5 2 1 2159
0 421 7 1 2 2120 2161
0 422 5 1 1 421
0 423 7 2 2 2117 422
0 424 5 2 1 2163
0 425 7 1 2 2106 2164
0 426 5 1 1 425
0 427 7 1 2 2108 2165
0 428 5 1 1 427
0 429 7 5 2 426 428
0 430 5 3 1 2167
0 431 7 1 2 2087 2172
0 432 5 2 1 431
0 433 7 1 2 2084 2168
0 434 5 1 1 433
0 435 7 2 2 2175 434
0 436 5 1 1 2177
0 437 7 3 2 2146 2149
0 438 5 2 1 2179
0 439 7 1 2 2152 2180
0 440 5 1 1 439
0 441 7 1 2 2154 2182
0 442 5 1 1 441
0 443 7 4 2 440 442
0 444 5 3 1 2184
0 445 7 1 2 2178 2188
0 446 5 2 1 445
0 447 7 2 2 2176 2191
0 448 5 1 1 2193
0 449 7 3 2 2133 2136
0 450 5 2 1 2195
0 451 7 1 2 2156 2198
0 452 5 1 1 451
0 453 7 1 2 2158 2196
0 454 5 1 1 453
0 455 7 4 2 452 454
0 456 5 4 1 2200
0 457 7 2 2 1911 1913
0 458 5 1 1 2208
0 459 7 1 2 1766 2209
0 460 5 1 1 459
0 461 7 1 2 1828 458
0 462 5 1 1 461
0 463 7 2 2 460 462
0 464 5 3 1 2210
0 465 7 1 2 1798 2212
0 466 5 3 1 465
0 467 7 1 2 95 2211
0 468 5 3 1 467
0 469 7 3 2 2215 2218
0 470 5 2 1 2221
0 471 7 1 2 2103 2166
0 472 5 1 1 471
0 473 7 2 2 2100 472
0 474 5 2 1 2226
0 475 7 1 2 2222 2227
0 476 5 1 1 475
0 477 7 1 2 2224 2228
0 478 5 1 1 477
0 479 7 4 2 476 478
0 480 5 2 1 2230
0 481 7 1 2 2189 2234
0 482 5 2 1 481
0 483 7 1 2 2185 2231
0 484 5 1 1 483
0 485 7 2 2 2236 484
0 486 5 1 1 2238
0 487 7 1 2 2201 2239
0 488 5 2 1 487
0 489 7 1 2 2204 486
0 490 5 1 1 489
0 491 7 2 2 2240 490
0 492 5 1 1 2242
0 493 7 1 2 448 2243
0 494 5 2 1 493
0 495 7 3 2 2121 2118
0 496 5 2 1 2246
0 497 7 1 2 2249 2160
0 498 5 1 1 497
0 499 7 1 2 2247 2162
0 500 5 1 1 499
0 501 7 5 2 498 500
0 502 5 3 1 2251
0 503 7 3 2 1943 1946
0 504 5 2 1 2259
0 505 7 1 2 2056 2262
0 506 5 1 1 505
0 507 7 1 2 2058 2260
0 508 5 1 1 507
0 509 7 4 2 506 508
0 510 5 3 1 2264
0 511 7 1 2 2252 2265
0 512 5 2 1 511
0 513 7 1 2 2256 2268
0 514 5 1 1 513
0 515 7 2 2 2271 514
0 516 5 1 1 2273
0 517 7 1 2 2274 2088
0 518 5 2 1 517
0 519 7 2 2 2272 2275
0 520 5 1 1 2277
0 521 7 1 2 436 2186
0 522 5 1 1 521
0 523 7 2 2 2192 522
0 524 5 1 1 2279
0 525 7 1 2 520 2280
0 526 5 2 1 525
0 527 7 3 2 1958 1961
0 528 5 2 1 2283
0 529 7 1 2 2052 2286
0 530 5 1 1 529
0 531 7 1 2 2054 2284
0 532 5 1 1 531
0 533 7 4 2 530 532
0 534 5 3 1 2288
0 535 7 1 2 2202 2289
0 536 5 2 1 535
0 537 7 1 2 2205 2292
0 538 5 1 1 537
0 539 7 2 2 2295 538
0 540 5 1 1 2297
0 541 7 1 2 2266 2298
0 542 5 2 1 541
0 543 7 2 2 2296 2299
0 544 5 1 1 2301
0 545 7 1 2 516 2085
0 546 5 1 1 545
0 547 7 2 2 2276 546
0 548 5 1 1 2303
0 549 7 1 2 544 2304
0 550 5 2 1 549
0 551 7 3 2 1973 1976
0 552 5 2 1 2307
0 553 7 1 2 2048 2310
0 554 5 1 1 553
0 555 7 1 2 2050 2308
0 556 5 1 1 555
0 557 7 4 2 554 556
0 558 5 3 1 2312
0 559 7 1 2 2190 2313
0 560 5 2 1 559
0 561 7 1 2 2187 2316
0 562 5 1 1 561
0 563 7 2 2 2319 562
0 564 5 1 1 2321
0 565 7 1 2 2290 2322
0 566 5 2 1 565
0 567 7 2 2 2320 2323
0 568 5 1 1 2325
0 569 7 1 2 2269 540
0 570 5 1 1 569
0 571 7 2 2 2300 570
0 572 5 1 1 2327
0 573 7 1 2 568 2328
0 574 5 2 1 573
0 575 7 3 2 1988 1991
0 576 5 2 1 2331
0 577 7 1 2 2044 2334
0 578 5 1 1 577
0 579 7 1 2 2046 2332
0 580 5 1 1 579
0 581 7 4 2 578 580
0 582 5 3 1 2336
0 583 7 1 2 2089 2337
0 584 5 2 1 583
0 585 7 1 2 2086 2340
0 586 5 1 1 585
0 587 7 2 2 2343 586
0 588 5 1 1 2345
0 589 7 1 2 2314 2346
0 590 5 2 1 589
0 591 7 2 2 2344 2347
0 592 5 1 1 2349
0 593 7 1 2 2293 564
0 594 5 1 1 593
0 595 7 2 2 2324 594
0 596 5 1 1 2351
0 597 7 1 2 592 2352
0 598 5 2 1 597
0 599 7 3 2 2001 2004
0 600 5 2 1 2355
0 601 7 1 2 2040 2358
0 602 5 1 1 601
0 603 7 1 2 2042 2356
0 604 5 1 1 603
0 605 7 4 2 602 604
0 606 5 4 1 2360
0 607 7 1 2 2267 2361
0 608 5 2 1 607
0 609 7 1 2 2270 2364
0 610 5 1 1 609
0 611 7 2 2 2368 610
0 612 5 1 1 2370
0 613 7 1 2 2338 2371
0 614 5 2 1 613
0 615 7 2 2 2369 2372
0 616 5 1 1 2374
0 617 7 1 2 2317 588
0 618 5 1 1 617
0 619 7 2 2 2348 618
0 620 5 1 1 2376
0 621 7 1 2 616 2377
0 622 5 2 1 621
0 623 7 3 2 2013 2016
0 624 5 2 1 2380
0 625 7 1 2 2036 2381
0 626 5 1 1 625
0 627 7 1 2 2038 2383
0 628 5 1 1 627
0 629 7 4 2 626 628
0 630 5 3 1 2385
0 631 7 1 2 2291 2389
0 632 5 2 1 631
0 633 7 1 2 2294 2386
0 634 5 1 1 633
0 635 7 2 2 2392 634
0 636 5 1 1 2394
0 637 7 1 2 2362 2395
0 638 5 2 1 637
0 639 7 2 2 2393 2396
0 640 5 1 1 2398
0 641 7 1 2 2341 612
0 642 5 1 1 641
0 643 7 2 2 2373 642
0 644 5 1 1 2400
0 645 7 1 2 640 2401
0 646 5 2 1 645
0 647 7 3 2 2023 2026
0 648 5 2 1 2404
0 649 7 1 2 2031 2405
0 650 5 1 1 649
0 651 7 1 2 2033 2407
0 652 5 1 1 651
0 653 7 4 2 650 652
0 654 5 2 1 2409
0 655 7 1 2 2315 2413
0 656 5 2 1 655
0 657 7 1 2 2318 2410
0 658 5 1 1 657
0 659 7 2 2 2415 658
0 660 5 1 1 2417
0 661 7 1 2 2390 2418
0 662 5 2 1 661
0 663 7 2 2 2416 2419
0 664 5 1 1 2421
0 665 7 1 2 2365 636
0 666 5 1 1 665
0 667 7 2 2 2397 666
0 668 5 1 1 2423
0 669 7 1 2 664 2424
0 670 5 2 1 669
0 671 7 2 2 2339 2414
0 672 5 2 1 2427
0 673 7 1 2 2387 660
0 674 5 1 1 673
0 675 7 2 2 2420 674
0 676 5 1 1 2431
0 677 7 1 2 2428 2432
0 678 5 2 1 677
0 679 7 1 2 2429 676
0 680 5 1 1 679
0 681 7 2 2 2433 680
0 682 5 1 1 2435
0 683 7 3 2 82 2029
0 684 5 2 1 2437
0 685 7 3 2 2034 2440
0 686 5 5 1 2442
0 687 7 1 2 2342 2411
0 688 5 1 1 687
0 689 7 2 2 2430 688
0 690 5 2 1 2450
0 691 7 1 2 2366 2452
0 692 5 1 1 691
0 693 7 2 2 2445 692
0 694 5 1 1 2454
0 695 7 1 2 2436 2455
0 696 5 2 1 695
0 697 7 2 2 2434 2456
0 698 5 1 1 2458
0 699 7 1 2 2422 668
0 700 5 1 1 699
0 701 7 2 2 2425 700
0 702 5 1 1 2460
0 703 7 1 2 698 2461
0 704 5 2 1 703
0 705 7 2 2 2426 2462
0 706 5 1 1 2464
0 707 7 1 2 2399 644
0 708 5 1 1 707
0 709 7 2 2 2402 708
0 710 5 1 1 2466
0 711 7 1 2 706 2467
0 712 5 2 1 711
0 713 7 2 2 2403 2468
0 714 5 1 1 2470
0 715 7 1 2 2375 620
0 716 5 1 1 715
0 717 7 2 2 2378 716
0 718 5 1 1 2472
0 719 7 1 2 714 2473
0 720 5 2 1 719
0 721 7 2 2 2379 2474
0 722 5 1 1 2476
0 723 7 1 2 2350 596
0 724 5 1 1 723
0 725 7 2 2 2353 724
0 726 5 1 1 2478
0 727 7 1 2 722 2479
0 728 5 2 1 727
0 729 7 2 2 2354 2480
0 730 5 1 1 2482
0 731 7 1 2 2326 572
0 732 5 1 1 731
0 733 7 2 2 2329 732
0 734 5 1 1 2484
0 735 7 1 2 730 2485
0 736 5 2 1 735
0 737 7 2 2 2330 2486
0 738 5 1 1 2488
0 739 7 1 2 2302 548
0 740 5 1 1 739
0 741 7 2 2 2305 740
0 742 5 1 1 2490
0 743 7 1 2 738 2491
0 744 5 2 1 743
0 745 7 2 2 2306 2492
0 746 5 1 1 2494
0 747 7 1 2 2278 524
0 748 5 1 1 747
0 749 7 2 2 2281 748
0 750 5 1 1 2496
0 751 7 1 2 746 2497
0 752 5 2 1 751
0 753 7 2 2 2282 2498
0 754 5 1 1 2500
0 755 7 1 2 2194 492
0 756 5 1 1 755
0 757 7 2 2 2244 756
0 758 5 1 1 2502
0 759 7 1 2 754 2503
0 760 5 2 1 759
0 761 7 3 2 2245 2504
0 762 5 2 1 2506
0 763 7 2 2 2237 2241
0 764 5 1 1 2511
0 765 7 2 2 1917 1919
0 766 5 1 1 2513
0 767 7 1 2 1768 766
0 768 5 1 1 767
0 769 7 1 2 1830 2514
0 770 5 1 1 769
0 771 7 4 2 768 770
0 772 5 3 1 2515
0 773 7 1 2 1800 2516
0 774 5 3 1 773
0 775 7 1 2 96 2519
0 776 5 3 1 775
0 777 7 3 2 2522 2525
0 778 5 2 1 2528
0 779 7 1 2 2216 2229
0 780 5 1 1 779
0 781 7 2 2 2219 780
0 782 5 2 1 2533
0 783 7 1 2 2529 2535
0 784 5 1 1 783
0 785 7 1 2 2531 2534
0 786 5 1 1 785
0 787 7 2 2 784 786
0 788 5 2 1 2537
0 789 7 1 2 2203 2538
0 790 5 2 1 789
0 791 7 1 2 2206 2539
0 792 5 1 1 791
0 793 7 2 2 2541 792
0 794 5 1 1 2543
0 795 7 1 2 2253 2544
0 796 5 2 1 795
0 797 7 1 2 2257 794
0 798 5 1 1 797
0 799 7 2 2 2545 798
0 800 5 1 1 2547
0 801 7 1 2 764 2548
0 802 5 2 1 801
0 803 7 2 2 2512 800
0 804 5 2 1 2551
0 805 7 2 2 2549 2553
0 806 5 1 1 2555
0 807 7 1 2 2507 806
0 808 5 1 1 807
0 809 7 1 2 2509 2556
0 810 5 1 1 809
0 811 7 1 2 808 810
0 812 5 1 1 811
0 813 7 1 2 1927 812
0 814 5 1 1 813
0 815 7 2 2 1925 1832
0 816 5 1 1 2557
0 817 7 1 2 1923 2558
0 818 5 1 1 817
0 819 7 1 2 1921 816
0 820 5 1 1 819
0 821 7 4 2 818 820
0 822 5 3 1 2559
0 823 7 1 2 2501 758
0 824 5 1 1 823
0 825 7 2 2 2505 824
0 826 5 1 1 2566
0 827 7 1 2 2560 2567
0 828 5 1 1 827
0 829 7 1 2 2495 750
0 830 5 1 1 829
0 831 7 2 2 2499 830
0 832 5 1 1 2568
0 833 7 1 2 2517 2569
0 834 5 1 1 833
0 835 7 1 2 2520 832
0 836 5 1 1 835
0 837 7 1 2 2489 742
0 838 5 1 1 837
0 839 7 2 2 2493 838
0 840 5 1 1 2570
0 841 7 1 2 2483 734
0 842 5 1 1 841
0 843 7 2 2 2487 842
0 844 5 1 1 2572
0 845 7 1 2 2097 2573
0 846 5 1 1 845
0 847 7 1 2 2094 844
0 848 5 1 1 847
0 849 7 1 2 2477 726
0 850 5 1 1 849
0 851 7 2 2 2481 850
0 852 5 1 1 2574
0 853 7 1 2 2471 718
0 854 5 1 1 853
0 855 7 2 2 2475 854
0 856 5 1 1 2576
0 857 7 1 2 2130 2577
0 858 5 1 1 857
0 859 7 1 2 2127 856
0 860 5 1 1 859
0 861 7 1 2 2465 710
0 862 5 1 1 861
0 863 7 2 2 2469 862
0 864 5 1 1 2578
0 865 7 1 2 2459 702
0 866 5 1 1 865
0 867 7 2 2 2463 866
0 868 5 1 1 2580
0 869 7 1 2 2070 2581
0 870 5 1 1 869
0 871 7 1 2 2067 868
0 872 5 1 1 871
0 873 7 1 2 682 694
0 874 5 1 1 873
0 875 7 2 2 2457 874
0 876 5 1 1 2582
0 877 7 1 2 1940 2583
0 878 5 1 1 877
0 879 7 1 2 1937 876
0 880 5 1 1 879
0 881 7 2 2 2367 2446
0 882 5 2 1 2584
0 883 7 1 2 2451 2586
0 884 5 1 1 883
0 885 7 1 2 2453 2585
0 886 5 1 1 885
0 887 7 2 2 884 886
0 888 5 1 1 2588
0 889 7 1 2 1955 888
0 890 5 1 1 889
0 891 7 1 2 1952 2589
0 892 5 1 1 891
0 893 7 1 2 2363 2443
0 894 5 1 1 893
0 895 7 2 2 2587 894
0 896 5 1 1 2590
0 897 7 1 2 1967 2591
0 898 5 1 1 897
0 899 7 1 2 1982 2388
0 900 5 1 1 899
0 901 7 1 2 1985 2391
0 902 5 1 1 901
0 903 7 2 2 2011 2447
0 904 5 1 1 2592
0 905 7 1 2 1997 904
0 906 5 2 1 905
0 907 7 1 2 1999 2593
0 908 5 2 1 907
0 909 7 1 2 2412 2596
0 910 5 1 1 909
0 911 7 1 2 2594 910
0 912 5 1 1 911
0 913 7 1 2 902 912
0 914 5 1 1 913
0 915 7 1 2 900 914
0 916 7 1 2 898 915
0 917 5 1 1 916
0 918 7 1 2 1970 896
0 919 5 1 1 918
0 920 7 1 2 917 919
0 921 5 1 1 920
0 922 7 1 2 892 921
0 923 5 1 1 922
0 924 7 1 2 890 923
0 925 5 1 1 924
0 926 7 1 2 880 925
0 927 5 1 1 926
0 928 7 1 2 878 927
0 929 5 1 1 928
0 930 7 1 2 872 929
0 931 5 1 1 930
0 932 7 2 2 870 931
0 933 5 1 1 2598
0 934 7 1 2 2579 933
0 935 5 1 1 934
0 936 7 1 2 864 2599
0 937 5 1 1 936
0 938 7 1 2 2143 937
0 939 5 1 1 938
0 940 7 1 2 935 939
0 941 5 1 1 940
0 942 7 1 2 860 941
0 943 5 1 1 942
0 944 7 2 2 858 943
0 945 5 1 1 2600
0 946 7 1 2 2575 945
0 947 5 1 1 946
0 948 7 1 2 852 2601
0 949 5 1 1 948
0 950 7 1 2 2115 949
0 951 5 1 1 950
0 952 7 1 2 947 951
0 953 5 1 1 952
0 954 7 1 2 848 953
0 955 5 1 1 954
0 956 7 2 2 846 955
0 957 5 1 1 2602
0 958 7 1 2 2571 957
0 959 5 1 1 958
0 960 7 1 2 840 2603
0 961 5 1 1 960
0 962 7 1 2 2213 961
0 963 5 1 1 962
0 964 7 1 2 959 963
0 965 5 1 1 964
0 966 7 1 2 836 965
0 967 5 1 1 966
0 968 7 1 2 834 967
0 969 7 1 2 828 968
0 970 5 1 1 969
0 971 7 1 2 2563 826
0 972 5 1 1 971
0 973 7 1 2 970 972
0 974 7 1 2 814 973
0 975 5 1 1 974
0 976 7 1 2 1802 2561
0 977 5 3 1 976
0 978 7 1 2 97 2564
0 979 5 3 1 978
0 980 7 3 2 2604 2607
0 981 5 2 1 2610
0 982 7 1 2 2523 2536
0 983 5 1 1 982
0 984 7 2 2 2526 983
0 985 5 2 1 2615
0 986 7 1 2 2611 2617
0 987 5 1 1 986
0 988 7 1 2 2613 2616
0 989 5 1 1 988
0 990 7 2 2 987 989
0 991 5 2 1 2619
0 992 7 1 2 2254 2620
0 993 5 2 1 992
0 994 7 1 2 2258 2621
0 995 5 2 1 994
0 996 7 2 2 2623 2625
0 997 5 1 1 2627
0 998 7 2 2 2542 2546
0 999 5 1 1 2629
0 1000 7 1 2 2173 2630
0 1001 5 1 1 1000
0 1002 7 1 2 2169 999
0 1003 5 1 1 1002
0 1004 7 2 2 1001 1003
0 1005 5 1 1 2631
0 1006 7 1 2 997 2632
0 1007 5 1 1 1006
0 1008 7 1 2 2628 1005
0 1009 5 1 1 1008
0 1010 7 1 2 1007 1009
0 1011 5 1 1 1010
0 1012 7 1 2 2508 2552
0 1013 5 1 1 1012
0 1014 7 1 2 1930 1013
0 1015 5 1 1 1014
0 1016 7 1 2 2510 2554
0 1017 5 1 1 1016
0 1018 7 2 2 98 1928
0 1019 5 3 1 2633
0 1020 7 1 2 2605 2618
0 1021 5 1 1 1020
0 1022 7 1 2 2608 1021
0 1023 5 2 1 1022
0 1024 7 1 2 1804 1931
0 1025 5 3 1 1024
0 1026 7 1 2 2638 2640
0 1027 5 1 1 1026
0 1028 7 2 2 2635 1027
0 1029 5 1 1 2643
0 1030 7 1 2 2634 2639
0 1031 5 1 1 1030
0 1032 7 1 2 2170 2207
0 1033 5 1 1 1032
0 1034 7 1 2 2255 1033
0 1035 5 1 1 1034
0 1036 7 1 2 2232 1035
0 1037 7 1 2 2540 1036
0 1038 7 1 2 2622 1037
0 1039 7 1 2 1031 1038
0 1040 7 1 2 1029 1039
0 1041 7 1 2 2550 1040
0 1042 7 1 2 2171 2624
0 1043 5 1 1 1042
0 1044 7 1 2 2174 2626
0 1045 5 1 1 1044
0 1046 7 2 2 1043 1045
0 1047 5 1 1 2645
0 1048 7 1 2 2233 2646
0 1049 5 1 1 1048
0 1050 7 1 2 2235 1047
0 1051 5 1 1 1050
0 1052 7 1 2 1049 1051
0 1053 7 1 2 1041 1052
0 1054 7 1 2 1017 1053
0 1055 7 1 2 1015 1054
0 1056 7 1 2 1011 1055
0 1057 7 1 2 975 1056
0 1058 5 1 1 1057
0 1059 7 1 2 2027 2438
0 1060 5 1 1 1059
0 1061 7 2 2 2024 1060
0 1062 5 2 1 2647
0 1063 7 1 2 2017 2649
0 1064 5 1 1 1063
0 1065 7 2 2 2014 1064
0 1066 5 2 1 2651
0 1067 7 1 2 2005 2653
0 1068 5 1 1 1067
0 1069 7 2 2 2002 1068
0 1070 5 2 1 2655
0 1071 7 1 2 1992 2657
0 1072 5 1 1 1071
0 1073 7 2 2 1989 1072
0 1074 5 2 1 2659
0 1075 7 1 2 1977 2661
0 1076 5 1 1 1075
0 1077 7 2 2 1974 1076
0 1078 5 2 1 2663
0 1079 7 1 2 1962 2665
0 1080 5 1 1 1079
0 1081 7 2 2 1959 1080
0 1082 5 2 1 2667
0 1083 7 1 2 1947 2669
0 1084 5 1 1 1083
0 1085 7 2 2 1944 1084
0 1086 5 2 1 2671
0 1087 7 1 2 2077 2673
0 1088 5 1 1 1087
0 1089 7 2 2 2074 1088
0 1090 5 2 1 2675
0 1091 7 1 2 2150 2677
0 1092 5 1 1 1091
0 1093 7 2 2 2147 1092
0 1094 5 2 1 2679
0 1095 7 1 2 2137 2681
0 1096 5 1 1 1095
0 1097 7 2 2 2134 1096
0 1098 5 2 1 2683
0 1099 7 1 2 2122 2685
0 1100 5 1 1 1099
0 1101 7 2 2 2119 1100
0 1102 5 2 1 2687
0 1103 7 1 2 2107 2688
0 1104 5 1 1 1103
0 1105 7 1 2 2109 2689
0 1106 5 1 1 1105
0 1107 7 4 2 1104 1106
0 1108 5 3 1 2691
0 1109 7 1 2 2080 2672
0 1110 5 1 1 1109
0 1111 7 1 2 2082 2674
0 1112 5 1 1 1111
0 1113 7 4 2 1110 1112
0 1114 5 3 1 2698
0 1115 7 1 2 2692 2699
0 1116 5 2 1 1115
0 1117 7 1 2 2695 2702
0 1118 5 1 1 1117
0 1119 7 2 2 2705 1118
0 1120 5 1 1 2707
0 1121 7 1 2 2181 2676
0 1122 5 1 1 1121
0 1123 7 1 2 2183 2678
0 1124 5 1 1 1123
0 1125 7 4 2 1122 1124
0 1126 5 3 1 2709
0 1127 7 1 2 2708 2710
0 1128 5 2 1 1127
0 1129 7 2 2 2706 2716
0 1130 5 1 1 2718
0 1131 7 1 2 2104 2690
0 1132 5 1 1 1131
0 1133 7 2 2 2101 1132
0 1134 5 2 1 2720
0 1135 7 1 2 2223 2721
0 1136 5 1 1 1135
0 1137 7 1 2 2225 2722
0 1138 5 1 1 1137
0 1139 7 3 2 1136 1138
0 1140 5 3 1 2724
0 1141 7 1 2 2711 2725
0 1142 5 2 1 1141
0 1143 7 1 2 2713 2727
0 1144 5 1 1 1143
0 1145 7 2 2 2730 1144
0 1146 5 1 1 2732
0 1147 7 1 2 2199 2680
0 1148 5 1 1 1147
0 1149 7 1 2 2197 2682
0 1150 5 1 1 1149
0 1151 7 4 2 1148 1150
0 1152 5 3 1 2734
0 1153 7 1 2 2733 2738
0 1154 5 2 1 1153
0 1155 7 1 2 1146 2735
0 1156 5 1 1 1155
0 1157 7 2 2 2741 1156
0 1158 5 1 1 2743
0 1159 7 1 2 1130 2744
0 1160 5 2 1 1159
0 1161 7 1 2 2250 2684
0 1162 5 1 1 1161
0 1163 7 1 2 2248 2686
0 1164 5 1 1 1163
0 1165 7 4 2 1162 1164
0 1166 5 3 1 2747
0 1167 7 1 2 2263 2668
0 1168 5 1 1 1167
0 1169 7 1 2 2261 2670
0 1170 5 1 1 1169
0 1171 7 4 2 1168 1170
0 1172 5 3 1 2754
0 1173 7 1 2 2751 2758
0 1174 5 2 1 1173
0 1175 7 1 2 2748 2755
0 1176 5 1 1 1175
0 1177 7 2 2 2761 1176
0 1178 5 1 1 2763
0 1179 7 1 2 2700 2764
0 1180 5 2 1 1179
0 1181 7 2 2 2762 2765
0 1182 5 1 1 2767
0 1183 7 1 2 1120 2714
0 1184 5 1 1 1183
0 1185 7 2 2 2717 1184
0 1186 5 1 1 2769
0 1187 7 1 2 1182 2770
0 1188 5 2 1 1187
0 1189 7 1 2 2287 2664
0 1190 5 1 1 1189
0 1191 7 1 2 2285 2666
0 1192 5 1 1 1191
0 1193 7 4 2 1190 1192
0 1194 5 3 1 2773
0 1195 7 1 2 2739 2777
0 1196 5 2 1 1195
0 1197 7 1 2 2736 2774
0 1198 5 1 1 1197
0 1199 7 2 2 2780 1198
0 1200 5 1 1 2782
0 1201 7 1 2 2759 2783
0 1202 5 2 1 1201
0 1203 7 2 2 2781 2784
0 1204 5 1 1 2786
0 1205 7 1 2 2703 1178
0 1206 5 1 1 1205
0 1207 7 2 2 2766 1206
0 1208 5 1 1 2788
0 1209 7 1 2 1204 2789
0 1210 5 2 1 1209
0 1211 7 1 2 2311 2660
0 1212 5 1 1 1211
0 1213 7 1 2 2309 2662
0 1214 5 1 1 1213
0 1215 7 4 2 1212 1214
0 1216 5 3 1 2792
0 1217 7 1 2 2712 2796
0 1218 5 2 1 1217
0 1219 7 1 2 2715 2793
0 1220 5 1 1 1219
0 1221 7 2 2 2799 1220
0 1222 5 1 1 2801
0 1223 7 1 2 2778 2802
0 1224 5 2 1 1223
0 1225 7 2 2 2800 2803
0 1226 5 1 1 2805
0 1227 7 1 2 2756 1200
0 1228 5 1 1 1227
0 1229 7 2 2 2785 1228
0 1230 5 1 1 2807
0 1231 7 1 2 1226 2808
0 1232 5 2 1 1231
0 1233 7 1 2 2335 2656
0 1234 5 1 1 1233
0 1235 7 1 2 2333 2658
0 1236 5 1 1 1235
0 1237 7 4 2 1234 1236
0 1238 5 3 1 2811
0 1239 7 1 2 2701 2815
0 1240 5 2 1 1239
0 1241 7 1 2 2704 2812
0 1242 5 1 1 1241
0 1243 7 2 2 2818 1242
0 1244 5 1 1 2820
0 1245 7 1 2 2797 2821
0 1246 5 2 1 1245
0 1247 7 2 2 2819 2822
0 1248 5 1 1 2824
0 1249 7 1 2 2775 1222
0 1250 5 1 1 1249
0 1251 7 2 2 2804 1250
0 1252 5 1 1 2826
0 1253 7 1 2 1248 2827
0 1254 5 2 1 1253
0 1255 7 1 2 2359 2652
0 1256 5 1 1 1255
0 1257 7 1 2 2357 2654
0 1258 5 1 1 1257
0 1259 7 5 2 1256 1258
0 1260 5 3 1 2830
0 1261 7 1 2 2760 2835
0 1262 5 2 1 1261
0 1263 7 1 2 2757 2831
0 1264 5 1 1 1263
0 1265 7 2 2 2838 1264
0 1266 5 1 1 2840
0 1267 7 1 2 2816 2841
0 1268 5 2 1 1267
0 1269 7 2 2 2839 2842
0 1270 5 1 1 2844
0 1271 7 1 2 2794 1244
0 1272 5 1 1 1271
0 1273 7 2 2 2823 1272
0 1274 5 1 1 2846
0 1275 7 1 2 1270 2847
0 1276 5 2 1 1275
0 1277 7 1 2 2384 2648
0 1278 5 1 1 1277
0 1279 7 1 2 2382 2650
0 1280 5 1 1 1279
0 1281 7 4 2 1278 1280
0 1282 5 3 1 2850
0 1283 7 1 2 2779 2854
0 1284 5 2 1 1283
0 1285 7 1 2 2776 2851
0 1286 5 1 1 1285
0 1287 7 2 2 2857 1286
0 1288 5 1 1 2859
0 1289 7 1 2 2836 2860
0 1290 5 2 1 1289
0 1291 7 2 2 2858 2861
0 1292 5 1 1 2863
0 1293 7 1 2 2813 1266
0 1294 5 1 1 1293
0 1295 7 2 2 2843 1294
0 1296 5 1 1 2865
0 1297 7 1 2 1292 2866
0 1298 5 2 1 1297
0 1299 7 1 2 2406 2441
0 1300 5 1 1 1299
0 1301 7 1 2 2408 2439
0 1302 5 1 1 1301
0 1303 7 3 2 1300 1302
0 1304 5 3 1 2869
0 1305 7 1 2 2798 2870
0 1306 5 2 1 1305
0 1307 7 1 2 2795 2872
0 1308 5 1 1 1307
0 1309 7 2 2 2875 1308
0 1310 5 1 1 2877
0 1311 7 1 2 2855 2878
0 1312 5 2 1 1311
0 1313 7 2 2 2876 2879
0 1314 5 1 1 2881
0 1315 7 1 2 2832 1288
0 1316 5 1 1 1315
0 1317 7 2 2 2862 1316
0 1318 5 1 1 2883
0 1319 7 1 2 1314 2884
0 1320 5 2 1 1319
0 1321 7 2 2 2817 2871
0 1322 5 2 1 2887
0 1323 7 1 2 2852 1310
0 1324 5 1 1 1323
0 1325 7 2 2 2880 1324
0 1326 5 1 1 2891
0 1327 7 1 2 2888 2892
0 1328 5 2 1 1327
0 1329 7 1 2 2889 1326
0 1330 5 1 1 1329
0 1331 7 2 2 2893 1330
0 1332 5 1 1 2895
0 1333 7 1 2 2814 2873
0 1334 5 1 1 1333
0 1335 7 2 2 2890 1334
0 1336 5 2 1 2897
0 1337 7 1 2 2833 2899
0 1338 5 1 1 1337
0 1339 7 2 2 2448 1338
0 1340 5 1 1 2901
0 1341 7 1 2 2896 2902
0 1342 5 2 1 1341
0 1343 7 2 2 2894 2903
0 1344 5 1 1 2905
0 1345 7 1 2 2882 1318
0 1346 5 1 1 1345
0 1347 7 2 2 2885 1346
0 1348 5 1 1 2907
0 1349 7 1 2 1344 2908
0 1350 5 2 1 1349
0 1351 7 2 2 2886 2909
0 1352 5 1 1 2911
0 1353 7 1 2 2864 1296
0 1354 5 1 1 1353
0 1355 7 2 2 2867 1354
0 1356 5 1 1 2913
0 1357 7 1 2 1352 2914
0 1358 5 2 1 1357
0 1359 7 2 2 2868 2915
0 1360 5 1 1 2917
0 1361 7 1 2 2845 1274
0 1362 5 1 1 1361
0 1363 7 2 2 2848 1362
0 1364 5 1 1 2919
0 1365 7 1 2 1360 2920
0 1366 5 2 1 1365
0 1367 7 2 2 2849 2921
0 1368 5 1 1 2923
0 1369 7 1 2 2825 1252
0 1370 5 1 1 1369
0 1371 7 2 2 2828 1370
0 1372 5 1 1 2925
0 1373 7 1 2 1368 2926
0 1374 5 2 1 1373
0 1375 7 2 2 2829 2927
0 1376 5 1 1 2929
0 1377 7 1 2 2806 1230
0 1378 5 1 1 1377
0 1379 7 2 2 2809 1378
0 1380 5 1 1 2931
0 1381 7 1 2 1376 2932
0 1382 5 2 1 1381
0 1383 7 2 2 2810 2933
0 1384 5 1 1 2935
0 1385 7 1 2 2787 1208
0 1386 5 1 1 1385
0 1387 7 2 2 2790 1386
0 1388 5 1 1 2937
0 1389 7 1 2 1384 2938
0 1390 5 2 1 1389
0 1391 7 2 2 2791 2939
0 1392 5 1 1 2941
0 1393 7 1 2 2768 1186
0 1394 5 1 1 1393
0 1395 7 2 2 2771 1394
0 1396 5 1 1 2943
0 1397 7 1 2 1392 2944
0 1398 5 2 1 1397
0 1399 7 2 2 2772 2945
0 1400 5 1 1 2947
0 1401 7 1 2 2719 1158
0 1402 5 1 1 1401
0 1403 7 2 2 2745 1402
0 1404 5 1 1 2949
0 1405 7 1 2 1400 2950
0 1406 5 2 1 1405
0 1407 7 2 2 2746 2951
0 1408 5 1 1 2953
0 1409 7 2 2 2731 2742
0 1410 5 1 1 2955
0 1411 7 1 2 2217 2723
0 1412 5 1 1 1411
0 1413 7 2 2 2220 1412
0 1414 5 2 1 2957
0 1415 7 1 2 2530 2958
0 1416 5 1 1 1415
0 1417 7 1 2 2532 2959
0 1418 5 1 1 1417
0 1419 7 4 2 1416 1418
0 1420 5 3 1 2961
0 1421 7 1 2 2740 2962
0 1422 5 2 1 1421
0 1423 7 1 2 2737 2965
0 1424 5 1 1 1423
0 1425 7 2 2 2968 1424
0 1426 5 1 1 2970
0 1427 7 1 2 2752 2971
0 1428 5 2 1 1427
0 1429 7 1 2 2749 1426
0 1430 5 1 1 1429
0 1431 7 2 2 2972 1430
0 1432 5 1 1 2974
0 1433 7 1 2 1410 2975
0 1434 5 2 1 1433
0 1435 7 1 2 2956 1432
0 1436 5 1 1 1435
0 1437 7 2 2 2976 1436
0 1438 5 1 1 2978
0 1439 7 1 2 1408 2979
0 1440 5 2 1 1439
0 1441 7 1 2 2954 1438
0 1442 5 1 1 1441
0 1443 7 2 2 2980 1442
0 1444 5 1 1 2982
0 1445 7 1 2 1932 2983
0 1446 5 1 1 1445
0 1447 7 1 2 2524 2960
0 1448 5 1 1 1447
0 1449 7 2 2 2527 1448
0 1450 5 2 1 2984
0 1451 7 1 2 2606 2986
0 1452 5 1 1 1451
0 1453 7 2 2 2609 1452
0 1454 5 2 1 2988
0 1455 7 1 2 2641 2990
0 1456 5 1 1 1455
0 1457 7 4 2 2636 1456
0 1458 5 2 1 2992
0 1459 7 1 2 2612 2987
0 1460 5 1 1 1459
0 1461 7 1 2 2614 2985
0 1462 5 1 1 1461
0 1463 7 3 2 1460 1462
0 1464 5 2 1 2998
0 1465 7 1 2 2996 3001
0 1466 5 2 1 1465
0 1467 7 1 2 2993 2999
0 1468 5 1 1 1467
0 1469 7 3 2 3003 1468
0 1470 5 2 1 3005
0 1471 7 1 2 2963 3006
0 1472 5 2 1 1471
0 1473 7 2 2 3004 3010
0 1474 5 1 1 3012
0 1475 7 2 2 2637 2642
0 1476 5 1 1 3014
0 1477 7 1 2 2991 3015
0 1478 5 1 1 1477
0 1479 7 1 2 2989 1476
0 1480 5 1 1 1479
0 1481 7 3 2 1478 1480
0 1482 5 2 1 3016
0 1483 7 1 2 3017 3007
0 1484 5 1 1 1483
0 1485 7 1 2 3019 3008
0 1486 5 1 1 1485
0 1487 7 2 2 1484 1486
0 1488 5 1 1 3021
0 1489 7 1 2 3013 3022
0 1490 7 1 2 2964 2997
0 1491 5 2 1 1490
0 1492 7 1 2 2966 2994
0 1493 5 1 1 1492
0 1494 7 2 2 3023 1493
0 1495 5 1 1 3025
0 1496 7 1 2 2726 3026
0 1497 5 2 1 1496
0 1498 7 2 2 3024 3027
0 1499 5 1 1 3029
0 1500 7 2 2 2969 2973
0 1501 5 1 1 3031
0 1502 7 1 2 2753 3002
0 1503 5 2 1 1502
0 1504 7 1 2 2750 3000
0 1505 5 1 1 1504
0 1506 7 2 2 3033 1505
0 1507 5 1 1 3035
0 1508 7 1 2 2693 3036
0 1509 5 1 1 1508
0 1510 7 1 2 2696 1507
0 1511 5 1 1 1510
0 1512 7 2 2 1509 1511
0 1513 5 1 1 3037
0 1514 7 1 2 1501 3038
0 1515 5 2 1 1514
0 1516 7 1 2 3032 1513
0 1517 5 1 1 1516
0 1518 7 1 2 3039 1517
0 1519 5 1 1 1518
0 1520 7 1 2 3030 1519
0 1521 7 1 2 1489 1520
0 1522 7 2 2 2728 1495
0 1523 5 1 1 3041
0 1524 7 2 2 2967 3009
0 1525 5 1 1 3043
0 1526 7 1 2 3042 3044
0 1527 7 1 2 3040 1526
0 1528 7 2 2 2697 3018
0 1529 5 1 1 3045
0 1530 7 1 2 2644 3034
0 1531 7 1 2 2995 1530
0 1532 7 1 2 3046 1531
0 1533 7 1 2 2977 1532
0 1534 7 1 2 2981 1533
0 1535 7 1 2 1527 1534
0 1536 7 1 2 1521 1535
0 1537 7 1 2 1446 1536
0 1538 7 1 2 1929 1444
0 1539 5 1 1 1538
0 1540 7 1 2 2942 1396
0 1541 5 1 1 1540
0 1542 7 2 2 2946 1541
0 1543 5 1 1 3047
0 1544 7 1 2 2518 3048
0 1545 5 1 1 1544
0 1546 7 1 2 2521 1543
0 1547 5 1 1 1546
0 1548 7 1 2 2936 1388
0 1549 5 1 1 1548
0 1550 7 2 2 2940 1549
0 1551 5 1 1 3049
0 1552 7 1 2 2930 1380
0 1553 5 1 1 1552
0 1554 7 2 2 2934 1553
0 1555 5 1 1 3051
0 1556 7 1 2 2098 3052
0 1557 5 1 1 1556
0 1558 7 1 2 2095 1555
0 1559 5 1 1 1558
0 1560 7 1 2 2924 1372
0 1561 5 1 1 1560
0 1562 7 2 2 2928 1561
0 1563 5 1 1 3053
0 1564 7 1 2 2918 1364
0 1565 5 1 1 1564
0 1566 7 2 2 2922 1565
0 1567 5 1 1 3055
0 1568 7 1 2 2131 3056
0 1569 5 1 1 1568
0 1570 7 1 2 2128 1567
0 1571 5 1 1 1570
0 1572 7 1 2 2912 1356
0 1573 5 1 1 1572
0 1574 7 2 2 2916 1573
0 1575 5 1 1 3057
0 1576 7 1 2 2906 1348
0 1577 5 1 1 1576
0 1578 7 2 2 2910 1577
0 1579 5 1 1 3059
0 1580 7 1 2 2071 3060
0 1581 5 1 1 1580
0 1582 7 1 2 2068 1579
0 1583 5 1 1 1582
0 1584 7 1 2 1332 1340
0 1585 5 1 1 1584
0 1586 7 2 2 2904 1585
0 1587 5 1 1 3061
0 1588 7 1 2 1941 3062
0 1589 5 1 1 1588
0 1590 7 1 2 1938 1587
0 1591 5 1 1 1590
0 1592 7 2 2 2449 2834
0 1593 5 2 1 3063
0 1594 7 1 2 2898 3065
0 1595 5 1 1 1594
0 1596 7 1 2 2900 3064
0 1597 5 1 1 1596
0 1598 7 2 2 1595 1597
0 1599 5 1 1 3067
0 1600 7 1 2 1956 1599
0 1601 5 1 1 1600
0 1602 7 1 2 1953 3068
0 1603 5 1 1 1602
0 1604 7 1 2 2444 2837
0 1605 5 1 1 1604
0 1606 7 2 2 3066 1605
0 1607 5 1 1 3069
0 1608 7 1 2 1971 1607
0 1609 5 1 1 1608
0 1610 7 1 2 1968 3070
0 1611 5 1 1 1610
0 1612 7 1 2 1986 2856
0 1613 5 1 1 1612
0 1614 7 1 2 1983 2853
0 1615 5 1 1 1614
0 1616 7 1 2 2597 2874
0 1617 5 1 1 1616
0 1618 7 1 2 2595 1617
0 1619 7 1 2 1615 1618
0 1620 5 1 1 1619
0 1621 7 1 2 1613 1620
0 1622 5 1 1 1621
0 1623 7 1 2 1611 1622
0 1624 5 1 1 1623
0 1625 7 1 2 1609 1624
0 1626 5 1 1 1625
0 1627 7 1 2 1603 1626
0 1628 5 1 1 1627
0 1629 7 1 2 1601 1628
0 1630 5 1 1 1629
0 1631 7 1 2 1591 1630
0 1632 5 1 1 1631
0 1633 7 1 2 1589 1632
0 1634 5 1 1 1633
0 1635 7 1 2 1583 1634
0 1636 5 1 1 1635
0 1637 7 2 2 1581 1636
0 1638 5 1 1 3071
0 1639 7 1 2 3058 1638
0 1640 5 1 1 1639
0 1641 7 1 2 1575 3072
0 1642 5 1 1 1641
0 1643 7 1 2 2144 1642
0 1644 5 1 1 1643
0 1645 7 1 2 1640 1644
0 1646 5 1 1 1645
0 1647 7 1 2 1571 1646
0 1648 5 1 1 1647
0 1649 7 2 2 1569 1648
0 1650 5 1 1 3073
0 1651 7 1 2 3054 1650
0 1652 5 1 1 1651
0 1653 7 1 2 1563 3074
0 1654 5 1 1 1653
0 1655 7 1 2 2116 1654
0 1656 5 1 1 1655
0 1657 7 1 2 1652 1656
0 1658 5 1 1 1657
0 1659 7 1 2 1559 1658
0 1660 5 1 1 1659
0 1661 7 2 2 1557 1660
0 1662 5 1 1 3075
0 1663 7 1 2 3050 1662
0 1664 5 1 1 1663
0 1665 7 1 2 1551 3076
0 1666 5 1 1 1665
0 1667 7 1 2 2214 1666
0 1668 5 1 1 1667
0 1669 7 1 2 1664 1668
0 1670 5 1 1 1669
0 1671 7 1 2 1547 1670
0 1672 5 1 1 1671
0 1673 7 1 2 1545 1672
0 1674 5 1 1 1673
0 1675 7 1 2 2948 1404
0 1676 5 1 1 1675
0 1677 7 2 2 2952 1676
0 1678 5 1 1 3077
0 1679 7 1 2 2565 1678
0 1680 5 1 1 1679
0 1681 7 1 2 1674 1680
0 1682 5 1 1 1681
0 1683 7 1 2 2562 3078
0 1684 5 1 1 1683
0 1685 7 1 2 1682 1684
0 1686 5 1 1 1685
0 1687 7 1 2 1539 1686
0 1688 5 1 1 1687
0 1689 7 1 2 3011 1525
0 1690 7 1 2 1499 1689
0 1691 5 1 1 1690
0 1692 7 1 2 2694 3020
0 1693 5 1 1 1692
0 1694 7 1 2 2729 1693
0 1695 5 1 1 1694
0 1696 7 1 2 1695 1529
0 1697 7 1 2 3028 1696
0 1698 7 1 2 1523 1697
0 1699 5 1 1 1698
0 1700 7 1 2 1474 1488
0 1701 5 1 1 1700
0 1702 7 1 2 1699 1701
0 1703 7 1 2 1691 1702
0 1704 7 1 2 1688 1703
0 1705 7 1 2 1537 1704
0 1706 5 1 1 1705
0 1707 7 1 2 1058 1706
3 3999 5 0 1 1707
