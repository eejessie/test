1 0 0 8 0
2 32 1 0
2 1983 1 0
2 1984 1 0
2 1985 1 0
2 1986 1 0
2 1987 1 0
2 1988 1 0
2 1989 1 0
1 1 0 10 0
2 1990 1 1
2 1991 1 1
2 1992 1 1
2 1993 1 1
2 1994 1 1
2 1995 1 1
2 1996 1 1
2 1997 1 1
2 1998 1 1
2 1999 1 1
1 2 0 10 0
2 2000 1 2
2 2001 1 2
2 2002 1 2
2 2003 1 2
2 2004 1 2
2 2005 1 2
2 2006 1 2
2 2007 1 2
2 2008 1 2
2 2009 1 2
1 3 0 11 0
2 2010 1 3
2 2011 1 3
2 2012 1 3
2 2013 1 3
2 2014 1 3
2 2015 1 3
2 2016 1 3
2 2017 1 3
2 2018 1 3
2 2019 1 3
2 2020 1 3
1 4 0 10 0
2 2021 1 4
2 2022 1 4
2 2023 1 4
2 2024 1 4
2 2025 1 4
2 2026 1 4
2 2027 1 4
2 2028 1 4
2 2029 1 4
2 2030 1 4
1 5 0 11 0
2 2031 1 5
2 2032 1 5
2 2033 1 5
2 2034 1 5
2 2035 1 5
2 2036 1 5
2 2037 1 5
2 2038 1 5
2 2039 1 5
2 2040 1 5
2 2041 1 5
1 6 0 10 0
2 2042 1 6
2 2043 1 6
2 2044 1 6
2 2045 1 6
2 2046 1 6
2 2047 1 6
2 2048 1 6
2 2049 1 6
2 2050 1 6
2 2051 1 6
1 7 0 10 0
2 2052 1 7
2 2053 1 7
2 2054 1 7
2 2055 1 7
2 2056 1 7
2 2057 1 7
2 2058 1 7
2 2059 1 7
2 2060 1 7
2 2061 1 7
1 8 0 10 0
2 2062 1 8
2 2063 1 8
2 2064 1 8
2 2065 1 8
2 2066 1 8
2 2067 1 8
2 2068 1 8
2 2069 1 8
2 2070 1 8
2 2071 1 8
1 9 0 10 0
2 2072 1 9
2 2073 1 9
2 2074 1 9
2 2075 1 9
2 2076 1 9
2 2077 1 9
2 2078 1 9
2 2079 1 9
2 2080 1 9
2 2081 1 9
1 10 0 11 0
2 2082 1 10
2 2083 1 10
2 2084 1 10
2 2085 1 10
2 2086 1 10
2 2087 1 10
2 2088 1 10
2 2089 1 10
2 2090 1 10
2 2091 1 10
2 2092 1 10
1 11 0 10 0
2 2093 1 11
2 2094 1 11
2 2095 1 11
2 2096 1 11
2 2097 1 11
2 2098 1 11
2 2099 1 11
2 2100 1 11
2 2101 1 11
2 2102 1 11
1 12 0 10 0
2 2103 1 12
2 2104 1 12
2 2105 1 12
2 2106 1 12
2 2107 1 12
2 2108 1 12
2 2109 1 12
2 2110 1 12
2 2111 1 12
2 2112 1 12
1 13 0 10 0
2 2113 1 13
2 2114 1 13
2 2115 1 13
2 2116 1 13
2 2117 1 13
2 2118 1 13
2 2119 1 13
2 2120 1 13
2 2121 1 13
2 2122 1 13
1 14 0 10 0
2 2123 1 14
2 2124 1 14
2 2125 1 14
2 2126 1 14
2 2127 1 14
2 2128 1 14
2 2129 1 14
2 2130 1 14
2 2131 1 14
2 2132 1 14
1 15 0 10 0
2 2133 1 15
2 2134 1 15
2 2135 1 15
2 2136 1 15
2 2137 1 15
2 2138 1 15
2 2139 1 15
2 2140 1 15
2 2141 1 15
2 2142 1 15
1 16 0 3 0
2 2143 1 16
2 2144 1 16
2 2145 1 16
1 17 0 3 0
2 2146 1 17
2 2147 1 17
2 2148 1 17
1 18 0 3 0
2 2149 1 18
2 2150 1 18
2 2151 1 18
1 19 0 3 0
2 2152 1 19
2 2153 1 19
2 2154 1 19
1 20 0 3 0
2 2155 1 20
2 2156 1 20
2 2157 1 20
1 21 0 3 0
2 2158 1 21
2 2159 1 21
2 2160 1 21
1 22 0 3 0
2 2161 1 22
2 2162 1 22
2 2163 1 22
1 23 0 3 0
2 2164 1 23
2 2165 1 23
2 2166 1 23
1 24 0 3 0
2 2167 1 24
2 2168 1 24
2 2169 1 24
1 25 0 3 0
2 2170 1 25
2 2171 1 25
2 2172 1 25
1 26 0 3 0
2 2173 1 26
2 2174 1 26
2 2175 1 26
1 27 0 3 0
2 2176 1 27
2 2177 1 27
2 2178 1 27
1 28 0 4 0
2 2179 1 28
2 2180 1 28
2 2181 1 28
2 2182 1 28
1 29 0 3 0
2 2183 1 29
2 2184 1 29
2 2185 1 29
1 30 0 4 0
2 2186 1 30
2 2187 1 30
2 2188 1 30
2 2189 1 30
1 31 0 4 0
2 2190 1 31
2 2191 1 31
2 2192 1 31
2 2193 1 31
2 2194 1 33
2 2195 1 33
2 2196 1 34
2 2197 1 34
2 2198 1 35
2 2199 1 35
2 2200 1 36
2 2201 1 36
2 2202 1 37
2 2203 1 37
2 2204 1 38
2 2205 1 38
2 2206 1 39
2 2207 1 39
2 2208 1 40
2 2209 1 40
2 2210 1 41
2 2211 1 41
2 2212 1 42
2 2213 1 42
2 2214 1 43
2 2215 1 43
2 2216 1 44
2 2217 1 44
2 2218 1 45
2 2219 1 45
2 2220 1 46
2 2221 1 46
2 2222 1 47
2 2223 1 47
2 2224 1 48
2 2225 1 48
2 2226 1 48
2 2227 1 49
2 2228 1 49
2 2229 1 49
2 2230 1 50
2 2231 1 50
2 2232 1 50
2 2233 1 51
2 2234 1 51
2 2235 1 51
2 2236 1 52
2 2237 1 52
2 2238 1 52
2 2239 1 53
2 2240 1 53
2 2241 1 53
2 2242 1 54
2 2243 1 54
2 2244 1 54
2 2245 1 55
2 2246 1 55
2 2247 1 55
2 2248 1 56
2 2249 1 56
2 2250 1 56
2 2251 1 57
2 2252 1 57
2 2253 1 57
2 2254 1 58
2 2255 1 58
2 2256 1 58
2 2257 1 59
2 2258 1 59
2 2259 1 59
2 2260 1 60
2 2261 1 60
2 2262 1 60
2 2263 1 60
2 2264 1 61
2 2265 1 61
2 2266 1 61
2 2267 1 62
2 2268 1 62
2 2269 1 63
2 2270 1 63
2 2271 1 64
2 2272 1 64
2 2273 1 66
2 2274 1 66
2 2275 1 66
2 2276 1 68
2 2277 1 68
2 2278 1 74
2 2279 1 74
2 2280 1 76
2 2281 1 76
2 2282 1 81
2 2283 1 81
2 2284 1 84
2 2285 1 84
2 2286 1 87
2 2287 1 87
2 2288 1 89
2 2289 1 89
2 2290 1 90
2 2291 1 90
2 2292 1 95
2 2293 1 95
2 2294 1 98
2 2295 1 98
2 2296 1 103
2 2297 1 103
2 2298 1 104
2 2299 1 104
2 2300 1 105
2 2301 1 105
2 2302 1 108
2 2303 1 108
2 2304 1 111
2 2305 1 111
2 2306 1 113
2 2307 1 113
2 2308 1 114
2 2309 1 114
2 2310 1 119
2 2311 1 119
2 2312 1 122
2 2313 1 122
2 2314 1 127
2 2315 1 127
2 2316 1 127
2 2317 1 129
2 2318 1 129
2 2319 1 132
2 2320 1 132
2 2321 1 135
2 2322 1 135
2 2323 1 137
2 2324 1 137
2 2325 1 138
2 2326 1 138
2 2327 1 143
2 2328 1 143
2 2329 1 146
2 2330 1 146
2 2331 1 151
2 2332 1 151
2 2333 1 151
2 2334 1 153
2 2335 1 153
2 2336 1 156
2 2337 1 156
2 2338 1 159
2 2339 1 159
2 2340 1 161
2 2341 1 161
2 2342 1 162
2 2343 1 162
2 2344 1 167
2 2345 1 167
2 2346 1 170
2 2347 1 170
2 2348 1 175
2 2349 1 175
2 2350 1 175
2 2351 1 177
2 2352 1 177
2 2353 1 180
2 2354 1 180
2 2355 1 183
2 2356 1 183
2 2357 1 185
2 2358 1 185
2 2359 1 186
2 2360 1 186
2 2361 1 191
2 2362 1 191
2 2363 1 194
2 2364 1 194
2 2365 1 199
2 2366 1 199
2 2367 1 199
2 2368 1 201
2 2369 1 201
2 2370 1 204
2 2371 1 204
2 2372 1 207
2 2373 1 207
2 2374 1 209
2 2375 1 209
2 2376 1 210
2 2377 1 210
2 2378 1 215
2 2379 1 215
2 2380 1 218
2 2381 1 218
2 2382 1 223
2 2383 1 223
2 2384 1 223
2 2385 1 225
2 2386 1 225
2 2387 1 228
2 2388 1 228
2 2389 1 231
2 2390 1 231
2 2391 1 233
2 2392 1 233
2 2393 1 234
2 2394 1 234
2 2395 1 239
2 2396 1 239
2 2397 1 242
2 2398 1 242
2 2399 1 247
2 2400 1 247
2 2401 1 247
2 2402 1 249
2 2403 1 249
2 2404 1 252
2 2405 1 252
2 2406 1 255
2 2407 1 255
2 2408 1 257
2 2409 1 257
2 2410 1 258
2 2411 1 258
2 2412 1 263
2 2413 1 263
2 2414 1 266
2 2415 1 266
2 2416 1 271
2 2417 1 271
2 2418 1 271
2 2419 1 273
2 2420 1 273
2 2421 1 276
2 2422 1 276
2 2423 1 279
2 2424 1 279
2 2425 1 281
2 2426 1 281
2 2427 1 282
2 2428 1 282
2 2429 1 287
2 2430 1 287
2 2431 1 290
2 2432 1 290
2 2433 1 295
2 2434 1 295
2 2435 1 295
2 2436 1 297
2 2437 1 297
2 2438 1 300
2 2439 1 300
2 2440 1 303
2 2441 1 303
2 2442 1 305
2 2443 1 305
2 2444 1 306
2 2445 1 306
2 2446 1 311
2 2447 1 311
2 2448 1 314
2 2449 1 314
2 2450 1 319
2 2451 1 319
2 2452 1 319
2 2453 1 321
2 2454 1 321
2 2455 1 324
2 2456 1 324
2 2457 1 327
2 2458 1 327
2 2459 1 329
2 2460 1 329
2 2461 1 330
2 2462 1 330
2 2463 1 335
2 2464 1 335
2 2465 1 338
2 2466 1 338
2 2467 1 343
2 2468 1 343
2 2469 1 343
2 2470 1 345
2 2471 1 345
2 2472 1 348
2 2473 1 348
2 2474 1 351
2 2475 1 351
2 2476 1 353
2 2477 1 353
2 2478 1 354
2 2479 1 354
2 2480 1 359
2 2481 1 359
2 2482 1 362
2 2483 1 362
2 2484 1 367
2 2485 1 367
2 2486 1 367
2 2487 1 369
2 2488 1 369
2 2489 1 372
2 2490 1 372
2 2491 1 375
2 2492 1 375
2 2493 1 377
2 2494 1 377
2 2495 1 378
2 2496 1 378
2 2497 1 383
2 2498 1 383
2 2499 1 386
2 2500 1 386
2 2501 1 391
2 2502 1 391
2 2503 1 391
2 2504 1 393
2 2505 1 393
2 2506 1 396
2 2507 1 396
2 2508 1 399
2 2509 1 399
2 2510 1 401
2 2511 1 401
2 2512 1 402
2 2513 1 402
2 2514 1 407
2 2515 1 407
2 2516 1 410
2 2517 1 410
2 2518 1 415
2 2519 1 415
2 2520 1 415
2 2521 1 417
2 2522 1 417
2 2523 1 420
2 2524 1 420
2 2525 1 423
2 2526 1 423
2 2527 1 425
2 2528 1 425
2 2529 1 426
2 2530 1 426
2 2531 1 431
2 2532 1 431
2 2533 1 434
2 2534 1 434
2 2535 1 439
2 2536 1 439
2 2537 1 439
2 2538 1 441
2 2539 1 441
2 2540 1 444
2 2541 1 444
2 2542 1 447
2 2543 1 447
2 2544 1 449
2 2545 1 449
2 2546 1 450
2 2547 1 450
2 2548 1 455
2 2549 1 455
2 2550 1 458
2 2551 1 458
2 2552 1 463
2 2553 1 463
2 2554 1 463
2 2555 1 465
2 2556 1 465
2 2557 1 468
2 2558 1 468
2 2559 1 471
2 2560 1 471
2 2561 1 473
2 2562 1 473
2 2563 1 474
2 2564 1 474
2 2565 1 479
2 2566 1 479
2 2567 1 482
2 2568 1 482
2 2569 1 487
2 2570 1 487
2 2571 1 487
2 2572 1 489
2 2573 1 489
2 2574 1 492
2 2575 1 492
2 2576 1 495
2 2577 1 495
2 2578 1 497
2 2579 1 497
2 2580 1 498
2 2581 1 498
2 2582 1 503
2 2583 1 503
2 2584 1 506
2 2585 1 506
2 2586 1 511
2 2587 1 511
2 2588 1 511
2 2589 1 513
2 2590 1 513
2 2591 1 516
2 2592 1 516
2 2593 1 519
2 2594 1 519
2 2595 1 521
2 2596 1 521
2 2597 1 522
2 2598 1 522
2 2599 1 527
2 2600 1 527
2 2601 1 530
2 2602 1 530
2 2603 1 535
2 2604 1 535
2 2605 1 535
2 2606 1 537
2 2607 1 537
2 2608 1 540
2 2609 1 540
2 2610 1 543
2 2611 1 543
2 2612 1 545
2 2613 1 545
2 2614 1 546
2 2615 1 546
2 2616 1 551
2 2617 1 551
2 2618 1 554
2 2619 1 554
2 2620 1 559
2 2621 1 559
2 2622 1 559
2 2623 1 561
2 2624 1 561
2 2625 1 564
2 2626 1 564
2 2627 1 567
2 2628 1 567
2 2629 1 569
2 2630 1 569
2 2631 1 570
2 2632 1 570
2 2633 1 575
2 2634 1 575
2 2635 1 578
2 2636 1 578
2 2637 1 583
2 2638 1 583
2 2639 1 583
2 2640 1 585
2 2641 1 585
2 2642 1 588
2 2643 1 588
2 2644 1 591
2 2645 1 591
2 2646 1 593
2 2647 1 593
2 2648 1 594
2 2649 1 594
2 2650 1 599
2 2651 1 599
2 2652 1 602
2 2653 1 602
2 2654 1 607
2 2655 1 607
2 2656 1 607
2 2657 1 609
2 2658 1 609
2 2659 1 612
2 2660 1 612
2 2661 1 615
2 2662 1 615
2 2663 1 617
2 2664 1 617
2 2665 1 618
2 2666 1 618
2 2667 1 623
2 2668 1 623
2 2669 1 626
2 2670 1 626
2 2671 1 631
2 2672 1 631
2 2673 1 631
2 2674 1 633
2 2675 1 633
2 2676 1 636
2 2677 1 636
2 2678 1 639
2 2679 1 639
2 2680 1 641
2 2681 1 641
2 2682 1 642
2 2683 1 642
2 2684 1 647
2 2685 1 647
2 2686 1 650
2 2687 1 650
2 2688 1 655
2 2689 1 655
2 2690 1 655
2 2691 1 657
2 2692 1 657
2 2693 1 660
2 2694 1 660
2 2695 1 663
2 2696 1 663
2 2697 1 665
2 2698 1 665
2 2699 1 666
2 2700 1 666
2 2701 1 671
2 2702 1 671
2 2703 1 674
2 2704 1 674
2 2705 1 679
2 2706 1 679
2 2707 1 679
2 2708 1 681
2 2709 1 681
2 2710 1 686
2 2711 1 686
2 2712 1 687
2 2713 1 687
2 2714 1 687
2 2715 1 688
2 2716 1 688
2 2717 1 689
2 2718 1 689
2 2719 1 690
2 2720 1 690
2 2721 1 695
2 2722 1 695
2 2723 1 698
2 2724 1 698
2 2725 1 703
2 2726 1 703
2 2727 1 703
2 2728 1 711
2 2729 1 711
2 2730 1 714
2 2731 1 714
2 2732 1 717
2 2733 1 717
2 2734 1 728
2 2735 1 728
2 2736 1 739
2 2737 1 739
2 2738 1 741
2 2739 1 741
2 2740 1 743
2 2741 1 743
2 2742 1 746
2 2743 1 746
2 2744 1 747
2 2745 1 747
2 2746 1 751
2 2747 1 751
2 2748 1 754
2 2749 1 754
2 2750 1 755
2 2751 1 755
2 2752 1 757
2 2753 1 757
2 2754 1 758
2 2755 1 758
2 2756 1 759
2 2757 1 759
2 2758 1 761
2 2759 1 761
2 2760 1 766
2 2761 1 766
2 2762 1 767
2 2763 1 767
2 2764 1 770
2 2765 1 770
2 2766 1 773
2 2767 1 773
2 2768 1 776
2 2769 1 776
2 2770 1 777
2 2771 1 777
2 2772 1 781
2 2773 1 781
2 2774 1 784
2 2775 1 784
2 2776 1 785
2 2777 1 785
2 2778 1 787
2 2779 1 787
2 2780 1 790
2 2781 1 790
2 2782 1 791
2 2783 1 791
2 2784 1 795
2 2785 1 795
2 2786 1 798
2 2787 1 798
2 2788 1 799
2 2789 1 799
2 2790 1 803
2 2791 1 803
2 2792 1 806
2 2793 1 806
2 2794 1 807
2 2795 1 807
2 2796 1 811
2 2797 1 811
2 2798 1 814
2 2799 1 814
2 2800 1 815
2 2801 1 815
2 2802 1 817
2 2803 1 817
2 2804 1 819
2 2805 1 819
2 2806 1 821
2 2807 1 821
2 2808 1 827
2 2809 1 827
2 2810 1 830
2 2811 1 830
2 2812 1 830
2 2813 1 833
2 2814 1 833
2 2815 1 836
2 2816 1 836
2 2817 1 837
2 2818 1 837
2 2819 1 841
2 2820 1 841
2 2821 1 844
2 2822 1 844
2 2823 1 845
2 2824 1 845
2 2825 1 849
2 2826 1 849
2 2827 1 852
2 2828 1 852
2 2829 1 853
2 2830 1 853
2 2831 1 857
2 2832 1 857
2 2833 1 860
2 2834 1 860
2 2835 1 861
2 2836 1 861
2 2837 1 863
2 2838 1 863
2 2839 1 865
2 2840 1 865
2 2841 1 867
2 2842 1 867
2 2843 1 868
2 2844 1 868
2 2845 1 869
2 2846 1 869
2 2847 1 870
2 2848 1 870
2 2849 1 872
2 2850 1 872
2 2851 1 873
2 2852 1 873
2 2853 1 877
2 2854 1 877
2 2855 1 880
2 2856 1 880
2 2857 1 881
2 2858 1 881
2 2859 1 885
2 2860 1 885
2 2861 1 888
2 2862 1 888
2 2863 1 889
2 2864 1 889
2 2865 1 893
2 2866 1 893
2 2867 1 896
2 2868 1 896
2 2869 1 897
2 2870 1 897
2 2871 1 901
2 2872 1 901
2 2873 1 904
2 2874 1 904
2 2875 1 905
2 2876 1 905
2 2877 1 909
2 2878 1 909
2 2879 1 912
2 2880 1 912
2 2881 1 913
2 2882 1 913
2 2883 1 917
2 2884 1 917
2 2885 1 920
2 2886 1 920
2 2887 1 921
2 2888 1 921
2 2889 1 925
2 2890 1 925
2 2891 1 928
2 2892 1 928
2 2893 1 929
2 2894 1 929
2 2895 1 931
2 2896 1 931
2 2897 1 934
2 2898 1 934
2 2899 1 937
2 2900 1 937
2 2901 1 941
2 2902 1 941
2 2903 1 944
2 2904 1 944
2 2905 1 945
2 2906 1 945
2 2907 1 949
2 2908 1 949
2 2909 1 952
2 2910 1 952
2 2911 1 953
2 2912 1 953
2 2913 1 955
2 2914 1 955
2 2915 1 958
2 2916 1 958
2 2917 1 959
2 2918 1 959
2 2919 1 961
2 2920 1 961
2 2921 1 967
2 2922 1 967
2 2923 1 970
2 2924 1 970
2 2925 1 973
2 2926 1 973
2 2927 1 976
2 2928 1 976
2 2929 1 979
2 2930 1 979
2 2931 1 983
2 2932 1 983
2 2933 1 986
2 2934 1 986
2 2935 1 987
2 2936 1 987
2 2937 1 991
2 2938 1 991
2 2939 1 994
2 2940 1 994
2 2941 1 995
2 2942 1 995
2 2943 1 997
2 2944 1 997
2 2945 1 1000
2 2946 1 1000
2 2947 1 1003
2 2948 1 1003
2 2949 1 1007
2 2950 1 1007
2 2951 1 1010
2 2952 1 1010
2 2953 1 1011
2 2954 1 1011
2 2955 1 1015
2 2956 1 1015
2 2957 1 1018
2 2958 1 1018
2 2959 1 1019
2 2960 1 1019
2 2961 1 1023
2 2962 1 1023
2 2963 1 1026
2 2964 1 1026
2 2965 1 1027
2 2966 1 1027
2 2967 1 1031
2 2968 1 1031
2 2969 1 1034
2 2970 1 1034
2 2971 1 1035
2 2972 1 1035
2 2973 1 1039
2 2974 1 1039
2 2975 1 1042
2 2976 1 1042
2 2977 1 1043
2 2978 1 1043
2 2979 1 1045
2 2980 1 1045
2 2981 1 1047
2 2982 1 1047
2 2983 1 1049
2 2984 1 1049
2 2985 1 1051
2 2986 1 1051
2 2987 1 1052
2 2988 1 1052
2 2989 1 1053
2 2990 1 1053
2 2991 1 1054
2 2992 1 1054
2 2993 1 1055
2 2994 1 1055
2 2995 1 1056
2 2996 1 1056
2 2997 1 1057
2 2998 1 1057
2 2999 1 1058
2 3000 1 1058
2 3001 1 1060
2 3002 1 1060
2 3003 1 1063
2 3004 1 1063
2 3005 1 1067
2 3006 1 1067
2 3007 1 1070
2 3008 1 1070
2 3009 1 1071
2 3010 1 1071
2 3011 1 1075
2 3012 1 1075
2 3013 1 1078
2 3014 1 1078
2 3015 1 1079
2 3016 1 1079
2 3017 1 1081
2 3018 1 1081
2 3019 1 1084
2 3020 1 1084
2 3021 1 1087
2 3022 1 1087
2 3023 1 1091
2 3024 1 1091
2 3025 1 1094
2 3026 1 1094
2 3027 1 1095
2 3028 1 1095
2 3029 1 1099
2 3030 1 1099
2 3031 1 1102
2 3032 1 1102
2 3033 1 1103
2 3034 1 1103
2 3035 1 1107
2 3036 1 1107
2 3037 1 1110
2 3038 1 1110
2 3039 1 1111
2 3040 1 1111
2 3041 1 1115
2 3042 1 1115
2 3043 1 1118
2 3044 1 1118
2 3045 1 1119
2 3046 1 1119
2 3047 1 1121
2 3048 1 1121
2 3049 1 1124
2 3050 1 1124
2 3051 1 1125
2 3052 1 1125
2 3053 1 1129
2 3054 1 1129
2 3055 1 1132
2 3056 1 1132
2 3057 1 1133
2 3058 1 1133
2 3059 1 1137
2 3060 1 1137
2 3061 1 1140
2 3062 1 1140
2 3063 1 1143
2 3064 1 1143
2 3065 1 1147
2 3066 1 1147
2 3067 1 1150
2 3068 1 1150
2 3069 1 1151
2 3070 1 1151
2 3071 1 1153
2 3072 1 1153
2 3073 1 1156
2 3074 1 1156
2 3075 1 1157
2 3076 1 1157
2 3077 1 1161
2 3078 1 1161
2 3079 1 1164
2 3080 1 1164
2 3081 1 1165
2 3082 1 1165
2 3083 1 1169
2 3084 1 1169
2 3085 1 1172
2 3086 1 1172
2 3087 1 1173
2 3088 1 1173
2 3089 1 1177
2 3090 1 1177
2 3091 1 1180
2 3092 1 1180
2 3093 1 1181
2 3094 1 1181
2 3095 1 1185
2 3096 1 1185
2 3097 1 1188
2 3098 1 1188
2 3099 1 1189
2 3100 1 1189
2 3101 1 1193
2 3102 1 1193
2 3103 1 1196
2 3104 1 1196
2 3105 1 1197
2 3106 1 1197
2 3107 1 1199
2 3108 1 1199
2 3109 1 1205
2 3110 1 1205
2 3111 1 1208
2 3112 1 1208
2 3113 1 1211
2 3114 1 1211
2 3115 1 1214
2 3116 1 1214
2 3117 1 1217
2 3118 1 1217
2 3119 1 1221
2 3120 1 1221
2 3121 1 1224
2 3122 1 1224
2 3123 1 1225
2 3124 1 1225
2 3125 1 1229
2 3126 1 1229
2 3127 1 1232
2 3128 1 1232
2 3129 1 1233
2 3130 1 1233
2 3131 1 1237
2 3132 1 1237
2 3133 1 1240
2 3134 1 1240
2 3135 1 1241
2 3136 1 1241
2 3137 1 1245
2 3138 1 1245
2 3139 1 1248
2 3140 1 1248
2 3141 1 1249
2 3142 1 1249
2 3143 1 1253
2 3144 1 1253
2 3145 1 1256
2 3146 1 1256
2 3147 1 1257
2 3148 1 1257
2 3149 1 1261
2 3150 1 1261
2 3151 1 1264
2 3152 1 1264
2 3153 1 1265
2 3154 1 1265
2 3155 1 1269
2 3156 1 1269
2 3157 1 1272
2 3158 1 1272
2 3159 1 1273
2 3160 1 1273
2 3161 1 1275
2 3162 1 1275
2 3163 1 1278
2 3164 1 1278
2 3165 1 1281
2 3166 1 1281
2 3167 1 1285
2 3168 1 1285
2 3169 1 1288
2 3170 1 1288
2 3171 1 1289
2 3172 1 1289
2 3173 1 1293
2 3174 1 1293
2 3175 1 1296
2 3176 1 1296
2 3177 1 1297
2 3178 1 1297
2 3179 1 1301
2 3180 1 1301
2 3181 1 1304
2 3182 1 1304
2 3183 1 1305
2 3184 1 1305
2 3185 1 1309
2 3186 1 1309
2 3187 1 1312
2 3188 1 1312
2 3189 1 1313
2 3190 1 1313
2 3191 1 1319
2 3192 1 1319
2 3193 1 1322
2 3194 1 1322
2 3195 1 1323
2 3196 1 1323
2 3197 1 1327
2 3198 1 1327
2 3199 1 1330
2 3200 1 1330
2 3201 1 1331
2 3202 1 1331
2 3203 1 1335
2 3204 1 1335
2 3205 1 1338
2 3206 1 1338
2 3207 1 1339
2 3208 1 1339
2 3209 1 1343
2 3210 1 1343
2 3211 1 1346
2 3212 1 1346
2 3213 1 1347
2 3214 1 1347
2 3215 1 1349
2 3216 1 1349
2 3217 1 1352
2 3218 1 1352
2 3219 1 1355
2 3220 1 1355
2 3221 1 1359
2 3222 1 1359
2 3223 1 1362
2 3224 1 1362
2 3225 1 1363
2 3226 1 1363
2 3227 1 1367
2 3228 1 1367
2 3229 1 1370
2 3230 1 1370
2 3231 1 1373
2 3232 1 1373
2 3233 1 1375
2 3234 1 1375
2 3235 1 1377
2 3236 1 1377
2 3237 1 1379
2 3238 1 1379
2 3239 1 1381
2 3240 1 1381
2 3241 1 1383
2 3242 1 1383
2 3243 1 1385
2 3244 1 1385
2 3245 1 1386
2 3246 1 1386
2 3247 1 1387
2 3248 1 1387
2 3249 1 1387
2 3250 1 1390
2 3251 1 1390
2 3252 1 1393
2 3253 1 1393
2 3254 1 1401
2 3255 1 1401
2 3256 1 1404
2 3257 1 1404
2 3258 1 1405
2 3259 1 1405
2 3260 1 1409
2 3261 1 1409
2 3262 1 1412
2 3263 1 1412
2 3264 1 1415
2 3265 1 1415
2 3266 1 1417
2 3267 1 1417
2 3268 1 1419
2 3269 1 1419
2 3270 1 1421
2 3271 1 1421
2 3272 1 1422
2 3273 1 1422
2 3274 1 1424
2 3275 1 1424
2 3276 1 1425
2 3277 1 1425
2 3278 1 1429
2 3279 1 1429
2 3280 1 1432
2 3281 1 1432
2 3282 1 1433
2 3283 1 1433
2 3284 1 1437
2 3285 1 1437
2 3286 1 1440
2 3287 1 1440
2 3288 1 1441
2 3289 1 1441
2 3290 1 1445
2 3291 1 1445
2 3292 1 1448
2 3293 1 1448
2 3294 1 1449
2 3295 1 1449
2 3296 1 1453
2 3297 1 1453
2 3298 1 1456
2 3299 1 1456
2 3300 1 1457
2 3301 1 1457
2 3302 1 1461
2 3303 1 1461
2 3304 1 1464
2 3305 1 1464
2 3306 1 1465
2 3307 1 1465
2 3308 1 1469
2 3309 1 1469
2 3310 1 1472
2 3311 1 1472
2 3312 1 1473
2 3313 1 1473
2 3314 1 1477
2 3315 1 1477
2 3316 1 1480
2 3317 1 1480
2 3318 1 1481
2 3319 1 1481
2 3320 1 1485
2 3321 1 1485
2 3322 1 1488
2 3323 1 1488
2 3324 1 1489
2 3325 1 1489
2 3326 1 1493
2 3327 1 1493
2 3328 1 1496
2 3329 1 1496
2 3330 1 1497
2 3331 1 1497
2 3332 1 1501
2 3333 1 1501
2 3334 1 1504
2 3335 1 1504
2 3336 1 1505
2 3337 1 1505
2 3338 1 1509
2 3339 1 1509
2 3340 1 1512
2 3341 1 1512
2 3342 1 1513
2 3343 1 1513
2 3344 1 1515
2 3345 1 1515
2 3346 1 1520
2 3347 1 1520
2 3348 1 1523
2 3349 1 1523
2 3350 1 1526
2 3351 1 1526
2 3352 1 1529
2 3353 1 1529
2 3354 1 1532
2 3355 1 1532
2 3356 1 1532
2 3357 1 1533
2 3358 1 1533
2 3359 1 1535
2 3360 1 1535
2 3361 1 1537
2 3362 1 1537
2 3363 1 1539
2 3364 1 1539
2 3365 1 1540
2 3366 1 1540
2 3367 1 1545
2 3368 1 1545
2 3369 1 1548
2 3370 1 1548
2 3371 1 1548
2 3372 1 1550
2 3373 1 1550
2 3374 1 1550
2 3375 1 1550
2 3376 1 1553
2 3377 1 1553
2 3378 1 1556
2 3379 1 1556
2 3380 1 1556
2 3381 1 1556
2 3382 1 1558
2 3383 1 1558
2 3384 1 1558
2 3385 1 1561
2 3386 1 1561
2 3387 1 1564
2 3388 1 1564
2 3389 1 1564
2 3390 1 1564
2 3391 1 1566
2 3392 1 1566
2 3393 1 1566
2 3394 1 1566
2 3395 1 1569
2 3396 1 1569
2 3397 1 1572
2 3398 1 1572
2 3399 1 1572
2 3400 1 1574
2 3401 1 1574
2 3402 1 1574
2 3403 1 1577
2 3404 1 1577
2 3405 1 1580
2 3406 1 1580
2 3407 1 1580
2 3408 1 1581
2 3409 1 1581
2 3410 1 1582
2 3411 1 1582
2 3412 1 1583
2 3413 1 1583
2 3414 1 1583
2 3415 1 1583
2 3416 1 1586
2 3417 1 1586
2 3418 1 1589
2 3419 1 1589
2 3420 1 1589
2 3421 1 1591
2 3422 1 1591
2 3423 1 1591
2 3424 1 1591
2 3425 1 1594
2 3426 1 1594
2 3427 1 1597
2 3428 1 1597
2 3429 1 1597
2 3430 1 1599
2 3431 1 1599
2 3432 1 1599
2 3433 1 1599
2 3434 1 1602
2 3435 1 1602
2 3436 1 1605
2 3437 1 1605
2 3438 1 1605
2 3439 1 1607
2 3440 1 1607
2 3441 1 1607
2 3442 1 1607
2 3443 1 1610
2 3444 1 1610
2 3445 1 1613
2 3446 1 1613
2 3447 1 1613
2 3448 1 1613
2 3449 1 1615
2 3450 1 1615
2 3451 1 1615
2 3452 1 1615
2 3453 1 1618
2 3454 1 1618
2 3455 1 1621
2 3456 1 1621
2 3457 1 1621
2 3458 1 1621
2 3459 1 1623
2 3460 1 1623
2 3461 1 1623
2 3462 1 1623
2 3463 1 1626
2 3464 1 1626
2 3465 1 1629
2 3466 1 1629
2 3467 1 1629
2 3468 1 1629
2 3469 1 1631
2 3470 1 1631
2 3471 1 1631
2 3472 1 1634
2 3473 1 1634
2 3474 1 1637
2 3475 1 1637
2 3476 1 1637
2 3477 1 1639
2 3478 1 1639
2 3479 1 1639
2 3480 1 1639
2 3481 1 1642
2 3482 1 1642
2 3483 1 1645
2 3484 1 1645
2 3485 1 1647
2 3486 1 1647
2 3487 1 1648
2 3488 1 1648
2 3489 1 1652
2 3490 1 1652
2 3491 1 1655
2 3492 1 1655
2 3493 1 1655
2 3494 1 1658
2 3495 1 1658
2 3496 1 1658
2 3497 1 1662
2 3498 1 1662
2 3499 1 1664
2 3500 1 1664
2 3501 1 1666
2 3502 1 1666
2 3503 1 1667
2 3504 1 1667
2 3505 1 1670
2 3506 1 1670
2 3507 1 1671
2 3508 1 1671
2 3509 1 1674
2 3510 1 1674
2 3511 1 1675
2 3512 1 1675
2 3513 1 1678
2 3514 1 1678
2 3515 1 1679
2 3516 1 1679
2 3517 1 1682
2 3518 1 1682
2 3519 1 1682
2 3520 1 1688
2 3521 1 1688
2 3522 1 1690
2 3523 1 1690
2 3524 1 1696
2 3525 1 1696
2 3526 1 1697
2 3527 1 1697
2 3528 1 1700
2 3529 1 1700
2 3530 1 1701
2 3531 1 1701
2 3532 1 1703
2 3533 1 1703
2 3534 1 1703
2 3535 1 1704
2 3536 1 1704
2 3537 1 1707
2 3538 1 1707
2 3539 1 1707
2 3540 1 1711
2 3541 1 1711
2 3542 1 1714
2 3543 1 1714
2 3544 1 1714
2 3545 1 1715
2 3546 1 1715
2 3547 1 1716
2 3548 1 1716
2 3549 1 1719
2 3550 1 1719
2 3551 1 1720
2 3552 1 1720
2 3553 1 1722
2 3554 1 1722
2 3555 1 1723
2 3556 1 1723
2 3557 1 1726
2 3558 1 1726
2 3559 1 1728
2 3560 1 1728
2 3561 1 1730
2 3562 1 1730
2 3563 1 1731
2 3564 1 1731
2 3565 1 1734
2 3566 1 1734
2 3567 1 1735
2 3568 1 1735
2 3569 1 1738
2 3570 1 1738
2 3571 1 1739
2 3572 1 1739
2 3573 1 1742
2 3574 1 1742
2 3575 1 1743
2 3576 1 1743
2 3577 1 1746
2 3578 1 1746
2 3579 1 1747
2 3580 1 1747
2 3581 1 1750
2 3582 1 1750
2 3583 1 1750
2 3584 1 1751
2 3585 1 1751
2 3586 1 1754
2 3587 1 1754
2 3588 1 1756
2 3589 1 1756
2 3590 1 1757
2 3591 1 1757
2 3592 1 1758
2 3593 1 1758
2 3594 1 1758
2 3595 1 1759
2 3596 1 1759
2 3597 1 1762
2 3598 1 1762
2 3599 1 1763
2 3600 1 1763
2 3601 1 1768
2 3602 1 1768
2 3603 1 1768
2 3604 1 1769
2 3605 1 1769
2 3606 1 1774
2 3607 1 1774
2 3608 1 1774
2 3609 1 1775
2 3610 1 1775
2 3611 1 1782
2 3612 1 1782
2 3613 1 1782
2 3614 1 1783
2 3615 1 1783
2 3616 1 1786
2 3617 1 1786
2 3618 1 1786
2 3619 1 1787
2 3620 1 1787
2 3621 1 1794
2 3622 1 1794
2 3623 1 1794
2 3624 1 1795
2 3625 1 1795
2 3626 1 1800
2 3627 1 1800
2 3628 1 1801
2 3629 1 1801
2 3630 1 1804
2 3631 1 1804
2 3632 1 1805
2 3633 1 1805
2 3634 1 1810
2 3635 1 1810
2 3636 1 1811
2 3637 1 1811
2 3638 1 1814
2 3639 1 1814
2 3640 1 1815
2 3641 1 1815
2 3642 1 1853
2 3643 1 1853
2 3644 1 1855
2 3645 1 1855
2 3646 1 1868
2 3647 1 1868
2 3648 1 1870
2 3649 1 1870
2 3650 1 1871
2 3651 1 1871
0 33 5 2 1 1990
0 34 5 2 1 2000
0 35 5 2 1 2010
0 36 5 2 1 2021
0 37 5 2 1 2031
0 38 5 2 1 2042
0 39 5 2 1 2052
0 40 5 2 1 2062
0 41 5 2 1 2072
0 42 5 2 1 2082
0 43 5 2 1 2093
0 44 5 2 1 2103
0 45 5 2 1 2113
0 46 5 2 1 2123
0 47 5 2 1 2133
0 48 5 3 1 2143
0 49 5 3 1 2146
0 50 5 3 1 2149
0 51 5 3 1 2152
0 52 5 3 1 2155
0 53 5 3 1 2158
0 54 5 3 1 2161
0 55 5 3 1 2164
0 56 5 3 1 2167
0 57 5 3 1 2170
0 58 5 3 1 2173
0 59 5 3 1 2176
0 60 5 4 1 2179
0 61 5 3 1 2183
0 62 5 2 1 2186
0 63 5 2 1 2190
0 64 7 2 2 2264 2267
0 65 5 1 1 2271
0 66 7 3 2 2191 2272
0 67 5 1 1 2273
0 68 7 2 2 2265 2192
0 69 5 1 1 2276
0 70 7 1 2 65 2277
0 71 5 1 1 70
0 72 7 1 2 2184 2269
0 73 5 1 1 72
0 74 7 2 2 71 73
0 75 5 1 1 2278
0 76 7 2 2 2260 2279
0 77 5 1 1 2280
0 78 7 1 2 2187 69
0 79 7 1 2 77 78
0 80 5 1 1 79
0 81 7 2 2 67 80
0 82 5 1 1 2282
0 83 7 1 2 2261 82
0 84 5 2 1 83
0 85 7 1 2 2180 2283
0 86 5 1 1 85
0 87 7 2 2 2284 86
0 88 5 1 1 2286
0 89 7 2 2 2257 2287
0 90 5 2 1 2288
0 91 7 1 2 75 2285
0 92 5 1 1 91
0 93 7 1 2 2262 2274
0 94 5 1 1 93
0 95 7 2 2 92 94
0 96 5 1 1 2292
0 97 7 1 2 2290 96
0 98 5 2 1 97
0 99 7 1 2 2188 2281
0 100 5 1 1 99
0 101 7 1 2 2181 2275
0 102 5 1 1 101
0 103 7 2 2 100 102
0 104 5 2 1 2296
0 105 7 2 2 2294 2297
0 106 5 1 1 2300
0 107 7 1 2 2258 106
0 108 5 2 1 107
0 109 7 1 2 2177 2301
0 110 5 1 1 109
0 111 7 2 2 2302 110
0 112 5 1 1 2304
0 113 7 2 2 2254 2305
0 114 5 2 1 2306
0 115 7 1 2 88 2303
0 116 5 1 1 115
0 117 7 1 2 2289 2298
0 118 5 1 1 117
0 119 7 2 2 116 118
0 120 5 1 1 2310
0 121 7 1 2 2308 120
0 122 5 2 1 121
0 123 7 1 2 2291 2299
0 124 5 1 1 123
0 125 7 1 2 2293 124
0 126 5 1 1 125
0 127 7 3 2 2295 126
0 128 5 1 1 2314
0 129 7 2 2 2312 128
0 130 5 1 1 2317
0 131 7 1 2 2255 130
0 132 5 2 1 131
0 133 7 1 2 2174 2318
0 134 5 1 1 133
0 135 7 2 2 2319 134
0 136 5 1 1 2321
0 137 7 2 2 2251 2322
0 138 5 2 1 2323
0 139 7 1 2 112 2320
0 140 5 1 1 139
0 141 7 1 2 2307 2315
0 142 5 1 1 141
0 143 7 2 2 140 142
0 144 5 1 1 2327
0 145 7 1 2 2325 144
0 146 5 2 1 145
0 147 7 1 2 2309 2316
0 148 5 1 1 147
0 149 7 1 2 2311 148
0 150 5 1 1 149
0 151 7 3 2 2313 150
0 152 5 1 1 2331
0 153 7 2 2 2329 152
0 154 5 1 1 2334
0 155 7 1 2 2252 154
0 156 5 2 1 155
0 157 7 1 2 2171 2335
0 158 5 1 1 157
0 159 7 2 2 2336 158
0 160 5 1 1 2338
0 161 7 2 2 2248 2339
0 162 5 2 1 2340
0 163 7 1 2 136 2337
0 164 5 1 1 163
0 165 7 1 2 2324 2332
0 166 5 1 1 165
0 167 7 2 2 164 166
0 168 5 1 1 2344
0 169 7 1 2 2342 168
0 170 5 2 1 169
0 171 7 1 2 2326 2333
0 172 5 1 1 171
0 173 7 1 2 2328 172
0 174 5 1 1 173
0 175 7 3 2 2330 174
0 176 5 1 1 2348
0 177 7 2 2 2346 176
0 178 5 1 1 2351
0 179 7 1 2 2249 178
0 180 5 2 1 179
0 181 7 1 2 2168 2352
0 182 5 1 1 181
0 183 7 2 2 2353 182
0 184 5 1 1 2355
0 185 7 2 2 2245 2356
0 186 5 2 1 2357
0 187 7 1 2 160 2354
0 188 5 1 1 187
0 189 7 1 2 2341 2349
0 190 5 1 1 189
0 191 7 2 2 188 190
0 192 5 1 1 2361
0 193 7 1 2 2359 192
0 194 5 2 1 193
0 195 7 1 2 2343 2350
0 196 5 1 1 195
0 197 7 1 2 2345 196
0 198 5 1 1 197
0 199 7 3 2 2347 198
0 200 5 1 1 2365
0 201 7 2 2 2363 200
0 202 5 1 1 2368
0 203 7 1 2 2246 202
0 204 5 2 1 203
0 205 7 1 2 2165 2369
0 206 5 1 1 205
0 207 7 2 2 2370 206
0 208 5 1 1 2372
0 209 7 2 2 2242 2373
0 210 5 2 1 2374
0 211 7 1 2 184 2371
0 212 5 1 1 211
0 213 7 1 2 2358 2366
0 214 5 1 1 213
0 215 7 2 2 212 214
0 216 5 1 1 2378
0 217 7 1 2 2376 216
0 218 5 2 1 217
0 219 7 1 2 2360 2367
0 220 5 1 1 219
0 221 7 1 2 2362 220
0 222 5 1 1 221
0 223 7 3 2 2364 222
0 224 5 1 1 2382
0 225 7 2 2 2380 224
0 226 5 1 1 2385
0 227 7 1 2 2243 226
0 228 5 2 1 227
0 229 7 1 2 2162 2386
0 230 5 1 1 229
0 231 7 2 2 2387 230
0 232 5 1 1 2389
0 233 7 2 2 2239 2390
0 234 5 2 1 2391
0 235 7 1 2 208 2388
0 236 5 1 1 235
0 237 7 1 2 2375 2383
0 238 5 1 1 237
0 239 7 2 2 236 238
0 240 5 1 1 2395
0 241 7 1 2 2393 240
0 242 5 2 1 241
0 243 7 1 2 2377 2384
0 244 5 1 1 243
0 245 7 1 2 2379 244
0 246 5 1 1 245
0 247 7 3 2 2381 246
0 248 5 1 1 2399
0 249 7 2 2 2397 248
0 250 5 1 1 2402
0 251 7 1 2 2240 250
0 252 5 2 1 251
0 253 7 1 2 2159 2403
0 254 5 1 1 253
0 255 7 2 2 2404 254
0 256 5 1 1 2406
0 257 7 2 2 2236 2407
0 258 5 2 1 2408
0 259 7 1 2 232 2405
0 260 5 1 1 259
0 261 7 1 2 2392 2400
0 262 5 1 1 261
0 263 7 2 2 260 262
0 264 5 1 1 2412
0 265 7 1 2 2410 264
0 266 5 2 1 265
0 267 7 1 2 2394 2401
0 268 5 1 1 267
0 269 7 1 2 2396 268
0 270 5 1 1 269
0 271 7 3 2 2398 270
0 272 5 1 1 2416
0 273 7 2 2 2414 272
0 274 5 1 1 2419
0 275 7 1 2 2237 274
0 276 5 2 1 275
0 277 7 1 2 2156 2420
0 278 5 1 1 277
0 279 7 2 2 2421 278
0 280 5 1 1 2423
0 281 7 2 2 2233 2424
0 282 5 2 1 2425
0 283 7 1 2 256 2422
0 284 5 1 1 283
0 285 7 1 2 2409 2417
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 2429
0 289 7 1 2 2427 288
0 290 5 2 1 289
0 291 7 1 2 2411 2418
0 292 5 1 1 291
0 293 7 1 2 2413 292
0 294 5 1 1 293
0 295 7 3 2 2415 294
0 296 5 1 1 2433
0 297 7 2 2 2431 296
0 298 5 1 1 2436
0 299 7 1 2 2234 298
0 300 5 2 1 299
0 301 7 1 2 2153 2437
0 302 5 1 1 301
0 303 7 2 2 2438 302
0 304 5 1 1 2440
0 305 7 2 2 2230 2441
0 306 5 2 1 2442
0 307 7 1 2 280 2439
0 308 5 1 1 307
0 309 7 1 2 2426 2434
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 2446
0 313 7 1 2 2444 312
0 314 5 2 1 313
0 315 7 1 2 2428 2435
0 316 5 1 1 315
0 317 7 1 2 2430 316
0 318 5 1 1 317
0 319 7 3 2 2432 318
0 320 5 1 1 2450
0 321 7 2 2 2448 320
0 322 5 1 1 2453
0 323 7 1 2 2231 322
0 324 5 2 1 323
0 325 7 1 2 2150 2454
0 326 5 1 1 325
0 327 7 2 2 2455 326
0 328 5 1 1 2457
0 329 7 2 2 2227 2458
0 330 5 2 1 2459
0 331 7 1 2 304 2456
0 332 5 1 1 331
0 333 7 1 2 2443 2451
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 2463
0 337 7 1 2 2461 336
0 338 5 2 1 337
0 339 7 1 2 2445 2452
0 340 5 1 1 339
0 341 7 1 2 2447 340
0 342 5 1 1 341
0 343 7 3 2 2449 342
0 344 5 1 1 2467
0 345 7 2 2 2465 344
0 346 5 1 1 2470
0 347 7 1 2 2228 346
0 348 5 2 1 347
0 349 7 1 2 2147 2471
0 350 5 1 1 349
0 351 7 2 2 2472 350
0 352 5 1 1 2474
0 353 7 2 2 2224 2475
0 354 5 2 1 2476
0 355 7 1 2 328 2473
0 356 5 1 1 355
0 357 7 1 2 2460 2468
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 2480
0 361 7 1 2 2478 360
0 362 5 2 1 361
0 363 7 1 2 2462 2469
0 364 5 1 1 363
0 365 7 1 2 2464 364
0 366 5 1 1 365
0 367 7 3 2 2466 366
0 368 5 1 1 2484
0 369 7 2 2 2482 368
0 370 5 1 1 2487
0 371 7 1 2 2225 370
0 372 5 2 1 371
0 373 7 1 2 2144 2488
0 374 5 1 1 373
0 375 7 2 2 2489 374
0 376 5 1 1 2491
0 377 7 2 2 2222 2492
0 378 5 2 1 2493
0 379 7 1 2 352 2490
0 380 5 1 1 379
0 381 7 1 2 2477 2485
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 2497
0 385 7 1 2 2495 384
0 386 5 2 1 385
0 387 7 1 2 2479 2486
0 388 5 1 1 387
0 389 7 1 2 2481 388
0 390 5 1 1 389
0 391 7 3 2 2483 390
0 392 5 1 1 2501
0 393 7 2 2 2499 392
0 394 5 1 1 2504
0 395 7 1 2 2223 394
0 396 5 2 1 395
0 397 7 1 2 2134 2505
0 398 5 1 1 397
0 399 7 2 2 2506 398
0 400 5 1 1 2508
0 401 7 2 2 2220 2509
0 402 5 2 1 2510
0 403 7 1 2 376 2507
0 404 5 1 1 403
0 405 7 1 2 2494 2502
0 406 5 1 1 405
0 407 7 2 2 404 406
0 408 5 1 1 2514
0 409 7 1 2 2512 408
0 410 5 2 1 409
0 411 7 1 2 2496 2503
0 412 5 1 1 411
0 413 7 1 2 2498 412
0 414 5 1 1 413
0 415 7 3 2 2500 414
0 416 5 1 1 2518
0 417 7 2 2 2516 416
0 418 5 1 1 2521
0 419 7 1 2 2221 418
0 420 5 2 1 419
0 421 7 1 2 2124 2522
0 422 5 1 1 421
0 423 7 2 2 2523 422
0 424 5 1 1 2525
0 425 7 2 2 2218 2526
0 426 5 2 1 2527
0 427 7 1 2 400 2524
0 428 5 1 1 427
0 429 7 1 2 2511 2519
0 430 5 1 1 429
0 431 7 2 2 428 430
0 432 5 1 1 2531
0 433 7 1 2 2529 432
0 434 5 2 1 433
0 435 7 1 2 2513 2520
0 436 5 1 1 435
0 437 7 1 2 2515 436
0 438 5 1 1 437
0 439 7 3 2 2517 438
0 440 5 1 1 2535
0 441 7 2 2 2533 440
0 442 5 1 1 2538
0 443 7 1 2 2219 442
0 444 5 2 1 443
0 445 7 1 2 2114 2539
0 446 5 1 1 445
0 447 7 2 2 2540 446
0 448 5 1 1 2542
0 449 7 2 2 2216 2543
0 450 5 2 1 2544
0 451 7 1 2 424 2541
0 452 5 1 1 451
0 453 7 1 2 2528 2536
0 454 5 1 1 453
0 455 7 2 2 452 454
0 456 5 1 1 2548
0 457 7 1 2 2546 456
0 458 5 2 1 457
0 459 7 1 2 2530 2537
0 460 5 1 1 459
0 461 7 1 2 2532 460
0 462 5 1 1 461
0 463 7 3 2 2534 462
0 464 5 1 1 2552
0 465 7 2 2 2550 464
0 466 5 1 1 2555
0 467 7 1 2 2217 466
0 468 5 2 1 467
0 469 7 1 2 2104 2556
0 470 5 1 1 469
0 471 7 2 2 2557 470
0 472 5 1 1 2559
0 473 7 2 2 2214 2560
0 474 5 2 1 2561
0 475 7 1 2 448 2558
0 476 5 1 1 475
0 477 7 1 2 2545 2553
0 478 5 1 1 477
0 479 7 2 2 476 478
0 480 5 1 1 2565
0 481 7 1 2 2563 480
0 482 5 2 1 481
0 483 7 1 2 2547 2554
0 484 5 1 1 483
0 485 7 1 2 2549 484
0 486 5 1 1 485
0 487 7 3 2 2551 486
0 488 5 1 1 2569
0 489 7 2 2 2567 488
0 490 5 1 1 2572
0 491 7 1 2 2215 490
0 492 5 2 1 491
0 493 7 1 2 2094 2573
0 494 5 1 1 493
0 495 7 2 2 2574 494
0 496 5 1 1 2576
0 497 7 2 2 2212 2577
0 498 5 2 1 2578
0 499 7 1 2 472 2575
0 500 5 1 1 499
0 501 7 1 2 2562 2570
0 502 5 1 1 501
0 503 7 2 2 500 502
0 504 5 1 1 2582
0 505 7 1 2 2580 504
0 506 5 2 1 505
0 507 7 1 2 2564 2571
0 508 5 1 1 507
0 509 7 1 2 2566 508
0 510 5 1 1 509
0 511 7 3 2 2568 510
0 512 5 1 1 2586
0 513 7 2 2 2584 512
0 514 5 1 1 2589
0 515 7 1 2 2213 514
0 516 5 2 1 515
0 517 7 1 2 2083 2590
0 518 5 1 1 517
0 519 7 2 2 2591 518
0 520 5 1 1 2593
0 521 7 2 2 2210 2594
0 522 5 2 1 2595
0 523 7 1 2 496 2592
0 524 5 1 1 523
0 525 7 1 2 2579 2587
0 526 5 1 1 525
0 527 7 2 2 524 526
0 528 5 1 1 2599
0 529 7 1 2 2597 528
0 530 5 2 1 529
0 531 7 1 2 2581 2588
0 532 5 1 1 531
0 533 7 1 2 2583 532
0 534 5 1 1 533
0 535 7 3 2 2585 534
0 536 5 1 1 2603
0 537 7 2 2 2601 536
0 538 5 1 1 2606
0 539 7 1 2 2211 538
0 540 5 2 1 539
0 541 7 1 2 2073 2607
0 542 5 1 1 541
0 543 7 2 2 2608 542
0 544 5 1 1 2610
0 545 7 2 2 2208 2611
0 546 5 2 1 2612
0 547 7 1 2 520 2609
0 548 5 1 1 547
0 549 7 1 2 2596 2604
0 550 5 1 1 549
0 551 7 2 2 548 550
0 552 5 1 1 2616
0 553 7 1 2 2614 552
0 554 5 2 1 553
0 555 7 1 2 2598 2605
0 556 5 1 1 555
0 557 7 1 2 2600 556
0 558 5 1 1 557
0 559 7 3 2 2602 558
0 560 5 1 1 2620
0 561 7 2 2 2618 560
0 562 5 1 1 2623
0 563 7 1 2 2209 562
0 564 5 2 1 563
0 565 7 1 2 2063 2624
0 566 5 1 1 565
0 567 7 2 2 2625 566
0 568 5 1 1 2627
0 569 7 2 2 2206 2628
0 570 5 2 1 2629
0 571 7 1 2 544 2626
0 572 5 1 1 571
0 573 7 1 2 2613 2621
0 574 5 1 1 573
0 575 7 2 2 572 574
0 576 5 1 1 2633
0 577 7 1 2 2631 576
0 578 5 2 1 577
0 579 7 1 2 2615 2622
0 580 5 1 1 579
0 581 7 1 2 2617 580
0 582 5 1 1 581
0 583 7 3 2 2619 582
0 584 5 1 1 2637
0 585 7 2 2 2635 584
0 586 5 1 1 2640
0 587 7 1 2 2207 586
0 588 5 2 1 587
0 589 7 1 2 2053 2641
0 590 5 1 1 589
0 591 7 2 2 2642 590
0 592 5 1 1 2644
0 593 7 2 2 2204 2645
0 594 5 2 1 2646
0 595 7 1 2 568 2643
0 596 5 1 1 595
0 597 7 1 2 2630 2638
0 598 5 1 1 597
0 599 7 2 2 596 598
0 600 5 1 1 2650
0 601 7 1 2 2648 600
0 602 5 2 1 601
0 603 7 1 2 2632 2639
0 604 5 1 1 603
0 605 7 1 2 2634 604
0 606 5 1 1 605
0 607 7 3 2 2636 606
0 608 5 1 1 2654
0 609 7 2 2 2652 608
0 610 5 1 1 2657
0 611 7 1 2 2205 610
0 612 5 2 1 611
0 613 7 1 2 2043 2658
0 614 5 1 1 613
0 615 7 2 2 2659 614
0 616 5 1 1 2661
0 617 7 2 2 2202 2662
0 618 5 2 1 2663
0 619 7 1 2 592 2660
0 620 5 1 1 619
0 621 7 1 2 2647 2655
0 622 5 1 1 621
0 623 7 2 2 620 622
0 624 5 1 1 2667
0 625 7 1 2 2665 624
0 626 5 2 1 625
0 627 7 1 2 2649 2656
0 628 5 1 1 627
0 629 7 1 2 2651 628
0 630 5 1 1 629
0 631 7 3 2 2653 630
0 632 5 1 1 2671
0 633 7 2 2 2669 632
0 634 5 1 1 2674
0 635 7 1 2 2203 634
0 636 5 2 1 635
0 637 7 1 2 2032 2675
0 638 5 1 1 637
0 639 7 2 2 2676 638
0 640 5 1 1 2678
0 641 7 2 2 2200 2679
0 642 5 2 1 2680
0 643 7 1 2 616 2677
0 644 5 1 1 643
0 645 7 1 2 2664 2672
0 646 5 1 1 645
0 647 7 2 2 644 646
0 648 5 1 1 2684
0 649 7 1 2 2682 648
0 650 5 2 1 649
0 651 7 1 2 2666 2673
0 652 5 1 1 651
0 653 7 1 2 2668 652
0 654 5 1 1 653
0 655 7 3 2 2670 654
0 656 5 1 1 2688
0 657 7 2 2 2686 656
0 658 5 1 1 2691
0 659 7 1 2 2201 658
0 660 5 2 1 659
0 661 7 1 2 2022 2692
0 662 5 1 1 661
0 663 7 2 2 2693 662
0 664 5 1 1 2695
0 665 7 2 2 2198 2696
0 666 5 2 1 2697
0 667 7 1 2 640 2694
0 668 5 1 1 667
0 669 7 1 2 2681 2689
0 670 5 1 1 669
0 671 7 2 2 668 670
0 672 5 1 1 2701
0 673 7 1 2 2699 672
0 674 5 2 1 673
0 675 7 1 2 2683 2690
0 676 5 1 1 675
0 677 7 1 2 2685 676
0 678 5 1 1 677
0 679 7 3 2 2687 678
0 680 5 1 1 2705
0 681 7 2 2 2703 680
0 682 5 1 1 2708
0 683 7 1 2 2011 2709
0 684 5 1 1 683
0 685 7 1 2 2199 682
0 686 5 2 1 685
0 687 7 3 2 684 2710
0 688 5 2 1 2712
0 689 7 2 2 2196 2713
0 690 5 2 1 2717
0 691 7 1 2 664 2711
0 692 5 1 1 691
0 693 7 1 2 2698 2706
0 694 5 1 1 693
0 695 7 2 2 692 694
0 696 5 1 1 2721
0 697 7 1 2 2719 696
0 698 5 2 1 697
0 699 7 1 2 2700 2707
0 700 5 1 1 699
0 701 7 1 2 2702 700
0 702 5 1 1 701
0 703 7 3 2 2704 702
0 704 5 1 1 2725
0 705 7 1 2 2720 2726
0 706 5 1 1 705
0 707 7 1 2 2722 706
0 708 5 1 1 707
0 709 7 1 2 2723 708
0 710 5 1 1 709
0 711 7 2 2 2724 704
0 712 5 1 1 2728
0 713 7 1 2 2197 712
0 714 5 2 1 713
0 715 7 1 2 2001 2729
0 716 5 1 1 715
0 717 7 2 2 2730 716
0 718 7 1 2 2194 2732
0 719 5 1 1 718
0 720 7 1 2 2715 2731
0 721 5 1 1 720
0 722 7 1 2 2718 2727
0 723 5 1 1 722
0 724 7 1 2 721 723
0 725 5 1 1 724
0 726 7 1 2 719 725
0 727 5 1 1 726
0 728 7 2 2 710 727
0 729 5 1 1 2734
0 730 7 1 2 2195 2714
0 731 5 1 1 730
0 732 7 1 2 2735 731
0 733 5 1 1 732
0 734 7 1 2 1991 2716
0 735 5 1 1 734
0 736 7 1 2 729 735
0 737 5 1 1 736
0 738 7 1 2 2733 737
0 739 7 2 2 733 738
0 740 5 1 1 2736
0 741 7 2 2 2023 2135
0 742 5 1 1 2738
0 743 7 2 2 2054 2105
0 744 5 1 1 2740
0 745 7 1 2 2739 2741
0 746 5 2 1 745
0 747 7 2 2 2044 2115
0 748 5 1 1 2744
0 749 7 1 2 742 744
0 750 5 1 1 749
0 751 7 2 2 750 2742
0 752 5 1 1 2746
0 753 7 1 2 2745 2747
0 754 5 2 1 753
0 755 7 2 2 2743 2748
0 756 5 1 1 2750
0 757 7 2 2 2045 2125
0 758 5 2 1 2752
0 759 7 2 2 2055 2116
0 760 5 1 1 2756
0 761 7 2 2 2033 2136
0 762 5 1 1 2758
0 763 7 1 2 760 762
0 764 5 1 1 763
0 765 7 1 2 2757 2759
0 766 5 2 1 765
0 767 7 2 2 764 2760
0 768 5 1 1 2762
0 769 7 1 2 2753 2763
0 770 5 2 1 769
0 771 7 1 2 2754 768
0 772 5 1 1 771
0 773 7 2 2 2764 772
0 774 5 1 1 2766
0 775 7 1 2 756 2767
0 776 5 2 1 775
0 777 7 2 2 2034 2126
0 778 5 1 1 2770
0 779 7 1 2 748 752
0 780 5 1 1 779
0 781 7 2 2 2749 780
0 782 5 1 1 2772
0 783 7 1 2 2771 2773
0 784 5 2 1 783
0 785 7 2 2 2012 2137
0 786 5 1 1 2776
0 787 7 2 2 2056 2095
0 788 5 1 1 2778
0 789 7 1 2 2777 2779
0 790 5 2 1 789
0 791 7 2 2 2046 2106
0 792 5 1 1 2782
0 793 7 1 2 786 788
0 794 5 1 1 793
0 795 7 2 2 794 2780
0 796 5 1 1 2784
0 797 7 1 2 2783 2785
0 798 5 2 1 797
0 799 7 2 2 2781 2786
0 800 5 1 1 2788
0 801 7 1 2 778 782
0 802 5 1 1 801
0 803 7 2 2 2774 802
0 804 5 1 1 2790
0 805 7 1 2 800 2791
0 806 5 2 1 805
0 807 7 2 2 2775 2792
0 808 5 1 1 2794
0 809 7 1 2 2751 774
0 810 5 1 1 809
0 811 7 2 2 2768 810
0 812 5 1 1 2796
0 813 7 1 2 808 2797
0 814 5 2 1 813
0 815 7 2 2 2769 2798
0 816 5 1 1 2800
0 817 7 2 2 2761 2765
0 818 5 1 1 2802
0 819 7 2 2 2047 2138
0 820 5 1 1 2804
0 821 7 2 2 2057 2127
0 822 5 1 1 2806
0 823 7 1 2 820 2807
0 824 5 1 1 823
0 825 7 1 2 2805 822
0 826 5 1 1 825
0 827 7 2 2 824 826
0 828 5 1 1 2808
0 829 7 1 2 818 828
0 830 5 3 1 829
0 831 7 1 2 2803 2809
0 832 5 1 1 831
0 833 7 2 2 2810 832
0 834 5 1 1 2813
0 835 7 1 2 816 2814
0 836 5 2 1 835
0 837 7 2 2 2024 2128
0 838 5 1 1 2817
0 839 7 1 2 792 796
0 840 5 1 1 839
0 841 7 2 2 2787 840
0 842 5 1 1 2819
0 843 7 1 2 2818 2820
0 844 5 2 1 843
0 845 7 2 2 2035 2117
0 846 5 1 1 2823
0 847 7 1 2 838 842
0 848 5 1 1 847
0 849 7 2 2 2821 848
0 850 5 1 1 2825
0 851 7 1 2 2824 2826
0 852 5 2 1 851
0 853 7 2 2 2822 2827
0 854 5 1 1 2829
0 855 7 1 2 2789 804
0 856 5 1 1 855
0 857 7 2 2 2793 856
0 858 5 1 1 2831
0 859 7 1 2 854 2832
0 860 5 2 1 859
0 861 7 2 2 2002 2139
0 862 5 1 1 2835
0 863 7 2 2 2058 2064
0 864 5 1 1 2837
0 865 7 2 2 2048 2074
0 866 5 1 1 2839
0 867 7 2 2 2838 2840
0 868 5 2 1 2841
0 869 7 2 2 2084 2842
0 870 5 2 1 2845
0 871 7 1 2 2836 2846
0 872 5 2 1 871
0 873 7 2 2 2059 2085
0 874 5 1 1 2851
0 875 7 1 2 862 2847
0 876 5 1 1 875
0 877 7 2 2 2849 876
0 878 5 1 1 2853
0 879 7 1 2 2852 2854
0 880 5 2 1 879
0 881 7 2 2 2850 2855
0 882 5 1 1 2857
0 883 7 1 2 846 850
0 884 5 1 1 883
0 885 7 2 2 2828 884
0 886 5 1 1 2859
0 887 7 1 2 882 2860
0 888 5 2 1 887
0 889 7 2 2 2036 2107
0 890 5 1 1 2863
0 891 7 1 2 874 878
0 892 5 1 1 891
0 893 7 2 2 2856 892
0 894 5 1 1 2865
0 895 7 1 2 2864 2866
0 896 5 2 1 895
0 897 7 2 2 2049 2096
0 898 5 1 1 2869
0 899 7 1 2 890 894
0 900 5 1 1 899
0 901 7 2 2 2867 900
0 902 5 1 1 2871
0 903 7 1 2 2870 2872
0 904 5 2 1 903
0 905 7 2 2 2868 2873
0 906 5 1 1 2875
0 907 7 1 2 2858 886
0 908 5 1 1 907
0 909 7 2 2 2861 908
0 910 5 1 1 2877
0 911 7 1 2 906 2878
0 912 5 2 1 911
0 913 7 2 2 2862 2879
0 914 5 1 1 2881
0 915 7 1 2 2830 858
0 916 5 1 1 915
0 917 7 2 2 2833 916
0 918 5 1 1 2883
0 919 7 1 2 914 2884
0 920 5 2 1 919
0 921 7 2 2 2834 2885
0 922 5 1 1 2887
0 923 7 1 2 2795 812
0 924 5 1 1 923
0 925 7 2 2 2799 924
0 926 5 1 1 2889
0 927 7 1 2 922 2890
0 928 5 2 1 927
0 929 7 2 2 2013 2129
0 930 5 1 1 2893
0 931 7 2 2 2025 2118
0 932 5 1 1 2895
0 933 7 1 2 2894 2896
0 934 5 2 1 933
0 935 7 1 2 898 902
0 936 5 1 1 935
0 937 7 2 2 2874 936
0 938 5 1 1 2899
0 939 7 1 2 930 932
0 940 5 1 1 939
0 941 7 2 2 2897 940
0 942 5 1 1 2901
0 943 7 1 2 2900 2902
0 944 5 2 1 943
0 945 7 2 2 2898 2903
0 946 5 1 1 2905
0 947 7 1 2 2876 910
0 948 5 1 1 947
0 949 7 2 2 2880 948
0 950 5 1 1 2907
0 951 7 1 2 946 2908
0 952 5 2 1 951
0 953 7 2 2 2037 2097
0 954 5 1 1 2911
0 955 7 2 2 2003 2130
0 956 5 1 1 2913
0 957 7 1 2 2912 2914
0 958 5 2 1 957
0 959 7 2 2 1992 2140
0 960 5 1 1 2917
0 961 7 2 2 2026 2108
0 962 5 1 1 2919
0 963 7 1 2 2050 2086
0 964 5 1 1 963
0 965 7 1 2 2843 964
0 966 5 1 1 965
0 967 7 2 2 2848 966
0 968 5 1 1 2921
0 969 7 1 2 2920 2922
0 970 5 2 1 969
0 971 7 1 2 962 968
0 972 5 1 1 971
0 973 7 2 2 2923 972
0 974 5 1 1 2925
0 975 7 1 2 2918 2926
0 976 5 2 1 975
0 977 7 1 2 960 974
0 978 5 1 1 977
0 979 7 2 2 2927 978
0 980 5 1 1 2929
0 981 7 1 2 954 956
0 982 5 1 1 981
0 983 7 2 2 2915 982
0 984 5 1 1 2931
0 985 7 1 2 2930 2932
0 986 5 2 1 985
0 987 7 2 2 2916 2933
0 988 5 1 1 2935
0 989 7 1 2 938 942
0 990 5 1 1 989
0 991 7 2 2 2904 990
0 992 5 1 1 2937
0 993 7 1 2 988 2938
0 994 5 2 1 993
0 995 7 2 2 2060 2075
0 996 5 1 1 2941
0 997 7 2 2 2014 2119
0 998 5 1 1 2943
0 999 7 1 2 2942 2944
0 1000 5 2 1 999
0 1001 7 1 2 980 984
0 1002 5 1 1 1001
0 1003 7 2 2 2934 1002
0 1004 5 1 1 2947
0 1005 7 1 2 996 998
0 1006 5 1 1 1005
0 1007 7 2 2 2945 1006
0 1008 5 1 1 2949
0 1009 7 1 2 2948 2950
0 1010 5 2 1 1009
0 1011 7 2 2 2946 2951
0 1012 5 1 1 2953
0 1013 7 1 2 2936 992
0 1014 5 1 1 1013
0 1015 7 2 2 2939 1014
0 1016 5 1 1 2955
0 1017 7 1 2 1012 2956
0 1018 5 2 1 1017
0 1019 7 2 2 2940 2957
0 1020 5 1 1 2959
0 1021 7 1 2 2906 950
0 1022 5 1 1 1021
0 1023 7 2 2 2909 1022
0 1024 5 1 1 2961
0 1025 7 1 2 1020 2962
0 1026 5 2 1 1025
0 1027 7 2 2 2910 2963
0 1028 5 1 1 2965
0 1029 7 1 2 2882 918
0 1030 5 1 1 1029
0 1031 7 2 2 2886 1030
0 1032 5 1 1 2967
0 1033 7 1 2 1028 2968
0 1034 5 2 1 1033
0 1035 7 2 2 2924 2928
0 1036 5 1 1 2971
0 1037 7 1 2 2954 1016
0 1038 5 1 1 1037
0 1039 7 2 2 2958 1038
0 1040 5 1 1 2973
0 1041 7 1 2 1036 2974
0 1042 5 2 1 1041
0 1043 7 2 2 2015 2109
0 1044 5 1 1 2977
0 1045 7 2 2 2027 2076
0 1046 5 1 1 2979
0 1047 7 2 2 32 2098
0 1048 5 1 1 2981
0 1049 7 2 2 2004 2077
0 1050 5 1 1 2983
0 1051 7 2 2 2982 2984
0 1052 5 2 1 2985
0 1053 7 2 2 2016 2986
0 1054 5 2 1 2989
0 1055 7 2 2 2980 2990
0 1056 5 2 1 2993
0 1057 7 2 2 2038 2994
0 1058 5 2 1 2997
0 1059 7 1 2 2978 2998
0 1060 5 2 1 1059
0 1061 7 1 2 1044 2999
0 1062 5 1 1 1061
0 1063 7 2 2 3001 1062
0 1064 5 1 1 3003
0 1065 7 1 2 864 866
0 1066 5 1 1 1065
0 1067 7 2 2 2844 1066
0 1068 5 1 1 3005
0 1069 7 1 2 3004 3006
0 1070 5 2 1 1069
0 1071 7 2 2 3002 3007
0 1072 5 1 1 3009
0 1073 7 1 2 1004 1008
0 1074 5 1 1 1073
0 1075 7 2 2 2952 1074
0 1076 5 1 1 3011
0 1077 7 1 2 1072 3012
0 1078 5 2 1 1077
0 1079 7 2 2 2005 2120
0 1080 5 1 1 3015
0 1081 7 2 2 1983 2141
0 1082 5 1 1 3017
0 1083 7 1 2 3016 3018
0 1084 5 2 1 1083
0 1085 7 1 2 1064 1068
0 1086 5 1 1 1085
0 1087 7 2 2 3008 1086
0 1088 5 1 1 3021
0 1089 7 1 2 1080 1082
0 1090 5 1 1 1089
0 1091 7 2 2 3019 1090
0 1092 5 1 1 3023
0 1093 7 1 2 3022 3024
0 1094 5 2 1 1093
0 1095 7 2 2 3020 3025
0 1096 5 1 1 3027
0 1097 7 1 2 3010 1076
0 1098 5 1 1 1097
0 1099 7 2 2 3013 1098
0 1100 5 1 1 3029
0 1101 7 1 2 1096 3030
0 1102 5 2 1 1101
0 1103 7 2 2 3014 3031
0 1104 5 1 1 3033
0 1105 7 1 2 2972 1040
0 1106 5 1 1 1105
0 1107 7 2 2 2975 1106
0 1108 5 1 1 3035
0 1109 7 1 2 1104 3036
0 1110 5 2 1 1109
0 1111 7 2 2 2976 3037
0 1112 5 1 1 3039
0 1113 7 1 2 2960 1024
0 1114 5 1 1 1113
0 1115 7 2 2 2964 1114
0 1116 5 1 1 3041
0 1117 7 1 2 1112 3042
0 1118 5 2 1 1117
0 1119 7 2 2 2039 2087
0 1120 5 1 1 3045
0 1121 7 2 2 2028 2099
0 1122 5 1 1 3047
0 1123 7 1 2 3046 3048
0 1124 5 2 1 1123
0 1125 7 2 2 1993 2131
0 1126 5 1 1 3051
0 1127 7 1 2 1120 1122
0 1128 5 1 1 1127
0 1129 7 2 2 3049 1128
0 1130 5 1 1 3053
0 1131 7 1 2 3052 3054
0 1132 5 2 1 1131
0 1133 7 2 2 3050 3055
0 1134 5 1 1 3057
0 1135 7 1 2 3028 1100
0 1136 5 1 1 1135
0 1137 7 2 2 3032 1136
0 1138 5 1 1 3059
0 1139 7 1 2 1134 3060
0 1140 5 2 1 1139
0 1141 7 1 2 1126 1130
0 1142 5 1 1 1141
0 1143 7 2 2 3056 1142
0 1144 5 1 1 3063
0 1145 7 1 2 1088 1092
0 1146 5 1 1 1145
0 1147 7 2 2 3026 1146
0 1148 5 1 1 3065
0 1149 7 1 2 3064 3066
0 1150 5 2 1 1149
0 1151 7 2 2 2017 2100
0 1152 5 1 1 3069
0 1153 7 2 2 2006 2110
0 1154 5 1 1 3071
0 1155 7 1 2 3070 3072
0 1156 5 2 1 1155
0 1157 7 2 2 1994 2121
0 1158 5 1 1 3075
0 1159 7 1 2 1152 1154
0 1160 5 1 1 1159
0 1161 7 2 2 3073 1160
0 1162 5 1 1 3077
0 1163 7 1 2 3076 3078
0 1164 5 2 1 1163
0 1165 7 2 2 3074 3079
0 1166 5 1 1 3081
0 1167 7 1 2 1144 1148
0 1168 5 1 1 1167
0 1169 7 2 2 3067 1168
0 1170 5 1 1 3083
0 1171 7 1 2 1166 3084
0 1172 5 2 1 1171
0 1173 7 2 2 3068 3085
0 1174 5 1 1 3087
0 1175 7 1 2 3058 1138
0 1176 5 1 1 1175
0 1177 7 2 2 3061 1176
0 1178 5 1 1 3089
0 1179 7 1 2 1174 3090
0 1180 5 2 1 1179
0 1181 7 2 2 3062 3091
0 1182 5 1 1 3093
0 1183 7 1 2 3034 1108
0 1184 5 1 1 1183
0 1185 7 2 2 3038 1184
0 1186 5 1 1 3095
0 1187 7 1 2 1182 3096
0 1188 5 2 1 1187
0 1189 7 2 2 1984 2132
0 1190 5 1 1 3099
0 1191 7 1 2 1158 1162
0 1192 5 1 1 1191
0 1193 7 2 2 3080 1192
0 1194 5 1 1 3101
0 1195 7 1 2 3100 3102
0 1196 5 2 1 1195
0 1197 7 2 2 2051 2065
0 1198 5 1 1 3105
0 1199 7 2 2 2029 2088
0 1200 5 1 1 3107
0 1201 7 1 2 2040 2078
0 1202 5 1 1 1201
0 1203 7 1 2 2995 1202
0 1204 5 1 1 1203
0 1205 7 2 2 3000 1204
0 1206 5 1 1 3109
0 1207 7 1 2 3108 3110
0 1208 5 2 1 1207
0 1209 7 1 2 1200 1206
0 1210 5 1 1 1209
0 1211 7 2 2 3111 1210
0 1212 5 1 1 3113
0 1213 7 1 2 3106 3114
0 1214 5 2 1 1213
0 1215 7 1 2 1198 1212
0 1216 5 1 1 1215
0 1217 7 2 2 3115 1216
0 1218 5 1 1 3117
0 1219 7 1 2 1190 1194
0 1220 5 1 1 1219
0 1221 7 2 2 3103 1220
0 1222 5 1 1 3119
0 1223 7 1 2 3118 3120
0 1224 5 2 1 1223
0 1225 7 2 2 3104 3121
0 1226 5 1 1 3123
0 1227 7 1 2 3082 1170
0 1228 5 1 1 1227
0 1229 7 2 2 3086 1228
0 1230 5 1 1 3125
0 1231 7 1 2 1226 3126
0 1232 5 2 1 1231
0 1233 7 2 2 3112 3116
0 1234 5 1 1 3129
0 1235 7 1 2 3124 1230
0 1236 5 1 1 1235
0 1237 7 2 2 3127 1236
0 1238 5 1 1 3131
0 1239 7 1 2 1234 3132
0 1240 5 2 1 1239
0 1241 7 2 2 3128 3133
0 1242 5 1 1 3135
0 1243 7 1 2 3088 1178
0 1244 5 1 1 1243
0 1245 7 2 2 3092 1244
0 1246 5 1 1 3137
0 1247 7 1 2 1242 3138
0 1248 5 2 1 1247
0 1249 7 2 2 2018 2089
0 1250 5 1 1 3141
0 1251 7 1 2 1046 2991
0 1252 5 1 1 1251
0 1253 7 2 2 2996 1252
0 1254 5 1 1 3143
0 1255 7 1 2 3142 3144
0 1256 5 2 1 1255
0 1257 7 2 2 2041 2066
0 1258 5 1 1 3147
0 1259 7 1 2 1250 1254
0 1260 5 1 1 1259
0 1261 7 2 2 3145 1260
0 1262 5 1 1 3149
0 1263 7 1 2 3148 3150
0 1264 5 2 1 1263
0 1265 7 2 2 3146 3151
0 1266 5 1 1 3153
0 1267 7 1 2 1218 1222
0 1268 5 1 1 1267
0 1269 7 2 2 3122 1268
0 1270 5 1 1 3155
0 1271 7 1 2 1266 3156
0 1272 5 2 1 1271
0 1273 7 2 2 1985 2122
0 1274 5 1 1 3159
0 1275 7 2 2 2007 2101
0 1276 5 1 1 3161
0 1277 7 1 2 3160 3162
0 1278 5 2 1 1277
0 1279 7 1 2 1258 1262
0 1280 5 1 1 1279
0 1281 7 2 2 3152 1280
0 1282 5 1 1 3165
0 1283 7 1 2 1274 1276
0 1284 5 1 1 1283
0 1285 7 2 2 3163 1284
0 1286 5 1 1 3167
0 1287 7 1 2 3166 3168
0 1288 5 2 1 1287
0 1289 7 2 2 3164 3169
0 1290 5 1 1 3171
0 1291 7 1 2 3154 1270
0 1292 5 1 1 1291
0 1293 7 2 2 3157 1292
0 1294 5 1 1 3173
0 1295 7 1 2 1290 3174
0 1296 5 2 1 1295
0 1297 7 2 2 3158 3175
0 1298 5 1 1 3177
0 1299 7 1 2 3130 1238
0 1300 5 1 1 1299
0 1301 7 2 2 3134 1300
0 1302 5 1 1 3179
0 1303 7 1 2 1298 3180
0 1304 5 2 1 1303
0 1305 7 2 2 1995 2111
0 1306 5 1 1 3183
0 1307 7 1 2 1282 1286
0 1308 5 1 1 1307
0 1309 7 2 2 3170 1308
0 1310 5 1 1 3185
0 1311 7 1 2 3184 3186
0 1312 5 2 1 1311
0 1313 7 2 2 2008 2090
0 1314 5 1 1 3189
0 1315 7 1 2 2019 2079
0 1316 5 1 1 1315
0 1317 7 1 2 2987 1316
0 1318 5 1 1 1317
0 1319 7 2 2 2992 1318
0 1320 5 1 1 3191
0 1321 7 1 2 3190 3192
0 1322 5 2 1 1321
0 1323 7 2 2 2030 2067
0 1324 5 1 1 3195
0 1325 7 1 2 1314 1320
0 1326 5 1 1 1325
0 1327 7 2 2 3193 1326
0 1328 5 1 1 3197
0 1329 7 1 2 3196 3198
0 1330 5 2 1 1329
0 1331 7 2 2 3194 3199
0 1332 5 1 1 3201
0 1333 7 1 2 1306 1310
0 1334 5 1 1 1333
0 1335 7 2 2 3187 1334
0 1336 5 1 1 3203
0 1337 7 1 2 1332 3204
0 1338 5 2 1 1337
0 1339 7 2 2 3188 3205
0 1340 5 1 1 3207
0 1341 7 1 2 3172 1294
0 1342 5 1 1 1341
0 1343 7 2 2 3176 1342
0 1344 5 1 1 3209
0 1345 7 1 2 1340 3210
0 1346 5 2 1 1345
0 1347 7 2 2 1986 2112
0 1348 5 1 1 3213
0 1349 7 2 2 1996 2102
0 1350 5 1 1 3215
0 1351 7 1 2 3214 3216
0 1352 5 2 1 1351
0 1353 7 1 2 1324 1328
0 1354 5 1 1 1353
0 1355 7 2 2 3200 1354
0 1356 5 1 1 3219
0 1357 7 1 2 1348 1350
0 1358 5 1 1 1357
0 1359 7 2 2 3217 1358
0 1360 5 1 1 3221
0 1361 7 1 2 3220 3222
0 1362 5 2 1 1361
0 1363 7 2 2 3218 3223
0 1364 5 1 1 3225
0 1365 7 1 2 3202 1336
0 1366 5 1 1 1365
0 1367 7 2 2 3206 1366
0 1368 5 1 1 3227
0 1369 7 1 2 1364 3228
0 1370 5 2 1 1369
0 1371 7 1 2 1356 1360
0 1372 5 1 1 1371
0 1373 7 2 2 3224 1372
0 1374 5 1 1 3231
0 1375 7 2 2 1997 2091
0 1376 5 1 1 3233
0 1377 7 2 2 2020 2068
0 1378 5 1 1 3235
0 1379 7 2 2 3234 3236
0 1380 5 1 1 3237
0 1381 7 2 2 1998 2080
0 1382 5 1 1 3239
0 1383 7 2 2 1987 2092
0 1384 5 1 1 3241
0 1385 7 2 2 3240 3242
0 1386 5 2 1 3243
0 1387 7 3 2 1380 3245
0 1388 5 1 1 3247
0 1389 7 1 2 3232 1388
0 1390 5 2 1 1389
0 1391 7 1 2 1048 1050
0 1392 5 1 1 1391
0 1393 7 2 2 2988 1392
0 1394 5 1 1 3252
0 1395 7 1 2 1376 1378
0 1396 5 1 1 1395
0 1397 7 1 2 3248 1396
0 1398 5 1 1 1397
0 1399 7 1 2 3238 3244
0 1400 5 1 1 1399
0 1401 7 2 2 1398 1400
0 1402 5 1 1 3254
0 1403 7 1 2 3253 1402
0 1404 5 2 1 1403
0 1405 7 2 2 2009 2069
0 1406 5 1 1 3258
0 1407 7 1 2 1382 1384
0 1408 5 1 1 1407
0 1409 7 2 2 3246 1408
0 1410 5 1 1 3260
0 1411 7 1 2 3259 3261
0 1412 5 2 1 1411
0 1413 7 1 2 1406 1410
0 1414 5 1 1 1413
0 1415 7 2 2 3262 1414
0 1416 5 1 1 3264
0 1417 7 2 2 1988 2081
0 1418 5 1 1 3266
0 1419 7 2 2 1999 2070
0 1420 5 1 1 3268
0 1421 7 2 2 3267 3269
0 1422 5 2 1 3270
0 1423 7 1 2 3265 3271
0 1424 5 2 1 1423
0 1425 7 2 2 3263 3274
0 1426 5 1 1 3276
0 1427 7 1 2 1394 3255
0 1428 5 1 1 1427
0 1429 7 2 2 3256 1428
0 1430 5 1 1 3278
0 1431 7 1 2 1426 3279
0 1432 5 2 1 1431
0 1433 7 2 2 3257 3280
0 1434 5 1 1 3282
0 1435 7 1 2 1374 3249
0 1436 5 1 1 1435
0 1437 7 2 2 3250 1436
0 1438 5 1 1 3284
0 1439 7 1 2 1434 3285
0 1440 5 2 1 1439
0 1441 7 2 2 3251 3286
0 1442 5 1 1 3288
0 1443 7 1 2 3226 1368
0 1444 5 1 1 1443
0 1445 7 2 2 3229 1444
0 1446 5 1 1 3290
0 1447 7 1 2 1442 3291
0 1448 5 2 1 1447
0 1449 7 2 2 3230 3292
0 1450 5 1 1 3294
0 1451 7 1 2 3208 1344
0 1452 5 1 1 1451
0 1453 7 2 2 3211 1452
0 1454 5 1 1 3296
0 1455 7 1 2 1450 3297
0 1456 5 2 1 1455
0 1457 7 2 2 3212 3298
0 1458 5 1 1 3300
0 1459 7 1 2 3178 1302
0 1460 5 1 1 1459
0 1461 7 2 2 3181 1460
0 1462 5 1 1 3302
0 1463 7 1 2 1458 3303
0 1464 5 2 1 1463
0 1465 7 2 2 3182 3304
0 1466 5 1 1 3306
0 1467 7 1 2 3136 1246
0 1468 5 1 1 1467
0 1469 7 2 2 3139 1468
0 1470 5 1 1 3308
0 1471 7 1 2 1466 3309
0 1472 5 2 1 1471
0 1473 7 2 2 3140 3310
0 1474 5 1 1 3312
0 1475 7 1 2 3094 1186
0 1476 5 1 1 1475
0 1477 7 2 2 3097 1476
0 1478 5 1 1 3314
0 1479 7 1 2 1474 3315
0 1480 5 2 1 1479
0 1481 7 2 2 3098 3316
0 1482 5 1 1 3318
0 1483 7 1 2 3040 1116
0 1484 5 1 1 1483
0 1485 7 2 2 3043 1484
0 1486 5 1 1 3320
0 1487 7 1 2 1482 3321
0 1488 5 2 1 1487
0 1489 7 2 2 3044 3322
0 1490 5 1 1 3324
0 1491 7 1 2 2966 1032
0 1492 5 1 1 1491
0 1493 7 2 2 2969 1492
0 1494 5 1 1 3326
0 1495 7 1 2 1490 3327
0 1496 5 2 1 1495
0 1497 7 2 2 2970 3328
0 1498 5 1 1 3330
0 1499 7 1 2 2888 926
0 1500 5 1 1 1499
0 1501 7 2 2 2891 1500
0 1502 5 1 1 3332
0 1503 7 1 2 1498 3333
0 1504 5 2 1 1503
0 1505 7 2 2 2892 3334
0 1506 5 1 1 3336
0 1507 7 1 2 2801 834
0 1508 5 1 1 1507
0 1509 7 2 2 2815 1508
0 1510 5 1 1 3338
0 1511 7 1 2 1506 3339
0 1512 5 2 1 1511
0 1513 7 2 2 2816 3340
0 1514 5 1 1 3342
0 1515 7 2 2 2061 2142
0 1516 5 1 1 3344
0 1517 7 1 2 2755 2811
0 1518 5 1 1 1517
0 1519 7 1 2 3345 1518
0 1520 5 2 1 1519
0 1521 7 1 2 2812 1516
0 1522 5 1 1 1521
0 1523 7 2 2 3346 1522
0 1524 5 1 1 3348
0 1525 7 1 2 1514 3349
0 1526 5 2 1 1525
0 1527 7 1 2 3343 1524
0 1528 5 1 1 1527
0 1529 7 2 2 3350 1528
0 1530 5 1 1 3352
0 1531 7 1 2 2189 1530
0 1532 5 3 1 1531
0 1533 7 2 2 3347 3351
0 1534 5 1 1 3357
0 1535 7 2 2 2193 3358
0 1536 5 1 1 3359
0 1537 7 2 2 3354 1536
0 1538 5 1 1 3361
0 1539 7 2 2 2270 1534
0 1540 5 2 1 3363
0 1541 7 1 2 1538 3365
0 1542 5 1 1 1541
0 1543 7 1 2 3337 1510
0 1544 5 1 1 1543
0 1545 7 2 2 3341 1544
0 1546 5 1 1 3367
0 1547 7 1 2 2185 1546
0 1548 5 3 1 1547
0 1549 7 1 2 2266 3368
0 1550 5 4 1 1549
0 1551 7 1 2 3331 1502
0 1552 5 1 1 1551
0 1553 7 2 2 3335 1552
0 1554 5 1 1 3376
0 1555 7 1 2 2182 1554
0 1556 5 4 1 1555
0 1557 7 1 2 2263 3377
0 1558 5 3 1 1557
0 1559 7 1 2 3325 1494
0 1560 5 1 1 1559
0 1561 7 2 2 3329 1560
0 1562 5 1 1 3385
0 1563 7 1 2 2178 1562
0 1564 5 4 1 1563
0 1565 7 1 2 2259 3386
0 1566 5 4 1 1565
0 1567 7 1 2 3319 1486
0 1568 5 1 1 1567
0 1569 7 2 2 3323 1568
0 1570 5 1 1 3395
0 1571 7 1 2 2175 1570
0 1572 5 3 1 1571
0 1573 7 1 2 2256 3396
0 1574 5 3 1 1573
0 1575 7 1 2 3313 1478
0 1576 5 1 1 1575
0 1577 7 2 2 3317 1576
0 1578 5 1 1 3403
0 1579 7 1 2 2253 3404
0 1580 5 3 1 1579
0 1581 7 2 2 3400 3405
0 1582 7 2 2 2172 1578
0 1583 5 4 1 3410
0 1584 7 1 2 3307 1470
0 1585 5 1 1 1584
0 1586 7 2 2 3311 1585
0 1587 5 1 1 3416
0 1588 7 1 2 2169 1587
0 1589 5 3 1 1588
0 1590 7 1 2 2250 3417
0 1591 5 4 1 1590
0 1592 7 1 2 3301 1462
0 1593 5 1 1 1592
0 1594 7 2 2 3305 1593
0 1595 5 1 1 3425
0 1596 7 1 2 2166 1595
0 1597 5 3 1 1596
0 1598 7 1 2 2247 3426
0 1599 5 4 1 1598
0 1600 7 1 2 3295 1454
0 1601 5 1 1 1600
0 1602 7 2 2 3299 1601
0 1603 5 1 1 3434
0 1604 7 1 2 2163 1603
0 1605 5 3 1 1604
0 1606 7 1 2 2244 3435
0 1607 5 4 1 1606
0 1608 7 1 2 3289 1446
0 1609 5 1 1 1608
0 1610 7 2 2 3293 1609
0 1611 5 1 1 3443
0 1612 7 1 2 2160 1611
0 1613 5 4 1 1612
0 1614 7 1 2 2241 3444
0 1615 5 4 1 1614
0 1616 7 1 2 3283 1438
0 1617 5 1 1 1616
0 1618 7 2 2 3287 1617
0 1619 5 1 1 3453
0 1620 7 1 2 2157 1619
0 1621 5 4 1 1620
0 1622 7 1 2 2238 3454
0 1623 5 4 1 1622
0 1624 7 1 2 3277 1430
0 1625 5 1 1 1624
0 1626 7 2 2 3281 1625
0 1627 5 1 1 3463
0 1628 7 1 2 2154 1627
0 1629 5 4 1 1628
0 1630 7 1 2 2235 3464
0 1631 5 3 1 1630
0 1632 7 1 2 1416 3272
0 1633 5 1 1 1632
0 1634 7 2 2 3275 1633
0 1635 5 1 1 3472
0 1636 7 1 2 2232 3473
0 1637 5 3 1 1636
0 1638 7 1 2 2151 1635
0 1639 5 4 1 1638
0 1640 7 1 2 1418 1420
0 1641 5 1 1 1640
0 1642 7 2 2 3273 1641
0 1643 5 1 1 3481
0 1644 7 1 2 2229 3482
0 1645 5 2 1 1644
0 1646 7 1 2 2148 1643
0 1647 5 2 1 1646
0 1648 7 2 2 1989 2071
0 1649 5 1 1 3487
0 1650 7 1 2 2145 1649
0 1651 5 1 1 1650
0 1652 7 2 2 3485 1651
0 1653 5 1 1 3489
0 1654 7 1 2 3483 1653
0 1655 5 3 1 1654
0 1656 7 1 2 3477 3491
0 1657 5 1 1 1656
0 1658 7 3 2 3474 1657
0 1659 5 1 1 3494
0 1660 7 1 2 3469 3495
0 1661 5 1 1 1660
0 1662 7 2 2 3465 1661
0 1663 5 1 1 3497
0 1664 7 2 2 3459 1663
0 1665 5 1 1 3499
0 1666 7 2 2 3455 1665
0 1667 5 2 1 3501
0 1668 7 1 2 3449 3503
0 1669 5 1 1 1668
0 1670 7 2 2 3445 1669
0 1671 5 2 1 3505
0 1672 7 1 2 3439 3507
0 1673 5 1 1 1672
0 1674 7 2 2 3436 1673
0 1675 5 2 1 3509
0 1676 7 1 2 3430 3511
0 1677 5 1 1 1676
0 1678 7 2 2 3427 1677
0 1679 5 2 1 3513
0 1680 7 1 2 3421 3515
0 1681 5 1 1 1680
0 1682 7 3 2 3418 1681
0 1683 5 1 1 3517
0 1684 7 1 2 3412 3518
0 1685 5 1 1 1684
0 1686 7 1 2 3408 1685
0 1687 5 1 1 1686
0 1688 7 2 2 3397 1687
0 1689 5 1 1 3520
0 1690 7 2 2 3391 1689
0 1691 5 1 1 3522
0 1692 7 1 2 3387 1691
0 1693 5 1 1 1692
0 1694 7 1 2 3382 1693
0 1695 5 1 1 1694
0 1696 7 2 2 3378 1695
0 1697 5 2 1 3524
0 1698 7 1 2 3372 3526
0 1699 5 1 1 1698
0 1700 7 2 2 3369 1699
0 1701 5 2 1 3528
0 1702 7 1 2 2268 3353
0 1703 5 3 1 1702
0 1704 7 2 2 3532 3366
0 1705 7 1 2 3530 3535
0 1706 5 1 1 1705
0 1707 7 3 2 1542 1706
0 1708 5 1 1 3537
0 1709 7 1 2 3533 3360
0 1710 5 1 1 1709
0 1711 7 2 2 3392 3383
0 1712 7 1 2 2226 3488
0 1713 5 1 1 1712
0 1714 7 3 2 3484 1713
0 1715 5 2 1 3542
0 1716 7 2 2 3486 3545
0 1717 7 1 2 3478 3547
0 1718 5 1 1 1717
0 1719 7 2 2 3470 3475
0 1720 7 2 2 1718 3549
0 1721 5 1 1 3551
0 1722 7 2 2 3466 1721
0 1723 5 2 1 3553
0 1724 7 1 2 3460 3555
0 1725 5 1 1 1724
0 1726 7 2 2 3456 1725
0 1727 5 1 1 3557
0 1728 7 2 2 3450 1727
0 1729 5 1 1 3559
0 1730 7 2 2 3446 1729
0 1731 5 2 1 3561
0 1732 7 1 2 3440 3563
0 1733 5 1 1 1732
0 1734 7 2 2 3437 1733
0 1735 5 2 1 3565
0 1736 7 1 2 3431 3567
0 1737 5 1 1 1736
0 1738 7 2 2 3428 1737
0 1739 5 2 1 3569
0 1740 7 1 2 3422 3571
0 1741 5 1 1 1740
0 1742 7 2 2 3419 1741
0 1743 5 2 1 3573
0 1744 7 1 2 3406 3575
0 1745 5 1 1 1744
0 1746 7 2 2 3413 1745
0 1747 5 2 1 3577
0 1748 7 1 2 3401 3579
0 1749 5 1 1 1748
0 1750 7 3 2 3398 1749
0 1751 5 2 1 3581
0 1752 7 1 2 3582 3388
0 1753 5 1 1 1752
0 1754 7 2 2 3540 1753
0 1755 5 1 1 3586
0 1756 7 2 2 3379 1755
0 1757 5 2 1 3588
0 1758 7 3 2 3370 3373
0 1759 5 2 1 3592
0 1760 7 1 2 3589 3593
0 1761 5 1 1 1760
0 1762 7 2 2 3393 3389
0 1763 5 2 1 3597
0 1764 7 1 2 3584 3599
0 1765 5 1 1 1764
0 1766 7 1 2 3583 3598
0 1767 5 1 1 1766
0 1768 7 3 2 3399 3402
0 1769 5 2 1 3601
0 1770 7 1 2 3578 3602
0 1771 5 1 1 1770
0 1772 7 1 2 3580 3604
0 1773 5 1 1 1772
0 1774 7 3 2 3414 3407
0 1775 5 2 1 3606
0 1776 7 1 2 3576 3607
0 1777 5 1 1 1776
0 1778 7 1 2 3574 3609
0 1779 5 1 1 1778
0 1780 7 1 2 1777 1779
0 1781 5 1 1 1780
0 1782 7 3 2 3420 3423
0 1783 5 2 1 3611
0 1784 7 1 2 3572 3612
0 1785 5 1 1 1784
0 1786 7 3 2 3429 3432
0 1787 5 2 1 3616
0 1788 7 1 2 3566 3619
0 1789 5 1 1 1788
0 1790 7 1 2 3568 3617
0 1791 5 1 1 1790
0 1792 7 1 2 1789 1791
0 1793 5 1 1 1792
0 1794 7 3 2 3438 3441
0 1795 5 2 1 3621
0 1796 7 1 2 3562 3622
0 1797 5 1 1 1796
0 1798 7 1 2 3447 3560
0 1799 5 1 1 1798
0 1800 7 2 2 3448 3451
0 1801 5 2 1 3626
0 1802 7 1 2 3558 3628
0 1803 5 1 1 1802
0 1804 7 2 2 3457 3461
0 1805 5 2 1 3630
0 1806 7 1 2 3554 3631
0 1807 5 1 1 1806
0 1808 7 1 2 3467 3552
0 1809 5 1 1 1808
0 1810 7 2 2 3468 3471
0 1811 5 2 1 3634
0 1812 7 1 2 3479 3636
0 1813 5 1 1 1812
0 1814 7 2 2 3480 3476
0 1815 5 2 1 3638
0 1816 7 1 2 3548 3640
0 1817 5 1 1 1816
0 1818 7 1 2 3543 3490
0 1819 5 1 1 1818
0 1820 7 1 2 1817 1819
0 1821 7 1 2 1813 1820
0 1822 7 1 2 1809 1821
0 1823 5 1 1 1822
0 1824 7 1 2 3556 3632
0 1825 5 1 1 1824
0 1826 7 1 2 1823 1825
0 1827 7 1 2 1807 1826
0 1828 5 1 1 1827
0 1829 7 1 2 1803 1828
0 1830 7 1 2 1799 1829
0 1831 5 1 1 1830
0 1832 7 1 2 3564 3624
0 1833 5 1 1 1832
0 1834 7 1 2 1831 1833
0 1835 7 1 2 1797 1834
0 1836 7 1 2 1793 1835
0 1837 5 1 1 1836
0 1838 7 1 2 3570 3614
0 1839 5 1 1 1838
0 1840 7 1 2 1837 1839
0 1841 7 1 2 1785 1840
0 1842 5 1 1 1841
0 1843 7 1 2 1781 1842
0 1844 7 1 2 1773 1843
0 1845 7 1 2 1771 1844
0 1846 7 1 2 1767 1845
0 1847 7 1 2 1765 1846
0 1848 7 1 2 1761 1847
0 1849 7 1 2 3590 3595
0 1850 5 1 1 1849
0 1851 7 1 2 3394 3585
0 1852 5 1 1 1851
0 1853 7 2 2 3380 3384
0 1854 5 1 1 3642
0 1855 7 2 2 3390 1854
0 1856 5 1 1 3644
0 1857 7 1 2 1852 3645
0 1858 5 1 1 1857
0 1859 7 1 2 3381 3587
0 1860 5 1 1 1859
0 1861 7 1 2 1858 1860
0 1862 5 1 1 1861
0 1863 7 1 2 1850 1862
0 1864 7 1 2 1848 1863
0 1865 7 1 2 1710 1864
0 1866 7 1 2 3591 3374
0 1867 5 1 1 1866
0 1868 7 2 2 3371 1867
0 1869 5 1 1 3646
0 1870 7 2 2 3534 3355
0 1871 5 2 1 3648
0 1872 7 1 2 1869 3650
0 1873 5 1 1 1872
0 1874 7 1 2 3647 3362
0 1875 5 1 1 1874
0 1876 7 1 2 1873 1875
0 1877 7 1 2 1865 1876
0 1878 7 1 2 1708 1877
0 1879 5 1 1 1878
0 1880 7 1 2 3356 3364
0 1881 5 1 1 1880
0 1882 7 1 2 3596 3525
0 1883 5 1 1 1882
0 1884 7 1 2 3594 3527
0 1885 5 1 1 1884
0 1886 7 1 2 3643 3523
0 1887 5 1 1 1886
0 1888 7 1 2 3600 3521
0 1889 5 1 1 1888
0 1890 7 1 2 3411 3603
0 1891 5 1 1 1890
0 1892 7 1 2 3415 3605
0 1893 5 1 1 1892
0 1894 7 1 2 3610 1683
0 1895 5 1 1 1894
0 1896 7 1 2 3608 3519
0 1897 5 1 1 1896
0 1898 7 1 2 1895 1897
0 1899 5 1 1 1898
0 1900 7 1 2 3620 3510
0 1901 5 1 1 1900
0 1902 7 1 2 3618 3512
0 1903 5 1 1 1902
0 1904 7 1 2 3625 3506
0 1905 5 1 1 1904
0 1906 7 1 2 3627 3502
0 1907 5 1 1 1906
0 1908 7 1 2 3458 3500
0 1909 5 1 1 1908
0 1910 7 1 2 3633 3498
0 1911 5 1 1 1910
0 1912 7 1 2 3637 3496
0 1913 5 1 1 1912
0 1914 7 1 2 3635 1659
0 1915 5 1 1 1914
0 1916 7 1 2 3639 3492
0 1917 5 1 1 1916
0 1918 7 1 2 3546 3493
0 1919 5 1 1 1918
0 1920 7 1 2 3641 1919
0 1921 5 1 1 1920
0 1922 7 1 2 1917 1921
0 1923 7 1 2 1915 1922
0 1924 7 1 2 1913 1923
0 1925 5 1 1 1924
0 1926 7 1 2 1911 1925
0 1927 7 1 2 1909 1926
0 1928 5 1 1 1927
0 1929 7 1 2 3629 3504
0 1930 5 1 1 1929
0 1931 7 1 2 1928 1930
0 1932 7 1 2 1907 1931
0 1933 5 1 1 1932
0 1934 7 1 2 3623 3508
0 1935 5 1 1 1934
0 1936 7 1 2 1933 1935
0 1937 7 1 2 1905 1936
0 1938 7 1 2 1903 1937
0 1939 7 1 2 1901 1938
0 1940 5 1 1 1939
0 1941 7 1 2 3613 3516
0 1942 5 1 1 1941
0 1943 7 1 2 3615 3514
0 1944 5 1 1 1943
0 1945 7 1 2 1942 1944
0 1946 5 1 1 1945
0 1947 7 1 2 1940 1946
0 1948 5 1 1 1947
0 1949 7 1 2 1899 1948
0 1950 7 1 2 1893 1949
0 1951 7 1 2 1891 1950
0 1952 7 1 2 1889 1951
0 1953 7 1 2 1856 1952
0 1954 7 1 2 1887 1953
0 1955 7 1 2 1885 1954
0 1956 7 1 2 1883 1955
0 1957 7 1 2 1881 1956
0 1958 7 1 2 3651 3529
0 1959 5 1 1 1958
0 1960 7 1 2 3649 3531
0 1961 5 1 1 1960
0 1962 7 1 2 1959 1961
0 1963 7 1 2 1957 1962
0 1964 7 1 2 3538 1963
0 1965 5 1 1 1964
0 1966 7 1 2 1879 1965
0 1967 7 1 2 2737 1966
0 1968 5 1 1 1967
0 1969 7 1 2 3544 3550
0 1970 7 1 2 3462 1969
0 1971 7 1 2 3452 1970
0 1972 7 1 2 3442 1971
0 1973 7 1 2 3433 1972
0 1974 7 1 2 3424 1973
0 1975 7 1 2 3409 1974
0 1976 7 1 2 3541 1975
0 1977 7 1 2 3375 1976
0 1978 7 1 2 3536 1977
0 1979 7 1 2 3539 1978
0 1980 5 1 1 1979
0 1981 7 1 2 740 1980
0 1982 5 1 1 1981
3 4099 7 0 2 1968 1982
