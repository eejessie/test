1 0 0 8 0
2 32 1 0
2 1259 1 0
2 1260 1 0
2 1261 1 0
2 1262 1 0
2 1263 1 0
2 1264 1 0
2 1265 1 0
1 1 0 8 0
2 1266 1 1
2 1267 1 1
2 1268 1 1
2 1269 1 1
2 1270 1 1
2 1271 1 1
2 1272 1 1
2 1273 1 1
1 2 0 8 0
2 1274 1 2
2 1275 1 2
2 1276 1 2
2 1277 1 2
2 1278 1 2
2 1279 1 2
2 1280 1 2
2 1281 1 2
1 3 0 9 0
2 1282 1 3
2 1283 1 3
2 1284 1 3
2 1285 1 3
2 1286 1 3
2 1287 1 3
2 1288 1 3
2 1289 1 3
2 1290 1 3
1 4 0 8 0
2 1291 1 4
2 1292 1 4
2 1293 1 4
2 1294 1 4
2 1295 1 4
2 1296 1 4
2 1297 1 4
2 1298 1 4
1 5 0 9 0
2 1299 1 5
2 1300 1 5
2 1301 1 5
2 1302 1 5
2 1303 1 5
2 1304 1 5
2 1305 1 5
2 1306 1 5
2 1307 1 5
1 6 0 8 0
2 1308 1 6
2 1309 1 6
2 1310 1 6
2 1311 1 6
2 1312 1 6
2 1313 1 6
2 1314 1 6
2 1315 1 6
1 7 0 8 0
2 1316 1 7
2 1317 1 7
2 1318 1 7
2 1319 1 7
2 1320 1 7
2 1321 1 7
2 1322 1 7
2 1323 1 7
1 8 0 8 0
2 1324 1 8
2 1325 1 8
2 1326 1 8
2 1327 1 8
2 1328 1 8
2 1329 1 8
2 1330 1 8
2 1331 1 8
1 9 0 8 0
2 1332 1 9
2 1333 1 9
2 1334 1 9
2 1335 1 9
2 1336 1 9
2 1337 1 9
2 1338 1 9
2 1339 1 9
1 10 0 9 0
2 1340 1 10
2 1341 1 10
2 1342 1 10
2 1343 1 10
2 1344 1 10
2 1345 1 10
2 1346 1 10
2 1347 1 10
2 1348 1 10
1 11 0 8 0
2 1349 1 11
2 1350 1 11
2 1351 1 11
2 1352 1 11
2 1353 1 11
2 1354 1 11
2 1355 1 11
2 1356 1 11
1 12 0 8 0
2 1357 1 12
2 1358 1 12
2 1359 1 12
2 1360 1 12
2 1361 1 12
2 1362 1 12
2 1363 1 12
2 1364 1 12
1 13 0 8 0
2 1365 1 13
2 1366 1 13
2 1367 1 13
2 1368 1 13
2 1369 1 13
2 1370 1 13
2 1371 1 13
2 1372 1 13
1 14 0 8 0
2 1373 1 14
2 1374 1 14
2 1375 1 14
2 1376 1 14
2 1377 1 14
2 1378 1 14
2 1379 1 14
2 1380 1 14
1 15 0 8 0
2 1381 1 15
2 1382 1 15
2 1383 1 15
2 1384 1 15
2 1385 1 15
2 1386 1 15
2 1387 1 15
2 1388 1 15
1 16 0 2 0
2 1389 1 16
2 1390 1 16
1 17 0 2 0
2 1391 1 17
2 1392 1 17
1 18 0 2 0
2 1393 1 18
2 1394 1 18
1 19 0 2 0
2 1395 1 19
2 1396 1 19
1 20 0 2 0
2 1397 1 20
2 1398 1 20
1 21 0 2 0
2 1399 1 21
2 1400 1 21
1 22 0 2 0
2 1401 1 22
2 1402 1 22
1 23 0 2 0
2 1403 1 23
2 1404 1 23
1 24 0 2 0
2 1405 1 24
2 1406 1 24
1 25 0 2 0
2 1407 1 25
2 1408 1 25
1 26 0 2 0
2 1409 1 26
2 1410 1 26
1 27 0 2 0
2 1411 1 27
2 1412 1 27
1 28 0 2 0
2 1413 1 28
2 1414 1 28
1 29 0 2 0
2 1415 1 29
2 1416 1 29
1 30 0 2 0
2 1417 1 30
2 1418 1 30
1 31 0 2 0
2 1419 1 31
2 1420 1 31
2 1421 1 49
2 1422 1 49
2 1423 1 51
2 1424 1 51
2 1425 1 52
2 1426 1 52
2 1427 1 53
2 1428 1 53
2 1429 1 55
2 1430 1 55
2 1431 1 58
2 1432 1 58
2 1433 1 61
2 1434 1 61
2 1435 1 64
2 1436 1 64
2 1437 1 65
2 1438 1 65
2 1439 1 67
2 1440 1 67
2 1441 1 69
2 1442 1 69
2 1443 1 75
2 1444 1 75
2 1445 1 78
2 1446 1 78
2 1447 1 78
2 1448 1 82
2 1449 1 82
2 1450 1 83
2 1451 1 83
2 1452 1 85
2 1453 1 85
2 1454 1 88
2 1455 1 88
2 1456 1 89
2 1457 1 89
2 1458 1 93
2 1459 1 93
2 1460 1 96
2 1461 1 96
2 1462 1 97
2 1463 1 97
2 1464 1 101
2 1465 1 101
2 1466 1 104
2 1467 1 104
2 1468 1 105
2 1469 1 105
2 1470 1 109
2 1471 1 109
2 1472 1 112
2 1473 1 112
2 1474 1 113
2 1475 1 113
2 1476 1 115
2 1477 1 115
2 1478 1 118
2 1479 1 118
2 1480 1 119
2 1481 1 119
2 1482 1 123
2 1483 1 123
2 1484 1 126
2 1485 1 126
2 1486 1 127
2 1487 1 127
2 1488 1 131
2 1489 1 131
2 1490 1 134
2 1491 1 134
2 1492 1 135
2 1493 1 135
2 1494 1 139
2 1495 1 139
2 1496 1 142
2 1497 1 142
2 1498 1 143
2 1499 1 143
2 1500 1 147
2 1501 1 147
2 1502 1 150
2 1503 1 150
2 1504 1 151
2 1505 1 151
2 1506 1 155
2 1507 1 155
2 1508 1 158
2 1509 1 158
2 1510 1 159
2 1511 1 159
2 1512 1 163
2 1513 1 163
2 1514 1 166
2 1515 1 166
2 1516 1 167
2 1517 1 167
2 1518 1 171
2 1519 1 171
2 1520 1 174
2 1521 1 174
2 1522 1 175
2 1523 1 175
2 1524 1 177
2 1525 1 177
2 1526 1 179
2 1527 1 179
2 1528 1 181
2 1529 1 181
2 1530 1 182
2 1531 1 182
2 1532 1 183
2 1533 1 183
2 1534 1 184
2 1535 1 184
2 1536 1 186
2 1537 1 186
2 1538 1 187
2 1539 1 187
2 1540 1 191
2 1541 1 191
2 1542 1 194
2 1543 1 194
2 1544 1 195
2 1545 1 195
2 1546 1 199
2 1547 1 199
2 1548 1 202
2 1549 1 202
2 1550 1 203
2 1551 1 203
2 1552 1 207
2 1553 1 207
2 1554 1 210
2 1555 1 210
2 1556 1 211
2 1557 1 211
2 1558 1 215
2 1559 1 215
2 1560 1 218
2 1561 1 218
2 1562 1 219
2 1563 1 219
2 1564 1 223
2 1565 1 223
2 1566 1 226
2 1567 1 226
2 1568 1 227
2 1569 1 227
2 1570 1 231
2 1571 1 231
2 1572 1 234
2 1573 1 234
2 1574 1 235
2 1575 1 235
2 1576 1 239
2 1577 1 239
2 1578 1 242
2 1579 1 242
2 1580 1 243
2 1581 1 243
2 1582 1 245
2 1583 1 245
2 1584 1 248
2 1585 1 248
2 1586 1 251
2 1587 1 251
2 1588 1 255
2 1589 1 255
2 1590 1 258
2 1591 1 258
2 1592 1 259
2 1593 1 259
2 1594 1 263
2 1595 1 263
2 1596 1 266
2 1597 1 266
2 1598 1 267
2 1599 1 267
2 1600 1 269
2 1601 1 269
2 1602 1 272
2 1603 1 272
2 1604 1 273
2 1605 1 273
2 1606 1 275
2 1607 1 275
2 1608 1 281
2 1609 1 281
2 1610 1 284
2 1611 1 284
2 1612 1 287
2 1613 1 287
2 1614 1 290
2 1615 1 290
2 1616 1 293
2 1617 1 293
2 1618 1 297
2 1619 1 297
2 1620 1 300
2 1621 1 300
2 1622 1 301
2 1623 1 301
2 1624 1 305
2 1625 1 305
2 1626 1 308
2 1627 1 308
2 1628 1 309
2 1629 1 309
2 1630 1 311
2 1631 1 311
2 1632 1 314
2 1633 1 314
2 1634 1 317
2 1635 1 317
2 1636 1 321
2 1637 1 321
2 1638 1 324
2 1639 1 324
2 1640 1 325
2 1641 1 325
2 1642 1 329
2 1643 1 329
2 1644 1 332
2 1645 1 332
2 1646 1 333
2 1647 1 333
2 1648 1 337
2 1649 1 337
2 1650 1 340
2 1651 1 340
2 1652 1 341
2 1653 1 341
2 1654 1 345
2 1655 1 345
2 1656 1 348
2 1657 1 348
2 1658 1 349
2 1659 1 349
2 1660 1 353
2 1661 1 353
2 1662 1 356
2 1663 1 356
2 1664 1 357
2 1665 1 357
2 1666 1 359
2 1667 1 359
2 1668 1 362
2 1669 1 362
2 1670 1 363
2 1671 1 363
2 1672 1 367
2 1673 1 367
2 1674 1 370
2 1675 1 370
2 1676 1 371
2 1677 1 371
2 1678 1 373
2 1679 1 373
2 1680 1 375
2 1681 1 375
2 1682 1 378
2 1683 1 378
2 1684 1 379
2 1685 1 379
2 1686 1 381
2 1687 1 381
2 1688 1 383
2 1689 1 383
2 1690 1 385
2 1691 1 385
2 1692 1 387
2 1693 1 387
2 1694 1 388
2 1695 1 388
2 1696 1 389
2 1697 1 389
2 1698 1 390
2 1699 1 390
2 1700 1 391
2 1701 1 391
2 1702 1 392
2 1703 1 392
2 1704 1 393
2 1705 1 393
2 1706 1 394
2 1707 1 394
2 1708 1 396
2 1709 1 396
2 1710 1 399
2 1711 1 399
2 1712 1 403
2 1713 1 403
2 1714 1 406
2 1715 1 406
2 1716 1 409
2 1717 1 409
2 1718 1 413
2 1719 1 413
2 1720 1 416
2 1721 1 416
2 1722 1 417
2 1723 1 417
2 1724 1 420
2 1725 1 420
2 1726 1 421
2 1727 1 421
2 1728 1 425
2 1729 1 425
2 1730 1 428
2 1731 1 428
2 1732 1 429
2 1733 1 429
2 1734 1 433
2 1735 1 433
2 1736 1 436
2 1737 1 436
2 1738 1 437
2 1739 1 437
2 1740 1 441
2 1741 1 441
2 1742 1 444
2 1743 1 444
2 1744 1 447
2 1745 1 447
2 1746 1 451
2 1747 1 451
2 1748 1 454
2 1749 1 454
2 1750 1 457
2 1751 1 457
2 1752 1 461
2 1753 1 461
2 1754 1 464
2 1755 1 464
2 1756 1 465
2 1757 1 465
2 1758 1 467
2 1759 1 467
2 1760 1 470
2 1761 1 470
2 1762 1 471
2 1763 1 471
2 1764 1 475
2 1765 1 475
2 1766 1 478
2 1767 1 478
2 1768 1 479
2 1769 1 479
2 1770 1 483
2 1771 1 483
2 1772 1 486
2 1773 1 486
2 1774 1 487
2 1775 1 487
2 1776 1 491
2 1777 1 491
2 1778 1 494
2 1779 1 494
2 1780 1 495
2 1781 1 495
2 1782 1 499
2 1783 1 499
2 1784 1 502
2 1785 1 502
2 1786 1 503
2 1787 1 503
2 1788 1 507
2 1789 1 507
2 1790 1 510
2 1791 1 510
2 1792 1 511
2 1793 1 511
2 1794 1 513
2 1795 1 513
2 1796 1 519
2 1797 1 519
2 1798 1 522
2 1799 1 522
2 1800 1 525
2 1801 1 525
2 1802 1 528
2 1803 1 528
2 1804 1 531
2 1805 1 531
2 1806 1 535
2 1807 1 535
2 1808 1 538
2 1809 1 538
2 1810 1 539
2 1811 1 539
2 1812 1 543
2 1813 1 543
2 1814 1 546
2 1815 1 546
2 1816 1 547
2 1817 1 547
2 1818 1 551
2 1819 1 551
2 1820 1 554
2 1821 1 554
2 1822 1 555
2 1823 1 555
2 1824 1 559
2 1825 1 559
2 1826 1 562
2 1827 1 562
2 1828 1 563
2 1829 1 563
2 1830 1 567
2 1831 1 567
2 1832 1 570
2 1833 1 570
2 1834 1 571
2 1835 1 571
2 1836 1 575
2 1837 1 575
2 1838 1 578
2 1839 1 578
2 1840 1 579
2 1841 1 579
2 1842 1 583
2 1843 1 583
2 1844 1 586
2 1845 1 586
2 1846 1 587
2 1847 1 587
2 1848 1 589
2 1849 1 589
2 1850 1 592
2 1851 1 592
2 1852 1 595
2 1853 1 595
2 1854 1 599
2 1855 1 599
2 1856 1 602
2 1857 1 602
2 1858 1 603
2 1859 1 603
2 1860 1 607
2 1861 1 607
2 1862 1 610
2 1863 1 610
2 1864 1 611
2 1865 1 611
2 1866 1 615
2 1867 1 615
2 1868 1 618
2 1869 1 618
2 1870 1 619
2 1871 1 619
2 1872 1 623
2 1873 1 623
2 1874 1 626
2 1875 1 626
2 1876 1 627
2 1877 1 627
2 1878 1 633
2 1879 1 633
2 1880 1 636
2 1881 1 636
2 1882 1 637
2 1883 1 637
2 1884 1 641
2 1885 1 641
2 1886 1 644
2 1887 1 644
2 1888 1 645
2 1889 1 645
2 1890 1 649
2 1891 1 649
2 1892 1 652
2 1893 1 652
2 1894 1 653
2 1895 1 653
2 1896 1 657
2 1897 1 657
2 1898 1 660
2 1899 1 660
2 1900 1 661
2 1901 1 661
2 1902 1 663
2 1903 1 663
2 1904 1 666
2 1905 1 666
2 1906 1 669
2 1907 1 669
2 1908 1 673
2 1909 1 673
2 1910 1 676
2 1911 1 676
2 1912 1 677
2 1913 1 677
2 1914 1 681
2 1915 1 681
2 1916 1 684
2 1917 1 684
2 1918 1 687
2 1919 1 687
2 1920 1 689
2 1921 1 689
2 1922 1 691
2 1923 1 691
2 1924 1 693
2 1925 1 693
2 1926 1 695
2 1927 1 695
2 1928 1 697
2 1929 1 697
2 1930 1 699
2 1931 1 699
2 1932 1 700
2 1933 1 700
2 1934 1 701
2 1935 1 701
2 1936 1 701
2 1937 1 704
2 1938 1 704
2 1939 1 707
2 1940 1 707
2 1941 1 715
2 1942 1 715
2 1943 1 718
2 1944 1 718
2 1945 1 719
2 1946 1 719
2 1947 1 723
2 1948 1 723
2 1949 1 726
2 1950 1 726
2 1951 1 729
2 1952 1 729
2 1953 1 731
2 1954 1 731
2 1955 1 733
2 1956 1 733
2 1957 1 735
2 1958 1 735
2 1959 1 736
2 1960 1 736
2 1961 1 738
2 1962 1 738
2 1963 1 739
2 1964 1 739
2 1965 1 743
2 1966 1 743
2 1967 1 746
2 1968 1 746
2 1969 1 747
2 1970 1 747
2 1971 1 751
2 1972 1 751
2 1973 1 754
2 1974 1 754
2 1975 1 755
2 1976 1 755
2 1977 1 759
2 1978 1 759
2 1979 1 762
2 1980 1 762
2 1981 1 763
2 1982 1 763
2 1983 1 767
2 1984 1 767
2 1985 1 770
2 1986 1 770
2 1987 1 771
2 1988 1 771
2 1989 1 775
2 1990 1 775
2 1991 1 778
2 1992 1 778
2 1993 1 779
2 1994 1 779
2 1995 1 783
2 1996 1 783
2 1997 1 786
2 1998 1 786
2 1999 1 787
2 2000 1 787
2 2001 1 791
2 2002 1 791
2 2003 1 794
2 2004 1 794
2 2005 1 795
2 2006 1 795
2 2007 1 799
2 2008 1 799
2 2009 1 802
2 2010 1 802
2 2011 1 803
2 2012 1 803
2 2013 1 807
2 2014 1 807
2 2015 1 810
2 2016 1 810
2 2017 1 811
2 2018 1 811
2 2019 1 815
2 2020 1 815
2 2021 1 818
2 2022 1 818
2 2023 1 819
2 2024 1 819
2 2025 1 823
2 2026 1 823
2 2027 1 826
2 2028 1 826
2 2029 1 827
2 2030 1 827
2 2031 1 831
2 2032 1 831
2 2033 1 834
2 2034 1 834
2 2035 1 835
2 2036 1 835
2 2037 1 837
2 2038 1 837
2 2039 1 838
2 2040 1 838
2 2041 1 839
2 2042 1 839
2 2043 1 840
2 2044 1 840
2 2045 1 843
2 2046 1 843
2 2047 1 846
2 2048 1 846
2 2049 1 846
2 2050 1 849
2 2051 1 849
2 2052 1 852
2 2053 1 852
2 2054 1 852
2 2055 1 854
2 2056 1 854
2 2057 1 854
2 2058 1 857
2 2059 1 857
2 2060 1 860
2 2061 1 860
2 2062 1 860
2 2063 1 860
2 2064 1 862
2 2065 1 862
2 2066 1 862
2 2067 1 865
2 2068 1 865
2 2069 1 868
2 2070 1 868
2 2071 1 868
2 2072 1 870
2 2073 1 870
2 2074 1 870
2 2075 1 870
2 2076 1 873
2 2077 1 873
2 2078 1 876
2 2079 1 876
2 2080 1 876
2 2081 1 876
2 2082 1 878
2 2083 1 878
2 2084 1 878
2 2085 1 881
2 2086 1 881
2 2087 1 884
2 2088 1 884
2 2089 1 884
2 2090 1 884
2 2091 1 886
2 2092 1 886
2 2093 1 886
2 2094 1 889
2 2095 1 889
2 2096 1 892
2 2097 1 892
2 2098 1 892
2 2099 1 892
2 2100 1 894
2 2101 1 894
2 2102 1 894
2 2103 1 897
2 2104 1 897
2 2105 1 900
2 2106 1 900
2 2107 1 900
2 2108 1 902
2 2109 1 902
2 2110 1 902
2 2111 1 905
2 2112 1 905
2 2113 1 908
2 2114 1 908
2 2115 1 908
2 2116 1 910
2 2117 1 910
2 2118 1 910
2 2119 1 913
2 2120 1 913
2 2121 1 916
2 2122 1 916
2 2123 1 916
2 2124 1 916
2 2125 1 916
2 2126 1 918
2 2127 1 918
2 2128 1 918
2 2129 1 918
2 2130 1 921
2 2131 1 921
2 2132 1 923
2 2133 1 923
2 2134 1 924
2 2135 1 924
2 2136 1 924
2 2137 1 925
2 2138 1 925
2 2139 1 926
2 2140 1 926
2 2141 1 926
2 2142 1 926
2 2143 1 929
2 2144 1 929
2 2145 1 932
2 2146 1 932
2 2147 1 932
2 2148 1 934
2 2149 1 934
2 2150 1 934
2 2151 1 937
2 2152 1 937
2 2153 1 940
2 2154 1 940
2 2155 1 940
2 2156 1 940
2 2157 1 942
2 2158 1 942
2 2159 1 942
2 2160 1 945
2 2161 1 945
2 2162 1 948
2 2163 1 948
2 2164 1 950
2 2165 1 950
2 2166 1 951
2 2167 1 951
2 2168 1 956
2 2169 1 956
2 2170 1 961
2 2171 1 961
2 2172 1 964
2 2173 1 964
2 2174 1 964
2 2175 1 971
2 2176 1 971
2 2177 1 975
2 2178 1 975
2 2179 1 976
2 2180 1 976
2 2181 1 979
2 2182 1 979
2 2183 1 980
2 2184 1 980
2 2185 1 983
2 2186 1 983
2 2187 1 986
2 2188 1 986
2 2189 1 990
2 2190 1 990
2 2191 1 998
2 2192 1 998
2 2193 1 1001
2 2194 1 1001
2 2195 1 1002
2 2196 1 1002
2 2197 1 1004
2 2198 1 1004
2 2199 1 1004
2 2200 1 1007
2 2201 1 1007
2 2202 1 1011
2 2203 1 1011
2 2204 1 1013
2 2205 1 1013
2 2206 1 1013
2 2207 1 1014
2 2208 1 1014
2 2209 1 1023
2 2210 1 1023
2 2211 1 1023
2 2212 1 1024
2 2213 1 1024
2 2214 1 1029
2 2215 1 1029
2 2216 1 1030
2 2217 1 1030
2 2218 1 1033
2 2219 1 1033
2 2220 1 1033
2 2221 1 1039
2 2222 1 1039
2 2223 1 1039
2 2224 1 1045
2 2225 1 1045
2 2226 1 1046
2 2227 1 1046
2 2228 1 1049
2 2229 1 1049
2 2230 1 1050
2 2231 1 1050
2 2232 1 1059
2 2233 1 1059
2 2234 1 1059
2 2235 1 1059
2 2236 1 1060
2 2237 1 1060
2 2238 1 1071
2 2239 1 1071
2 2240 1 1071
2 2241 1 1072
2 2242 1 1072
2 2243 1 1078
2 2244 1 1078
2 2245 1 1083
2 2246 1 1083
2 2247 1 1084
2 2248 1 1084
2 2249 1 1086
2 2250 1 1086
2 2251 1 1094
2 2252 1 1094
2 2253 1 1094
2 2254 1 1095
2 2255 1 1095
2 2256 1 1116
2 2257 1 1116
2 2258 1 1117
2 2259 1 1117
2 2260 1 1120
2 2261 1 1120
2 2262 1 1123
2 2263 1 1123
2 2264 1 1129
2 2265 1 1129
2 2266 1 1132
2 2267 1 1132
2 2268 1 1133
2 2269 1 1133
2 2270 1 1136
2 2271 1 1136
2 2272 1 1138
2 2273 1 1138
2 2274 1 1140
2 2275 1 1140
2 2276 1 1141
2 2277 1 1141
2 2278 1 1144
2 2279 1 1144
2 2280 1 1145
2 2281 1 1145
2 2282 1 1148
2 2283 1 1148
2 2284 1 1149
2 2285 1 1149
2 2286 1 1152
2 2287 1 1152
2 2288 1 1153
2 2289 1 1153
2 2290 1 1156
2 2291 1 1156
2 2292 1 1157
2 2293 1 1157
2 2294 1 1160
2 2295 1 1160
2 2296 1 1161
2 2297 1 1161
2 2298 1 1164
2 2299 1 1164
0 33 5 1 1 1389
0 34 5 1 1 1391
0 35 5 1 1 1393
0 36 5 1 1 1395
0 37 5 1 1 1397
0 38 5 1 1 1399
0 39 5 1 1 1401
0 40 5 1 1 1403
0 41 5 1 1 1405
0 42 5 1 1 1407
0 43 5 1 1 1409
0 44 5 1 1 1411
0 45 5 1 1 1413
0 46 5 1 1 1415
0 47 5 1 1 1417
0 48 5 1 1 1419
0 49 7 2 2 1316 1381
0 50 5 1 1 1421
0 51 7 2 2 1308 1373
0 52 5 2 1 1423
0 53 7 2 2 1299 1382
0 54 5 1 1 1427
0 55 7 2 2 1317 1365
0 56 5 1 1 1429
0 57 7 1 2 1428 1430
0 58 5 2 1 57
0 59 7 1 2 54 56
0 60 5 1 1 59
0 61 7 2 2 1431 60
0 62 5 1 1 1433
0 63 7 1 2 1424 1434
0 64 5 2 1 63
0 65 7 2 2 1432 1435
0 66 5 1 1 1437
0 67 7 2 2 1309 1383
0 68 5 1 1 1439
0 69 7 2 2 1318 1374
0 70 5 1 1 1441
0 71 7 1 2 68 1442
0 72 5 1 1 71
0 73 7 1 2 1440 70
0 74 5 1 1 73
0 75 7 2 2 72 74
0 76 5 1 1 1443
0 77 7 1 2 66 76
0 78 5 3 1 77
0 79 7 1 2 1425 1445
0 80 5 1 1 79
0 81 7 1 2 1422 80
0 82 5 2 1 81
0 83 7 2 2 1291 1384
0 84 5 1 1 1450
0 85 7 2 2 1319 1357
0 86 5 1 1 1452
0 87 7 1 2 1451 1453
0 88 5 2 1 87
0 89 7 2 2 1310 1366
0 90 5 1 1 1456
0 91 7 1 2 84 86
0 92 5 1 1 91
0 93 7 2 2 1454 92
0 94 5 1 1 1458
0 95 7 1 2 1457 1459
0 96 5 2 1 95
0 97 7 2 2 1455 1460
0 98 5 1 1 1462
0 99 7 1 2 1426 62
0 100 5 1 1 99
0 101 7 2 2 1436 100
0 102 5 1 1 1464
0 103 7 1 2 98 1465
0 104 5 2 1 103
0 105 7 2 2 1300 1375
0 106 5 1 1 1468
0 107 7 1 2 90 94
0 108 5 1 1 107
0 109 7 2 2 1461 108
0 110 5 1 1 1470
0 111 7 1 2 1469 1471
0 112 5 2 1 111
0 113 7 2 2 1282 1385
0 114 5 1 1 1474
0 115 7 2 2 1320 1349
0 116 5 1 1 1476
0 117 7 1 2 1475 1477
0 118 5 2 1 117
0 119 7 2 2 1311 1358
0 120 5 1 1 1480
0 121 7 1 2 114 116
0 122 5 1 1 121
0 123 7 2 2 1478 122
0 124 5 1 1 1482
0 125 7 1 2 1481 1483
0 126 5 2 1 125
0 127 7 2 2 1479 1484
0 128 5 1 1 1486
0 129 7 1 2 106 110
0 130 5 1 1 129
0 131 7 2 2 1472 130
0 132 5 1 1 1488
0 133 7 1 2 128 1489
0 134 5 2 1 133
0 135 7 2 2 1473 1490
0 136 5 1 1 1492
0 137 7 1 2 1463 102
0 138 5 1 1 137
0 139 7 2 2 1466 138
0 140 5 1 1 1494
0 141 7 1 2 136 1495
0 142 5 2 1 141
0 143 7 2 2 1467 1496
0 144 5 1 1 1498
0 145 7 1 2 1438 1444
0 146 5 1 1 145
0 147 7 2 2 1446 146
0 148 5 1 1 1500
0 149 7 1 2 144 1501
0 150 5 2 1 149
0 151 7 2 2 1292 1376
0 152 5 1 1 1504
0 153 7 1 2 120 124
0 154 5 1 1 153
0 155 7 2 2 1485 154
0 156 5 1 1 1506
0 157 7 1 2 1505 1507
0 158 5 2 1 157
0 159 7 2 2 1301 1367
0 160 5 1 1 1510
0 161 7 1 2 152 156
0 162 5 1 1 161
0 163 7 2 2 1508 162
0 164 5 1 1 1512
0 165 7 1 2 1511 1513
0 166 5 2 1 165
0 167 7 2 2 1509 1514
0 168 5 1 1 1516
0 169 7 1 2 1487 132
0 170 5 1 1 169
0 171 7 2 2 1491 170
0 172 5 1 1 1518
0 173 7 1 2 168 1519
0 174 5 2 1 173
0 175 7 2 2 1274 1386
0 176 5 1 1 1522
0 177 7 2 2 1321 1324
0 178 5 1 1 1524
0 179 7 2 2 1312 1332
0 180 5 1 1 1526
0 181 7 2 2 1525 1527
0 182 5 2 1 1528
0 183 7 2 2 1340 1529
0 184 5 2 1 1532
0 185 7 1 2 1523 1533
0 186 5 2 1 185
0 187 7 2 2 1322 1341
0 188 5 1 1 1538
0 189 7 1 2 176 1534
0 190 5 1 1 189
0 191 7 2 2 1536 190
0 192 5 1 1 1540
0 193 7 1 2 1539 1541
0 194 5 2 1 193
0 195 7 2 2 1537 1542
0 196 5 1 1 1544
0 197 7 1 2 160 164
0 198 5 1 1 197
0 199 7 2 2 1515 198
0 200 5 1 1 1546
0 201 7 1 2 196 1547
0 202 5 2 1 201
0 203 7 2 2 1302 1359
0 204 5 1 1 1550
0 205 7 1 2 188 192
0 206 5 1 1 205
0 207 7 2 2 1543 206
0 208 5 1 1 1552
0 209 7 1 2 1551 1553
0 210 5 2 1 209
0 211 7 2 2 1313 1350
0 212 5 1 1 1556
0 213 7 1 2 204 208
0 214 5 1 1 213
0 215 7 2 2 1554 214
0 216 5 1 1 1558
0 217 7 1 2 1557 1559
0 218 5 2 1 217
0 219 7 2 2 1555 1560
0 220 5 1 1 1562
0 221 7 1 2 1545 200
0 222 5 1 1 221
0 223 7 2 2 1548 222
0 224 5 1 1 1564
0 225 7 1 2 220 1565
0 226 5 2 1 225
0 227 7 2 2 1549 1566
0 228 5 1 1 1568
0 229 7 1 2 1517 172
0 230 5 1 1 229
0 231 7 2 2 1520 230
0 232 5 1 1 1570
0 233 7 1 2 228 1571
0 234 5 2 1 233
0 235 7 2 2 1521 1572
0 236 5 1 1 1574
0 237 7 1 2 1493 140
0 238 5 1 1 237
0 239 7 2 2 1497 238
0 240 5 1 1 1576
0 241 7 1 2 236 1577
0 242 5 2 1 241
0 243 7 2 2 1283 1377
0 244 5 1 1 1580
0 245 7 2 2 1293 1368
0 246 5 1 1 1582
0 247 7 1 2 1581 1583
0 248 5 2 1 247
0 249 7 1 2 212 216
0 250 5 1 1 249
0 251 7 2 2 1561 250
0 252 5 1 1 1586
0 253 7 1 2 244 246
0 254 5 1 1 253
0 255 7 2 2 1584 254
0 256 5 1 1 1588
0 257 7 1 2 1587 1589
0 258 5 2 1 257
0 259 7 2 2 1585 1590
0 260 5 1 1 1592
0 261 7 1 2 1563 224
0 262 5 1 1 261
0 263 7 2 2 1567 262
0 264 5 1 1 1594
0 265 7 1 2 260 1595
0 266 5 2 1 265
0 267 7 2 2 1303 1351
0 268 5 1 1 1598
0 269 7 2 2 1275 1378
0 270 5 1 1 1600
0 271 7 1 2 1599 1601
0 272 5 2 1 271
0 273 7 2 2 1266 1387
0 274 5 1 1 1604
0 275 7 2 2 1294 1360
0 276 5 1 1 1606
0 277 7 1 2 1314 1342
0 278 5 1 1 277
0 279 7 1 2 1530 278
0 280 5 1 1 279
0 281 7 2 2 1535 280
0 282 5 1 1 1608
0 283 7 1 2 1607 1609
0 284 5 2 1 283
0 285 7 1 2 276 282
0 286 5 1 1 285
0 287 7 2 2 1610 286
0 288 5 1 1 1612
0 289 7 1 2 1605 1613
0 290 5 2 1 289
0 291 7 1 2 274 288
0 292 5 1 1 291
0 293 7 2 2 1614 292
0 294 5 1 1 1616
0 295 7 1 2 268 270
0 296 5 1 1 295
0 297 7 2 2 1602 296
0 298 5 1 1 1618
0 299 7 1 2 1617 1619
0 300 5 2 1 299
0 301 7 2 2 1603 1620
0 302 5 1 1 1622
0 303 7 1 2 252 256
0 304 5 1 1 303
0 305 7 2 2 1591 304
0 306 5 1 1 1624
0 307 7 1 2 302 1625
0 308 5 2 1 307
0 309 7 2 2 1323 1333
0 310 5 1 1 1628
0 311 7 2 2 1284 1369
0 312 5 1 1 1630
0 313 7 1 2 1629 1631
0 314 5 2 1 313
0 315 7 1 2 294 298
0 316 5 1 1 315
0 317 7 2 2 1621 316
0 318 5 1 1 1634
0 319 7 1 2 310 312
0 320 5 1 1 319
0 321 7 2 2 1632 320
0 322 5 1 1 1636
0 323 7 1 2 1635 1637
0 324 5 2 1 323
0 325 7 2 2 1633 1638
0 326 5 1 1 1640
0 327 7 1 2 1623 306
0 328 5 1 1 327
0 329 7 2 2 1626 328
0 330 5 1 1 1642
0 331 7 1 2 326 1643
0 332 5 2 1 331
0 333 7 2 2 1627 1644
0 334 5 1 1 1646
0 335 7 1 2 1593 264
0 336 5 1 1 335
0 337 7 2 2 1596 336
0 338 5 1 1 1648
0 339 7 1 2 334 1649
0 340 5 2 1 339
0 341 7 2 2 1597 1650
0 342 5 1 1 1652
0 343 7 1 2 1569 232
0 344 5 1 1 343
0 345 7 2 2 1573 344
0 346 5 1 1 1654
0 347 7 1 2 342 1655
0 348 5 2 1 347
0 349 7 2 2 1611 1615
0 350 5 1 1 1658
0 351 7 1 2 1641 330
0 352 5 1 1 351
0 353 7 2 2 1645 352
0 354 5 1 1 1660
0 355 7 1 2 350 1661
0 356 5 2 1 355
0 357 7 2 2 1304 1343
0 358 5 1 1 1664
0 359 7 2 2 1295 1352
0 360 5 1 1 1666
0 361 7 1 2 1665 1667
0 362 5 2 1 361
0 363 7 2 2 1267 1379
0 364 5 1 1 1670
0 365 7 1 2 358 360
0 366 5 1 1 365
0 367 7 2 2 1668 366
0 368 5 1 1 1672
0 369 7 1 2 1671 1673
0 370 5 2 1 369
0 371 7 2 2 1669 1674
0 372 5 1 1 1676
0 373 7 2 2 1276 1370
0 374 5 1 1 1678
0 375 7 2 2 32 1388
0 376 5 1 1 1680
0 377 7 1 2 1679 1681
0 378 5 2 1 377
0 379 7 2 2 1285 1361
0 380 5 1 1 1684
0 381 7 2 2 1296 1334
0 382 5 1 1 1686
0 383 7 2 2 1259 1353
0 384 5 1 1 1688
0 385 7 2 2 1277 1335
0 386 5 1 1 1690
0 387 7 2 2 1689 1691
0 388 5 2 1 1692
0 389 7 2 2 1286 1693
0 390 5 2 1 1696
0 391 7 2 2 1687 1697
0 392 5 2 1 1700
0 393 7 2 2 1305 1701
0 394 5 2 1 1704
0 395 7 1 2 1685 1705
0 396 5 2 1 395
0 397 7 1 2 380 1706
0 398 5 1 1 397
0 399 7 2 2 1708 398
0 400 5 1 1 1710
0 401 7 1 2 178 180
0 402 5 1 1 401
0 403 7 2 2 1531 402
0 404 5 1 1 1712
0 405 7 1 2 1711 1713
0 406 5 2 1 405
0 407 7 1 2 400 404
0 408 5 1 1 407
0 409 7 2 2 1714 408
0 410 5 1 1 1716
0 411 7 1 2 374 376
0 412 5 1 1 411
0 413 7 2 2 1682 412
0 414 5 1 1 1718
0 415 7 1 2 1717 1719
0 416 5 2 1 415
0 417 7 2 2 1683 1720
0 418 5 1 1 1722
0 419 7 1 2 372 418
0 420 5 2 1 419
0 421 7 2 2 1709 1715
0 422 5 1 1 1726
0 423 7 1 2 1677 1723
0 424 5 1 1 423
0 425 7 2 2 1724 424
0 426 5 1 1 1728
0 427 7 1 2 422 1729
0 428 5 2 1 427
0 429 7 2 2 1725 1730
0 430 5 1 1 1732
0 431 7 1 2 1659 354
0 432 5 1 1 431
0 433 7 2 2 1662 432
0 434 5 1 1 1734
0 435 7 1 2 430 1735
0 436 5 2 1 435
0 437 7 2 2 1663 1736
0 438 5 1 1 1738
0 439 7 1 2 1647 338
0 440 5 1 1 439
0 441 7 2 2 1651 440
0 442 5 1 1 1740
0 443 7 1 2 438 1741
0 444 5 2 1 443
0 445 7 1 2 318 322
0 446 5 1 1 445
0 447 7 2 2 1639 446
0 448 5 1 1 1744
0 449 7 1 2 1727 426
0 450 5 1 1 449
0 451 7 2 2 1731 450
0 452 5 1 1 1746
0 453 7 1 2 1745 1747
0 454 5 2 1 453
0 455 7 1 2 364 368
0 456 5 1 1 455
0 457 7 2 2 1675 456
0 458 5 1 1 1750
0 459 7 1 2 410 414
0 460 5 1 1 459
0 461 7 2 2 1721 460
0 462 5 1 1 1752
0 463 7 1 2 1751 1753
0 464 5 2 1 463
0 465 7 2 2 1287 1354
0 466 5 1 1 1756
0 467 7 2 2 1278 1362
0 468 5 1 1 1758
0 469 7 1 2 1757 1759
0 470 5 2 1 469
0 471 7 2 2 1268 1371
0 472 5 1 1 1762
0 473 7 1 2 466 468
0 474 5 1 1 473
0 475 7 2 2 1760 474
0 476 5 1 1 1764
0 477 7 1 2 1763 1765
0 478 5 2 1 477
0 479 7 2 2 1761 1766
0 480 5 1 1 1768
0 481 7 1 2 458 462
0 482 5 1 1 481
0 483 7 2 2 1754 482
0 484 5 1 1 1770
0 485 7 1 2 480 1771
0 486 5 2 1 485
0 487 7 2 2 1755 1772
0 488 5 1 1 1774
0 489 7 1 2 448 452
0 490 5 1 1 489
0 491 7 2 2 1748 490
0 492 5 1 1 1776
0 493 7 1 2 488 1777
0 494 5 2 1 493
0 495 7 2 2 1749 1778
0 496 5 1 1 1780
0 497 7 1 2 1733 434
0 498 5 1 1 497
0 499 7 2 2 1737 498
0 500 5 1 1 1782
0 501 7 1 2 496 1783
0 502 5 2 1 501
0 503 7 2 2 1260 1380
0 504 5 1 1 1786
0 505 7 1 2 472 476
0 506 5 1 1 505
0 507 7 2 2 1767 506
0 508 5 1 1 1788
0 509 7 1 2 1787 1789
0 510 5 2 1 509
0 511 7 2 2 1315 1325
0 512 5 1 1 1792
0 513 7 2 2 1297 1344
0 514 5 1 1 1794
0 515 7 1 2 1306 1336
0 516 5 1 1 515
0 517 7 1 2 1702 516
0 518 5 1 1 517
0 519 7 2 2 1707 518
0 520 5 1 1 1796
0 521 7 1 2 1795 1797
0 522 5 2 1 521
0 523 7 1 2 514 520
0 524 5 1 1 523
0 525 7 2 2 1798 524
0 526 5 1 1 1800
0 527 7 1 2 1793 1801
0 528 5 2 1 527
0 529 7 1 2 512 526
0 530 5 1 1 529
0 531 7 2 2 1802 530
0 532 5 1 1 1804
0 533 7 1 2 504 508
0 534 5 1 1 533
0 535 7 2 2 1790 534
0 536 5 1 1 1806
0 537 7 1 2 1805 1807
0 538 5 2 1 537
0 539 7 2 2 1791 1808
0 540 5 1 1 1810
0 541 7 1 2 1769 484
0 542 5 1 1 541
0 543 7 2 2 1773 542
0 544 5 1 1 1812
0 545 7 1 2 540 1813
0 546 5 2 1 545
0 547 7 2 2 1799 1803
0 548 5 1 1 1816
0 549 7 1 2 1811 544
0 550 5 1 1 549
0 551 7 2 2 1814 550
0 552 5 1 1 1818
0 553 7 1 2 548 1819
0 554 5 2 1 553
0 555 7 2 2 1815 1820
0 556 5 1 1 1822
0 557 7 1 2 1775 492
0 558 5 1 1 557
0 559 7 2 2 1779 558
0 560 5 1 1 1824
0 561 7 1 2 556 1825
0 562 5 2 1 561
0 563 7 2 2 1288 1345
0 564 5 1 1 1828
0 565 7 1 2 382 1698
0 566 5 1 1 565
0 567 7 2 2 1703 566
0 568 5 1 1 1830
0 569 7 1 2 1829 1831
0 570 5 2 1 569
0 571 7 2 2 1307 1326
0 572 5 1 1 1834
0 573 7 1 2 564 568
0 574 5 1 1 573
0 575 7 2 2 1832 574
0 576 5 1 1 1836
0 577 7 1 2 1835 1837
0 578 5 2 1 577
0 579 7 2 2 1833 1838
0 580 5 1 1 1840
0 581 7 1 2 532 536
0 582 5 1 1 581
0 583 7 2 2 1809 582
0 584 5 1 1 1842
0 585 7 1 2 580 1843
0 586 5 2 1 585
0 587 7 2 2 1279 1355
0 588 5 1 1 1846
0 589 7 2 2 1261 1372
0 590 5 1 1 1848
0 591 7 1 2 1847 1849
0 592 5 2 1 591
0 593 7 1 2 572 576
0 594 5 1 1 593
0 595 7 2 2 1839 594
0 596 5 1 1 1852
0 597 7 1 2 588 590
0 598 5 1 1 597
0 599 7 2 2 1850 598
0 600 5 1 1 1854
0 601 7 1 2 1853 1855
0 602 5 2 1 601
0 603 7 2 2 1851 1856
0 604 5 1 1 1858
0 605 7 1 2 1841 584
0 606 5 1 1 605
0 607 7 2 2 1844 606
0 608 5 1 1 1860
0 609 7 1 2 604 1861
0 610 5 2 1 609
0 611 7 2 2 1845 1862
0 612 5 1 1 1864
0 613 7 1 2 1817 552
0 614 5 1 1 613
0 615 7 2 2 1821 614
0 616 5 1 1 1866
0 617 7 1 2 612 1867
0 618 5 2 1 617
0 619 7 2 2 1269 1363
0 620 5 1 1 1870
0 621 7 1 2 596 600
0 622 5 1 1 621
0 623 7 2 2 1857 622
0 624 5 1 1 1872
0 625 7 1 2 1871 1873
0 626 5 2 1 625
0 627 7 2 2 1280 1346
0 628 5 1 1 1876
0 629 7 1 2 1289 1337
0 630 5 1 1 629
0 631 7 1 2 1694 630
0 632 5 1 1 631
0 633 7 2 2 1699 632
0 634 5 1 1 1878
0 635 7 1 2 1877 1879
0 636 5 2 1 635
0 637 7 2 2 1298 1327
0 638 5 1 1 1882
0 639 7 1 2 628 634
0 640 5 1 1 639
0 641 7 2 2 1880 640
0 642 5 1 1 1884
0 643 7 1 2 1883 1885
0 644 5 2 1 643
0 645 7 2 2 1881 1886
0 646 5 1 1 1888
0 647 7 1 2 620 624
0 648 5 1 1 647
0 649 7 2 2 1874 648
0 650 5 1 1 1890
0 651 7 1 2 646 1891
0 652 5 2 1 651
0 653 7 2 2 1875 1892
0 654 5 1 1 1894
0 655 7 1 2 1859 608
0 656 5 1 1 655
0 657 7 2 2 1863 656
0 658 5 1 1 1896
0 659 7 1 2 654 1897
0 660 5 2 1 659
0 661 7 2 2 1262 1364
0 662 5 1 1 1900
0 663 7 2 2 1270 1356
0 664 5 1 1 1902
0 665 7 1 2 1901 1903
0 666 5 2 1 665
0 667 7 1 2 638 642
0 668 5 1 1 667
0 669 7 2 2 1887 668
0 670 5 1 1 1906
0 671 7 1 2 662 664
0 672 5 1 1 671
0 673 7 2 2 1904 672
0 674 5 1 1 1908
0 675 7 1 2 1907 1909
0 676 5 2 1 675
0 677 7 2 2 1905 1910
0 678 5 1 1 1912
0 679 7 1 2 1889 650
0 680 5 1 1 679
0 681 7 2 2 1893 680
0 682 5 1 1 1914
0 683 7 1 2 678 1915
0 684 5 2 1 683
0 685 7 1 2 670 674
0 686 5 1 1 685
0 687 7 2 2 1911 686
0 688 5 1 1 1918
0 689 7 2 2 1271 1347
0 690 5 1 1 1920
0 691 7 2 2 1290 1328
0 692 5 1 1 1922
0 693 7 2 2 1921 1923
0 694 5 1 1 1924
0 695 7 2 2 1272 1338
0 696 5 1 1 1926
0 697 7 2 2 1263 1348
0 698 5 1 1 1928
0 699 7 2 2 1927 1929
0 700 5 2 1 1930
0 701 7 3 2 694 1932
0 702 5 1 1 1934
0 703 7 1 2 1919 702
0 704 5 2 1 703
0 705 7 1 2 384 386
0 706 5 1 1 705
0 707 7 2 2 1695 706
0 708 5 1 1 1939
0 709 7 1 2 690 692
0 710 5 1 1 709
0 711 7 1 2 1935 710
0 712 5 1 1 711
0 713 7 1 2 1925 1931
0 714 5 1 1 713
0 715 7 2 2 712 714
0 716 5 1 1 1941
0 717 7 1 2 1940 716
0 718 5 2 1 717
0 719 7 2 2 1281 1329
0 720 5 1 1 1945
0 721 7 1 2 696 698
0 722 5 1 1 721
0 723 7 2 2 1933 722
0 724 5 1 1 1947
0 725 7 1 2 1946 1948
0 726 5 2 1 725
0 727 7 1 2 720 724
0 728 5 1 1 727
0 729 7 2 2 1949 728
0 730 5 1 1 1951
0 731 7 2 2 1264 1339
0 732 5 1 1 1953
0 733 7 2 2 1273 1330
0 734 5 1 1 1955
0 735 7 2 2 1954 1956
0 736 5 2 1 1957
0 737 7 1 2 1952 1958
0 738 5 2 1 737
0 739 7 2 2 1950 1961
0 740 5 1 1 1963
0 741 7 1 2 708 1942
0 742 5 1 1 741
0 743 7 2 2 1943 742
0 744 5 1 1 1965
0 745 7 1 2 740 1966
0 746 5 2 1 745
0 747 7 2 2 1944 1967
0 748 5 1 1 1969
0 749 7 1 2 688 1936
0 750 5 1 1 749
0 751 7 2 2 1937 750
0 752 5 1 1 1971
0 753 7 1 2 748 1972
0 754 5 2 1 753
0 755 7 2 2 1938 1973
0 756 5 1 1 1975
0 757 7 1 2 1913 682
0 758 5 1 1 757
0 759 7 2 2 1916 758
0 760 5 1 1 1977
0 761 7 1 2 756 1978
0 762 5 2 1 761
0 763 7 2 2 1917 1979
0 764 5 1 1 1981
0 765 7 1 2 1895 658
0 766 5 1 1 765
0 767 7 2 2 1898 766
0 768 5 1 1 1983
0 769 7 1 2 764 1984
0 770 5 2 1 769
0 771 7 2 2 1899 1985
0 772 5 1 1 1987
0 773 7 1 2 1865 616
0 774 5 1 1 773
0 775 7 2 2 1868 774
0 776 5 1 1 1989
0 777 7 1 2 772 1990
0 778 5 2 1 777
0 779 7 2 2 1869 1991
0 780 5 1 1 1993
0 781 7 1 2 1823 560
0 782 5 1 1 781
0 783 7 2 2 1826 782
0 784 5 1 1 1995
0 785 7 1 2 780 1996
0 786 5 2 1 785
0 787 7 2 2 1827 1997
0 788 5 1 1 1999
0 789 7 1 2 1781 500
0 790 5 1 1 789
0 791 7 2 2 1784 790
0 792 5 1 1 2001
0 793 7 1 2 788 2002
0 794 5 2 1 793
0 795 7 2 2 1785 2003
0 796 5 1 1 2005
0 797 7 1 2 1739 442
0 798 5 1 1 797
0 799 7 2 2 1742 798
0 800 5 1 1 2007
0 801 7 1 2 796 2008
0 802 5 2 1 801
0 803 7 2 2 1743 2009
0 804 5 1 1 2011
0 805 7 1 2 1653 346
0 806 5 1 1 805
0 807 7 2 2 1656 806
0 808 5 1 1 2013
0 809 7 1 2 804 2014
0 810 5 2 1 809
0 811 7 2 2 1657 2015
0 812 5 1 1 2017
0 813 7 1 2 1575 240
0 814 5 1 1 813
0 815 7 2 2 1578 814
0 816 5 1 1 2019
0 817 7 1 2 812 2020
0 818 5 2 1 817
0 819 7 2 2 1579 2021
0 820 5 1 1 2023
0 821 7 1 2 1499 148
0 822 5 1 1 821
0 823 7 2 2 1502 822
0 824 5 1 1 2025
0 825 7 1 2 820 2026
0 826 5 2 1 825
0 827 7 2 2 1503 2027
0 828 5 1 1 2029
0 829 7 1 2 50 1447
0 830 5 1 1 829
0 831 7 2 2 1448 830
0 832 5 1 1 2031
0 833 7 1 2 828 2032
0 834 5 2 1 833
0 835 7 2 2 1449 2033
0 836 5 1 1 2035
0 837 7 2 2 1420 2036
0 838 5 2 1 2037
0 839 7 2 2 48 836
0 840 5 2 1 2041
0 841 7 1 2 2030 832
0 842 5 1 1 841
0 843 7 2 2 2034 842
0 844 5 1 1 2045
0 845 7 1 2 1418 844
0 846 5 3 1 845
0 847 7 1 2 2024 824
0 848 5 1 1 847
0 849 7 2 2 2028 848
0 850 5 1 1 2050
0 851 7 1 2 1416 850
0 852 5 3 1 851
0 853 7 1 2 46 2051
0 854 5 3 1 853
0 855 7 1 2 2018 816
0 856 5 1 1 855
0 857 7 2 2 2022 856
0 858 5 1 1 2058
0 859 7 1 2 1414 858
0 860 5 4 1 859
0 861 7 1 2 45 2059
0 862 5 3 1 861
0 863 7 1 2 2012 808
0 864 5 1 1 863
0 865 7 2 2 2016 864
0 866 5 1 1 2067
0 867 7 1 2 44 2068
0 868 5 3 1 867
0 869 7 1 2 1412 866
0 870 5 4 1 869
0 871 7 1 2 2006 800
0 872 5 1 1 871
0 873 7 2 2 2010 872
0 874 5 1 1 2076
0 875 7 1 2 1410 874
0 876 5 4 1 875
0 877 7 1 2 43 2077
0 878 5 3 1 877
0 879 7 1 2 2000 792
0 880 5 1 1 879
0 881 7 2 2 2004 880
0 882 5 1 1 2085
0 883 7 1 2 1408 882
0 884 5 4 1 883
0 885 7 1 2 42 2086
0 886 5 3 1 885
0 887 7 1 2 1994 784
0 888 5 1 1 887
0 889 7 2 2 1998 888
0 890 5 1 1 2094
0 891 7 1 2 1406 890
0 892 5 4 1 891
0 893 7 1 2 41 2095
0 894 5 3 1 893
0 895 7 1 2 1988 776
0 896 5 1 1 895
0 897 7 2 2 1992 896
0 898 5 1 1 2103
0 899 7 1 2 1404 898
0 900 5 3 1 899
0 901 7 1 2 40 2104
0 902 5 3 1 901
0 903 7 1 2 1982 768
0 904 5 1 1 903
0 905 7 2 2 1986 904
0 906 5 1 1 2111
0 907 7 1 2 1402 906
0 908 5 3 1 907
0 909 7 1 2 39 2112
0 910 5 3 1 909
0 911 7 1 2 1976 760
0 912 5 1 1 911
0 913 7 2 2 1980 912
0 914 5 1 1 2119
0 915 7 1 2 1400 914
0 916 5 5 1 915
0 917 7 1 2 38 2120
0 918 5 4 1 917
0 919 7 1 2 1970 752
0 920 5 1 1 919
0 921 7 2 2 1974 920
0 922 5 1 1 2130
0 923 7 2 2 37 2131
0 924 5 3 1 2132
0 925 7 2 2 1398 922
0 926 5 4 1 2137
0 927 7 1 2 1964 744
0 928 5 1 1 927
0 929 7 2 2 1968 928
0 930 5 1 1 2143
0 931 7 1 2 1396 930
0 932 5 3 1 931
0 933 7 1 2 36 2144
0 934 5 3 1 933
0 935 7 1 2 730 1959
0 936 5 1 1 935
0 937 7 2 2 1962 936
0 938 5 1 1 2151
0 939 7 1 2 1394 938
0 940 5 4 1 939
0 941 7 1 2 35 2152
0 942 5 3 1 941
0 943 7 1 2 732 734
0 944 5 1 1 943
0 945 7 2 2 1960 944
0 946 5 1 1 2160
0 947 7 1 2 34 2161
0 948 5 2 1 947
0 949 7 1 2 1392 946
0 950 5 2 1 949
0 951 7 2 2 1265 1331
0 952 5 1 1 2166
0 953 7 1 2 1390 952
0 954 5 1 1 953
0 955 7 1 2 2164 954
0 956 5 2 1 955
0 957 7 1 2 2162 2168
0 958 7 1 2 2157 957
0 959 5 1 1 958
0 960 7 1 2 2153 959
0 961 5 2 1 960
0 962 7 1 2 2148 2170
0 963 5 1 1 962
0 964 7 3 2 2145 963
0 965 5 1 1 2172
0 966 7 1 2 2139 2173
0 967 5 1 1 966
0 968 7 1 2 2134 967
0 969 7 1 2 2126 968
0 970 5 1 1 969
0 971 7 2 2 2121 970
0 972 5 1 1 2175
0 973 7 1 2 2116 972
0 974 5 1 1 973
0 975 7 2 2 2113 974
0 976 5 2 1 2177
0 977 7 1 2 2108 2179
0 978 5 1 1 977
0 979 7 2 2 2105 978
0 980 5 2 1 2181
0 981 7 1 2 2100 2183
0 982 5 1 1 981
0 983 7 2 2 2096 982
0 984 5 1 1 2185
0 985 7 1 2 2091 984
0 986 5 2 1 985
0 987 7 1 2 2087 2187
0 988 5 1 1 987
0 989 7 1 2 2082 988
0 990 5 2 1 989
0 991 7 1 2 2078 2189
0 992 7 1 2 2072 991
0 993 5 1 1 992
0 994 7 1 2 2069 993
0 995 7 1 2 2064 994
0 996 5 1 1 995
0 997 7 1 2 2060 996
0 998 5 2 1 997
0 999 7 1 2 2055 2191
0 1000 5 1 1 999
0 1001 7 2 2 2052 1000
0 1002 5 2 1 2193
0 1003 7 1 2 47 2046
0 1004 5 3 1 1003
0 1005 7 1 2 2195 2197
0 1006 5 1 1 1005
0 1007 7 2 2 2047 1006
0 1008 5 1 1 2200
0 1009 7 1 2 2043 1008
0 1010 5 1 1 1009
0 1011 7 2 2 2039 1010
0 1012 5 1 1 2202
0 1013 7 3 2 2048 2198
0 1014 5 2 1 2204
0 1015 7 1 2 2196 2207
0 1016 5 1 1 1015
0 1017 7 1 2 2194 2205
0 1018 5 1 1 1017
0 1019 7 1 2 1016 1018
0 1020 5 1 1 1019
0 1021 7 1 2 2042 2201
0 1022 5 1 1 1021
0 1023 7 3 2 2053 2056
0 1024 5 2 1 2209
0 1025 7 1 2 2061 2212
0 1026 5 1 1 1025
0 1027 7 1 2 2192 2210
0 1028 5 1 1 1027
0 1029 7 2 2 2062 2065
0 1030 5 2 1 2214
0 1031 7 1 2 2073 2216
0 1032 5 1 1 1031
0 1033 7 3 2 2070 2074
0 1034 5 1 1 2218
0 1035 7 1 2 2190 2219
0 1036 5 1 1 1035
0 1037 7 1 2 2079 1036
0 1038 5 1 1 1037
0 1039 7 3 2 2080 2083
0 1040 5 1 1 2221
0 1041 7 1 2 2188 2222
0 1042 5 1 1 1041
0 1043 7 1 2 2088 1042
0 1044 5 1 1 1043
0 1045 7 2 2 2089 2092
0 1046 5 2 1 2224
0 1047 7 1 2 2186 2226
0 1048 5 1 1 1047
0 1049 7 2 2 2097 2101
0 1050 5 2 1 2228
0 1051 7 1 2 2182 2230
0 1052 5 1 1 1051
0 1053 7 1 2 2184 2229
0 1054 5 1 1 1053
0 1055 7 1 2 1052 1054
0 1056 5 1 1 1055
0 1057 7 1 2 2133 2174
0 1058 5 1 1 1057
0 1059 7 4 2 2114 2117
0 1060 5 2 1 2232
0 1061 7 1 2 2122 2233
0 1062 5 1 1 1061
0 1063 7 1 2 1058 1062
0 1064 5 1 1 1063
0 1065 7 1 2 2127 2236
0 1066 5 1 1 1065
0 1067 7 1 2 2176 2234
0 1068 5 1 1 1067
0 1069 7 1 2 2138 965
0 1070 5 1 1 1069
0 1071 7 3 2 2146 2149
0 1072 5 2 1 2238
0 1073 7 1 2 2154 2241
0 1074 5 1 1 1073
0 1075 7 1 2 2171 2239
0 1076 5 1 1 1075
0 1077 7 1 2 2155 2158
0 1078 5 2 1 1077
0 1079 7 1 2 33 2167
0 1080 5 1 1 1079
0 1081 7 1 2 2163 1080
0 1082 5 1 1 1081
0 1083 7 2 2 2165 1082
0 1084 5 2 1 2245
0 1085 7 1 2 2243 2246
0 1086 5 2 1 1085
0 1087 7 1 2 1076 2249
0 1088 7 1 2 1074 1087
0 1089 5 1 1 1088
0 1090 7 1 2 1070 1089
0 1091 7 1 2 1068 1090
0 1092 7 1 2 1066 1091
0 1093 7 1 2 1064 1092
0 1094 7 3 2 2106 2109
0 1095 5 2 1 2251
0 1096 7 1 2 2178 2252
0 1097 5 1 1 1096
0 1098 7 1 2 2180 2254
0 1099 5 1 1 1098
0 1100 7 1 2 1097 1099
0 1101 7 1 2 1093 1100
0 1102 7 1 2 1056 1101
0 1103 5 1 1 1102
0 1104 7 1 2 1048 1103
0 1105 7 1 2 1044 1104
0 1106 7 1 2 1038 1105
0 1107 7 1 2 1032 1106
0 1108 7 1 2 1028 1107
0 1109 7 1 2 1026 1108
0 1110 7 1 2 1022 1109
0 1111 7 1 2 1020 1110
0 1112 7 1 2 2203 1111
0 1113 5 1 1 1112
0 1114 7 1 2 2159 2247
0 1115 5 1 1 1114
0 1116 7 2 2 2156 1115
0 1117 5 2 1 2256
0 1118 7 1 2 2150 2258
0 1119 5 1 1 1118
0 1120 7 2 2 2147 1119
0 1121 5 1 1 2260
0 1122 7 1 2 2135 1121
0 1123 5 2 1 1122
0 1124 7 1 2 2140 2262
0 1125 5 1 1 1124
0 1126 7 1 2 2128 1125
0 1127 5 1 1 1126
0 1128 7 1 2 2123 1127
0 1129 5 2 1 1128
0 1130 7 1 2 2118 2264
0 1131 5 1 1 1130
0 1132 7 2 2 2115 1131
0 1133 5 2 1 2266
0 1134 7 1 2 2110 2268
0 1135 5 1 1 1134
0 1136 7 2 2 2107 1135
0 1137 5 1 1 2270
0 1138 7 2 2 2102 1137
0 1139 5 1 1 2272
0 1140 7 2 2 2098 1139
0 1141 5 2 1 2274
0 1142 7 1 2 2093 2276
0 1143 5 1 1 1142
0 1144 7 2 2 2090 1143
0 1145 5 2 1 2278
0 1146 7 1 2 2084 2280
0 1147 5 1 1 1146
0 1148 7 2 2 2081 1147
0 1149 5 2 1 2282
0 1150 7 1 2 2071 2284
0 1151 5 1 1 1150
0 1152 7 2 2 2075 1151
0 1153 5 2 1 2286
0 1154 7 1 2 2066 2288
0 1155 5 1 1 1154
0 1156 7 2 2 2063 1155
0 1157 5 2 1 2290
0 1158 7 1 2 2057 2292
0 1159 5 1 1 1158
0 1160 7 2 2 2054 1159
0 1161 5 2 1 2294
0 1162 7 1 2 2199 2296
0 1163 5 1 1 1162
0 1164 7 2 2 2049 1163
0 1165 5 1 1 2298
0 1166 7 1 2 2040 1165
0 1167 5 1 1 1166
0 1168 7 1 2 2038 2299
0 1169 5 1 1 1168
0 1170 7 1 2 1167 1169
0 1171 5 1 1 1170
0 1172 7 1 2 2206 2297
0 1173 5 1 1 1172
0 1174 7 1 2 2208 2295
0 1175 5 1 1 1174
0 1176 7 1 2 1173 1175
0 1177 5 1 1 1176
0 1178 7 1 2 2215 2287
0 1179 5 1 1 1178
0 1180 7 1 2 2217 2289
0 1181 5 1 1 1180
0 1182 7 1 2 2220 2285
0 1183 5 1 1 1182
0 1184 7 1 2 1034 2283
0 1185 5 1 1 1184
0 1186 7 1 2 1183 1185
0 1187 5 1 1 1186
0 1188 7 1 2 1040 2281
0 1189 5 1 1 1188
0 1190 7 1 2 2223 2279
0 1191 5 1 1 1190
0 1192 7 1 2 2225 2277
0 1193 5 1 1 1192
0 1194 7 1 2 2227 2275
0 1195 5 1 1 1194
0 1196 7 1 2 1193 1195
0 1197 5 1 1 1196
0 1198 7 1 2 2099 2273
0 1199 5 1 1 1198
0 1200 7 1 2 2231 2271
0 1201 5 1 1 1200
0 1202 7 1 2 2255 2267
0 1203 5 1 1 1202
0 1204 7 1 2 2253 2269
0 1205 5 1 1 1204
0 1206 7 1 2 2124 2237
0 1207 5 1 1 1206
0 1208 7 1 2 2235 2265
0 1209 5 1 1 1208
0 1210 7 1 2 2125 2263
0 1211 7 1 2 2129 1210
0 1212 5 1 1 1211
0 1213 7 1 2 2141 1212
0 1214 5 1 1 1213
0 1215 7 1 2 2136 2142
0 1216 5 1 1 1215
0 1217 7 1 2 2261 1216
0 1218 5 1 1 1217
0 1219 7 1 2 2240 2257
0 1220 5 1 1 1219
0 1221 7 1 2 2169 2244
0 1222 5 1 1 1221
0 1223 7 1 2 2248 1222
0 1224 5 1 1 1223
0 1225 7 1 2 2250 1224
0 1226 5 1 1 1225
0 1227 7 1 2 2242 2259
0 1228 5 1 1 1227
0 1229 7 1 2 1226 1228
0 1230 7 1 2 1220 1229
0 1231 5 1 1 1230
0 1232 7 1 2 1218 1231
0 1233 7 1 2 1214 1232
0 1234 7 1 2 1209 1233
0 1235 7 1 2 1207 1234
0 1236 7 1 2 1205 1235
0 1237 7 1 2 1203 1236
0 1238 7 1 2 1201 1237
0 1239 7 1 2 1199 1238
0 1240 5 1 1 1239
0 1241 7 1 2 1197 1240
0 1242 7 1 2 1191 1241
0 1243 7 1 2 1189 1242
0 1244 7 1 2 1187 1243
0 1245 7 1 2 1181 1244
0 1246 7 1 2 1179 1245
0 1247 7 1 2 2044 1246
0 1248 7 1 2 2213 2293
0 1249 5 1 1 1248
0 1250 7 1 2 2211 2291
0 1251 5 1 1 1250
0 1252 7 1 2 1249 1251
0 1253 7 1 2 1247 1252
0 1254 7 1 2 1177 1253
0 1255 7 1 2 1012 1254
0 1256 7 1 2 1171 1255
0 1257 5 1 1 1256
0 1258 7 1 2 1113 1257
3 4299 5 0 1 1258
