1 0 0 8 0
2 16 1 0
2 17 1 0
2 18 1 0
2 19 1 0
2 20 1 0
2 21 1 0
2 22 1 0
2 23 1 0
1 1 0 8 0
2 24 1 1
2 25 1 1
2 26 1 1
2 27 1 1
2 28 1 1
2 29 1 1
2 30 1 1
2 31 1 1
1 2 0 8 0
2 32 1 2
2 41 1 2
2 64 1 2
2 103 1 2
2 156 1 2
2 227 1 2
2 314 1 2
2 417 1 2
1 3 0 9 0
2 520 1 3
2 615 1 3
2 696 1 3
2 761 1 3
2 810 1 3
2 843 1 3
2 860 1 3
2 862 1 3
2 863 1 3
1 4 0 8 0
2 864 1 4
2 865 1 4
2 866 1 4
2 867 1 4
2 868 1 4
2 869 1 4
2 870 1 4
2 871 1 4
1 5 0 9 0
2 872 1 5
2 873 1 5
2 874 1 5
2 875 1 5
2 876 1 5
2 877 1 5
2 878 1 5
2 879 1 5
2 880 1 5
1 6 0 8 0
2 881 1 6
2 882 1 6
2 883 1 6
2 884 1 6
2 885 1 6
2 886 1 6
2 887 1 6
2 888 1 6
1 7 0 8 0
2 889 1 7
2 890 1 7
2 891 1 7
2 892 1 7
2 893 1 7
2 894 1 7
2 895 1 7
2 896 1 7
1 8 0 8 0
2 897 1 8
2 898 1 8
2 899 1 8
2 900 1 8
2 901 1 8
2 902 1 8
2 903 1 8
2 904 1 8
1 9 0 8 0
2 905 1 9
2 906 1 9
2 907 1 9
2 908 1 9
2 909 1 9
2 910 1 9
2 911 1 9
2 912 1 9
1 10 0 9 0
2 913 1 10
2 914 1 10
2 915 1 10
2 916 1 10
2 917 1 10
2 918 1 10
2 919 1 10
2 920 1 10
2 921 1 10
1 11 0 8 0
2 922 1 11
2 923 1 11
2 924 1 11
2 925 1 11
2 926 1 11
2 927 1 11
2 928 1 11
2 929 1 11
1 12 0 8 0
2 930 1 12
2 931 1 12
2 932 1 12
2 933 1 12
2 934 1 12
2 935 1 12
2 936 1 12
2 937 1 12
1 13 0 8 0
2 938 1 13
2 939 1 13
2 940 1 13
2 941 1 13
2 942 1 13
2 943 1 13
2 944 1 13
2 945 1 13
1 14 0 8 0
2 946 1 14
2 947 1 14
2 948 1 14
2 949 1 14
2 950 1 14
2 951 1 14
2 952 1 14
2 953 1 14
1 15 0 8 0
2 954 1 15
2 955 1 15
2 956 1 15
2 957 1 15
2 958 1 15
2 959 1 15
2 960 1 15
2 961 1 15
2 962 1 33
2 963 1 33
2 964 1 35
2 965 1 35
2 966 1 39
2 967 1 39
2 968 1 40
2 969 1 40
2 970 1 42
2 971 1 42
2 972 1 44
2 973 1 44
2 974 1 46
2 975 1 46
2 976 1 50
2 977 1 50
2 978 1 51
2 979 1 51
2 980 1 52
2 981 1 52
2 982 1 55
2 983 1 55
2 984 1 58
2 985 1 58
2 986 1 61
2 987 1 61
2 988 1 65
2 989 1 65
2 990 1 67
2 991 1 67
2 992 1 69
2 993 1 69
2 994 1 73
2 995 1 73
2 996 1 74
2 997 1 74
2 998 1 75
2 999 1 75
2 1000 1 77
2 1001 1 77
2 1002 1 79
2 1003 1 79
2 1004 1 81
2 1005 1 81
2 1006 1 83
2 1007 1 83
2 1008 1 84
2 1009 1 84
2 1010 1 91
2 1011 1 91
2 1012 1 94
2 1013 1 94
2 1014 1 97
2 1015 1 97
2 1016 1 100
2 1017 1 100
2 1018 1 104
2 1019 1 104
2 1020 1 106
2 1021 1 106
2 1022 1 108
2 1023 1 108
2 1024 1 114
2 1025 1 114
2 1026 1 115
2 1027 1 115
2 1028 1 116
2 1029 1 116
2 1030 1 119
2 1031 1 119
2 1032 1 122
2 1033 1 122
2 1034 1 125
2 1035 1 125
2 1036 1 128
2 1037 1 128
2 1038 1 130
2 1039 1 130
2 1040 1 132
2 1041 1 132
2 1042 1 137
2 1043 1 137
2 1044 1 138
2 1045 1 138
2 1046 1 141
2 1047 1 141
2 1048 1 144
2 1049 1 144
2 1050 1 147
2 1051 1 147
2 1052 1 150
2 1053 1 150
2 1054 1 153
2 1055 1 153
2 1056 1 157
2 1057 1 157
2 1058 1 159
2 1059 1 159
2 1060 1 161
2 1061 1 161
2 1062 1 163
2 1063 1 163
2 1064 1 165
2 1065 1 165
2 1066 1 167
2 1067 1 167
2 1068 1 169
2 1069 1 169
2 1070 1 171
2 1071 1 171
2 1072 1 172
2 1073 1 172
2 1074 1 175
2 1075 1 175
2 1076 1 178
2 1077 1 178
2 1078 1 181
2 1079 1 181
2 1080 1 184
2 1081 1 184
2 1082 1 187
2 1083 1 187
2 1084 1 189
2 1085 1 189
2 1086 1 191
2 1087 1 191
2 1088 1 196
2 1089 1 196
2 1090 1 197
2 1091 1 197
2 1092 1 200
2 1093 1 200
2 1094 1 203
2 1095 1 203
2 1096 1 206
2 1097 1 206
2 1098 1 209
2 1099 1 209
2 1100 1 212
2 1101 1 212
2 1102 1 215
2 1103 1 215
2 1104 1 218
2 1105 1 218
2 1106 1 221
2 1107 1 221
2 1108 1 224
2 1109 1 224
2 1110 1 228
2 1111 1 228
2 1112 1 230
2 1113 1 230
2 1114 1 232
2 1115 1 232
2 1116 1 234
2 1117 1 234
2 1118 1 236
2 1119 1 236
2 1120 1 238
2 1121 1 238
2 1122 1 244
2 1123 1 244
2 1124 1 245
2 1125 1 245
2 1126 1 246
2 1127 1 246
2 1128 1 249
2 1129 1 249
2 1130 1 252
2 1131 1 252
2 1132 1 255
2 1133 1 255
2 1134 1 258
2 1135 1 258
2 1136 1 260
2 1137 1 260
2 1138 1 262
2 1139 1 262
2 1140 1 264
2 1141 1 264
2 1142 1 266
2 1143 1 266
2 1144 1 271
2 1145 1 271
2 1146 1 272
2 1147 1 272
2 1148 1 275
2 1149 1 275
2 1150 1 278
2 1151 1 278
2 1152 1 281
2 1153 1 281
2 1154 1 284
2 1155 1 284
2 1156 1 287
2 1157 1 287
2 1158 1 290
2 1159 1 290
2 1160 1 293
2 1161 1 293
2 1162 1 296
2 1163 1 296
2 1164 1 299
2 1165 1 299
2 1166 1 302
2 1167 1 302
2 1168 1 305
2 1169 1 305
2 1170 1 308
2 1171 1 308
2 1172 1 311
2 1173 1 311
2 1174 1 315
2 1175 1 315
2 1176 1 317
2 1177 1 317
2 1178 1 319
2 1179 1 319
2 1180 1 321
2 1181 1 321
2 1182 1 323
2 1183 1 323
2 1184 1 325
2 1185 1 325
2 1186 1 327
2 1187 1 327
2 1188 1 329
2 1189 1 329
2 1190 1 334
2 1191 1 334
2 1192 1 335
2 1193 1 335
2 1194 1 338
2 1195 1 338
2 1196 1 341
2 1197 1 341
2 1198 1 343
2 1199 1 343
2 1200 1 346
2 1201 1 346
2 1202 1 349
2 1203 1 349
2 1204 1 351
2 1205 1 351
2 1206 1 353
2 1207 1 353
2 1208 1 357
2 1209 1 357
2 1210 1 358
2 1211 1 358
2 1212 1 359
2 1213 1 359
2 1214 1 362
2 1215 1 362
2 1216 1 365
2 1217 1 365
2 1218 1 367
2 1219 1 367
2 1220 1 369
2 1221 1 369
2 1222 1 374
2 1223 1 374
2 1224 1 375
2 1225 1 375
2 1226 1 378
2 1227 1 378
2 1228 1 381
2 1229 1 381
2 1230 1 384
2 1231 1 384
2 1232 1 387
2 1233 1 387
2 1234 1 390
2 1235 1 390
2 1236 1 393
2 1237 1 393
2 1238 1 396
2 1239 1 396
2 1240 1 399
2 1241 1 399
2 1242 1 402
2 1243 1 402
2 1244 1 405
2 1245 1 405
2 1246 1 408
2 1247 1 408
2 1248 1 411
2 1249 1 411
2 1250 1 414
2 1251 1 414
2 1252 1 418
2 1253 1 418
2 1254 1 420
2 1255 1 420
2 1256 1 422
2 1257 1 422
2 1258 1 424
2 1259 1 424
2 1260 1 426
2 1261 1 426
2 1262 1 432
2 1263 1 432
2 1264 1 433
2 1265 1 433
2 1266 1 434
2 1267 1 434
2 1268 1 437
2 1269 1 437
2 1270 1 440
2 1271 1 440
2 1272 1 443
2 1273 1 443
2 1274 1 446
2 1275 1 446
2 1276 1 448
2 1277 1 448
2 1278 1 450
2 1279 1 450
2 1280 1 455
2 1281 1 455
2 1282 1 456
2 1283 1 456
2 1284 1 459
2 1285 1 459
2 1286 1 462
2 1287 1 462
2 1288 1 464
2 1289 1 464
2 1290 1 466
2 1291 1 466
2 1292 1 471
2 1293 1 471
2 1294 1 472
2 1295 1 472
2 1296 1 475
2 1297 1 475
2 1298 1 478
2 1299 1 478
2 1300 1 480
2 1301 1 480
2 1302 1 482
2 1303 1 482
2 1304 1 484
2 1305 1 484
2 1306 1 487
2 1307 1 487
2 1308 1 490
2 1309 1 490
2 1310 1 493
2 1311 1 493
2 1312 1 496
2 1313 1 496
2 1314 1 499
2 1315 1 499
2 1316 1 502
2 1317 1 502
2 1318 1 505
2 1319 1 505
2 1320 1 508
2 1321 1 508
2 1322 1 511
2 1323 1 511
2 1324 1 514
2 1325 1 514
2 1326 1 517
2 1327 1 517
2 1328 1 521
2 1329 1 521
2 1330 1 523
2 1331 1 523
2 1332 1 525
2 1333 1 525
2 1334 1 527
2 1335 1 527
2 1336 1 529
2 1337 1 529
2 1338 1 531
2 1339 1 531
2 1340 1 533
2 1341 1 533
2 1342 1 535
2 1343 1 535
2 1344 1 537
2 1345 1 537
2 1346 1 539
2 1347 1 539
2 1348 1 542
2 1349 1 542
2 1350 1 545
2 1351 1 545
2 1352 1 548
2 1353 1 548
2 1354 1 551
2 1355 1 551
2 1356 1 554
2 1357 1 554
2 1358 1 557
2 1359 1 557
2 1360 1 560
2 1361 1 560
2 1362 1 563
2 1363 1 563
2 1364 1 565
2 1365 1 565
2 1366 1 567
2 1367 1 567
2 1368 1 572
2 1369 1 572
2 1370 1 573
2 1371 1 573
2 1372 1 576
2 1373 1 576
2 1374 1 579
2 1375 1 579
2 1376 1 582
2 1377 1 582
2 1378 1 585
2 1379 1 585
2 1380 1 588
2 1381 1 588
2 1382 1 591
2 1383 1 591
2 1384 1 594
2 1385 1 594
2 1386 1 597
2 1387 1 597
2 1388 1 600
2 1389 1 600
2 1390 1 603
2 1391 1 603
2 1392 1 606
2 1393 1 606
2 1394 1 609
2 1395 1 609
2 1396 1 612
2 1397 1 612
2 1398 1 616
2 1399 1 616
2 1400 1 618
2 1401 1 618
2 1402 1 620
2 1403 1 620
2 1404 1 622
2 1405 1 622
2 1406 1 624
2 1407 1 624
2 1408 1 626
2 1409 1 626
2 1410 1 628
2 1411 1 628
2 1412 1 630
2 1413 1 630
2 1414 1 632
2 1415 1 632
2 1416 1 634
2 1417 1 634
2 1418 1 636
2 1419 1 636
2 1420 1 641
2 1421 1 641
2 1422 1 642
2 1423 1 642
2 1424 1 645
2 1425 1 645
2 1426 1 648
2 1427 1 648
2 1428 1 651
2 1429 1 651
2 1430 1 654
2 1431 1 654
2 1432 1 657
2 1433 1 657
2 1434 1 660
2 1435 1 660
2 1436 1 663
2 1437 1 663
2 1438 1 666
2 1439 1 666
2 1440 1 669
2 1441 1 669
2 1442 1 672
2 1443 1 672
2 1444 1 675
2 1445 1 675
2 1446 1 678
2 1447 1 678
2 1448 1 681
2 1449 1 681
2 1450 1 684
2 1451 1 684
2 1452 1 687
2 1453 1 687
2 1454 1 690
2 1455 1 690
2 1456 1 693
2 1457 1 693
2 1458 1 697
2 1459 1 697
2 1460 1 699
2 1461 1 699
2 1462 1 701
2 1463 1 701
2 1464 1 703
2 1465 1 703
2 1466 1 705
2 1467 1 705
2 1468 1 707
2 1469 1 707
2 1470 1 709
2 1471 1 709
2 1472 1 711
2 1473 1 711
2 1474 1 713
2 1475 1 713
2 1476 1 718
2 1477 1 718
2 1478 1 719
2 1479 1 719
2 1480 1 722
2 1481 1 722
2 1482 1 725
2 1483 1 725
2 1484 1 728
2 1485 1 728
2 1486 1 731
2 1487 1 731
2 1488 1 734
2 1489 1 734
2 1490 1 737
2 1491 1 737
2 1492 1 740
2 1493 1 740
2 1494 1 743
2 1495 1 743
2 1496 1 746
2 1497 1 746
2 1498 1 749
2 1499 1 749
2 1500 1 752
2 1501 1 752
2 1502 1 755
2 1503 1 755
2 1504 1 758
2 1505 1 758
2 1506 1 762
2 1507 1 762
2 1508 1 764
2 1509 1 764
2 1510 1 766
2 1511 1 766
2 1512 1 768
2 1513 1 768
2 1514 1 770
2 1515 1 770
2 1516 1 771
2 1517 1 771
2 1518 1 772
2 1519 1 772
2 1520 1 774
2 1521 1 774
2 1522 1 779
2 1523 1 779
2 1524 1 780
2 1525 1 780
2 1526 1 783
2 1527 1 783
2 1528 1 786
2 1529 1 786
2 1530 1 789
2 1531 1 789
2 1532 1 792
2 1533 1 792
2 1534 1 795
2 1535 1 795
2 1536 1 798
2 1537 1 798
2 1538 1 801
2 1539 1 801
2 1540 1 804
2 1541 1 804
2 1542 1 807
2 1543 1 807
2 1544 1 811
2 1545 1 811
2 1546 1 813
2 1547 1 813
2 1548 1 815
2 1549 1 815
2 1550 1 817
2 1551 1 817
2 1552 1 819
2 1553 1 819
2 1554 1 825
2 1555 1 825
2 1556 1 828
2 1557 1 828
2 1558 1 828
2 1559 1 831
2 1560 1 831
2 1561 1 834
2 1562 1 834
2 1563 1 837
2 1564 1 837
2 1565 1 840
2 1566 1 840
2 1567 1 844
2 1568 1 844
2 1569 1 846
2 1570 1 846
2 1571 1 853
2 1572 1 853
2 1573 1 854
2 1574 1 854
2 1575 1 857
2 1576 1 857
3 1784 7 0 2 16 897
0 33 7 2 2 17 905
0 34 5 1 1 962
0 35 7 2 2 24 898
0 36 5 1 1 964
0 37 7 1 2 34 36
0 38 5 1 1 37
0 39 7 2 2 963 965
0 40 5 2 1 966
3 1785 7 0 2 38 968
0 42 7 2 2 32 899
0 43 5 1 1 970
0 44 7 2 2 25 906
0 45 5 1 1 972
0 46 7 2 2 18 913
0 47 5 1 1 974
0 48 7 1 2 45 47
0 49 5 1 1 48
0 50 7 2 2 973 975
0 51 5 2 1 976
0 52 7 2 2 49 978
0 53 5 1 1 980
0 54 7 1 2 971 981
0 55 5 2 1 54
0 56 7 1 2 43 53
0 57 5 1 1 56
0 58 7 2 2 982 57
0 59 5 1 1 984
0 60 7 1 2 967 985
0 61 5 2 1 60
0 62 7 1 2 969 59
0 63 5 1 1 62
3 1786 7 0 2 986 63
0 65 7 2 2 983 987
0 66 5 1 1 988
0 67 7 2 2 19 922
0 68 5 1 1 990
0 69 7 2 2 41 907
0 70 5 1 1 992
0 71 7 1 2 68 70
0 72 5 1 1 71
0 73 7 2 2 991 993
0 74 5 2 1 994
0 75 7 2 2 72 996
0 76 5 1 1 998
0 77 7 2 2 26 914
0 78 5 1 1 1000
0 79 7 2 2 520 900
0 80 5 1 1 1002
0 81 7 2 2 1001 1003
0 82 5 1 1 1004
0 83 7 2 2 979 82
0 84 5 2 1 1006
0 85 7 1 2 977 1005
0 86 5 1 1 85
0 87 7 1 2 1008 86
0 88 5 1 1 87
0 89 7 1 2 78 80
0 90 5 1 1 89
0 91 7 2 2 88 90
0 92 5 1 1 1010
0 93 7 1 2 999 1011
0 94 5 2 1 93
0 95 7 1 2 76 92
0 96 5 1 1 95
0 97 7 2 2 1012 96
0 98 5 1 1 1014
0 99 7 1 2 66 1015
0 100 5 2 1 99
0 101 7 1 2 989 98
0 102 5 1 1 101
3 1787 7 0 2 1016 102
0 104 7 2 2 1013 1017
0 105 5 1 1 1018
0 106 7 2 2 864 901
0 107 5 1 1 1020
0 108 7 2 2 64 915
0 109 5 1 1 1022
0 110 7 1 2 615 908
0 111 5 1 1 110
0 112 7 1 2 997 111
0 113 5 1 1 112
0 114 7 2 2 696 995
0 115 5 2 1 1024
0 116 7 2 2 113 1026
0 117 5 1 1 1028
0 118 7 1 2 1023 1029
0 119 5 2 1 118
0 120 7 1 2 109 117
0 121 5 1 1 120
0 122 7 2 2 1030 121
0 123 5 1 1 1032
0 124 7 1 2 1021 1033
0 125 5 2 1 124
0 126 7 1 2 107 123
0 127 5 1 1 126
0 128 7 2 2 1034 127
0 129 5 1 1 1036
0 130 7 2 2 20 930
0 131 5 1 1 1038
0 132 7 2 2 27 923
0 133 5 1 1 1040
0 134 7 1 2 131 133
0 135 5 1 1 134
0 136 7 1 2 1039 1041
0 137 5 2 1 136
0 138 7 2 2 135 1042
0 139 5 1 1 1044
0 140 7 1 2 1037 1045
0 141 5 2 1 140
0 142 7 1 2 129 139
0 143 5 1 1 142
0 144 7 2 2 1046 143
0 145 5 1 1 1048
0 146 7 1 2 1009 1049
0 147 5 2 1 146
0 148 7 1 2 1007 145
0 149 5 1 1 148
0 150 7 2 2 1050 149
0 151 5 1 1 1052
0 152 7 1 2 105 1053
0 153 5 2 1 152
0 154 7 1 2 1019 151
0 155 5 1 1 154
3 1788 7 0 2 1054 155
0 157 7 2 2 1051 1055
0 158 5 1 1 1056
0 159 7 2 2 1043 1047
0 160 5 1 1 1058
0 161 7 2 2 1031 1035
0 162 5 1 1 1060
0 163 7 2 2 28 931
0 164 5 1 1 1062
0 165 7 2 2 872 902
0 166 5 1 1 1064
0 167 7 2 2 761 916
0 168 5 1 1 1066
0 169 7 2 2 865 909
0 170 5 1 1 1068
0 171 7 2 2 1025 1069
0 172 5 2 1 1070
0 173 7 1 2 1027 170
0 174 5 1 1 173
0 175 7 2 2 1072 174
0 176 5 1 1 1074
0 177 7 1 2 1067 1075
0 178 5 2 1 177
0 179 7 1 2 168 176
0 180 5 1 1 179
0 181 7 2 2 1076 180
0 182 5 1 1 1078
0 183 7 1 2 1065 1079
0 184 5 2 1 183
0 185 7 1 2 166 182
0 186 5 1 1 185
0 187 7 2 2 1080 186
0 188 5 1 1 1082
0 189 7 2 2 103 924
0 190 5 1 1 1084
0 191 7 2 2 21 938
0 192 5 1 1 1086
0 193 7 1 2 190 192
0 194 5 1 1 193
0 195 7 1 2 1085 1087
0 196 5 2 1 195
0 197 7 2 2 194 1088
0 198 5 1 1 1090
0 199 7 1 2 1083 1091
0 200 5 2 1 199
0 201 7 1 2 188 198
0 202 5 1 1 201
0 203 7 2 2 1092 202
0 204 5 1 1 1094
0 205 7 1 2 1063 1095
0 206 5 2 1 205
0 207 7 1 2 164 204
0 208 5 1 1 207
0 209 7 2 2 1096 208
0 210 5 1 1 1098
0 211 7 1 2 162 1099
0 212 5 2 1 211
0 213 7 1 2 1061 210
0 214 5 1 1 213
0 215 7 2 2 1100 214
0 216 5 1 1 1102
0 217 7 1 2 160 1103
0 218 5 2 1 217
0 219 7 1 2 1059 216
0 220 5 1 1 219
0 221 7 2 2 1104 220
0 222 5 1 1 1106
0 223 7 1 2 158 1107
0 224 5 2 1 223
0 225 7 1 2 1057 222
0 226 5 1 1 225
3 1789 7 0 2 1108 226
0 228 7 2 2 1105 1109
0 229 5 1 1 1110
0 230 7 2 2 1097 1101
0 231 5 1 1 1112
0 232 7 2 2 1089 1093
0 233 5 1 1 1114
0 234 7 2 2 1077 1081
0 235 5 1 1 1116
0 236 7 2 2 881 903
0 237 5 1 1 1118
0 238 7 2 2 866 917
0 239 5 1 1 1120
0 240 7 1 2 873 910
0 241 5 1 1 240
0 242 7 1 2 1073 241
0 243 5 1 1 242
0 244 7 2 2 874 1071
0 245 5 2 1 1122
0 246 7 2 2 243 1124
0 247 5 1 1 1126
0 248 7 1 2 1121 1127
0 249 5 2 1 248
0 250 7 1 2 239 247
0 251 5 1 1 250
0 252 7 2 2 1128 251
0 253 5 1 1 1130
0 254 7 1 2 1119 1131
0 255 5 2 1 254
0 256 7 1 2 237 253
0 257 5 1 1 256
0 258 7 2 2 1132 257
0 259 5 1 1 1134
0 260 7 2 2 22 946
0 261 5 1 1 1136
0 262 7 2 2 29 939
0 263 5 1 1 1138
0 264 7 2 2 156 932
0 265 5 1 1 1140
0 266 7 2 2 810 925
0 267 5 1 1 1142
0 268 7 1 2 265 267
0 269 5 1 1 268
0 270 7 1 2 1141 1143
0 271 5 2 1 270
0 272 7 2 2 269 1144
0 273 5 1 1 1146
0 274 7 1 2 1139 1147
0 275 5 2 1 274
0 276 7 1 2 263 273
0 277 5 1 1 276
0 278 7 2 2 1148 277
0 279 5 1 1 1150
0 280 7 1 2 1137 1151
0 281 5 2 1 280
0 282 7 1 2 261 279
0 283 5 1 1 282
0 284 7 2 2 1152 283
0 285 5 1 1 1154
0 286 7 1 2 1135 1155
0 287 5 2 1 286
0 288 7 1 2 259 285
0 289 5 1 1 288
0 290 7 2 2 1156 289
0 291 5 1 1 1158
0 292 7 1 2 235 1159
0 293 5 2 1 292
0 294 7 1 2 1117 291
0 295 5 1 1 294
0 296 7 2 2 1160 295
0 297 5 1 1 1162
0 298 7 1 2 233 1163
0 299 5 2 1 298
0 300 7 1 2 1115 297
0 301 5 1 1 300
0 302 7 2 2 1164 301
0 303 5 1 1 1166
0 304 7 1 2 231 1167
0 305 5 2 1 304
0 306 7 1 2 1113 303
0 307 5 1 1 306
0 308 7 2 2 1168 307
0 309 5 1 1 1170
0 310 7 1 2 229 1171
0 311 5 2 1 310
0 312 7 1 2 1111 309
0 313 5 1 1 312
3 1790 7 0 2 1172 313
0 315 7 2 2 1169 1173
0 316 5 1 1 1174
0 317 7 2 2 1161 1165
0 318 5 1 1 1176
0 319 7 2 2 1129 1133
0 320 5 1 1 1178
0 321 7 2 2 1153 1157
0 322 5 1 1 1180
0 323 7 2 2 1145 1149
0 324 5 1 1 1182
0 325 7 2 2 30 947
0 326 5 1 1 1184
0 327 7 2 2 875 918
0 328 5 1 1 1186
0 329 7 2 2 867 926
0 330 5 1 1 1188
0 331 7 1 2 328 330
0 332 5 1 1 331
0 333 7 1 2 1187 1189
0 334 5 2 1 333
0 335 7 2 2 332 1190
0 336 5 1 1 1192
0 337 7 1 2 1185 1193
0 338 5 2 1 337
0 339 7 1 2 326 336
0 340 5 1 1 339
0 341 7 2 2 1194 340
0 342 5 1 1 1196
0 343 7 2 2 843 933
0 344 5 1 1 1198
0 345 7 1 2 1123 1199
0 346 5 2 1 345
0 347 7 1 2 1125 344
0 348 5 1 1 347
0 349 7 2 2 1200 348
0 350 5 1 1 1202
0 351 7 2 2 889 904
0 352 5 1 1 1204
0 353 7 2 2 882 911
0 354 5 1 1 1206
0 355 7 1 2 352 354
0 356 5 1 1 355
0 357 7 2 2 1205 1207
0 358 5 2 1 1208
0 359 7 2 2 356 1210
0 360 5 1 1 1212
0 361 7 1 2 1203 1213
0 362 5 2 1 361
0 363 7 1 2 350 360
0 364 5 1 1 363
0 365 7 2 2 1214 364
0 366 5 1 1 1216
0 367 7 2 2 227 940
0 368 5 1 1 1218
0 369 7 2 2 23 954
0 370 5 1 1 1220
0 371 7 1 2 368 370
0 372 5 1 1 371
0 373 7 1 2 1219 1221
0 374 5 2 1 373
0 375 7 2 2 372 1222
0 376 5 1 1 1224
0 377 7 1 2 1217 1225
0 378 5 2 1 377
0 379 7 1 2 366 376
0 380 5 1 1 379
0 381 7 2 2 1226 380
0 382 5 1 1 1228
0 383 7 1 2 1197 1229
0 384 5 2 1 383
0 385 7 1 2 342 382
0 386 5 1 1 385
0 387 7 2 2 1230 386
0 388 5 1 1 1232
0 389 7 1 2 324 1233
0 390 5 2 1 389
0 391 7 1 2 1183 388
0 392 5 1 1 391
0 393 7 2 2 1234 392
0 394 5 1 1 1236
0 395 7 1 2 322 1237
0 396 5 2 1 395
0 397 7 1 2 1181 394
0 398 5 1 1 397
0 399 7 2 2 1238 398
0 400 5 1 1 1240
0 401 7 1 2 320 1241
0 402 5 2 1 401
0 403 7 1 2 1179 400
0 404 5 1 1 403
0 405 7 2 2 1242 404
0 406 5 1 1 1244
0 407 7 1 2 318 1245
0 408 5 2 1 407
0 409 7 1 2 1177 406
0 410 5 1 1 409
0 411 7 2 2 1246 410
0 412 5 1 1 1248
0 413 7 1 2 316 1249
0 414 5 2 1 413
0 415 7 1 2 1175 412
0 416 5 1 1 415
3 1791 7 0 2 1250 416
0 418 7 2 2 1247 1251
0 419 5 1 1 1252
0 420 7 2 2 1239 1243
0 421 5 1 1 1254
0 422 7 2 2 1231 1235
0 423 5 1 1 1256
0 424 7 2 2 31 955
0 425 5 1 1 1258
0 426 7 2 2 868 934
0 427 5 1 1 1260
0 428 7 1 2 883 919
0 429 5 1 1 428
0 430 7 1 2 1211 429
0 431 5 1 1 430
0 432 7 2 2 920 1209
0 433 5 2 1 1262
0 434 7 2 2 431 1264
0 435 5 1 1 1266
0 436 7 1 2 1261 1267
0 437 5 2 1 436
0 438 7 1 2 427 435
0 439 5 1 1 438
0 440 7 2 2 1268 439
0 441 5 1 1 1270
0 442 7 1 2 1259 1271
0 443 5 2 1 442
0 444 7 1 2 425 441
0 445 5 1 1 444
0 446 7 2 2 1272 445
0 447 5 1 1 1274
0 448 7 2 2 876 927
0 449 5 1 1 1276
0 450 7 2 2 314 948
0 451 5 1 1 1278
0 452 7 1 2 449 451
0 453 5 1 1 452
0 454 7 1 2 1277 1279
0 455 5 2 1 454
0 456 7 2 2 453 1280
0 457 5 1 1 1282
0 458 7 1 2 1275 1283
0 459 5 2 1 458
0 460 7 1 2 447 457
0 461 5 1 1 460
0 462 7 2 2 1284 461
0 463 5 1 1 1286
0 464 7 2 2 890 912
0 465 5 1 1 1288
0 466 7 2 2 860 941
0 467 5 1 1 1290
0 468 7 1 2 465 467
0 469 5 1 1 468
0 470 7 1 2 1289 1291
0 471 5 2 1 470
0 472 7 2 2 469 1292
0 473 5 1 1 1294
0 474 7 1 2 1287 1295
0 475 5 2 1 474
0 476 7 1 2 463 473
0 477 5 1 1 476
0 478 7 2 2 1296 477
0 479 5 1 1 1298
0 480 7 2 2 1201 1215
0 481 5 1 1 1300
0 482 7 2 2 1191 1195
0 483 5 1 1 1302
0 484 7 2 2 1223 1227
0 485 5 1 1 1304
0 486 7 1 2 483 485
0 487 5 2 1 486
0 488 7 1 2 1303 1305
0 489 5 1 1 488
0 490 7 2 2 1306 489
0 491 5 1 1 1308
0 492 7 1 2 481 1309
0 493 5 2 1 492
0 494 7 1 2 1301 491
0 495 5 1 1 494
0 496 7 2 2 1310 495
0 497 5 1 1 1312
0 498 7 1 2 1299 1313
0 499 5 2 1 498
0 500 7 1 2 479 497
0 501 5 1 1 500
0 502 7 2 2 1314 501
0 503 5 1 1 1316
0 504 7 1 2 423 1317
0 505 5 2 1 504
0 506 7 1 2 1257 503
0 507 5 1 1 506
0 508 7 2 2 1318 507
0 509 5 1 1 1320
0 510 7 1 2 421 1321
0 511 5 2 1 510
0 512 7 1 2 1255 509
0 513 5 1 1 512
0 514 7 2 2 1322 513
0 515 5 1 1 1324
0 516 7 1 2 419 1325
0 517 5 2 1 516
0 518 7 1 2 1253 515
0 519 5 1 1 518
3 1792 7 0 2 1326 519
0 521 7 2 2 1323 1327
0 522 5 1 1 1328
0 523 7 2 2 1315 1319
0 524 5 1 1 1330
0 525 7 2 2 1307 1311
0 526 5 1 1 1332
0 527 7 2 2 1269 1273
0 528 5 1 1 1334
0 529 7 2 2 1293 1297
0 530 5 1 1 1336
0 531 7 2 2 1281 1285
0 532 5 1 1 1338
0 533 7 2 2 884 928
0 534 5 1 1 1340
0 535 7 2 2 877 935
0 536 5 1 1 1342
0 537 7 2 2 891 921
0 538 5 1 1 1344
0 539 7 2 2 417 956
0 540 5 1 1 1346
0 541 7 1 2 1263 1347
0 542 5 2 1 541
0 543 7 1 2 1265 540
0 544 5 1 1 543
0 545 7 2 2 1348 544
0 546 5 1 1 1350
0 547 7 1 2 1345 1351
0 548 5 2 1 547
0 549 7 1 2 538 546
0 550 5 1 1 549
0 551 7 2 2 1352 550
0 552 5 1 1 1354
0 553 7 1 2 1343 1355
0 554 5 2 1 553
0 555 7 1 2 536 552
0 556 5 1 1 555
0 557 7 2 2 1356 556
0 558 5 1 1 1358
0 559 7 1 2 1341 1359
0 560 5 2 1 559
0 561 7 1 2 534 558
0 562 5 1 1 561
0 563 7 2 2 1360 562
0 564 5 1 1 1362
0 565 7 2 2 862 949
0 566 5 1 1 1364
0 567 7 2 2 869 942
0 568 5 1 1 1366
0 569 7 1 2 566 568
0 570 5 1 1 569
0 571 7 1 2 1365 1367
0 572 5 2 1 571
0 573 7 2 2 570 1368
0 574 5 1 1 1370
0 575 7 1 2 1363 1371
0 576 5 2 1 575
0 577 7 1 2 564 574
0 578 5 1 1 577
0 579 7 2 2 1372 578
0 580 5 1 1 1374
0 581 7 1 2 532 1375
0 582 5 2 1 581
0 583 7 1 2 1339 580
0 584 5 1 1 583
0 585 7 2 2 1376 584
0 586 5 1 1 1378
0 587 7 1 2 530 1379
0 588 5 2 1 587
0 589 7 1 2 1337 586
0 590 5 1 1 589
0 591 7 2 2 1380 590
0 592 5 1 1 1382
0 593 7 1 2 528 1383
0 594 5 2 1 593
0 595 7 1 2 1335 592
0 596 5 1 1 595
0 597 7 2 2 1384 596
0 598 5 1 1 1386
0 599 7 1 2 526 1387
0 600 5 2 1 599
0 601 7 1 2 1333 598
0 602 5 1 1 601
0 603 7 2 2 1388 602
0 604 5 1 1 1390
0 605 7 1 2 524 1391
0 606 5 2 1 605
0 607 7 1 2 1331 604
0 608 5 1 1 607
0 609 7 2 2 1392 608
0 610 5 1 1 1394
0 611 7 1 2 522 1395
0 612 5 2 1 611
0 613 7 1 2 1329 610
0 614 5 1 1 613
3 1793 7 0 2 1396 614
0 616 7 2 2 1393 1397
0 617 5 1 1 1398
0 618 7 2 2 1385 1389
0 619 5 1 1 1400
0 620 7 2 2 1377 1381
0 621 5 1 1 1402
0 622 7 2 2 1369 1373
0 623 5 1 1 1404
0 624 7 2 2 1357 1361
0 625 5 1 1 1406
0 626 7 2 2 1349 1353
0 627 5 1 1 1408
0 628 7 2 2 878 943
0 629 5 1 1 1410
0 630 7 2 2 870 950
0 631 5 1 1 1412
0 632 7 2 2 885 936
0 633 5 1 1 1414
0 634 7 2 2 863 957
0 635 5 1 1 1416
0 636 7 2 2 892 929
0 637 5 1 1 1418
0 638 7 1 2 635 637
0 639 5 1 1 638
0 640 7 1 2 1417 1419
0 641 5 2 1 640
0 642 7 2 2 639 1420
0 643 5 1 1 1422
0 644 7 1 2 1415 1423
0 645 5 2 1 644
0 646 7 1 2 633 643
0 647 5 1 1 646
0 648 7 2 2 1424 647
0 649 5 1 1 1426
0 650 7 1 2 1413 1427
0 651 5 2 1 650
0 652 7 1 2 631 649
0 653 5 1 1 652
0 654 7 2 2 1428 653
0 655 5 1 1 1430
0 656 7 1 2 1411 1431
0 657 5 2 1 656
0 658 7 1 2 629 655
0 659 5 1 1 658
0 660 7 2 2 1432 659
0 661 5 1 1 1434
0 662 7 1 2 627 1435
0 663 5 2 1 662
0 664 7 1 2 1409 661
0 665 5 1 1 664
0 666 7 2 2 1436 665
0 667 5 1 1 1438
0 668 7 1 2 625 1439
0 669 5 2 1 668
0 670 7 1 2 1407 667
0 671 5 1 1 670
0 672 7 2 2 1440 671
0 673 5 1 1 1442
0 674 7 1 2 623 1443
0 675 5 2 1 674
0 676 7 1 2 1405 673
0 677 5 1 1 676
0 678 7 2 2 1444 677
0 679 5 1 1 1446
0 680 7 1 2 621 1447
0 681 5 2 1 680
0 682 7 1 2 1403 679
0 683 5 1 1 682
0 684 7 2 2 1448 683
0 685 5 1 1 1450
0 686 7 1 2 619 1451
0 687 5 2 1 686
0 688 7 1 2 1401 685
0 689 5 1 1 688
0 690 7 2 2 1452 689
0 691 5 1 1 1454
0 692 7 1 2 617 1455
0 693 5 2 1 692
0 694 7 1 2 1399 691
0 695 5 1 1 694
3 1794 7 0 2 1456 695
0 697 7 2 2 1453 1457
0 698 5 1 1 1458
0 699 7 2 2 1445 1449
0 700 5 1 1 1460
0 701 7 2 2 1437 1441
0 702 5 1 1 1462
0 703 7 2 2 1429 1433
0 704 5 1 1 1464
0 705 7 2 2 1421 1425
0 706 5 1 1 1466
0 707 7 2 2 879 951
0 708 5 1 1 1468
0 709 7 2 2 886 944
0 710 5 1 1 1470
0 711 7 2 2 871 958
0 712 5 1 1 1472
0 713 7 2 2 893 937
0 714 5 1 1 1474
0 715 7 1 2 712 714
0 716 5 1 1 715
0 717 7 1 2 1473 1475
0 718 5 2 1 717
0 719 7 2 2 716 1476
0 720 5 1 1 1478
0 721 7 1 2 1471 1479
0 722 5 2 1 721
0 723 7 1 2 710 720
0 724 5 1 1 723
0 725 7 2 2 1480 724
0 726 5 1 1 1482
0 727 7 1 2 1469 1483
0 728 5 2 1 727
0 729 7 1 2 708 726
0 730 5 1 1 729
0 731 7 2 2 1484 730
0 732 5 1 1 1486
0 733 7 1 2 706 1487
0 734 5 2 1 733
0 735 7 1 2 1467 732
0 736 5 1 1 735
0 737 7 2 2 1488 736
0 738 5 1 1 1490
0 739 7 1 2 704 1491
0 740 5 2 1 739
0 741 7 1 2 1465 738
0 742 5 1 1 741
0 743 7 2 2 1492 742
0 744 5 1 1 1494
0 745 7 1 2 702 1495
0 746 5 2 1 745
0 747 7 1 2 1463 744
0 748 5 1 1 747
0 749 7 2 2 1496 748
0 750 5 1 1 1498
0 751 7 1 2 700 1499
0 752 5 2 1 751
0 753 7 1 2 1461 750
0 754 5 1 1 753
0 755 7 2 2 1500 754
0 756 5 1 1 1502
0 757 7 1 2 698 1503
0 758 5 2 1 757
0 759 7 1 2 1459 756
0 760 5 1 1 759
3 1795 7 0 2 1504 760
0 762 7 2 2 1501 1505
0 763 5 1 1 1506
0 764 7 2 2 1493 1497
0 765 5 1 1 1508
0 766 7 2 2 1485 1489
0 767 5 1 1 1510
0 768 7 2 2 1477 1481
0 769 5 1 1 1512
0 770 7 2 2 887 952
0 771 5 2 1 1514
0 772 7 2 2 894 945
0 773 5 1 1 1518
0 774 7 2 2 880 959
0 775 5 1 1 1520
0 776 7 1 2 773 775
0 777 5 1 1 776
0 778 7 1 2 1519 1521
0 779 5 2 1 778
0 780 7 2 2 777 1522
0 781 5 1 1 1524
0 782 7 1 2 1515 1525
0 783 5 2 1 782
0 784 7 1 2 1516 781
0 785 5 1 1 784
0 786 7 2 2 1526 785
0 787 5 1 1 1528
0 788 7 1 2 769 1529
0 789 5 2 1 788
0 790 7 1 2 1513 787
0 791 5 1 1 790
0 792 7 2 2 1530 791
0 793 5 1 1 1532
0 794 7 1 2 767 1533
0 795 5 2 1 794
0 796 7 1 2 1511 793
0 797 5 1 1 796
0 798 7 2 2 1534 797
0 799 5 1 1 1536
0 800 7 1 2 765 1537
0 801 5 2 1 800
0 802 7 1 2 1509 799
0 803 5 1 1 802
0 804 7 2 2 1538 803
0 805 5 1 1 1540
0 806 7 1 2 763 1541
0 807 5 2 1 806
0 808 7 1 2 1507 805
0 809 5 1 1 808
3 1796 7 0 2 1542 809
0 811 7 2 2 1539 1543
0 812 5 1 1 1544
0 813 7 2 2 1531 1535
0 814 5 1 1 1546
0 815 7 2 2 1523 1527
0 816 5 1 1 1548
0 817 7 2 2 888 960
0 818 5 1 1 1550
0 819 7 2 2 895 953
0 820 5 1 1 1552
0 821 7 1 2 818 1553
0 822 5 1 1 821
0 823 7 1 2 1551 820
0 824 5 1 1 823
0 825 7 2 2 822 824
0 826 5 1 1 1554
0 827 7 1 2 816 826
0 828 5 3 1 827
0 829 7 1 2 1549 1555
0 830 5 1 1 829
0 831 7 2 2 1556 830
0 832 5 1 1 1559
0 833 7 1 2 814 1560
0 834 5 2 1 833
0 835 7 1 2 1547 832
0 836 5 1 1 835
0 837 7 2 2 1561 836
0 838 5 1 1 1563
0 839 7 1 2 812 1564
0 840 5 2 1 839
0 841 7 1 2 1545 838
0 842 5 1 1 841
3 1797 7 0 2 1565 842
0 844 7 2 2 1562 1566
0 845 5 1 1 1567
0 846 7 2 2 896 961
0 847 5 1 1 1569
0 848 7 1 2 1557 847
0 849 5 1 1 848
0 850 7 1 2 1517 1558
0 851 5 1 1 850
0 852 7 1 2 1570 851
0 853 5 2 1 852
0 854 7 2 2 849 1571
0 855 5 1 1 1573
0 856 7 1 2 845 1574
0 857 5 2 1 856
0 858 7 1 2 1568 855
0 859 5 1 1 858
3 1798 7 0 2 1575 859
0 861 7 1 2 1572 1576
3 1799 5 0 1 861
