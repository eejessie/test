1 0 0 92 0
2 25 1 0
2 26 1 0
2 61251 1 0
2 61252 1 0
2 61253 1 0
2 61254 1 0
2 61255 1 0
2 61256 1 0
2 61257 1 0
2 61258 1 0
2 61259 1 0
2 61260 1 0
2 61261 1 0
2 61262 1 0
2 61263 1 0
2 61264 1 0
2 61265 1 0
2 61266 1 0
2 61267 1 0
2 61268 1 0
2 61269 1 0
2 61270 1 0
2 61271 1 0
2 61272 1 0
2 61273 1 0
2 61274 1 0
2 61275 1 0
2 61276 1 0
2 61277 1 0
2 61278 1 0
2 61279 1 0
2 61280 1 0
2 61281 1 0
2 61282 1 0
2 61283 1 0
2 61284 1 0
2 61285 1 0
2 61286 1 0
2 61287 1 0
2 61288 1 0
2 61289 1 0
2 61290 1 0
2 61291 1 0
2 61292 1 0
2 61293 1 0
2 61294 1 0
2 61295 1 0
2 61296 1 0
2 61297 1 0
2 61298 1 0
2 61299 1 0
2 61300 1 0
2 61301 1 0
2 61302 1 0
2 61303 1 0
2 61304 1 0
2 61305 1 0
2 61306 1 0
2 61307 1 0
2 61308 1 0
2 61309 1 0
2 61310 1 0
2 61311 1 0
2 61312 1 0
2 61313 1 0
2 61314 1 0
2 61315 1 0
2 61316 1 0
2 61317 1 0
2 61318 1 0
2 61319 1 0
2 61320 1 0
2 61321 1 0
2 61322 1 0
2 61323 1 0
2 61324 1 0
2 61325 1 0
2 61326 1 0
2 61327 1 0
2 61328 1 0
2 61329 1 0
2 61330 1 0
2 61331 1 0
2 61332 1 0
2 61333 1 0
2 61334 1 0
2 61335 1 0
2 61336 1 0
2 61337 1 0
2 61338 1 0
2 61339 1 0
2 61340 1 0
1 1 0 83 0
2 61341 1 1
2 61342 1 1
2 61343 1 1
2 61344 1 1
2 61345 1 1
2 61346 1 1
2 61347 1 1
2 61348 1 1
2 61349 1 1
2 61350 1 1
2 61351 1 1
2 61352 1 1
2 61353 1 1
2 61354 1 1
2 61355 1 1
2 61356 1 1
2 61357 1 1
2 61358 1 1
2 61359 1 1
2 61360 1 1
2 61361 1 1
2 61362 1 1
2 61363 1 1
2 61364 1 1
2 61365 1 1
2 61366 1 1
2 61367 1 1
2 61368 1 1
2 61369 1 1
2 61370 1 1
2 61371 1 1
2 61372 1 1
2 61373 1 1
2 61374 1 1
2 61375 1 1
2 61376 1 1
2 61377 1 1
2 61378 1 1
2 61379 1 1
2 61380 1 1
2 61381 1 1
2 61382 1 1
2 61383 1 1
2 61384 1 1
2 61385 1 1
2 61386 1 1
2 61387 1 1
2 61388 1 1
2 61389 1 1
2 61390 1 1
2 61391 1 1
2 61392 1 1
2 61393 1 1
2 61394 1 1
2 61395 1 1
2 61396 1 1
2 61397 1 1
2 61398 1 1
2 61399 1 1
2 61400 1 1
2 61401 1 1
2 61402 1 1
2 61403 1 1
2 61404 1 1
2 61405 1 1
2 61406 1 1
2 61407 1 1
2 61408 1 1
2 61409 1 1
2 61410 1 1
2 61411 1 1
2 61412 1 1
2 61413 1 1
2 61414 1 1
2 61415 1 1
2 61416 1 1
2 61417 1 1
2 61418 1 1
2 61419 1 1
2 61420 1 1
2 61421 1 1
2 61422 1 1
2 61423 1 1
1 2 0 272 0
2 61424 1 2
2 61425 1 2
2 61426 1 2
2 61427 1 2
2 61428 1 2
2 61429 1 2
2 61430 1 2
2 61431 1 2
2 61432 1 2
2 61433 1 2
2 61434 1 2
2 61435 1 2
2 61436 1 2
2 61437 1 2
2 61438 1 2
2 61439 1 2
2 61440 1 2
2 61441 1 2
2 61442 1 2
2 61443 1 2
2 61444 1 2
2 61445 1 2
2 61446 1 2
2 61447 1 2
2 61448 1 2
2 61449 1 2
2 61450 1 2
2 61451 1 2
2 61452 1 2
2 61453 1 2
2 61454 1 2
2 61455 1 2
2 61456 1 2
2 61457 1 2
2 61458 1 2
2 61459 1 2
2 61460 1 2
2 61461 1 2
2 61462 1 2
2 61463 1 2
2 61464 1 2
2 61465 1 2
2 61466 1 2
2 61467 1 2
2 61468 1 2
2 61469 1 2
2 61470 1 2
2 61471 1 2
2 61472 1 2
2 61473 1 2
2 61474 1 2
2 61475 1 2
2 61476 1 2
2 61477 1 2
2 61478 1 2
2 61479 1 2
2 61480 1 2
2 61481 1 2
2 61482 1 2
2 61483 1 2
2 61484 1 2
2 61485 1 2
2 61486 1 2
2 61487 1 2
2 61488 1 2
2 61489 1 2
2 61490 1 2
2 61491 1 2
2 61492 1 2
2 61493 1 2
2 61494 1 2
2 61495 1 2
2 61496 1 2
2 61497 1 2
2 61498 1 2
2 61499 1 2
2 61500 1 2
2 61501 1 2
2 61502 1 2
2 61503 1 2
2 61504 1 2
2 61505 1 2
2 61506 1 2
2 61507 1 2
2 61508 1 2
2 61509 1 2
2 61510 1 2
2 61511 1 2
2 61512 1 2
2 61513 1 2
2 61514 1 2
2 61515 1 2
2 61516 1 2
2 61517 1 2
2 61518 1 2
2 61519 1 2
2 61520 1 2
2 61521 1 2
2 61522 1 2
2 61523 1 2
2 61524 1 2
2 61525 1 2
2 61526 1 2
2 61527 1 2
2 61528 1 2
2 61529 1 2
2 61530 1 2
2 61531 1 2
2 61532 1 2
2 61533 1 2
2 61534 1 2
2 61535 1 2
2 61536 1 2
2 61537 1 2
2 61538 1 2
2 61539 1 2
2 61540 1 2
2 61541 1 2
2 61542 1 2
2 61543 1 2
2 61544 1 2
2 61545 1 2
2 61546 1 2
2 61547 1 2
2 61548 1 2
2 61549 1 2
2 61550 1 2
2 61551 1 2
2 61552 1 2
2 61553 1 2
2 61554 1 2
2 61555 1 2
2 61556 1 2
2 61557 1 2
2 61558 1 2
2 61559 1 2
2 61560 1 2
2 61561 1 2
2 61562 1 2
2 61563 1 2
2 61564 1 2
2 61565 1 2
2 61566 1 2
2 61567 1 2
2 61568 1 2
2 61569 1 2
2 61570 1 2
2 61571 1 2
2 61572 1 2
2 61573 1 2
2 61574 1 2
2 61575 1 2
2 61576 1 2
2 61577 1 2
2 61578 1 2
2 61579 1 2
2 61580 1 2
2 61581 1 2
2 61582 1 2
2 61583 1 2
2 61584 1 2
2 61585 1 2
2 61586 1 2
2 61587 1 2
2 61588 1 2
2 61589 1 2
2 61590 1 2
2 61591 1 2
2 61592 1 2
2 61593 1 2
2 61594 1 2
2 61595 1 2
2 61596 1 2
2 61597 1 2
2 61598 1 2
2 61599 1 2
2 61600 1 2
2 61601 1 2
2 61602 1 2
2 61603 1 2
2 61604 1 2
2 61605 1 2
2 61606 1 2
2 61607 1 2
2 61608 1 2
2 61609 1 2
2 61610 1 2
2 61611 1 2
2 61612 1 2
2 61613 1 2
2 61614 1 2
2 61615 1 2
2 61616 1 2
2 61617 1 2
2 61618 1 2
2 61619 1 2
2 61620 1 2
2 61621 1 2
2 61622 1 2
2 61623 1 2
2 61624 1 2
2 61625 1 2
2 61626 1 2
2 61627 1 2
2 61628 1 2
2 61629 1 2
2 61630 1 2
2 61631 1 2
2 61632 1 2
2 61633 1 2
2 61634 1 2
2 61635 1 2
2 61636 1 2
2 61637 1 2
2 61638 1 2
2 61639 1 2
2 61640 1 2
2 61641 1 2
2 61642 1 2
2 61643 1 2
2 61644 1 2
2 61645 1 2
2 61646 1 2
2 61647 1 2
2 61648 1 2
2 61649 1 2
2 61650 1 2
2 61651 1 2
2 61652 1 2
2 61653 1 2
2 61654 1 2
2 61655 1 2
2 61656 1 2
2 61657 1 2
2 61658 1 2
2 61659 1 2
2 61660 1 2
2 61661 1 2
2 61662 1 2
2 61663 1 2
2 61664 1 2
2 61665 1 2
2 61666 1 2
2 61667 1 2
2 61668 1 2
2 61669 1 2
2 61670 1 2
2 61671 1 2
2 61672 1 2
2 61673 1 2
2 61674 1 2
2 61675 1 2
2 61676 1 2
2 61677 1 2
2 61678 1 2
2 61679 1 2
2 61680 1 2
2 61681 1 2
2 61682 1 2
2 61683 1 2
2 61684 1 2
2 61685 1 2
2 61686 1 2
2 61687 1 2
2 61688 1 2
2 61689 1 2
2 61690 1 2
2 61691 1 2
2 61692 1 2
2 61693 1 2
2 61694 1 2
2 61695 1 2
1 3 0 244 0
2 61696 1 3
2 61697 1 3
2 61698 1 3
2 61699 1 3
2 61700 1 3
2 61701 1 3
2 61702 1 3
2 61703 1 3
2 61704 1 3
2 61705 1 3
2 61706 1 3
2 61707 1 3
2 61708 1 3
2 61709 1 3
2 61710 1 3
2 61711 1 3
2 61712 1 3
2 61713 1 3
2 61714 1 3
2 61715 1 3
2 61716 1 3
2 61717 1 3
2 61718 1 3
2 61719 1 3
2 61720 1 3
2 61721 1 3
2 61722 1 3
2 61723 1 3
2 61724 1 3
2 61725 1 3
2 61726 1 3
2 61727 1 3
2 61728 1 3
2 61729 1 3
2 61730 1 3
2 61731 1 3
2 61732 1 3
2 61733 1 3
2 61734 1 3
2 61735 1 3
2 61736 1 3
2 61737 1 3
2 61738 1 3
2 61739 1 3
2 61740 1 3
2 61741 1 3
2 61742 1 3
2 61743 1 3
2 61744 1 3
2 61745 1 3
2 61746 1 3
2 61747 1 3
2 61748 1 3
2 61749 1 3
2 61750 1 3
2 61751 1 3
2 61752 1 3
2 61753 1 3
2 61754 1 3
2 61755 1 3
2 61756 1 3
2 61757 1 3
2 61758 1 3
2 61759 1 3
2 61760 1 3
2 61761 1 3
2 61762 1 3
2 61763 1 3
2 61764 1 3
2 61765 1 3
2 61766 1 3
2 61767 1 3
2 61768 1 3
2 61769 1 3
2 61770 1 3
2 61771 1 3
2 61772 1 3
2 61773 1 3
2 61774 1 3
2 61775 1 3
2 61776 1 3
2 61777 1 3
2 61778 1 3
2 61779 1 3
2 61780 1 3
2 61781 1 3
2 61782 1 3
2 61783 1 3
2 61784 1 3
2 61785 1 3
2 61786 1 3
2 61787 1 3
2 61788 1 3
2 61789 1 3
2 61790 1 3
2 61791 1 3
2 61792 1 3
2 61793 1 3
2 61794 1 3
2 61795 1 3
2 61796 1 3
2 61797 1 3
2 61798 1 3
2 61799 1 3
2 61800 1 3
2 61801 1 3
2 61802 1 3
2 61803 1 3
2 61804 1 3
2 61805 1 3
2 61806 1 3
2 61807 1 3
2 61808 1 3
2 61809 1 3
2 61810 1 3
2 61811 1 3
2 61812 1 3
2 61813 1 3
2 61814 1 3
2 61815 1 3
2 61816 1 3
2 61817 1 3
2 61818 1 3
2 61819 1 3
2 61820 1 3
2 61821 1 3
2 61822 1 3
2 61823 1 3
2 61824 1 3
2 61825 1 3
2 61826 1 3
2 61827 1 3
2 61828 1 3
2 61829 1 3
2 61830 1 3
2 61831 1 3
2 61832 1 3
2 61833 1 3
2 61834 1 3
2 61835 1 3
2 61836 1 3
2 61837 1 3
2 61838 1 3
2 61839 1 3
2 61840 1 3
2 61841 1 3
2 61842 1 3
2 61843 1 3
2 61844 1 3
2 61845 1 3
2 61846 1 3
2 61847 1 3
2 61848 1 3
2 61849 1 3
2 61850 1 3
2 61851 1 3
2 61852 1 3
2 61853 1 3
2 61854 1 3
2 61855 1 3
2 61856 1 3
2 61857 1 3
2 61858 1 3
2 61859 1 3
2 61860 1 3
2 61861 1 3
2 61862 1 3
2 61863 1 3
2 61864 1 3
2 61865 1 3
2 61866 1 3
2 61867 1 3
2 61868 1 3
2 61869 1 3
2 61870 1 3
2 61871 1 3
2 61872 1 3
2 61873 1 3
2 61874 1 3
2 61875 1 3
2 61876 1 3
2 61877 1 3
2 61878 1 3
2 61879 1 3
2 61880 1 3
2 61881 1 3
2 61882 1 3
2 61883 1 3
2 61884 1 3
2 61885 1 3
2 61886 1 3
2 61887 1 3
2 61888 1 3
2 61889 1 3
2 61890 1 3
2 61891 1 3
2 61892 1 3
2 61893 1 3
2 61894 1 3
2 61895 1 3
2 61896 1 3
2 61897 1 3
2 61898 1 3
2 61899 1 3
2 61900 1 3
2 61901 1 3
2 61902 1 3
2 61903 1 3
2 61904 1 3
2 61905 1 3
2 61906 1 3
2 61907 1 3
2 61908 1 3
2 61909 1 3
2 61910 1 3
2 61911 1 3
2 61912 1 3
2 61913 1 3
2 61914 1 3
2 61915 1 3
2 61916 1 3
2 61917 1 3
2 61918 1 3
2 61919 1 3
2 61920 1 3
2 61921 1 3
2 61922 1 3
2 61923 1 3
2 61924 1 3
2 61925 1 3
2 61926 1 3
2 61927 1 3
2 61928 1 3
2 61929 1 3
2 61930 1 3
2 61931 1 3
2 61932 1 3
2 61933 1 3
2 61934 1 3
2 61935 1 3
2 61936 1 3
2 61937 1 3
2 61938 1 3
2 61939 1 3
1 4 0 331 0
2 61940 1 4
2 61941 1 4
2 61942 1 4
2 61943 1 4
2 61944 1 4
2 61945 1 4
2 61946 1 4
2 61947 1 4
2 61948 1 4
2 61949 1 4
2 61950 1 4
2 61951 1 4
2 61952 1 4
2 61953 1 4
2 61954 1 4
2 61955 1 4
2 61956 1 4
2 61957 1 4
2 61958 1 4
2 61959 1 4
2 61960 1 4
2 61961 1 4
2 61962 1 4
2 61963 1 4
2 61964 1 4
2 61965 1 4
2 61966 1 4
2 61967 1 4
2 61968 1 4
2 61969 1 4
2 61970 1 4
2 61971 1 4
2 61972 1 4
2 61973 1 4
2 61974 1 4
2 61975 1 4
2 61976 1 4
2 61977 1 4
2 61978 1 4
2 61979 1 4
2 61980 1 4
2 61981 1 4
2 61982 1 4
2 61983 1 4
2 61984 1 4
2 61985 1 4
2 61986 1 4
2 61987 1 4
2 61988 1 4
2 61989 1 4
2 61990 1 4
2 61991 1 4
2 61992 1 4
2 61993 1 4
2 61994 1 4
2 61995 1 4
2 61996 1 4
2 61997 1 4
2 61998 1 4
2 61999 1 4
2 62000 1 4
2 62001 1 4
2 62002 1 4
2 62003 1 4
2 62004 1 4
2 62005 1 4
2 62006 1 4
2 62007 1 4
2 62008 1 4
2 62009 1 4
2 62010 1 4
2 62011 1 4
2 62012 1 4
2 62013 1 4
2 62014 1 4
2 62015 1 4
2 62016 1 4
2 62017 1 4
2 62018 1 4
2 62019 1 4
2 62020 1 4
2 62021 1 4
2 62022 1 4
2 62023 1 4
2 62024 1 4
2 62025 1 4
2 62026 1 4
2 62027 1 4
2 62028 1 4
2 62029 1 4
2 62030 1 4
2 62031 1 4
2 62032 1 4
2 62033 1 4
2 62034 1 4
2 62035 1 4
2 62036 1 4
2 62037 1 4
2 62038 1 4
2 62039 1 4
2 62040 1 4
2 62041 1 4
2 62042 1 4
2 62043 1 4
2 62044 1 4
2 62045 1 4
2 62046 1 4
2 62047 1 4
2 62048 1 4
2 62049 1 4
2 62050 1 4
2 62051 1 4
2 62052 1 4
2 62053 1 4
2 62054 1 4
2 62055 1 4
2 62056 1 4
2 62057 1 4
2 62058 1 4
2 62059 1 4
2 62060 1 4
2 62061 1 4
2 62062 1 4
2 62063 1 4
2 62064 1 4
2 62065 1 4
2 62066 1 4
2 62067 1 4
2 62068 1 4
2 62069 1 4
2 62070 1 4
2 62071 1 4
2 62072 1 4
2 62073 1 4
2 62074 1 4
2 62075 1 4
2 62076 1 4
2 62077 1 4
2 62078 1 4
2 62079 1 4
2 62080 1 4
2 62081 1 4
2 62082 1 4
2 62083 1 4
2 62084 1 4
2 62085 1 4
2 62086 1 4
2 62087 1 4
2 62088 1 4
2 62089 1 4
2 62090 1 4
2 62091 1 4
2 62092 1 4
2 62093 1 4
2 62094 1 4
2 62095 1 4
2 62096 1 4
2 62097 1 4
2 62098 1 4
2 62099 1 4
2 62100 1 4
2 62101 1 4
2 62102 1 4
2 62103 1 4
2 62104 1 4
2 62105 1 4
2 62106 1 4
2 62107 1 4
2 62108 1 4
2 62109 1 4
2 62110 1 4
2 62111 1 4
2 62112 1 4
2 62113 1 4
2 62114 1 4
2 62115 1 4
2 62116 1 4
2 62117 1 4
2 62118 1 4
2 62119 1 4
2 62120 1 4
2 62121 1 4
2 62122 1 4
2 62123 1 4
2 62124 1 4
2 62125 1 4
2 62126 1 4
2 62127 1 4
2 62128 1 4
2 62129 1 4
2 62130 1 4
2 62131 1 4
2 62132 1 4
2 62133 1 4
2 62134 1 4
2 62135 1 4
2 62136 1 4
2 62137 1 4
2 62138 1 4
2 62139 1 4
2 62140 1 4
2 62141 1 4
2 62142 1 4
2 62143 1 4
2 62144 1 4
2 62145 1 4
2 62146 1 4
2 62147 1 4
2 62148 1 4
2 62149 1 4
2 62150 1 4
2 62151 1 4
2 62152 1 4
2 62153 1 4
2 62154 1 4
2 62155 1 4
2 62156 1 4
2 62157 1 4
2 62158 1 4
2 62159 1 4
2 62160 1 4
2 62161 1 4
2 62162 1 4
2 62163 1 4
2 62164 1 4
2 62165 1 4
2 62166 1 4
2 62167 1 4
2 62168 1 4
2 62169 1 4
2 62170 1 4
2 62171 1 4
2 62172 1 4
2 62173 1 4
2 62174 1 4
2 62175 1 4
2 62176 1 4
2 62177 1 4
2 62178 1 4
2 62179 1 4
2 62180 1 4
2 62181 1 4
2 62182 1 4
2 62183 1 4
2 62184 1 4
2 62185 1 4
2 62186 1 4
2 62187 1 4
2 62188 1 4
2 62189 1 4
2 62190 1 4
2 62191 1 4
2 62192 1 4
2 62193 1 4
2 62194 1 4
2 62195 1 4
2 62196 1 4
2 62197 1 4
2 62198 1 4
2 62199 1 4
2 62200 1 4
2 62201 1 4
2 62202 1 4
2 62203 1 4
2 62204 1 4
2 62205 1 4
2 62206 1 4
2 62207 1 4
2 62208 1 4
2 62209 1 4
2 62210 1 4
2 62211 1 4
2 62212 1 4
2 62213 1 4
2 62214 1 4
2 62215 1 4
2 62216 1 4
2 62217 1 4
2 62218 1 4
2 62219 1 4
2 62220 1 4
2 62221 1 4
2 62222 1 4
2 62223 1 4
2 62224 1 4
2 62225 1 4
2 62226 1 4
2 62227 1 4
2 62228 1 4
2 62229 1 4
2 62230 1 4
2 62231 1 4
2 62232 1 4
2 62233 1 4
2 62234 1 4
2 62235 1 4
2 62236 1 4
2 62237 1 4
2 62238 1 4
2 62239 1 4
2 62240 1 4
2 62241 1 4
2 62242 1 4
2 62243 1 4
2 62244 1 4
2 62245 1 4
2 62246 1 4
2 62247 1 4
2 62248 1 4
2 62249 1 4
2 62250 1 4
2 62251 1 4
2 62252 1 4
2 62253 1 4
2 62254 1 4
2 62255 1 4
2 62256 1 4
2 62257 1 4
2 62258 1 4
2 62259 1 4
2 62260 1 4
2 62261 1 4
2 62262 1 4
2 62263 1 4
2 62264 1 4
2 62265 1 4
2 62266 1 4
2 62267 1 4
2 62268 1 4
2 62269 1 4
2 62270 1 4
1 5 0 189 0
2 62271 1 5
2 62272 1 5
2 62273 1 5
2 62274 1 5
2 62275 1 5
2 62276 1 5
2 62277 1 5
2 62278 1 5
2 62279 1 5
2 62280 1 5
2 62281 1 5
2 62282 1 5
2 62283 1 5
2 62284 1 5
2 62285 1 5
2 62286 1 5
2 62287 1 5
2 62288 1 5
2 62289 1 5
2 62290 1 5
2 62291 1 5
2 62292 1 5
2 62293 1 5
2 62294 1 5
2 62295 1 5
2 62296 1 5
2 62297 1 5
2 62298 1 5
2 62299 1 5
2 62300 1 5
2 62301 1 5
2 62302 1 5
2 62303 1 5
2 62304 1 5
2 62305 1 5
2 62306 1 5
2 62307 1 5
2 62308 1 5
2 62309 1 5
2 62310 1 5
2 62311 1 5
2 62312 1 5
2 62313 1 5
2 62314 1 5
2 62315 1 5
2 62316 1 5
2 62317 1 5
2 62318 1 5
2 62319 1 5
2 62320 1 5
2 62321 1 5
2 62322 1 5
2 62323 1 5
2 62324 1 5
2 62325 1 5
2 62326 1 5
2 62327 1 5
2 62328 1 5
2 62329 1 5
2 62330 1 5
2 62331 1 5
2 62332 1 5
2 62333 1 5
2 62334 1 5
2 62335 1 5
2 62336 1 5
2 62337 1 5
2 62338 1 5
2 62339 1 5
2 62340 1 5
2 62341 1 5
2 62342 1 5
2 62343 1 5
2 62344 1 5
2 62345 1 5
2 62346 1 5
2 62347 1 5
2 62348 1 5
2 62349 1 5
2 62350 1 5
2 62351 1 5
2 62352 1 5
2 62353 1 5
2 62354 1 5
2 62355 1 5
2 62356 1 5
2 62357 1 5
2 62358 1 5
2 62359 1 5
2 62360 1 5
2 62361 1 5
2 62362 1 5
2 62363 1 5
2 62364 1 5
2 62365 1 5
2 62366 1 5
2 62367 1 5
2 62368 1 5
2 62369 1 5
2 62370 1 5
2 62371 1 5
2 62372 1 5
2 62373 1 5
2 62374 1 5
2 62375 1 5
2 62376 1 5
2 62377 1 5
2 62378 1 5
2 62379 1 5
2 62380 1 5
2 62381 1 5
2 62382 1 5
2 62383 1 5
2 62384 1 5
2 62385 1 5
2 62386 1 5
2 62387 1 5
2 62388 1 5
2 62389 1 5
2 62390 1 5
2 62391 1 5
2 62392 1 5
2 62393 1 5
2 62394 1 5
2 62395 1 5
2 62396 1 5
2 62397 1 5
2 62398 1 5
2 62399 1 5
2 62400 1 5
2 62401 1 5
2 62402 1 5
2 62403 1 5
2 62404 1 5
2 62405 1 5
2 62406 1 5
2 62407 1 5
2 62408 1 5
2 62409 1 5
2 62410 1 5
2 62411 1 5
2 62412 1 5
2 62413 1 5
2 62414 1 5
2 62415 1 5
2 62416 1 5
2 62417 1 5
2 62418 1 5
2 62419 1 5
2 62420 1 5
2 62421 1 5
2 62422 1 5
2 62423 1 5
2 62424 1 5
2 62425 1 5
2 62426 1 5
2 62427 1 5
2 62428 1 5
2 62429 1 5
2 62430 1 5
2 62431 1 5
2 62432 1 5
2 62433 1 5
2 62434 1 5
2 62435 1 5
2 62436 1 5
2 62437 1 5
2 62438 1 5
2 62439 1 5
2 62440 1 5
2 62441 1 5
2 62442 1 5
2 62443 1 5
2 62444 1 5
2 62445 1 5
2 62446 1 5
2 62447 1 5
2 62448 1 5
2 62449 1 5
2 62450 1 5
2 62451 1 5
2 62452 1 5
2 62453 1 5
2 62454 1 5
2 62455 1 5
2 62456 1 5
2 62457 1 5
2 62458 1 5
2 62459 1 5
1 6 0 235 0
2 62460 1 6
2 62461 1 6
2 62462 1 6
2 62463 1 6
2 62464 1 6
2 62465 1 6
2 62466 1 6
2 62467 1 6
2 62468 1 6
2 62469 1 6
2 62470 1 6
2 62471 1 6
2 62472 1 6
2 62473 1 6
2 62474 1 6
2 62475 1 6
2 62476 1 6
2 62477 1 6
2 62478 1 6
2 62479 1 6
2 62480 1 6
2 62481 1 6
2 62482 1 6
2 62483 1 6
2 62484 1 6
2 62485 1 6
2 62486 1 6
2 62487 1 6
2 62488 1 6
2 62489 1 6
2 62490 1 6
2 62491 1 6
2 62492 1 6
2 62493 1 6
2 62494 1 6
2 62495 1 6
2 62496 1 6
2 62497 1 6
2 62498 1 6
2 62499 1 6
2 62500 1 6
2 62501 1 6
2 62502 1 6
2 62503 1 6
2 62504 1 6
2 62505 1 6
2 62506 1 6
2 62507 1 6
2 62508 1 6
2 62509 1 6
2 62510 1 6
2 62511 1 6
2 62512 1 6
2 62513 1 6
2 62514 1 6
2 62515 1 6
2 62516 1 6
2 62517 1 6
2 62518 1 6
2 62519 1 6
2 62520 1 6
2 62521 1 6
2 62522 1 6
2 62523 1 6
2 62524 1 6
2 62525 1 6
2 62526 1 6
2 62527 1 6
2 62528 1 6
2 62529 1 6
2 62530 1 6
2 62531 1 6
2 62532 1 6
2 62533 1 6
2 62534 1 6
2 62535 1 6
2 62536 1 6
2 62537 1 6
2 62538 1 6
2 62539 1 6
2 62540 1 6
2 62541 1 6
2 62542 1 6
2 62543 1 6
2 62544 1 6
2 62545 1 6
2 62546 1 6
2 62547 1 6
2 62548 1 6
2 62549 1 6
2 62550 1 6
2 62551 1 6
2 62552 1 6
2 62553 1 6
2 62554 1 6
2 62555 1 6
2 62556 1 6
2 62557 1 6
2 62558 1 6
2 62559 1 6
2 62560 1 6
2 62561 1 6
2 62562 1 6
2 62563 1 6
2 62564 1 6
2 62565 1 6
2 62566 1 6
2 62567 1 6
2 62568 1 6
2 62569 1 6
2 62570 1 6
2 62571 1 6
2 62572 1 6
2 62573 1 6
2 62574 1 6
2 62575 1 6
2 62576 1 6
2 62577 1 6
2 62578 1 6
2 62579 1 6
2 62580 1 6
2 62581 1 6
2 62582 1 6
2 62583 1 6
2 62584 1 6
2 62585 1 6
2 62586 1 6
2 62587 1 6
2 62588 1 6
2 62589 1 6
2 62590 1 6
2 62591 1 6
2 62592 1 6
2 62593 1 6
2 62594 1 6
2 62595 1 6
2 62596 1 6
2 62597 1 6
2 62598 1 6
2 62599 1 6
2 62600 1 6
2 62601 1 6
2 62602 1 6
2 62603 1 6
2 62604 1 6
2 62605 1 6
2 62606 1 6
2 62607 1 6
2 62608 1 6
2 62609 1 6
2 62610 1 6
2 62611 1 6
2 62612 1 6
2 62613 1 6
2 62614 1 6
2 62615 1 6
2 62616 1 6
2 62617 1 6
2 62618 1 6
2 62619 1 6
2 62620 1 6
2 62621 1 6
2 62622 1 6
2 62623 1 6
2 62624 1 6
2 62625 1 6
2 62626 1 6
2 62627 1 6
2 62628 1 6
2 62629 1 6
2 62630 1 6
2 62631 1 6
2 62632 1 6
2 62633 1 6
2 62634 1 6
2 62635 1 6
2 62636 1 6
2 62637 1 6
2 62638 1 6
2 62639 1 6
2 62640 1 6
2 62641 1 6
2 62642 1 6
2 62643 1 6
2 62644 1 6
2 62645 1 6
2 62646 1 6
2 62647 1 6
2 62648 1 6
2 62649 1 6
2 62650 1 6
2 62651 1 6
2 62652 1 6
2 62653 1 6
2 62654 1 6
2 62655 1 6
2 62656 1 6
2 62657 1 6
2 62658 1 6
2 62659 1 6
2 62660 1 6
2 62661 1 6
2 62662 1 6
2 62663 1 6
2 62664 1 6
2 62665 1 6
2 62666 1 6
2 62667 1 6
2 62668 1 6
2 62669 1 6
2 62670 1 6
2 62671 1 6
2 62672 1 6
2 62673 1 6
2 62674 1 6
2 62675 1 6
2 62676 1 6
2 62677 1 6
2 62678 1 6
2 62679 1 6
2 62680 1 6
2 62681 1 6
2 62682 1 6
2 62683 1 6
2 62684 1 6
2 62685 1 6
2 62686 1 6
2 62687 1 6
2 62688 1 6
2 62689 1 6
2 62690 1 6
2 62691 1 6
2 62692 1 6
2 62693 1 6
2 62694 1 6
1 7 0 243 0
2 62695 1 7
2 62696 1 7
2 62697 1 7
2 62698 1 7
2 62699 1 7
2 62700 1 7
2 62701 1 7
2 62702 1 7
2 62703 1 7
2 62704 1 7
2 62705 1 7
2 62706 1 7
2 62707 1 7
2 62708 1 7
2 62709 1 7
2 62710 1 7
2 62711 1 7
2 62712 1 7
2 62713 1 7
2 62714 1 7
2 62715 1 7
2 62716 1 7
2 62717 1 7
2 62718 1 7
2 62719 1 7
2 62720 1 7
2 62721 1 7
2 62722 1 7
2 62723 1 7
2 62724 1 7
2 62725 1 7
2 62726 1 7
2 62727 1 7
2 62728 1 7
2 62729 1 7
2 62730 1 7
2 62731 1 7
2 62732 1 7
2 62733 1 7
2 62734 1 7
2 62735 1 7
2 62736 1 7
2 62737 1 7
2 62738 1 7
2 62739 1 7
2 62740 1 7
2 62741 1 7
2 62742 1 7
2 62743 1 7
2 62744 1 7
2 62745 1 7
2 62746 1 7
2 62747 1 7
2 62748 1 7
2 62749 1 7
2 62750 1 7
2 62751 1 7
2 62752 1 7
2 62753 1 7
2 62754 1 7
2 62755 1 7
2 62756 1 7
2 62757 1 7
2 62758 1 7
2 62759 1 7
2 62760 1 7
2 62761 1 7
2 62762 1 7
2 62763 1 7
2 62764 1 7
2 62765 1 7
2 62766 1 7
2 62767 1 7
2 62768 1 7
2 62769 1 7
2 62770 1 7
2 62771 1 7
2 62772 1 7
2 62773 1 7
2 62774 1 7
2 62775 1 7
2 62776 1 7
2 62777 1 7
2 62778 1 7
2 62779 1 7
2 62780 1 7
2 62781 1 7
2 62782 1 7
2 62783 1 7
2 62784 1 7
2 62785 1 7
2 62786 1 7
2 62787 1 7
2 62788 1 7
2 62789 1 7
2 62790 1 7
2 62791 1 7
2 62792 1 7
2 62793 1 7
2 62794 1 7
2 62795 1 7
2 62796 1 7
2 62797 1 7
2 62798 1 7
2 62799 1 7
2 62800 1 7
2 62801 1 7
2 62802 1 7
2 62803 1 7
2 62804 1 7
2 62805 1 7
2 62806 1 7
2 62807 1 7
2 62808 1 7
2 62809 1 7
2 62810 1 7
2 62811 1 7
2 62812 1 7
2 62813 1 7
2 62814 1 7
2 62815 1 7
2 62816 1 7
2 62817 1 7
2 62818 1 7
2 62819 1 7
2 62820 1 7
2 62821 1 7
2 62822 1 7
2 62823 1 7
2 62824 1 7
2 62825 1 7
2 62826 1 7
2 62827 1 7
2 62828 1 7
2 62829 1 7
2 62830 1 7
2 62831 1 7
2 62832 1 7
2 62833 1 7
2 62834 1 7
2 62835 1 7
2 62836 1 7
2 62837 1 7
2 62838 1 7
2 62839 1 7
2 62840 1 7
2 62841 1 7
2 62842 1 7
2 62843 1 7
2 62844 1 7
2 62845 1 7
2 62846 1 7
2 62847 1 7
2 62848 1 7
2 62849 1 7
2 62850 1 7
2 62851 1 7
2 62852 1 7
2 62853 1 7
2 62854 1 7
2 62855 1 7
2 62856 1 7
2 62857 1 7
2 62858 1 7
2 62859 1 7
2 62860 1 7
2 62861 1 7
2 62862 1 7
2 62863 1 7
2 62864 1 7
2 62865 1 7
2 62866 1 7
2 62867 1 7
2 62868 1 7
2 62869 1 7
2 62870 1 7
2 62871 1 7
2 62872 1 7
2 62873 1 7
2 62874 1 7
2 62875 1 7
2 62876 1 7
2 62877 1 7
2 62878 1 7
2 62879 1 7
2 62880 1 7
2 62881 1 7
2 62882 1 7
2 62883 1 7
2 62884 1 7
2 62885 1 7
2 62886 1 7
2 62887 1 7
2 62888 1 7
2 62889 1 7
2 62890 1 7
2 62891 1 7
2 62892 1 7
2 62893 1 7
2 62894 1 7
2 62895 1 7
2 62896 1 7
2 62897 1 7
2 62898 1 7
2 62899 1 7
2 62900 1 7
2 62901 1 7
2 62902 1 7
2 62903 1 7
2 62904 1 7
2 62905 1 7
2 62906 1 7
2 62907 1 7
2 62908 1 7
2 62909 1 7
2 62910 1 7
2 62911 1 7
2 62912 1 7
2 62913 1 7
2 62914 1 7
2 62915 1 7
2 62916 1 7
2 62917 1 7
2 62918 1 7
2 62919 1 7
2 62920 1 7
2 62921 1 7
2 62922 1 7
2 62923 1 7
2 62924 1 7
2 62925 1 7
2 62926 1 7
2 62927 1 7
2 62928 1 7
2 62929 1 7
2 62930 1 7
2 62931 1 7
2 62932 1 7
2 62933 1 7
2 62934 1 7
2 62935 1 7
2 62936 1 7
2 62937 1 7
1 8 0 55 0
2 62938 1 8
2 62939 1 8
2 62940 1 8
2 62941 1 8
2 62942 1 8
2 62943 1 8
2 62944 1 8
2 62945 1 8
2 62946 1 8
2 62947 1 8
2 62948 1 8
2 62949 1 8
2 62950 1 8
2 62951 1 8
2 62952 1 8
2 62953 1 8
2 62954 1 8
2 62955 1 8
2 62956 1 8
2 62957 1 8
2 62958 1 8
2 62959 1 8
2 62960 1 8
2 62961 1 8
2 62962 1 8
2 62963 1 8
2 62964 1 8
2 62965 1 8
2 62966 1 8
2 62967 1 8
2 62968 1 8
2 62969 1 8
2 62970 1 8
2 62971 1 8
2 62972 1 8
2 62973 1 8
2 62974 1 8
2 62975 1 8
2 62976 1 8
2 62977 1 8
2 62978 1 8
2 62979 1 8
2 62980 1 8
2 62981 1 8
2 62982 1 8
2 62983 1 8
2 62984 1 8
2 62985 1 8
2 62986 1 8
2 62987 1 8
2 62988 1 8
2 62989 1 8
2 62990 1 8
2 62991 1 8
2 62992 1 8
1 9 0 52 0
2 62993 1 9
2 62994 1 9
2 62995 1 9
2 62996 1 9
2 62997 1 9
2 62998 1 9
2 62999 1 9
2 63000 1 9
2 63001 1 9
2 63002 1 9
2 63003 1 9
2 63004 1 9
2 63005 1 9
2 63006 1 9
2 63007 1 9
2 63008 1 9
2 63009 1 9
2 63010 1 9
2 63011 1 9
2 63012 1 9
2 63013 1 9
2 63014 1 9
2 63015 1 9
2 63016 1 9
2 63017 1 9
2 63018 1 9
2 63019 1 9
2 63020 1 9
2 63021 1 9
2 63022 1 9
2 63023 1 9
2 63024 1 9
2 63025 1 9
2 63026 1 9
2 63027 1 9
2 63028 1 9
2 63029 1 9
2 63030 1 9
2 63031 1 9
2 63032 1 9
2 63033 1 9
2 63034 1 9
2 63035 1 9
2 63036 1 9
2 63037 1 9
2 63038 1 9
2 63039 1 9
2 63040 1 9
2 63041 1 9
2 63042 1 9
2 63043 1 9
2 63044 1 9
1 10 0 171 0
2 63045 1 10
2 63046 1 10
2 63047 1 10
2 63048 1 10
2 63049 1 10
2 63050 1 10
2 63051 1 10
2 63052 1 10
2 63053 1 10
2 63054 1 10
2 63055 1 10
2 63056 1 10
2 63057 1 10
2 63058 1 10
2 63059 1 10
2 63060 1 10
2 63061 1 10
2 63062 1 10
2 63063 1 10
2 63064 1 10
2 63065 1 10
2 63066 1 10
2 63067 1 10
2 63068 1 10
2 63069 1 10
2 63070 1 10
2 63071 1 10
2 63072 1 10
2 63073 1 10
2 63074 1 10
2 63075 1 10
2 63076 1 10
2 63077 1 10
2 63078 1 10
2 63079 1 10
2 63080 1 10
2 63081 1 10
2 63082 1 10
2 63083 1 10
2 63084 1 10
2 63085 1 10
2 63086 1 10
2 63087 1 10
2 63088 1 10
2 63089 1 10
2 63090 1 10
2 63091 1 10
2 63092 1 10
2 63093 1 10
2 63094 1 10
2 63095 1 10
2 63096 1 10
2 63097 1 10
2 63098 1 10
2 63099 1 10
2 63100 1 10
2 63101 1 10
2 63102 1 10
2 63103 1 10
2 63104 1 10
2 63105 1 10
2 63106 1 10
2 63107 1 10
2 63108 1 10
2 63109 1 10
2 63110 1 10
2 63111 1 10
2 63112 1 10
2 63113 1 10
2 63114 1 10
2 63115 1 10
2 63116 1 10
2 63117 1 10
2 63118 1 10
2 63119 1 10
2 63120 1 10
2 63121 1 10
2 63122 1 10
2 63123 1 10
2 63124 1 10
2 63125 1 10
2 63126 1 10
2 63127 1 10
2 63128 1 10
2 63129 1 10
2 63130 1 10
2 63131 1 10
2 63132 1 10
2 63133 1 10
2 63134 1 10
2 63135 1 10
2 63136 1 10
2 63137 1 10
2 63138 1 10
2 63139 1 10
2 63140 1 10
2 63141 1 10
2 63142 1 10
2 63143 1 10
2 63144 1 10
2 63145 1 10
2 63146 1 10
2 63147 1 10
2 63148 1 10
2 63149 1 10
2 63150 1 10
2 63151 1 10
2 63152 1 10
2 63153 1 10
2 63154 1 10
2 63155 1 10
2 63156 1 10
2 63157 1 10
2 63158 1 10
2 63159 1 10
2 63160 1 10
2 63161 1 10
2 63162 1 10
2 63163 1 10
2 63164 1 10
2 63165 1 10
2 63166 1 10
2 63167 1 10
2 63168 1 10
2 63169 1 10
2 63170 1 10
2 63171 1 10
2 63172 1 10
2 63173 1 10
2 63174 1 10
2 63175 1 10
2 63176 1 10
2 63177 1 10
2 63178 1 10
2 63179 1 10
2 63180 1 10
2 63181 1 10
2 63182 1 10
2 63183 1 10
2 63184 1 10
2 63185 1 10
2 63186 1 10
2 63187 1 10
2 63188 1 10
2 63189 1 10
2 63190 1 10
2 63191 1 10
2 63192 1 10
2 63193 1 10
2 63194 1 10
2 63195 1 10
2 63196 1 10
2 63197 1 10
2 63198 1 10
2 63199 1 10
2 63200 1 10
2 63201 1 10
2 63202 1 10
2 63203 1 10
2 63204 1 10
2 63205 1 10
2 63206 1 10
2 63207 1 10
2 63208 1 10
2 63209 1 10
2 63210 1 10
2 63211 1 10
2 63212 1 10
2 63213 1 10
2 63214 1 10
2 63215 1 10
1 11 0 201 0
2 63216 1 11
2 63217 1 11
2 63218 1 11
2 63219 1 11
2 63220 1 11
2 63221 1 11
2 63222 1 11
2 63223 1 11
2 63224 1 11
2 63225 1 11
2 63226 1 11
2 63227 1 11
2 63228 1 11
2 63229 1 11
2 63230 1 11
2 63231 1 11
2 63232 1 11
2 63233 1 11
2 63234 1 11
2 63235 1 11
2 63236 1 11
2 63237 1 11
2 63238 1 11
2 63239 1 11
2 63240 1 11
2 63241 1 11
2 63242 1 11
2 63243 1 11
2 63244 1 11
2 63245 1 11
2 63246 1 11
2 63247 1 11
2 63248 1 11
2 63249 1 11
2 63250 1 11
2 63251 1 11
2 63252 1 11
2 63253 1 11
2 63254 1 11
2 63255 1 11
2 63256 1 11
2 63257 1 11
2 63258 1 11
2 63259 1 11
2 63260 1 11
2 63261 1 11
2 63262 1 11
2 63263 1 11
2 63264 1 11
2 63265 1 11
2 63266 1 11
2 63267 1 11
2 63268 1 11
2 63269 1 11
2 63270 1 11
2 63271 1 11
2 63272 1 11
2 63273 1 11
2 63274 1 11
2 63275 1 11
2 63276 1 11
2 63277 1 11
2 63278 1 11
2 63279 1 11
2 63280 1 11
2 63281 1 11
2 63282 1 11
2 63283 1 11
2 63284 1 11
2 63285 1 11
2 63286 1 11
2 63287 1 11
2 63288 1 11
2 63289 1 11
2 63290 1 11
2 63291 1 11
2 63292 1 11
2 63293 1 11
2 63294 1 11
2 63295 1 11
2 63296 1 11
2 63297 1 11
2 63298 1 11
2 63299 1 11
2 63300 1 11
2 63301 1 11
2 63302 1 11
2 63303 1 11
2 63304 1 11
2 63305 1 11
2 63306 1 11
2 63307 1 11
2 63308 1 11
2 63309 1 11
2 63310 1 11
2 63311 1 11
2 63312 1 11
2 63313 1 11
2 63314 1 11
2 63315 1 11
2 63316 1 11
2 63317 1 11
2 63318 1 11
2 63319 1 11
2 63320 1 11
2 63321 1 11
2 63322 1 11
2 63323 1 11
2 63324 1 11
2 63325 1 11
2 63326 1 11
2 63327 1 11
2 63328 1 11
2 63329 1 11
2 63330 1 11
2 63331 1 11
2 63332 1 11
2 63333 1 11
2 63334 1 11
2 63335 1 11
2 63336 1 11
2 63337 1 11
2 63338 1 11
2 63339 1 11
2 63340 1 11
2 63341 1 11
2 63342 1 11
2 63343 1 11
2 63344 1 11
2 63345 1 11
2 63346 1 11
2 63347 1 11
2 63348 1 11
2 63349 1 11
2 63350 1 11
2 63351 1 11
2 63352 1 11
2 63353 1 11
2 63354 1 11
2 63355 1 11
2 63356 1 11
2 63357 1 11
2 63358 1 11
2 63359 1 11
2 63360 1 11
2 63361 1 11
2 63362 1 11
2 63363 1 11
2 63364 1 11
2 63365 1 11
2 63366 1 11
2 63367 1 11
2 63368 1 11
2 63369 1 11
2 63370 1 11
2 63371 1 11
2 63372 1 11
2 63373 1 11
2 63374 1 11
2 63375 1 11
2 63376 1 11
2 63377 1 11
2 63378 1 11
2 63379 1 11
2 63380 1 11
2 63381 1 11
2 63382 1 11
2 63383 1 11
2 63384 1 11
2 63385 1 11
2 63386 1 11
2 63387 1 11
2 63388 1 11
2 63389 1 11
2 63390 1 11
2 63391 1 11
2 63392 1 11
2 63393 1 11
2 63394 1 11
2 63395 1 11
2 63396 1 11
2 63397 1 11
2 63398 1 11
2 63399 1 11
2 63400 1 11
2 63401 1 11
2 63402 1 11
2 63403 1 11
2 63404 1 11
2 63405 1 11
2 63406 1 11
2 63407 1 11
2 63408 1 11
2 63409 1 11
2 63410 1 11
2 63411 1 11
2 63412 1 11
2 63413 1 11
2 63414 1 11
2 63415 1 11
2 63416 1 11
1 12 0 239 0
2 63417 1 12
2 63418 1 12
2 63419 1 12
2 63420 1 12
2 63421 1 12
2 63422 1 12
2 63423 1 12
2 63424 1 12
2 63425 1 12
2 63426 1 12
2 63427 1 12
2 63428 1 12
2 63429 1 12
2 63430 1 12
2 63431 1 12
2 63432 1 12
2 63433 1 12
2 63434 1 12
2 63435 1 12
2 63436 1 12
2 63437 1 12
2 63438 1 12
2 63439 1 12
2 63440 1 12
2 63441 1 12
2 63442 1 12
2 63443 1 12
2 63444 1 12
2 63445 1 12
2 63446 1 12
2 63447 1 12
2 63448 1 12
2 63449 1 12
2 63450 1 12
2 63451 1 12
2 63452 1 12
2 63453 1 12
2 63454 1 12
2 63455 1 12
2 63456 1 12
2 63457 1 12
2 63458 1 12
2 63459 1 12
2 63460 1 12
2 63461 1 12
2 63462 1 12
2 63463 1 12
2 63464 1 12
2 63465 1 12
2 63466 1 12
2 63467 1 12
2 63468 1 12
2 63469 1 12
2 63470 1 12
2 63471 1 12
2 63472 1 12
2 63473 1 12
2 63474 1 12
2 63475 1 12
2 63476 1 12
2 63477 1 12
2 63478 1 12
2 63479 1 12
2 63480 1 12
2 63481 1 12
2 63482 1 12
2 63483 1 12
2 63484 1 12
2 63485 1 12
2 63486 1 12
2 63487 1 12
2 63488 1 12
2 63489 1 12
2 63490 1 12
2 63491 1 12
2 63492 1 12
2 63493 1 12
2 63494 1 12
2 63495 1 12
2 63496 1 12
2 63497 1 12
2 63498 1 12
2 63499 1 12
2 63500 1 12
2 63501 1 12
2 63502 1 12
2 63503 1 12
2 63504 1 12
2 63505 1 12
2 63506 1 12
2 63507 1 12
2 63508 1 12
2 63509 1 12
2 63510 1 12
2 63511 1 12
2 63512 1 12
2 63513 1 12
2 63514 1 12
2 63515 1 12
2 63516 1 12
2 63517 1 12
2 63518 1 12
2 63519 1 12
2 63520 1 12
2 63521 1 12
2 63522 1 12
2 63523 1 12
2 63524 1 12
2 63525 1 12
2 63526 1 12
2 63527 1 12
2 63528 1 12
2 63529 1 12
2 63530 1 12
2 63531 1 12
2 63532 1 12
2 63533 1 12
2 63534 1 12
2 63535 1 12
2 63536 1 12
2 63537 1 12
2 63538 1 12
2 63539 1 12
2 63540 1 12
2 63541 1 12
2 63542 1 12
2 63543 1 12
2 63544 1 12
2 63545 1 12
2 63546 1 12
2 63547 1 12
2 63548 1 12
2 63549 1 12
2 63550 1 12
2 63551 1 12
2 63552 1 12
2 63553 1 12
2 63554 1 12
2 63555 1 12
2 63556 1 12
2 63557 1 12
2 63558 1 12
2 63559 1 12
2 63560 1 12
2 63561 1 12
2 63562 1 12
2 63563 1 12
2 63564 1 12
2 63565 1 12
2 63566 1 12
2 63567 1 12
2 63568 1 12
2 63569 1 12
2 63570 1 12
2 63571 1 12
2 63572 1 12
2 63573 1 12
2 63574 1 12
2 63575 1 12
2 63576 1 12
2 63577 1 12
2 63578 1 12
2 63579 1 12
2 63580 1 12
2 63581 1 12
2 63582 1 12
2 63583 1 12
2 63584 1 12
2 63585 1 12
2 63586 1 12
2 63587 1 12
2 63588 1 12
2 63589 1 12
2 63590 1 12
2 63591 1 12
2 63592 1 12
2 63593 1 12
2 63594 1 12
2 63595 1 12
2 63596 1 12
2 63597 1 12
2 63598 1 12
2 63599 1 12
2 63600 1 12
2 63601 1 12
2 63602 1 12
2 63603 1 12
2 63604 1 12
2 63605 1 12
2 63606 1 12
2 63607 1 12
2 63608 1 12
2 63609 1 12
2 63610 1 12
2 63611 1 12
2 63612 1 12
2 63613 1 12
2 63614 1 12
2 63615 1 12
2 63616 1 12
2 63617 1 12
2 63618 1 12
2 63619 1 12
2 63620 1 12
2 63621 1 12
2 63622 1 12
2 63623 1 12
2 63624 1 12
2 63625 1 12
2 63626 1 12
2 63627 1 12
2 63628 1 12
2 63629 1 12
2 63630 1 12
2 63631 1 12
2 63632 1 12
2 63633 1 12
2 63634 1 12
2 63635 1 12
2 63636 1 12
2 63637 1 12
2 63638 1 12
2 63639 1 12
2 63640 1 12
2 63641 1 12
2 63642 1 12
2 63643 1 12
2 63644 1 12
2 63645 1 12
2 63646 1 12
2 63647 1 12
2 63648 1 12
2 63649 1 12
2 63650 1 12
2 63651 1 12
2 63652 1 12
2 63653 1 12
2 63654 1 12
2 63655 1 12
1 13 0 208 0
2 63656 1 13
2 63657 1 13
2 63658 1 13
2 63659 1 13
2 63660 1 13
2 63661 1 13
2 63662 1 13
2 63663 1 13
2 63664 1 13
2 63665 1 13
2 63666 1 13
2 63667 1 13
2 63668 1 13
2 63669 1 13
2 63670 1 13
2 63671 1 13
2 63672 1 13
2 63673 1 13
2 63674 1 13
2 63675 1 13
2 63676 1 13
2 63677 1 13
2 63678 1 13
2 63679 1 13
2 63680 1 13
2 63681 1 13
2 63682 1 13
2 63683 1 13
2 63684 1 13
2 63685 1 13
2 63686 1 13
2 63687 1 13
2 63688 1 13
2 63689 1 13
2 63690 1 13
2 63691 1 13
2 63692 1 13
2 63693 1 13
2 63694 1 13
2 63695 1 13
2 63696 1 13
2 63697 1 13
2 63698 1 13
2 63699 1 13
2 63700 1 13
2 63701 1 13
2 63702 1 13
2 63703 1 13
2 63704 1 13
2 63705 1 13
2 63706 1 13
2 63707 1 13
2 63708 1 13
2 63709 1 13
2 63710 1 13
2 63711 1 13
2 63712 1 13
2 63713 1 13
2 63714 1 13
2 63715 1 13
2 63716 1 13
2 63717 1 13
2 63718 1 13
2 63719 1 13
2 63720 1 13
2 63721 1 13
2 63722 1 13
2 63723 1 13
2 63724 1 13
2 63725 1 13
2 63726 1 13
2 63727 1 13
2 63728 1 13
2 63729 1 13
2 63730 1 13
2 63731 1 13
2 63732 1 13
2 63733 1 13
2 63734 1 13
2 63735 1 13
2 63736 1 13
2 63737 1 13
2 63738 1 13
2 63739 1 13
2 63740 1 13
2 63741 1 13
2 63742 1 13
2 63743 1 13
2 63744 1 13
2 63745 1 13
2 63746 1 13
2 63747 1 13
2 63748 1 13
2 63749 1 13
2 63750 1 13
2 63751 1 13
2 63752 1 13
2 63753 1 13
2 63754 1 13
2 63755 1 13
2 63756 1 13
2 63757 1 13
2 63758 1 13
2 63759 1 13
2 63760 1 13
2 63761 1 13
2 63762 1 13
2 63763 1 13
2 63764 1 13
2 63765 1 13
2 63766 1 13
2 63767 1 13
2 63768 1 13
2 63769 1 13
2 63770 1 13
2 63771 1 13
2 63772 1 13
2 63773 1 13
2 63774 1 13
2 63775 1 13
2 63776 1 13
2 63777 1 13
2 63778 1 13
2 63779 1 13
2 63780 1 13
2 63781 1 13
2 63782 1 13
2 63783 1 13
2 63784 1 13
2 63785 1 13
2 63786 1 13
2 63787 1 13
2 63788 1 13
2 63789 1 13
2 63790 1 13
2 63791 1 13
2 63792 1 13
2 63793 1 13
2 63794 1 13
2 63795 1 13
2 63796 1 13
2 63797 1 13
2 63798 1 13
2 63799 1 13
2 63800 1 13
2 63801 1 13
2 63802 1 13
2 63803 1 13
2 63804 1 13
2 63805 1 13
2 63806 1 13
2 63807 1 13
2 63808 1 13
2 63809 1 13
2 63810 1 13
2 63811 1 13
2 63812 1 13
2 63813 1 13
2 63814 1 13
2 63815 1 13
2 63816 1 13
2 63817 1 13
2 63818 1 13
2 63819 1 13
2 63820 1 13
2 63821 1 13
2 63822 1 13
2 63823 1 13
2 63824 1 13
2 63825 1 13
2 63826 1 13
2 63827 1 13
2 63828 1 13
2 63829 1 13
2 63830 1 13
2 63831 1 13
2 63832 1 13
2 63833 1 13
2 63834 1 13
2 63835 1 13
2 63836 1 13
2 63837 1 13
2 63838 1 13
2 63839 1 13
2 63840 1 13
2 63841 1 13
2 63842 1 13
2 63843 1 13
2 63844 1 13
2 63845 1 13
2 63846 1 13
2 63847 1 13
2 63848 1 13
2 63849 1 13
2 63850 1 13
2 63851 1 13
2 63852 1 13
2 63853 1 13
2 63854 1 13
2 63855 1 13
2 63856 1 13
2 63857 1 13
2 63858 1 13
2 63859 1 13
2 63860 1 13
2 63861 1 13
2 63862 1 13
2 63863 1 13
1 14 0 154 0
2 63864 1 14
2 63865 1 14
2 63866 1 14
2 63867 1 14
2 63868 1 14
2 63869 1 14
2 63870 1 14
2 63871 1 14
2 63872 1 14
2 63873 1 14
2 63874 1 14
2 63875 1 14
2 63876 1 14
2 63877 1 14
2 63878 1 14
2 63879 1 14
2 63880 1 14
2 63881 1 14
2 63882 1 14
2 63883 1 14
2 63884 1 14
2 63885 1 14
2 63886 1 14
2 63887 1 14
2 63888 1 14
2 63889 1 14
2 63890 1 14
2 63891 1 14
2 63892 1 14
2 63893 1 14
2 63894 1 14
2 63895 1 14
2 63896 1 14
2 63897 1 14
2 63898 1 14
2 63899 1 14
2 63900 1 14
2 63901 1 14
2 63902 1 14
2 63903 1 14
2 63904 1 14
2 63905 1 14
2 63906 1 14
2 63907 1 14
2 63908 1 14
2 63909 1 14
2 63910 1 14
2 63911 1 14
2 63912 1 14
2 63913 1 14
2 63914 1 14
2 63915 1 14
2 63916 1 14
2 63917 1 14
2 63918 1 14
2 63919 1 14
2 63920 1 14
2 63921 1 14
2 63922 1 14
2 63923 1 14
2 63924 1 14
2 63925 1 14
2 63926 1 14
2 63927 1 14
2 63928 1 14
2 63929 1 14
2 63930 1 14
2 63931 1 14
2 63932 1 14
2 63933 1 14
2 63934 1 14
2 63935 1 14
2 63936 1 14
2 63937 1 14
2 63938 1 14
2 63939 1 14
2 63940 1 14
2 63941 1 14
2 63942 1 14
2 63943 1 14
2 63944 1 14
2 63945 1 14
2 63946 1 14
2 63947 1 14
2 63948 1 14
2 63949 1 14
2 63950 1 14
2 63951 1 14
2 63952 1 14
2 63953 1 14
2 63954 1 14
2 63955 1 14
2 63956 1 14
2 63957 1 14
2 63958 1 14
2 63959 1 14
2 63960 1 14
2 63961 1 14
2 63962 1 14
2 63963 1 14
2 63964 1 14
2 63965 1 14
2 63966 1 14
2 63967 1 14
2 63968 1 14
2 63969 1 14
2 63970 1 14
2 63971 1 14
2 63972 1 14
2 63973 1 14
2 63974 1 14
2 63975 1 14
2 63976 1 14
2 63977 1 14
2 63978 1 14
2 63979 1 14
2 63980 1 14
2 63981 1 14
2 63982 1 14
2 63983 1 14
2 63984 1 14
2 63985 1 14
2 63986 1 14
2 63987 1 14
2 63988 1 14
2 63989 1 14
2 63990 1 14
2 63991 1 14
2 63992 1 14
2 63993 1 14
2 63994 1 14
2 63995 1 14
2 63996 1 14
2 63997 1 14
2 63998 1 14
2 63999 1 14
2 64000 1 14
2 64001 1 14
2 64002 1 14
2 64003 1 14
2 64004 1 14
2 64005 1 14
2 64006 1 14
2 64007 1 14
2 64008 1 14
2 64009 1 14
2 64010 1 14
2 64011 1 14
2 64012 1 14
2 64013 1 14
2 64014 1 14
2 64015 1 14
2 64016 1 14
2 64017 1 14
1 15 0 222 0
2 64018 1 15
2 64019 1 15
2 64020 1 15
2 64021 1 15
2 64022 1 15
2 64023 1 15
2 64024 1 15
2 64025 1 15
2 64026 1 15
2 64027 1 15
2 64028 1 15
2 64029 1 15
2 64030 1 15
2 64031 1 15
2 64032 1 15
2 64033 1 15
2 64034 1 15
2 64035 1 15
2 64036 1 15
2 64037 1 15
2 64038 1 15
2 64039 1 15
2 64040 1 15
2 64041 1 15
2 64042 1 15
2 64043 1 15
2 64044 1 15
2 64045 1 15
2 64046 1 15
2 64047 1 15
2 64048 1 15
2 64049 1 15
2 64050 1 15
2 64051 1 15
2 64052 1 15
2 64053 1 15
2 64054 1 15
2 64055 1 15
2 64056 1 15
2 64057 1 15
2 64058 1 15
2 64059 1 15
2 64060 1 15
2 64061 1 15
2 64062 1 15
2 64063 1 15
2 64064 1 15
2 64065 1 15
2 64066 1 15
2 64067 1 15
2 64068 1 15
2 64069 1 15
2 64070 1 15
2 64071 1 15
2 64072 1 15
2 64073 1 15
2 64074 1 15
2 64075 1 15
2 64076 1 15
2 64077 1 15
2 64078 1 15
2 64079 1 15
2 64080 1 15
2 64081 1 15
2 64082 1 15
2 64083 1 15
2 64084 1 15
2 64085 1 15
2 64086 1 15
2 64087 1 15
2 64088 1 15
2 64089 1 15
2 64090 1 15
2 64091 1 15
2 64092 1 15
2 64093 1 15
2 64094 1 15
2 64095 1 15
2 64096 1 15
2 64097 1 15
2 64098 1 15
2 64099 1 15
2 64100 1 15
2 64101 1 15
2 64102 1 15
2 64103 1 15
2 64104 1 15
2 64105 1 15
2 64106 1 15
2 64107 1 15
2 64108 1 15
2 64109 1 15
2 64110 1 15
2 64111 1 15
2 64112 1 15
2 64113 1 15
2 64114 1 15
2 64115 1 15
2 64116 1 15
2 64117 1 15
2 64118 1 15
2 64119 1 15
2 64120 1 15
2 64121 1 15
2 64122 1 15
2 64123 1 15
2 64124 1 15
2 64125 1 15
2 64126 1 15
2 64127 1 15
2 64128 1 15
2 64129 1 15
2 64130 1 15
2 64131 1 15
2 64132 1 15
2 64133 1 15
2 64134 1 15
2 64135 1 15
2 64136 1 15
2 64137 1 15
2 64138 1 15
2 64139 1 15
2 64140 1 15
2 64141 1 15
2 64142 1 15
2 64143 1 15
2 64144 1 15
2 64145 1 15
2 64146 1 15
2 64147 1 15
2 64148 1 15
2 64149 1 15
2 64150 1 15
2 64151 1 15
2 64152 1 15
2 64153 1 15
2 64154 1 15
2 64155 1 15
2 64156 1 15
2 64157 1 15
2 64158 1 15
2 64159 1 15
2 64160 1 15
2 64161 1 15
2 64162 1 15
2 64163 1 15
2 64164 1 15
2 64165 1 15
2 64166 1 15
2 64167 1 15
2 64168 1 15
2 64169 1 15
2 64170 1 15
2 64171 1 15
2 64172 1 15
2 64173 1 15
2 64174 1 15
2 64175 1 15
2 64176 1 15
2 64177 1 15
2 64178 1 15
2 64179 1 15
2 64180 1 15
2 64181 1 15
2 64182 1 15
2 64183 1 15
2 64184 1 15
2 64185 1 15
2 64186 1 15
2 64187 1 15
2 64188 1 15
2 64189 1 15
2 64190 1 15
2 64191 1 15
2 64192 1 15
2 64193 1 15
2 64194 1 15
2 64195 1 15
2 64196 1 15
2 64197 1 15
2 64198 1 15
2 64199 1 15
2 64200 1 15
2 64201 1 15
2 64202 1 15
2 64203 1 15
2 64204 1 15
2 64205 1 15
2 64206 1 15
2 64207 1 15
2 64208 1 15
2 64209 1 15
2 64210 1 15
2 64211 1 15
2 64212 1 15
2 64213 1 15
2 64214 1 15
2 64215 1 15
2 64216 1 15
2 64217 1 15
2 64218 1 15
2 64219 1 15
2 64220 1 15
2 64221 1 15
2 64222 1 15
2 64223 1 15
2 64224 1 15
2 64225 1 15
2 64226 1 15
2 64227 1 15
2 64228 1 15
2 64229 1 15
2 64230 1 15
2 64231 1 15
2 64232 1 15
2 64233 1 15
2 64234 1 15
2 64235 1 15
2 64236 1 15
2 64237 1 15
2 64238 1 15
2 64239 1 15
1 16 0 71 0
2 64240 1 16
2 64241 1 16
2 64242 1 16
2 64243 1 16
2 64244 1 16
2 64245 1 16
2 64246 1 16
2 64247 1 16
2 64248 1 16
2 64249 1 16
2 64250 1 16
2 64251 1 16
2 64252 1 16
2 64253 1 16
2 64254 1 16
2 64255 1 16
2 64256 1 16
2 64257 1 16
2 64258 1 16
2 64259 1 16
2 64260 1 16
2 64261 1 16
2 64262 1 16
2 64263 1 16
2 64264 1 16
2 64265 1 16
2 64266 1 16
2 64267 1 16
2 64268 1 16
2 64269 1 16
2 64270 1 16
2 64271 1 16
2 64272 1 16
2 64273 1 16
2 64274 1 16
2 64275 1 16
2 64276 1 16
2 64277 1 16
2 64278 1 16
2 64279 1 16
2 64280 1 16
2 64281 1 16
2 64282 1 16
2 64283 1 16
2 64284 1 16
2 64285 1 16
2 64286 1 16
2 64287 1 16
2 64288 1 16
2 64289 1 16
2 64290 1 16
2 64291 1 16
2 64292 1 16
2 64293 1 16
2 64294 1 16
2 64295 1 16
2 64296 1 16
2 64297 1 16
2 64298 1 16
2 64299 1 16
2 64300 1 16
2 64301 1 16
2 64302 1 16
2 64303 1 16
2 64304 1 16
2 64305 1 16
2 64306 1 16
2 64307 1 16
2 64308 1 16
2 64309 1 16
2 64310 1 16
1 17 0 115 0
2 64311 1 17
2 64312 1 17
2 64313 1 17
2 64314 1 17
2 64315 1 17
2 64316 1 17
2 64317 1 17
2 64318 1 17
2 64319 1 17
2 64320 1 17
2 64321 1 17
2 64322 1 17
2 64323 1 17
2 64324 1 17
2 64325 1 17
2 64326 1 17
2 64327 1 17
2 64328 1 17
2 64329 1 17
2 64330 1 17
2 64331 1 17
2 64332 1 17
2 64333 1 17
2 64334 1 17
2 64335 1 17
2 64336 1 17
2 64337 1 17
2 64338 1 17
2 64339 1 17
2 64340 1 17
2 64341 1 17
2 64342 1 17
2 64343 1 17
2 64344 1 17
2 64345 1 17
2 64346 1 17
2 64347 1 17
2 64348 1 17
2 64349 1 17
2 64350 1 17
2 64351 1 17
2 64352 1 17
2 64353 1 17
2 64354 1 17
2 64355 1 17
2 64356 1 17
2 64357 1 17
2 64358 1 17
2 64359 1 17
2 64360 1 17
2 64361 1 17
2 64362 1 17
2 64363 1 17
2 64364 1 17
2 64365 1 17
2 64366 1 17
2 64367 1 17
2 64368 1 17
2 64369 1 17
2 64370 1 17
2 64371 1 17
2 64372 1 17
2 64373 1 17
2 64374 1 17
2 64375 1 17
2 64376 1 17
2 64377 1 17
2 64378 1 17
2 64379 1 17
2 64380 1 17
2 64381 1 17
2 64382 1 17
2 64383 1 17
2 64384 1 17
2 64385 1 17
2 64386 1 17
2 64387 1 17
2 64388 1 17
2 64389 1 17
2 64390 1 17
2 64391 1 17
2 64392 1 17
2 64393 1 17
2 64394 1 17
2 64395 1 17
2 64396 1 17
2 64397 1 17
2 64398 1 17
2 64399 1 17
2 64400 1 17
2 64401 1 17
2 64402 1 17
2 64403 1 17
2 64404 1 17
2 64405 1 17
2 64406 1 17
2 64407 1 17
2 64408 1 17
2 64409 1 17
2 64410 1 17
2 64411 1 17
2 64412 1 17
2 64413 1 17
2 64414 1 17
2 64415 1 17
2 64416 1 17
2 64417 1 17
2 64418 1 17
2 64419 1 17
2 64420 1 17
2 64421 1 17
2 64422 1 17
2 64423 1 17
2 64424 1 17
2 64425 1 17
1 18 0 183 0
2 64426 1 18
2 64427 1 18
2 64428 1 18
2 64429 1 18
2 64430 1 18
2 64431 1 18
2 64432 1 18
2 64433 1 18
2 64434 1 18
2 64435 1 18
2 64436 1 18
2 64437 1 18
2 64438 1 18
2 64439 1 18
2 64440 1 18
2 64441 1 18
2 64442 1 18
2 64443 1 18
2 64444 1 18
2 64445 1 18
2 64446 1 18
2 64447 1 18
2 64448 1 18
2 64449 1 18
2 64450 1 18
2 64451 1 18
2 64452 1 18
2 64453 1 18
2 64454 1 18
2 64455 1 18
2 64456 1 18
2 64457 1 18
2 64458 1 18
2 64459 1 18
2 64460 1 18
2 64461 1 18
2 64462 1 18
2 64463 1 18
2 64464 1 18
2 64465 1 18
2 64466 1 18
2 64467 1 18
2 64468 1 18
2 64469 1 18
2 64470 1 18
2 64471 1 18
2 64472 1 18
2 64473 1 18
2 64474 1 18
2 64475 1 18
2 64476 1 18
2 64477 1 18
2 64478 1 18
2 64479 1 18
2 64480 1 18
2 64481 1 18
2 64482 1 18
2 64483 1 18
2 64484 1 18
2 64485 1 18
2 64486 1 18
2 64487 1 18
2 64488 1 18
2 64489 1 18
2 64490 1 18
2 64491 1 18
2 64492 1 18
2 64493 1 18
2 64494 1 18
2 64495 1 18
2 64496 1 18
2 64497 1 18
2 64498 1 18
2 64499 1 18
2 64500 1 18
2 64501 1 18
2 64502 1 18
2 64503 1 18
2 64504 1 18
2 64505 1 18
2 64506 1 18
2 64507 1 18
2 64508 1 18
2 64509 1 18
2 64510 1 18
2 64511 1 18
2 64512 1 18
2 64513 1 18
2 64514 1 18
2 64515 1 18
2 64516 1 18
2 64517 1 18
2 64518 1 18
2 64519 1 18
2 64520 1 18
2 64521 1 18
2 64522 1 18
2 64523 1 18
2 64524 1 18
2 64525 1 18
2 64526 1 18
2 64527 1 18
2 64528 1 18
2 64529 1 18
2 64530 1 18
2 64531 1 18
2 64532 1 18
2 64533 1 18
2 64534 1 18
2 64535 1 18
2 64536 1 18
2 64537 1 18
2 64538 1 18
2 64539 1 18
2 64540 1 18
2 64541 1 18
2 64542 1 18
2 64543 1 18
2 64544 1 18
2 64545 1 18
2 64546 1 18
2 64547 1 18
2 64548 1 18
2 64549 1 18
2 64550 1 18
2 64551 1 18
2 64552 1 18
2 64553 1 18
2 64554 1 18
2 64555 1 18
2 64556 1 18
2 64557 1 18
2 64558 1 18
2 64559 1 18
2 64560 1 18
2 64561 1 18
2 64562 1 18
2 64563 1 18
2 64564 1 18
2 64565 1 18
2 64566 1 18
2 64567 1 18
2 64568 1 18
2 64569 1 18
2 64570 1 18
2 64571 1 18
2 64572 1 18
2 64573 1 18
2 64574 1 18
2 64575 1 18
2 64576 1 18
2 64577 1 18
2 64578 1 18
2 64579 1 18
2 64580 1 18
2 64581 1 18
2 64582 1 18
2 64583 1 18
2 64584 1 18
2 64585 1 18
2 64586 1 18
2 64587 1 18
2 64588 1 18
2 64589 1 18
2 64590 1 18
2 64591 1 18
2 64592 1 18
2 64593 1 18
2 64594 1 18
2 64595 1 18
2 64596 1 18
2 64597 1 18
2 64598 1 18
2 64599 1 18
2 64600 1 18
2 64601 1 18
2 64602 1 18
2 64603 1 18
2 64604 1 18
2 64605 1 18
2 64606 1 18
2 64607 1 18
2 64608 1 18
1 19 0 210 0
2 64609 1 19
2 64610 1 19
2 64611 1 19
2 64612 1 19
2 64613 1 19
2 64614 1 19
2 64615 1 19
2 64616 1 19
2 64617 1 19
2 64618 1 19
2 64619 1 19
2 64620 1 19
2 64621 1 19
2 64622 1 19
2 64623 1 19
2 64624 1 19
2 64625 1 19
2 64626 1 19
2 64627 1 19
2 64628 1 19
2 64629 1 19
2 64630 1 19
2 64631 1 19
2 64632 1 19
2 64633 1 19
2 64634 1 19
2 64635 1 19
2 64636 1 19
2 64637 1 19
2 64638 1 19
2 64639 1 19
2 64640 1 19
2 64641 1 19
2 64642 1 19
2 64643 1 19
2 64644 1 19
2 64645 1 19
2 64646 1 19
2 64647 1 19
2 64648 1 19
2 64649 1 19
2 64650 1 19
2 64651 1 19
2 64652 1 19
2 64653 1 19
2 64654 1 19
2 64655 1 19
2 64656 1 19
2 64657 1 19
2 64658 1 19
2 64659 1 19
2 64660 1 19
2 64661 1 19
2 64662 1 19
2 64663 1 19
2 64664 1 19
2 64665 1 19
2 64666 1 19
2 64667 1 19
2 64668 1 19
2 64669 1 19
2 64670 1 19
2 64671 1 19
2 64672 1 19
2 64673 1 19
2 64674 1 19
2 64675 1 19
2 64676 1 19
2 64677 1 19
2 64678 1 19
2 64679 1 19
2 64680 1 19
2 64681 1 19
2 64682 1 19
2 64683 1 19
2 64684 1 19
2 64685 1 19
2 64686 1 19
2 64687 1 19
2 64688 1 19
2 64689 1 19
2 64690 1 19
2 64691 1 19
2 64692 1 19
2 64693 1 19
2 64694 1 19
2 64695 1 19
2 64696 1 19
2 64697 1 19
2 64698 1 19
2 64699 1 19
2 64700 1 19
2 64701 1 19
2 64702 1 19
2 64703 1 19
2 64704 1 19
2 64705 1 19
2 64706 1 19
2 64707 1 19
2 64708 1 19
2 64709 1 19
2 64710 1 19
2 64711 1 19
2 64712 1 19
2 64713 1 19
2 64714 1 19
2 64715 1 19
2 64716 1 19
2 64717 1 19
2 64718 1 19
2 64719 1 19
2 64720 1 19
2 64721 1 19
2 64722 1 19
2 64723 1 19
2 64724 1 19
2 64725 1 19
2 64726 1 19
2 64727 1 19
2 64728 1 19
2 64729 1 19
2 64730 1 19
2 64731 1 19
2 64732 1 19
2 64733 1 19
2 64734 1 19
2 64735 1 19
2 64736 1 19
2 64737 1 19
2 64738 1 19
2 64739 1 19
2 64740 1 19
2 64741 1 19
2 64742 1 19
2 64743 1 19
2 64744 1 19
2 64745 1 19
2 64746 1 19
2 64747 1 19
2 64748 1 19
2 64749 1 19
2 64750 1 19
2 64751 1 19
2 64752 1 19
2 64753 1 19
2 64754 1 19
2 64755 1 19
2 64756 1 19
2 64757 1 19
2 64758 1 19
2 64759 1 19
2 64760 1 19
2 64761 1 19
2 64762 1 19
2 64763 1 19
2 64764 1 19
2 64765 1 19
2 64766 1 19
2 64767 1 19
2 64768 1 19
2 64769 1 19
2 64770 1 19
2 64771 1 19
2 64772 1 19
2 64773 1 19
2 64774 1 19
2 64775 1 19
2 64776 1 19
2 64777 1 19
2 64778 1 19
2 64779 1 19
2 64780 1 19
2 64781 1 19
2 64782 1 19
2 64783 1 19
2 64784 1 19
2 64785 1 19
2 64786 1 19
2 64787 1 19
2 64788 1 19
2 64789 1 19
2 64790 1 19
2 64791 1 19
2 64792 1 19
2 64793 1 19
2 64794 1 19
2 64795 1 19
2 64796 1 19
2 64797 1 19
2 64798 1 19
2 64799 1 19
2 64800 1 19
2 64801 1 19
2 64802 1 19
2 64803 1 19
2 64804 1 19
2 64805 1 19
2 64806 1 19
2 64807 1 19
2 64808 1 19
2 64809 1 19
2 64810 1 19
2 64811 1 19
2 64812 1 19
2 64813 1 19
2 64814 1 19
2 64815 1 19
2 64816 1 19
2 64817 1 19
2 64818 1 19
1 20 0 189 0
2 64819 1 20
2 64820 1 20
2 64821 1 20
2 64822 1 20
2 64823 1 20
2 64824 1 20
2 64825 1 20
2 64826 1 20
2 64827 1 20
2 64828 1 20
2 64829 1 20
2 64830 1 20
2 64831 1 20
2 64832 1 20
2 64833 1 20
2 64834 1 20
2 64835 1 20
2 64836 1 20
2 64837 1 20
2 64838 1 20
2 64839 1 20
2 64840 1 20
2 64841 1 20
2 64842 1 20
2 64843 1 20
2 64844 1 20
2 64845 1 20
2 64846 1 20
2 64847 1 20
2 64848 1 20
2 64849 1 20
2 64850 1 20
2 64851 1 20
2 64852 1 20
2 64853 1 20
2 64854 1 20
2 64855 1 20
2 64856 1 20
2 64857 1 20
2 64858 1 20
2 64859 1 20
2 64860 1 20
2 64861 1 20
2 64862 1 20
2 64863 1 20
2 64864 1 20
2 64865 1 20
2 64866 1 20
2 64867 1 20
2 64868 1 20
2 64869 1 20
2 64870 1 20
2 64871 1 20
2 64872 1 20
2 64873 1 20
2 64874 1 20
2 64875 1 20
2 64876 1 20
2 64877 1 20
2 64878 1 20
2 64879 1 20
2 64880 1 20
2 64881 1 20
2 64882 1 20
2 64883 1 20
2 64884 1 20
2 64885 1 20
2 64886 1 20
2 64887 1 20
2 64888 1 20
2 64889 1 20
2 64890 1 20
2 64891 1 20
2 64892 1 20
2 64893 1 20
2 64894 1 20
2 64895 1 20
2 64896 1 20
2 64897 1 20
2 64898 1 20
2 64899 1 20
2 64900 1 20
2 64901 1 20
2 64902 1 20
2 64903 1 20
2 64904 1 20
2 64905 1 20
2 64906 1 20
2 64907 1 20
2 64908 1 20
2 64909 1 20
2 64910 1 20
2 64911 1 20
2 64912 1 20
2 64913 1 20
2 64914 1 20
2 64915 1 20
2 64916 1 20
2 64917 1 20
2 64918 1 20
2 64919 1 20
2 64920 1 20
2 64921 1 20
2 64922 1 20
2 64923 1 20
2 64924 1 20
2 64925 1 20
2 64926 1 20
2 64927 1 20
2 64928 1 20
2 64929 1 20
2 64930 1 20
2 64931 1 20
2 64932 1 20
2 64933 1 20
2 64934 1 20
2 64935 1 20
2 64936 1 20
2 64937 1 20
2 64938 1 20
2 64939 1 20
2 64940 1 20
2 64941 1 20
2 64942 1 20
2 64943 1 20
2 64944 1 20
2 64945 1 20
2 64946 1 20
2 64947 1 20
2 64948 1 20
2 64949 1 20
2 64950 1 20
2 64951 1 20
2 64952 1 20
2 64953 1 20
2 64954 1 20
2 64955 1 20
2 64956 1 20
2 64957 1 20
2 64958 1 20
2 64959 1 20
2 64960 1 20
2 64961 1 20
2 64962 1 20
2 64963 1 20
2 64964 1 20
2 64965 1 20
2 64966 1 20
2 64967 1 20
2 64968 1 20
2 64969 1 20
2 64970 1 20
2 64971 1 20
2 64972 1 20
2 64973 1 20
2 64974 1 20
2 64975 1 20
2 64976 1 20
2 64977 1 20
2 64978 1 20
2 64979 1 20
2 64980 1 20
2 64981 1 20
2 64982 1 20
2 64983 1 20
2 64984 1 20
2 64985 1 20
2 64986 1 20
2 64987 1 20
2 64988 1 20
2 64989 1 20
2 64990 1 20
2 64991 1 20
2 64992 1 20
2 64993 1 20
2 64994 1 20
2 64995 1 20
2 64996 1 20
2 64997 1 20
2 64998 1 20
2 64999 1 20
2 65000 1 20
2 65001 1 20
2 65002 1 20
2 65003 1 20
2 65004 1 20
2 65005 1 20
2 65006 1 20
2 65007 1 20
1 21 0 256 0
2 65008 1 21
2 65009 1 21
2 65010 1 21
2 65011 1 21
2 65012 1 21
2 65013 1 21
2 65014 1 21
2 65015 1 21
2 65016 1 21
2 65017 1 21
2 65018 1 21
2 65019 1 21
2 65020 1 21
2 65021 1 21
2 65022 1 21
2 65023 1 21
2 65024 1 21
2 65025 1 21
2 65026 1 21
2 65027 1 21
2 65028 1 21
2 65029 1 21
2 65030 1 21
2 65031 1 21
2 65032 1 21
2 65033 1 21
2 65034 1 21
2 65035 1 21
2 65036 1 21
2 65037 1 21
2 65038 1 21
2 65039 1 21
2 65040 1 21
2 65041 1 21
2 65042 1 21
2 65043 1 21
2 65044 1 21
2 65045 1 21
2 65046 1 21
2 65047 1 21
2 65048 1 21
2 65049 1 21
2 65050 1 21
2 65051 1 21
2 65052 1 21
2 65053 1 21
2 65054 1 21
2 65055 1 21
2 65056 1 21
2 65057 1 21
2 65058 1 21
2 65059 1 21
2 65060 1 21
2 65061 1 21
2 65062 1 21
2 65063 1 21
2 65064 1 21
2 65065 1 21
2 65066 1 21
2 65067 1 21
2 65068 1 21
2 65069 1 21
2 65070 1 21
2 65071 1 21
2 65072 1 21
2 65073 1 21
2 65074 1 21
2 65075 1 21
2 65076 1 21
2 65077 1 21
2 65078 1 21
2 65079 1 21
2 65080 1 21
2 65081 1 21
2 65082 1 21
2 65083 1 21
2 65084 1 21
2 65085 1 21
2 65086 1 21
2 65087 1 21
2 65088 1 21
2 65089 1 21
2 65090 1 21
2 65091 1 21
2 65092 1 21
2 65093 1 21
2 65094 1 21
2 65095 1 21
2 65096 1 21
2 65097 1 21
2 65098 1 21
2 65099 1 21
2 65100 1 21
2 65101 1 21
2 65102 1 21
2 65103 1 21
2 65104 1 21
2 65105 1 21
2 65106 1 21
2 65107 1 21
2 65108 1 21
2 65109 1 21
2 65110 1 21
2 65111 1 21
2 65112 1 21
2 65113 1 21
2 65114 1 21
2 65115 1 21
2 65116 1 21
2 65117 1 21
2 65118 1 21
2 65119 1 21
2 65120 1 21
2 65121 1 21
2 65122 1 21
2 65123 1 21
2 65124 1 21
2 65125 1 21
2 65126 1 21
2 65127 1 21
2 65128 1 21
2 65129 1 21
2 65130 1 21
2 65131 1 21
2 65132 1 21
2 65133 1 21
2 65134 1 21
2 65135 1 21
2 65136 1 21
2 65137 1 21
2 65138 1 21
2 65139 1 21
2 65140 1 21
2 65141 1 21
2 65142 1 21
2 65143 1 21
2 65144 1 21
2 65145 1 21
2 65146 1 21
2 65147 1 21
2 65148 1 21
2 65149 1 21
2 65150 1 21
2 65151 1 21
2 65152 1 21
2 65153 1 21
2 65154 1 21
2 65155 1 21
2 65156 1 21
2 65157 1 21
2 65158 1 21
2 65159 1 21
2 65160 1 21
2 65161 1 21
2 65162 1 21
2 65163 1 21
2 65164 1 21
2 65165 1 21
2 65166 1 21
2 65167 1 21
2 65168 1 21
2 65169 1 21
2 65170 1 21
2 65171 1 21
2 65172 1 21
2 65173 1 21
2 65174 1 21
2 65175 1 21
2 65176 1 21
2 65177 1 21
2 65178 1 21
2 65179 1 21
2 65180 1 21
2 65181 1 21
2 65182 1 21
2 65183 1 21
2 65184 1 21
2 65185 1 21
2 65186 1 21
2 65187 1 21
2 65188 1 21
2 65189 1 21
2 65190 1 21
2 65191 1 21
2 65192 1 21
2 65193 1 21
2 65194 1 21
2 65195 1 21
2 65196 1 21
2 65197 1 21
2 65198 1 21
2 65199 1 21
2 65200 1 21
2 65201 1 21
2 65202 1 21
2 65203 1 21
2 65204 1 21
2 65205 1 21
2 65206 1 21
2 65207 1 21
2 65208 1 21
2 65209 1 21
2 65210 1 21
2 65211 1 21
2 65212 1 21
2 65213 1 21
2 65214 1 21
2 65215 1 21
2 65216 1 21
2 65217 1 21
2 65218 1 21
2 65219 1 21
2 65220 1 21
2 65221 1 21
2 65222 1 21
2 65223 1 21
2 65224 1 21
2 65225 1 21
2 65226 1 21
2 65227 1 21
2 65228 1 21
2 65229 1 21
2 65230 1 21
2 65231 1 21
2 65232 1 21
2 65233 1 21
2 65234 1 21
2 65235 1 21
2 65236 1 21
2 65237 1 21
2 65238 1 21
2 65239 1 21
2 65240 1 21
2 65241 1 21
2 65242 1 21
2 65243 1 21
2 65244 1 21
2 65245 1 21
2 65246 1 21
2 65247 1 21
2 65248 1 21
2 65249 1 21
2 65250 1 21
2 65251 1 21
2 65252 1 21
2 65253 1 21
2 65254 1 21
2 65255 1 21
2 65256 1 21
2 65257 1 21
2 65258 1 21
2 65259 1 21
2 65260 1 21
2 65261 1 21
2 65262 1 21
2 65263 1 21
1 22 0 356 0
2 65264 1 22
2 65265 1 22
2 65266 1 22
2 65267 1 22
2 65268 1 22
2 65269 1 22
2 65270 1 22
2 65271 1 22
2 65272 1 22
2 65273 1 22
2 65274 1 22
2 65275 1 22
2 65276 1 22
2 65277 1 22
2 65278 1 22
2 65279 1 22
2 65280 1 22
2 65281 1 22
2 65282 1 22
2 65283 1 22
2 65284 1 22
2 65285 1 22
2 65286 1 22
2 65287 1 22
2 65288 1 22
2 65289 1 22
2 65290 1 22
2 65291 1 22
2 65292 1 22
2 65293 1 22
2 65294 1 22
2 65295 1 22
2 65296 1 22
2 65297 1 22
2 65298 1 22
2 65299 1 22
2 65300 1 22
2 65301 1 22
2 65302 1 22
2 65303 1 22
2 65304 1 22
2 65305 1 22
2 65306 1 22
2 65307 1 22
2 65308 1 22
2 65309 1 22
2 65310 1 22
2 65311 1 22
2 65312 1 22
2 65313 1 22
2 65314 1 22
2 65315 1 22
2 65316 1 22
2 65317 1 22
2 65318 1 22
2 65319 1 22
2 65320 1 22
2 65321 1 22
2 65322 1 22
2 65323 1 22
2 65324 1 22
2 65325 1 22
2 65326 1 22
2 65327 1 22
2 65328 1 22
2 65329 1 22
2 65330 1 22
2 65331 1 22
2 65332 1 22
2 65333 1 22
2 65334 1 22
2 65335 1 22
2 65336 1 22
2 65337 1 22
2 65338 1 22
2 65339 1 22
2 65340 1 22
2 65341 1 22
2 65342 1 22
2 65343 1 22
2 65344 1 22
2 65345 1 22
2 65346 1 22
2 65347 1 22
2 65348 1 22
2 65349 1 22
2 65350 1 22
2 65351 1 22
2 65352 1 22
2 65353 1 22
2 65354 1 22
2 65355 1 22
2 65356 1 22
2 65357 1 22
2 65358 1 22
2 65359 1 22
2 65360 1 22
2 65361 1 22
2 65362 1 22
2 65363 1 22
2 65364 1 22
2 65365 1 22
2 65366 1 22
2 65367 1 22
2 65368 1 22
2 65369 1 22
2 65370 1 22
2 65371 1 22
2 65372 1 22
2 65373 1 22
2 65374 1 22
2 65375 1 22
2 65376 1 22
2 65377 1 22
2 65378 1 22
2 65379 1 22
2 65380 1 22
2 65381 1 22
2 65382 1 22
2 65383 1 22
2 65384 1 22
2 65385 1 22
2 65386 1 22
2 65387 1 22
2 65388 1 22
2 65389 1 22
2 65390 1 22
2 65391 1 22
2 65392 1 22
2 65393 1 22
2 65394 1 22
2 65395 1 22
2 65396 1 22
2 65397 1 22
2 65398 1 22
2 65399 1 22
2 65400 1 22
2 65401 1 22
2 65402 1 22
2 65403 1 22
2 65404 1 22
2 65405 1 22
2 65406 1 22
2 65407 1 22
2 65408 1 22
2 65409 1 22
2 65410 1 22
2 65411 1 22
2 65412 1 22
2 65413 1 22
2 65414 1 22
2 65415 1 22
2 65416 1 22
2 65417 1 22
2 65418 1 22
2 65419 1 22
2 65420 1 22
2 65421 1 22
2 65422 1 22
2 65423 1 22
2 65424 1 22
2 65425 1 22
2 65426 1 22
2 65427 1 22
2 65428 1 22
2 65429 1 22
2 65430 1 22
2 65431 1 22
2 65432 1 22
2 65433 1 22
2 65434 1 22
2 65435 1 22
2 65436 1 22
2 65437 1 22
2 65438 1 22
2 65439 1 22
2 65440 1 22
2 65441 1 22
2 65442 1 22
2 65443 1 22
2 65444 1 22
2 65445 1 22
2 65446 1 22
2 65447 1 22
2 65448 1 22
2 65449 1 22
2 65450 1 22
2 65451 1 22
2 65452 1 22
2 65453 1 22
2 65454 1 22
2 65455 1 22
2 65456 1 22
2 65457 1 22
2 65458 1 22
2 65459 1 22
2 65460 1 22
2 65461 1 22
2 65462 1 22
2 65463 1 22
2 65464 1 22
2 65465 1 22
2 65466 1 22
2 65467 1 22
2 65468 1 22
2 65469 1 22
2 65470 1 22
2 65471 1 22
2 65472 1 22
2 65473 1 22
2 65474 1 22
2 65475 1 22
2 65476 1 22
2 65477 1 22
2 65478 1 22
2 65479 1 22
2 65480 1 22
2 65481 1 22
2 65482 1 22
2 65483 1 22
2 65484 1 22
2 65485 1 22
2 65486 1 22
2 65487 1 22
2 65488 1 22
2 65489 1 22
2 65490 1 22
2 65491 1 22
2 65492 1 22
2 65493 1 22
2 65494 1 22
2 65495 1 22
2 65496 1 22
2 65497 1 22
2 65498 1 22
2 65499 1 22
2 65500 1 22
2 65501 1 22
2 65502 1 22
2 65503 1 22
2 65504 1 22
2 65505 1 22
2 65506 1 22
2 65507 1 22
2 65508 1 22
2 65509 1 22
2 65510 1 22
2 65511 1 22
2 65512 1 22
2 65513 1 22
2 65514 1 22
2 65515 1 22
2 65516 1 22
2 65517 1 22
2 65518 1 22
2 65519 1 22
2 65520 1 22
2 65521 1 22
2 65522 1 22
2 65523 1 22
2 65524 1 22
2 65525 1 22
2 65526 1 22
2 65527 1 22
2 65528 1 22
2 65529 1 22
2 65530 1 22
2 65531 1 22
2 65532 1 22
2 65533 1 22
2 65534 1 22
2 65535 1 22
2 65536 1 22
2 65537 1 22
2 65538 1 22
2 65539 1 22
2 65540 1 22
2 65541 1 22
2 65542 1 22
2 65543 1 22
2 65544 1 22
2 65545 1 22
2 65546 1 22
2 65547 1 22
2 65548 1 22
2 65549 1 22
2 65550 1 22
2 65551 1 22
2 65552 1 22
2 65553 1 22
2 65554 1 22
2 65555 1 22
2 65556 1 22
2 65557 1 22
2 65558 1 22
2 65559 1 22
2 65560 1 22
2 65561 1 22
2 65562 1 22
2 65563 1 22
2 65564 1 22
2 65565 1 22
2 65566 1 22
2 65567 1 22
2 65568 1 22
2 65569 1 22
2 65570 1 22
2 65571 1 22
2 65572 1 22
2 65573 1 22
2 65574 1 22
2 65575 1 22
2 65576 1 22
2 65577 1 22
2 65578 1 22
2 65579 1 22
2 65580 1 22
2 65581 1 22
2 65582 1 22
2 65583 1 22
2 65584 1 22
2 65585 1 22
2 65586 1 22
2 65587 1 22
2 65588 1 22
2 65589 1 22
2 65590 1 22
2 65591 1 22
2 65592 1 22
2 65593 1 22
2 65594 1 22
2 65595 1 22
2 65596 1 22
2 65597 1 22
2 65598 1 22
2 65599 1 22
2 65600 1 22
2 65601 1 22
2 65602 1 22
2 65603 1 22
2 65604 1 22
2 65605 1 22
2 65606 1 22
2 65607 1 22
2 65608 1 22
2 65609 1 22
2 65610 1 22
2 65611 1 22
2 65612 1 22
2 65613 1 22
2 65614 1 22
2 65615 1 22
2 65616 1 22
2 65617 1 22
2 65618 1 22
2 65619 1 22
1 23 0 273 0
2 65620 1 23
2 65621 1 23
2 65622 1 23
2 65623 1 23
2 65624 1 23
2 65625 1 23
2 65626 1 23
2 65627 1 23
2 65628 1 23
2 65629 1 23
2 65630 1 23
2 65631 1 23
2 65632 1 23
2 65633 1 23
2 65634 1 23
2 65635 1 23
2 65636 1 23
2 65637 1 23
2 65638 1 23
2 65639 1 23
2 65640 1 23
2 65641 1 23
2 65642 1 23
2 65643 1 23
2 65644 1 23
2 65645 1 23
2 65646 1 23
2 65647 1 23
2 65648 1 23
2 65649 1 23
2 65650 1 23
2 65651 1 23
2 65652 1 23
2 65653 1 23
2 65654 1 23
2 65655 1 23
2 65656 1 23
2 65657 1 23
2 65658 1 23
2 65659 1 23
2 65660 1 23
2 65661 1 23
2 65662 1 23
2 65663 1 23
2 65664 1 23
2 65665 1 23
2 65666 1 23
2 65667 1 23
2 65668 1 23
2 65669 1 23
2 65670 1 23
2 65671 1 23
2 65672 1 23
2 65673 1 23
2 65674 1 23
2 65675 1 23
2 65676 1 23
2 65677 1 23
2 65678 1 23
2 65679 1 23
2 65680 1 23
2 65681 1 23
2 65682 1 23
2 65683 1 23
2 65684 1 23
2 65685 1 23
2 65686 1 23
2 65687 1 23
2 65688 1 23
2 65689 1 23
2 65690 1 23
2 65691 1 23
2 65692 1 23
2 65693 1 23
2 65694 1 23
2 65695 1 23
2 65696 1 23
2 65697 1 23
2 65698 1 23
2 65699 1 23
2 65700 1 23
2 65701 1 23
2 65702 1 23
2 65703 1 23
2 65704 1 23
2 65705 1 23
2 65706 1 23
2 65707 1 23
2 65708 1 23
2 65709 1 23
2 65710 1 23
2 65711 1 23
2 65712 1 23
2 65713 1 23
2 65714 1 23
2 65715 1 23
2 65716 1 23
2 65717 1 23
2 65718 1 23
2 65719 1 23
2 65720 1 23
2 65721 1 23
2 65722 1 23
2 65723 1 23
2 65724 1 23
2 65725 1 23
2 65726 1 23
2 65727 1 23
2 65728 1 23
2 65729 1 23
2 65730 1 23
2 65731 1 23
2 65732 1 23
2 65733 1 23
2 65734 1 23
2 65735 1 23
2 65736 1 23
2 65737 1 23
2 65738 1 23
2 65739 1 23
2 65740 1 23
2 65741 1 23
2 65742 1 23
2 65743 1 23
2 65744 1 23
2 65745 1 23
2 65746 1 23
2 65747 1 23
2 65748 1 23
2 65749 1 23
2 65750 1 23
2 65751 1 23
2 65752 1 23
2 65753 1 23
2 65754 1 23
2 65755 1 23
2 65756 1 23
2 65757 1 23
2 65758 1 23
2 65759 1 23
2 65760 1 23
2 65761 1 23
2 65762 1 23
2 65763 1 23
2 65764 1 23
2 65765 1 23
2 65766 1 23
2 65767 1 23
2 65768 1 23
2 65769 1 23
2 65770 1 23
2 65771 1 23
2 65772 1 23
2 65773 1 23
2 65774 1 23
2 65775 1 23
2 65776 1 23
2 65777 1 23
2 65778 1 23
2 65779 1 23
2 65780 1 23
2 65781 1 23
2 65782 1 23
2 65783 1 23
2 65784 1 23
2 65785 1 23
2 65786 1 23
2 65787 1 23
2 65788 1 23
2 65789 1 23
2 65790 1 23
2 65791 1 23
2 65792 1 23
2 65793 1 23
2 65794 1 23
2 65795 1 23
2 65796 1 23
2 65797 1 23
2 65798 1 23
2 65799 1 23
2 65800 1 23
2 65801 1 23
2 65802 1 23
2 65803 1 23
2 65804 1 23
2 65805 1 23
2 65806 1 23
2 65807 1 23
2 65808 1 23
2 65809 1 23
2 65810 1 23
2 65811 1 23
2 65812 1 23
2 65813 1 23
2 65814 1 23
2 65815 1 23
2 65816 1 23
2 65817 1 23
2 65818 1 23
2 65819 1 23
2 65820 1 23
2 65821 1 23
2 65822 1 23
2 65823 1 23
2 65824 1 23
2 65825 1 23
2 65826 1 23
2 65827 1 23
2 65828 1 23
2 65829 1 23
2 65830 1 23
2 65831 1 23
2 65832 1 23
2 65833 1 23
2 65834 1 23
2 65835 1 23
2 65836 1 23
2 65837 1 23
2 65838 1 23
2 65839 1 23
2 65840 1 23
2 65841 1 23
2 65842 1 23
2 65843 1 23
2 65844 1 23
2 65845 1 23
2 65846 1 23
2 65847 1 23
2 65848 1 23
2 65849 1 23
2 65850 1 23
2 65851 1 23
2 65852 1 23
2 65853 1 23
2 65854 1 23
2 65855 1 23
2 65856 1 23
2 65857 1 23
2 65858 1 23
2 65859 1 23
2 65860 1 23
2 65861 1 23
2 65862 1 23
2 65863 1 23
2 65864 1 23
2 65865 1 23
2 65866 1 23
2 65867 1 23
2 65868 1 23
2 65869 1 23
2 65870 1 23
2 65871 1 23
2 65872 1 23
2 65873 1 23
2 65874 1 23
2 65875 1 23
2 65876 1 23
2 65877 1 23
2 65878 1 23
2 65879 1 23
2 65880 1 23
2 65881 1 23
2 65882 1 23
2 65883 1 23
2 65884 1 23
2 65885 1 23
2 65886 1 23
2 65887 1 23
2 65888 1 23
2 65889 1 23
2 65890 1 23
2 65891 1 23
2 65892 1 23
1 24 0 176 0
2 65893 1 24
2 65894 1 24
2 65895 1 24
2 65896 1 24
2 65897 1 24
2 65898 1 24
2 65899 1 24
2 65900 1 24
2 65901 1 24
2 65902 1 24
2 65903 1 24
2 65904 1 24
2 65905 1 24
2 65906 1 24
2 65907 1 24
2 65908 1 24
2 65909 1 24
2 65910 1 24
2 65911 1 24
2 65912 1 24
2 65913 1 24
2 65914 1 24
2 65915 1 24
2 65916 1 24
2 65917 1 24
2 65918 1 24
2 65919 1 24
2 65920 1 24
2 65921 1 24
2 65922 1 24
2 65923 1 24
2 65924 1 24
2 65925 1 24
2 65926 1 24
2 65927 1 24
2 65928 1 24
2 65929 1 24
2 65930 1 24
2 65931 1 24
2 65932 1 24
2 65933 1 24
2 65934 1 24
2 65935 1 24
2 65936 1 24
2 65937 1 24
2 65938 1 24
2 65939 1 24
2 65940 1 24
2 65941 1 24
2 65942 1 24
2 65943 1 24
2 65944 1 24
2 65945 1 24
2 65946 1 24
2 65947 1 24
2 65948 1 24
2 65949 1 24
2 65950 1 24
2 65951 1 24
2 65952 1 24
2 65953 1 24
2 65954 1 24
2 65955 1 24
2 65956 1 24
2 65957 1 24
2 65958 1 24
2 65959 1 24
2 65960 1 24
2 65961 1 24
2 65962 1 24
2 65963 1 24
2 65964 1 24
2 65965 1 24
2 65966 1 24
2 65967 1 24
2 65968 1 24
2 65969 1 24
2 65970 1 24
2 65971 1 24
2 65972 1 24
2 65973 1 24
2 65974 1 24
2 65975 1 24
2 65976 1 24
2 65977 1 24
2 65978 1 24
2 65979 1 24
2 65980 1 24
2 65981 1 24
2 65982 1 24
2 65983 1 24
2 65984 1 24
2 65985 1 24
2 65986 1 24
2 65987 1 24
2 65988 1 24
2 65989 1 24
2 65990 1 24
2 65991 1 24
2 65992 1 24
2 65993 1 24
2 65994 1 24
2 65995 1 24
2 65996 1 24
2 65997 1 24
2 65998 1 24
2 65999 1 24
2 66000 1 24
2 66001 1 24
2 66002 1 24
2 66003 1 24
2 66004 1 24
2 66005 1 24
2 66006 1 24
2 66007 1 24
2 66008 1 24
2 66009 1 24
2 66010 1 24
2 66011 1 24
2 66012 1 24
2 66013 1 24
2 66014 1 24
2 66015 1 24
2 66016 1 24
2 66017 1 24
2 66018 1 24
2 66019 1 24
2 66020 1 24
2 66021 1 24
2 66022 1 24
2 66023 1 24
2 66024 1 24
2 66025 1 24
2 66026 1 24
2 66027 1 24
2 66028 1 24
2 66029 1 24
2 66030 1 24
2 66031 1 24
2 66032 1 24
2 66033 1 24
2 66034 1 24
2 66035 1 24
2 66036 1 24
2 66037 1 24
2 66038 1 24
2 66039 1 24
2 66040 1 24
2 66041 1 24
2 66042 1 24
2 66043 1 24
2 66044 1 24
2 66045 1 24
2 66046 1 24
2 66047 1 24
2 66048 1 24
2 66049 1 24
2 66050 1 24
2 66051 1 24
2 66052 1 24
2 66053 1 24
2 66054 1 24
2 66055 1 24
2 66056 1 24
2 66057 1 24
2 66058 1 24
2 66059 1 24
2 66060 1 24
2 66061 1 24
2 66062 1 24
2 66063 1 24
2 66064 1 24
2 66065 1 24
2 66066 1 24
2 66067 1 24
2 66068 1 24
2 66069 1 27
2 66070 1 27
2 66071 1 27
2 66072 1 27
2 66073 1 27
2 66074 1 27
2 66075 1 27
2 66076 1 27
2 66077 1 27
2 66078 1 27
2 66079 1 27
2 66080 1 27
2 66081 1 27
2 66082 1 27
2 66083 1 27
2 66084 1 27
2 66085 1 27
2 66086 1 27
2 66087 1 27
2 66088 1 27
2 66089 1 27
2 66090 1 27
2 66091 1 27
2 66092 1 27
2 66093 1 27
2 66094 1 27
2 66095 1 27
2 66096 1 27
2 66097 1 27
2 66098 1 27
2 66099 1 27
2 66100 1 27
2 66101 1 27
2 66102 1 27
2 66103 1 27
2 66104 1 27
2 66105 1 27
2 66106 1 27
2 66107 1 27
2 66108 1 27
2 66109 1 27
2 66110 1 27
2 66111 1 27
2 66112 1 27
2 66113 1 27
2 66114 1 27
2 66115 1 27
2 66116 1 27
2 66117 1 27
2 66118 1 27
2 66119 1 27
2 66120 1 27
2 66121 1 27
2 66122 1 27
2 66123 1 27
2 66124 1 27
2 66125 1 27
2 66126 1 27
2 66127 1 27
2 66128 1 27
2 66129 1 27
2 66130 1 27
2 66131 1 27
2 66132 1 27
2 66133 1 27
2 66134 1 27
2 66135 1 27
2 66136 1 27
2 66137 1 27
2 66138 1 27
2 66139 1 27
2 66140 1 27
2 66141 1 27
2 66142 1 27
2 66143 1 27
2 66144 1 27
2 66145 1 27
2 66146 1 27
2 66147 1 27
2 66148 1 27
2 66149 1 27
2 66150 1 27
2 66151 1 27
2 66152 1 27
2 66153 1 27
2 66154 1 27
2 66155 1 27
2 66156 1 27
2 66157 1 27
2 66158 1 27
2 66159 1 27
2 66160 1 27
2 66161 1 27
2 66162 1 27
2 66163 1 27
2 66164 1 27
2 66165 1 27
2 66166 1 27
2 66167 1 27
2 66168 1 27
2 66169 1 27
2 66170 1 27
2 66171 1 27
2 66172 1 27
2 66173 1 27
2 66174 1 27
2 66175 1 27
2 66176 1 27
2 66177 1 27
2 66178 1 27
2 66179 1 27
2 66180 1 27
2 66181 1 27
2 66182 1 27
2 66183 1 27
2 66184 1 27
2 66185 1 27
2 66186 1 27
2 66187 1 27
2 66188 1 27
2 66189 1 27
2 66190 1 27
2 66191 1 27
2 66192 1 27
2 66193 1 27
2 66194 1 27
2 66195 1 27
2 66196 1 27
2 66197 1 27
2 66198 1 27
2 66199 1 27
2 66200 1 27
2 66201 1 27
2 66202 1 27
2 66203 1 27
2 66204 1 27
2 66205 1 28
2 66206 1 28
2 66207 1 28
2 66208 1 28
2 66209 1 28
2 66210 1 28
2 66211 1 28
2 66212 1 28
2 66213 1 28
2 66214 1 28
2 66215 1 28
2 66216 1 28
2 66217 1 28
2 66218 1 28
2 66219 1 28
2 66220 1 28
2 66221 1 28
2 66222 1 28
2 66223 1 28
2 66224 1 28
2 66225 1 28
2 66226 1 28
2 66227 1 28
2 66228 1 28
2 66229 1 28
2 66230 1 28
2 66231 1 28
2 66232 1 28
2 66233 1 28
2 66234 1 28
2 66235 1 28
2 66236 1 28
2 66237 1 28
2 66238 1 28
2 66239 1 28
2 66240 1 28
2 66241 1 28
2 66242 1 28
2 66243 1 28
2 66244 1 28
2 66245 1 28
2 66246 1 28
2 66247 1 28
2 66248 1 28
2 66249 1 28
2 66250 1 28
2 66251 1 28
2 66252 1 28
2 66253 1 28
2 66254 1 28
2 66255 1 28
2 66256 1 28
2 66257 1 28
2 66258 1 28
2 66259 1 28
2 66260 1 28
2 66261 1 28
2 66262 1 28
2 66263 1 28
2 66264 1 28
2 66265 1 28
2 66266 1 28
2 66267 1 28
2 66268 1 28
2 66269 1 28
2 66270 1 28
2 66271 1 28
2 66272 1 28
2 66273 1 28
2 66274 1 28
2 66275 1 28
2 66276 1 28
2 66277 1 28
2 66278 1 28
2 66279 1 28
2 66280 1 28
2 66281 1 28
2 66282 1 28
2 66283 1 28
2 66284 1 28
2 66285 1 28
2 66286 1 28
2 66287 1 28
2 66288 1 28
2 66289 1 28
2 66290 1 28
2 66291 1 28
2 66292 1 28
2 66293 1 28
2 66294 1 28
2 66295 1 28
2 66296 1 28
2 66297 1 28
2 66298 1 28
2 66299 1 28
2 66300 1 28
2 66301 1 28
2 66302 1 28
2 66303 1 28
2 66304 1 28
2 66305 1 28
2 66306 1 28
2 66307 1 28
2 66308 1 28
2 66309 1 28
2 66310 1 28
2 66311 1 28
2 66312 1 28
2 66313 1 28
2 66314 1 28
2 66315 1 28
2 66316 1 28
2 66317 1 28
2 66318 1 28
2 66319 1 28
2 66320 1 28
2 66321 1 28
2 66322 1 28
2 66323 1 28
2 66324 1 28
2 66325 1 28
2 66326 1 28
2 66327 1 28
2 66328 1 28
2 66329 1 28
2 66330 1 28
2 66331 1 28
2 66332 1 28
2 66333 1 28
2 66334 1 28
2 66335 1 28
2 66336 1 28
2 66337 1 28
2 66338 1 29
2 66339 1 29
2 66340 1 29
2 66341 1 29
2 66342 1 29
2 66343 1 29
2 66344 1 29
2 66345 1 29
2 66346 1 29
2 66347 1 29
2 66348 1 29
2 66349 1 29
2 66350 1 29
2 66351 1 29
2 66352 1 29
2 66353 1 29
2 66354 1 29
2 66355 1 29
2 66356 1 29
2 66357 1 29
2 66358 1 29
2 66359 1 29
2 66360 1 29
2 66361 1 29
2 66362 1 29
2 66363 1 29
2 66364 1 29
2 66365 1 29
2 66366 1 29
2 66367 1 29
2 66368 1 29
2 66369 1 29
2 66370 1 29
2 66371 1 29
2 66372 1 29
2 66373 1 29
2 66374 1 29
2 66375 1 29
2 66376 1 29
2 66377 1 29
2 66378 1 29
2 66379 1 29
2 66380 1 29
2 66381 1 29
2 66382 1 29
2 66383 1 29
2 66384 1 29
2 66385 1 29
2 66386 1 29
2 66387 1 29
2 66388 1 29
2 66389 1 29
2 66390 1 29
2 66391 1 29
2 66392 1 29
2 66393 1 29
2 66394 1 29
2 66395 1 29
2 66396 1 29
2 66397 1 29
2 66398 1 29
2 66399 1 29
2 66400 1 29
2 66401 1 29
2 66402 1 29
2 66403 1 29
2 66404 1 29
2 66405 1 29
2 66406 1 29
2 66407 1 29
2 66408 1 29
2 66409 1 29
2 66410 1 29
2 66411 1 29
2 66412 1 29
2 66413 1 29
2 66414 1 29
2 66415 1 29
2 66416 1 29
2 66417 1 29
2 66418 1 29
2 66419 1 29
2 66420 1 29
2 66421 1 29
2 66422 1 29
2 66423 1 29
2 66424 1 29
2 66425 1 29
2 66426 1 29
2 66427 1 29
2 66428 1 29
2 66429 1 29
2 66430 1 29
2 66431 1 29
2 66432 1 29
2 66433 1 29
2 66434 1 29
2 66435 1 29
2 66436 1 29
2 66437 1 29
2 66438 1 29
2 66439 1 29
2 66440 1 29
2 66441 1 29
2 66442 1 29
2 66443 1 29
2 66444 1 29
2 66445 1 29
2 66446 1 29
2 66447 1 29
2 66448 1 29
2 66449 1 29
2 66450 1 29
2 66451 1 29
2 66452 1 29
2 66453 1 29
2 66454 1 29
2 66455 1 29
2 66456 1 29
2 66457 1 29
2 66458 1 29
2 66459 1 29
2 66460 1 29
2 66461 1 29
2 66462 1 29
2 66463 1 29
2 66464 1 29
2 66465 1 29
2 66466 1 29
2 66467 1 29
2 66468 1 29
2 66469 1 29
2 66470 1 29
2 66471 1 29
2 66472 1 29
2 66473 1 29
2 66474 1 29
2 66475 1 29
2 66476 1 29
2 66477 1 29
2 66478 1 29
2 66479 1 29
2 66480 1 29
2 66481 1 29
2 66482 1 29
2 66483 1 29
2 66484 1 29
2 66485 1 29
2 66486 1 29
2 66487 1 29
2 66488 1 29
2 66489 1 29
2 66490 1 29
2 66491 1 29
2 66492 1 29
2 66493 1 29
2 66494 1 29
2 66495 1 29
2 66496 1 29
2 66497 1 29
2 66498 1 29
2 66499 1 29
2 66500 1 29
2 66501 1 29
2 66502 1 29
2 66503 1 29
2 66504 1 29
2 66505 1 29
2 66506 1 29
2 66507 1 29
2 66508 1 29
2 66509 1 29
2 66510 1 29
2 66511 1 29
2 66512 1 29
2 66513 1 29
2 66514 1 29
2 66515 1 29
2 66516 1 29
2 66517 1 29
2 66518 1 29
2 66519 1 29
2 66520 1 29
2 66521 1 29
2 66522 1 29
2 66523 1 29
2 66524 1 29
2 66525 1 29
2 66526 1 29
2 66527 1 29
2 66528 1 29
2 66529 1 29
2 66530 1 29
2 66531 1 29
2 66532 1 29
2 66533 1 29
2 66534 1 29
2 66535 1 29
2 66536 1 29
2 66537 1 29
2 66538 1 29
2 66539 1 29
2 66540 1 29
2 66541 1 29
2 66542 1 29
2 66543 1 29
2 66544 1 29
2 66545 1 29
2 66546 1 29
2 66547 1 29
2 66548 1 29
2 66549 1 29
2 66550 1 29
2 66551 1 29
2 66552 1 29
2 66553 1 29
2 66554 1 29
2 66555 1 29
2 66556 1 29
2 66557 1 29
2 66558 1 29
2 66559 1 29
2 66560 1 29
2 66561 1 29
2 66562 1 29
2 66563 1 29
2 66564 1 29
2 66565 1 29
2 66566 1 29
2 66567 1 29
2 66568 1 29
2 66569 1 29
2 66570 1 29
2 66571 1 29
2 66572 1 29
2 66573 1 29
2 66574 1 29
2 66575 1 29
2 66576 1 30
2 66577 1 30
2 66578 1 30
2 66579 1 30
2 66580 1 30
2 66581 1 30
2 66582 1 30
2 66583 1 30
2 66584 1 30
2 66585 1 30
2 66586 1 30
2 66587 1 30
2 66588 1 30
2 66589 1 30
2 66590 1 30
2 66591 1 30
2 66592 1 30
2 66593 1 30
2 66594 1 30
2 66595 1 30
2 66596 1 30
2 66597 1 30
2 66598 1 30
2 66599 1 30
2 66600 1 30
2 66601 1 30
2 66602 1 30
2 66603 1 30
2 66604 1 30
2 66605 1 30
2 66606 1 30
2 66607 1 30
2 66608 1 30
2 66609 1 30
2 66610 1 30
2 66611 1 30
2 66612 1 30
2 66613 1 30
2 66614 1 30
2 66615 1 30
2 66616 1 30
2 66617 1 30
2 66618 1 30
2 66619 1 30
2 66620 1 30
2 66621 1 30
2 66622 1 30
2 66623 1 30
2 66624 1 30
2 66625 1 30
2 66626 1 30
2 66627 1 30
2 66628 1 30
2 66629 1 30
2 66630 1 30
2 66631 1 30
2 66632 1 30
2 66633 1 30
2 66634 1 30
2 66635 1 30
2 66636 1 30
2 66637 1 30
2 66638 1 30
2 66639 1 30
2 66640 1 30
2 66641 1 30
2 66642 1 30
2 66643 1 30
2 66644 1 30
2 66645 1 30
2 66646 1 30
2 66647 1 30
2 66648 1 30
2 66649 1 30
2 66650 1 30
2 66651 1 30
2 66652 1 30
2 66653 1 30
2 66654 1 30
2 66655 1 30
2 66656 1 30
2 66657 1 30
2 66658 1 30
2 66659 1 30
2 66660 1 30
2 66661 1 30
2 66662 1 30
2 66663 1 30
2 66664 1 30
2 66665 1 30
2 66666 1 30
2 66667 1 30
2 66668 1 30
2 66669 1 30
2 66670 1 30
2 66671 1 30
2 66672 1 30
2 66673 1 30
2 66674 1 30
2 66675 1 30
2 66676 1 30
2 66677 1 30
2 66678 1 30
2 66679 1 30
2 66680 1 30
2 66681 1 30
2 66682 1 30
2 66683 1 30
2 66684 1 30
2 66685 1 30
2 66686 1 30
2 66687 1 30
2 66688 1 30
2 66689 1 30
2 66690 1 30
2 66691 1 30
2 66692 1 30
2 66693 1 30
2 66694 1 30
2 66695 1 30
2 66696 1 30
2 66697 1 30
2 66698 1 30
2 66699 1 30
2 66700 1 30
2 66701 1 30
2 66702 1 30
2 66703 1 30
2 66704 1 30
2 66705 1 30
2 66706 1 30
2 66707 1 30
2 66708 1 30
2 66709 1 30
2 66710 1 30
2 66711 1 30
2 66712 1 30
2 66713 1 30
2 66714 1 30
2 66715 1 30
2 66716 1 30
2 66717 1 30
2 66718 1 30
2 66719 1 30
2 66720 1 30
2 66721 1 30
2 66722 1 30
2 66723 1 30
2 66724 1 30
2 66725 1 30
2 66726 1 30
2 66727 1 30
2 66728 1 30
2 66729 1 30
2 66730 1 30
2 66731 1 30
2 66732 1 30
2 66733 1 30
2 66734 1 30
2 66735 1 30
2 66736 1 30
2 66737 1 30
2 66738 1 30
2 66739 1 30
2 66740 1 30
2 66741 1 30
2 66742 1 30
2 66743 1 30
2 66744 1 30
2 66745 1 30
2 66746 1 30
2 66747 1 30
2 66748 1 30
2 66749 1 30
2 66750 1 30
2 66751 1 30
2 66752 1 30
2 66753 1 30
2 66754 1 30
2 66755 1 30
2 66756 1 30
2 66757 1 30
2 66758 1 30
2 66759 1 30
2 66760 1 30
2 66761 1 30
2 66762 1 30
2 66763 1 30
2 66764 1 30
2 66765 1 30
2 66766 1 30
2 66767 1 30
2 66768 1 30
2 66769 1 30
2 66770 1 30
2 66771 1 30
2 66772 1 30
2 66773 1 30
2 66774 1 30
2 66775 1 30
2 66776 1 30
2 66777 1 30
2 66778 1 30
2 66779 1 30
2 66780 1 30
2 66781 1 30
2 66782 1 30
2 66783 1 30
2 66784 1 30
2 66785 1 30
2 66786 1 30
2 66787 1 30
2 66788 1 30
2 66789 1 30
2 66790 1 30
2 66791 1 30
2 66792 1 30
2 66793 1 30
2 66794 1 30
2 66795 1 30
2 66796 1 30
2 66797 1 30
2 66798 1 30
2 66799 1 31
2 66800 1 31
2 66801 1 31
2 66802 1 31
2 66803 1 31
2 66804 1 31
2 66805 1 31
2 66806 1 31
2 66807 1 31
2 66808 1 31
2 66809 1 31
2 66810 1 31
2 66811 1 31
2 66812 1 31
2 66813 1 31
2 66814 1 31
2 66815 1 31
2 66816 1 31
2 66817 1 31
2 66818 1 31
2 66819 1 31
2 66820 1 31
2 66821 1 31
2 66822 1 31
2 66823 1 31
2 66824 1 31
2 66825 1 31
2 66826 1 31
2 66827 1 31
2 66828 1 31
2 66829 1 31
2 66830 1 31
2 66831 1 31
2 66832 1 31
2 66833 1 31
2 66834 1 31
2 66835 1 31
2 66836 1 31
2 66837 1 31
2 66838 1 31
2 66839 1 31
2 66840 1 31
2 66841 1 31
2 66842 1 31
2 66843 1 31
2 66844 1 31
2 66845 1 31
2 66846 1 31
2 66847 1 31
2 66848 1 31
2 66849 1 31
2 66850 1 31
2 66851 1 31
2 66852 1 31
2 66853 1 31
2 66854 1 31
2 66855 1 31
2 66856 1 31
2 66857 1 31
2 66858 1 31
2 66859 1 31
2 66860 1 31
2 66861 1 31
2 66862 1 31
2 66863 1 31
2 66864 1 31
2 66865 1 31
2 66866 1 31
2 66867 1 31
2 66868 1 31
2 66869 1 31
2 66870 1 31
2 66871 1 31
2 66872 1 31
2 66873 1 31
2 66874 1 31
2 66875 1 31
2 66876 1 31
2 66877 1 31
2 66878 1 31
2 66879 1 31
2 66880 1 31
2 66881 1 31
2 66882 1 31
2 66883 1 31
2 66884 1 31
2 66885 1 31
2 66886 1 31
2 66887 1 31
2 66888 1 31
2 66889 1 31
2 66890 1 31
2 66891 1 31
2 66892 1 31
2 66893 1 31
2 66894 1 31
2 66895 1 31
2 66896 1 31
2 66897 1 31
2 66898 1 31
2 66899 1 31
2 66900 1 31
2 66901 1 31
2 66902 1 31
2 66903 1 31
2 66904 1 31
2 66905 1 31
2 66906 1 31
2 66907 1 31
2 66908 1 31
2 66909 1 31
2 66910 1 31
2 66911 1 31
2 66912 1 31
2 66913 1 31
2 66914 1 31
2 66915 1 31
2 66916 1 31
2 66917 1 31
2 66918 1 31
2 66919 1 31
2 66920 1 31
2 66921 1 31
2 66922 1 31
2 66923 1 31
2 66924 1 31
2 66925 1 31
2 66926 1 31
2 66927 1 31
2 66928 1 31
2 66929 1 31
2 66930 1 31
2 66931 1 31
2 66932 1 31
2 66933 1 31
2 66934 1 31
2 66935 1 31
2 66936 1 31
2 66937 1 31
2 66938 1 31
2 66939 1 31
2 66940 1 31
2 66941 1 31
2 66942 1 31
2 66943 1 31
2 66944 1 31
2 66945 1 31
2 66946 1 31
2 66947 1 31
2 66948 1 31
2 66949 1 31
2 66950 1 31
2 66951 1 31
2 66952 1 31
2 66953 1 31
2 66954 1 31
2 66955 1 31
2 66956 1 31
2 66957 1 31
2 66958 1 31
2 66959 1 31
2 66960 1 31
2 66961 1 31
2 66962 1 31
2 66963 1 31
2 66964 1 31
2 66965 1 31
2 66966 1 31
2 66967 1 31
2 66968 1 31
2 66969 1 31
2 66970 1 31
2 66971 1 31
2 66972 1 31
2 66973 1 31
2 66974 1 31
2 66975 1 31
2 66976 1 31
2 66977 1 31
2 66978 1 31
2 66979 1 31
2 66980 1 31
2 66981 1 31
2 66982 1 31
2 66983 1 31
2 66984 1 31
2 66985 1 31
2 66986 1 31
2 66987 1 31
2 66988 1 31
2 66989 1 31
2 66990 1 31
2 66991 1 31
2 66992 1 31
2 66993 1 31
2 66994 1 31
2 66995 1 31
2 66996 1 31
2 66997 1 31
2 66998 1 31
2 66999 1 31
2 67000 1 31
2 67001 1 31
2 67002 1 31
2 67003 1 31
2 67004 1 31
2 67005 1 31
2 67006 1 31
2 67007 1 31
2 67008 1 31
2 67009 1 31
2 67010 1 31
2 67011 1 31
2 67012 1 31
2 67013 1 31
2 67014 1 31
2 67015 1 31
2 67016 1 31
2 67017 1 31
2 67018 1 31
2 67019 1 31
2 67020 1 31
2 67021 1 31
2 67022 1 31
2 67023 1 31
2 67024 1 31
2 67025 1 31
2 67026 1 31
2 67027 1 31
2 67028 1 31
2 67029 1 31
2 67030 1 31
2 67031 1 31
2 67032 1 31
2 67033 1 31
2 67034 1 31
2 67035 1 31
2 67036 1 31
2 67037 1 31
2 67038 1 31
2 67039 1 31
2 67040 1 31
2 67041 1 31
2 67042 1 31
2 67043 1 31
2 67044 1 31
2 67045 1 31
2 67046 1 31
2 67047 1 31
2 67048 1 31
2 67049 1 31
2 67050 1 31
2 67051 1 31
2 67052 1 31
2 67053 1 31
2 67054 1 31
2 67055 1 31
2 67056 1 31
2 67057 1 31
2 67058 1 31
2 67059 1 31
2 67060 1 31
2 67061 1 31
2 67062 1 31
2 67063 1 31
2 67064 1 31
2 67065 1 31
2 67066 1 31
2 67067 1 31
2 67068 1 31
2 67069 1 31
2 67070 1 31
2 67071 1 31
2 67072 1 31
2 67073 1 31
2 67074 1 31
2 67075 1 31
2 67076 1 31
2 67077 1 31
2 67078 1 31
2 67079 1 31
2 67080 1 31
2 67081 1 31
2 67082 1 31
2 67083 1 31
2 67084 1 31
2 67085 1 31
2 67086 1 31
2 67087 1 31
2 67088 1 31
2 67089 1 31
2 67090 1 31
2 67091 1 31
2 67092 1 31
2 67093 1 31
2 67094 1 31
2 67095 1 31
2 67096 1 31
2 67097 1 31
2 67098 1 31
2 67099 1 31
2 67100 1 31
2 67101 1 32
2 67102 1 32
2 67103 1 32
2 67104 1 32
2 67105 1 32
2 67106 1 32
2 67107 1 32
2 67108 1 32
2 67109 1 32
2 67110 1 32
2 67111 1 32
2 67112 1 32
2 67113 1 32
2 67114 1 32
2 67115 1 32
2 67116 1 32
2 67117 1 32
2 67118 1 32
2 67119 1 32
2 67120 1 32
2 67121 1 32
2 67122 1 32
2 67123 1 32
2 67124 1 32
2 67125 1 32
2 67126 1 32
2 67127 1 32
2 67128 1 32
2 67129 1 32
2 67130 1 32
2 67131 1 32
2 67132 1 32
2 67133 1 32
2 67134 1 32
2 67135 1 32
2 67136 1 32
2 67137 1 32
2 67138 1 32
2 67139 1 32
2 67140 1 32
2 67141 1 32
2 67142 1 32
2 67143 1 32
2 67144 1 32
2 67145 1 32
2 67146 1 32
2 67147 1 32
2 67148 1 32
2 67149 1 32
2 67150 1 32
2 67151 1 32
2 67152 1 32
2 67153 1 32
2 67154 1 32
2 67155 1 32
2 67156 1 32
2 67157 1 32
2 67158 1 32
2 67159 1 32
2 67160 1 32
2 67161 1 32
2 67162 1 32
2 67163 1 32
2 67164 1 32
2 67165 1 32
2 67166 1 32
2 67167 1 32
2 67168 1 32
2 67169 1 32
2 67170 1 32
2 67171 1 32
2 67172 1 32
2 67173 1 32
2 67174 1 32
2 67175 1 32
2 67176 1 32
2 67177 1 32
2 67178 1 32
2 67179 1 32
2 67180 1 32
2 67181 1 32
2 67182 1 32
2 67183 1 32
2 67184 1 32
2 67185 1 32
2 67186 1 32
2 67187 1 32
2 67188 1 32
2 67189 1 32
2 67190 1 32
2 67191 1 32
2 67192 1 32
2 67193 1 32
2 67194 1 32
2 67195 1 32
2 67196 1 32
2 67197 1 32
2 67198 1 32
2 67199 1 32
2 67200 1 32
2 67201 1 32
2 67202 1 32
2 67203 1 32
2 67204 1 32
2 67205 1 32
2 67206 1 32
2 67207 1 32
2 67208 1 32
2 67209 1 32
2 67210 1 32
2 67211 1 32
2 67212 1 32
2 67213 1 32
2 67214 1 32
2 67215 1 32
2 67216 1 32
2 67217 1 32
2 67218 1 32
2 67219 1 32
2 67220 1 32
2 67221 1 32
2 67222 1 32
2 67223 1 32
2 67224 1 32
2 67225 1 32
2 67226 1 32
2 67227 1 32
2 67228 1 32
2 67229 1 32
2 67230 1 32
2 67231 1 32
2 67232 1 32
2 67233 1 32
2 67234 1 32
2 67235 1 32
2 67236 1 32
2 67237 1 32
2 67238 1 32
2 67239 1 32
2 67240 1 32
2 67241 1 32
2 67242 1 32
2 67243 1 32
2 67244 1 32
2 67245 1 32
2 67246 1 32
2 67247 1 32
2 67248 1 32
2 67249 1 32
2 67250 1 32
2 67251 1 32
2 67252 1 32
2 67253 1 32
2 67254 1 32
2 67255 1 32
2 67256 1 32
2 67257 1 32
2 67258 1 32
2 67259 1 32
2 67260 1 32
2 67261 1 32
2 67262 1 32
2 67263 1 32
2 67264 1 32
2 67265 1 32
2 67266 1 32
2 67267 1 32
2 67268 1 32
2 67269 1 32
2 67270 1 32
2 67271 1 32
2 67272 1 32
2 67273 1 32
2 67274 1 32
2 67275 1 32
2 67276 1 32
2 67277 1 32
2 67278 1 32
2 67279 1 32
2 67280 1 32
2 67281 1 32
2 67282 1 32
2 67283 1 32
2 67284 1 32
2 67285 1 32
2 67286 1 32
2 67287 1 32
2 67288 1 32
2 67289 1 32
2 67290 1 32
2 67291 1 32
2 67292 1 32
2 67293 1 32
2 67294 1 32
2 67295 1 32
2 67296 1 32
2 67297 1 32
2 67298 1 32
2 67299 1 32
2 67300 1 32
2 67301 1 32
2 67302 1 32
2 67303 1 32
2 67304 1 32
2 67305 1 32
2 67306 1 32
2 67307 1 32
2 67308 1 32
2 67309 1 32
2 67310 1 32
2 67311 1 32
2 67312 1 32
2 67313 1 32
2 67314 1 32
2 67315 1 32
2 67316 1 32
2 67317 1 32
2 67318 1 33
2 67319 1 33
2 67320 1 33
2 67321 1 33
2 67322 1 33
2 67323 1 33
2 67324 1 33
2 67325 1 33
2 67326 1 33
2 67327 1 33
2 67328 1 33
2 67329 1 33
2 67330 1 33
2 67331 1 33
2 67332 1 33
2 67333 1 33
2 67334 1 33
2 67335 1 33
2 67336 1 33
2 67337 1 33
2 67338 1 33
2 67339 1 33
2 67340 1 33
2 67341 1 33
2 67342 1 33
2 67343 1 33
2 67344 1 33
2 67345 1 33
2 67346 1 33
2 67347 1 33
2 67348 1 33
2 67349 1 33
2 67350 1 33
2 67351 1 33
2 67352 1 33
2 67353 1 33
2 67354 1 33
2 67355 1 33
2 67356 1 33
2 67357 1 33
2 67358 1 33
2 67359 1 33
2 67360 1 33
2 67361 1 33
2 67362 1 33
2 67363 1 33
2 67364 1 33
2 67365 1 33
2 67366 1 33
2 67367 1 33
2 67368 1 33
2 67369 1 33
2 67370 1 33
2 67371 1 33
2 67372 1 33
2 67373 1 33
2 67374 1 33
2 67375 1 33
2 67376 1 33
2 67377 1 33
2 67378 1 33
2 67379 1 33
2 67380 1 33
2 67381 1 33
2 67382 1 33
2 67383 1 33
2 67384 1 33
2 67385 1 33
2 67386 1 33
2 67387 1 33
2 67388 1 33
2 67389 1 33
2 67390 1 33
2 67391 1 33
2 67392 1 33
2 67393 1 33
2 67394 1 33
2 67395 1 33
2 67396 1 33
2 67397 1 33
2 67398 1 33
2 67399 1 33
2 67400 1 33
2 67401 1 33
2 67402 1 33
2 67403 1 33
2 67404 1 33
2 67405 1 33
2 67406 1 33
2 67407 1 33
2 67408 1 33
2 67409 1 33
2 67410 1 33
2 67411 1 33
2 67412 1 33
2 67413 1 33
2 67414 1 33
2 67415 1 33
2 67416 1 33
2 67417 1 33
2 67418 1 33
2 67419 1 33
2 67420 1 33
2 67421 1 33
2 67422 1 33
2 67423 1 33
2 67424 1 33
2 67425 1 33
2 67426 1 33
2 67427 1 33
2 67428 1 33
2 67429 1 33
2 67430 1 33
2 67431 1 33
2 67432 1 33
2 67433 1 33
2 67434 1 33
2 67435 1 33
2 67436 1 33
2 67437 1 33
2 67438 1 33
2 67439 1 33
2 67440 1 33
2 67441 1 33
2 67442 1 33
2 67443 1 33
2 67444 1 33
2 67445 1 33
2 67446 1 33
2 67447 1 33
2 67448 1 33
2 67449 1 33
2 67450 1 33
2 67451 1 33
2 67452 1 33
2 67453 1 33
2 67454 1 33
2 67455 1 33
2 67456 1 33
2 67457 1 33
2 67458 1 33
2 67459 1 33
2 67460 1 33
2 67461 1 33
2 67462 1 33
2 67463 1 33
2 67464 1 33
2 67465 1 33
2 67466 1 33
2 67467 1 33
2 67468 1 33
2 67469 1 33
2 67470 1 33
2 67471 1 33
2 67472 1 33
2 67473 1 33
2 67474 1 33
2 67475 1 33
2 67476 1 33
2 67477 1 33
2 67478 1 33
2 67479 1 33
2 67480 1 33
2 67481 1 33
2 67482 1 33
2 67483 1 33
2 67484 1 33
2 67485 1 33
2 67486 1 33
2 67487 1 33
2 67488 1 33
2 67489 1 33
2 67490 1 33
2 67491 1 33
2 67492 1 33
2 67493 1 33
2 67494 1 33
2 67495 1 33
2 67496 1 33
2 67497 1 33
2 67498 1 33
2 67499 1 33
2 67500 1 33
2 67501 1 33
2 67502 1 33
2 67503 1 33
2 67504 1 33
2 67505 1 33
2 67506 1 33
2 67507 1 33
2 67508 1 33
2 67509 1 33
2 67510 1 33
2 67511 1 33
2 67512 1 33
2 67513 1 33
2 67514 1 33
2 67515 1 33
2 67516 1 33
2 67517 1 33
2 67518 1 33
2 67519 1 33
2 67520 1 33
2 67521 1 33
2 67522 1 33
2 67523 1 33
2 67524 1 33
2 67525 1 33
2 67526 1 33
2 67527 1 33
2 67528 1 33
2 67529 1 33
2 67530 1 33
2 67531 1 33
2 67532 1 33
2 67533 1 33
2 67534 1 33
2 67535 1 33
2 67536 1 33
2 67537 1 33
2 67538 1 33
2 67539 1 33
2 67540 1 33
2 67541 1 33
2 67542 1 33
2 67543 1 33
2 67544 1 33
2 67545 1 33
2 67546 1 33
2 67547 1 34
2 67548 1 34
2 67549 1 34
2 67550 1 34
2 67551 1 34
2 67552 1 34
2 67553 1 34
2 67554 1 34
2 67555 1 34
2 67556 1 34
2 67557 1 34
2 67558 1 34
2 67559 1 34
2 67560 1 34
2 67561 1 34
2 67562 1 34
2 67563 1 34
2 67564 1 34
2 67565 1 34
2 67566 1 34
2 67567 1 34
2 67568 1 34
2 67569 1 34
2 67570 1 34
2 67571 1 34
2 67572 1 34
2 67573 1 34
2 67574 1 34
2 67575 1 34
2 67576 1 34
2 67577 1 34
2 67578 1 34
2 67579 1 34
2 67580 1 34
2 67581 1 34
2 67582 1 34
2 67583 1 34
2 67584 1 34
2 67585 1 34
2 67586 1 34
2 67587 1 34
2 67588 1 34
2 67589 1 34
2 67590 1 34
2 67591 1 34
2 67592 1 34
2 67593 1 34
2 67594 1 34
2 67595 1 34
2 67596 1 34
2 67597 1 34
2 67598 1 34
2 67599 1 34
2 67600 1 34
2 67601 1 34
2 67602 1 34
2 67603 1 34
2 67604 1 34
2 67605 1 34
2 67606 1 34
2 67607 1 34
2 67608 1 34
2 67609 1 34
2 67610 1 34
2 67611 1 34
2 67612 1 34
2 67613 1 34
2 67614 1 34
2 67615 1 34
2 67616 1 34
2 67617 1 34
2 67618 1 34
2 67619 1 34
2 67620 1 34
2 67621 1 34
2 67622 1 34
2 67623 1 34
2 67624 1 34
2 67625 1 34
2 67626 1 34
2 67627 1 34
2 67628 1 34
2 67629 1 34
2 67630 1 34
2 67631 1 34
2 67632 1 34
2 67633 1 34
2 67634 1 34
2 67635 1 34
2 67636 1 34
2 67637 1 34
2 67638 1 34
2 67639 1 34
2 67640 1 34
2 67641 1 34
2 67642 1 34
2 67643 1 34
2 67644 1 34
2 67645 1 34
2 67646 1 34
2 67647 1 34
2 67648 1 34
2 67649 1 34
2 67650 1 34
2 67651 1 34
2 67652 1 34
2 67653 1 34
2 67654 1 34
2 67655 1 34
2 67656 1 34
2 67657 1 34
2 67658 1 34
2 67659 1 34
2 67660 1 34
2 67661 1 34
2 67662 1 34
2 67663 1 34
2 67664 1 34
2 67665 1 34
2 67666 1 34
2 67667 1 34
2 67668 1 34
2 67669 1 34
2 67670 1 34
2 67671 1 34
2 67672 1 34
2 67673 1 34
2 67674 1 34
2 67675 1 34
2 67676 1 34
2 67677 1 34
2 67678 1 34
2 67679 1 34
2 67680 1 34
2 67681 1 34
2 67682 1 34
2 67683 1 34
2 67684 1 34
2 67685 1 34
2 67686 1 34
2 67687 1 34
2 67688 1 34
2 67689 1 34
2 67690 1 34
2 67691 1 34
2 67692 1 34
2 67693 1 34
2 67694 1 34
2 67695 1 34
2 67696 1 34
2 67697 1 34
2 67698 1 34
2 67699 1 34
2 67700 1 34
2 67701 1 34
2 67702 1 34
2 67703 1 34
2 67704 1 34
2 67705 1 34
2 67706 1 34
2 67707 1 34
2 67708 1 34
2 67709 1 34
2 67710 1 34
2 67711 1 34
2 67712 1 34
2 67713 1 34
2 67714 1 34
2 67715 1 34
2 67716 1 34
2 67717 1 34
2 67718 1 34
2 67719 1 34
2 67720 1 34
2 67721 1 34
2 67722 1 34
2 67723 1 34
2 67724 1 34
2 67725 1 34
2 67726 1 34
2 67727 1 34
2 67728 1 34
2 67729 1 34
2 67730 1 34
2 67731 1 34
2 67732 1 34
2 67733 1 34
2 67734 1 34
2 67735 1 34
2 67736 1 34
2 67737 1 34
2 67738 1 34
2 67739 1 34
2 67740 1 34
2 67741 1 34
2 67742 1 34
2 67743 1 34
2 67744 1 34
2 67745 1 34
2 67746 1 34
2 67747 1 34
2 67748 1 34
2 67749 1 34
2 67750 1 34
2 67751 1 34
2 67752 1 34
2 67753 1 34
2 67754 1 34
2 67755 1 34
2 67756 1 34
2 67757 1 34
2 67758 1 34
2 67759 1 34
2 67760 1 35
2 67761 1 35
2 67762 1 35
2 67763 1 35
2 67764 1 35
2 67765 1 35
2 67766 1 35
2 67767 1 35
2 67768 1 35
2 67769 1 35
2 67770 1 35
2 67771 1 35
2 67772 1 35
2 67773 1 35
2 67774 1 35
2 67775 1 35
2 67776 1 35
2 67777 1 35
2 67778 1 35
2 67779 1 35
2 67780 1 35
2 67781 1 35
2 67782 1 35
2 67783 1 35
2 67784 1 35
2 67785 1 35
2 67786 1 35
2 67787 1 35
2 67788 1 35
2 67789 1 35
2 67790 1 35
2 67791 1 35
2 67792 1 35
2 67793 1 35
2 67794 1 35
2 67795 1 35
2 67796 1 35
2 67797 1 35
2 67798 1 35
2 67799 1 35
2 67800 1 35
2 67801 1 35
2 67802 1 35
2 67803 1 35
2 67804 1 35
2 67805 1 35
2 67806 1 35
2 67807 1 35
2 67808 1 35
2 67809 1 35
2 67810 1 35
2 67811 1 35
2 67812 1 35
2 67813 1 35
2 67814 1 35
2 67815 1 35
2 67816 1 35
2 67817 1 35
2 67818 1 35
2 67819 1 35
2 67820 1 35
2 67821 1 35
2 67822 1 35
2 67823 1 35
2 67824 1 35
2 67825 1 35
2 67826 1 35
2 67827 1 35
2 67828 1 35
2 67829 1 35
2 67830 1 35
2 67831 1 35
2 67832 1 35
2 67833 1 35
2 67834 1 35
2 67835 1 35
2 67836 1 35
2 67837 1 36
2 67838 1 36
2 67839 1 36
2 67840 1 36
2 67841 1 36
2 67842 1 36
2 67843 1 36
2 67844 1 36
2 67845 1 36
2 67846 1 36
2 67847 1 36
2 67848 1 36
2 67849 1 36
2 67850 1 36
2 67851 1 36
2 67852 1 36
2 67853 1 36
2 67854 1 36
2 67855 1 36
2 67856 1 36
2 67857 1 36
2 67858 1 36
2 67859 1 36
2 67860 1 36
2 67861 1 36
2 67862 1 36
2 67863 1 36
2 67864 1 36
2 67865 1 36
2 67866 1 36
2 67867 1 36
2 67868 1 36
2 67869 1 36
2 67870 1 36
2 67871 1 36
2 67872 1 36
2 67873 1 36
2 67874 1 36
2 67875 1 36
2 67876 1 36
2 67877 1 36
2 67878 1 36
2 67879 1 36
2 67880 1 36
2 67881 1 36
2 67882 1 36
2 67883 1 36
2 67884 1 36
2 67885 1 36
2 67886 1 36
2 67887 1 36
2 67888 1 36
2 67889 1 36
2 67890 1 36
2 67891 1 36
2 67892 1 36
2 67893 1 36
2 67894 1 36
2 67895 1 36
2 67896 1 36
2 67897 1 36
2 67898 1 36
2 67899 1 36
2 67900 1 36
2 67901 1 36
2 67902 1 36
2 67903 1 36
2 67904 1 36
2 67905 1 36
2 67906 1 36
2 67907 1 36
2 67908 1 36
2 67909 1 37
2 67910 1 37
2 67911 1 37
2 67912 1 37
2 67913 1 37
2 67914 1 37
2 67915 1 37
2 67916 1 37
2 67917 1 37
2 67918 1 37
2 67919 1 37
2 67920 1 37
2 67921 1 37
2 67922 1 37
2 67923 1 37
2 67924 1 37
2 67925 1 37
2 67926 1 37
2 67927 1 37
2 67928 1 37
2 67929 1 37
2 67930 1 37
2 67931 1 37
2 67932 1 37
2 67933 1 37
2 67934 1 37
2 67935 1 37
2 67936 1 37
2 67937 1 37
2 67938 1 37
2 67939 1 37
2 67940 1 37
2 67941 1 37
2 67942 1 37
2 67943 1 37
2 67944 1 37
2 67945 1 37
2 67946 1 37
2 67947 1 37
2 67948 1 37
2 67949 1 37
2 67950 1 37
2 67951 1 37
2 67952 1 37
2 67953 1 37
2 67954 1 37
2 67955 1 37
2 67956 1 37
2 67957 1 37
2 67958 1 37
2 67959 1 37
2 67960 1 37
2 67961 1 37
2 67962 1 37
2 67963 1 37
2 67964 1 37
2 67965 1 37
2 67966 1 37
2 67967 1 37
2 67968 1 37
2 67969 1 37
2 67970 1 37
2 67971 1 37
2 67972 1 37
2 67973 1 37
2 67974 1 37
2 67975 1 37
2 67976 1 37
2 67977 1 37
2 67978 1 37
2 67979 1 37
2 67980 1 37
2 67981 1 37
2 67982 1 37
2 67983 1 37
2 67984 1 37
2 67985 1 37
2 67986 1 37
2 67987 1 37
2 67988 1 37
2 67989 1 37
2 67990 1 37
2 67991 1 37
2 67992 1 37
2 67993 1 37
2 67994 1 37
2 67995 1 37
2 67996 1 37
2 67997 1 37
2 67998 1 37
2 67999 1 37
2 68000 1 37
2 68001 1 37
2 68002 1 37
2 68003 1 37
2 68004 1 37
2 68005 1 37
2 68006 1 37
2 68007 1 37
2 68008 1 37
2 68009 1 37
2 68010 1 37
2 68011 1 37
2 68012 1 37
2 68013 1 37
2 68014 1 37
2 68015 1 37
2 68016 1 37
2 68017 1 37
2 68018 1 37
2 68019 1 37
2 68020 1 37
2 68021 1 37
2 68022 1 37
2 68023 1 37
2 68024 1 37
2 68025 1 37
2 68026 1 37
2 68027 1 37
2 68028 1 37
2 68029 1 37
2 68030 1 37
2 68031 1 37
2 68032 1 37
2 68033 1 37
2 68034 1 37
2 68035 1 37
2 68036 1 37
2 68037 1 37
2 68038 1 37
2 68039 1 37
2 68040 1 37
2 68041 1 37
2 68042 1 37
2 68043 1 37
2 68044 1 37
2 68045 1 37
2 68046 1 37
2 68047 1 37
2 68048 1 37
2 68049 1 37
2 68050 1 37
2 68051 1 37
2 68052 1 37
2 68053 1 37
2 68054 1 38
2 68055 1 38
2 68056 1 38
2 68057 1 38
2 68058 1 38
2 68059 1 38
2 68060 1 38
2 68061 1 38
2 68062 1 38
2 68063 1 38
2 68064 1 38
2 68065 1 38
2 68066 1 38
2 68067 1 38
2 68068 1 38
2 68069 1 38
2 68070 1 38
2 68071 1 38
2 68072 1 38
2 68073 1 38
2 68074 1 38
2 68075 1 38
2 68076 1 38
2 68077 1 38
2 68078 1 38
2 68079 1 38
2 68080 1 38
2 68081 1 38
2 68082 1 38
2 68083 1 38
2 68084 1 38
2 68085 1 38
2 68086 1 38
2 68087 1 38
2 68088 1 38
2 68089 1 38
2 68090 1 38
2 68091 1 38
2 68092 1 38
2 68093 1 38
2 68094 1 38
2 68095 1 38
2 68096 1 38
2 68097 1 38
2 68098 1 38
2 68099 1 38
2 68100 1 38
2 68101 1 38
2 68102 1 38
2 68103 1 38
2 68104 1 38
2 68105 1 38
2 68106 1 38
2 68107 1 38
2 68108 1 38
2 68109 1 38
2 68110 1 38
2 68111 1 38
2 68112 1 38
2 68113 1 38
2 68114 1 38
2 68115 1 38
2 68116 1 38
2 68117 1 38
2 68118 1 38
2 68119 1 38
2 68120 1 38
2 68121 1 38
2 68122 1 38
2 68123 1 38
2 68124 1 38
2 68125 1 38
2 68126 1 38
2 68127 1 38
2 68128 1 38
2 68129 1 38
2 68130 1 38
2 68131 1 38
2 68132 1 38
2 68133 1 38
2 68134 1 38
2 68135 1 38
2 68136 1 38
2 68137 1 38
2 68138 1 38
2 68139 1 38
2 68140 1 38
2 68141 1 38
2 68142 1 38
2 68143 1 38
2 68144 1 38
2 68145 1 38
2 68146 1 38
2 68147 1 38
2 68148 1 38
2 68149 1 38
2 68150 1 38
2 68151 1 38
2 68152 1 38
2 68153 1 38
2 68154 1 38
2 68155 1 38
2 68156 1 38
2 68157 1 38
2 68158 1 38
2 68159 1 38
2 68160 1 38
2 68161 1 38
2 68162 1 38
2 68163 1 38
2 68164 1 38
2 68165 1 38
2 68166 1 38
2 68167 1 38
2 68168 1 38
2 68169 1 38
2 68170 1 38
2 68171 1 38
2 68172 1 38
2 68173 1 38
2 68174 1 38
2 68175 1 38
2 68176 1 38
2 68177 1 38
2 68178 1 38
2 68179 1 38
2 68180 1 38
2 68181 1 38
2 68182 1 38
2 68183 1 38
2 68184 1 38
2 68185 1 38
2 68186 1 38
2 68187 1 38
2 68188 1 38
2 68189 1 38
2 68190 1 38
2 68191 1 38
2 68192 1 38
2 68193 1 38
2 68194 1 38
2 68195 1 38
2 68196 1 38
2 68197 1 38
2 68198 1 38
2 68199 1 38
2 68200 1 38
2 68201 1 38
2 68202 1 38
2 68203 1 38
2 68204 1 38
2 68205 1 38
2 68206 1 38
2 68207 1 38
2 68208 1 38
2 68209 1 38
2 68210 1 38
2 68211 1 38
2 68212 1 38
2 68213 1 38
2 68214 1 38
2 68215 1 38
2 68216 1 38
2 68217 1 38
2 68218 1 38
2 68219 1 38
2 68220 1 38
2 68221 1 38
2 68222 1 38
2 68223 1 38
2 68224 1 38
2 68225 1 38
2 68226 1 38
2 68227 1 38
2 68228 1 38
2 68229 1 38
2 68230 1 38
2 68231 1 38
2 68232 1 38
2 68233 1 38
2 68234 1 38
2 68235 1 38
2 68236 1 38
2 68237 1 38
2 68238 1 38
2 68239 1 38
2 68240 1 38
2 68241 1 38
2 68242 1 38
2 68243 1 38
2 68244 1 38
2 68245 1 38
2 68246 1 38
2 68247 1 38
2 68248 1 38
2 68249 1 38
2 68250 1 38
2 68251 1 39
2 68252 1 39
2 68253 1 39
2 68254 1 39
2 68255 1 39
2 68256 1 39
2 68257 1 39
2 68258 1 39
2 68259 1 39
2 68260 1 39
2 68261 1 39
2 68262 1 39
2 68263 1 39
2 68264 1 39
2 68265 1 39
2 68266 1 39
2 68267 1 39
2 68268 1 39
2 68269 1 39
2 68270 1 39
2 68271 1 39
2 68272 1 39
2 68273 1 39
2 68274 1 39
2 68275 1 39
2 68276 1 39
2 68277 1 39
2 68278 1 39
2 68279 1 39
2 68280 1 39
2 68281 1 39
2 68282 1 39
2 68283 1 39
2 68284 1 39
2 68285 1 39
2 68286 1 39
2 68287 1 39
2 68288 1 39
2 68289 1 39
2 68290 1 39
2 68291 1 39
2 68292 1 39
2 68293 1 39
2 68294 1 39
2 68295 1 39
2 68296 1 39
2 68297 1 39
2 68298 1 39
2 68299 1 39
2 68300 1 39
2 68301 1 39
2 68302 1 39
2 68303 1 39
2 68304 1 39
2 68305 1 39
2 68306 1 39
2 68307 1 39
2 68308 1 39
2 68309 1 39
2 68310 1 39
2 68311 1 39
2 68312 1 39
2 68313 1 39
2 68314 1 39
2 68315 1 39
2 68316 1 39
2 68317 1 39
2 68318 1 39
2 68319 1 39
2 68320 1 39
2 68321 1 39
2 68322 1 39
2 68323 1 39
2 68324 1 39
2 68325 1 39
2 68326 1 39
2 68327 1 39
2 68328 1 39
2 68329 1 39
2 68330 1 39
2 68331 1 39
2 68332 1 39
2 68333 1 39
2 68334 1 39
2 68335 1 39
2 68336 1 39
2 68337 1 39
2 68338 1 39
2 68339 1 39
2 68340 1 39
2 68341 1 39
2 68342 1 39
2 68343 1 39
2 68344 1 39
2 68345 1 39
2 68346 1 39
2 68347 1 39
2 68348 1 39
2 68349 1 39
2 68350 1 39
2 68351 1 39
2 68352 1 39
2 68353 1 39
2 68354 1 39
2 68355 1 39
2 68356 1 39
2 68357 1 39
2 68358 1 39
2 68359 1 39
2 68360 1 39
2 68361 1 39
2 68362 1 39
2 68363 1 39
2 68364 1 39
2 68365 1 39
2 68366 1 39
2 68367 1 39
2 68368 1 39
2 68369 1 39
2 68370 1 39
2 68371 1 39
2 68372 1 39
2 68373 1 39
2 68374 1 39
2 68375 1 39
2 68376 1 39
2 68377 1 39
2 68378 1 39
2 68379 1 39
2 68380 1 39
2 68381 1 39
2 68382 1 39
2 68383 1 39
2 68384 1 39
2 68385 1 39
2 68386 1 39
2 68387 1 39
2 68388 1 39
2 68389 1 39
2 68390 1 39
2 68391 1 39
2 68392 1 39
2 68393 1 39
2 68394 1 39
2 68395 1 39
2 68396 1 39
2 68397 1 39
2 68398 1 39
2 68399 1 39
2 68400 1 39
2 68401 1 39
2 68402 1 39
2 68403 1 39
2 68404 1 39
2 68405 1 39
2 68406 1 39
2 68407 1 39
2 68408 1 39
2 68409 1 39
2 68410 1 39
2 68411 1 39
2 68412 1 39
2 68413 1 39
2 68414 1 39
2 68415 1 39
2 68416 1 39
2 68417 1 39
2 68418 1 39
2 68419 1 39
2 68420 1 39
2 68421 1 39
2 68422 1 39
2 68423 1 39
2 68424 1 39
2 68425 1 39
2 68426 1 39
2 68427 1 39
2 68428 1 39
2 68429 1 39
2 68430 1 39
2 68431 1 39
2 68432 1 39
2 68433 1 39
2 68434 1 39
2 68435 1 39
2 68436 1 39
2 68437 1 39
2 68438 1 39
2 68439 1 39
2 68440 1 39
2 68441 1 39
2 68442 1 39
2 68443 1 39
2 68444 1 39
2 68445 1 39
2 68446 1 39
2 68447 1 39
2 68448 1 39
2 68449 1 39
2 68450 1 39
2 68451 1 39
2 68452 1 39
2 68453 1 39
2 68454 1 39
2 68455 1 39
2 68456 1 39
2 68457 1 39
2 68458 1 39
2 68459 1 39
2 68460 1 39
2 68461 1 39
2 68462 1 39
2 68463 1 39
2 68464 1 39
2 68465 1 39
2 68466 1 39
2 68467 1 39
2 68468 1 39
2 68469 1 39
2 68470 1 39
2 68471 1 39
2 68472 1 39
2 68473 1 39
2 68474 1 39
2 68475 1 39
2 68476 1 39
2 68477 1 39
2 68478 1 39
2 68479 1 39
2 68480 1 39
2 68481 1 39
2 68482 1 39
2 68483 1 39
2 68484 1 39
2 68485 1 39
2 68486 1 39
2 68487 1 39
2 68488 1 39
2 68489 1 39
2 68490 1 39
2 68491 1 39
2 68492 1 39
2 68493 1 39
2 68494 1 39
2 68495 1 39
2 68496 1 39
2 68497 1 40
2 68498 1 40
2 68499 1 40
2 68500 1 40
2 68501 1 40
2 68502 1 40
2 68503 1 40
2 68504 1 40
2 68505 1 40
2 68506 1 40
2 68507 1 40
2 68508 1 40
2 68509 1 40
2 68510 1 40
2 68511 1 40
2 68512 1 40
2 68513 1 40
2 68514 1 40
2 68515 1 40
2 68516 1 40
2 68517 1 40
2 68518 1 40
2 68519 1 40
2 68520 1 40
2 68521 1 40
2 68522 1 40
2 68523 1 40
2 68524 1 40
2 68525 1 40
2 68526 1 40
2 68527 1 40
2 68528 1 40
2 68529 1 40
2 68530 1 40
2 68531 1 40
2 68532 1 40
2 68533 1 40
2 68534 1 40
2 68535 1 40
2 68536 1 40
2 68537 1 40
2 68538 1 40
2 68539 1 40
2 68540 1 40
2 68541 1 40
2 68542 1 40
2 68543 1 40
2 68544 1 40
2 68545 1 40
2 68546 1 40
2 68547 1 40
2 68548 1 40
2 68549 1 40
2 68550 1 40
2 68551 1 40
2 68552 1 40
2 68553 1 40
2 68554 1 40
2 68555 1 40
2 68556 1 40
2 68557 1 40
2 68558 1 40
2 68559 1 40
2 68560 1 40
2 68561 1 40
2 68562 1 40
2 68563 1 40
2 68564 1 40
2 68565 1 40
2 68566 1 40
2 68567 1 40
2 68568 1 40
2 68569 1 40
2 68570 1 40
2 68571 1 40
2 68572 1 40
2 68573 1 40
2 68574 1 40
2 68575 1 40
2 68576 1 40
2 68577 1 40
2 68578 1 40
2 68579 1 40
2 68580 1 40
2 68581 1 40
2 68582 1 40
2 68583 1 40
2 68584 1 40
2 68585 1 40
2 68586 1 40
2 68587 1 40
2 68588 1 40
2 68589 1 40
2 68590 1 40
2 68591 1 40
2 68592 1 40
2 68593 1 40
2 68594 1 40
2 68595 1 40
2 68596 1 40
2 68597 1 40
2 68598 1 40
2 68599 1 40
2 68600 1 40
2 68601 1 40
2 68602 1 40
2 68603 1 40
2 68604 1 40
2 68605 1 40
2 68606 1 40
2 68607 1 40
2 68608 1 40
2 68609 1 40
2 68610 1 40
2 68611 1 40
2 68612 1 40
2 68613 1 40
2 68614 1 40
2 68615 1 40
2 68616 1 40
2 68617 1 40
2 68618 1 40
2 68619 1 40
2 68620 1 40
2 68621 1 40
2 68622 1 40
2 68623 1 40
2 68624 1 40
2 68625 1 40
2 68626 1 40
2 68627 1 40
2 68628 1 40
2 68629 1 40
2 68630 1 40
2 68631 1 40
2 68632 1 40
2 68633 1 40
2 68634 1 40
2 68635 1 40
2 68636 1 40
2 68637 1 40
2 68638 1 40
2 68639 1 40
2 68640 1 40
2 68641 1 40
2 68642 1 40
2 68643 1 40
2 68644 1 40
2 68645 1 40
2 68646 1 40
2 68647 1 40
2 68648 1 40
2 68649 1 40
2 68650 1 40
2 68651 1 40
2 68652 1 40
2 68653 1 40
2 68654 1 40
2 68655 1 40
2 68656 1 40
2 68657 1 40
2 68658 1 40
2 68659 1 40
2 68660 1 40
2 68661 1 40
2 68662 1 40
2 68663 1 40
2 68664 1 40
2 68665 1 40
2 68666 1 40
2 68667 1 40
2 68668 1 40
2 68669 1 40
2 68670 1 40
2 68671 1 40
2 68672 1 40
2 68673 1 40
2 68674 1 40
2 68675 1 40
2 68676 1 40
2 68677 1 40
2 68678 1 40
2 68679 1 40
2 68680 1 40
2 68681 1 40
2 68682 1 40
2 68683 1 40
2 68684 1 40
2 68685 1 40
2 68686 1 40
2 68687 1 40
2 68688 1 40
2 68689 1 40
2 68690 1 40
2 68691 1 40
2 68692 1 40
2 68693 1 40
2 68694 1 40
2 68695 1 40
2 68696 1 40
2 68697 1 40
2 68698 1 40
2 68699 1 40
2 68700 1 40
2 68701 1 40
2 68702 1 40
2 68703 1 40
2 68704 1 40
2 68705 1 40
2 68706 1 40
2 68707 1 40
2 68708 1 40
2 68709 1 40
2 68710 1 40
2 68711 1 40
2 68712 1 40
2 68713 1 40
2 68714 1 40
2 68715 1 40
2 68716 1 40
2 68717 1 40
2 68718 1 40
2 68719 1 40
2 68720 1 40
2 68721 1 40
2 68722 1 40
2 68723 1 40
2 68724 1 40
2 68725 1 40
2 68726 1 40
2 68727 1 40
2 68728 1 40
2 68729 1 40
2 68730 1 40
2 68731 1 40
2 68732 1 40
2 68733 1 41
2 68734 1 41
2 68735 1 41
2 68736 1 41
2 68737 1 41
2 68738 1 41
2 68739 1 41
2 68740 1 41
2 68741 1 41
2 68742 1 41
2 68743 1 41
2 68744 1 41
2 68745 1 41
2 68746 1 41
2 68747 1 41
2 68748 1 41
2 68749 1 41
2 68750 1 41
2 68751 1 41
2 68752 1 41
2 68753 1 41
2 68754 1 41
2 68755 1 41
2 68756 1 41
2 68757 1 41
2 68758 1 41
2 68759 1 41
2 68760 1 41
2 68761 1 41
2 68762 1 41
2 68763 1 41
2 68764 1 41
2 68765 1 41
2 68766 1 41
2 68767 1 41
2 68768 1 41
2 68769 1 41
2 68770 1 41
2 68771 1 41
2 68772 1 41
2 68773 1 41
2 68774 1 41
2 68775 1 41
2 68776 1 41
2 68777 1 41
2 68778 1 41
2 68779 1 41
2 68780 1 41
2 68781 1 41
2 68782 1 41
2 68783 1 41
2 68784 1 41
2 68785 1 41
2 68786 1 41
2 68787 1 41
2 68788 1 41
2 68789 1 41
2 68790 1 41
2 68791 1 41
2 68792 1 41
2 68793 1 41
2 68794 1 41
2 68795 1 41
2 68796 1 41
2 68797 1 41
2 68798 1 41
2 68799 1 41
2 68800 1 41
2 68801 1 41
2 68802 1 41
2 68803 1 41
2 68804 1 41
2 68805 1 41
2 68806 1 41
2 68807 1 41
2 68808 1 41
2 68809 1 41
2 68810 1 41
2 68811 1 41
2 68812 1 41
2 68813 1 41
2 68814 1 41
2 68815 1 41
2 68816 1 41
2 68817 1 41
2 68818 1 41
2 68819 1 41
2 68820 1 41
2 68821 1 41
2 68822 1 41
2 68823 1 41
2 68824 1 41
2 68825 1 41
2 68826 1 41
2 68827 1 41
2 68828 1 41
2 68829 1 41
2 68830 1 41
2 68831 1 41
2 68832 1 41
2 68833 1 41
2 68834 1 41
2 68835 1 41
2 68836 1 41
2 68837 1 41
2 68838 1 41
2 68839 1 41
2 68840 1 41
2 68841 1 41
2 68842 1 41
2 68843 1 41
2 68844 1 41
2 68845 1 41
2 68846 1 41
2 68847 1 41
2 68848 1 41
2 68849 1 41
2 68850 1 41
2 68851 1 41
2 68852 1 41
2 68853 1 41
2 68854 1 41
2 68855 1 41
2 68856 1 41
2 68857 1 41
2 68858 1 41
2 68859 1 41
2 68860 1 41
2 68861 1 41
2 68862 1 41
2 68863 1 41
2 68864 1 41
2 68865 1 41
2 68866 1 41
2 68867 1 41
2 68868 1 41
2 68869 1 41
2 68870 1 41
2 68871 1 41
2 68872 1 41
2 68873 1 41
2 68874 1 41
2 68875 1 41
2 68876 1 41
2 68877 1 41
2 68878 1 41
2 68879 1 41
2 68880 1 41
2 68881 1 41
2 68882 1 41
2 68883 1 41
2 68884 1 41
2 68885 1 41
2 68886 1 41
2 68887 1 41
2 68888 1 42
2 68889 1 42
2 68890 1 42
2 68891 1 42
2 68892 1 42
2 68893 1 42
2 68894 1 42
2 68895 1 42
2 68896 1 42
2 68897 1 42
2 68898 1 42
2 68899 1 42
2 68900 1 42
2 68901 1 42
2 68902 1 42
2 68903 1 42
2 68904 1 42
2 68905 1 42
2 68906 1 42
2 68907 1 42
2 68908 1 42
2 68909 1 42
2 68910 1 42
2 68911 1 42
2 68912 1 42
2 68913 1 42
2 68914 1 42
2 68915 1 42
2 68916 1 42
2 68917 1 42
2 68918 1 42
2 68919 1 42
2 68920 1 42
2 68921 1 42
2 68922 1 42
2 68923 1 42
2 68924 1 42
2 68925 1 42
2 68926 1 42
2 68927 1 42
2 68928 1 42
2 68929 1 42
2 68930 1 42
2 68931 1 42
2 68932 1 42
2 68933 1 42
2 68934 1 42
2 68935 1 42
2 68936 1 42
2 68937 1 42
2 68938 1 42
2 68939 1 42
2 68940 1 42
2 68941 1 42
2 68942 1 42
2 68943 1 42
2 68944 1 42
2 68945 1 42
2 68946 1 42
2 68947 1 42
2 68948 1 42
2 68949 1 42
2 68950 1 42
2 68951 1 42
2 68952 1 42
2 68953 1 42
2 68954 1 42
2 68955 1 42
2 68956 1 42
2 68957 1 42
2 68958 1 42
2 68959 1 42
2 68960 1 42
2 68961 1 42
2 68962 1 42
2 68963 1 42
2 68964 1 42
2 68965 1 42
2 68966 1 42
2 68967 1 42
2 68968 1 42
2 68969 1 42
2 68970 1 42
2 68971 1 42
2 68972 1 42
2 68973 1 42
2 68974 1 42
2 68975 1 42
2 68976 1 42
2 68977 1 42
2 68978 1 42
2 68979 1 42
2 68980 1 42
2 68981 1 42
2 68982 1 42
2 68983 1 42
2 68984 1 42
2 68985 1 42
2 68986 1 42
2 68987 1 42
2 68988 1 42
2 68989 1 42
2 68990 1 42
2 68991 1 42
2 68992 1 42
2 68993 1 42
2 68994 1 42
2 68995 1 42
2 68996 1 42
2 68997 1 42
2 68998 1 42
2 68999 1 42
2 69000 1 42
2 69001 1 42
2 69002 1 42
2 69003 1 42
2 69004 1 42
2 69005 1 42
2 69006 1 42
2 69007 1 42
2 69008 1 42
2 69009 1 42
2 69010 1 42
2 69011 1 42
2 69012 1 42
2 69013 1 42
2 69014 1 42
2 69015 1 42
2 69016 1 42
2 69017 1 42
2 69018 1 42
2 69019 1 42
2 69020 1 42
2 69021 1 42
2 69022 1 42
2 69023 1 42
2 69024 1 42
2 69025 1 42
2 69026 1 42
2 69027 1 42
2 69028 1 42
2 69029 1 42
2 69030 1 42
2 69031 1 42
2 69032 1 42
2 69033 1 42
2 69034 1 42
2 69035 1 42
2 69036 1 42
2 69037 1 42
2 69038 1 42
2 69039 1 42
2 69040 1 42
2 69041 1 42
2 69042 1 42
2 69043 1 42
2 69044 1 42
2 69045 1 42
2 69046 1 42
2 69047 1 42
2 69048 1 42
2 69049 1 42
2 69050 1 42
2 69051 1 42
2 69052 1 42
2 69053 1 42
2 69054 1 42
2 69055 1 42
2 69056 1 42
2 69057 1 42
2 69058 1 42
2 69059 1 42
2 69060 1 42
2 69061 1 42
2 69062 1 42
2 69063 1 42
2 69064 1 42
2 69065 1 42
2 69066 1 42
2 69067 1 42
2 69068 1 42
2 69069 1 42
2 69070 1 42
2 69071 1 42
2 69072 1 42
2 69073 1 42
2 69074 1 42
2 69075 1 42
2 69076 1 42
2 69077 1 42
2 69078 1 42
2 69079 1 42
2 69080 1 42
2 69081 1 42
2 69082 1 42
2 69083 1 42
2 69084 1 43
2 69085 1 43
2 69086 1 43
2 69087 1 43
2 69088 1 43
2 69089 1 43
2 69090 1 43
2 69091 1 43
2 69092 1 43
2 69093 1 43
2 69094 1 43
2 69095 1 43
2 69096 1 43
2 69097 1 43
2 69098 1 43
2 69099 1 43
2 69100 1 43
2 69101 1 43
2 69102 1 43
2 69103 1 43
2 69104 1 43
2 69105 1 43
2 69106 1 43
2 69107 1 43
2 69108 1 43
2 69109 1 43
2 69110 1 43
2 69111 1 43
2 69112 1 43
2 69113 1 43
2 69114 1 43
2 69115 1 43
2 69116 1 43
2 69117 1 43
2 69118 1 43
2 69119 1 43
2 69120 1 43
2 69121 1 43
2 69122 1 43
2 69123 1 43
2 69124 1 43
2 69125 1 43
2 69126 1 43
2 69127 1 43
2 69128 1 43
2 69129 1 43
2 69130 1 43
2 69131 1 43
2 69132 1 43
2 69133 1 43
2 69134 1 43
2 69135 1 43
2 69136 1 43
2 69137 1 43
2 69138 1 43
2 69139 1 43
2 69140 1 43
2 69141 1 43
2 69142 1 43
2 69143 1 43
2 69144 1 43
2 69145 1 43
2 69146 1 43
2 69147 1 43
2 69148 1 43
2 69149 1 43
2 69150 1 43
2 69151 1 43
2 69152 1 43
2 69153 1 43
2 69154 1 43
2 69155 1 43
2 69156 1 44
2 69157 1 44
2 69158 1 44
2 69159 1 44
2 69160 1 44
2 69161 1 44
2 69162 1 44
2 69163 1 44
2 69164 1 44
2 69165 1 44
2 69166 1 44
2 69167 1 44
2 69168 1 44
2 69169 1 44
2 69170 1 44
2 69171 1 44
2 69172 1 44
2 69173 1 44
2 69174 1 44
2 69175 1 44
2 69176 1 44
2 69177 1 44
2 69178 1 44
2 69179 1 44
2 69180 1 44
2 69181 1 44
2 69182 1 44
2 69183 1 44
2 69184 1 44
2 69185 1 44
2 69186 1 44
2 69187 1 44
2 69188 1 44
2 69189 1 44
2 69190 1 44
2 69191 1 44
2 69192 1 44
2 69193 1 44
2 69194 1 44
2 69195 1 44
2 69196 1 44
2 69197 1 44
2 69198 1 44
2 69199 1 44
2 69200 1 44
2 69201 1 44
2 69202 1 44
2 69203 1 44
2 69204 1 44
2 69205 1 44
2 69206 1 44
2 69207 1 44
2 69208 1 44
2 69209 1 44
2 69210 1 44
2 69211 1 44
2 69212 1 44
2 69213 1 44
2 69214 1 44
2 69215 1 44
2 69216 1 44
2 69217 1 44
2 69218 1 44
2 69219 1 44
2 69220 1 44
2 69221 1 44
2 69222 1 44
2 69223 1 44
2 69224 1 44
2 69225 1 44
2 69226 1 44
2 69227 1 44
2 69228 1 44
2 69229 1 44
2 69230 1 44
2 69231 1 44
2 69232 1 44
2 69233 1 44
2 69234 1 44
2 69235 1 44
2 69236 1 44
2 69237 1 44
2 69238 1 44
2 69239 1 44
2 69240 1 44
2 69241 1 44
2 69242 1 44
2 69243 1 44
2 69244 1 44
2 69245 1 44
2 69246 1 44
2 69247 1 44
2 69248 1 44
2 69249 1 44
2 69250 1 44
2 69251 1 44
2 69252 1 44
2 69253 1 44
2 69254 1 44
2 69255 1 44
2 69256 1 44
2 69257 1 44
2 69258 1 44
2 69259 1 44
2 69260 1 44
2 69261 1 44
2 69262 1 44
2 69263 1 44
2 69264 1 44
2 69265 1 44
2 69266 1 44
2 69267 1 44
2 69268 1 44
2 69269 1 44
2 69270 1 44
2 69271 1 44
2 69272 1 44
2 69273 1 44
2 69274 1 44
2 69275 1 44
2 69276 1 45
2 69277 1 45
2 69278 1 45
2 69279 1 45
2 69280 1 45
2 69281 1 45
2 69282 1 45
2 69283 1 45
2 69284 1 45
2 69285 1 45
2 69286 1 45
2 69287 1 45
2 69288 1 45
2 69289 1 45
2 69290 1 45
2 69291 1 45
2 69292 1 45
2 69293 1 45
2 69294 1 45
2 69295 1 45
2 69296 1 45
2 69297 1 45
2 69298 1 45
2 69299 1 45
2 69300 1 45
2 69301 1 45
2 69302 1 45
2 69303 1 45
2 69304 1 45
2 69305 1 45
2 69306 1 45
2 69307 1 45
2 69308 1 45
2 69309 1 45
2 69310 1 45
2 69311 1 45
2 69312 1 45
2 69313 1 45
2 69314 1 45
2 69315 1 45
2 69316 1 45
2 69317 1 45
2 69318 1 45
2 69319 1 45
2 69320 1 45
2 69321 1 45
2 69322 1 45
2 69323 1 45
2 69324 1 45
2 69325 1 45
2 69326 1 45
2 69327 1 45
2 69328 1 45
2 69329 1 45
2 69330 1 45
2 69331 1 45
2 69332 1 45
2 69333 1 45
2 69334 1 45
2 69335 1 45
2 69336 1 45
2 69337 1 45
2 69338 1 45
2 69339 1 45
2 69340 1 45
2 69341 1 45
2 69342 1 45
2 69343 1 45
2 69344 1 45
2 69345 1 45
2 69346 1 45
2 69347 1 45
2 69348 1 45
2 69349 1 45
2 69350 1 45
2 69351 1 45
2 69352 1 45
2 69353 1 45
2 69354 1 45
2 69355 1 45
2 69356 1 45
2 69357 1 45
2 69358 1 45
2 69359 1 45
2 69360 1 45
2 69361 1 45
2 69362 1 45
2 69363 1 45
2 69364 1 45
2 69365 1 45
2 69366 1 45
2 69367 1 45
2 69368 1 45
2 69369 1 45
2 69370 1 45
2 69371 1 45
2 69372 1 45
2 69373 1 45
2 69374 1 45
2 69375 1 45
2 69376 1 45
2 69377 1 45
2 69378 1 45
2 69379 1 45
2 69380 1 45
2 69381 1 45
2 69382 1 45
2 69383 1 45
2 69384 1 45
2 69385 1 45
2 69386 1 45
2 69387 1 45
2 69388 1 45
2 69389 1 45
2 69390 1 45
2 69391 1 45
2 69392 1 45
2 69393 1 45
2 69394 1 45
2 69395 1 45
2 69396 1 45
2 69397 1 45
2 69398 1 45
2 69399 1 45
2 69400 1 45
2 69401 1 45
2 69402 1 45
2 69403 1 45
2 69404 1 45
2 69405 1 45
2 69406 1 45
2 69407 1 45
2 69408 1 45
2 69409 1 45
2 69410 1 45
2 69411 1 45
2 69412 1 45
2 69413 1 45
2 69414 1 45
2 69415 1 45
2 69416 1 45
2 69417 1 45
2 69418 1 45
2 69419 1 45
2 69420 1 45
2 69421 1 45
2 69422 1 45
2 69423 1 45
2 69424 1 45
2 69425 1 45
2 69426 1 45
2 69427 1 45
2 69428 1 45
2 69429 1 45
2 69430 1 45
2 69431 1 45
2 69432 1 45
2 69433 1 45
2 69434 1 45
2 69435 1 45
2 69436 1 45
2 69437 1 45
2 69438 1 45
2 69439 1 45
2 69440 1 45
2 69441 1 45
2 69442 1 45
2 69443 1 45
2 69444 1 45
2 69445 1 45
2 69446 1 45
2 69447 1 45
2 69448 1 45
2 69449 1 45
2 69450 1 45
2 69451 1 45
2 69452 1 45
2 69453 1 45
2 69454 1 45
2 69455 1 45
2 69456 1 45
2 69457 1 45
2 69458 1 45
2 69459 1 45
2 69460 1 46
2 69461 1 46
2 69462 1 46
2 69463 1 46
2 69464 1 46
2 69465 1 46
2 69466 1 46
2 69467 1 46
2 69468 1 46
2 69469 1 46
2 69470 1 46
2 69471 1 46
2 69472 1 46
2 69473 1 46
2 69474 1 46
2 69475 1 46
2 69476 1 46
2 69477 1 46
2 69478 1 46
2 69479 1 46
2 69480 1 46
2 69481 1 46
2 69482 1 46
2 69483 1 46
2 69484 1 46
2 69485 1 46
2 69486 1 46
2 69487 1 46
2 69488 1 46
2 69489 1 46
2 69490 1 46
2 69491 1 46
2 69492 1 46
2 69493 1 46
2 69494 1 46
2 69495 1 46
2 69496 1 46
2 69497 1 46
2 69498 1 46
2 69499 1 46
2 69500 1 46
2 69501 1 46
2 69502 1 46
2 69503 1 46
2 69504 1 46
2 69505 1 46
2 69506 1 46
2 69507 1 46
2 69508 1 46
2 69509 1 46
2 69510 1 46
2 69511 1 46
2 69512 1 46
2 69513 1 46
2 69514 1 46
2 69515 1 46
2 69516 1 46
2 69517 1 46
2 69518 1 46
2 69519 1 46
2 69520 1 46
2 69521 1 46
2 69522 1 46
2 69523 1 46
2 69524 1 46
2 69525 1 46
2 69526 1 46
2 69527 1 46
2 69528 1 46
2 69529 1 46
2 69530 1 46
2 69531 1 46
2 69532 1 46
2 69533 1 46
2 69534 1 46
2 69535 1 46
2 69536 1 46
2 69537 1 46
2 69538 1 46
2 69539 1 46
2 69540 1 46
2 69541 1 46
2 69542 1 46
2 69543 1 46
2 69544 1 46
2 69545 1 46
2 69546 1 46
2 69547 1 46
2 69548 1 46
2 69549 1 46
2 69550 1 46
2 69551 1 46
2 69552 1 46
2 69553 1 46
2 69554 1 46
2 69555 1 46
2 69556 1 46
2 69557 1 46
2 69558 1 46
2 69559 1 46
2 69560 1 46
2 69561 1 46
2 69562 1 46
2 69563 1 46
2 69564 1 46
2 69565 1 46
2 69566 1 46
2 69567 1 46
2 69568 1 46
2 69569 1 46
2 69570 1 46
2 69571 1 46
2 69572 1 46
2 69573 1 46
2 69574 1 46
2 69575 1 46
2 69576 1 46
2 69577 1 46
2 69578 1 46
2 69579 1 46
2 69580 1 46
2 69581 1 46
2 69582 1 46
2 69583 1 46
2 69584 1 46
2 69585 1 46
2 69586 1 46
2 69587 1 46
2 69588 1 46
2 69589 1 46
2 69590 1 46
2 69591 1 46
2 69592 1 46
2 69593 1 46
2 69594 1 46
2 69595 1 46
2 69596 1 46
2 69597 1 46
2 69598 1 46
2 69599 1 46
2 69600 1 46
2 69601 1 46
2 69602 1 46
2 69603 1 46
2 69604 1 46
2 69605 1 46
2 69606 1 46
2 69607 1 46
2 69608 1 46
2 69609 1 46
2 69610 1 46
2 69611 1 46
2 69612 1 46
2 69613 1 46
2 69614 1 46
2 69615 1 46
2 69616 1 46
2 69617 1 46
2 69618 1 46
2 69619 1 46
2 69620 1 46
2 69621 1 46
2 69622 1 46
2 69623 1 46
2 69624 1 46
2 69625 1 46
2 69626 1 46
2 69627 1 46
2 69628 1 46
2 69629 1 46
2 69630 1 46
2 69631 1 46
2 69632 1 46
2 69633 1 46
2 69634 1 46
2 69635 1 46
2 69636 1 46
2 69637 1 46
2 69638 1 46
2 69639 1 46
2 69640 1 46
2 69641 1 46
2 69642 1 46
2 69643 1 46
2 69644 1 46
2 69645 1 46
2 69646 1 46
2 69647 1 46
2 69648 1 46
2 69649 1 46
2 69650 1 46
2 69651 1 46
2 69652 1 46
2 69653 1 46
2 69654 1 46
2 69655 1 47
2 69656 1 47
2 69657 1 47
2 69658 1 47
2 69659 1 47
2 69660 1 47
2 69661 1 47
2 69662 1 47
2 69663 1 47
2 69664 1 47
2 69665 1 47
2 69666 1 47
2 69667 1 47
2 69668 1 47
2 69669 1 47
2 69670 1 47
2 69671 1 47
2 69672 1 47
2 69673 1 47
2 69674 1 47
2 69675 1 47
2 69676 1 47
2 69677 1 47
2 69678 1 47
2 69679 1 47
2 69680 1 47
2 69681 1 47
2 69682 1 47
2 69683 1 47
2 69684 1 47
2 69685 1 47
2 69686 1 47
2 69687 1 47
2 69688 1 47
2 69689 1 47
2 69690 1 47
2 69691 1 47
2 69692 1 47
2 69693 1 47
2 69694 1 47
2 69695 1 47
2 69696 1 47
2 69697 1 47
2 69698 1 47
2 69699 1 47
2 69700 1 47
2 69701 1 47
2 69702 1 47
2 69703 1 47
2 69704 1 47
2 69705 1 47
2 69706 1 47
2 69707 1 47
2 69708 1 47
2 69709 1 47
2 69710 1 47
2 69711 1 47
2 69712 1 47
2 69713 1 47
2 69714 1 47
2 69715 1 47
2 69716 1 47
2 69717 1 47
2 69718 1 47
2 69719 1 47
2 69720 1 47
2 69721 1 47
2 69722 1 47
2 69723 1 47
2 69724 1 47
2 69725 1 47
2 69726 1 47
2 69727 1 47
2 69728 1 47
2 69729 1 47
2 69730 1 47
2 69731 1 47
2 69732 1 47
2 69733 1 47
2 69734 1 47
2 69735 1 47
2 69736 1 47
2 69737 1 47
2 69738 1 47
2 69739 1 47
2 69740 1 47
2 69741 1 47
2 69742 1 47
2 69743 1 47
2 69744 1 47
2 69745 1 47
2 69746 1 47
2 69747 1 47
2 69748 1 47
2 69749 1 47
2 69750 1 47
2 69751 1 47
2 69752 1 47
2 69753 1 47
2 69754 1 47
2 69755 1 47
2 69756 1 47
2 69757 1 47
2 69758 1 47
2 69759 1 47
2 69760 1 47
2 69761 1 47
2 69762 1 47
2 69763 1 47
2 69764 1 47
2 69765 1 47
2 69766 1 47
2 69767 1 47
2 69768 1 47
2 69769 1 47
2 69770 1 47
2 69771 1 47
2 69772 1 47
2 69773 1 47
2 69774 1 47
2 69775 1 47
2 69776 1 47
2 69777 1 47
2 69778 1 47
2 69779 1 47
2 69780 1 47
2 69781 1 47
2 69782 1 47
2 69783 1 47
2 69784 1 47
2 69785 1 47
2 69786 1 47
2 69787 1 47
2 69788 1 47
2 69789 1 47
2 69790 1 47
2 69791 1 47
2 69792 1 47
2 69793 1 47
2 69794 1 47
2 69795 1 47
2 69796 1 47
2 69797 1 47
2 69798 1 47
2 69799 1 47
2 69800 1 47
2 69801 1 47
2 69802 1 47
2 69803 1 47
2 69804 1 47
2 69805 1 47
2 69806 1 47
2 69807 1 47
2 69808 1 47
2 69809 1 47
2 69810 1 47
2 69811 1 47
2 69812 1 47
2 69813 1 47
2 69814 1 47
2 69815 1 47
2 69816 1 47
2 69817 1 47
2 69818 1 47
2 69819 1 47
2 69820 1 47
2 69821 1 47
2 69822 1 47
2 69823 1 47
2 69824 1 47
2 69825 1 47
2 69826 1 47
2 69827 1 47
2 69828 1 47
2 69829 1 47
2 69830 1 47
2 69831 1 47
2 69832 1 47
2 69833 1 47
2 69834 1 47
2 69835 1 47
2 69836 1 47
2 69837 1 47
2 69838 1 47
2 69839 1 47
2 69840 1 47
2 69841 1 47
2 69842 1 47
2 69843 1 47
2 69844 1 47
2 69845 1 47
2 69846 1 47
2 69847 1 47
2 69848 1 47
2 69849 1 47
2 69850 1 47
2 69851 1 47
2 69852 1 47
2 69853 1 47
2 69854 1 47
2 69855 1 47
2 69856 1 47
2 69857 1 47
2 69858 1 47
2 69859 1 47
2 69860 1 47
2 69861 1 47
2 69862 1 47
2 69863 1 47
2 69864 1 47
2 69865 1 47
2 69866 1 47
2 69867 1 47
2 69868 1 47
2 69869 1 47
2 69870 1 47
2 69871 1 47
2 69872 1 47
2 69873 1 47
2 69874 1 47
2 69875 1 47
2 69876 1 48
2 69877 1 48
2 69878 1 48
2 69879 1 48
2 69880 1 48
2 69881 1 48
2 69882 1 48
2 69883 1 48
2 69884 1 48
2 69885 1 48
2 69886 1 48
2 69887 1 48
2 69888 1 48
2 69889 1 48
2 69890 1 48
2 69891 1 48
2 69892 1 48
2 69893 1 48
2 69894 1 48
2 69895 1 48
2 69896 1 48
2 69897 1 48
2 69898 1 48
2 69899 1 48
2 69900 1 48
2 69901 1 48
2 69902 1 48
2 69903 1 48
2 69904 1 48
2 69905 1 48
2 69906 1 48
2 69907 1 48
2 69908 1 48
2 69909 1 48
2 69910 1 48
2 69911 1 48
2 69912 1 48
2 69913 1 48
2 69914 1 48
2 69915 1 48
2 69916 1 48
2 69917 1 48
2 69918 1 48
2 69919 1 48
2 69920 1 48
2 69921 1 48
2 69922 1 48
2 69923 1 48
2 69924 1 48
2 69925 1 48
2 69926 1 48
2 69927 1 48
2 69928 1 48
2 69929 1 48
2 69930 1 48
2 69931 1 48
2 69932 1 48
2 69933 1 48
2 69934 1 48
2 69935 1 48
2 69936 1 48
2 69937 1 48
2 69938 1 48
2 69939 1 48
2 69940 1 48
2 69941 1 48
2 69942 1 48
2 69943 1 48
2 69944 1 48
2 69945 1 48
2 69946 1 48
2 69947 1 48
2 69948 1 48
2 69949 1 48
2 69950 1 48
2 69951 1 48
2 69952 1 48
2 69953 1 48
2 69954 1 48
2 69955 1 48
2 69956 1 48
2 69957 1 48
2 69958 1 48
2 69959 1 48
2 69960 1 48
2 69961 1 48
2 69962 1 48
2 69963 1 48
2 69964 1 48
2 69965 1 48
2 69966 1 48
2 69967 1 48
2 69968 1 48
2 69969 1 48
2 69970 1 48
2 69971 1 48
2 69972 1 48
2 69973 1 48
2 69974 1 48
2 69975 1 48
2 69976 1 48
2 69977 1 48
2 69978 1 48
2 69979 1 48
2 69980 1 48
2 69981 1 48
2 69982 1 48
2 69983 1 48
2 69984 1 48
2 69985 1 48
2 69986 1 48
2 69987 1 48
2 69988 1 48
2 69989 1 48
2 69990 1 48
2 69991 1 48
2 69992 1 48
2 69993 1 48
2 69994 1 48
2 69995 1 48
2 69996 1 48
2 69997 1 48
2 69998 1 48
2 69999 1 48
2 70000 1 48
2 70001 1 48
2 70002 1 48
2 70003 1 48
2 70004 1 48
2 70005 1 48
2 70006 1 48
2 70007 1 48
2 70008 1 48
2 70009 1 48
2 70010 1 48
2 70011 1 48
2 70012 1 48
2 70013 1 48
2 70014 1 48
2 70015 1 48
2 70016 1 48
2 70017 1 48
2 70018 1 48
2 70019 1 48
2 70020 1 48
2 70021 1 48
2 70022 1 48
2 70023 1 48
2 70024 1 48
2 70025 1 48
2 70026 1 48
2 70027 1 48
2 70028 1 48
2 70029 1 48
2 70030 1 48
2 70031 1 48
2 70032 1 48
2 70033 1 48
2 70034 1 48
2 70035 1 48
2 70036 1 48
2 70037 1 48
2 70038 1 48
2 70039 1 48
2 70040 1 48
2 70041 1 48
2 70042 1 48
2 70043 1 48
2 70044 1 48
2 70045 1 48
2 70046 1 48
2 70047 1 48
2 70048 1 48
2 70049 1 48
2 70050 1 48
2 70051 1 48
2 70052 1 48
2 70053 1 48
2 70054 1 48
2 70055 1 48
2 70056 1 48
2 70057 1 48
2 70058 1 48
2 70059 1 48
2 70060 1 48
2 70061 1 48
2 70062 1 48
2 70063 1 48
2 70064 1 48
2 70065 1 48
2 70066 1 48
2 70067 1 48
2 70068 1 48
2 70069 1 48
2 70070 1 48
2 70071 1 48
2 70072 1 48
2 70073 1 48
2 70074 1 48
2 70075 1 48
2 70076 1 48
2 70077 1 48
2 70078 1 48
2 70079 1 48
2 70080 1 48
2 70081 1 48
2 70082 1 48
2 70083 1 48
2 70084 1 48
2 70085 1 48
2 70086 1 48
2 70087 1 48
2 70088 1 48
2 70089 1 48
2 70090 1 48
2 70091 1 48
2 70092 1 48
2 70093 1 48
2 70094 1 48
2 70095 1 48
2 70096 1 48
2 70097 1 48
2 70098 1 48
2 70099 1 48
2 70100 1 48
2 70101 1 48
2 70102 1 48
2 70103 1 48
2 70104 1 48
2 70105 1 48
2 70106 1 48
2 70107 1 48
2 70108 1 48
2 70109 1 48
2 70110 1 48
2 70111 1 48
2 70112 1 48
2 70113 1 48
2 70114 1 48
2 70115 1 48
2 70116 1 48
2 70117 1 48
2 70118 1 48
2 70119 1 48
2 70120 1 48
2 70121 1 48
2 70122 1 48
2 70123 1 48
2 70124 1 48
2 70125 1 48
2 70126 1 48
2 70127 1 48
2 70128 1 48
2 70129 1 48
2 70130 1 48
2 70131 1 48
2 70132 1 48
2 70133 1 48
2 70134 1 48
2 70135 1 48
2 70136 1 48
2 70137 1 48
2 70138 1 48
2 70139 1 48
2 70140 1 48
2 70141 1 48
2 70142 1 48
2 70143 1 48
2 70144 1 48
2 70145 1 48
2 70146 1 48
2 70147 1 48
2 70148 1 48
2 70149 1 48
2 70150 1 48
2 70151 1 48
2 70152 1 48
2 70153 1 48
2 70154 1 48
2 70155 1 48
2 70156 1 48
2 70157 1 48
2 70158 1 48
2 70159 1 48
2 70160 1 48
2 70161 1 48
2 70162 1 48
2 70163 1 48
2 70164 1 48
2 70165 1 48
2 70166 1 48
2 70167 1 48
2 70168 1 48
2 70169 1 48
2 70170 1 48
2 70171 1 48
2 70172 1 48
2 70173 1 48
2 70174 1 48
2 70175 1 48
2 70176 1 48
2 70177 1 48
2 70178 1 48
2 70179 1 48
2 70180 1 48
2 70181 1 48
2 70182 1 49
2 70183 1 49
2 70184 1 49
2 70185 1 49
2 70186 1 49
2 70187 1 49
2 70188 1 49
2 70189 1 49
2 70190 1 49
2 70191 1 49
2 70192 1 49
2 70193 1 49
2 70194 1 49
2 70195 1 49
2 70196 1 49
2 70197 1 49
2 70198 1 49
2 70199 1 49
2 70200 1 49
2 70201 1 49
2 70202 1 49
2 70203 1 49
2 70204 1 49
2 70205 1 49
2 70206 1 49
2 70207 1 49
2 70208 1 49
2 70209 1 49
2 70210 1 49
2 70211 1 49
2 70212 1 49
2 70213 1 49
2 70214 1 49
2 70215 1 49
2 70216 1 49
2 70217 1 49
2 70218 1 49
2 70219 1 49
2 70220 1 49
2 70221 1 49
2 70222 1 49
2 70223 1 49
2 70224 1 49
2 70225 1 49
2 70226 1 49
2 70227 1 49
2 70228 1 49
2 70229 1 49
2 70230 1 49
2 70231 1 49
2 70232 1 49
2 70233 1 49
2 70234 1 49
2 70235 1 49
2 70236 1 49
2 70237 1 49
2 70238 1 49
2 70239 1 49
2 70240 1 49
2 70241 1 49
2 70242 1 49
2 70243 1 49
2 70244 1 49
2 70245 1 49
2 70246 1 49
2 70247 1 49
2 70248 1 49
2 70249 1 49
2 70250 1 49
2 70251 1 49
2 70252 1 49
2 70253 1 49
2 70254 1 49
2 70255 1 49
2 70256 1 49
2 70257 1 49
2 70258 1 49
2 70259 1 49
2 70260 1 49
2 70261 1 49
2 70262 1 49
2 70263 1 49
2 70264 1 49
2 70265 1 49
2 70266 1 49
2 70267 1 49
2 70268 1 49
2 70269 1 49
2 70270 1 49
2 70271 1 49
2 70272 1 49
2 70273 1 49
2 70274 1 49
2 70275 1 49
2 70276 1 49
2 70277 1 49
2 70278 1 49
2 70279 1 49
2 70280 1 49
2 70281 1 49
2 70282 1 49
2 70283 1 49
2 70284 1 49
2 70285 1 49
2 70286 1 49
2 70287 1 49
2 70288 1 49
2 70289 1 49
2 70290 1 49
2 70291 1 49
2 70292 1 49
2 70293 1 49
2 70294 1 49
2 70295 1 49
2 70296 1 49
2 70297 1 49
2 70298 1 49
2 70299 1 49
2 70300 1 49
2 70301 1 49
2 70302 1 49
2 70303 1 49
2 70304 1 49
2 70305 1 49
2 70306 1 49
2 70307 1 49
2 70308 1 49
2 70309 1 49
2 70310 1 49
2 70311 1 49
2 70312 1 49
2 70313 1 49
2 70314 1 49
2 70315 1 49
2 70316 1 49
2 70317 1 49
2 70318 1 49
2 70319 1 49
2 70320 1 49
2 70321 1 49
2 70322 1 49
2 70323 1 49
2 70324 1 49
2 70325 1 49
2 70326 1 49
2 70327 1 49
2 70328 1 49
2 70329 1 49
2 70330 1 49
2 70331 1 49
2 70332 1 49
2 70333 1 49
2 70334 1 49
2 70335 1 49
2 70336 1 49
2 70337 1 49
2 70338 1 49
2 70339 1 49
2 70340 1 49
2 70341 1 49
2 70342 1 49
2 70343 1 49
2 70344 1 49
2 70345 1 49
2 70346 1 49
2 70347 1 49
2 70348 1 49
2 70349 1 49
2 70350 1 49
2 70351 1 49
2 70352 1 49
2 70353 1 49
2 70354 1 49
2 70355 1 49
2 70356 1 49
2 70357 1 49
2 70358 1 49
2 70359 1 49
2 70360 1 49
2 70361 1 49
2 70362 1 49
2 70363 1 49
2 70364 1 49
2 70365 1 49
2 70366 1 49
2 70367 1 49
2 70368 1 49
2 70369 1 49
2 70370 1 49
2 70371 1 49
2 70372 1 49
2 70373 1 49
2 70374 1 49
2 70375 1 49
2 70376 1 49
2 70377 1 49
2 70378 1 49
2 70379 1 49
2 70380 1 49
2 70381 1 49
2 70382 1 49
2 70383 1 49
2 70384 1 49
2 70385 1 49
2 70386 1 49
2 70387 1 49
2 70388 1 49
2 70389 1 49
2 70390 1 49
2 70391 1 49
2 70392 1 49
2 70393 1 49
2 70394 1 49
2 70395 1 49
2 70396 1 49
2 70397 1 49
2 70398 1 49
2 70399 1 49
2 70400 1 49
2 70401 1 49
2 70402 1 49
2 70403 1 49
2 70404 1 49
2 70405 1 49
2 70406 1 49
2 70407 1 49
2 70408 1 49
2 70409 1 49
2 70410 1 49
2 70411 1 49
2 70412 1 49
2 70413 1 49
2 70414 1 49
2 70415 1 49
2 70416 1 49
2 70417 1 49
2 70418 1 49
2 70419 1 49
2 70420 1 49
2 70421 1 49
2 70422 1 49
2 70423 1 49
2 70424 1 49
2 70425 1 49
2 70426 1 49
2 70427 1 49
2 70428 1 49
2 70429 1 49
2 70430 1 49
2 70431 1 49
2 70432 1 49
2 70433 1 49
2 70434 1 49
2 70435 1 49
2 70436 1 49
2 70437 1 49
2 70438 1 49
2 70439 1 49
2 70440 1 49
2 70441 1 49
2 70442 1 49
2 70443 1 49
2 70444 1 49
2 70445 1 49
2 70446 1 49
2 70447 1 49
2 70448 1 49
2 70449 1 49
2 70450 1 49
2 70451 1 49
2 70452 1 49
2 70453 1 49
2 70454 1 49
2 70455 1 49
2 70456 1 49
2 70457 1 49
2 70458 1 49
2 70459 1 49
2 70460 1 49
2 70461 1 49
2 70462 1 49
2 70463 1 49
2 70464 1 49
2 70465 1 49
2 70466 1 49
2 70467 1 49
2 70468 1 49
2 70469 1 49
2 70470 1 49
2 70471 1 49
2 70472 1 49
2 70473 1 49
2 70474 1 49
2 70475 1 49
2 70476 1 49
2 70477 1 49
2 70478 1 49
2 70479 1 49
2 70480 1 49
2 70481 1 49
2 70482 1 49
2 70483 1 49
2 70484 1 49
2 70485 1 49
2 70486 1 49
2 70487 1 49
2 70488 1 49
2 70489 1 49
2 70490 1 49
2 70491 1 49
2 70492 1 49
2 70493 1 49
2 70494 1 49
2 70495 1 49
2 70496 1 49
2 70497 1 49
2 70498 1 49
2 70499 1 49
2 70500 1 49
2 70501 1 49
2 70502 1 49
2 70503 1 49
2 70504 1 49
2 70505 1 49
2 70506 1 49
2 70507 1 49
2 70508 1 49
2 70509 1 49
2 70510 1 49
2 70511 1 49
2 70512 1 49
2 70513 1 49
2 70514 1 49
2 70515 1 49
2 70516 1 49
2 70517 1 49
2 70518 1 49
2 70519 1 49
2 70520 1 49
2 70521 1 49
2 70522 1 49
2 70523 1 49
2 70524 1 49
2 70525 1 49
2 70526 1 49
2 70527 1 49
2 70528 1 49
2 70529 1 49
2 70530 1 49
2 70531 1 49
2 70532 1 49
2 70533 1 49
2 70534 1 49
2 70535 1 49
2 70536 1 49
2 70537 1 49
2 70538 1 49
2 70539 1 49
2 70540 1 49
2 70541 1 49
2 70542 1 49
2 70543 1 49
2 70544 1 49
2 70545 1 49
2 70546 1 49
2 70547 1 49
2 70548 1 49
2 70549 1 49
2 70550 1 49
2 70551 1 49
2 70552 1 49
2 70553 1 49
2 70554 1 49
2 70555 1 49
2 70556 1 49
2 70557 1 49
2 70558 1 50
2 70559 1 50
2 70560 1 50
2 70561 1 50
2 70562 1 50
2 70563 1 50
2 70564 1 50
2 70565 1 50
2 70566 1 50
2 70567 1 50
2 70568 1 50
2 70569 1 50
2 70570 1 50
2 70571 1 50
2 70572 1 50
2 70573 1 50
2 70574 1 50
2 70575 1 50
2 70576 1 50
2 70577 1 50
2 70578 1 50
2 70579 1 50
2 70580 1 50
2 70581 1 50
2 70582 1 50
2 70583 1 50
2 70584 1 50
2 70585 1 50
2 70586 1 50
2 70587 1 50
2 70588 1 50
2 70589 1 50
2 70590 1 50
2 70591 1 50
2 70592 1 50
2 70593 1 50
2 70594 1 50
2 70595 1 50
2 70596 1 50
2 70597 1 50
2 70598 1 50
2 70599 1 50
2 70600 1 50
2 70601 1 50
2 70602 1 50
2 70603 1 50
2 70604 1 50
2 70605 1 50
2 70606 1 50
2 70607 1 50
2 70608 1 50
2 70609 1 50
2 70610 1 50
2 70611 1 50
2 70612 1 50
2 70613 1 50
2 70614 1 50
2 70615 1 50
2 70616 1 50
2 70617 1 50
2 70618 1 50
2 70619 1 50
2 70620 1 50
2 70621 1 50
2 70622 1 50
2 70623 1 50
2 70624 1 50
2 70625 1 50
2 70626 1 50
2 70627 1 50
2 70628 1 50
2 70629 1 50
2 70630 1 50
2 70631 1 50
2 70632 1 50
2 70633 1 50
2 70634 1 50
2 70635 1 50
2 70636 1 50
2 70637 1 50
2 70638 1 50
2 70639 1 50
2 70640 1 50
2 70641 1 50
2 70642 1 50
2 70643 1 50
2 70644 1 50
2 70645 1 50
2 70646 1 50
2 70647 1 50
2 70648 1 50
2 70649 1 50
2 70650 1 50
2 70651 1 50
2 70652 1 50
2 70653 1 50
2 70654 1 50
2 70655 1 50
2 70656 1 50
2 70657 1 50
2 70658 1 50
2 70659 1 50
2 70660 1 50
2 70661 1 50
2 70662 1 50
2 70663 1 50
2 70664 1 50
2 70665 1 50
2 70666 1 50
2 70667 1 50
2 70668 1 50
2 70669 1 50
2 70670 1 50
2 70671 1 50
2 70672 1 50
2 70673 1 50
2 70674 1 50
2 70675 1 50
2 70676 1 50
2 70677 1 50
2 70678 1 50
2 70679 1 50
2 70680 1 50
2 70681 1 50
2 70682 1 50
2 70683 1 50
2 70684 1 50
2 70685 1 50
2 70686 1 50
2 70687 1 50
2 70688 1 50
2 70689 1 50
2 70690 1 50
2 70691 1 50
2 70692 1 50
2 70693 1 50
2 70694 1 50
2 70695 1 50
2 70696 1 50
2 70697 1 50
2 70698 1 50
2 70699 1 50
2 70700 1 50
2 70701 1 50
2 70702 1 50
2 70703 1 50
2 70704 1 50
2 70705 1 50
2 70706 1 50
2 70707 1 50
2 70708 1 50
2 70709 1 50
2 70710 1 50
2 70711 1 50
2 70712 1 50
2 70713 1 50
2 70714 1 50
2 70715 1 50
2 70716 1 50
2 70717 1 50
2 70718 1 50
2 70719 1 50
2 70720 1 50
2 70721 1 50
2 70722 1 50
2 70723 1 50
2 70724 1 50
2 70725 1 50
2 70726 1 50
2 70727 1 50
2 70728 1 50
2 70729 1 50
2 70730 1 50
2 70731 1 50
2 70732 1 50
2 70733 1 50
2 70734 1 50
2 70735 1 50
2 70736 1 50
2 70737 1 50
2 70738 1 50
2 70739 1 50
2 70740 1 50
2 70741 1 50
2 70742 1 50
2 70743 1 50
2 70744 1 50
2 70745 1 50
2 70746 1 50
2 70747 1 50
2 70748 1 50
2 70749 1 50
2 70750 1 50
2 70751 1 50
2 70752 1 50
2 70753 1 50
2 70754 1 50
2 70755 1 50
2 70756 1 50
2 70757 1 50
2 70758 1 50
2 70759 1 50
2 70760 1 50
2 70761 1 50
2 70762 1 50
2 70763 1 50
2 70764 1 50
2 70765 1 50
2 70766 1 50
2 70767 1 50
2 70768 1 50
2 70769 1 50
2 70770 1 50
2 70771 1 50
2 70772 1 50
2 70773 1 50
2 70774 1 50
2 70775 1 50
2 70776 1 50
2 70777 1 50
2 70778 1 50
2 70779 1 50
2 70780 1 50
2 70781 1 50
2 70782 1 50
2 70783 1 50
2 70784 1 50
2 70785 1 50
2 70786 1 50
2 70787 1 50
2 70788 1 50
2 70789 1 50
2 70790 1 50
2 70791 1 50
2 70792 1 50
2 70793 1 50
2 70794 1 50
2 70795 1 50
2 70796 1 50
2 70797 1 50
2 70798 1 50
2 70799 1 50
2 70800 1 50
2 70801 1 50
2 70802 1 50
2 70803 1 50
2 70804 1 50
2 70805 1 50
2 70806 1 51
2 70807 1 51
2 70808 1 51
2 70809 1 51
2 70810 1 51
2 70811 1 51
2 70812 1 51
2 70813 1 51
2 70814 1 51
2 70815 1 51
2 70816 1 51
2 70817 1 51
2 70818 1 51
2 70819 1 51
2 70820 1 51
2 70821 1 51
2 70822 1 51
2 70823 1 51
2 70824 1 51
2 70825 1 51
2 70826 1 51
2 70827 1 51
2 70828 1 51
2 70829 1 51
2 70830 1 51
2 70831 1 51
2 70832 1 51
2 70833 1 51
2 70834 1 51
2 70835 1 51
2 70836 1 51
2 70837 1 51
2 70838 1 51
2 70839 1 51
2 70840 1 51
2 70841 1 51
2 70842 1 51
2 70843 1 51
2 70844 1 51
2 70845 1 51
2 70846 1 51
2 70847 1 51
2 70848 1 51
2 70849 1 51
2 70850 1 51
2 70851 1 51
2 70852 1 51
2 70853 1 51
2 70854 1 51
2 70855 1 51
2 70856 1 51
2 70857 1 51
2 70858 1 51
2 70859 1 51
2 70860 1 51
2 70861 1 51
2 70862 1 51
2 70863 1 51
2 70864 1 51
2 70865 1 51
2 70866 1 51
2 70867 1 51
2 70868 1 51
2 70869 1 51
2 70870 1 51
2 70871 1 51
2 70872 1 51
2 70873 1 51
2 70874 1 51
2 70875 1 51
2 70876 1 51
2 70877 1 51
2 70878 1 51
2 70879 1 51
2 70880 1 51
2 70881 1 51
2 70882 1 51
2 70883 1 51
2 70884 1 51
2 70885 1 51
2 70886 1 51
2 70887 1 51
2 70888 1 51
2 70889 1 51
2 70890 1 51
2 70891 1 51
2 70892 1 51
2 70893 1 51
2 70894 1 51
2 70895 1 51
2 70896 1 51
2 70897 1 51
2 70898 1 51
2 70899 1 51
2 70900 1 51
2 70901 1 51
2 70902 1 51
2 70903 1 51
2 70904 1 51
2 70905 1 51
2 70906 1 51
2 70907 1 51
2 70908 1 51
2 70909 1 51
2 70910 1 51
2 70911 1 51
2 70912 1 51
2 70913 1 51
2 70914 1 51
2 70915 1 51
2 70916 1 51
2 70917 1 51
2 70918 1 51
2 70919 1 51
2 70920 1 51
2 70921 1 51
2 70922 1 51
2 70923 1 51
2 70924 1 51
2 70925 1 51
2 70926 1 51
2 70927 1 51
2 70928 1 51
2 70929 1 51
2 70930 1 51
2 70931 1 51
2 70932 1 51
2 70933 1 51
2 70934 1 51
2 70935 1 51
2 70936 1 51
2 70937 1 51
2 70938 1 51
2 70939 1 51
2 70940 1 51
2 70941 1 51
2 70942 1 51
2 70943 1 51
2 70944 1 51
2 70945 1 51
2 70946 1 51
2 70947 1 51
2 70948 1 51
2 70949 1 51
2 70950 1 51
2 70951 1 51
2 70952 1 51
2 70953 1 51
2 70954 1 51
2 70955 1 51
2 70956 1 51
2 70957 1 51
2 70958 1 51
2 70959 1 51
2 70960 1 51
2 70961 1 51
2 70962 1 51
2 70963 1 51
2 70964 1 51
2 70965 1 51
2 70966 1 51
2 70967 1 51
2 70968 1 51
2 70969 1 51
2 70970 1 51
2 70971 1 51
2 70972 1 51
2 70973 1 51
2 70974 1 51
2 70975 1 51
2 70976 1 51
2 70977 1 51
2 70978 1 51
2 70979 1 51
2 70980 1 51
2 70981 1 51
2 70982 1 51
2 70983 1 51
2 70984 1 51
2 70985 1 52
2 70986 1 52
2 70987 1 52
2 70988 1 52
2 70989 1 52
2 70990 1 52
2 70991 1 52
2 70992 1 52
2 70993 1 52
2 70994 1 52
2 70995 1 52
2 70996 1 52
2 70997 1 52
2 70998 1 52
2 70999 1 52
2 71000 1 53
2 71001 1 53
2 71002 1 53
2 71003 1 53
2 71004 1 53
2 71005 1 54
2 71006 1 54
2 71007 1 55
2 71008 1 55
2 71009 1 56
2 71010 1 56
2 71011 1 56
2 71012 1 56
2 71013 1 56
2 71014 1 56
2 71015 1 56
2 71016 1 56
2 71017 1 56
2 71018 1 56
2 71019 1 56
2 71020 1 56
2 71021 1 56
2 71022 1 56
2 71023 1 57
2 71024 1 57
2 71025 1 57
2 71026 1 57
2 71027 1 57
2 71028 1 58
2 71029 1 58
2 71030 1 58
2 71031 1 58
2 71032 1 58
2 71033 1 58
2 71034 1 58
2 71035 1 58
2 71036 1 58
2 71037 1 58
2 71038 1 58
2 71039 1 58
2 71040 1 58
2 71041 1 58
2 71042 1 58
2 71043 1 58
2 71044 1 58
2 71045 1 58
2 71046 1 58
2 71047 1 58
2 71048 1 58
2 71049 1 58
2 71050 1 58
2 71051 1 58
2 71052 1 58
2 71053 1 58
2 71054 1 58
2 71055 1 58
2 71056 1 58
2 71057 1 58
2 71058 1 58
2 71059 1 58
2 71060 1 58
2 71061 1 58
2 71062 1 58
2 71063 1 58
2 71064 1 58
2 71065 1 58
2 71066 1 58
2 71067 1 58
2 71068 1 58
2 71069 1 58
2 71070 1 58
2 71071 1 58
2 71072 1 58
2 71073 1 58
2 71074 1 58
2 71075 1 58
2 71076 1 58
2 71077 1 58
2 71078 1 58
2 71079 1 58
2 71080 1 58
2 71081 1 58
2 71082 1 58
2 71083 1 58
2 71084 1 58
2 71085 1 58
2 71086 1 58
2 71087 1 58
2 71088 1 58
2 71089 1 59
2 71090 1 59
2 71091 1 59
2 71092 1 59
2 71093 1 59
2 71094 1 59
2 71095 1 59
2 71096 1 59
2 71097 1 60
2 71098 1 60
2 71099 1 63
2 71100 1 63
2 71101 1 63
2 71102 1 63
2 71103 1 63
2 71104 1 63
2 71105 1 70
2 71106 1 70
2 71107 1 70
2 71108 1 70
2 71109 1 70
2 71110 1 70
2 71111 1 70
2 71112 1 70
2 71113 1 70
2 71114 1 70
2 71115 1 70
2 71116 1 70
2 71117 1 71
2 71118 1 71
2 71119 1 72
2 71120 1 72
2 71121 1 72
2 71122 1 72
2 71123 1 72
2 71124 1 72
2 71125 1 72
2 71126 1 72
2 71127 1 72
2 71128 1 72
2 71129 1 72
2 71130 1 72
2 71131 1 72
2 71132 1 72
2 71133 1 72
2 71134 1 73
2 71135 1 73
2 71136 1 74
2 71137 1 74
2 71138 1 75
2 71139 1 75
2 71140 1 75
2 71141 1 75
2 71142 1 75
2 71143 1 75
2 71144 1 75
2 71145 1 75
2 71146 1 75
2 71147 1 75
2 71148 1 75
2 71149 1 75
2 71150 1 75
2 71151 1 75
2 71152 1 75
2 71153 1 75
2 71154 1 75
2 71155 1 75
2 71156 1 75
2 71157 1 75
2 71158 1 75
2 71159 1 75
2 71160 1 75
2 71161 1 75
2 71162 1 75
2 71163 1 75
2 71164 1 75
2 71165 1 75
2 71166 1 75
2 71167 1 75
2 71168 1 75
2 71169 1 75
2 71170 1 75
2 71171 1 75
2 71172 1 75
2 71173 1 75
2 71174 1 75
2 71175 1 75
2 71176 1 75
2 71177 1 75
2 71178 1 75
2 71179 1 75
2 71180 1 75
2 71181 1 75
2 71182 1 75
2 71183 1 75
2 71184 1 75
2 71185 1 76
2 71186 1 76
2 71187 1 76
2 71188 1 76
2 71189 1 76
2 71190 1 76
2 71191 1 76
2 71192 1 76
2 71193 1 76
2 71194 1 76
2 71195 1 76
2 71196 1 76
2 71197 1 76
2 71198 1 76
2 71199 1 76
2 71200 1 76
2 71201 1 76
2 71202 1 76
2 71203 1 76
2 71204 1 76
2 71205 1 76
2 71206 1 76
2 71207 1 76
2 71208 1 76
2 71209 1 76
2 71210 1 76
2 71211 1 76
2 71212 1 76
2 71213 1 76
2 71214 1 76
2 71215 1 76
2 71216 1 76
2 71217 1 76
2 71218 1 76
2 71219 1 76
2 71220 1 76
2 71221 1 76
2 71222 1 76
2 71223 1 76
2 71224 1 76
2 71225 1 76
2 71226 1 76
2 71227 1 76
2 71228 1 76
2 71229 1 76
2 71230 1 76
2 71231 1 76
2 71232 1 76
2 71233 1 76
2 71234 1 76
2 71235 1 76
2 71236 1 76
2 71237 1 76
2 71238 1 76
2 71239 1 76
2 71240 1 76
2 71241 1 76
2 71242 1 76
2 71243 1 76
2 71244 1 76
2 71245 1 76
2 71246 1 76
2 71247 1 76
2 71248 1 76
2 71249 1 76
2 71250 1 76
2 71251 1 76
2 71252 1 76
2 71253 1 76
2 71254 1 76
2 71255 1 76
2 71256 1 76
2 71257 1 76
2 71258 1 76
2 71259 1 76
2 71260 1 76
2 71261 1 76
2 71262 1 76
2 71263 1 76
2 71264 1 76
2 71265 1 76
2 71266 1 76
2 71267 1 76
2 71268 1 76
2 71269 1 76
2 71270 1 76
2 71271 1 76
2 71272 1 76
2 71273 1 76
2 71274 1 76
2 71275 1 76
2 71276 1 76
2 71277 1 77
2 71278 1 77
2 71279 1 77
2 71280 1 77
2 71281 1 77
2 71282 1 77
2 71283 1 77
2 71284 1 77
2 71285 1 77
2 71286 1 77
2 71287 1 77
2 71288 1 77
2 71289 1 77
2 71290 1 77
2 71291 1 77
2 71292 1 77
2 71293 1 77
2 71294 1 77
2 71295 1 77
2 71296 1 77
2 71297 1 77
2 71298 1 77
2 71299 1 77
2 71300 1 77
2 71301 1 77
2 71302 1 77
2 71303 1 77
2 71304 1 77
2 71305 1 77
2 71306 1 77
2 71307 1 77
2 71308 1 77
2 71309 1 77
2 71310 1 77
2 71311 1 77
2 71312 1 77
2 71313 1 77
2 71314 1 77
2 71315 1 77
2 71316 1 77
2 71317 1 77
2 71318 1 77
2 71319 1 77
2 71320 1 77
2 71321 1 77
2 71322 1 77
2 71323 1 77
2 71324 1 77
2 71325 1 77
2 71326 1 77
2 71327 1 77
2 71328 1 77
2 71329 1 77
2 71330 1 77
2 71331 1 77
2 71332 1 77
2 71333 1 77
2 71334 1 77
2 71335 1 77
2 71336 1 77
2 71337 1 77
2 71338 1 77
2 71339 1 77
2 71340 1 77
2 71341 1 77
2 71342 1 77
2 71343 1 77
2 71344 1 77
2 71345 1 77
2 71346 1 77
2 71347 1 77
2 71348 1 77
2 71349 1 77
2 71350 1 77
2 71351 1 77
2 71352 1 77
2 71353 1 77
2 71354 1 77
2 71355 1 77
2 71356 1 77
2 71357 1 77
2 71358 1 77
2 71359 1 77
2 71360 1 77
2 71361 1 77
2 71362 1 77
2 71363 1 77
2 71364 1 77
2 71365 1 77
2 71366 1 77
2 71367 1 77
2 71368 1 77
2 71369 1 77
2 71370 1 77
2 71371 1 77
2 71372 1 77
2 71373 1 77
2 71374 1 77
2 71375 1 77
2 71376 1 77
2 71377 1 77
2 71378 1 77
2 71379 1 77
2 71380 1 77
2 71381 1 77
2 71382 1 77
2 71383 1 77
2 71384 1 77
2 71385 1 77
2 71386 1 77
2 71387 1 77
2 71388 1 77
2 71389 1 77
2 71390 1 77
2 71391 1 77
2 71392 1 77
2 71393 1 77
2 71394 1 77
2 71395 1 77
2 71396 1 77
2 71397 1 77
2 71398 1 77
2 71399 1 77
2 71400 1 77
2 71401 1 77
2 71402 1 77
2 71403 1 77
2 71404 1 77
2 71405 1 78
2 71406 1 78
2 71407 1 78
2 71408 1 78
2 71409 1 78
2 71410 1 78
2 71411 1 78
2 71412 1 78
2 71413 1 78
2 71414 1 78
2 71415 1 78
2 71416 1 78
2 71417 1 78
2 71418 1 78
2 71419 1 78
2 71420 1 78
2 71421 1 78
2 71422 1 78
2 71423 1 78
2 71424 1 78
2 71425 1 78
2 71426 1 78
2 71427 1 78
2 71428 1 78
2 71429 1 78
2 71430 1 78
2 71431 1 78
2 71432 1 78
2 71433 1 78
2 71434 1 78
2 71435 1 78
2 71436 1 78
2 71437 1 78
2 71438 1 78
2 71439 1 78
2 71440 1 78
2 71441 1 78
2 71442 1 78
2 71443 1 78
2 71444 1 78
2 71445 1 78
2 71446 1 78
2 71447 1 78
2 71448 1 78
2 71449 1 78
2 71450 1 78
2 71451 1 78
2 71452 1 78
2 71453 1 78
2 71454 1 78
2 71455 1 78
2 71456 1 79
2 71457 1 79
2 71458 1 80
2 71459 1 80
2 71460 1 80
2 71461 1 80
2 71462 1 87
2 71463 1 87
2 71464 1 87
2 71465 1 87
2 71466 1 87
2 71467 1 87
2 71468 1 87
2 71469 1 88
2 71470 1 88
2 71471 1 88
2 71472 1 91
2 71473 1 91
2 71474 1 91
2 71475 1 91
2 71476 1 91
2 71477 1 91
2 71478 1 91
2 71479 1 91
2 71480 1 91
2 71481 1 91
2 71482 1 91
2 71483 1 91
2 71484 1 91
2 71485 1 91
2 71486 1 92
2 71487 1 92
2 71488 1 92
2 71489 1 92
2 71490 1 92
2 71491 1 92
2 71492 1 92
2 71493 1 92
2 71494 1 92
2 71495 1 92
2 71496 1 92
2 71497 1 92
2 71498 1 92
2 71499 1 93
2 71500 1 93
2 71501 1 93
2 71502 1 93
2 71503 1 93
2 71504 1 93
2 71505 1 93
2 71506 1 93
2 71507 1 93
2 71508 1 93
2 71509 1 94
2 71510 1 94
2 71511 1 94
2 71512 1 94
2 71513 1 94
2 71514 1 94
2 71515 1 94
2 71516 1 94
2 71517 1 94
2 71518 1 94
2 71519 1 94
2 71520 1 94
2 71521 1 94
2 71522 1 94
2 71523 1 94
2 71524 1 94
2 71525 1 94
2 71526 1 94
2 71527 1 94
2 71528 1 94
2 71529 1 94
2 71530 1 94
2 71531 1 94
2 71532 1 94
2 71533 1 94
2 71534 1 94
2 71535 1 94
2 71536 1 94
2 71537 1 94
2 71538 1 94
2 71539 1 94
2 71540 1 94
2 71541 1 94
2 71542 1 94
2 71543 1 94
2 71544 1 94
2 71545 1 94
2 71546 1 94
2 71547 1 94
2 71548 1 94
2 71549 1 94
2 71550 1 94
2 71551 1 95
2 71552 1 95
2 71553 1 95
2 71554 1 95
2 71555 1 95
2 71556 1 95
2 71557 1 95
2 71558 1 95
2 71559 1 95
2 71560 1 95
2 71561 1 95
2 71562 1 95
2 71563 1 95
2 71564 1 95
2 71565 1 95
2 71566 1 95
2 71567 1 95
2 71568 1 95
2 71569 1 95
2 71570 1 95
2 71571 1 95
2 71572 1 95
2 71573 1 95
2 71574 1 95
2 71575 1 95
2 71576 1 95
2 71577 1 95
2 71578 1 95
2 71579 1 95
2 71580 1 95
2 71581 1 95
2 71582 1 95
2 71583 1 95
2 71584 1 95
2 71585 1 95
2 71586 1 95
2 71587 1 95
2 71588 1 95
2 71589 1 95
2 71590 1 95
2 71591 1 95
2 71592 1 95
2 71593 1 95
2 71594 1 95
2 71595 1 95
2 71596 1 95
2 71597 1 95
2 71598 1 95
2 71599 1 95
2 71600 1 95
2 71601 1 95
2 71602 1 95
2 71603 1 95
2 71604 1 95
2 71605 1 95
2 71606 1 95
2 71607 1 95
2 71608 1 95
2 71609 1 95
2 71610 1 95
2 71611 1 96
2 71612 1 96
2 71613 1 96
2 71614 1 96
2 71615 1 97
2 71616 1 97
2 71617 1 97
2 71618 1 97
2 71619 1 97
2 71620 1 97
2 71621 1 98
2 71622 1 98
2 71623 1 98
2 71624 1 99
2 71625 1 99
2 71626 1 100
2 71627 1 100
2 71628 1 100
2 71629 1 102
2 71630 1 102
2 71631 1 102
2 71632 1 102
2 71633 1 102
2 71634 1 102
2 71635 1 102
2 71636 1 102
2 71637 1 102
2 71638 1 102
2 71639 1 109
2 71640 1 109
2 71641 1 109
2 71642 1 109
2 71643 1 109
2 71644 1 109
2 71645 1 109
2 71646 1 109
2 71647 1 109
2 71648 1 109
2 71649 1 109
2 71650 1 109
2 71651 1 109
2 71652 1 109
2 71653 1 109
2 71654 1 109
2 71655 1 109
2 71656 1 109
2 71657 1 110
2 71658 1 110
2 71659 1 110
2 71660 1 110
2 71661 1 110
2 71662 1 111
2 71663 1 111
2 71664 1 111
2 71665 1 111
2 71666 1 111
2 71667 1 111
2 71668 1 111
2 71669 1 111
2 71670 1 111
2 71671 1 111
2 71672 1 111
2 71673 1 111
2 71674 1 111
2 71675 1 111
2 71676 1 111
2 71677 1 111
2 71678 1 111
2 71679 1 111
2 71680 1 111
2 71681 1 113
2 71682 1 113
2 71683 1 114
2 71684 1 114
2 71685 1 115
2 71686 1 115
2 71687 1 115
2 71688 1 115
2 71689 1 115
2 71690 1 115
2 71691 1 115
2 71692 1 115
2 71693 1 115
2 71694 1 115
2 71695 1 115
2 71696 1 116
2 71697 1 116
2 71698 1 116
2 71699 1 116
2 71700 1 116
2 71701 1 116
2 71702 1 125
2 71703 1 125
2 71704 1 125
2 71705 1 125
2 71706 1 125
2 71707 1 126
2 71708 1 126
2 71709 1 126
2 71710 1 126
2 71711 1 126
2 71712 1 126
2 71713 1 128
2 71714 1 128
2 71715 1 128
2 71716 1 128
2 71717 1 128
2 71718 1 128
2 71719 1 128
2 71720 1 128
2 71721 1 128
2 71722 1 128
2 71723 1 128
2 71724 1 128
2 71725 1 128
2 71726 1 128
2 71727 1 128
2 71728 1 128
2 71729 1 128
2 71730 1 128
2 71731 1 128
2 71732 1 128
2 71733 1 128
2 71734 1 128
2 71735 1 128
2 71736 1 128
2 71737 1 128
2 71738 1 128
2 71739 1 128
2 71740 1 128
2 71741 1 128
2 71742 1 128
2 71743 1 128
2 71744 1 128
2 71745 1 128
2 71746 1 128
2 71747 1 128
2 71748 1 128
2 71749 1 128
2 71750 1 128
2 71751 1 128
2 71752 1 128
2 71753 1 129
2 71754 1 129
2 71755 1 129
2 71756 1 129
2 71757 1 129
2 71758 1 130
2 71759 1 130
2 71760 1 130
2 71761 1 131
2 71762 1 131
2 71763 1 131
2 71764 1 133
2 71765 1 133
2 71766 1 133
2 71767 1 134
2 71768 1 134
2 71769 1 134
2 71770 1 134
2 71771 1 134
2 71772 1 134
2 71773 1 134
2 71774 1 134
2 71775 1 134
2 71776 1 134
2 71777 1 134
2 71778 1 134
2 71779 1 134
2 71780 1 134
2 71781 1 134
2 71782 1 134
2 71783 1 134
2 71784 1 134
2 71785 1 134
2 71786 1 134
2 71787 1 135
2 71788 1 135
2 71789 1 142
2 71790 1 142
2 71791 1 142
2 71792 1 142
2 71793 1 142
2 71794 1 142
2 71795 1 142
2 71796 1 142
2 71797 1 142
2 71798 1 142
2 71799 1 142
2 71800 1 142
2 71801 1 142
2 71802 1 142
2 71803 1 142
2 71804 1 142
2 71805 1 142
2 71806 1 142
2 71807 1 142
2 71808 1 142
2 71809 1 142
2 71810 1 142
2 71811 1 142
2 71812 1 142
2 71813 1 142
2 71814 1 142
2 71815 1 142
2 71816 1 142
2 71817 1 142
2 71818 1 142
2 71819 1 142
2 71820 1 142
2 71821 1 142
2 71822 1 142
2 71823 1 142
2 71824 1 142
2 71825 1 142
2 71826 1 142
2 71827 1 142
2 71828 1 142
2 71829 1 142
2 71830 1 142
2 71831 1 142
2 71832 1 142
2 71833 1 142
2 71834 1 142
2 71835 1 142
2 71836 1 142
2 71837 1 142
2 71838 1 142
2 71839 1 142
2 71840 1 142
2 71841 1 142
2 71842 1 142
2 71843 1 142
2 71844 1 142
2 71845 1 142
2 71846 1 142
2 71847 1 142
2 71848 1 142
2 71849 1 142
2 71850 1 142
2 71851 1 142
2 71852 1 142
2 71853 1 142
2 71854 1 142
2 71855 1 142
2 71856 1 142
2 71857 1 142
2 71858 1 142
2 71859 1 142
2 71860 1 142
2 71861 1 142
2 71862 1 142
2 71863 1 142
2 71864 1 142
2 71865 1 142
2 71866 1 142
2 71867 1 142
2 71868 1 142
2 71869 1 142
2 71870 1 142
2 71871 1 142
2 71872 1 142
2 71873 1 142
2 71874 1 142
2 71875 1 142
2 71876 1 142
2 71877 1 142
2 71878 1 142
2 71879 1 142
2 71880 1 142
2 71881 1 142
2 71882 1 142
2 71883 1 142
2 71884 1 142
2 71885 1 142
2 71886 1 143
2 71887 1 143
2 71888 1 143
2 71889 1 143
2 71890 1 143
2 71891 1 143
2 71892 1 143
2 71893 1 143
2 71894 1 143
2 71895 1 143
2 71896 1 143
2 71897 1 143
2 71898 1 143
2 71899 1 143
2 71900 1 143
2 71901 1 143
2 71902 1 143
2 71903 1 143
2 71904 1 143
2 71905 1 143
2 71906 1 143
2 71907 1 143
2 71908 1 143
2 71909 1 143
2 71910 1 143
2 71911 1 143
2 71912 1 143
2 71913 1 143
2 71914 1 143
2 71915 1 143
2 71916 1 143
2 71917 1 143
2 71918 1 143
2 71919 1 143
2 71920 1 143
2 71921 1 143
2 71922 1 143
2 71923 1 143
2 71924 1 143
2 71925 1 143
2 71926 1 143
2 71927 1 143
2 71928 1 143
2 71929 1 143
2 71930 1 143
2 71931 1 143
2 71932 1 143
2 71933 1 143
2 71934 1 143
2 71935 1 143
2 71936 1 143
2 71937 1 143
2 71938 1 143
2 71939 1 143
2 71940 1 143
2 71941 1 143
2 71942 1 143
2 71943 1 143
2 71944 1 143
2 71945 1 143
2 71946 1 143
2 71947 1 143
2 71948 1 143
2 71949 1 143
2 71950 1 143
2 71951 1 143
2 71952 1 143
2 71953 1 143
2 71954 1 143
2 71955 1 143
2 71956 1 143
2 71957 1 143
2 71958 1 143
2 71959 1 143
2 71960 1 143
2 71961 1 143
2 71962 1 143
2 71963 1 143
2 71964 1 143
2 71965 1 143
2 71966 1 143
2 71967 1 143
2 71968 1 143
2 71969 1 143
2 71970 1 143
2 71971 1 143
2 71972 1 143
2 71973 1 143
2 71974 1 143
2 71975 1 143
2 71976 1 143
2 71977 1 143
2 71978 1 143
2 71979 1 143
2 71980 1 143
2 71981 1 143
2 71982 1 143
2 71983 1 143
2 71984 1 143
2 71985 1 143
2 71986 1 143
2 71987 1 143
2 71988 1 143
2 71989 1 143
2 71990 1 143
2 71991 1 143
2 71992 1 143
2 71993 1 143
2 71994 1 143
2 71995 1 143
2 71996 1 144
2 71997 1 144
2 71998 1 144
2 71999 1 144
2 72000 1 144
2 72001 1 144
2 72002 1 144
2 72003 1 144
2 72004 1 144
2 72005 1 144
2 72006 1 144
2 72007 1 144
2 72008 1 144
2 72009 1 144
2 72010 1 144
2 72011 1 144
2 72012 1 144
2 72013 1 144
2 72014 1 144
2 72015 1 144
2 72016 1 144
2 72017 1 144
2 72018 1 144
2 72019 1 144
2 72020 1 144
2 72021 1 144
2 72022 1 144
2 72023 1 144
2 72024 1 144
2 72025 1 144
2 72026 1 144
2 72027 1 144
2 72028 1 144
2 72029 1 144
2 72030 1 144
2 72031 1 144
2 72032 1 144
2 72033 1 144
2 72034 1 144
2 72035 1 144
2 72036 1 144
2 72037 1 144
2 72038 1 144
2 72039 1 144
2 72040 1 144
2 72041 1 144
2 72042 1 144
2 72043 1 144
2 72044 1 144
2 72045 1 144
2 72046 1 144
2 72047 1 144
2 72048 1 144
2 72049 1 144
2 72050 1 144
2 72051 1 144
2 72052 1 144
2 72053 1 144
2 72054 1 144
2 72055 1 144
2 72056 1 144
2 72057 1 144
2 72058 1 144
2 72059 1 144
2 72060 1 144
2 72061 1 144
2 72062 1 144
2 72063 1 144
2 72064 1 144
2 72065 1 144
2 72066 1 144
2 72067 1 144
2 72068 1 144
2 72069 1 144
2 72070 1 144
2 72071 1 144
2 72072 1 144
2 72073 1 144
2 72074 1 144
2 72075 1 144
2 72076 1 144
2 72077 1 144
2 72078 1 144
2 72079 1 144
2 72080 1 144
2 72081 1 144
2 72082 1 144
2 72083 1 144
2 72084 1 144
2 72085 1 144
2 72086 1 144
2 72087 1 144
2 72088 1 144
2 72089 1 144
2 72090 1 144
2 72091 1 144
2 72092 1 144
2 72093 1 144
2 72094 1 144
2 72095 1 145
2 72096 1 145
2 72097 1 145
2 72098 1 145
2 72099 1 145
2 72100 1 145
2 72101 1 145
2 72102 1 145
2 72103 1 145
2 72104 1 145
2 72105 1 145
2 72106 1 145
2 72107 1 145
2 72108 1 145
2 72109 1 145
2 72110 1 145
2 72111 1 145
2 72112 1 145
2 72113 1 145
2 72114 1 145
2 72115 1 145
2 72116 1 145
2 72117 1 145
2 72118 1 145
2 72119 1 145
2 72120 1 145
2 72121 1 145
2 72122 1 145
2 72123 1 145
2 72124 1 145
2 72125 1 145
2 72126 1 145
2 72127 1 145
2 72128 1 145
2 72129 1 145
2 72130 1 145
2 72131 1 145
2 72132 1 145
2 72133 1 145
2 72134 1 145
2 72135 1 145
2 72136 1 145
2 72137 1 145
2 72138 1 145
2 72139 1 145
2 72140 1 145
2 72141 1 145
2 72142 1 145
2 72143 1 145
2 72144 1 145
2 72145 1 145
2 72146 1 145
2 72147 1 145
2 72148 1 145
2 72149 1 145
2 72150 1 145
2 72151 1 145
2 72152 1 145
2 72153 1 145
2 72154 1 145
2 72155 1 145
2 72156 1 145
2 72157 1 145
2 72158 1 145
2 72159 1 145
2 72160 1 145
2 72161 1 145
2 72162 1 145
2 72163 1 145
2 72164 1 145
2 72165 1 145
2 72166 1 145
2 72167 1 145
2 72168 1 145
2 72169 1 145
2 72170 1 145
2 72171 1 145
2 72172 1 145
2 72173 1 145
2 72174 1 145
2 72175 1 145
2 72176 1 145
2 72177 1 145
2 72178 1 145
2 72179 1 145
2 72180 1 145
2 72181 1 145
2 72182 1 145
2 72183 1 145
2 72184 1 145
2 72185 1 145
2 72186 1 145
2 72187 1 145
2 72188 1 145
2 72189 1 145
2 72190 1 145
2 72191 1 145
2 72192 1 145
2 72193 1 145
2 72194 1 145
2 72195 1 145
2 72196 1 145
2 72197 1 145
2 72198 1 145
2 72199 1 145
2 72200 1 145
2 72201 1 145
2 72202 1 145
2 72203 1 145
2 72204 1 145
2 72205 1 145
2 72206 1 145
2 72207 1 145
2 72208 1 145
2 72209 1 145
2 72210 1 145
2 72211 1 145
2 72212 1 145
2 72213 1 145
2 72214 1 145
2 72215 1 145
2 72216 1 145
2 72217 1 145
2 72218 1 146
2 72219 1 146
2 72220 1 146
2 72221 1 146
2 72222 1 146
2 72223 1 146
2 72224 1 146
2 72225 1 146
2 72226 1 146
2 72227 1 146
2 72228 1 146
2 72229 1 146
2 72230 1 146
2 72231 1 146
2 72232 1 147
2 72233 1 147
2 72234 1 148
2 72235 1 148
2 72236 1 149
2 72237 1 149
2 72238 1 149
2 72239 1 150
2 72240 1 150
2 72241 1 150
2 72242 1 150
2 72243 1 150
2 72244 1 150
2 72245 1 150
2 72246 1 150
2 72247 1 150
2 72248 1 150
2 72249 1 150
2 72250 1 150
2 72251 1 150
2 72252 1 150
2 72253 1 152
2 72254 1 152
2 72255 1 152
2 72256 1 152
2 72257 1 152
2 72258 1 152
2 72259 1 152
2 72260 1 152
2 72261 1 152
2 72262 1 152
2 72263 1 152
2 72264 1 152
2 72265 1 152
2 72266 1 152
2 72267 1 152
2 72268 1 152
2 72269 1 152
2 72270 1 152
2 72271 1 152
2 72272 1 152
2 72273 1 152
2 72274 1 152
2 72275 1 152
2 72276 1 152
2 72277 1 152
2 72278 1 152
2 72279 1 152
2 72280 1 152
2 72281 1 152
2 72282 1 153
2 72283 1 153
2 72284 1 154
2 72285 1 154
2 72286 1 154
2 72287 1 154
2 72288 1 154
2 72289 1 154
2 72290 1 154
2 72291 1 154
2 72292 1 154
2 72293 1 154
2 72294 1 154
2 72295 1 154
2 72296 1 155
2 72297 1 155
2 72298 1 155
2 72299 1 155
2 72300 1 155
2 72301 1 155
2 72302 1 155
2 72303 1 155
2 72304 1 155
2 72305 1 155
2 72306 1 156
2 72307 1 156
2 72308 1 156
2 72309 1 156
2 72310 1 158
2 72311 1 158
2 72312 1 158
2 72313 1 158
2 72314 1 158
2 72315 1 158
2 72316 1 158
2 72317 1 158
2 72318 1 158
2 72319 1 158
2 72320 1 158
2 72321 1 158
2 72322 1 158
2 72323 1 158
2 72324 1 158
2 72325 1 158
2 72326 1 158
2 72327 1 158
2 72328 1 158
2 72329 1 158
2 72330 1 158
2 72331 1 160
2 72332 1 160
2 72333 1 160
2 72334 1 160
2 72335 1 160
2 72336 1 160
2 72337 1 160
2 72338 1 160
2 72339 1 160
2 72340 1 161
2 72341 1 161
2 72342 1 161
2 72343 1 161
2 72344 1 161
2 72345 1 161
2 72346 1 161
2 72347 1 161
2 72348 1 161
2 72349 1 161
2 72350 1 161
2 72351 1 161
2 72352 1 161
2 72353 1 162
2 72354 1 162
2 72355 1 163
2 72356 1 163
2 72357 1 173
2 72358 1 173
2 72359 1 173
2 72360 1 173
2 72361 1 173
2 72362 1 173
2 72363 1 173
2 72364 1 173
2 72365 1 173
2 72366 1 173
2 72367 1 173
2 72368 1 173
2 72369 1 173
2 72370 1 173
2 72371 1 173
2 72372 1 173
2 72373 1 173
2 72374 1 173
2 72375 1 173
2 72376 1 173
2 72377 1 173
2 72378 1 173
2 72379 1 175
2 72380 1 175
2 72381 1 175
2 72382 1 175
2 72383 1 175
2 72384 1 175
2 72385 1 175
2 72386 1 175
2 72387 1 175
2 72388 1 175
2 72389 1 175
2 72390 1 175
2 72391 1 175
2 72392 1 177
2 72393 1 177
2 72394 1 177
2 72395 1 178
2 72396 1 178
2 72397 1 178
2 72398 1 178
2 72399 1 178
2 72400 1 179
2 72401 1 179
2 72402 1 179
2 72403 1 182
2 72404 1 182
2 72405 1 185
2 72406 1 185
2 72407 1 185
2 72408 1 185
2 72409 1 185
2 72410 1 185
2 72411 1 185
2 72412 1 185
2 72413 1 185
2 72414 1 185
2 72415 1 185
2 72416 1 187
2 72417 1 187
2 72418 1 187
2 72419 1 187
2 72420 1 187
2 72421 1 187
2 72422 1 187
2 72423 1 187
2 72424 1 187
2 72425 1 187
2 72426 1 187
2 72427 1 187
2 72428 1 189
2 72429 1 189
2 72430 1 189
2 72431 1 189
2 72432 1 190
2 72433 1 190
2 72434 1 190
2 72435 1 195
2 72436 1 195
2 72437 1 195
2 72438 1 195
2 72439 1 195
2 72440 1 195
2 72441 1 195
2 72442 1 195
2 72443 1 195
2 72444 1 195
2 72445 1 195
2 72446 1 195
2 72447 1 195
2 72448 1 195
2 72449 1 195
2 72450 1 195
2 72451 1 195
2 72452 1 195
2 72453 1 195
2 72454 1 195
2 72455 1 195
2 72456 1 195
2 72457 1 195
2 72458 1 195
2 72459 1 195
2 72460 1 195
2 72461 1 195
2 72462 1 195
2 72463 1 195
2 72464 1 195
2 72465 1 195
2 72466 1 195
2 72467 1 195
2 72468 1 195
2 72469 1 195
2 72470 1 195
2 72471 1 195
2 72472 1 195
2 72473 1 195
2 72474 1 195
2 72475 1 195
2 72476 1 195
2 72477 1 195
2 72478 1 196
2 72479 1 196
2 72480 1 196
2 72481 1 196
2 72482 1 197
2 72483 1 197
2 72484 1 197
2 72485 1 197
2 72486 1 198
2 72487 1 198
2 72488 1 198
2 72489 1 198
2 72490 1 198
2 72491 1 198
2 72492 1 198
2 72493 1 198
2 72494 1 199
2 72495 1 199
2 72496 1 199
2 72497 1 199
2 72498 1 199
2 72499 1 199
2 72500 1 199
2 72501 1 199
2 72502 1 199
2 72503 1 199
2 72504 1 199
2 72505 1 199
2 72506 1 199
2 72507 1 199
2 72508 1 199
2 72509 1 199
2 72510 1 199
2 72511 1 199
2 72512 1 199
2 72513 1 199
2 72514 1 199
2 72515 1 199
2 72516 1 199
2 72517 1 199
2 72518 1 199
2 72519 1 199
2 72520 1 199
2 72521 1 199
2 72522 1 199
2 72523 1 199
2 72524 1 199
2 72525 1 199
2 72526 1 199
2 72527 1 199
2 72528 1 199
2 72529 1 199
2 72530 1 199
2 72531 1 199
2 72532 1 199
2 72533 1 199
2 72534 1 199
2 72535 1 199
2 72536 1 199
2 72537 1 199
2 72538 1 199
2 72539 1 199
2 72540 1 199
2 72541 1 199
2 72542 1 199
2 72543 1 199
2 72544 1 199
2 72545 1 199
2 72546 1 199
2 72547 1 199
2 72548 1 199
2 72549 1 199
2 72550 1 199
2 72551 1 199
2 72552 1 199
2 72553 1 199
2 72554 1 199
2 72555 1 199
2 72556 1 199
2 72557 1 199
2 72558 1 199
2 72559 1 199
2 72560 1 199
2 72561 1 199
2 72562 1 199
2 72563 1 199
2 72564 1 199
2 72565 1 199
2 72566 1 199
2 72567 1 199
2 72568 1 199
2 72569 1 199
2 72570 1 199
2 72571 1 199
2 72572 1 199
2 72573 1 199
2 72574 1 199
2 72575 1 199
2 72576 1 199
2 72577 1 199
2 72578 1 199
2 72579 1 199
2 72580 1 199
2 72581 1 199
2 72582 1 199
2 72583 1 199
2 72584 1 199
2 72585 1 199
2 72586 1 199
2 72587 1 199
2 72588 1 199
2 72589 1 199
2 72590 1 199
2 72591 1 199
2 72592 1 199
2 72593 1 199
2 72594 1 199
2 72595 1 199
2 72596 1 199
2 72597 1 199
2 72598 1 199
2 72599 1 200
2 72600 1 200
2 72601 1 200
2 72602 1 200
2 72603 1 200
2 72604 1 200
2 72605 1 200
2 72606 1 200
2 72607 1 200
2 72608 1 200
2 72609 1 200
2 72610 1 200
2 72611 1 200
2 72612 1 200
2 72613 1 200
2 72614 1 200
2 72615 1 200
2 72616 1 200
2 72617 1 200
2 72618 1 200
2 72619 1 200
2 72620 1 200
2 72621 1 200
2 72622 1 200
2 72623 1 200
2 72624 1 200
2 72625 1 200
2 72626 1 200
2 72627 1 200
2 72628 1 200
2 72629 1 200
2 72630 1 200
2 72631 1 200
2 72632 1 200
2 72633 1 200
2 72634 1 200
2 72635 1 200
2 72636 1 200
2 72637 1 200
2 72638 1 200
2 72639 1 200
2 72640 1 200
2 72641 1 200
2 72642 1 200
2 72643 1 200
2 72644 1 200
2 72645 1 200
2 72646 1 200
2 72647 1 200
2 72648 1 200
2 72649 1 200
2 72650 1 200
2 72651 1 200
2 72652 1 200
2 72653 1 200
2 72654 1 200
2 72655 1 200
2 72656 1 200
2 72657 1 200
2 72658 1 200
2 72659 1 200
2 72660 1 200
2 72661 1 200
2 72662 1 200
2 72663 1 200
2 72664 1 200
2 72665 1 200
2 72666 1 200
2 72667 1 200
2 72668 1 200
2 72669 1 200
2 72670 1 200
2 72671 1 200
2 72672 1 200
2 72673 1 200
2 72674 1 200
2 72675 1 200
2 72676 1 200
2 72677 1 200
2 72678 1 200
2 72679 1 200
2 72680 1 200
2 72681 1 200
2 72682 1 200
2 72683 1 200
2 72684 1 200
2 72685 1 200
2 72686 1 201
2 72687 1 201
2 72688 1 201
2 72689 1 201
2 72690 1 201
2 72691 1 201
2 72692 1 201
2 72693 1 201
2 72694 1 201
2 72695 1 201
2 72696 1 201
2 72697 1 201
2 72698 1 201
2 72699 1 201
2 72700 1 201
2 72701 1 201
2 72702 1 201
2 72703 1 201
2 72704 1 201
2 72705 1 201
2 72706 1 201
2 72707 1 201
2 72708 1 201
2 72709 1 201
2 72710 1 201
2 72711 1 201
2 72712 1 201
2 72713 1 201
2 72714 1 202
2 72715 1 202
2 72716 1 202
2 72717 1 202
2 72718 1 202
2 72719 1 202
2 72720 1 202
2 72721 1 202
2 72722 1 202
2 72723 1 202
2 72724 1 202
2 72725 1 202
2 72726 1 202
2 72727 1 202
2 72728 1 202
2 72729 1 202
2 72730 1 203
2 72731 1 203
2 72732 1 203
2 72733 1 203
2 72734 1 204
2 72735 1 204
2 72736 1 205
2 72737 1 205
2 72738 1 206
2 72739 1 206
2 72740 1 206
2 72741 1 206
2 72742 1 213
2 72743 1 213
2 72744 1 213
2 72745 1 213
2 72746 1 213
2 72747 1 213
2 72748 1 213
2 72749 1 213
2 72750 1 213
2 72751 1 213
2 72752 1 213
2 72753 1 214
2 72754 1 214
2 72755 1 214
2 72756 1 215
2 72757 1 215
2 72758 1 215
2 72759 1 215
2 72760 1 215
2 72761 1 216
2 72762 1 216
2 72763 1 216
2 72764 1 216
2 72765 1 216
2 72766 1 216
2 72767 1 216
2 72768 1 217
2 72769 1 217
2 72770 1 218
2 72771 1 218
2 72772 1 218
2 72773 1 218
2 72774 1 218
2 72775 1 218
2 72776 1 218
2 72777 1 218
2 72778 1 218
2 72779 1 218
2 72780 1 218
2 72781 1 218
2 72782 1 218
2 72783 1 218
2 72784 1 218
2 72785 1 218
2 72786 1 218
2 72787 1 218
2 72788 1 218
2 72789 1 218
2 72790 1 218
2 72791 1 218
2 72792 1 218
2 72793 1 218
2 72794 1 218
2 72795 1 218
2 72796 1 218
2 72797 1 218
2 72798 1 218
2 72799 1 218
2 72800 1 218
2 72801 1 218
2 72802 1 218
2 72803 1 218
2 72804 1 218
2 72805 1 218
2 72806 1 218
2 72807 1 218
2 72808 1 218
2 72809 1 218
2 72810 1 218
2 72811 1 218
2 72812 1 219
2 72813 1 219
2 72814 1 219
2 72815 1 219
2 72816 1 219
2 72817 1 219
2 72818 1 219
2 72819 1 219
2 72820 1 219
2 72821 1 219
2 72822 1 219
2 72823 1 219
2 72824 1 219
2 72825 1 219
2 72826 1 219
2 72827 1 219
2 72828 1 219
2 72829 1 219
2 72830 1 219
2 72831 1 219
2 72832 1 219
2 72833 1 219
2 72834 1 219
2 72835 1 219
2 72836 1 219
2 72837 1 219
2 72838 1 219
2 72839 1 219
2 72840 1 219
2 72841 1 220
2 72842 1 220
2 72843 1 221
2 72844 1 221
2 72845 1 227
2 72846 1 227
2 72847 1 227
2 72848 1 227
2 72849 1 227
2 72850 1 227
2 72851 1 227
2 72852 1 227
2 72853 1 227
2 72854 1 227
2 72855 1 227
2 72856 1 227
2 72857 1 227
2 72858 1 227
2 72859 1 227
2 72860 1 227
2 72861 1 227
2 72862 1 227
2 72863 1 227
2 72864 1 227
2 72865 1 227
2 72866 1 227
2 72867 1 228
2 72868 1 228
2 72869 1 228
2 72870 1 228
2 72871 1 228
2 72872 1 228
2 72873 1 228
2 72874 1 228
2 72875 1 229
2 72876 1 229
2 72877 1 229
2 72878 1 229
2 72879 1 229
2 72880 1 229
2 72881 1 229
2 72882 1 229
2 72883 1 229
2 72884 1 229
2 72885 1 231
2 72886 1 231
2 72887 1 231
2 72888 1 231
2 72889 1 231
2 72890 1 231
2 72891 1 232
2 72892 1 232
2 72893 1 232
2 72894 1 232
2 72895 1 233
2 72896 1 233
2 72897 1 233
2 72898 1 233
2 72899 1 233
2 72900 1 233
2 72901 1 233
2 72902 1 233
2 72903 1 233
2 72904 1 234
2 72905 1 234
2 72906 1 234
2 72907 1 234
2 72908 1 234
2 72909 1 234
2 72910 1 234
2 72911 1 234
2 72912 1 234
2 72913 1 234
2 72914 1 234
2 72915 1 234
2 72916 1 234
2 72917 1 234
2 72918 1 234
2 72919 1 234
2 72920 1 234
2 72921 1 234
2 72922 1 234
2 72923 1 234
2 72924 1 234
2 72925 1 234
2 72926 1 234
2 72927 1 235
2 72928 1 235
2 72929 1 235
2 72930 1 235
2 72931 1 235
2 72932 1 235
2 72933 1 235
2 72934 1 235
2 72935 1 236
2 72936 1 236
2 72937 1 251
2 72938 1 251
2 72939 1 251
2 72940 1 251
2 72941 1 251
2 72942 1 251
2 72943 1 251
2 72944 1 251
2 72945 1 251
2 72946 1 251
2 72947 1 252
2 72948 1 252
2 72949 1 252
2 72950 1 252
2 72951 1 252
2 72952 1 253
2 72953 1 253
2 72954 1 253
2 72955 1 253
2 72956 1 254
2 72957 1 254
2 72958 1 254
2 72959 1 254
2 72960 1 254
2 72961 1 254
2 72962 1 254
2 72963 1 254
2 72964 1 254
2 72965 1 254
2 72966 1 254
2 72967 1 254
2 72968 1 254
2 72969 1 254
2 72970 1 254
2 72971 1 254
2 72972 1 254
2 72973 1 254
2 72974 1 254
2 72975 1 254
2 72976 1 254
2 72977 1 254
2 72978 1 254
2 72979 1 254
2 72980 1 254
2 72981 1 254
2 72982 1 254
2 72983 1 254
2 72984 1 254
2 72985 1 254
2 72986 1 254
2 72987 1 254
2 72988 1 254
2 72989 1 254
2 72990 1 254
2 72991 1 254
2 72992 1 254
2 72993 1 254
2 72994 1 254
2 72995 1 254
2 72996 1 254
2 72997 1 254
2 72998 1 254
2 72999 1 254
2 73000 1 254
2 73001 1 254
2 73002 1 254
2 73003 1 254
2 73004 1 254
2 73005 1 254
2 73006 1 254
2 73007 1 254
2 73008 1 254
2 73009 1 254
2 73010 1 254
2 73011 1 254
2 73012 1 254
2 73013 1 254
2 73014 1 254
2 73015 1 254
2 73016 1 254
2 73017 1 254
2 73018 1 254
2 73019 1 254
2 73020 1 254
2 73021 1 254
2 73022 1 254
2 73023 1 254
2 73024 1 254
2 73025 1 254
2 73026 1 254
2 73027 1 254
2 73028 1 254
2 73029 1 254
2 73030 1 254
2 73031 1 254
2 73032 1 254
2 73033 1 254
2 73034 1 254
2 73035 1 254
2 73036 1 254
2 73037 1 254
2 73038 1 254
2 73039 1 254
2 73040 1 254
2 73041 1 254
2 73042 1 254
2 73043 1 254
2 73044 1 254
2 73045 1 254
2 73046 1 254
2 73047 1 254
2 73048 1 254
2 73049 1 254
2 73050 1 254
2 73051 1 255
2 73052 1 255
2 73053 1 255
2 73054 1 255
2 73055 1 255
2 73056 1 255
2 73057 1 255
2 73058 1 255
2 73059 1 255
2 73060 1 255
2 73061 1 255
2 73062 1 255
2 73063 1 255
2 73064 1 255
2 73065 1 255
2 73066 1 255
2 73067 1 255
2 73068 1 255
2 73069 1 255
2 73070 1 255
2 73071 1 255
2 73072 1 255
2 73073 1 255
2 73074 1 255
2 73075 1 255
2 73076 1 255
2 73077 1 255
2 73078 1 255
2 73079 1 255
2 73080 1 255
2 73081 1 255
2 73082 1 255
2 73083 1 255
2 73084 1 255
2 73085 1 255
2 73086 1 255
2 73087 1 255
2 73088 1 255
2 73089 1 255
2 73090 1 255
2 73091 1 255
2 73092 1 255
2 73093 1 255
2 73094 1 255
2 73095 1 255
2 73096 1 256
2 73097 1 256
2 73098 1 257
2 73099 1 257
2 73100 1 257
2 73101 1 257
2 73102 1 257
2 73103 1 258
2 73104 1 258
2 73105 1 258
2 73106 1 258
2 73107 1 260
2 73108 1 260
2 73109 1 260
2 73110 1 260
2 73111 1 260
2 73112 1 260
2 73113 1 260
2 73114 1 260
2 73115 1 260
2 73116 1 260
2 73117 1 260
2 73118 1 260
2 73119 1 260
2 73120 1 260
2 73121 1 260
2 73122 1 260
2 73123 1 260
2 73124 1 260
2 73125 1 260
2 73126 1 260
2 73127 1 260
2 73128 1 260
2 73129 1 260
2 73130 1 260
2 73131 1 260
2 73132 1 260
2 73133 1 260
2 73134 1 260
2 73135 1 260
2 73136 1 260
2 73137 1 260
2 73138 1 260
2 73139 1 260
2 73140 1 260
2 73141 1 260
2 73142 1 261
2 73143 1 261
2 73144 1 261
2 73145 1 261
2 73146 1 261
2 73147 1 261
2 73148 1 263
2 73149 1 263
2 73150 1 263
2 73151 1 263
2 73152 1 263
2 73153 1 263
2 73154 1 263
2 73155 1 263
2 73156 1 263
2 73157 1 263
2 73158 1 263
2 73159 1 263
2 73160 1 263
2 73161 1 263
2 73162 1 263
2 73163 1 263
2 73164 1 263
2 73165 1 263
2 73166 1 263
2 73167 1 263
2 73168 1 263
2 73169 1 263
2 73170 1 263
2 73171 1 265
2 73172 1 265
2 73173 1 265
2 73174 1 265
2 73175 1 268
2 73176 1 268
2 73177 1 268
2 73178 1 268
2 73179 1 268
2 73180 1 271
2 73181 1 271
2 73182 1 271
2 73183 1 271
2 73184 1 271
2 73185 1 271
2 73186 1 271
2 73187 1 271
2 73188 1 271
2 73189 1 271
2 73190 1 271
2 73191 1 271
2 73192 1 271
2 73193 1 271
2 73194 1 271
2 73195 1 271
2 73196 1 271
2 73197 1 271
2 73198 1 271
2 73199 1 271
2 73200 1 271
2 73201 1 271
2 73202 1 271
2 73203 1 271
2 73204 1 271
2 73205 1 271
2 73206 1 271
2 73207 1 271
2 73208 1 271
2 73209 1 271
2 73210 1 271
2 73211 1 271
2 73212 1 271
2 73213 1 271
2 73214 1 271
2 73215 1 271
2 73216 1 271
2 73217 1 271
2 73218 1 271
2 73219 1 271
2 73220 1 271
2 73221 1 271
2 73222 1 271
2 73223 1 271
2 73224 1 271
2 73225 1 271
2 73226 1 271
2 73227 1 271
2 73228 1 271
2 73229 1 271
2 73230 1 271
2 73231 1 271
2 73232 1 271
2 73233 1 272
2 73234 1 272
2 73235 1 272
2 73236 1 272
2 73237 1 272
2 73238 1 272
2 73239 1 272
2 73240 1 272
2 73241 1 272
2 73242 1 272
2 73243 1 272
2 73244 1 272
2 73245 1 272
2 73246 1 272
2 73247 1 272
2 73248 1 272
2 73249 1 272
2 73250 1 272
2 73251 1 272
2 73252 1 272
2 73253 1 272
2 73254 1 272
2 73255 1 272
2 73256 1 272
2 73257 1 272
2 73258 1 272
2 73259 1 272
2 73260 1 272
2 73261 1 272
2 73262 1 272
2 73263 1 272
2 73264 1 272
2 73265 1 272
2 73266 1 272
2 73267 1 272
2 73268 1 272
2 73269 1 272
2 73270 1 273
2 73271 1 273
2 73272 1 274
2 73273 1 274
2 73274 1 276
2 73275 1 276
2 73276 1 283
2 73277 1 283
2 73278 1 283
2 73279 1 283
2 73280 1 283
2 73281 1 283
2 73282 1 283
2 73283 1 283
2 73284 1 283
2 73285 1 283
2 73286 1 283
2 73287 1 283
2 73288 1 283
2 73289 1 283
2 73290 1 283
2 73291 1 283
2 73292 1 283
2 73293 1 283
2 73294 1 283
2 73295 1 283
2 73296 1 283
2 73297 1 283
2 73298 1 283
2 73299 1 283
2 73300 1 283
2 73301 1 283
2 73302 1 283
2 73303 1 283
2 73304 1 283
2 73305 1 283
2 73306 1 283
2 73307 1 283
2 73308 1 283
2 73309 1 283
2 73310 1 283
2 73311 1 283
2 73312 1 283
2 73313 1 283
2 73314 1 283
2 73315 1 283
2 73316 1 283
2 73317 1 283
2 73318 1 283
2 73319 1 283
2 73320 1 283
2 73321 1 283
2 73322 1 283
2 73323 1 283
2 73324 1 283
2 73325 1 283
2 73326 1 283
2 73327 1 283
2 73328 1 283
2 73329 1 283
2 73330 1 283
2 73331 1 283
2 73332 1 283
2 73333 1 283
2 73334 1 283
2 73335 1 283
2 73336 1 283
2 73337 1 283
2 73338 1 283
2 73339 1 283
2 73340 1 283
2 73341 1 283
2 73342 1 283
2 73343 1 283
2 73344 1 283
2 73345 1 283
2 73346 1 283
2 73347 1 283
2 73348 1 283
2 73349 1 283
2 73350 1 283
2 73351 1 283
2 73352 1 283
2 73353 1 283
2 73354 1 283
2 73355 1 283
2 73356 1 283
2 73357 1 283
2 73358 1 283
2 73359 1 283
2 73360 1 283
2 73361 1 283
2 73362 1 283
2 73363 1 283
2 73364 1 283
2 73365 1 283
2 73366 1 283
2 73367 1 284
2 73368 1 284
2 73369 1 284
2 73370 1 284
2 73371 1 284
2 73372 1 284
2 73373 1 284
2 73374 1 284
2 73375 1 284
2 73376 1 284
2 73377 1 284
2 73378 1 284
2 73379 1 284
2 73380 1 284
2 73381 1 284
2 73382 1 284
2 73383 1 284
2 73384 1 284
2 73385 1 284
2 73386 1 284
2 73387 1 284
2 73388 1 284
2 73389 1 284
2 73390 1 284
2 73391 1 284
2 73392 1 284
2 73393 1 284
2 73394 1 284
2 73395 1 284
2 73396 1 284
2 73397 1 284
2 73398 1 284
2 73399 1 284
2 73400 1 284
2 73401 1 284
2 73402 1 284
2 73403 1 284
2 73404 1 284
2 73405 1 284
2 73406 1 284
2 73407 1 284
2 73408 1 284
2 73409 1 284
2 73410 1 284
2 73411 1 284
2 73412 1 284
2 73413 1 284
2 73414 1 284
2 73415 1 284
2 73416 1 284
2 73417 1 284
2 73418 1 284
2 73419 1 284
2 73420 1 284
2 73421 1 284
2 73422 1 284
2 73423 1 284
2 73424 1 284
2 73425 1 284
2 73426 1 284
2 73427 1 284
2 73428 1 284
2 73429 1 284
2 73430 1 284
2 73431 1 284
2 73432 1 284
2 73433 1 284
2 73434 1 284
2 73435 1 284
2 73436 1 284
2 73437 1 284
2 73438 1 284
2 73439 1 284
2 73440 1 284
2 73441 1 284
2 73442 1 284
2 73443 1 284
2 73444 1 284
2 73445 1 284
2 73446 1 284
2 73447 1 284
2 73448 1 284
2 73449 1 284
2 73450 1 284
2 73451 1 284
2 73452 1 284
2 73453 1 284
2 73454 1 284
2 73455 1 284
2 73456 1 284
2 73457 1 284
2 73458 1 284
2 73459 1 284
2 73460 1 284
2 73461 1 284
2 73462 1 284
2 73463 1 284
2 73464 1 284
2 73465 1 284
2 73466 1 284
2 73467 1 284
2 73468 1 284
2 73469 1 284
2 73470 1 284
2 73471 1 284
2 73472 1 284
2 73473 1 284
2 73474 1 284
2 73475 1 284
2 73476 1 284
2 73477 1 284
2 73478 1 284
2 73479 1 284
2 73480 1 284
2 73481 1 284
2 73482 1 284
2 73483 1 284
2 73484 1 284
2 73485 1 284
2 73486 1 284
2 73487 1 284
2 73488 1 284
2 73489 1 284
2 73490 1 284
2 73491 1 284
2 73492 1 284
2 73493 1 284
2 73494 1 284
2 73495 1 284
2 73496 1 284
2 73497 1 284
2 73498 1 284
2 73499 1 284
2 73500 1 284
2 73501 1 284
2 73502 1 284
2 73503 1 284
2 73504 1 284
2 73505 1 284
2 73506 1 284
2 73507 1 284
2 73508 1 284
2 73509 1 284
2 73510 1 284
2 73511 1 284
2 73512 1 284
2 73513 1 284
2 73514 1 284
2 73515 1 284
2 73516 1 284
2 73517 1 284
2 73518 1 284
2 73519 1 284
2 73520 1 284
2 73521 1 284
2 73522 1 284
2 73523 1 285
2 73524 1 285
2 73525 1 285
2 73526 1 286
2 73527 1 286
2 73528 1 286
2 73529 1 286
2 73530 1 287
2 73531 1 287
2 73532 1 287
2 73533 1 287
2 73534 1 287
2 73535 1 287
2 73536 1 287
2 73537 1 287
2 73538 1 287
2 73539 1 287
2 73540 1 287
2 73541 1 287
2 73542 1 287
2 73543 1 287
2 73544 1 287
2 73545 1 287
2 73546 1 287
2 73547 1 287
2 73548 1 287
2 73549 1 287
2 73550 1 287
2 73551 1 287
2 73552 1 287
2 73553 1 287
2 73554 1 287
2 73555 1 287
2 73556 1 287
2 73557 1 287
2 73558 1 287
2 73559 1 287
2 73560 1 288
2 73561 1 288
2 73562 1 288
2 73563 1 288
2 73564 1 288
2 73565 1 288
2 73566 1 288
2 73567 1 288
2 73568 1 288
2 73569 1 288
2 73570 1 288
2 73571 1 288
2 73572 1 288
2 73573 1 288
2 73574 1 288
2 73575 1 288
2 73576 1 288
2 73577 1 288
2 73578 1 288
2 73579 1 288
2 73580 1 288
2 73581 1 288
2 73582 1 288
2 73583 1 288
2 73584 1 288
2 73585 1 288
2 73586 1 288
2 73587 1 288
2 73588 1 288
2 73589 1 288
2 73590 1 288
2 73591 1 288
2 73592 1 288
2 73593 1 295
2 73594 1 295
2 73595 1 295
2 73596 1 295
2 73597 1 295
2 73598 1 295
2 73599 1 295
2 73600 1 295
2 73601 1 295
2 73602 1 295
2 73603 1 295
2 73604 1 295
2 73605 1 295
2 73606 1 295
2 73607 1 295
2 73608 1 295
2 73609 1 295
2 73610 1 295
2 73611 1 295
2 73612 1 295
2 73613 1 295
2 73614 1 295
2 73615 1 295
2 73616 1 295
2 73617 1 295
2 73618 1 297
2 73619 1 297
2 73620 1 297
2 73621 1 297
2 73622 1 297
2 73623 1 297
2 73624 1 297
2 73625 1 297
2 73626 1 297
2 73627 1 297
2 73628 1 298
2 73629 1 298
2 73630 1 299
2 73631 1 299
2 73632 1 299
2 73633 1 300
2 73634 1 300
2 73635 1 300
2 73636 1 302
2 73637 1 302
2 73638 1 302
2 73639 1 302
2 73640 1 302
2 73641 1 302
2 73642 1 302
2 73643 1 302
2 73644 1 302
2 73645 1 302
2 73646 1 302
2 73647 1 302
2 73648 1 302
2 73649 1 302
2 73650 1 302
2 73651 1 302
2 73652 1 302
2 73653 1 302
2 73654 1 302
2 73655 1 302
2 73656 1 302
2 73657 1 302
2 73658 1 304
2 73659 1 304
2 73660 1 305
2 73661 1 305
2 73662 1 305
2 73663 1 305
2 73664 1 305
2 73665 1 305
2 73666 1 305
2 73667 1 319
2 73668 1 319
2 73669 1 319
2 73670 1 319
2 73671 1 319
2 73672 1 319
2 73673 1 321
2 73674 1 321
2 73675 1 322
2 73676 1 322
2 73677 1 322
2 73678 1 322
2 73679 1 322
2 73680 1 322
2 73681 1 322
2 73682 1 322
2 73683 1 322
2 73684 1 322
2 73685 1 322
2 73686 1 322
2 73687 1 322
2 73688 1 322
2 73689 1 322
2 73690 1 322
2 73691 1 322
2 73692 1 322
2 73693 1 323
2 73694 1 323
2 73695 1 323
2 73696 1 323
2 73697 1 323
2 73698 1 323
2 73699 1 323
2 73700 1 323
2 73701 1 323
2 73702 1 323
2 73703 1 324
2 73704 1 324
2 73705 1 324
2 73706 1 324
2 73707 1 335
2 73708 1 335
2 73709 1 335
2 73710 1 335
2 73711 1 335
2 73712 1 335
2 73713 1 335
2 73714 1 335
2 73715 1 335
2 73716 1 335
2 73717 1 335
2 73718 1 335
2 73719 1 336
2 73720 1 336
2 73721 1 336
2 73722 1 337
2 73723 1 337
2 73724 1 339
2 73725 1 339
2 73726 1 339
2 73727 1 339
2 73728 1 339
2 73729 1 339
2 73730 1 339
2 73731 1 339
2 73732 1 341
2 73733 1 341
2 73734 1 346
2 73735 1 346
2 73736 1 346
2 73737 1 346
2 73738 1 346
2 73739 1 346
2 73740 1 346
2 73741 1 346
2 73742 1 346
2 73743 1 346
2 73744 1 346
2 73745 1 346
2 73746 1 346
2 73747 1 346
2 73748 1 346
2 73749 1 348
2 73750 1 348
2 73751 1 348
2 73752 1 348
2 73753 1 348
2 73754 1 348
2 73755 1 348
2 73756 1 348
2 73757 1 349
2 73758 1 349
2 73759 1 349
2 73760 1 360
2 73761 1 360
2 73762 1 360
2 73763 1 360
2 73764 1 360
2 73765 1 360
2 73766 1 360
2 73767 1 360
2 73768 1 360
2 73769 1 360
2 73770 1 360
2 73771 1 360
2 73772 1 360
2 73773 1 360
2 73774 1 360
2 73775 1 360
2 73776 1 360
2 73777 1 360
2 73778 1 360
2 73779 1 360
2 73780 1 360
2 73781 1 360
2 73782 1 360
2 73783 1 360
2 73784 1 360
2 73785 1 361
2 73786 1 361
2 73787 1 361
2 73788 1 361
2 73789 1 362
2 73790 1 362
2 73791 1 365
2 73792 1 365
2 73793 1 365
2 73794 1 374
2 73795 1 374
2 73796 1 377
2 73797 1 377
2 73798 1 377
2 73799 1 377
2 73800 1 377
2 73801 1 377
2 73802 1 377
2 73803 1 377
2 73804 1 377
2 73805 1 377
2 73806 1 377
2 73807 1 377
2 73808 1 377
2 73809 1 377
2 73810 1 377
2 73811 1 377
2 73812 1 377
2 73813 1 377
2 73814 1 377
2 73815 1 377
2 73816 1 377
2 73817 1 379
2 73818 1 379
2 73819 1 379
2 73820 1 379
2 73821 1 379
2 73822 1 379
2 73823 1 379
2 73824 1 379
2 73825 1 379
2 73826 1 379
2 73827 1 379
2 73828 1 379
2 73829 1 379
2 73830 1 379
2 73831 1 379
2 73832 1 379
2 73833 1 379
2 73834 1 379
2 73835 1 379
2 73836 1 379
2 73837 1 379
2 73838 1 379
2 73839 1 379
2 73840 1 380
2 73841 1 380
2 73842 1 380
2 73843 1 380
2 73844 1 380
2 73845 1 380
2 73846 1 380
2 73847 1 380
2 73848 1 380
2 73849 1 380
2 73850 1 380
2 73851 1 380
2 73852 1 380
2 73853 1 380
2 73854 1 380
2 73855 1 380
2 73856 1 380
2 73857 1 380
2 73858 1 380
2 73859 1 382
2 73860 1 382
2 73861 1 382
2 73862 1 382
2 73863 1 382
2 73864 1 382
2 73865 1 382
2 73866 1 382
2 73867 1 384
2 73868 1 384
2 73869 1 384
2 73870 1 388
2 73871 1 388
2 73872 1 395
2 73873 1 395
2 73874 1 395
2 73875 1 396
2 73876 1 396
2 73877 1 396
2 73878 1 396
2 73879 1 396
2 73880 1 396
2 73881 1 396
2 73882 1 396
2 73883 1 397
2 73884 1 397
2 73885 1 397
2 73886 1 397
2 73887 1 397
2 73888 1 397
2 73889 1 398
2 73890 1 398
2 73891 1 400
2 73892 1 400
2 73893 1 403
2 73894 1 403
2 73895 1 403
2 73896 1 403
2 73897 1 403
2 73898 1 403
2 73899 1 403
2 73900 1 410
2 73901 1 410
2 73902 1 410
2 73903 1 410
2 73904 1 410
2 73905 1 410
2 73906 1 410
2 73907 1 410
2 73908 1 410
2 73909 1 410
2 73910 1 410
2 73911 1 410
2 73912 1 410
2 73913 1 410
2 73914 1 410
2 73915 1 410
2 73916 1 410
2 73917 1 410
2 73918 1 410
2 73919 1 410
2 73920 1 410
2 73921 1 410
2 73922 1 410
2 73923 1 410
2 73924 1 410
2 73925 1 411
2 73926 1 411
2 73927 1 411
2 73928 1 412
2 73929 1 412
2 73930 1 412
2 73931 1 412
2 73932 1 412
2 73933 1 412
2 73934 1 412
2 73935 1 412
2 73936 1 412
2 73937 1 413
2 73938 1 413
2 73939 1 413
2 73940 1 413
2 73941 1 413
2 73942 1 413
2 73943 1 413
2 73944 1 413
2 73945 1 413
2 73946 1 413
2 73947 1 413
2 73948 1 413
2 73949 1 413
2 73950 1 413
2 73951 1 413
2 73952 1 413
2 73953 1 413
2 73954 1 413
2 73955 1 413
2 73956 1 414
2 73957 1 414
2 73958 1 414
2 73959 1 414
2 73960 1 414
2 73961 1 414
2 73962 1 414
2 73963 1 414
2 73964 1 414
2 73965 1 414
2 73966 1 414
2 73967 1 414
2 73968 1 415
2 73969 1 415
2 73970 1 416
2 73971 1 416
2 73972 1 416
2 73973 1 416
2 73974 1 416
2 73975 1 418
2 73976 1 418
2 73977 1 419
2 73978 1 419
2 73979 1 419
2 73980 1 426
2 73981 1 426
2 73982 1 426
2 73983 1 426
2 73984 1 426
2 73985 1 426
2 73986 1 426
2 73987 1 426
2 73988 1 426
2 73989 1 426
2 73990 1 426
2 73991 1 426
2 73992 1 426
2 73993 1 426
2 73994 1 426
2 73995 1 426
2 73996 1 426
2 73997 1 426
2 73998 1 427
2 73999 1 427
2 74000 1 427
2 74001 1 427
2 74002 1 427
2 74003 1 427
2 74004 1 428
2 74005 1 428
2 74006 1 428
2 74007 1 428
2 74008 1 428
2 74009 1 428
2 74010 1 428
2 74011 1 428
2 74012 1 429
2 74013 1 429
2 74014 1 429
2 74015 1 429
2 74016 1 431
2 74017 1 431
2 74018 1 432
2 74019 1 432
2 74020 1 443
2 74021 1 443
2 74022 1 443
2 74023 1 443
2 74024 1 443
2 74025 1 443
2 74026 1 443
2 74027 1 443
2 74028 1 443
2 74029 1 443
2 74030 1 443
2 74031 1 443
2 74032 1 443
2 74033 1 443
2 74034 1 443
2 74035 1 443
2 74036 1 443
2 74037 1 443
2 74038 1 443
2 74039 1 443
2 74040 1 443
2 74041 1 443
2 74042 1 443
2 74043 1 444
2 74044 1 444
2 74045 1 444
2 74046 1 444
2 74047 1 445
2 74048 1 445
2 74049 1 445
2 74050 1 445
2 74051 1 445
2 74052 1 446
2 74053 1 446
2 74054 1 446
2 74055 1 446
2 74056 1 446
2 74057 1 446
2 74058 1 447
2 74059 1 447
2 74060 1 447
2 74061 1 447
2 74062 1 447
2 74063 1 447
2 74064 1 447
2 74065 1 447
2 74066 1 447
2 74067 1 447
2 74068 1 447
2 74069 1 447
2 74070 1 447
2 74071 1 447
2 74072 1 447
2 74073 1 447
2 74074 1 447
2 74075 1 447
2 74076 1 447
2 74077 1 447
2 74078 1 447
2 74079 1 447
2 74080 1 447
2 74081 1 447
2 74082 1 447
2 74083 1 447
2 74084 1 447
2 74085 1 447
2 74086 1 447
2 74087 1 447
2 74088 1 447
2 74089 1 447
2 74090 1 447
2 74091 1 447
2 74092 1 447
2 74093 1 447
2 74094 1 447
2 74095 1 447
2 74096 1 447
2 74097 1 447
2 74098 1 448
2 74099 1 448
2 74100 1 448
2 74101 1 448
2 74102 1 448
2 74103 1 448
2 74104 1 448
2 74105 1 448
2 74106 1 448
2 74107 1 448
2 74108 1 448
2 74109 1 448
2 74110 1 448
2 74111 1 448
2 74112 1 448
2 74113 1 448
2 74114 1 448
2 74115 1 448
2 74116 1 448
2 74117 1 448
2 74118 1 448
2 74119 1 448
2 74120 1 448
2 74121 1 448
2 74122 1 448
2 74123 1 448
2 74124 1 448
2 74125 1 448
2 74126 1 448
2 74127 1 448
2 74128 1 448
2 74129 1 448
2 74130 1 448
2 74131 1 448
2 74132 1 448
2 74133 1 448
2 74134 1 448
2 74135 1 449
2 74136 1 449
2 74137 1 449
2 74138 1 449
2 74139 1 449
2 74140 1 449
2 74141 1 450
2 74142 1 450
2 74143 1 450
2 74144 1 450
2 74145 1 450
2 74146 1 455
2 74147 1 455
2 74148 1 455
2 74149 1 455
2 74150 1 455
2 74151 1 455
2 74152 1 455
2 74153 1 455
2 74154 1 455
2 74155 1 455
2 74156 1 455
2 74157 1 455
2 74158 1 455
2 74159 1 455
2 74160 1 455
2 74161 1 455
2 74162 1 455
2 74163 1 455
2 74164 1 456
2 74165 1 456
2 74166 1 456
2 74167 1 456
2 74168 1 465
2 74169 1 465
2 74170 1 465
2 74171 1 465
2 74172 1 465
2 74173 1 465
2 74174 1 465
2 74175 1 465
2 74176 1 465
2 74177 1 465
2 74178 1 465
2 74179 1 465
2 74180 1 465
2 74181 1 465
2 74182 1 465
2 74183 1 465
2 74184 1 465
2 74185 1 465
2 74186 1 465
2 74187 1 465
2 74188 1 465
2 74189 1 465
2 74190 1 465
2 74191 1 466
2 74192 1 466
2 74193 1 466
2 74194 1 467
2 74195 1 467
2 74196 1 467
2 74197 1 467
2 74198 1 467
2 74199 1 467
2 74200 1 467
2 74201 1 467
2 74202 1 467
2 74203 1 467
2 74204 1 467
2 74205 1 467
2 74206 1 467
2 74207 1 468
2 74208 1 468
2 74209 1 468
2 74210 1 469
2 74211 1 469
2 74212 1 469
2 74213 1 469
2 74214 1 469
2 74215 1 469
2 74216 1 469
2 74217 1 469
2 74218 1 469
2 74219 1 469
2 74220 1 469
2 74221 1 469
2 74222 1 469
2 74223 1 469
2 74224 1 469
2 74225 1 469
2 74226 1 469
2 74227 1 469
2 74228 1 469
2 74229 1 469
2 74230 1 469
2 74231 1 470
2 74232 1 470
2 74233 1 470
2 74234 1 470
2 74235 1 470
2 74236 1 470
2 74237 1 470
2 74238 1 470
2 74239 1 470
2 74240 1 470
2 74241 1 470
2 74242 1 470
2 74243 1 471
2 74244 1 471
2 74245 1 472
2 74246 1 472
2 74247 1 472
2 74248 1 472
2 74249 1 472
2 74250 1 472
2 74251 1 472
2 74252 1 472
2 74253 1 473
2 74254 1 473
2 74255 1 473
2 74256 1 473
2 74257 1 473
2 74258 1 473
2 74259 1 473
2 74260 1 473
2 74261 1 473
2 74262 1 473
2 74263 1 473
2 74264 1 473
2 74265 1 473
2 74266 1 473
2 74267 1 473
2 74268 1 473
2 74269 1 473
2 74270 1 473
2 74271 1 473
2 74272 1 473
2 74273 1 473
2 74274 1 473
2 74275 1 473
2 74276 1 473
2 74277 1 473
2 74278 1 473
2 74279 1 473
2 74280 1 473
2 74281 1 473
2 74282 1 474
2 74283 1 474
2 74284 1 475
2 74285 1 475
2 74286 1 475
2 74287 1 475
2 74288 1 475
2 74289 1 475
2 74290 1 475
2 74291 1 475
2 74292 1 475
2 74293 1 475
2 74294 1 475
2 74295 1 476
2 74296 1 476
2 74297 1 484
2 74298 1 484
2 74299 1 484
2 74300 1 484
2 74301 1 484
2 74302 1 484
2 74303 1 484
2 74304 1 484
2 74305 1 484
2 74306 1 484
2 74307 1 484
2 74308 1 484
2 74309 1 484
2 74310 1 484
2 74311 1 484
2 74312 1 484
2 74313 1 484
2 74314 1 484
2 74315 1 484
2 74316 1 484
2 74317 1 484
2 74318 1 484
2 74319 1 484
2 74320 1 484
2 74321 1 484
2 74322 1 484
2 74323 1 484
2 74324 1 484
2 74325 1 484
2 74326 1 484
2 74327 1 484
2 74328 1 484
2 74329 1 484
2 74330 1 484
2 74331 1 484
2 74332 1 484
2 74333 1 484
2 74334 1 484
2 74335 1 484
2 74336 1 484
2 74337 1 484
2 74338 1 484
2 74339 1 484
2 74340 1 484
2 74341 1 484
2 74342 1 485
2 74343 1 485
2 74344 1 485
2 74345 1 485
2 74346 1 485
2 74347 1 485
2 74348 1 485
2 74349 1 485
2 74350 1 485
2 74351 1 485
2 74352 1 485
2 74353 1 485
2 74354 1 485
2 74355 1 485
2 74356 1 485
2 74357 1 485
2 74358 1 485
2 74359 1 485
2 74360 1 485
2 74361 1 485
2 74362 1 485
2 74363 1 485
2 74364 1 485
2 74365 1 485
2 74366 1 485
2 74367 1 485
2 74368 1 485
2 74369 1 485
2 74370 1 485
2 74371 1 485
2 74372 1 485
2 74373 1 485
2 74374 1 485
2 74375 1 485
2 74376 1 485
2 74377 1 485
2 74378 1 485
2 74379 1 485
2 74380 1 485
2 74381 1 485
2 74382 1 485
2 74383 1 485
2 74384 1 485
2 74385 1 485
2 74386 1 485
2 74387 1 485
2 74388 1 485
2 74389 1 485
2 74390 1 486
2 74391 1 486
2 74392 1 486
2 74393 1 486
2 74394 1 489
2 74395 1 489
2 74396 1 489
2 74397 1 489
2 74398 1 489
2 74399 1 489
2 74400 1 489
2 74401 1 489
2 74402 1 489
2 74403 1 489
2 74404 1 489
2 74405 1 489
2 74406 1 489
2 74407 1 489
2 74408 1 489
2 74409 1 490
2 74410 1 490
2 74411 1 495
2 74412 1 495
2 74413 1 496
2 74414 1 496
2 74415 1 496
2 74416 1 496
2 74417 1 496
2 74418 1 496
2 74419 1 496
2 74420 1 496
2 74421 1 496
2 74422 1 499
2 74423 1 499
2 74424 1 499
2 74425 1 499
2 74426 1 499
2 74427 1 499
2 74428 1 499
2 74429 1 499
2 74430 1 499
2 74431 1 499
2 74432 1 499
2 74433 1 499
2 74434 1 499
2 74435 1 499
2 74436 1 499
2 74437 1 499
2 74438 1 499
2 74439 1 499
2 74440 1 499
2 74441 1 499
2 74442 1 499
2 74443 1 499
2 74444 1 499
2 74445 1 505
2 74446 1 505
2 74447 1 505
2 74448 1 505
2 74449 1 505
2 74450 1 505
2 74451 1 505
2 74452 1 505
2 74453 1 505
2 74454 1 505
2 74455 1 505
2 74456 1 505
2 74457 1 505
2 74458 1 505
2 74459 1 514
2 74460 1 514
2 74461 1 514
2 74462 1 514
2 74463 1 514
2 74464 1 514
2 74465 1 514
2 74466 1 514
2 74467 1 514
2 74468 1 514
2 74469 1 514
2 74470 1 514
2 74471 1 514
2 74472 1 514
2 74473 1 514
2 74474 1 514
2 74475 1 514
2 74476 1 515
2 74477 1 515
2 74478 1 515
2 74479 1 515
2 74480 1 516
2 74481 1 516
2 74482 1 516
2 74483 1 517
2 74484 1 517
2 74485 1 518
2 74486 1 518
2 74487 1 518
2 74488 1 518
2 74489 1 518
2 74490 1 518
2 74491 1 518
2 74492 1 518
2 74493 1 518
2 74494 1 518
2 74495 1 518
2 74496 1 518
2 74497 1 518
2 74498 1 519
2 74499 1 519
2 74500 1 527
2 74501 1 527
2 74502 1 527
2 74503 1 527
2 74504 1 528
2 74505 1 528
2 74506 1 528
2 74507 1 528
2 74508 1 528
2 74509 1 529
2 74510 1 529
2 74511 1 529
2 74512 1 529
2 74513 1 529
2 74514 1 529
2 74515 1 529
2 74516 1 530
2 74517 1 530
2 74518 1 530
2 74519 1 530
2 74520 1 530
2 74521 1 530
2 74522 1 532
2 74523 1 532
2 74524 1 532
2 74525 1 532
2 74526 1 532
2 74527 1 533
2 74528 1 533
2 74529 1 533
2 74530 1 533
2 74531 1 533
2 74532 1 533
2 74533 1 533
2 74534 1 533
2 74535 1 535
2 74536 1 535
2 74537 1 536
2 74538 1 536
2 74539 1 536
2 74540 1 536
2 74541 1 536
2 74542 1 536
2 74543 1 536
2 74544 1 536
2 74545 1 536
2 74546 1 536
2 74547 1 536
2 74548 1 536
2 74549 1 536
2 74550 1 536
2 74551 1 536
2 74552 1 536
2 74553 1 536
2 74554 1 536
2 74555 1 537
2 74556 1 537
2 74557 1 537
2 74558 1 538
2 74559 1 538
2 74560 1 539
2 74561 1 539
2 74562 1 539
2 74563 1 539
2 74564 1 539
2 74565 1 539
2 74566 1 539
2 74567 1 539
2 74568 1 539
2 74569 1 539
2 74570 1 539
2 74571 1 539
2 74572 1 539
2 74573 1 540
2 74574 1 540
2 74575 1 540
2 74576 1 540
2 74577 1 540
2 74578 1 540
2 74579 1 540
2 74580 1 540
2 74581 1 540
2 74582 1 540
2 74583 1 540
2 74584 1 540
2 74585 1 540
2 74586 1 540
2 74587 1 541
2 74588 1 541
2 74589 1 544
2 74590 1 544
2 74591 1 544
2 74592 1 544
2 74593 1 544
2 74594 1 544
2 74595 1 544
2 74596 1 547
2 74597 1 547
2 74598 1 547
2 74599 1 547
2 74600 1 547
2 74601 1 547
2 74602 1 547
2 74603 1 547
2 74604 1 547
2 74605 1 547
2 74606 1 547
2 74607 1 549
2 74608 1 549
2 74609 1 549
2 74610 1 549
2 74611 1 549
2 74612 1 549
2 74613 1 549
2 74614 1 549
2 74615 1 549
2 74616 1 549
2 74617 1 549
2 74618 1 549
2 74619 1 549
2 74620 1 549
2 74621 1 549
2 74622 1 549
2 74623 1 549
2 74624 1 549
2 74625 1 549
2 74626 1 549
2 74627 1 549
2 74628 1 549
2 74629 1 549
2 74630 1 549
2 74631 1 549
2 74632 1 549
2 74633 1 550
2 74634 1 550
2 74635 1 550
2 74636 1 550
2 74637 1 551
2 74638 1 551
2 74639 1 551
2 74640 1 551
2 74641 1 551
2 74642 1 551
2 74643 1 554
2 74644 1 554
2 74645 1 559
2 74646 1 559
2 74647 1 559
2 74648 1 559
2 74649 1 559
2 74650 1 559
2 74651 1 559
2 74652 1 559
2 74653 1 559
2 74654 1 559
2 74655 1 559
2 74656 1 559
2 74657 1 559
2 74658 1 559
2 74659 1 559
2 74660 1 559
2 74661 1 559
2 74662 1 559
2 74663 1 559
2 74664 1 559
2 74665 1 559
2 74666 1 559
2 74667 1 559
2 74668 1 560
2 74669 1 560
2 74670 1 560
2 74671 1 561
2 74672 1 561
2 74673 1 561
2 74674 1 561
2 74675 1 561
2 74676 1 561
2 74677 1 561
2 74678 1 561
2 74679 1 561
2 74680 1 561
2 74681 1 561
2 74682 1 561
2 74683 1 561
2 74684 1 561
2 74685 1 562
2 74686 1 562
2 74687 1 563
2 74688 1 563
2 74689 1 563
2 74690 1 564
2 74691 1 564
2 74692 1 573
2 74693 1 573
2 74694 1 573
2 74695 1 574
2 74696 1 574
2 74697 1 575
2 74698 1 575
2 74699 1 575
2 74700 1 575
2 74701 1 575
2 74702 1 575
2 74703 1 575
2 74704 1 575
2 74705 1 575
2 74706 1 575
2 74707 1 575
2 74708 1 575
2 74709 1 575
2 74710 1 575
2 74711 1 575
2 74712 1 575
2 74713 1 576
2 74714 1 576
2 74715 1 576
2 74716 1 577
2 74717 1 577
2 74718 1 577
2 74719 1 583
2 74720 1 583
2 74721 1 584
2 74722 1 584
2 74723 1 584
2 74724 1 584
2 74725 1 584
2 74726 1 584
2 74727 1 584
2 74728 1 584
2 74729 1 585
2 74730 1 585
2 74731 1 585
2 74732 1 585
2 74733 1 585
2 74734 1 585
2 74735 1 585
2 74736 1 585
2 74737 1 585
2 74738 1 586
2 74739 1 586
2 74740 1 587
2 74741 1 587
2 74742 1 588
2 74743 1 588
2 74744 1 590
2 74745 1 590
2 74746 1 590
2 74747 1 590
2 74748 1 590
2 74749 1 590
2 74750 1 590
2 74751 1 590
2 74752 1 590
2 74753 1 590
2 74754 1 590
2 74755 1 591
2 74756 1 591
2 74757 1 591
2 74758 1 591
2 74759 1 591
2 74760 1 591
2 74761 1 591
2 74762 1 591
2 74763 1 591
2 74764 1 591
2 74765 1 591
2 74766 1 591
2 74767 1 591
2 74768 1 591
2 74769 1 591
2 74770 1 591
2 74771 1 591
2 74772 1 591
2 74773 1 591
2 74774 1 591
2 74775 1 591
2 74776 1 591
2 74777 1 591
2 74778 1 591
2 74779 1 591
2 74780 1 591
2 74781 1 591
2 74782 1 591
2 74783 1 591
2 74784 1 591
2 74785 1 591
2 74786 1 591
2 74787 1 591
2 74788 1 591
2 74789 1 591
2 74790 1 591
2 74791 1 591
2 74792 1 591
2 74793 1 591
2 74794 1 591
2 74795 1 591
2 74796 1 591
2 74797 1 591
2 74798 1 591
2 74799 1 591
2 74800 1 591
2 74801 1 591
2 74802 1 591
2 74803 1 591
2 74804 1 591
2 74805 1 591
2 74806 1 591
2 74807 1 591
2 74808 1 591
2 74809 1 591
2 74810 1 591
2 74811 1 591
2 74812 1 591
2 74813 1 591
2 74814 1 591
2 74815 1 591
2 74816 1 591
2 74817 1 591
2 74818 1 591
2 74819 1 591
2 74820 1 591
2 74821 1 591
2 74822 1 591
2 74823 1 591
2 74824 1 591
2 74825 1 591
2 74826 1 591
2 74827 1 591
2 74828 1 591
2 74829 1 591
2 74830 1 592
2 74831 1 592
2 74832 1 592
2 74833 1 592
2 74834 1 592
2 74835 1 592
2 74836 1 592
2 74837 1 592
2 74838 1 592
2 74839 1 592
2 74840 1 592
2 74841 1 592
2 74842 1 592
2 74843 1 592
2 74844 1 592
2 74845 1 592
2 74846 1 592
2 74847 1 592
2 74848 1 592
2 74849 1 592
2 74850 1 592
2 74851 1 592
2 74852 1 594
2 74853 1 594
2 74854 1 594
2 74855 1 594
2 74856 1 594
2 74857 1 594
2 74858 1 594
2 74859 1 594
2 74860 1 594
2 74861 1 594
2 74862 1 594
2 74863 1 594
2 74864 1 594
2 74865 1 594
2 74866 1 594
2 74867 1 594
2 74868 1 594
2 74869 1 594
2 74870 1 594
2 74871 1 594
2 74872 1 595
2 74873 1 595
2 74874 1 599
2 74875 1 599
2 74876 1 599
2 74877 1 599
2 74878 1 599
2 74879 1 599
2 74880 1 599
2 74881 1 599
2 74882 1 599
2 74883 1 599
2 74884 1 599
2 74885 1 599
2 74886 1 599
2 74887 1 599
2 74888 1 599
2 74889 1 599
2 74890 1 599
2 74891 1 599
2 74892 1 599
2 74893 1 599
2 74894 1 599
2 74895 1 600
2 74896 1 600
2 74897 1 600
2 74898 1 600
2 74899 1 600
2 74900 1 601
2 74901 1 601
2 74902 1 601
2 74903 1 601
2 74904 1 601
2 74905 1 601
2 74906 1 602
2 74907 1 602
2 74908 1 602
2 74909 1 603
2 74910 1 603
2 74911 1 604
2 74912 1 604
2 74913 1 604
2 74914 1 604
2 74915 1 604
2 74916 1 604
2 74917 1 604
2 74918 1 605
2 74919 1 605
2 74920 1 605
2 74921 1 605
2 74922 1 605
2 74923 1 605
2 74924 1 605
2 74925 1 605
2 74926 1 605
2 74927 1 605
2 74928 1 605
2 74929 1 605
2 74930 1 613
2 74931 1 613
2 74932 1 613
2 74933 1 613
2 74934 1 613
2 74935 1 613
2 74936 1 613
2 74937 1 613
2 74938 1 613
2 74939 1 613
2 74940 1 613
2 74941 1 613
2 74942 1 613
2 74943 1 615
2 74944 1 615
2 74945 1 615
2 74946 1 622
2 74947 1 622
2 74948 1 622
2 74949 1 622
2 74950 1 622
2 74951 1 622
2 74952 1 622
2 74953 1 622
2 74954 1 622
2 74955 1 622
2 74956 1 624
2 74957 1 624
2 74958 1 625
2 74959 1 625
2 74960 1 638
2 74961 1 638
2 74962 1 638
2 74963 1 638
2 74964 1 638
2 74965 1 638
2 74966 1 638
2 74967 1 638
2 74968 1 638
2 74969 1 638
2 74970 1 638
2 74971 1 638
2 74972 1 638
2 74973 1 638
2 74974 1 638
2 74975 1 638
2 74976 1 638
2 74977 1 639
2 74978 1 639
2 74979 1 639
2 74980 1 639
2 74981 1 639
2 74982 1 639
2 74983 1 639
2 74984 1 639
2 74985 1 639
2 74986 1 639
2 74987 1 639
2 74988 1 639
2 74989 1 639
2 74990 1 639
2 74991 1 639
2 74992 1 639
2 74993 1 639
2 74994 1 639
2 74995 1 639
2 74996 1 640
2 74997 1 640
2 74998 1 640
2 74999 1 640
2 75000 1 640
2 75001 1 640
2 75002 1 640
2 75003 1 641
2 75004 1 641
2 75005 1 642
2 75006 1 642
2 75007 1 649
2 75008 1 649
2 75009 1 649
2 75010 1 649
2 75011 1 649
2 75012 1 649
2 75013 1 649
2 75014 1 657
2 75015 1 657
2 75016 1 657
2 75017 1 657
2 75018 1 658
2 75019 1 658
2 75020 1 658
2 75021 1 658
2 75022 1 658
2 75023 1 658
2 75024 1 658
2 75025 1 658
2 75026 1 658
2 75027 1 658
2 75028 1 658
2 75029 1 658
2 75030 1 658
2 75031 1 658
2 75032 1 658
2 75033 1 658
2 75034 1 658
2 75035 1 658
2 75036 1 658
2 75037 1 658
2 75038 1 658
2 75039 1 658
2 75040 1 660
2 75041 1 660
2 75042 1 667
2 75043 1 667
2 75044 1 667
2 75045 1 667
2 75046 1 667
2 75047 1 667
2 75048 1 667
2 75049 1 667
2 75050 1 667
2 75051 1 667
2 75052 1 667
2 75053 1 667
2 75054 1 667
2 75055 1 667
2 75056 1 667
2 75057 1 667
2 75058 1 669
2 75059 1 669
2 75060 1 673
2 75061 1 673
2 75062 1 673
2 75063 1 673
2 75064 1 674
2 75065 1 674
2 75066 1 674
2 75067 1 684
2 75068 1 684
2 75069 1 684
2 75070 1 684
2 75071 1 684
2 75072 1 684
2 75073 1 684
2 75074 1 684
2 75075 1 684
2 75076 1 684
2 75077 1 686
2 75078 1 686
2 75079 1 687
2 75080 1 687
2 75081 1 687
2 75082 1 688
2 75083 1 688
2 75084 1 697
2 75085 1 697
2 75086 1 697
2 75087 1 697
2 75088 1 697
2 75089 1 697
2 75090 1 697
2 75091 1 697
2 75092 1 697
2 75093 1 697
2 75094 1 697
2 75095 1 697
2 75096 1 697
2 75097 1 697
2 75098 1 697
2 75099 1 697
2 75100 1 697
2 75101 1 697
2 75102 1 699
2 75103 1 699
2 75104 1 699
2 75105 1 699
2 75106 1 699
2 75107 1 699
2 75108 1 699
2 75109 1 699
2 75110 1 699
2 75111 1 699
2 75112 1 699
2 75113 1 699
2 75114 1 699
2 75115 1 699
2 75116 1 699
2 75117 1 700
2 75118 1 700
2 75119 1 700
2 75120 1 701
2 75121 1 701
2 75122 1 701
2 75123 1 701
2 75124 1 702
2 75125 1 702
2 75126 1 702
2 75127 1 702
2 75128 1 702
2 75129 1 702
2 75130 1 702
2 75131 1 702
2 75132 1 702
2 75133 1 702
2 75134 1 702
2 75135 1 702
2 75136 1 702
2 75137 1 702
2 75138 1 702
2 75139 1 702
2 75140 1 702
2 75141 1 702
2 75142 1 702
2 75143 1 702
2 75144 1 702
2 75145 1 702
2 75146 1 702
2 75147 1 702
2 75148 1 702
2 75149 1 702
2 75150 1 702
2 75151 1 702
2 75152 1 702
2 75153 1 702
2 75154 1 702
2 75155 1 702
2 75156 1 702
2 75157 1 702
2 75158 1 702
2 75159 1 702
2 75160 1 702
2 75161 1 702
2 75162 1 702
2 75163 1 702
2 75164 1 702
2 75165 1 702
2 75166 1 702
2 75167 1 702
2 75168 1 702
2 75169 1 702
2 75170 1 702
2 75171 1 702
2 75172 1 702
2 75173 1 702
2 75174 1 702
2 75175 1 702
2 75176 1 703
2 75177 1 703
2 75178 1 703
2 75179 1 703
2 75180 1 703
2 75181 1 703
2 75182 1 703
2 75183 1 703
2 75184 1 703
2 75185 1 703
2 75186 1 703
2 75187 1 703
2 75188 1 703
2 75189 1 710
2 75190 1 710
2 75191 1 710
2 75192 1 710
2 75193 1 710
2 75194 1 717
2 75195 1 717
2 75196 1 717
2 75197 1 717
2 75198 1 717
2 75199 1 717
2 75200 1 717
2 75201 1 718
2 75202 1 718
2 75203 1 718
2 75204 1 718
2 75205 1 719
2 75206 1 719
2 75207 1 719
2 75208 1 721
2 75209 1 721
2 75210 1 721
2 75211 1 721
2 75212 1 721
2 75213 1 728
2 75214 1 728
2 75215 1 728
2 75216 1 728
2 75217 1 728
2 75218 1 728
2 75219 1 728
2 75220 1 728
2 75221 1 728
2 75222 1 728
2 75223 1 728
2 75224 1 728
2 75225 1 728
2 75226 1 729
2 75227 1 729
2 75228 1 729
2 75229 1 740
2 75230 1 740
2 75231 1 740
2 75232 1 740
2 75233 1 740
2 75234 1 740
2 75235 1 740
2 75236 1 740
2 75237 1 740
2 75238 1 740
2 75239 1 741
2 75240 1 741
2 75241 1 742
2 75242 1 742
2 75243 1 742
2 75244 1 742
2 75245 1 742
2 75246 1 742
2 75247 1 750
2 75248 1 750
2 75249 1 750
2 75250 1 750
2 75251 1 750
2 75252 1 750
2 75253 1 750
2 75254 1 750
2 75255 1 750
2 75256 1 750
2 75257 1 750
2 75258 1 750
2 75259 1 750
2 75260 1 751
2 75261 1 751
2 75262 1 751
2 75263 1 751
2 75264 1 751
2 75265 1 751
2 75266 1 752
2 75267 1 752
2 75268 1 752
2 75269 1 752
2 75270 1 752
2 75271 1 752
2 75272 1 752
2 75273 1 752
2 75274 1 752
2 75275 1 753
2 75276 1 753
2 75277 1 753
2 75278 1 754
2 75279 1 754
2 75280 1 754
2 75281 1 754
2 75282 1 754
2 75283 1 754
2 75284 1 754
2 75285 1 754
2 75286 1 754
2 75287 1 754
2 75288 1 754
2 75289 1 754
2 75290 1 754
2 75291 1 754
2 75292 1 754
2 75293 1 754
2 75294 1 754
2 75295 1 754
2 75296 1 754
2 75297 1 755
2 75298 1 755
2 75299 1 758
2 75300 1 758
2 75301 1 767
2 75302 1 767
2 75303 1 767
2 75304 1 767
2 75305 1 767
2 75306 1 767
2 75307 1 767
2 75308 1 767
2 75309 1 767
2 75310 1 767
2 75311 1 768
2 75312 1 768
2 75313 1 769
2 75314 1 769
2 75315 1 769
2 75316 1 769
2 75317 1 769
2 75318 1 769
2 75319 1 769
2 75320 1 769
2 75321 1 769
2 75322 1 769
2 75323 1 769
2 75324 1 769
2 75325 1 769
2 75326 1 769
2 75327 1 769
2 75328 1 769
2 75329 1 769
2 75330 1 769
2 75331 1 770
2 75332 1 770
2 75333 1 773
2 75334 1 773
2 75335 1 773
2 75336 1 773
2 75337 1 778
2 75338 1 778
2 75339 1 778
2 75340 1 778
2 75341 1 778
2 75342 1 778
2 75343 1 778
2 75344 1 778
2 75345 1 796
2 75346 1 796
2 75347 1 796
2 75348 1 796
2 75349 1 796
2 75350 1 796
2 75351 1 796
2 75352 1 796
2 75353 1 796
2 75354 1 796
2 75355 1 796
2 75356 1 796
2 75357 1 797
2 75358 1 797
2 75359 1 797
2 75360 1 797
2 75361 1 798
2 75362 1 798
2 75363 1 798
2 75364 1 798
2 75365 1 799
2 75366 1 799
2 75367 1 799
2 75368 1 799
2 75369 1 802
2 75370 1 802
2 75371 1 802
2 75372 1 802
2 75373 1 802
2 75374 1 802
2 75375 1 802
2 75376 1 802
2 75377 1 804
2 75378 1 804
2 75379 1 804
2 75380 1 804
2 75381 1 804
2 75382 1 804
2 75383 1 806
2 75384 1 806
2 75385 1 806
2 75386 1 809
2 75387 1 809
2 75388 1 809
2 75389 1 809
2 75390 1 809
2 75391 1 816
2 75392 1 816
2 75393 1 816
2 75394 1 816
2 75395 1 816
2 75396 1 816
2 75397 1 816
2 75398 1 816
2 75399 1 816
2 75400 1 816
2 75401 1 816
2 75402 1 816
2 75403 1 816
2 75404 1 816
2 75405 1 816
2 75406 1 816
2 75407 1 816
2 75408 1 816
2 75409 1 816
2 75410 1 816
2 75411 1 816
2 75412 1 816
2 75413 1 816
2 75414 1 816
2 75415 1 816
2 75416 1 816
2 75417 1 816
2 75418 1 816
2 75419 1 816
2 75420 1 816
2 75421 1 816
2 75422 1 816
2 75423 1 816
2 75424 1 816
2 75425 1 816
2 75426 1 816
2 75427 1 816
2 75428 1 816
2 75429 1 817
2 75430 1 817
2 75431 1 817
2 75432 1 817
2 75433 1 817
2 75434 1 817
2 75435 1 817
2 75436 1 818
2 75437 1 818
2 75438 1 818
2 75439 1 819
2 75440 1 819
2 75441 1 821
2 75442 1 821
2 75443 1 839
2 75444 1 839
2 75445 1 839
2 75446 1 839
2 75447 1 839
2 75448 1 839
2 75449 1 839
2 75450 1 839
2 75451 1 839
2 75452 1 839
2 75453 1 839
2 75454 1 839
2 75455 1 839
2 75456 1 839
2 75457 1 839
2 75458 1 839
2 75459 1 841
2 75460 1 841
2 75461 1 841
2 75462 1 842
2 75463 1 842
2 75464 1 842
2 75465 1 842
2 75466 1 842
2 75467 1 842
2 75468 1 842
2 75469 1 842
2 75470 1 842
2 75471 1 842
2 75472 1 842
2 75473 1 842
2 75474 1 842
2 75475 1 842
2 75476 1 842
2 75477 1 842
2 75478 1 842
2 75479 1 842
2 75480 1 842
2 75481 1 842
2 75482 1 842
2 75483 1 842
2 75484 1 842
2 75485 1 842
2 75486 1 842
2 75487 1 842
2 75488 1 842
2 75489 1 842
2 75490 1 842
2 75491 1 843
2 75492 1 843
2 75493 1 846
2 75494 1 846
2 75495 1 846
2 75496 1 846
2 75497 1 847
2 75498 1 847
2 75499 1 847
2 75500 1 847
2 75501 1 849
2 75502 1 849
2 75503 1 849
2 75504 1 849
2 75505 1 849
2 75506 1 849
2 75507 1 849
2 75508 1 849
2 75509 1 849
2 75510 1 849
2 75511 1 849
2 75512 1 849
2 75513 1 849
2 75514 1 849
2 75515 1 849
2 75516 1 849
2 75517 1 849
2 75518 1 849
2 75519 1 851
2 75520 1 851
2 75521 1 851
2 75522 1 851
2 75523 1 851
2 75524 1 851
2 75525 1 851
2 75526 1 851
2 75527 1 851
2 75528 1 851
2 75529 1 851
2 75530 1 851
2 75531 1 851
2 75532 1 851
2 75533 1 851
2 75534 1 851
2 75535 1 851
2 75536 1 852
2 75537 1 852
2 75538 1 852
2 75539 1 852
2 75540 1 852
2 75541 1 852
2 75542 1 852
2 75543 1 852
2 75544 1 852
2 75545 1 852
2 75546 1 852
2 75547 1 852
2 75548 1 852
2 75549 1 852
2 75550 1 852
2 75551 1 852
2 75552 1 852
2 75553 1 852
2 75554 1 852
2 75555 1 852
2 75556 1 852
2 75557 1 852
2 75558 1 852
2 75559 1 852
2 75560 1 852
2 75561 1 854
2 75562 1 854
2 75563 1 867
2 75564 1 867
2 75565 1 867
2 75566 1 868
2 75567 1 868
2 75568 1 869
2 75569 1 869
2 75570 1 869
2 75571 1 869
2 75572 1 869
2 75573 1 869
2 75574 1 869
2 75575 1 869
2 75576 1 869
2 75577 1 869
2 75578 1 869
2 75579 1 869
2 75580 1 870
2 75581 1 870
2 75582 1 870
2 75583 1 871
2 75584 1 871
2 75585 1 871
2 75586 1 879
2 75587 1 879
2 75588 1 881
2 75589 1 881
2 75590 1 881
2 75591 1 881
2 75592 1 881
2 75593 1 881
2 75594 1 881
2 75595 1 881
2 75596 1 881
2 75597 1 881
2 75598 1 881
2 75599 1 881
2 75600 1 881
2 75601 1 881
2 75602 1 882
2 75603 1 882
2 75604 1 883
2 75605 1 883
2 75606 1 886
2 75607 1 886
2 75608 1 886
2 75609 1 886
2 75610 1 890
2 75611 1 890
2 75612 1 890
2 75613 1 890
2 75614 1 890
2 75615 1 892
2 75616 1 892
2 75617 1 901
2 75618 1 901
2 75619 1 901
2 75620 1 901
2 75621 1 901
2 75622 1 901
2 75623 1 901
2 75624 1 901
2 75625 1 901
2 75626 1 901
2 75627 1 902
2 75628 1 902
2 75629 1 903
2 75630 1 903
2 75631 1 903
2 75632 1 904
2 75633 1 904
2 75634 1 904
2 75635 1 904
2 75636 1 905
2 75637 1 905
2 75638 1 905
2 75639 1 905
2 75640 1 905
2 75641 1 905
2 75642 1 905
2 75643 1 905
2 75644 1 905
2 75645 1 905
2 75646 1 905
2 75647 1 907
2 75648 1 907
2 75649 1 907
2 75650 1 907
2 75651 1 907
2 75652 1 911
2 75653 1 911
2 75654 1 911
2 75655 1 911
2 75656 1 911
2 75657 1 911
2 75658 1 912
2 75659 1 912
2 75660 1 912
2 75661 1 912
2 75662 1 912
2 75663 1 912
2 75664 1 912
2 75665 1 912
2 75666 1 912
2 75667 1 912
2 75668 1 912
2 75669 1 913
2 75670 1 913
2 75671 1 913
2 75672 1 913
2 75673 1 913
2 75674 1 913
2 75675 1 913
2 75676 1 913
2 75677 1 913
2 75678 1 913
2 75679 1 914
2 75680 1 914
2 75681 1 914
2 75682 1 914
2 75683 1 914
2 75684 1 914
2 75685 1 914
2 75686 1 914
2 75687 1 914
2 75688 1 914
2 75689 1 914
2 75690 1 922
2 75691 1 922
2 75692 1 922
2 75693 1 922
2 75694 1 922
2 75695 1 922
2 75696 1 922
2 75697 1 922
2 75698 1 922
2 75699 1 922
2 75700 1 922
2 75701 1 922
2 75702 1 922
2 75703 1 922
2 75704 1 922
2 75705 1 922
2 75706 1 922
2 75707 1 922
2 75708 1 922
2 75709 1 922
2 75710 1 922
2 75711 1 922
2 75712 1 922
2 75713 1 923
2 75714 1 923
2 75715 1 923
2 75716 1 923
2 75717 1 932
2 75718 1 932
2 75719 1 932
2 75720 1 932
2 75721 1 932
2 75722 1 932
2 75723 1 932
2 75724 1 932
2 75725 1 932
2 75726 1 932
2 75727 1 932
2 75728 1 932
2 75729 1 932
2 75730 1 932
2 75731 1 932
2 75732 1 932
2 75733 1 932
2 75734 1 932
2 75735 1 932
2 75736 1 932
2 75737 1 932
2 75738 1 932
2 75739 1 932
2 75740 1 933
2 75741 1 933
2 75742 1 933
2 75743 1 933
2 75744 1 933
2 75745 1 933
2 75746 1 933
2 75747 1 933
2 75748 1 933
2 75749 1 934
2 75750 1 934
2 75751 1 937
2 75752 1 937
2 75753 1 937
2 75754 1 937
2 75755 1 937
2 75756 1 937
2 75757 1 937
2 75758 1 937
2 75759 1 937
2 75760 1 937
2 75761 1 937
2 75762 1 937
2 75763 1 937
2 75764 1 937
2 75765 1 937
2 75766 1 937
2 75767 1 937
2 75768 1 937
2 75769 1 937
2 75770 1 937
2 75771 1 937
2 75772 1 937
2 75773 1 937
2 75774 1 937
2 75775 1 937
2 75776 1 937
2 75777 1 937
2 75778 1 937
2 75779 1 937
2 75780 1 937
2 75781 1 937
2 75782 1 937
2 75783 1 937
2 75784 1 937
2 75785 1 937
2 75786 1 937
2 75787 1 937
2 75788 1 937
2 75789 1 937
2 75790 1 937
2 75791 1 937
2 75792 1 937
2 75793 1 938
2 75794 1 938
2 75795 1 938
2 75796 1 938
2 75797 1 938
2 75798 1 938
2 75799 1 938
2 75800 1 938
2 75801 1 938
2 75802 1 938
2 75803 1 938
2 75804 1 938
2 75805 1 938
2 75806 1 938
2 75807 1 938
2 75808 1 938
2 75809 1 938
2 75810 1 938
2 75811 1 938
2 75812 1 938
2 75813 1 938
2 75814 1 938
2 75815 1 938
2 75816 1 938
2 75817 1 938
2 75818 1 938
2 75819 1 938
2 75820 1 938
2 75821 1 938
2 75822 1 938
2 75823 1 938
2 75824 1 939
2 75825 1 939
2 75826 1 939
2 75827 1 939
2 75828 1 939
2 75829 1 941
2 75830 1 941
2 75831 1 941
2 75832 1 942
2 75833 1 942
2 75834 1 944
2 75835 1 944
2 75836 1 944
2 75837 1 944
2 75838 1 944
2 75839 1 944
2 75840 1 944
2 75841 1 947
2 75842 1 947
2 75843 1 947
2 75844 1 947
2 75845 1 947
2 75846 1 947
2 75847 1 947
2 75848 1 947
2 75849 1 947
2 75850 1 947
2 75851 1 947
2 75852 1 947
2 75853 1 947
2 75854 1 947
2 75855 1 947
2 75856 1 947
2 75857 1 947
2 75858 1 947
2 75859 1 947
2 75860 1 947
2 75861 1 947
2 75862 1 947
2 75863 1 947
2 75864 1 949
2 75865 1 949
2 75866 1 949
2 75867 1 961
2 75868 1 961
2 75869 1 961
2 75870 1 961
2 75871 1 961
2 75872 1 961
2 75873 1 961
2 75874 1 961
2 75875 1 961
2 75876 1 961
2 75877 1 961
2 75878 1 961
2 75879 1 961
2 75880 1 961
2 75881 1 961
2 75882 1 961
2 75883 1 961
2 75884 1 961
2 75885 1 963
2 75886 1 963
2 75887 1 963
2 75888 1 963
2 75889 1 963
2 75890 1 964
2 75891 1 964
2 75892 1 964
2 75893 1 964
2 75894 1 964
2 75895 1 964
2 75896 1 964
2 75897 1 964
2 75898 1 964
2 75899 1 964
2 75900 1 964
2 75901 1 964
2 75902 1 964
2 75903 1 964
2 75904 1 965
2 75905 1 965
2 75906 1 980
2 75907 1 980
2 75908 1 981
2 75909 1 981
2 75910 1 981
2 75911 1 982
2 75912 1 982
2 75913 1 982
2 75914 1 982
2 75915 1 982
2 75916 1 982
2 75917 1 982
2 75918 1 982
2 75919 1 982
2 75920 1 982
2 75921 1 982
2 75922 1 982
2 75923 1 983
2 75924 1 983
2 75925 1 983
2 75926 1 984
2 75927 1 984
2 75928 1 984
2 75929 1 985
2 75930 1 985
2 75931 1 985
2 75932 1 986
2 75933 1 986
2 75934 1 986
2 75935 1 986
2 75936 1 986
2 75937 1 986
2 75938 1 986
2 75939 1 986
2 75940 1 986
2 75941 1 986
2 75942 1 986
2 75943 1 986
2 75944 1 986
2 75945 1 986
2 75946 1 986
2 75947 1 986
2 75948 1 986
2 75949 1 986
2 75950 1 986
2 75951 1 986
2 75952 1 986
2 75953 1 986
2 75954 1 986
2 75955 1 986
2 75956 1 986
2 75957 1 986
2 75958 1 986
2 75959 1 986
2 75960 1 986
2 75961 1 986
2 75962 1 986
2 75963 1 986
2 75964 1 986
2 75965 1 986
2 75966 1 986
2 75967 1 986
2 75968 1 986
2 75969 1 986
2 75970 1 986
2 75971 1 986
2 75972 1 986
2 75973 1 987
2 75974 1 987
2 75975 1 987
2 75976 1 987
2 75977 1 987
2 75978 1 987
2 75979 1 987
2 75980 1 989
2 75981 1 989
2 75982 1 989
2 75983 1 989
2 75984 1 990
2 75985 1 990
2 75986 1 991
2 75987 1 991
2 75988 1 1003
2 75989 1 1003
2 75990 1 1004
2 75991 1 1004
2 75992 1 1004
2 75993 1 1004
2 75994 1 1004
2 75995 1 1004
2 75996 1 1004
2 75997 1 1004
2 75998 1 1004
2 75999 1 1004
2 76000 1 1004
2 76001 1 1004
2 76002 1 1004
2 76003 1 1004
2 76004 1 1004
2 76005 1 1004
2 76006 1 1004
2 76007 1 1004
2 76008 1 1004
2 76009 1 1004
2 76010 1 1004
2 76011 1 1004
2 76012 1 1004
2 76013 1 1006
2 76014 1 1006
2 76015 1 1006
2 76016 1 1006
2 76017 1 1006
2 76018 1 1007
2 76019 1 1007
2 76020 1 1008
2 76021 1 1008
2 76022 1 1008
2 76023 1 1008
2 76024 1 1008
2 76025 1 1008
2 76026 1 1008
2 76027 1 1008
2 76028 1 1019
2 76029 1 1019
2 76030 1 1019
2 76031 1 1019
2 76032 1 1019
2 76033 1 1019
2 76034 1 1019
2 76035 1 1019
2 76036 1 1019
2 76037 1 1019
2 76038 1 1019
2 76039 1 1019
2 76040 1 1019
2 76041 1 1019
2 76042 1 1019
2 76043 1 1019
2 76044 1 1019
2 76045 1 1019
2 76046 1 1019
2 76047 1 1019
2 76048 1 1019
2 76049 1 1019
2 76050 1 1019
2 76051 1 1019
2 76052 1 1019
2 76053 1 1019
2 76054 1 1019
2 76055 1 1019
2 76056 1 1019
2 76057 1 1019
2 76058 1 1019
2 76059 1 1019
2 76060 1 1019
2 76061 1 1019
2 76062 1 1019
2 76063 1 1021
2 76064 1 1021
2 76065 1 1021
2 76066 1 1021
2 76067 1 1021
2 76068 1 1021
2 76069 1 1021
2 76070 1 1021
2 76071 1 1021
2 76072 1 1021
2 76073 1 1021
2 76074 1 1021
2 76075 1 1021
2 76076 1 1021
2 76077 1 1021
2 76078 1 1021
2 76079 1 1021
2 76080 1 1021
2 76081 1 1021
2 76082 1 1021
2 76083 1 1021
2 76084 1 1021
2 76085 1 1021
2 76086 1 1021
2 76087 1 1021
2 76088 1 1021
2 76089 1 1021
2 76090 1 1021
2 76091 1 1021
2 76092 1 1021
2 76093 1 1021
2 76094 1 1021
2 76095 1 1021
2 76096 1 1021
2 76097 1 1021
2 76098 1 1021
2 76099 1 1021
2 76100 1 1023
2 76101 1 1023
2 76102 1 1023
2 76103 1 1024
2 76104 1 1024
2 76105 1 1024
2 76106 1 1024
2 76107 1 1024
2 76108 1 1024
2 76109 1 1024
2 76110 1 1024
2 76111 1 1024
2 76112 1 1024
2 76113 1 1024
2 76114 1 1024
2 76115 1 1024
2 76116 1 1024
2 76117 1 1024
2 76118 1 1024
2 76119 1 1024
2 76120 1 1024
2 76121 1 1024
2 76122 1 1024
2 76123 1 1024
2 76124 1 1024
2 76125 1 1024
2 76126 1 1024
2 76127 1 1024
2 76128 1 1024
2 76129 1 1024
2 76130 1 1024
2 76131 1 1024
2 76132 1 1024
2 76133 1 1024
2 76134 1 1024
2 76135 1 1024
2 76136 1 1024
2 76137 1 1024
2 76138 1 1024
2 76139 1 1024
2 76140 1 1024
2 76141 1 1024
2 76142 1 1024
2 76143 1 1024
2 76144 1 1024
2 76145 1 1024
2 76146 1 1024
2 76147 1 1024
2 76148 1 1024
2 76149 1 1024
2 76150 1 1024
2 76151 1 1024
2 76152 1 1024
2 76153 1 1024
2 76154 1 1024
2 76155 1 1024
2 76156 1 1024
2 76157 1 1024
2 76158 1 1024
2 76159 1 1024
2 76160 1 1024
2 76161 1 1024
2 76162 1 1024
2 76163 1 1024
2 76164 1 1024
2 76165 1 1024
2 76166 1 1024
2 76167 1 1024
2 76168 1 1024
2 76169 1 1024
2 76170 1 1024
2 76171 1 1024
2 76172 1 1024
2 76173 1 1024
2 76174 1 1024
2 76175 1 1024
2 76176 1 1024
2 76177 1 1024
2 76178 1 1024
2 76179 1 1024
2 76180 1 1024
2 76181 1 1024
2 76182 1 1024
2 76183 1 1024
2 76184 1 1024
2 76185 1 1024
2 76186 1 1024
2 76187 1 1024
2 76188 1 1024
2 76189 1 1024
2 76190 1 1024
2 76191 1 1024
2 76192 1 1024
2 76193 1 1024
2 76194 1 1024
2 76195 1 1024
2 76196 1 1024
2 76197 1 1024
2 76198 1 1024
2 76199 1 1024
2 76200 1 1024
2 76201 1 1025
2 76202 1 1025
2 76203 1 1025
2 76204 1 1025
2 76205 1 1027
2 76206 1 1027
2 76207 1 1027
2 76208 1 1027
2 76209 1 1027
2 76210 1 1027
2 76211 1 1027
2 76212 1 1027
2 76213 1 1027
2 76214 1 1027
2 76215 1 1027
2 76216 1 1028
2 76217 1 1028
2 76218 1 1028
2 76219 1 1029
2 76220 1 1029
2 76221 1 1029
2 76222 1 1029
2 76223 1 1030
2 76224 1 1030
2 76225 1 1030
2 76226 1 1031
2 76227 1 1031
2 76228 1 1031
2 76229 1 1031
2 76230 1 1034
2 76231 1 1034
2 76232 1 1039
2 76233 1 1039
2 76234 1 1039
2 76235 1 1039
2 76236 1 1039
2 76237 1 1039
2 76238 1 1040
2 76239 1 1040
2 76240 1 1040
2 76241 1 1040
2 76242 1 1040
2 76243 1 1040
2 76244 1 1040
2 76245 1 1040
2 76246 1 1040
2 76247 1 1040
2 76248 1 1040
2 76249 1 1040
2 76250 1 1040
2 76251 1 1040
2 76252 1 1040
2 76253 1 1040
2 76254 1 1040
2 76255 1 1040
2 76256 1 1040
2 76257 1 1042
2 76258 1 1042
2 76259 1 1042
2 76260 1 1044
2 76261 1 1044
2 76262 1 1045
2 76263 1 1045
2 76264 1 1046
2 76265 1 1046
2 76266 1 1050
2 76267 1 1050
2 76268 1 1050
2 76269 1 1050
2 76270 1 1050
2 76271 1 1050
2 76272 1 1050
2 76273 1 1050
2 76274 1 1050
2 76275 1 1050
2 76276 1 1050
2 76277 1 1050
2 76278 1 1050
2 76279 1 1050
2 76280 1 1050
2 76281 1 1050
2 76282 1 1050
2 76283 1 1050
2 76284 1 1051
2 76285 1 1051
2 76286 1 1051
2 76287 1 1051
2 76288 1 1062
2 76289 1 1062
2 76290 1 1062
2 76291 1 1062
2 76292 1 1062
2 76293 1 1062
2 76294 1 1062
2 76295 1 1062
2 76296 1 1062
2 76297 1 1063
2 76298 1 1063
2 76299 1 1063
2 76300 1 1063
2 76301 1 1063
2 76302 1 1065
2 76303 1 1065
2 76304 1 1069
2 76305 1 1069
2 76306 1 1069
2 76307 1 1069
2 76308 1 1069
2 76309 1 1069
2 76310 1 1069
2 76311 1 1069
2 76312 1 1069
2 76313 1 1069
2 76314 1 1069
2 76315 1 1069
2 76316 1 1069
2 76317 1 1069
2 76318 1 1069
2 76319 1 1069
2 76320 1 1069
2 76321 1 1069
2 76322 1 1069
2 76323 1 1069
2 76324 1 1069
2 76325 1 1069
2 76326 1 1069
2 76327 1 1069
2 76328 1 1069
2 76329 1 1069
2 76330 1 1069
2 76331 1 1070
2 76332 1 1070
2 76333 1 1070
2 76334 1 1070
2 76335 1 1070
2 76336 1 1070
2 76337 1 1071
2 76338 1 1071
2 76339 1 1071
2 76340 1 1071
2 76341 1 1071
2 76342 1 1071
2 76343 1 1071
2 76344 1 1071
2 76345 1 1071
2 76346 1 1071
2 76347 1 1071
2 76348 1 1071
2 76349 1 1071
2 76350 1 1071
2 76351 1 1071
2 76352 1 1071
2 76353 1 1071
2 76354 1 1072
2 76355 1 1072
2 76356 1 1072
2 76357 1 1072
2 76358 1 1073
2 76359 1 1073
2 76360 1 1073
2 76361 1 1073
2 76362 1 1073
2 76363 1 1073
2 76364 1 1073
2 76365 1 1073
2 76366 1 1073
2 76367 1 1073
2 76368 1 1073
2 76369 1 1073
2 76370 1 1073
2 76371 1 1073
2 76372 1 1073
2 76373 1 1073
2 76374 1 1073
2 76375 1 1073
2 76376 1 1073
2 76377 1 1074
2 76378 1 1074
2 76379 1 1074
2 76380 1 1074
2 76381 1 1074
2 76382 1 1074
2 76383 1 1085
2 76384 1 1085
2 76385 1 1085
2 76386 1 1085
2 76387 1 1085
2 76388 1 1085
2 76389 1 1085
2 76390 1 1085
2 76391 1 1085
2 76392 1 1096
2 76393 1 1096
2 76394 1 1099
2 76395 1 1099
2 76396 1 1099
2 76397 1 1099
2 76398 1 1099
2 76399 1 1099
2 76400 1 1099
2 76401 1 1099
2 76402 1 1099
2 76403 1 1099
2 76404 1 1099
2 76405 1 1099
2 76406 1 1107
2 76407 1 1107
2 76408 1 1108
2 76409 1 1108
2 76410 1 1108
2 76411 1 1108
2 76412 1 1108
2 76413 1 1110
2 76414 1 1110
2 76415 1 1111
2 76416 1 1111
2 76417 1 1111
2 76418 1 1111
2 76419 1 1111
2 76420 1 1113
2 76421 1 1113
2 76422 1 1113
2 76423 1 1113
2 76424 1 1114
2 76425 1 1114
2 76426 1 1114
2 76427 1 1131
2 76428 1 1131
2 76429 1 1131
2 76430 1 1131
2 76431 1 1131
2 76432 1 1131
2 76433 1 1131
2 76434 1 1131
2 76435 1 1131
2 76436 1 1131
2 76437 1 1131
2 76438 1 1139
2 76439 1 1139
2 76440 1 1139
2 76441 1 1139
2 76442 1 1139
2 76443 1 1139
2 76444 1 1139
2 76445 1 1139
2 76446 1 1139
2 76447 1 1139
2 76448 1 1139
2 76449 1 1140
2 76450 1 1140
2 76451 1 1140
2 76452 1 1140
2 76453 1 1140
2 76454 1 1140
2 76455 1 1140
2 76456 1 1140
2 76457 1 1140
2 76458 1 1140
2 76459 1 1140
2 76460 1 1140
2 76461 1 1140
2 76462 1 1140
2 76463 1 1140
2 76464 1 1140
2 76465 1 1140
2 76466 1 1140
2 76467 1 1140
2 76468 1 1140
2 76469 1 1140
2 76470 1 1140
2 76471 1 1140
2 76472 1 1140
2 76473 1 1140
2 76474 1 1141
2 76475 1 1141
2 76476 1 1141
2 76477 1 1141
2 76478 1 1141
2 76479 1 1142
2 76480 1 1142
2 76481 1 1142
2 76482 1 1143
2 76483 1 1143
2 76484 1 1144
2 76485 1 1144
2 76486 1 1145
2 76487 1 1145
2 76488 1 1145
2 76489 1 1145
2 76490 1 1145
2 76491 1 1145
2 76492 1 1146
2 76493 1 1146
2 76494 1 1146
2 76495 1 1146
2 76496 1 1147
2 76497 1 1147
2 76498 1 1151
2 76499 1 1151
2 76500 1 1154
2 76501 1 1154
2 76502 1 1154
2 76503 1 1157
2 76504 1 1157
2 76505 1 1157
2 76506 1 1157
2 76507 1 1157
2 76508 1 1157
2 76509 1 1157
2 76510 1 1158
2 76511 1 1158
2 76512 1 1158
2 76513 1 1161
2 76514 1 1161
2 76515 1 1161
2 76516 1 1162
2 76517 1 1162
2 76518 1 1162
2 76519 1 1162
2 76520 1 1162
2 76521 1 1162
2 76522 1 1162
2 76523 1 1162
2 76524 1 1162
2 76525 1 1162
2 76526 1 1162
2 76527 1 1162
2 76528 1 1162
2 76529 1 1162
2 76530 1 1162
2 76531 1 1163
2 76532 1 1163
2 76533 1 1163
2 76534 1 1163
2 76535 1 1163
2 76536 1 1163
2 76537 1 1163
2 76538 1 1163
2 76539 1 1163
2 76540 1 1163
2 76541 1 1163
2 76542 1 1168
2 76543 1 1168
2 76544 1 1168
2 76545 1 1168
2 76546 1 1168
2 76547 1 1168
2 76548 1 1168
2 76549 1 1168
2 76550 1 1168
2 76551 1 1168
2 76552 1 1168
2 76553 1 1168
2 76554 1 1168
2 76555 1 1168
2 76556 1 1168
2 76557 1 1168
2 76558 1 1168
2 76559 1 1168
2 76560 1 1168
2 76561 1 1168
2 76562 1 1168
2 76563 1 1168
2 76564 1 1168
2 76565 1 1168
2 76566 1 1168
2 76567 1 1168
2 76568 1 1169
2 76569 1 1169
2 76570 1 1169
2 76571 1 1169
2 76572 1 1169
2 76573 1 1169
2 76574 1 1169
2 76575 1 1169
2 76576 1 1169
2 76577 1 1169
2 76578 1 1169
2 76579 1 1169
2 76580 1 1169
2 76581 1 1169
2 76582 1 1170
2 76583 1 1170
2 76584 1 1178
2 76585 1 1178
2 76586 1 1178
2 76587 1 1178
2 76588 1 1178
2 76589 1 1178
2 76590 1 1178
2 76591 1 1178
2 76592 1 1178
2 76593 1 1179
2 76594 1 1179
2 76595 1 1179
2 76596 1 1179
2 76597 1 1179
2 76598 1 1179
2 76599 1 1179
2 76600 1 1179
2 76601 1 1179
2 76602 1 1180
2 76603 1 1180
2 76604 1 1181
2 76605 1 1181
2 76606 1 1181
2 76607 1 1181
2 76608 1 1181
2 76609 1 1182
2 76610 1 1182
2 76611 1 1183
2 76612 1 1183
2 76613 1 1183
2 76614 1 1183
2 76615 1 1183
2 76616 1 1183
2 76617 1 1185
2 76618 1 1185
2 76619 1 1185
2 76620 1 1185
2 76621 1 1185
2 76622 1 1185
2 76623 1 1185
2 76624 1 1185
2 76625 1 1185
2 76626 1 1185
2 76627 1 1186
2 76628 1 1186
2 76629 1 1187
2 76630 1 1187
2 76631 1 1190
2 76632 1 1190
2 76633 1 1190
2 76634 1 1190
2 76635 1 1191
2 76636 1 1191
2 76637 1 1191
2 76638 1 1191
2 76639 1 1191
2 76640 1 1204
2 76641 1 1204
2 76642 1 1204
2 76643 1 1204
2 76644 1 1204
2 76645 1 1204
2 76646 1 1204
2 76647 1 1204
2 76648 1 1204
2 76649 1 1204
2 76650 1 1204
2 76651 1 1204
2 76652 1 1204
2 76653 1 1205
2 76654 1 1205
2 76655 1 1205
2 76656 1 1210
2 76657 1 1210
2 76658 1 1211
2 76659 1 1211
2 76660 1 1211
2 76661 1 1211
2 76662 1 1211
2 76663 1 1211
2 76664 1 1211
2 76665 1 1211
2 76666 1 1211
2 76667 1 1211
2 76668 1 1211
2 76669 1 1211
2 76670 1 1211
2 76671 1 1211
2 76672 1 1211
2 76673 1 1211
2 76674 1 1211
2 76675 1 1211
2 76676 1 1211
2 76677 1 1211
2 76678 1 1211
2 76679 1 1211
2 76680 1 1211
2 76681 1 1215
2 76682 1 1215
2 76683 1 1215
2 76684 1 1215
2 76685 1 1215
2 76686 1 1215
2 76687 1 1215
2 76688 1 1215
2 76689 1 1215
2 76690 1 1215
2 76691 1 1215
2 76692 1 1215
2 76693 1 1215
2 76694 1 1215
2 76695 1 1215
2 76696 1 1215
2 76697 1 1215
2 76698 1 1215
2 76699 1 1215
2 76700 1 1215
2 76701 1 1215
2 76702 1 1215
2 76703 1 1215
2 76704 1 1215
2 76705 1 1215
2 76706 1 1215
2 76707 1 1215
2 76708 1 1215
2 76709 1 1215
2 76710 1 1215
2 76711 1 1215
2 76712 1 1215
2 76713 1 1215
2 76714 1 1215
2 76715 1 1215
2 76716 1 1215
2 76717 1 1215
2 76718 1 1215
2 76719 1 1215
2 76720 1 1215
2 76721 1 1215
2 76722 1 1215
2 76723 1 1215
2 76724 1 1215
2 76725 1 1215
2 76726 1 1215
2 76727 1 1215
2 76728 1 1215
2 76729 1 1215
2 76730 1 1217
2 76731 1 1217
2 76732 1 1217
2 76733 1 1217
2 76734 1 1217
2 76735 1 1217
2 76736 1 1217
2 76737 1 1219
2 76738 1 1219
2 76739 1 1219
2 76740 1 1219
2 76741 1 1219
2 76742 1 1219
2 76743 1 1219
2 76744 1 1219
2 76745 1 1219
2 76746 1 1220
2 76747 1 1220
2 76748 1 1220
2 76749 1 1220
2 76750 1 1221
2 76751 1 1221
2 76752 1 1221
2 76753 1 1221
2 76754 1 1223
2 76755 1 1223
2 76756 1 1224
2 76757 1 1224
2 76758 1 1224
2 76759 1 1224
2 76760 1 1224
2 76761 1 1224
2 76762 1 1224
2 76763 1 1224
2 76764 1 1224
2 76765 1 1224
2 76766 1 1225
2 76767 1 1225
2 76768 1 1237
2 76769 1 1237
2 76770 1 1237
2 76771 1 1237
2 76772 1 1237
2 76773 1 1237
2 76774 1 1237
2 76775 1 1237
2 76776 1 1237
2 76777 1 1237
2 76778 1 1237
2 76779 1 1237
2 76780 1 1237
2 76781 1 1237
2 76782 1 1237
2 76783 1 1237
2 76784 1 1237
2 76785 1 1237
2 76786 1 1237
2 76787 1 1237
2 76788 1 1237
2 76789 1 1237
2 76790 1 1238
2 76791 1 1238
2 76792 1 1238
2 76793 1 1238
2 76794 1 1238
2 76795 1 1241
2 76796 1 1241
2 76797 1 1241
2 76798 1 1241
2 76799 1 1241
2 76800 1 1241
2 76801 1 1241
2 76802 1 1241
2 76803 1 1241
2 76804 1 1241
2 76805 1 1241
2 76806 1 1241
2 76807 1 1241
2 76808 1 1245
2 76809 1 1245
2 76810 1 1245
2 76811 1 1245
2 76812 1 1245
2 76813 1 1245
2 76814 1 1245
2 76815 1 1245
2 76816 1 1245
2 76817 1 1245
2 76818 1 1245
2 76819 1 1245
2 76820 1 1245
2 76821 1 1245
2 76822 1 1245
2 76823 1 1245
2 76824 1 1245
2 76825 1 1245
2 76826 1 1245
2 76827 1 1245
2 76828 1 1245
2 76829 1 1245
2 76830 1 1247
2 76831 1 1247
2 76832 1 1247
2 76833 1 1247
2 76834 1 1248
2 76835 1 1248
2 76836 1 1253
2 76837 1 1253
2 76838 1 1253
2 76839 1 1253
2 76840 1 1253
2 76841 1 1253
2 76842 1 1253
2 76843 1 1253
2 76844 1 1253
2 76845 1 1253
2 76846 1 1253
2 76847 1 1253
2 76848 1 1253
2 76849 1 1253
2 76850 1 1253
2 76851 1 1253
2 76852 1 1253
2 76853 1 1253
2 76854 1 1253
2 76855 1 1261
2 76856 1 1261
2 76857 1 1262
2 76858 1 1262
2 76859 1 1262
2 76860 1 1262
2 76861 1 1262
2 76862 1 1263
2 76863 1 1263
2 76864 1 1263
2 76865 1 1263
2 76866 1 1263
2 76867 1 1263
2 76868 1 1263
2 76869 1 1263
2 76870 1 1264
2 76871 1 1264
2 76872 1 1272
2 76873 1 1272
2 76874 1 1272
2 76875 1 1272
2 76876 1 1272
2 76877 1 1272
2 76878 1 1272
2 76879 1 1272
2 76880 1 1272
2 76881 1 1272
2 76882 1 1272
2 76883 1 1272
2 76884 1 1272
2 76885 1 1272
2 76886 1 1272
2 76887 1 1272
2 76888 1 1272
2 76889 1 1272
2 76890 1 1272
2 76891 1 1272
2 76892 1 1272
2 76893 1 1272
2 76894 1 1272
2 76895 1 1272
2 76896 1 1272
2 76897 1 1272
2 76898 1 1272
2 76899 1 1272
2 76900 1 1272
2 76901 1 1272
2 76902 1 1272
2 76903 1 1272
2 76904 1 1272
2 76905 1 1272
2 76906 1 1272
2 76907 1 1272
2 76908 1 1272
2 76909 1 1272
2 76910 1 1272
2 76911 1 1272
2 76912 1 1272
2 76913 1 1274
2 76914 1 1274
2 76915 1 1274
2 76916 1 1274
2 76917 1 1274
2 76918 1 1274
2 76919 1 1274
2 76920 1 1275
2 76921 1 1275
2 76922 1 1275
2 76923 1 1275
2 76924 1 1275
2 76925 1 1276
2 76926 1 1276
2 76927 1 1276
2 76928 1 1276
2 76929 1 1276
2 76930 1 1276
2 76931 1 1276
2 76932 1 1276
2 76933 1 1276
2 76934 1 1276
2 76935 1 1276
2 76936 1 1276
2 76937 1 1276
2 76938 1 1276
2 76939 1 1276
2 76940 1 1276
2 76941 1 1276
2 76942 1 1276
2 76943 1 1276
2 76944 1 1276
2 76945 1 1276
2 76946 1 1276
2 76947 1 1276
2 76948 1 1276
2 76949 1 1276
2 76950 1 1276
2 76951 1 1276
2 76952 1 1276
2 76953 1 1276
2 76954 1 1276
2 76955 1 1276
2 76956 1 1276
2 76957 1 1276
2 76958 1 1277
2 76959 1 1277
2 76960 1 1277
2 76961 1 1277
2 76962 1 1277
2 76963 1 1278
2 76964 1 1278
2 76965 1 1278
2 76966 1 1278
2 76967 1 1278
2 76968 1 1279
2 76969 1 1279
2 76970 1 1279
2 76971 1 1281
2 76972 1 1281
2 76973 1 1281
2 76974 1 1281
2 76975 1 1281
2 76976 1 1281
2 76977 1 1281
2 76978 1 1281
2 76979 1 1283
2 76980 1 1283
2 76981 1 1283
2 76982 1 1286
2 76983 1 1286
2 76984 1 1287
2 76985 1 1287
2 76986 1 1287
2 76987 1 1287
2 76988 1 1288
2 76989 1 1288
2 76990 1 1288
2 76991 1 1288
2 76992 1 1288
2 76993 1 1288
2 76994 1 1288
2 76995 1 1288
2 76996 1 1288
2 76997 1 1288
2 76998 1 1288
2 76999 1 1288
2 77000 1 1288
2 77001 1 1288
2 77002 1 1289
2 77003 1 1289
2 77004 1 1289
2 77005 1 1298
2 77006 1 1298
2 77007 1 1298
2 77008 1 1301
2 77009 1 1301
2 77010 1 1301
2 77011 1 1301
2 77012 1 1301
2 77013 1 1301
2 77014 1 1301
2 77015 1 1301
2 77016 1 1301
2 77017 1 1301
2 77018 1 1301
2 77019 1 1302
2 77020 1 1302
2 77021 1 1302
2 77022 1 1302
2 77023 1 1302
2 77024 1 1302
2 77025 1 1302
2 77026 1 1302
2 77027 1 1302
2 77028 1 1302
2 77029 1 1302
2 77030 1 1302
2 77031 1 1306
2 77032 1 1306
2 77033 1 1306
2 77034 1 1306
2 77035 1 1306
2 77036 1 1306
2 77037 1 1306
2 77038 1 1306
2 77039 1 1306
2 77040 1 1306
2 77041 1 1306
2 77042 1 1306
2 77043 1 1306
2 77044 1 1306
2 77045 1 1306
2 77046 1 1307
2 77047 1 1307
2 77048 1 1307
2 77049 1 1307
2 77050 1 1307
2 77051 1 1308
2 77052 1 1308
2 77053 1 1309
2 77054 1 1309
2 77055 1 1311
2 77056 1 1311
2 77057 1 1314
2 77058 1 1314
2 77059 1 1314
2 77060 1 1314
2 77061 1 1314
2 77062 1 1314
2 77063 1 1314
2 77064 1 1314
2 77065 1 1315
2 77066 1 1315
2 77067 1 1315
2 77068 1 1315
2 77069 1 1315
2 77070 1 1315
2 77071 1 1315
2 77072 1 1316
2 77073 1 1316
2 77074 1 1317
2 77075 1 1317
2 77076 1 1318
2 77077 1 1318
2 77078 1 1325
2 77079 1 1325
2 77080 1 1325
2 77081 1 1325
2 77082 1 1325
2 77083 1 1325
2 77084 1 1325
2 77085 1 1325
2 77086 1 1325
2 77087 1 1325
2 77088 1 1325
2 77089 1 1325
2 77090 1 1325
2 77091 1 1325
2 77092 1 1325
2 77093 1 1325
2 77094 1 1325
2 77095 1 1325
2 77096 1 1325
2 77097 1 1325
2 77098 1 1325
2 77099 1 1325
2 77100 1 1325
2 77101 1 1325
2 77102 1 1325
2 77103 1 1326
2 77104 1 1326
2 77105 1 1326
2 77106 1 1326
2 77107 1 1327
2 77108 1 1327
2 77109 1 1329
2 77110 1 1329
2 77111 1 1329
2 77112 1 1329
2 77113 1 1329
2 77114 1 1329
2 77115 1 1329
2 77116 1 1330
2 77117 1 1330
2 77118 1 1330
2 77119 1 1330
2 77120 1 1330
2 77121 1 1330
2 77122 1 1330
2 77123 1 1340
2 77124 1 1340
2 77125 1 1340
2 77126 1 1340
2 77127 1 1340
2 77128 1 1340
2 77129 1 1340
2 77130 1 1340
2 77131 1 1340
2 77132 1 1340
2 77133 1 1340
2 77134 1 1341
2 77135 1 1341
2 77136 1 1341
2 77137 1 1341
2 77138 1 1341
2 77139 1 1343
2 77140 1 1343
2 77141 1 1344
2 77142 1 1344
2 77143 1 1344
2 77144 1 1344
2 77145 1 1344
2 77146 1 1344
2 77147 1 1344
2 77148 1 1344
2 77149 1 1344
2 77150 1 1344
2 77151 1 1344
2 77152 1 1344
2 77153 1 1344
2 77154 1 1344
2 77155 1 1344
2 77156 1 1344
2 77157 1 1344
2 77158 1 1344
2 77159 1 1345
2 77160 1 1345
2 77161 1 1345
2 77162 1 1345
2 77163 1 1346
2 77164 1 1346
2 77165 1 1346
2 77166 1 1346
2 77167 1 1346
2 77168 1 1346
2 77169 1 1346
2 77170 1 1346
2 77171 1 1346
2 77172 1 1346
2 77173 1 1346
2 77174 1 1346
2 77175 1 1346
2 77176 1 1347
2 77177 1 1347
2 77178 1 1355
2 77179 1 1355
2 77180 1 1355
2 77181 1 1355
2 77182 1 1355
2 77183 1 1355
2 77184 1 1355
2 77185 1 1355
2 77186 1 1355
2 77187 1 1355
2 77188 1 1355
2 77189 1 1355
2 77190 1 1355
2 77191 1 1355
2 77192 1 1355
2 77193 1 1355
2 77194 1 1355
2 77195 1 1355
2 77196 1 1355
2 77197 1 1355
2 77198 1 1355
2 77199 1 1355
2 77200 1 1355
2 77201 1 1355
2 77202 1 1355
2 77203 1 1355
2 77204 1 1355
2 77205 1 1355
2 77206 1 1355
2 77207 1 1355
2 77208 1 1355
2 77209 1 1355
2 77210 1 1356
2 77211 1 1356
2 77212 1 1356
2 77213 1 1357
2 77214 1 1357
2 77215 1 1366
2 77216 1 1366
2 77217 1 1366
2 77218 1 1366
2 77219 1 1366
2 77220 1 1366
2 77221 1 1366
2 77222 1 1366
2 77223 1 1366
2 77224 1 1366
2 77225 1 1366
2 77226 1 1366
2 77227 1 1366
2 77228 1 1366
2 77229 1 1366
2 77230 1 1366
2 77231 1 1366
2 77232 1 1366
2 77233 1 1366
2 77234 1 1366
2 77235 1 1366
2 77236 1 1366
2 77237 1 1366
2 77238 1 1366
2 77239 1 1366
2 77240 1 1366
2 77241 1 1366
2 77242 1 1366
2 77243 1 1366
2 77244 1 1366
2 77245 1 1366
2 77246 1 1366
2 77247 1 1366
2 77248 1 1366
2 77249 1 1366
2 77250 1 1366
2 77251 1 1366
2 77252 1 1366
2 77253 1 1366
2 77254 1 1366
2 77255 1 1366
2 77256 1 1366
2 77257 1 1366
2 77258 1 1366
2 77259 1 1366
2 77260 1 1366
2 77261 1 1366
2 77262 1 1366
2 77263 1 1366
2 77264 1 1366
2 77265 1 1366
2 77266 1 1366
2 77267 1 1366
2 77268 1 1367
2 77269 1 1367
2 77270 1 1367
2 77271 1 1367
2 77272 1 1367
2 77273 1 1368
2 77274 1 1368
2 77275 1 1368
2 77276 1 1368
2 77277 1 1368
2 77278 1 1369
2 77279 1 1369
2 77280 1 1369
2 77281 1 1370
2 77282 1 1370
2 77283 1 1370
2 77284 1 1371
2 77285 1 1371
2 77286 1 1371
2 77287 1 1373
2 77288 1 1373
2 77289 1 1380
2 77290 1 1380
2 77291 1 1380
2 77292 1 1380
2 77293 1 1380
2 77294 1 1380
2 77295 1 1380
2 77296 1 1380
2 77297 1 1380
2 77298 1 1380
2 77299 1 1380
2 77300 1 1380
2 77301 1 1380
2 77302 1 1380
2 77303 1 1380
2 77304 1 1380
2 77305 1 1380
2 77306 1 1380
2 77307 1 1380
2 77308 1 1380
2 77309 1 1381
2 77310 1 1381
2 77311 1 1381
2 77312 1 1382
2 77313 1 1382
2 77314 1 1382
2 77315 1 1382
2 77316 1 1382
2 77317 1 1382
2 77318 1 1382
2 77319 1 1382
2 77320 1 1382
2 77321 1 1382
2 77322 1 1382
2 77323 1 1382
2 77324 1 1389
2 77325 1 1389
2 77326 1 1389
2 77327 1 1389
2 77328 1 1389
2 77329 1 1389
2 77330 1 1389
2 77331 1 1389
2 77332 1 1389
2 77333 1 1389
2 77334 1 1389
2 77335 1 1389
2 77336 1 1389
2 77337 1 1389
2 77338 1 1389
2 77339 1 1390
2 77340 1 1390
2 77341 1 1390
2 77342 1 1391
2 77343 1 1391
2 77344 1 1391
2 77345 1 1391
2 77346 1 1391
2 77347 1 1391
2 77348 1 1391
2 77349 1 1391
2 77350 1 1391
2 77351 1 1391
2 77352 1 1392
2 77353 1 1392
2 77354 1 1392
2 77355 1 1392
2 77356 1 1392
2 77357 1 1392
2 77358 1 1392
2 77359 1 1392
2 77360 1 1392
2 77361 1 1392
2 77362 1 1393
2 77363 1 1393
2 77364 1 1393
2 77365 1 1398
2 77366 1 1398
2 77367 1 1406
2 77368 1 1406
2 77369 1 1417
2 77370 1 1417
2 77371 1 1417
2 77372 1 1417
2 77373 1 1417
2 77374 1 1417
2 77375 1 1417
2 77376 1 1417
2 77377 1 1417
2 77378 1 1417
2 77379 1 1417
2 77380 1 1417
2 77381 1 1417
2 77382 1 1417
2 77383 1 1417
2 77384 1 1417
2 77385 1 1417
2 77386 1 1426
2 77387 1 1426
2 77388 1 1426
2 77389 1 1426
2 77390 1 1426
2 77391 1 1426
2 77392 1 1426
2 77393 1 1426
2 77394 1 1426
2 77395 1 1426
2 77396 1 1426
2 77397 1 1426
2 77398 1 1426
2 77399 1 1426
2 77400 1 1426
2 77401 1 1429
2 77402 1 1429
2 77403 1 1429
2 77404 1 1429
2 77405 1 1429
2 77406 1 1429
2 77407 1 1429
2 77408 1 1429
2 77409 1 1429
2 77410 1 1429
2 77411 1 1429
2 77412 1 1429
2 77413 1 1429
2 77414 1 1429
2 77415 1 1430
2 77416 1 1430
2 77417 1 1430
2 77418 1 1430
2 77419 1 1430
2 77420 1 1432
2 77421 1 1432
2 77422 1 1432
2 77423 1 1432
2 77424 1 1433
2 77425 1 1433
2 77426 1 1441
2 77427 1 1441
2 77428 1 1441
2 77429 1 1441
2 77430 1 1441
2 77431 1 1441
2 77432 1 1441
2 77433 1 1441
2 77434 1 1441
2 77435 1 1441
2 77436 1 1441
2 77437 1 1441
2 77438 1 1441
2 77439 1 1441
2 77440 1 1441
2 77441 1 1441
2 77442 1 1441
2 77443 1 1441
2 77444 1 1441
2 77445 1 1441
2 77446 1 1442
2 77447 1 1442
2 77448 1 1443
2 77449 1 1443
2 77450 1 1443
2 77451 1 1443
2 77452 1 1443
2 77453 1 1443
2 77454 1 1444
2 77455 1 1444
2 77456 1 1444
2 77457 1 1444
2 77458 1 1444
2 77459 1 1444
2 77460 1 1455
2 77461 1 1455
2 77462 1 1455
2 77463 1 1455
2 77464 1 1455
2 77465 1 1455
2 77466 1 1455
2 77467 1 1455
2 77468 1 1455
2 77469 1 1455
2 77470 1 1455
2 77471 1 1455
2 77472 1 1455
2 77473 1 1455
2 77474 1 1455
2 77475 1 1455
2 77476 1 1455
2 77477 1 1455
2 77478 1 1455
2 77479 1 1457
2 77480 1 1457
2 77481 1 1461
2 77482 1 1461
2 77483 1 1461
2 77484 1 1461
2 77485 1 1461
2 77486 1 1468
2 77487 1 1468
2 77488 1 1468
2 77489 1 1468
2 77490 1 1468
2 77491 1 1468
2 77492 1 1468
2 77493 1 1468
2 77494 1 1468
2 77495 1 1468
2 77496 1 1468
2 77497 1 1468
2 77498 1 1468
2 77499 1 1468
2 77500 1 1468
2 77501 1 1468
2 77502 1 1468
2 77503 1 1469
2 77504 1 1469
2 77505 1 1469
2 77506 1 1470
2 77507 1 1470
2 77508 1 1470
2 77509 1 1470
2 77510 1 1470
2 77511 1 1473
2 77512 1 1473
2 77513 1 1473
2 77514 1 1473
2 77515 1 1473
2 77516 1 1473
2 77517 1 1474
2 77518 1 1474
2 77519 1 1474
2 77520 1 1474
2 77521 1 1474
2 77522 1 1474
2 77523 1 1474
2 77524 1 1474
2 77525 1 1474
2 77526 1 1474
2 77527 1 1474
2 77528 1 1474
2 77529 1 1474
2 77530 1 1474
2 77531 1 1475
2 77532 1 1475
2 77533 1 1475
2 77534 1 1476
2 77535 1 1476
2 77536 1 1476
2 77537 1 1476
2 77538 1 1477
2 77539 1 1477
2 77540 1 1477
2 77541 1 1484
2 77542 1 1484
2 77543 1 1484
2 77544 1 1484
2 77545 1 1484
2 77546 1 1484
2 77547 1 1484
2 77548 1 1484
2 77549 1 1484
2 77550 1 1484
2 77551 1 1485
2 77552 1 1485
2 77553 1 1485
2 77554 1 1485
2 77555 1 1485
2 77556 1 1485
2 77557 1 1485
2 77558 1 1485
2 77559 1 1485
2 77560 1 1485
2 77561 1 1485
2 77562 1 1496
2 77563 1 1496
2 77564 1 1496
2 77565 1 1499
2 77566 1 1499
2 77567 1 1499
2 77568 1 1499
2 77569 1 1499
2 77570 1 1499
2 77571 1 1499
2 77572 1 1499
2 77573 1 1499
2 77574 1 1499
2 77575 1 1499
2 77576 1 1499
2 77577 1 1499
2 77578 1 1499
2 77579 1 1499
2 77580 1 1499
2 77581 1 1499
2 77582 1 1500
2 77583 1 1500
2 77584 1 1500
2 77585 1 1500
2 77586 1 1501
2 77587 1 1501
2 77588 1 1520
2 77589 1 1520
2 77590 1 1520
2 77591 1 1521
2 77592 1 1521
2 77593 1 1521
2 77594 1 1521
2 77595 1 1521
2 77596 1 1521
2 77597 1 1521
2 77598 1 1521
2 77599 1 1521
2 77600 1 1521
2 77601 1 1521
2 77602 1 1521
2 77603 1 1521
2 77604 1 1521
2 77605 1 1521
2 77606 1 1523
2 77607 1 1523
2 77608 1 1523
2 77609 1 1523
2 77610 1 1523
2 77611 1 1523
2 77612 1 1523
2 77613 1 1523
2 77614 1 1523
2 77615 1 1523
2 77616 1 1523
2 77617 1 1523
2 77618 1 1524
2 77619 1 1524
2 77620 1 1525
2 77621 1 1525
2 77622 1 1525
2 77623 1 1525
2 77624 1 1525
2 77625 1 1525
2 77626 1 1529
2 77627 1 1529
2 77628 1 1529
2 77629 1 1529
2 77630 1 1529
2 77631 1 1529
2 77632 1 1529
2 77633 1 1530
2 77634 1 1530
2 77635 1 1530
2 77636 1 1532
2 77637 1 1532
2 77638 1 1533
2 77639 1 1533
2 77640 1 1533
2 77641 1 1533
2 77642 1 1533
2 77643 1 1533
2 77644 1 1533
2 77645 1 1533
2 77646 1 1534
2 77647 1 1534
2 77648 1 1538
2 77649 1 1538
2 77650 1 1538
2 77651 1 1558
2 77652 1 1558
2 77653 1 1558
2 77654 1 1558
2 77655 1 1558
2 77656 1 1558
2 77657 1 1558
2 77658 1 1558
2 77659 1 1558
2 77660 1 1558
2 77661 1 1558
2 77662 1 1558
2 77663 1 1558
2 77664 1 1558
2 77665 1 1558
2 77666 1 1558
2 77667 1 1558
2 77668 1 1558
2 77669 1 1558
2 77670 1 1558
2 77671 1 1558
2 77672 1 1558
2 77673 1 1558
2 77674 1 1559
2 77675 1 1559
2 77676 1 1559
2 77677 1 1559
2 77678 1 1559
2 77679 1 1560
2 77680 1 1560
2 77681 1 1560
2 77682 1 1560
2 77683 1 1560
2 77684 1 1560
2 77685 1 1560
2 77686 1 1560
2 77687 1 1560
2 77688 1 1561
2 77689 1 1561
2 77690 1 1561
2 77691 1 1561
2 77692 1 1561
2 77693 1 1561
2 77694 1 1562
2 77695 1 1562
2 77696 1 1564
2 77697 1 1564
2 77698 1 1564
2 77699 1 1564
2 77700 1 1566
2 77701 1 1566
2 77702 1 1567
2 77703 1 1567
2 77704 1 1567
2 77705 1 1567
2 77706 1 1567
2 77707 1 1567
2 77708 1 1567
2 77709 1 1567
2 77710 1 1569
2 77711 1 1569
2 77712 1 1570
2 77713 1 1570
2 77714 1 1570
2 77715 1 1570
2 77716 1 1570
2 77717 1 1570
2 77718 1 1570
2 77719 1 1570
2 77720 1 1570
2 77721 1 1571
2 77722 1 1571
2 77723 1 1572
2 77724 1 1572
2 77725 1 1572
2 77726 1 1572
2 77727 1 1572
2 77728 1 1572
2 77729 1 1573
2 77730 1 1573
2 77731 1 1573
2 77732 1 1573
2 77733 1 1573
2 77734 1 1573
2 77735 1 1573
2 77736 1 1573
2 77737 1 1573
2 77738 1 1574
2 77739 1 1574
2 77740 1 1585
2 77741 1 1585
2 77742 1 1585
2 77743 1 1585
2 77744 1 1585
2 77745 1 1585
2 77746 1 1586
2 77747 1 1586
2 77748 1 1586
2 77749 1 1586
2 77750 1 1586
2 77751 1 1586
2 77752 1 1586
2 77753 1 1586
2 77754 1 1586
2 77755 1 1586
2 77756 1 1586
2 77757 1 1588
2 77758 1 1588
2 77759 1 1595
2 77760 1 1595
2 77761 1 1595
2 77762 1 1595
2 77763 1 1595
2 77764 1 1595
2 77765 1 1595
2 77766 1 1595
2 77767 1 1595
2 77768 1 1595
2 77769 1 1596
2 77770 1 1596
2 77771 1 1597
2 77772 1 1597
2 77773 1 1598
2 77774 1 1598
2 77775 1 1598
2 77776 1 1599
2 77777 1 1599
2 77778 1 1600
2 77779 1 1600
2 77780 1 1607
2 77781 1 1607
2 77782 1 1607
2 77783 1 1608
2 77784 1 1608
2 77785 1 1611
2 77786 1 1611
2 77787 1 1611
2 77788 1 1611
2 77789 1 1611
2 77790 1 1622
2 77791 1 1622
2 77792 1 1622
2 77793 1 1622
2 77794 1 1622
2 77795 1 1622
2 77796 1 1622
2 77797 1 1622
2 77798 1 1622
2 77799 1 1622
2 77800 1 1622
2 77801 1 1622
2 77802 1 1622
2 77803 1 1623
2 77804 1 1623
2 77805 1 1626
2 77806 1 1626
2 77807 1 1626
2 77808 1 1626
2 77809 1 1626
2 77810 1 1626
2 77811 1 1626
2 77812 1 1626
2 77813 1 1626
2 77814 1 1626
2 77815 1 1626
2 77816 1 1626
2 77817 1 1626
2 77818 1 1626
2 77819 1 1626
2 77820 1 1626
2 77821 1 1626
2 77822 1 1626
2 77823 1 1626
2 77824 1 1626
2 77825 1 1626
2 77826 1 1626
2 77827 1 1627
2 77828 1 1627
2 77829 1 1628
2 77830 1 1628
2 77831 1 1628
2 77832 1 1628
2 77833 1 1628
2 77834 1 1628
2 77835 1 1628
2 77836 1 1629
2 77837 1 1629
2 77838 1 1629
2 77839 1 1629
2 77840 1 1629
2 77841 1 1629
2 77842 1 1629
2 77843 1 1629
2 77844 1 1629
2 77845 1 1631
2 77846 1 1631
2 77847 1 1634
2 77848 1 1634
2 77849 1 1634
2 77850 1 1634
2 77851 1 1634
2 77852 1 1634
2 77853 1 1634
2 77854 1 1634
2 77855 1 1634
2 77856 1 1636
2 77857 1 1636
2 77858 1 1636
2 77859 1 1636
2 77860 1 1636
2 77861 1 1636
2 77862 1 1637
2 77863 1 1637
2 77864 1 1644
2 77865 1 1644
2 77866 1 1647
2 77867 1 1647
2 77868 1 1647
2 77869 1 1647
2 77870 1 1647
2 77871 1 1647
2 77872 1 1647
2 77873 1 1647
2 77874 1 1647
2 77875 1 1657
2 77876 1 1657
2 77877 1 1657
2 77878 1 1657
2 77879 1 1657
2 77880 1 1657
2 77881 1 1658
2 77882 1 1658
2 77883 1 1658
2 77884 1 1658
2 77885 1 1659
2 77886 1 1659
2 77887 1 1660
2 77888 1 1660
2 77889 1 1669
2 77890 1 1669
2 77891 1 1669
2 77892 1 1676
2 77893 1 1676
2 77894 1 1677
2 77895 1 1677
2 77896 1 1677
2 77897 1 1677
2 77898 1 1677
2 77899 1 1677
2 77900 1 1677
2 77901 1 1677
2 77902 1 1677
2 77903 1 1677
2 77904 1 1677
2 77905 1 1677
2 77906 1 1678
2 77907 1 1678
2 77908 1 1678
2 77909 1 1679
2 77910 1 1679
2 77911 1 1679
2 77912 1 1679
2 77913 1 1692
2 77914 1 1692
2 77915 1 1692
2 77916 1 1693
2 77917 1 1693
2 77918 1 1693
2 77919 1 1693
2 77920 1 1693
2 77921 1 1693
2 77922 1 1693
2 77923 1 1693
2 77924 1 1693
2 77925 1 1693
2 77926 1 1693
2 77927 1 1705
2 77928 1 1705
2 77929 1 1705
2 77930 1 1705
2 77931 1 1705
2 77932 1 1705
2 77933 1 1705
2 77934 1 1705
2 77935 1 1705
2 77936 1 1705
2 77937 1 1706
2 77938 1 1706
2 77939 1 1706
2 77940 1 1706
2 77941 1 1706
2 77942 1 1706
2 77943 1 1706
2 77944 1 1706
2 77945 1 1706
2 77946 1 1706
2 77947 1 1706
2 77948 1 1706
2 77949 1 1706
2 77950 1 1706
2 77951 1 1706
2 77952 1 1706
2 77953 1 1706
2 77954 1 1706
2 77955 1 1706
2 77956 1 1707
2 77957 1 1707
2 77958 1 1708
2 77959 1 1708
2 77960 1 1708
2 77961 1 1714
2 77962 1 1714
2 77963 1 1714
2 77964 1 1714
2 77965 1 1714
2 77966 1 1714
2 77967 1 1714
2 77968 1 1714
2 77969 1 1714
2 77970 1 1714
2 77971 1 1714
2 77972 1 1715
2 77973 1 1715
2 77974 1 1715
2 77975 1 1716
2 77976 1 1716
2 77977 1 1720
2 77978 1 1720
2 77979 1 1720
2 77980 1 1720
2 77981 1 1720
2 77982 1 1720
2 77983 1 1720
2 77984 1 1721
2 77985 1 1721
2 77986 1 1723
2 77987 1 1723
2 77988 1 1723
2 77989 1 1723
2 77990 1 1723
2 77991 1 1723
2 77992 1 1723
2 77993 1 1723
2 77994 1 1724
2 77995 1 1724
2 77996 1 1724
2 77997 1 1724
2 77998 1 1724
2 77999 1 1724
2 78000 1 1724
2 78001 1 1724
2 78002 1 1724
2 78003 1 1724
2 78004 1 1724
2 78005 1 1724
2 78006 1 1724
2 78007 1 1724
2 78008 1 1724
2 78009 1 1724
2 78010 1 1724
2 78011 1 1724
2 78012 1 1725
2 78013 1 1725
2 78014 1 1725
2 78015 1 1739
2 78016 1 1739
2 78017 1 1739
2 78018 1 1739
2 78019 1 1739
2 78020 1 1752
2 78021 1 1752
2 78022 1 1752
2 78023 1 1752
2 78024 1 1752
2 78025 1 1752
2 78026 1 1752
2 78027 1 1752
2 78028 1 1752
2 78029 1 1752
2 78030 1 1752
2 78031 1 1752
2 78032 1 1754
2 78033 1 1754
2 78034 1 1754
2 78035 1 1754
2 78036 1 1754
2 78037 1 1754
2 78038 1 1754
2 78039 1 1754
2 78040 1 1754
2 78041 1 1754
2 78042 1 1754
2 78043 1 1754
2 78044 1 1754
2 78045 1 1754
2 78046 1 1754
2 78047 1 1755
2 78048 1 1755
2 78049 1 1758
2 78050 1 1758
2 78051 1 1758
2 78052 1 1758
2 78053 1 1758
2 78054 1 1758
2 78055 1 1758
2 78056 1 1758
2 78057 1 1758
2 78058 1 1758
2 78059 1 1758
2 78060 1 1758
2 78061 1 1758
2 78062 1 1758
2 78063 1 1758
2 78064 1 1758
2 78065 1 1758
2 78066 1 1758
2 78067 1 1758
2 78068 1 1758
2 78069 1 1758
2 78070 1 1758
2 78071 1 1758
2 78072 1 1758
2 78073 1 1758
2 78074 1 1758
2 78075 1 1758
2 78076 1 1758
2 78077 1 1758
2 78078 1 1758
2 78079 1 1758
2 78080 1 1758
2 78081 1 1758
2 78082 1 1758
2 78083 1 1758
2 78084 1 1758
2 78085 1 1758
2 78086 1 1758
2 78087 1 1758
2 78088 1 1759
2 78089 1 1759
2 78090 1 1759
2 78091 1 1759
2 78092 1 1760
2 78093 1 1760
2 78094 1 1760
2 78095 1 1760
2 78096 1 1760
2 78097 1 1768
2 78098 1 1768
2 78099 1 1768
2 78100 1 1768
2 78101 1 1768
2 78102 1 1768
2 78103 1 1768
2 78104 1 1768
2 78105 1 1768
2 78106 1 1768
2 78107 1 1768
2 78108 1 1768
2 78109 1 1768
2 78110 1 1768
2 78111 1 1768
2 78112 1 1768
2 78113 1 1768
2 78114 1 1768
2 78115 1 1768
2 78116 1 1768
2 78117 1 1768
2 78118 1 1768
2 78119 1 1769
2 78120 1 1769
2 78121 1 1769
2 78122 1 1769
2 78123 1 1769
2 78124 1 1769
2 78125 1 1769
2 78126 1 1770
2 78127 1 1770
2 78128 1 1770
2 78129 1 1770
2 78130 1 1770
2 78131 1 1770
2 78132 1 1770
2 78133 1 1770
2 78134 1 1771
2 78135 1 1771
2 78136 1 1771
2 78137 1 1776
2 78138 1 1776
2 78139 1 1776
2 78140 1 1783
2 78141 1 1783
2 78142 1 1783
2 78143 1 1783
2 78144 1 1783
2 78145 1 1783
2 78146 1 1783
2 78147 1 1783
2 78148 1 1783
2 78149 1 1783
2 78150 1 1783
2 78151 1 1783
2 78152 1 1783
2 78153 1 1783
2 78154 1 1784
2 78155 1 1784
2 78156 1 1785
2 78157 1 1785
2 78158 1 1785
2 78159 1 1786
2 78160 1 1786
2 78161 1 1794
2 78162 1 1794
2 78163 1 1796
2 78164 1 1796
2 78165 1 1796
2 78166 1 1796
2 78167 1 1797
2 78168 1 1797
2 78169 1 1798
2 78170 1 1798
2 78171 1 1799
2 78172 1 1799
2 78173 1 1799
2 78174 1 1799
2 78175 1 1809
2 78176 1 1809
2 78177 1 1809
2 78178 1 1809
2 78179 1 1809
2 78180 1 1809
2 78181 1 1809
2 78182 1 1810
2 78183 1 1810
2 78184 1 1810
2 78185 1 1810
2 78186 1 1810
2 78187 1 1810
2 78188 1 1810
2 78189 1 1810
2 78190 1 1810
2 78191 1 1810
2 78192 1 1810
2 78193 1 1810
2 78194 1 1810
2 78195 1 1810
2 78196 1 1810
2 78197 1 1810
2 78198 1 1810
2 78199 1 1810
2 78200 1 1810
2 78201 1 1810
2 78202 1 1810
2 78203 1 1810
2 78204 1 1810
2 78205 1 1811
2 78206 1 1811
2 78207 1 1811
2 78208 1 1811
2 78209 1 1811
2 78210 1 1811
2 78211 1 1811
2 78212 1 1811
2 78213 1 1811
2 78214 1 1811
2 78215 1 1811
2 78216 1 1811
2 78217 1 1811
2 78218 1 1811
2 78219 1 1811
2 78220 1 1812
2 78221 1 1812
2 78222 1 1812
2 78223 1 1812
2 78224 1 1812
2 78225 1 1812
2 78226 1 1812
2 78227 1 1813
2 78228 1 1813
2 78229 1 1817
2 78230 1 1817
2 78231 1 1817
2 78232 1 1817
2 78233 1 1817
2 78234 1 1817
2 78235 1 1817
2 78236 1 1817
2 78237 1 1817
2 78238 1 1817
2 78239 1 1817
2 78240 1 1817
2 78241 1 1817
2 78242 1 1817
2 78243 1 1817
2 78244 1 1819
2 78245 1 1819
2 78246 1 1819
2 78247 1 1819
2 78248 1 1819
2 78249 1 1820
2 78250 1 1820
2 78251 1 1820
2 78252 1 1820
2 78253 1 1823
2 78254 1 1823
2 78255 1 1832
2 78256 1 1832
2 78257 1 1832
2 78258 1 1832
2 78259 1 1832
2 78260 1 1832
2 78261 1 1832
2 78262 1 1832
2 78263 1 1832
2 78264 1 1832
2 78265 1 1832
2 78266 1 1832
2 78267 1 1832
2 78268 1 1832
2 78269 1 1832
2 78270 1 1832
2 78271 1 1832
2 78272 1 1832
2 78273 1 1832
2 78274 1 1832
2 78275 1 1834
2 78276 1 1834
2 78277 1 1834
2 78278 1 1834
2 78279 1 1834
2 78280 1 1834
2 78281 1 1834
2 78282 1 1834
2 78283 1 1834
2 78284 1 1834
2 78285 1 1834
2 78286 1 1834
2 78287 1 1834
2 78288 1 1834
2 78289 1 1841
2 78290 1 1841
2 78291 1 1841
2 78292 1 1841
2 78293 1 1842
2 78294 1 1842
2 78295 1 1842
2 78296 1 1844
2 78297 1 1844
2 78298 1 1844
2 78299 1 1844
2 78300 1 1844
2 78301 1 1844
2 78302 1 1845
2 78303 1 1845
2 78304 1 1852
2 78305 1 1852
2 78306 1 1852
2 78307 1 1852
2 78308 1 1852
2 78309 1 1852
2 78310 1 1852
2 78311 1 1852
2 78312 1 1852
2 78313 1 1852
2 78314 1 1852
2 78315 1 1852
2 78316 1 1852
2 78317 1 1852
2 78318 1 1852
2 78319 1 1853
2 78320 1 1853
2 78321 1 1853
2 78322 1 1853
2 78323 1 1853
2 78324 1 1853
2 78325 1 1853
2 78326 1 1853
2 78327 1 1853
2 78328 1 1853
2 78329 1 1853
2 78330 1 1853
2 78331 1 1853
2 78332 1 1853
2 78333 1 1853
2 78334 1 1853
2 78335 1 1853
2 78336 1 1853
2 78337 1 1853
2 78338 1 1853
2 78339 1 1853
2 78340 1 1853
2 78341 1 1853
2 78342 1 1853
2 78343 1 1853
2 78344 1 1853
2 78345 1 1853
2 78346 1 1853
2 78347 1 1853
2 78348 1 1853
2 78349 1 1853
2 78350 1 1853
2 78351 1 1853
2 78352 1 1853
2 78353 1 1853
2 78354 1 1853
2 78355 1 1853
2 78356 1 1853
2 78357 1 1854
2 78358 1 1854
2 78359 1 1854
2 78360 1 1854
2 78361 1 1854
2 78362 1 1855
2 78363 1 1855
2 78364 1 1855
2 78365 1 1857
2 78366 1 1857
2 78367 1 1864
2 78368 1 1864
2 78369 1 1864
2 78370 1 1864
2 78371 1 1876
2 78372 1 1876
2 78373 1 1876
2 78374 1 1876
2 78375 1 1876
2 78376 1 1876
2 78377 1 1876
2 78378 1 1876
2 78379 1 1876
2 78380 1 1876
2 78381 1 1876
2 78382 1 1876
2 78383 1 1877
2 78384 1 1877
2 78385 1 1878
2 78386 1 1878
2 78387 1 1878
2 78388 1 1878
2 78389 1 1878
2 78390 1 1879
2 78391 1 1879
2 78392 1 1882
2 78393 1 1882
2 78394 1 1882
2 78395 1 1882
2 78396 1 1882
2 78397 1 1882
2 78398 1 1882
2 78399 1 1882
2 78400 1 1882
2 78401 1 1882
2 78402 1 1883
2 78403 1 1883
2 78404 1 1899
2 78405 1 1899
2 78406 1 1899
2 78407 1 1899
2 78408 1 1899
2 78409 1 1899
2 78410 1 1899
2 78411 1 1899
2 78412 1 1899
2 78413 1 1899
2 78414 1 1899
2 78415 1 1899
2 78416 1 1899
2 78417 1 1899
2 78418 1 1899
2 78419 1 1899
2 78420 1 1899
2 78421 1 1899
2 78422 1 1901
2 78423 1 1901
2 78424 1 1903
2 78425 1 1903
2 78426 1 1903
2 78427 1 1903
2 78428 1 1903
2 78429 1 1903
2 78430 1 1903
2 78431 1 1903
2 78432 1 1903
2 78433 1 1903
2 78434 1 1903
2 78435 1 1904
2 78436 1 1904
2 78437 1 1904
2 78438 1 1904
2 78439 1 1904
2 78440 1 1904
2 78441 1 1904
2 78442 1 1904
2 78443 1 1904
2 78444 1 1904
2 78445 1 1904
2 78446 1 1904
2 78447 1 1904
2 78448 1 1904
2 78449 1 1904
2 78450 1 1904
2 78451 1 1904
2 78452 1 1904
2 78453 1 1904
2 78454 1 1905
2 78455 1 1905
2 78456 1 1917
2 78457 1 1917
2 78458 1 1917
2 78459 1 1917
2 78460 1 1917
2 78461 1 1917
2 78462 1 1917
2 78463 1 1917
2 78464 1 1917
2 78465 1 1917
2 78466 1 1917
2 78467 1 1917
2 78468 1 1917
2 78469 1 1917
2 78470 1 1917
2 78471 1 1917
2 78472 1 1917
2 78473 1 1917
2 78474 1 1917
2 78475 1 1917
2 78476 1 1917
2 78477 1 1917
2 78478 1 1917
2 78479 1 1917
2 78480 1 1917
2 78481 1 1917
2 78482 1 1917
2 78483 1 1917
2 78484 1 1917
2 78485 1 1917
2 78486 1 1917
2 78487 1 1917
2 78488 1 1918
2 78489 1 1918
2 78490 1 1918
2 78491 1 1918
2 78492 1 1918
2 78493 1 1918
2 78494 1 1918
2 78495 1 1918
2 78496 1 1918
2 78497 1 1918
2 78498 1 1918
2 78499 1 1918
2 78500 1 1918
2 78501 1 1918
2 78502 1 1918
2 78503 1 1918
2 78504 1 1918
2 78505 1 1918
2 78506 1 1918
2 78507 1 1918
2 78508 1 1918
2 78509 1 1918
2 78510 1 1918
2 78511 1 1918
2 78512 1 1918
2 78513 1 1918
2 78514 1 1918
2 78515 1 1918
2 78516 1 1918
2 78517 1 1918
2 78518 1 1918
2 78519 1 1918
2 78520 1 1918
2 78521 1 1918
2 78522 1 1918
2 78523 1 1918
2 78524 1 1919
2 78525 1 1919
2 78526 1 1926
2 78527 1 1926
2 78528 1 1926
2 78529 1 1926
2 78530 1 1926
2 78531 1 1926
2 78532 1 1926
2 78533 1 1926
2 78534 1 1926
2 78535 1 1926
2 78536 1 1926
2 78537 1 1926
2 78538 1 1926
2 78539 1 1926
2 78540 1 1926
2 78541 1 1926
2 78542 1 1926
2 78543 1 1926
2 78544 1 1926
2 78545 1 1926
2 78546 1 1926
2 78547 1 1926
2 78548 1 1926
2 78549 1 1926
2 78550 1 1926
2 78551 1 1926
2 78552 1 1926
2 78553 1 1926
2 78554 1 1926
2 78555 1 1926
2 78556 1 1926
2 78557 1 1926
2 78558 1 1926
2 78559 1 1926
2 78560 1 1926
2 78561 1 1926
2 78562 1 1926
2 78563 1 1926
2 78564 1 1926
2 78565 1 1926
2 78566 1 1926
2 78567 1 1926
2 78568 1 1926
2 78569 1 1926
2 78570 1 1926
2 78571 1 1926
2 78572 1 1926
2 78573 1 1928
2 78574 1 1928
2 78575 1 1928
2 78576 1 1929
2 78577 1 1929
2 78578 1 1929
2 78579 1 1932
2 78580 1 1932
2 78581 1 1932
2 78582 1 1932
2 78583 1 1932
2 78584 1 1932
2 78585 1 1932
2 78586 1 1932
2 78587 1 1932
2 78588 1 1932
2 78589 1 1932
2 78590 1 1932
2 78591 1 1932
2 78592 1 1932
2 78593 1 1932
2 78594 1 1932
2 78595 1 1932
2 78596 1 1932
2 78597 1 1932
2 78598 1 1932
2 78599 1 1932
2 78600 1 1932
2 78601 1 1932
2 78602 1 1932
2 78603 1 1932
2 78604 1 1932
2 78605 1 1932
2 78606 1 1932
2 78607 1 1932
2 78608 1 1932
2 78609 1 1932
2 78610 1 1932
2 78611 1 1932
2 78612 1 1932
2 78613 1 1932
2 78614 1 1932
2 78615 1 1932
2 78616 1 1932
2 78617 1 1932
2 78618 1 1932
2 78619 1 1932
2 78620 1 1932
2 78621 1 1932
2 78622 1 1932
2 78623 1 1932
2 78624 1 1932
2 78625 1 1932
2 78626 1 1934
2 78627 1 1934
2 78628 1 1934
2 78629 1 1934
2 78630 1 1934
2 78631 1 1934
2 78632 1 1935
2 78633 1 1935
2 78634 1 1935
2 78635 1 1942
2 78636 1 1942
2 78637 1 1942
2 78638 1 1943
2 78639 1 1943
2 78640 1 1943
2 78641 1 1950
2 78642 1 1950
2 78643 1 1950
2 78644 1 1950
2 78645 1 1950
2 78646 1 1950
2 78647 1 1950
2 78648 1 1950
2 78649 1 1950
2 78650 1 1950
2 78651 1 1950
2 78652 1 1950
2 78653 1 1950
2 78654 1 1950
2 78655 1 1950
2 78656 1 1950
2 78657 1 1950
2 78658 1 1950
2 78659 1 1950
2 78660 1 1950
2 78661 1 1950
2 78662 1 1950
2 78663 1 1951
2 78664 1 1951
2 78665 1 1952
2 78666 1 1952
2 78667 1 1952
2 78668 1 1953
2 78669 1 1953
2 78670 1 1953
2 78671 1 1953
2 78672 1 1953
2 78673 1 1953
2 78674 1 1953
2 78675 1 1953
2 78676 1 1953
2 78677 1 1953
2 78678 1 1953
2 78679 1 1953
2 78680 1 1953
2 78681 1 1953
2 78682 1 1953
2 78683 1 1953
2 78684 1 1953
2 78685 1 1953
2 78686 1 1954
2 78687 1 1954
2 78688 1 1954
2 78689 1 1954
2 78690 1 1954
2 78691 1 1954
2 78692 1 1954
2 78693 1 1954
2 78694 1 1954
2 78695 1 1954
2 78696 1 1954
2 78697 1 1954
2 78698 1 1954
2 78699 1 1954
2 78700 1 1954
2 78701 1 1954
2 78702 1 1954
2 78703 1 1954
2 78704 1 1962
2 78705 1 1962
2 78706 1 1962
2 78707 1 1963
2 78708 1 1963
2 78709 1 1963
2 78710 1 1963
2 78711 1 1963
2 78712 1 1963
2 78713 1 1963
2 78714 1 1963
2 78715 1 1963
2 78716 1 1963
2 78717 1 1963
2 78718 1 1963
2 78719 1 1963
2 78720 1 1963
2 78721 1 1963
2 78722 1 1970
2 78723 1 1970
2 78724 1 1970
2 78725 1 1970
2 78726 1 1970
2 78727 1 1970
2 78728 1 1970
2 78729 1 1970
2 78730 1 1970
2 78731 1 1970
2 78732 1 1970
2 78733 1 1970
2 78734 1 1970
2 78735 1 1970
2 78736 1 1970
2 78737 1 1970
2 78738 1 1971
2 78739 1 1971
2 78740 1 1972
2 78741 1 1972
2 78742 1 1972
2 78743 1 1973
2 78744 1 1973
2 78745 1 1974
2 78746 1 1974
2 78747 1 1974
2 78748 1 1974
2 78749 1 1974
2 78750 1 1974
2 78751 1 1974
2 78752 1 1974
2 78753 1 1974
2 78754 1 1974
2 78755 1 1974
2 78756 1 1974
2 78757 1 1974
2 78758 1 1974
2 78759 1 1974
2 78760 1 1974
2 78761 1 1974
2 78762 1 1974
2 78763 1 1974
2 78764 1 1975
2 78765 1 1975
2 78766 1 1983
2 78767 1 1983
2 78768 1 1983
2 78769 1 1983
2 78770 1 1983
2 78771 1 1983
2 78772 1 1983
2 78773 1 1984
2 78774 1 1984
2 78775 1 1984
2 78776 1 1984
2 78777 1 1984
2 78778 1 1984
2 78779 1 1984
2 78780 1 1984
2 78781 1 1984
2 78782 1 1984
2 78783 1 1986
2 78784 1 1986
2 78785 1 1988
2 78786 1 1988
2 78787 1 1989
2 78788 1 1989
2 78789 1 1989
2 78790 1 1989
2 78791 1 1989
2 78792 1 1989
2 78793 1 1989
2 78794 1 1989
2 78795 1 1989
2 78796 1 1989
2 78797 1 1989
2 78798 1 1989
2 78799 1 1989
2 78800 1 1989
2 78801 1 1998
2 78802 1 1998
2 78803 1 1998
2 78804 1 1998
2 78805 1 1998
2 78806 1 1998
2 78807 1 1998
2 78808 1 1998
2 78809 1 1998
2 78810 1 1998
2 78811 1 1998
2 78812 1 1999
2 78813 1 1999
2 78814 1 1999
2 78815 1 1999
2 78816 1 2000
2 78817 1 2000
2 78818 1 2002
2 78819 1 2002
2 78820 1 2002
2 78821 1 2002
2 78822 1 2002
2 78823 1 2002
2 78824 1 2002
2 78825 1 2002
2 78826 1 2002
2 78827 1 2002
2 78828 1 2002
2 78829 1 2002
2 78830 1 2002
2 78831 1 2002
2 78832 1 2002
2 78833 1 2002
2 78834 1 2011
2 78835 1 2011
2 78836 1 2011
2 78837 1 2011
2 78838 1 2011
2 78839 1 2011
2 78840 1 2011
2 78841 1 2011
2 78842 1 2011
2 78843 1 2011
2 78844 1 2011
2 78845 1 2011
2 78846 1 2011
2 78847 1 2011
2 78848 1 2011
2 78849 1 2011
2 78850 1 2011
2 78851 1 2011
2 78852 1 2011
2 78853 1 2011
2 78854 1 2011
2 78855 1 2011
2 78856 1 2012
2 78857 1 2012
2 78858 1 2013
2 78859 1 2013
2 78860 1 2013
2 78861 1 2013
2 78862 1 2013
2 78863 1 2013
2 78864 1 2013
2 78865 1 2013
2 78866 1 2013
2 78867 1 2013
2 78868 1 2013
2 78869 1 2013
2 78870 1 2013
2 78871 1 2013
2 78872 1 2013
2 78873 1 2013
2 78874 1 2013
2 78875 1 2013
2 78876 1 2013
2 78877 1 2013
2 78878 1 2013
2 78879 1 2013
2 78880 1 2013
2 78881 1 2013
2 78882 1 2013
2 78883 1 2013
2 78884 1 2013
2 78885 1 2013
2 78886 1 2013
2 78887 1 2013
2 78888 1 2013
2 78889 1 2013
2 78890 1 2013
2 78891 1 2013
2 78892 1 2013
2 78893 1 2013
2 78894 1 2013
2 78895 1 2013
2 78896 1 2013
2 78897 1 2013
2 78898 1 2014
2 78899 1 2014
2 78900 1 2014
2 78901 1 2014
2 78902 1 2014
2 78903 1 2014
2 78904 1 2015
2 78905 1 2015
2 78906 1 2015
2 78907 1 2015
2 78908 1 2015
2 78909 1 2015
2 78910 1 2015
2 78911 1 2015
2 78912 1 2015
2 78913 1 2015
2 78914 1 2015
2 78915 1 2015
2 78916 1 2015
2 78917 1 2015
2 78918 1 2015
2 78919 1 2015
2 78920 1 2015
2 78921 1 2015
2 78922 1 2015
2 78923 1 2015
2 78924 1 2015
2 78925 1 2015
2 78926 1 2015
2 78927 1 2015
2 78928 1 2015
2 78929 1 2015
2 78930 1 2015
2 78931 1 2015
2 78932 1 2015
2 78933 1 2015
2 78934 1 2015
2 78935 1 2015
2 78936 1 2015
2 78937 1 2015
2 78938 1 2015
2 78939 1 2015
2 78940 1 2017
2 78941 1 2017
2 78942 1 2018
2 78943 1 2018
2 78944 1 2018
2 78945 1 2018
2 78946 1 2018
2 78947 1 2018
2 78948 1 2018
2 78949 1 2018
2 78950 1 2018
2 78951 1 2018
2 78952 1 2018
2 78953 1 2018
2 78954 1 2018
2 78955 1 2018
2 78956 1 2018
2 78957 1 2018
2 78958 1 2018
2 78959 1 2018
2 78960 1 2018
2 78961 1 2018
2 78962 1 2018
2 78963 1 2018
2 78964 1 2018
2 78965 1 2021
2 78966 1 2021
2 78967 1 2021
2 78968 1 2021
2 78969 1 2021
2 78970 1 2021
2 78971 1 2021
2 78972 1 2021
2 78973 1 2023
2 78974 1 2023
2 78975 1 2023
2 78976 1 2027
2 78977 1 2027
2 78978 1 2030
2 78979 1 2030
2 78980 1 2030
2 78981 1 2030
2 78982 1 2030
2 78983 1 2030
2 78984 1 2030
2 78985 1 2030
2 78986 1 2031
2 78987 1 2031
2 78988 1 2031
2 78989 1 2031
2 78990 1 2031
2 78991 1 2031
2 78992 1 2031
2 78993 1 2032
2 78994 1 2032
2 78995 1 2035
2 78996 1 2035
2 78997 1 2035
2 78998 1 2035
2 78999 1 2035
2 79000 1 2036
2 79001 1 2036
2 79002 1 2036
2 79003 1 2036
2 79004 1 2036
2 79005 1 2036
2 79006 1 2036
2 79007 1 2036
2 79008 1 2038
2 79009 1 2038
2 79010 1 2038
2 79011 1 2038
2 79012 1 2038
2 79013 1 2038
2 79014 1 2038
2 79015 1 2038
2 79016 1 2038
2 79017 1 2038
2 79018 1 2039
2 79019 1 2039
2 79020 1 2039
2 79021 1 2039
2 79022 1 2040
2 79023 1 2040
2 79024 1 2041
2 79025 1 2041
2 79026 1 2041
2 79027 1 2041
2 79028 1 2041
2 79029 1 2041
2 79030 1 2041
2 79031 1 2041
2 79032 1 2041
2 79033 1 2050
2 79034 1 2050
2 79035 1 2050
2 79036 1 2050
2 79037 1 2051
2 79038 1 2051
2 79039 1 2051
2 79040 1 2052
2 79041 1 2052
2 79042 1 2052
2 79043 1 2052
2 79044 1 2053
2 79045 1 2053
2 79046 1 2053
2 79047 1 2053
2 79048 1 2055
2 79049 1 2055
2 79050 1 2055
2 79051 1 2055
2 79052 1 2055
2 79053 1 2055
2 79054 1 2055
2 79055 1 2055
2 79056 1 2056
2 79057 1 2056
2 79058 1 2056
2 79059 1 2060
2 79060 1 2060
2 79061 1 2060
2 79062 1 2060
2 79063 1 2060
2 79064 1 2060
2 79065 1 2060
2 79066 1 2060
2 79067 1 2060
2 79068 1 2060
2 79069 1 2060
2 79070 1 2060
2 79071 1 2060
2 79072 1 2060
2 79073 1 2060
2 79074 1 2060
2 79075 1 2060
2 79076 1 2060
2 79077 1 2060
2 79078 1 2060
2 79079 1 2060
2 79080 1 2060
2 79081 1 2060
2 79082 1 2060
2 79083 1 2060
2 79084 1 2060
2 79085 1 2060
2 79086 1 2060
2 79087 1 2060
2 79088 1 2060
2 79089 1 2060
2 79090 1 2060
2 79091 1 2060
2 79092 1 2060
2 79093 1 2060
2 79094 1 2060
2 79095 1 2060
2 79096 1 2060
2 79097 1 2061
2 79098 1 2061
2 79099 1 2061
2 79100 1 2061
2 79101 1 2061
2 79102 1 2061
2 79103 1 2061
2 79104 1 2061
2 79105 1 2061
2 79106 1 2061
2 79107 1 2061
2 79108 1 2061
2 79109 1 2061
2 79110 1 2062
2 79111 1 2062
2 79112 1 2062
2 79113 1 2063
2 79114 1 2063
2 79115 1 2063
2 79116 1 2063
2 79117 1 2063
2 79118 1 2063
2 79119 1 2063
2 79120 1 2063
2 79121 1 2063
2 79122 1 2063
2 79123 1 2063
2 79124 1 2063
2 79125 1 2063
2 79126 1 2063
2 79127 1 2063
2 79128 1 2063
2 79129 1 2063
2 79130 1 2063
2 79131 1 2063
2 79132 1 2063
2 79133 1 2063
2 79134 1 2063
2 79135 1 2063
2 79136 1 2063
2 79137 1 2063
2 79138 1 2063
2 79139 1 2063
2 79140 1 2063
2 79141 1 2063
2 79142 1 2063
2 79143 1 2063
2 79144 1 2063
2 79145 1 2063
2 79146 1 2064
2 79147 1 2064
2 79148 1 2064
2 79149 1 2064
2 79150 1 2064
2 79151 1 2064
2 79152 1 2064
2 79153 1 2064
2 79154 1 2064
2 79155 1 2064
2 79156 1 2064
2 79157 1 2064
2 79158 1 2065
2 79159 1 2065
2 79160 1 2065
2 79161 1 2067
2 79162 1 2067
2 79163 1 2067
2 79164 1 2067
2 79165 1 2067
2 79166 1 2067
2 79167 1 2067
2 79168 1 2067
2 79169 1 2067
2 79170 1 2067
2 79171 1 2067
2 79172 1 2067
2 79173 1 2067
2 79174 1 2067
2 79175 1 2067
2 79176 1 2067
2 79177 1 2067
2 79178 1 2067
2 79179 1 2067
2 79180 1 2067
2 79181 1 2067
2 79182 1 2067
2 79183 1 2067
2 79184 1 2067
2 79185 1 2067
2 79186 1 2067
2 79187 1 2067
2 79188 1 2067
2 79189 1 2067
2 79190 1 2067
2 79191 1 2067
2 79192 1 2067
2 79193 1 2067
2 79194 1 2067
2 79195 1 2067
2 79196 1 2067
2 79197 1 2067
2 79198 1 2067
2 79199 1 2067
2 79200 1 2068
2 79201 1 2068
2 79202 1 2068
2 79203 1 2069
2 79204 1 2069
2 79205 1 2069
2 79206 1 2069
2 79207 1 2069
2 79208 1 2069
2 79209 1 2079
2 79210 1 2079
2 79211 1 2079
2 79212 1 2079
2 79213 1 2079
2 79214 1 2079
2 79215 1 2079
2 79216 1 2080
2 79217 1 2080
2 79218 1 2080
2 79219 1 2080
2 79220 1 2080
2 79221 1 2080
2 79222 1 2080
2 79223 1 2080
2 79224 1 2080
2 79225 1 2080
2 79226 1 2080
2 79227 1 2082
2 79228 1 2082
2 79229 1 2082
2 79230 1 2082
2 79231 1 2082
2 79232 1 2082
2 79233 1 2083
2 79234 1 2083
2 79235 1 2083
2 79236 1 2083
2 79237 1 2083
2 79238 1 2083
2 79239 1 2083
2 79240 1 2083
2 79241 1 2083
2 79242 1 2083
2 79243 1 2083
2 79244 1 2084
2 79245 1 2084
2 79246 1 2084
2 79247 1 2093
2 79248 1 2093
2 79249 1 2093
2 79250 1 2093
2 79251 1 2093
2 79252 1 2093
2 79253 1 2093
2 79254 1 2093
2 79255 1 2093
2 79256 1 2093
2 79257 1 2093
2 79258 1 2093
2 79259 1 2093
2 79260 1 2093
2 79261 1 2093
2 79262 1 2093
2 79263 1 2093
2 79264 1 2093
2 79265 1 2093
2 79266 1 2093
2 79267 1 2093
2 79268 1 2093
2 79269 1 2093
2 79270 1 2093
2 79271 1 2093
2 79272 1 2093
2 79273 1 2093
2 79274 1 2094
2 79275 1 2094
2 79276 1 2095
2 79277 1 2095
2 79278 1 2095
2 79279 1 2095
2 79280 1 2095
2 79281 1 2095
2 79282 1 2095
2 79283 1 2095
2 79284 1 2096
2 79285 1 2096
2 79286 1 2097
2 79287 1 2097
2 79288 1 2097
2 79289 1 2097
2 79290 1 2097
2 79291 1 2097
2 79292 1 2106
2 79293 1 2106
2 79294 1 2106
2 79295 1 2106
2 79296 1 2106
2 79297 1 2106
2 79298 1 2106
2 79299 1 2106
2 79300 1 2106
2 79301 1 2106
2 79302 1 2107
2 79303 1 2107
2 79304 1 2107
2 79305 1 2110
2 79306 1 2110
2 79307 1 2110
2 79308 1 2110
2 79309 1 2110
2 79310 1 2119
2 79311 1 2119
2 79312 1 2132
2 79313 1 2132
2 79314 1 2141
2 79315 1 2141
2 79316 1 2141
2 79317 1 2142
2 79318 1 2142
2 79319 1 2142
2 79320 1 2142
2 79321 1 2142
2 79322 1 2144
2 79323 1 2144
2 79324 1 2144
2 79325 1 2155
2 79326 1 2155
2 79327 1 2155
2 79328 1 2155
2 79329 1 2168
2 79330 1 2168
2 79331 1 2168
2 79332 1 2168
2 79333 1 2168
2 79334 1 2168
2 79335 1 2168
2 79336 1 2168
2 79337 1 2168
2 79338 1 2168
2 79339 1 2168
2 79340 1 2168
2 79341 1 2168
2 79342 1 2168
2 79343 1 2168
2 79344 1 2168
2 79345 1 2168
2 79346 1 2168
2 79347 1 2168
2 79348 1 2168
2 79349 1 2168
2 79350 1 2168
2 79351 1 2168
2 79352 1 2168
2 79353 1 2168
2 79354 1 2168
2 79355 1 2168
2 79356 1 2168
2 79357 1 2168
2 79358 1 2168
2 79359 1 2168
2 79360 1 2168
2 79361 1 2168
2 79362 1 2168
2 79363 1 2168
2 79364 1 2168
2 79365 1 2168
2 79366 1 2168
2 79367 1 2168
2 79368 1 2168
2 79369 1 2168
2 79370 1 2168
2 79371 1 2168
2 79372 1 2168
2 79373 1 2168
2 79374 1 2168
2 79375 1 2168
2 79376 1 2168
2 79377 1 2168
2 79378 1 2168
2 79379 1 2168
2 79380 1 2168
2 79381 1 2168
2 79382 1 2168
2 79383 1 2168
2 79384 1 2168
2 79385 1 2169
2 79386 1 2169
2 79387 1 2169
2 79388 1 2169
2 79389 1 2169
2 79390 1 2170
2 79391 1 2170
2 79392 1 2170
2 79393 1 2170
2 79394 1 2170
2 79395 1 2170
2 79396 1 2170
2 79397 1 2170
2 79398 1 2171
2 79399 1 2171
2 79400 1 2171
2 79401 1 2178
2 79402 1 2178
2 79403 1 2178
2 79404 1 2178
2 79405 1 2178
2 79406 1 2195
2 79407 1 2195
2 79408 1 2196
2 79409 1 2196
2 79410 1 2196
2 79411 1 2196
2 79412 1 2196
2 79413 1 2196
2 79414 1 2196
2 79415 1 2196
2 79416 1 2196
2 79417 1 2196
2 79418 1 2196
2 79419 1 2196
2 79420 1 2196
2 79421 1 2196
2 79422 1 2196
2 79423 1 2196
2 79424 1 2196
2 79425 1 2196
2 79426 1 2196
2 79427 1 2196
2 79428 1 2196
2 79429 1 2196
2 79430 1 2196
2 79431 1 2196
2 79432 1 2196
2 79433 1 2196
2 79434 1 2196
2 79435 1 2196
2 79436 1 2196
2 79437 1 2196
2 79438 1 2196
2 79439 1 2196
2 79440 1 2196
2 79441 1 2196
2 79442 1 2196
2 79443 1 2196
2 79444 1 2196
2 79445 1 2196
2 79446 1 2196
2 79447 1 2196
2 79448 1 2196
2 79449 1 2196
2 79450 1 2196
2 79451 1 2196
2 79452 1 2196
2 79453 1 2196
2 79454 1 2196
2 79455 1 2196
2 79456 1 2196
2 79457 1 2196
2 79458 1 2196
2 79459 1 2196
2 79460 1 2196
2 79461 1 2196
2 79462 1 2197
2 79463 1 2197
2 79464 1 2197
2 79465 1 2197
2 79466 1 2197
2 79467 1 2197
2 79468 1 2198
2 79469 1 2198
2 79470 1 2198
2 79471 1 2198
2 79472 1 2198
2 79473 1 2198
2 79474 1 2198
2 79475 1 2198
2 79476 1 2198
2 79477 1 2198
2 79478 1 2198
2 79479 1 2198
2 79480 1 2200
2 79481 1 2200
2 79482 1 2208
2 79483 1 2208
2 79484 1 2214
2 79485 1 2214
2 79486 1 2215
2 79487 1 2215
2 79488 1 2215
2 79489 1 2215
2 79490 1 2215
2 79491 1 2215
2 79492 1 2215
2 79493 1 2215
2 79494 1 2216
2 79495 1 2216
2 79496 1 2219
2 79497 1 2219
2 79498 1 2219
2 79499 1 2219
2 79500 1 2219
2 79501 1 2219
2 79502 1 2219
2 79503 1 2219
2 79504 1 2219
2 79505 1 2219
2 79506 1 2219
2 79507 1 2220
2 79508 1 2220
2 79509 1 2220
2 79510 1 2220
2 79511 1 2220
2 79512 1 2220
2 79513 1 2220
2 79514 1 2220
2 79515 1 2220
2 79516 1 2220
2 79517 1 2220
2 79518 1 2220
2 79519 1 2220
2 79520 1 2232
2 79521 1 2232
2 79522 1 2232
2 79523 1 2232
2 79524 1 2232
2 79525 1 2238
2 79526 1 2238
2 79527 1 2238
2 79528 1 2238
2 79529 1 2238
2 79530 1 2238
2 79531 1 2238
2 79532 1 2238
2 79533 1 2238
2 79534 1 2238
2 79535 1 2238
2 79536 1 2238
2 79537 1 2238
2 79538 1 2238
2 79539 1 2239
2 79540 1 2239
2 79541 1 2239
2 79542 1 2239
2 79543 1 2239
2 79544 1 2239
2 79545 1 2239
2 79546 1 2239
2 79547 1 2239
2 79548 1 2239
2 79549 1 2239
2 79550 1 2240
2 79551 1 2240
2 79552 1 2248
2 79553 1 2248
2 79554 1 2248
2 79555 1 2248
2 79556 1 2248
2 79557 1 2250
2 79558 1 2250
2 79559 1 2250
2 79560 1 2252
2 79561 1 2252
2 79562 1 2252
2 79563 1 2252
2 79564 1 2261
2 79565 1 2261
2 79566 1 2262
2 79567 1 2262
2 79568 1 2262
2 79569 1 2262
2 79570 1 2262
2 79571 1 2262
2 79572 1 2270
2 79573 1 2270
2 79574 1 2270
2 79575 1 2270
2 79576 1 2270
2 79577 1 2270
2 79578 1 2270
2 79579 1 2270
2 79580 1 2270
2 79581 1 2270
2 79582 1 2270
2 79583 1 2274
2 79584 1 2274
2 79585 1 2295
2 79586 1 2295
2 79587 1 2297
2 79588 1 2297
2 79589 1 2297
2 79590 1 2297
2 79591 1 2297
2 79592 1 2297
2 79593 1 2297
2 79594 1 2305
2 79595 1 2305
2 79596 1 2305
2 79597 1 2305
2 79598 1 2305
2 79599 1 2305
2 79600 1 2305
2 79601 1 2305
2 79602 1 2305
2 79603 1 2305
2 79604 1 2305
2 79605 1 2305
2 79606 1 2305
2 79607 1 2305
2 79608 1 2305
2 79609 1 2305
2 79610 1 2305
2 79611 1 2305
2 79612 1 2305
2 79613 1 2305
2 79614 1 2307
2 79615 1 2307
2 79616 1 2320
2 79617 1 2320
2 79618 1 2320
2 79619 1 2320
2 79620 1 2320
2 79621 1 2320
2 79622 1 2320
2 79623 1 2320
2 79624 1 2322
2 79625 1 2322
2 79626 1 2322
2 79627 1 2322
2 79628 1 2322
2 79629 1 2322
2 79630 1 2322
2 79631 1 2322
2 79632 1 2322
2 79633 1 2324
2 79634 1 2324
2 79635 1 2348
2 79636 1 2348
2 79637 1 2348
2 79638 1 2348
2 79639 1 2348
2 79640 1 2348
2 79641 1 2348
2 79642 1 2348
2 79643 1 2348
2 79644 1 2348
2 79645 1 2348
2 79646 1 2348
2 79647 1 2348
2 79648 1 2349
2 79649 1 2349
2 79650 1 2349
2 79651 1 2374
2 79652 1 2374
2 79653 1 2374
2 79654 1 2374
2 79655 1 2374
2 79656 1 2374
2 79657 1 2374
2 79658 1 2374
2 79659 1 2374
2 79660 1 2374
2 79661 1 2375
2 79662 1 2375
2 79663 1 2375
2 79664 1 2375
2 79665 1 2375
2 79666 1 2375
2 79667 1 2384
2 79668 1 2384
2 79669 1 2384
2 79670 1 2384
2 79671 1 2384
2 79672 1 2391
2 79673 1 2391
2 79674 1 2392
2 79675 1 2392
2 79676 1 2392
2 79677 1 2392
2 79678 1 2392
2 79679 1 2392
2 79680 1 2392
2 79681 1 2392
2 79682 1 2392
2 79683 1 2392
2 79684 1 2392
2 79685 1 2392
2 79686 1 2392
2 79687 1 2393
2 79688 1 2393
2 79689 1 2393
2 79690 1 2393
2 79691 1 2393
2 79692 1 2394
2 79693 1 2394
2 79694 1 2394
2 79695 1 2394
2 79696 1 2394
2 79697 1 2394
2 79698 1 2394
2 79699 1 2394
2 79700 1 2394
2 79701 1 2394
2 79702 1 2394
2 79703 1 2395
2 79704 1 2395
2 79705 1 2397
2 79706 1 2397
2 79707 1 2418
2 79708 1 2418
2 79709 1 2418
2 79710 1 2418
2 79711 1 2419
2 79712 1 2419
2 79713 1 2419
2 79714 1 2419
2 79715 1 2421
2 79716 1 2421
2 79717 1 2421
2 79718 1 2421
2 79719 1 2421
2 79720 1 2421
2 79721 1 2421
2 79722 1 2421
2 79723 1 2421
2 79724 1 2422
2 79725 1 2422
2 79726 1 2426
2 79727 1 2426
2 79728 1 2430
2 79729 1 2430
2 79730 1 2434
2 79731 1 2434
2 79732 1 2434
2 79733 1 2434
2 79734 1 2434
2 79735 1 2434
2 79736 1 2434
2 79737 1 2434
2 79738 1 2434
2 79739 1 2434
2 79740 1 2434
2 79741 1 2435
2 79742 1 2435
2 79743 1 2435
2 79744 1 2435
2 79745 1 2435
2 79746 1 2435
2 79747 1 2435
2 79748 1 2435
2 79749 1 2435
2 79750 1 2435
2 79751 1 2435
2 79752 1 2435
2 79753 1 2435
2 79754 1 2435
2 79755 1 2435
2 79756 1 2435
2 79757 1 2435
2 79758 1 2435
2 79759 1 2436
2 79760 1 2436
2 79761 1 2436
2 79762 1 2436
2 79763 1 2444
2 79764 1 2444
2 79765 1 2444
2 79766 1 2444
2 79767 1 2444
2 79768 1 2444
2 79769 1 2444
2 79770 1 2444
2 79771 1 2444
2 79772 1 2444
2 79773 1 2444
2 79774 1 2444
2 79775 1 2444
2 79776 1 2444
2 79777 1 2444
2 79778 1 2444
2 79779 1 2444
2 79780 1 2444
2 79781 1 2444
2 79782 1 2444
2 79783 1 2444
2 79784 1 2445
2 79785 1 2445
2 79786 1 2445
2 79787 1 2445
2 79788 1 2445
2 79789 1 2446
2 79790 1 2446
2 79791 1 2453
2 79792 1 2453
2 79793 1 2453
2 79794 1 2453
2 79795 1 2453
2 79796 1 2453
2 79797 1 2453
2 79798 1 2453
2 79799 1 2453
2 79800 1 2453
2 79801 1 2453
2 79802 1 2454
2 79803 1 2454
2 79804 1 2454
2 79805 1 2454
2 79806 1 2454
2 79807 1 2454
2 79808 1 2454
2 79809 1 2454
2 79810 1 2454
2 79811 1 2457
2 79812 1 2457
2 79813 1 2457
2 79814 1 2457
2 79815 1 2458
2 79816 1 2458
2 79817 1 2458
2 79818 1 2458
2 79819 1 2458
2 79820 1 2458
2 79821 1 2458
2 79822 1 2458
2 79823 1 2458
2 79824 1 2459
2 79825 1 2459
2 79826 1 2466
2 79827 1 2466
2 79828 1 2466
2 79829 1 2466
2 79830 1 2466
2 79831 1 2466
2 79832 1 2466
2 79833 1 2466
2 79834 1 2466
2 79835 1 2467
2 79836 1 2467
2 79837 1 2467
2 79838 1 2467
2 79839 1 2467
2 79840 1 2468
2 79841 1 2468
2 79842 1 2468
2 79843 1 2470
2 79844 1 2470
2 79845 1 2470
2 79846 1 2470
2 79847 1 2470
2 79848 1 2477
2 79849 1 2477
2 79850 1 2477
2 79851 1 2477
2 79852 1 2477
2 79853 1 2477
2 79854 1 2477
2 79855 1 2477
2 79856 1 2477
2 79857 1 2477
2 79858 1 2477
2 79859 1 2477
2 79860 1 2477
2 79861 1 2477
2 79862 1 2478
2 79863 1 2478
2 79864 1 2478
2 79865 1 2478
2 79866 1 2478
2 79867 1 2478
2 79868 1 2478
2 79869 1 2478
2 79870 1 2478
2 79871 1 2480
2 79872 1 2480
2 79873 1 2481
2 79874 1 2481
2 79875 1 2481
2 79876 1 2481
2 79877 1 2490
2 79878 1 2490
2 79879 1 2490
2 79880 1 2490
2 79881 1 2502
2 79882 1 2502
2 79883 1 2516
2 79884 1 2516
2 79885 1 2516
2 79886 1 2516
2 79887 1 2516
2 79888 1 2516
2 79889 1 2516
2 79890 1 2517
2 79891 1 2517
2 79892 1 2517
2 79893 1 2517
2 79894 1 2517
2 79895 1 2517
2 79896 1 2517
2 79897 1 2517
2 79898 1 2517
2 79899 1 2517
2 79900 1 2517
2 79901 1 2517
2 79902 1 2517
2 79903 1 2517
2 79904 1 2517
2 79905 1 2517
2 79906 1 2517
2 79907 1 2517
2 79908 1 2517
2 79909 1 2517
2 79910 1 2517
2 79911 1 2517
2 79912 1 2517
2 79913 1 2517
2 79914 1 2517
2 79915 1 2517
2 79916 1 2518
2 79917 1 2518
2 79918 1 2518
2 79919 1 2518
2 79920 1 2518
2 79921 1 2518
2 79922 1 2518
2 79923 1 2523
2 79924 1 2523
2 79925 1 2523
2 79926 1 2523
2 79927 1 2523
2 79928 1 2523
2 79929 1 2524
2 79930 1 2524
2 79931 1 2532
2 79932 1 2532
2 79933 1 2532
2 79934 1 2532
2 79935 1 2532
2 79936 1 2532
2 79937 1 2532
2 79938 1 2532
2 79939 1 2532
2 79940 1 2532
2 79941 1 2532
2 79942 1 2532
2 79943 1 2533
2 79944 1 2533
2 79945 1 2533
2 79946 1 2534
2 79947 1 2534
2 79948 1 2535
2 79949 1 2535
2 79950 1 2535
2 79951 1 2535
2 79952 1 2535
2 79953 1 2535
2 79954 1 2535
2 79955 1 2535
2 79956 1 2535
2 79957 1 2535
2 79958 1 2535
2 79959 1 2535
2 79960 1 2535
2 79961 1 2535
2 79962 1 2535
2 79963 1 2535
2 79964 1 2535
2 79965 1 2536
2 79966 1 2536
2 79967 1 2536
2 79968 1 2536
2 79969 1 2536
2 79970 1 2536
2 79971 1 2536
2 79972 1 2537
2 79973 1 2537
2 79974 1 2537
2 79975 1 2538
2 79976 1 2538
2 79977 1 2552
2 79978 1 2552
2 79979 1 2552
2 79980 1 2552
2 79981 1 2552
2 79982 1 2552
2 79983 1 2556
2 79984 1 2556
2 79985 1 2556
2 79986 1 2556
2 79987 1 2556
2 79988 1 2576
2 79989 1 2576
2 79990 1 2576
2 79991 1 2576
2 79992 1 2576
2 79993 1 2576
2 79994 1 2576
2 79995 1 2577
2 79996 1 2577
2 79997 1 2577
2 79998 1 2577
2 79999 1 2577
2 80000 1 2577
2 80001 1 2577
2 80002 1 2577
2 80003 1 2577
2 80004 1 2577
2 80005 1 2577
2 80006 1 2577
2 80007 1 2577
2 80008 1 2577
2 80009 1 2577
2 80010 1 2577
2 80011 1 2577
2 80012 1 2577
2 80013 1 2577
2 80014 1 2577
2 80015 1 2577
2 80016 1 2578
2 80017 1 2578
2 80018 1 2578
2 80019 1 2581
2 80020 1 2581
2 80021 1 2582
2 80022 1 2582
2 80023 1 2582
2 80024 1 2582
2 80025 1 2582
2 80026 1 2582
2 80027 1 2582
2 80028 1 2582
2 80029 1 2582
2 80030 1 2582
2 80031 1 2582
2 80032 1 2582
2 80033 1 2582
2 80034 1 2582
2 80035 1 2582
2 80036 1 2582
2 80037 1 2582
2 80038 1 2583
2 80039 1 2583
2 80040 1 2583
2 80041 1 2583
2 80042 1 2583
2 80043 1 2583
2 80044 1 2583
2 80045 1 2583
2 80046 1 2583
2 80047 1 2583
2 80048 1 2583
2 80049 1 2583
2 80050 1 2583
2 80051 1 2583
2 80052 1 2583
2 80053 1 2583
2 80054 1 2583
2 80055 1 2584
2 80056 1 2584
2 80057 1 2584
2 80058 1 2584
2 80059 1 2584
2 80060 1 2584
2 80061 1 2584
2 80062 1 2592
2 80063 1 2592
2 80064 1 2592
2 80065 1 2592
2 80066 1 2592
2 80067 1 2592
2 80068 1 2592
2 80069 1 2592
2 80070 1 2592
2 80071 1 2592
2 80072 1 2592
2 80073 1 2593
2 80074 1 2593
2 80075 1 2593
2 80076 1 2594
2 80077 1 2594
2 80078 1 2594
2 80079 1 2594
2 80080 1 2594
2 80081 1 2594
2 80082 1 2601
2 80083 1 2601
2 80084 1 2601
2 80085 1 2601
2 80086 1 2601
2 80087 1 2601
2 80088 1 2601
2 80089 1 2601
2 80090 1 2601
2 80091 1 2601
2 80092 1 2601
2 80093 1 2601
2 80094 1 2609
2 80095 1 2609
2 80096 1 2609
2 80097 1 2609
2 80098 1 2609
2 80099 1 2609
2 80100 1 2609
2 80101 1 2609
2 80102 1 2609
2 80103 1 2609
2 80104 1 2611
2 80105 1 2611
2 80106 1 2611
2 80107 1 2611
2 80108 1 2611
2 80109 1 2612
2 80110 1 2612
2 80111 1 2613
2 80112 1 2613
2 80113 1 2613
2 80114 1 2613
2 80115 1 2613
2 80116 1 2613
2 80117 1 2613
2 80118 1 2613
2 80119 1 2613
2 80120 1 2617
2 80121 1 2617
2 80122 1 2620
2 80123 1 2620
2 80124 1 2620
2 80125 1 2620
2 80126 1 2620
2 80127 1 2620
2 80128 1 2620
2 80129 1 2620
2 80130 1 2620
2 80131 1 2620
2 80132 1 2620
2 80133 1 2620
2 80134 1 2620
2 80135 1 2620
2 80136 1 2620
2 80137 1 2620
2 80138 1 2620
2 80139 1 2620
2 80140 1 2620
2 80141 1 2620
2 80142 1 2620
2 80143 1 2620
2 80144 1 2620
2 80145 1 2621
2 80146 1 2621
2 80147 1 2621
2 80148 1 2621
2 80149 1 2621
2 80150 1 2621
2 80151 1 2621
2 80152 1 2621
2 80153 1 2621
2 80154 1 2623
2 80155 1 2623
2 80156 1 2625
2 80157 1 2625
2 80158 1 2632
2 80159 1 2632
2 80160 1 2635
2 80161 1 2635
2 80162 1 2635
2 80163 1 2635
2 80164 1 2635
2 80165 1 2635
2 80166 1 2635
2 80167 1 2635
2 80168 1 2635
2 80169 1 2635
2 80170 1 2635
2 80171 1 2635
2 80172 1 2635
2 80173 1 2635
2 80174 1 2636
2 80175 1 2636
2 80176 1 2637
2 80177 1 2637
2 80178 1 2644
2 80179 1 2644
2 80180 1 2644
2 80181 1 2645
2 80182 1 2645
2 80183 1 2645
2 80184 1 2645
2 80185 1 2645
2 80186 1 2645
2 80187 1 2645
2 80188 1 2645
2 80189 1 2645
2 80190 1 2645
2 80191 1 2645
2 80192 1 2646
2 80193 1 2646
2 80194 1 2646
2 80195 1 2646
2 80196 1 2646
2 80197 1 2646
2 80198 1 2646
2 80199 1 2646
2 80200 1 2646
2 80201 1 2646
2 80202 1 2646
2 80203 1 2646
2 80204 1 2646
2 80205 1 2646
2 80206 1 2646
2 80207 1 2646
2 80208 1 2646
2 80209 1 2646
2 80210 1 2646
2 80211 1 2646
2 80212 1 2646
2 80213 1 2646
2 80214 1 2647
2 80215 1 2647
2 80216 1 2659
2 80217 1 2659
2 80218 1 2659
2 80219 1 2659
2 80220 1 2659
2 80221 1 2659
2 80222 1 2659
2 80223 1 2659
2 80224 1 2659
2 80225 1 2659
2 80226 1 2659
2 80227 1 2659
2 80228 1 2659
2 80229 1 2659
2 80230 1 2661
2 80231 1 2661
2 80232 1 2661
2 80233 1 2661
2 80234 1 2661
2 80235 1 2661
2 80236 1 2665
2 80237 1 2665
2 80238 1 2669
2 80239 1 2669
2 80240 1 2669
2 80241 1 2669
2 80242 1 2669
2 80243 1 2669
2 80244 1 2669
2 80245 1 2669
2 80246 1 2669
2 80247 1 2669
2 80248 1 2669
2 80249 1 2669
2 80250 1 2670
2 80251 1 2670
2 80252 1 2670
2 80253 1 2678
2 80254 1 2678
2 80255 1 2686
2 80256 1 2686
2 80257 1 2686
2 80258 1 2686
2 80259 1 2686
2 80260 1 2686
2 80261 1 2686
2 80262 1 2686
2 80263 1 2686
2 80264 1 2687
2 80265 1 2687
2 80266 1 2689
2 80267 1 2689
2 80268 1 2689
2 80269 1 2689
2 80270 1 2689
2 80271 1 2689
2 80272 1 2689
2 80273 1 2689
2 80274 1 2691
2 80275 1 2691
2 80276 1 2691
2 80277 1 2700
2 80278 1 2700
2 80279 1 2700
2 80280 1 2700
2 80281 1 2700
2 80282 1 2700
2 80283 1 2700
2 80284 1 2700
2 80285 1 2700
2 80286 1 2700
2 80287 1 2700
2 80288 1 2702
2 80289 1 2702
2 80290 1 2702
2 80291 1 2702
2 80292 1 2702
2 80293 1 2702
2 80294 1 2702
2 80295 1 2702
2 80296 1 2702
2 80297 1 2702
2 80298 1 2702
2 80299 1 2702
2 80300 1 2702
2 80301 1 2702
2 80302 1 2702
2 80303 1 2702
2 80304 1 2702
2 80305 1 2702
2 80306 1 2702
2 80307 1 2702
2 80308 1 2702
2 80309 1 2702
2 80310 1 2702
2 80311 1 2702
2 80312 1 2704
2 80313 1 2704
2 80314 1 2704
2 80315 1 2707
2 80316 1 2707
2 80317 1 2707
2 80318 1 2715
2 80319 1 2715
2 80320 1 2715
2 80321 1 2715
2 80322 1 2715
2 80323 1 2715
2 80324 1 2715
2 80325 1 2715
2 80326 1 2715
2 80327 1 2715
2 80328 1 2715
2 80329 1 2715
2 80330 1 2716
2 80331 1 2716
2 80332 1 2716
2 80333 1 2716
2 80334 1 2717
2 80335 1 2717
2 80336 1 2721
2 80337 1 2721
2 80338 1 2736
2 80339 1 2736
2 80340 1 2736
2 80341 1 2736
2 80342 1 2736
2 80343 1 2736
2 80344 1 2736
2 80345 1 2736
2 80346 1 2736
2 80347 1 2736
2 80348 1 2736
2 80349 1 2736
2 80350 1 2736
2 80351 1 2736
2 80352 1 2736
2 80353 1 2737
2 80354 1 2737
2 80355 1 2737
2 80356 1 2738
2 80357 1 2738
2 80358 1 2738
2 80359 1 2738
2 80360 1 2740
2 80361 1 2740
2 80362 1 2740
2 80363 1 2742
2 80364 1 2742
2 80365 1 2745
2 80366 1 2745
2 80367 1 2747
2 80368 1 2747
2 80369 1 2747
2 80370 1 2749
2 80371 1 2749
2 80372 1 2750
2 80373 1 2750
2 80374 1 2752
2 80375 1 2752
2 80376 1 2760
2 80377 1 2760
2 80378 1 2760
2 80379 1 2761
2 80380 1 2761
2 80381 1 2761
2 80382 1 2761
2 80383 1 2761
2 80384 1 2761
2 80385 1 2761
2 80386 1 2761
2 80387 1 2761
2 80388 1 2761
2 80389 1 2762
2 80390 1 2762
2 80391 1 2762
2 80392 1 2762
2 80393 1 2763
2 80394 1 2763
2 80395 1 2766
2 80396 1 2766
2 80397 1 2766
2 80398 1 2766
2 80399 1 2766
2 80400 1 2766
2 80401 1 2768
2 80402 1 2768
2 80403 1 2776
2 80404 1 2776
2 80405 1 2776
2 80406 1 2776
2 80407 1 2776
2 80408 1 2776
2 80409 1 2776
2 80410 1 2776
2 80411 1 2776
2 80412 1 2776
2 80413 1 2776
2 80414 1 2776
2 80415 1 2777
2 80416 1 2777
2 80417 1 2777
2 80418 1 2777
2 80419 1 2778
2 80420 1 2778
2 80421 1 2778
2 80422 1 2778
2 80423 1 2781
2 80424 1 2781
2 80425 1 2784
2 80426 1 2784
2 80427 1 2784
2 80428 1 2791
2 80429 1 2791
2 80430 1 2791
2 80431 1 2791
2 80432 1 2793
2 80433 1 2793
2 80434 1 2793
2 80435 1 2793
2 80436 1 2793
2 80437 1 2793
2 80438 1 2793
2 80439 1 2793
2 80440 1 2793
2 80441 1 2793
2 80442 1 2793
2 80443 1 2793
2 80444 1 2793
2 80445 1 2807
2 80446 1 2807
2 80447 1 2807
2 80448 1 2807
2 80449 1 2807
2 80450 1 2808
2 80451 1 2808
2 80452 1 2808
2 80453 1 2809
2 80454 1 2809
2 80455 1 2809
2 80456 1 2809
2 80457 1 2809
2 80458 1 2809
2 80459 1 2809
2 80460 1 2809
2 80461 1 2810
2 80462 1 2810
2 80463 1 2810
2 80464 1 2828
2 80465 1 2828
2 80466 1 2828
2 80467 1 2828
2 80468 1 2828
2 80469 1 2828
2 80470 1 2828
2 80471 1 2828
2 80472 1 2828
2 80473 1 2828
2 80474 1 2828
2 80475 1 2828
2 80476 1 2828
2 80477 1 2828
2 80478 1 2829
2 80479 1 2829
2 80480 1 2830
2 80481 1 2830
2 80482 1 2830
2 80483 1 2830
2 80484 1 2830
2 80485 1 2830
2 80486 1 2830
2 80487 1 2830
2 80488 1 2830
2 80489 1 2830
2 80490 1 2831
2 80491 1 2831
2 80492 1 2831
2 80493 1 2835
2 80494 1 2835
2 80495 1 2835
2 80496 1 2835
2 80497 1 2835
2 80498 1 2835
2 80499 1 2835
2 80500 1 2835
2 80501 1 2835
2 80502 1 2835
2 80503 1 2836
2 80504 1 2836
2 80505 1 2836
2 80506 1 2836
2 80507 1 2836
2 80508 1 2836
2 80509 1 2836
2 80510 1 2850
2 80511 1 2850
2 80512 1 2850
2 80513 1 2850
2 80514 1 2850
2 80515 1 2850
2 80516 1 2851
2 80517 1 2851
2 80518 1 2851
2 80519 1 2851
2 80520 1 2851
2 80521 1 2851
2 80522 1 2854
2 80523 1 2854
2 80524 1 2855
2 80525 1 2855
2 80526 1 2856
2 80527 1 2856
2 80528 1 2864
2 80529 1 2864
2 80530 1 2864
2 80531 1 2864
2 80532 1 2864
2 80533 1 2864
2 80534 1 2865
2 80535 1 2865
2 80536 1 2865
2 80537 1 2865
2 80538 1 2865
2 80539 1 2865
2 80540 1 2866
2 80541 1 2866
2 80542 1 2866
2 80543 1 2866
2 80544 1 2866
2 80545 1 2867
2 80546 1 2867
2 80547 1 2867
2 80548 1 2867
2 80549 1 2867
2 80550 1 2867
2 80551 1 2867
2 80552 1 2867
2 80553 1 2868
2 80554 1 2868
2 80555 1 2868
2 80556 1 2868
2 80557 1 2868
2 80558 1 2868
2 80559 1 2868
2 80560 1 2868
2 80561 1 2868
2 80562 1 2869
2 80563 1 2869
2 80564 1 2869
2 80565 1 2869
2 80566 1 2871
2 80567 1 2871
2 80568 1 2871
2 80569 1 2871
2 80570 1 2871
2 80571 1 2871
2 80572 1 2871
2 80573 1 2871
2 80574 1 2871
2 80575 1 2871
2 80576 1 2871
2 80577 1 2871
2 80578 1 2871
2 80579 1 2871
2 80580 1 2871
2 80581 1 2871
2 80582 1 2871
2 80583 1 2871
2 80584 1 2871
2 80585 1 2871
2 80586 1 2871
2 80587 1 2871
2 80588 1 2871
2 80589 1 2871
2 80590 1 2871
2 80591 1 2871
2 80592 1 2871
2 80593 1 2871
2 80594 1 2871
2 80595 1 2871
2 80596 1 2871
2 80597 1 2871
2 80598 1 2875
2 80599 1 2875
2 80600 1 2875
2 80601 1 2883
2 80602 1 2883
2 80603 1 2883
2 80604 1 2883
2 80605 1 2883
2 80606 1 2883
2 80607 1 2883
2 80608 1 2883
2 80609 1 2883
2 80610 1 2883
2 80611 1 2883
2 80612 1 2884
2 80613 1 2884
2 80614 1 2884
2 80615 1 2884
2 80616 1 2884
2 80617 1 2884
2 80618 1 2884
2 80619 1 2884
2 80620 1 2890
2 80621 1 2890
2 80622 1 2890
2 80623 1 2890
2 80624 1 2890
2 80625 1 2890
2 80626 1 2890
2 80627 1 2890
2 80628 1 2890
2 80629 1 2890
2 80630 1 2890
2 80631 1 2890
2 80632 1 2890
2 80633 1 2890
2 80634 1 2890
2 80635 1 2897
2 80636 1 2897
2 80637 1 2897
2 80638 1 2900
2 80639 1 2900
2 80640 1 2900
2 80641 1 2908
2 80642 1 2908
2 80643 1 2908
2 80644 1 2908
2 80645 1 2908
2 80646 1 2908
2 80647 1 2908
2 80648 1 2908
2 80649 1 2908
2 80650 1 2908
2 80651 1 2908
2 80652 1 2908
2 80653 1 2908
2 80654 1 2908
2 80655 1 2908
2 80656 1 2908
2 80657 1 2909
2 80658 1 2909
2 80659 1 2909
2 80660 1 2909
2 80661 1 2910
2 80662 1 2910
2 80663 1 2910
2 80664 1 2911
2 80665 1 2911
2 80666 1 2918
2 80667 1 2918
2 80668 1 2918
2 80669 1 2918
2 80670 1 2918
2 80671 1 2918
2 80672 1 2918
2 80673 1 2918
2 80674 1 2918
2 80675 1 2919
2 80676 1 2919
2 80677 1 2919
2 80678 1 2919
2 80679 1 2919
2 80680 1 2919
2 80681 1 2919
2 80682 1 2919
2 80683 1 2919
2 80684 1 2919
2 80685 1 2920
2 80686 1 2920
2 80687 1 2927
2 80688 1 2927
2 80689 1 2927
2 80690 1 2927
2 80691 1 2927
2 80692 1 2927
2 80693 1 2927
2 80694 1 2927
2 80695 1 2927
2 80696 1 2928
2 80697 1 2928
2 80698 1 2932
2 80699 1 2932
2 80700 1 2932
2 80701 1 2932
2 80702 1 2932
2 80703 1 2932
2 80704 1 2932
2 80705 1 2932
2 80706 1 2932
2 80707 1 2932
2 80708 1 2932
2 80709 1 2932
2 80710 1 2932
2 80711 1 2932
2 80712 1 2932
2 80713 1 2932
2 80714 1 2932
2 80715 1 2933
2 80716 1 2933
2 80717 1 2933
2 80718 1 2933
2 80719 1 2934
2 80720 1 2934
2 80721 1 2942
2 80722 1 2942
2 80723 1 2942
2 80724 1 2942
2 80725 1 2942
2 80726 1 2942
2 80727 1 2942
2 80728 1 2942
2 80729 1 2942
2 80730 1 2942
2 80731 1 2942
2 80732 1 2942
2 80733 1 2942
2 80734 1 2942
2 80735 1 2942
2 80736 1 2943
2 80737 1 2943
2 80738 1 2943
2 80739 1 2943
2 80740 1 2943
2 80741 1 2943
2 80742 1 2943
2 80743 1 2943
2 80744 1 2943
2 80745 1 2943
2 80746 1 2943
2 80747 1 2943
2 80748 1 2943
2 80749 1 2943
2 80750 1 2944
2 80751 1 2944
2 80752 1 2945
2 80753 1 2945
2 80754 1 2945
2 80755 1 2945
2 80756 1 2945
2 80757 1 2945
2 80758 1 2953
2 80759 1 2953
2 80760 1 2953
2 80761 1 2953
2 80762 1 2953
2 80763 1 2953
2 80764 1 2953
2 80765 1 2955
2 80766 1 2955
2 80767 1 2955
2 80768 1 2955
2 80769 1 2955
2 80770 1 2955
2 80771 1 2955
2 80772 1 2955
2 80773 1 2955
2 80774 1 2955
2 80775 1 2955
2 80776 1 2956
2 80777 1 2956
2 80778 1 2968
2 80779 1 2968
2 80780 1 2968
2 80781 1 2968
2 80782 1 2968
2 80783 1 2968
2 80784 1 2968
2 80785 1 2968
2 80786 1 2968
2 80787 1 2968
2 80788 1 2968
2 80789 1 2968
2 80790 1 2968
2 80791 1 2968
2 80792 1 2968
2 80793 1 2968
2 80794 1 2968
2 80795 1 2968
2 80796 1 2968
2 80797 1 2968
2 80798 1 2969
2 80799 1 2969
2 80800 1 2969
2 80801 1 2969
2 80802 1 2969
2 80803 1 2969
2 80804 1 2969
2 80805 1 2969
2 80806 1 2969
2 80807 1 2969
2 80808 1 2969
2 80809 1 2973
2 80810 1 2973
2 80811 1 2974
2 80812 1 2974
2 80813 1 2974
2 80814 1 2974
2 80815 1 2974
2 80816 1 2983
2 80817 1 2983
2 80818 1 2984
2 80819 1 2984
2 80820 1 2984
2 80821 1 2984
2 80822 1 2984
2 80823 1 2984
2 80824 1 2984
2 80825 1 2984
2 80826 1 2984
2 80827 1 2984
2 80828 1 2985
2 80829 1 2985
2 80830 1 2985
2 80831 1 2994
2 80832 1 2994
2 80833 1 2994
2 80834 1 2994
2 80835 1 2994
2 80836 1 2994
2 80837 1 2994
2 80838 1 2994
2 80839 1 2994
2 80840 1 2994
2 80841 1 2994
2 80842 1 2995
2 80843 1 2995
2 80844 1 2996
2 80845 1 2996
2 80846 1 2996
2 80847 1 2996
2 80848 1 2996
2 80849 1 2996
2 80850 1 2996
2 80851 1 2996
2 80852 1 2996
2 80853 1 2996
2 80854 1 2996
2 80855 1 2997
2 80856 1 2997
2 80857 1 2997
2 80858 1 2997
2 80859 1 2997
2 80860 1 2997
2 80861 1 2997
2 80862 1 2997
2 80863 1 2997
2 80864 1 3006
2 80865 1 3006
2 80866 1 3006
2 80867 1 3006
2 80868 1 3006
2 80869 1 3006
2 80870 1 3006
2 80871 1 3006
2 80872 1 3006
2 80873 1 3006
2 80874 1 3006
2 80875 1 3006
2 80876 1 3006
2 80877 1 3006
2 80878 1 3006
2 80879 1 3006
2 80880 1 3007
2 80881 1 3007
2 80882 1 3007
2 80883 1 3009
2 80884 1 3009
2 80885 1 3010
2 80886 1 3010
2 80887 1 3019
2 80888 1 3019
2 80889 1 3019
2 80890 1 3019
2 80891 1 3020
2 80892 1 3020
2 80893 1 3029
2 80894 1 3029
2 80895 1 3029
2 80896 1 3029
2 80897 1 3029
2 80898 1 3029
2 80899 1 3029
2 80900 1 3032
2 80901 1 3032
2 80902 1 3035
2 80903 1 3035
2 80904 1 3035
2 80905 1 3035
2 80906 1 3035
2 80907 1 3035
2 80908 1 3035
2 80909 1 3035
2 80910 1 3035
2 80911 1 3035
2 80912 1 3035
2 80913 1 3035
2 80914 1 3036
2 80915 1 3036
2 80916 1 3036
2 80917 1 3037
2 80918 1 3037
2 80919 1 3037
2 80920 1 3037
2 80921 1 3037
2 80922 1 3037
2 80923 1 3037
2 80924 1 3037
2 80925 1 3037
2 80926 1 3037
2 80927 1 3037
2 80928 1 3037
2 80929 1 3037
2 80930 1 3037
2 80931 1 3037
2 80932 1 3037
2 80933 1 3037
2 80934 1 3037
2 80935 1 3037
2 80936 1 3037
2 80937 1 3037
2 80938 1 3037
2 80939 1 3037
2 80940 1 3037
2 80941 1 3037
2 80942 1 3037
2 80943 1 3037
2 80944 1 3038
2 80945 1 3038
2 80946 1 3038
2 80947 1 3038
2 80948 1 3038
2 80949 1 3038
2 80950 1 3038
2 80951 1 3038
2 80952 1 3038
2 80953 1 3038
2 80954 1 3039
2 80955 1 3039
2 80956 1 3047
2 80957 1 3047
2 80958 1 3047
2 80959 1 3047
2 80960 1 3047
2 80961 1 3047
2 80962 1 3047
2 80963 1 3047
2 80964 1 3047
2 80965 1 3047
2 80966 1 3047
2 80967 1 3047
2 80968 1 3047
2 80969 1 3047
2 80970 1 3047
2 80971 1 3047
2 80972 1 3047
2 80973 1 3047
2 80974 1 3047
2 80975 1 3047
2 80976 1 3047
2 80977 1 3047
2 80978 1 3047
2 80979 1 3047
2 80980 1 3047
2 80981 1 3047
2 80982 1 3047
2 80983 1 3047
2 80984 1 3047
2 80985 1 3047
2 80986 1 3047
2 80987 1 3047
2 80988 1 3047
2 80989 1 3047
2 80990 1 3047
2 80991 1 3047
2 80992 1 3047
2 80993 1 3047
2 80994 1 3047
2 80995 1 3047
2 80996 1 3047
2 80997 1 3047
2 80998 1 3047
2 80999 1 3047
2 81000 1 3047
2 81001 1 3047
2 81002 1 3047
2 81003 1 3048
2 81004 1 3048
2 81005 1 3048
2 81006 1 3049
2 81007 1 3049
2 81008 1 3049
2 81009 1 3049
2 81010 1 3049
2 81011 1 3049
2 81012 1 3049
2 81013 1 3049
2 81014 1 3050
2 81015 1 3050
2 81016 1 3050
2 81017 1 3050
2 81018 1 3050
2 81019 1 3050
2 81020 1 3051
2 81021 1 3051
2 81022 1 3055
2 81023 1 3055
2 81024 1 3055
2 81025 1 3055
2 81026 1 3055
2 81027 1 3055
2 81028 1 3055
2 81029 1 3056
2 81030 1 3056
2 81031 1 3057
2 81032 1 3057
2 81033 1 3057
2 81034 1 3058
2 81035 1 3058
2 81036 1 3059
2 81037 1 3059
2 81038 1 3059
2 81039 1 3059
2 81040 1 3059
2 81041 1 3059
2 81042 1 3059
2 81043 1 3059
2 81044 1 3059
2 81045 1 3059
2 81046 1 3059
2 81047 1 3059
2 81048 1 3059
2 81049 1 3059
2 81050 1 3059
2 81051 1 3059
2 81052 1 3059
2 81053 1 3059
2 81054 1 3059
2 81055 1 3059
2 81056 1 3059
2 81057 1 3059
2 81058 1 3059
2 81059 1 3060
2 81060 1 3060
2 81061 1 3060
2 81062 1 3060
2 81063 1 3061
2 81064 1 3061
2 81065 1 3061
2 81066 1 3062
2 81067 1 3062
2 81068 1 3065
2 81069 1 3065
2 81070 1 3065
2 81071 1 3065
2 81072 1 3065
2 81073 1 3065
2 81074 1 3066
2 81075 1 3066
2 81076 1 3081
2 81077 1 3081
2 81078 1 3081
2 81079 1 3081
2 81080 1 3081
2 81081 1 3081
2 81082 1 3081
2 81083 1 3081
2 81084 1 3081
2 81085 1 3081
2 81086 1 3081
2 81087 1 3081
2 81088 1 3081
2 81089 1 3081
2 81090 1 3081
2 81091 1 3081
2 81092 1 3081
2 81093 1 3081
2 81094 1 3081
2 81095 1 3081
2 81096 1 3081
2 81097 1 3081
2 81098 1 3081
2 81099 1 3081
2 81100 1 3081
2 81101 1 3081
2 81102 1 3081
2 81103 1 3081
2 81104 1 3081
2 81105 1 3081
2 81106 1 3081
2 81107 1 3081
2 81108 1 3081
2 81109 1 3081
2 81110 1 3081
2 81111 1 3081
2 81112 1 3081
2 81113 1 3081
2 81114 1 3081
2 81115 1 3081
2 81116 1 3082
2 81117 1 3082
2 81118 1 3082
2 81119 1 3083
2 81120 1 3083
2 81121 1 3083
2 81122 1 3083
2 81123 1 3083
2 81124 1 3083
2 81125 1 3083
2 81126 1 3083
2 81127 1 3083
2 81128 1 3083
2 81129 1 3083
2 81130 1 3083
2 81131 1 3083
2 81132 1 3083
2 81133 1 3085
2 81134 1 3085
2 81135 1 3085
2 81136 1 3107
2 81137 1 3107
2 81138 1 3108
2 81139 1 3108
2 81140 1 3109
2 81141 1 3109
2 81142 1 3121
2 81143 1 3121
2 81144 1 3121
2 81145 1 3129
2 81146 1 3129
2 81147 1 3129
2 81148 1 3129
2 81149 1 3129
2 81150 1 3129
2 81151 1 3129
2 81152 1 3129
2 81153 1 3129
2 81154 1 3130
2 81155 1 3130
2 81156 1 3131
2 81157 1 3131
2 81158 1 3136
2 81159 1 3136
2 81160 1 3136
2 81161 1 3136
2 81162 1 3136
2 81163 1 3136
2 81164 1 3137
2 81165 1 3137
2 81166 1 3138
2 81167 1 3138
2 81168 1 3139
2 81169 1 3139
2 81170 1 3141
2 81171 1 3141
2 81172 1 3141
2 81173 1 3141
2 81174 1 3143
2 81175 1 3143
2 81176 1 3147
2 81177 1 3147
2 81178 1 3147
2 81179 1 3159
2 81180 1 3159
2 81181 1 3159
2 81182 1 3159
2 81183 1 3159
2 81184 1 3161
2 81185 1 3161
2 81186 1 3161
2 81187 1 3176
2 81188 1 3176
2 81189 1 3176
2 81190 1 3176
2 81191 1 3180
2 81192 1 3180
2 81193 1 3180
2 81194 1 3181
2 81195 1 3181
2 81196 1 3189
2 81197 1 3189
2 81198 1 3189
2 81199 1 3189
2 81200 1 3189
2 81201 1 3190
2 81202 1 3190
2 81203 1 3190
2 81204 1 3190
2 81205 1 3190
2 81206 1 3191
2 81207 1 3191
2 81208 1 3191
2 81209 1 3191
2 81210 1 3191
2 81211 1 3191
2 81212 1 3191
2 81213 1 3191
2 81214 1 3191
2 81215 1 3191
2 81216 1 3191
2 81217 1 3192
2 81218 1 3192
2 81219 1 3192
2 81220 1 3193
2 81221 1 3193
2 81222 1 3204
2 81223 1 3204
2 81224 1 3205
2 81225 1 3205
2 81226 1 3207
2 81227 1 3207
2 81228 1 3229
2 81229 1 3229
2 81230 1 3229
2 81231 1 3231
2 81232 1 3231
2 81233 1 3237
2 81234 1 3237
2 81235 1 3237
2 81236 1 3237
2 81237 1 3237
2 81238 1 3238
2 81239 1 3238
2 81240 1 3238
2 81241 1 3238
2 81242 1 3238
2 81243 1 3238
2 81244 1 3238
2 81245 1 3238
2 81246 1 3238
2 81247 1 3238
2 81248 1 3238
2 81249 1 3238
2 81250 1 3238
2 81251 1 3238
2 81252 1 3238
2 81253 1 3238
2 81254 1 3253
2 81255 1 3253
2 81256 1 3253
2 81257 1 3253
2 81258 1 3253
2 81259 1 3253
2 81260 1 3253
2 81261 1 3253
2 81262 1 3253
2 81263 1 3253
2 81264 1 3253
2 81265 1 3253
2 81266 1 3253
2 81267 1 3253
2 81268 1 3253
2 81269 1 3253
2 81270 1 3255
2 81271 1 3255
2 81272 1 3255
2 81273 1 3255
2 81274 1 3255
2 81275 1 3255
2 81276 1 3255
2 81277 1 3255
2 81278 1 3255
2 81279 1 3255
2 81280 1 3255
2 81281 1 3255
2 81282 1 3255
2 81283 1 3255
2 81284 1 3255
2 81285 1 3255
2 81286 1 3255
2 81287 1 3255
2 81288 1 3256
2 81289 1 3256
2 81290 1 3257
2 81291 1 3257
2 81292 1 3257
2 81293 1 3257
2 81294 1 3257
2 81295 1 3257
2 81296 1 3257
2 81297 1 3257
2 81298 1 3257
2 81299 1 3257
2 81300 1 3257
2 81301 1 3257
2 81302 1 3257
2 81303 1 3257
2 81304 1 3257
2 81305 1 3257
2 81306 1 3257
2 81307 1 3257
2 81308 1 3257
2 81309 1 3257
2 81310 1 3258
2 81311 1 3258
2 81312 1 3258
2 81313 1 3260
2 81314 1 3260
2 81315 1 3260
2 81316 1 3260
2 81317 1 3260
2 81318 1 3260
2 81319 1 3263
2 81320 1 3263
2 81321 1 3263
2 81322 1 3263
2 81323 1 3263
2 81324 1 3263
2 81325 1 3263
2 81326 1 3263
2 81327 1 3263
2 81328 1 3263
2 81329 1 3263
2 81330 1 3263
2 81331 1 3264
2 81332 1 3264
2 81333 1 3264
2 81334 1 3264
2 81335 1 3265
2 81336 1 3265
2 81337 1 3265
2 81338 1 3265
2 81339 1 3265
2 81340 1 3265
2 81341 1 3265
2 81342 1 3265
2 81343 1 3265
2 81344 1 3265
2 81345 1 3265
2 81346 1 3265
2 81347 1 3265
2 81348 1 3265
2 81349 1 3266
2 81350 1 3266
2 81351 1 3273
2 81352 1 3273
2 81353 1 3273
2 81354 1 3273
2 81355 1 3273
2 81356 1 3273
2 81357 1 3273
2 81358 1 3273
2 81359 1 3273
2 81360 1 3273
2 81361 1 3274
2 81362 1 3274
2 81363 1 3274
2 81364 1 3282
2 81365 1 3282
2 81366 1 3282
2 81367 1 3282
2 81368 1 3282
2 81369 1 3282
2 81370 1 3282
2 81371 1 3282
2 81372 1 3282
2 81373 1 3282
2 81374 1 3282
2 81375 1 3283
2 81376 1 3283
2 81377 1 3283
2 81378 1 3285
2 81379 1 3285
2 81380 1 3295
2 81381 1 3295
2 81382 1 3295
2 81383 1 3295
2 81384 1 3298
2 81385 1 3298
2 81386 1 3298
2 81387 1 3298
2 81388 1 3298
2 81389 1 3298
2 81390 1 3298
2 81391 1 3298
2 81392 1 3298
2 81393 1 3298
2 81394 1 3298
2 81395 1 3298
2 81396 1 3298
2 81397 1 3301
2 81398 1 3301
2 81399 1 3301
2 81400 1 3301
2 81401 1 3301
2 81402 1 3301
2 81403 1 3301
2 81404 1 3302
2 81405 1 3302
2 81406 1 3302
2 81407 1 3302
2 81408 1 3302
2 81409 1 3302
2 81410 1 3302
2 81411 1 3302
2 81412 1 3302
2 81413 1 3302
2 81414 1 3302
2 81415 1 3302
2 81416 1 3302
2 81417 1 3302
2 81418 1 3302
2 81419 1 3302
2 81420 1 3302
2 81421 1 3302
2 81422 1 3302
2 81423 1 3303
2 81424 1 3303
2 81425 1 3303
2 81426 1 3303
2 81427 1 3303
2 81428 1 3304
2 81429 1 3304
2 81430 1 3311
2 81431 1 3311
2 81432 1 3311
2 81433 1 3311
2 81434 1 3311
2 81435 1 3311
2 81436 1 3311
2 81437 1 3311
2 81438 1 3311
2 81439 1 3311
2 81440 1 3311
2 81441 1 3311
2 81442 1 3311
2 81443 1 3311
2 81444 1 3311
2 81445 1 3311
2 81446 1 3311
2 81447 1 3311
2 81448 1 3311
2 81449 1 3311
2 81450 1 3311
2 81451 1 3311
2 81452 1 3311
2 81453 1 3311
2 81454 1 3311
2 81455 1 3311
2 81456 1 3311
2 81457 1 3311
2 81458 1 3311
2 81459 1 3311
2 81460 1 3311
2 81461 1 3311
2 81462 1 3311
2 81463 1 3311
2 81464 1 3313
2 81465 1 3313
2 81466 1 3326
2 81467 1 3326
2 81468 1 3326
2 81469 1 3326
2 81470 1 3326
2 81471 1 3326
2 81472 1 3326
2 81473 1 3326
2 81474 1 3326
2 81475 1 3326
2 81476 1 3326
2 81477 1 3326
2 81478 1 3326
2 81479 1 3326
2 81480 1 3327
2 81481 1 3327
2 81482 1 3328
2 81483 1 3328
2 81484 1 3328
2 81485 1 3328
2 81486 1 3328
2 81487 1 3328
2 81488 1 3328
2 81489 1 3328
2 81490 1 3328
2 81491 1 3328
2 81492 1 3328
2 81493 1 3328
2 81494 1 3329
2 81495 1 3329
2 81496 1 3332
2 81497 1 3332
2 81498 1 3332
2 81499 1 3332
2 81500 1 3333
2 81501 1 3333
2 81502 1 3333
2 81503 1 3333
2 81504 1 3341
2 81505 1 3341
2 81506 1 3341
2 81507 1 3342
2 81508 1 3342
2 81509 1 3343
2 81510 1 3343
2 81511 1 3344
2 81512 1 3344
2 81513 1 3344
2 81514 1 3344
2 81515 1 3344
2 81516 1 3344
2 81517 1 3344
2 81518 1 3344
2 81519 1 3344
2 81520 1 3344
2 81521 1 3344
2 81522 1 3344
2 81523 1 3345
2 81524 1 3345
2 81525 1 3345
2 81526 1 3346
2 81527 1 3346
2 81528 1 3346
2 81529 1 3346
2 81530 1 3346
2 81531 1 3346
2 81532 1 3346
2 81533 1 3346
2 81534 1 3346
2 81535 1 3346
2 81536 1 3346
2 81537 1 3346
2 81538 1 3346
2 81539 1 3355
2 81540 1 3355
2 81541 1 3355
2 81542 1 3355
2 81543 1 3355
2 81544 1 3355
2 81545 1 3355
2 81546 1 3355
2 81547 1 3355
2 81548 1 3355
2 81549 1 3355
2 81550 1 3355
2 81551 1 3355
2 81552 1 3355
2 81553 1 3355
2 81554 1 3355
2 81555 1 3355
2 81556 1 3355
2 81557 1 3355
2 81558 1 3355
2 81559 1 3355
2 81560 1 3355
2 81561 1 3356
2 81562 1 3356
2 81563 1 3356
2 81564 1 3359
2 81565 1 3359
2 81566 1 3359
2 81567 1 3359
2 81568 1 3359
2 81569 1 3359
2 81570 1 3360
2 81571 1 3360
2 81572 1 3360
2 81573 1 3367
2 81574 1 3367
2 81575 1 3368
2 81576 1 3368
2 81577 1 3368
2 81578 1 3368
2 81579 1 3368
2 81580 1 3368
2 81581 1 3368
2 81582 1 3368
2 81583 1 3368
2 81584 1 3368
2 81585 1 3368
2 81586 1 3368
2 81587 1 3368
2 81588 1 3368
2 81589 1 3368
2 81590 1 3368
2 81591 1 3368
2 81592 1 3368
2 81593 1 3368
2 81594 1 3368
2 81595 1 3368
2 81596 1 3368
2 81597 1 3368
2 81598 1 3368
2 81599 1 3368
2 81600 1 3369
2 81601 1 3369
2 81602 1 3369
2 81603 1 3376
2 81604 1 3376
2 81605 1 3377
2 81606 1 3377
2 81607 1 3377
2 81608 1 3377
2 81609 1 3377
2 81610 1 3377
2 81611 1 3377
2 81612 1 3377
2 81613 1 3377
2 81614 1 3377
2 81615 1 3377
2 81616 1 3377
2 81617 1 3377
2 81618 1 3377
2 81619 1 3377
2 81620 1 3377
2 81621 1 3377
2 81622 1 3377
2 81623 1 3377
2 81624 1 3377
2 81625 1 3377
2 81626 1 3377
2 81627 1 3377
2 81628 1 3377
2 81629 1 3377
2 81630 1 3377
2 81631 1 3377
2 81632 1 3377
2 81633 1 3377
2 81634 1 3377
2 81635 1 3377
2 81636 1 3377
2 81637 1 3377
2 81638 1 3377
2 81639 1 3377
2 81640 1 3377
2 81641 1 3377
2 81642 1 3377
2 81643 1 3377
2 81644 1 3377
2 81645 1 3378
2 81646 1 3378
2 81647 1 3378
2 81648 1 3378
2 81649 1 3378
2 81650 1 3378
2 81651 1 3378
2 81652 1 3378
2 81653 1 3378
2 81654 1 3378
2 81655 1 3378
2 81656 1 3378
2 81657 1 3378
2 81658 1 3378
2 81659 1 3378
2 81660 1 3378
2 81661 1 3379
2 81662 1 3379
2 81663 1 3379
2 81664 1 3379
2 81665 1 3379
2 81666 1 3379
2 81667 1 3379
2 81668 1 3379
2 81669 1 3379
2 81670 1 3379
2 81671 1 3379
2 81672 1 3379
2 81673 1 3379
2 81674 1 3379
2 81675 1 3380
2 81676 1 3380
2 81677 1 3388
2 81678 1 3388
2 81679 1 3388
2 81680 1 3388
2 81681 1 3388
2 81682 1 3388
2 81683 1 3389
2 81684 1 3389
2 81685 1 3390
2 81686 1 3390
2 81687 1 3390
2 81688 1 3391
2 81689 1 3391
2 81690 1 3391
2 81691 1 3391
2 81692 1 3391
2 81693 1 3391
2 81694 1 3391
2 81695 1 3391
2 81696 1 3391
2 81697 1 3391
2 81698 1 3391
2 81699 1 3391
2 81700 1 3391
2 81701 1 3391
2 81702 1 3391
2 81703 1 3391
2 81704 1 3391
2 81705 1 3398
2 81706 1 3398
2 81707 1 3398
2 81708 1 3398
2 81709 1 3398
2 81710 1 3398
2 81711 1 3398
2 81712 1 3398
2 81713 1 3398
2 81714 1 3398
2 81715 1 3398
2 81716 1 3406
2 81717 1 3406
2 81718 1 3409
2 81719 1 3409
2 81720 1 3409
2 81721 1 3409
2 81722 1 3409
2 81723 1 3409
2 81724 1 3409
2 81725 1 3409
2 81726 1 3409
2 81727 1 3409
2 81728 1 3409
2 81729 1 3409
2 81730 1 3409
2 81731 1 3409
2 81732 1 3409
2 81733 1 3409
2 81734 1 3409
2 81735 1 3409
2 81736 1 3409
2 81737 1 3409
2 81738 1 3409
2 81739 1 3409
2 81740 1 3409
2 81741 1 3409
2 81742 1 3409
2 81743 1 3409
2 81744 1 3409
2 81745 1 3409
2 81746 1 3411
2 81747 1 3411
2 81748 1 3412
2 81749 1 3412
2 81750 1 3412
2 81751 1 3412
2 81752 1 3412
2 81753 1 3412
2 81754 1 3412
2 81755 1 3412
2 81756 1 3412
2 81757 1 3412
2 81758 1 3412
2 81759 1 3412
2 81760 1 3412
2 81761 1 3412
2 81762 1 3412
2 81763 1 3412
2 81764 1 3412
2 81765 1 3412
2 81766 1 3412
2 81767 1 3412
2 81768 1 3412
2 81769 1 3412
2 81770 1 3412
2 81771 1 3412
2 81772 1 3412
2 81773 1 3412
2 81774 1 3412
2 81775 1 3412
2 81776 1 3412
2 81777 1 3412
2 81778 1 3412
2 81779 1 3412
2 81780 1 3412
2 81781 1 3412
2 81782 1 3412
2 81783 1 3412
2 81784 1 3413
2 81785 1 3413
2 81786 1 3414
2 81787 1 3414
2 81788 1 3416
2 81789 1 3416
2 81790 1 3416
2 81791 1 3416
2 81792 1 3416
2 81793 1 3416
2 81794 1 3423
2 81795 1 3423
2 81796 1 3423
2 81797 1 3423
2 81798 1 3423
2 81799 1 3424
2 81800 1 3424
2 81801 1 3425
2 81802 1 3425
2 81803 1 3425
2 81804 1 3425
2 81805 1 3425
2 81806 1 3425
2 81807 1 3425
2 81808 1 3425
2 81809 1 3425
2 81810 1 3425
2 81811 1 3425
2 81812 1 3425
2 81813 1 3425
2 81814 1 3425
2 81815 1 3425
2 81816 1 3425
2 81817 1 3425
2 81818 1 3425
2 81819 1 3425
2 81820 1 3425
2 81821 1 3425
2 81822 1 3425
2 81823 1 3425
2 81824 1 3425
2 81825 1 3425
2 81826 1 3425
2 81827 1 3425
2 81828 1 3425
2 81829 1 3425
2 81830 1 3425
2 81831 1 3425
2 81832 1 3425
2 81833 1 3425
2 81834 1 3433
2 81835 1 3433
2 81836 1 3433
2 81837 1 3433
2 81838 1 3433
2 81839 1 3433
2 81840 1 3433
2 81841 1 3433
2 81842 1 3433
2 81843 1 3433
2 81844 1 3433
2 81845 1 3433
2 81846 1 3433
2 81847 1 3433
2 81848 1 3433
2 81849 1 3433
2 81850 1 3433
2 81851 1 3433
2 81852 1 3434
2 81853 1 3434
2 81854 1 3434
2 81855 1 3435
2 81856 1 3435
2 81857 1 3435
2 81858 1 3435
2 81859 1 3435
2 81860 1 3435
2 81861 1 3435
2 81862 1 3441
2 81863 1 3441
2 81864 1 3441
2 81865 1 3441
2 81866 1 3442
2 81867 1 3442
2 81868 1 3443
2 81869 1 3443
2 81870 1 3443
2 81871 1 3443
2 81872 1 3443
2 81873 1 3443
2 81874 1 3443
2 81875 1 3451
2 81876 1 3451
2 81877 1 3451
2 81878 1 3451
2 81879 1 3451
2 81880 1 3451
2 81881 1 3451
2 81882 1 3452
2 81883 1 3452
2 81884 1 3454
2 81885 1 3454
2 81886 1 3455
2 81887 1 3455
2 81888 1 3455
2 81889 1 3455
2 81890 1 3455
2 81891 1 3455
2 81892 1 3455
2 81893 1 3455
2 81894 1 3455
2 81895 1 3455
2 81896 1 3455
2 81897 1 3456
2 81898 1 3456
2 81899 1 3456
2 81900 1 3456
2 81901 1 3456
2 81902 1 3460
2 81903 1 3460
2 81904 1 3469
2 81905 1 3469
2 81906 1 3469
2 81907 1 3469
2 81908 1 3469
2 81909 1 3469
2 81910 1 3469
2 81911 1 3469
2 81912 1 3469
2 81913 1 3469
2 81914 1 3469
2 81915 1 3469
2 81916 1 3469
2 81917 1 3469
2 81918 1 3469
2 81919 1 3469
2 81920 1 3469
2 81921 1 3469
2 81922 1 3469
2 81923 1 3469
2 81924 1 3469
2 81925 1 3469
2 81926 1 3469
2 81927 1 3469
2 81928 1 3469
2 81929 1 3469
2 81930 1 3469
2 81931 1 3469
2 81932 1 3469
2 81933 1 3469
2 81934 1 3469
2 81935 1 3469
2 81936 1 3469
2 81937 1 3469
2 81938 1 3469
2 81939 1 3469
2 81940 1 3469
2 81941 1 3469
2 81942 1 3469
2 81943 1 3469
2 81944 1 3469
2 81945 1 3469
2 81946 1 3469
2 81947 1 3469
2 81948 1 3469
2 81949 1 3469
2 81950 1 3469
2 81951 1 3469
2 81952 1 3469
2 81953 1 3469
2 81954 1 3469
2 81955 1 3469
2 81956 1 3469
2 81957 1 3469
2 81958 1 3469
2 81959 1 3469
2 81960 1 3469
2 81961 1 3469
2 81962 1 3469
2 81963 1 3469
2 81964 1 3469
2 81965 1 3469
2 81966 1 3469
2 81967 1 3469
2 81968 1 3469
2 81969 1 3469
2 81970 1 3469
2 81971 1 3469
2 81972 1 3469
2 81973 1 3470
2 81974 1 3470
2 81975 1 3471
2 81976 1 3471
2 81977 1 3471
2 81978 1 3471
2 81979 1 3471
2 81980 1 3471
2 81981 1 3471
2 81982 1 3471
2 81983 1 3471
2 81984 1 3471
2 81985 1 3471
2 81986 1 3471
2 81987 1 3471
2 81988 1 3471
2 81989 1 3471
2 81990 1 3471
2 81991 1 3471
2 81992 1 3471
2 81993 1 3471
2 81994 1 3471
2 81995 1 3471
2 81996 1 3471
2 81997 1 3471
2 81998 1 3471
2 81999 1 3471
2 82000 1 3471
2 82001 1 3471
2 82002 1 3471
2 82003 1 3471
2 82004 1 3471
2 82005 1 3471
2 82006 1 3471
2 82007 1 3471
2 82008 1 3471
2 82009 1 3471
2 82010 1 3471
2 82011 1 3471
2 82012 1 3471
2 82013 1 3471
2 82014 1 3473
2 82015 1 3473
2 82016 1 3476
2 82017 1 3476
2 82018 1 3476
2 82019 1 3476
2 82020 1 3476
2 82021 1 3476
2 82022 1 3476
2 82023 1 3476
2 82024 1 3476
2 82025 1 3480
2 82026 1 3480
2 82027 1 3480
2 82028 1 3480
2 82029 1 3487
2 82030 1 3487
2 82031 1 3487
2 82032 1 3487
2 82033 1 3489
2 82034 1 3489
2 82035 1 3489
2 82036 1 3489
2 82037 1 3489
2 82038 1 3489
2 82039 1 3489
2 82040 1 3489
2 82041 1 3489
2 82042 1 3490
2 82043 1 3490
2 82044 1 3498
2 82045 1 3498
2 82046 1 3498
2 82047 1 3498
2 82048 1 3498
2 82049 1 3498
2 82050 1 3498
2 82051 1 3498
2 82052 1 3498
2 82053 1 3498
2 82054 1 3498
2 82055 1 3498
2 82056 1 3498
2 82057 1 3498
2 82058 1 3498
2 82059 1 3498
2 82060 1 3499
2 82061 1 3499
2 82062 1 3501
2 82063 1 3501
2 82064 1 3501
2 82065 1 3501
2 82066 1 3501
2 82067 1 3502
2 82068 1 3502
2 82069 1 3511
2 82070 1 3511
2 82071 1 3511
2 82072 1 3511
2 82073 1 3514
2 82074 1 3514
2 82075 1 3514
2 82076 1 3514
2 82077 1 3514
2 82078 1 3514
2 82079 1 3514
2 82080 1 3514
2 82081 1 3514
2 82082 1 3514
2 82083 1 3515
2 82084 1 3515
2 82085 1 3515
2 82086 1 3515
2 82087 1 3523
2 82088 1 3523
2 82089 1 3524
2 82090 1 3524
2 82091 1 3524
2 82092 1 3524
2 82093 1 3524
2 82094 1 3524
2 82095 1 3524
2 82096 1 3524
2 82097 1 3524
2 82098 1 3534
2 82099 1 3534
2 82100 1 3534
2 82101 1 3534
2 82102 1 3534
2 82103 1 3534
2 82104 1 3534
2 82105 1 3534
2 82106 1 3534
2 82107 1 3534
2 82108 1 3534
2 82109 1 3534
2 82110 1 3534
2 82111 1 3534
2 82112 1 3534
2 82113 1 3534
2 82114 1 3534
2 82115 1 3534
2 82116 1 3534
2 82117 1 3534
2 82118 1 3534
2 82119 1 3534
2 82120 1 3534
2 82121 1 3534
2 82122 1 3534
2 82123 1 3534
2 82124 1 3534
2 82125 1 3534
2 82126 1 3535
2 82127 1 3535
2 82128 1 3535
2 82129 1 3535
2 82130 1 3535
2 82131 1 3535
2 82132 1 3535
2 82133 1 3535
2 82134 1 3535
2 82135 1 3535
2 82136 1 3535
2 82137 1 3535
2 82138 1 3535
2 82139 1 3535
2 82140 1 3535
2 82141 1 3535
2 82142 1 3535
2 82143 1 3535
2 82144 1 3535
2 82145 1 3536
2 82146 1 3536
2 82147 1 3537
2 82148 1 3537
2 82149 1 3537
2 82150 1 3537
2 82151 1 3537
2 82152 1 3537
2 82153 1 3537
2 82154 1 3537
2 82155 1 3537
2 82156 1 3537
2 82157 1 3537
2 82158 1 3537
2 82159 1 3537
2 82160 1 3537
2 82161 1 3537
2 82162 1 3538
2 82163 1 3538
2 82164 1 3538
2 82165 1 3538
2 82166 1 3538
2 82167 1 3538
2 82168 1 3538
2 82169 1 3538
2 82170 1 3538
2 82171 1 3538
2 82172 1 3538
2 82173 1 3538
2 82174 1 3538
2 82175 1 3538
2 82176 1 3538
2 82177 1 3538
2 82178 1 3542
2 82179 1 3542
2 82180 1 3542
2 82181 1 3543
2 82182 1 3543
2 82183 1 3543
2 82184 1 3543
2 82185 1 3543
2 82186 1 3543
2 82187 1 3543
2 82188 1 3547
2 82189 1 3547
2 82190 1 3547
2 82191 1 3547
2 82192 1 3547
2 82193 1 3547
2 82194 1 3547
2 82195 1 3547
2 82196 1 3547
2 82197 1 3547
2 82198 1 3547
2 82199 1 3547
2 82200 1 3547
2 82201 1 3547
2 82202 1 3547
2 82203 1 3549
2 82204 1 3549
2 82205 1 3549
2 82206 1 3549
2 82207 1 3549
2 82208 1 3549
2 82209 1 3549
2 82210 1 3549
2 82211 1 3549
2 82212 1 3549
2 82213 1 3549
2 82214 1 3550
2 82215 1 3550
2 82216 1 3562
2 82217 1 3562
2 82218 1 3562
2 82219 1 3562
2 82220 1 3562
2 82221 1 3563
2 82222 1 3563
2 82223 1 3570
2 82224 1 3570
2 82225 1 3571
2 82226 1 3571
2 82227 1 3571
2 82228 1 3571
2 82229 1 3571
2 82230 1 3571
2 82231 1 3571
2 82232 1 3571
2 82233 1 3571
2 82234 1 3571
2 82235 1 3571
2 82236 1 3571
2 82237 1 3571
2 82238 1 3571
2 82239 1 3571
2 82240 1 3571
2 82241 1 3571
2 82242 1 3571
2 82243 1 3571
2 82244 1 3571
2 82245 1 3571
2 82246 1 3572
2 82247 1 3572
2 82248 1 3572
2 82249 1 3572
2 82250 1 3572
2 82251 1 3572
2 82252 1 3573
2 82253 1 3573
2 82254 1 3581
2 82255 1 3581
2 82256 1 3581
2 82257 1 3582
2 82258 1 3582
2 82259 1 3582
2 82260 1 3584
2 82261 1 3584
2 82262 1 3584
2 82263 1 3587
2 82264 1 3587
2 82265 1 3587
2 82266 1 3587
2 82267 1 3587
2 82268 1 3587
2 82269 1 3587
2 82270 1 3592
2 82271 1 3592
2 82272 1 3592
2 82273 1 3592
2 82274 1 3592
2 82275 1 3592
2 82276 1 3592
2 82277 1 3592
2 82278 1 3592
2 82279 1 3592
2 82280 1 3592
2 82281 1 3592
2 82282 1 3592
2 82283 1 3592
2 82284 1 3592
2 82285 1 3592
2 82286 1 3592
2 82287 1 3592
2 82288 1 3592
2 82289 1 3592
2 82290 1 3592
2 82291 1 3592
2 82292 1 3592
2 82293 1 3593
2 82294 1 3593
2 82295 1 3593
2 82296 1 3593
2 82297 1 3593
2 82298 1 3593
2 82299 1 3602
2 82300 1 3602
2 82301 1 3602
2 82302 1 3603
2 82303 1 3603
2 82304 1 3603
2 82305 1 3603
2 82306 1 3603
2 82307 1 3603
2 82308 1 3603
2 82309 1 3603
2 82310 1 3603
2 82311 1 3603
2 82312 1 3604
2 82313 1 3604
2 82314 1 3604
2 82315 1 3604
2 82316 1 3604
2 82317 1 3607
2 82318 1 3607
2 82319 1 3607
2 82320 1 3607
2 82321 1 3607
2 82322 1 3607
2 82323 1 3607
2 82324 1 3607
2 82325 1 3607
2 82326 1 3607
2 82327 1 3607
2 82328 1 3607
2 82329 1 3607
2 82330 1 3607
2 82331 1 3607
2 82332 1 3607
2 82333 1 3607
2 82334 1 3607
2 82335 1 3607
2 82336 1 3607
2 82337 1 3607
2 82338 1 3607
2 82339 1 3607
2 82340 1 3607
2 82341 1 3607
2 82342 1 3607
2 82343 1 3607
2 82344 1 3607
2 82345 1 3607
2 82346 1 3607
2 82347 1 3607
2 82348 1 3607
2 82349 1 3615
2 82350 1 3615
2 82351 1 3615
2 82352 1 3615
2 82353 1 3615
2 82354 1 3616
2 82355 1 3616
2 82356 1 3617
2 82357 1 3617
2 82358 1 3617
2 82359 1 3617
2 82360 1 3617
2 82361 1 3622
2 82362 1 3622
2 82363 1 3622
2 82364 1 3622
2 82365 1 3622
2 82366 1 3622
2 82367 1 3622
2 82368 1 3622
2 82369 1 3622
2 82370 1 3622
2 82371 1 3622
2 82372 1 3622
2 82373 1 3622
2 82374 1 3622
2 82375 1 3622
2 82376 1 3622
2 82377 1 3622
2 82378 1 3622
2 82379 1 3622
2 82380 1 3622
2 82381 1 3622
2 82382 1 3622
2 82383 1 3622
2 82384 1 3622
2 82385 1 3622
2 82386 1 3623
2 82387 1 3623
2 82388 1 3623
2 82389 1 3624
2 82390 1 3624
2 82391 1 3624
2 82392 1 3624
2 82393 1 3624
2 82394 1 3624
2 82395 1 3624
2 82396 1 3624
2 82397 1 3624
2 82398 1 3624
2 82399 1 3625
2 82400 1 3625
2 82401 1 3625
2 82402 1 3625
2 82403 1 3625
2 82404 1 3633
2 82405 1 3633
2 82406 1 3633
2 82407 1 3633
2 82408 1 3633
2 82409 1 3633
2 82410 1 3633
2 82411 1 3633
2 82412 1 3633
2 82413 1 3633
2 82414 1 3633
2 82415 1 3633
2 82416 1 3635
2 82417 1 3635
2 82418 1 3635
2 82419 1 3635
2 82420 1 3635
2 82421 1 3635
2 82422 1 3635
2 82423 1 3635
2 82424 1 3635
2 82425 1 3636
2 82426 1 3636
2 82427 1 3636
2 82428 1 3636
2 82429 1 3636
2 82430 1 3636
2 82431 1 3636
2 82432 1 3637
2 82433 1 3637
2 82434 1 3637
2 82435 1 3637
2 82436 1 3637
2 82437 1 3637
2 82438 1 3637
2 82439 1 3637
2 82440 1 3637
2 82441 1 3637
2 82442 1 3637
2 82443 1 3637
2 82444 1 3637
2 82445 1 3637
2 82446 1 3637
2 82447 1 3637
2 82448 1 3646
2 82449 1 3646
2 82450 1 3646
2 82451 1 3646
2 82452 1 3647
2 82453 1 3647
2 82454 1 3647
2 82455 1 3648
2 82456 1 3648
2 82457 1 3648
2 82458 1 3648
2 82459 1 3648
2 82460 1 3648
2 82461 1 3650
2 82462 1 3650
2 82463 1 3651
2 82464 1 3651
2 82465 1 3651
2 82466 1 3651
2 82467 1 3651
2 82468 1 3651
2 82469 1 3651
2 82470 1 3651
2 82471 1 3651
2 82472 1 3651
2 82473 1 3653
2 82474 1 3653
2 82475 1 3659
2 82476 1 3659
2 82477 1 3659
2 82478 1 3660
2 82479 1 3660
2 82480 1 3667
2 82481 1 3667
2 82482 1 3667
2 82483 1 3667
2 82484 1 3667
2 82485 1 3667
2 82486 1 3669
2 82487 1 3669
2 82488 1 3669
2 82489 1 3669
2 82490 1 3669
2 82491 1 3669
2 82492 1 3670
2 82493 1 3670
2 82494 1 3670
2 82495 1 3673
2 82496 1 3673
2 82497 1 3673
2 82498 1 3673
2 82499 1 3673
2 82500 1 3673
2 82501 1 3673
2 82502 1 3674
2 82503 1 3674
2 82504 1 3674
2 82505 1 3675
2 82506 1 3675
2 82507 1 3682
2 82508 1 3682
2 82509 1 3682
2 82510 1 3682
2 82511 1 3682
2 82512 1 3682
2 82513 1 3682
2 82514 1 3682
2 82515 1 3690
2 82516 1 3690
2 82517 1 3690
2 82518 1 3702
2 82519 1 3702
2 82520 1 3702
2 82521 1 3702
2 82522 1 3702
2 82523 1 3702
2 82524 1 3702
2 82525 1 3702
2 82526 1 3702
2 82527 1 3702
2 82528 1 3702
2 82529 1 3702
2 82530 1 3702
2 82531 1 3703
2 82532 1 3703
2 82533 1 3703
2 82534 1 3704
2 82535 1 3704
2 82536 1 3704
2 82537 1 3704
2 82538 1 3705
2 82539 1 3705
2 82540 1 3705
2 82541 1 3705
2 82542 1 3705
2 82543 1 3705
2 82544 1 3705
2 82545 1 3705
2 82546 1 3705
2 82547 1 3705
2 82548 1 3705
2 82549 1 3705
2 82550 1 3705
2 82551 1 3705
2 82552 1 3705
2 82553 1 3706
2 82554 1 3706
2 82555 1 3706
2 82556 1 3706
2 82557 1 3706
2 82558 1 3707
2 82559 1 3707
2 82560 1 3708
2 82561 1 3708
2 82562 1 3708
2 82563 1 3708
2 82564 1 3708
2 82565 1 3708
2 82566 1 3712
2 82567 1 3712
2 82568 1 3712
2 82569 1 3712
2 82570 1 3715
2 82571 1 3715
2 82572 1 3715
2 82573 1 3715
2 82574 1 3715
2 82575 1 3715
2 82576 1 3715
2 82577 1 3715
2 82578 1 3715
2 82579 1 3715
2 82580 1 3715
2 82581 1 3715
2 82582 1 3715
2 82583 1 3715
2 82584 1 3715
2 82585 1 3715
2 82586 1 3716
2 82587 1 3716
2 82588 1 3717
2 82589 1 3717
2 82590 1 3717
2 82591 1 3717
2 82592 1 3722
2 82593 1 3722
2 82594 1 3722
2 82595 1 3722
2 82596 1 3722
2 82597 1 3722
2 82598 1 3722
2 82599 1 3722
2 82600 1 3722
2 82601 1 3722
2 82602 1 3722
2 82603 1 3722
2 82604 1 3722
2 82605 1 3722
2 82606 1 3722
2 82607 1 3722
2 82608 1 3722
2 82609 1 3722
2 82610 1 3723
2 82611 1 3723
2 82612 1 3723
2 82613 1 3723
2 82614 1 3723
2 82615 1 3723
2 82616 1 3723
2 82617 1 3723
2 82618 1 3723
2 82619 1 3723
2 82620 1 3723
2 82621 1 3723
2 82622 1 3723
2 82623 1 3723
2 82624 1 3723
2 82625 1 3723
2 82626 1 3723
2 82627 1 3723
2 82628 1 3723
2 82629 1 3723
2 82630 1 3723
2 82631 1 3723
2 82632 1 3723
2 82633 1 3723
2 82634 1 3723
2 82635 1 3723
2 82636 1 3723
2 82637 1 3723
2 82638 1 3723
2 82639 1 3724
2 82640 1 3724
2 82641 1 3724
2 82642 1 3732
2 82643 1 3732
2 82644 1 3732
2 82645 1 3732
2 82646 1 3732
2 82647 1 3732
2 82648 1 3732
2 82649 1 3732
2 82650 1 3732
2 82651 1 3734
2 82652 1 3734
2 82653 1 3734
2 82654 1 3734
2 82655 1 3734
2 82656 1 3734
2 82657 1 3734
2 82658 1 3734
2 82659 1 3734
2 82660 1 3734
2 82661 1 3734
2 82662 1 3734
2 82663 1 3734
2 82664 1 3734
2 82665 1 3734
2 82666 1 3734
2 82667 1 3734
2 82668 1 3734
2 82669 1 3734
2 82670 1 3734
2 82671 1 3734
2 82672 1 3734
2 82673 1 3734
2 82674 1 3734
2 82675 1 3734
2 82676 1 3734
2 82677 1 3735
2 82678 1 3735
2 82679 1 3735
2 82680 1 3735
2 82681 1 3735
2 82682 1 3735
2 82683 1 3735
2 82684 1 3735
2 82685 1 3735
2 82686 1 3736
2 82687 1 3736
2 82688 1 3737
2 82689 1 3737
2 82690 1 3738
2 82691 1 3738
2 82692 1 3738
2 82693 1 3738
2 82694 1 3738
2 82695 1 3741
2 82696 1 3741
2 82697 1 3741
2 82698 1 3741
2 82699 1 3741
2 82700 1 3741
2 82701 1 3741
2 82702 1 3741
2 82703 1 3741
2 82704 1 3741
2 82705 1 3741
2 82706 1 3741
2 82707 1 3741
2 82708 1 3741
2 82709 1 3742
2 82710 1 3742
2 82711 1 3743
2 82712 1 3743
2 82713 1 3743
2 82714 1 3743
2 82715 1 3743
2 82716 1 3743
2 82717 1 3743
2 82718 1 3743
2 82719 1 3743
2 82720 1 3744
2 82721 1 3744
2 82722 1 3744
2 82723 1 3744
2 82724 1 3752
2 82725 1 3752
2 82726 1 3752
2 82727 1 3752
2 82728 1 3752
2 82729 1 3752
2 82730 1 3752
2 82731 1 3752
2 82732 1 3752
2 82733 1 3752
2 82734 1 3752
2 82735 1 3752
2 82736 1 3752
2 82737 1 3752
2 82738 1 3752
2 82739 1 3752
2 82740 1 3752
2 82741 1 3752
2 82742 1 3752
2 82743 1 3752
2 82744 1 3752
2 82745 1 3752
2 82746 1 3752
2 82747 1 3752
2 82748 1 3752
2 82749 1 3752
2 82750 1 3752
2 82751 1 3752
2 82752 1 3753
2 82753 1 3753
2 82754 1 3753
2 82755 1 3754
2 82756 1 3754
2 82757 1 3754
2 82758 1 3754
2 82759 1 3754
2 82760 1 3754
2 82761 1 3754
2 82762 1 3754
2 82763 1 3755
2 82764 1 3755
2 82765 1 3755
2 82766 1 3755
2 82767 1 3756
2 82768 1 3756
2 82769 1 3756
2 82770 1 3757
2 82771 1 3757
2 82772 1 3757
2 82773 1 3757
2 82774 1 3757
2 82775 1 3757
2 82776 1 3757
2 82777 1 3757
2 82778 1 3757
2 82779 1 3757
2 82780 1 3757
2 82781 1 3757
2 82782 1 3757
2 82783 1 3757
2 82784 1 3757
2 82785 1 3757
2 82786 1 3757
2 82787 1 3757
2 82788 1 3757
2 82789 1 3757
2 82790 1 3757
2 82791 1 3758
2 82792 1 3758
2 82793 1 3758
2 82794 1 3758
2 82795 1 3758
2 82796 1 3767
2 82797 1 3767
2 82798 1 3767
2 82799 1 3767
2 82800 1 3768
2 82801 1 3768
2 82802 1 3769
2 82803 1 3769
2 82804 1 3769
2 82805 1 3769
2 82806 1 3769
2 82807 1 3769
2 82808 1 3769
2 82809 1 3769
2 82810 1 3769
2 82811 1 3769
2 82812 1 3769
2 82813 1 3769
2 82814 1 3769
2 82815 1 3769
2 82816 1 3769
2 82817 1 3770
2 82818 1 3770
2 82819 1 3770
2 82820 1 3771
2 82821 1 3771
2 82822 1 3771
2 82823 1 3771
2 82824 1 3771
2 82825 1 3771
2 82826 1 3775
2 82827 1 3775
2 82828 1 3777
2 82829 1 3777
2 82830 1 3780
2 82831 1 3780
2 82832 1 3786
2 82833 1 3786
2 82834 1 3786
2 82835 1 3786
2 82836 1 3786
2 82837 1 3786
2 82838 1 3786
2 82839 1 3786
2 82840 1 3786
2 82841 1 3786
2 82842 1 3786
2 82843 1 3786
2 82844 1 3786
2 82845 1 3786
2 82846 1 3786
2 82847 1 3786
2 82848 1 3786
2 82849 1 3786
2 82850 1 3786
2 82851 1 3786
2 82852 1 3786
2 82853 1 3786
2 82854 1 3786
2 82855 1 3786
2 82856 1 3786
2 82857 1 3786
2 82858 1 3786
2 82859 1 3787
2 82860 1 3787
2 82861 1 3787
2 82862 1 3787
2 82863 1 3787
2 82864 1 3787
2 82865 1 3787
2 82866 1 3795
2 82867 1 3795
2 82868 1 3795
2 82869 1 3795
2 82870 1 3795
2 82871 1 3795
2 82872 1 3795
2 82873 1 3795
2 82874 1 3798
2 82875 1 3798
2 82876 1 3798
2 82877 1 3798
2 82878 1 3798
2 82879 1 3798
2 82880 1 3798
2 82881 1 3798
2 82882 1 3798
2 82883 1 3798
2 82884 1 3798
2 82885 1 3799
2 82886 1 3799
2 82887 1 3800
2 82888 1 3800
2 82889 1 3800
2 82890 1 3800
2 82891 1 3800
2 82892 1 3800
2 82893 1 3801
2 82894 1 3801
2 82895 1 3801
2 82896 1 3801
2 82897 1 3801
2 82898 1 3801
2 82899 1 3801
2 82900 1 3806
2 82901 1 3806
2 82902 1 3806
2 82903 1 3806
2 82904 1 3806
2 82905 1 3806
2 82906 1 3806
2 82907 1 3807
2 82908 1 3807
2 82909 1 3817
2 82910 1 3817
2 82911 1 3817
2 82912 1 3817
2 82913 1 3817
2 82914 1 3817
2 82915 1 3817
2 82916 1 3817
2 82917 1 3818
2 82918 1 3818
2 82919 1 3818
2 82920 1 3818
2 82921 1 3818
2 82922 1 3818
2 82923 1 3818
2 82924 1 3818
2 82925 1 3819
2 82926 1 3819
2 82927 1 3820
2 82928 1 3820
2 82929 1 3820
2 82930 1 3820
2 82931 1 3821
2 82932 1 3821
2 82933 1 3821
2 82934 1 3836
2 82935 1 3836
2 82936 1 3836
2 82937 1 3836
2 82938 1 3836
2 82939 1 3836
2 82940 1 3836
2 82941 1 3836
2 82942 1 3838
2 82943 1 3838
2 82944 1 3839
2 82945 1 3839
2 82946 1 3839
2 82947 1 3839
2 82948 1 3843
2 82949 1 3843
2 82950 1 3843
2 82951 1 3843
2 82952 1 3843
2 82953 1 3844
2 82954 1 3844
2 82955 1 3850
2 82956 1 3850
2 82957 1 3856
2 82958 1 3856
2 82959 1 3856
2 82960 1 3864
2 82961 1 3864
2 82962 1 3864
2 82963 1 3864
2 82964 1 3864
2 82965 1 3864
2 82966 1 3864
2 82967 1 3864
2 82968 1 3864
2 82969 1 3864
2 82970 1 3864
2 82971 1 3864
2 82972 1 3866
2 82973 1 3866
2 82974 1 3866
2 82975 1 3866
2 82976 1 3866
2 82977 1 3870
2 82978 1 3870
2 82979 1 3871
2 82980 1 3871
2 82981 1 3872
2 82982 1 3872
2 82983 1 3872
2 82984 1 3872
2 82985 1 3872
2 82986 1 3872
2 82987 1 3872
2 82988 1 3872
2 82989 1 3872
2 82990 1 3872
2 82991 1 3872
2 82992 1 3872
2 82993 1 3872
2 82994 1 3872
2 82995 1 3872
2 82996 1 3872
2 82997 1 3872
2 82998 1 3872
2 82999 1 3872
2 83000 1 3873
2 83001 1 3873
2 83002 1 3873
2 83003 1 3882
2 83004 1 3882
2 83005 1 3884
2 83006 1 3884
2 83007 1 3884
2 83008 1 3884
2 83009 1 3884
2 83010 1 3884
2 83011 1 3884
2 83012 1 3884
2 83013 1 3885
2 83014 1 3885
2 83015 1 3888
2 83016 1 3888
2 83017 1 3888
2 83018 1 3889
2 83019 1 3889
2 83020 1 3898
2 83021 1 3898
2 83022 1 3899
2 83023 1 3899
2 83024 1 3899
2 83025 1 3902
2 83026 1 3902
2 83027 1 3902
2 83028 1 3902
2 83029 1 3902
2 83030 1 3902
2 83031 1 3902
2 83032 1 3902
2 83033 1 3902
2 83034 1 3902
2 83035 1 3902
2 83036 1 3902
2 83037 1 3902
2 83038 1 3902
2 83039 1 3902
2 83040 1 3902
2 83041 1 3902
2 83042 1 3902
2 83043 1 3902
2 83044 1 3902
2 83045 1 3902
2 83046 1 3902
2 83047 1 3902
2 83048 1 3902
2 83049 1 3902
2 83050 1 3902
2 83051 1 3902
2 83052 1 3902
2 83053 1 3902
2 83054 1 3902
2 83055 1 3902
2 83056 1 3902
2 83057 1 3902
2 83058 1 3902
2 83059 1 3902
2 83060 1 3902
2 83061 1 3902
2 83062 1 3902
2 83063 1 3902
2 83064 1 3902
2 83065 1 3902
2 83066 1 3902
2 83067 1 3902
2 83068 1 3902
2 83069 1 3902
2 83070 1 3902
2 83071 1 3904
2 83072 1 3904
2 83073 1 3904
2 83074 1 3905
2 83075 1 3905
2 83076 1 3905
2 83077 1 3905
2 83078 1 3905
2 83079 1 3905
2 83080 1 3905
2 83081 1 3905
2 83082 1 3905
2 83083 1 3905
2 83084 1 3905
2 83085 1 3905
2 83086 1 3905
2 83087 1 3905
2 83088 1 3905
2 83089 1 3905
2 83090 1 3905
2 83091 1 3905
2 83092 1 3905
2 83093 1 3905
2 83094 1 3905
2 83095 1 3905
2 83096 1 3905
2 83097 1 3905
2 83098 1 3905
2 83099 1 3905
2 83100 1 3905
2 83101 1 3905
2 83102 1 3905
2 83103 1 3905
2 83104 1 3905
2 83105 1 3905
2 83106 1 3905
2 83107 1 3905
2 83108 1 3905
2 83109 1 3905
2 83110 1 3905
2 83111 1 3905
2 83112 1 3905
2 83113 1 3905
2 83114 1 3905
2 83115 1 3905
2 83116 1 3905
2 83117 1 3905
2 83118 1 3905
2 83119 1 3905
2 83120 1 3905
2 83121 1 3905
2 83122 1 3905
2 83123 1 3905
2 83124 1 3905
2 83125 1 3905
2 83126 1 3905
2 83127 1 3905
2 83128 1 3905
2 83129 1 3905
2 83130 1 3905
2 83131 1 3905
2 83132 1 3905
2 83133 1 3905
2 83134 1 3905
2 83135 1 3905
2 83136 1 3905
2 83137 1 3905
2 83138 1 3905
2 83139 1 3905
2 83140 1 3905
2 83141 1 3905
2 83142 1 3905
2 83143 1 3905
2 83144 1 3905
2 83145 1 3905
2 83146 1 3905
2 83147 1 3905
2 83148 1 3905
2 83149 1 3905
2 83150 1 3905
2 83151 1 3905
2 83152 1 3905
2 83153 1 3905
2 83154 1 3905
2 83155 1 3905
2 83156 1 3905
2 83157 1 3905
2 83158 1 3905
2 83159 1 3905
2 83160 1 3905
2 83161 1 3905
2 83162 1 3905
2 83163 1 3905
2 83164 1 3905
2 83165 1 3905
2 83166 1 3905
2 83167 1 3905
2 83168 1 3905
2 83169 1 3905
2 83170 1 3906
2 83171 1 3906
2 83172 1 3906
2 83173 1 3906
2 83174 1 3906
2 83175 1 3906
2 83176 1 3906
2 83177 1 3906
2 83178 1 3913
2 83179 1 3913
2 83180 1 3925
2 83181 1 3925
2 83182 1 3925
2 83183 1 3925
2 83184 1 3925
2 83185 1 3928
2 83186 1 3928
2 83187 1 3928
2 83188 1 3928
2 83189 1 3928
2 83190 1 3929
2 83191 1 3929
2 83192 1 3929
2 83193 1 3930
2 83194 1 3930
2 83195 1 3930
2 83196 1 3930
2 83197 1 3944
2 83198 1 3944
2 83199 1 3944
2 83200 1 3944
2 83201 1 3945
2 83202 1 3945
2 83203 1 3945
2 83204 1 3945
2 83205 1 3945
2 83206 1 3945
2 83207 1 3945
2 83208 1 3945
2 83209 1 3945
2 83210 1 3945
2 83211 1 3945
2 83212 1 3945
2 83213 1 3945
2 83214 1 3945
2 83215 1 3945
2 83216 1 3945
2 83217 1 3947
2 83218 1 3947
2 83219 1 3947
2 83220 1 3947
2 83221 1 3947
2 83222 1 3947
2 83223 1 3947
2 83224 1 3947
2 83225 1 3947
2 83226 1 3947
2 83227 1 3947
2 83228 1 3947
2 83229 1 3948
2 83230 1 3948
2 83231 1 3949
2 83232 1 3949
2 83233 1 3949
2 83234 1 3949
2 83235 1 3952
2 83236 1 3952
2 83237 1 3956
2 83238 1 3956
2 83239 1 3961
2 83240 1 3961
2 83241 1 3961
2 83242 1 3963
2 83243 1 3963
2 83244 1 3968
2 83245 1 3968
2 83246 1 3968
2 83247 1 3968
2 83248 1 3968
2 83249 1 3969
2 83250 1 3969
2 83251 1 3969
2 83252 1 3977
2 83253 1 3977
2 83254 1 3980
2 83255 1 3980
2 83256 1 3982
2 83257 1 3982
2 83258 1 3983
2 83259 1 3983
2 83260 1 3983
2 83261 1 3983
2 83262 1 3987
2 83263 1 3987
2 83264 1 3987
2 83265 1 3988
2 83266 1 3988
2 83267 1 3988
2 83268 1 3988
2 83269 1 3988
2 83270 1 3988
2 83271 1 3988
2 83272 1 3989
2 83273 1 3989
2 83274 1 3997
2 83275 1 3997
2 83276 1 3997
2 83277 1 4000
2 83278 1 4000
2 83279 1 4000
2 83280 1 4000
2 83281 1 4000
2 83282 1 4000
2 83283 1 4000
2 83284 1 4000
2 83285 1 4000
2 83286 1 4000
2 83287 1 4000
2 83288 1 4000
2 83289 1 4000
2 83290 1 4000
2 83291 1 4000
2 83292 1 4000
2 83293 1 4000
2 83294 1 4000
2 83295 1 4000
2 83296 1 4001
2 83297 1 4001
2 83298 1 4001
2 83299 1 4001
2 83300 1 4001
2 83301 1 4009
2 83302 1 4009
2 83303 1 4009
2 83304 1 4009
2 83305 1 4009
2 83306 1 4009
2 83307 1 4009
2 83308 1 4010
2 83309 1 4010
2 83310 1 4010
2 83311 1 4011
2 83312 1 4011
2 83313 1 4013
2 83314 1 4013
2 83315 1 4013
2 83316 1 4013
2 83317 1 4013
2 83318 1 4014
2 83319 1 4014
2 83320 1 4016
2 83321 1 4016
2 83322 1 4016
2 83323 1 4016
2 83324 1 4019
2 83325 1 4019
2 83326 1 4019
2 83327 1 4019
2 83328 1 4019
2 83329 1 4019
2 83330 1 4019
2 83331 1 4019
2 83332 1 4019
2 83333 1 4019
2 83334 1 4019
2 83335 1 4019
2 83336 1 4019
2 83337 1 4019
2 83338 1 4019
2 83339 1 4019
2 83340 1 4019
2 83341 1 4019
2 83342 1 4019
2 83343 1 4019
2 83344 1 4019
2 83345 1 4019
2 83346 1 4019
2 83347 1 4021
2 83348 1 4021
2 83349 1 4021
2 83350 1 4021
2 83351 1 4021
2 83352 1 4021
2 83353 1 4021
2 83354 1 4021
2 83355 1 4021
2 83356 1 4021
2 83357 1 4021
2 83358 1 4021
2 83359 1 4021
2 83360 1 4021
2 83361 1 4021
2 83362 1 4021
2 83363 1 4033
2 83364 1 4033
2 83365 1 4033
2 83366 1 4033
2 83367 1 4033
2 83368 1 4034
2 83369 1 4034
2 83370 1 4034
2 83371 1 4034
2 83372 1 4034
2 83373 1 4034
2 83374 1 4042
2 83375 1 4042
2 83376 1 4042
2 83377 1 4042
2 83378 1 4042
2 83379 1 4042
2 83380 1 4042
2 83381 1 4042
2 83382 1 4042
2 83383 1 4042
2 83384 1 4042
2 83385 1 4042
2 83386 1 4042
2 83387 1 4042
2 83388 1 4042
2 83389 1 4042
2 83390 1 4044
2 83391 1 4044
2 83392 1 4044
2 83393 1 4044
2 83394 1 4044
2 83395 1 4044
2 83396 1 4044
2 83397 1 4044
2 83398 1 4044
2 83399 1 4045
2 83400 1 4045
2 83401 1 4054
2 83402 1 4054
2 83403 1 4054
2 83404 1 4054
2 83405 1 4054
2 83406 1 4054
2 83407 1 4054
2 83408 1 4054
2 83409 1 4054
2 83410 1 4054
2 83411 1 4054
2 83412 1 4054
2 83413 1 4054
2 83414 1 4054
2 83415 1 4054
2 83416 1 4054
2 83417 1 4054
2 83418 1 4054
2 83419 1 4054
2 83420 1 4054
2 83421 1 4054
2 83422 1 4054
2 83423 1 4054
2 83424 1 4054
2 83425 1 4054
2 83426 1 4055
2 83427 1 4055
2 83428 1 4056
2 83429 1 4056
2 83430 1 4070
2 83431 1 4070
2 83432 1 4070
2 83433 1 4070
2 83434 1 4073
2 83435 1 4073
2 83436 1 4073
2 83437 1 4073
2 83438 1 4073
2 83439 1 4073
2 83440 1 4073
2 83441 1 4077
2 83442 1 4077
2 83443 1 4080
2 83444 1 4080
2 83445 1 4091
2 83446 1 4091
2 83447 1 4092
2 83448 1 4092
2 83449 1 4092
2 83450 1 4093
2 83451 1 4093
2 83452 1 4093
2 83453 1 4093
2 83454 1 4093
2 83455 1 4093
2 83456 1 4093
2 83457 1 4093
2 83458 1 4093
2 83459 1 4093
2 83460 1 4100
2 83461 1 4100
2 83462 1 4108
2 83463 1 4108
2 83464 1 4108
2 83465 1 4108
2 83466 1 4108
2 83467 1 4108
2 83468 1 4108
2 83469 1 4109
2 83470 1 4109
2 83471 1 4109
2 83472 1 4109
2 83473 1 4109
2 83474 1 4109
2 83475 1 4110
2 83476 1 4110
2 83477 1 4111
2 83478 1 4111
2 83479 1 4114
2 83480 1 4114
2 83481 1 4117
2 83482 1 4117
2 83483 1 4123
2 83484 1 4123
2 83485 1 4123
2 83486 1 4123
2 83487 1 4124
2 83488 1 4124
2 83489 1 4132
2 83490 1 4132
2 83491 1 4132
2 83492 1 4141
2 83493 1 4141
2 83494 1 4141
2 83495 1 4141
2 83496 1 4141
2 83497 1 4141
2 83498 1 4141
2 83499 1 4141
2 83500 1 4141
2 83501 1 4142
2 83502 1 4142
2 83503 1 4142
2 83504 1 4143
2 83505 1 4143
2 83506 1 4143
2 83507 1 4150
2 83508 1 4150
2 83509 1 4150
2 83510 1 4150
2 83511 1 4150
2 83512 1 4152
2 83513 1 4152
2 83514 1 4152
2 83515 1 4155
2 83516 1 4155
2 83517 1 4155
2 83518 1 4155
2 83519 1 4155
2 83520 1 4155
2 83521 1 4155
2 83522 1 4155
2 83523 1 4155
2 83524 1 4155
2 83525 1 4155
2 83526 1 4156
2 83527 1 4156
2 83528 1 4167
2 83529 1 4167
2 83530 1 4167
2 83531 1 4167
2 83532 1 4167
2 83533 1 4167
2 83534 1 4167
2 83535 1 4168
2 83536 1 4168
2 83537 1 4168
2 83538 1 4168
2 83539 1 4168
2 83540 1 4168
2 83541 1 4168
2 83542 1 4168
2 83543 1 4168
2 83544 1 4168
2 83545 1 4168
2 83546 1 4168
2 83547 1 4168
2 83548 1 4168
2 83549 1 4168
2 83550 1 4168
2 83551 1 4168
2 83552 1 4168
2 83553 1 4177
2 83554 1 4177
2 83555 1 4177
2 83556 1 4177
2 83557 1 4177
2 83558 1 4177
2 83559 1 4177
2 83560 1 4177
2 83561 1 4178
2 83562 1 4178
2 83563 1 4186
2 83564 1 4186
2 83565 1 4186
2 83566 1 4186
2 83567 1 4186
2 83568 1 4186
2 83569 1 4186
2 83570 1 4187
2 83571 1 4187
2 83572 1 4187
2 83573 1 4188
2 83574 1 4188
2 83575 1 4189
2 83576 1 4189
2 83577 1 4189
2 83578 1 4189
2 83579 1 4189
2 83580 1 4189
2 83581 1 4189
2 83582 1 4189
2 83583 1 4189
2 83584 1 4189
2 83585 1 4189
2 83586 1 4189
2 83587 1 4189
2 83588 1 4189
2 83589 1 4189
2 83590 1 4189
2 83591 1 4189
2 83592 1 4189
2 83593 1 4189
2 83594 1 4189
2 83595 1 4189
2 83596 1 4189
2 83597 1 4189
2 83598 1 4189
2 83599 1 4189
2 83600 1 4189
2 83601 1 4189
2 83602 1 4190
2 83603 1 4190
2 83604 1 4203
2 83605 1 4203
2 83606 1 4203
2 83607 1 4203
2 83608 1 4204
2 83609 1 4204
2 83610 1 4204
2 83611 1 4204
2 83612 1 4205
2 83613 1 4205
2 83614 1 4205
2 83615 1 4205
2 83616 1 4205
2 83617 1 4205
2 83618 1 4205
2 83619 1 4205
2 83620 1 4205
2 83621 1 4206
2 83622 1 4206
2 83623 1 4206
2 83624 1 4209
2 83625 1 4209
2 83626 1 4209
2 83627 1 4209
2 83628 1 4209
2 83629 1 4209
2 83630 1 4209
2 83631 1 4209
2 83632 1 4209
2 83633 1 4209
2 83634 1 4209
2 83635 1 4209
2 83636 1 4210
2 83637 1 4210
2 83638 1 4211
2 83639 1 4211
2 83640 1 4212
2 83641 1 4212
2 83642 1 4212
2 83643 1 4213
2 83644 1 4213
2 83645 1 4213
2 83646 1 4213
2 83647 1 4213
2 83648 1 4213
2 83649 1 4213
2 83650 1 4213
2 83651 1 4213
2 83652 1 4213
2 83653 1 4213
2 83654 1 4217
2 83655 1 4217
2 83656 1 4217
2 83657 1 4217
2 83658 1 4220
2 83659 1 4220
2 83660 1 4220
2 83661 1 4220
2 83662 1 4220
2 83663 1 4221
2 83664 1 4221
2 83665 1 4221
2 83666 1 4221
2 83667 1 4221
2 83668 1 4228
2 83669 1 4228
2 83670 1 4229
2 83671 1 4229
2 83672 1 4229
2 83673 1 4229
2 83674 1 4229
2 83675 1 4229
2 83676 1 4229
2 83677 1 4229
2 83678 1 4229
2 83679 1 4229
2 83680 1 4229
2 83681 1 4229
2 83682 1 4229
2 83683 1 4230
2 83684 1 4230
2 83685 1 4238
2 83686 1 4238
2 83687 1 4238
2 83688 1 4238
2 83689 1 4238
2 83690 1 4238
2 83691 1 4238
2 83692 1 4238
2 83693 1 4238
2 83694 1 4238
2 83695 1 4239
2 83696 1 4239
2 83697 1 4242
2 83698 1 4242
2 83699 1 4242
2 83700 1 4243
2 83701 1 4243
2 83702 1 4243
2 83703 1 4253
2 83704 1 4253
2 83705 1 4253
2 83706 1 4253
2 83707 1 4253
2 83708 1 4253
2 83709 1 4253
2 83710 1 4261
2 83711 1 4261
2 83712 1 4262
2 83713 1 4262
2 83714 1 4262
2 83715 1 4262
2 83716 1 4262
2 83717 1 4262
2 83718 1 4262
2 83719 1 4262
2 83720 1 4263
2 83721 1 4263
2 83722 1 4263
2 83723 1 4263
2 83724 1 4264
2 83725 1 4264
2 83726 1 4267
2 83727 1 4267
2 83728 1 4267
2 83729 1 4267
2 83730 1 4267
2 83731 1 4267
2 83732 1 4268
2 83733 1 4268
2 83734 1 4268
2 83735 1 4268
2 83736 1 4268
2 83737 1 4268
2 83738 1 4268
2 83739 1 4268
2 83740 1 4268
2 83741 1 4268
2 83742 1 4268
2 83743 1 4268
2 83744 1 4268
2 83745 1 4268
2 83746 1 4269
2 83747 1 4269
2 83748 1 4276
2 83749 1 4276
2 83750 1 4276
2 83751 1 4285
2 83752 1 4285
2 83753 1 4285
2 83754 1 4285
2 83755 1 4285
2 83756 1 4285
2 83757 1 4285
2 83758 1 4285
2 83759 1 4285
2 83760 1 4285
2 83761 1 4285
2 83762 1 4285
2 83763 1 4286
2 83764 1 4286
2 83765 1 4287
2 83766 1 4287
2 83767 1 4287
2 83768 1 4287
2 83769 1 4287
2 83770 1 4287
2 83771 1 4288
2 83772 1 4288
2 83773 1 4289
2 83774 1 4289
2 83775 1 4297
2 83776 1 4297
2 83777 1 4298
2 83778 1 4298
2 83779 1 4300
2 83780 1 4300
2 83781 1 4300
2 83782 1 4300
2 83783 1 4300
2 83784 1 4300
2 83785 1 4300
2 83786 1 4301
2 83787 1 4301
2 83788 1 4308
2 83789 1 4308
2 83790 1 4316
2 83791 1 4316
2 83792 1 4316
2 83793 1 4316
2 83794 1 4316
2 83795 1 4316
2 83796 1 4316
2 83797 1 4316
2 83798 1 4316
2 83799 1 4316
2 83800 1 4316
2 83801 1 4316
2 83802 1 4316
2 83803 1 4316
2 83804 1 4316
2 83805 1 4316
2 83806 1 4316
2 83807 1 4316
2 83808 1 4316
2 83809 1 4316
2 83810 1 4316
2 83811 1 4316
2 83812 1 4316
2 83813 1 4316
2 83814 1 4316
2 83815 1 4316
2 83816 1 4316
2 83817 1 4316
2 83818 1 4316
2 83819 1 4316
2 83820 1 4316
2 83821 1 4316
2 83822 1 4316
2 83823 1 4316
2 83824 1 4316
2 83825 1 4316
2 83826 1 4317
2 83827 1 4317
2 83828 1 4317
2 83829 1 4317
2 83830 1 4317
2 83831 1 4317
2 83832 1 4317
2 83833 1 4317
2 83834 1 4317
2 83835 1 4317
2 83836 1 4317
2 83837 1 4317
2 83838 1 4317
2 83839 1 4318
2 83840 1 4318
2 83841 1 4318
2 83842 1 4319
2 83843 1 4319
2 83844 1 4319
2 83845 1 4319
2 83846 1 4319
2 83847 1 4322
2 83848 1 4322
2 83849 1 4322
2 83850 1 4322
2 83851 1 4322
2 83852 1 4326
2 83853 1 4326
2 83854 1 4341
2 83855 1 4341
2 83856 1 4341
2 83857 1 4344
2 83858 1 4344
2 83859 1 4345
2 83860 1 4345
2 83861 1 4345
2 83862 1 4345
2 83863 1 4345
2 83864 1 4345
2 83865 1 4345
2 83866 1 4345
2 83867 1 4345
2 83868 1 4346
2 83869 1 4346
2 83870 1 4346
2 83871 1 4346
2 83872 1 4347
2 83873 1 4347
2 83874 1 4355
2 83875 1 4355
2 83876 1 4355
2 83877 1 4355
2 83878 1 4355
2 83879 1 4355
2 83880 1 4356
2 83881 1 4356
2 83882 1 4359
2 83883 1 4359
2 83884 1 4359
2 83885 1 4367
2 83886 1 4367
2 83887 1 4367
2 83888 1 4367
2 83889 1 4367
2 83890 1 4367
2 83891 1 4367
2 83892 1 4367
2 83893 1 4367
2 83894 1 4368
2 83895 1 4368
2 83896 1 4368
2 83897 1 4376
2 83898 1 4376
2 83899 1 4376
2 83900 1 4376
2 83901 1 4376
2 83902 1 4376
2 83903 1 4376
2 83904 1 4376
2 83905 1 4376
2 83906 1 4376
2 83907 1 4376
2 83908 1 4376
2 83909 1 4378
2 83910 1 4378
2 83911 1 4378
2 83912 1 4378
2 83913 1 4378
2 83914 1 4378
2 83915 1 4379
2 83916 1 4379
2 83917 1 4379
2 83918 1 4379
2 83919 1 4379
2 83920 1 4379
2 83921 1 4381
2 83922 1 4381
2 83923 1 4381
2 83924 1 4381
2 83925 1 4381
2 83926 1 4381
2 83927 1 4381
2 83928 1 4381
2 83929 1 4381
2 83930 1 4382
2 83931 1 4382
2 83932 1 4384
2 83933 1 4384
2 83934 1 4392
2 83935 1 4392
2 83936 1 4400
2 83937 1 4400
2 83938 1 4400
2 83939 1 4400
2 83940 1 4400
2 83941 1 4401
2 83942 1 4401
2 83943 1 4409
2 83944 1 4409
2 83945 1 4413
2 83946 1 4413
2 83947 1 4413
2 83948 1 4413
2 83949 1 4413
2 83950 1 4413
2 83951 1 4413
2 83952 1 4413
2 83953 1 4413
2 83954 1 4413
2 83955 1 4413
2 83956 1 4413
2 83957 1 4413
2 83958 1 4413
2 83959 1 4413
2 83960 1 4413
2 83961 1 4413
2 83962 1 4413
2 83963 1 4413
2 83964 1 4413
2 83965 1 4413
2 83966 1 4413
2 83967 1 4413
2 83968 1 4413
2 83969 1 4413
2 83970 1 4413
2 83971 1 4413
2 83972 1 4413
2 83973 1 4414
2 83974 1 4414
2 83975 1 4414
2 83976 1 4421
2 83977 1 4421
2 83978 1 4422
2 83979 1 4422
2 83980 1 4432
2 83981 1 4432
2 83982 1 4432
2 83983 1 4432
2 83984 1 4432
2 83985 1 4432
2 83986 1 4432
2 83987 1 4432
2 83988 1 4432
2 83989 1 4432
2 83990 1 4433
2 83991 1 4433
2 83992 1 4433
2 83993 1 4450
2 83994 1 4450
2 83995 1 4450
2 83996 1 4450
2 83997 1 4450
2 83998 1 4450
2 83999 1 4450
2 84000 1 4450
2 84001 1 4450
2 84002 1 4451
2 84003 1 4451
2 84004 1 4451
2 84005 1 4451
2 84006 1 4451
2 84007 1 4451
2 84008 1 4451
2 84009 1 4451
2 84010 1 4451
2 84011 1 4451
2 84012 1 4451
2 84013 1 4451
2 84014 1 4451
2 84015 1 4451
2 84016 1 4451
2 84017 1 4451
2 84018 1 4451
2 84019 1 4451
2 84020 1 4451
2 84021 1 4451
2 84022 1 4451
2 84023 1 4451
2 84024 1 4451
2 84025 1 4451
2 84026 1 4452
2 84027 1 4452
2 84028 1 4453
2 84029 1 4453
2 84030 1 4453
2 84031 1 4453
2 84032 1 4454
2 84033 1 4454
2 84034 1 4454
2 84035 1 4454
2 84036 1 4454
2 84037 1 4454
2 84038 1 4454
2 84039 1 4454
2 84040 1 4454
2 84041 1 4456
2 84042 1 4456
2 84043 1 4456
2 84044 1 4457
2 84045 1 4457
2 84046 1 4465
2 84047 1 4465
2 84048 1 4465
2 84049 1 4465
2 84050 1 4465
2 84051 1 4465
2 84052 1 4466
2 84053 1 4466
2 84054 1 4466
2 84055 1 4466
2 84056 1 4466
2 84057 1 4466
2 84058 1 4466
2 84059 1 4466
2 84060 1 4466
2 84061 1 4466
2 84062 1 4467
2 84063 1 4467
2 84064 1 4467
2 84065 1 4470
2 84066 1 4470
2 84067 1 4470
2 84068 1 4470
2 84069 1 4470
2 84070 1 4470
2 84071 1 4470
2 84072 1 4470
2 84073 1 4470
2 84074 1 4470
2 84075 1 4470
2 84076 1 4470
2 84077 1 4470
2 84078 1 4470
2 84079 1 4470
2 84080 1 4470
2 84081 1 4470
2 84082 1 4470
2 84083 1 4470
2 84084 1 4470
2 84085 1 4470
2 84086 1 4471
2 84087 1 4471
2 84088 1 4471
2 84089 1 4471
2 84090 1 4471
2 84091 1 4471
2 84092 1 4471
2 84093 1 4471
2 84094 1 4471
2 84095 1 4471
2 84096 1 4478
2 84097 1 4478
2 84098 1 4478
2 84099 1 4491
2 84100 1 4491
2 84101 1 4491
2 84102 1 4491
2 84103 1 4491
2 84104 1 4491
2 84105 1 4491
2 84106 1 4491
2 84107 1 4491
2 84108 1 4493
2 84109 1 4493
2 84110 1 4511
2 84111 1 4511
2 84112 1 4511
2 84113 1 4529
2 84114 1 4529
2 84115 1 4529
2 84116 1 4529
2 84117 1 4529
2 84118 1 4530
2 84119 1 4530
2 84120 1 4530
2 84121 1 4530
2 84122 1 4530
2 84123 1 4530
2 84124 1 4530
2 84125 1 4530
2 84126 1 4530
2 84127 1 4530
2 84128 1 4530
2 84129 1 4530
2 84130 1 4530
2 84131 1 4530
2 84132 1 4532
2 84133 1 4532
2 84134 1 4532
2 84135 1 4533
2 84136 1 4533
2 84137 1 4533
2 84138 1 4534
2 84139 1 4534
2 84140 1 4539
2 84141 1 4539
2 84142 1 4543
2 84143 1 4543
2 84144 1 4543
2 84145 1 4543
2 84146 1 4543
2 84147 1 4543
2 84148 1 4543
2 84149 1 4543
2 84150 1 4543
2 84151 1 4543
2 84152 1 4543
2 84153 1 4544
2 84154 1 4544
2 84155 1 4546
2 84156 1 4546
2 84157 1 4546
2 84158 1 4546
2 84159 1 4546
2 84160 1 4546
2 84161 1 4546
2 84162 1 4546
2 84163 1 4546
2 84164 1 4546
2 84165 1 4546
2 84166 1 4546
2 84167 1 4546
2 84168 1 4546
2 84169 1 4547
2 84170 1 4547
2 84171 1 4547
2 84172 1 4547
2 84173 1 4547
2 84174 1 4548
2 84175 1 4548
2 84176 1 4548
2 84177 1 4548
2 84178 1 4548
2 84179 1 4556
2 84180 1 4556
2 84181 1 4557
2 84182 1 4557
2 84183 1 4557
2 84184 1 4557
2 84185 1 4557
2 84186 1 4557
2 84187 1 4558
2 84188 1 4558
2 84189 1 4558
2 84190 1 4558
2 84191 1 4558
2 84192 1 4572
2 84193 1 4572
2 84194 1 4572
2 84195 1 4572
2 84196 1 4572
2 84197 1 4572
2 84198 1 4572
2 84199 1 4572
2 84200 1 4572
2 84201 1 4574
2 84202 1 4574
2 84203 1 4574
2 84204 1 4575
2 84205 1 4575
2 84206 1 4581
2 84207 1 4581
2 84208 1 4581
2 84209 1 4581
2 84210 1 4581
2 84211 1 4581
2 84212 1 4581
2 84213 1 4581
2 84214 1 4582
2 84215 1 4582
2 84216 1 4582
2 84217 1 4582
2 84218 1 4582
2 84219 1 4590
2 84220 1 4590
2 84221 1 4590
2 84222 1 4593
2 84223 1 4593
2 84224 1 4593
2 84225 1 4593
2 84226 1 4593
2 84227 1 4593
2 84228 1 4593
2 84229 1 4593
2 84230 1 4593
2 84231 1 4593
2 84232 1 4593
2 84233 1 4593
2 84234 1 4595
2 84235 1 4595
2 84236 1 4595
2 84237 1 4598
2 84238 1 4598
2 84239 1 4598
2 84240 1 4598
2 84241 1 4598
2 84242 1 4603
2 84243 1 4603
2 84244 1 4603
2 84245 1 4603
2 84246 1 4603
2 84247 1 4603
2 84248 1 4603
2 84249 1 4604
2 84250 1 4604
2 84251 1 4604
2 84252 1 4604
2 84253 1 4604
2 84254 1 4604
2 84255 1 4605
2 84256 1 4605
2 84257 1 4605
2 84258 1 4605
2 84259 1 4605
2 84260 1 4605
2 84261 1 4605
2 84262 1 4616
2 84263 1 4616
2 84264 1 4616
2 84265 1 4616
2 84266 1 4616
2 84267 1 4616
2 84268 1 4617
2 84269 1 4617
2 84270 1 4617
2 84271 1 4618
2 84272 1 4618
2 84273 1 4619
2 84274 1 4619
2 84275 1 4619
2 84276 1 4619
2 84277 1 4619
2 84278 1 4619
2 84279 1 4619
2 84280 1 4619
2 84281 1 4619
2 84282 1 4620
2 84283 1 4620
2 84284 1 4621
2 84285 1 4621
2 84286 1 4621
2 84287 1 4621
2 84288 1 4621
2 84289 1 4630
2 84290 1 4630
2 84291 1 4630
2 84292 1 4630
2 84293 1 4630
2 84294 1 4631
2 84295 1 4631
2 84296 1 4631
2 84297 1 4632
2 84298 1 4632
2 84299 1 4632
2 84300 1 4632
2 84301 1 4632
2 84302 1 4632
2 84303 1 4632
2 84304 1 4632
2 84305 1 4632
2 84306 1 4632
2 84307 1 4632
2 84308 1 4632
2 84309 1 4633
2 84310 1 4633
2 84311 1 4633
2 84312 1 4633
2 84313 1 4633
2 84314 1 4633
2 84315 1 4633
2 84316 1 4633
2 84317 1 4633
2 84318 1 4633
2 84319 1 4633
2 84320 1 4633
2 84321 1 4633
2 84322 1 4633
2 84323 1 4633
2 84324 1 4633
2 84325 1 4633
2 84326 1 4633
2 84327 1 4636
2 84328 1 4636
2 84329 1 4637
2 84330 1 4637
2 84331 1 4637
2 84332 1 4637
2 84333 1 4637
2 84334 1 4637
2 84335 1 4637
2 84336 1 4637
2 84337 1 4637
2 84338 1 4637
2 84339 1 4637
2 84340 1 4644
2 84341 1 4644
2 84342 1 4644
2 84343 1 4644
2 84344 1 4644
2 84345 1 4644
2 84346 1 4646
2 84347 1 4646
2 84348 1 4647
2 84349 1 4647
2 84350 1 4654
2 84351 1 4654
2 84352 1 4654
2 84353 1 4654
2 84354 1 4662
2 84355 1 4662
2 84356 1 4662
2 84357 1 4662
2 84358 1 4662
2 84359 1 4662
2 84360 1 4662
2 84361 1 4662
2 84362 1 4662
2 84363 1 4662
2 84364 1 4662
2 84365 1 4662
2 84366 1 4662
2 84367 1 4662
2 84368 1 4662
2 84369 1 4662
2 84370 1 4662
2 84371 1 4662
2 84372 1 4663
2 84373 1 4663
2 84374 1 4663
2 84375 1 4663
2 84376 1 4664
2 84377 1 4664
2 84378 1 4664
2 84379 1 4664
2 84380 1 4664
2 84381 1 4664
2 84382 1 4664
2 84383 1 4664
2 84384 1 4664
2 84385 1 4664
2 84386 1 4664
2 84387 1 4664
2 84388 1 4664
2 84389 1 4664
2 84390 1 4664
2 84391 1 4664
2 84392 1 4665
2 84393 1 4665
2 84394 1 4665
2 84395 1 4665
2 84396 1 4665
2 84397 1 4665
2 84398 1 4673
2 84399 1 4673
2 84400 1 4673
2 84401 1 4673
2 84402 1 4673
2 84403 1 4673
2 84404 1 4673
2 84405 1 4673
2 84406 1 4673
2 84407 1 4673
2 84408 1 4673
2 84409 1 4673
2 84410 1 4673
2 84411 1 4673
2 84412 1 4673
2 84413 1 4673
2 84414 1 4673
2 84415 1 4673
2 84416 1 4673
2 84417 1 4673
2 84418 1 4673
2 84419 1 4673
2 84420 1 4673
2 84421 1 4676
2 84422 1 4676
2 84423 1 4676
2 84424 1 4676
2 84425 1 4676
2 84426 1 4676
2 84427 1 4676
2 84428 1 4676
2 84429 1 4677
2 84430 1 4677
2 84431 1 4677
2 84432 1 4677
2 84433 1 4677
2 84434 1 4677
2 84435 1 4677
2 84436 1 4677
2 84437 1 4677
2 84438 1 4677
2 84439 1 4677
2 84440 1 4677
2 84441 1 4690
2 84442 1 4690
2 84443 1 4690
2 84444 1 4690
2 84445 1 4690
2 84446 1 4690
2 84447 1 4690
2 84448 1 4690
2 84449 1 4690
2 84450 1 4690
2 84451 1 4690
2 84452 1 4690
2 84453 1 4691
2 84454 1 4691
2 84455 1 4691
2 84456 1 4691
2 84457 1 4691
2 84458 1 4691
2 84459 1 4692
2 84460 1 4692
2 84461 1 4700
2 84462 1 4700
2 84463 1 4700
2 84464 1 4700
2 84465 1 4700
2 84466 1 4700
2 84467 1 4700
2 84468 1 4700
2 84469 1 4700
2 84470 1 4701
2 84471 1 4701
2 84472 1 4701
2 84473 1 4701
2 84474 1 4701
2 84475 1 4701
2 84476 1 4701
2 84477 1 4704
2 84478 1 4704
2 84479 1 4704
2 84480 1 4704
2 84481 1 4704
2 84482 1 4704
2 84483 1 4704
2 84484 1 4704
2 84485 1 4704
2 84486 1 4704
2 84487 1 4704
2 84488 1 4704
2 84489 1 4704
2 84490 1 4704
2 84491 1 4706
2 84492 1 4706
2 84493 1 4711
2 84494 1 4711
2 84495 1 4711
2 84496 1 4711
2 84497 1 4711
2 84498 1 4711
2 84499 1 4711
2 84500 1 4711
2 84501 1 4711
2 84502 1 4711
2 84503 1 4711
2 84504 1 4711
2 84505 1 4712
2 84506 1 4712
2 84507 1 4712
2 84508 1 4721
2 84509 1 4721
2 84510 1 4721
2 84511 1 4721
2 84512 1 4721
2 84513 1 4721
2 84514 1 4721
2 84515 1 4721
2 84516 1 4721
2 84517 1 4722
2 84518 1 4722
2 84519 1 4723
2 84520 1 4723
2 84521 1 4723
2 84522 1 4723
2 84523 1 4723
2 84524 1 4723
2 84525 1 4723
2 84526 1 4723
2 84527 1 4723
2 84528 1 4723
2 84529 1 4723
2 84530 1 4723
2 84531 1 4723
2 84532 1 4725
2 84533 1 4725
2 84534 1 4725
2 84535 1 4725
2 84536 1 4733
2 84537 1 4733
2 84538 1 4733
2 84539 1 4734
2 84540 1 4734
2 84541 1 4735
2 84542 1 4735
2 84543 1 4735
2 84544 1 4735
2 84545 1 4735
2 84546 1 4748
2 84547 1 4748
2 84548 1 4748
2 84549 1 4749
2 84550 1 4749
2 84551 1 4749
2 84552 1 4752
2 84553 1 4752
2 84554 1 4758
2 84555 1 4758
2 84556 1 4758
2 84557 1 4758
2 84558 1 4758
2 84559 1 4758
2 84560 1 4758
2 84561 1 4758
2 84562 1 4758
2 84563 1 4758
2 84564 1 4759
2 84565 1 4759
2 84566 1 4759
2 84567 1 4759
2 84568 1 4759
2 84569 1 4759
2 84570 1 4759
2 84571 1 4759
2 84572 1 4759
2 84573 1 4760
2 84574 1 4760
2 84575 1 4760
2 84576 1 4760
2 84577 1 4760
2 84578 1 4760
2 84579 1 4760
2 84580 1 4761
2 84581 1 4761
2 84582 1 4761
2 84583 1 4761
2 84584 1 4766
2 84585 1 4766
2 84586 1 4766
2 84587 1 4766
2 84588 1 4766
2 84589 1 4766
2 84590 1 4766
2 84591 1 4766
2 84592 1 4766
2 84593 1 4766
2 84594 1 4766
2 84595 1 4767
2 84596 1 4767
2 84597 1 4767
2 84598 1 4767
2 84599 1 4767
2 84600 1 4767
2 84601 1 4767
2 84602 1 4767
2 84603 1 4767
2 84604 1 4767
2 84605 1 4767
2 84606 1 4767
2 84607 1 4767
2 84608 1 4767
2 84609 1 4767
2 84610 1 4768
2 84611 1 4768
2 84612 1 4770
2 84613 1 4770
2 84614 1 4770
2 84615 1 4771
2 84616 1 4771
2 84617 1 4771
2 84618 1 4771
2 84619 1 4771
2 84620 1 4771
2 84621 1 4771
2 84622 1 4771
2 84623 1 4773
2 84624 1 4773
2 84625 1 4773
2 84626 1 4787
2 84627 1 4787
2 84628 1 4803
2 84629 1 4803
2 84630 1 4803
2 84631 1 4803
2 84632 1 4803
2 84633 1 4808
2 84634 1 4808
2 84635 1 4808
2 84636 1 4811
2 84637 1 4811
2 84638 1 4811
2 84639 1 4812
2 84640 1 4812
2 84641 1 4812
2 84642 1 4812
2 84643 1 4812
2 84644 1 4812
2 84645 1 4812
2 84646 1 4817
2 84647 1 4817
2 84648 1 4817
2 84649 1 4817
2 84650 1 4817
2 84651 1 4817
2 84652 1 4817
2 84653 1 4817
2 84654 1 4817
2 84655 1 4817
2 84656 1 4817
2 84657 1 4817
2 84658 1 4817
2 84659 1 4817
2 84660 1 4817
2 84661 1 4817
2 84662 1 4817
2 84663 1 4817
2 84664 1 4817
2 84665 1 4817
2 84666 1 4817
2 84667 1 4818
2 84668 1 4818
2 84669 1 4818
2 84670 1 4818
2 84671 1 4818
2 84672 1 4818
2 84673 1 4818
2 84674 1 4818
2 84675 1 4818
2 84676 1 4819
2 84677 1 4819
2 84678 1 4821
2 84679 1 4821
2 84680 1 4822
2 84681 1 4822
2 84682 1 4822
2 84683 1 4822
2 84684 1 4822
2 84685 1 4822
2 84686 1 4837
2 84687 1 4837
2 84688 1 4837
2 84689 1 4837
2 84690 1 4838
2 84691 1 4838
2 84692 1 4840
2 84693 1 4840
2 84694 1 4843
2 84695 1 4843
2 84696 1 4843
2 84697 1 4844
2 84698 1 4844
2 84699 1 4847
2 84700 1 4847
2 84701 1 4856
2 84702 1 4856
2 84703 1 4856
2 84704 1 4856
2 84705 1 4856
2 84706 1 4857
2 84707 1 4857
2 84708 1 4858
2 84709 1 4858
2 84710 1 4858
2 84711 1 4858
2 84712 1 4858
2 84713 1 4858
2 84714 1 4858
2 84715 1 4858
2 84716 1 4860
2 84717 1 4860
2 84718 1 4860
2 84719 1 4860
2 84720 1 4861
2 84721 1 4861
2 84722 1 4864
2 84723 1 4864
2 84724 1 4866
2 84725 1 4866
2 84726 1 4867
2 84727 1 4867
2 84728 1 4870
2 84729 1 4870
2 84730 1 4872
2 84731 1 4872
2 84732 1 4872
2 84733 1 4872
2 84734 1 4874
2 84735 1 4874
2 84736 1 4875
2 84737 1 4875
2 84738 1 4875
2 84739 1 4875
2 84740 1 4875
2 84741 1 4875
2 84742 1 4876
2 84743 1 4876
2 84744 1 4876
2 84745 1 4880
2 84746 1 4880
2 84747 1 4880
2 84748 1 4880
2 84749 1 4887
2 84750 1 4887
2 84751 1 4889
2 84752 1 4889
2 84753 1 4889
2 84754 1 4889
2 84755 1 4889
2 84756 1 4889
2 84757 1 4896
2 84758 1 4896
2 84759 1 4896
2 84760 1 4896
2 84761 1 4897
2 84762 1 4897
2 84763 1 4897
2 84764 1 4897
2 84765 1 4897
2 84766 1 4897
2 84767 1 4897
2 84768 1 4897
2 84769 1 4898
2 84770 1 4898
2 84771 1 4901
2 84772 1 4901
2 84773 1 4915
2 84774 1 4915
2 84775 1 4916
2 84776 1 4916
2 84777 1 4920
2 84778 1 4920
2 84779 1 4920
2 84780 1 4920
2 84781 1 4920
2 84782 1 4920
2 84783 1 4920
2 84784 1 4920
2 84785 1 4920
2 84786 1 4920
2 84787 1 4920
2 84788 1 4920
2 84789 1 4920
2 84790 1 4920
2 84791 1 4920
2 84792 1 4920
2 84793 1 4920
2 84794 1 4920
2 84795 1 4920
2 84796 1 4920
2 84797 1 4920
2 84798 1 4920
2 84799 1 4920
2 84800 1 4920
2 84801 1 4920
2 84802 1 4920
2 84803 1 4920
2 84804 1 4920
2 84805 1 4921
2 84806 1 4921
2 84807 1 4922
2 84808 1 4922
2 84809 1 4922
2 84810 1 4922
2 84811 1 4922
2 84812 1 4923
2 84813 1 4923
2 84814 1 4930
2 84815 1 4930
2 84816 1 4930
2 84817 1 4930
2 84818 1 4930
2 84819 1 4930
2 84820 1 4930
2 84821 1 4931
2 84822 1 4931
2 84823 1 4931
2 84824 1 4931
2 84825 1 4942
2 84826 1 4942
2 84827 1 4942
2 84828 1 4942
2 84829 1 4942
2 84830 1 4943
2 84831 1 4943
2 84832 1 4943
2 84833 1 4946
2 84834 1 4946
2 84835 1 4946
2 84836 1 4946
2 84837 1 4955
2 84838 1 4955
2 84839 1 4955
2 84840 1 4955
2 84841 1 4956
2 84842 1 4956
2 84843 1 4956
2 84844 1 4956
2 84845 1 4957
2 84846 1 4957
2 84847 1 4960
2 84848 1 4960
2 84849 1 4960
2 84850 1 4960
2 84851 1 4960
2 84852 1 4960
2 84853 1 4961
2 84854 1 4961
2 84855 1 4968
2 84856 1 4968
2 84857 1 4968
2 84858 1 4968
2 84859 1 4968
2 84860 1 4968
2 84861 1 4968
2 84862 1 4968
2 84863 1 4968
2 84864 1 4968
2 84865 1 4968
2 84866 1 4968
2 84867 1 4968
2 84868 1 4979
2 84869 1 4979
2 84870 1 4979
2 84871 1 4979
2 84872 1 4981
2 84873 1 4981
2 84874 1 4981
2 84875 1 4990
2 84876 1 4990
2 84877 1 4990
2 84878 1 4991
2 84879 1 4991
2 84880 1 4991
2 84881 1 4999
2 84882 1 4999
2 84883 1 4999
2 84884 1 4999
2 84885 1 4999
2 84886 1 5000
2 84887 1 5000
2 84888 1 5000
2 84889 1 5000
2 84890 1 5000
2 84891 1 5000
2 84892 1 5000
2 84893 1 5013
2 84894 1 5013
2 84895 1 5013
2 84896 1 5013
2 84897 1 5014
2 84898 1 5014
2 84899 1 5015
2 84900 1 5015
2 84901 1 5016
2 84902 1 5016
2 84903 1 5016
2 84904 1 5016
2 84905 1 5016
2 84906 1 5016
2 84907 1 5016
2 84908 1 5016
2 84909 1 5017
2 84910 1 5017
2 84911 1 5017
2 84912 1 5018
2 84913 1 5018
2 84914 1 5018
2 84915 1 5025
2 84916 1 5025
2 84917 1 5025
2 84918 1 5027
2 84919 1 5027
2 84920 1 5027
2 84921 1 5027
2 84922 1 5027
2 84923 1 5027
2 84924 1 5027
2 84925 1 5027
2 84926 1 5028
2 84927 1 5028
2 84928 1 5028
2 84929 1 5028
2 84930 1 5035
2 84931 1 5035
2 84932 1 5035
2 84933 1 5036
2 84934 1 5036
2 84935 1 5036
2 84936 1 5043
2 84937 1 5043
2 84938 1 5043
2 84939 1 5046
2 84940 1 5046
2 84941 1 5047
2 84942 1 5047
2 84943 1 5047
2 84944 1 5047
2 84945 1 5047
2 84946 1 5047
2 84947 1 5047
2 84948 1 5047
2 84949 1 5047
2 84950 1 5056
2 84951 1 5056
2 84952 1 5056
2 84953 1 5056
2 84954 1 5057
2 84955 1 5057
2 84956 1 5057
2 84957 1 5058
2 84958 1 5058
2 84959 1 5059
2 84960 1 5059
2 84961 1 5059
2 84962 1 5059
2 84963 1 5059
2 84964 1 5060
2 84965 1 5060
2 84966 1 5065
2 84967 1 5065
2 84968 1 5065
2 84969 1 5065
2 84970 1 5065
2 84971 1 5068
2 84972 1 5068
2 84973 1 5068
2 84974 1 5068
2 84975 1 5070
2 84976 1 5070
2 84977 1 5070
2 84978 1 5070
2 84979 1 5070
2 84980 1 5072
2 84981 1 5072
2 84982 1 5072
2 84983 1 5073
2 84984 1 5073
2 84985 1 5073
2 84986 1 5073
2 84987 1 5073
2 84988 1 5073
2 84989 1 5073
2 84990 1 5073
2 84991 1 5073
2 84992 1 5096
2 84993 1 5096
2 84994 1 5096
2 84995 1 5096
2 84996 1 5098
2 84997 1 5098
2 84998 1 5098
2 84999 1 5098
2 85000 1 5098
2 85001 1 5099
2 85002 1 5099
2 85003 1 5099
2 85004 1 5099
2 85005 1 5099
2 85006 1 5124
2 85007 1 5124
2 85008 1 5124
2 85009 1 5124
2 85010 1 5124
2 85011 1 5124
2 85012 1 5124
2 85013 1 5124
2 85014 1 5124
2 85015 1 5124
2 85016 1 5126
2 85017 1 5126
2 85018 1 5126
2 85019 1 5129
2 85020 1 5129
2 85021 1 5129
2 85022 1 5129
2 85023 1 5129
2 85024 1 5130
2 85025 1 5130
2 85026 1 5130
2 85027 1 5130
2 85028 1 5130
2 85029 1 5130
2 85030 1 5130
2 85031 1 5130
2 85032 1 5130
2 85033 1 5130
2 85034 1 5130
2 85035 1 5131
2 85036 1 5131
2 85037 1 5131
2 85038 1 5141
2 85039 1 5141
2 85040 1 5142
2 85041 1 5142
2 85042 1 5144
2 85043 1 5144
2 85044 1 5149
2 85045 1 5149
2 85046 1 5157
2 85047 1 5157
2 85048 1 5167
2 85049 1 5167
2 85050 1 5167
2 85051 1 5167
2 85052 1 5167
2 85053 1 5167
2 85054 1 5167
2 85055 1 5168
2 85056 1 5168
2 85057 1 5169
2 85058 1 5169
2 85059 1 5169
2 85060 1 5172
2 85061 1 5172
2 85062 1 5172
2 85063 1 5172
2 85064 1 5172
2 85065 1 5179
2 85066 1 5179
2 85067 1 5179
2 85068 1 5179
2 85069 1 5179
2 85070 1 5179
2 85071 1 5179
2 85072 1 5179
2 85073 1 5179
2 85074 1 5179
2 85075 1 5179
2 85076 1 5179
2 85077 1 5179
2 85078 1 5179
2 85079 1 5180
2 85080 1 5180
2 85081 1 5180
2 85082 1 5180
2 85083 1 5180
2 85084 1 5180
2 85085 1 5180
2 85086 1 5180
2 85087 1 5180
2 85088 1 5180
2 85089 1 5181
2 85090 1 5181
2 85091 1 5189
2 85092 1 5189
2 85093 1 5190
2 85094 1 5190
2 85095 1 5190
2 85096 1 5190
2 85097 1 5202
2 85098 1 5202
2 85099 1 5202
2 85100 1 5202
2 85101 1 5202
2 85102 1 5202
2 85103 1 5202
2 85104 1 5202
2 85105 1 5202
2 85106 1 5202
2 85107 1 5202
2 85108 1 5212
2 85109 1 5212
2 85110 1 5212
2 85111 1 5213
2 85112 1 5213
2 85113 1 5230
2 85114 1 5230
2 85115 1 5231
2 85116 1 5231
2 85117 1 5231
2 85118 1 5232
2 85119 1 5232
2 85120 1 5232
2 85121 1 5232
2 85122 1 5232
2 85123 1 5232
2 85124 1 5232
2 85125 1 5232
2 85126 1 5232
2 85127 1 5232
2 85128 1 5232
2 85129 1 5232
2 85130 1 5232
2 85131 1 5232
2 85132 1 5233
2 85133 1 5233
2 85134 1 5233
2 85135 1 5233
2 85136 1 5233
2 85137 1 5233
2 85138 1 5234
2 85139 1 5234
2 85140 1 5234
2 85141 1 5234
2 85142 1 5244
2 85143 1 5244
2 85144 1 5244
2 85145 1 5245
2 85146 1 5245
2 85147 1 5245
2 85148 1 5245
2 85149 1 5245
2 85150 1 5247
2 85151 1 5247
2 85152 1 5250
2 85153 1 5250
2 85154 1 5254
2 85155 1 5254
2 85156 1 5255
2 85157 1 5255
2 85158 1 5255
2 85159 1 5255
2 85160 1 5255
2 85161 1 5256
2 85162 1 5256
2 85163 1 5256
2 85164 1 5258
2 85165 1 5258
2 85166 1 5259
2 85167 1 5259
2 85168 1 5262
2 85169 1 5262
2 85170 1 5262
2 85171 1 5264
2 85172 1 5264
2 85173 1 5264
2 85174 1 5264
2 85175 1 5264
2 85176 1 5272
2 85177 1 5272
2 85178 1 5272
2 85179 1 5274
2 85180 1 5274
2 85181 1 5276
2 85182 1 5276
2 85183 1 5276
2 85184 1 5276
2 85185 1 5276
2 85186 1 5276
2 85187 1 5276
2 85188 1 5276
2 85189 1 5276
2 85190 1 5276
2 85191 1 5276
2 85192 1 5276
2 85193 1 5276
2 85194 1 5277
2 85195 1 5277
2 85196 1 5278
2 85197 1 5278
2 85198 1 5278
2 85199 1 5278
2 85200 1 5291
2 85201 1 5291
2 85202 1 5291
2 85203 1 5293
2 85204 1 5293
2 85205 1 5293
2 85206 1 5293
2 85207 1 5298
2 85208 1 5298
2 85209 1 5298
2 85210 1 5298
2 85211 1 5301
2 85212 1 5301
2 85213 1 5301
2 85214 1 5301
2 85215 1 5301
2 85216 1 5301
2 85217 1 5302
2 85218 1 5302
2 85219 1 5302
2 85220 1 5302
2 85221 1 5302
2 85222 1 5304
2 85223 1 5304
2 85224 1 5307
2 85225 1 5307
2 85226 1 5307
2 85227 1 5308
2 85228 1 5308
2 85229 1 5308
2 85230 1 5320
2 85231 1 5320
2 85232 1 5320
2 85233 1 5321
2 85234 1 5321
2 85235 1 5321
2 85236 1 5321
2 85237 1 5325
2 85238 1 5325
2 85239 1 5330
2 85240 1 5330
2 85241 1 5330
2 85242 1 5330
2 85243 1 5330
2 85244 1 5331
2 85245 1 5331
2 85246 1 5331
2 85247 1 5331
2 85248 1 5331
2 85249 1 5331
2 85250 1 5331
2 85251 1 5331
2 85252 1 5331
2 85253 1 5331
2 85254 1 5331
2 85255 1 5332
2 85256 1 5332
2 85257 1 5332
2 85258 1 5332
2 85259 1 5332
2 85260 1 5334
2 85261 1 5334
2 85262 1 5334
2 85263 1 5334
2 85264 1 5334
2 85265 1 5334
2 85266 1 5334
2 85267 1 5334
2 85268 1 5334
2 85269 1 5334
2 85270 1 5342
2 85271 1 5342
2 85272 1 5342
2 85273 1 5343
2 85274 1 5343
2 85275 1 5348
2 85276 1 5348
2 85277 1 5348
2 85278 1 5348
2 85279 1 5355
2 85280 1 5355
2 85281 1 5355
2 85282 1 5355
2 85283 1 5355
2 85284 1 5356
2 85285 1 5356
2 85286 1 5356
2 85287 1 5356
2 85288 1 5356
2 85289 1 5356
2 85290 1 5357
2 85291 1 5357
2 85292 1 5357
2 85293 1 5358
2 85294 1 5358
2 85295 1 5358
2 85296 1 5359
2 85297 1 5359
2 85298 1 5370
2 85299 1 5370
2 85300 1 5373
2 85301 1 5373
2 85302 1 5374
2 85303 1 5374
2 85304 1 5382
2 85305 1 5382
2 85306 1 5382
2 85307 1 5383
2 85308 1 5383
2 85309 1 5383
2 85310 1 5383
2 85311 1 5384
2 85312 1 5384
2 85313 1 5386
2 85314 1 5386
2 85315 1 5386
2 85316 1 5394
2 85317 1 5394
2 85318 1 5394
2 85319 1 5394
2 85320 1 5394
2 85321 1 5402
2 85322 1 5402
2 85323 1 5402
2 85324 1 5402
2 85325 1 5402
2 85326 1 5402
2 85327 1 5402
2 85328 1 5402
2 85329 1 5403
2 85330 1 5403
2 85331 1 5403
2 85332 1 5403
2 85333 1 5403
2 85334 1 5403
2 85335 1 5403
2 85336 1 5403
2 85337 1 5406
2 85338 1 5406
2 85339 1 5406
2 85340 1 5406
2 85341 1 5407
2 85342 1 5407
2 85343 1 5408
2 85344 1 5408
2 85345 1 5409
2 85346 1 5409
2 85347 1 5409
2 85348 1 5411
2 85349 1 5411
2 85350 1 5418
2 85351 1 5418
2 85352 1 5418
2 85353 1 5418
2 85354 1 5418
2 85355 1 5418
2 85356 1 5418
2 85357 1 5418
2 85358 1 5418
2 85359 1 5418
2 85360 1 5418
2 85361 1 5420
2 85362 1 5420
2 85363 1 5420
2 85364 1 5420
2 85365 1 5420
2 85366 1 5421
2 85367 1 5421
2 85368 1 5430
2 85369 1 5430
2 85370 1 5431
2 85371 1 5431
2 85372 1 5433
2 85373 1 5433
2 85374 1 5439
2 85375 1 5439
2 85376 1 5440
2 85377 1 5440
2 85378 1 5440
2 85379 1 5440
2 85380 1 5440
2 85381 1 5440
2 85382 1 5440
2 85383 1 5440
2 85384 1 5440
2 85385 1 5440
2 85386 1 5441
2 85387 1 5441
2 85388 1 5441
2 85389 1 5457
2 85390 1 5457
2 85391 1 5457
2 85392 1 5470
2 85393 1 5470
2 85394 1 5470
2 85395 1 5470
2 85396 1 5471
2 85397 1 5471
2 85398 1 5471
2 85399 1 5472
2 85400 1 5472
2 85401 1 5472
2 85402 1 5478
2 85403 1 5478
2 85404 1 5478
2 85405 1 5478
2 85406 1 5478
2 85407 1 5478
2 85408 1 5478
2 85409 1 5478
2 85410 1 5494
2 85411 1 5494
2 85412 1 5494
2 85413 1 5494
2 85414 1 5494
2 85415 1 5494
2 85416 1 5494
2 85417 1 5494
2 85418 1 5494
2 85419 1 5494
2 85420 1 5494
2 85421 1 5494
2 85422 1 5494
2 85423 1 5494
2 85424 1 5494
2 85425 1 5494
2 85426 1 5494
2 85427 1 5496
2 85428 1 5496
2 85429 1 5496
2 85430 1 5496
2 85431 1 5496
2 85432 1 5496
2 85433 1 5513
2 85434 1 5513
2 85435 1 5521
2 85436 1 5521
2 85437 1 5536
2 85438 1 5536
2 85439 1 5543
2 85440 1 5543
2 85441 1 5543
2 85442 1 5543
2 85443 1 5544
2 85444 1 5544
2 85445 1 5544
2 85446 1 5557
2 85447 1 5557
2 85448 1 5557
2 85449 1 5557
2 85450 1 5558
2 85451 1 5558
2 85452 1 5558
2 85453 1 5558
2 85454 1 5559
2 85455 1 5559
2 85456 1 5559
2 85457 1 5559
2 85458 1 5560
2 85459 1 5560
2 85460 1 5561
2 85461 1 5561
2 85462 1 5564
2 85463 1 5564
2 85464 1 5564
2 85465 1 5564
2 85466 1 5571
2 85467 1 5571
2 85468 1 5577
2 85469 1 5577
2 85470 1 5577
2 85471 1 5577
2 85472 1 5577
2 85473 1 5577
2 85474 1 5577
2 85475 1 5577
2 85476 1 5577
2 85477 1 5577
2 85478 1 5577
2 85479 1 5577
2 85480 1 5579
2 85481 1 5579
2 85482 1 5591
2 85483 1 5591
2 85484 1 5591
2 85485 1 5593
2 85486 1 5593
2 85487 1 5615
2 85488 1 5615
2 85489 1 5615
2 85490 1 5615
2 85491 1 5615
2 85492 1 5615
2 85493 1 5623
2 85494 1 5623
2 85495 1 5623
2 85496 1 5623
2 85497 1 5623
2 85498 1 5623
2 85499 1 5632
2 85500 1 5632
2 85501 1 5632
2 85502 1 5632
2 85503 1 5632
2 85504 1 5635
2 85505 1 5635
2 85506 1 5635
2 85507 1 5643
2 85508 1 5643
2 85509 1 5643
2 85510 1 5656
2 85511 1 5656
2 85512 1 5656
2 85513 1 5659
2 85514 1 5659
2 85515 1 5659
2 85516 1 5659
2 85517 1 5659
2 85518 1 5659
2 85519 1 5662
2 85520 1 5662
2 85521 1 5662
2 85522 1 5665
2 85523 1 5665
2 85524 1 5666
2 85525 1 5666
2 85526 1 5666
2 85527 1 5666
2 85528 1 5666
2 85529 1 5667
2 85530 1 5667
2 85531 1 5680
2 85532 1 5680
2 85533 1 5680
2 85534 1 5680
2 85535 1 5680
2 85536 1 5683
2 85537 1 5683
2 85538 1 5683
2 85539 1 5697
2 85540 1 5697
2 85541 1 5704
2 85542 1 5704
2 85543 1 5704
2 85544 1 5704
2 85545 1 5704
2 85546 1 5704
2 85547 1 5705
2 85548 1 5705
2 85549 1 5705
2 85550 1 5705
2 85551 1 5705
2 85552 1 5705
2 85553 1 5706
2 85554 1 5706
2 85555 1 5706
2 85556 1 5706
2 85557 1 5706
2 85558 1 5706
2 85559 1 5707
2 85560 1 5707
2 85561 1 5707
2 85562 1 5707
2 85563 1 5707
2 85564 1 5707
2 85565 1 5707
2 85566 1 5707
2 85567 1 5707
2 85568 1 5707
2 85569 1 5707
2 85570 1 5707
2 85571 1 5707
2 85572 1 5707
2 85573 1 5707
2 85574 1 5707
2 85575 1 5707
2 85576 1 5707
2 85577 1 5714
2 85578 1 5714
2 85579 1 5714
2 85580 1 5716
2 85581 1 5716
2 85582 1 5716
2 85583 1 5716
2 85584 1 5716
2 85585 1 5716
2 85586 1 5716
2 85587 1 5716
2 85588 1 5717
2 85589 1 5717
2 85590 1 5717
2 85591 1 5717
2 85592 1 5717
2 85593 1 5717
2 85594 1 5721
2 85595 1 5721
2 85596 1 5729
2 85597 1 5729
2 85598 1 5729
2 85599 1 5738
2 85600 1 5738
2 85601 1 5738
2 85602 1 5739
2 85603 1 5739
2 85604 1 5739
2 85605 1 5739
2 85606 1 5740
2 85607 1 5740
2 85608 1 5742
2 85609 1 5742
2 85610 1 5753
2 85611 1 5753
2 85612 1 5754
2 85613 1 5754
2 85614 1 5754
2 85615 1 5754
2 85616 1 5755
2 85617 1 5755
2 85618 1 5756
2 85619 1 5756
2 85620 1 5764
2 85621 1 5764
2 85622 1 5765
2 85623 1 5765
2 85624 1 5766
2 85625 1 5766
2 85626 1 5767
2 85627 1 5767
2 85628 1 5770
2 85629 1 5770
2 85630 1 5770
2 85631 1 5770
2 85632 1 5770
2 85633 1 5771
2 85634 1 5771
2 85635 1 5782
2 85636 1 5782
2 85637 1 5782
2 85638 1 5782
2 85639 1 5782
2 85640 1 5782
2 85641 1 5782
2 85642 1 5782
2 85643 1 5782
2 85644 1 5782
2 85645 1 5782
2 85646 1 5782
2 85647 1 5782
2 85648 1 5783
2 85649 1 5783
2 85650 1 5783
2 85651 1 5792
2 85652 1 5792
2 85653 1 5792
2 85654 1 5792
2 85655 1 5792
2 85656 1 5792
2 85657 1 5792
2 85658 1 5793
2 85659 1 5793
2 85660 1 5793
2 85661 1 5793
2 85662 1 5796
2 85663 1 5796
2 85664 1 5796
2 85665 1 5796
2 85666 1 5796
2 85667 1 5797
2 85668 1 5797
2 85669 1 5797
2 85670 1 5805
2 85671 1 5805
2 85672 1 5806
2 85673 1 5806
2 85674 1 5813
2 85675 1 5813
2 85676 1 5813
2 85677 1 5816
2 85678 1 5816
2 85679 1 5824
2 85680 1 5824
2 85681 1 5824
2 85682 1 5824
2 85683 1 5824
2 85684 1 5824
2 85685 1 5824
2 85686 1 5824
2 85687 1 5825
2 85688 1 5825
2 85689 1 5826
2 85690 1 5826
2 85691 1 5826
2 85692 1 5826
2 85693 1 5827
2 85694 1 5827
2 85695 1 5828
2 85696 1 5828
2 85697 1 5829
2 85698 1 5829
2 85699 1 5829
2 85700 1 5829
2 85701 1 5829
2 85702 1 5832
2 85703 1 5832
2 85704 1 5832
2 85705 1 5832
2 85706 1 5832
2 85707 1 5832
2 85708 1 5832
2 85709 1 5832
2 85710 1 5832
2 85711 1 5832
2 85712 1 5832
2 85713 1 5832
2 85714 1 5832
2 85715 1 5832
2 85716 1 5834
2 85717 1 5834
2 85718 1 5835
2 85719 1 5835
2 85720 1 5845
2 85721 1 5845
2 85722 1 5845
2 85723 1 5845
2 85724 1 5845
2 85725 1 5845
2 85726 1 5845
2 85727 1 5845
2 85728 1 5845
2 85729 1 5845
2 85730 1 5845
2 85731 1 5860
2 85732 1 5860
2 85733 1 5860
2 85734 1 5861
2 85735 1 5861
2 85736 1 5861
2 85737 1 5861
2 85738 1 5861
2 85739 1 5861
2 85740 1 5866
2 85741 1 5866
2 85742 1 5866
2 85743 1 5866
2 85744 1 5868
2 85745 1 5868
2 85746 1 5868
2 85747 1 5868
2 85748 1 5868
2 85749 1 5869
2 85750 1 5869
2 85751 1 5871
2 85752 1 5871
2 85753 1 5871
2 85754 1 5871
2 85755 1 5879
2 85756 1 5879
2 85757 1 5879
2 85758 1 5879
2 85759 1 5879
2 85760 1 5880
2 85761 1 5880
2 85762 1 5880
2 85763 1 5880
2 85764 1 5880
2 85765 1 5880
2 85766 1 5880
2 85767 1 5880
2 85768 1 5882
2 85769 1 5882
2 85770 1 5882
2 85771 1 5882
2 85772 1 5890
2 85773 1 5890
2 85774 1 5890
2 85775 1 5890
2 85776 1 5890
2 85777 1 5892
2 85778 1 5892
2 85779 1 5897
2 85780 1 5897
2 85781 1 5905
2 85782 1 5905
2 85783 1 5905
2 85784 1 5906
2 85785 1 5906
2 85786 1 5923
2 85787 1 5923
2 85788 1 5924
2 85789 1 5924
2 85790 1 5924
2 85791 1 5924
2 85792 1 5925
2 85793 1 5925
2 85794 1 5939
2 85795 1 5939
2 85796 1 5939
2 85797 1 5946
2 85798 1 5946
2 85799 1 5946
2 85800 1 5953
2 85801 1 5953
2 85802 1 5953
2 85803 1 5953
2 85804 1 5953
2 85805 1 5960
2 85806 1 5960
2 85807 1 5967
2 85808 1 5967
2 85809 1 5980
2 85810 1 5980
2 85811 1 5980
2 85812 1 5980
2 85813 1 5980
2 85814 1 5980
2 85815 1 5980
2 85816 1 5980
2 85817 1 5980
2 85818 1 5981
2 85819 1 5981
2 85820 1 5981
2 85821 1 5981
2 85822 1 5982
2 85823 1 5982
2 85824 1 5982
2 85825 1 5982
2 85826 1 5982
2 85827 1 5982
2 85828 1 5982
2 85829 1 5982
2 85830 1 5982
2 85831 1 5984
2 85832 1 5984
2 85833 1 5984
2 85834 1 5987
2 85835 1 5987
2 85836 1 5987
2 85837 1 5987
2 85838 1 5987
2 85839 1 5987
2 85840 1 5987
2 85841 1 5987
2 85842 1 5987
2 85843 1 5987
2 85844 1 5987
2 85845 1 5987
2 85846 1 5987
2 85847 1 5987
2 85848 1 5987
2 85849 1 5987
2 85850 1 5988
2 85851 1 5988
2 85852 1 5989
2 85853 1 5989
2 85854 1 5992
2 85855 1 5992
2 85856 1 5999
2 85857 1 5999
2 85858 1 5999
2 85859 1 5999
2 85860 1 5999
2 85861 1 6005
2 85862 1 6005
2 85863 1 6005
2 85864 1 6013
2 85865 1 6013
2 85866 1 6013
2 85867 1 6013
2 85868 1 6015
2 85869 1 6015
2 85870 1 6015
2 85871 1 6015
2 85872 1 6015
2 85873 1 6018
2 85874 1 6018
2 85875 1 6018
2 85876 1 6018
2 85877 1 6018
2 85878 1 6018
2 85879 1 6018
2 85880 1 6018
2 85881 1 6018
2 85882 1 6025
2 85883 1 6025
2 85884 1 6025
2 85885 1 6025
2 85886 1 6035
2 85887 1 6035
2 85888 1 6035
2 85889 1 6035
2 85890 1 6035
2 85891 1 6035
2 85892 1 6035
2 85893 1 6035
2 85894 1 6035
2 85895 1 6035
2 85896 1 6035
2 85897 1 6035
2 85898 1 6035
2 85899 1 6035
2 85900 1 6036
2 85901 1 6036
2 85902 1 6036
2 85903 1 6036
2 85904 1 6037
2 85905 1 6037
2 85906 1 6037
2 85907 1 6038
2 85908 1 6038
2 85909 1 6038
2 85910 1 6046
2 85911 1 6046
2 85912 1 6046
2 85913 1 6046
2 85914 1 6046
2 85915 1 6046
2 85916 1 6046
2 85917 1 6046
2 85918 1 6046
2 85919 1 6046
2 85920 1 6046
2 85921 1 6047
2 85922 1 6047
2 85923 1 6048
2 85924 1 6048
2 85925 1 6048
2 85926 1 6048
2 85927 1 6048
2 85928 1 6052
2 85929 1 6052
2 85930 1 6052
2 85931 1 6052
2 85932 1 6053
2 85933 1 6053
2 85934 1 6066
2 85935 1 6066
2 85936 1 6066
2 85937 1 6067
2 85938 1 6067
2 85939 1 6067
2 85940 1 6067
2 85941 1 6067
2 85942 1 6067
2 85943 1 6067
2 85944 1 6075
2 85945 1 6075
2 85946 1 6075
2 85947 1 6076
2 85948 1 6076
2 85949 1 6076
2 85950 1 6076
2 85951 1 6078
2 85952 1 6078
2 85953 1 6078
2 85954 1 6078
2 85955 1 6080
2 85956 1 6080
2 85957 1 6088
2 85958 1 6088
2 85959 1 6088
2 85960 1 6088
2 85961 1 6088
2 85962 1 6088
2 85963 1 6088
2 85964 1 6088
2 85965 1 6088
2 85966 1 6091
2 85967 1 6091
2 85968 1 6091
2 85969 1 6091
2 85970 1 6091
2 85971 1 6091
2 85972 1 6091
2 85973 1 6091
2 85974 1 6092
2 85975 1 6092
2 85976 1 6093
2 85977 1 6093
2 85978 1 6093
2 85979 1 6102
2 85980 1 6102
2 85981 1 6111
2 85982 1 6111
2 85983 1 6112
2 85984 1 6112
2 85985 1 6112
2 85986 1 6112
2 85987 1 6116
2 85988 1 6116
2 85989 1 6116
2 85990 1 6137
2 85991 1 6137
2 85992 1 6137
2 85993 1 6138
2 85994 1 6138
2 85995 1 6139
2 85996 1 6139
2 85997 1 6140
2 85998 1 6140
2 85999 1 6161
2 86000 1 6161
2 86001 1 6161
2 86002 1 6161
2 86003 1 6161
2 86004 1 6161
2 86005 1 6161
2 86006 1 6161
2 86007 1 6161
2 86008 1 6161
2 86009 1 6163
2 86010 1 6163
2 86011 1 6163
2 86012 1 6164
2 86013 1 6164
2 86014 1 6174
2 86015 1 6174
2 86016 1 6174
2 86017 1 6174
2 86018 1 6174
2 86019 1 6174
2 86020 1 6174
2 86021 1 6174
2 86022 1 6174
2 86023 1 6179
2 86024 1 6179
2 86025 1 6179
2 86026 1 6192
2 86027 1 6192
2 86028 1 6192
2 86029 1 6192
2 86030 1 6192
2 86031 1 6192
2 86032 1 6192
2 86033 1 6192
2 86034 1 6192
2 86035 1 6192
2 86036 1 6192
2 86037 1 6192
2 86038 1 6193
2 86039 1 6193
2 86040 1 6193
2 86041 1 6193
2 86042 1 6193
2 86043 1 6193
2 86044 1 6193
2 86045 1 6193
2 86046 1 6193
2 86047 1 6193
2 86048 1 6197
2 86049 1 6197
2 86050 1 6197
2 86051 1 6197
2 86052 1 6197
2 86053 1 6197
2 86054 1 6197
2 86055 1 6197
2 86056 1 6197
2 86057 1 6197
2 86058 1 6197
2 86059 1 6197
2 86060 1 6197
2 86061 1 6197
2 86062 1 6197
2 86063 1 6197
2 86064 1 6197
2 86065 1 6197
2 86066 1 6197
2 86067 1 6197
2 86068 1 6197
2 86069 1 6197
2 86070 1 6206
2 86071 1 6206
2 86072 1 6206
2 86073 1 6213
2 86074 1 6213
2 86075 1 6213
2 86076 1 6228
2 86077 1 6228
2 86078 1 6229
2 86079 1 6229
2 86080 1 6232
2 86081 1 6232
2 86082 1 6232
2 86083 1 6232
2 86084 1 6232
2 86085 1 6232
2 86086 1 6232
2 86087 1 6233
2 86088 1 6233
2 86089 1 6233
2 86090 1 6255
2 86091 1 6255
2 86092 1 6255
2 86093 1 6255
2 86094 1 6255
2 86095 1 6255
2 86096 1 6255
2 86097 1 6255
2 86098 1 6255
2 86099 1 6256
2 86100 1 6256
2 86101 1 6257
2 86102 1 6257
2 86103 1 6257
2 86104 1 6260
2 86105 1 6260
2 86106 1 6260
2 86107 1 6260
2 86108 1 6260
2 86109 1 6262
2 86110 1 6262
2 86111 1 6270
2 86112 1 6270
2 86113 1 6273
2 86114 1 6273
2 86115 1 6273
2 86116 1 6286
2 86117 1 6286
2 86118 1 6286
2 86119 1 6286
2 86120 1 6287
2 86121 1 6287
2 86122 1 6288
2 86123 1 6288
2 86124 1 6288
2 86125 1 6288
2 86126 1 6289
2 86127 1 6289
2 86128 1 6289
2 86129 1 6296
2 86130 1 6296
2 86131 1 6296
2 86132 1 6296
2 86133 1 6296
2 86134 1 6296
2 86135 1 6296
2 86136 1 6296
2 86137 1 6296
2 86138 1 6296
2 86139 1 6296
2 86140 1 6296
2 86141 1 6296
2 86142 1 6296
2 86143 1 6296
2 86144 1 6296
2 86145 1 6296
2 86146 1 6303
2 86147 1 6303
2 86148 1 6303
2 86149 1 6306
2 86150 1 6306
2 86151 1 6306
2 86152 1 6306
2 86153 1 6318
2 86154 1 6318
2 86155 1 6318
2 86156 1 6319
2 86157 1 6319
2 86158 1 6319
2 86159 1 6319
2 86160 1 6319
2 86161 1 6319
2 86162 1 6319
2 86163 1 6319
2 86164 1 6320
2 86165 1 6320
2 86166 1 6320
2 86167 1 6327
2 86168 1 6327
2 86169 1 6327
2 86170 1 6327
2 86171 1 6327
2 86172 1 6327
2 86173 1 6327
2 86174 1 6327
2 86175 1 6327
2 86176 1 6327
2 86177 1 6327
2 86178 1 6327
2 86179 1 6329
2 86180 1 6329
2 86181 1 6338
2 86182 1 6338
2 86183 1 6338
2 86184 1 6338
2 86185 1 6346
2 86186 1 6346
2 86187 1 6346
2 86188 1 6346
2 86189 1 6346
2 86190 1 6346
2 86191 1 6346
2 86192 1 6346
2 86193 1 6346
2 86194 1 6348
2 86195 1 6348
2 86196 1 6348
2 86197 1 6348
2 86198 1 6348
2 86199 1 6348
2 86200 1 6348
2 86201 1 6349
2 86202 1 6349
2 86203 1 6358
2 86204 1 6358
2 86205 1 6358
2 86206 1 6361
2 86207 1 6361
2 86208 1 6361
2 86209 1 6361
2 86210 1 6361
2 86211 1 6361
2 86212 1 6361
2 86213 1 6362
2 86214 1 6362
2 86215 1 6364
2 86216 1 6364
2 86217 1 6364
2 86218 1 6364
2 86219 1 6367
2 86220 1 6367
2 86221 1 6370
2 86222 1 6370
2 86223 1 6378
2 86224 1 6378
2 86225 1 6385
2 86226 1 6385
2 86227 1 6398
2 86228 1 6398
2 86229 1 6398
2 86230 1 6398
2 86231 1 6398
2 86232 1 6403
2 86233 1 6403
2 86234 1 6404
2 86235 1 6404
2 86236 1 6404
2 86237 1 6404
2 86238 1 6404
2 86239 1 6404
2 86240 1 6404
2 86241 1 6407
2 86242 1 6407
2 86243 1 6407
2 86244 1 6407
2 86245 1 6418
2 86246 1 6418
2 86247 1 6420
2 86248 1 6420
2 86249 1 6420
2 86250 1 6421
2 86251 1 6421
2 86252 1 6421
2 86253 1 6421
2 86254 1 6434
2 86255 1 6434
2 86256 1 6439
2 86257 1 6439
2 86258 1 6439
2 86259 1 6439
2 86260 1 6439
2 86261 1 6439
2 86262 1 6439
2 86263 1 6458
2 86264 1 6458
2 86265 1 6472
2 86266 1 6472
2 86267 1 6472
2 86268 1 6472
2 86269 1 6472
2 86270 1 6472
2 86271 1 6472
2 86272 1 6473
2 86273 1 6473
2 86274 1 6473
2 86275 1 6485
2 86276 1 6485
2 86277 1 6487
2 86278 1 6487
2 86279 1 6487
2 86280 1 6487
2 86281 1 6487
2 86282 1 6505
2 86283 1 6505
2 86284 1 6505
2 86285 1 6505
2 86286 1 6505
2 86287 1 6505
2 86288 1 6506
2 86289 1 6506
2 86290 1 6506
2 86291 1 6506
2 86292 1 6506
2 86293 1 6515
2 86294 1 6515
2 86295 1 6520
2 86296 1 6520
2 86297 1 6520
2 86298 1 6528
2 86299 1 6528
2 86300 1 6528
2 86301 1 6528
2 86302 1 6528
2 86303 1 6528
2 86304 1 6528
2 86305 1 6528
2 86306 1 6528
2 86307 1 6528
2 86308 1 6528
2 86309 1 6528
2 86310 1 6528
2 86311 1 6528
2 86312 1 6528
2 86313 1 6528
2 86314 1 6528
2 86315 1 6528
2 86316 1 6528
2 86317 1 6529
2 86318 1 6529
2 86319 1 6529
2 86320 1 6538
2 86321 1 6538
2 86322 1 6557
2 86323 1 6557
2 86324 1 6559
2 86325 1 6559
2 86326 1 6559
2 86327 1 6560
2 86328 1 6560
2 86329 1 6560
2 86330 1 6567
2 86331 1 6567
2 86332 1 6567
2 86333 1 6567
2 86334 1 6567
2 86335 1 6567
2 86336 1 6567
2 86337 1 6572
2 86338 1 6572
2 86339 1 6573
2 86340 1 6573
2 86341 1 6573
2 86342 1 6576
2 86343 1 6576
2 86344 1 6577
2 86345 1 6577
2 86346 1 6577
2 86347 1 6577
2 86348 1 6577
2 86349 1 6577
2 86350 1 6577
2 86351 1 6577
2 86352 1 6577
2 86353 1 6577
2 86354 1 6577
2 86355 1 6580
2 86356 1 6580
2 86357 1 6580
2 86358 1 6580
2 86359 1 6581
2 86360 1 6581
2 86361 1 6592
2 86362 1 6592
2 86363 1 6601
2 86364 1 6601
2 86365 1 6604
2 86366 1 6604
2 86367 1 6604
2 86368 1 6605
2 86369 1 6605
2 86370 1 6605
2 86371 1 6605
2 86372 1 6605
2 86373 1 6606
2 86374 1 6606
2 86375 1 6614
2 86376 1 6614
2 86377 1 6614
2 86378 1 6614
2 86379 1 6614
2 86380 1 6614
2 86381 1 6614
2 86382 1 6614
2 86383 1 6614
2 86384 1 6614
2 86385 1 6614
2 86386 1 6622
2 86387 1 6622
2 86388 1 6625
2 86389 1 6625
2 86390 1 6625
2 86391 1 6625
2 86392 1 6625
2 86393 1 6625
2 86394 1 6625
2 86395 1 6626
2 86396 1 6626
2 86397 1 6626
2 86398 1 6639
2 86399 1 6639
2 86400 1 6639
2 86401 1 6639
2 86402 1 6639
2 86403 1 6639
2 86404 1 6639
2 86405 1 6639
2 86406 1 6639
2 86407 1 6639
2 86408 1 6639
2 86409 1 6639
2 86410 1 6639
2 86411 1 6640
2 86412 1 6640
2 86413 1 6641
2 86414 1 6641
2 86415 1 6641
2 86416 1 6641
2 86417 1 6650
2 86418 1 6650
2 86419 1 6650
2 86420 1 6650
2 86421 1 6654
2 86422 1 6654
2 86423 1 6654
2 86424 1 6654
2 86425 1 6657
2 86426 1 6657
2 86427 1 6657
2 86428 1 6657
2 86429 1 6657
2 86430 1 6666
2 86431 1 6666
2 86432 1 6666
2 86433 1 6666
2 86434 1 6666
2 86435 1 6666
2 86436 1 6666
2 86437 1 6666
2 86438 1 6666
2 86439 1 6667
2 86440 1 6667
2 86441 1 6669
2 86442 1 6669
2 86443 1 6674
2 86444 1 6674
2 86445 1 6674
2 86446 1 6674
2 86447 1 6674
2 86448 1 6674
2 86449 1 6674
2 86450 1 6683
2 86451 1 6683
2 86452 1 6683
2 86453 1 6683
2 86454 1 6683
2 86455 1 6683
2 86456 1 6683
2 86457 1 6683
2 86458 1 6695
2 86459 1 6695
2 86460 1 6695
2 86461 1 6695
2 86462 1 6695
2 86463 1 6696
2 86464 1 6696
2 86465 1 6696
2 86466 1 6698
2 86467 1 6698
2 86468 1 6699
2 86469 1 6699
2 86470 1 6699
2 86471 1 6699
2 86472 1 6699
2 86473 1 6701
2 86474 1 6701
2 86475 1 6701
2 86476 1 6706
2 86477 1 6706
2 86478 1 6706
2 86479 1 6706
2 86480 1 6706
2 86481 1 6706
2 86482 1 6713
2 86483 1 6713
2 86484 1 6716
2 86485 1 6716
2 86486 1 6716
2 86487 1 6716
2 86488 1 6716
2 86489 1 6716
2 86490 1 6716
2 86491 1 6716
2 86492 1 6717
2 86493 1 6717
2 86494 1 6717
2 86495 1 6717
2 86496 1 6717
2 86497 1 6725
2 86498 1 6725
2 86499 1 6725
2 86500 1 6725
2 86501 1 6725
2 86502 1 6726
2 86503 1 6726
2 86504 1 6726
2 86505 1 6726
2 86506 1 6726
2 86507 1 6726
2 86508 1 6726
2 86509 1 6726
2 86510 1 6726
2 86511 1 6727
2 86512 1 6727
2 86513 1 6728
2 86514 1 6728
2 86515 1 6729
2 86516 1 6729
2 86517 1 6737
2 86518 1 6737
2 86519 1 6738
2 86520 1 6738
2 86521 1 6741
2 86522 1 6741
2 86523 1 6741
2 86524 1 6753
2 86525 1 6753
2 86526 1 6753
2 86527 1 6753
2 86528 1 6753
2 86529 1 6753
2 86530 1 6753
2 86531 1 6763
2 86532 1 6763
2 86533 1 6763
2 86534 1 6775
2 86535 1 6775
2 86536 1 6775
2 86537 1 6777
2 86538 1 6777
2 86539 1 6777
2 86540 1 6777
2 86541 1 6786
2 86542 1 6786
2 86543 1 6787
2 86544 1 6787
2 86545 1 6792
2 86546 1 6792
2 86547 1 6792
2 86548 1 6792
2 86549 1 6792
2 86550 1 6792
2 86551 1 6792
2 86552 1 6792
2 86553 1 6792
2 86554 1 6792
2 86555 1 6793
2 86556 1 6793
2 86557 1 6793
2 86558 1 6793
2 86559 1 6793
2 86560 1 6801
2 86561 1 6801
2 86562 1 6802
2 86563 1 6802
2 86564 1 6804
2 86565 1 6804
2 86566 1 6807
2 86567 1 6807
2 86568 1 6807
2 86569 1 6807
2 86570 1 6807
2 86571 1 6807
2 86572 1 6807
2 86573 1 6807
2 86574 1 6807
2 86575 1 6807
2 86576 1 6807
2 86577 1 6807
2 86578 1 6807
2 86579 1 6807
2 86580 1 6807
2 86581 1 6808
2 86582 1 6808
2 86583 1 6808
2 86584 1 6808
2 86585 1 6809
2 86586 1 6809
2 86587 1 6813
2 86588 1 6813
2 86589 1 6821
2 86590 1 6821
2 86591 1 6824
2 86592 1 6824
2 86593 1 6825
2 86594 1 6825
2 86595 1 6846
2 86596 1 6846
2 86597 1 6846
2 86598 1 6846
2 86599 1 6846
2 86600 1 6846
2 86601 1 6846
2 86602 1 6846
2 86603 1 6846
2 86604 1 6846
2 86605 1 6846
2 86606 1 6846
2 86607 1 6846
2 86608 1 6846
2 86609 1 6846
2 86610 1 6846
2 86611 1 6846
2 86612 1 6846
2 86613 1 6846
2 86614 1 6846
2 86615 1 6846
2 86616 1 6846
2 86617 1 6846
2 86618 1 6846
2 86619 1 6846
2 86620 1 6847
2 86621 1 6847
2 86622 1 6847
2 86623 1 6847
2 86624 1 6848
2 86625 1 6848
2 86626 1 6848
2 86627 1 6848
2 86628 1 6848
2 86629 1 6848
2 86630 1 6848
2 86631 1 6848
2 86632 1 6848
2 86633 1 6848
2 86634 1 6848
2 86635 1 6848
2 86636 1 6848
2 86637 1 6848
2 86638 1 6856
2 86639 1 6856
2 86640 1 6856
2 86641 1 6857
2 86642 1 6857
2 86643 1 6865
2 86644 1 6865
2 86645 1 6865
2 86646 1 6865
2 86647 1 6865
2 86648 1 6865
2 86649 1 6865
2 86650 1 6865
2 86651 1 6865
2 86652 1 6865
2 86653 1 6865
2 86654 1 6865
2 86655 1 6865
2 86656 1 6865
2 86657 1 6865
2 86658 1 6865
2 86659 1 6866
2 86660 1 6866
2 86661 1 6866
2 86662 1 6866
2 86663 1 6870
2 86664 1 6870
2 86665 1 6870
2 86666 1 6881
2 86667 1 6881
2 86668 1 6884
2 86669 1 6884
2 86670 1 6884
2 86671 1 6884
2 86672 1 6884
2 86673 1 6884
2 86674 1 6884
2 86675 1 6884
2 86676 1 6893
2 86677 1 6893
2 86678 1 6893
2 86679 1 6893
2 86680 1 6893
2 86681 1 6893
2 86682 1 6893
2 86683 1 6894
2 86684 1 6894
2 86685 1 6895
2 86686 1 6895
2 86687 1 6903
2 86688 1 6903
2 86689 1 6913
2 86690 1 6913
2 86691 1 6914
2 86692 1 6914
2 86693 1 6914
2 86694 1 6914
2 86695 1 6914
2 86696 1 6914
2 86697 1 6914
2 86698 1 6914
2 86699 1 6914
2 86700 1 6914
2 86701 1 6914
2 86702 1 6914
2 86703 1 6914
2 86704 1 6914
2 86705 1 6914
2 86706 1 6914
2 86707 1 6914
2 86708 1 6914
2 86709 1 6914
2 86710 1 6915
2 86711 1 6915
2 86712 1 6916
2 86713 1 6916
2 86714 1 6917
2 86715 1 6917
2 86716 1 6918
2 86717 1 6918
2 86718 1 6927
2 86719 1 6927
2 86720 1 6927
2 86721 1 6927
2 86722 1 6928
2 86723 1 6928
2 86724 1 6928
2 86725 1 6928
2 86726 1 6928
2 86727 1 6928
2 86728 1 6928
2 86729 1 6928
2 86730 1 6929
2 86731 1 6929
2 86732 1 6929
2 86733 1 6929
2 86734 1 6929
2 86735 1 6929
2 86736 1 6929
2 86737 1 6929
2 86738 1 6930
2 86739 1 6930
2 86740 1 6930
2 86741 1 6930
2 86742 1 6930
2 86743 1 6931
2 86744 1 6931
2 86745 1 6936
2 86746 1 6936
2 86747 1 6941
2 86748 1 6941
2 86749 1 6944
2 86750 1 6944
2 86751 1 6945
2 86752 1 6945
2 86753 1 6957
2 86754 1 6957
2 86755 1 6957
2 86756 1 6957
2 86757 1 6957
2 86758 1 6957
2 86759 1 6957
2 86760 1 6957
2 86761 1 6957
2 86762 1 6957
2 86763 1 6957
2 86764 1 6957
2 86765 1 6957
2 86766 1 6957
2 86767 1 6957
2 86768 1 6957
2 86769 1 6957
2 86770 1 6958
2 86771 1 6958
2 86772 1 6958
2 86773 1 6959
2 86774 1 6959
2 86775 1 6959
2 86776 1 6967
2 86777 1 6967
2 86778 1 6972
2 86779 1 6972
2 86780 1 6987
2 86781 1 6987
2 86782 1 6988
2 86783 1 6988
2 86784 1 6995
2 86785 1 6995
2 86786 1 6999
2 86787 1 6999
2 86788 1 6999
2 86789 1 6999
2 86790 1 6999
2 86791 1 7002
2 86792 1 7002
2 86793 1 7002
2 86794 1 7002
2 86795 1 7002
2 86796 1 7002
2 86797 1 7002
2 86798 1 7002
2 86799 1 7002
2 86800 1 7002
2 86801 1 7002
2 86802 1 7002
2 86803 1 7010
2 86804 1 7010
2 86805 1 7010
2 86806 1 7010
2 86807 1 7010
2 86808 1 7030
2 86809 1 7030
2 86810 1 7035
2 86811 1 7035
2 86812 1 7035
2 86813 1 7035
2 86814 1 7035
2 86815 1 7035
2 86816 1 7035
2 86817 1 7035
2 86818 1 7035
2 86819 1 7037
2 86820 1 7037
2 86821 1 7055
2 86822 1 7055
2 86823 1 7055
2 86824 1 7062
2 86825 1 7062
2 86826 1 7062
2 86827 1 7075
2 86828 1 7075
2 86829 1 7076
2 86830 1 7076
2 86831 1 7076
2 86832 1 7076
2 86833 1 7076
2 86834 1 7076
2 86835 1 7076
2 86836 1 7076
2 86837 1 7076
2 86838 1 7076
2 86839 1 7076
2 86840 1 7076
2 86841 1 7076
2 86842 1 7076
2 86843 1 7076
2 86844 1 7076
2 86845 1 7076
2 86846 1 7078
2 86847 1 7078
2 86848 1 7078
2 86849 1 7079
2 86850 1 7079
2 86851 1 7095
2 86852 1 7095
2 86853 1 7095
2 86854 1 7096
2 86855 1 7096
2 86856 1 7098
2 86857 1 7098
2 86858 1 7103
2 86859 1 7103
2 86860 1 7103
2 86861 1 7103
2 86862 1 7103
2 86863 1 7109
2 86864 1 7109
2 86865 1 7109
2 86866 1 7109
2 86867 1 7109
2 86868 1 7109
2 86869 1 7109
2 86870 1 7109
2 86871 1 7109
2 86872 1 7109
2 86873 1 7109
2 86874 1 7118
2 86875 1 7118
2 86876 1 7118
2 86877 1 7118
2 86878 1 7118
2 86879 1 7118
2 86880 1 7118
2 86881 1 7119
2 86882 1 7119
2 86883 1 7122
2 86884 1 7122
2 86885 1 7123
2 86886 1 7123
2 86887 1 7123
2 86888 1 7123
2 86889 1 7123
2 86890 1 7123
2 86891 1 7124
2 86892 1 7124
2 86893 1 7124
2 86894 1 7125
2 86895 1 7125
2 86896 1 7125
2 86897 1 7125
2 86898 1 7125
2 86899 1 7126
2 86900 1 7126
2 86901 1 7126
2 86902 1 7131
2 86903 1 7131
2 86904 1 7139
2 86905 1 7139
2 86906 1 7140
2 86907 1 7140
2 86908 1 7140
2 86909 1 7151
2 86910 1 7151
2 86911 1 7151
2 86912 1 7157
2 86913 1 7157
2 86914 1 7157
2 86915 1 7157
2 86916 1 7169
2 86917 1 7169
2 86918 1 7169
2 86919 1 7170
2 86920 1 7170
2 86921 1 7171
2 86922 1 7171
2 86923 1 7171
2 86924 1 7171
2 86925 1 7171
2 86926 1 7171
2 86927 1 7171
2 86928 1 7171
2 86929 1 7171
2 86930 1 7171
2 86931 1 7171
2 86932 1 7171
2 86933 1 7171
2 86934 1 7171
2 86935 1 7171
2 86936 1 7171
2 86937 1 7171
2 86938 1 7184
2 86939 1 7184
2 86940 1 7184
2 86941 1 7184
2 86942 1 7184
2 86943 1 7184
2 86944 1 7184
2 86945 1 7184
2 86946 1 7184
2 86947 1 7184
2 86948 1 7184
2 86949 1 7184
2 86950 1 7184
2 86951 1 7184
2 86952 1 7184
2 86953 1 7184
2 86954 1 7184
2 86955 1 7184
2 86956 1 7184
2 86957 1 7184
2 86958 1 7184
2 86959 1 7184
2 86960 1 7184
2 86961 1 7184
2 86962 1 7184
2 86963 1 7184
2 86964 1 7184
2 86965 1 7184
2 86966 1 7184
2 86967 1 7184
2 86968 1 7184
2 86969 1 7184
2 86970 1 7184
2 86971 1 7184
2 86972 1 7184
2 86973 1 7184
2 86974 1 7184
2 86975 1 7184
2 86976 1 7184
2 86977 1 7184
2 86978 1 7184
2 86979 1 7184
2 86980 1 7184
2 86981 1 7184
2 86982 1 7184
2 86983 1 7184
2 86984 1 7184
2 86985 1 7184
2 86986 1 7184
2 86987 1 7184
2 86988 1 7184
2 86989 1 7184
2 86990 1 7184
2 86991 1 7184
2 86992 1 7184
2 86993 1 7184
2 86994 1 7184
2 86995 1 7184
2 86996 1 7184
2 86997 1 7184
2 86998 1 7184
2 86999 1 7184
2 87000 1 7184
2 87001 1 7184
2 87002 1 7184
2 87003 1 7184
2 87004 1 7184
2 87005 1 7184
2 87006 1 7184
2 87007 1 7184
2 87008 1 7184
2 87009 1 7184
2 87010 1 7184
2 87011 1 7185
2 87012 1 7185
2 87013 1 7185
2 87014 1 7185
2 87015 1 7185
2 87016 1 7186
2 87017 1 7186
2 87018 1 7186
2 87019 1 7186
2 87020 1 7186
2 87021 1 7186
2 87022 1 7186
2 87023 1 7187
2 87024 1 7187
2 87025 1 7187
2 87026 1 7187
2 87027 1 7188
2 87028 1 7188
2 87029 1 7191
2 87030 1 7191
2 87031 1 7191
2 87032 1 7193
2 87033 1 7193
2 87034 1 7201
2 87035 1 7201
2 87036 1 7202
2 87037 1 7202
2 87038 1 7202
2 87039 1 7202
2 87040 1 7202
2 87041 1 7203
2 87042 1 7203
2 87043 1 7203
2 87044 1 7204
2 87045 1 7204
2 87046 1 7205
2 87047 1 7205
2 87048 1 7206
2 87049 1 7206
2 87050 1 7206
2 87051 1 7213
2 87052 1 7213
2 87053 1 7217
2 87054 1 7217
2 87055 1 7225
2 87056 1 7225
2 87057 1 7225
2 87058 1 7226
2 87059 1 7226
2 87060 1 7226
2 87061 1 7226
2 87062 1 7226
2 87063 1 7226
2 87064 1 7226
2 87065 1 7226
2 87066 1 7226
2 87067 1 7226
2 87068 1 7226
2 87069 1 7226
2 87070 1 7226
2 87071 1 7226
2 87072 1 7226
2 87073 1 7226
2 87074 1 7235
2 87075 1 7235
2 87076 1 7235
2 87077 1 7236
2 87078 1 7236
2 87079 1 7236
2 87080 1 7236
2 87081 1 7239
2 87082 1 7239
2 87083 1 7239
2 87084 1 7252
2 87085 1 7252
2 87086 1 7252
2 87087 1 7252
2 87088 1 7253
2 87089 1 7253
2 87090 1 7253
2 87091 1 7253
2 87092 1 7253
2 87093 1 7253
2 87094 1 7253
2 87095 1 7253
2 87096 1 7253
2 87097 1 7253
2 87098 1 7253
2 87099 1 7254
2 87100 1 7254
2 87101 1 7257
2 87102 1 7257
2 87103 1 7258
2 87104 1 7258
2 87105 1 7258
2 87106 1 7258
2 87107 1 7258
2 87108 1 7258
2 87109 1 7258
2 87110 1 7258
2 87111 1 7258
2 87112 1 7258
2 87113 1 7258
2 87114 1 7258
2 87115 1 7258
2 87116 1 7258
2 87117 1 7266
2 87118 1 7266
2 87119 1 7275
2 87120 1 7275
2 87121 1 7276
2 87122 1 7276
2 87123 1 7279
2 87124 1 7279
2 87125 1 7279
2 87126 1 7279
2 87127 1 7279
2 87128 1 7280
2 87129 1 7280
2 87130 1 7282
2 87131 1 7282
2 87132 1 7282
2 87133 1 7282
2 87134 1 7282
2 87135 1 7282
2 87136 1 7283
2 87137 1 7283
2 87138 1 7284
2 87139 1 7284
2 87140 1 7284
2 87141 1 7284
2 87142 1 7284
2 87143 1 7284
2 87144 1 7284
2 87145 1 7303
2 87146 1 7303
2 87147 1 7304
2 87148 1 7304
2 87149 1 7304
2 87150 1 7304
2 87151 1 7305
2 87152 1 7305
2 87153 1 7305
2 87154 1 7305
2 87155 1 7305
2 87156 1 7306
2 87157 1 7306
2 87158 1 7307
2 87159 1 7307
2 87160 1 7324
2 87161 1 7324
2 87162 1 7324
2 87163 1 7328
2 87164 1 7328
2 87165 1 7328
2 87166 1 7328
2 87167 1 7328
2 87168 1 7328
2 87169 1 7329
2 87170 1 7329
2 87171 1 7329
2 87172 1 7329
2 87173 1 7329
2 87174 1 7335
2 87175 1 7335
2 87176 1 7335
2 87177 1 7335
2 87178 1 7361
2 87179 1 7361
2 87180 1 7361
2 87181 1 7361
2 87182 1 7369
2 87183 1 7369
2 87184 1 7369
2 87185 1 7369
2 87186 1 7369
2 87187 1 7370
2 87188 1 7370
2 87189 1 7373
2 87190 1 7373
2 87191 1 7373
2 87192 1 7374
2 87193 1 7374
2 87194 1 7394
2 87195 1 7394
2 87196 1 7394
2 87197 1 7394
2 87198 1 7394
2 87199 1 7394
2 87200 1 7394
2 87201 1 7394
2 87202 1 7394
2 87203 1 7394
2 87204 1 7394
2 87205 1 7394
2 87206 1 7394
2 87207 1 7394
2 87208 1 7394
2 87209 1 7394
2 87210 1 7394
2 87211 1 7394
2 87212 1 7394
2 87213 1 7395
2 87214 1 7395
2 87215 1 7410
2 87216 1 7410
2 87217 1 7418
2 87218 1 7418
2 87219 1 7418
2 87220 1 7418
2 87221 1 7418
2 87222 1 7419
2 87223 1 7419
2 87224 1 7431
2 87225 1 7431
2 87226 1 7443
2 87227 1 7443
2 87228 1 7443
2 87229 1 7443
2 87230 1 7444
2 87231 1 7444
2 87232 1 7448
2 87233 1 7448
2 87234 1 7448
2 87235 1 7448
2 87236 1 7448
2 87237 1 7448
2 87238 1 7448
2 87239 1 7449
2 87240 1 7449
2 87241 1 7449
2 87242 1 7449
2 87243 1 7449
2 87244 1 7452
2 87245 1 7452
2 87246 1 7452
2 87247 1 7452
2 87248 1 7452
2 87249 1 7452
2 87250 1 7452
2 87251 1 7452
2 87252 1 7452
2 87253 1 7452
2 87254 1 7452
2 87255 1 7452
2 87256 1 7452
2 87257 1 7452
2 87258 1 7455
2 87259 1 7455
2 87260 1 7461
2 87261 1 7461
2 87262 1 7461
2 87263 1 7461
2 87264 1 7461
2 87265 1 7461
2 87266 1 7473
2 87267 1 7473
2 87268 1 7473
2 87269 1 7474
2 87270 1 7474
2 87271 1 7474
2 87272 1 7476
2 87273 1 7476
2 87274 1 7486
2 87275 1 7486
2 87276 1 7486
2 87277 1 7486
2 87278 1 7486
2 87279 1 7486
2 87280 1 7499
2 87281 1 7499
2 87282 1 7500
2 87283 1 7500
2 87284 1 7503
2 87285 1 7503
2 87286 1 7503
2 87287 1 7511
2 87288 1 7511
2 87289 1 7520
2 87290 1 7520
2 87291 1 7521
2 87292 1 7521
2 87293 1 7530
2 87294 1 7530
2 87295 1 7530
2 87296 1 7530
2 87297 1 7530
2 87298 1 7530
2 87299 1 7530
2 87300 1 7532
2 87301 1 7532
2 87302 1 7540
2 87303 1 7540
2 87304 1 7540
2 87305 1 7540
2 87306 1 7540
2 87307 1 7540
2 87308 1 7540
2 87309 1 7540
2 87310 1 7540
2 87311 1 7540
2 87312 1 7540
2 87313 1 7540
2 87314 1 7540
2 87315 1 7540
2 87316 1 7540
2 87317 1 7541
2 87318 1 7541
2 87319 1 7541
2 87320 1 7541
2 87321 1 7541
2 87322 1 7541
2 87323 1 7541
2 87324 1 7541
2 87325 1 7541
2 87326 1 7541
2 87327 1 7541
2 87328 1 7541
2 87329 1 7541
2 87330 1 7541
2 87331 1 7541
2 87332 1 7541
2 87333 1 7541
2 87334 1 7542
2 87335 1 7542
2 87336 1 7542
2 87337 1 7542
2 87338 1 7542
2 87339 1 7542
2 87340 1 7545
2 87341 1 7545
2 87342 1 7552
2 87343 1 7552
2 87344 1 7552
2 87345 1 7552
2 87346 1 7552
2 87347 1 7552
2 87348 1 7563
2 87349 1 7563
2 87350 1 7564
2 87351 1 7564
2 87352 1 7564
2 87353 1 7564
2 87354 1 7564
2 87355 1 7564
2 87356 1 7564
2 87357 1 7564
2 87358 1 7564
2 87359 1 7564
2 87360 1 7564
2 87361 1 7564
2 87362 1 7564
2 87363 1 7564
2 87364 1 7564
2 87365 1 7564
2 87366 1 7564
2 87367 1 7564
2 87368 1 7564
2 87369 1 7564
2 87370 1 7564
2 87371 1 7564
2 87372 1 7564
2 87373 1 7564
2 87374 1 7564
2 87375 1 7564
2 87376 1 7564
2 87377 1 7564
2 87378 1 7564
2 87379 1 7564
2 87380 1 7564
2 87381 1 7564
2 87382 1 7564
2 87383 1 7564
2 87384 1 7565
2 87385 1 7565
2 87386 1 7565
2 87387 1 7565
2 87388 1 7568
2 87389 1 7568
2 87390 1 7568
2 87391 1 7568
2 87392 1 7568
2 87393 1 7568
2 87394 1 7568
2 87395 1 7569
2 87396 1 7569
2 87397 1 7570
2 87398 1 7570
2 87399 1 7570
2 87400 1 7570
2 87401 1 7570
2 87402 1 7570
2 87403 1 7570
2 87404 1 7570
2 87405 1 7570
2 87406 1 7570
2 87407 1 7570
2 87408 1 7570
2 87409 1 7570
2 87410 1 7570
2 87411 1 7570
2 87412 1 7570
2 87413 1 7578
2 87414 1 7578
2 87415 1 7578
2 87416 1 7578
2 87417 1 7578
2 87418 1 7578
2 87419 1 7578
2 87420 1 7578
2 87421 1 7578
2 87422 1 7578
2 87423 1 7579
2 87424 1 7579
2 87425 1 7579
2 87426 1 7579
2 87427 1 7579
2 87428 1 7579
2 87429 1 7579
2 87430 1 7587
2 87431 1 7587
2 87432 1 7596
2 87433 1 7596
2 87434 1 7596
2 87435 1 7596
2 87436 1 7596
2 87437 1 7596
2 87438 1 7596
2 87439 1 7596
2 87440 1 7596
2 87441 1 7596
2 87442 1 7596
2 87443 1 7615
2 87444 1 7615
2 87445 1 7615
2 87446 1 7616
2 87447 1 7616
2 87448 1 7616
2 87449 1 7616
2 87450 1 7616
2 87451 1 7616
2 87452 1 7617
2 87453 1 7617
2 87454 1 7617
2 87455 1 7629
2 87456 1 7629
2 87457 1 7629
2 87458 1 7629
2 87459 1 7629
2 87460 1 7630
2 87461 1 7630
2 87462 1 7630
2 87463 1 7630
2 87464 1 7630
2 87465 1 7630
2 87466 1 7630
2 87467 1 7630
2 87468 1 7630
2 87469 1 7630
2 87470 1 7630
2 87471 1 7631
2 87472 1 7631
2 87473 1 7631
2 87474 1 7631
2 87475 1 7631
2 87476 1 7631
2 87477 1 7636
2 87478 1 7636
2 87479 1 7636
2 87480 1 7636
2 87481 1 7636
2 87482 1 7636
2 87483 1 7636
2 87484 1 7636
2 87485 1 7636
2 87486 1 7636
2 87487 1 7637
2 87488 1 7637
2 87489 1 7638
2 87490 1 7638
2 87491 1 7638
2 87492 1 7638
2 87493 1 7638
2 87494 1 7638
2 87495 1 7638
2 87496 1 7638
2 87497 1 7638
2 87498 1 7638
2 87499 1 7638
2 87500 1 7638
2 87501 1 7638
2 87502 1 7638
2 87503 1 7638
2 87504 1 7646
2 87505 1 7646
2 87506 1 7646
2 87507 1 7646
2 87508 1 7647
2 87509 1 7647
2 87510 1 7648
2 87511 1 7648
2 87512 1 7656
2 87513 1 7656
2 87514 1 7666
2 87515 1 7666
2 87516 1 7666
2 87517 1 7666
2 87518 1 7666
2 87519 1 7674
2 87520 1 7674
2 87521 1 7674
2 87522 1 7678
2 87523 1 7678
2 87524 1 7678
2 87525 1 7678
2 87526 1 7686
2 87527 1 7686
2 87528 1 7686
2 87529 1 7696
2 87530 1 7696
2 87531 1 7697
2 87532 1 7697
2 87533 1 7704
2 87534 1 7704
2 87535 1 7704
2 87536 1 7715
2 87537 1 7715
2 87538 1 7719
2 87539 1 7719
2 87540 1 7719
2 87541 1 7720
2 87542 1 7720
2 87543 1 7720
2 87544 1 7720
2 87545 1 7720
2 87546 1 7720
2 87547 1 7721
2 87548 1 7721
2 87549 1 7729
2 87550 1 7729
2 87551 1 7729
2 87552 1 7730
2 87553 1 7730
2 87554 1 7731
2 87555 1 7731
2 87556 1 7731
2 87557 1 7731
2 87558 1 7731
2 87559 1 7731
2 87560 1 7731
2 87561 1 7731
2 87562 1 7731
2 87563 1 7731
2 87564 1 7732
2 87565 1 7732
2 87566 1 7732
2 87567 1 7732
2 87568 1 7733
2 87569 1 7733
2 87570 1 7733
2 87571 1 7733
2 87572 1 7733
2 87573 1 7733
2 87574 1 7733
2 87575 1 7733
2 87576 1 7733
2 87577 1 7744
2 87578 1 7744
2 87579 1 7744
2 87580 1 7748
2 87581 1 7748
2 87582 1 7748
2 87583 1 7748
2 87584 1 7751
2 87585 1 7751
2 87586 1 7752
2 87587 1 7752
2 87588 1 7752
2 87589 1 7760
2 87590 1 7760
2 87591 1 7760
2 87592 1 7760
2 87593 1 7769
2 87594 1 7769
2 87595 1 7773
2 87596 1 7773
2 87597 1 7773
2 87598 1 7773
2 87599 1 7791
2 87600 1 7791
2 87601 1 7791
2 87602 1 7791
2 87603 1 7791
2 87604 1 7791
2 87605 1 7791
2 87606 1 7791
2 87607 1 7792
2 87608 1 7792
2 87609 1 7792
2 87610 1 7792
2 87611 1 7792
2 87612 1 7794
2 87613 1 7794
2 87614 1 7794
2 87615 1 7794
2 87616 1 7794
2 87617 1 7794
2 87618 1 7794
2 87619 1 7794
2 87620 1 7794
2 87621 1 7794
2 87622 1 7794
2 87623 1 7794
2 87624 1 7794
2 87625 1 7794
2 87626 1 7794
2 87627 1 7794
2 87628 1 7794
2 87629 1 7801
2 87630 1 7801
2 87631 1 7801
2 87632 1 7809
2 87633 1 7809
2 87634 1 7828
2 87635 1 7828
2 87636 1 7828
2 87637 1 7828
2 87638 1 7828
2 87639 1 7828
2 87640 1 7828
2 87641 1 7828
2 87642 1 7828
2 87643 1 7828
2 87644 1 7828
2 87645 1 7828
2 87646 1 7828
2 87647 1 7828
2 87648 1 7828
2 87649 1 7828
2 87650 1 7828
2 87651 1 7828
2 87652 1 7829
2 87653 1 7829
2 87654 1 7829
2 87655 1 7829
2 87656 1 7829
2 87657 1 7829
2 87658 1 7829
2 87659 1 7829
2 87660 1 7829
2 87661 1 7830
2 87662 1 7830
2 87663 1 7830
2 87664 1 7830
2 87665 1 7830
2 87666 1 7830
2 87667 1 7831
2 87668 1 7831
2 87669 1 7831
2 87670 1 7833
2 87671 1 7833
2 87672 1 7833
2 87673 1 7833
2 87674 1 7833
2 87675 1 7833
2 87676 1 7833
2 87677 1 7834
2 87678 1 7834
2 87679 1 7834
2 87680 1 7834
2 87681 1 7834
2 87682 1 7834
2 87683 1 7834
2 87684 1 7834
2 87685 1 7834
2 87686 1 7834
2 87687 1 7834
2 87688 1 7834
2 87689 1 7834
2 87690 1 7848
2 87691 1 7848
2 87692 1 7848
2 87693 1 7848
2 87694 1 7850
2 87695 1 7850
2 87696 1 7850
2 87697 1 7850
2 87698 1 7850
2 87699 1 7853
2 87700 1 7853
2 87701 1 7853
2 87702 1 7853
2 87703 1 7853
2 87704 1 7853
2 87705 1 7853
2 87706 1 7854
2 87707 1 7854
2 87708 1 7854
2 87709 1 7854
2 87710 1 7854
2 87711 1 7854
2 87712 1 7854
2 87713 1 7854
2 87714 1 7854
2 87715 1 7854
2 87716 1 7854
2 87717 1 7854
2 87718 1 7854
2 87719 1 7854
2 87720 1 7854
2 87721 1 7854
2 87722 1 7854
2 87723 1 7854
2 87724 1 7854
2 87725 1 7854
2 87726 1 7854
2 87727 1 7854
2 87728 1 7854
2 87729 1 7854
2 87730 1 7854
2 87731 1 7854
2 87732 1 7854
2 87733 1 7854
2 87734 1 7854
2 87735 1 7854
2 87736 1 7854
2 87737 1 7854
2 87738 1 7854
2 87739 1 7854
2 87740 1 7854
2 87741 1 7854
2 87742 1 7854
2 87743 1 7854
2 87744 1 7854
2 87745 1 7854
2 87746 1 7854
2 87747 1 7854
2 87748 1 7854
2 87749 1 7854
2 87750 1 7854
2 87751 1 7854
2 87752 1 7854
2 87753 1 7854
2 87754 1 7854
2 87755 1 7854
2 87756 1 7854
2 87757 1 7854
2 87758 1 7854
2 87759 1 7854
2 87760 1 7854
2 87761 1 7854
2 87762 1 7854
2 87763 1 7855
2 87764 1 7855
2 87765 1 7855
2 87766 1 7856
2 87767 1 7856
2 87768 1 7856
2 87769 1 7856
2 87770 1 7856
2 87771 1 7856
2 87772 1 7858
2 87773 1 7858
2 87774 1 7858
2 87775 1 7858
2 87776 1 7865
2 87777 1 7865
2 87778 1 7865
2 87779 1 7865
2 87780 1 7865
2 87781 1 7865
2 87782 1 7865
2 87783 1 7865
2 87784 1 7865
2 87785 1 7865
2 87786 1 7865
2 87787 1 7865
2 87788 1 7865
2 87789 1 7865
2 87790 1 7865
2 87791 1 7865
2 87792 1 7865
2 87793 1 7865
2 87794 1 7865
2 87795 1 7865
2 87796 1 7865
2 87797 1 7865
2 87798 1 7865
2 87799 1 7865
2 87800 1 7865
2 87801 1 7865
2 87802 1 7865
2 87803 1 7865
2 87804 1 7865
2 87805 1 7865
2 87806 1 7865
2 87807 1 7865
2 87808 1 7865
2 87809 1 7865
2 87810 1 7865
2 87811 1 7865
2 87812 1 7865
2 87813 1 7865
2 87814 1 7865
2 87815 1 7865
2 87816 1 7865
2 87817 1 7865
2 87818 1 7865
2 87819 1 7872
2 87820 1 7872
2 87821 1 7872
2 87822 1 7873
2 87823 1 7873
2 87824 1 7873
2 87825 1 7873
2 87826 1 7873
2 87827 1 7873
2 87828 1 7873
2 87829 1 7881
2 87830 1 7881
2 87831 1 7881
2 87832 1 7881
2 87833 1 7881
2 87834 1 7881
2 87835 1 7881
2 87836 1 7881
2 87837 1 7881
2 87838 1 7881
2 87839 1 7881
2 87840 1 7881
2 87841 1 7881
2 87842 1 7881
2 87843 1 7881
2 87844 1 7881
2 87845 1 7881
2 87846 1 7881
2 87847 1 7881
2 87848 1 7882
2 87849 1 7882
2 87850 1 7882
2 87851 1 7885
2 87852 1 7885
2 87853 1 7885
2 87854 1 7885
2 87855 1 7885
2 87856 1 7885
2 87857 1 7885
2 87858 1 7885
2 87859 1 7885
2 87860 1 7885
2 87861 1 7898
2 87862 1 7898
2 87863 1 7911
2 87864 1 7911
2 87865 1 7911
2 87866 1 7911
2 87867 1 7911
2 87868 1 7911
2 87869 1 7912
2 87870 1 7912
2 87871 1 7912
2 87872 1 7912
2 87873 1 7912
2 87874 1 7912
2 87875 1 7913
2 87876 1 7913
2 87877 1 7913
2 87878 1 7913
2 87879 1 7913
2 87880 1 7930
2 87881 1 7930
2 87882 1 7930
2 87883 1 7932
2 87884 1 7932
2 87885 1 7932
2 87886 1 7932
2 87887 1 7932
2 87888 1 7933
2 87889 1 7933
2 87890 1 7933
2 87891 1 7939
2 87892 1 7939
2 87893 1 7939
2 87894 1 7939
2 87895 1 7939
2 87896 1 7939
2 87897 1 7939
2 87898 1 7939
2 87899 1 7948
2 87900 1 7948
2 87901 1 7948
2 87902 1 7948
2 87903 1 7948
2 87904 1 7950
2 87905 1 7950
2 87906 1 7953
2 87907 1 7953
2 87908 1 7954
2 87909 1 7954
2 87910 1 7954
2 87911 1 7955
2 87912 1 7955
2 87913 1 7965
2 87914 1 7965
2 87915 1 7975
2 87916 1 7975
2 87917 1 7975
2 87918 1 7978
2 87919 1 7978
2 87920 1 7993
2 87921 1 7993
2 87922 1 7993
2 87923 1 7993
2 87924 1 7993
2 87925 1 7993
2 87926 1 7993
2 87927 1 7993
2 87928 1 7993
2 87929 1 7994
2 87930 1 7994
2 87931 1 7994
2 87932 1 7997
2 87933 1 7997
2 87934 1 7997
2 87935 1 7997
2 87936 1 7998
2 87937 1 7998
2 87938 1 7998
2 87939 1 7998
2 87940 1 7998
2 87941 1 7998
2 87942 1 7998
2 87943 1 7998
2 87944 1 7998
2 87945 1 8005
2 87946 1 8005
2 87947 1 8005
2 87948 1 8005
2 87949 1 8005
2 87950 1 8005
2 87951 1 8005
2 87952 1 8005
2 87953 1 8005
2 87954 1 8006
2 87955 1 8006
2 87956 1 8006
2 87957 1 8006
2 87958 1 8006
2 87959 1 8006
2 87960 1 8006
2 87961 1 8007
2 87962 1 8007
2 87963 1 8007
2 87964 1 8014
2 87965 1 8014
2 87966 1 8015
2 87967 1 8015
2 87968 1 8015
2 87969 1 8016
2 87970 1 8016
2 87971 1 8016
2 87972 1 8016
2 87973 1 8016
2 87974 1 8016
2 87975 1 8035
2 87976 1 8035
2 87977 1 8049
2 87978 1 8049
2 87979 1 8055
2 87980 1 8055
2 87981 1 8057
2 87982 1 8057
2 87983 1 8058
2 87984 1 8058
2 87985 1 8058
2 87986 1 8058
2 87987 1 8067
2 87988 1 8067
2 87989 1 8067
2 87990 1 8068
2 87991 1 8068
2 87992 1 8068
2 87993 1 8080
2 87994 1 8080
2 87995 1 8102
2 87996 1 8102
2 87997 1 8102
2 87998 1 8114
2 87999 1 8114
2 88000 1 8116
2 88001 1 8116
2 88002 1 8122
2 88003 1 8122
2 88004 1 8126
2 88005 1 8126
2 88006 1 8127
2 88007 1 8127
2 88008 1 8144
2 88009 1 8144
2 88010 1 8145
2 88011 1 8145
2 88012 1 8146
2 88013 1 8146
2 88014 1 8147
2 88015 1 8147
2 88016 1 8156
2 88017 1 8156
2 88018 1 8168
2 88019 1 8168
2 88020 1 8168
2 88021 1 8171
2 88022 1 8171
2 88023 1 8200
2 88024 1 8200
2 88025 1 8206
2 88026 1 8206
2 88027 1 8207
2 88028 1 8207
2 88029 1 8207
2 88030 1 8207
2 88031 1 8207
2 88032 1 8207
2 88033 1 8207
2 88034 1 8238
2 88035 1 8238
2 88036 1 8248
2 88037 1 8248
2 88038 1 8248
2 88039 1 8248
2 88040 1 8248
2 88041 1 8248
2 88042 1 8248
2 88043 1 8248
2 88044 1 8248
2 88045 1 8248
2 88046 1 8261
2 88047 1 8261
2 88048 1 8269
2 88049 1 8269
2 88050 1 8269
2 88051 1 8269
2 88052 1 8269
2 88053 1 8271
2 88054 1 8271
2 88055 1 8271
2 88056 1 8280
2 88057 1 8280
2 88058 1 8280
2 88059 1 8289
2 88060 1 8289
2 88061 1 8289
2 88062 1 8293
2 88063 1 8293
2 88064 1 8311
2 88065 1 8311
2 88066 1 8313
2 88067 1 8313
2 88068 1 8313
2 88069 1 8313
2 88070 1 8322
2 88071 1 8322
2 88072 1 8322
2 88073 1 8322
2 88074 1 8324
2 88075 1 8324
2 88076 1 8324
2 88077 1 8324
2 88078 1 8324
2 88079 1 8324
2 88080 1 8324
2 88081 1 8325
2 88082 1 8325
2 88083 1 8333
2 88084 1 8333
2 88085 1 8333
2 88086 1 8341
2 88087 1 8341
2 88088 1 8342
2 88089 1 8342
2 88090 1 8343
2 88091 1 8343
2 88092 1 8343
2 88093 1 8343
2 88094 1 8343
2 88095 1 8343
2 88096 1 8343
2 88097 1 8343
2 88098 1 8343
2 88099 1 8343
2 88100 1 8343
2 88101 1 8343
2 88102 1 8343
2 88103 1 8343
2 88104 1 8343
2 88105 1 8343
2 88106 1 8343
2 88107 1 8343
2 88108 1 8343
2 88109 1 8352
2 88110 1 8352
2 88111 1 8352
2 88112 1 8353
2 88113 1 8353
2 88114 1 8358
2 88115 1 8358
2 88116 1 8358
2 88117 1 8358
2 88118 1 8358
2 88119 1 8358
2 88120 1 8358
2 88121 1 8358
2 88122 1 8358
2 88123 1 8358
2 88124 1 8358
2 88125 1 8358
2 88126 1 8358
2 88127 1 8358
2 88128 1 8358
2 88129 1 8358
2 88130 1 8358
2 88131 1 8358
2 88132 1 8358
2 88133 1 8359
2 88134 1 8359
2 88135 1 8371
2 88136 1 8371
2 88137 1 8371
2 88138 1 8371
2 88139 1 8371
2 88140 1 8371
2 88141 1 8371
2 88142 1 8372
2 88143 1 8372
2 88144 1 8372
2 88145 1 8372
2 88146 1 8372
2 88147 1 8372
2 88148 1 8372
2 88149 1 8372
2 88150 1 8376
2 88151 1 8376
2 88152 1 8384
2 88153 1 8384
2 88154 1 8384
2 88155 1 8392
2 88156 1 8392
2 88157 1 8403
2 88158 1 8403
2 88159 1 8407
2 88160 1 8407
2 88161 1 8407
2 88162 1 8407
2 88163 1 8428
2 88164 1 8428
2 88165 1 8428
2 88166 1 8428
2 88167 1 8428
2 88168 1 8428
2 88169 1 8428
2 88170 1 8428
2 88171 1 8428
2 88172 1 8428
2 88173 1 8429
2 88174 1 8429
2 88175 1 8429
2 88176 1 8429
2 88177 1 8429
2 88178 1 8429
2 88179 1 8429
2 88180 1 8429
2 88181 1 8432
2 88182 1 8432
2 88183 1 8432
2 88184 1 8432
2 88185 1 8432
2 88186 1 8432
2 88187 1 8432
2 88188 1 8432
2 88189 1 8432
2 88190 1 8432
2 88191 1 8432
2 88192 1 8432
2 88193 1 8432
2 88194 1 8432
2 88195 1 8432
2 88196 1 8432
2 88197 1 8432
2 88198 1 8432
2 88199 1 8432
2 88200 1 8434
2 88201 1 8434
2 88202 1 8434
2 88203 1 8434
2 88204 1 8434
2 88205 1 8438
2 88206 1 8438
2 88207 1 8446
2 88208 1 8446
2 88209 1 8456
2 88210 1 8456
2 88211 1 8456
2 88212 1 8456
2 88213 1 8456
2 88214 1 8456
2 88215 1 8456
2 88216 1 8457
2 88217 1 8457
2 88218 1 8464
2 88219 1 8464
2 88220 1 8464
2 88221 1 8464
2 88222 1 8464
2 88223 1 8464
2 88224 1 8464
2 88225 1 8464
2 88226 1 8464
2 88227 1 8464
2 88228 1 8465
2 88229 1 8465
2 88230 1 8472
2 88231 1 8472
2 88232 1 8472
2 88233 1 8472
2 88234 1 8472
2 88235 1 8472
2 88236 1 8472
2 88237 1 8474
2 88238 1 8474
2 88239 1 8484
2 88240 1 8484
2 88241 1 8484
2 88242 1 8484
2 88243 1 8484
2 88244 1 8484
2 88245 1 8484
2 88246 1 8484
2 88247 1 8484
2 88248 1 8484
2 88249 1 8484
2 88250 1 8484
2 88251 1 8484
2 88252 1 8484
2 88253 1 8484
2 88254 1 8484
2 88255 1 8484
2 88256 1 8484
2 88257 1 8496
2 88258 1 8496
2 88259 1 8496
2 88260 1 8496
2 88261 1 8496
2 88262 1 8496
2 88263 1 8502
2 88264 1 8502
2 88265 1 8508
2 88266 1 8508
2 88267 1 8508
2 88268 1 8515
2 88269 1 8515
2 88270 1 8523
2 88271 1 8523
2 88272 1 8523
2 88273 1 8523
2 88274 1 8523
2 88275 1 8523
2 88276 1 8523
2 88277 1 8524
2 88278 1 8524
2 88279 1 8524
2 88280 1 8524
2 88281 1 8524
2 88282 1 8524
2 88283 1 8525
2 88284 1 8525
2 88285 1 8525
2 88286 1 8525
2 88287 1 8525
2 88288 1 8525
2 88289 1 8534
2 88290 1 8534
2 88291 1 8535
2 88292 1 8535
2 88293 1 8535
2 88294 1 8535
2 88295 1 8535
2 88296 1 8535
2 88297 1 8535
2 88298 1 8535
2 88299 1 8535
2 88300 1 8535
2 88301 1 8535
2 88302 1 8535
2 88303 1 8535
2 88304 1 8552
2 88305 1 8552
2 88306 1 8552
2 88307 1 8553
2 88308 1 8553
2 88309 1 8560
2 88310 1 8560
2 88311 1 8564
2 88312 1 8564
2 88313 1 8567
2 88314 1 8567
2 88315 1 8581
2 88316 1 8581
2 88317 1 8581
2 88318 1 8581
2 88319 1 8582
2 88320 1 8582
2 88321 1 8583
2 88322 1 8583
2 88323 1 8583
2 88324 1 8583
2 88325 1 8584
2 88326 1 8584
2 88327 1 8605
2 88328 1 8605
2 88329 1 8605
2 88330 1 8608
2 88331 1 8608
2 88332 1 8608
2 88333 1 8608
2 88334 1 8609
2 88335 1 8609
2 88336 1 8609
2 88337 1 8609
2 88338 1 8610
2 88339 1 8610
2 88340 1 8621
2 88341 1 8621
2 88342 1 8622
2 88343 1 8622
2 88344 1 8632
2 88345 1 8632
2 88346 1 8645
2 88347 1 8645
2 88348 1 8645
2 88349 1 8645
2 88350 1 8645
2 88351 1 8645
2 88352 1 8645
2 88353 1 8646
2 88354 1 8646
2 88355 1 8647
2 88356 1 8647
2 88357 1 8647
2 88358 1 8647
2 88359 1 8648
2 88360 1 8648
2 88361 1 8651
2 88362 1 8651
2 88363 1 8666
2 88364 1 8666
2 88365 1 8669
2 88366 1 8669
2 88367 1 8669
2 88368 1 8669
2 88369 1 8669
2 88370 1 8669
2 88371 1 8669
2 88372 1 8672
2 88373 1 8672
2 88374 1 8673
2 88375 1 8673
2 88376 1 8673
2 88377 1 8674
2 88378 1 8674
2 88379 1 8674
2 88380 1 8674
2 88381 1 8674
2 88382 1 8674
2 88383 1 8674
2 88384 1 8674
2 88385 1 8684
2 88386 1 8684
2 88387 1 8684
2 88388 1 8687
2 88389 1 8687
2 88390 1 8687
2 88391 1 8688
2 88392 1 8688
2 88393 1 8689
2 88394 1 8689
2 88395 1 8689
2 88396 1 8702
2 88397 1 8702
2 88398 1 8702
2 88399 1 8703
2 88400 1 8703
2 88401 1 8706
2 88402 1 8706
2 88403 1 8706
2 88404 1 8707
2 88405 1 8707
2 88406 1 8721
2 88407 1 8721
2 88408 1 8722
2 88409 1 8722
2 88410 1 8722
2 88411 1 8735
2 88412 1 8735
2 88413 1 8735
2 88414 1 8735
2 88415 1 8735
2 88416 1 8737
2 88417 1 8737
2 88418 1 8737
2 88419 1 8737
2 88420 1 8737
2 88421 1 8737
2 88422 1 8737
2 88423 1 8737
2 88424 1 8737
2 88425 1 8737
2 88426 1 8737
2 88427 1 8738
2 88428 1 8738
2 88429 1 8740
2 88430 1 8740
2 88431 1 8745
2 88432 1 8745
2 88433 1 8750
2 88434 1 8750
2 88435 1 8759
2 88436 1 8759
2 88437 1 8760
2 88438 1 8760
2 88439 1 8760
2 88440 1 8760
2 88441 1 8761
2 88442 1 8761
2 88443 1 8762
2 88444 1 8762
2 88445 1 8762
2 88446 1 8762
2 88447 1 8772
2 88448 1 8772
2 88449 1 8772
2 88450 1 8772
2 88451 1 8772
2 88452 1 8772
2 88453 1 8781
2 88454 1 8781
2 88455 1 8794
2 88456 1 8794
2 88457 1 8794
2 88458 1 8795
2 88459 1 8795
2 88460 1 8795
2 88461 1 8795
2 88462 1 8795
2 88463 1 8795
2 88464 1 8795
2 88465 1 8795
2 88466 1 8795
2 88467 1 8795
2 88468 1 8795
2 88469 1 8795
2 88470 1 8795
2 88471 1 8795
2 88472 1 8795
2 88473 1 8805
2 88474 1 8805
2 88475 1 8806
2 88476 1 8806
2 88477 1 8806
2 88478 1 8809
2 88479 1 8809
2 88480 1 8814
2 88481 1 8814
2 88482 1 8814
2 88483 1 8818
2 88484 1 8818
2 88485 1 8821
2 88486 1 8821
2 88487 1 8827
2 88488 1 8827
2 88489 1 8833
2 88490 1 8833
2 88491 1 8833
2 88492 1 8833
2 88493 1 8833
2 88494 1 8833
2 88495 1 8833
2 88496 1 8834
2 88497 1 8834
2 88498 1 8834
2 88499 1 8834
2 88500 1 8835
2 88501 1 8835
2 88502 1 8835
2 88503 1 8835
2 88504 1 8835
2 88505 1 8835
2 88506 1 8835
2 88507 1 8835
2 88508 1 8835
2 88509 1 8835
2 88510 1 8835
2 88511 1 8835
2 88512 1 8835
2 88513 1 8835
2 88514 1 8835
2 88515 1 8835
2 88516 1 8835
2 88517 1 8836
2 88518 1 8836
2 88519 1 8838
2 88520 1 8838
2 88521 1 8839
2 88522 1 8839
2 88523 1 8839
2 88524 1 8839
2 88525 1 8856
2 88526 1 8856
2 88527 1 8857
2 88528 1 8857
2 88529 1 8857
2 88530 1 8857
2 88531 1 8857
2 88532 1 8857
2 88533 1 8857
2 88534 1 8857
2 88535 1 8857
2 88536 1 8857
2 88537 1 8857
2 88538 1 8857
2 88539 1 8857
2 88540 1 8858
2 88541 1 8858
2 88542 1 8858
2 88543 1 8858
2 88544 1 8859
2 88545 1 8859
2 88546 1 8859
2 88547 1 8860
2 88548 1 8860
2 88549 1 8861
2 88550 1 8861
2 88551 1 8861
2 88552 1 8861
2 88553 1 8861
2 88554 1 8869
2 88555 1 8869
2 88556 1 8869
2 88557 1 8869
2 88558 1 8870
2 88559 1 8870
2 88560 1 8870
2 88561 1 8870
2 88562 1 8870
2 88563 1 8889
2 88564 1 8889
2 88565 1 8906
2 88566 1 8906
2 88567 1 8906
2 88568 1 8906
2 88569 1 8907
2 88570 1 8907
2 88571 1 8916
2 88572 1 8916
2 88573 1 8924
2 88574 1 8924
2 88575 1 8924
2 88576 1 8924
2 88577 1 8928
2 88578 1 8928
2 88579 1 8937
2 88580 1 8937
2 88581 1 8937
2 88582 1 8938
2 88583 1 8938
2 88584 1 8941
2 88585 1 8941
2 88586 1 8952
2 88587 1 8952
2 88588 1 8952
2 88589 1 8952
2 88590 1 8952
2 88591 1 8952
2 88592 1 8953
2 88593 1 8953
2 88594 1 8963
2 88595 1 8963
2 88596 1 8966
2 88597 1 8966
2 88598 1 8966
2 88599 1 8974
2 88600 1 8974
2 88601 1 8979
2 88602 1 8979
2 88603 1 8982
2 88604 1 8982
2 88605 1 8983
2 88606 1 8983
2 88607 1 8983
2 88608 1 8983
2 88609 1 8984
2 88610 1 8984
2 88611 1 8990
2 88612 1 8990
2 88613 1 9002
2 88614 1 9002
2 88615 1 9006
2 88616 1 9006
2 88617 1 9006
2 88618 1 9006
2 88619 1 9008
2 88620 1 9008
2 88621 1 9008
2 88622 1 9008
2 88623 1 9008
2 88624 1 9008
2 88625 1 9008
2 88626 1 9008
2 88627 1 9008
2 88628 1 9022
2 88629 1 9022
2 88630 1 9027
2 88631 1 9027
2 88632 1 9027
2 88633 1 9027
2 88634 1 9030
2 88635 1 9030
2 88636 1 9030
2 88637 1 9030
2 88638 1 9030
2 88639 1 9030
2 88640 1 9030
2 88641 1 9030
2 88642 1 9030
2 88643 1 9037
2 88644 1 9037
2 88645 1 9037
2 88646 1 9052
2 88647 1 9052
2 88648 1 9052
2 88649 1 9052
2 88650 1 9052
2 88651 1 9053
2 88652 1 9053
2 88653 1 9062
2 88654 1 9062
2 88655 1 9062
2 88656 1 9062
2 88657 1 9063
2 88658 1 9063
2 88659 1 9075
2 88660 1 9075
2 88661 1 9088
2 88662 1 9088
2 88663 1 9095
2 88664 1 9095
2 88665 1 9095
2 88666 1 9095
2 88667 1 9095
2 88668 1 9095
2 88669 1 9095
2 88670 1 9095
2 88671 1 9095
2 88672 1 9095
2 88673 1 9095
2 88674 1 9095
2 88675 1 9095
2 88676 1 9095
2 88677 1 9095
2 88678 1 9095
2 88679 1 9104
2 88680 1 9104
2 88681 1 9104
2 88682 1 9104
2 88683 1 9112
2 88684 1 9112
2 88685 1 9112
2 88686 1 9112
2 88687 1 9112
2 88688 1 9112
2 88689 1 9112
2 88690 1 9112
2 88691 1 9113
2 88692 1 9113
2 88693 1 9113
2 88694 1 9114
2 88695 1 9114
2 88696 1 9114
2 88697 1 9114
2 88698 1 9114
2 88699 1 9114
2 88700 1 9115
2 88701 1 9115
2 88702 1 9123
2 88703 1 9123
2 88704 1 9123
2 88705 1 9123
2 88706 1 9123
2 88707 1 9125
2 88708 1 9125
2 88709 1 9125
2 88710 1 9125
2 88711 1 9135
2 88712 1 9135
2 88713 1 9135
2 88714 1 9135
2 88715 1 9135
2 88716 1 9135
2 88717 1 9136
2 88718 1 9136
2 88719 1 9136
2 88720 1 9136
2 88721 1 9136
2 88722 1 9143
2 88723 1 9143
2 88724 1 9143
2 88725 1 9143
2 88726 1 9146
2 88727 1 9146
2 88728 1 9152
2 88729 1 9152
2 88730 1 9152
2 88731 1 9152
2 88732 1 9152
2 88733 1 9152
2 88734 1 9152
2 88735 1 9152
2 88736 1 9152
2 88737 1 9152
2 88738 1 9152
2 88739 1 9153
2 88740 1 9153
2 88741 1 9176
2 88742 1 9176
2 88743 1 9177
2 88744 1 9177
2 88745 1 9178
2 88746 1 9178
2 88747 1 9178
2 88748 1 9178
2 88749 1 9178
2 88750 1 9188
2 88751 1 9188
2 88752 1 9188
2 88753 1 9190
2 88754 1 9190
2 88755 1 9190
2 88756 1 9190
2 88757 1 9190
2 88758 1 9190
2 88759 1 9190
2 88760 1 9190
2 88761 1 9191
2 88762 1 9191
2 88763 1 9227
2 88764 1 9227
2 88765 1 9227
2 88766 1 9227
2 88767 1 9227
2 88768 1 9227
2 88769 1 9227
2 88770 1 9227
2 88771 1 9227
2 88772 1 9227
2 88773 1 9227
2 88774 1 9239
2 88775 1 9239
2 88776 1 9239
2 88777 1 9239
2 88778 1 9239
2 88779 1 9242
2 88780 1 9242
2 88781 1 9242
2 88782 1 9254
2 88783 1 9254
2 88784 1 9254
2 88785 1 9254
2 88786 1 9254
2 88787 1 9264
2 88788 1 9264
2 88789 1 9264
2 88790 1 9264
2 88791 1 9276
2 88792 1 9276
2 88793 1 9276
2 88794 1 9285
2 88795 1 9285
2 88796 1 9285
2 88797 1 9285
2 88798 1 9285
2 88799 1 9285
2 88800 1 9285
2 88801 1 9308
2 88802 1 9308
2 88803 1 9319
2 88804 1 9319
2 88805 1 9320
2 88806 1 9320
2 88807 1 9320
2 88808 1 9320
2 88809 1 9323
2 88810 1 9323
2 88811 1 9323
2 88812 1 9331
2 88813 1 9331
2 88814 1 9331
2 88815 1 9331
2 88816 1 9332
2 88817 1 9332
2 88818 1 9332
2 88819 1 9332
2 88820 1 9332
2 88821 1 9332
2 88822 1 9332
2 88823 1 9332
2 88824 1 9332
2 88825 1 9341
2 88826 1 9341
2 88827 1 9341
2 88828 1 9341
2 88829 1 9341
2 88830 1 9341
2 88831 1 9342
2 88832 1 9342
2 88833 1 9347
2 88834 1 9347
2 88835 1 9347
2 88836 1 9355
2 88837 1 9355
2 88838 1 9355
2 88839 1 9355
2 88840 1 9409
2 88841 1 9409
2 88842 1 9409
2 88843 1 9417
2 88844 1 9417
2 88845 1 9426
2 88846 1 9426
2 88847 1 9429
2 88848 1 9429
2 88849 1 9429
2 88850 1 9430
2 88851 1 9430
2 88852 1 9430
2 88853 1 9430
2 88854 1 9430
2 88855 1 9430
2 88856 1 9430
2 88857 1 9430
2 88858 1 9430
2 88859 1 9431
2 88860 1 9431
2 88861 1 9433
2 88862 1 9433
2 88863 1 9433
2 88864 1 9437
2 88865 1 9437
2 88866 1 9439
2 88867 1 9439
2 88868 1 9439
2 88869 1 9439
2 88870 1 9452
2 88871 1 9452
2 88872 1 9452
2 88873 1 9452
2 88874 1 9452
2 88875 1 9452
2 88876 1 9452
2 88877 1 9452
2 88878 1 9452
2 88879 1 9452
2 88880 1 9458
2 88881 1 9458
2 88882 1 9474
2 88883 1 9474
2 88884 1 9475
2 88885 1 9475
2 88886 1 9476
2 88887 1 9476
2 88888 1 9476
2 88889 1 9476
2 88890 1 9477
2 88891 1 9477
2 88892 1 9477
2 88893 1 9491
2 88894 1 9491
2 88895 1 9499
2 88896 1 9499
2 88897 1 9499
2 88898 1 9499
2 88899 1 9499
2 88900 1 9499
2 88901 1 9499
2 88902 1 9499
2 88903 1 9499
2 88904 1 9500
2 88905 1 9500
2 88906 1 9500
2 88907 1 9503
2 88908 1 9503
2 88909 1 9510
2 88910 1 9510
2 88911 1 9510
2 88912 1 9510
2 88913 1 9510
2 88914 1 9510
2 88915 1 9510
2 88916 1 9510
2 88917 1 9510
2 88918 1 9510
2 88919 1 9510
2 88920 1 9510
2 88921 1 9510
2 88922 1 9510
2 88923 1 9518
2 88924 1 9518
2 88925 1 9518
2 88926 1 9526
2 88927 1 9526
2 88928 1 9541
2 88929 1 9541
2 88930 1 9541
2 88931 1 9541
2 88932 1 9546
2 88933 1 9546
2 88934 1 9546
2 88935 1 9546
2 88936 1 9546
2 88937 1 9554
2 88938 1 9554
2 88939 1 9554
2 88940 1 9554
2 88941 1 9554
2 88942 1 9554
2 88943 1 9554
2 88944 1 9554
2 88945 1 9554
2 88946 1 9554
2 88947 1 9554
2 88948 1 9554
2 88949 1 9554
2 88950 1 9554
2 88951 1 9554
2 88952 1 9554
2 88953 1 9554
2 88954 1 9554
2 88955 1 9554
2 88956 1 9554
2 88957 1 9554
2 88958 1 9558
2 88959 1 9558
2 88960 1 9570
2 88961 1 9570
2 88962 1 9578
2 88963 1 9578
2 88964 1 9578
2 88965 1 9578
2 88966 1 9578
2 88967 1 9578
2 88968 1 9578
2 88969 1 9578
2 88970 1 9578
2 88971 1 9578
2 88972 1 9578
2 88973 1 9578
2 88974 1 9578
2 88975 1 9578
2 88976 1 9578
2 88977 1 9578
2 88978 1 9578
2 88979 1 9578
2 88980 1 9578
2 88981 1 9579
2 88982 1 9579
2 88983 1 9579
2 88984 1 9579
2 88985 1 9580
2 88986 1 9580
2 88987 1 9580
2 88988 1 9592
2 88989 1 9592
2 88990 1 9594
2 88991 1 9594
2 88992 1 9600
2 88993 1 9600
2 88994 1 9600
2 88995 1 9604
2 88996 1 9604
2 88997 1 9604
2 88998 1 9604
2 88999 1 9604
2 89000 1 9604
2 89001 1 9604
2 89002 1 9604
2 89003 1 9604
2 89004 1 9612
2 89005 1 9612
2 89006 1 9618
2 89007 1 9618
2 89008 1 9621
2 89009 1 9621
2 89010 1 9621
2 89011 1 9621
2 89012 1 9630
2 89013 1 9630
2 89014 1 9630
2 89015 1 9630
2 89016 1 9645
2 89017 1 9645
2 89018 1 9645
2 89019 1 9645
2 89020 1 9653
2 89021 1 9653
2 89022 1 9653
2 89023 1 9653
2 89024 1 9654
2 89025 1 9654
2 89026 1 9654
2 89027 1 9654
2 89028 1 9656
2 89029 1 9656
2 89030 1 9672
2 89031 1 9672
2 89032 1 9680
2 89033 1 9680
2 89034 1 9681
2 89035 1 9681
2 89036 1 9682
2 89037 1 9682
2 89038 1 9683
2 89039 1 9683
2 89040 1 9691
2 89041 1 9691
2 89042 1 9692
2 89043 1 9692
2 89044 1 9701
2 89045 1 9701
2 89046 1 9708
2 89047 1 9708
2 89048 1 9709
2 89049 1 9709
2 89050 1 9710
2 89051 1 9710
2 89052 1 9714
2 89053 1 9714
2 89054 1 9714
2 89055 1 9721
2 89056 1 9721
2 89057 1 9721
2 89058 1 9721
2 89059 1 9721
2 89060 1 9722
2 89061 1 9722
2 89062 1 9722
2 89063 1 9722
2 89064 1 9723
2 89065 1 9723
2 89066 1 9726
2 89067 1 9726
2 89068 1 9726
2 89069 1 9726
2 89070 1 9727
2 89071 1 9727
2 89072 1 9727
2 89073 1 9730
2 89074 1 9730
2 89075 1 9730
2 89076 1 9737
2 89077 1 9737
2 89078 1 9737
2 89079 1 9737
2 89080 1 9737
2 89081 1 9737
2 89082 1 9737
2 89083 1 9737
2 89084 1 9737
2 89085 1 9737
2 89086 1 9737
2 89087 1 9737
2 89088 1 9737
2 89089 1 9737
2 89090 1 9737
2 89091 1 9738
2 89092 1 9738
2 89093 1 9769
2 89094 1 9769
2 89095 1 9769
2 89096 1 9784
2 89097 1 9784
2 89098 1 9792
2 89099 1 9792
2 89100 1 9811
2 89101 1 9811
2 89102 1 9825
2 89103 1 9825
2 89104 1 9825
2 89105 1 9825
2 89106 1 9825
2 89107 1 9825
2 89108 1 9825
2 89109 1 9825
2 89110 1 9825
2 89111 1 9825
2 89112 1 9825
2 89113 1 9825
2 89114 1 9828
2 89115 1 9828
2 89116 1 9838
2 89117 1 9838
2 89118 1 9838
2 89119 1 9839
2 89120 1 9839
2 89121 1 9839
2 89122 1 9839
2 89123 1 9839
2 89124 1 9856
2 89125 1 9856
2 89126 1 9864
2 89127 1 9864
2 89128 1 9872
2 89129 1 9872
2 89130 1 9874
2 89131 1 9874
2 89132 1 9874
2 89133 1 9874
2 89134 1 9874
2 89135 1 9888
2 89136 1 9888
2 89137 1 9888
2 89138 1 9893
2 89139 1 9893
2 89140 1 9894
2 89141 1 9894
2 89142 1 9914
2 89143 1 9914
2 89144 1 9914
2 89145 1 9917
2 89146 1 9917
2 89147 1 9918
2 89148 1 9918
2 89149 1 9918
2 89150 1 9932
2 89151 1 9932
2 89152 1 9942
2 89153 1 9942
2 89154 1 9984
2 89155 1 9984
2 89156 1 9985
2 89157 1 9985
2 89158 1 10008
2 89159 1 10008
2 89160 1 10008
2 89161 1 10008
2 89162 1 10008
2 89163 1 10008
2 89164 1 10008
2 89165 1 10008
2 89166 1 10008
2 89167 1 10008
2 89168 1 10008
2 89169 1 10008
2 89170 1 10008
2 89171 1 10008
2 89172 1 10010
2 89173 1 10010
2 89174 1 10011
2 89175 1 10011
2 89176 1 10020
2 89177 1 10020
2 89178 1 10020
2 89179 1 10021
2 89180 1 10021
2 89181 1 10021
2 89182 1 10021
2 89183 1 10021
2 89184 1 10035
2 89185 1 10035
2 89186 1 10035
2 89187 1 10035
2 89188 1 10038
2 89189 1 10038
2 89190 1 10045
2 89191 1 10045
2 89192 1 10052
2 89193 1 10052
2 89194 1 10053
2 89195 1 10053
2 89196 1 10060
2 89197 1 10060
2 89198 1 10062
2 89199 1 10062
2 89200 1 10062
2 89201 1 10062
2 89202 1 10062
2 89203 1 10062
2 89204 1 10062
2 89205 1 10070
2 89206 1 10070
2 89207 1 10070
2 89208 1 10070
2 89209 1 10070
2 89210 1 10070
2 89211 1 10070
2 89212 1 10078
2 89213 1 10078
2 89214 1 10078
2 89215 1 10078
2 89216 1 10079
2 89217 1 10079
2 89218 1 10090
2 89219 1 10090
2 89220 1 10091
2 89221 1 10091
2 89222 1 10092
2 89223 1 10092
2 89224 1 10101
2 89225 1 10101
2 89226 1 10101
2 89227 1 10122
2 89228 1 10122
2 89229 1 10133
2 89230 1 10133
2 89231 1 10133
2 89232 1 10133
2 89233 1 10133
2 89234 1 10136
2 89235 1 10136
2 89236 1 10136
2 89237 1 10141
2 89238 1 10141
2 89239 1 10158
2 89240 1 10158
2 89241 1 10158
2 89242 1 10161
2 89243 1 10161
2 89244 1 10184
2 89245 1 10184
2 89246 1 10186
2 89247 1 10186
2 89248 1 10218
2 89249 1 10218
2 89250 1 10218
2 89251 1 10218
2 89252 1 10221
2 89253 1 10221
2 89254 1 10221
2 89255 1 10235
2 89256 1 10235
2 89257 1 10235
2 89258 1 10235
2 89259 1 10235
2 89260 1 10235
2 89261 1 10235
2 89262 1 10235
2 89263 1 10235
2 89264 1 10235
2 89265 1 10235
2 89266 1 10235
2 89267 1 10235
2 89268 1 10235
2 89269 1 10235
2 89270 1 10235
2 89271 1 10235
2 89272 1 10235
2 89273 1 10235
2 89274 1 10235
2 89275 1 10235
2 89276 1 10236
2 89277 1 10236
2 89278 1 10237
2 89279 1 10237
2 89280 1 10242
2 89281 1 10242
2 89282 1 10242
2 89283 1 10242
2 89284 1 10242
2 89285 1 10242
2 89286 1 10242
2 89287 1 10242
2 89288 1 10242
2 89289 1 10243
2 89290 1 10243
2 89291 1 10243
2 89292 1 10243
2 89293 1 10251
2 89294 1 10251
2 89295 1 10251
2 89296 1 10252
2 89297 1 10252
2 89298 1 10252
2 89299 1 10252
2 89300 1 10252
2 89301 1 10252
2 89302 1 10252
2 89303 1 10252
2 89304 1 10252
2 89305 1 10252
2 89306 1 10252
2 89307 1 10252
2 89308 1 10255
2 89309 1 10255
2 89310 1 10255
2 89311 1 10255
2 89312 1 10256
2 89313 1 10256
2 89314 1 10275
2 89315 1 10275
2 89316 1 10276
2 89317 1 10276
2 89318 1 10276
2 89319 1 10280
2 89320 1 10280
2 89321 1 10292
2 89322 1 10292
2 89323 1 10305
2 89324 1 10305
2 89325 1 10305
2 89326 1 10306
2 89327 1 10306
2 89328 1 10314
2 89329 1 10314
2 89330 1 10314
2 89331 1 10314
2 89332 1 10326
2 89333 1 10326
2 89334 1 10330
2 89335 1 10330
2 89336 1 10330
2 89337 1 10330
2 89338 1 10330
2 89339 1 10338
2 89340 1 10338
2 89341 1 10357
2 89342 1 10357
2 89343 1 10364
2 89344 1 10364
2 89345 1 10364
2 89346 1 10364
2 89347 1 10364
2 89348 1 10364
2 89349 1 10368
2 89350 1 10368
2 89351 1 10371
2 89352 1 10371
2 89353 1 10371
2 89354 1 10372
2 89355 1 10372
2 89356 1 10373
2 89357 1 10373
2 89358 1 10373
2 89359 1 10381
2 89360 1 10381
2 89361 1 10381
2 89362 1 10381
2 89363 1 10381
2 89364 1 10381
2 89365 1 10381
2 89366 1 10381
2 89367 1 10382
2 89368 1 10382
2 89369 1 10382
2 89370 1 10382
2 89371 1 10387
2 89372 1 10387
2 89373 1 10409
2 89374 1 10409
2 89375 1 10409
2 89376 1 10410
2 89377 1 10410
2 89378 1 10410
2 89379 1 10423
2 89380 1 10423
2 89381 1 10423
2 89382 1 10423
2 89383 1 10423
2 89384 1 10423
2 89385 1 10431
2 89386 1 10431
2 89387 1 10441
2 89388 1 10441
2 89389 1 10442
2 89390 1 10442
2 89391 1 10443
2 89392 1 10443
2 89393 1 10443
2 89394 1 10443
2 89395 1 10444
2 89396 1 10444
2 89397 1 10466
2 89398 1 10466
2 89399 1 10466
2 89400 1 10489
2 89401 1 10489
2 89402 1 10490
2 89403 1 10490
2 89404 1 10490
2 89405 1 10497
2 89406 1 10497
2 89407 1 10497
2 89408 1 10498
2 89409 1 10498
2 89410 1 10498
2 89411 1 10498
2 89412 1 10505
2 89413 1 10505
2 89414 1 10516
2 89415 1 10516
2 89416 1 10531
2 89417 1 10531
2 89418 1 10531
2 89419 1 10533
2 89420 1 10533
2 89421 1 10541
2 89422 1 10541
2 89423 1 10556
2 89424 1 10556
2 89425 1 10556
2 89426 1 10559
2 89427 1 10559
2 89428 1 10559
2 89429 1 10559
2 89430 1 10559
2 89431 1 10560
2 89432 1 10560
2 89433 1 10560
2 89434 1 10570
2 89435 1 10570
2 89436 1 10570
2 89437 1 10570
2 89438 1 10573
2 89439 1 10573
2 89440 1 10583
2 89441 1 10583
2 89442 1 10583
2 89443 1 10583
2 89444 1 10583
2 89445 1 10583
2 89446 1 10592
2 89447 1 10592
2 89448 1 10593
2 89449 1 10593
2 89450 1 10595
2 89451 1 10595
2 89452 1 10609
2 89453 1 10609
2 89454 1 10609
2 89455 1 10609
2 89456 1 10609
2 89457 1 10621
2 89458 1 10621
2 89459 1 10621
2 89460 1 10621
2 89461 1 10621
2 89462 1 10623
2 89463 1 10623
2 89464 1 10629
2 89465 1 10629
2 89466 1 10629
2 89467 1 10629
2 89468 1 10629
2 89469 1 10629
2 89470 1 10630
2 89471 1 10630
2 89472 1 10630
2 89473 1 10630
2 89474 1 10630
2 89475 1 10630
2 89476 1 10632
2 89477 1 10632
2 89478 1 10633
2 89479 1 10633
2 89480 1 10633
2 89481 1 10633
2 89482 1 10633
2 89483 1 10633
2 89484 1 10633
2 89485 1 10633
2 89486 1 10634
2 89487 1 10634
2 89488 1 10640
2 89489 1 10640
2 89490 1 10640
2 89491 1 10640
2 89492 1 10643
2 89493 1 10643
2 89494 1 10653
2 89495 1 10653
2 89496 1 10653
2 89497 1 10653
2 89498 1 10653
2 89499 1 10653
2 89500 1 10653
2 89501 1 10653
2 89502 1 10653
2 89503 1 10653
2 89504 1 10654
2 89505 1 10654
2 89506 1 10654
2 89507 1 10654
2 89508 1 10654
2 89509 1 10654
2 89510 1 10654
2 89511 1 10654
2 89512 1 10654
2 89513 1 10654
2 89514 1 10654
2 89515 1 10654
2 89516 1 10654
2 89517 1 10654
2 89518 1 10654
2 89519 1 10654
2 89520 1 10654
2 89521 1 10654
2 89522 1 10654
2 89523 1 10654
2 89524 1 10654
2 89525 1 10654
2 89526 1 10655
2 89527 1 10655
2 89528 1 10655
2 89529 1 10664
2 89530 1 10664
2 89531 1 10664
2 89532 1 10665
2 89533 1 10665
2 89534 1 10691
2 89535 1 10691
2 89536 1 10691
2 89537 1 10691
2 89538 1 10692
2 89539 1 10692
2 89540 1 10692
2 89541 1 10693
2 89542 1 10693
2 89543 1 10723
2 89544 1 10723
2 89545 1 10732
2 89546 1 10732
2 89547 1 10738
2 89548 1 10738
2 89549 1 10738
2 89550 1 10738
2 89551 1 10738
2 89552 1 10752
2 89553 1 10752
2 89554 1 10752
2 89555 1 10753
2 89556 1 10753
2 89557 1 10753
2 89558 1 10754
2 89559 1 10754
2 89560 1 10756
2 89561 1 10756
2 89562 1 10756
2 89563 1 10756
2 89564 1 10756
2 89565 1 10756
2 89566 1 10756
2 89567 1 10761
2 89568 1 10761
2 89569 1 10761
2 89570 1 10761
2 89571 1 10761
2 89572 1 10761
2 89573 1 10770
2 89574 1 10770
2 89575 1 10770
2 89576 1 10770
2 89577 1 10770
2 89578 1 10771
2 89579 1 10771
2 89580 1 10771
2 89581 1 10771
2 89582 1 10787
2 89583 1 10787
2 89584 1 10802
2 89585 1 10802
2 89586 1 10811
2 89587 1 10811
2 89588 1 10811
2 89589 1 10812
2 89590 1 10812
2 89591 1 10814
2 89592 1 10814
2 89593 1 10815
2 89594 1 10815
2 89595 1 10815
2 89596 1 10815
2 89597 1 10815
2 89598 1 10815
2 89599 1 10815
2 89600 1 10816
2 89601 1 10816
2 89602 1 10824
2 89603 1 10824
2 89604 1 10827
2 89605 1 10827
2 89606 1 10837
2 89607 1 10837
2 89608 1 10837
2 89609 1 10845
2 89610 1 10845
2 89611 1 10846
2 89612 1 10846
2 89613 1 10851
2 89614 1 10851
2 89615 1 10853
2 89616 1 10853
2 89617 1 10853
2 89618 1 10877
2 89619 1 10877
2 89620 1 10877
2 89621 1 10884
2 89622 1 10884
2 89623 1 10884
2 89624 1 10884
2 89625 1 10887
2 89626 1 10887
2 89627 1 10893
2 89628 1 10893
2 89629 1 10902
2 89630 1 10902
2 89631 1 10902
2 89632 1 10902
2 89633 1 10903
2 89634 1 10903
2 89635 1 10904
2 89636 1 10904
2 89637 1 10904
2 89638 1 10904
2 89639 1 10919
2 89640 1 10919
2 89641 1 10919
2 89642 1 10920
2 89643 1 10920
2 89644 1 10921
2 89645 1 10921
2 89646 1 10927
2 89647 1 10927
2 89648 1 10928
2 89649 1 10928
2 89650 1 10928
2 89651 1 10928
2 89652 1 10928
2 89653 1 10928
2 89654 1 10940
2 89655 1 10940
2 89656 1 10944
2 89657 1 10944
2 89658 1 10963
2 89659 1 10963
2 89660 1 10971
2 89661 1 10971
2 89662 1 10980
2 89663 1 10980
2 89664 1 10981
2 89665 1 10981
2 89666 1 10982
2 89667 1 10982
2 89668 1 10982
2 89669 1 10982
2 89670 1 10982
2 89671 1 10982
2 89672 1 10982
2 89673 1 10982
2 89674 1 10983
2 89675 1 10983
2 89676 1 10998
2 89677 1 10998
2 89678 1 11001
2 89679 1 11001
2 89680 1 11001
2 89681 1 11009
2 89682 1 11009
2 89683 1 11019
2 89684 1 11019
2 89685 1 11024
2 89686 1 11024
2 89687 1 11024
2 89688 1 11037
2 89689 1 11037
2 89690 1 11054
2 89691 1 11054
2 89692 1 11061
2 89693 1 11061
2 89694 1 11073
2 89695 1 11073
2 89696 1 11073
2 89697 1 11073
2 89698 1 11074
2 89699 1 11074
2 89700 1 11075
2 89701 1 11075
2 89702 1 11075
2 89703 1 11075
2 89704 1 11075
2 89705 1 11075
2 89706 1 11079
2 89707 1 11079
2 89708 1 11080
2 89709 1 11080
2 89710 1 11100
2 89711 1 11100
2 89712 1 11100
2 89713 1 11101
2 89714 1 11101
2 89715 1 11105
2 89716 1 11105
2 89717 1 11111
2 89718 1 11111
2 89719 1 11111
2 89720 1 11111
2 89721 1 11111
2 89722 1 11111
2 89723 1 11111
2 89724 1 11111
2 89725 1 11111
2 89726 1 11111
2 89727 1 11121
2 89728 1 11121
2 89729 1 11127
2 89730 1 11127
2 89731 1 11127
2 89732 1 11128
2 89733 1 11128
2 89734 1 11128
2 89735 1 11128
2 89736 1 11139
2 89737 1 11139
2 89738 1 11139
2 89739 1 11147
2 89740 1 11147
2 89741 1 11170
2 89742 1 11170
2 89743 1 11170
2 89744 1 11180
2 89745 1 11180
2 89746 1 11180
2 89747 1 11182
2 89748 1 11182
2 89749 1 11182
2 89750 1 11201
2 89751 1 11201
2 89752 1 11210
2 89753 1 11210
2 89754 1 11210
2 89755 1 11226
2 89756 1 11226
2 89757 1 11226
2 89758 1 11234
2 89759 1 11234
2 89760 1 11234
2 89761 1 11234
2 89762 1 11234
2 89763 1 11250
2 89764 1 11250
2 89765 1 11251
2 89766 1 11251
2 89767 1 11265
2 89768 1 11265
2 89769 1 11265
2 89770 1 11265
2 89771 1 11269
2 89772 1 11269
2 89773 1 11275
2 89774 1 11275
2 89775 1 11282
2 89776 1 11282
2 89777 1 11282
2 89778 1 11282
2 89779 1 11282
2 89780 1 11282
2 89781 1 11282
2 89782 1 11282
2 89783 1 11282
2 89784 1 11282
2 89785 1 11284
2 89786 1 11284
2 89787 1 11292
2 89788 1 11292
2 89789 1 11293
2 89790 1 11293
2 89791 1 11293
2 89792 1 11294
2 89793 1 11294
2 89794 1 11294
2 89795 1 11294
2 89796 1 11308
2 89797 1 11308
2 89798 1 11310
2 89799 1 11310
2 89800 1 11312
2 89801 1 11312
2 89802 1 11318
2 89803 1 11318
2 89804 1 11319
2 89805 1 11319
2 89806 1 11319
2 89807 1 11331
2 89808 1 11331
2 89809 1 11331
2 89810 1 11332
2 89811 1 11332
2 89812 1 11332
2 89813 1 11332
2 89814 1 11338
2 89815 1 11338
2 89816 1 11353
2 89817 1 11353
2 89818 1 11353
2 89819 1 11353
2 89820 1 11369
2 89821 1 11369
2 89822 1 11369
2 89823 1 11369
2 89824 1 11370
2 89825 1 11370
2 89826 1 11371
2 89827 1 11371
2 89828 1 11371
2 89829 1 11371
2 89830 1 11380
2 89831 1 11380
2 89832 1 11388
2 89833 1 11388
2 89834 1 11415
2 89835 1 11415
2 89836 1 11430
2 89837 1 11430
2 89838 1 11430
2 89839 1 11450
2 89840 1 11450
2 89841 1 11450
2 89842 1 11459
2 89843 1 11459
2 89844 1 11461
2 89845 1 11461
2 89846 1 11462
2 89847 1 11462
2 89848 1 11462
2 89849 1 11494
2 89850 1 11494
2 89851 1 11494
2 89852 1 11498
2 89853 1 11498
2 89854 1 11498
2 89855 1 11498
2 89856 1 11506
2 89857 1 11506
2 89858 1 11506
2 89859 1 11506
2 89860 1 11519
2 89861 1 11519
2 89862 1 11520
2 89863 1 11520
2 89864 1 11527
2 89865 1 11527
2 89866 1 11527
2 89867 1 11527
2 89868 1 11538
2 89869 1 11538
2 89870 1 11538
2 89871 1 11548
2 89872 1 11548
2 89873 1 11559
2 89874 1 11559
2 89875 1 11559
2 89876 1 11560
2 89877 1 11560
2 89878 1 11567
2 89879 1 11567
2 89880 1 11567
2 89881 1 11567
2 89882 1 11567
2 89883 1 11568
2 89884 1 11568
2 89885 1 11587
2 89886 1 11587
2 89887 1 11587
2 89888 1 11587
2 89889 1 11587
2 89890 1 11587
2 89891 1 11590
2 89892 1 11590
2 89893 1 11590
2 89894 1 11590
2 89895 1 11590
2 89896 1 11590
2 89897 1 11603
2 89898 1 11603
2 89899 1 11608
2 89900 1 11608
2 89901 1 11608
2 89902 1 11608
2 89903 1 11608
2 89904 1 11618
2 89905 1 11618
2 89906 1 11618
2 89907 1 11618
2 89908 1 11636
2 89909 1 11636
2 89910 1 11639
2 89911 1 11639
2 89912 1 11639
2 89913 1 11639
2 89914 1 11639
2 89915 1 11639
2 89916 1 11639
2 89917 1 11639
2 89918 1 11639
2 89919 1 11639
2 89920 1 11639
2 89921 1 11647
2 89922 1 11647
2 89923 1 11647
2 89924 1 11647
2 89925 1 11647
2 89926 1 11673
2 89927 1 11673
2 89928 1 11692
2 89929 1 11692
2 89930 1 11692
2 89931 1 11692
2 89932 1 11692
2 89933 1 11692
2 89934 1 11692
2 89935 1 11692
2 89936 1 11692
2 89937 1 11692
2 89938 1 11692
2 89939 1 11692
2 89940 1 11692
2 89941 1 11692
2 89942 1 11696
2 89943 1 11696
2 89944 1 11696
2 89945 1 11696
2 89946 1 11696
2 89947 1 11696
2 89948 1 11697
2 89949 1 11697
2 89950 1 11697
2 89951 1 11697
2 89952 1 11697
2 89953 1 11697
2 89954 1 11698
2 89955 1 11698
2 89956 1 11698
2 89957 1 11698
2 89958 1 11721
2 89959 1 11721
2 89960 1 11734
2 89961 1 11734
2 89962 1 11759
2 89963 1 11759
2 89964 1 11768
2 89965 1 11768
2 89966 1 11794
2 89967 1 11794
2 89968 1 11794
2 89969 1 11806
2 89970 1 11806
2 89971 1 11806
2 89972 1 11806
2 89973 1 11823
2 89974 1 11823
2 89975 1 11823
2 89976 1 11835
2 89977 1 11835
2 89978 1 11835
2 89979 1 11835
2 89980 1 11835
2 89981 1 11835
2 89982 1 11835
2 89983 1 11835
2 89984 1 11835
2 89985 1 11836
2 89986 1 11836
2 89987 1 11843
2 89988 1 11843
2 89989 1 11851
2 89990 1 11851
2 89991 1 11851
2 89992 1 11890
2 89993 1 11890
2 89994 1 11900
2 89995 1 11900
2 89996 1 11911
2 89997 1 11911
2 89998 1 11912
2 89999 1 11912
2 90000 1 11929
2 90001 1 11929
2 90002 1 11929
2 90003 1 11929
2 90004 1 11929
2 90005 1 11929
2 90006 1 11929
2 90007 1 11929
2 90008 1 11929
2 90009 1 11929
2 90010 1 11929
2 90011 1 11929
2 90012 1 11930
2 90013 1 11930
2 90014 1 11930
2 90015 1 11941
2 90016 1 11941
2 90017 1 11941
2 90018 1 11965
2 90019 1 11965
2 90020 1 11980
2 90021 1 11980
2 90022 1 11981
2 90023 1 11981
2 90024 1 11981
2 90025 1 11981
2 90026 1 11981
2 90027 1 11981
2 90028 1 11981
2 90029 1 11981
2 90030 1 11981
2 90031 1 11981
2 90032 1 11981
2 90033 1 11981
2 90034 1 11983
2 90035 1 11983
2 90036 1 11983
2 90037 1 11983
2 90038 1 11983
2 90039 1 11984
2 90040 1 11984
2 90041 1 11988
2 90042 1 11988
2 90043 1 11988
2 90044 1 11988
2 90045 1 11988
2 90046 1 11992
2 90047 1 11992
2 90048 1 11992
2 90049 1 12006
2 90050 1 12006
2 90051 1 12006
2 90052 1 12007
2 90053 1 12007
2 90054 1 12007
2 90055 1 12007
2 90056 1 12008
2 90057 1 12008
2 90058 1 12009
2 90059 1 12009
2 90060 1 12010
2 90061 1 12010
2 90062 1 12010
2 90063 1 12022
2 90064 1 12022
2 90065 1 12022
2 90066 1 12022
2 90067 1 12044
2 90068 1 12044
2 90069 1 12045
2 90070 1 12045
2 90071 1 12051
2 90072 1 12051
2 90073 1 12051
2 90074 1 12051
2 90075 1 12051
2 90076 1 12051
2 90077 1 12059
2 90078 1 12059
2 90079 1 12059
2 90080 1 12062
2 90081 1 12062
2 90082 1 12062
2 90083 1 12069
2 90084 1 12069
2 90085 1 12069
2 90086 1 12069
2 90087 1 12069
2 90088 1 12069
2 90089 1 12069
2 90090 1 12070
2 90091 1 12070
2 90092 1 12070
2 90093 1 12078
2 90094 1 12078
2 90095 1 12092
2 90096 1 12092
2 90097 1 12092
2 90098 1 12104
2 90099 1 12104
2 90100 1 12104
2 90101 1 12104
2 90102 1 12112
2 90103 1 12112
2 90104 1 12112
2 90105 1 12112
2 90106 1 12112
2 90107 1 12112
2 90108 1 12122
2 90109 1 12122
2 90110 1 12123
2 90111 1 12123
2 90112 1 12136
2 90113 1 12136
2 90114 1 12136
2 90115 1 12136
2 90116 1 12144
2 90117 1 12144
2 90118 1 12144
2 90119 1 12144
2 90120 1 12144
2 90121 1 12144
2 90122 1 12144
2 90123 1 12144
2 90124 1 12144
2 90125 1 12144
2 90126 1 12170
2 90127 1 12170
2 90128 1 12170
2 90129 1 12175
2 90130 1 12175
2 90131 1 12179
2 90132 1 12179
2 90133 1 12191
2 90134 1 12191
2 90135 1 12191
2 90136 1 12191
2 90137 1 12191
2 90138 1 12191
2 90139 1 12192
2 90140 1 12192
2 90141 1 12213
2 90142 1 12213
2 90143 1 12213
2 90144 1 12227
2 90145 1 12227
2 90146 1 12236
2 90147 1 12236
2 90148 1 12250
2 90149 1 12250
2 90150 1 12250
2 90151 1 12250
2 90152 1 12254
2 90153 1 12254
2 90154 1 12256
2 90155 1 12256
2 90156 1 12274
2 90157 1 12274
2 90158 1 12303
2 90159 1 12303
2 90160 1 12303
2 90161 1 12336
2 90162 1 12336
2 90163 1 12348
2 90164 1 12348
2 90165 1 12350
2 90166 1 12350
2 90167 1 12351
2 90168 1 12351
2 90169 1 12361
2 90170 1 12361
2 90171 1 12361
2 90172 1 12361
2 90173 1 12361
2 90174 1 12361
2 90175 1 12362
2 90176 1 12362
2 90177 1 12363
2 90178 1 12363
2 90179 1 12363
2 90180 1 12363
2 90181 1 12364
2 90182 1 12364
2 90183 1 12366
2 90184 1 12366
2 90185 1 12366
2 90186 1 12366
2 90187 1 12366
2 90188 1 12366
2 90189 1 12366
2 90190 1 12366
2 90191 1 12366
2 90192 1 12366
2 90193 1 12366
2 90194 1 12366
2 90195 1 12366
2 90196 1 12366
2 90197 1 12366
2 90198 1 12366
2 90199 1 12366
2 90200 1 12366
2 90201 1 12366
2 90202 1 12366
2 90203 1 12366
2 90204 1 12366
2 90205 1 12366
2 90206 1 12366
2 90207 1 12366
2 90208 1 12366
2 90209 1 12366
2 90210 1 12366
2 90211 1 12366
2 90212 1 12366
2 90213 1 12366
2 90214 1 12366
2 90215 1 12366
2 90216 1 12366
2 90217 1 12366
2 90218 1 12366
2 90219 1 12367
2 90220 1 12367
2 90221 1 12367
2 90222 1 12367
2 90223 1 12367
2 90224 1 12368
2 90225 1 12368
2 90226 1 12371
2 90227 1 12371
2 90228 1 12371
2 90229 1 12388
2 90230 1 12388
2 90231 1 12388
2 90232 1 12388
2 90233 1 12388
2 90234 1 12388
2 90235 1 12388
2 90236 1 12388
2 90237 1 12388
2 90238 1 12388
2 90239 1 12388
2 90240 1 12388
2 90241 1 12388
2 90242 1 12388
2 90243 1 12388
2 90244 1 12388
2 90245 1 12388
2 90246 1 12388
2 90247 1 12388
2 90248 1 12388
2 90249 1 12397
2 90250 1 12397
2 90251 1 12412
2 90252 1 12412
2 90253 1 12415
2 90254 1 12415
2 90255 1 12418
2 90256 1 12418
2 90257 1 12418
2 90258 1 12418
2 90259 1 12418
2 90260 1 12418
2 90261 1 12418
2 90262 1 12418
2 90263 1 12418
2 90264 1 12418
2 90265 1 12418
2 90266 1 12418
2 90267 1 12418
2 90268 1 12418
2 90269 1 12418
2 90270 1 12418
2 90271 1 12418
2 90272 1 12418
2 90273 1 12418
2 90274 1 12418
2 90275 1 12418
2 90276 1 12418
2 90277 1 12418
2 90278 1 12418
2 90279 1 12418
2 90280 1 12418
2 90281 1 12418
2 90282 1 12418
2 90283 1 12418
2 90284 1 12418
2 90285 1 12420
2 90286 1 12420
2 90287 1 12421
2 90288 1 12421
2 90289 1 12424
2 90290 1 12424
2 90291 1 12424
2 90292 1 12425
2 90293 1 12425
2 90294 1 12425
2 90295 1 12428
2 90296 1 12428
2 90297 1 12437
2 90298 1 12437
2 90299 1 12440
2 90300 1 12440
2 90301 1 12440
2 90302 1 12447
2 90303 1 12447
2 90304 1 12452
2 90305 1 12452
2 90306 1 12470
2 90307 1 12470
2 90308 1 12470
2 90309 1 12470
2 90310 1 12485
2 90311 1 12485
2 90312 1 12485
2 90313 1 12485
2 90314 1 12485
2 90315 1 12485
2 90316 1 12485
2 90317 1 12488
2 90318 1 12488
2 90319 1 12488
2 90320 1 12488
2 90321 1 12488
2 90322 1 12488
2 90323 1 12488
2 90324 1 12488
2 90325 1 12489
2 90326 1 12489
2 90327 1 12490
2 90328 1 12490
2 90329 1 12512
2 90330 1 12512
2 90331 1 12522
2 90332 1 12522
2 90333 1 12528
2 90334 1 12528
2 90335 1 12529
2 90336 1 12529
2 90337 1 12530
2 90338 1 12530
2 90339 1 12547
2 90340 1 12547
2 90341 1 12547
2 90342 1 12547
2 90343 1 12547
2 90344 1 12547
2 90345 1 12547
2 90346 1 12547
2 90347 1 12547
2 90348 1 12547
2 90349 1 12547
2 90350 1 12547
2 90351 1 12547
2 90352 1 12547
2 90353 1 12547
2 90354 1 12547
2 90355 1 12551
2 90356 1 12551
2 90357 1 12551
2 90358 1 12560
2 90359 1 12560
2 90360 1 12567
2 90361 1 12567
2 90362 1 12587
2 90363 1 12587
2 90364 1 12597
2 90365 1 12597
2 90366 1 12610
2 90367 1 12610
2 90368 1 12612
2 90369 1 12612
2 90370 1 12625
2 90371 1 12625
2 90372 1 12625
2 90373 1 12625
2 90374 1 12625
2 90375 1 12625
2 90376 1 12625
2 90377 1 12625
2 90378 1 12625
2 90379 1 12625
2 90380 1 12626
2 90381 1 12626
2 90382 1 12645
2 90383 1 12645
2 90384 1 12648
2 90385 1 12648
2 90386 1 12659
2 90387 1 12659
2 90388 1 12659
2 90389 1 12659
2 90390 1 12660
2 90391 1 12660
2 90392 1 12668
2 90393 1 12668
2 90394 1 12678
2 90395 1 12678
2 90396 1 12698
2 90397 1 12698
2 90398 1 12699
2 90399 1 12699
2 90400 1 12706
2 90401 1 12706
2 90402 1 12724
2 90403 1 12724
2 90404 1 12729
2 90405 1 12729
2 90406 1 12729
2 90407 1 12736
2 90408 1 12736
2 90409 1 12736
2 90410 1 12753
2 90411 1 12753
2 90412 1 12754
2 90413 1 12754
2 90414 1 12770
2 90415 1 12770
2 90416 1 12783
2 90417 1 12783
2 90418 1 12783
2 90419 1 12803
2 90420 1 12803
2 90421 1 12803
2 90422 1 12803
2 90423 1 12803
2 90424 1 12817
2 90425 1 12817
2 90426 1 12838
2 90427 1 12838
2 90428 1 12838
2 90429 1 12845
2 90430 1 12845
2 90431 1 12847
2 90432 1 12847
2 90433 1 12868
2 90434 1 12868
2 90435 1 12871
2 90436 1 12871
2 90437 1 12871
2 90438 1 12878
2 90439 1 12878
2 90440 1 12878
2 90441 1 12878
2 90442 1 12878
2 90443 1 12878
2 90444 1 12878
2 90445 1 12879
2 90446 1 12879
2 90447 1 12880
2 90448 1 12880
2 90449 1 12893
2 90450 1 12893
2 90451 1 12893
2 90452 1 12903
2 90453 1 12903
2 90454 1 12903
2 90455 1 12903
2 90456 1 12911
2 90457 1 12911
2 90458 1 12911
2 90459 1 12915
2 90460 1 12915
2 90461 1 12929
2 90462 1 12929
2 90463 1 12937
2 90464 1 12937
2 90465 1 12965
2 90466 1 12965
2 90467 1 12965
2 90468 1 12965
2 90469 1 12965
2 90470 1 12965
2 90471 1 12966
2 90472 1 12966
2 90473 1 12975
2 90474 1 12975
2 90475 1 12975
2 90476 1 12975
2 90477 1 12975
2 90478 1 12975
2 90479 1 12975
2 90480 1 12975
2 90481 1 12975
2 90482 1 12976
2 90483 1 12976
2 90484 1 12976
2 90485 1 12977
2 90486 1 12977
2 90487 1 12977
2 90488 1 12977
2 90489 1 12986
2 90490 1 12986
2 90491 1 12986
2 90492 1 12990
2 90493 1 12990
2 90494 1 12991
2 90495 1 12991
2 90496 1 12992
2 90497 1 12992
2 90498 1 13009
2 90499 1 13009
2 90500 1 13012
2 90501 1 13012
2 90502 1 13012
2 90503 1 13012
2 90504 1 13013
2 90505 1 13013
2 90506 1 13013
2 90507 1 13014
2 90508 1 13014
2 90509 1 13044
2 90510 1 13044
2 90511 1 13057
2 90512 1 13057
2 90513 1 13057
2 90514 1 13057
2 90515 1 13059
2 90516 1 13059
2 90517 1 13059
2 90518 1 13059
2 90519 1 13059
2 90520 1 13062
2 90521 1 13062
2 90522 1 13069
2 90523 1 13069
2 90524 1 13069
2 90525 1 13069
2 90526 1 13070
2 90527 1 13070
2 90528 1 13070
2 90529 1 13070
2 90530 1 13070
2 90531 1 13071
2 90532 1 13071
2 90533 1 13079
2 90534 1 13079
2 90535 1 13079
2 90536 1 13079
2 90537 1 13088
2 90538 1 13088
2 90539 1 13088
2 90540 1 13088
2 90541 1 13096
2 90542 1 13096
2 90543 1 13096
2 90544 1 13104
2 90545 1 13104
2 90546 1 13108
2 90547 1 13108
2 90548 1 13114
2 90549 1 13114
2 90550 1 13116
2 90551 1 13116
2 90552 1 13135
2 90553 1 13135
2 90554 1 13135
2 90555 1 13135
2 90556 1 13136
2 90557 1 13136
2 90558 1 13150
2 90559 1 13150
2 90560 1 13150
2 90561 1 13150
2 90562 1 13151
2 90563 1 13151
2 90564 1 13151
2 90565 1 13152
2 90566 1 13152
2 90567 1 13152
2 90568 1 13152
2 90569 1 13152
2 90570 1 13152
2 90571 1 13152
2 90572 1 13155
2 90573 1 13155
2 90574 1 13155
2 90575 1 13178
2 90576 1 13178
2 90577 1 13179
2 90578 1 13179
2 90579 1 13179
2 90580 1 13179
2 90581 1 13179
2 90582 1 13180
2 90583 1 13180
2 90584 1 13180
2 90585 1 13180
2 90586 1 13180
2 90587 1 13180
2 90588 1 13180
2 90589 1 13180
2 90590 1 13180
2 90591 1 13180
2 90592 1 13180
2 90593 1 13190
2 90594 1 13190
2 90595 1 13190
2 90596 1 13190
2 90597 1 13190
2 90598 1 13190
2 90599 1 13190
2 90600 1 13190
2 90601 1 13190
2 90602 1 13190
2 90603 1 13190
2 90604 1 13190
2 90605 1 13190
2 90606 1 13190
2 90607 1 13190
2 90608 1 13190
2 90609 1 13190
2 90610 1 13190
2 90611 1 13190
2 90612 1 13190
2 90613 1 13190
2 90614 1 13190
2 90615 1 13190
2 90616 1 13190
2 90617 1 13190
2 90618 1 13190
2 90619 1 13190
2 90620 1 13190
2 90621 1 13190
2 90622 1 13190
2 90623 1 13190
2 90624 1 13190
2 90625 1 13190
2 90626 1 13190
2 90627 1 13190
2 90628 1 13190
2 90629 1 13190
2 90630 1 13190
2 90631 1 13190
2 90632 1 13190
2 90633 1 13191
2 90634 1 13191
2 90635 1 13191
2 90636 1 13191
2 90637 1 13191
2 90638 1 13192
2 90639 1 13192
2 90640 1 13192
2 90641 1 13192
2 90642 1 13192
2 90643 1 13192
2 90644 1 13192
2 90645 1 13192
2 90646 1 13192
2 90647 1 13194
2 90648 1 13194
2 90649 1 13194
2 90650 1 13194
2 90651 1 13194
2 90652 1 13194
2 90653 1 13194
2 90654 1 13194
2 90655 1 13194
2 90656 1 13194
2 90657 1 13194
2 90658 1 13194
2 90659 1 13194
2 90660 1 13194
2 90661 1 13194
2 90662 1 13194
2 90663 1 13194
2 90664 1 13194
2 90665 1 13194
2 90666 1 13194
2 90667 1 13194
2 90668 1 13194
2 90669 1 13194
2 90670 1 13194
2 90671 1 13194
2 90672 1 13194
2 90673 1 13194
2 90674 1 13194
2 90675 1 13194
2 90676 1 13194
2 90677 1 13194
2 90678 1 13194
2 90679 1 13194
2 90680 1 13194
2 90681 1 13194
2 90682 1 13194
2 90683 1 13194
2 90684 1 13194
2 90685 1 13194
2 90686 1 13194
2 90687 1 13194
2 90688 1 13194
2 90689 1 13194
2 90690 1 13194
2 90691 1 13194
2 90692 1 13195
2 90693 1 13195
2 90694 1 13195
2 90695 1 13196
2 90696 1 13196
2 90697 1 13199
2 90698 1 13199
2 90699 1 13199
2 90700 1 13199
2 90701 1 13199
2 90702 1 13199
2 90703 1 13199
2 90704 1 13199
2 90705 1 13199
2 90706 1 13199
2 90707 1 13199
2 90708 1 13199
2 90709 1 13199
2 90710 1 13199
2 90711 1 13199
2 90712 1 13199
2 90713 1 13199
2 90714 1 13199
2 90715 1 13199
2 90716 1 13199
2 90717 1 13199
2 90718 1 13199
2 90719 1 13199
2 90720 1 13199
2 90721 1 13199
2 90722 1 13199
2 90723 1 13199
2 90724 1 13199
2 90725 1 13199
2 90726 1 13199
2 90727 1 13199
2 90728 1 13199
2 90729 1 13199
2 90730 1 13199
2 90731 1 13199
2 90732 1 13199
2 90733 1 13199
2 90734 1 13199
2 90735 1 13199
2 90736 1 13199
2 90737 1 13199
2 90738 1 13199
2 90739 1 13203
2 90740 1 13203
2 90741 1 13203
2 90742 1 13203
2 90743 1 13206
2 90744 1 13206
2 90745 1 13206
2 90746 1 13206
2 90747 1 13230
2 90748 1 13230
2 90749 1 13230
2 90750 1 13231
2 90751 1 13231
2 90752 1 13232
2 90753 1 13232
2 90754 1 13232
2 90755 1 13232
2 90756 1 13232
2 90757 1 13252
2 90758 1 13252
2 90759 1 13252
2 90760 1 13252
2 90761 1 13253
2 90762 1 13253
2 90763 1 13253
2 90764 1 13253
2 90765 1 13253
2 90766 1 13253
2 90767 1 13253
2 90768 1 13253
2 90769 1 13253
2 90770 1 13253
2 90771 1 13253
2 90772 1 13253
2 90773 1 13253
2 90774 1 13253
2 90775 1 13253
2 90776 1 13253
2 90777 1 13253
2 90778 1 13253
2 90779 1 13253
2 90780 1 13253
2 90781 1 13253
2 90782 1 13253
2 90783 1 13254
2 90784 1 13254
2 90785 1 13261
2 90786 1 13261
2 90787 1 13261
2 90788 1 13261
2 90789 1 13262
2 90790 1 13262
2 90791 1 13262
2 90792 1 13275
2 90793 1 13275
2 90794 1 13275
2 90795 1 13275
2 90796 1 13275
2 90797 1 13275
2 90798 1 13276
2 90799 1 13276
2 90800 1 13276
2 90801 1 13284
2 90802 1 13284
2 90803 1 13284
2 90804 1 13293
2 90805 1 13293
2 90806 1 13301
2 90807 1 13301
2 90808 1 13301
2 90809 1 13301
2 90810 1 13301
2 90811 1 13302
2 90812 1 13302
2 90813 1 13309
2 90814 1 13309
2 90815 1 13310
2 90816 1 13310
2 90817 1 13310
2 90818 1 13310
2 90819 1 13319
2 90820 1 13319
2 90821 1 13319
2 90822 1 13331
2 90823 1 13331
2 90824 1 13331
2 90825 1 13331
2 90826 1 13331
2 90827 1 13339
2 90828 1 13339
2 90829 1 13359
2 90830 1 13359
2 90831 1 13360
2 90832 1 13360
2 90833 1 13369
2 90834 1 13369
2 90835 1 13374
2 90836 1 13374
2 90837 1 13391
2 90838 1 13391
2 90839 1 13391
2 90840 1 13399
2 90841 1 13399
2 90842 1 13399
2 90843 1 13399
2 90844 1 13406
2 90845 1 13406
2 90846 1 13406
2 90847 1 13406
2 90848 1 13406
2 90849 1 13406
2 90850 1 13408
2 90851 1 13408
2 90852 1 13424
2 90853 1 13424
2 90854 1 13425
2 90855 1 13425
2 90856 1 13426
2 90857 1 13426
2 90858 1 13426
2 90859 1 13426
2 90860 1 13426
2 90861 1 13426
2 90862 1 13426
2 90863 1 13426
2 90864 1 13426
2 90865 1 13426
2 90866 1 13426
2 90867 1 13426
2 90868 1 13426
2 90869 1 13426
2 90870 1 13426
2 90871 1 13426
2 90872 1 13427
2 90873 1 13427
2 90874 1 13427
2 90875 1 13427
2 90876 1 13427
2 90877 1 13427
2 90878 1 13427
2 90879 1 13427
2 90880 1 13427
2 90881 1 13427
2 90882 1 13427
2 90883 1 13427
2 90884 1 13427
2 90885 1 13436
2 90886 1 13436
2 90887 1 13436
2 90888 1 13436
2 90889 1 13436
2 90890 1 13442
2 90891 1 13442
2 90892 1 13442
2 90893 1 13442
2 90894 1 13443
2 90895 1 13443
2 90896 1 13443
2 90897 1 13450
2 90898 1 13450
2 90899 1 13450
2 90900 1 13452
2 90901 1 13452
2 90902 1 13452
2 90903 1 13452
2 90904 1 13452
2 90905 1 13452
2 90906 1 13452
2 90907 1 13452
2 90908 1 13452
2 90909 1 13464
2 90910 1 13464
2 90911 1 13473
2 90912 1 13473
2 90913 1 13473
2 90914 1 13473
2 90915 1 13473
2 90916 1 13479
2 90917 1 13479
2 90918 1 13479
2 90919 1 13499
2 90920 1 13499
2 90921 1 13499
2 90922 1 13499
2 90923 1 13501
2 90924 1 13501
2 90925 1 13501
2 90926 1 13523
2 90927 1 13523
2 90928 1 13523
2 90929 1 13548
2 90930 1 13548
2 90931 1 13548
2 90932 1 13548
2 90933 1 13548
2 90934 1 13548
2 90935 1 13548
2 90936 1 13548
2 90937 1 13548
2 90938 1 13548
2 90939 1 13565
2 90940 1 13565
2 90941 1 13584
2 90942 1 13584
2 90943 1 13584
2 90944 1 13590
2 90945 1 13590
2 90946 1 13598
2 90947 1 13598
2 90948 1 13598
2 90949 1 13598
2 90950 1 13598
2 90951 1 13598
2 90952 1 13599
2 90953 1 13599
2 90954 1 13599
2 90955 1 13600
2 90956 1 13600
2 90957 1 13600
2 90958 1 13600
2 90959 1 13600
2 90960 1 13600
2 90961 1 13600
2 90962 1 13600
2 90963 1 13600
2 90964 1 13601
2 90965 1 13601
2 90966 1 13601
2 90967 1 13601
2 90968 1 13602
2 90969 1 13602
2 90970 1 13602
2 90971 1 13607
2 90972 1 13607
2 90973 1 13614
2 90974 1 13614
2 90975 1 13614
2 90976 1 13614
2 90977 1 13614
2 90978 1 13614
2 90979 1 13614
2 90980 1 13614
2 90981 1 13614
2 90982 1 13614
2 90983 1 13614
2 90984 1 13615
2 90985 1 13615
2 90986 1 13615
2 90987 1 13615
2 90988 1 13615
2 90989 1 13615
2 90990 1 13615
2 90991 1 13615
2 90992 1 13615
2 90993 1 13615
2 90994 1 13615
2 90995 1 13615
2 90996 1 13615
2 90997 1 13615
2 90998 1 13615
2 90999 1 13615
2 91000 1 13615
2 91001 1 13615
2 91002 1 13615
2 91003 1 13615
2 91004 1 13616
2 91005 1 13616
2 91006 1 13616
2 91007 1 13616
2 91008 1 13616
2 91009 1 13616
2 91010 1 13616
2 91011 1 13616
2 91012 1 13624
2 91013 1 13624
2 91014 1 13624
2 91015 1 13627
2 91016 1 13627
2 91017 1 13627
2 91018 1 13627
2 91019 1 13627
2 91020 1 13627
2 91021 1 13627
2 91022 1 13627
2 91023 1 13627
2 91024 1 13627
2 91025 1 13627
2 91026 1 13627
2 91027 1 13627
2 91028 1 13627
2 91029 1 13627
2 91030 1 13627
2 91031 1 13627
2 91032 1 13627
2 91033 1 13627
2 91034 1 13627
2 91035 1 13627
2 91036 1 13627
2 91037 1 13627
2 91038 1 13627
2 91039 1 13627
2 91040 1 13628
2 91041 1 13628
2 91042 1 13628
2 91043 1 13629
2 91044 1 13629
2 91045 1 13629
2 91046 1 13629
2 91047 1 13629
2 91048 1 13630
2 91049 1 13630
2 91050 1 13637
2 91051 1 13637
2 91052 1 13638
2 91053 1 13638
2 91054 1 13638
2 91055 1 13647
2 91056 1 13647
2 91057 1 13648
2 91058 1 13648
2 91059 1 13648
2 91060 1 13648
2 91061 1 13649
2 91062 1 13649
2 91063 1 13649
2 91064 1 13657
2 91065 1 13657
2 91066 1 13657
2 91067 1 13657
2 91068 1 13690
2 91069 1 13690
2 91070 1 13691
2 91071 1 13691
2 91072 1 13693
2 91073 1 13693
2 91074 1 13698
2 91075 1 13698
2 91076 1 13709
2 91077 1 13709
2 91078 1 13710
2 91079 1 13710
2 91080 1 13710
2 91081 1 13712
2 91082 1 13712
2 91083 1 13715
2 91084 1 13715
2 91085 1 13715
2 91086 1 13715
2 91087 1 13715
2 91088 1 13715
2 91089 1 13715
2 91090 1 13715
2 91091 1 13715
2 91092 1 13715
2 91093 1 13715
2 91094 1 13715
2 91095 1 13715
2 91096 1 13715
2 91097 1 13715
2 91098 1 13716
2 91099 1 13716
2 91100 1 13723
2 91101 1 13723
2 91102 1 13723
2 91103 1 13723
2 91104 1 13723
2 91105 1 13723
2 91106 1 13723
2 91107 1 13723
2 91108 1 13723
2 91109 1 13723
2 91110 1 13723
2 91111 1 13724
2 91112 1 13724
2 91113 1 13724
2 91114 1 13726
2 91115 1 13726
2 91116 1 13739
2 91117 1 13739
2 91118 1 13744
2 91119 1 13744
2 91120 1 13752
2 91121 1 13752
2 91122 1 13752
2 91123 1 13752
2 91124 1 13752
2 91125 1 13752
2 91126 1 13752
2 91127 1 13761
2 91128 1 13761
2 91129 1 13761
2 91130 1 13762
2 91131 1 13762
2 91132 1 13769
2 91133 1 13769
2 91134 1 13808
2 91135 1 13808
2 91136 1 13808
2 91137 1 13811
2 91138 1 13811
2 91139 1 13829
2 91140 1 13829
2 91141 1 13829
2 91142 1 13840
2 91143 1 13840
2 91144 1 13840
2 91145 1 13841
2 91146 1 13841
2 91147 1 13841
2 91148 1 13841
2 91149 1 13841
2 91150 1 13841
2 91151 1 13841
2 91152 1 13841
2 91153 1 13841
2 91154 1 13860
2 91155 1 13860
2 91156 1 13860
2 91157 1 13860
2 91158 1 13861
2 91159 1 13861
2 91160 1 13861
2 91161 1 13861
2 91162 1 13861
2 91163 1 13861
2 91164 1 13861
2 91165 1 13861
2 91166 1 13864
2 91167 1 13864
2 91168 1 13865
2 91169 1 13865
2 91170 1 13865
2 91171 1 13883
2 91172 1 13883
2 91173 1 13884
2 91174 1 13884
2 91175 1 13885
2 91176 1 13885
2 91177 1 13909
2 91178 1 13909
2 91179 1 13918
2 91180 1 13918
2 91181 1 13918
2 91182 1 13919
2 91183 1 13919
2 91184 1 13919
2 91185 1 13919
2 91186 1 13919
2 91187 1 13919
2 91188 1 13919
2 91189 1 13919
2 91190 1 13919
2 91191 1 13919
2 91192 1 13919
2 91193 1 13919
2 91194 1 13919
2 91195 1 13919
2 91196 1 13919
2 91197 1 13920
2 91198 1 13920
2 91199 1 13920
2 91200 1 13920
2 91201 1 13921
2 91202 1 13921
2 91203 1 13931
2 91204 1 13931
2 91205 1 13941
2 91206 1 13941
2 91207 1 13941
2 91208 1 13941
2 91209 1 13941
2 91210 1 13942
2 91211 1 13942
2 91212 1 13942
2 91213 1 13942
2 91214 1 13942
2 91215 1 13942
2 91216 1 13943
2 91217 1 13943
2 91218 1 13955
2 91219 1 13955
2 91220 1 13955
2 91221 1 13955
2 91222 1 13956
2 91223 1 13956
2 91224 1 13959
2 91225 1 13959
2 91226 1 13975
2 91227 1 13975
2 91228 1 13975
2 91229 1 13975
2 91230 1 13975
2 91231 1 13975
2 91232 1 13978
2 91233 1 13978
2 91234 1 13978
2 91235 1 13979
2 91236 1 13979
2 91237 1 13988
2 91238 1 13988
2 91239 1 14007
2 91240 1 14007
2 91241 1 14012
2 91242 1 14012
2 91243 1 14012
2 91244 1 14013
2 91245 1 14013
2 91246 1 14013
2 91247 1 14013
2 91248 1 14013
2 91249 1 14015
2 91250 1 14015
2 91251 1 14015
2 91252 1 14015
2 91253 1 14016
2 91254 1 14016
2 91255 1 14016
2 91256 1 14016
2 91257 1 14016
2 91258 1 14016
2 91259 1 14016
2 91260 1 14016
2 91261 1 14016
2 91262 1 14034
2 91263 1 14034
2 91264 1 14034
2 91265 1 14034
2 91266 1 14060
2 91267 1 14060
2 91268 1 14060
2 91269 1 14060
2 91270 1 14060
2 91271 1 14060
2 91272 1 14073
2 91273 1 14073
2 91274 1 14073
2 91275 1 14073
2 91276 1 14088
2 91277 1 14088
2 91278 1 14088
2 91279 1 14088
2 91280 1 14088
2 91281 1 14088
2 91282 1 14088
2 91283 1 14088
2 91284 1 14088
2 91285 1 14088
2 91286 1 14089
2 91287 1 14089
2 91288 1 14100
2 91289 1 14100
2 91290 1 14118
2 91291 1 14118
2 91292 1 14132
2 91293 1 14132
2 91294 1 14132
2 91295 1 14134
2 91296 1 14134
2 91297 1 14134
2 91298 1 14137
2 91299 1 14137
2 91300 1 14137
2 91301 1 14137
2 91302 1 14137
2 91303 1 14137
2 91304 1 14137
2 91305 1 14137
2 91306 1 14137
2 91307 1 14137
2 91308 1 14137
2 91309 1 14137
2 91310 1 14137
2 91311 1 14137
2 91312 1 14137
2 91313 1 14137
2 91314 1 14150
2 91315 1 14150
2 91316 1 14160
2 91317 1 14160
2 91318 1 14161
2 91319 1 14161
2 91320 1 14161
2 91321 1 14161
2 91322 1 14161
2 91323 1 14161
2 91324 1 14161
2 91325 1 14166
2 91326 1 14166
2 91327 1 14167
2 91328 1 14167
2 91329 1 14167
2 91330 1 14167
2 91331 1 14167
2 91332 1 14167
2 91333 1 14179
2 91334 1 14179
2 91335 1 14185
2 91336 1 14185
2 91337 1 14186
2 91338 1 14186
2 91339 1 14197
2 91340 1 14197
2 91341 1 14197
2 91342 1 14197
2 91343 1 14197
2 91344 1 14197
2 91345 1 14197
2 91346 1 14197
2 91347 1 14197
2 91348 1 14197
2 91349 1 14197
2 91350 1 14197
2 91351 1 14197
2 91352 1 14197
2 91353 1 14197
2 91354 1 14197
2 91355 1 14198
2 91356 1 14198
2 91357 1 14198
2 91358 1 14198
2 91359 1 14207
2 91360 1 14207
2 91361 1 14207
2 91362 1 14207
2 91363 1 14207
2 91364 1 14207
2 91365 1 14208
2 91366 1 14208
2 91367 1 14208
2 91368 1 14208
2 91369 1 14208
2 91370 1 14208
2 91371 1 14208
2 91372 1 14208
2 91373 1 14208
2 91374 1 14208
2 91375 1 14208
2 91376 1 14208
2 91377 1 14208
2 91378 1 14210
2 91379 1 14210
2 91380 1 14210
2 91381 1 14210
2 91382 1 14210
2 91383 1 14210
2 91384 1 14210
2 91385 1 14210
2 91386 1 14212
2 91387 1 14212
2 91388 1 14212
2 91389 1 14212
2 91390 1 14212
2 91391 1 14212
2 91392 1 14212
2 91393 1 14212
2 91394 1 14212
2 91395 1 14229
2 91396 1 14229
2 91397 1 14237
2 91398 1 14237
2 91399 1 14238
2 91400 1 14238
2 91401 1 14257
2 91402 1 14257
2 91403 1 14260
2 91404 1 14260
2 91405 1 14262
2 91406 1 14262
2 91407 1 14263
2 91408 1 14263
2 91409 1 14273
2 91410 1 14273
2 91411 1 14273
2 91412 1 14276
2 91413 1 14276
2 91414 1 14277
2 91415 1 14277
2 91416 1 14277
2 91417 1 14277
2 91418 1 14290
2 91419 1 14290
2 91420 1 14291
2 91421 1 14291
2 91422 1 14291
2 91423 1 14291
2 91424 1 14291
2 91425 1 14291
2 91426 1 14291
2 91427 1 14291
2 91428 1 14291
2 91429 1 14291
2 91430 1 14291
2 91431 1 14291
2 91432 1 14291
2 91433 1 14291
2 91434 1 14291
2 91435 1 14291
2 91436 1 14291
2 91437 1 14291
2 91438 1 14291
2 91439 1 14291
2 91440 1 14291
2 91441 1 14292
2 91442 1 14292
2 91443 1 14292
2 91444 1 14314
2 91445 1 14314
2 91446 1 14314
2 91447 1 14314
2 91448 1 14314
2 91449 1 14316
2 91450 1 14316
2 91451 1 14316
2 91452 1 14316
2 91453 1 14316
2 91454 1 14316
2 91455 1 14331
2 91456 1 14331
2 91457 1 14331
2 91458 1 14342
2 91459 1 14342
2 91460 1 14342
2 91461 1 14342
2 91462 1 14343
2 91463 1 14343
2 91464 1 14351
2 91465 1 14351
2 91466 1 14351
2 91467 1 14353
2 91468 1 14353
2 91469 1 14358
2 91470 1 14358
2 91471 1 14359
2 91472 1 14359
2 91473 1 14365
2 91474 1 14365
2 91475 1 14365
2 91476 1 14365
2 91477 1 14366
2 91478 1 14366
2 91479 1 14369
2 91480 1 14369
2 91481 1 14371
2 91482 1 14371
2 91483 1 14371
2 91484 1 14371
2 91485 1 14371
2 91486 1 14379
2 91487 1 14379
2 91488 1 14379
2 91489 1 14379
2 91490 1 14391
2 91491 1 14391
2 91492 1 14406
2 91493 1 14406
2 91494 1 14407
2 91495 1 14407
2 91496 1 14416
2 91497 1 14416
2 91498 1 14416
2 91499 1 14417
2 91500 1 14417
2 91501 1 14422
2 91502 1 14422
2 91503 1 14428
2 91504 1 14428
2 91505 1 14440
2 91506 1 14440
2 91507 1 14440
2 91508 1 14440
2 91509 1 14440
2 91510 1 14448
2 91511 1 14448
2 91512 1 14448
2 91513 1 14448
2 91514 1 14448
2 91515 1 14448
2 91516 1 14448
2 91517 1 14448
2 91518 1 14448
2 91519 1 14448
2 91520 1 14448
2 91521 1 14448
2 91522 1 14457
2 91523 1 14457
2 91524 1 14458
2 91525 1 14458
2 91526 1 14458
2 91527 1 14458
2 91528 1 14470
2 91529 1 14470
2 91530 1 14470
2 91531 1 14473
2 91532 1 14473
2 91533 1 14474
2 91534 1 14474
2 91535 1 14474
2 91536 1 14474
2 91537 1 14474
2 91538 1 14483
2 91539 1 14483
2 91540 1 14483
2 91541 1 14483
2 91542 1 14483
2 91543 1 14484
2 91544 1 14484
2 91545 1 14484
2 91546 1 14491
2 91547 1 14491
2 91548 1 14491
2 91549 1 14494
2 91550 1 14494
2 91551 1 14508
2 91552 1 14508
2 91553 1 14508
2 91554 1 14508
2 91555 1 14517
2 91556 1 14517
2 91557 1 14517
2 91558 1 14519
2 91559 1 14519
2 91560 1 14519
2 91561 1 14520
2 91562 1 14520
2 91563 1 14520
2 91564 1 14521
2 91565 1 14521
2 91566 1 14521
2 91567 1 14529
2 91568 1 14529
2 91569 1 14554
2 91570 1 14554
2 91571 1 14554
2 91572 1 14557
2 91573 1 14557
2 91574 1 14561
2 91575 1 14561
2 91576 1 14570
2 91577 1 14570
2 91578 1 14570
2 91579 1 14570
2 91580 1 14570
2 91581 1 14570
2 91582 1 14570
2 91583 1 14571
2 91584 1 14571
2 91585 1 14571
2 91586 1 14571
2 91587 1 14571
2 91588 1 14571
2 91589 1 14571
2 91590 1 14580
2 91591 1 14580
2 91592 1 14581
2 91593 1 14581
2 91594 1 14584
2 91595 1 14584
2 91596 1 14593
2 91597 1 14593
2 91598 1 14593
2 91599 1 14609
2 91600 1 14609
2 91601 1 14609
2 91602 1 14609
2 91603 1 14609
2 91604 1 14609
2 91605 1 14609
2 91606 1 14609
2 91607 1 14619
2 91608 1 14619
2 91609 1 14634
2 91610 1 14634
2 91611 1 14634
2 91612 1 14635
2 91613 1 14635
2 91614 1 14635
2 91615 1 14635
2 91616 1 14635
2 91617 1 14637
2 91618 1 14637
2 91619 1 14639
2 91620 1 14639
2 91621 1 14639
2 91622 1 14640
2 91623 1 14640
2 91624 1 14640
2 91625 1 14647
2 91626 1 14647
2 91627 1 14647
2 91628 1 14648
2 91629 1 14648
2 91630 1 14648
2 91631 1 14648
2 91632 1 14649
2 91633 1 14649
2 91634 1 14649
2 91635 1 14649
2 91636 1 14649
2 91637 1 14649
2 91638 1 14658
2 91639 1 14658
2 91640 1 14659
2 91641 1 14659
2 91642 1 14680
2 91643 1 14680
2 91644 1 14683
2 91645 1 14683
2 91646 1 14683
2 91647 1 14683
2 91648 1 14683
2 91649 1 14683
2 91650 1 14683
2 91651 1 14696
2 91652 1 14696
2 91653 1 14710
2 91654 1 14710
2 91655 1 14722
2 91656 1 14722
2 91657 1 14722
2 91658 1 14722
2 91659 1 14730
2 91660 1 14730
2 91661 1 14730
2 91662 1 14730
2 91663 1 14730
2 91664 1 14731
2 91665 1 14731
2 91666 1 14731
2 91667 1 14732
2 91668 1 14732
2 91669 1 14732
2 91670 1 14732
2 91671 1 14737
2 91672 1 14737
2 91673 1 14737
2 91674 1 14737
2 91675 1 14737
2 91676 1 14757
2 91677 1 14757
2 91678 1 14757
2 91679 1 14757
2 91680 1 14785
2 91681 1 14785
2 91682 1 14785
2 91683 1 14785
2 91684 1 14785
2 91685 1 14787
2 91686 1 14787
2 91687 1 14787
2 91688 1 14787
2 91689 1 14787
2 91690 1 14787
2 91691 1 14787
2 91692 1 14787
2 91693 1 14787
2 91694 1 14787
2 91695 1 14787
2 91696 1 14787
2 91697 1 14787
2 91698 1 14787
2 91699 1 14787
2 91700 1 14787
2 91701 1 14787
2 91702 1 14787
2 91703 1 14787
2 91704 1 14788
2 91705 1 14788
2 91706 1 14789
2 91707 1 14789
2 91708 1 14792
2 91709 1 14792
2 91710 1 14793
2 91711 1 14793
2 91712 1 14793
2 91713 1 14796
2 91714 1 14796
2 91715 1 14804
2 91716 1 14804
2 91717 1 14805
2 91718 1 14805
2 91719 1 14805
2 91720 1 14805
2 91721 1 14814
2 91722 1 14814
2 91723 1 14814
2 91724 1 14814
2 91725 1 14814
2 91726 1 14824
2 91727 1 14824
2 91728 1 14824
2 91729 1 14825
2 91730 1 14825
2 91731 1 14827
2 91732 1 14827
2 91733 1 14827
2 91734 1 14827
2 91735 1 14830
2 91736 1 14830
2 91737 1 14837
2 91738 1 14837
2 91739 1 14837
2 91740 1 14838
2 91741 1 14838
2 91742 1 14855
2 91743 1 14855
2 91744 1 14855
2 91745 1 14858
2 91746 1 14858
2 91747 1 14858
2 91748 1 14858
2 91749 1 14858
2 91750 1 14866
2 91751 1 14866
2 91752 1 14866
2 91753 1 14869
2 91754 1 14869
2 91755 1 14869
2 91756 1 14870
2 91757 1 14870
2 91758 1 14876
2 91759 1 14876
2 91760 1 14884
2 91761 1 14884
2 91762 1 14884
2 91763 1 14884
2 91764 1 14884
2 91765 1 14892
2 91766 1 14892
2 91767 1 14892
2 91768 1 14892
2 91769 1 14901
2 91770 1 14901
2 91771 1 14901
2 91772 1 14901
2 91773 1 14901
2 91774 1 14903
2 91775 1 14903
2 91776 1 14913
2 91777 1 14913
2 91778 1 14913
2 91779 1 14913
2 91780 1 14913
2 91781 1 14918
2 91782 1 14918
2 91783 1 14919
2 91784 1 14919
2 91785 1 14919
2 91786 1 14919
2 91787 1 14930
2 91788 1 14930
2 91789 1 14930
2 91790 1 14936
2 91791 1 14936
2 91792 1 14936
2 91793 1 14936
2 91794 1 14945
2 91795 1 14945
2 91796 1 14946
2 91797 1 14946
2 91798 1 14946
2 91799 1 14946
2 91800 1 14946
2 91801 1 14947
2 91802 1 14947
2 91803 1 14956
2 91804 1 14956
2 91805 1 14956
2 91806 1 14956
2 91807 1 14959
2 91808 1 14959
2 91809 1 14959
2 91810 1 14959
2 91811 1 14959
2 91812 1 14959
2 91813 1 14959
2 91814 1 14959
2 91815 1 14959
2 91816 1 14959
2 91817 1 14961
2 91818 1 14961
2 91819 1 14962
2 91820 1 14962
2 91821 1 14962
2 91822 1 14972
2 91823 1 14972
2 91824 1 14972
2 91825 1 14972
2 91826 1 14972
2 91827 1 14972
2 91828 1 14972
2 91829 1 14972
2 91830 1 14972
2 91831 1 14972
2 91832 1 14972
2 91833 1 14972
2 91834 1 14973
2 91835 1 14973
2 91836 1 14973
2 91837 1 14973
2 91838 1 14983
2 91839 1 14983
2 91840 1 14984
2 91841 1 14984
2 91842 1 14984
2 91843 1 14984
2 91844 1 14984
2 91845 1 14984
2 91846 1 14984
2 91847 1 14984
2 91848 1 14984
2 91849 1 14984
2 91850 1 14984
2 91851 1 14984
2 91852 1 14984
2 91853 1 14985
2 91854 1 14985
2 91855 1 14987
2 91856 1 14987
2 91857 1 14987
2 91858 1 14987
2 91859 1 14987
2 91860 1 14987
2 91861 1 14987
2 91862 1 14987
2 91863 1 14987
2 91864 1 14987
2 91865 1 14987
2 91866 1 14987
2 91867 1 14987
2 91868 1 14987
2 91869 1 14987
2 91870 1 14987
2 91871 1 14987
2 91872 1 14987
2 91873 1 14987
2 91874 1 14987
2 91875 1 14988
2 91876 1 14988
2 91877 1 14988
2 91878 1 14988
2 91879 1 14988
2 91880 1 14988
2 91881 1 14988
2 91882 1 14988
2 91883 1 14988
2 91884 1 14988
2 91885 1 14989
2 91886 1 14989
2 91887 1 14989
2 91888 1 14989
2 91889 1 14990
2 91890 1 14990
2 91891 1 14990
2 91892 1 14990
2 91893 1 14990
2 91894 1 14998
2 91895 1 14998
2 91896 1 14999
2 91897 1 14999
2 91898 1 15001
2 91899 1 15001
2 91900 1 15001
2 91901 1 15001
2 91902 1 15008
2 91903 1 15008
2 91904 1 15009
2 91905 1 15009
2 91906 1 15013
2 91907 1 15013
2 91908 1 15013
2 91909 1 15021
2 91910 1 15021
2 91911 1 15031
2 91912 1 15031
2 91913 1 15043
2 91914 1 15043
2 91915 1 15057
2 91916 1 15057
2 91917 1 15058
2 91918 1 15058
2 91919 1 15058
2 91920 1 15058
2 91921 1 15059
2 91922 1 15059
2 91923 1 15068
2 91924 1 15068
2 91925 1 15083
2 91926 1 15083
2 91927 1 15098
2 91928 1 15098
2 91929 1 15098
2 91930 1 15099
2 91931 1 15099
2 91932 1 15100
2 91933 1 15100
2 91934 1 15110
2 91935 1 15110
2 91936 1 15114
2 91937 1 15114
2 91938 1 15128
2 91939 1 15128
2 91940 1 15128
2 91941 1 15128
2 91942 1 15128
2 91943 1 15128
2 91944 1 15128
2 91945 1 15128
2 91946 1 15128
2 91947 1 15128
2 91948 1 15128
2 91949 1 15129
2 91950 1 15129
2 91951 1 15129
2 91952 1 15129
2 91953 1 15129
2 91954 1 15129
2 91955 1 15129
2 91956 1 15131
2 91957 1 15131
2 91958 1 15131
2 91959 1 15131
2 91960 1 15134
2 91961 1 15134
2 91962 1 15134
2 91963 1 15134
2 91964 1 15134
2 91965 1 15134
2 91966 1 15138
2 91967 1 15138
2 91968 1 15138
2 91969 1 15150
2 91970 1 15150
2 91971 1 15150
2 91972 1 15153
2 91973 1 15153
2 91974 1 15153
2 91975 1 15153
2 91976 1 15153
2 91977 1 15153
2 91978 1 15153
2 91979 1 15153
2 91980 1 15153
2 91981 1 15154
2 91982 1 15154
2 91983 1 15154
2 91984 1 15154
2 91985 1 15154
2 91986 1 15155
2 91987 1 15155
2 91988 1 15155
2 91989 1 15155
2 91990 1 15165
2 91991 1 15165
2 91992 1 15173
2 91993 1 15173
2 91994 1 15173
2 91995 1 15173
2 91996 1 15173
2 91997 1 15190
2 91998 1 15190
2 91999 1 15190
2 92000 1 15191
2 92001 1 15191
2 92002 1 15192
2 92003 1 15192
2 92004 1 15209
2 92005 1 15209
2 92006 1 15213
2 92007 1 15213
2 92008 1 15213
2 92009 1 15213
2 92010 1 15214
2 92011 1 15214
2 92012 1 15214
2 92013 1 15214
2 92014 1 15214
2 92015 1 15214
2 92016 1 15214
2 92017 1 15214
2 92018 1 15234
2 92019 1 15234
2 92020 1 15234
2 92021 1 15234
2 92022 1 15234
2 92023 1 15234
2 92024 1 15234
2 92025 1 15234
2 92026 1 15238
2 92027 1 15238
2 92028 1 15238
2 92029 1 15238
2 92030 1 15247
2 92031 1 15247
2 92032 1 15248
2 92033 1 15248
2 92034 1 15248
2 92035 1 15248
2 92036 1 15258
2 92037 1 15258
2 92038 1 15258
2 92039 1 15259
2 92040 1 15259
2 92041 1 15259
2 92042 1 15259
2 92043 1 15260
2 92044 1 15260
2 92045 1 15260
2 92046 1 15260
2 92047 1 15264
2 92048 1 15264
2 92049 1 15264
2 92050 1 15264
2 92051 1 15264
2 92052 1 15264
2 92053 1 15264
2 92054 1 15265
2 92055 1 15265
2 92056 1 15266
2 92057 1 15266
2 92058 1 15270
2 92059 1 15270
2 92060 1 15273
2 92061 1 15273
2 92062 1 15291
2 92063 1 15291
2 92064 1 15291
2 92065 1 15291
2 92066 1 15291
2 92067 1 15291
2 92068 1 15291
2 92069 1 15291
2 92070 1 15334
2 92071 1 15334
2 92072 1 15334
2 92073 1 15343
2 92074 1 15343
2 92075 1 15343
2 92076 1 15352
2 92077 1 15352
2 92078 1 15364
2 92079 1 15364
2 92080 1 15364
2 92081 1 15367
2 92082 1 15367
2 92083 1 15368
2 92084 1 15368
2 92085 1 15401
2 92086 1 15401
2 92087 1 15401
2 92088 1 15444
2 92089 1 15444
2 92090 1 15444
2 92091 1 15444
2 92092 1 15445
2 92093 1 15445
2 92094 1 15452
2 92095 1 15452
2 92096 1 15452
2 92097 1 15452
2 92098 1 15452
2 92099 1 15452
2 92100 1 15452
2 92101 1 15452
2 92102 1 15452
2 92103 1 15452
2 92104 1 15453
2 92105 1 15453
2 92106 1 15466
2 92107 1 15466
2 92108 1 15467
2 92109 1 15467
2 92110 1 15489
2 92111 1 15489
2 92112 1 15489
2 92113 1 15489
2 92114 1 15489
2 92115 1 15489
2 92116 1 15489
2 92117 1 15489
2 92118 1 15489
2 92119 1 15489
2 92120 1 15489
2 92121 1 15489
2 92122 1 15490
2 92123 1 15490
2 92124 1 15490
2 92125 1 15490
2 92126 1 15498
2 92127 1 15498
2 92128 1 15502
2 92129 1 15502
2 92130 1 15502
2 92131 1 15503
2 92132 1 15503
2 92133 1 15511
2 92134 1 15511
2 92135 1 15511
2 92136 1 15511
2 92137 1 15513
2 92138 1 15513
2 92139 1 15527
2 92140 1 15527
2 92141 1 15528
2 92142 1 15528
2 92143 1 15531
2 92144 1 15531
2 92145 1 15531
2 92146 1 15545
2 92147 1 15545
2 92148 1 15545
2 92149 1 15554
2 92150 1 15554
2 92151 1 15554
2 92152 1 15554
2 92153 1 15555
2 92154 1 15555
2 92155 1 15563
2 92156 1 15563
2 92157 1 15563
2 92158 1 15583
2 92159 1 15583
2 92160 1 15583
2 92161 1 15583
2 92162 1 15584
2 92163 1 15584
2 92164 1 15598
2 92165 1 15598
2 92166 1 15598
2 92167 1 15598
2 92168 1 15598
2 92169 1 15598
2 92170 1 15598
2 92171 1 15598
2 92172 1 15598
2 92173 1 15598
2 92174 1 15598
2 92175 1 15598
2 92176 1 15598
2 92177 1 15598
2 92178 1 15598
2 92179 1 15598
2 92180 1 15598
2 92181 1 15598
2 92182 1 15598
2 92183 1 15598
2 92184 1 15598
2 92185 1 15598
2 92186 1 15598
2 92187 1 15604
2 92188 1 15604
2 92189 1 15604
2 92190 1 15604
2 92191 1 15604
2 92192 1 15604
2 92193 1 15604
2 92194 1 15604
2 92195 1 15604
2 92196 1 15604
2 92197 1 15604
2 92198 1 15604
2 92199 1 15604
2 92200 1 15604
2 92201 1 15604
2 92202 1 15604
2 92203 1 15604
2 92204 1 15606
2 92205 1 15606
2 92206 1 15606
2 92207 1 15606
2 92208 1 15607
2 92209 1 15607
2 92210 1 15607
2 92211 1 15607
2 92212 1 15607
2 92213 1 15607
2 92214 1 15607
2 92215 1 15607
2 92216 1 15607
2 92217 1 15607
2 92218 1 15607
2 92219 1 15607
2 92220 1 15607
2 92221 1 15607
2 92222 1 15608
2 92223 1 15608
2 92224 1 15608
2 92225 1 15620
2 92226 1 15620
2 92227 1 15624
2 92228 1 15624
2 92229 1 15624
2 92230 1 15624
2 92231 1 15624
2 92232 1 15631
2 92233 1 15631
2 92234 1 15631
2 92235 1 15646
2 92236 1 15646
2 92237 1 15646
2 92238 1 15646
2 92239 1 15646
2 92240 1 15648
2 92241 1 15648
2 92242 1 15650
2 92243 1 15650
2 92244 1 15677
2 92245 1 15677
2 92246 1 15677
2 92247 1 15677
2 92248 1 15677
2 92249 1 15684
2 92250 1 15684
2 92251 1 15692
2 92252 1 15692
2 92253 1 15710
2 92254 1 15710
2 92255 1 15717
2 92256 1 15717
2 92257 1 15717
2 92258 1 15725
2 92259 1 15725
2 92260 1 15733
2 92261 1 15733
2 92262 1 15733
2 92263 1 15733
2 92264 1 15733
2 92265 1 15733
2 92266 1 15735
2 92267 1 15735
2 92268 1 15736
2 92269 1 15736
2 92270 1 15747
2 92271 1 15747
2 92272 1 15747
2 92273 1 15760
2 92274 1 15760
2 92275 1 15760
2 92276 1 15769
2 92277 1 15769
2 92278 1 15771
2 92279 1 15771
2 92280 1 15771
2 92281 1 15771
2 92282 1 15771
2 92283 1 15798
2 92284 1 15798
2 92285 1 15798
2 92286 1 15798
2 92287 1 15799
2 92288 1 15799
2 92289 1 15799
2 92290 1 15799
2 92291 1 15799
2 92292 1 15809
2 92293 1 15809
2 92294 1 15809
2 92295 1 15810
2 92296 1 15810
2 92297 1 15811
2 92298 1 15811
2 92299 1 15812
2 92300 1 15812
2 92301 1 15826
2 92302 1 15826
2 92303 1 15837
2 92304 1 15837
2 92305 1 15837
2 92306 1 15838
2 92307 1 15838
2 92308 1 15841
2 92309 1 15841
2 92310 1 15841
2 92311 1 15849
2 92312 1 15849
2 92313 1 15869
2 92314 1 15869
2 92315 1 15894
2 92316 1 15894
2 92317 1 15901
2 92318 1 15901
2 92319 1 15909
2 92320 1 15909
2 92321 1 15909
2 92322 1 15909
2 92323 1 15909
2 92324 1 15911
2 92325 1 15911
2 92326 1 15911
2 92327 1 15912
2 92328 1 15912
2 92329 1 15912
2 92330 1 15912
2 92331 1 15912
2 92332 1 15914
2 92333 1 15914
2 92334 1 15925
2 92335 1 15925
2 92336 1 15928
2 92337 1 15928
2 92338 1 15934
2 92339 1 15934
2 92340 1 15934
2 92341 1 15934
2 92342 1 15934
2 92343 1 15948
2 92344 1 15948
2 92345 1 15948
2 92346 1 15948
2 92347 1 15948
2 92348 1 15948
2 92349 1 15948
2 92350 1 15948
2 92351 1 15950
2 92352 1 15950
2 92353 1 15958
2 92354 1 15958
2 92355 1 15965
2 92356 1 15965
2 92357 1 15965
2 92358 1 15965
2 92359 1 15965
2 92360 1 15965
2 92361 1 15965
2 92362 1 15965
2 92363 1 15982
2 92364 1 15982
2 92365 1 15999
2 92366 1 15999
2 92367 1 16012
2 92368 1 16012
2 92369 1 16027
2 92370 1 16027
2 92371 1 16027
2 92372 1 16027
2 92373 1 16028
2 92374 1 16028
2 92375 1 16028
2 92376 1 16028
2 92377 1 16029
2 92378 1 16029
2 92379 1 16031
2 92380 1 16031
2 92381 1 16040
2 92382 1 16040
2 92383 1 16040
2 92384 1 16048
2 92385 1 16048
2 92386 1 16080
2 92387 1 16080
2 92388 1 16080
2 92389 1 16087
2 92390 1 16087
2 92391 1 16088
2 92392 1 16088
2 92393 1 16095
2 92394 1 16095
2 92395 1 16103
2 92396 1 16103
2 92397 1 16103
2 92398 1 16103
2 92399 1 16103
2 92400 1 16103
2 92401 1 16103
2 92402 1 16103
2 92403 1 16103
2 92404 1 16104
2 92405 1 16104
2 92406 1 16105
2 92407 1 16105
2 92408 1 16106
2 92409 1 16106
2 92410 1 16106
2 92411 1 16107
2 92412 1 16107
2 92413 1 16114
2 92414 1 16114
2 92415 1 16140
2 92416 1 16140
2 92417 1 16140
2 92418 1 16140
2 92419 1 16140
2 92420 1 16140
2 92421 1 16146
2 92422 1 16146
2 92423 1 16156
2 92424 1 16156
2 92425 1 16157
2 92426 1 16157
2 92427 1 16157
2 92428 1 16162
2 92429 1 16162
2 92430 1 16190
2 92431 1 16190
2 92432 1 16190
2 92433 1 16190
2 92434 1 16191
2 92435 1 16191
2 92436 1 16191
2 92437 1 16191
2 92438 1 16191
2 92439 1 16192
2 92440 1 16192
2 92441 1 16193
2 92442 1 16193
2 92443 1 16193
2 92444 1 16196
2 92445 1 16196
2 92446 1 16196
2 92447 1 16196
2 92448 1 16204
2 92449 1 16204
2 92450 1 16225
2 92451 1 16225
2 92452 1 16225
2 92453 1 16227
2 92454 1 16227
2 92455 1 16227
2 92456 1 16227
2 92457 1 16227
2 92458 1 16227
2 92459 1 16227
2 92460 1 16227
2 92461 1 16227
2 92462 1 16230
2 92463 1 16230
2 92464 1 16230
2 92465 1 16230
2 92466 1 16230
2 92467 1 16230
2 92468 1 16230
2 92469 1 16230
2 92470 1 16230
2 92471 1 16230
2 92472 1 16230
2 92473 1 16230
2 92474 1 16230
2 92475 1 16230
2 92476 1 16230
2 92477 1 16230
2 92478 1 16230
2 92479 1 16230
2 92480 1 16230
2 92481 1 16230
2 92482 1 16230
2 92483 1 16230
2 92484 1 16230
2 92485 1 16230
2 92486 1 16230
2 92487 1 16230
2 92488 1 16230
2 92489 1 16230
2 92490 1 16230
2 92491 1 16230
2 92492 1 16230
2 92493 1 16230
2 92494 1 16230
2 92495 1 16230
2 92496 1 16230
2 92497 1 16243
2 92498 1 16243
2 92499 1 16243
2 92500 1 16264
2 92501 1 16264
2 92502 1 16264
2 92503 1 16264
2 92504 1 16272
2 92505 1 16272
2 92506 1 16283
2 92507 1 16283
2 92508 1 16312
2 92509 1 16312
2 92510 1 16313
2 92511 1 16313
2 92512 1 16331
2 92513 1 16331
2 92514 1 16331
2 92515 1 16331
2 92516 1 16331
2 92517 1 16332
2 92518 1 16332
2 92519 1 16343
2 92520 1 16343
2 92521 1 16343
2 92522 1 16345
2 92523 1 16345
2 92524 1 16345
2 92525 1 16363
2 92526 1 16363
2 92527 1 16372
2 92528 1 16372
2 92529 1 16397
2 92530 1 16397
2 92531 1 16397
2 92532 1 16397
2 92533 1 16400
2 92534 1 16400
2 92535 1 16400
2 92536 1 16400
2 92537 1 16408
2 92538 1 16408
2 92539 1 16408
2 92540 1 16408
2 92541 1 16408
2 92542 1 16408
2 92543 1 16424
2 92544 1 16424
2 92545 1 16424
2 92546 1 16424
2 92547 1 16424
2 92548 1 16424
2 92549 1 16424
2 92550 1 16424
2 92551 1 16424
2 92552 1 16424
2 92553 1 16424
2 92554 1 16424
2 92555 1 16424
2 92556 1 16424
2 92557 1 16424
2 92558 1 16424
2 92559 1 16424
2 92560 1 16424
2 92561 1 16424
2 92562 1 16424
2 92563 1 16426
2 92564 1 16426
2 92565 1 16429
2 92566 1 16429
2 92567 1 16433
2 92568 1 16433
2 92569 1 16444
2 92570 1 16444
2 92571 1 16444
2 92572 1 16444
2 92573 1 16444
2 92574 1 16444
2 92575 1 16455
2 92576 1 16455
2 92577 1 16459
2 92578 1 16459
2 92579 1 16459
2 92580 1 16469
2 92581 1 16469
2 92582 1 16469
2 92583 1 16469
2 92584 1 16500
2 92585 1 16500
2 92586 1 16504
2 92587 1 16504
2 92588 1 16504
2 92589 1 16506
2 92590 1 16506
2 92591 1 16506
2 92592 1 16507
2 92593 1 16507
2 92594 1 16520
2 92595 1 16520
2 92596 1 16521
2 92597 1 16521
2 92598 1 16528
2 92599 1 16528
2 92600 1 16528
2 92601 1 16528
2 92602 1 16528
2 92603 1 16535
2 92604 1 16535
2 92605 1 16537
2 92606 1 16537
2 92607 1 16542
2 92608 1 16542
2 92609 1 16556
2 92610 1 16556
2 92611 1 16558
2 92612 1 16558
2 92613 1 16564
2 92614 1 16564
2 92615 1 16564
2 92616 1 16564
2 92617 1 16564
2 92618 1 16572
2 92619 1 16572
2 92620 1 16572
2 92621 1 16600
2 92622 1 16600
2 92623 1 16603
2 92624 1 16603
2 92625 1 16605
2 92626 1 16605
2 92627 1 16620
2 92628 1 16620
2 92629 1 16620
2 92630 1 16629
2 92631 1 16629
2 92632 1 16629
2 92633 1 16629
2 92634 1 16629
2 92635 1 16629
2 92636 1 16629
2 92637 1 16630
2 92638 1 16630
2 92639 1 16630
2 92640 1 16630
2 92641 1 16630
2 92642 1 16630
2 92643 1 16630
2 92644 1 16630
2 92645 1 16630
2 92646 1 16630
2 92647 1 16630
2 92648 1 16630
2 92649 1 16630
2 92650 1 16630
2 92651 1 16630
2 92652 1 16630
2 92653 1 16630
2 92654 1 16630
2 92655 1 16630
2 92656 1 16630
2 92657 1 16630
2 92658 1 16630
2 92659 1 16631
2 92660 1 16631
2 92661 1 16631
2 92662 1 16632
2 92663 1 16632
2 92664 1 16632
2 92665 1 16641
2 92666 1 16641
2 92667 1 16641
2 92668 1 16641
2 92669 1 16641
2 92670 1 16641
2 92671 1 16641
2 92672 1 16641
2 92673 1 16641
2 92674 1 16641
2 92675 1 16641
2 92676 1 16641
2 92677 1 16641
2 92678 1 16641
2 92679 1 16642
2 92680 1 16642
2 92681 1 16643
2 92682 1 16643
2 92683 1 16646
2 92684 1 16646
2 92685 1 16646
2 92686 1 16646
2 92687 1 16653
2 92688 1 16653
2 92689 1 16653
2 92690 1 16662
2 92691 1 16662
2 92692 1 16670
2 92693 1 16670
2 92694 1 16670
2 92695 1 16673
2 92696 1 16673
2 92697 1 16673
2 92698 1 16673
2 92699 1 16673
2 92700 1 16673
2 92701 1 16673
2 92702 1 16673
2 92703 1 16673
2 92704 1 16673
2 92705 1 16673
2 92706 1 16673
2 92707 1 16673
2 92708 1 16673
2 92709 1 16673
2 92710 1 16673
2 92711 1 16673
2 92712 1 16673
2 92713 1 16673
2 92714 1 16673
2 92715 1 16673
2 92716 1 16673
2 92717 1 16673
2 92718 1 16674
2 92719 1 16674
2 92720 1 16683
2 92721 1 16683
2 92722 1 16684
2 92723 1 16684
2 92724 1 16693
2 92725 1 16693
2 92726 1 16693
2 92727 1 16693
2 92728 1 16693
2 92729 1 16698
2 92730 1 16698
2 92731 1 16698
2 92732 1 16698
2 92733 1 16698
2 92734 1 16723
2 92735 1 16723
2 92736 1 16723
2 92737 1 16723
2 92738 1 16726
2 92739 1 16726
2 92740 1 16726
2 92741 1 16726
2 92742 1 16726
2 92743 1 16726
2 92744 1 16726
2 92745 1 16731
2 92746 1 16731
2 92747 1 16740
2 92748 1 16740
2 92749 1 16741
2 92750 1 16741
2 92751 1 16759
2 92752 1 16759
2 92753 1 16760
2 92754 1 16760
2 92755 1 16771
2 92756 1 16771
2 92757 1 16771
2 92758 1 16773
2 92759 1 16773
2 92760 1 16785
2 92761 1 16785
2 92762 1 16785
2 92763 1 16792
2 92764 1 16792
2 92765 1 16792
2 92766 1 16792
2 92767 1 16792
2 92768 1 16792
2 92769 1 16792
2 92770 1 16792
2 92771 1 16792
2 92772 1 16792
2 92773 1 16792
2 92774 1 16792
2 92775 1 16792
2 92776 1 16792
2 92777 1 16792
2 92778 1 16792
2 92779 1 16792
2 92780 1 16792
2 92781 1 16792
2 92782 1 16792
2 92783 1 16792
2 92784 1 16792
2 92785 1 16792
2 92786 1 16792
2 92787 1 16792
2 92788 1 16792
2 92789 1 16792
2 92790 1 16792
2 92791 1 16792
2 92792 1 16792
2 92793 1 16792
2 92794 1 16792
2 92795 1 16792
2 92796 1 16792
2 92797 1 16792
2 92798 1 16792
2 92799 1 16792
2 92800 1 16792
2 92801 1 16792
2 92802 1 16792
2 92803 1 16792
2 92804 1 16792
2 92805 1 16792
2 92806 1 16792
2 92807 1 16792
2 92808 1 16792
2 92809 1 16792
2 92810 1 16792
2 92811 1 16792
2 92812 1 16792
2 92813 1 16792
2 92814 1 16792
2 92815 1 16792
2 92816 1 16792
2 92817 1 16792
2 92818 1 16792
2 92819 1 16792
2 92820 1 16792
2 92821 1 16792
2 92822 1 16792
2 92823 1 16792
2 92824 1 16793
2 92825 1 16793
2 92826 1 16793
2 92827 1 16793
2 92828 1 16793
2 92829 1 16794
2 92830 1 16794
2 92831 1 16795
2 92832 1 16795
2 92833 1 16795
2 92834 1 16795
2 92835 1 16795
2 92836 1 16795
2 92837 1 16795
2 92838 1 16795
2 92839 1 16795
2 92840 1 16795
2 92841 1 16795
2 92842 1 16795
2 92843 1 16795
2 92844 1 16795
2 92845 1 16795
2 92846 1 16796
2 92847 1 16796
2 92848 1 16796
2 92849 1 16796
2 92850 1 16796
2 92851 1 16796
2 92852 1 16796
2 92853 1 16796
2 92854 1 16796
2 92855 1 16796
2 92856 1 16796
2 92857 1 16796
2 92858 1 16796
2 92859 1 16796
2 92860 1 16796
2 92861 1 16796
2 92862 1 16808
2 92863 1 16808
2 92864 1 16808
2 92865 1 16808
2 92866 1 16808
2 92867 1 16809
2 92868 1 16809
2 92869 1 16810
2 92870 1 16810
2 92871 1 16810
2 92872 1 16811
2 92873 1 16811
2 92874 1 16811
2 92875 1 16811
2 92876 1 16819
2 92877 1 16819
2 92878 1 16827
2 92879 1 16827
2 92880 1 16830
2 92881 1 16830
2 92882 1 16830
2 92883 1 16842
2 92884 1 16842
2 92885 1 16842
2 92886 1 16842
2 92887 1 16843
2 92888 1 16843
2 92889 1 16846
2 92890 1 16846
2 92891 1 16850
2 92892 1 16850
2 92893 1 16850
2 92894 1 16850
2 92895 1 16858
2 92896 1 16858
2 92897 1 16858
2 92898 1 16864
2 92899 1 16864
2 92900 1 16881
2 92901 1 16881
2 92902 1 16881
2 92903 1 16881
2 92904 1 16884
2 92905 1 16884
2 92906 1 16884
2 92907 1 16884
2 92908 1 16884
2 92909 1 16884
2 92910 1 16884
2 92911 1 16884
2 92912 1 16884
2 92913 1 16884
2 92914 1 16894
2 92915 1 16894
2 92916 1 16900
2 92917 1 16900
2 92918 1 16909
2 92919 1 16909
2 92920 1 16909
2 92921 1 16909
2 92922 1 16909
2 92923 1 16909
2 92924 1 16918
2 92925 1 16918
2 92926 1 16918
2 92927 1 16924
2 92928 1 16924
2 92929 1 16927
2 92930 1 16927
2 92931 1 16930
2 92932 1 16930
2 92933 1 16937
2 92934 1 16937
2 92935 1 16937
2 92936 1 16937
2 92937 1 16937
2 92938 1 16937
2 92939 1 16938
2 92940 1 16938
2 92941 1 16939
2 92942 1 16939
2 92943 1 16939
2 92944 1 16939
2 92945 1 16939
2 92946 1 16939
2 92947 1 16939
2 92948 1 16939
2 92949 1 16942
2 92950 1 16942
2 92951 1 16947
2 92952 1 16947
2 92953 1 16947
2 92954 1 16965
2 92955 1 16965
2 92956 1 16965
2 92957 1 16965
2 92958 1 16965
2 92959 1 16965
2 92960 1 16965
2 92961 1 16965
2 92962 1 16965
2 92963 1 16965
2 92964 1 16965
2 92965 1 16965
2 92966 1 16965
2 92967 1 16967
2 92968 1 16967
2 92969 1 16967
2 92970 1 16967
2 92971 1 16968
2 92972 1 16968
2 92973 1 16968
2 92974 1 16968
2 92975 1 16968
2 92976 1 16968
2 92977 1 16968
2 92978 1 16976
2 92979 1 16976
2 92980 1 16976
2 92981 1 16976
2 92982 1 16976
2 92983 1 16978
2 92984 1 16978
2 92985 1 16990
2 92986 1 16990
2 92987 1 16990
2 92988 1 16990
2 92989 1 16992
2 92990 1 16992
2 92991 1 16995
2 92992 1 16995
2 92993 1 16995
2 92994 1 16995
2 92995 1 17004
2 92996 1 17004
2 92997 1 17004
2 92998 1 17004
2 92999 1 17005
2 93000 1 17005
2 93001 1 17005
2 93002 1 17005
2 93003 1 17005
2 93004 1 17005
2 93005 1 17005
2 93006 1 17005
2 93007 1 17005
2 93008 1 17006
2 93009 1 17006
2 93010 1 17006
2 93011 1 17006
2 93012 1 17007
2 93013 1 17007
2 93014 1 17008
2 93015 1 17008
2 93016 1 17008
2 93017 1 17008
2 93018 1 17008
2 93019 1 17008
2 93020 1 17008
2 93021 1 17008
2 93022 1 17008
2 93023 1 17008
2 93024 1 17009
2 93025 1 17009
2 93026 1 17009
2 93027 1 17009
2 93028 1 17010
2 93029 1 17010
2 93030 1 17010
2 93031 1 17010
2 93032 1 17019
2 93033 1 17019
2 93034 1 17019
2 93035 1 17019
2 93036 1 17019
2 93037 1 17019
2 93038 1 17019
2 93039 1 17019
2 93040 1 17019
2 93041 1 17019
2 93042 1 17019
2 93043 1 17019
2 93044 1 17019
2 93045 1 17019
2 93046 1 17019
2 93047 1 17019
2 93048 1 17019
2 93049 1 17020
2 93050 1 17020
2 93051 1 17027
2 93052 1 17027
2 93053 1 17028
2 93054 1 17028
2 93055 1 17028
2 93056 1 17028
2 93057 1 17028
2 93058 1 17028
2 93059 1 17028
2 93060 1 17028
2 93061 1 17029
2 93062 1 17029
2 93063 1 17029
2 93064 1 17029
2 93065 1 17029
2 93066 1 17033
2 93067 1 17033
2 93068 1 17033
2 93069 1 17034
2 93070 1 17034
2 93071 1 17034
2 93072 1 17044
2 93073 1 17044
2 93074 1 17046
2 93075 1 17046
2 93076 1 17046
2 93077 1 17047
2 93078 1 17047
2 93079 1 17047
2 93080 1 17047
2 93081 1 17047
2 93082 1 17047
2 93083 1 17047
2 93084 1 17051
2 93085 1 17051
2 93086 1 17051
2 93087 1 17051
2 93088 1 17053
2 93089 1 17053
2 93090 1 17053
2 93091 1 17053
2 93092 1 17053
2 93093 1 17053
2 93094 1 17053
2 93095 1 17053
2 93096 1 17053
2 93097 1 17053
2 93098 1 17053
2 93099 1 17053
2 93100 1 17053
2 93101 1 17053
2 93102 1 17053
2 93103 1 17053
2 93104 1 17053
2 93105 1 17053
2 93106 1 17053
2 93107 1 17053
2 93108 1 17053
2 93109 1 17053
2 93110 1 17053
2 93111 1 17053
2 93112 1 17053
2 93113 1 17053
2 93114 1 17053
2 93115 1 17053
2 93116 1 17053
2 93117 1 17053
2 93118 1 17053
2 93119 1 17053
2 93120 1 17053
2 93121 1 17053
2 93122 1 17053
2 93123 1 17053
2 93124 1 17053
2 93125 1 17053
2 93126 1 17053
2 93127 1 17053
2 93128 1 17053
2 93129 1 17053
2 93130 1 17053
2 93131 1 17053
2 93132 1 17053
2 93133 1 17053
2 93134 1 17053
2 93135 1 17053
2 93136 1 17053
2 93137 1 17053
2 93138 1 17053
2 93139 1 17053
2 93140 1 17053
2 93141 1 17053
2 93142 1 17053
2 93143 1 17053
2 93144 1 17053
2 93145 1 17054
2 93146 1 17054
2 93147 1 17054
2 93148 1 17054
2 93149 1 17054
2 93150 1 17054
2 93151 1 17062
2 93152 1 17062
2 93153 1 17062
2 93154 1 17062
2 93155 1 17062
2 93156 1 17062
2 93157 1 17062
2 93158 1 17073
2 93159 1 17073
2 93160 1 17073
2 93161 1 17074
2 93162 1 17074
2 93163 1 17074
2 93164 1 17074
2 93165 1 17074
2 93166 1 17074
2 93167 1 17074
2 93168 1 17074
2 93169 1 17075
2 93170 1 17075
2 93171 1 17075
2 93172 1 17075
2 93173 1 17075
2 93174 1 17075
2 93175 1 17075
2 93176 1 17076
2 93177 1 17076
2 93178 1 17085
2 93179 1 17085
2 93180 1 17085
2 93181 1 17085
2 93182 1 17085
2 93183 1 17086
2 93184 1 17086
2 93185 1 17086
2 93186 1 17101
2 93187 1 17101
2 93188 1 17102
2 93189 1 17102
2 93190 1 17112
2 93191 1 17112
2 93192 1 17112
2 93193 1 17112
2 93194 1 17112
2 93195 1 17112
2 93196 1 17112
2 93197 1 17112
2 93198 1 17120
2 93199 1 17120
2 93200 1 17123
2 93201 1 17123
2 93202 1 17129
2 93203 1 17129
2 93204 1 17129
2 93205 1 17129
2 93206 1 17138
2 93207 1 17138
2 93208 1 17155
2 93209 1 17155
2 93210 1 17159
2 93211 1 17159
2 93212 1 17199
2 93213 1 17199
2 93214 1 17199
2 93215 1 17199
2 93216 1 17209
2 93217 1 17209
2 93218 1 17209
2 93219 1 17209
2 93220 1 17209
2 93221 1 17211
2 93222 1 17211
2 93223 1 17211
2 93224 1 17219
2 93225 1 17219
2 93226 1 17224
2 93227 1 17224
2 93228 1 17228
2 93229 1 17228
2 93230 1 17228
2 93231 1 17231
2 93232 1 17231
2 93233 1 17251
2 93234 1 17251
2 93235 1 17251
2 93236 1 17251
2 93237 1 17258
2 93238 1 17258
2 93239 1 17258
2 93240 1 17270
2 93241 1 17270
2 93242 1 17271
2 93243 1 17271
2 93244 1 17271
2 93245 1 17283
2 93246 1 17283
2 93247 1 17283
2 93248 1 17283
2 93249 1 17284
2 93250 1 17284
2 93251 1 17285
2 93252 1 17285
2 93253 1 17285
2 93254 1 17286
2 93255 1 17286
2 93256 1 17286
2 93257 1 17286
2 93258 1 17301
2 93259 1 17301
2 93260 1 17358
2 93261 1 17358
2 93262 1 17358
2 93263 1 17359
2 93264 1 17359
2 93265 1 17378
2 93266 1 17378
2 93267 1 17379
2 93268 1 17379
2 93269 1 17382
2 93270 1 17382
2 93271 1 17391
2 93272 1 17391
2 93273 1 17399
2 93274 1 17399
2 93275 1 17399
2 93276 1 17403
2 93277 1 17403
2 93278 1 17403
2 93279 1 17403
2 93280 1 17403
2 93281 1 17403
2 93282 1 17403
2 93283 1 17405
2 93284 1 17405
2 93285 1 17417
2 93286 1 17417
2 93287 1 17417
2 93288 1 17417
2 93289 1 17417
2 93290 1 17417
2 93291 1 17417
2 93292 1 17417
2 93293 1 17417
2 93294 1 17417
2 93295 1 17417
2 93296 1 17417
2 93297 1 17417
2 93298 1 17418
2 93299 1 17418
2 93300 1 17436
2 93301 1 17436
2 93302 1 17436
2 93303 1 17436
2 93304 1 17437
2 93305 1 17437
2 93306 1 17444
2 93307 1 17444
2 93308 1 17444
2 93309 1 17444
2 93310 1 17444
2 93311 1 17468
2 93312 1 17468
2 93313 1 17476
2 93314 1 17476
2 93315 1 17477
2 93316 1 17477
2 93317 1 17486
2 93318 1 17486
2 93319 1 17486
2 93320 1 17512
2 93321 1 17512
2 93322 1 17513
2 93323 1 17513
2 93324 1 17524
2 93325 1 17524
2 93326 1 17532
2 93327 1 17532
2 93328 1 17548
2 93329 1 17548
2 93330 1 17548
2 93331 1 17548
2 93332 1 17548
2 93333 1 17548
2 93334 1 17548
2 93335 1 17548
2 93336 1 17550
2 93337 1 17550
2 93338 1 17559
2 93339 1 17559
2 93340 1 17562
2 93341 1 17562
2 93342 1 17562
2 93343 1 17579
2 93344 1 17579
2 93345 1 17582
2 93346 1 17582
2 93347 1 17594
2 93348 1 17594
2 93349 1 17632
2 93350 1 17632
2 93351 1 17640
2 93352 1 17640
2 93353 1 17663
2 93354 1 17663
2 93355 1 17665
2 93356 1 17665
2 93357 1 17665
2 93358 1 17665
2 93359 1 17666
2 93360 1 17666
2 93361 1 17667
2 93362 1 17667
2 93363 1 17682
2 93364 1 17682
2 93365 1 17682
2 93366 1 17682
2 93367 1 17704
2 93368 1 17704
2 93369 1 17743
2 93370 1 17743
2 93371 1 17743
2 93372 1 17743
2 93373 1 17743
2 93374 1 17765
2 93375 1 17765
2 93376 1 17765
2 93377 1 17765
2 93378 1 17765
2 93379 1 17777
2 93380 1 17777
2 93381 1 17777
2 93382 1 17780
2 93383 1 17780
2 93384 1 17780
2 93385 1 17780
2 93386 1 17780
2 93387 1 17781
2 93388 1 17781
2 93389 1 17794
2 93390 1 17794
2 93391 1 17800
2 93392 1 17800
2 93393 1 17801
2 93394 1 17801
2 93395 1 17801
2 93396 1 17815
2 93397 1 17815
2 93398 1 17815
2 93399 1 17815
2 93400 1 17824
2 93401 1 17824
2 93402 1 17824
2 93403 1 17827
2 93404 1 17827
2 93405 1 17836
2 93406 1 17836
2 93407 1 17836
2 93408 1 17836
2 93409 1 17838
2 93410 1 17838
2 93411 1 17838
2 93412 1 17838
2 93413 1 17845
2 93414 1 17845
2 93415 1 17846
2 93416 1 17846
2 93417 1 17851
2 93418 1 17851
2 93419 1 17860
2 93420 1 17860
2 93421 1 17860
2 93422 1 17860
2 93423 1 17861
2 93424 1 17861
2 93425 1 17861
2 93426 1 17861
2 93427 1 17861
2 93428 1 17869
2 93429 1 17869
2 93430 1 17870
2 93431 1 17870
2 93432 1 17870
2 93433 1 17879
2 93434 1 17879
2 93435 1 17883
2 93436 1 17883
2 93437 1 17883
2 93438 1 17909
2 93439 1 17909
2 93440 1 17909
2 93441 1 17911
2 93442 1 17911
2 93443 1 17911
2 93444 1 17913
2 93445 1 17913
2 93446 1 17930
2 93447 1 17930
2 93448 1 17933
2 93449 1 17933
2 93450 1 17949
2 93451 1 17949
2 93452 1 17949
2 93453 1 17960
2 93454 1 17960
2 93455 1 17960
2 93456 1 17960
2 93457 1 17965
2 93458 1 17965
2 93459 1 17966
2 93460 1 17966
2 93461 1 18000
2 93462 1 18000
2 93463 1 18000
2 93464 1 18001
2 93465 1 18001
2 93466 1 18001
2 93467 1 18026
2 93468 1 18026
2 93469 1 18028
2 93470 1 18028
2 93471 1 18035
2 93472 1 18035
2 93473 1 18035
2 93474 1 18035
2 93475 1 18048
2 93476 1 18048
2 93477 1 18057
2 93478 1 18057
2 93479 1 18057
2 93480 1 18057
2 93481 1 18064
2 93482 1 18064
2 93483 1 18064
2 93484 1 18064
2 93485 1 18065
2 93486 1 18065
2 93487 1 18065
2 93488 1 18065
2 93489 1 18065
2 93490 1 18066
2 93491 1 18066
2 93492 1 18068
2 93493 1 18068
2 93494 1 18068
2 93495 1 18068
2 93496 1 18068
2 93497 1 18068
2 93498 1 18069
2 93499 1 18069
2 93500 1 18093
2 93501 1 18093
2 93502 1 18093
2 93503 1 18094
2 93504 1 18094
2 93505 1 18116
2 93506 1 18116
2 93507 1 18121
2 93508 1 18121
2 93509 1 18121
2 93510 1 18121
2 93511 1 18123
2 93512 1 18123
2 93513 1 18123
2 93514 1 18123
2 93515 1 18123
2 93516 1 18124
2 93517 1 18124
2 93518 1 18124
2 93519 1 18132
2 93520 1 18132
2 93521 1 18132
2 93522 1 18132
2 93523 1 18133
2 93524 1 18133
2 93525 1 18141
2 93526 1 18141
2 93527 1 18141
2 93528 1 18141
2 93529 1 18141
2 93530 1 18142
2 93531 1 18142
2 93532 1 18144
2 93533 1 18144
2 93534 1 18152
2 93535 1 18152
2 93536 1 18153
2 93537 1 18153
2 93538 1 18155
2 93539 1 18155
2 93540 1 18159
2 93541 1 18159
2 93542 1 18159
2 93543 1 18159
2 93544 1 18159
2 93545 1 18161
2 93546 1 18161
2 93547 1 18161
2 93548 1 18161
2 93549 1 18163
2 93550 1 18163
2 93551 1 18163
2 93552 1 18163
2 93553 1 18163
2 93554 1 18163
2 93555 1 18163
2 93556 1 18163
2 93557 1 18164
2 93558 1 18164
2 93559 1 18167
2 93560 1 18167
2 93561 1 18167
2 93562 1 18168
2 93563 1 18168
2 93564 1 18168
2 93565 1 18168
2 93566 1 18168
2 93567 1 18168
2 93568 1 18168
2 93569 1 18168
2 93570 1 18168
2 93571 1 18168
2 93572 1 18168
2 93573 1 18169
2 93574 1 18169
2 93575 1 18169
2 93576 1 18169
2 93577 1 18169
2 93578 1 18170
2 93579 1 18170
2 93580 1 18171
2 93581 1 18171
2 93582 1 18171
2 93583 1 18171
2 93584 1 18171
2 93585 1 18171
2 93586 1 18185
2 93587 1 18185
2 93588 1 18185
2 93589 1 18185
2 93590 1 18185
2 93591 1 18185
2 93592 1 18185
2 93593 1 18185
2 93594 1 18185
2 93595 1 18185
2 93596 1 18185
2 93597 1 18185
2 93598 1 18185
2 93599 1 18185
2 93600 1 18185
2 93601 1 18185
2 93602 1 18185
2 93603 1 18185
2 93604 1 18185
2 93605 1 18185
2 93606 1 18185
2 93607 1 18185
2 93608 1 18185
2 93609 1 18185
2 93610 1 18185
2 93611 1 18185
2 93612 1 18185
2 93613 1 18186
2 93614 1 18186
2 93615 1 18186
2 93616 1 18186
2 93617 1 18186
2 93618 1 18186
2 93619 1 18186
2 93620 1 18186
2 93621 1 18188
2 93622 1 18188
2 93623 1 18195
2 93624 1 18195
2 93625 1 18195
2 93626 1 18195
2 93627 1 18195
2 93628 1 18195
2 93629 1 18195
2 93630 1 18195
2 93631 1 18195
2 93632 1 18195
2 93633 1 18195
2 93634 1 18196
2 93635 1 18196
2 93636 1 18196
2 93637 1 18197
2 93638 1 18197
2 93639 1 18197
2 93640 1 18198
2 93641 1 18198
2 93642 1 18198
2 93643 1 18198
2 93644 1 18198
2 93645 1 18198
2 93646 1 18211
2 93647 1 18211
2 93648 1 18211
2 93649 1 18217
2 93650 1 18217
2 93651 1 18230
2 93652 1 18230
2 93653 1 18230
2 93654 1 18231
2 93655 1 18231
2 93656 1 18231
2 93657 1 18239
2 93658 1 18239
2 93659 1 18239
2 93660 1 18239
2 93661 1 18239
2 93662 1 18282
2 93663 1 18282
2 93664 1 18282
2 93665 1 18296
2 93666 1 18296
2 93667 1 18296
2 93668 1 18305
2 93669 1 18305
2 93670 1 18305
2 93671 1 18306
2 93672 1 18306
2 93673 1 18313
2 93674 1 18313
2 93675 1 18313
2 93676 1 18313
2 93677 1 18314
2 93678 1 18314
2 93679 1 18314
2 93680 1 18329
2 93681 1 18329
2 93682 1 18330
2 93683 1 18330
2 93684 1 18330
2 93685 1 18330
2 93686 1 18330
2 93687 1 18331
2 93688 1 18331
2 93689 1 18331
2 93690 1 18332
2 93691 1 18332
2 93692 1 18332
2 93693 1 18333
2 93694 1 18333
2 93695 1 18333
2 93696 1 18333
2 93697 1 18333
2 93698 1 18333
2 93699 1 18333
2 93700 1 18333
2 93701 1 18333
2 93702 1 18334
2 93703 1 18334
2 93704 1 18347
2 93705 1 18347
2 93706 1 18348
2 93707 1 18348
2 93708 1 18348
2 93709 1 18351
2 93710 1 18351
2 93711 1 18351
2 93712 1 18351
2 93713 1 18351
2 93714 1 18351
2 93715 1 18351
2 93716 1 18352
2 93717 1 18352
2 93718 1 18368
2 93719 1 18368
2 93720 1 18369
2 93721 1 18369
2 93722 1 18369
2 93723 1 18370
2 93724 1 18370
2 93725 1 18370
2 93726 1 18370
2 93727 1 18401
2 93728 1 18401
2 93729 1 18401
2 93730 1 18401
2 93731 1 18405
2 93732 1 18405
2 93733 1 18405
2 93734 1 18405
2 93735 1 18405
2 93736 1 18405
2 93737 1 18405
2 93738 1 18405
2 93739 1 18405
2 93740 1 18405
2 93741 1 18405
2 93742 1 18418
2 93743 1 18418
2 93744 1 18440
2 93745 1 18440
2 93746 1 18440
2 93747 1 18440
2 93748 1 18440
2 93749 1 18440
2 93750 1 18440
2 93751 1 18440
2 93752 1 18440
2 93753 1 18440
2 93754 1 18440
2 93755 1 18440
2 93756 1 18440
2 93757 1 18442
2 93758 1 18442
2 93759 1 18442
2 93760 1 18442
2 93761 1 18442
2 93762 1 18442
2 93763 1 18442
2 93764 1 18442
2 93765 1 18444
2 93766 1 18444
2 93767 1 18444
2 93768 1 18444
2 93769 1 18444
2 93770 1 18445
2 93771 1 18445
2 93772 1 18445
2 93773 1 18445
2 93774 1 18445
2 93775 1 18445
2 93776 1 18445
2 93777 1 18445
2 93778 1 18445
2 93779 1 18445
2 93780 1 18445
2 93781 1 18445
2 93782 1 18445
2 93783 1 18445
2 93784 1 18445
2 93785 1 18445
2 93786 1 18445
2 93787 1 18445
2 93788 1 18445
2 93789 1 18445
2 93790 1 18445
2 93791 1 18445
2 93792 1 18445
2 93793 1 18445
2 93794 1 18445
2 93795 1 18445
2 93796 1 18445
2 93797 1 18445
2 93798 1 18445
2 93799 1 18445
2 93800 1 18445
2 93801 1 18445
2 93802 1 18445
2 93803 1 18445
2 93804 1 18445
2 93805 1 18445
2 93806 1 18445
2 93807 1 18445
2 93808 1 18445
2 93809 1 18445
2 93810 1 18445
2 93811 1 18445
2 93812 1 18445
2 93813 1 18445
2 93814 1 18445
2 93815 1 18445
2 93816 1 18445
2 93817 1 18445
2 93818 1 18445
2 93819 1 18445
2 93820 1 18445
2 93821 1 18445
2 93822 1 18445
2 93823 1 18445
2 93824 1 18445
2 93825 1 18445
2 93826 1 18445
2 93827 1 18445
2 93828 1 18445
2 93829 1 18445
2 93830 1 18445
2 93831 1 18445
2 93832 1 18445
2 93833 1 18445
2 93834 1 18445
2 93835 1 18445
2 93836 1 18445
2 93837 1 18445
2 93838 1 18445
2 93839 1 18445
2 93840 1 18445
2 93841 1 18445
2 93842 1 18445
2 93843 1 18445
2 93844 1 18446
2 93845 1 18446
2 93846 1 18446
2 93847 1 18446
2 93848 1 18449
2 93849 1 18449
2 93850 1 18449
2 93851 1 18449
2 93852 1 18449
2 93853 1 18449
2 93854 1 18449
2 93855 1 18449
2 93856 1 18449
2 93857 1 18449
2 93858 1 18449
2 93859 1 18449
2 93860 1 18449
2 93861 1 18449
2 93862 1 18449
2 93863 1 18449
2 93864 1 18449
2 93865 1 18449
2 93866 1 18449
2 93867 1 18449
2 93868 1 18449
2 93869 1 18449
2 93870 1 18449
2 93871 1 18449
2 93872 1 18449
2 93873 1 18449
2 93874 1 18449
2 93875 1 18449
2 93876 1 18449
2 93877 1 18449
2 93878 1 18449
2 93879 1 18449
2 93880 1 18449
2 93881 1 18449
2 93882 1 18449
2 93883 1 18449
2 93884 1 18449
2 93885 1 18449
2 93886 1 18449
2 93887 1 18449
2 93888 1 18449
2 93889 1 18449
2 93890 1 18450
2 93891 1 18450
2 93892 1 18450
2 93893 1 18450
2 93894 1 18450
2 93895 1 18450
2 93896 1 18450
2 93897 1 18450
2 93898 1 18450
2 93899 1 18450
2 93900 1 18450
2 93901 1 18450
2 93902 1 18450
2 93903 1 18450
2 93904 1 18450
2 93905 1 18450
2 93906 1 18450
2 93907 1 18450
2 93908 1 18450
2 93909 1 18450
2 93910 1 18450
2 93911 1 18450
2 93912 1 18450
2 93913 1 18450
2 93914 1 18450
2 93915 1 18450
2 93916 1 18450
2 93917 1 18450
2 93918 1 18450
2 93919 1 18450
2 93920 1 18450
2 93921 1 18450
2 93922 1 18450
2 93923 1 18450
2 93924 1 18450
2 93925 1 18450
2 93926 1 18451
2 93927 1 18451
2 93928 1 18451
2 93929 1 18451
2 93930 1 18452
2 93931 1 18452
2 93932 1 18453
2 93933 1 18453
2 93934 1 18453
2 93935 1 18454
2 93936 1 18454
2 93937 1 18455
2 93938 1 18455
2 93939 1 18455
2 93940 1 18455
2 93941 1 18455
2 93942 1 18455
2 93943 1 18459
2 93944 1 18459
2 93945 1 18462
2 93946 1 18462
2 93947 1 18462
2 93948 1 18462
2 93949 1 18462
2 93950 1 18462
2 93951 1 18462
2 93952 1 18462
2 93953 1 18462
2 93954 1 18469
2 93955 1 18469
2 93956 1 18475
2 93957 1 18475
2 93958 1 18483
2 93959 1 18483
2 93960 1 18491
2 93961 1 18491
2 93962 1 18491
2 93963 1 18492
2 93964 1 18492
2 93965 1 18492
2 93966 1 18492
2 93967 1 18492
2 93968 1 18499
2 93969 1 18499
2 93970 1 18502
2 93971 1 18502
2 93972 1 18504
2 93973 1 18504
2 93974 1 18504
2 93975 1 18504
2 93976 1 18504
2 93977 1 18504
2 93978 1 18504
2 93979 1 18504
2 93980 1 18507
2 93981 1 18507
2 93982 1 18514
2 93983 1 18514
2 93984 1 18527
2 93985 1 18527
2 93986 1 18527
2 93987 1 18532
2 93988 1 18532
2 93989 1 18550
2 93990 1 18550
2 93991 1 18550
2 93992 1 18554
2 93993 1 18554
2 93994 1 18592
2 93995 1 18592
2 93996 1 18612
2 93997 1 18612
2 93998 1 18614
2 93999 1 18614
2 94000 1 18614
2 94001 1 18614
2 94002 1 18614
2 94003 1 18616
2 94004 1 18616
2 94005 1 18617
2 94006 1 18617
2 94007 1 18625
2 94008 1 18625
2 94009 1 18625
2 94010 1 18625
2 94011 1 18627
2 94012 1 18627
2 94013 1 18628
2 94014 1 18628
2 94015 1 18633
2 94016 1 18633
2 94017 1 18636
2 94018 1 18636
2 94019 1 18636
2 94020 1 18636
2 94021 1 18636
2 94022 1 18645
2 94023 1 18645
2 94024 1 18645
2 94025 1 18645
2 94026 1 18645
2 94027 1 18645
2 94028 1 18645
2 94029 1 18645
2 94030 1 18645
2 94031 1 18645
2 94032 1 18645
2 94033 1 18646
2 94034 1 18646
2 94035 1 18646
2 94036 1 18646
2 94037 1 18665
2 94038 1 18665
2 94039 1 18665
2 94040 1 18666
2 94041 1 18666
2 94042 1 18666
2 94043 1 18666
2 94044 1 18667
2 94045 1 18667
2 94046 1 18677
2 94047 1 18677
2 94048 1 18677
2 94049 1 18677
2 94050 1 18677
2 94051 1 18677
2 94052 1 18677
2 94053 1 18677
2 94054 1 18677
2 94055 1 18677
2 94056 1 18677
2 94057 1 18679
2 94058 1 18679
2 94059 1 18679
2 94060 1 18698
2 94061 1 18698
2 94062 1 18718
2 94063 1 18718
2 94064 1 18720
2 94065 1 18720
2 94066 1 18725
2 94067 1 18725
2 94068 1 18725
2 94069 1 18725
2 94070 1 18725
2 94071 1 18725
2 94072 1 18732
2 94073 1 18732
2 94074 1 18740
2 94075 1 18740
2 94076 1 18743
2 94077 1 18743
2 94078 1 18744
2 94079 1 18744
2 94080 1 18745
2 94081 1 18745
2 94082 1 18749
2 94083 1 18749
2 94084 1 18765
2 94085 1 18765
2 94086 1 18765
2 94087 1 18772
2 94088 1 18772
2 94089 1 18772
2 94090 1 18772
2 94091 1 18772
2 94092 1 18787
2 94093 1 18787
2 94094 1 18788
2 94095 1 18788
2 94096 1 18802
2 94097 1 18802
2 94098 1 18802
2 94099 1 18803
2 94100 1 18803
2 94101 1 18804
2 94102 1 18804
2 94103 1 18808
2 94104 1 18808
2 94105 1 18812
2 94106 1 18812
2 94107 1 18813
2 94108 1 18813
2 94109 1 18819
2 94110 1 18819
2 94111 1 18820
2 94112 1 18820
2 94113 1 18820
2 94114 1 18820
2 94115 1 18820
2 94116 1 18820
2 94117 1 18820
2 94118 1 18820
2 94119 1 18820
2 94120 1 18820
2 94121 1 18820
2 94122 1 18820
2 94123 1 18820
2 94124 1 18820
2 94125 1 18820
2 94126 1 18820
2 94127 1 18820
2 94128 1 18820
2 94129 1 18820
2 94130 1 18820
2 94131 1 18820
2 94132 1 18820
2 94133 1 18820
2 94134 1 18820
2 94135 1 18820
2 94136 1 18820
2 94137 1 18820
2 94138 1 18820
2 94139 1 18820
2 94140 1 18820
2 94141 1 18821
2 94142 1 18821
2 94143 1 18823
2 94144 1 18823
2 94145 1 18823
2 94146 1 18826
2 94147 1 18826
2 94148 1 18826
2 94149 1 18826
2 94150 1 18836
2 94151 1 18836
2 94152 1 18836
2 94153 1 18837
2 94154 1 18837
2 94155 1 18847
2 94156 1 18847
2 94157 1 18847
2 94158 1 18848
2 94159 1 18848
2 94160 1 18856
2 94161 1 18856
2 94162 1 18890
2 94163 1 18890
2 94164 1 18891
2 94165 1 18891
2 94166 1 18897
2 94167 1 18897
2 94168 1 18907
2 94169 1 18907
2 94170 1 18915
2 94171 1 18915
2 94172 1 18915
2 94173 1 18938
2 94174 1 18938
2 94175 1 18958
2 94176 1 18958
2 94177 1 18959
2 94178 1 18959
2 94179 1 18980
2 94180 1 18980
2 94181 1 18986
2 94182 1 18986
2 94183 1 18997
2 94184 1 18997
2 94185 1 18997
2 94186 1 18997
2 94187 1 18998
2 94188 1 18998
2 94189 1 18998
2 94190 1 18998
2 94191 1 18998
2 94192 1 19017
2 94193 1 19017
2 94194 1 19018
2 94195 1 19018
2 94196 1 19025
2 94197 1 19025
2 94198 1 19025
2 94199 1 19062
2 94200 1 19062
2 94201 1 19062
2 94202 1 19062
2 94203 1 19066
2 94204 1 19066
2 94205 1 19066
2 94206 1 19066
2 94207 1 19066
2 94208 1 19066
2 94209 1 19066
2 94210 1 19066
2 94211 1 19066
2 94212 1 19066
2 94213 1 19066
2 94214 1 19066
2 94215 1 19066
2 94216 1 19066
2 94217 1 19066
2 94218 1 19074
2 94219 1 19074
2 94220 1 19085
2 94221 1 19085
2 94222 1 19110
2 94223 1 19110
2 94224 1 19110
2 94225 1 19116
2 94226 1 19116
2 94227 1 19121
2 94228 1 19121
2 94229 1 19123
2 94230 1 19123
2 94231 1 19136
2 94232 1 19136
2 94233 1 19136
2 94234 1 19136
2 94235 1 19136
2 94236 1 19136
2 94237 1 19136
2 94238 1 19136
2 94239 1 19136
2 94240 1 19145
2 94241 1 19145
2 94242 1 19154
2 94243 1 19154
2 94244 1 19154
2 94245 1 19158
2 94246 1 19158
2 94247 1 19178
2 94248 1 19178
2 94249 1 19178
2 94250 1 19180
2 94251 1 19180
2 94252 1 19192
2 94253 1 19192
2 94254 1 19199
2 94255 1 19199
2 94256 1 19204
2 94257 1 19204
2 94258 1 19204
2 94259 1 19204
2 94260 1 19205
2 94261 1 19205
2 94262 1 19228
2 94263 1 19228
2 94264 1 19231
2 94265 1 19231
2 94266 1 19232
2 94267 1 19232
2 94268 1 19234
2 94269 1 19234
2 94270 1 19234
2 94271 1 19234
2 94272 1 19238
2 94273 1 19238
2 94274 1 19238
2 94275 1 19238
2 94276 1 19238
2 94277 1 19238
2 94278 1 19238
2 94279 1 19241
2 94280 1 19241
2 94281 1 19257
2 94282 1 19257
2 94283 1 19258
2 94284 1 19258
2 94285 1 19258
2 94286 1 19282
2 94287 1 19282
2 94288 1 19282
2 94289 1 19282
2 94290 1 19283
2 94291 1 19283
2 94292 1 19288
2 94293 1 19288
2 94294 1 19288
2 94295 1 19300
2 94296 1 19300
2 94297 1 19300
2 94298 1 19311
2 94299 1 19311
2 94300 1 19314
2 94301 1 19314
2 94302 1 19314
2 94303 1 19321
2 94304 1 19321
2 94305 1 19331
2 94306 1 19331
2 94307 1 19337
2 94308 1 19337
2 94309 1 19344
2 94310 1 19344
2 94311 1 19372
2 94312 1 19372
2 94313 1 19372
2 94314 1 19385
2 94315 1 19385
2 94316 1 19405
2 94317 1 19405
2 94318 1 19408
2 94319 1 19408
2 94320 1 19409
2 94321 1 19409
2 94322 1 19409
2 94323 1 19409
2 94324 1 19409
2 94325 1 19409
2 94326 1 19423
2 94327 1 19423
2 94328 1 19443
2 94329 1 19443
2 94330 1 19455
2 94331 1 19455
2 94332 1 19458
2 94333 1 19458
2 94334 1 19484
2 94335 1 19484
2 94336 1 19484
2 94337 1 19484
2 94338 1 19484
2 94339 1 19484
2 94340 1 19484
2 94341 1 19497
2 94342 1 19497
2 94343 1 19497
2 94344 1 19497
2 94345 1 19499
2 94346 1 19499
2 94347 1 19510
2 94348 1 19510
2 94349 1 19539
2 94350 1 19539
2 94351 1 19539
2 94352 1 19539
2 94353 1 19539
2 94354 1 19539
2 94355 1 19539
2 94356 1 19539
2 94357 1 19539
2 94358 1 19539
2 94359 1 19539
2 94360 1 19539
2 94361 1 19539
2 94362 1 19539
2 94363 1 19539
2 94364 1 19539
2 94365 1 19539
2 94366 1 19539
2 94367 1 19539
2 94368 1 19539
2 94369 1 19539
2 94370 1 19539
2 94371 1 19539
2 94372 1 19539
2 94373 1 19539
2 94374 1 19539
2 94375 1 19539
2 94376 1 19539
2 94377 1 19539
2 94378 1 19539
2 94379 1 19539
2 94380 1 19539
2 94381 1 19539
2 94382 1 19539
2 94383 1 19539
2 94384 1 19539
2 94385 1 19539
2 94386 1 19539
2 94387 1 19539
2 94388 1 19539
2 94389 1 19539
2 94390 1 19539
2 94391 1 19539
2 94392 1 19539
2 94393 1 19540
2 94394 1 19540
2 94395 1 19540
2 94396 1 19540
2 94397 1 19540
2 94398 1 19540
2 94399 1 19540
2 94400 1 19540
2 94401 1 19540
2 94402 1 19540
2 94403 1 19540
2 94404 1 19540
2 94405 1 19540
2 94406 1 19540
2 94407 1 19540
2 94408 1 19540
2 94409 1 19540
2 94410 1 19542
2 94411 1 19542
2 94412 1 19555
2 94413 1 19555
2 94414 1 19579
2 94415 1 19579
2 94416 1 19579
2 94417 1 19579
2 94418 1 19579
2 94419 1 19580
2 94420 1 19580
2 94421 1 19580
2 94422 1 19594
2 94423 1 19594
2 94424 1 19594
2 94425 1 19609
2 94426 1 19609
2 94427 1 19620
2 94428 1 19620
2 94429 1 19620
2 94430 1 19622
2 94431 1 19622
2 94432 1 19622
2 94433 1 19622
2 94434 1 19622
2 94435 1 19623
2 94436 1 19623
2 94437 1 19623
2 94438 1 19623
2 94439 1 19631
2 94440 1 19631
2 94441 1 19634
2 94442 1 19634
2 94443 1 19636
2 94444 1 19636
2 94445 1 19645
2 94446 1 19645
2 94447 1 19645
2 94448 1 19648
2 94449 1 19648
2 94450 1 19648
2 94451 1 19648
2 94452 1 19648
2 94453 1 19648
2 94454 1 19657
2 94455 1 19657
2 94456 1 19657
2 94457 1 19657
2 94458 1 19657
2 94459 1 19663
2 94460 1 19663
2 94461 1 19679
2 94462 1 19679
2 94463 1 19696
2 94464 1 19696
2 94465 1 19696
2 94466 1 19696
2 94467 1 19696
2 94468 1 19696
2 94469 1 19696
2 94470 1 19715
2 94471 1 19715
2 94472 1 19717
2 94473 1 19717
2 94474 1 19717
2 94475 1 19717
2 94476 1 19736
2 94477 1 19736
2 94478 1 19737
2 94479 1 19737
2 94480 1 19738
2 94481 1 19738
2 94482 1 19738
2 94483 1 19753
2 94484 1 19753
2 94485 1 19761
2 94486 1 19761
2 94487 1 19769
2 94488 1 19769
2 94489 1 19769
2 94490 1 19772
2 94491 1 19772
2 94492 1 19790
2 94493 1 19790
2 94494 1 19798
2 94495 1 19798
2 94496 1 19798
2 94497 1 19799
2 94498 1 19799
2 94499 1 19799
2 94500 1 19799
2 94501 1 19799
2 94502 1 19818
2 94503 1 19818
2 94504 1 19818
2 94505 1 19818
2 94506 1 19827
2 94507 1 19827
2 94508 1 19827
2 94509 1 19827
2 94510 1 19828
2 94511 1 19828
2 94512 1 19835
2 94513 1 19835
2 94514 1 19853
2 94515 1 19853
2 94516 1 19854
2 94517 1 19854
2 94518 1 19854
2 94519 1 19856
2 94520 1 19856
2 94521 1 19856
2 94522 1 19856
2 94523 1 19857
2 94524 1 19857
2 94525 1 19860
2 94526 1 19860
2 94527 1 19861
2 94528 1 19861
2 94529 1 19861
2 94530 1 19861
2 94531 1 19861
2 94532 1 19861
2 94533 1 19861
2 94534 1 19861
2 94535 1 19866
2 94536 1 19866
2 94537 1 19866
2 94538 1 19885
2 94539 1 19885
2 94540 1 19885
2 94541 1 19886
2 94542 1 19886
2 94543 1 19932
2 94544 1 19932
2 94545 1 19940
2 94546 1 19940
2 94547 1 19940
2 94548 1 19951
2 94549 1 19951
2 94550 1 19952
2 94551 1 19952
2 94552 1 19952
2 94553 1 19997
2 94554 1 19997
2 94555 1 19997
2 94556 1 19997
2 94557 1 20019
2 94558 1 20019
2 94559 1 20019
2 94560 1 20022
2 94561 1 20022
2 94562 1 20026
2 94563 1 20026
2 94564 1 20027
2 94565 1 20027
2 94566 1 20027
2 94567 1 20035
2 94568 1 20035
2 94569 1 20060
2 94570 1 20060
2 94571 1 20062
2 94572 1 20062
2 94573 1 20062
2 94574 1 20062
2 94575 1 20080
2 94576 1 20080
2 94577 1 20081
2 94578 1 20081
2 94579 1 20097
2 94580 1 20097
2 94581 1 20097
2 94582 1 20103
2 94583 1 20103
2 94584 1 20103
2 94585 1 20103
2 94586 1 20104
2 94587 1 20104
2 94588 1 20104
2 94589 1 20134
2 94590 1 20134
2 94591 1 20134
2 94592 1 20134
2 94593 1 20134
2 94594 1 20135
2 94595 1 20135
2 94596 1 20135
2 94597 1 20135
2 94598 1 20135
2 94599 1 20138
2 94600 1 20138
2 94601 1 20138
2 94602 1 20138
2 94603 1 20138
2 94604 1 20138
2 94605 1 20138
2 94606 1 20138
2 94607 1 20138
2 94608 1 20138
2 94609 1 20138
2 94610 1 20138
2 94611 1 20138
2 94612 1 20138
2 94613 1 20138
2 94614 1 20138
2 94615 1 20138
2 94616 1 20138
2 94617 1 20138
2 94618 1 20138
2 94619 1 20139
2 94620 1 20139
2 94621 1 20145
2 94622 1 20145
2 94623 1 20145
2 94624 1 20145
2 94625 1 20146
2 94626 1 20146
2 94627 1 20146
2 94628 1 20154
2 94629 1 20154
2 94630 1 20154
2 94631 1 20154
2 94632 1 20154
2 94633 1 20154
2 94634 1 20154
2 94635 1 20154
2 94636 1 20154
2 94637 1 20154
2 94638 1 20154
2 94639 1 20154
2 94640 1 20154
2 94641 1 20154
2 94642 1 20155
2 94643 1 20155
2 94644 1 20163
2 94645 1 20163
2 94646 1 20173
2 94647 1 20173
2 94648 1 20173
2 94649 1 20173
2 94650 1 20173
2 94651 1 20173
2 94652 1 20179
2 94653 1 20179
2 94654 1 20179
2 94655 1 20179
2 94656 1 20187
2 94657 1 20187
2 94658 1 20188
2 94659 1 20188
2 94660 1 20188
2 94661 1 20208
2 94662 1 20208
2 94663 1 20209
2 94664 1 20209
2 94665 1 20209
2 94666 1 20210
2 94667 1 20210
2 94668 1 20210
2 94669 1 20210
2 94670 1 20222
2 94671 1 20222
2 94672 1 20222
2 94673 1 20229
2 94674 1 20229
2 94675 1 20237
2 94676 1 20237
2 94677 1 20243
2 94678 1 20243
2 94679 1 20243
2 94680 1 20243
2 94681 1 20243
2 94682 1 20243
2 94683 1 20253
2 94684 1 20253
2 94685 1 20272
2 94686 1 20272
2 94687 1 20293
2 94688 1 20293
2 94689 1 20293
2 94690 1 20301
2 94691 1 20301
2 94692 1 20301
2 94693 1 20301
2 94694 1 20301
2 94695 1 20301
2 94696 1 20303
2 94697 1 20303
2 94698 1 20306
2 94699 1 20306
2 94700 1 20307
2 94701 1 20307
2 94702 1 20307
2 94703 1 20307
2 94704 1 20307
2 94705 1 20307
2 94706 1 20307
2 94707 1 20307
2 94708 1 20307
2 94709 1 20307
2 94710 1 20307
2 94711 1 20307
2 94712 1 20307
2 94713 1 20307
2 94714 1 20310
2 94715 1 20310
2 94716 1 20310
2 94717 1 20310
2 94718 1 20310
2 94719 1 20310
2 94720 1 20310
2 94721 1 20311
2 94722 1 20311
2 94723 1 20311
2 94724 1 20311
2 94725 1 20311
2 94726 1 20311
2 94727 1 20311
2 94728 1 20319
2 94729 1 20319
2 94730 1 20320
2 94731 1 20320
2 94732 1 20320
2 94733 1 20320
2 94734 1 20320
2 94735 1 20320
2 94736 1 20320
2 94737 1 20320
2 94738 1 20320
2 94739 1 20320
2 94740 1 20320
2 94741 1 20320
2 94742 1 20320
2 94743 1 20321
2 94744 1 20321
2 94745 1 20321
2 94746 1 20321
2 94747 1 20321
2 94748 1 20321
2 94749 1 20321
2 94750 1 20321
2 94751 1 20321
2 94752 1 20321
2 94753 1 20321
2 94754 1 20335
2 94755 1 20335
2 94756 1 20336
2 94757 1 20336
2 94758 1 20336
2 94759 1 20336
2 94760 1 20336
2 94761 1 20336
2 94762 1 20336
2 94763 1 20344
2 94764 1 20344
2 94765 1 20344
2 94766 1 20344
2 94767 1 20344
2 94768 1 20344
2 94769 1 20344
2 94770 1 20344
2 94771 1 20345
2 94772 1 20345
2 94773 1 20346
2 94774 1 20346
2 94775 1 20346
2 94776 1 20358
2 94777 1 20358
2 94778 1 20360
2 94779 1 20360
2 94780 1 20364
2 94781 1 20364
2 94782 1 20365
2 94783 1 20365
2 94784 1 20365
2 94785 1 20365
2 94786 1 20365
2 94787 1 20365
2 94788 1 20366
2 94789 1 20366
2 94790 1 20366
2 94791 1 20376
2 94792 1 20376
2 94793 1 20379
2 94794 1 20379
2 94795 1 20379
2 94796 1 20399
2 94797 1 20399
2 94798 1 20402
2 94799 1 20402
2 94800 1 20418
2 94801 1 20418
2 94802 1 20418
2 94803 1 20425
2 94804 1 20425
2 94805 1 20447
2 94806 1 20447
2 94807 1 20447
2 94808 1 20459
2 94809 1 20459
2 94810 1 20463
2 94811 1 20463
2 94812 1 20463
2 94813 1 20463
2 94814 1 20495
2 94815 1 20495
2 94816 1 20495
2 94817 1 20495
2 94818 1 20538
2 94819 1 20538
2 94820 1 20538
2 94821 1 20538
2 94822 1 20538
2 94823 1 20538
2 94824 1 20538
2 94825 1 20538
2 94826 1 20538
2 94827 1 20539
2 94828 1 20539
2 94829 1 20539
2 94830 1 20539
2 94831 1 20539
2 94832 1 20540
2 94833 1 20540
2 94834 1 20540
2 94835 1 20540
2 94836 1 20577
2 94837 1 20577
2 94838 1 20578
2 94839 1 20578
2 94840 1 20580
2 94841 1 20580
2 94842 1 20584
2 94843 1 20584
2 94844 1 20593
2 94845 1 20593
2 94846 1 20607
2 94847 1 20607
2 94848 1 20607
2 94849 1 20607
2 94850 1 20607
2 94851 1 20607
2 94852 1 20607
2 94853 1 20607
2 94854 1 20607
2 94855 1 20607
2 94856 1 20607
2 94857 1 20607
2 94858 1 20607
2 94859 1 20621
2 94860 1 20621
2 94861 1 20622
2 94862 1 20622
2 94863 1 20623
2 94864 1 20623
2 94865 1 20623
2 94866 1 20623
2 94867 1 20623
2 94868 1 20624
2 94869 1 20624
2 94870 1 20624
2 94871 1 20626
2 94872 1 20626
2 94873 1 20626
2 94874 1 20626
2 94875 1 20626
2 94876 1 20626
2 94877 1 20626
2 94878 1 20626
2 94879 1 20626
2 94880 1 20626
2 94881 1 20628
2 94882 1 20628
2 94883 1 20628
2 94884 1 20628
2 94885 1 20632
2 94886 1 20632
2 94887 1 20632
2 94888 1 20635
2 94889 1 20635
2 94890 1 20635
2 94891 1 20648
2 94892 1 20648
2 94893 1 20648
2 94894 1 20650
2 94895 1 20650
2 94896 1 20667
2 94897 1 20667
2 94898 1 20667
2 94899 1 20667
2 94900 1 20667
2 94901 1 20667
2 94902 1 20667
2 94903 1 20676
2 94904 1 20676
2 94905 1 20687
2 94906 1 20687
2 94907 1 20689
2 94908 1 20689
2 94909 1 20689
2 94910 1 20692
2 94911 1 20692
2 94912 1 20692
2 94913 1 20692
2 94914 1 20692
2 94915 1 20692
2 94916 1 20692
2 94917 1 20692
2 94918 1 20694
2 94919 1 20694
2 94920 1 20711
2 94921 1 20711
2 94922 1 20738
2 94923 1 20738
2 94924 1 20739
2 94925 1 20739
2 94926 1 20756
2 94927 1 20756
2 94928 1 20777
2 94929 1 20777
2 94930 1 20777
2 94931 1 20800
2 94932 1 20800
2 94933 1 20809
2 94934 1 20809
2 94935 1 20816
2 94936 1 20816
2 94937 1 20816
2 94938 1 20816
2 94939 1 20816
2 94940 1 20816
2 94941 1 20816
2 94942 1 20816
2 94943 1 20816
2 94944 1 20816
2 94945 1 20816
2 94946 1 20816
2 94947 1 20816
2 94948 1 20816
2 94949 1 20816
2 94950 1 20816
2 94951 1 20817
2 94952 1 20817
2 94953 1 20817
2 94954 1 20817
2 94955 1 20820
2 94956 1 20820
2 94957 1 20820
2 94958 1 20829
2 94959 1 20829
2 94960 1 20857
2 94961 1 20857
2 94962 1 20857
2 94963 1 20878
2 94964 1 20878
2 94965 1 20878
2 94966 1 20899
2 94967 1 20899
2 94968 1 20915
2 94969 1 20915
2 94970 1 20916
2 94971 1 20916
2 94972 1 20930
2 94973 1 20930
2 94974 1 20962
2 94975 1 20962
2 94976 1 20972
2 94977 1 20972
2 94978 1 20972
2 94979 1 20972
2 94980 1 20972
2 94981 1 20980
2 94982 1 20980
2 94983 1 20980
2 94984 1 20980
2 94985 1 20980
2 94986 1 20983
2 94987 1 20983
2 94988 1 20992
2 94989 1 20992
2 94990 1 21011
2 94991 1 21011
2 94992 1 21022
2 94993 1 21022
2 94994 1 21022
2 94995 1 21022
2 94996 1 21022
2 94997 1 21022
2 94998 1 21022
2 94999 1 21022
2 95000 1 21022
2 95001 1 21022
2 95002 1 21023
2 95003 1 21023
2 95004 1 21025
2 95005 1 21025
2 95006 1 21031
2 95007 1 21031
2 95008 1 21032
2 95009 1 21032
2 95010 1 21032
2 95011 1 21039
2 95012 1 21039
2 95013 1 21056
2 95014 1 21056
2 95015 1 21056
2 95016 1 21056
2 95017 1 21059
2 95018 1 21059
2 95019 1 21062
2 95020 1 21062
2 95021 1 21062
2 95022 1 21062
2 95023 1 21062
2 95024 1 21062
2 95025 1 21062
2 95026 1 21063
2 95027 1 21063
2 95028 1 21070
2 95029 1 21070
2 95030 1 21082
2 95031 1 21082
2 95032 1 21082
2 95033 1 21082
2 95034 1 21093
2 95035 1 21093
2 95036 1 21111
2 95037 1 21111
2 95038 1 21111
2 95039 1 21114
2 95040 1 21114
2 95041 1 21114
2 95042 1 21114
2 95043 1 21114
2 95044 1 21115
2 95045 1 21115
2 95046 1 21115
2 95047 1 21119
2 95048 1 21119
2 95049 1 21119
2 95050 1 21136
2 95051 1 21136
2 95052 1 21136
2 95053 1 21145
2 95054 1 21145
2 95055 1 21151
2 95056 1 21151
2 95057 1 21184
2 95058 1 21184
2 95059 1 21186
2 95060 1 21186
2 95061 1 21186
2 95062 1 21187
2 95063 1 21187
2 95064 1 21190
2 95065 1 21190
2 95066 1 21190
2 95067 1 21213
2 95068 1 21213
2 95069 1 21216
2 95070 1 21216
2 95071 1 21216
2 95072 1 21217
2 95073 1 21217
2 95074 1 21237
2 95075 1 21237
2 95076 1 21244
2 95077 1 21244
2 95078 1 21245
2 95079 1 21245
2 95080 1 21246
2 95081 1 21246
2 95082 1 21255
2 95083 1 21255
2 95084 1 21257
2 95085 1 21257
2 95086 1 21292
2 95087 1 21292
2 95088 1 21323
2 95089 1 21323
2 95090 1 21323
2 95091 1 21354
2 95092 1 21354
2 95093 1 21354
2 95094 1 21354
2 95095 1 21354
2 95096 1 21354
2 95097 1 21354
2 95098 1 21354
2 95099 1 21354
2 95100 1 21362
2 95101 1 21362
2 95102 1 21362
2 95103 1 21362
2 95104 1 21362
2 95105 1 21362
2 95106 1 21371
2 95107 1 21371
2 95108 1 21371
2 95109 1 21371
2 95110 1 21371
2 95111 1 21371
2 95112 1 21371
2 95113 1 21371
2 95114 1 21371
2 95115 1 21371
2 95116 1 21371
2 95117 1 21371
2 95118 1 21372
2 95119 1 21372
2 95120 1 21372
2 95121 1 21372
2 95122 1 21380
2 95123 1 21380
2 95124 1 21391
2 95125 1 21391
2 95126 1 21391
2 95127 1 21392
2 95128 1 21392
2 95129 1 21392
2 95130 1 21392
2 95131 1 21402
2 95132 1 21402
2 95133 1 21402
2 95134 1 21402
2 95135 1 21409
2 95136 1 21409
2 95137 1 21425
2 95138 1 21425
2 95139 1 21434
2 95140 1 21434
2 95141 1 21443
2 95142 1 21443
2 95143 1 21443
2 95144 1 21446
2 95145 1 21446
2 95146 1 21446
2 95147 1 21446
2 95148 1 21446
2 95149 1 21446
2 95150 1 21446
2 95151 1 21446
2 95152 1 21446
2 95153 1 21446
2 95154 1 21446
2 95155 1 21447
2 95156 1 21447
2 95157 1 21447
2 95158 1 21456
2 95159 1 21456
2 95160 1 21464
2 95161 1 21464
2 95162 1 21464
2 95163 1 21476
2 95164 1 21476
2 95165 1 21476
2 95166 1 21476
2 95167 1 21476
2 95168 1 21476
2 95169 1 21476
2 95170 1 21486
2 95171 1 21486
2 95172 1 21486
2 95173 1 21486
2 95174 1 21487
2 95175 1 21487
2 95176 1 21488
2 95177 1 21488
2 95178 1 21489
2 95179 1 21489
2 95180 1 21490
2 95181 1 21490
2 95182 1 21490
2 95183 1 21490
2 95184 1 21491
2 95185 1 21491
2 95186 1 21491
2 95187 1 21501
2 95188 1 21501
2 95189 1 21501
2 95190 1 21502
2 95191 1 21502
2 95192 1 21502
2 95193 1 21503
2 95194 1 21503
2 95195 1 21503
2 95196 1 21503
2 95197 1 21503
2 95198 1 21503
2 95199 1 21519
2 95200 1 21519
2 95201 1 21544
2 95202 1 21544
2 95203 1 21544
2 95204 1 21544
2 95205 1 21544
2 95206 1 21554
2 95207 1 21554
2 95208 1 21569
2 95209 1 21569
2 95210 1 21569
2 95211 1 21569
2 95212 1 21570
2 95213 1 21570
2 95214 1 21573
2 95215 1 21573
2 95216 1 21576
2 95217 1 21576
2 95218 1 21576
2 95219 1 21594
2 95220 1 21594
2 95221 1 21594
2 95222 1 21646
2 95223 1 21646
2 95224 1 21646
2 95225 1 21654
2 95226 1 21654
2 95227 1 21654
2 95228 1 21655
2 95229 1 21655
2 95230 1 21657
2 95231 1 21657
2 95232 1 21673
2 95233 1 21673
2 95234 1 21673
2 95235 1 21687
2 95236 1 21687
2 95237 1 21697
2 95238 1 21697
2 95239 1 21716
2 95240 1 21716
2 95241 1 21724
2 95242 1 21724
2 95243 1 21724
2 95244 1 21725
2 95245 1 21725
2 95246 1 21725
2 95247 1 21730
2 95248 1 21730
2 95249 1 21735
2 95250 1 21735
2 95251 1 21735
2 95252 1 21735
2 95253 1 21735
2 95254 1 21735
2 95255 1 21735
2 95256 1 21736
2 95257 1 21736
2 95258 1 21736
2 95259 1 21736
2 95260 1 21736
2 95261 1 21736
2 95262 1 21736
2 95263 1 21736
2 95264 1 21746
2 95265 1 21746
2 95266 1 21746
2 95267 1 21755
2 95268 1 21755
2 95269 1 21771
2 95270 1 21771
2 95271 1 21771
2 95272 1 21778
2 95273 1 21778
2 95274 1 21788
2 95275 1 21788
2 95276 1 21788
2 95277 1 21788
2 95278 1 21789
2 95279 1 21789
2 95280 1 21802
2 95281 1 21802
2 95282 1 21802
2 95283 1 21802
2 95284 1 21802
2 95285 1 21802
2 95286 1 21802
2 95287 1 21802
2 95288 1 21802
2 95289 1 21802
2 95290 1 21807
2 95291 1 21807
2 95292 1 21807
2 95293 1 21807
2 95294 1 21807
2 95295 1 21807
2 95296 1 21808
2 95297 1 21808
2 95298 1 21816
2 95299 1 21816
2 95300 1 21816
2 95301 1 21817
2 95302 1 21817
2 95303 1 21817
2 95304 1 21817
2 95305 1 21817
2 95306 1 21817
2 95307 1 21817
2 95308 1 21818
2 95309 1 21818
2 95310 1 21818
2 95311 1 21819
2 95312 1 21819
2 95313 1 21819
2 95314 1 21819
2 95315 1 21819
2 95316 1 21819
2 95317 1 21819
2 95318 1 21819
2 95319 1 21819
2 95320 1 21819
2 95321 1 21819
2 95322 1 21833
2 95323 1 21833
2 95324 1 21854
2 95325 1 21854
2 95326 1 21855
2 95327 1 21855
2 95328 1 21855
2 95329 1 21878
2 95330 1 21878
2 95331 1 21878
2 95332 1 21878
2 95333 1 21892
2 95334 1 21892
2 95335 1 21894
2 95336 1 21894
2 95337 1 21894
2 95338 1 21894
2 95339 1 21894
2 95340 1 21894
2 95341 1 21894
2 95342 1 21894
2 95343 1 21894
2 95344 1 21894
2 95345 1 21894
2 95346 1 21894
2 95347 1 21894
2 95348 1 21894
2 95349 1 21894
2 95350 1 21894
2 95351 1 21894
2 95352 1 21894
2 95353 1 21894
2 95354 1 21913
2 95355 1 21913
2 95356 1 21953
2 95357 1 21953
2 95358 1 21953
2 95359 1 21958
2 95360 1 21958
2 95361 1 21959
2 95362 1 21959
2 95363 1 22019
2 95364 1 22019
2 95365 1 22019
2 95366 1 22019
2 95367 1 22027
2 95368 1 22027
2 95369 1 22027
2 95370 1 22027
2 95371 1 22027
2 95372 1 22027
2 95373 1 22028
2 95374 1 22028
2 95375 1 22029
2 95376 1 22029
2 95377 1 22029
2 95378 1 22030
2 95379 1 22030
2 95380 1 22030
2 95381 1 22034
2 95382 1 22034
2 95383 1 22034
2 95384 1 22046
2 95385 1 22046
2 95386 1 22049
2 95387 1 22049
2 95388 1 22049
2 95389 1 22049
2 95390 1 22049
2 95391 1 22049
2 95392 1 22049
2 95393 1 22051
2 95394 1 22051
2 95395 1 22051
2 95396 1 22051
2 95397 1 22051
2 95398 1 22051
2 95399 1 22066
2 95400 1 22066
2 95401 1 22081
2 95402 1 22081
2 95403 1 22090
2 95404 1 22090
2 95405 1 22102
2 95406 1 22102
2 95407 1 22105
2 95408 1 22105
2 95409 1 22105
2 95410 1 22105
2 95411 1 22105
2 95412 1 22105
2 95413 1 22105
2 95414 1 22132
2 95415 1 22132
2 95416 1 22132
2 95417 1 22132
2 95418 1 22132
2 95419 1 22133
2 95420 1 22133
2 95421 1 22150
2 95422 1 22150
2 95423 1 22157
2 95424 1 22157
2 95425 1 22157
2 95426 1 22157
2 95427 1 22157
2 95428 1 22157
2 95429 1 22157
2 95430 1 22157
2 95431 1 22159
2 95432 1 22159
2 95433 1 22162
2 95434 1 22162
2 95435 1 22173
2 95436 1 22173
2 95437 1 22181
2 95438 1 22181
2 95439 1 22182
2 95440 1 22182
2 95441 1 22184
2 95442 1 22184
2 95443 1 22189
2 95444 1 22189
2 95445 1 22189
2 95446 1 22189
2 95447 1 22189
2 95448 1 22189
2 95449 1 22189
2 95450 1 22189
2 95451 1 22190
2 95452 1 22190
2 95453 1 22190
2 95454 1 22199
2 95455 1 22199
2 95456 1 22228
2 95457 1 22228
2 95458 1 22245
2 95459 1 22245
2 95460 1 22245
2 95461 1 22245
2 95462 1 22303
2 95463 1 22303
2 95464 1 22304
2 95465 1 22304
2 95466 1 22304
2 95467 1 22314
2 95468 1 22314
2 95469 1 22314
2 95470 1 22334
2 95471 1 22334
2 95472 1 22335
2 95473 1 22335
2 95474 1 22335
2 95475 1 22349
2 95476 1 22349
2 95477 1 22349
2 95478 1 22349
2 95479 1 22359
2 95480 1 22359
2 95481 1 22359
2 95482 1 22359
2 95483 1 22367
2 95484 1 22367
2 95485 1 22367
2 95486 1 22367
2 95487 1 22368
2 95488 1 22368
2 95489 1 22396
2 95490 1 22396
2 95491 1 22421
2 95492 1 22421
2 95493 1 22421
2 95494 1 22424
2 95495 1 22424
2 95496 1 22424
2 95497 1 22454
2 95498 1 22454
2 95499 1 22462
2 95500 1 22462
2 95501 1 22462
2 95502 1 22462
2 95503 1 22463
2 95504 1 22463
2 95505 1 22465
2 95506 1 22465
2 95507 1 22465
2 95508 1 22465
2 95509 1 22475
2 95510 1 22475
2 95511 1 22483
2 95512 1 22483
2 95513 1 22494
2 95514 1 22494
2 95515 1 22495
2 95516 1 22495
2 95517 1 22503
2 95518 1 22503
2 95519 1 22504
2 95520 1 22504
2 95521 1 22508
2 95522 1 22508
2 95523 1 22521
2 95524 1 22521
2 95525 1 22532
2 95526 1 22532
2 95527 1 22546
2 95528 1 22546
2 95529 1 22554
2 95530 1 22554
2 95531 1 22556
2 95532 1 22556
2 95533 1 22585
2 95534 1 22585
2 95535 1 22616
2 95536 1 22616
2 95537 1 22631
2 95538 1 22631
2 95539 1 22664
2 95540 1 22664
2 95541 1 22686
2 95542 1 22686
2 95543 1 22686
2 95544 1 22687
2 95545 1 22687
2 95546 1 22687
2 95547 1 22687
2 95548 1 22687
2 95549 1 22700
2 95550 1 22700
2 95551 1 22727
2 95552 1 22727
2 95553 1 22727
2 95554 1 22731
2 95555 1 22731
2 95556 1 22739
2 95557 1 22739
2 95558 1 22739
2 95559 1 22754
2 95560 1 22754
2 95561 1 22762
2 95562 1 22762
2 95563 1 22773
2 95564 1 22773
2 95565 1 22773
2 95566 1 22773
2 95567 1 22773
2 95568 1 22774
2 95569 1 22774
2 95570 1 22783
2 95571 1 22783
2 95572 1 22784
2 95573 1 22784
2 95574 1 22789
2 95575 1 22789
2 95576 1 22806
2 95577 1 22806
2 95578 1 22814
2 95579 1 22814
2 95580 1 22819
2 95581 1 22819
2 95582 1 22837
2 95583 1 22837
2 95584 1 22858
2 95585 1 22858
2 95586 1 22858
2 95587 1 22859
2 95588 1 22859
2 95589 1 22859
2 95590 1 22881
2 95591 1 22881
2 95592 1 22881
2 95593 1 22881
2 95594 1 22883
2 95595 1 22883
2 95596 1 22888
2 95597 1 22888
2 95598 1 22888
2 95599 1 22888
2 95600 1 22888
2 95601 1 22898
2 95602 1 22898
2 95603 1 22929
2 95604 1 22929
2 95605 1 22931
2 95606 1 22931
2 95607 1 22947
2 95608 1 22947
2 95609 1 22947
2 95610 1 22965
2 95611 1 22965
2 95612 1 22973
2 95613 1 22973
2 95614 1 22978
2 95615 1 22978
2 95616 1 22990
2 95617 1 22990
2 95618 1 23001
2 95619 1 23001
2 95620 1 23009
2 95621 1 23009
2 95622 1 23009
2 95623 1 23009
2 95624 1 23009
2 95625 1 23010
2 95626 1 23010
2 95627 1 23012
2 95628 1 23012
2 95629 1 23023
2 95630 1 23023
2 95631 1 23023
2 95632 1 23029
2 95633 1 23029
2 95634 1 23034
2 95635 1 23034
2 95636 1 23047
2 95637 1 23047
2 95638 1 23080
2 95639 1 23080
2 95640 1 23081
2 95641 1 23081
2 95642 1 23081
2 95643 1 23081
2 95644 1 23086
2 95645 1 23086
2 95646 1 23086
2 95647 1 23086
2 95648 1 23089
2 95649 1 23089
2 95650 1 23090
2 95651 1 23090
2 95652 1 23090
2 95653 1 23098
2 95654 1 23098
2 95655 1 23108
2 95656 1 23108
2 95657 1 23117
2 95658 1 23117
2 95659 1 23117
2 95660 1 23117
2 95661 1 23118
2 95662 1 23118
2 95663 1 23118
2 95664 1 23118
2 95665 1 23122
2 95666 1 23122
2 95667 1 23122
2 95668 1 23122
2 95669 1 23122
2 95670 1 23129
2 95671 1 23129
2 95672 1 23175
2 95673 1 23175
2 95674 1 23196
2 95675 1 23196
2 95676 1 23196
2 95677 1 23200
2 95678 1 23200
2 95679 1 23201
2 95680 1 23201
2 95681 1 23207
2 95682 1 23207
2 95683 1 23207
2 95684 1 23207
2 95685 1 23207
2 95686 1 23208
2 95687 1 23208
2 95688 1 23208
2 95689 1 23208
2 95690 1 23222
2 95691 1 23222
2 95692 1 23244
2 95693 1 23244
2 95694 1 23287
2 95695 1 23287
2 95696 1 23315
2 95697 1 23315
2 95698 1 23317
2 95699 1 23317
2 95700 1 23319
2 95701 1 23319
2 95702 1 23321
2 95703 1 23321
2 95704 1 23328
2 95705 1 23328
2 95706 1 23328
2 95707 1 23329
2 95708 1 23329
2 95709 1 23329
2 95710 1 23329
2 95711 1 23329
2 95712 1 23329
2 95713 1 23329
2 95714 1 23329
2 95715 1 23329
2 95716 1 23329
2 95717 1 23330
2 95718 1 23330
2 95719 1 23338
2 95720 1 23338
2 95721 1 23348
2 95722 1 23348
2 95723 1 23352
2 95724 1 23352
2 95725 1 23354
2 95726 1 23354
2 95727 1 23372
2 95728 1 23372
2 95729 1 23375
2 95730 1 23375
2 95731 1 23383
2 95732 1 23383
2 95733 1 23389
2 95734 1 23389
2 95735 1 23390
2 95736 1 23390
2 95737 1 23390
2 95738 1 23407
2 95739 1 23407
2 95740 1 23410
2 95741 1 23410
2 95742 1 23410
2 95743 1 23411
2 95744 1 23411
2 95745 1 23421
2 95746 1 23421
2 95747 1 23424
2 95748 1 23424
2 95749 1 23433
2 95750 1 23433
2 95751 1 23448
2 95752 1 23448
2 95753 1 23451
2 95754 1 23451
2 95755 1 23461
2 95756 1 23461
2 95757 1 23515
2 95758 1 23515
2 95759 1 23516
2 95760 1 23516
2 95761 1 23520
2 95762 1 23520
2 95763 1 23529
2 95764 1 23529
2 95765 1 23529
2 95766 1 23529
2 95767 1 23531
2 95768 1 23531
2 95769 1 23545
2 95770 1 23545
2 95771 1 23552
2 95772 1 23552
2 95773 1 23580
2 95774 1 23580
2 95775 1 23608
2 95776 1 23608
2 95777 1 23608
2 95778 1 23608
2 95779 1 23608
2 95780 1 23608
2 95781 1 23609
2 95782 1 23609
2 95783 1 23610
2 95784 1 23610
2 95785 1 23615
2 95786 1 23615
2 95787 1 23618
2 95788 1 23618
2 95789 1 23632
2 95790 1 23632
2 95791 1 23633
2 95792 1 23633
2 95793 1 23633
2 95794 1 23634
2 95795 1 23634
2 95796 1 23635
2 95797 1 23635
2 95798 1 23636
2 95799 1 23636
2 95800 1 23650
2 95801 1 23650
2 95802 1 23650
2 95803 1 23650
2 95804 1 23654
2 95805 1 23654
2 95806 1 23654
2 95807 1 23666
2 95808 1 23666
2 95809 1 23666
2 95810 1 23684
2 95811 1 23684
2 95812 1 23697
2 95813 1 23697
2 95814 1 23710
2 95815 1 23710
2 95816 1 23721
2 95817 1 23721
2 95818 1 23721
2 95819 1 23747
2 95820 1 23747
2 95821 1 23765
2 95822 1 23765
2 95823 1 23765
2 95824 1 23778
2 95825 1 23778
2 95826 1 23778
2 95827 1 23778
2 95828 1 23778
2 95829 1 23779
2 95830 1 23779
2 95831 1 23786
2 95832 1 23786
2 95833 1 23797
2 95834 1 23797
2 95835 1 23797
2 95836 1 23797
2 95837 1 23797
2 95838 1 23800
2 95839 1 23800
2 95840 1 23800
2 95841 1 23800
2 95842 1 23801
2 95843 1 23801
2 95844 1 23801
2 95845 1 23843
2 95846 1 23843
2 95847 1 23856
2 95848 1 23856
2 95849 1 23891
2 95850 1 23891
2 95851 1 23891
2 95852 1 23902
2 95853 1 23902
2 95854 1 23902
2 95855 1 23902
2 95856 1 23927
2 95857 1 23927
2 95858 1 23927
2 95859 1 23945
2 95860 1 23945
2 95861 1 23946
2 95862 1 23946
2 95863 1 23946
2 95864 1 23946
2 95865 1 23946
2 95866 1 23946
2 95867 1 23989
2 95868 1 23989
2 95869 1 23989
2 95870 1 23989
2 95871 1 23989
2 95872 1 23991
2 95873 1 23991
2 95874 1 24005
2 95875 1 24005
2 95876 1 24005
2 95877 1 24008
2 95878 1 24008
2 95879 1 24008
2 95880 1 24008
2 95881 1 24008
2 95882 1 24008
2 95883 1 24008
2 95884 1 24009
2 95885 1 24009
2 95886 1 24009
2 95887 1 24009
2 95888 1 24009
2 95889 1 24028
2 95890 1 24028
2 95891 1 24029
2 95892 1 24029
2 95893 1 24044
2 95894 1 24044
2 95895 1 24047
2 95896 1 24047
2 95897 1 24075
2 95898 1 24075
2 95899 1 24075
2 95900 1 24075
2 95901 1 24075
2 95902 1 24075
2 95903 1 24076
2 95904 1 24076
2 95905 1 24076
2 95906 1 24077
2 95907 1 24077
2 95908 1 24080
2 95909 1 24080
2 95910 1 24086
2 95911 1 24086
2 95912 1 24096
2 95913 1 24096
2 95914 1 24096
2 95915 1 24107
2 95916 1 24107
2 95917 1 24108
2 95918 1 24108
2 95919 1 24117
2 95920 1 24117
2 95921 1 24117
2 95922 1 24132
2 95923 1 24132
2 95924 1 24176
2 95925 1 24176
2 95926 1 24177
2 95927 1 24177
2 95928 1 24203
2 95929 1 24203
2 95930 1 24203
2 95931 1 24204
2 95932 1 24204
2 95933 1 24204
2 95934 1 24232
2 95935 1 24232
2 95936 1 24237
2 95937 1 24237
2 95938 1 24247
2 95939 1 24247
2 95940 1 24247
2 95941 1 24248
2 95942 1 24248
2 95943 1 24261
2 95944 1 24261
2 95945 1 24271
2 95946 1 24271
2 95947 1 24278
2 95948 1 24278
2 95949 1 24281
2 95950 1 24281
2 95951 1 24281
2 95952 1 24281
2 95953 1 24282
2 95954 1 24282
2 95955 1 24282
2 95956 1 24282
2 95957 1 24282
2 95958 1 24289
2 95959 1 24289
2 95960 1 24297
2 95961 1 24297
2 95962 1 24298
2 95963 1 24298
2 95964 1 24299
2 95965 1 24299
2 95966 1 24307
2 95967 1 24307
2 95968 1 24322
2 95969 1 24322
2 95970 1 24330
2 95971 1 24330
2 95972 1 24339
2 95973 1 24339
2 95974 1 24340
2 95975 1 24340
2 95976 1 24340
2 95977 1 24340
2 95978 1 24342
2 95979 1 24342
2 95980 1 24342
2 95981 1 24362
2 95982 1 24362
2 95983 1 24363
2 95984 1 24363
2 95985 1 24385
2 95986 1 24385
2 95987 1 24386
2 95988 1 24386
2 95989 1 24386
2 95990 1 24386
2 95991 1 24386
2 95992 1 24386
2 95993 1 24386
2 95994 1 24422
2 95995 1 24422
2 95996 1 24428
2 95997 1 24428
2 95998 1 24432
2 95999 1 24432
2 96000 1 24433
2 96001 1 24433
2 96002 1 24434
2 96003 1 24434
2 96004 1 24456
2 96005 1 24456
2 96006 1 24470
2 96007 1 24470
2 96008 1 24496
2 96009 1 24496
2 96010 1 24550
2 96011 1 24550
2 96012 1 24565
2 96013 1 24565
2 96014 1 24571
2 96015 1 24571
2 96016 1 24607
2 96017 1 24607
2 96018 1 24611
2 96019 1 24611
2 96020 1 24624
2 96021 1 24624
2 96022 1 24637
2 96023 1 24637
2 96024 1 24637
2 96025 1 24648
2 96026 1 24648
2 96027 1 24654
2 96028 1 24654
2 96029 1 24671
2 96030 1 24671
2 96031 1 24679
2 96032 1 24679
2 96033 1 24691
2 96034 1 24691
2 96035 1 24706
2 96036 1 24706
2 96037 1 24746
2 96038 1 24746
2 96039 1 24746
2 96040 1 24746
2 96041 1 24746
2 96042 1 24746
2 96043 1 24746
2 96044 1 24746
2 96045 1 24746
2 96046 1 24746
2 96047 1 24746
2 96048 1 24767
2 96049 1 24767
2 96050 1 24779
2 96051 1 24779
2 96052 1 24780
2 96053 1 24780
2 96054 1 24787
2 96055 1 24787
2 96056 1 24798
2 96057 1 24798
2 96058 1 24817
2 96059 1 24817
2 96060 1 24818
2 96061 1 24818
2 96062 1 24818
2 96063 1 24818
2 96064 1 24818
2 96065 1 24818
2 96066 1 24822
2 96067 1 24822
2 96068 1 24823
2 96069 1 24823
2 96070 1 24823
2 96071 1 24823
2 96072 1 24824
2 96073 1 24824
2 96074 1 24824
2 96075 1 24824
2 96076 1 24824
2 96077 1 24824
2 96078 1 24824
2 96079 1 24833
2 96080 1 24833
2 96081 1 24837
2 96082 1 24837
2 96083 1 24837
2 96084 1 24837
2 96085 1 24837
2 96086 1 24845
2 96087 1 24845
2 96088 1 24845
2 96089 1 24845
2 96090 1 24846
2 96091 1 24846
2 96092 1 24847
2 96093 1 24847
2 96094 1 24847
2 96095 1 24847
2 96096 1 24862
2 96097 1 24862
2 96098 1 24862
2 96099 1 24862
2 96100 1 24862
2 96101 1 24862
2 96102 1 24862
2 96103 1 24862
2 96104 1 24862
2 96105 1 24862
2 96106 1 24862
2 96107 1 24862
2 96108 1 24862
2 96109 1 24871
2 96110 1 24871
2 96111 1 24871
2 96112 1 24871
2 96113 1 24871
2 96114 1 24871
2 96115 1 24880
2 96116 1 24880
2 96117 1 24880
2 96118 1 24880
2 96119 1 24880
2 96120 1 24898
2 96121 1 24898
2 96122 1 24898
2 96123 1 24898
2 96124 1 24898
2 96125 1 24899
2 96126 1 24899
2 96127 1 24926
2 96128 1 24926
2 96129 1 24929
2 96130 1 24929
2 96131 1 24955
2 96132 1 24955
2 96133 1 24955
2 96134 1 24955
2 96135 1 24955
2 96136 1 24955
2 96137 1 24959
2 96138 1 24959
2 96139 1 24959
2 96140 1 24959
2 96141 1 24959
2 96142 1 24959
2 96143 1 24959
2 96144 1 24959
2 96145 1 24959
2 96146 1 24959
2 96147 1 24983
2 96148 1 24983
2 96149 1 24986
2 96150 1 24986
2 96151 1 24990
2 96152 1 24990
2 96153 1 24992
2 96154 1 24992
2 96155 1 24992
2 96156 1 24992
2 96157 1 24992
2 96158 1 25001
2 96159 1 25001
2 96160 1 25001
2 96161 1 25002
2 96162 1 25002
2 96163 1 25019
2 96164 1 25019
2 96165 1 25048
2 96166 1 25048
2 96167 1 25048
2 96168 1 25052
2 96169 1 25052
2 96170 1 25052
2 96171 1 25052
2 96172 1 25052
2 96173 1 25064
2 96174 1 25064
2 96175 1 25064
2 96176 1 25064
2 96177 1 25064
2 96178 1 25064
2 96179 1 25066
2 96180 1 25066
2 96181 1 25066
2 96182 1 25066
2 96183 1 25066
2 96184 1 25066
2 96185 1 25067
2 96186 1 25067
2 96187 1 25067
2 96188 1 25075
2 96189 1 25075
2 96190 1 25078
2 96191 1 25078
2 96192 1 25079
2 96193 1 25079
2 96194 1 25079
2 96195 1 25079
2 96196 1 25090
2 96197 1 25090
2 96198 1 25093
2 96199 1 25093
2 96200 1 25093
2 96201 1 25093
2 96202 1 25093
2 96203 1 25093
2 96204 1 25093
2 96205 1 25093
2 96206 1 25096
2 96207 1 25096
2 96208 1 25107
2 96209 1 25107
2 96210 1 25107
2 96211 1 25107
2 96212 1 25115
2 96213 1 25115
2 96214 1 25124
2 96215 1 25124
2 96216 1 25124
2 96217 1 25125
2 96218 1 25125
2 96219 1 25125
2 96220 1 25140
2 96221 1 25140
2 96222 1 25143
2 96223 1 25143
2 96224 1 25145
2 96225 1 25145
2 96226 1 25170
2 96227 1 25170
2 96228 1 25170
2 96229 1 25171
2 96230 1 25171
2 96231 1 25176
2 96232 1 25176
2 96233 1 25179
2 96234 1 25179
2 96235 1 25181
2 96236 1 25181
2 96237 1 25181
2 96238 1 25181
2 96239 1 25181
2 96240 1 25181
2 96241 1 25181
2 96242 1 25192
2 96243 1 25192
2 96244 1 25207
2 96245 1 25207
2 96246 1 25207
2 96247 1 25207
2 96248 1 25207
2 96249 1 25207
2 96250 1 25220
2 96251 1 25220
2 96252 1 25232
2 96253 1 25232
2 96254 1 25245
2 96255 1 25245
2 96256 1 25245
2 96257 1 25245
2 96258 1 25246
2 96259 1 25246
2 96260 1 25247
2 96261 1 25247
2 96262 1 25256
2 96263 1 25256
2 96264 1 25268
2 96265 1 25268
2 96266 1 25268
2 96267 1 25268
2 96268 1 25291
2 96269 1 25291
2 96270 1 25295
2 96271 1 25295
2 96272 1 25296
2 96273 1 25296
2 96274 1 25296
2 96275 1 25298
2 96276 1 25298
2 96277 1 25298
2 96278 1 25298
2 96279 1 25301
2 96280 1 25301
2 96281 1 25311
2 96282 1 25311
2 96283 1 25311
2 96284 1 25311
2 96285 1 25324
2 96286 1 25324
2 96287 1 25325
2 96288 1 25325
2 96289 1 25325
2 96290 1 25325
2 96291 1 25334
2 96292 1 25334
2 96293 1 25334
2 96294 1 25372
2 96295 1 25372
2 96296 1 25372
2 96297 1 25373
2 96298 1 25373
2 96299 1 25378
2 96300 1 25378
2 96301 1 25378
2 96302 1 25381
2 96303 1 25381
2 96304 1 25381
2 96305 1 25381
2 96306 1 25389
2 96307 1 25389
2 96308 1 25392
2 96309 1 25392
2 96310 1 25392
2 96311 1 25400
2 96312 1 25400
2 96313 1 25406
2 96314 1 25406
2 96315 1 25409
2 96316 1 25409
2 96317 1 25478
2 96318 1 25478
2 96319 1 25488
2 96320 1 25488
2 96321 1 25555
2 96322 1 25555
2 96323 1 25555
2 96324 1 25555
2 96325 1 25576
2 96326 1 25576
2 96327 1 25622
2 96328 1 25622
2 96329 1 25624
2 96330 1 25624
2 96331 1 25652
2 96332 1 25652
2 96333 1 25652
2 96334 1 25667
2 96335 1 25667
2 96336 1 25667
2 96337 1 25668
2 96338 1 25668
2 96339 1 25669
2 96340 1 25669
2 96341 1 25687
2 96342 1 25687
2 96343 1 25687
2 96344 1 25687
2 96345 1 25687
2 96346 1 25709
2 96347 1 25709
2 96348 1 25710
2 96349 1 25710
2 96350 1 25726
2 96351 1 25726
2 96352 1 25726
2 96353 1 25730
2 96354 1 25730
2 96355 1 25764
2 96356 1 25764
2 96357 1 25786
2 96358 1 25786
2 96359 1 25786
2 96360 1 25786
2 96361 1 25786
2 96362 1 25786
2 96363 1 25787
2 96364 1 25787
2 96365 1 25788
2 96366 1 25788
2 96367 1 25800
2 96368 1 25800
2 96369 1 25813
2 96370 1 25813
2 96371 1 25814
2 96372 1 25814
2 96373 1 25815
2 96374 1 25815
2 96375 1 25838
2 96376 1 25838
2 96377 1 25866
2 96378 1 25866
2 96379 1 25867
2 96380 1 25867
2 96381 1 25867
2 96382 1 25872
2 96383 1 25872
2 96384 1 25907
2 96385 1 25907
2 96386 1 25907
2 96387 1 25907
2 96388 1 25911
2 96389 1 25911
2 96390 1 25911
2 96391 1 25911
2 96392 1 25911
2 96393 1 25911
2 96394 1 25911
2 96395 1 25911
2 96396 1 25918
2 96397 1 25918
2 96398 1 25933
2 96399 1 25933
2 96400 1 25937
2 96401 1 25937
2 96402 1 25938
2 96403 1 25938
2 96404 1 25948
2 96405 1 25948
2 96406 1 25949
2 96407 1 25949
2 96408 1 25949
2 96409 1 25972
2 96410 1 25972
2 96411 1 25976
2 96412 1 25976
2 96413 1 25976
2 96414 1 25976
2 96415 1 25976
2 96416 1 25976
2 96417 1 25977
2 96418 1 25977
2 96419 1 25977
2 96420 1 25977
2 96421 1 25995
2 96422 1 25995
2 96423 1 25998
2 96424 1 25998
2 96425 1 26005
2 96426 1 26005
2 96427 1 26011
2 96428 1 26011
2 96429 1 26012
2 96430 1 26012
2 96431 1 26012
2 96432 1 26015
2 96433 1 26015
2 96434 1 26015
2 96435 1 26015
2 96436 1 26015
2 96437 1 26015
2 96438 1 26018
2 96439 1 26018
2 96440 1 26034
2 96441 1 26034
2 96442 1 26038
2 96443 1 26038
2 96444 1 26039
2 96445 1 26039
2 96446 1 26039
2 96447 1 26039
2 96448 1 26039
2 96449 1 26039
2 96450 1 26039
2 96451 1 26039
2 96452 1 26039
2 96453 1 26039
2 96454 1 26039
2 96455 1 26065
2 96456 1 26065
2 96457 1 26065
2 96458 1 26066
2 96459 1 26066
2 96460 1 26066
2 96461 1 26079
2 96462 1 26079
2 96463 1 26079
2 96464 1 26106
2 96465 1 26106
2 96466 1 26114
2 96467 1 26114
2 96468 1 26119
2 96469 1 26119
2 96470 1 26119
2 96471 1 26124
2 96472 1 26124
2 96473 1 26145
2 96474 1 26145
2 96475 1 26145
2 96476 1 26145
2 96477 1 26145
2 96478 1 26146
2 96479 1 26146
2 96480 1 26181
2 96481 1 26181
2 96482 1 26187
2 96483 1 26187
2 96484 1 26187
2 96485 1 26187
2 96486 1 26187
2 96487 1 26195
2 96488 1 26195
2 96489 1 26207
2 96490 1 26207
2 96491 1 26207
2 96492 1 26207
2 96493 1 26208
2 96494 1 26208
2 96495 1 26209
2 96496 1 26209
2 96497 1 26209
2 96498 1 26209
2 96499 1 26209
2 96500 1 26209
2 96501 1 26209
2 96502 1 26212
2 96503 1 26212
2 96504 1 26212
2 96505 1 26212
2 96506 1 26215
2 96507 1 26215
2 96508 1 26215
2 96509 1 26215
2 96510 1 26216
2 96511 1 26216
2 96512 1 26217
2 96513 1 26217
2 96514 1 26217
2 96515 1 26221
2 96516 1 26221
2 96517 1 26221
2 96518 1 26221
2 96519 1 26221
2 96520 1 26221
2 96521 1 26221
2 96522 1 26230
2 96523 1 26230
2 96524 1 26230
2 96525 1 26230
2 96526 1 26230
2 96527 1 26230
2 96528 1 26231
2 96529 1 26231
2 96530 1 26231
2 96531 1 26231
2 96532 1 26231
2 96533 1 26244
2 96534 1 26244
2 96535 1 26262
2 96536 1 26262
2 96537 1 26263
2 96538 1 26263
2 96539 1 26263
2 96540 1 26263
2 96541 1 26263
2 96542 1 26263
2 96543 1 26277
2 96544 1 26277
2 96545 1 26284
2 96546 1 26284
2 96547 1 26284
2 96548 1 26284
2 96549 1 26284
2 96550 1 26284
2 96551 1 26284
2 96552 1 26289
2 96553 1 26289
2 96554 1 26289
2 96555 1 26309
2 96556 1 26309
2 96557 1 26309
2 96558 1 26309
2 96559 1 26328
2 96560 1 26328
2 96561 1 26331
2 96562 1 26331
2 96563 1 26332
2 96564 1 26332
2 96565 1 26334
2 96566 1 26334
2 96567 1 26334
2 96568 1 26334
2 96569 1 26342
2 96570 1 26342
2 96571 1 26358
2 96572 1 26358
2 96573 1 26371
2 96574 1 26371
2 96575 1 26372
2 96576 1 26372
2 96577 1 26383
2 96578 1 26383
2 96579 1 26383
2 96580 1 26384
2 96581 1 26384
2 96582 1 26385
2 96583 1 26385
2 96584 1 26407
2 96585 1 26407
2 96586 1 26407
2 96587 1 26407
2 96588 1 26407
2 96589 1 26407
2 96590 1 26407
2 96591 1 26407
2 96592 1 26407
2 96593 1 26407
2 96594 1 26408
2 96595 1 26408
2 96596 1 26409
2 96597 1 26409
2 96598 1 26412
2 96599 1 26412
2 96600 1 26431
2 96601 1 26431
2 96602 1 26440
2 96603 1 26440
2 96604 1 26448
2 96605 1 26448
2 96606 1 26448
2 96607 1 26469
2 96608 1 26469
2 96609 1 26501
2 96610 1 26501
2 96611 1 26512
2 96612 1 26512
2 96613 1 26533
2 96614 1 26533
2 96615 1 26541
2 96616 1 26541
2 96617 1 26541
2 96618 1 26541
2 96619 1 26541
2 96620 1 26541
2 96621 1 26541
2 96622 1 26541
2 96623 1 26550
2 96624 1 26550
2 96625 1 26551
2 96626 1 26551
2 96627 1 26564
2 96628 1 26564
2 96629 1 26564
2 96630 1 26564
2 96631 1 26580
2 96632 1 26580
2 96633 1 26585
2 96634 1 26585
2 96635 1 26593
2 96636 1 26593
2 96637 1 26596
2 96638 1 26596
2 96639 1 26597
2 96640 1 26597
2 96641 1 26600
2 96642 1 26600
2 96643 1 26659
2 96644 1 26659
2 96645 1 26659
2 96646 1 26666
2 96647 1 26666
2 96648 1 26666
2 96649 1 26666
2 96650 1 26666
2 96651 1 26666
2 96652 1 26669
2 96653 1 26669
2 96654 1 26691
2 96655 1 26691
2 96656 1 26691
2 96657 1 26692
2 96658 1 26692
2 96659 1 26701
2 96660 1 26701
2 96661 1 26708
2 96662 1 26708
2 96663 1 26708
2 96664 1 26709
2 96665 1 26709
2 96666 1 26710
2 96667 1 26710
2 96668 1 26711
2 96669 1 26711
2 96670 1 26711
2 96671 1 26724
2 96672 1 26724
2 96673 1 26724
2 96674 1 26724
2 96675 1 26737
2 96676 1 26737
2 96677 1 26740
2 96678 1 26740
2 96679 1 26740
2 96680 1 26740
2 96681 1 26740
2 96682 1 26740
2 96683 1 26740
2 96684 1 26740
2 96685 1 26752
2 96686 1 26752
2 96687 1 26752
2 96688 1 26752
2 96689 1 26753
2 96690 1 26753
2 96691 1 26754
2 96692 1 26754
2 96693 1 26761
2 96694 1 26761
2 96695 1 26761
2 96696 1 26761
2 96697 1 26783
2 96698 1 26783
2 96699 1 26783
2 96700 1 26796
2 96701 1 26796
2 96702 1 26796
2 96703 1 26808
2 96704 1 26808
2 96705 1 26815
2 96706 1 26815
2 96707 1 26816
2 96708 1 26816
2 96709 1 26818
2 96710 1 26818
2 96711 1 26818
2 96712 1 26818
2 96713 1 26820
2 96714 1 26820
2 96715 1 26835
2 96716 1 26835
2 96717 1 26848
2 96718 1 26848
2 96719 1 26852
2 96720 1 26852
2 96721 1 26857
2 96722 1 26857
2 96723 1 26857
2 96724 1 26857
2 96725 1 26858
2 96726 1 26858
2 96727 1 26858
2 96728 1 26875
2 96729 1 26875
2 96730 1 26875
2 96731 1 26875
2 96732 1 26876
2 96733 1 26876
2 96734 1 26903
2 96735 1 26903
2 96736 1 26909
2 96737 1 26909
2 96738 1 26909
2 96739 1 26909
2 96740 1 26909
2 96741 1 26909
2 96742 1 26909
2 96743 1 26909
2 96744 1 26909
2 96745 1 26920
2 96746 1 26920
2 96747 1 26970
2 96748 1 26970
2 96749 1 27011
2 96750 1 27011
2 96751 1 27028
2 96752 1 27028
2 96753 1 27047
2 96754 1 27047
2 96755 1 27047
2 96756 1 27047
2 96757 1 27051
2 96758 1 27051
2 96759 1 27059
2 96760 1 27059
2 96761 1 27069
2 96762 1 27069
2 96763 1 27081
2 96764 1 27081
2 96765 1 27081
2 96766 1 27081
2 96767 1 27090
2 96768 1 27090
2 96769 1 27101
2 96770 1 27101
2 96771 1 27101
2 96772 1 27101
2 96773 1 27101
2 96774 1 27102
2 96775 1 27102
2 96776 1 27102
2 96777 1 27102
2 96778 1 27103
2 96779 1 27103
2 96780 1 27104
2 96781 1 27104
2 96782 1 27104
2 96783 1 27112
2 96784 1 27112
2 96785 1 27116
2 96786 1 27116
2 96787 1 27116
2 96788 1 27128
2 96789 1 27128
2 96790 1 27145
2 96791 1 27145
2 96792 1 27150
2 96793 1 27150
2 96794 1 27150
2 96795 1 27150
2 96796 1 27150
2 96797 1 27164
2 96798 1 27164
2 96799 1 27199
2 96800 1 27199
2 96801 1 27207
2 96802 1 27207
2 96803 1 27207
2 96804 1 27207
2 96805 1 27217
2 96806 1 27217
2 96807 1 27226
2 96808 1 27226
2 96809 1 27233
2 96810 1 27233
2 96811 1 27251
2 96812 1 27251
2 96813 1 27277
2 96814 1 27277
2 96815 1 27285
2 96816 1 27285
2 96817 1 27285
2 96818 1 27294
2 96819 1 27294
2 96820 1 27311
2 96821 1 27311
2 96822 1 27311
2 96823 1 27312
2 96824 1 27312
2 96825 1 27342
2 96826 1 27342
2 96827 1 27342
2 96828 1 27342
2 96829 1 27394
2 96830 1 27394
2 96831 1 27394
2 96832 1 27394
2 96833 1 27394
2 96834 1 27394
2 96835 1 27394
2 96836 1 27395
2 96837 1 27395
2 96838 1 27395
2 96839 1 27398
2 96840 1 27398
2 96841 1 27415
2 96842 1 27415
2 96843 1 27415
2 96844 1 27415
2 96845 1 27423
2 96846 1 27423
2 96847 1 27454
2 96848 1 27454
2 96849 1 27454
2 96850 1 27455
2 96851 1 27455
2 96852 1 27468
2 96853 1 27468
2 96854 1 27468
2 96855 1 27475
2 96856 1 27475
2 96857 1 27475
2 96858 1 27475
2 96859 1 27475
2 96860 1 27484
2 96861 1 27484
2 96862 1 27484
2 96863 1 27486
2 96864 1 27486
2 96865 1 27486
2 96866 1 27500
2 96867 1 27500
2 96868 1 27581
2 96869 1 27581
2 96870 1 27591
2 96871 1 27591
2 96872 1 27591
2 96873 1 27591
2 96874 1 27619
2 96875 1 27619
2 96876 1 27634
2 96877 1 27634
2 96878 1 27634
2 96879 1 27634
2 96880 1 27646
2 96881 1 27646
2 96882 1 27646
2 96883 1 27646
2 96884 1 27655
2 96885 1 27655
2 96886 1 27662
2 96887 1 27662
2 96888 1 27682
2 96889 1 27682
2 96890 1 27682
2 96891 1 27682
2 96892 1 27682
2 96893 1 27682
2 96894 1 27682
2 96895 1 27684
2 96896 1 27684
2 96897 1 27684
2 96898 1 27693
2 96899 1 27693
2 96900 1 27693
2 96901 1 27693
2 96902 1 27693
2 96903 1 27693
2 96904 1 27694
2 96905 1 27694
2 96906 1 27697
2 96907 1 27697
2 96908 1 27697
2 96909 1 27698
2 96910 1 27698
2 96911 1 27698
2 96912 1 27698
2 96913 1 27723
2 96914 1 27723
2 96915 1 27724
2 96916 1 27724
2 96917 1 27736
2 96918 1 27736
2 96919 1 27736
2 96920 1 27736
2 96921 1 27736
2 96922 1 27768
2 96923 1 27768
2 96924 1 27768
2 96925 1 27780
2 96926 1 27780
2 96927 1 27781
2 96928 1 27781
2 96929 1 27781
2 96930 1 27781
2 96931 1 27781
2 96932 1 27782
2 96933 1 27782
2 96934 1 27783
2 96935 1 27783
2 96936 1 27783
2 96937 1 27801
2 96938 1 27801
2 96939 1 27801
2 96940 1 27801
2 96941 1 27801
2 96942 1 27801
2 96943 1 27801
2 96944 1 27801
2 96945 1 27801
2 96946 1 27801
2 96947 1 27801
2 96948 1 27801
2 96949 1 27801
2 96950 1 27801
2 96951 1 27801
2 96952 1 27801
2 96953 1 27802
2 96954 1 27802
2 96955 1 27802
2 96956 1 27803
2 96957 1 27803
2 96958 1 27803
2 96959 1 27803
2 96960 1 27803
2 96961 1 27803
2 96962 1 27803
2 96963 1 27803
2 96964 1 27803
2 96965 1 27803
2 96966 1 27803
2 96967 1 27803
2 96968 1 27803
2 96969 1 27803
2 96970 1 27803
2 96971 1 27803
2 96972 1 27803
2 96973 1 27803
2 96974 1 27803
2 96975 1 27803
2 96976 1 27803
2 96977 1 27803
2 96978 1 27803
2 96979 1 27803
2 96980 1 27803
2 96981 1 27803
2 96982 1 27803
2 96983 1 27821
2 96984 1 27821
2 96985 1 27831
2 96986 1 27831
2 96987 1 27861
2 96988 1 27861
2 96989 1 27861
2 96990 1 27862
2 96991 1 27862
2 96992 1 27911
2 96993 1 27911
2 96994 1 27921
2 96995 1 27921
2 96996 1 27931
2 96997 1 27931
2 96998 1 27931
2 96999 1 27931
2 97000 1 27931
2 97001 1 27931
2 97002 1 27931
2 97003 1 27948
2 97004 1 27948
2 97005 1 27949
2 97006 1 27949
2 97007 1 27949
2 97008 1 27960
2 97009 1 27960
2 97010 1 27973
2 97011 1 27973
2 97012 1 27973
2 97013 1 27973
2 97014 1 27973
2 97015 1 27973
2 97016 1 27973
2 97017 1 27973
2 97018 1 27973
2 97019 1 27973
2 97020 1 27974
2 97021 1 27974
2 97022 1 27974
2 97023 1 27974
2 97024 1 27976
2 97025 1 27976
2 97026 1 28002
2 97027 1 28002
2 97028 1 28003
2 97029 1 28003
2 97030 1 28003
2 97031 1 28003
2 97032 1 28003
2 97033 1 28007
2 97034 1 28007
2 97035 1 28017
2 97036 1 28017
2 97037 1 28017
2 97038 1 28017
2 97039 1 28017
2 97040 1 28017
2 97041 1 28031
2 97042 1 28031
2 97043 1 28032
2 97044 1 28032
2 97045 1 28032
2 97046 1 28037
2 97047 1 28037
2 97048 1 28040
2 97049 1 28040
2 97050 1 28064
2 97051 1 28064
2 97052 1 28085
2 97053 1 28085
2 97054 1 28086
2 97055 1 28086
2 97056 1 28087
2 97057 1 28087
2 97058 1 28087
2 97059 1 28087
2 97060 1 28088
2 97061 1 28088
2 97062 1 28093
2 97063 1 28093
2 97064 1 28101
2 97065 1 28101
2 97066 1 28134
2 97067 1 28134
2 97068 1 28135
2 97069 1 28135
2 97070 1 28136
2 97071 1 28136
2 97072 1 28150
2 97073 1 28150
2 97074 1 28192
2 97075 1 28192
2 97076 1 28197
2 97077 1 28197
2 97078 1 28197
2 97079 1 28197
2 97080 1 28197
2 97081 1 28240
2 97082 1 28240
2 97083 1 28240
2 97084 1 28240
2 97085 1 28250
2 97086 1 28250
2 97087 1 28278
2 97088 1 28278
2 97089 1 28280
2 97090 1 28280
2 97091 1 28289
2 97092 1 28289
2 97093 1 28289
2 97094 1 28289
2 97095 1 28289
2 97096 1 28289
2 97097 1 28298
2 97098 1 28298
2 97099 1 28298
2 97100 1 28301
2 97101 1 28301
2 97102 1 28301
2 97103 1 28332
2 97104 1 28332
2 97105 1 28332
2 97106 1 28332
2 97107 1 28336
2 97108 1 28336
2 97109 1 28337
2 97110 1 28337
2 97111 1 28337
2 97112 1 28337
2 97113 1 28337
2 97114 1 28346
2 97115 1 28346
2 97116 1 28366
2 97117 1 28366
2 97118 1 28366
2 97119 1 28367
2 97120 1 28367
2 97121 1 28367
2 97122 1 28368
2 97123 1 28368
2 97124 1 28368
2 97125 1 28416
2 97126 1 28416
2 97127 1 28433
2 97128 1 28433
2 97129 1 28453
2 97130 1 28453
2 97131 1 28455
2 97132 1 28455
2 97133 1 28464
2 97134 1 28464
2 97135 1 28464
2 97136 1 28464
2 97137 1 28481
2 97138 1 28481
2 97139 1 28481
2 97140 1 28481
2 97141 1 28490
2 97142 1 28490
2 97143 1 28499
2 97144 1 28499
2 97145 1 28512
2 97146 1 28512
2 97147 1 28512
2 97148 1 28512
2 97149 1 28513
2 97150 1 28513
2 97151 1 28514
2 97152 1 28514
2 97153 1 28517
2 97154 1 28517
2 97155 1 28538
2 97156 1 28538
2 97157 1 28538
2 97158 1 28538
2 97159 1 28549
2 97160 1 28549
2 97161 1 28549
2 97162 1 28549
2 97163 1 28557
2 97164 1 28557
2 97165 1 28557
2 97166 1 28558
2 97167 1 28558
2 97168 1 28560
2 97169 1 28560
2 97170 1 28560
2 97171 1 28560
2 97172 1 28560
2 97173 1 28560
2 97174 1 28569
2 97175 1 28569
2 97176 1 28618
2 97177 1 28618
2 97178 1 28619
2 97179 1 28619
2 97180 1 28627
2 97181 1 28627
2 97182 1 28655
2 97183 1 28655
2 97184 1 28656
2 97185 1 28656
2 97186 1 28660
2 97187 1 28660
2 97188 1 28668
2 97189 1 28668
2 97190 1 28669
2 97191 1 28669
2 97192 1 28678
2 97193 1 28678
2 97194 1 28678
2 97195 1 28678
2 97196 1 28680
2 97197 1 28680
2 97198 1 28689
2 97199 1 28689
2 97200 1 28691
2 97201 1 28691
2 97202 1 28691
2 97203 1 28695
2 97204 1 28695
2 97205 1 28705
2 97206 1 28705
2 97207 1 28705
2 97208 1 28706
2 97209 1 28706
2 97210 1 28706
2 97211 1 28731
2 97212 1 28731
2 97213 1 28740
2 97214 1 28740
2 97215 1 28762
2 97216 1 28762
2 97217 1 28773
2 97218 1 28773
2 97219 1 28822
2 97220 1 28822
2 97221 1 28822
2 97222 1 28833
2 97223 1 28833
2 97224 1 28833
2 97225 1 28836
2 97226 1 28836
2 97227 1 28836
2 97228 1 28844
2 97229 1 28844
2 97230 1 28844
2 97231 1 28885
2 97232 1 28885
2 97233 1 28885
2 97234 1 28888
2 97235 1 28888
2 97236 1 28908
2 97237 1 28908
2 97238 1 28908
2 97239 1 28937
2 97240 1 28937
2 97241 1 28937
2 97242 1 28937
2 97243 1 28937
2 97244 1 28941
2 97245 1 28941
2 97246 1 28966
2 97247 1 28966
2 97248 1 28989
2 97249 1 28989
2 97250 1 28994
2 97251 1 28994
2 97252 1 29050
2 97253 1 29050
2 97254 1 29100
2 97255 1 29100
2 97256 1 29100
2 97257 1 29105
2 97258 1 29105
2 97259 1 29160
2 97260 1 29160
2 97261 1 29160
2 97262 1 29164
2 97263 1 29164
2 97264 1 29165
2 97265 1 29165
2 97266 1 29168
2 97267 1 29168
2 97268 1 29176
2 97269 1 29176
2 97270 1 29176
2 97271 1 29193
2 97272 1 29193
2 97273 1 29194
2 97274 1 29194
2 97275 1 29205
2 97276 1 29205
2 97277 1 29205
2 97278 1 29213
2 97279 1 29213
2 97280 1 29240
2 97281 1 29240
2 97282 1 29240
2 97283 1 29241
2 97284 1 29241
2 97285 1 29241
2 97286 1 29261
2 97287 1 29261
2 97288 1 29261
2 97289 1 29261
2 97290 1 29261
2 97291 1 29261
2 97292 1 29267
2 97293 1 29267
2 97294 1 29267
2 97295 1 29275
2 97296 1 29275
2 97297 1 29279
2 97298 1 29279
2 97299 1 29305
2 97300 1 29305
2 97301 1 29320
2 97302 1 29320
2 97303 1 29340
2 97304 1 29340
2 97305 1 29340
2 97306 1 29340
2 97307 1 29340
2 97308 1 29340
2 97309 1 29340
2 97310 1 29340
2 97311 1 29340
2 97312 1 29340
2 97313 1 29340
2 97314 1 29340
2 97315 1 29340
2 97316 1 29340
2 97317 1 29340
2 97318 1 29340
2 97319 1 29340
2 97320 1 29340
2 97321 1 29340
2 97322 1 29340
2 97323 1 29340
2 97324 1 29340
2 97325 1 29340
2 97326 1 29340
2 97327 1 29340
2 97328 1 29348
2 97329 1 29348
2 97330 1 29348
2 97331 1 29351
2 97332 1 29351
2 97333 1 29358
2 97334 1 29358
2 97335 1 29358
2 97336 1 29359
2 97337 1 29359
2 97338 1 29359
2 97339 1 29359
2 97340 1 29359
2 97341 1 29359
2 97342 1 29375
2 97343 1 29375
2 97344 1 29397
2 97345 1 29397
2 97346 1 29397
2 97347 1 29397
2 97348 1 29397
2 97349 1 29398
2 97350 1 29398
2 97351 1 29398
2 97352 1 29398
2 97353 1 29398
2 97354 1 29408
2 97355 1 29408
2 97356 1 29408
2 97357 1 29408
2 97358 1 29408
2 97359 1 29408
2 97360 1 29409
2 97361 1 29409
2 97362 1 29409
2 97363 1 29419
2 97364 1 29419
2 97365 1 29420
2 97366 1 29420
2 97367 1 29420
2 97368 1 29420
2 97369 1 29420
2 97370 1 29420
2 97371 1 29420
2 97372 1 29438
2 97373 1 29438
2 97374 1 29450
2 97375 1 29450
2 97376 1 29469
2 97377 1 29469
2 97378 1 29469
2 97379 1 29469
2 97380 1 29469
2 97381 1 29469
2 97382 1 29469
2 97383 1 29470
2 97384 1 29470
2 97385 1 29470
2 97386 1 29472
2 97387 1 29472
2 97388 1 29472
2 97389 1 29483
2 97390 1 29483
2 97391 1 29483
2 97392 1 29484
2 97393 1 29484
2 97394 1 29489
2 97395 1 29489
2 97396 1 29490
2 97397 1 29490
2 97398 1 29490
2 97399 1 29491
2 97400 1 29491
2 97401 1 29491
2 97402 1 29496
2 97403 1 29496
2 97404 1 29499
2 97405 1 29499
2 97406 1 29500
2 97407 1 29500
2 97408 1 29500
2 97409 1 29500
2 97410 1 29517
2 97411 1 29517
2 97412 1 29518
2 97413 1 29518
2 97414 1 29520
2 97415 1 29520
2 97416 1 29520
2 97417 1 29520
2 97418 1 29520
2 97419 1 29520
2 97420 1 29520
2 97421 1 29520
2 97422 1 29520
2 97423 1 29520
2 97424 1 29520
2 97425 1 29520
2 97426 1 29520
2 97427 1 29521
2 97428 1 29521
2 97429 1 29529
2 97430 1 29529
2 97431 1 29529
2 97432 1 29542
2 97433 1 29542
2 97434 1 29542
2 97435 1 29542
2 97436 1 29542
2 97437 1 29542
2 97438 1 29543
2 97439 1 29543
2 97440 1 29545
2 97441 1 29545
2 97442 1 29550
2 97443 1 29550
2 97444 1 29550
2 97445 1 29550
2 97446 1 29550
2 97447 1 29550
2 97448 1 29556
2 97449 1 29556
2 97450 1 29556
2 97451 1 29556
2 97452 1 29564
2 97453 1 29564
2 97454 1 29564
2 97455 1 29565
2 97456 1 29565
2 97457 1 29565
2 97458 1 29565
2 97459 1 29565
2 97460 1 29565
2 97461 1 29565
2 97462 1 29565
2 97463 1 29565
2 97464 1 29566
2 97465 1 29566
2 97466 1 29566
2 97467 1 29566
2 97468 1 29566
2 97469 1 29567
2 97470 1 29567
2 97471 1 29570
2 97472 1 29570
2 97473 1 29573
2 97474 1 29573
2 97475 1 29574
2 97476 1 29574
2 97477 1 29589
2 97478 1 29589
2 97479 1 29589
2 97480 1 29589
2 97481 1 29606
2 97482 1 29606
2 97483 1 29607
2 97484 1 29607
2 97485 1 29625
2 97486 1 29625
2 97487 1 29625
2 97488 1 29636
2 97489 1 29636
2 97490 1 29636
2 97491 1 29636
2 97492 1 29636
2 97493 1 29638
2 97494 1 29638
2 97495 1 29649
2 97496 1 29649
2 97497 1 29662
2 97498 1 29662
2 97499 1 29664
2 97500 1 29664
2 97501 1 29664
2 97502 1 29664
2 97503 1 29664
2 97504 1 29664
2 97505 1 29664
2 97506 1 29664
2 97507 1 29665
2 97508 1 29665
2 97509 1 29668
2 97510 1 29668
2 97511 1 29684
2 97512 1 29684
2 97513 1 29688
2 97514 1 29688
2 97515 1 29688
2 97516 1 29688
2 97517 1 29693
2 97518 1 29693
2 97519 1 29693
2 97520 1 29693
2 97521 1 29696
2 97522 1 29696
2 97523 1 29697
2 97524 1 29697
2 97525 1 29697
2 97526 1 29697
2 97527 1 29697
2 97528 1 29697
2 97529 1 29697
2 97530 1 29703
2 97531 1 29703
2 97532 1 29704
2 97533 1 29704
2 97534 1 29707
2 97535 1 29707
2 97536 1 29749
2 97537 1 29749
2 97538 1 29750
2 97539 1 29750
2 97540 1 29750
2 97541 1 29750
2 97542 1 29751
2 97543 1 29751
2 97544 1 29751
2 97545 1 29751
2 97546 1 29752
2 97547 1 29752
2 97548 1 29752
2 97549 1 29755
2 97550 1 29755
2 97551 1 29755
2 97552 1 29755
2 97553 1 29756
2 97554 1 29756
2 97555 1 29764
2 97556 1 29764
2 97557 1 29765
2 97558 1 29765
2 97559 1 29765
2 97560 1 29773
2 97561 1 29773
2 97562 1 29778
2 97563 1 29778
2 97564 1 29778
2 97565 1 29778
2 97566 1 29778
2 97567 1 29778
2 97568 1 29778
2 97569 1 29778
2 97570 1 29779
2 97571 1 29779
2 97572 1 29779
2 97573 1 29779
2 97574 1 29779
2 97575 1 29779
2 97576 1 29779
2 97577 1 29779
2 97578 1 29784
2 97579 1 29784
2 97580 1 29785
2 97581 1 29785
2 97582 1 29785
2 97583 1 29785
2 97584 1 29785
2 97585 1 29785
2 97586 1 29785
2 97587 1 29785
2 97588 1 29785
2 97589 1 29785
2 97590 1 29785
2 97591 1 29785
2 97592 1 29785
2 97593 1 29785
2 97594 1 29785
2 97595 1 29786
2 97596 1 29786
2 97597 1 29787
2 97598 1 29787
2 97599 1 29787
2 97600 1 29791
2 97601 1 29791
2 97602 1 29791
2 97603 1 29791
2 97604 1 29791
2 97605 1 29791
2 97606 1 29791
2 97607 1 29799
2 97608 1 29799
2 97609 1 29799
2 97610 1 29799
2 97611 1 29799
2 97612 1 29799
2 97613 1 29799
2 97614 1 29799
2 97615 1 29799
2 97616 1 29799
2 97617 1 29799
2 97618 1 29799
2 97619 1 29799
2 97620 1 29799
2 97621 1 29799
2 97622 1 29799
2 97623 1 29799
2 97624 1 29810
2 97625 1 29810
2 97626 1 29810
2 97627 1 29810
2 97628 1 29810
2 97629 1 29810
2 97630 1 29810
2 97631 1 29810
2 97632 1 29810
2 97633 1 29810
2 97634 1 29810
2 97635 1 29810
2 97636 1 29810
2 97637 1 29810
2 97638 1 29810
2 97639 1 29810
2 97640 1 29811
2 97641 1 29811
2 97642 1 29826
2 97643 1 29826
2 97644 1 29826
2 97645 1 29826
2 97646 1 29826
2 97647 1 29826
2 97648 1 29826
2 97649 1 29826
2 97650 1 29826
2 97651 1 29826
2 97652 1 29826
2 97653 1 29826
2 97654 1 29826
2 97655 1 29826
2 97656 1 29827
2 97657 1 29827
2 97658 1 29827
2 97659 1 29827
2 97660 1 29827
2 97661 1 29827
2 97662 1 29827
2 97663 1 29827
2 97664 1 29827
2 97665 1 29827
2 97666 1 29827
2 97667 1 29827
2 97668 1 29827
2 97669 1 29827
2 97670 1 29827
2 97671 1 29827
2 97672 1 29827
2 97673 1 29827
2 97674 1 29827
2 97675 1 29827
2 97676 1 29827
2 97677 1 29827
2 97678 1 29827
2 97679 1 29827
2 97680 1 29827
2 97681 1 29827
2 97682 1 29827
2 97683 1 29827
2 97684 1 29827
2 97685 1 29827
2 97686 1 29827
2 97687 1 29827
2 97688 1 29827
2 97689 1 29828
2 97690 1 29828
2 97691 1 29829
2 97692 1 29829
2 97693 1 29829
2 97694 1 29838
2 97695 1 29838
2 97696 1 29839
2 97697 1 29839
2 97698 1 29839
2 97699 1 29845
2 97700 1 29845
2 97701 1 29848
2 97702 1 29848
2 97703 1 29862
2 97704 1 29862
2 97705 1 29870
2 97706 1 29870
2 97707 1 29870
2 97708 1 29870
2 97709 1 29870
2 97710 1 29870
2 97711 1 29870
2 97712 1 29870
2 97713 1 29870
2 97714 1 29870
2 97715 1 29870
2 97716 1 29870
2 97717 1 29870
2 97718 1 29870
2 97719 1 29870
2 97720 1 29870
2 97721 1 29870
2 97722 1 29870
2 97723 1 29870
2 97724 1 29870
2 97725 1 29870
2 97726 1 29870
2 97727 1 29870
2 97728 1 29870
2 97729 1 29870
2 97730 1 29870
2 97731 1 29870
2 97732 1 29870
2 97733 1 29870
2 97734 1 29871
2 97735 1 29871
2 97736 1 29871
2 97737 1 29871
2 97738 1 29871
2 97739 1 29871
2 97740 1 29871
2 97741 1 29871
2 97742 1 29871
2 97743 1 29871
2 97744 1 29871
2 97745 1 29871
2 97746 1 29871
2 97747 1 29871
2 97748 1 29871
2 97749 1 29871
2 97750 1 29871
2 97751 1 29871
2 97752 1 29871
2 97753 1 29871
2 97754 1 29871
2 97755 1 29871
2 97756 1 29872
2 97757 1 29872
2 97758 1 29888
2 97759 1 29888
2 97760 1 29893
2 97761 1 29893
2 97762 1 29893
2 97763 1 29904
2 97764 1 29904
2 97765 1 29913
2 97766 1 29913
2 97767 1 29916
2 97768 1 29916
2 97769 1 29934
2 97770 1 29934
2 97771 1 29947
2 97772 1 29947
2 97773 1 29947
2 97774 1 29947
2 97775 1 29947
2 97776 1 29947
2 97777 1 29947
2 97778 1 29947
2 97779 1 29948
2 97780 1 29948
2 97781 1 29948
2 97782 1 29948
2 97783 1 29950
2 97784 1 29950
2 97785 1 29956
2 97786 1 29956
2 97787 1 29956
2 97788 1 29956
2 97789 1 29956
2 97790 1 29956
2 97791 1 29956
2 97792 1 29956
2 97793 1 29956
2 97794 1 29956
2 97795 1 29956
2 97796 1 29956
2 97797 1 29956
2 97798 1 29966
2 97799 1 29966
2 97800 1 29968
2 97801 1 29968
2 97802 1 29972
2 97803 1 29972
2 97804 1 29972
2 97805 1 29972
2 97806 1 29972
2 97807 1 29972
2 97808 1 29975
2 97809 1 29975
2 97810 1 29982
2 97811 1 29982
2 97812 1 29982
2 97813 1 29983
2 97814 1 29983
2 97815 1 29990
2 97816 1 29990
2 97817 1 29990
2 97818 1 29990
2 97819 1 29990
2 97820 1 29991
2 97821 1 29991
2 97822 1 29992
2 97823 1 29992
2 97824 1 29992
2 97825 1 29992
2 97826 1 29993
2 97827 1 29993
2 97828 1 29998
2 97829 1 29998
2 97830 1 30015
2 97831 1 30015
2 97832 1 30033
2 97833 1 30033
2 97834 1 30035
2 97835 1 30035
2 97836 1 30042
2 97837 1 30042
2 97838 1 30042
2 97839 1 30078
2 97840 1 30078
2 97841 1 30100
2 97842 1 30100
2 97843 1 30107
2 97844 1 30107
2 97845 1 30107
2 97846 1 30118
2 97847 1 30118
2 97848 1 30118
2 97849 1 30118
2 97850 1 30120
2 97851 1 30120
2 97852 1 30124
2 97853 1 30124
2 97854 1 30124
2 97855 1 30139
2 97856 1 30139
2 97857 1 30139
2 97858 1 30163
2 97859 1 30163
2 97860 1 30163
2 97861 1 30164
2 97862 1 30164
2 97863 1 30165
2 97864 1 30165
2 97865 1 30191
2 97866 1 30191
2 97867 1 30191
2 97868 1 30191
2 97869 1 30191
2 97870 1 30191
2 97871 1 30222
2 97872 1 30222
2 97873 1 30230
2 97874 1 30230
2 97875 1 30230
2 97876 1 30230
2 97877 1 30252
2 97878 1 30252
2 97879 1 30265
2 97880 1 30265
2 97881 1 30265
2 97882 1 30265
2 97883 1 30265
2 97884 1 30265
2 97885 1 30266
2 97886 1 30266
2 97887 1 30267
2 97888 1 30267
2 97889 1 30270
2 97890 1 30270
2 97891 1 30280
2 97892 1 30280
2 97893 1 30281
2 97894 1 30281
2 97895 1 30289
2 97896 1 30289
2 97897 1 30305
2 97898 1 30305
2 97899 1 30332
2 97900 1 30332
2 97901 1 30337
2 97902 1 30337
2 97903 1 30339
2 97904 1 30339
2 97905 1 30339
2 97906 1 30339
2 97907 1 30348
2 97908 1 30348
2 97909 1 30360
2 97910 1 30360
2 97911 1 30361
2 97912 1 30361
2 97913 1 30366
2 97914 1 30366
2 97915 1 30376
2 97916 1 30376
2 97917 1 30376
2 97918 1 30376
2 97919 1 30376
2 97920 1 30383
2 97921 1 30383
2 97922 1 30386
2 97923 1 30386
2 97924 1 30388
2 97925 1 30388
2 97926 1 30389
2 97927 1 30389
2 97928 1 30408
2 97929 1 30408
2 97930 1 30419
2 97931 1 30419
2 97932 1 30427
2 97933 1 30427
2 97934 1 30434
2 97935 1 30434
2 97936 1 30482
2 97937 1 30482
2 97938 1 30485
2 97939 1 30485
2 97940 1 30507
2 97941 1 30507
2 97942 1 30507
2 97943 1 30508
2 97944 1 30508
2 97945 1 30508
2 97946 1 30510
2 97947 1 30510
2 97948 1 30510
2 97949 1 30517
2 97950 1 30517
2 97951 1 30520
2 97952 1 30520
2 97953 1 30526
2 97954 1 30526
2 97955 1 30537
2 97956 1 30537
2 97957 1 30538
2 97958 1 30538
2 97959 1 30546
2 97960 1 30546
2 97961 1 30570
2 97962 1 30570
2 97963 1 30570
2 97964 1 30571
2 97965 1 30571
2 97966 1 30600
2 97967 1 30600
2 97968 1 30634
2 97969 1 30634
2 97970 1 30654
2 97971 1 30654
2 97972 1 30664
2 97973 1 30664
2 97974 1 30664
2 97975 1 30672
2 97976 1 30672
2 97977 1 30677
2 97978 1 30677
2 97979 1 30688
2 97980 1 30688
2 97981 1 30688
2 97982 1 30688
2 97983 1 30688
2 97984 1 30688
2 97985 1 30688
2 97986 1 30688
2 97987 1 30688
2 97988 1 30688
2 97989 1 30688
2 97990 1 30688
2 97991 1 30688
2 97992 1 30688
2 97993 1 30688
2 97994 1 30688
2 97995 1 30688
2 97996 1 30688
2 97997 1 30688
2 97998 1 30688
2 97999 1 30688
2 98000 1 30688
2 98001 1 30688
2 98002 1 30689
2 98003 1 30689
2 98004 1 30689
2 98005 1 30689
2 98006 1 30689
2 98007 1 30689
2 98008 1 30689
2 98009 1 30689
2 98010 1 30689
2 98011 1 30689
2 98012 1 30689
2 98013 1 30689
2 98014 1 30689
2 98015 1 30689
2 98016 1 30689
2 98017 1 30689
2 98018 1 30689
2 98019 1 30689
2 98020 1 30689
2 98021 1 30689
2 98022 1 30689
2 98023 1 30689
2 98024 1 30689
2 98025 1 30689
2 98026 1 30689
2 98027 1 30689
2 98028 1 30689
2 98029 1 30689
2 98030 1 30689
2 98031 1 30696
2 98032 1 30696
2 98033 1 30723
2 98034 1 30723
2 98035 1 30723
2 98036 1 30723
2 98037 1 30723
2 98038 1 30723
2 98039 1 30723
2 98040 1 30723
2 98041 1 30723
2 98042 1 30723
2 98043 1 30723
2 98044 1 30723
2 98045 1 30723
2 98046 1 30724
2 98047 1 30724
2 98048 1 30724
2 98049 1 30724
2 98050 1 30724
2 98051 1 30724
2 98052 1 30724
2 98053 1 30725
2 98054 1 30725
2 98055 1 30725
2 98056 1 30726
2 98057 1 30726
2 98058 1 30731
2 98059 1 30731
2 98060 1 30742
2 98061 1 30742
2 98062 1 30760
2 98063 1 30760
2 98064 1 30760
2 98065 1 30760
2 98066 1 30770
2 98067 1 30770
2 98068 1 30777
2 98069 1 30777
2 98070 1 30777
2 98071 1 30777
2 98072 1 30778
2 98073 1 30778
2 98074 1 30778
2 98075 1 30778
2 98076 1 30778
2 98077 1 30779
2 98078 1 30779
2 98079 1 30779
2 98080 1 30779
2 98081 1 30779
2 98082 1 30779
2 98083 1 30787
2 98084 1 30787
2 98085 1 30787
2 98086 1 30787
2 98087 1 30787
2 98088 1 30787
2 98089 1 30787
2 98090 1 30787
2 98091 1 30787
2 98092 1 30787
2 98093 1 30787
2 98094 1 30790
2 98095 1 30790
2 98096 1 30856
2 98097 1 30856
2 98098 1 30866
2 98099 1 30866
2 98100 1 30866
2 98101 1 30866
2 98102 1 30866
2 98103 1 30866
2 98104 1 30866
2 98105 1 30866
2 98106 1 30866
2 98107 1 30866
2 98108 1 30866
2 98109 1 30866
2 98110 1 30866
2 98111 1 30866
2 98112 1 30866
2 98113 1 30866
2 98114 1 30867
2 98115 1 30867
2 98116 1 30867
2 98117 1 30867
2 98118 1 30868
2 98119 1 30868
2 98120 1 30876
2 98121 1 30876
2 98122 1 30876
2 98123 1 30876
2 98124 1 30876
2 98125 1 30877
2 98126 1 30877
2 98127 1 30877
2 98128 1 30878
2 98129 1 30878
2 98130 1 30888
2 98131 1 30888
2 98132 1 30889
2 98133 1 30889
2 98134 1 30889
2 98135 1 30897
2 98136 1 30897
2 98137 1 30897
2 98138 1 30898
2 98139 1 30898
2 98140 1 30898
2 98141 1 30898
2 98142 1 30898
2 98143 1 30898
2 98144 1 30900
2 98145 1 30900
2 98146 1 30901
2 98147 1 30901
2 98148 1 30902
2 98149 1 30902
2 98150 1 30924
2 98151 1 30924
2 98152 1 30924
2 98153 1 30924
2 98154 1 30924
2 98155 1 30924
2 98156 1 30924
2 98157 1 30925
2 98158 1 30925
2 98159 1 30929
2 98160 1 30929
2 98161 1 30929
2 98162 1 30929
2 98163 1 30929
2 98164 1 30944
2 98165 1 30944
2 98166 1 30944
2 98167 1 30944
2 98168 1 30944
2 98169 1 30945
2 98170 1 30945
2 98171 1 30945
2 98172 1 30946
2 98173 1 30946
2 98174 1 30946
2 98175 1 30949
2 98176 1 30949
2 98177 1 30950
2 98178 1 30950
2 98179 1 30950
2 98180 1 30950
2 98181 1 30950
2 98182 1 30950
2 98183 1 30950
2 98184 1 30950
2 98185 1 30951
2 98186 1 30951
2 98187 1 30951
2 98188 1 30952
2 98189 1 30952
2 98190 1 30952
2 98191 1 30952
2 98192 1 30960
2 98193 1 30960
2 98194 1 30960
2 98195 1 30960
2 98196 1 30960
2 98197 1 30960
2 98198 1 30961
2 98199 1 30961
2 98200 1 30961
2 98201 1 30961
2 98202 1 30972
2 98203 1 30972
2 98204 1 30972
2 98205 1 30984
2 98206 1 30984
2 98207 1 30984
2 98208 1 30984
2 98209 1 30984
2 98210 1 30984
2 98211 1 30984
2 98212 1 30985
2 98213 1 30985
2 98214 1 30985
2 98215 1 30985
2 98216 1 31007
2 98217 1 31007
2 98218 1 31007
2 98219 1 31007
2 98220 1 31008
2 98221 1 31008
2 98222 1 31009
2 98223 1 31009
2 98224 1 31009
2 98225 1 31025
2 98226 1 31025
2 98227 1 31033
2 98228 1 31033
2 98229 1 31044
2 98230 1 31044
2 98231 1 31048
2 98232 1 31048
2 98233 1 31059
2 98234 1 31059
2 98235 1 31087
2 98236 1 31087
2 98237 1 31088
2 98238 1 31088
2 98239 1 31103
2 98240 1 31103
2 98241 1 31115
2 98242 1 31115
2 98243 1 31142
2 98244 1 31142
2 98245 1 31142
2 98246 1 31142
2 98247 1 31142
2 98248 1 31167
2 98249 1 31167
2 98250 1 31167
2 98251 1 31181
2 98252 1 31181
2 98253 1 31181
2 98254 1 31196
2 98255 1 31196
2 98256 1 31196
2 98257 1 31196
2 98258 1 31197
2 98259 1 31197
2 98260 1 31205
2 98261 1 31205
2 98262 1 31206
2 98263 1 31206
2 98264 1 31213
2 98265 1 31213
2 98266 1 31253
2 98267 1 31253
2 98268 1 31261
2 98269 1 31261
2 98270 1 31295
2 98271 1 31295
2 98272 1 31304
2 98273 1 31304
2 98274 1 31304
2 98275 1 31304
2 98276 1 31330
2 98277 1 31330
2 98278 1 31345
2 98279 1 31345
2 98280 1 31345
2 98281 1 31361
2 98282 1 31361
2 98283 1 31375
2 98284 1 31375
2 98285 1 31375
2 98286 1 31424
2 98287 1 31424
2 98288 1 31476
2 98289 1 31476
2 98290 1 31476
2 98291 1 31476
2 98292 1 31477
2 98293 1 31477
2 98294 1 31477
2 98295 1 31477
2 98296 1 31477
2 98297 1 31477
2 98298 1 31477
2 98299 1 31477
2 98300 1 31477
2 98301 1 31477
2 98302 1 31477
2 98303 1 31477
2 98304 1 31477
2 98305 1 31477
2 98306 1 31477
2 98307 1 31477
2 98308 1 31477
2 98309 1 31477
2 98310 1 31477
2 98311 1 31477
2 98312 1 31477
2 98313 1 31477
2 98314 1 31477
2 98315 1 31477
2 98316 1 31477
2 98317 1 31477
2 98318 1 31477
2 98319 1 31477
2 98320 1 31477
2 98321 1 31477
2 98322 1 31477
2 98323 1 31477
2 98324 1 31477
2 98325 1 31477
2 98326 1 31477
2 98327 1 31477
2 98328 1 31477
2 98329 1 31477
2 98330 1 31477
2 98331 1 31477
2 98332 1 31477
2 98333 1 31490
2 98334 1 31490
2 98335 1 31503
2 98336 1 31503
2 98337 1 31504
2 98338 1 31504
2 98339 1 31504
2 98340 1 31504
2 98341 1 31504
2 98342 1 31504
2 98343 1 31505
2 98344 1 31505
2 98345 1 31508
2 98346 1 31508
2 98347 1 31508
2 98348 1 31511
2 98349 1 31511
2 98350 1 31512
2 98351 1 31512
2 98352 1 31522
2 98353 1 31522
2 98354 1 31524
2 98355 1 31524
2 98356 1 31525
2 98357 1 31525
2 98358 1 31525
2 98359 1 31525
2 98360 1 31537
2 98361 1 31537
2 98362 1 31537
2 98363 1 31537
2 98364 1 31538
2 98365 1 31538
2 98366 1 31539
2 98367 1 31539
2 98368 1 31539
2 98369 1 31539
2 98370 1 31540
2 98371 1 31540
2 98372 1 31548
2 98373 1 31548
2 98374 1 31548
2 98375 1 31566
2 98376 1 31566
2 98377 1 31568
2 98378 1 31568
2 98379 1 31592
2 98380 1 31592
2 98381 1 31592
2 98382 1 31592
2 98383 1 31592
2 98384 1 31592
2 98385 1 31592
2 98386 1 31593
2 98387 1 31593
2 98388 1 31595
2 98389 1 31595
2 98390 1 31595
2 98391 1 31598
2 98392 1 31598
2 98393 1 31598
2 98394 1 31598
2 98395 1 31598
2 98396 1 31598
2 98397 1 31598
2 98398 1 31598
2 98399 1 31598
2 98400 1 31601
2 98401 1 31601
2 98402 1 31601
2 98403 1 31601
2 98404 1 31601
2 98405 1 31601
2 98406 1 31601
2 98407 1 31602
2 98408 1 31602
2 98409 1 31602
2 98410 1 31602
2 98411 1 31603
2 98412 1 31603
2 98413 1 31606
2 98414 1 31606
2 98415 1 31606
2 98416 1 31606
2 98417 1 31606
2 98418 1 31606
2 98419 1 31606
2 98420 1 31607
2 98421 1 31607
2 98422 1 31607
2 98423 1 31607
2 98424 1 31607
2 98425 1 31607
2 98426 1 31608
2 98427 1 31608
2 98428 1 31611
2 98429 1 31611
2 98430 1 31616
2 98431 1 31616
2 98432 1 31619
2 98433 1 31619
2 98434 1 31620
2 98435 1 31620
2 98436 1 31620
2 98437 1 31620
2 98438 1 31620
2 98439 1 31620
2 98440 1 31620
2 98441 1 31628
2 98442 1 31628
2 98443 1 31629
2 98444 1 31629
2 98445 1 31629
2 98446 1 31632
2 98447 1 31632
2 98448 1 31640
2 98449 1 31640
2 98450 1 31640
2 98451 1 31640
2 98452 1 31640
2 98453 1 31641
2 98454 1 31641
2 98455 1 31641
2 98456 1 31641
2 98457 1 31648
2 98458 1 31648
2 98459 1 31663
2 98460 1 31663
2 98461 1 31663
2 98462 1 31663
2 98463 1 31663
2 98464 1 31664
2 98465 1 31664
2 98466 1 31675
2 98467 1 31675
2 98468 1 31676
2 98469 1 31676
2 98470 1 31676
2 98471 1 31676
2 98472 1 31676
2 98473 1 31676
2 98474 1 31676
2 98475 1 31676
2 98476 1 31676
2 98477 1 31676
2 98478 1 31676
2 98479 1 31676
2 98480 1 31685
2 98481 1 31685
2 98482 1 31685
2 98483 1 31689
2 98484 1 31689
2 98485 1 31698
2 98486 1 31698
2 98487 1 31699
2 98488 1 31699
2 98489 1 31699
2 98490 1 31700
2 98491 1 31700
2 98492 1 31700
2 98493 1 31716
2 98494 1 31716
2 98495 1 31716
2 98496 1 31716
2 98497 1 31716
2 98498 1 31716
2 98499 1 31719
2 98500 1 31719
2 98501 1 31728
2 98502 1 31728
2 98503 1 31728
2 98504 1 31728
2 98505 1 31735
2 98506 1 31735
2 98507 1 31735
2 98508 1 31735
2 98509 1 31741
2 98510 1 31741
2 98511 1 31741
2 98512 1 31741
2 98513 1 31741
2 98514 1 31744
2 98515 1 31744
2 98516 1 31752
2 98517 1 31752
2 98518 1 31766
2 98519 1 31766
2 98520 1 31766
2 98521 1 31766
2 98522 1 31766
2 98523 1 31766
2 98524 1 31766
2 98525 1 31766
2 98526 1 31766
2 98527 1 31766
2 98528 1 31766
2 98529 1 31766
2 98530 1 31766
2 98531 1 31766
2 98532 1 31766
2 98533 1 31767
2 98534 1 31767
2 98535 1 31774
2 98536 1 31774
2 98537 1 31774
2 98538 1 31774
2 98539 1 31774
2 98540 1 31774
2 98541 1 31774
2 98542 1 31785
2 98543 1 31785
2 98544 1 31790
2 98545 1 31790
2 98546 1 31790
2 98547 1 31790
2 98548 1 31790
2 98549 1 31790
2 98550 1 31792
2 98551 1 31792
2 98552 1 31797
2 98553 1 31797
2 98554 1 31799
2 98555 1 31799
2 98556 1 31799
2 98557 1 31799
2 98558 1 31800
2 98559 1 31800
2 98560 1 31800
2 98561 1 31803
2 98562 1 31803
2 98563 1 31803
2 98564 1 31803
2 98565 1 31803
2 98566 1 31804
2 98567 1 31804
2 98568 1 31804
2 98569 1 31808
2 98570 1 31808
2 98571 1 31808
2 98572 1 31809
2 98573 1 31809
2 98574 1 31809
2 98575 1 31809
2 98576 1 31809
2 98577 1 31809
2 98578 1 31809
2 98579 1 31818
2 98580 1 31818
2 98581 1 31819
2 98582 1 31819
2 98583 1 31819
2 98584 1 31819
2 98585 1 31819
2 98586 1 31819
2 98587 1 31820
2 98588 1 31820
2 98589 1 31824
2 98590 1 31824
2 98591 1 31824
2 98592 1 31824
2 98593 1 31825
2 98594 1 31825
2 98595 1 31825
2 98596 1 31825
2 98597 1 31826
2 98598 1 31826
2 98599 1 31834
2 98600 1 31834
2 98601 1 31834
2 98602 1 31834
2 98603 1 31834
2 98604 1 31852
2 98605 1 31852
2 98606 1 31855
2 98607 1 31855
2 98608 1 31857
2 98609 1 31857
2 98610 1 31858
2 98611 1 31858
2 98612 1 31858
2 98613 1 31858
2 98614 1 31861
2 98615 1 31861
2 98616 1 31861
2 98617 1 31870
2 98618 1 31870
2 98619 1 31870
2 98620 1 31870
2 98621 1 31870
2 98622 1 31870
2 98623 1 31870
2 98624 1 31870
2 98625 1 31870
2 98626 1 31870
2 98627 1 31874
2 98628 1 31874
2 98629 1 31874
2 98630 1 31874
2 98631 1 31874
2 98632 1 31888
2 98633 1 31888
2 98634 1 31891
2 98635 1 31891
2 98636 1 31891
2 98637 1 31891
2 98638 1 31899
2 98639 1 31899
2 98640 1 31902
2 98641 1 31902
2 98642 1 31902
2 98643 1 31913
2 98644 1 31913
2 98645 1 31913
2 98646 1 31913
2 98647 1 31913
2 98648 1 31913
2 98649 1 31913
2 98650 1 31913
2 98651 1 31917
2 98652 1 31917
2 98653 1 31917
2 98654 1 31917
2 98655 1 31917
2 98656 1 31917
2 98657 1 31917
2 98658 1 31917
2 98659 1 31917
2 98660 1 31917
2 98661 1 31917
2 98662 1 31918
2 98663 1 31918
2 98664 1 31919
2 98665 1 31919
2 98666 1 31923
2 98667 1 31923
2 98668 1 31923
2 98669 1 31923
2 98670 1 31923
2 98671 1 31923
2 98672 1 31923
2 98673 1 31923
2 98674 1 31923
2 98675 1 31923
2 98676 1 31923
2 98677 1 31934
2 98678 1 31934
2 98679 1 31934
2 98680 1 31934
2 98681 1 31934
2 98682 1 31934
2 98683 1 31934
2 98684 1 31934
2 98685 1 31934
2 98686 1 31934
2 98687 1 31934
2 98688 1 31934
2 98689 1 31936
2 98690 1 31936
2 98691 1 31957
2 98692 1 31957
2 98693 1 31970
2 98694 1 31970
2 98695 1 31970
2 98696 1 31970
2 98697 1 31971
2 98698 1 31971
2 98699 1 31971
2 98700 1 31971
2 98701 1 31971
2 98702 1 31980
2 98703 1 31980
2 98704 1 31988
2 98705 1 31988
2 98706 1 31988
2 98707 1 31999
2 98708 1 31999
2 98709 1 31999
2 98710 1 31999
2 98711 1 32003
2 98712 1 32003
2 98713 1 32003
2 98714 1 32003
2 98715 1 32004
2 98716 1 32004
2 98717 1 32004
2 98718 1 32005
2 98719 1 32005
2 98720 1 32013
2 98721 1 32013
2 98722 1 32015
2 98723 1 32015
2 98724 1 32015
2 98725 1 32015
2 98726 1 32015
2 98727 1 32023
2 98728 1 32023
2 98729 1 32024
2 98730 1 32024
2 98731 1 32024
2 98732 1 32024
2 98733 1 32024
2 98734 1 32024
2 98735 1 32034
2 98736 1 32034
2 98737 1 32034
2 98738 1 32034
2 98739 1 32034
2 98740 1 32035
2 98741 1 32035
2 98742 1 32035
2 98743 1 32036
2 98744 1 32036
2 98745 1 32037
2 98746 1 32037
2 98747 1 32037
2 98748 1 32037
2 98749 1 32037
2 98750 1 32042
2 98751 1 32042
2 98752 1 32057
2 98753 1 32057
2 98754 1 32057
2 98755 1 32059
2 98756 1 32059
2 98757 1 32062
2 98758 1 32062
2 98759 1 32062
2 98760 1 32075
2 98761 1 32075
2 98762 1 32075
2 98763 1 32076
2 98764 1 32076
2 98765 1 32089
2 98766 1 32089
2 98767 1 32106
2 98768 1 32106
2 98769 1 32106
2 98770 1 32106
2 98771 1 32106
2 98772 1 32106
2 98773 1 32107
2 98774 1 32107
2 98775 1 32121
2 98776 1 32121
2 98777 1 32124
2 98778 1 32124
2 98779 1 32124
2 98780 1 32126
2 98781 1 32126
2 98782 1 32131
2 98783 1 32131
2 98784 1 32147
2 98785 1 32147
2 98786 1 32153
2 98787 1 32153
2 98788 1 32170
2 98789 1 32170
2 98790 1 32173
2 98791 1 32173
2 98792 1 32178
2 98793 1 32178
2 98794 1 32194
2 98795 1 32194
2 98796 1 32196
2 98797 1 32196
2 98798 1 32196
2 98799 1 32196
2 98800 1 32196
2 98801 1 32197
2 98802 1 32197
2 98803 1 32198
2 98804 1 32198
2 98805 1 32199
2 98806 1 32199
2 98807 1 32200
2 98808 1 32200
2 98809 1 32200
2 98810 1 32200
2 98811 1 32200
2 98812 1 32200
2 98813 1 32203
2 98814 1 32203
2 98815 1 32206
2 98816 1 32206
2 98817 1 32211
2 98818 1 32211
2 98819 1 32218
2 98820 1 32218
2 98821 1 32219
2 98822 1 32219
2 98823 1 32221
2 98824 1 32221
2 98825 1 32222
2 98826 1 32222
2 98827 1 32223
2 98828 1 32223
2 98829 1 32223
2 98830 1 32223
2 98831 1 32232
2 98832 1 32232
2 98833 1 32232
2 98834 1 32244
2 98835 1 32244
2 98836 1 32244
2 98837 1 32245
2 98838 1 32245
2 98839 1 32253
2 98840 1 32253
2 98841 1 32282
2 98842 1 32282
2 98843 1 32282
2 98844 1 32282
2 98845 1 32291
2 98846 1 32291
2 98847 1 32291
2 98848 1 32293
2 98849 1 32293
2 98850 1 32293
2 98851 1 32303
2 98852 1 32303
2 98853 1 32304
2 98854 1 32304
2 98855 1 32314
2 98856 1 32314
2 98857 1 32314
2 98858 1 32348
2 98859 1 32348
2 98860 1 32366
2 98861 1 32366
2 98862 1 32374
2 98863 1 32374
2 98864 1 32377
2 98865 1 32377
2 98866 1 32380
2 98867 1 32380
2 98868 1 32380
2 98869 1 32380
2 98870 1 32398
2 98871 1 32398
2 98872 1 32403
2 98873 1 32403
2 98874 1 32403
2 98875 1 32403
2 98876 1 32403
2 98877 1 32404
2 98878 1 32404
2 98879 1 32416
2 98880 1 32416
2 98881 1 32416
2 98882 1 32416
2 98883 1 32416
2 98884 1 32416
2 98885 1 32416
2 98886 1 32416
2 98887 1 32416
2 98888 1 32416
2 98889 1 32416
2 98890 1 32416
2 98891 1 32416
2 98892 1 32416
2 98893 1 32416
2 98894 1 32416
2 98895 1 32416
2 98896 1 32416
2 98897 1 32416
2 98898 1 32416
2 98899 1 32416
2 98900 1 32430
2 98901 1 32430
2 98902 1 32438
2 98903 1 32438
2 98904 1 32438
2 98905 1 32460
2 98906 1 32460
2 98907 1 32461
2 98908 1 32461
2 98909 1 32464
2 98910 1 32464
2 98911 1 32464
2 98912 1 32464
2 98913 1 32465
2 98914 1 32465
2 98915 1 32473
2 98916 1 32473
2 98917 1 32473
2 98918 1 32473
2 98919 1 32473
2 98920 1 32474
2 98921 1 32474
2 98922 1 32493
2 98923 1 32493
2 98924 1 32536
2 98925 1 32536
2 98926 1 32537
2 98927 1 32537
2 98928 1 32546
2 98929 1 32546
2 98930 1 32546
2 98931 1 32558
2 98932 1 32558
2 98933 1 32567
2 98934 1 32567
2 98935 1 32578
2 98936 1 32578
2 98937 1 32578
2 98938 1 32578
2 98939 1 32578
2 98940 1 32578
2 98941 1 32587
2 98942 1 32587
2 98943 1 32626
2 98944 1 32626
2 98945 1 32646
2 98946 1 32646
2 98947 1 32647
2 98948 1 32647
2 98949 1 32700
2 98950 1 32700
2 98951 1 32700
2 98952 1 32703
2 98953 1 32703
2 98954 1 32706
2 98955 1 32706
2 98956 1 32706
2 98957 1 32706
2 98958 1 32706
2 98959 1 32725
2 98960 1 32725
2 98961 1 32725
2 98962 1 32728
2 98963 1 32728
2 98964 1 32728
2 98965 1 32728
2 98966 1 32733
2 98967 1 32733
2 98968 1 32741
2 98969 1 32741
2 98970 1 32743
2 98971 1 32743
2 98972 1 32761
2 98973 1 32761
2 98974 1 32761
2 98975 1 32761
2 98976 1 32761
2 98977 1 32788
2 98978 1 32788
2 98979 1 32788
2 98980 1 32788
2 98981 1 32788
2 98982 1 32788
2 98983 1 32788
2 98984 1 32788
2 98985 1 32789
2 98986 1 32789
2 98987 1 32789
2 98988 1 32789
2 98989 1 32800
2 98990 1 32800
2 98991 1 32801
2 98992 1 32801
2 98993 1 32832
2 98994 1 32832
2 98995 1 32832
2 98996 1 32832
2 98997 1 32832
2 98998 1 32832
2 98999 1 32833
2 99000 1 32833
2 99001 1 32834
2 99002 1 32834
2 99003 1 32848
2 99004 1 32848
2 99005 1 32849
2 99006 1 32849
2 99007 1 32849
2 99008 1 32849
2 99009 1 32857
2 99010 1 32857
2 99011 1 32857
2 99012 1 32858
2 99013 1 32858
2 99014 1 32859
2 99015 1 32859
2 99016 1 32859
2 99017 1 32859
2 99018 1 32859
2 99019 1 32859
2 99020 1 32859
2 99021 1 32859
2 99022 1 32859
2 99023 1 32859
2 99024 1 32859
2 99025 1 32859
2 99026 1 32859
2 99027 1 32859
2 99028 1 32859
2 99029 1 32859
2 99030 1 32859
2 99031 1 32861
2 99032 1 32861
2 99033 1 32861
2 99034 1 32869
2 99035 1 32869
2 99036 1 32869
2 99037 1 32869
2 99038 1 32869
2 99039 1 32869
2 99040 1 32869
2 99041 1 32869
2 99042 1 32878
2 99043 1 32878
2 99044 1 32878
2 99045 1 32878
2 99046 1 32878
2 99047 1 32878
2 99048 1 32878
2 99049 1 32878
2 99050 1 32878
2 99051 1 32878
2 99052 1 32878
2 99053 1 32878
2 99054 1 32878
2 99055 1 32878
2 99056 1 32878
2 99057 1 32878
2 99058 1 32878
2 99059 1 32879
2 99060 1 32879
2 99061 1 32886
2 99062 1 32886
2 99063 1 32886
2 99064 1 32917
2 99065 1 32917
2 99066 1 32917
2 99067 1 32918
2 99068 1 32918
2 99069 1 32918
2 99070 1 32919
2 99071 1 32919
2 99072 1 32919
2 99073 1 32919
2 99074 1 32919
2 99075 1 32930
2 99076 1 32930
2 99077 1 32930
2 99078 1 32931
2 99079 1 32931
2 99080 1 32939
2 99081 1 32939
2 99082 1 32948
2 99083 1 32948
2 99084 1 32949
2 99085 1 32949
2 99086 1 32958
2 99087 1 32958
2 99088 1 32958
2 99089 1 32958
2 99090 1 32958
2 99091 1 32958
2 99092 1 32958
2 99093 1 32959
2 99094 1 32959
2 99095 1 32965
2 99096 1 32965
2 99097 1 32965
2 99098 1 32965
2 99099 1 32965
2 99100 1 32965
2 99101 1 32965
2 99102 1 32965
2 99103 1 32973
2 99104 1 32973
2 99105 1 32973
2 99106 1 32973
2 99107 1 32973
2 99108 1 32973
2 99109 1 32973
2 99110 1 32973
2 99111 1 32973
2 99112 1 32979
2 99113 1 32979
2 99114 1 32979
2 99115 1 32979
2 99116 1 32979
2 99117 1 32980
2 99118 1 32980
2 99119 1 32980
2 99120 1 32980
2 99121 1 32980
2 99122 1 32980
2 99123 1 32980
2 99124 1 32980
2 99125 1 32980
2 99126 1 32980
2 99127 1 32990
2 99128 1 32990
2 99129 1 32990
2 99130 1 32994
2 99131 1 32994
2 99132 1 32994
2 99133 1 32994
2 99134 1 32994
2 99135 1 32998
2 99136 1 32998
2 99137 1 33000
2 99138 1 33000
2 99139 1 33000
2 99140 1 33006
2 99141 1 33006
2 99142 1 33015
2 99143 1 33015
2 99144 1 33026
2 99145 1 33026
2 99146 1 33026
2 99147 1 33027
2 99148 1 33027
2 99149 1 33027
2 99150 1 33027
2 99151 1 33027
2 99152 1 33027
2 99153 1 33027
2 99154 1 33027
2 99155 1 33027
2 99156 1 33027
2 99157 1 33042
2 99158 1 33042
2 99159 1 33042
2 99160 1 33043
2 99161 1 33043
2 99162 1 33043
2 99163 1 33047
2 99164 1 33047
2 99165 1 33047
2 99166 1 33047
2 99167 1 33047
2 99168 1 33047
2 99169 1 33047
2 99170 1 33047
2 99171 1 33047
2 99172 1 33047
2 99173 1 33048
2 99174 1 33048
2 99175 1 33068
2 99176 1 33068
2 99177 1 33068
2 99178 1 33069
2 99179 1 33069
2 99180 1 33078
2 99181 1 33078
2 99182 1 33078
2 99183 1 33082
2 99184 1 33082
2 99185 1 33092
2 99186 1 33092
2 99187 1 33092
2 99188 1 33101
2 99189 1 33101
2 99190 1 33101
2 99191 1 33101
2 99192 1 33102
2 99193 1 33102
2 99194 1 33102
2 99195 1 33102
2 99196 1 33102
2 99197 1 33104
2 99198 1 33104
2 99199 1 33105
2 99200 1 33105
2 99201 1 33115
2 99202 1 33115
2 99203 1 33115
2 99204 1 33115
2 99205 1 33115
2 99206 1 33115
2 99207 1 33115
2 99208 1 33115
2 99209 1 33116
2 99210 1 33116
2 99211 1 33116
2 99212 1 33116
2 99213 1 33117
2 99214 1 33117
2 99215 1 33118
2 99216 1 33118
2 99217 1 33120
2 99218 1 33120
2 99219 1 33132
2 99220 1 33132
2 99221 1 33132
2 99222 1 33132
2 99223 1 33133
2 99224 1 33133
2 99225 1 33133
2 99226 1 33133
2 99227 1 33133
2 99228 1 33134
2 99229 1 33134
2 99230 1 33134
2 99231 1 33143
2 99232 1 33143
2 99233 1 33146
2 99234 1 33146
2 99235 1 33160
2 99236 1 33160
2 99237 1 33183
2 99238 1 33183
2 99239 1 33183
2 99240 1 33200
2 99241 1 33200
2 99242 1 33201
2 99243 1 33201
2 99244 1 33204
2 99245 1 33204
2 99246 1 33204
2 99247 1 33205
2 99248 1 33205
2 99249 1 33208
2 99250 1 33208
2 99251 1 33208
2 99252 1 33208
2 99253 1 33211
2 99254 1 33211
2 99255 1 33211
2 99256 1 33211
2 99257 1 33211
2 99258 1 33211
2 99259 1 33212
2 99260 1 33212
2 99261 1 33212
2 99262 1 33213
2 99263 1 33213
2 99264 1 33213
2 99265 1 33222
2 99266 1 33222
2 99267 1 33242
2 99268 1 33242
2 99269 1 33251
2 99270 1 33251
2 99271 1 33252
2 99272 1 33252
2 99273 1 33269
2 99274 1 33269
2 99275 1 33269
2 99276 1 33269
2 99277 1 33269
2 99278 1 33269
2 99279 1 33277
2 99280 1 33277
2 99281 1 33286
2 99282 1 33286
2 99283 1 33286
2 99284 1 33295
2 99285 1 33295
2 99286 1 33296
2 99287 1 33296
2 99288 1 33296
2 99289 1 33296
2 99290 1 33308
2 99291 1 33308
2 99292 1 33325
2 99293 1 33325
2 99294 1 33325
2 99295 1 33327
2 99296 1 33327
2 99297 1 33327
2 99298 1 33327
2 99299 1 33341
2 99300 1 33341
2 99301 1 33341
2 99302 1 33341
2 99303 1 33341
2 99304 1 33342
2 99305 1 33342
2 99306 1 33342
2 99307 1 33342
2 99308 1 33342
2 99309 1 33345
2 99310 1 33345
2 99311 1 33345
2 99312 1 33346
2 99313 1 33346
2 99314 1 33346
2 99315 1 33353
2 99316 1 33353
2 99317 1 33353
2 99318 1 33353
2 99319 1 33353
2 99320 1 33354
2 99321 1 33354
2 99322 1 33374
2 99323 1 33374
2 99324 1 33378
2 99325 1 33378
2 99326 1 33378
2 99327 1 33378
2 99328 1 33378
2 99329 1 33378
2 99330 1 33378
2 99331 1 33379
2 99332 1 33379
2 99333 1 33379
2 99334 1 33379
2 99335 1 33396
2 99336 1 33396
2 99337 1 33396
2 99338 1 33404
2 99339 1 33404
2 99340 1 33407
2 99341 1 33407
2 99342 1 33407
2 99343 1 33407
2 99344 1 33407
2 99345 1 33416
2 99346 1 33416
2 99347 1 33439
2 99348 1 33439
2 99349 1 33442
2 99350 1 33442
2 99351 1 33443
2 99352 1 33443
2 99353 1 33443
2 99354 1 33444
2 99355 1 33444
2 99356 1 33458
2 99357 1 33458
2 99358 1 33461
2 99359 1 33461
2 99360 1 33475
2 99361 1 33475
2 99362 1 33475
2 99363 1 33477
2 99364 1 33477
2 99365 1 33477
2 99366 1 33477
2 99367 1 33477
2 99368 1 33477
2 99369 1 33477
2 99370 1 33477
2 99371 1 33477
2 99372 1 33477
2 99373 1 33477
2 99374 1 33478
2 99375 1 33478
2 99376 1 33478
2 99377 1 33478
2 99378 1 33478
2 99379 1 33478
2 99380 1 33484
2 99381 1 33484
2 99382 1 33484
2 99383 1 33484
2 99384 1 33484
2 99385 1 33484
2 99386 1 33484
2 99387 1 33484
2 99388 1 33484
2 99389 1 33484
2 99390 1 33484
2 99391 1 33498
2 99392 1 33498
2 99393 1 33498
2 99394 1 33499
2 99395 1 33499
2 99396 1 33509
2 99397 1 33509
2 99398 1 33509
2 99399 1 33547
2 99400 1 33547
2 99401 1 33561
2 99402 1 33561
2 99403 1 33568
2 99404 1 33568
2 99405 1 33589
2 99406 1 33589
2 99407 1 33589
2 99408 1 33590
2 99409 1 33590
2 99410 1 33590
2 99411 1 33590
2 99412 1 33590
2 99413 1 33611
2 99414 1 33611
2 99415 1 33611
2 99416 1 33612
2 99417 1 33612
2 99418 1 33612
2 99419 1 33612
2 99420 1 33612
2 99421 1 33612
2 99422 1 33612
2 99423 1 33622
2 99424 1 33622
2 99425 1 33622
2 99426 1 33632
2 99427 1 33632
2 99428 1 33632
2 99429 1 33641
2 99430 1 33641
2 99431 1 33650
2 99432 1 33650
2 99433 1 33653
2 99434 1 33653
2 99435 1 33670
2 99436 1 33670
2 99437 1 33670
2 99438 1 33675
2 99439 1 33675
2 99440 1 33675
2 99441 1 33675
2 99442 1 33677
2 99443 1 33677
2 99444 1 33686
2 99445 1 33686
2 99446 1 33686
2 99447 1 33696
2 99448 1 33696
2 99449 1 33696
2 99450 1 33697
2 99451 1 33697
2 99452 1 33701
2 99453 1 33701
2 99454 1 33701
2 99455 1 33701
2 99456 1 33702
2 99457 1 33702
2 99458 1 33702
2 99459 1 33710
2 99460 1 33710
2 99461 1 33718
2 99462 1 33718
2 99463 1 33718
2 99464 1 33718
2 99465 1 33733
2 99466 1 33733
2 99467 1 33762
2 99468 1 33762
2 99469 1 33764
2 99470 1 33764
2 99471 1 33764
2 99472 1 33769
2 99473 1 33769
2 99474 1 33797
2 99475 1 33797
2 99476 1 33805
2 99477 1 33805
2 99478 1 33805
2 99479 1 33822
2 99480 1 33822
2 99481 1 33828
2 99482 1 33828
2 99483 1 33828
2 99484 1 33828
2 99485 1 33828
2 99486 1 33828
2 99487 1 33828
2 99488 1 33828
2 99489 1 33828
2 99490 1 33828
2 99491 1 33828
2 99492 1 33828
2 99493 1 33828
2 99494 1 33828
2 99495 1 33828
2 99496 1 33828
2 99497 1 33828
2 99498 1 33828
2 99499 1 33828
2 99500 1 33828
2 99501 1 33828
2 99502 1 33828
2 99503 1 33828
2 99504 1 33828
2 99505 1 33828
2 99506 1 33828
2 99507 1 33828
2 99508 1 33828
2 99509 1 33828
2 99510 1 33828
2 99511 1 33828
2 99512 1 33828
2 99513 1 33828
2 99514 1 33828
2 99515 1 33828
2 99516 1 33828
2 99517 1 33828
2 99518 1 33828
2 99519 1 33829
2 99520 1 33829
2 99521 1 33829
2 99522 1 33830
2 99523 1 33830
2 99524 1 33830
2 99525 1 33839
2 99526 1 33839
2 99527 1 33839
2 99528 1 33839
2 99529 1 33841
2 99530 1 33841
2 99531 1 33844
2 99532 1 33844
2 99533 1 33844
2 99534 1 33844
2 99535 1 33844
2 99536 1 33844
2 99537 1 33844
2 99538 1 33852
2 99539 1 33852
2 99540 1 33852
2 99541 1 33852
2 99542 1 33885
2 99543 1 33885
2 99544 1 33885
2 99545 1 33885
2 99546 1 33885
2 99547 1 33885
2 99548 1 33886
2 99549 1 33886
2 99550 1 33886
2 99551 1 33887
2 99552 1 33887
2 99553 1 33890
2 99554 1 33890
2 99555 1 33901
2 99556 1 33901
2 99557 1 33915
2 99558 1 33915
2 99559 1 33928
2 99560 1 33928
2 99561 1 33928
2 99562 1 33930
2 99563 1 33930
2 99564 1 33931
2 99565 1 33931
2 99566 1 33931
2 99567 1 33931
2 99568 1 33935
2 99569 1 33935
2 99570 1 33944
2 99571 1 33944
2 99572 1 33959
2 99573 1 33959
2 99574 1 33964
2 99575 1 33964
2 99576 1 33964
2 99577 1 33964
2 99578 1 33964
2 99579 1 33964
2 99580 1 33964
2 99581 1 33964
2 99582 1 33964
2 99583 1 33964
2 99584 1 33964
2 99585 1 33964
2 99586 1 33964
2 99587 1 33966
2 99588 1 33966
2 99589 1 33969
2 99590 1 33969
2 99591 1 33969
2 99592 1 33969
2 99593 1 33969
2 99594 1 33969
2 99595 1 33969
2 99596 1 33969
2 99597 1 33969
2 99598 1 33969
2 99599 1 33969
2 99600 1 33969
2 99601 1 33969
2 99602 1 33969
2 99603 1 33969
2 99604 1 33969
2 99605 1 33969
2 99606 1 33970
2 99607 1 33970
2 99608 1 33970
2 99609 1 33970
2 99610 1 33970
2 99611 1 33970
2 99612 1 33970
2 99613 1 33972
2 99614 1 33972
2 99615 1 33989
2 99616 1 33989
2 99617 1 33989
2 99618 1 33989
2 99619 1 33989
2 99620 1 33989
2 99621 1 33990
2 99622 1 33990
2 99623 1 33990
2 99624 1 33991
2 99625 1 33991
2 99626 1 33991
2 99627 1 33991
2 99628 1 33991
2 99629 1 33991
2 99630 1 33991
2 99631 1 34000
2 99632 1 34000
2 99633 1 34001
2 99634 1 34001
2 99635 1 34001
2 99636 1 34001
2 99637 1 34013
2 99638 1 34013
2 99639 1 34013
2 99640 1 34022
2 99641 1 34022
2 99642 1 34022
2 99643 1 34022
2 99644 1 34028
2 99645 1 34028
2 99646 1 34028
2 99647 1 34028
2 99648 1 34028
2 99649 1 34028
2 99650 1 34028
2 99651 1 34028
2 99652 1 34028
2 99653 1 34028
2 99654 1 34028
2 99655 1 34028
2 99656 1 34028
2 99657 1 34028
2 99658 1 34028
2 99659 1 34028
2 99660 1 34028
2 99661 1 34028
2 99662 1 34028
2 99663 1 34028
2 99664 1 34028
2 99665 1 34028
2 99666 1 34028
2 99667 1 34028
2 99668 1 34028
2 99669 1 34028
2 99670 1 34028
2 99671 1 34028
2 99672 1 34028
2 99673 1 34028
2 99674 1 34028
2 99675 1 34029
2 99676 1 34029
2 99677 1 34037
2 99678 1 34037
2 99679 1 34037
2 99680 1 34046
2 99681 1 34046
2 99682 1 34047
2 99683 1 34047
2 99684 1 34055
2 99685 1 34055
2 99686 1 34059
2 99687 1 34059
2 99688 1 34060
2 99689 1 34060
2 99690 1 34060
2 99691 1 34060
2 99692 1 34060
2 99693 1 34060
2 99694 1 34060
2 99695 1 34060
2 99696 1 34068
2 99697 1 34068
2 99698 1 34068
2 99699 1 34068
2 99700 1 34068
2 99701 1 34068
2 99702 1 34068
2 99703 1 34068
2 99704 1 34076
2 99705 1 34076
2 99706 1 34076
2 99707 1 34076
2 99708 1 34076
2 99709 1 34077
2 99710 1 34077
2 99711 1 34078
2 99712 1 34078
2 99713 1 34086
2 99714 1 34086
2 99715 1 34086
2 99716 1 34097
2 99717 1 34097
2 99718 1 34114
2 99719 1 34114
2 99720 1 34114
2 99721 1 34114
2 99722 1 34114
2 99723 1 34114
2 99724 1 34114
2 99725 1 34114
2 99726 1 34114
2 99727 1 34114
2 99728 1 34114
2 99729 1 34114
2 99730 1 34115
2 99731 1 34115
2 99732 1 34115
2 99733 1 34115
2 99734 1 34116
2 99735 1 34116
2 99736 1 34118
2 99737 1 34118
2 99738 1 34119
2 99739 1 34119
2 99740 1 34119
2 99741 1 34119
2 99742 1 34119
2 99743 1 34119
2 99744 1 34119
2 99745 1 34119
2 99746 1 34119
2 99747 1 34119
2 99748 1 34127
2 99749 1 34127
2 99750 1 34127
2 99751 1 34127
2 99752 1 34127
2 99753 1 34127
2 99754 1 34127
2 99755 1 34127
2 99756 1 34127
2 99757 1 34128
2 99758 1 34128
2 99759 1 34129
2 99760 1 34129
2 99761 1 34129
2 99762 1 34129
2 99763 1 34143
2 99764 1 34143
2 99765 1 34143
2 99766 1 34152
2 99767 1 34152
2 99768 1 34152
2 99769 1 34152
2 99770 1 34152
2 99771 1 34153
2 99772 1 34153
2 99773 1 34153
2 99774 1 34164
2 99775 1 34164
2 99776 1 34164
2 99777 1 34165
2 99778 1 34165
2 99779 1 34174
2 99780 1 34174
2 99781 1 34175
2 99782 1 34175
2 99783 1 34175
2 99784 1 34175
2 99785 1 34175
2 99786 1 34175
2 99787 1 34175
2 99788 1 34180
2 99789 1 34180
2 99790 1 34182
2 99791 1 34182
2 99792 1 34182
2 99793 1 34182
2 99794 1 34206
2 99795 1 34206
2 99796 1 34206
2 99797 1 34206
2 99798 1 34206
2 99799 1 34217
2 99800 1 34217
2 99801 1 34222
2 99802 1 34222
2 99803 1 34224
2 99804 1 34224
2 99805 1 34239
2 99806 1 34239
2 99807 1 34239
2 99808 1 34239
2 99809 1 34239
2 99810 1 34239
2 99811 1 34239
2 99812 1 34256
2 99813 1 34256
2 99814 1 34257
2 99815 1 34257
2 99816 1 34258
2 99817 1 34258
2 99818 1 34267
2 99819 1 34267
2 99820 1 34271
2 99821 1 34271
2 99822 1 34274
2 99823 1 34274
2 99824 1 34274
2 99825 1 34274
2 99826 1 34274
2 99827 1 34282
2 99828 1 34282
2 99829 1 34282
2 99830 1 34282
2 99831 1 34282
2 99832 1 34282
2 99833 1 34282
2 99834 1 34288
2 99835 1 34288
2 99836 1 34290
2 99837 1 34290
2 99838 1 34300
2 99839 1 34300
2 99840 1 34300
2 99841 1 34308
2 99842 1 34308
2 99843 1 34308
2 99844 1 34308
2 99845 1 34317
2 99846 1 34317
2 99847 1 34317
2 99848 1 34317
2 99849 1 34317
2 99850 1 34325
2 99851 1 34325
2 99852 1 34330
2 99853 1 34330
2 99854 1 34330
2 99855 1 34333
2 99856 1 34333
2 99857 1 34333
2 99858 1 34366
2 99859 1 34366
2 99860 1 34373
2 99861 1 34373
2 99862 1 34373
2 99863 1 34373
2 99864 1 34373
2 99865 1 34373
2 99866 1 34387
2 99867 1 34387
2 99868 1 34387
2 99869 1 34388
2 99870 1 34388
2 99871 1 34388
2 99872 1 34388
2 99873 1 34412
2 99874 1 34412
2 99875 1 34416
2 99876 1 34416
2 99877 1 34417
2 99878 1 34417
2 99879 1 34418
2 99880 1 34418
2 99881 1 34449
2 99882 1 34449
2 99883 1 34457
2 99884 1 34457
2 99885 1 34458
2 99886 1 34458
2 99887 1 34499
2 99888 1 34499
2 99889 1 34522
2 99890 1 34522
2 99891 1 34525
2 99892 1 34525
2 99893 1 34525
2 99894 1 34540
2 99895 1 34540
2 99896 1 34540
2 99897 1 34549
2 99898 1 34549
2 99899 1 34549
2 99900 1 34559
2 99901 1 34559
2 99902 1 34559
2 99903 1 34572
2 99904 1 34572
2 99905 1 34573
2 99906 1 34573
2 99907 1 34573
2 99908 1 34576
2 99909 1 34576
2 99910 1 34576
2 99911 1 34577
2 99912 1 34577
2 99913 1 34584
2 99914 1 34584
2 99915 1 34584
2 99916 1 34584
2 99917 1 34585
2 99918 1 34585
2 99919 1 34585
2 99920 1 34593
2 99921 1 34593
2 99922 1 34601
2 99923 1 34601
2 99924 1 34610
2 99925 1 34610
2 99926 1 34610
2 99927 1 34610
2 99928 1 34610
2 99929 1 34619
2 99930 1 34619
2 99931 1 34623
2 99932 1 34623
2 99933 1 34623
2 99934 1 34634
2 99935 1 34634
2 99936 1 34642
2 99937 1 34642
2 99938 1 34650
2 99939 1 34650
2 99940 1 34654
2 99941 1 34654
2 99942 1 34655
2 99943 1 34655
2 99944 1 34655
2 99945 1 34659
2 99946 1 34659
2 99947 1 34659
2 99948 1 34672
2 99949 1 34672
2 99950 1 34672
2 99951 1 34698
2 99952 1 34698
2 99953 1 34698
2 99954 1 34700
2 99955 1 34700
2 99956 1 34701
2 99957 1 34701
2 99958 1 34709
2 99959 1 34709
2 99960 1 34709
2 99961 1 34718
2 99962 1 34718
2 99963 1 34729
2 99964 1 34729
2 99965 1 34729
2 99966 1 34729
2 99967 1 34729
2 99968 1 34729
2 99969 1 34729
2 99970 1 34729
2 99971 1 34729
2 99972 1 34730
2 99973 1 34730
2 99974 1 34739
2 99975 1 34739
2 99976 1 34739
2 99977 1 34744
2 99978 1 34744
2 99979 1 34762
2 99980 1 34762
2 99981 1 34762
2 99982 1 34794
2 99983 1 34794
2 99984 1 34794
2 99985 1 34794
2 99986 1 34795
2 99987 1 34795
2 99988 1 34795
2 99989 1 34795
2 99990 1 34795
2 99991 1 34795
2 99992 1 34796
2 99993 1 34796
2 99994 1 34799
2 99995 1 34799
2 99996 1 34808
2 99997 1 34808
2 99998 1 34808
2 99999 1 34808
2 100000 1 34808
2 100001 1 34808
2 100002 1 34808
2 100003 1 34808
2 100004 1 34808
2 100005 1 34808
2 100006 1 34808
2 100007 1 34808
2 100008 1 34808
2 100009 1 34808
2 100010 1 34808
2 100011 1 34808
2 100012 1 34808
2 100013 1 34808
2 100014 1 34808
2 100015 1 34808
2 100016 1 34808
2 100017 1 34808
2 100018 1 34808
2 100019 1 34808
2 100020 1 34808
2 100021 1 34808
2 100022 1 34808
2 100023 1 34808
2 100024 1 34808
2 100025 1 34808
2 100026 1 34808
2 100027 1 34808
2 100028 1 34808
2 100029 1 34812
2 100030 1 34812
2 100031 1 34812
2 100032 1 34812
2 100033 1 34812
2 100034 1 34820
2 100035 1 34820
2 100036 1 34820
2 100037 1 34820
2 100038 1 34820
2 100039 1 34832
2 100040 1 34832
2 100041 1 34832
2 100042 1 34832
2 100043 1 34834
2 100044 1 34834
2 100045 1 34834
2 100046 1 34834
2 100047 1 34837
2 100048 1 34837
2 100049 1 34849
2 100050 1 34849
2 100051 1 34853
2 100052 1 34853
2 100053 1 34859
2 100054 1 34859
2 100055 1 34863
2 100056 1 34863
2 100057 1 34883
2 100058 1 34883
2 100059 1 34926
2 100060 1 34926
2 100061 1 34926
2 100062 1 34926
2 100063 1 34935
2 100064 1 34935
2 100065 1 34935
2 100066 1 34936
2 100067 1 34936
2 100068 1 34957
2 100069 1 34957
2 100070 1 34957
2 100071 1 34971
2 100072 1 34971
2 100073 1 34971
2 100074 1 34971
2 100075 1 34971
2 100076 1 34971
2 100077 1 34972
2 100078 1 34972
2 100079 1 34972
2 100080 1 34972
2 100081 1 34973
2 100082 1 34973
2 100083 1 34973
2 100084 1 34977
2 100085 1 34977
2 100086 1 34983
2 100087 1 34983
2 100088 1 34983
2 100089 1 34983
2 100090 1 34983
2 100091 1 34986
2 100092 1 34986
2 100093 1 34986
2 100094 1 34986
2 100095 1 34986
2 100096 1 34986
2 100097 1 34986
2 100098 1 34986
2 100099 1 34986
2 100100 1 34986
2 100101 1 35002
2 100102 1 35002
2 100103 1 35020
2 100104 1 35020
2 100105 1 35040
2 100106 1 35040
2 100107 1 35040
2 100108 1 35041
2 100109 1 35041
2 100110 1 35044
2 100111 1 35044
2 100112 1 35044
2 100113 1 35044
2 100114 1 35044
2 100115 1 35045
2 100116 1 35045
2 100117 1 35065
2 100118 1 35065
2 100119 1 35065
2 100120 1 35065
2 100121 1 35065
2 100122 1 35075
2 100123 1 35075
2 100124 1 35075
2 100125 1 35075
2 100126 1 35075
2 100127 1 35087
2 100128 1 35087
2 100129 1 35088
2 100130 1 35088
2 100131 1 35108
2 100132 1 35108
2 100133 1 35108
2 100134 1 35108
2 100135 1 35109
2 100136 1 35109
2 100137 1 35118
2 100138 1 35118
2 100139 1 35122
2 100140 1 35122
2 100141 1 35122
2 100142 1 35122
2 100143 1 35122
2 100144 1 35122
2 100145 1 35123
2 100146 1 35123
2 100147 1 35140
2 100148 1 35140
2 100149 1 35141
2 100150 1 35141
2 100151 1 35149
2 100152 1 35149
2 100153 1 35149
2 100154 1 35149
2 100155 1 35149
2 100156 1 35150
2 100157 1 35150
2 100158 1 35154
2 100159 1 35154
2 100160 1 35154
2 100161 1 35169
2 100162 1 35169
2 100163 1 35169
2 100164 1 35169
2 100165 1 35176
2 100166 1 35176
2 100167 1 35177
2 100168 1 35177
2 100169 1 35202
2 100170 1 35202
2 100171 1 35205
2 100172 1 35205
2 100173 1 35251
2 100174 1 35251
2 100175 1 35252
2 100176 1 35252
2 100177 1 35274
2 100178 1 35274
2 100179 1 35282
2 100180 1 35282
2 100181 1 35304
2 100182 1 35304
2 100183 1 35328
2 100184 1 35328
2 100185 1 35329
2 100186 1 35329
2 100187 1 35329
2 100188 1 35344
2 100189 1 35344
2 100190 1 35344
2 100191 1 35344
2 100192 1 35348
2 100193 1 35348
2 100194 1 35358
2 100195 1 35358
2 100196 1 35365
2 100197 1 35365
2 100198 1 35372
2 100199 1 35372
2 100200 1 35372
2 100201 1 35396
2 100202 1 35396
2 100203 1 35396
2 100204 1 35396
2 100205 1 35396
2 100206 1 35396
2 100207 1 35396
2 100208 1 35404
2 100209 1 35404
2 100210 1 35404
2 100211 1 35405
2 100212 1 35405
2 100213 1 35415
2 100214 1 35415
2 100215 1 35429
2 100216 1 35429
2 100217 1 35429
2 100218 1 35430
2 100219 1 35430
2 100220 1 35430
2 100221 1 35452
2 100222 1 35452
2 100223 1 35452
2 100224 1 35483
2 100225 1 35483
2 100226 1 35483
2 100227 1 35483
2 100228 1 35483
2 100229 1 35483
2 100230 1 35483
2 100231 1 35483
2 100232 1 35483
2 100233 1 35483
2 100234 1 35483
2 100235 1 35483
2 100236 1 35483
2 100237 1 35483
2 100238 1 35483
2 100239 1 35483
2 100240 1 35483
2 100241 1 35483
2 100242 1 35483
2 100243 1 35483
2 100244 1 35483
2 100245 1 35483
2 100246 1 35483
2 100247 1 35483
2 100248 1 35483
2 100249 1 35483
2 100250 1 35483
2 100251 1 35483
2 100252 1 35483
2 100253 1 35483
2 100254 1 35484
2 100255 1 35484
2 100256 1 35484
2 100257 1 35490
2 100258 1 35490
2 100259 1 35492
2 100260 1 35492
2 100261 1 35492
2 100262 1 35492
2 100263 1 35493
2 100264 1 35493
2 100265 1 35493
2 100266 1 35500
2 100267 1 35500
2 100268 1 35500
2 100269 1 35504
2 100270 1 35504
2 100271 1 35515
2 100272 1 35515
2 100273 1 35528
2 100274 1 35528
2 100275 1 35528
2 100276 1 35528
2 100277 1 35528
2 100278 1 35528
2 100279 1 35528
2 100280 1 35528
2 100281 1 35530
2 100282 1 35530
2 100283 1 35530
2 100284 1 35530
2 100285 1 35531
2 100286 1 35531
2 100287 1 35531
2 100288 1 35531
2 100289 1 35531
2 100290 1 35531
2 100291 1 35531
2 100292 1 35538
2 100293 1 35538
2 100294 1 35539
2 100295 1 35539
2 100296 1 35539
2 100297 1 35555
2 100298 1 35555
2 100299 1 35555
2 100300 1 35555
2 100301 1 35555
2 100302 1 35555
2 100303 1 35560
2 100304 1 35560
2 100305 1 35560
2 100306 1 35561
2 100307 1 35561
2 100308 1 35561
2 100309 1 35577
2 100310 1 35577
2 100311 1 35593
2 100312 1 35593
2 100313 1 35594
2 100314 1 35594
2 100315 1 35602
2 100316 1 35602
2 100317 1 35602
2 100318 1 35603
2 100319 1 35603
2 100320 1 35612
2 100321 1 35612
2 100322 1 35630
2 100323 1 35630
2 100324 1 35630
2 100325 1 35667
2 100326 1 35667
2 100327 1 35671
2 100328 1 35671
2 100329 1 35675
2 100330 1 35675
2 100331 1 35685
2 100332 1 35685
2 100333 1 35690
2 100334 1 35690
2 100335 1 35690
2 100336 1 35690
2 100337 1 35690
2 100338 1 35700
2 100339 1 35700
2 100340 1 35719
2 100341 1 35719
2 100342 1 35729
2 100343 1 35729
2 100344 1 35737
2 100345 1 35737
2 100346 1 35737
2 100347 1 35738
2 100348 1 35738
2 100349 1 35750
2 100350 1 35750
2 100351 1 35772
2 100352 1 35772
2 100353 1 35772
2 100354 1 35773
2 100355 1 35773
2 100356 1 35774
2 100357 1 35774
2 100358 1 35774
2 100359 1 35774
2 100360 1 35774
2 100361 1 35775
2 100362 1 35775
2 100363 1 35775
2 100364 1 35775
2 100365 1 35775
2 100366 1 35775
2 100367 1 35775
2 100368 1 35775
2 100369 1 35812
2 100370 1 35812
2 100371 1 35821
2 100372 1 35821
2 100373 1 35840
2 100374 1 35840
2 100375 1 35841
2 100376 1 35841
2 100377 1 35841
2 100378 1 35843
2 100379 1 35843
2 100380 1 35862
2 100381 1 35862
2 100382 1 35870
2 100383 1 35870
2 100384 1 35870
2 100385 1 35878
2 100386 1 35878
2 100387 1 35879
2 100388 1 35879
2 100389 1 35885
2 100390 1 35885
2 100391 1 35902
2 100392 1 35902
2 100393 1 35906
2 100394 1 35906
2 100395 1 35906
2 100396 1 35906
2 100397 1 35907
2 100398 1 35907
2 100399 1 35915
2 100400 1 35915
2 100401 1 35938
2 100402 1 35938
2 100403 1 35957
2 100404 1 35957
2 100405 1 35957
2 100406 1 35957
2 100407 1 35957
2 100408 1 35957
2 100409 1 35957
2 100410 1 35957
2 100411 1 35957
2 100412 1 35957
2 100413 1 35957
2 100414 1 35957
2 100415 1 35957
2 100416 1 35958
2 100417 1 35958
2 100418 1 35958
2 100419 1 35958
2 100420 1 35958
2 100421 1 35958
2 100422 1 35958
2 100423 1 35962
2 100424 1 35962
2 100425 1 35968
2 100426 1 35968
2 100427 1 35968
2 100428 1 35991
2 100429 1 35991
2 100430 1 36020
2 100431 1 36020
2 100432 1 36020
2 100433 1 36020
2 100434 1 36021
2 100435 1 36021
2 100436 1 36027
2 100437 1 36027
2 100438 1 36027
2 100439 1 36027
2 100440 1 36042
2 100441 1 36042
2 100442 1 36043
2 100443 1 36043
2 100444 1 36062
2 100445 1 36062
2 100446 1 36066
2 100447 1 36066
2 100448 1 36066
2 100449 1 36081
2 100450 1 36081
2 100451 1 36091
2 100452 1 36091
2 100453 1 36102
2 100454 1 36102
2 100455 1 36103
2 100456 1 36103
2 100457 1 36104
2 100458 1 36104
2 100459 1 36104
2 100460 1 36106
2 100461 1 36106
2 100462 1 36143
2 100463 1 36143
2 100464 1 36187
2 100465 1 36187
2 100466 1 36187
2 100467 1 36188
2 100468 1 36188
2 100469 1 36200
2 100470 1 36200
2 100471 1 36200
2 100472 1 36203
2 100473 1 36203
2 100474 1 36203
2 100475 1 36218
2 100476 1 36218
2 100477 1 36218
2 100478 1 36218
2 100479 1 36222
2 100480 1 36222
2 100481 1 36222
2 100482 1 36243
2 100483 1 36243
2 100484 1 36246
2 100485 1 36246
2 100486 1 36247
2 100487 1 36247
2 100488 1 36248
2 100489 1 36248
2 100490 1 36259
2 100491 1 36259
2 100492 1 36260
2 100493 1 36260
2 100494 1 36260
2 100495 1 36260
2 100496 1 36272
2 100497 1 36272
2 100498 1 36272
2 100499 1 36272
2 100500 1 36273
2 100501 1 36273
2 100502 1 36274
2 100503 1 36274
2 100504 1 36274
2 100505 1 36287
2 100506 1 36287
2 100507 1 36287
2 100508 1 36287
2 100509 1 36287
2 100510 1 36288
2 100511 1 36288
2 100512 1 36291
2 100513 1 36291
2 100514 1 36291
2 100515 1 36291
2 100516 1 36291
2 100517 1 36327
2 100518 1 36327
2 100519 1 36327
2 100520 1 36327
2 100521 1 36327
2 100522 1 36342
2 100523 1 36342
2 100524 1 36344
2 100525 1 36344
2 100526 1 36344
2 100527 1 36351
2 100528 1 36351
2 100529 1 36352
2 100530 1 36352
2 100531 1 36354
2 100532 1 36354
2 100533 1 36363
2 100534 1 36363
2 100535 1 36371
2 100536 1 36371
2 100537 1 36378
2 100538 1 36378
2 100539 1 36378
2 100540 1 36378
2 100541 1 36379
2 100542 1 36379
2 100543 1 36389
2 100544 1 36389
2 100545 1 36391
2 100546 1 36391
2 100547 1 36400
2 100548 1 36400
2 100549 1 36400
2 100550 1 36400
2 100551 1 36400
2 100552 1 36400
2 100553 1 36400
2 100554 1 36400
2 100555 1 36400
2 100556 1 36410
2 100557 1 36410
2 100558 1 36410
2 100559 1 36410
2 100560 1 36411
2 100561 1 36411
2 100562 1 36411
2 100563 1 36411
2 100564 1 36419
2 100565 1 36419
2 100566 1 36420
2 100567 1 36420
2 100568 1 36429
2 100569 1 36429
2 100570 1 36454
2 100571 1 36454
2 100572 1 36454
2 100573 1 36454
2 100574 1 36454
2 100575 1 36454
2 100576 1 36454
2 100577 1 36454
2 100578 1 36454
2 100579 1 36454
2 100580 1 36454
2 100581 1 36455
2 100582 1 36455
2 100583 1 36455
2 100584 1 36455
2 100585 1 36473
2 100586 1 36473
2 100587 1 36475
2 100588 1 36475
2 100589 1 36475
2 100590 1 36475
2 100591 1 36475
2 100592 1 36475
2 100593 1 36475
2 100594 1 36475
2 100595 1 36475
2 100596 1 36475
2 100597 1 36478
2 100598 1 36478
2 100599 1 36478
2 100600 1 36478
2 100601 1 36482
2 100602 1 36482
2 100603 1 36482
2 100604 1 36482
2 100605 1 36482
2 100606 1 36486
2 100607 1 36486
2 100608 1 36486
2 100609 1 36496
2 100610 1 36496
2 100611 1 36496
2 100612 1 36504
2 100613 1 36504
2 100614 1 36506
2 100615 1 36506
2 100616 1 36507
2 100617 1 36507
2 100618 1 36528
2 100619 1 36528
2 100620 1 36528
2 100621 1 36528
2 100622 1 36528
2 100623 1 36528
2 100624 1 36528
2 100625 1 36528
2 100626 1 36528
2 100627 1 36528
2 100628 1 36528
2 100629 1 36535
2 100630 1 36535
2 100631 1 36535
2 100632 1 36535
2 100633 1 36536
2 100634 1 36536
2 100635 1 36536
2 100636 1 36536
2 100637 1 36536
2 100638 1 36536
2 100639 1 36536
2 100640 1 36536
2 100641 1 36536
2 100642 1 36546
2 100643 1 36546
2 100644 1 36553
2 100645 1 36553
2 100646 1 36563
2 100647 1 36563
2 100648 1 36563
2 100649 1 36578
2 100650 1 36578
2 100651 1 36587
2 100652 1 36587
2 100653 1 36588
2 100654 1 36588
2 100655 1 36599
2 100656 1 36599
2 100657 1 36600
2 100658 1 36600
2 100659 1 36615
2 100660 1 36615
2 100661 1 36616
2 100662 1 36616
2 100663 1 36616
2 100664 1 36616
2 100665 1 36616
2 100666 1 36616
2 100667 1 36626
2 100668 1 36626
2 100669 1 36626
2 100670 1 36629
2 100671 1 36629
2 100672 1 36629
2 100673 1 36629
2 100674 1 36629
2 100675 1 36629
2 100676 1 36629
2 100677 1 36629
2 100678 1 36629
2 100679 1 36629
2 100680 1 36629
2 100681 1 36629
2 100682 1 36629
2 100683 1 36630
2 100684 1 36630
2 100685 1 36630
2 100686 1 36630
2 100687 1 36630
2 100688 1 36630
2 100689 1 36630
2 100690 1 36630
2 100691 1 36630
2 100692 1 36630
2 100693 1 36630
2 100694 1 36630
2 100695 1 36630
2 100696 1 36630
2 100697 1 36630
2 100698 1 36630
2 100699 1 36630
2 100700 1 36634
2 100701 1 36634
2 100702 1 36634
2 100703 1 36634
2 100704 1 36634
2 100705 1 36634
2 100706 1 36635
2 100707 1 36635
2 100708 1 36655
2 100709 1 36655
2 100710 1 36660
2 100711 1 36660
2 100712 1 36660
2 100713 1 36660
2 100714 1 36672
2 100715 1 36672
2 100716 1 36672
2 100717 1 36680
2 100718 1 36680
2 100719 1 36680
2 100720 1 36700
2 100721 1 36700
2 100722 1 36701
2 100723 1 36701
2 100724 1 36701
2 100725 1 36701
2 100726 1 36702
2 100727 1 36702
2 100728 1 36711
2 100729 1 36711
2 100730 1 36718
2 100731 1 36718
2 100732 1 36719
2 100733 1 36719
2 100734 1 36734
2 100735 1 36734
2 100736 1 36734
2 100737 1 36734
2 100738 1 36747
2 100739 1 36747
2 100740 1 36747
2 100741 1 36747
2 100742 1 36779
2 100743 1 36779
2 100744 1 36792
2 100745 1 36792
2 100746 1 36793
2 100747 1 36793
2 100748 1 36793
2 100749 1 36826
2 100750 1 36826
2 100751 1 36827
2 100752 1 36827
2 100753 1 36827
2 100754 1 36829
2 100755 1 36829
2 100756 1 36829
2 100757 1 36831
2 100758 1 36831
2 100759 1 36832
2 100760 1 36832
2 100761 1 36832
2 100762 1 36832
2 100763 1 36832
2 100764 1 36832
2 100765 1 36833
2 100766 1 36833
2 100767 1 36833
2 100768 1 36833
2 100769 1 36836
2 100770 1 36836
2 100771 1 36836
2 100772 1 36839
2 100773 1 36839
2 100774 1 36857
2 100775 1 36857
2 100776 1 36857
2 100777 1 36857
2 100778 1 36866
2 100779 1 36866
2 100780 1 36866
2 100781 1 36878
2 100782 1 36878
2 100783 1 36886
2 100784 1 36886
2 100785 1 36900
2 100786 1 36900
2 100787 1 36904
2 100788 1 36904
2 100789 1 36915
2 100790 1 36915
2 100791 1 36915
2 100792 1 36915
2 100793 1 36915
2 100794 1 36915
2 100795 1 36915
2 100796 1 36915
2 100797 1 36927
2 100798 1 36927
2 100799 1 36935
2 100800 1 36935
2 100801 1 36935
2 100802 1 36943
2 100803 1 36943
2 100804 1 36943
2 100805 1 36944
2 100806 1 36944
2 100807 1 36944
2 100808 1 36944
2 100809 1 36944
2 100810 1 36944
2 100811 1 36944
2 100812 1 36944
2 100813 1 36944
2 100814 1 36944
2 100815 1 36944
2 100816 1 36944
2 100817 1 36947
2 100818 1 36947
2 100819 1 36964
2 100820 1 36964
2 100821 1 36966
2 100822 1 36966
2 100823 1 36966
2 100824 1 36966
2 100825 1 36966
2 100826 1 36966
2 100827 1 36972
2 100828 1 36972
2 100829 1 36972
2 100830 1 36973
2 100831 1 36973
2 100832 1 36984
2 100833 1 36984
2 100834 1 36992
2 100835 1 36992
2 100836 1 36992
2 100837 1 36992
2 100838 1 37005
2 100839 1 37005
2 100840 1 37013
2 100841 1 37013
2 100842 1 37013
2 100843 1 37013
2 100844 1 37013
2 100845 1 37014
2 100846 1 37014
2 100847 1 37016
2 100848 1 37016
2 100849 1 37017
2 100850 1 37017
2 100851 1 37029
2 100852 1 37029
2 100853 1 37029
2 100854 1 37033
2 100855 1 37033
2 100856 1 37039
2 100857 1 37039
2 100858 1 37054
2 100859 1 37054
2 100860 1 37061
2 100861 1 37061
2 100862 1 37075
2 100863 1 37075
2 100864 1 37075
2 100865 1 37090
2 100866 1 37090
2 100867 1 37124
2 100868 1 37124
2 100869 1 37124
2 100870 1 37132
2 100871 1 37132
2 100872 1 37158
2 100873 1 37158
2 100874 1 37158
2 100875 1 37159
2 100876 1 37159
2 100877 1 37159
2 100878 1 37159
2 100879 1 37159
2 100880 1 37159
2 100881 1 37161
2 100882 1 37161
2 100883 1 37161
2 100884 1 37164
2 100885 1 37164
2 100886 1 37187
2 100887 1 37187
2 100888 1 37205
2 100889 1 37205
2 100890 1 37206
2 100891 1 37206
2 100892 1 37206
2 100893 1 37212
2 100894 1 37212
2 100895 1 37213
2 100896 1 37213
2 100897 1 37213
2 100898 1 37213
2 100899 1 37213
2 100900 1 37214
2 100901 1 37214
2 100902 1 37214
2 100903 1 37214
2 100904 1 37214
2 100905 1 37214
2 100906 1 37214
2 100907 1 37214
2 100908 1 37214
2 100909 1 37216
2 100910 1 37216
2 100911 1 37216
2 100912 1 37236
2 100913 1 37236
2 100914 1 37266
2 100915 1 37266
2 100916 1 37267
2 100917 1 37267
2 100918 1 37287
2 100919 1 37287
2 100920 1 37291
2 100921 1 37291
2 100922 1 37298
2 100923 1 37298
2 100924 1 37306
2 100925 1 37306
2 100926 1 37306
2 100927 1 37306
2 100928 1 37306
2 100929 1 37338
2 100930 1 37338
2 100931 1 37443
2 100932 1 37443
2 100933 1 37446
2 100934 1 37446
2 100935 1 37446
2 100936 1 37457
2 100937 1 37457
2 100938 1 37465
2 100939 1 37465
2 100940 1 37466
2 100941 1 37466
2 100942 1 37466
2 100943 1 37510
2 100944 1 37510
2 100945 1 37513
2 100946 1 37513
2 100947 1 37513
2 100948 1 37525
2 100949 1 37525
2 100950 1 37528
2 100951 1 37528
2 100952 1 37577
2 100953 1 37577
2 100954 1 37577
2 100955 1 37594
2 100956 1 37594
2 100957 1 37594
2 100958 1 37603
2 100959 1 37603
2 100960 1 37635
2 100961 1 37635
2 100962 1 37638
2 100963 1 37638
2 100964 1 37722
2 100965 1 37722
2 100966 1 37723
2 100967 1 37723
2 100968 1 37751
2 100969 1 37751
2 100970 1 37812
2 100971 1 37812
2 100972 1 37812
2 100973 1 37813
2 100974 1 37813
2 100975 1 37886
2 100976 1 37886
2 100977 1 37916
2 100978 1 37916
2 100979 1 37916
2 100980 1 37917
2 100981 1 37917
2 100982 1 37931
2 100983 1 37931
2 100984 1 37932
2 100985 1 37932
2 100986 1 37933
2 100987 1 37933
2 100988 1 37933
2 100989 1 37933
2 100990 1 37933
2 100991 1 37933
2 100992 1 37933
2 100993 1 37933
2 100994 1 37933
2 100995 1 37933
2 100996 1 37935
2 100997 1 37935
2 100998 1 37941
2 100999 1 37941
2 101000 1 37942
2 101001 1 37942
2 101002 1 37963
2 101003 1 37963
2 101004 1 37998
2 101005 1 37998
2 101006 1 38026
2 101007 1 38026
2 101008 1 38085
2 101009 1 38085
2 101010 1 38085
2 101011 1 38104
2 101012 1 38104
2 101013 1 38105
2 101014 1 38105
2 101015 1 38114
2 101016 1 38114
2 101017 1 38115
2 101018 1 38115
2 101019 1 38124
2 101020 1 38124
2 101021 1 38131
2 101022 1 38131
2 101023 1 38131
2 101024 1 38132
2 101025 1 38132
2 101026 1 38150
2 101027 1 38150
2 101028 1 38152
2 101029 1 38152
2 101030 1 38168
2 101031 1 38168
2 101032 1 38194
2 101033 1 38194
2 101034 1 38194
2 101035 1 38194
2 101036 1 38194
2 101037 1 38194
2 101038 1 38194
2 101039 1 38197
2 101040 1 38197
2 101041 1 38197
2 101042 1 38204
2 101043 1 38204
2 101044 1 38217
2 101045 1 38217
2 101046 1 38217
2 101047 1 38232
2 101048 1 38232
2 101049 1 38232
2 101050 1 38232
2 101051 1 38236
2 101052 1 38236
2 101053 1 38248
2 101054 1 38248
2 101055 1 38248
2 101056 1 38248
2 101057 1 38275
2 101058 1 38275
2 101059 1 38275
2 101060 1 38276
2 101061 1 38276
2 101062 1 38276
2 101063 1 38276
2 101064 1 38276
2 101065 1 38280
2 101066 1 38280
2 101067 1 38286
2 101068 1 38286
2 101069 1 38300
2 101070 1 38300
2 101071 1 38301
2 101072 1 38301
2 101073 1 38305
2 101074 1 38305
2 101075 1 38317
2 101076 1 38317
2 101077 1 38318
2 101078 1 38318
2 101079 1 38318
2 101080 1 38365
2 101081 1 38365
2 101082 1 38384
2 101083 1 38384
2 101084 1 38407
2 101085 1 38407
2 101086 1 38431
2 101087 1 38431
2 101088 1 38431
2 101089 1 38432
2 101090 1 38432
2 101091 1 38457
2 101092 1 38457
2 101093 1 38471
2 101094 1 38471
2 101095 1 38616
2 101096 1 38616
2 101097 1 38616
2 101098 1 38627
2 101099 1 38627
2 101100 1 38628
2 101101 1 38628
2 101102 1 38667
2 101103 1 38667
2 101104 1 38669
2 101105 1 38669
2 101106 1 38684
2 101107 1 38684
2 101108 1 38684
2 101109 1 38736
2 101110 1 38736
2 101111 1 38748
2 101112 1 38748
2 101113 1 38748
2 101114 1 38748
2 101115 1 38749
2 101116 1 38749
2 101117 1 38749
2 101118 1 38750
2 101119 1 38750
2 101120 1 38767
2 101121 1 38767
2 101122 1 38784
2 101123 1 38784
2 101124 1 38785
2 101125 1 38785
2 101126 1 38786
2 101127 1 38786
2 101128 1 38788
2 101129 1 38788
2 101130 1 38824
2 101131 1 38824
2 101132 1 38841
2 101133 1 38841
2 101134 1 38842
2 101135 1 38842
2 101136 1 38871
2 101137 1 38871
2 101138 1 38888
2 101139 1 38888
2 101140 1 38929
2 101141 1 38929
2 101142 1 38973
2 101143 1 38973
2 101144 1 38977
2 101145 1 38977
2 101146 1 38977
2 101147 1 38984
2 101148 1 38984
2 101149 1 38984
2 101150 1 39015
2 101151 1 39015
2 101152 1 39023
2 101153 1 39023
2 101154 1 39051
2 101155 1 39051
2 101156 1 39067
2 101157 1 39067
2 101158 1 39101
2 101159 1 39101
2 101160 1 39153
2 101161 1 39153
2 101162 1 39153
2 101163 1 39162
2 101164 1 39162
2 101165 1 39210
2 101166 1 39210
2 101167 1 39210
2 101168 1 39218
2 101169 1 39218
2 101170 1 39224
2 101171 1 39224
2 101172 1 39225
2 101173 1 39225
2 101174 1 39226
2 101175 1 39226
2 101176 1 39255
2 101177 1 39255
2 101178 1 39255
2 101179 1 39255
2 101180 1 39256
2 101181 1 39256
2 101182 1 39272
2 101183 1 39272
2 101184 1 39272
2 101185 1 39370
2 101186 1 39370
2 101187 1 39373
2 101188 1 39373
2 101189 1 39402
2 101190 1 39402
2 101191 1 39423
2 101192 1 39423
2 101193 1 39450
2 101194 1 39450
2 101195 1 39450
2 101196 1 39450
2 101197 1 39454
2 101198 1 39454
2 101199 1 39473
2 101200 1 39473
2 101201 1 39473
2 101202 1 39482
2 101203 1 39482
2 101204 1 39563
2 101205 1 39563
2 101206 1 39581
2 101207 1 39581
2 101208 1 39596
2 101209 1 39596
2 101210 1 39608
2 101211 1 39608
2 101212 1 39627
2 101213 1 39627
2 101214 1 39631
2 101215 1 39631
2 101216 1 39672
2 101217 1 39672
2 101218 1 39722
2 101219 1 39722
2 101220 1 39724
2 101221 1 39724
2 101222 1 39736
2 101223 1 39736
2 101224 1 39756
2 101225 1 39756
2 101226 1 39855
2 101227 1 39855
2 101228 1 39917
2 101229 1 39917
2 101230 1 39932
2 101231 1 39932
2 101232 1 39953
2 101233 1 39953
2 101234 1 40030
2 101235 1 40030
2 101236 1 40033
2 101237 1 40033
2 101238 1 40082
2 101239 1 40082
2 101240 1 40171
2 101241 1 40171
2 101242 1 40172
2 101243 1 40172
2 101244 1 40179
2 101245 1 40179
2 101246 1 40189
2 101247 1 40189
2 101248 1 40189
2 101249 1 40230
2 101250 1 40230
2 101251 1 40232
2 101252 1 40232
2 101253 1 40318
2 101254 1 40318
2 101255 1 40321
2 101256 1 40321
2 101257 1 40330
2 101258 1 40330
2 101259 1 40330
2 101260 1 40332
2 101261 1 40332
2 101262 1 40381
2 101263 1 40381
2 101264 1 40381
2 101265 1 40381
2 101266 1 40389
2 101267 1 40389
2 101268 1 40404
2 101269 1 40404
2 101270 1 40404
2 101271 1 40404
2 101272 1 40416
2 101273 1 40416
2 101274 1 40417
2 101275 1 40417
2 101276 1 40425
2 101277 1 40425
2 101278 1 40425
2 101279 1 40429
2 101280 1 40429
2 101281 1 40433
2 101282 1 40433
2 101283 1 40540
2 101284 1 40540
2 101285 1 40560
2 101286 1 40560
2 101287 1 40575
2 101288 1 40575
2 101289 1 40585
2 101290 1 40585
2 101291 1 40593
2 101292 1 40593
2 101293 1 40606
2 101294 1 40606
2 101295 1 40619
2 101296 1 40619
2 101297 1 40631
2 101298 1 40631
2 101299 1 40632
2 101300 1 40632
2 101301 1 40642
2 101302 1 40642
2 101303 1 40642
2 101304 1 40706
2 101305 1 40706
2 101306 1 40801
2 101307 1 40801
2 101308 1 40870
2 101309 1 40870
2 101310 1 40870
2 101311 1 40897
2 101312 1 40897
2 101313 1 40907
2 101314 1 40907
2 101315 1 40913
2 101316 1 40913
2 101317 1 40913
2 101318 1 40913
2 101319 1 40913
2 101320 1 40913
2 101321 1 40913
2 101322 1 40913
2 101323 1 40913
2 101324 1 40913
2 101325 1 40913
2 101326 1 40913
2 101327 1 40913
2 101328 1 40914
2 101329 1 40914
2 101330 1 40923
2 101331 1 40923
2 101332 1 40923
2 101333 1 40923
2 101334 1 40924
2 101335 1 40924
2 101336 1 40944
2 101337 1 40944
2 101338 1 40958
2 101339 1 40958
2 101340 1 41024
2 101341 1 41024
2 101342 1 41059
2 101343 1 41059
2 101344 1 41063
2 101345 1 41063
2 101346 1 41069
2 101347 1 41069
2 101348 1 41071
2 101349 1 41071
2 101350 1 41095
2 101351 1 41095
2 101352 1 41095
2 101353 1 41102
2 101354 1 41102
2 101355 1 41153
2 101356 1 41153
2 101357 1 41185
2 101358 1 41185
2 101359 1 41185
2 101360 1 41186
2 101361 1 41186
2 101362 1 41186
2 101363 1 41186
2 101364 1 41204
2 101365 1 41204
2 101366 1 41218
2 101367 1 41218
2 101368 1 41218
2 101369 1 41222
2 101370 1 41222
2 101371 1 41222
2 101372 1 41222
2 101373 1 41232
2 101374 1 41232
2 101375 1 41235
2 101376 1 41235
2 101377 1 41254
2 101378 1 41254
2 101379 1 41265
2 101380 1 41265
2 101381 1 41266
2 101382 1 41266
2 101383 1 41266
2 101384 1 41278
2 101385 1 41278
2 101386 1 41335
2 101387 1 41335
2 101388 1 41343
2 101389 1 41343
2 101390 1 41343
2 101391 1 41343
2 101392 1 41343
2 101393 1 41344
2 101394 1 41344
2 101395 1 41375
2 101396 1 41375
2 101397 1 41378
2 101398 1 41378
2 101399 1 41404
2 101400 1 41404
2 101401 1 41412
2 101402 1 41412
2 101403 1 41450
2 101404 1 41450
2 101405 1 41476
2 101406 1 41476
2 101407 1 41592
2 101408 1 41592
2 101409 1 41635
2 101410 1 41635
2 101411 1 41639
2 101412 1 41639
2 101413 1 41639
2 101414 1 41639
2 101415 1 41657
2 101416 1 41657
2 101417 1 41657
2 101418 1 41658
2 101419 1 41658
2 101420 1 41665
2 101421 1 41665
2 101422 1 41694
2 101423 1 41694
2 101424 1 41694
2 101425 1 41694
2 101426 1 41694
2 101427 1 41703
2 101428 1 41703
2 101429 1 41709
2 101430 1 41709
2 101431 1 41714
2 101432 1 41714
2 101433 1 41714
2 101434 1 41737
2 101435 1 41737
2 101436 1 41737
2 101437 1 41740
2 101438 1 41740
2 101439 1 41740
2 101440 1 41740
2 101441 1 41740
2 101442 1 41740
2 101443 1 41740
2 101444 1 41740
2 101445 1 41740
2 101446 1 41740
2 101447 1 41740
2 101448 1 41740
2 101449 1 41740
2 101450 1 41752
2 101451 1 41752
2 101452 1 41752
2 101453 1 41752
2 101454 1 41761
2 101455 1 41761
2 101456 1 41774
2 101457 1 41774
2 101458 1 41774
2 101459 1 41783
2 101460 1 41783
2 101461 1 41783
2 101462 1 41795
2 101463 1 41795
2 101464 1 41796
2 101465 1 41796
2 101466 1 41807
2 101467 1 41807
2 101468 1 41807
2 101469 1 41824
2 101470 1 41824
2 101471 1 41826
2 101472 1 41826
2 101473 1 41849
2 101474 1 41849
2 101475 1 41849
2 101476 1 41887
2 101477 1 41887
2 101478 1 41888
2 101479 1 41888
2 101480 1 41892
2 101481 1 41892
2 101482 1 41903
2 101483 1 41903
2 101484 1 41920
2 101485 1 41920
2 101486 1 41931
2 101487 1 41931
2 101488 1 42040
2 101489 1 42040
2 101490 1 42076
2 101491 1 42076
2 101492 1 42084
2 101493 1 42084
2 101494 1 42086
2 101495 1 42086
2 101496 1 42086
2 101497 1 42094
2 101498 1 42094
2 101499 1 42110
2 101500 1 42110
2 101501 1 42110
2 101502 1 42162
2 101503 1 42162
2 101504 1 42164
2 101505 1 42164
2 101506 1 42202
2 101507 1 42202
2 101508 1 42202
2 101509 1 42203
2 101510 1 42203
2 101511 1 42203
2 101512 1 42203
2 101513 1 42203
2 101514 1 42203
2 101515 1 42203
2 101516 1 42204
2 101517 1 42204
2 101518 1 42209
2 101519 1 42209
2 101520 1 42225
2 101521 1 42225
2 101522 1 42240
2 101523 1 42240
2 101524 1 42240
2 101525 1 42244
2 101526 1 42244
2 101527 1 42244
2 101528 1 42244
2 101529 1 42244
2 101530 1 42244
2 101531 1 42244
2 101532 1 42244
2 101533 1 42245
2 101534 1 42245
2 101535 1 42273
2 101536 1 42273
2 101537 1 42273
2 101538 1 42282
2 101539 1 42282
2 101540 1 42282
2 101541 1 42282
2 101542 1 42282
2 101543 1 42282
2 101544 1 42285
2 101545 1 42285
2 101546 1 42285
2 101547 1 42285
2 101548 1 42285
2 101549 1 42285
2 101550 1 42285
2 101551 1 42286
2 101552 1 42286
2 101553 1 42286
2 101554 1 42287
2 101555 1 42287
2 101556 1 42305
2 101557 1 42305
2 101558 1 42305
2 101559 1 42306
2 101560 1 42306
2 101561 1 42307
2 101562 1 42307
2 101563 1 42307
2 101564 1 42318
2 101565 1 42318
2 101566 1 42338
2 101567 1 42338
2 101568 1 42340
2 101569 1 42340
2 101570 1 42343
2 101571 1 42343
2 101572 1 42343
2 101573 1 42343
2 101574 1 42347
2 101575 1 42347
2 101576 1 42347
2 101577 1 42347
2 101578 1 42347
2 101579 1 42360
2 101580 1 42360
2 101581 1 42381
2 101582 1 42381
2 101583 1 42381
2 101584 1 42382
2 101585 1 42382
2 101586 1 42382
2 101587 1 42385
2 101588 1 42385
2 101589 1 42385
2 101590 1 42385
2 101591 1 42386
2 101592 1 42386
2 101593 1 42393
2 101594 1 42393
2 101595 1 42394
2 101596 1 42394
2 101597 1 42414
2 101598 1 42414
2 101599 1 42440
2 101600 1 42440
2 101601 1 42440
2 101602 1 42441
2 101603 1 42441
2 101604 1 42441
2 101605 1 42441
2 101606 1 42441
2 101607 1 42441
2 101608 1 42441
2 101609 1 42441
2 101610 1 42441
2 101611 1 42441
2 101612 1 42447
2 101613 1 42447
2 101614 1 42447
2 101615 1 42450
2 101616 1 42450
2 101617 1 42451
2 101618 1 42451
2 101619 1 42452
2 101620 1 42452
2 101621 1 42464
2 101622 1 42464
2 101623 1 42464
2 101624 1 42467
2 101625 1 42467
2 101626 1 42474
2 101627 1 42474
2 101628 1 42482
2 101629 1 42482
2 101630 1 42482
2 101631 1 42483
2 101632 1 42483
2 101633 1 42484
2 101634 1 42484
2 101635 1 42484
2 101636 1 42487
2 101637 1 42487
2 101638 1 42490
2 101639 1 42490
2 101640 1 42491
2 101641 1 42491
2 101642 1 42493
2 101643 1 42493
2 101644 1 42528
2 101645 1 42528
2 101646 1 42528
2 101647 1 42539
2 101648 1 42539
2 101649 1 42544
2 101650 1 42544
2 101651 1 42544
2 101652 1 42544
2 101653 1 42544
2 101654 1 42544
2 101655 1 42545
2 101656 1 42545
2 101657 1 42552
2 101658 1 42552
2 101659 1 42552
2 101660 1 42556
2 101661 1 42556
2 101662 1 42566
2 101663 1 42566
2 101664 1 42580
2 101665 1 42580
2 101666 1 42585
2 101667 1 42585
2 101668 1 42585
2 101669 1 42585
2 101670 1 42585
2 101671 1 42598
2 101672 1 42598
2 101673 1 42598
2 101674 1 42599
2 101675 1 42599
2 101676 1 42600
2 101677 1 42600
2 101678 1 42611
2 101679 1 42611
2 101680 1 42624
2 101681 1 42624
2 101682 1 42658
2 101683 1 42658
2 101684 1 42658
2 101685 1 42659
2 101686 1 42659
2 101687 1 42687
2 101688 1 42687
2 101689 1 42687
2 101690 1 42687
2 101691 1 42698
2 101692 1 42698
2 101693 1 42708
2 101694 1 42708
2 101695 1 42708
2 101696 1 42708
2 101697 1 42708
2 101698 1 42708
2 101699 1 42708
2 101700 1 42709
2 101701 1 42709
2 101702 1 42709
2 101703 1 42724
2 101704 1 42724
2 101705 1 42744
2 101706 1 42744
2 101707 1 42744
2 101708 1 42754
2 101709 1 42754
2 101710 1 42766
2 101711 1 42766
2 101712 1 42767
2 101713 1 42767
2 101714 1 42785
2 101715 1 42785
2 101716 1 42785
2 101717 1 42786
2 101718 1 42786
2 101719 1 42790
2 101720 1 42790
2 101721 1 42798
2 101722 1 42798
2 101723 1 42799
2 101724 1 42799
2 101725 1 42807
2 101726 1 42807
2 101727 1 42841
2 101728 1 42841
2 101729 1 42849
2 101730 1 42849
2 101731 1 42849
2 101732 1 42855
2 101733 1 42855
2 101734 1 42903
2 101735 1 42903
2 101736 1 42911
2 101737 1 42911
2 101738 1 43036
2 101739 1 43036
2 101740 1 43037
2 101741 1 43037
2 101742 1 43037
2 101743 1 43042
2 101744 1 43042
2 101745 1 43048
2 101746 1 43048
2 101747 1 43056
2 101748 1 43056
2 101749 1 43056
2 101750 1 43075
2 101751 1 43075
2 101752 1 43078
2 101753 1 43078
2 101754 1 43084
2 101755 1 43084
2 101756 1 43087
2 101757 1 43087
2 101758 1 43088
2 101759 1 43088
2 101760 1 43107
2 101761 1 43107
2 101762 1 43107
2 101763 1 43120
2 101764 1 43120
2 101765 1 43133
2 101766 1 43133
2 101767 1 43144
2 101768 1 43144
2 101769 1 43145
2 101770 1 43145
2 101771 1 43156
2 101772 1 43156
2 101773 1 43156
2 101774 1 43157
2 101775 1 43157
2 101776 1 43177
2 101777 1 43177
2 101778 1 43177
2 101779 1 43186
2 101780 1 43186
2 101781 1 43186
2 101782 1 43211
2 101783 1 43211
2 101784 1 43236
2 101785 1 43236
2 101786 1 43269
2 101787 1 43269
2 101788 1 43269
2 101789 1 43282
2 101790 1 43282
2 101791 1 43282
2 101792 1 43282
2 101793 1 43283
2 101794 1 43283
2 101795 1 43285
2 101796 1 43285
2 101797 1 43285
2 101798 1 43285
2 101799 1 43285
2 101800 1 43286
2 101801 1 43286
2 101802 1 43295
2 101803 1 43295
2 101804 1 43297
2 101805 1 43297
2 101806 1 43299
2 101807 1 43299
2 101808 1 43299
2 101809 1 43302
2 101810 1 43302
2 101811 1 43316
2 101812 1 43316
2 101813 1 43316
2 101814 1 43316
2 101815 1 43317
2 101816 1 43317
2 101817 1 43317
2 101818 1 43317
2 101819 1 43317
2 101820 1 43328
2 101821 1 43328
2 101822 1 43329
2 101823 1 43329
2 101824 1 43352
2 101825 1 43352
2 101826 1 43411
2 101827 1 43411
2 101828 1 43427
2 101829 1 43427
2 101830 1 43440
2 101831 1 43440
2 101832 1 43455
2 101833 1 43455
2 101834 1 43455
2 101835 1 43455
2 101836 1 43455
2 101837 1 43455
2 101838 1 43456
2 101839 1 43456
2 101840 1 43456
2 101841 1 43459
2 101842 1 43459
2 101843 1 43459
2 101844 1 43459
2 101845 1 43459
2 101846 1 43459
2 101847 1 43459
2 101848 1 43462
2 101849 1 43462
2 101850 1 43479
2 101851 1 43479
2 101852 1 43499
2 101853 1 43499
2 101854 1 43521
2 101855 1 43521
2 101856 1 43521
2 101857 1 43521
2 101858 1 43537
2 101859 1 43537
2 101860 1 43537
2 101861 1 43546
2 101862 1 43546
2 101863 1 43546
2 101864 1 43546
2 101865 1 43562
2 101866 1 43562
2 101867 1 43574
2 101868 1 43574
2 101869 1 43574
2 101870 1 43577
2 101871 1 43577
2 101872 1 43577
2 101873 1 43602
2 101874 1 43602
2 101875 1 43602
2 101876 1 43602
2 101877 1 43651
2 101878 1 43651
2 101879 1 43651
2 101880 1 43652
2 101881 1 43652
2 101882 1 43660
2 101883 1 43660
2 101884 1 43670
2 101885 1 43670
2 101886 1 43677
2 101887 1 43677
2 101888 1 43677
2 101889 1 43678
2 101890 1 43678
2 101891 1 43693
2 101892 1 43693
2 101893 1 43693
2 101894 1 43710
2 101895 1 43710
2 101896 1 43718
2 101897 1 43718
2 101898 1 43721
2 101899 1 43721
2 101900 1 43723
2 101901 1 43723
2 101902 1 43724
2 101903 1 43724
2 101904 1 43769
2 101905 1 43769
2 101906 1 43773
2 101907 1 43773
2 101908 1 43773
2 101909 1 43779
2 101910 1 43779
2 101911 1 43779
2 101912 1 43790
2 101913 1 43790
2 101914 1 43790
2 101915 1 43790
2 101916 1 43793
2 101917 1 43793
2 101918 1 43820
2 101919 1 43820
2 101920 1 43820
2 101921 1 43822
2 101922 1 43822
2 101923 1 43830
2 101924 1 43830
2 101925 1 43837
2 101926 1 43837
2 101927 1 43837
2 101928 1 43837
2 101929 1 43837
2 101930 1 43850
2 101931 1 43850
2 101932 1 43850
2 101933 1 43850
2 101934 1 43879
2 101935 1 43879
2 101936 1 43879
2 101937 1 43880
2 101938 1 43880
2 101939 1 43894
2 101940 1 43894
2 101941 1 43917
2 101942 1 43917
2 101943 1 43925
2 101944 1 43925
2 101945 1 44013
2 101946 1 44013
2 101947 1 44013
2 101948 1 44013
2 101949 1 44013
2 101950 1 44013
2 101951 1 44013
2 101952 1 44013
2 101953 1 44022
2 101954 1 44022
2 101955 1 44040
2 101956 1 44040
2 101957 1 44045
2 101958 1 44045
2 101959 1 44048
2 101960 1 44048
2 101961 1 44048
2 101962 1 44051
2 101963 1 44051
2 101964 1 44051
2 101965 1 44051
2 101966 1 44057
2 101967 1 44057
2 101968 1 44064
2 101969 1 44064
2 101970 1 44078
2 101971 1 44078
2 101972 1 44086
2 101973 1 44086
2 101974 1 44099
2 101975 1 44099
2 101976 1 44100
2 101977 1 44100
2 101978 1 44136
2 101979 1 44136
2 101980 1 44136
2 101981 1 44142
2 101982 1 44142
2 101983 1 44172
2 101984 1 44172
2 101985 1 44183
2 101986 1 44183
2 101987 1 44183
2 101988 1 44203
2 101989 1 44203
2 101990 1 44237
2 101991 1 44237
2 101992 1 44239
2 101993 1 44239
2 101994 1 44279
2 101995 1 44279
2 101996 1 44325
2 101997 1 44325
2 101998 1 44350
2 101999 1 44350
2 102000 1 44350
2 102001 1 44362
2 102002 1 44362
2 102003 1 44365
2 102004 1 44365
2 102005 1 44372
2 102006 1 44372
2 102007 1 44384
2 102008 1 44384
2 102009 1 44384
2 102010 1 44386
2 102011 1 44386
2 102012 1 44397
2 102013 1 44397
2 102014 1 44412
2 102015 1 44412
2 102016 1 44414
2 102017 1 44414
2 102018 1 44418
2 102019 1 44418
2 102020 1 44418
2 102021 1 44418
2 102022 1 44418
2 102023 1 44420
2 102024 1 44420
2 102025 1 44426
2 102026 1 44426
2 102027 1 44427
2 102028 1 44427
2 102029 1 44427
2 102030 1 44427
2 102031 1 44448
2 102032 1 44448
2 102033 1 44448
2 102034 1 44449
2 102035 1 44449
2 102036 1 44521
2 102037 1 44521
2 102038 1 44528
2 102039 1 44528
2 102040 1 44614
2 102041 1 44614
2 102042 1 44636
2 102043 1 44636
2 102044 1 44659
2 102045 1 44659
2 102046 1 44659
2 102047 1 44660
2 102048 1 44660
2 102049 1 44681
2 102050 1 44681
2 102051 1 44699
2 102052 1 44699
2 102053 1 44700
2 102054 1 44700
2 102055 1 44702
2 102056 1 44702
2 102057 1 44757
2 102058 1 44757
2 102059 1 44788
2 102060 1 44788
2 102061 1 44842
2 102062 1 44842
2 102063 1 44856
2 102064 1 44856
2 102065 1 44908
2 102066 1 44908
2 102067 1 44928
2 102068 1 44928
2 102069 1 44931
2 102070 1 44931
2 102071 1 44931
2 102072 1 44976
2 102073 1 44976
2 102074 1 44976
2 102075 1 44976
2 102076 1 44979
2 102077 1 44979
2 102078 1 44983
2 102079 1 44983
2 102080 1 45006
2 102081 1 45006
2 102082 1 45006
2 102083 1 45006
2 102084 1 45037
2 102085 1 45037
2 102086 1 45037
2 102087 1 45037
2 102088 1 45058
2 102089 1 45058
2 102090 1 45058
2 102091 1 45089
2 102092 1 45089
2 102093 1 45094
2 102094 1 45094
2 102095 1 45095
2 102096 1 45095
2 102097 1 45104
2 102098 1 45104
2 102099 1 45126
2 102100 1 45126
2 102101 1 45134
2 102102 1 45134
2 102103 1 45135
2 102104 1 45135
2 102105 1 45135
2 102106 1 45135
2 102107 1 45161
2 102108 1 45161
2 102109 1 45188
2 102110 1 45188
2 102111 1 45227
2 102112 1 45227
2 102113 1 45248
2 102114 1 45248
2 102115 1 45248
2 102116 1 45255
2 102117 1 45255
2 102118 1 45308
2 102119 1 45308
2 102120 1 45392
2 102121 1 45392
2 102122 1 45393
2 102123 1 45393
2 102124 1 45396
2 102125 1 45396
2 102126 1 45412
2 102127 1 45412
2 102128 1 45438
2 102129 1 45438
2 102130 1 45440
2 102131 1 45440
2 102132 1 45450
2 102133 1 45450
2 102134 1 45482
2 102135 1 45482
2 102136 1 45499
2 102137 1 45499
2 102138 1 45519
2 102139 1 45519
2 102140 1 45521
2 102141 1 45521
2 102142 1 45521
2 102143 1 45531
2 102144 1 45531
2 102145 1 45532
2 102146 1 45532
2 102147 1 45558
2 102148 1 45558
2 102149 1 45560
2 102150 1 45560
2 102151 1 45574
2 102152 1 45574
2 102153 1 45574
2 102154 1 45575
2 102155 1 45575
2 102156 1 45588
2 102157 1 45588
2 102158 1 45607
2 102159 1 45607
2 102160 1 45615
2 102161 1 45615
2 102162 1 45621
2 102163 1 45621
2 102164 1 45621
2 102165 1 45659
2 102166 1 45659
2 102167 1 45699
2 102168 1 45699
2 102169 1 45710
2 102170 1 45710
2 102171 1 45711
2 102172 1 45711
2 102173 1 45713
2 102174 1 45713
2 102175 1 45731
2 102176 1 45731
2 102177 1 45753
2 102178 1 45753
2 102179 1 45784
2 102180 1 45784
2 102181 1 45789
2 102182 1 45789
2 102183 1 45806
2 102184 1 45806
2 102185 1 45807
2 102186 1 45807
2 102187 1 45823
2 102188 1 45823
2 102189 1 45823
2 102190 1 45823
2 102191 1 45823
2 102192 1 45823
2 102193 1 45852
2 102194 1 45852
2 102195 1 45856
2 102196 1 45856
2 102197 1 45856
2 102198 1 45856
2 102199 1 45870
2 102200 1 45870
2 102201 1 45870
2 102202 1 45870
2 102203 1 45870
2 102204 1 45870
2 102205 1 45870
2 102206 1 45870
2 102207 1 45870
2 102208 1 45870
2 102209 1 45870
2 102210 1 45884
2 102211 1 45884
2 102212 1 45884
2 102213 1 45884
2 102214 1 45893
2 102215 1 45893
2 102216 1 45893
2 102217 1 45893
2 102218 1 45940
2 102219 1 45940
2 102220 1 45948
2 102221 1 45948
2 102222 1 45960
2 102223 1 45960
2 102224 1 45961
2 102225 1 45961
2 102226 1 45966
2 102227 1 45966
2 102228 1 45977
2 102229 1 45977
2 102230 1 45977
2 102231 1 45977
2 102232 1 45977
2 102233 1 45977
2 102234 1 45978
2 102235 1 45978
2 102236 1 45980
2 102237 1 45980
2 102238 1 45981
2 102239 1 45981
2 102240 1 45988
2 102241 1 45988
2 102242 1 46014
2 102243 1 46014
2 102244 1 46014
2 102245 1 46014
2 102246 1 46014
2 102247 1 46015
2 102248 1 46015
2 102249 1 46063
2 102250 1 46063
2 102251 1 46074
2 102252 1 46074
2 102253 1 46082
2 102254 1 46082
2 102255 1 46088
2 102256 1 46088
2 102257 1 46100
2 102258 1 46100
2 102259 1 46100
2 102260 1 46100
2 102261 1 46100
2 102262 1 46100
2 102263 1 46108
2 102264 1 46108
2 102265 1 46108
2 102266 1 46112
2 102267 1 46112
2 102268 1 46112
2 102269 1 46115
2 102270 1 46115
2 102271 1 46115
2 102272 1 46140
2 102273 1 46140
2 102274 1 46154
2 102275 1 46154
2 102276 1 46155
2 102277 1 46155
2 102278 1 46156
2 102279 1 46156
2 102280 1 46156
2 102281 1 46159
2 102282 1 46159
2 102283 1 46159
2 102284 1 46159
2 102285 1 46159
2 102286 1 46159
2 102287 1 46159
2 102288 1 46159
2 102289 1 46159
2 102290 1 46159
2 102291 1 46160
2 102292 1 46160
2 102293 1 46163
2 102294 1 46163
2 102295 1 46163
2 102296 1 46185
2 102297 1 46185
2 102298 1 46185
2 102299 1 46186
2 102300 1 46186
2 102301 1 46186
2 102302 1 46192
2 102303 1 46192
2 102304 1 46201
2 102305 1 46201
2 102306 1 46201
2 102307 1 46201
2 102308 1 46201
2 102309 1 46201
2 102310 1 46211
2 102311 1 46211
2 102312 1 46222
2 102313 1 46222
2 102314 1 46222
2 102315 1 46230
2 102316 1 46230
2 102317 1 46230
2 102318 1 46230
2 102319 1 46268
2 102320 1 46268
2 102321 1 46268
2 102322 1 46269
2 102323 1 46269
2 102324 1 46301
2 102325 1 46301
2 102326 1 46301
2 102327 1 46310
2 102328 1 46310
2 102329 1 46310
2 102330 1 46323
2 102331 1 46323
2 102332 1 46348
2 102333 1 46348
2 102334 1 46357
2 102335 1 46357
2 102336 1 46390
2 102337 1 46390
2 102338 1 46391
2 102339 1 46391
2 102340 1 46427
2 102341 1 46427
2 102342 1 46439
2 102343 1 46439
2 102344 1 46483
2 102345 1 46483
2 102346 1 46634
2 102347 1 46634
2 102348 1 46651
2 102349 1 46651
2 102350 1 46663
2 102351 1 46663
2 102352 1 46674
2 102353 1 46674
2 102354 1 46674
2 102355 1 46713
2 102356 1 46713
2 102357 1 46722
2 102358 1 46722
2 102359 1 46742
2 102360 1 46742
2 102361 1 46743
2 102362 1 46743
2 102363 1 46743
2 102364 1 46743
2 102365 1 46757
2 102366 1 46757
2 102367 1 46773
2 102368 1 46773
2 102369 1 46806
2 102370 1 46806
2 102371 1 46806
2 102372 1 46806
2 102373 1 46820
2 102374 1 46820
2 102375 1 46826
2 102376 1 46826
2 102377 1 46826
2 102378 1 46826
2 102379 1 46845
2 102380 1 46845
2 102381 1 46854
2 102382 1 46854
2 102383 1 46854
2 102384 1 46854
2 102385 1 46871
2 102386 1 46871
2 102387 1 46884
2 102388 1 46884
2 102389 1 46884
2 102390 1 46885
2 102391 1 46885
2 102392 1 46885
2 102393 1 46928
2 102394 1 46928
2 102395 1 46967
2 102396 1 46967
2 102397 1 46976
2 102398 1 46976
2 102399 1 46976
2 102400 1 46978
2 102401 1 46978
2 102402 1 46980
2 102403 1 46980
2 102404 1 46980
2 102405 1 46998
2 102406 1 46998
2 102407 1 46998
2 102408 1 46998
2 102409 1 47003
2 102410 1 47003
2 102411 1 47023
2 102412 1 47023
2 102413 1 47033
2 102414 1 47033
2 102415 1 47052
2 102416 1 47052
2 102417 1 47072
2 102418 1 47072
2 102419 1 47098
2 102420 1 47098
2 102421 1 47105
2 102422 1 47105
2 102423 1 47117
2 102424 1 47117
2 102425 1 47126
2 102426 1 47126
2 102427 1 47160
2 102428 1 47160
2 102429 1 47194
2 102430 1 47194
2 102431 1 47204
2 102432 1 47204
2 102433 1 47219
2 102434 1 47219
2 102435 1 47221
2 102436 1 47221
2 102437 1 47229
2 102438 1 47229
2 102439 1 47264
2 102440 1 47264
2 102441 1 47291
2 102442 1 47291
2 102443 1 47304
2 102444 1 47304
2 102445 1 47324
2 102446 1 47324
2 102447 1 47324
2 102448 1 47378
2 102449 1 47378
2 102450 1 47386
2 102451 1 47386
2 102452 1 47415
2 102453 1 47415
2 102454 1 47422
2 102455 1 47422
2 102456 1 47423
2 102457 1 47423
2 102458 1 47430
2 102459 1 47430
2 102460 1 47460
2 102461 1 47460
2 102462 1 47472
2 102463 1 47472
2 102464 1 47478
2 102465 1 47478
2 102466 1 47480
2 102467 1 47480
2 102468 1 47486
2 102469 1 47486
2 102470 1 47526
2 102471 1 47526
2 102472 1 47526
2 102473 1 47534
2 102474 1 47534
2 102475 1 47537
2 102476 1 47537
2 102477 1 47537
2 102478 1 47538
2 102479 1 47538
2 102480 1 47538
2 102481 1 47538
2 102482 1 47546
2 102483 1 47546
2 102484 1 47548
2 102485 1 47548
2 102486 1 47560
2 102487 1 47560
2 102488 1 47580
2 102489 1 47580
2 102490 1 47625
2 102491 1 47625
2 102492 1 47643
2 102493 1 47643
2 102494 1 47652
2 102495 1 47652
2 102496 1 47663
2 102497 1 47663
2 102498 1 47694
2 102499 1 47694
2 102500 1 47726
2 102501 1 47726
2 102502 1 47729
2 102503 1 47729
2 102504 1 47747
2 102505 1 47747
2 102506 1 47757
2 102507 1 47757
2 102508 1 47762
2 102509 1 47762
2 102510 1 47763
2 102511 1 47763
2 102512 1 47768
2 102513 1 47768
2 102514 1 47782
2 102515 1 47782
2 102516 1 47786
2 102517 1 47786
2 102518 1 47799
2 102519 1 47799
2 102520 1 47873
2 102521 1 47873
2 102522 1 47876
2 102523 1 47876
2 102524 1 47884
2 102525 1 47884
2 102526 1 47894
2 102527 1 47894
2 102528 1 47894
2 102529 1 47926
2 102530 1 47926
2 102531 1 47997
2 102532 1 47997
2 102533 1 48005
2 102534 1 48005
2 102535 1 48006
2 102536 1 48006
2 102537 1 48006
2 102538 1 48009
2 102539 1 48009
2 102540 1 48017
2 102541 1 48017
2 102542 1 48140
2 102543 1 48140
2 102544 1 48145
2 102545 1 48145
2 102546 1 48238
2 102547 1 48238
2 102548 1 48242
2 102549 1 48242
2 102550 1 48244
2 102551 1 48244
2 102552 1 48260
2 102553 1 48260
2 102554 1 48260
2 102555 1 48283
2 102556 1 48283
2 102557 1 48287
2 102558 1 48287
2 102559 1 48288
2 102560 1 48288
2 102561 1 48296
2 102562 1 48296
2 102563 1 48296
2 102564 1 48303
2 102565 1 48303
2 102566 1 48307
2 102567 1 48307
2 102568 1 48316
2 102569 1 48316
2 102570 1 48316
2 102571 1 48323
2 102572 1 48323
2 102573 1 48329
2 102574 1 48329
2 102575 1 48358
2 102576 1 48358
2 102577 1 48358
2 102578 1 48365
2 102579 1 48365
2 102580 1 48368
2 102581 1 48368
2 102582 1 48369
2 102583 1 48369
2 102584 1 48386
2 102585 1 48386
2 102586 1 48397
2 102587 1 48397
2 102588 1 48397
2 102589 1 48397
2 102590 1 48400
2 102591 1 48400
2 102592 1 48425
2 102593 1 48425
2 102594 1 48426
2 102595 1 48426
2 102596 1 48434
2 102597 1 48434
2 102598 1 48434
2 102599 1 48434
2 102600 1 48435
2 102601 1 48435
2 102602 1 48454
2 102603 1 48454
2 102604 1 48457
2 102605 1 48457
2 102606 1 48465
2 102607 1 48465
2 102608 1 48473
2 102609 1 48473
2 102610 1 48477
2 102611 1 48477
2 102612 1 48477
2 102613 1 48477
2 102614 1 48478
2 102615 1 48478
2 102616 1 48478
2 102617 1 48478
2 102618 1 48481
2 102619 1 48481
2 102620 1 48482
2 102621 1 48482
2 102622 1 48520
2 102623 1 48520
2 102624 1 48520
2 102625 1 48561
2 102626 1 48561
2 102627 1 48564
2 102628 1 48564
2 102629 1 48569
2 102630 1 48569
2 102631 1 48569
2 102632 1 48573
2 102633 1 48573
2 102634 1 48573
2 102635 1 48573
2 102636 1 48573
2 102637 1 48573
2 102638 1 48573
2 102639 1 48596
2 102640 1 48596
2 102641 1 48633
2 102642 1 48633
2 102643 1 48679
2 102644 1 48679
2 102645 1 48696
2 102646 1 48696
2 102647 1 48696
2 102648 1 48696
2 102649 1 48704
2 102650 1 48704
2 102651 1 48704
2 102652 1 48705
2 102653 1 48705
2 102654 1 48712
2 102655 1 48712
2 102656 1 48712
2 102657 1 48733
2 102658 1 48733
2 102659 1 48733
2 102660 1 48738
2 102661 1 48738
2 102662 1 48752
2 102663 1 48752
2 102664 1 48752
2 102665 1 48752
2 102666 1 48772
2 102667 1 48772
2 102668 1 48772
2 102669 1 48799
2 102670 1 48799
2 102671 1 48819
2 102672 1 48819
2 102673 1 48851
2 102674 1 48851
2 102675 1 48855
2 102676 1 48855
2 102677 1 48855
2 102678 1 48855
2 102679 1 48855
2 102680 1 48855
2 102681 1 48856
2 102682 1 48856
2 102683 1 48857
2 102684 1 48857
2 102685 1 48862
2 102686 1 48862
2 102687 1 48862
2 102688 1 48862
2 102689 1 48862
2 102690 1 48862
2 102691 1 48865
2 102692 1 48865
2 102693 1 48896
2 102694 1 48896
2 102695 1 48928
2 102696 1 48928
2 102697 1 48947
2 102698 1 48947
2 102699 1 48947
2 102700 1 48953
2 102701 1 48953
2 102702 1 48956
2 102703 1 48956
2 102704 1 48956
2 102705 1 48969
2 102706 1 48969
2 102707 1 48982
2 102708 1 48982
2 102709 1 49001
2 102710 1 49001
2 102711 1 49020
2 102712 1 49020
2 102713 1 49028
2 102714 1 49028
2 102715 1 49031
2 102716 1 49031
2 102717 1 49033
2 102718 1 49033
2 102719 1 49038
2 102720 1 49038
2 102721 1 49067
2 102722 1 49067
2 102723 1 49084
2 102724 1 49084
2 102725 1 49109
2 102726 1 49109
2 102727 1 49144
2 102728 1 49144
2 102729 1 49157
2 102730 1 49157
2 102731 1 49166
2 102732 1 49166
2 102733 1 49173
2 102734 1 49173
2 102735 1 49199
2 102736 1 49199
2 102737 1 49199
2 102738 1 49204
2 102739 1 49204
2 102740 1 49211
2 102741 1 49211
2 102742 1 49211
2 102743 1 49225
2 102744 1 49225
2 102745 1 49232
2 102746 1 49232
2 102747 1 49250
2 102748 1 49250
2 102749 1 49279
2 102750 1 49279
2 102751 1 49281
2 102752 1 49281
2 102753 1 49310
2 102754 1 49310
2 102755 1 49310
2 102756 1 49329
2 102757 1 49329
2 102758 1 49329
2 102759 1 49329
2 102760 1 49329
2 102761 1 49329
2 102762 1 49329
2 102763 1 49329
2 102764 1 49329
2 102765 1 49332
2 102766 1 49332
2 102767 1 49332
2 102768 1 49342
2 102769 1 49342
2 102770 1 49355
2 102771 1 49355
2 102772 1 49355
2 102773 1 49357
2 102774 1 49357
2 102775 1 49369
2 102776 1 49369
2 102777 1 49434
2 102778 1 49434
2 102779 1 49434
2 102780 1 49435
2 102781 1 49435
2 102782 1 49436
2 102783 1 49436
2 102784 1 49470
2 102785 1 49470
2 102786 1 49497
2 102787 1 49497
2 102788 1 49498
2 102789 1 49498
2 102790 1 49515
2 102791 1 49515
2 102792 1 49519
2 102793 1 49519
2 102794 1 49521
2 102795 1 49521
2 102796 1 49558
2 102797 1 49558
2 102798 1 49567
2 102799 1 49567
2 102800 1 49567
2 102801 1 49580
2 102802 1 49580
2 102803 1 49581
2 102804 1 49581
2 102805 1 49588
2 102806 1 49588
2 102807 1 49653
2 102808 1 49653
2 102809 1 49702
2 102810 1 49702
2 102811 1 49703
2 102812 1 49703
2 102813 1 49703
2 102814 1 49703
2 102815 1 49740
2 102816 1 49740
2 102817 1 49751
2 102818 1 49751
2 102819 1 49751
2 102820 1 49751
2 102821 1 49772
2 102822 1 49772
2 102823 1 49772
2 102824 1 49772
2 102825 1 49772
2 102826 1 49772
2 102827 1 49788
2 102828 1 49788
2 102829 1 49788
2 102830 1 49789
2 102831 1 49789
2 102832 1 49789
2 102833 1 49789
2 102834 1 49789
2 102835 1 49789
2 102836 1 49803
2 102837 1 49803
2 102838 1 49818
2 102839 1 49818
2 102840 1 49818
2 102841 1 49818
2 102842 1 49833
2 102843 1 49833
2 102844 1 49833
2 102845 1 49864
2 102846 1 49864
2 102847 1 49878
2 102848 1 49878
2 102849 1 49896
2 102850 1 49896
2 102851 1 49896
2 102852 1 49897
2 102853 1 49897
2 102854 1 49919
2 102855 1 49919
2 102856 1 49930
2 102857 1 49930
2 102858 1 49975
2 102859 1 49975
2 102860 1 49975
2 102861 1 49983
2 102862 1 49983
2 102863 1 49995
2 102864 1 49995
2 102865 1 50060
2 102866 1 50060
2 102867 1 50064
2 102868 1 50064
2 102869 1 50083
2 102870 1 50083
2 102871 1 50097
2 102872 1 50097
2 102873 1 50103
2 102874 1 50103
2 102875 1 50105
2 102876 1 50105
2 102877 1 50126
2 102878 1 50126
2 102879 1 50127
2 102880 1 50127
2 102881 1 50144
2 102882 1 50144
2 102883 1 50149
2 102884 1 50149
2 102885 1 50169
2 102886 1 50169
2 102887 1 50177
2 102888 1 50177
2 102889 1 50179
2 102890 1 50179
2 102891 1 50179
2 102892 1 50180
2 102893 1 50180
2 102894 1 50235
2 102895 1 50235
2 102896 1 50238
2 102897 1 50238
2 102898 1 50238
2 102899 1 50238
2 102900 1 50238
2 102901 1 50361
2 102902 1 50361
2 102903 1 50373
2 102904 1 50373
2 102905 1 50381
2 102906 1 50381
2 102907 1 50393
2 102908 1 50393
2 102909 1 50425
2 102910 1 50425
2 102911 1 50559
2 102912 1 50559
2 102913 1 50566
2 102914 1 50566
2 102915 1 50574
2 102916 1 50574
2 102917 1 50581
2 102918 1 50581
2 102919 1 50613
2 102920 1 50613
2 102921 1 50634
2 102922 1 50634
2 102923 1 50649
2 102924 1 50649
2 102925 1 50652
2 102926 1 50652
2 102927 1 50675
2 102928 1 50675
2 102929 1 50678
2 102930 1 50678
2 102931 1 50678
2 102932 1 50678
2 102933 1 50685
2 102934 1 50685
2 102935 1 50685
2 102936 1 50698
2 102937 1 50698
2 102938 1 50839
2 102939 1 50839
2 102940 1 50992
2 102941 1 50992
2 102942 1 51031
2 102943 1 51031
2 102944 1 51125
2 102945 1 51125
2 102946 1 51126
2 102947 1 51126
2 102948 1 51127
2 102949 1 51127
2 102950 1 51130
2 102951 1 51130
2 102952 1 51159
2 102953 1 51159
2 102954 1 51159
2 102955 1 51159
2 102956 1 51159
2 102957 1 51164
2 102958 1 51164
2 102959 1 51165
2 102960 1 51165
2 102961 1 51167
2 102962 1 51167
2 102963 1 51167
2 102964 1 51167
2 102965 1 51169
2 102966 1 51169
2 102967 1 51213
2 102968 1 51213
2 102969 1 51261
2 102970 1 51261
2 102971 1 51263
2 102972 1 51263
2 102973 1 51296
2 102974 1 51296
2 102975 1 51332
2 102976 1 51332
2 102977 1 51334
2 102978 1 51334
2 102979 1 51343
2 102980 1 51343
2 102981 1 51343
2 102982 1 51343
2 102983 1 51352
2 102984 1 51352
2 102985 1 51353
2 102986 1 51353
2 102987 1 51360
2 102988 1 51360
2 102989 1 51373
2 102990 1 51373
2 102991 1 51374
2 102992 1 51374
2 102993 1 51374
2 102994 1 51374
2 102995 1 51374
2 102996 1 51427
2 102997 1 51427
2 102998 1 51427
2 102999 1 51428
2 103000 1 51428
2 103001 1 51436
2 103002 1 51436
2 103003 1 51437
2 103004 1 51437
2 103005 1 51470
2 103006 1 51470
2 103007 1 51470
2 103008 1 51470
2 103009 1 51470
2 103010 1 51470
2 103011 1 51472
2 103012 1 51472
2 103013 1 51484
2 103014 1 51484
2 103015 1 51484
2 103016 1 51494
2 103017 1 51494
2 103018 1 51494
2 103019 1 51495
2 103020 1 51495
2 103021 1 51511
2 103022 1 51511
2 103023 1 51511
2 103024 1 51529
2 103025 1 51529
2 103026 1 51543
2 103027 1 51543
2 103028 1 51551
2 103029 1 51551
2 103030 1 51553
2 103031 1 51553
2 103032 1 51556
2 103033 1 51556
2 103034 1 51556
2 103035 1 51556
2 103036 1 51559
2 103037 1 51559
2 103038 1 51561
2 103039 1 51561
2 103040 1 51581
2 103041 1 51581
2 103042 1 51595
2 103043 1 51595
2 103044 1 51613
2 103045 1 51613
2 103046 1 51614
2 103047 1 51614
2 103048 1 51614
2 103049 1 51627
2 103050 1 51627
2 103051 1 51627
2 103052 1 51629
2 103053 1 51629
2 103054 1 51643
2 103055 1 51643
2 103056 1 51646
2 103057 1 51646
2 103058 1 51662
2 103059 1 51662
2 103060 1 51665
2 103061 1 51665
2 103062 1 51670
2 103063 1 51670
2 103064 1 51693
2 103065 1 51693
2 103066 1 51693
2 103067 1 51704
2 103068 1 51704
2 103069 1 51715
2 103070 1 51715
2 103071 1 51715
2 103072 1 51720
2 103073 1 51720
2 103074 1 51722
2 103075 1 51722
2 103076 1 51748
2 103077 1 51748
2 103078 1 51751
2 103079 1 51751
2 103080 1 51760
2 103081 1 51760
2 103082 1 51760
2 103083 1 51760
2 103084 1 51760
2 103085 1 51796
2 103086 1 51796
2 103087 1 51796
2 103088 1 51844
2 103089 1 51844
2 103090 1 51859
2 103091 1 51859
2 103092 1 51867
2 103093 1 51867
2 103094 1 51936
2 103095 1 51936
2 103096 1 51937
2 103097 1 51937
2 103098 1 51938
2 103099 1 51938
2 103100 1 51946
2 103101 1 51946
2 103102 1 51968
2 103103 1 51968
2 103104 1 52042
2 103105 1 52042
2 103106 1 52042
2 103107 1 52045
2 103108 1 52045
2 103109 1 52057
2 103110 1 52057
2 103111 1 52057
2 103112 1 52069
2 103113 1 52069
2 103114 1 52071
2 103115 1 52071
2 103116 1 52074
2 103117 1 52074
2 103118 1 52074
2 103119 1 52082
2 103120 1 52082
2 103121 1 52138
2 103122 1 52138
2 103123 1 52196
2 103124 1 52196
2 103125 1 52196
2 103126 1 52198
2 103127 1 52198
2 103128 1 52201
2 103129 1 52201
2 103130 1 52234
2 103131 1 52234
2 103132 1 52239
2 103133 1 52239
2 103134 1 52259
2 103135 1 52259
2 103136 1 52259
2 103137 1 52259
2 103138 1 52259
2 103139 1 52259
2 103140 1 52259
2 103141 1 52259
2 103142 1 52263
2 103143 1 52263
2 103144 1 52263
2 103145 1 52284
2 103146 1 52284
2 103147 1 52299
2 103148 1 52299
2 103149 1 52308
2 103150 1 52308
2 103151 1 52308
2 103152 1 52315
2 103153 1 52315
2 103154 1 52315
2 103155 1 52315
2 103156 1 52369
2 103157 1 52369
2 103158 1 52369
2 103159 1 52371
2 103160 1 52371
2 103161 1 52375
2 103162 1 52375
2 103163 1 52418
2 103164 1 52418
2 103165 1 52438
2 103166 1 52438
2 103167 1 52479
2 103168 1 52479
2 103169 1 52494
2 103170 1 52494
2 103171 1 52494
2 103172 1 52498
2 103173 1 52498
2 103174 1 52498
2 103175 1 52506
2 103176 1 52506
2 103177 1 52506
2 103178 1 52507
2 103179 1 52507
2 103180 1 52509
2 103181 1 52509
2 103182 1 52517
2 103183 1 52517
2 103184 1 52531
2 103185 1 52531
2 103186 1 52531
2 103187 1 52547
2 103188 1 52547
2 103189 1 52575
2 103190 1 52575
2 103191 1 52577
2 103192 1 52577
2 103193 1 52581
2 103194 1 52581
2 103195 1 52581
2 103196 1 52588
2 103197 1 52588
2 103198 1 52603
2 103199 1 52603
2 103200 1 52603
2 103201 1 52603
2 103202 1 52603
2 103203 1 52604
2 103204 1 52604
2 103205 1 52629
2 103206 1 52629
2 103207 1 52640
2 103208 1 52640
2 103209 1 52653
2 103210 1 52653
2 103211 1 52660
2 103212 1 52660
2 103213 1 52674
2 103214 1 52674
2 103215 1 52689
2 103216 1 52689
2 103217 1 52689
2 103218 1 52689
2 103219 1 52689
2 103220 1 52731
2 103221 1 52731
2 103222 1 52780
2 103223 1 52780
2 103224 1 52780
2 103225 1 52780
2 103226 1 52780
2 103227 1 52783
2 103228 1 52783
2 103229 1 52783
2 103230 1 52791
2 103231 1 52791
2 103232 1 52791
2 103233 1 52791
2 103234 1 52791
2 103235 1 52791
2 103236 1 52791
2 103237 1 52791
2 103238 1 52791
2 103239 1 52836
2 103240 1 52836
2 103241 1 52843
2 103242 1 52843
2 103243 1 52854
2 103244 1 52854
2 103245 1 52898
2 103246 1 52898
2 103247 1 52898
2 103248 1 52900
2 103249 1 52900
2 103250 1 52916
2 103251 1 52916
2 103252 1 52999
2 103253 1 52999
2 103254 1 52999
2 103255 1 52999
2 103256 1 52999
2 103257 1 53009
2 103258 1 53009
2 103259 1 53040
2 103260 1 53040
2 103261 1 53048
2 103262 1 53048
2 103263 1 53051
2 103264 1 53051
2 103265 1 53121
2 103266 1 53121
2 103267 1 53121
2 103268 1 53135
2 103269 1 53135
2 103270 1 53138
2 103271 1 53138
2 103272 1 53142
2 103273 1 53142
2 103274 1 53160
2 103275 1 53160
2 103276 1 53164
2 103277 1 53164
2 103278 1 53164
2 103279 1 53164
2 103280 1 53204
2 103281 1 53204
2 103282 1 53215
2 103283 1 53215
2 103284 1 53269
2 103285 1 53269
2 103286 1 53289
2 103287 1 53289
2 103288 1 53337
2 103289 1 53337
2 103290 1 53337
2 103291 1 53360
2 103292 1 53360
2 103293 1 53360
2 103294 1 53363
2 103295 1 53363
2 103296 1 53367
2 103297 1 53367
2 103298 1 53370
2 103299 1 53370
2 103300 1 53385
2 103301 1 53385
2 103302 1 53388
2 103303 1 53388
2 103304 1 53390
2 103305 1 53390
2 103306 1 53404
2 103307 1 53404
2 103308 1 53404
2 103309 1 53406
2 103310 1 53406
2 103311 1 53424
2 103312 1 53424
2 103313 1 53424
2 103314 1 53474
2 103315 1 53474
2 103316 1 53476
2 103317 1 53476
2 103318 1 53476
2 103319 1 53478
2 103320 1 53478
2 103321 1 53504
2 103322 1 53504
2 103323 1 53505
2 103324 1 53505
2 103325 1 53505
2 103326 1 53509
2 103327 1 53509
2 103328 1 53514
2 103329 1 53514
2 103330 1 53521
2 103331 1 53521
2 103332 1 53521
2 103333 1 53536
2 103334 1 53536
2 103335 1 53536
2 103336 1 53551
2 103337 1 53551
2 103338 1 53553
2 103339 1 53553
2 103340 1 53555
2 103341 1 53555
2 103342 1 53592
2 103343 1 53592
2 103344 1 53603
2 103345 1 53603
2 103346 1 53623
2 103347 1 53623
2 103348 1 53623
2 103349 1 53648
2 103350 1 53648
2 103351 1 53716
2 103352 1 53716
2 103353 1 53744
2 103354 1 53744
2 103355 1 53756
2 103356 1 53756
2 103357 1 53782
2 103358 1 53782
2 103359 1 53815
2 103360 1 53815
2 103361 1 53815
2 103362 1 53846
2 103363 1 53846
2 103364 1 53858
2 103365 1 53858
2 103366 1 53912
2 103367 1 53912
2 103368 1 53945
2 103369 1 53945
2 103370 1 53945
2 103371 1 53947
2 103372 1 53947
2 103373 1 53947
2 103374 1 53983
2 103375 1 53983
2 103376 1 54014
2 103377 1 54014
2 103378 1 54076
2 103379 1 54076
2 103380 1 54132
2 103381 1 54132
2 103382 1 54132
2 103383 1 54171
2 103384 1 54171
2 103385 1 54197
2 103386 1 54197
2 103387 1 54261
2 103388 1 54261
2 103389 1 54261
2 103390 1 54375
2 103391 1 54375
2 103392 1 54385
2 103393 1 54385
2 103394 1 54387
2 103395 1 54387
2 103396 1 54389
2 103397 1 54389
2 103398 1 54390
2 103399 1 54390
2 103400 1 54394
2 103401 1 54394
2 103402 1 54433
2 103403 1 54433
2 103404 1 54438
2 103405 1 54438
2 103406 1 54447
2 103407 1 54447
2 103408 1 54457
2 103409 1 54457
2 103410 1 54490
2 103411 1 54490
2 103412 1 54492
2 103413 1 54492
2 103414 1 54492
2 103415 1 54492
2 103416 1 54493
2 103417 1 54493
2 103418 1 54508
2 103419 1 54508
2 103420 1 54518
2 103421 1 54518
2 103422 1 54599
2 103423 1 54599
2 103424 1 54612
2 103425 1 54612
2 103426 1 54634
2 103427 1 54634
2 103428 1 54636
2 103429 1 54636
2 103430 1 54712
2 103431 1 54712
2 103432 1 54712
2 103433 1 54737
2 103434 1 54737
2 103435 1 54752
2 103436 1 54752
2 103437 1 54767
2 103438 1 54767
2 103439 1 54767
2 103440 1 54771
2 103441 1 54771
2 103442 1 54833
2 103443 1 54833
2 103444 1 54849
2 103445 1 54849
2 103446 1 54850
2 103447 1 54850
2 103448 1 54892
2 103449 1 54892
2 103450 1 54905
2 103451 1 54905
2 103452 1 54981
2 103453 1 54981
2 103454 1 55005
2 103455 1 55005
2 103456 1 55030
2 103457 1 55030
2 103458 1 55044
2 103459 1 55044
2 103460 1 55044
2 103461 1 55065
2 103462 1 55065
2 103463 1 55065
2 103464 1 55095
2 103465 1 55095
2 103466 1 55153
2 103467 1 55153
2 103468 1 55153
2 103469 1 55154
2 103470 1 55154
2 103471 1 55154
2 103472 1 55218
2 103473 1 55218
2 103474 1 55228
2 103475 1 55228
2 103476 1 55231
2 103477 1 55231
2 103478 1 55241
2 103479 1 55241
2 103480 1 55249
2 103481 1 55249
2 103482 1 55250
2 103483 1 55250
2 103484 1 55255
2 103485 1 55255
2 103486 1 55255
2 103487 1 55258
2 103488 1 55258
2 103489 1 55258
2 103490 1 55265
2 103491 1 55265
2 103492 1 55266
2 103493 1 55266
2 103494 1 55266
2 103495 1 55266
2 103496 1 55266
2 103497 1 55266
2 103498 1 55266
2 103499 1 55266
2 103500 1 55266
2 103501 1 55266
2 103502 1 55271
2 103503 1 55271
2 103504 1 55271
2 103505 1 55273
2 103506 1 55273
2 103507 1 55289
2 103508 1 55289
2 103509 1 55311
2 103510 1 55311
2 103511 1 55312
2 103512 1 55312
2 103513 1 55313
2 103514 1 55313
2 103515 1 55333
2 103516 1 55333
2 103517 1 55333
2 103518 1 55351
2 103519 1 55351
2 103520 1 55373
2 103521 1 55373
2 103522 1 55390
2 103523 1 55390
2 103524 1 55445
2 103525 1 55445
2 103526 1 55457
2 103527 1 55457
2 103528 1 55531
2 103529 1 55531
2 103530 1 55579
2 103531 1 55579
2 103532 1 55604
2 103533 1 55604
2 103534 1 55611
2 103535 1 55611
2 103536 1 55612
2 103537 1 55612
2 103538 1 55615
2 103539 1 55615
2 103540 1 55618
2 103541 1 55618
2 103542 1 55645
2 103543 1 55645
2 103544 1 55672
2 103545 1 55672
2 103546 1 55687
2 103547 1 55687
2 103548 1 55688
2 103549 1 55688
2 103550 1 55688
2 103551 1 55695
2 103552 1 55695
2 103553 1 55695
2 103554 1 55697
2 103555 1 55697
2 103556 1 55701
2 103557 1 55701
2 103558 1 55708
2 103559 1 55708
2 103560 1 55723
2 103561 1 55723
2 103562 1 55732
2 103563 1 55732
2 103564 1 55745
2 103565 1 55745
2 103566 1 55790
2 103567 1 55790
2 103568 1 55816
2 103569 1 55816
2 103570 1 55825
2 103571 1 55825
2 103572 1 55833
2 103573 1 55833
2 103574 1 55841
2 103575 1 55841
2 103576 1 55862
2 103577 1 55862
2 103578 1 55891
2 103579 1 55891
2 103580 1 55891
2 103581 1 55894
2 103582 1 55894
2 103583 1 55909
2 103584 1 55909
2 103585 1 55921
2 103586 1 55921
2 103587 1 55924
2 103588 1 55924
2 103589 1 55947
2 103590 1 55947
2 103591 1 55957
2 103592 1 55957
2 103593 1 55968
2 103594 1 55968
2 103595 1 55976
2 103596 1 55976
2 103597 1 56038
2 103598 1 56038
2 103599 1 56068
2 103600 1 56068
2 103601 1 56084
2 103602 1 56084
2 103603 1 56122
2 103604 1 56122
2 103605 1 56173
2 103606 1 56173
2 103607 1 56173
2 103608 1 56190
2 103609 1 56190
2 103610 1 56227
2 103611 1 56227
2 103612 1 56346
2 103613 1 56346
2 103614 1 56365
2 103615 1 56365
2 103616 1 56404
2 103617 1 56404
2 103618 1 56577
2 103619 1 56577
2 103620 1 56599
2 103621 1 56599
2 103622 1 56603
2 103623 1 56603
2 103624 1 56611
2 103625 1 56611
2 103626 1 56612
2 103627 1 56612
2 103628 1 56627
2 103629 1 56627
2 103630 1 56638
2 103631 1 56638
2 103632 1 56638
2 103633 1 56642
2 103634 1 56642
2 103635 1 56659
2 103636 1 56659
2 103637 1 56708
2 103638 1 56708
2 103639 1 56708
2 103640 1 56711
2 103641 1 56711
2 103642 1 56736
2 103643 1 56736
2 103644 1 56823
2 103645 1 56823
2 103646 1 56823
2 103647 1 56987
2 103648 1 56987
2 103649 1 56987
2 103650 1 57056
2 103651 1 57056
2 103652 1 57122
2 103653 1 57122
2 103654 1 57122
2 103655 1 57159
2 103656 1 57159
2 103657 1 57168
2 103658 1 57168
2 103659 1 57168
2 103660 1 57191
2 103661 1 57191
2 103662 1 57192
2 103663 1 57192
2 103664 1 57201
2 103665 1 57201
2 103666 1 57295
2 103667 1 57295
2 103668 1 57303
2 103669 1 57303
2 103670 1 57384
2 103671 1 57384
2 103672 1 57416
2 103673 1 57416
2 103674 1 57545
2 103675 1 57545
2 103676 1 57609
2 103677 1 57609
2 103678 1 57680
2 103679 1 57680
2 103680 1 57688
2 103681 1 57688
2 103682 1 57710
2 103683 1 57710
2 103684 1 57710
2 103685 1 57798
2 103686 1 57798
2 103687 1 57829
2 103688 1 57829
2 103689 1 57850
2 103690 1 57850
2 103691 1 57887
2 103692 1 57887
2 103693 1 57918
2 103694 1 57918
2 103695 1 57957
2 103696 1 57957
2 103697 1 57957
2 103698 1 57976
2 103699 1 57976
2 103700 1 57976
2 103701 1 58265
2 103702 1 58265
2 103703 1 58273
2 103704 1 58273
2 103705 1 58273
2 103706 1 58299
2 103707 1 58299
2 103708 1 58334
2 103709 1 58334
2 103710 1 58334
2 103711 1 58404
2 103712 1 58404
2 103713 1 58418
2 103714 1 58418
2 103715 1 58433
2 103716 1 58433
2 103717 1 58479
2 103718 1 58479
2 103719 1 58479
2 103720 1 58487
2 103721 1 58487
2 103722 1 58488
2 103723 1 58488
2 103724 1 58508
2 103725 1 58508
2 103726 1 58525
2 103727 1 58525
2 103728 1 58573
2 103729 1 58573
2 103730 1 58581
2 103731 1 58581
2 103732 1 58590
2 103733 1 58590
2 103734 1 58636
2 103735 1 58636
2 103736 1 58639
2 103737 1 58639
2 103738 1 58664
2 103739 1 58664
2 103740 1 58673
2 103741 1 58673
2 103742 1 58709
2 103743 1 58709
2 103744 1 58744
2 103745 1 58744
2 103746 1 58744
2 103747 1 58760
2 103748 1 58760
2 103749 1 58776
2 103750 1 58776
2 103751 1 58783
2 103752 1 58783
2 103753 1 58788
2 103754 1 58788
2 103755 1 58793
2 103756 1 58793
2 103757 1 58793
2 103758 1 58895
2 103759 1 58895
2 103760 1 58957
2 103761 1 58957
2 103762 1 59046
2 103763 1 59046
2 103764 1 59068
2 103765 1 59068
2 103766 1 59099
2 103767 1 59099
2 103768 1 59100
2 103769 1 59100
2 103770 1 59154
2 103771 1 59154
2 103772 1 59155
2 103773 1 59155
2 103774 1 59190
2 103775 1 59190
2 103776 1 59315
2 103777 1 59315
2 103778 1 59408
2 103779 1 59408
2 103780 1 59539
2 103781 1 59539
2 103782 1 59570
2 103783 1 59570
2 103784 1 59668
2 103785 1 59668
2 103786 1 59720
2 103787 1 59720
2 103788 1 59729
2 103789 1 59729
2 103790 1 59922
2 103791 1 59922
2 103792 1 60003
2 103793 1 60003
2 103794 1 60099
2 103795 1 60099
2 103796 1 60160
2 103797 1 60160
2 103798 1 60163
2 103799 1 60163
2 103800 1 60297
2 103801 1 60297
2 103802 1 60318
2 103803 1 60318
2 103804 1 60380
2 103805 1 60380
2 103806 1 60494
2 103807 1 60494
2 103808 1 60507
2 103809 1 60507
2 103810 1 60563
2 103811 1 60563
2 103812 1 60577
2 103813 1 60577
2 103814 1 60633
2 103815 1 60633
2 103816 1 60679
2 103817 1 60679
2 103818 1 60694
2 103819 1 60694
2 103820 1 60749
2 103821 1 60749
2 103822 1 60833
2 103823 1 60833
2 103824 1 60934
2 103825 1 60934
2 103826 1 60956
2 103827 1 60956
2 103828 1 61060
2 103829 1 61060
2 103830 1 61091
2 103831 1 61091
2 103832 1 61118
2 103833 1 61118
0 27 5 136 1 25
0 28 5 133 1 61341
0 29 5 238 1 61424
0 30 5 223 1 61696
0 31 5 302 1 61940
0 32 5 217 1 62271
0 33 5 229 1 62460
0 34 5 213 1 62695
0 35 5 77 1 62938
0 36 5 72 1 62993
0 37 5 145 1 63045
0 38 5 197 1 63216
0 39 5 246 1 63417
0 40 5 236 1 63656
0 41 5 155 1 63864
0 42 5 196 1 64018
0 43 5 72 1 64240
0 44 5 120 1 64311
0 45 5 184 1 64426
0 46 5 195 1 64609
0 47 5 221 1 64819
0 48 5 306 1 65008
0 49 5 376 1 65264
0 50 5 248 1 65620
0 51 5 179 1 65893
0 52 7 15 2 66576 62461
0 53 7 5 2 68888 69655
0 54 7 2 2 70985 71000
0 55 5 2 1 71005
0 56 7 14 2 67547 68733
0 57 5 5 1 71009
0 58 7 61 2 61697 64820
0 59 5 8 1 71028
0 60 7 2 2 66577 71001
0 61 5 1 1 71097
0 62 7 1 2 71089 61
0 63 5 6 1 62
0 64 7 1 2 71023 71099
0 65 5 1 1 64
0 66 7 1 2 71007 65
0 67 5 1 1 66
0 68 7 1 2 70558 67
0 69 5 1 1 68
0 70 7 12 2 67548 64019
0 71 5 2 1 71105
0 72 7 15 2 62696 68889
0 73 5 2 1 71119
0 74 7 2 2 71117 71134
0 75 5 47 1 71136
0 76 7 92 2 67318 68734
0 77 5 128 1 71185
0 78 7 51 2 66578 69656
0 79 5 2 1 71405
0 80 7 4 2 71277 71406
0 81 7 1 2 71138 71458
0 82 5 1 1 81
0 83 7 1 2 69 82
0 84 5 1 1 83
0 85 7 1 2 68497 84
0 86 5 1 1 85
0 87 7 7 2 67549 69657
0 88 7 3 2 66579 71462
0 89 5 1 1 71469
0 90 7 1 2 71090 89
0 91 5 14 1 90
0 92 7 13 2 62272 68498
0 93 5 10 1 71486
0 94 7 42 2 68735 65621
0 95 5 60 1 71509
0 96 7 4 2 62273 71551
0 97 5 6 1 71611
0 98 7 3 2 63657 71615
0 99 5 2 1 71621
0 100 7 3 2 71499 71624
0 101 5 1 1 71626
0 102 7 10 2 68499 64020
0 103 7 1 2 70559 71629
0 104 5 1 1 103
0 105 7 1 2 71627 104
0 106 5 1 1 105
0 107 7 1 2 71472 106
0 108 5 1 1 107
0 109 7 18 2 68890 65622
0 110 5 5 1 71639
0 111 7 19 2 62462 67550
0 112 5 1 1 71662
0 113 7 2 2 71640 71663
0 114 5 2 1 71681
0 115 7 11 2 69658 65894
0 116 7 6 2 66580 63865
0 117 7 1 2 71685 71696
0 118 7 1 2 71682 117
0 119 5 1 1 118
0 120 7 1 2 108 119
0 121 7 1 2 86 120
0 122 5 1 1 121
0 123 7 1 2 65265 122
0 124 5 1 1 123
0 125 7 5 2 63658 64821
0 126 7 6 2 70806 71278
0 127 5 1 1 71707
0 128 7 40 2 70182 70560
0 129 5 5 1 71713
0 130 7 3 2 64021 71714
0 131 7 3 2 71708 71758
0 132 5 1 1 71761
0 133 7 3 2 71702 71762
0 134 7 20 2 66581 62274
0 135 7 2 2 62697 71767
0 136 7 1 2 71764 71787
0 137 5 1 1 136
0 138 7 1 2 124 137
0 139 5 1 1 138
0 140 7 1 2 61941 139
0 141 5 1 1 140
0 142 7 97 2 62275 63659
0 143 5 110 1 71789
0 144 7 99 2 64022 70807
0 145 5 123 1 71996
0 146 7 14 2 66799 62698
0 147 5 2 1 72218
0 148 7 2 2 71997 72219
0 149 5 3 1 72234
0 150 7 14 2 67551 63866
0 151 5 1 1 72239
0 152 7 29 2 70561 65895
0 153 5 2 1 72253
0 154 7 12 2 68891 72254
0 155 5 10 1 72284
0 156 7 4 2 72240 72285
0 157 5 1 1 72306
0 158 7 21 2 68736 64023
0 159 5 1 1 72310
0 160 7 9 2 70808 72311
0 161 7 13 2 62699 65623
0 162 5 2 1 72340
0 163 7 2 2 72331 72341
0 164 5 1 1 72355
0 165 7 1 2 157 164
0 166 5 1 1 165
0 167 7 1 2 67319 166
0 168 5 1 1 167
0 169 7 1 2 72236 168
0 170 5 1 1 169
0 171 7 1 2 65266 170
0 172 5 1 1 171
0 173 7 22 2 68737 65267
0 174 5 1 1 72357
0 175 7 13 2 62463 65624
0 176 5 1 1 72379
0 177 7 3 2 72358 72380
0 178 5 5 1 72392
0 179 7 3 2 66800 71552
0 180 5 1 1 72400
0 181 7 1 2 72395 180
0 182 5 2 1 181
0 183 7 1 2 71139 72403
0 184 5 1 1 183
0 185 7 11 2 67552 70183
0 186 5 1 1 72405
0 187 7 12 2 68892 70562
0 188 5 1 1 72416
0 189 7 4 2 63867 72417
0 190 5 3 1 72428
0 191 7 1 2 186 72432
0 192 5 1 1 191
0 193 7 1 2 66801 192
0 194 5 1 1 193
0 195 7 43 2 70184 65625
0 196 5 4 1 72435
0 197 7 4 2 68738 72436
0 198 5 8 1 72482
0 199 7 105 2 68893 65896
0 200 5 87 1 72494
0 201 7 28 2 67320 67553
0 202 5 16 1 72686
0 203 7 4 2 72495 72687
0 204 5 2 1 72730
0 205 7 2 2 72483 72731
0 206 5 4 1 72736
0 207 7 1 2 194 72738
0 208 7 1 2 184 207
0 209 7 1 2 172 208
0 210 5 1 1 209
0 211 7 1 2 71407 210
0 212 5 1 1 211
0 213 7 11 2 68739 68894
0 214 5 3 1 72742
0 215 7 5 2 70563 72753
0 216 7 7 2 67321 65897
0 217 5 2 1 72761
0 218 7 42 2 62700 64024
0 219 5 29 1 72770
0 220 7 2 2 65268 72812
0 221 7 2 2 72762 72841
0 222 5 1 1 72843
0 223 7 1 2 61942 222
0 224 5 1 1 223
0 225 7 1 2 72756 224
0 226 5 1 1 225
0 227 7 22 2 66802 70185
0 228 5 8 1 72845
0 229 7 10 2 65898 71641
0 230 5 1 1 72875
0 231 7 6 2 68740 70186
0 232 7 4 2 67322 72885
0 233 5 9 1 72891
0 234 7 23 2 62464 62701
0 235 5 8 1 72904
0 236 7 2 2 65269 72905
0 237 5 1 1 72935
0 238 7 1 2 72895 237
0 239 5 1 1 238
0 240 7 1 2 72876 239
0 241 5 1 1 240
0 242 7 1 2 72867 241
0 243 7 1 2 226 242
0 244 5 1 1 243
0 245 7 1 2 71029 244
0 246 5 1 1 245
0 247 7 1 2 212 246
0 248 5 1 1 247
0 249 7 1 2 71790 248
0 250 5 1 1 249
0 251 7 10 2 67101 63660
0 252 5 5 1 72937
0 253 7 4 2 71500 72947
0 254 5 95 1 72952
0 255 7 45 2 65270 70564
0 256 5 2 1 73051
0 257 7 5 2 63868 73052
0 258 5 4 1 73098
0 259 7 1 2 72486 73103
0 260 5 35 1 259
0 261 7 6 2 62465 71140
0 262 5 1 1 73142
0 263 7 23 2 67323 62702
0 264 5 1 1 73148
0 265 7 4 2 71998 73149
0 266 5 1 1 73171
0 267 7 1 2 262 266
0 268 5 5 1 267
0 269 7 1 2 73107 73175
0 270 5 1 1 269
0 271 7 53 2 63869 70565
0 272 5 37 1 73180
0 273 7 2 2 73181 72732
0 274 5 2 1 73270
0 275 7 1 2 73272 72237
0 276 5 2 1 275
0 277 7 1 2 70187 73274
0 278 5 1 1 277
0 279 7 1 2 270 278
0 280 5 1 1 279
0 281 7 1 2 71408 280
0 282 5 1 1 281
0 283 7 91 2 62466 63870
0 284 5 156 1 73276
0 285 7 3 2 73053 73277
0 286 5 4 1 73523
0 287 7 30 2 62703 70809
0 288 5 33 1 73530
0 289 7 1 2 73531 72484
0 290 5 1 1 289
0 291 7 1 2 73526 290
0 292 5 1 1 291
0 293 7 1 2 64025 292
0 294 5 1 1 293
0 295 7 25 2 63871 70188
0 296 5 1 1 73593
0 297 7 10 2 70566 73594
0 298 5 2 1 73618
0 299 7 3 2 72496 73619
0 300 7 3 2 67324 73630
0 301 5 1 1 73633
0 302 7 22 2 70189 65899
0 303 5 1 1 73636
0 304 7 2 2 71642 73637
0 305 5 7 1 73658
0 306 7 1 2 73104 73660
0 307 5 1 1 306
0 308 7 1 2 72906 307
0 309 5 1 1 308
0 310 7 1 2 301 309
0 311 7 1 2 294 310
0 312 5 1 1 311
0 313 7 1 2 71030 312
0 314 5 1 1 313
0 315 7 1 2 282 314
0 316 5 1 1 315
0 317 7 1 2 72956 316
0 318 5 1 1 317
0 319 7 6 2 66803 71999
0 320 5 1 1 73667
0 321 7 2 2 71715 73668
0 322 7 18 2 68500 63872
0 323 7 10 2 66582 62704
0 324 7 4 2 69659 73693
0 325 5 1 1 73703
0 326 7 1 2 73675 73704
0 327 7 1 2 73673 326
0 328 5 1 1 327
0 329 7 1 2 318 328
0 330 7 1 2 250 329
0 331 7 1 2 141 330
0 332 5 1 1 331
0 333 7 1 2 63418 332
0 334 5 1 1 333
0 335 7 12 2 62467 63419
0 336 5 3 1 73707
0 337 7 2 2 73719 73674
0 338 5 1 1 73722
0 339 7 8 2 68251 68895
0 340 7 1 2 61943 73724
0 341 5 2 1 340
0 342 7 1 2 338 73732
0 343 5 1 1 342
0 344 7 1 2 63873 343
0 345 5 1 1 344
0 346 7 15 2 61944 68896
0 347 5 1 1 73734
0 348 7 8 2 68252 70567
0 349 5 3 1 73749
0 350 7 1 2 73757 72396
0 351 5 1 1 350
0 352 7 1 2 73735 351
0 353 5 1 1 352
0 354 7 1 2 345 353
0 355 5 1 1 354
0 356 7 1 2 62705 355
0 357 5 1 1 356
0 358 7 1 2 71106 72393
0 359 5 1 1 358
0 360 7 25 2 64026 70568
0 361 5 4 1 73760
0 362 7 2 2 68741 73785
0 363 5 1 1 73789
0 364 7 1 2 71118 188
0 365 5 3 1 364
0 366 7 1 2 68253 73791
0 367 7 1 2 363 366
0 368 5 1 1 367
0 369 7 1 2 359 368
0 370 5 1 1 369
0 371 7 1 2 61945 370
0 372 5 1 1 371
0 373 7 1 2 357 372
0 374 5 2 1 373
0 375 7 1 2 63661 73794
0 376 5 1 1 375
0 377 7 21 2 61946 68501
0 378 5 1 1 73796
0 379 7 23 2 62706 68254
0 380 7 19 2 70190 70810
0 381 5 1 1 73840
0 382 7 8 2 64027 73841
0 383 7 1 2 73817 73859
0 384 5 3 1 383
0 385 7 1 2 73108 73143
0 386 5 1 1 385
0 387 7 1 2 73867 386
0 388 5 2 1 387
0 389 7 1 2 73797 73870
0 390 5 1 1 389
0 391 7 1 2 376 390
0 392 5 1 1 391
0 393 7 1 2 62276 392
0 394 5 1 1 393
0 395 7 3 2 68502 73182
0 396 5 8 1 73872
0 397 7 6 2 63662 71510
0 398 5 2 1 73883
0 399 7 1 2 73875 73889
0 400 5 2 1 399
0 401 7 1 2 73144 73891
0 402 5 1 1 401
0 403 7 7 2 63663 72000
0 404 7 1 2 73893 73818
0 405 5 1 1 404
0 406 7 1 2 402 405
0 407 5 1 1 406
0 408 7 1 2 67102 407
0 409 5 1 1 408
0 410 7 25 2 68255 68503
0 411 5 3 1 73900
0 412 7 9 2 62707 70569
0 413 5 19 1 73928
0 414 7 12 2 63874 64028
0 415 5 2 1 73956
0 416 7 5 2 70811 73957
0 417 5 1 1 73970
0 418 7 2 2 73929 73971
0 419 5 3 1 73975
0 420 7 1 2 73901 73976
0 421 5 1 1 420
0 422 7 1 2 409 421
0 423 5 1 1 422
0 424 7 1 2 70191 423
0 425 5 1 1 424
0 426 7 18 2 63664 65271
0 427 5 6 1 73980
0 428 7 8 2 67103 62468
0 429 7 4 2 63875 74004
0 430 5 1 1 74012
0 431 7 2 2 70570 71141
0 432 7 2 2 74013 74016
0 433 7 1 2 73981 74018
0 434 5 1 1 433
0 435 7 1 2 425 434
0 436 5 1 1 435
0 437 7 1 2 61947 436
0 438 5 1 1 437
0 439 7 1 2 394 438
0 440 5 1 1 439
0 441 7 1 2 71409 440
0 442 5 1 1 441
0 443 7 23 2 68256 63665
0 444 5 4 1 74020
0 445 7 5 2 62277 74021
0 446 5 6 1 74047
0 447 7 40 2 67554 68897
0 448 5 37 1 74058
0 449 7 6 2 65272 74098
0 450 7 5 2 62469 72957
0 451 7 1 2 74135 74141
0 452 5 1 1 451
0 453 7 1 2 74052 452
0 454 5 1 1 453
0 455 7 18 2 61698 61948
0 456 7 4 2 64822 74146
0 457 7 1 2 73183 74164
0 458 7 1 2 454 457
0 459 5 1 1 458
0 460 7 1 2 442 459
0 461 7 1 2 334 460
0 462 5 1 1 461
0 463 7 1 2 63046 462
0 464 5 1 1 463
0 465 7 23 2 70571 70812
0 466 5 3 1 74168
0 467 7 13 2 70192 74169
0 468 7 3 2 71279 74194
0 469 7 21 2 61949 67909
0 470 7 12 2 62708 69660
0 471 7 2 2 74210 74231
0 472 7 8 2 61699 64029
0 473 7 29 2 63420 63666
0 474 5 2 1 74253
0 475 7 11 2 62278 74254
0 476 5 2 1 74284
0 477 7 1 2 74245 74285
0 478 7 1 2 74243 477
0 479 7 1 2 74207 478
0 480 5 1 1 479
0 481 7 1 2 66338 480
0 482 7 1 2 464 481
0 483 5 1 1 482
0 484 7 45 2 66804 68257
0 485 5 48 1 74297
0 486 7 4 2 62470 74342
0 487 7 1 2 71142 74390
0 488 5 1 1 487
0 489 7 15 2 67325 63421
0 490 7 2 2 70813 74394
0 491 5 1 1 74409
0 492 7 1 2 72771 74410
0 493 5 1 1 492
0 494 7 1 2 488 493
0 495 5 2 1 494
0 496 7 9 2 70193 72958
0 497 7 1 2 74411 74413
0 498 5 1 1 497
0 499 7 23 2 67555 63422
0 500 5 1 1 74422
0 501 7 1 2 62279 73145
0 502 5 1 1 501
0 503 7 1 2 500 502
0 504 5 1 1 503
0 505 7 14 2 61950 63667
0 506 5 1 1 74445
0 507 7 1 2 65273 74446
0 508 7 1 2 504 507
0 509 5 1 1 508
0 510 7 1 2 498 509
0 511 5 1 1 510
0 512 7 1 2 68742 511
0 513 5 1 1 512
0 514 7 17 2 61951 67556
0 515 5 4 1 74459
0 516 7 3 2 72497 74460
0 517 5 2 1 74480
0 518 7 13 2 63876 65274
0 519 7 2 2 73708 74485
0 520 5 1 1 74498
0 521 7 1 2 74481 74499
0 522 5 1 1 521
0 523 7 1 2 513 522
0 524 5 1 1 523
0 525 7 1 2 71410 524
0 526 5 1 1 525
0 527 7 4 2 62471 72498
0 528 5 5 1 74500
0 529 7 7 2 68743 72001
0 530 5 6 1 74509
0 531 7 1 2 74504 74516
0 532 5 5 1 531
0 533 7 8 2 68504 70194
0 534 5 1 1 74527
0 535 7 2 2 534 73998
0 536 5 18 1 74535
0 537 7 3 2 62280 74537
0 538 5 2 1 74555
0 539 7 13 2 63668 70195
0 540 5 14 1 74560
0 541 7 2 2 67104 74561
0 542 5 1 1 74587
0 543 7 1 2 74558 542
0 544 5 7 1 543
0 545 7 1 2 74522 74589
0 546 5 1 1 545
0 547 7 11 2 63423 68898
0 548 5 1 1 74596
0 549 7 26 2 65275 65900
0 550 5 4 1 74607
0 551 7 6 2 74597 74608
0 552 5 1 1 74637
0 553 7 1 2 71280 74638
0 554 5 2 1 553
0 555 7 1 2 546 74643
0 556 5 1 1 555
0 557 7 1 2 62709 556
0 558 5 1 1 557
0 559 7 23 2 63424 65276
0 560 5 3 1 74645
0 561 7 14 2 63669 68744
0 562 5 2 1 74671
0 563 7 3 2 72499 73278
0 564 5 2 1 74687
0 565 7 1 2 74685 74690
0 566 5 1 1 565
0 567 7 1 2 74646 566
0 568 5 1 1 567
0 569 7 1 2 558 568
0 570 5 1 1 569
0 571 7 1 2 61952 570
0 572 5 1 1 571
0 573 7 3 2 62710 74523
0 574 5 2 1 74692
0 575 7 16 2 63425 70196
0 576 5 3 1 74697
0 577 7 3 2 72959 74698
0 578 7 1 2 74693 74716
0 579 5 1 1 578
0 580 7 1 2 64823 579
0 581 7 1 2 572 580
0 582 5 1 1 581
0 583 7 2 2 74059 73638
0 584 5 8 1 74719
0 585 7 9 2 62711 65277
0 586 5 2 1 74729
0 587 7 2 2 72002 74730
0 588 5 2 1 74740
0 589 7 1 2 74721 74742
0 590 5 11 1 589
0 591 7 75 2 67105 68505
0 592 5 22 1 74755
0 593 7 1 2 63426 74830
0 594 5 20 1 593
0 595 7 2 2 67326 74852
0 596 5 1 1 74872
0 597 7 1 2 74744 74873
0 598 5 1 1 597
0 599 7 21 2 63427 68506
0 600 5 5 1 74874
0 601 7 6 2 67106 74875
0 602 5 3 1 74900
0 603 7 2 2 74043 74906
0 604 5 7 1 74909
0 605 7 12 2 67557 65278
0 606 5 1 1 74918
0 607 7 1 2 74911 74919
0 608 5 1 1 607
0 609 7 1 2 598 608
0 610 5 1 1 609
0 611 7 1 2 68745 610
0 612 5 1 1 611
0 613 7 13 2 67558 68258
0 614 5 1 1 74930
0 615 7 3 2 67327 74931
0 616 7 1 2 73982 74943
0 617 5 1 1 616
0 618 7 1 2 612 617
0 619 5 1 1 618
0 620 7 1 2 66805 619
0 621 5 1 1 620
0 622 7 10 2 67107 67559
0 623 5 1 1 74946
0 624 7 2 2 61953 74947
0 625 7 2 2 73902 72359
0 626 7 1 2 74956 74958
0 627 5 1 1 626
0 628 7 1 2 69661 627
0 629 7 1 2 621 628
0 630 5 1 1 629
0 631 7 1 2 61700 630
0 632 7 1 2 582 631
0 633 5 1 1 632
0 634 7 1 2 526 633
0 635 5 1 1 634
0 636 7 1 2 65626 635
0 637 5 1 1 636
0 638 7 17 2 64824 70572
0 639 7 19 2 70814 72772
0 640 5 7 1 74977
0 641 7 2 2 74528 74978
0 642 5 2 1 75003
0 643 7 1 2 67108 75004
0 644 5 1 1 643
0 645 7 1 2 74053 644
0 646 5 1 1 645
0 647 7 1 2 61954 646
0 648 5 1 1 647
0 649 7 7 2 67328 72500
0 650 5 1 1 75007
0 651 7 1 2 75008 74717
0 652 5 1 1 651
0 653 7 1 2 648 652
0 654 5 1 1 653
0 655 7 1 2 63877 654
0 656 5 1 1 655
0 657 7 4 2 73842 72907
0 658 7 22 2 61955 67109
0 659 5 1 1 75018
0 660 7 2 2 71630 75019
0 661 7 1 2 75014 75040
0 662 5 1 1 661
0 663 7 1 2 656 662
0 664 5 1 1 663
0 665 7 1 2 74960 664
0 666 5 1 1 665
0 667 7 16 2 68259 69662
0 668 5 1 1 75042
0 669 7 2 2 74756 75043
0 670 5 1 1 75058
0 671 7 1 2 75059 73172
0 672 5 1 1 671
0 673 7 4 2 63878 64825
0 674 7 3 2 70573 75060
0 675 7 1 2 74286 75064
0 676 5 1 1 675
0 677 7 1 2 672 676
0 678 5 1 1 677
0 679 7 1 2 66806 678
0 680 5 1 1 679
0 681 7 1 2 61701 680
0 682 7 1 2 666 681
0 683 5 1 1 682
0 684 7 10 2 62712 63670
0 685 7 1 2 75067 73669
0 686 5 2 1 685
0 687 7 3 2 68507 65901
0 688 7 2 2 74423 75079
0 689 5 1 1 75082
0 690 7 1 2 68899 75083
0 691 5 1 1 690
0 692 7 1 2 75077 691
0 693 5 1 1 692
0 694 7 1 2 70197 73720
0 695 7 1 2 693 694
0 696 5 1 1 695
0 697 7 18 2 66807 63428
0 698 5 1 1 75084
0 699 7 15 2 61956 68260
0 700 5 3 1 75102
0 701 7 4 2 698 75117
0 702 5 52 1 75120
0 703 7 13 2 63671 68900
0 704 7 1 2 75124 75176
0 705 5 1 1 704
0 706 7 1 2 696 705
0 707 5 1 1 706
0 708 7 1 2 70574 707
0 709 5 1 1 708
0 710 7 5 2 63672 75125
0 711 7 1 2 71143 75189
0 712 5 1 1 711
0 713 7 1 2 709 712
0 714 5 1 1 713
0 715 7 1 2 63879 714
0 716 5 1 1 715
0 717 7 7 2 63673 70575
0 718 5 4 1 75194
0 719 7 3 2 68901 75195
0 720 5 1 1 75205
0 721 7 5 2 68508 72003
0 722 7 1 2 70198 75208
0 723 5 1 1 722
0 724 7 1 2 720 723
0 725 5 1 1 724
0 726 7 1 2 62713 725
0 727 5 1 1 726
0 728 7 13 2 67560 63674
0 729 7 3 2 64030 75213
0 730 7 1 2 70576 75226
0 731 5 1 1 730
0 732 7 1 2 727 731
0 733 5 1 1 732
0 734 7 1 2 75126 733
0 735 5 1 1 734
0 736 7 1 2 716 735
0 737 5 1 1 736
0 738 7 1 2 69663 737
0 739 5 1 1 738
0 740 7 10 2 61957 62714
0 741 5 2 1 75229
0 742 7 6 2 63429 75230
0 743 5 1 1 75241
0 744 7 1 2 75242 71765
0 745 5 1 1 744
0 746 7 1 2 739 745
0 747 5 1 1 746
0 748 7 1 2 62281 747
0 749 5 1 1 748
0 750 7 13 2 69664 70199
0 751 7 6 2 61958 74005
0 752 7 9 2 68509 70577
0 753 5 3 1 75266
0 754 7 19 2 63880 68902
0 755 7 2 2 75267 75278
0 756 7 1 2 75260 75297
0 757 5 1 1 756
0 758 7 2 2 72948 73876
0 759 5 1 1 75299
0 760 7 1 2 72004 75127
0 761 7 1 2 759 760
0 762 5 1 1 761
0 763 7 1 2 757 762
0 764 5 1 1 763
0 765 7 1 2 62715 764
0 766 5 1 1 765
0 767 7 10 2 61959 64031
0 768 5 2 1 75301
0 769 7 18 2 62472 68510
0 770 5 2 1 75313
0 771 7 1 2 75302 75314
0 772 5 1 1 771
0 773 7 4 2 68903 74255
0 774 7 1 2 72763 75333
0 775 5 1 1 774
0 776 7 1 2 772 775
0 777 5 1 1 776
0 778 7 8 2 67110 70578
0 779 5 1 1 75337
0 780 7 1 2 75338 72241
0 781 7 1 2 777 780
0 782 5 1 1 781
0 783 7 1 2 766 782
0 784 5 1 1 783
0 785 7 1 2 75247 784
0 786 5 1 1 785
0 787 7 1 2 66583 786
0 788 7 1 2 749 787
0 789 5 1 1 788
0 790 7 1 2 683 789
0 791 5 1 1 790
0 792 7 1 2 637 791
0 793 5 1 1 792
0 794 7 1 2 67910 793
0 795 5 1 1 794
0 796 7 12 2 67911 69665
0 797 7 4 2 63430 73798
0 798 7 4 2 68746 72688
0 799 5 4 1 75361
0 800 7 1 2 75357 75365
0 801 5 1 1 800
0 802 7 8 2 63881 72908
0 803 5 1 1 75369
0 804 7 6 2 63431 72960
0 805 5 1 1 75377
0 806 7 3 2 61960 72961
0 807 5 1 1 75383
0 808 7 1 2 805 807
0 809 5 5 1 808
0 810 7 1 2 75370 75386
0 811 5 1 1 810
0 812 7 1 2 801 811
0 813 5 1 1 812
0 814 7 1 2 66584 813
0 815 5 1 1 814
0 816 7 38 2 61702 66808
0 817 7 7 2 68261 68747
0 818 5 3 1 75429
0 819 7 2 2 62716 75430
0 820 5 1 1 75439
0 821 7 2 2 74948 75080
0 822 5 1 1 75441
0 823 7 1 2 63882 75442
0 824 5 1 1 823
0 825 7 1 2 820 824
0 826 5 1 1 825
0 827 7 1 2 67329 826
0 828 5 1 1 827
0 829 7 1 2 73903 71024
0 830 5 1 1 829
0 831 7 1 2 828 830
0 832 5 1 1 831
0 833 7 1 2 75391 832
0 834 5 1 1 833
0 835 7 1 2 815 834
0 836 5 1 1 835
0 837 7 1 2 70579 836
0 838 5 1 1 837
0 839 7 16 2 62717 63432
0 840 5 1 1 75443
0 841 7 3 2 68511 75444
0 842 7 29 2 66585 61961
0 843 7 2 2 71281 75462
0 844 7 1 2 75459 75491
0 845 5 1 1 844
0 846 7 4 2 68262 75392
0 847 7 4 2 62718 73676
0 848 5 1 1 75497
0 849 7 18 2 67330 63675
0 850 5 1 1 75501
0 851 7 17 2 67561 65902
0 852 5 25 1 75519
0 853 7 1 2 75502 75520
0 854 5 2 1 853
0 855 7 1 2 848 75561
0 856 5 1 1 855
0 857 7 1 2 75493 856
0 858 5 1 1 857
0 859 7 1 2 845 858
0 860 7 1 2 838 859
0 861 5 1 1 860
0 862 7 1 2 75345 861
0 863 5 1 1 862
0 864 7 1 2 67111 73873
0 865 5 1 1 864
0 866 7 1 2 74044 865
0 867 5 3 1 866
0 868 7 2 2 67331 75563
0 869 7 12 2 66809 63047
0 870 7 3 2 64826 75568
0 871 7 3 2 66586 65903
0 872 7 1 2 75580 75583
0 873 7 1 2 75566 872
0 874 5 1 1 873
0 875 7 1 2 863 874
0 876 5 1 1 875
0 877 7 1 2 68904 876
0 878 5 1 1 877
0 879 7 2 2 61962 71473
0 880 5 1 1 75586
0 881 7 14 2 66587 67332
0 882 7 2 2 69666 75588
0 883 5 2 1 75602
0 884 7 1 2 75604 71091
0 885 5 1 1 884
0 886 7 4 2 71282 73532
0 887 5 1 1 75606
0 888 7 1 2 885 75607
0 889 5 1 1 888
0 890 7 5 2 66588 73279
0 891 7 1 2 71463 75610
0 892 5 2 1 891
0 893 7 1 2 889 75615
0 894 5 1 1 893
0 895 7 1 2 73761 894
0 896 5 1 1 895
0 897 7 1 2 880 896
0 898 5 1 1 897
0 899 7 1 2 63433 898
0 900 5 1 1 899
0 901 7 10 2 62719 64827
0 902 5 2 1 75617
0 903 7 3 2 61703 75618
0 904 5 4 1 75629
0 905 7 11 2 70580 72005
0 906 5 1 1 75636
0 907 7 5 2 71283 75637
0 908 5 1 1 75647
0 909 7 1 2 75630 75648
0 910 5 1 1 909
0 911 7 6 2 62473 73184
0 912 5 11 1 75652
0 913 7 10 2 64032 69667
0 914 7 11 2 66589 67562
0 915 7 1 2 75669 75679
0 916 7 1 2 75653 915
0 917 5 1 1 916
0 918 7 1 2 910 917
0 919 5 1 1 918
0 920 7 1 2 61963 919
0 921 5 1 1 920
0 922 7 23 2 61704 67563
0 923 7 4 2 66810 75044
0 924 5 1 1 75713
0 925 7 1 2 75690 75714
0 926 5 1 1 925
0 927 7 1 2 921 926
0 928 7 1 2 900 927
0 929 5 1 1 928
0 930 7 1 2 72962 929
0 931 5 1 1 930
0 932 7 23 2 70581 71284
0 933 5 9 1 75717
0 934 7 2 2 63434 75718
0 935 7 1 2 74165 75749
0 936 5 1 1 935
0 937 7 42 2 61964 63435
0 938 5 31 1 75751
0 939 7 5 2 66590 75752
0 940 5 1 1 75824
0 941 7 3 2 61705 74298
0 942 5 2 1 75829
0 943 7 1 2 940 75832
0 944 5 7 1 943
0 945 7 1 2 71553 75834
0 946 5 1 1 945
0 947 7 23 2 61965 62474
0 948 5 1 1 75841
0 949 7 3 2 66591 75842
0 950 7 1 2 63436 75864
0 951 5 1 1 950
0 952 7 1 2 946 951
0 953 5 1 1 952
0 954 7 1 2 69668 71107
0 955 7 1 2 953 954
0 956 5 1 1 955
0 957 7 1 2 936 956
0 958 5 1 1 957
0 959 7 1 2 68512 958
0 960 5 1 1 959
0 961 7 18 2 66811 67564
0 962 5 1 1 75867
0 963 7 5 2 61706 75868
0 964 7 14 2 67333 70582
0 965 5 2 1 75890
0 966 7 1 2 75670 75431
0 967 7 1 2 75891 966
0 968 7 1 2 75885 967
0 969 5 1 1 968
0 970 7 1 2 960 969
0 971 7 1 2 931 970
0 972 5 1 1 971
0 973 7 1 2 67912 972
0 974 5 1 1 973
0 975 7 1 2 878 974
0 976 5 1 1 975
0 977 7 1 2 65279 976
0 978 5 1 1 977
0 979 7 1 2 68263 73983
0 980 5 2 1 979
0 981 7 3 2 65904 72743
0 982 7 12 2 68264 70200
0 983 5 3 1 75911
0 984 7 3 2 67112 74538
0 985 5 3 1 75926
0 986 7 41 2 68513 65280
0 987 5 7 1 75932
0 988 7 1 2 62282 75933
0 989 5 4 1 988
0 990 7 2 2 75929 75980
0 991 5 2 1 75984
0 992 7 1 2 75923 75985
0 993 5 1 1 992
0 994 7 1 2 75908 993
0 995 5 1 1 994
0 996 7 1 2 75906 995
0 997 5 1 1 996
0 998 7 1 2 67334 997
0 999 5 1 1 998
0 1000 7 1 2 74901 72360
0 1001 5 1 1 1000
0 1002 7 1 2 999 1001
0 1003 5 2 1 1002
0 1004 7 23 2 63048 64828
0 1005 5 1 1 75990
0 1006 7 5 2 66592 75991
0 1007 5 2 1 76013
0 1008 7 8 2 66812 65627
0 1009 7 1 2 76014 76020
0 1010 7 1 2 75988 1009
0 1011 5 1 1 1010
0 1012 7 1 2 61425 1011
0 1013 7 1 2 978 1012
0 1014 7 1 2 795 1013
0 1015 5 1 1 1014
0 1016 7 1 2 69876 1015
0 1017 7 1 2 483 1016
0 1018 5 1 1 1017
0 1019 7 35 2 61426 67913
0 1020 5 1 1 76028
0 1021 7 37 2 66339 63049
0 1022 5 1 1 76063
0 1023 7 3 2 1020 1022
0 1024 5 98 1 76100
0 1025 7 4 2 65009 75393
0 1026 5 1 1 76201
0 1027 7 11 2 68265 63883
0 1028 5 3 1 76205
0 1029 7 4 2 70583 76206
0 1030 5 3 1 76219
0 1031 7 4 2 67335 73109
0 1032 5 1 1 76226
0 1033 7 1 2 72501 76227
0 1034 5 2 1 1033
0 1035 7 1 2 76223 76230
0 1036 5 1 1 1035
0 1037 7 1 2 76202 1036
0 1038 5 1 1 1037
0 1039 7 6 2 63437 75463
0 1040 7 19 2 68905 65281
0 1041 5 1 1 76238
0 1042 7 3 2 65905 72381
0 1043 5 1 1 76257
0 1044 7 2 2 76239 76258
0 1045 5 2 1 76260
0 1046 7 2 2 67565 76261
0 1047 5 1 1 76264
0 1048 7 1 2 63884 76265
0 1049 5 1 1 1048
0 1050 7 18 2 62720 71285
0 1051 5 4 1 76266
0 1052 7 1 2 65010 76267
0 1053 5 1 1 1052
0 1054 7 1 2 1049 1053
0 1055 5 1 1 1054
0 1056 7 1 2 76232 1055
0 1057 5 1 1 1056
0 1058 7 1 2 1038 1057
0 1059 5 1 1 1058
0 1060 7 1 2 62283 1059
0 1061 5 1 1 1060
0 1062 7 9 2 61707 65011
0 1063 7 5 2 65628 74694
0 1064 5 1 1 76297
0 1065 7 2 2 75912 76298
0 1066 5 1 1 76302
0 1067 7 1 2 73819 75649
0 1068 5 1 1 1067
0 1069 7 27 2 65629 65906
0 1070 5 6 1 76304
0 1071 7 17 2 68906 76305
0 1072 5 4 1 76337
0 1073 7 19 2 63438 68748
0 1074 7 6 2 67336 76358
0 1075 7 1 2 76338 76377
0 1076 5 1 1 1075
0 1077 7 1 2 1068 1076
0 1078 5 1 1 1077
0 1079 7 1 2 65282 1078
0 1080 5 1 1 1079
0 1081 7 1 2 1066 1080
0 1082 5 1 1 1081
0 1083 7 1 2 67113 1082
0 1084 5 1 1 1083
0 1085 7 9 2 65283 75128
0 1086 7 1 2 71616 76383
0 1087 5 1 1 1086
0 1088 7 1 2 1084 1087
0 1089 5 1 1 1088
0 1090 7 1 2 76288 1089
0 1091 5 1 1 1090
0 1092 7 1 2 1061 1091
0 1093 5 1 1 1092
0 1094 7 1 2 63676 1093
0 1095 5 1 1 1094
0 1096 7 2 2 65630 74524
0 1097 7 1 2 75020 76392
0 1098 5 1 1 1097
0 1099 7 12 2 62284 68266
0 1100 5 1 1 76394
0 1101 7 1 2 76395 75650
0 1102 5 1 1 1101
0 1103 7 1 2 1098 1102
0 1104 5 1 1 1103
0 1105 7 1 2 62721 1104
0 1106 5 1 1 1105
0 1107 7 2 2 67114 73233
0 1108 5 5 1 76406
0 1109 7 1 2 75129 76408
0 1110 5 2 1 1109
0 1111 7 5 2 65631 76359
0 1112 5 1 1 76415
0 1113 7 4 2 62285 68907
0 1114 7 3 2 65907 76420
0 1115 5 1 1 76424
0 1116 7 1 2 67337 76425
0 1117 5 1 1 1116
0 1118 7 1 2 659 1117
0 1119 5 1 1 1118
0 1120 7 1 2 76416 1119
0 1121 5 1 1 1120
0 1122 7 1 2 76413 1121
0 1123 7 1 2 1106 1122
0 1124 5 1 1 1123
0 1125 7 1 2 65284 1124
0 1126 5 1 1 1125
0 1127 7 1 2 62286 76303
0 1128 5 1 1 1127
0 1129 7 1 2 1126 1128
0 1130 5 1 1 1129
0 1131 7 11 2 61708 68514
0 1132 7 1 2 65012 76427
0 1133 7 1 2 1130 1132
0 1134 5 1 1 1133
0 1135 7 1 2 1095 1134
0 1136 5 1 1 1135
0 1137 7 1 2 76103 1136
0 1138 5 1 1 1137
0 1139 7 11 2 68267 71886
0 1140 5 25 1 76438
0 1141 7 5 2 66813 71887
0 1142 5 3 1 76474
0 1143 7 2 2 76449 76479
0 1144 5 2 1 76482
0 1145 7 6 2 74343 76483
0 1146 7 4 2 62722 71554
0 1147 5 2 1 76492
0 1148 7 1 2 64033 76493
0 1149 5 1 1 1148
0 1150 7 1 2 73234 1149
0 1151 5 2 1 1150
0 1152 7 1 2 62475 76498
0 1153 5 1 1 1152
0 1154 7 3 2 72773 73185
0 1155 5 1 1 76500
0 1156 7 1 2 1153 1155
0 1157 5 7 1 1156
0 1158 7 3 2 70201 76503
0 1159 7 1 2 76486 76510
0 1160 5 1 1 1159
0 1161 7 3 2 65632 72813
0 1162 5 15 1 76513
0 1163 7 11 2 71791 75753
0 1164 7 1 2 76516 76531
0 1165 5 1 1 1164
0 1166 7 1 2 1160 1165
0 1167 5 1 1 1166
0 1168 7 26 2 66340 66593
0 1169 7 14 2 65013 70815
0 1170 7 2 2 63050 76568
0 1171 7 1 2 76542 76582
0 1172 7 1 2 1167 1171
0 1173 5 1 1 1172
0 1174 7 1 2 1138 1173
0 1175 5 1 1 1174
0 1176 7 1 2 69669 1175
0 1177 5 1 1 1176
0 1178 7 9 2 61427 64829
0 1179 7 9 2 68908 70202
0 1180 5 2 1 76593
0 1181 7 5 2 72255 76594
0 1182 5 2 1 76604
0 1183 7 6 2 67338 63885
0 1184 5 1 1 76611
0 1185 7 10 2 66814 63677
0 1186 5 2 1 76617
0 1187 7 2 2 76612 76618
0 1188 7 1 2 76605 76629
0 1189 5 1 1 1188
0 1190 7 4 2 61966 75934
0 1191 5 5 1 76631
0 1192 7 1 2 76632 76299
0 1193 5 1 1 1192
0 1194 7 1 2 1189 1193
0 1195 5 1 1 1194
0 1196 7 1 2 67115 1195
0 1197 5 1 1 1196
0 1198 7 1 2 63678 73110
0 1199 5 1 1 1198
0 1200 7 1 2 75268 73595
0 1201 5 1 1 1200
0 1202 7 1 2 1199 1201
0 1203 5 1 1 1202
0 1204 7 13 2 62287 67339
0 1205 7 3 2 66815 72502
0 1206 7 1 2 76640 76653
0 1207 7 1 2 1203 1206
0 1208 5 1 1 1207
0 1209 7 1 2 1197 1208
0 1210 5 2 1 1209
0 1211 7 23 2 66594 63051
0 1212 7 1 2 65014 76658
0 1213 7 1 2 76656 1212
0 1214 5 1 1 1213
0 1215 7 49 2 65285 65633
0 1216 5 1 1 76681
0 1217 7 7 2 65908 71286
0 1218 5 1 1 76730
0 1219 7 9 2 67566 73367
0 1220 5 4 1 76737
0 1221 7 4 2 76731 76746
0 1222 5 1 1 76750
0 1223 7 2 2 76682 76751
0 1224 7 10 2 61709 62288
0 1225 7 2 2 76756 74211
0 1226 7 1 2 75334 76766
0 1227 7 1 2 76754 1226
0 1228 5 1 1 1227
0 1229 7 1 2 1214 1228
0 1230 5 1 1 1229
0 1231 7 1 2 76584 1230
0 1232 5 1 1 1231
0 1233 7 1 2 69460 1232
0 1234 7 1 2 1177 1233
0 1235 7 1 2 1018 1234
0 1236 5 1 1 1235
0 1237 7 22 2 69670 65286
0 1238 7 5 2 66595 76768
0 1239 7 1 2 74876 76790
0 1240 5 1 1 1239
0 1241 7 13 2 65287 72963
0 1242 5 1 1 76795
0 1243 7 1 2 61710 76796
0 1244 5 1 1 1243
0 1245 7 22 2 62289 63439
0 1246 5 1 1 76808
0 1247 7 4 2 66596 76809
0 1248 7 2 2 64034 74562
0 1249 7 1 2 76830 76834
0 1250 5 1 1 1249
0 1251 7 1 2 1244 1250
0 1252 5 1 1 1251
0 1253 7 19 2 64830 70816
0 1254 7 1 2 62723 76836
0 1255 7 1 2 1252 1254
0 1256 5 1 1 1255
0 1257 7 1 2 1240 1256
0 1258 5 1 1 1257
0 1259 7 1 2 69877 1258
0 1260 5 1 1 1259
0 1261 7 2 2 70817 76450
0 1262 7 5 2 70203 71031
0 1263 7 8 2 62724 65015
0 1264 5 2 1 76862
0 1265 7 1 2 76857 76863
0 1266 7 1 2 76855 1265
0 1267 5 1 1 1266
0 1268 7 1 2 1260 1267
0 1269 5 1 1 1268
0 1270 7 1 2 61967 1269
0 1271 5 1 1 1270
0 1272 7 41 2 69878 65288
0 1273 5 1 1 76872
0 1274 7 7 2 68515 76873
0 1275 5 5 1 76913
0 1276 7 33 2 65016 70204
0 1277 5 5 1 76925
0 1278 7 5 2 63679 76926
0 1279 5 3 1 76963
0 1280 7 1 2 76920 76968
0 1281 5 8 1 1280
0 1282 7 1 2 62290 76971
0 1283 5 3 1 1282
0 1284 7 1 2 72938 76874
0 1285 5 1 1 1284
0 1286 7 2 2 76979 1285
0 1287 5 4 1 76982
0 1288 7 14 2 61711 62725
0 1289 7 3 2 76837 76988
0 1290 5 1 1 77002
0 1291 7 1 2 63440 77003
0 1292 7 1 2 76984 1291
0 1293 5 1 1 1292
0 1294 7 1 2 1271 1293
0 1295 5 1 1 1294
0 1296 7 1 2 70584 1295
0 1297 5 1 1 1296
0 1298 7 3 2 66597 74232
0 1299 5 1 1 77005
0 1300 7 1 2 71092 1299
0 1301 5 11 1 1300
0 1302 7 12 2 70818 73762
0 1303 5 1 1 77019
0 1304 7 1 2 74344 76985
0 1305 5 1 1 1304
0 1306 7 15 2 61968 65017
0 1307 5 5 1 77031
0 1308 7 2 2 77032 74699
0 1309 5 2 1 77051
0 1310 7 1 2 1305 77053
0 1311 5 2 1 1310
0 1312 7 1 2 77020 77055
0 1313 5 1 1 1312
0 1314 7 8 2 65018 71888
0 1315 5 7 1 77057
0 1316 7 2 2 65634 74639
0 1317 5 2 1 77072
0 1318 7 2 2 77065 77073
0 1319 7 1 2 61969 77076
0 1320 5 1 1 1319
0 1321 7 1 2 1313 1320
0 1322 5 1 1 1321
0 1323 7 1 2 77008 1322
0 1324 5 1 1 1323
0 1325 7 25 2 61970 64831
0 1326 7 4 2 68909 71792
0 1327 7 2 2 77078 77103
0 1328 5 1 1 77107
0 1329 7 7 2 61712 69879
0 1330 7 7 2 65289 76306
0 1331 5 1 1 77116
0 1332 7 1 2 77109 77117
0 1333 7 1 2 77108 1332
0 1334 5 1 1 1333
0 1335 7 1 2 1324 1334
0 1336 7 1 2 1297 1335
0 1337 5 1 1 1336
0 1338 7 1 2 63052 1337
0 1339 5 1 1 1338
0 1340 7 11 2 69880 70585
0 1341 7 5 2 77123 73843
0 1342 7 1 2 63680 75671
0 1343 7 2 2 77134 1342
0 1344 7 18 2 61971 62291
0 1345 7 4 2 62726 77141
0 1346 7 13 2 67914 63441
0 1347 7 2 2 61713 77163
0 1348 7 1 2 77159 77176
0 1349 7 1 2 77139 1348
0 1350 5 1 1 1349
0 1351 7 1 2 1339 1350
0 1352 5 1 1 1351
0 1353 7 1 2 61428 1352
0 1354 5 1 1 1353
0 1355 7 32 2 66341 61714
0 1356 7 3 2 61972 77178
0 1357 7 2 2 62292 75445
0 1358 7 1 2 63053 77213
0 1359 7 1 2 77210 1358
0 1360 7 1 2 77140 1359
0 1361 5 1 1 1360
0 1362 7 1 2 1354 1361
0 1363 5 1 1 1362
0 1364 7 1 2 71287 1363
0 1365 5 1 1 1364
0 1366 7 53 2 61429 63054
0 1367 5 5 1 77215
0 1368 7 5 2 63886 72503
0 1369 5 3 1 77273
0 1370 7 3 2 75892 77274
0 1371 5 3 1 77281
0 1372 7 1 2 63442 77282
0 1373 5 2 1 1372
0 1374 7 1 2 74345 76300
0 1375 5 1 1 1374
0 1376 7 1 2 77287 1375
0 1377 5 1 1 1376
0 1378 7 1 2 65290 1377
0 1379 5 1 1 1378
0 1380 7 20 2 63443 63887
0 1381 5 3 1 77289
0 1382 7 12 2 66816 70586
0 1383 7 1 2 77290 77312
0 1384 5 1 1 1383
0 1385 7 1 2 1379 1384
0 1386 5 1 1 1385
0 1387 7 1 2 69881 1386
0 1388 5 1 1 1387
0 1389 7 15 2 65019 70587
0 1390 5 3 1 77324
0 1391 7 10 2 68910 74609
0 1392 7 10 2 63888 65635
0 1393 5 3 1 77352
0 1394 7 1 2 77342 77353
0 1395 5 1 1 1394
0 1396 7 1 2 77339 1395
0 1397 5 1 1 1396
0 1398 7 2 2 73709 1397
0 1399 5 1 1 77365
0 1400 7 1 2 61973 77366
0 1401 5 1 1 1400
0 1402 7 1 2 1388 1401
0 1403 5 1 1 1402
0 1404 7 1 2 62293 1403
0 1405 5 1 1 1404
0 1406 7 2 2 76875 71617
0 1407 7 1 2 75754 77367
0 1408 5 1 1 1407
0 1409 7 1 2 1405 1408
0 1410 5 1 1 1409
0 1411 7 1 2 63681 1410
0 1412 5 1 1 1411
0 1413 7 1 2 73280 72877
0 1414 5 1 1 1413
0 1415 7 1 2 71501 1414
0 1416 5 1 1 1415
0 1417 7 17 2 61974 69882
0 1418 5 1 1 77369
0 1419 7 1 2 77370 74647
0 1420 7 1 2 1416 1419
0 1421 5 1 1 1420
0 1422 7 1 2 1412 1421
0 1423 5 1 1 1422
0 1424 7 1 2 71411 1423
0 1425 5 1 1 1424
0 1426 7 15 2 66817 69671
0 1427 7 1 2 77386 75989
0 1428 5 1 1 1427
0 1429 7 14 2 63444 64832
0 1430 7 5 2 68749 70819
0 1431 5 1 1 77415
0 1432 7 4 2 67116 64035
0 1433 7 2 2 61975 77420
0 1434 5 1 1 77424
0 1435 7 1 2 71793 74136
0 1436 5 1 1 1435
0 1437 7 1 2 1434 1436
0 1438 5 1 1 1437
0 1439 7 1 2 77416 1438
0 1440 5 1 1 1439
0 1441 7 20 2 62294 62476
0 1442 5 2 1 77426
0 1443 7 6 2 63682 77427
0 1444 7 6 2 65909 76240
0 1445 7 1 2 77448 77454
0 1446 5 1 1 1445
0 1447 7 1 2 1440 1446
0 1448 5 1 1 1447
0 1449 7 1 2 77401 1448
0 1450 5 1 1 1449
0 1451 7 1 2 1428 1450
0 1452 5 1 1 1451
0 1453 7 1 2 65636 1452
0 1454 5 1 1 1453
0 1455 7 19 2 67340 68268
0 1456 5 1 1 77460
0 1457 7 2 2 72504 76769
0 1458 5 1 1 77479
0 1459 7 1 2 77461 77480
0 1460 5 1 1 1459
0 1461 7 5 2 64036 76838
0 1462 7 1 2 76810 77481
0 1463 5 1 1 1462
0 1464 7 1 2 1460 1463
0 1465 5 1 1 1464
0 1466 7 1 2 66818 1465
0 1467 5 1 1 1466
0 1468 7 17 2 70820 74099
0 1469 5 3 1 77486
0 1470 7 5 2 77487 74346
0 1471 7 1 2 74014 77506
0 1472 5 1 1 1471
0 1473 7 6 2 63445 76641
0 1474 7 14 2 65910 72814
0 1475 5 3 1 77517
0 1476 7 4 2 70588 77518
0 1477 5 3 1 77534
0 1478 7 1 2 77511 77535
0 1479 5 1 1 1478
0 1480 7 1 2 1472 1479
0 1481 5 1 1 1480
0 1482 7 1 2 65291 1481
0 1483 5 1 1 1482
0 1484 7 10 2 62295 70205
0 1485 5 11 1 77541
0 1486 7 1 2 75103 77542
0 1487 5 1 1 1486
0 1488 7 1 2 1483 1487
0 1489 5 1 1 1488
0 1490 7 1 2 64833 1489
0 1491 5 1 1 1490
0 1492 7 1 2 1467 1491
0 1493 5 1 1 1492
0 1494 7 1 2 63683 1493
0 1495 5 1 1 1494
0 1496 7 3 2 64834 77428
0 1497 7 1 2 77507 77562
0 1498 5 1 1 1497
0 1499 7 17 2 67117 67341
0 1500 7 4 2 66819 77565
0 1501 7 2 2 71686 72418
0 1502 7 1 2 77582 77586
0 1503 5 1 1 1502
0 1504 7 1 2 1498 1503
0 1505 5 1 1 1504
0 1506 7 1 2 63889 1505
0 1507 5 1 1 1506
0 1508 7 1 2 76839 75243
0 1509 5 1 1 1508
0 1510 7 1 2 1507 1509
0 1511 5 1 1 1510
0 1512 7 1 2 75935 1511
0 1513 5 1 1 1512
0 1514 7 1 2 69883 1513
0 1515 7 1 2 1495 1514
0 1516 7 1 2 1454 1515
0 1517 5 1 1 1516
0 1518 7 1 2 69672 76657
0 1519 5 1 1 1518
0 1520 7 3 2 74100 76840
0 1521 7 15 2 62477 63684
0 1522 5 1 1 77591
0 1523 7 12 2 62296 63890
0 1524 5 2 1 77606
0 1525 7 6 2 77592 77607
0 1526 5 1 1 77620
0 1527 7 1 2 77621 74700
0 1528 5 1 1 1527
0 1529 7 7 2 62478 73596
0 1530 5 3 1 77626
0 1531 7 1 2 77633 74295
0 1532 5 2 1 1531
0 1533 7 8 2 61976 76451
0 1534 5 2 1 77638
0 1535 7 1 2 77636 77639
0 1536 5 1 1 1535
0 1537 7 1 2 1528 1536
0 1538 5 3 1 1537
0 1539 7 1 2 77588 77648
0 1540 5 1 1 1539
0 1541 7 1 2 65020 1540
0 1542 7 1 2 1519 1541
0 1543 5 1 1 1542
0 1544 7 1 2 61715 1543
0 1545 7 1 2 1517 1544
0 1546 5 1 1 1545
0 1547 7 1 2 1425 1546
0 1548 5 1 1 1547
0 1549 7 1 2 77216 1548
0 1550 5 1 1 1549
0 1551 7 1 2 64610 1550
0 1552 7 1 2 1365 1551
0 1553 5 1 1 1552
0 1554 7 1 2 1236 1553
0 1555 5 1 1 1554
0 1556 7 1 2 64427 1555
0 1557 5 1 1 1556
0 1558 7 23 2 66820 69884
0 1559 5 5 1 77651
0 1560 7 9 2 69673 70589
0 1561 7 6 2 66598 77679
0 1562 5 2 1 77688
0 1563 7 1 2 77694 75632
0 1564 5 4 1 1563
0 1565 7 1 2 72964 77696
0 1566 5 2 1 1565
0 1567 7 8 2 64835 76989
0 1568 7 1 2 73677 77702
0 1569 5 2 1 1568
0 1570 7 9 2 63685 73281
0 1571 5 2 1 77712
0 1572 7 6 2 68516 73368
0 1573 5 9 1 77723
0 1574 7 2 2 71412 77729
0 1575 7 1 2 77721 77738
0 1576 5 1 1 1575
0 1577 7 1 2 77710 1576
0 1578 5 1 1 1577
0 1579 7 1 2 70590 1578
0 1580 5 1 1 1579
0 1581 7 1 2 77700 1580
0 1582 5 1 1 1581
0 1583 7 1 2 70206 1582
0 1584 5 1 1 1583
0 1585 7 6 2 63686 71768
0 1586 7 11 2 65637 71288
0 1587 5 1 1 77746
0 1588 7 2 2 69674 77747
0 1589 7 1 2 77740 77757
0 1590 5 1 1 1589
0 1591 7 1 2 1584 1590
0 1592 5 1 1 1591
0 1593 7 1 2 70821 1592
0 1594 5 1 1 1593
0 1595 7 10 2 62297 67567
0 1596 5 2 1 77759
0 1597 7 2 2 61716 77760
0 1598 7 3 2 63687 71555
0 1599 5 2 1 77773
0 1600 7 2 2 64836 77774
0 1601 7 1 2 77771 77778
0 1602 5 1 1 1601
0 1603 7 1 2 1594 1602
0 1604 5 1 1 1603
0 1605 7 1 2 64037 1604
0 1606 5 1 1 1605
0 1607 7 3 2 71120 71032
0 1608 5 2 1 77780
0 1609 7 1 2 71556 77781
0 1610 5 1 1 1609
0 1611 7 5 2 69675 72256
0 1612 7 1 2 71697 77785
0 1613 5 1 1 1612
0 1614 7 1 2 1610 1613
0 1615 5 1 1 1614
0 1616 7 1 2 71794 1615
0 1617 5 1 1 1616
0 1618 7 1 2 1606 1617
0 1619 5 1 1 1618
0 1620 7 1 2 77652 1619
0 1621 5 1 1 1620
0 1622 7 13 2 62298 62727
0 1623 5 2 1 77790
0 1624 7 1 2 77791 71766
0 1625 5 1 1 1624
0 1626 7 22 2 65638 70822
0 1627 5 2 1 77805
0 1628 7 7 2 64038 77806
0 1629 5 9 1 77829
0 1630 7 1 2 72282 77836
0 1631 5 2 1 1630
0 1632 7 1 2 62479 77845
0 1633 5 1 1 1632
0 1634 7 9 2 62299 65639
0 1635 5 1 1 77847
0 1636 7 6 2 63891 72257
0 1637 5 2 1 77856
0 1638 7 1 2 1635 77862
0 1639 7 1 2 1633 1638
0 1640 5 1 1 1639
0 1641 7 1 2 68517 1640
0 1642 5 1 1 1641
0 1643 7 1 2 75503 71511
0 1644 5 2 1 1643
0 1645 7 1 2 70591 74517
0 1646 5 1 1 1645
0 1647 7 9 2 68518 65640
0 1648 5 1 1 77866
0 1649 7 1 2 67118 1648
0 1650 7 1 2 1646 1649
0 1651 5 1 1 1650
0 1652 7 1 2 77864 1651
0 1653 7 1 2 1642 1652
0 1654 5 1 1 1653
0 1655 7 1 2 65292 1654
0 1656 5 1 1 1655
0 1657 7 6 2 74757 73369
0 1658 5 4 1 77875
0 1659 7 2 2 77021 77876
0 1660 5 2 1 77885
0 1661 7 1 2 1656 77887
0 1662 5 1 1 1661
0 1663 7 1 2 69676 1662
0 1664 5 1 1 1663
0 1665 7 1 2 1625 1664
0 1666 5 1 1 1665
0 1667 7 1 2 66599 1666
0 1668 5 1 1 1667
0 1669 7 3 2 64039 71557
0 1670 5 1 1 77889
0 1671 7 1 2 68519 77890
0 1672 5 1 1 1671
0 1673 7 1 2 67568 1672
0 1674 7 1 2 71628 1673
0 1675 5 1 1 1674
0 1676 7 2 2 65293 71033
0 1677 7 12 2 68520 68911
0 1678 7 3 2 65641 71186
0 1679 5 4 1 77906
0 1680 7 1 2 77894 77909
0 1681 5 1 1 1680
0 1682 7 1 2 62728 1681
0 1683 5 1 1 1682
0 1684 7 1 2 77892 1683
0 1685 7 1 2 1675 1684
0 1686 5 1 1 1685
0 1687 7 1 2 1668 1686
0 1688 5 1 1 1687
0 1689 7 1 2 69885 1688
0 1690 5 1 1 1689
0 1691 7 1 2 71889 73628
0 1692 5 3 1 1691
0 1693 7 11 2 62480 65021
0 1694 7 1 2 77782 77916
0 1695 7 1 2 77913 1694
0 1696 5 1 1 1695
0 1697 7 1 2 1690 1696
0 1698 5 1 1 1697
0 1699 7 1 2 61977 1698
0 1700 5 1 1 1699
0 1701 7 1 2 1621 1700
0 1702 5 1 1 1701
0 1703 7 1 2 63446 1702
0 1704 5 1 1 1703
0 1705 7 10 2 66821 70823
0 1706 7 19 2 64040 70207
0 1707 5 2 1 77937
0 1708 7 3 2 77927 77938
0 1709 5 1 1 77958
0 1710 7 1 2 77959 72242
0 1711 5 1 1 1710
0 1712 7 1 2 73733 1711
0 1713 5 1 1 1712
0 1714 7 11 2 62481 70592
0 1715 5 3 1 77961
0 1716 7 2 2 71769 77962
0 1717 7 1 2 1713 77975
0 1718 5 1 1 1717
0 1719 7 1 2 62482 71558
0 1720 5 7 1 1719
0 1721 7 2 2 65294 77977
0 1722 5 1 1 77984
0 1723 7 8 2 70593 72599
0 1724 5 18 1 77986
0 1725 7 3 2 67569 77994
0 1726 7 1 2 75494 78012
0 1727 7 1 2 77985 1726
0 1728 5 1 1 1727
0 1729 7 1 2 1718 1728
0 1730 5 1 1 1729
0 1731 7 1 2 63688 1730
0 1732 5 1 1 1731
0 1733 7 1 2 75830 72737
0 1734 5 1 1 1733
0 1735 7 1 2 1732 1734
0 1736 5 1 1 1735
0 1737 7 1 2 69677 1736
0 1738 5 1 1 1737
0 1739 7 5 2 61978 72909
0 1740 7 1 2 67119 78015
0 1741 7 1 2 76858 75298
0 1742 7 1 2 1740 1741
0 1743 5 1 1 1742
0 1744 7 1 2 1738 1743
0 1745 5 1 1 1744
0 1746 7 1 2 69886 1745
0 1747 5 1 1 1746
0 1748 7 1 2 1704 1747
0 1749 5 1 1 1748
0 1750 7 1 2 64611 1749
0 1751 5 1 1 1750
0 1752 7 12 2 62483 64041
0 1753 5 1 1 78020
0 1754 7 15 2 65022 65911
0 1755 7 2 2 78032 75231
0 1756 7 1 2 78021 78047
0 1757 5 1 1 1756
0 1758 7 39 2 63447 69887
0 1759 5 4 1 78049
0 1760 7 5 2 66822 78050
0 1761 5 1 1 78092
0 1762 7 1 2 67342 78093
0 1763 5 1 1 1762
0 1764 7 1 2 1757 1763
0 1765 5 1 1 1764
0 1766 7 1 2 74758 1765
0 1767 5 1 1 1766
0 1768 7 22 2 68269 69888
0 1769 5 7 1 78097
0 1770 7 8 2 64042 65023
0 1771 7 3 2 70824 78126
0 1772 7 1 2 77429 78134
0 1773 5 1 1 1772
0 1774 7 1 2 78119 1773
0 1775 5 1 1 1774
0 1776 7 3 2 66823 75214
0 1777 7 1 2 1775 78137
0 1778 5 1 1 1777
0 1779 7 1 2 1767 1778
0 1780 5 1 1 1779
0 1781 7 1 2 68750 1780
0 1782 5 1 1 1781
0 1783 7 14 2 63689 69889
0 1784 5 2 1 78140
0 1785 7 3 2 66824 77462
0 1786 7 2 2 78141 78156
0 1787 5 1 1 78159
0 1788 7 1 2 67570 78160
0 1789 5 1 1 1788
0 1790 7 1 2 1782 1789
0 1791 5 1 1 1790
0 1792 7 1 2 65642 1791
0 1793 5 1 1 1792
0 1794 7 2 2 72764 75177
0 1795 5 1 1 78161
0 1796 7 4 2 67120 70825
0 1797 5 2 1 78163
0 1798 7 2 2 73763 78164
0 1799 5 4 1 78169
0 1800 7 1 2 1795 78171
0 1801 5 1 1 1800
0 1802 7 1 2 74932 77653
0 1803 7 1 2 1801 1802
0 1804 5 1 1 1803
0 1805 7 1 2 1793 1804
0 1806 5 1 1 1805
0 1807 7 1 2 65295 1806
0 1808 5 1 1 1807
0 1809 7 7 2 68270 75869
0 1810 7 23 2 69890 65643
0 1811 7 15 2 68912 73639
0 1812 5 7 1 78205
0 1813 7 2 2 71187 78206
0 1814 5 1 1 78227
0 1815 7 1 2 78182 78228
0 1816 5 1 1 1815
0 1817 7 15 2 68521 69891
0 1818 5 1 1 78229
0 1819 7 5 2 67121 78230
0 1820 5 4 1 78244
0 1821 7 1 2 76969 78249
0 1822 5 1 1 1821
0 1823 7 2 2 70826 1822
0 1824 7 1 2 73764 78253
0 1825 5 1 1 1824
0 1826 7 1 2 1816 1825
0 1827 5 1 1 1826
0 1828 7 1 2 78175 1827
0 1829 5 1 1 1828
0 1830 7 1 2 1808 1829
0 1831 5 1 1 1830
0 1832 7 20 2 66600 69461
0 1833 5 1 1 78255
0 1834 7 14 2 64837 78256
0 1835 7 1 2 1831 78275
0 1836 5 1 1 1835
0 1837 7 1 2 1751 1836
0 1838 5 1 1 1837
0 1839 7 1 2 66342 1838
0 1840 5 1 1 1839
0 1841 7 4 2 65644 72361
0 1842 7 3 2 74424 78289
0 1843 5 1 1 78293
0 1844 7 6 2 68271 72006
0 1845 5 2 1 78296
0 1846 7 1 2 73150 78297
0 1847 5 1 1 1846
0 1848 7 1 2 1843 1847
0 1849 5 1 1 1848
0 1850 7 1 2 74759 1849
0 1851 5 1 1 1850
0 1852 7 15 2 65645 72095
0 1853 5 38 1 78304
0 1854 7 5 2 62729 78319
0 1855 5 3 1 78357
0 1856 7 1 2 73790 78358
0 1857 5 2 1 1856
0 1858 7 1 2 75215 77995
0 1859 5 1 1 1858
0 1860 7 1 2 78365 1859
0 1861 5 1 1 1860
0 1862 7 1 2 65296 1861
0 1863 5 1 1 1862
0 1864 7 4 2 72505 71512
0 1865 5 1 1 78367
0 1866 7 1 2 72406 78368
0 1867 5 1 1 1866
0 1868 7 1 2 1863 1867
0 1869 5 1 1 1868
0 1870 7 1 2 77463 1869
0 1871 5 1 1 1870
0 1872 7 1 2 1851 1871
0 1873 5 1 1 1872
0 1874 7 1 2 69892 1873
0 1875 5 1 1 1874
0 1876 7 12 2 67571 70594
0 1877 5 2 1 78371
0 1878 7 5 2 63448 75936
0 1879 5 2 1 78385
0 1880 7 1 2 78372 78386
0 1881 5 1 1 1880
0 1882 7 10 2 68751 76683
0 1883 5 2 1 78392
0 1884 7 1 2 62300 78393
0 1885 5 1 1 1884
0 1886 7 1 2 75924 1885
0 1887 5 1 1 1886
0 1888 7 1 2 73533 75504
0 1889 7 1 2 1887 1888
0 1890 5 1 1 1889
0 1891 7 1 2 1881 1890
0 1892 5 1 1 1891
0 1893 7 1 2 78127 1892
0 1894 5 1 1 1893
0 1895 7 1 2 1875 1894
0 1896 5 1 1 1895
0 1897 7 1 2 66825 1896
0 1898 5 1 1 1897
0 1899 7 18 2 65024 65297
0 1900 5 1 1 78404
0 1901 7 2 2 73799 78405
0 1902 5 1 1 78422
0 1903 7 11 2 67572 65646
0 1904 5 19 1 78424
0 1905 7 2 2 74006 78425
0 1906 5 1 1 78454
0 1907 7 1 2 72312 78455
0 1908 5 1 1 1907
0 1909 7 1 2 76494 73725
0 1910 5 1 1 1909
0 1911 7 1 2 1908 1910
0 1912 5 1 1 1911
0 1913 7 1 2 78423 1912
0 1914 5 1 1 1913
0 1915 7 1 2 1898 1914
0 1916 5 1 1 1915
0 1917 7 32 2 64612 64838
0 1918 7 36 2 61430 66601
0 1919 7 2 2 78456 78488
0 1920 7 1 2 1916 78524
0 1921 5 1 1 1920
0 1922 7 1 2 1840 1921
0 1923 5 1 1 1922
0 1924 7 1 2 67915 1923
0 1925 5 1 1 1924
0 1926 7 47 2 64839 69893
0 1927 5 1 1 78526
0 1928 7 3 2 63449 78527
0 1929 5 3 1 78573
0 1930 7 1 2 73151 78574
0 1931 5 1 1 1930
0 1932 7 47 2 69678 65025
0 1933 5 1 1 78579
0 1934 7 6 2 66826 78580
0 1935 5 3 1 78626
0 1936 7 1 2 78627 71664
0 1937 5 1 1 1936
0 1938 7 1 2 1931 1937
0 1939 5 1 1 1938
0 1940 7 1 2 61717 1939
0 1941 5 1 1 1940
0 1942 7 3 2 71464 70986
0 1943 5 3 1 78635
0 1944 7 1 2 78051 78636
0 1945 5 1 1 1944
0 1946 7 1 2 1941 1945
0 1947 5 1 1 1946
0 1948 7 1 2 67916 1947
0 1949 5 1 1 1948
0 1950 7 22 2 66827 67343
0 1951 5 2 1 78641
0 1952 7 3 2 66602 78642
0 1953 7 18 2 64840 65026
0 1954 7 18 2 62730 63055
0 1955 7 1 2 78668 78686
0 1956 7 1 2 78665 1955
0 1957 5 1 1 1956
0 1958 7 1 2 1949 1957
0 1959 5 1 1 1958
0 1960 7 1 2 70827 1959
0 1961 5 1 1 1960
0 1962 7 3 2 61718 71665
0 1963 7 15 2 67917 64841
0 1964 7 1 2 78052 78707
0 1965 7 1 2 78704 1964
0 1966 5 1 1 1965
0 1967 7 1 2 64043 1966
0 1968 7 1 2 1961 1967
0 1969 5 1 1 1968
0 1970 7 16 2 69894 74347
0 1971 5 2 1 78722
0 1972 7 3 2 64842 78723
0 1973 5 2 1 78740
0 1974 7 19 2 62484 67918
0 1975 7 2 2 78745 76990
0 1976 7 1 2 78741 78764
0 1977 5 1 1 1976
0 1978 7 1 2 68913 1977
0 1979 5 1 1 1978
0 1980 7 1 2 64613 1979
0 1981 7 1 2 1969 1980
0 1982 5 1 1 1981
0 1983 7 7 2 67919 64044
0 1984 7 10 2 67573 69462
0 1985 5 1 1 78773
0 1986 7 2 2 78766 78774
0 1987 5 1 1 78783
0 1988 7 2 2 64843 76569
0 1989 7 14 2 66828 62485
0 1990 7 1 2 66603 78787
0 1991 7 1 2 78785 1990
0 1992 7 1 2 78784 1991
0 1993 5 1 1 1992
0 1994 7 1 2 1982 1993
0 1995 5 1 1 1994
0 1996 7 1 2 66343 1995
0 1997 5 1 1 1996
0 1998 7 11 2 64614 70828
0 1999 7 4 2 64045 64844
0 2000 7 2 2 78801 78812
0 2001 7 1 2 67920 73152
0 2002 7 16 2 66829 65027
0 2003 7 1 2 78489 78818
0 2004 7 1 2 2001 2003
0 2005 7 1 2 78816 2004
0 2006 5 1 1 2005
0 2007 7 1 2 1997 2006
0 2008 5 1 1 2007
0 2009 7 1 2 72965 2008
0 2010 5 1 1 2009
0 2011 7 22 2 66604 64845
0 2012 5 2 1 78834
0 2013 7 40 2 63056 64615
0 2014 5 6 1 78858
0 2015 7 36 2 67921 69463
0 2016 5 1 1 78904
0 2017 7 2 2 78898 2016
0 2018 5 23 1 78940
0 2019 7 1 2 78835 78942
0 2020 5 1 1 2019
0 2021 7 8 2 67922 64616
0 2022 5 1 1 78965
0 2023 7 3 2 69679 78966
0 2024 7 1 2 61719 78973
0 2025 5 1 1 2024
0 2026 7 1 2 2020 2025
0 2027 5 2 1 2026
0 2028 7 1 2 66344 78976
0 2029 5 1 1 2028
0 2030 7 8 2 66605 64617
0 2031 7 7 2 64846 78978
0 2032 7 2 2 76029 78986
0 2033 5 1 1 78993
0 2034 7 1 2 2029 2033
0 2035 5 5 1 2034
0 2036 7 8 2 63690 65028
0 2037 5 1 1 79000
0 2038 7 10 2 62301 79001
0 2039 5 4 1 79008
0 2040 7 2 2 79018 78250
0 2041 5 9 1 79022
0 2042 7 1 2 75870 75009
0 2043 7 1 2 79024 2042
0 2044 7 1 2 78995 2043
0 2045 5 1 1 2044
0 2046 7 1 2 2010 2045
0 2047 5 1 1 2046
0 2048 7 1 2 73111 2047
0 2049 5 1 1 2048
0 2050 7 4 2 77325 73597
0 2051 5 3 1 79033
0 2052 7 4 2 72362 78183
0 2053 5 4 1 79040
0 2054 7 1 2 79037 79044
0 2055 5 8 1 2054
0 2056 7 3 2 72506 72966
0 2057 7 1 2 67344 79056
0 2058 7 1 2 78996 2057
0 2059 5 1 1 2058
0 2060 7 38 2 69464 64847
0 2061 7 13 2 66606 79059
0 2062 5 3 1 79097
0 2063 7 33 2 64618 69680
0 2064 7 12 2 61720 79113
0 2065 5 3 1 79146
0 2066 7 1 2 79110 79158
0 2067 5 39 1 2066
0 2068 7 3 2 70829 79161
0 2069 7 6 2 67122 75315
0 2070 5 1 1 79203
0 2071 7 1 2 66345 78767
0 2072 7 1 2 79204 2071
0 2073 7 1 2 79200 2072
0 2074 5 1 1 2073
0 2075 7 1 2 2059 2074
0 2076 5 1 1 2075
0 2077 7 1 2 67574 2076
0 2078 5 1 1 2077
0 2079 7 7 2 70830 76104
0 2080 7 11 2 67123 62731
0 2081 5 1 1 79216
0 2082 7 6 2 68522 79217
0 2083 7 11 2 67345 64046
0 2084 5 3 1 79233
0 2085 7 1 2 79234 78987
0 2086 7 1 2 79227 2085
0 2087 7 1 2 79209 2086
0 2088 5 1 1 2087
0 2089 7 1 2 2078 2088
0 2090 5 1 1 2089
0 2091 7 1 2 66830 2090
0 2092 5 1 1 2091
0 2093 7 27 2 66346 61979
0 2094 7 2 2 77430 79247
0 2095 7 8 2 67923 63691
0 2096 7 2 2 62732 79276
0 2097 7 6 2 61721 68914
0 2098 7 1 2 78457 79286
0 2099 7 1 2 79284 2098
0 2100 7 1 2 79274 2099
0 2101 5 1 1 2100
0 2102 7 1 2 2092 2101
0 2103 5 1 1 2102
0 2104 7 1 2 79048 2103
0 2105 5 1 1 2104
0 2106 7 10 2 65029 65647
0 2107 7 3 2 68523 79292
0 2108 7 1 2 75261 79302
0 2109 5 1 1 2108
0 2110 7 5 2 68272 77124
0 2111 5 1 1 79305
0 2112 7 1 2 79306 78643
0 2113 5 1 1 2112
0 2114 7 1 2 2109 2113
0 2115 5 1 1 2114
0 2116 7 1 2 71144 2115
0 2117 5 1 1 2116
0 2118 7 1 2 79019 78120
0 2119 5 2 1 2118
0 2120 7 1 2 73173 79310
0 2121 5 1 1 2120
0 2122 7 1 2 78245 74425
0 2123 5 1 1 2122
0 2124 7 1 2 2121 2123
0 2125 5 1 1 2124
0 2126 7 1 2 76021 2125
0 2127 5 1 1 2126
0 2128 7 1 2 2117 2127
0 2129 5 1 1 2128
0 2130 7 1 2 68752 2129
0 2131 5 1 1 2130
0 2132 7 2 2 77996 77654
0 2133 5 1 1 79312
0 2134 7 1 2 77464 75216
0 2135 7 1 2 79313 2134
0 2136 5 1 1 2135
0 2137 7 1 2 2131 2136
0 2138 5 1 1 2137
0 2139 7 1 2 65298 2138
0 2140 5 1 1 2139
0 2141 7 3 2 68273 78644
0 2142 7 5 2 67575 72744
0 2143 5 1 1 79317
0 2144 7 3 2 78184 73640
0 2145 7 1 2 79318 79322
0 2146 5 1 1 2145
0 2147 7 1 2 72774 78254
0 2148 5 1 1 2147
0 2149 7 1 2 2146 2148
0 2150 5 1 1 2149
0 2151 7 1 2 79314 2150
0 2152 5 1 1 2151
0 2153 7 1 2 2140 2152
0 2154 5 1 1 2153
0 2155 7 4 2 78458 76543
0 2156 7 1 2 63057 79325
0 2157 7 1 2 2154 2156
0 2158 5 1 1 2157
0 2159 7 1 2 69276 2158
0 2160 7 1 2 2105 2159
0 2161 7 1 2 2049 2160
0 2162 7 1 2 1925 2161
0 2163 5 1 1 2162
0 2164 7 1 2 1557 2163
0 2165 5 1 1 2164
0 2166 7 1 2 63217 2165
0 2167 5 1 1 2166
0 2168 7 56 2 64428 69465
0 2169 7 5 2 69895 79329
0 2170 7 8 2 72007 73930
0 2171 5 3 1 79390
0 2172 7 1 2 76613 79391
0 2173 5 1 1 2172
0 2174 7 1 2 74476 2173
0 2175 5 1 1 2174
0 2176 7 1 2 76811 2175
0 2177 5 1 1 2176
0 2178 7 5 2 62302 73186
0 2179 7 1 2 74348 79401
0 2180 5 1 1 2179
0 2181 7 1 2 75793 2180
0 2182 5 1 1 2181
0 2183 7 1 2 71145 2182
0 2184 5 1 1 2183
0 2185 7 1 2 75755 72419
0 2186 5 1 1 2185
0 2187 7 1 2 2184 2186
0 2188 5 1 1 2187
0 2189 7 1 2 62486 2188
0 2190 5 1 1 2189
0 2191 7 1 2 2177 2190
0 2192 5 1 1 2191
0 2193 7 1 2 79385 2192
0 2194 5 1 1 2193
0 2195 7 2 2 65648 72927
0 2196 7 54 2 69277 64619
0 2197 7 6 2 65030 79408
0 2198 7 12 2 67124 68753
0 2199 5 1 1 79468
0 2200 7 2 2 74299 79469
0 2201 7 1 2 79462 79480
0 2202 7 1 2 79406 2201
0 2203 5 1 1 2202
0 2204 7 1 2 2194 2203
0 2205 5 1 1 2204
0 2206 7 1 2 65299 2205
0 2207 5 1 1 2206
0 2208 7 2 2 76409 71618
0 2209 7 1 2 61980 79482
0 2210 5 1 1 2209
0 2211 7 1 2 62303 76417
0 2212 5 1 1 2211
0 2213 7 1 2 2210 2212
0 2214 5 2 1 2213
0 2215 7 8 2 62487 68915
0 2216 5 2 1 79486
0 2217 7 1 2 79484 79487
0 2218 5 1 1 2217
0 2219 7 11 2 67346 71513
0 2220 5 13 1 79496
0 2221 7 1 2 76812 79497
0 2222 5 1 1 2221
0 2223 7 1 2 76414 2222
0 2224 5 1 1 2223
0 2225 7 1 2 72008 2224
0 2226 5 1 1 2225
0 2227 7 1 2 62733 2226
0 2228 7 1 2 2218 2227
0 2229 5 1 1 2228
0 2230 7 1 2 78022 79485
0 2231 5 1 1 2230
0 2232 7 5 2 72258 75279
0 2233 7 1 2 77512 79520
0 2234 5 1 1 2233
0 2235 7 1 2 67576 2234
0 2236 7 1 2 2231 2235
0 2237 5 1 1 2236
0 2238 7 14 2 64429 69896
0 2239 7 11 2 69466 70208
0 2240 7 2 2 79525 79539
0 2241 7 1 2 2237 79550
0 2242 7 1 2 2229 2241
0 2243 5 1 1 2242
0 2244 7 1 2 2207 2243
0 2245 5 1 1 2244
0 2246 7 1 2 68524 2245
0 2247 5 1 1 2246
0 2248 7 5 2 62734 76927
0 2249 5 1 1 79552
0 2250 7 3 2 77022 79553
0 2251 5 1 1 79557
0 2252 7 4 2 76307 76876
0 2253 5 1 1 79560
0 2254 7 1 2 67577 75280
0 2255 7 1 2 79561 2254
0 2256 5 1 1 2255
0 2257 7 1 2 2251 2256
0 2258 5 1 1 2257
0 2259 7 1 2 62488 2258
0 2260 5 1 1 2259
0 2261 7 2 2 77326 73844
0 2262 7 6 2 62735 73958
0 2263 5 1 1 79566
0 2264 7 1 2 79564 79567
0 2265 5 1 1 2264
0 2266 7 1 2 2260 2265
0 2267 5 1 1 2266
0 2268 7 1 2 75756 2267
0 2269 5 1 1 2268
0 2270 7 11 2 67125 69897
0 2271 7 1 2 65300 73176
0 2272 5 1 1 2271
0 2273 7 1 2 72689 78207
0 2274 5 2 1 2273
0 2275 7 1 2 2272 79583
0 2276 5 1 1 2275
0 2277 7 1 2 79572 2276
0 2278 5 1 1 2277
0 2279 7 1 2 62304 77033
0 2280 5 1 1 2279
0 2281 7 1 2 2278 2280
0 2282 5 1 1 2281
0 2283 7 1 2 70595 2282
0 2284 5 1 1 2283
0 2285 7 1 2 1047 76870
0 2286 5 1 1 2285
0 2287 7 1 2 77142 2286
0 2288 5 1 1 2287
0 2289 7 1 2 2284 2288
0 2290 5 1 1 2289
0 2291 7 1 2 63892 2290
0 2292 5 1 1 2291
0 2293 7 1 2 67578 77368
0 2294 5 1 1 2293
0 2295 7 2 2 62489 78435
0 2296 5 1 1 79585
0 2297 7 7 2 62305 65031
0 2298 5 1 1 79587
0 2299 7 1 2 79586 79588
0 2300 5 1 1 2299
0 2301 7 1 2 2294 2300
0 2302 5 1 1 2301
0 2303 7 1 2 61981 2302
0 2304 5 1 1 2303
0 2305 7 20 2 69898 70209
0 2306 5 1 1 79594
0 2307 7 2 2 67126 79595
0 2308 5 1 1 79614
0 2309 7 1 2 71514 73177
0 2310 5 1 1 2309
0 2311 7 1 2 72238 2310
0 2312 5 1 1 2311
0 2313 7 1 2 79615 2312
0 2314 5 1 1 2313
0 2315 7 1 2 2304 2314
0 2316 7 1 2 2292 2315
0 2317 5 1 1 2316
0 2318 7 1 2 63450 2317
0 2319 5 1 1 2318
0 2320 7 8 2 64047 76570
0 2321 5 1 1 79616
0 2322 7 9 2 71289 71716
0 2323 5 1 1 79624
0 2324 7 2 2 79617 79625
0 2325 7 1 2 77160 79633
0 2326 5 1 1 2325
0 2327 7 1 2 62306 73795
0 2328 5 1 1 2327
0 2329 7 1 2 75021 73871
0 2330 5 1 1 2329
0 2331 7 1 2 2328 2330
0 2332 5 1 1 2331
0 2333 7 1 2 69899 2332
0 2334 5 1 1 2333
0 2335 7 1 2 2326 2334
0 2336 7 1 2 2319 2335
0 2337 5 1 1 2336
0 2338 7 1 2 63692 2337
0 2339 5 1 1 2338
0 2340 7 1 2 2269 2339
0 2341 5 1 1 2340
0 2342 7 1 2 79330 2341
0 2343 5 1 1 2342
0 2344 7 1 2 2247 2343
0 2345 5 1 1 2344
0 2346 7 1 2 69681 2345
0 2347 5 1 1 2346
0 2348 7 13 2 64848 79409
0 2349 7 3 2 68274 74529
0 2350 5 1 1 79648
0 2351 7 1 2 75505 78394
0 2352 5 1 1 2351
0 2353 7 1 2 2350 2352
0 2354 5 1 1 2353
0 2355 7 1 2 62307 2354
0 2356 5 1 1 2355
0 2357 7 1 2 850 75300
0 2358 5 1 1 2357
0 2359 7 1 2 75913 2358
0 2360 5 1 1 2359
0 2361 7 1 2 2356 2360
0 2362 5 1 1 2361
0 2363 7 1 2 65032 2362
0 2364 5 1 1 2363
0 2365 7 1 2 74831 78402
0 2366 5 1 1 2365
0 2367 7 1 2 69900 77465
0 2368 7 1 2 2366 2367
0 2369 5 1 1 2368
0 2370 7 1 2 2364 2369
0 2371 5 1 1 2370
0 2372 7 1 2 72009 2371
0 2373 5 1 1 2372
0 2374 7 10 2 68916 71188
0 2375 7 6 2 69901 73054
0 2376 7 1 2 68275 79661
0 2377 7 1 2 79651 2376
0 2378 5 1 1 2377
0 2379 7 1 2 2373 2378
0 2380 5 1 1 2379
0 2381 7 1 2 62736 2380
0 2382 5 1 1 2381
0 2383 7 1 2 2037 78251
0 2384 5 5 1 2383
0 2385 7 1 2 79667 78294
0 2386 5 1 1 2385
0 2387 7 1 2 2382 2386
0 2388 5 1 1 2387
0 2389 7 1 2 66831 2388
0 2390 5 1 1 2389
0 2391 7 2 2 67127 74282
0 2392 7 13 2 64048 65649
0 2393 5 5 1 79674
0 2394 7 11 2 62490 68754
0 2395 5 2 1 79692
0 2396 7 1 2 79675 79693
0 2397 5 2 1 2396
0 2398 7 1 2 68525 79705
0 2399 5 1 1 2398
0 2400 7 1 2 79672 2399
0 2401 5 1 1 2400
0 2402 7 1 2 68276 74832
0 2403 7 1 2 77776 2402
0 2404 5 1 1 2403
0 2405 7 1 2 2401 2404
0 2406 5 1 1 2405
0 2407 7 1 2 78406 74461
0 2408 7 1 2 2406 2407
0 2409 5 1 1 2408
0 2410 7 1 2 2390 2409
0 2411 5 1 1 2410
0 2412 7 1 2 79635 2411
0 2413 5 1 1 2412
0 2414 7 1 2 2347 2413
0 2415 5 1 1 2414
0 2416 7 1 2 61722 2415
0 2417 5 1 1 2416
0 2418 7 4 2 66832 71795
0 2419 5 4 1 79707
0 2420 7 1 2 76635 79711
0 2421 5 9 1 2420
0 2422 7 2 2 71146 71559
0 2423 5 1 1 79724
0 2424 7 1 2 72433 2423
0 2425 5 1 1 2424
0 2426 7 2 2 79331 77110
0 2427 7 1 2 63451 79726
0 2428 7 1 2 2425 2427
0 2429 5 1 1 2428
0 2430 7 2 2 72010 72382
0 2431 5 1 1 79728
0 2432 7 1 2 77863 2431
0 2433 5 1 1 2432
0 2434 7 11 2 66607 68277
0 2435 7 18 2 64620 65033
0 2436 7 4 2 69278 79741
0 2437 7 1 2 79730 79759
0 2438 7 1 2 2433 2437
0 2439 5 1 1 2438
0 2440 7 1 2 2429 2439
0 2441 5 1 1 2440
0 2442 7 1 2 69682 2441
0 2443 5 1 1 2442
0 2444 7 21 2 61723 68278
0 2445 7 5 2 78669 79410
0 2446 7 2 2 79763 79784
0 2447 7 1 2 79789 79725
0 2448 5 1 1 2447
0 2449 7 1 2 2443 2448
0 2450 5 1 1 2449
0 2451 7 1 2 79715 2450
0 2452 5 1 1 2451
0 2453 7 11 2 66608 69279
0 2454 7 9 2 68917 64849
0 2455 7 1 2 79802 76532
0 2456 5 1 1 2455
0 2457 7 4 2 72011 73598
0 2458 7 9 2 66833 68526
0 2459 7 2 2 79815 75045
0 2460 7 1 2 79811 79824
0 2461 5 1 1 2460
0 2462 7 1 2 2456 2461
0 2463 5 1 1 2462
0 2464 7 1 2 62491 2463
0 2465 5 1 1 2464
0 2466 7 9 2 68279 64049
0 2467 7 5 2 70831 79826
0 2468 7 3 2 68527 77387
0 2469 5 1 1 79840
0 2470 7 5 2 61982 75068
0 2471 7 1 2 75061 79843
0 2472 5 1 1 2471
0 2473 7 1 2 2469 2472
0 2474 5 1 1 2473
0 2475 7 1 2 62308 2474
0 2476 5 1 1 2475
0 2477 7 14 2 63693 69683
0 2478 7 9 2 63893 77431
0 2479 5 1 1 79862
0 2480 7 2 2 66834 2479
0 2481 5 4 1 79871
0 2482 7 1 2 79848 79872
0 2483 5 1 1 2482
0 2484 7 1 2 2476 2483
0 2485 5 1 1 2484
0 2486 7 1 2 70210 2485
0 2487 5 1 1 2486
0 2488 7 1 2 174 77730
0 2489 5 1 1 2488
0 2490 7 4 2 67128 69684
0 2491 7 1 2 61983 79877
0 2492 7 1 2 2489 2491
0 2493 5 1 1 2492
0 2494 7 1 2 2487 2493
0 2495 5 1 1 2494
0 2496 7 1 2 79835 2495
0 2497 5 1 1 2496
0 2498 7 1 2 2465 2497
0 2499 5 1 1 2498
0 2500 7 1 2 65034 2499
0 2501 5 1 1 2500
0 2502 7 2 2 78528 74648
0 2503 7 1 2 73800 79488
0 2504 7 1 2 79881 2503
0 2505 5 1 1 2504
0 2506 7 1 2 2501 2505
0 2507 5 1 1 2506
0 2508 7 1 2 70596 2507
0 2509 5 1 1 2508
0 2510 7 1 2 76619 73972
0 2511 5 1 1 2510
0 2512 7 1 2 76636 2511
0 2513 5 1 1 2512
0 2514 7 1 2 62309 2513
0 2515 5 1 1 2514
0 2516 7 7 2 62310 71290
0 2517 5 26 1 79883
0 2518 7 7 2 65301 79890
0 2519 7 1 2 74447 79916
0 2520 5 1 1 2519
0 2521 7 1 2 2515 2520
0 2522 5 1 1 2521
0 2523 7 6 2 68280 65650
0 2524 5 2 1 79923
0 2525 7 1 2 78581 79924
0 2526 7 1 2 2522 2525
0 2527 5 1 1 2526
0 2528 7 1 2 2509 2527
0 2529 5 1 1 2528
0 2530 7 1 2 64621 2529
0 2531 5 1 1 2530
0 2532 7 12 2 64850 65302
0 2533 7 3 2 79293 79931
0 2534 7 2 2 72928 79943
0 2535 7 17 2 66835 67129
0 2536 7 7 2 68528 69467
0 2537 7 3 2 79965 75432
0 2538 7 2 2 79948 79972
0 2539 7 1 2 79946 79975
0 2540 5 1 1 2539
0 2541 7 1 2 2531 2540
0 2542 5 1 1 2541
0 2543 7 1 2 79791 2542
0 2544 5 1 1 2543
0 2545 7 1 2 2452 2544
0 2546 7 1 2 2417 2545
0 2547 5 1 1 2546
0 2548 7 1 2 76105 2547
0 2549 5 1 1 2548
0 2550 7 1 2 75638 74944
0 2551 5 1 1 2550
0 2552 7 6 2 70832 71108
0 2553 5 1 1 79977
0 2554 7 1 2 62492 2553
0 2555 5 1 1 2554
0 2556 7 5 2 65651 74760
0 2557 7 1 2 1456 79983
0 2558 7 1 2 2555 2557
0 2559 5 1 1 2558
0 2560 7 1 2 2551 2559
0 2561 5 1 1 2560
0 2562 7 1 2 78859 2561
0 2563 5 1 1 2562
0 2564 7 1 2 74912 75010
0 2565 5 1 1 2564
0 2566 7 1 2 75209 73750
0 2567 5 1 1 2566
0 2568 7 1 2 2565 2567
0 2569 5 1 1 2568
0 2570 7 1 2 78905 2569
0 2571 5 1 1 2570
0 2572 7 1 2 2563 2571
0 2573 5 1 1 2572
0 2574 7 1 2 68755 2573
0 2575 5 1 1 2574
0 2576 7 7 2 73370 75740
0 2577 5 21 1 79988
0 2578 7 3 2 68529 79995
0 2579 5 1 1 80016
0 2580 7 1 2 72953 2579
0 2581 5 2 1 2580
0 2582 7 17 2 67924 68281
0 2583 7 17 2 69468 65912
0 2584 7 7 2 68918 80038
0 2585 7 1 2 80021 80055
0 2586 7 1 2 80019 2585
0 2587 5 1 1 2586
0 2588 7 1 2 2575 2587
0 2589 5 1 1 2588
0 2590 7 1 2 66836 2589
0 2591 5 1 1 2590
0 2592 7 11 2 62493 70833
0 2593 5 3 1 80062
0 2594 7 6 2 65652 71147
0 2595 7 1 2 80063 80076
0 2596 5 1 1 2595
0 2597 7 1 2 61984 75011
0 2598 5 1 1 2597
0 2599 7 1 2 2596 2598
0 2600 5 1 1 2599
0 2601 7 12 2 67130 67925
0 2602 7 1 2 80082 79973
0 2603 7 1 2 2600 2602
0 2604 5 1 1 2603
0 2605 7 1 2 2591 2604
0 2606 5 1 1 2605
0 2607 7 1 2 69685 2606
0 2608 5 1 1 2607
0 2609 7 10 2 68919 69469
0 2610 5 1 1 80094
0 2611 7 5 2 65913 78906
0 2612 5 2 1 80104
0 2613 7 9 2 63058 68920
0 2614 5 1 1 80111
0 2615 7 1 2 80109 2614
0 2616 5 1 1 2615
0 2617 7 2 2 2610 2616
0 2618 7 1 2 62737 80120
0 2619 5 1 1 2618
0 2620 7 23 2 67579 63059
0 2621 7 9 2 64050 64622
0 2622 7 1 2 80122 80145
0 2623 5 2 1 2622
0 2624 7 1 2 2619 80154
0 2625 5 2 1 2624
0 2626 7 1 2 62311 73892
0 2627 5 1 1 2626
0 2628 7 1 2 72939 73187
0 2629 5 1 1 2628
0 2630 7 1 2 74895 2629
0 2631 7 1 2 2627 2630
0 2632 5 2 1 2631
0 2633 7 1 2 80156 80158
0 2634 5 1 1 2633
0 2635 7 14 2 68921 64623
0 2636 7 2 2 76308 80160
0 2637 7 2 2 77291 80123
0 2638 7 1 2 80174 80176
0 2639 5 1 1 2638
0 2640 7 1 2 2634 2639
0 2641 5 1 1 2640
0 2642 7 1 2 62494 2641
0 2643 5 1 1 2642
0 2644 7 3 2 65914 71560
0 2645 7 11 2 64051 69470
0 2646 7 22 2 62738 67926
0 2647 7 2 2 80192 74877
0 2648 7 1 2 80181 80214
0 2649 7 1 2 80178 2648
0 2650 5 1 1 2649
0 2651 7 1 2 2643 2650
0 2652 5 1 1 2651
0 2653 7 1 2 77079 2652
0 2654 5 1 1 2653
0 2655 7 1 2 2608 2654
0 2656 5 1 1 2655
0 2657 7 1 2 65303 2656
0 2658 5 1 1 2657
0 2659 7 14 2 67580 67927
0 2660 5 1 1 80216
0 2661 7 6 2 67581 64624
0 2662 5 1 1 80230
0 2663 7 1 2 2662 80110
0 2664 5 1 1 2663
0 2665 7 2 2 2660 2664
0 2666 7 1 2 73801 71515
0 2667 7 1 2 80236 2666
0 2668 5 1 1 2667
0 2669 7 12 2 69471 70834
0 2670 7 3 2 73188 80238
0 2671 7 1 2 75871 79277
0 2672 7 1 2 80250 2671
0 2673 5 1 1 2672
0 2674 7 1 2 2668 2673
0 2675 5 1 1 2674
0 2676 7 1 2 62495 2675
0 2677 5 1 1 2676
0 2678 7 2 2 70835 78860
0 2679 7 1 2 73931 76630
0 2680 7 1 2 80253 2679
0 2681 5 1 1 2680
0 2682 7 1 2 2677 2681
0 2683 5 1 1 2682
0 2684 7 1 2 64052 2683
0 2685 5 1 1 2684
0 2686 7 9 2 64625 65653
0 2687 7 2 2 78687 80255
0 2688 5 1 1 80264
0 2689 7 8 2 61985 68756
0 2690 5 1 1 80266
0 2691 7 3 2 68922 80267
0 2692 7 1 2 80274 75316
0 2693 7 1 2 80265 2692
0 2694 5 1 1 2693
0 2695 7 1 2 2685 2694
0 2696 5 1 1 2695
0 2697 7 1 2 64851 77543
0 2698 7 1 2 2696 2697
0 2699 5 1 1 2698
0 2700 7 11 2 61986 70597
0 2701 5 1 1 80277
0 2702 7 24 2 64852 70211
0 2703 7 1 2 73282 80288
0 2704 7 3 2 80278 2703
0 2705 7 1 2 68530 80312
0 2706 5 1 1 2705
0 2707 7 3 2 64853 72437
0 2708 7 1 2 74448 79694
0 2709 7 1 2 80315 2708
0 2710 5 1 1 2709
0 2711 7 1 2 2706 2710
0 2712 5 1 1 2711
0 2713 7 1 2 80157 2712
0 2714 5 1 1 2713
0 2715 7 12 2 64626 70598
0 2716 7 4 2 63060 71109
0 2717 7 2 2 80318 80330
0 2718 5 1 1 80334
0 2719 7 1 2 70836 2718
0 2720 5 1 1 2719
0 2721 7 2 2 78907 76595
0 2722 5 1 1 80336
0 2723 7 1 2 65915 2722
0 2724 5 1 1 2723
0 2725 7 1 2 79825 2724
0 2726 7 1 2 2720 2725
0 2727 5 1 1 2726
0 2728 7 1 2 2714 2727
0 2729 5 1 1 2728
0 2730 7 1 2 67131 2729
0 2731 5 1 1 2730
0 2732 7 1 2 69902 2731
0 2733 7 1 2 2699 2732
0 2734 7 1 2 2658 2733
0 2735 5 1 1 2734
0 2736 7 15 2 69686 70837
0 2737 7 3 2 69472 80022
0 2738 7 4 2 72967 73112
0 2739 5 1 1 80356
0 2740 7 3 2 70599 74761
0 2741 7 1 2 73599 80360
0 2742 5 2 1 2741
0 2743 7 1 2 2739 80363
0 2744 5 1 1 2743
0 2745 7 2 2 80353 2744
0 2746 5 1 1 80365
0 2747 7 3 2 77848 74672
0 2748 5 1 1 80367
0 2749 7 2 2 65304 80368
0 2750 5 2 1 80370
0 2751 7 1 2 80364 80372
0 2752 5 2 1 2751
0 2753 7 1 2 64627 75569
0 2754 7 1 2 80374 2753
0 2755 5 1 1 2754
0 2756 7 1 2 2746 2755
0 2757 5 1 1 2756
0 2758 7 1 2 80338 2757
0 2759 5 1 1 2758
0 2760 7 3 2 63061 78459
0 2761 7 10 2 70212 73189
0 2762 7 4 2 71796 80379
0 2763 5 2 1 80389
0 2764 7 1 2 68282 80393
0 2765 5 1 1 2764
0 2766 7 6 2 77914 2765
0 2767 5 1 1 80395
0 2768 7 2 2 61987 80396
0 2769 5 1 1 80401
0 2770 7 1 2 80376 80402
0 2771 5 1 1 2770
0 2772 7 1 2 2759 2771
0 2773 5 1 1 2772
0 2774 7 1 2 67582 2773
0 2775 5 1 1 2774
0 2776 7 12 2 63062 63452
0 2777 7 4 2 64628 80403
0 2778 7 4 2 70838 71561
0 2779 5 1 1 80419
0 2780 7 1 2 70213 75201
0 2781 7 2 2 80420 2780
0 2782 7 1 2 80415 80423
0 2783 5 1 1 2782
0 2784 7 3 2 67928 80039
0 2785 7 1 2 80397 80425
0 2786 5 1 1 2785
0 2787 7 1 2 2783 2786
0 2788 5 1 1 2787
0 2789 7 1 2 62739 2788
0 2790 5 1 1 2789
0 2791 7 4 2 68283 74563
0 2792 5 1 1 80428
0 2793 7 13 2 62312 67929
0 2794 7 1 2 80432 80251
0 2795 7 1 2 80429 2794
0 2796 5 1 1 2795
0 2797 7 1 2 2790 2796
0 2798 5 1 1 2797
0 2799 7 1 2 77080 2798
0 2800 5 1 1 2799
0 2801 7 1 2 2775 2800
0 2802 5 1 1 2801
0 2803 7 1 2 64053 2802
0 2804 5 1 1 2803
0 2805 7 1 2 80377 80398
0 2806 5 1 1 2805
0 2807 7 5 2 65305 77807
0 2808 7 3 2 67930 80445
0 2809 7 8 2 68757 69473
0 2810 7 3 2 68531 80453
0 2811 7 1 2 79878 80461
0 2812 7 1 2 80450 2811
0 2813 5 1 1 2812
0 2814 7 1 2 2806 2813
0 2815 5 1 1 2814
0 2816 7 1 2 61988 2815
0 2817 5 1 1 2816
0 2818 7 1 2 80339 80366
0 2819 5 1 1 2818
0 2820 7 1 2 2817 2819
0 2821 5 1 1 2820
0 2822 7 1 2 71121 2821
0 2823 5 1 1 2822
0 2824 7 1 2 2804 2823
0 2825 5 1 1 2824
0 2826 7 1 2 62496 2825
0 2827 5 1 1 2826
0 2828 7 14 2 63694 64054
0 2829 7 2 2 80433 75232
0 2830 7 10 2 63453 69474
0 2831 7 3 2 64854 80480
0 2832 7 1 2 80179 80490
0 2833 7 1 2 80478 2832
0 2834 5 1 1 2833
0 2835 7 10 2 70839 71717
0 2836 7 7 2 63063 69687
0 2837 7 1 2 74300 80503
0 2838 7 1 2 80231 2837
0 2839 7 1 2 80493 2838
0 2840 5 1 1 2839
0 2841 7 1 2 2834 2840
0 2842 5 1 1 2841
0 2843 7 1 2 80464 2842
0 2844 5 1 1 2843
0 2845 7 1 2 65035 2844
0 2846 7 1 2 2827 2845
0 2847 5 1 1 2846
0 2848 7 1 2 2735 2847
0 2849 5 1 1 2848
0 2850 7 6 2 65306 78460
0 2851 7 6 2 63695 65916
0 2852 7 1 2 80404 80516
0 2853 7 1 2 80510 2852
0 2854 7 2 2 67583 71643
0 2855 5 2 1 80522
0 2856 7 2 2 75843 77608
0 2857 7 1 2 80523 80526
0 2858 7 1 2 2853 2857
0 2859 5 1 1 2858
0 2860 7 1 2 2849 2859
0 2861 5 1 1 2860
0 2862 7 1 2 66347 2861
0 2863 5 1 1 2862
0 2864 7 6 2 64055 74170
0 2865 5 6 1 80528
0 2866 7 5 2 65307 80534
0 2867 5 8 1 80540
0 2868 7 9 2 71753 80545
0 2869 7 4 2 69688 74762
0 2870 7 1 2 77046 77674
0 2871 5 32 1 2870
0 2872 7 1 2 80562 80566
0 2873 7 1 2 80553 2872
0 2874 5 1 1 2873
0 2875 7 3 2 69903 79803
0 2876 7 1 2 80598 71612
0 2877 7 1 2 79844 2876
0 2878 5 1 1 2877
0 2879 7 1 2 2874 2878
0 2880 5 1 1 2879
0 2881 7 1 2 67931 2880
0 2882 5 1 1 2881
0 2883 7 11 2 63064 68758
0 2884 7 8 2 68532 79949
0 2885 7 1 2 80601 80612
0 2886 7 1 2 79947 2885
0 2887 5 1 1 2886
0 2888 7 1 2 2882 2887
0 2889 5 1 1 2888
0 2890 7 15 2 61431 68284
0 2891 7 1 2 64629 80620
0 2892 7 1 2 2889 2891
0 2893 5 1 1 2892
0 2894 7 1 2 66609 2893
0 2895 7 1 2 2863 2894
0 2896 5 1 1 2895
0 2897 7 3 2 61432 80023
0 2898 7 1 2 80567 80635
0 2899 5 1 1 2898
0 2900 7 3 2 66348 78645
0 2901 7 1 2 78185 80602
0 2902 7 1 2 80638 2901
0 2903 5 1 1 2902
0 2904 7 1 2 2899 2903
0 2905 5 1 1 2904
0 2906 7 1 2 65308 2905
0 2907 5 1 1 2906
0 2908 7 16 2 67347 63065
0 2909 7 4 2 66349 80641
0 2910 7 3 2 70214 78819
0 2911 7 2 2 73190 80661
0 2912 7 1 2 80657 80664
0 2913 5 1 1 2912
0 2914 7 1 2 2907 2913
0 2915 5 1 1 2914
0 2916 7 1 2 74763 2915
0 2917 5 1 1 2916
0 2918 7 9 2 66350 78746
0 2919 7 10 2 69904 71718
0 2920 7 2 2 76533 80675
0 2921 7 1 2 80666 80685
0 2922 5 1 1 2921
0 2923 7 1 2 2917 2922
0 2924 5 1 1 2923
0 2925 7 1 2 73534 2924
0 2926 5 1 1 2925
0 2927 7 9 2 68759 69905
0 2928 7 2 2 68285 80687
0 2929 5 1 1 80696
0 2930 7 1 2 80697 80658
0 2931 5 1 1 2930
0 2932 7 17 2 63454 65036
0 2933 5 4 1 80698
0 2934 7 2 2 68533 76030
0 2935 5 1 1 80719
0 2936 7 1 2 80699 80720
0 2937 5 1 1 2936
0 2938 7 1 2 2931 2937
0 2939 5 1 1 2938
0 2940 7 1 2 66837 2939
0 2941 5 1 1 2940
0 2942 7 15 2 66351 62497
0 2943 7 14 2 63066 68286
0 2944 7 2 2 80721 80736
0 2945 7 6 2 63894 65037
0 2946 7 1 2 72968 80752
0 2947 7 1 2 80750 2946
0 2948 5 1 1 2947
0 2949 7 1 2 2941 2948
0 2950 5 1 1 2949
0 2951 7 1 2 73055 2950
0 2952 5 1 1 2951
0 2953 7 7 2 65654 72969
0 2954 5 1 1 80758
0 2955 7 11 2 68760 65038
0 2956 7 2 2 70215 80765
0 2957 7 1 2 80751 80776
0 2958 7 1 2 80759 2957
0 2959 5 1 1 2958
0 2960 7 1 2 2952 2959
0 2961 5 1 1 2960
0 2962 7 1 2 67584 2961
0 2963 5 1 1 2962
0 2964 7 1 2 2926 2963
0 2965 5 1 1 2964
0 2966 7 1 2 64056 2965
0 2967 5 1 1 2966
0 2968 7 20 2 61433 67585
0 2969 7 11 2 67932 68534
0 2970 7 1 2 80778 80798
0 2971 7 1 2 80568 2970
0 2972 5 1 1 2971
0 2973 7 2 2 71644 80766
0 2974 7 5 2 66352 78688
0 2975 5 1 1 80811
0 2976 7 1 2 77593 80812
0 2977 7 1 2 80809 2976
0 2978 5 1 1 2977
0 2979 7 1 2 2972 2978
0 2980 5 1 1 2979
0 2981 7 1 2 70216 2980
0 2982 5 1 1 2981
0 2983 7 2 2 65039 73056
0 2984 7 10 2 63067 63696
0 2985 7 3 2 62740 80818
0 2986 7 1 2 75281 80722
0 2987 7 1 2 80828 2986
0 2988 7 1 2 80816 2987
0 2989 5 1 1 2988
0 2990 7 1 2 2982 2989
0 2991 5 1 1 2990
0 2992 7 1 2 67132 2991
0 2993 5 1 1 2992
0 2994 7 11 2 66353 62313
0 2995 7 2 2 72910 80831
0 2996 7 11 2 63068 68535
0 2997 7 9 2 68923 65040
0 2998 7 1 2 80844 80855
0 2999 7 1 2 80842 2998
0 3000 7 1 2 73113 2999
0 3001 5 1 1 3000
0 3002 7 1 2 2993 3001
0 3003 5 1 1 3002
0 3004 7 1 2 68287 3003
0 3005 5 1 1 3004
0 3006 7 16 2 68536 65041
0 3007 7 3 2 66354 75022
0 3008 7 1 2 80864 80880
0 3009 7 2 2 62498 78689
0 3010 7 2 2 71645 72363
0 3011 7 1 2 80883 80885
0 3012 7 1 2 3008 3011
0 3013 5 1 1 3012
0 3014 7 1 2 3005 3013
0 3015 7 1 2 2967 3014
0 3016 5 1 1 3015
0 3017 7 1 2 64630 3016
0 3018 5 1 1 3017
0 3019 7 4 2 63697 72364
0 3020 5 2 1 80887
0 3021 7 1 2 73999 72487
0 3022 5 1 1 3021
0 3023 7 1 2 67348 3022
0 3024 5 1 1 3023
0 3025 7 1 2 80891 3024
0 3026 5 1 1 3025
0 3027 7 1 2 72507 3026
0 3028 5 1 1 3027
0 3029 7 7 2 67133 74573
0 3030 5 1 1 80893
0 3031 7 1 2 75639 80894
0 3032 5 2 1 3031
0 3033 7 1 2 3028 80900
0 3034 5 1 1 3033
0 3035 7 12 2 68288 69475
0 3036 7 3 2 69906 80902
0 3037 7 27 2 66355 67586
0 3038 7 10 2 66838 67933
0 3039 7 2 2 80917 80944
0 3040 7 1 2 80914 80954
0 3041 7 1 2 3034 3040
0 3042 5 1 1 3041
0 3043 7 1 2 3018 3042
0 3044 5 1 1 3043
0 3045 7 1 2 64855 3044
0 3046 5 1 1 3045
0 3047 7 47 2 66356 67934
0 3048 5 3 1 80956
0 3049 7 8 2 69689 80957
0 3050 7 6 2 65042 76684
0 3051 7 2 2 79976 81014
0 3052 5 1 1 81020
0 3053 7 1 2 72929 81021
0 3054 5 1 1 3053
0 3055 7 7 2 67587 69907
0 3056 5 2 1 81022
0 3057 7 3 2 66839 81023
0 3058 5 2 1 81031
0 3059 7 23 2 68289 65043
0 3060 5 4 1 81036
0 3061 7 3 2 61989 81037
0 3062 5 2 1 81063
0 3063 7 1 2 81034 81066
0 3064 5 1 1 3063
0 3065 7 6 2 63895 64631
0 3066 7 2 2 80465 81068
0 3067 7 1 2 80494 77432
0 3068 7 1 2 81074 3067
0 3069 7 1 2 3064 3068
0 3070 5 1 1 3069
0 3071 7 1 2 3054 3070
0 3072 5 1 1 3071
0 3073 7 1 2 81006 3072
0 3074 5 1 1 3073
0 3075 7 1 2 61724 3074
0 3076 7 1 2 3046 3075
0 3077 5 1 1 3076
0 3078 7 1 2 69280 3077
0 3079 7 1 2 2896 3078
0 3080 5 1 1 3079
0 3081 7 40 2 64430 77217
0 3082 5 3 1 81076
0 3083 7 14 2 61990 64632
0 3084 7 1 2 76928 77023
0 3085 5 3 1 3084
0 3086 7 1 2 77074 81133
0 3087 5 1 1 3086
0 3088 7 1 2 76268 3087
0 3089 5 1 1 3088
0 3090 7 1 2 1399 3089
0 3091 5 1 1 3090
0 3092 7 1 2 71797 3091
0 3093 5 1 1 3092
0 3094 7 1 2 75446 79634
0 3095 5 1 1 3094
0 3096 7 1 2 3093 3095
0 3097 5 1 1 3096
0 3098 7 1 2 81119 3097
0 3099 5 1 1 3098
0 3100 7 1 2 3052 3099
0 3101 5 1 1 3100
0 3102 7 1 2 69690 3101
0 3103 5 1 1 3102
0 3104 7 1 2 68537 1112
0 3105 5 1 1 3104
0 3106 7 1 2 79673 3105
0 3107 5 2 1 3106
0 3108 7 2 2 68538 76410
0 3109 5 2 1 81138
0 3110 7 1 2 63698 77997
0 3111 7 1 2 77978 3110
0 3112 5 1 1 3111
0 3113 7 1 2 81140 3112
0 3114 5 1 1 3113
0 3115 7 1 2 68290 3114
0 3116 5 1 1 3115
0 3117 7 1 2 81136 3116
0 3118 5 1 1 3117
0 3119 7 1 2 66840 3118
0 3120 5 1 1 3119
0 3121 7 3 2 74764 75104
0 3122 5 1 1 81142
0 3123 7 1 2 81143 71516
0 3124 5 1 1 3123
0 3125 7 1 2 3120 3124
0 3126 5 1 1 3125
0 3127 7 1 2 79060 3126
0 3128 5 1 1 3127
0 3129 7 9 2 69691 81120
0 3130 7 2 2 76309 75282
0 3131 5 2 1 81154
0 3132 7 1 2 75275 81156
0 3133 5 1 1 3132
0 3134 7 1 2 63455 3133
0 3135 5 1 1 3134
0 3136 7 6 2 68539 70840
0 3137 5 2 1 81158
0 3138 7 2 2 73765 81159
0 3139 5 2 1 81166
0 3140 7 1 2 76310 75178
0 3141 5 4 1 3140
0 3142 7 1 2 81168 81170
0 3143 5 2 1 3142
0 3144 7 1 2 62314 81174
0 3145 5 1 1 3144
0 3146 7 1 2 76311 74598
0 3147 5 3 1 3146
0 3148 7 1 2 75339 73894
0 3149 5 1 1 3148
0 3150 7 1 2 81176 3149
0 3151 7 1 2 3145 3150
0 3152 5 1 1 3151
0 3153 7 1 2 62741 3152
0 3154 5 1 1 3153
0 3155 7 1 2 3135 3154
0 3156 5 1 1 3155
0 3157 7 1 2 62499 3156
0 3158 5 1 1 3157
0 3159 7 5 2 63456 65917
0 3160 7 1 2 81179 75283
0 3161 5 3 1 3160
0 3162 7 1 2 71798 74510
0 3163 5 1 1 3162
0 3164 7 1 2 81184 3163
0 3165 5 1 1 3164
0 3166 7 1 2 72342 3165
0 3167 5 1 1 3166
0 3168 7 1 2 3158 3167
0 3169 5 1 1 3168
0 3170 7 1 2 81145 3169
0 3171 5 1 1 3170
0 3172 7 1 2 3128 3171
0 3173 5 1 1 3172
0 3174 7 1 2 65309 3173
0 3175 5 1 1 3174
0 3176 7 4 2 74765 78646
0 3177 7 1 2 80040 79804
0 3178 7 1 2 81187 3177
0 3179 5 1 1 3178
0 3180 7 3 2 70841 72970
0 3181 7 2 2 69692 75233
0 3182 7 1 2 80146 81194
0 3183 7 1 2 81191 3182
0 3184 5 1 1 3183
0 3185 7 1 2 3179 3184
0 3186 5 1 1 3185
0 3187 7 1 2 73114 3186
0 3188 5 1 1 3187
0 3189 7 5 2 66841 68761
0 3190 7 5 2 77466 81196
0 3191 7 11 2 64856 65918
0 3192 7 3 2 69476 81206
0 3193 7 2 2 71646 81217
0 3194 7 1 2 81201 81220
0 3195 5 1 1 3194
0 3196 7 1 2 62500 81175
0 3197 5 1 1 3196
0 3198 7 1 2 73678 75640
0 3199 5 1 1 3198
0 3200 7 1 2 3197 3199
0 3201 5 1 1 3200
0 3202 7 1 2 67134 3201
0 3203 5 1 1 3202
0 3204 7 2 2 76312 79489
0 3205 5 2 1 81222
0 3206 7 1 2 71487 81223
0 3207 5 2 1 3206
0 3208 7 1 2 3203 81226
0 3209 5 1 1 3208
0 3210 7 1 2 81121 74233
0 3211 7 1 2 3209 3210
0 3212 5 1 1 3211
0 3213 7 1 2 3195 3212
0 3214 5 1 1 3213
0 3215 7 1 2 70217 3214
0 3216 5 1 1 3215
0 3217 7 1 2 3188 3216
0 3218 7 1 2 3175 3217
0 3219 5 1 1 3218
0 3220 7 1 2 69908 3219
0 3221 5 1 1 3220
0 3222 7 1 2 3103 3221
0 3223 5 1 1 3222
0 3224 7 1 2 61725 3223
0 3225 5 1 1 3224
0 3226 7 1 2 79009 73710
0 3227 5 1 1 3226
0 3228 7 1 2 63457 76929
0 3229 5 3 1 3228
0 3230 7 1 2 76983 81228
0 3231 5 2 1 3230
0 3232 7 1 2 72012 76269
0 3233 7 1 2 81231 3232
0 3234 5 1 1 3233
0 3235 7 1 2 3227 3234
0 3236 5 1 1 3235
0 3237 7 5 2 64857 75464
0 3238 7 16 2 69477 70600
0 3239 7 1 2 81233 81238
0 3240 7 1 2 3236 3239
0 3241 5 1 1 3240
0 3242 7 1 2 3225 3241
0 3243 5 1 1 3242
0 3244 7 1 2 81077 3243
0 3245 5 1 1 3244
0 3246 7 1 2 68054 3245
0 3247 7 1 2 3080 3246
0 3248 7 1 2 2549 3247
0 3249 5 1 1 3248
0 3250 7 1 2 66069 3249
0 3251 7 1 2 2167 3250
0 3252 5 1 1 3251
0 3253 7 16 2 64633 76106
0 3254 7 1 2 78088 668
0 3255 7 18 2 68055 64858
0 3256 5 2 1 81270
0 3257 7 20 2 63218 65044
0 3258 5 3 1 81290
0 3259 7 1 2 81288 81310
0 3260 7 6 2 3254 3259
0 3261 7 1 2 81254 81313
0 3262 5 1 1 3261
0 3263 7 12 2 67588 68056
0 3264 7 4 2 80958 81319
0 3265 7 14 2 69478 69909
0 3266 7 2 2 75046 81335
0 3267 7 1 2 81331 81349
0 3268 5 1 1 3267
0 3269 7 1 2 3262 3268
0 3270 5 1 1 3269
0 3271 7 1 2 67349 3270
0 3272 5 1 1 3271
0 3273 7 10 2 69693 69910
0 3274 7 3 2 68291 81351
0 3275 7 1 2 80454 81332
0 3276 7 1 2 81361 3275
0 3277 5 1 1 3276
0 3278 7 1 2 3272 3277
0 3279 5 1 1 3278
0 3280 7 1 2 66610 3279
0 3281 5 1 1 3280
0 3282 7 11 2 68057 69479
0 3283 7 3 2 81364 78098
0 3284 7 1 2 71034 73371
0 3285 7 2 2 81375 3284
0 3286 5 1 1 81378
0 3287 7 1 2 80959 81379
0 3288 5 1 1 3287
0 3289 7 1 2 3281 3288
0 3290 5 1 1 3289
0 3291 7 1 2 69281 3290
0 3292 5 1 1 3291
0 3293 7 1 2 68058 79061
0 3294 5 1 1 3293
0 3295 7 4 2 63219 79114
0 3296 5 1 1 81380
0 3297 7 1 2 3294 3296
0 3298 5 13 1 3297
0 3299 7 1 2 81384 80124
0 3300 5 1 1 3299
0 3301 7 7 2 69480 73372
0 3302 7 19 2 63220 69694
0 3303 7 5 2 67935 81404
0 3304 5 2 1 81423
0 3305 7 1 2 81397 81424
0 3306 5 1 1 3305
0 3307 7 1 2 3300 3306
0 3308 5 1 1 3307
0 3309 7 1 2 61726 3308
0 3310 5 1 1 3309
0 3311 7 34 2 66611 63221
0 3312 5 1 1 81430
0 3313 7 2 2 81431 79062
0 3314 5 1 1 81464
0 3315 7 1 2 81465 80125
0 3316 5 1 1 3315
0 3317 7 1 2 3310 3316
0 3318 5 1 1 3317
0 3319 7 1 2 79526 80621
0 3320 7 1 2 3318 3319
0 3321 5 1 1 3320
0 3322 7 1 2 3292 3321
0 3323 5 1 1 3322
0 3324 7 1 2 70218 3323
0 3325 5 1 1 3324
0 3326 7 14 2 63069 69481
0 3327 5 2 1 81466
0 3328 7 12 2 64431 81467
0 3329 5 2 1 81482
0 3330 7 1 2 71189 80622
0 3331 7 1 2 81483 3330
0 3332 7 4 2 61727 81320
0 3333 7 4 2 65310 78582
0 3334 7 1 2 81496 81500
0 3335 7 1 2 3331 3334
0 3336 5 1 1 3335
0 3337 7 1 2 3325 3336
0 3338 5 1 1 3337
0 3339 7 1 2 66070 3338
0 3340 5 1 1 3339
0 3341 7 3 2 26 76544
0 3342 7 2 2 79742 79932
0 3343 7 2 2 81504 81507
0 3344 7 12 2 67350 67936
0 3345 7 3 2 81321 81511
0 3346 7 13 2 68762 64432
0 3347 7 1 2 68292 81526
0 3348 7 1 2 81523 3347
0 3349 7 1 2 81509 3348
0 3350 5 1 1 3349
0 3351 7 1 2 3340 3350
0 3352 5 1 1 3351
0 3353 7 1 2 66842 3352
0 3354 5 1 1 3353
0 3355 7 22 2 68059 68293
0 3356 7 3 2 67351 81539
0 3357 7 1 2 79760 81561
0 3358 5 1 1 3357
0 3359 7 6 2 64433 81336
0 3360 7 3 2 63222 76360
0 3361 7 1 2 81564 81570
0 3362 5 1 1 3361
0 3363 7 1 2 3358 3362
0 3364 5 1 1 3363
0 3365 7 1 2 66612 3364
0 3366 5 1 1 3365
0 3367 7 2 2 79332 80688
0 3368 7 25 2 68060 63458
0 3369 7 3 2 61728 81575
0 3370 7 1 2 81573 81600
0 3371 5 1 1 3370
0 3372 7 1 2 3366 3371
0 3373 5 1 1 3372
0 3374 7 1 2 76107 3373
0 3375 5 1 1 3374
0 3376 7 2 2 69911 79411
0 3377 7 40 2 63223 63459
0 3378 7 16 2 66613 67937
0 3379 7 14 2 66357 67352
0 3380 7 2 2 81645 81661
0 3381 7 1 2 81605 81675
0 3382 7 1 2 81603 3381
0 3383 5 1 1 3382
0 3384 7 1 2 3375 3383
0 3385 5 1 1 3384
0 3386 7 1 2 69695 3385
0 3387 5 1 1 3386
0 3388 7 6 2 61729 63460
0 3389 7 2 2 61434 81677
0 3390 7 3 2 64634 78529
0 3391 7 17 2 63224 64434
0 3392 7 1 2 81688 80126
0 3393 7 1 2 81685 3392
0 3394 7 1 2 81683 3393
0 3395 5 1 1 3394
0 3396 7 1 2 3387 3395
0 3397 5 1 1 3396
0 3398 7 11 2 66071 61991
0 3399 7 1 2 70219 81705
0 3400 7 1 2 3397 3399
0 3401 5 1 1 3400
0 3402 7 1 2 3354 3401
0 3403 5 1 1 3402
0 3404 7 1 2 65655 3403
0 3405 5 1 1 3404
0 3406 7 2 2 66843 80217
0 3407 7 1 2 81716 81376
0 3408 5 1 1 3407
0 3409 7 28 2 67938 63225
0 3410 7 1 2 78053 81718
0 3411 5 2 1 3410
0 3412 7 36 2 63070 68061
0 3413 7 2 2 81038 81748
0 3414 5 2 1 81784
0 3415 7 1 2 81746 81786
0 3416 5 6 1 3415
0 3417 7 1 2 81788 81122
0 3418 5 1 1 3417
0 3419 7 1 2 3408 3418
0 3420 5 1 1 3419
0 3421 7 1 2 71413 3420
0 3422 5 1 1 3421
0 3423 7 5 2 66844 69482
0 3424 7 2 2 81794 79764
0 3425 7 33 2 67939 68062
0 3426 7 1 2 81801 78530
0 3427 7 1 2 81799 3426
0 3428 5 1 1 3427
0 3429 7 1 2 3422 3428
0 3430 5 1 1 3429
0 3431 7 1 2 66358 3430
0 3432 5 1 1 3431
0 3433 7 18 2 61435 68063
0 3434 7 3 2 79731 81834
0 3435 7 7 2 65045 79115
0 3436 7 1 2 74212 81855
0 3437 7 1 2 81852 3436
0 3438 5 1 1 3437
0 3439 7 1 2 3432 3438
0 3440 5 1 1 3439
0 3441 7 4 2 68763 69282
0 3442 7 2 2 70220 81862
0 3443 7 7 2 66072 67353
0 3444 7 1 2 81866 81868
0 3445 7 1 2 3440 3444
0 3446 5 1 1 3445
0 3447 7 1 2 3405 3446
0 3448 5 1 1 3447
0 3449 7 1 2 71890 3448
0 3450 5 1 1 3449
0 3451 7 7 2 67354 69283
0 3452 7 2 2 74766 79063
0 3453 7 1 2 66845 81882
0 3454 5 2 1 3453
0 3455 7 11 2 63699 64635
0 3456 7 5 2 61992 69696
0 3457 7 1 2 81886 81897
0 3458 5 1 1 3457
0 3459 7 1 2 81884 3458
0 3460 5 2 1 3459
0 3461 7 1 2 66614 81902
0 3462 5 1 1 3461
0 3463 7 1 2 79147 80613
0 3464 5 1 1 3463
0 3465 7 1 2 3462 3464
0 3466 5 1 1 3465
0 3467 7 1 2 76108 3466
0 3468 5 1 1 3467
0 3469 7 69 2 66359 69483
0 3470 5 2 1 81904
0 3471 7 39 2 61730 69697
0 3472 5 1 1 81975
0 3473 7 2 2 81905 81976
0 3474 7 1 2 67940 82014
0 3475 5 1 1 3474
0 3476 7 9 2 66615 78461
0 3477 7 1 2 77218 82016
0 3478 5 1 1 3477
0 3479 7 1 2 3475 3478
0 3480 5 4 1 3479
0 3481 7 1 2 80614 82025
0 3482 5 1 1 3481
0 3483 7 1 2 3468 3482
0 3484 5 1 1 3483
0 3485 7 1 2 81039 3484
0 3486 5 1 1 3485
0 3487 7 4 2 66616 75570
0 3488 7 1 2 67135 82029
0 3489 7 9 2 64636 81352
0 3490 7 2 2 66360 74878
0 3491 7 1 2 82033 82042
0 3492 7 1 2 3488 3491
0 3493 5 1 1 3492
0 3494 7 1 2 3486 3493
0 3495 5 1 1 3494
0 3496 7 1 2 81875 3495
0 3497 5 1 1 3496
0 3498 7 16 2 61731 67136
0 3499 7 2 2 82044 79816
0 3500 7 1 2 61436 82060
0 3501 7 5 2 65046 75047
0 3502 7 2 2 79333 80127
0 3503 5 1 1 82067
0 3504 7 1 2 82062 82068
0 3505 7 1 2 3500 3504
0 3506 5 1 1 3505
0 3507 7 1 2 3497 3506
0 3508 5 1 1 3507
0 3509 7 1 2 66073 3508
0 3510 5 1 1 3509
0 3511 7 4 2 66846 74949
0 3512 7 1 2 68540 80024
0 3513 7 1 2 82069 3512
0 3514 7 10 2 64435 64859
0 3515 7 4 2 79743 82073
0 3516 7 1 2 81505 82083
0 3517 7 1 2 3513 3516
0 3518 5 1 1 3517
0 3519 7 1 2 3510 3518
0 3520 5 1 1 3519
0 3521 7 1 2 68064 3520
0 3522 5 1 1 3521
0 3523 7 2 2 69912 81719
0 3524 7 9 2 66074 66361
0 3525 7 1 2 79792 74395
0 3526 7 1 2 82089 3525
0 3527 7 1 2 82087 3526
0 3528 7 1 2 81903 3527
0 3529 5 1 1 3528
0 3530 7 1 2 3522 3529
0 3531 5 1 1 3530
0 3532 7 1 2 73235 3531
0 3533 5 1 1 3532
0 3534 7 28 2 66362 69284
0 3535 7 19 2 63226 68541
0 3536 7 2 2 82126 76361
0 3537 7 15 2 66617 67137
0 3538 7 16 2 64860 65656
0 3539 7 1 2 82147 82162
0 3540 7 1 2 82145 3539
0 3541 5 1 1 3540
0 3542 7 3 2 63700 79884
0 3543 5 7 1 82178
0 3544 7 1 2 68294 77881
0 3545 7 1 2 82181 3544
0 3546 5 1 1 3545
0 3547 7 15 2 67138 63461
0 3548 5 1 1 82188
0 3549 7 11 2 68542 82189
0 3550 5 2 1 82203
0 3551 7 1 2 71190 82204
0 3552 5 1 1 3551
0 3553 7 1 2 3546 3552
0 3554 5 1 1 3553
0 3555 7 1 2 68065 71474
0 3556 7 1 2 3554 3555
0 3557 5 1 1 3556
0 3558 7 1 2 3541 3557
0 3559 5 1 1 3558
0 3560 7 1 2 82098 3559
0 3561 5 1 1 3560
0 3562 7 5 2 63701 73373
0 3563 7 2 2 65657 82216
0 3564 5 1 1 82221
0 3565 7 1 2 71502 3564
0 3566 5 1 1 3565
0 3567 7 1 2 68295 3566
0 3568 5 1 1 3567
0 3569 7 1 2 81137 3568
0 3570 5 2 1 3569
0 3571 7 21 2 64436 69698
0 3572 7 6 2 61437 63227
0 3573 7 2 2 82225 82246
0 3574 7 1 2 61732 82252
0 3575 7 1 2 82223 3574
0 3576 5 1 1 3575
0 3577 7 1 2 3561 3576
0 3578 5 1 1 3577
0 3579 7 1 2 67941 3578
0 3580 5 1 1 3579
0 3581 7 3 2 71191 72971
0 3582 5 3 1 82254
0 3583 7 1 2 74045 82257
0 3584 5 3 1 3583
0 3585 7 1 2 81432 82260
0 3586 5 1 1 3585
0 3587 7 7 2 68066 63702
0 3588 7 1 2 79765 82263
0 3589 5 1 1 3588
0 3590 7 1 2 3586 3589
0 3591 5 1 1 3590
0 3592 7 23 2 67589 64437
0 3593 7 6 2 77219 82270
0 3594 5 1 1 82293
0 3595 7 1 2 82163 82294
0 3596 7 1 2 3591 3595
0 3597 5 1 1 3596
0 3598 7 1 2 3580 3597
0 3599 5 1 1 3598
0 3600 7 1 2 69484 3599
0 3601 5 1 1 3600
0 3602 7 3 2 64438 72972
0 3603 7 10 2 61438 67355
0 3604 7 5 2 82302 80128
0 3605 7 1 2 82299 82312
0 3606 5 1 1 3605
0 3607 7 32 2 69285 80960
0 3608 5 1 1 82317
0 3609 7 1 2 82318 82205
0 3610 5 1 1 3609
0 3611 7 1 2 3606 3610
0 3612 5 1 1 3611
0 3613 7 1 2 68764 3612
0 3614 5 1 1 3613
0 3615 7 5 2 63703 64439
0 3616 7 2 2 68296 82349
0 3617 7 5 2 61439 80129
0 3618 7 1 2 82354 82356
0 3619 5 1 1 3618
0 3620 7 1 2 3614 3619
0 3621 5 1 1 3620
0 3622 7 25 2 61733 63228
0 3623 5 3 1 82361
0 3624 7 10 2 69699 65658
0 3625 7 5 2 64637 82389
0 3626 7 1 2 82362 82399
0 3627 7 1 2 3621 3626
0 3628 5 1 1 3627
0 3629 7 1 2 3601 3628
0 3630 5 1 1 3629
0 3631 7 1 2 69913 3630
0 3632 5 1 1 3631
0 3633 7 12 2 67139 68297
0 3634 5 1 1 82404
0 3635 7 9 2 68067 68543
0 3636 7 7 2 82405 82416
0 3637 7 16 2 69286 65659
0 3638 7 1 2 80767 82432
0 3639 7 1 2 82425 3638
0 3640 7 1 2 82026 3639
0 3641 5 1 1 3640
0 3642 7 1 2 3632 3641
0 3643 5 1 1 3642
0 3644 7 1 2 66847 3643
0 3645 5 1 1 3644
0 3646 7 4 2 81689 80481
0 3647 7 3 2 61734 72690
0 3648 7 6 2 68765 79294
0 3649 7 1 2 82452 82455
0 3650 5 2 1 3649
0 3651 7 10 2 66618 69914
0 3652 5 1 1 82463
0 3653 7 2 2 61993 82464
0 3654 5 1 1 82473
0 3655 7 1 2 82461 3654
0 3656 5 1 1 3655
0 3657 7 1 2 72973 3656
0 3658 5 1 1 3657
0 3659 7 3 2 65660 80689
0 3660 7 2 2 66619 74449
0 3661 7 1 2 82475 82478
0 3662 5 1 1 3661
0 3663 7 1 2 3658 3662
0 3664 5 1 1 3663
0 3665 7 1 2 82448 3664
0 3666 5 1 1 3665
0 3667 7 6 2 68544 75844
0 3668 5 1 1 82480
0 3669 7 6 2 68298 71562
0 3670 5 3 1 82486
0 3671 7 1 2 82481 82487
0 3672 5 1 1 3671
0 3673 7 7 2 63462 65661
0 3674 5 3 1 82495
0 3675 7 2 2 63704 78647
0 3676 7 1 2 82496 82505
0 3677 5 1 1 3676
0 3678 7 1 2 3672 3677
0 3679 5 1 1 3678
0 3680 7 1 2 66620 3679
0 3681 5 1 1 3680
0 3682 7 8 2 68299 74767
0 3683 7 1 2 75394 71517
0 3684 7 1 2 82507 3683
0 3685 5 1 1 3684
0 3686 7 1 2 3681 3685
0 3687 5 1 1 3686
0 3688 7 1 2 79463 3687
0 3689 5 1 1 3688
0 3690 7 3 2 63463 74147
0 3691 7 1 2 81565 82515
0 3692 7 1 2 101 3691
0 3693 5 1 1 3692
0 3694 7 1 2 3689 3693
0 3695 5 1 1 3694
0 3696 7 1 2 68068 3695
0 3697 5 1 1 3696
0 3698 7 1 2 3666 3697
0 3699 5 1 1 3698
0 3700 7 1 2 69700 3699
0 3701 5 1 1 3700
0 3702 7 13 2 68545 68766
0 3703 5 3 1 82518
0 3704 7 4 2 67140 82519
0 3705 7 15 2 63229 64638
0 3706 7 5 2 78054 82538
0 3707 5 2 1 82553
0 3708 7 6 2 65047 81540
0 3709 7 1 2 69485 82560
0 3710 5 1 1 3709
0 3711 7 1 2 82558 3710
0 3712 5 4 1 3711
0 3713 7 1 2 82534 82566
0 3714 5 1 1 3713
0 3715 7 16 2 67356 63230
0 3716 7 2 2 69915 82570
0 3717 7 4 2 68300 81887
0 3718 7 1 2 82586 82588
0 3719 5 1 1 3718
0 3720 7 1 2 3714 3719
0 3721 5 1 1 3720
0 3722 7 18 2 69287 64861
0 3723 7 29 2 66621 66848
0 3724 7 3 2 82592 82610
0 3725 7 1 2 65662 82639
0 3726 7 1 2 3721 3725
0 3727 5 1 1 3726
0 3728 7 1 2 3701 3727
0 3729 5 1 1 3728
0 3730 7 1 2 76109 3729
0 3731 5 1 1 3730
0 3732 7 9 2 64639 80779
0 3733 5 1 1 82642
0 3734 7 26 2 63071 63231
0 3735 7 9 2 61994 64440
0 3736 7 2 2 82651 82677
0 3737 7 2 2 82643 82686
0 3738 7 5 2 65663 76452
0 3739 7 1 2 82688 82690
0 3740 5 1 1 3739
0 3741 7 14 2 66363 66849
0 3742 7 2 2 67942 82695
0 3743 7 9 2 68069 73904
0 3744 7 4 2 69288 81239
0 3745 7 1 2 82711 82720
0 3746 7 1 2 82709 3745
0 3747 5 1 1 3746
0 3748 7 1 2 3740 3747
0 3749 5 1 1 3748
0 3750 7 1 2 71035 3749
0 3751 5 1 1 3750
0 3752 7 28 2 66622 68070
0 3753 5 3 1 82724
0 3754 7 8 2 67943 80918
0 3755 7 4 2 82725 82755
0 3756 7 3 2 66850 73905
0 3757 7 21 2 69486 69701
0 3758 7 5 2 69289 82770
0 3759 7 1 2 70601 82791
0 3760 7 1 2 82767 3759
0 3761 7 1 2 82763 3760
0 3762 5 1 1 3761
0 3763 7 1 2 3751 3762
0 3764 5 1 1 3763
0 3765 7 1 2 71291 3764
0 3766 5 1 1 3765
0 3767 7 4 2 67357 81802
0 3768 7 2 2 82796 80881
0 3769 7 15 2 69290 69487
0 3770 7 3 2 64862 82802
0 3771 7 6 2 68301 82520
0 3772 7 1 2 82817 82820
0 3773 7 1 2 82800 3772
0 3774 5 1 1 3773
0 3775 7 2 2 76813 77594
0 3776 5 1 1 82826
0 3777 7 2 2 78462 80130
0 3778 7 1 2 82827 82828
0 3779 5 1 1 3778
0 3780 7 2 2 73802 79470
0 3781 7 1 2 80903 75346
0 3782 7 1 2 82830 3781
0 3783 5 1 1 3782
0 3784 7 1 2 3779 3783
0 3785 5 1 1 3784
0 3786 7 27 2 61440 64441
0 3787 7 7 2 63232 65664
0 3788 7 1 2 82832 82859
0 3789 7 1 2 3785 3788
0 3790 5 1 1 3789
0 3791 7 1 2 3774 3790
0 3792 5 1 1 3791
0 3793 7 1 2 61735 3792
0 3794 5 1 1 3793
0 3795 7 8 2 64640 81606
0 3796 7 1 2 73283 82866
0 3797 5 1 1 3796
0 3798 7 11 2 67141 68071
0 3799 7 2 2 82874 80904
0 3800 7 6 2 67358 71010
0 3801 5 7 1 82887
0 3802 7 1 2 82885 82888
0 3803 5 1 1 3802
0 3804 7 1 2 3797 3803
0 3805 5 1 1 3804
0 3806 7 7 2 69291 69702
0 3807 7 2 2 68546 82900
0 3808 7 1 2 76545 74213
0 3809 7 1 2 82907 3808
0 3810 7 1 2 3805 3809
0 3811 5 1 1 3810
0 3812 7 1 2 3794 3811
0 3813 7 1 2 3766 3812
0 3814 5 1 1 3813
0 3815 7 1 2 69916 3814
0 3816 5 1 1 3815
0 3817 7 8 2 61441 74148
0 3818 7 8 2 63233 74256
0 3819 7 2 2 82909 82917
0 3820 7 4 2 62315 80131
0 3821 7 3 2 64442 78463
0 3822 7 1 2 77748 82931
0 3823 7 1 2 82927 3822
0 3824 7 1 2 82925 3823
0 3825 5 1 1 3824
0 3826 7 1 2 3816 3825
0 3827 7 1 2 3731 3826
0 3828 7 1 2 3645 3827
0 3829 5 1 1 3828
0 3830 7 1 2 66075 3829
0 3831 5 1 1 3830
0 3832 7 1 2 3533 3831
0 3833 5 1 1 3832
0 3834 7 1 2 65311 3833
0 3835 5 1 1 3834
0 3836 7 8 2 69292 69917
0 3837 7 1 2 68547 81541
0 3838 7 2 2 82934 3837
0 3839 7 4 2 80919 80083
0 3840 7 1 2 66623 82944
0 3841 7 1 2 82942 3840
0 3842 5 1 1 3841
0 3843 7 5 2 66624 63464
0 3844 7 2 2 69918 82948
0 3845 5 1 1 82953
0 3846 7 1 2 3845 82462
0 3847 5 1 1 3846
0 3848 7 1 2 76064 3847
0 3849 5 1 1 3848
0 3850 7 2 2 75691 82303
0 3851 7 1 2 67944 82456
0 3852 7 1 2 82955 3851
0 3853 5 1 1 3852
0 3854 7 1 2 3849 3853
0 3855 5 1 1 3854
0 3856 7 3 2 64443 71799
0 3857 7 1 2 63234 82957
0 3858 7 1 2 3855 3857
0 3859 5 1 1 3858
0 3860 7 1 2 3842 3859
0 3861 5 1 1 3860
0 3862 7 1 2 69488 3861
0 3863 5 1 1 3862
0 3864 7 12 2 65048 71800
0 3865 5 1 1 82960
0 3866 7 5 2 69919 74768
0 3867 5 1 1 82972
0 3868 7 1 2 3867 78121
0 3869 7 1 2 3865 3868
0 3870 5 2 1 3869
0 3871 7 2 2 82571 71518
0 3872 7 19 2 64444 64641
0 3873 7 3 2 77220 75692
0 3874 7 1 2 82981 83000
0 3875 7 1 2 82979 3874
0 3876 7 1 2 82977 3875
0 3877 5 1 1 3876
0 3878 7 1 2 3863 3877
0 3879 5 1 1 3878
0 3880 7 1 2 70221 3879
0 3881 5 1 1 3880
0 3882 7 2 2 66364 81789
0 3883 5 1 1 83003
0 3884 7 8 2 68072 81040
0 3885 7 2 2 76031 83005
0 3886 5 1 1 83013
0 3887 7 1 2 3883 3886
0 3888 5 3 1 3887
0 3889 7 2 2 71770 77595
0 3890 7 1 2 79412 71563
0 3891 7 1 2 83018 3890
0 3892 7 1 2 83015 3891
0 3893 5 1 1 3892
0 3894 7 1 2 3881 3893
0 3895 5 1 1 3894
0 3896 7 1 2 69703 3895
0 3897 5 1 1 3896
0 3898 7 2 2 69489 80289
0 3899 7 3 2 80961 82045
0 3900 7 1 2 82943 83022
0 3901 5 1 1 3900
0 3902 7 46 2 61736 68073
0 3903 5 1 1 83025
0 3904 7 3 2 3903 3312
0 3905 5 96 1 83071
0 3906 7 8 2 69920 83074
0 3907 7 1 2 74853 83170
0 3908 5 1 1 3907
0 3909 7 1 2 81291 77741
0 3910 5 1 1 3909
0 3911 7 1 2 3908 3910
0 3912 5 1 1 3911
0 3913 7 2 2 65665 81527
0 3914 7 1 2 82313 83178
0 3915 7 1 2 3912 3914
0 3916 5 1 1 3915
0 3917 7 1 2 3901 3916
0 3918 5 1 1 3917
0 3919 7 1 2 83020 3918
0 3920 5 1 1 3919
0 3921 7 1 2 3897 3920
0 3922 5 1 1 3921
0 3923 7 1 2 66851 3922
0 3924 5 1 1 3923
0 3925 7 5 2 68767 64863
0 3926 7 1 2 78142 76642
0 3927 7 1 2 83180 3926
0 3928 7 5 2 67590 72438
0 3929 5 3 1 83185
0 3930 7 4 2 63072 77179
0 3931 7 1 2 83193 82449
0 3932 7 1 2 83186 3931
0 3933 7 1 2 3927 3932
0 3934 5 1 1 3933
0 3935 7 1 2 3924 3934
0 3936 5 1 1 3935
0 3937 7 1 2 66076 3936
0 3938 5 1 1 3937
0 3939 7 1 2 3835 3938
0 3940 7 1 2 3450 3939
0 3941 5 1 1 3940
0 3942 7 1 2 72096 3941
0 3943 5 1 1 3942
0 3944 7 4 2 66077 63465
0 3945 7 16 2 69921 65919
0 3946 5 1 1 83201
0 3947 7 12 2 63235 68924
0 3948 7 2 2 83202 83217
0 3949 7 4 2 67591 78908
0 3950 5 1 1 83231
0 3951 7 1 2 78899 3950
0 3952 5 2 1 3951
0 3953 7 1 2 81977 83235
0 3954 5 1 1 3953
0 3955 7 1 2 79064 76659
0 3956 5 2 1 3955
0 3957 7 1 2 3954 83237
0 3958 5 1 1 3957
0 3959 7 1 2 64445 3958
0 3960 5 1 1 3959
0 3961 7 3 2 69293 80218
0 3962 7 1 2 82017 83239
0 3963 5 2 1 3962
0 3964 7 1 2 3960 83242
0 3965 5 1 1 3964
0 3966 7 1 2 61442 3965
0 3967 5 1 1 3966
0 3968 7 5 2 82099 78464
0 3969 7 3 2 83244 76660
0 3970 5 1 1 83249
0 3971 7 1 2 67592 83250
0 3972 5 1 1 3971
0 3973 7 1 2 3967 3972
0 3974 5 1 1 3973
0 3975 7 1 2 83229 3974
0 3976 5 1 1 3975
0 3977 7 2 2 80219 79413
0 3978 5 1 1 83252
0 3979 7 1 2 81494 3978
0 3980 5 2 1 3979
0 3981 7 1 2 61443 83254
0 3982 5 2 1 3981
0 3983 7 4 2 63073 79414
0 3984 7 1 2 80920 83258
0 3985 5 1 1 3984
0 3986 7 1 2 83256 3985
0 3987 5 3 1 3986
0 3988 7 7 2 69922 72508
0 3989 7 2 2 71036 83265
0 3990 7 1 2 68074 83272
0 3991 7 1 2 83262 3990
0 3992 5 1 1 3991
0 3993 7 1 2 3976 3992
0 3994 5 1 1 3993
0 3995 7 1 2 83197 3994
0 3996 5 1 1 3995
0 3997 7 3 2 67945 78465
0 3998 7 1 2 81506 83274
0 3999 5 1 1 3998
0 4000 7 19 2 61444 61737
0 4001 7 5 2 66078 83277
0 4002 7 1 2 69490 80504
0 4003 7 1 2 83296 4002
0 4004 5 1 1 4003
0 4005 7 1 2 3999 4004
0 4006 5 1 1 4005
0 4007 7 1 2 64446 4006
0 4008 5 1 1 4007
0 4009 7 7 2 66079 67593
0 4010 7 3 2 69294 83301
0 4011 7 2 2 69704 77180
0 4012 5 1 1 83311
0 4013 7 5 2 64864 78490
0 4014 5 2 1 83313
0 4015 7 1 2 4012 83318
0 4016 5 4 1 4015
0 4017 7 1 2 83320 78943
0 4018 5 1 1 4017
0 4019 7 23 2 61738 64642
0 4020 5 1 1 83324
0 4021 7 16 2 69705 83325
0 4022 7 1 2 76032 83347
0 4023 5 1 1 4022
0 4024 7 1 2 76065 78276
0 4025 5 1 1 4024
0 4026 7 1 2 4023 4025
0 4027 7 1 2 4018 4026
0 4028 5 1 1 4027
0 4029 7 1 2 83308 4028
0 4030 5 1 1 4029
0 4031 7 1 2 4008 4030
0 4032 5 1 1 4031
0 4033 7 5 2 62501 72600
0 4034 5 6 1 83363
0 4035 7 1 2 83006 83368
0 4036 7 1 2 4032 4035
0 4037 5 1 1 4036
0 4038 7 1 2 3996 4037
0 4039 5 1 1 4038
0 4040 7 1 2 74769 4039
0 4041 5 1 1 4040
0 4042 7 16 2 68075 64643
0 4043 5 1 1 83374
0 4044 7 9 2 63466 69295
0 4045 7 2 2 78670 83390
0 4046 7 1 2 83375 83399
0 4047 5 1 1 4046
0 4048 7 1 2 81690 81350
0 4049 5 1 1 4048
0 4050 7 1 2 4047 4049
0 4051 5 1 1 4050
0 4052 7 1 2 61445 4051
0 4053 5 1 1 4052
0 4054 7 25 2 63236 68302
0 4055 7 2 2 66365 83401
0 4056 7 2 2 79116 82935
0 4057 7 1 2 83426 83428
0 4058 5 1 1 4057
0 4059 7 1 2 4053 4058
0 4060 5 1 1 4059
0 4061 7 1 2 67946 4060
0 4062 5 1 1 4061
0 4063 7 1 2 76066 81576
0 4064 7 1 2 79785 4063
0 4065 5 1 1 4064
0 4066 7 1 2 4062 4065
0 4067 5 1 1 4066
0 4068 7 1 2 67594 4067
0 4069 5 1 1 4068
0 4070 7 4 2 63237 80700
0 4071 7 1 2 83430 75347
0 4072 5 1 1 4071
0 4073 7 7 2 63074 81542
0 4074 7 1 2 78531 83434
0 4075 5 1 1 4074
0 4076 7 1 2 4072 4075
0 4077 5 2 1 4076
0 4078 7 1 2 61446 83441
0 4079 5 1 1 4078
0 4080 7 2 2 76067 81607
0 4081 7 1 2 78583 83443
0 4082 5 1 1 4081
0 4083 7 1 2 4079 4082
0 4084 5 1 1 4083
0 4085 7 1 2 79334 4084
0 4086 5 1 1 4085
0 4087 7 1 2 4069 4086
0 4088 5 1 1 4087
0 4089 7 1 2 61739 4088
0 4090 5 1 1 4089
0 4091 7 2 2 67595 81720
0 4092 7 3 2 69491 78532
0 4093 7 10 2 66366 68303
0 4094 7 1 2 79793 83450
0 4095 7 1 2 83447 4094
0 4096 7 1 2 83445 4095
0 4097 5 1 1 4096
0 4098 7 1 2 4090 4097
0 4099 5 1 1 4098
0 4100 7 2 2 66080 63705
0 4101 7 1 2 72509 83460
0 4102 7 1 2 4099 4101
0 4103 5 1 1 4102
0 4104 7 1 2 4041 4103
0 4105 5 1 1 4104
0 4106 7 1 2 66852 4105
0 4107 5 1 1 4106
0 4108 7 7 2 65920 73736
0 4109 7 6 2 68548 69706
0 4110 7 2 2 67142 83469
0 4111 5 2 1 83475
0 4112 7 1 2 1927 83477
0 4113 5 1 1 4112
0 4114 7 2 2 1818 4113
0 4115 7 1 2 63467 83479
0 4116 5 1 1 4115
0 4117 7 2 2 78584 74022
0 4118 5 1 1 83481
0 4119 7 1 2 4116 4118
0 4120 5 1 1 4119
0 4121 7 1 2 61740 4120
0 4122 5 1 1 4121
0 4123 7 4 2 69923 75680
0 4124 7 2 2 79849 83483
0 4125 5 1 1 83487
0 4126 7 1 2 63468 83488
0 4127 5 1 1 4126
0 4128 7 1 2 4122 4127
0 4129 5 1 1 4128
0 4130 7 1 2 76110 4129
0 4131 5 1 1 4130
0 4132 7 3 2 67596 82046
0 4133 7 1 2 69924 83470
0 4134 7 1 2 80636 4133
0 4135 7 1 2 83489 4134
0 4136 5 1 1 4135
0 4137 7 1 2 4131 4136
0 4138 5 1 1 4137
0 4139 7 1 2 69492 4138
0 4140 5 1 1 4139
0 4141 7 9 2 63469 64644
0 4142 7 3 2 83492 80819
0 4143 7 3 2 78491 81353
0 4144 7 1 2 83501 83504
0 4145 5 1 1 4144
0 4146 7 1 2 4140 4145
0 4147 5 1 1 4146
0 4148 7 1 2 63238 4147
0 4149 5 1 1 4148
0 4150 7 5 2 66367 80132
0 4151 5 1 1 83507
0 4152 7 3 2 63470 79850
0 4153 7 1 2 83508 83512
0 4154 5 1 1 4153
0 4155 7 11 2 63471 69707
0 4156 7 2 2 79278 83515
0 4157 7 1 2 67597 83526
0 4158 5 1 1 4157
0 4159 7 1 2 75992 82508
0 4160 5 1 1 4159
0 4161 7 1 2 4158 4160
0 4162 5 1 1 4161
0 4163 7 1 2 61447 4162
0 4164 5 1 1 4163
0 4165 7 1 2 4154 4164
0 4166 5 1 1 4165
0 4167 7 7 2 61741 69493
0 4168 7 18 2 68076 69925
0 4169 5 1 1 83535
0 4170 7 1 2 83528 83536
0 4171 7 1 2 4166 4170
0 4172 5 1 1 4171
0 4173 7 1 2 4149 4172
0 4174 5 1 1 4173
0 4175 7 1 2 64447 4174
0 4176 5 1 1 4175
0 4177 7 8 2 63706 69296
0 4178 7 2 2 78466 83553
0 4179 7 1 2 75693 83561
0 4180 7 1 2 83016 4179
0 4181 5 1 1 4180
0 4182 7 1 2 4176 4181
0 4183 5 1 1 4182
0 4184 7 1 2 83462 4183
0 4185 5 1 1 4184
0 4186 7 7 2 63472 82652
0 4187 7 3 2 83563 82958
0 4188 5 2 1 83570
0 4189 7 27 2 64645 69926
0 4190 7 2 2 76841 83575
0 4191 7 1 2 83278 79235
0 4192 7 1 2 83602 4191
0 4193 7 1 2 83571 4192
0 4194 5 1 1 4193
0 4195 7 1 2 4185 4194
0 4196 5 1 1 4195
0 4197 7 1 2 66081 4196
0 4198 5 1 1 4197
0 4199 7 1 2 4107 4198
0 4200 5 1 1 4199
0 4201 7 1 2 65312 4200
0 4202 5 1 1 4201
0 4203 7 4 2 66853 74564
0 4204 5 4 1 83604
0 4205 7 9 2 61995 74770
0 4206 5 3 1 83612
0 4207 7 1 2 83608 83621
0 4208 5 1 1 4207
0 4209 7 12 2 69297 78467
0 4210 7 2 2 81041 83624
0 4211 5 2 1 83636
0 4212 7 3 2 69494 81354
0 4213 7 11 2 63473 64448
0 4214 7 1 2 83640 83643
0 4215 5 1 1 4214
0 4216 7 1 2 83638 4215
0 4217 5 4 1 4216
0 4218 7 1 2 83026 83654
0 4219 5 1 1 4218
0 4220 7 5 2 81337 82226
0 4221 7 5 2 66625 81608
0 4222 7 1 2 83658 83663
0 4223 5 1 1 4222
0 4224 7 1 2 4219 4223
0 4225 5 1 1 4224
0 4226 7 1 2 76111 4225
0 4227 5 1 1 4226
0 4228 7 2 2 64646 83391
0 4229 7 13 2 63239 69927
0 4230 7 2 2 83670 78708
0 4231 7 1 2 77181 83683
0 4232 7 1 2 83668 4231
0 4233 5 1 1 4232
0 4234 7 1 2 4227 4233
0 4235 5 1 1 4234
0 4236 7 1 2 4208 4235
0 4237 5 1 1 4236
0 4238 7 10 2 76112 83075
0 4239 7 2 2 70222 83685
0 4240 7 1 2 74450 83695
0 4241 5 1 1 4240
0 4242 7 3 2 66854 83279
0 4243 7 3 2 82127 80084
0 4244 7 1 2 83697 83700
0 4245 5 1 1 4244
0 4246 7 1 2 4241 4245
0 4247 5 1 1 4246
0 4248 7 1 2 75048 81566
0 4249 7 1 2 4247 4248
0 4250 5 1 1 4249
0 4251 7 1 2 4237 4250
0 4252 5 1 1 4251
0 4253 7 7 2 66082 62742
0 4254 7 1 2 72013 83703
0 4255 7 1 2 4252 4254
0 4256 5 1 1 4255
0 4257 7 1 2 4202 4256
0 4258 5 1 1 4257
0 4259 7 1 2 73236 4258
0 4260 5 1 1 4259
0 4261 7 2 2 82100 71414
0 4262 7 8 2 73237 77979
0 4263 5 4 1 83712
0 4264 7 2 2 65921 83713
0 4265 7 1 2 80337 83724
0 4266 5 1 1 4265
0 4267 7 6 2 70223 71292
0 4268 5 14 1 83726
0 4269 7 2 2 70842 83732
0 4270 7 1 2 80335 83746
0 4271 5 1 1 4270
0 4272 7 1 2 4266 4271
0 4273 5 1 1 4272
0 4274 7 1 2 83710 4273
0 4275 5 1 1 4274
0 4276 7 3 2 62743 80603
0 4277 7 1 2 80319 83748
0 4278 5 1 1 4277
0 4279 7 1 2 72407 80105
0 4280 5 1 1 4279
0 4281 7 1 2 4278 4280
0 4282 5 1 1 4281
0 4283 7 1 2 66368 4282
0 4284 5 1 1 4283
0 4285 7 12 2 68768 70602
0 4286 5 2 1 83751
0 4287 7 6 2 62744 64647
0 4288 5 2 1 83765
0 4289 7 2 2 76033 83766
0 4290 5 1 1 83773
0 4291 7 1 2 83752 83774
0 4292 5 1 1 4291
0 4293 7 1 2 4284 4292
0 4294 5 1 1 4293
0 4295 7 1 2 67359 4294
0 4296 5 1 1 4295
0 4297 7 2 2 65922 73238
0 4298 7 2 2 67598 83775
0 4299 5 1 1 83777
0 4300 7 7 2 67947 70224
0 4301 7 2 2 81906 83779
0 4302 7 1 2 83778 83786
0 4303 5 1 1 4302
0 4304 7 1 2 4296 4303
0 4305 5 1 1 4304
0 4306 7 1 2 69298 4305
0 4307 5 1 1 4306
0 4308 7 2 2 79335 73641
0 4309 7 1 2 77221 75658
0 4310 7 1 2 83788 4309
0 4311 5 1 1 4310
0 4312 7 1 2 4307 4311
0 4313 5 1 1 4312
0 4314 7 1 2 68925 4313
0 4315 5 1 1 4314
0 4316 7 36 2 63075 64449
0 4317 7 13 2 61448 83790
0 4318 5 3 1 83826
0 4319 7 5 2 82101 80220
0 4320 5 1 1 83842
0 4321 7 1 2 83839 4320
0 4322 5 5 1 4321
0 4323 7 1 2 81398 72439
0 4324 7 1 2 83847 4323
0 4325 5 1 1 4324
0 4326 7 2 2 81662 72313
0 4327 7 1 2 78373 83259
0 4328 7 1 2 83852 4327
0 4329 5 1 1 4328
0 4330 7 1 2 4325 4329
0 4331 7 1 2 4315 4330
0 4332 5 1 1 4331
0 4333 7 1 2 71037 4332
0 4334 5 1 1 4333
0 4335 7 1 2 4275 4334
0 4336 5 1 1 4335
0 4337 7 1 2 74301 4336
0 4338 5 1 1 4337
0 4339 7 1 2 73239 74745
0 4340 5 1 1 4339
0 4341 7 3 2 72440 71011
0 4342 5 1 1 83854
0 4343 7 1 2 4340 4342
0 4344 5 2 1 4343
0 4345 7 9 2 61742 76113
0 4346 7 4 2 69708 75757
0 4347 7 2 2 79336 83868
0 4348 5 1 1 83872
0 4349 7 1 2 83859 83873
0 4350 7 1 2 83857 4349
0 4351 5 1 1 4350
0 4352 7 1 2 68077 4351
0 4353 7 1 2 4338 4352
0 4354 5 1 1 4353
0 4355 7 6 2 70225 77998
0 4356 5 2 1 83874
0 4357 7 1 2 79162 82833
0 4358 5 1 1 4357
0 4359 7 3 2 66626 83245
0 4360 5 1 1 83882
0 4361 7 1 2 67599 83883
0 4362 5 1 1 4361
0 4363 7 1 2 4358 4362
0 4364 5 1 1 4363
0 4365 7 1 2 83875 4364
0 4366 5 1 1 4365
0 4367 7 9 2 68769 64648
0 4368 7 3 2 82593 83885
0 4369 7 1 2 76546 83894
0 4370 7 1 2 74017 4369
0 4371 5 1 1 4370
0 4372 7 1 2 4366 4371
0 4373 5 1 1 4372
0 4374 7 1 2 80642 4373
0 4375 5 1 1 4374
0 4376 7 12 2 78979 82594
0 4377 5 1 1 83897
0 4378 7 6 2 82227 83529
0 4379 5 6 1 83909
0 4380 7 1 2 4377 83915
0 4381 5 9 1 4380
0 4382 7 2 2 70226 78013
0 4383 5 1 1 83930
0 4384 7 2 2 70603 72745
0 4385 5 1 1 83932
0 4386 7 1 2 62745 83933
0 4387 5 1 1 4386
0 4388 7 1 2 4383 4387
0 4389 5 1 1 4388
0 4390 7 1 2 83921 4389
0 4391 5 1 1 4390
0 4392 7 2 2 82228 81240
0 4393 7 1 2 75694 72314
0 4394 7 1 2 83934 4393
0 4395 5 1 1 4394
0 4396 7 1 2 4391 4395
0 4397 5 1 1 4396
0 4398 7 1 2 61449 4397
0 4399 5 1 1 4398
0 4400 7 5 2 69299 80921
0 4401 7 2 2 79163 83936
0 4402 5 1 1 83941
0 4403 7 1 2 83876 83942
0 4404 5 1 1 4403
0 4405 7 1 2 4399 4404
0 4406 5 1 1 4405
0 4407 7 1 2 67360 4406
0 4408 5 1 1 4407
0 4409 7 2 2 80922 79415
0 4410 5 1 1 83943
0 4411 7 1 2 78208 83944
0 4412 5 1 1 4411
0 4413 7 28 2 69495 82834
0 4414 5 3 1 83945
0 4415 7 1 2 83946 74746
0 4416 5 1 1 4415
0 4417 7 1 2 4412 4416
0 4418 5 1 1 4417
0 4419 7 1 2 81978 4418
0 4420 5 1 1 4419
0 4421 7 2 2 79794 80290
0 4422 7 2 2 66369 74060
0 4423 7 1 2 80041 83978
0 4424 7 1 2 83976 4423
0 4425 5 1 1 4424
0 4426 7 1 2 4420 4425
0 4427 5 1 1 4426
0 4428 7 1 2 73240 4427
0 4429 5 1 1 4428
0 4430 7 1 2 82102 79164
0 4431 5 1 1 4430
0 4432 7 10 2 64450 82771
0 4433 7 3 2 83280 83980
0 4434 5 1 1 83990
0 4435 7 1 2 4431 4434
0 4436 5 1 1 4435
0 4437 7 1 2 83855 4436
0 4438 5 1 1 4437
0 4439 7 1 2 4429 4438
0 4440 7 1 2 4408 4439
0 4441 5 1 1 4440
0 4442 7 1 2 67948 4441
0 4443 5 1 1 4442
0 4444 7 1 2 4375 4443
0 4445 5 1 1 4444
0 4446 7 1 2 74302 4445
0 4447 5 1 1 4446
0 4448 7 1 2 81484 83858
0 4449 5 1 1 4448
0 4450 7 9 2 67949 79416
0 4451 7 24 2 65313 70843
0 4452 5 2 1 84002
0 4453 7 4 2 73766 84003
0 4454 5 9 1 84028
0 4455 7 1 2 72488 84032
0 4456 5 3 1 4455
0 4457 7 2 2 67361 84041
0 4458 5 1 1 84044
0 4459 7 1 2 83993 84045
0 4460 5 1 1 4459
0 4461 7 1 2 4449 4460
0 4462 5 1 1 4461
0 4463 7 1 2 71415 4462
0 4464 5 1 1 4463
0 4465 7 6 2 69496 73642
0 4466 7 10 2 68926 64451
0 4467 7 3 2 63076 84052
0 4468 7 1 2 84046 84062
0 4469 5 1 1 4468
0 4470 7 21 2 67950 69300
0 4471 7 10 2 64649 84065
0 4472 7 1 2 74747 84086
0 4473 5 1 1 4472
0 4474 7 1 2 4469 4473
0 4475 5 1 1 4474
0 4476 7 1 2 73241 4475
0 4477 5 1 1 4476
0 4478 7 3 2 65666 72886
0 4479 7 1 2 83255 84096
0 4480 5 1 1 4479
0 4481 7 1 2 4477 4480
0 4482 5 1 1 4481
0 4483 7 1 2 71038 4482
0 4484 5 1 1 4483
0 4485 7 1 2 4464 4484
0 4486 5 1 1 4485
0 4487 7 1 2 66370 4486
0 4488 5 1 1 4487
0 4489 7 1 2 71416 74748
0 4490 5 1 1 4489
0 4491 7 9 2 81207 79287
0 4492 5 1 1 84099
0 4493 7 2 2 70227 84100
0 4494 5 1 1 84108
0 4495 7 1 2 4490 4494
0 4496 5 1 1 4495
0 4497 7 1 2 73242 4496
0 4498 5 1 1 4497
0 4499 7 1 2 71475 84097
0 4500 5 1 1 4499
0 4501 7 1 2 4498 4500
0 4502 5 1 1 4501
0 4503 7 1 2 78909 4502
0 4504 5 1 1 4503
0 4505 7 1 2 71417 83877
0 4506 5 1 1 4505
0 4507 7 1 2 70604 84101
0 4508 5 1 1 4507
0 4509 7 1 2 4506 4508
0 4510 5 1 1 4509
0 4511 7 3 2 63077 83886
0 4512 7 1 2 4510 84110
0 4513 5 1 1 4512
0 4514 7 1 2 4504 4513
0 4515 5 1 1 4514
0 4516 7 1 2 82835 4515
0 4517 5 1 1 4516
0 4518 7 1 2 4488 4517
0 4519 5 1 1 4518
0 4520 7 1 2 75758 4519
0 4521 5 1 1 4520
0 4522 7 1 2 63240 4521
0 4523 7 1 2 4447 4522
0 4524 5 1 1 4523
0 4525 7 1 2 4354 4524
0 4526 5 1 1 4525
0 4527 7 1 2 69928 4526
0 4528 5 1 1 4527
0 4529 7 5 2 70228 75130
0 4530 7 14 2 63241 69497
0 4531 5 1 1 84118
0 4532 7 3 2 84119 82229
0 4533 5 3 1 84132
0 4534 7 2 2 82595 80232
0 4535 7 1 2 68078 84138
0 4536 5 1 1 4535
0 4537 7 1 2 84135 4536
0 4538 5 1 1 4537
0 4539 7 2 2 84113 4538
0 4540 5 1 1 84140
0 4541 7 1 2 72510 84141
0 4542 5 1 1 4541
0 4543 7 11 2 68079 79417
0 4544 7 2 2 76842 84142
0 4545 5 1 1 84153
0 4546 7 14 2 68304 65314
0 4547 5 5 1 84155
0 4548 7 5 2 61996 72775
0 4549 7 1 2 84156 84174
0 4550 7 1 2 84154 4549
0 4551 5 1 1 4550
0 4552 7 1 2 4542 4551
0 4553 5 1 1 4552
0 4554 7 1 2 73243 4553
0 4555 5 1 1 4554
0 4556 7 2 2 78648 77343
0 4557 7 6 2 69709 79418
0 4558 7 5 2 67600 81543
0 4559 7 1 2 84181 84187
0 4560 7 1 2 84179 4559
0 4561 5 1 1 4560
0 4562 7 1 2 4540 4561
0 4563 5 1 1 4562
0 4564 7 1 2 71519 4563
0 4565 5 1 1 4564
0 4566 7 1 2 4555 4565
0 4567 5 1 1 4566
0 4568 7 1 2 61743 4567
0 4569 5 1 1 4568
0 4570 7 1 2 81146 84042
0 4571 5 1 1 4570
0 4572 7 9 2 66855 65315
0 4573 5 1 1 84192
0 4574 7 3 2 76313 84193
0 4575 7 2 2 79065 84201
0 4576 5 1 1 84204
0 4577 7 1 2 79319 84205
0 4578 5 1 1 4577
0 4579 7 1 2 4571 4578
0 4580 5 1 1 4579
0 4581 7 8 2 68305 69301
0 4582 7 5 2 68080 75589
0 4583 7 1 2 84206 84214
0 4584 7 1 2 4580 4583
0 4585 5 1 1 4584
0 4586 7 1 2 4569 4585
0 4587 5 1 1 4586
0 4588 7 1 2 76114 4587
0 4589 5 1 1 4588
0 4590 7 3 2 80962 75695
0 4591 7 1 2 82792 84219
0 4592 5 1 1 4591
0 4593 7 12 2 67601 69302
0 4594 5 1 1 84222
0 4595 7 3 2 82018 84223
0 4596 5 1 1 84234
0 4597 7 1 2 83916 4596
0 4598 5 5 1 4597
0 4599 7 1 2 77222 84237
0 4600 5 1 1 4599
0 4601 7 1 2 4592 4600
0 4602 5 1 1 4601
0 4603 7 7 2 65923 76685
0 4604 7 6 2 66856 81544
0 4605 7 7 2 67362 72746
0 4606 7 1 2 84249 84255
0 4607 7 1 2 84242 4606
0 4608 7 1 2 4602 4607
0 4609 5 1 1 4608
0 4610 7 1 2 65049 4609
0 4611 7 1 2 4589 4610
0 4612 5 1 1 4611
0 4613 7 1 2 66083 4612
0 4614 7 1 2 4528 4613
0 4615 5 1 1 4614
0 4616 7 6 2 64865 76686
0 4617 7 3 2 78033 84262
0 4618 7 2 2 80161 81528
0 4619 7 9 2 61251 67363
0 4620 7 2 2 74303 84273
0 4621 7 5 2 80963 82726
0 4622 7 1 2 84282 84284
0 4623 7 1 2 84271 4622
0 4624 7 1 2 84268 4623
0 4625 5 1 1 4624
0 4626 7 1 2 4615 4625
0 4627 5 1 1 4626
0 4628 7 1 2 71891 4627
0 4629 5 1 1 4628
0 4630 7 5 2 70229 71564
0 4631 5 3 1 84289
0 4632 7 12 2 62746 72014
0 4633 5 18 1 84297
0 4634 7 1 2 78533 84298
0 4635 5 1 1 4634
0 4636 7 2 2 72511 78585
0 4637 7 11 2 67602 68549
0 4638 7 1 2 84327 84329
0 4639 5 1 1 4638
0 4640 7 1 2 4635 4639
0 4641 5 1 1 4640
0 4642 7 1 2 83326 4641
0 4643 5 1 1 4642
0 4644 7 6 2 67603 65050
0 4645 5 1 1 84340
0 4646 7 2 2 72512 84341
0 4647 7 2 2 68550 79098
0 4648 7 1 2 84346 84348
0 4649 5 1 1 4648
0 4650 7 1 2 4643 4649
0 4651 5 1 1 4650
0 4652 7 1 2 76115 4651
0 4653 5 1 1 4652
0 4654 7 4 2 65924 80856
0 4655 7 1 2 84350 84330
0 4656 7 1 2 82027 4655
0 4657 5 1 1 4656
0 4658 7 1 2 4653 4657
0 4659 5 1 1 4658
0 4660 7 1 2 69303 4659
0 4661 5 1 1 4660
0 4662 7 18 2 62747 72601
0 4663 5 4 1 84354
0 4664 7 16 2 72097 84372
0 4665 7 6 2 65051 84376
0 4666 7 1 2 80845 83991
0 4667 7 1 2 84392 4666
0 4668 5 1 1 4667
0 4669 7 1 2 4661 4668
0 4670 5 1 1 4669
0 4671 7 1 2 66084 4670
0 4672 5 1 1 4671
0 4673 7 23 2 66371 64650
0 4674 5 1 1 84398
0 4675 7 1 2 84399 78709
0 4676 7 8 2 61252 66627
0 4677 7 12 2 68551 64452
0 4678 7 1 2 84421 84429
0 4679 7 1 2 4675 4678
0 4680 7 1 2 84393 4679
0 4681 5 1 1 4680
0 4682 7 1 2 4672 4681
0 4683 5 1 1 4682
0 4684 7 1 2 68081 4683
0 4685 5 1 1 4684
0 4686 7 1 2 76034 83922
0 4687 5 1 1 4686
0 4688 7 1 2 3970 4687
0 4689 5 1 1 4688
0 4690 7 12 2 69929 70844
0 4691 7 6 2 63242 64057
0 4692 7 2 2 84441 84453
0 4693 7 1 2 84459 83704
0 4694 7 1 2 4689 4693
0 4695 5 1 1 4694
0 4696 7 1 2 4685 4695
0 4697 5 1 1 4696
0 4698 7 1 2 67143 4697
0 4699 5 1 1 4698
0 4700 7 9 2 61744 67951
0 4701 7 7 2 61450 84461
0 4702 7 1 2 84133 84470
0 4703 5 1 1 4702
0 4704 7 14 2 64866 83076
0 4705 5 1 1 84477
0 4706 7 2 2 79419 84478
0 4707 7 1 2 76116 84491
0 4708 5 1 1 4707
0 4709 7 1 2 4703 4708
0 4710 5 1 1 4709
0 4711 7 12 2 64058 69930
0 4712 7 3 2 84493 81160
0 4713 7 1 2 83705 84505
0 4714 7 1 2 4710 4713
0 4715 5 1 1 4714
0 4716 7 1 2 4699 4715
0 4717 5 1 1 4716
0 4718 7 1 2 79315 4717
0 4719 5 1 1 4718
0 4720 7 1 2 83297 83603
0 4721 7 9 2 64059 64453
0 4722 7 2 2 68552 84508
0 4723 7 13 2 61997 63243
0 4724 5 1 1 84519
0 4725 7 4 2 80405 84520
0 4726 7 1 2 84517 84532
0 4727 7 1 2 4720 4726
0 4728 5 1 1 4727
0 4729 7 1 2 4719 4728
0 4730 5 1 1 4729
0 4731 7 1 2 84294 4730
0 4732 5 1 1 4731
0 4733 7 3 2 83887 84430
0 4734 7 2 2 79944 84536
0 4735 7 5 2 61253 68306
0 4736 7 1 2 79950 84541
0 4737 7 1 2 84285 4736
0 4738 7 1 2 84539 4737
0 4739 5 1 1 4738
0 4740 7 1 2 4732 4739
0 4741 7 1 2 4629 4740
0 4742 7 1 2 4260 4741
0 4743 7 1 2 3943 4742
0 4744 7 1 2 3252 4743
0 4745 5 1 1 4744
0 4746 7 1 2 69156 4745
0 4747 5 1 1 4746
0 4748 7 3 2 63896 74101
0 4749 5 3 1 84546
0 4750 7 1 2 67364 84549
0 4751 5 1 1 4750
0 4752 7 2 2 63707 2143
0 4753 5 1 1 84552
0 4754 7 1 2 4751 84553
0 4755 5 1 1 4754
0 4756 7 1 2 73643 4755
0 4757 5 1 1 4756
0 4758 7 10 2 62748 63897
0 4759 5 9 1 84554
0 4760 7 7 2 62502 84555
0 4761 5 4 1 84573
0 4762 7 1 2 64060 84574
0 4763 5 1 1 4762
0 4764 7 1 2 67144 4763
0 4765 5 1 1 4764
0 4766 7 11 2 65316 73374
0 4767 5 15 1 84584
0 4768 7 2 2 84595 77731
0 4769 5 1 1 84610
0 4770 7 3 2 63708 71293
0 4771 5 8 1 84612
0 4772 7 1 2 70230 84613
0 4773 5 3 1 4772
0 4774 7 1 2 72815 84623
0 4775 5 1 1 4774
0 4776 7 1 2 84611 4775
0 4777 7 1 2 4765 4776
0 4778 5 1 1 4777
0 4779 7 1 2 70845 4778
0 4780 5 1 1 4779
0 4781 7 1 2 4757 4780
0 4782 5 1 1 4781
0 4783 7 1 2 77655 4782
0 4784 5 1 1 4783
0 4785 7 1 2 76972 72776
0 4786 5 1 1 4785
0 4787 7 2 2 65317 78663
0 4788 7 1 2 68553 84626
0 4789 5 1 1 4788
0 4790 7 1 2 72868 4789
0 4791 5 1 1 4790
0 4792 7 1 2 69931 4791
0 4793 5 1 1 4792
0 4794 7 1 2 4786 4793
0 4795 5 1 1 4794
0 4796 7 1 2 67145 65925
0 4797 7 1 2 4795 4796
0 4798 5 1 1 4797
0 4799 7 1 2 4784 4798
0 4800 5 1 1 4799
0 4801 7 1 2 65667 4800
0 4802 5 1 1 4801
0 4803 7 5 2 68770 74574
0 4804 5 1 1 84628
0 4805 7 1 2 67365 84629
0 4806 5 1 1 4805
0 4807 7 1 2 75973 4806
0 4808 5 3 1 4807
0 4809 7 1 2 70846 84633
0 4810 5 1 1 4809
0 4811 7 3 2 74061 72259
0 4812 5 7 1 84636
0 4813 7 1 2 78167 84639
0 4814 5 1 1 4813
0 4815 7 1 2 84624 4814
0 4816 5 1 1 4815
0 4817 7 21 2 67604 72513
0 4818 5 9 1 84646
0 4819 7 2 2 75340 84647
0 4820 5 1 1 84676
0 4821 7 2 2 62316 74565
0 4822 5 6 1 84678
0 4823 7 1 2 76331 73375
0 4824 7 1 2 74996 4823
0 4825 7 1 2 84680 4824
0 4826 5 1 1 4825
0 4827 7 1 2 4820 4826
0 4828 7 1 2 4816 4827
0 4829 7 1 2 4810 4828
0 4830 5 1 1 4829
0 4831 7 1 2 77656 4830
0 4832 5 1 1 4831
0 4833 7 1 2 4802 4832
0 4834 5 1 1 4833
0 4835 7 1 2 68307 4834
0 4836 5 1 1 4835
0 4837 7 4 2 67366 74062
0 4838 5 2 1 84686
0 4839 7 1 2 70231 84690
0 4840 5 2 1 4839
0 4841 7 1 2 83753 84692
0 4842 5 1 1 4841
0 4843 7 3 2 65318 82497
0 4844 5 2 1 84694
0 4845 7 1 2 4842 84697
0 4846 5 1 1 4845
0 4847 7 2 2 79817 79573
0 4848 5 1 1 84699
0 4849 7 1 2 65926 84700
0 4850 7 1 2 4846 4849
0 4851 5 1 1 4850
0 4852 7 1 2 4836 4851
0 4853 5 1 1 4852
0 4854 7 1 2 83027 4853
0 4855 5 1 1 4854
0 4856 7 5 2 62317 72911
0 4857 5 2 1 84701
0 4858 7 8 2 68082 64061
0 4859 5 1 1 84708
0 4860 7 4 2 63898 74257
0 4861 7 2 2 84709 84716
0 4862 7 1 2 84702 84720
0 4863 5 1 1 4862
0 4864 7 2 2 67605 83754
0 4865 5 1 1 84722
0 4866 7 2 2 78162 84723
0 4867 5 2 1 84724
0 4868 7 1 2 66857 84725
0 4869 5 1 1 4868
0 4870 7 2 2 63474 77895
0 4871 5 1 1 84728
0 4872 7 4 2 65927 71192
0 4873 5 1 1 84730
0 4874 7 2 2 73376 76284
0 4875 7 6 2 127 84734
0 4876 5 3 1 84736
0 4877 7 1 2 68927 84737
0 4878 5 1 1 4877
0 4879 7 1 2 4873 4878
0 4880 5 4 1 4879
0 4881 7 1 2 71801 84745
0 4882 5 1 1 4881
0 4883 7 1 2 4871 4882
0 4884 5 1 1 4883
0 4885 7 1 2 66858 4884
0 4886 5 1 1 4885
0 4887 7 2 2 66859 74599
0 4888 5 1 1 84749
0 4889 7 6 2 64062 73820
0 4890 7 1 2 80517 84751
0 4891 5 1 1 4890
0 4892 7 1 2 4888 4891
0 4893 5 1 1 4892
0 4894 7 1 2 67146 4893
0 4895 5 1 1 4894
0 4896 7 4 2 62503 73821
0 4897 7 8 2 64063 65928
0 4898 5 2 1 84761
0 4899 7 1 2 73679 84762
0 4900 7 1 2 84757 4899
0 4901 5 2 1 4900
0 4902 7 1 2 4895 84771
0 4903 7 1 2 4886 4902
0 4904 5 1 1 4903
0 4905 7 1 2 65668 4904
0 4906 5 1 1 4905
0 4907 7 1 2 4869 4906
0 4908 5 1 1 4907
0 4909 7 1 2 63244 4908
0 4910 5 1 1 4909
0 4911 7 1 2 4863 4910
0 4912 5 1 1 4911
0 4913 7 1 2 65052 4912
0 4914 5 1 1 4913
0 4915 7 2 2 70847 79891
0 4916 7 2 2 80466 81577
0 4917 5 1 1 84775
0 4918 7 1 2 84773 84776
0 4919 5 1 1 4918
0 4920 7 28 2 66860 63245
0 4921 7 2 2 68928 84777
0 4922 7 5 2 65929 74854
0 4923 7 2 2 84807 73377
0 4924 7 1 2 84805 84812
0 4925 5 1 1 4924
0 4926 7 1 2 4919 4925
0 4927 5 1 1 4926
0 4928 7 1 2 67606 4927
0 4929 5 1 1 4928
0 4930 7 7 2 63246 68771
0 4931 7 4 2 78649 84814
0 4932 7 1 2 84808 84821
0 4933 5 1 1 4932
0 4934 7 1 2 4929 4933
0 4935 5 1 1 4934
0 4936 7 1 2 78186 4935
0 4937 5 1 1 4936
0 4938 7 1 2 4914 4937
0 4939 5 1 1 4938
0 4940 7 1 2 70232 4939
0 4941 5 1 1 4940
0 4942 7 5 2 73600 77917
0 4943 5 3 1 84825
0 4944 7 1 2 76517 84826
0 4945 5 1 1 4944
0 4946 7 4 2 62749 84494
0 4947 7 1 2 84833 77118
0 4948 5 1 1 4947
0 4949 7 1 2 4945 4948
0 4950 5 1 1 4949
0 4951 7 1 2 68083 76453
0 4952 7 1 2 4950 4951
0 4953 5 1 1 4952
0 4954 7 1 2 70233 71657
0 4955 5 4 1 4954
0 4956 7 4 2 68084 70848
0 4957 7 2 2 78055 84841
0 4958 7 1 2 84837 84845
0 4959 5 1 1 4958
0 4960 7 6 2 65053 72441
0 4961 7 2 2 63247 73726
0 4962 7 1 2 84847 84853
0 4963 5 1 1 4962
0 4964 7 1 2 4959 4963
0 4965 5 1 1 4964
0 4966 7 1 2 71892 4965
0 4967 5 1 1 4966
0 4968 7 13 2 67147 63248
0 4969 7 1 2 74879 84855
0 4970 7 1 2 80857 76687
0 4971 7 1 2 4969 4970
0 4972 5 1 1 4971
0 4973 7 1 2 4967 4972
0 4974 7 1 2 4953 4973
0 4975 5 1 1 4974
0 4976 7 1 2 61998 4975
0 4977 5 1 1 4976
0 4978 7 1 2 77827 72296
0 4979 5 4 1 4978
0 4980 7 1 2 67607 84868
0 4981 5 3 1 4980
0 4982 7 1 2 71658 82179
0 4983 5 1 1 4982
0 4984 7 1 2 70849 4983
0 4985 5 1 1 4984
0 4986 7 1 2 84872 4985
0 4987 5 1 1 4986
0 4988 7 1 2 68308 4987
0 4989 5 1 1 4988
0 4990 7 3 2 67367 84331
0 4991 7 3 2 72260 72747
0 4992 5 1 1 84878
0 4993 7 1 2 84875 84879
0 4994 5 1 1 4993
0 4995 7 1 2 81164 84640
0 4996 5 1 1 4995
0 4997 7 1 2 71193 4996
0 4998 5 1 1 4997
0 4999 7 5 2 70605 74102
0 5000 5 7 1 84881
0 5001 7 1 2 75081 79929
0 5002 7 1 2 84886 5001
0 5003 5 1 1 5002
0 5004 7 1 2 4998 5003
0 5005 5 1 1 5004
0 5006 7 1 2 67148 5005
0 5007 5 1 1 5006
0 5008 7 1 2 4994 5007
0 5009 7 1 2 4989 5008
0 5010 5 1 1 5009
0 5011 7 1 2 69932 5010
0 5012 5 1 1 5011
0 5013 7 4 2 67368 70850
0 5014 5 2 1 84893
0 5015 7 2 2 84894 72315
0 5016 5 8 1 84899
0 5017 7 3 2 84641 84901
0 5018 5 3 1 84909
0 5019 7 1 2 79010 84912
0 5020 5 1 1 5019
0 5021 7 1 2 5012 5020
0 5022 5 1 1 5021
0 5023 7 1 2 65319 5022
0 5024 5 1 1 5023
0 5025 7 3 2 69933 72261
0 5026 5 1 1 84915
0 5027 7 8 2 62750 73767
0 5028 5 4 1 84918
0 5029 7 1 2 84442 84926
0 5030 5 1 1 5029
0 5031 7 1 2 5026 5030
0 5032 5 1 1 5031
0 5033 7 1 2 74855 5032
0 5034 5 1 1 5033
0 5035 7 3 2 70606 72098
0 5036 5 3 1 84930
0 5037 7 1 2 82961 84931
0 5038 5 1 1 5037
0 5039 7 1 2 5034 5038
0 5040 5 1 1 5039
0 5041 7 1 2 65320 5040
0 5042 5 1 1 5041
0 5043 7 3 2 70851 73937
0 5044 5 1 1 84936
0 5045 7 1 2 5044 84933
0 5046 5 2 1 5045
0 5047 7 9 2 69934 71893
0 5048 5 1 1 84941
0 5049 7 1 2 68309 84942
0 5050 7 1 2 84939 5049
0 5051 5 1 1 5050
0 5052 7 1 2 5042 5051
0 5053 5 1 1 5052
0 5054 7 1 2 73378 5053
0 5055 5 1 1 5054
0 5056 7 4 2 76285 75741
0 5057 7 3 2 71802 78436
0 5058 5 2 1 84954
0 5059 7 5 2 68310 70852
0 5060 5 2 1 84959
0 5061 7 1 2 84957 84960
0 5062 7 1 2 82182 5061
0 5063 7 1 2 84950 5062
0 5064 5 1 1 5063
0 5065 7 5 2 68554 71194
0 5066 5 1 1 84966
0 5067 7 1 2 63475 5066
0 5068 5 4 1 5067
0 5069 7 1 2 1246 82183
0 5070 7 5 2 84971 5069
0 5071 5 1 1 84975
0 5072 7 3 2 70607 75536
0 5073 5 9 1 84980
0 5074 7 1 2 68929 76332
0 5075 7 1 2 84983 5074
0 5076 7 1 2 84976 5075
0 5077 5 1 1 5076
0 5078 7 1 2 5064 5077
0 5079 5 1 1 5078
0 5080 7 1 2 69935 5079
0 5081 5 1 1 5080
0 5082 7 1 2 5055 5081
0 5083 7 1 2 5024 5082
0 5084 5 1 1 5083
0 5085 7 1 2 84778 5084
0 5086 5 1 1 5085
0 5087 7 1 2 4977 5086
0 5088 7 1 2 4941 5087
0 5089 5 1 1 5088
0 5090 7 1 2 66628 5089
0 5091 5 1 1 5090
0 5092 7 1 2 4855 5091
0 5093 5 1 1 5092
0 5094 7 1 2 67952 5093
0 5095 5 1 1 5094
0 5096 7 4 2 72514 80768
0 5097 7 1 2 84992 82712
0 5098 7 5 2 66629 79951
0 5099 7 5 2 67369 80133
0 5100 7 1 2 84996 85001
0 5101 7 1 2 5097 5100
0 5102 5 1 1 5101
0 5103 7 1 2 5095 5102
0 5104 5 1 1 5103
0 5105 7 1 2 82103 5104
0 5106 5 1 1 5105
0 5107 7 1 2 77544 73751
0 5108 5 1 1 5107
0 5109 7 1 2 65321 2081
0 5110 5 1 1 5109
0 5111 7 1 2 61999 74713
0 5112 7 1 2 5110 5111
0 5113 5 1 1 5112
0 5114 7 1 2 5108 5113
0 5115 5 1 1 5114
0 5116 7 1 2 68085 5115
0 5117 5 1 1 5116
0 5118 7 1 2 82572 79481
0 5119 5 1 1 5118
0 5120 7 1 2 5117 5119
0 5121 5 1 1 5120
0 5122 7 1 2 61745 5121
0 5123 5 1 1 5122
0 5124 7 10 2 62504 68086
0 5125 5 1 1 85006
0 5126 7 3 2 73601 85007
0 5127 7 1 2 79766 85016
0 5128 5 1 1 5127
0 5129 7 5 2 66630 84521
0 5130 7 11 2 67149 65322
0 5131 5 3 1 85024
0 5132 7 1 2 85019 85025
0 5133 5 1 1 5132
0 5134 7 1 2 5128 5133
0 5135 5 1 1 5134
0 5136 7 1 2 78437 5135
0 5137 5 1 1 5136
0 5138 7 1 2 65054 5137
0 5139 7 1 2 5123 5138
0 5140 5 1 1 5139
0 5141 7 2 2 67150 83077
0 5142 7 2 2 73244 1216
0 5143 7 1 2 77980 85040
0 5144 5 2 1 5143
0 5145 7 1 2 74668 85042
0 5146 5 1 1 5145
0 5147 7 1 2 85038 5146
0 5148 5 1 1 5147
0 5149 7 2 2 72365 75893
0 5150 5 1 1 85044
0 5151 7 1 2 81433 85045
0 5152 5 1 1 5151
0 5153 7 1 2 5148 5152
0 5154 5 1 1 5153
0 5155 7 1 2 66861 5154
0 5156 5 1 1 5155
0 5157 7 2 2 84157 75023
0 5158 5 1 1 85046
0 5159 7 1 2 83028 85047
0 5160 5 1 1 5159
0 5161 7 1 2 69936 5160
0 5162 7 1 2 5156 5161
0 5163 5 1 1 5162
0 5164 7 1 2 68555 5163
0 5165 7 1 2 5140 5164
0 5166 5 1 1 5165
0 5167 7 7 2 67370 69937
0 5168 7 2 2 85048 83755
0 5169 7 3 2 61746 81545
0 5170 5 1 1 85057
0 5171 7 1 2 63476 85035
0 5172 5 5 1 5171
0 5173 7 1 2 81434 85060
0 5174 5 1 1 5173
0 5175 7 1 2 5170 5174
0 5176 5 1 1 5175
0 5177 7 1 2 85055 5176
0 5178 5 1 1 5177
0 5179 7 14 2 65669 73379
0 5180 5 10 1 85065
0 5181 7 2 2 79767 83537
0 5182 5 1 1 85089
0 5183 7 1 2 81435 79311
0 5184 5 1 1 5183
0 5185 7 1 2 5182 5184
0 5186 5 1 1 5185
0 5187 7 1 2 85066 5186
0 5188 5 1 1 5187
0 5189 7 2 2 74673 75894
0 5190 5 4 1 85091
0 5191 7 1 2 65055 81436
0 5192 7 1 2 85092 5191
0 5193 5 1 1 5192
0 5194 7 1 2 5188 5193
0 5195 5 1 1 5194
0 5196 7 1 2 70234 5195
0 5197 5 1 1 5196
0 5198 7 1 2 5178 5197
0 5199 5 1 1 5198
0 5200 7 1 2 66862 5199
0 5201 5 1 1 5200
0 5202 7 11 2 61747 70235
0 5203 7 1 2 75024 85097
0 5204 7 1 2 83007 5203
0 5205 5 1 1 5204
0 5206 7 1 2 5201 5205
0 5207 7 1 2 5166 5206
0 5208 5 1 1 5207
0 5209 7 1 2 65930 5208
0 5210 5 1 1 5209
0 5211 7 1 2 63249 74304
0 5212 5 3 1 5211
0 5213 7 2 2 63477 84842
0 5214 5 1 1 85111
0 5215 7 1 2 85108 5214
0 5216 5 1 1 5215
0 5217 7 1 2 85067 5216
0 5218 5 1 1 5217
0 5219 7 1 2 68311 84822
0 5220 5 1 1 5219
0 5221 7 1 2 5218 5220
0 5222 5 1 1 5221
0 5223 7 1 2 80865 83490
0 5224 7 1 2 5222 5223
0 5225 5 1 1 5224
0 5226 7 1 2 5210 5225
0 5227 5 1 1 5226
0 5228 7 1 2 61451 5227
0 5229 5 1 1 5228
0 5230 7 2 2 70236 85079
0 5231 5 3 1 85113
0 5232 7 14 2 62318 63250
0 5233 7 6 2 63709 85118
0 5234 7 4 2 69938 77182
0 5235 7 1 2 81180 606
0 5236 7 1 2 85138 5235
0 5237 7 1 2 85132 5236
0 5238 7 1 2 85115 5237
0 5239 5 1 1 5238
0 5240 7 1 2 5229 5239
0 5241 5 1 1 5240
0 5242 7 1 2 68930 5241
0 5243 5 1 1 5242
0 5244 7 3 2 68087 75465
0 5245 7 5 2 73845 73768
0 5246 5 1 1 85145
0 5247 7 2 2 63899 80546
0 5248 5 1 1 85150
0 5249 7 1 2 62505 85151
0 5250 5 2 1 5249
0 5251 7 1 2 5246 85152
0 5252 5 1 1 5251
0 5253 7 1 2 62751 5252
0 5254 5 2 1 5253
0 5255 7 5 2 71719 73284
0 5256 5 3 1 85156
0 5257 7 1 2 85154 85161
0 5258 5 2 1 5257
0 5259 7 2 2 76454 85164
0 5260 7 1 2 85142 85166
0 5261 5 1 1 5260
0 5262 7 3 2 68772 84984
0 5263 5 1 1 85168
0 5264 7 5 2 61748 83402
0 5265 7 1 2 81188 85171
0 5266 7 1 2 85169 5265
0 5267 5 1 1 5266
0 5268 7 1 2 5261 5267
0 5269 5 1 1 5268
0 5270 7 1 2 65056 5269
0 5271 5 1 1 5270
0 5272 7 3 2 62000 84596
0 5273 5 1 1 85176
0 5274 7 2 2 77551 85177
0 5275 5 1 1 85179
0 5276 7 13 2 62752 68088
0 5277 7 2 2 71631 85181
0 5278 7 4 2 69939 74171
0 5279 7 1 2 66631 85196
0 5280 7 1 2 85194 5279
0 5281 7 1 2 85180 5280
0 5282 5 1 1 5281
0 5283 7 1 2 5271 5282
0 5284 5 1 1 5283
0 5285 7 1 2 61452 5284
0 5286 5 1 1 5285
0 5287 7 1 2 5243 5286
0 5288 5 1 1 5287
0 5289 7 1 2 63078 5288
0 5290 5 1 1 5289
0 5291 7 3 2 63478 77066
0 5292 5 1 1 85200
0 5293 7 4 2 62319 78143
0 5294 5 1 1 85203
0 5295 7 1 2 77067 85204
0 5296 5 1 1 5295
0 5297 7 1 2 5292 5296
0 5298 5 4 1 5297
0 5299 7 1 2 65323 85207
0 5300 5 1 1 5299
0 5301 7 6 2 62506 73680
0 5302 5 5 1 85211
0 5303 7 1 2 79596 85212
0 5304 5 2 1 5303
0 5305 7 1 2 5300 85222
0 5306 5 1 1 5305
0 5307 7 3 2 65931 83218
0 5308 7 3 2 62001 78438
0 5309 7 1 2 85227 84471
0 5310 7 1 2 85224 5309
0 5311 7 1 2 5306 5310
0 5312 5 1 1 5311
0 5313 7 1 2 5290 5312
0 5314 5 1 1 5313
0 5315 7 1 2 64454 5314
0 5316 5 1 1 5315
0 5317 7 1 2 64867 5316
0 5318 7 1 2 5106 5317
0 5319 5 1 1 5318
0 5320 7 3 2 68089 71894
0 5321 7 4 2 67151 75395
0 5322 7 1 2 72816 85116
0 5323 5 1 1 5322
0 5324 7 1 2 71195 84887
0 5325 5 2 1 5324
0 5326 7 1 2 5323 85237
0 5327 5 1 1 5326
0 5328 7 1 2 85233 5327
0 5329 5 1 1 5328
0 5330 7 5 2 67152 73380
0 5331 5 11 1 85239
0 5332 7 5 2 70608 85244
0 5333 5 1 1 85255
0 5334 7 10 2 66632 70237
0 5335 7 1 2 74063 85260
0 5336 7 1 2 85256 5335
0 5337 5 1 1 5336
0 5338 7 1 2 5329 5337
0 5339 5 1 1 5338
0 5340 7 1 2 65932 5339
0 5341 5 1 1 5340
0 5342 7 3 2 71196 72817
0 5343 5 2 1 85270
0 5344 7 1 2 70238 85273
0 5345 5 1 1 5344
0 5346 7 1 2 85234 5345
0 5347 5 1 1 5346
0 5348 7 4 2 70239 71148
0 5349 7 1 2 75611 85275
0 5350 5 1 1 5349
0 5351 7 1 2 5347 5350
0 5352 5 1 1 5351
0 5353 7 1 2 65670 5352
0 5354 5 1 1 5353
0 5355 7 5 2 62507 74103
0 5356 5 6 1 85279
0 5357 7 3 2 63900 85280
0 5358 5 3 1 85290
0 5359 7 2 2 75396 85026
0 5360 5 1 1 85296
0 5361 7 1 2 85293 85297
0 5362 5 1 1 5361
0 5363 7 1 2 5354 5362
0 5364 7 1 2 5341 5363
0 5365 5 1 1 5364
0 5366 7 1 2 68556 5365
0 5367 5 1 1 5366
0 5368 7 1 2 85261 74482
0 5369 5 1 1 5368
0 5370 7 2 2 84377 79989
0 5371 5 1 1 85298
0 5372 7 1 2 77910 5371
0 5373 5 2 1 5372
0 5374 7 2 2 65324 85300
0 5375 7 1 2 75397 85302
0 5376 5 1 1 5375
0 5377 7 1 2 5369 5376
0 5378 7 1 2 5367 5377
0 5379 5 1 1 5378
0 5380 7 1 2 85230 5379
0 5381 5 1 1 5380
0 5382 7 3 2 77999 78362
0 5383 5 4 1 85304
0 5384 7 2 2 68773 85305
0 5385 5 1 1 85311
0 5386 7 3 2 82573 82611
0 5387 7 1 2 74771 85313
0 5388 7 1 2 85312 5387
0 5389 5 1 1 5388
0 5390 7 1 2 5381 5389
0 5391 5 1 1 5390
0 5392 7 1 2 63079 5391
0 5393 5 1 1 5392
0 5394 7 5 2 71803 82363
0 5395 7 1 2 80193 85316
0 5396 7 1 2 77455 5395
0 5397 5 1 1 5396
0 5398 7 1 2 5393 5397
0 5399 5 1 1 5398
0 5400 7 1 2 65057 5399
0 5401 5 1 1 5400
0 5402 7 8 2 63251 84462
0 5403 7 8 2 64064 73938
0 5404 5 1 1 85329
0 5405 7 1 2 71135 5404
0 5406 5 4 1 5405
0 5407 7 2 2 73381 85337
0 5408 5 2 1 85341
0 5409 7 3 2 65671 71110
0 5410 5 1 1 85345
0 5411 7 2 2 62753 84838
0 5412 5 1 1 85348
0 5413 7 1 2 5410 5412
0 5414 7 1 2 85343 5413
0 5415 5 1 1 5414
0 5416 7 1 2 69940 5415
0 5417 5 1 1 5416
0 5418 7 11 2 62754 68774
0 5419 5 1 1 85350
0 5420 7 5 2 67371 85351
0 5421 7 2 2 73769 85361
0 5422 5 1 1 85366
0 5423 7 1 2 73846 85367
0 5424 5 1 1 5423
0 5425 7 1 2 5417 5424
0 5426 5 1 1 5425
0 5427 7 1 2 71895 5426
0 5428 5 1 1 5427
0 5429 7 1 2 70240 76354
0 5430 5 2 1 5429
0 5431 7 2 2 1041 85368
0 5432 7 1 2 67608 85370
0 5433 5 2 1 5432
0 5434 7 1 2 73786 74137
0 5435 5 1 1 5434
0 5436 7 1 2 85372 5435
0 5437 5 1 1 5436
0 5438 7 1 2 73382 5437
0 5439 5 2 1 5438
0 5440 7 10 2 64065 65325
0 5441 5 3 1 85376
0 5442 7 1 2 85386 84642
0 5443 5 1 1 5442
0 5444 7 1 2 71197 5443
0 5445 5 1 1 5444
0 5446 7 1 2 83733 80077
0 5447 5 1 1 5446
0 5448 7 1 2 5445 5447
0 5449 7 1 2 85374 5448
0 5450 5 1 1 5449
0 5451 7 1 2 69941 5450
0 5452 5 1 1 5451
0 5453 7 1 2 5428 5452
0 5454 5 1 1 5453
0 5455 7 1 2 66863 5454
0 5456 5 1 1 5455
0 5457 7 3 2 76241 83203
0 5458 5 1 1 85389
0 5459 7 1 2 74772 74462
0 5460 7 1 2 85390 5459
0 5461 5 1 1 5460
0 5462 7 1 2 5456 5461
0 5463 5 1 1 5462
0 5464 7 1 2 85321 5463
0 5465 5 1 1 5464
0 5466 7 1 2 5401 5465
0 5467 5 1 1 5466
0 5468 7 1 2 68312 5467
0 5469 5 1 1 5468
0 5470 7 4 2 65933 76877
0 5471 7 3 2 74064 85392
0 5472 5 3 1 85396
0 5473 7 1 2 85399 76871
0 5474 5 1 1 5473
0 5475 7 1 2 63479 5474
0 5476 5 1 1 5475
0 5477 7 1 2 72297 79687
0 5478 5 8 1 5477
0 5479 7 1 2 85402 75362
0 5480 5 1 1 5479
0 5481 7 1 2 85375 5480
0 5482 5 1 1 5481
0 5483 7 1 2 69942 5482
0 5484 5 1 1 5483
0 5485 7 1 2 5476 5484
0 5486 5 1 1 5485
0 5487 7 1 2 75398 83701
0 5488 7 1 2 5486 5487
0 5489 5 1 1 5488
0 5490 7 1 2 5469 5489
0 5491 5 1 1 5490
0 5492 7 1 2 61453 5491
0 5493 5 1 1 5492
0 5494 7 17 2 66372 63252
0 5495 5 1 1 85410
0 5496 7 6 2 69943 84585
0 5497 7 1 2 76831 85427
0 5498 5 1 1 5497
0 5499 7 1 2 84848 85235
0 5500 5 1 1 5499
0 5501 7 1 2 5498 5500
0 5502 5 1 1 5501
0 5503 7 1 2 71149 5502
0 5504 5 1 1 5503
0 5505 7 1 2 74722 85387
0 5506 5 1 1 5505
0 5507 7 1 2 85068 5506
0 5508 5 1 1 5507
0 5509 7 1 2 72232 5508
0 5510 5 1 1 5509
0 5511 7 1 2 63480 5510
0 5512 5 1 1 5511
0 5513 7 2 2 71720 84752
0 5514 5 1 1 85433
0 5515 7 1 2 70853 85434
0 5516 5 1 1 5515
0 5517 7 1 2 69944 5516
0 5518 7 1 2 5512 5517
0 5519 5 1 1 5518
0 5520 7 1 2 65326 84927
0 5521 5 2 1 5520
0 5522 7 1 2 70854 74349
0 5523 7 1 2 73285 5522
0 5524 7 1 2 85435 5523
0 5525 5 1 1 5524
0 5526 7 1 2 65058 743
0 5527 7 1 2 5525 5526
0 5528 5 1 1 5527
0 5529 7 1 2 71771 5528
0 5530 7 1 2 5519 5529
0 5531 5 1 1 5530
0 5532 7 1 2 5504 5531
0 5533 5 1 1 5532
0 5534 7 1 2 63080 5533
0 5535 5 1 1 5534
0 5536 7 2 2 78056 85165
0 5537 7 1 2 76767 85437
0 5538 5 1 1 5537
0 5539 7 1 2 5535 5538
0 5540 5 1 1 5539
0 5541 7 1 2 63710 5540
0 5542 5 1 1 5541
0 5543 7 4 2 63901 75845
0 5544 7 3 2 80701 85439
0 5545 7 1 2 70855 76661
0 5546 7 1 2 85436 5545
0 5547 7 1 2 85443 5546
0 5548 5 1 1 5547
0 5549 7 1 2 5542 5548
0 5550 5 1 1 5549
0 5551 7 1 2 85411 5550
0 5552 5 1 1 5551
0 5553 7 1 2 5493 5552
0 5554 5 1 1 5553
0 5555 7 1 2 64455 5554
0 5556 5 1 1 5555
0 5557 7 4 2 67372 65672
0 5558 5 4 1 85446
0 5559 7 4 2 72366 85447
0 5560 5 2 1 85454
0 5561 7 2 2 65673 83734
0 5562 5 1 1 85460
0 5563 7 1 2 84597 5562
0 5564 5 4 1 5563
0 5565 7 1 2 68557 85462
0 5566 5 1 1 5565
0 5567 7 1 2 85458 5566
0 5568 5 1 1 5567
0 5569 7 1 2 67153 5568
0 5570 5 1 1 5569
0 5571 7 2 2 84967 76688
0 5572 5 1 1 85466
0 5573 7 1 2 5570 5572
0 5574 5 1 1 5573
0 5575 7 1 2 76289 5574
0 5576 5 1 1 5575
0 5577 7 12 2 70609 73383
0 5578 5 1 1 85468
0 5579 7 2 2 85469 84681
0 5580 5 1 1 85480
0 5581 7 1 2 72442 82184
0 5582 5 1 1 5581
0 5583 7 1 2 5580 5582
0 5584 5 1 1 5583
0 5585 7 1 2 83484 5584
0 5586 5 1 1 5585
0 5587 7 1 2 5576 5586
0 5588 5 1 1 5587
0 5589 7 1 2 68313 5588
0 5590 5 1 1 5589
0 5591 7 3 2 76878 84332
0 5592 7 1 2 83763 82502
0 5593 5 2 1 5592
0 5594 7 1 2 82148 85485
0 5595 7 1 2 85482 5594
0 5596 5 1 1 5595
0 5597 7 1 2 5590 5596
0 5598 5 1 1 5597
0 5599 7 1 2 66864 5598
0 5600 5 1 1 5599
0 5601 7 1 2 78664 84158
0 5602 7 1 2 79984 5601
0 5603 7 1 2 83485 5602
0 5604 5 1 1 5603
0 5605 7 1 2 5600 5604
0 5606 5 1 1 5605
0 5607 7 1 2 72099 5606
0 5608 5 1 1 5607
0 5609 7 1 2 67154 84627
0 5610 5 1 1 5609
0 5611 7 1 2 72869 5610
0 5612 5 1 1 5611
0 5613 7 1 2 83204 5612
0 5614 5 1 1 5613
0 5615 7 6 2 70856 76930
0 5616 5 1 1 85487
0 5617 7 1 2 75371 85488
0 5618 5 1 1 5617
0 5619 7 1 2 5614 5618
0 5620 5 1 1 5619
0 5621 7 1 2 66633 5620
0 5622 5 1 1 5621
0 5623 7 6 2 65934 73384
0 5624 7 1 2 67609 77552
0 5625 7 1 2 85493 5624
0 5626 7 1 2 76203 5625
0 5627 5 1 1 5626
0 5628 7 1 2 5622 5627
0 5629 5 1 1 5628
0 5630 7 1 2 68931 5629
0 5631 5 1 1 5630
0 5632 7 5 2 66634 70857
0 5633 7 1 2 84495 85499
0 5634 5 1 1 5633
0 5635 7 3 2 65327 82047
0 5636 7 1 2 65059 85504
0 5637 5 1 1 5636
0 5638 7 1 2 5634 5637
0 5639 5 1 1 5638
0 5640 7 1 2 73385 5639
0 5641 5 1 1 5640
0 5642 7 1 2 79892 77553
0 5643 7 3 2 83735 5642
0 5644 5 1 1 85507
0 5645 7 1 2 65060 75696
0 5646 7 1 2 85508 5645
0 5647 5 1 1 5646
0 5648 7 1 2 5641 5647
0 5649 5 1 1 5648
0 5650 7 1 2 66865 5649
0 5651 5 1 1 5650
0 5652 7 1 2 5631 5651
0 5653 5 1 1 5652
0 5654 7 1 2 65674 5653
0 5655 5 1 1 5654
0 5656 7 3 2 72015 77554
0 5657 7 1 2 75466 85510
0 5658 5 1 1 5657
0 5659 7 6 2 68775 77566
0 5660 5 1 1 85513
0 5661 7 1 2 71198 72515
0 5662 5 3 1 5661
0 5663 7 1 2 62320 85519
0 5664 5 1 1 5663
0 5665 7 2 2 63902 83364
0 5666 5 5 1 85522
0 5667 7 2 2 67610 85524
0 5668 7 1 2 5664 85529
0 5669 5 1 1 5668
0 5670 7 1 2 5660 5669
0 5671 5 1 1 5670
0 5672 7 1 2 65328 75399
0 5673 7 1 2 5671 5672
0 5674 5 1 1 5673
0 5675 7 1 2 5658 5674
0 5676 5 1 1 5675
0 5677 7 1 2 65061 5676
0 5678 5 1 1 5677
0 5679 7 1 2 72298 74518
0 5680 5 5 1 5679
0 5681 7 1 2 67373 85531
0 5682 5 1 1 5681
0 5683 7 3 2 70858 77421
0 5684 5 1 1 85536
0 5685 7 1 2 4992 5684
0 5686 7 1 2 5682 5685
0 5687 5 1 1 5686
0 5688 7 1 2 66635 77657
0 5689 7 1 2 5687 5688
0 5690 5 1 1 5689
0 5691 7 1 2 5678 5690
0 5692 7 1 2 5655 5691
0 5693 5 1 1 5692
0 5694 7 1 2 68558 5693
0 5695 5 1 1 5694
0 5696 7 1 2 79893 72443
0 5697 5 2 1 5696
0 5698 7 1 2 77555 85470
0 5699 5 1 1 5698
0 5700 7 1 2 85539 5699
0 5701 5 1 1 5700
0 5702 7 1 2 72516 5701
0 5703 5 1 1 5702
0 5704 7 6 2 67374 73245
0 5705 5 6 1 85541
0 5706 7 6 2 71565 85547
0 5707 5 18 1 85553
0 5708 7 1 2 85511 85559
0 5709 5 1 1 5708
0 5710 7 1 2 5703 5709
0 5711 5 1 1 5710
0 5712 7 1 2 82465 5711
0 5713 5 1 1 5712
0 5714 7 3 2 1670 2779
0 5715 5 1 1 85577
0 5716 7 8 2 73246 85578
0 5717 5 6 1 85580
0 5718 7 1 2 67375 85581
0 5719 5 1 1 5718
0 5720 7 1 2 1865 5719
0 5721 5 2 1 5720
0 5722 7 1 2 85505 84342
0 5723 7 1 2 85594 5722
0 5724 5 1 1 5723
0 5725 7 1 2 5713 5724
0 5726 5 1 1 5725
0 5727 7 1 2 66866 5726
0 5728 5 1 1 5727
0 5729 7 3 2 66636 75025
0 5730 7 1 2 65329 79618
0 5731 7 1 2 85596 5730
0 5732 5 1 1 5731
0 5733 7 1 2 5728 5732
0 5734 7 1 2 5695 5733
0 5735 5 1 1 5734
0 5736 7 1 2 68314 5735
0 5737 5 1 1 5736
0 5738 7 3 2 76747 85080
0 5739 5 4 1 85599
0 5740 7 2 2 78439 85600
0 5741 5 1 1 85606
0 5742 7 2 2 72016 5741
0 5743 5 1 1 85608
0 5744 7 1 2 82962 85609
0 5745 5 1 1 5744
0 5746 7 1 2 74773 83266
0 5747 7 1 2 85486 5746
0 5748 5 1 1 5747
0 5749 7 1 2 5745 5748
0 5750 5 1 1 5749
0 5751 7 1 2 66867 5750
0 5752 5 1 1 5751
0 5753 7 2 2 67376 72017
0 5754 5 4 1 85610
0 5755 7 2 2 71520 85611
0 5756 5 2 1 85616
0 5757 7 1 2 77058 74426
0 5758 7 1 2 85617 5757
0 5759 5 1 1 5758
0 5760 7 1 2 5752 5759
0 5761 5 1 1 5760
0 5762 7 1 2 65330 5761
0 5763 5 1 1 5762
0 5764 7 2 2 66868 77545
0 5765 5 2 1 85620
0 5766 7 2 2 77567 76362
0 5767 5 2 1 85624
0 5768 7 1 2 85622 85626
0 5769 5 1 1 5768
0 5770 7 5 2 67611 72018
0 5771 5 2 1 85628
0 5772 7 1 2 79303 85629
0 5773 7 1 2 5769 5772
0 5774 5 1 1 5773
0 5775 7 1 2 5763 5774
0 5776 5 1 1 5775
0 5777 7 1 2 66637 5776
0 5778 5 1 1 5777
0 5779 7 1 2 5737 5778
0 5780 7 1 2 5608 5779
0 5781 5 1 1 5780
0 5782 7 13 2 66373 68090
0 5783 7 3 2 84066 85635
0 5784 7 1 2 5781 85648
0 5785 5 1 1 5784
0 5786 7 1 2 69710 5785
0 5787 7 1 2 5556 5786
0 5788 5 1 1 5787
0 5789 7 1 2 69498 5788
0 5790 7 1 2 5319 5789
0 5791 5 1 1 5790
0 5792 7 7 2 69304 65331
0 5793 7 4 2 79744 85651
0 5794 7 1 2 73906 85658
0 5795 5 1 1 5794
0 5796 7 5 2 63903 79337
0 5797 7 3 2 69945 74258
0 5798 7 1 2 75846 85667
0 5799 7 1 2 85662 5798
0 5800 5 1 1 5799
0 5801 7 1 2 5795 5800
0 5802 5 1 1 5801
0 5803 7 1 2 62321 5802
0 5804 5 1 1 5803
0 5805 7 2 2 76207 75317
0 5806 5 2 1 85670
0 5807 7 1 2 85659 85671
0 5808 5 1 1 5807
0 5809 7 1 2 5804 5808
0 5810 5 1 1 5809
0 5811 7 1 2 73932 5810
0 5812 5 1 1 5811
0 5813 7 3 2 70241 78440
0 5814 5 1 1 85674
0 5815 7 1 2 71199 5814
0 5816 5 2 1 5815
0 5817 7 1 2 74575 78426
0 5818 5 1 1 5817
0 5819 7 1 2 85677 5818
0 5820 5 1 1 5819
0 5821 7 1 2 68315 5820
0 5822 5 1 1 5821
0 5823 7 1 2 63481 75974
0 5824 5 8 1 5823
0 5825 7 2 2 68316 74576
0 5826 5 4 1 85687
0 5827 7 2 2 62322 85689
0 5828 5 2 1 85693
0 5829 7 5 2 85679 85695
0 5830 7 1 2 85602 85697
0 5831 5 1 1 5830
0 5832 7 14 2 67377 68559
0 5833 5 1 1 85702
0 5834 7 2 2 85703 72367
0 5835 5 2 1 85716
0 5836 7 1 2 68317 78427
0 5837 5 1 1 5836
0 5838 7 1 2 85718 5837
0 5839 5 1 1 5838
0 5840 7 1 2 67155 5839
0 5841 5 1 1 5840
0 5842 7 1 2 5831 5841
0 5843 7 1 2 5822 5842
0 5844 5 1 1 5843
0 5845 7 11 2 66869 69305
0 5846 7 1 2 85720 83576
0 5847 7 1 2 5844 5846
0 5848 5 1 1 5847
0 5849 7 1 2 5812 5848
0 5850 5 1 1 5849
0 5851 7 1 2 70859 5850
0 5852 5 1 1 5851
0 5853 7 1 2 82206 85660
0 5854 7 1 2 84951 5853
0 5855 5 1 1 5854
0 5856 7 1 2 5852 5855
0 5857 5 1 1 5856
0 5858 7 1 2 64066 5857
0 5859 5 1 1 5858
0 5860 7 3 2 63904 75537
0 5861 5 6 1 85731
0 5862 7 1 2 68560 85734
0 5863 5 1 1 5862
0 5864 7 1 2 62508 5863
0 5865 5 1 1 5864
0 5866 7 4 2 68776 65935
0 5867 5 1 1 85740
0 5868 7 5 2 67612 85741
0 5869 5 2 1 85744
0 5870 7 1 2 63711 85749
0 5871 5 4 1 5870
0 5872 7 1 2 68318 85751
0 5873 7 1 2 5865 5872
0 5874 5 1 1 5873
0 5875 7 1 2 85742 84876
0 5876 5 1 1 5875
0 5877 7 1 2 63482 5876
0 5878 5 1 1 5877
0 5879 7 5 2 62509 75538
0 5880 5 8 1 85755
0 5881 7 1 2 63905 85756
0 5882 5 4 1 5881
0 5883 7 1 2 77556 85768
0 5884 7 1 2 5878 5883
0 5885 5 1 1 5884
0 5886 7 1 2 5874 5885
0 5887 5 1 1 5886
0 5888 7 1 2 77125 5887
0 5889 5 1 1 5888
0 5890 7 5 2 62323 75069
0 5891 5 1 1 85772
0 5892 7 2 2 65062 75659
0 5893 5 1 1 85777
0 5894 7 1 2 85773 85778
0 5895 5 1 1 5894
0 5896 7 1 2 62510 82531
0 5897 5 2 1 5896
0 5898 7 1 2 70610 85779
0 5899 7 1 2 85752 5898
0 5900 5 1 1 5899
0 5901 7 1 2 689 5900
0 5902 5 1 1 5901
0 5903 7 1 2 69946 5902
0 5904 5 1 1 5903
0 5905 7 3 2 65675 74880
0 5906 5 2 1 85781
0 5907 7 1 2 62755 85782
0 5908 5 1 1 5907
0 5909 7 1 2 5904 5908
0 5910 5 1 1 5909
0 5911 7 1 2 67156 5910
0 5912 5 1 1 5911
0 5913 7 1 2 5895 5912
0 5914 5 1 1 5913
0 5915 7 1 2 65332 5914
0 5916 5 1 1 5915
0 5917 7 1 2 5889 5916
0 5918 5 1 1 5917
0 5919 7 1 2 68932 5918
0 5920 5 1 1 5919
0 5921 7 1 2 79662 84813
0 5922 5 1 1 5921
0 5923 7 2 2 70611 83205
0 5924 7 4 2 68319 73386
0 5925 5 2 1 85788
0 5926 7 1 2 85786 85789
0 5927 5 1 1 5926
0 5928 7 1 2 74649 76864
0 5929 5 1 1 5928
0 5930 7 1 2 5927 5929
0 5931 5 1 1 5930
0 5932 7 1 2 71896 5931
0 5933 5 1 1 5932
0 5934 7 1 2 5922 5933
0 5935 7 1 2 5920 5934
0 5936 5 1 1 5935
0 5937 7 1 2 66870 5936
0 5938 5 1 1 5937
0 5939 7 3 2 68777 71647
0 5940 7 1 2 74396 85794
0 5941 5 1 1 5940
0 5942 7 1 2 75118 5941
0 5943 5 1 1 5942
0 5944 7 1 2 71897 5943
0 5945 5 1 1 5944
0 5946 7 3 2 68561 71648
0 5947 7 1 2 82190 85797
0 5948 5 1 1 5947
0 5949 7 1 2 5945 5948
0 5950 5 1 1 5949
0 5951 7 1 2 65063 5950
0 5952 5 1 1 5951
0 5953 7 5 2 68320 75026
0 5954 7 1 2 85800 85798
0 5955 5 1 1 5954
0 5956 7 1 2 5952 5955
0 5957 5 1 1 5956
0 5958 7 1 2 65333 5957
0 5959 5 1 1 5958
0 5960 7 2 2 74881 77568
0 5961 7 1 2 80810 85805
0 5962 5 1 1 5961
0 5963 7 1 2 5959 5962
0 5964 5 1 1 5963
0 5965 7 1 2 62756 5964
0 5966 5 1 1 5965
0 5967 7 2 2 78374 83463
0 5968 7 1 2 80866 85027
0 5969 7 1 2 85807 5968
0 5970 5 1 1 5969
0 5971 7 1 2 5966 5970
0 5972 7 1 2 5938 5971
0 5973 5 1 1 5972
0 5974 7 1 2 79420 5973
0 5975 5 1 1 5974
0 5976 7 1 2 5859 5975
0 5977 5 1 1 5976
0 5978 7 1 2 64868 5977
0 5979 5 1 1 5978
0 5980 7 9 2 67378 74674
0 5981 5 4 1 85809
0 5982 7 9 2 62757 69947
0 5983 5 1 1 85822
0 5984 7 3 2 72019 85823
0 5985 7 1 2 85810 85831
0 5986 5 1 1 5985
0 5987 7 16 2 65936 74065
0 5988 5 2 1 85834
0 5989 7 2 2 62002 77068
0 5990 5 1 1 85852
0 5991 7 1 2 5294 5990
0 5992 5 2 1 5991
0 5993 7 1 2 85835 85854
0 5994 5 1 1 5993
0 5995 7 1 2 5986 5994
0 5996 5 1 1 5995
0 5997 7 1 2 70612 5996
0 5998 5 1 1 5997
0 5999 7 5 2 62758 71898
0 6000 5 1 1 85856
0 6001 7 1 2 85857 77371
0 6002 5 1 1 6001
0 6003 7 1 2 5998 6002
0 6004 5 1 1 6003
0 6005 7 3 2 65334 82772
0 6006 7 1 2 83644 85861
0 6007 7 1 2 6004 6006
0 6008 5 1 1 6007
0 6009 7 1 2 5979 6008
0 6010 5 1 1 6009
0 6011 7 1 2 66638 6010
0 6012 5 1 1 6011
0 6013 7 4 2 72020 73822
0 6014 5 1 1 85864
0 6015 7 5 2 67379 83756
0 6016 7 1 2 85865 85868
0 6017 5 1 1 6016
0 6018 7 9 2 68933 78034
0 6019 7 1 2 74427 85873
0 6020 5 1 1 6019
0 6021 7 1 2 6017 6020
0 6022 5 1 1 6021
0 6023 7 1 2 83898 6022
0 6024 5 1 1 6023
0 6025 7 4 2 67380 79338
0 6026 7 1 2 73770 80340
0 6027 7 1 2 80769 76991
0 6028 7 1 2 6026 6027
0 6029 7 1 2 85882 6028
0 6030 5 1 1 6029
0 6031 7 1 2 6024 6030
0 6032 5 1 1 6031
0 6033 7 1 2 66871 6032
0 6034 5 1 1 6033
0 6035 7 14 2 69306 65937
0 6036 7 4 2 65064 78468
0 6037 7 3 2 85886 85900
0 6038 7 3 2 66639 74463
0 6039 7 1 2 73727 85907
0 6040 7 1 2 85904 6039
0 6041 5 1 1 6040
0 6042 7 1 2 6034 6041
0 6043 5 1 1 6042
0 6044 7 1 2 71899 6043
0 6045 5 1 1 6044
0 6046 7 11 2 61749 67381
0 6047 7 2 2 85910 71012
0 6048 7 5 2 69499 82390
0 6049 7 1 2 84509 85923
0 6050 7 1 2 85921 6049
0 6051 5 1 1 6050
0 6052 7 4 2 67157 65676
0 6053 5 2 1 85928
0 6054 7 1 2 72517 73939
0 6055 7 1 2 85932 6054
0 6056 7 1 2 83714 6055
0 6057 7 1 2 84238 6056
0 6058 5 1 1 6057
0 6059 7 1 2 6051 6058
0 6060 5 1 1 6059
0 6061 7 1 2 76620 6060
0 6062 5 1 1 6061
0 6063 7 1 2 65065 6062
0 6064 5 1 1 6063
0 6065 7 1 2 71804 75467
0 6066 5 3 1 6065
0 6067 7 7 2 68562 72518
0 6068 7 1 2 61750 85937
0 6069 5 1 1 6068
0 6070 7 1 2 85934 6069
0 6071 5 1 1 6070
0 6072 7 1 2 64869 78441
0 6073 7 1 2 6071 6072
0 6074 5 1 1 6073
0 6075 7 3 2 67613 85403
0 6076 5 4 1 85944
0 6077 7 1 2 62759 71649
0 6078 5 4 1 6077
0 6079 7 1 2 85947 85951
0 6080 5 2 1 6079
0 6081 7 1 2 66640 83471
0 6082 7 1 2 85955 6081
0 6083 5 1 1 6082
0 6084 7 1 2 6074 6083
0 6085 5 1 1 6084
0 6086 7 1 2 73286 6085
0 6087 5 1 1 6086
0 6088 7 9 2 65938 71900
0 6089 7 1 2 85957 75587
0 6090 5 1 1 6089
0 6091 7 8 2 63712 79894
0 6092 5 2 1 85966
0 6093 7 3 2 65677 71418
0 6094 5 1 1 85976
0 6095 7 1 2 62760 85977
0 6096 7 1 2 85967 6095
0 6097 5 1 1 6096
0 6098 7 1 2 6090 6097
0 6099 5 1 1 6098
0 6100 7 1 2 68934 6099
0 6101 5 1 1 6100
0 6102 7 2 2 80467 75681
0 6103 7 1 2 85979 82391
0 6104 7 1 2 79895 6103
0 6105 5 1 1 6104
0 6106 7 1 2 6101 6105
0 6107 7 1 2 6087 6106
0 6108 5 1 1 6107
0 6109 7 1 2 69500 6108
0 6110 5 1 1 6109
0 6111 7 2 2 73287 84955
0 6112 7 4 2 81979 81123
0 6113 5 1 1 85983
0 6114 7 1 2 85981 85984
0 6115 5 1 1 6114
0 6116 7 3 2 78802 75672
0 6117 7 1 2 85987 79845
0 6118 5 1 1 6117
0 6119 7 1 2 79066 85938
0 6120 5 1 1 6119
0 6121 7 1 2 6118 6120
0 6122 5 1 1 6121
0 6123 7 1 2 61751 6122
0 6124 5 1 1 6123
0 6125 7 1 2 77482 79846
0 6126 5 1 1 6125
0 6127 7 1 2 83472 84648
0 6128 5 1 1 6127
0 6129 7 1 2 6126 6128
0 6130 5 1 1 6129
0 6131 7 1 2 78257 6130
0 6132 5 1 1 6131
0 6133 7 1 2 6124 6132
0 6134 5 1 1 6133
0 6135 7 1 2 62324 6134
0 6136 5 1 1 6135
0 6137 7 3 2 69501 71200
0 6138 7 2 2 71901 84299
0 6139 5 2 1 85993
0 6140 7 2 2 63713 84649
0 6141 5 1 1 85997
0 6142 7 1 2 85995 6141
0 6143 5 1 1 6142
0 6144 7 1 2 71419 6143
0 6145 5 1 1 6144
0 6146 7 1 2 63714 84102
0 6147 5 1 1 6146
0 6148 7 1 2 6145 6147
0 6149 5 1 1 6148
0 6150 7 1 2 85990 6149
0 6151 5 1 1 6150
0 6152 7 1 2 6136 6151
0 6153 5 1 1 6152
0 6154 7 1 2 70613 6153
0 6155 5 1 1 6154
0 6156 7 1 2 6115 6155
0 6157 7 1 2 6110 6156
0 6158 5 1 1 6157
0 6159 7 1 2 63483 6158
0 6160 5 1 1 6159
0 6161 7 10 2 62761 68563
0 6162 7 1 2 62511 75284
0 6163 7 3 2 85999 6162
0 6164 5 2 1 86009
0 6165 7 1 2 75468 85924
0 6166 7 1 2 86010 6165
0 6167 5 1 1 6166
0 6168 7 1 2 6160 6167
0 6169 5 1 1 6168
0 6170 7 1 2 64456 6169
0 6171 5 1 1 6170
0 6172 7 1 2 74856 84746
0 6173 5 1 1 6172
0 6174 7 9 2 72100 71902
0 6175 7 1 2 68321 86014
0 6176 5 1 1 6175
0 6177 7 1 2 6173 6176
0 6178 5 1 1 6177
0 6179 7 3 2 79421 82164
0 6180 7 1 2 82612 86023
0 6181 7 1 2 6178 6180
0 6182 5 1 1 6181
0 6183 7 1 2 69948 6182
0 6184 7 1 2 6171 6183
0 6185 5 1 1 6184
0 6186 7 1 2 6064 6185
0 6187 5 1 1 6186
0 6188 7 1 2 6045 6187
0 6189 5 1 1 6188
0 6190 7 1 2 70242 6189
0 6191 5 1 1 6190
0 6192 7 12 2 61752 64457
0 6193 7 10 2 63484 64067
0 6194 7 1 2 67614 86038
0 6195 7 1 2 85069 6194
0 6196 5 1 1 6195
0 6197 7 22 2 62003 65335
0 6198 5 1 1 86048
0 6199 7 1 2 68935 86049
0 6200 7 1 2 79930 6199
0 6201 5 1 1 6200
0 6202 7 1 2 6196 6201
0 6203 5 1 1 6202
0 6204 7 1 2 68564 6203
0 6205 5 1 1 6204
0 6206 7 3 2 68936 73057
0 6207 7 1 2 76378 86070
0 6208 5 1 1 6207
0 6209 7 1 2 6205 6208
0 6210 5 1 1 6209
0 6211 7 1 2 67158 6210
0 6212 5 1 1 6211
0 6213 7 3 2 70614 76455
0 6214 7 1 2 76242 84972
0 6215 7 1 2 86073 6214
0 6216 5 1 1 6215
0 6217 7 1 2 6212 6216
0 6218 5 1 1 6217
0 6219 7 1 2 65939 6218
0 6220 5 1 1 6219
0 6221 7 1 2 79218 74023
0 6222 7 1 2 84029 6221
0 6223 5 1 1 6222
0 6224 7 1 2 6220 6223
0 6225 5 1 1 6224
0 6226 7 1 2 78586 6225
0 6227 5 1 1 6226
0 6228 7 2 2 72021 79219
0 6229 5 2 1 86076
0 6230 7 1 2 1115 86078
0 6231 5 1 1 6230
0 6232 7 7 2 65336 78534
0 6233 7 3 2 70615 74259
0 6234 7 1 2 86080 86087
0 6235 7 1 2 6231 6234
0 6236 5 1 1 6235
0 6237 7 1 2 6227 6236
0 6238 5 1 1 6237
0 6239 7 1 2 69502 6238
0 6240 5 1 1 6239
0 6241 7 1 2 74172 81888
0 6242 7 1 2 83516 6241
0 6243 7 1 2 84834 80527
0 6244 7 1 2 6242 6243
0 6245 5 1 1 6244
0 6246 7 1 2 6240 6245
0 6247 5 1 1 6246
0 6248 7 1 2 86026 6247
0 6249 5 1 1 6248
0 6250 7 1 2 6191 6249
0 6251 7 1 2 6012 6250
0 6252 5 1 1 6251
0 6253 7 1 2 63253 6252
0 6254 5 1 1 6253
0 6255 7 9 2 69949 82773
0 6256 7 2 2 82678 86090
0 6257 5 3 1 86099
0 6258 7 1 2 83639 86101
0 6259 5 1 1 6258
0 6260 7 5 2 62325 75179
0 6261 5 1 1 86104
0 6262 7 2 2 65337 72262
0 6263 7 1 2 86105 86109
0 6264 5 1 1 6263
0 6265 7 1 2 71659 85213
0 6266 7 1 2 83878 6265
0 6267 5 1 1 6266
0 6268 7 1 2 6264 6267
0 6269 5 1 1 6268
0 6270 7 2 2 67615 83078
0 6271 7 1 2 6269 86111
0 6272 5 1 1 6271
0 6273 7 3 2 70860 73058
0 6274 7 1 2 83029 75318
0 6275 7 1 2 79568 6274
0 6276 7 1 2 86113 6275
0 6277 5 1 1 6276
0 6278 7 1 2 6272 6277
0 6279 5 1 1 6278
0 6280 7 1 2 6259 6279
0 6281 5 1 1 6280
0 6282 7 1 2 74723 74738
0 6283 5 1 1 6282
0 6284 7 1 2 76439 6283
0 6285 5 1 1 6284
0 6286 7 4 2 67159 84333
0 6287 5 2 1 86116
0 6288 7 4 2 72263 76243
0 6289 5 3 1 86122
0 6290 7 1 2 86117 86123
0 6291 5 1 1 6290
0 6292 7 1 2 6285 6291
0 6293 5 1 1 6292
0 6294 7 1 2 79636 6293
0 6295 5 1 1 6294
0 6296 7 17 2 69711 79339
0 6297 7 1 2 86129 85167
0 6298 5 1 1 6297
0 6299 7 1 2 6295 6298
0 6300 5 1 1 6299
0 6301 7 1 2 61753 6300
0 6302 5 1 1 6301
0 6303 7 3 2 76456 73288
0 6304 7 1 2 74961 86146
0 6305 5 1 1 6304
0 6306 7 4 2 71903 78305
0 6307 7 1 2 75049 86149
0 6308 5 1 1 6307
0 6309 7 1 2 6305 6308
0 6310 5 1 1 6309
0 6311 7 1 2 85262 79422
0 6312 7 1 2 6310 6311
0 6313 5 1 1 6312
0 6314 7 1 2 6302 6313
0 6315 5 1 1 6314
0 6316 7 1 2 62004 6315
0 6317 5 1 1 6316
0 6318 7 3 2 65338 71150
0 6319 7 8 2 68565 64870
0 6320 7 3 2 82048 86156
0 6321 7 1 2 86153 86164
0 6322 5 1 1 6321
0 6323 7 1 2 71420 85630
0 6324 5 1 1 6323
0 6325 7 1 2 77783 6324
0 6326 5 1 1 6325
0 6327 7 12 2 71201 71904
0 6328 5 1 1 86167
0 6329 7 2 2 70243 74833
0 6330 5 1 1 86179
0 6331 7 1 2 86168 6330
0 6332 7 1 2 6326 6331
0 6333 5 1 1 6332
0 6334 7 1 2 6322 6333
0 6335 5 1 1 6334
0 6336 7 1 2 65678 6335
0 6337 5 1 1 6336
0 6338 7 4 2 68566 77569
0 6339 7 1 2 72316 77893
0 6340 7 1 2 86181 6339
0 6341 5 1 1 6340
0 6342 7 1 2 6337 6341
0 6343 5 1 1 6342
0 6344 7 1 2 63485 6343
0 6345 5 1 1 6344
0 6346 7 9 2 68322 75937
0 6347 5 1 1 86185
0 6348 7 7 2 62762 74173
0 6349 5 2 1 86194
0 6350 7 1 2 76757 78813
0 6351 7 1 2 86195 6350
0 6352 7 1 2 86186 6351
0 6353 5 1 1 6352
0 6354 7 1 2 6345 6353
0 6355 5 1 1 6354
0 6356 7 1 2 64651 6355
0 6357 5 1 1 6356
0 6358 7 3 2 61754 83493
0 6359 7 1 2 86203 75619
0 6360 5 1 1 6359
0 6361 7 7 2 71650 75521
0 6362 5 2 1 86206
0 6363 7 1 2 5385 86213
0 6364 5 4 1 6363
0 6365 7 1 2 67382 86215
0 6366 5 1 1 6365
0 6367 7 2 2 71651 85745
0 6368 5 1 1 86219
0 6369 7 1 2 6366 6368
0 6370 5 2 1 6369
0 6371 7 1 2 68323 79165
0 6372 7 1 2 86221 6371
0 6373 5 1 1 6372
0 6374 7 1 2 6360 6373
0 6375 5 1 1 6374
0 6376 7 1 2 71905 6375
0 6377 5 1 1 6376
0 6378 7 2 2 79166 82509
0 6379 7 1 2 85850 79996
0 6380 5 1 1 6379
0 6381 7 1 2 86223 6380
0 6382 5 1 1 6381
0 6383 7 1 2 84309 86224
0 6384 5 1 1 6383
0 6385 7 2 2 61755 77792
0 6386 7 1 2 78469 75180
0 6387 7 1 2 86225 6386
0 6388 5 1 1 6387
0 6389 7 1 2 6384 6388
0 6390 5 1 1 6389
0 6391 7 1 2 75660 6390
0 6392 5 1 1 6391
0 6393 7 1 2 6382 6392
0 6394 7 1 2 6377 6393
0 6395 5 1 1 6394
0 6396 7 1 2 65339 6395
0 6397 5 1 1 6396
0 6398 7 5 2 70244 79117
0 6399 7 1 2 72101 82949
0 6400 7 1 2 86227 6399
0 6401 5 1 1 6400
0 6402 7 1 2 63906 650
0 6403 5 2 1 6402
0 6404 7 7 2 83369 86232
0 6405 7 1 2 67616 86234
0 6406 5 1 1 6405
0 6407 7 4 2 71202 72102
0 6408 5 1 1 86241
0 6409 7 1 2 6406 6408
0 6410 5 1 1 6409
0 6411 7 1 2 79167 73907
0 6412 7 1 2 6410 6411
0 6413 5 1 1 6412
0 6414 7 1 2 6401 6413
0 6415 5 1 1 6414
0 6416 7 1 2 65679 6415
0 6417 5 1 1 6416
0 6418 7 2 2 63486 80291
0 6419 5 1 1 86245
0 6420 7 3 2 68324 71203
0 6421 5 4 1 86247
0 6422 7 1 2 83473 86248
0 6423 5 1 1 6422
0 6424 7 1 2 6419 6423
0 6425 5 1 1 6424
0 6426 7 1 2 83327 84650
0 6427 7 1 2 6425 6426
0 6428 5 1 1 6427
0 6429 7 1 2 6417 6428
0 6430 5 1 1 6429
0 6431 7 1 2 67160 6430
0 6432 5 1 1 6431
0 6433 7 1 2 71039 84651
0 6434 5 2 1 6433
0 6435 7 1 2 71421 78306
0 6436 5 1 1 6435
0 6437 7 1 2 86254 6436
0 6438 5 1 1 6437
0 6439 7 7 2 68567 64652
0 6440 7 1 2 86256 74701
0 6441 7 1 2 6438 6440
0 6442 5 1 1 6441
0 6443 7 1 2 6432 6442
0 6444 7 1 2 6397 6443
0 6445 5 1 1 6444
0 6446 7 1 2 66872 6445
0 6447 5 1 1 6446
0 6448 7 1 2 6357 6447
0 6449 5 1 1 6448
0 6450 7 1 2 69307 6449
0 6451 5 1 1 6450
0 6452 7 1 2 6317 6451
0 6453 5 1 1 6452
0 6454 7 1 2 65066 6453
0 6455 5 1 1 6454
0 6456 7 1 2 83935 85855
0 6457 5 1 1 6456
0 6458 7 2 2 78535 79423
0 6459 7 1 2 86263 80615
0 6460 5 1 1 6459
0 6461 7 1 2 6457 6460
0 6462 5 1 1 6461
0 6463 7 1 2 75522 6462
0 6464 5 1 1 6463
0 6465 7 1 2 86000 79952
0 6466 7 1 2 86024 6465
0 6467 5 1 1 6466
0 6468 7 1 2 6464 6467
0 6469 5 1 1 6468
0 6470 7 1 2 68937 6469
0 6471 5 1 1 6470
0 6472 7 7 2 62005 71906
0 6473 5 3 1 86265
0 6474 7 1 2 85811 75641
0 6475 5 1 1 6474
0 6476 7 1 2 86272 6475
0 6477 5 1 1 6476
0 6478 7 1 2 86130 85824
0 6479 7 1 2 6477 6478
0 6480 5 1 1 6479
0 6481 7 1 2 6471 6480
0 6482 5 1 1 6481
0 6483 7 1 2 65340 6482
0 6484 5 1 1 6483
0 6485 7 2 2 75181 85362
0 6486 5 1 1 86275
0 6487 7 5 2 69950 72444
0 6488 7 1 2 86131 86277
0 6489 7 1 2 86276 6488
0 6490 5 1 1 6489
0 6491 7 1 2 6484 6490
0 6492 5 1 1 6491
0 6493 7 1 2 61756 6492
0 6494 5 1 1 6493
0 6495 7 1 2 75341 72519
0 6496 5 1 1 6495
0 6497 7 1 2 85618 6496
0 6498 5 1 1 6497
0 6499 7 1 2 75217 6498
0 6500 5 1 1 6499
0 6501 7 1 2 62006 86150
0 6502 5 1 1 6501
0 6503 7 1 2 6500 6502
0 6504 5 1 1 6503
0 6505 7 6 2 64653 79795
0 6506 7 5 2 70245 78536
0 6507 7 1 2 86282 86288
0 6508 7 1 2 6504 6507
0 6509 5 1 1 6508
0 6510 7 1 2 6494 6509
0 6511 5 1 1 6510
0 6512 7 1 2 63487 6511
0 6513 5 1 1 6512
0 6514 7 1 2 75285 72383
0 6515 5 2 1 6514
0 6516 7 1 2 78172 86293
0 6517 5 1 1 6516
0 6518 7 1 2 86100 6517
0 6519 5 1 1 6518
0 6520 7 3 2 70616 79424
0 6521 7 1 2 81202 77483
0 6522 7 1 2 86295 6521
0 6523 5 1 1 6522
0 6524 7 1 2 6519 6523
0 6525 5 1 1 6524
0 6526 7 1 2 68568 6525
0 6527 5 1 1 6526
0 6528 7 19 2 64068 69308
0 6529 7 3 2 86298 78470
0 6530 7 1 2 83757 84961
0 6531 7 1 2 77583 6530
0 6532 7 1 2 86317 6531
0 6533 5 1 1 6532
0 6534 7 1 2 6527 6533
0 6535 5 1 1 6534
0 6536 7 1 2 70246 6535
0 6537 5 1 1 6536
0 6538 7 2 2 68325 77896
0 6539 7 1 2 79425 75027
0 6540 7 1 2 84263 6539
0 6541 7 1 2 86320 6540
0 6542 5 1 1 6541
0 6543 7 1 2 6537 6542
0 6544 5 1 1 6543
0 6545 7 1 2 76992 6544
0 6546 5 1 1 6545
0 6547 7 1 2 6513 6546
0 6548 7 1 2 6455 6547
0 6549 5 1 1 6548
0 6550 7 1 2 68091 6549
0 6551 5 1 1 6550
0 6552 7 1 2 6281 6551
0 6553 7 1 2 6254 6552
0 6554 5 1 1 6553
0 6555 7 1 2 76117 6554
0 6556 5 1 1 6555
0 6557 7 2 2 78587 73289
0 6558 5 1 1 86322
0 6559 7 3 2 62007 78537
0 6560 5 3 1 86324
0 6561 7 1 2 84598 86325
0 6562 5 1 1 6561
0 6563 7 1 2 6558 6562
0 6564 5 1 1 6563
0 6565 7 1 2 79392 6564
0 6566 5 1 1 6565
0 6567 7 7 2 69712 76931
0 6568 7 1 2 62008 86330
0 6569 5 1 1 6568
0 6570 7 1 2 6566 6569
0 6571 5 1 1 6570
0 6572 7 2 2 63488 82350
0 6573 7 3 2 85119 86337
0 6574 7 1 2 6571 86339
0 6575 5 1 1 6574
0 6576 7 2 2 75975 3030
0 6577 5 11 1 86342
0 6578 7 1 2 86344 86222
0 6579 5 1 1 6578
0 6580 7 4 2 65341 74774
0 6581 7 2 2 62512 85851
0 6582 5 1 1 86359
0 6583 7 1 2 73191 86360
0 6584 5 1 1 6583
0 6585 7 1 2 74997 6584
0 6586 5 1 1 6585
0 6587 7 1 2 79997 6586
0 6588 5 1 1 6587
0 6589 7 1 2 86355 6588
0 6590 5 1 1 6589
0 6591 7 1 2 6579 6590
0 6592 5 2 1 6591
0 6593 7 1 2 65067 82596
0 6594 7 1 2 84250 6593
0 6595 7 1 2 86361 6594
0 6596 5 1 1 6595
0 6597 7 1 2 6575 6596
0 6598 5 1 1 6597
0 6599 7 1 2 66641 6598
0 6600 5 1 1 6599
0 6601 7 2 2 77508 75065
0 6602 7 1 2 62513 86363
0 6603 5 1 1 6602
0 6604 7 3 2 66873 71002
0 6605 7 5 2 65940 85070
0 6606 7 2 2 86365 86368
0 6607 5 1 1 86373
0 6608 7 1 2 70247 86374
0 6609 5 1 1 6608
0 6610 7 1 2 6603 6609
0 6611 5 1 1 6610
0 6612 7 1 2 62326 6611
0 6613 5 1 1 6612
0 6614 7 11 2 67383 70248
0 6615 7 1 2 77388 86375
0 6616 7 1 2 84880 6615
0 6617 5 1 1 6616
0 6618 7 1 2 6613 6617
0 6619 5 1 1 6618
0 6620 7 1 2 65068 6619
0 6621 5 1 1 6620
0 6622 7 2 2 62009 80535
0 6623 5 1 1 86386
0 6624 7 1 2 76333 77402
0 6625 7 7 2 62327 65342
0 6626 5 3 1 86388
0 6627 7 1 2 86389 73940
0 6628 7 1 2 6624 6627
0 6629 7 1 2 86387 6628
0 6630 5 1 1 6629
0 6631 7 1 2 6621 6630
0 6632 5 1 1 6631
0 6633 7 1 2 63715 6632
0 6634 5 1 1 6633
0 6635 7 1 2 77589 85444
0 6636 5 1 1 6635
0 6637 7 1 2 63489 86343
0 6638 5 1 1 6637
0 6639 7 13 2 68778 72520
0 6640 5 2 1 86398
0 6641 7 4 2 67384 69713
0 6642 7 1 2 77658 86413
0 6643 7 1 2 86399 6642
0 6644 7 1 2 6638 6643
0 6645 5 1 1 6644
0 6646 7 1 2 6636 6645
0 6647 5 1 1 6646
0 6648 7 1 2 70617 6647
0 6649 5 1 1 6648
0 6650 7 4 2 70249 85071
0 6651 7 1 2 74857 86417
0 6652 5 1 1 6651
0 6653 7 1 2 75938 82191
0 6654 5 4 1 6653
0 6655 7 1 2 6652 86421
0 6656 5 1 1 6655
0 6657 7 5 2 68938 83206
0 6658 7 1 2 77389 86425
0 6659 7 1 2 6656 6658
0 6660 5 1 1 6659
0 6661 7 1 2 6649 6660
0 6662 7 1 2 6634 6661
0 6663 5 1 1 6662
0 6664 7 1 2 63254 6663
0 6665 5 1 1 6664
0 6666 7 9 2 62763 70250
0 6667 5 2 1 86430
0 6668 7 1 2 86431 79619
0 6669 5 2 1 6668
0 6670 7 1 2 552 86441
0 6671 5 1 1 6670
0 6672 7 1 2 71805 6671
0 6673 5 1 1 6672
0 6674 7 7 2 84599 77557
0 6675 7 1 2 78231 86443
0 6676 5 1 1 6675
0 6677 7 1 2 81229 6676
0 6678 5 1 1 6677
0 6679 7 1 2 74979 6678
0 6680 5 1 1 6679
0 6681 7 1 2 6673 6680
0 6682 5 1 1 6681
0 6683 7 8 2 68092 70618
0 6684 7 1 2 81898 86450
0 6685 7 1 2 6682 6684
0 6686 5 1 1 6685
0 6687 7 1 2 6665 6686
0 6688 5 1 1 6687
0 6689 7 1 2 86027 6688
0 6690 5 1 1 6689
0 6691 7 1 2 6600 6690
0 6692 5 1 1 6691
0 6693 7 1 2 61454 6692
0 6694 5 1 1 6693
0 6695 7 5 2 69309 85636
0 6696 7 3 2 68779 73059
0 6697 5 1 1 86463
0 6698 7 2 2 73096 72489
0 6699 5 5 1 86466
0 6700 7 1 2 67385 86468
0 6701 5 3 1 6700
0 6702 7 1 2 6697 86473
0 6703 5 1 1 6702
0 6704 7 1 2 82963 6703
0 6705 5 1 1 6704
0 6706 7 6 2 69951 76689
0 6707 7 1 2 82207 86476
0 6708 5 1 1 6707
0 6709 7 1 2 6705 6708
0 6710 5 1 1 6709
0 6711 7 1 2 72103 6710
0 6712 5 1 1 6711
0 6713 7 2 2 74539 72264
0 6714 7 1 2 68939 86482
0 6715 5 1 1 6714
0 6716 7 8 2 64069 84004
0 6717 5 5 1 86484
0 6718 7 1 2 63716 75661
0 6719 7 1 2 86485 6718
0 6720 5 1 1 6719
0 6721 7 1 2 6715 6720
0 6722 5 1 1 6721
0 6723 7 1 2 67617 6722
0 6724 5 1 1 6723
0 6725 7 5 2 65343 73247
0 6726 5 9 1 86497
0 6727 7 2 2 77981 86498
0 6728 5 2 1 86511
0 6729 7 2 2 72022 86512
0 6730 5 1 1 86515
0 6731 7 1 2 63717 86516
0 6732 5 1 1 6731
0 6733 7 1 2 6724 6732
0 6734 5 1 1 6733
0 6735 7 1 2 79589 6734
0 6736 5 1 1 6735
0 6737 7 2 2 75342 74610
0 6738 7 2 2 67618 77897
0 6739 7 1 2 86517 86519
0 6740 5 1 1 6739
0 6741 7 3 2 68780 77467
0 6742 7 1 2 72023 86521
0 6743 5 1 1 6742
0 6744 7 1 2 6740 6743
0 6745 5 1 1 6744
0 6746 7 1 2 84943 6745
0 6747 5 1 1 6746
0 6748 7 1 2 6736 6747
0 6749 7 1 2 6712 6748
0 6750 5 1 1 6749
0 6751 7 1 2 77390 6750
0 6752 5 1 1 6751
0 6753 7 7 2 70251 76457
0 6754 7 1 2 85440 86524
0 6755 5 1 1 6754
0 6756 7 1 2 84600 75642
0 6757 7 1 2 76487 6756
0 6758 5 1 1 6757
0 6759 7 1 2 6755 6758
0 6760 5 1 1 6759
0 6761 7 1 2 76865 6760
0 6762 5 1 1 6761
0 6763 7 3 2 71806 74650
0 6764 5 1 1 86531
0 6765 7 1 2 85808 86532
0 6766 5 1 1 6765
0 6767 7 1 2 6762 6766
0 6768 5 1 1 6767
0 6769 7 1 2 64871 6768
0 6770 5 1 1 6769
0 6771 7 1 2 6752 6770
0 6772 5 1 1 6771
0 6773 7 1 2 66642 6772
0 6774 5 1 1 6773
0 6775 7 3 2 84005 79676
0 6776 5 1 1 86534
0 6777 7 4 2 68326 78538
0 6778 7 1 2 74775 75697
0 6779 7 1 2 86537 6778
0 6780 7 1 2 86535 6779
0 6781 5 1 1 6780
0 6782 7 1 2 6774 6781
0 6783 5 1 1 6782
0 6784 7 1 2 86458 6783
0 6785 5 1 1 6784
0 6786 7 2 2 83030 73737
0 6787 7 2 2 76770 83207
0 6788 7 1 2 86541 86543
0 6789 5 1 1 6788
0 6790 7 1 2 1933 86327
0 6791 5 1 1 6790
0 6792 7 10 2 70252 73290
0 6793 5 5 1 86545
0 6794 7 1 2 86546 83664
0 6795 7 1 2 6791 6794
0 6796 5 1 1 6795
0 6797 7 1 2 6789 6796
0 6798 5 1 1 6797
0 6799 7 1 2 71807 6798
0 6800 5 1 1 6799
0 6801 7 2 2 73602 75319
0 6802 5 2 1 86560
0 6803 7 1 2 74669 86562
0 6804 5 2 1 6803
0 6805 7 1 2 83538 86564
0 6806 5 1 1 6805
0 6807 7 15 2 63255 65344
0 6808 7 4 2 65069 74776
0 6809 7 2 2 86566 86581
0 6810 5 1 1 86585
0 6811 7 1 2 6806 6810
0 6812 5 1 1 6811
0 6813 7 2 2 71687 74149
0 6814 7 1 2 68940 86587
0 6815 7 1 2 6812 6814
0 6816 5 1 1 6815
0 6817 7 1 2 6800 6816
0 6818 5 1 1 6817
0 6819 7 1 2 82836 6818
0 6820 5 1 1 6819
0 6821 7 2 2 66374 71772
0 6822 7 1 2 63907 83554
0 6823 7 1 2 86589 6822
0 6824 7 2 2 64872 76932
0 6825 7 2 2 62514 81578
0 6826 7 1 2 86591 86593
0 6827 7 1 2 6823 6826
0 6828 5 1 1 6827
0 6829 7 1 2 6820 6828
0 6830 5 1 1 6829
0 6831 7 1 2 78442 6830
0 6832 5 1 1 6831
0 6833 7 1 2 6785 6832
0 6834 7 1 2 6694 6833
0 6835 5 1 1 6834
0 6836 7 1 2 63081 6835
0 6837 5 1 1 6836
0 6838 7 1 2 66874 74556
0 6839 5 1 1 6838
0 6840 7 1 2 86345 76379
0 6841 5 1 1 6840
0 6842 7 1 2 6839 6841
0 6843 5 1 1 6842
0 6844 7 1 2 65680 6843
0 6845 5 1 1 6844
0 6846 7 25 2 66875 62328
0 6847 5 4 1 86595
0 6848 7 14 2 63718 86596
0 6849 5 1 1 86624
0 6850 7 1 2 86625 84586
0 6851 5 1 1 6850
0 6852 7 1 2 6845 6851
0 6853 5 1 1 6852
0 6854 7 1 2 67619 6853
0 6855 5 1 1 6854
0 6856 7 3 2 63719 76690
0 6857 7 2 2 73387 86638
0 6858 5 1 1 86641
0 6859 7 1 2 86597 86642
0 6860 5 1 1 6859
0 6861 7 1 2 6855 6860
0 6862 5 1 1 6861
0 6863 7 1 2 64070 6862
0 6864 5 1 1 6863
0 6865 7 16 2 62515 68327
0 6866 7 4 2 63908 86643
0 6867 5 1 1 86659
0 6868 7 1 2 86620 6867
0 6869 5 1 1 6868
0 6870 7 3 2 68569 72445
0 6871 5 1 1 86663
0 6872 7 1 2 71122 86664
0 6873 7 1 2 6869 6872
0 6874 5 1 1 6873
0 6875 7 1 2 6864 6874
0 6876 5 1 1 6875
0 6877 7 1 2 64873 82104
0 6878 7 1 2 6876 6877
0 6879 5 1 1 6878
0 6880 7 1 2 62764 80547
0 6881 5 2 1 6880
0 6882 7 1 2 71754 86666
0 6883 5 1 1 6882
0 6884 7 8 2 61455 62010
0 6885 7 1 2 86668 82230
0 6886 7 1 2 86147 6885
0 6887 7 1 2 6883 6886
0 6888 5 1 1 6887
0 6889 7 1 2 6879 6888
0 6890 5 1 1 6889
0 6891 7 1 2 63082 6890
0 6892 5 1 1 6891
0 6893 7 7 2 71907 75131
0 6894 7 2 2 70861 85652
0 6895 7 2 2 64874 76035
0 6896 7 1 2 86683 86685
0 6897 7 1 2 86676 6896
0 6898 5 1 1 6897
0 6899 7 1 2 6892 6898
0 6900 5 1 1 6899
0 6901 7 1 2 65070 6900
0 6902 5 1 1 6901
0 6903 7 2 2 84053 77143
0 6904 7 1 2 77223 74611
0 6905 7 1 2 79851 75447
0 6906 7 1 2 6904 6905
0 6907 7 1 2 86687 6906
0 6908 5 1 1 6907
0 6909 7 1 2 6902 6908
0 6910 5 1 1 6909
0 6911 7 1 2 83079 6910
0 6912 5 1 1 6911
0 6913 7 2 2 77837 72299
0 6914 5 19 1 86689
0 6915 7 2 2 67620 86691
0 6916 5 2 1 86710
0 6917 7 2 2 70253 78307
0 6918 5 2 1 86714
0 6919 7 1 2 86492 86716
0 6920 5 1 1 6919
0 6921 7 1 2 71204 6920
0 6922 5 1 1 6921
0 6923 7 1 2 86712 6922
0 6924 5 1 1 6923
0 6925 7 1 2 84625 6924
0 6926 5 1 1 6925
0 6927 7 4 2 68781 72104
0 6928 5 8 1 86718
0 6929 7 8 2 67386 72105
0 6930 5 5 1 86730
0 6931 7 2 2 84667 86738
0 6932 5 1 1 86743
0 6933 7 1 2 86722 86744
0 6934 5 1 1 6933
0 6935 7 1 2 70619 6934
0 6936 5 2 1 6935
0 6937 7 1 2 5743 86745
0 6938 5 1 1 6937
0 6939 7 1 2 67161 6938
0 6940 5 1 1 6939
0 6941 7 2 2 78320 79398
0 6942 7 1 2 74577 86747
0 6943 5 1 1 6942
0 6944 7 2 2 72521 83187
0 6945 5 2 1 86749
0 6946 7 1 2 6943 86751
0 6947 5 1 1 6946
0 6948 7 1 2 73388 6947
0 6949 5 1 1 6948
0 6950 7 1 2 6940 6949
0 6951 7 1 2 6926 6950
0 6952 5 1 1 6951
0 6953 7 1 2 69714 83671
0 6954 7 1 2 82696 6953
0 6955 7 1 2 6952 6954
0 6956 5 1 1 6955
0 6957 7 17 2 61456 67162
0 6958 7 3 2 62011 86753
0 6959 7 3 2 81271 80867
0 6960 7 1 2 75539 86773
0 6961 7 1 2 86770 6960
0 6962 5 1 1 6961
0 6963 7 1 2 6956 6962
0 6964 5 1 1 6963
0 6965 7 1 2 68328 6964
0 6966 5 1 1 6965
0 6967 7 2 2 73291 76488
0 6968 7 1 2 75620 86776
0 6969 5 1 1 6968
0 6970 7 1 2 70620 79896
0 6971 5 1 1 6970
0 6972 7 2 2 62329 85072
0 6973 5 1 1 86778
0 6974 7 1 2 6971 6973
0 6975 5 1 1 6974
0 6976 7 1 2 72522 6975
0 6977 5 1 1 6976
0 6978 7 1 2 85619 6977
0 6979 5 1 1 6978
0 6980 7 1 2 79852 75872
0 6981 7 1 2 6979 6980
0 6982 5 1 1 6981
0 6983 7 1 2 6969 6982
0 6984 5 1 1 6983
0 6985 7 1 2 65071 6984
0 6986 5 1 1 6985
0 6987 7 2 2 65681 84747
0 6988 7 2 2 81355 86780
0 6989 7 1 2 80616 86782
0 6990 5 1 1 6989
0 6991 7 1 2 6986 6990
0 6992 5 1 1 6991
0 6993 7 1 2 70254 6992
0 6994 5 1 1 6993
0 6995 7 2 2 69952 77391
0 6996 7 1 2 67163 84634
0 6997 5 1 1 6996
0 6998 7 1 2 85719 6997
0 6999 5 5 1 6998
0 7000 7 1 2 86692 86786
0 7001 5 1 1 7000
0 7002 7 12 2 70862 85377
0 7003 7 1 2 86791 77877
0 7004 5 1 1 7003
0 7005 7 1 2 7001 7004
0 7006 5 1 1 7005
0 7007 7 1 2 67621 7006
0 7008 5 1 1 7007
0 7009 7 1 2 77838 84934
0 7010 5 5 1 7009
0 7011 7 1 2 73389 86803
0 7012 5 1 1 7011
0 7013 7 1 2 84902 7012
0 7014 5 1 1 7013
0 7015 7 1 2 86356 7014
0 7016 5 1 1 7015
0 7017 7 1 2 7008 7016
0 7018 5 1 1 7017
0 7019 7 1 2 86784 7018
0 7020 5 1 1 7019
0 7021 7 1 2 6994 7020
0 7022 5 1 1 7021
0 7023 7 1 2 85412 7022
0 7024 5 1 1 7023
0 7025 7 1 2 6966 7024
0 7026 5 1 1 7025
0 7027 7 1 2 61757 7026
0 7028 5 1 1 7027
0 7029 7 1 2 61457 81272
0 7030 5 2 1 7029
0 7031 7 1 2 75673 85413
0 7032 5 1 1 7031
0 7033 7 1 2 86808 7032
0 7034 5 1 1 7033
0 7035 7 9 2 65072 76458
0 7036 5 1 1 86810
0 7037 7 2 2 70863 75469
0 7038 7 1 2 86547 86819
0 7039 7 1 2 86811 7038
0 7040 7 1 2 7034 7039
0 7041 5 1 1 7040
0 7042 7 1 2 7028 7041
0 7043 5 1 1 7042
0 7044 7 1 2 84067 7043
0 7045 5 1 1 7044
0 7046 7 1 2 6912 7045
0 7047 7 1 2 6837 7046
0 7048 5 1 1 7047
0 7049 7 1 2 64654 7048
0 7050 5 1 1 7049
0 7051 7 1 2 84136 4545
0 7052 5 1 1 7051
0 7053 7 1 2 85330 7052
0 7054 5 1 1 7053
0 7055 7 3 2 62765 83219
0 7056 7 1 2 83981 86821
0 7057 5 1 1 7056
0 7058 7 1 2 7054 7057
0 7059 5 1 1 7058
0 7060 7 1 2 74702 7059
0 7061 5 1 1 7060
0 7062 7 3 2 74066 84243
0 7063 5 1 1 86824
0 7064 7 1 2 84779 79637
0 7065 7 1 2 86825 7064
0 7066 5 1 1 7065
0 7067 7 1 2 7061 7066
0 7068 5 1 1 7067
0 7069 7 1 2 73390 7068
0 7070 5 1 1 7069
0 7071 7 1 2 84522 82271
0 7072 7 1 2 80095 7071
0 7073 7 1 2 77786 7072
0 7074 5 1 1 7073
0 7075 7 2 2 176 75904
0 7076 5 17 1 86827
0 7077 7 1 2 72106 86829
0 7078 5 3 1 7077
0 7079 7 2 2 70864 84952
0 7080 7 1 2 64071 86849
0 7081 5 1 1 7080
0 7082 7 1 2 86846 7081
0 7083 5 1 1 7082
0 7084 7 1 2 77403 84143
0 7085 7 1 2 7083 7084
0 7086 5 1 1 7085
0 7087 7 1 2 7074 7086
0 7088 5 1 1 7087
0 7089 7 1 2 70255 7088
0 7090 5 1 1 7089
0 7091 7 1 2 7070 7090
0 7092 5 1 1 7091
0 7093 7 1 2 69953 7092
0 7094 5 1 1 7093
0 7095 7 3 2 66876 71721
0 7096 5 2 1 86851
0 7097 7 1 2 74397 76691
0 7098 5 2 1 7097
0 7099 7 1 2 86854 86856
0 7100 5 1 1 7099
0 7101 7 1 2 68782 7100
0 7102 5 1 1 7101
0 7103 7 5 2 65682 86644
0 7104 5 1 1 86858
0 7105 7 1 2 70256 86859
0 7106 5 1 1 7105
0 7107 7 1 2 7102 7106
0 7108 5 1 1 7107
0 7109 7 11 2 68093 69310
0 7110 7 1 2 72107 86863
0 7111 7 1 2 81856 7110
0 7112 7 1 2 7108 7111
0 7113 5 1 1 7112
0 7114 7 1 2 7094 7113
0 7115 5 1 1 7114
0 7116 7 1 2 66643 7115
0 7117 5 1 1 7116
0 7118 7 7 2 69503 86028
0 7119 7 2 2 83539 80279
0 7120 5 1 1 86881
0 7121 7 1 2 74749 86882
0 7122 5 2 1 7121
0 7123 7 6 2 70621 72777
0 7124 5 3 1 86885
0 7125 7 5 2 70257 74104
0 7126 7 3 2 86891 86894
0 7127 7 1 2 66877 86899
0 7128 5 1 1 7127
0 7129 7 1 2 77075 7128
0 7130 5 1 1 7129
0 7131 7 2 2 73391 7130
0 7132 5 1 1 86902
0 7133 7 1 2 81292 86903
0 7134 5 1 1 7133
0 7135 7 1 2 86883 7134
0 7136 5 1 1 7135
0 7137 7 1 2 69715 7136
0 7138 5 1 1 7137
0 7139 7 2 2 78539 73644
0 7140 7 3 2 83220 75448
0 7141 7 1 2 86904 86906
0 7142 5 1 1 7141
0 7143 7 1 2 7138 7142
0 7144 5 1 1 7143
0 7145 7 1 2 86874 7144
0 7146 5 1 1 7145
0 7147 7 1 2 7117 7146
0 7148 5 1 1 7147
0 7149 7 1 2 66375 7148
0 7150 5 1 1 7149
0 7151 7 3 2 65941 78443
0 7152 7 1 2 86228 86542
0 7153 7 1 2 86909 7152
0 7154 5 1 1 7153
0 7155 7 1 2 84806 86369
0 7156 5 1 1 7155
0 7157 7 4 2 62012 85182
0 7158 7 1 2 75643 86912
0 7159 5 1 1 7158
0 7160 7 1 2 7156 7159
0 7161 5 1 1 7160
0 7162 7 1 2 65345 79168
0 7163 7 1 2 7161 7162
0 7164 5 1 1 7163
0 7165 7 1 2 7154 7164
0 7166 5 1 1 7165
0 7167 7 1 2 69954 7166
0 7168 5 1 1 7167
0 7169 7 3 2 65073 73645
0 7170 7 2 2 68094 73728
0 7171 7 17 2 62766 69504
0 7172 5 1 1 86921
0 7173 7 1 2 86922 71040
0 7174 7 1 2 86919 7173
0 7175 7 1 2 86916 7174
0 7176 5 1 1 7175
0 7177 7 1 2 7168 7176
0 7178 5 1 1 7177
0 7179 7 1 2 82837 7178
0 7180 5 1 1 7179
0 7181 7 1 2 63083 7180
0 7182 7 1 2 7150 7181
0 7183 5 1 1 7182
0 7184 7 73 2 61458 64655
0 7185 5 5 1 86938
0 7186 7 7 2 66878 68941
0 7187 7 4 2 62767 83080
0 7188 7 2 2 65074 87023
0 7189 7 1 2 87016 87027
0 7190 5 1 1 7189
0 7191 7 3 2 78057 82727
0 7192 5 1 1 87029
0 7193 7 2 2 72024 84580
0 7194 5 1 1 87032
0 7195 7 1 2 87030 87033
0 7196 5 1 1 7195
0 7197 7 1 2 7190 7196
0 7198 5 1 1 7197
0 7199 7 1 2 65683 7198
0 7200 5 1 1 7199
0 7201 7 2 2 62516 71025
0 7202 5 5 1 87034
0 7203 7 3 2 72025 84564
0 7204 5 2 1 87041
0 7205 7 2 2 87036 87042
0 7206 5 3 1 87046
0 7207 7 1 2 87031 87047
0 7208 5 1 1 7207
0 7209 7 1 2 7200 7208
0 7210 5 1 1 7209
0 7211 7 1 2 86939 7210
0 7212 5 1 1 7211
0 7213 7 2 2 69955 83494
0 7214 7 1 2 81835 86830
0 7215 7 1 2 87051 7214
0 7216 5 1 1 7215
0 7217 7 2 2 66376 78820
0 7218 7 1 2 84120 85471
0 7219 7 1 2 87053 7218
0 7220 5 1 1 7219
0 7221 7 1 2 7216 7220
0 7222 5 1 1 7221
0 7223 7 1 2 66644 7222
0 7224 5 1 1 7223
0 7225 7 3 2 68783 83031
0 7226 7 16 2 69505 65075
0 7227 7 1 2 70622 87058
0 7228 7 1 2 82697 7227
0 7229 7 1 2 87055 7228
0 7230 5 1 1 7229
0 7231 7 1 2 7224 7230
0 7232 5 1 1 7231
0 7233 7 1 2 72108 7232
0 7234 5 1 1 7233
0 7235 7 3 2 69506 76547
0 7236 7 4 2 73392 85331
0 7237 7 1 2 84846 87077
0 7238 5 1 1 7237
0 7239 7 3 2 66879 81293
0 7240 5 1 1 87081
0 7241 7 1 2 84913 87082
0 7242 5 1 1 7241
0 7243 7 1 2 7238 7242
0 7244 5 1 1 7243
0 7245 7 1 2 87074 7244
0 7246 5 1 1 7245
0 7247 7 1 2 7234 7246
0 7248 7 1 2 7212 7247
0 7249 5 1 1 7248
0 7250 7 1 2 64875 7249
0 7251 5 1 1 7250
0 7252 7 4 2 61758 78650
0 7253 7 11 2 63256 70623
0 7254 7 2 2 64656 87088
0 7255 7 1 2 87084 87099
0 7256 5 1 1 7255
0 7257 7 2 2 66645 81546
0 7258 7 14 2 63909 69507
0 7259 7 1 2 65684 87103
0 7260 7 1 2 87101 7259
0 7261 5 1 1 7260
0 7262 7 1 2 7256 7261
0 7263 5 1 1 7262
0 7264 7 1 2 66377 7263
0 7265 5 1 1 7264
0 7266 7 2 2 61459 70987
0 7267 7 1 2 83376 79925
0 7268 7 1 2 87117 7267
0 7269 5 1 1 7268
0 7270 7 1 2 7265 7269
0 7271 5 1 1 7270
0 7272 7 1 2 72109 7271
0 7273 5 1 1 7272
0 7274 7 1 2 72930 73248
0 7275 5 2 1 7274
0 7276 7 2 2 72714 87119
0 7277 5 1 1 87121
0 7278 7 1 2 71566 87122
0 7279 5 5 1 7278
0 7280 7 2 2 70865 87123
0 7281 5 1 1 87128
0 7282 7 6 2 66880 64657
0 7283 7 2 2 82364 87130
0 7284 7 7 2 66378 64072
0 7285 7 1 2 87136 87138
0 7286 7 1 2 87129 7285
0 7287 5 1 1 7286
0 7288 7 1 2 7273 7287
0 7289 5 1 1 7288
0 7290 7 1 2 78588 7289
0 7291 5 1 1 7290
0 7292 7 1 2 70258 7291
0 7293 7 1 2 7251 7292
0 7294 5 1 1 7293
0 7295 7 1 2 86783 87137
0 7296 5 1 1 7295
0 7297 7 1 2 83403 79620
0 7298 5 1 1 7297
0 7299 7 1 2 7120 7298
0 7300 5 1 1 7299
0 7301 7 1 2 73292 7300
0 7302 5 1 1 7301
0 7303 7 2 2 85284 84550
0 7304 5 4 1 87145
0 7305 7 5 2 73393 87146
0 7306 5 2 1 87151
0 7307 7 2 2 66881 83208
0 7308 7 1 2 87152 87158
0 7309 5 1 1 7308
0 7310 7 1 2 80702 84256
0 7311 5 1 1 7310
0 7312 7 1 2 7309 7311
0 7313 5 1 1 7312
0 7314 7 1 2 82860 7313
0 7315 5 1 1 7314
0 7316 7 1 2 7302 7315
0 7317 5 1 1 7316
0 7318 7 1 2 78277 7317
0 7319 5 1 1 7318
0 7320 7 1 2 7296 7319
0 7321 5 1 1 7320
0 7322 7 1 2 66379 7321
0 7323 5 1 1 7322
0 7324 7 3 2 68784 78589
0 7325 7 1 2 86731 81579
0 7326 7 1 2 87160 7325
0 7327 5 1 1 7326
0 7328 7 6 2 64876 73394
0 7329 7 5 2 67622 83221
0 7330 7 1 2 87169 87159
0 7331 7 1 2 87163 7330
0 7332 5 1 1 7331
0 7333 7 1 2 7327 7332
0 7334 5 1 1 7333
0 7335 7 4 2 61460 65685
0 7336 7 1 2 78980 87174
0 7337 7 1 2 7334 7336
0 7338 5 1 1 7337
0 7339 7 1 2 65346 7338
0 7340 7 1 2 7323 7339
0 7341 5 1 1 7340
0 7342 7 1 2 69311 7341
0 7343 7 1 2 7294 7342
0 7344 5 1 1 7343
0 7345 7 1 2 76022 85276
0 7346 5 1 1 7345
0 7347 7 1 2 7132 7346
0 7348 5 1 1 7347
0 7349 7 1 2 81294 7348
0 7350 5 1 1 7349
0 7351 7 1 2 86884 7350
0 7352 5 1 1 7351
0 7353 7 1 2 61759 7352
0 7354 5 1 1 7353
0 7355 7 1 2 84652 80280
0 7356 5 1 1 7355
0 7357 7 1 2 63490 85342
0 7358 5 1 1 7357
0 7359 7 1 2 7356 7358
0 7360 5 1 1 7359
0 7361 7 4 2 66646 83672
0 7362 7 1 2 70259 87178
0 7363 7 1 2 7360 7362
0 7364 5 1 1 7363
0 7365 7 1 2 7354 7364
0 7366 5 1 1 7365
0 7367 7 1 2 69716 7366
0 7368 5 1 1 7367
0 7369 7 5 2 62768 74350
0 7370 5 2 1 87182
0 7371 7 1 2 2701 87187
0 7372 5 1 1 7371
0 7373 7 3 2 65942 79597
0 7374 7 2 2 71041 83222
0 7375 7 1 2 87189 87192
0 7376 7 1 2 7372 7375
0 7377 5 1 1 7376
0 7378 7 1 2 7368 7377
0 7379 5 1 1 7378
0 7380 7 1 2 83947 7379
0 7381 5 1 1 7380
0 7382 7 1 2 67953 7381
0 7383 7 1 2 7344 7382
0 7384 5 1 1 7383
0 7385 7 1 2 72974 7384
0 7386 7 1 2 7183 7385
0 7387 5 1 1 7386
0 7388 7 1 2 7050 7387
0 7389 7 1 2 6556 7388
0 7390 7 1 2 5791 7389
0 7391 5 1 1 7390
0 7392 7 1 2 61254 7391
0 7393 5 1 1 7392
0 7394 7 19 2 67623 63257
0 7395 7 2 2 79340 71688
0 7396 7 1 2 87194 87213
0 7397 5 1 1 7396
0 7398 7 1 2 84144 82165
0 7399 5 1 1 7398
0 7400 7 1 2 7397 7399
0 7401 5 1 1 7400
0 7402 7 1 2 66647 7401
0 7403 5 1 1 7402
0 7404 7 1 2 81497 87214
0 7405 5 1 1 7404
0 7406 7 1 2 7403 7405
0 7407 5 1 1 7406
0 7408 7 1 2 68942 7407
0 7409 5 1 1 7408
0 7410 7 2 2 69312 76314
0 7411 7 1 2 68095 78988
0 7412 7 1 2 87215 7411
0 7413 5 1 1 7412
0 7414 7 1 2 7409 7413
0 7415 5 1 1 7414
0 7416 7 1 2 70260 7415
0 7417 5 1 1 7416
0 7418 7 5 2 65347 74174
0 7419 7 2 2 78471 87217
0 7420 7 1 2 86299 82728
0 7421 7 1 2 87222 7420
0 7422 5 1 1 7421
0 7423 7 1 2 7417 7422
0 7424 5 1 1 7423
0 7425 7 1 2 76118 7424
0 7426 5 1 1 7425
0 7427 7 1 2 84033 86717
0 7428 5 1 1 7427
0 7429 7 1 2 79169 7428
0 7430 5 1 1 7429
0 7431 7 2 2 73535 78278
0 7432 5 1 1 87224
0 7433 7 1 2 85378 87225
0 7434 5 1 1 7433
0 7435 7 1 2 7430 7434
0 7436 5 1 1 7435
0 7437 7 1 2 85649 7436
0 7438 5 1 1 7437
0 7439 7 1 2 7426 7438
0 7440 5 1 1 7439
0 7441 7 1 2 72975 7440
0 7442 5 1 1 7441
0 7443 7 4 2 64073 74777
0 7444 7 2 2 74195 87226
0 7445 5 1 1 87230
0 7446 7 1 2 78997 87231
0 7447 5 1 1 7446
0 7448 7 7 2 64658 72110
0 7449 7 5 2 61760 75348
0 7450 5 1 1 87239
0 7451 7 1 2 76018 7450
0 7452 5 14 1 7451
0 7453 7 1 2 66380 87244
0 7454 5 1 1 7453
0 7455 7 2 2 76036 78836
0 7456 5 1 1 87258
0 7457 7 1 2 7454 7456
0 7458 5 1 1 7457
0 7459 7 1 2 87232 7458
0 7460 5 1 1 7459
0 7461 7 6 2 67954 76548
0 7462 7 1 2 81218 87260
0 7463 5 1 1 7462
0 7464 7 1 2 7460 7463
0 7465 5 1 1 7464
0 7466 7 1 2 65348 82691
0 7467 7 1 2 7465 7466
0 7468 5 1 1 7467
0 7469 7 1 2 7447 7468
0 7470 5 1 1 7469
0 7471 7 1 2 69313 7470
0 7472 5 1 1 7471
0 7473 7 3 2 76119 84653
0 7474 7 3 2 79341 76771
0 7475 7 1 2 76459 87269
0 7476 7 2 2 87266 7475
0 7477 5 1 1 87272
0 7478 7 1 2 61761 87273
0 7479 5 1 1 7478
0 7480 7 1 2 7472 7479
0 7481 5 1 1 7480
0 7482 7 1 2 68096 7481
0 7483 5 1 1 7482
0 7484 7 1 2 63491 80468
0 7485 7 1 2 74196 7484
0 7486 7 6 2 66381 80434
0 7487 7 1 2 83625 87274
0 7488 7 1 2 7485 7487
0 7489 5 1 1 7488
0 7490 7 1 2 7477 7489
0 7491 5 1 1 7490
0 7492 7 1 2 81437 7491
0 7493 5 1 1 7492
0 7494 7 1 2 7483 7493
0 7495 7 1 2 7442 7494
0 7496 5 1 1 7495
0 7497 7 1 2 69956 7496
0 7498 5 1 1 7497
0 7499 7 2 2 86754 84334
0 7500 7 2 2 74612 79805
0 7501 7 1 2 87280 87282
0 7502 5 1 1 7501
0 7503 7 3 2 70624 75248
0 7504 7 1 2 87284 87139
0 7505 7 1 2 76856 7504
0 7506 5 1 1 7505
0 7507 7 1 2 7502 7506
0 7508 5 1 1 7507
0 7509 7 1 2 83081 7508
0 7510 5 1 1 7509
0 7511 7 2 2 64877 76518
0 7512 7 1 2 81836 85500
0 7513 7 1 2 86525 7512
0 7514 7 1 2 87287 7513
0 7515 5 1 1 7514
0 7516 7 1 2 7510 7515
0 7517 5 1 1 7516
0 7518 7 1 2 64659 7517
0 7519 5 1 1 7518
0 7520 7 2 2 70625 86526
0 7521 7 2 2 72778 78279
0 7522 5 1 1 87291
0 7523 7 1 2 85637 87292
0 7524 7 1 2 87289 7523
0 7525 5 1 1 7524
0 7526 7 1 2 7519 7525
0 7527 5 1 1 7526
0 7528 7 1 2 69314 7527
0 7529 5 1 1 7528
0 7530 7 7 2 67164 82128
0 7531 5 1 1 87293
0 7532 7 2 2 77456 87294
0 7533 5 1 1 87300
0 7534 7 1 2 83992 87301
0 7535 5 1 1 7534
0 7536 7 1 2 7529 7535
0 7537 5 1 1 7536
0 7538 7 1 2 65076 7537
0 7539 5 1 1 7538
0 7540 7 15 2 69717 83082
0 7541 7 17 2 61461 79342
0 7542 5 6 1 87317
0 7543 7 1 2 85836 87318
0 7544 5 1 1 7543
0 7545 7 2 2 65686 82105
0 7546 7 1 2 87233 87340
0 7547 5 1 1 7546
0 7548 7 1 2 7544 7547
0 7549 5 1 1 7548
0 7550 7 1 2 87302 7549
0 7551 5 1 1 7550
0 7552 7 6 2 68097 76549
0 7553 7 1 2 82818 78308
0 7554 7 1 2 87342 7553
0 7555 5 1 1 7554
0 7556 7 1 2 7551 7555
0 7557 5 1 1 7556
0 7558 7 1 2 86533 7557
0 7559 5 1 1 7558
0 7560 7 1 2 67955 7559
0 7561 7 1 2 7539 7560
0 7562 5 1 1 7561
0 7563 7 2 2 81973 87011
0 7564 5 34 1 87348
0 7565 7 4 2 69718 87350
0 7566 7 1 2 82049 80868
0 7567 5 1 1 7566
0 7568 7 7 2 74260 71773
0 7569 5 2 1 87388
0 7570 7 16 2 66382 62769
0 7571 5 1 1 87397
0 7572 7 1 2 87389 7571
0 7573 5 1 1 7572
0 7574 7 1 2 7567 7573
0 7575 5 1 1 7574
0 7576 7 1 2 87384 7575
0 7577 5 1 1 7576
0 7578 7 10 2 65077 79067
0 7579 7 7 2 66648 68570
0 7580 7 1 2 86755 87423
0 7581 7 1 2 87413 7580
0 7582 5 1 1 7581
0 7583 7 1 2 7577 7582
0 7584 5 1 1 7583
0 7585 7 1 2 64458 7584
0 7586 5 1 1 7585
0 7587 7 2 2 83626 86582
0 7588 5 1 1 87430
0 7589 7 1 2 66383 75682
0 7590 7 1 2 87431 7589
0 7591 5 1 1 7590
0 7592 7 1 2 7586 7591
0 7593 5 1 1 7592
0 7594 7 1 2 63258 7593
0 7595 5 1 1 7594
0 7596 7 11 2 63492 71808
0 7597 5 1 1 87432
0 7598 7 1 2 86132 87433
0 7599 5 1 1 7598
0 7600 7 1 2 7588 7599
0 7601 5 1 1 7600
0 7602 7 1 2 61762 7601
0 7603 5 1 1 7602
0 7604 7 1 2 76832 83562
0 7605 5 1 1 7604
0 7606 7 1 2 7603 7605
0 7607 5 1 1 7606
0 7608 7 1 2 66384 81322
0 7609 7 1 2 7607 7608
0 7610 5 1 1 7609
0 7611 7 1 2 7595 7610
0 7612 5 1 1 7611
0 7613 7 1 2 77457 7612
0 7614 5 1 1 7613
0 7615 7 3 2 70261 86812
0 7616 7 6 2 66649 64074
0 7617 7 3 2 87446 74234
0 7618 5 1 1 87452
0 7619 7 1 2 70866 81691
0 7620 7 1 2 87351 7619
0 7621 7 1 2 87453 7620
0 7622 7 1 2 87443 7621
0 7623 5 1 1 7622
0 7624 7 1 2 63084 7623
0 7625 7 1 2 7614 7624
0 7626 5 1 1 7625
0 7627 7 1 2 7562 7626
0 7628 5 1 1 7627
0 7629 7 5 2 67165 76550
0 7630 7 11 2 69315 65078
0 7631 7 6 2 65349 72111
0 7632 5 1 1 87471
0 7633 7 1 2 87460 87472
0 7634 7 1 2 87455 7633
0 7635 5 1 1 7634
0 7636 7 10 2 61462 62770
0 7637 7 2 2 87477 74246
0 7638 7 15 2 64459 70262
0 7639 7 1 2 84443 87489
0 7640 7 1 2 87487 7639
0 7641 5 1 1 7640
0 7642 7 1 2 7635 7641
0 7643 5 1 1 7642
0 7644 7 1 2 65687 7643
0 7645 5 1 1 7644
0 7646 7 4 2 84054 87190
0 7647 7 2 2 67166 73941
0 7648 5 2 1 87508
0 7649 7 1 2 83281 87510
0 7650 7 1 2 87504 7649
0 7651 5 1 1 7650
0 7652 7 1 2 7645 7651
0 7653 5 1 1 7652
0 7654 7 1 2 68571 7653
0 7655 5 1 1 7654
0 7656 7 2 2 63493 76879
0 7657 5 1 1 87512
0 7658 7 1 2 81059 86390
0 7659 5 1 1 7658
0 7660 7 1 2 2308 7659
0 7661 5 1 1 7660
0 7662 7 1 2 63720 7661
0 7663 5 1 1 7662
0 7664 7 1 2 7657 7663
0 7665 5 1 1 7664
0 7666 7 5 2 65943 84055
0 7667 7 1 2 83282 87514
0 7668 7 1 2 7665 7667
0 7669 5 1 1 7668
0 7670 7 1 2 7655 7669
0 7671 5 1 1 7670
0 7672 7 1 2 81721 79068
0 7673 5 1 1 7672
0 7674 7 3 2 63085 83377
0 7675 7 1 2 69719 87519
0 7676 5 1 1 7675
0 7677 7 1 2 7673 7676
0 7678 5 4 1 7677
0 7679 7 1 2 7671 87522
0 7680 5 1 1 7679
0 7681 7 1 2 7628 7680
0 7682 7 1 2 7498 7681
0 7683 5 1 1 7682
0 7684 7 1 2 62013 7683
0 7685 5 1 1 7684
0 7686 7 3 2 84006 76519
0 7687 5 1 1 87526
0 7688 7 1 2 76037 87527
0 7689 5 1 1 7688
0 7690 7 1 2 70263 87267
0 7691 5 1 1 7690
0 7692 7 1 2 7689 7691
0 7693 5 1 1 7692
0 7694 7 1 2 84479 7693
0 7695 5 1 1 7694
0 7696 7 2 2 75674 82729
0 7697 7 2 2 73060 79210
0 7698 7 1 2 87529 87531
0 7699 5 1 1 7698
0 7700 7 1 2 7695 7699
0 7701 5 1 1 7700
0 7702 7 1 2 81042 7701
0 7703 5 1 1 7702
0 7704 7 3 2 77404 84496
0 7705 5 1 1 87533
0 7706 7 1 2 82730 87534
0 7707 7 1 2 87532 7706
0 7708 5 1 1 7707
0 7709 7 1 2 7703 7708
0 7710 5 1 1 7709
0 7711 7 1 2 72976 7710
0 7712 5 1 1 7711
0 7713 7 1 2 87447 77680
0 7714 5 1 1 7713
0 7715 7 2 2 61763 87288
0 7716 5 1 1 87536
0 7717 7 1 2 7714 7716
0 7718 5 1 1 7717
0 7719 7 3 2 74778 80025
0 7720 7 6 2 68098 87538
0 7721 7 2 2 61463 87541
0 7722 7 1 2 85489 87547
0 7723 7 1 2 7718 7722
0 7724 5 1 1 7723
0 7725 7 1 2 7712 7724
0 7726 5 1 1 7725
0 7727 7 1 2 69316 7726
0 7728 5 1 1 7727
0 7729 7 3 2 62330 78492
0 7730 7 2 2 86331 87549
0 7731 7 10 2 62771 63259
0 7732 7 4 2 87554 80406
0 7733 7 9 2 63721 70867
0 7734 7 1 2 87568 84510
0 7735 7 1 2 87564 7734
0 7736 7 1 2 87552 7735
0 7737 5 1 1 7736
0 7738 7 1 2 7728 7737
0 7739 5 1 1 7738
0 7740 7 1 2 64660 7739
0 7741 5 1 1 7740
0 7742 7 1 2 61464 81790
0 7743 5 1 1 7742
0 7744 7 3 2 63260 78058
0 7745 7 1 2 76068 87577
0 7746 5 1 1 7745
0 7747 7 1 2 7743 7746
0 7748 5 4 1 7747
0 7749 7 1 2 74414 87580
0 7750 5 1 1 7749
0 7751 7 2 2 63261 76880
0 7752 7 3 2 74261 80832
0 7753 7 1 2 63086 87586
0 7754 7 1 2 87584 7753
0 7755 5 1 1 7754
0 7756 7 1 2 7750 7755
0 7757 5 1 1 7756
0 7758 7 1 2 71476 7757
0 7759 5 1 1 7758
0 7760 7 4 2 61764 70626
0 7761 7 1 2 86432 86157
0 7762 7 1 2 87589 7761
0 7763 7 1 2 87581 7762
0 7764 5 1 1 7763
0 7765 7 1 2 7759 7764
0 7766 5 1 1 7765
0 7767 7 1 2 72523 7766
0 7768 5 1 1 7767
0 7769 7 2 2 72026 86433
0 7770 7 1 2 76428 82166
0 7771 7 1 2 87582 7770
0 7772 5 1 1 7771
0 7773 7 4 2 63722 78590
0 7774 7 1 2 83564 87595
0 7775 7 1 2 86590 7774
0 7776 5 1 1 7775
0 7777 7 1 2 7772 7776
0 7778 5 1 1 7777
0 7779 7 1 2 87593 7778
0 7780 5 1 1 7779
0 7781 7 1 2 7768 7780
0 7782 5 1 1 7781
0 7783 7 1 2 64460 7782
0 7784 5 1 1 7783
0 7785 7 1 2 70627 82063
0 7786 5 1 1 7785
0 7787 7 1 2 7705 7786
0 7788 5 1 1 7787
0 7789 7 1 2 62772 7788
0 7790 5 1 1 7789
0 7791 7 8 2 68329 78591
0 7792 5 5 1 87599
0 7793 7 1 2 87607 78576
0 7794 5 17 1 7793
0 7795 7 1 2 73771 87612
0 7796 5 1 1 7795
0 7797 7 1 2 7790 7796
0 7798 5 1 1 7797
0 7799 7 1 2 84843 7798
0 7800 5 1 1 7799
0 7801 7 3 2 78671 83404
0 7802 5 1 1 87629
0 7803 7 1 2 87630 86886
0 7804 5 1 1 7803
0 7805 7 1 2 7800 7804
0 7806 5 1 1 7805
0 7807 7 1 2 76797 7806
0 7808 5 1 1 7807
0 7809 7 2 2 84882 85490
0 7810 5 1 1 87632
0 7811 7 1 2 80563 81547
0 7812 7 1 2 87633 7811
0 7813 5 1 1 7812
0 7814 7 1 2 7808 7813
0 7815 5 1 1 7814
0 7816 7 1 2 80964 79796
0 7817 7 1 2 7815 7816
0 7818 5 1 1 7817
0 7819 7 1 2 7784 7818
0 7820 5 1 1 7819
0 7821 7 1 2 69508 7820
0 7822 5 1 1 7821
0 7823 7 1 2 7741 7822
0 7824 7 1 2 7685 7823
0 7825 5 1 1 7824
0 7826 7 1 2 61255 7825
0 7827 5 1 1 7826
0 7828 7 18 2 63262 63723
0 7829 7 9 2 87634 80407
0 7830 7 6 2 62331 87652
0 7831 7 3 2 84444 87285
0 7832 7 1 2 61765 80182
0 7833 7 7 2 62014 69317
0 7834 7 13 2 66085 61465
0 7835 7 1 2 87670 87677
0 7836 7 1 2 7832 7835
0 7837 7 1 2 87667 7836
0 7838 7 1 2 87661 7837
0 7839 5 1 1 7838
0 7840 7 1 2 7827 7839
0 7841 5 1 1 7840
0 7842 7 1 2 71294 7841
0 7843 5 1 1 7842
0 7844 7 1 2 7393 7843
0 7845 5 1 1 7844
0 7846 7 1 2 64312 7845
0 7847 5 1 1 7846
0 7848 7 4 2 61466 82731
0 7849 5 1 1 87690
0 7850 7 5 2 66385 82365
0 7851 5 1 1 87694
0 7852 7 1 2 7849 7851
0 7853 5 7 1 7852
0 7854 7 57 2 61256 64313
0 7855 5 3 1 87706
0 7856 7 6 2 65688 87707
0 7857 5 1 1 87766
0 7858 7 4 2 69157 81869
0 7859 7 1 2 73249 87772
0 7860 5 1 1 7859
0 7861 7 1 2 7857 7860
0 7862 5 1 1 7861
0 7863 7 1 2 72112 7862
0 7864 5 1 1 7863
0 7865 7 43 2 66086 69158
0 7866 7 1 2 79498 87776
0 7867 5 1 1 7866
0 7868 7 1 2 7864 7867
0 7869 5 1 1 7868
0 7870 7 1 2 74651 7869
0 7871 5 1 1 7870
0 7872 7 3 2 66087 74175
0 7873 7 7 2 64075 69159
0 7874 7 1 2 74933 87822
0 7875 7 1 2 87819 7874
0 7876 5 1 1 7875
0 7877 7 1 2 7871 7876
0 7878 5 1 1 7877
0 7879 7 1 2 68572 7878
0 7880 5 1 1 7879
0 7881 7 19 2 69160 70628
0 7882 7 3 2 83302 87829
0 7883 7 1 2 83736 87848
0 7884 5 1 1 7883
0 7885 7 10 2 68785 64314
0 7886 7 1 2 84274 87851
0 7887 5 1 1 7886
0 7888 7 1 2 7884 7887
0 7889 5 1 1 7888
0 7890 7 1 2 79836 7889
0 7891 5 1 1 7890
0 7892 7 1 2 7880 7891
0 7893 5 1 1 7892
0 7894 7 1 2 67167 7893
0 7895 5 1 1 7894
0 7896 7 1 2 84635 87849
0 7897 5 1 1 7896
0 7898 7 2 2 68573 87852
0 7899 7 1 2 84275 87861
0 7900 5 1 1 7899
0 7901 7 1 2 7897 7900
0 7902 5 1 1 7901
0 7903 7 1 2 79837 7902
0 7904 5 1 1 7903
0 7905 7 1 2 7895 7904
0 7906 5 1 1 7905
0 7907 7 1 2 69720 7906
0 7908 5 1 1 7907
0 7909 7 1 2 71722 73536
0 7910 7 1 2 78814 7909
0 7911 7 6 2 62332 75506
0 7912 7 6 2 63910 69161
0 7913 7 5 2 66088 87869
0 7914 5 1 1 87875
0 7915 7 1 2 87863 87876
0 7916 7 1 2 7910 7915
0 7917 5 1 1 7916
0 7918 7 1 2 7908 7917
0 7919 5 1 1 7918
0 7920 7 1 2 66882 7919
0 7921 5 1 1 7920
0 7922 7 1 2 64076 80159
0 7923 5 1 1 7922
0 7924 7 1 2 76339 77292
0 7925 5 1 1 7924
0 7926 7 1 2 7923 7925
0 7927 5 1 1 7926
0 7928 7 1 2 65350 7927
0 7929 5 1 1 7928
0 7930 7 3 2 72954 73877
0 7931 5 1 1 87880
0 7932 7 5 2 72977 71567
0 7933 5 3 1 87883
0 7934 7 1 2 77939 87888
0 7935 7 1 2 7931 7934
0 7936 5 1 1 7935
0 7937 7 1 2 7929 7936
0 7938 5 1 1 7937
0 7939 7 8 2 67624 64878
0 7940 7 1 2 75847 87891
0 7941 7 1 2 87777 7940
0 7942 7 1 2 7938 7941
0 7943 5 1 1 7942
0 7944 7 1 2 7921 7943
0 7945 5 1 1 7944
0 7946 7 1 2 84087 7945
0 7947 5 1 1 7946
0 7948 7 5 2 68574 75132
0 7949 5 1 1 87899
0 7950 7 2 2 67168 87900
0 7951 7 1 2 71465 87904
0 7952 5 1 1 7951
0 7953 7 2 2 72691 71521
0 7954 5 3 1 87906
0 7955 7 2 2 64879 87908
0 7956 7 1 2 77640 87911
0 7957 5 1 1 7956
0 7958 7 1 2 7952 7957
0 7959 5 1 1 7958
0 7960 7 1 2 87708 7959
0 7961 5 1 1 7960
0 7962 7 1 2 66883 74913
0 7963 5 1 1 7962
0 7964 7 1 2 7963 3122
0 7965 5 2 1 7964
0 7966 7 1 2 87913 73250
0 7967 5 1 1 7966
0 7968 7 1 2 66884 75567
0 7969 5 1 1 7968
0 7970 7 1 2 7967 7969
0 7971 5 1 1 7970
0 7972 7 1 2 71466 7971
0 7973 5 1 1 7972
0 7974 7 1 2 84565 87037
0 7975 5 3 1 7974
0 7976 7 1 2 63494 87915
0 7977 5 1 1 7976
0 7978 7 2 2 77793 77596
0 7979 5 1 1 87918
0 7980 7 1 2 7977 7979
0 7981 5 1 1 7980
0 7982 7 1 2 62015 82167
0 7983 7 1 2 7981 7982
0 7984 5 1 1 7983
0 7985 7 1 2 7973 7984
0 7986 5 1 1 7985
0 7987 7 1 2 87778 7986
0 7988 5 1 1 7987
0 7989 7 1 2 7961 7988
0 7990 5 1 1 7989
0 7991 7 1 2 65944 7990
0 7992 5 1 1 7991
0 7993 7 9 2 69162 65689
0 7994 7 3 2 68786 87920
0 7995 7 1 2 83198 87929
0 7996 5 1 1 7995
0 7997 7 4 2 61257 62773
0 7998 7 9 2 64315 73395
0 7999 7 1 2 87932 87936
0 8000 5 1 1 7999
0 8001 7 1 2 7996 8000
0 8002 5 1 1 8001
0 8003 7 1 2 74779 8002
0 8004 5 1 1 8003
0 8005 7 9 2 70629 73293
0 8006 5 7 1 87945
0 8007 7 3 2 64316 87933
0 8008 7 1 2 87954 87961
0 8009 5 1 1 8008
0 8010 7 1 2 76496 76407
0 8011 5 1 1 8010
0 8012 7 1 2 68575 8011
0 8013 5 1 1 8012
0 8014 7 2 2 62774 83758
0 8015 5 3 1 87964
0 8016 7 6 2 63724 65690
0 8017 5 1 1 87969
0 8018 7 1 2 87966 8017
0 8019 5 1 1 8018
0 8020 7 1 2 67387 8019
0 8021 5 1 1 8020
0 8022 7 1 2 71625 8021
0 8023 7 1 2 8013 8022
0 8024 5 1 1 8023
0 8025 7 1 2 87779 8024
0 8026 5 1 1 8025
0 8027 7 1 2 8009 8026
0 8028 5 1 1 8027
0 8029 7 1 2 68330 8028
0 8030 5 1 1 8029
0 8031 7 1 2 8004 8030
0 8032 5 1 1 8031
0 8033 7 1 2 66885 8032
0 8034 5 1 1 8033
0 8035 7 2 2 74780 75433
0 8036 7 1 2 81706 87921
0 8037 7 1 2 87975 8036
0 8038 5 1 1 8037
0 8039 7 1 2 8034 8038
0 8040 5 1 1 8039
0 8041 7 1 2 69721 8040
0 8042 5 1 1 8041
0 8043 7 1 2 7992 8042
0 8044 5 1 1 8043
0 8045 7 1 2 68943 8044
0 8046 5 1 1 8045
0 8047 7 1 2 73560 82224
0 8048 5 1 1 8047
0 8049 7 2 2 67169 75662
0 8050 5 1 1 87977
0 8051 7 1 2 8050 77732
0 8052 5 1 1 8051
0 8053 7 1 2 73537 8052
0 8054 5 1 1 8053
0 8055 7 2 2 63911 84335
0 8056 5 1 1 87979
0 8057 7 2 2 65691 73561
0 8058 5 4 1 87981
0 8059 7 1 2 84615 73942
0 8060 7 1 2 87983 8059
0 8061 5 1 1 8060
0 8062 7 1 2 8056 8061
0 8063 7 1 2 8054 8062
0 8064 5 1 1 8063
0 8065 7 1 2 68331 8064
0 8066 5 1 1 8065
0 8067 7 3 2 62775 77808
0 8068 5 3 1 87987
0 8069 7 1 2 67388 82535
0 8070 7 1 2 87988 8069
0 8071 5 1 1 8070
0 8072 7 1 2 8066 8071
0 8073 5 1 1 8072
0 8074 7 1 2 64077 8073
0 8075 5 1 1 8074
0 8076 7 1 2 8048 8075
0 8077 5 1 1 8076
0 8078 7 1 2 87780 8077
0 8079 5 1 1 8078
0 8080 7 2 2 68787 74858
0 8081 7 1 2 85404 87993
0 8082 5 1 1 8081
0 8083 7 1 2 71908 79827
0 8084 5 1 1 8083
0 8085 7 1 2 8082 8084
0 8086 5 1 1 8085
0 8087 7 1 2 67625 8086
0 8088 5 1 1 8087
0 8089 7 1 2 71909 74105
0 8090 7 1 2 73787 8089
0 8091 5 1 1 8090
0 8092 7 1 2 62776 85795
0 8093 5 1 1 8092
0 8094 7 1 2 8091 8093
0 8095 5 1 1 8094
0 8096 7 1 2 68332 8095
0 8097 5 1 1 8096
0 8098 7 1 2 8088 8097
0 8099 5 1 1 8098
0 8100 7 1 2 67389 8099
0 8101 5 1 1 8100
0 8102 7 3 2 68788 79677
0 8103 5 1 1 87995
0 8104 7 1 2 71137 8103
0 8105 5 1 1 8104
0 8106 7 1 2 76440 73251
0 8107 7 1 2 8105 8106
0 8108 5 1 1 8107
0 8109 7 1 2 8101 8108
0 8110 5 1 1 8109
0 8111 7 1 2 87709 8110
0 8112 5 1 1 8111
0 8113 7 1 2 73538 87227
0 8114 5 2 1 8113
0 8115 7 1 2 84888 74998
0 8116 5 2 1 8115
0 8117 7 1 2 86169 86892
0 8118 7 1 2 88000 8117
0 8119 5 1 1 8118
0 8120 7 1 2 87998 8119
0 8121 5 1 1 8120
0 8122 7 2 2 68333 87781
0 8123 7 1 2 88002 87955
0 8124 7 1 2 8121 8123
0 8125 5 1 1 8124
0 8126 7 2 2 8112 8125
0 8127 7 2 2 64078 87124
0 8128 5 1 1 88006
0 8129 7 1 2 6000 8128
0 8130 5 1 1 8129
0 8131 7 1 2 68334 8130
0 8132 5 1 1 8131
0 8133 7 1 2 74781 87078
0 8134 5 1 1 8133
0 8135 7 1 2 8132 8134
0 8136 5 1 1 8135
0 8137 7 1 2 87710 8136
0 8138 5 1 1 8137
0 8139 7 1 2 88004 8138
0 8140 7 1 2 8079 8139
0 8141 5 1 1 8140
0 8142 7 1 2 77392 8141
0 8143 5 1 1 8142
0 8144 7 2 2 62016 87782
0 8145 7 2 2 73562 75050
0 8146 7 2 2 65692 79471
0 8147 5 2 1 88012
0 8148 7 1 2 88010 88013
0 8149 5 1 1 8148
0 8150 7 1 2 73711 74962
0 8151 5 1 1 8150
0 8152 7 1 2 8149 8151
0 8153 5 1 1 8152
0 8154 7 1 2 68576 8153
0 8155 5 1 1 8154
0 8156 7 2 2 76843 79678
0 8157 7 1 2 71809 85352
0 8158 7 1 2 88016 8157
0 8159 5 1 1 8158
0 8160 7 1 2 8155 8159
0 8161 5 1 1 8160
0 8162 7 1 2 88008 8161
0 8163 5 1 1 8162
0 8164 7 1 2 65351 8163
0 8165 7 1 2 8143 8164
0 8166 7 1 2 8046 8165
0 8167 5 1 1 8166
0 8168 7 3 2 72524 87711
0 8169 7 1 2 74859 88018
0 8170 5 1 1 8169
0 8171 7 2 2 76441 87783
0 8172 5 1 1 88021
0 8173 7 1 2 8170 8172
0 8174 5 1 1 8173
0 8175 7 1 2 67626 8174
0 8176 5 1 1 8175
0 8177 7 1 2 86015 88003
0 8178 5 1 1 8177
0 8179 7 1 2 8176 8178
0 8180 5 1 1 8179
0 8181 7 1 2 65693 8180
0 8182 5 1 1 8181
0 8183 7 1 2 84654 88022
0 8184 5 1 1 8183
0 8185 7 1 2 8182 8184
0 8186 5 1 1 8185
0 8187 7 1 2 73396 8186
0 8188 5 1 1 8187
0 8189 7 1 2 69163 83303
0 8190 7 1 2 72878 8189
0 8191 7 1 2 84977 8190
0 8192 5 1 1 8191
0 8193 7 1 2 8188 8192
0 8194 7 1 2 88005 8193
0 8195 5 1 1 8194
0 8196 7 1 2 77393 8195
0 8197 5 1 1 8196
0 8198 7 1 2 78170 87784
0 8199 5 1 1 8198
0 8200 7 2 2 86693 87712
0 8201 5 1 1 88023
0 8202 7 1 2 8199 8201
0 8203 5 1 1 8202
0 8204 7 1 2 76270 8203
0 8205 5 1 1 8204
0 8206 7 2 2 61258 73294
0 8207 7 7 2 68944 64317
0 8208 7 1 2 86910 88027
0 8209 7 1 2 88025 8208
0 8210 5 1 1 8209
0 8211 7 1 2 8205 8210
0 8212 5 1 1 8211
0 8213 7 1 2 68577 8212
0 8214 5 1 1 8213
0 8215 7 1 2 87909 88019
0 8216 5 1 1 8215
0 8217 7 1 2 76301 87785
0 8218 5 1 1 8217
0 8219 7 1 2 8216 8218
0 8220 5 1 1 8219
0 8221 7 1 2 72978 8220
0 8222 5 1 1 8221
0 8223 7 1 2 8214 8222
0 8224 5 1 1 8223
0 8225 7 1 2 77081 8224
0 8226 5 1 1 8225
0 8227 7 1 2 70264 8226
0 8228 7 1 2 8197 8227
0 8229 5 1 1 8228
0 8230 7 1 2 81485 8229
0 8231 7 1 2 8167 8230
0 8232 5 1 1 8231
0 8233 7 1 2 7947 8232
0 8234 5 1 1 8233
0 8235 7 1 2 69957 8234
0 8236 5 1 1 8235
0 8237 7 1 2 68335 73629
0 8238 5 2 1 8237
0 8239 7 1 2 77082 88034
0 8240 5 1 1 8239
0 8241 7 1 2 77928 72368
0 8242 7 1 2 82392 8241
0 8243 5 1 1 8242
0 8244 7 1 2 8240 8243
0 8245 5 1 1 8244
0 8246 7 1 2 77433 8245
0 8247 5 1 1 8246
0 8248 7 10 2 69722 74305
0 8249 7 1 2 80495 88036
0 8250 5 1 1 8249
0 8251 7 1 2 8247 8250
0 8252 5 1 1 8251
0 8253 7 1 2 63725 8252
0 8254 5 1 1 8253
0 8255 7 1 2 63495 80313
0 8256 5 1 1 8255
0 8257 7 1 2 8254 8256
0 8258 5 1 1 8257
0 8259 7 1 2 67627 8258
0 8260 5 1 1 8259
0 8261 7 2 2 77405 72912
0 8262 7 1 2 62017 88046
0 8263 7 1 2 80424 8262
0 8264 5 1 1 8263
0 8265 7 1 2 8260 8264
0 8266 5 1 1 8265
0 8267 7 1 2 78128 8266
0 8268 5 1 1 8267
0 8269 7 5 2 64880 74262
0 8270 5 1 1 88048
0 8271 7 3 2 62018 77434
0 8272 7 1 2 63912 88053
0 8273 7 1 2 88049 8272
0 8274 7 1 2 86826 8273
0 8275 5 1 1 8274
0 8276 7 1 2 8268 8275
0 8277 5 1 1 8276
0 8278 7 1 2 84088 8277
0 8279 5 1 1 8278
0 8280 7 3 2 79069 84056
0 8281 7 1 2 63087 76534
0 8282 7 1 2 88056 8281
0 8283 7 1 2 76755 8282
0 8284 5 1 1 8283
0 8285 7 1 2 8279 8284
0 8286 5 1 1 8285
0 8287 7 1 2 87786 8286
0 8288 5 1 1 8287
0 8289 7 3 2 72113 72979
0 8290 7 1 2 67956 79761
0 8291 7 1 2 88059 8290
0 8292 5 1 1 8291
0 8293 7 2 2 81468 84511
0 8294 5 1 1 88062
0 8295 7 1 2 70868 77468
0 8296 7 1 2 85858 8295
0 8297 7 1 2 88063 8296
0 8298 5 1 1 8297
0 8299 7 1 2 8292 8298
0 8300 5 1 1 8299
0 8301 7 1 2 70630 8300
0 8302 5 1 1 8301
0 8303 7 1 2 76643 79279
0 8304 7 1 2 78309 8303
0 8305 7 1 2 79762 8304
0 8306 5 1 1 8305
0 8307 7 1 2 8302 8306
0 8308 5 1 1 8307
0 8309 7 1 2 70265 8308
0 8310 5 1 1 8309
0 8311 7 2 2 80064 84919
0 8312 5 1 1 88064
0 8313 7 4 2 62333 79280
0 8314 7 1 2 88066 78321
0 8315 7 1 2 85661 8314
0 8316 7 1 2 8312 8315
0 8317 5 1 1 8316
0 8318 7 1 2 8310 8317
0 8319 5 1 1 8318
0 8320 7 1 2 69723 8319
0 8321 5 1 1 8320
0 8322 7 4 2 80799 84207
0 8323 7 1 2 72525 88070
0 8324 7 7 2 67170 72692
0 8325 5 2 1 88074
0 8326 7 1 2 87414 88075
0 8327 7 1 2 8323 8326
0 8328 5 1 1 8327
0 8329 7 1 2 8321 8328
0 8330 5 1 1 8329
0 8331 7 1 2 68789 8330
0 8332 5 1 1 8331
0 8333 7 3 2 67171 75449
0 8334 5 1 1 88083
0 8335 7 1 2 77849 85277
0 8336 5 1 1 8335
0 8337 7 1 2 8334 8336
0 8338 5 1 1 8337
0 8339 7 1 2 81486 8338
0 8340 5 1 1 8339
0 8341 7 2 2 72265 76421
0 8342 5 2 1 88086
0 8343 7 19 2 64661 70266
0 8344 7 1 2 88090 83240
0 8345 7 1 2 88087 8344
0 8346 5 1 1 8345
0 8347 7 1 2 8340 8346
0 8348 5 1 1 8347
0 8349 7 1 2 68578 8348
0 8350 5 1 1 8349
0 8351 7 1 2 70631 6932
0 8352 5 3 1 8351
0 8353 7 2 2 70869 85332
0 8354 7 1 2 2296 88112
0 8355 5 1 1 8354
0 8356 7 1 2 88109 8355
0 8357 5 1 1 8356
0 8358 7 19 2 64662 65352
0 8359 7 2 2 83555 88114
0 8360 7 1 2 80435 88133
0 8361 7 1 2 8357 8360
0 8362 5 1 1 8361
0 8363 7 1 2 8350 8362
0 8364 5 1 1 8363
0 8365 7 1 2 78592 8364
0 8366 5 1 1 8365
0 8367 7 1 2 8332 8366
0 8368 5 1 1 8367
0 8369 7 1 2 66886 8368
0 8370 5 1 1 8369
0 8371 7 7 2 71295 72114
0 8372 7 8 2 69724 76692
0 8373 7 1 2 74782 88142
0 8374 7 1 2 88135 8373
0 8375 5 1 1 8374
0 8376 7 2 2 84601 74963
0 8377 7 1 2 76460 74980
0 8378 7 1 2 88150 8377
0 8379 5 1 1 8378
0 8380 7 1 2 8375 8379
0 8381 5 1 1 8380
0 8382 7 1 2 65079 8381
0 8383 5 1 1 8382
0 8384 7 3 2 74263 77761
0 8385 7 1 2 79507 87283
0 8386 7 1 2 88152 8385
0 8387 5 1 1 8386
0 8388 7 1 2 8383 8387
0 8389 5 1 1 8388
0 8390 7 1 2 84089 8389
0 8391 5 1 1 8390
0 8392 7 2 2 69509 74613
0 8393 7 1 2 74287 84063
0 8394 7 1 2 88155 8393
0 8395 7 1 2 87912 8394
0 8396 5 1 1 8395
0 8397 7 1 2 8391 8396
0 8398 5 1 1 8397
0 8399 7 1 2 62019 8398
0 8400 5 1 1 8399
0 8401 7 1 2 84310 86555
0 8402 5 1 1 8401
0 8403 7 2 2 77164 79426
0 8404 7 1 2 88157 88151
0 8405 7 1 2 8402 8404
0 8406 5 1 1 8405
0 8407 7 4 2 74614 86133
0 8408 7 1 2 73823 80112
0 8409 7 1 2 88159 8408
0 8410 5 1 1 8409
0 8411 7 1 2 8406 8410
0 8412 5 1 1 8411
0 8413 7 1 2 82964 8412
0 8414 5 1 1 8413
0 8415 7 1 2 8400 8414
0 8416 7 1 2 8370 8415
0 8417 5 1 1 8416
0 8418 7 1 2 87713 8417
0 8419 5 1 1 8418
0 8420 7 1 2 8288 8419
0 8421 7 1 2 8236 8420
0 8422 5 1 1 8421
0 8423 7 1 2 87699 8422
0 8424 5 1 1 8423
0 8425 7 1 2 7847 8424
0 8426 7 1 2 4747 8425
0 8427 5 1 1 8426
0 8428 7 10 2 61342 62939
0 8429 7 8 2 62994 88163
0 8430 7 1 2 8427 88173
0 8431 5 1 1 8430
0 8432 7 19 2 69510 76120
0 8433 5 1 1 88181
0 8434 7 5 2 65080 83032
0 8435 7 1 2 62334 75196
0 8436 7 1 2 88200 8435
0 8437 5 1 1 8436
0 8438 7 2 2 72818 83083
0 8439 7 1 2 76914 71660
0 8440 7 1 2 88205 8439
0 8441 5 1 1 8440
0 8442 7 1 2 8437 8441
0 8443 5 1 1 8442
0 8444 7 1 2 88182 8443
0 8445 5 1 1 8444
0 8446 7 2 2 77224 79663
0 8447 7 1 2 78981 82129
0 8448 7 1 2 88207 8447
0 8449 5 1 1 8448
0 8450 7 1 2 8445 8449
0 8451 5 1 1 8450
0 8452 7 1 2 63496 8451
0 8453 5 1 1 8452
0 8454 7 1 2 83084 81232
0 8455 5 1 1 8454
0 8456 7 7 2 68579 82875
0 8457 7 2 2 61766 79598
0 8458 7 1 2 88209 88216
0 8459 5 1 1 8458
0 8460 7 1 2 8455 8459
0 8461 5 1 1 8460
0 8462 7 1 2 61467 8461
0 8463 5 1 1 8462
0 8464 7 10 2 76814 87635
0 8465 7 2 2 70267 88218
0 8466 7 1 2 85139 88228
0 8467 5 1 1 8466
0 8468 7 1 2 8463 8467
0 8469 5 1 1 8468
0 8470 7 1 2 64663 8469
0 8471 5 1 1 8470
0 8472 7 7 2 70268 81907
0 8473 5 1 1 88230
0 8474 7 2 2 83085 86813
0 8475 5 1 1 88237
0 8476 7 1 2 88231 88238
0 8477 5 1 1 8476
0 8478 7 1 2 8471 8477
0 8479 5 1 1 8478
0 8480 7 1 2 77024 8479
0 8481 5 1 1 8480
0 8482 7 1 2 78232 81908
0 8483 5 1 1 8482
0 8484 7 18 2 64664 65945
0 8485 7 1 2 87175 88239
0 8486 7 1 2 77069 8485
0 8487 5 1 1 8486
0 8488 7 1 2 8483 8487
0 8489 5 1 1 8488
0 8490 7 1 2 76244 8489
0 8491 5 1 1 8490
0 8492 7 1 2 79011 81909
0 8493 5 1 1 8492
0 8494 7 1 2 8491 8493
0 8495 5 1 1 8494
0 8496 7 6 2 63497 83086
0 8497 7 1 2 8495 88257
0 8498 5 1 1 8497
0 8499 7 1 2 63088 8498
0 8500 7 1 2 8481 8499
0 8501 5 1 1 8500
0 8502 7 2 2 76881 77898
0 8503 5 1 1 88263
0 8504 7 1 2 79020 8503
0 8505 5 1 1 8504
0 8506 7 1 2 83087 8505
0 8507 5 1 1 8506
0 8508 7 3 2 61767 84710
0 8509 7 1 2 88265 79565
0 8510 5 1 1 8509
0 8511 7 1 2 8507 8510
0 8512 5 1 1 8511
0 8513 7 1 2 69511 8512
0 8514 5 1 1 8513
0 8515 7 2 2 77126 88091
0 8516 7 1 2 72027 88268
0 8517 7 1 2 85317 8516
0 8518 5 1 1 8517
0 8519 7 1 2 8514 8518
0 8520 5 1 1 8519
0 8521 7 1 2 63498 8520
0 8522 5 1 1 8521
0 8523 7 7 2 68099 87059
0 8524 7 6 2 61768 63726
0 8525 7 6 2 62335 64079
0 8526 7 1 2 88277 88283
0 8527 7 1 2 80496 8526
0 8528 7 1 2 88270 8527
0 8529 5 1 1 8528
0 8530 7 1 2 8522 8529
0 8531 5 1 1 8530
0 8532 7 1 2 61468 8531
0 8533 5 1 1 8532
0 8534 7 2 2 77183 85120
0 8535 7 13 2 63727 69512
0 8536 7 1 2 78059 88291
0 8537 7 1 2 88289 8536
0 8538 7 1 2 85146 8537
0 8539 5 1 1 8538
0 8540 7 1 2 67957 8539
0 8541 7 1 2 8533 8540
0 8542 5 1 1 8541
0 8543 7 1 2 62777 8542
0 8544 7 1 2 8501 8543
0 8545 5 1 1 8544
0 8546 7 1 2 8453 8545
0 8547 5 1 1 8546
0 8548 7 1 2 62020 8547
0 8549 5 1 1 8548
0 8550 7 1 2 78861 82954
0 8551 5 1 1 8550
0 8552 7 3 2 61769 81043
0 8553 5 2 1 88304
0 8554 7 1 2 78910 88305
0 8555 5 1 1 8554
0 8556 7 1 2 8551 8555
0 8557 5 1 1 8556
0 8558 7 1 2 61469 8557
0 8559 5 1 1 8558
0 8560 7 2 2 68336 87060
0 8561 7 1 2 83194 88309
0 8562 5 1 1 8561
0 8563 7 1 2 8559 8562
0 8564 5 2 1 8563
0 8565 7 1 2 76798 88311
0 8566 5 1 1 8565
0 8567 7 2 2 79012 87352
0 8568 5 1 1 88313
0 8569 7 1 2 80408 85263
0 8570 7 1 2 88314 8569
0 8571 5 1 1 8570
0 8572 7 1 2 8566 8571
0 8573 5 1 1 8572
0 8574 7 1 2 87555 80529
0 8575 7 1 2 8573 8574
0 8576 5 1 1 8575
0 8577 7 1 2 8549 8576
0 8578 5 1 1 8577
0 8579 7 1 2 64461 8578
0 8580 5 1 1 8579
0 8581 7 4 2 65353 84378
0 8582 7 2 2 70632 88315
0 8583 7 4 2 69958 74306
0 8584 7 2 2 81365 80800
0 8585 7 1 2 66386 88325
0 8586 7 1 2 88321 8585
0 8587 7 1 2 88319 8586
0 8588 5 1 1 8587
0 8589 7 1 2 72266 79716
0 8590 5 1 1 8589
0 8591 7 1 2 77830 86626
0 8592 5 1 1 8591
0 8593 7 1 2 8590 8592
0 8594 5 1 1 8593
0 8595 7 1 2 64665 83017
0 8596 7 1 2 8594 8595
0 8597 5 1 1 8596
0 8598 7 1 2 8588 8597
0 8599 5 1 1 8598
0 8600 7 1 2 79797 8599
0 8601 5 1 1 8600
0 8602 7 1 2 69725 8601
0 8603 7 1 2 8580 8602
0 8604 5 1 1 8603
0 8605 7 3 2 65694 85208
0 8606 7 1 2 88327 82689
0 8607 5 1 1 8606
0 8608 7 4 2 69513 81803
0 8609 7 4 2 66387 68580
0 8610 7 2 2 88334 85721
0 8611 7 1 2 88338 79307
0 8612 7 1 2 88330 8611
0 8613 5 1 1 8612
0 8614 7 1 2 8607 8613
0 8615 5 1 1 8614
0 8616 7 1 2 72115 8615
0 8617 5 1 1 8616
0 8618 7 1 2 82106 77165
0 8619 7 1 2 71151 8618
0 8620 5 1 1 8619
0 8621 7 2 2 70870 84883
0 8622 7 2 2 62336 83827
0 8623 7 1 2 88340 88342
0 8624 5 1 1 8623
0 8625 7 1 2 8620 8624
0 8626 5 1 1 8625
0 8627 7 1 2 68581 8626
0 8628 5 1 1 8627
0 8629 7 1 2 77488 75343
0 8630 5 1 1 8629
0 8631 7 1 2 72526 77850
0 8632 5 2 1 8631
0 8633 7 1 2 8630 88344
0 8634 5 1 1 8633
0 8635 7 1 2 63728 8634
0 8636 5 1 1 8635
0 8637 7 1 2 8636 81177
0 8638 5 1 1 8637
0 8639 7 1 2 81078 8638
0 8640 5 1 1 8639
0 8641 7 1 2 8628 8640
0 8642 5 1 1 8641
0 8643 7 1 2 64666 8642
0 8644 5 1 1 8643
0 8645 7 7 2 61470 64080
0 8646 7 2 2 80194 88346
0 8647 7 4 2 70633 72980
0 8648 7 2 2 70871 88355
0 8649 7 1 2 88353 88359
0 8650 5 1 1 8649
0 8651 7 2 2 63499 76121
0 8652 7 1 2 62778 76340
0 8653 5 1 1 8652
0 8654 7 1 2 75276 8653
0 8655 5 1 1 8654
0 8656 7 1 2 88361 8655
0 8657 5 1 1 8656
0 8658 7 1 2 8650 8657
0 8659 5 1 1 8658
0 8660 7 1 2 79343 8659
0 8661 5 1 1 8660
0 8662 7 1 2 8644 8661
0 8663 5 1 1 8662
0 8664 7 1 2 62021 8663
0 8665 5 1 1 8664
0 8666 7 2 2 62779 78911
0 8667 5 1 1 88363
0 8668 7 1 2 78900 8667
0 8669 5 7 1 8668
0 8670 7 1 2 68945 83771
0 8671 5 1 1 8670
0 8672 7 2 2 88365 8671
0 8673 7 3 2 61471 70634
0 8674 7 8 2 64462 70872
0 8675 7 1 2 88374 88377
0 8676 7 1 2 75378 8675
0 8677 7 1 2 88372 8676
0 8678 5 1 1 8677
0 8679 7 1 2 8665 8678
0 8680 5 1 1 8679
0 8681 7 1 2 69959 8680
0 8682 5 1 1 8681
0 8683 7 1 2 69514 76101
0 8684 5 3 1 8683
0 8685 7 1 2 77268 7172
0 8686 5 1 1 8685
0 8687 7 3 2 88385 8686
0 8688 7 2 2 65946 88388
0 8689 7 3 2 65695 71810
0 8690 7 1 2 82679 74600
0 8691 7 1 2 88393 8690
0 8692 7 1 2 88391 8691
0 8693 5 1 1 8692
0 8694 7 1 2 8682 8693
0 8695 5 1 1 8694
0 8696 7 1 2 63263 8695
0 8697 5 1 1 8696
0 8698 7 1 2 8617 8697
0 8699 5 1 1 8698
0 8700 7 1 2 65354 8699
0 8701 5 1 1 8700
0 8702 7 3 2 74106 76461
0 8703 7 2 2 65081 78862
0 8704 7 1 2 88396 88399
0 8705 5 1 1 8704
0 8706 7 3 2 67172 80195
0 8707 7 2 2 80183 78233
0 8708 7 1 2 88401 88404
0 8709 5 1 1 8708
0 8710 7 1 2 8705 8709
0 8711 5 1 1 8710
0 8712 7 1 2 61472 8711
0 8713 5 1 1 8712
0 8714 7 1 2 76069 79220
0 8715 7 1 2 88405 8714
0 8716 5 1 1 8715
0 8717 7 1 2 8713 8716
0 8718 5 1 1 8717
0 8719 7 1 2 62022 8718
0 8720 5 1 1 8719
0 8721 7 2 2 77225 76815
0 8722 7 3 2 63729 79745
0 8723 7 1 2 74107 88408
0 8724 7 1 2 88406 8723
0 8725 5 1 1 8724
0 8726 7 1 2 8720 8725
0 8727 5 1 1 8726
0 8728 7 1 2 81692 80497
0 8729 7 1 2 8727 8728
0 8730 5 1 1 8729
0 8731 7 1 2 8701 8730
0 8732 5 1 1 8731
0 8733 7 1 2 61770 8732
0 8734 5 1 1 8733
0 8735 7 5 2 62780 75470
0 8736 7 1 2 76921 79021
0 8737 5 11 1 8736
0 8738 7 2 2 63500 88416
0 8739 5 1 1 88427
0 8740 7 2 2 80965 85887
0 8741 7 1 2 88428 88429
0 8742 5 1 1 8741
0 8743 7 1 2 69960 75927
0 8744 5 1 1 8743
0 8745 7 2 2 76980 8744
0 8746 5 1 1 88431
0 8747 7 1 2 74176 8746
0 8748 5 1 1 8747
0 8749 7 1 2 80703 74197
0 8750 5 2 1 8749
0 8751 7 1 2 8748 88433
0 8752 5 1 1 8751
0 8753 7 1 2 83828 8752
0 8754 5 1 1 8753
0 8755 7 1 2 8742 8754
0 8756 5 1 1 8755
0 8757 7 1 2 68100 8756
0 8758 5 1 1 8757
0 8759 7 2 2 71811 76122
0 8760 7 4 2 64463 70635
0 8761 7 2 2 70873 88437
0 8762 7 4 2 79599 81609
0 8763 7 1 2 88441 88443
0 8764 7 1 2 88435 8763
0 8765 5 1 1 8764
0 8766 7 1 2 8758 8765
0 8767 5 1 1 8766
0 8768 7 1 2 69515 8767
0 8769 5 1 1 8768
0 8770 7 1 2 81116 3608
0 8771 5 1 1 8770
0 8772 7 6 2 70636 79600
0 8773 7 1 2 88447 78803
0 8774 7 1 2 88219 8773
0 8775 7 1 2 8771 8774
0 8776 5 1 1 8775
0 8777 7 1 2 8769 8776
0 8778 5 1 1 8777
0 8779 7 1 2 64081 8778
0 8780 5 1 1 8779
0 8781 7 2 2 83829 81366
0 8782 7 1 2 77077 88453
0 8783 5 1 1 8782
0 8784 7 1 2 8780 8783
0 8785 5 1 1 8784
0 8786 7 1 2 88411 8785
0 8787 5 1 1 8786
0 8788 7 1 2 64881 8787
0 8789 7 1 2 8734 8788
0 8790 5 1 1 8789
0 8791 7 1 2 69164 8790
0 8792 7 1 2 8604 8791
0 8793 5 1 1 8792
0 8794 7 3 2 76758 86669
0 8795 7 15 2 64318 69516
0 8796 7 1 2 88458 86300
0 8797 7 1 2 88455 8796
0 8798 7 1 2 87653 8797
0 8799 7 1 2 87668 8798
0 8800 5 1 1 8799
0 8801 7 1 2 8793 8800
0 8802 5 1 1 8801
0 8803 7 1 2 71296 8802
0 8804 5 1 1 8803
0 8805 7 2 2 62781 80869
0 8806 7 3 2 61473 82149
0 8807 7 1 2 88473 88475
0 8808 5 1 1 8807
0 8809 7 2 2 71812 77184
0 8810 7 1 2 77293 88478
0 8811 5 1 1 8810
0 8812 7 1 2 8808 8811
0 8813 5 1 1 8812
0 8814 7 3 2 63264 75848
0 8815 7 1 2 8813 88480
0 8816 5 1 1 8815
0 8817 7 1 2 5891 77309
0 8818 5 2 1 8817
0 8819 7 1 2 62023 88483
0 8820 5 1 1 8819
0 8821 7 2 2 76816 75070
0 8822 5 1 1 88485
0 8823 7 1 2 8820 8822
0 8824 5 1 1 8823
0 8825 7 1 2 62517 8824
0 8826 5 1 1 8825
0 8827 7 2 2 63730 75759
0 8828 5 1 1 88487
0 8829 7 1 2 8826 8828
0 8830 5 1 1 8829
0 8831 7 1 2 77185 8830
0 8832 5 1 1 8831
0 8833 7 7 2 71297 72981
0 8834 5 4 1 88489
0 8835 7 17 2 68582 82406
0 8836 5 2 1 88500
0 8837 7 1 2 71910 88517
0 8838 7 2 2 88496 8837
0 8839 7 4 2 66887 78493
0 8840 7 1 2 88519 88521
0 8841 5 1 1 8840
0 8842 7 1 2 63265 8841
0 8843 7 1 2 8832 8842
0 8844 5 1 1 8843
0 8845 7 1 2 83283 87914
0 8846 5 1 1 8845
0 8847 7 1 2 68101 8846
0 8848 5 1 1 8847
0 8849 7 1 2 69961 8848
0 8850 7 1 2 8844 8849
0 8851 5 1 1 8850
0 8852 7 1 2 8816 8851
0 8853 5 1 1 8852
0 8854 7 1 2 64464 8853
0 8855 5 1 1 8854
0 8856 7 2 2 79897 84616
0 8857 7 13 2 71911 88525
0 8858 7 4 2 65082 88527
0 8859 7 3 2 69318 81548
0 8860 7 2 2 88540 88544
0 8861 7 5 2 67628 82613
0 8862 7 1 2 66388 88549
0 8863 7 1 2 88547 8862
0 8864 5 1 1 8863
0 8865 7 1 2 8855 8864
0 8866 5 1 1 8865
0 8867 7 1 2 69517 8866
0 8868 5 1 1 8867
0 8869 7 4 2 61474 76759
0 8870 7 5 2 62518 63266
0 8871 7 1 2 82351 88558
0 8872 7 1 2 88554 8871
0 8873 5 1 1 8872
0 8874 7 1 2 88339 74950
0 8875 7 1 2 83088 8874
0 8876 5 1 1 8875
0 8877 7 1 2 8873 8876
0 8878 5 1 1 8877
0 8879 7 1 2 63501 8878
0 8880 5 1 1 8879
0 8881 7 1 2 79798 80923
0 8882 7 1 2 72982 8881
0 8883 7 1 2 84823 8882
0 8884 5 1 1 8883
0 8885 7 1 2 8880 8884
0 8886 5 1 1 8885
0 8887 7 1 2 69962 8886
0 8888 5 1 1 8887
0 8889 7 2 2 77186 75190
0 8890 5 1 1 88563
0 8891 7 1 2 82614 80623
0 8892 7 1 2 88528 8891
0 8893 5 1 1 8892
0 8894 7 1 2 8890 8893
0 8895 5 1 1 8894
0 8896 7 1 2 81323 87461
0 8897 7 1 2 8895 8896
0 8898 5 1 1 8897
0 8899 7 1 2 8888 8898
0 8900 5 1 1 8899
0 8901 7 1 2 64667 8900
0 8902 5 1 1 8901
0 8903 7 1 2 63089 8902
0 8904 7 1 2 8868 8903
0 8905 5 1 1 8904
0 8906 7 4 2 66888 80905
0 8907 7 2 2 88541 88565
0 8908 5 1 1 88569
0 8909 7 1 2 73295 81124
0 8910 7 1 2 85201 8909
0 8911 5 1 1 8910
0 8912 7 1 2 8908 8911
0 8913 5 1 1 8912
0 8914 7 1 2 68102 8913
0 8915 5 1 1 8914
0 8916 7 2 2 84780 88520
0 8917 5 1 1 88571
0 8918 7 1 2 83577 88572
0 8919 5 1 1 8918
0 8920 7 1 2 8915 8919
0 8921 5 1 1 8920
0 8922 7 1 2 66650 8921
0 8923 5 1 1 8922
0 8924 7 4 2 64668 83033
0 8925 7 1 2 75085 79668
0 8926 5 1 1 8925
0 8927 7 1 2 79002 75105
0 8928 5 2 1 8927
0 8929 7 1 2 8926 88577
0 8930 5 1 1 8929
0 8931 7 1 2 88573 8930
0 8932 5 1 1 8931
0 8933 7 1 2 8923 8932
0 8934 5 1 1 8933
0 8935 7 1 2 61475 8934
0 8936 5 1 1 8935
0 8937 7 3 2 69963 85414
0 8938 7 2 2 69518 82615
0 8939 7 1 2 82261 88582
0 8940 5 1 1 8939
0 8941 7 2 2 63502 81889
0 8942 7 1 2 74150 88584
0 8943 5 1 1 8942
0 8944 7 1 2 8940 8943
0 8945 5 1 1 8944
0 8946 7 1 2 88579 8945
0 8947 5 1 1 8946
0 8948 7 1 2 8936 8947
0 8949 5 1 1 8948
0 8950 7 1 2 84224 8949
0 8951 5 1 1 8950
0 8952 7 6 2 61476 63503
0 8953 7 2 2 88278 88586
0 8954 7 1 2 88592 84523
0 8955 7 1 2 81567 8954
0 8956 5 1 1 8955
0 8957 7 1 2 67958 8956
0 8958 7 1 2 8951 8957
0 8959 5 1 1 8958
0 8960 7 1 2 65947 8959
0 8961 7 1 2 8905 8960
0 8962 5 1 1 8961
0 8963 7 2 2 63267 81890
0 8964 7 1 2 85049 88594
0 8965 5 1 1 8964
0 8966 7 3 2 88271 74783
0 8967 5 1 1 88596
0 8968 7 1 2 73397 88597
0 8969 5 1 1 8968
0 8970 7 1 2 8965 8969
0 8971 5 1 1 8970
0 8972 7 1 2 68337 8971
0 8973 5 1 1 8972
0 8974 7 2 2 83578 84815
0 8975 7 1 2 82208 88599
0 8976 5 1 1 8975
0 8977 7 1 2 8973 8976
0 8978 5 1 1 8977
0 8979 7 2 2 82107 82616
0 8980 7 1 2 8978 88601
0 8981 5 1 1 8980
0 8982 7 2 2 86864 88501
0 8983 7 4 2 65083 73398
0 8984 7 2 2 66889 88605
0 8985 7 1 2 78982 88609
0 8986 7 1 2 88603 8985
0 8987 5 1 1 8986
0 8988 7 1 2 82255 88583
0 8989 5 1 1 8988
0 8990 7 2 2 61771 77435
0 8991 7 1 2 88585 88611
0 8992 5 1 1 8991
0 8993 7 1 2 8989 8992
0 8994 5 1 1 8993
0 8995 7 1 2 79527 87195
0 8996 7 1 2 8994 8995
0 8997 5 1 1 8996
0 8998 7 1 2 8987 8997
0 8999 5 1 1 8998
0 9000 7 1 2 61477 8999
0 9001 5 1 1 9000
0 9002 7 2 2 88292 79528
0 9003 7 1 2 80780 74307
0 9004 7 1 2 88613 9003
0 9005 5 1 1 9004
0 9006 7 4 2 67173 72913
0 9007 5 1 1 88615
0 9008 7 9 2 66389 68790
0 9009 7 1 2 73803 88619
0 9010 7 1 2 88616 9009
0 9011 7 1 2 79464 9010
0 9012 5 1 1 9011
0 9013 7 1 2 9005 9012
0 9014 5 1 1 9013
0 9015 7 1 2 83089 9014
0 9016 5 1 1 9015
0 9017 7 1 2 9001 9016
0 9018 7 1 2 8981 9017
0 9019 5 1 1 9018
0 9020 7 1 2 63090 9019
0 9021 5 1 1 9020
0 9022 7 2 2 78060 85415
0 9023 5 1 1 88628
0 9024 7 1 2 61478 83008
0 9025 5 1 1 9024
0 9026 7 1 2 9023 9025
0 9027 5 4 1 9026
0 9028 7 1 2 81399 88630
0 9029 5 1 1 9028
0 9030 7 9 2 61479 68791
0 9031 7 1 2 88634 82554
0 9032 5 1 1 9031
0 9033 7 1 2 9029 9032
0 9034 5 1 1 9033
0 9035 7 1 2 74784 9034
0 9036 5 1 1 9035
0 9037 7 3 2 61480 83579
0 9038 7 1 2 82574 74024
0 9039 7 1 2 88643 9038
0 9040 5 1 1 9039
0 9041 7 1 2 9036 9040
0 9042 5 1 1 9041
0 9043 7 1 2 85722 81646
0 9044 7 1 2 9042 9043
0 9045 5 1 1 9044
0 9046 7 1 2 64882 9045
0 9047 7 1 2 9021 9046
0 9048 7 1 2 8962 9047
0 9049 5 1 1 9048
0 9050 7 1 2 73908 9007
0 9051 5 1 1 9050
0 9052 7 5 2 65084 82366
0 9053 7 2 2 9051 88646
0 9054 7 1 2 74860 88651
0 9055 5 1 1 9054
0 9056 7 1 2 77070 73296
0 9057 5 1 1 9056
0 9058 7 1 2 78154 9057
0 9059 5 1 1 9058
0 9060 7 1 2 88258 9059
0 9061 5 1 1 9060
0 9062 7 4 2 61772 84856
0 9063 7 2 2 69964 73909
0 9064 5 1 1 88657
0 9065 7 1 2 88653 88658
0 9066 5 1 1 9065
0 9067 7 1 2 9061 9066
0 9068 5 1 1 9067
0 9069 7 1 2 67629 9068
0 9070 5 1 1 9069
0 9071 7 1 2 9055 9070
0 9072 5 1 1 9071
0 9073 7 1 2 62024 9072
0 9074 5 1 1 9073
0 9075 7 2 2 63268 75400
0 9076 7 1 2 74914 81024
0 9077 5 1 1 9076
0 9078 7 1 2 65085 74264
0 9079 5 1 1 9078
0 9080 7 1 2 9077 9079
0 9081 5 1 1 9080
0 9082 7 1 2 88659 9081
0 9083 5 1 1 9082
0 9084 7 1 2 9074 9083
0 9085 5 1 1 9084
0 9086 7 1 2 65948 9085
0 9087 5 1 1 9086
0 9088 7 2 2 78144 83405
0 9089 7 1 2 87085 88661
0 9090 5 1 1 9089
0 9091 7 1 2 9087 9090
0 9092 5 1 1 9091
0 9093 7 1 2 83791 9092
0 9094 5 1 1 9093
0 9095 7 16 2 62025 68103
0 9096 7 1 2 68338 84706
0 9097 5 1 1 9096
0 9098 7 1 2 88663 9097
0 9099 5 1 1 9098
0 9100 7 1 2 9099 85109
0 9101 5 1 1 9100
0 9102 7 1 2 78145 9101
0 9103 5 1 1 9102
0 9104 7 4 2 65086 73563
0 9105 7 1 2 82130 88679
0 9106 7 1 2 77513 9105
0 9107 5 1 1 9106
0 9108 7 1 2 9103 9107
0 9109 5 1 1 9108
0 9110 7 1 2 83792 9109
0 9111 5 1 1 9110
0 9112 7 8 2 68583 69319
0 9113 7 3 2 68339 88683
0 9114 7 6 2 67630 81804
0 9115 7 2 2 88691 88694
0 9116 7 1 2 78651 78035
0 9117 7 1 2 88700 9116
0 9118 5 1 1 9117
0 9119 7 1 2 9111 9118
0 9120 5 1 1 9119
0 9121 7 1 2 61773 9120
0 9122 5 1 1 9121
0 9123 7 5 2 69320 81805
0 9124 7 1 2 78122 77047
0 9125 5 4 1 9124
0 9126 7 1 2 73539 70988
0 9127 7 1 2 88707 9126
0 9128 5 1 1 9127
0 9129 7 1 2 65087 75495
0 9130 5 1 1 9129
0 9131 7 1 2 9128 9130
0 9132 5 1 1 9131
0 9133 7 1 2 88702 9132
0 9134 5 1 1 9133
0 9135 7 6 2 69965 75133
0 9136 7 5 2 83793 82367
0 9137 7 1 2 88711 88717
0 9138 5 1 1 9137
0 9139 7 1 2 9134 9138
0 9140 5 1 1 9139
0 9141 7 1 2 68584 9140
0 9142 5 1 1 9141
0 9143 7 4 2 81806 74308
0 9144 7 1 2 85888 88722
0 9145 5 1 1 9144
0 9146 7 2 2 82352 83565
0 9147 5 1 1 88726
0 9148 7 1 2 9145 9147
0 9149 5 1 1 9148
0 9150 7 1 2 67631 9149
0 9151 5 1 1 9150
0 9152 7 11 2 64465 65949
0 9153 7 2 2 87654 88728
0 9154 5 1 1 88739
0 9155 7 1 2 9151 9154
0 9156 5 1 1 9155
0 9157 7 1 2 65088 85911
0 9158 7 1 2 9156 9157
0 9159 5 1 1 9158
0 9160 7 1 2 9142 9159
0 9161 5 1 1 9160
0 9162 7 1 2 67174 9161
0 9163 5 1 1 9162
0 9164 7 1 2 75794 84707
0 9165 5 1 1 9164
0 9166 7 1 2 78146 83794
0 9167 7 1 2 74351 81438
0 9168 7 1 2 9166 9167
0 9169 7 1 2 9165 9168
0 9170 5 1 1 9169
0 9171 7 1 2 9163 9170
0 9172 7 1 2 9122 9171
0 9173 5 1 1 9172
0 9174 7 1 2 68792 9173
0 9175 5 1 1 9174
0 9176 7 2 2 61774 85760
0 9177 7 2 2 67175 88684
0 9178 7 5 2 68340 81807
0 9179 7 1 2 78821 88745
0 9180 7 1 2 88743 9179
0 9181 7 1 2 88741 9180
0 9182 5 1 1 9181
0 9183 7 1 2 9175 9182
0 9184 7 1 2 9094 9183
0 9185 5 1 1 9184
0 9186 7 1 2 66390 9185
0 9187 5 1 1 9186
0 9188 7 3 2 62519 74428
0 9189 5 1 1 88750
0 9190 7 8 2 63913 69966
0 9191 7 2 2 65950 88753
0 9192 7 1 2 88751 88761
0 9193 5 1 1 9192
0 9194 7 1 2 62782 80690
0 9195 5 1 1 9194
0 9196 7 1 2 77310 9195
0 9197 5 1 1 9196
0 9198 7 1 2 77436 9197
0 9199 5 1 1 9198
0 9200 7 1 2 78089 9199
0 9201 5 1 1 9200
0 9202 7 1 2 63731 85735
0 9203 7 1 2 9201 9202
0 9204 5 1 1 9203
0 9205 7 1 2 9193 9204
0 9206 5 1 1 9205
0 9207 7 1 2 83090 9206
0 9208 5 1 1 9207
0 9209 7 1 2 84809 88652
0 9210 5 1 1 9209
0 9211 7 1 2 9208 9210
0 9212 5 1 1 9211
0 9213 7 1 2 62026 9212
0 9214 5 1 1 9213
0 9215 7 1 2 66890 80518
0 9216 5 1 1 9215
0 9217 7 1 2 82258 9216
0 9218 5 1 1 9217
0 9219 7 1 2 81610 73564
0 9220 7 1 2 76290 9219
0 9221 7 1 2 9218 9220
0 9222 5 1 1 9221
0 9223 7 1 2 9214 9222
0 9224 5 1 1 9223
0 9225 7 1 2 67959 9224
0 9226 5 1 1 9225
0 9227 7 11 2 61775 63091
0 9228 7 1 2 73565 88763
0 9229 7 1 2 84251 9228
0 9230 7 1 2 88542 9229
0 9231 5 1 1 9230
0 9232 7 1 2 9226 9231
0 9233 5 1 1 9232
0 9234 7 1 2 82838 9233
0 9235 5 1 1 9234
0 9236 7 1 2 69519 9235
0 9237 7 1 2 9187 9236
0 9238 5 1 1 9237
0 9239 7 5 2 80801 81549
0 9240 7 1 2 87462 88774
0 9241 5 1 1 9240
0 9242 7 3 2 64466 82653
0 9243 7 1 2 81025 88779
0 9244 7 1 2 85812 9243
0 9245 5 1 1 9244
0 9246 7 1 2 9241 9245
0 9247 5 1 1 9246
0 9248 7 1 2 85240 9247
0 9249 5 1 1 9248
0 9250 7 1 2 62337 84968
0 9251 5 1 1 9250
0 9252 7 1 2 74046 9251
0 9253 5 1 1 9252
0 9254 7 5 2 67632 82654
0 9255 7 1 2 79529 88782
0 9256 7 1 2 9253 9255
0 9257 5 1 1 9256
0 9258 7 1 2 9249 9257
0 9259 5 1 1 9258
0 9260 7 1 2 61481 9259
0 9261 5 1 1 9260
0 9262 7 1 2 83435 88606
0 9263 5 1 1 9262
0 9264 7 4 2 67960 81611
0 9265 7 1 2 80691 88787
0 9266 5 1 1 9265
0 9267 7 1 2 9263 9266
0 9268 5 1 1 9267
0 9269 7 1 2 82108 74785
0 9270 7 1 2 9268 9269
0 9271 5 1 1 9270
0 9272 7 1 2 9261 9271
0 9273 5 1 1 9272
0 9274 7 1 2 66891 9273
0 9275 5 1 1 9274
0 9276 7 3 2 68104 75849
0 9277 7 1 2 88484 88791
0 9278 5 1 1 9277
0 9279 7 1 2 8917 9278
0 9280 5 1 1 9279
0 9281 7 1 2 69967 9280
0 9282 5 1 1 9281
0 9283 7 1 2 84857 88474
0 9284 5 1 1 9283
0 9285 7 7 2 62338 82264
0 9286 7 1 2 77294 88794
0 9287 5 1 1 9286
0 9288 7 1 2 9284 9287
0 9289 5 1 1 9288
0 9290 7 1 2 75850 9289
0 9291 5 1 1 9290
0 9292 7 1 2 9282 9291
0 9293 5 1 1 9292
0 9294 7 1 2 83795 9293
0 9295 5 1 1 9294
0 9296 7 1 2 81717 88548
0 9297 5 1 1 9296
0 9298 7 1 2 9295 9297
0 9299 5 1 1 9298
0 9300 7 1 2 61482 9299
0 9301 5 1 1 9300
0 9302 7 1 2 82088 82262
0 9303 5 1 1 9302
0 9304 7 1 2 88543 83436
0 9305 5 1 1 9304
0 9306 7 1 2 9303 9305
0 9307 5 1 1 9306
0 9308 7 2 2 85723 80924
0 9309 7 1 2 9307 88801
0 9310 5 1 1 9309
0 9311 7 1 2 9301 9310
0 9312 5 1 1 9311
0 9313 7 1 2 65951 9312
0 9314 5 1 1 9313
0 9315 7 1 2 9275 9314
0 9316 5 1 1 9315
0 9317 7 1 2 61776 9316
0 9318 5 1 1 9317
0 9319 7 2 2 69968 88587
0 9320 7 4 2 80802 86865
0 9321 7 1 2 77584 88805
0 9322 5 1 1 9321
0 9323 7 3 2 65952 73297
0 9324 5 1 1 88809
0 9325 7 1 2 82687 88810
0 9326 5 1 1 9325
0 9327 7 1 2 9322 9326
0 9328 5 1 1 9327
0 9329 7 1 2 88803 9328
0 9330 5 1 1 9329
0 9331 7 4 2 68105 76123
0 9332 7 9 2 65089 75134
0 9333 7 1 2 88812 88816
0 9334 5 1 1 9333
0 9335 7 1 2 74214 88629
0 9336 5 1 1 9335
0 9337 7 1 2 9334 9336
0 9338 5 1 1 9337
0 9339 7 1 2 81876 9338
0 9340 5 1 1 9339
0 9341 7 6 2 69969 75760
0 9342 5 2 1 88825
0 9343 7 1 2 77311 5983
0 9344 5 1 1 9343
0 9345 7 1 2 62027 9344
0 9346 5 1 1 9345
0 9347 7 3 2 62783 78061
0 9348 5 1 1 88833
0 9349 7 1 2 9346 9348
0 9350 5 1 1 9349
0 9351 7 1 2 77437 9350
0 9352 5 1 1 9351
0 9353 7 1 2 88831 9352
0 9354 5 1 1 9353
0 9355 7 4 2 77226 88729
0 9356 5 1 1 88836
0 9357 7 1 2 63269 88837
0 9358 7 1 2 9354 9357
0 9359 5 1 1 9358
0 9360 7 1 2 9340 9359
0 9361 5 1 1 9360
0 9362 7 1 2 63732 9361
0 9363 5 1 1 9362
0 9364 7 1 2 9330 9363
0 9365 5 1 1 9364
0 9366 7 1 2 66651 9365
0 9367 5 1 1 9366
0 9368 7 1 2 64669 9367
0 9369 7 1 2 9318 9368
0 9370 5 1 1 9369
0 9371 7 1 2 9238 9370
0 9372 5 1 1 9371
0 9373 7 1 2 69726 9372
0 9374 5 1 1 9373
0 9375 7 1 2 68946 9374
0 9376 7 1 2 9049 9375
0 9377 5 1 1 9376
0 9378 7 1 2 85774 85988
0 9379 5 1 1 9378
0 9380 7 1 2 9379 81885
0 9381 5 1 1 9380
0 9382 7 1 2 66652 9381
0 9383 5 1 1 9382
0 9384 7 1 2 71813 77590
0 9385 5 1 1 9384
0 9386 7 1 2 67176 79841
0 9387 5 1 1 9386
0 9388 7 1 2 9385 9387
0 9389 5 1 1 9388
0 9390 7 1 2 83328 9389
0 9391 5 1 1 9390
0 9392 7 1 2 9383 9391
0 9393 5 1 1 9392
0 9394 7 1 2 61483 9393
0 9395 5 1 1 9394
0 9396 7 1 2 77438 85980
0 9397 5 1 1 9396
0 9398 7 1 2 73566 82061
0 9399 5 1 1 9398
0 9400 7 1 2 9397 9399
0 9401 5 1 1 9400
0 9402 7 1 2 66391 82774
0 9403 7 1 2 9401 9402
0 9404 5 1 1 9403
0 9405 7 1 2 9395 9404
0 9406 5 1 1 9405
0 9407 7 1 2 63504 9406
0 9408 5 1 1 9407
0 9409 7 3 2 63733 77187
0 9410 7 1 2 81795 88840
0 9411 7 1 2 88011 9410
0 9412 5 1 1 9411
0 9413 7 1 2 9408 9412
0 9414 5 1 1 9413
0 9415 7 1 2 69970 9414
0 9416 5 1 1 9415
0 9417 7 2 2 75086 78593
0 9418 5 1 1 88843
0 9419 7 1 2 77188 88293
0 9420 7 1 2 88844 9419
0 9421 5 1 1 9420
0 9422 7 1 2 9416 9421
0 9423 5 1 1 9422
0 9424 7 1 2 63092 9423
0 9425 5 1 1 9424
0 9426 7 2 2 75401 74861
0 9427 5 1 1 88845
0 9428 7 1 2 87395 9427
0 9429 5 3 1 9428
0 9430 7 9 2 63093 64082
0 9431 7 2 2 88850 87398
0 9432 5 1 1 88859
0 9433 7 3 2 81338 80341
0 9434 7 1 2 88860 88861
0 9435 7 1 2 88847 9434
0 9436 5 1 1 9435
0 9437 7 2 2 75571 83580
0 9438 5 1 1 88864
0 9439 7 4 2 69520 77166
0 9440 7 1 2 65090 88866
0 9441 5 1 1 9440
0 9442 7 1 2 9438 9441
0 9443 5 1 1 9442
0 9444 7 1 2 81980 9443
0 9445 5 1 1 9444
0 9446 7 1 2 82030 83448
0 9447 5 1 1 9446
0 9448 7 1 2 9445 9447
0 9449 5 1 1 9448
0 9450 7 1 2 61484 9449
0 9451 5 1 1 9450
0 9452 7 10 2 66392 88764
0 9453 7 1 2 78594 80482
0 9454 7 1 2 88870 9453
0 9455 5 1 1 9454
0 9456 7 1 2 9451 9455
0 9457 5 1 1 9456
0 9458 7 2 2 65953 72983
0 9459 7 1 2 67633 88880
0 9460 7 1 2 9457 9459
0 9461 5 1 1 9460
0 9462 7 1 2 9436 9461
0 9463 5 1 1 9462
0 9464 7 1 2 67390 9463
0 9465 5 1 1 9464
0 9466 7 1 2 78912 88593
0 9467 7 1 2 78628 9466
0 9468 5 1 1 9467
0 9469 7 1 2 9465 9468
0 9470 7 1 2 9425 9469
0 9471 5 1 1 9470
0 9472 7 1 2 63270 9471
0 9473 5 1 1 9472
0 9474 7 2 2 63734 78540
0 9475 5 2 1 88882
0 9476 7 4 2 65954 72693
0 9477 5 3 1 88886
0 9478 7 1 2 74834 88890
0 9479 5 1 1 9478
0 9480 7 1 2 69727 77059
0 9481 7 1 2 9479 9480
0 9482 5 1 1 9481
0 9483 7 1 2 88884 9482
0 9484 5 1 1 9483
0 9485 7 1 2 68341 9484
0 9486 5 1 1 9485
0 9487 7 1 2 77406 82973
0 9488 5 1 1 9487
0 9489 7 1 2 9486 9488
0 9490 5 1 1 9489
0 9491 7 2 2 81749 81796
0 9492 7 1 2 83284 88893
0 9493 7 1 2 9490 9492
0 9494 5 1 1 9493
0 9495 7 1 2 9473 9494
0 9496 5 1 1 9495
0 9497 7 1 2 64467 9496
0 9498 5 1 1 9497
0 9499 7 9 2 62784 64468
0 9500 7 3 2 84121 88895
0 9501 7 1 2 80342 88904
0 9502 5 1 1 9501
0 9503 7 2 2 62520 81324
0 9504 7 1 2 83627 88907
0 9505 5 1 1 9504
0 9506 7 1 2 9502 9505
0 9507 5 1 1 9506
0 9508 7 1 2 61777 9507
0 9509 5 1 1 9508
0 9510 7 14 2 63271 69321
0 9511 7 1 2 88909 71666
0 9512 7 1 2 82019 9511
0 9513 5 1 1 9512
0 9514 7 1 2 9509 9513
0 9515 5 1 1 9514
0 9516 7 1 2 64083 9515
0 9517 5 1 1 9516
0 9518 7 3 2 81612 86134
0 9519 5 1 1 88923
0 9520 7 1 2 61778 88924
0 9521 5 1 1 9520
0 9522 7 1 2 9517 9521
0 9523 5 1 1 9522
0 9524 7 1 2 76124 9523
0 9525 5 1 1 9524
0 9526 7 2 2 64084 87556
0 9527 7 1 2 81079 79201
0 9528 5 1 1 9527
0 9529 7 1 2 80042 82597
0 9530 7 1 2 76551 78747
0 9531 7 1 2 9529 9530
0 9532 5 1 1 9531
0 9533 7 1 2 9528 9532
0 9534 5 1 1 9533
0 9535 7 1 2 88926 9534
0 9536 5 1 1 9535
0 9537 7 1 2 9525 9536
0 9538 5 1 1 9537
0 9539 7 1 2 65091 9538
0 9540 5 1 1 9539
0 9541 7 4 2 69728 73567
0 9542 7 1 2 85416 88928
0 9543 5 1 1 9542
0 9544 7 1 2 86809 9543
0 9545 5 1 1 9544
0 9546 7 5 2 64469 88765
0 9547 7 1 2 80915 88932
0 9548 7 1 2 9545 9547
0 9549 5 1 1 9548
0 9550 7 1 2 9540 9549
0 9551 5 1 1 9550
0 9552 7 1 2 74786 9551
0 9553 5 1 1 9552
0 9554 7 21 2 68106 69729
0 9555 5 1 1 88937
0 9556 7 1 2 71667 88938
0 9557 5 1 1 9556
0 9558 7 2 2 87557 76844
0 9559 5 1 1 88958
0 9560 7 1 2 9557 9559
0 9561 5 1 1 9560
0 9562 7 1 2 61779 9561
0 9563 5 1 1 9562
0 9564 7 1 2 63272 78637
0 9565 5 1 1 9564
0 9566 7 1 2 9563 9565
0 9567 5 1 1 9566
0 9568 7 1 2 83796 9567
0 9569 5 1 1 9568
0 9570 7 2 2 80196 70989
0 9571 7 1 2 81208 86866
0 9572 7 1 2 88960 9571
0 9573 5 1 1 9572
0 9574 7 1 2 9569 9573
0 9575 5 1 1 9574
0 9576 7 1 2 88284 9575
0 9577 5 1 1 9576
0 9578 7 19 2 63273 64883
0 9579 5 4 1 88962
0 9580 7 3 2 61780 88963
0 9581 5 1 1 88985
0 9582 7 1 2 83091 88929
0 9583 5 1 1 9582
0 9584 7 1 2 9581 9583
0 9585 5 1 1 9584
0 9586 7 1 2 64470 80409
0 9587 7 1 2 9585 9586
0 9588 5 1 1 9587
0 9589 7 1 2 66393 9588
0 9590 7 1 2 9577 9589
0 9591 5 1 1 9590
0 9592 7 2 2 63505 73568
0 9593 5 1 1 88988
0 9594 7 2 2 78023 77762
0 9595 5 1 1 88990
0 9596 7 1 2 9593 9595
0 9597 5 1 1 9596
0 9598 7 1 2 87303 9597
0 9599 5 1 1 9598
0 9600 7 3 2 81678 88964
0 9601 5 1 1 88992
0 9602 7 1 2 9599 9601
0 9603 5 1 1 9602
0 9604 7 9 2 67961 64471
0 9605 7 1 2 9603 88995
0 9606 5 1 1 9605
0 9607 7 1 2 61485 9606
0 9608 5 1 1 9607
0 9609 7 1 2 69971 9608
0 9610 7 1 2 9591 9609
0 9611 5 1 1 9610
0 9612 7 2 2 81693 83860
0 9613 7 1 2 87600 89004
0 9614 5 1 1 9613
0 9615 7 1 2 69521 9614
0 9616 7 1 2 9611 9615
0 9617 5 1 1 9616
0 9618 7 2 2 80026 84225
0 9619 7 1 2 78672 89006
0 9620 5 1 1 9619
0 9621 7 4 2 72028 77794
0 9622 5 1 1 89008
0 9623 7 1 2 79530 80505
0 9624 7 1 2 89009 9623
0 9625 5 1 1 9624
0 9626 7 1 2 9620 9625
0 9627 5 1 1 9626
0 9628 7 1 2 61781 9627
0 9629 5 1 1 9628
0 9630 7 4 2 69322 81647
0 9631 7 1 2 78541 88991
0 9632 5 1 1 9631
0 9633 7 1 2 67391 87601
0 9634 5 1 1 9633
0 9635 7 1 2 9632 9634
0 9636 5 1 1 9635
0 9637 7 1 2 89012 9636
0 9638 5 1 1 9637
0 9639 7 1 2 9629 9638
0 9640 5 1 1 9639
0 9641 7 1 2 68107 9640
0 9642 5 1 1 9641
0 9643 7 1 2 68342 9622
0 9644 5 1 1 9643
0 9645 7 4 2 69730 83797
0 9646 7 1 2 87179 89016
0 9647 7 1 2 9644 9646
0 9648 5 1 1 9647
0 9649 7 1 2 9642 9648
0 9650 5 1 1 9649
0 9651 7 1 2 61486 9650
0 9652 5 1 1 9651
0 9653 7 4 2 67634 71042
0 9654 5 4 1 89020
0 9655 7 1 2 75605 89024
0 9656 5 2 1 9655
0 9657 7 1 2 69323 89028
0 9658 7 1 2 83004 9657
0 9659 5 1 1 9658
0 9660 7 1 2 64670 9659
0 9661 7 1 2 9652 9660
0 9662 5 1 1 9661
0 9663 7 1 2 63735 9662
0 9664 7 1 2 9617 9663
0 9665 5 1 1 9664
0 9666 7 1 2 9553 9665
0 9667 5 1 1 9666
0 9668 7 1 2 62028 9667
0 9669 5 1 1 9668
0 9670 7 1 2 74902 85050
0 9671 5 1 1 9670
0 9672 7 2 2 62339 71668
0 9673 7 1 2 65092 89030
0 9674 7 1 2 73895 9673
0 9675 5 1 1 9674
0 9676 7 1 2 9671 9675
0 9677 5 1 1 9676
0 9678 7 1 2 66653 9677
0 9679 5 1 1 9678
0 9680 7 2 2 62785 80065
0 9681 5 2 1 89032
0 9682 7 2 2 65093 89034
0 9683 7 2 2 74787 79768
0 9684 5 1 1 89038
0 9685 7 1 2 89036 89039
0 9686 5 1 1 9685
0 9687 7 1 2 9679 9686
0 9688 5 1 1 9687
0 9689 7 1 2 86940 9688
0 9690 5 1 1 9689
0 9691 7 2 2 82407 79966
0 9692 7 2 2 65094 77189
0 9693 7 1 2 89035 89042
0 9694 7 1 2 89040 9693
0 9695 5 1 1 9694
0 9696 7 1 2 9690 9695
0 9697 5 1 1 9696
0 9698 7 1 2 67962 9697
0 9699 5 1 1 9698
0 9700 7 1 2 78863 88502
0 9701 7 2 2 89037 9700
0 9702 7 1 2 77190 89044
0 9703 5 1 1 9702
0 9704 7 1 2 9699 9703
0 9705 5 1 1 9704
0 9706 7 1 2 68108 9705
0 9707 5 1 1 9706
0 9708 7 2 2 67635 74025
0 9709 5 2 1 89046
0 9710 7 2 2 74788 81181
0 9711 5 1 1 89050
0 9712 7 1 2 89048 9711
0 9713 5 1 1 9712
0 9714 7 3 2 81722 77191
0 9715 7 1 2 83581 89052
0 9716 7 1 2 9713 9715
0 9717 5 1 1 9716
0 9718 7 1 2 69731 9717
0 9719 7 1 2 9707 9718
0 9720 5 1 1 9719
0 9721 7 5 2 62786 78864
0 9722 5 4 1 89055
0 9723 7 2 2 62521 78913
0 9724 5 1 1 89064
0 9725 7 1 2 89060 9724
0 9726 5 4 1 9725
0 9727 7 3 2 72931 89066
0 9728 7 1 2 81439 89070
0 9729 5 1 1 9728
0 9730 7 3 2 61782 73153
0 9731 7 1 2 87520 89073
0 9732 5 1 1 9731
0 9733 7 1 2 9729 9732
0 9734 5 1 1 9733
0 9735 7 1 2 66394 9734
0 9736 5 1 1 9735
0 9737 7 15 2 61487 78967
0 9738 5 2 1 89076
0 9739 7 1 2 82575 73694
0 9740 7 1 2 89077 9739
0 9741 5 1 1 9740
0 9742 7 1 2 9736 9741
0 9743 5 1 1 9742
0 9744 7 1 2 79025 9743
0 9745 5 1 1 9744
0 9746 7 1 2 78099 83686
0 9747 5 1 1 9746
0 9748 7 1 2 81808 79003
0 9749 7 1 2 88555 9748
0 9750 5 1 1 9749
0 9751 7 1 2 9747 9750
0 9752 5 1 1 9751
0 9753 7 1 2 64671 73154
0 9754 7 1 2 9752 9753
0 9755 5 1 1 9754
0 9756 7 1 2 9745 9755
0 9757 5 1 1 9756
0 9758 7 1 2 72029 9757
0 9759 5 1 1 9758
0 9760 7 1 2 79669 86204
0 9761 5 1 1 9760
0 9762 7 1 2 80906 82150
0 9763 7 1 2 80870 9762
0 9764 5 1 1 9763
0 9765 7 1 2 9761 9764
0 9766 5 1 1 9765
0 9767 7 1 2 67636 9766
0 9768 5 1 1 9767
0 9769 7 3 2 74789 79732
0 9770 7 1 2 87061 80073
0 9771 7 1 2 89093 9770
0 9772 5 1 1 9771
0 9773 7 1 2 9768 9772
0 9774 5 1 1 9773
0 9775 7 1 2 76125 9774
0 9776 5 1 1 9775
0 9777 7 1 2 78494 89045
0 9778 5 1 1 9777
0 9779 7 1 2 9776 9778
0 9780 5 1 1 9779
0 9781 7 1 2 68109 9780
0 9782 5 1 1 9781
0 9783 7 1 2 82131 83582
0 9784 7 2 2 88989 9783
0 9785 7 1 2 63094 82151
0 9786 7 1 2 89096 9785
0 9787 5 1 1 9786
0 9788 7 1 2 80074 82209
0 9789 5 1 1 9788
0 9790 7 1 2 89049 9789
0 9791 5 1 1 9790
0 9792 7 2 2 69972 81648
0 9793 7 1 2 84122 89098
0 9794 7 1 2 9791 9793
0 9795 5 1 1 9794
0 9796 7 1 2 9787 9795
0 9797 5 1 1 9796
0 9798 7 1 2 66395 9797
0 9799 5 1 1 9798
0 9800 7 1 2 81649 86756
0 9801 7 1 2 89097 9800
0 9802 5 1 1 9801
0 9803 7 1 2 64884 9802
0 9804 7 1 2 9799 9803
0 9805 7 1 2 9782 9804
0 9806 7 1 2 9759 9805
0 9807 5 1 1 9806
0 9808 7 1 2 66892 9807
0 9809 7 1 2 9720 9808
0 9810 5 1 1 9809
0 9811 7 2 2 68343 71632
0 9812 7 1 2 88862 74007
0 9813 7 1 2 89100 9812
0 9814 7 1 2 82764 9813
0 9815 5 1 1 9814
0 9816 7 1 2 9810 9815
0 9817 5 1 1 9816
0 9818 7 1 2 69324 9817
0 9819 5 1 1 9818
0 9820 7 1 2 9669 9819
0 9821 7 1 2 9498 9820
0 9822 5 1 1 9821
0 9823 7 1 2 68793 9822
0 9824 5 1 1 9823
0 9825 7 12 2 68110 65095
0 9826 7 1 2 62340 72768
0 9827 5 1 1 9826
0 9828 7 2 2 63736 9827
0 9829 5 1 1 89114
0 9830 7 1 2 71422 89115
0 9831 5 1 1 9830
0 9832 7 1 2 71043 85994
0 9833 5 1 1 9832
0 9834 7 1 2 9831 9833
0 9835 5 1 1 9834
0 9836 7 1 2 62029 9835
0 9837 5 1 1 9836
0 9838 7 3 2 67392 73569
0 9839 5 5 1 89116
0 9840 7 1 2 75402 80564
0 9841 7 1 2 89117 9840
0 9842 5 1 1 9841
0 9843 7 1 2 9837 9842
0 9844 5 1 1 9843
0 9845 7 1 2 89102 9844
0 9846 5 1 1 9845
0 9847 7 1 2 73570 88883
0 9848 7 1 2 85314 9847
0 9849 5 1 1 9848
0 9850 7 1 2 9846 9849
0 9851 5 1 1 9850
0 9852 7 1 2 67963 9851
0 9853 5 1 1 9852
0 9854 7 1 2 67177 78822
0 9855 7 1 2 78837 9854
0 9856 7 2 2 68585 81750
0 9857 7 1 2 89118 89124
0 9858 7 1 2 9855 9857
0 9859 5 1 1 9858
0 9860 7 1 2 9853 9859
0 9861 5 1 1 9860
0 9862 7 1 2 69325 9861
0 9863 5 1 1 9862
0 9864 7 2 2 81694 80820
0 9865 7 1 2 86785 89126
0 9866 7 1 2 88742 9865
0 9867 5 1 1 9866
0 9868 7 1 2 9863 9867
0 9869 5 1 1 9868
0 9870 7 1 2 68344 9869
0 9871 5 1 1 9870
0 9872 7 2 2 78542 74429
0 9873 5 1 1 89128
0 9874 7 5 2 63737 76760
0 9875 7 1 2 82655 88730
0 9876 7 1 2 89130 9875
0 9877 7 1 2 89129 9876
0 9878 5 1 1 9877
0 9879 7 1 2 72030 78595
0 9880 7 1 2 87671 87424
0 9881 7 1 2 9879 9880
0 9882 7 1 2 88746 9881
0 9883 5 1 1 9882
0 9884 7 1 2 9878 9883
0 9885 5 1 1 9884
0 9886 7 1 2 62522 9885
0 9887 5 1 1 9886
0 9888 7 3 2 75471 78596
0 9889 5 1 1 89135
0 9890 7 1 2 68111 88071
0 9891 7 1 2 89136 9890
0 9892 5 1 1 9891
0 9893 7 2 2 88378 84497
0 9894 7 2 2 61783 81613
0 9895 7 1 2 75993 75507
0 9896 7 1 2 89140 9895
0 9897 7 1 2 89138 9896
0 9898 5 1 1 9897
0 9899 7 1 2 9892 9898
0 9900 5 1 1 9899
0 9901 7 1 2 62341 9900
0 9902 5 1 1 9901
0 9903 7 1 2 82617 83392
0 9904 7 1 2 71689 9903
0 9905 7 1 2 82797 9904
0 9906 7 1 2 79670 9905
0 9907 5 1 1 9906
0 9908 7 1 2 9902 9907
0 9909 7 1 2 9887 9908
0 9910 7 1 2 9871 9909
0 9911 5 1 1 9910
0 9912 7 1 2 61488 9911
0 9913 5 1 1 9912
0 9914 7 3 2 61784 78597
0 9915 7 1 2 88210 89142
0 9916 5 1 1 9915
0 9917 7 2 2 87180 71703
0 9918 5 3 1 89145
0 9919 7 1 2 9916 89147
0 9920 5 1 1 9919
0 9921 7 1 2 68345 73571
0 9922 7 1 2 9920 9921
0 9923 5 1 1 9922
0 9924 7 1 2 66654 78598
0 9925 7 1 2 81182 82265
0 9926 7 1 2 9924 9925
0 9927 5 1 1 9926
0 9928 7 1 2 9923 9927
0 9929 5 1 1 9928
0 9930 7 1 2 63095 9929
0 9931 5 1 1 9930
0 9932 7 2 2 81723 75698
0 9933 7 1 2 78100 79853
0 9934 7 1 2 89150 9933
0 9935 5 1 1 9934
0 9936 7 1 2 9931 9935
0 9937 5 1 1 9936
0 9938 7 1 2 78652 9937
0 9939 5 1 1 9938
0 9940 7 1 2 71044 85859
0 9941 5 1 1 9940
0 9942 7 2 2 69732 70990
0 9943 5 1 1 89152
0 9944 7 1 2 68586 89153
0 9945 5 1 1 9944
0 9946 7 1 2 9941 9945
0 9947 5 1 1 9946
0 9948 7 1 2 72031 9947
0 9949 5 1 1 9948
0 9950 7 1 2 71503 9829
0 9951 5 1 1 9950
0 9952 7 1 2 71423 9951
0 9953 5 1 1 9952
0 9954 7 1 2 9949 9953
0 9955 5 1 1 9954
0 9956 7 1 2 62030 81791
0 9957 7 1 2 9955 9956
0 9958 5 1 1 9957
0 9959 7 1 2 9939 9958
0 9960 5 1 1 9959
0 9961 7 1 2 82109 9960
0 9962 5 1 1 9961
0 9963 7 1 2 64672 9962
0 9964 7 1 2 9913 9963
0 9965 5 1 1 9964
0 9966 7 1 2 83034 83480
0 9967 5 1 1 9966
0 9968 7 1 2 89148 9967
0 9969 5 1 1 9968
0 9970 7 1 2 61489 85761
0 9971 7 1 2 9969 9970
0 9972 5 1 1 9971
0 9973 7 1 2 73572 75508
0 9974 5 1 1 9973
0 9975 7 1 2 85996 9974
0 9976 5 1 1 9975
0 9977 7 1 2 83673 83312
0 9978 7 1 2 9976 9977
0 9979 5 1 1 9978
0 9980 7 1 2 9972 9979
0 9981 5 1 1 9980
0 9982 7 1 2 64472 9981
0 9983 5 1 1 9982
0 9984 7 2 2 82876 87425
0 9985 7 2 2 64885 73573
0 9986 7 1 2 81663 87463
0 9987 7 1 2 89156 9986
0 9988 7 1 2 89154 9987
0 9989 5 1 1 9988
0 9990 7 1 2 9983 9989
0 9991 5 1 1 9990
0 9992 7 1 2 63096 9991
0 9993 5 1 1 9992
0 9994 7 1 2 80925 89146
0 9995 5 1 1 9994
0 9996 7 1 2 88211 88680
0 9997 7 1 2 83321 9996
0 9998 5 1 1 9997
0 9999 7 1 2 9995 9998
0 10000 5 1 1 9999
0 10001 7 1 2 67393 84068
0 10002 7 1 2 10000 10001
0 10003 5 1 1 10002
0 10004 7 1 2 9993 10003
0 10005 5 1 1 10004
0 10006 7 1 2 68346 10005
0 10007 5 1 1 10006
0 10008 7 14 2 66396 67178
0 10009 7 1 2 81650 85704
0 10010 7 2 2 89158 10009
0 10011 7 2 2 78062 88965
0 10012 7 1 2 85889 89174
0 10013 7 1 2 89172 10012
0 10014 5 1 1 10013
0 10015 7 1 2 10007 10014
0 10016 5 1 1 10015
0 10017 7 1 2 66893 10016
0 10018 5 1 1 10017
0 10019 7 1 2 87024 82231
0 10020 7 3 2 72032 88826
0 10021 7 5 2 71912 76126
0 10022 7 1 2 89176 89179
0 10023 7 1 2 10019 10022
0 10024 5 1 1 10023
0 10025 7 1 2 69522 10024
0 10026 7 1 2 10018 10025
0 10027 5 1 1 10026
0 10028 7 1 2 9965 10027
0 10029 5 1 1 10028
0 10030 7 1 2 9824 10029
0 10031 7 1 2 9377 10030
0 10032 5 1 1 10031
0 10033 7 1 2 65355 10032
0 10034 5 1 1 10033
0 10035 7 4 2 82598 83378
0 10036 5 1 1 89184
0 10037 7 1 2 10036 84137
0 10038 5 2 1 10037
0 10039 7 1 2 62031 89188
0 10040 5 1 1 10039
0 10041 7 1 2 9519 10040
0 10042 5 1 1 10041
0 10043 7 1 2 71669 10042
0 10044 5 1 1 10043
0 10045 7 2 2 74235 84895
0 10046 7 1 2 82450 89190
0 10047 5 1 1 10046
0 10048 7 1 2 10044 10047
0 10049 5 1 1 10048
0 10050 7 1 2 69973 10049
0 10051 5 1 1 10050
0 10052 7 2 2 76845 79465
0 10053 7 2 2 82576 72220
0 10054 7 1 2 89192 89194
0 10055 5 1 1 10054
0 10056 7 1 2 10051 10055
0 10057 5 1 1 10056
0 10058 7 1 2 66655 10057
0 10059 5 1 1 10058
0 10060 7 2 2 74352 71670
0 10061 5 1 1 89196
0 10062 7 7 2 63506 70874
0 10063 5 1 1 89198
0 10064 7 1 2 73155 89199
0 10065 5 1 1 10064
0 10066 7 1 2 10061 10065
0 10067 5 1 1 10066
0 10068 7 1 2 83540 10067
0 10069 5 1 1 10068
0 10070 7 7 2 65096 83406
0 10071 5 1 1 89205
0 10072 7 1 2 73540 89206
0 10073 5 1 1 10072
0 10074 7 1 2 10069 10073
0 10075 5 1 1 10074
0 10076 7 1 2 69733 10075
0 10077 5 1 1 10076
0 10078 7 4 2 64886 84445
0 10079 7 2 2 62787 81614
0 10080 7 1 2 89212 89216
0 10081 5 1 1 10080
0 10082 7 1 2 10077 10081
0 10083 5 1 1 10082
0 10084 7 1 2 86875 10083
0 10085 5 1 1 10084
0 10086 7 1 2 10059 10085
0 10087 5 1 1 10086
0 10088 7 1 2 67964 10087
0 10089 5 1 1 10088
0 10090 7 2 2 61785 88896
0 10091 7 2 2 81125 89218
0 10092 7 2 2 69734 84446
0 10093 7 1 2 81751 89222
0 10094 7 1 2 89220 10093
0 10095 5 1 1 10094
0 10096 7 1 2 61490 10095
0 10097 7 1 2 10089 10096
0 10098 5 1 1 10097
0 10099 7 1 2 88933 78724
0 10100 5 1 1 10099
0 10101 7 3 2 68347 76571
0 10102 7 1 2 89013 89224
0 10103 5 1 1 10102
0 10104 7 1 2 10100 10103
0 10105 5 1 1 10104
0 10106 7 1 2 71467 10105
0 10107 5 1 1 10106
0 10108 7 1 2 85890 78543
0 10109 7 1 2 73695 74215
0 10110 7 1 2 10108 10109
0 10111 5 1 1 10110
0 10112 7 1 2 10107 10111
0 10113 5 1 1 10112
0 10114 7 1 2 69523 10113
0 10115 5 1 1 10114
0 10116 7 1 2 79790 80134
0 10117 5 1 1 10116
0 10118 7 1 2 10115 10117
0 10119 5 1 1 10118
0 10120 7 1 2 62523 10119
0 10121 5 1 1 10120
0 10122 7 2 2 80343 79386
0 10123 7 1 2 80410 89074
0 10124 7 1 2 89227 10123
0 10125 5 1 1 10124
0 10126 7 1 2 10121 10125
0 10127 5 1 1 10126
0 10128 7 1 2 68112 10127
0 10129 5 1 1 10128
0 10130 7 1 2 66656 80344
0 10131 5 1 1 10130
0 10132 7 1 2 71093 10131
0 10133 5 5 1 10132
0 10134 7 1 2 71671 89229
0 10135 5 1 1 10134
0 10136 7 3 2 67394 73541
0 10137 5 1 1 89234
0 10138 7 1 2 71045 89235
0 10139 5 1 1 10138
0 10140 7 1 2 10135 10139
0 10141 5 2 1 10140
0 10142 7 1 2 88158 89237
0 10143 5 1 1 10142
0 10144 7 1 2 78638 1290
0 10145 5 1 1 10144
0 10146 7 1 2 74353 10145
0 10147 5 1 1 10146
0 10148 7 1 2 82950 89191
0 10149 5 1 1 10148
0 10150 7 1 2 10147 10149
0 10151 5 1 1 10150
0 10152 7 1 2 81487 10151
0 10153 5 1 1 10152
0 10154 7 1 2 10143 10153
0 10155 5 1 1 10154
0 10156 7 1 2 69974 10155
0 10157 5 1 1 10156
0 10158 7 3 2 64473 78690
0 10159 7 1 2 80907 89239
0 10160 5 1 1 10159
0 10161 7 2 2 67637 78788
0 10162 7 1 2 89242 83994
0 10163 5 1 1 10162
0 10164 7 1 2 10160 10163
0 10165 5 1 1 10164
0 10166 7 1 2 81981 10165
0 10167 5 1 1 10166
0 10168 7 1 2 89071 82640
0 10169 5 1 1 10168
0 10170 7 1 2 10167 10169
0 10171 5 1 1 10170
0 10172 7 1 2 76572 10171
0 10173 5 1 1 10172
0 10174 7 1 2 10157 10173
0 10175 5 1 1 10174
0 10176 7 1 2 63274 10175
0 10177 5 1 1 10176
0 10178 7 1 2 66397 10177
0 10179 7 1 2 10129 10178
0 10180 5 1 1 10179
0 10181 7 1 2 64085 10180
0 10182 7 1 2 10098 10181
0 10183 5 1 1 10182
0 10184 7 2 2 74354 83171
0 10185 5 1 1 89244
0 10186 7 2 2 83982 89245
0 10187 5 1 1 89246
0 10188 7 1 2 79786 85058
0 10189 5 1 1 10188
0 10190 7 1 2 10187 10189
0 10191 5 1 1 10190
0 10192 7 1 2 63097 10191
0 10193 5 1 1 10192
0 10194 7 1 2 89141 81686
0 10195 5 1 1 10194
0 10196 7 1 2 82775 76573
0 10197 7 1 2 87102 10196
0 10198 5 1 1 10197
0 10199 7 1 2 10195 10198
0 10200 5 1 1 10199
0 10201 7 1 2 84069 10200
0 10202 5 1 1 10201
0 10203 7 1 2 10193 10202
0 10204 5 1 1 10203
0 10205 7 1 2 66398 10204
0 10206 5 1 1 10205
0 10207 7 1 2 76038 89247
0 10208 5 1 1 10207
0 10209 7 1 2 10206 10208
0 10210 5 1 1 10209
0 10211 7 1 2 62524 71123
0 10212 7 1 2 10210 10211
0 10213 5 1 1 10212
0 10214 7 1 2 10183 10213
0 10215 5 1 1 10214
0 10216 7 1 2 68794 10215
0 10217 5 1 1 10216
0 10218 7 4 2 69524 78599
0 10219 7 1 2 83427 89248
0 10220 5 1 1 10219
0 10221 7 3 2 79070 85417
0 10222 5 1 1 89252
0 10223 7 1 2 74355 89253
0 10224 5 1 1 10223
0 10225 7 1 2 81147 81837
0 10226 5 1 1 10225
0 10227 7 1 2 10224 10226
0 10228 5 1 1 10227
0 10229 7 1 2 69975 10228
0 10230 5 1 1 10229
0 10231 7 1 2 10220 10230
0 10232 5 1 1 10231
0 10233 7 1 2 63098 10232
0 10234 5 1 1 10233
0 10235 7 21 2 61491 69525
0 10236 5 2 1 89255
0 10237 7 2 2 87613 89256
0 10238 7 1 2 81724 89278
0 10239 5 1 1 10238
0 10240 7 1 2 10234 10239
0 10241 5 1 1 10240
0 10242 7 9 2 61786 62525
0 10243 7 4 2 62788 89280
0 10244 7 1 2 87515 89289
0 10245 7 1 2 10241 10244
0 10246 5 1 1 10245
0 10247 7 1 2 10217 10246
0 10248 5 1 1 10247
0 10249 7 1 2 72984 10248
0 10250 5 1 1 10249
0 10251 7 3 2 63914 72602
0 10252 5 12 1 89293
0 10253 7 1 2 89021 89296
0 10254 5 1 1 10253
0 10255 7 4 2 63915 72033
0 10256 5 2 1 89308
0 10257 7 1 2 75603 89312
0 10258 5 1 1 10257
0 10259 7 1 2 10254 10258
0 10260 5 1 1 10259
0 10261 7 1 2 71913 88631
0 10262 7 1 2 10260 10261
0 10263 5 1 1 10262
0 10264 7 1 2 89309 88047
0 10265 5 1 1 10264
0 10266 7 1 2 670 10265
0 10267 5 1 1 10266
0 10268 7 1 2 78495 89103
0 10269 7 1 2 10267 10268
0 10270 5 1 1 10269
0 10271 7 1 2 10263 10270
0 10272 5 1 1 10271
0 10273 7 1 2 81126 10272
0 10274 5 1 1 10273
0 10275 7 2 2 69526 83451
0 10276 7 3 2 89297 84944
0 10277 5 1 1 89316
0 10278 7 1 2 89314 89317
0 10279 5 1 1 10278
0 10280 7 2 2 62342 74675
0 10281 7 1 2 85874 89319
0 10282 5 1 1 10281
0 10283 7 1 2 63738 86411
0 10284 5 1 1 10283
0 10285 7 1 2 68348 10284
0 10286 5 1 1 10285
0 10287 7 1 2 62343 10286
0 10288 5 1 1 10287
0 10289 7 1 2 68587 86400
0 10290 5 1 1 10289
0 10291 7 1 2 63507 10290
0 10292 5 2 1 10291
0 10293 7 1 2 69976 89321
0 10294 7 1 2 10288 10293
0 10295 5 1 1 10294
0 10296 7 1 2 10282 10295
0 10297 5 1 1 10296
0 10298 7 1 2 67395 87353
0 10299 7 1 2 10297 10298
0 10300 5 1 1 10299
0 10301 7 1 2 10279 10300
0 10302 5 1 1 10301
0 10303 7 1 2 81440 10302
0 10304 5 1 1 10303
0 10305 7 3 2 77060 89298
0 10306 7 2 2 64673 88588
0 10307 5 1 1 89326
0 10308 7 1 2 89323 89327
0 10309 5 1 1 10308
0 10310 7 1 2 71914 85525
0 10311 5 1 1 10310
0 10312 7 1 2 10311 85520
0 10313 5 1 1 10312
0 10314 7 4 2 66399 69977
0 10315 7 1 2 80908 89328
0 10316 7 1 2 10313 10315
0 10317 5 1 1 10316
0 10318 7 1 2 10309 10317
0 10319 5 1 1 10318
0 10320 7 1 2 83035 10319
0 10321 5 1 1 10320
0 10322 7 1 2 10304 10321
0 10323 5 1 1 10322
0 10324 7 1 2 67638 10323
0 10325 5 1 1 10324
0 10326 7 2 2 73399 86016
0 10327 7 1 2 80916 85638
0 10328 7 1 2 89332 10327
0 10329 5 1 1 10328
0 10330 7 5 2 64086 75071
0 10331 7 1 2 78804 89334
0 10332 7 1 2 88632 10331
0 10333 5 1 1 10332
0 10334 7 1 2 10329 10333
0 10335 5 1 1 10334
0 10336 7 1 2 61787 10335
0 10337 5 1 1 10336
0 10338 7 2 2 78983 80624
0 10339 7 1 2 82587 86017
0 10340 7 1 2 89339 10339
0 10341 5 1 1 10340
0 10342 7 1 2 64887 10341
0 10343 7 1 2 10337 10342
0 10344 7 1 2 10325 10343
0 10345 5 1 1 10344
0 10346 7 1 2 63739 85521
0 10347 5 1 1 10346
0 10348 7 1 2 68349 10347
0 10349 5 1 1 10348
0 10350 7 1 2 62344 10349
0 10351 5 1 1 10350
0 10352 7 1 2 68350 89299
0 10353 5 1 1 10352
0 10354 7 1 2 62526 10353
0 10355 5 1 1 10354
0 10356 7 1 2 89322 10355
0 10357 7 2 2 10351 10356
0 10358 7 1 2 69978 89341
0 10359 5 1 1 10358
0 10360 7 1 2 87864 84993
0 10361 5 1 1 10360
0 10362 7 1 2 10359 10361
0 10363 5 1 1 10362
0 10364 7 6 2 64674 82368
0 10365 7 1 2 80926 89343
0 10366 7 1 2 10363 10365
0 10367 5 1 1 10366
0 10368 7 2 2 63508 79746
0 10369 7 1 2 82304 89349
0 10370 5 1 1 10369
0 10371 7 3 2 67639 78101
0 10372 5 2 1 89351
0 10373 7 3 2 81910 73400
0 10374 5 1 1 89356
0 10375 7 1 2 89352 89357
0 10376 5 1 1 10375
0 10377 7 1 2 10370 10376
0 10378 5 1 1 10377
0 10379 7 1 2 86018 10378
0 10380 5 1 1 10379
0 10381 7 8 2 66400 68947
0 10382 7 4 2 69527 89359
0 10383 5 1 1 89367
0 10384 7 1 2 71915 85494
0 10385 7 1 2 89368 10384
0 10386 5 1 1 10385
0 10387 7 2 2 67179 86257
0 10388 7 1 2 61492 89371
0 10389 5 1 1 10388
0 10390 7 1 2 10386 10389
0 10391 5 1 1 10390
0 10392 7 1 2 78102 10391
0 10393 5 1 1 10392
0 10394 7 1 2 10380 10393
0 10395 5 1 1 10394
0 10396 7 1 2 82732 10395
0 10397 5 1 1 10396
0 10398 7 1 2 69735 10397
0 10399 7 1 2 10367 10398
0 10400 5 1 1 10399
0 10401 7 1 2 66894 10400
0 10402 7 1 2 10345 10401
0 10403 5 1 1 10402
0 10404 7 1 2 10274 10403
0 10405 5 1 1 10404
0 10406 7 1 2 69326 10405
0 10407 5 1 1 10406
0 10408 7 1 2 76291 83407
0 10409 5 3 1 10408
0 10410 7 3 2 78063 83092
0 10411 7 1 2 84311 89376
0 10412 5 1 1 10411
0 10413 7 1 2 89373 10412
0 10414 5 1 1 10413
0 10415 7 1 2 62032 10414
0 10416 5 1 1 10415
0 10417 7 1 2 75403 83431
0 10418 5 1 1 10417
0 10419 7 1 2 10416 10418
0 10420 5 1 1 10419
0 10421 7 1 2 71916 10420
0 10422 5 1 1 10421
0 10423 7 6 2 63740 76644
0 10424 7 1 2 88660 89379
0 10425 7 1 2 84394 10424
0 10426 5 1 1 10425
0 10427 7 1 2 10422 10426
0 10428 5 1 1 10427
0 10429 7 1 2 68795 10428
0 10430 5 1 1 10429
0 10431 7 2 2 70875 83172
0 10432 7 1 2 89335 89385
0 10433 5 1 1 10432
0 10434 7 1 2 79288 81295
0 10435 7 1 2 85958 10434
0 10436 5 1 1 10435
0 10437 7 1 2 10433 10436
0 10438 5 1 1 10437
0 10439 7 1 2 75135 10438
0 10440 5 1 1 10439
0 10441 7 2 2 68948 74430
0 10442 7 2 2 77372 89387
0 10443 7 4 2 71917 83093
0 10444 7 2 2 65955 89391
0 10445 7 1 2 89389 89395
0 10446 5 1 1 10445
0 10447 7 1 2 10440 10446
0 10448 7 1 2 10430 10447
0 10449 5 1 1 10448
0 10450 7 1 2 69736 10449
0 10451 5 1 1 10450
0 10452 7 1 2 88966 82516
0 10453 7 1 2 89318 10452
0 10454 5 1 1 10453
0 10455 7 1 2 10451 10454
0 10456 5 1 1 10455
0 10457 7 1 2 83948 10456
0 10458 5 1 1 10457
0 10459 7 1 2 10407 10458
0 10460 5 1 1 10459
0 10461 7 1 2 67965 10460
0 10462 5 1 1 10461
0 10463 7 1 2 67640 88939
0 10464 5 1 1 10463
0 10465 7 1 2 88981 10464
0 10466 5 3 1 10465
0 10467 7 1 2 75761 89397
0 10468 5 1 1 10467
0 10469 7 1 2 78176 81405
0 10470 5 1 1 10469
0 10471 7 1 2 10468 10470
0 10472 5 1 1 10471
0 10473 7 1 2 72527 10472
0 10474 5 1 1 10473
0 10475 7 1 2 77083 81571
0 10476 5 1 1 10475
0 10477 7 1 2 10474 10476
0 10478 5 1 1 10477
0 10479 7 1 2 61788 10478
0 10480 5 1 1 10479
0 10481 7 1 2 81406 84655
0 10482 7 1 2 76233 10481
0 10483 5 1 1 10482
0 10484 7 1 2 10480 10483
0 10485 5 1 1 10484
0 10486 7 1 2 79344 10485
0 10487 5 1 1 10486
0 10488 7 1 2 83628 75590
0 10489 5 2 1 10488
0 10490 7 3 2 61789 82232
0 10491 7 1 2 81400 89402
0 10492 5 1 1 10491
0 10493 7 1 2 89400 10492
0 10494 5 1 1 10493
0 10495 7 1 2 74309 10494
0 10496 5 1 1 10495
0 10497 7 3 2 68796 69737
0 10498 7 4 2 79345 89405
0 10499 7 1 2 75825 89408
0 10500 5 1 1 10499
0 10501 7 1 2 10496 10500
0 10502 5 1 1 10501
0 10503 7 1 2 63275 10502
0 10504 5 1 1 10503
0 10505 7 2 2 83036 75762
0 10506 7 1 2 89409 89412
0 10507 5 1 1 10506
0 10508 7 1 2 10504 10507
0 10509 5 1 1 10508
0 10510 7 1 2 84312 10509
0 10511 5 1 1 10510
0 10512 7 1 2 10487 10511
0 10513 5 1 1 10512
0 10514 7 1 2 69979 10513
0 10515 5 1 1 10514
0 10516 7 2 2 84145 86249
0 10517 7 1 2 89137 89414
0 10518 5 1 1 10517
0 10519 7 1 2 10515 10518
0 10520 5 1 1 10519
0 10521 7 1 2 71918 10520
0 10522 5 1 1 10521
0 10523 7 1 2 63276 89324
0 10524 5 1 1 10523
0 10525 7 1 2 82266 85832
0 10526 5 1 1 10525
0 10527 7 1 2 10524 10526
0 10528 5 1 1 10527
0 10529 7 1 2 61790 10528
0 10530 5 1 1 10529
0 10531 7 3 2 73542 87448
0 10532 5 1 1 89416
0 10533 7 2 2 69980 89417
0 10534 5 1 1 89419
0 10535 7 1 2 87636 89420
0 10536 5 1 1 10535
0 10537 7 1 2 10530 10536
0 10538 5 1 1 10537
0 10539 7 1 2 79346 10538
0 10540 5 1 1 10539
0 10541 7 2 2 83379 87464
0 10542 7 1 2 75591 86019
0 10543 7 1 2 89421 10542
0 10544 5 1 1 10543
0 10545 7 1 2 10540 10544
0 10546 5 1 1 10545
0 10547 7 1 2 69738 10546
0 10548 5 1 1 10547
0 10549 7 1 2 75699 89185
0 10550 7 1 2 89325 10549
0 10551 5 1 1 10550
0 10552 7 1 2 10548 10551
0 10553 5 1 1 10552
0 10554 7 1 2 75136 10553
0 10555 5 1 1 10554
0 10556 7 3 2 69981 83923
0 10557 7 1 2 84810 89423
0 10558 5 1 1 10557
0 10559 7 5 2 64888 79799
0 10560 7 3 2 88240 89426
0 10561 5 1 1 89431
0 10562 7 1 2 83917 10561
0 10563 5 1 1 10562
0 10564 7 1 2 82965 10563
0 10565 5 1 1 10564
0 10566 7 1 2 10558 10565
0 10567 5 1 1 10566
0 10568 7 1 2 66895 10567
0 10569 5 1 1 10568
0 10570 7 4 2 66657 71690
0 10571 5 1 1 89434
0 10572 7 1 2 71094 10571
0 10573 5 2 1 10572
0 10574 7 1 2 76817 88614
0 10575 7 1 2 89438 10574
0 10576 5 1 1 10575
0 10577 7 1 2 10569 10576
0 10578 5 1 1 10577
0 10579 7 1 2 74067 10578
0 10580 5 1 1 10579
0 10581 7 1 2 78632 78577
0 10582 5 1 1 10581
0 10583 7 6 2 64474 80043
0 10584 7 1 2 89131 89440
0 10585 7 1 2 10582 10584
0 10586 5 1 1 10585
0 10587 7 1 2 10580 10586
0 10588 5 1 1 10587
0 10589 7 1 2 63277 85271
0 10590 7 1 2 10588 10589
0 10591 5 1 1 10590
0 10592 7 2 2 89186 76993
0 10593 7 2 2 65097 74026
0 10594 5 1 1 89448
0 10595 7 2 2 64087 77929
0 10596 5 1 1 89450
0 10597 7 1 2 89449 89451
0 10598 7 1 2 89446 10597
0 10599 5 1 1 10598
0 10600 7 1 2 10591 10599
0 10601 7 1 2 10555 10600
0 10602 7 1 2 10522 10601
0 10603 5 1 1 10602
0 10604 7 1 2 66401 10603
0 10605 5 1 1 10604
0 10606 7 1 2 61791 81385
0 10607 5 1 1 10606
0 10608 7 1 2 10607 3314
0 10609 5 5 1 10608
0 10610 7 1 2 67396 89452
0 10611 5 1 1 10610
0 10612 7 1 2 81367 84103
0 10613 5 1 1 10612
0 10614 7 1 2 10611 10613
0 10615 5 1 1 10614
0 10616 7 1 2 74310 10615
0 10617 5 1 1 10616
0 10618 7 1 2 69739 83495
0 10619 7 1 2 85020 10618
0 10620 5 1 1 10619
0 10621 7 5 2 74311 83037
0 10622 5 1 1 89457
0 10623 7 2 2 79071 89458
0 10624 5 1 1 89462
0 10625 7 1 2 10620 10624
0 10626 5 1 1 10625
0 10627 7 1 2 68797 10626
0 10628 5 1 1 10627
0 10629 7 6 2 67641 72116
0 10630 5 6 1 89464
0 10631 7 1 2 74312 81386
0 10632 5 2 1 10631
0 10633 7 8 2 63509 84524
0 10634 7 2 2 78472 89478
0 10635 5 1 1 89486
0 10636 7 1 2 89476 10635
0 10637 5 1 1 10636
0 10638 7 1 2 61792 10637
0 10639 5 1 1 10638
0 10640 7 4 2 66896 83408
0 10641 5 1 1 89488
0 10642 7 1 2 79099 89489
0 10643 5 2 1 10642
0 10644 7 1 2 10639 89492
0 10645 5 1 1 10644
0 10646 7 1 2 89465 10645
0 10647 5 1 1 10646
0 10648 7 1 2 10628 10647
0 10649 7 1 2 10617 10648
0 10650 5 1 1 10649
0 10651 7 1 2 71919 10650
0 10652 5 1 1 10651
0 10653 7 10 2 72603 89470
0 10654 5 22 1 89494
0 10655 7 3 2 66897 71205
0 10656 7 1 2 74862 89526
0 10657 7 1 2 89504 10656
0 10658 7 1 2 89453 10657
0 10659 5 1 1 10658
0 10660 7 1 2 10652 10659
0 10661 5 1 1 10660
0 10662 7 1 2 69982 10661
0 10663 5 1 1 10662
0 10664 7 3 2 76645 74676
0 10665 5 2 1 89529
0 10666 7 1 2 84781 89530
0 10667 7 1 2 79170 10666
0 10668 7 1 2 84395 10667
0 10669 5 1 1 10668
0 10670 7 1 2 10663 10669
0 10671 5 1 1 10670
0 10672 7 1 2 82839 10671
0 10673 5 1 1 10672
0 10674 7 1 2 10605 10673
0 10675 5 1 1 10674
0 10676 7 1 2 63099 10675
0 10677 5 1 1 10676
0 10678 7 1 2 10462 10677
0 10679 7 1 2 10250 10678
0 10680 5 1 1 10679
0 10681 7 1 2 70269 10680
0 10682 5 1 1 10681
0 10683 7 1 2 73804 83655
0 10684 5 1 1 10683
0 10685 7 1 2 81203 86264
0 10686 5 1 1 10685
0 10687 7 1 2 10684 10686
0 10688 5 1 1 10687
0 10689 7 1 2 74981 10688
0 10690 5 1 1 10689
0 10691 7 4 2 68798 79427
0 10692 7 3 2 73910 89534
0 10693 7 2 2 66898 72694
0 10694 7 1 2 84328 89541
0 10695 7 1 2 89538 10694
0 10696 5 1 1 10695
0 10697 7 1 2 10690 10696
0 10698 5 1 1 10697
0 10699 7 1 2 61793 10698
0 10700 5 1 1 10699
0 10701 7 1 2 68588 74934
0 10702 7 1 2 84994 10701
0 10703 7 1 2 82819 78666
0 10704 7 1 2 10702 10703
0 10705 5 1 1 10704
0 10706 7 1 2 10700 10705
0 10707 5 1 1 10706
0 10708 7 1 2 68113 10707
0 10709 5 1 1 10708
0 10710 7 1 2 78157 83895
0 10711 5 1 1 10710
0 10712 7 1 2 86135 75358
0 10713 5 1 1 10712
0 10714 7 1 2 10711 10713
0 10715 5 1 1 10714
0 10716 7 1 2 83674 89418
0 10717 7 1 2 10715 10716
0 10718 5 1 1 10717
0 10719 7 1 2 10709 10718
0 10720 5 1 1 10719
0 10721 7 1 2 67180 10720
0 10722 5 1 1 10721
0 10723 7 2 2 66899 73156
0 10724 7 1 2 89543 82821
0 10725 7 1 2 86318 10724
0 10726 7 1 2 89386 10725
0 10727 5 1 1 10726
0 10728 7 1 2 10722 10727
0 10729 5 1 1 10728
0 10730 7 1 2 76127 10729
0 10731 5 1 1 10730
0 10732 7 2 2 76070 84617
0 10733 5 1 1 89545
0 10734 7 1 2 68351 72221
0 10735 7 1 2 86136 10734
0 10736 7 1 2 89546 10735
0 10737 5 1 1 10736
0 10738 7 5 2 67966 87399
0 10739 7 1 2 88685 89547
0 10740 5 1 1 10739
0 10741 7 1 2 68799 83830
0 10742 5 1 1 10741
0 10743 7 1 2 10740 10742
0 10744 5 1 1 10743
0 10745 7 1 2 83496 77084
0 10746 7 1 2 10744 10745
0 10747 5 1 1 10746
0 10748 7 1 2 10737 10747
0 10749 5 1 1 10748
0 10750 7 1 2 84460 10749
0 10751 5 1 1 10750
0 10752 7 3 2 68949 85891
0 10753 7 3 2 66402 80221
0 10754 7 2 2 89552 89555
0 10755 5 1 1 89558
0 10756 7 7 2 64475 89505
0 10757 7 1 2 77227 89560
0 10758 5 1 1 10757
0 10759 7 1 2 10755 10758
0 10760 5 1 1 10759
0 10761 7 6 2 68800 78653
0 10762 7 1 2 89249 89567
0 10763 7 1 2 82713 10762
0 10764 7 1 2 10760 10763
0 10765 5 1 1 10764
0 10766 7 1 2 10751 10765
0 10767 5 1 1 10766
0 10768 7 1 2 67181 10767
0 10769 5 1 1 10768
0 10770 7 5 2 62033 77407
0 10771 5 4 1 89573
0 10772 7 1 2 86941 89574
0 10773 5 1 1 10772
0 10774 7 1 2 86923 75051
0 10775 7 1 2 80639 10774
0 10776 5 1 1 10775
0 10777 7 1 2 10773 10776
0 10778 5 1 1 10777
0 10779 7 1 2 84816 80846
0 10780 7 1 2 89139 10779
0 10781 7 1 2 10778 10780
0 10782 5 1 1 10781
0 10783 7 1 2 10769 10782
0 10784 5 1 1 10783
0 10785 7 1 2 61794 10784
0 10786 5 1 1 10785
0 10787 7 2 2 77228 82426
0 10788 7 1 2 88550 79652
0 10789 7 1 2 89582 10788
0 10790 7 1 2 85905 10789
0 10791 5 1 1 10790
0 10792 7 1 2 10786 10791
0 10793 7 1 2 10731 10792
0 10794 7 1 2 10682 10793
0 10795 7 1 2 10034 10794
0 10796 5 1 1 10795
0 10797 7 1 2 65696 10796
0 10798 5 1 1 10797
0 10799 7 1 2 82192 86401
0 10800 5 1 1 10799
0 10801 7 1 2 1100 10800
0 10802 5 2 1 10801
0 10803 7 1 2 62034 89584
0 10804 5 1 1 10803
0 10805 7 1 2 75087 76411
0 10806 5 1 1 10805
0 10807 7 1 2 10804 10806
0 10808 5 1 1 10807
0 10809 7 1 2 81725 10808
0 10810 5 1 1 10809
0 10811 7 3 2 72819 85495
0 10812 5 2 1 89586
0 10813 7 1 2 87156 89589
0 10814 5 2 1 10813
0 10815 7 7 2 67182 63100
0 10816 7 2 2 68114 89593
0 10817 7 1 2 74313 89600
0 10818 7 1 2 89591 10817
0 10819 5 1 1 10818
0 10820 7 1 2 10810 10819
0 10821 5 1 1 10820
0 10822 7 1 2 89143 10821
0 10823 5 1 1 10822
0 10824 7 2 2 69740 80436
0 10825 7 1 2 89602 74412
0 10826 5 1 1 10825
0 10827 7 2 2 67183 75012
0 10828 5 1 1 89604
0 10829 7 1 2 63510 10828
0 10830 5 1 1 10829
0 10831 7 1 2 75581 10830
0 10832 5 1 1 10831
0 10833 7 1 2 10826 10832
0 10834 5 1 1 10833
0 10835 7 1 2 63916 10834
0 10836 5 1 1 10835
0 10837 7 3 2 74216 83517
0 10838 5 1 1 89606
0 10839 7 1 2 71152 89607
0 10840 5 1 1 10839
0 10841 7 1 2 10836 10840
0 10842 5 1 1 10841
0 10843 7 1 2 70637 10842
0 10844 5 1 1 10843
0 10845 7 2 2 72034 85353
0 10846 5 2 1 89609
0 10847 7 1 2 62345 84313
0 10848 5 1 1 10847
0 10849 7 1 2 89611 10848
0 10850 5 1 1 10849
0 10851 7 2 2 62035 10850
0 10852 5 1 1 89613
0 10853 7 3 2 69741 77167
0 10854 7 1 2 89614 89615
0 10855 5 1 1 10854
0 10856 7 1 2 66900 89585
0 10857 5 1 1 10856
0 10858 7 1 2 86402 85801
0 10859 5 1 1 10858
0 10860 7 1 2 10857 10859
0 10861 5 1 1 10860
0 10862 7 1 2 75994 10861
0 10863 5 1 1 10862
0 10864 7 1 2 10855 10863
0 10865 7 1 2 10844 10864
0 10866 5 1 1 10865
0 10867 7 1 2 68115 10866
0 10868 5 1 1 10867
0 10869 7 1 2 63278 80437
0 10870 7 1 2 89575 10869
0 10871 5 1 1 10870
0 10872 7 1 2 61795 10871
0 10873 7 1 2 10868 10872
0 10874 5 1 1 10873
0 10875 7 1 2 80281 85008
0 10876 5 1 1 10875
0 10877 7 3 2 66901 84858
0 10878 7 1 2 86403 89618
0 10879 5 1 1 10878
0 10880 7 1 2 10876 10879
0 10881 5 1 1 10880
0 10882 7 1 2 75995 10881
0 10883 5 1 1 10882
0 10884 7 4 2 69742 81726
0 10885 7 1 2 71153 79873
0 10886 5 1 1 10885
0 10887 7 2 2 62346 73157
0 10888 7 1 2 89310 89625
0 10889 5 1 1 10888
0 10890 7 1 2 10886 10889
0 10891 5 1 1 10890
0 10892 7 1 2 70638 10891
0 10893 5 2 1 10892
0 10894 7 1 2 89627 10852
0 10895 5 1 1 10894
0 10896 7 1 2 89621 10895
0 10897 5 1 1 10896
0 10898 7 1 2 10883 10897
0 10899 5 1 1 10898
0 10900 7 1 2 63511 10899
0 10901 5 1 1 10900
0 10902 7 4 2 62036 80438
0 10903 7 2 2 77963 89629
0 10904 7 4 2 63917 69743
0 10905 7 1 2 63279 89635
0 10906 7 1 2 71154 10905
0 10907 7 1 2 89633 10906
0 10908 5 1 1 10907
0 10909 7 1 2 66658 10908
0 10910 7 1 2 10901 10909
0 10911 5 1 1 10910
0 10912 7 1 2 69983 10911
0 10913 7 1 2 10874 10912
0 10914 5 1 1 10913
0 10915 7 1 2 10823 10914
0 10916 5 1 1 10915
0 10917 7 1 2 64476 10916
0 10918 5 1 1 10917
0 10919 7 3 2 62789 86723
0 10920 5 2 1 89639
0 10921 7 2 2 67397 89300
0 10922 7 1 2 89642 89644
0 10923 5 1 1 10922
0 10924 7 1 2 68801 84656
0 10925 5 1 1 10924
0 10926 7 1 2 10923 10925
0 10927 5 2 1 10926
0 10928 7 6 2 82877 80027
0 10929 7 1 2 65098 82641
0 10930 7 1 2 89648 10929
0 10931 7 1 2 89646 10930
0 10932 5 1 1 10931
0 10933 7 1 2 10918 10932
0 10934 5 1 1 10933
0 10935 7 1 2 68589 10934
0 10936 5 1 1 10935
0 10937 7 1 2 66902 83442
0 10938 5 1 1 10937
0 10939 7 1 2 73192 73178
0 10940 5 2 1 10939
0 10941 7 1 2 62037 84314
0 10942 5 1 1 10941
0 10943 7 1 2 89654 10942
0 10944 5 2 1 10943
0 10945 7 1 2 88940 89656
0 10946 5 1 1 10945
0 10947 7 1 2 64889 84525
0 10948 5 1 1 10947
0 10949 7 1 2 10946 10948
0 10950 5 1 1 10949
0 10951 7 1 2 78064 10950
0 10952 5 1 1 10951
0 10953 7 1 2 87602 84526
0 10954 5 1 1 10953
0 10955 7 1 2 10952 10954
0 10956 5 1 1 10955
0 10957 7 1 2 67967 10956
0 10958 5 1 1 10957
0 10959 7 1 2 10938 10958
0 10960 5 1 1 10959
0 10961 7 1 2 61796 10960
0 10962 5 1 1 10961
0 10963 7 2 2 69744 81615
0 10964 7 1 2 89099 89658
0 10965 7 1 2 89657 10964
0 10966 5 1 1 10965
0 10967 7 1 2 10962 10966
0 10968 5 1 1 10967
0 10969 7 1 2 63741 10968
0 10970 5 1 1 10969
0 10971 7 2 2 62790 89608
0 10972 5 1 1 89660
0 10973 7 1 2 83173 72332
0 10974 7 1 2 89661 10973
0 10975 5 1 1 10974
0 10976 7 1 2 10970 10975
0 10977 5 1 1 10976
0 10978 7 1 2 67184 10977
0 10979 5 1 1 10978
0 10980 7 2 2 61797 86598
0 10981 7 2 2 82577 89662
0 10982 7 8 2 67968 63918
0 10983 7 2 2 72286 89666
0 10984 7 1 2 89674 87596
0 10985 7 1 2 89664 10984
0 10986 5 1 1 10985
0 10987 7 1 2 10979 10986
0 10988 5 1 1 10987
0 10989 7 1 2 64477 10988
0 10990 5 1 1 10989
0 10991 7 1 2 10936 10990
0 10992 5 1 1 10991
0 10993 7 1 2 65356 10992
0 10994 5 1 1 10993
0 10995 7 1 2 88654 84995
0 10996 5 1 1 10995
0 10997 7 1 2 63742 77618
0 10998 5 2 1 10997
0 10999 7 1 2 81141 89676
0 11000 5 1 1 10999
0 11001 7 3 2 70876 83094
0 11002 7 1 2 84835 89678
0 11003 7 1 2 11000 11002
0 11004 5 1 1 11003
0 11005 7 1 2 10996 11004
0 11006 5 1 1 11005
0 11007 7 1 2 70270 11006
0 11008 5 1 1 11007
0 11009 7 2 2 70639 83174
0 11010 7 1 2 63919 86106
0 11011 7 1 2 89681 11010
0 11012 5 1 1 11011
0 11013 7 1 2 11008 11012
0 11014 5 1 1 11013
0 11015 7 1 2 69745 11014
0 11016 5 1 1 11015
0 11017 7 1 2 88754 74964
0 11018 7 1 2 85318 11017
0 11019 5 2 1 11018
0 11020 7 1 2 11016 89683
0 11021 5 1 1 11020
0 11022 7 1 2 75137 11021
0 11023 5 1 1 11022
0 11024 7 3 2 73543 71633
0 11025 5 1 1 89685
0 11026 7 1 2 74724 11025
0 11027 5 1 1 11026
0 11028 7 1 2 80268 11027
0 11029 5 1 1 11028
0 11030 7 1 2 75509 72243
0 11031 7 1 2 76606 11030
0 11032 5 1 1 11031
0 11033 7 1 2 11029 11032
0 11034 5 1 1 11033
0 11035 7 1 2 67185 11034
0 11036 5 1 1 11035
0 11037 7 2 2 67642 71488
0 11038 7 1 2 89688 73634
0 11039 5 1 1 11038
0 11040 7 1 2 11036 11039
0 11041 5 1 1 11040
0 11042 7 1 2 63512 11041
0 11043 5 1 1 11042
0 11044 7 1 2 71814 84556
0 11045 7 1 2 73723 11044
0 11046 5 1 1 11045
0 11047 7 1 2 11043 11046
0 11048 5 1 1 11047
0 11049 7 1 2 87304 11048
0 11050 5 1 1 11049
0 11051 7 1 2 75510 73193
0 11052 5 1 1 11051
0 11053 7 1 2 2690 11052
0 11054 5 2 1 11053
0 11055 7 1 2 67186 89690
0 11056 5 1 1 11055
0 11057 7 1 2 76646 73874
0 11058 5 1 1 11057
0 11059 7 1 2 11056 11058
0 11060 5 1 1 11059
0 11061 7 2 2 70271 81616
0 11062 7 1 2 84104 89692
0 11063 7 1 2 11060 11062
0 11064 5 1 1 11063
0 11065 7 1 2 11050 11064
0 11066 5 1 1 11065
0 11067 7 1 2 69984 11066
0 11068 5 1 1 11067
0 11069 7 1 2 11023 11068
0 11070 5 1 1 11069
0 11071 7 1 2 67969 11070
0 11072 5 1 1 11071
0 11073 7 4 2 68116 74265
0 11074 5 2 1 89694
0 11075 7 6 2 75472 77439
0 11076 7 1 2 77327 89700
0 11077 7 1 2 89695 11076
0 11078 5 1 1 11077
0 11079 7 2 2 66659 82578
0 11080 5 2 1 89706
0 11081 7 1 2 83038 73401
0 11082 5 1 1 11081
0 11083 7 1 2 89708 11082
0 11084 5 1 1 11083
0 11085 7 1 2 82408 87017
0 11086 7 1 2 87191 11085
0 11087 7 1 2 11084 11086
0 11088 5 1 1 11087
0 11089 7 1 2 11078 11088
0 11090 5 1 1 11089
0 11091 7 1 2 75996 11090
0 11092 5 1 1 11091
0 11093 7 1 2 11072 11092
0 11094 5 1 1 11093
0 11095 7 1 2 64478 11094
0 11096 5 1 1 11095
0 11097 7 1 2 61493 11096
0 11098 7 1 2 10994 11097
0 11099 5 1 1 11098
0 11100 7 3 2 69985 82233
0 11101 7 2 2 71206 84682
0 11102 5 1 1 89713
0 11103 7 1 2 71155 89714
0 11104 5 1 1 11103
0 11105 7 2 2 76245 73681
0 11106 5 1 1 89715
0 11107 7 1 2 11104 11106
0 11108 5 1 1 11107
0 11109 7 1 2 63280 11108
0 11110 5 1 1 11109
0 11111 7 10 2 62347 68117
0 11112 7 1 2 75072 89717
0 11113 7 1 2 79812 11112
0 11114 5 1 1 11113
0 11115 7 1 2 11110 11114
0 11116 5 1 1 11115
0 11117 7 1 2 70640 11116
0 11118 5 1 1 11117
0 11119 7 1 2 74951 78209
0 11120 5 1 1 11119
0 11121 7 2 2 84300 86346
0 11122 5 1 1 89727
0 11123 7 1 2 11120 11122
0 11124 5 1 1 11123
0 11125 7 1 2 73402 11124
0 11126 5 1 1 11125
0 11127 7 3 2 65357 84315
0 11128 5 4 1 89729
0 11129 7 1 2 72985 89730
0 11130 5 1 1 11129
0 11131 7 1 2 11126 11130
0 11132 5 1 1 11131
0 11133 7 1 2 63281 11132
0 11134 5 1 1 11133
0 11135 7 1 2 11118 11134
0 11136 5 1 1 11135
0 11137 7 1 2 61798 11136
0 11138 5 1 1 11137
0 11139 7 3 2 87637 71774
0 11140 7 1 2 80498 89736
0 11141 7 1 2 79569 11140
0 11142 5 1 1 11141
0 11143 7 1 2 11138 11142
0 11144 5 1 1 11143
0 11145 7 1 2 89710 11144
0 11146 5 1 1 11145
0 11147 7 2 2 75939 89104
0 11148 7 1 2 82599 82152
0 11149 7 1 2 89739 11148
0 11150 7 1 2 89647 11149
0 11151 5 1 1 11150
0 11152 7 1 2 11146 11151
0 11153 5 1 1 11152
0 11154 7 1 2 66903 11153
0 11155 5 1 1 11154
0 11156 7 1 2 63920 75206
0 11157 5 1 1 11156
0 11158 7 1 2 75005 11157
0 11159 5 1 1 11158
0 11160 7 1 2 62348 11159
0 11161 5 1 1 11160
0 11162 7 1 2 89677 73878
0 11163 5 1 1 11162
0 11164 7 1 2 11163 87594
0 11165 5 1 1 11164
0 11166 7 1 2 11161 11165
0 11167 5 1 1 11166
0 11168 7 1 2 83095 11167
0 11169 5 1 1 11168
0 11170 7 3 2 65358 71013
0 11171 5 1 1 89741
0 11172 7 1 2 88655 85939
0 11173 7 1 2 89742 11172
0 11174 5 1 1 11173
0 11175 7 1 2 11169 11174
0 11176 5 1 1 11175
0 11177 7 1 2 69986 11176
0 11178 5 1 1 11177
0 11179 7 1 2 73646 72748
0 11180 5 3 1 11179
0 11181 7 1 2 74000 89744
0 11182 5 3 1 11181
0 11183 7 1 2 67187 89747
0 11184 5 1 1 11183
0 11185 7 1 2 75981 11184
0 11186 5 1 1 11185
0 11187 7 1 2 88647 11186
0 11188 5 1 1 11187
0 11189 7 1 2 11178 11188
0 11190 5 1 1 11189
0 11191 7 1 2 69746 11190
0 11192 5 1 1 11191
0 11193 7 1 2 89684 11192
0 11194 5 1 1 11193
0 11195 7 1 2 82680 11194
0 11196 5 1 1 11195
0 11197 7 1 2 11155 11196
0 11198 5 1 1 11197
0 11199 7 1 2 68352 11198
0 11200 5 1 1 11199
0 11201 7 2 2 63921 64479
0 11202 7 1 2 82482 86154
0 11203 5 1 1 11202
0 11204 7 1 2 83605 73174
0 11205 5 1 1 11204
0 11206 7 1 2 11203 11205
0 11207 5 1 1 11206
0 11208 7 1 2 83175 11207
0 11209 5 1 1 11208
0 11210 7 3 2 70272 75473
0 11211 5 1 1 89752
0 11212 7 1 2 80066 89753
0 11213 5 1 1 11212
0 11214 7 1 2 61799 84180
0 11215 5 1 1 11214
0 11216 7 1 2 11213 11215
0 11217 5 1 1 11216
0 11218 7 1 2 63282 79004
0 11219 7 1 2 11217 11218
0 11220 5 1 1 11219
0 11221 7 1 2 11209 11220
0 11222 5 1 1 11221
0 11223 7 1 2 69747 11222
0 11224 5 1 1 11223
0 11225 7 1 2 61800 88481
0 11226 7 3 2 69987 86158
0 11227 7 1 2 74138 89755
0 11228 7 1 2 11225 11227
0 11229 5 1 1 11228
0 11230 7 1 2 11224 11229
0 11231 5 1 1 11230
0 11232 7 1 2 62349 11231
0 11233 5 1 1 11232
0 11234 7 5 2 64890 74108
0 11235 7 1 2 62038 77597
0 11236 7 1 2 89758 11235
0 11237 5 1 1 11236
0 11238 7 1 2 69748 89542
0 11239 7 1 2 85940 11238
0 11240 5 1 1 11239
0 11241 7 1 2 11237 11240
0 11242 5 1 1 11241
0 11243 7 1 2 83675 85506
0 11244 7 1 2 11242 11243
0 11245 5 1 1 11244
0 11246 7 1 2 11233 11245
0 11247 5 1 1 11246
0 11248 7 1 2 70641 11247
0 11249 5 1 1 11248
0 11250 7 2 2 80469 89701
0 11251 7 2 2 76933 80345
0 11252 7 1 2 87558 89765
0 11253 7 1 2 89763 11252
0 11254 5 1 1 11253
0 11255 7 1 2 11249 11254
0 11256 5 1 1 11255
0 11257 7 1 2 89750 11256
0 11258 5 1 1 11257
0 11259 7 1 2 11200 11258
0 11260 5 1 1 11259
0 11261 7 1 2 63101 11260
0 11262 5 1 1 11261
0 11263 7 1 2 83541 74566
0 11264 5 1 1 11263
0 11265 7 4 2 68590 78407
0 11266 7 1 2 63283 89767
0 11267 5 1 1 11266
0 11268 7 1 2 11264 11267
0 11269 5 2 1 11268
0 11270 7 1 2 89771 79863
0 11271 5 1 1 11270
0 11272 7 1 2 74578 79574
0 11273 5 1 1 11272
0 11274 7 1 2 76970 11273
0 11275 5 2 1 11274
0 11276 7 1 2 83409 89773
0 11277 5 1 1 11276
0 11278 7 1 2 11271 11277
0 11279 5 1 1 11278
0 11280 7 1 2 77025 11279
0 11281 5 1 1 11280
0 11282 7 10 2 70273 73403
0 11283 5 1 1 89775
0 11284 7 2 2 68353 84859
0 11285 7 1 2 89785 86426
0 11286 7 1 2 89776 11285
0 11287 5 1 1 11286
0 11288 7 1 2 11281 11287
0 11289 5 1 1 11288
0 11290 7 1 2 64891 11289
0 11291 5 1 1 11290
0 11292 7 2 2 79472 86376
0 11293 5 3 1 89787
0 11294 7 4 2 68591 85245
0 11295 5 1 1 89792
0 11296 7 1 2 65359 89793
0 11297 5 1 1 11296
0 11298 7 1 2 89789 11297
0 11299 5 1 1 11298
0 11300 7 1 2 72117 75052
0 11301 7 1 2 83542 11300
0 11302 7 1 2 11299 11301
0 11303 5 1 1 11302
0 11304 7 1 2 11291 11303
0 11305 5 1 1 11304
0 11306 7 1 2 66660 11305
0 11307 5 1 1 11306
0 11308 7 2 2 72035 74579
0 11309 5 1 1 89796
0 11310 7 2 2 70642 89797
0 11311 5 1 1 89798
0 11312 7 2 2 73404 78210
0 11313 5 1 1 89800
0 11314 7 1 2 11311 11313
0 11315 5 1 1 11314
0 11316 7 1 2 78544 11315
0 11317 5 1 1 11316
0 11318 7 2 2 80871 76772
0 11319 5 3 1 89802
0 11320 7 1 2 86235 89803
0 11321 5 1 1 11320
0 11322 7 1 2 11317 11321
0 11323 5 1 1 11322
0 11324 7 1 2 82878 79769
0 11325 7 1 2 11323 11324
0 11326 5 1 1 11325
0 11327 7 1 2 11307 11326
0 11328 5 1 1 11327
0 11329 7 1 2 67643 11328
0 11330 5 1 1 11329
0 11331 7 3 2 61801 72118
0 11332 7 4 2 64892 79601
0 11333 5 1 1 89810
0 11334 7 1 2 89804 11333
0 11335 5 1 1 11334
0 11336 7 1 2 85514 11335
0 11337 5 1 1 11336
0 11338 7 2 2 65360 85246
0 11339 7 1 2 89756 89814
0 11340 5 1 1 11339
0 11341 7 1 2 11337 11340
0 11342 5 1 1 11341
0 11343 7 1 2 89807 11342
0 11344 5 1 1 11343
0 11345 7 1 2 75940 80530
0 11346 5 1 1 11345
0 11347 7 1 2 77570 78211
0 11348 5 1 1 11347
0 11349 7 1 2 11346 11348
0 11350 5 1 1 11349
0 11351 7 1 2 68802 11350
0 11352 5 1 1 11351
0 11353 7 4 2 72528 75941
0 11354 7 1 2 85247 89816
0 11355 5 1 1 11354
0 11356 7 1 2 11352 11355
0 11357 5 1 1 11356
0 11358 7 1 2 69988 71424
0 11359 7 1 2 11357 11358
0 11360 5 1 1 11359
0 11361 7 1 2 11344 11360
0 11362 5 1 1 11361
0 11363 7 1 2 81550 11362
0 11364 5 1 1 11363
0 11365 7 1 2 11330 11364
0 11366 5 1 1 11365
0 11367 7 1 2 66904 11366
0 11368 5 1 1 11367
0 11369 7 4 2 70877 71156
0 11370 7 2 2 77328 89820
0 11371 7 4 2 70991 89636
0 11372 7 1 2 62350 89826
0 11373 7 1 2 89824 11372
0 11374 5 1 1 11373
0 11375 7 1 2 72119 71477
0 11376 5 1 1 11375
0 11377 7 1 2 68950 89435
0 11378 5 1 1 11377
0 11379 7 1 2 11376 11378
0 11380 5 2 1 11379
0 11381 7 1 2 77373 85515
0 11382 7 1 2 89830 11381
0 11383 5 1 1 11382
0 11384 7 1 2 11374 11383
0 11385 5 1 1 11384
0 11386 7 1 2 75942 11385
0 11387 5 1 1 11386
0 11388 7 2 2 76964 73298
0 11389 5 1 1 89832
0 11390 7 1 2 78838 77144
0 11391 7 1 2 77026 11390
0 11392 7 1 2 89833 11391
0 11393 5 1 1 11392
0 11394 7 1 2 11387 11393
0 11395 5 1 1 11394
0 11396 7 1 2 81551 11395
0 11397 5 1 1 11396
0 11398 7 1 2 11368 11397
0 11399 5 1 1 11398
0 11400 7 1 2 84070 11399
0 11401 5 1 1 11400
0 11402 7 1 2 87638 88551
0 11403 5 1 1 11402
0 11404 7 1 2 61802 82417
0 11405 7 1 2 73275 11404
0 11406 5 1 1 11405
0 11407 7 1 2 11403 11406
0 11408 5 1 1 11407
0 11409 7 1 2 62351 11408
0 11410 5 1 1 11409
0 11411 7 1 2 74686 73879
0 11412 5 1 1 11411
0 11413 7 1 2 72235 11412
0 11414 5 1 1 11413
0 11415 7 2 2 65956 89691
0 11416 7 1 2 74068 89834
0 11417 5 1 1 11416
0 11418 7 1 2 75078 11417
0 11419 5 1 1 11418
0 11420 7 1 2 67188 11419
0 11421 5 1 1 11420
0 11422 7 1 2 11414 11421
0 11423 5 1 1 11422
0 11424 7 1 2 83096 11423
0 11425 5 1 1 11424
0 11426 7 1 2 11410 11425
0 11427 5 1 1 11426
0 11428 7 1 2 69749 11427
0 11429 5 1 1 11428
0 11430 7 3 2 87639 71046
0 11431 7 1 2 86599 89836
0 11432 5 1 1 11431
0 11433 7 1 2 67189 87193
0 11434 7 1 2 89835 11433
0 11435 5 1 1 11434
0 11436 7 1 2 11432 11435
0 11437 7 1 2 11429 11436
0 11438 5 1 1 11437
0 11439 7 1 2 70274 11438
0 11440 5 1 1 11439
0 11441 7 1 2 79708 72429
0 11442 5 1 1 11441
0 11443 7 1 2 85354 81161
0 11444 7 1 2 77425 11443
0 11445 5 1 1 11444
0 11446 7 1 2 11442 11445
0 11447 5 1 1 11446
0 11448 7 1 2 87305 11447
0 11449 5 1 1 11448
0 11450 7 3 2 86600 73194
0 11451 5 1 1 89839
0 11452 7 1 2 89837 89840
0 11453 5 1 1 11452
0 11454 7 1 2 11449 11453
0 11455 7 1 2 11440 11454
0 11456 5 1 1 11455
0 11457 7 1 2 83798 11456
0 11458 5 1 1 11457
0 11459 7 2 2 62039 77763
0 11460 5 1 1 89842
0 11461 7 2 2 62791 77417
0 11462 5 3 1 89844
0 11463 7 1 2 89846 78383
0 11464 5 1 1 11463
0 11465 7 1 2 62040 11464
0 11466 5 1 1 11465
0 11467 7 1 2 72932 89119
0 11468 7 1 2 79402 11467
0 11469 5 1 1 11468
0 11470 7 1 2 11466 11469
0 11471 5 1 1 11470
0 11472 7 1 2 64088 11471
0 11473 5 1 1 11472
0 11474 7 1 2 11460 11473
0 11475 5 1 1 11474
0 11476 7 1 2 68592 11475
0 11477 5 1 1 11476
0 11478 7 1 2 74477 89655
0 11479 5 1 1 11478
0 11480 7 1 2 63743 11479
0 11481 5 1 1 11480
0 11482 7 1 2 72333 75234
0 11483 5 1 1 11482
0 11484 7 1 2 11481 11483
0 11485 5 1 1 11484
0 11486 7 1 2 67190 11485
0 11487 5 1 1 11486
0 11488 7 1 2 11477 11487
0 11489 5 1 1 11488
0 11490 7 1 2 83799 83097
0 11491 7 1 2 11489 11490
0 11492 5 1 1 11491
0 11493 7 1 2 75523 79953
0 11494 7 3 2 84817 11493
0 11495 5 1 1 89849
0 11496 7 1 2 61803 89850
0 11497 5 1 1 11496
0 11498 7 4 2 70643 83098
0 11499 7 1 2 62792 79874
0 11500 7 1 2 89852 11499
0 11501 5 1 1 11500
0 11502 7 1 2 11497 11501
0 11503 5 1 1 11502
0 11504 7 1 2 83800 11503
0 11505 5 1 1 11504
0 11506 7 4 2 68803 85892
0 11507 7 1 2 82798 89856
0 11508 7 1 2 84997 11507
0 11509 5 1 1 11508
0 11510 7 1 2 11505 11509
0 11511 5 1 1 11510
0 11512 7 1 2 77899 11511
0 11513 5 1 1 11512
0 11514 7 1 2 69750 11513
0 11515 7 1 2 11492 11514
0 11516 5 1 1 11515
0 11517 7 1 2 88718 79875
0 11518 5 1 1 11517
0 11519 7 2 2 66661 74217
0 11520 7 2 2 85893 84711
0 11521 7 1 2 89860 89862
0 11522 5 1 1 11521
0 11523 7 1 2 11518 11522
0 11524 5 1 1 11523
0 11525 7 1 2 68593 11524
0 11526 5 1 1 11525
0 11527 7 4 2 67191 82656
0 11528 7 1 2 86029 77713
0 11529 7 1 2 89864 11528
0 11530 5 1 1 11529
0 11531 7 1 2 11526 11530
0 11532 5 1 1 11531
0 11533 7 1 2 62793 11532
0 11534 5 1 1 11533
0 11535 7 1 2 62352 75562
0 11536 7 1 2 85217 11535
0 11537 5 1 1 11536
0 11538 7 3 2 63102 84454
0 11539 7 1 2 74835 86030
0 11540 7 1 2 85248 11539
0 11541 7 1 2 89868 11540
0 11542 7 1 2 11537 11541
0 11543 5 1 1 11542
0 11544 7 1 2 11534 11543
0 11545 5 1 1 11544
0 11546 7 1 2 70644 11545
0 11547 5 1 1 11546
0 11548 7 2 2 88766 84527
0 11549 7 1 2 89871 82300
0 11550 5 1 1 11549
0 11551 7 1 2 64893 11550
0 11552 7 1 2 11547 11551
0 11553 5 1 1 11552
0 11554 7 1 2 65361 11553
0 11555 7 1 2 11516 11554
0 11556 5 1 1 11555
0 11557 7 1 2 89017 75384
0 11558 5 1 1 11557
0 11559 7 3 2 79818 79473
0 11560 7 2 2 82600 81512
0 11561 7 1 2 89873 89876
0 11562 5 1 1 11561
0 11563 7 1 2 11558 11562
0 11564 5 1 1 11563
0 11565 7 1 2 83099 11564
0 11566 5 1 1 11565
0 11567 7 5 2 66662 71207
0 11568 7 2 2 69751 89878
0 11569 7 1 2 88806 82070
0 11570 7 1 2 89883 11569
0 11571 5 1 1 11570
0 11572 7 1 2 11566 11571
0 11573 5 1 1 11572
0 11574 7 1 2 65362 11573
0 11575 5 1 1 11574
0 11576 7 1 2 71425 89127
0 11577 7 1 2 85621 11576
0 11578 5 1 1 11577
0 11579 7 1 2 11575 11578
0 11580 5 1 1 11579
0 11581 7 1 2 72120 11580
0 11582 5 1 1 11581
0 11583 7 1 2 69989 11582
0 11584 7 1 2 11556 11583
0 11585 7 1 2 11458 11584
0 11586 5 1 1 11585
0 11587 7 6 2 83801 81407
0 11588 7 1 2 66905 89748
0 11589 5 1 1 11588
0 11590 7 6 2 72529 72369
0 11591 7 1 2 73805 89891
0 11592 5 1 1 11591
0 11593 7 1 2 11589 11592
0 11594 5 1 1 11593
0 11595 7 1 2 67192 11594
0 11596 5 1 1 11595
0 11597 7 1 2 81139 84194
0 11598 5 1 1 11597
0 11599 7 1 2 11596 11598
0 11600 5 1 1 11599
0 11601 7 1 2 61804 11600
0 11602 5 1 1 11601
0 11603 7 2 2 70275 77622
0 11604 5 1 1 89897
0 11605 7 1 2 66906 11604
0 11606 5 1 1 11605
0 11607 7 1 2 71920 86556
0 11608 5 5 1 11607
0 11609 7 1 2 85501 76520
0 11610 7 1 2 89899 11609
0 11611 7 1 2 11606 11610
0 11612 5 1 1 11611
0 11613 7 1 2 11602 11612
0 11614 5 1 1 11613
0 11615 7 1 2 89885 11614
0 11616 5 1 1 11615
0 11617 7 1 2 66663 88703
0 11618 7 4 2 64894 72267
0 11619 7 1 2 89904 84175
0 11620 7 1 2 11617 11619
0 11621 7 1 2 89900 11620
0 11622 5 1 1 11621
0 11623 7 1 2 65099 11622
0 11624 7 1 2 11616 11623
0 11625 5 1 1 11624
0 11626 7 1 2 63513 11625
0 11627 7 1 2 11586 11626
0 11628 5 1 1 11627
0 11629 7 1 2 66403 11628
0 11630 7 1 2 11401 11629
0 11631 7 1 2 11262 11630
0 11632 5 1 1 11631
0 11633 7 1 2 69528 11632
0 11634 7 1 2 11099 11633
0 11635 5 1 1 11634
0 11636 7 2 2 66404 84528
0 11637 7 1 2 75644 89908
0 11638 5 1 1 11637
0 11639 7 11 2 66907 68118
0 11640 7 1 2 86757 89910
0 11641 7 1 2 86719 11640
0 11642 5 1 1 11641
0 11643 7 1 2 11638 11642
0 11644 5 1 1 11643
0 11645 7 1 2 67398 11644
0 11646 5 1 1 11645
0 11647 7 5 2 62353 70645
0 11648 5 1 1 89921
0 11649 7 1 2 89922 79978
0 11650 5 1 1 11649
0 11651 7 1 2 347 11650
0 11652 5 1 1 11651
0 11653 7 1 2 85418 73299
0 11654 7 1 2 11652 11653
0 11655 5 1 1 11654
0 11656 7 1 2 11646 11655
0 11657 5 1 1 11656
0 11658 7 1 2 69752 11657
0 11659 5 1 1 11658
0 11660 7 1 2 88792 73792
0 11661 5 1 1 11660
0 11662 7 1 2 68951 89851
0 11663 5 1 1 11662
0 11664 7 1 2 11661 11663
0 11665 5 1 1 11664
0 11666 7 1 2 76585 11665
0 11667 5 1 1 11666
0 11668 7 1 2 11659 11667
0 11669 5 1 1 11668
0 11670 7 1 2 66664 11669
0 11671 5 1 1 11670
0 11672 7 1 2 77769 89612
0 11673 5 2 1 11672
0 11674 7 1 2 62041 89926
0 11675 5 1 1 11674
0 11676 7 1 2 89628 11675
0 11677 5 1 1 11676
0 11678 7 1 2 85419 11677
0 11679 5 1 1 11678
0 11680 7 1 2 68119 88635
0 11681 7 1 2 79954 11680
0 11682 7 1 2 84657 11681
0 11683 5 1 1 11682
0 11684 7 1 2 11679 11683
0 11685 5 1 1 11684
0 11686 7 1 2 71047 11685
0 11687 5 1 1 11686
0 11688 7 1 2 11671 11687
0 11689 5 1 1 11688
0 11690 7 1 2 68594 11689
0 11691 5 1 1 11690
0 11692 7 14 2 63744 63922
0 11693 5 1 1 89928
0 11694 7 1 2 89238 89929
0 11695 5 1 1 11694
0 11696 7 6 2 70878 73405
0 11697 5 6 1 89942
0 11698 7 4 2 69753 75474
0 11699 5 1 1 89954
0 11700 7 1 2 89943 89955
0 11701 5 1 1 11700
0 11702 7 1 2 11695 11701
0 11703 5 1 1 11702
0 11704 7 1 2 70646 11703
0 11705 5 1 1 11704
0 11706 7 1 2 77004 80269
0 11707 5 1 1 11706
0 11708 7 1 2 11705 11707
0 11709 5 1 1 11708
0 11710 7 1 2 64089 11709
0 11711 5 1 1 11710
0 11712 7 1 2 72914 72430
0 11713 5 1 1 11712
0 11714 7 1 2 74478 11713
0 11715 5 1 1 11714
0 11716 7 1 2 64895 88279
0 11717 7 1 2 11715 11716
0 11718 5 1 1 11717
0 11719 7 1 2 11711 11718
0 11720 5 1 1 11719
0 11721 7 2 2 67193 85420
0 11722 7 1 2 11720 89958
0 11723 5 1 1 11722
0 11724 7 1 2 11691 11723
0 11725 5 1 1 11724
0 11726 7 1 2 67970 11725
0 11727 5 1 1 11726
0 11728 7 1 2 85228 85009
0 11729 5 1 1 11728
0 11730 7 1 2 11495 11729
0 11731 5 1 1 11730
0 11732 7 1 2 66665 11731
0 11733 5 1 1 11732
0 11734 7 2 2 83039 79955
0 11735 7 1 2 85746 89960
0 11736 5 1 1 11735
0 11737 7 1 2 11733 11736
0 11738 5 1 1 11737
0 11739 7 1 2 68952 11738
0 11740 5 1 1 11739
0 11741 7 1 2 67644 84712
0 11742 7 1 2 75865 11741
0 11743 5 1 1 11742
0 11744 7 1 2 11740 11743
0 11745 5 1 1 11744
0 11746 7 1 2 76071 86159
0 11747 7 1 2 11745 11746
0 11748 5 1 1 11747
0 11749 7 1 2 11727 11748
0 11750 5 1 1 11749
0 11751 7 1 2 65363 11750
0 11752 5 1 1 11751
0 11753 7 1 2 77739 1522
0 11754 5 1 1 11753
0 11755 7 1 2 11754 77711
0 11756 5 1 1 11755
0 11757 7 1 2 70647 11756
0 11758 5 1 1 11757
0 11759 7 2 2 62354 68804
0 11760 5 1 1 89962
0 11761 7 1 2 77697 89963
0 11762 5 1 1 11761
0 11763 7 1 2 77701 11762
0 11764 7 1 2 11758 11763
0 11765 5 1 1 11764
0 11766 7 1 2 84782 11765
0 11767 5 1 1 11766
0 11768 7 2 2 62355 77598
0 11769 7 1 2 83040 77085
0 11770 7 1 2 73933 11769
0 11771 7 1 2 89964 11770
0 11772 5 1 1 11771
0 11773 7 1 2 11767 11772
0 11774 5 1 1 11773
0 11775 7 1 2 70276 11774
0 11776 5 1 1 11775
0 11777 7 1 2 71426 85472
0 11778 5 1 1 11777
0 11779 7 1 2 68805 77703
0 11780 5 1 1 11779
0 11781 7 1 2 11778 11780
0 11782 5 1 1 11781
0 11783 7 1 2 82132 75028
0 11784 7 1 2 11782 11783
0 11785 5 1 1 11784
0 11786 7 1 2 11776 11785
0 11787 5 1 1 11786
0 11788 7 1 2 72036 11787
0 11789 5 1 1 11788
0 11790 7 1 2 71427 86732
0 11791 5 1 1 11790
0 11792 7 1 2 86255 11791
0 11793 5 1 1 11792
0 11794 7 3 2 70277 84818
0 11795 7 1 2 75029 89966
0 11796 7 1 2 11793 11795
0 11797 5 1 1 11796
0 11798 7 1 2 11789 11797
0 11799 5 1 1 11798
0 11800 7 1 2 80966 11799
0 11801 5 1 1 11800
0 11802 7 1 2 11752 11801
0 11803 5 1 1 11802
0 11804 7 1 2 69327 11803
0 11805 5 1 1 11804
0 11806 7 4 2 70648 85959
0 11807 7 1 2 80275 89969
0 11808 5 1 1 11807
0 11809 7 1 2 76647 72317
0 11810 5 1 1 11809
0 11811 7 1 2 74109 74015
0 11812 5 1 1 11811
0 11813 7 1 2 11810 11812
0 11814 5 1 1 11813
0 11815 7 1 2 70879 11814
0 11816 5 1 1 11815
0 11817 7 1 2 76648 77536
0 11818 5 1 1 11817
0 11819 7 1 2 11816 11818
0 11820 5 1 1 11819
0 11821 7 1 2 63745 11820
0 11822 5 1 1 11821
0 11823 7 3 2 62042 70880
0 11824 5 1 1 89973
0 11825 7 1 2 86001 89974
0 11826 5 1 1 11825
0 11827 7 1 2 11822 11826
0 11828 5 1 1 11827
0 11829 7 1 2 65364 11828
0 11830 5 1 1 11829
0 11831 7 1 2 11808 11830
0 11832 5 1 1 11831
0 11833 7 1 2 71048 11832
0 11834 5 1 1 11833
0 11835 7 9 2 67194 70278
0 11836 5 2 1 89976
0 11837 7 1 2 89977 75909
0 11838 5 1 1 11837
0 11839 7 1 2 1242 11838
0 11840 5 1 1 11839
0 11841 7 1 2 62043 11840
0 11842 5 1 1 11841
0 11843 7 2 2 73195 77344
0 11844 5 1 1 89987
0 11845 7 1 2 87865 89988
0 11846 5 1 1 11845
0 11847 7 1 2 11842 11846
0 11848 5 1 1 11847
0 11849 7 1 2 66666 11848
0 11850 5 1 1 11849
0 11851 7 3 2 61805 74790
0 11852 7 1 2 89892 89989
0 11853 5 1 1 11852
0 11854 7 1 2 73196 77742
0 11855 5 1 1 11854
0 11856 7 1 2 11853 11855
0 11857 5 1 1 11856
0 11858 7 1 2 66908 11857
0 11859 5 1 1 11858
0 11860 7 1 2 11850 11859
0 11861 5 1 1 11860
0 11862 7 1 2 69754 11861
0 11863 5 1 1 11862
0 11864 7 1 2 11834 11863
0 11865 5 1 1 11864
0 11866 7 1 2 63284 11865
0 11867 5 1 1 11866
0 11868 7 1 2 73061 88941
0 11869 7 1 2 73806 89281
0 11870 7 1 2 11868 11869
0 11871 5 1 1 11870
0 11872 7 1 2 11867 11871
0 11873 5 1 1 11872
0 11874 7 1 2 81080 11873
0 11875 5 1 1 11874
0 11876 7 1 2 69990 11875
0 11877 7 1 2 11805 11876
0 11878 5 1 1 11877
0 11879 7 1 2 75197 89702
0 11880 5 1 1 11879
0 11881 7 1 2 79956 85098
0 11882 7 1 2 85747 11881
0 11883 5 1 1 11882
0 11884 7 1 2 11880 11883
0 11885 5 1 1 11884
0 11886 7 1 2 68953 76128
0 11887 7 1 2 11885 11886
0 11888 5 1 1 11887
0 11889 7 1 2 75943 75886
0 11890 5 2 1 11889
0 11891 7 1 2 62794 81165
0 11892 5 1 1 11891
0 11893 7 1 2 89754 87035
0 11894 7 1 2 11892 11893
0 11895 5 1 1 11894
0 11896 7 1 2 89992 11895
0 11897 5 1 1 11896
0 11898 7 1 2 70649 11897
0 11899 5 1 1 11898
0 11900 7 2 2 75218 89703
0 11901 5 1 1 89994
0 11902 7 1 2 11899 11901
0 11903 5 1 1 11902
0 11904 7 1 2 61494 78768
0 11905 7 1 2 11903 11904
0 11906 5 1 1 11905
0 11907 7 1 2 11888 11906
0 11908 5 1 1 11907
0 11909 7 1 2 68120 11908
0 11910 5 1 1 11909
0 11911 7 2 2 82133 78496
0 11912 7 2 2 73772 74920
0 11913 5 1 1 89998
0 11914 7 1 2 89999 80945
0 11915 7 1 2 89996 11914
0 11916 5 1 1 11915
0 11917 7 1 2 11910 11916
0 11918 5 1 1 11917
0 11919 7 1 2 69328 11918
0 11920 5 1 1 11919
0 11921 7 1 2 77489 82840
0 11922 7 1 2 89872 11921
0 11923 7 1 2 89901 11922
0 11924 5 1 1 11923
0 11925 7 1 2 11920 11924
0 11926 5 1 1 11925
0 11927 7 1 2 64896 11926
0 11928 5 1 1 11927
0 11929 7 12 2 61495 62356
0 11930 7 3 2 75851 90000
0 11931 7 1 2 83802 79854
0 11932 7 1 2 90012 11931
0 11933 7 1 2 89853 11932
0 11934 5 1 1 11933
0 11935 7 1 2 65100 11934
0 11936 7 1 2 11928 11935
0 11937 5 1 1 11936
0 11938 7 1 2 63514 11937
0 11939 7 1 2 11878 11938
0 11940 5 1 1 11939
0 11941 7 3 2 64897 73603
0 11942 7 1 2 85775 90015
0 11943 5 1 1 11942
0 11944 7 1 2 85705 76773
0 11945 5 1 1 11944
0 11946 7 1 2 11943 11945
0 11947 5 1 1 11946
0 11948 7 1 2 62044 11947
0 11949 5 1 1 11948
0 11950 7 1 2 66909 75249
0 11951 7 1 2 77722 11950
0 11952 7 1 2 77882 11951
0 11953 5 1 1 11952
0 11954 7 1 2 11949 11953
0 11955 5 1 1 11954
0 11956 7 1 2 66667 11955
0 11957 5 1 1 11956
0 11958 7 1 2 75404 86002
0 11959 7 1 2 90016 11958
0 11960 5 1 1 11959
0 11961 7 1 2 11957 11960
0 11962 5 1 1 11961
0 11963 7 1 2 78135 11962
0 11964 5 1 1 11963
0 11965 7 2 2 80599 84630
0 11966 7 1 2 75405 73158
0 11967 7 1 2 90018 11966
0 11968 5 1 1 11967
0 11969 7 1 2 11964 11968
0 11970 5 1 1 11969
0 11971 7 1 2 68121 11970
0 11972 5 1 1 11971
0 11973 7 1 2 66668 89195
0 11974 7 1 2 90019 11973
0 11975 5 1 1 11974
0 11976 7 1 2 11972 11975
0 11977 5 1 1 11976
0 11978 7 1 2 76129 11977
0 11979 5 1 1 11978
0 11980 7 2 2 62527 77192
0 11981 7 12 2 62357 63103
0 11982 7 1 2 90020 90022
0 11983 7 5 2 64898 78408
0 11984 7 2 2 63923 82418
0 11985 7 1 2 90034 90039
0 11986 7 1 2 11982 11985
0 11987 5 1 1 11986
0 11988 7 5 2 76039 82733
0 11989 5 1 1 90041
0 11990 7 1 2 80346 90042
0 11991 5 1 1 11990
0 11992 7 3 2 76072 83100
0 11993 5 1 1 90046
0 11994 7 1 2 64899 90047
0 11995 5 1 1 11994
0 11996 7 1 2 11991 11995
0 11997 5 1 1 11996
0 11998 7 1 2 69991 74580
0 11999 7 1 2 89527 11998
0 12000 7 1 2 11997 11999
0 12001 5 1 1 12000
0 12002 7 1 2 11987 12001
0 12003 5 1 1 12002
0 12004 7 1 2 67645 12003
0 12005 5 1 1 12004
0 12006 7 3 2 62358 78748
0 12007 7 4 2 66405 74151
0 12008 7 2 2 90049 90052
0 12009 7 2 2 68122 75250
0 12010 5 3 1 90058
0 12011 7 1 2 80753 87569
0 12012 7 1 2 90059 12011
0 12013 7 1 2 90056 12012
0 12014 5 1 1 12013
0 12015 7 1 2 12005 12014
0 12016 5 1 1 12015
0 12017 7 1 2 64090 12016
0 12018 5 1 1 12017
0 12019 7 1 2 78147 81408
0 12020 7 1 2 89861 12019
0 12021 5 1 1 12020
0 12022 7 4 2 63104 83041
0 12023 7 1 2 90035 90063
0 12024 7 1 2 75498 12023
0 12025 5 1 1 12024
0 12026 7 1 2 12021 12025
0 12027 5 1 1 12026
0 12028 7 1 2 80723 76422
0 12029 7 1 2 12027 12028
0 12030 5 1 1 12029
0 12031 7 1 2 12018 12030
0 12032 7 1 2 11979 12031
0 12033 5 1 1 12032
0 12034 7 1 2 70650 12033
0 12035 5 1 1 12034
0 12036 7 1 2 77795 77960
0 12037 5 1 1 12036
0 12038 7 1 2 86050 89927
0 12039 5 1 1 12038
0 12040 7 1 2 12037 12039
0 12041 5 1 1 12040
0 12042 7 1 2 68595 12041
0 12043 5 1 1 12042
0 12044 7 2 2 66910 77940
0 12045 5 2 1 90067
0 12046 7 1 2 87570 85355
0 12047 7 1 2 90068 12046
0 12048 5 1 1 12047
0 12049 7 1 2 12043 12048
0 12050 5 1 1 12049
0 12051 7 6 2 64900 76130
0 12052 7 1 2 88201 90071
0 12053 7 1 2 12050 12052
0 12054 5 1 1 12053
0 12055 7 1 2 12035 12054
0 12056 5 1 1 12055
0 12057 7 1 2 68354 12056
0 12058 5 1 1 12057
0 12059 7 3 2 66669 73159
0 12060 7 1 2 76586 90077
0 12061 5 1 1 12060
0 12062 7 3 2 66406 71672
0 12063 7 1 2 81982 90080
0 12064 5 1 1 12063
0 12065 7 1 2 12061 12064
0 12066 5 1 1 12065
0 12067 7 1 2 12066 89772
0 12068 5 1 1 12067
0 12069 7 7 2 69755 79602
0 12070 7 3 2 87640 76552
0 12071 7 1 2 71673 90090
0 12072 7 1 2 90083 12071
0 12073 5 1 1 12072
0 12074 7 1 2 12068 12073
0 12075 5 1 1 12074
0 12076 7 1 2 67971 12075
0 12077 5 1 1 12076
0 12078 7 2 2 67399 78691
0 12079 7 1 2 82134 76553
0 12080 7 1 2 90036 12079
0 12081 7 1 2 90093 12080
0 12082 5 1 1 12081
0 12083 7 1 2 12077 12082
0 12084 5 1 1 12083
0 12085 7 1 2 79403 73670
0 12086 7 1 2 12084 12085
0 12087 5 1 1 12086
0 12088 7 1 2 12058 12087
0 12089 5 1 1 12088
0 12090 7 1 2 69329 12089
0 12091 5 1 1 12090
0 12092 7 3 2 83452 85183
0 12093 7 1 2 87465 72318
0 12094 7 1 2 90095 12093
0 12095 5 1 1 12094
0 12096 7 1 2 61496 87641
0 12097 7 1 2 79531 12096
0 12098 7 1 2 85291 12097
0 12099 5 1 1 12098
0 12100 7 1 2 12095 12099
0 12101 5 1 1 12100
0 12102 7 1 2 65365 12101
0 12103 5 1 1 12102
0 12104 7 4 2 69330 82521
0 12105 7 1 2 78129 90096
0 12106 7 1 2 90098 12105
0 12107 5 1 1 12106
0 12108 7 1 2 12103 12107
0 12109 5 1 1 12108
0 12110 7 1 2 62045 12109
0 12111 5 1 1 12110
0 12112 7 6 2 65101 71723
0 12113 5 1 1 90102
0 12114 7 1 2 73682 90103
0 12115 5 1 1 12114
0 12116 7 1 2 69992 85688
0 12117 5 1 1 12116
0 12118 7 1 2 12115 12117
0 12119 5 1 1 12118
0 12120 7 1 2 67400 12119
0 12121 5 1 1 12120
0 12122 7 2 2 76934 74027
0 12123 5 2 1 90108
0 12124 7 1 2 12121 90110
0 12125 5 1 1 12124
0 12126 7 1 2 86301 85184
0 12127 7 1 2 82698 12126
0 12128 7 1 2 12125 12127
0 12129 5 1 1 12128
0 12130 7 1 2 12111 12129
0 12131 5 1 1 12130
0 12132 7 1 2 70881 12131
0 12133 5 1 1 12132
0 12134 7 1 2 62046 89749
0 12135 5 1 1 12134
0 12136 7 4 2 64091 73062
0 12137 5 1 1 90112
0 12138 7 1 2 77714 90113
0 12139 5 1 1 12138
0 12140 7 1 2 12135 12139
0 12141 5 1 1 12140
0 12142 7 1 2 65102 12141
0 12143 5 1 1 12142
0 12144 7 10 2 66911 64092
0 12145 7 1 2 90116 85056
0 12146 5 1 1 12145
0 12147 7 1 2 12143 12146
0 12148 5 1 1 12147
0 12149 7 1 2 67646 12148
0 12150 5 1 1 12149
0 12151 7 1 2 77715 78409
0 12152 5 1 1 12151
0 12153 7 1 2 85051 81197
0 12154 5 1 1 12153
0 12155 7 1 2 12152 12154
0 12156 5 1 1 12155
0 12157 7 1 2 62795 72420
0 12158 7 1 2 12156 12157
0 12159 5 1 1 12158
0 12160 7 1 2 12150 12159
0 12161 5 1 1 12160
0 12162 7 1 2 86867 83453
0 12163 7 1 2 12161 12162
0 12164 5 1 1 12163
0 12165 7 1 2 12133 12164
0 12166 5 1 1 12165
0 12167 7 1 2 61806 12166
0 12168 5 1 1 12167
0 12169 7 1 2 65366 89301
0 12170 7 3 2 89643 12169
0 12171 5 1 1 90126
0 12172 7 1 2 80872 81838
0 12173 7 1 2 90127 12172
0 12174 5 1 1 12173
0 12175 7 2 2 11309 4385
0 12176 5 1 1 90129
0 12177 7 1 2 62796 90130
0 12178 5 1 1 12177
0 12179 7 2 2 70651 72319
0 12180 5 1 1 90131
0 12181 7 1 2 67647 78220
0 12182 7 1 2 12180 12181
0 12183 5 1 1 12182
0 12184 7 1 2 88580 12183
0 12185 7 1 2 12178 12184
0 12186 5 1 1 12185
0 12187 7 1 2 12174 12186
0 12188 5 1 1 12187
0 12189 7 1 2 67401 12188
0 12190 5 1 1 12189
0 12191 7 6 2 68596 74615
0 12192 7 2 2 74069 88636
0 12193 7 1 2 89105 90139
0 12194 7 1 2 90133 12193
0 12195 5 1 1 12194
0 12196 7 1 2 12190 12195
0 12197 5 1 1 12196
0 12198 7 1 2 85724 79733
0 12199 7 1 2 12197 12198
0 12200 5 1 1 12199
0 12201 7 1 2 12168 12200
0 12202 5 1 1 12201
0 12203 7 1 2 64901 12202
0 12204 5 1 1 12203
0 12205 7 1 2 75406 90128
0 12206 5 1 1 12205
0 12207 7 1 2 75475 77027
0 12208 5 1 1 12207
0 12209 7 1 2 12206 12208
0 12210 5 1 1 12209
0 12211 7 1 2 68597 12210
0 12212 5 1 1 12211
0 12213 7 3 2 70279 86720
0 12214 5 1 1 90141
0 12215 7 1 2 84034 12214
0 12216 5 1 1 12215
0 12217 7 1 2 75476 12216
0 12218 5 1 1 12217
0 12219 7 1 2 12212 12218
0 12220 5 1 1 12219
0 12221 7 1 2 67402 12220
0 12222 5 1 1 12221
0 12223 7 1 2 62047 84631
0 12224 5 1 1 12223
0 12225 7 1 2 83609 12224
0 12226 5 1 1 12225
0 12227 7 2 2 74177 87449
0 12228 7 1 2 12226 90144
0 12229 5 1 1 12228
0 12230 7 1 2 79819 75700
0 12231 7 1 2 89893 12230
0 12232 5 1 1 12231
0 12233 7 1 2 12229 12232
0 12234 7 1 2 12222 12233
0 12235 5 1 1 12234
0 12236 7 2 2 87466 85639
0 12237 7 1 2 12235 90146
0 12238 5 1 1 12237
0 12239 7 1 2 87086 82247
0 12240 7 1 2 87505 12239
0 12241 5 1 1 12240
0 12242 7 1 2 12238 12241
0 12243 5 1 1 12242
0 12244 7 1 2 75053 12243
0 12245 5 1 1 12244
0 12246 7 1 2 12204 12245
0 12247 5 1 1 12246
0 12248 7 1 2 63105 12247
0 12249 5 1 1 12248
0 12250 7 4 2 61497 65103
0 12251 7 1 2 90148 85143
0 12252 7 1 2 89799 12251
0 12253 5 1 1 12252
0 12254 7 2 2 61498 89740
0 12255 5 1 1 90152
0 12256 7 2 2 70280 88581
0 12257 5 1 1 90154
0 12258 7 1 2 12255 12257
0 12259 5 1 1 12258
0 12260 7 1 2 75407 85837
0 12261 7 1 2 12259 12260
0 12262 5 1 1 12261
0 12263 7 1 2 12253 12262
0 12264 5 1 1 12263
0 12265 7 1 2 73406 12264
0 12266 5 1 1 12265
0 12267 7 1 2 74581 81032
0 12268 5 1 1 12267
0 12269 7 1 2 12268 1902
0 12270 5 1 1 12269
0 12271 7 1 2 90145 12270
0 12272 5 1 1 12271
0 12273 7 1 2 75944 75408
0 12274 5 2 1 12273
0 12275 7 1 2 11211 90156
0 12276 5 1 1 12275
0 12277 7 1 2 72121 12276
0 12278 5 1 1 12277
0 12279 7 1 2 12278 89993
0 12280 5 1 1 12279
0 12281 7 1 2 65104 12280
0 12282 5 1 1 12281
0 12283 7 1 2 73773 84447
0 12284 7 1 2 88552 12283
0 12285 5 1 1 12284
0 12286 7 1 2 12282 12285
0 12287 5 1 1 12286
0 12288 7 1 2 71208 12287
0 12289 5 1 1 12288
0 12290 7 1 2 12272 12289
0 12291 5 1 1 12290
0 12292 7 1 2 81839 12291
0 12293 5 1 1 12292
0 12294 7 1 2 12266 12293
0 12295 5 1 1 12294
0 12296 7 1 2 69756 12295
0 12297 5 1 1 12296
0 12298 7 1 2 78654 83176
0 12299 7 1 2 12176 12298
0 12300 5 1 1 12299
0 12301 7 1 2 75976 4804
0 12302 5 1 1 12301
0 12303 7 3 2 68123 74152
0 12304 7 1 2 79621 90158
0 12305 7 1 2 12302 12304
0 12306 5 1 1 12305
0 12307 7 1 2 12300 12306
0 12308 5 1 1 12307
0 12309 7 1 2 62797 12308
0 12310 5 1 1 12309
0 12311 7 1 2 66912 78234
0 12312 5 1 1 12311
0 12313 7 1 2 85875 80270
0 12314 5 1 1 12313
0 12315 7 1 2 12312 12314
0 12316 5 1 1 12315
0 12317 7 1 2 83042 12316
0 12318 5 1 1 12317
0 12319 7 1 2 78667 83230
0 12320 5 1 1 12319
0 12321 7 1 2 12318 12320
0 12322 5 1 1 12321
0 12323 7 1 2 72408 12322
0 12324 5 1 1 12323
0 12325 7 1 2 12310 12324
0 12326 5 1 1 12325
0 12327 7 1 2 76587 12326
0 12328 5 1 1 12327
0 12329 7 1 2 12297 12328
0 12330 5 1 1 12329
0 12331 7 1 2 68355 12330
0 12332 5 1 1 12331
0 12333 7 1 2 78600 80067
0 12334 7 1 2 73197 86567
0 12335 7 1 2 12333 12334
0 12336 7 2 2 66407 75409
0 12337 7 1 2 90161 75227
0 12338 7 1 2 12335 12337
0 12339 5 1 1 12338
0 12340 7 1 2 12332 12339
0 12341 5 1 1 12340
0 12342 7 1 2 84071 12341
0 12343 5 1 1 12342
0 12344 7 1 2 12249 12343
0 12345 5 1 1 12344
0 12346 7 1 2 67195 12345
0 12347 5 1 1 12346
0 12348 7 2 2 63106 74028
0 12349 7 1 2 82248 90163
0 12350 7 2 2 78545 87490
0 12351 7 2 2 62359 74153
0 12352 7 1 2 90165 90167
0 12353 7 1 2 12349 12352
0 12354 5 1 1 12353
0 12355 7 1 2 12347 12354
0 12356 7 1 2 12091 12355
0 12357 7 1 2 11940 12356
0 12358 5 1 1 12357
0 12359 7 1 2 64675 12358
0 12360 5 1 1 12359
0 12361 7 6 2 61807 81727
0 12362 5 2 1 90169
0 12363 7 4 2 66670 81752
0 12364 5 2 1 90177
0 12365 7 1 2 90175 90181
0 12366 5 36 1 12365
0 12367 7 5 2 62360 69529
0 12368 7 2 2 82841 90219
0 12369 7 1 2 82476 90224
0 12370 5 1 1 12369
0 12371 7 3 2 65105 77964
0 12372 7 1 2 83393 84400
0 12373 7 1 2 90226 12372
0 12374 5 1 1 12373
0 12375 7 1 2 12370 12374
0 12376 5 1 1 12375
0 12377 7 1 2 70281 77086
0 12378 7 1 2 12376 12377
0 12379 5 1 1 12378
0 12380 7 1 2 63515 85459
0 12381 5 1 1 12380
0 12382 7 1 2 87978 12381
0 12383 5 1 1 12382
0 12384 7 1 2 68356 85463
0 12385 5 1 1 12384
0 12386 7 1 2 12383 12385
0 12387 5 1 1 12386
0 12388 7 20 2 61499 66913
0 12389 7 1 2 83659 90229
0 12390 7 1 2 12387 12389
0 12391 5 1 1 12390
0 12392 7 1 2 12379 12391
0 12393 5 1 1 12392
0 12394 7 1 2 62798 12393
0 12395 5 1 1 12394
0 12396 7 1 2 62528 79049
0 12397 5 2 1 12396
0 12398 7 1 2 2111 90249
0 12399 5 1 1 12398
0 12400 7 1 2 79308 83737
0 12401 5 1 1 12400
0 12402 7 1 2 62361 12401
0 12403 5 1 1 12402
0 12404 7 1 2 79118 88802
0 12405 7 1 2 12403 12404
0 12406 7 1 2 12399 12405
0 12407 5 1 1 12406
0 12408 7 1 2 12395 12407
0 12409 5 1 1 12408
0 12410 7 1 2 70882 12409
0 12411 5 1 1 12410
0 12412 7 2 2 62362 73115
0 12413 5 1 1 90251
0 12414 7 1 2 73198 89978
0 12415 5 2 1 12414
0 12416 7 1 2 12413 90253
0 12417 5 1 1 12416
0 12418 7 30 2 66408 79428
0 12419 5 1 1 90255
0 12420 7 2 2 77087 90256
0 12421 7 2 2 62529 90285
0 12422 7 1 2 12417 90287
0 12423 5 1 1 12422
0 12424 7 3 2 68357 90230
0 12425 7 3 2 83983 90289
0 12426 7 1 2 83738 71568
0 12427 7 1 2 90292 12426
0 12428 5 2 1 12427
0 12429 7 1 2 12423 90295
0 12430 5 1 1 12429
0 12431 7 1 2 81026 12430
0 12432 5 1 1 12431
0 12433 7 1 2 12411 12432
0 12434 5 1 1 12433
0 12435 7 1 2 64093 12434
0 12436 5 1 1 12435
0 12437 7 2 2 76315 80292
0 12438 7 1 2 78016 90297
0 12439 5 1 1 12438
0 12440 7 3 2 77394 84159
0 12441 5 1 1 90299
0 12442 7 1 2 12439 12441
0 12443 5 1 1 12442
0 12444 7 1 2 62363 12443
0 12445 5 1 1 12444
0 12446 7 1 2 71569 4299
0 12447 5 2 1 12446
0 12448 7 1 2 66914 84169
0 12449 7 1 2 85061 12448
0 12450 5 1 1 12449
0 12451 7 1 2 5158 12450
0 12452 5 2 1 12451
0 12453 7 1 2 90302 90304
0 12454 5 1 1 12453
0 12455 7 1 2 67196 73116
0 12456 5 1 1 12455
0 12457 7 1 2 75925 12456
0 12458 5 1 1 12457
0 12459 7 1 2 75524 12458
0 12460 5 1 1 12459
0 12461 7 1 2 72478 87967
0 12462 5 1 1 12461
0 12463 7 1 2 68358 12462
0 12464 5 1 1 12463
0 12465 7 1 2 12460 12464
0 12466 5 1 1 12465
0 12467 7 1 2 67403 12466
0 12468 5 1 1 12467
0 12469 7 1 2 73252 76497
0 12470 5 4 1 12469
0 12471 7 1 2 84160 90306
0 12472 5 1 1 12471
0 12473 7 1 2 12468 12472
0 12474 5 1 1 12473
0 12475 7 1 2 66915 12474
0 12476 5 1 1 12475
0 12477 7 1 2 12454 12476
0 12478 5 1 1 12477
0 12479 7 1 2 69757 12478
0 12480 5 1 1 12479
0 12481 7 1 2 12445 12480
0 12482 5 1 1 12481
0 12483 7 1 2 83949 12482
0 12484 5 1 1 12483
0 12485 7 7 2 69331 84401
0 12486 7 1 2 62799 80314
0 12487 5 1 1 12486
0 12488 7 8 2 67404 65367
0 12489 5 2 1 90317
0 12490 7 2 2 73253 90318
0 12491 5 1 1 90327
0 12492 7 1 2 69758 75088
0 12493 7 1 2 90328 12492
0 12494 5 1 1 12493
0 12495 7 1 2 12487 12494
0 12496 5 1 1 12495
0 12497 7 1 2 67197 12496
0 12498 5 1 1 12497
0 12499 7 1 2 75852 75621
0 12500 7 1 2 90252 12499
0 12501 5 1 1 12500
0 12502 7 1 2 12498 12501
0 12503 5 1 1 12502
0 12504 7 1 2 90310 12503
0 12505 5 1 1 12504
0 12506 7 1 2 12484 12505
0 12507 5 1 1 12506
0 12508 7 1 2 68954 12507
0 12509 5 1 1 12508
0 12510 7 1 2 68806 90305
0 12511 5 1 1 12510
0 12512 7 2 2 77469 72846
0 12513 5 1 1 90329
0 12514 7 1 2 12511 12513
0 12515 5 1 1 12514
0 12516 7 1 2 65697 12515
0 12517 5 1 1 12516
0 12518 7 1 2 86601 84161
0 12519 5 1 1 12518
0 12520 7 1 2 12517 12519
0 12521 5 1 1 12520
0 12522 7 2 2 73574 83950
0 12523 5 1 1 90331
0 12524 7 1 2 12521 90332
0 12525 5 1 1 12524
0 12526 7 1 2 74191 77571
0 12527 7 1 2 90257 12526
0 12528 7 2 2 65368 75089
0 12529 7 2 2 63924 76334
0 12530 5 2 1 90335
0 12531 7 1 2 90333 90337
0 12532 7 1 2 12527 12531
0 12533 5 1 1 12532
0 12534 7 1 2 12525 12533
0 12535 5 1 1 12534
0 12536 7 1 2 69759 12535
0 12537 5 1 1 12536
0 12538 7 1 2 12509 12537
0 12539 5 1 1 12538
0 12540 7 1 2 69993 12539
0 12541 5 1 1 12540
0 12542 7 1 2 12436 12541
0 12543 5 1 1 12542
0 12544 7 1 2 68598 12543
0 12545 5 1 1 12544
0 12546 7 1 2 89985 86395
0 12547 5 16 1 12546
0 12548 7 1 2 71157 80692
0 12549 7 1 2 90339 12548
0 12550 5 1 1 12549
0 12551 7 3 2 74616 75286
0 12552 7 1 2 62364 74431
0 12553 7 1 2 90355 12552
0 12554 5 1 1 12553
0 12555 7 1 2 12550 12554
0 12556 5 1 1 12555
0 12557 7 1 2 63746 12556
0 12558 5 1 1 12557
0 12559 7 1 2 85400 86442
0 12560 5 2 1 12559
0 12561 7 1 2 77295 90358
0 12562 5 1 1 12561
0 12563 7 1 2 12558 12562
0 12564 5 1 1 12563
0 12565 7 1 2 77088 12564
0 12566 5 1 1 12565
0 12567 7 2 2 78601 86792
0 12568 7 1 2 79709 71014
0 12569 7 1 2 90360 12568
0 12570 5 1 1 12569
0 12571 7 1 2 12566 12570
0 12572 5 1 1 12571
0 12573 7 1 2 90258 12572
0 12574 5 1 1 12573
0 12575 7 1 2 85825 90340
0 12576 5 1 1 12575
0 12577 7 1 2 77296 86391
0 12578 5 1 1 12577
0 12579 7 1 2 12576 12578
0 12580 5 1 1 12579
0 12581 7 1 2 63747 12580
0 12582 5 1 1 12581
0 12583 7 1 2 88755 74652
0 12584 5 1 1 12583
0 12585 7 1 2 12582 12584
0 12586 5 1 1 12585
0 12587 7 2 2 86670 79072
0 12588 7 1 2 87516 90362
0 12589 7 1 2 12586 12588
0 12590 5 1 1 12589
0 12591 7 1 2 12574 12590
0 12592 5 1 1 12591
0 12593 7 1 2 62530 12592
0 12594 5 1 1 12593
0 12595 7 1 2 84316 90300
0 12596 5 1 1 12595
0 12597 7 2 2 73544 75303
0 12598 5 1 1 90364
0 12599 7 1 2 64902 90341
0 12600 7 1 2 90365 12599
0 12601 5 1 1 12600
0 12602 7 1 2 12596 12601
0 12603 5 1 1 12602
0 12604 7 1 2 63748 12603
0 12605 5 1 1 12604
0 12606 7 1 2 62800 85512
0 12607 5 1 1 12606
0 12608 7 1 2 74725 12607
0 12609 5 1 1 12608
0 12610 7 2 2 67405 12609
0 12611 5 1 1 90366
0 12612 7 2 2 70282 84317
0 12613 5 1 1 90368
0 12614 7 1 2 67198 90369
0 12615 5 1 1 12614
0 12616 7 1 2 12611 12615
0 12617 5 1 1 12616
0 12618 7 1 2 88037 12617
0 12619 5 1 1 12618
0 12620 7 1 2 12605 12619
0 12621 5 1 1 12620
0 12622 7 1 2 68807 12621
0 12623 5 1 1 12622
0 12624 7 1 2 74001 89986
0 12625 5 10 1 12624
0 12626 7 2 2 74999 6582
0 12627 5 1 1 90380
0 12628 7 1 2 90370 90381
0 12629 5 1 1 12628
0 12630 7 1 2 84301 85028
0 12631 5 1 1 12630
0 12632 7 1 2 12629 12631
0 12633 5 1 1 12632
0 12634 7 1 2 88038 12633
0 12635 5 1 1 12634
0 12636 7 1 2 12623 12635
0 12637 5 1 1 12636
0 12638 7 1 2 61500 81568
0 12639 7 1 2 12637 12638
0 12640 5 1 1 12639
0 12641 7 1 2 12594 12640
0 12642 5 1 1 12641
0 12643 7 1 2 65698 12642
0 12644 5 1 1 12643
0 12645 7 2 2 67199 74750
0 12646 5 1 1 90382
0 12647 7 1 2 73984 85838
0 12648 5 2 1 12647
0 12649 7 1 2 12646 90384
0 12650 5 1 1 12649
0 12651 7 1 2 73407 12650
0 12652 5 1 1 12651
0 12653 7 1 2 72940 89731
0 12654 5 1 1 12653
0 12655 7 1 2 12652 12654
0 12656 5 1 1 12655
0 12657 7 1 2 83951 12656
0 12658 5 1 1 12657
0 12659 7 4 2 70883 86302
0 12660 7 2 2 80927 80320
0 12661 7 1 2 90386 90390
0 12662 7 1 2 85509 12661
0 12663 5 1 1 12662
0 12664 7 1 2 12658 12663
0 12665 5 1 1 12664
0 12666 7 1 2 69994 12665
0 12667 5 1 1 12666
0 12668 7 2 2 63749 86303
0 12669 7 1 2 79747 80928
0 12670 7 1 2 74198 12669
0 12671 7 1 2 90392 12670
0 12672 5 1 1 12671
0 12673 7 1 2 12667 12672
0 12674 5 1 1 12673
0 12675 7 1 2 75054 12674
0 12676 5 1 1 12675
0 12677 7 1 2 76649 77135
0 12678 7 2 2 80470 84557
0 12679 7 1 2 83246 90394
0 12680 7 1 2 12677 12679
0 12681 5 1 1 12680
0 12682 7 1 2 12676 12681
0 12683 5 1 1 12682
0 12684 7 1 2 66916 12683
0 12685 5 1 1 12684
0 12686 7 1 2 78655 80625
0 12687 7 1 2 77558 12686
0 12688 7 1 2 89410 12687
0 12689 5 1 1 12688
0 12690 7 1 2 73300 83556
0 12691 7 1 2 80511 12690
0 12692 7 1 2 80882 12691
0 12693 5 1 1 12692
0 12694 7 1 2 12689 12693
0 12695 5 1 1 12694
0 12696 7 1 2 69995 12695
0 12697 5 1 1 12696
0 12698 7 2 2 79638 87444
0 12699 7 2 2 73301 79248
0 12700 7 1 2 90396 90398
0 12701 5 1 1 12700
0 12702 7 1 2 12697 12701
0 12703 5 1 1 12702
0 12704 7 1 2 70652 12703
0 12705 5 1 1 12704
0 12706 7 2 2 62365 73712
0 12707 7 1 2 83557 79249
0 12708 7 1 2 85901 12707
0 12709 7 1 2 90400 12708
0 12710 5 1 1 12709
0 12711 7 1 2 12705 12710
0 12712 5 1 1 12711
0 12713 7 1 2 71158 12712
0 12714 5 1 1 12713
0 12715 7 1 2 12685 12714
0 12716 7 1 2 12644 12715
0 12717 7 1 2 12545 12716
0 12718 5 1 1 12717
0 12719 7 1 2 90183 12718
0 12720 5 1 1 12719
0 12721 7 1 2 65106 79404
0 12722 5 1 1 12721
0 12723 7 1 2 78123 12722
0 12724 5 2 1 12723
0 12725 7 1 2 67406 90402
0 12726 5 1 1 12725
0 12727 7 1 2 2929 12726
0 12728 5 1 1 12727
0 12729 7 3 2 63285 79171
0 12730 7 1 2 12728 90404
0 12731 5 1 1 12730
0 12732 7 1 2 12731 3286
0 12733 5 1 1 12732
0 12734 7 1 2 65957 12733
0 12735 5 1 1 12734
0 12736 7 3 2 69760 81368
0 12737 7 1 2 66671 78103
0 12738 7 1 2 79898 12737
0 12739 7 1 2 90407 12738
0 12740 5 1 1 12739
0 12741 7 1 2 12735 12740
0 12742 5 1 1 12741
0 12743 7 1 2 67648 12742
0 12744 5 1 1 12743
0 12745 7 1 2 79899 81377
0 12746 7 1 2 89439 12745
0 12747 5 1 1 12746
0 12748 7 1 2 12744 12747
0 12749 5 1 1 12748
0 12750 7 1 2 68955 12749
0 12751 5 1 1 12750
0 12752 7 1 2 77028 78673
0 12753 7 2 2 62531 87196
0 12754 7 2 2 63925 82153
0 12755 7 1 2 90410 90412
0 12756 7 1 2 12752 12755
0 12757 5 1 1 12756
0 12758 7 1 2 81552 83209
0 12759 7 1 2 79900 12758
0 12760 7 1 2 71478 12759
0 12761 5 1 1 12760
0 12762 7 1 2 12757 12761
0 12763 5 1 1 12762
0 12764 7 1 2 69530 12763
0 12765 5 1 1 12764
0 12766 7 1 2 12751 12765
0 12767 5 1 1 12766
0 12768 7 1 2 66917 12767
0 12769 5 1 1 12768
0 12770 7 2 2 72122 83583
0 12771 7 1 2 71209 89479
0 12772 7 1 2 90414 12771
0 12773 5 1 1 12772
0 12774 7 1 2 73302 82886
0 12775 7 1 2 89825 12774
0 12776 5 1 1 12775
0 12777 7 1 2 12773 12776
0 12778 5 1 1 12777
0 12779 7 1 2 69761 12778
0 12780 5 1 1 12779
0 12781 7 1 2 81273 75030
0 12782 7 1 2 87104 12781
0 12783 7 3 2 62532 72779
0 12784 5 1 1 90416
0 12785 7 1 2 90417 84916
0 12786 7 1 2 12782 12785
0 12787 5 1 1 12786
0 12788 7 1 2 12780 12787
0 12789 5 1 1 12788
0 12790 7 1 2 66672 12789
0 12791 5 1 1 12790
0 12792 7 1 2 74154 87892
0 12793 7 1 2 82555 12792
0 12794 7 1 2 86404 12793
0 12795 5 1 1 12794
0 12796 7 1 2 12791 12795
0 12797 7 1 2 12769 12796
0 12798 5 1 1 12797
0 12799 7 1 2 84072 12798
0 12800 5 1 1 12799
0 12801 7 1 2 82951 89010
0 12802 5 1 1 12801
0 12803 7 5 2 74070 85496
0 12804 5 1 1 90419
0 12805 7 1 2 79770 90420
0 12806 5 1 1 12805
0 12807 7 1 2 12802 12806
0 12808 5 1 1 12807
0 12809 7 1 2 66918 12808
0 12810 5 1 1 12809
0 12811 7 1 2 76833 73271
0 12812 5 1 1 12811
0 12813 7 1 2 12810 12812
0 12814 5 1 1 12813
0 12815 7 1 2 69762 12814
0 12816 5 1 1 12815
0 12817 7 2 2 62366 85912
0 12818 7 1 2 77408 90424
0 12819 7 1 2 79521 12818
0 12820 5 1 1 12819
0 12821 7 1 2 12816 12820
0 12822 5 1 1 12821
0 12823 7 1 2 81339 88780
0 12824 7 1 2 12822 12823
0 12825 5 1 1 12824
0 12826 7 1 2 12800 12825
0 12827 5 1 1 12826
0 12828 7 1 2 66409 12827
0 12829 5 1 1 12828
0 12830 7 1 2 90403 90405
0 12831 5 1 1 12830
0 12832 7 1 2 79073 85090
0 12833 5 1 1 12832
0 12834 7 1 2 12831 12833
0 12835 5 1 1 12834
0 12836 7 1 2 67407 12835
0 12837 5 1 1 12836
0 12838 7 3 2 78546 80455
0 12839 7 1 2 85059 90426
0 12840 5 1 1 12839
0 12841 7 1 2 12837 12840
0 12842 5 1 1 12841
0 12843 7 1 2 66919 12842
0 12844 5 1 1 12843
0 12845 7 2 2 75477 81617
0 12846 5 1 1 90429
0 12847 7 2 2 79119 80693
0 12848 7 1 2 90430 90431
0 12849 5 1 1 12848
0 12850 7 1 2 12844 12849
0 12851 5 1 1 12850
0 12852 7 1 2 83803 72530
0 12853 7 1 2 12851 12852
0 12854 5 1 1 12853
0 12855 7 1 2 69996 73774
0 12856 7 1 2 75612 12855
0 12857 5 1 1 12856
0 12858 7 1 2 88307 12857
0 12859 5 1 1 12858
0 12860 7 1 2 74464 80085
0 12861 7 1 2 89187 12860
0 12862 7 1 2 12859 12861
0 12863 5 1 1 12862
0 12864 7 1 2 12854 12863
0 12865 5 1 1 12864
0 12866 7 1 2 61501 12865
0 12867 5 1 1 12866
0 12868 7 2 2 72222 79236
0 12869 7 1 2 89193 90433
0 12870 5 1 1 12869
0 12871 7 3 2 71159 83660
0 12872 7 1 2 75853 90435
0 12873 5 1 1 12872
0 12874 7 1 2 12870 12873
0 12875 5 1 1 12874
0 12876 7 1 2 67200 12875
0 12877 5 1 1 12876
0 12878 7 7 2 68956 72695
0 12879 5 2 1 90438
0 12880 7 2 2 85906 90439
0 12881 7 1 2 86602 90447
0 12882 5 1 1 12881
0 12883 7 1 2 12877 12882
0 12884 5 1 1 12883
0 12885 7 1 2 73199 12884
0 12886 5 1 1 12885
0 12887 7 1 2 75763 89411
0 12888 5 1 1 12887
0 12889 7 1 2 83629 78158
0 12890 5 1 1 12889
0 12891 7 1 2 12888 12890
0 12892 5 1 1 12891
0 12893 7 3 2 74071 83210
0 12894 7 1 2 12892 90449
0 12895 5 1 1 12894
0 12896 7 1 2 12886 12895
0 12897 5 1 1 12896
0 12898 7 1 2 66673 12897
0 12899 5 1 1 12898
0 12900 7 1 2 62048 87614
0 12901 5 1 1 12900
0 12902 7 1 2 9418 12901
0 12903 5 4 1 12902
0 12904 7 1 2 68808 79289
0 12905 7 1 2 89441 12904
0 12906 7 1 2 90452 12905
0 12907 5 1 1 12906
0 12908 7 1 2 63286 12907
0 12909 7 1 2 12899 12908
0 12910 5 1 1 12909
0 12911 7 3 2 83530 82272
0 12912 7 1 2 72531 78065
0 12913 7 1 2 90456 12912
0 12914 5 1 1 12913
0 12915 7 2 2 66674 84208
0 12916 7 1 2 79748 86733
0 12917 7 1 2 90459 12916
0 12918 5 1 1 12917
0 12919 7 1 2 12914 12918
0 12920 5 1 1 12919
0 12921 7 1 2 68809 12920
0 12922 5 1 1 12921
0 12923 7 1 2 74019 79727
0 12924 5 1 1 12923
0 12925 7 1 2 12922 12924
0 12926 5 1 1 12925
0 12927 7 1 2 69763 12926
0 12928 5 1 1 12927
0 12929 7 2 2 74072 79771
0 12930 7 1 2 85902 89857
0 12931 7 1 2 90461 12930
0 12932 5 1 1 12931
0 12933 7 1 2 12928 12932
0 12934 5 1 1 12933
0 12935 7 1 2 62049 12934
0 12936 5 1 1 12935
0 12937 7 2 2 75410 76363
0 12938 7 1 2 90463 84351
0 12939 7 1 2 84139 12938
0 12940 5 1 1 12939
0 12941 7 1 2 68124 12940
0 12942 7 1 2 12936 12941
0 12943 5 1 1 12942
0 12944 7 1 2 76131 12943
0 12945 7 1 2 12910 12944
0 12946 5 1 1 12945
0 12947 7 1 2 12867 12946
0 12948 7 1 2 12829 12947
0 12949 5 1 1 12948
0 12950 7 1 2 74540 12949
0 12951 5 1 1 12950
0 12952 7 1 2 83043 77446
0 12953 5 1 1 12952
0 12954 7 1 2 89709 12953
0 12955 5 1 1 12954
0 12956 7 1 2 12955 85866
0 12957 5 1 1 12956
0 12958 7 1 2 82579 71698
0 12959 7 1 2 84677 12958
0 12960 5 1 1 12959
0 12961 7 1 2 12957 12960
0 12962 5 1 1 12961
0 12963 7 1 2 66920 12962
0 12964 5 1 1 12963
0 12965 7 6 2 66675 77145
0 12966 7 2 2 73775 72244
0 12967 5 1 1 90471
0 12968 7 1 2 85010 90472
0 12969 7 1 2 90465 12968
0 12970 5 1 1 12969
0 12971 7 1 2 12964 12970
0 12972 5 1 1 12971
0 12973 7 1 2 84073 12972
0 12974 5 1 1 12973
0 12975 7 9 2 62533 63107
0 12976 7 3 2 62367 90473
0 12977 7 4 2 63287 63926
0 12978 7 1 2 86031 90485
0 12979 7 1 2 90482 12978
0 12980 7 1 2 77509 12979
0 12981 5 1 1 12980
0 12982 7 1 2 12974 12981
0 12983 5 1 1 12982
0 12984 7 1 2 64903 12983
0 12985 5 1 1 12984
0 12986 7 3 2 80028 82734
0 12987 7 1 2 77803 90387
0 12988 7 1 2 90489 12987
0 12989 5 1 1 12988
0 12990 7 2 2 61808 90486
0 12991 7 2 2 67201 80643
0 12992 7 2 2 68957 88731
0 12993 7 1 2 90494 90496
0 12994 7 1 2 90492 12993
0 12995 5 1 1 12994
0 12996 7 1 2 12989 12995
0 12997 5 1 1 12996
0 12998 7 1 2 66921 77681
0 12999 7 1 2 12997 12998
0 13000 5 1 1 12999
0 13001 7 1 2 12985 13000
0 13002 5 1 1 13001
0 13003 7 1 2 61502 13002
0 13004 5 1 1 13003
0 13005 7 1 2 67202 72307
0 13006 5 1 1 13005
0 13007 7 1 2 6014 13006
0 13008 5 1 1 13007
0 13009 7 2 2 88967 76662
0 13010 7 1 2 13008 90498
0 13011 5 1 1 13010
0 13012 7 4 2 63108 81274
0 13013 5 3 1 90500
0 13014 7 2 2 72037 90501
0 13015 5 1 1 90507
0 13016 7 1 2 73824 90508
0 13017 5 1 1 13016
0 13018 7 1 2 67203 87197
0 13019 7 1 2 89667 13018
0 13020 7 1 2 77587 13019
0 13021 5 1 1 13020
0 13022 7 1 2 13017 13021
0 13023 5 1 1 13022
0 13024 7 1 2 61809 13023
0 13025 5 1 1 13024
0 13026 7 1 2 13011 13025
0 13027 5 1 1 13026
0 13028 7 1 2 85725 81664
0 13029 7 1 2 13027 13028
0 13030 5 1 1 13029
0 13031 7 1 2 13004 13030
0 13032 5 1 1 13031
0 13033 7 1 2 64676 13032
0 13034 5 1 1 13033
0 13035 7 1 2 77585 87170
0 13036 5 1 1 13035
0 13037 7 1 2 62368 78024
0 13038 7 1 2 86913 13037
0 13039 5 1 1 13038
0 13040 7 1 2 13036 13039
0 13041 5 1 1 13040
0 13042 7 1 2 82319 13041
0 13043 5 1 1 13042
0 13044 7 2 2 86758 78656
0 13045 7 1 2 83804 83223
0 13046 7 1 2 90509 13045
0 13047 5 1 1 13046
0 13048 7 1 2 13043 13047
0 13049 5 1 1 13048
0 13050 7 1 2 79100 77857
0 13051 7 1 2 13049 13050
0 13052 5 1 1 13051
0 13053 7 1 2 13034 13052
0 13054 5 1 1 13053
0 13055 7 1 2 76973 13054
0 13056 5 1 1 13055
0 13057 7 4 2 71815 78094
0 13058 5 1 1 90511
0 13059 7 5 2 66410 84463
0 13060 7 1 2 78473 88910
0 13061 7 1 2 90515 13060
0 13062 5 2 1 13061
0 13063 7 1 2 86137 83687
0 13064 5 1 1 13063
0 13065 7 1 2 90520 13064
0 13066 5 1 1 13065
0 13067 7 1 2 71160 13066
0 13068 5 1 1 13067
0 13069 7 4 2 67972 68958
0 13070 7 5 2 66411 90522
0 13071 7 2 2 88911 79120
0 13072 7 1 2 70992 90531
0 13073 7 1 2 90526 13072
0 13074 5 1 1 13073
0 13075 7 1 2 13068 13074
0 13076 5 1 1 13075
0 13077 7 1 2 90512 13076
0 13078 5 1 1 13077
0 13079 7 4 2 61503 81651
0 13080 7 1 2 77796 74451
0 13081 7 1 2 80600 13080
0 13082 7 1 2 90533 13081
0 13083 5 1 1 13082
0 13084 7 1 2 71161 71049
0 13085 5 1 1 13084
0 13086 7 1 2 13085 71008
0 13087 5 1 1 13086
0 13088 7 4 2 65107 76132
0 13089 7 1 2 79717 90537
0 13090 7 1 2 13087 13089
0 13091 5 1 1 13090
0 13092 7 1 2 13083 13091
0 13093 5 1 1 13092
0 13094 7 1 2 79429 13093
0 13095 5 1 1 13094
0 13096 7 3 2 63750 77146
0 13097 7 1 2 83861 90541
0 13098 7 1 2 90436 13097
0 13099 5 1 1 13098
0 13100 7 1 2 68125 13099
0 13101 7 1 2 13095 13100
0 13102 5 1 1 13101
0 13103 7 1 2 90157 85935
0 13104 5 2 1 13103
0 13105 7 1 2 76073 90544
0 13106 5 1 1 13105
0 13107 7 1 2 62050 78497
0 13108 7 2 2 88067 13107
0 13109 5 1 1 90546
0 13110 7 1 2 13106 13109
0 13111 5 1 1 13110
0 13112 7 1 2 90437 13111
0 13113 5 1 1 13112
0 13114 7 2 2 68959 78410
0 13115 7 1 2 79430 90548
0 13116 7 2 2 80803 87478
0 13117 7 1 2 90550 81234
0 13118 7 1 2 13115 13117
0 13119 5 1 1 13118
0 13120 7 1 2 63288 13119
0 13121 7 1 2 13113 13120
0 13122 5 1 1 13121
0 13123 7 1 2 68359 13122
0 13124 7 1 2 13102 13123
0 13125 5 1 1 13124
0 13126 7 1 2 13078 13125
0 13127 5 1 1 13126
0 13128 7 1 2 71570 13127
0 13129 5 1 1 13128
0 13130 7 1 2 81618 76554
0 13131 7 1 2 78749 79431
0 13132 7 1 2 83211 13131
0 13133 7 1 2 13130 13132
0 13134 5 1 1 13133
0 13135 7 4 2 69332 88241
0 13136 7 2 2 68126 70993
0 13137 7 1 2 90552 90556
0 13138 5 1 1 13137
0 13139 7 1 2 86876 87089
0 13140 5 1 1 13139
0 13141 7 1 2 13138 13140
0 13142 5 1 1 13141
0 13143 7 1 2 68360 90538
0 13144 7 1 2 13142 13143
0 13145 5 1 1 13144
0 13146 7 1 2 13134 13145
0 13147 5 1 1 13146
0 13148 7 1 2 89637 13147
0 13149 5 1 1 13148
0 13150 7 4 2 66412 81241
0 13151 5 3 1 90558
0 13152 7 7 2 70884 86942
0 13153 5 1 1 90565
0 13154 7 1 2 90562 13153
0 13155 5 3 1 13154
0 13156 7 1 2 83805 74247
0 13157 7 1 2 89175 13156
0 13158 7 1 2 90572 13157
0 13159 5 1 1 13158
0 13160 7 1 2 13149 13159
0 13161 5 1 1 13160
0 13162 7 1 2 79718 13161
0 13163 5 1 1 13162
0 13164 7 1 2 13129 13163
0 13165 7 1 2 13056 13164
0 13166 7 1 2 12951 13165
0 13167 7 1 2 12720 13166
0 13168 7 1 2 12360 13167
0 13169 7 1 2 11635 13168
0 13170 7 1 2 10798 13169
0 13171 5 1 1 13170
0 13172 7 1 2 69165 13171
0 13173 5 1 1 13172
0 13174 7 1 2 8804 13173
0 13175 5 1 1 13174
0 13176 7 1 2 61259 13175
0 13177 5 1 1 13176
0 13178 7 2 2 61810 73303
0 13179 7 5 2 69166 82803
0 13180 7 11 2 63751 81619
0 13181 7 1 2 90577 90582
0 13182 7 1 2 90575 13181
0 13183 7 1 2 75304 90023
0 13184 7 1 2 87678 13183
0 13185 7 1 2 87669 13184
0 13186 7 1 2 13182 13185
0 13187 5 1 1 13186
0 13188 7 1 2 13177 13187
0 13189 5 1 1 13188
0 13190 7 40 2 61343 62995
0 13191 5 5 1 90593
0 13192 7 9 2 67760 90594
0 13193 5 1 1 90638
0 13194 7 45 2 66205 67837
0 13195 5 3 1 90647
0 13196 7 2 2 62940 90648
0 13197 5 1 1 90695
0 13198 7 1 2 13193 13197
0 13199 5 42 1 13198
0 13200 7 1 2 13189 90697
0 13201 5 1 1 13200
0 13202 7 1 2 88432 81230
0 13203 5 4 1 13202
0 13204 7 1 2 81369 90739
0 13205 5 1 1 13204
0 13206 7 4 2 62369 81620
0 13207 7 1 2 78148 88092
0 13208 7 1 2 90743 13207
0 13209 5 1 1 13208
0 13210 7 1 2 13205 13209
0 13211 5 1 1 13210
0 13212 7 1 2 63109 13211
0 13213 5 1 1 13212
0 13214 7 1 2 88294 80439
0 13215 7 1 2 88444 13214
0 13216 5 1 1 13215
0 13217 7 1 2 13213 13216
0 13218 5 1 1 13217
0 13219 7 1 2 82234 13218
0 13220 5 1 1 13219
0 13221 7 1 2 81728 90397
0 13222 5 1 1 13221
0 13223 7 1 2 13220 13222
0 13224 5 1 1 13223
0 13225 7 1 2 62051 13224
0 13226 5 1 1 13225
0 13227 7 1 2 68127 76799
0 13228 7 1 2 83656 13227
0 13229 5 1 1 13228
0 13230 7 3 2 68361 79603
0 13231 5 2 1 90747
0 13232 7 5 2 64904 79347
0 13233 7 1 2 90752 85133
0 13234 7 1 2 90748 13233
0 13235 5 1 1 13234
0 13236 7 1 2 13229 13235
0 13237 5 1 1 13236
0 13238 7 1 2 63110 13237
0 13239 5 1 1 13238
0 13240 7 1 2 13226 13239
0 13241 5 1 1 13240
0 13242 7 1 2 66413 13241
0 13243 5 1 1 13242
0 13244 7 1 2 78914 90740
0 13245 5 1 1 13244
0 13246 7 1 2 78865 87445
0 13247 5 1 1 13246
0 13248 7 1 2 13245 13247
0 13249 5 1 1 13248
0 13250 7 1 2 62052 13249
0 13251 5 1 1 13250
0 13252 7 4 2 67973 69997
0 13253 7 22 2 69531 65369
0 13254 7 2 2 75379 90761
0 13255 7 1 2 90757 90783
0 13256 5 1 1 13255
0 13257 7 1 2 13251 13256
0 13258 5 1 1 13257
0 13259 7 1 2 68128 13258
0 13260 5 1 1 13259
0 13261 7 4 2 80440 90583
0 13262 5 3 1 90785
0 13263 7 1 2 88093 77374
0 13264 7 1 2 90786 13263
0 13265 5 1 1 13264
0 13266 7 1 2 13260 13265
0 13267 5 1 1 13266
0 13268 7 1 2 69764 82842
0 13269 7 1 2 13267 13268
0 13270 5 1 1 13269
0 13271 7 1 2 13243 13270
0 13272 5 1 1 13271
0 13273 7 1 2 76271 13272
0 13274 5 1 1 13273
0 13275 7 6 2 68129 63927
0 13276 7 3 2 62053 90792
0 13277 7 1 2 80667 84182
0 13278 7 1 2 90798 13277
0 13279 7 1 2 90741 13278
0 13280 5 1 1 13279
0 13281 7 1 2 61811 13280
0 13282 7 1 2 13274 13281
0 13283 5 1 1 13282
0 13284 7 3 2 70283 79250
0 13285 7 1 2 85214 79575
0 13286 5 1 1 13285
0 13287 7 1 2 86814 76272
0 13288 5 1 1 13287
0 13289 7 1 2 13286 13288
0 13290 5 1 1 13289
0 13291 7 1 2 78866 13290
0 13292 5 1 1 13291
0 13293 7 2 2 67204 78750
0 13294 7 1 2 78235 87105
0 13295 7 1 2 90804 13294
0 13296 5 1 1 13295
0 13297 7 1 2 13292 13296
0 13298 5 1 1 13297
0 13299 7 1 2 68130 13298
0 13300 5 1 1 13299
0 13301 7 5 2 77297 77449
0 13302 7 2 2 81729 83584
0 13303 7 1 2 90806 90811
0 13304 5 1 1 13303
0 13305 7 1 2 13300 13304
0 13306 5 1 1 13305
0 13307 7 1 2 69333 13306
0 13308 5 1 1 13307
0 13309 7 2 2 88295 83645
0 13310 7 4 2 69998 71298
0 13311 7 1 2 87559 90024
0 13312 7 1 2 90815 13311
0 13313 7 1 2 90813 13312
0 13314 5 1 1 13313
0 13315 7 1 2 13308 13314
0 13316 5 1 1 13315
0 13317 7 1 2 64905 13316
0 13318 5 1 1 13317
0 13319 7 3 2 79348 83474
0 13320 7 1 2 82657 79221
0 13321 7 1 2 90816 13320
0 13322 7 1 2 90819 13321
0 13323 5 1 1 13322
0 13324 7 1 2 13318 13323
0 13325 5 1 1 13324
0 13326 7 1 2 90801 13325
0 13327 5 1 1 13326
0 13328 7 1 2 80813 87631
0 13329 5 1 1 13328
0 13330 7 1 2 87608 78743
0 13331 5 5 1 13330
0 13332 7 1 2 63928 88813
0 13333 7 1 2 90822 13332
0 13334 5 1 1 13333
0 13335 7 1 2 13329 13334
0 13336 5 1 1 13335
0 13337 7 1 2 62534 13336
0 13338 5 1 1 13337
0 13339 7 2 2 82658 87400
0 13340 7 1 2 78674 76208
0 13341 7 1 2 90827 13340
0 13342 5 1 1 13341
0 13343 7 1 2 13338 13342
0 13344 5 1 1 13343
0 13345 7 1 2 72986 13344
0 13346 5 1 1 13345
0 13347 7 1 2 68131 90453
0 13348 5 1 1 13347
0 13349 7 1 2 84783 86538
0 13350 5 1 1 13349
0 13351 7 1 2 13348 13350
0 13352 5 1 1 13351
0 13353 7 1 2 89180 13352
0 13354 5 1 1 13353
0 13355 7 1 2 13346 13354
0 13356 5 1 1 13355
0 13357 7 1 2 79432 13356
0 13358 5 1 1 13357
0 13359 7 2 2 81695 86091
0 13360 7 2 2 76133 74356
0 13361 7 1 2 72987 76273
0 13362 7 1 2 90831 13361
0 13363 7 1 2 90829 13362
0 13364 5 1 1 13363
0 13365 7 1 2 13358 13364
0 13366 5 1 1 13365
0 13367 7 1 2 65370 13366
0 13368 5 1 1 13367
0 13369 7 2 2 69334 73304
0 13370 7 1 2 81275 89372
0 13371 7 1 2 90833 13370
0 13372 5 1 1 13371
0 13373 7 1 2 76818 71704
0 13374 5 2 1 13373
0 13375 7 1 2 83478 90835
0 13376 5 1 1 13375
0 13377 7 1 2 71299 88905
0 13378 7 1 2 13376 13377
0 13379 5 1 1 13378
0 13380 7 1 2 13372 13379
0 13381 5 1 1 13380
0 13382 7 1 2 79604 13381
0 13383 5 1 1 13382
0 13384 7 1 2 88604 81857
0 13385 5 1 1 13384
0 13386 7 1 2 13383 13385
0 13387 5 1 1 13386
0 13388 7 1 2 62054 13387
0 13389 5 1 1 13388
0 13390 7 1 2 74008 82714
0 13391 7 3 2 63929 79433
0 13392 7 1 2 86332 90837
0 13393 7 1 2 13390 13392
0 13394 5 1 1 13393
0 13395 7 1 2 13389 13394
0 13396 5 1 1 13395
0 13397 7 1 2 67974 13396
0 13398 5 1 1 13397
0 13399 7 4 2 69999 82539
0 13400 7 1 2 87434 90840
0 13401 5 1 1 13400
0 13402 7 1 2 76462 88272
0 13403 5 1 1 13402
0 13404 7 1 2 13401 13403
0 13405 5 1 1 13404
0 13406 7 6 2 62055 71300
0 13407 5 1 1 90844
0 13408 7 2 2 86434 82074
0 13409 7 1 2 63111 90850
0 13410 7 1 2 90845 13409
0 13411 7 1 2 13405 13410
0 13412 5 1 1 13411
0 13413 7 1 2 13398 13412
0 13414 5 1 1 13413
0 13415 7 1 2 61504 13414
0 13416 5 1 1 13415
0 13417 7 1 2 66676 13416
0 13418 7 1 2 13368 13417
0 13419 7 1 2 13327 13418
0 13420 5 1 1 13419
0 13421 7 1 2 62941 13420
0 13422 7 1 2 13283 13421
0 13423 5 1 1 13422
0 13424 7 2 2 88456 86092
0 13425 7 2 2 70284 90852
0 13426 7 16 2 63930 69335
0 13427 7 13 2 62535 67761
0 13428 7 1 2 90856 90872
0 13429 7 1 2 87655 13428
0 13430 7 1 2 90854 13429
0 13431 5 1 1 13430
0 13432 7 1 2 13423 13431
0 13433 5 1 1 13432
0 13434 7 1 2 64319 13433
0 13435 5 1 1 13434
0 13436 7 5 2 72988 73305
0 13437 5 1 1 90885
0 13438 7 1 2 74896 13437
0 13439 5 1 1 13438
0 13440 7 1 2 76882 13439
0 13441 5 1 1 13440
0 13442 7 4 2 76463 77637
0 13443 7 3 2 65108 90890
0 13444 5 1 1 90894
0 13445 7 1 2 13441 13444
0 13446 5 1 1 13445
0 13447 7 1 2 80506 82843
0 13448 7 1 2 13446 13447
0 13449 5 1 1 13448
0 13450 7 3 2 78149 80293
0 13451 5 1 1 90897
0 13452 7 9 2 62536 69336
0 13453 7 1 2 77298 90900
0 13454 7 1 2 87275 13453
0 13455 7 1 2 90898 13454
0 13456 5 1 1 13455
0 13457 7 1 2 13449 13456
0 13458 5 1 1 13457
0 13459 7 1 2 83101 13458
0 13460 5 1 1 13459
0 13461 7 1 2 63112 88212
0 13462 5 1 1 13461
0 13463 7 1 2 90789 13462
0 13464 5 2 1 13463
0 13465 7 1 2 81983 90909
0 13466 5 1 1 13465
0 13467 7 1 2 88220 76015
0 13468 5 1 1 13467
0 13469 7 1 2 13466 13468
0 13470 5 1 1 13469
0 13471 7 1 2 61505 13470
0 13472 5 1 1 13471
0 13473 7 5 2 81621 77193
0 13474 7 1 2 79855 90025
0 13475 7 1 2 90911 13474
0 13476 5 1 1 13475
0 13477 7 1 2 13472 13476
0 13478 5 1 1 13477
0 13479 7 3 2 62537 79532
0 13480 7 1 2 73604 90916
0 13481 7 1 2 13478 13480
0 13482 5 1 1 13481
0 13483 7 1 2 13460 13482
0 13484 5 1 1 13483
0 13485 7 1 2 64677 13484
0 13486 5 1 1 13485
0 13487 7 1 2 73306 90742
0 13488 5 1 1 13487
0 13489 7 1 2 8739 13488
0 13490 5 1 1 13489
0 13491 7 1 2 76016 13490
0 13492 5 1 1 13491
0 13493 7 1 2 90895 87240
0 13494 5 1 1 13493
0 13495 7 1 2 13492 13494
0 13496 5 1 1 13495
0 13497 7 1 2 68132 13496
0 13498 5 1 1 13497
0 13499 7 4 2 61812 75945
0 13500 5 1 1 90919
0 13501 7 3 2 63516 74567
0 13502 7 1 2 66677 90923
0 13503 5 1 1 13502
0 13504 7 1 2 13500 13503
0 13505 5 1 1 13504
0 13506 7 1 2 62370 13505
0 13507 5 1 1 13506
0 13508 7 1 2 61813 75928
0 13509 5 1 1 13508
0 13510 7 1 2 13507 13509
0 13511 5 1 1 13510
0 13512 7 1 2 73307 13511
0 13513 5 1 1 13512
0 13514 7 1 2 63517 90920
0 13515 5 1 1 13514
0 13516 7 1 2 13513 13515
0 13517 5 1 1 13516
0 13518 7 1 2 13517 83684
0 13519 5 1 1 13518
0 13520 7 1 2 61506 13519
0 13521 7 1 2 13498 13520
0 13522 5 1 1 13521
0 13523 7 3 2 63113 89106
0 13524 5 1 1 90926
0 13525 7 1 2 81747 13524
0 13526 5 1 1 13525
0 13527 7 1 2 71816 13526
0 13528 5 1 1 13527
0 13529 7 1 2 80704 81753
0 13530 5 1 1 13529
0 13531 7 1 2 13528 13530
0 13532 5 1 1 13531
0 13533 7 1 2 69765 13532
0 13534 5 1 1 13533
0 13535 7 1 2 89865 89757
0 13536 5 1 1 13535
0 13537 7 1 2 13534 13536
0 13538 5 1 1 13537
0 13539 7 1 2 61814 13538
0 13540 5 1 1 13539
0 13541 7 1 2 78066 75997
0 13542 7 1 2 89737 13541
0 13543 5 1 1 13542
0 13544 7 1 2 13540 13543
0 13545 5 1 1 13544
0 13546 7 1 2 86548 13545
0 13547 5 1 1 13546
0 13548 7 10 2 63752 89718
0 13549 7 1 2 65109 81679
0 13550 7 1 2 80507 13549
0 13551 7 1 2 90929 13550
0 13552 5 1 1 13551
0 13553 7 1 2 66414 13552
0 13554 7 1 2 13547 13553
0 13555 5 1 1 13554
0 13556 7 1 2 79349 13555
0 13557 7 1 2 13522 13556
0 13558 5 1 1 13557
0 13559 7 1 2 13486 13558
0 13560 5 1 1 13559
0 13561 7 1 2 62056 13560
0 13562 5 1 1 13561
0 13563 7 1 2 69766 88312
0 13564 5 1 1 13563
0 13565 7 2 2 78547 80483
0 13566 7 1 2 84472 90939
0 13567 5 1 1 13566
0 13568 7 1 2 13564 13567
0 13569 5 1 1 13568
0 13570 7 1 2 76800 13569
0 13571 5 1 1 13570
0 13572 7 1 2 87553 83502
0 13573 5 1 1 13572
0 13574 7 1 2 13571 13573
0 13575 5 1 1 13574
0 13576 7 1 2 81696 73308
0 13577 7 1 2 13575 13576
0 13578 5 1 1 13577
0 13579 7 1 2 13562 13578
0 13580 5 1 1 13579
0 13581 7 1 2 62801 13580
0 13582 5 1 1 13581
0 13583 7 1 2 89866 86081
0 13584 7 3 2 63518 82982
0 13585 7 1 2 82910 90941
0 13586 7 1 2 13583 13585
0 13587 5 1 1 13586
0 13588 7 1 2 13582 13587
0 13589 5 1 1 13588
0 13590 7 2 2 69167 13589
0 13591 5 1 1 90944
0 13592 7 1 2 67762 90945
0 13593 5 1 1 13592
0 13594 7 1 2 13435 13593
0 13595 5 1 1 13594
0 13596 7 1 2 90595 13595
0 13597 5 1 1 13596
0 13598 7 6 2 66206 62942
0 13599 7 3 2 67838 90946
0 13600 7 9 2 63114 64320
0 13601 7 4 2 88912 90955
0 13602 7 3 2 63519 90964
0 13603 7 1 2 77716 90968
0 13604 7 1 2 90855 13603
0 13605 5 1 1 13604
0 13606 7 1 2 13591 13605
0 13607 5 2 1 13606
0 13608 7 1 2 90952 90971
0 13609 5 1 1 13608
0 13610 7 1 2 13597 13609
0 13611 5 1 1 13610
0 13612 7 1 2 61260 13611
0 13613 5 1 1 13612
0 13614 7 11 2 62943 62996
0 13615 7 20 2 66089 61344
0 13616 7 8 2 90973 90984
0 13617 5 1 1 91004
0 13618 7 1 2 91005 90972
0 13619 5 1 1 13618
0 13620 7 1 2 13613 13619
0 13621 5 1 1 13620
0 13622 7 1 2 78322 13621
0 13623 5 1 1 13622
0 13624 7 3 2 61261 90698
0 13625 5 1 1 91012
0 13626 7 1 2 13625 13617
0 13627 5 25 1 13626
0 13628 7 3 2 72989 76134
0 13629 7 5 2 70285 72268
0 13630 7 2 2 85913 91043
0 13631 7 1 2 84134 75287
0 13632 7 1 2 91048 13631
0 13633 5 1 1 13632
0 13634 7 1 2 67408 75631
0 13635 5 1 1 13634
0 13636 7 1 2 78639 13635
0 13637 5 2 1 13636
0 13638 7 3 2 70885 79434
0 13639 7 1 2 84713 91052
0 13640 7 1 2 73117 13639
0 13641 7 1 2 91050 13640
0 13642 5 1 1 13641
0 13643 7 1 2 13633 13642
0 13644 5 1 1 13643
0 13645 7 1 2 65110 13644
0 13646 5 1 1 13645
0 13647 7 2 2 81409 90457
0 13648 7 4 2 70000 71210
0 13649 7 3 2 76316 76246
0 13650 7 1 2 91057 91061
0 13651 7 1 2 91055 13650
0 13652 5 1 1 13651
0 13653 7 1 2 13646 13652
0 13654 5 1 1 13653
0 13655 7 1 2 91040 13654
0 13656 5 1 1 13655
0 13657 7 4 2 72038 77354
0 13658 5 1 1 91064
0 13659 7 1 2 76791 91065
0 13660 5 1 1 13659
0 13661 7 1 2 84105 73118
0 13662 5 1 1 13661
0 13663 7 1 2 13660 13662
0 13664 5 1 1 13663
0 13665 7 1 2 67409 13664
0 13666 5 1 1 13665
0 13667 7 1 2 62538 76792
0 13668 7 1 2 81155 13667
0 13669 5 1 1 13668
0 13670 7 1 2 13666 13669
0 13671 5 1 1 13670
0 13672 7 1 2 79967 82936
0 13673 7 1 2 82945 13672
0 13674 7 1 2 13671 13673
0 13675 5 1 1 13674
0 13676 7 1 2 61507 72039
0 13677 7 1 2 74791 13676
0 13678 7 1 2 83995 13677
0 13679 7 1 2 79050 13678
0 13680 7 1 2 91051 13679
0 13681 5 1 1 13680
0 13682 7 1 2 13675 13681
0 13683 5 1 1 13682
0 13684 7 1 2 68133 13683
0 13685 5 1 1 13684
0 13686 7 1 2 13656 13685
0 13687 5 1 1 13686
0 13688 7 1 2 91015 13687
0 13689 5 1 1 13688
0 13690 7 2 2 91016 76693
0 13691 7 2 2 64906 89808
0 13692 7 1 2 84373 91070
0 13693 5 2 1 13692
0 13694 7 1 2 71428 85839
0 13695 5 1 1 13694
0 13696 7 1 2 91072 13695
0 13697 5 1 1 13696
0 13698 7 2 2 61508 72990
0 13699 7 1 2 68134 80644
0 13700 7 1 2 81574 13699
0 13701 7 1 2 91074 13700
0 13702 7 1 2 13697 13701
0 13703 7 1 2 91068 13702
0 13704 5 1 1 13703
0 13705 7 1 2 13689 13704
0 13706 5 1 1 13705
0 13707 7 1 2 69168 13706
0 13708 5 1 1 13707
0 13709 7 2 2 84007 73934
0 13710 5 3 1 91076
0 13711 7 1 2 83190 91078
0 13712 5 2 1 13711
0 13713 7 1 2 63753 91081
0 13714 5 1 1 13713
0 13715 7 15 2 70286 71921
0 13716 5 2 1 91083
0 13717 7 1 2 86196 91084
0 13718 5 1 1 13717
0 13719 7 1 2 13714 13718
0 13720 5 1 1 13719
0 13721 7 1 2 65111 13720
0 13722 5 1 1 13721
0 13723 7 11 2 67649 70886
0 13724 5 3 1 91100
0 13725 7 1 2 78187 91101
0 13726 7 2 2 86347 13725
0 13727 5 1 1 91114
0 13728 7 1 2 13722 13727
0 13729 5 1 1 13728
0 13730 7 1 2 64094 13729
0 13731 5 1 1 13730
0 13732 7 1 2 63754 71124
0 13733 7 1 2 84849 13732
0 13734 5 1 1 13733
0 13735 7 1 2 13731 13734
0 13736 5 1 1 13735
0 13737 7 1 2 78867 13736
0 13738 5 1 1 13737
0 13739 7 2 2 71922 72820
0 13740 7 1 2 65371 91116
0 13741 5 1 1 13740
0 13742 7 1 2 86120 13741
0 13743 5 1 1 13742
0 13744 7 2 2 70001 78915
0 13745 7 1 2 77809 91118
0 13746 7 1 2 13743 13745
0 13747 5 1 1 13746
0 13748 7 1 2 13738 13747
0 13749 5 1 1 13748
0 13750 7 1 2 81441 13749
0 13751 5 1 1 13750
0 13752 7 7 2 70887 71923
0 13753 7 1 2 84920 91120
0 13754 5 1 1 13753
0 13755 7 1 2 63755 80078
0 13756 5 1 1 13755
0 13757 7 1 2 13754 13756
0 13758 5 1 1 13757
0 13759 7 1 2 78868 13758
0 13760 5 1 1 13759
0 13761 7 3 2 72269 80096
0 13762 7 2 2 67975 91127
0 13763 7 1 2 75219 91130
0 13764 5 1 1 13763
0 13765 7 1 2 13760 13764
0 13766 5 1 1 13765
0 13767 7 1 2 70287 13766
0 13768 5 1 1 13767
0 13769 7 2 2 80321 84008
0 13770 7 1 2 63115 89336
0 13771 7 1 2 91132 13770
0 13772 5 1 1 13771
0 13773 7 1 2 13768 13772
0 13774 5 1 1 13773
0 13775 7 1 2 65112 13774
0 13776 5 1 1 13775
0 13777 7 1 2 70888 71652
0 13778 5 1 1 13777
0 13779 7 1 2 84873 13778
0 13780 5 1 1 13779
0 13781 7 1 2 71924 13780
0 13782 5 1 1 13781
0 13783 7 1 2 76335 74836
0 13784 5 1 1 13783
0 13785 7 1 2 72955 78168
0 13786 5 1 1 13785
0 13787 7 1 2 13784 13786
0 13788 5 1 1 13787
0 13789 7 1 2 13782 13788
0 13790 5 1 1 13789
0 13791 7 1 2 65372 13790
0 13792 5 1 1 13791
0 13793 7 1 2 74633 75000
0 13794 7 1 2 79985 13793
0 13795 5 1 1 13794
0 13796 7 1 2 13792 13795
0 13797 5 1 1 13796
0 13798 7 1 2 91119 13797
0 13799 5 1 1 13798
0 13800 7 1 2 13776 13799
0 13801 5 1 1 13800
0 13802 7 1 2 83044 13801
0 13803 5 1 1 13802
0 13804 7 1 2 13751 13803
0 13805 5 1 1 13804
0 13806 7 1 2 66415 13805
0 13807 5 1 1 13806
0 13808 7 3 2 84839 80548
0 13809 7 1 2 63756 91134
0 13810 5 1 1 13809
0 13811 7 2 2 64095 91121
0 13812 7 1 2 71724 91137
0 13813 5 1 1 13812
0 13814 7 1 2 13810 13813
0 13815 5 1 1 13814
0 13816 7 1 2 13815 87028
0 13817 5 1 1 13816
0 13818 7 1 2 64096 81442
0 13819 7 1 2 91115 13818
0 13820 5 1 1 13819
0 13821 7 1 2 13817 13820
0 13822 5 1 1 13821
0 13823 7 1 2 89078 13822
0 13824 5 1 1 13823
0 13825 7 1 2 13807 13824
0 13826 5 1 1 13825
0 13827 7 1 2 68810 13826
0 13828 5 1 1 13827
0 13829 7 3 2 76935 81242
0 13830 7 1 2 61815 81809
0 13831 7 1 2 91139 13830
0 13832 5 1 1 13831
0 13833 7 1 2 76663 76694
0 13834 7 1 2 88600 13833
0 13835 5 1 1 13834
0 13836 7 1 2 13832 13835
0 13837 5 1 1 13836
0 13838 7 1 2 66416 13837
0 13839 5 1 1 13838
0 13840 7 3 2 63289 76040
0 13841 7 9 2 65699 76883
0 13842 5 1 1 91145
0 13843 7 1 2 66678 83888
0 13844 7 1 2 91146 13843
0 13845 7 1 2 91142 13844
0 13846 5 1 1 13845
0 13847 7 1 2 13839 13846
0 13848 5 1 1 13847
0 13849 7 1 2 88060 13848
0 13850 5 1 1 13849
0 13851 7 1 2 89329 76429
0 13852 7 1 2 88331 13851
0 13853 7 1 2 86518 13852
0 13854 5 1 1 13853
0 13855 7 1 2 13850 13854
0 13856 7 1 2 13828 13855
0 13857 5 1 1 13856
0 13858 7 1 2 67410 13857
0 13859 5 1 1 13858
0 13860 7 4 2 65373 78236
0 13861 7 8 2 70889 78916
0 13862 5 1 1 91158
0 13863 7 1 2 91154 91159
0 13864 5 2 1 13863
0 13865 7 3 2 64678 76936
0 13866 7 1 2 63116 80471
0 13867 7 1 2 91168 13866
0 13868 5 1 1 13867
0 13869 7 1 2 91166 13868
0 13870 5 1 1 13869
0 13871 7 1 2 67650 13870
0 13872 5 1 1 13871
0 13873 7 1 2 91169 80829
0 13874 5 1 1 13873
0 13875 7 1 2 91167 13874
0 13876 5 1 1 13875
0 13877 7 1 2 68960 13876
0 13878 5 1 1 13877
0 13879 7 1 2 13872 13878
0 13880 5 1 1 13879
0 13881 7 1 2 83102 13880
0 13882 5 1 1 13881
0 13883 7 2 2 66679 87198
0 13884 7 2 2 72040 78869
0 13885 5 2 1 91173
0 13886 7 1 2 91155 91174
0 13887 7 1 2 91171 13886
0 13888 5 1 1 13887
0 13889 7 1 2 13882 13888
0 13890 5 1 1 13889
0 13891 7 1 2 65700 13890
0 13892 5 1 1 13891
0 13893 7 1 2 76974 81498
0 13894 7 1 2 91131 13893
0 13895 5 1 1 13894
0 13896 7 1 2 13892 13895
0 13897 5 1 1 13896
0 13898 7 1 2 67205 13897
0 13899 5 1 1 13898
0 13900 7 1 2 88332 80873
0 13901 7 1 2 76607 77772
0 13902 7 1 2 13900 13901
0 13903 5 1 1 13902
0 13904 7 1 2 13899 13903
0 13905 5 1 1 13904
0 13906 7 1 2 66417 13905
0 13907 5 1 1 13906
0 13908 7 1 2 76915 88476
0 13909 7 2 2 78805 79679
0 13910 7 1 2 83446 91177
0 13911 7 1 2 13908 13910
0 13912 5 1 1 13911
0 13913 7 1 2 13907 13912
0 13914 7 1 2 13859 13913
0 13915 5 1 1 13914
0 13916 7 1 2 64907 13915
0 13917 5 1 1 13916
0 13918 7 3 2 66680 88942
0 13919 7 15 2 69532 65701
0 13920 7 4 2 82522 91182
0 13921 7 2 2 70002 91197
0 13922 7 1 2 82946 91201
0 13923 5 1 1 13922
0 13924 7 1 2 65113 80322
0 13925 7 1 2 91041 13924
0 13926 5 1 1 13925
0 13927 7 1 2 13923 13926
0 13928 5 1 1 13927
0 13929 7 1 2 72123 13928
0 13930 5 1 1 13929
0 13931 7 2 2 65702 82756
0 13932 7 1 2 88296 91203
0 13933 5 1 1 13932
0 13934 7 1 2 74837 84958
0 13935 7 1 2 81255 13934
0 13936 5 1 1 13935
0 13937 7 1 2 13933 13936
0 13938 5 1 1 13937
0 13939 7 1 2 78136 13938
0 13940 5 1 1 13939
0 13941 7 5 2 66418 80086
0 13942 7 6 2 70003 76317
0 13943 7 2 2 68599 80097
0 13944 7 1 2 91210 91216
0 13945 7 1 2 91205 13944
0 13946 5 1 1 13945
0 13947 7 1 2 13940 13946
0 13948 5 1 1 13947
0 13949 7 1 2 68811 13948
0 13950 5 1 1 13949
0 13951 7 1 2 13930 13950
0 13952 5 1 1 13951
0 13953 7 1 2 67411 13952
0 13954 5 1 1 13953
0 13955 7 4 2 80184 77810
0 13956 7 2 2 89159 79281
0 13957 7 1 2 91218 91222
0 13958 5 1 1 13957
0 13959 7 2 2 71489 77831
0 13960 5 1 1 91224
0 13961 7 1 2 72941 86694
0 13962 5 1 1 13961
0 13963 7 1 2 13960 13962
0 13964 5 1 1 13963
0 13965 7 1 2 81256 13964
0 13966 5 1 1 13965
0 13967 7 1 2 13958 13966
0 13968 5 1 1 13967
0 13969 7 1 2 84343 13968
0 13970 5 1 1 13969
0 13971 7 1 2 13954 13970
0 13972 5 1 1 13971
0 13973 7 1 2 70288 13972
0 13974 5 1 1 13973
0 13975 7 6 2 69533 81665
0 13976 7 1 2 74792 72334
0 13977 5 1 1 13976
0 13978 7 3 2 67206 77867
0 13979 5 2 1 91232
0 13980 7 1 2 71925 91235
0 13981 7 1 2 89506 13980
0 13982 7 1 2 87889 13981
0 13983 5 1 1 13982
0 13984 7 1 2 13977 13983
0 13985 5 1 1 13984
0 13986 7 1 2 91226 13985
0 13987 5 1 1 13986
0 13988 7 2 2 72270 80162
0 13989 7 1 2 87281 91237
0 13990 5 1 1 13989
0 13991 7 1 2 13987 13990
0 13992 5 1 1 13991
0 13993 7 1 2 65374 90758
0 13994 7 1 2 13992 13993
0 13995 5 1 1 13994
0 13996 7 1 2 13974 13995
0 13997 5 1 1 13996
0 13998 7 1 2 91179 13997
0 13999 5 1 1 13998
0 14000 7 1 2 13917 13999
0 14001 5 1 1 14000
0 14002 7 1 2 69337 14001
0 14003 5 1 1 14002
0 14004 7 1 2 85338 84480
0 14005 5 1 1 14004
0 14006 7 1 2 84937 87530
0 14007 5 2 1 14006
0 14008 7 1 2 14005 91239
0 14009 5 1 1 14008
0 14010 7 1 2 78870 14009
0 14011 5 1 1 14010
0 14012 7 3 2 70653 84379
0 14013 5 5 1 91241
0 14014 7 1 2 77839 91244
0 14015 5 4 1 14014
0 14016 7 9 2 67976 82735
0 14017 7 1 2 82776 91253
0 14018 7 1 2 91249 14017
0 14019 5 1 1 14018
0 14020 7 1 2 14011 14019
0 14021 5 1 1 14020
0 14022 7 1 2 66419 14021
0 14023 5 1 1 14022
0 14024 7 1 2 71125 84481
0 14025 5 1 1 14024
0 14026 7 1 2 91240 14025
0 14027 5 1 1 14026
0 14028 7 1 2 89079 14027
0 14029 5 1 1 14028
0 14030 7 1 2 14023 14029
0 14031 5 1 1 14030
0 14032 7 1 2 69338 14031
0 14033 5 1 1 14032
0 14034 7 4 2 81754 78498
0 14035 7 1 2 86138 91262
0 14036 7 1 2 85339 14035
0 14037 5 1 1 14036
0 14038 7 1 2 14033 14037
0 14039 5 1 1 14038
0 14040 7 1 2 76937 14039
0 14041 5 1 1 14040
0 14042 7 1 2 67651 81425
0 14043 5 1 1 14042
0 14044 7 1 2 90504 14043
0 14045 5 1 1 14044
0 14046 7 1 2 61509 14045
0 14047 5 1 1 14046
0 14048 7 1 2 81410 83509
0 14049 5 1 1 14048
0 14050 7 1 2 14047 14049
0 14051 5 1 1 14050
0 14052 7 1 2 64480 14051
0 14053 5 1 1 14052
0 14054 7 1 2 82601 81333
0 14055 5 1 1 14054
0 14056 7 1 2 14053 14055
0 14057 5 1 1 14056
0 14058 7 1 2 61816 14057
0 14059 5 1 1 14058
0 14060 7 6 2 61510 81755
0 14061 7 1 2 75683 82235
0 14062 7 1 2 91266 14061
0 14063 5 1 1 14062
0 14064 7 1 2 14059 14063
0 14065 5 1 1 14064
0 14066 7 1 2 91147 80056
0 14067 7 1 2 14065 14066
0 14068 5 1 1 14067
0 14069 7 1 2 14041 14068
0 14070 5 1 1 14069
0 14071 7 1 2 72991 14070
0 14072 5 1 1 14071
0 14073 7 4 2 68961 70890
0 14074 5 1 1 91272
0 14075 7 1 2 90502 91273
0 14076 5 1 1 14075
0 14077 7 1 2 81426 84763
0 14078 5 1 1 14077
0 14079 7 1 2 14076 14078
0 14080 5 1 1 14079
0 14081 7 1 2 61511 14080
0 14082 5 1 1 14081
0 14083 7 1 2 76074 71691
0 14084 7 1 2 84455 14083
0 14085 5 1 1 14084
0 14086 7 1 2 14082 14085
0 14087 5 1 1 14086
0 14088 7 10 2 64481 65114
0 14089 7 2 2 70289 91276
0 14090 7 1 2 91286 87970
0 14091 7 1 2 14087 14090
0 14092 5 1 1 14091
0 14093 7 1 2 78548 86684
0 14094 5 1 1 14093
0 14095 7 1 2 69339 83267
0 14096 7 1 2 80316 14095
0 14097 5 1 1 14096
0 14098 7 1 2 14094 14097
0 14099 5 1 1 14098
0 14100 7 2 2 67977 82419
0 14101 7 1 2 89160 91288
0 14102 7 1 2 14099 14101
0 14103 5 1 1 14102
0 14104 7 1 2 14092 14103
0 14105 5 1 1 14104
0 14106 7 1 2 67652 14105
0 14107 5 1 1 14106
0 14108 7 1 2 70891 73788
0 14109 7 1 2 89161 14108
0 14110 7 1 2 88807 86082
0 14111 7 1 2 14109 14110
0 14112 5 1 1 14111
0 14113 7 1 2 14107 14112
0 14114 5 1 1 14113
0 14115 7 1 2 61817 14114
0 14116 5 1 1 14115
0 14117 7 1 2 81810 76916
0 14118 7 2 2 77811 77422
0 14119 7 1 2 83711 91290
0 14120 7 1 2 14117 14119
0 14121 5 1 1 14120
0 14122 7 1 2 14116 14121
0 14123 5 1 1 14122
0 14124 7 1 2 69534 14123
0 14125 5 1 1 14124
0 14126 7 1 2 14072 14125
0 14127 5 1 1 14126
0 14128 7 1 2 73408 14127
0 14129 5 1 1 14128
0 14130 7 1 2 91263 79558
0 14131 5 1 1 14130
0 14132 7 3 2 61512 90184
0 14133 5 1 1 91292
0 14134 7 3 2 82659 77194
0 14135 5 1 1 91295
0 14136 7 1 2 14133 14135
0 14137 5 16 1 14136
0 14138 7 1 2 76884 85956
0 14139 7 1 2 91298 14138
0 14140 5 1 1 14139
0 14141 7 1 2 14131 14140
0 14142 5 1 1 14141
0 14143 7 1 2 71926 14142
0 14144 5 1 1 14143
0 14145 7 1 2 85388 85952
0 14146 5 1 1 14145
0 14147 7 1 2 82974 14146
0 14148 7 1 2 91299 14147
0 14149 5 1 1 14148
0 14150 7 2 2 71661 83931
0 14151 5 1 1 91314
0 14152 7 1 2 79005 91264
0 14153 7 1 2 91315 14152
0 14154 5 1 1 14153
0 14155 7 1 2 14149 14154
0 14156 7 1 2 14144 14155
0 14157 5 1 1 14156
0 14158 7 1 2 69767 14157
0 14159 5 1 1 14158
0 14160 7 2 2 77329 80519
0 14161 7 7 2 61513 68962
0 14162 7 1 2 81756 91318
0 14163 7 1 2 91316 14162
0 14164 7 1 2 76859 14163
0 14165 5 1 1 14164
0 14166 7 2 2 71050 84945
0 14167 7 6 2 68135 65375
0 14168 7 1 2 77229 91327
0 14169 7 1 2 72287 14168
0 14170 7 1 2 91325 14169
0 14171 5 1 1 14170
0 14172 7 1 2 14165 14171
0 14173 7 1 2 14159 14172
0 14174 5 1 1 14173
0 14175 7 1 2 71211 14174
0 14176 5 1 1 14175
0 14177 7 1 2 91156 91300
0 14178 5 1 1 14177
0 14179 7 2 2 61514 76664
0 14180 7 1 2 68136 76965
0 14181 7 1 2 91333 14180
0 14182 5 1 1 14181
0 14183 7 1 2 14178 14182
0 14184 5 1 1 14183
0 14185 7 2 2 67207 71162
0 14186 5 2 1 91335
0 14187 7 1 2 91336 82393
0 14188 7 1 2 14184 14187
0 14189 5 1 1 14188
0 14190 7 1 2 14176 14189
0 14191 5 1 1 14190
0 14192 7 1 2 79350 14191
0 14193 5 1 1 14192
0 14194 7 1 2 14129 14193
0 14195 7 1 2 14003 14194
0 14196 5 1 1 14195
0 14197 7 16 2 61345 90974
0 14198 7 4 2 87714 91339
0 14199 7 1 2 14196 91355
0 14200 5 1 1 14199
0 14201 7 1 2 13708 14200
0 14202 5 1 1 14201
0 14203 7 1 2 75795 14202
0 14204 5 1 1 14203
0 14205 7 1 2 90168 86093
0 14206 7 1 2 84717 14205
0 14207 7 6 2 62539 67839
0 14208 7 13 2 61262 66207
0 14209 7 1 2 91359 91365
0 14210 7 8 2 61515 67763
0 14211 5 1 1 91378
0 14212 7 9 2 69169 69340
0 14213 7 1 2 91379 91386
0 14214 7 1 2 14209 14213
0 14215 7 1 2 64097 82660
0 14216 7 1 2 80499 14215
0 14217 7 1 2 14214 14216
0 14218 7 1 2 14206 14217
0 14219 5 1 1 14218
0 14220 7 1 2 14204 14219
0 14221 7 1 2 13623 14220
0 14222 7 1 2 13201 14221
0 14223 7 1 2 8431 14222
0 14224 5 1 1 14223
0 14225 7 1 2 64241 14224
0 14226 5 1 1 14225
0 14227 7 1 2 80087 79540
0 14228 5 1 1 14227
0 14229 7 2 2 62802 74486
0 14230 5 1 1 91395
0 14231 7 1 2 78871 91396
0 14232 5 1 1 14231
0 14233 7 1 2 14228 14232
0 14234 5 1 1 14233
0 14235 7 1 2 62540 14234
0 14236 5 1 1 14235
0 14237 7 2 2 62371 81513
0 14238 7 2 2 70290 80456
0 14239 7 1 2 91397 91399
0 14240 5 1 1 14239
0 14241 7 1 2 14236 14240
0 14242 5 1 1 14241
0 14243 7 1 2 68600 14242
0 14244 5 1 1 14243
0 14245 7 1 2 89056 90371
0 14246 5 1 1 14245
0 14247 7 1 2 78917 74588
0 14248 5 1 1 14247
0 14249 7 1 2 14246 14248
0 14250 5 1 1 14249
0 14251 7 1 2 71212 14250
0 14252 5 1 1 14251
0 14253 7 1 2 14244 14252
0 14254 5 1 1 14253
0 14255 7 1 2 65703 14254
0 14256 5 1 1 14255
0 14257 7 2 2 77965 73683
0 14258 5 1 1 91401
0 14259 7 1 2 88497 14258
0 14260 5 2 1 14259
0 14261 7 1 2 75525 91403
0 14262 5 2 1 14261
0 14263 7 2 2 67208 75511
0 14264 5 1 1 91407
0 14265 7 1 2 62372 77724
0 14266 5 1 1 14265
0 14267 7 1 2 14264 14266
0 14268 5 1 1 14267
0 14269 7 1 2 62803 14268
0 14270 5 1 1 14269
0 14271 7 1 2 91405 14270
0 14272 5 1 1 14271
0 14273 7 3 2 65376 78872
0 14274 7 1 2 14272 91409
0 14275 5 1 1 14274
0 14276 7 2 2 70654 80044
0 14277 7 4 2 70291 71015
0 14278 5 1 1 91414
0 14279 7 1 2 67978 77572
0 14280 7 1 2 91415 14279
0 14281 7 1 2 91412 14280
0 14282 5 1 1 14281
0 14283 7 1 2 14275 14282
0 14284 7 1 2 14256 14283
0 14285 5 1 1 14284
0 14286 7 1 2 66420 14285
0 14287 5 1 1 14286
0 14288 7 1 2 73409 75986
0 14289 5 1 1 14288
0 14290 7 2 2 74002 91098
0 14291 5 21 1 91418
0 14292 7 3 2 79499 91420
0 14293 5 1 1 91441
0 14294 7 1 2 14289 14293
0 14295 5 1 1 14294
0 14296 7 1 2 62804 14295
0 14297 5 1 1 14296
0 14298 7 1 2 71301 75987
0 14299 5 1 1 14298
0 14300 7 1 2 75946 87946
0 14301 5 1 1 14300
0 14302 7 1 2 14299 14301
0 14303 5 1 1 14302
0 14304 7 1 2 75526 14303
0 14305 5 1 1 14304
0 14306 7 1 2 14297 14305
0 14307 5 1 1 14306
0 14308 7 1 2 89080 14307
0 14309 5 1 1 14308
0 14310 7 1 2 14287 14309
0 14311 5 1 1 14310
0 14312 7 1 2 69341 14311
0 14313 5 1 1 14312
0 14314 7 5 2 80781 79351
0 14315 5 1 1 91444
0 14316 7 6 2 63117 70892
0 14317 7 1 2 73985 91449
0 14318 7 1 2 91445 14317
0 14319 5 1 1 14318
0 14320 7 1 2 78375 80106
0 14321 5 1 1 14320
0 14322 7 1 2 2688 14321
0 14323 5 1 1 14322
0 14324 7 1 2 82110 74530
0 14325 7 1 2 14323 14324
0 14326 5 1 1 14325
0 14327 7 1 2 14319 14326
0 14328 5 1 1 14327
0 14329 7 1 2 79901 14328
0 14330 5 1 1 14329
0 14331 7 3 2 69535 84009
0 14332 7 1 2 77230 77764
0 14333 7 1 2 84431 14332
0 14334 7 1 2 91455 14333
0 14335 5 1 1 14334
0 14336 7 1 2 14330 14335
0 14337 7 1 2 14313 14336
0 14338 5 1 1 14337
0 14339 7 1 2 68362 14338
0 14340 5 1 1 14339
0 14341 7 1 2 90762 85002
0 14342 7 4 2 64482 86759
0 14343 7 2 2 63520 82523
0 14344 7 1 2 91458 91462
0 14345 7 1 2 14341 14344
0 14346 5 1 1 14345
0 14347 7 1 2 14340 14346
0 14348 5 1 1 14347
0 14349 7 1 2 68137 14348
0 14350 5 1 1 14349
0 14351 7 3 2 80323 83937
0 14352 5 1 1 91464
0 14353 7 2 2 67979 91465
0 14354 7 1 2 84602 91467
0 14355 5 1 1 14354
0 14356 7 1 2 70655 88389
0 14357 5 1 1 14356
0 14358 7 2 2 70292 76075
0 14359 7 2 2 69536 91469
0 14360 5 1 1 91471
0 14361 7 1 2 14357 14360
0 14362 5 1 1 14361
0 14363 7 1 2 71302 14362
0 14364 5 1 1 14363
0 14365 7 4 2 67980 81243
0 14366 5 2 1 91473
0 14367 7 1 2 78901 91477
0 14368 5 1 1 14367
0 14369 7 2 2 61516 14368
0 14370 5 1 1 91479
0 14371 7 5 2 66421 81469
0 14372 5 1 1 91481
0 14373 7 1 2 78444 91482
0 14374 5 1 1 14373
0 14375 7 1 2 14370 14374
0 14376 5 1 1 14375
0 14377 7 1 2 84603 14376
0 14378 5 1 1 14377
0 14379 7 4 2 78751 87479
0 14380 7 1 2 87106 91486
0 14381 5 1 1 14380
0 14382 7 1 2 14378 14381
0 14383 7 1 2 14364 14382
0 14384 5 1 1 14383
0 14385 7 1 2 64483 14384
0 14386 5 1 1 14385
0 14387 7 1 2 14355 14386
0 14388 5 1 1 14387
0 14389 7 1 2 65958 14388
0 14390 5 1 1 14389
0 14391 7 2 2 80197 80724
0 14392 7 1 2 90857 80256
0 14393 7 1 2 91490 14392
0 14394 5 1 1 14393
0 14395 7 1 2 14390 14394
0 14396 5 1 1 14395
0 14397 7 1 2 88221 14396
0 14398 5 1 1 14397
0 14399 7 1 2 14350 14398
0 14400 5 1 1 14399
0 14401 7 1 2 61818 14400
0 14402 5 1 1 14401
0 14403 7 1 2 78944 83938
0 14404 5 1 1 14403
0 14405 7 1 2 83257 14404
0 14406 5 2 1 14405
0 14407 7 2 2 68812 74617
0 14408 7 1 2 82210 89707
0 14409 7 1 2 91494 14408
0 14410 7 1 2 91492 14409
0 14411 5 1 1 14410
0 14412 7 1 2 14402 14411
0 14413 5 1 1 14412
0 14414 7 1 2 70004 14413
0 14415 5 1 1 14414
0 14416 7 3 2 66681 65377
0 14417 7 2 2 67653 82427
0 14418 7 1 2 89535 91499
0 14419 5 1 1 14418
0 14420 7 1 2 79352 87971
0 14421 7 1 2 90744 14420
0 14422 5 2 1 14421
0 14423 7 1 2 14419 91501
0 14424 5 1 1 14423
0 14425 7 1 2 61517 14424
0 14426 5 1 1 14425
0 14427 7 1 2 82428 80457
0 14428 5 2 1 14427
0 14429 7 1 2 88222 80257
0 14430 5 1 1 14429
0 14431 7 1 2 91503 14430
0 14432 5 1 1 14431
0 14433 7 1 2 83939 14432
0 14434 5 1 1 14433
0 14435 7 1 2 14426 14434
0 14436 5 1 1 14435
0 14437 7 1 2 67412 14436
0 14438 5 1 1 14437
0 14439 7 1 2 83973 4410
0 14440 5 5 1 14439
0 14441 7 1 2 81622 80369
0 14442 7 1 2 91505 14441
0 14443 5 1 1 14442
0 14444 7 1 2 14438 14443
0 14445 5 1 1 14444
0 14446 7 1 2 63118 14445
0 14447 5 1 1 14446
0 14448 7 12 2 61518 69342
0 14449 7 1 2 82409 91510
0 14450 7 1 2 88695 14449
0 14451 7 1 2 91198 14450
0 14452 5 1 1 14451
0 14453 7 1 2 14447 14452
0 14454 5 1 1 14453
0 14455 7 1 2 91496 14454
0 14456 5 1 1 14455
0 14457 7 2 2 89257 87590
0 14458 7 4 2 62373 81757
0 14459 7 1 2 74029 87491
0 14460 7 1 2 91524 14459
0 14461 7 1 2 91522 14460
0 14462 5 1 1 14461
0 14463 7 1 2 14456 14462
0 14464 5 1 1 14463
0 14465 7 1 2 78036 14464
0 14466 5 1 1 14465
0 14467 7 1 2 64908 14466
0 14468 7 1 2 14415 14467
0 14469 5 1 1 14468
0 14470 7 3 2 66422 78775
0 14471 5 1 1 91528
0 14472 7 1 2 87012 14471
0 14473 5 2 1 14472
0 14474 7 5 2 72992 85073
0 14475 7 1 2 79772 91533
0 14476 5 1 1 14475
0 14477 7 1 2 87390 79508
0 14478 5 1 1 14477
0 14479 7 1 2 14476 14478
0 14480 5 1 1 14479
0 14481 7 1 2 91531 14480
0 14482 5 1 1 14481
0 14483 7 5 2 62805 78499
0 14484 7 3 2 76819 81891
0 14485 7 1 2 91538 91543
0 14486 5 1 1 14485
0 14487 7 1 2 14482 14486
0 14488 5 1 1 14487
0 14489 7 1 2 63290 14488
0 14490 5 1 1 14489
0 14491 7 3 2 66423 76761
0 14492 7 1 2 86088 91546
0 14493 5 1 1 14492
0 14494 7 2 2 66682 80626
0 14495 7 1 2 91534 91549
0 14496 5 1 1 14495
0 14497 7 1 2 14493 14496
0 14498 5 1 1 14497
0 14499 7 1 2 69537 81325
0 14500 7 1 2 14498 14499
0 14501 5 1 1 14500
0 14502 7 1 2 14490 14501
0 14503 5 1 1 14502
0 14504 7 1 2 70005 14503
0 14505 5 1 1 14504
0 14506 7 1 2 63757 88014
0 14507 5 1 1 14506
0 14508 7 4 2 63521 87062
0 14509 7 1 2 71619 91551
0 14510 7 1 2 87700 14509
0 14511 7 1 2 14507 14510
0 14512 5 1 1 14511
0 14513 7 1 2 14505 14512
0 14514 5 1 1 14513
0 14515 7 1 2 63119 14514
0 14516 5 1 1 14515
0 14517 7 3 2 77061 76364
0 14518 5 1 1 91555
0 14519 7 3 2 72993 73410
0 14520 5 3 1 91558
0 14521 7 3 2 67654 91559
0 14522 5 1 1 91564
0 14523 7 1 2 78104 91565
0 14524 5 1 1 14523
0 14525 7 1 2 14518 14524
0 14526 5 1 1 14525
0 14527 7 1 2 65704 14526
0 14528 5 1 1 14527
0 14529 7 2 2 80705 74793
0 14530 5 1 1 91567
0 14531 7 1 2 14528 14530
0 14532 5 1 1 14531
0 14533 7 1 2 63291 14532
0 14534 5 1 1 14533
0 14535 7 1 2 83543 78376
0 14536 7 1 2 87435 14535
0 14537 5 1 1 14536
0 14538 7 1 2 14534 14537
0 14539 5 1 1 14538
0 14540 7 1 2 61819 14539
0 14541 5 1 1 14540
0 14542 7 1 2 83676 78377
0 14543 7 1 2 87391 14542
0 14544 5 1 1 14543
0 14545 7 1 2 14541 14544
0 14546 5 1 1 14545
0 14547 7 1 2 69538 76041
0 14548 7 1 2 14546 14547
0 14549 5 1 1 14548
0 14550 7 1 2 14516 14549
0 14551 5 1 1 14550
0 14552 7 1 2 65959 14551
0 14553 5 1 1 14552
0 14554 7 3 2 74266 73411
0 14555 5 1 1 91569
0 14556 7 1 2 63292 80833
0 14557 7 2 2 91570 14556
0 14558 5 1 1 91572
0 14559 7 1 2 76665 91573
0 14560 5 1 1 14559
0 14561 7 2 2 74794 79926
0 14562 7 1 2 91301 91574
0 14563 5 1 1 14562
0 14564 7 1 2 14560 14563
0 14565 5 1 1 14564
0 14566 7 1 2 62806 81340
0 14567 7 1 2 14565 14566
0 14568 5 1 1 14567
0 14569 7 1 2 74952 76583
0 14570 7 7 2 64679 83285
0 14571 7 7 2 63293 74882
0 14572 7 1 2 91576 91583
0 14573 7 1 2 14569 14572
0 14574 5 1 1 14573
0 14575 7 1 2 14568 14574
0 14576 7 1 2 14553 14575
0 14577 5 1 1 14576
0 14578 7 1 2 64484 14577
0 14579 5 1 1 14578
0 14580 7 2 2 61820 82540
0 14581 5 2 1 91590
0 14582 7 1 2 91317 91591
0 14583 5 1 1 14582
0 14584 7 2 2 75592 80458
0 14585 7 1 2 82420 78188
0 14586 7 1 2 91594 14585
0 14587 5 1 1 14586
0 14588 7 1 2 14583 14587
0 14589 5 1 1 14588
0 14590 7 1 2 62374 14589
0 14591 5 1 1 14590
0 14592 7 1 2 85818 75331
0 14593 5 3 1 14592
0 14594 7 1 2 82879 91183
0 14595 7 1 2 82466 14594
0 14596 7 1 2 91596 14595
0 14597 5 1 1 14596
0 14598 7 1 2 14591 14597
0 14599 5 1 1 14598
0 14600 7 1 2 67655 14599
0 14601 5 1 1 14600
0 14602 7 1 2 89155 81401
0 14603 7 1 2 85787 14602
0 14604 5 1 1 14603
0 14605 7 1 2 14601 14604
0 14606 5 1 1 14605
0 14607 7 1 2 68363 14606
0 14608 5 1 1 14607
0 14609 7 8 2 65705 88529
0 14610 5 1 1 91599
0 14611 7 1 2 61821 87560
0 14612 7 1 2 89350 14611
0 14613 7 1 2 91600 14612
0 14614 5 1 1 14613
0 14615 7 1 2 14608 14614
0 14616 5 1 1 14615
0 14617 7 1 2 66424 14616
0 14618 5 1 1 14617
0 14619 7 2 2 82410 86258
0 14620 7 1 2 80782 82736
0 14621 7 1 2 84917 14620
0 14622 7 1 2 91607 14621
0 14623 5 1 1 14622
0 14624 7 1 2 14618 14623
0 14625 5 1 1 14624
0 14626 7 1 2 84074 14625
0 14627 5 1 1 14626
0 14628 7 1 2 14579 14627
0 14629 5 1 1 14628
0 14630 7 1 2 70293 14629
0 14631 5 1 1 14630
0 14632 7 1 2 81296 91535
0 14633 5 1 1 14632
0 14634 7 3 2 62807 73200
0 14635 5 5 1 91609
0 14636 7 1 2 62541 90307
0 14637 5 2 1 14636
0 14638 7 1 2 91612 91617
0 14639 5 3 1 14638
0 14640 7 3 2 70006 91619
0 14641 7 1 2 90930 91622
0 14642 5 1 1 14641
0 14643 7 1 2 14633 14642
0 14644 5 1 1 14643
0 14645 7 1 2 63522 14644
0 14646 5 1 1 14645
0 14647 7 3 2 65115 71571
0 14648 7 4 2 85548 91625
0 14649 7 6 2 63758 76396
0 14650 5 1 1 91632
0 14651 7 1 2 63294 91633
0 14652 7 1 2 91628 14651
0 14653 5 1 1 14652
0 14654 7 1 2 14646 14653
0 14655 5 1 1 14654
0 14656 7 1 2 78873 14655
0 14657 5 1 1 14656
0 14658 7 2 2 88297 91620
0 14659 7 2 2 89207 91638
0 14660 7 1 2 80441 91640
0 14661 5 1 1 14660
0 14662 7 1 2 14657 14661
0 14663 5 1 1 14662
0 14664 7 1 2 61822 14663
0 14665 5 1 1 14664
0 14666 7 1 2 89738 80416
0 14667 7 1 2 91623 14666
0 14668 5 1 1 14667
0 14669 7 1 2 14665 14668
0 14670 5 1 1 14669
0 14671 7 1 2 61519 14670
0 14672 5 1 1 14671
0 14673 7 1 2 62375 83195
0 14674 7 1 2 91641 14673
0 14675 5 1 1 14674
0 14676 7 1 2 14672 14675
0 14677 5 1 1 14676
0 14678 7 1 2 88732 14677
0 14679 5 1 1 14678
0 14680 7 2 2 79353 85914
0 14681 7 1 2 82146 91642
0 14682 5 1 1 14681
0 14683 7 7 2 69343 70656
0 14684 7 1 2 68138 78984
0 14685 7 1 2 91644 14684
0 14686 7 1 2 89047 14685
0 14687 5 1 1 14686
0 14688 7 1 2 14682 14687
0 14689 5 1 1 14688
0 14690 7 1 2 76135 14689
0 14691 5 1 1 14690
0 14692 7 1 2 68364 75202
0 14693 5 1 1 14692
0 14694 7 1 2 83843 14693
0 14695 5 1 1 14694
0 14696 7 2 2 68365 84618
0 14697 5 1 1 91651
0 14698 7 1 2 81081 14697
0 14699 5 1 1 14698
0 14700 7 1 2 14695 14699
0 14701 5 1 1 14700
0 14702 7 1 2 89344 84973
0 14703 7 1 2 14701 14702
0 14704 5 1 1 14703
0 14705 7 1 2 14691 14704
0 14706 5 1 1 14705
0 14707 7 1 2 67209 14706
0 14708 5 1 1 14707
0 14709 7 1 2 67210 77972
0 14710 5 2 1 14709
0 14711 7 1 2 71026 91653
0 14712 5 1 1 14711
0 14713 7 1 2 62376 85450
0 14714 5 1 1 14713
0 14715 7 1 2 91613 14714
0 14716 7 1 2 14712 14715
0 14717 5 1 1 14716
0 14718 7 1 2 68601 14717
0 14719 5 1 1 14718
0 14720 7 1 2 85093 14719
0 14721 5 1 1 14720
0 14722 7 4 2 83831 89345
0 14723 7 1 2 68366 91655
0 14724 7 1 2 14721 14723
0 14725 5 1 1 14724
0 14726 7 1 2 14708 14725
0 14727 5 1 1 14726
0 14728 7 1 2 70007 14727
0 14729 5 1 1 14728
0 14730 7 5 2 64680 71303
0 14731 7 3 2 70657 91659
0 14732 7 4 2 81697 80411
0 14733 7 1 2 91664 91667
0 14734 5 1 1 14733
0 14735 7 1 2 79354 80645
0 14736 5 1 1 14735
0 14737 7 5 2 69344 80258
0 14738 7 1 2 80222 91671
0 14739 5 1 1 14738
0 14740 7 1 2 14736 14739
0 14741 5 1 1 14740
0 14742 7 1 2 81553 79474
0 14743 7 1 2 14741 14742
0 14744 5 1 1 14743
0 14745 7 1 2 14734 14744
0 14746 5 1 1 14745
0 14747 7 1 2 68602 14746
0 14748 5 1 1 14747
0 14749 7 1 2 80259 81529
0 14750 7 1 2 87656 14749
0 14751 5 1 1 14750
0 14752 7 1 2 61520 14751
0 14753 7 1 2 14748 14752
0 14754 5 1 1 14753
0 14755 7 1 2 82867 91404
0 14756 5 1 1 14755
0 14757 7 4 2 67211 81554
0 14758 7 1 2 91199 91676
0 14759 5 1 1 14758
0 14760 7 1 2 14756 14759
0 14761 5 1 1 14760
0 14762 7 1 2 83241 14761
0 14763 5 1 1 14762
0 14764 7 1 2 68139 88076
0 14765 7 1 2 89539 14764
0 14766 5 1 1 14765
0 14767 7 1 2 63295 90814
0 14768 7 1 2 86779 14767
0 14769 5 1 1 14768
0 14770 7 1 2 14766 14769
0 14771 5 1 1 14770
0 14772 7 1 2 63120 14771
0 14773 5 1 1 14772
0 14774 7 1 2 66425 14773
0 14775 7 1 2 14763 14774
0 14776 5 1 1 14775
0 14777 7 1 2 76292 14776
0 14778 7 1 2 14754 14777
0 14779 5 1 1 14778
0 14780 7 1 2 14729 14779
0 14781 5 1 1 14780
0 14782 7 1 2 65960 14781
0 14783 5 1 1 14782
0 14784 7 1 2 72949 85218
0 14785 5 5 1 14784
0 14786 7 1 2 80715 78124
0 14787 5 19 1 14786
0 14788 7 2 2 65961 91685
0 14789 7 2 2 81029 91704
0 14790 7 1 2 91656 91706
0 14791 5 1 1 14790
0 14792 7 2 2 68140 73696
0 14793 7 3 2 80967 91708
0 14794 7 1 2 77812 81341
0 14795 7 1 2 84209 14794
0 14796 7 2 2 91710 14795
0 14797 5 1 1 91713
0 14798 7 1 2 14791 14797
0 14799 5 1 1 14798
0 14800 7 1 2 91680 14799
0 14801 5 1 1 14800
0 14802 7 1 2 62377 73412
0 14803 5 1 1 14802
0 14804 7 2 2 62542 77355
0 14805 5 4 1 91715
0 14806 7 1 2 14803 91717
0 14807 5 1 1 14806
0 14808 7 1 2 68603 14807
0 14809 5 1 1 14808
0 14810 7 1 2 67413 71622
0 14811 5 1 1 14810
0 14812 7 1 2 14809 14811
0 14813 5 1 1 14812
0 14814 7 5 2 69345 80198
0 14815 7 1 2 79749 90912
0 14816 7 1 2 91721 14815
0 14817 7 1 2 14813 14816
0 14818 5 1 1 14817
0 14819 7 1 2 14801 14818
0 14820 7 1 2 14783 14819
0 14821 5 1 1 14820
0 14822 7 1 2 65378 14821
0 14823 5 1 1 14822
0 14824 7 3 2 67656 72271
0 14825 5 2 1 91726
0 14826 7 1 2 72353 91729
0 14827 5 4 1 14826
0 14828 7 1 2 83688 90807
0 14829 5 1 1 14828
0 14830 7 2 2 91085 91302
0 14831 7 1 2 86522 91735
0 14832 5 1 1 14831
0 14833 7 1 2 14829 14832
0 14834 5 1 1 14833
0 14835 7 1 2 79387 14834
0 14836 5 1 1 14835
0 14837 7 3 2 68367 81730
0 14838 7 2 2 89930 91737
0 14839 7 1 2 79435 77918
0 14840 7 1 2 91547 14839
0 14841 7 1 2 91740 14840
0 14842 5 1 1 14841
0 14843 7 1 2 14836 14842
0 14844 5 1 1 14843
0 14845 7 1 2 91731 14844
0 14846 5 1 1 14845
0 14847 7 1 2 69768 14846
0 14848 7 1 2 14823 14847
0 14849 7 1 2 14679 14848
0 14850 7 1 2 14631 14849
0 14851 5 1 1 14850
0 14852 7 1 2 67764 14851
0 14853 7 1 2 14469 14852
0 14854 5 1 1 14853
0 14855 7 3 2 67212 62944
0 14856 7 1 2 81530 91742
0 14857 7 1 2 88775 14856
0 14858 7 5 2 74618 79295
0 14859 7 1 2 79326 91745
0 14860 7 1 2 14857 14859
0 14861 5 1 1 14860
0 14862 7 1 2 14854 14861
0 14863 5 1 1 14862
0 14864 7 1 2 90649 14863
0 14865 5 1 1 14864
0 14866 7 3 2 86259 85653
0 14867 7 1 2 84188 91750
0 14868 5 1 1 14867
0 14869 7 3 2 70294 79355
0 14870 7 2 2 81623 91753
0 14871 5 1 1 91756
0 14872 7 1 2 14868 14871
0 14873 5 1 1 14872
0 14874 7 1 2 61521 14873
0 14875 5 1 1 14874
0 14876 7 2 2 85640 74935
0 14877 7 1 2 88686 90763
0 14878 7 1 2 91758 14877
0 14879 5 1 1 14878
0 14880 7 1 2 14875 14879
0 14881 5 1 1 14880
0 14882 7 1 2 67981 14881
0 14883 5 1 1 14882
0 14884 7 5 2 66426 82661
0 14885 7 1 2 80484 87492
0 14886 7 1 2 91760 14885
0 14887 5 1 1 14886
0 14888 7 1 2 14883 14887
0 14889 5 1 1 14888
0 14890 7 1 2 72765 14889
0 14891 5 1 1 14890
0 14892 7 4 2 82111 88115
0 14893 5 1 1 91765
0 14894 7 1 2 80199 82918
0 14895 7 1 2 91766 14894
0 14896 5 1 1 14895
0 14897 7 1 2 14891 14896
0 14898 5 1 1 14897
0 14899 7 1 2 78602 14898
0 14900 5 1 1 14899
0 14901 7 5 2 87401 79436
0 14902 5 1 1 91769
0 14903 7 2 2 81758 74030
0 14904 7 1 2 86083 91774
0 14905 7 1 2 91770 14904
0 14906 5 1 1 14905
0 14907 7 1 2 14900 14906
0 14908 5 1 1 14907
0 14909 7 1 2 67213 14908
0 14910 5 1 1 14909
0 14911 7 1 2 74531 88183
0 14912 5 1 1 14911
0 14913 7 5 2 61522 63759
0 14914 7 1 2 91410 91776
0 14915 5 1 1 14914
0 14916 7 1 2 14912 14915
0 14917 5 1 1 14916
0 14918 7 2 2 69769 78037
0 14919 7 4 2 67414 64485
0 14920 7 1 2 81624 91783
0 14921 7 1 2 91781 14920
0 14922 7 1 2 14917 14921
0 14923 5 1 1 14922
0 14924 7 1 2 14910 14923
0 14925 5 1 1 14924
0 14926 7 1 2 61823 14925
0 14927 5 1 1 14926
0 14928 7 1 2 89018 74703
0 14929 5 1 1 14928
0 14930 7 3 2 67657 80029
0 14931 7 1 2 88744 79933
0 14932 7 1 2 91787 14931
0 14933 5 1 1 14932
0 14934 7 1 2 14929 14933
0 14935 5 1 1 14934
0 14936 7 4 2 67415 78500
0 14937 7 1 2 88273 85960
0 14938 7 1 2 91790 14937
0 14939 7 1 2 14935 14938
0 14940 5 1 1 14939
0 14941 7 1 2 14927 14940
0 14942 5 1 1 14941
0 14943 7 1 2 67765 14942
0 14944 5 1 1 14943
0 14945 7 2 2 88776 87456
0 14946 7 5 2 67416 62945
0 14947 7 2 2 79934 91796
0 14948 7 1 2 78038 82983
0 14949 7 1 2 91801 14948
0 14950 7 1 2 91794 14949
0 14951 5 1 1 14950
0 14952 7 1 2 14944 14951
0 14953 5 1 1 14952
0 14954 7 1 2 90650 14953
0 14955 5 1 1 14954
0 14956 7 4 2 67766 62997
0 14957 7 1 2 81514 84432
0 14958 7 1 2 91803 14957
0 14959 7 10 2 61346 66683
0 14960 5 1 1 91807
0 14961 7 2 2 89162 91808
0 14962 7 3 2 64909 74619
0 14963 7 1 2 81044 83380
0 14964 7 1 2 91819 14963
0 14965 7 1 2 91817 14964
0 14966 7 1 2 14958 14965
0 14967 5 1 1 14966
0 14968 7 1 2 14955 14967
0 14969 5 1 1 14968
0 14970 7 1 2 73254 14969
0 14971 5 1 1 14970
0 14972 7 12 2 67982 81555
0 14973 7 4 2 87457 91822
0 14974 7 1 2 90639 84537
0 14975 7 1 2 84269 14974
0 14976 7 1 2 91834 14975
0 14977 5 1 1 14976
0 14978 7 1 2 14971 14977
0 14979 7 1 2 14865 14978
0 14980 5 1 1 14979
0 14981 7 1 2 64321 14980
0 14982 5 1 1 14981
0 14983 7 2 2 81556 84270
0 14984 7 13 2 69170 82984
0 14985 7 2 2 66684 77573
0 14986 7 1 2 91840 91853
0 14987 7 20 2 67767 67840
0 14988 7 10 2 66208 66427
0 14989 7 4 2 91855 91875
0 14990 7 5 2 67983 82524
0 14991 7 1 2 91885 91889
0 14992 7 1 2 14986 14991
0 14993 7 1 2 91838 14992
0 14994 5 1 1 14993
0 14995 7 1 2 61263 14994
0 14996 7 1 2 14982 14995
0 14997 5 1 1 14996
0 14998 7 2 2 70658 82844
0 14999 7 2 2 80847 91894
0 15000 5 1 1 91896
0 15001 7 4 2 69346 72994
0 15002 7 1 2 82757 91898
0 15003 5 1 1 15002
0 15004 7 1 2 15000 15003
0 15005 5 1 1 15004
0 15006 7 1 2 71304 15005
0 15007 5 1 1 15006
0 15008 7 2 2 80968 90901
0 15009 7 2 2 72245 91902
0 15010 5 1 1 91904
0 15011 7 1 2 75269 91905
0 15012 5 1 1 15011
0 15013 7 3 2 83806 91777
0 15014 7 1 2 85560 91906
0 15015 5 1 1 15014
0 15016 7 1 2 15012 15015
0 15017 7 1 2 15007 15016
0 15018 5 1 1 15017
0 15019 7 1 2 65116 15018
0 15020 5 1 1 15019
0 15021 7 2 2 74795 91058
0 15022 5 1 1 91909
0 15023 7 1 2 83848 91910
0 15024 5 1 1 15023
0 15025 7 1 2 15020 15024
0 15026 5 1 1 15025
0 15027 7 1 2 65962 15026
0 15028 5 1 1 15027
0 15029 7 1 2 77865 91561
0 15030 5 1 1 15029
0 15031 7 2 2 62808 15030
0 15032 5 1 1 91911
0 15033 7 1 2 80969 87467
0 15034 7 1 2 91912 15033
0 15035 5 1 1 15034
0 15036 7 1 2 15028 15035
0 15037 5 1 1 15036
0 15038 7 1 2 64681 15037
0 15039 5 1 1 15038
0 15040 7 1 2 79013 85074
0 15041 5 1 1 15040
0 15042 7 1 2 15022 15041
0 15043 5 2 1 15042
0 15044 7 1 2 76076 91913
0 15045 5 1 1 15044
0 15046 7 1 2 82305 79576
0 15047 7 1 2 91890 15046
0 15048 5 1 1 15047
0 15049 7 1 2 15045 15048
0 15050 5 1 1 15049
0 15051 7 1 2 89442 15050
0 15052 5 1 1 15051
0 15053 7 1 2 15039 15052
0 15054 5 1 1 15053
0 15055 7 1 2 81411 15054
0 15056 5 1 1 15055
0 15057 7 2 2 78549 79968
0 15058 7 4 2 80783 81759
0 15059 7 2 2 77574 81531
0 15060 7 1 2 91917 91921
0 15061 7 1 2 91915 15060
0 15062 5 1 1 15061
0 15063 7 1 2 63523 15062
0 15064 7 1 2 15056 15063
0 15065 5 1 1 15064
0 15066 7 1 2 91406 15032
0 15067 5 1 1 15066
0 15068 7 2 2 76136 81276
0 15069 7 1 2 15067 91923
0 15070 5 1 1 15069
0 15071 7 1 2 87642 82947
0 15072 7 1 2 77787 15071
0 15073 5 1 1 15072
0 15074 7 1 2 15070 15073
0 15075 5 1 1 15074
0 15076 7 1 2 69347 15075
0 15077 5 1 1 15076
0 15078 7 1 2 77804 5333
0 15079 5 1 1 15078
0 15080 7 1 2 68604 15079
0 15081 5 1 1 15080
0 15082 7 1 2 74796 73943
0 15083 5 2 1 15082
0 15084 7 1 2 71305 71927
0 15085 7 1 2 91925 15084
0 15086 5 1 1 15085
0 15087 7 1 2 85094 15086
0 15088 7 1 2 15081 15087
0 15089 5 1 1 15088
0 15090 7 1 2 88838 81412
0 15091 7 1 2 15089 15090
0 15092 5 1 1 15091
0 15093 7 1 2 15077 15092
0 15094 5 1 1 15093
0 15095 7 1 2 64682 15094
0 15096 5 1 1 15095
0 15097 7 1 2 71504 85974
0 15098 5 3 1 15097
0 15099 7 2 2 81277 91450
0 15100 5 2 1 91930
0 15101 7 1 2 91446 91931
0 15102 7 1 2 91927 15101
0 15103 5 1 1 15102
0 15104 7 1 2 15096 15103
0 15105 5 1 1 15104
0 15106 7 1 2 70008 15105
0 15107 5 1 1 15106
0 15108 7 1 2 71213 91493
0 15109 5 1 1 15108
0 15110 7 2 2 80223 82433
0 15111 7 1 2 87354 91934
0 15112 5 1 1 15111
0 15113 7 1 2 15109 15112
0 15114 5 2 1 15113
0 15115 7 1 2 89107 71692
0 15116 7 1 2 77878 15115
0 15117 7 1 2 91936 15116
0 15118 5 1 1 15117
0 15119 7 1 2 68368 15118
0 15120 7 1 2 15107 15119
0 15121 5 1 1 15120
0 15122 7 1 2 61824 15121
0 15123 7 1 2 15065 15122
0 15124 5 1 1 15123
0 15125 7 1 2 61523 78945
0 15126 5 1 1 15125
0 15127 7 1 2 14372 15126
0 15128 5 11 1 15127
0 15129 7 7 2 67214 71214
0 15130 5 1 1 91949
0 15131 7 4 2 82715 91950
0 15132 7 1 2 91938 91956
0 15133 5 1 1 15132
0 15134 7 6 2 66428 90026
0 15135 7 1 2 74267 82541
0 15136 7 1 2 91960 15135
0 15137 5 1 1 15136
0 15138 7 3 2 82716 80088
0 15139 5 1 1 91966
0 15140 7 1 2 89258 91967
0 15141 5 1 1 15140
0 15142 7 1 2 15137 15141
0 15143 5 1 1 15142
0 15144 7 1 2 85075 15143
0 15145 5 1 1 15144
0 15146 7 1 2 15133 15145
0 15147 5 1 1 15146
0 15148 7 1 2 65117 15147
0 15149 5 1 1 15148
0 15150 7 3 2 66429 78946
0 15151 5 1 1 91969
0 15152 7 1 2 89091 15151
0 15153 5 9 1 15152
0 15154 7 5 2 70009 81625
0 15155 7 4 2 85706 79475
0 15156 5 1 1 91986
0 15157 7 1 2 91981 91987
0 15158 7 1 2 91972 15157
0 15159 5 1 1 15158
0 15160 7 1 2 15149 15159
0 15161 5 1 1 15160
0 15162 7 1 2 64910 15161
0 15163 5 1 1 15162
0 15164 7 1 2 76137 86451
0 15165 7 2 2 63760 82411
0 15166 7 1 2 82034 91990
0 15167 7 1 2 15164 15166
0 15168 5 1 1 15167
0 15169 7 1 2 15163 15168
0 15170 5 1 1 15169
0 15171 7 1 2 84226 15170
0 15172 5 1 1 15171
0 15173 7 5 2 64911 77231
0 15174 7 1 2 82451 91992
0 15175 7 1 2 91914 15174
0 15176 5 1 1 15175
0 15177 7 1 2 15172 15176
0 15178 5 1 1 15177
0 15179 7 1 2 75584 15178
0 15180 5 1 1 15179
0 15181 7 1 2 82253 91707
0 15182 5 1 1 15181
0 15183 7 1 2 82602 78189
0 15184 7 1 2 90097 15183
0 15185 5 1 1 15184
0 15186 7 1 2 15182 15185
0 15187 5 1 1 15186
0 15188 7 1 2 63121 15187
0 15189 5 1 1 15188
0 15190 7 3 2 69770 79296
0 15191 7 2 2 80970 88913
0 15192 7 2 2 75450 92000
0 15193 7 1 2 91997 92002
0 15194 5 1 1 15193
0 15195 7 1 2 15189 15194
0 15196 5 1 1 15195
0 15197 7 1 2 83329 15196
0 15198 5 1 1 15197
0 15199 7 1 2 69771 91714
0 15200 5 1 1 15199
0 15201 7 1 2 15198 15200
0 15202 5 1 1 15201
0 15203 7 1 2 91681 15202
0 15204 5 1 1 15203
0 15205 7 1 2 65379 15204
0 15206 7 1 2 15180 15205
0 15207 7 1 2 15124 15206
0 15208 5 1 1 15207
0 15209 7 2 2 82236 91303
0 15210 5 1 1 92004
0 15211 7 1 2 80760 92005
0 15212 5 1 1 15211
0 15213 7 4 2 64912 83045
0 15214 7 8 2 66430 84075
0 15215 7 1 2 92006 92010
0 15216 5 1 1 15215
0 15217 7 1 2 15210 15216
0 15218 5 1 1 15217
0 15219 7 1 2 71928 85869
0 15220 7 1 2 15218 15219
0 15221 5 1 1 15220
0 15222 7 1 2 15212 15221
0 15223 5 1 1 15222
0 15224 7 1 2 85790 15223
0 15225 5 1 1 15224
0 15226 7 1 2 64486 89923
0 15227 7 1 2 83513 15226
0 15228 7 1 2 83689 15227
0 15229 5 1 1 15228
0 15230 7 1 2 15225 15229
0 15231 5 1 1 15230
0 15232 7 1 2 69539 15231
0 15233 5 1 1 15232
0 15234 7 8 2 66431 69772
0 15235 7 1 2 78258 92018
0 15236 7 1 2 83572 15235
0 15237 5 1 1 15236
0 15238 7 4 2 81840 84464
0 15239 5 1 1 92026
0 15240 7 1 2 88503 79639
0 15241 7 1 2 92027 15240
0 15242 5 1 1 15241
0 15243 7 1 2 15237 15242
0 15244 5 1 1 15243
0 15245 7 1 2 71306 15244
0 15246 5 1 1 15245
0 15247 7 2 2 82369 87276
0 15248 7 4 2 64683 74965
0 15249 7 1 2 63761 83394
0 15250 7 1 2 92032 15249
0 15251 7 1 2 92030 15250
0 15252 5 1 1 15251
0 15253 7 1 2 15246 15252
0 15254 7 1 2 15233 15253
0 15255 5 1 1 15254
0 15256 7 1 2 67658 15255
0 15257 5 1 1 15256
0 15258 7 3 2 79121 78501
0 15259 5 4 1 92036
0 15260 7 4 2 61825 79074
0 15261 7 1 2 66432 92043
0 15262 5 1 1 15261
0 15263 7 1 2 92039 15262
0 15264 5 7 1 15263
0 15265 7 2 2 67215 80224
0 15266 7 2 2 84210 82421
0 15267 7 1 2 92054 92056
0 15268 5 1 1 15267
0 15269 7 1 2 83573 15268
0 15270 5 2 1 15269
0 15271 7 1 2 70659 92058
0 15272 5 1 1 15271
0 15273 7 2 2 87643 83646
0 15274 7 1 2 90027 82893
0 15275 7 1 2 92060 15274
0 15276 5 1 1 15275
0 15277 7 1 2 15272 15276
0 15278 5 1 1 15277
0 15279 7 1 2 92047 15278
0 15280 5 1 1 15279
0 15281 7 1 2 88993 82959
0 15282 7 1 2 91480 15281
0 15283 5 1 1 15282
0 15284 7 1 2 80761 91657
0 15285 5 1 1 15284
0 15286 7 1 2 82154 88808
0 15287 7 1 2 90559 15286
0 15288 5 1 1 15287
0 15289 7 1 2 15285 15288
0 15290 5 1 1 15289
0 15291 7 8 2 69773 73413
0 15292 7 1 2 68369 92062
0 15293 7 1 2 15290 15292
0 15294 5 1 1 15293
0 15295 7 1 2 15283 15294
0 15296 7 1 2 15280 15295
0 15297 7 1 2 15257 15296
0 15298 5 1 1 15297
0 15299 7 1 2 65963 15298
0 15300 5 1 1 15299
0 15301 7 1 2 76994 89886
0 15302 7 1 2 88530 15301
0 15303 5 1 1 15302
0 15304 7 1 2 82259 2070
0 15305 5 1 1 15304
0 15306 7 1 2 88704 71479
0 15307 7 1 2 15305 15306
0 15308 5 1 1 15307
0 15309 7 1 2 15303 15308
0 15310 5 1 1 15309
0 15311 7 1 2 66433 15310
0 15312 5 1 1 15311
0 15313 7 1 2 85860 82237
0 15314 7 1 2 88526 15313
0 15315 7 1 2 91293 15314
0 15316 5 1 1 15315
0 15317 7 1 2 15312 15316
0 15318 5 1 1 15317
0 15319 7 1 2 69540 15318
0 15320 5 1 1 15319
0 15321 7 1 2 89163 80848
0 15322 5 1 1 15321
0 15323 7 1 2 71215 89181
0 15324 5 1 1 15323
0 15325 7 1 2 15322 15324
0 15326 5 1 1 15325
0 15327 7 1 2 89447 15326
0 15328 5 1 1 15327
0 15329 7 1 2 15320 15328
0 15330 5 1 1 15329
0 15331 7 1 2 65706 15330
0 15332 5 1 1 15331
0 15333 7 1 2 85241 75622
0 15334 7 3 2 64684 88687
0 15335 7 1 2 92070 92028
0 15336 7 1 2 15333 15335
0 15337 5 1 1 15336
0 15338 7 1 2 15332 15337
0 15339 5 1 1 15338
0 15340 7 1 2 68370 15339
0 15341 5 1 1 15340
0 15342 7 1 2 87657 83984
0 15343 7 3 2 66434 73414
0 15344 5 1 1 92073
0 15345 7 1 2 71788 92074
0 15346 7 1 2 15342 15345
0 15347 5 1 1 15346
0 15348 7 1 2 70010 15347
0 15349 7 1 2 15341 15348
0 15350 7 1 2 15300 15349
0 15351 5 1 1 15350
0 15352 7 2 2 82112 80200
0 15353 5 1 1 92076
0 15354 7 1 2 91601 92077
0 15355 5 1 1 15354
0 15356 7 1 2 78165 84433
0 15357 7 1 2 82357 15356
0 15358 5 1 1 15357
0 15359 7 1 2 15355 15358
0 15360 5 1 1 15359
0 15361 7 1 2 86205 81413
0 15362 7 1 2 15360 15361
0 15363 5 1 1 15362
0 15364 7 3 2 71929 85561
0 15365 5 1 1 92078
0 15366 7 1 2 74838 15365
0 15367 5 2 1 15366
0 15368 7 2 2 80485 82238
0 15369 7 1 2 91265 92083
0 15370 5 1 1 15369
0 15371 7 1 2 88925 83862
0 15372 5 1 1 15371
0 15373 7 1 2 15370 15372
0 15374 5 1 1 15373
0 15375 7 1 2 92081 15374
0 15376 5 1 1 15375
0 15377 7 1 2 91267 90753
0 15378 5 1 1 15377
0 15379 7 1 2 82758 90532
0 15380 5 1 1 15379
0 15381 7 1 2 15378 15380
0 15382 5 1 1 15381
0 15383 7 1 2 89132 73752
0 15384 7 1 2 15382 15383
0 15385 5 1 1 15384
0 15386 7 1 2 15376 15385
0 15387 5 1 1 15386
0 15388 7 1 2 65964 15387
0 15389 5 1 1 15388
0 15390 7 1 2 65118 15389
0 15391 7 1 2 15363 15390
0 15392 5 1 1 15391
0 15393 7 1 2 15351 15392
0 15394 5 1 1 15393
0 15395 7 1 2 70295 15394
0 15396 5 1 1 15395
0 15397 7 1 2 15208 15396
0 15398 5 1 1 15397
0 15399 7 1 2 78603 91536
0 15400 5 1 1 15399
0 15401 7 3 2 71817 78550
0 15402 5 1 1 92085
0 15403 7 1 2 79998 92086
0 15404 5 1 1 15403
0 15405 7 1 2 15400 15404
0 15406 5 1 1 15405
0 15407 7 1 2 78874 15406
0 15408 5 1 1 15407
0 15409 7 1 2 79075 88068
0 15410 7 1 2 91624 15409
0 15411 5 1 1 15410
0 15412 7 1 2 15408 15411
0 15413 5 1 1 15412
0 15414 7 1 2 63524 15413
0 15415 5 1 1 15414
0 15416 7 1 2 88366 79999
0 15417 5 1 1 15416
0 15418 7 1 2 73309 91474
0 15419 5 1 1 15418
0 15420 7 1 2 15417 15419
0 15421 5 1 1 15420
0 15422 7 1 2 62378 83482
0 15423 7 1 2 15421 15422
0 15424 5 1 1 15423
0 15425 7 1 2 15415 15424
0 15426 5 1 1 15425
0 15427 7 1 2 61524 15426
0 15428 5 1 1 15427
0 15429 7 1 2 87615 91961
0 15430 7 1 2 91639 15429
0 15431 5 1 1 15430
0 15432 7 1 2 15428 15431
0 15433 5 1 1 15432
0 15434 7 1 2 82370 15433
0 15435 5 1 1 15434
0 15436 7 1 2 78875 90308
0 15437 5 1 1 15436
0 15438 7 1 2 72246 91475
0 15439 5 1 1 15438
0 15440 7 1 2 15437 15439
0 15441 5 1 1 15440
0 15442 7 1 2 61525 15441
0 15443 5 1 1 15442
0 15444 7 4 2 63122 63931
0 15445 7 2 2 81244 92088
0 15446 7 1 2 80929 92092
0 15447 5 1 1 15446
0 15448 7 1 2 15443 15447
0 15449 5 1 1 15448
0 15450 7 1 2 62543 15449
0 15451 5 1 1 15450
0 15452 7 10 2 61526 78692
0 15453 7 2 2 64685 73201
0 15454 7 1 2 92094 92104
0 15455 5 1 1 15454
0 15456 7 1 2 15451 15455
0 15457 5 1 1 15456
0 15458 7 1 2 71818 81356
0 15459 7 1 2 88259 15458
0 15460 7 1 2 15457 15459
0 15461 5 1 1 15460
0 15462 7 1 2 15435 15461
0 15463 5 1 1 15462
0 15464 7 1 2 65965 15463
0 15465 5 1 1 15464
0 15466 7 2 2 65707 83690
0 15467 7 2 2 76820 77717
0 15468 5 1 1 92108
0 15469 7 1 2 81342 74236
0 15470 7 1 2 92109 15469
0 15471 7 1 2 92106 15470
0 15472 5 1 1 15471
0 15473 7 1 2 15465 15472
0 15474 5 1 1 15473
0 15475 7 1 2 64487 15474
0 15476 5 1 1 15475
0 15477 7 1 2 62379 81892
0 15478 7 1 2 80725 90858
0 15479 7 1 2 15477 15478
0 15480 7 1 2 90170 15479
0 15481 7 1 2 87616 91732
0 15482 7 1 2 15480 15481
0 15483 5 1 1 15482
0 15484 7 1 2 15476 15483
0 15485 7 1 2 15398 15484
0 15486 5 1 1 15485
0 15487 7 1 2 64322 15486
0 15488 5 1 1 15487
0 15489 7 12 2 69171 64686
0 15490 7 4 2 81532 92110
0 15491 7 1 2 89173 92122
0 15492 7 1 2 91839 15491
0 15493 5 1 1 15492
0 15494 7 1 2 15488 15493
0 15495 5 1 1 15494
0 15496 7 1 2 90699 15495
0 15497 5 1 1 15496
0 15498 7 2 2 89164 91823
0 15499 7 1 2 90099 80239
0 15500 7 1 2 92126 15499
0 15501 5 1 1 15500
0 15502 7 3 2 64488 88242
0 15503 7 2 2 77609 91778
0 15504 7 1 2 83566 92131
0 15505 7 1 2 92128 15504
0 15506 5 1 1 15505
0 15507 7 1 2 15501 15506
0 15508 5 1 1 15507
0 15509 7 1 2 67417 15508
0 15510 5 1 1 15509
0 15511 7 4 2 62544 87561
0 15512 7 1 2 83647 87107
0 15513 7 2 2 91042 15512
0 15514 7 1 2 92133 92137
0 15515 5 1 1 15514
0 15516 7 1 2 15510 15515
0 15517 5 1 1 15516
0 15518 7 1 2 66685 15517
0 15519 5 1 1 15518
0 15520 7 1 2 76995 85011
0 15521 7 1 2 92138 15520
0 15522 5 1 1 15521
0 15523 7 1 2 15519 15522
0 15524 5 1 1 15523
0 15525 7 1 2 70660 15524
0 15526 5 1 1 15525
0 15527 7 2 2 80930 80240
0 15528 5 2 1 92139
0 15529 7 1 2 63932 92140
0 15530 5 1 1 15529
0 15531 7 3 2 61527 72915
0 15532 7 1 2 88243 92143
0 15533 5 1 1 15532
0 15534 7 1 2 15530 15533
0 15535 5 1 1 15534
0 15536 7 1 2 66686 90028
0 15537 7 1 2 82861 15536
0 15538 7 1 2 86338 15537
0 15539 7 1 2 15535 15538
0 15540 5 1 1 15539
0 15541 7 1 2 15526 15540
0 15542 5 1 1 15541
0 15543 7 1 2 70011 15542
0 15544 5 1 1 15543
0 15545 7 3 2 72995 73202
0 15546 7 1 2 89053 79466
0 15547 7 1 2 84758 15546
0 15548 7 1 2 92146 15547
0 15549 5 1 1 15548
0 15550 7 1 2 15544 15549
0 15551 5 1 1 15550
0 15552 7 1 2 70296 15551
0 15553 5 1 1 15552
0 15554 7 4 2 65380 87355
0 15555 7 2 2 85915 80770
0 15556 7 1 2 76318 92153
0 15557 7 1 2 92149 15556
0 15558 7 1 2 92059 15557
0 15559 5 1 1 15558
0 15560 7 1 2 69774 15559
0 15561 7 1 2 15553 15560
0 15562 5 1 1 15561
0 15563 7 3 2 71775 74677
0 15564 7 1 2 85003 91746
0 15565 7 1 2 92155 15564
0 15566 5 1 1 15565
0 15567 7 1 2 79605 78765
0 15568 7 1 2 92147 15567
0 15569 5 1 1 15568
0 15570 7 1 2 15566 15569
0 15571 5 1 1 15570
0 15572 7 1 2 81626 84402
0 15573 7 1 2 15571 15572
0 15574 5 1 1 15573
0 15575 7 1 2 88477 79974
0 15576 7 1 2 81524 91747
0 15577 7 1 2 15575 15576
0 15578 5 1 1 15577
0 15579 7 1 2 15574 15578
0 15580 5 1 1 15579
0 15581 7 1 2 69348 15580
0 15582 5 1 1 15581
0 15583 7 4 2 70012 83330
0 15584 7 2 2 70297 86831
0 15585 7 1 2 92158 92162
0 15586 5 1 1 15585
0 15587 7 1 2 69541 89879
0 15588 7 1 2 81015 15587
0 15589 5 1 1 15588
0 15590 7 1 2 15586 15589
0 15591 5 1 1 15590
0 15592 7 1 2 88740 90001
0 15593 7 1 2 15591 15592
0 15594 5 1 1 15593
0 15595 7 1 2 64913 15594
0 15596 7 1 2 15582 15595
0 15597 5 1 1 15596
0 15598 7 23 2 67768 69172
0 15599 7 1 2 90651 92164
0 15600 7 1 2 15597 15599
0 15601 7 1 2 15562 15600
0 15602 5 1 1 15601
0 15603 7 1 2 89094 81508
0 15604 7 17 2 61347 66435
0 15605 5 1 1 92187
0 15606 7 4 2 90975 92188
0 15607 7 14 2 64323 64489
0 15608 7 3 2 81811 92208
0 15609 7 1 2 92204 92222
0 15610 7 1 2 15603 15609
0 15611 7 1 2 83725 15610
0 15612 5 1 1 15611
0 15613 7 1 2 66090 15612
0 15614 7 1 2 15602 15613
0 15615 7 1 2 15497 15614
0 15616 5 1 1 15615
0 15617 7 1 2 68963 15616
0 15618 7 1 2 14997 15617
0 15619 5 1 1 15618
0 15620 7 2 2 63762 79990
0 15621 5 1 1 92225
0 15622 7 1 2 87695 92226
0 15623 5 1 1 15622
0 15624 7 5 2 68141 78502
0 15625 7 1 2 80017 92227
0 15626 5 1 1 15625
0 15627 7 1 2 15623 15626
0 15628 5 1 1 15627
0 15629 7 1 2 67216 15628
0 15630 5 1 1 15629
0 15631 7 3 2 68605 79991
0 15632 5 1 1 92232
0 15633 7 1 2 88290 92233
0 15634 5 1 1 15633
0 15635 7 1 2 15630 15634
0 15636 5 1 1 15635
0 15637 7 1 2 64687 15636
0 15638 5 1 1 15637
0 15639 7 1 2 85641 78259
0 15640 7 1 2 91537 15639
0 15641 5 1 1 15640
0 15642 7 1 2 15638 15641
0 15643 5 1 1 15642
0 15644 7 1 2 65381 15643
0 15645 5 1 1 15644
0 15646 7 5 2 70298 83715
0 15647 5 1 1 92235
0 15648 7 2 2 67217 92236
0 15649 5 1 1 92240
0 15650 7 2 2 83381 78503
0 15651 5 1 1 92242
0 15652 7 1 2 68606 92243
0 15653 7 1 2 92241 15652
0 15654 5 1 1 15653
0 15655 7 1 2 15645 15654
0 15656 5 1 1 15655
0 15657 7 1 2 84076 15656
0 15658 5 1 1 15657
0 15659 7 1 2 71307 76430
0 15660 7 1 2 82862 15659
0 15661 7 1 2 92150 15660
0 15662 5 1 1 15661
0 15663 7 1 2 80459 86452
0 15664 7 1 2 91791 15663
0 15665 7 1 2 86348 15664
0 15666 5 1 1 15665
0 15667 7 1 2 15662 15666
0 15668 5 1 1 15667
0 15669 7 1 2 89240 15668
0 15670 5 1 1 15669
0 15671 7 1 2 15658 15670
0 15672 5 1 1 15671
0 15673 7 1 2 70893 15672
0 15674 5 1 1 15673
0 15675 7 1 2 83807 85991
0 15676 5 1 1 15675
0 15677 7 5 2 69349 78806
0 15678 7 1 2 80804 92244
0 15679 5 1 1 15678
0 15680 7 1 2 15676 15679
0 15681 5 1 1 15680
0 15682 7 1 2 92228 15681
0 15683 5 1 1 15682
0 15684 7 2 2 68813 81666
0 15685 7 1 2 90171 92245
0 15686 7 1 2 92249 15685
0 15687 5 1 1 15686
0 15688 7 1 2 15683 15687
0 15689 5 1 1 15688
0 15690 7 1 2 67218 15689
0 15691 5 1 1 15690
0 15692 7 2 2 88620 92246
0 15693 5 1 1 92251
0 15694 7 1 2 85707 90172
0 15695 7 1 2 92252 15694
0 15696 5 1 1 15695
0 15697 7 1 2 15691 15696
0 15698 5 1 1 15697
0 15699 7 1 2 70299 15698
0 15700 5 1 1 15699
0 15701 7 1 2 70894 91751
0 15702 7 1 2 92031 15701
0 15703 5 1 1 15702
0 15704 7 1 2 15700 15703
0 15705 5 1 1 15704
0 15706 7 1 2 65708 15705
0 15707 5 1 1 15706
0 15708 7 1 2 90178 86665
0 15709 5 1 1 15708
0 15710 7 2 2 63763 74620
0 15711 7 1 2 85322 92253
0 15712 5 1 1 15711
0 15713 7 1 2 15709 15712
0 15714 5 1 1 15713
0 15715 7 1 2 82845 15714
0 15716 5 1 1 15715
0 15717 7 3 2 69350 77813
0 15718 7 1 2 73986 84286
0 15719 7 1 2 92255 15718
0 15720 5 1 1 15719
0 15721 7 1 2 15716 15720
0 15722 5 1 1 15721
0 15723 7 1 2 69542 15722
0 15724 5 1 1 15723
0 15725 7 2 2 61826 87644
0 15726 7 1 2 90311 92258
0 15727 7 1 2 80451 15726
0 15728 5 1 1 15727
0 15729 7 1 2 15724 15728
0 15730 5 1 1 15729
0 15731 7 1 2 79902 15730
0 15732 5 1 1 15731
0 15733 7 6 2 68142 76666
0 15734 5 1 1 92260
0 15735 7 2 2 87319 92261
0 15736 5 2 1 92266
0 15737 7 1 2 70895 82320
0 15738 7 1 2 4020 1833
0 15739 5 1 1 15738
0 15740 7 1 2 83072 15739
0 15741 7 1 2 15737 15740
0 15742 5 1 1 15741
0 15743 7 1 2 92268 15742
0 15744 5 1 1 15743
0 15745 7 1 2 76801 15744
0 15746 5 1 1 15745
0 15747 7 3 2 80089 87691
0 15748 7 1 2 73847 92071
0 15749 7 1 2 92270 15748
0 15750 5 1 1 15749
0 15751 7 1 2 15746 15750
0 15752 5 1 1 15751
0 15753 7 1 2 73415 15752
0 15754 5 1 1 15753
0 15755 7 1 2 15732 15754
0 15756 7 1 2 15707 15755
0 15757 5 1 1 15756
0 15758 7 1 2 67659 15757
0 15759 5 1 1 15758
0 15760 7 3 2 69543 76695
0 15761 7 1 2 78504 84434
0 15762 7 1 2 91525 15761
0 15763 7 1 2 92273 15762
0 15764 5 1 1 15763
0 15765 7 1 2 68371 15764
0 15766 7 1 2 15759 15765
0 15767 7 1 2 15674 15766
0 15768 5 1 1 15767
0 15769 7 2 2 80000 84090
0 15770 5 1 1 92276
0 15771 7 5 2 64490 81245
0 15772 7 1 2 78693 92278
0 15773 5 1 1 15772
0 15774 7 1 2 15770 15773
0 15775 5 1 1 15774
0 15776 7 1 2 81162 15775
0 15777 5 1 1 15776
0 15778 7 1 2 83808 88298
0 15779 7 1 2 85603 15778
0 15780 5 1 1 15779
0 15781 7 1 2 15777 15780
0 15782 5 1 1 15781
0 15783 7 1 2 62380 15782
0 15784 5 1 1 15783
0 15785 7 1 2 72942 92277
0 15786 5 1 1 15785
0 15787 7 1 2 62809 81488
0 15788 7 1 2 91402 15787
0 15789 5 1 1 15788
0 15790 7 1 2 15786 15789
0 15791 5 1 1 15790
0 15792 7 1 2 70896 15791
0 15793 5 1 1 15792
0 15794 7 1 2 15784 15793
0 15795 5 1 1 15794
0 15796 7 1 2 81443 15795
0 15797 5 1 1 15796
0 15798 7 4 2 67984 72996
0 15799 7 5 2 69351 70897
0 15800 7 1 2 88574 92287
0 15801 7 1 2 80001 15800
0 15802 7 1 2 92283 15801
0 15803 5 1 1 15802
0 15804 7 1 2 15797 15803
0 15805 5 1 1 15804
0 15806 7 1 2 66436 15805
0 15807 5 1 1 15806
0 15808 7 1 2 72950 11295
0 15809 5 3 1 15808
0 15810 7 2 2 78807 78505
0 15811 7 2 2 78694 87090
0 15812 7 2 2 64491 92297
0 15813 7 1 2 92295 92299
0 15814 7 1 2 92292 15813
0 15815 5 1 1 15814
0 15816 7 1 2 15807 15815
0 15817 5 1 1 15816
0 15818 7 1 2 70300 15817
0 15819 5 1 1 15818
0 15820 7 1 2 81444 73063
0 15821 5 1 1 15820
0 15822 7 1 2 83103 77749
0 15823 5 1 1 15822
0 15824 7 1 2 15821 15823
0 15825 5 1 1 15824
0 15826 7 2 2 83809 75073
0 15827 7 1 2 78808 90002
0 15828 7 1 2 92301 15827
0 15829 7 1 2 15825 15828
0 15830 5 1 1 15829
0 15831 7 1 2 63525 15830
0 15832 7 1 2 15819 15831
0 15833 5 1 1 15832
0 15834 7 1 2 64098 15833
0 15835 7 1 2 15768 15834
0 15836 5 1 1 15835
0 15837 7 3 2 66687 78752
0 15838 7 2 2 86868 92303
0 15839 7 1 2 76220 92306
0 15840 5 1 1 15839
0 15841 7 3 2 65709 85916
0 15842 7 1 2 68814 91668
0 15843 7 1 2 92308 15842
0 15844 5 1 1 15843
0 15845 7 1 2 15840 15844
0 15846 5 1 1 15845
0 15847 7 1 2 61528 15846
0 15848 5 1 1 15847
0 15849 7 2 2 68815 82434
0 15850 7 1 2 67418 80225
0 15851 7 1 2 90913 15850
0 15852 7 1 2 92311 15851
0 15853 5 1 1 15852
0 15854 7 1 2 15848 15853
0 15855 5 1 1 15854
0 15856 7 1 2 88116 15855
0 15857 5 1 1 15856
0 15858 7 1 2 77362 4865
0 15859 5 1 1 15858
0 15860 7 1 2 79734 84047
0 15861 7 1 2 85650 15860
0 15862 7 1 2 15859 15861
0 15863 5 1 1 15862
0 15864 7 1 2 15857 15863
0 15865 5 1 1 15864
0 15866 7 1 2 68607 15865
0 15867 5 1 1 15866
0 15868 7 1 2 88094 90859
0 15869 7 2 2 89854 15868
0 15870 7 1 2 66437 77168
0 15871 7 1 2 77599 15870
0 15872 7 1 2 92313 15871
0 15873 5 1 1 15872
0 15874 7 1 2 15867 15873
0 15875 5 1 1 15874
0 15876 7 1 2 67219 15875
0 15877 5 1 1 15876
0 15878 7 1 2 63526 75320
0 15879 7 1 2 87277 15878
0 15880 7 1 2 92314 15879
0 15881 5 1 1 15880
0 15882 7 1 2 70013 15881
0 15883 7 1 2 15877 15882
0 15884 7 1 2 15836 15883
0 15885 5 1 1 15884
0 15886 7 1 2 70301 77814
0 15887 5 1 1 15886
0 15888 7 1 2 62810 90132
0 15889 5 1 1 15888
0 15890 7 1 2 15887 15889
0 15891 5 1 1 15890
0 15892 7 1 2 81082 15891
0 15893 5 1 1 15892
0 15894 7 2 2 86304 72446
0 15895 7 1 2 89556 92315
0 15896 5 1 1 15895
0 15897 7 1 2 15893 15896
0 15898 5 1 1 15897
0 15899 7 1 2 68608 15898
0 15900 5 1 1 15899
0 15901 7 2 2 80931 81515
0 15902 7 1 2 68816 92316
0 15903 7 1 2 92317 15902
0 15904 5 1 1 15903
0 15905 7 1 2 15900 15904
0 15906 5 1 1 15905
0 15907 7 1 2 63527 15906
0 15908 5 1 1 15907
0 15909 7 5 2 68964 73416
0 15910 5 1 1 92319
0 15911 7 3 2 76748 15910
0 15912 7 5 2 71308 92324
0 15913 5 1 1 92327
0 15914 7 2 2 73848 92328
0 15915 5 1 1 92332
0 15916 7 1 2 82321 74031
0 15917 7 1 2 92333 15916
0 15918 5 1 1 15917
0 15919 7 1 2 15908 15918
0 15920 5 1 1 15919
0 15921 7 1 2 67220 15920
0 15922 5 1 1 15921
0 15923 7 1 2 68609 15915
0 15924 5 1 1 15923
0 15925 7 2 2 71674 77356
0 15926 5 1 1 92334
0 15927 7 1 2 64099 92335
0 15928 5 2 1 15927
0 15929 7 1 2 63764 92336
0 15930 5 1 1 15929
0 15931 7 1 2 76397 15930
0 15932 7 1 2 15924 15931
0 15933 5 1 1 15932
0 15934 7 5 2 71216 71111
0 15935 5 1 1 92338
0 15936 7 1 2 70302 85783
0 15937 7 1 2 92339 15936
0 15938 5 1 1 15937
0 15939 7 1 2 15933 15938
0 15940 5 1 1 15939
0 15941 7 1 2 82322 15940
0 15942 5 1 1 15941
0 15943 7 1 2 15922 15942
0 15944 5 1 1 15943
0 15945 7 1 2 64688 15944
0 15946 5 1 1 15945
0 15947 7 1 2 88394 84512
0 15948 7 8 2 62545 73545
0 15949 5 1 1 92343
0 15950 7 2 2 80030 89259
0 15951 7 1 2 92344 92351
0 15952 7 1 2 15947 15951
0 15953 5 1 1 15952
0 15954 7 1 2 15946 15953
0 15955 5 1 1 15954
0 15956 7 1 2 63296 15955
0 15957 5 1 1 15956
0 15958 7 2 2 65966 75220
0 15959 7 1 2 82868 92353
0 15960 5 1 1 15959
0 15961 7 1 2 91504 15960
0 15962 5 1 1 15961
0 15963 7 1 2 61529 15962
0 15964 5 1 1 15963
0 15965 7 8 2 66438 80185
0 15966 5 1 1 92355
0 15967 7 1 2 85736 90584
0 15968 7 1 2 92356 15967
0 15969 5 1 1 15968
0 15970 7 1 2 15964 15969
0 15971 5 1 1 15970
0 15972 7 1 2 83810 15971
0 15973 5 1 1 15972
0 15974 7 1 2 80462 84189
0 15975 5 1 1 15974
0 15976 7 1 2 80147 82919
0 15977 5 1 1 15976
0 15978 7 1 2 15975 15977
0 15979 5 1 1 15978
0 15980 7 1 2 67221 15979
0 15981 5 1 1 15980
0 15982 7 2 2 67660 74678
0 15983 5 1 1 92363
0 15984 7 1 2 71505 15983
0 15985 5 1 1 15984
0 15986 7 1 2 82542 86039
0 15987 7 1 2 15985 15986
0 15988 5 1 1 15987
0 15989 7 1 2 15981 15988
0 15990 5 1 1 15989
0 15991 7 1 2 82323 15990
0 15992 5 1 1 15991
0 15993 7 1 2 15973 15992
0 15994 5 1 1 15993
0 15995 7 1 2 67419 15994
0 15996 5 1 1 15995
0 15997 7 1 2 77725 11760
0 15998 5 1 1 15997
0 15999 7 2 2 80971 86305
0 16000 7 1 2 71930 84566
0 16001 7 1 2 92365 16000
0 16002 7 1 2 15998 16001
0 16003 5 1 1 16002
0 16004 7 1 2 81083 74839
0 16005 7 1 2 85753 16004
0 16006 5 1 1 16005
0 16007 7 1 2 16003 16006
0 16008 5 1 1 16007
0 16009 7 1 2 64689 16008
0 16010 5 1 1 16009
0 16011 7 1 2 62381 85750
0 16012 5 2 1 16011
0 16013 7 1 2 79356 76077
0 16014 7 1 2 80472 16013
0 16015 7 1 2 92367 16014
0 16016 5 1 1 16015
0 16017 7 1 2 16010 16016
0 16018 5 1 1 16017
0 16019 7 1 2 81627 16018
0 16020 5 1 1 16019
0 16021 7 1 2 15996 16020
0 16022 5 1 1 16021
0 16023 7 1 2 65710 16022
0 16024 5 1 1 16023
0 16025 7 1 2 79222 91897
0 16026 5 1 1 16025
0 16027 7 4 2 68817 73160
0 16028 7 4 2 74178 92369
0 16029 5 2 1 92373
0 16030 7 1 2 71931 92374
0 16031 5 2 1 16030
0 16032 7 1 2 14522 92379
0 16033 5 1 1 16032
0 16034 7 1 2 82324 16033
0 16035 5 1 1 16034
0 16036 7 1 2 16026 16035
0 16037 5 1 1 16036
0 16038 7 1 2 64100 16037
0 16039 5 1 1 16038
0 16040 7 3 2 65967 79903
0 16041 7 1 2 81084 75221
0 16042 7 1 2 92381 16041
0 16043 5 1 1 16042
0 16044 7 1 2 16039 16043
0 16045 5 1 1 16044
0 16046 7 1 2 64690 16045
0 16047 5 1 1 16046
0 16048 7 2 2 76078 80186
0 16049 7 1 2 73417 92384
0 16050 7 1 2 82301 16049
0 16051 5 1 1 16050
0 16052 7 1 2 16047 16051
0 16053 5 1 1 16052
0 16054 7 1 2 81628 16053
0 16055 5 1 1 16054
0 16056 7 1 2 16024 16055
0 16057 5 1 1 16056
0 16058 7 1 2 65382 16057
0 16059 5 1 1 16058
0 16060 7 1 2 15957 16059
0 16061 5 1 1 16060
0 16062 7 1 2 61827 16061
0 16063 5 1 1 16062
0 16064 7 1 2 822 14610
0 16065 5 1 1 16064
0 16066 7 1 2 63528 16065
0 16067 5 1 1 16066
0 16068 7 1 2 88490 84753
0 16069 5 1 1 16068
0 16070 7 1 2 16067 16069
0 16071 5 1 1 16070
0 16072 7 1 2 70303 92267
0 16073 7 1 2 16071 16072
0 16074 5 1 1 16073
0 16075 7 1 2 65119 16074
0 16076 7 1 2 16063 16075
0 16077 5 1 1 16076
0 16078 7 1 2 15885 16077
0 16079 5 1 1 16078
0 16080 7 3 2 81557 79437
0 16081 7 1 2 76885 88007
0 16082 5 1 1 16081
0 16083 7 1 2 84830 16082
0 16084 5 1 1 16083
0 16085 7 1 2 72997 16084
0 16086 5 1 1 16085
0 16087 7 2 2 71112 91421
0 16088 7 2 2 71217 78190
0 16089 7 1 2 92389 92391
0 16090 5 1 1 16089
0 16091 7 1 2 16086 16090
0 16092 5 1 1 16091
0 16093 7 1 2 85502 16092
0 16094 5 1 1 16093
0 16095 7 2 2 76293 76696
0 16096 7 1 2 67661 91988
0 16097 7 1 2 92393 16096
0 16098 5 1 1 16097
0 16099 7 1 2 16094 16098
0 16100 5 1 1 16099
0 16101 7 1 2 92386 16100
0 16102 5 1 1 16101
0 16103 7 9 2 63933 70898
0 16104 5 2 1 92395
0 16105 7 2 2 62546 92396
0 16106 5 3 1 92406
0 16107 7 2 2 65383 92408
0 16108 7 1 2 73546 85870
0 16109 5 1 1 16108
0 16110 7 1 2 77770 16109
0 16111 5 1 1 16110
0 16112 7 1 2 92411 16111
0 16113 5 1 1 16112
0 16114 7 2 2 71218 72409
0 16115 5 1 1 92413
0 16116 7 1 2 86396 16115
0 16117 5 1 1 16116
0 16118 7 1 2 65711 16117
0 16119 5 1 1 16118
0 16120 7 1 2 83191 92377
0 16121 5 1 1 16120
0 16122 7 1 2 67222 16121
0 16123 5 1 1 16122
0 16124 7 1 2 16119 16123
0 16125 7 1 2 16113 16124
0 16126 5 1 1 16125
0 16127 7 1 2 70014 16126
0 16128 5 1 1 16127
0 16129 7 1 2 79885 79554
0 16130 5 1 1 16129
0 16131 7 1 2 16128 16130
0 16132 5 1 1 16131
0 16133 7 1 2 64101 16132
0 16134 5 1 1 16133
0 16135 7 1 2 74208 79590
0 16136 5 1 1 16135
0 16137 7 1 2 68372 16136
0 16138 7 1 2 16134 16137
0 16139 5 1 1 16138
0 16140 7 6 2 65384 85052
0 16141 7 1 2 79476 92415
0 16142 5 1 1 16141
0 16143 7 1 2 76958 16142
0 16144 5 1 1 16143
0 16145 7 1 2 62382 79509
0 16146 5 2 1 16145
0 16147 7 1 2 84985 92421
0 16148 7 1 2 16144 16147
0 16149 5 1 1 16148
0 16150 7 1 2 63529 16149
0 16151 5 1 1 16150
0 16152 7 1 2 68610 16151
0 16153 7 1 2 16139 16152
0 16154 5 1 1 16153
0 16155 7 1 2 71113 85428
0 16156 5 2 1 16155
0 16157 7 3 2 71309 74179
0 16158 5 1 1 92425
0 16159 7 1 2 72821 16158
0 16160 5 1 1 16159
0 16161 7 1 2 71219 74192
0 16162 5 2 1 16161
0 16163 7 1 2 76938 92428
0 16164 7 1 2 16160 16163
0 16165 5 1 1 16164
0 16166 7 1 2 92423 16165
0 16167 5 1 1 16166
0 16168 7 1 2 63765 16167
0 16169 5 1 1 16168
0 16170 7 1 2 64102 91059
0 16171 7 1 2 91082 16170
0 16172 5 1 1 16171
0 16173 7 1 2 16169 16172
0 16174 5 1 1 16173
0 16175 7 1 2 68373 16174
0 16176 5 1 1 16175
0 16177 7 1 2 84850 76380
0 16178 5 1 1 16177
0 16179 7 1 2 16176 16178
0 16180 5 1 1 16179
0 16181 7 1 2 67223 16180
0 16182 5 1 1 16181
0 16183 7 1 2 91066 76866
0 16184 7 1 2 74048 16183
0 16185 5 1 1 16184
0 16186 7 1 2 82371 16185
0 16187 7 1 2 16182 16186
0 16188 7 1 2 16154 16187
0 16189 5 1 1 16188
0 16190 7 4 2 71310 72041
0 16191 5 5 1 92430
0 16192 7 2 2 75742 92434
0 16193 5 3 1 92439
0 16194 7 1 2 74590 92441
0 16195 5 1 1 16194
0 16196 7 4 2 83739 85036
0 16197 7 1 2 70661 73896
0 16198 7 1 2 92444 16197
0 16199 5 1 1 16198
0 16200 7 1 2 16195 16199
0 16201 5 1 1 16200
0 16202 7 1 2 62811 16201
0 16203 5 1 1 16202
0 16204 7 2 2 63766 73959
0 16205 7 1 2 77765 72384
0 16206 7 1 2 92448 16205
0 16207 5 1 1 16206
0 16208 7 1 2 16203 16207
0 16209 5 1 1 16208
0 16210 7 1 2 78067 16209
0 16211 5 1 1 16210
0 16212 7 1 2 82386 16211
0 16213 5 1 1 16212
0 16214 7 1 2 79357 82752
0 16215 7 1 2 16213 16214
0 16216 7 1 2 16189 16215
0 16217 5 1 1 16216
0 16218 7 1 2 16102 16217
0 16219 5 1 1 16218
0 16220 7 1 2 76138 16219
0 16221 5 1 1 16220
0 16222 7 1 2 69775 16221
0 16223 7 1 2 16079 16222
0 16224 5 1 1 16223
0 16225 7 3 2 66091 90700
0 16226 5 1 1 92450
0 16227 7 9 2 91366 91856
0 16228 5 1 1 92453
0 16229 7 1 2 16226 16228
0 16230 5 35 1 16229
0 16231 7 1 2 62383 84986
0 16232 7 1 2 91907 91982
0 16233 7 1 2 16231 16232
0 16234 5 1 1 16233
0 16235 7 1 2 81760 89225
0 16236 5 1 1 16235
0 16237 7 1 2 81731 88834
0 16238 5 1 1 16237
0 16239 7 1 2 16236 16238
0 16240 5 1 1 16239
0 16241 7 1 2 66439 16240
0 16242 5 1 1 16241
0 16243 7 3 2 61530 81812
0 16244 7 1 2 89226 92497
0 16245 5 1 1 16244
0 16246 7 1 2 16242 16245
0 16247 5 1 1 16246
0 16248 7 1 2 75719 91899
0 16249 7 1 2 16247 16248
0 16250 5 1 1 16249
0 16251 7 1 2 16234 16250
0 16252 5 1 1 16251
0 16253 7 1 2 70304 16252
0 16254 5 1 1 16253
0 16255 7 1 2 81813 79577
0 16256 7 1 2 91511 16255
0 16257 7 1 2 86187 92426
0 16258 7 1 2 16256 16257
0 16259 5 1 1 16258
0 16260 7 1 2 16254 16259
0 16261 5 1 1 16260
0 16262 7 1 2 64691 16261
0 16263 5 1 1 16262
0 16264 7 4 2 84619 77883
0 16265 7 1 2 70662 92500
0 16266 5 1 1 16265
0 16267 7 1 2 88498 16266
0 16268 5 1 1 16267
0 16269 7 1 2 73547 88788
0 16270 7 1 2 16268 16269
0 16271 5 1 1 16270
0 16272 7 2 2 88531 79927
0 16273 7 1 2 67662 81761
0 16274 7 1 2 92504 16273
0 16275 5 1 1 16274
0 16276 7 1 2 16271 16275
0 16277 5 1 1 16276
0 16278 7 1 2 70305 16277
0 16279 5 1 1 16278
0 16280 7 1 2 86197 90787
0 16281 5 1 1 16280
0 16282 7 1 2 73944 91560
0 16283 5 2 1 16282
0 16284 7 1 2 92380 92506
0 16285 5 1 1 16284
0 16286 7 1 2 83437 16285
0 16287 5 1 1 16286
0 16288 7 1 2 16281 16287
0 16289 5 1 1 16288
0 16290 7 1 2 65385 16289
0 16291 5 1 1 16290
0 16292 7 1 2 81762 86188
0 16293 5 1 1 16292
0 16294 7 1 2 90790 16293
0 16295 5 1 1 16294
0 16296 7 1 2 73310 16295
0 16297 5 1 1 16296
0 16298 7 1 2 81763 84162
0 16299 7 1 2 85968 16298
0 16300 5 1 1 16299
0 16301 7 1 2 16297 16300
0 16302 5 1 1 16301
0 16303 7 1 2 78428 16302
0 16304 5 1 1 16303
0 16305 7 1 2 16291 16304
0 16306 7 1 2 16279 16305
0 16307 5 1 1 16306
0 16308 7 1 2 79438 16307
0 16309 5 1 1 16308
0 16310 7 1 2 82928 92061
0 16311 5 1 1 16310
0 16312 7 2 2 73911 82435
0 16313 7 2 2 80201 82880
0 16314 7 1 2 92508 92510
0 16315 5 1 1 16314
0 16316 7 1 2 16311 16315
0 16317 5 1 1 16316
0 16318 7 1 2 84048 16317
0 16319 5 1 1 16318
0 16320 7 1 2 66440 16319
0 16321 7 1 2 16309 16320
0 16322 5 1 1 16321
0 16323 7 1 2 91677 91752
0 16324 5 1 1 16323
0 16325 7 1 2 91502 16324
0 16326 5 1 1 16325
0 16327 7 1 2 71311 16326
0 16328 5 1 1 16327
0 16329 7 1 2 72943 91757
0 16330 5 1 1 16329
0 16331 7 5 2 65386 71932
0 16332 5 2 1 92512
0 16333 7 1 2 89415 92513
0 16334 5 1 1 16333
0 16335 7 1 2 16330 16334
0 16336 5 1 1 16335
0 16337 7 1 2 70663 16336
0 16338 5 1 1 16337
0 16339 7 1 2 16328 16338
0 16340 5 1 1 16339
0 16341 7 1 2 80202 16340
0 16342 5 1 1 16341
0 16343 7 3 2 70664 89777
0 16344 5 1 1 92519
0 16345 7 3 2 80821 83648
0 16346 7 1 2 82543 92522
0 16347 7 1 2 92520 16346
0 16348 5 1 1 16347
0 16349 7 1 2 16342 16348
0 16350 5 1 1 16349
0 16351 7 1 2 70899 16350
0 16352 5 1 1 16351
0 16353 7 1 2 78753 76697
0 16354 7 1 2 87980 16353
0 16355 7 1 2 92387 16354
0 16356 5 1 1 16355
0 16357 7 1 2 61531 16356
0 16358 7 1 2 16352 16357
0 16359 5 1 1 16358
0 16360 7 1 2 70015 16359
0 16361 7 1 2 16322 16360
0 16362 5 1 1 16361
0 16363 7 2 2 91053 92501
0 16364 7 1 2 80203 92525
0 16365 5 1 1 16364
0 16366 7 1 2 88491 81489
0 16367 5 1 1 16366
0 16368 7 1 2 16365 16367
0 16369 5 1 1 16368
0 16370 7 1 2 61532 16369
0 16371 5 1 1 16370
0 16372 7 2 2 63123 87402
0 16373 7 1 2 92526 92527
0 16374 5 1 1 16373
0 16375 7 1 2 16371 16374
0 16376 5 1 1 16375
0 16377 7 1 2 70306 16376
0 16378 5 1 1 16377
0 16379 7 1 2 77797 88134
0 16380 7 1 2 79211 16379
0 16381 5 1 1 16380
0 16382 7 1 2 16378 16381
0 16383 5 1 1 16382
0 16384 7 1 2 77330 81558
0 16385 7 1 2 16383 16384
0 16386 5 1 1 16385
0 16387 7 1 2 16362 16386
0 16388 5 1 1 16387
0 16389 7 1 2 64103 16388
0 16390 5 1 1 16389
0 16391 7 1 2 16263 16390
0 16392 5 1 1 16391
0 16393 7 1 2 61828 16392
0 16394 5 1 1 16393
0 16395 7 1 2 76139 82567
0 16396 5 1 1 16395
0 16397 7 4 2 66441 78918
0 16398 7 1 2 87578 92529
0 16399 5 1 1 16398
0 16400 7 4 2 68374 79750
0 16401 7 1 2 91268 92533
0 16402 5 1 1 16401
0 16403 7 1 2 16399 16402
0 16404 7 1 2 16396 16403
0 16405 5 1 1 16404
0 16406 7 1 2 84227 16405
0 16407 5 1 1 16406
0 16408 7 6 2 63124 70016
0 16409 7 1 2 81629 92537
0 16410 7 1 2 87320 16409
0 16411 5 1 1 16410
0 16412 7 1 2 16407 16411
0 16413 5 1 1 16412
0 16414 7 1 2 82155 85467
0 16415 7 1 2 16413 16414
0 16416 5 1 1 16415
0 16417 7 1 2 64914 16416
0 16418 7 1 2 16394 16417
0 16419 5 1 1 16418
0 16420 7 1 2 92462 16419
0 16421 7 1 2 16224 16420
0 16422 5 1 1 16421
0 16423 7 1 2 83009 84538
0 16424 7 20 2 62998 67985
0 16425 5 1 1 92543
0 16426 7 2 2 90985 92544
0 16427 7 1 2 87458 91802
0 16428 7 1 2 92563 16427
0 16429 7 2 2 16423 16428
0 16430 5 1 1 92565
0 16431 7 1 2 65712 92566
0 16432 5 1 1 16431
0 16433 7 2 2 67420 91835
0 16434 7 1 2 91013 84540
0 16435 7 1 2 92567 16434
0 16436 5 1 1 16435
0 16437 7 1 2 16432 16436
0 16438 7 1 2 16422 16437
0 16439 5 1 1 16438
0 16440 7 1 2 64324 16439
0 16441 5 1 1 16440
0 16442 7 1 2 80726 83253
0 16443 5 1 1 16442
0 16444 7 6 2 67421 69544
0 16445 5 1 1 92569
0 16446 7 1 2 77269 16445
0 16447 5 1 1 16446
0 16448 7 1 2 88897 16447
0 16449 7 1 2 88386 16448
0 16450 5 1 1 16449
0 16451 7 1 2 16443 16450
0 16452 5 1 1 16451
0 16453 7 1 2 63934 16452
0 16454 5 1 1 16453
0 16455 7 2 2 63125 82985
0 16456 7 1 2 92144 92575
0 16457 5 1 1 16456
0 16458 7 1 2 16454 16457
0 16459 5 3 1 16458
0 16460 7 1 2 90585 92577
0 16461 5 1 1 16460
0 16462 7 1 2 88696 82306
0 16463 7 1 2 89540 16462
0 16464 5 1 1 16463
0 16465 7 1 2 16461 16464
0 16466 5 1 1 16465
0 16467 7 1 2 64104 16466
0 16468 5 1 1 16467
0 16469 7 4 2 68818 82804
0 16470 7 1 2 85708 83454
0 16471 7 1 2 88697 16470
0 16472 7 1 2 92580 16471
0 16473 5 1 1 16472
0 16474 7 1 2 16468 16473
0 16475 5 1 1 16474
0 16476 7 1 2 67224 16475
0 16477 5 1 1 16476
0 16478 7 1 2 88285 91584
0 16479 7 1 2 92578 16478
0 16480 5 1 1 16479
0 16481 7 1 2 16477 16480
0 16482 5 1 1 16481
0 16483 7 1 2 66688 16482
0 16484 5 1 1 16483
0 16485 7 1 2 75380 88266
0 16486 7 1 2 92579 16485
0 16487 5 1 1 16486
0 16488 7 1 2 16484 16487
0 16489 5 1 1 16488
0 16490 7 1 2 70900 16489
0 16491 5 1 1 16490
0 16492 7 1 2 89061 1987
0 16493 5 1 1 16492
0 16494 7 1 2 61533 16493
0 16495 5 1 1 16494
0 16496 7 1 2 81911 80331
0 16497 5 1 1 16496
0 16498 7 1 2 16495 16497
0 16499 5 1 1 16498
0 16500 7 2 2 83104 90886
0 16501 5 1 1 92584
0 16502 7 1 2 16499 92585
0 16503 5 1 1 16502
0 16504 7 3 2 67422 72320
0 16505 7 1 2 69545 92586
0 16506 7 3 2 63126 87645
0 16507 7 2 2 76555 77766
0 16508 7 1 2 92589 92592
0 16509 7 1 2 16505 16508
0 16510 5 1 1 16509
0 16511 7 1 2 16503 16510
0 16512 5 1 1 16511
0 16513 7 1 2 83649 16512
0 16514 5 1 1 16513
0 16515 7 1 2 16491 16514
0 16516 5 1 1 16515
0 16517 7 1 2 69776 16516
0 16518 5 1 1 16517
0 16519 7 1 2 83952 86739
0 16520 5 2 1 16519
0 16521 7 2 2 66442 79237
0 16522 7 1 2 92247 92596
0 16523 5 1 1 16522
0 16524 7 1 2 92594 16523
0 16525 5 1 1 16524
0 16526 7 1 2 62812 16525
0 16527 5 1 1 16526
0 16528 7 5 2 64692 86306
0 16529 7 1 2 90081 92598
0 16530 5 1 1 16529
0 16531 7 1 2 16527 16530
0 16532 5 1 1 16531
0 16533 7 1 2 63935 16532
0 16534 5 1 1 16533
0 16535 7 2 2 72780 80068
0 16536 7 1 2 87321 92603
0 16537 5 2 1 16536
0 16538 7 1 2 16534 92605
0 16539 5 1 1 16538
0 16540 7 1 2 92284 16539
0 16541 5 1 1 16540
0 16542 7 2 2 63127 88244
0 16543 5 1 1 92607
0 16544 7 1 2 71819 80784
0 16545 7 1 2 91784 16544
0 16546 7 1 2 92608 16545
0 16547 5 1 1 16546
0 16548 7 1 2 16541 16547
0 16549 5 1 1 16548
0 16550 7 1 2 88994 16549
0 16551 5 1 1 16550
0 16552 7 1 2 16518 16551
0 16553 5 1 1 16552
0 16554 7 1 2 70665 16553
0 16555 5 1 1 16554
0 16556 7 2 2 63530 72042
0 16557 7 1 2 66689 85121
0 16558 7 2 2 73884 16557
0 16559 5 1 1 92611
0 16560 7 1 2 16501 16559
0 16561 5 1 1 16560
0 16562 7 1 2 74237 16561
0 16563 5 1 1 16562
0 16564 7 5 2 64915 73255
0 16565 7 1 2 67423 85319
0 16566 7 1 2 92613 16565
0 16567 5 1 1 16566
0 16568 7 1 2 16563 16567
0 16569 5 1 1 16568
0 16570 7 1 2 81085 16569
0 16571 5 1 1 16570
0 16572 7 3 2 72998 83105
0 16573 7 1 2 82394 90860
0 16574 7 1 2 91491 16573
0 16575 7 1 2 92618 16574
0 16576 5 1 1 16575
0 16577 7 1 2 16571 16576
0 16578 5 1 1 16577
0 16579 7 1 2 64693 16578
0 16580 5 1 1 16579
0 16581 7 1 2 71776 80822
0 16582 7 1 2 71522 92019
0 16583 7 1 2 16581 16582
0 16584 5 1 1 16583
0 16585 7 1 2 84473 75062
0 16586 7 1 2 74142 16585
0 16587 5 1 1 16586
0 16588 7 1 2 16584 16587
0 16589 5 1 1 16588
0 16590 7 1 2 88906 16589
0 16591 5 1 1 16590
0 16592 7 1 2 16580 16591
0 16593 5 1 1 16592
0 16594 7 1 2 92609 16593
0 16595 5 1 1 16594
0 16596 7 1 2 16555 16595
0 16597 5 1 1 16596
0 16598 7 1 2 70017 16597
0 16599 5 1 1 16598
0 16600 7 2 2 62547 91466
0 16601 5 1 1 92621
0 16602 7 1 2 67424 90259
0 16603 5 2 1 16602
0 16604 7 1 2 83974 92623
0 16605 5 2 1 16604
0 16606 7 1 2 73548 85451
0 16607 7 1 2 92625 16606
0 16608 5 1 1 16607
0 16609 7 1 2 16601 16608
0 16610 5 1 1 16609
0 16611 7 1 2 64105 16610
0 16612 5 1 1 16611
0 16613 7 1 2 92145 92279
0 16614 5 1 1 16613
0 16615 7 1 2 16612 16614
0 16616 5 1 1 16615
0 16617 7 1 2 63936 16616
0 16618 5 1 1 16617
0 16619 7 1 2 87322 88065
0 16620 5 3 1 16619
0 16621 7 1 2 16618 92627
0 16622 5 1 1 16621
0 16623 7 1 2 81984 89208
0 16624 7 1 2 92285 16623
0 16625 7 1 2 16622 16624
0 16626 5 1 1 16625
0 16627 7 1 2 16599 16626
0 16628 5 1 1 16627
0 16629 7 7 2 69173 90652
0 16630 7 22 2 66092 67769
0 16631 5 3 1 92637
0 16632 7 3 2 70307 92638
0 16633 7 1 2 92630 92662
0 16634 7 1 2 16628 16633
0 16635 5 1 1 16634
0 16636 7 1 2 16441 16635
0 16637 7 1 2 15619 16636
0 16638 5 1 1 16637
0 16639 7 1 2 66922 16638
0 16640 5 1 1 16639
0 16641 7 14 2 64325 92463
0 16642 7 2 2 90104 82908
0 16643 7 2 2 80972 75831
0 16644 7 1 2 92679 92681
0 16645 5 1 1 16644
0 16646 7 4 2 70018 75411
0 16647 7 1 2 82168 92683
0 16648 5 1 1 16647
0 16649 7 1 2 78411 89956
0 16650 5 1 1 16649
0 16651 7 1 2 16648 16650
0 16652 5 1 1 16651
0 16653 7 3 2 82846 91451
0 16654 5 1 1 92687
0 16655 7 1 2 74268 92688
0 16656 7 1 2 16652 16655
0 16657 5 1 1 16656
0 16658 7 1 2 16645 16657
0 16659 5 1 1 16658
0 16660 7 1 2 63297 16659
0 16661 5 1 1 16660
0 16662 7 2 2 67986 81580
0 16663 7 1 2 90053 92690
0 16664 7 1 2 92680 16663
0 16665 5 1 1 16664
0 16666 7 1 2 16661 16665
0 16667 5 1 1 16666
0 16668 7 1 2 62384 16667
0 16669 5 1 1 16668
0 16670 7 3 2 68143 75764
0 16671 5 1 1 92692
0 16672 7 1 2 85110 16671
0 16673 5 23 1 16672
0 16674 7 2 2 69352 71725
0 16675 7 1 2 87597 83023
0 16676 7 1 2 92718 16675
0 16677 7 1 2 92695 16676
0 16678 5 1 1 16677
0 16679 7 1 2 16669 16678
0 16680 5 1 1 16679
0 16681 7 1 2 64694 16680
0 16682 5 1 1 16681
0 16683 7 2 2 66923 91836
0 16684 7 2 2 80347 81246
0 16685 7 1 2 69353 76917
0 16686 7 1 2 92722 16685
0 16687 7 1 2 92720 16686
0 16688 5 1 1 16687
0 16689 7 1 2 16682 16688
0 16690 5 1 1 16689
0 16691 7 1 2 71312 16690
0 16692 5 1 1 16691
0 16693 7 5 2 86943 71051
0 16694 5 1 1 92724
0 16695 7 1 2 91669 92725
0 16696 7 1 2 85257 16695
0 16697 5 1 1 16696
0 16698 7 5 2 69777 82805
0 16699 7 1 2 85076 92729
0 16700 7 1 2 91837 16699
0 16701 5 1 1 16700
0 16702 7 1 2 16697 16701
0 16703 5 1 1 16702
0 16704 7 1 2 68611 16703
0 16705 5 1 1 16704
0 16706 7 1 2 67225 74966
0 16707 7 1 2 91577 16706
0 16708 7 1 2 88727 16707
0 16709 5 1 1 16708
0 16710 7 1 2 16705 16709
0 16711 5 1 1 16710
0 16712 7 1 2 70308 16711
0 16713 5 1 1 16712
0 16714 7 1 2 65387 74967
0 16715 7 1 2 88556 16714
0 16716 7 1 2 90942 92590
0 16717 7 1 2 16715 16716
0 16718 5 1 1 16717
0 16719 7 1 2 16713 16718
0 16720 5 1 1 16719
0 16721 7 1 2 66924 16720
0 16722 5 1 1 16721
0 16723 7 4 2 71777 89931
0 16724 7 1 2 71726 92734
0 16725 5 1 1 16724
0 16726 7 7 2 68612 76698
0 16727 7 1 2 61829 92738
0 16728 5 1 1 16727
0 16729 7 1 2 16725 16728
0 16730 5 1 1 16729
0 16731 7 2 2 61534 90474
0 16732 7 1 2 64492 92745
0 16733 7 1 2 89487 16732
0 16734 7 1 2 16730 16733
0 16735 5 1 1 16734
0 16736 7 1 2 16722 16735
0 16737 5 1 1 16736
0 16738 7 1 2 70019 16737
0 16739 5 1 1 16738
0 16740 7 2 2 85122 80412
0 16741 7 2 2 82911 92747
0 16742 7 1 2 73064 82075
0 16743 7 1 2 88409 16742
0 16744 7 1 2 92749 16743
0 16745 5 1 1 16744
0 16746 7 1 2 16739 16745
0 16747 5 1 1 16746
0 16748 7 1 2 70901 16747
0 16749 5 1 1 16748
0 16750 7 1 2 16692 16749
0 16751 5 1 1 16750
0 16752 7 1 2 92665 16751
0 16753 5 1 1 16752
0 16754 7 1 2 62057 81314
0 16755 5 1 1 16754
0 16756 7 1 2 84784 87617
0 16757 5 1 1 16756
0 16758 7 1 2 16755 16757
0 16759 5 2 1 16758
0 16760 7 2 2 74415 92751
0 16761 5 1 1 92753
0 16762 7 1 2 86603 90586
0 16763 7 1 2 86084 16762
0 16764 5 1 1 16763
0 16765 7 1 2 16761 16764
0 16766 5 1 1 16765
0 16767 7 1 2 75720 16766
0 16768 5 1 1 16767
0 16769 7 1 2 90887 92752
0 16770 5 1 1 16769
0 16771 7 3 2 65713 86604
0 16772 5 1 1 92755
0 16773 7 2 2 63767 83181
0 16774 7 1 2 91983 92758
0 16775 7 1 2 92756 16774
0 16776 5 1 1 16775
0 16777 7 1 2 16770 16776
0 16778 5 1 1 16777
0 16779 7 1 2 70309 16778
0 16780 5 1 1 16779
0 16781 7 1 2 16768 16780
0 16782 5 1 1 16781
0 16783 7 1 2 90566 16782
0 16784 5 1 1 16783
0 16785 7 3 2 62548 81912
0 16786 5 1 1 92760
0 16787 7 1 2 73203 92761
0 16788 7 1 2 92754 16787
0 16789 5 1 1 16788
0 16790 7 1 2 16784 16789
0 16791 5 1 1 16790
0 16792 7 61 2 69174 64493
0 16793 7 5 2 61830 67770
0 16794 7 2 2 92763 92824
0 16795 7 15 2 66093 66209
0 16796 7 16 2 67841 63128
0 16797 5 1 1 92846
0 16798 7 1 2 92831 92847
0 16799 7 1 2 92829 16798
0 16800 7 1 2 16791 16799
0 16801 5 1 1 16800
0 16802 7 1 2 16753 16801
0 16803 5 1 1 16802
0 16804 7 1 2 74110 16803
0 16805 5 1 1 16804
0 16806 7 1 2 85992 91736
0 16807 5 1 1 16806
0 16808 7 5 2 65388 71572
0 16809 7 2 2 85549 92862
0 16810 5 3 1 92867
0 16811 7 4 2 77232 82372
0 16812 7 1 2 86260 92872
0 16813 7 1 2 92868 16812
0 16814 5 1 1 16813
0 16815 7 1 2 16807 16814
0 16816 5 1 1 16815
0 16817 7 1 2 65120 16816
0 16818 5 1 1 16817
0 16819 7 2 2 82525 90495
0 16820 7 1 2 87585 91578
0 16821 7 1 2 92876 16820
0 16822 5 1 1 16821
0 16823 7 1 2 16818 16822
0 16824 5 1 1 16823
0 16825 7 1 2 69778 16824
0 16826 5 1 1 16825
0 16827 7 2 2 82526 90764
0 16828 7 1 2 91854 92878
0 16829 5 1 1 16828
0 16830 7 3 2 64695 80002
0 16831 7 1 2 89133 92880
0 16832 5 1 1 16831
0 16833 7 1 2 16829 16832
0 16834 5 1 1 16833
0 16835 7 1 2 83677 91993
0 16836 7 1 2 16834 16835
0 16837 5 1 1 16836
0 16838 7 1 2 16826 16837
0 16839 5 1 1 16838
0 16840 7 1 2 63531 16839
0 16841 5 1 1 16840
0 16842 7 4 2 67425 68144
0 16843 7 2 2 67226 92883
0 16844 7 1 2 92879 92887
0 16845 5 1 1 16844
0 16846 7 2 2 85134 92881
0 16847 5 1 1 92889
0 16848 7 1 2 16845 16847
0 16849 5 1 1 16848
0 16850 7 4 2 63129 83286
0 16851 7 1 2 87603 92891
0 16852 7 1 2 16849 16851
0 16853 5 1 1 16852
0 16854 7 1 2 16841 16853
0 16855 5 1 1 16854
0 16856 7 1 2 64494 16855
0 16857 5 1 1 16856
0 16858 7 3 2 77127 75251
0 16859 7 1 2 68613 82806
0 16860 7 1 2 92895 16859
0 16861 7 1 2 92568 16860
0 16862 5 1 1 16861
0 16863 7 1 2 16857 16862
0 16864 5 2 1 16863
0 16865 7 1 2 66094 92898
0 16866 5 1 1 16865
0 16867 7 1 2 88777 91922
0 16868 7 1 2 81510 16867
0 16869 5 1 1 16868
0 16870 7 1 2 16866 16869
0 16871 5 1 1 16870
0 16872 7 1 2 90701 16871
0 16873 5 1 1 16872
0 16874 7 1 2 92454 92899
0 16875 5 1 1 16874
0 16876 7 1 2 16430 16875
0 16877 7 1 2 16873 16876
0 16878 5 1 1 16877
0 16879 7 1 2 67663 16878
0 16880 5 1 1 16879
0 16881 7 4 2 66443 90185
0 16882 5 1 1 92900
0 16883 7 1 2 11989 16882
0 16884 5 10 1 16883
0 16885 7 1 2 76802 92904
0 16886 5 1 1 16885
0 16887 7 1 2 85264 86760
0 16888 7 1 2 91289 16887
0 16889 5 1 1 16888
0 16890 7 1 2 16886 16889
0 16891 5 1 1 16890
0 16892 7 1 2 79122 16891
0 16893 5 1 1 16892
0 16894 7 2 2 81370 80294
0 16895 7 1 2 80973 89990
0 16896 7 1 2 92914 16895
0 16897 5 1 1 16896
0 16898 7 1 2 16893 16897
0 16899 5 1 1 16898
0 16900 7 2 2 70666 82937
0 16901 7 1 2 77470 92916
0 16902 7 1 2 92464 16901
0 16903 7 1 2 16899 16902
0 16904 5 1 1 16903
0 16905 7 1 2 16880 16904
0 16906 5 1 1 16905
0 16907 7 1 2 64326 16906
0 16908 5 1 1 16907
0 16909 7 6 2 66690 77233
0 16910 7 1 2 82561 92918
0 16911 5 1 1 16910
0 16912 7 1 2 76140 89377
0 16913 5 1 1 16912
0 16914 7 1 2 16911 16913
0 16915 5 1 1 16914
0 16916 7 1 2 64916 16915
0 16917 5 1 1 16916
0 16918 7 3 2 76079 81985
0 16919 5 1 1 92924
0 16920 7 1 2 83010 92925
0 16921 5 1 1 16920
0 16922 7 1 2 16917 16921
0 16923 5 1 1 16922
0 16924 7 2 2 89536 16923
0 16925 7 1 2 86182 92927
0 16926 5 1 1 16925
0 16927 7 2 2 69779 92905
0 16928 7 1 2 68375 72999
0 16929 7 1 2 81604 16928
0 16930 7 2 2 92929 16929
0 16931 7 1 2 62549 92931
0 16932 5 1 1 16931
0 16933 7 1 2 16926 16932
0 16934 5 1 1 16933
0 16935 7 1 2 66095 16934
0 16936 5 1 1 16935
0 16937 7 6 2 64696 78675
0 16938 7 2 2 90490 92933
0 16939 7 8 2 61264 66444
0 16940 7 1 2 92939 92941
0 16941 5 1 1 16940
0 16942 7 2 2 81792 82777
0 16943 7 1 2 83298 92949
0 16944 5 1 1 16943
0 16945 7 1 2 16941 16944
0 16946 5 1 1 16945
0 16947 7 3 2 73418 82273
0 16948 7 1 2 74797 92951
0 16949 7 1 2 16946 16948
0 16950 5 1 1 16949
0 16951 7 1 2 16936 16950
0 16952 5 1 1 16951
0 16953 7 1 2 90702 16952
0 16954 5 1 1 16953
0 16955 7 1 2 83287 92455
0 16956 7 1 2 92950 16955
0 16957 5 1 1 16956
0 16958 7 1 2 82090 88174
0 16959 7 1 2 92940 16958
0 16960 5 1 1 16959
0 16961 7 1 2 16957 16960
0 16962 5 1 1 16961
0 16963 7 1 2 92952 16962
0 16964 5 1 1 16963
0 16965 7 13 2 61265 67771
0 16966 5 1 1 92954
0 16967 7 4 2 67426 67842
0 16968 7 7 2 66210 92967
0 16969 7 1 2 92955 92971
0 16970 7 1 2 92928 16969
0 16971 5 1 1 16970
0 16972 7 1 2 16964 16971
0 16973 5 1 1 16972
0 16974 7 1 2 74798 16973
0 16975 5 1 1 16974
0 16976 7 5 2 67843 91367
0 16977 5 1 1 92978
0 16978 7 2 2 90873 92979
0 16979 7 1 2 92983 92932
0 16980 5 1 1 16979
0 16981 7 1 2 16975 16980
0 16982 7 1 2 16954 16981
0 16983 5 1 1 16982
0 16984 7 1 2 64327 16983
0 16985 5 1 1 16984
0 16986 7 1 2 87349 78856
0 16987 5 1 1 16986
0 16988 7 1 2 3472 89276
0 16989 5 1 1 16988
0 16990 7 4 2 16987 16989
0 16991 5 1 1 92985
0 16992 7 2 2 64495 78068
0 16993 7 1 2 88783 92989
0 16994 5 1 1 16993
0 16995 7 4 2 65121 71220
0 16996 7 1 2 67987 88545
0 16997 7 1 2 92991 16996
0 16998 5 1 1 16997
0 16999 7 1 2 16994 16998
0 17000 5 1 1 16999
0 17001 7 1 2 77879 17000
0 17002 7 1 2 92666 17001
0 17003 5 1 1 17002
0 17004 7 4 2 67427 67772
0 17005 7 9 2 67664 67844
0 17006 7 4 2 92995 92999
0 17007 7 2 2 87658 93008
0 17008 7 10 2 68819 69175
0 17009 7 4 2 66096 93014
0 17010 7 4 2 66211 62385
0 17011 7 1 2 91277 93028
0 17012 7 1 2 93024 17011
0 17013 7 1 2 93012 17012
0 17014 5 1 1 17013
0 17015 7 1 2 17003 17014
0 17016 5 1 1 17015
0 17017 7 1 2 92986 17016
0 17018 5 1 1 17017
0 17019 7 17 2 64697 92764
0 17020 7 2 2 68820 82091
0 17021 7 1 2 81525 93049
0 17022 7 1 2 93032 17021
0 17023 7 1 2 78676 89095
0 17024 7 1 2 90703 17023
0 17025 7 1 2 17022 17024
0 17026 5 1 1 17025
0 17027 7 2 2 67227 67773
0 17028 7 8 2 67845 64496
0 17029 7 5 2 67428 69176
0 17030 7 1 2 93053 93061
0 17031 7 1 2 93051 17030
0 17032 7 1 2 88698 82822
0 17033 7 3 2 66212 66691
0 17034 7 3 2 92942 93066
0 17035 7 1 2 92934 93069
0 17036 7 1 2 17032 17035
0 17037 7 1 2 17031 17036
0 17038 5 1 1 17037
0 17039 7 1 2 65389 17038
0 17040 7 1 2 17026 17039
0 17041 7 1 2 17018 17040
0 17042 7 1 2 16985 17041
0 17043 5 1 1 17042
0 17044 7 2 2 67774 63768
0 17045 7 1 2 78705 93072
0 17046 7 3 2 64917 92765
0 17047 7 7 2 63130 81630
0 17048 7 1 2 93074 93077
0 17049 7 1 2 17045 17048
0 17050 5 1 1 17049
0 17051 7 4 2 62946 68376
0 17052 7 1 2 84215 93084
0 17053 7 57 2 64328 69354
0 17054 7 6 2 69780 93088
0 17055 7 1 2 91891 93145
0 17056 7 1 2 17052 17055
0 17057 5 1 1 17056
0 17058 7 1 2 17050 17057
0 17059 5 1 1 17058
0 17060 7 1 2 62386 17059
0 17061 5 1 1 17060
0 17062 7 7 2 62947 67988
0 17063 5 1 1 93151
0 17064 7 1 2 82412 82737
0 17065 7 1 2 93152 17064
0 17066 7 1 2 93146 17065
0 17067 7 1 2 91597 17066
0 17068 5 1 1 17067
0 17069 7 1 2 17061 17068
0 17070 5 1 1 17069
0 17071 7 1 2 83585 17070
0 17072 5 1 1 17071
0 17073 7 3 2 77062 79358
0 17074 7 8 2 63532 64329
0 17075 7 7 2 67665 62948
0 17076 7 2 2 93161 93169
0 17077 7 1 2 92063 93176
0 17078 7 1 2 90186 17077
0 17079 7 1 2 93158 17078
0 17080 5 1 1 17079
0 17081 7 1 2 17072 17080
0 17082 5 1 1 17081
0 17083 7 1 2 90653 17082
0 17084 5 1 1 17083
0 17085 7 5 2 63533 73419
0 17086 7 3 2 93159 93178
0 17087 7 1 2 89151 93183
0 17088 5 1 1 17087
0 17089 7 1 2 62550 83586
0 17090 7 1 2 88072 17089
0 17091 5 1 1 17090
0 17092 7 1 2 74032 83996
0 17093 7 1 2 91060 17092
0 17094 5 1 1 17093
0 17095 7 1 2 17091 17094
0 17096 5 1 1 17095
0 17097 7 1 2 67228 17096
0 17098 5 1 1 17097
0 17099 7 1 2 80135 93184
0 17100 5 1 1 17099
0 17101 7 2 2 83587 81863
0 17102 7 2 2 91398 93186
0 17103 7 1 2 73912 93188
0 17104 5 1 1 17103
0 17105 7 1 2 17100 17104
0 17106 7 1 2 17098 17105
0 17107 5 1 1 17106
0 17108 7 1 2 82738 17107
0 17109 5 1 1 17108
0 17110 7 1 2 17088 17109
0 17111 5 1 1 17110
0 17112 7 8 2 64330 69781
0 17113 7 1 2 90640 93190
0 17114 7 1 2 17111 17113
0 17115 5 1 1 17114
0 17116 7 1 2 17084 17115
0 17117 5 1 1 17116
0 17118 7 1 2 61535 17117
0 17119 5 1 1 17118
0 17120 7 2 2 75701 83567
0 17121 7 1 2 93160 93198
0 17122 5 1 1 17121
0 17123 7 2 2 83588 84211
0 17124 7 1 2 82256 93200
0 17125 7 1 2 90187 17124
0 17126 5 1 1 17125
0 17127 7 1 2 17122 17126
0 17128 5 1 1 17127
0 17129 7 4 2 64331 90704
0 17130 7 1 2 73420 92020
0 17131 7 1 2 93202 17130
0 17132 7 1 2 17128 17131
0 17133 5 1 1 17132
0 17134 7 1 2 17119 17133
0 17135 5 1 1 17134
0 17136 7 1 2 66097 17135
0 17137 5 1 1 17136
0 17138 7 2 2 64497 71933
0 17139 7 1 2 80785 91552
0 17140 7 1 2 93206 17139
0 17141 5 1 1 17140
0 17142 7 1 2 73000 83455
0 17143 7 1 2 93187 17142
0 17144 5 1 1 17143
0 17145 7 1 2 17141 17144
0 17146 5 1 1 17145
0 17147 7 1 2 67429 17146
0 17148 5 1 1 17147
0 17149 7 1 2 91447 91556
0 17150 5 1 1 17149
0 17151 7 1 2 17148 17150
0 17152 5 1 1 17151
0 17153 7 1 2 90188 17152
0 17154 5 1 1 17153
0 17155 7 2 2 64498 90914
0 17156 7 1 2 87063 73421
0 17157 7 1 2 80136 17156
0 17158 7 1 2 93208 17157
0 17159 5 2 1 17158
0 17160 7 1 2 90043 93201
0 17161 7 1 2 91598 17160
0 17162 5 1 1 17161
0 17163 7 1 2 93210 17162
0 17164 5 1 1 17163
0 17165 7 1 2 67229 17164
0 17166 5 1 1 17165
0 17167 7 1 2 81853 93189
0 17168 5 1 1 17167
0 17169 7 1 2 93211 17168
0 17170 5 1 1 17169
0 17171 7 1 2 68614 17170
0 17172 5 1 1 17171
0 17173 7 1 2 17166 17172
0 17174 7 1 2 17154 17173
0 17175 5 1 1 17174
0 17176 7 1 2 92456 93191
0 17177 7 1 2 17175 17176
0 17178 5 1 1 17177
0 17179 7 1 2 70310 17178
0 17180 7 1 2 17137 17179
0 17181 5 1 1 17180
0 17182 7 1 2 65714 17181
0 17183 7 1 2 17043 17182
0 17184 5 1 1 17183
0 17185 7 1 2 16908 17184
0 17186 5 1 1 17185
0 17187 7 1 2 72124 17186
0 17188 5 1 1 17187
0 17189 7 1 2 66925 17188
0 17190 5 1 1 17189
0 17191 7 1 2 71313 88390
0 17192 5 1 1 17191
0 17193 7 1 2 88184 73311
0 17194 5 1 1 17193
0 17195 7 1 2 17192 17194
0 17196 5 1 1 17195
0 17197 7 1 2 76426 17196
0 17198 5 1 1 17197
0 17199 7 4 2 62813 76042
0 17200 7 1 2 79541 85537
0 17201 7 1 2 93212 17200
0 17202 5 1 1 17201
0 17203 7 1 2 17198 17202
0 17204 5 1 1 17203
0 17205 7 1 2 81315 17204
0 17206 5 1 1 17205
0 17207 7 1 2 74640 86944
0 17208 5 1 1 17207
0 17209 7 5 2 66445 80241
0 17210 5 1 1 93216
0 17211 7 3 2 77941 73825
0 17212 7 1 2 93217 93221
0 17213 5 1 1 17212
0 17214 7 1 2 17208 17213
0 17215 5 1 1 17214
0 17216 7 1 2 71221 17215
0 17217 5 1 1 17216
0 17218 7 1 2 72532 72247
0 17219 5 2 1 17218
0 17220 7 1 2 74739 93224
0 17221 5 1 1 17220
0 17222 7 1 2 62551 17221
0 17223 5 1 1 17222
0 17224 7 2 2 74726 17223
0 17225 7 1 2 74731 86724
0 17226 5 1 1 17225
0 17227 7 1 2 93226 17226
0 17228 5 3 1 17227
0 17229 7 1 2 81913 93228
0 17230 5 1 1 17229
0 17231 7 2 2 80163 76752
0 17232 7 1 2 61536 93231
0 17233 5 1 1 17232
0 17234 7 1 2 17230 17233
0 17235 5 1 1 17234
0 17236 7 1 2 76398 17235
0 17237 5 1 1 17236
0 17238 7 1 2 17217 17237
0 17239 5 1 1 17238
0 17240 7 1 2 70020 17239
0 17241 5 1 1 17240
0 17242 7 1 2 85491 88084
0 17243 7 1 2 92357 17242
0 17244 5 1 1 17243
0 17245 7 1 2 17241 17244
0 17246 5 1 1 17245
0 17247 7 1 2 63131 17246
0 17248 5 1 1 17247
0 17249 7 1 2 70021 93229
0 17250 5 1 1 17249
0 17251 7 4 2 73312 74982
0 17252 7 1 2 76939 93233
0 17253 5 1 1 17252
0 17254 7 1 2 17250 17253
0 17255 5 1 1 17254
0 17256 7 1 2 62387 17255
0 17257 5 1 1 17256
0 17258 7 3 2 84448 77942
0 17259 7 1 2 85363 93237
0 17260 5 1 1 17259
0 17261 7 1 2 17257 17260
0 17262 5 1 1 17261
0 17263 7 1 2 92352 17262
0 17264 5 1 1 17263
0 17265 7 1 2 17248 17264
0 17266 5 1 1 17265
0 17267 7 1 2 68145 17266
0 17268 5 1 1 17267
0 17269 7 1 2 77440 90828
0 17270 7 2 2 63534 73960
0 17271 7 3 2 88095 84449
0 17272 7 1 2 93240 93242
0 17273 7 1 2 17269 17272
0 17274 5 1 1 17273
0 17275 7 1 2 17268 17274
0 17276 5 1 1 17275
0 17277 7 1 2 69782 17276
0 17278 5 1 1 17277
0 17279 7 1 2 17206 17278
0 17280 5 1 1 17279
0 17281 7 1 2 64499 17280
0 17282 5 1 1 17281
0 17283 7 4 2 85894 80233
0 17284 7 2 2 90527 93245
0 17285 7 3 2 69783 76886
0 17286 7 4 2 63535 82881
0 17287 7 1 2 93251 93254
0 17288 5 1 1 17287
0 17289 7 1 2 62388 84604
0 17290 7 1 2 81316 17289
0 17291 5 1 1 17290
0 17292 7 1 2 17288 17291
0 17293 5 1 1 17292
0 17294 7 1 2 93249 17293
0 17295 5 1 1 17294
0 17296 7 1 2 61831 17295
0 17297 7 1 2 17282 17296
0 17298 5 1 1 17297
0 17299 7 1 2 83997 85397
0 17300 5 1 1 17299
0 17301 7 2 2 88898 91452
0 17302 7 1 2 87064 77943
0 17303 7 1 2 93258 17302
0 17304 5 1 1 17303
0 17305 7 1 2 17300 17304
0 17306 5 1 1 17305
0 17307 7 1 2 82193 17306
0 17308 5 1 1 17307
0 17309 7 1 2 14230 93227
0 17310 5 1 1 17309
0 17311 7 1 2 62389 17310
0 17312 5 1 1 17311
0 17313 7 1 2 73860 92370
0 17314 5 1 1 17313
0 17315 7 1 2 17312 17314
0 17316 5 1 1 17315
0 17317 7 1 2 79388 80737
0 17318 7 1 2 17316 17317
0 17319 5 1 1 17318
0 17320 7 1 2 17308 17319
0 17321 5 1 1 17320
0 17322 7 1 2 66446 17321
0 17323 5 1 1 17322
0 17324 7 1 2 78876 74641
0 17325 5 1 1 17324
0 17326 7 1 2 91160 93222
0 17327 5 1 1 17326
0 17328 7 1 2 17325 17327
0 17329 5 1 1 17328
0 17330 7 1 2 71222 17329
0 17331 5 1 1 17330
0 17332 7 1 2 63132 93232
0 17333 5 1 1 17332
0 17334 7 1 2 78919 93230
0 17335 5 1 1 17334
0 17336 7 1 2 17333 17335
0 17337 5 1 1 17336
0 17338 7 1 2 76399 17337
0 17339 5 1 1 17338
0 17340 7 1 2 17331 17339
0 17341 5 1 1 17340
0 17342 7 1 2 70022 17341
0 17343 5 1 1 17342
0 17344 7 1 2 64698 78695
0 17345 7 1 2 78130 17344
0 17346 7 1 2 77514 17345
0 17347 5 1 1 17346
0 17348 7 1 2 17343 17347
0 17349 5 1 1 17348
0 17350 7 1 2 82847 17349
0 17351 5 1 1 17350
0 17352 7 1 2 17323 17351
0 17353 5 1 1 17352
0 17354 7 1 2 81414 17353
0 17355 5 1 1 17354
0 17356 7 1 2 81045 81278
0 17357 7 1 2 79813 17356
0 17358 7 3 2 61537 77441
0 17359 7 2 2 80204 79439
0 17360 5 1 1 93263
0 17361 7 1 2 93260 93264
0 17362 7 1 2 17357 17361
0 17363 5 1 1 17362
0 17364 7 1 2 66692 17363
0 17365 7 1 2 17355 17364
0 17366 5 1 1 17365
0 17367 7 1 2 63769 17366
0 17368 7 1 2 17298 17367
0 17369 5 1 1 17368
0 17370 7 1 2 82527 90367
0 17371 5 1 1 17370
0 17372 7 1 2 74751 91951
0 17373 5 1 1 17372
0 17374 7 1 2 17371 17373
0 17375 5 1 1 17374
0 17376 7 1 2 88185 17375
0 17377 5 1 1 17376
0 17378 7 2 2 67230 84567
0 17379 5 2 1 93265
0 17380 7 1 2 87038 93266
0 17381 5 1 1 17380
0 17382 7 2 2 86945 80113
0 17383 7 1 2 90134 93269
0 17384 7 1 2 17381 17383
0 17385 5 1 1 17384
0 17386 7 1 2 17377 17385
0 17387 5 1 1 17386
0 17388 7 1 2 83106 17387
0 17389 5 1 1 17388
0 17390 7 1 2 85961 80646
0 17391 7 2 2 78506 80164
0 17392 7 1 2 89967 93271
0 17393 7 1 2 17390 17392
0 17394 5 1 1 17393
0 17395 7 1 2 17389 17394
0 17396 5 1 1 17395
0 17397 7 1 2 69784 17396
0 17398 5 1 1 17397
0 17399 7 3 2 80045 89360
0 17400 5 1 1 93273
0 17401 7 1 2 72887 93274
0 17402 5 1 1 17401
0 17403 7 7 2 64699 88347
0 17404 5 1 1 93276
0 17405 7 2 2 84010 93277
0 17406 5 1 1 93283
0 17407 7 1 2 17402 17406
0 17408 5 1 1 17407
0 17409 7 1 2 71934 17408
0 17410 5 1 1 17409
0 17411 7 1 2 90567 87228
0 17412 5 1 1 17411
0 17413 7 1 2 17410 17412
0 17414 5 1 1 17413
0 17415 7 1 2 67430 17414
0 17416 5 1 1 17415
0 17417 7 13 2 65390 71314
0 17418 5 2 1 93285
0 17419 7 1 2 85941 93286
0 17420 5 1 1 17419
0 17421 7 1 2 80895 74511
0 17422 5 1 1 17421
0 17423 7 1 2 17420 17422
0 17424 5 1 1 17423
0 17425 7 1 2 86946 17424
0 17426 5 1 1 17425
0 17427 7 1 2 17416 17426
0 17428 5 1 1 17427
0 17429 7 1 2 82373 75998
0 17430 7 1 2 17428 17429
0 17431 5 1 1 17430
0 17432 7 1 2 17398 17431
0 17433 5 1 1 17432
0 17434 7 1 2 64500 17433
0 17435 5 1 1 17434
0 17436 7 4 2 73161 72321
0 17437 5 2 1 93300
0 17438 7 1 2 91122 93301
0 17439 5 1 1 17438
0 17440 7 1 2 84336 74688
0 17441 5 1 1 17440
0 17442 7 1 2 17439 17441
0 17443 5 1 1 17442
0 17444 7 5 2 79440 79935
0 17445 7 1 2 89054 93306
0 17446 7 1 2 17443 17445
0 17447 5 1 1 17446
0 17448 7 1 2 17435 17447
0 17449 5 1 1 17448
0 17450 7 1 2 78069 17449
0 17451 5 1 1 17450
0 17452 7 1 2 71223 83288
0 17453 7 1 2 85962 17452
0 17454 7 1 2 88057 17453
0 17455 5 1 1 17454
0 17456 7 1 2 64501 92987
0 17457 5 1 1 17456
0 17458 7 1 2 4360 17457
0 17459 5 1 1 17458
0 17460 7 1 2 74983 77623
0 17461 7 1 2 17459 17460
0 17462 5 1 1 17461
0 17463 7 1 2 17455 17462
0 17464 5 1 1 17463
0 17465 7 1 2 70311 17464
0 17466 5 1 1 17465
0 17467 7 1 2 88688 77704
0 17468 7 2 2 81667 83889
0 17469 7 1 2 85538 93311
0 17470 7 1 2 17467 17469
0 17471 5 1 1 17470
0 17472 7 1 2 17466 17471
0 17473 5 1 1 17472
0 17474 7 1 2 81793 17473
0 17475 5 1 1 17474
0 17476 7 2 2 71224 92011
0 17477 5 2 1 93313
0 17478 7 1 2 91123 93314
0 17479 5 1 1 17478
0 17480 7 1 2 80849 91459
0 17481 5 1 1 17480
0 17482 7 1 2 17479 17481
0 17483 5 1 1 17482
0 17484 7 1 2 72781 17483
0 17485 5 1 1 17484
0 17486 7 3 2 71315 81086
0 17487 5 1 1 93317
0 17488 7 1 2 15010 17487
0 17489 5 1 1 17488
0 17490 7 1 2 85942 17489
0 17491 5 1 1 17490
0 17492 7 1 2 17485 17491
0 17493 5 1 1 17492
0 17494 7 1 2 79751 76774
0 17495 7 1 2 85172 17494
0 17496 7 1 2 17493 17495
0 17497 5 1 1 17496
0 17498 7 1 2 17475 17497
0 17499 7 1 2 17451 17498
0 17500 7 1 2 17369 17499
0 17501 5 1 1 17500
0 17502 7 1 2 70667 17501
0 17503 5 1 1 17502
0 17504 7 1 2 77868 80417
0 17505 5 1 1 17504
0 17506 7 1 2 78920 91634
0 17507 5 1 1 17506
0 17508 7 1 2 17505 17507
0 17509 5 1 1 17508
0 17510 7 1 2 75608 17509
0 17511 5 1 1 17510
0 17512 7 2 2 62390 77869
0 17513 5 2 1 93320
0 17514 7 1 2 75527 85813
0 17515 5 1 1 17514
0 17516 7 1 2 93322 17515
0 17517 5 1 1 17516
0 17518 7 1 2 88867 17517
0 17519 5 1 1 17518
0 17520 7 1 2 17511 17519
0 17521 5 1 1 17520
0 17522 7 1 2 64106 17521
0 17523 5 1 1 17522
0 17524 7 2 2 86003 80418
0 17525 5 1 1 93324
0 17526 7 1 2 74689 93325
0 17527 5 1 1 17526
0 17528 7 1 2 17523 17527
0 17529 5 1 1 17528
0 17530 7 1 2 83544 17529
0 17531 5 1 1 17530
0 17532 7 2 2 65968 80738
0 17533 7 1 2 81893 93326
0 17534 5 1 1 17533
0 17535 7 1 2 76319 78877
0 17536 5 1 1 17535
0 17537 7 1 2 71225 83232
0 17538 5 1 1 17537
0 17539 7 1 2 17536 17538
0 17540 5 1 1 17539
0 17541 7 1 2 74883 73422
0 17542 7 1 2 17540 17541
0 17543 5 1 1 17542
0 17544 7 1 2 17534 17543
0 17545 5 1 1 17544
0 17546 7 1 2 67231 17545
0 17547 5 1 1 17546
0 17548 7 8 2 68377 65969
0 17549 5 1 1 93328
0 17550 7 2 2 78878 93329
0 17551 7 1 2 85219 15621
0 17552 5 1 1 17551
0 17553 7 1 2 93336 17552
0 17554 5 1 1 17553
0 17555 7 1 2 17547 17554
0 17556 5 1 1 17555
0 17557 7 1 2 68965 17556
0 17558 5 1 1 17557
0 17559 7 2 2 64700 80739
0 17560 5 1 1 93338
0 17561 7 1 2 62391 85554
0 17562 5 3 1 17561
0 17563 7 1 2 92354 93340
0 17564 5 1 1 17563
0 17565 7 1 2 93323 17564
0 17566 5 1 1 17565
0 17567 7 1 2 93339 17566
0 17568 5 1 1 17567
0 17569 7 1 2 17558 17568
0 17570 5 1 1 17569
0 17571 7 1 2 81297 17570
0 17572 5 1 1 17571
0 17573 7 1 2 17531 17572
0 17574 5 1 1 17573
0 17575 7 1 2 61538 17574
0 17576 5 1 1 17575
0 17577 7 1 2 62392 84742
0 17578 5 1 1 17577
0 17579 7 2 2 74033 79680
0 17580 7 1 2 17578 93343
0 17581 5 1 1 17580
0 17582 7 2 2 77900 75363
0 17583 5 1 1 93345
0 17584 7 1 2 82194 93346
0 17585 5 1 1 17584
0 17586 7 1 2 17581 17585
0 17587 5 1 1 17586
0 17588 7 1 2 81298 17587
0 17589 5 1 1 17588
0 17590 7 1 2 85784 14650
0 17591 5 1 1 17590
0 17592 7 1 2 75609 17591
0 17593 5 1 1 17592
0 17594 7 2 2 68615 76821
0 17595 7 1 2 84987 93347
0 17596 5 1 1 17595
0 17597 7 1 2 17593 17596
0 17598 5 1 1 17597
0 17599 7 1 2 64107 83545
0 17600 7 1 2 17598 17599
0 17601 5 1 1 17600
0 17602 7 1 2 17589 17601
0 17603 5 1 1 17602
0 17604 7 1 2 91483 17603
0 17605 5 1 1 17604
0 17606 7 1 2 17576 17605
0 17607 5 1 1 17606
0 17608 7 1 2 69785 17607
0 17609 5 1 1 17608
0 17610 7 1 2 82429 80098
0 17611 5 1 1 17610
0 17612 7 1 2 80520 82869
0 17613 5 1 1 17612
0 17614 7 1 2 17611 17613
0 17615 5 1 1 17614
0 17616 7 1 2 63133 17615
0 17617 5 1 1 17616
0 17618 7 1 2 88299 91274
0 17619 7 1 2 88789 17618
0 17620 5 1 1 17619
0 17621 7 1 2 17617 17620
0 17622 5 1 1 17621
0 17623 7 1 2 68821 17622
0 17624 5 1 1 17623
0 17625 7 1 2 88245 87972
0 17626 7 1 2 93078 17625
0 17627 5 1 1 17626
0 17628 7 1 2 17624 17627
0 17629 5 1 1 17628
0 17630 7 1 2 67666 17629
0 17631 5 1 1 17630
0 17632 7 2 2 78879 83224
0 17633 7 1 2 74269 83776
0 17634 7 1 2 93349 17633
0 17635 5 1 1 17634
0 17636 7 1 2 17631 17635
0 17637 5 1 1 17636
0 17638 7 1 2 67431 17637
0 17639 5 1 1 17638
0 17640 7 2 2 65970 74679
0 17641 7 1 2 72822 93351
0 17642 5 1 1 17641
0 17643 7 1 2 71506 17642
0 17644 5 1 1 17643
0 17645 7 1 2 65715 17644
0 17646 5 1 1 17645
0 17647 7 1 2 77901 88811
0 17648 5 1 1 17647
0 17649 7 1 2 17646 17648
0 17650 5 1 1 17649
0 17651 7 1 2 78880 81631
0 17652 7 1 2 17650 17651
0 17653 5 1 1 17652
0 17654 7 1 2 17639 17653
0 17655 5 1 1 17654
0 17656 7 1 2 70023 76588
0 17657 7 1 2 17655 17656
0 17658 5 1 1 17657
0 17659 7 1 2 17609 17658
0 17660 5 1 1 17659
0 17661 7 1 2 64502 17660
0 17662 5 1 1 17661
0 17663 7 2 2 80974 91672
0 17664 7 1 2 85220 85975
0 17665 5 4 1 17664
0 17666 7 2 2 71163 87618
0 17667 7 2 2 63298 93359
0 17668 5 1 1 93361
0 17669 7 1 2 93355 93362
0 17670 5 1 1 17669
0 17671 7 1 2 89223 89696
0 17672 7 1 2 92340 17671
0 17673 5 1 1 17672
0 17674 7 1 2 17670 17673
0 17675 5 1 1 17674
0 17676 7 1 2 93353 17675
0 17677 5 1 1 17676
0 17678 7 1 2 17662 17677
0 17679 5 1 1 17678
0 17680 7 1 2 65391 17679
0 17681 5 1 1 17680
0 17682 7 4 2 66447 80205
0 17683 7 1 2 91673 93363
0 17684 5 1 1 17683
0 17685 7 1 2 64503 88392
0 17686 5 1 1 17685
0 17687 7 1 2 17684 17686
0 17688 5 1 1 17687
0 17689 7 1 2 68966 17688
0 17690 5 1 1 17689
0 17691 7 1 2 91204 92599
0 17692 5 1 1 17691
0 17693 7 1 2 17690 17692
0 17694 5 1 1 17693
0 17695 7 1 2 63937 17694
0 17696 5 1 1 17695
0 17697 7 1 2 79359 77815
0 17698 7 1 2 88354 17697
0 17699 5 1 1 17698
0 17700 7 1 2 17696 17699
0 17701 5 1 1 17700
0 17702 7 1 2 81317 17701
0 17703 5 1 1 17702
0 17704 7 2 2 86947 78696
0 17705 5 1 1 93367
0 17706 7 1 2 72533 93368
0 17707 5 1 1 17706
0 17708 7 1 2 88186 80079
0 17709 5 1 1 17708
0 17710 7 1 2 17707 17709
0 17711 5 1 1 17710
0 17712 7 1 2 63938 17711
0 17713 5 1 1 17712
0 17714 7 1 2 91178 92095
0 17715 5 1 1 17714
0 17716 7 1 2 17713 17715
0 17717 5 1 1 17716
0 17718 7 1 2 81559 89711
0 17719 7 1 2 17717 17718
0 17720 5 1 1 17719
0 17721 7 1 2 17703 17720
0 17722 5 1 1 17721
0 17723 7 1 2 62552 17722
0 17724 5 1 1 17723
0 17725 7 1 2 78921 81318
0 17726 5 1 1 17725
0 17727 7 1 2 83438 82035
0 17728 5 1 1 17727
0 17729 7 1 2 17726 17728
0 17730 5 1 1 17729
0 17731 7 1 2 87176 88899
0 17732 7 1 2 73973 17731
0 17733 7 1 2 17730 17732
0 17734 5 1 1 17733
0 17735 7 1 2 17724 17734
0 17736 5 1 1 17735
0 17737 7 1 2 71820 17736
0 17738 5 1 1 17737
0 17739 7 1 2 17681 17738
0 17740 5 1 1 17739
0 17741 7 1 2 61832 17740
0 17742 5 1 1 17741
0 17743 7 5 2 66693 81415
0 17744 5 1 1 93369
0 17745 7 1 2 88246 90003
0 17746 5 1 1 17745
0 17747 7 1 2 92141 17746
0 17748 5 1 1 17747
0 17749 7 1 2 92320 17748
0 17750 5 1 1 17749
0 17751 7 1 2 81914 84774
0 17752 5 1 1 17751
0 17753 7 1 2 17750 17752
0 17754 5 1 1 17753
0 17755 7 1 2 74653 17754
0 17756 5 1 1 17755
0 17757 7 1 2 73313 89369
0 17758 5 1 1 17757
0 17759 7 1 2 86948 92431
0 17760 5 1 1 17759
0 17761 7 1 2 17758 17760
0 17762 5 1 1 17761
0 17763 7 1 2 62814 17762
0 17764 5 1 1 17763
0 17765 7 5 2 62553 73961
0 17766 5 1 1 93374
0 17767 7 1 2 91529 93375
0 17768 5 1 1 17767
0 17769 7 1 2 17764 17768
0 17770 5 1 1 17769
0 17771 7 1 2 76400 17770
0 17772 5 1 1 17771
0 17773 7 1 2 17756 17772
0 17774 5 1 1 17773
0 17775 7 1 2 65716 17774
0 17776 5 1 1 17775
0 17777 7 3 2 70902 93287
0 17778 7 1 2 92358 93379
0 17779 5 1 1 17778
0 17780 7 5 2 61539 75288
0 17781 7 2 2 88247 93382
0 17782 5 1 1 93387
0 17783 7 1 2 62554 93388
0 17784 5 1 1 17783
0 17785 7 1 2 17779 17784
0 17786 5 1 1 17785
0 17787 7 1 2 62393 73826
0 17788 7 1 2 17786 17787
0 17789 5 1 1 17788
0 17790 7 1 2 17776 17789
0 17791 5 1 1 17790
0 17792 7 1 2 63134 17791
0 17793 5 1 1 17792
0 17794 7 2 2 63939 71653
0 17795 5 1 1 93389
0 17796 7 1 2 86493 17795
0 17797 5 1 1 17796
0 17798 7 1 2 62555 17797
0 17799 5 1 1 17798
0 17800 7 2 2 72043 74487
0 17801 5 3 1 93391
0 17802 7 1 2 17799 93393
0 17803 5 1 1 17802
0 17804 7 1 2 62815 17803
0 17805 5 1 1 17804
0 17806 7 1 2 92337 17805
0 17807 5 1 1 17806
0 17808 7 1 2 90220 80637
0 17809 7 1 2 17807 17808
0 17810 5 1 1 17809
0 17811 7 1 2 17793 17810
0 17812 5 1 1 17811
0 17813 7 1 2 64504 17812
0 17814 5 1 1 17813
0 17815 7 4 2 66448 72696
0 17816 7 1 2 76365 92600
0 17817 7 1 2 93396 17816
0 17818 7 1 2 80452 17817
0 17819 5 1 1 17818
0 17820 7 1 2 17814 17819
0 17821 5 1 1 17820
0 17822 7 1 2 63770 17821
0 17823 5 1 1 17822
0 17824 7 3 2 69546 80834
0 17825 5 1 1 93400
0 17826 7 1 2 61540 91660
0 17827 5 2 1 17826
0 17828 7 1 2 16786 93403
0 17829 5 1 1 17828
0 17830 7 1 2 73549 17829
0 17831 5 1 1 17830
0 17832 7 1 2 17825 17831
0 17833 5 1 1 17832
0 17834 7 1 2 79681 17833
0 17835 5 1 1 17834
0 17836 7 4 2 61541 88248
0 17837 5 1 1 93405
0 17838 7 4 2 71126 73314
0 17839 7 1 2 93406 93409
0 17840 5 1 1 17839
0 17841 7 1 2 17835 17840
0 17842 5 1 1 17841
0 17843 7 1 2 63135 17842
0 17844 5 1 1 17843
0 17845 7 2 2 61542 80442
0 17846 7 2 2 65717 80187
0 17847 7 1 2 93413 93415
0 17848 5 1 1 17847
0 17849 7 1 2 17844 17848
0 17850 5 1 1 17849
0 17851 7 2 2 75947 83650
0 17852 7 1 2 17850 93417
0 17853 5 1 1 17852
0 17854 7 1 2 17823 17853
0 17855 5 1 1 17854
0 17856 7 1 2 70024 17855
0 17857 5 1 1 17856
0 17858 7 1 2 77851 87571
0 17859 7 1 2 91484 17858
0 17860 7 4 2 65122 75451
0 17861 7 5 2 63940 84513
0 17862 7 1 2 93419 93423
0 17863 7 1 2 17859 17862
0 17864 5 1 1 17863
0 17865 7 1 2 17857 17864
0 17866 5 1 1 17865
0 17867 7 1 2 93370 17866
0 17868 5 1 1 17867
0 17869 7 2 2 71226 74073
0 17870 5 3 1 93428
0 17871 7 1 2 92048 93430
0 17872 5 1 1 17871
0 17873 7 1 2 16694 17872
0 17874 5 1 1 17873
0 17875 7 1 2 79014 72823
0 17876 7 1 2 17874 17875
0 17877 5 1 1 17876
0 17878 7 1 2 72824 86949
0 17879 5 2 1 17878
0 17880 7 1 2 67667 92359
0 17881 5 1 1 17880
0 17882 7 1 2 93433 17881
0 17883 5 3 1 17882
0 17884 7 1 2 91326 85562
0 17885 7 1 2 93435 17884
0 17886 5 1 1 17885
0 17887 7 1 2 17877 17886
0 17888 5 1 1 17887
0 17889 7 1 2 65971 17888
0 17890 5 1 1 17889
0 17891 7 1 2 81915 85294
0 17892 5 1 1 17891
0 17893 7 1 2 89948 79688
0 17894 5 1 1 17893
0 17895 7 1 2 86950 17894
0 17896 5 1 1 17895
0 17897 7 1 2 17892 17896
0 17898 5 1 1 17897
0 17899 7 1 2 82966 17898
0 17900 5 1 1 17899
0 17901 7 1 2 81916 78191
0 17902 7 1 2 71164 17901
0 17903 7 1 2 88532 17902
0 17904 5 1 1 17903
0 17905 7 1 2 17900 17904
0 17906 5 1 1 17905
0 17907 7 1 2 71429 17906
0 17908 5 1 1 17907
0 17909 7 3 2 65718 71052
0 17910 5 1 1 93438
0 17911 7 3 2 88410 90004
0 17912 5 1 1 93441
0 17913 7 2 2 70025 72322
0 17914 5 1 1 93444
0 17915 7 1 2 71935 91227
0 17916 7 1 2 93445 17915
0 17917 5 1 1 17916
0 17918 7 1 2 17912 17917
0 17919 5 1 1 17918
0 17920 7 1 2 93439 17919
0 17921 5 1 1 17920
0 17922 7 1 2 17908 17921
0 17923 7 1 2 17890 17922
0 17924 5 1 1 17923
0 17925 7 1 2 63536 17924
0 17926 5 1 1 17925
0 17927 7 1 2 81917 85595
0 17928 5 1 1 17927
0 17929 7 1 2 70668 77531
0 17930 5 2 1 17929
0 17931 7 1 2 81918 93446
0 17932 5 1 1 17931
0 17933 7 2 2 70903 84889
0 17934 7 1 2 86951 93448
0 17935 5 1 1 17934
0 17936 7 1 2 17932 17935
0 17937 5 1 1 17936
0 17938 7 1 2 74799 17937
0 17939 5 1 1 17938
0 17940 7 1 2 17928 17939
0 17941 5 1 1 17940
0 17942 7 1 2 76442 89144
0 17943 7 1 2 17941 17942
0 17944 5 1 1 17943
0 17945 7 1 2 17926 17944
0 17946 5 1 1 17945
0 17947 7 1 2 63299 17946
0 17948 5 1 1 17947
0 17949 7 3 2 78070 77195
0 17950 7 1 2 80080 93450
0 17951 5 1 1 17950
0 17952 7 1 2 81046 78507
0 17953 7 1 2 78000 17952
0 17954 5 1 1 17953
0 17955 7 1 2 17951 17954
0 17956 5 1 1 17955
0 17957 7 1 2 88533 17956
0 17958 5 1 1 17957
0 17959 7 1 2 85249 77733
0 17960 5 4 1 17959
0 17961 7 1 2 71654 93453
0 17962 5 1 1 17961
0 17963 7 1 2 86121 17962
0 17964 5 1 1 17963
0 17965 7 2 2 65972 81047
0 17966 7 2 2 17964 93457
0 17967 7 1 2 78508 93459
0 17968 5 1 1 17967
0 17969 7 1 2 17958 17968
0 17970 5 1 1 17969
0 17971 7 1 2 90408 17970
0 17972 5 1 1 17971
0 17973 7 1 2 17948 17972
0 17974 5 1 1 17973
0 17975 7 1 2 63136 17974
0 17976 5 1 1 17975
0 17977 7 1 2 71165 89378
0 17978 5 1 1 17977
0 17979 7 1 2 89374 17978
0 17980 5 1 1 17979
0 17981 7 1 2 65719 17980
0 17982 5 1 1 17981
0 17983 7 1 2 85876 85173
0 17984 5 1 1 17983
0 17985 7 1 2 17982 17984
0 17986 5 1 1 17985
0 17987 7 1 2 88534 17986
0 17988 5 1 1 17987
0 17989 7 1 2 82374 93460
0 17990 5 1 1 17989
0 17991 7 1 2 17988 17990
0 17992 5 1 1 17991
0 17993 7 1 2 76043 82778
0 17994 7 1 2 17992 17993
0 17995 5 1 1 17994
0 17996 7 1 2 17976 17995
0 17997 5 1 1 17996
0 17998 7 1 2 64505 17997
0 17999 5 1 1 17998
0 18000 7 3 2 67668 81581
0 18001 7 3 2 80348 84498
0 18002 7 1 2 93461 93464
0 18003 5 1 1 18002
0 18004 7 1 2 17668 18003
0 18005 5 1 1 18004
0 18006 7 1 2 61833 18005
0 18007 5 1 1 18006
0 18008 7 1 2 81445 74432
0 18009 7 1 2 93465 18008
0 18010 5 1 1 18009
0 18011 7 1 2 18007 18010
0 18012 5 1 1 18011
0 18013 7 1 2 86170 18012
0 18014 5 1 1 18013
0 18015 7 1 2 82135 82050
0 18016 7 1 2 93360 18015
0 18017 5 1 1 18016
0 18018 7 1 2 18014 18017
0 18019 5 1 1 18018
0 18020 7 1 2 93354 18019
0 18021 5 1 1 18020
0 18022 7 1 2 17999 18021
0 18023 5 1 1 18022
0 18024 7 1 2 70312 18023
0 18025 5 1 1 18024
0 18026 7 2 2 76940 82779
0 18027 7 1 2 76443 93467
0 18028 7 2 2 85563 18027
0 18029 7 1 2 67989 93469
0 18030 5 1 1 18029
0 18031 7 1 2 89805 15402
0 18032 5 1 1 18031
0 18033 7 1 2 68378 18032
0 18034 5 1 1 18033
0 18035 7 4 2 76887 74884
0 18036 5 1 1 93471
0 18037 7 1 2 64918 93472
0 18038 5 1 1 18037
0 18039 7 1 2 18034 18038
0 18040 5 1 1 18039
0 18041 7 1 2 78881 80003
0 18042 7 1 2 18040 18041
0 18043 5 1 1 18042
0 18044 7 1 2 18030 18043
0 18045 5 1 1 18044
0 18046 7 1 2 63300 18045
0 18047 5 1 1 18046
0 18048 7 2 2 83497 79856
0 18049 5 1 1 93475
0 18050 7 1 2 91526 93476
0 18051 7 1 2 91629 18050
0 18052 5 1 1 18051
0 18053 7 1 2 18047 18052
0 18054 5 1 1 18053
0 18055 7 1 2 61543 18054
0 18056 5 1 1 18055
0 18057 7 4 2 63301 76080
0 18058 7 1 2 93470 93477
0 18059 5 1 1 18058
0 18060 7 1 2 18056 18059
0 18061 5 1 1 18060
0 18062 7 1 2 82274 18061
0 18063 5 1 1 18062
0 18064 7 4 2 70026 73001
0 18065 7 5 2 62556 76699
0 18066 5 2 1 93485
0 18067 7 1 2 86474 93490
0 18068 5 6 1 18067
0 18069 7 2 2 93481 93492
0 18070 7 1 2 68146 93498
0 18071 5 1 1 18070
0 18072 7 1 2 81299 79500
0 18073 7 1 2 86357 18072
0 18074 5 1 1 18073
0 18075 7 1 2 18071 18074
0 18076 5 1 1 18075
0 18077 7 1 2 89616 18076
0 18078 5 1 1 18077
0 18079 7 1 2 75999 86477
0 18080 7 1 2 91957 18079
0 18081 5 1 1 18080
0 18082 7 1 2 18078 18081
0 18083 5 1 1 18082
0 18084 7 1 2 90260 18083
0 18085 5 1 1 18084
0 18086 7 1 2 18063 18085
0 18087 5 1 1 18086
0 18088 7 1 2 61834 18087
0 18089 5 1 1 18088
0 18090 7 1 2 82870 92012
0 18091 7 1 2 93499 18090
0 18092 5 1 1 18091
0 18093 7 3 2 70313 92079
0 18094 5 2 1 93500
0 18095 7 1 2 81785 91448
0 18096 7 1 2 93501 18095
0 18097 5 1 1 18096
0 18098 7 1 2 18092 18097
0 18099 5 1 1 18098
0 18100 7 1 2 71430 18099
0 18101 5 1 1 18100
0 18102 7 1 2 18089 18101
0 18103 5 1 1 18102
0 18104 7 1 2 72125 18103
0 18105 5 1 1 18104
0 18106 7 1 2 18025 18105
0 18107 7 1 2 17868 18106
0 18108 7 1 2 17742 18107
0 18109 7 1 2 17503 18108
0 18110 5 1 1 18109
0 18111 7 1 2 92667 18110
0 18112 5 1 1 18111
0 18113 7 1 2 73827 92442
0 18114 5 1 1 18113
0 18115 7 1 2 86207 93179
0 18116 5 2 1 18115
0 18117 7 1 2 18114 93505
0 18118 5 1 1 18117
0 18119 7 1 2 92668 18118
0 18120 5 1 1 18119
0 18121 7 4 2 68379 73204
0 18122 5 1 1 93507
0 18123 7 5 2 69177 92639
0 18124 7 3 2 90654 93511
0 18125 7 1 2 93508 93516
0 18126 7 1 2 73179 18125
0 18127 5 1 1 18126
0 18128 7 1 2 18120 18127
0 18129 5 1 1 18128
0 18130 7 1 2 70314 18129
0 18131 5 1 1 18130
0 18132 7 4 2 73423 74654
0 18133 7 2 2 92669 93519
0 18134 5 1 1 93523
0 18135 7 1 2 71114 93524
0 18136 5 1 1 18135
0 18137 7 1 2 18131 18136
0 18138 5 1 1 18137
0 18139 7 1 2 70027 18138
0 18140 5 1 1 18139
0 18141 7 5 2 71316 92465
0 18142 7 2 2 64332 93525
0 18143 5 1 1 93530
0 18144 7 2 2 62816 78131
0 18145 7 1 2 74704 93532
0 18146 7 1 2 93531 18145
0 18147 5 1 1 18146
0 18148 7 1 2 18140 18147
0 18149 5 1 1 18148
0 18150 7 1 2 88187 18149
0 18151 5 1 1 18150
0 18152 7 2 2 72534 92466
0 18153 7 2 2 71227 74921
0 18154 5 1 1 93536
0 18155 7 2 2 85117 18154
0 18156 7 1 2 93162 93538
0 18157 7 1 2 93534 18156
0 18158 5 1 1 18157
0 18159 7 5 2 72044 73205
0 18160 5 1 1 93540
0 18161 7 4 2 86725 78323
0 18162 5 1 1 93545
0 18163 7 8 2 71573 93546
0 18164 5 2 1 93549
0 18165 7 1 2 62557 93550
0 18166 5 1 1 18165
0 18167 7 3 2 18160 18166
0 18168 5 11 1 93559
0 18169 7 5 2 67846 68380
0 18170 7 2 2 69178 93573
0 18171 7 6 2 66213 62817
0 18172 7 1 2 92663 93580
0 18173 7 1 2 93578 18172
0 18174 7 1 2 93562 18173
0 18175 5 1 1 18174
0 18176 7 1 2 18158 18175
0 18177 5 1 1 18176
0 18178 7 1 2 77234 83589
0 18179 7 1 2 18177 18178
0 18180 5 1 1 18179
0 18181 7 1 2 18151 18180
0 18182 5 1 1 18181
0 18183 7 1 2 64506 18182
0 18184 5 1 1 18183
0 18185 7 27 2 62949 64333
0 18186 5 8 1 93586
0 18187 7 1 2 74655 87125
0 18188 5 2 1 18187
0 18189 7 1 2 84290 86645
0 18190 5 1 1 18189
0 18191 7 1 2 93621 18190
0 18192 5 1 1 18191
0 18193 7 1 2 93587 18192
0 18194 5 1 1 18193
0 18195 7 11 2 64334 70669
0 18196 7 3 2 62950 93623
0 18197 5 3 1 93634
0 18198 7 6 2 69179 90874
0 18199 7 1 2 78445 73945
0 18200 7 1 2 93640 18199
0 18201 5 1 1 18200
0 18202 7 1 2 93637 18201
0 18203 5 1 1 18202
0 18204 7 1 2 63941 75914
0 18205 7 1 2 18203 18204
0 18206 5 1 1 18205
0 18207 7 1 2 18194 18206
0 18208 5 1 1 18207
0 18209 7 1 2 90655 18208
0 18210 5 1 1 18209
0 18211 7 3 2 71317 75915
0 18212 5 1 1 93646
0 18213 7 1 2 85081 93647
0 18214 5 1 1 18213
0 18215 7 1 2 93622 18214
0 18216 5 1 1 18215
0 18217 7 2 2 64335 18216
0 18218 7 1 2 90641 93649
0 18219 5 1 1 18218
0 18220 7 1 2 18210 18219
0 18221 5 1 1 18220
0 18222 7 1 2 66098 18221
0 18223 5 1 1 18222
0 18224 7 1 2 92457 93650
0 18225 5 1 1 18224
0 18226 7 1 2 18223 18225
0 18227 5 1 1 18226
0 18228 7 1 2 72045 18227
0 18229 5 1 1 18228
0 18230 7 3 2 73605 86646
0 18231 5 3 1 93651
0 18232 7 1 2 70670 93652
0 18233 7 1 2 92670 18232
0 18234 5 1 1 18233
0 18235 7 1 2 18229 18234
0 18236 5 1 1 18235
0 18237 7 1 2 70028 18236
0 18238 5 1 1 18237
0 18239 7 5 2 63942 64336
0 18240 7 1 2 73713 93657
0 18241 7 1 2 85492 18240
0 18242 7 1 2 92467 18241
0 18243 5 1 1 18242
0 18244 7 1 2 18238 18243
0 18245 5 1 1 18244
0 18246 7 1 2 80975 79441
0 18247 7 1 2 18245 18246
0 18248 5 1 1 18247
0 18249 7 1 2 18184 18248
0 18250 5 1 1 18249
0 18251 7 1 2 83107 18250
0 18252 5 1 1 18251
0 18253 7 1 2 90765 87140
0 18254 5 1 1 18253
0 18255 7 1 2 86952 72879
0 18256 5 1 1 18255
0 18257 7 1 2 18254 18256
0 18258 5 1 1 18257
0 18259 7 1 2 83811 18258
0 18260 5 1 1 18259
0 18261 7 1 2 82325 88117
0 18262 7 1 2 85340 18261
0 18263 5 1 1 18262
0 18264 7 1 2 18260 18263
0 18265 5 1 1 18264
0 18266 7 1 2 73424 18265
0 18267 5 1 1 18266
0 18268 7 1 2 93288 93250
0 18269 5 1 1 18268
0 18270 7 1 2 18267 18269
0 18271 5 1 1 18270
0 18272 7 1 2 83410 18271
0 18273 5 1 1 18272
0 18274 7 1 2 80206 92601
0 18275 5 1 1 18274
0 18276 7 1 2 70671 81490
0 18277 5 1 1 18276
0 18278 7 1 2 18275 18277
0 18279 5 1 1 18278
0 18280 7 1 2 66449 18279
0 18281 5 1 1 18280
0 18282 7 3 2 79360 76044
0 18283 5 1 1 93662
0 18284 7 1 2 70672 93663
0 18285 5 1 1 18284
0 18286 7 1 2 18281 18285
0 18287 5 1 1 18286
0 18288 7 1 2 83727 85112
0 18289 7 1 2 18287 18288
0 18290 5 1 1 18289
0 18291 7 1 2 18273 18290
0 18292 5 1 1 18291
0 18293 7 1 2 65123 18292
0 18294 5 1 1 18293
0 18295 7 1 2 88348 85393
0 18296 7 3 2 67669 79361
0 18297 7 1 2 92691 93665
0 18298 7 1 2 18295 18297
0 18299 5 1 1 18298
0 18300 7 1 2 18294 18299
0 18301 5 1 1 18300
0 18302 7 1 2 92671 18301
0 18303 5 1 1 18302
0 18304 7 1 2 79494 85612
0 18305 5 3 1 18304
0 18306 7 2 2 79442 93668
0 18307 7 1 2 66450 93671
0 18308 5 1 1 18307
0 18309 7 1 2 92595 18308
0 18310 5 1 1 18309
0 18311 7 1 2 70673 18310
0 18312 5 1 1 18311
0 18313 7 4 2 62558 72046
0 18314 5 3 1 93673
0 18315 7 1 2 87323 93674
0 18316 5 1 1 18315
0 18317 7 1 2 18312 18316
0 18318 5 1 1 18317
0 18319 7 1 2 62818 18318
0 18320 5 1 1 18319
0 18321 7 1 2 64108 92622
0 18322 5 1 1 18321
0 18323 7 1 2 18320 18322
0 18324 5 1 1 18323
0 18325 7 1 2 63943 18324
0 18326 5 1 1 18325
0 18327 7 1 2 92628 18326
0 18328 5 1 1 18327
0 18329 7 2 2 70315 18328
0 18330 7 5 2 67847 68147
0 18331 7 3 2 67775 67990
0 18332 7 3 2 93682 93687
0 18333 7 9 2 63537 69180
0 18334 7 2 2 65124 93693
0 18335 7 1 2 92832 93702
0 18336 7 1 2 93690 18335
0 18337 7 1 2 93680 18336
0 18338 5 1 1 18337
0 18339 7 1 2 18303 18338
0 18340 5 1 1 18339
0 18341 7 1 2 61835 18340
0 18342 5 1 1 18341
0 18343 7 1 2 18252 18342
0 18344 5 1 1 18343
0 18345 7 1 2 69786 18344
0 18346 5 1 1 18345
0 18347 7 2 2 73425 92468
0 18348 7 3 2 64701 76888
0 18349 7 1 2 92003 93706
0 18350 5 1 1 18349
0 18351 7 7 2 70316 76320
0 18352 5 2 1 93709
0 18353 7 1 2 79362 93710
0 18354 7 1 2 87583 18353
0 18355 5 1 1 18354
0 18356 7 1 2 18350 18355
0 18357 5 1 1 18356
0 18358 7 1 2 68967 18357
0 18359 5 1 1 18358
0 18360 7 1 2 81632 73946
0 18361 7 1 2 92366 18360
0 18362 7 1 2 93707 18361
0 18363 5 1 1 18362
0 18364 7 1 2 18359 18363
0 18365 5 1 1 18364
0 18366 7 1 2 93704 18365
0 18367 5 1 1 18366
0 18368 7 2 2 74621 89388
0 18369 5 3 1 93718
0 18370 7 4 2 70317 78324
0 18371 7 1 2 73828 93723
0 18372 5 1 1 18371
0 18373 7 1 2 93720 18372
0 18374 5 1 1 18373
0 18375 7 1 2 70029 18374
0 18376 5 1 1 18375
0 18377 7 1 2 88434 18376
0 18378 5 1 1 18377
0 18379 7 1 2 84091 18378
0 18380 5 1 1 18379
0 18381 7 1 2 88851 83651
0 18382 7 1 2 91140 18381
0 18383 5 1 1 18382
0 18384 7 1 2 18380 18383
0 18385 5 1 1 18384
0 18386 7 1 2 66451 18385
0 18387 5 1 1 18386
0 18388 7 1 2 90105 86040
0 18389 7 1 2 93664 18388
0 18390 5 1 1 18389
0 18391 7 1 2 18387 18390
0 18392 5 1 1 18391
0 18393 7 1 2 93526 18392
0 18394 5 1 1 18393
0 18395 7 1 2 68968 91161
0 18396 5 1 1 18395
0 18397 7 1 2 16543 18396
0 18398 5 1 1 18397
0 18399 7 1 2 67670 18398
0 18400 5 1 1 18399
0 18401 7 4 2 88249 80114
0 18402 5 1 1 93727
0 18403 7 1 2 18400 18402
0 18404 5 1 1 18403
0 18405 7 11 2 64507 65392
0 18406 7 1 2 88804 93731
0 18407 7 1 2 92469 18406
0 18408 7 1 2 18404 18407
0 18409 5 1 1 18408
0 18410 7 1 2 18394 18409
0 18411 5 1 1 18410
0 18412 7 1 2 63302 18411
0 18413 5 1 1 18412
0 18414 7 1 2 18367 18413
0 18415 5 1 1 18414
0 18416 7 1 2 64337 18415
0 18417 5 1 1 18416
0 18418 7 2 2 70030 93517
0 18419 7 1 2 91738 93742
0 18420 7 1 2 93681 18419
0 18421 5 1 1 18420
0 18422 7 1 2 18417 18421
0 18423 5 1 1 18422
0 18424 7 1 2 71053 18423
0 18425 5 1 1 18424
0 18426 7 1 2 18346 18425
0 18427 5 1 1 18426
0 18428 7 1 2 73002 18427
0 18429 5 1 1 18428
0 18430 7 1 2 62058 18429
0 18431 7 1 2 18112 18430
0 18432 5 1 1 18431
0 18433 7 1 2 17190 18432
0 18434 5 1 1 18433
0 18435 7 1 2 16805 18434
0 18436 7 1 2 16640 18435
0 18437 5 1 1 18436
0 18438 7 1 2 69084 18437
0 18439 5 1 1 18438
0 18440 7 13 2 61348 67848
0 18441 5 1 1 93744
0 18442 7 8 2 66214 62999
0 18443 5 1 1 93757
0 18444 7 5 2 18441 18443
0 18445 5 74 1 93765
0 18446 7 4 2 66099 62951
0 18447 5 1 1 93844
0 18448 7 1 2 16966 18447
0 18449 5 42 1 18448
0 18450 7 36 2 64242 69181
0 18451 7 4 2 68381 72604
0 18452 5 2 1 93926
0 18453 7 3 2 62059 65720
0 18454 5 2 1 93932
0 18455 7 6 2 70674 72847
0 18456 7 1 2 62559 93937
0 18457 5 1 1 18456
0 18458 7 1 2 93935 18457
0 18459 5 2 1 18458
0 18460 7 1 2 77610 93943
0 18461 5 1 1 18460
0 18462 7 9 2 62060 70318
0 18463 7 1 2 85473 93945
0 18464 5 1 1 18463
0 18465 7 1 2 18461 18464
0 18466 5 1 1 18465
0 18467 7 1 2 63771 18466
0 18468 5 1 1 18467
0 18469 7 2 2 73620 82483
0 18470 5 1 1 93954
0 18471 7 1 2 18468 18470
0 18472 5 1 1 18471
0 18473 7 1 2 93927 18472
0 18474 5 1 1 18473
0 18475 7 2 2 72749 80446
0 18476 7 1 2 62061 77450
0 18477 7 1 2 93956 18476
0 18478 5 1 1 18477
0 18479 7 1 2 18474 18478
0 18480 5 1 1 18479
0 18481 7 1 2 62819 18480
0 18482 5 1 1 18481
0 18483 7 2 2 74452 76401
0 18484 5 1 1 93958
0 18485 7 1 2 79522 93959
0 18486 5 1 1 18485
0 18487 7 1 2 87919 93957
0 18488 5 1 1 18487
0 18489 7 1 2 71936 89801
0 18490 5 1 1 18489
0 18491 7 3 2 68616 72916
0 18492 7 5 2 65393 72605
0 18493 5 1 1 93963
0 18494 7 1 2 93960 93964
0 18495 5 1 1 18494
0 18496 7 1 2 65721 18495
0 18497 7 1 2 18490 18496
0 18498 5 1 1 18497
0 18499 7 2 2 68617 90319
0 18500 5 1 1 93968
0 18501 7 1 2 73426 80896
0 18502 5 2 1 18501
0 18503 7 1 2 18500 93970
0 18504 5 8 1 18503
0 18505 7 1 2 72782 93972
0 18506 5 1 1 18505
0 18507 7 2 2 68618 90356
0 18508 5 1 1 93980
0 18509 7 1 2 70675 18508
0 18510 7 1 2 18506 18509
0 18511 5 1 1 18510
0 18512 7 1 2 18498 18511
0 18513 5 1 1 18512
0 18514 7 2 2 65973 91422
0 18515 7 1 2 79653 93982
0 18516 5 1 1 18515
0 18517 7 1 2 62062 18516
0 18518 7 1 2 18513 18517
0 18519 5 1 1 18518
0 18520 7 1 2 71755 71613
0 18521 5 1 1 18520
0 18522 7 1 2 16344 18521
0 18523 5 1 1 18522
0 18524 7 1 2 63772 18523
0 18525 5 1 1 18524
0 18526 7 1 2 68619 85157
0 18527 5 3 1 18526
0 18528 7 1 2 18525 93984
0 18529 5 1 1 18528
0 18530 7 1 2 84355 18529
0 18531 5 1 1 18530
0 18532 7 2 2 71821 72535
0 18533 5 1 1 93987
0 18534 7 1 2 86502 93988
0 18535 5 1 1 18534
0 18536 7 1 2 66926 18535
0 18537 7 1 2 18531 18536
0 18538 5 1 1 18537
0 18539 7 1 2 18519 18538
0 18540 5 1 1 18539
0 18541 7 1 2 18488 18540
0 18542 5 1 1 18541
0 18543 7 1 2 63538 18542
0 18544 5 1 1 18543
0 18545 7 1 2 18486 18544
0 18546 7 1 2 18482 18545
0 18547 5 1 1 18546
0 18548 7 1 2 63303 18547
0 18549 5 1 1 18548
0 18550 7 3 2 77718 89719
0 18551 5 1 1 93989
0 18552 7 1 2 86895 93990
0 18553 5 1 1 18552
0 18554 7 2 2 63304 93973
0 18555 7 1 2 62820 93992
0 18556 5 1 1 18555
0 18557 7 1 2 18553 18556
0 18558 5 1 1 18557
0 18559 7 1 2 89200 80282
0 18560 7 1 2 18558 18559
0 18561 5 1 1 18560
0 18562 7 1 2 18549 18561
0 18563 5 1 1 18562
0 18564 7 1 2 66452 18563
0 18565 5 1 1 18564
0 18566 7 1 2 84356 73065
0 18567 5 1 1 18566
0 18568 7 1 2 89745 18567
0 18569 5 1 1 18568
0 18570 7 1 2 68620 18569
0 18571 5 1 1 18570
0 18572 7 1 2 86405 90372
0 18573 5 1 1 18572
0 18574 7 1 2 18571 18573
0 18575 5 1 1 18574
0 18576 7 1 2 67432 18575
0 18577 5 1 1 18576
0 18578 7 1 2 62821 74582
0 18579 7 1 2 77987 18578
0 18580 5 1 1 18579
0 18581 7 1 2 73661 18580
0 18582 5 1 1 18581
0 18583 7 1 2 67232 18582
0 18584 5 1 1 18583
0 18585 7 1 2 77902 93711
0 18586 5 1 1 18585
0 18587 7 1 2 18584 18586
0 18588 5 1 1 18587
0 18589 7 1 2 73427 18588
0 18590 5 1 1 18589
0 18591 7 1 2 74519 77278
0 18592 5 2 1 18591
0 18593 7 1 2 65394 75270
0 18594 7 1 2 93994 18593
0 18595 5 1 1 18594
0 18596 7 1 2 18590 18595
0 18597 7 1 2 18577 18596
0 18598 5 1 1 18597
0 18599 7 1 2 68382 18598
0 18600 5 1 1 18599
0 18601 7 1 2 89894 85806
0 18602 5 1 1 18601
0 18603 7 1 2 18600 18602
0 18604 5 1 1 18603
0 18605 7 1 2 66927 18604
0 18606 5 1 1 18605
0 18607 7 1 2 67233 84170
0 18608 5 1 1 18607
0 18609 7 1 2 74536 18608
0 18610 5 1 1 18609
0 18611 7 1 2 68822 85680
0 18612 7 2 2 18610 18611
0 18613 5 1 1 93996
0 18614 7 5 2 65722 71937
0 18615 5 1 1 93998
0 18616 7 2 2 68383 93999
0 18617 5 2 1 94003
0 18618 7 1 2 70319 94004
0 18619 5 1 1 18618
0 18620 7 1 2 18613 18619
0 18621 5 1 1 18620
0 18622 7 1 2 67433 18621
0 18623 5 1 1 18622
0 18624 7 1 2 75948 73206
0 18625 5 4 1 18624
0 18626 7 1 2 72490 94007
0 18627 5 2 1 18626
0 18628 7 2 2 71938 94011
0 18629 5 1 1 94013
0 18630 7 1 2 68384 94014
0 18631 5 1 1 18630
0 18632 7 1 2 18623 18631
0 18633 5 2 1 18632
0 18634 7 1 2 66928 94015
0 18635 5 1 1 18634
0 18636 7 5 2 75949 75031
0 18637 5 1 1 94017
0 18638 7 1 2 86523 94018
0 18639 5 1 1 18638
0 18640 7 1 2 18635 18639
0 18641 5 1 1 18640
0 18642 7 1 2 72126 18641
0 18643 5 1 1 18642
0 18644 7 1 2 74505 85613
0 18645 5 11 1 18644
0 18646 7 4 2 63944 76700
0 18647 5 1 1 94033
0 18648 7 1 2 80617 94034
0 18649 7 1 2 94022 18648
0 18650 5 1 1 18649
0 18651 7 1 2 18643 18650
0 18652 5 1 1 18651
0 18653 7 1 2 67671 18652
0 18654 5 1 1 18653
0 18655 7 1 2 79654 90135
0 18656 7 1 2 85802 18655
0 18657 5 1 1 18656
0 18658 7 1 2 18654 18657
0 18659 7 1 2 18606 18658
0 18660 5 1 1 18659
0 18661 7 1 2 81841 18660
0 18662 5 1 1 18661
0 18663 7 1 2 89333 93946
0 18664 5 1 1 18663
0 18665 7 3 2 73428 92435
0 18666 5 4 1 94037
0 18667 7 2 2 65395 71822
0 18668 7 1 2 85526 94044
0 18669 7 1 2 94040 18668
0 18670 5 1 1 18669
0 18671 7 1 2 18664 18670
0 18672 5 1 1 18671
0 18673 7 1 2 65723 18672
0 18674 5 1 1 18673
0 18675 7 1 2 86605 86503
0 18676 5 1 1 18675
0 18677 7 11 2 62063 67434
0 18678 7 1 2 72370 94046
0 18679 5 3 1 18678
0 18680 7 1 2 18676 94057
0 18681 5 1 1 18680
0 18682 7 1 2 63773 18681
0 18683 5 1 1 18682
0 18684 7 1 2 71228 91086
0 18685 5 1 1 18684
0 18686 7 1 2 94008 18685
0 18687 5 1 1 18686
0 18688 7 1 2 62064 18687
0 18689 5 1 1 18688
0 18690 7 1 2 18683 18689
0 18691 5 1 1 18690
0 18692 7 1 2 72127 18691
0 18693 5 1 1 18692
0 18694 7 1 2 18674 18693
0 18695 5 1 1 18694
0 18696 7 1 2 63539 18695
0 18697 5 1 1 18696
0 18698 7 2 2 89932 77147
0 18699 7 1 2 79238 80447
0 18700 5 1 1 18699
0 18701 7 1 2 72128 73753
0 18702 5 1 1 18701
0 18703 7 1 2 18700 18702
0 18704 5 1 1 18703
0 18705 7 1 2 94060 18704
0 18706 5 1 1 18705
0 18707 7 1 2 18697 18706
0 18708 5 1 1 18707
0 18709 7 1 2 63305 80932
0 18710 7 1 2 18708 18709
0 18711 5 1 1 18710
0 18712 7 1 2 18662 18711
0 18713 7 1 2 18565 18712
0 18714 5 1 1 18713
0 18715 7 1 2 63137 18714
0 18716 5 1 1 18715
0 18717 7 1 2 62394 90325
0 18718 5 2 1 18717
0 18719 7 1 2 93180 94062
0 18720 5 2 1 18719
0 18721 7 1 2 93654 94064
0 18722 5 1 1 18721
0 18723 7 1 2 62065 18722
0 18724 5 1 1 18723
0 18725 7 6 2 63945 78789
0 18726 7 1 2 74705 94066
0 18727 5 1 1 18726
0 18728 7 1 2 18724 18727
0 18729 5 1 1 18728
0 18730 7 1 2 68621 18729
0 18731 5 1 1 18730
0 18732 7 2 2 82195 84587
0 18733 5 1 1 94072
0 18734 7 1 2 62066 94073
0 18735 5 1 1 18734
0 18736 7 1 2 18731 18735
0 18737 5 1 1 18736
0 18738 7 1 2 70676 18737
0 18739 5 1 1 18738
0 18740 7 2 2 63540 76701
0 18741 7 1 2 82484 94074
0 18742 5 1 1 18741
0 18743 7 2 2 66929 77442
0 18744 7 2 2 73606 73754
0 18745 5 2 1 94078
0 18746 7 1 2 94076 94079
0 18747 5 1 1 18746
0 18748 7 1 2 70677 11283
0 18749 5 2 1 18748
0 18750 7 1 2 65724 77619
0 18751 5 1 1 18750
0 18752 7 1 2 75138 18751
0 18753 7 1 2 94082 18752
0 18754 5 1 1 18753
0 18755 7 1 2 18747 18754
0 18756 5 1 1 18755
0 18757 7 1 2 63774 18756
0 18758 5 1 1 18757
0 18759 7 1 2 18742 18758
0 18760 7 1 2 18739 18759
0 18761 5 1 1 18760
0 18762 7 1 2 84357 18761
0 18763 5 1 1 18762
0 18764 7 1 2 72371 74398
0 18765 5 3 1 18764
0 18766 7 1 2 62395 76221
0 18767 5 1 1 18766
0 18768 7 1 2 94084 18767
0 18769 5 1 1 18768
0 18770 7 1 2 62067 18769
0 18771 5 1 1 18770
0 18772 7 5 2 70678 77299
0 18773 7 1 2 86606 94087
0 18774 5 1 1 18773
0 18775 7 1 2 18771 18774
0 18776 5 1 1 18775
0 18777 7 1 2 63775 18776
0 18778 5 1 1 18777
0 18779 7 1 2 93503 94009
0 18780 5 1 1 18779
0 18781 7 1 2 75765 18780
0 18782 5 1 1 18781
0 18783 7 1 2 18778 18782
0 18784 5 1 1 18783
0 18785 7 1 2 89507 18784
0 18786 5 1 1 18785
0 18787 7 2 2 72047 94035
0 18788 7 2 2 62396 75222
0 18789 5 1 1 94094
0 18790 7 1 2 94047 94095
0 18791 7 1 2 94092 18790
0 18792 5 1 1 18791
0 18793 7 1 2 18786 18792
0 18794 7 1 2 18763 18793
0 18795 5 1 1 18794
0 18796 7 1 2 91143 18795
0 18797 5 1 1 18796
0 18798 7 1 2 18716 18797
0 18799 5 1 1 18798
0 18800 7 1 2 79800 18799
0 18801 5 1 1 18800
0 18802 7 3 2 68823 78001
0 18803 7 2 2 67435 94096
0 18804 5 2 1 94099
0 18805 7 1 2 72129 75743
0 18806 7 1 2 85604 18805
0 18807 5 1 1 18806
0 18808 7 2 2 94101 18807
0 18809 5 1 1 94103
0 18810 7 1 2 63776 94104
0 18811 5 1 1 18810
0 18812 7 2 2 63946 91242
0 18813 5 2 1 94105
0 18814 7 1 2 68622 94107
0 18815 5 1 1 18814
0 18816 7 1 2 65396 18815
0 18817 7 1 2 18811 18816
0 18818 5 1 1 18817
0 18819 7 2 2 77503 72825
0 18820 5 30 1 94109
0 18821 7 2 2 70679 93974
0 18822 5 1 1 94141
0 18823 7 3 2 76702 75321
0 18824 5 1 1 94143
0 18825 7 1 2 18822 18824
0 18826 5 4 1 18825
0 18827 7 1 2 94111 94146
0 18828 5 1 1 18827
0 18829 7 1 2 91087 85301
0 18830 5 1 1 18829
0 18831 7 1 2 18828 18830
0 18832 7 1 2 18818 18831
0 18833 5 1 1 18832
0 18834 7 1 2 88705 18833
0 18835 5 1 1 18834
0 18836 7 3 2 85123 80823
0 18837 7 2 2 88438 73607
0 18838 7 1 2 94150 94153
0 18839 7 1 2 12627 18838
0 18840 5 1 1 18839
0 18841 7 1 2 18835 18840
0 18842 5 1 1 18841
0 18843 7 1 2 61544 18842
0 18844 5 1 1 18843
0 18845 7 1 2 81764 94147
0 18846 5 1 1 18845
0 18847 7 3 2 73207 74568
0 18848 7 2 2 85124 78754
0 18849 7 1 2 94155 94158
0 18850 5 1 1 18849
0 18851 7 1 2 18846 18850
0 18852 5 1 1 18851
0 18853 7 1 2 94112 18852
0 18854 5 1 1 18853
0 18855 7 1 2 85819 73880
0 18856 5 2 1 18855
0 18857 7 1 2 65397 94160
0 18858 5 1 1 18857
0 18859 7 1 2 93504 18858
0 18860 5 1 1 18859
0 18861 7 1 2 67672 18860
0 18862 5 1 1 18861
0 18863 7 1 2 6858 18862
0 18864 5 1 1 18863
0 18865 7 1 2 72130 18864
0 18866 5 1 1 18865
0 18867 7 1 2 91423 94100
0 18868 5 1 1 18867
0 18869 7 1 2 85448 91088
0 18870 5 1 1 18869
0 18871 7 1 2 18629 18870
0 18872 5 1 1 18871
0 18873 7 1 2 72536 18872
0 18874 5 1 1 18873
0 18875 7 1 2 18868 18874
0 18876 7 1 2 18866 18875
0 18877 5 1 1 18876
0 18878 7 1 2 81765 18877
0 18879 5 1 1 18878
0 18880 7 1 2 18854 18879
0 18881 5 1 1 18880
0 18882 7 1 2 82113 18881
0 18883 5 1 1 18882
0 18884 7 1 2 18844 18883
0 18885 5 1 1 18884
0 18886 7 1 2 75766 18885
0 18887 5 1 1 18886
0 18888 7 1 2 89778 94113
0 18889 5 1 1 18888
0 18890 7 2 2 63947 89508
0 18891 7 2 2 62397 94162
0 18892 5 1 1 94164
0 18893 7 1 2 18889 18892
0 18894 5 1 1 18893
0 18895 7 1 2 70680 18894
0 18896 5 1 1 18895
0 18897 7 2 2 72606 84558
0 18898 5 1 1 94166
0 18899 7 1 2 93677 18898
0 18900 5 1 1 18899
0 18901 7 1 2 77852 18900
0 18902 5 1 1 18901
0 18903 7 1 2 18896 18902
0 18904 5 1 1 18903
0 18905 7 1 2 63777 18904
0 18906 5 1 1 18905
0 18907 7 2 2 75271 94114
0 18908 5 1 1 94168
0 18909 7 1 2 77627 94169
0 18910 5 1 1 18909
0 18911 7 1 2 18906 18910
0 18912 5 1 1 18911
0 18913 7 1 2 68148 18912
0 18914 5 1 1 18913
0 18915 7 3 2 82136 85029
0 18916 7 1 2 18809 94170
0 18917 5 1 1 18916
0 18918 7 1 2 18914 18917
0 18919 5 1 1 18918
0 18920 7 1 2 68385 18919
0 18921 5 1 1 18920
0 18922 7 1 2 72697 88795
0 18923 7 1 2 94093 18922
0 18924 5 1 1 18923
0 18925 7 1 2 62068 18924
0 18926 7 1 2 18921 18925
0 18927 5 1 1 18926
0 18928 7 1 2 76224 85627
0 18929 5 1 1 18928
0 18930 7 1 2 72131 18929
0 18931 5 1 1 18930
0 18932 7 1 2 91291 76614
0 18933 5 1 1 18932
0 18934 7 1 2 18931 18933
0 18935 5 1 1 18934
0 18936 7 1 2 67673 18935
0 18937 5 1 1 18936
0 18938 7 2 2 72537 76366
0 18939 5 1 1 94173
0 18940 7 1 2 77575 94174
0 18941 5 1 1 18940
0 18942 7 1 2 73758 1906
0 18943 5 1 1 18942
0 18944 7 1 2 93995 18943
0 18945 5 1 1 18944
0 18946 7 1 2 18941 18945
0 18947 7 1 2 18937 18946
0 18948 5 1 1 18947
0 18949 7 1 2 65398 18948
0 18950 5 1 1 18949
0 18951 7 1 2 75916 85299
0 18952 5 1 1 18951
0 18953 7 1 2 18950 18952
0 18954 5 1 1 18953
0 18955 7 1 2 68623 18954
0 18956 5 1 1 18955
0 18957 7 1 2 75512 72372
0 18958 5 2 1 18957
0 18959 7 2 2 15649 94175
0 18960 5 1 1 94177
0 18961 7 1 2 89509 18960
0 18962 5 1 1 18961
0 18963 7 1 2 85530 86639
0 18964 5 1 1 18963
0 18965 7 1 2 18962 18964
0 18966 5 1 1 18965
0 18967 7 1 2 68386 18966
0 18968 5 1 1 18967
0 18969 7 1 2 18956 18968
0 18970 5 1 1 18969
0 18971 7 1 2 63306 18970
0 18972 5 1 1 18971
0 18973 7 1 2 71727 86647
0 18974 5 1 1 18973
0 18975 7 1 2 82503 18974
0 18976 5 1 1 18975
0 18977 7 1 2 77611 18976
0 18978 5 1 1 18977
0 18979 7 1 2 85474 74706
0 18980 5 2 1 18979
0 18981 7 1 2 18978 94179
0 18982 5 1 1 18981
0 18983 7 1 2 63778 18982
0 18984 5 1 1 18983
0 18985 7 1 2 74885 85158
0 18986 5 2 1 18985
0 18987 7 1 2 18984 94181
0 18988 5 1 1 18987
0 18989 7 1 2 68149 18988
0 18990 5 1 1 18989
0 18991 7 1 2 83411 94142
0 18992 5 1 1 18991
0 18993 7 1 2 18990 18992
0 18994 5 1 1 18993
0 18995 7 1 2 84358 18994
0 18996 5 1 1 18995
0 18997 7 4 2 74270 89720
0 18998 5 5 1 94183
0 18999 7 1 2 94106 94184
0 19000 5 1 1 18999
0 19001 7 1 2 66930 19000
0 19002 7 1 2 18996 19001
0 19003 7 1 2 18972 19002
0 19004 5 1 1 19003
0 19005 7 1 2 69355 76141
0 19006 7 1 2 19004 19005
0 19007 7 1 2 18927 19006
0 19008 5 1 1 19007
0 19009 7 1 2 18887 19008
0 19010 5 1 1 19009
0 19011 7 1 2 61836 19010
0 19012 5 1 1 19011
0 19013 7 1 2 18801 19012
0 19014 5 1 1 19013
0 19015 7 1 2 70031 19014
0 19016 5 1 1 19015
0 19017 7 2 2 71523 90373
0 19018 5 2 1 94192
0 19019 7 1 2 85542 91424
0 19020 5 1 1 19019
0 19021 7 1 2 94194 19020
0 19022 5 1 1 19021
0 19023 7 1 2 66931 19022
0 19024 5 1 1 19023
0 19025 7 3 2 90320 79477
0 19026 7 1 2 73807 94196
0 19027 5 1 1 19026
0 19028 7 1 2 19024 19027
0 19029 5 1 1 19028
0 19030 7 1 2 63541 19029
0 19031 5 1 1 19030
0 19032 7 1 2 11451 94058
0 19033 5 1 1 19032
0 19034 7 1 2 63779 19033
0 19035 5 1 1 19034
0 19036 7 1 2 85550 88015
0 19037 5 1 1 19036
0 19038 7 1 2 62069 91089
0 19039 7 1 2 19037 19038
0 19040 5 1 1 19039
0 19041 7 1 2 19035 19040
0 19042 5 1 1 19041
0 19043 7 1 2 68387 19042
0 19044 5 1 1 19043
0 19045 7 1 2 71823 88887
0 19046 5 1 1 19045
0 19047 7 1 2 66932 74897
0 19048 7 1 2 19046 19047
0 19049 5 1 1 19048
0 19050 7 1 2 62070 73925
0 19051 5 1 1 19050
0 19052 7 1 2 73119 19051
0 19053 7 1 2 19049 19052
0 19054 5 1 1 19053
0 19055 7 1 2 19044 19054
0 19056 7 1 2 19031 19055
0 19057 5 1 1 19056
0 19058 7 1 2 68969 19057
0 19059 5 1 1 19058
0 19060 7 1 2 75090 91442
0 19061 5 1 1 19060
0 19062 7 4 2 79992 91425
0 19063 7 1 2 63542 94199
0 19064 5 1 1 19063
0 19065 7 1 2 74054 78390
0 19066 5 15 1 19065
0 19067 7 1 2 73208 94203
0 19068 5 1 1 19067
0 19069 7 1 2 19064 19068
0 19070 5 1 1 19069
0 19071 7 1 2 66933 19070
0 19072 5 1 1 19071
0 19073 7 1 2 62071 94016
0 19074 5 2 1 19073
0 19075 7 1 2 19072 94218
0 19076 5 1 1 19075
0 19077 7 1 2 65974 19076
0 19078 5 1 1 19077
0 19079 7 1 2 19061 19078
0 19080 7 1 2 19059 19079
0 19081 5 1 1 19080
0 19082 7 1 2 61837 19081
0 19083 5 1 1 19082
0 19084 7 1 2 63543 11171
0 19085 5 2 1 19084
0 19086 7 1 2 65725 75412
0 19087 7 1 2 94220 19086
0 19088 5 1 1 19087
0 19089 7 1 2 66694 74433
0 19090 7 1 2 80380 19089
0 19091 5 1 1 19090
0 19092 7 1 2 19088 19091
0 19093 5 1 1 19092
0 19094 7 1 2 62560 19093
0 19095 5 1 1 19094
0 19096 7 1 2 75496 77357
0 19097 5 1 1 19096
0 19098 7 1 2 19095 19097
0 19099 5 1 1 19098
0 19100 7 1 2 62398 19099
0 19101 5 1 1 19100
0 19102 7 1 2 79773 803
0 19103 7 1 2 86852 19102
0 19104 5 1 1 19103
0 19105 7 1 2 19101 19104
0 19106 5 1 1 19105
0 19107 7 1 2 63780 19106
0 19108 5 1 1 19107
0 19109 7 1 2 63544 623
0 19110 5 3 1 19109
0 19111 7 1 2 86549 94222
0 19112 5 1 1 19111
0 19113 7 1 2 94065 19112
0 19114 5 1 1 19113
0 19115 7 1 2 68624 19114
0 19116 5 2 1 19115
0 19117 7 1 2 18733 94225
0 19118 5 1 1 19117
0 19119 7 1 2 70681 19118
0 19120 5 1 1 19119
0 19121 7 2 2 73714 76703
0 19122 7 1 2 68625 94227
0 19123 5 2 1 19122
0 19124 7 1 2 19120 94229
0 19125 5 1 1 19124
0 19126 7 1 2 75413 19125
0 19127 5 1 1 19126
0 19128 7 1 2 19108 19127
0 19129 5 1 1 19128
0 19130 7 1 2 72048 19129
0 19131 5 1 1 19130
0 19132 7 1 2 63545 80390
0 19133 5 1 1 19132
0 19134 7 1 2 2769 19133
0 19135 5 1 1 19134
0 19136 7 9 2 66695 68970
0 19137 7 1 2 92345 94231
0 19138 7 1 2 19135 19137
0 19139 5 1 1 19138
0 19140 7 1 2 19131 19139
0 19141 7 1 2 19083 19140
0 19142 5 1 1 19141
0 19143 7 1 2 76081 19142
0 19144 5 1 1 19143
0 19145 7 2 2 76381 91426
0 19146 5 1 1 94240
0 19147 7 1 2 66934 94241
0 19148 5 1 1 19147
0 19149 7 1 2 94219 19148
0 19150 5 1 1 19149
0 19151 7 1 2 72132 19150
0 19152 5 1 1 19151
0 19153 7 1 2 78025 84011
0 19154 5 3 1 19153
0 19155 7 1 2 67436 78212
0 19156 5 1 1 19155
0 19157 7 1 2 94242 19156
0 19158 5 2 1 19157
0 19159 7 1 2 77767 94245
0 19160 5 1 1 19159
0 19161 7 1 2 74656 93678
0 19162 5 1 1 19161
0 19163 7 1 2 19160 19162
0 19164 5 1 1 19163
0 19165 7 1 2 68824 19164
0 19166 5 1 1 19165
0 19167 7 1 2 79886 78298
0 19168 5 1 1 19167
0 19169 7 1 2 74399 87473
0 19170 5 1 1 19169
0 19171 7 1 2 19168 19170
0 19172 7 1 2 19166 19171
0 19173 5 1 1 19172
0 19174 7 1 2 63781 19173
0 19175 5 1 1 19174
0 19176 7 1 2 86734 91090
0 19177 5 1 1 19176
0 19178 7 3 2 65399 75322
0 19179 7 1 2 72049 94247
0 19180 5 2 1 19179
0 19181 7 1 2 19177 94250
0 19182 5 1 1 19181
0 19183 7 1 2 63546 19182
0 19184 5 1 1 19183
0 19185 7 1 2 76367 91091
0 19186 7 1 2 93679 19185
0 19187 5 1 1 19186
0 19188 7 1 2 65726 19187
0 19189 7 1 2 19184 19188
0 19190 7 1 2 19175 19189
0 19191 5 1 1 19190
0 19192 7 2 2 73429 85062
0 19193 5 1 1 94252
0 19194 7 1 2 614 19193
0 19195 5 1 1 19194
0 19196 7 1 2 85690 19195
0 19197 5 1 1 19196
0 19198 7 1 2 94226 19197
0 19199 5 2 1 19198
0 19200 7 1 2 72050 94254
0 19201 5 1 1 19200
0 19202 7 1 2 72133 94204
0 19203 5 1 1 19202
0 19204 7 4 2 62399 72698
0 19205 7 2 2 75182 94256
0 19206 5 1 1 94260
0 19207 7 1 2 74622 94261
0 19208 5 1 1 19207
0 19209 7 1 2 19203 19208
0 19210 5 1 1 19209
0 19211 7 1 2 63948 19210
0 19212 5 1 1 19211
0 19213 7 1 2 70682 19212
0 19214 7 1 2 19201 19213
0 19215 5 1 1 19214
0 19216 7 1 2 66935 19215
0 19217 7 1 2 19191 19216
0 19218 5 1 1 19217
0 19219 7 1 2 19152 19218
0 19220 5 1 1 19219
0 19221 7 1 2 67991 83289
0 19222 7 1 2 19220 19221
0 19223 5 1 1 19222
0 19224 7 1 2 19144 19223
0 19225 5 1 1 19224
0 19226 7 1 2 63307 19225
0 19227 5 1 1 19226
0 19228 7 2 2 85709 71016
0 19229 5 1 1 94262
0 19230 7 1 2 91062 94263
0 19231 5 2 1 19230
0 19232 7 2 2 65400 86216
0 19233 5 1 1 94266
0 19234 7 4 2 85369 86667
0 19235 5 1 1 94268
0 19236 7 1 2 68825 94269
0 19237 5 1 1 19236
0 19238 7 7 2 65401 78002
0 19239 5 1 1 94272
0 19240 7 1 2 78363 94273
0 19241 5 2 1 19240
0 19242 7 1 2 19237 94279
0 19243 5 1 1 19242
0 19244 7 1 2 67437 19243
0 19245 5 1 1 19244
0 19246 7 1 2 19233 19245
0 19247 5 1 1 19246
0 19248 7 1 2 68626 19247
0 19249 5 1 1 19248
0 19250 7 1 2 76341 93537
0 19251 5 1 1 19250
0 19252 7 1 2 19249 19251
0 19253 5 1 1 19252
0 19254 7 1 2 67234 19253
0 19255 5 1 1 19254
0 19256 7 1 2 94264 19255
0 19257 5 2 1 19256
0 19258 7 3 2 75572 80627
0 19259 7 1 2 94281 94283
0 19260 5 1 1 19259
0 19261 7 1 2 72051 93944
0 19262 5 1 1 19261
0 19263 7 1 2 62072 84932
0 19264 5 1 1 19263
0 19265 7 1 2 19262 19264
0 19266 5 1 1 19265
0 19267 7 1 2 88436 77300
0 19268 7 1 2 19266 19267
0 19269 5 1 1 19268
0 19270 7 1 2 19260 19269
0 19271 5 1 1 19270
0 19272 7 1 2 83046 19271
0 19273 5 1 1 19272
0 19274 7 1 2 19227 19273
0 19275 5 1 1 19274
0 19276 7 1 2 87468 19275
0 19277 5 1 1 19276
0 19278 7 1 2 19016 19277
0 19279 5 1 1 19278
0 19280 7 1 2 69547 19279
0 19281 5 1 1 19280
0 19282 7 4 2 65727 79904
0 19283 5 2 1 94286
0 19284 7 1 2 63782 94083
0 19285 7 1 2 94290 19284
0 19286 5 1 1 19285
0 19287 7 1 2 93985 19286
0 19288 5 3 1 19287
0 19289 7 1 2 72052 94292
0 19290 5 1 1 19289
0 19291 7 1 2 71824 77858
0 19292 5 1 1 19291
0 19293 7 1 2 19290 19292
0 19294 5 1 1 19293
0 19295 7 1 2 83108 19294
0 19296 5 1 1 19295
0 19297 7 1 2 77982 18162
0 19298 5 1 1 19297
0 19299 7 1 2 79510 19298
0 19300 5 3 1 19299
0 19301 7 1 2 94171 94295
0 19302 5 1 1 19301
0 19303 7 1 2 88796 72431
0 19304 5 1 1 19303
0 19305 7 1 2 19302 19304
0 19306 5 1 1 19305
0 19307 7 1 2 61838 19306
0 19308 5 1 1 19307
0 19309 7 1 2 19296 19308
0 19310 5 1 1 19309
0 19311 7 2 2 61545 80740
0 19312 7 1 2 19310 94298
0 19313 5 1 1 19312
0 19314 7 3 2 63783 78310
0 19315 5 1 1 94300
0 19316 7 1 2 78173 19315
0 19317 5 1 1 19316
0 19318 7 1 2 73430 19317
0 19319 5 1 1 19318
0 19320 7 1 2 73890 81169
0 19321 5 2 1 19320
0 19322 7 1 2 67438 94303
0 19323 5 1 1 19322
0 19324 7 1 2 68627 79729
0 19325 5 1 1 19324
0 19326 7 1 2 72134 94161
0 19327 5 1 1 19326
0 19328 7 1 2 19325 19327
0 19329 7 1 2 19323 19328
0 19330 7 1 2 19319 19329
0 19331 5 2 1 19330
0 19332 7 1 2 83047 94305
0 19333 5 1 1 19332
0 19334 7 1 2 5833 85258
0 19335 5 1 1 19334
0 19336 7 1 2 65728 75332
0 19337 5 2 1 19336
0 19338 7 1 2 72053 94307
0 19339 7 1 2 19335 19338
0 19340 5 1 1 19339
0 19341 7 1 2 75513 93557
0 19342 5 1 1 19341
0 19343 7 1 2 72283 79495
0 19344 5 2 1 19343
0 19345 7 1 2 73684 94309
0 19346 5 1 1 19345
0 19347 7 1 2 19342 19346
0 19348 7 1 2 19340 19347
0 19349 5 1 1 19348
0 19350 7 1 2 81446 19349
0 19351 5 1 1 19350
0 19352 7 1 2 19333 19351
0 19353 5 1 1 19352
0 19354 7 1 2 65402 19353
0 19355 5 1 1 19354
0 19356 7 1 2 86151 87056
0 19357 5 1 1 19356
0 19358 7 1 2 67439 89392
0 19359 7 1 2 93558 19358
0 19360 5 1 1 19359
0 19361 7 1 2 19357 19360
0 19362 5 1 1 19361
0 19363 7 1 2 70320 19362
0 19364 5 1 1 19363
0 19365 7 1 2 83109 77886
0 19366 5 1 1 19365
0 19367 7 1 2 19364 19366
0 19368 7 1 2 19355 19367
0 19369 5 1 1 19368
0 19370 7 1 2 77235 19369
0 19371 5 1 1 19370
0 19372 7 3 2 62561 89495
0 19373 5 1 1 94311
0 19374 7 1 2 80391 94312
0 19375 7 1 2 91304 19374
0 19376 5 1 1 19375
0 19377 7 1 2 19371 19376
0 19378 5 1 1 19377
0 19379 7 1 2 63547 19378
0 19380 5 1 1 19379
0 19381 7 1 2 19313 19380
0 19382 5 1 1 19381
0 19383 7 1 2 77375 19382
0 19384 5 1 1 19383
0 19385 7 2 2 71939 94296
0 19386 7 1 2 75414 94314
0 19387 5 1 1 19386
0 19388 7 1 2 75239 83019
0 19389 7 1 2 93541 19388
0 19390 5 1 1 19389
0 19391 7 1 2 19387 19390
0 19392 5 1 1 19391
0 19393 7 1 2 70321 19392
0 19394 5 1 1 19393
0 19395 7 1 2 65403 94306
0 19396 5 1 1 19395
0 19397 7 1 2 77888 19396
0 19398 5 1 1 19397
0 19399 7 1 2 75415 19398
0 19400 5 1 1 19399
0 19401 7 1 2 19394 19400
0 19402 5 1 1 19401
0 19403 7 1 2 63548 19402
0 19404 5 1 1 19403
0 19405 7 2 2 77853 84614
0 19406 5 1 1 94316
0 19407 7 1 2 94221 94317
0 19408 5 2 1 19407
0 19409 7 6 2 63949 75323
0 19410 7 1 2 94223 94320
0 19411 5 1 1 19410
0 19412 7 1 2 74034 84581
0 19413 5 1 1 19412
0 19414 7 1 2 19411 19413
0 19415 5 1 1 19414
0 19416 7 1 2 71728 19415
0 19417 5 1 1 19416
0 19418 7 1 2 94318 19417
0 19419 5 1 1 19418
0 19420 7 1 2 72054 19419
0 19421 5 1 1 19420
0 19422 7 1 2 75528 76228
0 19423 5 2 1 19422
0 19424 7 1 2 76225 94326
0 19425 5 1 1 19424
0 19426 7 1 2 68971 19425
0 19427 5 1 1 19426
0 19428 7 1 2 68388 77859
0 19429 5 1 1 19428
0 19430 7 1 2 19427 19429
0 19431 5 1 1 19430
0 19432 7 1 2 71825 19431
0 19433 5 1 1 19432
0 19434 7 1 2 19421 19433
0 19435 5 1 1 19434
0 19436 7 1 2 75416 19435
0 19437 5 1 1 19436
0 19438 7 1 2 19404 19437
0 19439 5 1 1 19438
0 19440 7 1 2 63308 19439
0 19441 5 1 1 19440
0 19442 7 1 2 73897 85099
0 19443 7 2 2 89841 19442
0 19444 7 1 2 86594 94328
0 19445 5 1 1 19444
0 19446 7 1 2 65125 19445
0 19447 7 1 2 19441 19446
0 19448 5 1 1 19447
0 19449 7 1 2 72248 73861
0 19450 5 1 1 19449
0 19451 7 1 2 548 19450
0 19452 5 1 1 19451
0 19453 7 1 2 77976 19452
0 19454 5 1 1 19453
0 19455 7 2 2 73431 78003
0 19456 5 1 1 94330
0 19457 7 1 2 76355 19456
0 19458 5 2 1 19457
0 19459 7 1 2 79774 74922
0 19460 7 1 2 94332 19459
0 19461 5 1 1 19460
0 19462 7 1 2 19454 19461
0 19463 5 1 1 19462
0 19464 7 1 2 66936 19463
0 19465 5 1 1 19464
0 19466 7 1 2 71778 72323
0 19467 7 1 2 88752 19466
0 19468 7 1 2 80448 19467
0 19469 5 1 1 19468
0 19470 7 1 2 19465 19469
0 19471 5 1 1 19470
0 19472 7 1 2 63784 19471
0 19473 5 1 1 19472
0 19474 7 1 2 74863 71524
0 19475 5 1 1 19474
0 19476 7 1 2 76464 19475
0 19477 5 1 1 19476
0 19478 7 1 2 72538 19477
0 19479 5 1 1 19478
0 19480 7 1 2 94005 19479
0 19481 5 1 1 19480
0 19482 7 1 2 70322 19481
0 19483 5 1 1 19482
0 19484 7 7 2 70683 84683
0 19485 7 1 2 72324 84962
0 19486 5 1 1 19485
0 19487 7 1 2 67235 93981
0 19488 5 1 1 19487
0 19489 7 1 2 19486 19488
0 19490 5 1 1 19489
0 19491 7 1 2 94334 19490
0 19492 5 1 1 19491
0 19493 7 1 2 19483 19492
0 19494 5 1 1 19493
0 19495 7 1 2 67440 19494
0 19496 5 1 1 19495
0 19497 7 4 2 70323 73256
0 19498 7 1 2 85579 94341
0 19499 5 2 1 19498
0 19500 7 1 2 84035 94345
0 19501 5 1 1 19500
0 19502 7 1 2 71940 19501
0 19503 5 1 1 19502
0 19504 7 1 2 75344 75210
0 19505 5 1 1 19504
0 19506 7 1 2 19503 19505
0 19507 5 1 1 19506
0 19508 7 1 2 68389 19507
0 19509 5 1 1 19508
0 19510 7 2 2 78290 93675
0 19511 5 1 1 94347
0 19512 7 1 2 74800 94348
0 19513 5 1 1 19512
0 19514 7 1 2 19509 19513
0 19515 7 1 2 19496 19514
0 19516 5 1 1 19515
0 19517 7 1 2 75887 19516
0 19518 5 1 1 19517
0 19519 7 1 2 19473 19518
0 19520 5 1 1 19519
0 19521 7 1 2 63309 19520
0 19522 5 1 1 19521
0 19523 7 1 2 88908 94329
0 19524 5 1 1 19523
0 19525 7 1 2 70032 19524
0 19526 7 1 2 19522 19525
0 19527 5 1 1 19526
0 19528 7 1 2 77236 19527
0 19529 7 1 2 19448 19528
0 19530 5 1 1 19529
0 19531 7 1 2 19384 19530
0 19532 5 1 1 19531
0 19533 7 1 2 79443 19532
0 19534 5 1 1 19533
0 19535 7 1 2 19281 19534
0 19536 5 1 1 19535
0 19537 7 1 2 93890 19536
0 19538 5 1 1 19537
0 19539 7 44 2 69085 64338
0 19540 7 17 2 64508 94349
0 19541 7 1 2 72410 91275
0 19542 5 2 1 19541
0 19543 7 1 2 65404 84921
0 19544 5 1 1 19543
0 19545 7 1 2 94410 19544
0 19546 5 1 1 19545
0 19547 7 1 2 67236 19546
0 19548 5 1 1 19547
0 19549 7 1 2 72783 94036
0 19550 5 1 1 19549
0 19551 7 1 2 19548 19550
0 19552 5 1 1 19551
0 19553 7 1 2 90189 19552
0 19554 5 1 1 19553
0 19555 7 2 2 78026 72343
0 19556 5 1 1 94412
0 19557 7 1 2 94108 19556
0 19558 5 1 1 19557
0 19559 7 1 2 65405 85323
0 19560 7 1 2 19558 19559
0 19561 5 1 1 19560
0 19562 7 1 2 19554 19561
0 19563 5 1 1 19562
0 19564 7 1 2 68628 19563
0 19565 5 1 1 19564
0 19566 7 1 2 89510 93341
0 19567 5 1 1 19566
0 19568 7 1 2 79511 19567
0 19569 5 1 1 19568
0 19570 7 1 2 73987 85324
0 19571 7 1 2 19569 19570
0 19572 5 1 1 19571
0 19573 7 1 2 19565 19572
0 19574 5 1 1 19573
0 19575 7 1 2 65126 19574
0 19576 5 1 1 19575
0 19577 7 1 2 71634 75015
0 19578 5 1 1 19577
0 19579 7 5 2 72539 72715
0 19580 5 3 1 94414
0 19581 7 1 2 71826 94415
0 19582 5 1 1 19581
0 19583 7 1 2 19578 19582
0 19584 5 1 1 19583
0 19585 7 1 2 63950 19584
0 19586 5 1 1 19585
0 19587 7 1 2 73647 77104
0 19588 5 1 1 19587
0 19589 7 1 2 19586 19588
0 19590 5 1 1 19589
0 19591 7 1 2 70684 19590
0 19592 5 1 1 19591
0 19593 7 1 2 73432 887
0 19594 5 3 1 19593
0 19595 7 1 2 64109 94422
0 19596 5 1 1 19595
0 19597 7 1 2 92409 19596
0 19598 5 1 1 19597
0 19599 7 1 2 88395 19598
0 19600 5 1 1 19599
0 19601 7 1 2 19592 19600
0 19602 5 1 1 19601
0 19603 7 1 2 83110 19602
0 19604 5 1 1 19603
0 19605 7 1 2 89466 83716
0 19606 5 1 1 19605
0 19607 7 1 2 94102 19606
0 19608 5 1 1 19607
0 19609 7 2 2 75950 19608
0 19610 7 1 2 88656 94425
0 19611 5 1 1 19610
0 19612 7 1 2 19604 19611
0 19613 5 1 1 19612
0 19614 7 1 2 90759 19613
0 19615 5 1 1 19614
0 19616 7 1 2 19576 19615
0 19617 5 1 1 19616
0 19618 7 1 2 68390 19617
0 19619 5 1 1 19618
0 19620 7 3 2 70324 79905
0 19621 5 1 1 94427
0 19622 7 5 2 62562 74488
0 19623 5 4 1 94430
0 19624 7 1 2 19621 94435
0 19625 5 1 1 19624
0 19626 7 1 2 72607 19625
0 19627 5 1 1 19626
0 19628 7 1 2 86793 76274
0 19629 5 1 1 19628
0 19630 7 1 2 19627 19629
0 19631 5 2 1 19630
0 19632 7 1 2 65729 94439
0 19633 5 1 1 19632
0 19634 7 2 2 63951 72716
0 19635 5 1 1 94441
0 19636 7 2 2 85030 19635
0 19637 5 1 1 94443
0 19638 7 1 2 83740 72288
0 19639 7 1 2 19637 19638
0 19640 5 1 1 19639
0 19641 7 1 2 19633 19640
0 19642 5 1 1 19641
0 19643 7 1 2 68629 19642
0 19644 5 1 1 19643
0 19645 7 3 2 65730 72608
0 19646 5 1 1 94445
0 19647 7 1 2 72300 19646
0 19648 5 6 1 19647
0 19649 7 1 2 89788 94448
0 19650 5 1 1 19649
0 19651 7 1 2 19644 19650
0 19652 5 1 1 19651
0 19653 7 1 2 70033 19652
0 19654 5 1 1 19653
0 19655 7 1 2 84396 77612
0 19656 5 1 1 19655
0 19657 7 5 2 70034 74623
0 19658 7 1 2 84257 94454
0 19659 5 1 1 19658
0 19660 7 1 2 70685 19659
0 19661 7 1 2 19656 19660
0 19662 5 1 1 19661
0 19663 7 2 2 72609 79906
0 19664 5 1 1 94459
0 19665 7 1 2 76889 94460
0 19666 5 1 1 19665
0 19667 7 1 2 79887 93533
0 19668 5 1 1 19667
0 19669 7 1 2 65731 19668
0 19670 7 1 2 19666 19669
0 19671 5 1 1 19670
0 19672 7 1 2 63785 19671
0 19673 7 1 2 19662 19672
0 19674 5 1 1 19673
0 19675 7 1 2 19654 19674
0 19676 5 1 1 19675
0 19677 7 1 2 68150 19676
0 19678 5 1 1 19677
0 19679 7 2 2 80858 86370
0 19680 7 1 2 94172 94461
0 19681 5 1 1 19680
0 19682 7 1 2 19678 19681
0 19683 5 1 1 19682
0 19684 7 1 2 61839 19683
0 19685 5 1 1 19684
0 19686 7 1 2 86568 85943
0 19687 5 1 1 19686
0 19688 7 1 2 85185 77600
0 19689 7 1 2 79814 19688
0 19690 5 1 1 19689
0 19691 7 1 2 19687 19690
0 19692 5 1 1 19691
0 19693 7 1 2 62400 19692
0 19694 5 1 1 19693
0 19695 7 1 2 71229 90374
0 19696 5 7 1 19695
0 19697 7 1 2 72717 74489
0 19698 5 1 1 19697
0 19699 7 1 2 72896 19698
0 19700 5 1 1 19699
0 19701 7 1 2 68630 19700
0 19702 5 1 1 19701
0 19703 7 1 2 94463 19702
0 19704 5 1 1 19703
0 19705 7 1 2 85225 19704
0 19706 5 1 1 19705
0 19707 7 1 2 19694 19706
0 19708 5 1 1 19707
0 19709 7 1 2 70686 19708
0 19710 5 1 1 19709
0 19711 7 1 2 68631 94440
0 19712 5 1 1 19711
0 19713 7 1 2 67237 75977
0 19714 7 1 2 83741 19713
0 19715 5 2 1 19714
0 19716 7 1 2 94176 94470
0 19717 5 4 1 19716
0 19718 7 1 2 72610 94472
0 19719 5 1 1 19718
0 19720 7 1 2 19712 19719
0 19721 5 1 1 19720
0 19722 7 1 2 82863 19721
0 19723 5 1 1 19722
0 19724 7 1 2 19710 19723
0 19725 5 1 1 19724
0 19726 7 1 2 82467 19725
0 19727 5 1 1 19726
0 19728 7 1 2 19685 19727
0 19729 5 1 1 19728
0 19730 7 1 2 77169 19729
0 19731 5 1 1 19730
0 19732 7 1 2 19619 19731
0 19733 5 1 1 19732
0 19734 7 1 2 66453 19733
0 19735 5 1 1 19734
0 19736 7 2 2 77490 93289
0 19737 5 2 1 94476
0 19738 7 3 2 65127 78509
0 19739 7 1 2 87542 94480
0 19740 7 1 2 94477 19739
0 19741 5 1 1 19740
0 19742 7 1 2 62073 19741
0 19743 7 1 2 19735 19742
0 19744 5 1 1 19743
0 19745 7 1 2 80706 87965
0 19746 5 1 1 19745
0 19747 7 1 2 68391 86278
0 19748 5 1 1 19747
0 19749 7 1 2 19746 19748
0 19750 5 1 1 19749
0 19751 7 1 2 67238 19750
0 19752 5 1 1 19751
0 19753 7 2 2 71318 93420
0 19754 5 1 1 94483
0 19755 7 1 2 76704 94484
0 19756 5 1 1 19755
0 19757 7 1 2 19752 19756
0 19758 5 1 1 19757
0 19759 7 1 2 68632 19758
0 19760 5 1 1 19759
0 19761 7 2 2 72344 77919
0 19762 7 1 2 74049 94485
0 19763 5 1 1 19762
0 19764 7 1 2 19760 19763
0 19765 5 1 1 19764
0 19766 7 1 2 63310 19765
0 19767 5 1 1 19766
0 19768 7 1 2 68826 73575
0 19769 5 3 1 19768
0 19770 7 1 2 78192 94487
0 19771 5 1 1 19770
0 19772 7 2 2 65128 73550
0 19773 7 1 2 73621 94490
0 19774 5 1 1 19773
0 19775 7 1 2 19771 19774
0 19776 5 1 1 19775
0 19777 7 1 2 62563 19776
0 19778 5 1 1 19777
0 19779 7 1 2 88756 87989
0 19780 5 1 1 19779
0 19781 7 1 2 19778 19780
0 19782 5 1 1 19781
0 19783 7 1 2 94185 19782
0 19784 5 1 1 19783
0 19785 7 1 2 19767 19784
0 19786 5 1 1 19785
0 19787 7 1 2 64110 19786
0 19788 5 1 1 19787
0 19789 7 1 2 79907 89511
0 19790 5 2 1 19789
0 19791 7 1 2 79512 94492
0 19792 5 1 1 19791
0 19793 7 1 2 65406 81300
0 19794 7 1 2 19792 19793
0 19795 5 1 1 19794
0 19796 7 1 2 62564 84869
0 19797 5 1 1 19796
0 19798 7 3 2 62822 72540
0 19799 5 5 1 94494
0 19800 7 1 2 70687 94495
0 19801 5 1 1 19800
0 19802 7 1 2 19797 19801
0 19803 5 1 1 19802
0 19804 7 1 2 83546 77613
0 19805 7 1 2 19803 19804
0 19806 5 1 1 19805
0 19807 7 1 2 19795 19806
0 19808 5 1 1 19807
0 19809 7 1 2 63786 19808
0 19810 5 1 1 19809
0 19811 7 1 2 82137 80754
0 19812 7 1 2 88320 19811
0 19813 5 1 1 19812
0 19814 7 1 2 19810 19813
0 19815 5 1 1 19814
0 19816 7 1 2 63549 19815
0 19817 5 1 1 19816
0 19818 7 4 2 68392 80755
0 19819 7 1 2 85135 94502
0 19820 7 1 2 91243 19819
0 19821 5 1 1 19820
0 19822 7 1 2 19817 19821
0 19823 7 1 2 19788 19822
0 19824 5 1 1 19823
0 19825 7 1 2 61840 19824
0 19826 5 1 1 19825
0 19827 7 4 2 62823 86695
0 19828 5 2 1 94506
0 19829 7 1 2 62565 94449
0 19830 5 1 1 19829
0 19831 7 1 2 94510 19830
0 19832 5 1 1 19831
0 19833 7 1 2 70035 19832
0 19834 5 1 1 19833
0 19835 7 2 2 74180 79555
0 19836 7 1 2 78027 94512
0 19837 5 1 1 19836
0 19838 7 1 2 19834 19837
0 19839 5 1 1 19838
0 19840 7 1 2 63952 19839
0 19841 5 1 1 19840
0 19842 7 1 2 84450 94413
0 19843 5 1 1 19842
0 19844 7 1 2 19841 19843
0 19845 5 1 1 19844
0 19846 7 1 2 71779 82920
0 19847 7 1 2 19845 19846
0 19848 5 1 1 19847
0 19849 7 1 2 19826 19848
0 19850 5 1 1 19849
0 19851 7 1 2 66454 19850
0 19852 5 1 1 19851
0 19853 7 2 2 89302 83370
0 19854 5 3 1 94514
0 19855 7 1 2 84318 94515
0 19856 5 4 1 19855
0 19857 7 2 2 70688 94519
0 19858 7 1 2 82468 94523
0 19859 5 1 1 19858
0 19860 7 2 2 89471 77988
0 19861 5 8 1 94525
0 19862 7 1 2 92154 94527
0 19863 5 1 1 19862
0 19864 7 1 2 19859 19863
0 19865 5 1 1 19864
0 19866 7 3 2 86761 82422
0 19867 5 1 1 94535
0 19868 7 1 2 84163 94536
0 19869 7 1 2 19865 19868
0 19870 5 1 1 19869
0 19871 7 1 2 19852 19870
0 19872 5 1 1 19871
0 19873 7 1 2 67992 19872
0 19874 5 1 1 19873
0 19875 7 1 2 68633 94442
0 19876 5 1 1 19875
0 19877 7 1 2 85820 19876
0 19878 5 1 1 19877
0 19879 7 1 2 76890 19878
0 19880 5 1 1 19879
0 19881 7 1 2 76981 19880
0 19882 5 1 1 19881
0 19883 7 1 2 72541 19882
0 19884 5 1 1 19883
0 19885 7 3 2 76574 77944
0 19886 5 2 1 94538
0 19887 7 1 2 73315 86004
0 19888 7 1 2 94539 19887
0 19889 5 1 1 19888
0 19890 7 1 2 19884 19889
0 19891 5 1 1 19890
0 19892 7 1 2 70689 19891
0 19893 5 1 1 19892
0 19894 7 1 2 72611 93356
0 19895 5 1 1 19894
0 19896 7 1 2 71319 89686
0 19897 5 1 1 19896
0 19898 7 1 2 19895 19897
0 19899 5 1 1 19898
0 19900 7 1 2 91148 19899
0 19901 5 1 1 19900
0 19902 7 1 2 19893 19901
0 19903 5 1 1 19902
0 19904 7 1 2 68393 19903
0 19905 5 1 1 19904
0 19906 7 1 2 86171 94450
0 19907 5 1 1 19906
0 19908 7 1 2 74801 93449
0 19909 5 1 1 19908
0 19910 7 1 2 19907 19909
0 19911 5 1 1 19910
0 19912 7 1 2 70325 19911
0 19913 5 1 1 19912
0 19914 7 1 2 90114 79228
0 19915 5 1 1 19914
0 19916 7 1 2 19913 19915
0 19917 5 1 1 19916
0 19918 7 1 2 80707 19917
0 19919 5 1 1 19918
0 19920 7 1 2 19905 19919
0 19921 5 1 1 19920
0 19922 7 1 2 92906 19921
0 19923 5 1 1 19922
0 19924 7 1 2 74490 93421
0 19925 5 1 1 19924
0 19926 7 1 2 75917 79578
0 19927 5 1 1 19926
0 19928 7 1 2 19925 19927
0 19929 5 1 1 19928
0 19930 7 1 2 87450 19929
0 19931 5 1 1 19930
0 19932 7 2 2 61841 77576
0 19933 7 1 2 81048 72373
0 19934 7 1 2 94543 19933
0 19935 5 1 1 19934
0 19936 7 1 2 19931 19935
0 19937 5 1 1 19936
0 19938 7 1 2 65732 19937
0 19939 5 1 1 19938
0 19940 7 3 2 68394 82051
0 19941 7 1 2 92992 94545
0 19942 7 1 2 88316 19941
0 19943 5 1 1 19942
0 19944 7 1 2 19939 19943
0 19945 5 1 1 19944
0 19946 7 1 2 88335 81766
0 19947 7 1 2 19945 19946
0 19948 5 1 1 19947
0 19949 7 1 2 63787 88790
0 19950 5 1 1 19949
0 19951 7 2 2 81767 88504
0 19952 5 3 1 94548
0 19953 7 1 2 66455 94550
0 19954 7 1 2 19950 19953
0 19955 5 1 1 19954
0 19956 7 1 2 61546 15139
0 19957 5 1 1 19956
0 19958 7 1 2 89512 92394
0 19959 7 1 2 19957 19958
0 19960 7 1 2 19955 19959
0 19961 5 1 1 19960
0 19962 7 1 2 71635 90749
0 19963 7 1 2 92271 19962
0 19964 5 1 1 19963
0 19965 7 1 2 19961 19964
0 19966 5 1 1 19965
0 19967 7 1 2 73433 19966
0 19968 5 1 1 19967
0 19969 7 1 2 66937 19968
0 19970 7 1 2 19948 19969
0 19971 7 1 2 19923 19970
0 19972 7 1 2 19874 19971
0 19973 5 1 1 19972
0 19974 7 1 2 64702 19973
0 19975 7 1 2 19744 19974
0 19976 5 1 1 19975
0 19977 7 1 2 89933 94491
0 19978 5 1 1 19977
0 19979 7 1 2 76922 19978
0 19980 5 1 1 19979
0 19981 7 1 2 88286 19980
0 19982 5 1 1 19981
0 19983 7 1 2 63788 82894
0 19984 5 1 1 19983
0 19985 7 1 2 67239 84582
0 19986 7 1 2 19984 19985
0 19987 5 1 1 19986
0 19988 7 1 2 19229 19987
0 19989 5 1 1 19988
0 19990 7 1 2 70326 19989
0 19991 5 1 1 19990
0 19992 7 1 2 75951 92346
0 19993 5 1 1 19992
0 19994 7 1 2 64111 19993
0 19995 7 1 2 19991 19994
0 19996 5 1 1 19995
0 19997 7 4 2 70327 88535
0 19998 5 1 1 94553
0 19999 7 1 2 62824 94554
0 20000 5 1 1 19999
0 20001 7 1 2 70904 74923
0 20002 7 1 2 82217 20001
0 20003 5 1 1 20002
0 20004 7 1 2 68972 20003
0 20005 7 1 2 20000 20004
0 20006 5 1 1 20005
0 20007 7 1 2 19996 20006
0 20008 5 1 1 20007
0 20009 7 1 2 87572 79917
0 20010 5 1 1 20009
0 20011 7 1 2 20008 20010
0 20012 5 1 1 20011
0 20013 7 1 2 70036 20012
0 20014 5 1 1 20013
0 20015 7 1 2 19982 20014
0 20016 5 1 1 20015
0 20017 7 1 2 66938 20016
0 20018 5 1 1 20017
0 20019 7 3 2 84380 73434
0 20020 5 1 1 94557
0 20021 7 1 2 71320 20020
0 20022 5 2 1 20021
0 20023 7 1 2 71941 94560
0 20024 5 1 1 20023
0 20025 7 1 2 74840 20024
0 20026 5 2 1 20025
0 20027 7 3 2 62074 76941
0 20028 5 1 1 94564
0 20029 7 1 2 94562 94565
0 20030 5 1 1 20029
0 20031 7 1 2 20018 20030
0 20032 5 1 1 20031
0 20033 7 1 2 65733 20032
0 20034 5 1 1 20033
0 20035 7 2 2 70690 86349
0 20036 7 1 2 89568 84836
0 20037 7 1 2 94567 20036
0 20038 5 1 1 20037
0 20039 7 1 2 76247 80874
0 20040 7 1 2 89843 20039
0 20041 5 1 1 20040
0 20042 7 1 2 20038 20041
0 20043 5 1 1 20042
0 20044 7 1 2 70905 20043
0 20045 5 1 1 20044
0 20046 7 1 2 76867 93542
0 20047 5 1 1 20046
0 20048 7 1 2 74953 86427
0 20049 5 1 1 20048
0 20050 7 1 2 20047 20049
0 20051 5 1 1 20050
0 20052 7 1 2 62566 20051
0 20053 5 1 1 20052
0 20054 7 1 2 71166 73435
0 20055 5 1 1 20054
0 20056 7 1 2 93225 20055
0 20057 5 1 1 20056
0 20058 7 1 2 67240 20057
0 20059 5 1 1 20058
0 20060 7 2 2 75529 84258
0 20061 7 1 2 70691 94569
0 20062 5 4 1 20061
0 20063 7 1 2 20059 94571
0 20064 5 1 1 20063
0 20065 7 1 2 70037 20064
0 20066 5 1 1 20065
0 20067 7 1 2 20053 20066
0 20068 5 1 1 20067
0 20069 7 1 2 66939 20068
0 20070 5 1 1 20069
0 20071 7 1 2 85250 94493
0 20072 5 1 1 20071
0 20073 7 1 2 77034 20072
0 20074 5 1 1 20073
0 20075 7 1 2 20070 20074
0 20076 5 1 1 20075
0 20077 7 1 2 68634 20076
0 20078 5 1 1 20077
0 20079 7 1 2 62075 84397
0 20080 5 2 1 20079
0 20081 7 2 2 74074 77659
0 20082 7 1 2 72272 94577
0 20083 5 1 1 20082
0 20084 7 1 2 94575 20083
0 20085 5 1 1 20084
0 20086 7 1 2 91952 20085
0 20087 5 1 1 20086
0 20088 7 1 2 20078 20087
0 20089 5 1 1 20088
0 20090 7 1 2 70328 20089
0 20091 5 1 1 20090
0 20092 7 1 2 20045 20091
0 20093 7 1 2 20034 20092
0 20094 5 1 1 20093
0 20095 7 1 2 68395 20094
0 20096 5 1 1 20095
0 20097 7 3 2 71490 91102
0 20098 7 1 2 76248 94579
0 20099 5 1 1 20098
0 20100 7 1 2 74075 85564
0 20101 5 1 1 20100
0 20102 7 1 2 77911 20101
0 20103 5 4 1 20102
0 20104 7 3 2 71942 94582
0 20105 5 1 1 94586
0 20106 7 1 2 77519 92082
0 20107 5 1 1 20106
0 20108 7 1 2 91236 20107
0 20109 7 1 2 20105 20108
0 20110 5 1 1 20109
0 20111 7 1 2 70329 20110
0 20112 5 1 1 20111
0 20113 7 1 2 20099 20112
0 20114 5 1 1 20113
0 20115 7 1 2 65129 75091
0 20116 7 1 2 20114 20115
0 20117 5 1 1 20116
0 20118 7 1 2 20096 20117
0 20119 5 1 1 20118
0 20120 7 1 2 66696 20119
0 20121 5 1 1 20120
0 20122 7 1 2 76204 82510
0 20123 7 1 2 85303 20122
0 20124 5 1 1 20123
0 20125 7 1 2 20121 20124
0 20126 5 1 1 20125
0 20127 7 1 2 78922 85642
0 20128 7 1 2 20126 20127
0 20129 5 1 1 20128
0 20130 7 1 2 19976 20129
0 20131 5 1 1 20130
0 20132 7 1 2 94393 20131
0 20133 5 1 1 20132
0 20134 7 5 2 67993 69086
0 20135 7 5 2 92209 94589
0 20136 7 1 2 84403 94594
0 20137 5 1 1 20136
0 20138 7 20 2 69356 93891
0 20139 7 2 2 91939 94599
0 20140 5 1 1 94619
0 20141 7 1 2 20137 20140
0 20142 5 1 1 20141
0 20143 7 1 2 65734 20142
0 20144 5 1 1 20143
0 20145 7 4 2 92129 94350
0 20146 7 3 2 90523 94621
0 20147 5 1 1 94625
0 20148 7 1 2 66456 94626
0 20149 5 1 1 20148
0 20150 7 1 2 20144 20149
0 20151 5 1 1 20150
0 20152 7 1 2 91463 20151
0 20153 5 1 1 20152
0 20154 7 14 2 64243 69357
0 20155 7 2 2 87830 94628
0 20156 7 1 2 79838 94642
0 20157 7 1 2 91940 20156
0 20158 5 1 1 20157
0 20159 7 1 2 20153 20158
0 20160 5 1 1 20159
0 20161 7 1 2 67241 20160
0 20162 5 1 1 20161
0 20163 7 2 2 84212 93892
0 20164 7 1 2 94304 94644
0 20165 7 1 2 91941 20164
0 20166 5 1 1 20165
0 20167 7 1 2 20162 20166
0 20168 5 1 1 20167
0 20169 7 1 2 67441 20168
0 20170 5 1 1 20169
0 20171 7 1 2 74910 79993
0 20172 5 1 1 20171
0 20173 7 6 2 64703 77237
0 20174 7 1 2 73926 80004
0 20175 5 1 1 20174
0 20176 7 1 2 94646 20175
0 20177 7 1 2 20172 20176
0 20178 5 1 1 20177
0 20179 7 4 2 76142 73436
0 20180 7 1 2 74915 91184
0 20181 7 1 2 94652 20180
0 20182 5 1 1 20181
0 20183 7 1 2 20178 20182
0 20184 5 1 1 20183
0 20185 7 1 2 94600 20184
0 20186 5 1 1 20185
0 20187 7 2 2 82759 94394
0 20188 7 3 2 64704 73437
0 20189 7 1 2 74903 75744
0 20190 7 1 2 94658 20189
0 20191 7 1 2 94656 20190
0 20192 5 1 1 20191
0 20193 7 1 2 20186 20192
0 20194 5 1 1 20193
0 20195 7 1 2 72135 20194
0 20196 5 1 1 20195
0 20197 7 1 2 70692 2199
0 20198 5 1 1 20197
0 20199 7 1 2 78299 94308
0 20200 7 1 2 20198 20199
0 20201 7 1 2 94620 20200
0 20202 5 1 1 20201
0 20203 7 1 2 20196 20202
0 20204 7 1 2 20170 20203
0 20205 5 1 1 20204
0 20206 7 1 2 65407 20205
0 20207 5 1 1 20206
0 20208 7 2 2 80531 73438
0 20209 7 3 2 68635 64244
0 20210 7 4 2 69182 94663
0 20211 7 1 2 69358 82413
0 20212 7 1 2 94666 20211
0 20213 7 1 2 94661 20212
0 20214 7 1 2 91942 20213
0 20215 5 1 1 20214
0 20216 7 1 2 20207 20215
0 20217 5 1 1 20216
0 20218 7 1 2 63311 20217
0 20219 5 1 1 20218
0 20220 7 1 2 77832 78947
0 20221 5 1 1 20220
0 20222 7 3 2 72136 71574
0 20223 7 1 2 78882 94670
0 20224 5 1 1 20223
0 20225 7 1 2 20221 20224
0 20226 5 1 1 20225
0 20227 7 1 2 61547 20226
0 20228 5 1 1 20227
0 20229 7 2 2 77816 81919
0 20230 5 1 1 94673
0 20231 7 1 2 88852 94674
0 20232 5 1 1 20231
0 20233 7 1 2 20228 20232
0 20234 5 1 1 20233
0 20235 7 1 2 62567 20234
0 20236 5 1 1 20235
0 20237 7 2 2 61548 63953
0 20238 7 1 2 78883 94675
0 20239 7 1 2 86804 20238
0 20240 5 1 1 20239
0 20241 7 1 2 20236 20240
0 20242 5 1 1 20241
0 20243 7 6 2 64245 91387
0 20244 7 1 2 94186 94677
0 20245 7 1 2 20242 20244
0 20246 5 1 1 20245
0 20247 7 1 2 20219 20246
0 20248 5 1 1 20247
0 20249 7 1 2 61842 20248
0 20250 5 1 1 20249
0 20251 7 1 2 83111 87587
0 20252 5 1 1 20251
0 20253 7 2 2 86172 87701
0 20254 5 1 1 94683
0 20255 7 1 2 68396 94684
0 20256 5 1 1 20255
0 20257 7 1 2 20252 20256
0 20258 5 1 1 20257
0 20259 7 1 2 70693 20258
0 20260 5 1 1 20259
0 20261 7 1 2 88505 75366
0 20262 7 1 2 92229 20261
0 20263 5 1 1 20262
0 20264 7 1 2 20260 20263
0 20265 5 1 1 20264
0 20266 7 1 2 72542 20265
0 20267 5 1 1 20266
0 20268 7 1 2 74802 87692
0 20269 5 1 1 20268
0 20270 7 1 2 20254 20269
0 20271 5 1 1 20270
0 20272 7 2 2 65735 79828
0 20273 7 1 2 20271 94685
0 20274 5 1 1 20273
0 20275 7 1 2 20267 20274
0 20276 5 1 1 20275
0 20277 7 1 2 67994 20276
0 20278 5 1 1 20277
0 20279 7 1 2 80741 86173
0 20280 7 1 2 87343 20279
0 20281 7 1 2 85405 20280
0 20282 5 1 1 20281
0 20283 7 1 2 20278 20282
0 20284 5 1 1 20283
0 20285 7 1 2 94395 20284
0 20286 5 1 1 20285
0 20287 7 1 2 79775 94315
0 20288 5 1 1 20287
0 20289 7 1 2 65736 87392
0 20290 5 1 1 20289
0 20291 7 1 2 20288 20290
0 20292 5 1 1 20291
0 20293 7 3 2 88914 93893
0 20294 7 1 2 77238 94687
0 20295 7 1 2 20292 20294
0 20296 5 1 1 20295
0 20297 7 1 2 20286 20296
0 20298 5 1 1 20297
0 20299 7 1 2 64705 20298
0 20300 5 1 1 20299
0 20301 7 6 2 64706 83112
0 20302 5 1 1 94690
0 20303 7 2 2 74283 86148
0 20304 5 1 1 94696
0 20305 7 1 2 14555 20304
0 20306 5 2 1 20305
0 20307 7 14 2 77239 94601
0 20308 7 1 2 94698 94700
0 20309 5 1 1 20308
0 20310 7 7 2 66457 64509
0 20311 7 7 2 94351 94714
0 20312 7 1 2 80207 94721
0 20313 7 1 2 94697 20312
0 20314 5 1 1 20313
0 20315 7 1 2 20309 20314
0 20316 5 1 1 20315
0 20317 7 1 2 94691 20316
0 20318 5 1 1 20317
0 20319 7 2 2 76143 94699
0 20320 7 13 2 64246 69548
0 20321 7 11 2 91388 94730
0 20322 7 1 2 83048 94743
0 20323 7 1 2 94728 20322
0 20324 5 1 1 20323
0 20325 7 1 2 20318 20324
0 20326 5 1 1 20325
0 20327 7 1 2 73776 20326
0 20328 5 1 1 20327
0 20329 7 1 2 91602 92907
0 20330 5 1 1 20329
0 20331 7 1 2 77726 92272
0 20332 5 1 1 20331
0 20333 7 1 2 20330 20332
0 20334 5 1 1 20333
0 20335 7 2 2 64339 82986
0 20336 7 7 2 68397 69087
0 20337 7 1 2 94754 94756
0 20338 7 1 2 20334 20337
0 20339 5 1 1 20338
0 20340 7 1 2 20328 20339
0 20341 5 1 1 20340
0 20342 7 1 2 70906 20341
0 20343 5 1 1 20342
0 20344 7 8 2 68827 64247
0 20345 7 2 2 67442 94763
0 20346 7 3 2 69183 82436
0 20347 7 1 2 83412 83531
0 20348 7 1 2 94773 20347
0 20349 7 1 2 94771 20348
0 20350 7 1 2 89182 20349
0 20351 5 1 1 20350
0 20352 7 1 2 20343 20351
0 20353 7 1 2 20300 20352
0 20354 5 1 1 20353
0 20355 7 1 2 70330 20354
0 20356 5 1 1 20355
0 20357 7 1 2 71321 77846
0 20358 5 2 1 20357
0 20359 7 1 2 72137 73316
0 20360 5 2 1 20359
0 20361 7 1 2 84036 94778
0 20362 7 1 2 94776 20361
0 20363 5 1 1 20362
0 20364 7 2 2 78510 90029
0 20365 7 6 2 63789 69184
0 20366 7 3 2 94629 94782
0 20367 7 1 2 82871 94788
0 20368 7 1 2 94780 20367
0 20369 7 1 2 20363 20368
0 20370 5 1 1 20369
0 20371 7 1 2 20356 20370
0 20372 7 1 2 20250 20371
0 20373 5 1 1 20372
0 20374 7 1 2 80569 20373
0 20375 5 1 1 20374
0 20376 7 2 2 69359 80859
0 20377 7 1 2 76556 94791
0 20378 5 1 1 20377
0 20379 7 3 2 61549 89282
0 20380 7 1 2 84499 87493
0 20381 7 1 2 94793 20380
0 20382 5 1 1 20381
0 20383 7 1 2 20378 20382
0 20384 5 1 1 20383
0 20385 7 1 2 70907 75452
0 20386 7 1 2 20384 20385
0 20387 5 1 1 20386
0 20388 7 1 2 82114 82469
0 20389 7 1 2 86648 20388
0 20390 7 1 2 89513 20389
0 20391 5 1 1 20390
0 20392 7 1 2 20387 20391
0 20393 5 1 1 20392
0 20394 7 1 2 71827 20393
0 20395 5 1 1 20394
0 20396 7 1 2 63550 83486
0 20397 5 1 1 20396
0 20398 7 1 2 88308 20397
0 20399 5 2 1 20398
0 20400 7 1 2 72138 94796
0 20401 5 1 1 20400
0 20402 7 2 2 66697 72543
0 20403 7 1 2 78071 94798
0 20404 5 1 1 20403
0 20405 7 1 2 20401 20404
0 20406 5 1 1 20405
0 20407 7 1 2 68636 80727
0 20408 7 1 2 85654 20407
0 20409 7 1 2 20406 20408
0 20410 5 1 1 20409
0 20411 7 1 2 20395 20410
0 20412 5 1 1 20411
0 20413 7 1 2 62076 20412
0 20414 5 1 1 20413
0 20415 7 1 2 71828 94797
0 20416 5 1 1 20415
0 20417 7 1 2 80716 89354
0 20418 5 3 1 20417
0 20419 7 1 2 90921 94800
0 20420 5 1 1 20419
0 20421 7 1 2 20416 20420
0 20422 5 1 1 20421
0 20423 7 1 2 72139 20422
0 20424 5 1 1 20423
0 20425 7 2 2 75952 79776
0 20426 5 1 1 94803
0 20427 7 1 2 87396 20426
0 20428 5 1 1 20427
0 20429 7 1 2 83268 20428
0 20430 5 1 1 20429
0 20431 7 1 2 20424 20430
0 20432 5 1 1 20431
0 20433 7 1 2 82699 90902
0 20434 7 1 2 20432 20433
0 20435 5 1 1 20434
0 20436 7 1 2 20414 20435
0 20437 5 1 1 20436
0 20438 7 1 2 63138 20437
0 20439 5 1 1 20438
0 20440 7 1 2 70038 85908
0 20441 5 1 1 20440
0 20442 7 1 2 1026 20441
0 20443 5 1 1 20442
0 20444 7 1 2 94205 20443
0 20445 5 1 1 20444
0 20446 7 1 2 77048 81035
0 20447 5 3 1 20446
0 20448 7 1 2 94804 94805
0 20449 5 1 1 20448
0 20450 7 1 2 75684 90513
0 20451 5 1 1 20450
0 20452 7 1 2 20449 20451
0 20453 7 1 2 20445 20452
0 20454 5 1 1 20453
0 20455 7 1 2 72140 20454
0 20456 5 1 1 20455
0 20457 7 1 2 62077 94206
0 20458 5 1 1 20457
0 20459 7 2 2 66940 76822
0 20460 7 1 2 63790 94808
0 20461 5 1 1 20460
0 20462 7 1 2 20458 20461
0 20463 5 4 1 20462
0 20464 7 1 2 66698 94810
0 20465 5 1 1 20464
0 20466 7 1 2 75417 86189
0 20467 5 1 1 20466
0 20468 7 1 2 20465 20467
0 20469 5 1 1 20468
0 20470 7 1 2 83269 20469
0 20471 5 1 1 20470
0 20472 7 1 2 20456 20471
0 20473 5 1 1 20472
0 20474 7 1 2 78755 91512
0 20475 7 1 2 20473 20474
0 20476 5 1 1 20475
0 20477 7 1 2 20439 20476
0 20478 5 1 1 20477
0 20479 7 1 2 63312 20478
0 20480 5 1 1 20479
0 20481 7 1 2 71829 94801
0 20482 5 1 1 20481
0 20483 7 1 2 63551 85483
0 20484 5 1 1 20483
0 20485 7 1 2 20482 20484
0 20486 5 1 1 20485
0 20487 7 1 2 62078 20486
0 20488 5 1 1 20487
0 20489 7 1 2 77660 88153
0 20490 5 1 1 20489
0 20491 7 1 2 20488 20490
0 20492 5 1 1 20491
0 20493 7 1 2 83863 20492
0 20494 5 1 1 20493
0 20495 7 4 2 63139 78511
0 20496 7 1 2 76918 78177
0 20497 7 1 2 94814 20496
0 20498 5 1 1 20497
0 20499 7 1 2 20494 20498
0 20500 5 1 1 20499
0 20501 7 1 2 72141 20500
0 20502 5 1 1 20501
0 20503 7 1 2 83864 94811
0 20504 5 1 1 20503
0 20505 7 1 2 75953 82618
0 20506 7 1 2 94299 20505
0 20507 5 1 1 20506
0 20508 7 1 2 20504 20507
0 20509 5 1 1 20508
0 20510 7 1 2 83270 20509
0 20511 5 1 1 20510
0 20512 7 1 2 20502 20511
0 20513 5 1 1 20512
0 20514 7 1 2 62568 86869
0 20515 7 1 2 20513 20514
0 20516 5 1 1 20515
0 20517 7 1 2 20480 20516
0 20518 5 1 1 20517
0 20519 7 1 2 69549 20518
0 20520 5 1 1 20519
0 20521 7 1 2 88662 90466
0 20522 5 1 1 20521
0 20523 7 1 2 81311 1418
0 20524 5 1 1 20523
0 20525 7 1 2 61843 4724
0 20526 7 1 2 20524 20525
0 20527 7 1 2 94207 20526
0 20528 5 1 1 20527
0 20529 7 1 2 20522 20528
0 20530 5 1 1 20529
0 20531 7 1 2 72142 20530
0 20532 5 1 1 20531
0 20533 7 1 2 82138 76234
0 20534 7 1 2 85394 20533
0 20535 5 1 1 20534
0 20536 7 1 2 20532 20535
0 20537 5 1 1 20536
0 20538 7 9 2 63140 69360
0 20539 7 5 2 61550 62569
0 20540 7 4 2 64707 94827
0 20541 7 1 2 94818 94832
0 20542 7 1 2 20537 20541
0 20543 5 1 1 20542
0 20544 7 1 2 20520 20543
0 20545 5 1 1 20544
0 20546 7 1 2 93894 20545
0 20547 5 1 1 20546
0 20548 7 1 2 70039 86914
0 20549 5 1 1 20548
0 20550 7 1 2 7240 20549
0 20551 5 1 1 20550
0 20552 7 1 2 61844 20551
0 20553 5 1 1 20552
0 20554 7 1 2 87181 75235
0 20555 5 1 1 20554
0 20556 7 1 2 20553 20555
0 20557 5 1 1 20556
0 20558 7 1 2 65975 20557
0 20559 5 1 1 20558
0 20560 7 1 2 75702 87083
0 20561 5 1 1 20560
0 20562 7 1 2 20559 20561
0 20563 5 1 1 20562
0 20564 7 1 2 68973 20563
0 20565 5 1 1 20564
0 20566 7 1 2 63313 78039
0 20567 7 1 2 75888 20566
0 20568 5 1 1 20567
0 20569 7 1 2 20565 20568
0 20570 5 1 1 20569
0 20571 7 1 2 94208 20570
0 20572 5 1 1 20571
0 20573 7 1 2 72223 86428
0 20574 5 1 1 20573
0 20575 7 1 2 94576 20574
0 20576 5 1 1 20575
0 20577 7 2 2 82139 84164
0 20578 5 2 1 94836
0 20579 7 1 2 94187 94838
0 20580 5 2 1 20579
0 20581 7 1 2 61845 94840
0 20582 7 1 2 20576 20581
0 20583 5 1 1 20582
0 20584 7 2 2 81447 75092
0 20585 7 1 2 85776 83271
0 20586 7 1 2 94842 20585
0 20587 5 1 1 20586
0 20588 7 1 2 20583 20587
0 20589 7 1 2 20572 20588
0 20590 5 1 1 20589
0 20591 7 1 2 67995 20590
0 20592 5 1 1 20591
0 20593 7 2 2 86321 94455
0 20594 7 1 2 75573 91709
0 20595 7 1 2 94844 20594
0 20596 5 1 1 20595
0 20597 7 1 2 20592 20596
0 20598 5 1 1 20597
0 20599 7 1 2 66458 20598
0 20600 5 1 1 20599
0 20601 7 1 2 67996 85186
0 20602 7 1 2 88522 20601
0 20603 7 1 2 94845 20602
0 20604 5 1 1 20603
0 20605 7 1 2 20600 20604
0 20606 5 1 1 20605
0 20607 7 13 2 82987 94352
0 20608 7 1 2 62570 94846
0 20609 7 1 2 20606 20608
0 20610 5 1 1 20609
0 20611 7 1 2 20547 20610
0 20612 5 1 1 20611
0 20613 7 1 2 71575 20612
0 20614 5 1 1 20613
0 20615 7 1 2 20375 20614
0 20616 7 1 2 20133 20615
0 20617 7 1 2 19538 20616
0 20618 5 1 1 20617
0 20619 7 1 2 69787 20618
0 20620 5 1 1 20619
0 20621 7 2 2 63314 81049
0 20622 5 2 1 94859
0 20623 7 5 2 68151 78072
0 20624 5 3 1 94863
0 20625 7 1 2 94861 94868
0 20626 5 10 1 20625
0 20627 7 1 2 62079 94871
0 20628 5 4 1 20627
0 20629 7 1 2 84785 91686
0 20630 5 1 1 20629
0 20631 7 1 2 94881 20630
0 20632 5 3 1 20631
0 20633 7 1 2 64919 94885
0 20634 5 1 1 20633
0 20635 7 3 2 66941 81326
0 20636 7 1 2 81362 94888
0 20637 5 1 1 20636
0 20638 7 1 2 20634 20637
0 20639 5 1 1 20638
0 20640 7 1 2 69550 20639
0 20641 5 1 1 20640
0 20642 7 1 2 89480 82036
0 20643 5 1 1 20642
0 20644 7 1 2 20641 20643
0 20645 5 1 1 20644
0 20646 7 1 2 66699 20645
0 20647 5 1 1 20646
0 20648 7 3 2 69788 88664
0 20649 5 1 1 94891
0 20650 7 2 2 83498 94892
0 20651 5 1 1 94894
0 20652 7 1 2 89477 20651
0 20653 5 1 1 20652
0 20654 7 1 2 77111 20653
0 20655 5 1 1 20654
0 20656 7 1 2 20647 20655
0 20657 5 1 1 20656
0 20658 7 1 2 67997 20657
0 20659 5 1 1 20658
0 20660 7 1 2 88943 79735
0 20661 7 1 2 88865 20660
0 20662 5 1 1 20661
0 20663 7 1 2 20659 20662
0 20664 5 1 1 20663
0 20665 7 1 2 66459 20664
0 20666 5 1 1 20665
0 20667 7 7 2 70040 79123
0 20668 7 1 2 80946 81854
0 20669 7 1 2 94896 20668
0 20670 5 1 1 20669
0 20671 7 1 2 20666 20670
0 20672 5 1 1 20671
0 20673 7 1 2 73439 85371
0 20674 7 1 2 20672 20673
0 20675 5 1 1 20674
0 20676 7 2 2 69789 71322
0 20677 7 1 2 83011 82031
0 20678 5 1 1 20677
0 20679 7 1 2 74218 3652
0 20680 7 1 2 83113 20679
0 20681 7 1 2 91687 20680
0 20682 5 1 1 20681
0 20683 7 1 2 20678 20682
0 20684 5 1 1 20683
0 20685 7 1 2 94903 20684
0 20686 5 1 1 20685
0 20687 7 2 2 74314 81768
0 20688 5 1 1 94905
0 20689 7 3 2 81633 74219
0 20690 5 1 1 94907
0 20691 7 1 2 20688 20690
0 20692 5 8 1 20691
0 20693 7 1 2 61846 94910
0 20694 5 2 1 20693
0 20695 7 1 2 75767 92262
0 20696 5 1 1 20695
0 20697 7 1 2 94918 20696
0 20698 5 1 1 20697
0 20699 7 1 2 65130 20698
0 20700 5 1 1 20699
0 20701 7 1 2 83439 82474
0 20702 5 1 1 20701
0 20703 7 1 2 20700 20702
0 20704 5 1 1 20703
0 20705 7 1 2 75623 20704
0 20706 5 1 1 20705
0 20707 7 1 2 20686 20706
0 20708 5 1 1 20707
0 20709 7 1 2 72612 20708
0 20710 5 1 1 20709
0 20711 7 2 2 69790 80208
0 20712 7 1 2 61847 94920
0 20713 5 1 1 20712
0 20714 7 1 2 76019 20713
0 20715 5 1 1 20714
0 20716 7 1 2 88665 91688
0 20717 7 1 2 20715 20716
0 20718 5 1 1 20717
0 20719 7 1 2 65131 77009
0 20720 7 1 2 94911 20719
0 20721 5 1 1 20720
0 20722 7 1 2 20718 20721
0 20723 5 1 1 20722
0 20724 7 1 2 72055 20723
0 20725 5 1 1 20724
0 20726 7 1 2 20710 20725
0 20727 5 1 1 20726
0 20728 7 1 2 71729 20727
0 20729 5 1 1 20728
0 20730 7 1 2 90176 15734
0 20731 5 1 1 20730
0 20732 7 1 2 69791 20731
0 20733 7 1 2 94462 20732
0 20734 5 1 1 20733
0 20735 7 1 2 72056 77010
0 20736 5 1 1 20735
0 20737 7 1 2 72613 71459
0 20738 5 2 1 20737
0 20739 7 2 2 72614 71054
0 20740 5 1 1 94924
0 20741 7 1 2 62825 94925
0 20742 5 1 1 20741
0 20743 7 1 2 94922 20742
0 20744 7 1 2 20736 20743
0 20745 5 1 1 20744
0 20746 7 1 2 81732 80676
0 20747 7 1 2 20745 20746
0 20748 5 1 1 20747
0 20749 7 1 2 20734 20748
0 20750 5 1 1 20749
0 20751 7 1 2 75139 20750
0 20752 5 1 1 20751
0 20753 7 1 2 75140 75663
0 20754 7 1 2 87241 20753
0 20755 5 1 1 20754
0 20756 7 2 2 64920 94528
0 20757 7 1 2 75093 76667
0 20758 7 1 2 94926 20757
0 20759 5 1 1 20758
0 20760 7 1 2 20755 20759
0 20761 5 1 1 20760
0 20762 7 1 2 63315 20761
0 20763 5 1 1 20762
0 20764 7 1 2 75141 92064
0 20765 7 1 2 92263 20764
0 20766 5 1 1 20765
0 20767 7 1 2 65132 20766
0 20768 7 1 2 20763 20767
0 20769 5 1 1 20768
0 20770 7 1 2 82032 83413
0 20771 5 1 1 20770
0 20772 7 1 2 94919 20771
0 20773 5 1 1 20772
0 20774 7 1 2 94927 20773
0 20775 5 1 1 20774
0 20776 7 1 2 72544 82895
0 20777 5 3 1 20776
0 20778 7 1 2 89949 94928
0 20779 5 1 1 20778
0 20780 7 1 2 71431 94912
0 20781 5 1 1 20780
0 20782 7 1 2 87242 92696
0 20783 5 1 1 20782
0 20784 7 1 2 20781 20783
0 20785 5 1 1 20784
0 20786 7 1 2 20779 20785
0 20787 5 1 1 20786
0 20788 7 1 2 70041 20787
0 20789 7 1 2 20775 20788
0 20790 5 1 1 20789
0 20791 7 1 2 65408 20790
0 20792 7 1 2 20769 20791
0 20793 5 1 1 20792
0 20794 7 1 2 20752 20793
0 20795 7 1 2 20729 20794
0 20796 5 1 1 20795
0 20797 7 1 2 64708 20796
0 20798 5 1 1 20797
0 20799 7 1 2 84026 73662
0 20800 5 2 1 20799
0 20801 7 1 2 75106 94931
0 20802 5 1 1 20801
0 20803 7 1 2 84750 93712
0 20804 5 1 1 20803
0 20805 7 1 2 20802 20804
0 20806 5 1 1 20805
0 20807 7 1 2 73440 20806
0 20808 5 1 1 20807
0 20809 7 2 2 83728 77313
0 20810 7 1 2 79829 94933
0 20811 5 1 1 20810
0 20812 7 1 2 20808 20811
0 20813 5 1 1 20812
0 20814 7 1 2 88202 20813
0 20815 5 1 1 20814
0 20816 7 16 2 78090 81060
0 20817 7 4 2 77520 93431
0 20818 5 1 1 94951
0 20819 7 1 2 89950 20818
0 20820 5 3 1 20819
0 20821 7 1 2 81448 94955
0 20822 5 1 1 20821
0 20823 7 1 2 83049 89944
0 20824 5 1 1 20823
0 20825 7 1 2 20822 20824
0 20826 5 1 1 20825
0 20827 7 1 2 84195 20826
0 20828 5 1 1 20827
0 20829 7 2 2 85265 90846
0 20830 5 1 1 94958
0 20831 7 1 2 72615 86453
0 20832 7 1 2 94959 20831
0 20833 5 1 1 20832
0 20834 7 1 2 20828 20833
0 20835 5 1 1 20834
0 20836 7 1 2 94935 20835
0 20837 5 1 1 20836
0 20838 7 1 2 20815 20837
0 20839 5 1 1 20838
0 20840 7 1 2 64921 20839
0 20841 5 1 1 20840
0 20842 7 1 2 79736 85187
0 20843 7 1 2 90117 20842
0 20844 7 1 2 86333 92429
0 20845 7 1 2 20843 20844
0 20846 5 1 1 20845
0 20847 7 1 2 20841 20846
0 20848 5 1 1 20847
0 20849 7 1 2 78923 20848
0 20850 5 1 1 20849
0 20851 7 1 2 20798 20850
0 20852 5 1 1 20851
0 20853 7 1 2 66460 20852
0 20854 5 1 1 20853
0 20855 7 1 2 78924 94956
0 20856 5 1 1 20855
0 20857 7 3 2 64709 94529
0 20858 7 1 2 63141 94960
0 20859 5 1 1 20858
0 20860 7 1 2 20856 20859
0 20861 5 1 1 20860
0 20862 7 1 2 86051 20861
0 20863 5 1 1 20862
0 20864 7 1 2 71323 78925
0 20865 5 1 1 20864
0 20866 7 1 2 89062 91175
0 20867 7 1 2 20865 20866
0 20868 5 1 1 20867
0 20869 7 1 2 72616 93938
0 20870 7 1 2 20868 20869
0 20871 5 1 1 20870
0 20872 7 1 2 20863 20871
0 20873 5 1 1 20872
0 20874 7 1 2 66461 20873
0 20875 5 1 1 20874
0 20876 7 1 2 86052 77521
0 20877 5 1 1 20876
0 20878 7 3 2 74111 71730
0 20879 7 1 2 77930 94963
0 20880 5 1 1 20879
0 20881 7 1 2 20877 20880
0 20882 5 1 1 20881
0 20883 7 1 2 89081 20882
0 20884 5 1 1 20883
0 20885 7 1 2 20875 20884
0 20886 5 1 1 20885
0 20887 7 1 2 78839 20886
0 20888 5 1 1 20887
0 20889 7 1 2 79124 72848
0 20890 7 1 2 90516 20889
0 20891 7 1 2 94524 20890
0 20892 5 1 1 20891
0 20893 7 1 2 20888 20892
0 20894 5 1 1 20893
0 20895 7 1 2 94872 20894
0 20896 5 1 1 20895
0 20897 7 1 2 85877 82498
0 20898 5 1 1 20897
0 20899 7 2 2 65409 78105
0 20900 7 1 2 70908 94966
0 20901 5 1 1 20900
0 20902 7 1 2 20898 20901
0 20903 5 1 1 20902
0 20904 7 1 2 66942 20903
0 20905 5 1 1 20904
0 20906 7 1 2 76342 81064
0 20907 5 1 1 20906
0 20908 7 1 2 20905 20907
0 20909 5 1 1 20908
0 20910 7 1 2 73441 20909
0 20911 5 1 1 20910
0 20912 7 1 2 81134 5458
0 20913 5 1 1 20912
0 20914 7 1 2 62826 20913
0 20915 5 2 1 20914
0 20916 7 2 2 70042 72617
0 20917 5 1 1 94970
0 20918 7 1 2 71324 1900
0 20919 7 1 2 20917 20918
0 20920 7 1 2 83880 20919
0 20921 5 1 1 20920
0 20922 7 1 2 94968 20921
0 20923 5 1 1 20922
0 20924 7 1 2 74315 20923
0 20925 5 1 1 20924
0 20926 7 1 2 20911 20925
0 20927 5 1 1 20926
0 20928 7 1 2 88944 20927
0 20929 5 1 1 20928
0 20930 7 2 2 65410 84786
0 20931 7 1 2 77522 94972
0 20932 5 1 1 20931
0 20933 7 1 2 74112 88666
0 20934 7 1 2 74199 20933
0 20935 5 1 1 20934
0 20936 7 1 2 20932 20935
0 20937 5 1 1 20936
0 20938 7 1 2 64922 91689
0 20939 7 1 2 20937 20938
0 20940 5 1 1 20939
0 20941 7 1 2 20929 20940
0 20942 5 1 1 20941
0 20943 7 1 2 66700 20942
0 20944 5 1 1 20943
0 20945 7 1 2 72826 85395
0 20946 5 1 1 20945
0 20947 7 1 2 7810 20946
0 20948 5 1 1 20947
0 20949 7 1 2 74316 92007
0 20950 7 1 2 20948 20949
0 20951 5 1 1 20950
0 20952 7 1 2 20944 20951
0 20953 5 1 1 20952
0 20954 7 1 2 89082 20953
0 20955 5 1 1 20954
0 20956 7 1 2 20896 20955
0 20957 7 1 2 20854 20956
0 20958 7 1 2 20675 20957
0 20959 5 1 1 20958
0 20960 7 1 2 94396 20959
0 20961 5 1 1 20960
0 20962 7 2 2 87403 80046
0 20963 5 1 1 94974
0 20964 7 1 2 74357 94975
0 20965 5 1 1 20964
0 20966 7 1 2 62080 82644
0 20967 5 1 1 20966
0 20968 7 1 2 20965 20967
0 20969 5 1 1 20968
0 20970 7 1 2 78551 20969
0 20971 5 1 1 20970
0 20972 7 5 2 65133 75796
0 20973 7 1 2 91103 94976
0 20974 7 1 2 87385 20973
0 20975 5 1 1 20974
0 20976 7 1 2 20971 20975
0 20977 5 1 1 20976
0 20978 7 1 2 63142 20977
0 20979 5 1 1 20978
0 20980 7 5 2 78604 75797
0 20981 5 1 1 94981
0 20982 7 1 2 78578 20981
0 20983 5 2 1 20982
0 20984 7 1 2 80786 91162
0 20985 7 1 2 94986 20984
0 20986 5 1 1 20985
0 20987 7 1 2 20979 20986
0 20988 5 1 1 20987
0 20989 7 1 2 61848 20988
0 20990 5 1 1 20989
0 20991 7 1 2 83590 83518
0 20992 5 2 1 20991
0 20993 7 1 2 79076 94977
0 20994 5 1 1 20993
0 20995 7 1 2 94988 20994
0 20996 5 1 1 20995
0 20997 7 1 2 91104 92919
0 20998 7 1 2 20996 20997
0 20999 5 1 1 20998
0 21000 7 1 2 20990 20999
0 21001 5 1 1 21000
0 21002 7 1 2 63316 21001
0 21003 5 1 1 21002
0 21004 7 1 2 82358 94864
0 21005 7 1 2 79202 21004
0 21006 5 1 1 21005
0 21007 7 1 2 21003 21006
0 21008 5 1 1 21007
0 21009 7 1 2 62571 21008
0 21010 5 1 1 21009
0 21011 7 2 2 81634 91579
0 21012 7 1 2 89213 90094
0 21013 7 1 2 94990 21012
0 21014 5 1 1 21013
0 21015 7 1 2 21010 21014
0 21016 5 1 1 21015
0 21017 7 1 2 73120 21016
0 21018 5 1 1 21017
0 21019 7 1 2 62081 91690
0 21020 5 1 1 21019
0 21021 7 1 2 1761 21020
0 21022 5 10 1 21021
0 21023 7 2 2 82375 75624
0 21024 5 1 1 95002
0 21025 7 2 2 83114 77682
0 21026 5 1 1 95004
0 21027 7 1 2 21024 21026
0 21028 5 1 1 21027
0 21029 7 1 2 64710 21028
0 21030 5 1 1 21029
0 21031 7 2 2 74968 78260
0 21032 5 3 1 95006
0 21033 7 1 2 68152 95007
0 21034 5 1 1 21033
0 21035 7 1 2 21030 21034
0 21036 5 1 1 21035
0 21037 7 1 2 63143 21036
0 21038 5 1 1 21037
0 21039 7 2 2 81986 81247
0 21040 7 1 2 81814 95011
0 21041 5 1 1 21040
0 21042 7 1 2 21038 21041
0 21043 5 1 1 21042
0 21044 7 1 2 61551 21043
0 21045 5 1 1 21044
0 21046 7 1 2 88945 81248
0 21047 7 1 2 88871 21046
0 21048 5 1 1 21047
0 21049 7 1 2 21045 21048
0 21050 5 1 1 21049
0 21051 7 1 2 94992 21050
0 21052 5 1 1 21051
0 21053 7 1 2 81987 78948
0 21054 5 1 1 21053
0 21055 7 1 2 83238 21054
0 21056 5 4 1 21055
0 21057 7 1 2 61552 95013
0 21058 5 1 1 21057
0 21059 7 2 2 69551 92926
0 21060 5 1 1 95017
0 21061 7 1 2 21058 21060
0 21062 5 7 1 21061
0 21063 7 2 2 89209 95019
0 21064 7 1 2 77314 95026
0 21065 5 1 1 21064
0 21066 7 1 2 21052 21065
0 21067 5 1 1 21066
0 21068 7 1 2 70909 21067
0 21069 5 1 1 21068
0 21070 7 2 2 62827 88188
0 21071 7 1 2 88712 95005
0 21072 7 1 2 95028 21071
0 21073 5 1 1 21072
0 21074 7 1 2 21069 21073
0 21075 5 1 1 21074
0 21076 7 1 2 70331 21075
0 21077 5 1 1 21076
0 21078 7 1 2 21018 21077
0 21079 5 1 1 21078
0 21080 7 1 2 64112 21079
0 21081 5 1 1 21080
0 21082 7 4 2 69792 76144
0 21083 7 1 2 88648 80541
0 21084 5 1 1 21083
0 21085 7 1 2 77128 86435
0 21086 7 1 2 89679 21085
0 21087 5 1 1 21086
0 21088 7 1 2 21084 21087
0 21089 5 1 1 21088
0 21090 7 1 2 95030 21089
0 21091 5 1 1 21090
0 21092 7 1 2 63317 78677
0 21093 7 2 2 94815 21092
0 21094 7 1 2 80542 95034
0 21095 5 1 1 21094
0 21096 7 1 2 21091 21095
0 21097 5 1 1 21096
0 21098 7 1 2 69552 21097
0 21099 5 1 1 21098
0 21100 7 1 2 80536 78412
0 21101 7 1 2 81381 92892
0 21102 7 1 2 21100 21101
0 21103 5 1 1 21102
0 21104 7 1 2 21099 21103
0 21105 5 1 1 21104
0 21106 7 1 2 75142 21105
0 21107 5 1 1 21106
0 21108 7 1 2 61849 92697
0 21109 5 1 1 21108
0 21110 7 1 2 12846 21109
0 21111 5 3 1 21110
0 21112 7 1 2 89514 95036
0 21113 5 1 1 21112
0 21114 7 5 2 61850 65737
0 21115 7 3 2 65976 75798
0 21116 7 1 2 87199 79655
0 21117 7 1 2 95044 21116
0 21118 5 1 1 21117
0 21119 7 3 2 62082 81582
0 21120 5 1 1 95047
0 21121 7 1 2 10641 21120
0 21122 7 1 2 21118 21121
0 21123 5 1 1 21122
0 21124 7 1 2 95039 21123
0 21125 5 1 1 21124
0 21126 7 1 2 21113 21125
0 21127 5 1 1 21126
0 21128 7 1 2 69793 21127
0 21129 5 1 1 21128
0 21130 7 1 2 89481 91071
0 21131 5 1 1 21130
0 21132 7 1 2 21129 21131
0 21133 5 1 1 21132
0 21134 7 1 2 65411 21133
0 21135 5 1 1 21134
0 21136 7 3 2 63318 74601
0 21137 7 1 2 67674 75063
0 21138 7 1 2 95050 21137
0 21139 7 1 2 91049 21138
0 21140 5 1 1 21139
0 21141 7 1 2 21135 21140
0 21142 5 1 1 21141
0 21143 7 1 2 70043 21142
0 21144 5 1 1 21143
0 21145 7 2 2 76368 76705
0 21146 5 1 1 95053
0 21147 7 1 2 75799 80381
0 21148 5 1 1 21147
0 21149 7 1 2 21146 21148
0 21150 5 1 1 21149
0 21151 7 2 2 78040 21150
0 21152 7 1 2 87200 79290
0 21153 7 1 2 86414 21152
0 21154 7 1 2 95055 21153
0 21155 5 1 1 21154
0 21156 7 1 2 21144 21155
0 21157 5 1 1 21156
0 21158 7 1 2 69553 21157
0 21159 5 1 1 21158
0 21160 7 1 2 77270 21159
0 21161 5 1 1 21160
0 21162 7 1 2 80537 92698
0 21163 5 1 1 21162
0 21164 7 1 2 82580 75800
0 21165 7 1 2 86220 21164
0 21166 5 1 1 21165
0 21167 7 1 2 21163 21166
0 21168 5 1 1 21167
0 21169 7 1 2 65412 21168
0 21170 5 1 1 21169
0 21171 7 1 2 73635 93462
0 21172 5 1 1 21171
0 21173 7 1 2 21170 21172
0 21174 5 1 1 21173
0 21175 7 1 2 70044 21174
0 21176 5 1 1 21175
0 21177 7 1 2 72699 83225
0 21178 7 1 2 95056 21177
0 21179 5 1 1 21178
0 21180 7 1 2 21176 21179
0 21181 5 1 1 21180
0 21182 7 1 2 79172 21181
0 21183 5 1 1 21182
0 21184 7 2 2 89025 6094
0 21185 5 1 1 95057
0 21186 7 3 2 75768 82544
0 21187 5 2 1 95059
0 21188 7 1 2 21185 95060
0 21189 5 1 1 21188
0 21190 7 3 2 81371 74317
0 21191 5 1 1 95064
0 21192 7 1 2 89831 95065
0 21193 5 1 1 21192
0 21194 7 1 2 21189 21193
0 21195 5 1 1 21194
0 21196 7 1 2 76891 21195
0 21197 5 1 1 21196
0 21198 7 1 2 77240 21197
0 21199 7 1 2 21183 21198
0 21200 5 1 1 21199
0 21201 7 1 2 81003 21200
0 21202 7 1 2 21161 21201
0 21203 5 1 1 21202
0 21204 7 1 2 21107 21203
0 21205 7 1 2 21081 21204
0 21206 5 1 1 21205
0 21207 7 1 2 94602 21206
0 21208 5 1 1 21207
0 21209 7 1 2 20961 21208
0 21210 5 1 1 21209
0 21211 7 1 2 73003 21210
0 21212 5 1 1 21211
0 21213 7 2 2 70332 72784
0 21214 7 1 2 77148 94503
0 21215 5 1 1 21214
0 21216 7 3 2 66943 91691
0 21217 5 2 1 95069
0 21218 7 1 2 77614 95070
0 21219 5 1 1 21218
0 21220 7 1 2 21215 21219
0 21221 5 1 1 21220
0 21222 7 1 2 77601 21221
0 21223 5 1 1 21222
0 21224 7 1 2 94321 94993
0 21225 5 1 1 21224
0 21226 7 1 2 21223 21225
0 21227 5 1 1 21226
0 21228 7 1 2 76082 21227
0 21229 5 1 1 21228
0 21230 7 1 2 63791 94653
0 21231 7 1 2 94994 21230
0 21232 5 1 1 21231
0 21233 7 1 2 21229 21232
0 21234 5 1 1 21233
0 21235 7 1 2 95067 21234
0 21236 5 1 1 21235
0 21237 7 2 2 71830 91692
0 21238 5 1 1 95074
0 21239 7 1 2 18036 21238
0 21240 5 1 1 21239
0 21241 7 1 2 62083 21240
0 21242 5 1 1 21241
0 21243 7 1 2 13058 21242
0 21244 5 2 1 21243
0 21245 7 2 2 71325 76145
0 21246 7 2 2 89515 95078
0 21247 7 1 2 95076 95080
0 21248 5 1 1 21247
0 21249 7 1 2 79015 75094
0 21250 5 1 1 21249
0 21251 7 1 2 78106 73808
0 21252 5 1 1 21251
0 21253 7 1 2 21250 21252
0 21254 5 1 1 21253
0 21255 7 2 2 73317 21254
0 21256 5 1 1 95082
0 21257 7 2 2 63792 75107
0 21258 7 1 2 70045 73442
0 21259 7 1 2 95084 21258
0 21260 5 1 1 21259
0 21261 7 1 2 21256 21260
0 21262 5 1 1 21261
0 21263 7 1 2 70910 86896
0 21264 7 1 2 21262 21263
0 21265 5 1 1 21264
0 21266 7 1 2 88827 94115
0 21267 7 1 2 93975 21266
0 21268 5 1 1 21267
0 21269 7 1 2 21265 21268
0 21270 5 1 1 21269
0 21271 7 1 2 76146 21270
0 21272 5 1 1 21271
0 21273 7 1 2 21248 21272
0 21274 7 1 2 21236 21273
0 21275 5 1 1 21274
0 21276 7 1 2 66701 21275
0 21277 5 1 1 21276
0 21278 7 1 2 85266 94729
0 21279 5 1 1 21278
0 21280 7 1 2 86762 84465
0 21281 7 1 2 86190 21280
0 21282 5 1 1 21281
0 21283 7 1 2 21279 21282
0 21284 5 1 1 21283
0 21285 7 1 2 77491 80570
0 21286 7 1 2 21284 21285
0 21287 5 1 1 21286
0 21288 7 1 2 21277 21287
0 21289 5 1 1 21288
0 21290 7 1 2 64711 21289
0 21291 5 1 1 21290
0 21292 7 2 2 68637 83742
0 21293 7 1 2 72933 94444
0 21294 5 1 1 21293
0 21295 7 1 2 95086 21294
0 21296 5 1 1 21295
0 21297 7 1 2 94464 21296
0 21298 5 1 1 21297
0 21299 7 1 2 88828 21298
0 21300 5 1 1 21299
0 21301 7 1 2 65413 84735
0 21302 5 1 1 21301
0 21303 7 1 2 71831 94995
0 21304 7 1 2 21302 21303
0 21305 5 1 1 21304
0 21306 7 1 2 21300 21305
0 21307 5 1 1 21306
0 21308 7 1 2 80057 87261
0 21309 7 1 2 21307 21308
0 21310 5 1 1 21309
0 21311 7 1 2 21291 21310
0 21312 5 1 1 21311
0 21313 7 1 2 94397 21312
0 21314 5 1 1 21313
0 21315 7 1 2 63552 89774
0 21316 5 1 1 21315
0 21317 7 1 2 70046 80430
0 21318 5 1 1 21317
0 21319 7 1 2 21316 21318
0 21320 5 1 1 21319
0 21321 7 1 2 62084 21320
0 21322 5 1 1 21321
0 21323 7 3 2 66944 74271
0 21324 7 1 2 79606 95088
0 21325 5 1 1 21324
0 21326 7 1 2 21322 21325
0 21327 5 1 1 21326
0 21328 7 1 2 73443 21327
0 21329 5 1 1 21328
0 21330 7 1 2 93473 94048
0 21331 5 1 1 21330
0 21332 7 1 2 77071 78155
0 21333 7 1 2 75143 21332
0 21334 5 1 1 21333
0 21335 7 1 2 80708 73809
0 21336 5 1 1 21335
0 21337 7 1 2 78150 86607
0 21338 7 1 2 840 21337
0 21339 5 1 1 21338
0 21340 7 1 2 21336 21339
0 21341 7 1 2 21334 21340
0 21342 5 1 1 21341
0 21343 7 1 2 86550 21342
0 21344 5 1 1 21343
0 21345 7 1 2 21331 21344
0 21346 7 1 2 21329 21345
0 21347 5 1 1 21346
0 21348 7 1 2 72057 21347
0 21349 5 1 1 21348
0 21350 7 1 2 88136 95077
0 21351 5 1 1 21350
0 21352 7 1 2 21349 21351
0 21353 5 1 1 21352
0 21354 7 9 2 89260 94678
0 21355 5 1 1 95091
0 21356 7 1 2 76668 95092
0 21357 7 1 2 21353 21356
0 21358 5 1 1 21357
0 21359 7 1 2 68153 21358
0 21360 7 1 2 21314 21359
0 21361 5 1 1 21360
0 21362 7 6 2 93895 94819
0 21363 7 1 2 80047 95100
0 21364 5 1 1 21363
0 21365 7 1 2 81516 94847
0 21366 5 1 1 21365
0 21367 7 1 2 21364 21366
0 21368 5 1 1 21367
0 21369 7 1 2 86053 21368
0 21370 5 1 1 21369
0 21371 7 12 2 69088 92210
0 21372 7 4 2 88096 95106
0 21373 7 1 2 67998 94067
0 21374 7 1 2 95118 21373
0 21375 5 1 1 21374
0 21376 7 1 2 21370 21375
0 21377 5 1 1 21376
0 21378 7 1 2 77112 21377
0 21379 5 1 1 21378
0 21380 7 2 2 65134 82988
0 21381 7 1 2 80604 94353
0 21382 7 1 2 84998 21381
0 21383 7 1 2 95122 21382
0 21384 5 1 1 21383
0 21385 7 1 2 21379 21384
0 21386 5 1 1 21385
0 21387 7 1 2 63553 21386
0 21388 5 1 1 21387
0 21389 7 1 2 85100 87108
0 21390 7 1 2 90475 21389
0 21391 7 3 2 69185 70047
0 21392 7 4 2 94630 95124
0 21393 7 1 2 65977 75032
0 21394 7 1 2 95127 21393
0 21395 7 1 2 21390 21394
0 21396 5 1 1 21395
0 21397 7 1 2 21388 21396
0 21398 5 1 1 21397
0 21399 7 1 2 64113 21398
0 21400 5 1 1 21399
0 21401 7 1 2 66945 77634
0 21402 5 4 1 21401
0 21403 7 1 2 62085 90326
0 21404 5 1 1 21403
0 21405 7 1 2 89201 92159
0 21406 7 1 2 21404 21405
0 21407 7 1 2 95131 21406
0 21408 5 1 1 21407
0 21409 7 2 2 65978 93290
0 21410 7 1 2 81050 73738
0 21411 7 1 2 78261 21410
0 21412 7 1 2 95135 21411
0 21413 5 1 1 21412
0 21414 7 1 2 21408 21413
0 21415 5 1 1 21414
0 21416 7 1 2 94595 21415
0 21417 5 1 1 21416
0 21418 7 1 2 21400 21417
0 21419 5 1 1 21418
0 21420 7 1 2 62828 21419
0 21421 5 1 1 21420
0 21422 7 1 2 85251 78262
0 21423 7 1 2 93458 21422
0 21424 5 1 1 21423
0 21425 7 2 2 83499 77113
0 21426 7 1 2 71326 73576
0 21427 7 1 2 95137 21426
0 21428 5 1 1 21427
0 21429 7 1 2 21424 21428
0 21430 5 1 1 21429
0 21431 7 1 2 68974 21430
0 21432 5 1 1 21431
0 21433 7 1 2 67675 76732
0 21434 5 2 1 21433
0 21435 7 1 2 85614 95139
0 21436 5 1 1 21435
0 21437 7 1 2 95138 21436
0 21438 5 1 1 21437
0 21439 7 1 2 21432 21438
0 21440 5 1 1 21439
0 21441 7 1 2 94596 21440
0 21442 5 1 1 21441
0 21443 7 3 2 69186 69554
0 21444 7 1 2 63554 77114
0 21445 7 1 2 95141 21444
0 21446 7 11 2 63144 64248
0 21447 7 3 2 69361 95144
0 21448 7 1 2 88137 95155
0 21449 7 1 2 21445 21448
0 21450 5 1 1 21449
0 21451 7 1 2 21442 21450
0 21452 5 1 1 21451
0 21453 7 1 2 86054 21452
0 21454 5 1 1 21453
0 21455 7 1 2 77177 93243
0 21456 7 2 2 78790 73962
0 21457 7 1 2 95107 95158
0 21458 7 1 2 21455 21457
0 21459 5 1 1 21458
0 21460 7 1 2 68638 21459
0 21461 7 1 2 21454 21460
0 21462 7 1 2 21421 21461
0 21463 5 1 1 21462
0 21464 7 3 2 64712 78041
0 21465 7 1 2 78178 95108
0 21466 7 1 2 95160 21465
0 21467 5 1 1 21466
0 21468 7 1 2 84500 73608
0 21469 7 1 2 75244 21468
0 21470 7 1 2 94744 21469
0 21471 5 1 1 21470
0 21472 7 1 2 21467 21471
0 21473 5 1 1 21472
0 21474 7 1 2 66702 21473
0 21475 5 1 1 21474
0 21476 7 7 2 63954 64249
0 21477 7 1 2 77945 91105
0 21478 7 1 2 95163 21477
0 21479 7 1 2 90578 92684
0 21480 7 1 2 21478 21479
0 21481 5 1 1 21480
0 21482 7 1 2 21475 21481
0 21483 5 1 1 21482
0 21484 7 1 2 63145 21483
0 21485 5 1 1 21484
0 21486 7 4 2 70333 72618
0 21487 5 2 1 95170
0 21488 7 2 2 89472 95171
0 21489 7 2 2 83331 74220
0 21490 7 4 2 63955 69089
0 21491 7 3 2 92211 95180
0 21492 7 1 2 81051 95184
0 21493 7 1 2 95178 21492
0 21494 7 1 2 95176 21493
0 21495 5 1 1 21494
0 21496 7 1 2 21485 21495
0 21497 5 1 1 21496
0 21498 7 1 2 62572 21497
0 21499 5 1 1 21498
0 21500 7 1 2 72249 95161
0 21501 7 3 2 63146 69090
0 21502 7 3 2 92212 95187
0 21503 7 6 2 68398 82619
0 21504 7 1 2 95190 95193
0 21505 7 1 2 21500 21504
0 21506 5 1 1 21505
0 21507 7 1 2 21499 21506
0 21508 5 1 1 21507
0 21509 7 1 2 62401 21508
0 21510 5 1 1 21509
0 21511 7 1 2 76892 90425
0 21512 7 1 2 80177 94603
0 21513 7 1 2 21511 21512
0 21514 5 1 1 21513
0 21515 7 1 2 86608 87916
0 21516 5 1 1 21515
0 21517 7 1 2 94059 21516
0 21518 5 1 1 21517
0 21519 7 2 2 65135 92213
0 21520 7 1 2 79737 94590
0 21521 7 1 2 95199 21520
0 21522 7 1 2 21518 21521
0 21523 5 1 1 21522
0 21524 7 1 2 21514 21523
0 21525 5 1 1 21524
0 21526 7 1 2 80048 21525
0 21527 5 1 1 21526
0 21528 7 1 2 82620 80742
0 21529 7 1 2 88681 21528
0 21530 7 1 2 79888 94848
0 21531 7 1 2 21529 21530
0 21532 5 1 1 21531
0 21533 7 1 2 21527 21532
0 21534 5 1 1 21533
0 21535 7 1 2 68975 21534
0 21536 5 1 1 21535
0 21537 7 1 2 63793 21536
0 21538 7 1 2 21510 21537
0 21539 5 1 1 21538
0 21540 7 1 2 21463 21539
0 21541 5 1 1 21540
0 21542 7 1 2 66462 21541
0 21543 5 1 1 21542
0 21544 7 5 2 81470 94679
0 21545 5 1 1 95201
0 21546 7 1 2 84012 95202
0 21547 5 1 1 21546
0 21548 7 1 2 88402 94849
0 21549 5 1 1 21548
0 21550 7 1 2 21547 21549
0 21551 5 1 1 21550
0 21552 7 1 2 94049 21551
0 21553 5 1 1 21552
0 21554 7 2 2 73849 90579
0 21555 7 1 2 94068 95145
0 21556 7 1 2 95206 21555
0 21557 5 1 1 21556
0 21558 7 1 2 21553 21557
0 21559 5 1 1 21558
0 21560 7 1 2 68639 21559
0 21561 5 1 1 21560
0 21562 7 1 2 78138 95146
0 21563 7 1 2 95207 21562
0 21564 5 1 1 21563
0 21565 7 1 2 21561 21564
0 21566 5 1 1 21565
0 21567 7 1 2 64114 21566
0 21568 5 1 1 21567
0 21569 7 4 2 67999 94850
0 21570 7 2 2 67676 95208
0 21571 5 1 1 95212
0 21572 7 1 2 21545 21571
0 21573 5 2 1 21572
0 21574 7 1 2 88138 95214
0 21575 5 1 1 21574
0 21576 7 3 2 68976 76733
0 21577 5 1 1 95216
0 21578 7 1 2 95209 95217
0 21579 5 1 1 21578
0 21580 7 1 2 21575 21579
0 21581 5 1 1 21580
0 21582 7 1 2 86627 21581
0 21583 5 1 1 21582
0 21584 7 1 2 21568 21583
0 21585 5 1 1 21584
0 21586 7 1 2 68399 21585
0 21587 5 1 1 21586
0 21588 7 1 2 73862 79205
0 21589 5 1 1 21588
0 21590 7 1 2 89380 77458
0 21591 5 1 1 21590
0 21592 7 1 2 21589 21591
0 21593 5 1 1 21592
0 21594 7 3 2 66946 63956
0 21595 5 1 1 95219
0 21596 7 1 2 80137 95220
0 21597 7 1 2 94745 21596
0 21598 7 1 2 21593 21597
0 21599 5 1 1 21598
0 21600 7 1 2 21587 21599
0 21601 5 1 1 21600
0 21602 7 1 2 66703 21601
0 21603 5 1 1 21602
0 21604 7 1 2 68400 73551
0 21605 5 1 1 21604
0 21606 7 1 2 112 21605
0 21607 5 1 1 21606
0 21608 7 1 2 71832 21607
0 21609 5 1 1 21608
0 21610 7 1 2 9189 21609
0 21611 5 1 1 21610
0 21612 7 1 2 63957 21611
0 21613 5 1 1 21612
0 21614 7 1 2 80069 75460
0 21615 5 1 1 21614
0 21616 7 1 2 21613 21615
0 21617 5 1 1 21616
0 21618 7 1 2 62086 21617
0 21619 5 1 1 21618
0 21620 7 1 2 77301 87573
0 21621 7 1 2 89626 21620
0 21622 5 1 1 21621
0 21623 7 1 2 21619 21622
0 21624 5 1 1 21623
0 21625 7 1 2 85101 80148
0 21626 7 1 2 95101 21625
0 21627 7 1 2 21624 21626
0 21628 5 1 1 21627
0 21629 7 1 2 21603 21628
0 21630 5 1 1 21629
0 21631 7 1 2 65136 21630
0 21632 5 1 1 21631
0 21633 7 1 2 71833 89072
0 21634 5 1 1 21633
0 21635 7 1 2 17525 21634
0 21636 5 1 1 21635
0 21637 7 1 2 77931 21636
0 21638 5 1 1 21637
0 21639 7 1 2 86261 80138
0 21640 7 1 2 75262 21639
0 21641 5 1 1 21640
0 21642 7 1 2 21638 21641
0 21643 5 1 1 21642
0 21644 7 1 2 77946 21643
0 21645 5 1 1 21644
0 21646 7 3 2 69555 87474
0 21647 7 1 2 77170 73810
0 21648 7 1 2 95222 21647
0 21649 5 1 1 21648
0 21650 7 1 2 21645 21649
0 21651 5 1 1 21650
0 21652 7 1 2 63958 21651
0 21653 5 1 1 21652
0 21654 7 3 2 62573 72143
0 21655 5 2 1 95225
0 21656 7 1 2 78926 95226
0 21657 5 2 1 21656
0 21658 7 1 2 80155 95230
0 21659 5 1 1 21658
0 21660 7 1 2 76633 21659
0 21661 5 1 1 21660
0 21662 7 1 2 80473 87131
0 21663 7 1 2 82929 21662
0 21664 5 1 1 21663
0 21665 7 1 2 21661 21664
0 21666 5 1 1 21665
0 21667 7 1 2 63555 21666
0 21668 5 1 1 21667
0 21669 7 1 2 21653 21668
0 21670 5 1 1 21669
0 21671 7 1 2 61851 21670
0 21672 5 1 1 21671
0 21673 7 3 2 75478 89965
0 21674 7 1 2 77171 87109
0 21675 7 1 2 95177 21674
0 21676 7 1 2 95232 21675
0 21677 5 1 1 21676
0 21678 7 1 2 21672 21677
0 21679 5 1 1 21678
0 21680 7 1 2 95128 21679
0 21681 5 1 1 21680
0 21682 7 1 2 61553 21681
0 21683 7 1 2 21632 21682
0 21684 5 1 1 21683
0 21685 7 1 2 21543 21684
0 21686 5 1 1 21685
0 21687 7 2 2 81894 73609
0 21688 7 1 2 86226 95235
0 21689 5 1 1 21688
0 21690 7 1 2 68640 75593
0 21691 7 1 2 90766 21690
0 21692 5 1 1 21691
0 21693 7 1 2 21689 21692
0 21694 5 1 1 21693
0 21695 7 1 2 94701 21694
0 21696 5 1 1 21695
0 21697 7 2 2 78756 80835
0 21698 7 1 2 89934 85102
0 21699 7 1 2 94851 21698
0 21700 7 1 2 95237 21699
0 21701 5 1 1 21700
0 21702 7 1 2 21696 21701
0 21703 5 1 1 21702
0 21704 7 1 2 70911 21703
0 21705 5 1 1 21704
0 21706 7 1 2 88841 77546
0 21707 7 1 2 84575 21706
0 21708 7 1 2 95210 21707
0 21709 5 1 1 21708
0 21710 7 1 2 21705 21709
0 21711 5 1 1 21710
0 21712 7 1 2 64115 21711
0 21713 5 1 1 21712
0 21714 7 1 2 89817 78263
0 21715 5 1 1 21714
0 21716 7 2 2 83767 89935
0 21717 7 1 2 73850 89283
0 21718 7 1 2 95239 21717
0 21719 5 1 1 21718
0 21720 7 1 2 21715 21719
0 21721 5 1 1 21720
0 21722 7 1 2 62402 21721
0 21723 5 1 1 21722
0 21724 7 3 2 69556 94232
0 21725 7 3 2 65414 84620
0 21726 5 1 1 95244
0 21727 7 1 2 77727 76286
0 21728 5 1 1 21727
0 21729 7 1 2 65979 21728
0 21730 7 2 2 95245 21729
0 21731 7 1 2 95241 95247
0 21732 5 1 1 21731
0 21733 7 1 2 21723 21732
0 21734 5 1 1 21733
0 21735 7 7 2 64510 80976
0 21736 7 8 2 94354 95249
0 21737 7 1 2 21734 95256
0 21738 5 1 1 21737
0 21739 7 1 2 21713 21738
0 21740 5 1 1 21739
0 21741 7 1 2 66947 21740
0 21742 5 1 1 21741
0 21743 7 1 2 79282 77211
0 21744 7 1 2 95119 21743
0 21745 5 1 1 21744
0 21746 7 3 2 82156 90231
0 21747 7 1 2 69557 74583
0 21748 7 1 2 95102 21747
0 21749 7 1 2 95264 21748
0 21750 5 1 1 21749
0 21751 7 1 2 21745 21750
0 21752 5 1 1 21751
0 21753 7 1 2 70912 21752
0 21754 5 1 1 21753
0 21755 7 2 2 62087 80209
0 21756 7 1 2 88842 95267
0 21757 7 1 2 95120 21756
0 21758 5 1 1 21757
0 21759 7 1 2 21754 21758
0 21760 5 1 1 21759
0 21761 7 1 2 64116 21760
0 21762 5 1 1 21761
0 21763 7 1 2 80210 87574
0 21764 7 1 2 90054 21763
0 21765 7 1 2 95121 21764
0 21766 5 1 1 21765
0 21767 7 1 2 21762 21766
0 21768 5 1 1 21767
0 21769 7 1 2 73444 21768
0 21770 5 1 1 21769
0 21771 7 3 2 64713 74155
0 21772 7 1 2 73851 75499
0 21773 5 1 1 21772
0 21774 7 1 2 18789 21773
0 21775 5 1 1 21774
0 21776 7 1 2 94702 21775
0 21777 5 1 1 21776
0 21778 7 2 2 80668 95185
0 21779 5 1 1 95272
0 21780 7 1 2 74532 75540
0 21781 7 1 2 95273 21780
0 21782 5 1 1 21781
0 21783 7 1 2 21777 21782
0 21784 5 1 1 21783
0 21785 7 1 2 64117 21784
0 21786 5 1 1 21785
0 21787 7 1 2 75324 93364
0 21788 7 4 2 63959 94355
0 21789 7 2 2 64511 73852
0 21790 7 1 2 95274 95278
0 21791 7 1 2 21787 21790
0 21792 5 1 1 21791
0 21793 7 1 2 21786 21792
0 21794 5 1 1 21793
0 21795 7 1 2 95269 21794
0 21796 5 1 1 21795
0 21797 7 1 2 21770 21796
0 21798 7 1 2 21742 21797
0 21799 5 1 1 21798
0 21800 7 1 2 94936 21799
0 21801 5 1 1 21800
0 21802 7 10 2 64118 69091
0 21803 7 1 2 82157 95280
0 21804 7 1 2 91892 21803
0 21805 7 1 2 95200 21804
0 21806 5 1 1 21805
0 21807 7 6 2 68977 93896
0 21808 7 2 2 69362 88767
0 21809 7 1 2 85205 95296
0 21810 7 1 2 95290 21809
0 21811 5 1 1 21810
0 21812 7 1 2 21806 21811
0 21813 5 1 1 21812
0 21814 7 1 2 62829 21813
0 21815 5 1 1 21814
0 21816 7 3 2 71327 84381
0 21817 7 7 2 64340 65137
0 21818 7 3 2 93732 95301
0 21819 7 11 2 68641 69092
0 21820 7 1 2 81652 95311
0 21821 7 1 2 95308 21820
0 21822 7 1 2 95298 21821
0 21823 5 1 1 21822
0 21824 7 1 2 21815 21823
0 21825 5 1 1 21824
0 21826 7 1 2 61554 21825
0 21827 5 1 1 21826
0 21828 7 1 2 89768 76669
0 21829 5 1 1 21828
0 21830 7 1 2 85206 84466
0 21831 5 1 1 21830
0 21832 7 1 2 21829 21831
0 21833 5 2 1 21832
0 21834 7 1 2 94722 95299
0 21835 7 1 2 95322 21834
0 21836 5 1 1 21835
0 21837 7 1 2 21827 21836
0 21838 5 1 1 21837
0 21839 7 1 2 64714 21838
0 21840 5 1 1 21839
0 21841 7 1 2 61555 95323
0 21842 5 1 1 21841
0 21843 7 1 2 88479 92538
0 21844 5 1 1 21843
0 21845 7 1 2 21842 21844
0 21846 5 1 1 21845
0 21847 7 1 2 88139 94746
0 21848 7 1 2 21846 21847
0 21849 5 1 1 21848
0 21850 7 1 2 21840 21849
0 21851 5 1 1 21850
0 21852 7 1 2 75144 21851
0 21853 5 1 1 21852
0 21854 7 2 2 70048 89496
0 21855 7 3 2 63556 77196
0 21856 7 1 2 95326 95211
0 21857 7 1 2 95324 21856
0 21858 5 1 1 21857
0 21859 7 1 2 79839 94481
0 21860 7 1 2 95203 21859
0 21861 5 1 1 21860
0 21862 7 1 2 21858 21861
0 21863 5 1 1 21862
0 21864 7 1 2 62088 80897
0 21865 5 1 1 21864
0 21866 7 1 2 83610 21865
0 21867 5 1 1 21866
0 21868 7 1 2 73445 21867
0 21869 7 1 2 21863 21868
0 21870 5 1 1 21869
0 21871 7 1 2 63319 21870
0 21872 7 1 2 21853 21871
0 21873 7 1 2 21801 21872
0 21874 7 1 2 21686 21873
0 21875 5 1 1 21874
0 21876 7 1 2 21361 21875
0 21877 5 1 1 21876
0 21878 7 4 2 68401 75574
0 21879 7 1 2 80875 95329
0 21880 5 1 1 21879
0 21881 7 1 2 89630 85668
0 21882 5 1 1 21881
0 21883 7 1 2 21880 21882
0 21884 5 1 1 21883
0 21885 7 1 2 73318 21884
0 21886 5 1 1 21885
0 21887 7 1 2 88610 90164
0 21888 5 1 1 21887
0 21889 7 1 2 21886 21888
0 21890 5 1 1 21889
0 21891 7 1 2 70334 21890
0 21892 5 2 1 21891
0 21893 7 1 2 81067 95072
0 21894 5 19 1 21893
0 21895 7 1 2 67443 86350
0 21896 5 1 1 21895
0 21897 7 1 2 65415 79478
0 21898 5 1 1 21897
0 21899 7 1 2 21896 21898
0 21900 5 1 1 21899
0 21901 7 1 2 95335 21900
0 21902 5 1 1 21901
0 21903 7 1 2 80571 87976
0 21904 5 1 1 21903
0 21905 7 1 2 21902 21904
0 21906 5 1 1 21905
0 21907 7 1 2 63147 21906
0 21908 5 1 1 21907
0 21909 7 1 2 95333 21908
0 21910 5 1 1 21909
0 21911 7 1 2 66463 21910
0 21912 5 1 1 21911
0 21913 7 2 2 65138 85691
0 21914 7 1 2 85063 95354
0 21915 5 1 1 21914
0 21916 7 1 2 78107 80898
0 21917 5 1 1 21916
0 21918 7 1 2 21915 21917
0 21919 5 1 1 21918
0 21920 7 1 2 66948 21919
0 21921 5 1 1 21920
0 21922 7 1 2 78413 85803
0 21923 5 1 1 21922
0 21924 7 1 2 21921 21923
0 21925 5 1 1 21924
0 21926 7 1 2 73446 21925
0 21927 5 1 1 21926
0 21928 7 1 2 70335 3548
0 21929 5 1 1 21928
0 21930 7 1 2 95071 21929
0 21931 5 1 1 21930
0 21932 7 1 2 75108 78414
0 21933 5 1 1 21932
0 21934 7 1 2 21931 21933
0 21935 5 1 1 21934
0 21936 7 1 2 85710 21935
0 21937 5 1 1 21936
0 21938 7 1 2 21927 21937
0 21939 5 1 1 21938
0 21940 7 1 2 76045 21939
0 21941 5 1 1 21940
0 21942 7 1 2 21912 21941
0 21943 5 1 1 21942
0 21944 7 1 2 72785 21943
0 21945 5 1 1 21944
0 21946 7 1 2 77661 86191
0 21947 7 1 2 95081 21946
0 21948 5 1 1 21947
0 21949 7 1 2 21945 21948
0 21950 5 1 1 21949
0 21951 7 1 2 94398 21950
0 21952 5 1 1 21951
0 21953 7 3 2 91278 94356
0 21954 7 1 2 74113 80031
0 21955 7 1 2 95356 21954
0 21956 7 1 2 93976 21955
0 21957 5 1 1 21956
0 21958 7 2 2 74272 93897
0 21959 7 2 2 70336 82938
0 21960 7 1 2 90030 95361
0 21961 7 1 2 95359 21960
0 21962 7 1 2 92329 21961
0 21963 5 1 1 21962
0 21964 7 1 2 21957 21963
0 21965 5 1 1 21964
0 21966 7 1 2 62089 21965
0 21967 5 1 1 21966
0 21968 7 1 2 80899 94937
0 21969 5 1 1 21968
0 21970 7 1 2 90111 21969
0 21971 5 1 1 21970
0 21972 7 1 2 73447 21971
0 21973 5 1 1 21972
0 21974 7 1 2 81052 77628
0 21975 5 1 1 21974
0 21976 7 1 2 90321 94938
0 21977 5 1 1 21976
0 21978 7 1 2 21975 21977
0 21979 5 1 1 21978
0 21980 7 1 2 68642 21979
0 21981 5 1 1 21980
0 21982 7 1 2 21973 21981
0 21983 5 1 1 21982
0 21984 7 1 2 74114 80947
0 21985 7 1 2 94399 21984
0 21986 7 1 2 21983 21985
0 21987 5 1 1 21986
0 21988 7 1 2 21967 21987
0 21989 5 1 1 21988
0 21990 7 1 2 61556 21989
0 21991 5 1 1 21990
0 21992 7 1 2 63148 93977
0 21993 7 1 2 95336 21992
0 21994 5 1 1 21993
0 21995 7 1 2 95334 21994
0 21996 5 1 1 21995
0 21997 7 1 2 74115 94723
0 21998 7 1 2 21996 21997
0 21999 5 1 1 21998
0 22000 7 1 2 21991 21999
0 22001 5 1 1 22000
0 22002 7 1 2 70913 22001
0 22003 5 1 1 22002
0 22004 7 1 2 64715 22003
0 22005 7 1 2 21952 22004
0 22006 5 1 1 22005
0 22007 7 1 2 77345 76615
0 22008 5 1 1 22007
0 22009 7 1 2 78302 22008
0 22010 5 1 1 22009
0 22011 7 1 2 74954 22010
0 22012 5 1 1 22011
0 22013 7 1 2 84165 88140
0 22014 5 1 1 22013
0 22015 7 1 2 22012 22014
0 22016 5 1 1 22015
0 22017 7 1 2 68643 22016
0 22018 5 1 1 22017
0 22019 7 4 2 72325 84013
0 22020 5 1 1 95363
0 22021 7 1 2 74945 95364
0 22022 5 1 1 22021
0 22023 7 1 2 22018 22022
0 22024 5 1 1 22023
0 22025 7 1 2 94703 22024
0 22026 5 1 1 22025
0 22027 7 6 2 67444 68978
0 22028 7 2 2 88621 95367
0 22029 7 3 2 68000 94357
0 22030 7 3 2 65980 87494
0 22031 7 1 2 95375 95378
0 22032 7 1 2 95373 22031
0 22033 5 1 1 22032
0 22034 7 3 2 91513 93898
0 22035 7 1 2 80332 95381
0 22036 7 1 2 83747 22035
0 22037 5 1 1 22036
0 22038 7 1 2 22033 22037
0 22039 5 1 1 22038
0 22040 7 1 2 76444 22039
0 22041 5 1 1 22040
0 22042 7 1 2 22026 22041
0 22043 5 1 1 22042
0 22044 7 1 2 70049 22043
0 22045 5 1 1 22044
0 22046 7 2 2 68402 75183
0 22047 7 1 2 87278 95384
0 22048 5 1 1 22047
0 22049 7 7 2 63557 71943
0 22050 5 1 1 95386
0 22051 7 6 2 66464 81517
0 22052 7 1 2 72750 95393
0 22053 7 1 2 95387 22052
0 22054 5 1 1 22053
0 22055 7 1 2 22048 22054
0 22056 5 1 1 22055
0 22057 7 1 2 86917 95109
0 22058 7 1 2 22056 22057
0 22059 5 1 1 22058
0 22060 7 1 2 22045 22059
0 22061 5 1 1 22060
0 22062 7 1 2 66949 22061
0 22063 5 1 1 22062
0 22064 7 1 2 71944 88622
0 22065 7 1 2 78213 22064
0 22066 7 2 2 74221 77471
0 22067 7 1 2 95357 95399
0 22068 7 1 2 22065 22067
0 22069 5 1 1 22068
0 22070 7 1 2 69558 22069
0 22071 7 1 2 22063 22070
0 22072 5 1 1 22071
0 22073 7 1 2 83115 22072
0 22074 7 1 2 22006 22073
0 22075 5 1 1 22074
0 22076 7 1 2 21877 22075
0 22077 5 1 1 22076
0 22078 7 1 2 70694 22077
0 22079 5 1 1 22078
0 22080 7 1 2 65416 94313
0 22081 5 2 1 22080
0 22082 7 1 2 72897 95401
0 22083 5 1 1 22082
0 22084 7 1 2 68644 22083
0 22085 5 1 1 22084
0 22086 7 1 2 94465 22085
0 22087 5 1 1 22086
0 22088 7 1 2 70050 22087
0 22089 5 1 1 22088
0 22090 7 2 2 74116 71709
0 22091 5 1 1 95403
0 22092 7 1 2 2263 22091
0 22093 5 1 1 22092
0 22094 7 1 2 82967 22093
0 22095 5 1 1 22094
0 22096 7 1 2 22089 22095
0 22097 5 1 1 22096
0 22098 7 1 2 75835 22097
0 22099 5 1 1 22098
0 22100 7 1 2 89764 93422
0 22101 5 1 1 22100
0 22102 7 2 2 77728 77346
0 22103 7 1 2 82052 95405
0 22104 5 1 1 22103
0 22105 7 7 2 77532 87147
0 22106 5 1 1 95407
0 22107 7 1 2 77743 95408
0 22108 5 1 1 22107
0 22109 7 1 2 22104 22108
0 22110 5 1 1 22109
0 22111 7 1 2 70051 22110
0 22112 5 1 1 22111
0 22113 7 1 2 85281 84014
0 22114 5 1 1 22113
0 22115 7 1 2 72898 22114
0 22116 5 1 1 22115
0 22117 7 1 2 68645 22116
0 22118 5 1 1 22117
0 22119 7 1 2 89790 22118
0 22120 5 1 1 22119
0 22121 7 1 2 76294 22120
0 22122 5 1 1 22121
0 22123 7 1 2 22112 22122
0 22124 5 1 1 22123
0 22125 7 1 2 75145 22124
0 22126 5 1 1 22125
0 22127 7 1 2 22101 22126
0 22128 7 1 2 22099 22127
0 22129 5 1 1 22128
0 22130 7 1 2 66465 22129
0 22131 5 1 1 22130
0 22132 7 5 2 71945 84114
0 22133 5 2 1 95414
0 22134 7 1 2 76295 95415
0 22135 5 1 1 22134
0 22136 7 1 2 70052 75836
0 22137 7 1 2 91427 22136
0 22138 5 1 1 22137
0 22139 7 1 2 22135 22138
0 22140 5 1 1 22139
0 22141 7 1 2 66466 22140
0 22142 5 1 1 22141
0 22143 7 1 2 81053 75954
0 22144 7 1 2 95265 22143
0 22145 5 1 1 22144
0 22146 7 1 2 22142 22145
0 22147 5 1 1 22146
0 22148 7 1 2 94558 22147
0 22149 5 1 1 22148
0 22150 7 2 2 78512 78415
0 22151 7 1 2 77472 89874
0 22152 7 1 2 95421 22151
0 22153 5 1 1 22152
0 22154 7 1 2 22149 22153
0 22155 7 1 2 22131 22154
0 22156 5 1 1 22155
0 22157 7 8 2 69093 64512
0 22158 7 1 2 68154 64341
0 22159 7 2 2 95423 22158
0 22160 7 1 2 22156 95431
0 22161 5 1 1 22160
0 22162 7 2 2 83290 94604
0 22163 7 1 2 81185 17914
0 22164 5 1 1 22163
0 22165 7 1 2 77443 22164
0 22166 5 1 1 22165
0 22167 7 1 2 78073 89303
0 22168 5 1 1 22167
0 22169 7 1 2 22166 22168
0 22170 5 1 1 22169
0 22171 7 1 2 95433 22170
0 22172 5 1 1 22171
0 22173 7 2 2 79738 94724
0 22174 7 1 2 72144 88607
0 22175 7 1 2 95435 22174
0 22176 5 1 1 22175
0 22177 7 1 2 22172 22176
0 22178 5 1 1 22177
0 22179 7 1 2 63794 22178
0 22180 5 1 1 22179
0 22181 7 2 2 76557 94400
0 22182 7 2 2 74803 95437
0 22183 7 1 2 86726 86740
0 22184 5 2 1 22183
0 22185 7 1 2 91693 95441
0 22186 7 1 2 95439 22185
0 22187 5 1 1 22186
0 22188 7 1 2 88762 90903
0 22189 7 8 2 68979 64250
0 22190 7 3 2 69187 95443
0 22191 7 1 2 81684 95451
0 22192 7 1 2 22188 22191
0 22193 5 1 1 22192
0 22194 7 1 2 22187 22193
0 22195 7 1 2 22180 22194
0 22196 5 1 1 22195
0 22197 7 1 2 67677 22196
0 22198 5 1 1 22197
0 22199 7 2 2 65139 86236
0 22200 5 1 1 95454
0 22201 7 1 2 95440 95455
0 22202 5 1 1 22201
0 22203 7 1 2 91124 87488
0 22204 7 1 2 95129 22203
0 22205 5 1 1 22204
0 22206 7 1 2 22202 22205
0 22207 5 1 1 22206
0 22208 7 1 2 63558 22207
0 22209 5 1 1 22208
0 22210 7 1 2 79579 86237
0 22211 5 1 1 22210
0 22212 7 1 2 77920 94116
0 22213 5 1 1 22212
0 22214 7 1 2 68646 22213
0 22215 7 1 2 22211 22214
0 22216 5 1 1 22215
0 22217 7 1 2 63795 22200
0 22218 5 1 1 22217
0 22219 7 1 2 95436 22218
0 22220 7 1 2 22216 22219
0 22221 5 1 1 22220
0 22222 7 1 2 22209 22221
0 22223 7 1 2 22198 22222
0 22224 5 1 1 22223
0 22225 7 1 2 62090 22224
0 22226 5 1 1 22225
0 22227 7 1 2 88557 74512
0 22228 7 2 2 74273 73162
0 22229 7 1 2 95130 95456
0 22230 7 1 2 22227 22229
0 22231 5 1 1 22230
0 22232 7 1 2 74886 79580
0 22233 7 1 2 89592 22232
0 22234 5 1 1 22233
0 22235 7 1 2 82218 22106
0 22236 5 1 1 22235
0 22237 7 1 2 75325 94117
0 22238 5 1 1 22237
0 22239 7 1 2 22236 22238
0 22240 5 1 1 22239
0 22241 7 1 2 94939 22240
0 22242 5 1 1 22241
0 22243 7 1 2 22234 22242
0 22244 5 1 1 22243
0 22245 7 4 2 66467 82621
0 22246 7 1 2 94401 95458
0 22247 7 1 2 22244 22246
0 22248 5 1 1 22247
0 22249 7 1 2 22231 22248
0 22250 7 1 2 22226 22249
0 22251 5 1 1 22250
0 22252 7 1 2 65417 22251
0 22253 5 1 1 22252
0 22254 7 1 2 74318 82968
0 22255 7 1 2 95409 22254
0 22256 5 1 1 22255
0 22257 7 1 2 91092 95337
0 22258 7 1 2 94561 22257
0 22259 5 1 1 22258
0 22260 7 1 2 22256 22259
0 22261 5 1 1 22260
0 22262 7 1 2 95438 22261
0 22263 5 1 1 22262
0 22264 7 1 2 74035 85833
0 22265 5 1 1 22264
0 22266 7 1 2 79622 77734
0 22267 5 1 1 22266
0 22268 7 1 2 62830 22267
0 22269 5 1 1 22268
0 22270 7 1 2 67678 10277
0 22271 5 1 1 22270
0 22272 7 1 2 63559 22271
0 22273 7 1 2 22269 22272
0 22274 5 1 1 22273
0 22275 7 1 2 22265 22274
0 22276 5 1 1 22275
0 22277 7 1 2 70337 22276
0 22278 5 1 1 22277
0 22279 7 1 2 84506 88085
0 22280 5 1 1 22279
0 22281 7 1 2 22278 22280
0 22282 5 1 1 22281
0 22283 7 1 2 62091 22282
0 22284 5 1 1 22283
0 22285 7 1 2 74274 72224
0 22286 7 1 2 93238 22285
0 22287 5 1 1 22286
0 22288 7 1 2 22284 22287
0 22289 5 1 1 22288
0 22290 7 1 2 95434 22289
0 22291 5 1 1 22290
0 22292 7 1 2 22263 22291
0 22293 7 1 2 22253 22292
0 22294 5 1 1 22293
0 22295 7 1 2 63320 22294
0 22296 5 1 1 22295
0 22297 7 1 2 22161 22296
0 22298 5 1 1 22297
0 22299 7 1 2 63149 22298
0 22300 5 1 1 22299
0 22301 7 1 2 87702 94996
0 22302 5 1 1 22301
0 22303 7 2 2 65140 83116
0 22304 7 3 2 68403 95462
0 22305 5 1 1 95464
0 22306 7 1 2 90232 95465
0 22307 5 1 1 22306
0 22308 7 1 2 22302 22307
0 22309 5 1 1 22308
0 22310 7 1 2 82180 22309
0 22311 5 1 1 22310
0 22312 7 1 2 62092 88633
0 22313 5 1 1 22312
0 22314 7 3 2 68155 90233
0 22315 7 1 2 94940 95467
0 22316 5 1 1 22315
0 22317 7 1 2 22313 22316
0 22318 5 1 1 22317
0 22319 7 1 2 61852 22318
0 22320 5 1 1 22319
0 22321 7 1 2 78513 94886
0 22322 5 1 1 22321
0 22323 7 1 2 22320 22322
0 22324 5 1 1 22323
0 22325 7 1 2 94248 22324
0 22326 5 1 1 22325
0 22327 7 1 2 22311 22326
0 22328 5 1 1 22327
0 22329 7 1 2 77492 22328
0 22330 5 1 1 22329
0 22331 7 1 2 66704 92699
0 22332 5 1 1 22331
0 22333 7 1 2 10622 22332
0 22334 5 2 1 22333
0 22335 7 3 2 73448 91428
0 22336 7 1 2 77523 95472
0 22337 5 1 1 22336
0 22338 7 1 2 75982 22337
0 22339 5 1 1 22338
0 22340 7 1 2 95470 22339
0 22341 5 1 1 22340
0 22342 7 1 2 63560 89961
0 22343 7 1 2 95406 22342
0 22344 5 1 1 22343
0 22345 7 1 2 22341 22344
0 22346 5 1 1 22345
0 22347 7 1 2 61557 22346
0 22348 5 1 1 22347
0 22349 7 4 2 68647 85379
0 22350 7 1 2 78017 90915
0 22351 7 1 2 95475 22350
0 22352 5 1 1 22351
0 22353 7 1 2 22348 22352
0 22354 5 1 1 22353
0 22355 7 1 2 70053 22354
0 22356 5 1 1 22355
0 22357 7 1 2 89587 95422
0 22358 5 1 1 22357
0 22359 7 4 2 64119 77197
0 22360 7 1 2 77798 90817
0 22361 7 1 2 95479 22360
0 22362 5 1 1 22361
0 22363 7 1 2 22358 22362
0 22364 5 1 1 22363
0 22365 7 1 2 63796 22364
0 22366 5 1 1 22365
0 22367 7 4 2 72827 73648
0 22368 7 2 2 93454 95483
0 22369 5 1 1 95487
0 22370 7 1 2 75983 22369
0 22371 5 1 1 22370
0 22372 7 1 2 94482 22371
0 22373 5 1 1 22372
0 22374 7 1 2 22366 22373
0 22375 5 1 1 22374
0 22376 7 1 2 63321 22375
0 22377 5 1 1 22376
0 22378 7 1 2 83050 90149
0 22379 7 1 2 95488 22378
0 22380 5 1 1 22379
0 22381 7 1 2 22377 22380
0 22382 5 1 1 22381
0 22383 7 1 2 75146 22382
0 22384 5 1 1 22383
0 22385 7 1 2 22356 22384
0 22386 7 1 2 22330 22385
0 22387 5 1 1 22386
0 22388 7 1 2 64513 22387
0 22389 5 1 1 22388
0 22390 7 1 2 88602 78416
0 22391 7 1 2 82823 92888
0 22392 7 1 2 22390 22391
0 22393 5 1 1 22392
0 22394 7 1 2 85140 74707
0 22395 5 1 1 22394
0 22396 7 2 2 65418 91694
0 22397 7 1 2 68648 78514
0 22398 7 1 2 95489 22397
0 22399 5 1 1 22398
0 22400 7 1 2 22395 22399
0 22401 5 1 1 22400
0 22402 7 1 2 67242 22401
0 22403 5 1 1 22402
0 22404 7 1 2 74541 93451
0 22405 5 1 1 22404
0 22406 7 1 2 22403 22405
0 22407 5 1 1 22406
0 22408 7 1 2 62093 22407
0 22409 5 1 1 22408
0 22410 7 1 2 93474 95266
0 22411 5 1 1 22410
0 22412 7 1 2 22409 22411
0 22413 5 1 1 22412
0 22414 7 1 2 63322 92953
0 22415 7 1 2 22413 22414
0 22416 5 1 1 22415
0 22417 7 1 2 22393 22416
0 22418 5 1 1 22417
0 22419 7 1 2 72145 22418
0 22420 5 1 1 22419
0 22421 7 3 2 81698 75769
0 22422 7 1 2 88217 95491
0 22423 5 1 1 22422
0 22424 7 3 2 66705 75873
0 22425 7 1 2 88546 89769
0 22426 7 1 2 95494 22425
0 22427 5 1 1 22426
0 22428 7 1 2 22423 22427
0 22429 5 1 1 22428
0 22430 7 1 2 66468 22429
0 22431 5 1 1 22430
0 22432 7 1 2 89997 93733
0 22433 7 1 2 94997 22432
0 22434 5 1 1 22433
0 22435 7 1 2 22431 22434
0 22436 5 1 1 22435
0 22437 7 1 2 67243 22436
0 22438 5 1 1 22437
0 22439 7 1 2 74542 85141
0 22440 7 1 2 95492 22439
0 22441 5 1 1 22440
0 22442 7 1 2 22438 22441
0 22443 5 1 1 22442
0 22444 7 1 2 86238 22443
0 22445 5 1 1 22444
0 22446 7 1 2 22420 22445
0 22447 7 1 2 22389 22446
0 22448 5 1 1 22447
0 22449 7 1 2 95376 22448
0 22450 5 1 1 22449
0 22451 7 1 2 64716 22450
0 22452 7 1 2 22300 22451
0 22453 5 1 1 22452
0 22454 7 2 2 67244 95368
0 22455 5 1 1 95497
0 22456 7 1 2 73577 93455
0 22457 5 1 1 22456
0 22458 7 1 2 22455 22457
0 22459 5 1 1 22458
0 22460 7 1 2 94704 22459
0 22461 5 1 1 22460
0 22462 7 4 2 61558 80115
0 22463 7 2 2 94605 95499
0 22464 5 1 1 95503
0 22465 7 4 2 92214 95281
0 22466 7 1 2 95394 95505
0 22467 5 1 1 22466
0 22468 7 1 2 22464 22467
0 22469 5 1 1 22468
0 22470 7 1 2 71946 85737
0 22471 7 1 2 22469 22470
0 22472 5 1 1 22471
0 22473 7 1 2 91206 95506
0 22474 5 1 1 22473
0 22475 7 2 2 80647 91389
0 22476 7 1 2 61559 95444
0 22477 7 1 2 95509 22476
0 22478 5 1 1 22477
0 22479 7 1 2 22474 22478
0 22480 5 1 1 22479
0 22481 7 1 2 85754 22480
0 22482 5 1 1 22481
0 22483 7 2 2 84764 95110
0 22484 7 1 2 80933 91893
0 22485 7 1 2 95511 22484
0 22486 5 1 1 22485
0 22487 7 1 2 22482 22486
0 22488 7 1 2 22472 22487
0 22489 7 1 2 22461 22488
0 22490 5 1 1 22489
0 22491 7 1 2 68404 22490
0 22492 5 1 1 22491
0 22493 7 1 2 84228 95291
0 22494 7 2 2 65981 80850
0 22495 7 2 2 77577 88637
0 22496 7 1 2 95513 95515
0 22497 7 1 2 22493 22496
0 22498 5 1 1 22497
0 22499 7 1 2 22492 22498
0 22500 5 1 1 22499
0 22501 7 1 2 89911 22500
0 22502 5 1 1 22501
0 22503 7 2 2 72700 86406
0 22504 5 2 1 95517
0 22505 7 1 2 80824 80836
0 22506 7 1 2 95518 22505
0 22507 5 1 1 22506
0 22508 7 2 2 62094 72146
0 22509 7 1 2 73449 95521
0 22510 7 1 2 89183 22509
0 22511 5 1 1 22510
0 22512 7 1 2 22507 22511
0 22513 5 1 1 22512
0 22514 7 1 2 81635 94606
0 22515 7 1 2 22513 22514
0 22516 5 1 1 22515
0 22517 7 1 2 22502 22516
0 22518 5 1 1 22517
0 22519 7 1 2 70054 22518
0 22520 5 1 1 22519
0 22521 7 2 2 89165 80948
0 22522 7 1 2 76575 81583
0 22523 7 1 2 84435 94358
0 22524 7 1 2 22522 22523
0 22525 7 1 2 95523 22524
0 22526 5 1 1 22525
0 22527 7 1 2 22520 22526
0 22528 5 1 1 22527
0 22529 7 1 2 85103 22528
0 22530 5 1 1 22529
0 22531 7 1 2 69559 22530
0 22532 7 2 2 82662 94607
0 22533 7 1 2 1814 91419
0 22534 5 1 1 22533
0 22535 7 1 2 78108 85527
0 22536 7 1 2 22534 22535
0 22537 5 1 1 22536
0 22538 7 1 2 68828 79026
0 22539 7 1 2 94246 22538
0 22540 5 1 1 22539
0 22541 7 1 2 22537 22540
0 22542 5 1 1 22541
0 22543 7 1 2 95525 22542
0 22544 5 1 1 22543
0 22545 7 1 2 68156 69094
0 22546 7 2 2 95309 22545
0 22547 7 1 2 87539 95527
0 22548 7 1 2 95442 22547
0 22549 5 1 1 22548
0 22550 7 1 2 22544 22549
0 22551 5 1 1 22550
0 22552 7 1 2 67679 22551
0 22553 5 1 1 22552
0 22554 7 2 2 65419 95312
0 22555 7 1 2 80090 92215
0 22556 7 2 2 95529 22555
0 22557 7 1 2 82562 95531
0 22558 7 1 2 86239 22557
0 22559 5 1 1 22558
0 22560 7 1 2 22553 22559
0 22561 5 1 1 22560
0 22562 7 1 2 66950 22561
0 22563 5 1 1 22562
0 22564 7 1 2 87469 93899
0 22565 7 1 2 83568 22564
0 22566 7 1 2 94019 22565
0 22567 7 1 2 94038 22566
0 22568 5 1 1 22567
0 22569 7 1 2 22563 22568
0 22570 5 1 1 22569
0 22571 7 1 2 61560 22570
0 22572 5 1 1 22571
0 22573 7 1 2 92436 95473
0 22574 5 1 1 22573
0 22575 7 1 2 94251 22574
0 22576 5 1 1 22575
0 22577 7 1 2 70055 22576
0 22578 5 1 1 22577
0 22579 7 1 2 79016 92432
0 22580 5 1 1 22579
0 22581 7 1 2 22578 22580
0 22582 5 1 1 22581
0 22583 7 1 2 94705 22582
0 22584 5 1 1 22583
0 22585 7 2 2 88417 73319
0 22586 5 1 1 95533
0 22587 7 1 2 70338 78246
0 22588 5 1 1 22587
0 22589 7 1 2 22586 22588
0 22590 5 1 1 22589
0 22591 7 1 2 72619 22590
0 22592 5 1 1 22591
0 22593 7 1 2 70914 75500
0 22594 5 1 1 22593
0 22595 7 1 2 72951 22594
0 22596 5 1 1 22595
0 22597 7 1 2 65420 22596
0 22598 5 1 1 22597
0 22599 7 1 2 84738 91429
0 22600 5 1 1 22599
0 22601 7 1 2 22598 22600
0 22602 5 1 1 22601
0 22603 7 1 2 84501 22602
0 22604 5 1 1 22603
0 22605 7 1 2 22592 22604
0 22606 5 1 1 22605
0 22607 7 1 2 95257 22606
0 22608 5 1 1 22607
0 22609 7 1 2 22584 22608
0 22610 5 1 1 22609
0 22611 7 1 2 92700 22610
0 22612 5 1 1 22611
0 22613 7 1 2 73450 89467
0 22614 5 1 1 22613
0 22615 7 1 2 71328 22614
0 22616 5 2 1 22615
0 22617 7 1 2 89166 95313
0 22618 7 1 2 95310 22617
0 22619 7 1 2 94913 22618
0 22620 7 1 2 95535 22619
0 22621 5 1 1 22620
0 22622 7 1 2 22612 22621
0 22623 7 1 2 22572 22622
0 22624 5 1 1 22623
0 22625 7 1 2 66706 22624
0 22626 5 1 1 22625
0 22627 7 1 2 74841 84743
0 22628 5 1 1 22627
0 22629 7 1 2 91093 22628
0 22630 5 1 1 22629
0 22631 7 2 2 73552 74491
0 22632 5 1 1 95537
0 22633 7 1 2 68649 95538
0 22634 5 1 1 22633
0 22635 7 1 2 22630 22634
0 22636 5 1 1 22635
0 22637 7 1 2 88267 22636
0 22638 5 1 1 22637
0 22639 7 1 2 72620 86444
0 22640 5 1 1 22639
0 22641 7 1 2 70339 84739
0 22642 5 1 1 22641
0 22643 7 1 2 22632 22642
0 22644 5 1 1 22643
0 22645 7 1 2 64120 22644
0 22646 5 1 1 22645
0 22647 7 1 2 22640 22646
0 22648 5 1 1 22647
0 22649 7 1 2 68650 22648
0 22650 5 1 1 22649
0 22651 7 1 2 85037 84744
0 22652 5 1 1 22651
0 22653 7 1 2 64121 90375
0 22654 7 1 2 22652 22653
0 22655 5 1 1 22654
0 22656 7 1 2 22650 22655
0 22657 5 1 1 22656
0 22658 7 1 2 81449 22657
0 22659 5 1 1 22658
0 22660 7 1 2 22638 22659
0 22661 5 1 1 22660
0 22662 7 1 2 95258 22661
0 22663 5 1 1 22662
0 22664 7 2 2 72147 91430
0 22665 7 1 2 73451 95539
0 22666 5 1 1 22665
0 22667 7 1 2 72899 94243
0 22668 5 1 1 22667
0 22669 7 1 2 68651 22668
0 22670 5 1 1 22669
0 22671 7 1 2 94466 22670
0 22672 7 1 2 22666 22671
0 22673 5 1 1 22672
0 22674 7 1 2 81450 94706
0 22675 7 1 2 22673 22674
0 22676 5 1 1 22675
0 22677 7 1 2 65141 22676
0 22678 7 1 2 22663 22677
0 22679 5 1 1 22678
0 22680 7 1 2 71710 94707
0 22681 5 1 1 22680
0 22682 7 1 2 21779 22681
0 22683 5 1 1 22682
0 22684 7 1 2 64122 22683
0 22685 5 1 1 22684
0 22686 7 3 2 62574 95181
0 22687 7 5 2 64342 70915
0 22688 7 1 2 95250 95544
0 22689 7 1 2 95541 22688
0 22690 5 1 1 22689
0 22691 7 1 2 22685 22690
0 22692 5 1 1 22691
0 22693 7 1 2 71780 82267
0 22694 7 1 2 22692 22693
0 22695 5 1 1 22694
0 22696 7 1 2 89134 73963
0 22697 7 1 2 79212 22696
0 22698 5 1 1 22697
0 22699 7 1 2 66707 84588
0 22700 7 2 2 86763 80851
0 22701 7 1 2 92437 95549
0 22702 7 1 2 22699 22701
0 22703 5 1 1 22702
0 22704 7 1 2 22698 22703
0 22705 5 1 1 22704
0 22706 7 1 2 94608 22705
0 22707 5 1 1 22706
0 22708 7 1 2 76558 95532
0 22709 7 1 2 95536 22708
0 22710 5 1 1 22709
0 22711 7 1 2 22707 22710
0 22712 5 1 1 22711
0 22713 7 1 2 63323 22712
0 22714 5 1 1 22713
0 22715 7 1 2 70056 22714
0 22716 7 1 2 22695 22715
0 22717 5 1 1 22716
0 22718 7 1 2 75147 22717
0 22719 7 1 2 22679 22718
0 22720 5 1 1 22719
0 22721 7 1 2 22626 22720
0 22722 7 1 2 22531 22721
0 22723 5 1 1 22722
0 22724 7 1 2 65738 22723
0 22725 7 1 2 22453 22724
0 22726 5 1 1 22725
0 22727 7 3 2 80934 94852
0 22728 5 1 1 95551
0 22729 7 1 2 95338 95552
0 22730 5 1 1 22729
0 22731 7 2 2 64251 90290
0 22732 7 1 2 82807 95125
0 22733 7 1 2 95554 22732
0 22734 5 1 1 22733
0 22735 7 1 2 22730 22734
0 22736 5 1 1 22735
0 22737 7 1 2 72148 22736
0 22738 5 1 1 22737
0 22739 7 3 2 65982 95339
0 22740 7 1 2 89361 94853
0 22741 7 1 2 95556 22740
0 22742 5 1 1 22741
0 22743 7 1 2 22738 22742
0 22744 5 1 1 22743
0 22745 7 1 2 63150 22744
0 22746 5 1 1 22745
0 22747 7 1 2 93436 94597
0 22748 7 1 2 95557 22747
0 22749 5 1 1 22748
0 22750 7 1 2 22746 22749
0 22751 5 1 1 22750
0 22752 7 1 2 68829 22751
0 22753 5 1 1 22752
0 22754 7 2 2 66951 80049
0 22755 7 1 2 89353 95559
0 22756 7 1 2 95504 22755
0 22757 5 1 1 22756
0 22758 7 1 2 22753 22757
0 22759 5 1 1 22758
0 22760 7 1 2 67445 22759
0 22761 5 1 1 22760
0 22762 7 2 2 61561 75874
0 22763 7 1 2 78109 86407
0 22764 7 1 2 95561 22763
0 22765 7 1 2 95204 22764
0 22766 5 1 1 22765
0 22767 7 1 2 22761 22766
0 22768 5 1 1 22767
0 22769 7 1 2 71947 22768
0 22770 5 1 1 22769
0 22771 7 1 2 84451 78697
0 22772 7 1 2 90013 22771
0 22773 7 5 2 79444 93900
0 22774 7 2 2 80474 77302
0 22775 7 1 2 95563 95568
0 22776 7 1 2 22772 22775
0 22777 5 1 1 22776
0 22778 7 1 2 22770 22777
0 22779 5 1 1 22778
0 22780 7 1 2 70340 22779
0 22781 5 1 1 22780
0 22782 7 1 2 68830 74434
0 22783 7 2 2 81518 22782
0 22784 7 2 2 79969 89167
0 22785 5 1 1 95572
0 22786 7 1 2 95570 95573
0 22787 5 1 1 22786
0 22788 7 1 2 85821 85221
0 22789 5 2 1 22788
0 22790 7 1 2 81257 93330
0 22791 7 1 2 95574 22790
0 22792 5 1 1 22791
0 22793 7 1 2 22787 22792
0 22794 5 1 1 22793
0 22795 7 1 2 66952 22794
0 22796 5 1 1 22795
0 22797 7 1 2 74222 83456
0 22798 7 1 2 80463 22797
0 22799 7 1 2 88077 22798
0 22800 5 1 1 22799
0 22801 7 1 2 22796 22800
0 22802 5 1 1 22801
0 22803 7 1 2 94402 22802
0 22804 5 1 1 22803
0 22805 7 1 2 82219 93331
0 22806 7 2 2 80139 90234
0 22807 7 1 2 94747 95576
0 22808 7 1 2 22805 22807
0 22809 5 1 1 22808
0 22810 7 1 2 22804 22809
0 22811 5 1 1 22810
0 22812 7 1 2 68980 22811
0 22813 5 1 1 22812
0 22814 7 2 2 86764 74887
0 22815 7 1 2 90580 94772
0 22816 7 1 2 95578 22815
0 22817 5 1 1 22816
0 22818 7 1 2 21355 22728
0 22819 5 2 1 22818
0 22820 7 1 2 77735 91652
0 22821 7 1 2 95580 22820
0 22822 5 1 1 22821
0 22823 7 1 2 22817 22822
0 22824 5 1 1 22823
0 22825 7 1 2 63151 22824
0 22826 5 1 1 22825
0 22827 7 1 2 86953 75326
0 22828 7 1 2 91788 22827
0 22829 7 1 2 95186 22828
0 22830 5 1 1 22829
0 22831 7 1 2 22826 22830
0 22832 5 1 1 22831
0 22833 7 1 2 66953 22832
0 22834 5 1 1 22833
0 22835 7 1 2 68652 94764
0 22836 7 1 2 90581 22835
0 22837 7 2 2 67446 80743
0 22838 7 1 2 86771 95582
0 22839 7 1 2 22836 22838
0 22840 5 1 1 22839
0 22841 7 1 2 22834 22840
0 22842 7 1 2 22813 22841
0 22843 5 1 1 22842
0 22844 7 1 2 72149 22843
0 22845 5 1 1 22844
0 22846 7 1 2 89569 91779
0 22847 7 1 2 91789 22846
0 22848 7 1 2 94622 22847
0 22849 5 1 1 22848
0 22850 7 1 2 22845 22849
0 22851 5 1 1 22850
0 22852 7 1 2 76893 22851
0 22853 5 1 1 22852
0 22854 7 1 2 22781 22853
0 22855 5 1 1 22854
0 22856 7 1 2 83117 22855
0 22857 5 1 1 22856
0 22858 7 3 2 73320 94209
0 22859 5 3 1 95584
0 22860 7 1 2 61562 95215
0 22861 5 1 1 22860
0 22862 7 1 2 83510 94854
0 22863 5 1 1 22862
0 22864 7 1 2 22861 22863
0 22865 5 1 1 22864
0 22866 7 1 2 95585 22865
0 22867 5 1 1 22866
0 22868 7 1 2 91431 95093
0 22869 5 1 1 22868
0 22870 7 1 2 73988 95553
0 22871 5 1 1 22870
0 22872 7 1 2 22869 22871
0 22873 5 1 1 22872
0 22874 7 1 2 74400 80605
0 22875 7 1 2 22873 22874
0 22876 5 1 1 22875
0 22877 7 1 2 22867 22876
0 22878 5 1 1 22877
0 22879 7 1 2 72150 22878
0 22880 5 1 1 22879
0 22881 7 4 2 88733 94359
0 22882 7 1 2 74401 80888
0 22883 5 2 1 22882
0 22884 7 1 2 95587 95594
0 22885 5 1 1 22884
0 22886 7 1 2 81258 22885
0 22887 5 1 1 22886
0 22888 7 5 2 66469 86924
0 22889 5 1 1 95596
0 22890 7 1 2 68001 95597
0 22891 7 1 2 95586 22890
0 22892 5 1 1 22891
0 22893 7 1 2 22887 22892
0 22894 5 1 1 22893
0 22895 7 1 2 68981 22894
0 22896 5 1 1 22895
0 22897 7 1 2 87013 15966
0 22898 5 2 1 22897
0 22899 7 1 2 73989 95601
0 22900 7 1 2 95571 22899
0 22901 5 1 1 22900
0 22902 7 1 2 22896 22901
0 22903 5 1 1 22902
0 22904 7 1 2 95590 22903
0 22905 5 1 1 22904
0 22906 7 1 2 22880 22905
0 22907 5 1 1 22906
0 22908 7 1 2 63324 22907
0 22909 5 1 1 22908
0 22910 7 1 2 89561 91943
0 22911 5 1 1 22910
0 22912 7 1 2 64717 89559
0 22913 5 1 1 22912
0 22914 7 1 2 22911 22913
0 22915 5 1 1 22914
0 22916 7 1 2 65421 94360
0 22917 7 1 2 91958 22916
0 22918 7 1 2 22915 22917
0 22919 5 1 1 22918
0 22920 7 1 2 22909 22919
0 22921 5 1 1 22920
0 22922 7 1 2 66708 22921
0 22923 5 1 1 22922
0 22924 7 1 2 76147 77524
0 22925 5 1 1 22924
0 22926 7 1 2 80935 80116
0 22927 5 1 1 22926
0 22928 7 1 2 22925 22927
0 22929 5 2 1 22928
0 22930 7 1 2 94755 95530
0 22931 7 2 2 95603 22930
0 22932 7 1 2 81680 89721
0 22933 7 1 2 95605 22932
0 22934 5 1 1 22933
0 22935 7 1 2 22923 22934
0 22936 5 1 1 22935
0 22937 7 1 2 65142 22936
0 22938 5 1 1 22937
0 22939 7 1 2 84605 95205
0 22940 5 1 1 22939
0 22941 7 1 2 73321 95213
0 22942 5 1 1 22941
0 22943 7 1 2 22940 22942
0 22944 5 1 1 22943
0 22945 7 1 2 66470 22944
0 22946 5 1 1 22945
0 22947 7 3 2 63960 78757
0 22948 7 1 2 95094 95607
0 22949 5 1 1 22948
0 22950 7 1 2 22946 22949
0 22951 5 1 1 22950
0 22952 7 1 2 72151 22951
0 22953 5 1 1 22952
0 22954 7 1 2 80669 95591
0 22955 5 1 1 22954
0 22956 7 1 2 92096 94609
0 22957 5 1 1 22956
0 22958 7 1 2 22955 22957
0 22959 5 1 1 22958
0 22960 7 1 2 63961 80165
0 22961 7 1 2 22959 22960
0 22962 5 1 1 22961
0 22963 7 1 2 22953 22962
0 22964 5 1 1 22963
0 22965 7 2 2 74275 83678
0 22966 7 1 2 76762 95610
0 22967 7 1 2 22964 22966
0 22968 5 1 1 22967
0 22969 7 1 2 22938 22968
0 22970 5 1 1 22969
0 22971 7 1 2 66954 22970
0 22972 5 1 1 22971
0 22973 7 2 2 68002 82158
0 22974 7 1 2 84969 95111
0 22975 7 1 2 95612 22974
0 22976 7 1 2 88317 22975
0 22977 5 1 1 22976
0 22978 7 2 2 62831 84015
0 22979 5 1 1 95614
0 22980 7 1 2 151 22979
0 22981 5 1 1 22980
0 22982 7 1 2 62403 22981
0 22983 5 1 1 22982
0 22984 7 1 2 73553 72888
0 22985 5 1 1 22984
0 22986 7 1 2 22983 22985
0 22987 5 1 1 22986
0 22988 7 1 2 64123 22987
0 22989 5 1 1 22988
0 22990 7 2 2 62404 72411
0 22991 5 1 1 95616
0 22992 7 1 2 22989 22991
0 22993 5 1 1 22992
0 22994 7 1 2 88768 94789
0 22995 7 1 2 22993 22994
0 22996 5 1 1 22995
0 22997 7 1 2 22977 22996
0 22998 5 1 1 22997
0 22999 7 1 2 63325 22998
0 23000 5 1 1 22999
0 23001 7 2 2 89562 95275
0 23002 7 1 2 88797 92304
0 23003 7 1 2 95618 23002
0 23004 5 1 1 23003
0 23005 7 1 2 23000 23004
0 23006 5 1 1 23005
0 23007 7 1 2 61563 23006
0 23008 5 1 1 23007
0 23009 7 5 2 67447 72374
0 23010 5 2 1 95620
0 23011 7 1 2 87295 95621
0 23012 5 2 1 23011
0 23013 7 1 2 18551 95627
0 23014 5 1 1 23013
0 23015 7 1 2 76559 95191
0 23016 7 1 2 89516 23015
0 23017 7 1 2 23014 23016
0 23018 5 1 1 23017
0 23019 7 1 2 23008 23018
0 23020 5 1 1 23019
0 23021 7 1 2 64718 23020
0 23022 5 1 1 23021
0 23023 7 3 2 87853 95424
0 23024 7 1 2 80977 87296
0 23025 7 1 2 95629 23024
0 23026 7 1 2 72844 23025
0 23027 5 1 1 23026
0 23028 7 1 2 72152 94708
0 23029 5 2 1 23028
0 23030 7 1 2 67680 95632
0 23031 5 1 1 23030
0 23032 7 1 2 90528 95592
0 23033 5 1 1 23032
0 23034 7 2 2 95633 23033
0 23035 5 1 1 95634
0 23036 7 1 2 93991 23035
0 23037 7 1 2 23031 23036
0 23038 5 1 1 23037
0 23039 7 1 2 23027 23038
0 23040 5 1 1 23039
0 23041 7 1 2 78264 23040
0 23042 5 1 1 23041
0 23043 7 1 2 23022 23042
0 23044 5 1 1 23043
0 23045 7 1 2 63561 23044
0 23046 5 1 1 23045
0 23047 7 2 2 72828 93432
0 23048 7 1 2 81920 95636
0 23049 5 1 1 23048
0 23050 7 1 2 93434 23049
0 23051 5 1 1 23050
0 23052 7 1 2 65983 23051
0 23053 5 1 1 23052
0 23054 7 1 2 72621 89358
0 23055 5 1 1 23054
0 23056 7 1 2 23053 23055
0 23057 5 1 1 23056
0 23058 7 1 2 83051 89979
0 23059 7 1 2 23057 23058
0 23060 5 1 1 23059
0 23061 7 1 2 90357 87075
0 23062 7 1 2 92134 23061
0 23063 5 1 1 23062
0 23064 7 1 2 23060 23063
0 23065 5 1 1 23064
0 23066 7 1 2 68653 23065
0 23067 5 1 1 23066
0 23068 7 1 2 90091 88156
0 23069 7 1 2 92341 23068
0 23070 5 1 1 23069
0 23071 7 1 2 23067 23070
0 23072 5 1 1 23071
0 23073 7 1 2 80032 94403
0 23074 7 1 2 23072 23073
0 23075 5 1 1 23074
0 23076 7 1 2 23046 23075
0 23077 5 1 1 23076
0 23078 7 1 2 80572 23077
0 23079 5 1 1 23078
0 23080 7 2 2 83332 91514
0 23081 7 4 2 64124 64252
0 23082 7 1 2 94783 95640
0 23083 7 1 2 90483 23082
0 23084 7 1 2 95638 23083
0 23085 5 1 1 23084
0 23086 7 4 2 64343 65422
0 23087 7 1 2 80805 95644
0 23088 7 1 2 85883 23087
0 23089 7 2 2 68982 69095
0 23090 7 3 2 68831 95648
0 23091 7 1 2 87459 95650
0 23092 7 1 2 23088 23091
0 23093 5 1 1 23092
0 23094 7 1 2 23085 23093
0 23095 5 1 1 23094
0 23096 7 1 2 63562 23095
0 23097 5 1 1 23096
0 23098 7 2 2 61564 81519
0 23099 7 1 2 93352 95653
0 23100 5 1 1 23099
0 23101 7 1 2 10733 2935
0 23102 5 1 1 23101
0 23103 7 1 2 72153 77736
0 23104 7 1 2 23102 23103
0 23105 5 1 1 23104
0 23106 7 1 2 23100 23105
0 23107 5 1 1 23106
0 23108 7 2 2 65423 79739
0 23109 7 1 2 94855 95655
0 23110 7 1 2 23107 23109
0 23111 5 1 1 23110
0 23112 7 1 2 23097 23111
0 23113 5 1 1 23112
0 23114 7 1 2 67681 23113
0 23115 5 1 1 23114
0 23116 7 1 2 71948 94748
0 23117 7 4 2 70341 72154
0 23118 7 4 2 82307 80606
0 23119 7 1 2 95657 95661
0 23120 7 1 2 23116 23119
0 23121 5 1 1 23120
0 23122 7 5 2 69560 72155
0 23123 7 1 2 95103 95665
0 23124 5 1 1 23123
0 23125 7 1 2 20147 23124
0 23126 5 1 1 23125
0 23127 7 1 2 61565 23126
0 23128 5 1 1 23127
0 23129 7 2 2 68983 76083
0 23130 5 1 1 95670
0 23131 7 1 2 94623 95671
0 23132 5 1 1 23131
0 23133 7 1 2 23128 23132
0 23134 5 1 1 23133
0 23135 7 1 2 77737 95246
0 23136 7 1 2 23134 23135
0 23137 5 1 1 23136
0 23138 7 1 2 23121 23137
0 23139 5 1 1 23138
0 23140 7 1 2 68405 23139
0 23141 5 1 1 23140
0 23142 7 1 2 94765 95579
0 23143 7 1 2 95510 23142
0 23144 7 1 2 95223 23143
0 23145 5 1 1 23144
0 23146 7 1 2 23141 23145
0 23147 5 1 1 23146
0 23148 7 1 2 66709 23147
0 23149 5 1 1 23148
0 23150 7 1 2 23115 23149
0 23151 5 1 1 23150
0 23152 7 1 2 63326 23151
0 23153 5 1 1 23152
0 23154 7 1 2 83052 76402
0 23155 7 1 2 95606 23154
0 23156 5 1 1 23155
0 23157 7 1 2 65143 23156
0 23158 7 1 2 23153 23157
0 23159 5 1 1 23158
0 23160 7 1 2 84216 95112
0 23161 7 1 2 95604 23160
0 23162 5 1 1 23161
0 23163 7 1 2 85421 85917
0 23164 7 1 2 94598 23163
0 23165 7 1 2 89517 23164
0 23166 5 1 1 23165
0 23167 7 1 2 23162 23166
0 23168 5 1 1 23167
0 23169 7 1 2 64719 23168
0 23170 5 1 1 23169
0 23171 7 1 2 82765 95512
0 23172 5 1 1 23171
0 23173 7 1 2 72156 94610
0 23174 7 1 2 91305 23173
0 23175 5 2 1 23174
0 23176 7 1 2 23172 95672
0 23177 5 1 1 23176
0 23178 7 1 2 92570 23177
0 23179 5 1 1 23178
0 23180 7 1 2 23170 23179
0 23181 5 1 1 23180
0 23182 7 1 2 91432 23181
0 23183 5 1 1 23182
0 23184 7 1 2 71949 74752
0 23185 5 1 1 23184
0 23186 7 1 2 90385 87999
0 23187 7 1 2 23185 23186
0 23188 5 1 1 23187
0 23189 7 1 2 89346 94709
0 23190 7 1 2 23188 23189
0 23191 5 1 1 23190
0 23192 7 1 2 23183 23191
0 23193 5 1 1 23192
0 23194 7 1 2 68832 23193
0 23195 5 1 1 23194
0 23196 7 3 2 78758 82739
0 23197 7 1 2 75289 95113
0 23198 7 1 2 95674 23197
0 23199 5 1 1 23198
0 23200 7 2 2 63327 64253
0 23201 7 2 2 87823 95677
0 23202 7 1 2 71329 95297
0 23203 7 1 2 95679 23202
0 23204 5 1 1 23203
0 23205 7 1 2 23199 23204
0 23206 5 1 1 23205
0 23207 7 5 2 61566 80234
0 23208 5 4 1 95681
0 23209 7 1 2 20963 95686
0 23210 5 1 1 23209
0 23211 7 1 2 23206 23210
0 23212 5 1 1 23211
0 23213 7 1 2 90190 95581
0 23214 5 1 1 23213
0 23215 7 1 2 91296 94749
0 23216 5 1 1 23215
0 23217 7 1 2 23214 23216
0 23218 5 1 1 23217
0 23219 7 1 2 72157 23218
0 23220 5 1 1 23219
0 23221 7 1 2 76046 72829
0 23222 5 2 1 23221
0 23223 7 1 2 23130 95690
0 23224 5 1 1 23223
0 23225 7 1 2 82740 23224
0 23226 5 1 1 23225
0 23227 7 1 2 89362 85325
0 23228 5 1 1 23227
0 23229 7 1 2 23226 23228
0 23230 5 1 1 23229
0 23231 7 1 2 94624 23230
0 23232 5 1 1 23231
0 23233 7 1 2 23220 23232
0 23234 5 1 1 23233
0 23235 7 1 2 73322 23234
0 23236 5 1 1 23235
0 23237 7 1 2 23212 23236
0 23238 5 1 1 23237
0 23239 7 1 2 75955 23238
0 23240 5 1 1 23239
0 23241 7 1 2 63563 23240
0 23242 7 1 2 23195 23241
0 23243 5 1 1 23242
0 23244 7 2 2 62405 70994
0 23245 7 1 2 81815 95692
0 23246 7 1 2 95619 23245
0 23247 5 1 1 23246
0 23248 7 1 2 71167 77615
0 23249 5 1 1 23248
0 23250 7 1 2 70342 89610
0 23251 5 1 1 23250
0 23252 7 1 2 23249 23251
0 23253 5 1 1 23252
0 23254 7 1 2 88769 94688
0 23255 7 1 2 23253 23254
0 23256 5 1 1 23255
0 23257 7 1 2 23247 23256
0 23258 5 1 1 23257
0 23259 7 1 2 61567 23258
0 23260 5 1 1 23259
0 23261 7 1 2 80728 95114
0 23262 7 1 2 90191 23261
0 23263 7 1 2 94165 23262
0 23264 5 1 1 23263
0 23265 7 1 2 23260 23264
0 23266 5 1 1 23265
0 23267 7 1 2 64720 23266
0 23268 5 1 1 23267
0 23269 7 1 2 72545 95115
0 23270 7 1 2 91711 23269
0 23271 5 1 1 23270
0 23272 7 1 2 95673 23271
0 23273 5 1 1 23272
0 23274 7 1 2 73323 90221
0 23275 7 1 2 23273 23274
0 23276 5 1 1 23275
0 23277 7 1 2 23268 23276
0 23278 5 1 1 23277
0 23279 7 1 2 63797 23278
0 23280 5 1 1 23279
0 23281 7 1 2 77525 91973
0 23282 5 1 1 23281
0 23283 7 1 2 74076 81259
0 23284 5 1 1 23283
0 23285 7 1 2 23282 23284
0 23286 5 1 1 23285
0 23287 7 2 2 82140 82159
0 23288 7 1 2 94404 95622
0 23289 7 1 2 95694 23288
0 23290 7 1 2 23286 23289
0 23291 5 1 1 23290
0 23292 7 1 2 68406 23291
0 23293 7 1 2 23280 23292
0 23294 5 1 1 23293
0 23295 7 1 2 23243 23294
0 23296 5 1 1 23295
0 23297 7 1 2 70057 23296
0 23298 5 1 1 23297
0 23299 7 1 2 62095 23298
0 23300 7 1 2 23159 23299
0 23301 5 1 1 23300
0 23302 7 1 2 23079 23301
0 23303 7 1 2 22972 23302
0 23304 7 1 2 22857 23303
0 23305 7 1 2 22726 23304
0 23306 7 1 2 22079 23305
0 23307 5 1 1 23306
0 23308 7 1 2 64923 23307
0 23309 5 1 1 23308
0 23310 7 1 2 21212 23309
0 23311 7 1 2 20620 23310
0 23312 5 1 1 23311
0 23313 7 1 2 93848 23312
0 23314 5 1 1 23313
0 23315 7 2 2 67245 76343
0 23316 7 1 2 73685 95696
0 23317 5 2 1 23316
0 23318 7 1 2 71950 94118
0 23319 5 2 1 23318
0 23320 7 1 2 779 95700
0 23321 5 2 1 23320
0 23322 7 1 2 68407 95702
0 23323 5 1 1 23322
0 23324 7 1 2 95698 23323
0 23325 5 1 1 23324
0 23326 7 1 2 88203 23325
0 23327 5 1 1 23326
0 23328 7 3 2 84374 78311
0 23329 5 10 1 95704
0 23330 7 2 2 68408 95707
0 23331 5 1 1 95717
0 23332 7 1 2 72546 77870
0 23333 7 1 2 75436 23332
0 23334 5 1 1 23333
0 23335 7 1 2 23331 23334
0 23336 5 1 1 23335
0 23337 7 1 2 67246 23336
0 23338 5 2 1 23337
0 23339 7 1 2 73913 94119
0 23340 5 1 1 23339
0 23341 7 1 2 95719 23340
0 23342 5 1 1 23341
0 23343 7 1 2 65144 23342
0 23344 5 1 1 23343
0 23345 7 1 2 70058 88506
0 23346 7 1 2 72880 23345
0 23347 5 1 1 23346
0 23348 7 2 2 63328 23347
0 23349 7 1 2 23344 95721
0 23350 5 1 1 23349
0 23351 7 1 2 88328 77275
0 23352 5 2 1 23351
0 23353 7 1 2 67247 76521
0 23354 5 2 1 23353
0 23355 7 1 2 71951 77493
0 23356 5 1 1 23355
0 23357 7 1 2 95725 23356
0 23358 5 1 1 23357
0 23359 7 1 2 78074 23358
0 23360 5 1 1 23359
0 23361 7 1 2 68157 23360
0 23362 7 1 2 95723 23361
0 23363 5 1 1 23362
0 23364 7 1 2 66710 23363
0 23365 7 1 2 23350 23364
0 23366 5 1 1 23365
0 23367 7 1 2 23327 23366
0 23368 5 1 1 23367
0 23369 7 1 2 64924 23368
0 23370 5 1 1 23369
0 23371 7 1 2 73881 81171
0 23372 5 2 1 23371
0 23373 7 1 2 68409 95727
0 23374 5 1 1 23373
0 23375 7 2 2 73554 71525
0 23376 5 1 1 95729
0 23377 7 1 2 87229 95730
0 23378 5 1 1 23377
0 23379 7 1 2 23374 23378
0 23380 5 1 1 23379
0 23381 7 1 2 71432 89108
0 23382 7 1 2 23380 23381
0 23383 5 2 1 23382
0 23384 7 1 2 23370 95731
0 23385 5 1 1 23384
0 23386 7 1 2 62096 23385
0 23387 5 1 1 23386
0 23388 7 1 2 82717 72326
0 23389 7 2 2 66711 79223
0 23390 7 3 2 77817 81357
0 23391 7 1 2 95733 95735
0 23392 7 1 2 23388 23391
0 23393 5 1 1 23392
0 23394 7 1 2 23387 23393
0 23395 5 1 1 23394
0 23396 7 1 2 61568 23395
0 23397 5 1 1 23396
0 23398 7 1 2 70059 74513
0 23399 5 1 1 23398
0 23400 7 1 2 81186 23399
0 23401 5 1 1 23400
0 23402 7 1 2 71834 23401
0 23403 5 1 1 23402
0 23404 7 1 2 77303 86429
0 23405 5 1 1 23404
0 23406 7 1 2 23403 23405
0 23407 5 2 1 23406
0 23408 7 1 2 68158 95738
0 23409 5 1 1 23408
0 23410 7 3 2 80876 84860
0 23411 5 2 1 95740
0 23412 7 1 2 72335 95741
0 23413 5 1 1 23412
0 23414 7 1 2 23409 23413
0 23415 5 1 1 23414
0 23416 7 1 2 62832 23415
0 23417 5 1 1 23416
0 23418 7 1 2 74804 94941
0 23419 5 1 1 23418
0 23420 7 1 2 10594 23419
0 23421 5 2 1 23420
0 23422 7 1 2 63329 95745
0 23423 5 1 1 23422
0 23424 7 2 2 78151 81584
0 23425 5 1 1 95747
0 23426 7 1 2 23423 23425
0 23427 5 1 1 23426
0 23428 7 1 2 72547 23427
0 23429 5 1 1 23428
0 23430 7 1 2 23417 23429
0 23431 5 1 1 23430
0 23432 7 1 2 65739 23431
0 23433 5 2 1 23432
0 23434 7 1 2 10071 94869
0 23435 5 1 1 23434
0 23436 7 1 2 73209 23435
0 23437 5 1 1 23436
0 23438 7 1 2 78359 94865
0 23439 5 1 1 23438
0 23440 7 1 2 23437 23439
0 23441 5 1 1 23440
0 23442 7 1 2 68654 23441
0 23443 5 1 1 23442
0 23444 7 1 2 95749 23443
0 23445 5 1 1 23444
0 23446 7 1 2 69794 23445
0 23447 5 1 1 23446
0 23448 7 2 2 71952 95708
0 23449 7 1 2 78075 95751
0 23450 5 1 1 23449
0 23451 7 2 2 95724 23450
0 23452 5 1 1 95753
0 23453 7 1 2 88968 23452
0 23454 5 1 1 23453
0 23455 7 1 2 23447 23454
0 23456 5 1 1 23455
0 23457 7 1 2 61853 23456
0 23458 5 1 1 23457
0 23459 7 1 2 65740 95739
0 23460 5 1 1 23459
0 23461 7 2 2 63564 78325
0 23462 7 1 2 78237 95755
0 23463 5 1 1 23462
0 23464 7 1 2 23460 23463
0 23465 5 1 1 23464
0 23466 7 1 2 62833 23465
0 23467 5 1 1 23466
0 23468 7 1 2 78076 95728
0 23469 5 1 1 23468
0 23470 7 1 2 23467 23469
0 23471 5 1 1 23470
0 23472 7 1 2 93371 23471
0 23473 5 1 1 23472
0 23474 7 1 2 23458 23473
0 23475 5 1 1 23474
0 23476 7 1 2 79251 23475
0 23477 5 1 1 23476
0 23478 7 1 2 23397 23477
0 23479 5 1 1 23478
0 23480 7 1 2 68003 23479
0 23481 5 1 1 23480
0 23482 7 1 2 71953 95718
0 23483 5 1 1 23482
0 23484 7 1 2 95699 23483
0 23485 5 1 1 23484
0 23486 7 1 2 88204 23485
0 23487 5 1 1 23486
0 23488 7 1 2 73914 95709
0 23489 5 1 1 23488
0 23490 7 1 2 95720 23489
0 23491 5 1 1 23490
0 23492 7 1 2 65145 23491
0 23493 5 1 1 23492
0 23494 7 1 2 95722 23493
0 23495 5 1 1 23494
0 23496 7 1 2 68159 95754
0 23497 5 1 1 23496
0 23498 7 1 2 66712 23497
0 23499 7 1 2 23495 23498
0 23500 5 1 1 23499
0 23501 7 1 2 23487 23500
0 23502 5 1 1 23501
0 23503 7 1 2 64925 23502
0 23504 5 1 1 23503
0 23505 7 1 2 95732 23504
0 23506 5 1 1 23505
0 23507 7 1 2 63152 79252
0 23508 7 1 2 23506 23507
0 23509 5 1 1 23508
0 23510 7 1 2 23481 23509
0 23511 5 1 1 23510
0 23512 7 1 2 64721 23511
0 23513 5 1 1 23512
0 23514 7 1 2 74898 19206
0 23515 5 2 1 23514
0 23516 7 2 2 81921 77689
0 23517 7 1 2 95757 95759
0 23518 5 1 1 23517
0 23519 7 1 2 71835 80005
0 23520 5 2 1 23519
0 23521 7 1 2 88397 92726
0 23522 7 1 2 95761 23521
0 23523 5 1 1 23522
0 23524 7 1 2 23518 23523
0 23525 5 1 1 23524
0 23526 7 1 2 70916 23525
0 23527 5 1 1 23526
0 23528 7 1 2 62406 76356
0 23529 5 4 1 23528
0 23530 7 1 2 63798 95763
0 23531 5 2 1 23530
0 23532 7 1 2 73882 95767
0 23533 5 1 1 23532
0 23534 7 1 2 63565 23533
0 23535 5 1 1 23534
0 23536 7 1 2 63799 77284
0 23537 5 1 1 23536
0 23538 7 1 2 62407 73927
0 23539 7 1 2 23537 23538
0 23540 5 1 1 23539
0 23541 7 1 2 23535 23540
0 23542 5 1 1 23541
0 23543 7 1 2 71433 23542
0 23544 5 1 1 23543
0 23545 7 2 2 62834 71636
0 23546 5 1 1 95769
0 23547 7 1 2 95726 23546
0 23548 5 1 1 23547
0 23549 7 1 2 63566 23548
0 23550 5 1 1 23549
0 23551 7 1 2 72786 73257
0 23552 5 2 1 23551
0 23553 7 1 2 77538 95771
0 23554 5 1 1 23553
0 23555 7 1 2 89381 23554
0 23556 5 1 1 23555
0 23557 7 1 2 23550 23556
0 23558 5 1 1 23557
0 23559 7 1 2 71055 23558
0 23560 5 1 1 23559
0 23561 7 1 2 23544 23560
0 23562 5 1 1 23561
0 23563 7 1 2 86954 23562
0 23564 5 1 1 23563
0 23565 7 1 2 23527 23564
0 23566 5 1 1 23565
0 23567 7 1 2 65146 23566
0 23568 5 1 1 23567
0 23569 7 1 2 74904 89370
0 23570 7 1 2 91211 23569
0 23571 7 1 2 71480 23570
0 23572 5 1 1 23571
0 23573 7 1 2 23568 23572
0 23574 5 1 1 23573
0 23575 7 1 2 68160 23574
0 23576 5 1 1 23575
0 23577 7 1 2 65147 95703
0 23578 5 1 1 23577
0 23579 7 1 2 76344 78247
0 23580 5 2 1 23579
0 23581 7 1 2 23578 95773
0 23582 5 1 1 23581
0 23583 7 1 2 78525 23582
0 23584 5 1 1 23583
0 23585 7 1 2 81172 87881
0 23586 5 1 1 23585
0 23587 7 1 2 65148 23586
0 23588 5 1 1 23587
0 23589 7 1 2 95774 23588
0 23590 5 1 1 23589
0 23591 7 1 2 79173 23590
0 23592 5 1 1 23591
0 23593 7 1 2 63962 76576
0 23594 7 1 2 84349 23593
0 23595 5 1 1 23594
0 23596 7 1 2 23592 23595
0 23597 5 1 1 23596
0 23598 7 1 2 66471 23597
0 23599 5 1 1 23598
0 23600 7 1 2 23584 23599
0 23601 5 1 1 23600
0 23602 7 1 2 81636 23601
0 23603 5 1 1 23602
0 23604 7 1 2 23576 23603
0 23605 5 1 1 23604
0 23606 7 1 2 68004 23605
0 23607 5 1 1 23606
0 23608 7 6 2 64722 76084
0 23609 7 2 2 73258 94120
0 23610 5 2 1 95781
0 23611 7 1 2 72301 95783
0 23612 5 1 1 23611
0 23613 7 1 2 95775 23612
0 23614 5 1 1 23613
0 23615 7 2 2 86955 94121
0 23616 5 1 1 95785
0 23617 7 1 2 73259 95786
0 23618 5 2 1 23617
0 23619 7 1 2 68984 88623
0 23620 5 1 1 23619
0 23621 7 1 2 87356 23620
0 23622 7 1 2 77537 23621
0 23623 5 1 1 23622
0 23624 7 1 2 95787 23623
0 23625 5 1 1 23624
0 23626 7 1 2 68005 23625
0 23627 5 1 1 23626
0 23628 7 1 2 23614 23627
0 23629 5 1 1 23628
0 23630 7 1 2 67448 23629
0 23631 5 1 1 23630
0 23632 7 2 2 89473 94446
0 23633 5 3 1 95789
0 23634 7 2 2 72302 95791
0 23635 5 2 1 95794
0 23636 7 2 2 76148 95796
0 23637 5 1 1 95798
0 23638 7 1 2 83890 95799
0 23639 5 1 1 23638
0 23640 7 1 2 23631 23639
0 23641 5 1 1 23640
0 23642 7 1 2 81451 23641
0 23643 5 1 1 23642
0 23644 7 1 2 77494 85565
0 23645 5 1 1 23644
0 23646 7 1 2 93304 23645
0 23647 5 1 1 23646
0 23648 7 1 2 76085 23647
0 23649 5 1 1 23648
0 23650 7 4 2 68006 68833
0 23651 5 1 1 95800
0 23652 7 1 2 15344 23651
0 23653 5 1 1 23652
0 23654 7 3 2 76522 78004
0 23655 7 1 2 81004 95804
0 23656 7 1 2 23653 23655
0 23657 5 1 1 23656
0 23658 7 1 2 23649 23657
0 23659 5 1 1 23658
0 23660 7 1 2 88575 23659
0 23661 5 1 1 23660
0 23662 7 1 2 23643 23661
0 23663 5 1 1 23662
0 23664 7 1 2 64926 23663
0 23665 5 1 1 23664
0 23666 7 3 2 79125 81668
0 23667 7 1 2 79523 95807
0 23668 7 1 2 90192 23667
0 23669 5 1 1 23668
0 23670 7 1 2 23665 23669
0 23671 5 1 1 23670
0 23672 7 1 2 79027 23671
0 23673 5 1 1 23672
0 23674 7 1 2 88345 87882
0 23675 5 1 1 23674
0 23676 7 1 2 91180 23675
0 23677 5 1 1 23676
0 23678 7 1 2 84482 95752
0 23679 5 1 1 23678
0 23680 7 1 2 23677 23679
0 23681 5 1 1 23680
0 23682 7 1 2 65149 23681
0 23683 5 1 1 23682
0 23684 7 2 2 79806 91212
0 23685 7 1 2 95695 95810
0 23686 5 1 1 23685
0 23687 7 1 2 23683 23686
0 23688 5 1 1 23687
0 23689 7 1 2 63567 95776
0 23690 7 1 2 23688 23689
0 23691 5 1 1 23690
0 23692 7 1 2 23673 23691
0 23693 7 1 2 23607 23692
0 23694 5 1 1 23693
0 23695 7 1 2 66955 23694
0 23696 5 1 1 23695
0 23697 7 2 2 76321 82581
0 23698 7 1 2 76369 80860
0 23699 7 1 2 95812 23698
0 23700 5 1 1 23699
0 23701 7 1 2 94882 23700
0 23702 5 1 1 23701
0 23703 7 1 2 81007 23702
0 23704 5 1 1 23703
0 23705 7 1 2 77495 83014
0 23706 5 1 1 23705
0 23707 7 1 2 81733 78725
0 23708 5 1 1 23707
0 23709 7 1 2 81787 23708
0 23710 5 2 1 23709
0 23711 7 1 2 66472 94122
0 23712 7 1 2 95814 23711
0 23713 5 1 1 23712
0 23714 7 1 2 23706 23713
0 23715 5 1 1 23714
0 23716 7 1 2 64927 23715
0 23717 5 1 1 23716
0 23718 7 1 2 68161 78726
0 23719 5 1 1 23718
0 23720 7 1 2 94862 23719
0 23721 5 3 1 23720
0 23722 7 1 2 84302 81008
0 23723 7 1 2 95816 23722
0 23724 5 1 1 23723
0 23725 7 1 2 23717 23724
0 23726 5 1 1 23725
0 23727 7 1 2 73210 23726
0 23728 5 1 1 23727
0 23729 7 1 2 23704 23728
0 23730 5 1 1 23729
0 23731 7 1 2 83333 23730
0 23732 5 1 1 23731
0 23733 7 1 2 68410 73977
0 23734 5 1 1 23733
0 23735 7 1 2 89622 23734
0 23736 5 1 1 23735
0 23737 7 1 2 81769 75066
0 23738 7 1 2 94123 23737
0 23739 5 1 1 23738
0 23740 7 1 2 23736 23739
0 23741 5 1 1 23740
0 23742 7 1 2 62097 23741
0 23743 5 1 1 23742
0 23744 7 1 2 72158 90505
0 23745 5 1 1 23744
0 23746 7 1 2 90506 81428
0 23747 5 2 1 23746
0 23748 7 1 2 84359 95819
0 23749 7 1 2 23745 23748
0 23750 5 1 1 23749
0 23751 7 1 2 13015 23750
0 23752 5 1 1 23751
0 23753 7 1 2 94088 23752
0 23754 5 1 1 23753
0 23755 7 1 2 23743 23754
0 23756 5 1 1 23755
0 23757 7 1 2 66473 23756
0 23758 5 1 1 23757
0 23759 7 1 2 86364 92498
0 23760 5 1 1 23759
0 23761 7 1 2 23758 23760
0 23762 5 1 1 23761
0 23763 7 1 2 64723 23762
0 23764 5 1 1 23763
0 23765 7 3 2 66474 80486
0 23766 5 1 1 95821
0 23767 7 1 2 88667 78710
0 23768 7 1 2 95822 23767
0 23769 5 1 1 23768
0 23770 7 1 2 70060 23769
0 23771 7 1 2 23764 23770
0 23772 5 1 1 23771
0 23773 7 1 2 62098 87523
0 23774 5 1 1 23773
0 23775 7 1 2 75675 84844
0 23776 7 1 2 78949 23775
0 23777 5 1 1 23776
0 23778 7 5 2 64724 72622
0 23779 7 2 2 63153 88969
0 23780 7 1 2 95824 95829
0 23781 5 1 1 23780
0 23782 7 1 2 23777 23781
0 23783 5 1 1 23782
0 23784 7 1 2 62835 23783
0 23785 5 1 1 23784
0 23786 7 2 2 76846 82545
0 23787 7 1 2 88853 95831
0 23788 5 1 1 23787
0 23789 7 1 2 23785 23788
0 23790 5 1 1 23789
0 23791 7 1 2 73211 23790
0 23792 5 1 1 23791
0 23793 7 1 2 23774 23792
0 23794 5 1 1 23793
0 23795 7 1 2 66475 23794
0 23796 5 1 1 23795
0 23797 7 5 2 62836 88946
0 23798 5 1 1 95833
0 23799 7 1 2 88982 23798
0 23800 5 4 1 23799
0 23801 7 3 2 70917 73212
0 23802 7 1 2 68985 75627
0 23803 5 1 1 23802
0 23804 7 1 2 95842 23803
0 23805 7 1 2 95838 23804
0 23806 5 1 1 23805
0 23807 7 1 2 20649 23806
0 23808 5 1 1 23807
0 23809 7 1 2 89083 23808
0 23810 5 1 1 23809
0 23811 7 1 2 23796 23810
0 23812 5 1 1 23811
0 23813 7 1 2 68411 23812
0 23814 5 1 1 23813
0 23815 7 1 2 76370 79807
0 23816 7 1 2 95813 23815
0 23817 7 1 2 91974 23816
0 23818 5 1 1 23817
0 23819 7 1 2 65150 23818
0 23820 7 1 2 23814 23819
0 23821 5 1 1 23820
0 23822 7 1 2 66713 23821
0 23823 7 1 2 23772 23822
0 23824 5 1 1 23823
0 23825 7 1 2 23732 23824
0 23826 5 1 1 23825
0 23827 7 1 2 73004 23826
0 23828 5 1 1 23827
0 23829 7 1 2 90336 94873
0 23830 5 1 1 23829
0 23831 7 1 2 73935 94866
0 23832 5 1 1 23831
0 23833 7 1 2 23830 23832
0 23834 5 1 1 23833
0 23835 7 1 2 68655 23834
0 23836 5 1 1 23835
0 23837 7 1 2 95750 23836
0 23838 5 1 1 23837
0 23839 7 1 2 64928 23838
0 23840 5 1 1 23839
0 23841 7 1 2 65151 74181
0 23842 5 1 1 23841
0 23843 7 2 2 67248 74077
0 23844 5 1 1 95845
0 23845 7 1 2 91213 95846
0 23846 5 1 1 23845
0 23847 7 1 2 23842 23846
0 23848 5 1 1 23847
0 23849 7 1 2 88947 73915
0 23850 7 1 2 23848 23849
0 23851 5 1 1 23850
0 23852 7 1 2 23840 23851
0 23853 5 1 1 23852
0 23854 7 1 2 66714 23853
0 23855 5 1 1 23854
0 23856 7 2 2 83053 88507
0 23857 7 1 2 95811 95847
0 23858 5 1 1 23857
0 23859 7 1 2 23855 23858
0 23860 5 1 1 23859
0 23861 7 1 2 78927 79253
0 23862 7 1 2 23860 23861
0 23863 5 1 1 23862
0 23864 7 1 2 23828 23863
0 23865 7 1 2 23696 23864
0 23866 7 1 2 23513 23865
0 23867 5 1 1 23866
0 23868 7 1 2 64514 23867
0 23869 5 1 1 23868
0 23870 7 1 2 85711 87161
0 23871 5 1 1 23870
0 23872 7 1 2 88885 23871
0 23873 5 1 1 23872
0 23874 7 1 2 61854 23873
0 23875 5 1 1 23874
0 23876 7 1 2 4125 23875
0 23877 5 1 1 23876
0 23878 7 1 2 68162 23877
0 23879 5 1 1 23878
0 23880 7 1 2 89149 23879
0 23881 5 1 1 23880
0 23882 7 1 2 68007 23881
0 23883 5 1 1 23882
0 23884 7 1 2 86160 92264
0 23885 7 1 2 92993 23884
0 23886 5 1 1 23885
0 23887 7 1 2 23883 23886
0 23888 5 1 1 23887
0 23889 7 1 2 95764 23888
0 23890 5 1 1 23889
0 23891 7 3 2 63330 76847
0 23892 5 1 1 95849
0 23893 7 1 2 68986 95834
0 23894 5 1 1 23893
0 23895 7 1 2 23892 23894
0 23896 5 1 1 23895
0 23897 7 1 2 71230 23896
0 23898 5 1 1 23897
0 23899 7 1 2 68163 71003
0 23900 5 1 1 23899
0 23901 7 1 2 88983 23900
0 23902 5 4 1 23901
0 23903 7 1 2 73686 95852
0 23904 5 1 1 23903
0 23905 7 1 2 23898 23904
0 23906 5 1 1 23905
0 23907 7 1 2 70695 23906
0 23908 5 1 1 23907
0 23909 7 1 2 91125 95835
0 23910 5 1 1 23909
0 23911 7 1 2 87201 89905
0 23912 5 1 1 23911
0 23913 7 1 2 23910 23912
0 23914 5 1 1 23913
0 23915 7 1 2 73452 23914
0 23916 5 1 1 23915
0 23917 7 1 2 68164 79224
0 23918 7 1 2 75203 80349
0 23919 7 1 2 23917 23918
0 23920 5 1 1 23919
0 23921 7 1 2 23916 23920
0 23922 5 1 1 23921
0 23923 7 1 2 64125 23922
0 23924 5 1 1 23923
0 23925 7 1 2 73687 95850
0 23926 5 1 1 23925
0 23927 7 3 2 67449 73777
0 23928 5 1 1 95856
0 23929 7 1 2 68834 95857
0 23930 5 1 1 23929
0 23931 7 1 2 71507 23930
0 23932 5 1 1 23931
0 23933 7 1 2 89398 23932
0 23934 5 1 1 23933
0 23935 7 1 2 23926 23934
0 23936 7 1 2 23924 23935
0 23937 7 1 2 23908 23936
0 23938 5 1 1 23937
0 23939 7 1 2 66715 23938
0 23940 5 1 1 23939
0 23941 7 1 2 67249 90338
0 23942 5 1 1 23941
0 23943 7 1 2 68656 23942
0 23944 5 1 1 23943
0 23945 7 2 2 67450 77418
0 23946 5 6 1 95859
0 23947 7 1 2 64126 84740
0 23948 5 1 1 23947
0 23949 7 1 2 95861 23948
0 23950 5 1 1 23949
0 23951 7 1 2 70696 23950
0 23952 5 1 1 23951
0 23953 7 1 2 23944 23952
0 23954 5 1 1 23953
0 23955 7 1 2 92008 23954
0 23956 5 1 1 23955
0 23957 7 1 2 23940 23956
0 23958 5 1 1 23957
0 23959 7 1 2 90760 23958
0 23960 5 1 1 23959
0 23961 7 1 2 23890 23960
0 23962 5 1 1 23961
0 23963 7 1 2 66476 23962
0 23964 5 1 1 23963
0 23965 7 1 2 86774 95801
0 23966 7 1 2 91792 23965
0 23967 7 1 2 95765 23966
0 23968 5 1 1 23967
0 23969 7 1 2 23964 23968
0 23970 5 1 1 23969
0 23971 7 1 2 79363 23970
0 23972 5 1 1 23971
0 23973 7 1 2 76047 91727
0 23974 5 1 1 23973
0 23975 7 1 2 23637 23974
0 23976 5 1 1 23975
0 23977 7 1 2 73453 23976
0 23978 5 1 1 23977
0 23979 7 1 2 76086 75272
0 23980 5 1 1 23979
0 23981 7 1 2 67250 76149
0 23982 7 1 2 95710 23981
0 23983 5 1 1 23982
0 23984 7 1 2 23980 23983
0 23985 7 1 2 23978 23984
0 23986 5 1 1 23985
0 23987 7 1 2 84483 23986
0 23988 5 1 1 23987
0 23989 7 5 2 67451 72623
0 23990 5 1 1 95867
0 23991 7 2 2 68835 23990
0 23992 5 1 1 95872
0 23993 7 1 2 70697 11693
0 23994 7 1 2 23992 23993
0 23995 5 1 1 23994
0 23996 7 1 2 71508 95768
0 23997 7 1 2 23995 23996
0 23998 5 1 1 23997
0 23999 7 1 2 92930 23998
0 24000 5 1 1 23999
0 24001 7 1 2 23988 24000
0 24002 5 1 1 24001
0 24003 7 1 2 70061 24002
0 24004 5 1 1 24003
0 24005 7 3 2 61569 87245
0 24006 5 1 1 95874
0 24007 7 1 2 16919 24006
0 24008 5 7 1 24007
0 24009 7 5 2 68165 71231
0 24010 7 1 2 80877 95884
0 24011 7 1 2 95766 24010
0 24012 7 1 2 95877 24011
0 24013 5 1 1 24012
0 24014 7 1 2 24004 24013
0 24015 5 1 1 24014
0 24016 7 1 2 64515 24015
0 24017 5 1 1 24016
0 24018 7 1 2 86214 87511
0 24019 5 1 1 24018
0 24020 7 1 2 81676 81864
0 24021 7 1 2 86775 24020
0 24022 7 1 2 24019 24021
0 24023 5 1 1 24022
0 24024 7 1 2 24017 24023
0 24025 5 1 1 24024
0 24026 7 1 2 64725 24025
0 24027 5 1 1 24026
0 24028 7 2 2 68166 65741
0 24029 7 2 2 64929 78042
0 24030 7 1 2 89594 93272
0 24031 7 1 2 95891 24030
0 24032 5 1 1 24031
0 24033 7 1 2 82053 85878
0 24034 5 1 1 24033
0 24035 7 1 2 10534 24034
0 24036 5 1 1 24035
0 24037 7 1 2 78928 92021
0 24038 7 1 2 24036 24037
0 24039 5 1 1 24038
0 24040 7 1 2 24032 24039
0 24041 5 1 1 24040
0 24042 7 1 2 95889 24041
0 24043 5 1 1 24042
0 24044 7 2 2 83118 78474
0 24045 7 1 2 95325 95893
0 24046 5 1 1 24045
0 24047 7 2 2 68167 79174
0 24048 7 1 2 84352 85929
0 24049 7 1 2 95895 24048
0 24050 5 1 1 24049
0 24051 7 1 2 24046 24050
0 24052 5 1 1 24051
0 24053 7 1 2 76150 24052
0 24054 5 1 1 24053
0 24055 7 1 2 24043 24054
0 24056 5 1 1 24055
0 24057 7 1 2 64516 24056
0 24058 5 1 1 24057
0 24059 7 1 2 82766 79787
0 24060 7 1 2 95697 24059
0 24061 5 1 1 24060
0 24062 7 1 2 24058 24061
0 24063 5 1 1 24062
0 24064 7 1 2 84621 24063
0 24065 5 1 1 24064
0 24066 7 1 2 24027 24065
0 24067 7 1 2 23972 24066
0 24068 5 1 1 24067
0 24069 7 1 2 74319 24068
0 24070 5 1 1 24069
0 24071 7 1 2 23869 24070
0 24072 5 1 1 24071
0 24073 7 1 2 69188 24072
0 24074 5 1 1 24073
0 24075 7 6 2 64344 82808
0 24076 7 3 2 80140 95897
0 24077 5 2 1 95903
0 24078 7 1 2 68836 95904
0 24079 5 1 1 24078
0 24080 7 2 2 80806 91841
0 24081 5 1 1 95908
0 24082 7 1 2 24079 24081
0 24083 5 1 1 24082
0 24084 7 1 2 67452 24083
0 24085 5 1 1 24084
0 24086 7 2 2 91842 95802
0 24087 5 1 1 95910
0 24088 7 1 2 95906 24087
0 24089 5 1 1 24088
0 24090 7 1 2 68657 24089
0 24091 5 1 1 24090
0 24092 7 1 2 24085 24091
0 24093 5 1 1 24092
0 24094 7 1 2 81988 24093
0 24095 5 1 1 24094
0 24096 7 3 2 78950 92766
0 24097 7 1 2 87426 87164
0 24098 7 1 2 95912 24097
0 24099 5 1 1 24098
0 24100 7 1 2 24095 24099
0 24101 5 1 1 24100
0 24102 7 1 2 61570 24101
0 24103 5 1 1 24102
0 24104 7 1 2 64517 95014
0 24105 5 1 1 24104
0 24106 7 1 2 83243 24105
0 24107 5 2 1 24106
0 24108 7 2 2 68658 69189
0 24109 7 1 2 92075 95917
0 24110 7 1 2 95915 24109
0 24111 5 1 1 24110
0 24112 7 1 2 24103 24111
0 24113 5 1 1 24112
0 24114 7 1 2 67251 24113
0 24115 5 1 1 24114
0 24116 7 1 2 82780 85004
0 24117 7 3 2 69363 83291
0 24118 7 1 2 87862 95919
0 24119 7 1 2 24116 24118
0 24120 5 1 1 24119
0 24121 7 1 2 24115 24120
0 24122 5 1 1 24121
0 24123 7 1 2 65152 24122
0 24124 5 1 1 24123
0 24125 7 1 2 68008 92049
0 24126 5 1 1 24125
0 24127 7 1 2 66477 71434
0 24128 7 1 2 83236 24127
0 24129 5 1 1 24128
0 24130 7 1 2 24126 24129
0 24131 5 1 1 24130
0 24132 7 2 2 79533 73454
0 24133 7 1 2 94784 95922
0 24134 7 1 2 24131 24133
0 24135 5 1 1 24134
0 24136 7 1 2 24124 24135
0 24137 5 1 1 24136
0 24138 7 1 2 68412 24137
0 24139 5 1 1 24138
0 24140 7 1 2 79671 81260
0 24141 5 1 1 24140
0 24142 7 1 2 78238 78776
0 24143 7 1 2 91207 24142
0 24144 5 1 1 24143
0 24145 7 1 2 24141 24144
0 24146 5 1 1 24145
0 24147 7 1 2 71435 24146
0 24148 5 1 1 24147
0 24149 7 1 2 83024 91916
0 24150 5 1 1 24149
0 24151 7 1 2 24148 24150
0 24152 5 1 1 24151
0 24153 7 1 2 81533 93694
0 24154 7 1 2 24152 24153
0 24155 5 1 1 24154
0 24156 7 1 2 24139 24155
0 24157 5 1 1 24156
0 24158 7 1 2 66956 24157
0 24159 5 1 1 24158
0 24160 7 1 2 79077 82511
0 24161 5 1 1 24160
0 24162 7 1 2 18049 24161
0 24163 5 1 1 24162
0 24164 7 1 2 61855 24163
0 24165 5 1 1 24164
0 24166 7 1 2 83476 74936
0 24167 5 1 1 24166
0 24168 7 1 2 8270 24167
0 24169 5 1 1 24168
0 24170 7 1 2 78265 24169
0 24171 5 1 1 24170
0 24172 7 1 2 24165 24171
0 24173 5 1 1 24172
0 24174 7 1 2 68009 24173
0 24175 5 1 1 24174
0 24176 7 2 2 66716 79126
0 24177 7 2 2 74805 80744
0 24178 7 1 2 95924 95926
0 24179 5 1 1 24178
0 24180 7 1 2 24175 24179
0 24181 5 1 1 24180
0 24182 7 1 2 70062 24181
0 24183 5 1 1 24182
0 24184 7 1 2 76670 81858
0 24185 7 1 2 74916 24184
0 24186 5 1 1 24185
0 24187 7 1 2 24183 24186
0 24188 5 1 1 24187
0 24189 7 1 2 66478 24188
0 24190 5 1 1 24189
0 24191 7 1 2 79127 90534
0 24192 7 1 2 95746 24191
0 24193 5 1 1 24192
0 24194 7 1 2 24190 24193
0 24195 5 1 1 24194
0 24196 7 1 2 80271 92767
0 24197 7 1 2 24195 24196
0 24198 5 1 1 24197
0 24199 7 1 2 24159 24198
0 24200 5 1 1 24199
0 24201 7 1 2 68168 24200
0 24202 5 1 1 24201
0 24203 7 3 2 63331 69190
0 24204 7 3 2 95251 95928
0 24205 7 1 2 76627 83622
0 24206 5 1 1 24205
0 24207 7 1 2 91695 24206
0 24208 5 1 1 24207
0 24209 7 1 2 82211 77662
0 24210 5 1 1 24209
0 24211 7 1 2 88578 24210
0 24212 7 1 2 24208 24211
0 24213 5 1 1 24212
0 24214 7 1 2 68837 24213
0 24215 5 1 1 24214
0 24216 7 1 2 1787 24215
0 24217 5 1 1 24216
0 24218 7 1 2 79175 24217
0 24219 5 1 1 24218
0 24220 7 1 2 75479 74276
0 24221 7 1 2 90432 24220
0 24222 5 1 1 24221
0 24223 7 1 2 24219 24222
0 24224 5 1 1 24223
0 24225 7 1 2 95931 24224
0 24226 5 1 1 24225
0 24227 7 1 2 24202 24226
0 24228 5 1 1 24227
0 24229 7 1 2 78005 24228
0 24230 5 1 1 24229
0 24231 7 1 2 71954 92701
0 24232 5 2 1 24231
0 24233 7 1 2 90793 94124
0 24234 7 1 2 75387 24233
0 24235 5 1 1 24234
0 24236 7 1 2 95934 24235
0 24237 5 2 1 24236
0 24238 7 1 2 69795 95936
0 24239 5 1 1 24238
0 24240 7 1 2 88223 81209
0 24241 7 1 2 85285 24240
0 24242 5 1 1 24241
0 24243 7 1 2 24239 24242
0 24244 5 1 1 24243
0 24245 7 1 2 70698 24244
0 24246 5 1 1 24245
0 24247 7 3 2 62837 79682
0 24248 5 2 1 95938
0 24249 7 1 2 65984 95939
0 24250 5 1 1 24249
0 24251 7 1 2 95862 24250
0 24252 5 1 1 24251
0 24253 7 1 2 88970 74288
0 24254 7 1 2 24252 24253
0 24255 5 1 1 24254
0 24256 7 1 2 24246 24255
0 24257 5 1 1 24256
0 24258 7 1 2 61856 24257
0 24259 5 1 1 24258
0 24260 7 1 2 89474 95868
0 24261 5 2 1 24260
0 24262 7 1 2 77840 95943
0 24263 5 1 1 24262
0 24264 7 1 2 89659 92156
0 24265 7 1 2 24263 24264
0 24266 5 1 1 24265
0 24267 7 1 2 24259 24266
0 24268 5 1 1 24267
0 24269 7 1 2 66479 24268
0 24270 5 1 1 24269
0 24271 7 2 2 70699 95937
0 24272 7 1 2 83314 95945
0 24273 5 1 1 24272
0 24274 7 1 2 24270 24273
0 24275 5 1 1 24274
0 24276 7 1 2 63154 24275
0 24277 5 1 1 24276
0 24278 7 2 2 69796 84360
0 24279 7 1 2 88848 95947
0 24280 5 1 1 24279
0 24281 7 4 2 61857 76848
0 24282 5 5 1 95949
0 24283 7 1 2 87436 95950
0 24284 5 1 1 24283
0 24285 7 1 2 24280 24284
0 24286 5 1 1 24285
0 24287 7 1 2 65742 24286
0 24288 5 1 1 24287
0 24289 7 2 2 70918 72830
0 24290 7 1 2 76763 88050
0 24291 7 1 2 95958 24290
0 24292 5 1 1 24291
0 24293 7 1 2 24288 24292
0 24294 5 1 1 24293
0 24295 7 1 2 85422 24294
0 24296 5 1 1 24295
0 24297 7 2 2 72624 82395
0 24298 7 2 2 74864 95960
0 24299 7 2 2 66717 72225
0 24300 7 1 2 81842 95964
0 24301 7 1 2 95962 24300
0 24302 5 1 1 24301
0 24303 7 1 2 24296 24302
0 24304 5 1 1 24303
0 24305 7 1 2 63155 24304
0 24306 5 1 1 24305
0 24307 7 2 2 62838 81734
0 24308 7 1 2 83698 95966
0 24309 7 1 2 95963 24308
0 24310 5 1 1 24309
0 24311 7 1 2 24306 24310
0 24312 5 1 1 24311
0 24313 7 1 2 73455 24312
0 24314 5 1 1 24313
0 24315 7 1 2 74842 79570
0 24316 5 1 1 24315
0 24317 7 1 2 68413 24316
0 24318 5 1 1 24317
0 24319 7 1 2 91126 24318
0 24320 5 1 1 24319
0 24321 7 1 2 68838 72831
0 24322 5 2 1 24321
0 24323 7 1 2 65985 95968
0 24324 7 1 2 82692 24323
0 24325 5 1 1 24324
0 24326 7 1 2 24320 24325
0 24327 5 1 1 24326
0 24328 7 1 2 62099 24327
0 24329 5 1 1 24328
0 24330 7 2 2 84559 86041
0 24331 7 1 2 81192 95970
0 24332 5 1 1 24331
0 24333 7 1 2 24329 24332
0 24334 5 1 1 24333
0 24335 7 1 2 64930 24334
0 24336 5 1 1 24335
0 24337 7 1 2 74320 94125
0 24338 5 1 1 24337
0 24339 7 2 2 68839 94126
0 24340 5 4 1 95972
0 24341 7 1 2 67453 95973
0 24342 5 3 1 24341
0 24343 7 1 2 81178 95978
0 24344 5 1 1 24343
0 24345 7 1 2 66957 24344
0 24346 5 1 1 24345
0 24347 7 1 2 76345 75109
0 24348 5 1 1 24347
0 24349 7 1 2 24346 24348
0 24350 5 1 1 24349
0 24351 7 1 2 74806 24350
0 24352 5 1 1 24351
0 24353 7 1 2 24338 24352
0 24354 5 1 1 24353
0 24355 7 1 2 69797 82185
0 24356 7 1 2 24354 24355
0 24357 5 1 1 24356
0 24358 7 1 2 24336 24357
0 24359 5 1 1 24358
0 24360 7 1 2 91306 24359
0 24361 5 1 1 24360
0 24362 7 2 2 76000 90235
0 24363 7 2 2 84643 95863
0 24364 5 1 1 95983
0 24365 7 1 2 73456 84940
0 24366 5 1 1 24365
0 24367 7 1 2 95984 24366
0 24368 5 1 1 24367
0 24369 7 1 2 74865 24368
0 24370 5 1 1 24369
0 24371 7 1 2 63800 76523
0 24372 5 1 1 24371
0 24373 7 1 2 84963 24372
0 24374 5 1 1 24373
0 24375 7 1 2 65986 85785
0 24376 5 1 1 24375
0 24377 7 1 2 67252 10063
0 24378 7 1 2 24376 24377
0 24379 5 1 1 24378
0 24380 7 1 2 24374 24379
0 24381 7 1 2 24370 24380
0 24382 5 1 1 24381
0 24383 7 1 2 95981 24382
0 24384 5 1 1 24383
0 24385 7 2 2 65743 86765
0 24386 7 7 2 68414 64931
0 24387 7 1 2 95514 95987
0 24388 7 1 2 95985 24387
0 24389 5 1 1 24388
0 24390 7 1 2 81157 95701
0 24391 5 1 1 24390
0 24392 7 1 2 76465 95031
0 24393 7 1 2 24391 24392
0 24394 5 1 1 24393
0 24395 7 1 2 24389 24394
0 24396 5 1 1 24395
0 24397 7 1 2 62100 24396
0 24398 5 1 1 24397
0 24399 7 1 2 24384 24398
0 24400 5 1 1 24399
0 24401 7 1 2 83119 24400
0 24402 5 1 1 24401
0 24403 7 1 2 61571 87243
0 24404 7 1 2 95946 24403
0 24405 5 1 1 24404
0 24406 7 1 2 24402 24405
0 24407 7 1 2 24361 24406
0 24408 7 1 2 24314 24407
0 24409 7 1 2 24277 24408
0 24410 5 1 1 24409
0 24411 7 1 2 70063 24410
0 24412 5 1 1 24411
0 24413 7 1 2 93509 94127
0 24414 5 1 1 24413
0 24415 7 1 2 93506 24414
0 24416 5 1 1 24415
0 24417 7 1 2 73005 24416
0 24418 5 1 1 24417
0 24419 7 1 2 78326 86677
0 24420 5 1 1 24419
0 24421 7 1 2 76749 80006
0 24422 5 2 1 24421
0 24423 7 1 2 86609 73898
0 24424 7 1 2 95994 24423
0 24425 5 1 1 24424
0 24426 7 1 2 24420 24425
0 24427 7 1 2 24418 24426
0 24428 5 2 1 24427
0 24429 7 1 2 95035 95996
0 24430 5 1 1 24429
0 24431 7 1 2 81301 95997
0 24432 5 2 1 24431
0 24433 7 2 2 75770 89722
0 24434 7 2 2 76346 89936
0 24435 7 1 2 96000 96002
0 24436 5 1 1 24435
0 24437 7 1 2 95998 24436
0 24438 5 1 1 24437
0 24439 7 1 2 61858 24438
0 24440 5 1 1 24439
0 24441 7 1 2 85125 75826
0 24442 7 1 2 96003 24441
0 24443 5 1 1 24442
0 24444 7 1 2 24440 24443
0 24445 5 1 1 24444
0 24446 7 1 2 76151 24445
0 24447 5 1 1 24446
0 24448 7 1 2 71955 86208
0 24449 5 1 1 24448
0 24450 7 1 2 91926 24449
0 24451 5 1 1 24450
0 24452 7 1 2 73457 24451
0 24453 5 1 1 24452
0 24454 7 1 2 15156 24453
0 24455 5 1 1 24454
0 24456 7 2 2 77241 75418
0 24457 7 1 2 82563 96004
0 24458 7 1 2 24455 24457
0 24459 5 1 1 24458
0 24460 7 1 2 24447 24459
0 24461 5 1 1 24460
0 24462 7 1 2 69798 24461
0 24463 5 1 1 24462
0 24464 7 1 2 24430 24463
0 24465 7 1 2 24412 24464
0 24466 5 1 1 24465
0 24467 7 1 2 69561 24466
0 24468 5 1 1 24467
0 24469 7 1 2 71232 95388
0 24470 5 2 1 24469
0 24471 7 1 2 79712 96006
0 24472 5 1 1 24471
0 24473 7 1 2 65153 24472
0 24474 7 1 2 95020 24473
0 24475 5 1 1 24474
0 24476 7 1 2 77242 82037
0 24477 7 1 2 88849 24476
0 24478 5 1 1 24477
0 24479 7 1 2 24475 24478
0 24480 5 1 1 24479
0 24481 7 1 2 67682 24480
0 24482 5 1 1 24481
0 24483 7 1 2 87393 80659
0 24484 5 1 1 24483
0 24485 7 1 2 88846 94654
0 24486 5 1 1 24485
0 24487 7 1 2 24484 24486
0 24488 5 1 1 24487
0 24489 7 1 2 86094 24488
0 24490 5 1 1 24489
0 24491 7 1 2 24482 24490
0 24492 5 1 1 24491
0 24493 7 1 2 63332 24492
0 24494 5 1 1 24493
0 24495 7 1 2 77884 85792
0 24496 5 2 1 24495
0 24497 7 1 2 88894 83505
0 24498 7 1 2 96008 24497
0 24499 5 1 1 24498
0 24500 7 1 2 24494 24499
0 24501 5 1 1 24500
0 24502 7 1 2 86696 24501
0 24503 5 1 1 24502
0 24504 7 1 2 85188 92397
0 24505 7 1 2 75388 24504
0 24506 5 1 1 24505
0 24507 7 1 2 95935 24506
0 24508 5 1 1 24507
0 24509 7 1 2 70700 24508
0 24510 5 1 1 24509
0 24511 7 1 2 89975 95389
0 24512 5 1 1 24511
0 24513 7 1 2 63963 84981
0 24514 7 1 2 75389 24513
0 24515 5 1 1 24514
0 24516 7 1 2 24512 24515
0 24517 5 1 1 24516
0 24518 7 1 2 68169 24517
0 24519 5 1 1 24518
0 24520 7 1 2 73947 96009
0 24521 5 1 1 24520
0 24522 7 1 2 5071 24521
0 24523 5 1 1 24522
0 24524 7 1 2 63333 77932
0 24525 7 1 2 24523 24524
0 24526 5 1 1 24525
0 24527 7 1 2 24519 24526
0 24528 5 1 1 24527
0 24529 7 1 2 64127 24528
0 24530 5 1 1 24529
0 24531 7 1 2 24510 24530
0 24532 5 1 1 24531
0 24533 7 1 2 70064 24532
0 24534 5 1 1 24533
0 24535 7 1 2 95999 24534
0 24536 5 1 1 24535
0 24537 7 1 2 77243 79148
0 24538 7 1 2 24536 24537
0 24539 5 1 1 24538
0 24540 7 1 2 24503 24539
0 24541 7 1 2 24468 24540
0 24542 5 1 1 24541
0 24543 7 1 2 93089 24542
0 24544 5 1 1 24543
0 24545 7 1 2 83054 71576
0 24546 5 1 1 24545
0 24547 7 1 2 63964 81452
0 24548 5 1 1 24547
0 24549 7 1 2 24546 24548
0 24550 5 2 1 24549
0 24551 7 1 2 75349 96010
0 24552 5 1 1 24551
0 24553 7 1 2 90179 78446
0 24554 5 1 1 24553
0 24555 7 1 2 62839 85326
0 24556 5 1 1 24555
0 24557 7 1 2 24554 24556
0 24558 5 1 1 24557
0 24559 7 1 2 64932 24558
0 24560 5 1 1 24559
0 24561 7 1 2 24552 24560
0 24562 5 1 1 24561
0 24563 7 1 2 61572 24562
0 24564 5 1 1 24563
0 24565 7 2 2 66718 89638
0 24566 5 1 1 96012
0 24567 7 1 2 75633 24566
0 24568 5 1 1 24567
0 24569 7 1 2 63334 24568
0 24570 5 1 1 24569
0 24571 7 2 2 69799 71577
0 24572 7 1 2 83055 96014
0 24573 5 1 1 24572
0 24574 7 1 2 24570 24573
0 24575 5 1 1 24574
0 24576 7 1 2 76087 24575
0 24577 5 1 1 24576
0 24578 7 1 2 24564 24577
0 24579 5 1 1 24578
0 24580 7 1 2 72058 24579
0 24581 5 1 1 24580
0 24582 7 1 2 63965 86454
0 24583 7 1 2 95878 24582
0 24584 5 1 1 24583
0 24585 7 1 2 24581 24584
0 24586 5 1 1 24585
0 24587 7 1 2 69562 24586
0 24588 5 1 1 24587
0 24589 7 1 2 79149 91269
0 24590 7 1 2 93551 24589
0 24591 5 1 1 24590
0 24592 7 1 2 24588 24591
0 24593 5 1 1 24592
0 24594 7 1 2 78727 24593
0 24595 5 1 1 24594
0 24596 7 1 2 93552 95027
0 24597 5 1 1 24596
0 24598 7 1 2 24595 24597
0 24599 5 1 1 24598
0 24600 7 1 2 73006 24599
0 24601 5 1 1 24600
0 24602 7 1 2 61859 95853
0 24603 5 1 1 24602
0 24604 7 1 2 68987 93372
0 24605 5 1 1 24604
0 24606 7 1 2 24603 24605
0 24607 5 2 1 24606
0 24608 7 1 2 76152 96016
0 24609 5 1 1 24608
0 24610 7 1 2 90180 76589
0 24611 5 2 1 24610
0 24612 7 1 2 24609 96018
0 24613 5 1 1 24612
0 24614 7 1 2 70065 76466
0 24615 7 1 2 24613 24614
0 24616 5 1 1 24615
0 24617 7 1 2 88260 77105
0 24618 7 1 2 95032 24617
0 24619 5 1 1 24618
0 24620 7 1 2 24616 24619
0 24621 5 1 1 24620
0 24622 7 1 2 62101 24621
0 24623 5 1 1 24622
0 24624 7 2 2 82663 80837
0 24625 7 1 2 85669 96020
0 24626 7 1 2 71100 24625
0 24627 5 1 1 24626
0 24628 7 1 2 24623 24627
0 24629 5 1 1 24628
0 24630 7 1 2 65987 91185
0 24631 7 1 2 24629 24630
0 24632 5 1 1 24631
0 24633 7 1 2 24601 24632
0 24634 5 1 1 24633
0 24635 7 1 2 93090 24634
0 24636 5 1 1 24635
0 24637 7 3 2 87884 93547
0 24638 7 1 2 78728 96022
0 24639 5 1 1 24638
0 24640 7 1 2 88329 83464
0 24641 5 1 1 24640
0 24642 7 1 2 24639 24641
0 24643 5 1 1 24642
0 24644 7 1 2 64933 24643
0 24645 5 1 1 24644
0 24646 7 1 2 68415 96023
0 24647 5 1 1 24646
0 24648 7 2 2 76322 83613
0 24649 5 1 1 96025
0 24650 7 1 2 68988 96026
0 24651 5 1 1 24650
0 24652 7 1 2 24647 24651
0 24653 5 1 1 24652
0 24654 7 2 2 65154 24653
0 24655 7 1 2 74238 96027
0 24656 5 1 1 24655
0 24657 7 1 2 24645 24656
0 24658 5 1 1 24657
0 24659 7 1 2 66719 24658
0 24660 5 1 1 24659
0 24661 7 1 2 83073 24660
0 24662 5 1 1 24661
0 24663 7 1 2 64934 96028
0 24664 5 1 1 24663
0 24665 7 1 2 82753 24664
0 24666 5 1 1 24665
0 24667 7 1 2 95777 24666
0 24668 7 1 2 24662 24667
0 24669 5 1 1 24668
0 24670 7 1 2 89375 10185
0 24671 5 2 1 24670
0 24672 7 1 2 66480 96029
0 24673 5 1 1 24672
0 24674 7 1 2 83012 78515
0 24675 5 1 1 24674
0 24676 7 1 2 24673 24675
0 24677 5 1 1 24676
0 24678 7 1 2 92148 24677
0 24679 5 2 1 24678
0 24680 7 1 2 88708 94537
0 24681 5 1 1 24680
0 24682 7 1 2 85209 89909
0 24683 5 1 1 24682
0 24684 7 1 2 24681 24683
0 24685 5 1 1 24684
0 24686 7 1 2 66720 24685
0 24687 5 1 1 24686
0 24688 7 1 2 68170 85210
0 24689 5 1 1 24688
0 24690 7 1 2 95743 24689
0 24691 5 2 1 24690
0 24692 7 1 2 90055 96033
0 24693 5 1 1 24692
0 24694 7 1 2 24687 24693
0 24695 5 1 1 24694
0 24696 7 1 2 72881 24695
0 24697 5 1 1 24696
0 24698 7 1 2 96031 24697
0 24699 5 1 1 24698
0 24700 7 1 2 64726 24699
0 24701 5 1 1 24700
0 24702 7 1 2 81343 88508
0 24703 7 1 2 85796 87344
0 24704 7 1 2 24702 24703
0 24705 5 1 1 24704
0 24706 7 2 2 88310 82741
0 24707 5 1 1 96035
0 24708 7 1 2 64727 96030
0 24709 5 1 1 24708
0 24710 7 1 2 24707 24709
0 24711 5 1 1 24710
0 24712 7 1 2 66481 24711
0 24713 5 1 1 24712
0 24714 7 1 2 92230 92534
0 24715 5 1 1 24714
0 24716 7 1 2 24713 24715
0 24717 5 1 1 24716
0 24718 7 1 2 77891 81193
0 24719 7 1 2 24717 24718
0 24720 5 1 1 24719
0 24721 7 1 2 24705 24720
0 24722 7 1 2 24701 24721
0 24723 5 1 1 24722
0 24724 7 1 2 62840 24723
0 24725 5 1 1 24724
0 24726 7 1 2 88360 96036
0 24727 5 1 1 24726
0 24728 7 1 2 88261 80175
0 24729 7 1 2 85853 24728
0 24730 5 1 1 24729
0 24731 7 1 2 24727 24730
0 24732 5 1 1 24731
0 24733 7 1 2 63966 24732
0 24734 5 1 1 24733
0 24735 7 1 2 64728 75359
0 24736 7 1 2 89682 24735
0 24737 5 1 1 24736
0 24738 7 1 2 24734 24737
0 24739 5 1 1 24738
0 24740 7 1 2 66482 24739
0 24741 5 1 1 24740
0 24742 7 1 2 69800 24741
0 24743 7 1 2 24725 24742
0 24744 5 1 1 24743
0 24745 7 1 2 87014 22889
0 24746 5 11 1 24745
0 24747 7 1 2 75480 96034
0 24748 5 1 1 24747
0 24749 7 1 2 70066 95848
0 24750 5 1 1 24749
0 24751 7 1 2 24748 24750
0 24752 5 1 1 24751
0 24753 7 1 2 96037 24752
0 24754 5 1 1 24753
0 24755 7 1 2 82742 87110
0 24756 5 1 1 24755
0 24757 7 1 2 91592 24756
0 24758 5 1 1 24757
0 24759 7 1 2 85202 24758
0 24760 5 1 1 24759
0 24761 7 1 2 85320 83591
0 24762 5 1 1 24761
0 24763 7 1 2 24760 24762
0 24764 5 1 1 24763
0 24765 7 1 2 66483 24764
0 24766 5 1 1 24765
0 24767 7 2 2 61573 82054
0 24768 7 1 2 83382 80878
0 24769 7 1 2 96048 24768
0 24770 5 1 1 24769
0 24771 7 1 2 24766 24770
0 24772 5 1 1 24771
0 24773 7 1 2 62102 24772
0 24774 5 1 1 24773
0 24775 7 1 2 24754 24774
0 24776 5 1 1 24775
0 24777 7 1 2 72882 24776
0 24778 5 1 1 24777
0 24779 7 2 2 88356 95817
0 24780 7 2 2 69563 96050
0 24781 7 1 2 66484 71699
0 24782 7 1 2 96052 24781
0 24783 5 1 1 24782
0 24784 7 1 2 82743 78729
0 24785 5 1 1 24784
0 24786 7 1 2 22305 24785
0 24787 5 2 1 24786
0 24788 7 1 2 90568 87885
0 24789 7 1 2 96054 24788
0 24790 5 1 1 24789
0 24791 7 1 2 24783 24790
0 24792 5 1 1 24791
0 24793 7 1 2 74117 24792
0 24794 5 1 1 24793
0 24795 7 1 2 82744 81249
0 24796 7 1 2 75360 24795
0 24797 5 1 1 24796
0 24798 7 2 2 61860 74358
0 24799 7 1 2 82546 96056
0 24800 7 1 2 96024 24799
0 24801 5 1 1 24800
0 24802 7 1 2 24797 24801
0 24803 5 1 1 24802
0 24804 7 1 2 89330 24803
0 24805 5 1 1 24804
0 24806 7 1 2 64935 24805
0 24807 7 1 2 24794 24806
0 24808 7 1 2 24778 24807
0 24809 5 1 1 24808
0 24810 7 1 2 68010 24809
0 24811 7 1 2 24744 24810
0 24812 5 1 1 24811
0 24813 7 1 2 24669 24812
0 24814 5 1 1 24813
0 24815 7 1 2 92768 24814
0 24816 5 1 1 24815
0 24817 7 2 2 63801 85895
0 24818 7 6 2 64345 64729
0 24819 7 1 2 79808 96060
0 24820 7 1 2 96058 24819
0 24821 7 1 2 92750 24820
0 24822 5 2 1 24821
0 24823 7 4 2 69191 69801
0 24824 7 7 2 79364 96068
0 24825 7 1 2 78193 72327
0 24826 7 1 2 96072 24825
0 24827 7 1 2 91795 24826
0 24828 5 1 1 24827
0 24829 7 1 2 96066 24828
0 24830 5 1 1 24829
0 24831 7 1 2 67683 24830
0 24832 5 1 1 24831
0 24833 7 2 2 80324 91279
0 24834 7 1 2 79740 87870
0 24835 7 1 2 96079 24834
0 24836 5 1 1 24835
0 24837 7 5 2 88459 82939
0 24838 7 1 2 76495 96057
0 24839 7 1 2 96081 24838
0 24840 5 1 1 24839
0 24841 7 1 2 24836 24840
0 24842 5 1 1 24841
0 24843 7 1 2 73007 24842
0 24844 5 1 1 24843
0 24845 7 4 2 67253 64518
0 24846 7 2 2 80272 96086
0 24847 7 4 2 66721 69192
0 24848 7 1 2 86262 79297
0 24849 7 1 2 96092 24848
0 24850 7 1 2 96090 24849
0 24851 5 1 1 24850
0 24852 7 1 2 24844 24851
0 24853 5 1 1 24852
0 24854 7 1 2 68171 24853
0 24855 5 1 1 24854
0 24856 7 1 2 78730 71700
0 24857 5 1 1 24856
0 24858 7 1 2 70701 88306
0 24859 5 1 1 24858
0 24860 7 1 2 24857 24859
0 24861 5 1 1 24860
0 24862 7 13 2 69564 93091
0 24863 7 1 2 73008 87562
0 24864 7 1 2 96096 24863
0 24865 7 1 2 24861 24864
0 24866 5 1 1 24865
0 24867 7 1 2 24855 24866
0 24868 5 1 1 24867
0 24869 7 1 2 66485 24868
0 24870 5 1 1 24869
0 24871 7 6 2 62841 64346
0 24872 7 1 2 95639 96109
0 24873 7 1 2 96051 24872
0 24874 5 1 1 24873
0 24875 7 1 2 63156 24874
0 24876 7 1 2 24870 24875
0 24877 5 1 1 24876
0 24878 7 1 2 79254 87579
0 24879 5 1 1 24878
0 24880 7 5 2 68172 68840
0 24881 7 1 2 88709 96115
0 24882 7 1 2 95986 24881
0 24883 5 1 1 24882
0 24884 7 1 2 24879 24883
0 24885 5 1 1 24884
0 24886 7 1 2 66722 24885
0 24887 5 1 1 24886
0 24888 7 1 2 84861 82457
0 24889 5 1 1 24888
0 24890 7 1 2 94870 24889
0 24891 5 1 1 24890
0 24892 7 1 2 77212 24891
0 24893 5 1 1 24892
0 24894 7 1 2 24887 24893
0 24895 5 1 1 24894
0 24896 7 1 2 68659 24895
0 24897 5 1 1 24896
0 24898 7 5 2 65744 83120
0 24899 7 2 2 71836 79255
0 24900 7 1 2 80694 96125
0 24901 7 1 2 96120 24900
0 24902 5 1 1 24901
0 24903 7 1 2 96032 24902
0 24904 7 1 2 24897 24903
0 24905 5 1 1 24904
0 24906 7 1 2 93033 24905
0 24907 5 1 1 24906
0 24908 7 1 2 78731 96011
0 24909 5 1 1 24908
0 24910 7 1 2 88649 73755
0 24911 5 1 1 24910
0 24912 7 1 2 24909 24911
0 24913 5 1 1 24912
0 24914 7 1 2 86925 93092
0 24915 7 1 2 91075 24914
0 24916 7 1 2 24913 24915
0 24917 5 1 1 24916
0 24918 7 1 2 68011 24917
0 24919 7 1 2 24907 24918
0 24920 5 1 1 24919
0 24921 7 1 2 24877 24920
0 24922 5 1 1 24921
0 24923 7 1 2 69802 24922
0 24924 5 1 1 24923
0 24925 7 1 2 74899 2748
0 24926 5 2 1 24925
0 24927 7 1 2 78929 96127
0 24928 5 1 1 24927
0 24929 7 2 2 89057 87886
0 24930 5 1 1 96129
0 24931 7 1 2 24928 24930
0 24932 5 1 1 24931
0 24933 7 1 2 83547 24932
0 24934 5 1 1 24933
0 24935 7 1 2 80771 91186
0 24936 7 1 2 83702 24935
0 24937 5 1 1 24936
0 24938 7 1 2 24934 24937
0 24939 5 1 1 24938
0 24940 7 1 2 62103 24939
0 24941 5 1 1 24940
0 24942 7 1 2 94874 96130
0 24943 5 1 1 24942
0 24944 7 1 2 66723 24943
0 24945 7 1 2 24941 24944
0 24946 5 1 1 24945
0 24947 7 1 2 83768 87887
0 24948 7 1 2 95815 24947
0 24949 5 1 1 24948
0 24950 7 1 2 89649 91202
0 24951 5 1 1 24950
0 24952 7 1 2 61861 24951
0 24953 7 1 2 24949 24952
0 24954 5 1 1 24953
0 24955 7 6 2 69193 94715
0 24956 7 1 2 24954 96131
0 24957 7 1 2 24946 24956
0 24958 5 1 1 24957
0 24959 7 10 2 69364 90956
0 24960 7 1 2 91539 96137
0 24961 7 1 2 96053 24960
0 24962 5 1 1 24961
0 24963 7 1 2 64936 24962
0 24964 7 1 2 24958 24963
0 24965 5 1 1 24964
0 24966 7 1 2 72625 24965
0 24967 7 1 2 24924 24966
0 24968 5 1 1 24967
0 24969 7 1 2 24832 24968
0 24970 7 1 2 24816 24969
0 24971 7 1 2 24636 24970
0 24972 5 1 1 24971
0 24973 7 1 2 62575 24972
0 24974 5 1 1 24973
0 24975 7 1 2 88778 87824
0 24976 7 1 2 83661 95459
0 24977 7 1 2 24975 24976
0 24978 5 1 1 24977
0 24979 7 1 2 96067 24978
0 24980 5 1 1 24979
0 24981 7 1 2 67684 24980
0 24982 5 1 1 24981
0 24983 7 2 2 69194 84436
0 24984 7 1 2 70067 92702
0 24985 5 1 1 24984
0 24986 7 2 2 75148 81302
0 24987 5 1 1 96149
0 24988 7 1 2 24985 24987
0 24989 5 1 1 24988
0 24990 7 2 2 79078 87451
0 24991 5 1 1 96151
0 24992 7 5 2 69803 72626
0 24993 7 1 2 83334 96153
0 24994 5 1 1 24993
0 24995 7 1 2 24991 24994
0 24996 5 1 1 24995
0 24997 7 1 2 24989 24996
0 24998 5 1 1 24997
0 24999 7 1 2 89482 95825
0 25000 5 1 1 24999
0 25001 7 3 2 66958 80099
0 25002 7 2 2 68173 73829
0 25003 7 1 2 96158 96161
0 25004 5 1 1 25003
0 25005 7 1 2 25000 25004
0 25006 5 1 1 25005
0 25007 7 1 2 71436 25006
0 25008 5 1 1 25007
0 25009 7 1 2 64128 89463
0 25010 5 1 1 25009
0 25011 7 1 2 25008 25010
0 25012 5 1 1 25011
0 25013 7 1 2 70068 25012
0 25014 5 1 1 25013
0 25015 7 1 2 24998 25014
0 25016 5 1 1 25015
0 25017 7 1 2 80978 25016
0 25018 5 1 1 25017
0 25019 7 2 2 76153 95826
0 25020 5 1 1 96163
0 25021 7 1 2 91181 96164
0 25022 7 1 2 95340 25021
0 25023 5 1 1 25022
0 25024 7 1 2 25018 25023
0 25025 5 1 1 25024
0 25026 7 1 2 96147 25025
0 25027 5 1 1 25026
0 25028 7 1 2 24982 25027
0 25029 5 1 1 25028
0 25030 7 1 2 71578 25029
0 25031 5 1 1 25030
0 25032 7 1 2 65424 25031
0 25033 7 1 2 24974 25032
0 25034 7 1 2 24544 25033
0 25035 7 1 2 24230 25034
0 25036 7 1 2 24074 25035
0 25037 5 1 1 25036
0 25038 7 1 2 79256 93034
0 25039 7 1 2 91630 25038
0 25040 5 1 1 25039
0 25041 7 1 2 61574 86660
0 25042 7 1 2 96082 25041
0 25043 5 1 1 25042
0 25044 7 1 2 25040 25043
0 25045 5 1 1 25044
0 25046 7 1 2 84361 25045
0 25047 5 1 1 25046
0 25048 7 3 2 92111 94716
0 25049 5 1 1 96165
0 25050 7 1 2 93563 96166
0 25051 5 1 1 25050
0 25052 7 5 2 61575 82809
0 25053 7 1 2 77966 93658
0 25054 7 1 2 96168 25053
0 25055 5 1 1 25054
0 25056 7 1 2 25051 25055
0 25057 5 1 1 25056
0 25058 7 1 2 77035 25057
0 25059 5 1 1 25058
0 25060 7 1 2 25047 25059
0 25061 5 1 1 25060
0 25062 7 1 2 63157 25061
0 25063 5 1 1 25062
0 25064 7 6 2 88996 92112
0 25065 5 1 1 96173
0 25066 7 6 2 88460 94820
0 25067 5 3 1 96179
0 25068 7 1 2 25065 96185
0 25069 5 1 1 25068
0 25070 7 1 2 61576 25069
0 25071 5 1 1 25070
0 25072 7 1 2 76088 93035
0 25073 5 1 1 25072
0 25074 7 1 2 25071 25073
0 25075 5 2 1 25074
0 25076 7 1 2 94998 96188
0 25077 5 1 1 25076
0 25078 7 2 2 82848 81127
0 25079 7 4 2 68012 69195
0 25080 7 1 2 74118 76577
0 25081 7 1 2 96192 25080
0 25082 7 1 2 96190 25081
0 25083 7 1 2 83720 25082
0 25084 5 1 1 25083
0 25085 7 1 2 25077 25084
0 25086 7 1 2 25063 25085
0 25087 5 1 1 25086
0 25088 7 1 2 62408 25087
0 25089 5 1 1 25088
0 25090 7 2 2 68841 83365
0 25091 5 1 1 96196
0 25092 7 1 2 74695 25091
0 25093 5 8 1 25092
0 25094 7 1 2 96198 96174
0 25095 5 1 1 25094
0 25096 7 2 2 88461 92288
0 25097 7 1 2 80333 96206
0 25098 5 1 1 25097
0 25099 7 1 2 25095 25098
0 25100 5 1 1 25099
0 25101 7 1 2 65745 25100
0 25102 5 1 1 25101
0 25103 7 1 2 72548 88439
0 25104 7 1 2 89668 92113
0 25105 7 1 2 25103 25104
0 25106 5 1 1 25105
0 25107 7 4 2 63158 82810
0 25108 7 1 2 72059 87854
0 25109 7 1 2 96208 25108
0 25110 5 1 1 25109
0 25111 7 1 2 25106 25110
0 25112 5 1 1 25111
0 25113 7 1 2 67454 25112
0 25114 5 1 1 25113
0 25115 7 2 2 78777 94821
0 25116 7 1 2 72273 88028
0 25117 7 1 2 96212 25116
0 25118 5 1 1 25117
0 25119 7 1 2 25114 25118
0 25120 7 1 2 25102 25119
0 25121 5 1 1 25120
0 25122 7 1 2 61577 25121
0 25123 5 1 1 25122
0 25124 7 3 2 65746 96199
0 25125 5 3 1 96214
0 25126 7 1 2 77285 96217
0 25127 5 1 1 25126
0 25128 7 1 2 91970 92769
0 25129 7 1 2 25127 25128
0 25130 5 1 1 25129
0 25131 7 1 2 25123 25130
0 25132 5 1 1 25131
0 25133 7 1 2 63568 25132
0 25134 5 1 1 25133
0 25135 7 1 2 82681 87922
0 25136 7 1 2 91975 25135
0 25137 7 1 2 96200 25136
0 25138 5 1 1 25137
0 25139 7 1 2 25134 25138
0 25140 5 2 1 25139
0 25141 7 1 2 67254 96220
0 25142 5 1 1 25141
0 25143 7 2 2 69565 86697
0 25144 7 1 2 76371 93093
0 25145 7 2 2 96222 25144
0 25146 7 1 2 82314 96224
0 25147 5 1 1 25146
0 25148 7 1 2 25142 25147
0 25149 5 1 1 25148
0 25150 7 1 2 70069 25149
0 25151 5 1 1 25150
0 25152 7 1 2 25089 25151
0 25153 5 1 1 25152
0 25154 7 1 2 63802 25153
0 25155 5 1 1 25154
0 25156 7 1 2 62409 96221
0 25157 5 1 1 25156
0 25158 7 1 2 80211 91843
0 25159 5 1 1 25158
0 25160 7 1 2 96186 25159
0 25161 5 1 1 25160
0 25162 7 1 2 61578 25161
0 25163 5 1 1 25162
0 25164 7 1 2 87404 95913
0 25165 5 1 1 25164
0 25166 7 1 2 25163 25165
0 25167 5 1 1 25166
0 25168 7 1 2 70702 94041
0 25169 5 1 1 25168
0 25170 7 3 2 78028 92398
0 25171 5 2 1 96226
0 25172 7 1 2 25169 96229
0 25173 5 1 1 25172
0 25174 7 1 2 25167 25173
0 25175 5 1 1 25174
0 25176 7 2 2 63967 92770
0 25177 7 1 2 91971 96231
0 25178 5 1 1 25177
0 25179 7 2 2 78698 95898
0 25180 5 1 1 96233
0 25181 7 7 2 68013 92771
0 25182 7 1 2 81069 96235
0 25183 5 1 1 25182
0 25184 7 1 2 25180 25183
0 25185 5 1 1 25184
0 25186 7 1 2 61579 25185
0 25187 5 1 1 25186
0 25188 7 1 2 25178 25187
0 25189 5 1 1 25188
0 25190 7 1 2 62576 25189
0 25191 5 1 1 25190
0 25192 7 2 2 88462 90861
0 25193 7 1 2 92097 96242
0 25194 5 1 1 25193
0 25195 7 1 2 25191 25194
0 25196 5 1 1 25195
0 25197 7 1 2 77989 25196
0 25198 5 1 1 25197
0 25199 7 1 2 25175 25198
0 25200 5 1 1 25199
0 25201 7 1 2 75033 25200
0 25202 5 1 1 25201
0 25203 7 1 2 25157 25202
0 25204 5 1 1 25203
0 25205 7 1 2 78239 25204
0 25206 5 1 1 25205
0 25207 7 6 2 65155 75771
0 25208 7 1 2 77496 76154
0 25209 5 1 1 25208
0 25210 7 1 2 9432 25209
0 25211 5 1 1 25210
0 25212 7 1 2 80007 25211
0 25213 5 1 1 25212
0 25214 7 1 2 76089 87947
0 25215 5 1 1 25214
0 25216 7 1 2 25213 25215
0 25217 5 1 1 25216
0 25218 7 1 2 93036 25217
0 25219 5 1 1 25218
0 25220 7 2 2 77244 73324
0 25221 7 1 2 88463 91645
0 25222 7 1 2 96250 25221
0 25223 5 1 1 25222
0 25224 7 1 2 25219 25223
0 25225 5 1 1 25224
0 25226 7 1 2 96244 25225
0 25227 5 1 1 25226
0 25228 7 1 2 66724 25227
0 25229 7 1 2 25206 25228
0 25230 7 1 2 25155 25229
0 25231 5 1 1 25230
0 25232 7 2 2 79752 96236
0 25233 7 1 2 77497 80018
0 25234 5 1 1 25233
0 25235 7 1 2 76347 77602
0 25236 5 1 1 25235
0 25237 7 1 2 25234 25236
0 25238 5 1 1 25237
0 25239 7 1 2 67255 25238
0 25240 5 1 1 25239
0 25241 7 1 2 81227 25240
0 25242 5 1 1 25241
0 25243 7 1 2 68416 25242
0 25244 5 1 1 25243
0 25245 7 4 2 86610 74036
0 25246 5 2 1 96254
0 25247 7 2 2 81198 95805
0 25248 5 1 1 96260
0 25249 7 1 2 73009 96261
0 25250 5 1 1 25249
0 25251 7 1 2 96258 25250
0 25252 7 1 2 25244 25251
0 25253 5 1 1 25252
0 25254 7 1 2 96252 25253
0 25255 5 1 1 25254
0 25256 7 2 2 65747 84811
0 25257 7 1 2 81199 80648
0 25258 7 1 2 96083 25257
0 25259 7 1 2 96262 25258
0 25260 5 1 1 25259
0 25261 7 1 2 25255 25260
0 25262 5 1 1 25261
0 25263 7 1 2 61580 25262
0 25264 5 1 1 25263
0 25265 7 1 2 68842 77315
0 25266 5 1 1 25265
0 25267 7 1 2 7104 25266
0 25268 5 4 1 25267
0 25269 7 1 2 79057 96264
0 25270 5 1 1 25269
0 25271 7 1 2 25270 96259
0 25272 5 1 1 25271
0 25273 7 1 2 88400 25272
0 25274 5 1 1 25273
0 25275 7 1 2 81344 80091
0 25276 7 1 2 82768 25275
0 25277 5 1 1 25276
0 25278 7 1 2 25274 25277
0 25279 5 1 1 25278
0 25280 7 1 2 96132 25279
0 25281 5 1 1 25280
0 25282 7 1 2 61862 25281
0 25283 7 1 2 25264 25282
0 25284 5 1 1 25283
0 25285 7 1 2 25231 25284
0 25286 5 1 1 25285
0 25287 7 1 2 64937 25286
0 25288 5 1 1 25287
0 25289 7 1 2 63968 85307
0 25290 5 1 1 25289
0 25291 7 2 2 79399 25290
0 25292 5 1 1 96268
0 25293 7 1 2 62577 25292
0 25294 5 1 1 25293
0 25295 7 2 2 73978 25294
0 25296 5 3 1 96270
0 25297 7 1 2 66959 96271
0 25298 5 4 1 25297
0 25299 7 1 2 74807 96275
0 25300 5 1 1 25299
0 25301 7 2 2 80762 96201
0 25302 5 1 1 96279
0 25303 7 1 2 25300 25302
0 25304 5 1 1 25303
0 25305 7 1 2 65156 25304
0 25306 5 1 1 25305
0 25307 7 1 2 4848 25306
0 25308 5 1 1 25307
0 25309 7 1 2 89340 25308
0 25310 5 1 1 25309
0 25311 7 4 2 65748 74359
0 25312 7 1 2 96202 96281
0 25313 5 1 1 25312
0 25314 7 1 2 77288 25313
0 25315 5 1 1 25314
0 25316 7 1 2 73010 25315
0 25317 5 1 1 25316
0 25318 7 1 2 83614 96272
0 25319 5 1 1 25318
0 25320 7 1 2 25317 25319
0 25321 5 1 1 25320
0 25322 7 1 2 83335 25321
0 25323 5 1 1 25322
0 25324 7 2 2 71233 76348
0 25325 5 4 1 96285
0 25326 7 1 2 74843 96287
0 25327 5 1 1 25326
0 25328 7 1 2 78778 95194
0 25329 7 1 2 25327 25328
0 25330 5 1 1 25329
0 25331 7 1 2 70070 25330
0 25332 7 1 2 25323 25331
0 25333 5 1 1 25332
0 25334 7 3 2 77641 80008
0 25335 5 1 1 96291
0 25336 7 1 2 83336 96292
0 25337 5 1 1 25336
0 25338 7 1 2 66725 80909
0 25339 7 1 2 87890 25338
0 25340 7 1 2 80020 25339
0 25341 5 1 1 25340
0 25342 7 1 2 25337 25341
0 25343 5 1 1 25342
0 25344 7 1 2 72787 25343
0 25345 5 1 1 25344
0 25346 7 1 2 83337 77642
0 25347 5 1 1 25346
0 25348 7 1 2 88509 78266
0 25349 5 1 1 25348
0 25350 7 1 2 25347 25349
0 25351 5 1 1 25350
0 25352 7 1 2 87948 25351
0 25353 5 1 1 25352
0 25354 7 1 2 25345 25353
0 25355 5 1 1 25354
0 25356 7 1 2 70919 25355
0 25357 5 1 1 25356
0 25358 7 1 2 87949 95270
0 25359 7 1 2 88398 25358
0 25360 5 1 1 25359
0 25361 7 1 2 65157 25360
0 25362 7 1 2 25357 25361
0 25363 5 1 1 25362
0 25364 7 1 2 66486 25363
0 25365 7 1 2 25333 25364
0 25366 5 1 1 25365
0 25367 7 1 2 25310 25366
0 25368 5 1 1 25367
0 25369 7 1 2 92772 25368
0 25370 5 1 1 25369
0 25371 7 1 2 73721 13407
0 25372 5 3 1 25371
0 25373 7 2 2 65749 96294
0 25374 5 1 1 96297
0 25375 7 1 2 63569 75895
0 25376 5 1 1 25375
0 25377 7 1 2 25374 25376
0 25378 5 3 1 25377
0 25379 7 1 2 72549 96299
0 25380 5 1 1 25379
0 25381 7 4 2 68843 74402
0 25382 5 1 1 96302
0 25383 7 1 2 72060 96303
0 25384 5 1 1 25383
0 25385 7 1 2 25380 25384
0 25386 5 1 1 25385
0 25387 7 1 2 73011 25386
0 25388 5 1 1 25387
0 25389 7 2 2 83615 93564
0 25390 5 1 1 96306
0 25391 7 1 2 62410 75191
0 25392 5 3 1 25391
0 25393 7 1 2 25390 96308
0 25394 7 1 2 25388 25393
0 25395 5 1 1 25394
0 25396 7 1 2 70071 25395
0 25397 5 1 1 25396
0 25398 7 1 2 74296 93560
0 25399 5 1 1 25398
0 25400 7 2 2 77643 25399
0 25401 5 1 1 96311
0 25402 7 1 2 65158 96312
0 25403 5 1 1 25402
0 25404 7 1 2 80717 79023
0 25405 5 1 1 25404
0 25406 7 2 2 62104 80009
0 25407 7 1 2 25405 96313
0 25408 5 1 1 25407
0 25409 7 2 2 77719 79591
0 25410 5 1 1 96315
0 25411 7 1 2 71234 93482
0 25412 5 1 1 25411
0 25413 7 1 2 25410 25412
0 25414 5 1 1 25413
0 25415 7 1 2 63570 25414
0 25416 5 1 1 25415
0 25417 7 1 2 25408 25416
0 25418 5 1 1 25417
0 25419 7 1 2 84362 25418
0 25420 5 1 1 25419
0 25421 7 1 2 25403 25420
0 25422 7 1 2 25397 25421
0 25423 5 1 1 25422
0 25424 7 1 2 83292 96097
0 25425 7 1 2 25423 25424
0 25426 5 1 1 25425
0 25427 7 1 2 68014 25426
0 25428 7 1 2 25370 25427
0 25429 5 1 1 25428
0 25430 7 1 2 90236 94233
0 25431 7 1 2 96263 25430
0 25432 5 1 1 25431
0 25433 7 1 2 75381 77198
0 25434 7 1 2 89497 25433
0 25435 5 1 1 25434
0 25436 7 1 2 25432 25435
0 25437 5 1 1 25436
0 25438 7 1 2 68844 25437
0 25439 5 1 1 25438
0 25440 7 1 2 72421 95327
0 25441 7 1 2 88881 25440
0 25442 5 1 1 25441
0 25443 7 1 2 25439 25442
0 25444 5 1 1 25443
0 25445 7 1 2 67455 25444
0 25446 5 1 1 25445
0 25447 7 1 2 81173 18908
0 25448 5 1 1 25447
0 25449 7 1 2 71330 25448
0 25450 5 1 1 25449
0 25451 7 1 2 94322 95711
0 25452 5 1 1 25451
0 25453 7 1 2 25450 25452
0 25454 5 1 1 25453
0 25455 7 1 2 62105 25454
0 25456 5 1 1 25455
0 25457 7 1 2 76259 75335
0 25458 5 1 1 25457
0 25459 7 1 2 25456 25458
0 25460 5 1 1 25459
0 25461 7 1 2 67256 25460
0 25462 5 1 1 25461
0 25463 7 1 2 72550 71491
0 25464 7 1 2 96298 25463
0 25465 5 1 1 25464
0 25466 7 1 2 96309 25465
0 25467 7 1 2 25462 25466
0 25468 5 1 1 25467
0 25469 7 1 2 77199 25468
0 25470 5 1 1 25469
0 25471 7 1 2 25446 25470
0 25472 5 1 1 25471
0 25473 7 1 2 70072 25472
0 25474 5 1 1 25473
0 25475 7 1 2 15468 25335
0 25476 5 1 1 25475
0 25477 7 1 2 84363 25476
0 25478 5 2 1 25477
0 25479 7 1 2 25401 96317
0 25480 5 1 1 25479
0 25481 7 1 2 89043 25480
0 25482 5 1 1 25481
0 25483 7 1 2 25474 25482
0 25484 5 1 1 25483
0 25485 7 1 2 69566 25484
0 25486 5 1 1 25485
0 25487 7 1 2 7036 78252
0 25488 5 2 1 25487
0 25489 7 1 2 75721 96319
0 25490 5 1 1 25489
0 25491 7 1 2 86815 73325
0 25492 5 1 1 25491
0 25493 7 1 2 25490 25492
0 25494 5 1 1 25493
0 25495 7 1 2 84364 25494
0 25496 5 1 1 25495
0 25497 7 1 2 79028 93565
0 25498 5 1 1 25497
0 25499 7 1 2 71837 78110
0 25500 5 1 1 25499
0 25501 7 1 2 25498 25500
0 25502 7 1 2 25496 25501
0 25503 5 1 1 25502
0 25504 7 1 2 62106 25503
0 25505 5 1 1 25504
0 25506 7 1 2 86711 91928
0 25507 5 1 1 25506
0 25508 7 1 2 74514 91408
0 25509 5 1 1 25508
0 25510 7 1 2 85712 74515
0 25511 5 1 1 25510
0 25512 7 1 2 76628 25511
0 25513 5 1 1 25512
0 25514 7 1 2 62411 25513
0 25515 5 1 1 25514
0 25516 7 1 2 25509 25515
0 25517 7 1 2 25507 25516
0 25518 5 1 1 25517
0 25519 7 1 2 70073 25518
0 25520 5 1 1 25519
0 25521 7 1 2 71956 93561
0 25522 5 1 1 25521
0 25523 7 1 2 77036 25522
0 25524 5 1 1 25523
0 25525 7 1 2 25520 25524
0 25526 5 1 1 25525
0 25527 7 1 2 63571 25526
0 25528 5 1 1 25527
0 25529 7 1 2 77451 91696
0 25530 7 1 2 94167 25529
0 25531 5 1 1 25530
0 25532 7 1 2 25528 25531
0 25533 7 1 2 25505 25532
0 25534 5 1 1 25533
0 25535 7 1 2 91580 25534
0 25536 5 1 1 25535
0 25537 7 1 2 25486 25536
0 25538 5 1 1 25537
0 25539 7 1 2 93094 25538
0 25540 5 1 1 25539
0 25541 7 1 2 83457 96093
0 25542 7 1 2 95123 25541
0 25543 7 1 2 96280 25542
0 25544 5 1 1 25543
0 25545 7 1 2 63159 25544
0 25546 7 1 2 25540 25545
0 25547 5 1 1 25546
0 25548 7 1 2 25429 25547
0 25549 5 1 1 25548
0 25550 7 1 2 69804 25549
0 25551 5 1 1 25550
0 25552 7 1 2 68174 25551
0 25553 7 1 2 25288 25552
0 25554 5 1 1 25553
0 25555 7 4 2 66960 74866
0 25556 5 1 1 96321
0 25557 7 1 2 79291 92022
0 25558 5 1 1 25557
0 25559 7 1 2 83319 25558
0 25560 5 1 1 25559
0 25561 7 1 2 96322 25560
0 25562 5 1 1 25561
0 25563 7 1 2 71101 87588
0 25564 5 1 1 25563
0 25565 7 1 2 25562 25564
0 25566 5 1 1 25565
0 25567 7 1 2 63160 25566
0 25568 5 1 1 25567
0 25569 7 1 2 74867 84474
0 25570 7 1 2 86366 25569
0 25571 5 1 1 25570
0 25572 7 1 2 25568 25571
0 25573 5 1 1 25572
0 25574 7 1 2 71235 25573
0 25575 5 1 1 25574
0 25576 7 2 2 76155 96295
0 25577 7 1 2 73012 71098
0 25578 7 1 2 96325 25577
0 25579 5 1 1 25578
0 25580 7 1 2 25575 25579
0 25581 5 1 1 25580
0 25582 7 1 2 65750 25581
0 25583 5 1 1 25582
0 25584 7 1 2 73013 89029
0 25585 5 1 1 25584
0 25586 7 1 2 82453 92759
0 25587 5 1 1 25586
0 25588 7 1 2 25585 25587
0 25589 5 1 1 25588
0 25590 7 1 2 88362 72422
0 25591 7 1 2 25589 25590
0 25592 5 1 1 25591
0 25593 7 1 2 25583 25592
0 25594 5 1 1 25593
0 25595 7 1 2 65988 25594
0 25596 5 1 1 25595
0 25597 7 1 2 3668 25382
0 25598 5 1 1 25597
0 25599 7 1 2 67257 82532
0 25600 7 1 2 25598 25599
0 25601 5 1 1 25600
0 25602 7 1 2 77515 82528
0 25603 5 1 1 25602
0 25604 7 1 2 25601 25603
0 25605 5 1 1 25604
0 25606 7 1 2 69805 25605
0 25607 5 1 1 25606
0 25608 7 1 2 77089 87437
0 25609 7 1 2 83721 25608
0 25610 5 1 1 25609
0 25611 7 1 2 25607 25610
0 25612 5 1 1 25611
0 25613 7 1 2 66726 25612
0 25614 5 1 1 25613
0 25615 7 1 2 88280 95988
0 25616 7 1 2 79864 25615
0 25617 5 1 1 25616
0 25618 7 1 2 25614 25617
0 25619 5 1 1 25618
0 25620 7 1 2 76156 25619
0 25621 5 1 1 25620
0 25622 7 2 2 77775 85551
0 25623 5 1 1 96327
0 25624 7 2 2 77200 77149
0 25625 7 1 2 89617 96329
0 25626 7 1 2 96328 25625
0 25627 5 1 1 25626
0 25628 7 1 2 25621 25627
0 25629 5 1 1 25628
0 25630 7 1 2 84365 25629
0 25631 5 1 1 25630
0 25632 7 1 2 75703 94287
0 25633 5 1 1 25632
0 25634 7 1 2 90467 80010
0 25635 5 1 1 25634
0 25636 7 1 2 25633 25635
0 25637 5 1 1 25636
0 25638 7 1 2 72061 25637
0 25639 5 1 1 25638
0 25640 7 1 2 90468 87950
0 25641 5 1 1 25640
0 25642 7 1 2 25639 25641
0 25643 5 1 1 25642
0 25644 7 1 2 63803 25643
0 25645 5 1 1 25644
0 25646 7 1 2 75704 91225
0 25647 5 1 1 25646
0 25648 7 1 2 25645 25647
0 25649 5 1 1 25648
0 25650 7 1 2 90072 25649
0 25651 5 1 1 25650
0 25652 7 3 2 69806 79283
0 25653 7 1 2 96330 96331
0 25654 7 1 2 93566 25653
0 25655 5 1 1 25654
0 25656 7 1 2 25651 25655
0 25657 5 1 1 25656
0 25658 7 1 2 63572 25657
0 25659 5 1 1 25658
0 25660 7 1 2 25631 25659
0 25661 7 1 2 25596 25660
0 25662 5 1 1 25661
0 25663 7 1 2 69567 25662
0 25664 5 1 1 25663
0 25665 7 1 2 85082 95410
0 25666 5 1 1 25665
0 25667 7 3 2 75664 25666
0 25668 5 2 1 96334
0 25669 7 2 2 64730 74277
0 25670 7 1 2 77150 96339
0 25671 7 1 2 95879 25670
0 25672 7 1 2 96337 25671
0 25673 5 1 1 25672
0 25674 7 1 2 70074 25673
0 25675 7 1 2 25664 25674
0 25676 5 1 1 25675
0 25677 7 1 2 74321 95015
0 25678 5 1 1 25677
0 25679 7 1 2 77690 87148
0 25680 5 1 1 25679
0 25681 7 1 2 64129 89827
0 25682 5 1 1 25681
0 25683 7 1 2 25680 25682
0 25684 5 1 1 25683
0 25685 7 1 2 63573 25684
0 25686 5 1 1 25685
0 25687 7 5 2 71331 72788
0 25688 5 1 1 96341
0 25689 7 1 2 84928 25688
0 25690 7 1 2 79994 25689
0 25691 5 1 1 25690
0 25692 7 1 2 74360 71056
0 25693 7 1 2 25691 25692
0 25694 5 1 1 25693
0 25695 7 1 2 25686 25694
0 25696 5 1 1 25695
0 25697 7 1 2 70920 25696
0 25698 5 1 1 25697
0 25699 7 1 2 75750 87454
0 25700 5 1 1 25699
0 25701 7 1 2 25698 25700
0 25702 5 1 1 25701
0 25703 7 1 2 78884 25702
0 25704 5 1 1 25703
0 25705 7 1 2 25678 25704
0 25706 5 1 1 25705
0 25707 7 1 2 61581 25706
0 25708 5 1 1 25707
0 25709 7 2 2 81471 92023
0 25710 7 2 2 66727 80011
0 25711 7 1 2 77510 96348
0 25712 5 1 1 25711
0 25713 7 1 2 75833 25712
0 25714 5 1 1 25713
0 25715 7 1 2 96346 25714
0 25716 5 1 1 25715
0 25717 7 1 2 25708 25716
0 25718 5 1 1 25717
0 25719 7 1 2 71838 25718
0 25720 5 1 1 25719
0 25721 7 1 2 73458 76514
0 25722 5 1 1 25721
0 25723 7 1 2 71332 92727
0 25724 7 1 2 25722 25723
0 25725 5 1 1 25724
0 25726 7 3 2 61582 76996
0 25727 7 1 2 80325 78815
0 25728 7 1 2 96350 25727
0 25729 5 1 1 25728
0 25730 7 2 2 74119 81922
0 25731 5 1 1 96353
0 25732 7 1 2 71460 85083
0 25733 7 1 2 96354 25732
0 25734 5 1 1 25733
0 25735 7 1 2 25729 25734
0 25736 7 1 2 25725 25735
0 25737 5 1 1 25736
0 25738 7 1 2 75772 91453
0 25739 7 1 2 25737 25738
0 25740 5 1 1 25739
0 25741 7 1 2 65159 25740
0 25742 7 1 2 25720 25741
0 25743 5 1 1 25742
0 25744 7 1 2 69365 25743
0 25745 7 1 2 25676 25744
0 25746 5 1 1 25745
0 25747 7 1 2 72159 71526
0 25748 5 1 1 25747
0 25749 7 1 2 62842 25748
0 25750 5 1 1 25749
0 25751 7 1 2 85582 25750
0 25752 5 1 1 25751
0 25753 7 1 2 62578 25752
0 25754 5 1 1 25753
0 25755 7 1 2 96269 25754
0 25756 5 1 1 25755
0 25757 7 1 2 90853 92523
0 25758 7 1 2 25756 25757
0 25759 5 1 1 25758
0 25760 7 1 2 25746 25759
0 25761 5 1 1 25760
0 25762 7 1 2 64347 25761
0 25763 5 1 1 25762
0 25764 7 2 2 78951 96286
0 25765 5 1 1 96355
0 25766 7 1 2 17560 25765
0 25767 5 1 1 25766
0 25768 7 1 2 82622 25767
0 25769 5 1 1 25768
0 25770 7 1 2 68417 96335
0 25771 5 1 1 25770
0 25772 7 1 2 95179 25771
0 25773 5 1 1 25772
0 25774 7 1 2 25769 25773
0 25775 5 1 1 25774
0 25776 7 1 2 63804 25775
0 25777 5 1 1 25776
0 25778 7 1 2 88367 86860
0 25779 5 1 1 25778
0 25780 7 1 2 77316 84111
0 25781 5 1 1 25780
0 25782 7 1 2 25779 25781
0 25783 5 1 1 25782
0 25784 7 1 2 72551 25783
0 25785 5 1 1 25784
0 25786 7 6 2 62579 71527
0 25787 5 2 1 96357
0 25788 7 2 2 72627 96358
0 25789 5 1 1 96365
0 25790 7 1 2 80354 96366
0 25791 5 1 1 25790
0 25792 7 1 2 25785 25791
0 25793 5 1 1 25792
0 25794 7 1 2 87427 25793
0 25795 5 1 1 25794
0 25796 7 1 2 25777 25795
0 25797 5 1 1 25796
0 25798 7 1 2 62412 25797
0 25799 5 1 1 25798
0 25800 7 2 2 81681 74223
0 25801 5 1 1 96367
0 25802 7 1 2 96338 96368
0 25803 5 1 1 25802
0 25804 7 1 2 80521 89595
0 25805 7 1 2 94234 25804
0 25806 7 1 2 96265 25805
0 25807 5 1 1 25806
0 25808 7 1 2 25803 25807
0 25809 5 1 1 25808
0 25810 7 1 2 64731 25809
0 25811 5 1 1 25810
0 25812 7 1 2 65751 89304
0 25813 7 2 2 84668 25812
0 25814 7 2 2 69568 74037
0 25815 7 2 2 78759 82160
0 25816 7 1 2 96371 96373
0 25817 7 1 2 96369 25816
0 25818 5 1 1 25817
0 25819 7 1 2 25811 25818
0 25820 7 1 2 25799 25819
0 25821 5 1 1 25820
0 25822 7 1 2 64938 25821
0 25823 5 1 1 25822
0 25824 7 1 2 73916 96203
0 25825 5 1 1 25824
0 25826 7 1 2 86408 82506
0 25827 5 1 1 25826
0 25828 7 1 2 25825 25827
0 25829 5 1 1 25828
0 25830 7 1 2 62413 25829
0 25831 5 1 1 25830
0 25832 7 1 2 91991 96204
0 25833 5 1 1 25832
0 25834 7 1 2 25831 25833
0 25835 5 1 1 25834
0 25836 7 1 2 95040 25835
0 25837 5 1 1 25836
0 25838 7 2 2 76467 76504
0 25839 7 1 2 86820 96375
0 25840 5 1 1 25839
0 25841 7 1 2 25837 25840
0 25842 5 1 1 25841
0 25843 7 1 2 78974 25842
0 25844 5 1 1 25843
0 25845 7 1 2 25823 25844
0 25846 5 1 1 25845
0 25847 7 1 2 66487 25846
0 25848 5 1 1 25847
0 25849 7 1 2 76349 86649
0 25850 5 1 1 25849
0 25851 7 1 2 25248 25850
0 25852 5 1 1 25851
0 25853 7 1 2 73014 25852
0 25854 5 1 1 25853
0 25855 7 1 2 63574 96288
0 25856 5 1 1 25855
0 25857 7 1 2 86628 25856
0 25858 5 1 1 25857
0 25859 7 1 2 25854 25858
0 25860 5 1 1 25859
0 25861 7 1 2 78994 25860
0 25862 5 1 1 25861
0 25863 7 1 2 65160 25862
0 25864 7 1 2 25848 25863
0 25865 5 1 1 25864
0 25866 7 2 2 65989 96323
0 25867 7 3 2 71528 95369
0 25868 5 1 1 96379
0 25869 7 1 2 91976 96380
0 25870 7 1 2 96377 25869
0 25871 5 1 1 25870
0 25872 7 2 2 68015 79257
0 25873 7 1 2 91544 96382
0 25874 7 1 2 96273 25873
0 25875 5 1 1 25874
0 25876 7 1 2 25871 25875
0 25877 5 1 1 25876
0 25878 7 1 2 66728 25877
0 25879 5 1 1 25878
0 25880 7 1 2 64732 80443
0 25881 7 1 2 88564 25880
0 25882 5 1 1 25881
0 25883 7 1 2 25879 25882
0 25884 5 1 1 25883
0 25885 7 1 2 64939 25884
0 25886 5 1 1 25885
0 25887 7 1 2 71693 83891
0 25888 7 1 2 85236 25887
0 25889 7 1 2 85799 95395
0 25890 7 1 2 25888 25889
0 25891 5 1 1 25890
0 25892 7 1 2 70075 25891
0 25893 7 1 2 25886 25892
0 25894 5 1 1 25893
0 25895 7 1 2 92773 25894
0 25896 7 1 2 25865 25895
0 25897 5 1 1 25896
0 25898 7 1 2 25763 25897
0 25899 5 1 1 25898
0 25900 7 1 2 63335 25899
0 25901 5 1 1 25900
0 25902 7 1 2 70343 25901
0 25903 7 1 2 25554 25902
0 25904 5 1 1 25903
0 25905 7 1 2 25037 25904
0 25906 5 1 1 25905
0 25907 7 4 2 80787 96138
0 25908 5 1 1 96384
0 25909 7 1 2 87994 96385
0 25910 5 1 1 25909
0 25911 7 8 2 80979 92774
0 25912 7 1 2 76445 96388
0 25913 5 1 1 25912
0 25914 7 1 2 25910 25913
0 25915 5 1 1 25914
0 25916 7 1 2 70344 25915
0 25917 5 1 1 25916
0 25918 7 2 2 66488 80033
0 25919 7 1 2 93734 94785
0 25920 7 1 2 96396 25919
0 25921 5 1 1 25920
0 25922 7 1 2 25917 25921
0 25923 5 1 1 25922
0 25924 7 1 2 67456 25923
0 25925 5 1 1 25924
0 25926 7 1 2 68418 80889
0 25927 7 1 2 96389 25926
0 25928 5 1 1 25927
0 25929 7 1 2 25925 25928
0 25930 5 1 1 25929
0 25931 7 1 2 65752 25930
0 25932 5 1 1 25931
0 25933 7 2 2 85475 85698
0 25934 5 1 1 96398
0 25935 7 1 2 96399 96386
0 25936 5 1 1 25935
0 25937 7 2 2 67258 69196
0 25938 7 2 2 88997 96400
0 25939 7 1 2 88336 75918
0 25940 7 1 2 96402 25939
0 25941 5 1 1 25940
0 25942 7 1 2 25936 25941
0 25943 7 1 2 25932 25942
0 25944 5 1 1 25943
0 25945 7 1 2 66961 25944
0 25946 5 1 1 25945
0 25947 7 1 2 75956 75110
0 25948 5 2 1 25947
0 25949 7 3 2 66962 85681
0 25950 5 1 1 96406
0 25951 7 1 2 84171 96407
0 25952 5 1 1 25951
0 25953 7 1 2 96404 25952
0 25954 5 1 1 25953
0 25955 7 1 2 67259 25954
0 25956 5 1 1 25955
0 25957 7 1 2 70345 82769
0 25958 5 1 1 25957
0 25959 7 1 2 25956 25958
0 25960 5 1 1 25959
0 25961 7 1 2 93015 95252
0 25962 5 1 1 25961
0 25963 7 1 2 25908 25962
0 25964 5 1 1 25963
0 25965 7 1 2 65753 25964
0 25966 7 1 2 25960 25965
0 25967 5 1 1 25966
0 25968 7 1 2 25946 25967
0 25969 5 1 1 25968
0 25970 7 1 2 71437 25969
0 25971 5 1 1 25970
0 25972 7 2 2 70346 82186
0 25973 5 1 1 96409
0 25974 7 1 2 74003 25973
0 25975 5 1 1 25974
0 25976 7 6 2 67685 69197
0 25977 7 4 2 64519 96411
0 25978 7 1 2 82169 96417
0 25979 7 1 2 92682 25978
0 25980 7 1 2 25975 25979
0 25981 5 1 1 25980
0 25982 7 1 2 25971 25981
0 25983 5 1 1 25982
0 25984 7 1 2 68175 25983
0 25985 5 1 1 25984
0 25986 7 1 2 87659 92593
0 25987 7 1 2 93147 25986
0 25988 7 1 2 93493 25987
0 25989 5 1 1 25988
0 25990 7 1 2 69569 25989
0 25991 7 1 2 25985 25990
0 25992 5 1 1 25991
0 25993 7 1 2 91099 93298
0 25994 5 1 1 25993
0 25995 7 2 2 76468 25994
0 25996 7 1 2 68176 96421
0 25997 5 1 1 25996
0 25998 7 2 2 84862 86192
0 25999 5 1 1 96423
0 26000 7 1 2 25997 25999
0 26001 5 1 1 26000
0 26002 7 1 2 62107 26001
0 26003 5 1 1 26002
0 26004 7 1 2 70347 84978
0 26005 5 2 1 26004
0 26006 7 1 2 86422 96425
0 26007 5 1 1 26006
0 26008 7 1 2 84787 26007
0 26009 5 1 1 26008
0 26010 7 1 2 26003 26009
0 26011 5 2 1 26010
0 26012 7 3 2 93192 94822
0 26013 7 1 2 96427 96429
0 26014 5 1 1 26013
0 26015 7 6 2 69198 65425
0 26016 7 1 2 67686 95989
0 26017 7 1 2 96432 26016
0 26018 7 2 2 64520 81816
0 26019 7 1 2 79206 96438
0 26020 7 1 2 26017 26019
0 26021 5 1 1 26020
0 26022 7 1 2 26014 26021
0 26023 5 1 1 26022
0 26024 7 1 2 61583 26023
0 26025 5 1 1 26024
0 26026 7 1 2 64940 74465
0 26027 7 1 2 95932 26026
0 26028 7 1 2 96422 26027
0 26029 5 1 1 26028
0 26030 7 1 2 26025 26029
0 26031 5 1 1 26030
0 26032 7 1 2 65754 26031
0 26033 5 1 1 26032
0 26034 7 2 2 63336 64348
0 26035 7 1 2 91515 96440
0 26036 7 1 2 92065 26035
0 26037 5 1 1 26036
0 26038 7 2 2 68177 64521
0 26039 7 11 2 69199 64941
0 26040 7 1 2 96442 96444
0 26041 7 1 2 93397 26040
0 26042 5 1 1 26041
0 26043 7 1 2 26037 26042
0 26044 5 1 1 26043
0 26045 7 1 2 85699 26044
0 26046 5 1 1 26045
0 26047 7 1 2 81534 96445
0 26048 7 1 2 84684 26047
0 26049 7 1 2 91759 26048
0 26050 5 1 1 26049
0 26051 7 1 2 26046 26050
0 26052 5 1 1 26051
0 26053 7 1 2 70703 75575
0 26054 7 1 2 26052 26053
0 26055 5 1 1 26054
0 26056 7 1 2 26033 26055
0 26057 5 1 1 26056
0 26058 7 1 2 61863 26057
0 26059 5 1 1 26058
0 26060 7 1 2 67457 85700
0 26061 5 1 1 26060
0 26062 7 1 2 84685 75434
0 26063 5 1 1 26062
0 26064 7 1 2 26061 26063
0 26065 5 3 1 26064
0 26066 7 3 2 74969 92775
0 26067 7 1 2 88553 91761
0 26068 7 1 2 96458 26067
0 26069 7 1 2 96455 26068
0 26070 5 1 1 26069
0 26071 7 1 2 64733 26070
0 26072 7 1 2 26059 26071
0 26073 5 1 1 26072
0 26074 7 1 2 70076 26073
0 26075 7 1 2 25992 26074
0 26076 5 1 1 26075
0 26077 7 1 2 81303 96266
0 26078 5 1 1 26077
0 26079 7 3 2 70077 96300
0 26080 7 1 2 68178 96461
0 26081 5 1 1 26080
0 26082 7 1 2 26078 26081
0 26083 5 1 1 26082
0 26084 7 1 2 66729 26083
0 26085 5 1 1 26084
0 26086 7 1 2 77331 75419
0 26087 7 1 2 96116 26086
0 26088 5 1 1 26087
0 26089 7 1 2 26085 26088
0 26090 5 1 1 26089
0 26091 7 1 2 63161 26090
0 26092 5 1 1 26091
0 26093 7 1 2 90173 96462
0 26094 5 1 1 26093
0 26095 7 1 2 26092 26094
0 26096 5 1 1 26095
0 26097 7 1 2 61584 26096
0 26098 5 1 1 26097
0 26099 7 1 2 88872 83679
0 26100 7 1 2 96301 26099
0 26101 5 1 1 26100
0 26102 7 1 2 26098 26101
0 26103 5 1 1 26102
0 26104 7 1 2 96098 26103
0 26105 5 1 1 26104
0 26106 7 2 2 84344 93037
0 26107 7 1 2 83691 96267
0 26108 7 1 2 96464 26107
0 26109 5 1 1 26108
0 26110 7 1 2 26105 26109
0 26111 5 1 1 26110
0 26112 7 1 2 70348 26111
0 26113 5 1 1 26112
0 26114 7 2 2 80936 95914
0 26115 5 1 1 96466
0 26116 7 1 2 80226 91844
0 26117 5 1 1 26116
0 26118 7 1 2 96187 26117
0 26119 5 3 1 26118
0 26120 7 1 2 61585 96468
0 26121 5 1 1 26120
0 26122 7 1 2 26115 26121
0 26123 5 1 1 26122
0 26124 7 2 2 80772 76706
0 26125 7 1 2 81453 74403
0 26126 7 1 2 96471 26125
0 26127 7 1 2 26123 26126
0 26128 5 1 1 26127
0 26129 7 1 2 64942 26128
0 26130 7 1 2 26113 26129
0 26131 5 1 1 26130
0 26132 7 1 2 67458 94085
0 26133 5 1 1 26132
0 26134 7 1 2 94647 26133
0 26135 5 1 1 26134
0 26136 7 1 2 8433 26135
0 26137 5 1 1 26136
0 26138 7 1 2 18212 94086
0 26139 5 1 1 26138
0 26140 7 1 2 81304 26139
0 26141 7 1 2 26137 26140
0 26142 5 1 1 26141
0 26143 7 1 2 77271 1985
0 26144 5 1 1 26143
0 26145 7 5 2 88387 26144
0 26146 7 2 2 70349 83548
0 26147 7 1 2 96296 96478
0 26148 7 1 2 96473 26147
0 26149 5 1 1 26148
0 26150 7 1 2 26142 26149
0 26151 5 1 1 26150
0 26152 7 1 2 61864 26151
0 26153 5 1 1 26152
0 26154 7 1 2 91270 94504
0 26155 5 1 1 26154
0 26156 7 1 2 70078 87202
0 26157 7 1 2 96326 26156
0 26158 5 1 1 26157
0 26159 7 1 2 26155 26158
0 26160 5 1 1 26159
0 26161 7 1 2 70350 78267
0 26162 7 1 2 26160 26161
0 26163 5 1 1 26162
0 26164 7 1 2 26153 26163
0 26165 5 1 1 26164
0 26166 7 1 2 65755 26165
0 26167 5 1 1 26166
0 26168 7 1 2 83338 91271
0 26169 5 1 1 26168
0 26170 7 1 2 88189 86112
0 26171 5 1 1 26170
0 26172 7 1 2 26169 26171
0 26173 5 1 1 26172
0 26174 7 1 2 88448 74404
0 26175 7 1 2 26173 26174
0 26176 5 1 1 26175
0 26177 7 1 2 26167 26176
0 26178 5 1 1 26177
0 26179 7 1 2 93095 26178
0 26180 5 1 1 26179
0 26181 7 2 2 76560 92776
0 26182 7 1 2 81817 76894
0 26183 7 1 2 80910 26182
0 26184 7 1 2 96480 26183
0 26185 5 1 1 26184
0 26186 7 1 2 77332 89968
0 26187 7 5 2 63162 93096
0 26188 7 1 2 91581 96482
0 26189 7 1 2 26186 26188
0 26190 5 1 1 26189
0 26191 7 1 2 26185 26190
0 26192 5 1 1 26191
0 26193 7 1 2 66963 26192
0 26194 5 1 1 26193
0 26195 7 2 2 66489 85918
0 26196 7 1 2 63337 96487
0 26197 7 1 2 78295 26196
0 26198 7 1 2 96253 26197
0 26199 5 1 1 26198
0 26200 7 1 2 69807 26199
0 26201 7 1 2 26194 26200
0 26202 7 1 2 26180 26201
0 26203 5 1 1 26202
0 26204 7 1 2 73015 26203
0 26205 7 1 2 26131 26204
0 26206 5 1 1 26205
0 26207 7 4 2 81989 96099
0 26208 5 2 1 96489
0 26209 7 7 2 82020 92777
0 26210 5 1 1 96495
0 26211 7 1 2 96493 26210
0 26212 5 4 1 26211
0 26213 7 1 2 96502 96428
0 26214 5 1 1 26213
0 26215 7 4 2 70351 82781
0 26216 7 2 2 71957 96506
0 26217 7 3 2 69366 96441
0 26218 7 1 2 76235 96512
0 26219 7 1 2 96510 26218
0 26220 5 1 1 26219
0 26221 7 7 2 83383 92778
0 26222 7 1 2 75149 86165
0 26223 5 1 1 26222
0 26224 7 1 2 79857 95195
0 26225 5 1 1 26224
0 26226 7 1 2 26223 26225
0 26227 5 1 1 26226
0 26228 7 1 2 96515 26227
0 26229 5 1 1 26228
0 26230 7 6 2 71333 76469
0 26231 7 5 2 88464 88915
0 26232 7 1 2 89957 96528
0 26233 7 1 2 96522 26232
0 26234 5 1 1 26233
0 26235 7 1 2 26229 26234
0 26236 5 1 1 26235
0 26237 7 1 2 65426 26236
0 26238 5 1 1 26237
0 26239 7 1 2 26220 26238
0 26240 7 1 2 26214 26239
0 26241 5 1 1 26240
0 26242 7 1 2 65756 26241
0 26243 5 1 1 26242
0 26244 7 2 2 75957 81279
0 26245 7 1 2 92123 96533
0 26246 5 1 1 26245
0 26247 7 1 2 85682 92066
0 26248 7 1 2 96529 26247
0 26249 5 1 1 26248
0 26250 7 1 2 26246 26249
0 26251 5 1 1 26250
0 26252 7 1 2 61865 26251
0 26253 5 1 1 26252
0 26254 7 1 2 81454 82529
0 26255 7 1 2 79936 26254
0 26256 7 1 2 91845 26255
0 26257 5 1 1 26256
0 26258 7 1 2 26253 26257
0 26259 5 1 1 26258
0 26260 7 1 2 67260 26259
0 26261 5 1 1 26260
0 26262 7 2 2 63338 82811
0 26263 7 6 2 68419 64349
0 26264 7 1 2 81990 96537
0 26265 7 1 2 96535 26264
0 26266 7 1 2 4769 26265
0 26267 5 1 1 26266
0 26268 7 1 2 26261 26267
0 26269 5 1 1 26268
0 26270 7 1 2 77317 26269
0 26271 5 1 1 26270
0 26272 7 1 2 26243 26271
0 26273 5 1 1 26272
0 26274 7 1 2 70079 26273
0 26275 5 1 1 26274
0 26276 7 1 2 81416 96100
0 26277 5 2 1 26276
0 26278 7 1 2 81280 93038
0 26279 5 1 1 26278
0 26280 7 1 2 96543 26279
0 26281 5 1 1 26280
0 26282 7 1 2 66730 26281
0 26283 5 1 1 26282
0 26284 7 7 2 88465 82901
0 26285 7 1 2 83056 96545
0 26286 5 1 1 26285
0 26287 7 1 2 26283 26286
0 26288 5 1 1 26287
0 26289 7 3 2 65757 93291
0 26290 5 1 1 96552
0 26291 7 1 2 62108 87438
0 26292 7 1 2 96553 26291
0 26293 7 1 2 26288 26292
0 26294 5 1 1 26293
0 26295 7 1 2 26275 26294
0 26296 5 1 1 26295
0 26297 7 1 2 67687 26296
0 26298 5 1 1 26297
0 26299 7 1 2 86250 94020
0 26300 5 1 1 26299
0 26301 7 1 2 95419 26300
0 26302 5 1 1 26301
0 26303 7 1 2 65758 26302
0 26304 5 1 1 26303
0 26305 7 1 2 79710 86464
0 26306 5 1 1 26305
0 26307 7 1 2 26304 26306
0 26308 5 1 1 26307
0 26309 7 4 2 82275 92114
0 26310 7 1 2 81281 96555
0 26311 5 1 1 26310
0 26312 7 1 2 96544 26311
0 26313 5 1 1 26312
0 26314 7 1 2 61866 26313
0 26315 5 1 1 26314
0 26316 7 1 2 87203 96496
0 26317 5 1 1 26316
0 26318 7 1 2 26315 26317
0 26319 5 1 1 26318
0 26320 7 1 2 26308 26319
0 26321 5 1 1 26320
0 26322 7 1 2 85136 95899
0 26323 7 1 2 86469 26322
0 26324 5 1 1 26323
0 26325 7 1 2 68660 84295
0 26326 5 1 1 26325
0 26327 7 1 2 78403 26326
0 26328 5 2 1 26327
0 26329 7 1 2 67261 96559
0 26330 5 1 1 26329
0 26331 7 2 2 75958 71529
0 26332 5 2 1 96561
0 26333 7 1 2 26330 96563
0 26334 5 4 1 26333
0 26335 7 1 2 74937 96516
0 26336 7 1 2 96565 26335
0 26337 5 1 1 26336
0 26338 7 1 2 26324 26337
0 26339 5 1 1 26338
0 26340 7 1 2 81991 26339
0 26341 5 1 1 26340
0 26342 7 2 2 68179 80911
0 26343 5 1 1 96569
0 26344 7 1 2 96566 96570
0 26345 5 1 1 26344
0 26346 7 1 2 83892 72447
0 26347 7 1 2 85137 26346
0 26348 5 1 1 26347
0 26349 7 1 2 26345 26348
0 26350 5 1 1 26349
0 26351 7 1 2 78840 96418
0 26352 7 1 2 26350 26351
0 26353 5 1 1 26352
0 26354 7 1 2 26341 26353
0 26355 5 1 1 26354
0 26356 7 1 2 67459 26355
0 26357 5 1 1 26356
0 26358 7 2 2 88510 92779
0 26359 7 1 2 81327 86499
0 26360 7 1 2 79176 26359
0 26361 7 1 2 96571 26360
0 26362 5 1 1 26361
0 26363 7 1 2 26357 26362
0 26364 5 1 1 26363
0 26365 7 1 2 66964 26364
0 26366 5 1 1 26365
0 26367 7 1 2 26321 26366
0 26368 5 1 1 26367
0 26369 7 1 2 65161 26368
0 26370 5 1 1 26369
0 26371 7 2 2 74156 93097
0 26372 7 2 2 88300 77409
0 26373 7 1 2 85126 96575
0 26374 7 1 2 96573 26373
0 26375 7 1 2 96554 26374
0 26376 5 1 1 26375
0 26377 7 1 2 26370 26376
0 26378 7 1 2 26298 26377
0 26379 5 1 1 26378
0 26380 7 1 2 76157 26379
0 26381 5 1 1 26380
0 26382 7 1 2 92920 93148
0 26383 5 3 1 26382
0 26384 7 2 2 66490 75705
0 26385 7 2 2 88998 96446
0 26386 7 1 2 96580 96582
0 26387 5 1 1 26386
0 26388 7 1 2 96577 26387
0 26389 5 1 1 26388
0 26390 7 1 2 88224 90847
0 26391 7 1 2 26389 26390
0 26392 5 1 1 26391
0 26393 7 1 2 88536 82295
0 26394 5 1 1 26393
0 26395 7 1 2 82326 77880
0 26396 5 1 1 26395
0 26397 7 1 2 26394 26396
0 26398 5 1 1 26397
0 26399 7 1 2 82623 96447
0 26400 7 1 2 82564 26399
0 26401 7 1 2 26398 26400
0 26402 5 1 1 26401
0 26403 7 1 2 26392 26402
0 26404 5 1 1 26403
0 26405 7 1 2 64734 26404
0 26406 5 1 1 26405
0 26407 7 10 2 90957 91516
0 26408 5 2 1 96584
0 26409 7 2 2 80937 96237
0 26410 5 1 1 96596
0 26411 7 1 2 96594 26410
0 26412 5 2 1 26411
0 26413 7 1 2 89459 89250
0 26414 7 1 2 88537 26413
0 26415 7 1 2 96598 26414
0 26416 5 1 1 26415
0 26417 7 1 2 26406 26416
0 26418 5 1 1 26417
0 26419 7 1 2 65759 26418
0 26420 5 1 1 26419
0 26421 7 1 2 88873 89382
0 26422 7 1 2 92033 26421
0 26423 5 1 1 26422
0 26424 7 1 2 73917 85242
0 26425 7 1 2 82028 26424
0 26426 5 1 1 26425
0 26427 7 1 2 26423 26426
0 26428 5 1 1 26427
0 26429 7 1 2 68180 26428
0 26430 5 1 1 26429
0 26431 7 2 2 62414 80649
0 26432 7 1 2 90092 92034
0 26433 7 1 2 96600 26432
0 26434 5 1 1 26433
0 26435 7 1 2 26430 26434
0 26436 5 1 1 26435
0 26437 7 1 2 82276 26436
0 26438 5 1 1 26437
0 26439 7 1 2 80034 92884
0 26440 7 2 2 90100 26439
0 26441 7 1 2 67262 79327
0 26442 7 1 2 96602 26441
0 26443 5 1 1 26442
0 26444 7 1 2 26438 26443
0 26445 5 1 1 26444
0 26446 7 1 2 69200 26445
0 26447 5 1 1 26446
0 26448 7 3 2 69367 87937
0 26449 7 1 2 81992 89261
0 26450 7 1 2 94549 26449
0 26451 7 1 2 96604 26450
0 26452 5 1 1 26451
0 26453 7 1 2 26447 26452
0 26454 5 1 1 26453
0 26455 7 1 2 78823 26454
0 26456 5 1 1 26455
0 26457 7 1 2 26420 26456
0 26458 5 1 1 26457
0 26459 7 1 2 65427 26458
0 26460 5 1 1 26459
0 26461 7 1 2 79889 89697
0 26462 5 1 1 26461
0 26463 7 1 2 86251 95742
0 26464 5 1 1 26463
0 26465 7 1 2 26462 26464
0 26466 5 1 1 26465
0 26467 7 1 2 65428 26466
0 26468 5 1 1 26467
0 26469 7 2 2 70352 76446
0 26470 7 1 2 81305 96607
0 26471 5 1 1 26470
0 26472 7 1 2 26468 26471
0 26473 5 1 1 26472
0 26474 7 1 2 62109 26473
0 26475 5 1 1 26474
0 26476 7 1 2 89532 22050
0 26477 5 1 1 26476
0 26478 7 1 2 81306 72849
0 26479 7 1 2 26477 26478
0 26480 5 1 1 26479
0 26481 7 1 2 26475 26480
0 26482 5 1 1 26481
0 26483 7 1 2 96585 26482
0 26484 5 1 1 26483
0 26485 7 1 2 75907 96426
0 26486 5 1 1 26485
0 26487 7 1 2 70080 26486
0 26488 5 1 1 26487
0 26489 7 1 2 87866 80777
0 26490 5 1 1 26489
0 26491 7 1 2 26488 26490
0 26492 5 1 1 26491
0 26493 7 1 2 75875 95933
0 26494 7 1 2 26492 26493
0 26495 5 1 1 26494
0 26496 7 1 2 26484 26495
0 26497 5 1 1 26496
0 26498 7 1 2 65760 26497
0 26499 5 1 1 26498
0 26500 7 1 2 73066 88608
0 26501 7 2 2 90237 93098
0 26502 7 1 2 94151 96609
0 26503 7 1 2 26500 26502
0 26504 5 1 1 26503
0 26505 7 1 2 26499 26504
0 26506 5 1 1 26505
0 26507 7 1 2 79177 26506
0 26508 5 1 1 26507
0 26509 7 1 2 82021 96419
0 26510 5 1 1 26509
0 26511 7 1 2 96494 26510
0 26512 5 2 1 26511
0 26513 7 1 2 77245 96611
0 26514 5 1 1 26513
0 26515 7 1 2 84220 96073
0 26516 5 1 1 26515
0 26517 7 1 2 26514 26516
0 26518 5 1 1 26517
0 26519 7 1 2 80618 82458
0 26520 7 1 2 81562 26519
0 26521 7 1 2 26518 26520
0 26522 5 1 1 26521
0 26523 7 1 2 26508 26522
0 26524 7 1 2 26460 26523
0 26525 7 1 2 26381 26524
0 26526 7 1 2 26206 26525
0 26527 7 1 2 26076 26526
0 26528 5 1 1 26527
0 26529 7 1 2 72160 26528
0 26530 5 1 1 26529
0 26531 7 1 2 84870 95905
0 26532 5 1 1 26531
0 26533 7 2 2 94128 96175
0 26534 5 1 1 96613
0 26535 7 1 2 65429 96614
0 26536 5 1 1 26535
0 26537 7 1 2 26532 26536
0 26538 5 1 1 26537
0 26539 7 1 2 68845 26538
0 26540 5 1 1 26539
0 26541 7 8 2 64522 96193
0 26542 7 1 2 88118 96615
0 26543 7 1 2 93447 26542
0 26544 7 1 2 95712 26543
0 26545 5 1 1 26544
0 26546 7 1 2 26540 26545
0 26547 5 1 1 26546
0 26548 7 1 2 61586 26547
0 26549 5 1 1 26548
0 26550 7 2 2 68989 73121
0 26551 5 2 1 96623
0 26552 7 1 2 72491 12137
0 26553 5 1 1 26552
0 26554 7 1 2 67688 26553
0 26555 5 1 1 26554
0 26556 7 1 2 96625 26555
0 26557 5 1 1 26556
0 26558 7 1 2 65990 26557
0 26559 5 1 1 26558
0 26560 7 1 2 72448 79320
0 26561 5 1 1 26560
0 26562 7 1 2 26559 26561
0 26563 5 1 1 26562
0 26564 7 4 2 69201 79365
0 26565 7 1 2 80980 96627
0 26566 7 1 2 26563 26565
0 26567 5 1 1 26566
0 26568 7 1 2 26549 26567
0 26569 5 1 1 26568
0 26570 7 1 2 71057 26569
0 26571 5 1 1 26570
0 26572 7 1 2 75530 96624
0 26573 5 1 1 26572
0 26574 7 1 2 72345 95365
0 26575 5 1 1 26574
0 26576 7 1 2 26573 26575
0 26577 5 1 1 26576
0 26578 7 1 2 81923 26577
0 26579 5 1 1 26578
0 26580 7 2 2 73067 88250
0 26581 7 1 2 93383 96631
0 26582 5 1 1 26581
0 26583 7 1 2 26579 26582
0 26584 5 1 1 26583
0 26585 7 2 2 69202 82239
0 26586 7 1 2 81653 96633
0 26587 7 1 2 26584 26586
0 26588 5 1 1 26587
0 26589 7 1 2 26571 26588
0 26590 5 1 1 26589
0 26591 7 1 2 68181 26590
0 26592 5 1 1 26591
0 26593 7 2 2 69570 84871
0 26594 7 1 2 78841 96635
0 26595 5 1 1 26594
0 26596 7 2 2 86698 83348
0 26597 5 2 1 96637
0 26598 7 1 2 26595 96639
0 26599 5 1 1 26598
0 26600 7 2 2 69368 87855
0 26601 7 1 2 77246 87204
0 26602 7 1 2 96641 26601
0 26603 7 1 2 26599 26602
0 26604 5 1 1 26603
0 26605 7 1 2 26592 26604
0 26606 5 1 1 26605
0 26607 7 1 2 74808 26606
0 26608 5 1 1 26607
0 26609 7 1 2 63339 96638
0 26610 5 1 1 26609
0 26611 7 1 2 84484 96636
0 26612 5 1 1 26611
0 26613 7 1 2 26610 26612
0 26614 5 1 1 26613
0 26615 7 1 2 67689 26614
0 26616 5 1 1 26615
0 26617 7 1 2 79809 91187
0 26618 7 1 2 89680 26617
0 26619 5 1 1 26618
0 26620 7 1 2 26616 26619
0 26621 5 1 1 26620
0 26622 7 1 2 72375 96586
0 26623 7 1 2 26621 26622
0 26624 5 1 1 26623
0 26625 7 1 2 26608 26624
0 26626 5 1 1 26625
0 26627 7 1 2 84946 26626
0 26628 5 1 1 26627
0 26629 7 1 2 90406 86699
0 26630 5 1 1 26629
0 26631 7 1 2 81282 87591
0 26632 7 1 2 80058 26631
0 26633 5 1 1 26632
0 26634 7 1 2 26630 26633
0 26635 5 1 1 26634
0 26636 7 1 2 63163 26635
0 26637 5 1 1 26636
0 26638 7 1 2 81417 78769
0 26639 7 1 2 80242 95041
0 26640 7 1 2 26638 26639
0 26641 5 1 1 26640
0 26642 7 1 2 26637 26641
0 26643 5 1 1 26642
0 26644 7 1 2 61587 26643
0 26645 5 1 1 26644
0 26646 7 1 2 80350 91297
0 26647 7 1 2 93416 26646
0 26648 5 1 1 26647
0 26649 7 1 2 26645 26648
0 26650 5 1 1 26649
0 26651 7 1 2 83558 95302
0 26652 7 1 2 91416 26651
0 26653 7 1 2 26650 26652
0 26654 5 1 1 26653
0 26655 7 1 2 26628 26654
0 26656 5 1 1 26655
0 26657 7 1 2 67460 26656
0 26658 5 1 1 26657
0 26659 7 3 2 77201 76001
0 26660 5 1 1 96643
0 26661 7 1 2 74078 75896
0 26662 5 1 1 26661
0 26663 7 1 2 62843 87996
0 26664 5 1 1 26663
0 26665 7 1 2 26662 26664
0 26666 5 6 1 26665
0 26667 7 1 2 96644 96646
0 26668 5 1 1 26667
0 26669 7 2 2 77498 71058
0 26670 5 1 1 96652
0 26671 7 1 2 71530 96653
0 26672 5 1 1 26671
0 26673 7 1 2 77539 95784
0 26674 5 1 1 26673
0 26675 7 1 2 71059 26674
0 26676 5 1 1 26675
0 26677 7 1 2 72289 96013
0 26678 5 1 1 26677
0 26679 7 1 2 26676 26678
0 26680 5 1 1 26679
0 26681 7 1 2 67461 26680
0 26682 5 1 1 26681
0 26683 7 1 2 26672 26682
0 26684 5 1 1 26683
0 26685 7 1 2 76158 26684
0 26686 5 1 1 26685
0 26687 7 1 2 26668 26686
0 26688 5 1 1 26687
0 26689 7 1 2 64735 26688
0 26690 5 1 1 26689
0 26691 7 3 2 69571 74182
0 26692 7 2 2 75350 94235
0 26693 7 1 2 93398 96657
0 26694 7 1 2 96654 26693
0 26695 5 1 1 26694
0 26696 7 1 2 26690 26695
0 26697 5 1 1 26696
0 26698 7 1 2 92780 26697
0 26699 5 1 1 26698
0 26700 7 1 2 85356 95869
0 26701 5 2 1 26700
0 26702 7 1 2 84382 85476
0 26703 5 1 1 26702
0 26704 7 1 2 96659 26703
0 26705 5 1 1 26704
0 26706 7 1 2 71438 26705
0 26707 5 1 1 26706
0 26708 7 3 2 64130 73459
0 26709 5 2 1 96661
0 26710 7 2 2 70921 96662
0 26711 5 3 1 96666
0 26712 7 1 2 72303 96668
0 26713 5 1 1 26712
0 26714 7 1 2 67690 26713
0 26715 5 1 1 26714
0 26716 7 1 2 70704 86735
0 26717 5 1 1 26716
0 26718 7 1 2 26715 26717
0 26719 5 1 1 26718
0 26720 7 1 2 71060 26719
0 26721 5 1 1 26720
0 26722 7 1 2 26707 26721
0 26723 5 1 1 26722
0 26724 7 4 2 89262 96139
0 26725 7 1 2 26723 96671
0 26726 5 1 1 26725
0 26727 7 1 2 26699 26726
0 26728 5 1 1 26727
0 26729 7 1 2 76942 26728
0 26730 5 1 1 26729
0 26731 7 1 2 90517 93075
0 26732 5 1 1 26731
0 26733 7 1 2 26732 96578
0 26734 5 1 1 26733
0 26735 7 1 2 89518 26734
0 26736 5 1 1 26735
0 26737 7 2 2 88770 76590
0 26738 7 1 2 93099 96675
0 26739 5 1 1 26738
0 26740 7 8 2 68990 69203
0 26741 7 1 2 71470 96677
0 26742 7 1 2 95253 26741
0 26743 5 1 1 26742
0 26744 7 1 2 26739 26743
0 26745 5 1 1 26744
0 26746 7 1 2 65991 26745
0 26747 5 1 1 26746
0 26748 7 1 2 26736 26747
0 26749 5 1 1 26748
0 26750 7 1 2 68846 26749
0 26751 5 1 1 26750
0 26752 7 4 2 68991 81210
0 26753 5 2 1 96685
0 26754 7 2 2 93100 96686
0 26755 7 1 2 83001 96691
0 26756 5 1 1 26755
0 26757 7 1 2 26751 26756
0 26758 5 1 1 26757
0 26759 7 1 2 67462 26758
0 26760 5 1 1 26759
0 26761 7 4 2 61588 88771
0 26762 7 1 2 71017 96693
0 26763 7 1 2 96692 26762
0 26764 5 1 1 26763
0 26765 7 1 2 26760 26764
0 26766 5 1 1 26765
0 26767 7 1 2 78194 90767
0 26768 7 1 2 26766 26767
0 26769 5 1 1 26768
0 26770 7 1 2 68182 26769
0 26771 7 1 2 26730 26770
0 26772 5 1 1 26771
0 26773 7 1 2 72274 93437
0 26774 5 1 1 26773
0 26775 7 1 2 95788 26774
0 26776 5 1 1 26775
0 26777 7 1 2 68016 26776
0 26778 5 1 1 26777
0 26779 7 1 2 95778 95782
0 26780 5 1 1 26779
0 26781 7 1 2 26778 26780
0 26782 5 1 1 26781
0 26783 7 3 2 82076 96094
0 26784 7 1 2 26782 96697
0 26785 5 1 1 26784
0 26786 7 1 2 77841 95974
0 26787 5 1 1 26786
0 26788 7 1 2 76159 96490
0 26789 7 1 2 26787 26788
0 26790 5 1 1 26789
0 26791 7 1 2 26785 26790
0 26792 5 1 1 26791
0 26793 7 1 2 76943 26792
0 26794 5 1 1 26793
0 26795 7 1 2 84183 86478
0 26796 7 3 2 68847 88029
0 26797 7 1 2 92893 96700
0 26798 7 1 2 26795 26797
0 26799 5 1 1 26798
0 26800 7 1 2 26794 26799
0 26801 5 1 1 26800
0 26802 7 1 2 67463 26801
0 26803 5 1 1 26802
0 26804 7 1 2 2253 94541
0 26805 5 1 1 26804
0 26806 7 1 2 68848 26805
0 26807 5 1 1 26806
0 26808 7 2 2 70353 86805
0 26809 7 1 2 65162 96703
0 26810 5 1 1 26809
0 26811 7 1 2 26807 26810
0 26812 5 1 1 26811
0 26813 7 1 2 67464 26812
0 26814 5 1 1 26813
0 26815 7 2 2 76944 86700
0 26816 5 2 1 96705
0 26817 7 1 2 72552 86479
0 26818 5 4 1 26817
0 26819 7 1 2 94542 96709
0 26820 5 2 1 26819
0 26821 7 1 2 73460 96713
0 26822 5 1 1 26821
0 26823 7 1 2 96707 26822
0 26824 5 1 1 26823
0 26825 7 1 2 67691 26824
0 26826 5 1 1 26825
0 26827 7 1 2 73863 82459
0 26828 5 1 1 26827
0 26829 7 1 2 26826 26828
0 26830 7 1 2 26814 26829
0 26831 5 1 1 26830
0 26832 7 1 2 96587 26831
0 26833 5 1 1 26832
0 26834 7 1 2 84383 79041
0 26835 5 2 1 26834
0 26836 7 1 2 72553 79034
0 26837 5 1 1 26836
0 26838 7 1 2 96715 26837
0 26839 5 1 1 26838
0 26840 7 1 2 92781 95396
0 26841 7 1 2 26839 26840
0 26842 5 1 1 26841
0 26843 7 1 2 26833 26842
0 26844 5 1 1 26843
0 26845 7 1 2 79178 26844
0 26846 5 1 1 26845
0 26847 7 1 2 79045 12113
0 26848 5 2 1 26847
0 26849 7 1 2 76090 96503
0 26850 5 1 1 26849
0 26851 7 1 2 84475 96546
0 26852 5 2 1 26851
0 26853 7 1 2 26850 96719
0 26854 5 1 1 26853
0 26855 7 1 2 96717 26854
0 26856 5 1 1 26855
0 26857 7 4 2 78475 79534
0 26858 7 3 2 69204 76707
0 26859 7 1 2 81654 88638
0 26860 7 1 2 96725 26859
0 26861 7 1 2 96721 26860
0 26862 5 1 1 26861
0 26863 7 1 2 26856 26862
0 26864 5 1 1 26863
0 26865 7 1 2 67465 26864
0 26866 5 1 1 26865
0 26867 7 1 2 83759 93101
0 26868 7 1 2 93468 26867
0 26869 7 1 2 83865 26868
0 26870 5 1 1 26869
0 26871 7 1 2 26866 26870
0 26872 5 1 1 26871
0 26873 7 1 2 89519 26872
0 26874 5 1 1 26873
0 26875 7 4 2 68849 92782
0 26876 7 2 2 82022 96728
0 26877 7 1 2 74120 96732
0 26878 5 1 1 26877
0 26879 7 1 2 64131 84568
0 26880 7 1 2 96491 26879
0 26881 5 1 1 26880
0 26882 7 1 2 26878 26881
0 26883 5 1 1 26882
0 26884 7 1 2 79213 26883
0 26885 5 1 1 26884
0 26886 7 1 2 83749 87141
0 26887 7 1 2 96497 26886
0 26888 5 1 1 26887
0 26889 7 1 2 26885 26888
0 26890 5 1 1 26889
0 26891 7 1 2 84851 26890
0 26892 5 1 1 26891
0 26893 7 1 2 63340 26892
0 26894 7 1 2 26874 26893
0 26895 7 1 2 26846 26894
0 26896 7 1 2 26803 26895
0 26897 5 1 1 26896
0 26898 7 1 2 73016 26897
0 26899 7 1 2 26772 26898
0 26900 5 1 1 26899
0 26901 7 1 2 88206 96180
0 26902 5 1 1 26901
0 26903 7 2 2 74121 93039
0 26904 7 1 2 68017 87057
0 26905 7 1 2 96734 26904
0 26906 5 1 1 26905
0 26907 7 1 2 26902 26906
0 26908 5 1 1 26907
0 26909 7 9 2 61589 70922
0 26910 7 1 2 86085 96736
0 26911 7 1 2 79986 26910
0 26912 7 1 2 26908 26911
0 26913 5 1 1 26912
0 26914 7 1 2 26900 26913
0 26915 7 1 2 26658 26914
0 26916 5 1 1 26915
0 26917 7 1 2 75801 26916
0 26918 5 1 1 26917
0 26919 7 1 2 84366 92024
0 26920 7 2 2 75382 26919
0 26921 5 1 1 96745
0 26922 7 1 2 87893 91319
0 26923 7 1 2 96378 26922
0 26924 5 1 1 26923
0 26925 7 1 2 26921 26924
0 26926 5 1 1 26925
0 26927 7 1 2 66731 26926
0 26928 5 1 1 26927
0 26929 7 1 2 77202 88154
0 26930 7 1 2 96687 26929
0 26931 5 1 1 26930
0 26932 7 1 2 26928 26931
0 26933 5 1 1 26932
0 26934 7 1 2 63341 26933
0 26935 5 1 1 26934
0 26936 7 1 2 83057 96746
0 26937 5 1 1 26936
0 26938 7 1 2 26935 26937
0 26939 5 1 1 26938
0 26940 7 1 2 63164 26939
0 26941 5 1 1 26940
0 26942 7 1 2 88589 75351
0 26943 7 1 2 84367 26942
0 26944 7 1 2 92619 26943
0 26945 5 1 1 26944
0 26946 7 1 2 26941 26945
0 26947 5 1 1 26946
0 26948 7 1 2 81345 26947
0 26949 5 1 1 26948
0 26950 7 1 2 81585 84507
0 26951 5 1 1 26950
0 26952 7 1 2 72554 81307
0 26953 7 1 2 78139 26952
0 26954 5 1 1 26953
0 26955 7 1 2 26951 26954
0 26956 5 1 1 26955
0 26957 7 1 2 62415 26956
0 26958 5 1 1 26957
0 26959 7 1 2 84502 87575
0 26960 7 1 2 93255 26959
0 26961 5 1 1 26960
0 26962 7 1 2 26958 26961
0 26963 5 1 1 26962
0 26964 7 1 2 95021 26963
0 26965 5 1 1 26964
0 26966 7 1 2 26949 26965
0 26967 5 1 1 26966
0 26968 7 1 2 70354 26967
0 26969 5 1 1 26968
0 26970 7 2 2 69808 90193
0 26971 7 1 2 74122 96747
0 26972 5 1 1 26971
0 26973 7 1 2 63165 84485
0 26974 5 1 1 26973
0 26975 7 1 2 26972 26974
0 26976 5 1 1 26975
0 26977 7 1 2 70923 26976
0 26978 5 1 1 26977
0 26979 7 1 2 72789 96748
0 26980 5 1 1 26979
0 26981 7 1 2 26978 26980
0 26982 5 1 1 26981
0 26983 7 1 2 61590 26982
0 26984 5 1 1 26983
0 26985 7 1 2 88874 81418
0 26986 7 1 2 89498 26985
0 26987 5 1 1 26986
0 26988 7 1 2 26984 26987
0 26989 5 1 1 26988
0 26990 7 1 2 69572 26989
0 26991 5 1 1 26990
0 26992 7 1 2 85989 92873
0 26993 5 1 1 26992
0 26994 7 1 2 26991 26993
0 26995 5 1 1 26994
0 26996 7 1 2 84947 26995
0 26997 5 1 1 26996
0 26998 7 1 2 82055 91217
0 26999 7 1 2 91782 91918
0 27000 7 1 2 26998 26999
0 27001 5 1 1 27000
0 27002 7 1 2 26997 27001
0 27003 5 1 1 27002
0 27004 7 1 2 74322 27003
0 27005 5 1 1 27004
0 27006 7 1 2 26969 27005
0 27007 5 1 1 27006
0 27008 7 1 2 93102 27007
0 27009 5 1 1 27008
0 27010 7 1 2 89475 95827
0 27011 7 2 2 90073 27010
0 27012 7 1 2 83058 96749
0 27013 5 1 1 27012
0 27014 7 1 2 89399 83787
0 27015 5 1 1 27014
0 27016 7 1 2 88971 94129
0 27017 5 1 1 27016
0 27018 7 1 2 90060 27017
0 27019 5 1 1 27018
0 27020 7 1 2 81261 27019
0 27021 5 1 1 27020
0 27022 7 1 2 27015 27021
0 27023 5 1 1 27022
0 27024 7 1 2 66732 27023
0 27025 5 1 1 27024
0 27026 7 1 2 27013 27025
0 27027 5 1 1 27026
0 27028 7 2 2 70081 92783
0 27029 7 1 2 71958 74323
0 27030 7 1 2 96751 27029
0 27031 7 1 2 27027 27030
0 27032 5 1 1 27031
0 27033 7 1 2 27009 27032
0 27034 5 1 1 27033
0 27035 7 1 2 65761 27034
0 27036 5 1 1 27035
0 27037 7 1 2 64943 71959
0 27038 7 1 2 81800 27037
0 27039 5 1 1 27038
0 27040 7 1 2 64132 79179
0 27041 7 1 2 74718 27040
0 27042 5 1 1 27041
0 27043 7 1 2 27039 27042
0 27044 5 1 1 27043
0 27045 7 1 2 68183 27044
0 27046 5 1 1 27045
0 27047 7 4 2 69809 80149
0 27048 7 1 2 61867 96753
0 27049 5 1 1 27048
0 27050 7 1 2 79111 27049
0 27051 5 2 1 27050
0 27052 7 1 2 83414 76475
0 27053 7 1 2 96757 27052
0 27054 5 1 1 27053
0 27055 7 1 2 27046 27054
0 27056 5 1 1 27055
0 27057 7 1 2 67692 27056
0 27058 5 1 1 27057
0 27059 7 2 2 74324 79079
0 27060 5 1 1 96759
0 27061 7 1 2 68992 96760
0 27062 7 1 2 89393 27061
0 27063 5 1 1 27062
0 27064 7 1 2 27058 27063
0 27065 5 1 1 27064
0 27066 7 1 2 70924 27065
0 27067 5 1 1 27066
0 27068 7 1 2 61868 81283
0 27069 5 2 1 27068
0 27070 7 1 2 66733 95854
0 27071 5 1 1 27070
0 27072 7 1 2 96761 27071
0 27073 5 1 1 27072
0 27074 7 1 2 88566 89970
0 27075 7 1 2 27073 27074
0 27076 5 1 1 27075
0 27077 7 1 2 27067 27076
0 27078 5 1 1 27077
0 27079 7 1 2 96140 27078
0 27080 5 1 1 27079
0 27081 7 4 2 70705 92784
0 27082 7 1 2 78179 83275
0 27083 7 1 2 96763 27082
0 27084 7 1 2 89396 27083
0 27085 5 1 1 27084
0 27086 7 1 2 27080 27085
0 27087 5 1 1 27086
0 27088 7 1 2 61591 27087
0 27089 5 1 1 27088
0 27090 7 2 2 75055 87018
0 27091 5 1 1 96767
0 27092 7 1 2 89971 96768
0 27093 5 1 1 27092
0 27094 7 1 2 74435 77484
0 27095 7 1 2 74416 27094
0 27096 5 1 1 27095
0 27097 7 1 2 27093 27096
0 27098 5 1 1 27097
0 27099 7 1 2 96530 27098
0 27100 5 1 1 27099
0 27101 7 5 2 68420 89912
0 27102 7 4 2 68993 92785
0 27103 7 2 2 96769 96774
0 27104 7 3 2 88251 74970
0 27105 7 1 2 71960 96780
0 27106 7 1 2 96778 27105
0 27107 5 1 1 27106
0 27108 7 1 2 27100 27107
0 27109 5 1 1 27108
0 27110 7 1 2 61869 27109
0 27111 5 1 1 27110
0 27112 7 2 2 64944 87091
0 27113 5 1 1 96783
0 27114 7 1 2 90061 27113
0 27115 5 1 1 27114
0 27116 7 3 2 88252 92786
0 27117 7 1 2 71961 82624
0 27118 7 1 2 73729 27117
0 27119 7 1 2 96785 27118
0 27120 7 1 2 27115 27119
0 27121 5 1 1 27120
0 27122 7 1 2 27111 27121
0 27123 5 1 1 27122
0 27124 7 1 2 76160 27123
0 27125 5 1 1 27124
0 27126 7 1 2 80295 83226
0 27127 5 1 1 27126
0 27128 7 2 2 64133 74971
0 27129 5 1 1 96788
0 27130 7 1 2 90062 27129
0 27131 5 1 1 27130
0 27132 7 1 2 67693 4859
0 27133 7 1 2 27131 27132
0 27134 5 1 1 27133
0 27135 7 1 2 27127 27134
0 27136 5 1 1 27135
0 27137 7 1 2 66734 27136
0 27138 5 1 1 27137
0 27139 7 1 2 81499 96789
0 27140 5 1 1 27139
0 27141 7 1 2 27138 27140
0 27142 5 1 1 27141
0 27143 7 1 2 85963 27142
0 27144 5 1 1 27143
0 27145 7 2 2 75211 95836
0 27146 7 1 2 82161 96790
0 27147 5 1 1 27146
0 27148 7 1 2 27144 27147
0 27149 5 1 1 27148
0 27150 7 5 2 83458 80949
0 27151 7 1 2 96628 96792
0 27152 7 1 2 27149 27151
0 27153 5 1 1 27152
0 27154 7 1 2 27125 27153
0 27155 7 1 2 27089 27154
0 27156 5 1 1 27155
0 27157 7 1 2 70082 27156
0 27158 5 1 1 27157
0 27159 7 1 2 27036 27158
0 27160 5 1 1 27159
0 27161 7 1 2 73461 27160
0 27162 5 1 1 27161
0 27163 7 1 2 72161 74634
0 27164 7 2 2 96101 27163
0 27165 7 1 2 82376 96797
0 27166 5 1 1 27165
0 27167 7 1 2 66735 78214
0 27168 7 1 2 96517 27167
0 27169 5 1 1 27168
0 27170 7 1 2 27166 27169
0 27171 5 1 1 27170
0 27172 7 1 2 63166 27171
0 27173 5 1 1 27172
0 27174 7 1 2 91254 84049
0 27175 7 1 2 96775 27174
0 27176 5 1 1 27175
0 27177 7 1 2 27173 27176
0 27178 5 1 1 27177
0 27179 7 1 2 66491 27178
0 27180 5 1 1 27179
0 27181 7 1 2 78221 95975
0 27182 5 1 1 27181
0 27183 7 1 2 90044 93040
0 27184 7 1 2 27182 27183
0 27185 5 1 1 27184
0 27186 7 1 2 27180 27185
0 27187 5 1 1 27186
0 27188 7 1 2 65762 27187
0 27189 5 1 1 27188
0 27190 7 1 2 61592 96798
0 27191 5 1 1 27190
0 27192 7 1 2 88624 91846
0 27193 7 1 2 89499 27192
0 27194 5 1 1 27193
0 27195 7 1 2 27191 27194
0 27196 5 1 1 27195
0 27197 7 1 2 65763 27196
0 27198 5 1 1 27197
0 27199 7 2 2 89363 96786
0 27200 5 1 1 96799
0 27201 7 1 2 83760 96800
0 27202 5 1 1 27201
0 27203 7 1 2 27198 27202
0 27204 5 1 1 27203
0 27205 7 1 2 90194 27204
0 27206 5 1 1 27205
0 27207 7 4 2 72275 92787
0 27208 7 1 2 94236 96117
0 27209 7 1 2 89084 27208
0 27210 7 1 2 96801 27209
0 27211 5 1 1 27210
0 27212 7 1 2 27206 27211
0 27213 7 1 2 27189 27212
0 27214 5 1 1 27213
0 27215 7 1 2 64945 27214
0 27216 5 1 1 27215
0 27217 7 2 2 69573 83692
0 27218 7 1 2 93103 96805
0 27219 5 1 1 27218
0 27220 7 1 2 90518 96518
0 27221 5 1 1 27220
0 27222 7 1 2 27219 27221
0 27223 5 1 1 27222
0 27224 7 1 2 65764 27223
0 27225 5 1 1 27224
0 27226 7 2 2 85643 84467
0 27227 7 1 2 92124 96807
0 27228 5 1 1 27227
0 27229 7 1 2 27225 27228
0 27230 5 1 1 27229
0 27231 7 1 2 72555 27230
0 27232 5 1 1 27231
0 27233 7 2 2 71531 93041
0 27234 5 1 1 96809
0 27235 7 1 2 96808 96810
0 27236 5 1 1 27235
0 27237 7 1 2 27232 27236
0 27238 5 1 1 27237
0 27239 7 1 2 75252 27238
0 27240 5 1 1 27239
0 27241 7 1 2 27216 27240
0 27242 5 1 1 27241
0 27243 7 1 2 75773 27242
0 27244 5 1 1 27243
0 27245 7 1 2 89500 89623
0 27246 5 1 1 27245
0 27247 7 1 2 91932 27246
0 27248 5 1 1 27247
0 27249 7 1 2 71236 27248
0 27250 5 1 1 27249
0 27251 7 2 2 69810 73649
0 27252 7 1 2 81735 96811
0 27253 5 1 1 27252
0 27254 7 1 2 91933 27253
0 27255 5 1 1 27254
0 27256 7 1 2 68994 27255
0 27257 5 1 1 27256
0 27258 7 1 2 74635 73578
0 27259 7 1 2 90503 27258
0 27260 5 1 1 27259
0 27261 7 1 2 27257 27260
0 27262 5 1 1 27261
0 27263 7 1 2 65765 27262
0 27264 5 1 1 27263
0 27265 7 1 2 27250 27264
0 27266 5 1 1 27265
0 27267 7 1 2 69574 27266
0 27268 5 1 1 27267
0 27269 7 1 2 82664 96754
0 27270 7 1 2 86850 27269
0 27271 5 1 1 27270
0 27272 7 1 2 27268 27271
0 27273 5 1 1 27272
0 27274 7 1 2 61593 27273
0 27275 5 1 1 27274
0 27276 7 1 2 73663 95979
0 27277 5 2 1 27276
0 27278 7 1 2 82782 91762
0 27279 7 1 2 96813 27278
0 27280 5 1 1 27279
0 27281 7 1 2 27275 27280
0 27282 5 1 1 27281
0 27283 7 1 2 93104 27282
0 27284 5 1 1 27283
0 27285 7 3 2 64523 93016
0 27286 7 1 2 92885 96815
0 27287 7 1 2 96750 27286
0 27288 5 1 1 27287
0 27289 7 1 2 61870 27288
0 27290 7 1 2 27284 27289
0 27291 5 1 1 27290
0 27292 7 1 2 73659 78952
0 27293 5 1 1 27292
0 27294 7 2 2 89063 91478
0 27295 5 1 1 96818
0 27296 7 1 2 91176 96819
0 27297 5 1 1 27296
0 27298 7 1 2 71237 72628
0 27299 7 1 2 27297 27298
0 27300 5 1 1 27299
0 27301 7 1 2 27293 27300
0 27302 5 1 1 27301
0 27303 7 1 2 96133 27302
0 27304 5 1 1 27303
0 27305 7 1 2 74636 78312
0 27306 5 1 1 27305
0 27307 7 1 2 84874 27306
0 27308 5 1 1 27307
0 27309 7 1 2 96181 27308
0 27310 5 1 1 27309
0 27311 7 3 2 69369 80243
0 27312 7 2 2 90958 96820
0 27313 5 1 1 96823
0 27314 7 1 2 26534 27313
0 27315 5 1 1 27314
0 27316 7 1 2 71238 27315
0 27317 5 1 1 27316
0 27318 7 1 2 78968 93713
0 27319 7 1 2 96776 27318
0 27320 5 1 1 27319
0 27321 7 1 2 27317 27320
0 27322 7 1 2 27310 27321
0 27323 5 1 1 27322
0 27324 7 1 2 61594 27323
0 27325 5 1 1 27324
0 27326 7 1 2 27304 27325
0 27327 5 1 1 27326
0 27328 7 1 2 88972 27327
0 27329 5 1 1 27328
0 27330 7 1 2 71168 92530
0 27331 5 1 1 27330
0 27332 7 1 2 25020 27331
0 27333 5 1 1 27332
0 27334 7 1 2 70706 27333
0 27335 5 1 1 27334
0 27336 7 1 2 91219 93365
0 27337 5 1 1 27336
0 27338 7 1 2 27335 27337
0 27339 5 1 1 27338
0 27340 7 1 2 71239 27339
0 27341 5 1 1 27340
0 27342 7 4 2 67694 76323
0 27343 5 1 1 96825
0 27344 7 1 2 88232 90524
0 27345 7 1 2 96826 27344
0 27346 5 1 1 27345
0 27347 7 1 2 27341 27346
0 27348 5 1 1 27347
0 27349 7 1 2 92788 27348
0 27350 5 1 1 27349
0 27351 7 1 2 96672 96814
0 27352 5 1 1 27351
0 27353 7 1 2 27350 27352
0 27354 5 1 1 27353
0 27355 7 1 2 88948 27354
0 27356 5 1 1 27355
0 27357 7 1 2 66736 27356
0 27358 7 1 2 27329 27357
0 27359 5 1 1 27358
0 27360 7 1 2 74325 27359
0 27361 7 1 2 27291 27360
0 27362 5 1 1 27361
0 27363 7 1 2 27244 27362
0 27364 5 1 1 27363
0 27365 7 1 2 70083 27364
0 27366 5 1 1 27365
0 27367 7 1 2 79128 90045
0 27368 5 1 1 27367
0 27369 7 1 2 66737 87524
0 27370 5 1 1 27369
0 27371 7 1 2 79129 85327
0 27372 5 1 1 27371
0 27373 7 1 2 27370 27372
0 27374 5 1 1 27373
0 27375 7 1 2 66492 27374
0 27376 5 1 1 27375
0 27377 7 1 2 27368 27376
0 27378 5 1 1 27377
0 27379 7 1 2 94097 27378
0 27380 5 1 1 27379
0 27381 7 1 2 63342 76350
0 27382 7 1 2 78998 27381
0 27383 5 1 1 27382
0 27384 7 1 2 27380 27383
0 27385 5 1 1 27384
0 27386 7 1 2 76945 92789
0 27387 7 1 2 75150 27386
0 27388 7 1 2 27385 27387
0 27389 5 1 1 27388
0 27390 7 1 2 27366 27389
0 27391 5 1 1 27390
0 27392 7 1 2 71962 27391
0 27393 5 1 1 27392
0 27394 7 7 2 68184 69205
0 27395 7 3 2 64524 96829
0 27396 7 1 2 82625 96356
0 27397 5 1 1 27396
0 27398 7 2 2 78969 95713
0 27399 5 1 1 96839
0 27400 7 1 2 74157 96840
0 27401 5 1 1 27400
0 27402 7 1 2 27397 27401
0 27403 5 1 1 27402
0 27404 7 1 2 96836 27403
0 27405 5 1 1 27404
0 27406 7 1 2 69370 80050
0 27407 7 1 2 87087 27406
0 27408 7 1 2 88784 96701
0 27409 7 1 2 27407 27408
0 27410 5 1 1 27409
0 27411 7 1 2 27405 27410
0 27412 5 1 1 27411
0 27413 7 1 2 68421 27412
0 27414 5 1 1 27413
0 27415 7 4 2 87205 80650
0 27416 7 1 2 66738 96841
0 27417 7 1 2 96225 27416
0 27418 5 1 1 27417
0 27419 7 1 2 27414 27418
0 27420 5 1 1 27419
0 27421 7 1 2 65163 27420
0 27422 5 1 1 27421
0 27423 7 2 2 83059 80035
0 27424 7 1 2 96735 96845
0 27425 5 1 1 27424
0 27426 7 1 2 80607 95370
0 27427 7 1 2 95900 27426
0 27428 7 1 2 96121 27427
0 27429 5 1 1 27428
0 27430 7 1 2 27425 27429
0 27431 5 1 1 27430
0 27432 7 1 2 70925 27431
0 27433 5 1 1 27432
0 27434 7 1 2 76524 93042
0 27435 7 1 2 96846 27434
0 27436 5 1 1 27435
0 27437 7 1 2 27433 27436
0 27438 5 1 1 27437
0 27439 7 1 2 77663 27438
0 27440 5 1 1 27439
0 27441 7 1 2 27422 27440
0 27442 5 1 1 27441
0 27443 7 1 2 74809 27442
0 27444 5 1 1 27443
0 27445 7 1 2 72290 91172
0 27446 5 1 1 27445
0 27447 7 1 2 95959 96122
0 27448 5 1 1 27447
0 27449 7 1 2 27446 27448
0 27450 5 1 1 27449
0 27451 7 1 2 81346 81204
0 27452 7 1 2 27450 27451
0 27453 5 1 1 27452
0 27454 7 3 2 75453 85441
0 27455 7 2 2 61871 80150
0 27456 7 1 2 76578 87092
0 27457 7 1 2 96850 27456
0 27458 7 1 2 96847 27457
0 27459 5 1 1 27458
0 27460 7 1 2 27453 27459
0 27461 5 1 1 27460
0 27462 7 1 2 96141 27461
0 27463 5 1 1 27462
0 27464 7 1 2 27444 27463
0 27465 5 1 1 27464
0 27466 7 1 2 64946 27465
0 27467 5 1 1 27466
0 27468 7 3 2 68995 88253
0 27469 7 1 2 96238 96852
0 27470 5 1 1 27469
0 27471 7 1 2 95907 27470
0 27472 5 1 1 27471
0 27473 7 1 2 96770 27472
0 27474 5 1 1 27473
0 27475 7 5 2 70926 93105
0 27476 7 1 2 87206 86042
0 27477 7 1 2 78953 27476
0 27478 7 1 2 96855 27477
0 27479 5 1 1 27478
0 27480 7 1 2 27474 27479
0 27481 5 1 1 27480
0 27482 7 1 2 86583 27481
0 27483 5 1 1 27482
0 27484 7 3 2 78885 83415
0 27485 5 1 1 96860
0 27486 7 3 2 64134 93106
0 27487 7 1 2 91106 77664
0 27488 7 1 2 96863 27487
0 27489 7 1 2 96861 27488
0 27490 5 1 1 27489
0 27491 7 1 2 27483 27490
0 27492 5 1 1 27491
0 27493 7 1 2 89406 92309
0 27494 7 1 2 27492 27493
0 27495 5 1 1 27494
0 27496 7 1 2 27467 27495
0 27497 5 1 1 27496
0 27498 7 1 2 61595 27497
0 27499 5 1 1 27498
0 27500 7 2 2 73462 78195
0 27501 7 1 2 72850 96866
0 27502 5 1 1 27501
0 27503 7 1 2 77333 96304
0 27504 5 1 1 27503
0 27505 7 1 2 27502 27504
0 27506 5 1 1 27505
0 27507 7 1 2 68661 27506
0 27508 5 1 1 27507
0 27509 7 1 2 73756 77665
0 27510 5 1 1 27509
0 27511 7 1 2 27508 27510
0 27512 5 1 1 27511
0 27513 7 1 2 67263 27512
0 27514 5 1 1 27513
0 27515 7 1 2 75277 85043
0 27516 5 1 1 27515
0 27517 7 1 2 88322 27516
0 27518 5 1 1 27517
0 27519 7 1 2 27514 27518
0 27520 5 1 1 27519
0 27521 7 1 2 61872 84658
0 27522 7 1 2 27520 27521
0 27523 5 1 1 27522
0 27524 7 1 2 72062 96293
0 27525 5 1 1 27524
0 27526 7 1 2 96318 27525
0 27527 5 1 1 27526
0 27528 7 1 2 65164 85267
0 27529 7 1 2 27527 27528
0 27530 5 1 1 27529
0 27531 7 1 2 27523 27530
0 27532 5 1 1 27531
0 27533 7 1 2 96588 27532
0 27534 5 1 1 27533
0 27535 7 1 2 84948 94098
0 27536 5 1 1 27535
0 27537 7 1 2 90227 84547
0 27538 5 1 1 27537
0 27539 7 1 2 27536 27538
0 27540 5 1 1 27539
0 27541 7 1 2 70355 27540
0 27542 5 1 1 27541
0 27543 7 1 2 71334 76357
0 27544 5 1 1 27543
0 27545 7 1 2 85306 27544
0 27546 5 1 1 27545
0 27547 7 1 2 82969 27546
0 27548 5 1 1 27547
0 27549 7 1 2 27542 27548
0 27550 5 1 1 27549
0 27551 7 1 2 63575 27550
0 27552 5 1 1 27551
0 27553 7 1 2 77921 86897
0 27554 5 1 1 27553
0 27555 7 1 2 78125 27554
0 27556 5 1 1 27555
0 27557 7 1 2 70707 27556
0 27558 5 1 1 27557
0 27559 7 1 2 70084 93928
0 27560 5 1 1 27559
0 27561 7 1 2 27558 27560
0 27562 5 1 1 27561
0 27563 7 1 2 63969 27562
0 27564 5 1 1 27563
0 27565 7 1 2 79309 72629
0 27566 5 1 1 27565
0 27567 7 1 2 27564 27566
0 27568 5 1 1 27567
0 27569 7 1 2 71839 27568
0 27570 5 1 1 27569
0 27571 7 1 2 27552 27570
0 27572 5 1 1 27571
0 27573 7 1 2 62110 27572
0 27574 5 1 1 27573
0 27575 7 1 2 90514 85588
0 27576 5 1 1 27575
0 27577 7 1 2 27574 27576
0 27578 5 1 1 27577
0 27579 7 1 2 66739 27578
0 27580 5 1 1 27579
0 27581 7 2 2 72630 83761
0 27582 5 1 1 96868
0 27583 7 1 2 83881 27582
0 27584 5 1 1 27583
0 27585 7 1 2 67466 27584
0 27586 5 1 1 27585
0 27587 7 1 2 94346 27586
0 27588 5 1 1 27587
0 27589 7 1 2 71963 27588
0 27590 5 1 1 27589
0 27591 7 4 2 65992 72449
0 27592 5 1 1 96870
0 27593 7 1 2 84259 96871
0 27594 5 1 1 27593
0 27595 7 1 2 27590 27594
0 27596 5 1 1 27595
0 27597 7 1 2 61873 88323
0 27598 7 1 2 27596 27597
0 27599 5 1 1 27598
0 27600 7 1 2 27580 27599
0 27601 5 1 1 27600
0 27602 7 1 2 96390 27601
0 27603 5 1 1 27602
0 27604 7 1 2 27534 27603
0 27605 5 1 1 27604
0 27606 7 1 2 81387 27605
0 27607 5 1 1 27606
0 27608 7 1 2 75245 96483
0 27609 7 1 2 87306 27608
0 27610 5 1 1 27609
0 27611 7 1 2 82626 71579
0 27612 7 1 2 91739 27611
0 27613 7 1 2 93076 27612
0 27614 5 1 1 27613
0 27615 7 1 2 27610 27614
0 27616 5 1 1 27615
0 27617 7 1 2 72631 27616
0 27618 5 1 1 27617
0 27619 7 2 2 92289 93193
0 27620 7 1 2 88854 75774
0 27621 7 1 2 96874 27620
0 27622 5 1 1 27621
0 27623 7 1 2 80950 76209
0 27624 7 1 2 96459 27623
0 27625 5 1 1 27624
0 27626 7 1 2 27622 27625
0 27627 5 1 1 27626
0 27628 7 1 2 81455 27627
0 27629 5 1 1 27628
0 27630 7 1 2 27618 27629
0 27631 5 1 1 27630
0 27632 7 1 2 66493 27631
0 27633 5 1 1 27632
0 27634 7 4 2 61596 83121
0 27635 7 1 2 62111 93163
0 27636 7 1 2 91722 27635
0 27637 7 1 2 96154 27636
0 27638 7 1 2 96876 27637
0 27639 5 1 1 27638
0 27640 7 1 2 69575 27639
0 27641 7 1 2 27633 27640
0 27642 5 1 1 27641
0 27643 7 1 2 96793 96634
0 27644 5 1 1 27643
0 27645 7 1 2 82603 90476
0 27646 7 4 2 64135 64350
0 27647 7 1 2 96737 96880
0 27648 7 1 2 27645 27647
0 27649 7 1 2 87183 27648
0 27650 5 1 1 27649
0 27651 7 1 2 27644 27650
0 27652 5 1 1 27651
0 27653 7 1 2 63970 27652
0 27654 5 1 1 27653
0 27655 7 2 2 92790 96155
0 27656 7 1 2 96794 96884
0 27657 5 1 1 27656
0 27658 7 1 2 27654 27657
0 27659 5 1 1 27658
0 27660 7 1 2 63343 27659
0 27661 5 1 1 27660
0 27662 7 2 2 62112 95519
0 27663 5 1 1 96886
0 27664 7 1 2 81586 92791
0 27665 7 1 2 81009 27664
0 27666 7 1 2 96887 27665
0 27667 5 1 1 27666
0 27668 7 1 2 27661 27667
0 27669 5 1 1 27668
0 27670 7 1 2 70708 27669
0 27671 5 1 1 27670
0 27672 7 1 2 75541 91994
0 27673 7 1 2 96513 27672
0 27674 5 1 1 27673
0 27675 7 1 2 81010 96837
0 27676 7 1 2 94520 27675
0 27677 5 1 1 27676
0 27678 7 1 2 27674 27677
0 27679 5 1 1 27678
0 27680 7 1 2 75775 27679
0 27681 5 1 1 27680
0 27682 7 7 2 68422 84788
0 27683 5 1 1 96888
0 27684 7 3 2 66494 89669
0 27685 7 1 2 96889 96895
0 27686 7 1 2 96885 27685
0 27687 5 1 1 27686
0 27688 7 1 2 27681 27687
0 27689 7 1 2 27671 27688
0 27690 5 1 1 27689
0 27691 7 1 2 61874 27690
0 27692 5 1 1 27691
0 27693 7 6 2 64525 85589
0 27694 7 2 2 69206 96898
0 27695 7 1 2 88723 96904
0 27696 5 1 1 27695
0 27697 7 3 2 69371 78327
0 27698 7 4 2 64351 81637
0 27699 7 1 2 62113 63167
0 27700 7 1 2 96909 27699
0 27701 7 1 2 96906 27700
0 27702 5 1 1 27701
0 27703 7 1 2 27696 27702
0 27704 5 1 1 27703
0 27705 7 1 2 61597 27704
0 27706 5 1 1 27705
0 27707 7 1 2 76091 84252
0 27708 7 1 2 96905 27707
0 27709 5 1 1 27708
0 27710 7 1 2 27706 27709
0 27711 5 1 1 27710
0 27712 7 1 2 71439 27711
0 27713 5 1 1 27712
0 27714 7 1 2 64736 27713
0 27715 7 1 2 27692 27714
0 27716 5 1 1 27715
0 27717 7 1 2 27642 27716
0 27718 5 1 1 27717
0 27719 7 1 2 65165 27718
0 27720 5 1 1 27719
0 27721 7 1 2 94843 96234
0 27722 5 1 1 27721
0 27723 7 2 2 75151 71580
0 27724 5 2 1 96913
0 27725 7 1 2 84468 96519
0 27726 7 1 2 96914 27725
0 27727 5 1 1 27726
0 27728 7 1 2 27722 27727
0 27729 5 1 1 27728
0 27730 7 1 2 72632 27729
0 27731 5 1 1 27730
0 27732 7 1 2 75152 73213
0 27733 7 1 2 88576 96616
0 27734 7 1 2 27732 27733
0 27735 5 1 1 27734
0 27736 7 5 2 66740 64352
0 27737 7 1 2 90118 96917
0 27738 7 1 2 93079 27737
0 27739 7 1 2 96821 27738
0 27740 5 1 1 27739
0 27741 7 1 2 27735 27740
0 27742 7 1 2 27731 27741
0 27743 5 1 1 27742
0 27744 7 1 2 69811 27743
0 27745 5 1 1 27744
0 27746 7 1 2 62114 25868
0 27747 5 1 1 27746
0 27748 7 1 2 92044 93080
0 27749 7 1 2 96856 27748
0 27750 7 1 2 27747 27749
0 27751 5 1 1 27750
0 27752 7 1 2 27745 27751
0 27753 5 1 1 27752
0 27754 7 1 2 66495 27753
0 27755 5 1 1 27754
0 27756 7 1 2 62580 89751
0 27757 7 1 2 96881 27756
0 27758 7 1 2 82912 87565
0 27759 7 1 2 92723 27758
0 27760 7 1 2 27757 27759
0 27761 5 1 1 27760
0 27762 7 1 2 70085 27761
0 27763 7 1 2 27755 27762
0 27764 5 1 1 27763
0 27765 7 1 2 71840 27764
0 27766 7 1 2 27720 27765
0 27767 5 1 1 27766
0 27768 7 3 2 69576 80351
0 27769 7 1 2 96864 96922
0 27770 7 1 2 93199 27769
0 27771 5 1 1 27770
0 27772 7 1 2 65993 96678
0 27773 7 1 2 84253 27772
0 27774 7 1 2 95916 27773
0 27775 5 1 1 27774
0 27776 7 1 2 27771 27775
0 27777 5 1 1 27776
0 27778 7 1 2 92994 27777
0 27779 5 1 1 27778
0 27780 7 2 2 68423 69207
0 27781 7 5 2 64526 96925
0 27782 7 2 2 81818 96927
0 27783 7 3 2 73697 90119
0 27784 7 1 2 88863 96934
0 27785 7 1 2 96932 27784
0 27786 5 1 1 27785
0 27787 7 1 2 27779 27786
0 27788 5 1 1 27787
0 27789 7 1 2 89168 77871
0 27790 7 1 2 27788 27789
0 27791 5 1 1 27790
0 27792 7 1 2 27767 27791
0 27793 7 1 2 27607 27792
0 27794 7 1 2 27499 27793
0 27795 7 1 2 27393 27794
0 27796 7 1 2 27162 27795
0 27797 7 1 2 26918 27796
0 27798 7 1 2 26530 27797
0 27799 7 1 2 25906 27798
0 27800 5 1 1 27799
0 27801 7 16 2 61266 62952
0 27802 5 3 1 96937
0 27803 7 27 2 64254 96938
0 27804 7 1 2 27800 96956
0 27805 5 1 1 27804
0 27806 7 1 2 72346 95061
0 27807 5 1 1 27806
0 27808 7 1 2 72276 80912
0 27809 7 1 2 94889 27808
0 27810 5 1 1 27809
0 27811 7 1 2 27807 27810
0 27812 5 1 1 27811
0 27813 7 1 2 71964 27812
0 27814 5 1 1 27813
0 27815 7 1 2 80763 95066
0 27816 5 1 1 27815
0 27817 7 1 2 27814 27816
0 27818 5 1 1 27817
0 27819 7 1 2 70356 27818
0 27820 5 1 1 27819
0 27821 7 2 2 86569 82499
0 27822 7 1 2 64737 79847
0 27823 7 1 2 96983 27822
0 27824 5 1 1 27823
0 27825 7 1 2 27820 27824
0 27826 5 1 1 27825
0 27827 7 1 2 68850 27826
0 27828 5 1 1 27827
0 27829 7 1 2 65430 75385
0 27830 5 1 1 27829
0 27831 7 2 2 62416 83606
0 27832 5 1 1 96985
0 27833 7 1 2 27830 27832
0 27834 5 1 1 27833
0 27835 7 1 2 62844 82872
0 27836 7 1 2 27834 27835
0 27837 5 1 1 27836
0 27838 7 1 2 27828 27837
0 27839 5 1 1 27838
0 27840 7 1 2 63168 27839
0 27841 5 1 1 27840
0 27842 7 1 2 71965 91728
0 27843 5 1 1 27842
0 27844 7 1 2 2954 27843
0 27845 5 1 1 27844
0 27846 7 1 2 91400 94908
0 27847 7 1 2 27845 27846
0 27848 5 1 1 27847
0 27849 7 1 2 27841 27848
0 27850 5 1 1 27849
0 27851 7 1 2 68996 27850
0 27852 5 1 1 27851
0 27853 7 1 2 73068 89058
0 27854 5 1 1 27853
0 27855 7 1 2 72450 83233
0 27856 5 1 1 27855
0 27857 7 1 2 27854 27856
0 27858 5 1 1 27857
0 27859 7 1 2 89483 27858
0 27860 5 1 1 27859
0 27861 7 3 2 69577 72451
0 27862 7 2 2 81770 75876
0 27863 7 1 2 68424 96990
0 27864 7 1 2 96987 27863
0 27865 5 1 1 27864
0 27866 7 1 2 27860 27865
0 27867 5 1 1 27866
0 27868 7 1 2 71966 27867
0 27869 5 1 1 27868
0 27870 7 1 2 81128 80361
0 27871 7 1 2 87566 27870
0 27872 5 1 1 27871
0 27873 7 1 2 27869 27872
0 27874 5 1 1 27873
0 27875 7 1 2 72336 27874
0 27876 5 1 1 27875
0 27877 7 1 2 27852 27876
0 27878 5 1 1 27877
0 27879 7 1 2 61598 27878
0 27880 5 1 1 27879
0 27881 7 1 2 85748 86266
0 27882 5 1 1 27881
0 27883 7 1 2 79713 27882
0 27884 5 1 1 27883
0 27885 7 1 2 68997 27884
0 27886 5 1 1 27885
0 27887 7 1 2 65994 86629
0 27888 5 1 1 27887
0 27889 7 1 2 27886 27888
0 27890 5 1 1 27889
0 27891 7 1 2 70709 27890
0 27892 5 1 1 27891
0 27893 7 1 2 80276 80764
0 27894 5 1 1 27893
0 27895 7 1 2 27892 27894
0 27896 5 1 1 27895
0 27897 7 1 2 81638 91472
0 27898 7 1 2 27896 27897
0 27899 5 1 1 27898
0 27900 7 1 2 27880 27899
0 27901 5 1 1 27900
0 27902 7 1 2 67467 27901
0 27903 5 1 1 27902
0 27904 7 1 2 5419 95140
0 27905 5 1 1 27904
0 27906 7 1 2 76637 83611
0 27907 5 1 1 27906
0 27908 7 1 2 68998 27907
0 27909 7 1 2 27905 27908
0 27910 5 1 1 27909
0 27911 7 2 2 76525 93292
0 27912 5 1 1 96992
0 27913 7 1 2 70927 76621
0 27914 7 1 2 96993 27913
0 27915 5 1 1 27914
0 27916 7 1 2 27910 27915
0 27917 5 1 1 27916
0 27918 7 1 2 86956 27917
0 27919 5 1 1 27918
0 27920 7 1 2 65766 79490
0 27921 5 2 1 27920
0 27922 7 1 2 86713 96994
0 27923 5 1 1 27922
0 27924 7 1 2 81924 83607
0 27925 7 1 2 27923 27924
0 27926 5 1 1 27925
0 27927 7 1 2 27919 27926
0 27928 5 1 1 27927
0 27929 7 1 2 62417 27928
0 27930 5 1 1 27929
0 27931 7 7 2 64738 86671
0 27932 7 1 2 80892 6871
0 27933 5 1 1 27932
0 27934 7 1 2 62845 27933
0 27935 5 1 1 27934
0 27936 7 1 2 75223 95136
0 27937 5 1 1 27936
0 27938 7 1 2 27935 27937
0 27939 5 1 1 27938
0 27940 7 1 2 68999 27939
0 27941 5 1 1 27940
0 27942 7 1 2 74533 85346
0 27943 5 1 1 27942
0 27944 7 1 2 27941 27943
0 27945 5 1 1 27944
0 27946 7 1 2 67264 27945
0 27947 5 1 1 27946
0 27948 7 2 2 74492 75327
0 27949 5 3 1 97003
0 27950 7 1 2 85945 97004
0 27951 5 1 1 27950
0 27952 7 1 2 27947 27951
0 27953 5 1 1 27952
0 27954 7 1 2 96996 27953
0 27955 5 1 1 27954
0 27956 7 1 2 27930 27955
0 27957 5 1 1 27956
0 27958 7 1 2 63576 27957
0 27959 5 1 1 27958
0 27960 7 2 2 90005 74453
0 27961 7 1 2 74938 80166
0 27962 7 1 2 91044 27961
0 27963 7 1 2 97008 27962
0 27964 5 1 1 27963
0 27965 7 1 2 27959 27964
0 27966 5 1 1 27965
0 27967 7 1 2 82665 27966
0 27968 5 1 1 27967
0 27969 7 1 2 27903 27968
0 27970 5 1 1 27969
0 27971 7 1 2 93107 27970
0 27972 5 1 1 27971
0 27973 7 10 2 71335 73069
0 27974 5 4 1 97010
0 27975 7 1 2 72492 97020
0 27976 5 2 1 27975
0 27977 7 1 2 74123 97024
0 27978 5 1 1 27977
0 27979 7 1 2 79239 94342
0 27980 5 1 1 27979
0 27981 7 1 2 27978 27980
0 27982 5 1 1 27981
0 27983 7 1 2 70928 27982
0 27984 5 1 1 27983
0 27985 7 1 2 77526 86832
0 27986 5 1 1 27985
0 27987 7 1 2 71683 27986
0 27988 5 1 1 27987
0 27989 7 1 2 70357 27988
0 27990 5 1 1 27989
0 27991 7 1 2 27984 27990
0 27992 5 1 1 27991
0 27993 7 1 2 79820 82849
0 27994 7 1 2 92115 27993
0 27995 7 1 2 89650 27994
0 27996 7 1 2 27992 27995
0 27997 5 1 1 27996
0 27998 7 1 2 27972 27997
0 27999 5 1 1 27998
0 28000 7 1 2 64947 27999
0 28001 5 1 1 28000
0 28002 7 2 2 88466 82240
0 28003 7 5 2 90745 91780
0 28004 7 1 2 62115 90477
0 28005 7 1 2 74984 28004
0 28006 7 1 2 73622 28005
0 28007 7 2 2 97028 28006
0 28008 7 1 2 97026 97033
0 28009 5 1 1 28008
0 28010 7 1 2 61875 28009
0 28011 7 1 2 28001 28010
0 28012 5 1 1 28011
0 28013 7 1 2 72162 91532
0 28014 5 1 1 28013
0 28015 7 1 2 17400 28014
0 28016 5 1 1 28015
0 28017 7 6 2 87662 93108
0 28018 7 1 2 28016 97035
0 28019 5 1 1 28018
0 28020 7 1 2 71018 92360
0 28021 5 1 1 28020
0 28022 7 1 2 17782 28021
0 28023 5 1 1 28022
0 28024 7 1 2 81819 96572
0 28025 7 1 2 28023 28024
0 28026 5 1 1 28025
0 28027 7 1 2 28019 28026
0 28028 5 1 1 28027
0 28029 7 1 2 70710 28028
0 28030 5 1 1 28029
0 28031 7 2 2 61599 74079
0 28032 7 3 2 82423 75435
0 28033 7 1 2 91188 97043
0 28034 7 1 2 97041 28033
0 28035 5 1 1 28034
0 28036 7 1 2 17404 25731
0 28037 5 2 1 28036
0 28038 7 1 2 65767 97046
0 28039 5 1 1 28038
0 28040 7 2 2 84569 93278
0 28041 5 1 1 97048
0 28042 7 1 2 28039 28041
0 28043 5 1 1 28042
0 28044 7 1 2 87646 89202
0 28045 7 1 2 28043 28044
0 28046 5 1 1 28045
0 28047 7 1 2 28035 28046
0 28048 5 1 1 28047
0 28049 7 1 2 62418 28048
0 28050 5 1 1 28049
0 28051 7 1 2 82882 80628
0 28052 7 1 2 71532 75184
0 28053 7 1 2 78779 28052
0 28054 7 1 2 28051 28053
0 28055 5 1 1 28054
0 28056 7 1 2 28050 28055
0 28057 5 1 1 28056
0 28058 7 1 2 96142 28057
0 28059 5 1 1 28058
0 28060 7 1 2 28030 28059
0 28061 5 1 1 28060
0 28062 7 1 2 66965 28061
0 28063 5 1 1 28062
0 28064 7 2 2 80788 78886
0 28065 7 1 2 91138 97050
0 28066 5 1 1 28065
0 28067 7 1 2 69000 96474
0 28068 5 1 1 28067
0 28069 7 1 2 65995 94648
0 28070 5 1 1 28069
0 28071 7 1 2 28068 28070
0 28072 5 1 1 28071
0 28073 7 1 2 73017 28072
0 28074 5 1 1 28073
0 28075 7 1 2 28066 28074
0 28076 5 1 1 28075
0 28077 7 1 2 84529 93109
0 28078 7 1 2 76418 28077
0 28079 7 1 2 28076 28078
0 28080 5 1 1 28079
0 28081 7 1 2 28063 28080
0 28082 5 1 1 28081
0 28083 7 1 2 70358 28082
0 28084 5 1 1 28083
0 28085 7 2 2 65431 93110
0 28086 7 2 2 84533 97052
0 28087 7 4 2 80244 87142
0 28088 7 2 2 73018 73948
0 28089 5 1 1 97060
0 28090 7 1 2 67695 73885
0 28091 5 1 1 28090
0 28092 7 1 2 28089 28091
0 28093 5 2 1 28092
0 28094 7 1 2 97056 97062
0 28095 5 1 1 28094
0 28096 7 1 2 71492 78328
0 28097 7 1 2 73979 28096
0 28098 5 1 1 28097
0 28099 7 1 2 84303 76412
0 28100 5 1 1 28099
0 28101 7 2 2 72163 85930
0 28102 5 1 1 97064
0 28103 7 1 2 71623 28102
0 28104 7 1 2 28100 28103
0 28105 5 1 1 28104
0 28106 7 1 2 28098 28105
0 28107 5 1 1 28106
0 28108 7 1 2 86957 28107
0 28109 5 1 1 28108
0 28110 7 1 2 28095 28109
0 28111 5 1 1 28110
0 28112 7 1 2 97054 28111
0 28113 5 1 1 28112
0 28114 7 1 2 28084 28113
0 28115 5 1 1 28114
0 28116 7 1 2 67468 28115
0 28117 5 1 1 28116
0 28118 7 1 2 74124 97036
0 28119 5 1 1 28118
0 28120 7 1 2 71637 92511
0 28121 7 1 2 96928 28120
0 28122 5 1 1 28121
0 28123 7 1 2 28119 28122
0 28124 5 1 1 28123
0 28125 7 1 2 68851 28124
0 28126 5 1 1 28125
0 28127 7 1 2 75290 86118
0 28128 7 1 2 96933 28127
0 28129 5 1 1 28128
0 28130 7 1 2 28126 28129
0 28131 5 1 1 28130
0 28132 7 1 2 70929 28131
0 28133 5 1 1 28132
0 28134 7 2 2 63971 65996
0 28135 5 2 1 97066
0 28136 7 2 2 62581 74080
0 28137 5 1 1 97070
0 28138 7 1 2 97068 28137
0 28139 5 1 1 28138
0 28140 7 1 2 97037 28139
0 28141 5 1 1 28140
0 28142 7 1 2 28133 28141
0 28143 5 1 1 28142
0 28144 7 1 2 81925 28143
0 28145 5 1 1 28144
0 28146 7 1 2 87044 95228
0 28147 5 1 1 28146
0 28148 7 1 2 97038 28147
0 28149 5 1 1 28148
0 28150 7 2 2 82718 96239
0 28151 7 1 2 79225 74525
0 28152 7 1 2 97072 28151
0 28153 5 1 1 28152
0 28154 7 1 2 28149 28153
0 28155 5 1 1 28154
0 28156 7 1 2 86958 28155
0 28157 5 1 1 28156
0 28158 7 1 2 28145 28157
0 28159 5 1 1 28158
0 28160 7 1 2 72851 28159
0 28161 5 1 1 28160
0 28162 7 1 2 71127 91682
0 28163 5 1 1 28162
0 28164 7 1 2 82533 93267
0 28165 5 1 1 28164
0 28166 7 1 2 64136 74844
0 28167 7 1 2 28165 28166
0 28168 5 1 1 28167
0 28169 7 1 2 28163 28168
0 28170 5 1 1 28169
0 28171 7 1 2 81926 28170
0 28172 5 1 1 28171
0 28173 7 1 2 73019 97049
0 28174 5 1 1 28173
0 28175 7 1 2 28172 28174
0 28176 5 1 1 28175
0 28177 7 1 2 70930 28176
0 28178 5 1 1 28177
0 28179 7 1 2 88061 94833
0 28180 5 1 1 28179
0 28181 7 1 2 28178 28180
0 28182 5 1 1 28181
0 28183 7 1 2 97055 28182
0 28184 5 1 1 28183
0 28185 7 1 2 28161 28184
0 28186 5 1 1 28185
0 28187 7 1 2 65768 28186
0 28188 5 1 1 28187
0 28189 7 1 2 71711 97047
0 28190 5 1 1 28189
0 28191 7 1 2 81070 94828
0 28192 5 2 1 28191
0 28193 7 1 2 28190 97074
0 28194 5 1 1 28193
0 28195 7 1 2 65432 28194
0 28196 5 1 1 28195
0 28197 7 5 2 69578 88625
0 28198 5 1 1 97076
0 28199 7 1 2 95484 97077
0 28200 5 1 1 28199
0 28201 7 1 2 28196 28200
0 28202 5 1 1 28201
0 28203 7 1 2 70711 28202
0 28204 5 1 1 28203
0 28205 7 1 2 14278 94436
0 28206 5 1 1 28205
0 28207 7 1 2 80151 96738
0 28208 7 1 2 28206 28207
0 28209 5 1 1 28208
0 28210 7 1 2 28204 28209
0 28211 5 1 1 28210
0 28212 7 1 2 86611 28211
0 28213 5 1 1 28212
0 28214 7 1 2 86959 85532
0 28215 5 1 1 28214
0 28216 7 1 2 72063 97078
0 28217 5 1 1 28216
0 28218 7 1 2 28215 28217
0 28219 5 1 1 28218
0 28220 7 1 2 85031 74466
0 28221 7 1 2 28219 28220
0 28222 5 1 1 28221
0 28223 7 1 2 28213 28222
0 28224 5 1 1 28223
0 28225 7 1 2 63805 28224
0 28226 5 1 1 28225
0 28227 7 1 2 71493 74467
0 28228 7 1 2 87357 28227
0 28229 7 1 2 95366 28228
0 28230 5 1 1 28229
0 28231 7 1 2 28226 28230
0 28232 5 1 1 28231
0 28233 7 1 2 90969 28232
0 28234 5 1 1 28233
0 28235 7 1 2 28188 28234
0 28236 7 1 2 28117 28235
0 28237 5 1 1 28236
0 28238 7 1 2 69812 28237
0 28239 5 1 1 28238
0 28240 7 4 2 78476 93111
0 28241 7 1 2 97034 97081
0 28242 5 1 1 28241
0 28243 7 1 2 66741 28242
0 28244 7 1 2 28239 28243
0 28245 5 1 1 28244
0 28246 7 1 2 70086 28245
0 28247 7 1 2 28012 28246
0 28248 5 1 1 28247
0 28249 7 1 2 64353 85896
0 28250 7 2 2 95022 28249
0 28251 7 1 2 74081 97085
0 28252 5 1 1 28251
0 28253 7 1 2 77504 96492
0 28254 5 1 1 28253
0 28255 7 1 2 89520 96498
0 28256 5 1 1 28255
0 28257 7 1 2 28254 28256
0 28258 5 1 1 28257
0 28259 7 1 2 76161 28258
0 28260 5 1 1 28259
0 28261 7 1 2 72164 96599
0 28262 5 1 1 28261
0 28263 7 1 2 72556 96391
0 28264 5 1 1 28263
0 28265 7 1 2 28262 28264
0 28266 5 1 1 28265
0 28267 7 1 2 79180 28266
0 28268 5 1 1 28267
0 28269 7 1 2 28260 28268
0 28270 5 1 1 28269
0 28271 7 1 2 71240 28270
0 28272 5 1 1 28271
0 28273 7 1 2 28252 28272
0 28274 5 1 1 28273
0 28275 7 1 2 86418 28274
0 28276 5 1 1 28275
0 28277 7 1 2 62582 84384
0 28278 5 2 1 28277
0 28279 7 1 2 96669 97087
0 28280 5 2 1 28279
0 28281 7 1 2 76162 97089
0 28282 5 1 1 28281
0 28283 7 1 2 76048 89845
0 28284 5 1 1 28283
0 28285 7 1 2 28282 28284
0 28286 5 1 1 28285
0 28287 7 1 2 64739 28286
0 28288 5 1 1 28287
0 28289 7 6 2 62846 65997
0 28290 5 1 1 97091
0 28291 7 1 2 79491 97092
0 28292 7 1 2 92531 28291
0 28293 5 1 1 28292
0 28294 7 1 2 28288 28293
0 28295 5 1 1 28294
0 28296 7 1 2 92792 28295
0 28297 5 1 1 28296
0 28298 7 3 2 85615 95229
0 28299 5 1 1 97097
0 28300 7 1 2 87045 97098
0 28301 5 3 1 28300
0 28302 7 1 2 96673 97100
0 28303 5 1 1 28302
0 28304 7 1 2 28297 28303
0 28305 5 1 1 28304
0 28306 7 1 2 78842 28305
0 28307 5 1 1 28306
0 28308 7 1 2 91944 93112
0 28309 7 1 2 97101 28308
0 28310 5 1 1 28309
0 28311 7 1 2 84404 96617
0 28312 7 1 2 97090 28311
0 28313 5 1 1 28312
0 28314 7 1 2 28310 28313
0 28315 5 1 1 28314
0 28316 7 1 2 81993 28315
0 28317 5 1 1 28316
0 28318 7 1 2 28307 28317
0 28319 5 1 1 28318
0 28320 7 1 2 65769 28319
0 28321 5 1 1 28320
0 28322 7 1 2 66742 78711
0 28323 7 1 2 96802 28322
0 28324 5 1 1 28323
0 28325 7 1 2 61876 88855
0 28326 7 1 2 96875 28325
0 28327 5 1 1 28326
0 28328 7 1 2 28324 28327
0 28329 5 1 1 28328
0 28330 7 1 2 67696 28329
0 28331 5 1 1 28330
0 28332 7 4 2 68018 96698
0 28333 7 1 2 85533 97103
0 28334 5 1 1 28333
0 28335 7 1 2 74520 84935
0 28336 5 2 1 28335
0 28337 7 5 2 81994 96143
0 28338 5 1 1 97109
0 28339 7 1 2 97107 97110
0 28340 5 1 1 28339
0 28341 7 1 2 28334 28340
0 28342 7 1 2 28331 28341
0 28343 5 1 1 28342
0 28344 7 1 2 86960 28343
0 28345 5 1 1 28344
0 28346 7 2 2 72754 77527
0 28347 7 1 2 97104 97114
0 28348 5 1 1 28347
0 28349 7 1 2 72165 97111
0 28350 5 1 1 28349
0 28351 7 1 2 28348 28350
0 28352 5 1 1 28351
0 28353 7 1 2 70712 28352
0 28354 5 1 1 28353
0 28355 7 1 2 87043 97112
0 28356 5 1 1 28355
0 28357 7 1 2 28354 28356
0 28358 5 1 1 28357
0 28359 7 1 2 81927 28358
0 28360 5 1 1 28359
0 28361 7 1 2 28345 28360
0 28362 5 1 1 28361
0 28363 7 1 2 67469 28362
0 28364 5 1 1 28363
0 28365 7 1 2 87048 88110
0 28366 5 3 1 28365
0 28367 7 3 2 88467 91517
0 28368 5 3 1 97119
0 28369 7 1 2 97116 97120
0 28370 5 1 1 28369
0 28371 7 1 2 91245 74521
0 28372 5 1 1 28371
0 28373 7 1 2 81669 93043
0 28374 7 1 2 28372 28373
0 28375 5 1 1 28374
0 28376 7 1 2 28370 28375
0 28377 5 1 1 28376
0 28378 7 1 2 87246 28377
0 28379 5 1 1 28378
0 28380 7 1 2 87358 75706
0 28381 7 1 2 96430 28380
0 28382 7 1 2 85534 28381
0 28383 5 1 1 28382
0 28384 7 1 2 28379 28383
0 28385 7 1 2 28364 28384
0 28386 7 1 2 28321 28385
0 28387 5 1 1 28386
0 28388 7 1 2 65433 28387
0 28389 5 1 1 28388
0 28390 7 1 2 28276 28389
0 28391 5 1 1 28390
0 28392 7 1 2 70087 28391
0 28393 5 1 1 28392
0 28394 7 1 2 96739 27295
0 28395 5 1 1 28394
0 28396 7 1 2 81250 80814
0 28397 5 1 1 28396
0 28398 7 1 2 28395 28397
0 28399 5 1 1 28398
0 28400 7 1 2 93113 28399
0 28401 5 1 1 28400
0 28402 7 1 2 66496 74183
0 28403 7 1 2 96176 28402
0 28404 5 1 1 28403
0 28405 7 1 2 28401 28404
0 28406 5 1 1 28405
0 28407 7 1 2 81995 28406
0 28408 5 1 1 28407
0 28409 7 1 2 74184 78843
0 28410 7 1 2 96189 28409
0 28411 5 1 1 28410
0 28412 7 1 2 28408 28411
0 28413 5 1 1 28412
0 28414 7 1 2 64137 28413
0 28415 5 1 1 28414
0 28416 7 2 2 64948 74185
0 28417 7 1 2 91540 96177
0 28418 7 1 2 97125 28417
0 28419 5 1 1 28418
0 28420 7 1 2 28415 28419
0 28421 5 1 1 28420
0 28422 7 1 2 71336 28421
0 28423 5 1 1 28422
0 28424 7 1 2 81655 92793
0 28425 7 1 2 89759 28424
0 28426 5 1 1 28425
0 28427 7 1 2 28338 28426
0 28428 5 1 1 28427
0 28429 7 1 2 90573 28428
0 28430 5 1 1 28429
0 28431 7 1 2 25049 97122
0 28432 5 1 1 28431
0 28433 7 2 2 87247 28432
0 28434 7 1 2 78329 97127
0 28435 5 1 1 28434
0 28436 7 1 2 95480 96484
0 28437 7 1 2 96923 28436
0 28438 5 1 1 28437
0 28439 7 1 2 28435 28438
0 28440 7 1 2 28430 28439
0 28441 5 1 1 28440
0 28442 7 1 2 73326 28441
0 28443 5 1 1 28442
0 28444 7 1 2 28423 28443
0 28445 5 1 1 28444
0 28446 7 1 2 76946 28445
0 28447 5 1 1 28446
0 28448 7 1 2 28393 28447
0 28449 5 1 1 28448
0 28450 7 1 2 73020 28449
0 28451 5 1 1 28450
0 28452 7 1 2 73327 85406
0 28453 5 2 1 28452
0 28454 7 1 2 76609 97129
0 28455 5 2 1 28454
0 28456 7 1 2 93442 97131
0 28457 5 1 1 28456
0 28458 7 1 2 86961 91094
0 28459 5 1 1 28458
0 28460 7 1 2 63806 92151
0 28461 5 1 1 28460
0 28462 7 1 2 28459 28461
0 28463 5 1 1 28462
0 28464 7 4 2 70088 86701
0 28465 7 1 2 71241 97133
0 28466 7 1 2 28463 28465
0 28467 5 1 1 28466
0 28468 7 1 2 28457 28467
0 28469 5 1 1 28468
0 28470 7 1 2 67697 28469
0 28471 5 1 1 28470
0 28472 7 1 2 65166 76324
0 28473 7 1 2 80475 87111
0 28474 7 1 2 28472 28473
0 28475 7 1 2 80843 28474
0 28476 5 1 1 28475
0 28477 7 1 2 28471 28476
0 28478 5 1 1 28477
0 28479 7 1 2 69813 28478
0 28480 5 1 1 28479
0 28481 7 4 2 80532 86289
0 28482 5 1 1 97137
0 28483 7 1 2 93261 95240
0 28484 7 1 2 97138 28483
0 28485 5 1 1 28484
0 28486 7 1 2 28480 28485
0 28487 5 1 1 28486
0 28488 7 1 2 61877 28487
0 28489 5 1 1 28488
0 28490 7 2 2 75685 82308
0 28491 7 1 2 90427 97141
0 28492 7 1 2 86702 28491
0 28493 7 1 2 91433 28492
0 28494 5 1 1 28493
0 28495 7 1 2 28489 28494
0 28496 5 1 1 28495
0 28497 7 1 2 63169 28496
0 28498 5 1 1 28497
0 28499 7 2 2 65434 97134
0 28500 7 1 2 80460 82956
0 28501 7 1 2 96332 28500
0 28502 7 1 2 97143 28501
0 28503 5 1 1 28502
0 28504 7 1 2 28498 28503
0 28505 5 1 1 28504
0 28506 7 1 2 93114 28505
0 28507 5 1 1 28506
0 28508 7 1 2 28451 28507
0 28509 5 1 1 28508
0 28510 7 1 2 92703 28509
0 28511 5 1 1 28510
0 28512 7 4 2 71337 93624
0 28513 7 2 2 78954 82902
0 28514 7 2 2 97145 97149
0 28515 7 1 2 74278 97151
0 28516 5 1 1 28515
0 28517 7 2 2 77473 92614
0 28518 7 1 2 95909 97153
0 28519 5 1 1 28518
0 28520 7 1 2 28516 28519
0 28521 5 1 1 28520
0 28522 7 1 2 67265 28521
0 28523 5 1 1 28522
0 28524 7 1 2 93348 97152
0 28525 5 1 1 28524
0 28526 7 1 2 28523 28525
0 28527 5 1 1 28526
0 28528 7 1 2 66966 28527
0 28529 5 1 1 28528
0 28530 7 1 2 80283 96538
0 28531 7 1 2 88492 28530
0 28532 7 1 2 97150 28531
0 28533 5 1 1 28532
0 28534 7 1 2 28529 28533
0 28535 5 1 1 28534
0 28536 7 1 2 61878 28535
0 28537 5 1 1 28536
0 28538 7 4 2 75153 75722
0 28539 7 1 2 79101 90959
0 28540 7 1 2 91900 28539
0 28541 7 1 2 97155 28540
0 28542 5 1 1 28541
0 28543 7 1 2 28537 28542
0 28544 5 1 1 28543
0 28545 7 1 2 70089 28544
0 28546 5 1 1 28545
0 28547 7 1 2 73021 80709
0 28548 7 1 2 75723 28547
0 28549 7 4 2 62116 96102
0 28550 7 1 2 87248 97159
0 28551 7 1 2 28548 28550
0 28552 5 1 1 28551
0 28553 7 1 2 28546 28552
0 28554 5 1 1 28553
0 28555 7 1 2 68185 28554
0 28556 5 1 1 28555
0 28557 7 3 2 87065 95990
0 28558 5 2 1 97163
0 28559 7 1 2 94989 97166
0 28560 5 6 1 28559
0 28561 7 1 2 66967 97168
0 28562 5 1 1 28561
0 28563 7 1 2 75111 82038
0 28564 5 1 1 28563
0 28565 7 1 2 28562 28564
0 28566 5 1 1 28565
0 28567 7 1 2 76671 28566
0 28568 5 1 1 28567
0 28569 7 2 2 81996 78824
0 28570 7 1 2 80355 97174
0 28571 5 1 1 28570
0 28572 7 1 2 28568 28571
0 28573 5 1 1 28572
0 28574 7 1 2 88916 93625
0 28575 7 1 2 88493 28574
0 28576 7 1 2 28573 28575
0 28577 5 1 1 28576
0 28578 7 1 2 28556 28577
0 28579 5 1 1 28578
0 28580 7 1 2 62847 28579
0 28581 5 1 1 28580
0 28582 7 1 2 84999 87923
0 28583 7 1 2 90917 78975
0 28584 7 1 2 97044 28583
0 28585 7 1 2 28582 28584
0 28586 5 1 1 28585
0 28587 7 1 2 28581 28586
0 28588 5 1 1 28587
0 28589 7 1 2 70359 28588
0 28590 5 1 1 28589
0 28591 7 1 2 63807 81358
0 28592 7 1 2 94823 28591
0 28593 7 1 2 97146 28592
0 28594 5 1 1 28593
0 28595 7 1 2 80879 78712
0 28596 7 1 2 92794 28595
0 28597 7 1 2 85543 28596
0 28598 5 1 1 28597
0 28599 7 1 2 28594 28598
0 28600 5 1 1 28599
0 28601 7 1 2 63577 28600
0 28602 5 1 1 28601
0 28603 7 1 2 78240 96618
0 28604 7 1 2 97154 28603
0 28605 5 1 1 28604
0 28606 7 1 2 28602 28605
0 28607 5 1 1 28606
0 28608 7 1 2 62419 28607
0 28609 5 1 1 28608
0 28610 7 1 2 75514 91697
0 28611 7 1 2 92615 96403
0 28612 7 1 2 28610 28611
0 28613 5 1 1 28612
0 28614 7 1 2 28609 28613
0 28615 5 1 1 28614
0 28616 7 1 2 66968 28615
0 28617 5 1 1 28616
0 28618 7 2 2 73022 73260
0 28619 7 2 2 78678 92795
0 28620 7 1 2 95400 97178
0 28621 7 1 2 97176 28620
0 28622 5 1 1 28621
0 28623 7 1 2 28617 28622
0 28624 5 1 1 28623
0 28625 7 1 2 63344 28624
0 28626 5 1 1 28625
0 28627 7 2 2 94050 96194
0 28628 7 1 2 82077 94867
0 28629 7 1 2 97180 28628
0 28630 7 1 2 97177 28629
0 28631 5 1 1 28630
0 28632 7 1 2 28626 28631
0 28633 5 1 1 28632
0 28634 7 1 2 73698 88119
0 28635 7 1 2 28633 28634
0 28636 5 1 1 28635
0 28637 7 1 2 61600 28636
0 28638 7 1 2 28590 28637
0 28639 5 1 1 28638
0 28640 7 1 2 82547 96583
0 28641 5 1 1 28640
0 28642 7 1 2 90409 96485
0 28643 5 1 1 28642
0 28644 7 1 2 28641 28643
0 28645 5 1 1 28644
0 28646 7 1 2 61879 28645
0 28647 5 1 1 28646
0 28648 7 1 2 81771 96499
0 28649 5 1 1 28648
0 28650 7 1 2 28647 28649
0 28651 5 1 1 28650
0 28652 7 1 2 93483 97156
0 28653 7 1 2 28651 28652
0 28654 5 1 1 28653
0 28655 7 2 2 87249 92704
0 28656 7 2 2 65167 85084
0 28657 7 1 2 88494 97184
0 28658 7 1 2 97182 28657
0 28659 5 1 1 28658
0 28660 7 2 2 64949 90195
0 28661 7 1 2 88713 90888
0 28662 7 1 2 97186 28661
0 28663 5 1 1 28662
0 28664 7 1 2 28659 28663
0 28665 5 1 1 28664
0 28666 7 1 2 93044 28665
0 28667 5 1 1 28666
0 28668 7 2 2 82793 87856
0 28669 7 2 2 85053 97188
0 28670 7 1 2 82627 87663
0 28671 7 1 2 97190 28670
0 28672 5 1 1 28671
0 28673 7 1 2 28667 28672
0 28674 7 1 2 28654 28673
0 28675 5 1 1 28674
0 28676 7 1 2 70360 28675
0 28677 5 1 1 28676
0 28678 7 4 2 64527 88120
0 28679 7 1 2 85566 97192
0 28680 7 2 2 69208 73023
0 28681 7 1 2 87250 97196
0 28682 7 1 2 28679 28681
0 28683 7 1 2 94887 28682
0 28684 5 1 1 28683
0 28685 7 1 2 28677 28684
0 28686 5 1 1 28685
0 28687 7 1 2 62848 28686
0 28688 5 1 1 28687
0 28689 7 2 2 73623 82039
0 28690 5 1 1 97198
0 28691 7 3 2 79080 76708
0 28692 7 1 2 80773 97200
0 28693 5 1 1 28692
0 28694 7 1 2 28690 28693
0 28695 5 2 1 28694
0 28696 7 1 2 81456 97203
0 28697 5 1 1 28696
0 28698 7 1 2 83339 90794
0 28699 7 1 2 92896 28698
0 28700 5 1 1 28699
0 28701 7 1 2 28697 28700
0 28702 5 1 1 28701
0 28703 7 1 2 75154 28702
0 28704 5 1 1 28703
0 28705 7 3 2 65435 92705
0 28706 7 3 2 65770 97205
0 28707 7 1 2 66743 90428
0 28708 7 1 2 97208 28707
0 28709 5 1 1 28708
0 28710 7 1 2 28704 28709
0 28711 5 1 1 28710
0 28712 7 1 2 74143 28711
0 28713 5 1 1 28712
0 28714 7 1 2 72452 73688
0 28715 7 1 2 85000 28714
0 28716 7 1 2 86095 81563
0 28717 7 1 2 28715 28716
0 28718 5 1 1 28717
0 28719 7 1 2 28713 28718
0 28720 5 1 1 28719
0 28721 7 1 2 96619 28720
0 28722 5 1 1 28721
0 28723 7 1 2 66497 28722
0 28724 7 1 2 28688 28723
0 28725 5 1 1 28724
0 28726 7 1 2 72633 28725
0 28727 7 1 2 28639 28726
0 28728 5 1 1 28727
0 28729 7 1 2 28511 28728
0 28730 7 1 2 85021 80491
0 28731 5 2 1 28730
0 28732 7 1 2 95062 21191
0 28733 5 1 1 28732
0 28734 7 1 2 81997 28733
0 28735 5 1 1 28734
0 28736 7 1 2 97211 28735
0 28737 5 1 1 28736
0 28738 7 1 2 61601 28737
0 28739 5 1 1 28738
0 28740 7 2 2 81899 95328
0 28741 7 1 2 84123 97213
0 28742 5 1 1 28741
0 28743 7 1 2 28739 28742
0 28744 5 1 1 28743
0 28745 7 1 2 78014 28744
0 28746 5 1 1 28745
0 28747 7 1 2 78313 81900
0 28748 7 1 2 94991 28747
0 28749 5 1 1 28748
0 28750 7 1 2 28746 28749
0 28751 5 1 1 28750
0 28752 7 1 2 74810 28751
0 28753 5 1 1 28752
0 28754 7 1 2 90587 92757
0 28755 7 1 2 95666 28754
0 28756 7 1 2 83322 28755
0 28757 5 1 1 28756
0 28758 7 1 2 28753 28757
0 28759 5 1 1 28758
0 28760 7 1 2 68852 28759
0 28761 5 1 1 28760
0 28762 7 2 2 76325 92988
0 28763 7 1 2 86612 87207
0 28764 7 1 2 75336 28763
0 28765 7 1 2 97215 28764
0 28766 5 1 1 28765
0 28767 7 1 2 28761 28766
0 28768 5 1 1 28767
0 28769 7 1 2 67470 28768
0 28770 5 1 1 28769
0 28771 7 1 2 84176 97126
0 28772 5 1 1 28771
0 28773 7 2 2 75877 78369
0 28774 7 1 2 69814 97217
0 28775 5 1 1 28774
0 28776 7 1 2 28772 28775
0 28777 5 1 1 28776
0 28778 7 1 2 83340 28777
0 28779 5 1 1 28778
0 28780 7 1 2 82628 71019
0 28781 7 1 2 81221 28780
0 28782 5 1 1 28781
0 28783 7 1 2 28779 28782
0 28784 5 1 1 28783
0 28785 7 1 2 61602 28784
0 28786 5 1 1 28785
0 28787 7 1 2 82015 97218
0 28788 5 1 1 28787
0 28789 7 1 2 28786 28788
0 28790 5 1 1 28789
0 28791 7 1 2 88225 28790
0 28792 5 1 1 28791
0 28793 7 1 2 28770 28792
0 28794 5 1 1 28793
0 28795 7 1 2 65436 28794
0 28796 5 1 1 28795
0 28797 7 1 2 72790 92502
0 28798 5 1 1 28797
0 28799 7 1 2 88499 28798
0 28800 5 1 1 28799
0 28801 7 1 2 76860 28800
0 28802 5 1 1 28801
0 28803 7 1 2 75676 73163
0 28804 7 1 2 92157 28803
0 28805 5 1 1 28804
0 28806 7 1 2 28802 28805
0 28807 5 1 1 28806
0 28808 7 1 2 70713 28807
0 28809 5 1 1 28808
0 28810 7 1 2 89828 74417
0 28811 5 1 1 28810
0 28812 7 1 2 28809 28811
0 28813 5 1 1 28812
0 28814 7 1 2 63345 89203
0 28815 7 1 2 96997 28814
0 28816 7 1 2 28813 28815
0 28817 5 1 1 28816
0 28818 7 1 2 28796 28817
0 28819 5 1 1 28818
0 28820 7 1 2 93115 28819
0 28821 5 1 1 28820
0 28822 7 3 2 74279 86570
0 28823 7 1 2 66498 76650
0 28824 7 1 2 76023 28823
0 28825 7 1 2 97219 28824
0 28826 7 1 2 84385 96733
0 28827 7 1 2 28825 28826
0 28828 5 1 1 28827
0 28829 7 1 2 28821 28828
0 28830 5 1 1 28829
0 28831 7 1 2 63170 28830
0 28832 5 1 1 28831
0 28833 7 3 2 82377 75776
0 28834 7 1 2 96547 97222
0 28835 5 1 1 28834
0 28836 7 3 2 72166 79181
0 28837 7 1 2 89913 96929
0 28838 7 1 2 97225 28837
0 28839 5 1 1 28838
0 28840 7 1 2 28835 28839
0 28841 5 1 1 28840
0 28842 7 1 2 65771 28841
0 28843 5 1 1 28842
0 28844 7 3 2 65998 82783
0 28845 7 1 2 95051 96574
0 28846 7 1 2 97228 28845
0 28847 5 1 1 28846
0 28848 7 1 2 28843 28847
0 28849 5 1 1 28848
0 28850 7 1 2 61603 28849
0 28851 5 1 1 28850
0 28852 7 1 2 83985 89809
0 28853 5 1 1 28852
0 28854 7 1 2 69001 89432
0 28855 5 1 1 28854
0 28856 7 1 2 28853 28855
0 28857 5 1 1 28856
0 28858 7 1 2 74326 85644
0 28859 7 1 2 87924 28858
0 28860 7 1 2 28857 28859
0 28861 5 1 1 28860
0 28862 7 1 2 28851 28861
0 28863 5 1 1 28862
0 28864 7 1 2 67698 28863
0 28865 5 1 1 28864
0 28866 7 1 2 96779 97216
0 28867 5 1 1 28866
0 28868 7 1 2 28865 28867
0 28869 5 1 1 28868
0 28870 7 1 2 80807 94197
0 28871 7 1 2 28869 28870
0 28872 5 1 1 28871
0 28873 7 1 2 28832 28872
0 28874 5 1 1 28873
0 28875 7 1 2 65168 28874
0 28876 5 1 1 28875
0 28877 7 1 2 86833 97105
0 28878 5 1 1 28877
0 28879 7 1 2 78706 96431
0 28880 5 1 1 28879
0 28881 7 1 2 28878 28880
0 28882 5 1 1 28881
0 28883 7 1 2 86962 28882
0 28884 5 1 1 28883
0 28885 7 3 2 79130 93116
0 28886 7 1 2 83002 97231
0 28887 5 1 1 28886
0 28888 7 2 2 81656 96460
0 28889 7 1 2 91228 97234
0 28890 5 1 1 28889
0 28891 7 1 2 28887 28890
0 28892 5 1 1 28891
0 28893 7 1 2 63972 28892
0 28894 5 1 1 28893
0 28895 7 1 2 28884 28894
0 28896 7 1 2 78378 97113
0 28897 5 1 1 28896
0 28898 7 1 2 82170 92796
0 28899 7 1 2 88961 28898
0 28900 5 1 1 28899
0 28901 7 1 2 28897 28900
0 28902 5 1 1 28901
0 28903 7 1 2 81928 28902
0 28904 5 1 1 28903
0 28905 7 1 2 64354 80789
0 28906 7 1 2 82721 28905
0 28907 5 1 1 28906
0 28908 7 3 2 64740 86834
0 28909 7 1 2 96134 97236
0 28910 5 1 1 28909
0 28911 7 1 2 28907 28910
0 28912 5 1 1 28911
0 28913 7 1 2 87251 28912
0 28914 5 1 1 28913
0 28915 7 1 2 28904 28914
0 28916 7 1 2 28895 28915
0 28917 5 1 1 28916
0 28918 7 1 2 65999 28917
0 28919 5 1 1 28918
0 28920 7 1 2 88190 86835
0 28921 5 1 1 28920
0 28922 7 1 2 92098 94659
0 28923 5 1 1 28922
0 28924 7 1 2 28921 28923
0 28925 5 1 1 28924
0 28926 7 1 2 93117 28925
0 28927 5 1 1 28926
0 28928 7 1 2 96597 97237
0 28929 5 1 1 28928
0 28930 7 1 2 28927 28929
0 28931 5 1 1 28930
0 28932 7 1 2 81998 28931
0 28933 5 1 1 28932
0 28934 7 1 2 80938 91847
0 28935 5 1 1 28934
0 28936 7 1 2 97123 28935
0 28937 5 5 1 28936
0 28938 7 1 2 63171 86836
0 28939 7 1 2 97239 28938
0 28940 5 1 1 28939
0 28941 7 2 2 82989 87925
0 28942 7 1 2 80790 78760
0 28943 7 1 2 97244 28942
0 28944 5 1 1 28943
0 28945 7 1 2 28940 28944
0 28946 5 1 1 28945
0 28947 7 1 2 78844 28946
0 28948 5 1 1 28947
0 28949 7 1 2 28933 28948
0 28950 7 1 2 28919 28949
0 28951 5 1 1 28950
0 28952 7 1 2 69002 28951
0 28953 5 1 1 28952
0 28954 7 1 2 85544 91848
0 28955 5 1 1 28954
0 28956 7 1 2 27234 28955
0 28957 5 1 1 28956
0 28958 7 1 2 66499 28957
0 28959 5 1 1 28958
0 28960 7 1 2 87126 97121
0 28961 5 1 1 28960
0 28962 7 1 2 28959 28961
0 28963 5 1 1 28962
0 28964 7 1 2 87252 28963
0 28965 5 1 1 28964
0 28966 7 2 2 78477 92797
0 28967 7 1 2 90535 97246
0 28968 7 1 2 85567 28967
0 28969 5 1 1 28968
0 28970 7 1 2 67471 83196
0 28971 7 1 2 97189 28970
0 28972 5 1 1 28971
0 28973 7 1 2 28969 28972
0 28974 7 1 2 28965 28973
0 28975 5 1 1 28974
0 28976 7 1 2 64138 28975
0 28977 5 1 1 28976
0 28978 7 1 2 82171 91541
0 28979 7 1 2 95911 28978
0 28980 5 1 1 28979
0 28981 7 1 2 28977 28980
0 28982 5 1 1 28981
0 28983 7 1 2 70931 28982
0 28984 5 1 1 28983
0 28985 7 1 2 82829 96481
0 28986 5 1 1 28985
0 28987 7 1 2 83323 96469
0 28988 5 1 1 28987
0 28989 7 2 2 96720 28988
0 28990 7 1 2 28986 97248
0 28991 5 1 1 28990
0 28992 7 1 2 86837 28991
0 28993 5 1 1 28992
0 28994 7 2 2 72701 92361
0 28995 5 1 1 97250
0 28996 7 1 2 97235 97251
0 28997 5 1 1 28996
0 28998 7 1 2 28993 28997
0 28999 5 1 1 28998
0 29000 7 1 2 66000 28999
0 29001 5 1 1 29000
0 29002 7 1 2 28984 29001
0 29003 7 1 2 28953 29002
0 29004 5 1 1 29003
0 29005 7 1 2 65437 29004
0 29006 5 1 1 29005
0 29007 7 1 2 76738 97086
0 29008 5 1 1 29007
0 29009 7 1 2 73555 97124
0 29010 5 1 1 29009
0 29011 7 1 2 97128 29010
0 29012 5 1 1 29011
0 29013 7 1 2 87359 73579
0 29014 7 1 2 97106 29013
0 29015 5 1 1 29014
0 29016 7 1 2 88875 96548
0 29017 5 1 1 29016
0 29018 7 1 2 29015 29017
0 29019 7 1 2 29012 29018
0 29020 5 1 1 29019
0 29021 7 1 2 71242 29020
0 29022 5 1 1 29021
0 29023 7 1 2 29008 29022
0 29024 5 1 1 29023
0 29025 7 1 2 69003 29024
0 29026 5 1 1 29025
0 29027 7 1 2 78845 96467
0 29028 5 1 1 29027
0 29029 7 1 2 97249 29028
0 29030 5 1 1 29029
0 29031 7 1 2 84731 29030
0 29032 5 1 1 29031
0 29033 7 1 2 29026 29032
0 29034 5 1 1 29033
0 29035 7 1 2 72453 29034
0 29036 5 1 1 29035
0 29037 7 1 2 29006 29036
0 29038 5 1 1 29037
0 29039 7 1 2 65169 29038
0 29040 5 1 1 29039
0 29041 7 1 2 86963 87537
0 29042 5 1 1 29041
0 29043 7 1 2 64139 95760
0 29044 5 1 1 29043
0 29045 7 1 2 29042 29044
0 29046 5 1 1 29045
0 29047 7 1 2 63172 71338
0 29048 7 1 2 29046 29047
0 29049 5 1 1 29048
0 29050 7 2 2 78761 84560
0 29051 7 1 2 82784 78516
0 29052 7 1 2 97252 29051
0 29053 5 1 1 29052
0 29054 7 1 2 29049 29053
0 29055 5 1 1 29054
0 29056 7 1 2 93118 29055
0 29057 5 1 1 29056
0 29058 7 1 2 71061 93045
0 29059 5 1 1 29058
0 29060 7 1 2 77006 91849
0 29061 5 1 1 29060
0 29062 7 1 2 29059 29061
0 29063 5 1 1 29062
0 29064 7 1 2 78770 29063
0 29065 5 1 1 29064
0 29066 7 1 2 73705 96182
0 29067 5 1 1 29066
0 29068 7 1 2 29065 29067
0 29069 5 1 1 29068
0 29070 7 1 2 66500 29069
0 29071 5 1 1 29070
0 29072 7 1 2 88856 78517
0 29073 7 1 2 97232 29072
0 29074 5 1 1 29073
0 29075 7 1 2 29071 29074
0 29076 5 1 1 29075
0 29077 7 1 2 80012 29076
0 29078 5 1 1 29077
0 29079 7 1 2 29057 29078
0 29080 5 1 1 29079
0 29081 7 1 2 70932 29080
0 29082 5 1 1 29081
0 29083 7 1 2 77011 96392
0 29084 5 1 1 29083
0 29085 7 1 2 96579 29084
0 29086 5 1 1 29085
0 29087 7 1 2 64741 75654
0 29088 7 1 2 29086 29087
0 29089 5 1 1 29088
0 29090 7 1 2 29082 29089
0 29091 5 1 1 29090
0 29092 7 1 2 79607 29091
0 29093 5 1 1 29092
0 29094 7 1 2 29040 29093
0 29095 5 1 1 29094
0 29096 7 1 2 63346 29095
0 29097 5 1 1 29096
0 29098 7 1 2 79182 96589
0 29099 5 1 1 29098
0 29100 7 3 2 77203 92798
0 29101 7 1 2 80212 79131
0 29102 7 1 2 97254 29101
0 29103 5 1 1 29102
0 29104 7 1 2 29099 29103
0 29105 5 2 1 29104
0 29106 7 1 2 78330 97257
0 29107 5 1 1 29106
0 29108 7 1 2 86964 73556
0 29109 5 1 1 29108
0 29110 7 1 2 84884 81929
0 29111 5 1 1 29110
0 29112 7 1 2 29109 29111
0 29113 5 1 1 29112
0 29114 7 1 2 68019 29113
0 29115 5 1 1 29114
0 29116 7 1 2 70714 95779
0 29117 5 1 1 29116
0 29118 7 1 2 29115 29117
0 29119 5 1 1 29118
0 29120 7 1 2 96699 29119
0 29121 5 1 1 29120
0 29122 7 1 2 29107 29121
0 29123 5 1 1 29122
0 29124 7 1 2 73328 29123
0 29125 5 1 1 29124
0 29126 7 1 2 61880 84576
0 29127 7 1 2 96549 29126
0 29128 5 1 1 29127
0 29129 7 1 2 64140 85555
0 29130 7 1 2 96504 29129
0 29131 5 1 1 29130
0 29132 7 1 2 29128 29131
0 29133 5 1 1 29132
0 29134 7 1 2 70933 29133
0 29135 5 1 1 29134
0 29136 7 1 2 89284 77683
0 29137 7 1 2 96243 29136
0 29138 5 1 1 29137
0 29139 7 1 2 29135 29138
0 29140 5 1 1 29139
0 29141 7 1 2 76163 29140
0 29142 5 1 1 29141
0 29143 7 1 2 64141 97258
0 29144 5 1 1 29143
0 29145 7 1 2 93213 96500
0 29146 5 1 1 29145
0 29147 7 1 2 29144 29146
0 29148 5 1 1 29147
0 29149 7 1 2 92427 29148
0 29150 5 1 1 29149
0 29151 7 1 2 29142 29150
0 29152 7 1 2 29125 29151
0 29153 5 1 1 29152
0 29154 7 1 2 96479 29153
0 29155 5 1 1 29154
0 29156 7 1 2 29097 29155
0 29157 5 1 1 29156
0 29158 7 1 2 73024 29157
0 29159 5 1 1 29158
0 29160 7 3 2 68853 94274
0 29161 7 1 2 87208 86183
0 29162 7 1 2 97259 29161
0 29163 5 1 1 29162
0 29164 7 2 2 64142 76326
0 29165 5 2 1 97262
0 29166 7 1 2 84027 97264
0 29167 5 1 1 29166
0 29168 7 2 2 73329 85189
0 29169 7 1 2 71841 97266
0 29170 7 1 2 29167 29169
0 29171 5 1 1 29170
0 29172 7 1 2 29163 29171
0 29173 5 1 1 29172
0 29174 7 1 2 70090 29173
0 29175 5 1 1 29174
0 29176 7 3 2 70715 72702
0 29177 7 1 2 84819 80861
0 29178 7 1 2 97268 29177
0 29179 7 1 2 93983 29178
0 29180 5 1 1 29179
0 29181 7 1 2 29175 29180
0 29182 5 1 1 29181
0 29183 7 1 2 61881 29182
0 29184 5 1 1 29183
0 29185 7 1 2 70091 84016
0 29186 7 1 2 92135 29185
0 29187 7 1 2 92735 29186
0 29188 5 1 1 29187
0 29189 7 1 2 29184 29188
0 29190 5 1 1 29189
0 29191 7 1 2 76164 29190
0 29192 5 1 1 29191
0 29193 7 2 2 71243 74543
0 29194 5 2 1 97271
0 29195 7 1 2 76049 97272
0 29196 5 1 1 29195
0 29197 7 1 2 75959 91962
0 29198 5 1 1 29197
0 29199 7 1 2 29196 29198
0 29200 5 1 1 29199
0 29201 7 1 2 91107 29200
0 29202 5 1 1 29201
0 29203 7 1 2 92254 92528
0 29204 5 1 1 29203
0 29205 7 3 2 61604 72703
0 29206 7 1 2 73853 95803
0 29207 7 1 2 97275 29206
0 29208 5 1 1 29207
0 29209 7 1 2 29204 29208
0 29210 5 1 1 29209
0 29211 7 1 2 67266 29210
0 29212 5 1 1 29211
0 29213 7 2 2 78699 80729
0 29214 7 1 2 74624 73689
0 29215 7 1 2 97278 29214
0 29216 5 1 1 29215
0 29217 7 1 2 29212 29216
0 29218 7 1 2 29202 29217
0 29219 5 1 1 29218
0 29220 7 1 2 88650 79683
0 29221 7 1 2 29219 29220
0 29222 5 1 1 29221
0 29223 7 1 2 29192 29222
0 29224 5 1 1 29223
0 29225 7 1 2 69579 29224
0 29226 5 1 1 29225
0 29227 7 1 2 73070 86077
0 29228 5 1 1 29227
0 29229 7 1 2 69004 90376
0 29230 7 1 2 91733 29229
0 29231 5 1 1 29230
0 29232 7 1 2 29228 29231
0 29233 5 1 1 29232
0 29234 7 1 2 71244 29233
0 29235 5 1 1 29234
0 29236 7 1 2 88088 97130
0 29237 5 1 1 29236
0 29238 7 1 2 67699 29237
0 29239 5 1 1 29238
0 29240 7 3 2 80533 92371
0 29241 5 3 1 97280
0 29242 7 1 2 65438 97283
0 29243 7 1 2 29239 29242
0 29244 5 1 1 29243
0 29245 7 1 2 62849 79656
0 29246 5 1 1 29245
0 29247 7 1 2 91337 29246
0 29248 5 1 1 29247
0 29249 7 1 2 65772 29248
0 29250 5 1 1 29249
0 29251 7 1 2 70361 94572
0 29252 7 1 2 29250 29251
0 29253 5 1 1 29252
0 29254 7 1 2 68662 29253
0 29255 7 1 2 29244 29254
0 29256 5 1 1 29255
0 29257 7 1 2 29235 29256
0 29258 5 1 1 29257
0 29259 7 1 2 65170 29258
0 29260 5 1 1 29259
0 29261 7 6 2 67267 85713
0 29262 7 1 2 81027 97286
0 29263 7 1 2 97260 29262
0 29264 5 1 1 29263
0 29265 7 1 2 29260 29264
0 29266 5 1 1 29265
0 29267 7 3 2 78887 82249
0 29268 7 1 2 61882 97292
0 29269 7 1 2 29266 29268
0 29270 5 1 1 29269
0 29271 7 1 2 29226 29270
0 29272 5 1 1 29271
0 29273 7 1 2 69815 29272
0 29274 5 1 1 29273
0 29275 7 2 2 61605 88973
0 29276 7 1 2 79865 92160
0 29277 7 1 2 85407 29276
0 29278 5 1 1 29277
0 29279 7 2 2 65439 87066
0 29280 7 1 2 89880 97297
0 29281 7 1 2 86703 29280
0 29282 5 1 1 29281
0 29283 7 1 2 29278 29282
0 29284 5 1 1 29283
0 29285 7 1 2 63808 29284
0 29286 5 1 1 29285
0 29287 7 1 2 71967 96706
0 29288 5 1 1 29287
0 29289 7 1 2 78248 94275
0 29290 5 1 1 29289
0 29291 7 1 2 29288 29290
0 29292 5 1 1 29291
0 29293 7 1 2 91595 29292
0 29294 5 1 1 29293
0 29295 7 1 2 29286 29294
0 29296 5 1 1 29295
0 29297 7 1 2 67700 29296
0 29298 5 1 1 29297
0 29299 7 1 2 70092 74544
0 29300 5 1 1 29299
0 29301 7 1 2 11389 29300
0 29302 5 1 1 29301
0 29303 7 1 2 62420 29302
0 29304 5 1 1 29303
0 29305 7 2 2 70362 95575
0 29306 5 1 1 97299
0 29307 7 1 2 70093 97300
0 29308 5 1 1 29307
0 29309 7 1 2 29304 29308
0 29310 5 1 1 29309
0 29311 7 1 2 86198 96851
0 29312 7 1 2 29310 29311
0 29313 5 1 1 29312
0 29314 7 1 2 29298 29313
0 29315 5 1 1 29314
0 29316 7 1 2 63173 29315
0 29317 5 1 1 29316
0 29318 7 1 2 69005 87112
0 29319 7 1 2 88612 29318
0 29320 7 2 2 70094 77818
0 29321 7 1 2 79285 97301
0 29322 7 1 2 29319 29321
0 29323 5 1 1 29322
0 29324 7 1 2 29317 29323
0 29325 5 1 1 29324
0 29326 7 1 2 97295 29325
0 29327 5 1 1 29326
0 29328 7 1 2 29274 29327
0 29329 5 1 1 29328
0 29330 7 1 2 93119 29329
0 29331 5 1 1 29330
0 29332 7 1 2 29159 29331
0 29333 5 1 1 29332
0 29334 7 1 2 75155 29333
0 29335 5 1 1 29334
0 29336 7 1 2 28876 29335
0 29337 7 1 2 28729 29336
0 29338 7 1 2 28248 29337
0 29339 5 1 1 29338
0 29340 7 25 2 69096 92640
0 29341 7 1 2 29339 97303
0 29342 5 1 1 29341
0 29343 7 1 2 27805 29342
0 29344 7 1 2 23314 29343
0 29345 5 1 1 29344
0 29346 7 1 2 93770 29345
0 29347 5 1 1 29346
0 29348 7 3 2 77973 87120
0 29349 7 1 2 78280 97328
0 29350 5 1 1 29349
0 29351 7 2 2 79132 86838
0 29352 7 1 2 61883 97331
0 29353 5 1 1 29352
0 29354 7 1 2 29350 29353
0 29355 5 1 1 29354
0 29356 7 1 2 92165 29355
0 29357 5 1 1 29356
0 29358 7 3 2 79081 82896
0 29359 7 6 2 66744 62953
0 29360 7 1 2 64355 97336
0 29361 7 1 2 97333 29360
0 29362 5 1 1 29361
0 29363 7 1 2 29357 29362
0 29364 5 1 1 29363
0 29365 7 1 2 69006 29364
0 29366 5 1 1 29365
0 29367 7 1 2 75707 92166
0 29368 7 1 2 97332 29367
0 29369 5 1 1 29368
0 29370 7 1 2 29366 29369
0 29371 5 1 1 29370
0 29372 7 1 2 66001 29371
0 29373 5 1 1 29372
0 29374 7 1 2 62850 71533
0 29375 5 2 1 29374
0 29376 7 1 2 75745 96663
0 29377 5 1 1 29376
0 29378 7 1 2 97342 29377
0 29379 5 1 1 29378
0 29380 7 1 2 70934 29379
0 29381 5 1 1 29380
0 29382 7 1 2 71684 29381
0 29383 5 1 1 29382
0 29384 7 1 2 83349 29383
0 29385 5 1 1 29384
0 29386 7 1 2 79102 72356
0 29387 5 1 1 29386
0 29388 7 1 2 29385 29387
0 29389 5 1 1 29388
0 29390 7 1 2 92167 29389
0 29391 5 1 1 29390
0 29392 7 1 2 29373 29391
0 29393 5 1 1 29392
0 29394 7 1 2 61606 29393
0 29395 5 1 1 29394
0 29396 7 1 2 77788 95142
0 29397 7 5 2 67701 67776
0 29398 7 5 2 67472 97344
0 29399 7 1 2 95481 97349
0 29400 7 1 2 29396 29399
0 29401 5 1 1 29400
0 29402 7 1 2 29395 29401
0 29403 5 1 1 29402
0 29404 7 1 2 64528 29403
0 29405 5 1 1 29404
0 29406 7 1 2 87079 93588
0 29407 5 1 1 29406
0 29408 7 6 2 67777 68854
0 29409 7 3 2 87926 97354
0 29410 7 1 2 73146 97360
0 29411 5 1 1 29410
0 29412 7 1 2 29407 29411
0 29413 5 1 1 29412
0 29414 7 1 2 83884 29413
0 29415 5 1 1 29414
0 29416 7 1 2 63174 29415
0 29417 7 1 2 29405 29416
0 29418 5 1 1 29417
0 29419 7 2 2 64950 95667
0 29420 7 7 2 62583 62954
0 29421 7 1 2 96918 97365
0 29422 7 1 2 97363 29421
0 29423 5 1 1 29422
0 29424 7 1 2 83350 93669
0 29425 5 1 1 29424
0 29426 7 1 2 66745 78029
0 29427 7 1 2 81219 29426
0 29428 5 1 1 29427
0 29429 7 1 2 29425 29428
0 29430 5 1 1 29429
0 29431 7 1 2 85357 92168
0 29432 7 1 2 29430 29431
0 29433 5 1 1 29432
0 29434 7 1 2 29423 29433
0 29435 5 1 1 29434
0 29436 7 1 2 65773 29435
0 29437 5 1 1 29436
0 29438 7 2 2 89906 95242
0 29439 5 1 1 97372
0 29440 7 1 2 93589 97373
0 29441 5 1 1 29440
0 29442 7 1 2 89285 87825
0 29443 7 1 2 97355 29442
0 29444 7 1 2 82400 29443
0 29445 5 1 1 29444
0 29446 7 1 2 29441 29445
0 29447 5 1 1 29446
0 29448 7 1 2 67702 29447
0 29449 5 1 1 29448
0 29450 7 2 2 79082 93590
0 29451 7 1 2 75594 97374
0 29452 7 1 2 97108 29451
0 29453 5 1 1 29452
0 29454 7 1 2 29449 29453
0 29455 7 1 2 29437 29454
0 29456 5 1 1 29455
0 29457 7 1 2 82115 29456
0 29458 5 1 1 29457
0 29459 7 1 2 77833 97356
0 29460 7 1 2 96074 96351
0 29461 7 1 2 29459 29460
0 29462 5 1 1 29461
0 29463 7 1 2 68020 29462
0 29464 7 1 2 29458 29463
0 29465 5 1 1 29464
0 29466 7 1 2 90656 29465
0 29467 7 1 2 29418 29466
0 29468 5 1 1 29467
0 29469 7 7 2 64356 64951
0 29470 7 3 2 66002 82897
0 29471 5 1 1 97383
0 29472 7 3 2 83812 91320
0 29473 7 1 2 97384 97386
0 29474 5 1 1 29473
0 29475 7 1 2 84910 86847
0 29476 5 1 1 29475
0 29477 7 1 2 82327 29476
0 29478 5 1 1 29477
0 29479 7 1 2 29474 29478
0 29480 5 1 1 29479
0 29481 7 1 2 69580 29480
0 29482 5 1 1 29481
0 29483 7 3 2 64143 76092
0 29484 7 2 2 79445 97389
0 29485 7 1 2 85605 97392
0 29486 5 1 1 29485
0 29487 7 1 2 29482 29486
0 29488 5 1 1 29487
0 29489 7 2 2 97376 29488
0 29490 7 3 2 66746 63000
0 29491 7 3 2 61349 67778
0 29492 7 1 2 97396 97399
0 29493 7 1 2 97394 29492
0 29494 5 1 1 29493
0 29495 7 1 2 29468 29494
0 29496 5 2 1 29495
0 29497 7 1 2 66100 97402
0 29498 5 1 1 29497
0 29499 7 2 2 66747 67779
0 29500 7 4 2 92980 97404
0 29501 5 1 1 97406
0 29502 7 1 2 97407 97395
0 29503 5 1 1 29502
0 29504 7 1 2 29498 29503
0 29505 5 1 1 29504
0 29506 7 1 2 65440 29505
0 29507 5 1 1 29506
0 29508 7 1 2 73463 88839
0 29509 5 1 1 29508
0 29510 7 1 2 93315 29509
0 29511 5 1 1 29510
0 29512 7 1 2 69007 29511
0 29513 5 1 1 29512
0 29514 7 1 2 89858 95397
0 29515 5 1 1 29514
0 29516 7 1 2 29513 29515
0 29517 5 2 1 29516
0 29518 7 2 2 80296 78268
0 29519 5 1 1 97412
0 29520 7 13 2 64357 65774
0 29521 7 2 2 97413 97414
0 29522 7 1 2 92470 97427
0 29523 7 1 2 97410 29522
0 29524 5 1 1 29523
0 29525 7 1 2 29507 29524
0 29526 5 1 1 29525
0 29527 7 1 2 66969 29526
0 29528 5 1 1 29527
0 29529 7 3 2 61884 89760
0 29530 5 1 1 97429
0 29531 7 1 2 7618 29530
0 29532 5 1 1 29531
0 29533 7 1 2 74200 90960
0 29534 7 1 2 96191 29533
0 29535 7 1 2 29532 29534
0 29536 7 1 2 92471 29535
0 29537 5 1 1 29536
0 29538 7 1 2 29528 29537
0 29539 5 1 1 29538
0 29540 7 1 2 69097 29539
0 29541 5 1 1 29540
0 29542 7 6 2 69209 70363
0 29543 7 2 2 70935 75305
0 29544 7 1 2 97432 97438
0 29545 7 2 2 91017 29544
0 29546 7 1 2 77698 97440
0 29547 5 1 1 29546
0 29548 7 1 2 61885 84276
0 29549 7 1 2 88175 29548
0 29550 7 6 2 65775 76775
0 29551 7 1 2 96702 97442
0 29552 7 1 2 29549 29551
0 29553 5 1 1 29552
0 29554 7 1 2 29547 29553
0 29555 5 1 1 29554
0 29556 7 4 2 64255 64742
0 29557 7 1 2 82328 97448
0 29558 7 1 2 29555 29557
0 29559 5 1 1 29558
0 29560 7 1 2 29541 29559
0 29561 5 1 1 29560
0 29562 7 1 2 63347 29561
0 29563 5 1 1 29562
0 29564 7 3 2 63973 87831
0 29565 7 9 2 66215 67780
0 29566 7 5 2 67849 97455
0 29567 7 2 2 81870 97464
0 29568 7 1 2 97452 97469
0 29569 5 1 1 29568
0 29570 7 2 2 18143 29569
0 29571 5 1 1 97471
0 29572 7 1 2 86915 73864
0 29573 5 2 1 29572
0 29574 7 2 2 76249 75531
0 29575 5 1 1 97475
0 29576 7 1 2 84789 97476
0 29577 5 1 1 29576
0 29578 7 1 2 97473 29577
0 29579 5 1 1 29578
0 29580 7 1 2 83899 29579
0 29581 5 1 1 29580
0 29582 7 1 2 75420 83227
0 29583 7 1 2 88160 29582
0 29584 5 1 1 29583
0 29585 7 1 2 29581 29584
0 29586 5 1 1 29585
0 29587 7 1 2 29571 29586
0 29588 5 1 1 29587
0 29589 7 4 2 67781 93017
0 29590 5 1 1 97477
0 29591 7 1 2 67703 89433
0 29592 5 1 1 29591
0 29593 7 1 2 88930 86877
0 29594 5 1 1 29593
0 29595 7 1 2 29592 29594
0 29596 5 1 1 29595
0 29597 7 1 2 97478 29596
0 29598 5 1 1 29597
0 29599 7 1 2 97337 97377
0 29600 7 1 2 93246 29599
0 29601 5 1 1 29600
0 29602 7 1 2 29598 29601
0 29603 5 1 1 29602
0 29604 7 1 2 67473 29603
0 29605 5 1 1 29604
0 29606 7 2 2 64358 84229
0 29607 7 2 2 64743 81211
0 29608 7 1 2 68855 97338
0 29609 7 1 2 97483 29608
0 29610 7 1 2 97481 29609
0 29611 5 1 1 29610
0 29612 7 1 2 29605 29611
0 29613 5 1 1 29612
0 29614 7 1 2 70364 29613
0 29615 5 1 1 29614
0 29616 7 1 2 89290 92169
0 29617 7 1 2 88161 29616
0 29618 5 1 1 29617
0 29619 7 1 2 29615 29618
0 29620 5 1 1 29619
0 29621 7 1 2 65776 29620
0 29622 5 1 1 29621
0 29623 7 1 2 80051 89403
0 29624 5 1 1 29623
0 29625 7 3 2 86283 87165
0 29626 5 1 1 97485
0 29627 7 1 2 29624 29626
0 29628 5 1 1 29627
0 29629 7 1 2 74732 93591
0 29630 7 1 2 29628 29629
0 29631 5 1 1 29630
0 29632 7 1 2 29622 29631
0 29633 5 1 1 29632
0 29634 7 1 2 90657 29633
0 29635 5 1 1 29634
0 29636 7 5 2 69581 76776
0 29637 7 1 2 89219 97488
0 29638 5 2 1 29637
0 29639 7 1 2 83188 97486
0 29640 5 1 1 29639
0 29641 7 1 2 97493 29640
0 29642 5 1 1 29641
0 29643 7 1 2 66003 29642
0 29644 5 1 1 29643
0 29645 7 1 2 74733 97487
0 29646 5 1 1 29645
0 29647 7 1 2 29644 29646
0 29648 5 1 1 29647
0 29649 7 2 2 64359 29648
0 29650 7 1 2 90642 97495
0 29651 5 1 1 29650
0 29652 7 1 2 29635 29651
0 29653 5 1 1 29652
0 29654 7 1 2 66101 29653
0 29655 5 1 1 29654
0 29656 7 1 2 92458 97496
0 29657 5 1 1 29656
0 29658 7 1 2 29655 29657
0 29659 5 1 1 29658
0 29660 7 1 2 69008 29659
0 29661 5 1 1 29660
0 29662 7 2 2 87930 97470
0 29663 5 1 1 97497
0 29664 7 8 2 61886 82785
0 29665 7 2 2 73650 82277
0 29666 7 1 2 97499 97507
0 29667 5 1 1 29666
0 29668 7 2 2 76849 88121
0 29669 7 1 2 86307 73699
0 29670 7 1 2 97509 29669
0 29671 5 1 1 29670
0 29672 7 1 2 29667 29671
0 29673 5 1 1 29672
0 29674 7 1 2 97498 29673
0 29675 5 1 1 29674
0 29676 7 1 2 29661 29675
0 29677 5 1 1 29676
0 29678 7 1 2 84790 29677
0 29679 5 1 1 29678
0 29680 7 1 2 29588 29679
0 29681 5 1 1 29680
0 29682 7 1 2 69098 29681
0 29683 5 1 1 29682
0 29684 7 2 2 64744 94631
0 29685 7 1 2 85190 97441
0 29686 5 1 1 29685
0 29687 7 1 2 62117 96289
0 29688 5 4 1 29687
0 29689 7 1 2 66970 72167
0 29690 5 1 1 29689
0 29691 7 1 2 62851 29690
0 29692 5 1 1 29691
0 29693 7 4 2 66102 90596
0 29694 5 1 1 97517
0 29695 7 1 2 16977 29694
0 29696 5 2 1 29695
0 29697 7 7 2 62955 69210
0 29698 7 1 2 97521 97523
0 29699 7 1 2 29692 29698
0 29700 7 1 2 97513 29699
0 29701 5 1 1 29700
0 29702 7 1 2 66971 92170
0 29703 5 2 1 29702
0 29704 7 2 2 62956 87857
0 29705 5 1 1 97532
0 29706 7 1 2 93613 29590
0 29707 5 2 1 29706
0 29708 7 1 2 67474 97534
0 29709 5 1 1 29708
0 29710 7 1 2 29705 29709
0 29711 5 1 1 29710
0 29712 7 1 2 86209 29711
0 29713 5 1 1 29712
0 29714 7 1 2 97530 29713
0 29715 5 1 1 29714
0 29716 7 1 2 61267 90597
0 29717 7 1 2 84319 29716
0 29718 7 1 2 29715 29717
0 29719 5 1 1 29718
0 29720 7 1 2 29701 29719
0 29721 5 1 1 29720
0 29722 7 1 2 86571 29721
0 29723 5 1 1 29722
0 29724 7 1 2 29686 29723
0 29725 5 1 1 29724
0 29726 7 1 2 64952 29725
0 29727 5 1 1 29726
0 29728 7 1 2 89914 96069
0 29729 7 1 2 91069 29728
0 29730 5 1 1 29729
0 29731 7 1 2 29727 29730
0 29732 5 1 1 29731
0 29733 7 1 2 66748 29732
0 29734 5 1 1 29733
0 29735 7 1 2 91328 96448
0 29736 7 1 2 75889 29735
0 29737 7 1 2 91018 29736
0 29738 5 1 1 29737
0 29739 7 1 2 29734 29738
0 29740 5 1 1 29739
0 29741 7 1 2 97511 29740
0 29742 5 1 1 29741
0 29743 7 1 2 29683 29742
0 29744 5 1 1 29743
0 29745 7 1 2 76165 29744
0 29746 5 1 1 29745
0 29747 7 1 2 66103 92799
0 29748 7 1 2 95662 29747
0 29749 5 2 1 29748
0 29750 7 4 2 61268 87938
0 29751 5 4 1 97538
0 29752 7 3 2 81871 93018
0 29753 5 1 1 97546
0 29754 7 1 2 97542 29753
0 29755 5 4 1 29754
0 29756 7 2 2 66004 97549
0 29757 5 1 1 97553
0 29758 7 1 2 82329 97554
0 29759 5 1 1 29758
0 29760 7 1 2 97536 29759
0 29761 5 1 1 29760
0 29762 7 1 2 69009 29761
0 29763 5 1 1 29762
0 29764 7 2 2 80651 87679
0 29765 7 3 2 69211 66005
0 29766 7 1 2 81535 97557
0 29767 7 1 2 97555 29766
0 29768 5 1 1 29767
0 29769 7 1 2 29763 29768
0 29770 5 1 1 29769
0 29771 7 1 2 67704 29770
0 29772 5 1 1 29771
0 29773 7 2 2 86409 92800
0 29774 7 1 2 97560 97556
0 29775 5 1 1 29774
0 29776 7 1 2 29772 29775
0 29777 5 1 1 29776
0 29778 7 8 2 69099 91857
0 29779 7 8 2 66216 66972
0 29780 7 1 2 82864 97570
0 29781 7 1 2 97562 29780
0 29782 7 1 2 29777 29781
0 29783 5 1 1 29782
0 29784 7 2 2 77029 88668
0 29785 7 15 2 62852 67782
0 29786 7 2 2 61607 97580
0 29787 7 3 2 61269 90658
0 29788 7 1 2 95192 97597
0 29789 7 1 2 97595 29788
0 29790 5 1 1 29789
0 29791 7 7 2 66501 62957
0 29792 7 1 2 92564 97600
0 29793 7 1 2 94611 29792
0 29794 5 1 1 29793
0 29795 7 1 2 29790 29794
0 29796 5 1 1 29795
0 29797 7 1 2 97578 29796
0 29798 5 1 1 29797
0 29799 7 17 2 61270 93901
0 29800 5 1 1 97607
0 29801 7 1 2 82330 97608
0 29802 5 1 1 29801
0 29803 7 1 2 66104 92099
0 29804 7 1 2 95116 29803
0 29805 5 1 1 29804
0 29806 7 1 2 29802 29805
0 29807 5 1 1 29806
0 29808 7 1 2 97579 29807
0 29809 5 1 1 29808
0 29810 7 16 2 66105 69100
0 29811 7 2 2 82700 97624
0 29812 7 1 2 88917 80227
0 29813 7 1 2 88030 29812
0 29814 7 1 2 97640 29813
0 29815 7 1 2 86371 29814
0 29816 5 1 1 29815
0 29817 7 1 2 29809 29816
0 29818 5 1 1 29817
0 29819 7 1 2 90705 29818
0 29820 5 1 1 29819
0 29821 7 1 2 29798 29820
0 29822 7 1 2 29783 29821
0 29823 5 1 1 29822
0 29824 7 1 2 70365 29823
0 29825 5 1 1 29824
0 29826 7 14 2 62958 64256
0 29827 7 33 2 90598 97642
0 29828 5 2 1 97656
0 29829 7 3 2 85726 80981
0 29830 5 1 1 97691
0 29831 7 1 2 83832 87907
0 29832 5 1 1 29831
0 29833 7 1 2 29830 29832
0 29834 5 1 1 29833
0 29835 7 1 2 72168 29834
0 29836 5 1 1 29835
0 29837 7 1 2 81087 97514
0 29838 5 2 1 29837
0 29839 7 3 2 80982 82437
0 29840 5 1 1 97696
0 29841 7 1 2 27663 97697
0 29842 5 1 1 29841
0 29843 7 1 2 97694 29842
0 29844 7 1 2 29836 29843
0 29845 5 2 1 29844
0 29846 7 1 2 87787 97699
0 29847 5 1 1 29846
0 29848 7 2 2 83849 92321
0 29849 5 1 1 97701
0 29850 7 1 2 93316 29849
0 29851 5 1 1 29850
0 29852 7 1 2 66006 87767
0 29853 7 1 2 29851 29852
0 29854 5 1 1 29853
0 29855 7 1 2 29847 29854
0 29856 5 1 1 29855
0 29857 7 1 2 97657 29856
0 29858 5 1 1 29857
0 29859 7 1 2 85897 72423
0 29860 7 1 2 87871 94591
0 29861 7 1 2 29859 29860
0 29862 7 2 2 93009 29861
0 29863 7 1 2 82092 97571
0 29864 7 1 2 97703 29863
0 29865 5 1 1 29864
0 29866 7 1 2 29858 29865
0 29867 5 1 1 29866
0 29868 7 1 2 86572 29867
0 29869 5 1 1 29868
0 29870 7 29 2 61271 64257
0 29871 7 22 2 69212 97705
0 29872 7 2 2 86573 97734
0 29873 7 1 2 90706 97756
0 29874 7 1 2 97700 29873
0 29875 5 1 1 29874
0 29876 7 1 2 29869 29875
0 29877 7 1 2 29825 29876
0 29878 5 1 1 29877
0 29879 7 1 2 79183 29878
0 29880 5 1 1 29879
0 29881 7 1 2 84057 96005
0 29882 7 1 2 86372 29881
0 29883 5 1 1 29882
0 29884 7 1 2 73949 92404
0 29885 5 1 1 29884
0 29886 7 1 2 62584 29885
0 29887 5 1 1 29886
0 29888 7 2 2 91614 29887
0 29889 5 1 1 97758
0 29890 7 1 2 64144 29889
0 29891 5 1 1 29890
0 29892 7 1 2 75665 29891
0 29893 5 3 1 29892
0 29894 7 1 2 87672 87262
0 29895 7 1 2 97760 29894
0 29896 5 1 1 29895
0 29897 7 1 2 29883 29896
0 29898 5 1 1 29897
0 29899 7 1 2 69582 29898
0 29900 5 1 1 29899
0 29901 7 1 2 70936 76050
0 29902 5 1 1 29901
0 29903 7 1 2 2975 29902
0 29904 5 2 1 29903
0 29905 7 1 2 75492 86296
0 29906 7 1 2 97763 29905
0 29907 5 1 1 29906
0 29908 7 1 2 29900 29907
0 29909 5 1 1 29908
0 29910 7 1 2 92672 29909
0 29911 5 1 1 29910
0 29912 7 1 2 79393 87324
0 29913 5 2 1 29912
0 29914 7 1 2 83953 78331
0 29915 5 1 1 29914
0 29916 7 2 2 79446 89364
0 29917 5 1 1 97767
0 29918 7 1 2 70716 97768
0 29919 5 1 1 29918
0 29920 7 1 2 29915 29919
0 29921 5 1 1 29920
0 29922 7 1 2 62853 29921
0 29923 5 1 1 29922
0 29924 7 1 2 86308 90391
0 29925 5 1 1 29924
0 29926 7 1 2 29923 29925
0 29927 5 1 1 29926
0 29928 7 1 2 63974 29927
0 29929 5 1 1 29928
0 29930 7 1 2 97765 29929
0 29931 5 1 1 29930
0 29932 7 1 2 63175 29931
0 29933 5 1 1 29932
0 29934 7 2 2 66502 90862
0 29935 7 1 2 80426 86887
0 29936 7 1 2 97769 29935
0 29937 5 1 1 29936
0 29938 7 1 2 29933 29937
0 29939 5 1 1 29938
0 29940 7 1 2 62585 29939
0 29941 5 1 1 29940
0 29942 7 1 2 92100 93424
0 29943 7 1 2 96655 29942
0 29944 5 1 1 29943
0 29945 7 1 2 29941 29944
0 29946 5 1 1 29945
0 29947 7 8 2 66217 62118
0 29948 7 4 2 66106 97771
0 29949 7 1 2 69213 91858
0 29950 7 2 2 97779 29949
0 29951 7 1 2 66749 97783
0 29952 7 1 2 29946 29951
0 29953 5 1 1 29952
0 29954 7 1 2 29911 29953
0 29955 5 1 1 29954
0 29956 7 13 2 69101 70366
0 29957 7 1 2 81284 97785
0 29958 7 1 2 29955 29957
0 29959 5 1 1 29958
0 29960 7 1 2 29880 29959
0 29961 7 1 2 29746 29960
0 29962 7 1 2 29563 29961
0 29963 5 1 1 29962
0 29964 7 1 2 73025 29963
0 29965 5 1 1 29964
0 29966 7 2 2 79184 91019
0 29967 7 1 2 75960 84791
0 29968 5 2 1 29967
0 29969 7 1 2 62119 90931
0 29970 5 1 1 29969
0 29971 7 1 2 97800 29970
0 29972 5 6 1 29971
0 29973 7 1 2 73214 97802
0 29974 5 1 1 29973
0 29975 7 2 2 66973 74545
0 29976 5 1 1 97808
0 29977 7 1 2 76638 72870
0 29978 5 1 1 29977
0 29979 7 1 2 67268 29978
0 29980 5 1 1 29979
0 29981 7 1 2 29976 29980
0 29982 5 3 1 29981
0 29983 7 2 2 63348 97810
0 29984 7 1 2 85583 97813
0 29985 5 1 1 29984
0 29986 7 1 2 29974 29985
0 29987 5 1 1 29986
0 29988 7 1 2 81088 29987
0 29989 5 1 1 29988
0 29990 7 5 2 68186 70367
0 29991 7 2 2 79714 378
0 29992 5 4 1 97820
0 29993 7 2 2 73330 97822
0 29994 5 1 1 97826
0 29995 7 1 2 73464 74454
0 29996 5 1 1 29995
0 29997 7 1 2 29994 29996
0 29998 5 2 1 29997
0 29999 7 1 2 97815 97828
0 30000 5 1 1 29999
0 30001 7 1 2 66974 93993
0 30002 5 1 1 30001
0 30003 7 1 2 30000 30002
0 30004 5 1 1 30003
0 30005 7 1 2 70717 30004
0 30006 5 1 1 30005
0 30007 7 1 2 84792 94144
0 30008 5 1 1 30007
0 30009 7 1 2 30006 30008
0 30010 5 1 1 30009
0 30011 7 1 2 72064 30010
0 30012 5 1 1 30011
0 30013 7 1 2 94297 97814
0 30014 5 1 1 30013
0 30015 7 2 2 71339 97803
0 30016 7 1 2 72169 85085
0 30017 7 1 2 97830 30016
0 30018 5 1 1 30017
0 30019 7 1 2 88287 88669
0 30020 7 1 2 87576 30019
0 30021 7 1 2 77750 30020
0 30022 5 1 1 30021
0 30023 7 1 2 30018 30022
0 30024 7 1 2 30014 30023
0 30025 7 1 2 30012 30024
0 30026 5 1 1 30025
0 30027 7 1 2 82331 30026
0 30028 5 1 1 30027
0 30029 7 1 2 29989 30028
0 30030 5 1 1 30029
0 30031 7 1 2 97798 30030
0 30032 5 1 1 30031
0 30033 7 2 2 64745 91020
0 30034 7 1 2 78791 80392
0 30035 5 2 1 30034
0 30036 7 1 2 62120 94293
0 30037 5 1 1 30036
0 30038 7 1 2 97834 30037
0 30039 5 1 1 30038
0 30040 7 1 2 75352 30039
0 30041 5 1 1 30040
0 30042 7 3 2 73261 86351
0 30043 7 1 2 76002 72226
0 30044 7 1 2 97836 30043
0 30045 5 1 1 30044
0 30046 7 1 2 30041 30045
0 30047 5 1 1 30046
0 30048 7 1 2 63349 30047
0 30049 5 1 1 30048
0 30050 7 1 2 77395 93978
0 30051 5 1 1 30050
0 30052 7 1 2 62854 90017
0 30053 7 1 2 97823 30052
0 30054 5 1 1 30053
0 30055 7 1 2 30051 30054
0 30056 5 1 1 30055
0 30057 7 1 2 70718 30056
0 30058 5 1 1 30057
0 30059 7 1 2 79842 93486
0 30060 5 1 1 30059
0 30061 7 1 2 86436 74455
0 30062 7 1 2 92616 30061
0 30063 5 1 1 30062
0 30064 7 1 2 30060 30063
0 30065 7 1 2 30058 30064
0 30066 5 1 1 30065
0 30067 7 1 2 81772 30066
0 30068 5 1 1 30067
0 30069 7 1 2 30049 30068
0 30070 5 1 1 30069
0 30071 7 1 2 66503 30070
0 30072 5 1 1 30071
0 30073 7 1 2 73215 97821
0 30074 5 1 1 30073
0 30075 7 1 2 73262 506
0 30076 5 1 1 30075
0 30077 7 1 2 70368 30076
0 30078 7 2 2 30074 30077
0 30079 7 1 2 68187 97839
0 30080 5 1 1 30079
0 30081 7 1 2 84793 97837
0 30082 5 1 1 30081
0 30083 7 1 2 30080 30082
0 30084 5 1 1 30083
0 30085 7 1 2 75625 30084
0 30086 5 1 1 30085
0 30087 7 1 2 66975 88949
0 30088 7 1 2 94148 30087
0 30089 5 1 1 30088
0 30090 7 1 2 30086 30089
0 30091 5 1 1 30090
0 30092 7 1 2 76051 30091
0 30093 5 1 1 30092
0 30094 7 1 2 30072 30093
0 30095 5 1 1 30094
0 30096 7 1 2 66750 30095
0 30097 5 1 1 30096
0 30098 7 1 2 81736 97840
0 30099 5 1 1 30098
0 30100 7 2 2 68188 97838
0 30101 7 1 2 75576 97841
0 30102 5 1 1 30101
0 30103 7 1 2 30099 30102
0 30104 5 1 1 30103
0 30105 7 1 2 66504 30104
0 30106 5 1 1 30105
0 30107 7 3 2 61608 80951
0 30108 7 1 2 97842 97843
0 30109 5 1 1 30108
0 30110 7 1 2 30106 30109
0 30111 5 1 1 30110
0 30112 7 1 2 77705 30111
0 30113 5 1 1 30112
0 30114 7 1 2 30097 30113
0 30115 5 1 1 30114
0 30116 7 1 2 70937 30115
0 30117 5 1 1 30116
0 30118 7 4 2 68189 75961
0 30119 7 1 2 75577 97846
0 30120 5 2 1 30119
0 30121 7 1 2 87647 89631
0 30122 5 1 1 30121
0 30123 7 1 2 97850 30122
0 30124 5 3 1 30123
0 30125 7 1 2 61887 97852
0 30126 5 1 1 30125
0 30127 7 1 2 76672 97804
0 30128 5 1 1 30127
0 30129 7 1 2 30126 30128
0 30130 5 1 1 30129
0 30131 7 1 2 66505 30130
0 30132 5 1 1 30131
0 30133 7 1 2 68190 90547
0 30134 5 1 1 30133
0 30135 7 1 2 30132 30134
0 30136 5 1 1 30135
0 30137 7 1 2 71581 30136
0 30138 5 1 1 30137
0 30139 7 3 2 65441 83122
0 30140 7 1 2 73690 97844
0 30141 7 1 2 97855 30140
0 30142 5 1 1 30141
0 30143 7 1 2 30138 30142
0 30144 5 1 1 30143
0 30145 7 1 2 87894 30144
0 30146 5 1 1 30145
0 30147 7 1 2 30117 30146
0 30148 5 1 1 30147
0 30149 7 1 2 64145 30148
0 30150 5 1 1 30149
0 30151 7 1 2 86161 89596
0 30152 7 1 2 94267 30151
0 30153 5 1 1 30152
0 30154 7 1 2 89937 89603
0 30155 7 1 2 94310 30154
0 30156 5 1 1 30155
0 30157 7 1 2 30153 30156
0 30158 5 1 1 30157
0 30159 7 1 2 62121 30158
0 30160 5 1 1 30159
0 30161 7 1 2 86217 91434
0 30162 5 1 1 30161
0 30163 7 3 2 70719 89716
0 30164 5 2 1 97858
0 30165 7 2 2 30162 97861
0 30166 5 1 1 97863
0 30167 7 1 2 75582 30166
0 30168 5 1 1 30167
0 30169 7 1 2 30160 30168
0 30170 5 1 1 30169
0 30171 7 1 2 66506 30170
0 30172 5 1 1 30171
0 30173 7 1 2 86218 97811
0 30174 5 1 1 30173
0 30175 7 1 2 66976 97859
0 30176 5 1 1 30175
0 30177 7 1 2 30174 30176
0 30178 5 1 1 30177
0 30179 7 1 2 86686 30178
0 30180 5 1 1 30179
0 30181 7 1 2 30172 30180
0 30182 5 1 1 30181
0 30183 7 1 2 63350 30182
0 30184 5 1 1 30183
0 30185 7 1 2 77396 90136
0 30186 5 1 1 30185
0 30187 7 1 2 1328 30186
0 30188 5 1 1 30187
0 30189 7 1 2 73216 30188
0 30190 5 1 1 30189
0 30191 7 6 2 65777 87475
0 30192 5 1 1 97865
0 30193 7 1 2 83616 97866
0 30194 5 1 1 30193
0 30195 7 1 2 68856 80538
0 30196 7 1 2 97812 30195
0 30197 5 1 1 30196
0 30198 7 1 2 30194 30197
0 30199 5 1 1 30198
0 30200 7 1 2 86415 30199
0 30201 5 1 1 30200
0 30202 7 1 2 30190 30201
0 30203 5 1 1 30202
0 30204 7 1 2 88814 30203
0 30205 5 1 1 30204
0 30206 7 1 2 30184 30205
0 30207 5 1 1 30206
0 30208 7 1 2 66751 30207
0 30209 5 1 1 30208
0 30210 7 1 2 66507 97853
0 30211 5 1 1 30210
0 30212 7 1 2 97847 97845
0 30213 5 1 1 30212
0 30214 7 1 2 30211 30213
0 30215 5 1 1 30214
0 30216 7 1 2 70995 71694
0 30217 5 1 1 30216
0 30218 7 1 2 77784 30217
0 30219 5 1 1 30218
0 30220 7 1 2 30215 30219
0 30221 5 1 1 30220
0 30222 7 2 2 76166 81289
0 30223 5 1 1 97871
0 30224 7 1 2 75628 5125
0 30225 5 1 1 30224
0 30226 7 1 2 65442 79821
0 30227 7 1 2 30225 30226
0 30228 7 1 2 97872 30227
0 30229 5 1 1 30228
0 30230 7 4 2 77799 79258
0 30231 7 1 2 81285 80825
0 30232 7 1 2 97873 30231
0 30233 5 1 1 30232
0 30234 7 1 2 30229 30233
0 30235 5 1 1 30234
0 30236 7 1 2 94237 30235
0 30237 5 1 1 30236
0 30238 7 1 2 30221 30237
0 30239 5 1 1 30238
0 30240 7 1 2 71582 30239
0 30241 5 1 1 30240
0 30242 7 1 2 74957 96534
0 30243 7 1 2 83866 30242
0 30244 7 1 2 85584 30243
0 30245 5 1 1 30244
0 30246 7 1 2 30241 30245
0 30247 7 1 2 30209 30246
0 30248 7 1 2 30150 30247
0 30249 5 1 1 30248
0 30250 7 1 2 69372 30249
0 30251 5 1 1 30250
0 30252 7 2 2 64529 84530
0 30253 7 1 2 79858 73217
0 30254 7 1 2 94781 30253
0 30255 7 1 2 97877 30254
0 30256 5 1 1 30255
0 30257 7 1 2 30251 30256
0 30258 5 1 1 30257
0 30259 7 1 2 97832 30258
0 30260 5 1 1 30259
0 30261 7 1 2 30032 30260
0 30262 5 1 1 30261
0 30263 7 1 2 93902 30262
0 30264 5 1 1 30263
0 30265 7 6 2 90707 97625
0 30266 7 2 2 80476 92399
0 30267 7 2 2 71781 72917
0 30268 7 1 2 97885 97887
0 30269 5 1 1 30268
0 30270 7 2 2 72557 86174
0 30271 7 1 2 61888 97889
0 30272 5 1 1 30271
0 30273 7 1 2 30269 30272
0 30274 5 1 1 30273
0 30275 7 1 2 66977 30274
0 30276 5 1 1 30275
0 30277 7 1 2 73974 93961
0 30278 5 1 1 30277
0 30279 7 1 2 18533 30278
0 30280 5 2 1 30279
0 30281 7 2 2 62122 97891
0 30282 5 1 1 97893
0 30283 7 1 2 66752 97894
0 30284 5 1 1 30283
0 30285 7 1 2 30276 30284
0 30286 5 1 1 30285
0 30287 7 1 2 71731 30286
0 30288 5 1 1 30287
0 30289 7 2 2 62123 94426
0 30290 7 1 2 82056 97895
0 30291 5 1 1 30290
0 30292 7 1 2 30288 30291
0 30293 5 1 1 30292
0 30294 7 1 2 78888 30293
0 30295 5 1 1 30294
0 30296 7 1 2 75962 72227
0 30297 7 1 2 74248 30296
0 30298 7 1 2 91163 77751
0 30299 7 1 2 30297 30298
0 30300 5 1 1 30299
0 30301 7 1 2 30295 30300
0 30302 5 1 1 30301
0 30303 7 1 2 61609 30302
0 30304 5 1 1 30303
0 30305 7 2 2 65443 75708
0 30306 7 1 2 92382 97897
0 30307 5 1 1 30306
0 30308 7 1 2 70369 95843
0 30309 7 1 2 97888 30308
0 30310 5 1 1 30309
0 30311 7 1 2 30307 30310
0 30312 5 1 1 30311
0 30313 7 1 2 66978 30312
0 30314 5 1 1 30313
0 30315 7 1 2 90469 91077
0 30316 5 1 1 30315
0 30317 7 1 2 30314 30316
0 30318 5 1 1 30317
0 30319 7 1 2 63809 30318
0 30320 5 1 1 30319
0 30321 7 1 2 80500 88412
0 30322 7 1 2 89794 30321
0 30323 5 1 1 30322
0 30324 7 1 2 30320 30323
0 30325 5 1 1 30324
0 30326 7 1 2 92385 30325
0 30327 5 1 1 30326
0 30328 7 1 2 30304 30327
0 30329 5 1 1 30328
0 30330 7 1 2 63351 30329
0 30331 5 1 1 30330
0 30332 7 2 2 86613 72918
0 30333 7 1 2 97899 97886
0 30334 5 1 1 30333
0 30335 7 1 2 30282 30334
0 30336 5 1 1 30335
0 30337 7 2 2 68191 30336
0 30338 5 1 1 97901
0 30339 7 4 2 64746 71732
0 30340 7 1 2 96694 97903
0 30341 7 1 2 97902 30340
0 30342 5 1 1 30341
0 30343 7 1 2 30331 30342
0 30344 5 1 1 30343
0 30345 7 1 2 64530 30344
0 30346 5 1 1 30345
0 30347 7 1 2 72558 93939
0 30348 5 2 1 30347
0 30349 7 1 2 73811 94276
0 30350 5 1 1 30349
0 30351 7 1 2 97907 30350
0 30352 5 1 1 30351
0 30353 7 1 2 67269 30352
0 30354 5 1 1 30353
0 30355 7 1 2 72291 97809
0 30356 5 1 1 30355
0 30357 7 1 2 30354 30356
0 30358 5 1 1 30357
0 30359 7 1 2 71245 30358
0 30360 5 2 1 30359
0 30361 7 2 2 66979 71494
0 30362 7 1 2 86124 97911
0 30363 5 1 1 30362
0 30364 7 1 2 97909 30363
0 30365 5 1 1 30364
0 30366 7 2 2 64747 88918
0 30367 7 1 2 84221 97913
0 30368 7 1 2 30365 30367
0 30369 5 1 1 30368
0 30370 7 1 2 30346 30369
0 30371 5 1 1 30370
0 30372 7 1 2 69816 30371
0 30373 5 1 1 30372
0 30374 7 1 2 79879 85717
0 30375 5 1 1 30374
0 30376 7 5 2 64953 71733
0 30377 7 1 2 71842 97915
0 30378 5 1 1 30377
0 30379 7 1 2 30375 30378
0 30380 5 1 1 30379
0 30381 7 1 2 62124 30380
0 30382 5 1 1 30381
0 30383 7 2 2 66980 76777
0 30384 7 1 2 70720 93268
0 30385 5 1 1 30384
0 30386 7 2 2 91618 30385
0 30387 5 1 1 97922
0 30388 7 2 2 68663 30387
0 30389 5 2 1 97924
0 30390 7 1 2 85095 97926
0 30391 5 1 1 30390
0 30392 7 1 2 97920 30391
0 30393 5 1 1 30392
0 30394 7 1 2 30382 30393
0 30395 5 1 1 30394
0 30396 7 1 2 86878 30395
0 30397 5 1 1 30396
0 30398 7 1 2 76639 86855
0 30399 5 1 1 30398
0 30400 7 1 2 67270 30399
0 30401 5 1 1 30400
0 30402 7 1 2 74546 77318
0 30403 5 1 1 30402
0 30404 7 1 2 30401 30403
0 30405 5 1 1 30404
0 30406 7 1 2 71246 30405
0 30407 5 1 1 30406
0 30408 7 2 2 70721 89815
0 30409 7 1 2 79822 97928
0 30410 5 1 1 30409
0 30411 7 1 2 30407 30410
0 30412 5 1 1 30411
0 30413 7 1 2 84235 30412
0 30414 5 1 1 30413
0 30415 7 1 2 30397 30414
0 30416 5 1 1 30415
0 30417 7 1 2 66007 30416
0 30418 5 1 1 30417
0 30419 7 2 2 75595 83896
0 30420 5 1 1 97930
0 30421 7 1 2 90458 92067
0 30422 5 1 1 30421
0 30423 7 1 2 30420 30422
0 30424 5 1 1 30423
0 30425 7 1 2 86055 30424
0 30426 5 1 1 30425
0 30427 7 2 2 79447 80297
0 30428 7 1 2 95965 97932
0 30429 5 1 1 30428
0 30430 7 1 2 30426 30429
0 30431 5 1 1 30430
0 30432 7 1 2 68664 30431
0 30433 5 1 1 30432
0 30434 7 2 2 85364 87132
0 30435 7 1 2 83977 97934
0 30436 5 1 1 30435
0 30437 7 1 2 30433 30436
0 30438 5 1 1 30437
0 30439 7 1 2 67271 30438
0 30440 5 1 1 30439
0 30441 7 1 2 74547 89427
0 30442 7 1 2 97935 30441
0 30443 5 1 1 30442
0 30444 7 1 2 30440 30443
0 30445 5 1 1 30444
0 30446 7 1 2 65778 30445
0 30447 5 1 1 30446
0 30448 7 1 2 30418 30447
0 30449 5 1 1 30448
0 30450 7 1 2 69010 30449
0 30451 5 1 1 30450
0 30452 7 1 2 83910 84988
0 30453 5 1 1 30452
0 30454 7 1 2 83900 87982
0 30455 5 1 1 30454
0 30456 7 1 2 30453 30455
0 30457 5 1 1 30456
0 30458 7 1 2 86056 30457
0 30459 5 1 1 30458
0 30460 7 1 2 74972 91054
0 30461 7 1 2 96935 30460
0 30462 5 1 1 30461
0 30463 7 1 2 30459 30462
0 30464 5 1 1 30463
0 30465 7 1 2 68665 30464
0 30466 5 1 1 30465
0 30467 7 1 2 69373 96936
0 30468 7 1 2 87223 30467
0 30469 5 1 1 30468
0 30470 7 1 2 30466 30469
0 30471 5 1 1 30470
0 30472 7 1 2 68857 30471
0 30473 5 1 1 30472
0 30474 7 1 2 62125 75709
0 30475 7 1 2 90820 30474
0 30476 7 1 2 84244 30475
0 30477 5 1 1 30476
0 30478 7 1 2 30473 30477
0 30479 5 1 1 30478
0 30480 7 1 2 67475 30479
0 30481 5 1 1 30480
0 30482 7 2 2 66753 90120
0 30483 7 1 2 97933 97936
0 30484 5 1 1 30483
0 30485 7 2 2 90768 81536
0 30486 7 1 2 86588 97938
0 30487 5 1 1 30486
0 30488 7 1 2 30484 30487
0 30489 5 1 1 30488
0 30490 7 1 2 65779 84337
0 30491 7 1 2 30489 30490
0 30492 5 1 1 30491
0 30493 7 1 2 30481 30492
0 30494 5 1 1 30493
0 30495 7 1 2 67272 30494
0 30496 5 1 1 30495
0 30497 7 1 2 92378 15926
0 30498 5 1 1 30497
0 30499 7 1 2 87428 90121
0 30500 7 1 2 93307 30499
0 30501 7 1 2 30498 30500
0 30502 5 1 1 30501
0 30503 7 1 2 63352 30502
0 30504 7 1 2 30496 30503
0 30505 7 1 2 30451 30504
0 30506 5 1 1 30505
0 30507 7 3 2 64531 75253
0 30508 7 3 2 83532 97940
0 30509 7 1 2 86630 73331
0 30510 5 3 1 30509
0 30511 7 1 2 85252 73812
0 30512 5 1 1 30511
0 30513 7 1 2 97946 30512
0 30514 5 1 1 30513
0 30515 7 1 2 97943 30514
0 30516 5 1 1 30515
0 30517 7 2 2 76431 91953
0 30518 5 1 1 97949
0 30519 7 1 2 77744 77629
0 30520 5 2 1 30519
0 30521 7 1 2 30518 97951
0 30522 5 1 1 30521
0 30523 7 1 2 66981 30522
0 30524 5 1 1 30523
0 30525 7 1 2 74559 29306
0 30526 5 2 1 30525
0 30527 7 1 2 75481 97953
0 30528 5 1 1 30527
0 30529 7 1 2 30524 30528
0 30530 5 1 1 30529
0 30531 7 1 2 79640 30530
0 30532 5 1 1 30531
0 30533 7 1 2 30516 30532
0 30534 5 1 1 30533
0 30535 7 1 2 74985 30534
0 30536 5 1 1 30535
0 30537 7 2 2 84606 79641
0 30538 7 2 2 71782 75224
0 30539 7 1 2 83465 97957
0 30540 7 1 2 97955 30539
0 30541 5 1 1 30540
0 30542 7 1 2 30536 30541
0 30543 5 1 1 30542
0 30544 7 1 2 70722 30543
0 30545 5 1 1 30544
0 30546 7 2 2 64748 82172
0 30547 7 1 2 64146 90863
0 30548 7 1 2 97959 30547
0 30549 7 1 2 89995 30548
0 30550 5 1 1 30549
0 30551 7 1 2 68192 30550
0 30552 7 1 2 30545 30551
0 30553 5 1 1 30552
0 30554 7 1 2 76167 30553
0 30555 7 1 2 30506 30554
0 30556 5 1 1 30555
0 30557 7 1 2 86536 97912
0 30558 5 1 1 30557
0 30559 7 1 2 97910 30558
0 30560 5 1 1 30559
0 30561 7 1 2 67705 30560
0 30562 5 1 1 30561
0 30563 7 1 2 75074 77423
0 30564 7 1 2 84202 30563
0 30565 5 1 1 30564
0 30566 7 1 2 30562 30565
0 30567 5 1 1 30566
0 30568 7 1 2 92001 30567
0 30569 5 1 1 30568
0 30570 7 3 2 74845 84622
0 30571 7 2 2 84794 77347
0 30572 5 1 1 97964
0 30573 7 1 2 97961 97965
0 30574 5 1 1 30573
0 30575 7 1 2 84795 97890
0 30576 5 1 1 30575
0 30577 7 1 2 30338 30576
0 30578 5 1 1 30577
0 30579 7 1 2 70370 30578
0 30580 5 1 1 30579
0 30581 7 1 2 30574 30580
0 30582 5 1 1 30581
0 30583 7 1 2 70723 30582
0 30584 5 1 1 30583
0 30585 7 1 2 84863 97896
0 30586 5 1 1 30585
0 30587 7 1 2 30584 30586
0 30588 5 1 1 30587
0 30589 7 1 2 81089 30588
0 30590 5 1 1 30589
0 30591 7 1 2 30569 30590
0 30592 5 1 1 30591
0 30593 7 1 2 69583 30592
0 30594 5 1 1 30593
0 30595 7 1 2 93318 96223
0 30596 5 1 1 30595
0 30597 7 1 2 80121 87341
0 30598 5 1 1 30597
0 30599 7 1 2 89443 95500
0 30600 5 2 1 30599
0 30601 7 1 2 30598 97966
0 30602 5 1 1 30601
0 30603 7 1 2 73332 30602
0 30604 5 1 1 30603
0 30605 7 1 2 30596 30604
0 30606 5 1 1 30605
0 30607 7 1 2 62855 30606
0 30608 5 1 1 30607
0 30609 7 1 2 87517 81251
0 30610 7 1 2 96251 30609
0 30611 5 1 1 30610
0 30612 7 1 2 30608 30611
0 30613 5 1 1 30612
0 30614 7 1 2 97805 30613
0 30615 5 1 1 30614
0 30616 7 1 2 94471 97273
0 30617 5 1 1 30616
0 30618 7 1 2 71115 30617
0 30619 5 1 1 30618
0 30620 7 1 2 67273 76250
0 30621 7 1 2 75075 30620
0 30622 5 1 1 30621
0 30623 7 1 2 30619 30622
0 30624 5 1 1 30623
0 30625 7 1 2 79448 76024
0 30626 7 1 2 91763 30625
0 30627 7 1 2 30624 30626
0 30628 5 1 1 30627
0 30629 7 1 2 66754 30628
0 30630 7 1 2 30615 30629
0 30631 7 1 2 30594 30630
0 30632 5 1 1 30631
0 30633 7 1 2 85964 80100
0 30634 7 2 2 95885 30633
0 30635 5 1 1 97968
0 30636 7 1 2 66982 97969
0 30637 5 1 1 30636
0 30638 7 1 2 64147 97829
0 30639 5 1 1 30638
0 30640 7 1 2 75372 97824
0 30641 5 1 1 30640
0 30642 7 1 2 30639 30641
0 30643 5 1 1 30642
0 30644 7 1 2 70938 82548
0 30645 7 1 2 30643 30644
0 30646 5 1 1 30645
0 30647 7 1 2 30637 30646
0 30648 5 1 1 30647
0 30649 7 1 2 81090 30648
0 30650 5 1 1 30649
0 30651 7 1 2 62126 92503
0 30652 5 1 1 30651
0 30653 7 1 2 97947 30652
0 30654 5 2 1 30653
0 30655 7 1 2 72065 81737
0 30656 7 1 2 91771 30655
0 30657 7 1 2 97970 30656
0 30658 5 1 1 30657
0 30659 7 1 2 30650 30658
0 30660 5 1 1 30659
0 30661 7 1 2 70371 30660
0 30662 5 1 1 30661
0 30663 7 1 2 81738 90393
0 30664 7 3 2 64749 84017
0 30665 7 1 2 97972 97874
0 30666 7 1 2 30663 30665
0 30667 5 1 1 30666
0 30668 7 1 2 30662 30667
0 30669 5 1 1 30668
0 30670 7 1 2 70724 30669
0 30671 5 1 1 30670
0 30672 7 2 2 65780 82990
0 30673 7 1 2 86672 94152
0 30674 7 1 2 97975 30673
0 30675 7 1 2 95404 30674
0 30676 5 1 1 30675
0 30677 7 2 2 61889 30676
0 30678 7 1 2 30671 97977
0 30679 5 1 1 30678
0 30680 7 1 2 64954 30679
0 30681 7 1 2 30632 30680
0 30682 5 1 1 30681
0 30683 7 1 2 30556 30682
0 30684 7 1 2 30373 30683
0 30685 5 1 1 30684
0 30686 7 1 2 97879 30685
0 30687 5 1 1 30686
0 30688 7 23 2 67783 69102
0 30689 7 29 2 90659 97979
0 30690 7 1 2 75034 94277
0 30691 5 1 1 30690
0 30692 7 1 2 97908 30691
0 30693 5 1 1 30692
0 30694 7 1 2 78999 30693
0 30695 5 1 1 30694
0 30696 7 2 2 76003 84405
0 30697 7 1 2 72454 98031
0 30698 7 1 2 97937 30697
0 30699 5 1 1 30698
0 30700 7 1 2 30695 30699
0 30701 5 1 1 30700
0 30702 7 1 2 98002 30701
0 30703 5 1 1 30702
0 30704 7 1 2 96640 29439
0 30705 5 1 1 30704
0 30706 7 1 2 80983 30705
0 30707 5 1 1 30706
0 30708 7 1 2 81005 94238
0 30709 7 1 2 96781 30708
0 30710 5 1 1 30709
0 30711 7 1 2 30707 30710
0 30712 5 1 1 30711
0 30713 7 1 2 77272 77559
0 30714 7 1 2 97658 30713
0 30715 7 1 2 30712 30714
0 30716 5 1 1 30715
0 30717 7 1 2 30703 30716
0 30718 5 1 1 30717
0 30719 7 1 2 69374 30718
0 30720 5 1 1 30719
0 30721 7 1 2 85408 97659
0 30722 5 1 1 30721
0 30723 7 13 2 69103 65444
0 30724 7 7 2 62127 67850
0 30725 7 3 2 97456 98046
0 30726 7 2 2 98033 98053
0 30727 5 1 1 98056
0 30728 7 1 2 66008 98057
0 30729 5 1 1 30728
0 30730 7 1 2 30722 30729
0 30731 5 2 1 30730
0 30732 7 1 2 78930 98058
0 30733 5 1 1 30732
0 30734 7 1 2 64750 95188
0 30735 7 1 2 87476 30734
0 30736 7 1 2 98054 30735
0 30737 5 1 1 30736
0 30738 7 1 2 30733 30737
0 30739 5 1 1 30738
0 30740 7 1 2 81999 30739
0 30741 5 1 1 30740
0 30742 7 2 2 75482 98003
0 30743 7 1 2 76004 95224
0 30744 7 1 2 98060 30743
0 30745 5 1 1 30744
0 30746 7 1 2 30741 30745
0 30747 5 1 1 30746
0 30748 7 1 2 61610 30747
0 30749 5 1 1 30748
0 30750 7 1 2 95018 98059
0 30751 5 1 1 30750
0 30752 7 1 2 30749 30751
0 30753 5 1 1 30752
0 30754 7 1 2 96087 30753
0 30755 5 1 1 30754
0 30756 7 1 2 30720 30755
0 30757 5 1 1 30756
0 30758 7 1 2 68858 30757
0 30759 5 1 1 30758
0 30760 7 4 2 98034 97465
0 30761 7 1 2 82682 97065
0 30762 7 1 2 98062 30761
0 30763 7 1 2 95023 30762
0 30764 5 1 1 30763
0 30765 7 1 2 30759 30764
0 30766 5 1 1 30765
0 30767 7 1 2 67476 30766
0 30768 5 1 1 30767
0 30769 7 1 2 66983 97944
0 30770 5 2 1 30769
0 30771 7 1 2 85597 93308
0 30772 5 1 1 30771
0 30773 7 1 2 98066 30772
0 30774 5 1 1 30773
0 30775 7 1 2 97660 30774
0 30776 5 1 1 30775
0 30777 7 4 2 66984 67851
0 30778 7 5 2 97457 98068
0 30779 7 6 2 69104 98072
0 30780 7 1 2 83901 98077
0 30781 7 1 2 97929 30780
0 30782 5 1 1 30781
0 30783 7 1 2 30776 30782
0 30784 5 1 1 30783
0 30785 7 1 2 66009 30784
0 30786 5 1 1 30785
0 30787 7 11 2 66218 61890
0 30788 5 1 1 98083
0 30789 7 1 2 96091 98084
0 30790 7 2 2 82396 90769
0 30791 7 1 2 98094 97563
0 30792 7 1 2 30789 30791
0 30793 5 1 1 30792
0 30794 7 1 2 30786 30793
0 30795 5 1 1 30794
0 30796 7 1 2 69011 30795
0 30797 5 1 1 30796
0 30798 7 1 2 74158 79479
0 30799 7 1 2 88162 30798
0 30800 5 1 1 30799
0 30801 7 1 2 82629 86319
0 30802 7 1 2 86445 30801
0 30803 5 1 1 30802
0 30804 7 1 2 30800 30803
0 30805 5 1 1 30804
0 30806 7 1 2 65781 98004
0 30807 7 1 2 30805 30806
0 30808 5 1 1 30807
0 30809 7 1 2 30797 30808
0 30810 5 1 1 30809
0 30811 7 1 2 76168 30810
0 30812 5 1 1 30811
0 30813 7 1 2 78846 91220
0 30814 5 1 1 30813
0 30815 7 1 2 82000 91238
0 30816 5 1 1 30815
0 30817 7 1 2 30814 30816
0 30818 5 1 1 30817
0 30819 7 1 2 62421 97692
0 30820 7 1 2 30818 30819
0 30821 5 1 1 30820
0 30822 7 1 2 83813 71534
0 30823 7 1 2 86772 30822
0 30824 7 1 2 97226 30823
0 30825 5 1 1 30824
0 30826 7 1 2 30821 30825
0 30827 5 1 1 30826
0 30828 7 1 2 98063 30827
0 30829 5 1 1 30828
0 30830 7 1 2 30812 30829
0 30831 7 1 2 30768 30830
0 30832 5 1 1 30831
0 30833 7 1 2 68666 30832
0 30834 5 1 1 30833
0 30835 7 1 2 83998 72424
0 30836 5 1 1 30835
0 30837 7 1 2 8294 30836
0 30838 5 1 1 30837
0 30839 7 1 2 82001 30838
0 30840 5 1 1 30839
0 30841 7 1 2 70725 82604
0 30842 7 1 2 94239 30841
0 30843 7 1 2 78955 30842
0 30844 5 1 1 30843
0 30845 7 1 2 30840 30844
0 30846 5 1 1 30845
0 30847 7 1 2 71247 30846
0 30848 5 1 1 30847
0 30849 7 1 2 88857 96088
0 30850 7 1 2 97500 30849
0 30851 5 1 1 30850
0 30852 7 1 2 30848 30851
0 30853 5 1 1 30852
0 30854 7 1 2 73990 30853
0 30855 5 1 1 30854
0 30856 7 2 2 70726 78977
0 30857 7 1 2 81867 95498
0 30858 7 1 2 98096 30857
0 30859 5 1 1 30858
0 30860 7 1 2 30855 30859
0 30861 5 1 1 30860
0 30862 7 1 2 98005 30861
0 30863 5 1 1 30862
0 30864 7 1 2 64532 95445
0 30865 7 1 2 96507 30864
0 30866 7 16 2 63001 63176
0 30867 7 4 2 62959 98098
0 30868 7 2 2 61350 82057
0 30869 7 1 2 98114 98118
0 30870 7 1 2 30865 30869
0 30871 5 1 1 30870
0 30872 7 1 2 30863 30871
0 30873 5 1 1 30872
0 30874 7 1 2 66985 30873
0 30875 5 1 1 30874
0 30876 7 5 2 63002 68859
0 30877 7 3 2 91797 98120
0 30878 7 2 2 61351 69012
0 30879 7 1 2 85032 94632
0 30880 7 1 2 98128 30879
0 30881 7 1 2 98125 30880
0 30882 7 1 2 98097 30881
0 30883 5 1 1 30882
0 30884 7 1 2 30875 30883
0 30885 5 1 1 30884
0 30886 7 1 2 66508 30885
0 30887 5 1 1 30886
0 30888 7 2 2 69013 76052
0 30889 7 3 2 74973 88122
0 30890 7 1 2 69375 89881
0 30891 7 1 2 98132 30890
0 30892 5 1 1 30891
0 30893 7 1 2 98067 30892
0 30894 5 1 1 30893
0 30895 7 1 2 97661 30894
0 30896 5 1 1 30895
0 30897 7 3 2 66219 82630
0 30898 7 6 2 68860 69105
0 30899 7 1 2 69376 98138
0 30900 7 2 2 98135 30899
0 30901 7 2 2 67477 91859
0 30902 7 2 2 88097 74974
0 30903 7 1 2 98146 98148
0 30904 7 1 2 98144 30903
0 30905 5 1 1 30904
0 30906 7 1 2 30896 30905
0 30907 5 1 1 30906
0 30908 7 1 2 67274 30907
0 30909 5 1 1 30908
0 30910 7 1 2 75515 91860
0 30911 7 1 2 98133 30910
0 30912 7 1 2 98145 30911
0 30913 5 1 1 30912
0 30914 7 1 2 30909 30913
0 30915 5 1 1 30914
0 30916 7 1 2 98130 30915
0 30917 5 1 1 30916
0 30918 7 1 2 30887 30917
0 30919 5 1 1 30918
0 30920 7 1 2 66010 30919
0 30921 5 1 1 30920
0 30922 7 1 2 69817 81520
0 30923 7 1 2 90976 30922
0 30924 7 7 2 64258 65445
0 30925 7 2 2 77419 98150
0 30926 7 1 2 98157 98119
0 30927 7 1 2 30923 30926
0 30928 5 1 1 30927
0 30929 7 5 2 69106 64955
0 30930 7 1 2 76673 98159
0 30931 7 1 2 98073 30930
0 30932 7 1 2 94473 30931
0 30933 5 1 1 30932
0 30934 7 1 2 30928 30933
0 30935 5 1 1 30934
0 30936 7 1 2 87143 91674
0 30937 7 1 2 30935 30936
0 30938 5 1 1 30937
0 30939 7 1 2 63353 30938
0 30940 7 1 2 30921 30939
0 30941 7 1 2 30834 30940
0 30942 5 1 1 30941
0 30943 7 1 2 82241 82536
0 30944 7 5 2 90977 95147
0 30945 7 3 2 61352 67478
0 30946 7 3 2 69584 98169
0 30947 7 1 2 98164 98172
0 30948 7 1 2 30943 30947
0 30949 5 2 1 30948
0 30950 7 8 2 63810 69107
0 30951 7 3 2 67784 98177
0 30952 7 4 2 90660 98185
0 30953 7 1 2 89632 98188
0 30954 7 1 2 97956 30953
0 30955 5 1 1 30954
0 30956 7 1 2 98175 30955
0 30957 5 1 1 30956
0 30958 7 1 2 70727 30957
0 30959 5 1 1 30958
0 30960 7 6 2 64259 90978
0 30961 7 4 2 61353 66986
0 30962 7 1 2 83814 98198
0 30963 7 1 2 98192 30962
0 30964 7 1 2 96511 30963
0 30965 5 1 1 30964
0 30966 7 1 2 30959 30965
0 30967 5 1 1 30966
0 30968 7 1 2 72559 30967
0 30969 5 1 1 30968
0 30970 7 1 2 77151 90864
0 30971 7 1 2 98178 30970
0 30972 7 3 2 91360 97458
0 30973 7 1 2 83276 98202
0 30974 7 1 2 30971 30973
0 30975 5 1 1 30974
0 30976 7 1 2 98176 30975
0 30977 5 1 1 30976
0 30978 7 1 2 79684 30977
0 30979 5 1 1 30978
0 30980 7 1 2 30969 30979
0 30981 5 1 1 30980
0 30982 7 1 2 61611 30981
0 30983 5 1 1 30982
0 30984 7 7 2 69108 64751
0 30985 7 4 2 82605 98205
0 30986 7 1 2 90031 74456
0 30987 7 1 2 91886 30986
0 30988 7 1 2 98212 30987
0 30989 7 1 2 97132 30988
0 30990 5 1 1 30989
0 30991 7 1 2 30983 30990
0 30992 5 1 1 30991
0 30993 7 1 2 66755 30992
0 30994 5 1 1 30993
0 30995 7 1 2 71248 91476
0 30996 5 1 1 30995
0 30997 7 1 2 62128 91411
0 30998 5 1 1 30997
0 30999 7 1 2 30996 30998
0 31000 5 1 1 30999
0 31001 7 1 2 66509 31000
0 31002 5 1 1 31001
0 31003 7 1 2 89085 86057
0 31004 5 1 1 31003
0 31005 7 1 2 31002 31004
0 31006 5 1 1 31005
0 31007 7 4 2 61354 67275
0 31008 7 2 2 90979 98216
0 31009 7 3 2 66011 95446
0 31010 7 1 2 71062 88689
0 31011 7 1 2 98222 31010
0 31012 7 1 2 98220 31011
0 31013 7 1 2 31006 31012
0 31014 5 1 1 31013
0 31015 7 1 2 68193 31014
0 31016 7 1 2 30994 31015
0 31017 5 1 1 31016
0 31018 7 1 2 67706 31017
0 31019 7 1 2 30942 31018
0 31020 5 1 1 31019
0 31021 7 1 2 97474 30572
0 31022 5 1 1 31021
0 31023 7 1 2 85253 31022
0 31024 5 1 1 31023
0 31025 7 2 2 63354 72228
0 31026 7 1 2 76251 76734
0 31027 7 1 2 98225 31026
0 31028 5 1 1 31027
0 31029 7 1 2 31024 31028
0 31030 5 1 1 31029
0 31031 7 1 2 70728 31030
0 31032 5 1 1 31031
0 31033 7 2 2 62129 86574
0 31034 7 1 2 85516 78006
0 31035 7 1 2 98227 31034
0 31036 5 1 1 31035
0 31037 7 1 2 31032 31036
0 31038 5 1 1 31037
0 31039 7 1 2 76169 31038
0 31040 5 1 1 31039
0 31041 7 1 2 77276 97279
0 31042 5 1 1 31041
0 31043 7 1 2 77842 77279
0 31044 5 2 1 31043
0 31045 7 1 2 62586 98229
0 31046 5 1 1 31045
0 31047 7 1 2 13658 31046
0 31048 5 2 1 31047
0 31049 7 1 2 93214 98231
0 31050 5 1 1 31049
0 31051 7 1 2 31042 31050
0 31052 5 1 1 31051
0 31053 7 1 2 94973 31052
0 31054 5 1 1 31053
0 31055 7 1 2 31040 31054
0 31056 5 1 1 31055
0 31057 7 1 2 69585 31056
0 31058 5 1 1 31057
0 31059 7 2 2 67276 82582
0 31060 7 1 2 97261 98233
0 31061 5 1 1 31060
0 31062 7 1 2 85147 97267
0 31063 5 1 1 31062
0 31064 7 1 2 31061 31063
0 31065 5 1 1 31064
0 31066 7 1 2 62130 31065
0 31067 5 1 1 31066
0 31068 7 1 2 84824 76608
0 31069 5 1 1 31068
0 31070 7 1 2 31067 31069
0 31071 5 1 1 31070
0 31072 7 1 2 94649 31071
0 31073 5 1 1 31072
0 31074 7 1 2 31058 31073
0 31075 5 1 1 31074
0 31076 7 1 2 68667 31075
0 31077 5 1 1 31076
0 31078 7 1 2 82583 89895
0 31079 5 1 1 31078
0 31080 7 1 2 89011 85017
0 31081 5 1 1 31080
0 31082 7 1 2 31079 31081
0 31083 5 1 1 31082
0 31084 7 1 2 88191 31083
0 31085 5 1 1 31084
0 31086 7 1 2 78700 93262
0 31087 7 2 2 64752 73854
0 31088 7 2 2 68194 73964
0 31089 7 1 2 98235 98237
0 31090 7 1 2 31086 31089
0 31091 5 1 1 31090
0 31092 7 1 2 31085 31091
0 31093 5 1 1 31092
0 31094 7 1 2 63811 31093
0 31095 5 1 1 31094
0 31096 7 1 2 78215 91954
0 31097 7 1 2 97293 31096
0 31098 5 1 1 31097
0 31099 7 1 2 31095 31098
0 31100 5 1 1 31099
0 31101 7 1 2 66987 31100
0 31102 5 1 1 31101
0 31103 7 2 2 73651 75185
0 31104 7 1 2 91527 96998
0 31105 7 1 2 98239 31104
0 31106 5 1 1 31105
0 31107 7 1 2 31102 31106
0 31108 5 1 1 31107
0 31109 7 1 2 70729 31108
0 31110 5 1 1 31109
0 31111 7 1 2 31077 31110
0 31112 5 1 1 31111
0 31113 7 1 2 61891 31112
0 31114 5 1 1 31113
0 31115 7 2 2 73652 80167
0 31116 7 1 2 97009 98241
0 31117 5 1 1 31116
0 31118 7 1 2 90770 96126
0 31119 5 1 1 31118
0 31120 7 1 2 87360 97827
0 31121 5 1 1 31120
0 31122 7 1 2 68668 90222
0 31123 7 1 2 79259 31122
0 31124 5 1 1 31123
0 31125 7 1 2 31121 31124
0 31126 5 1 1 31125
0 31127 7 1 2 70372 31126
0 31128 5 1 1 31127
0 31129 7 1 2 31119 31128
0 31130 5 1 1 31129
0 31131 7 1 2 74986 31130
0 31132 5 1 1 31131
0 31133 7 1 2 31117 31132
0 31134 5 1 1 31133
0 31135 7 1 2 76674 87093
0 31136 7 1 2 31134 31135
0 31137 5 1 1 31136
0 31138 7 1 2 31114 31137
0 31139 5 1 1 31138
0 31140 7 1 2 82242 31139
0 31141 5 1 1 31140
0 31142 7 5 2 69377 81262
0 31143 7 1 2 70373 97971
0 31144 5 1 1 31143
0 31145 7 1 2 62131 94045
0 31146 5 1 1 31145
0 31147 7 1 2 31144 31146
0 31148 5 1 1 31147
0 31149 7 1 2 98243 31148
0 31150 5 1 1 31149
0 31151 7 1 2 70374 85663
0 31152 7 1 2 92746 31151
0 31153 7 1 2 97825 31152
0 31154 5 1 1 31153
0 31155 7 1 2 31150 31154
0 31156 5 1 1 31155
0 31157 7 1 2 68195 31156
0 31158 5 1 1 31157
0 31159 7 1 2 88919 89570
0 31160 7 1 2 86352 31159
0 31161 7 1 2 81263 31160
0 31162 5 1 1 31161
0 31163 7 1 2 31158 31162
0 31164 5 1 1 31163
0 31165 7 1 2 72066 31164
0 31166 5 1 1 31165
0 31167 7 3 2 83833 80059
0 31168 7 1 2 98248 97831
0 31169 5 1 1 31168
0 31170 7 1 2 31166 31169
0 31171 5 1 1 31170
0 31172 7 1 2 62856 31171
0 31173 5 1 1 31172
0 31174 7 1 2 82268 85178
0 31175 5 1 1 31174
0 31176 7 1 2 97801 31175
0 31177 5 1 1 31176
0 31178 7 1 2 62422 31177
0 31179 5 1 1 31178
0 31180 7 1 2 72900 94437
0 31181 5 3 1 31180
0 31182 7 1 2 68669 98251
0 31183 5 1 1 31182
0 31184 7 1 2 94467 31183
0 31185 5 1 1 31184
0 31186 7 1 2 84796 31185
0 31187 5 1 1 31186
0 31188 7 1 2 31179 31187
0 31189 5 1 1 31188
0 31190 7 1 2 98249 31189
0 31191 5 1 1 31190
0 31192 7 1 2 31173 31191
0 31193 5 1 1 31192
0 31194 7 1 2 70730 31193
0 31195 5 1 1 31194
0 31196 7 4 2 84406 82438
0 31197 7 2 2 75291 98254
0 31198 5 1 1 98258
0 31199 7 1 2 83954 98230
0 31200 5 1 1 31199
0 31201 7 1 2 31198 31200
0 31202 5 1 1 31201
0 31203 7 1 2 63177 31202
0 31204 5 1 1 31203
0 31205 7 2 2 82116 78931
0 31206 7 2 2 77358 84765
0 31207 7 1 2 98260 98262
0 31208 5 1 1 31207
0 31209 7 1 2 31204 31208
0 31210 5 1 1 31209
0 31211 7 1 2 62587 31210
0 31212 5 1 1 31211
0 31213 7 2 2 82850 81472
0 31214 5 1 1 98264
0 31215 7 1 2 91067 98265
0 31216 5 1 1 31215
0 31217 7 1 2 31212 31216
0 31218 5 1 1 31217
0 31219 7 1 2 97806 31218
0 31220 5 1 1 31219
0 31221 7 1 2 80188 74625
0 31222 7 1 2 91223 31221
0 31223 5 1 1 31222
0 31224 7 1 2 65446 76093
0 31225 5 1 1 31224
0 31226 7 1 2 63812 31225
0 31227 5 1 1 31226
0 31228 7 1 2 67277 31227
0 31229 5 1 1 31228
0 31230 7 1 2 11102 31229
0 31231 5 1 1 31230
0 31232 7 1 2 69014 75978
0 31233 7 1 2 81264 31232
0 31234 7 1 2 31231 31233
0 31235 5 1 1 31234
0 31236 7 1 2 31223 31235
0 31237 5 1 1 31236
0 31238 7 1 2 84797 82439
0 31239 7 1 2 31237 31238
0 31240 5 1 1 31239
0 31241 7 1 2 31220 31240
0 31242 5 1 1 31241
0 31243 7 1 2 62857 31242
0 31244 5 1 1 31243
0 31245 7 1 2 72170 98244
0 31246 5 1 1 31245
0 31247 7 1 2 31246 31214
0 31248 5 1 1 31247
0 31249 7 1 2 65782 31248
0 31250 5 1 1 31249
0 31251 7 1 2 97967 31250
0 31252 5 1 1 31251
0 31253 7 2 2 84864 84970
0 31254 7 1 2 86058 98266
0 31255 7 1 2 31252 31254
0 31256 5 1 1 31255
0 31257 7 1 2 66756 31256
0 31258 7 1 2 31244 31257
0 31259 7 1 2 31195 31258
0 31260 5 1 1 31259
0 31261 7 2 2 92248 93302
0 31262 7 1 2 68021 88213
0 31263 7 1 2 98268 31262
0 31264 5 1 1 31263
0 31265 7 1 2 77499 88595
0 31266 7 1 2 79866 31265
0 31267 5 1 1 31266
0 31268 7 1 2 30635 31267
0 31269 5 1 1 31268
0 31270 7 1 2 70375 83815
0 31271 7 1 2 31269 31270
0 31272 5 1 1 31271
0 31273 7 1 2 31264 31272
0 31274 5 1 1 31273
0 31275 7 1 2 66988 31274
0 31276 5 1 1 31275
0 31277 7 1 2 64148 82220
0 31278 5 1 1 31277
0 31279 7 1 2 74125 85215
0 31280 5 1 1 31279
0 31281 7 1 2 31278 31280
0 31282 5 1 1 31281
0 31283 7 1 2 80254 31282
0 31284 5 1 1 31283
0 31285 7 1 2 86107 80107
0 31286 5 1 1 31285
0 31287 7 1 2 31284 31286
0 31288 5 1 1 31287
0 31289 7 1 2 84531 87495
0 31290 7 1 2 31288 31289
0 31291 5 1 1 31290
0 31292 7 1 2 61612 31291
0 31293 7 1 2 31276 31292
0 31294 5 1 1 31293
0 31295 7 2 2 87648 73610
0 31296 7 1 2 90050 98270
0 31297 5 1 1 31296
0 31298 7 1 2 68196 92877
0 31299 5 1 1 31298
0 31300 7 1 2 31297 31299
0 31301 5 1 1 31300
0 31302 7 1 2 66989 31301
0 31303 5 1 1 31302
0 31304 7 4 2 63355 74224
0 31305 7 1 2 98272 97954
0 31306 5 1 1 31305
0 31307 7 1 2 31303 31306
0 31308 5 1 1 31307
0 31309 7 1 2 83769 90388
0 31310 7 1 2 31308 31309
0 31311 5 1 1 31310
0 31312 7 1 2 84050 86688
0 31313 7 1 2 92591 31312
0 31314 5 1 1 31313
0 31315 7 1 2 66510 31314
0 31316 7 1 2 31311 31315
0 31317 5 1 1 31316
0 31318 7 1 2 70731 31317
0 31319 7 1 2 31294 31318
0 31320 5 1 1 31319
0 31321 7 1 2 97978 31320
0 31322 5 1 1 31321
0 31323 7 1 2 64956 31322
0 31324 7 1 2 31260 31323
0 31325 5 1 1 31324
0 31326 7 1 2 31141 31325
0 31327 5 1 1 31326
0 31328 7 1 2 98006 31327
0 31329 5 1 1 31328
0 31330 7 2 2 95379 95501
0 31331 5 1 1 98276
0 31332 7 1 2 71063 98277
0 31333 5 1 1 31332
0 31334 7 1 2 82332 71440
0 31335 7 1 2 86794 31334
0 31336 5 1 1 31335
0 31337 7 1 2 31333 31336
0 31338 5 1 1 31337
0 31339 7 1 2 76476 31338
0 31340 5 1 1 31339
0 31341 7 1 2 79657 89907
0 31342 7 1 2 95550 31341
0 31343 5 1 1 31342
0 31344 7 1 2 66990 75666
0 31345 5 3 1 31344
0 31346 7 1 2 70376 98278
0 31347 5 1 1 31346
0 31348 7 1 2 85155 31347
0 31349 5 1 1 31348
0 31350 7 1 2 71843 95033
0 31351 7 1 2 31349 31350
0 31352 5 1 1 31351
0 31353 7 1 2 31343 31352
0 31354 5 1 1 31353
0 31355 7 1 2 86032 31354
0 31356 5 1 1 31355
0 31357 7 1 2 31340 31356
0 31358 5 1 1 31357
0 31359 7 1 2 69586 31358
0 31360 5 1 1 31359
0 31361 7 2 2 71844 80298
0 31362 5 1 1 98281
0 31363 7 1 2 80565 97867
0 31364 5 1 1 31363
0 31365 7 1 2 31362 31364
0 31366 5 1 1 31365
0 31367 7 1 2 75483 98245
0 31368 7 1 2 31366 31367
0 31369 5 1 1 31368
0 31370 7 1 2 31360 31369
0 31371 5 1 1 31370
0 31372 7 1 2 68197 31371
0 31373 5 1 1 31372
0 31374 7 1 2 74569 89723
0 31375 5 3 1 31374
0 31376 7 1 2 77119 87297
0 31377 5 1 1 31376
0 31378 7 1 2 98283 31377
0 31379 5 1 1 31378
0 31380 7 1 2 62132 31379
0 31381 5 1 1 31380
0 31382 7 1 2 73097 27592
0 31383 5 1 1 31382
0 31384 7 1 2 63356 76477
0 31385 7 1 2 31383 31384
0 31386 5 1 1 31385
0 31387 7 1 2 31381 31386
0 31388 5 1 1 31387
0 31389 7 1 2 82333 31388
0 31390 5 1 1 31389
0 31391 7 1 2 71340 93724
0 31392 5 1 1 31391
0 31393 7 1 2 85153 31392
0 31394 5 1 1 31393
0 31395 7 1 2 62858 31394
0 31396 5 1 1 31395
0 31397 7 1 2 85162 31396
0 31398 5 1 1 31397
0 31399 7 1 2 90932 31398
0 31400 5 1 1 31399
0 31401 7 1 2 7533 98284
0 31402 5 1 1 31401
0 31403 7 1 2 62133 31402
0 31404 5 1 1 31403
0 31405 7 1 2 72871 5150
0 31406 5 1 1 31405
0 31407 7 1 2 71968 31406
0 31408 5 1 1 31407
0 31409 7 1 2 75273 91955
0 31410 5 1 1 31409
0 31411 7 1 2 31408 31410
0 31412 5 1 1 31411
0 31413 7 1 2 85226 31412
0 31414 5 1 1 31413
0 31415 7 1 2 31404 31414
0 31416 7 1 2 31400 31415
0 31417 5 1 1 31416
0 31418 7 1 2 81091 31417
0 31419 5 1 1 31418
0 31420 7 1 2 31390 31419
0 31421 5 1 1 31420
0 31422 7 1 2 79185 31421
0 31423 5 1 1 31422
0 31424 7 2 2 77397 89365
0 31425 7 1 2 71969 91675
0 31426 7 1 2 98286 31425
0 31427 5 1 1 31426
0 31428 7 1 2 71845 87480
0 31429 7 1 2 90754 31428
0 31430 7 1 2 92443 31429
0 31431 5 1 1 31430
0 31432 7 1 2 31427 31431
0 31433 5 1 1 31432
0 31434 7 1 2 70377 31433
0 31435 5 1 1 31434
0 31436 7 1 2 71655 83617
0 31437 5 1 1 31436
0 31438 7 1 2 71970 73671
0 31439 5 1 1 31438
0 31440 7 1 2 31437 31439
0 31441 5 1 1 31440
0 31442 7 1 2 90261 76778
0 31443 7 1 2 31441 31442
0 31444 5 1 1 31443
0 31445 7 1 2 31435 31444
0 31446 5 1 1 31445
0 31447 7 1 2 61892 31446
0 31448 5 1 1 31447
0 31449 7 1 2 74201 86139
0 31450 7 1 2 89337 87550
0 31451 7 1 2 31449 31450
0 31452 5 1 1 31451
0 31453 7 1 2 31448 31452
0 31454 5 1 1 31453
0 31455 7 1 2 81739 31454
0 31456 5 1 1 31455
0 31457 7 1 2 31423 31456
0 31458 7 1 2 31373 31457
0 31459 5 1 1 31458
0 31460 7 1 2 97662 31459
0 31461 5 1 1 31460
0 31462 7 1 2 31329 31461
0 31463 7 1 2 31020 31462
0 31464 5 1 1 31463
0 31465 7 1 2 61272 31464
0 31466 5 1 1 31465
0 31467 7 1 2 30687 31466
0 31468 5 1 1 31467
0 31469 7 1 2 64360 31468
0 31470 5 1 1 31469
0 31471 7 1 2 30264 31470
0 31472 7 1 2 29965 31471
0 31473 5 1 1 31472
0 31474 7 1 2 94942 31473
0 31475 5 1 1 31474
0 31476 7 4 2 14074 84769
0 31477 5 41 1 98288
0 31478 7 1 2 66991 92445
0 31479 5 1 1 31478
0 31480 7 1 2 68425 94428
0 31481 5 1 1 31480
0 31482 7 1 2 31479 31481
0 31483 5 1 1 31482
0 31484 7 1 2 63813 31483
0 31485 5 1 1 31484
0 31486 7 1 2 63578 86787
0 31487 5 1 1 31486
0 31488 7 1 2 73918 77630
0 31489 5 1 1 31488
0 31490 7 2 2 31487 31489
0 31491 5 1 1 98333
0 31492 7 1 2 31485 98334
0 31493 5 1 1 31492
0 31494 7 1 2 93592 31493
0 31495 5 1 1 31494
0 31496 7 1 2 90875 96433
0 31497 7 1 2 82831 31496
0 31498 5 1 1 31497
0 31499 7 1 2 31495 31498
0 31500 5 1 1 31499
0 31501 7 1 2 65783 31500
0 31502 5 1 1 31501
0 31503 7 2 2 65447 87939
0 31504 7 6 2 66992 62960
0 31505 7 2 2 71846 98337
0 31506 7 1 2 98335 98343
0 31507 5 1 1 31506
0 31508 7 3 2 66993 94210
0 31509 5 1 1 98345
0 31510 7 1 2 96405 31509
0 31511 5 2 1 31510
0 31512 7 2 2 71583 98348
0 31513 5 1 1 98350
0 31514 7 1 2 92171 98351
0 31515 5 1 1 31514
0 31516 7 1 2 31507 31515
0 31517 7 1 2 31502 31516
0 31518 5 1 1 31517
0 31519 7 1 2 90599 31518
0 31520 5 1 1 31519
0 31521 7 1 2 75263 96562
0 31522 5 2 1 31521
0 31523 7 1 2 31513 98352
0 31524 5 2 1 31523
0 31525 7 4 2 90661 97524
0 31526 7 1 2 98354 98356
0 31527 5 1 1 31526
0 31528 7 1 2 31520 31527
0 31529 5 1 1 31528
0 31530 7 1 2 78713 31529
0 31531 5 1 1 31530
0 31532 7 1 2 62588 80399
0 31533 5 1 1 31532
0 31534 7 1 2 71584 74289
0 31535 5 1 1 31534
0 31536 7 1 2 31533 31535
0 31537 5 4 1 31536
0 31538 7 2 2 92172 98360
0 31539 7 4 2 63178 93771
0 31540 7 2 2 74239 98366
0 31541 7 1 2 62134 98370
0 31542 7 1 2 98364 31541
0 31543 5 1 1 31542
0 31544 7 1 2 31531 31543
0 31545 5 1 1 31544
0 31546 7 1 2 61273 31545
0 31547 5 1 1 31546
0 31548 7 3 2 69214 93845
0 31549 7 1 2 79859 92848
0 31550 7 1 2 77214 31549
0 31551 5 1 1 31550
0 31552 7 1 2 84166 86162
0 31553 7 1 2 92545 31552
0 31554 5 1 1 31553
0 31555 7 1 2 31551 31554
0 31556 5 1 1 31555
0 31557 7 1 2 62135 31556
0 31558 5 1 1 31557
0 31559 7 1 2 64957 92546
0 31560 7 1 2 98346 31559
0 31561 5 1 1 31560
0 31562 7 1 2 31558 31561
0 31563 5 1 1 31562
0 31564 7 1 2 61355 31563
0 31565 5 1 1 31564
0 31566 7 2 2 77161 83514
0 31567 7 1 2 66220 98099
0 31568 7 2 2 98375 31567
0 31569 5 1 1 98377
0 31570 7 1 2 31565 31569
0 31571 5 1 1 31570
0 31572 7 1 2 71585 31571
0 31573 5 1 1 31572
0 31574 7 1 2 80400 98371
0 31575 5 1 1 31574
0 31576 7 1 2 82530 92547
0 31577 7 1 2 98217 31576
0 31578 7 1 2 84264 31577
0 31579 5 1 1 31578
0 31580 7 1 2 31575 31579
0 31581 5 1 1 31580
0 31582 7 1 2 75854 31581
0 31583 5 1 1 31582
0 31584 7 1 2 31573 31583
0 31585 5 1 1 31584
0 31586 7 1 2 98372 31585
0 31587 5 1 1 31586
0 31588 7 1 2 31547 31587
0 31589 5 1 1 31588
0 31590 7 1 2 83123 31589
0 31591 5 1 1 31590
0 31592 7 7 2 61893 67852
0 31593 7 2 2 82666 98379
0 31594 5 1 1 98386
0 31595 7 3 2 82745 92548
0 31596 5 1 1 98388
0 31597 7 1 2 31594 31596
0 31598 5 9 1 31597
0 31599 7 1 2 61356 98391
0 31600 5 1 1 31599
0 31601 7 7 2 61894 63003
0 31602 7 4 2 66221 98400
0 31603 7 2 2 82667 98407
0 31604 5 1 1 98411
0 31605 7 1 2 31600 31604
0 31606 5 7 1 31605
0 31607 7 6 2 69215 93849
0 31608 7 2 2 64958 98361
0 31609 5 1 1 98426
0 31610 7 1 2 74811 85358
0 31611 7 2 2 97443 31610
0 31612 5 1 1 98428
0 31613 7 1 2 62589 98429
0 31614 5 1 1 31613
0 31615 7 1 2 31609 31614
0 31616 5 2 1 31615
0 31617 7 1 2 98420 98430
0 31618 5 1 1 31617
0 31619 7 2 2 74812 87715
0 31620 7 7 2 62859 62961
0 31621 7 1 2 88143 98434
0 31622 7 1 2 98432 31621
0 31623 5 1 1 31622
0 31624 7 1 2 31618 31623
0 31625 5 1 1 31624
0 31626 7 1 2 62136 31625
0 31627 5 1 1 31626
0 31628 7 2 2 68670 93659
0 31629 7 3 2 69818 72455
0 31630 7 1 2 86650 98435
0 31631 7 1 2 98443 31630
0 31632 7 2 2 98441 31631
0 31633 5 1 1 98446
0 31634 7 1 2 61274 98447
0 31635 5 1 1 31634
0 31636 7 1 2 31627 31635
0 31637 5 1 1 31636
0 31638 7 1 2 98413 31637
0 31639 5 1 1 31638
0 31640 7 5 2 62962 67853
0 31641 7 4 2 81820 98448
0 31642 7 1 2 82512 98453
0 31643 5 1 1 31642
0 31644 7 1 2 93073 98100
0 31645 7 1 2 90746 31644
0 31646 5 1 1 31645
0 31647 7 1 2 31643 31646
0 31648 5 2 1 31647
0 31649 7 1 2 77012 98457
0 31650 5 1 1 31649
0 31651 7 1 2 78847 98454
0 31652 7 1 2 77644 31651
0 31653 5 1 1 31652
0 31654 7 1 2 31650 31653
0 31655 5 1 1 31654
0 31656 7 1 2 66222 31655
0 31657 5 1 1 31656
0 31658 7 1 2 88226 92849
0 31659 5 1 1 31658
0 31660 7 1 2 63004 87543
0 31661 5 1 1 31660
0 31662 7 1 2 31659 31661
0 31663 5 5 1 31662
0 31664 7 2 2 61357 98459
0 31665 5 1 1 98464
0 31666 7 1 2 67785 77013
0 31667 7 1 2 98465 31666
0 31668 5 1 1 31667
0 31669 7 1 2 31657 31668
0 31670 5 1 1 31669
0 31671 7 1 2 73624 31670
0 31672 5 1 1 31671
0 31673 7 1 2 90836 31612
0 31674 5 1 1 31673
0 31675 7 2 2 66223 97339
0 31676 7 12 2 67854 68022
0 31677 7 1 2 88670 98468
0 31678 7 1 2 98466 31677
0 31679 7 1 2 31674 31678
0 31680 5 1 1 31679
0 31681 7 1 2 31672 31680
0 31682 5 1 1 31681
0 31683 7 1 2 61275 31682
0 31684 5 1 1 31683
0 31685 7 3 2 90588 98101
0 31686 7 1 2 93029 98480
0 31687 5 1 1 31686
0 31688 7 1 2 31665 31687
0 31689 5 2 1 31688
0 31690 7 1 2 80382 93846
0 31691 7 1 2 77014 31690
0 31692 7 1 2 98483 31691
0 31693 5 1 1 31692
0 31694 7 1 2 31684 31693
0 31695 5 1 1 31694
0 31696 7 1 2 62590 31695
0 31697 5 1 1 31696
0 31698 7 2 2 75484 91368
0 31699 7 3 2 81587 98469
0 31700 7 3 2 62423 62963
0 31701 7 1 2 98487 98490
0 31702 7 1 2 98485 31701
0 31703 7 1 2 77779 31702
0 31704 5 1 1 31703
0 31705 7 1 2 31697 31704
0 31706 5 1 1 31705
0 31707 7 1 2 69216 31706
0 31708 5 1 1 31707
0 31709 7 1 2 31639 31708
0 31710 7 1 2 31591 31709
0 31711 5 1 1 31710
0 31712 7 1 2 64260 31711
0 31713 5 1 1 31712
0 31714 7 1 2 78857 16797
0 31715 5 1 1 31714
0 31716 7 6 2 66757 67855
0 31717 5 1 1 98493
0 31718 7 1 2 1005 31717
0 31719 7 2 2 31715 31718
0 31720 7 1 2 61358 98499
0 31721 5 1 1 31720
0 31722 7 1 2 80508 98408
0 31723 5 1 1 31722
0 31724 7 1 2 31721 31723
0 31725 5 1 1 31724
0 31726 7 1 2 67786 31725
0 31727 5 1 1 31726
0 31728 7 4 2 67856 78714
0 31729 7 1 2 98501 98467
0 31730 5 1 1 31729
0 31731 7 1 2 31727 31730
0 31732 5 1 1 31731
0 31733 7 1 2 66107 31732
0 31734 5 1 1 31733
0 31735 7 4 2 67787 84422
0 31736 7 1 2 66224 98502
0 31737 7 1 2 98505 31736
0 31738 5 1 1 31737
0 31739 7 1 2 31734 31738
0 31740 5 1 1 31739
0 31741 7 5 2 69109 97415
0 31742 7 1 2 79867 92706
0 31743 5 1 1 31742
0 31744 7 2 2 63357 75156
0 31745 7 1 2 79918 98514
0 31746 5 1 1 31745
0 31747 7 1 2 31743 31746
0 31748 5 1 1 31747
0 31749 7 1 2 63814 31748
0 31750 5 1 1 31749
0 31751 7 1 2 19998 97005
0 31752 5 2 1 31751
0 31753 7 1 2 98515 98516
0 31754 5 1 1 31753
0 31755 7 1 2 31750 31754
0 31756 5 1 1 31755
0 31757 7 1 2 98509 31756
0 31758 7 1 2 31740 31757
0 31759 5 1 1 31758
0 31760 7 1 2 31713 31759
0 31761 5 1 1 31760
0 31762 7 1 2 69378 31761
0 31763 5 1 1 31762
0 31764 7 1 2 84115 97304
0 31765 5 1 1 31764
0 31766 7 15 2 61276 97643
0 31767 5 2 1 98518
0 31768 7 1 2 74657 98519
0 31769 5 1 1 31768
0 31770 7 1 2 31765 31769
0 31771 5 1 1 31770
0 31772 7 1 2 71971 31771
0 31773 5 1 1 31772
0 31774 7 7 2 70378 75802
0 31775 7 1 2 63815 98535
0 31776 5 1 1 31775
0 31777 7 1 2 82214 31776
0 31778 5 1 1 31777
0 31779 7 1 2 96957 31778
0 31780 5 1 1 31779
0 31781 7 1 2 31773 31780
0 31782 5 1 1 31781
0 31783 7 1 2 85568 31782
0 31784 5 1 1 31783
0 31785 7 2 2 61277 98151
0 31786 7 1 2 98344 98542
0 31787 5 1 1 31786
0 31788 7 1 2 31784 31787
0 31789 5 1 1 31788
0 31790 7 6 2 63005 82668
0 31791 7 1 2 61895 64361
0 31792 7 2 2 98544 31791
0 31793 5 1 1 98550
0 31794 7 1 2 61359 98551
0 31795 7 1 2 31789 31794
0 31796 5 1 1 31795
0 31797 7 2 2 66225 98392
0 31798 5 1 1 98552
0 31799 7 4 2 81657 93683
0 31800 7 3 2 61360 98554
0 31801 5 1 1 98558
0 31802 7 1 2 31798 31801
0 31803 5 5 1 31802
0 31804 7 3 2 93850 94361
0 31805 7 1 2 85569 98566
0 31806 7 1 2 95416 31805
0 31807 5 1 1 31806
0 31808 7 3 2 98152 97525
0 31809 7 7 2 61278 66994
0 31810 7 1 2 75516 89924
0 31811 7 1 2 98572 31810
0 31812 7 1 2 98569 31811
0 31813 5 1 1 31812
0 31814 7 1 2 31807 31813
0 31815 5 1 1 31814
0 31816 7 1 2 98561 31815
0 31817 5 1 1 31816
0 31818 7 2 2 64362 70379
0 31819 7 6 2 69110 98579
0 31820 7 2 2 82719 98581
0 31821 7 1 2 85598 98470
0 31822 7 1 2 98587 31821
0 31823 5 1 1 31822
0 31824 7 4 2 69217 73071
0 31825 7 4 2 63006 63816
0 31826 7 2 2 95148 98593
0 31827 7 1 2 98589 98597
0 31828 7 1 2 89665 31827
0 31829 5 1 1 31828
0 31830 7 1 2 31823 31829
0 31831 5 1 1 31830
0 31832 7 1 2 61361 31831
0 31833 5 1 1 31832
0 31834 7 5 2 66226 67278
0 31835 7 1 2 75485 92549
0 31836 7 1 2 98599 31835
0 31837 7 1 2 98588 31836
0 31838 5 1 1 31837
0 31839 7 1 2 31833 31838
0 31840 5 1 1 31839
0 31841 7 1 2 93851 31840
0 31842 5 1 1 31841
0 31843 7 1 2 31817 31842
0 31844 7 1 2 31796 31843
0 31845 5 1 1 31844
0 31846 7 1 2 69819 82278
0 31847 7 1 2 31845 31846
0 31848 5 1 1 31847
0 31849 7 1 2 64753 31848
0 31850 7 1 2 31763 31849
0 31851 5 1 1 31850
0 31852 7 2 2 63358 98347
0 31853 5 1 1 98604
0 31854 7 1 2 62137 94841
0 31855 5 2 1 31854
0 31856 7 1 2 31853 98606
0 31857 5 2 1 31856
0 31858 7 4 2 97980 97416
0 31859 7 1 2 98608 98610
0 31860 5 1 1 31859
0 31861 7 3 2 68198 64261
0 31862 7 1 2 80284 98614
0 31863 7 1 2 97526 31862
0 31864 7 1 2 86527 31863
0 31865 5 1 1 31864
0 31866 7 1 2 31860 31865
0 31867 5 1 1 31866
0 31868 7 1 2 66108 31867
0 31869 5 1 1 31868
0 31870 7 10 2 62138 67788
0 31871 7 1 2 96830 98617
0 31872 7 1 2 86074 31871
0 31873 5 1 1 31872
0 31874 7 5 2 62964 63359
0 31875 7 1 2 73919 97417
0 31876 7 1 2 98627 31875
0 31877 5 1 1 31876
0 31878 7 1 2 31873 31877
0 31879 5 1 1 31878
0 31880 7 1 2 70380 97706
0 31881 7 1 2 31879 31880
0 31882 5 1 1 31881
0 31883 7 1 2 31869 31882
0 31884 5 1 1 31883
0 31885 7 1 2 63975 31884
0 31886 5 1 1 31885
0 31887 7 1 2 78395 87298
0 31888 5 2 1 31887
0 31889 7 1 2 94188 98632
0 31890 5 1 1 31889
0 31891 7 4 2 62139 64262
0 31892 7 1 2 98634 98421
0 31893 7 1 2 31890 31892
0 31894 5 1 1 31893
0 31895 7 1 2 31886 31894
0 31896 5 1 1 31895
0 31897 7 1 2 62591 31896
0 31898 5 1 1 31897
0 31899 7 2 2 76709 98628
0 31900 7 1 2 98638 98433
0 31901 5 1 1 31900
0 31902 7 3 2 63579 71586
0 31903 5 1 1 98640
0 31904 7 1 2 90933 98641
0 31905 7 1 2 98422 31904
0 31906 5 1 1 31905
0 31907 7 1 2 31901 31906
0 31908 5 1 1 31907
0 31909 7 1 2 98635 31908
0 31910 5 1 1 31909
0 31911 7 1 2 31898 31910
0 31912 5 1 1 31911
0 31913 7 8 2 62860 69379
0 31914 7 1 2 93772 98643
0 31915 7 1 2 31912 31914
0 31916 5 1 1 31915
0 31917 7 11 2 91340 97707
0 31918 5 2 1 98651
0 31919 7 2 2 86631 98652
0 31920 5 1 1 98664
0 31921 7 1 2 95390 98653
0 31922 5 1 1 31921
0 31923 7 11 2 69111 92472
0 31924 7 1 2 75192 98666
0 31925 5 1 1 31924
0 31926 7 1 2 31922 31925
0 31927 5 1 1 31926
0 31928 7 1 2 85570 31927
0 31929 5 1 1 31928
0 31930 7 1 2 31920 31929
0 31931 5 1 1 31930
0 31932 7 1 2 64363 31931
0 31933 5 1 1 31932
0 31934 7 12 2 64263 91021
0 31935 5 1 1 98677
0 31936 7 2 2 86614 75517
0 31937 7 1 2 87832 98689
0 31938 7 1 2 98678 31937
0 31939 5 1 1 31938
0 31940 7 1 2 31933 31939
0 31941 5 1 1 31940
0 31942 7 1 2 87209 93735
0 31943 7 1 2 31941 31942
0 31944 5 1 1 31943
0 31945 7 1 2 31916 31944
0 31946 5 1 1 31945
0 31947 7 1 2 87253 31946
0 31948 5 1 1 31947
0 31949 7 1 2 81457 85571
0 31950 5 1 1 31949
0 31951 7 1 2 61896 95886
0 31952 5 1 1 31951
0 31953 7 1 2 31950 31952
0 31954 5 1 1 31953
0 31955 7 1 2 86678 98007
0 31956 5 1 1 31955
0 31957 7 2 2 63817 75803
0 31958 7 1 2 97663 98691
0 31959 5 1 1 31958
0 31960 7 1 2 31956 31959
0 31961 5 1 1 31960
0 31962 7 1 2 61279 31961
0 31963 5 1 1 31962
0 31964 7 1 2 86679 97880
0 31965 5 1 1 31964
0 31966 7 1 2 31963 31965
0 31967 5 1 1 31966
0 31968 7 1 2 70381 31967
0 31969 5 1 1 31968
0 31970 7 4 2 62965 94664
0 31971 7 5 2 63007 63580
0 31972 7 1 2 61280 98697
0 31973 7 1 2 98218 31972
0 31974 7 1 2 98693 31973
0 31975 5 1 1 31974
0 31976 7 1 2 31969 31975
0 31977 5 1 1 31976
0 31978 7 1 2 31954 31977
0 31979 5 1 1 31978
0 31980 7 2 2 75157 92473
0 31981 7 1 2 69112 95042
0 31982 7 1 2 89779 31981
0 31983 7 1 2 85231 31982
0 31984 7 1 2 98702 31983
0 31985 5 1 1 31984
0 31986 7 1 2 31979 31985
0 31987 5 1 1 31986
0 31988 7 3 2 64959 92216
0 31989 7 1 2 80141 98704
0 31990 7 1 2 31987 31989
0 31991 5 1 1 31990
0 31992 7 1 2 69587 31991
0 31993 7 1 2 31948 31992
0 31994 5 1 1 31993
0 31995 7 1 2 31851 31994
0 31996 5 1 1 31995
0 31997 7 1 2 61613 31996
0 31998 5 1 1 31997
0 31999 7 4 2 91341 98153
0 32000 5 1 1 98707
0 32001 7 1 2 83124 98708
0 32002 5 1 1 32001
0 32003 7 4 2 67857 63976
0 32004 7 3 2 69113 93067
0 32005 7 2 2 98711 98715
0 32006 7 1 2 83416 90876
0 32007 7 1 2 98718 32006
0 32008 5 1 1 32007
0 32009 7 1 2 32002 32008
0 32010 5 1 1 32009
0 32011 7 1 2 76005 32010
0 32012 5 1 1 32011
0 32013 7 2 2 66227 69820
0 32014 7 1 2 85174 98720
0 32015 7 5 2 67789 98471
0 32016 7 1 2 95542 98722
0 32017 7 1 2 32014 32016
0 32018 5 1 1 32017
0 32019 7 1 2 32012 32018
0 32020 5 1 1 32019
0 32021 7 1 2 66995 32020
0 32022 5 1 1 32021
0 32023 7 2 2 69114 77304
0 32024 7 6 2 66228 62592
0 32025 7 1 2 88671 91861
0 32026 7 1 2 98729 32025
0 32027 7 1 2 98727 32026
0 32028 7 1 2 87254 32027
0 32029 5 1 1 32028
0 32030 7 1 2 32022 32029
0 32031 5 1 1 32030
0 32032 7 1 2 62424 32031
0 32033 5 1 1 32032
0 32034 7 5 2 64264 88164
0 32035 7 3 2 98102 98735
0 32036 7 2 2 84486 98740
0 32037 7 5 2 67479 75804
0 32038 5 1 1 98745
0 32039 7 1 2 68861 98746
0 32040 5 1 1 32039
0 32041 7 1 2 3634 32040
0 32042 5 2 1 32041
0 32043 7 1 2 70382 98750
0 32044 7 1 2 98743 32043
0 32045 5 1 1 32044
0 32046 7 1 2 32033 32045
0 32047 5 1 1 32046
0 32048 7 1 2 63818 32047
0 32049 5 1 1 32048
0 32050 7 1 2 31491 98744
0 32051 5 1 1 32050
0 32052 7 1 2 32049 32051
0 32053 5 1 1 32052
0 32054 7 1 2 64754 32053
0 32055 5 1 1 32054
0 32056 7 1 2 62425 75919
0 32057 5 3 1 32056
0 32058 7 1 2 62140 85033
0 32059 5 2 1 32058
0 32060 7 1 2 98752 98755
0 32061 5 1 1 32060
0 32062 7 3 2 61362 92550
0 32063 7 1 2 78848 98757
0 32064 7 1 2 32061 32063
0 32065 5 1 1 32064
0 32066 7 1 2 93655 98756
0 32067 5 1 1 32066
0 32068 7 1 2 82002 98367
0 32069 7 1 2 32067 32068
0 32070 5 1 1 32069
0 32071 7 1 2 32065 32070
0 32072 5 1 1 32071
0 32073 7 1 2 63360 32072
0 32074 5 1 1 32073
0 32075 7 3 2 62426 63008
0 32076 7 2 2 61363 98760
0 32077 7 1 2 88747 76861
0 32078 7 1 2 98763 32077
0 32079 5 1 1 32078
0 32080 7 1 2 32074 32079
0 32081 5 1 1 32080
0 32082 7 1 2 86926 98694
0 32083 7 1 2 32081 32082
0 32084 5 1 1 32083
0 32085 7 1 2 32055 32084
0 32086 5 1 1 32085
0 32087 7 1 2 65784 32086
0 32088 5 1 1 32087
0 32089 7 2 2 83125 73465
0 32090 7 1 2 98199 98491
0 32091 7 1 2 80512 32090
0 32092 7 1 2 98598 32091
0 32093 7 1 2 98765 32092
0 32094 5 1 1 32093
0 32095 7 1 2 32088 32094
0 32096 5 1 1 32095
0 32097 7 1 2 64364 32096
0 32098 5 1 1 32097
0 32099 7 1 2 68199 98362
0 32100 5 1 1 32099
0 32101 7 1 2 86575 79695
0 32102 7 1 2 91233 32101
0 32103 5 1 1 32102
0 32104 7 1 2 32100 32103
0 32105 5 1 1 32104
0 32106 7 6 2 69588 93773
0 32107 7 2 2 95149 97581
0 32108 7 1 2 74159 96070
0 32109 7 1 2 98773 32108
0 32110 7 1 2 98767 32109
0 32111 7 1 2 32105 32110
0 32112 5 1 1 32111
0 32113 7 1 2 32098 32112
0 32114 5 1 1 32113
0 32115 7 1 2 61281 32114
0 32116 5 1 1 32115
0 32117 7 1 2 2022 93766
0 32118 5 1 1 32117
0 32119 7 1 2 81480 90633
0 32120 5 1 1 32119
0 32121 7 2 2 32118 32120
0 32122 7 1 2 83060 98775
0 32123 5 1 1 32122
0 32124 7 3 2 63009 63361
0 32125 7 1 2 64755 91809
0 32126 7 2 2 98777 32125
0 32127 7 1 2 68023 98780
0 32128 5 1 1 32127
0 32129 7 1 2 32123 32128
0 32130 5 1 1 32129
0 32131 7 2 2 62593 88035
0 32132 5 1 1 98782
0 32133 7 1 2 31903 32132
0 32134 5 1 1 32133
0 32135 7 1 2 81195 32134
0 32136 7 1 2 32130 32135
0 32137 5 1 1 32136
0 32138 7 1 2 74327 76006
0 32139 7 1 2 71587 90600
0 32140 7 1 2 32138 32139
0 32141 7 1 2 94692 32140
0 32142 5 1 1 32141
0 32143 7 1 2 32137 32142
0 32144 5 1 1 32143
0 32145 7 1 2 71847 32144
0 32146 5 1 1 32145
0 32147 7 2 2 80383 81588
0 32148 5 1 1 98784
0 32149 7 1 2 78970 90601
0 32150 7 1 2 98785 32149
0 32151 5 1 1 32150
0 32152 7 1 2 98633 32148
0 32153 5 2 1 32152
0 32154 7 1 2 63179 98768
0 32155 7 1 2 98786 32154
0 32156 5 1 1 32155
0 32157 7 1 2 32151 32156
0 32158 5 1 1 32157
0 32159 7 1 2 74240 32158
0 32160 5 1 1 32159
0 32161 7 1 2 67279 86163
0 32162 7 1 2 90602 32161
0 32163 7 1 2 87521 78396
0 32164 7 1 2 32162 32163
0 32165 5 1 1 32164
0 32166 7 1 2 32160 32165
0 32167 5 1 1 32166
0 32168 7 1 2 61897 32167
0 32169 5 1 1 32168
0 32170 7 2 2 83519 83780
0 32171 7 1 2 91610 98788
0 32172 5 1 1 32171
0 32173 7 2 2 67280 80852
0 32174 7 1 2 76710 83182
0 32175 7 1 2 98790 32174
0 32176 5 1 1 32175
0 32177 7 1 2 32172 32176
0 32178 5 2 1 32177
0 32179 7 1 2 98781 98792
0 32180 5 1 1 32179
0 32181 7 1 2 32169 32180
0 32182 5 1 1 32181
0 32183 7 1 2 75855 32182
0 32184 5 1 1 32183
0 32185 7 1 2 32146 32184
0 32186 5 1 1 32185
0 32187 7 1 2 64265 98373
0 32188 7 1 2 32186 32187
0 32189 5 1 1 32188
0 32190 7 1 2 32116 32189
0 32191 5 1 1 32190
0 32192 7 1 2 69380 32191
0 32193 5 1 1 32192
0 32194 7 2 2 71588 97609
0 32195 5 1 1 98794
0 32196 7 5 2 97626 97418
0 32197 7 2 2 73333 98796
0 32198 5 2 1 98801
0 32199 7 2 2 32195 98803
0 32200 5 6 1 98805
0 32201 7 1 2 65448 98807
0 32202 5 1 1 32201
0 32203 7 2 2 79908 98797
0 32204 5 1 1 98813
0 32205 7 1 2 70383 98814
0 32206 5 2 1 32205
0 32207 7 1 2 32202 98815
0 32208 5 1 1 32207
0 32209 7 1 2 68671 32208
0 32210 5 1 1 32209
0 32211 7 2 2 94474 98798
0 32212 5 1 1 98817
0 32213 7 1 2 32210 32212
0 32214 5 1 1 32213
0 32215 7 1 2 76017 32214
0 32216 5 1 1 32215
0 32217 7 1 2 75930 89791
0 32218 7 2 2 97274 32217
0 32219 5 2 1 98819
0 32220 7 1 2 97006 98820
0 32221 5 2 1 32220
0 32222 7 2 2 65785 98823
0 32223 7 4 2 66109 61898
0 32224 7 1 2 75353 94362
0 32225 7 1 2 98827 32224
0 32226 7 1 2 98825 32225
0 32227 5 1 1 32226
0 32228 7 1 2 32216 32227
0 32229 5 1 1 32228
0 32230 7 1 2 64756 32229
0 32231 5 1 1 32230
0 32232 7 3 2 66110 68024
0 32233 7 1 2 77800 94363
0 32234 7 1 2 98831 32233
0 32235 7 1 2 79103 92739
0 32236 7 1 2 32234 32235
0 32237 5 1 1 32236
0 32238 7 1 2 32231 32237
0 32239 5 1 1 32238
0 32240 7 1 2 69381 32239
0 32241 5 1 1 32240
0 32242 7 1 2 66111 76764
0 32243 7 1 2 80853 32242
0 32244 7 3 2 67707 69115
0 32245 7 2 2 92217 98834
0 32246 7 1 2 85862 98837
0 32247 7 1 2 32243 32246
0 32248 5 1 1 32247
0 32249 7 1 2 32241 32248
0 32250 5 1 1 32249
0 32251 7 1 2 63362 32250
0 32252 5 1 1 32251
0 32253 7 2 2 78478 92863
0 32254 7 1 2 88690 90064
0 32255 7 1 2 97610 32254
0 32256 7 1 2 98839 32255
0 32257 5 1 1 32256
0 32258 7 1 2 32252 32257
0 32259 5 1 1 32258
0 32260 7 1 2 75158 32259
0 32261 5 1 1 32260
0 32262 7 1 2 64960 95330
0 32263 5 1 1 32262
0 32264 7 1 2 10972 32263
0 32265 5 1 1 32264
0 32266 7 1 2 71589 32265
0 32267 5 1 1 32266
0 32268 7 1 2 74244 98783
0 32269 5 1 1 32268
0 32270 7 1 2 32267 32269
0 32271 5 1 1 32270
0 32272 7 1 2 71848 32271
0 32273 5 1 1 32272
0 32274 7 1 2 75856 98793
0 32275 5 1 1 32274
0 32276 7 1 2 32273 32275
0 32277 5 1 1 32276
0 32278 7 1 2 83126 97735
0 32279 7 1 2 32277 32278
0 32280 5 1 1 32279
0 32281 7 1 2 77616 72385
0 32282 7 4 2 63819 64365
0 32283 7 1 2 97627 98841
0 32284 7 1 2 32281 32283
0 32285 7 1 2 97183 32284
0 32286 5 1 1 32285
0 32287 7 1 2 32280 32286
0 32288 5 1 1 32287
0 32289 7 1 2 79449 32288
0 32290 5 1 1 32289
0 32291 7 3 2 63820 64266
0 32292 7 1 2 89663 98845
0 32293 7 3 2 61282 73072
0 32294 7 1 2 96075 96842
0 32295 7 1 2 98848 32294
0 32296 7 1 2 32292 32295
0 32297 5 1 1 32296
0 32298 7 1 2 32290 32297
0 32299 7 1 2 32261 32298
0 32300 5 1 1 32299
0 32301 7 1 2 90708 32300
0 32302 5 1 1 32301
0 32303 7 2 2 67858 64757
0 32304 7 2 2 91369 98851
0 32305 7 1 2 95608 98853
0 32306 5 1 1 32305
0 32307 7 1 2 90032 83706
0 32308 7 1 2 98769 32307
0 32309 5 1 1 32308
0 32310 7 1 2 32306 32309
0 32311 5 1 1 32310
0 32312 7 1 2 65449 32311
0 32313 5 1 1 32312
0 32314 7 3 2 91370 98472
0 32315 7 1 2 88098 79909
0 32316 7 1 2 98855 32315
0 32317 5 1 1 32316
0 32318 7 1 2 32313 32317
0 32319 5 1 1 32318
0 32320 7 1 2 82003 32319
0 32321 5 1 1 32320
0 32322 7 1 2 86927 80444
0 32323 5 1 1 32322
0 32324 7 1 2 90478 81071
0 32325 5 1 1 32324
0 32326 7 1 2 32323 32325
0 32327 5 1 1 32326
0 32328 7 1 2 65450 32327
0 32329 5 1 1 32328
0 32330 7 1 2 78889 94429
0 32331 5 1 1 32330
0 32332 7 1 2 32329 32331
0 32333 5 1 1 32332
0 32334 7 1 2 78849 97598
0 32335 7 1 2 32333 32334
0 32336 5 1 1 32335
0 32337 7 1 2 32321 32336
0 32338 5 1 1 32337
0 32339 7 1 2 68672 32338
0 32340 5 1 1 32339
0 32341 7 1 2 87255 98854
0 32342 7 1 2 94475 32341
0 32343 5 1 1 32342
0 32344 7 1 2 32340 32343
0 32345 5 1 1 32344
0 32346 7 1 2 98611 32345
0 32347 5 1 1 32346
0 32348 7 2 2 94667 98840
0 32349 7 1 2 76675 91006
0 32350 7 1 2 98858 32349
0 32351 5 1 1 32350
0 32352 7 1 2 32347 32351
0 32353 5 1 1 32352
0 32354 7 1 2 63363 32353
0 32355 5 1 1 32354
0 32356 7 1 2 90065 91007
0 32357 7 1 2 98859 32356
0 32358 5 1 1 32357
0 32359 7 1 2 32355 32358
0 32360 5 1 1 32359
0 32361 7 1 2 69382 32360
0 32362 5 1 1 32361
0 32363 7 1 2 87210 76432
0 32364 7 1 2 92956 93030
0 32365 7 1 2 32363 32364
0 32366 7 2 2 92850 94364
0 32367 7 1 2 87270 98860
0 32368 7 1 2 32365 32367
0 32369 5 1 1 32368
0 32370 7 1 2 32362 32369
0 32371 5 1 1 32370
0 32372 7 1 2 75159 32371
0 32373 5 1 1 32372
0 32374 7 2 2 61283 93164
0 32375 7 1 2 92080 98862
0 32376 5 1 1 32375
0 32377 7 2 2 81872 87833
0 32378 5 1 1 98864
0 32379 7 1 2 87763 32378
0 32380 5 4 1 32379
0 32381 7 1 2 86632 98866
0 32382 5 1 1 32381
0 32383 7 1 2 32376 32382
0 32384 5 1 1 32383
0 32385 7 1 2 74924 32384
0 32386 5 1 1 32385
0 32387 7 1 2 71249 98692
0 32388 5 1 1 32387
0 32389 7 1 2 85672 32388
0 32390 5 1 1 32389
0 32391 7 1 2 70384 32390
0 32392 5 1 1 32391
0 32393 7 1 2 67281 85692
0 32394 7 1 2 84974 32393
0 32395 5 1 1 32394
0 32396 7 1 2 32392 32395
0 32397 5 1 1 32396
0 32398 7 2 2 65786 32397
0 32399 7 1 2 87716 98870
0 32400 5 1 1 32399
0 32401 7 1 2 32386 32400
0 32402 5 1 1 32401
0 32403 7 5 2 88165 98401
0 32404 7 2 2 94731 98872
0 32405 7 1 2 89887 98877
0 32406 7 1 2 32402 32405
0 32407 5 1 1 32406
0 32408 7 1 2 66511 32407
0 32409 7 1 2 32373 32408
0 32410 7 1 2 32302 32409
0 32411 7 1 2 32193 32410
0 32412 5 1 1 32411
0 32413 7 1 2 65171 32412
0 32414 7 1 2 31998 32413
0 32415 5 1 1 32414
0 32416 7 21 2 64366 97628
0 32417 7 1 2 76053 77015
0 32418 5 1 1 32417
0 32419 7 1 2 26660 32418
0 32420 5 1 1 32419
0 32421 7 1 2 68200 32420
0 32422 5 1 1 32421
0 32423 7 1 2 76561 95830
0 32424 5 1 1 32423
0 32425 7 1 2 32422 32424
0 32426 5 1 1 32425
0 32427 7 1 2 86446 32426
0 32428 5 1 1 32427
0 32429 7 1 2 11993 15239
0 32430 5 2 1 32429
0 32431 7 1 2 86377 83183
0 32432 7 1 2 98900 32431
0 32433 5 1 1 32432
0 32434 7 1 2 32428 32433
0 32435 5 1 1 32434
0 32436 7 1 2 65787 32435
0 32437 5 1 1 32436
0 32438 7 3 2 70385 87166
0 32439 7 1 2 61614 83061
0 32440 7 1 2 80092 32439
0 32441 7 1 2 98902 32440
0 32442 5 1 1 32441
0 32443 7 1 2 32437 32442
0 32444 5 1 1 32443
0 32445 7 1 2 98879 32444
0 32446 5 1 1 32445
0 32447 7 1 2 92864 98901
0 32448 5 1 1 32447
0 32449 7 1 2 83693 85871
0 32450 5 1 1 32449
0 32451 7 1 2 32448 32450
0 32452 5 1 1 32451
0 32453 7 1 2 96449 97708
0 32454 7 1 2 32452 32453
0 32455 5 1 1 32454
0 32456 7 1 2 32446 32455
0 32457 5 1 1 32456
0 32458 7 1 2 68673 32457
0 32459 5 1 1 32458
0 32460 7 2 2 63180 82093
0 32461 7 2 2 90377 98510
0 32462 7 1 2 98905 98907
0 32463 5 1 1 32462
0 32464 7 4 2 64267 87834
0 32465 7 2 2 77560 98909
0 32466 7 1 2 61284 76170
0 32467 7 1 2 98913 32466
0 32468 5 1 1 32467
0 32469 7 1 2 32463 32468
0 32470 5 1 1 32469
0 32471 7 1 2 71250 32470
0 32472 5 1 1 32471
0 32473 7 5 2 64367 76711
0 32474 7 2 2 98179 98915
0 32475 7 1 2 89597 82094
0 32476 7 1 2 98920 32475
0 32477 5 1 1 32476
0 32478 7 1 2 32472 32477
0 32479 5 1 1 32478
0 32480 7 1 2 83127 32479
0 32481 5 1 1 32480
0 32482 7 1 2 92029 98818
0 32483 5 1 1 32482
0 32484 7 1 2 32481 32483
0 32485 5 1 1 32484
0 32486 7 1 2 64961 32485
0 32487 5 1 1 32486
0 32488 7 1 2 32459 32487
0 32489 5 1 1 32488
0 32490 7 1 2 69383 32489
0 32491 5 1 1 32490
0 32492 7 1 2 61285 61615
0 32493 7 2 2 93903 32492
0 32494 7 1 2 75710 89888
0 32495 7 1 2 98922 32494
0 32496 7 1 2 85481 32495
0 32497 5 1 1 32496
0 32498 7 1 2 32491 32497
0 32499 5 1 1 32498
0 32500 7 1 2 64758 32499
0 32501 5 1 1 32500
0 32502 7 1 2 87680 97378
0 32503 7 1 2 98835 32502
0 32504 7 1 2 89394 32503
0 32505 7 1 2 92237 32504
0 32506 5 1 1 32505
0 32507 7 1 2 64962 80791
0 32508 7 1 2 98766 32507
0 32509 5 1 1 32508
0 32510 7 1 2 68862 81419
0 32511 7 1 2 96488 32510
0 32512 5 1 1 32511
0 32513 7 1 2 32509 32512
0 32514 5 1 1 32513
0 32515 7 1 2 94335 97611
0 32516 7 1 2 32514 32515
0 32517 5 1 1 32516
0 32518 7 1 2 32506 32517
0 32519 5 1 1 32518
0 32520 7 1 2 81491 32519
0 32521 5 1 1 32520
0 32522 7 1 2 32501 32521
0 32523 5 1 1 32522
0 32524 7 1 2 68426 32523
0 32525 5 1 1 32524
0 32526 7 1 2 88785 97941
0 32527 7 1 2 98880 32526
0 32528 5 1 1 32527
0 32529 7 1 2 81821 82606
0 32530 7 1 2 98808 32529
0 32531 5 1 1 32530
0 32532 7 1 2 32528 32531
0 32533 5 1 1 32532
0 32534 7 1 2 86965 32533
0 32535 5 1 1 32534
0 32536 7 2 2 66112 95425
0 32537 7 2 2 88468 98924
0 32538 7 1 2 75254 73466
0 32539 7 1 2 93478 32538
0 32540 7 1 2 98926 32539
0 32541 5 1 1 32540
0 32542 7 1 2 32535 32541
0 32543 5 1 1 32542
0 32544 7 1 2 87394 32543
0 32545 5 1 1 32544
0 32546 7 3 2 79450 93366
0 32547 7 1 2 98802 98928
0 32548 5 1 1 32547
0 32549 7 1 2 64533 88192
0 32550 7 1 2 98809 32549
0 32551 5 1 1 32550
0 32552 7 1 2 32548 32551
0 32553 5 1 1 32552
0 32554 7 1 2 71849 83520
0 32555 7 1 2 32553 32554
0 32556 5 1 1 32555
0 32557 7 1 2 81092 81883
0 32558 7 2 2 73073 72704
0 32559 7 1 2 97612 98931
0 32560 7 1 2 32557 32559
0 32561 5 1 1 32560
0 32562 7 1 2 32556 32561
0 32563 5 1 1 32562
0 32564 7 1 2 83128 32563
0 32565 5 1 1 32564
0 32566 7 1 2 75274 91460
0 32567 7 2 2 82004 88123
0 32568 7 1 2 96843 98933
0 32569 7 1 2 97736 32568
0 32570 7 1 2 32566 32569
0 32571 5 1 1 32570
0 32572 7 1 2 32565 32571
0 32573 7 1 2 32545 32572
0 32574 7 1 2 32525 32573
0 32575 5 1 1 32574
0 32576 7 1 2 66996 32575
0 32577 5 1 1 32576
0 32578 7 6 2 81707 94365
0 32579 7 1 2 91772 94211
0 32580 5 1 1 32579
0 32581 7 1 2 87325 91635
0 32582 5 1 1 32581
0 32583 7 1 2 32580 32582
0 32584 5 1 1 32583
0 32585 7 1 2 73334 32584
0 32586 5 1 1 32585
0 32587 7 2 2 83955 94555
0 32588 5 1 1 98941
0 32589 7 1 2 63581 98942
0 32590 5 1 1 32589
0 32591 7 1 2 32586 32590
0 32592 5 1 1 32591
0 32593 7 1 2 68025 32592
0 32594 5 1 1 32593
0 32595 7 1 2 66512 90479
0 32596 7 1 2 74050 32595
0 32597 7 1 2 85664 32596
0 32598 5 1 1 32597
0 32599 7 1 2 32594 32598
0 32600 5 1 1 32599
0 32601 7 1 2 83129 32600
0 32602 5 1 1 32601
0 32603 7 1 2 82645 95474
0 32604 5 1 1 32603
0 32605 7 1 2 88233 88538
0 32606 5 1 1 32605
0 32607 7 1 2 32604 32606
0 32608 5 1 1 32607
0 32609 7 1 2 83816 83665
0 32610 7 1 2 32608 32609
0 32611 5 1 1 32610
0 32612 7 1 2 32602 32611
0 32613 5 1 1 32612
0 32614 7 1 2 65788 32613
0 32615 5 1 1 32614
0 32616 7 1 2 78518 76372
0 32617 7 1 2 82991 32616
0 32618 7 1 2 96844 32617
0 32619 7 1 2 91435 32618
0 32620 5 1 1 32619
0 32621 7 1 2 32615 32620
0 32622 5 1 1 32621
0 32623 7 1 2 69821 32622
0 32624 5 1 1 32623
0 32625 7 1 2 80629 86025
0 32626 7 2 2 62594 81822
0 32627 7 1 2 92736 98943
0 32628 7 1 2 32625 32627
0 32629 5 1 1 32628
0 32630 7 1 2 32624 32629
0 32631 5 1 1 32630
0 32632 7 1 2 98935 32631
0 32633 5 1 1 32632
0 32634 7 1 2 83315 84092
0 32635 5 1 1 32634
0 32636 7 1 2 88876 83986
0 32637 5 1 1 32636
0 32638 7 1 2 32635 32637
0 32639 5 1 1 32638
0 32640 7 1 2 65451 98795
0 32641 5 1 1 32640
0 32642 7 1 2 98816 32641
0 32643 5 1 1 32642
0 32644 7 1 2 68674 32643
0 32645 5 1 1 32644
0 32646 7 2 2 71535 86378
0 32647 7 2 2 98945 98881
0 32648 7 1 2 67282 98947
0 32649 5 1 1 32648
0 32650 7 1 2 32645 32649
0 32651 5 1 1 32650
0 32652 7 1 2 32639 32651
0 32653 5 1 1 32652
0 32654 7 1 2 73991 95016
0 32655 5 1 1 32654
0 32656 7 1 2 71972 88772
0 32657 7 1 2 86229 32656
0 32658 5 1 1 32657
0 32659 7 1 2 32655 32658
0 32660 5 1 1 32659
0 32661 7 1 2 61616 32660
0 32662 5 1 1 32661
0 32663 7 1 2 88301 76779
0 32664 7 1 2 88877 32663
0 32665 5 1 1 32664
0 32666 7 1 2 32662 32665
0 32667 5 1 1 32666
0 32668 7 1 2 85077 32667
0 32669 5 1 1 32668
0 32670 7 1 2 79150 91436
0 32671 5 1 1 32670
0 32672 7 1 2 73992 79104
0 32673 5 1 1 32672
0 32674 7 1 2 32671 32673
0 32675 5 1 1 32674
0 32676 7 1 2 95663 32675
0 32677 5 1 1 32676
0 32678 7 1 2 32669 32677
0 32679 5 1 1 32678
0 32680 7 1 2 82279 32679
0 32681 5 1 1 32680
0 32682 7 1 2 86966 93357
0 32683 5 1 1 32682
0 32684 7 1 2 86005 93401
0 32685 5 1 1 32684
0 32686 7 1 2 32683 32685
0 32687 5 1 1 32686
0 32688 7 1 2 89014 84265
0 32689 7 1 2 32687 32688
0 32690 5 1 1 32689
0 32691 7 1 2 32681 32690
0 32692 5 1 1 32691
0 32693 7 1 2 98882 32692
0 32694 5 1 1 32693
0 32695 7 1 2 32653 32694
0 32696 5 1 1 32695
0 32697 7 1 2 92707 32696
0 32698 5 1 1 32697
0 32699 7 1 2 90254 74670
0 32700 5 3 1 32699
0 32701 7 1 2 62595 98949
0 32702 5 1 1 32701
0 32703 7 2 2 71590 74658
0 32704 5 1 1 98952
0 32705 7 1 2 32702 32704
0 32706 5 5 1 32705
0 32707 7 1 2 68675 98954
0 32708 5 1 1 32707
0 32709 7 1 2 77452 78291
0 32710 5 1 1 32709
0 32711 7 1 2 32708 32710
0 32712 5 1 1 32711
0 32713 7 1 2 87334 14902
0 32714 5 1 1 32713
0 32715 7 1 2 32712 32714
0 32716 5 1 1 32715
0 32717 7 1 2 89263 71614
0 32718 7 1 2 82355 32717
0 32719 5 1 1 32718
0 32720 7 1 2 32716 32719
0 32721 5 1 1 32720
0 32722 7 1 2 87307 32721
0 32723 5 1 1 32722
0 32724 7 1 2 72397 82492
0 32725 5 3 1 32724
0 32726 7 1 2 71850 98959
0 32727 5 1 1 32726
0 32728 7 4 2 68676 98950
0 32729 5 1 1 98962
0 32730 7 1 2 62596 98963
0 32731 5 1 1 32730
0 32732 7 1 2 32727 32731
0 32733 5 2 1 32732
0 32734 7 1 2 79642 87693
0 32735 7 1 2 98966 32734
0 32736 5 1 1 32735
0 32737 7 1 2 32723 32736
0 32738 5 1 1 32737
0 32739 7 1 2 62141 32738
0 32740 5 1 1 32739
0 32741 7 2 2 86967 77016
0 32742 5 1 1 98968
0 32743 7 2 2 69384 96118
0 32744 7 1 2 86358 86861
0 32745 7 1 2 98970 32744
0 32746 7 1 2 98969 32745
0 32747 5 1 1 32746
0 32748 7 1 2 32740 32747
0 32749 5 1 1 32748
0 32750 7 1 2 68026 32749
0 32751 5 1 1 32750
0 32752 7 1 2 83130 98967
0 32753 5 1 1 32752
0 32754 7 1 2 66758 91585
0 32755 7 1 2 92865 32754
0 32756 5 1 1 32755
0 32757 7 1 2 32753 32756
0 32758 5 1 1 32757
0 32759 7 1 2 62142 32758
0 32760 5 1 1 32759
0 32761 7 5 2 62427 88559
0 32762 7 1 2 66759 74280
0 32763 7 1 2 78397 32762
0 32764 7 1 2 98972 32763
0 32765 5 1 1 32764
0 32766 7 1 2 32760 32765
0 32767 5 1 1 32766
0 32768 7 1 2 81930 32767
0 32769 5 1 1 32768
0 32770 7 1 2 89925 80235
0 32771 7 1 2 91793 32770
0 32772 7 1 2 97220 32771
0 32773 5 1 1 32772
0 32774 7 1 2 32769 32773
0 32775 5 1 1 32774
0 32776 7 1 2 89019 32775
0 32777 5 1 1 32776
0 32778 7 1 2 32751 32777
0 32779 5 1 1 32778
0 32780 7 1 2 97737 32779
0 32781 5 1 1 32780
0 32782 7 1 2 32698 32781
0 32783 7 1 2 32633 32782
0 32784 7 1 2 32577 32783
0 32785 5 1 1 32784
0 32786 7 1 2 90709 32785
0 32787 5 1 1 32786
0 32788 7 8 2 64368 97981
0 32789 7 4 2 75160 79868
0 32790 5 1 1 98985
0 32791 7 1 2 75777 79919
0 32792 5 1 1 32791
0 32793 7 1 2 32790 32792
0 32794 5 1 1 32793
0 32795 7 1 2 63821 32794
0 32796 5 1 1 32795
0 32797 7 1 2 75778 98517
0 32798 5 1 1 32797
0 32799 7 1 2 32796 32798
0 32800 5 2 1 32799
0 32801 7 2 2 63364 93774
0 32802 7 1 2 83299 98991
0 32803 7 1 2 98989 32802
0 32804 5 1 1 32803
0 32805 7 1 2 63365 98069
0 32806 7 1 2 93070 32805
0 32807 5 1 1 32806
0 32808 7 1 2 66229 77204
0 32809 7 1 2 93684 98573
0 32810 7 1 2 32808 32809
0 32811 5 1 1 32810
0 32812 7 1 2 32807 32811
0 32813 5 1 1 32812
0 32814 7 1 2 68427 32813
0 32815 7 1 2 98824 32814
0 32816 5 1 1 32815
0 32817 7 1 2 32804 32816
0 32818 5 1 1 32817
0 32819 7 1 2 65789 32818
0 32820 5 1 1 32819
0 32821 7 1 2 75421 73467
0 32822 7 1 2 87681 32821
0 32823 7 1 2 93775 32822
0 32824 7 1 2 88229 32823
0 32825 5 1 1 32824
0 32826 7 1 2 32820 32825
0 32827 5 1 1 32826
0 32828 7 1 2 98977 32827
0 32829 5 1 1 32828
0 32830 7 1 2 97029 98380
0 32831 5 1 1 32830
0 32832 7 6 2 63010 68428
0 32833 7 2 2 83131 98993
0 32834 7 2 2 66513 75963
0 32835 7 1 2 98999 99001
0 32836 5 1 1 32835
0 32837 7 1 2 32831 32836
0 32838 5 1 1 32837
0 32839 7 1 2 71591 32838
0 32840 5 1 1 32839
0 32841 7 1 2 92250 94336
0 32842 7 1 2 99000 32841
0 32843 5 1 1 32842
0 32844 7 1 2 32840 32843
0 32845 5 1 1 32844
0 32846 7 1 2 66997 32845
0 32847 5 1 1 32846
0 32848 7 2 2 71592 94212
0 32849 7 4 2 67859 63366
0 32850 7 1 2 82913 99005
0 32851 7 1 2 99003 32850
0 32852 5 1 1 32851
0 32853 7 1 2 32847 32852
0 32854 5 1 1 32853
0 32855 7 1 2 61364 32854
0 32856 5 1 1 32855
0 32857 7 3 2 71593 94812
0 32858 5 2 1 99009
0 32859 7 17 2 66230 61617
0 32860 5 1 1 99014
0 32861 7 3 2 63011 99015
0 32862 7 1 2 82378 99031
0 32863 7 1 2 99010 32862
0 32864 5 1 1 32863
0 32865 7 1 2 32856 32864
0 32866 5 1 1 32865
0 32867 7 1 2 93847 32866
0 32868 5 1 1 32867
0 32869 7 8 2 61286 61899
0 32870 7 1 2 91380 99034
0 32871 7 1 2 98992 32870
0 32872 7 1 2 99011 32871
0 32873 5 1 1 32872
0 32874 7 1 2 32868 32873
0 32875 5 1 1 32874
0 32876 7 1 2 69218 32875
0 32877 5 1 1 32876
0 32878 7 17 2 93776 93852
0 32879 7 2 2 82379 90006
0 32880 7 1 2 74680 96434
0 32881 7 1 2 99059 32880
0 32882 7 1 2 99042 32881
0 32883 5 1 1 32882
0 32884 7 1 2 87429 90795
0 32885 7 1 2 92189 96110
0 32886 7 3 2 63012 70386
0 32887 7 1 2 96939 99061
0 32888 7 1 2 32885 32887
0 32889 7 1 2 32884 32888
0 32890 5 1 1 32889
0 32891 7 1 2 32883 32890
0 32892 5 1 1 32891
0 32893 7 1 2 96282 32892
0 32894 5 1 1 32893
0 32895 7 1 2 82914 95929
0 32896 7 1 2 99043 32895
0 32897 7 1 2 98964 32896
0 32898 5 1 1 32897
0 32899 7 1 2 32894 32898
0 32900 5 1 1 32899
0 32901 7 1 2 62597 32900
0 32902 5 1 1 32901
0 32903 7 1 2 66514 91329
0 32904 7 1 2 88413 32903
0 32905 7 1 2 91356 32904
0 32906 7 1 2 82693 32905
0 32907 5 1 1 32906
0 32908 7 1 2 32902 32907
0 32909 7 1 2 32877 32908
0 32910 5 1 1 32909
0 32911 7 1 2 64268 32910
0 32912 5 1 1 32911
0 32913 7 1 2 32829 32912
0 32914 5 1 1 32913
0 32915 7 1 2 64759 32914
0 32916 5 1 1 32915
0 32917 7 3 2 61900 62966
0 32918 7 3 2 64269 99064
0 32919 7 5 2 70387 74361
0 32920 7 1 2 92943 99070
0 32921 7 1 2 99067 32920
0 32922 5 1 1 32921
0 32923 7 1 2 84196 91550
0 32924 7 1 2 97305 32923
0 32925 5 1 1 32924
0 32926 7 1 2 32922 32925
0 32927 5 1 1 32926
0 32928 7 1 2 63367 32927
0 32929 5 1 1 32928
0 32930 7 3 2 67790 68201
0 32931 7 2 2 87682 99075
0 32932 7 1 2 76236 98035
0 32933 7 1 2 99078 32932
0 32934 5 1 1 32933
0 32935 7 1 2 32929 32934
0 32936 5 1 1 32935
0 32937 7 1 2 68677 32936
0 32938 5 1 1 32937
0 32939 7 2 2 69116 75161
0 32940 7 1 2 77745 99079
0 32941 7 1 2 99080 32940
0 32942 5 1 1 32941
0 32943 7 1 2 32938 32942
0 32944 5 1 1 32943
0 32945 7 1 2 93660 32944
0 32946 5 1 1 32945
0 32947 7 1 2 94766 96435
0 32948 7 2 2 93853 32947
0 32949 7 2 2 71783 81843
0 32950 7 1 2 74457 99084
0 32951 7 1 2 99082 32950
0 32952 5 1 1 32951
0 32953 7 1 2 32946 32952
0 32954 5 1 1 32953
0 32955 7 1 2 62598 32954
0 32956 5 1 1 32955
0 32957 7 1 2 90162 90589
0 32958 7 7 2 62428 67791
0 32959 7 2 2 66113 99086
0 32960 7 1 2 98582 99093
0 32961 7 1 2 32957 32960
0 32962 5 1 1 32961
0 32963 7 1 2 32956 32962
0 32964 5 1 1 32963
0 32965 7 8 2 62861 93777
0 32966 7 1 2 91189 99095
0 32967 7 1 2 32964 32966
0 32968 5 1 1 32967
0 32969 7 1 2 32916 32968
0 32970 5 1 1 32969
0 32971 7 1 2 69385 32970
0 32972 5 1 1 32971
0 32973 7 9 2 61618 67860
0 32974 5 1 1 99103
0 32975 7 1 2 67792 99104
0 32976 7 1 2 98716 32975
0 32977 7 1 2 97206 32976
0 32978 5 1 1 32977
0 32979 7 5 2 63013 92190
0 32980 7 10 2 64270 70388
0 32981 7 1 2 81682 99117
0 32982 7 1 2 98629 32981
0 32983 7 1 2 99112 32982
0 32984 5 1 1 32983
0 32985 7 1 2 32978 32984
0 32986 5 1 1 32985
0 32987 7 1 2 63822 32986
0 32988 5 1 1 32987
0 32989 7 1 2 88518 25556
0 32990 5 3 1 32989
0 32991 7 1 2 97664 99127
0 32992 5 1 1 32991
0 32993 7 1 2 91862 97786
0 32994 7 5 2 97572 32993
0 32995 5 1 1 99130
0 32996 7 1 2 76447 99131
0 32997 5 1 1 32996
0 32998 7 2 2 32992 32997
0 32999 5 1 1 99135
0 33000 7 3 2 65452 75805
0 33001 5 1 1 99137
0 33002 7 1 2 71973 99138
0 33003 7 1 2 97665 33002
0 33004 5 1 1 33003
0 33005 7 1 2 99136 33004
0 33006 5 2 1 33005
0 33007 7 1 2 96877 99140
0 33008 5 1 1 33007
0 33009 7 1 2 32988 33008
0 33010 5 1 1 33009
0 33011 7 1 2 85572 33010
0 33012 5 1 1 33011
0 33013 7 1 2 91548 97221
0 33014 5 1 1 33013
0 33015 7 2 2 85696 96408
0 33016 7 1 2 96878 99142
0 33017 5 1 1 33016
0 33018 7 1 2 33014 33017
0 33019 5 1 1 33018
0 33020 7 1 2 97666 33019
0 33021 5 1 1 33020
0 33022 7 1 2 33012 33021
0 33023 5 1 1 33022
0 33024 7 1 2 87717 33023
0 33025 5 1 1 33024
0 33026 7 3 2 64271 90603
0 33027 7 10 2 98374 99144
0 33028 5 1 1 99147
0 33029 7 1 2 90238 89855
0 33030 7 1 2 99148 33029
0 33031 7 1 2 96456 33030
0 33032 5 1 1 33031
0 33033 7 1 2 33025 33032
0 33034 5 1 1 33033
0 33035 7 1 2 93666 33034
0 33036 5 1 1 33035
0 33037 7 1 2 32972 33036
0 33038 5 1 1 33037
0 33039 7 1 2 63181 33038
0 33040 5 1 1 33039
0 33041 7 1 2 64272 87361
0 33042 7 3 2 62599 98436
0 33043 7 3 2 63977 90604
0 33044 7 1 2 99157 99160
0 33045 7 1 2 33041 33044
0 33046 5 1 1 33045
0 33047 7 10 2 63582 69117
0 33048 7 2 2 99016 99163
0 33049 7 1 2 64760 91863
0 33050 7 1 2 79910 33049
0 33051 7 1 2 99173 33050
0 33052 5 1 1 33051
0 33053 7 1 2 33046 33052
0 33054 5 1 1 33053
0 33055 7 1 2 70389 33054
0 33056 5 1 1 33055
0 33057 7 1 2 62862 93402
0 33058 5 1 1 33057
0 33059 7 1 2 97075 33058
0 33060 5 1 1 33059
0 33061 7 1 2 74659 98008
0 33062 7 1 2 33060 33061
0 33063 5 1 1 33062
0 33064 7 1 2 33056 33063
0 33065 5 1 1 33064
0 33066 7 1 2 62143 33065
0 33067 5 1 1 33066
0 33068 7 3 2 70390 87362
0 33069 7 2 2 95164 98437
0 33070 7 1 2 73715 90605
0 33071 7 1 2 99178 33070
0 33072 7 1 2 99175 33071
0 33073 5 1 1 33072
0 33074 7 1 2 33067 33073
0 33075 5 1 1 33074
0 33076 7 1 2 68678 33075
0 33077 5 1 1 33076
0 33078 7 3 2 63583 85969
0 33079 5 1 1 99180
0 33080 7 1 2 98009 99181
0 33081 5 1 1 33080
0 33082 7 2 2 62863 97667
0 33083 7 1 2 76470 99183
0 33084 5 1 1 33083
0 33085 7 1 2 33081 33084
0 33086 5 1 1 33085
0 33087 7 1 2 65453 33086
0 33088 5 1 1 33087
0 33089 7 1 2 82196 72892
0 33090 5 1 1 33089
0 33091 7 1 2 77720 76403
0 33092 5 3 1 33091
0 33093 7 1 2 33090 99185
0 33094 5 1 1 33093
0 33095 7 1 2 98010 33094
0 33096 5 1 1 33095
0 33097 7 1 2 33088 33096
0 33098 5 1 1 33097
0 33099 7 1 2 62144 33098
0 33100 5 1 1 33099
0 33101 7 4 2 66231 90877
0 33102 7 5 2 67861 69118
0 33103 7 1 2 86615 99192
0 33104 7 2 2 99188 33103
0 33105 7 2 2 84718 99197
0 33106 5 1 1 99199
0 33107 7 1 2 33100 33106
0 33108 5 1 1 33107
0 33109 7 1 2 86968 33108
0 33110 5 1 1 33109
0 33111 7 1 2 33077 33110
0 33112 5 1 1 33111
0 33113 7 1 2 87718 33112
0 33114 5 1 1 33113
0 33115 7 8 2 61365 61619
0 33116 7 4 2 66114 99201
0 33117 7 2 2 63014 93904
0 33118 7 2 2 99209 99213
0 33119 7 1 2 77152 97366
0 33120 7 2 2 80890 33119
0 33121 7 1 2 64761 99217
0 33122 7 1 2 99215 33121
0 33123 5 1 1 33122
0 33124 7 1 2 33114 33123
0 33125 5 1 1 33124
0 33126 7 1 2 65790 33125
0 33127 5 1 1 33126
0 33128 7 1 2 82485 98951
0 33129 5 1 1 33128
0 33130 7 1 2 99012 33129
0 33131 5 1 1 33130
0 33132 7 4 2 63015 64273
0 33133 7 5 2 61620 62967
0 33134 7 3 2 99219 99223
0 33135 7 1 2 90986 92116
0 33136 7 1 2 99228 33135
0 33137 7 1 2 33131 33136
0 33138 5 1 1 33137
0 33139 7 1 2 33127 33138
0 33140 5 1 1 33139
0 33141 7 1 2 66760 33140
0 33142 5 1 1 33141
0 33143 7 2 2 87719 98078
0 33144 7 1 2 63978 99231
0 33145 5 1 1 33144
0 33146 7 2 2 93905 98121
0 33147 7 1 2 90987 91743
0 33148 7 1 2 99233 33147
0 33149 5 1 1 33148
0 33150 7 1 2 33145 33149
0 33151 5 1 1 33150
0 33152 7 1 2 72386 33151
0 33153 5 1 1 33152
0 33154 7 1 2 72401 99149
0 33155 5 1 1 33154
0 33156 7 1 2 33153 33155
0 33157 5 1 1 33156
0 33158 7 1 2 65454 33157
0 33159 5 1 1 33158
0 33160 7 2 2 90988 98126
0 33161 7 1 2 98910 99235
0 33162 5 1 1 33161
0 33163 7 1 2 75667 92459
0 33164 7 1 2 98583 33163
0 33165 7 1 2 92422 33164
0 33166 5 1 1 33165
0 33167 7 1 2 33162 33166
0 33168 5 1 1 33167
0 33169 7 1 2 66998 33168
0 33170 5 1 1 33169
0 33171 7 1 2 33159 33170
0 33172 5 1 1 33171
0 33173 7 1 2 68679 33172
0 33174 5 1 1 33173
0 33175 7 1 2 92460 98908
0 33176 5 1 1 33175
0 33177 7 1 2 91008 98914
0 33178 5 1 1 33177
0 33179 7 1 2 33176 33178
0 33180 5 1 1 33179
0 33181 7 1 2 71251 33180
0 33182 5 1 1 33181
0 33183 7 3 2 91864 98600
0 33184 7 1 2 61287 99237
0 33185 7 1 2 98921 33184
0 33186 5 1 1 33185
0 33187 7 1 2 33182 33186
0 33188 5 1 1 33187
0 33189 7 1 2 66999 33188
0 33190 5 1 1 33189
0 33191 7 1 2 33174 33190
0 33192 5 1 1 33191
0 33193 7 1 2 86969 79777
0 33194 7 1 2 33192 33193
0 33195 5 1 1 33194
0 33196 7 1 2 33142 33195
0 33197 5 1 1 33196
0 33198 7 1 2 68202 33197
0 33199 5 1 1 33198
0 33200 7 2 2 82631 83417
0 33201 7 2 2 68680 74493
0 33202 5 1 1 99242
0 33203 7 1 2 6328 21726
0 33204 5 3 1 33203
0 33205 7 2 2 70732 99244
0 33206 5 1 1 99247
0 33207 7 1 2 33202 33206
0 33208 5 4 1 33207
0 33209 7 1 2 99150 99249
0 33210 5 1 1 33209
0 33211 7 6 2 69119 90662
0 33212 7 3 2 64369 92957
0 33213 7 3 2 99253 99259
0 33214 7 1 2 99262 98826
0 33215 5 1 1 33214
0 33216 7 1 2 33210 33215
0 33217 5 1 1 33216
0 33218 7 1 2 86970 33217
0 33219 5 1 1 33218
0 33220 7 1 2 86928 99087
0 33221 7 1 2 92981 33220
0 33222 7 2 2 65791 94366
0 33223 7 1 2 99265 99002
0 33224 7 1 2 33221 33223
0 33225 5 1 1 33224
0 33226 7 1 2 33219 33225
0 33227 5 1 1 33226
0 33228 7 1 2 99240 33227
0 33229 5 1 1 33228
0 33230 7 1 2 33199 33229
0 33231 5 1 1 33230
0 33232 7 1 2 84077 33231
0 33233 5 1 1 33232
0 33234 7 1 2 33040 33233
0 33235 5 1 1 33234
0 33236 7 1 2 64963 33235
0 33237 5 1 1 33236
0 33238 7 1 2 85442 92298
0 33239 7 1 2 98193 33238
0 33240 5 1 1 33239
0 33241 7 1 2 87968 77363
0 33242 5 2 1 33241
0 33243 7 1 2 69120 79316
0 33244 7 1 2 93691 33243
0 33245 7 1 2 99267 33244
0 33246 5 1 1 33245
0 33247 7 1 2 33240 33246
0 33248 5 1 1 33247
0 33249 7 1 2 89980 33248
0 33250 5 1 1 33249
0 33251 7 2 2 97644 98545
0 33252 7 2 2 75779 79513
0 33253 5 1 1 99271
0 33254 7 1 2 74734 99272
0 33255 7 1 2 99269 33254
0 33256 5 1 1 33255
0 33257 7 1 2 33250 33256
0 33258 5 1 1 33257
0 33259 7 1 2 66232 33258
0 33260 5 1 1 33259
0 33261 7 1 2 89651 98122
0 33262 7 1 2 93487 33261
0 33263 5 1 1 33262
0 33264 7 1 2 82669 98047
0 33265 7 1 2 98955 33264
0 33266 5 1 1 33265
0 33267 7 1 2 33263 33266
0 33268 5 1 1 33267
0 33269 7 6 2 61366 62864
0 33270 7 1 2 99273 97645
0 33271 7 1 2 33268 33270
0 33272 5 1 1 33271
0 33273 7 1 2 33260 33272
0 33274 5 1 1 33273
0 33275 7 1 2 66761 33274
0 33276 5 1 1 33275
0 33277 7 2 2 93778 98956
0 33278 7 1 2 88672 78701
0 33279 7 1 2 99068 33278
0 33280 7 1 2 99279 33279
0 33281 5 1 1 33280
0 33282 7 1 2 33276 33281
0 33283 5 1 1 33282
0 33284 7 1 2 66115 33283
0 33285 5 1 1 33284
0 33286 7 3 2 61288 62145
0 33287 7 1 2 83132 99281
0 33288 7 1 2 98774 33287
0 33289 7 1 2 99280 33288
0 33290 5 1 1 33289
0 33291 7 1 2 33285 33290
0 33292 5 1 1 33291
0 33293 7 1 2 69219 33292
0 33294 5 1 1 33293
0 33295 7 2 2 66116 73335
0 33296 7 4 2 62146 74660
0 33297 7 1 2 98546 99286
0 33298 7 1 2 99284 33297
0 33299 5 1 1 33298
0 33300 7 1 2 61289 67862
0 33301 7 1 2 88724 33300
0 33302 7 1 2 86447 33301
0 33303 5 1 1 33302
0 33304 7 1 2 33299 33303
0 33305 5 1 1 33304
0 33306 7 1 2 66762 33305
0 33307 5 1 1 33306
0 33308 7 2 2 61901 98103
0 33309 7 1 2 99290 99285
0 33310 7 1 2 97207 33309
0 33311 5 1 1 33310
0 33312 7 1 2 33307 33311
0 33313 5 1 1 33312
0 33314 7 1 2 66233 33313
0 33315 5 1 1 33314
0 33316 7 1 2 65455 90989
0 33317 7 1 2 91361 92089
0 33318 7 1 2 33316 33317
0 33319 7 1 2 95037 33318
0 33320 5 1 1 33319
0 33321 7 1 2 33315 33320
0 33322 5 1 1 33321
0 33323 7 1 2 97982 33322
0 33324 5 1 1 33323
0 33325 7 3 2 62968 93779
0 33326 7 1 2 62600 90066
0 33327 7 4 2 61290 95165
0 33328 7 1 2 99071 99295
0 33329 7 1 2 33326 33328
0 33330 7 1 2 99292 33329
0 33331 5 1 1 33330
0 33332 7 1 2 33324 33331
0 33333 5 1 1 33332
0 33334 7 1 2 65792 96111
0 33335 7 1 2 33333 33334
0 33336 5 1 1 33335
0 33337 7 1 2 33294 33336
0 33338 5 1 1 33337
0 33339 7 1 2 68681 33338
0 33340 5 1 1 33339
0 33341 7 5 2 64370 94757
0 33342 7 5 2 67793 63979
0 33343 7 1 2 99299 99304
0 33344 5 1 1 33343
0 33345 7 3 2 62969 65456
0 33346 7 3 2 68863 93906
0 33347 7 1 2 99309 99312
0 33348 5 1 1 33347
0 33349 7 1 2 33344 33348
0 33350 5 1 1 33349
0 33351 7 1 2 62147 33350
0 33352 5 1 1 33351
0 33353 7 5 2 67794 63584
0 33354 7 2 2 94367 95221
0 33355 7 1 2 99315 99320
0 33356 5 1 1 33355
0 33357 7 1 2 33352 33356
0 33358 5 1 1 33357
0 33359 7 1 2 66117 33358
0 33360 5 1 1 33359
0 33361 7 1 2 86059 97357
0 33362 7 1 2 97613 33361
0 33363 5 1 1 33362
0 33364 7 1 2 33360 33363
0 33365 5 1 1 33364
0 33366 7 1 2 83133 33365
0 33367 5 1 1 33366
0 33368 7 1 2 83666 99083
0 33369 5 1 1 33368
0 33370 7 1 2 33367 33369
0 33371 5 1 1 33370
0 33372 7 1 2 62601 33371
0 33373 5 1 1 33372
0 33374 7 2 2 96940 98154
0 33375 5 1 1 99322
0 33376 7 1 2 90159 99323
0 33377 5 1 1 33376
0 33378 7 7 2 66118 97983
0 33379 7 4 2 72852 99324
0 33380 5 1 1 99331
0 33381 7 1 2 83667 99332
0 33382 5 1 1 33381
0 33383 7 1 2 33377 33382
0 33384 5 1 1 33383
0 33385 7 1 2 64371 33384
0 33386 5 1 1 33385
0 33387 7 1 2 33373 33386
0 33388 5 1 1 33387
0 33389 7 1 2 71851 33388
0 33390 5 1 1 33389
0 33391 7 1 2 89413 93593
0 33392 7 1 2 98543 33391
0 33393 5 1 1 33392
0 33394 7 1 2 33390 33393
0 33395 5 1 1 33394
0 33396 7 3 2 65793 93780
0 33397 7 1 2 78702 99335
0 33398 7 1 2 33395 33397
0 33399 5 1 1 33398
0 33400 7 1 2 33340 33399
0 33401 5 1 1 33400
0 33402 7 1 2 61621 33401
0 33403 5 1 1 33402
0 33404 7 2 2 92982 98612
0 33405 7 1 2 94213 99338
0 33406 5 1 1 33405
0 33407 7 5 2 69220 71734
0 33408 7 1 2 74813 90990
0 33409 7 1 2 99340 33408
0 33410 7 1 2 98194 33409
0 33411 5 1 1 33410
0 33412 7 1 2 33406 33411
0 33413 5 1 1 33412
0 33414 7 1 2 63980 33413
0 33415 5 1 1 33414
0 33416 7 2 2 65457 96128
0 33417 7 1 2 99151 99345
0 33418 5 1 1 33417
0 33419 7 1 2 33415 33418
0 33420 5 1 1 33419
0 33421 7 1 2 62602 33420
0 33422 5 1 1 33421
0 33423 7 1 2 91009 94668
0 33424 7 1 2 98953 33423
0 33425 5 1 1 33424
0 33426 7 1 2 33422 33425
0 33427 5 1 1 33426
0 33428 7 1 2 62148 33427
0 33429 5 1 1 33428
0 33430 7 1 2 87768 99200
0 33431 5 1 1 33430
0 33432 7 1 2 33429 33431
0 33433 5 1 1 33432
0 33434 7 1 2 83134 33433
0 33435 5 1 1 33434
0 33436 7 1 2 65458 77646
0 33437 5 1 1 33436
0 33438 7 1 2 74362 85216
0 33439 5 2 1 33438
0 33440 7 1 2 70391 99347
0 33441 5 1 1 33440
0 33442 7 2 2 88166 99035
0 33443 7 3 2 63016 68203
0 33444 7 2 2 64274 99351
0 33445 7 1 2 97419 99354
0 33446 7 1 2 99349 33445
0 33447 7 1 2 33441 33446
0 33448 7 1 2 33437 33447
0 33449 5 1 1 33448
0 33450 7 1 2 33435 33449
0 33451 5 1 1 33450
0 33452 7 1 2 89548 33451
0 33453 5 1 1 33452
0 33454 7 1 2 33403 33453
0 33455 5 1 1 33454
0 33456 7 1 2 64762 33455
0 33457 5 1 1 33456
0 33458 7 2 2 67795 74888
0 33459 7 1 2 95276 99356
0 33460 5 1 1 33459
0 33461 7 2 2 62970 71852
0 33462 7 1 2 99313 99358
0 33463 5 1 1 33462
0 33464 7 1 2 33460 33463
0 33465 5 1 1 33464
0 33466 7 1 2 66119 33465
0 33467 5 1 1 33466
0 33468 7 1 2 74681 99088
0 33469 7 1 2 97614 33468
0 33470 5 1 1 33469
0 33471 7 1 2 33467 33470
0 33472 5 1 1 33471
0 33473 7 1 2 88673 33472
0 33474 5 1 1 33473
0 33475 7 3 2 68682 83418
0 33476 5 1 1 99360
0 33477 7 11 2 67000 67796
0 33478 7 6 2 66120 99363
0 33479 7 1 2 95277 99374
0 33480 7 1 2 99361 33479
0 33481 5 1 1 33480
0 33482 7 1 2 33474 33481
0 33483 5 1 1 33482
0 33484 7 11 2 76171 93781
0 33485 7 1 2 89291 92274
0 33486 7 1 2 99380 33485
0 33487 7 1 2 33483 33486
0 33488 5 1 1 33487
0 33489 7 1 2 69386 33488
0 33490 7 1 2 33457 33489
0 33491 5 1 1 33490
0 33492 7 1 2 71252 99141
0 33493 5 1 1 33492
0 33494 7 1 2 97668 99143
0 33495 5 1 1 33494
0 33496 7 1 2 33493 33495
0 33497 5 1 1 33496
0 33498 7 3 2 66515 91190
0 33499 5 2 1 99391
0 33500 7 1 2 95687 99394
0 33501 5 1 1 33500
0 33502 7 1 2 33497 33501
0 33503 5 1 1 33502
0 33504 7 1 2 74814 83459
0 33505 7 1 2 97573 33504
0 33506 7 1 2 96988 97564
0 33507 7 1 2 33505 33506
0 33508 5 1 1 33507
0 33509 7 3 2 66516 76712
0 33510 7 1 2 89041 99396
0 33511 7 1 2 97669 33510
0 33512 5 1 1 33511
0 33513 7 1 2 33508 33512
0 33514 7 1 2 33503 33513
0 33515 5 1 1 33514
0 33516 7 1 2 63368 33515
0 33517 5 1 1 33516
0 33518 7 1 2 68429 86576
0 33519 7 1 2 98079 33518
0 33520 5 1 1 33519
0 33521 7 1 2 81589 99118
0 33522 7 1 2 91342 33521
0 33523 5 1 1 33522
0 33524 7 1 2 33520 33523
0 33525 5 1 1 33524
0 33526 7 1 2 85814 95682
0 33527 7 1 2 33525 33526
0 33528 5 1 1 33527
0 33529 7 1 2 33517 33528
0 33530 5 1 1 33529
0 33531 7 1 2 87720 33530
0 33532 5 1 1 33531
0 33533 7 1 2 82646 75964
0 33534 5 1 1 33533
0 33535 7 1 2 68430 97079
0 33536 5 1 1 33535
0 33537 7 1 2 33534 33536
0 33538 5 1 1 33537
0 33539 7 1 2 67283 33538
0 33540 5 1 1 33539
0 33541 7 1 2 89315 84632
0 33542 5 1 1 33541
0 33543 7 1 2 33540 33542
0 33544 5 1 1 33543
0 33545 7 1 2 75897 33544
0 33546 5 1 1 33545
0 33547 7 2 2 88337 90771
0 33548 7 1 2 82488 99399
0 33549 5 1 1 33548
0 33550 7 1 2 33546 33549
0 33551 5 1 1 33550
0 33552 7 1 2 84798 99152
0 33553 7 1 2 33551 33552
0 33554 5 1 1 33553
0 33555 7 1 2 33532 33554
0 33556 5 1 1 33555
0 33557 7 1 2 63182 33556
0 33558 5 1 1 33557
0 33559 7 1 2 90239 96862
0 33560 5 1 1 33559
0 33561 7 2 2 76172 92708
0 33562 7 1 2 69589 99401
0 33563 5 1 1 33562
0 33564 7 1 2 33560 33563
0 33565 5 1 1 33564
0 33566 7 1 2 98189 33565
0 33567 5 1 1 33566
0 33568 7 2 2 61367 86971
0 33569 7 1 2 76484 99403
0 33570 7 1 2 99270 33569
0 33571 5 1 1 33570
0 33572 7 1 2 33567 33571
0 33573 5 1 1 33572
0 33574 7 1 2 65459 33573
0 33575 5 1 1 33574
0 33576 7 1 2 63369 32999
0 33577 5 1 1 33576
0 33578 7 1 2 68204 90924
0 33579 7 1 2 97670 33578
0 33580 5 1 1 33579
0 33581 7 1 2 33577 33580
0 33582 5 1 1 33581
0 33583 7 1 2 94650 33582
0 33584 5 1 1 33583
0 33585 7 1 2 33575 33584
0 33586 5 1 1 33585
0 33587 7 1 2 78429 33586
0 33588 5 1 1 33587
0 33589 7 3 2 64275 92191
0 33590 7 5 2 63017 69590
0 33591 7 1 2 75578 99408
0 33592 7 1 2 98630 33591
0 33593 7 1 2 99405 33592
0 33594 7 1 2 85701 33593
0 33595 5 1 1 33594
0 33596 7 1 2 33588 33595
0 33597 5 1 1 33596
0 33598 7 1 2 87721 33597
0 33599 5 1 1 33598
0 33600 7 1 2 96890 97051
0 33601 7 1 2 94337 33600
0 33602 7 1 2 99153 33601
0 33603 5 1 1 33602
0 33604 7 1 2 33599 33603
0 33605 5 1 1 33604
0 33606 7 1 2 73468 33605
0 33607 5 1 1 33606
0 33608 7 1 2 61902 33607
0 33609 7 1 2 33558 33608
0 33610 5 1 1 33609
0 33611 7 3 2 81823 93782
0 33612 7 7 2 64372 93854
0 33613 5 1 1 99416
0 33614 7 1 2 71974 80792
0 33615 7 1 2 83893 33614
0 33616 5 1 1 33615
0 33617 7 1 2 22785 33616
0 33618 5 1 1 33617
0 33619 7 1 2 77974 33618
0 33620 5 1 1 33619
0 33621 7 1 2 95688 28198
0 33622 5 3 1 33621
0 33623 7 1 2 74846 85452
0 33624 5 1 1 33623
0 33625 7 1 2 71975 33624
0 33626 7 1 2 99423 33625
0 33627 5 1 1 33626
0 33628 7 1 2 33620 33627
0 33629 5 1 1 33628
0 33630 7 1 2 99417 33629
0 33631 5 1 1 33630
0 33632 7 3 2 66121 87835
0 33633 7 1 2 67797 97287
0 33634 7 1 2 99426 33633
0 33635 7 1 2 99424 33634
0 33636 5 1 1 33635
0 33637 7 1 2 33631 33636
0 33638 5 1 1 33637
0 33639 7 1 2 70392 33638
0 33640 5 1 1 33639
0 33641 7 2 2 63823 93855
0 33642 7 1 2 82647 95645
0 33643 7 1 2 85573 33642
0 33644 7 1 2 99429 33643
0 33645 5 1 1 33644
0 33646 7 1 2 33640 33645
0 33647 5 1 1 33646
0 33648 7 1 2 69121 33647
0 33649 5 1 1 33648
0 33650 7 2 2 97709 97527
0 33651 7 1 2 71594 99400
0 33652 5 1 1 33651
0 33653 7 2 2 88626 92571
0 33654 5 1 1 99433
0 33655 7 1 2 82648 73469
0 33656 5 1 1 33655
0 33657 7 1 2 33654 33656
0 33658 5 1 1 33657
0 33659 7 1 2 94338 33658
0 33660 5 1 1 33659
0 33661 7 1 2 33652 33660
0 33662 5 1 1 33661
0 33663 7 1 2 99431 33662
0 33664 5 1 1 33663
0 33665 7 1 2 33649 33664
0 33666 5 1 1 33665
0 33667 7 1 2 67001 33666
0 33668 5 1 1 33667
0 33669 7 1 2 79696 99392
0 33670 5 3 1 33669
0 33671 7 1 2 80326 97276
0 33672 5 1 1 33671
0 33673 7 1 2 99435 33672
0 33674 5 1 1 33673
0 33675 7 4 2 61291 67284
0 33676 7 1 2 65460 99438
0 33677 7 2 2 98695 33676
0 33678 7 1 2 69221 99442
0 33679 7 1 2 33674 33678
0 33680 5 1 1 33679
0 33681 7 1 2 33668 33680
0 33682 5 1 1 33681
0 33683 7 1 2 68431 33682
0 33684 5 1 1 33683
0 33685 7 1 2 69222 88078
0 33686 7 3 2 64763 90240
0 33687 7 1 2 99444 98849
0 33688 7 1 2 98696 33687
0 33689 7 1 2 33685 33688
0 33690 5 1 1 33689
0 33691 7 1 2 33684 33690
0 33692 5 1 1 33691
0 33693 7 1 2 99413 33692
0 33694 5 1 1 33693
0 33695 7 1 2 32000 32995
0 33696 5 3 1 33695
0 33697 7 2 2 87722 99447
0 33698 5 1 1 99450
0 33699 7 1 2 67480 99451
0 33700 5 1 1 33699
0 33701 7 4 2 63018 97367
0 33702 7 3 2 90991 99452
0 33703 7 1 2 78398 93907
0 33704 7 1 2 99456 33703
0 33705 5 1 1 33704
0 33706 7 1 2 33700 33705
0 33707 5 1 1 33706
0 33708 7 1 2 81931 33707
0 33709 5 1 1 33708
0 33710 7 2 2 90663 99341
0 33711 7 1 2 78657 99325
0 33712 7 1 2 99459 33711
0 33713 5 1 1 33712
0 33714 7 1 2 33698 33713
0 33715 5 1 1 33714
0 33716 7 1 2 99425 33715
0 33717 5 1 1 33716
0 33718 7 4 2 64764 73074
0 33719 7 1 2 67481 93170
0 33720 7 1 2 99461 33719
0 33721 7 1 2 99216 33720
0 33722 5 1 1 33721
0 33723 7 1 2 33717 33722
0 33724 7 1 2 33709 33723
0 33725 5 1 1 33724
0 33726 7 1 2 87664 33725
0 33727 5 1 1 33726
0 33728 7 1 2 66763 33727
0 33729 7 1 2 33694 33728
0 33730 5 1 1 33729
0 33731 7 1 2 33610 33730
0 33732 5 1 1 33731
0 33733 7 2 2 80373 32729
0 33734 5 1 1 99465
0 33735 7 1 2 75857 33734
0 33736 5 1 1 33735
0 33737 7 1 2 99013 33736
0 33738 5 1 1 33737
0 33739 7 1 2 87788 33738
0 33740 5 1 1 33739
0 33741 7 1 2 33079 99348
0 33742 5 1 1 33741
0 33743 7 1 2 72456 87723
0 33744 7 1 2 33742 33743
0 33745 5 1 1 33744
0 33746 7 1 2 33740 33745
0 33747 5 1 1 33746
0 33748 7 1 2 97671 33747
0 33749 5 1 1 33748
0 33750 7 1 2 75780 94556
0 33751 5 1 1 33750
0 33752 7 1 2 63824 98986
0 33753 5 1 1 33752
0 33754 7 1 2 33751 33753
0 33755 5 1 1 33754
0 33756 7 1 2 99339 33755
0 33757 5 1 1 33756
0 33758 7 1 2 33749 33757
0 33759 5 1 1 33758
0 33760 7 1 2 88193 33759
0 33761 5 1 1 33760
0 33762 7 2 2 80984 99044
0 33763 5 1 1 99467
0 33764 7 3 2 92851 99017
0 33765 7 1 2 92958 99469
0 33766 5 1 1 33765
0 33767 7 1 2 33763 33766
0 33768 5 1 1 33767
0 33769 7 2 2 93165 98206
0 33770 7 1 2 74468 99472
0 33771 7 1 2 94200 33770
0 33772 7 1 2 33768 33771
0 33773 5 1 1 33772
0 33774 7 1 2 33761 33773
0 33775 5 1 1 33774
0 33776 7 1 2 83135 33775
0 33777 5 1 1 33776
0 33778 7 1 2 64534 33777
0 33779 7 1 2 33732 33778
0 33780 5 1 1 33779
0 33781 7 1 2 69822 33780
0 33782 7 1 2 33491 33781
0 33783 5 1 1 33782
0 33784 7 1 2 33237 33783
0 33785 7 1 2 32787 33784
0 33786 5 1 1 33785
0 33787 7 1 2 70095 33786
0 33788 5 1 1 33787
0 33789 7 1 2 82607 87962
0 33790 7 1 2 4531 14960
0 33791 5 1 1 33790
0 33792 7 1 2 4043 30788
0 33793 5 1 1 33792
0 33794 7 1 2 33791 33793
0 33795 7 1 2 33789 33794
0 33796 5 1 1 33795
0 33797 7 2 2 90992 96629
0 33798 7 1 2 87308 79697
0 33799 7 1 2 99474 33798
0 33800 5 1 1 33799
0 33801 7 1 2 33796 33800
0 33802 5 1 1 33801
0 33803 7 1 2 72457 33802
0 33804 5 1 1 33803
0 33805 7 3 2 70733 97856
0 33806 7 1 2 73336 90993
0 33807 7 1 2 96076 33806
0 33808 7 1 2 99476 33807
0 33809 5 1 1 33808
0 33810 7 1 2 33804 33809
0 33811 5 1 1 33810
0 33812 7 1 2 74363 33811
0 33813 5 1 1 33812
0 33814 7 1 2 88974 75711
0 33815 5 1 1 33814
0 33816 7 1 2 83136 92068
0 33817 5 1 1 33816
0 33818 7 1 2 33815 33817
0 33819 5 1 1 33818
0 33820 7 1 2 87724 33819
0 33821 5 1 1 33820
0 33822 7 2 2 85919 83304
0 33823 7 1 2 69223 96784
0 33824 7 1 2 99479 33823
0 33825 5 1 1 33824
0 33826 7 1 2 33821 33825
0 33827 5 1 1 33826
0 33828 7 38 2 61368 64535
0 33829 5 3 1 99481
0 33830 7 3 2 70393 99482
0 33831 5 1 1 99522
0 33832 7 1 2 80487 99523
0 33833 7 1 2 33827 33832
0 33834 5 1 1 33833
0 33835 7 1 2 33813 33834
0 33836 5 1 1 33835
0 33837 7 1 2 70096 33836
0 33838 5 1 1 33837
0 33839 7 4 2 61369 65172
0 33840 7 1 2 85793 98279
0 33841 5 2 1 33840
0 33842 7 1 2 87725 99529
0 33843 5 1 1 33842
0 33844 7 7 2 66122 62603
0 33845 7 1 2 68432 99531
0 33846 7 1 2 87931 33845
0 33847 5 1 1 33846
0 33848 7 1 2 33843 33847
0 33849 5 1 1 33848
0 33850 7 1 2 84492 33849
0 33851 5 1 1 33850
0 33852 7 4 2 66123 72705
0 33853 7 1 2 87836 99538
0 33854 5 1 1 33853
0 33855 7 1 2 97543 33854
0 33856 5 1 1 33855
0 33857 7 1 2 75806 33856
0 33858 5 1 1 33857
0 33859 7 1 2 98574 97420
0 33860 5 1 1 33859
0 33861 7 1 2 33858 33860
0 33862 5 1 1 33861
0 33863 7 1 2 82380 86140
0 33864 7 1 2 33862 33863
0 33865 5 1 1 33864
0 33866 7 1 2 33851 33865
0 33867 5 1 1 33866
0 33868 7 1 2 70394 33867
0 33869 5 1 1 33868
0 33870 7 1 2 64765 90904
0 33871 7 1 2 95991 33870
0 33872 7 1 2 87877 33871
0 33873 7 1 2 99477 33872
0 33874 5 1 1 33873
0 33875 7 1 2 33869 33874
0 33876 5 1 1 33875
0 33877 7 1 2 99525 33876
0 33878 5 1 1 33877
0 33879 7 1 2 33838 33878
0 33880 5 1 1 33879
0 33881 7 1 2 98195 33880
0 33882 5 1 1 33881
0 33883 7 1 2 97539 99287
0 33884 5 1 1 33883
0 33885 7 6 2 69224 99532
0 33886 7 3 2 73625 99542
0 33887 7 2 2 75162 99548
0 33888 5 1 1 99551
0 33889 7 1 2 33884 33888
0 33890 5 2 1 33889
0 33891 7 1 2 90830 99553
0 33892 5 1 1 33891
0 33893 7 1 2 79051 92709
0 33894 5 1 1 33893
0 33895 7 1 2 78292 96150
0 33896 5 1 1 33895
0 33897 7 1 2 33894 33896
0 33898 5 1 1 33897
0 33899 7 1 2 99543 33898
0 33900 5 1 1 33899
0 33901 7 2 2 65461 95341
0 33902 7 1 2 63370 97540
0 33903 7 1 2 99555 33902
0 33904 5 1 1 33903
0 33905 7 1 2 33900 33904
0 33906 5 1 1 33905
0 33907 7 1 2 79643 33906
0 33908 5 1 1 33907
0 33909 7 1 2 33892 33908
0 33910 5 1 1 33909
0 33911 7 1 2 66764 33910
0 33912 5 1 1 33911
0 33913 7 1 2 86141 99554
0 33914 5 1 1 33913
0 33915 7 2 2 96539 98575
0 33916 7 1 2 84589 79644
0 33917 7 1 2 99557 33916
0 33918 5 1 1 33917
0 33919 7 1 2 33914 33918
0 33920 5 1 1 33919
0 33921 7 1 2 70097 83062
0 33922 7 1 2 33920 33921
0 33923 5 1 1 33922
0 33924 7 1 2 33912 33923
0 33925 5 1 1 33924
0 33926 7 1 2 98011 33925
0 33927 5 1 1 33926
0 33928 7 3 2 61292 81590
0 33929 7 1 2 75596 93171
0 33930 7 2 2 99559 33929
0 33931 7 4 2 64536 93908
0 33932 7 1 2 99564 98149
0 33933 7 1 2 99562 33932
0 33934 5 1 1 33933
0 33935 7 2 2 83707 94368
0 33936 7 1 2 82794 92825
0 33937 7 1 2 99568 33936
0 33938 7 1 2 97209 33937
0 33939 5 1 1 33938
0 33940 7 1 2 33934 33939
0 33941 5 1 1 33940
0 33942 7 1 2 70098 33941
0 33943 5 1 1 33942
0 33944 7 2 2 73122 93856
0 33945 7 1 2 88560 76997
0 33946 7 1 2 89251 33945
0 33947 7 1 2 94645 33946
0 33948 7 1 2 99570 33947
0 33949 5 1 1 33948
0 33950 7 1 2 33943 33949
0 33951 5 1 1 33950
0 33952 7 1 2 93783 33951
0 33953 5 1 1 33952
0 33954 7 1 2 33927 33953
0 33955 7 1 2 33882 33954
0 33956 5 1 1 33955
0 33957 7 1 2 63183 33956
0 33958 5 1 1 33957
0 33959 7 2 2 87872 99533
0 33960 7 1 2 67863 73830
0 33961 7 1 2 92719 33960
0 33962 7 1 2 99572 33961
0 33963 5 1 1 33962
0 33964 7 13 2 62865 67864
0 33965 7 1 2 82440 99574
0 33966 5 2 1 33965
0 33967 7 1 2 62866 99587
0 33968 5 1 1 33967
0 33969 7 17 2 63019 64537
0 33970 5 7 1 99589
0 33971 7 1 2 99606 99588
0 33972 5 2 1 33971
0 33973 7 1 2 74661 87726
0 33974 7 1 2 99613 33973
0 33975 7 1 2 33968 33974
0 33976 5 1 1 33975
0 33977 7 1 2 33963 33976
0 33978 5 1 1 33977
0 33979 7 1 2 62149 33978
0 33980 5 1 1 33979
0 33981 7 1 2 83395 99575
0 33982 7 1 2 93940 33981
0 33983 7 1 2 99573 33982
0 33984 5 1 1 33983
0 33985 7 1 2 33980 33984
0 33986 5 1 1 33985
0 33987 7 1 2 66234 33986
0 33988 5 1 1 33987
0 33989 7 6 2 61293 61370
0 33990 7 3 2 64373 99615
0 33991 7 7 2 67865 63585
0 33992 7 1 2 74469 93736
0 33993 7 1 2 99624 33992
0 33994 7 1 2 99621 33993
0 33995 5 1 1 33994
0 33996 7 1 2 33988 33995
0 33997 5 1 1 33996
0 33998 7 1 2 83137 33997
0 33999 5 1 1 33998
0 34000 7 2 2 91390 92833
0 34001 7 4 2 67866 68864
0 34002 7 1 2 89286 99633
0 34003 7 1 2 99631 34002
0 34004 7 1 2 97210 34003
0 34005 5 1 1 34004
0 34006 7 1 2 33999 34005
0 34007 5 1 1 34006
0 34008 7 1 2 70099 34007
0 34009 5 1 1 34008
0 34010 7 1 2 87789 96359
0 34011 5 1 1 34010
0 34012 7 1 2 97544 34011
0 34013 5 3 1 34012
0 34014 7 1 2 76384 99637
0 34015 5 1 1 34014
0 34016 7 1 2 74328 99549
0 34017 5 1 1 34016
0 34018 7 1 2 34015 34017
0 34019 5 1 1 34018
0 34020 7 1 2 63371 34019
0 34021 5 1 1 34020
0 34022 7 4 2 94089 97433
0 34023 7 1 2 85012 81708
0 34024 7 1 2 99640 34023
0 34025 5 1 1 34024
0 34026 7 1 2 34021 34025
0 34027 5 1 1 34026
0 34028 7 31 2 67867 69387
0 34029 7 2 2 65173 99644
0 34030 7 1 2 98085 99675
0 34031 7 1 2 34027 34030
0 34032 5 1 1 34031
0 34033 7 1 2 34009 34032
0 34034 5 1 1 34033
0 34035 7 1 2 64766 34034
0 34036 5 1 1 34035
0 34037 7 3 2 79366 93685
0 34038 7 1 2 95196 99677
0 34039 7 1 2 99622 34038
0 34040 7 1 2 85429 34039
0 34041 5 1 1 34040
0 34042 7 1 2 34036 34041
0 34043 5 1 1 34042
0 34044 7 1 2 67798 34043
0 34045 5 1 1 34044
0 34046 7 2 2 83177 97193
0 34047 7 2 2 81709 93784
0 34048 7 1 2 93177 99682
0 34049 7 1 2 99680 34048
0 34050 5 1 1 34049
0 34051 7 1 2 34045 34050
0 34052 5 1 1 34051
0 34053 7 1 2 69122 34052
0 34054 5 1 1 34053
0 34055 7 2 2 72919 90994
0 34056 7 1 2 82441 98123
0 34057 7 1 2 99684 34056
0 34058 5 1 1 34057
0 34059 7 2 2 70734 91785
0 34060 7 8 2 61294 67708
0 34061 7 1 2 93785 99688
0 34062 7 1 2 99686 34061
0 34063 5 1 1 34062
0 34064 7 1 2 34058 34063
0 34065 5 1 1 34064
0 34066 7 1 2 70395 34065
0 34067 5 1 1 34066
0 34068 7 8 2 63020 69388
0 34069 7 1 2 73099 99696
0 34070 7 1 2 99685 34069
0 34071 5 1 1 34070
0 34072 7 1 2 34067 34071
0 34073 5 1 1 34072
0 34074 7 1 2 63586 34073
0 34075 5 1 1 34074
0 34076 7 5 2 62604 73123
0 34077 5 2 1 99704
0 34078 7 2 2 62867 97518
0 34079 7 1 2 87673 99711
0 34080 7 1 2 99705 34079
0 34081 5 1 1 34080
0 34082 7 1 2 34075 34081
0 34083 5 1 1 34082
0 34084 7 1 2 83063 34083
0 34085 5 1 1 34084
0 34086 7 3 2 74364 73124
0 34087 7 1 2 88920 70996
0 34088 7 1 2 99712 34087
0 34089 7 1 2 99713 34088
0 34090 5 1 1 34089
0 34091 7 1 2 34085 34090
0 34092 5 1 1 34091
0 34093 7 1 2 69225 34092
0 34094 5 1 1 34093
0 34095 7 1 2 83064 90606
0 34096 7 1 2 87727 34095
0 34097 7 2 2 65794 98644
0 34098 7 1 2 99072 99716
0 34099 7 1 2 34096 34098
0 34100 5 1 1 34099
0 34101 7 1 2 34094 34100
0 34102 5 1 1 34101
0 34103 7 1 2 83592 97646
0 34104 7 1 2 34102 34103
0 34105 5 1 1 34104
0 34106 7 1 2 34054 34105
0 34107 5 1 1 34106
0 34108 7 1 2 75354 34107
0 34109 5 1 1 34108
0 34110 7 1 2 33958 34109
0 34111 5 1 1 34110
0 34112 7 1 2 66517 34111
0 34113 5 1 1 34112
0 34114 7 12 2 61371 69389
0 34115 7 4 2 67799 99718
0 34116 7 2 2 99730 99706
0 34117 5 1 1 99734
0 34118 7 2 2 66235 71735
0 34119 7 10 2 62971 64538
0 34120 7 1 2 71020 99738
0 34121 7 1 2 99736 34120
0 34122 5 1 1 34121
0 34123 7 1 2 34117 34122
0 34124 5 1 1 34123
0 34125 7 1 2 86972 34124
0 34126 5 1 1 34125
0 34127 7 9 2 66236 64539
0 34128 7 2 2 91798 99748
0 34129 7 4 2 69591 71736
0 34130 7 1 2 80939 99759
0 34131 7 1 2 99757 34130
0 34132 5 1 1 34131
0 34133 7 1 2 34126 34132
0 34134 5 1 1 34133
0 34135 7 1 2 63587 34134
0 34136 5 1 1 34135
0 34137 7 1 2 96999 99735
0 34138 5 1 1 34137
0 34139 7 1 2 34136 34138
0 34140 5 1 1 34139
0 34141 7 1 2 61295 34140
0 34142 5 1 1 34141
0 34143 7 3 2 62972 69390
0 34144 7 1 2 90995 99763
0 34145 7 1 2 94834 34144
0 34146 7 1 2 99714 34145
0 34147 5 1 1 34146
0 34148 7 1 2 34142 34147
0 34149 5 1 1 34148
0 34150 7 1 2 69226 34149
0 34151 5 1 1 34150
0 34152 7 5 2 64374 96941
0 34153 7 3 2 72458 99766
0 34154 5 1 1 99771
0 34155 7 1 2 74365 99719
0 34156 7 1 2 95598 34155
0 34157 7 1 2 99772 34156
0 34158 5 1 1 34157
0 34159 7 1 2 34151 34158
0 34160 5 1 1 34159
0 34161 7 1 2 64276 34160
0 34162 5 1 1 34161
0 34163 7 1 2 84590 99210
0 34164 7 3 2 62150 99316
0 34165 7 2 2 79451 94369
0 34166 7 1 2 99774 99777
0 34167 7 1 2 34163 34166
0 34168 5 1 1 34167
0 34169 7 1 2 34162 34168
0 34170 5 1 1 34169
0 34171 7 1 2 64964 34170
0 34172 5 1 1 34171
0 34173 7 1 2 74329 76780
0 34174 7 2 2 94370 34173
0 34175 7 7 2 93857 99749
0 34176 7 1 2 3733 10374
0 34177 5 1 1 34176
0 34178 7 1 2 99781 34177
0 34179 5 1 1 34178
0 34180 7 2 2 86973 72347
0 34181 5 1 1 99788
0 34182 7 4 2 67800 69391
0 34183 7 1 2 90996 99790
0 34184 7 1 2 99789 34183
0 34185 5 1 1 34184
0 34186 7 1 2 34179 34185
0 34187 5 1 1 34186
0 34188 7 1 2 99779 34187
0 34189 5 1 1 34188
0 34190 7 1 2 34172 34189
0 34191 5 1 1 34190
0 34192 7 1 2 70100 34191
0 34193 5 1 1 34192
0 34194 7 1 2 99689 99342
0 34195 7 1 2 99758 34194
0 34196 5 1 1 34195
0 34197 7 1 2 98423 99707
0 34198 5 1 1 34197
0 34199 7 1 2 34154 34198
0 34200 5 1 1 34199
0 34201 7 1 2 73831 99720
0 34202 7 1 2 34200 34201
0 34203 5 1 1 34202
0 34204 7 1 2 34196 34203
0 34205 5 1 1 34204
0 34206 7 5 2 61622 64277
0 34207 7 1 2 75807 99794
0 34208 7 1 2 81859 34207
0 34209 7 1 2 34205 34208
0 34210 5 1 1 34209
0 34211 7 1 2 34193 34210
0 34212 5 1 1 34211
0 34213 7 1 2 98393 34212
0 34214 5 1 1 34213
0 34215 7 1 2 76385 98883
0 34216 5 1 1 34215
0 34217 7 2 2 98536 98911
0 34218 7 1 2 84277 99799
0 34219 5 1 1 34218
0 34220 7 1 2 34216 34219
0 34221 5 1 1 34220
0 34222 7 2 2 65174 34221
0 34223 5 1 1 99801
0 34224 7 2 2 76895 94371
0 34225 7 1 2 66124 74330
0 34226 7 1 2 99803 34225
0 34227 5 1 1 34226
0 34228 7 1 2 34223 34227
0 34229 5 1 1 34228
0 34230 7 1 2 63372 34229
0 34231 5 1 1 34230
0 34232 7 1 2 81591 81710
0 34233 7 1 2 99804 34232
0 34234 5 1 1 34233
0 34235 7 1 2 34231 34234
0 34236 5 1 1 34235
0 34237 7 1 2 78281 34236
0 34238 5 1 1 34237
0 34239 7 7 2 64278 69823
0 34240 7 1 2 86379 87837
0 34241 7 1 2 99805 34240
0 34242 7 1 2 92161 99560
0 34243 7 1 2 34241 34242
0 34244 5 1 1 34243
0 34245 7 1 2 34238 34244
0 34246 5 1 1 34245
0 34247 7 1 2 63184 34246
0 34248 5 1 1 34247
0 34249 7 1 2 81740 97501
0 34250 7 1 2 99802 34249
0 34251 5 1 1 34250
0 34252 7 1 2 34248 34251
0 34253 5 1 1 34252
0 34254 7 1 2 82280 34253
0 34255 5 1 1 34254
0 34256 7 2 2 73470 76386
0 34257 7 2 2 66125 66765
0 34258 7 2 2 94372 99814
0 34259 7 1 2 81741 79788
0 34260 7 1 2 99816 34259
0 34261 7 1 2 99812 34260
0 34262 5 1 1 34261
0 34263 7 1 2 34255 34262
0 34264 5 1 1 34263
0 34265 7 1 2 90710 34264
0 34266 5 1 1 34265
0 34267 7 2 2 79133 78732
0 34268 5 1 1 99818
0 34269 7 1 2 97167 34268
0 34270 5 1 1 34269
0 34271 7 2 2 93786 34270
0 34272 7 1 2 66766 99820
0 34273 5 1 1 34272
0 34274 7 5 2 64767 78605
0 34275 7 1 2 79778 93758
0 34276 7 1 2 99822 34275
0 34277 5 1 1 34276
0 34278 7 1 2 34273 34277
0 34279 5 1 1 34278
0 34280 7 1 2 62868 34279
0 34281 5 1 1 34280
0 34282 7 7 2 63021 64768
0 34283 7 1 2 98086 99827
0 34284 7 1 2 78742 34283
0 34285 5 1 1 34284
0 34286 7 1 2 34281 34285
0 34287 5 1 1 34286
0 34288 7 2 2 95166 98590
0 34289 5 1 1 99834
0 34290 7 2 2 65795 97434
0 34291 7 1 2 94767 99836
0 34292 5 1 1 34291
0 34293 7 1 2 34289 34292
0 34294 5 1 1 34293
0 34295 7 1 2 97368 34294
0 34296 7 1 2 34287 34295
0 34297 5 1 1 34296
0 34298 7 1 2 73471 83351
0 34299 5 1 1 34298
0 34300 7 3 2 86929 78850
0 34301 5 1 1 99838
0 34302 7 1 2 65796 99839
0 34303 5 1 1 34302
0 34304 7 1 2 34299 34303
0 34305 5 1 1 34304
0 34306 7 1 2 88817 34305
0 34307 5 1 1 34306
0 34308 7 4 2 81129 83521
0 34309 5 1 1 99841
0 34310 7 1 2 27060 34309
0 34311 5 1 1 34310
0 34312 7 1 2 72348 82470
0 34313 7 1 2 34311 34312
0 34314 5 1 1 34313
0 34315 7 1 2 34307 34314
0 34316 5 1 1 34315
0 34317 7 5 2 65462 93787
0 34318 7 1 2 99845 98978
0 34319 7 1 2 34316 34318
0 34320 5 1 1 34319
0 34321 7 1 2 34297 34320
0 34322 5 1 1 34321
0 34323 7 1 2 66126 34322
0 34324 5 1 1 34323
0 34325 7 2 2 63022 79134
0 34326 7 1 2 93085 95303
0 34327 7 1 2 98087 34326
0 34328 7 1 2 99850 34327
0 34329 5 1 1 34328
0 34330 7 3 2 90878 93019
0 34331 5 1 1 99852
0 34332 7 1 2 93614 34331
0 34333 5 3 1 34332
0 34334 7 1 2 97164 99855
0 34335 5 1 1 34334
0 34336 7 1 2 99853 99819
0 34337 5 1 1 34336
0 34338 7 1 2 34335 34337
0 34339 5 1 1 34338
0 34340 7 1 2 66767 93788
0 34341 7 1 2 34339 34340
0 34342 5 1 1 34341
0 34343 7 1 2 34329 34342
0 34344 5 1 1 34343
0 34345 7 1 2 72459 34344
0 34346 5 1 1 34345
0 34347 7 1 2 71701 90879
0 34348 7 1 2 98591 34347
0 34349 7 1 2 99821 34348
0 34350 5 1 1 34349
0 34351 7 1 2 34346 34350
0 34352 5 1 1 34351
0 34353 7 1 2 62869 97710
0 34354 7 1 2 34352 34353
0 34355 5 1 1 34354
0 34356 7 1 2 34324 34355
0 34357 5 1 1 34356
0 34358 7 1 2 63373 34357
0 34359 5 1 1 34358
0 34360 7 1 2 61296 99856
0 34361 5 1 1 34360
0 34362 7 1 2 93025 97369
0 34363 5 1 1 34362
0 34364 7 1 2 34361 34363
0 34365 5 1 1 34364
0 34366 7 2 2 63588 83352
0 34367 5 1 1 99858
0 34368 7 1 2 6113 34367
0 34369 5 1 1 34368
0 34370 7 1 2 99119 34369
0 34371 7 1 2 34365 34370
0 34372 5 1 1 34371
0 34373 7 6 2 69592 79937
0 34374 7 1 2 96919 99860
0 34375 5 1 1 34374
0 34376 7 1 2 83353 95646
0 34377 5 1 1 34376
0 34378 7 1 2 34375 34377
0 34379 5 1 1 34378
0 34380 7 1 2 75781 97306
0 34381 7 1 2 34379 34380
0 34382 5 1 1 34381
0 34383 7 1 2 34372 34382
0 34384 5 1 1 34383
0 34385 7 1 2 65797 34384
0 34386 5 1 1 34385
0 34387 7 3 2 77684 93858
0 34388 7 4 2 65463 74366
0 34389 7 1 2 64279 92117
0 34390 7 1 2 90576 34389
0 34391 7 1 2 99869 34390
0 34392 7 1 2 99866 34391
0 34393 5 1 1 34392
0 34394 7 1 2 34386 34393
0 34395 5 1 1 34394
0 34396 7 1 2 70101 34395
0 34397 5 1 1 34396
0 34398 7 1 2 79779 97711
0 34399 7 1 2 84852 34398
0 34400 7 1 2 97375 34399
0 34401 5 1 1 34400
0 34402 7 1 2 34397 34401
0 34403 5 1 1 34402
0 34404 7 1 2 68205 99096
0 34405 7 1 2 34403 34404
0 34406 5 1 1 34405
0 34407 7 1 2 34359 34406
0 34408 5 1 1 34407
0 34409 7 1 2 69392 34408
0 34410 5 1 1 34409
0 34411 7 1 2 86334 97449
0 34412 7 2 2 98873 34411
0 34413 5 1 1 99873
0 34414 7 1 2 67002 99874
0 34415 5 1 1 34414
0 34416 7 2 2 98537 97672
0 34417 5 2 1 99875
0 34418 7 2 2 66237 99364
0 34419 7 1 2 98036 99625
0 34420 7 1 2 99879 34419
0 34421 5 1 1 34420
0 34422 7 1 2 99877 34421
0 34423 5 1 1 34422
0 34424 7 1 2 65175 34423
0 34425 5 1 1 34424
0 34426 7 1 2 94967 98080
0 34427 5 1 1 34426
0 34428 7 1 2 34425 34427
0 34429 5 1 1 34428
0 34430 7 1 2 78282 34429
0 34431 5 1 1 34430
0 34432 7 1 2 34415 34431
0 34433 5 1 1 34432
0 34434 7 1 2 67482 34433
0 34435 5 1 1 34434
0 34436 7 1 2 83341 76373
0 34437 7 1 2 86290 34436
0 34438 7 1 2 97673 34437
0 34439 5 1 1 34438
0 34440 7 1 2 34435 34439
0 34441 5 1 1 34440
0 34442 7 1 2 87094 87790
0 34443 7 1 2 34441 34442
0 34444 5 1 1 34443
0 34445 7 1 2 87415 99876
0 34446 5 1 1 34445
0 34447 7 1 2 67801 97772
0 34448 7 1 2 98207 99626
0 34449 7 2 2 34447 34448
0 34450 7 1 2 93252 99881
0 34451 5 1 1 34450
0 34452 7 1 2 34446 34451
0 34453 5 1 1 34452
0 34454 7 1 2 83138 34453
0 34455 5 1 1 34454
0 34456 7 1 2 90772 98160
0 34457 7 2 2 91698 34456
0 34458 7 2 2 98494 97459
0 34459 7 1 2 99883 99885
0 34460 5 1 1 34459
0 34461 7 1 2 34460 34413
0 34462 5 1 1 34461
0 34463 7 1 2 84799 34462
0 34464 5 1 1 34463
0 34465 7 1 2 34455 34464
0 34466 5 1 1 34465
0 34467 7 1 2 87728 34466
0 34468 5 1 1 34467
0 34469 7 1 2 99861 98061
0 34470 5 1 1 34469
0 34471 7 1 2 88099 99806
0 34472 7 1 2 98874 34471
0 34473 5 1 1 34472
0 34474 7 1 2 34470 34473
0 34475 5 1 1 34474
0 34476 7 1 2 94875 98867
0 34477 7 1 2 34475 34476
0 34478 5 1 1 34477
0 34479 7 1 2 34468 34478
0 34480 7 1 2 34444 34479
0 34481 5 1 1 34480
0 34482 7 1 2 82281 34481
0 34483 5 1 1 34482
0 34484 7 1 2 63185 34483
0 34485 7 1 2 34410 34484
0 34486 5 1 1 34485
0 34487 7 1 2 74331 83630
0 34488 5 1 1 34487
0 34489 7 1 2 4348 34488
0 34490 5 1 1 34489
0 34491 7 1 2 83065 34490
0 34492 5 1 1 34491
0 34493 7 1 2 85022 92084
0 34494 5 1 1 34493
0 34495 7 1 2 34492 34494
0 34496 5 1 1 34495
0 34497 7 1 2 73472 34496
0 34498 5 1 1 34497
0 34499 7 2 2 86870 73832
0 34500 7 1 2 82632 82401
0 34501 7 1 2 99887 34500
0 34502 5 1 1 34501
0 34503 7 1 2 34498 34502
0 34504 5 1 1 34503
0 34505 7 1 2 87729 34504
0 34506 5 1 1 34505
0 34507 7 1 2 83902 99638
0 34508 5 1 1 34507
0 34509 7 1 2 86142 87838
0 34510 7 1 2 99480 34509
0 34511 5 1 1 34510
0 34512 7 1 2 34508 34511
0 34513 5 1 1 34512
0 34514 7 1 2 92710 34513
0 34515 5 1 1 34514
0 34516 7 1 2 34506 34515
0 34517 5 1 1 34516
0 34518 7 1 2 65464 34517
0 34519 5 1 1 34518
0 34520 7 1 2 66768 89189
0 34521 5 1 1 34520
0 34522 7 2 2 83066 83987
0 34523 5 1 1 99889
0 34524 7 1 2 34521 34523
0 34525 5 3 1 34524
0 34526 7 1 2 99891 99552
0 34527 5 1 1 34526
0 34528 7 1 2 34519 34527
0 34529 5 1 1 34528
0 34530 7 1 2 98012 34529
0 34531 5 1 1 34530
0 34532 7 1 2 70396 99639
0 34533 5 1 1 34532
0 34534 7 1 2 73100 99544
0 34535 5 1 1 34534
0 34536 7 1 2 34533 34535
0 34537 5 1 1 34536
0 34538 7 1 2 63589 34537
0 34539 5 1 1 34538
0 34540 7 3 2 69227 73125
0 34541 7 1 2 66127 75858
0 34542 7 1 2 99894 34541
0 34543 5 1 1 34542
0 34544 7 1 2 34539 34543
0 34545 5 1 1 34544
0 34546 7 1 2 83139 83988
0 34547 7 1 2 34545 34546
0 34548 5 1 1 34547
0 34549 7 3 2 74367 72460
0 34550 7 1 2 85191 84423
0 34551 7 1 2 97082 34550
0 34552 7 1 2 99897 34551
0 34553 5 1 1 34552
0 34554 7 1 2 34548 34553
0 34555 5 1 1 34554
0 34556 7 1 2 98196 34555
0 34557 5 1 1 34556
0 34558 7 1 2 93737 94890
0 34559 7 3 2 67868 92959
0 34560 7 1 2 95925 99300
0 34561 7 1 2 99900 34560
0 34562 7 1 2 34558 34561
0 34563 5 1 1 34562
0 34564 7 1 2 34557 34563
0 34565 5 1 1 34564
0 34566 7 1 2 61372 34565
0 34567 5 1 1 34566
0 34568 7 1 2 34531 34567
0 34569 5 1 1 34568
0 34570 7 1 2 70102 34569
0 34571 5 1 1 34570
0 34572 7 2 2 62605 64280
0 34573 7 3 2 69228 99903
0 34574 7 1 2 99905 99571
0 34575 5 1 1 34574
0 34576 7 3 2 66128 76713
0 34577 7 2 2 94373 98618
0 34578 7 1 2 99908 99911
0 34579 5 1 1 34578
0 34580 7 1 2 34575 34579
0 34581 5 1 1 34580
0 34582 7 1 2 65176 34581
0 34583 5 1 1 34582
0 34584 7 4 2 99365 97629
0 34585 7 3 2 64375 70103
0 34586 7 1 2 76714 99917
0 34587 7 1 2 99913 34586
0 34588 5 1 1 34587
0 34589 7 1 2 34583 34588
0 34590 5 1 1 34589
0 34591 7 1 2 68433 34590
0 34592 5 1 1 34591
0 34593 7 2 2 65177 98884
0 34594 7 1 2 84695 99366
0 34595 7 1 2 99920 34594
0 34596 5 1 1 34595
0 34597 7 1 2 34592 34596
0 34598 5 1 1 34597
0 34599 7 1 2 63374 34598
0 34600 5 1 1 34599
0 34601 7 2 2 86480 94374
0 34602 7 1 2 92641 92693
0 34603 7 1 2 99922 34602
0 34604 5 1 1 34603
0 34605 7 1 2 34600 34604
0 34606 5 1 1 34605
0 34607 7 1 2 76998 92730
0 34608 7 1 2 34606 34607
0 34609 5 1 1 34608
0 34610 7 5 2 77129 80299
0 34611 7 1 2 82992 93909
0 34612 7 1 2 99924 34611
0 34613 7 1 2 99563 34612
0 34614 5 1 1 34613
0 34615 7 1 2 34609 34614
0 34616 5 1 1 34615
0 34617 7 1 2 93789 34616
0 34618 5 1 1 34617
0 34619 7 2 2 76387 98013
0 34620 5 1 1 99929
0 34621 7 1 2 98868 99930
0 34622 5 1 1 34621
0 34623 7 3 2 91343 81873
0 34624 7 1 2 99931 99800
0 34625 5 1 1 34624
0 34626 7 1 2 34622 34625
0 34627 5 1 1 34626
0 34628 7 1 2 91056 34627
0 34629 5 1 1 34628
0 34630 7 1 2 99878 34620
0 34631 5 1 1 34630
0 34632 7 1 2 81458 34631
0 34633 5 1 1 34632
0 34634 7 2 2 83067 88176
0 34635 7 1 2 64281 98538
0 34636 7 1 2 99934 34635
0 34637 5 1 1 34636
0 34638 7 1 2 34633 34637
0 34639 5 1 1 34638
0 34640 7 1 2 73473 34639
0 34641 5 1 1 34640
0 34642 7 2 2 90980 98200
0 34643 7 1 2 99120 99936
0 34644 7 1 2 96123 34643
0 34645 5 1 1 34644
0 34646 7 1 2 34641 34645
0 34647 5 1 1 34646
0 34648 7 1 2 87730 34647
0 34649 5 1 1 34648
0 34650 7 2 2 73126 97674
0 34651 5 1 1 99938
0 34652 7 1 2 83140 99939
0 34653 5 1 1 34652
0 34654 7 2 2 71536 86060
0 34655 5 3 1 99940
0 34656 7 1 2 73611 77319
0 34657 5 1 1 34656
0 34658 7 1 2 99942 34657
0 34659 5 3 1 34658
0 34660 7 1 2 81459 98014
0 34661 7 1 2 99945 34660
0 34662 5 1 1 34661
0 34663 7 1 2 34653 34662
0 34664 5 1 1 34663
0 34665 7 1 2 68434 34664
0 34666 5 1 1 34665
0 34667 7 1 2 71737 90799
0 34668 5 1 1 34667
0 34669 7 1 2 84800 78399
0 34670 5 1 1 34669
0 34671 7 1 2 34668 34670
0 34672 5 3 1 34671
0 34673 7 1 2 99164 99886
0 34674 7 1 2 99948 34673
0 34675 5 1 1 34674
0 34676 7 1 2 34666 34675
0 34677 5 1 1 34676
0 34678 7 1 2 99545 34677
0 34679 5 1 1 34678
0 34680 7 1 2 34649 34679
0 34681 5 1 1 34680
0 34682 7 1 2 79645 34681
0 34683 5 1 1 34682
0 34684 7 1 2 34629 34683
0 34685 5 1 1 34684
0 34686 7 1 2 65178 34685
0 34687 5 1 1 34686
0 34688 7 1 2 68027 34687
0 34689 7 1 2 34618 34688
0 34690 7 1 2 34571 34689
0 34691 5 1 1 34690
0 34692 7 1 2 34486 34691
0 34693 5 1 1 34692
0 34694 7 1 2 34266 34693
0 34695 5 1 1 34694
0 34696 7 1 2 61623 34695
0 34697 5 1 1 34696
0 34698 7 3 2 75655 97738
0 34699 7 1 2 74368 99951
0 34700 5 2 1 34699
0 34701 7 2 2 73474 98936
0 34702 5 1 1 99956
0 34703 7 1 2 63590 99957
0 34704 5 1 1 34703
0 34705 7 1 2 99954 34704
0 34706 5 1 1 34705
0 34707 7 1 2 88194 34706
0 34708 5 1 1 34707
0 34709 7 3 2 69123 74470
0 34710 7 1 2 80413 87683
0 34711 7 1 2 96061 34710
0 34712 7 1 2 99958 34711
0 34713 5 1 1 34712
0 34714 7 1 2 34708 34713
0 34715 5 1 1 34714
0 34716 7 1 2 64540 34715
0 34717 5 1 1 34716
0 34718 7 2 2 63591 93933
0 34719 7 1 2 98885 99961
0 34720 5 1 1 34719
0 34721 7 1 2 99955 34720
0 34722 5 1 1 34721
0 34723 7 1 2 98929 34722
0 34724 5 1 1 34723
0 34725 7 1 2 34717 34724
0 34726 5 1 1 34725
0 34727 7 1 2 69824 34726
0 34728 5 1 1 34727
0 34729 7 9 2 66129 67003
0 34730 7 2 2 94758 99963
0 34731 7 1 2 97083 99972
0 34732 7 1 2 94655 34731
0 34733 5 1 1 34732
0 34734 7 1 2 34728 34733
0 34735 5 1 1 34734
0 34736 7 1 2 65465 34735
0 34737 5 1 1 34736
0 34738 7 1 2 81495 17360
0 34739 5 3 1 34738
0 34740 7 1 2 66518 99974
0 34741 5 1 1 34740
0 34742 7 1 2 18283 34741
0 34743 5 1 1 34742
0 34744 7 2 2 79698 97712
0 34745 7 1 2 96071 99898
0 34746 7 1 2 99977 34745
0 34747 7 1 2 34743 34746
0 34748 5 1 1 34747
0 34749 7 1 2 34737 34748
0 34750 5 1 1 34749
0 34751 7 1 2 70104 34750
0 34752 5 1 1 34751
0 34753 7 1 2 78679 86651
0 34754 7 1 2 97615 34753
0 34755 7 1 2 73127 34754
0 34756 7 1 2 98246 34755
0 34757 5 1 1 34756
0 34758 7 1 2 34752 34757
0 34759 5 1 1 34758
0 34760 7 1 2 83141 34759
0 34761 5 1 1 34760
0 34762 7 3 2 66130 95189
0 34763 7 1 2 86284 97379
0 34764 7 1 2 99979 34763
0 34765 7 1 2 99813 34764
0 34766 5 1 1 34765
0 34767 7 1 2 75898 95150
0 34768 7 1 2 99690 34767
0 34769 7 1 2 96630 98539
0 34770 7 1 2 34768 34769
0 34771 5 1 1 34770
0 34772 7 1 2 98832 99778
0 34773 7 1 2 76388 34772
0 34774 5 1 1 34773
0 34775 7 1 2 34771 34774
0 34776 5 1 1 34775
0 34777 7 1 2 61903 92069
0 34778 7 1 2 34776 34777
0 34779 5 1 1 34778
0 34780 7 1 2 34766 34779
0 34781 5 1 1 34780
0 34782 7 1 2 65179 85423
0 34783 7 1 2 34781 34782
0 34784 5 1 1 34783
0 34785 7 1 2 34761 34784
0 34786 5 1 1 34785
0 34787 7 1 2 90711 34786
0 34788 5 1 1 34787
0 34789 7 1 2 92826 98547
0 34790 5 1 1 34789
0 34791 7 1 2 62973 98555
0 34792 5 1 1 34791
0 34793 7 1 2 34790 34792
0 34794 5 4 1 34793
0 34795 7 6 2 61373 67709
0 34796 7 2 2 64541 99986
0 34797 7 1 2 66131 99780
0 34798 5 1 1 34797
0 34799 7 2 2 94768 96450
0 34800 7 1 2 61297 63592
0 34801 7 1 2 71738 34800
0 34802 7 1 2 99994 34801
0 34803 5 1 1 34802
0 34804 7 1 2 34798 34803
0 34805 5 1 1 34804
0 34806 7 1 2 99992 34805
0 34807 5 1 1 34806
0 34808 7 33 2 66238 69393
0 34809 7 1 2 74391 97713
0 34810 7 1 2 99895 34809
0 34811 5 1 1 34810
0 34812 7 5 2 62151 69124
0 34813 7 1 2 83199 100029
0 34814 7 1 2 98336 34813
0 34815 5 1 1 34814
0 34816 7 1 2 34811 34815
0 34817 5 1 1 34816
0 34818 7 1 2 64965 34817
0 34819 5 1 1 34818
0 34820 7 5 2 94375 99964
0 34821 7 1 2 73833 88144
0 34822 7 1 2 100034 34821
0 34823 5 1 1 34822
0 34824 7 1 2 34819 34823
0 34825 5 1 1 34824
0 34826 7 1 2 99996 34825
0 34827 5 1 1 34826
0 34828 7 1 2 34807 34827
0 34829 5 1 1 34828
0 34830 7 1 2 86974 34829
0 34831 5 1 1 34830
0 34832 7 4 2 79367 92192
0 34833 5 1 1 100039
0 34834 7 4 2 87940 97630
0 34835 7 1 2 90301 100043
0 34836 5 1 1 34835
0 34837 7 2 2 84278 93910
0 34838 7 1 2 74436 97916
0 34839 7 1 2 100047 34838
0 34840 5 1 1 34839
0 34841 7 1 2 34836 34840
0 34842 5 1 1 34841
0 34843 7 1 2 100040 34842
0 34844 5 1 1 34843
0 34845 7 1 2 34831 34844
0 34846 5 1 1 34845
0 34847 7 1 2 70105 34846
0 34848 5 1 1 34847
0 34849 7 2 2 90865 98730
0 34850 7 1 2 73075 73834
0 34851 7 1 2 100049 34850
0 34852 5 1 1 34851
0 34853 7 2 2 99987 99687
0 34854 5 1 1 100051
0 34855 7 1 2 67004 100052
0 34856 5 1 1 34855
0 34857 7 1 2 63593 34856
0 34858 5 1 1 34857
0 34859 7 2 2 66239 72920
0 34860 7 1 2 92312 100053
0 34861 5 1 1 34860
0 34862 7 1 2 34861 34854
0 34863 5 2 1 34862
0 34864 7 1 2 70397 100055
0 34865 7 1 2 34858 34864
0 34866 5 1 1 34865
0 34867 7 1 2 34852 34866
0 34868 5 1 1 34867
0 34869 7 1 2 81860 98923
0 34870 7 1 2 34868 34869
0 34871 5 1 1 34870
0 34872 7 1 2 34848 34871
0 34873 5 1 1 34872
0 34874 7 1 2 99982 34873
0 34875 5 1 1 34874
0 34876 7 1 2 34788 34875
0 34877 7 1 2 34697 34876
0 34878 7 1 2 34214 34877
0 34879 7 1 2 34113 34878
0 34880 5 1 1 34879
0 34881 7 1 2 73026 34880
0 34882 5 1 1 34881
0 34883 7 2 2 76210 99343
0 34884 7 1 2 100057 98203
0 34885 5 1 1 34884
0 34886 7 1 2 93203 93520
0 34887 5 1 1 34886
0 34888 7 1 2 34885 34887
0 34889 5 1 1 34888
0 34890 7 1 2 62152 34889
0 34891 5 1 1 34890
0 34892 7 1 2 78792 97466
0 34893 7 1 2 99641 34892
0 34894 5 1 1 34893
0 34895 7 1 2 34891 34894
0 34896 5 1 1 34895
0 34897 7 1 2 64966 34896
0 34898 5 1 1 34897
0 34899 7 1 2 72229 96540
0 34900 7 1 2 97444 34899
0 34901 7 1 2 90712 34900
0 34902 5 1 1 34901
0 34903 7 1 2 34898 34902
0 34904 5 1 1 34903
0 34905 7 1 2 69394 34904
0 34906 5 1 1 34905
0 34907 7 1 2 82282 93594
0 34908 7 1 2 88039 34907
0 34909 7 1 2 99846 34908
0 34910 5 1 1 34909
0 34911 7 1 2 34906 34910
0 34912 5 1 1 34911
0 34913 7 1 2 84407 34912
0 34914 5 1 1 34913
0 34915 7 1 2 83956 84591
0 34916 7 1 2 88040 34915
0 34917 7 1 2 93204 34916
0 34918 5 1 1 34917
0 34919 7 1 2 34914 34918
0 34920 5 1 1 34919
0 34921 7 1 2 73027 34920
0 34922 5 1 1 34921
0 34923 7 1 2 90262 98990
0 34924 5 1 1 34923
0 34925 7 1 2 63594 76739
0 34926 7 4 2 82851 79542
0 34927 5 1 1 100059
0 34928 7 1 2 86267 100060
0 34929 7 1 2 34925 34928
0 34930 5 1 1 34929
0 34931 7 1 2 34924 34930
0 34932 5 1 1 34931
0 34933 7 1 2 64967 34932
0 34934 5 1 1 34933
0 34935 7 3 2 69395 88124
0 34936 7 2 2 87405 94323
0 34937 7 1 2 100063 100066
0 34938 5 1 1 34937
0 34939 7 1 2 32588 34938
0 34940 5 1 1 34939
0 34941 7 1 2 88041 34940
0 34942 5 1 1 34941
0 34943 7 1 2 34934 34942
0 34944 5 1 1 34943
0 34945 7 1 2 65798 34944
0 34946 5 1 1 34945
0 34947 7 1 2 88639 77090
0 34948 7 1 2 72412 34947
0 34949 7 1 2 85884 95391
0 34950 7 1 2 34948 34949
0 34951 5 1 1 34950
0 34952 7 1 2 34946 34951
0 34953 5 1 1 34952
0 34954 7 1 2 90713 34953
0 34955 5 1 1 34954
0 34956 7 1 2 79135 75878
0 34957 7 3 2 68435 64542
0 34958 7 1 2 97601 100068
0 34959 7 1 2 34956 34958
0 34960 7 1 2 93790 34959
0 34961 7 1 2 94201 34960
0 34962 5 1 1 34961
0 34963 7 1 2 34955 34962
0 34964 5 1 1 34963
0 34965 7 1 2 64376 34964
0 34966 5 1 1 34965
0 34967 7 1 2 34922 34966
0 34968 5 1 1 34967
0 34969 7 1 2 69125 34968
0 34970 5 1 1 34969
0 34971 7 6 2 69229 97647
0 34972 7 4 2 66519 99828
0 34973 5 3 1 100077
0 34974 7 1 2 86930 99105
0 34975 5 1 1 34974
0 34976 7 1 2 100081 34975
0 34977 5 2 1 34976
0 34978 7 1 2 61374 100084
0 34979 5 1 1 34978
0 34980 7 1 2 86931 99032
0 34981 5 1 1 34980
0 34982 7 1 2 34979 34981
0 34983 5 5 1 34982
0 34984 7 1 2 100086 98965
0 34985 5 1 1 34984
0 34986 7 10 2 92193 99829
0 34987 7 1 2 80371 100091
0 34988 5 1 1 34987
0 34989 7 1 2 34985 34988
0 34990 5 1 1 34989
0 34991 7 1 2 62153 34990
0 34992 5 1 1 34991
0 34993 7 1 2 74369 80357
0 34994 7 1 2 100087 34993
0 34995 5 1 1 34994
0 34996 7 1 2 34992 34995
0 34997 5 1 1 34996
0 34998 7 1 2 62606 34997
0 34999 5 1 1 34998
0 35000 7 1 2 78387 100088
0 35001 5 1 1 35000
0 35002 7 2 2 90607 80838
0 35003 7 1 2 82589 100101
0 35004 5 1 1 35003
0 35005 7 1 2 35001 35004
0 35006 5 1 1 35005
0 35007 7 1 2 62154 35006
0 35008 5 1 1 35007
0 35009 7 1 2 67005 96340
0 35010 7 1 2 100102 35009
0 35011 5 1 1 35010
0 35012 7 1 2 35008 35011
0 35013 5 1 1 35012
0 35014 7 1 2 71595 35013
0 35015 5 1 1 35014
0 35016 7 1 2 34999 35015
0 35017 5 1 1 35016
0 35018 7 1 2 69396 35017
0 35019 5 1 1 35018
0 35020 7 2 2 79368 99202
0 35021 7 1 2 97269 98698
0 35022 7 1 2 100103 35021
0 35023 7 1 2 74418 35022
0 35024 5 1 1 35023
0 35025 7 1 2 35019 35024
0 35026 5 1 1 35025
0 35027 7 1 2 64968 35026
0 35028 5 1 1 35027
0 35029 7 1 2 90293 90608
0 35030 7 1 2 99250 35029
0 35031 5 1 1 35030
0 35032 7 1 2 35028 35031
0 35033 5 1 1 35032
0 35034 7 1 2 100071 35033
0 35035 5 1 1 35034
0 35036 7 1 2 34970 35035
0 35037 5 1 1 35036
0 35038 7 1 2 70106 35037
0 35039 5 1 1 35038
0 35040 7 3 2 62155 93000
0 35041 7 2 2 93502 94405
0 35042 7 1 2 100105 100108
0 35043 5 1 1 35042
0 35044 7 5 2 63023 69230
0 35045 7 2 2 94633 100110
0 35046 7 1 2 72921 100115
0 35047 7 1 2 80358 35046
0 35048 5 1 1 35047
0 35049 7 1 2 35043 35048
0 35050 5 1 1 35049
0 35051 7 1 2 68436 35050
0 35052 5 1 1 35051
0 35053 7 1 2 75879 99627
0 35054 7 1 2 100109 35053
0 35055 5 1 1 35054
0 35056 7 1 2 75264 98645
0 35057 7 1 2 92740 99234
0 35058 7 1 2 35056 35057
0 35059 5 1 1 35058
0 35060 7 1 2 35055 35059
0 35061 7 1 2 35052 35060
0 35062 5 1 1 35061
0 35063 7 1 2 61375 35062
0 35064 5 1 1 35063
0 35065 7 5 2 63024 64377
0 35066 7 1 2 99750 100117
0 35067 7 1 2 98836 35066
0 35068 7 1 2 83717 35067
0 35069 7 1 2 95417 35068
0 35070 5 1 1 35069
0 35071 7 1 2 35064 35070
0 35072 5 1 1 35071
0 35073 7 1 2 69825 35072
0 35074 5 1 1 35073
0 35075 7 5 2 61376 62156
0 35076 7 1 2 100122 100116
0 35077 7 1 2 98427 35076
0 35078 5 1 1 35077
0 35079 7 1 2 35074 35078
0 35080 5 1 1 35079
0 35081 7 1 2 79753 97602
0 35082 7 1 2 35080 35081
0 35083 5 1 1 35082
0 35084 7 1 2 66132 35083
0 35085 7 1 2 35039 35084
0 35086 5 1 1 35085
0 35087 7 2 2 79369 99224
0 35088 7 2 2 93194 100127
0 35089 7 1 2 98871 100129
0 35090 5 1 1 35089
0 35091 7 1 2 64969 98365
0 35092 5 1 1 35091
0 35093 7 1 2 79229 88145
0 35094 7 1 2 99857 35093
0 35095 5 1 1 35094
0 35096 7 1 2 35092 35095
0 35097 5 1 1 35096
0 35098 7 1 2 62157 35097
0 35099 5 1 1 35098
0 35100 7 1 2 31633 35099
0 35101 5 1 1 35100
0 35102 7 1 2 90263 35101
0 35103 5 1 1 35102
0 35104 7 1 2 35090 35103
0 35105 5 1 1 35104
0 35106 7 1 2 90609 35105
0 35107 5 1 1 35106
0 35108 7 4 2 67869 69231
0 35109 7 2 2 79452 100131
0 35110 7 1 2 97603 97773
0 35111 7 1 2 100135 35110
0 35112 7 1 2 98431 35111
0 35113 5 1 1 35112
0 35114 7 1 2 35107 35113
0 35115 5 1 1 35114
0 35116 7 1 2 65180 35115
0 35117 5 1 1 35116
0 35118 7 2 2 62607 97582
0 35119 7 1 2 96169 100137
0 35120 7 1 2 99715 35119
0 35121 5 1 1 35120
0 35122 7 6 2 62974 63595
0 35123 7 2 2 97904 100139
0 35124 7 1 2 80940 81537
0 35125 7 1 2 100145 35124
0 35126 5 1 1 35125
0 35127 7 1 2 35121 35126
0 35128 5 1 1 35127
0 35129 7 1 2 78552 35128
0 35130 5 1 1 35129
0 35131 7 1 2 70735 91280
0 35132 7 1 2 93172 35131
0 35133 7 1 2 95808 98540
0 35134 7 1 2 35132 35133
0 35135 5 1 1 35134
0 35136 7 1 2 35130 35135
0 35137 5 1 1 35136
0 35138 7 1 2 69232 35137
0 35139 5 1 1 35138
0 35140 7 2 2 83449 99899
0 35141 7 2 2 62870 93595
0 35142 7 1 2 91518 100149
0 35143 7 1 2 100147 35142
0 35144 5 1 1 35143
0 35145 7 1 2 35139 35144
0 35146 5 1 1 35145
0 35147 7 1 2 93791 35146
0 35148 5 1 1 35147
0 35149 7 5 2 69233 90714
0 35150 7 2 2 92280 97277
0 35151 5 1 1 100156
0 35152 7 1 2 63596 100157
0 35153 5 1 1 35152
0 35154 7 3 2 79453 80730
0 35155 7 1 2 74370 71537
0 35156 7 1 2 100158 35155
0 35157 5 1 1 35156
0 35158 7 1 2 35153 35157
0 35159 5 1 1 35158
0 35160 7 1 2 78553 35159
0 35161 5 1 1 35160
0 35162 7 1 2 75440 91998
0 35163 7 1 2 100159 35162
0 35164 5 1 1 35163
0 35165 7 1 2 35161 35164
0 35166 5 1 1 35165
0 35167 7 1 2 100151 35166
0 35168 5 1 1 35167
0 35169 7 4 2 90610 93596
0 35170 7 1 2 78606 99530
0 35171 5 1 1 35170
0 35172 7 1 2 9873 35171
0 35173 5 1 1 35172
0 35174 7 1 2 83957 35173
0 35175 5 1 1 35174
0 35176 7 2 2 78607 73835
0 35177 5 2 1 100165
0 35178 7 1 2 98255 100166
0 35179 5 1 1 35178
0 35180 7 1 2 35175 35179
0 35181 5 1 1 35180
0 35182 7 1 2 100161 35181
0 35183 5 1 1 35182
0 35184 7 1 2 35168 35183
0 35185 5 1 1 35184
0 35186 7 1 2 70398 35185
0 35187 5 1 1 35186
0 35188 7 1 2 78744 100167
0 35189 5 1 1 35188
0 35190 7 1 2 90312 73524
0 35191 7 1 2 100152 35190
0 35192 7 1 2 35189 35191
0 35193 5 1 1 35192
0 35194 7 1 2 35187 35193
0 35195 7 1 2 35148 35194
0 35196 5 1 1 35195
0 35197 7 1 2 73028 35196
0 35198 5 1 1 35197
0 35199 7 1 2 70399 430
0 35200 5 1 1 35199
0 35201 7 1 2 73813 84172
0 35202 7 2 2 35200 35201
0 35203 5 1 1 100169
0 35204 7 1 2 96310 35203
0 35205 5 2 1 35204
0 35206 7 1 2 83247 100171
0 35207 5 1 1 35206
0 35208 7 1 2 90294 99245
0 35209 5 1 1 35208
0 35210 7 1 2 35207 35209
0 35211 5 1 1 35210
0 35212 7 1 2 70736 35211
0 35213 5 1 1 35212
0 35214 7 1 2 90288 99346
0 35215 5 1 1 35214
0 35216 7 1 2 83248 94813
0 35217 5 1 1 35216
0 35218 7 1 2 73920 90241
0 35219 7 1 2 87271 35218
0 35220 5 1 1 35219
0 35221 7 1 2 35217 35220
0 35222 5 1 1 35221
0 35223 7 1 2 63981 35222
0 35224 5 1 1 35223
0 35225 7 1 2 35215 35224
0 35226 7 1 2 35213 35225
0 35227 5 1 1 35226
0 35228 7 1 2 98357 35227
0 35229 5 1 1 35228
0 35230 7 1 2 90286 98957
0 35231 5 1 1 35230
0 35232 7 1 2 90296 35231
0 35233 5 1 1 35232
0 35234 7 1 2 92173 35233
0 35235 5 1 1 35234
0 35236 7 1 2 67006 94253
0 35237 5 1 1 35236
0 35238 7 1 2 74371 5644
0 35239 5 1 1 35238
0 35240 7 1 2 65799 75808
0 35241 7 1 2 35239 35240
0 35242 5 1 1 35241
0 35243 7 1 2 35237 35242
0 35244 5 1 1 35243
0 35245 7 1 2 100130 35244
0 35246 5 1 1 35245
0 35247 7 1 2 35235 35246
0 35248 5 1 1 35247
0 35249 7 1 2 68683 35248
0 35250 5 1 1 35249
0 35251 7 2 2 82786 82852
0 35252 7 2 2 79501 93597
0 35253 5 1 1 100175
0 35254 7 1 2 85064 100176
0 35255 5 1 1 35254
0 35256 7 1 2 75905 93615
0 35257 5 1 1 35256
0 35258 7 1 2 68437 77561
0 35259 7 1 2 87956 35258
0 35260 7 1 2 35257 35259
0 35261 7 1 2 97535 35260
0 35262 5 1 1 35261
0 35263 7 1 2 35255 35262
0 35264 5 1 1 35263
0 35265 7 1 2 67007 35264
0 35266 5 1 1 35265
0 35267 7 1 2 82414 93598
0 35268 7 1 2 85455 35267
0 35269 5 1 1 35268
0 35270 7 1 2 35266 35269
0 35271 5 1 1 35270
0 35272 7 1 2 100173 35271
0 35273 5 1 1 35272
0 35274 7 2 2 69593 92218
0 35275 7 1 2 80793 100140
0 35276 7 1 2 100177 35275
0 35277 7 1 2 92238 35276
0 35278 5 1 1 35277
0 35279 7 1 2 75859 78400
0 35280 5 1 1 35279
0 35281 7 1 2 96915 35280
0 35282 5 2 1 35281
0 35283 7 1 2 69234 99089
0 35284 7 1 2 90313 35283
0 35285 7 1 2 100179 35284
0 35286 5 1 1 35285
0 35287 7 1 2 35278 35286
0 35288 5 1 1 35287
0 35289 7 1 2 71705 35288
0 35290 5 1 1 35289
0 35291 7 1 2 35273 35290
0 35292 7 1 2 35250 35291
0 35293 5 1 1 35292
0 35294 7 1 2 90611 35293
0 35295 5 1 1 35294
0 35296 7 1 2 35229 35295
0 35297 5 1 1 35296
0 35298 7 1 2 70107 35297
0 35299 5 1 1 35298
0 35300 7 1 2 85223 6764
0 35301 5 1 1 35300
0 35302 7 1 2 62158 35301
0 35303 5 1 1 35302
0 35304 7 2 2 74534 88757
0 35305 7 1 2 73716 100181
0 35306 5 1 1 35305
0 35307 7 1 2 35303 35306
0 35308 5 1 1 35307
0 35309 7 1 2 69594 82173
0 35310 7 1 2 91519 96112
0 35311 7 1 2 35309 35310
0 35312 7 1 2 35308 35311
0 35313 5 1 1 35312
0 35314 7 1 2 70108 96457
0 35315 5 1 1 35314
0 35316 7 1 2 89383 78417
0 35317 5 1 1 35316
0 35318 7 1 2 35315 35317
0 35319 5 1 1 35318
0 35320 7 1 2 82701 77685
0 35321 7 1 2 96556 35320
0 35322 7 1 2 35319 35321
0 35323 5 1 1 35322
0 35324 7 1 2 35313 35323
0 35325 5 1 1 35324
0 35326 7 1 2 62975 35325
0 35327 5 1 1 35326
0 35328 7 2 2 95918 97583
0 35329 7 3 2 70109 77091
0 35330 7 1 2 96170 100185
0 35331 7 1 2 100183 35330
0 35332 7 1 2 98958 35331
0 35333 5 1 1 35332
0 35334 7 1 2 35327 35333
0 35335 5 1 1 35334
0 35336 7 1 2 93792 35335
0 35337 5 1 1 35336
0 35338 7 1 2 35299 35337
0 35339 7 1 2 35198 35338
0 35340 7 1 2 35117 35339
0 35341 5 1 1 35340
0 35342 7 1 2 64282 35341
0 35343 5 1 1 35342
0 35344 7 4 2 82283 93793
0 35345 7 1 2 74847 100188
0 35346 7 1 2 95762 35345
0 35347 5 1 1 35346
0 35348 7 2 2 66240 82442
0 35349 5 1 1 100192
0 35350 7 1 2 99576 100193
0 35351 7 1 2 92293 35350
0 35352 5 1 1 35351
0 35353 7 1 2 35347 35352
0 35354 5 1 1 35353
0 35355 7 1 2 65466 35354
0 35356 5 1 1 35355
0 35357 7 1 2 91095 93794
0 35358 7 2 2 83718 35357
0 35359 7 1 2 82284 100194
0 35360 5 1 1 35359
0 35361 7 1 2 35356 35360
0 35362 5 1 1 35361
0 35363 7 1 2 78111 35362
0 35364 5 1 1 35363
0 35365 7 2 2 91281 100195
0 35366 7 1 2 74437 100196
0 35367 5 1 1 35366
0 35368 7 1 2 35364 35367
0 35369 5 1 1 35368
0 35370 7 1 2 67008 35369
0 35371 5 1 1 35370
0 35372 7 3 2 62159 74939
0 35373 7 1 2 100198 100197
0 35374 5 1 1 35373
0 35375 7 1 2 35371 35374
0 35376 5 1 1 35375
0 35377 7 1 2 69826 35376
0 35378 5 1 1 35377
0 35379 7 1 2 63597 98821
0 35380 5 1 1 35379
0 35381 7 1 2 95588 35380
0 35382 5 1 1 35381
0 35383 7 1 2 65800 35382
0 35384 5 1 1 35383
0 35385 7 1 2 73029 93521
0 35386 5 1 1 35385
0 35387 7 1 2 35384 35386
0 35388 5 1 1 35387
0 35389 7 1 2 62160 35388
0 35390 5 1 1 35389
0 35391 7 1 2 77305 87973
0 35392 7 1 2 94077 35391
0 35393 5 1 1 35392
0 35394 7 1 2 35390 35393
0 35395 5 1 1 35394
0 35396 7 7 2 69397 90664
0 35397 7 1 2 78554 100201
0 35398 7 1 2 35395 35397
0 35399 5 1 1 35398
0 35400 7 1 2 35378 35399
0 35401 5 1 1 35400
0 35402 7 1 2 84408 35401
0 35403 5 1 1 35402
0 35404 7 3 2 70400 94000
0 35405 7 2 2 77410 74471
0 35406 5 1 1 100211
0 35407 7 1 2 100208 100212
0 35408 5 1 1 35407
0 35409 7 1 2 76803 75715
0 35410 5 1 1 35409
0 35411 7 1 2 35408 35410
0 35412 5 1 1 35411
0 35413 7 1 2 73475 35412
0 35414 5 1 1 35413
0 35415 7 2 2 65801 88042
0 35416 5 1 1 100213
0 35417 7 1 2 35406 35416
0 35418 5 1 1 35417
0 35419 7 1 2 86175 35418
0 35420 5 1 1 35419
0 35421 7 1 2 74815 100214
0 35422 5 1 1 35421
0 35423 7 1 2 35420 35422
0 35424 5 1 1 35423
0 35425 7 1 2 70401 35424
0 35426 5 1 1 35425
0 35427 7 1 2 35414 35426
0 35428 5 1 1 35427
0 35429 7 3 2 67870 69595
0 35430 7 3 2 99018 100215
0 35431 7 1 2 79535 100218
0 35432 7 1 2 35428 35431
0 35433 5 1 1 35432
0 35434 7 1 2 35403 35433
0 35435 5 1 1 35434
0 35436 7 1 2 98979 35435
0 35437 5 1 1 35436
0 35438 7 1 2 61298 35437
0 35439 7 1 2 35343 35438
0 35440 5 1 1 35439
0 35441 7 1 2 90196 35440
0 35442 7 1 2 35086 35441
0 35443 5 1 1 35442
0 35444 7 1 2 90074 87905
0 35445 5 1 1 35444
0 35446 7 1 2 83527 97875
0 35447 5 1 1 35446
0 35448 7 1 2 35445 35447
0 35449 5 1 1 35448
0 35450 7 1 2 63025 35449
0 35451 5 1 1 35450
0 35452 7 3 2 61624 92852
0 35453 5 1 1 100221
0 35454 7 1 2 100222 98376
0 35455 5 1 1 35454
0 35456 7 1 2 35451 35455
0 35457 5 1 1 35456
0 35458 7 1 2 61377 35457
0 35459 5 1 1 35458
0 35460 7 1 2 61625 98378
0 35461 5 1 1 35460
0 35462 7 1 2 35459 35461
0 35463 5 1 1 35462
0 35464 7 1 2 94693 35463
0 35465 5 1 1 35464
0 35466 7 1 2 96576 97876
0 35467 7 1 2 98414 35466
0 35468 5 1 1 35467
0 35469 7 1 2 35465 35468
0 35470 5 1 1 35469
0 35471 7 1 2 94634 99310
0 35472 7 1 2 87769 35471
0 35473 7 1 2 35470 35472
0 35474 5 1 1 35473
0 35475 7 1 2 35443 35474
0 35476 7 1 2 34882 35475
0 35477 7 1 2 33788 35476
0 35478 7 1 2 32415 35477
0 35479 5 1 1 35478
0 35480 7 1 2 98292 35479
0 35481 5 1 1 35480
0 35482 7 1 2 71095 71456
0 35483 5 30 1 35482
0 35484 7 3 2 69398 93759
0 35485 7 1 2 86494 93716
0 35486 5 1 1 35485
0 35487 7 1 2 71253 35486
0 35488 5 1 1 35487
0 35489 7 1 2 67710 72425
0 35490 5 2 1 35489
0 35491 7 1 2 95941 100257
0 35492 5 4 1 35491
0 35493 7 3 2 66012 100259
0 35494 7 1 2 65467 100263
0 35495 5 1 1 35494
0 35496 7 1 2 35488 35495
0 35497 5 1 1 35496
0 35498 7 1 2 63598 35497
0 35499 5 1 1 35498
0 35500 7 3 2 70402 97761
0 35501 7 1 2 68438 100266
0 35502 5 1 1 35501
0 35503 7 1 2 35499 35502
0 35504 5 2 1 35503
0 35505 7 1 2 62161 100269
0 35506 5 1 1 35505
0 35507 7 1 2 75095 100267
0 35508 5 1 1 35507
0 35509 7 1 2 35506 35508
0 35510 5 1 1 35509
0 35511 7 1 2 100254 35510
0 35512 5 1 1 35511
0 35513 7 1 2 99645 100270
0 35514 5 1 1 35513
0 35515 7 2 2 81183 86155
0 35516 5 1 1 100271
0 35517 7 1 2 79626 93929
0 35518 5 1 1 35517
0 35519 7 1 2 74644 35518
0 35520 7 1 2 35516 35519
0 35521 5 1 1 35520
0 35522 7 1 2 99590 35521
0 35523 5 1 1 35522
0 35524 7 1 2 35514 35523
0 35525 5 1 1 35524
0 35526 7 1 2 62162 35525
0 35527 5 1 1 35526
0 35528 7 8 2 64543 72634
0 35529 7 1 2 63026 100273
0 35530 5 4 1 35529
0 35531 7 7 2 67871 64149
0 35532 7 1 2 100285 98646
0 35533 5 1 1 35532
0 35534 7 1 2 100281 35533
0 35535 5 1 1 35534
0 35536 7 1 2 75724 35535
0 35537 5 1 1 35536
0 35538 7 2 2 73337 78332
0 35539 5 3 1 100292
0 35540 7 1 2 99646 100293
0 35541 5 1 1 35540
0 35542 7 1 2 35537 35541
0 35543 5 1 1 35542
0 35544 7 1 2 70403 75096
0 35545 7 1 2 35543 35544
0 35546 5 1 1 35545
0 35547 7 1 2 35527 35546
0 35548 5 1 1 35547
0 35549 7 1 2 61378 35548
0 35550 5 1 1 35549
0 35551 7 1 2 35512 35550
0 35552 5 1 1 35551
0 35553 7 1 2 70110 35552
0 35554 5 1 1 35553
0 35555 7 6 2 69399 93795
0 35556 7 1 2 96227 100297
0 35557 5 1 1 35556
0 35558 7 1 2 92325 100298
0 35559 5 1 1 35558
0 35560 7 3 2 63027 88379
0 35561 5 3 1 100303
0 35562 7 1 2 61379 100304
0 35563 5 1 1 35562
0 35564 7 1 2 35559 35563
0 35565 5 1 1 35564
0 35566 7 1 2 75725 35565
0 35567 5 1 1 35566
0 35568 7 1 2 35557 35567
0 35569 5 1 1 35568
0 35570 7 1 2 77052 35569
0 35571 5 1 1 35570
0 35572 7 1 2 35554 35571
0 35573 5 1 1 35572
0 35574 7 1 2 67802 35573
0 35575 5 1 1 35574
0 35576 7 1 2 75782 77348
0 35577 5 2 1 35576
0 35578 7 1 2 77990 84116
0 35579 5 1 1 35578
0 35580 7 1 2 100309 35579
0 35581 5 1 1 35580
0 35582 7 1 2 70111 35581
0 35583 5 1 1 35582
0 35584 7 1 2 74202 96245
0 35585 5 1 1 35584
0 35586 7 1 2 35583 35585
0 35587 5 1 1 35586
0 35588 7 1 2 71341 35587
0 35589 5 1 1 35588
0 35590 7 1 2 77376 100272
0 35591 5 1 1 35590
0 35592 7 1 2 35589 35591
0 35593 5 2 1 35592
0 35594 7 2 2 98449 99751
0 35595 5 1 1 100313
0 35596 7 1 2 100311 100314
0 35597 5 1 1 35596
0 35598 7 1 2 35575 35597
0 35599 5 1 1 35598
0 35600 7 1 2 66133 35599
0 35601 5 1 1 35600
0 35602 7 3 2 67803 91371
0 35603 7 2 2 93054 100315
0 35604 5 1 1 100318
0 35605 7 1 2 100312 100319
0 35606 5 1 1 35605
0 35607 7 1 2 35601 35606
0 35608 5 1 1 35607
0 35609 7 1 2 84124 35608
0 35610 5 1 1 35609
0 35611 7 1 2 73868 93721
0 35612 5 2 1 35611
0 35613 7 1 2 67009 100320
0 35614 5 1 1 35613
0 35615 7 1 2 77349 100199
0 35616 5 1 1 35615
0 35617 7 1 2 35614 35616
0 35618 5 1 1 35617
0 35619 7 1 2 89422 93527
0 35620 7 1 2 35618 35619
0 35621 5 1 1 35620
0 35622 7 1 2 35610 35621
0 35623 5 1 1 35622
0 35624 7 1 2 64378 35623
0 35625 5 1 1 35624
0 35626 7 1 2 79038 96710
0 35627 5 1 1 35626
0 35628 7 1 2 72922 35627
0 35629 5 1 1 35628
0 35630 7 3 2 67483 83212
0 35631 7 1 2 11913 96626
0 35632 5 1 1 35631
0 35633 7 1 2 100322 35632
0 35634 5 1 1 35633
0 35635 7 1 2 35629 35634
0 35636 5 1 1 35635
0 35637 7 1 2 80488 99006
0 35638 7 1 2 35636 35637
0 35639 5 1 1 35638
0 35640 7 1 2 72560 86470
0 35641 5 1 1 35640
0 35642 7 1 2 95976 95942
0 35643 5 1 1 35642
0 35644 7 1 2 65468 35643
0 35645 5 1 1 35644
0 35646 7 1 2 35641 35645
0 35647 5 1 1 35646
0 35648 7 1 2 67484 35647
0 35649 5 1 1 35648
0 35650 7 1 2 76262 35649
0 35651 5 1 1 35650
0 35652 7 1 2 92535 99352
0 35653 7 1 2 35651 35652
0 35654 5 1 1 35653
0 35655 7 1 2 35639 35654
0 35656 5 1 1 35655
0 35657 7 1 2 62163 35656
0 35658 5 1 1 35657
0 35659 7 1 2 77922 84291
0 35660 5 1 1 35659
0 35661 7 1 2 73263 92416
0 35662 5 1 1 35661
0 35663 7 1 2 35660 35662
0 35664 5 1 1 35663
0 35665 7 1 2 68439 35664
0 35666 5 1 1 35665
0 35667 7 2 2 68865 78418
0 35668 7 1 2 74405 100325
0 35669 5 1 1 35668
0 35670 7 1 2 35666 35669
0 35671 5 2 1 35670
0 35672 7 1 2 77500 100327
0 35673 5 1 1 35672
0 35674 7 1 2 72304 95772
0 35675 5 2 1 35674
0 35676 7 1 2 65469 100329
0 35677 5 1 1 35676
0 35678 7 1 2 86410 72461
0 35679 5 1 1 35678
0 35680 7 1 2 35677 35679
0 35681 5 1 1 35680
0 35682 7 1 2 67485 35681
0 35683 5 1 1 35682
0 35684 7 1 2 76263 35683
0 35685 5 2 1 35684
0 35686 7 1 2 94943 100331
0 35687 5 1 1 35686
0 35688 7 1 2 35673 35687
0 35689 5 1 1 35688
0 35690 7 5 2 67010 63028
0 35691 7 1 2 83384 100333
0 35692 7 1 2 35689 35691
0 35693 5 1 1 35692
0 35694 7 1 2 35658 35693
0 35695 5 1 1 35694
0 35696 7 1 2 66241 35695
0 35697 5 1 1 35696
0 35698 7 1 2 67011 100328
0 35699 5 1 1 35698
0 35700 7 2 2 62164 77474
0 35701 5 1 1 100338
0 35702 7 1 2 100326 100339
0 35703 5 1 1 35702
0 35704 7 1 2 35699 35703
0 35705 5 1 1 35704
0 35706 7 1 2 77501 35705
0 35707 5 1 1 35706
0 35708 7 1 2 95342 100332
0 35709 5 1 1 35708
0 35710 7 1 2 35707 35709
0 35711 5 1 1 35710
0 35712 7 1 2 83385 93745
0 35713 7 1 2 35711 35712
0 35714 5 1 1 35713
0 35715 7 1 2 35697 35714
0 35716 5 1 1 35715
0 35717 7 1 2 64544 35716
0 35718 5 1 1 35717
0 35719 7 2 2 84146 90665
0 35720 7 1 2 264 98289
0 35721 5 1 1 35720
0 35722 7 1 2 65470 86741
0 35723 7 1 2 35721 35722
0 35724 5 1 1 35723
0 35725 7 1 2 79584 35724
0 35726 5 1 1 35725
0 35727 7 1 2 71538 35726
0 35728 5 1 1 35727
0 35729 7 2 2 72250 75013
0 35730 5 1 1 100342
0 35731 7 1 2 73076 100343
0 35732 5 1 1 35731
0 35733 7 1 2 35728 35732
0 35734 5 1 1 35733
0 35735 7 1 2 88818 35734
0 35736 5 1 1 35735
0 35737 7 3 2 70112 73128
0 35738 7 2 2 66013 100344
0 35739 7 1 2 74332 90440
0 35740 7 1 2 100347 35739
0 35741 5 1 1 35740
0 35742 7 1 2 35736 35741
0 35743 5 1 1 35742
0 35744 7 1 2 100340 35743
0 35745 5 1 1 35744
0 35746 7 1 2 35718 35745
0 35747 5 1 1 35746
0 35748 7 1 2 93512 35747
0 35749 5 1 1 35748
0 35750 7 2 2 70939 74139
0 35751 5 1 1 100349
0 35752 7 1 2 88819 96520
0 35753 7 1 2 100350 35752
0 35754 5 1 1 35753
0 35755 7 1 2 73653 96531
0 35756 7 1 2 89390 35755
0 35757 5 1 1 35756
0 35758 7 1 2 35754 35757
0 35759 5 1 1 35758
0 35760 7 1 2 93796 35759
0 35761 5 1 1 35760
0 35762 7 1 2 88031 99062
0 35763 7 1 2 99988 35762
0 35764 7 1 2 84147 35763
0 35765 7 1 2 95558 35764
0 35766 5 1 1 35765
0 35767 7 1 2 35761 35766
0 35768 5 1 1 35767
0 35769 7 1 2 65802 35768
0 35770 5 1 1 35769
0 35771 7 1 2 69015 75542
0 35772 5 3 1 35771
0 35773 7 2 2 84770 100351
0 35774 5 5 1 100354
0 35775 7 8 2 61380 64379
0 35776 7 1 2 100361 99353
0 35777 7 1 2 100064 35776
0 35778 7 1 2 88820 35777
0 35779 7 1 2 100356 35778
0 35780 5 1 1 35779
0 35781 7 1 2 35770 35780
0 35782 5 1 1 35781
0 35783 7 1 2 92642 35782
0 35784 5 1 1 35783
0 35785 7 1 2 76252 75543
0 35786 5 1 1 35785
0 35787 7 1 2 69016 83192
0 35788 5 1 1 35787
0 35789 7 1 2 66014 77956
0 35790 7 1 2 35788 35789
0 35791 5 1 1 35790
0 35792 7 1 2 35786 35791
0 35793 5 1 1 35792
0 35794 7 1 2 88821 35793
0 35795 5 1 1 35794
0 35796 7 1 2 74082 74333
0 35797 7 1 2 79323 35796
0 35798 5 1 1 35797
0 35799 7 1 2 35795 35798
0 35800 5 1 1 35799
0 35801 7 1 2 99418 100341
0 35802 7 1 2 35800 35801
0 35803 5 1 1 35802
0 35804 7 1 2 35784 35803
0 35805 5 1 1 35804
0 35806 7 1 2 73476 35805
0 35807 5 1 1 35806
0 35808 7 1 2 69126 35807
0 35809 7 1 2 35749 35808
0 35810 7 1 2 35625 35809
0 35811 5 1 1 35810
0 35812 7 2 2 81061 88832
0 35813 7 1 2 92322 95890
0 35814 7 1 2 93247 35813
0 35815 7 1 2 100369 35814
0 35816 5 1 1 35815
0 35817 7 1 2 74372 94516
0 35818 5 1 1 35817
0 35819 7 1 2 12598 35818
0 35820 5 1 1 35819
0 35821 7 2 2 69596 77130
0 35822 7 1 2 81699 100371
0 35823 7 1 2 35820 35822
0 35824 5 1 1 35823
0 35825 7 1 2 35816 35824
0 35826 5 1 1 35825
0 35827 7 1 2 93599 35826
0 35828 5 1 1 35827
0 35829 7 1 2 86871 96679
0 35830 7 1 2 76419 35829
0 35831 7 1 2 95162 97350
0 35832 7 1 2 35830 35831
0 35833 5 1 1 35832
0 35834 7 1 2 35828 35833
0 35835 5 1 1 35834
0 35836 7 1 2 90612 35835
0 35837 5 1 1 35836
0 35838 7 1 2 78043 72751
0 35839 7 1 2 91391 80260
0 35840 7 2 2 35838 35839
0 35841 7 3 2 66242 98450
0 35842 5 1 1 100375
0 35843 7 2 2 72706 81592
0 35844 7 1 2 100376 100378
0 35845 7 1 2 100373 35844
0 35846 5 1 1 35845
0 35847 7 1 2 35837 35846
0 35848 5 1 1 35847
0 35849 7 1 2 61299 35848
0 35850 5 1 1 35849
0 35851 7 1 2 91010 100379
0 35852 7 1 2 100374 35851
0 35853 5 1 1 35852
0 35854 7 1 2 35850 35853
0 35855 5 1 1 35854
0 35856 7 1 2 65471 35855
0 35857 5 1 1 35856
0 35858 7 1 2 68206 91799
0 35859 7 1 2 77120 35858
0 35860 7 1 2 84272 35859
0 35861 5 1 1 35860
0 35862 7 2 2 74203 82812
0 35863 7 1 2 84456 98619
0 35864 7 1 2 100380 35863
0 35865 5 1 1 35864
0 35866 7 1 2 35861 35865
0 35867 5 1 1 35866
0 35868 7 1 2 61300 35867
0 35869 5 1 1 35868
0 35870 7 3 2 62976 81711
0 35871 7 1 2 84457 100382
0 35872 7 1 2 100381 35871
0 35873 5 1 1 35872
0 35874 7 1 2 35869 35873
0 35875 5 1 1 35874
0 35876 7 1 2 93703 35875
0 35877 5 1 1 35876
0 35878 7 2 2 62977 79502
0 35879 7 2 2 69017 82993
0 35880 7 1 2 61301 91330
0 35881 7 1 2 95045 35880
0 35882 7 1 2 100387 35881
0 35883 7 1 2 100385 35882
0 35884 5 1 1 35883
0 35885 7 2 2 71739 78300
0 35886 5 1 1 100389
0 35887 7 1 2 84698 35886
0 35888 5 1 1 35887
0 35889 7 1 2 62165 35888
0 35890 5 1 1 35889
0 35891 7 1 2 86853 92610
0 35892 5 1 1 35891
0 35893 7 1 2 35890 35892
0 35894 5 1 1 35893
0 35895 7 1 2 93859 96536
0 35896 7 1 2 35894 35895
0 35897 5 1 1 35896
0 35898 7 1 2 35884 35897
0 35899 5 1 1 35898
0 35900 7 1 2 69235 35899
0 35901 5 1 1 35900
0 35902 7 2 2 75544 75726
0 35903 5 1 1 100391
0 35904 7 1 2 99870 100392
0 35905 5 1 1 35904
0 35906 7 4 2 70940 73264
0 35907 7 2 2 77983 100393
0 35908 5 1 1 100397
0 35909 7 1 2 74708 100398
0 35910 5 1 1 35909
0 35911 7 1 2 35905 35910
0 35912 5 1 1 35911
0 35913 7 1 2 64150 35912
0 35914 5 1 1 35913
0 35915 7 2 2 73077 94423
0 35916 5 1 1 100399
0 35917 7 1 2 74373 100400
0 35918 5 1 1 35917
0 35919 7 1 2 35914 35918
0 35920 5 1 1 35919
0 35921 7 1 2 96532 96942
0 35922 7 1 2 35920 35921
0 35923 5 1 1 35922
0 35924 7 1 2 35901 35923
0 35925 5 1 1 35924
0 35926 7 1 2 70113 35925
0 35927 5 1 1 35926
0 35928 7 1 2 35877 35927
0 35929 5 1 1 35928
0 35930 7 1 2 93797 35929
0 35931 5 1 1 35930
0 35932 7 1 2 64283 35931
0 35933 7 1 2 35857 35932
0 35934 5 1 1 35933
0 35935 7 1 2 76173 35934
0 35936 7 1 2 35811 35935
0 35937 5 1 1 35936
0 35938 7 2 2 63186 80261
0 35939 5 1 1 100401
0 35940 7 1 2 81402 78771
0 35941 5 1 1 35940
0 35942 7 1 2 35939 35941
0 35943 5 1 1 35942
0 35944 7 1 2 75163 35943
0 35945 5 1 1 35944
0 35946 7 1 2 78932 75112
0 35947 7 1 2 94952 35946
0 35948 5 1 1 35947
0 35949 7 1 2 35945 35948
0 35950 5 1 1 35949
0 35951 7 1 2 94725 35950
0 35952 5 1 1 35951
0 35953 7 1 2 63599 95520
0 35954 5 1 1 35953
0 35955 7 1 2 96283 35954
0 35956 5 1 1 35955
0 35957 7 13 2 62871 98293
0 35958 5 7 1 100403
0 35959 7 1 2 68440 100404
0 35960 5 1 1 35959
0 35961 7 1 2 85633 35960
0 35962 5 2 1 35961
0 35963 7 1 2 75809 87951
0 35964 7 1 2 100423 35963
0 35965 5 1 1 35964
0 35966 7 1 2 35956 35965
0 35967 5 1 1 35966
0 35968 7 3 2 69597 77247
0 35969 7 1 2 94612 100425
0 35970 7 1 2 35967 35969
0 35971 5 1 1 35970
0 35972 7 1 2 35952 35971
0 35973 5 1 1 35972
0 35974 7 1 2 65472 35973
0 35975 5 1 1 35974
0 35976 7 1 2 71342 95259
0 35977 5 1 1 35976
0 35978 7 1 2 64151 94710
0 35979 5 1 1 35978
0 35980 7 1 2 35977 35979
0 35981 5 1 1 35980
0 35982 7 1 2 77320 35981
0 35983 5 1 1 35982
0 35984 7 1 2 71539 73147
0 35985 7 1 2 94711 35984
0 35986 5 1 1 35985
0 35987 7 1 2 35983 35986
0 35988 5 1 1 35987
0 35989 7 1 2 70941 35988
0 35990 5 1 1 35989
0 35991 7 2 2 94680 94829
0 35992 7 1 2 83750 97263
0 35993 7 1 2 100428 35992
0 35994 5 1 1 35993
0 35995 7 1 2 35990 35994
0 35996 5 1 1 35995
0 35997 7 1 2 68441 35996
0 35998 5 1 1 35997
0 35999 7 1 2 88349 80608
0 36000 7 1 2 93911 35999
0 36001 7 1 2 89243 92256
0 36002 7 1 2 36000 36001
0 36003 5 1 1 36002
0 36004 7 1 2 35998 36003
0 36005 5 1 1 36004
0 36006 7 1 2 79543 36005
0 36007 5 1 1 36006
0 36008 7 1 2 35975 36007
0 36009 5 1 1 36008
0 36010 7 1 2 89109 36009
0 36011 5 1 1 36010
0 36012 7 1 2 88445 79524
0 36013 7 1 2 82315 95564
0 36014 7 1 2 36012 36013
0 36015 5 1 1 36014
0 36016 7 1 2 36011 36015
0 36017 5 1 1 36016
0 36018 7 1 2 93860 36017
0 36019 5 1 1 36018
0 36020 7 4 2 72277 72707
0 36021 5 2 1 100430
0 36022 7 1 2 96363 100434
0 36023 5 1 1 36022
0 36024 7 1 2 96393 36023
0 36025 5 1 1 36024
0 36026 7 1 2 62872 76327
0 36027 5 4 1 36026
0 36028 7 1 2 7281 100436
0 36029 5 1 1 36028
0 36030 7 1 2 96590 36029
0 36031 5 1 1 36030
0 36032 7 1 2 36025 36031
0 36033 5 1 1 36032
0 36034 7 1 2 86061 36033
0 36035 5 1 1 36034
0 36036 7 1 2 85762 84570
0 36037 5 1 1 36036
0 36038 7 1 2 70737 36037
0 36039 5 1 1 36038
0 36040 7 1 2 92410 36039
0 36041 5 1 1 36040
0 36042 7 2 2 61626 90961
0 36043 7 2 2 70404 85727
0 36044 7 1 2 100440 100442
0 36045 7 1 2 36041 36044
0 36046 5 1 1 36045
0 36047 7 1 2 36035 36046
0 36048 5 1 1 36047
0 36049 7 1 2 69598 36048
0 36050 5 1 1 36049
0 36051 7 1 2 78793 84292
0 36052 5 1 1 36051
0 36053 7 1 2 99943 36052
0 36054 5 1 1 36053
0 36055 7 1 2 80815 93046
0 36056 7 1 2 36054 36055
0 36057 5 1 1 36056
0 36058 7 1 2 36050 36057
0 36059 5 1 1 36058
0 36060 7 1 2 64152 36059
0 36061 5 1 1 36060
0 36062 7 2 2 63982 81932
0 36063 5 1 1 100444
0 36064 7 1 2 78794 86437
0 36065 5 1 1 36064
0 36066 7 3 2 74626 73739
0 36067 5 1 1 100446
0 36068 7 1 2 67486 100447
0 36069 5 1 1 36068
0 36070 7 1 2 36065 36069
0 36071 5 1 1 36070
0 36072 7 1 2 100445 36071
0 36073 5 1 1 36072
0 36074 7 1 2 74627 94051
0 36075 7 1 2 95683 36074
0 36076 5 1 1 36075
0 36077 7 1 2 36073 36076
0 36078 5 1 1 36077
0 36079 7 1 2 68028 36078
0 36080 5 1 1 36079
0 36081 7 2 2 66520 92090
0 36082 5 1 1 100449
0 36083 7 1 2 88100 78795
0 36084 7 1 2 100450 36083
0 36085 5 1 1 36084
0 36086 7 1 2 36080 36085
0 36087 5 1 1 36086
0 36088 7 1 2 92801 36087
0 36089 5 1 1 36088
0 36090 7 1 2 74472 77350
0 36091 5 2 1 36090
0 36092 7 1 2 72853 94424
0 36093 5 1 1 36092
0 36094 7 1 2 100451 36093
0 36095 5 1 1 36094
0 36096 7 1 2 96674 36095
0 36097 5 1 1 36096
0 36098 7 1 2 36089 36097
0 36099 5 1 1 36098
0 36100 7 1 2 70738 36099
0 36101 5 1 1 36100
0 36102 7 2 2 1431 94497
0 36103 5 2 1 100453
0 36104 7 3 2 80731 96620
0 36105 7 1 2 100455 100457
0 36106 5 2 1 36105
0 36107 7 1 2 71128 77248
0 36108 7 1 2 96857 36107
0 36109 5 1 1 36108
0 36110 7 1 2 100460 36109
0 36111 5 1 1 36110
0 36112 7 1 2 90773 93934
0 36113 7 1 2 36111 36112
0 36114 5 1 1 36113
0 36115 7 1 2 36101 36114
0 36116 7 1 2 36061 36115
0 36117 5 1 1 36116
0 36118 7 1 2 68442 36117
0 36119 5 1 1 36118
0 36120 7 1 2 89067 96135
0 36121 5 1 1 36120
0 36122 7 1 2 61627 96824
0 36123 5 1 1 36122
0 36124 7 1 2 36121 36123
0 36125 5 1 1 36124
0 36126 7 1 2 90122 95054
0 36127 7 1 2 36125 36126
0 36128 5 1 1 36127
0 36129 7 1 2 36119 36128
0 36130 5 1 1 36129
0 36131 7 1 2 97307 36130
0 36132 5 1 1 36131
0 36133 7 1 2 73218 85282
0 36134 5 1 1 36133
0 36135 7 1 2 68443 36134
0 36136 5 1 1 36135
0 36137 7 1 2 97515 36136
0 36138 5 1 1 36137
0 36139 7 1 2 75119 36138
0 36140 5 1 1 36139
0 36141 7 1 2 65473 36140
0 36142 5 1 1 36141
0 36143 7 2 2 72757 95485
0 36144 7 1 2 78658 100462
0 36145 5 1 1 36144
0 36146 7 1 2 36142 36145
0 36147 5 1 1 36146
0 36148 7 1 2 96394 36147
0 36149 5 1 1 36148
0 36150 7 1 2 1709 93722
0 36151 5 1 1 36150
0 36152 7 1 2 73477 36151
0 36153 5 1 1 36152
0 36154 7 1 2 75880 73865
0 36155 5 1 1 36154
0 36156 7 1 2 36153 36155
0 36157 5 1 1 36156
0 36158 7 1 2 65803 36157
0 36159 5 1 1 36158
0 36160 7 1 2 89528 73866
0 36161 5 1 1 36160
0 36162 7 1 2 36159 36161
0 36163 5 1 1 36162
0 36164 7 1 2 96591 36163
0 36165 5 1 1 36164
0 36166 7 1 2 36149 36165
0 36167 5 1 1 36166
0 36168 7 1 2 94732 96943
0 36169 7 1 2 36167 36168
0 36170 5 1 1 36169
0 36171 7 1 2 36132 36170
0 36172 5 1 1 36171
0 36173 7 1 2 68207 36172
0 36174 5 1 1 36173
0 36175 7 1 2 5715 100458
0 36176 5 1 1 36175
0 36177 7 1 2 92433 96592
0 36178 5 1 1 36177
0 36179 7 1 2 36176 36178
0 36180 5 1 1 36179
0 36181 7 1 2 62873 36180
0 36182 5 1 1 36181
0 36183 7 1 2 93553 100459
0 36184 5 1 1 36183
0 36185 7 1 2 36182 36184
0 36186 5 1 1 36185
0 36187 7 3 2 67804 81712
0 36188 7 2 2 63375 100464
0 36189 7 1 2 88101 99165
0 36190 7 1 2 100467 36189
0 36191 7 1 2 36186 36190
0 36192 5 1 1 36191
0 36193 7 1 2 65181 36192
0 36194 7 1 2 36174 36193
0 36195 5 1 1 36194
0 36196 7 1 2 64153 76740
0 36197 5 1 1 36196
0 36198 7 1 2 85953 36197
0 36199 5 1 1 36198
0 36200 7 3 2 78890 98520
0 36201 7 1 2 36199 100469
0 36202 5 1 1 36201
0 36203 7 3 2 74126 75727
0 36204 5 1 1 100472
0 36205 7 1 2 78933 99914
0 36206 7 1 2 100473 36205
0 36207 5 1 1 36206
0 36208 7 1 2 36202 36207
0 36209 5 1 1 36208
0 36210 7 1 2 70942 36209
0 36211 5 1 1 36210
0 36212 7 1 2 100264 100470
0 36213 5 1 1 36212
0 36214 7 1 2 36211 36213
0 36215 5 1 1 36214
0 36216 7 1 2 63600 36215
0 36217 5 1 1 36216
0 36218 7 4 2 65804 100405
0 36219 5 1 1 100475
0 36220 7 1 2 100476 100471
0 36221 5 1 1 36220
0 36222 7 3 2 67805 64154
0 36223 7 1 2 94759 100479
0 36224 7 1 2 98833 36223
0 36225 7 1 2 80252 36224
0 36226 5 1 1 36225
0 36227 7 1 2 36221 36226
0 36228 5 1 1 36227
0 36229 7 1 2 62166 36228
0 36230 5 1 1 36229
0 36231 7 1 2 36217 36230
0 36232 5 1 1 36231
0 36233 7 1 2 63376 36232
0 36234 5 1 1 36233
0 36235 7 1 2 91191 93327
0 36236 7 1 2 95887 99915
0 36237 7 1 2 36235 36236
0 36238 5 1 1 36237
0 36239 7 1 2 36234 36238
0 36240 5 1 1 36239
0 36241 7 1 2 70405 36240
0 36242 5 1 1 36241
0 36243 7 2 2 95151 96944
0 36244 7 1 2 92882 100482
0 36245 5 1 1 36244
0 36246 7 2 2 62874 85453
0 36247 5 2 1 100484
0 36248 7 2 2 87957 100486
0 36249 5 1 1 100488
0 36250 7 1 2 88868 97308
0 36251 7 1 2 100489 36250
0 36252 5 1 1 36251
0 36253 7 1 2 36245 36252
0 36254 5 1 1 36253
0 36255 7 1 2 64155 36254
0 36256 5 1 1 36255
0 36257 7 1 2 91665 100483
0 36258 5 1 1 36257
0 36259 7 2 2 66134 69018
0 36260 7 4 2 97984 100490
0 36261 7 1 2 77172 91192
0 36262 7 1 2 100492 36261
0 36263 5 1 1 36262
0 36264 7 1 2 36258 36263
0 36265 5 1 1 36264
0 36266 7 1 2 62875 36265
0 36267 5 1 1 36266
0 36268 7 1 2 36256 36267
0 36269 5 1 1 36268
0 36270 7 1 2 70943 36269
0 36271 5 1 1 36270
0 36272 7 4 2 64284 70739
0 36273 7 2 2 96945 100496
0 36274 5 3 1 100500
0 36275 7 1 2 78891 100501
0 36276 7 1 2 92330 36275
0 36277 5 1 1 36276
0 36278 7 1 2 36271 36277
0 36279 5 1 1 36278
0 36280 7 1 2 98228 36279
0 36281 5 1 1 36280
0 36282 7 1 2 36242 36281
0 36283 5 1 1 36282
0 36284 7 1 2 61628 93120
0 36285 7 1 2 36283 36284
0 36286 5 1 1 36285
0 36287 7 5 2 96946 99121
0 36288 5 2 1 100505
0 36289 7 1 2 96647 100506
0 36290 5 1 1 36289
0 36291 7 5 2 98037 100465
0 36292 5 1 1 100512
0 36293 7 1 2 74127 85545
0 36294 7 1 2 100513 36293
0 36295 5 1 1 36294
0 36296 7 1 2 36290 36295
0 36297 5 1 1 36296
0 36298 7 1 2 70944 36297
0 36299 5 1 1 36298
0 36300 7 1 2 67487 100330
0 36301 5 1 1 36300
0 36302 7 1 2 81224 36301
0 36303 5 1 1 36302
0 36304 7 1 2 100514 36303
0 36305 5 1 1 36304
0 36306 7 1 2 36299 36305
0 36307 5 1 1 36306
0 36308 7 1 2 63601 36307
0 36309 5 1 1 36308
0 36310 7 1 2 93947 98521
0 36311 7 1 2 96215 36310
0 36312 5 1 1 36311
0 36313 7 1 2 36309 36312
0 36314 5 1 1 36313
0 36315 7 1 2 82549 96395
0 36316 7 1 2 36314 36315
0 36317 5 1 1 36316
0 36318 7 1 2 70114 36317
0 36319 7 1 2 36286 36318
0 36320 5 1 1 36319
0 36321 7 1 2 36195 36320
0 36322 5 1 1 36321
0 36323 7 1 2 36019 36322
0 36324 5 1 1 36323
0 36325 7 1 2 93798 36324
0 36326 5 1 1 36325
0 36327 7 5 2 62876 99647
0 36328 5 1 1 100517
0 36329 7 1 2 66015 100518
0 36330 5 1 1 36329
0 36331 7 1 2 99607 36330
0 36332 5 1 1 36331
0 36333 7 1 2 81933 36332
0 36334 5 1 1 36333
0 36335 7 1 2 93407 99648
0 36336 5 1 1 36335
0 36337 7 1 2 36334 36336
0 36338 5 1 1 36337
0 36339 7 1 2 62608 36338
0 36340 5 1 1 36339
0 36341 7 1 2 81877 99577
0 36342 5 2 1 36341
0 36343 7 1 2 100522 99608
0 36344 5 3 1 36343
0 36345 7 1 2 90569 100524
0 36346 5 1 1 36345
0 36347 7 1 2 36340 36346
0 36348 5 1 1 36347
0 36349 7 1 2 64156 36348
0 36350 5 1 1 36349
0 36351 7 2 2 62877 99591
0 36352 5 2 1 100527
0 36353 7 1 2 79492 99649
0 36354 5 2 1 36353
0 36355 7 1 2 100529 100531
0 36356 5 1 1 36355
0 36357 7 1 2 90570 36356
0 36358 5 1 1 36357
0 36359 7 1 2 36350 36358
0 36360 5 1 1 36359
0 36361 7 1 2 88725 36360
0 36362 5 1 1 36361
0 36363 7 2 2 67872 84534
0 36364 5 1 1 100533
0 36365 7 1 2 80189 80732
0 36366 5 1 1 36365
0 36367 7 1 2 74128 90571
0 36368 5 1 1 36367
0 36369 7 1 2 36366 36368
0 36370 5 1 1 36369
0 36371 7 2 2 64545 36370
0 36372 7 1 2 100534 100535
0 36373 5 1 1 36372
0 36374 7 1 2 36362 36373
0 36375 5 1 1 36374
0 36376 7 1 2 66243 36375
0 36377 5 1 1 36376
0 36378 7 4 2 89120 15949
0 36379 7 2 2 64157 100537
0 36380 7 1 2 99650 100541
0 36381 5 1 1 36380
0 36382 7 1 2 70945 100528
0 36383 5 1 1 36382
0 36384 7 1 2 36381 36383
0 36385 5 1 1 36384
0 36386 7 1 2 66244 36385
0 36387 5 1 1 36386
0 36388 7 1 2 84514 93746
0 36389 5 2 1 36388
0 36390 7 1 2 63029 84515
0 36391 5 2 1 36390
0 36392 7 1 2 100545 100532
0 36393 5 1 1 36392
0 36394 7 1 2 66245 36393
0 36395 5 1 1 36394
0 36396 7 1 2 100543 36395
0 36397 5 1 1 36396
0 36398 7 1 2 75545 36397
0 36399 5 1 1 36398
0 36400 7 9 2 64546 93747
0 36401 5 1 1 100547
0 36402 7 1 2 73557 100548
0 36403 5 1 1 36402
0 36404 7 1 2 36399 36403
0 36405 7 1 2 36387 36404
0 36406 5 1 1 36405
0 36407 7 1 2 84409 36406
0 36408 5 1 1 36407
0 36409 7 1 2 84320 83371
0 36410 5 4 1 36409
0 36411 7 4 2 66246 100216
0 36412 7 1 2 82853 100560
0 36413 7 1 2 100556 36412
0 36414 5 1 1 36413
0 36415 7 1 2 36408 36414
0 36416 5 1 1 36415
0 36417 7 1 2 94914 36416
0 36418 5 1 1 36417
0 36419 7 2 2 67873 98201
0 36420 7 2 2 91824 100564
0 36421 5 1 1 100566
0 36422 7 1 2 100567 100536
0 36423 5 1 1 36422
0 36424 7 1 2 36418 36423
0 36425 7 1 2 36377 36424
0 36426 5 1 1 36425
0 36427 7 1 2 69236 36426
0 36428 5 1 1 36427
0 36429 7 2 2 70946 98770
0 36430 7 1 2 91520 96882
0 36431 7 1 2 94915 36430
0 36432 7 1 2 100568 36431
0 36433 5 1 1 36432
0 36434 7 1 2 36428 36433
0 36435 5 1 1 36434
0 36436 7 1 2 97985 36435
0 36437 5 1 1 36436
0 36438 7 1 2 61629 98776
0 36439 5 1 1 36438
0 36440 7 1 2 78956 99113
0 36441 5 1 1 36440
0 36442 7 1 2 36439 36441
0 36443 5 1 1 36442
0 36444 7 1 2 81328 94635
0 36445 7 1 2 95371 97528
0 36446 7 1 2 36444 36445
0 36447 7 1 2 95046 36446
0 36448 7 1 2 36443 36447
0 36449 5 1 1 36448
0 36450 7 1 2 36437 36449
0 36451 5 1 1 36450
0 36452 7 1 2 66135 36451
0 36453 5 1 1 36452
0 36454 7 11 2 89264 93799
0 36455 7 4 2 67806 63187
0 36456 7 1 2 100570 100581
0 36457 5 1 1 36456
0 36458 7 1 2 90715 91977
0 36459 5 1 1 36458
0 36460 7 1 2 36457 36459
0 36461 5 1 1 36460
0 36462 7 1 2 81329 75810
0 36463 7 1 2 91392 84279
0 36464 7 1 2 36462 36463
0 36465 7 1 2 98223 36464
0 36466 7 1 2 36461 36465
0 36467 5 1 1 36466
0 36468 7 1 2 36453 36467
0 36469 5 1 1 36468
0 36470 7 1 2 79052 36469
0 36471 5 1 1 36470
0 36472 7 1 2 14211 17063
0 36473 5 2 1 36472
0 36474 7 1 2 16425 32974
0 36475 7 10 2 100585 36474
0 36476 7 1 2 66136 100587
0 36477 5 1 1 36476
0 36478 7 4 2 66521 98473
0 36479 7 1 2 92960 100597
0 36480 5 1 1 36479
0 36481 7 1 2 36477 36480
0 36482 5 5 1 36481
0 36483 7 1 2 86839 96103
0 36484 7 1 2 100601 36483
0 36485 5 1 1 36484
0 36486 7 3 2 63030 83817
0 36487 7 1 2 84410 100606
0 36488 7 1 2 99427 97351
0 36489 7 1 2 36487 36488
0 36490 5 1 1 36489
0 36491 7 1 2 36485 36490
0 36492 5 1 1 36491
0 36493 7 1 2 78112 36492
0 36494 5 1 1 36493
0 36495 7 1 2 80660 83305
0 36496 7 3 2 91804 93695
0 36497 7 1 2 96080 100609
0 36498 7 1 2 36495 36497
0 36499 5 1 1 36498
0 36500 7 1 2 36494 36499
0 36501 5 1 1 36500
0 36502 7 1 2 66247 36501
0 36503 5 1 1 36502
0 36504 7 2 2 66137 98170
0 36505 7 1 2 67807 80941
0 36506 7 2 2 100612 36505
0 36507 7 2 2 64769 91699
0 36508 7 1 2 92853 96764
0 36509 7 1 2 100616 36508
0 36510 7 1 2 100614 36509
0 36511 5 1 1 36510
0 36512 7 1 2 36503 36511
0 36513 5 1 1 36512
0 36514 7 1 2 65474 36513
0 36515 5 1 1 36514
0 36516 7 1 2 68029 71540
0 36517 7 1 2 100132 36516
0 36518 7 1 2 91700 91754
0 36519 7 1 2 36517 36518
0 36520 7 1 2 100615 36519
0 36521 5 1 1 36520
0 36522 7 1 2 36515 36521
0 36523 5 1 1 36522
0 36524 7 1 2 67012 36523
0 36525 5 1 1 36524
0 36526 7 1 2 99462 98368
0 36527 5 1 1 36526
0 36528 7 11 2 61381 68030
0 36529 5 1 1 100618
0 36530 7 1 2 100619 99634
0 36531 7 1 2 96989 36530
0 36532 5 1 1 36531
0 36533 7 1 2 36527 36532
0 36534 5 1 1 36533
0 36535 7 4 2 66138 79260
0 36536 7 9 2 69237 65182
0 36537 7 1 2 100633 100069
0 36538 7 1 2 100629 36537
0 36539 7 1 2 97352 36538
0 36540 7 1 2 36534 36539
0 36541 5 1 1 36540
0 36542 7 1 2 36525 36541
0 36543 5 1 1 36542
0 36544 7 1 2 68208 36543
0 36545 5 1 1 36544
0 36546 7 2 2 81372 93121
0 36547 7 1 2 66248 100642
0 36548 7 1 2 88822 36547
0 36549 7 1 2 100602 36548
0 36550 5 1 1 36549
0 36551 7 1 2 74225 82095
0 36552 7 1 2 97400 36551
0 36553 7 2 2 92802 93001
0 36554 5 1 1 100644
0 36555 7 1 2 82556 100645
0 36556 7 1 2 36552 36555
0 36557 5 1 1 36556
0 36558 7 1 2 36550 36557
0 36559 5 1 1 36558
0 36560 7 1 2 93494 36559
0 36561 5 1 1 36560
0 36562 7 1 2 64547 90812
0 36563 7 3 2 79261 92834
0 36564 7 1 2 100610 100646
0 36565 7 1 2 98932 36564
0 36566 7 1 2 36562 36565
0 36567 5 1 1 36566
0 36568 7 1 2 69127 36567
0 36569 7 1 2 36561 36568
0 36570 7 1 2 36545 36569
0 36571 5 1 1 36570
0 36572 7 1 2 61302 100588
0 36573 5 1 1 36572
0 36574 7 1 2 87684 98115
0 36575 5 1 1 36574
0 36576 7 1 2 36573 36575
0 36577 5 1 1 36576
0 36578 7 2 2 69238 36577
0 36579 7 1 2 62167 82568
0 36580 5 1 1 36579
0 36581 7 1 2 89915 91553
0 36582 5 1 1 36581
0 36583 7 1 2 36580 36582
0 36584 5 1 1 36583
0 36585 7 1 2 99997 36584
0 36586 5 1 1 36585
0 36587 7 2 2 69599 79298
0 36588 7 2 2 81538 98171
0 36589 7 1 2 93463 100653
0 36590 7 1 2 100651 36589
0 36591 5 1 1 36590
0 36592 7 1 2 36586 36591
0 36593 5 1 1 36592
0 36594 7 1 2 100649 36593
0 36595 5 1 1 36594
0 36596 7 1 2 80774 92572
0 36597 7 1 2 97421 99764
0 36598 7 1 2 36596 36597
0 36599 7 2 2 61303 99019
0 36600 7 2 2 81773 98699
0 36601 7 1 2 100655 100657
0 36602 7 1 2 36598 36601
0 36603 5 1 1 36602
0 36604 7 1 2 36595 36603
0 36605 5 1 1 36604
0 36606 7 1 2 65475 36605
0 36607 5 1 1 36606
0 36608 7 1 2 82550 96463
0 36609 5 1 1 36608
0 36610 7 1 2 68209 86652
0 36611 7 1 2 100652 36610
0 36612 5 1 1 36611
0 36613 7 1 2 36609 36612
0 36614 5 1 1 36613
0 36615 7 2 2 70406 93122
0 36616 7 6 2 98104 99225
0 36617 7 1 2 91372 100661
0 36618 7 1 2 100659 36617
0 36619 7 1 2 36614 36618
0 36620 5 1 1 36619
0 36621 7 1 2 64285 36620
0 36622 7 1 2 36607 36621
0 36623 5 1 1 36622
0 36624 7 1 2 36571 36623
0 36625 5 1 1 36624
0 36626 7 3 2 66522 92551
0 36627 5 1 1 100667
0 36628 7 1 2 35453 36627
0 36629 5 13 1 36628
0 36630 7 17 2 69400 100362
0 36631 5 1 1 100683
0 36632 7 1 2 86471 100684
0 36633 5 1 1 36632
0 36634 7 6 2 66249 92803
0 36635 7 2 2 83856 100700
0 36636 5 1 1 100706
0 36637 7 1 2 36633 36636
0 36638 5 1 1 36637
0 36639 7 1 2 67488 36638
0 36640 5 1 1 36639
0 36641 7 1 2 93488 100685
0 36642 5 1 1 36641
0 36643 7 1 2 36640 36642
0 36644 5 1 1 36643
0 36645 7 1 2 97986 36644
0 36646 5 1 1 36645
0 36647 7 1 2 99721 98570
0 36648 5 1 1 36647
0 36649 7 1 2 36646 36648
0 36650 5 1 1 36649
0 36651 7 1 2 88823 36650
0 36652 5 1 1 36651
0 36653 7 1 2 67489 100707
0 36654 5 1 1 36653
0 36655 7 2 2 65476 86840
0 36656 7 1 2 100686 100708
0 36657 5 1 1 36656
0 36658 7 1 2 36654 36657
0 36659 5 1 1 36658
0 36660 7 4 2 69128 99367
0 36661 7 1 2 78113 100710
0 36662 7 1 2 36659 36661
0 36663 5 1 1 36662
0 36664 7 1 2 36652 36663
0 36665 5 1 1 36664
0 36666 7 1 2 66139 36665
0 36667 5 1 1 36666
0 36668 7 1 2 35253 97531
0 36669 5 1 1 36668
0 36670 7 1 2 99722 36669
0 36671 5 1 1 36670
0 36672 7 3 2 96412 99752
0 36673 5 1 1 100714
0 36674 7 1 2 100715 100386
0 36675 5 1 1 36674
0 36676 7 1 2 36671 36675
0 36677 5 1 1 36676
0 36678 7 1 2 63602 36677
0 36679 5 1 1 36678
0 36680 7 3 2 61382 69239
0 36681 7 1 2 75113 99791
0 36682 7 1 2 100717 36681
0 36683 5 1 1 36682
0 36684 7 1 2 36679 36683
0 36685 5 1 1 36684
0 36686 7 1 2 65477 36685
0 36687 5 1 1 36686
0 36688 7 1 2 86862 88167
0 36689 7 1 2 100660 36688
0 36690 5 1 1 36689
0 36691 7 1 2 36687 36690
0 36692 5 1 1 36691
0 36693 7 1 2 65183 97714
0 36694 7 1 2 36692 36693
0 36695 5 1 1 36694
0 36696 7 1 2 36667 36695
0 36697 5 1 1 36696
0 36698 7 1 2 81373 36697
0 36699 5 1 1 36698
0 36700 7 2 2 66250 71675
0 36701 7 4 2 64548 65805
0 36702 7 2 2 97987 100722
0 36703 7 1 2 100720 100726
0 36704 5 1 1 36703
0 36705 7 1 2 88168 94636
0 36706 5 1 1 36705
0 36707 7 1 2 36704 36706
0 36708 5 1 1 36707
0 36709 7 1 2 66140 36708
0 36710 5 1 1 36709
0 36711 7 2 2 64286 99616
0 36712 7 1 2 100728 99792
0 36713 5 1 1 36712
0 36714 7 1 2 36710 36713
0 36715 5 1 1 36714
0 36716 7 1 2 65478 36715
0 36717 5 1 1 36716
0 36718 7 2 2 92835 98139
0 36719 7 2 2 65806 87496
0 36720 7 1 2 100732 97353
0 36721 7 1 2 100730 36720
0 36722 5 1 1 36721
0 36723 7 1 2 36717 36722
0 36724 5 1 1 36723
0 36725 7 1 2 93696 36724
0 36726 5 1 1 36725
0 36727 7 1 2 77752 100507
0 36728 7 1 2 100687 36727
0 36729 5 1 1 36728
0 36730 7 1 2 36726 36729
0 36731 5 1 1 36730
0 36732 7 1 2 62168 36731
0 36733 5 1 1 36732
0 36734 7 4 2 69401 70407
0 36735 7 1 2 86841 100734
0 36736 7 1 2 98736 98863
0 36737 7 1 2 36735 36736
0 36738 5 1 1 36737
0 36739 7 1 2 36733 36738
0 36740 5 1 1 36739
0 36741 7 1 2 90841 36740
0 36742 5 1 1 36741
0 36743 7 1 2 36699 36742
0 36744 5 1 1 36743
0 36745 7 1 2 100670 36744
0 36746 5 1 1 36745
0 36747 7 4 2 88921 93166
0 36748 7 1 2 81347 100738
0 36749 5 1 1 36748
0 36750 7 1 2 79754 92804
0 36751 7 1 2 84190 36750
0 36752 5 1 1 36751
0 36753 7 1 2 36749 36752
0 36754 5 1 1 36753
0 36755 7 1 2 62169 36754
0 36756 5 1 1 36755
0 36757 7 1 2 75881 96838
0 36758 7 1 2 100617 36757
0 36759 5 1 1 36758
0 36760 7 1 2 36756 36759
0 36761 5 1 1 36760
0 36762 7 1 2 72387 36761
0 36763 5 1 1 36762
0 36764 7 1 2 94052 100739
0 36765 7 1 2 100372 36764
0 36766 5 1 1 36765
0 36767 7 1 2 36763 36766
0 36768 5 1 1 36767
0 36769 7 1 2 65479 36768
0 36770 5 1 1 36769
0 36771 7 1 2 92414 96831
0 36772 7 1 2 97976 36771
0 36773 7 1 2 95343 36772
0 36774 5 1 1 36773
0 36775 7 1 2 36770 36774
0 36776 5 1 1 36775
0 36777 7 1 2 97309 36776
0 36778 5 1 1 36777
0 36779 7 2 2 84280 94769
0 36780 7 1 2 83386 74925
0 36781 7 1 2 87927 99739
0 36782 7 1 2 36780 36781
0 36783 7 1 2 100742 36782
0 36784 7 1 2 100370 36783
0 36785 5 1 1 36784
0 36786 7 1 2 36778 36785
0 36787 5 1 1 36786
0 36788 7 1 2 93800 36787
0 36789 5 1 1 36788
0 36790 7 1 2 79370 76374
0 36791 7 1 2 97345 36790
0 36792 7 2 2 95930 99193
0 36793 7 3 2 92836 94053
0 36794 7 1 2 86279 100746
0 36795 7 1 2 100744 36794
0 36796 7 1 2 36791 36795
0 36797 5 1 1 36796
0 36798 7 1 2 95344 100153
0 36799 5 1 1 36798
0 36800 7 1 2 78196 87858
0 36801 7 1 2 88177 36800
0 36802 7 1 2 98747 36801
0 36803 5 1 1 36802
0 36804 7 1 2 36799 36803
0 36805 5 1 1 36804
0 36806 7 1 2 61304 36805
0 36807 5 1 1 36806
0 36808 7 1 2 97519 97529
0 36809 7 1 2 95345 36808
0 36810 5 1 1 36809
0 36811 7 1 2 36807 36810
0 36812 5 1 1 36811
0 36813 7 1 2 84148 98155
0 36814 7 1 2 36812 36813
0 36815 5 1 1 36814
0 36816 7 1 2 36797 36815
0 36817 7 1 2 36789 36816
0 36818 5 1 1 36817
0 36819 7 1 2 76174 36818
0 36820 5 1 1 36819
0 36821 7 1 2 36746 36820
0 36822 7 1 2 36625 36821
0 36823 5 1 1 36822
0 36824 7 1 2 72171 36823
0 36825 5 1 1 36824
0 36826 7 2 2 93600 97715
0 36827 7 3 2 61383 100671
0 36828 5 1 1 100751
0 36829 7 3 2 99020 98105
0 36830 5 1 1 100754
0 36831 7 2 2 36828 36830
0 36832 5 6 1 100757
0 36833 7 4 2 69402 100759
0 36834 7 1 2 96228 100765
0 36835 5 1 1 36834
0 36836 7 3 2 62609 63031
0 36837 7 1 2 64549 100769
0 36838 5 1 1 36837
0 36839 7 2 2 67874 90866
0 36840 5 1 1 100772
0 36841 7 1 2 62878 100773
0 36842 5 1 1 36841
0 36843 7 1 2 36838 36842
0 36844 5 1 1 36843
0 36845 7 1 2 61384 36844
0 36846 5 1 1 36845
0 36847 7 1 2 84561 100255
0 36848 5 1 1 36847
0 36849 7 1 2 36846 36848
0 36850 5 1 1 36849
0 36851 7 1 2 72635 36850
0 36852 5 1 1 36851
0 36853 7 1 2 84516 99161
0 36854 5 1 1 36853
0 36855 7 1 2 85286 73968
0 36856 5 1 1 36855
0 36857 7 4 2 70947 93801
0 36858 7 1 2 69403 100774
0 36859 7 1 2 36856 36858
0 36860 5 1 1 36859
0 36861 7 1 2 36854 36860
0 36862 7 1 2 36852 36861
0 36863 5 1 1 36862
0 36864 7 1 2 77249 36863
0 36865 5 1 1 36864
0 36866 7 3 2 67875 90905
0 36867 5 1 1 100778
0 36868 7 1 2 36867 100306
0 36869 5 1 1 36868
0 36870 7 1 2 77250 36869
0 36871 5 1 1 36870
0 36872 7 1 2 82334 100770
0 36873 5 1 1 36872
0 36874 7 1 2 36871 36873
0 36875 5 1 1 36874
0 36876 7 1 2 61385 36875
0 36877 5 1 1 36876
0 36878 7 2 2 66251 94830
0 36879 7 1 2 63188 99697
0 36880 7 1 2 100781 36879
0 36881 5 1 1 36880
0 36882 7 1 2 36877 36881
0 36883 5 1 1 36882
0 36884 7 1 2 95969 36883
0 36885 5 1 1 36884
0 36886 7 2 2 89670 92194
0 36887 7 1 2 72791 99698
0 36888 7 1 2 100783 36887
0 36889 5 1 1 36888
0 36890 7 1 2 36885 36889
0 36891 7 1 2 36865 36890
0 36892 5 1 1 36891
0 36893 7 1 2 70740 36892
0 36894 5 1 1 36893
0 36895 7 1 2 36835 36894
0 36896 5 1 1 36895
0 36897 7 1 2 100749 36896
0 36898 5 1 1 36897
0 36899 7 1 2 100647 97704
0 36900 5 2 1 36899
0 36901 7 1 2 65480 100785
0 36902 7 1 2 36898 36901
0 36903 5 1 1 36902
0 36904 7 2 2 61630 95152
0 36905 7 1 2 91011 96360
0 36906 5 1 1 36905
0 36907 7 1 2 91022 96648
0 36908 5 1 1 36907
0 36909 7 1 2 36906 36908
0 36910 5 1 1 36909
0 36911 7 1 2 92805 36910
0 36912 5 1 1 36911
0 36913 7 1 2 84583 99336
0 36914 5 1 1 36913
0 36915 7 8 2 66252 67490
0 36916 7 1 2 100789 98124
0 36917 5 1 1 36916
0 36918 7 1 2 36914 36917
0 36919 5 1 1 36918
0 36920 7 1 2 96865 96947
0 36921 7 1 2 36919 36920
0 36922 5 1 1 36921
0 36923 7 1 2 36912 36922
0 36924 5 1 1 36923
0 36925 7 1 2 70948 36924
0 36926 5 1 1 36925
0 36927 7 2 2 75899 97115
0 36928 5 1 1 100797
0 36929 7 1 2 159 94498
0 36930 5 1 1 36929
0 36931 7 1 2 72388 36930
0 36932 5 1 1 36931
0 36933 7 1 2 36928 36932
0 36934 5 1 1 36933
0 36935 7 3 2 90997 92806
0 36936 7 1 2 90981 100799
0 36937 7 1 2 36934 36936
0 36938 5 1 1 36937
0 36939 7 1 2 36926 36938
0 36940 5 1 1 36939
0 36941 7 1 2 100787 36940
0 36942 5 1 1 36941
0 36943 7 3 2 66253 69240
0 36944 7 12 2 64550 100802
0 36945 7 1 2 71129 72389
0 36946 5 1 1 36945
0 36947 7 2 2 72832 72758
0 36948 7 1 2 67491 100817
0 36949 5 1 1 36948
0 36950 7 1 2 36946 36949
0 36951 5 1 1 36950
0 36952 7 1 2 66016 36951
0 36953 5 1 1 36952
0 36954 7 1 2 25789 36953
0 36955 5 1 1 36954
0 36956 7 1 2 100805 36955
0 36957 5 1 1 36956
0 36958 7 1 2 84900 100688
0 36959 5 1 1 36958
0 36960 7 1 2 36957 36959
0 36961 5 1 1 36960
0 36962 7 1 2 96958 36961
0 36963 5 1 1 36962
0 36964 7 2 2 96729 100790
0 36965 5 1 1 100819
0 36966 7 6 2 61386 93123
0 36967 5 1 1 100821
0 36968 7 1 2 76741 100822
0 36969 5 1 1 36968
0 36970 7 1 2 36965 36969
0 36971 5 1 1 36970
0 36972 7 3 2 69129 65807
0 36973 7 2 2 92643 100827
0 36974 7 1 2 83466 100830
0 36975 7 1 2 36971 36974
0 36976 5 1 1 36975
0 36977 7 1 2 36963 36976
0 36978 5 1 1 36977
0 36979 7 1 2 100672 36978
0 36980 5 1 1 36979
0 36981 7 1 2 92837 99959
0 36982 7 1 2 96605 36981
0 36983 5 1 1 36982
0 36984 7 2 2 99274 99904
0 36985 7 1 2 61305 92807
0 36986 7 1 2 100832 36985
0 36987 5 1 1 36986
0 36988 7 1 2 36983 36987
0 36989 5 1 1 36988
0 36990 7 1 2 72561 36989
0 36991 5 1 1 36990
0 36992 7 4 2 99617 99565
0 36993 7 1 2 96197 100834
0 36994 5 1 1 36993
0 36995 7 1 2 36991 36994
0 36996 5 1 1 36995
0 36997 7 1 2 65808 36996
0 36998 5 1 1 36997
0 36999 7 1 2 100835 100798
0 37000 5 1 1 36999
0 37001 7 1 2 36998 37000
0 37002 5 1 1 37001
0 37003 7 1 2 100589 37002
0 37004 5 1 1 37003
0 37005 7 2 2 66254 84230
0 37006 5 1 1 100838
0 37007 7 1 2 100839 97550
0 37008 5 1 1 37007
0 37009 7 1 2 96730 100613
0 37010 5 1 1 37009
0 37011 7 1 2 37008 37010
0 37012 5 1 1 37011
0 37013 7 5 2 62170 91865
0 37014 7 2 2 69130 66017
0 37015 7 1 2 90529 100845
0 37016 7 2 2 100840 37015
0 37017 5 2 1 100847
0 37018 7 1 2 65809 100848
0 37019 7 1 2 37012 37018
0 37020 5 1 1 37019
0 37021 7 1 2 70408 37020
0 37022 7 1 2 37004 37021
0 37023 7 1 2 36980 37022
0 37024 7 1 2 36942 37023
0 37025 5 1 1 37024
0 37026 7 1 2 82569 37025
0 37027 7 1 2 36903 37026
0 37028 5 1 1 37027
0 37029 7 3 2 69241 91023
0 37030 7 1 2 62171 81093
0 37031 7 1 2 96216 37030
0 37032 5 1 1 37031
0 37033 7 2 2 77173 81670
0 37034 7 1 2 69404 100854
0 37035 7 1 2 72308 37034
0 37036 5 1 1 37035
0 37037 7 1 2 37032 37036
0 37038 5 1 1 37037
0 37039 7 2 2 79608 82551
0 37040 7 1 2 37038 100856
0 37041 5 1 1 37040
0 37042 7 1 2 90418 77860
0 37043 5 1 1 37042
0 37044 7 1 2 93936 37043
0 37045 5 1 1 37044
0 37046 7 1 2 82335 37045
0 37047 5 1 1 37046
0 37048 7 1 2 81094 96276
0 37049 5 1 1 37048
0 37050 7 1 2 37047 37049
0 37051 5 1 1 37050
0 37052 7 1 2 68444 37051
0 37053 5 1 1 37052
0 37054 7 2 2 82760 84260
0 37055 7 1 2 87216 100858
0 37056 5 1 1 37055
0 37057 7 1 2 37056 97695
0 37058 5 1 1 37057
0 37059 7 1 2 63603 37058
0 37060 5 1 1 37059
0 37061 7 2 2 69405 74186
0 37062 7 1 2 80955 93376
0 37063 7 1 2 100860 37062
0 37064 5 1 1 37063
0 37065 7 1 2 65481 37064
0 37066 7 1 2 37060 37065
0 37067 7 1 2 37053 37066
0 37068 5 1 1 37067
0 37069 7 1 2 67711 96361
0 37070 5 1 1 37069
0 37071 7 1 2 73759 37070
0 37072 5 1 1 37071
0 37073 7 1 2 77933 37072
0 37074 5 1 1 37073
0 37075 7 3 2 68866 76328
0 37076 7 1 2 84759 100862
0 37077 5 1 1 37076
0 37078 7 1 2 37074 37077
0 37079 5 1 1 37078
0 37080 7 1 2 82336 37079
0 37081 5 1 1 37080
0 37082 7 1 2 83818 90242
0 37083 7 1 2 100431 37082
0 37084 5 1 1 37083
0 37085 7 1 2 37081 37084
0 37086 5 1 1 37085
0 37087 7 1 2 64158 37086
0 37088 5 1 1 37087
0 37089 7 1 2 91111 97069
0 37090 5 2 1 37089
0 37091 7 1 2 80652 87019
0 37092 7 1 2 91895 37091
0 37093 7 1 2 100865 37092
0 37094 5 1 1 37093
0 37095 7 1 2 70409 37094
0 37096 7 1 2 37088 37095
0 37097 5 1 1 37096
0 37098 7 1 2 88274 37097
0 37099 7 1 2 37068 37098
0 37100 5 1 1 37099
0 37101 7 1 2 37041 37100
0 37102 5 1 1 37101
0 37103 7 1 2 100851 37102
0 37104 5 1 1 37103
0 37105 7 1 2 80985 85655
0 37106 7 1 2 88341 37105
0 37107 5 1 1 37106
0 37108 7 1 2 31331 37107
0 37109 5 1 1 37108
0 37110 7 1 2 71343 37109
0 37111 5 1 1 37110
0 37112 7 1 2 82337 84938
0 37113 5 1 1 37112
0 37114 7 1 2 81117 37113
0 37115 5 1 1 37114
0 37116 7 1 2 73478 37115
0 37117 5 1 1 37116
0 37118 7 1 2 77819 83844
0 37119 5 1 1 37118
0 37120 7 1 2 37117 37119
0 37121 5 1 1 37120
0 37122 7 1 2 64159 37121
0 37123 5 1 1 37122
0 37124 7 3 2 77251 88900
0 37125 5 1 1 100867
0 37126 7 1 2 78379 92013
0 37127 5 1 1 37126
0 37128 7 1 2 37125 37127
0 37129 5 1 1 37128
0 37130 7 1 2 72562 37129
0 37131 5 1 1 37130
0 37132 7 2 2 89549 82443
0 37133 5 1 1 100870
0 37134 7 1 2 3594 37133
0 37135 5 1 1 37134
0 37136 7 1 2 98294 37135
0 37137 5 1 1 37136
0 37138 7 1 2 81095 89945
0 37139 5 1 1 37138
0 37140 7 1 2 37137 37139
0 37141 7 1 2 37131 37140
0 37142 7 1 2 37123 37141
0 37143 5 1 1 37142
0 37144 7 1 2 70410 37143
0 37145 5 1 1 37144
0 37146 7 1 2 37111 37145
0 37147 5 1 1 37146
0 37148 7 1 2 90842 37147
0 37149 5 1 1 37148
0 37150 7 1 2 88275 84245
0 37151 7 1 2 97702 37150
0 37152 5 1 1 37151
0 37153 7 1 2 37149 37152
0 37154 5 1 1 37153
0 37155 7 1 2 63604 37154
0 37156 5 1 1 37155
0 37157 7 1 2 65482 93567
0 37158 5 3 1 37157
0 37159 7 6 2 65810 98295
0 37160 5 1 1 100875
0 37161 7 3 2 70411 100876
0 37162 5 1 1 100881
0 37163 7 1 2 75728 93965
0 37164 5 2 1 37163
0 37165 7 1 2 37162 100884
0 37166 5 1 1 37165
0 37167 7 1 2 62879 37166
0 37168 5 1 1 37167
0 37169 7 1 2 100872 37168
0 37170 5 1 1 37169
0 37171 7 1 2 82338 37170
0 37172 5 1 1 37171
0 37173 7 1 2 78222 84037
0 37174 5 1 1 37173
0 37175 7 1 2 62880 37174
0 37176 5 1 1 37175
0 37177 7 1 2 71344 78216
0 37178 5 1 1 37177
0 37179 7 1 2 76610 100885
0 37180 7 1 2 37178 37179
0 37181 7 1 2 37176 37180
0 37182 5 1 1 37181
0 37183 7 1 2 81096 37182
0 37184 5 1 1 37183
0 37185 7 1 2 37172 37184
0 37186 5 1 1 37185
0 37187 7 2 2 83680 81130
0 37188 7 1 2 37186 100886
0 37189 5 1 1 37188
0 37190 7 1 2 82710 92886
0 37191 7 1 2 92581 94540
0 37192 7 1 2 37190 37191
0 37193 5 1 1 37192
0 37194 7 1 2 37189 37193
0 37195 7 1 2 37156 37194
0 37196 5 1 1 37195
0 37197 7 1 2 91357 37196
0 37198 5 1 1 37197
0 37199 7 1 2 37104 37198
0 37200 5 1 1 37199
0 37201 7 1 2 64287 37200
0 37202 5 1 1 37201
0 37203 7 1 2 37028 37202
0 37204 7 1 2 36825 37203
0 37205 7 2 2 72636 83958
0 37206 5 3 1 100888
0 37207 7 1 2 90264 85333
0 37208 5 1 1 37207
0 37209 7 1 2 100890 37208
0 37210 5 1 1 37209
0 37211 7 1 2 73479 37210
0 37212 5 2 1 37211
0 37213 7 5 2 67712 98296
0 37214 5 9 1 100895
0 37215 7 1 2 94929 100900
0 37216 5 3 1 37215
0 37217 7 1 2 83959 100909
0 37218 5 1 1 37217
0 37219 7 1 2 100893 37218
0 37220 5 1 1 37219
0 37221 7 1 2 86062 37220
0 37222 5 1 1 37221
0 37223 7 1 2 90314 87149
0 37224 5 1 1 37223
0 37225 7 1 2 88380 89265
0 37226 7 1 2 85274 37225
0 37227 5 1 1 37226
0 37228 7 1 2 37224 37227
0 37229 5 1 1 37228
0 37230 7 1 2 93941 37229
0 37231 5 1 1 37230
0 37232 7 1 2 37222 37231
0 37233 5 1 1 37232
0 37234 7 1 2 68445 37233
0 37235 5 1 1 37234
0 37236 7 2 2 64551 80245
0 37237 7 1 2 97042 100912
0 37238 5 1 1 37237
0 37239 7 1 2 100894 37238
0 37240 5 1 1 37239
0 37241 7 1 2 90334 37240
0 37242 5 1 1 37241
0 37243 7 1 2 37235 37242
0 37244 5 1 1 37243
0 37245 7 1 2 63189 37244
0 37246 5 1 1 37245
0 37247 7 1 2 95864 100437
0 37248 5 1 1 37247
0 37249 7 1 2 64160 37248
0 37250 5 1 1 37249
0 37251 7 1 2 84644 37250
0 37252 5 1 1 37251
0 37253 7 1 2 86063 37252
0 37254 5 1 1 37253
0 37255 7 1 2 67013 100268
0 37256 5 1 1 37255
0 37257 7 1 2 37254 37256
0 37258 5 1 1 37257
0 37259 7 1 2 80913 92014
0 37260 7 1 2 37258 37259
0 37261 5 1 1 37260
0 37262 7 1 2 37246 37261
0 37263 5 1 1 37262
0 37264 7 1 2 68210 37263
0 37265 5 1 1 37264
0 37266 7 2 2 64770 82117
0 37267 7 2 2 71345 100914
0 37268 7 1 2 88001 100916
0 37269 5 1 1 37268
0 37270 7 1 2 37269 97766
0 37271 5 1 1 37270
0 37272 7 1 2 74709 98273
0 37273 7 1 2 37271 37272
0 37274 5 1 1 37273
0 37275 7 1 2 37265 37274
0 37276 5 1 1 37275
0 37277 7 1 2 65184 37276
0 37278 5 1 1 37277
0 37279 7 1 2 80640 79324
0 37280 7 1 2 91825 92582
0 37281 7 1 2 37279 37280
0 37282 5 1 1 37281
0 37283 7 1 2 37278 37282
0 37284 5 1 1 37283
0 37285 7 1 2 92673 37284
0 37286 5 1 1 37285
0 37287 7 2 2 89444 80884
0 37288 7 1 2 80630 73740
0 37289 7 1 2 100918 37288
0 37290 5 1 1 37289
0 37291 7 2 2 64771 71169
0 37292 7 1 2 82118 100920
0 37293 5 1 1 37292
0 37294 7 1 2 100891 37293
0 37295 5 1 1 37294
0 37296 7 1 2 63190 37295
0 37297 5 1 1 37296
0 37298 7 2 2 87144 91723
0 37299 5 1 1 100922
0 37300 7 1 2 80052 100923
0 37301 5 1 1 37300
0 37302 7 1 2 37297 37301
0 37303 5 1 1 37302
0 37304 7 1 2 62610 37303
0 37305 5 1 1 37304
0 37306 7 5 2 79371 74987
0 37307 7 1 2 77252 100924
0 37308 5 1 1 37307
0 37309 7 1 2 37305 37308
0 37310 5 1 1 37309
0 37311 7 1 2 68867 75164
0 37312 7 1 2 37310 37311
0 37313 5 1 1 37312
0 37314 7 1 2 37290 37313
0 37315 5 1 1 37314
0 37316 7 1 2 89110 37315
0 37317 5 1 1 37316
0 37318 7 1 2 74506 95944
0 37319 5 1 1 37318
0 37320 7 1 2 86975 37319
0 37321 5 1 1 37320
0 37322 7 1 2 80070 97080
0 37323 5 1 1 37322
0 37324 7 1 2 37321 37323
0 37325 5 1 1 37324
0 37326 7 1 2 92539 95493
0 37327 7 1 2 37325 37326
0 37328 5 1 1 37327
0 37329 7 1 2 37317 37328
0 37330 5 1 1 37329
0 37331 7 1 2 65811 37330
0 37332 5 1 1 37331
0 37333 7 1 2 77540 95977
0 37334 5 1 1 37333
0 37335 7 1 2 82557 37334
0 37336 5 1 1 37335
0 37337 7 1 2 77280 100901
0 37338 5 2 1 37337
0 37339 7 1 2 81252 82565
0 37340 7 1 2 100929 37339
0 37341 5 1 1 37340
0 37342 7 1 2 37336 37341
0 37343 5 1 1 37342
0 37344 7 1 2 63191 37343
0 37345 5 1 1 37344
0 37346 7 1 2 74602 81742
0 37347 7 1 2 81028 37346
0 37348 7 1 2 96656 37347
0 37349 5 1 1 37348
0 37350 7 1 2 37345 37349
0 37351 5 1 1 37350
0 37352 7 1 2 82854 94054
0 37353 7 1 2 37351 37352
0 37354 5 1 1 37353
0 37355 7 1 2 37332 37354
0 37356 5 1 1 37355
0 37357 7 1 2 65483 37356
0 37358 5 1 1 37357
0 37359 7 1 2 88373 89484
0 37360 5 1 1 37359
0 37361 7 1 2 72792 81473
0 37362 7 1 2 84254 37361
0 37363 5 1 1 37362
0 37364 7 1 2 37360 37363
0 37365 5 1 1 37364
0 37366 7 1 2 80421 37365
0 37367 5 1 1 37366
0 37368 7 1 2 86932 73219
0 37369 7 1 2 89916 80745
0 37370 7 1 2 37368 37369
0 37371 5 1 1 37370
0 37372 7 1 2 37367 37371
0 37373 5 1 1 37372
0 37374 7 1 2 91287 94831
0 37375 7 1 2 37373 37374
0 37376 5 1 1 37375
0 37377 7 1 2 37358 37376
0 37378 5 1 1 37377
0 37379 7 1 2 93518 37378
0 37380 5 1 1 37379
0 37381 7 1 2 37286 37380
0 37382 5 1 1 37381
0 37383 7 1 2 69131 37382
0 37384 5 1 1 37383
0 37385 7 1 2 94953 95260
0 37386 5 1 1 37385
0 37387 7 1 2 94774 100788
0 37388 5 1 1 37387
0 37389 7 1 2 37386 37388
0 37390 5 1 1 37389
0 37391 7 1 2 93861 37390
0 37392 5 1 1 37391
0 37393 7 1 2 72067 72934
0 37394 5 1 1 37393
0 37395 7 1 2 100416 37394
0 37396 5 1 1 37395
0 37397 7 1 2 96593 37396
0 37398 5 1 1 37397
0 37399 7 1 2 100461 37398
0 37400 5 1 1 37399
0 37401 7 1 2 65812 37400
0 37402 5 1 1 37401
0 37403 7 1 2 82761 96803
0 37404 5 1 1 37403
0 37405 7 1 2 77253 84571
0 37406 7 1 2 96858 37405
0 37407 5 1 1 37406
0 37408 7 1 2 37404 37407
0 37409 5 1 1 37408
0 37410 7 1 2 64161 37409
0 37411 5 1 1 37410
0 37412 7 1 2 89675 96136
0 37413 5 1 1 37412
0 37414 7 1 2 37411 37413
0 37415 5 1 1 37414
0 37416 7 1 2 67492 37415
0 37417 5 1 1 37416
0 37418 7 1 2 85535 96387
0 37419 5 1 1 37418
0 37420 7 1 2 37417 37419
0 37421 7 1 2 37402 37420
0 37422 5 1 1 37421
0 37423 7 1 2 97310 37422
0 37424 5 1 1 37423
0 37425 7 1 2 37392 37424
0 37426 5 1 1 37425
0 37427 7 1 2 65484 37426
0 37428 5 1 1 37427
0 37429 7 1 2 82359 96606
0 37430 5 1 1 37429
0 37431 7 1 2 95398 96816
0 37432 5 1 1 37431
0 37433 7 1 2 37430 37432
0 37434 5 1 1 37433
0 37435 7 1 2 93714 100493
0 37436 7 1 2 37434 37435
0 37437 5 1 1 37436
0 37438 7 1 2 37428 37437
0 37439 5 1 1 37438
0 37440 7 1 2 89917 37439
0 37441 5 1 1 37440
0 37442 7 1 2 84572 85287
0 37443 5 2 1 37442
0 37444 7 1 2 70949 87095
0 37445 7 1 2 83781 37444
0 37446 7 3 2 69406 87685
0 37447 7 1 2 100933 99912
0 37448 7 1 2 37445 37447
0 37449 7 1 2 100931 37448
0 37450 5 1 1 37449
0 37451 7 1 2 37441 37450
0 37452 5 1 1 37451
0 37453 7 1 2 69600 37452
0 37454 5 1 1 37453
0 37455 7 1 2 90243 97988
0 37456 7 1 2 96632 37455
0 37457 7 2 2 81824 92808
0 37458 7 1 2 99539 100936
0 37459 7 1 2 37456 37458
0 37460 5 1 1 37459
0 37461 7 1 2 37454 37460
0 37462 5 1 1 37461
0 37463 7 1 2 93802 37462
0 37464 5 1 1 37463
0 37465 7 2 2 68031 93124
0 37466 7 3 2 66523 100938
0 37467 7 1 2 99691 100940
0 37468 5 1 1 37467
0 37469 7 1 2 63983 87773
0 37470 7 1 2 83850 37469
0 37471 5 1 1 37470
0 37472 7 1 2 37468 37471
0 37473 5 1 1 37472
0 37474 7 1 2 70741 37473
0 37475 5 1 1 37474
0 37476 7 1 2 72349 99546
0 37477 5 1 1 37476
0 37478 7 1 2 87731 75367
0 37479 5 1 1 37478
0 37480 7 1 2 37477 37479
0 37481 5 1 1 37480
0 37482 7 1 2 81097 37481
0 37483 5 1 1 37482
0 37484 7 1 2 37475 37483
0 37485 5 1 1 37484
0 37486 7 1 2 65485 37485
0 37487 5 1 1 37486
0 37488 7 1 2 83845 97551
0 37489 5 1 1 37488
0 37490 7 1 2 37489 97537
0 37491 5 1 1 37490
0 37492 7 1 2 72462 37491
0 37493 5 1 1 37492
0 37494 7 1 2 37487 37493
0 37495 5 1 1 37494
0 37496 7 1 2 69019 37495
0 37497 5 1 1 37496
0 37498 7 1 2 82296 98869
0 37499 5 1 1 37498
0 37500 7 1 2 87732 100871
0 37501 5 1 1 37500
0 37502 7 1 2 37499 37501
0 37503 5 1 1 37502
0 37504 7 1 2 85380 37503
0 37505 5 1 1 37504
0 37506 7 1 2 37497 37505
0 37507 5 1 1 37506
0 37508 7 1 2 66018 37507
0 37509 5 1 1 37508
0 37510 7 2 2 67493 84018
0 37511 7 1 2 87850 97387
0 37512 5 1 1 37511
0 37513 7 3 2 61306 80986
0 37514 7 1 2 72328 93125
0 37515 7 1 2 100945 37514
0 37516 5 1 1 37515
0 37517 7 1 2 37512 37516
0 37518 5 1 1 37517
0 37519 7 1 2 100943 37518
0 37520 5 1 1 37519
0 37521 7 1 2 37509 37520
0 37522 5 1 1 37521
0 37523 7 1 2 98015 37522
0 37524 5 1 1 37523
0 37525 7 2 2 76715 99154
0 37526 7 1 2 82339 100948
0 37527 5 1 1 37526
0 37528 7 2 2 77254 93738
0 37529 7 1 2 94954 100950
0 37530 5 1 1 37529
0 37531 7 1 2 86752 22020
0 37532 5 1 1 37531
0 37533 7 1 2 67494 37532
0 37534 5 1 1 37533
0 37535 7 1 2 74083 86472
0 37536 5 1 1 37535
0 37537 7 1 2 85381 72350
0 37538 5 1 1 37537
0 37539 7 1 2 37536 37538
0 37540 5 1 1 37539
0 37541 7 1 2 66019 37540
0 37542 5 1 1 37541
0 37543 7 1 2 37534 37542
0 37544 5 1 1 37543
0 37545 7 1 2 82340 37544
0 37546 5 1 1 37545
0 37547 7 1 2 37530 37546
0 37548 5 1 1 37547
0 37549 7 1 2 98886 37548
0 37550 5 1 1 37549
0 37551 7 1 2 84078 97739
0 37552 7 1 2 99397 37551
0 37553 5 1 1 37552
0 37554 7 1 2 37550 37553
0 37555 5 1 1 37554
0 37556 7 1 2 90716 37555
0 37557 5 1 1 37556
0 37558 7 1 2 37527 37557
0 37559 7 1 2 37524 37558
0 37560 5 1 1 37559
0 37561 7 1 2 69601 89918
0 37562 7 1 2 37560 37561
0 37563 5 1 1 37562
0 37564 7 1 2 37464 37563
0 37565 5 1 1 37564
0 37566 7 1 2 94944 37565
0 37567 5 1 1 37566
0 37568 7 1 2 37384 37567
0 37569 7 1 2 37204 37568
0 37570 7 1 2 36471 37569
0 37571 7 1 2 36326 37570
0 37572 7 1 2 35937 37571
0 37573 5 1 1 37572
0 37574 7 1 2 73030 37573
0 37575 5 1 1 37574
0 37576 7 1 2 71254 72292
0 37577 5 3 1 37576
0 37578 7 1 2 67495 85170
0 37579 5 1 1 37578
0 37580 7 1 2 85933 37579
0 37581 5 1 1 37580
0 37582 7 1 2 64162 37581
0 37583 5 1 1 37582
0 37584 7 1 2 100952 37583
0 37585 5 1 1 37584
0 37586 7 1 2 63825 37585
0 37587 5 1 1 37586
0 37588 7 1 2 72563 97925
0 37589 5 1 1 37588
0 37590 7 1 2 37587 37589
0 37591 5 1 1 37590
0 37592 7 1 2 80710 37591
0 37593 5 1 1 37592
0 37594 7 3 2 63984 78197
0 37595 7 1 2 68684 85867
0 37596 7 1 2 100955 37595
0 37597 5 1 1 37596
0 37598 7 1 2 37593 37597
0 37599 5 1 1 37598
0 37600 7 1 2 67014 37599
0 37601 5 1 1 37600
0 37602 7 1 2 63605 80862
0 37603 5 2 1 37602
0 37604 7 1 2 70115 93332
0 37605 5 1 1 37604
0 37606 7 1 2 100958 37605
0 37607 5 1 1 37606
0 37608 7 1 2 67713 37607
0 37609 5 1 1 37608
0 37610 7 1 2 78114 78007
0 37611 5 1 1 37610
0 37612 7 1 2 37609 37611
0 37613 5 1 1 37612
0 37614 7 1 2 73814 85517
0 37615 7 1 2 37613 37614
0 37616 5 1 1 37615
0 37617 7 1 2 37601 37616
0 37618 5 1 1 37617
0 37619 7 1 2 65486 37618
0 37620 5 1 1 37619
0 37621 7 1 2 84353 96255
0 37622 7 1 2 91621 37621
0 37623 5 1 1 37622
0 37624 7 1 2 37620 37623
0 37625 5 1 1 37624
0 37626 7 1 2 68211 37625
0 37627 5 1 1 37626
0 37628 7 1 2 81205 86586
0 37629 7 1 2 94530 37628
0 37630 5 1 1 37629
0 37631 7 1 2 37627 37630
0 37632 5 1 1 37631
0 37633 7 1 2 95261 37632
0 37634 5 1 1 37633
0 37635 7 2 2 67015 90153
0 37636 7 1 2 77820 100960
0 37637 5 1 1 37636
0 37638 7 2 2 66020 79053
0 37639 7 1 2 63377 100962
0 37640 5 1 1 37639
0 37641 7 1 2 88449 90800
0 37642 5 1 1 37641
0 37643 7 1 2 37640 37642
0 37644 5 1 1 37643
0 37645 7 1 2 75076 80839
0 37646 7 1 2 37644 37645
0 37647 5 1 1 37646
0 37648 7 1 2 37637 37647
0 37649 5 1 1 37648
0 37650 7 1 2 64163 37649
0 37651 5 1 1 37650
0 37652 7 1 2 94671 100961
0 37653 5 1 1 37652
0 37654 7 1 2 37651 37653
0 37655 5 1 1 37654
0 37656 7 1 2 62611 37655
0 37657 5 1 1 37656
0 37658 7 1 2 95516 97848
0 37659 5 1 1 37658
0 37660 7 1 2 85424 84679
0 37661 5 1 1 37660
0 37662 7 1 2 37659 37661
0 37663 5 1 1 37662
0 37664 7 1 2 62172 37663
0 37665 5 1 1 37664
0 37666 7 1 2 86504 95087
0 37667 5 1 1 37666
0 37668 7 1 2 94468 37667
0 37669 5 1 1 37668
0 37670 7 1 2 95468 37669
0 37671 5 1 1 37670
0 37672 7 1 2 37665 37671
0 37673 5 1 1 37672
0 37674 7 1 2 72172 37673
0 37675 5 1 1 37674
0 37676 7 1 2 68685 84043
0 37677 5 1 1 37676
0 37678 7 1 2 94195 37677
0 37679 5 1 1 37678
0 37680 7 1 2 78659 81844
0 37681 7 1 2 37679 37680
0 37682 5 1 1 37681
0 37683 7 1 2 37675 37682
0 37684 5 1 1 37683
0 37685 7 1 2 65185 37684
0 37686 5 1 1 37685
0 37687 7 1 2 37657 37686
0 37688 5 1 1 37687
0 37689 7 1 2 63606 37688
0 37690 5 1 1 37689
0 37691 7 1 2 67714 100390
0 37692 5 1 1 37691
0 37693 7 1 2 68446 85556
0 37694 5 1 1 37693
0 37695 7 1 2 94327 37694
0 37696 5 1 1 37695
0 37697 7 1 2 69020 37696
0 37698 5 1 1 37697
0 37699 7 1 2 9324 94777
0 37700 5 1 1 37699
0 37701 7 1 2 68447 37700
0 37702 5 1 1 37701
0 37703 7 1 2 71676 72329
0 37704 7 1 2 80449 37703
0 37705 5 1 1 37704
0 37706 7 1 2 37702 37705
0 37707 7 1 2 37698 37706
0 37708 5 1 1 37707
0 37709 7 1 2 62429 37708
0 37710 5 1 1 37709
0 37711 7 1 2 37692 37710
0 37712 5 1 1 37711
0 37713 7 1 2 63826 37712
0 37714 5 1 1 37713
0 37715 7 1 2 73965 75328
0 37716 7 1 2 74204 37715
0 37717 7 1 2 94224 37716
0 37718 5 1 1 37717
0 37719 7 1 2 67016 37718
0 37720 7 1 2 37714 37719
0 37721 5 1 1 37720
0 37722 7 2 2 74009 71541
0 37723 5 2 1 100964
0 37724 7 1 2 100406 100965
0 37725 5 1 1 37724
0 37726 7 1 2 68448 85086
0 37727 7 1 2 88141 37726
0 37728 5 1 1 37727
0 37729 7 1 2 37725 37728
0 37730 5 1 1 37729
0 37731 7 1 2 65487 37730
0 37732 5 1 1 37731
0 37733 7 1 2 77475 90142
0 37734 5 1 1 37733
0 37735 7 1 2 37732 37734
0 37736 5 1 1 37735
0 37737 7 1 2 68686 37736
0 37738 5 1 1 37737
0 37739 7 1 2 77476 90378
0 37740 7 1 2 86721 37739
0 37741 5 1 1 37740
0 37742 7 1 2 62173 37741
0 37743 7 1 2 37738 37742
0 37744 5 1 1 37743
0 37745 7 1 2 68212 37744
0 37746 7 1 2 37721 37745
0 37747 5 1 1 37746
0 37748 7 1 2 68687 94270
0 37749 5 1 1 37748
0 37750 7 1 2 7063 37749
0 37751 5 2 1 37750
0 37752 7 1 2 71255 100968
0 37753 5 1 1 37752
0 37754 7 1 2 78430 89818
0 37755 5 1 1 37754
0 37756 7 1 2 37753 37755
0 37757 5 1 1 37756
0 37758 7 1 2 67285 37757
0 37759 5 1 1 37758
0 37760 7 1 2 94265 37759
0 37761 5 1 1 37760
0 37762 7 1 2 96891 37761
0 37763 5 1 1 37762
0 37764 7 1 2 37747 37763
0 37765 5 1 1 37764
0 37766 7 1 2 65186 37765
0 37767 5 1 1 37766
0 37768 7 1 2 72337 79207
0 37769 5 1 1 37768
0 37770 7 1 2 72564 74038
0 37771 5 1 1 37770
0 37772 7 1 2 37769 37771
0 37773 5 1 1 37772
0 37774 7 1 2 75882 37773
0 37775 5 1 1 37774
0 37776 7 1 2 67286 94055
0 37777 7 1 2 82824 37776
0 37778 5 1 1 37777
0 37779 7 1 2 37775 37778
0 37780 5 1 1 37779
0 37781 7 1 2 78198 91331
0 37782 7 1 2 37780 37781
0 37783 5 1 1 37782
0 37784 7 1 2 37767 37783
0 37785 5 1 1 37784
0 37786 7 1 2 61631 37785
0 37787 5 1 1 37786
0 37788 7 1 2 37690 37787
0 37789 5 1 1 37788
0 37790 7 1 2 63192 37789
0 37791 5 1 1 37790
0 37792 7 1 2 80677 98238
0 37793 5 1 1 37792
0 37794 7 1 2 65187 86822
0 37795 5 1 1 37794
0 37796 7 1 2 37793 37795
0 37797 5 1 1 37796
0 37798 7 1 2 63607 37797
0 37799 5 1 1 37798
0 37800 7 1 2 79054 86823
0 37801 5 1 1 37800
0 37802 7 1 2 37799 37801
0 37803 5 1 1 37802
0 37804 7 1 2 62612 37803
0 37805 5 1 1 37804
0 37806 7 1 2 86907 91626
0 37807 5 1 1 37806
0 37808 7 1 2 37805 37807
0 37809 5 1 1 37808
0 37810 7 1 2 71853 37809
0 37811 5 1 1 37810
0 37812 7 3 2 88561 75454
0 37813 7 2 2 73220 76596
0 37814 7 1 2 65188 100973
0 37815 7 1 2 100970 37814
0 37816 5 1 1 37815
0 37817 7 1 2 37811 37816
0 37818 5 1 1 37817
0 37819 7 1 2 74226 96740
0 37820 7 1 2 37818 37819
0 37821 5 1 1 37820
0 37822 7 1 2 37791 37821
0 37823 5 1 1 37822
0 37824 7 1 2 94613 37823
0 37825 5 1 1 37824
0 37826 7 1 2 37634 37825
0 37827 5 1 1 37826
0 37828 7 1 2 69602 37827
0 37829 5 1 1 37828
0 37830 7 1 2 79042 94712
0 37831 5 1 1 37830
0 37832 7 1 2 62430 91631
0 37833 7 1 2 94657 37832
0 37834 5 1 1 37833
0 37835 7 1 2 37831 37834
0 37836 5 1 1 37835
0 37837 7 1 2 63827 37836
0 37838 5 1 1 37837
0 37839 7 1 2 80695 94713
0 37840 7 1 2 100209 37839
0 37841 5 1 1 37840
0 37842 7 1 2 37838 37841
0 37843 5 1 1 37842
0 37844 7 1 2 72173 37843
0 37845 5 1 1 37844
0 37846 7 1 2 77903 94614
0 37847 7 1 2 88208 37846
0 37848 5 1 1 37847
0 37849 7 1 2 82970 95262
0 37850 7 1 2 95806 37849
0 37851 5 1 1 37850
0 37852 7 1 2 37848 37851
0 37853 5 1 1 37852
0 37854 7 1 2 71346 37853
0 37855 5 1 1 37854
0 37856 7 1 2 95593 96896
0 37857 5 1 1 37856
0 37858 7 1 2 88375 95104
0 37859 5 1 1 37858
0 37860 7 1 2 37857 37859
0 37861 5 1 1 37860
0 37862 7 1 2 86108 77923
0 37863 7 1 2 37861 37862
0 37864 5 1 1 37863
0 37865 7 1 2 37855 37864
0 37866 7 1 2 37845 37865
0 37867 5 1 1 37866
0 37868 7 1 2 62174 37867
0 37869 5 1 1 37868
0 37870 7 1 2 94257 94790
0 37871 7 1 2 95502 37870
0 37872 7 1 2 100348 37871
0 37873 5 1 1 37872
0 37874 7 1 2 37869 37873
0 37875 5 1 1 37874
0 37876 7 1 2 63378 37875
0 37877 5 1 1 37876
0 37878 7 1 2 85238 23844
0 37879 5 1 1 37878
0 37880 7 1 2 63828 37879
0 37881 5 1 1 37880
0 37882 7 1 2 79685 93962
0 37883 5 1 1 37882
0 37884 7 1 2 37881 37883
0 37885 5 1 1 37884
0 37886 7 2 2 76094 37885
0 37887 5 1 1 100975
0 37888 7 1 2 76054 93321
0 37889 5 1 1 37888
0 37890 7 1 2 37887 37889
0 37891 5 1 1 37890
0 37892 7 1 2 65488 89919
0 37893 7 1 2 95358 37892
0 37894 7 1 2 37891 37893
0 37895 5 1 1 37894
0 37896 7 1 2 63608 37895
0 37897 7 1 2 37877 37896
0 37898 5 1 1 37897
0 37899 7 1 2 88758 75207
0 37900 7 1 2 95526 37899
0 37901 5 1 1 37900
0 37902 7 1 2 81016 95314
0 37903 7 1 2 92223 37902
0 37904 5 1 1 37903
0 37905 7 1 2 37901 37904
0 37906 5 1 1 37905
0 37907 7 1 2 90007 37906
0 37908 5 1 1 37907
0 37909 7 1 2 95528 100976
0 37910 5 1 1 37909
0 37911 7 1 2 37908 37910
0 37912 5 1 1 37911
0 37913 7 1 2 62175 37912
0 37914 5 1 1 37913
0 37915 7 1 2 94486 95507
0 37916 7 3 2 63829 81774
0 37917 7 2 2 66524 86616
0 37918 7 1 2 100977 100980
0 37919 7 1 2 37915 37918
0 37920 5 1 1 37919
0 37921 7 1 2 68449 37920
0 37922 7 1 2 37914 37921
0 37923 5 1 1 37922
0 37924 7 1 2 64772 37923
0 37925 7 1 2 37898 37924
0 37926 5 1 1 37925
0 37927 7 1 2 37829 37926
0 37928 5 1 1 37927
0 37929 7 1 2 93862 37928
0 37930 5 1 1 37929
0 37931 7 2 2 74290 97311
0 37932 7 2 2 85634 100417
0 37933 5 10 1 100984
0 37934 7 1 2 65813 100986
0 37935 5 2 1 37934
0 37936 7 1 2 88111 96995
0 37937 7 1 2 100996 37936
0 37938 5 1 1 37937
0 37939 7 1 2 100982 37938
0 37940 5 1 1 37939
0 37941 7 2 2 85087 96523
0 37942 7 2 2 61307 98438
0 37943 7 1 2 95641 101000
0 37944 7 1 2 100998 37943
0 37945 5 1 1 37944
0 37946 7 1 2 37940 37945
0 37947 5 1 1 37946
0 37948 7 1 2 90965 37947
0 37949 5 1 1 37948
0 37950 7 1 2 74848 85590
0 37951 5 1 1 37950
0 37952 7 1 2 81825 84542
0 37953 7 1 2 93207 37952
0 37954 7 1 2 100072 37953
0 37955 7 1 2 37951 37954
0 37956 5 1 1 37955
0 37957 7 1 2 37949 37956
0 37958 5 1 1 37957
0 37959 7 1 2 93948 37958
0 37960 5 1 1 37959
0 37961 7 1 2 75097 85585
0 37962 5 1 1 37961
0 37963 7 2 2 70742 73921
0 37964 5 1 1 101002
0 37965 7 1 2 85292 101003
0 37966 5 1 1 37965
0 37967 7 1 2 37962 37966
0 37968 5 1 1 37967
0 37969 7 1 2 67287 37968
0 37970 5 1 1 37969
0 37971 7 1 2 74889 78008
0 37972 5 1 1 37971
0 37973 7 1 2 87867 95705
0 37974 5 1 1 37973
0 37975 7 1 2 37972 37974
0 37976 5 1 1 37975
0 37977 7 1 2 68868 37976
0 37978 5 1 1 37977
0 37979 7 1 2 76351 74890
0 37980 5 1 1 37979
0 37981 7 1 2 37978 37980
0 37982 5 1 1 37981
0 37983 7 1 2 67017 37982
0 37984 5 1 1 37983
0 37985 7 1 2 37970 37984
0 37986 5 1 1 37985
0 37987 7 1 2 100937 37986
0 37988 5 1 1 37987
0 37989 7 1 2 76505 97039
0 37990 5 1 1 37989
0 37991 7 1 2 37988 37990
0 37992 5 1 1 37991
0 37993 7 1 2 70412 37992
0 37994 5 1 1 37993
0 37995 7 1 2 63609 89305
0 37996 5 1 1 37995
0 37997 7 1 2 74696 37996
0 37998 5 2 1 37997
0 37999 7 1 2 65814 101004
0 38000 5 1 1 37999
0 38001 7 1 2 18939 38000
0 38002 5 1 1 38001
0 38003 7 1 2 67288 38002
0 38004 5 1 1 38003
0 38005 7 1 2 68450 72759
0 38006 5 1 1 38005
0 38007 7 1 2 38004 38006
0 38008 5 1 1 38007
0 38009 7 1 2 68688 38008
0 38010 5 1 1 38009
0 38011 7 1 2 74039 85586
0 38012 5 1 1 38011
0 38013 7 1 2 38010 38012
0 38014 5 1 1 38013
0 38015 7 1 2 88674 38014
0 38016 5 1 1 38015
0 38017 7 1 2 90934 100818
0 38018 5 1 1 38017
0 38019 7 1 2 83419 71542
0 38020 7 1 2 91117 38019
0 38021 5 1 1 38020
0 38022 7 1 2 38018 38021
0 38023 5 1 1 38022
0 38024 7 1 2 67496 38023
0 38025 5 1 1 38024
0 38026 7 2 2 63379 72833
0 38027 7 1 2 91575 101006
0 38028 5 1 1 38027
0 38029 7 1 2 73265 75186
0 38030 7 1 2 81593 38029
0 38031 5 1 1 38030
0 38032 7 1 2 38028 38031
0 38033 7 1 2 38025 38032
0 38034 5 1 1 38033
0 38035 7 1 2 66021 38034
0 38036 5 1 1 38035
0 38037 7 1 2 72760 81594
0 38038 5 1 1 38037
0 38039 7 1 2 80524 15130
0 38040 5 1 1 38039
0 38041 7 1 2 79911 83420
0 38042 7 1 2 38040 38041
0 38043 5 1 1 38042
0 38044 7 1 2 38038 38043
0 38045 5 1 1 38044
0 38046 7 1 2 68689 38045
0 38047 5 1 1 38046
0 38048 7 1 2 84854 88079
0 38049 5 1 1 38048
0 38050 7 1 2 89698 38049
0 38051 5 1 1 38050
0 38052 7 1 2 71543 38051
0 38053 5 1 1 38052
0 38054 7 1 2 38047 38053
0 38055 7 1 2 38036 38054
0 38056 5 1 1 38055
0 38057 7 1 2 67018 38056
0 38058 5 1 1 38057
0 38059 7 1 2 38016 38058
0 38060 5 1 1 38059
0 38061 7 1 2 65489 38060
0 38062 5 1 1 38061
0 38063 7 1 2 95706 98267
0 38064 5 1 1 38063
0 38065 7 1 2 88798 73221
0 38066 5 1 1 38065
0 38067 7 1 2 38064 38066
0 38068 5 1 1 38067
0 38069 7 1 2 74334 38068
0 38070 5 1 1 38069
0 38071 7 1 2 38062 38070
0 38072 5 1 1 38071
0 38073 7 1 2 96621 38072
0 38074 5 1 1 38073
0 38075 7 1 2 37994 38074
0 38076 5 1 1 38075
0 38077 7 1 2 96959 38076
0 38078 5 1 1 38077
0 38079 7 1 2 37960 38078
0 38080 5 1 1 38079
0 38081 7 1 2 81934 38080
0 38082 5 1 1 38081
0 38083 7 1 2 72174 96960
0 38084 5 1 1 38083
0 38085 7 3 2 72708 72338
0 38086 7 1 2 97312 101008
0 38087 5 1 1 38086
0 38088 7 1 2 38084 38087
0 38089 5 1 1 38088
0 38090 7 1 2 96608 38089
0 38091 5 1 1 38090
0 38092 7 1 2 72175 86252
0 38093 5 1 1 38092
0 38094 7 1 2 100418 38093
0 38095 5 1 1 38094
0 38096 7 1 2 99443 38095
0 38097 5 1 1 38096
0 38098 7 1 2 38091 38097
0 38099 5 1 1 38098
0 38100 7 1 2 96183 38099
0 38101 5 1 1 38100
0 38102 7 1 2 89847 97088
0 38103 5 1 1 38102
0 38104 7 2 2 70413 82994
0 38105 7 2 2 92174 97631
0 38106 7 1 2 87540 101013
0 38107 7 1 2 101011 38106
0 38108 7 1 2 38103 38107
0 38109 5 1 1 38108
0 38110 7 1 2 38101 38109
0 38111 5 1 1 38110
0 38112 7 1 2 65815 38111
0 38113 5 1 1 38112
0 38114 7 2 2 77947 95860
0 38115 5 2 1 101015
0 38116 7 1 2 67497 95486
0 38117 5 1 1 38116
0 38118 7 1 2 94478 38117
0 38119 5 1 1 38118
0 38120 7 1 2 70743 38119
0 38121 5 1 1 38120
0 38122 7 1 2 101017 38121
0 38123 5 1 1 38122
0 38124 7 2 2 74816 99326
0 38125 5 1 1 101019
0 38126 7 1 2 96178 101020
0 38127 7 1 2 38123 38126
0 38128 5 1 1 38127
0 38129 7 1 2 86795 98522
0 38130 5 1 1 38129
0 38131 7 3 2 67808 69021
0 38132 7 2 2 98140 101021
0 38133 7 1 2 91045 101024
0 38134 7 1 2 99540 38133
0 38135 5 1 1 38134
0 38136 7 1 2 38130 38135
0 38137 5 1 1 38136
0 38138 7 1 2 71976 96184
0 38139 7 1 2 38137 38138
0 38140 5 1 1 38139
0 38141 7 1 2 38128 38140
0 38142 5 1 1 38141
0 38143 7 1 2 68451 38142
0 38144 5 1 1 38143
0 38145 7 1 2 38113 38144
0 38146 5 1 1 38145
0 38147 7 1 2 68213 38146
0 38148 5 1 1 38147
0 38149 7 1 2 85948 37160
0 38150 5 2 1 38149
0 38151 7 1 2 73338 101026
0 38152 5 2 1 38151
0 38153 7 1 2 74727 7687
0 38154 5 1 1 38153
0 38155 7 1 2 71347 38154
0 38156 5 1 1 38155
0 38157 7 1 2 101028 38156
0 38158 5 1 1 38157
0 38159 7 1 2 78892 38158
0 38160 5 1 1 38159
0 38161 7 1 2 77821 80101
0 38162 7 1 2 97253 38161
0 38163 5 1 1 38162
0 38164 7 1 2 38160 38163
0 38165 5 1 1 38164
0 38166 7 1 2 100983 38165
0 38167 5 1 1 38166
0 38168 7 2 2 68032 80190
0 38169 5 1 1 101030
0 38170 7 1 2 80422 101031
0 38171 5 1 1 38170
0 38172 7 1 2 63193 92105
0 38173 5 1 1 38172
0 38174 7 1 2 38171 38173
0 38175 5 1 1 38174
0 38176 7 1 2 62613 38175
0 38177 5 1 1 38176
0 38178 7 1 2 78934 93543
0 38179 5 1 1 38178
0 38180 7 1 2 38177 38179
0 38181 5 1 1 38180
0 38182 7 1 2 86528 98523
0 38183 7 1 2 38181 38182
0 38184 5 1 1 38183
0 38185 7 1 2 38167 38184
0 38186 5 1 1 38185
0 38187 7 1 2 96514 38186
0 38188 5 1 1 38187
0 38189 7 1 2 38148 38188
0 38190 5 1 1 38189
0 38191 7 1 2 62176 38190
0 38192 5 1 1 38191
0 38193 7 1 2 33375 33380
0 38194 5 7 1 38193
0 38195 7 1 2 101032 101009
0 38196 5 1 1 38195
0 38197 7 3 2 97648 98576
0 38198 7 1 2 95658 101039
0 38199 5 1 1 38198
0 38200 7 1 2 38196 38199
0 38201 5 1 1 38200
0 38202 7 1 2 71977 38201
0 38203 5 1 1 38202
0 38204 7 2 2 63830 98038
0 38205 7 1 2 99375 101042
0 38206 5 1 1 38205
0 38207 7 1 2 74817 96961
0 38208 5 1 1 38207
0 38209 7 1 2 38206 38208
0 38210 5 1 1 38209
0 38211 7 1 2 101010 38210
0 38212 5 1 1 38211
0 38213 7 1 2 38203 38212
0 38214 5 1 1 38213
0 38215 7 1 2 63610 38214
0 38216 5 1 1 38215
0 38217 7 3 2 96948 98846
0 38218 7 1 2 76651 90143
0 38219 5 1 1 38218
0 38220 7 1 2 85631 92446
0 38221 5 1 1 38220
0 38222 7 1 2 38219 38221
0 38223 5 1 1 38222
0 38224 7 1 2 67019 38223
0 38225 5 1 1 38224
0 38226 7 1 2 74940 101016
0 38227 5 1 1 38226
0 38228 7 1 2 38225 38227
0 38229 5 1 1 38228
0 38230 7 1 2 101044 38229
0 38231 5 1 1 38230
0 38232 7 4 2 73339 100407
0 38233 5 1 1 101047
0 38234 7 1 2 79649 96962
0 38235 5 1 1 38234
0 38236 7 2 2 94214 97632
0 38237 7 1 2 99368 101051
0 38238 5 1 1 38237
0 38239 7 1 2 38235 38238
0 38240 5 1 1 38239
0 38241 7 1 2 101048 38240
0 38242 5 1 1 38241
0 38243 7 1 2 38231 38242
0 38244 7 1 2 38216 38243
0 38245 5 1 1 38244
0 38246 7 1 2 68214 38245
0 38247 5 1 1 38246
0 38248 7 4 2 93052 97633
0 38249 7 1 2 84338 95623
0 38250 7 1 2 101053 38249
0 38251 5 1 1 38250
0 38252 7 1 2 75001 98524
0 38253 7 1 2 86788 38252
0 38254 5 1 1 38253
0 38255 7 1 2 38251 38254
0 38256 5 1 1 38255
0 38257 7 1 2 96892 38256
0 38258 5 1 1 38257
0 38259 7 1 2 38247 38258
0 38260 5 1 1 38259
0 38261 7 1 2 65816 38260
0 38262 5 1 1 38261
0 38263 7 1 2 98533 38125
0 38264 5 1 1 38263
0 38265 7 1 2 71978 83421
0 38266 7 1 2 38264 38265
0 38267 5 1 1 38266
0 38268 7 1 2 75198 81595
0 38269 7 1 2 97313 38268
0 38270 5 1 1 38269
0 38271 7 1 2 38267 38270
0 38272 5 1 1 38271
0 38273 7 1 2 94570 38272
0 38274 5 1 1 38273
0 38275 7 3 2 74818 83422
0 38276 5 5 1 101057
0 38277 7 1 2 73899 89724
0 38278 5 1 1 38277
0 38279 7 1 2 101060 38278
0 38280 5 2 1 38279
0 38281 7 1 2 71256 101065
0 38282 5 1 1 38281
0 38283 7 1 2 70744 88799
0 38284 5 1 1 38283
0 38285 7 1 2 101061 38284
0 38286 5 2 1 38285
0 38287 7 1 2 85840 101067
0 38288 5 1 1 38287
0 38289 7 1 2 85232 95756
0 38290 5 1 1 38289
0 38291 7 1 2 38288 38290
0 38292 7 1 2 38282 38291
0 38293 5 1 1 38292
0 38294 7 1 2 96963 38293
0 38295 5 1 1 38294
0 38296 7 1 2 38274 38295
0 38297 5 1 1 38296
0 38298 7 1 2 65490 38297
0 38299 5 1 1 38298
0 38300 7 2 2 92996 98141
0 38301 7 2 2 74084 101069
0 38302 7 1 2 89972 83200
0 38303 7 1 2 101071 38302
0 38304 5 1 1 38303
0 38305 7 2 2 74040 96964
0 38306 5 1 1 101073
0 38307 7 1 2 62431 101074
0 38308 5 1 1 38307
0 38309 7 1 2 38304 38308
0 38310 5 1 1 38309
0 38311 7 1 2 97816 38310
0 38312 5 1 1 38311
0 38313 7 1 2 38299 38312
0 38314 5 1 1 38313
0 38315 7 1 2 67020 38314
0 38316 5 1 1 38315
0 38317 7 2 2 71979 86110
0 38318 7 3 2 64288 93173
0 38319 7 1 2 84261 101077
0 38320 7 1 2 99561 38319
0 38321 7 1 2 101075 38320
0 38322 5 1 1 38321
0 38323 7 1 2 38316 38322
0 38324 7 1 2 38262 38323
0 38325 5 1 1 38324
0 38326 7 1 2 69603 38325
0 38327 5 1 1 38326
0 38328 7 1 2 63831 98973
0 38329 7 1 2 99296 38328
0 38330 7 1 2 100146 38329
0 38331 5 1 1 38330
0 38332 7 1 2 38327 38331
0 38333 5 1 1 38332
0 38334 7 1 2 96144 38333
0 38335 5 1 1 38334
0 38336 7 1 2 38192 38335
0 38337 5 1 1 38336
0 38338 7 1 2 61632 38337
0 38339 5 1 1 38338
0 38340 7 1 2 89699 101062
0 38341 5 1 1 38340
0 38342 7 1 2 67021 38341
0 38343 5 1 1 38342
0 38344 7 1 2 68215 95085
0 38345 5 1 1 38344
0 38346 7 1 2 38343 38345
0 38347 5 1 1 38346
0 38348 7 1 2 72834 38347
0 38349 5 1 1 38348
0 38350 7 1 2 67289 88675
0 38351 7 1 2 84729 38350
0 38352 5 1 1 38351
0 38353 7 1 2 38349 38352
0 38354 5 1 1 38353
0 38355 7 1 2 66022 38354
0 38356 5 1 1 38355
0 38357 7 1 2 82141 73730
0 38358 7 1 2 82071 38357
0 38359 5 1 1 38358
0 38360 7 1 2 38356 38359
0 38361 5 1 1 38360
0 38362 7 1 2 76716 38361
0 38363 5 1 1 38362
0 38364 7 1 2 80285 79830
0 38365 7 2 2 79230 38364
0 38366 5 1 1 101080
0 38367 7 1 2 68216 101081
0 38368 5 1 1 38367
0 38369 7 1 2 38363 38368
0 38370 5 1 1 38369
0 38371 7 1 2 88999 93863
0 38372 7 1 2 38370 38371
0 38373 5 1 1 38372
0 38374 7 1 2 70414 94824
0 38375 7 1 2 87439 38374
0 38376 7 1 2 100357 38375
0 38377 7 1 2 100468 38376
0 38378 5 1 1 38377
0 38379 7 1 2 38373 38378
0 38380 5 1 1 38379
0 38381 7 1 2 98208 38380
0 38382 5 1 1 38381
0 38383 7 1 2 74849 92517
0 38384 5 2 1 38383
0 38385 7 1 2 83423 101082
0 38386 5 1 1 38385
0 38387 7 1 2 98285 38386
0 38388 5 1 1 38387
0 38389 7 1 2 86210 38388
0 38390 5 1 1 38389
0 38391 7 1 2 73950 101066
0 38392 5 1 1 38391
0 38393 7 1 2 72176 101068
0 38394 5 1 1 38393
0 38395 7 1 2 38392 38394
0 38396 5 1 1 38395
0 38397 7 1 2 65491 38396
0 38398 5 1 1 38397
0 38399 7 1 2 38390 38398
0 38400 5 1 1 38399
0 38401 7 1 2 96209 101040
0 38402 7 1 2 38400 38401
0 38403 5 1 1 38402
0 38404 7 1 2 64380 38403
0 38405 7 1 2 38382 38404
0 38406 5 1 1 38405
0 38407 7 2 2 74819 96893
0 38408 5 1 1 101084
0 38409 7 1 2 93153 99692
0 38410 7 1 2 97194 38409
0 38411 7 1 2 101085 38410
0 38412 5 1 1 38411
0 38413 7 1 2 65492 95089
0 38414 5 1 1 38413
0 38415 7 1 2 95420 38414
0 38416 5 1 1 38415
0 38417 7 1 2 68217 38416
0 38418 5 1 1 38417
0 38419 7 1 2 89619 86193
0 38420 5 1 1 38419
0 38421 7 1 2 38418 38420
0 38422 5 1 1 38421
0 38423 7 1 2 81474 82444
0 38424 7 1 2 93864 38423
0 38425 7 1 2 38422 38424
0 38426 5 1 1 38425
0 38427 7 1 2 38412 38426
0 38428 5 1 1 38427
0 38429 7 1 2 72177 38428
0 38430 5 1 1 38429
0 38431 7 3 2 74187 93865
0 38432 7 2 2 68218 86043
0 38433 7 1 2 74584 96210
0 38434 7 1 2 101089 38433
0 38435 7 1 2 101086 38434
0 38436 5 1 1 38435
0 38437 7 1 2 67809 96213
0 38438 5 1 1 38437
0 38439 7 1 2 82995 93154
0 38440 5 1 1 38439
0 38441 7 1 2 38438 38440
0 38442 5 1 1 38441
0 38443 7 1 2 61308 38442
0 38444 5 1 1 38443
0 38445 7 1 2 66141 93174
0 38446 7 1 2 96211 38445
0 38447 5 1 1 38446
0 38448 7 1 2 38444 38447
0 38449 5 1 1 38448
0 38450 7 1 2 94278 99362
0 38451 7 1 2 38449 38450
0 38452 5 1 1 38451
0 38453 7 1 2 38436 38452
0 38454 5 1 1 38453
0 38455 7 1 2 67290 38454
0 38456 5 1 1 38455
0 38457 7 2 2 80191 100735
0 38458 7 1 2 91775 101091
0 38459 7 1 2 101087 38458
0 38460 5 1 1 38459
0 38461 7 1 2 38456 38460
0 38462 5 1 1 38461
0 38463 7 1 2 67022 38462
0 38464 5 1 1 38463
0 38465 7 1 2 38430 38464
0 38466 5 1 1 38465
0 38467 7 1 2 64289 38466
0 38468 5 1 1 38467
0 38469 7 1 2 80036 99076
0 38470 7 1 2 75041 38469
0 38471 7 2 2 77822 88102
0 38472 7 1 2 98925 101093
0 38473 7 1 2 38470 38472
0 38474 5 1 1 38473
0 38475 7 1 2 69242 38474
0 38476 7 1 2 38468 38475
0 38477 5 1 1 38476
0 38478 7 1 2 61633 38477
0 38479 7 1 2 38406 38478
0 38480 5 1 1 38479
0 38481 7 1 2 75121 83623
0 38482 5 1 1 38481
0 38483 7 1 2 68219 7949
0 38484 7 1 2 38482 38483
0 38485 5 1 1 38484
0 38486 7 1 2 38408 38485
0 38487 5 1 1 38486
0 38488 7 1 2 93728 38487
0 38489 5 1 1 38488
0 38490 7 1 2 78957 101058
0 38491 5 1 1 38490
0 38492 7 1 2 83500 100978
0 38493 5 1 1 38492
0 38494 7 1 2 38491 38493
0 38495 5 1 1 38494
0 38496 7 1 2 67023 38495
0 38497 5 1 1 38496
0 38498 7 1 2 64773 75114
0 38499 7 1 2 100979 38498
0 38500 5 1 1 38499
0 38501 7 1 2 38497 38500
0 38502 5 1 1 38501
0 38503 7 1 2 72178 38502
0 38504 5 1 1 38503
0 38505 7 1 2 84714 80108
0 38506 7 1 2 95090 38505
0 38507 5 1 1 38506
0 38508 7 1 2 38504 38507
0 38509 5 1 1 38508
0 38510 7 1 2 67715 38509
0 38511 5 1 1 38510
0 38512 7 1 2 38489 38511
0 38513 5 1 1 38512
0 38514 7 1 2 99419 100828
0 38515 7 1 2 38513 38514
0 38516 5 1 1 38515
0 38517 7 1 2 84865 84543
0 38518 7 1 2 98338 38517
0 38519 7 1 2 78958 94669
0 38520 7 1 2 38518 38519
0 38521 7 1 2 94531 38520
0 38522 5 1 1 38521
0 38523 7 1 2 38516 38522
0 38524 5 1 1 38523
0 38525 7 1 2 65493 94717
0 38526 7 1 2 38524 38525
0 38527 5 1 1 38526
0 38528 7 1 2 38480 38527
0 38529 5 1 1 38528
0 38530 7 1 2 73480 38529
0 38531 5 1 1 38530
0 38532 7 1 2 38339 38531
0 38533 7 1 2 38082 38532
0 38534 5 1 1 38533
0 38535 7 1 2 65189 38534
0 38536 5 1 1 38535
0 38537 7 1 2 97093 98363
0 38538 5 1 1 38537
0 38539 7 1 2 65817 92400
0 38540 7 1 2 87440 38539
0 38541 5 1 1 38540
0 38542 7 1 2 38538 38541
0 38543 5 1 1 38542
0 38544 7 1 2 75306 94750
0 38545 7 1 2 38543 38544
0 38546 5 1 1 38545
0 38547 7 1 2 76535 94751
0 38548 7 1 2 83722 38547
0 38549 5 1 1 38548
0 38550 7 1 2 78180 88125
0 38551 7 1 2 95630 97288
0 38552 7 1 2 38550 38551
0 38553 5 1 1 38552
0 38554 7 1 2 38549 38553
0 38555 5 1 1 38554
0 38556 7 1 2 72179 38555
0 38557 5 1 1 38556
0 38558 7 1 2 80501 90401
0 38559 7 1 2 92449 94752
0 38560 7 1 2 38558 38559
0 38561 5 1 1 38560
0 38562 7 1 2 90322 78009
0 38563 7 1 2 91608 95631
0 38564 7 1 2 38562 38563
0 38565 5 1 1 38564
0 38566 7 1 2 38561 38565
0 38567 5 1 1 38566
0 38568 7 1 2 67024 38567
0 38569 5 1 1 38568
0 38570 7 1 2 38557 38569
0 38571 7 1 2 38546 38570
0 38572 5 1 1 38571
0 38573 7 1 2 63380 38572
0 38574 5 1 1 38573
0 38575 7 1 2 80013 96256
0 38576 5 1 1 38575
0 38577 7 1 2 76389 82187
0 38578 7 1 2 15632 38577
0 38579 5 1 1 38578
0 38580 7 1 2 38576 38579
0 38581 5 1 1 38580
0 38582 7 1 2 77528 38581
0 38583 5 1 1 38582
0 38584 7 1 2 73778 75455
0 38585 7 1 2 89875 38584
0 38586 5 1 1 38585
0 38587 7 1 2 74085 85557
0 38588 7 1 2 98349 38587
0 38589 5 1 1 38588
0 38590 7 1 2 38586 38589
0 38591 7 1 2 38583 38590
0 38592 5 1 1 38591
0 38593 7 1 2 83387 95117
0 38594 7 1 2 38592 38593
0 38595 5 1 1 38594
0 38596 7 1 2 38574 38595
0 38597 5 1 1 38596
0 38598 7 1 2 65190 38597
0 38599 5 1 1 38598
0 38600 7 1 2 62881 91495
0 38601 5 1 1 38600
0 38602 7 1 2 84964 38601
0 38603 5 1 1 38602
0 38604 7 1 2 71854 38603
0 38605 5 1 1 38604
0 38606 7 1 2 70950 78388
0 38607 5 1 1 38606
0 38608 7 1 2 38605 38607
0 38609 5 1 1 38608
0 38610 7 1 2 78030 38609
0 38611 5 1 1 38610
0 38612 7 1 2 19146 38611
0 38613 5 1 1 38612
0 38614 7 1 2 65818 38613
0 38615 5 1 1 38614
0 38616 7 3 2 67498 74662
0 38617 5 1 1 101095
0 38618 7 1 2 93656 38617
0 38619 5 1 1 38618
0 38620 7 1 2 81167 38619
0 38621 5 1 1 38620
0 38622 7 1 2 38615 38621
0 38623 5 1 1 38622
0 38624 7 1 2 84125 94681
0 38625 7 1 2 38623 38624
0 38626 5 1 1 38625
0 38627 7 2 2 65494 94532
0 38628 5 2 1 101098
0 38629 7 1 2 91959 94856
0 38630 7 1 2 101099 38629
0 38631 5 1 1 38630
0 38632 7 1 2 38626 38631
0 38633 5 1 1 38632
0 38634 7 1 2 77377 38633
0 38635 5 1 1 38634
0 38636 7 1 2 38599 38635
0 38637 5 1 1 38636
0 38638 7 1 2 93866 38637
0 38639 5 1 1 38638
0 38640 7 1 2 82975 93568
0 38641 5 1 1 38640
0 38642 7 1 2 77924 94090
0 38643 5 1 1 38642
0 38644 7 1 2 71855 78091
0 38645 7 1 2 5893 38644
0 38646 5 1 1 38645
0 38647 7 1 2 38643 38646
0 38648 7 1 2 38641 38647
0 38649 5 1 1 38648
0 38650 7 1 2 70415 38649
0 38651 5 1 1 38650
0 38652 7 1 2 79664 95392
0 38653 5 1 1 38652
0 38654 7 1 2 38651 38653
0 38655 5 1 1 38654
0 38656 7 1 2 97160 38655
0 38657 5 1 1 38656
0 38658 7 1 2 79957 92536
0 38659 7 1 2 93969 96731
0 38660 7 1 2 38658 38659
0 38661 5 1 1 38660
0 38662 7 1 2 38657 38661
0 38663 5 1 1 38662
0 38664 7 1 2 96965 38663
0 38665 5 1 1 38664
0 38666 7 1 2 72293 99317
0 38667 7 2 2 72709 74682
0 38668 5 1 1 101102
0 38669 7 2 2 81713 98039
0 38670 7 1 2 96084 101104
0 38671 7 1 2 101103 38670
0 38672 7 1 2 38666 38671
0 38673 5 1 1 38672
0 38674 7 1 2 38665 38673
0 38675 5 1 1 38674
0 38676 7 1 2 63381 38675
0 38677 5 1 1 38676
0 38678 7 1 2 72835 78825
0 38679 7 1 2 93086 97716
0 38680 7 1 2 38678 38679
0 38681 7 1 2 91850 38680
0 38682 7 1 2 86789 38681
0 38683 5 1 1 38682
0 38684 7 3 2 73340 97584
0 38685 7 1 2 75307 96085
0 38686 7 1 2 101106 38685
0 38687 7 1 2 101052 38686
0 38688 5 1 1 38687
0 38689 7 1 2 38683 38688
0 38690 5 1 1 38689
0 38691 7 1 2 63382 38690
0 38692 5 1 1 38691
0 38693 7 1 2 85272 82978
0 38694 5 1 1 38693
0 38695 7 1 2 89355 100959
0 38696 5 1 1 38695
0 38697 7 1 2 71980 38696
0 38698 5 1 1 38697
0 38699 7 1 2 38694 38698
0 38700 5 1 1 38699
0 38701 7 1 2 72854 38700
0 38702 5 1 1 38701
0 38703 7 1 2 88264 85804
0 38704 5 1 1 38703
0 38705 7 1 2 38702 38704
0 38706 5 1 1 38705
0 38707 7 1 2 96521 98525
0 38708 7 1 2 38706 38707
0 38709 5 1 1 38708
0 38710 7 1 2 38692 38709
0 38711 5 1 1 38710
0 38712 7 1 2 66023 38711
0 38713 5 1 1 38712
0 38714 7 1 2 81308 86790
0 38715 5 1 1 38714
0 38716 7 1 2 83549 96410
0 38717 5 1 1 38716
0 38718 7 1 2 38715 38717
0 38719 5 1 1 38718
0 38720 7 1 2 68452 38719
0 38721 5 1 1 38720
0 38722 7 1 2 71257 97817
0 38723 7 1 2 79029 38722
0 38724 5 1 1 38723
0 38725 7 1 2 38721 38724
0 38726 5 1 1 38725
0 38727 7 1 2 87020 97649
0 38728 7 1 2 99693 38727
0 38729 7 1 2 91851 38728
0 38730 7 1 2 38726 38729
0 38731 5 1 1 38730
0 38732 7 1 2 38713 38731
0 38733 5 1 1 38732
0 38734 7 1 2 65819 38733
0 38735 5 1 1 38734
0 38736 7 2 2 79609 93569
0 38737 7 1 2 76536 98526
0 38738 7 1 2 100643 38737
0 38739 7 1 2 101109 38738
0 38740 5 1 1 38739
0 38741 7 1 2 38735 38740
0 38742 7 1 2 38677 38741
0 38743 7 1 2 38639 38742
0 38744 5 1 1 38743
0 38745 7 1 2 76175 38744
0 38746 5 1 1 38745
0 38747 7 1 2 7531 94189
0 38748 5 4 1 38747
0 38749 7 3 2 75729 101111
0 38750 5 2 1 101115
0 38751 7 1 2 70951 101116
0 38752 5 1 1 38751
0 38753 7 1 2 76329 73691
0 38754 7 1 2 92136 38753
0 38755 5 1 1 38754
0 38756 7 1 2 38752 38755
0 38757 5 1 1 38756
0 38758 7 1 2 70416 38757
0 38759 5 1 1 38758
0 38760 7 1 2 86577 97094
0 38761 7 1 2 82694 38760
0 38762 5 1 1 38761
0 38763 7 1 2 38759 38762
0 38764 5 1 1 38763
0 38765 7 1 2 64164 38764
0 38766 5 1 1 38765
0 38767 7 2 2 71130 77823
0 38768 5 1 1 101120
0 38769 7 1 2 86565 101121
0 38770 5 1 1 38769
0 38771 7 1 2 65495 38768
0 38772 5 1 1 38771
0 38773 7 1 2 71856 74714
0 38774 7 1 2 38772 38773
0 38775 5 1 1 38774
0 38776 7 1 2 38770 38775
0 38777 5 1 1 38776
0 38778 7 1 2 63383 38777
0 38779 5 1 1 38778
0 38780 7 1 2 38766 38779
0 38781 5 1 1 38780
0 38782 7 1 2 62177 38781
0 38783 5 1 1 38782
0 38784 7 2 2 85815 85632
0 38785 5 2 1 101122
0 38786 7 2 2 70417 101123
0 38787 5 1 1 101126
0 38788 7 2 2 74585 89902
0 38789 7 1 2 100408 101128
0 38790 5 1 1 38789
0 38791 7 1 2 38787 38790
0 38792 5 1 1 38791
0 38793 7 1 2 65820 38792
0 38794 5 1 1 38793
0 38795 7 1 2 71740 84659
0 38796 5 1 1 38795
0 38797 7 1 2 62432 86486
0 38798 5 1 1 38797
0 38799 7 1 2 38796 38798
0 38800 5 1 1 38799
0 38801 7 1 2 85816 38800
0 38802 5 1 1 38801
0 38803 7 1 2 38794 38802
0 38804 5 1 1 38803
0 38805 7 1 2 81639 38804
0 38806 5 1 1 38805
0 38807 7 1 2 38783 38806
0 38808 5 1 1 38807
0 38809 7 1 2 96145 38808
0 38810 5 1 1 38809
0 38811 7 1 2 62178 96524
0 38812 5 1 1 38811
0 38813 7 1 2 3776 38812
0 38814 5 1 1 38813
0 38815 7 1 2 90966 38814
0 38816 5 1 1 38815
0 38817 7 1 2 65496 38816
0 38818 5 1 1 38817
0 38819 7 1 2 82415 85714
0 38820 7 1 2 88699 38819
0 38821 7 1 2 96817 38820
0 38822 5 1 1 38821
0 38823 7 1 2 89533 86273
0 38824 5 2 1 38823
0 38825 7 1 2 90970 101130
0 38826 5 1 1 38825
0 38827 7 1 2 70418 38826
0 38828 7 1 2 38822 38827
0 38829 5 1 1 38828
0 38830 7 1 2 65821 38829
0 38831 7 1 2 38818 38830
0 38832 5 1 1 38831
0 38833 7 1 2 85656 93626
0 38834 7 1 2 87868 38833
0 38835 7 1 2 93081 38834
0 38836 5 1 1 38835
0 38837 7 1 2 38832 38836
0 38838 5 1 1 38837
0 38839 7 1 2 72180 38838
0 38840 5 1 1 38839
0 38841 7 2 2 88748 86184
0 38842 7 2 2 87497 96680
0 38843 7 1 2 101134 100863
0 38844 7 1 2 101132 38843
0 38845 5 1 1 38844
0 38846 7 1 2 38840 38845
0 38847 7 1 2 38810 38846
0 38848 5 1 1 38847
0 38849 7 1 2 61634 38848
0 38850 5 1 1 38849
0 38851 7 1 2 88590 90967
0 38852 7 1 2 92514 38851
0 38853 5 1 1 38852
0 38854 7 1 2 87406 96240
0 38855 5 1 1 38854
0 38856 7 1 2 96595 38855
0 38857 5 1 1 38856
0 38858 7 1 2 77631 101112
0 38859 7 1 2 38857 38858
0 38860 5 1 1 38859
0 38861 7 1 2 38853 38860
0 38862 5 1 1 38861
0 38863 7 1 2 62179 38862
0 38864 5 1 1 38863
0 38865 7 1 2 87665 96610
0 38866 5 1 1 38865
0 38867 7 1 2 38864 38866
0 38868 5 1 1 38867
0 38869 7 1 2 78333 38868
0 38870 5 1 1 38869
0 38871 7 2 2 71981 72883
0 38872 7 1 2 81640 101136
0 38873 5 1 1 38872
0 38874 7 1 2 84304 101117
0 38875 5 1 1 38874
0 38876 7 1 2 38873 38875
0 38877 5 1 1 38876
0 38878 7 1 2 90802 96622
0 38879 7 1 2 38877 38878
0 38880 5 1 1 38879
0 38881 7 1 2 38870 38880
0 38882 7 1 2 38850 38881
0 38883 5 1 1 38882
0 38884 7 1 2 96966 38883
0 38885 5 1 1 38884
0 38886 7 1 2 97073 97868
0 38887 5 1 1 38886
0 38888 7 2 2 95052 96146
0 38889 7 1 2 91046 101138
0 38890 5 1 1 38889
0 38891 7 1 2 38887 38890
0 38892 5 1 1 38891
0 38893 7 1 2 67291 38892
0 38894 5 1 1 38893
0 38895 7 1 2 86483 101139
0 38896 5 1 1 38895
0 38897 7 1 2 38894 38896
0 38898 5 1 1 38897
0 38899 7 1 2 67716 38898
0 38900 5 1 1 38899
0 38901 7 1 2 77121 96777
0 38902 7 1 2 87544 38901
0 38903 5 1 1 38902
0 38904 7 1 2 38900 38903
0 38905 5 1 1 38904
0 38906 7 1 2 71258 38905
0 38907 5 1 1 38906
0 38908 7 1 2 72294 82930
0 38909 7 1 2 91586 97053
0 38910 7 1 2 38908 38909
0 38911 5 1 1 38910
0 38912 7 1 2 38907 38911
0 38913 5 1 1 38912
0 38914 7 1 2 86673 99327
0 38915 7 1 2 38913 38914
0 38916 5 1 1 38915
0 38917 7 1 2 38885 38916
0 38918 5 1 1 38917
0 38919 7 1 2 64774 38918
0 38920 5 1 1 38919
0 38921 7 1 2 91500 94857
0 38922 5 1 1 38921
0 38923 7 1 2 82921 94753
0 38924 5 1 1 38923
0 38925 7 1 2 38922 38924
0 38926 5 1 1 38925
0 38927 7 1 2 78314 38926
0 38928 5 1 1 38927
0 38929 7 2 2 87839 96822
0 38930 7 1 2 67292 81641
0 38931 7 1 2 95642 38930
0 38932 7 1 2 101140 38931
0 38933 5 1 1 38932
0 38934 7 1 2 38928 38933
0 38935 5 1 1 38934
0 38936 7 1 2 65497 38935
0 38937 5 1 1 38936
0 38938 7 1 2 74907 2792
0 38939 5 1 1 38938
0 38940 7 1 2 70952 82722
0 38941 7 1 2 95680 38940
0 38942 7 1 2 38939 38941
0 38943 5 1 1 38942
0 38944 7 1 2 38937 38943
0 38945 5 1 1 38944
0 38946 7 1 2 76176 38945
0 38947 5 1 1 38946
0 38948 7 1 2 89468 95263
0 38949 5 1 1 38948
0 38950 7 1 2 95635 38949
0 38951 5 1 1 38950
0 38952 7 1 2 69604 38951
0 38953 5 1 1 38952
0 38954 7 1 2 61635 94627
0 38955 5 1 1 38954
0 38956 7 1 2 38953 38955
0 38957 5 1 1 38956
0 38958 7 1 2 91678 92741
0 38959 7 1 2 38957 38958
0 38960 5 1 1 38959
0 38961 7 1 2 38947 38960
0 38962 5 1 1 38961
0 38963 7 1 2 62180 38962
0 38964 5 1 1 38963
0 38965 7 1 2 81775 78181
0 38966 7 1 2 86640 38965
0 38967 7 1 2 95095 38966
0 38968 5 1 1 38967
0 38969 7 1 2 38964 38968
0 38970 5 1 1 38969
0 38971 7 1 2 93867 38970
0 38972 5 1 1 38971
0 38973 7 2 2 97634 98620
0 38974 7 1 2 91063 101142
0 38975 5 1 1 38974
0 38976 7 1 2 73664 86495
0 38977 5 3 1 38976
0 38978 7 1 2 96967 101144
0 38979 5 1 1 38978
0 38980 7 1 2 38975 38979
0 38981 5 1 1 38980
0 38982 7 1 2 86976 38981
0 38983 5 1 1 38982
0 38984 7 3 2 69132 69605
0 38985 7 1 2 101022 101147
0 38986 7 1 2 84246 38985
0 38987 7 1 2 100630 38986
0 38988 5 1 1 38987
0 38989 7 1 2 38983 38988
0 38990 5 1 1 38989
0 38991 7 1 2 67717 38990
0 38992 5 1 1 38991
0 38993 7 1 2 88126 97717
0 38994 7 1 2 99226 38993
0 38995 7 1 2 77834 38994
0 38996 5 1 1 38995
0 38997 7 1 2 38992 38996
0 38998 5 1 1 38997
0 38999 7 1 2 97040 38998
0 39000 5 1 1 38999
0 39001 7 1 2 38972 39000
0 39002 5 1 1 39001
0 39003 7 1 2 73481 39002
0 39004 5 1 1 39003
0 39005 7 1 2 80746 96119
0 39006 7 1 2 88080 39005
0 39007 5 1 1 39006
0 39008 7 1 2 78762 92401
0 39009 7 1 2 86908 39008
0 39010 5 1 1 39009
0 39011 7 1 2 39007 39010
0 39012 5 1 1 39011
0 39013 7 1 2 61636 39012
0 39014 5 1 1 39013
0 39015 7 2 2 62433 89821
0 39016 5 1 1 101150
0 39017 7 1 2 83444 101151
0 39018 5 1 1 39017
0 39019 7 1 2 39014 39018
0 39020 5 1 1 39019
0 39021 7 1 2 93126 39020
0 39022 5 1 1 39021
0 39023 7 2 2 89563 93020
0 39024 7 1 2 81671 89652
0 39025 7 1 2 101152 39024
0 39026 5 1 1 39025
0 39027 7 1 2 39022 39026
0 39028 5 1 1 39027
0 39029 7 1 2 68690 39028
0 39030 5 1 1 39029
0 39031 7 1 2 72181 91963
0 39032 5 1 1 39031
0 39033 7 1 2 76055 79979
0 39034 5 1 1 39033
0 39035 7 1 2 39032 39034
0 39036 5 1 1 39035
0 39037 7 1 2 71259 93127
0 39038 7 1 2 90590 39037
0 39039 7 1 2 39036 39038
0 39040 5 1 1 39039
0 39041 7 1 2 39030 39040
0 39042 5 1 1 39041
0 39043 7 1 2 65822 39042
0 39044 5 1 1 39043
0 39045 7 1 2 90101 96541
0 39046 7 1 2 91919 39045
0 39047 7 1 2 89605 39046
0 39048 5 1 1 39047
0 39049 7 1 2 39044 39048
0 39050 5 1 1 39049
0 39051 7 2 2 90774 97989
0 39052 7 1 2 81714 101154
0 39053 7 1 2 39050 39052
0 39054 5 1 1 39053
0 39055 7 1 2 39004 39054
0 39056 7 1 2 38920 39055
0 39057 5 1 1 39056
0 39058 7 1 2 70116 39057
0 39059 5 1 1 39058
0 39060 7 1 2 38746 39059
0 39061 7 1 2 38536 39060
0 39062 7 1 2 37930 39061
0 39063 5 1 1 39062
0 39064 7 1 2 93803 39063
0 39065 5 1 1 39064
0 39066 7 1 2 73341 78447
0 39067 5 2 1 39066
0 39068 7 1 2 11648 101156
0 39069 5 1 1 39068
0 39070 7 1 2 68691 39069
0 39071 5 1 1 39070
0 39072 7 1 2 85096 39071
0 39073 5 1 1 39072
0 39074 7 1 2 76177 39073
0 39075 5 1 1 39074
0 39076 7 1 2 82222 91964
0 39077 5 1 1 39076
0 39078 7 1 2 39075 39077
0 39079 5 1 1 39078
0 39080 7 1 2 76896 39079
0 39081 5 1 1 39080
0 39082 7 1 2 90539 85982
0 39083 5 1 1 39082
0 39084 7 1 2 39081 39083
0 39085 5 1 1 39084
0 39086 7 1 2 69606 39085
0 39087 5 1 1 39086
0 39088 7 1 2 79755 90480
0 39089 7 1 2 92132 39088
0 39090 5 1 1 39089
0 39091 7 1 2 39087 39090
0 39092 5 1 1 39091
0 39093 7 1 2 64552 39092
0 39094 5 1 1 39093
0 39095 7 1 2 68692 92447
0 39096 5 1 1 39095
0 39097 7 1 2 94469 39096
0 39098 5 1 1 39097
0 39099 7 1 2 70117 39098
0 39100 5 1 1 39099
0 39101 7 2 2 65191 84607
0 39102 7 1 2 71857 101158
0 39103 5 1 1 39102
0 39104 7 1 2 39100 39103
0 39105 5 1 1 39104
0 39106 7 1 2 91468 39105
0 39107 5 1 1 39106
0 39108 7 1 2 39094 39107
0 39109 5 1 1 39108
0 39110 7 1 2 81642 39109
0 39111 5 1 1 39110
0 39112 7 1 2 86766 91170
0 39113 7 1 2 88701 39112
0 39114 5 1 1 39113
0 39115 7 1 2 63194 93443
0 39116 5 1 1 39115
0 39117 7 1 2 88418 95029
0 39118 5 1 1 39117
0 39119 7 1 2 39116 39118
0 39120 5 1 1 39119
0 39121 7 1 2 83652 87096
0 39122 7 1 2 39120 39121
0 39123 5 1 1 39122
0 39124 7 1 2 39114 39123
0 39125 5 1 1 39124
0 39126 7 1 2 71348 39125
0 39127 5 1 1 39126
0 39128 7 1 2 91141 83846
0 39129 5 1 1 39128
0 39130 7 1 2 85430 91937
0 39131 5 1 1 39130
0 39132 7 1 2 39129 39131
0 39133 5 1 1 39132
0 39134 7 1 2 82430 39133
0 39135 5 1 1 39134
0 39136 7 1 2 39127 39135
0 39137 7 1 2 39111 39136
0 39138 5 1 1 39137
0 39139 7 1 2 62181 39138
0 39140 5 1 1 39139
0 39141 7 1 2 74683 90775
0 39142 7 1 2 100855 39141
0 39143 5 1 1 39142
0 39144 7 1 2 74055 96007
0 39145 5 1 1 39144
0 39146 7 1 2 70419 81265
0 39147 7 1 2 39145 39146
0 39148 5 1 1 39147
0 39149 7 1 2 39143 39148
0 39150 5 1 1 39149
0 39151 7 1 2 86455 39150
0 39152 5 1 1 39151
0 39153 7 3 2 89169 90776
0 39154 7 1 2 67499 81743
0 39155 7 1 2 82825 39154
0 39156 7 1 2 101160 39155
0 39157 5 1 1 39156
0 39158 7 1 2 39152 39157
0 39159 5 1 1 39158
0 39160 7 1 2 84231 39159
0 39161 5 1 1 39160
0 39162 7 2 2 77603 76211
0 39163 5 1 1 101163
0 39164 7 1 2 78391 39163
0 39165 5 1 1 39164
0 39166 7 1 2 62434 39165
0 39167 5 1 1 39166
0 39168 7 1 2 95595 39167
0 39169 5 1 1 39168
0 39170 7 1 2 86456 39169
0 39171 5 1 1 39170
0 39172 7 1 2 74959 98234
0 39173 5 1 1 39172
0 39174 7 1 2 39171 39173
0 39175 5 1 1 39174
0 39176 7 1 2 83263 39175
0 39177 5 1 1 39176
0 39178 7 1 2 94091 94249
0 39179 5 1 1 39178
0 39180 7 1 2 62882 85558
0 39181 7 1 2 94215 39180
0 39182 5 1 1 39181
0 39183 7 1 2 39179 39182
0 39184 5 1 1 39183
0 39185 7 1 2 88454 39184
0 39186 5 1 1 39185
0 39187 7 1 2 39177 39186
0 39188 7 1 2 39161 39187
0 39189 5 1 1 39188
0 39190 7 1 2 78826 39189
0 39191 5 1 1 39190
0 39192 7 1 2 39140 39191
0 39193 5 1 1 39192
0 39194 7 1 2 69022 39193
0 39195 5 1 1 39194
0 39196 7 1 2 90777 80215
0 39197 5 1 1 39196
0 39198 7 1 2 88368 91636
0 39199 5 1 1 39198
0 39200 7 1 2 39197 39199
0 39201 5 1 1 39200
0 39202 7 1 2 66525 39201
0 39203 5 1 1 39202
0 39204 7 1 2 82590 93414
0 39205 5 1 1 39204
0 39206 7 1 2 39203 39205
0 39207 5 1 1 39206
0 39208 7 1 2 90834 39207
0 39209 5 1 1 39208
0 39210 7 3 2 65498 89266
0 39211 7 1 2 76742 92524
0 39212 7 1 2 101165 39211
0 39213 5 1 1 39212
0 39214 7 1 2 39209 39213
0 39215 5 1 1 39214
0 39216 7 1 2 84715 39215
0 39217 5 1 1 39216
0 39218 7 2 2 93312 94825
0 39219 5 1 1 101168
0 39220 7 1 2 67500 83999
0 39221 5 1 1 39220
0 39222 7 1 2 3503 39221
0 39223 5 1 1 39222
0 39224 7 2 2 61637 39223
0 39225 5 2 1 101170
0 39226 7 2 2 79372 85005
0 39227 5 1 1 101174
0 39228 7 1 2 63985 39227
0 39229 5 1 1 39228
0 39230 7 1 2 101171 39229
0 39231 5 1 1 39230
0 39232 7 1 2 39219 39231
0 39233 5 1 1 39232
0 39234 7 1 2 96424 39233
0 39235 5 1 1 39234
0 39236 7 1 2 39217 39235
0 39237 5 1 1 39236
0 39238 7 1 2 67025 39237
0 39239 5 1 1 39238
0 39240 7 1 2 78935 93223
0 39241 5 1 1 39240
0 39242 7 1 2 84112 101096
0 39243 5 1 1 39242
0 39244 7 1 2 39241 39243
0 39245 5 1 1 39244
0 39246 7 1 2 66526 39245
0 39247 5 1 1 39246
0 39248 7 1 2 76375 88127
0 39249 7 1 2 95654 39248
0 39250 5 1 1 39249
0 39251 7 1 2 39247 39250
0 39252 5 1 1 39251
0 39253 7 1 2 88214 39252
0 39254 5 1 1 39253
0 39255 7 4 2 63611 89938
0 39256 7 2 2 80152 101176
0 39257 7 1 2 85127 80670
0 39258 7 1 2 101180 39257
0 39259 5 1 1 39258
0 39260 7 1 2 39254 39259
0 39261 5 1 1 39260
0 39262 7 1 2 87674 39261
0 39263 5 1 1 39262
0 39264 7 1 2 39239 39263
0 39265 5 1 1 39264
0 39266 7 1 2 65823 39265
0 39267 5 1 1 39266
0 39268 7 1 2 75783 92890
0 39269 5 1 1 39268
0 39270 7 1 2 4917 101063
0 39271 5 1 1 39270
0 39272 7 3 2 78660 72376
0 39273 7 1 2 69607 101182
0 39274 7 1 2 39271 39273
0 39275 5 1 1 39274
0 39276 7 1 2 39269 39275
0 39277 5 1 1 39276
0 39278 7 1 2 64553 80142
0 39279 7 1 2 39277 39278
0 39280 5 1 1 39279
0 39281 7 1 2 89780 83618
0 39282 7 1 2 91826 92602
0 39283 7 1 2 39281 39282
0 39284 5 1 1 39283
0 39285 7 1 2 39280 39284
0 39286 5 1 1 39285
0 39287 7 1 2 61638 39286
0 39288 5 1 1 39287
0 39289 7 1 2 88692 99760
0 39290 7 1 2 82801 39289
0 39291 5 1 1 39290
0 39292 7 1 2 39288 39291
0 39293 7 1 2 39267 39292
0 39294 5 1 1 39293
0 39295 7 1 2 65192 39294
0 39296 5 1 1 39295
0 39297 7 1 2 91208 92509
0 39298 7 1 2 95888 39297
0 39299 5 1 1 39298
0 39300 7 1 2 78772 82922
0 39301 5 1 1 39300
0 39302 7 1 2 94551 39301
0 39303 5 1 1 39302
0 39304 7 1 2 61639 39303
0 39305 5 1 1 39304
0 39306 7 1 2 90591 97390
0 39307 5 1 1 39306
0 39308 7 1 2 39305 39307
0 39309 5 1 1 39308
0 39310 7 1 2 82285 85574
0 39311 7 1 2 39309 39310
0 39312 5 1 1 39311
0 39313 7 1 2 39299 39312
0 39314 5 1 1 39313
0 39315 7 1 2 69608 39314
0 39316 5 1 1 39315
0 39317 7 1 2 79454 79503
0 39318 7 1 2 87548 39317
0 39319 5 1 1 39318
0 39320 7 1 2 39316 39319
0 39321 5 1 1 39320
0 39322 7 1 2 65499 77378
0 39323 7 1 2 39321 39322
0 39324 5 1 1 39323
0 39325 7 1 2 39296 39324
0 39326 7 1 2 39195 39325
0 39327 5 1 1 39326
0 39328 7 1 2 66024 39327
0 39329 5 1 1 39328
0 39330 7 1 2 71858 85013
0 39331 7 1 2 85732 39330
0 39332 5 1 1 39331
0 39333 7 1 2 95628 39332
0 39334 5 1 1 39333
0 39335 7 1 2 74335 39334
0 39336 5 1 1 39335
0 39337 7 1 2 88676 82537
0 39338 7 1 2 101097 39337
0 39339 5 1 1 39338
0 39340 7 1 2 39336 39339
0 39341 5 1 1 39340
0 39342 7 1 2 63195 39341
0 39343 5 1 1 39342
0 39344 7 1 2 85733 88488
0 39345 7 1 2 94159 39344
0 39346 5 1 1 39345
0 39347 7 1 2 39343 39346
0 39348 5 1 1 39347
0 39349 7 1 2 64775 39348
0 39350 5 1 1 39349
0 39351 7 1 2 75920 75265
0 39352 5 1 1 39351
0 39353 7 1 2 94809 95615
0 39354 5 1 1 39353
0 39355 7 1 2 39352 39354
0 39356 5 1 1 39355
0 39357 7 1 2 88326 39356
0 39358 5 1 1 39357
0 39359 7 1 2 39350 39358
0 39360 5 1 1 39359
0 39361 7 1 2 65824 39360
0 39362 5 1 1 39361
0 39363 7 1 2 82799 81144
0 39364 7 1 2 99761 39363
0 39365 5 1 1 39364
0 39366 7 1 2 39362 39365
0 39367 5 1 1 39366
0 39368 7 1 2 69023 39367
0 39369 5 1 1 39368
0 39370 7 2 2 85518 94837
0 39371 7 1 2 78959 101185
0 39372 5 1 1 39371
0 39373 7 2 2 62614 80747
0 39374 7 1 2 63832 81072
0 39375 7 1 2 101187 39374
0 39376 5 1 1 39375
0 39377 7 1 2 68693 77174
0 39378 7 1 2 91456 39377
0 39379 5 1 1 39378
0 39380 7 1 2 39376 39379
0 39381 5 1 1 39380
0 39382 7 1 2 64165 89725
0 39383 7 1 2 39381 39382
0 39384 5 1 1 39383
0 39385 7 1 2 39372 39384
0 39386 5 1 1 39385
0 39387 7 1 2 67026 39386
0 39388 5 1 1 39387
0 39389 7 1 2 74227 98974
0 39390 7 1 2 101181 39389
0 39391 5 1 1 39390
0 39392 7 1 2 39388 39391
0 39393 5 1 1 39392
0 39394 7 1 2 78431 39393
0 39395 5 1 1 39394
0 39396 7 1 2 39369 39395
0 39397 5 1 1 39396
0 39398 7 1 2 82119 39397
0 39399 5 1 1 39398
0 39400 7 1 2 94216 96342
0 39401 5 1 1 39400
0 39402 7 2 2 69024 75225
0 39403 7 1 2 93522 101189
0 39404 5 1 1 39403
0 39405 7 1 2 39401 39404
0 39406 5 1 1 39405
0 39407 7 1 2 65825 39406
0 39408 5 1 1 39407
0 39409 7 1 2 62615 76501
0 39410 7 1 2 79650 39409
0 39411 5 1 1 39410
0 39412 7 1 2 39408 39411
0 39413 5 1 1 39412
0 39414 7 1 2 81776 39413
0 39415 5 1 1 39414
0 39416 7 1 2 71759 95967
0 39417 7 1 2 90808 39416
0 39418 5 1 1 39417
0 39419 7 1 2 39415 39418
0 39420 5 1 1 39419
0 39421 7 1 2 70953 39420
0 39422 5 1 1 39421
0 39423 7 2 2 65500 94583
0 39424 7 1 2 63384 95927
0 39425 7 1 2 101191 39424
0 39426 5 1 1 39425
0 39427 7 1 2 39422 39426
0 39428 5 1 1 39427
0 39429 7 1 2 79373 39428
0 39430 5 1 1 39429
0 39431 7 1 2 72836 101186
0 39432 5 1 1 39431
0 39433 7 1 2 82212 85278
0 39434 5 1 1 39433
0 39435 7 1 2 72837 74051
0 39436 7 1 2 85523 39435
0 39437 5 1 1 39436
0 39438 7 1 2 39434 39437
0 39439 5 1 1 39438
0 39440 7 1 2 68220 39439
0 39441 5 1 1 39440
0 39442 7 1 2 39432 39441
0 39443 5 1 1 39442
0 39444 7 1 2 84079 80262
0 39445 7 1 2 39443 39444
0 39446 5 1 1 39445
0 39447 7 1 2 67027 39446
0 39448 7 1 2 39430 39447
0 39449 5 1 1 39448
0 39450 7 4 2 70420 75546
0 39451 7 1 2 85791 101193
0 39452 5 1 1 39451
0 39453 7 1 2 74663 79504
0 39454 5 2 1 39453
0 39455 7 1 2 39452 101197
0 39456 5 1 1 39455
0 39457 7 1 2 84093 39456
0 39458 5 1 1 39457
0 39459 7 1 2 74438 80653
0 39460 7 1 2 97939 39459
0 39461 5 1 1 39460
0 39462 7 1 2 39458 39461
0 39463 5 1 1 39462
0 39464 7 1 2 88215 39463
0 39465 5 1 1 39464
0 39466 7 1 2 88786 82996
0 39467 7 1 2 90809 39466
0 39468 5 1 1 39467
0 39469 7 1 2 39465 39468
0 39470 5 1 1 39469
0 39471 7 1 2 69025 39470
0 39472 5 1 1 39471
0 39473 7 3 2 69026 80327
0 39474 7 1 2 80143 101199
0 39475 5 1 1 39474
0 39476 7 1 2 88364 77835
0 39477 5 1 1 39476
0 39478 7 1 2 39475 39477
0 39479 5 1 1 39478
0 39480 7 1 2 86340 39479
0 39481 5 1 1 39480
0 39482 7 2 2 81826 79455
0 39483 7 1 2 82513 101202
0 39484 7 1 2 87528 39483
0 39485 5 1 1 39484
0 39486 7 1 2 39481 39485
0 39487 5 1 1 39486
0 39488 7 1 2 71349 39487
0 39489 5 1 1 39488
0 39490 7 1 2 88749 80362
0 39491 7 1 2 98269 39490
0 39492 5 1 1 39491
0 39493 7 1 2 62182 39492
0 39494 7 1 2 39489 39493
0 39495 7 1 2 39472 39494
0 39496 5 1 1 39495
0 39497 7 1 2 61640 39496
0 39498 7 1 2 39449 39497
0 39499 5 1 1 39498
0 39500 7 1 2 39399 39499
0 39501 5 1 1 39500
0 39502 7 1 2 65193 39501
0 39503 5 1 1 39502
0 39504 7 1 2 79912 97391
0 39505 5 1 1 39504
0 39506 7 1 2 90525 96741
0 39507 7 1 2 76743 39506
0 39508 5 1 1 39507
0 39509 7 1 2 39505 39508
0 39510 5 1 1 39509
0 39511 7 1 2 63833 39510
0 39512 5 1 1 39511
0 39513 7 1 2 71350 76056
0 39514 5 1 1 39513
0 39515 7 1 2 36082 39514
0 39516 5 1 1 39515
0 39517 7 1 2 89687 39516
0 39518 5 1 1 39517
0 39519 7 1 2 39512 39518
0 39520 5 1 1 39519
0 39521 7 1 2 81643 39520
0 39522 5 1 1 39521
0 39523 7 1 2 89583 87153
0 39524 5 1 1 39523
0 39525 7 1 2 39522 39524
0 39526 5 1 1 39525
0 39527 7 1 2 64554 39526
0 39528 5 1 1 39527
0 39529 7 1 2 72838 89170
0 39530 7 1 2 96603 39529
0 39531 5 1 1 39530
0 39532 7 1 2 39528 39531
0 39533 5 1 1 39532
0 39534 7 1 2 76717 39533
0 39535 5 1 1 39534
0 39536 7 1 2 94190 33476
0 39537 5 1 1 39536
0 39538 7 1 2 87498 91487
0 39539 7 1 2 93544 39538
0 39540 7 1 2 39537 39539
0 39541 5 1 1 39540
0 39542 7 1 2 39535 39541
0 39543 5 1 1 39542
0 39544 7 1 2 69609 39543
0 39545 5 1 1 39544
0 39546 7 1 2 4151 95691
0 39547 5 1 1 39546
0 39548 7 1 2 77872 92388
0 39549 7 1 2 94198 39548
0 39550 7 1 2 39547 39549
0 39551 5 1 1 39550
0 39552 7 1 2 39545 39551
0 39553 5 1 1 39552
0 39554 7 1 2 77379 39553
0 39555 5 1 1 39554
0 39556 7 1 2 39503 39555
0 39557 7 1 2 39329 39556
0 39558 5 1 1 39557
0 39559 7 1 2 98667 39558
0 39560 5 1 1 39559
0 39561 7 1 2 86353 97135
0 39562 5 1 1 39561
0 39563 7 2 2 71741 85879
0 39564 7 1 2 63834 101204
0 39565 5 1 1 39564
0 39566 7 1 2 39562 39565
0 39567 5 1 1 39566
0 39568 7 1 2 75811 39567
0 39569 5 1 1 39568
0 39570 7 1 2 72295 91568
0 39571 5 1 1 39570
0 39572 7 1 2 88324 86704
0 39573 5 1 1 39572
0 39574 7 1 2 39571 39573
0 39575 7 1 2 39569 39574
0 39576 5 1 1 39575
0 39577 7 1 2 68869 39576
0 39578 5 1 1 39577
0 39579 7 1 2 74868 101145
0 39580 5 1 1 39579
0 39581 7 2 2 71982 78301
0 39582 5 1 1 101206
0 39583 7 1 2 39580 39582
0 39584 5 1 1 39583
0 39585 7 1 2 77666 39584
0 39586 5 1 1 39585
0 39587 7 1 2 39578 39586
0 39588 5 1 1 39587
0 39589 7 1 2 67718 39588
0 39590 5 1 1 39589
0 39591 7 1 2 70745 76448
0 39592 5 1 1 39591
0 39593 7 1 2 72182 86467
0 39594 7 1 2 39592 39593
0 39595 5 1 1 39594
0 39596 7 2 2 70118 96324
0 39597 7 1 2 72068 86505
0 39598 7 1 2 94006 39597
0 39599 5 1 1 39598
0 39600 7 1 2 101208 39599
0 39601 7 1 2 39595 39600
0 39602 5 1 1 39601
0 39603 7 1 2 39590 39602
0 39604 5 1 1 39603
0 39605 7 1 2 67501 39604
0 39606 5 1 1 39605
0 39607 7 1 2 64166 100394
0 39608 5 2 1 39607
0 39609 7 1 2 72305 101210
0 39610 5 1 1 39609
0 39611 7 1 2 71983 39610
0 39612 5 1 1 39611
0 39613 7 1 2 86126 39612
0 39614 5 1 1 39613
0 39615 7 1 2 67719 39614
0 39616 5 1 1 39615
0 39617 7 1 2 72339 94001
0 39618 5 1 1 39617
0 39619 7 1 2 86020 85041
0 39620 5 1 1 39619
0 39621 7 1 2 39618 39620
0 39622 7 1 2 39616 39621
0 39623 5 1 1 39622
0 39624 7 1 2 68453 39623
0 39625 5 1 1 39624
0 39626 7 1 2 67720 101146
0 39627 5 2 1 39626
0 39628 7 1 2 65501 86806
0 39629 5 1 1 39628
0 39630 7 1 2 101212 39629
0 39631 5 2 1 39630
0 39632 7 1 2 68870 101214
0 39633 5 1 1 39632
0 39634 7 1 2 79980 76718
0 39635 5 1 1 39634
0 39636 7 1 2 39633 39635
0 39637 7 1 2 39625 39636
0 39638 5 1 1 39637
0 39639 7 1 2 101209 39638
0 39640 5 1 1 39639
0 39641 7 1 2 68454 89689
0 39642 7 1 2 101205 39641
0 39643 5 1 1 39642
0 39644 7 1 2 39640 39643
0 39645 7 1 2 39606 39644
0 39646 5 1 1 39645
0 39647 7 1 2 68221 39646
0 39648 5 1 1 39647
0 39649 7 1 2 72842 91603
0 39650 5 1 1 39649
0 39651 7 1 2 84660 91989
0 39652 5 1 1 39651
0 39653 7 1 2 39650 39652
0 39654 5 1 1 39653
0 39655 7 1 2 81054 84801
0 39656 7 1 2 39654 39655
0 39657 5 1 1 39656
0 39658 7 1 2 39648 39657
0 39659 5 1 1 39658
0 39660 7 1 2 76095 39659
0 39661 5 1 1 39660
0 39662 7 1 2 90291 86362
0 39663 5 1 1 39662
0 39664 7 1 2 90399 87290
0 39665 5 1 1 39664
0 39666 7 1 2 39663 39665
0 39667 5 1 1 39666
0 39668 7 1 2 63385 39667
0 39669 5 1 1 39668
0 39670 7 1 2 76376 94568
0 39671 5 1 1 39670
0 39672 7 2 2 68871 75812
0 39673 7 1 2 70746 101216
0 39674 5 1 1 39673
0 39675 7 1 2 16772 39674
0 39676 5 1 1 39675
0 39677 7 1 2 74570 39676
0 39678 5 1 1 39677
0 39679 7 1 2 39671 39678
0 39680 5 1 1 39679
0 39681 7 1 2 67502 39680
0 39682 5 1 1 39681
0 39683 7 1 2 67028 73886
0 39684 5 1 1 39683
0 39685 7 1 2 37964 39684
0 39686 5 1 1 39685
0 39687 7 1 2 77547 39686
0 39688 5 1 1 39687
0 39689 7 1 2 39682 39688
0 39690 5 1 1 39689
0 39691 7 1 2 85841 39690
0 39692 5 1 1 39691
0 39693 7 1 2 68455 96986
0 39694 5 1 1 39693
0 39695 7 1 2 39692 39694
0 39696 5 1 1 39695
0 39697 7 1 2 81845 39696
0 39698 5 1 1 39697
0 39699 7 1 2 65194 39698
0 39700 7 1 2 39669 39699
0 39701 5 1 1 39700
0 39702 7 1 2 72463 84979
0 39703 5 1 1 39702
0 39704 7 1 2 25934 39703
0 39705 5 1 1 39704
0 39706 7 1 2 67029 39705
0 39707 5 1 1 39706
0 39708 7 1 2 88511 93495
0 39709 5 1 1 39708
0 39710 7 1 2 39707 39709
0 39711 5 1 1 39710
0 39712 7 1 2 72183 39711
0 39713 5 1 1 39712
0 39714 7 1 2 71984 96667
0 39715 5 1 1 39714
0 39716 7 1 2 86127 39715
0 39717 5 1 1 39716
0 39718 7 1 2 74336 39717
0 39719 5 1 1 39718
0 39720 7 1 2 86705 76485
0 39721 7 1 2 62183 95625
0 39722 5 2 1 39721
0 39723 7 1 2 63612 95626
0 39724 5 2 1 39723
0 39725 7 1 2 101218 101220
0 39726 7 1 2 39720 39725
0 39727 5 1 1 39726
0 39728 7 1 2 39719 39727
0 39729 5 1 1 39728
0 39730 7 1 2 67721 39729
0 39731 5 1 1 39730
0 39732 7 1 2 6776 101213
0 39733 5 1 1 39732
0 39734 7 1 2 73482 39733
0 39735 5 1 1 39734
0 39736 7 2 2 65826 74926
0 39737 5 1 1 101222
0 39738 7 1 2 85678 39737
0 39739 5 1 1 39738
0 39740 7 1 2 72069 39739
0 39741 5 1 1 39740
0 39742 7 1 2 94573 39741
0 39743 7 1 2 39735 39742
0 39744 5 1 1 39743
0 39745 7 1 2 99128 39744
0 39746 5 1 1 39745
0 39747 7 1 2 73483 76025
0 39748 7 1 2 101207 39747
0 39749 5 1 1 39748
0 39750 7 1 2 39746 39749
0 39751 7 1 2 39731 39750
0 39752 7 1 2 39713 39751
0 39753 5 1 1 39752
0 39754 7 1 2 81846 39753
0 39755 5 1 1 39754
0 39756 7 2 2 70421 85425
0 39757 7 1 2 62184 85965
0 39758 5 1 1 39757
0 39759 7 1 2 101124 39758
0 39760 5 1 1 39759
0 39761 7 1 2 65827 39760
0 39762 5 1 1 39761
0 39763 7 1 2 84726 39762
0 39764 5 1 1 39763
0 39765 7 1 2 63613 39764
0 39766 5 1 1 39765
0 39767 7 1 2 18484 39766
0 39768 5 1 1 39767
0 39769 7 1 2 101224 39768
0 39770 5 1 1 39769
0 39771 7 1 2 70119 39770
0 39772 7 1 2 39755 39771
0 39773 5 1 1 39772
0 39774 7 1 2 68033 39773
0 39775 7 1 2 39701 39774
0 39776 5 1 1 39775
0 39777 7 1 2 39661 39776
0 39778 5 1 1 39777
0 39779 7 1 2 64776 39778
0 39780 5 1 1 39779
0 39781 7 1 2 70747 76478
0 39782 5 1 1 39781
0 39783 7 1 2 24649 39782
0 39784 5 1 1 39783
0 39785 7 1 2 63614 39784
0 39786 5 1 1 39785
0 39787 7 1 2 84903 86746
0 39788 5 1 1 39787
0 39789 7 1 2 86633 39788
0 39790 5 1 1 39789
0 39791 7 1 2 39786 39790
0 39792 5 1 1 39791
0 39793 7 1 2 65502 39792
0 39794 5 1 1 39793
0 39795 7 1 2 76622 86242
0 39796 5 1 1 39795
0 39797 7 1 2 74941 75212
0 39798 5 1 1 39797
0 39799 7 1 2 39796 39798
0 39800 5 1 1 39799
0 39801 7 1 2 62435 39800
0 39802 5 1 1 39801
0 39803 7 1 2 84772 39802
0 39804 5 1 1 39803
0 39805 7 1 2 72464 39804
0 39806 5 1 1 39805
0 39807 7 1 2 39794 39806
0 39808 5 1 1 39807
0 39809 7 1 2 80987 88276
0 39810 7 1 2 39808 39809
0 39811 5 1 1 39810
0 39812 7 1 2 39780 39811
0 39813 5 1 1 39812
0 39814 7 1 2 69407 39813
0 39815 5 1 1 39814
0 39816 7 1 2 72872 86128
0 39817 5 1 1 39816
0 39818 7 1 2 68456 39817
0 39819 5 1 1 39818
0 39820 7 1 2 76654 86419
0 39821 5 1 1 39820
0 39822 7 1 2 39819 39821
0 39823 5 1 1 39822
0 39824 7 1 2 90150 39823
0 39825 5 1 1 39824
0 39826 7 1 2 79262 85438
0 39827 5 1 1 39826
0 39828 7 1 2 39825 39827
0 39829 5 1 1 39828
0 39830 7 1 2 62436 39829
0 39831 5 1 1 39830
0 39832 7 1 2 88350 75813
0 39833 7 1 2 73484 84345
0 39834 7 1 2 39832 39833
0 39835 7 1 2 96872 39834
0 39836 5 1 1 39835
0 39837 7 1 2 39831 39836
0 39838 5 1 1 39837
0 39839 7 1 2 63835 39838
0 39840 5 1 1 39839
0 39841 7 1 2 85243 85347
0 39842 5 1 1 39841
0 39843 7 1 2 71260 86071
0 39844 5 1 1 39843
0 39845 7 1 2 39842 39844
0 39846 5 1 1 39845
0 39847 7 1 2 63615 39846
0 39848 5 1 1 39847
0 39849 7 1 2 75035 86072
0 39850 5 1 1 39849
0 39851 7 1 2 39848 39850
0 39852 5 1 1 39851
0 39853 7 1 2 66025 39852
0 39854 5 1 1 39853
0 39855 7 2 2 73342 73836
0 39856 7 1 2 84030 101226
0 39857 5 1 1 39856
0 39858 7 1 2 39854 39857
0 39859 5 1 1 39858
0 39860 7 1 2 68694 39859
0 39861 5 1 1 39860
0 39862 7 1 2 85625 86125
0 39863 5 1 1 39862
0 39864 7 1 2 39861 39863
0 39865 5 1 1 39864
0 39866 7 1 2 90151 39865
0 39867 5 1 1 39866
0 39868 7 1 2 39840 39867
0 39869 5 1 1 39868
0 39870 7 1 2 81777 39869
0 39871 5 1 1 39870
0 39872 7 1 2 65828 94563
0 39873 5 1 1 39872
0 39874 7 1 2 68695 84551
0 39875 5 1 1 39874
0 39876 7 1 2 62616 39875
0 39877 5 1 1 39876
0 39878 7 1 2 67293 4753
0 39879 7 1 2 39877 39878
0 39880 5 1 1 39879
0 39881 7 1 2 17583 39880
0 39882 7 1 2 39873 39881
0 39883 5 1 1 39882
0 39884 7 1 2 65503 39883
0 39885 5 1 1 39884
0 39886 7 1 2 89588 79987
0 39887 5 1 1 39886
0 39888 7 1 2 39885 39887
0 39889 5 1 1 39888
0 39890 7 1 2 94284 39889
0 39891 5 1 1 39890
0 39892 7 1 2 91488 95844
0 39893 5 1 1 39892
0 39894 7 1 2 73485 86201
0 39895 5 1 1 39894
0 39896 7 1 2 91470 39895
0 39897 5 1 1 39896
0 39898 7 1 2 39893 39897
0 39899 5 1 1 39898
0 39900 7 1 2 64167 76489
0 39901 7 1 2 39899 39900
0 39902 5 1 1 39901
0 39903 7 1 2 39891 39902
0 39904 5 1 1 39903
0 39905 7 1 2 65195 39904
0 39906 5 1 1 39905
0 39907 7 1 2 85445 85675
0 39908 5 1 1 39907
0 39909 7 1 2 84031 75461
0 39910 5 1 1 39909
0 39911 7 1 2 62185 80431
0 39912 5 1 1 39911
0 39913 7 1 2 39910 39912
0 39914 5 1 1 39913
0 39915 7 1 2 70120 39914
0 39916 5 1 1 39915
0 39917 7 2 2 63836 80756
0 39918 7 1 2 74392 85676
0 39919 7 1 2 101228 39918
0 39920 5 1 1 39919
0 39921 7 1 2 39916 39920
0 39922 5 1 1 39921
0 39923 7 1 2 62437 39922
0 39924 5 1 1 39923
0 39925 7 1 2 39908 39924
0 39926 5 1 1 39925
0 39927 7 1 2 76178 39926
0 39928 5 1 1 39927
0 39929 7 1 2 84956 93653
0 39930 5 1 1 39929
0 39931 7 1 2 520 5275
0 39932 5 2 1 39931
0 39933 7 1 2 68696 101230
0 39934 5 1 1 39933
0 39935 7 1 2 99186 39934
0 39936 5 1 1 39935
0 39937 7 1 2 79394 39936
0 39938 5 1 1 39937
0 39939 7 1 2 39930 39938
0 39940 5 1 1 39939
0 39941 7 1 2 66527 92540
0 39942 7 1 2 39940 39941
0 39943 5 1 1 39942
0 39944 7 1 2 39928 39943
0 39945 7 1 2 39906 39944
0 39946 5 1 1 39945
0 39947 7 1 2 63386 39946
0 39948 5 1 1 39947
0 39949 7 1 2 39871 39948
0 39950 5 1 1 39949
0 39951 7 1 2 69610 39950
0 39952 5 1 1 39951
0 39953 7 2 2 65504 76480
0 39954 5 1 1 101232
0 39955 7 1 2 86563 39954
0 39956 5 1 1 39955
0 39957 7 1 2 78448 39956
0 39958 5 1 1 39957
0 39959 7 1 2 86180 18615
0 39960 7 1 2 25623 39959
0 39961 5 1 1 39960
0 39962 7 1 2 39958 39961
0 39963 5 1 1 39962
0 39964 7 1 2 63616 39963
0 39965 5 1 1 39964
0 39966 7 1 2 85229 101129
0 39967 5 1 1 39966
0 39968 7 1 2 39965 39967
0 39969 5 1 1 39968
0 39970 7 1 2 70121 39969
0 39971 5 1 1 39970
0 39972 7 1 2 73078 76537
0 39973 5 1 1 39972
0 39974 7 1 2 39971 39973
0 39975 5 1 1 39974
0 39976 7 1 2 72565 39975
0 39977 5 1 1 39976
0 39978 7 1 2 79559 74291
0 39979 5 1 1 39978
0 39980 7 1 2 39977 39979
0 39981 5 1 1 39980
0 39982 7 1 2 97294 39981
0 39983 5 1 1 39982
0 39984 7 1 2 39952 39983
0 39985 5 1 1 39984
0 39986 7 1 2 64555 39985
0 39987 5 1 1 39986
0 39988 7 1 2 90838 80671
0 39989 7 1 2 95048 39988
0 39990 5 1 1 39989
0 39991 7 1 2 78960 92694
0 39992 5 1 1 39991
0 39993 7 1 2 27485 39992
0 39994 5 1 1 39993
0 39995 7 1 2 61641 39994
0 39996 5 1 1 39995
0 39997 7 1 2 91485 95049
0 39998 5 1 1 39997
0 39999 7 1 2 39996 39998
0 40000 5 1 1 39999
0 40001 7 1 2 64556 76275
0 40002 7 1 2 40000 40001
0 40003 5 1 1 40002
0 40004 7 1 2 39990 40003
0 40005 5 1 1 40004
0 40006 7 1 2 71859 40005
0 40007 5 1 1 40006
0 40008 7 1 2 82142 79263
0 40009 7 1 2 90805 40008
0 40010 7 1 2 90839 40009
0 40011 5 1 1 40010
0 40012 7 1 2 40007 40011
0 40013 5 1 1 40012
0 40014 7 1 2 70422 40013
0 40015 5 1 1 40014
0 40016 7 1 2 66528 92515
0 40017 7 1 2 94916 40016
0 40018 5 1 1 40017
0 40019 7 1 2 76057 96771
0 40020 7 1 2 101083 40019
0 40021 5 1 1 40020
0 40022 7 1 2 40018 40021
0 40023 5 1 1 40022
0 40024 7 1 2 79456 40023
0 40025 5 1 1 40024
0 40026 7 1 2 40015 40025
0 40027 5 1 1 40026
0 40028 7 1 2 70122 40027
0 40029 5 1 1 40028
0 40030 7 2 2 85014 97770
0 40031 7 1 2 88512 101234
0 40032 5 1 1 40031
0 40033 7 2 2 82683 82250
0 40034 7 1 2 76471 76276
0 40035 7 1 2 101236 40034
0 40036 5 1 1 40035
0 40037 7 1 2 40032 40036
0 40038 5 1 1 40037
0 40039 7 1 2 87067 83782
0 40040 7 1 2 40038 40039
0 40041 5 1 1 40040
0 40042 7 1 2 40029 40041
0 40043 5 1 1 40042
0 40044 7 1 2 78334 40043
0 40045 5 1 1 40044
0 40046 7 1 2 82559 8967
0 40047 5 1 1 40046
0 40048 7 1 2 79264 40047
0 40049 5 1 1 40048
0 40050 7 1 2 88644 82431
0 40051 5 1 1 40050
0 40052 7 1 2 40049 40051
0 40053 5 1 1 40052
0 40054 7 1 2 91724 40053
0 40055 5 1 1 40054
0 40056 7 1 2 91920 93185
0 40057 5 1 1 40056
0 40058 7 1 2 40055 40057
0 40059 5 1 1 40058
0 40060 7 1 2 65829 40059
0 40061 5 1 1 40060
0 40062 7 1 2 87068 96443
0 40063 7 1 2 95577 40062
0 40064 5 1 1 40063
0 40065 7 1 2 77380 82865
0 40066 7 1 2 98930 40065
0 40067 5 1 1 40066
0 40068 7 1 2 40064 40067
0 40069 5 1 1 40068
0 40070 7 1 2 71860 40069
0 40071 5 1 1 40070
0 40072 7 1 2 81847 91557
0 40073 7 1 2 101175 40072
0 40074 5 1 1 40073
0 40075 7 1 2 40071 40074
0 40076 7 1 2 40061 40075
0 40077 5 1 1 40076
0 40078 7 1 2 65505 40077
0 40079 5 1 1 40078
0 40080 7 1 2 82297 91571
0 40081 5 1 1 40080
0 40082 7 2 2 74374 84080
0 40083 7 1 2 101238 100067
0 40084 5 1 1 40083
0 40085 7 1 2 40081 40084
0 40086 5 1 1 40085
0 40087 7 1 2 65830 40086
0 40088 5 1 1 40087
0 40089 7 1 2 74684 83653
0 40090 7 1 2 82316 40089
0 40091 5 1 1 40090
0 40092 7 1 2 40088 40091
0 40093 5 1 1 40092
0 40094 7 1 2 100857 40093
0 40095 5 1 1 40094
0 40096 7 1 2 40079 40095
0 40097 5 1 1 40096
0 40098 7 1 2 98297 40097
0 40099 5 1 1 40098
0 40100 7 1 2 9356 29840
0 40101 5 1 1 40100
0 40102 7 1 2 88570 101007
0 40103 5 1 1 40102
0 40104 7 1 2 90843 96525
0 40105 5 1 1 40104
0 40106 7 1 2 88598 86253
0 40107 5 1 1 40106
0 40108 7 1 2 40105 40107
0 40109 5 1 1 40108
0 40110 7 1 2 73741 40109
0 40111 5 1 1 40110
0 40112 7 1 2 40103 40111
0 40113 5 1 1 40112
0 40114 7 1 2 65506 40113
0 40115 5 1 1 40114
0 40116 7 1 2 74603 91096
0 40117 7 1 2 100887 40116
0 40118 5 1 1 40117
0 40119 7 1 2 40115 40118
0 40120 5 1 1 40119
0 40121 7 1 2 40101 40120
0 40122 5 1 1 40121
0 40123 7 1 2 40099 40122
0 40124 7 1 2 40045 40123
0 40125 7 1 2 74205 101090
0 40126 5 1 1 40125
0 40127 7 1 2 63387 77122
0 40128 5 1 1 40127
0 40129 7 1 2 40126 40128
0 40130 5 1 1 40129
0 40131 7 1 2 71861 40130
0 40132 5 1 1 40131
0 40133 7 1 2 66026 94075
0 40134 5 1 1 40133
0 40135 7 1 2 7445 40134
0 40136 5 1 1 40135
0 40137 7 1 2 63388 40136
0 40138 5 1 1 40137
0 40139 7 1 2 40132 40138
0 40140 5 1 1 40139
0 40141 7 1 2 83593 40140
0 40142 5 1 1 40141
0 40143 7 1 2 82883 79970
0 40144 7 1 2 91748 40143
0 40145 5 1 1 40144
0 40146 7 1 2 40142 40145
0 40147 5 1 1 40146
0 40148 7 1 2 84081 40147
0 40149 5 1 1 40148
0 40150 7 1 2 87069 86529
0 40151 7 1 2 92300 40150
0 40152 5 1 1 40151
0 40153 7 1 2 40149 40152
0 40154 5 1 1 40153
0 40155 7 1 2 66529 40154
0 40156 5 1 1 40155
0 40157 7 1 2 68697 97136
0 40158 5 1 1 40157
0 40159 7 1 2 65196 86075
0 40160 5 1 1 40159
0 40161 7 1 2 40158 40160
0 40162 5 1 1 40161
0 40163 7 1 2 81700 88103
0 40164 7 1 2 92101 40163
0 40165 7 1 2 40162 40164
0 40166 5 1 1 40165
0 40167 7 1 2 40156 40166
0 40168 5 1 1 40167
0 40169 7 1 2 62186 40168
0 40170 5 1 1 40169
0 40171 7 2 2 88254 91321
0 40172 5 2 1 101240
0 40173 7 1 2 78241 101241
0 40174 5 1 1 40173
0 40175 7 1 2 8568 40174
0 40176 5 1 1 40175
0 40177 7 1 2 91670 40176
0 40178 5 1 1 40177
0 40179 7 2 2 69408 87070
0 40180 7 1 2 71638 101244
0 40181 7 1 2 92127 40180
0 40182 5 1 1 40181
0 40183 7 1 2 40178 40182
0 40184 5 1 1 40183
0 40185 7 1 2 70748 40184
0 40186 5 1 1 40185
0 40187 7 1 2 68698 77255
0 40188 7 1 2 81644 40187
0 40189 7 3 2 64168 82997
0 40190 7 1 2 97302 101246
0 40191 7 1 2 40188 40190
0 40192 5 1 1 40191
0 40193 7 1 2 40186 40192
0 40194 5 1 1 40193
0 40195 7 1 2 86438 40194
0 40196 5 1 1 40195
0 40197 7 1 2 85391 92576
0 40198 7 1 2 97030 40197
0 40199 5 1 1 40198
0 40200 7 1 2 40196 40199
0 40201 7 1 2 40170 40200
0 40202 5 1 1 40201
0 40203 7 1 2 71351 40202
0 40204 5 1 1 40203
0 40205 7 1 2 73486 100969
0 40206 5 1 1 40205
0 40207 7 1 2 84890 90137
0 40208 5 1 1 40207
0 40209 7 1 2 78449 93725
0 40210 5 1 1 40209
0 40211 7 1 2 68699 40210
0 40212 5 1 1 40211
0 40213 7 1 2 1331 29575
0 40214 7 1 2 40212 40213
0 40215 5 1 1 40214
0 40216 7 1 2 71261 40215
0 40217 5 1 1 40216
0 40218 7 1 2 40208 40217
0 40219 7 1 2 40206 40218
0 40220 5 1 1 40219
0 40221 7 1 2 67294 40220
0 40222 5 1 1 40221
0 40223 7 1 2 90138 94584
0 40224 5 1 1 40223
0 40225 7 1 2 40222 40224
0 40226 5 1 1 40225
0 40227 7 1 2 84213 87054
0 40228 7 1 2 40226 40227
0 40229 5 1 1 40228
0 40230 7 2 2 88759 86653
0 40231 5 1 1 101249
0 40232 7 2 2 71862 101250
0 40233 5 1 1 101251
0 40234 7 1 2 70423 101252
0 40235 5 1 1 40234
0 40236 7 1 2 78242 101231
0 40237 5 1 1 40236
0 40238 7 1 2 20028 40231
0 40239 5 1 1 40238
0 40240 7 1 2 71863 40239
0 40241 5 1 1 40240
0 40242 7 1 2 77054 40241
0 40243 7 1 2 40237 40242
0 40244 5 1 1 40243
0 40245 7 1 2 77030 40244
0 40246 5 1 1 40245
0 40247 7 1 2 40235 40246
0 40248 5 1 1 40247
0 40249 7 1 2 62883 40248
0 40250 5 1 1 40249
0 40251 7 1 2 78152 77967
0 40252 7 1 2 77548 76212
0 40253 7 1 2 40251 40252
0 40254 5 1 1 40253
0 40255 7 1 2 40250 40254
0 40256 5 1 1 40255
0 40257 7 1 2 82855 40256
0 40258 5 1 1 40257
0 40259 7 1 2 63389 40258
0 40260 7 1 2 40229 40259
0 40261 5 1 1 40260
0 40262 7 1 2 79400 101157
0 40263 5 1 1 40262
0 40264 7 1 2 86674 92990
0 40265 7 1 2 40263 40264
0 40266 5 1 1 40265
0 40267 7 1 2 73487 86211
0 40268 5 1 1 40267
0 40269 7 1 2 63617 40268
0 40270 5 1 1 40269
0 40271 7 1 2 82120 78827
0 40272 7 1 2 40270 40271
0 40273 5 1 1 40272
0 40274 7 1 2 40266 40273
0 40275 5 1 1 40274
0 40276 7 1 2 70424 40275
0 40277 5 1 1 40276
0 40278 7 1 2 62617 86675
0 40279 7 1 2 75456 40278
0 40280 7 1 2 85197 93425
0 40281 7 1 2 40279 40280
0 40282 5 1 1 40281
0 40283 7 1 2 40277 40282
0 40284 5 1 1 40283
0 40285 7 1 2 71864 40284
0 40286 5 1 1 40285
0 40287 7 1 2 74439 87470
0 40288 7 1 2 95374 40287
0 40289 7 1 2 101076 40288
0 40290 5 1 1 40289
0 40291 7 1 2 68222 40290
0 40292 7 1 2 40286 40291
0 40293 5 1 1 40292
0 40294 7 1 2 78961 40293
0 40295 7 1 2 40261 40294
0 40296 5 1 1 40295
0 40297 7 1 2 40204 40296
0 40298 7 1 2 40124 40297
0 40299 7 1 2 39987 40298
0 40300 7 1 2 39815 40299
0 40301 5 1 1 40300
0 40302 7 1 2 98654 40301
0 40303 5 1 1 40302
0 40304 7 1 2 39560 40303
0 40305 5 1 1 40304
0 40306 7 1 2 64381 40305
0 40307 5 1 1 40306
0 40308 7 1 2 81935 98679
0 40309 5 1 1 40308
0 40310 7 1 2 64777 87686
0 40311 7 1 2 98016 40310
0 40312 7 1 2 93380 40311
0 40313 5 1 1 40312
0 40314 7 1 2 40309 40313
0 40315 5 1 1 40314
0 40316 7 1 2 76538 40315
0 40317 5 1 1 40316
0 40318 7 2 2 70425 91024
0 40319 7 1 2 7597 77647
0 40320 5 1 1 40319
0 40321 7 2 2 66530 73343
0 40322 7 1 2 94733 101255
0 40323 7 1 2 40320 40322
0 40324 7 1 2 101253 40323
0 40325 5 1 1 40324
0 40326 7 1 2 40317 40325
0 40327 5 1 1 40326
0 40328 7 1 2 70749 40327
0 40329 5 1 1 40328
0 40330 7 3 2 66142 99021
0 40331 7 1 2 76539 101257
0 40332 7 2 2 99194 97358
0 40333 7 1 2 101260 101094
0 40334 7 1 2 40331 40333
0 40335 5 1 1 40334
0 40336 7 1 2 40329 40335
0 40337 5 1 1 40336
0 40338 7 1 2 74129 40337
0 40339 5 1 1 40338
0 40340 7 1 2 67030 98994
0 40341 7 1 2 97650 40340
0 40342 7 1 2 98173 40341
0 40343 7 1 2 96567 40342
0 40344 5 1 1 40343
0 40345 7 1 2 91545 98621
0 40346 7 1 2 99254 40345
0 40347 7 1 2 92163 40346
0 40348 5 1 1 40347
0 40349 7 1 2 40344 40348
0 40350 5 1 1 40349
0 40351 7 1 2 66143 40350
0 40352 5 1 1 40351
0 40353 7 1 2 84283 94734
0 40354 7 1 2 90717 40353
0 40355 7 1 2 96568 40354
0 40356 5 1 1 40355
0 40357 7 1 2 40352 40356
0 40358 5 1 1 40357
0 40359 7 1 2 77529 40358
0 40360 5 1 1 40359
0 40361 7 1 2 90441 96560
0 40362 5 1 1 40361
0 40363 7 1 2 96564 40362
0 40364 5 1 1 40363
0 40365 7 1 2 67295 40364
0 40366 5 1 1 40365
0 40367 7 1 2 80886 84877
0 40368 5 1 1 40367
0 40369 7 1 2 40366 40368
0 40370 5 1 1 40369
0 40371 7 1 2 88567 98680
0 40372 7 1 2 40370 40371
0 40373 5 1 1 40372
0 40374 7 1 2 74440 72465
0 40375 7 1 2 80168 40374
0 40376 7 1 2 67876 77444
0 40377 7 1 2 98186 40376
0 40378 7 1 2 97780 40377
0 40379 7 1 2 40375 40378
0 40380 5 1 1 40379
0 40381 7 4 2 65507 91025
0 40382 7 1 2 73922 79958
0 40383 7 1 2 94735 40382
0 40384 7 1 2 19373 40383
0 40385 7 1 2 101262 40384
0 40386 5 1 1 40385
0 40387 7 1 2 72070 74571
0 40388 7 1 2 77516 40387
0 40389 7 2 2 91866 98209
0 40390 7 1 2 97781 101266
0 40391 7 1 2 40388 40390
0 40392 5 1 1 40391
0 40393 7 1 2 40386 40392
0 40394 5 1 1 40393
0 40395 7 1 2 73266 40394
0 40396 5 1 1 40395
0 40397 7 1 2 40380 40396
0 40398 7 1 2 40373 40397
0 40399 7 1 2 40360 40398
0 40400 5 1 1 40399
0 40401 7 1 2 61642 40400
0 40402 5 1 1 40401
0 40403 7 1 2 65508 75746
0 40404 5 4 1 40403
0 40405 7 1 2 69611 76823
0 40406 7 1 2 79265 98847
0 40407 7 1 2 40405 40406
0 40408 7 1 2 101268 40407
0 40409 7 1 2 91026 40408
0 40410 5 1 1 40409
0 40411 7 1 2 40402 40410
0 40412 7 1 2 40339 40411
0 40413 5 1 1 40412
0 40414 7 1 2 64557 40413
0 40415 5 1 1 40414
0 40416 7 2 2 79457 82702
0 40417 7 2 2 68457 98681
0 40418 7 1 2 101272 101274
0 40419 7 1 2 94282 40418
0 40420 5 1 1 40419
0 40421 7 1 2 40415 40420
0 40422 5 1 1 40421
0 40423 7 1 2 63390 40422
0 40424 5 1 1 40423
0 40425 7 3 2 67722 97067
0 40426 5 1 1 101276
0 40427 7 1 2 90265 101277
0 40428 5 1 1 40427
0 40429 7 2 2 69612 100866
0 40430 7 1 2 82856 101279
0 40431 5 1 1 40430
0 40432 7 1 2 40428 40431
0 40433 5 2 1 40432
0 40434 7 1 2 90323 101281
0 40435 5 1 1 40434
0 40436 7 1 2 90266 76213
0 40437 5 1 1 40436
0 40438 7 1 2 40435 40437
0 40439 5 1 1 40438
0 40440 7 1 2 71865 40439
0 40441 5 1 1 40440
0 40442 7 1 2 90867 88128
0 40443 7 1 2 82043 40442
0 40444 5 1 1 40443
0 40445 7 1 2 40441 40444
0 40446 5 1 1 40445
0 40447 7 1 2 77321 40446
0 40448 5 1 1 40447
0 40449 7 1 2 82857 80273
0 40450 7 1 2 90778 40449
0 40451 7 1 2 89051 40450
0 40452 5 1 1 40451
0 40453 7 1 2 40448 40452
0 40454 5 1 1 40453
0 40455 7 1 2 69027 40454
0 40456 5 1 1 40455
0 40457 7 1 2 94021 101005
0 40458 5 1 1 40457
0 40459 7 1 2 72889 98690
0 40460 7 1 2 89521 40459
0 40461 5 1 1 40460
0 40462 7 1 2 40458 40461
0 40463 5 1 1 40462
0 40464 7 1 2 83960 40463
0 40465 5 1 1 40464
0 40466 7 1 2 63618 95540
0 40467 5 1 1 40466
0 40468 7 1 2 94258 98240
0 40469 5 1 1 40468
0 40470 7 1 2 40467 40469
0 40471 5 1 1 40470
0 40472 7 1 2 81200 90315
0 40473 7 1 2 40471 40472
0 40474 5 1 1 40473
0 40475 7 1 2 40465 40474
0 40476 5 1 1 40475
0 40477 7 1 2 65831 40476
0 40478 5 1 1 40477
0 40479 7 1 2 88888 85382
0 40480 5 1 1 40479
0 40481 7 1 2 76216 40480
0 40482 5 1 1 40481
0 40483 7 1 2 90008 76623
0 40484 7 1 2 92281 40483
0 40485 7 1 2 40482 40484
0 40486 5 1 1 40485
0 40487 7 1 2 40478 40486
0 40488 7 1 2 40456 40487
0 40489 5 1 1 40488
0 40490 7 1 2 68223 98682
0 40491 7 1 2 40489 40490
0 40492 5 1 1 40491
0 40493 7 1 2 40424 40492
0 40494 5 1 1 40493
0 40495 7 1 2 63196 40494
0 40496 5 1 1 40495
0 40497 7 1 2 86021 84098
0 40498 5 1 1 40497
0 40499 7 1 2 97862 40498
0 40500 5 1 1 40499
0 40501 7 1 2 95469 40500
0 40502 5 1 1 40501
0 40503 7 1 2 75199 83228
0 40504 7 1 2 79275 40503
0 40505 5 1 1 40504
0 40506 7 1 2 40502 40505
0 40507 5 1 1 40506
0 40508 7 1 2 83669 40507
0 40509 5 1 1 40508
0 40510 7 1 2 78335 90891
0 40511 5 1 1 40510
0 40512 7 1 2 85148 96526
0 40513 5 1 1 40512
0 40514 7 1 2 40511 40513
0 40515 5 1 1 40514
0 40516 7 1 2 62884 40515
0 40517 5 1 1 40516
0 40518 7 1 2 87441 75730
0 40519 5 1 1 40518
0 40520 7 1 2 40517 40519
0 40521 5 1 1 40520
0 40522 7 1 2 101237 40521
0 40523 5 1 1 40522
0 40524 7 1 2 70750 94255
0 40525 5 1 1 40524
0 40526 7 1 2 94230 94319
0 40527 7 1 2 40525 40526
0 40528 5 1 1 40527
0 40529 7 1 2 77934 40528
0 40530 5 1 1 40529
0 40531 7 1 2 94080 99944
0 40532 5 1 1 40531
0 40533 7 1 2 79208 97095
0 40534 7 1 2 40532 40533
0 40535 5 1 1 40534
0 40536 7 1 2 40530 40535
0 40537 5 1 1 40536
0 40538 7 1 2 64169 40537
0 40539 5 1 1 40538
0 40540 7 2 2 62438 86654
0 40541 7 1 2 71596 101283
0 40542 5 1 1 40541
0 40543 7 1 2 86857 40542
0 40544 5 1 1 40543
0 40545 7 1 2 72184 40544
0 40546 5 1 1 40545
0 40547 7 1 2 79405 93333
0 40548 5 1 1 40547
0 40549 7 1 2 101198 40548
0 40550 7 1 2 40546 40549
0 40551 5 1 1 40550
0 40552 7 1 2 63837 40551
0 40553 5 1 1 40552
0 40554 7 1 2 76382 100210
0 40555 5 1 1 40554
0 40556 7 1 2 40553 40555
0 40557 5 1 1 40556
0 40558 7 1 2 67031 40557
0 40559 5 1 1 40558
0 40560 7 2 2 74820 101221
0 40561 7 1 2 84173 95522
0 40562 7 1 2 101285 40561
0 40563 5 1 1 40562
0 40564 7 1 2 40559 40563
0 40565 7 1 2 40539 40564
0 40566 5 1 1 40565
0 40567 7 1 2 86459 40566
0 40568 5 1 1 40567
0 40569 7 1 2 40523 40568
0 40570 5 1 1 40569
0 40571 7 1 2 69613 40570
0 40572 5 1 1 40571
0 40573 7 1 2 40509 40572
0 40574 5 1 1 40573
0 40575 7 2 2 68034 98683
0 40576 7 1 2 40574 101287
0 40577 5 1 1 40576
0 40578 7 1 2 40496 40577
0 40579 5 1 1 40578
0 40580 7 1 2 65197 40579
0 40581 5 1 1 40580
0 40582 7 1 2 92302 96001
0 40583 7 1 2 101110 40582
0 40584 5 1 1 40583
0 40585 7 2 2 71021 93715
0 40586 5 1 1 101289
0 40587 7 1 2 67503 101290
0 40588 5 1 1 40587
0 40589 7 1 2 18122 40588
0 40590 5 1 1 40589
0 40591 7 1 2 90935 40590
0 40592 5 1 1 40591
0 40593 7 2 2 78432 85743
0 40594 7 1 2 82584 88513
0 40595 7 1 2 101291 40594
0 40596 5 1 1 40595
0 40597 7 1 2 40592 40596
0 40598 5 1 1 40597
0 40599 7 1 2 80952 94792
0 40600 7 1 2 40598 40599
0 40601 5 1 1 40600
0 40602 7 1 2 40584 40601
0 40603 5 1 1 40602
0 40604 7 1 2 98684 40603
0 40605 5 1 1 40604
0 40606 7 2 2 69133 70123
0 40607 7 1 2 68224 73815
0 40608 7 1 2 101293 40607
0 40609 7 1 2 99238 40608
0 40610 5 1 1 40609
0 40611 7 1 2 67032 98778
0 40612 7 1 2 77063 40611
0 40613 7 1 2 98737 40612
0 40614 5 1 1 40613
0 40615 7 1 2 40610 40614
0 40616 5 1 1 40615
0 40617 7 1 2 89007 40616
0 40618 5 1 1 40617
0 40619 7 2 2 93055 97774
0 40620 7 1 2 90033 97990
0 40621 7 1 2 95611 40620
0 40622 7 1 2 101295 40621
0 40623 5 1 1 40622
0 40624 7 1 2 40618 40623
0 40625 5 1 1 40624
0 40626 7 1 2 66144 40625
0 40627 5 1 1 40626
0 40628 7 1 2 61387 91805
0 40629 5 1 1 40628
0 40630 7 1 2 35842 40629
0 40631 5 2 1 40630
0 40632 7 2 2 74337 80228
0 40633 7 1 2 88922 97718
0 40634 7 1 2 77064 40633
0 40635 7 1 2 101299 40634
0 40636 7 1 2 101297 40635
0 40637 5 1 1 40636
0 40638 7 1 2 40627 40637
0 40639 5 1 1 40638
0 40640 7 1 2 72566 40639
0 40641 5 1 1 40640
0 40642 7 3 2 69409 101288
0 40643 7 1 2 80619 94860
0 40644 7 1 2 101301 40643
0 40645 5 1 1 40644
0 40646 7 1 2 40641 40645
0 40647 5 1 1 40646
0 40648 7 1 2 71262 40647
0 40649 5 1 1 40648
0 40650 7 1 2 70124 82269
0 40651 5 1 1 40650
0 40652 7 1 2 95744 40651
0 40653 5 1 1 40652
0 40654 7 1 2 94637 101300
0 40655 7 1 2 40653 40654
0 40656 7 1 2 91027 40655
0 40657 5 1 1 40656
0 40658 7 1 2 40649 40657
0 40659 5 1 1 40658
0 40660 7 1 2 65832 85528
0 40661 7 1 2 40659 40660
0 40662 5 1 1 40661
0 40663 7 1 2 89786 92234
0 40664 5 1 1 40663
0 40665 7 1 2 73887 81596
0 40666 5 1 1 40665
0 40667 7 1 2 40664 40666
0 40668 5 1 1 40667
0 40669 7 1 2 78828 40668
0 40670 5 1 1 40669
0 40671 7 1 2 78199 75036
0 40672 7 1 2 97045 40671
0 40673 5 1 1 40672
0 40674 7 1 2 40670 40673
0 40675 5 1 1 40674
0 40676 7 1 2 101302 40675
0 40677 5 1 1 40676
0 40678 7 1 2 62439 77381
0 40679 7 1 2 100723 40678
0 40680 7 1 2 100731 40679
0 40681 7 1 2 93013 40680
0 40682 5 1 1 40681
0 40683 7 1 2 40677 40682
0 40684 5 1 1 40683
0 40685 7 1 2 72185 40684
0 40686 5 1 1 40685
0 40687 7 1 2 86240 101059
0 40688 5 1 1 40687
0 40689 7 1 2 90936 77283
0 40690 5 1 1 40689
0 40691 7 1 2 40688 40690
0 40692 5 1 1 40691
0 40693 7 1 2 65198 75883
0 40694 7 1 2 40692 40693
0 40695 7 1 2 101303 40694
0 40696 5 1 1 40695
0 40697 7 1 2 40686 40696
0 40698 7 1 2 40662 40697
0 40699 5 1 1 40698
0 40700 7 1 2 65509 40699
0 40701 5 1 1 40700
0 40702 7 1 2 40605 40701
0 40703 5 1 1 40702
0 40704 7 1 2 87363 40703
0 40705 5 1 1 40704
0 40706 7 2 2 64778 82670
0 40707 7 1 2 62885 96307
0 40708 5 1 1 40707
0 40709 7 1 2 72567 101131
0 40710 5 1 1 40709
0 40711 7 1 2 89469 89531
0 40712 5 1 1 40711
0 40713 7 1 2 40710 40712
0 40714 5 1 1 40713
0 40715 7 1 2 82500 40714
0 40716 5 1 1 40715
0 40717 7 1 2 40708 40716
0 40718 5 1 1 40717
0 40719 7 1 2 101304 40718
0 40720 5 1 1 40719
0 40721 7 1 2 88302 81597
0 40722 7 1 2 80479 40721
0 40723 7 1 2 93570 40722
0 40724 5 1 1 40723
0 40725 7 1 2 40720 40724
0 40726 5 1 1 40725
0 40727 7 1 2 64558 40726
0 40728 5 1 1 40727
0 40729 7 1 2 71985 94333
0 40730 5 1 1 40729
0 40731 7 1 2 96290 40730
0 40732 5 1 1 40731
0 40733 7 1 2 68458 40732
0 40734 5 1 1 40733
0 40735 7 1 2 78370 97289
0 40736 5 1 1 40735
0 40737 7 1 2 40734 40736
0 40738 5 1 1 40737
0 40739 7 1 2 67723 40738
0 40740 5 1 1 40739
0 40741 7 1 2 77477 86152
0 40742 5 1 1 40741
0 40743 7 1 2 40740 40742
0 40744 5 1 1 40743
0 40745 7 1 2 67033 40744
0 40746 5 1 1 40745
0 40747 7 1 2 79658 82514
0 40748 7 1 2 96827 40747
0 40749 5 1 1 40748
0 40750 7 1 2 40746 40749
0 40751 5 1 1 40750
0 40752 7 1 2 101203 40751
0 40753 5 1 1 40752
0 40754 7 1 2 40728 40753
0 40755 5 1 1 40754
0 40756 7 1 2 61643 40755
0 40757 5 1 1 40756
0 40758 7 1 2 80654 96772
0 40759 5 1 1 40758
0 40760 7 1 2 74228 81572
0 40761 5 1 1 40760
0 40762 7 1 2 40759 40761
0 40763 5 1 1 40762
0 40764 7 1 2 86022 40763
0 40765 5 1 1 40764
0 40766 7 1 2 89342 96991
0 40767 5 1 1 40766
0 40768 7 1 2 40765 40767
0 40769 5 1 1 40768
0 40770 7 1 2 65833 40769
0 40771 5 1 1 40770
0 40772 7 1 2 71986 94906
0 40773 7 1 2 90421 40772
0 40774 5 1 1 40773
0 40775 7 1 2 40771 40774
0 40776 5 1 1 40775
0 40777 7 1 2 90267 40776
0 40778 5 1 1 40777
0 40779 7 1 2 40757 40778
0 40780 5 1 1 40779
0 40781 7 1 2 70426 40780
0 40782 5 1 1 40781
0 40783 7 1 2 75115 80609
0 40784 7 1 2 87234 40783
0 40785 5 1 1 40784
0 40786 7 1 2 962 17549
0 40787 5 1 1 40786
0 40788 7 1 2 85757 72330
0 40789 7 1 2 40787 40788
0 40790 5 1 1 40789
0 40791 7 1 2 35701 40790
0 40792 5 1 1 40791
0 40793 7 1 2 78936 417
0 40794 7 1 2 40792 40793
0 40795 5 1 1 40794
0 40796 7 1 2 40785 40795
0 40797 5 1 1 40796
0 40798 7 1 2 74821 40797
0 40799 5 1 1 40798
0 40800 7 1 2 69028 85763
0 40801 5 2 1 40800
0 40802 7 1 2 73580 87039
0 40803 5 1 1 40802
0 40804 7 1 2 101306 40803
0 40805 5 1 1 40804
0 40806 7 1 2 81895 95331
0 40807 7 1 2 40805 40806
0 40808 5 1 1 40807
0 40809 7 1 2 40799 40808
0 40810 5 1 1 40809
0 40811 7 1 2 65834 40810
0 40812 5 1 1 40811
0 40813 7 1 2 73488 75884
0 40814 7 1 2 93729 40813
0 40815 7 1 2 75564 40814
0 40816 5 1 1 40815
0 40817 7 1 2 40812 40816
0 40818 5 1 1 40817
0 40819 7 1 2 66531 40818
0 40820 5 1 1 40819
0 40821 7 1 2 85842 75565
0 40822 5 1 1 40821
0 40823 7 1 2 68459 94301
0 40824 5 1 1 40823
0 40825 7 1 2 40822 40824
0 40826 5 1 1 40825
0 40827 7 1 2 67034 40826
0 40828 5 1 1 40827
0 40829 7 1 2 74822 84661
0 40830 7 1 2 93510 40829
0 40831 5 1 1 40830
0 40832 7 1 2 40828 40831
0 40833 5 1 1 40832
0 40834 7 1 2 67504 40833
0 40835 5 1 1 40834
0 40836 7 1 2 68460 76655
0 40837 7 1 2 92364 40836
0 40838 5 1 1 40837
0 40839 7 1 2 40835 40838
0 40840 5 1 1 40839
0 40841 7 1 2 89086 40840
0 40842 5 1 1 40841
0 40843 7 1 2 40820 40842
0 40844 5 1 1 40843
0 40845 7 1 2 68225 40844
0 40846 5 1 1 40845
0 40847 7 1 2 77904 75731
0 40848 5 1 1 40847
0 40849 7 1 2 68872 94302
0 40850 5 1 1 40849
0 40851 7 1 2 40848 40850
0 40852 5 1 1 40851
0 40853 7 1 2 82873 96383
0 40854 7 1 2 40852 40853
0 40855 5 1 1 40854
0 40856 7 1 2 40846 40855
0 40857 5 1 1 40856
0 40858 7 1 2 65510 40857
0 40859 5 1 1 40858
0 40860 7 1 2 66532 77153
0 40861 7 1 2 101200 40860
0 40862 7 1 2 91741 40861
0 40863 5 1 1 40862
0 40864 7 1 2 40859 40863
0 40865 5 1 1 40864
0 40866 7 1 2 69410 40865
0 40867 5 1 1 40866
0 40868 7 1 2 40782 40867
0 40869 5 1 1 40868
0 40870 7 3 2 64290 70125
0 40871 7 1 2 91028 101308
0 40872 7 1 2 40869 40871
0 40873 5 1 1 40872
0 40874 7 1 2 40705 40873
0 40875 7 1 2 40581 40874
0 40876 5 1 1 40875
0 40877 7 1 2 69243 40876
0 40878 5 1 1 40877
0 40879 7 1 2 81896 98741
0 40880 5 1 1 40879
0 40881 7 1 2 81163 81253
0 40882 7 1 2 93581 95282
0 40883 7 1 2 40881 40882
0 40884 7 1 2 98723 40883
0 40885 5 1 1 40884
0 40886 7 1 2 40880 40885
0 40887 5 1 1 40886
0 40888 7 1 2 85128 79536
0 40889 7 1 2 40887 40888
0 40890 5 1 1 40889
0 40891 7 1 2 86176 100358
0 40892 5 1 1 40891
0 40893 7 1 2 74823 98298
0 40894 5 1 1 40893
0 40895 7 1 2 40892 40894
0 40896 5 1 1 40895
0 40897 7 2 2 93686 94592
0 40898 7 1 2 79756 82445
0 40899 7 1 2 97460 40898
0 40900 7 1 2 101311 40899
0 40901 7 1 2 40896 40900
0 40902 5 1 1 40901
0 40903 7 1 2 40890 40902
0 40904 5 1 1 40903
0 40905 7 1 2 61644 40904
0 40906 5 1 1 40905
0 40907 7 2 2 68035 97675
0 40908 7 1 2 95668 101313
0 40909 5 1 1 40908
0 40910 7 1 2 64170 73581
0 40911 5 1 1 40910
0 40912 7 1 2 100352 40911
0 40913 5 13 1 40912
0 40914 7 2 2 64779 101315
0 40915 7 1 2 80610 97991
0 40916 7 1 2 92972 40915
0 40917 7 1 2 101328 40916
0 40918 5 1 1 40917
0 40919 7 1 2 40909 40918
0 40920 5 1 1 40919
0 40921 7 1 2 65835 40920
0 40922 5 1 1 40921
0 40923 7 4 2 93002 93688
0 40924 7 2 2 100791 101330
0 40925 7 1 2 91413 95651
0 40926 7 1 2 101334 40925
0 40927 5 1 1 40926
0 40928 7 1 2 40922 40927
0 40929 5 1 1 40928
0 40930 7 1 2 71987 40929
0 40931 5 1 1 40930
0 40932 7 1 2 95315 99239
0 40933 7 1 2 100402 40932
0 40934 7 1 2 101316 40933
0 40935 5 1 1 40934
0 40936 7 1 2 40931 40935
0 40937 5 1 1 40936
0 40938 7 1 2 90147 40937
0 40939 5 1 1 40938
0 40940 7 1 2 40906 40939
0 40941 5 1 1 40940
0 40942 7 1 2 61309 40941
0 40943 5 1 1 40942
0 40944 7 2 2 76179 100359
0 40945 5 1 1 101336
0 40946 7 1 2 64171 83511
0 40947 5 1 1 40946
0 40948 7 1 2 40945 40947
0 40949 5 1 1 40948
0 40950 7 1 2 80263 40949
0 40951 5 1 1 40950
0 40952 7 1 2 82762 91128
0 40953 5 1 1 40952
0 40954 7 1 2 40951 40953
0 40955 5 1 1 40954
0 40956 7 1 2 86177 40955
0 40957 5 1 1 40956
0 40958 7 2 2 71170 76096
0 40959 5 1 1 101338
0 40960 7 1 2 98290 40959
0 40961 5 1 1 40960
0 40962 7 1 2 81266 91234
0 40963 7 1 2 40961 40962
0 40964 5 1 1 40963
0 40965 7 1 2 40957 40964
0 40966 5 1 1 40965
0 40967 7 1 2 65199 86872
0 40968 7 1 2 40966 40967
0 40969 5 1 1 40968
0 40970 7 1 2 88351 71495
0 40971 7 1 2 81744 40970
0 40972 7 1 2 79389 86199
0 40973 7 1 2 40971 40972
0 40974 5 1 1 40973
0 40975 7 1 2 40969 40974
0 40976 5 1 1 40975
0 40977 7 1 2 97881 40976
0 40978 5 1 1 40977
0 40979 7 1 2 40943 40978
0 40980 5 1 1 40979
0 40981 7 1 2 70427 40980
0 40982 5 1 1 40981
0 40983 7 1 2 97284 101029
0 40984 5 1 1 40983
0 40985 7 1 2 68700 40984
0 40986 5 1 1 40985
0 40987 7 1 2 91338 15935
0 40988 5 1 1 40987
0 40989 7 1 2 63838 40988
0 40990 5 1 1 40989
0 40991 7 1 2 86012 40990
0 40992 5 1 1 40991
0 40993 7 1 2 65836 76097
0 40994 7 1 2 40992 40993
0 40995 5 1 1 40994
0 40996 7 1 2 85970 100877
0 40997 5 1 1 40996
0 40998 7 1 2 65837 75187
0 40999 5 1 1 40998
0 41000 7 1 2 78174 40999
0 41001 5 1 1 41000
0 41002 7 1 2 92372 41001
0 41003 5 1 1 41002
0 41004 7 1 2 40997 41003
0 41005 7 1 2 40995 41004
0 41006 7 1 2 40986 41005
0 41007 5 1 1 41006
0 41008 7 1 2 98247 41007
0 41009 5 1 1 41008
0 41010 7 1 2 80826 82309
0 41011 7 1 2 79321 41010
0 41012 7 1 2 100913 41011
0 41013 5 1 1 41012
0 41014 7 1 2 41009 41013
0 41015 5 1 1 41014
0 41016 7 1 2 89111 98040
0 41017 7 1 2 92474 41016
0 41018 7 1 2 41015 41017
0 41019 5 1 1 41018
0 41020 7 1 2 40982 41019
0 41021 5 1 1 41020
0 41022 7 1 2 64382 41021
0 41023 5 1 1 41022
0 41024 7 2 2 85587 91437
0 41025 5 1 1 101340
0 41026 7 1 2 94010 41025
0 41027 5 1 1 41026
0 41028 7 1 2 81098 41027
0 41029 5 1 1 41028
0 41030 7 1 2 15647 92869
0 41031 5 1 1 41030
0 41032 7 1 2 68701 41031
0 41033 5 1 1 41032
0 41034 7 1 2 94178 41033
0 41035 5 1 1 41034
0 41036 7 1 2 72186 82341
0 41037 7 1 2 41035 41036
0 41038 5 1 1 41037
0 41039 7 1 2 41029 41038
0 41040 5 1 1 41039
0 41041 7 1 2 89112 94736
0 41042 7 1 2 100852 41041
0 41043 7 1 2 41040 41042
0 41044 5 1 1 41043
0 41045 7 1 2 41023 41044
0 41046 5 1 1 41045
0 41047 7 1 2 75165 41046
0 41048 5 1 1 41047
0 41049 7 1 2 40878 41048
0 41050 7 1 2 40307 41049
0 41051 7 1 2 84321 89306
0 41052 5 1 1 41051
0 41053 7 1 2 65838 41052
0 41054 5 1 1 41053
0 41055 7 1 2 72568 90309
0 41056 5 1 1 41055
0 41057 7 1 2 41054 41056
0 41058 5 1 1 41057
0 41059 7 2 2 62618 41058
0 41060 5 1 1 101342
0 41061 7 1 2 63986 94507
0 41062 5 1 1 41061
0 41063 7 2 2 41060 41062
0 41064 5 1 1 101344
0 41065 7 1 2 88089 101345
0 41066 5 1 1 41065
0 41067 7 1 2 100951 41066
0 41068 5 1 1 41067
0 41069 7 2 2 62619 97096
0 41070 5 1 1 101346
0 41071 7 2 2 73966 101347
0 41072 5 1 1 101348
0 41073 7 1 2 39016 41072
0 41074 5 1 1 41073
0 41075 7 1 2 65839 41074
0 41076 5 1 1 41075
0 41077 7 1 2 67296 97762
0 41078 5 1 1 41077
0 41079 7 1 2 41076 41078
0 41080 5 1 1 41079
0 41081 7 1 2 65511 41080
0 41082 5 1 1 41081
0 41083 7 1 2 1043 84904
0 41084 5 1 1 41083
0 41085 7 1 2 89981 41084
0 41086 5 1 1 41085
0 41087 7 1 2 41082 41086
0 41088 5 1 1 41087
0 41089 7 1 2 82342 41088
0 41090 5 1 1 41089
0 41091 7 1 2 41068 41090
0 41092 5 1 1 41091
0 41093 7 1 2 68702 41092
0 41094 5 1 1 41093
0 41095 7 3 2 69411 72278
0 41096 5 1 1 101350
0 41097 7 1 2 101351 100859
0 41098 5 1 1 41097
0 41099 7 1 2 73793 84732
0 41100 5 1 1 41099
0 41101 7 1 2 76744 98299
0 41102 5 2 1 41101
0 41103 7 1 2 19664 101353
0 41104 5 1 1 41103
0 41105 7 1 2 65840 41104
0 41106 5 1 1 41105
0 41107 7 1 2 41100 41106
0 41108 5 1 1 41107
0 41109 7 1 2 81099 41108
0 41110 5 1 1 41109
0 41111 7 1 2 41098 41110
0 41112 5 1 1 41111
0 41113 7 1 2 73993 41112
0 41114 5 1 1 41113
0 41115 7 1 2 41094 41114
0 41116 5 1 1 41115
0 41117 7 1 2 69614 41116
0 41118 5 1 1 41117
0 41119 7 1 2 69412 99463
0 41120 7 1 2 87268 41119
0 41121 7 1 2 97962 41120
0 41122 5 1 1 41121
0 41123 7 1 2 41118 41122
0 41124 5 1 1 41123
0 41125 7 1 2 92475 41124
0 41126 5 1 1 41125
0 41127 7 1 2 68703 101049
0 41128 5 1 1 41127
0 41129 7 1 2 101125 41128
0 41130 5 1 1 41129
0 41131 7 1 2 65841 41130
0 41132 5 1 1 41131
0 41133 7 1 2 84727 41132
0 41134 5 1 1 41133
0 41135 7 1 2 100934 100582
0 41136 7 1 2 41134 41135
0 41137 5 1 1 41136
0 41138 7 1 2 67505 90303
0 41139 5 1 1 41138
0 41140 7 1 2 65842 92368
0 41141 5 1 1 41140
0 41142 7 1 2 41139 41141
0 41143 5 1 1 41142
0 41144 7 1 2 64172 41143
0 41145 5 1 1 41144
0 41146 7 1 2 100953 41145
0 41147 5 1 1 41146
0 41148 7 1 2 63839 41147
0 41149 5 1 1 41148
0 41150 7 1 2 72569 97923
0 41151 5 1 1 41150
0 41152 7 1 2 67297 75732
0 41153 5 2 1 41152
0 41154 7 1 2 72637 91718
0 41155 7 1 2 101355 41154
0 41156 5 1 1 41155
0 41157 7 1 2 68704 41156
0 41158 7 1 2 41151 41157
0 41159 5 1 1 41158
0 41160 7 1 2 41149 41159
0 41161 5 1 1 41160
0 41162 7 1 2 93868 95254
0 41163 7 1 2 41161 41162
0 41164 5 1 1 41163
0 41165 7 1 2 41137 41164
0 41166 5 1 1 41165
0 41167 7 1 2 90779 93804
0 41168 7 1 2 41166 41167
0 41169 5 1 1 41168
0 41170 7 1 2 41126 41169
0 41171 5 1 1 41170
0 41172 7 1 2 69134 41171
0 41173 5 1 1 41172
0 41174 7 1 2 90780 97651
0 41175 7 1 2 100760 41174
0 41176 5 1 1 41175
0 41177 7 1 2 73654 90666
0 41178 7 1 2 81267 41177
0 41179 7 1 2 101072 41178
0 41180 5 1 1 41179
0 41181 7 1 2 41176 41180
0 41182 5 1 1 41181
0 41183 7 1 2 91646 41182
0 41184 5 1 1 41183
0 41185 7 3 2 61388 100274
0 41186 5 4 1 101357
0 41187 7 1 2 98165 101166
0 41188 7 1 2 101358 41187
0 41189 5 1 1 41188
0 41190 7 1 2 41184 41189
0 41191 5 1 1 41190
0 41192 7 1 2 61310 41191
0 41193 5 1 1 41192
0 41194 7 1 2 83306 97787
0 41195 7 1 2 89553 41194
0 41196 7 1 2 85872 41195
0 41197 7 1 2 90718 81268
0 41198 7 1 2 41196 41197
0 41199 5 1 1 41198
0 41200 7 1 2 41193 41199
0 41201 5 1 1 41200
0 41202 7 1 2 71988 41201
0 41203 5 1 1 41202
0 41204 7 2 2 67298 97676
0 41205 5 1 1 101364
0 41206 7 1 2 68705 82723
0 41207 7 1 2 100946 41206
0 41208 7 1 2 101365 41207
0 41209 5 1 1 41208
0 41210 7 1 2 41203 41209
0 41211 7 1 2 41173 41210
0 41212 5 1 1 41211
0 41213 7 1 2 68461 41212
0 41214 5 1 1 41213
0 41215 7 1 2 67724 99651
0 41216 5 1 1 41215
0 41217 7 1 2 99609 41216
0 41218 5 3 1 41217
0 41219 7 1 2 66255 101366
0 41220 5 1 1 41219
0 41221 7 1 2 36401 41220
0 41222 5 4 1 41221
0 41223 7 1 2 93869 101369
0 41224 5 1 1 41223
0 41225 7 1 2 90643 83309
0 41226 5 1 1 41225
0 41227 7 1 2 41224 41226
0 41228 5 1 1 41227
0 41229 7 1 2 91978 41228
0 41230 5 1 1 41229
0 41231 7 1 2 69413 93767
0 41232 5 2 1 41231
0 41233 7 1 2 4594 90634
0 41234 5 1 1 41233
0 41235 7 2 2 101373 41234
0 41236 7 1 2 67810 101375
0 41237 5 1 1 41236
0 41238 7 1 2 35595 41237
0 41239 5 1 1 41238
0 41240 7 1 2 66145 41239
0 41241 5 1 1 41240
0 41242 7 1 2 35604 41241
0 41243 5 1 1 41242
0 41244 7 1 2 100426 41243
0 41245 5 1 1 41244
0 41246 7 1 2 41230 41245
0 41247 5 1 1 41246
0 41248 7 1 2 78010 41247
0 41249 5 1 1 41248
0 41250 7 1 2 80169 99381
0 41251 5 1 1 41250
0 41252 7 1 2 91979 93805
0 41253 5 1 1 41252
0 41254 7 2 2 67877 81475
0 41255 7 1 2 99022 101377
0 41256 5 1 1 41255
0 41257 7 1 2 41253 41256
0 41258 5 1 1 41257
0 41259 7 1 2 66027 41258
0 41260 5 1 1 41259
0 41261 7 1 2 41251 41260
0 41262 5 1 1 41261
0 41263 7 1 2 93870 41262
0 41264 5 1 1 41263
0 41265 7 2 2 90998 91381
0 41266 7 3 2 98106 101379
0 41267 5 1 1 101381
0 41268 7 1 2 80053 101382
0 41269 5 1 1 41268
0 41270 7 1 2 41264 41269
0 41271 5 1 1 41270
0 41272 7 1 2 82286 41271
0 41273 5 1 1 41272
0 41274 7 1 2 41249 41273
0 41275 5 1 1 41274
0 41276 7 1 2 71263 41275
0 41277 5 1 1 41276
0 41278 7 2 2 69615 92476
0 41279 7 1 2 77256 101384
0 41280 5 1 1 41279
0 41281 7 1 2 91980 99045
0 41282 5 1 1 41281
0 41283 7 1 2 41280 41282
0 41284 5 1 1 41283
0 41285 7 1 2 82287 78315
0 41286 7 1 2 41284 41285
0 41287 5 1 1 41286
0 41288 7 1 2 41277 41287
0 41289 5 1 1 41288
0 41290 7 1 2 73489 98041
0 41291 7 1 2 74905 41290
0 41292 7 1 2 41289 41291
0 41293 5 1 1 41292
0 41294 7 1 2 68226 41293
0 41295 7 1 2 41214 41294
0 41296 5 1 1 41295
0 41297 7 1 2 73105 93717
0 41298 5 1 1 41297
0 41299 7 1 2 62620 41298
0 41300 5 1 1 41299
0 41301 7 1 2 65512 97759
0 41302 5 1 1 41301
0 41303 7 1 2 70428 95865
0 41304 5 1 1 41303
0 41305 7 1 2 64173 41304
0 41306 7 1 2 41302 41305
0 41307 5 1 1 41306
0 41308 7 1 2 41300 41307
0 41309 5 1 1 41308
0 41310 7 1 2 97314 41309
0 41311 5 1 1 41310
0 41312 7 1 2 100502 41311
0 41313 5 1 1 41312
0 41314 7 1 2 76098 41313
0 41315 5 1 1 41314
0 41316 7 1 2 100831 101349
0 41317 5 1 1 41316
0 41318 7 1 2 100510 41317
0 41319 7 1 2 41315 41318
0 41320 5 1 1 41319
0 41321 7 1 2 88195 41320
0 41322 5 1 1 41321
0 41323 7 1 2 84637 99328
0 41324 5 1 1 41323
0 41325 7 1 2 98534 41324
0 41326 5 1 1 41325
0 41327 7 1 2 77257 88104
0 41328 7 1 2 41326 41327
0 41329 5 1 1 41328
0 41330 7 1 2 41322 41329
0 41331 5 1 1 41330
0 41332 7 1 2 93806 41331
0 41333 5 1 1 41332
0 41334 7 1 2 88105 96949
0 41335 7 2 2 99406 41334
0 41336 5 1 1 101386
0 41337 7 1 2 92552 101387
0 41338 5 1 1 41337
0 41339 7 1 2 41333 41338
0 41340 5 1 1 41339
0 41341 7 1 2 69414 41340
0 41342 5 1 1 41341
0 41343 7 5 2 88178 99122
0 41344 5 2 1 101388
0 41345 7 1 2 97011 98017
0 41346 5 1 1 41345
0 41347 7 1 2 97689 41346
0 41348 5 1 1 41347
0 41349 7 1 2 72638 41348
0 41350 5 1 1 41349
0 41351 7 1 2 101393 41350
0 41352 5 1 1 41351
0 41353 7 1 2 76099 41352
0 41354 5 1 1 41353
0 41355 7 1 2 99123 99227
0 41356 7 1 2 98758 41355
0 41357 5 1 1 41356
0 41358 7 1 2 41354 41357
0 41359 5 1 1 41358
0 41360 7 1 2 61311 41359
0 41361 5 1 1 41360
0 41362 7 1 2 66533 72639
0 41363 7 1 2 97012 41362
0 41364 7 1 2 99980 41363
0 41365 7 1 2 90719 41364
0 41366 5 1 1 41365
0 41367 7 1 2 41361 41366
0 41368 5 1 1 41367
0 41369 7 1 2 79374 41368
0 41370 5 1 1 41369
0 41371 7 1 2 41342 41370
0 41372 5 1 1 41371
0 41373 7 1 2 63619 41372
0 41374 5 1 1 41373
0 41375 7 2 2 74188 92477
0 41376 7 1 2 77948 87113
0 41377 7 1 2 95426 41376
0 41378 7 2 2 101395 41377
0 41379 7 1 2 86655 93215
0 41380 7 1 2 101397 41379
0 41381 5 1 1 41380
0 41382 7 1 2 41374 41381
0 41383 5 1 1 41382
0 41384 7 1 2 71866 41383
0 41385 5 1 1 41384
0 41386 7 1 2 74891 91489
0 41387 7 1 2 101398 41386
0 41388 5 1 1 41387
0 41389 7 1 2 63391 41388
0 41390 7 1 2 41385 41389
0 41391 5 1 1 41390
0 41392 7 1 2 64383 41391
0 41393 7 1 2 41296 41392
0 41394 5 1 1 41393
0 41395 7 1 2 80071 90667
0 41396 7 1 2 101054 41395
0 41397 5 1 1 41396
0 41398 7 1 2 31935 41397
0 41399 5 1 1 41398
0 41400 7 1 2 69029 41399
0 41401 5 1 1 41400
0 41402 7 1 2 80075 92644
0 41403 7 1 2 98601 41402
0 41404 7 2 2 69135 100286
0 41405 7 1 2 89121 101399
0 41406 7 1 2 41403 41405
0 41407 5 1 1 41406
0 41408 7 1 2 41401 41407
0 41409 5 1 1 41408
0 41410 7 1 2 86977 41409
0 41411 5 1 1 41410
0 41412 7 2 2 80054 100287
0 41413 7 1 2 80733 93582
0 41414 7 1 2 101401 41413
0 41415 7 1 2 101055 41414
0 41416 5 1 1 41415
0 41417 7 1 2 41411 41416
0 41418 5 1 1 41417
0 41419 7 1 2 73129 41418
0 41420 5 1 1 41419
0 41421 7 1 2 81936 79913
0 41422 5 1 1 41421
0 41423 7 1 2 68873 93408
0 41424 5 1 1 41423
0 41425 7 1 2 41422 41424
0 41426 5 1 1 41425
0 41427 7 1 2 65843 41426
0 41428 5 1 1 41427
0 41429 7 1 2 86767 87235
0 41430 5 1 1 41429
0 41431 7 1 2 41428 41430
0 41432 5 1 1 41431
0 41433 7 1 2 70429 41432
0 41434 5 1 1 41433
0 41435 7 1 2 70751 77635
0 41436 7 1 2 94063 41435
0 41437 5 1 1 41436
0 41438 7 1 2 93491 41437
0 41439 5 1 1 41438
0 41440 7 1 2 97057 41439
0 41441 5 1 1 41440
0 41442 7 1 2 41434 41441
0 41443 5 1 1 41442
0 41444 7 1 2 98685 41443
0 41445 5 1 1 41444
0 41446 7 1 2 41420 41445
0 41447 5 1 1 41446
0 41448 7 1 2 68706 41447
0 41449 5 1 1 41448
0 41450 7 2 2 88106 86768
0 41451 5 1 1 101403
0 41452 7 1 2 68874 101404
0 41453 5 1 1 41452
0 41454 7 1 2 73994 91229
0 41455 5 1 1 41454
0 41456 7 1 2 41453 41455
0 41457 5 1 1 41456
0 41458 7 1 2 72187 41457
0 41459 5 1 1 41458
0 41460 7 1 2 90379 99434
0 41461 5 1 1 41460
0 41462 7 1 2 41459 41461
0 41463 5 1 1 41462
0 41464 7 1 2 65844 41463
0 41465 5 1 1 41464
0 41466 7 1 2 94662 101161
0 41467 5 1 1 41466
0 41468 7 1 2 41465 41467
0 41469 5 1 1 41468
0 41470 7 1 2 98686 41469
0 41471 5 1 1 41470
0 41472 7 1 2 41449 41471
0 41473 5 1 1 41472
0 41474 7 1 2 68462 41473
0 41475 5 1 1 41474
0 41476 7 2 2 77861 93010
0 41477 7 1 2 75921 95316
0 41478 7 1 2 100491 98602
0 41479 7 1 2 41477 41478
0 41480 7 1 2 101405 41479
0 41481 5 1 1 41480
0 41482 7 1 2 74917 94770
0 41483 7 1 2 97869 41482
0 41484 7 1 2 91029 41483
0 41485 5 1 1 41484
0 41486 7 1 2 41481 41485
0 41487 5 1 1 41486
0 41488 7 1 2 87364 41487
0 41489 5 1 1 41488
0 41490 7 1 2 65845 81672
0 41491 7 1 2 94737 41490
0 41492 7 1 2 82213 89313
0 41493 7 1 2 41491 41492
0 41494 7 1 2 101263 41493
0 41495 5 1 1 41494
0 41496 7 1 2 41489 41495
0 41497 7 1 2 41475 41496
0 41498 5 1 1 41497
0 41499 7 1 2 68036 41498
0 41500 5 1 1 41499
0 41501 7 1 2 78316 93997
0 41502 5 1 1 41501
0 41503 7 1 2 68463 97860
0 41504 5 1 1 41503
0 41505 7 1 2 41502 41504
0 41506 5 1 1 41505
0 41507 7 1 2 66534 41506
0 41508 7 1 2 97833 41507
0 41509 5 1 1 41508
0 41510 7 1 2 63840 97870
0 41511 5 1 1 41510
0 41512 7 1 2 80901 41511
0 41513 5 1 1 41512
0 41514 7 1 2 73490 41513
0 41515 5 1 1 41514
0 41516 7 1 2 67506 94193
0 41517 5 1 1 41516
0 41518 7 1 2 72071 93489
0 41519 5 1 1 41518
0 41520 7 1 2 4458 41519
0 41521 5 1 1 41520
0 41522 7 1 2 68707 41521
0 41523 5 1 1 41522
0 41524 7 1 2 41517 41523
0 41525 7 1 2 41515 41524
0 41526 5 1 1 41525
0 41527 7 1 2 68464 41526
0 41528 5 1 1 41527
0 41529 7 1 2 82197 92742
0 41530 7 1 2 94039 41529
0 41531 5 1 1 41530
0 41532 7 1 2 41528 41531
0 41533 5 1 1 41532
0 41534 7 1 2 89267 99046
0 41535 7 1 2 41533 41534
0 41536 5 1 1 41535
0 41537 7 1 2 41509 41536
0 41538 5 1 1 41537
0 41539 7 1 2 95153 41538
0 41540 5 1 1 41539
0 41541 7 1 2 41500 41540
0 41542 5 1 1 41541
0 41543 7 1 2 68227 41542
0 41544 5 1 1 41543
0 41545 7 1 2 82504 94081
0 41546 5 1 1 41545
0 41547 7 1 2 77445 41546
0 41548 5 1 1 41547
0 41549 7 1 2 94180 41548
0 41550 5 1 1 41549
0 41551 7 1 2 63841 41550
0 41552 5 1 1 41551
0 41553 7 1 2 94182 41552
0 41554 5 1 1 41553
0 41555 7 1 2 72072 76180
0 41556 7 1 2 41554 41555
0 41557 5 1 1 41556
0 41558 7 1 2 72479 84038
0 41559 5 1 1 41558
0 41560 7 1 2 63842 80414
0 41561 7 1 2 80840 41560
0 41562 7 1 2 41559 41561
0 41563 5 1 1 41562
0 41564 7 1 2 41557 41563
0 41565 5 1 1 41564
0 41566 7 1 2 69616 41565
0 41567 5 1 1 41566
0 41568 7 1 2 90009 83503
0 41569 7 1 2 64174 303
0 41570 5 1 1 41569
0 41571 7 1 2 86506 41570
0 41572 7 1 2 41568 41571
0 41573 5 1 1 41572
0 41574 7 1 2 41567 41573
0 41575 5 1 1 41574
0 41576 7 1 2 99047 41575
0 41577 5 1 1 41576
0 41578 7 1 2 64780 76423
0 41579 7 1 2 86089 41578
0 41580 7 1 2 96897 41579
0 41581 7 1 2 91030 41580
0 41582 5 1 1 41581
0 41583 7 1 2 41577 41582
0 41584 5 1 1 41583
0 41585 7 1 2 95678 41584
0 41586 5 1 1 41585
0 41587 7 1 2 69415 41586
0 41588 7 1 2 41544 41587
0 41589 5 1 1 41588
0 41590 7 1 2 90720 87666
0 41591 5 1 1 41590
0 41592 7 2 2 93807 101137
0 41593 7 1 2 81827 93087
0 41594 7 1 2 101407 41593
0 41595 5 1 1 41594
0 41596 7 1 2 41591 41595
0 41597 5 1 1 41596
0 41598 7 1 2 61645 41597
0 41599 5 1 1 41598
0 41600 7 1 2 83440 97604
0 41601 7 1 2 101408 41600
0 41602 5 1 1 41601
0 41603 7 1 2 41599 41602
0 41604 5 1 1 41603
0 41605 7 1 2 70430 41604
0 41606 5 1 1 41605
0 41607 7 1 2 72570 82884
0 41608 7 1 2 100141 41607
0 41609 7 1 2 92743 41608
0 41610 7 1 2 99382 41609
0 41611 5 1 1 41610
0 41612 7 1 2 41606 41611
0 41613 5 1 1 41612
0 41614 7 1 2 61312 97450
0 41615 7 1 2 41613 41614
0 41616 5 1 1 41615
0 41617 7 1 2 88107 97031
0 41618 7 1 2 98742 41617
0 41619 5 1 1 41618
0 41620 7 1 2 88234 96370
0 41621 5 1 1 41620
0 41622 7 1 2 74130 74494
0 41623 7 1 2 90574 41622
0 41624 5 1 1 41623
0 41625 7 1 2 41621 41624
0 41626 5 1 1 41625
0 41627 7 1 2 62621 41626
0 41628 5 1 1 41627
0 41629 7 1 2 91230 100463
0 41630 5 1 1 41629
0 41631 7 1 2 41628 41630
0 41632 5 1 1 41631
0 41633 7 1 2 66256 98460
0 41634 5 1 1 41633
0 41635 7 2 2 80808 93748
0 41636 7 1 2 91679 101409
0 41637 5 1 1 41636
0 41638 7 1 2 41634 41637
0 41639 5 4 1 41638
0 41640 7 1 2 97992 101411
0 41641 7 1 2 41632 41640
0 41642 5 1 1 41641
0 41643 7 1 2 41619 41642
0 41644 5 1 1 41643
0 41645 7 1 2 66146 41644
0 41646 5 1 1 41645
0 41647 7 1 2 64559 41646
0 41648 7 1 2 41616 41647
0 41649 5 1 1 41648
0 41650 7 1 2 69244 41649
0 41651 7 1 2 41589 41650
0 41652 5 1 1 41651
0 41653 7 1 2 41394 41652
0 41654 5 1 1 41653
0 41655 7 1 2 80573 41654
0 41656 5 1 1 41655
0 41657 7 3 2 77334 83729
0 41658 5 2 1 101415
0 41659 7 1 2 76481 101416
0 41660 5 1 1 41659
0 41661 7 1 2 86621 85540
0 41662 5 1 1 41661
0 41663 7 1 2 63843 41662
0 41664 5 1 1 41663
0 41665 7 2 2 72466 94324
0 41666 5 1 1 101420
0 41667 7 1 2 1526 101233
0 41668 5 1 1 41667
0 41669 7 1 2 41666 41668
0 41670 7 1 2 41664 41669
0 41671 5 1 1 41670
0 41672 7 1 2 70126 41671
0 41673 5 1 1 41672
0 41674 7 1 2 41660 41673
0 41675 5 1 1 41674
0 41676 7 1 2 63620 41675
0 41677 5 1 1 41676
0 41678 7 1 2 79030 75733
0 41679 5 1 1 41678
0 41680 7 1 2 75329 100956
0 41681 5 1 1 41680
0 41682 7 1 2 41679 41681
0 41683 5 1 1 41682
0 41684 7 1 2 62187 41683
0 41685 5 1 1 41684
0 41686 7 1 2 40233 41685
0 41687 5 1 1 41686
0 41688 7 1 2 70431 41687
0 41689 5 1 1 41688
0 41690 7 1 2 41677 41689
0 41691 5 1 1 41690
0 41692 7 1 2 63392 41691
0 41693 5 1 1 41692
0 41694 7 5 2 71352 85114
0 41695 5 1 1 101422
0 41696 7 1 2 77154 95748
0 41697 7 1 2 101423 41696
0 41698 5 1 1 41697
0 41699 7 1 2 41693 41698
0 41700 5 1 1 41699
0 41701 7 1 2 99592 41700
0 41702 5 1 1 41701
0 41703 7 2 2 68228 90810
0 41704 5 1 1 101427
0 41705 7 1 2 41704 101118
0 41706 5 1 1 41705
0 41707 7 1 2 62188 41706
0 41708 5 1 1 41707
0 41709 7 2 2 90487 86656
0 41710 7 1 2 71867 101429
0 41711 5 1 1 41710
0 41712 7 1 2 41708 41711
0 41713 5 1 1 41712
0 41714 7 3 2 95362 41713
0 41715 7 1 2 99578 101431
0 41716 5 1 1 41715
0 41717 7 1 2 41702 41716
0 41718 5 1 1 41717
0 41719 7 1 2 77258 41718
0 41720 5 1 1 41719
0 41721 7 1 2 87407 92553
0 41722 7 1 2 101432 41721
0 41723 5 1 1 41722
0 41724 7 1 2 41720 41723
0 41725 5 1 1 41724
0 41726 7 1 2 61389 41725
0 41727 5 1 1 41726
0 41728 7 1 2 92102 93760
0 41729 7 1 2 101433 41728
0 41730 5 1 1 41729
0 41731 7 1 2 41727 41730
0 41732 5 1 1 41731
0 41733 7 1 2 64384 41732
0 41734 5 1 1 41733
0 41735 7 1 2 66257 100673
0 41736 5 1 1 41735
0 41737 7 3 2 80988 93749
0 41738 5 1 1 101434
0 41739 7 1 2 41736 41738
0 41740 5 13 1 41739
0 41741 7 1 2 90918 93949
0 41742 7 1 2 97453 41741
0 41743 7 1 2 101113 41742
0 41744 7 1 2 101437 41743
0 41745 5 1 1 41744
0 41746 7 1 2 41734 41745
0 41747 5 1 1 41746
0 41748 7 1 2 62978 41747
0 41749 5 1 1 41748
0 41750 7 1 2 79610 75860
0 41751 7 1 2 99305 41750
0 41752 7 4 2 98107 99203
0 41753 7 1 2 96765 101450
0 41754 7 1 2 41751 41753
0 41755 7 1 2 101114 41754
0 41756 5 1 1 41755
0 41757 7 1 2 41749 41756
0 41758 5 1 1 41757
0 41759 7 1 2 97451 41758
0 41760 5 1 1 41759
0 41761 7 2 2 70752 92175
0 41762 5 1 1 101454
0 41763 7 1 2 93616 41762
0 41764 5 1 1 41763
0 41765 7 1 2 90613 41764
0 41766 5 1 1 41765
0 41767 7 1 2 90953 87840
0 41768 5 1 1 41767
0 41769 7 1 2 41766 41768
0 41770 5 1 1 41769
0 41771 7 1 2 88800 99124
0 41772 7 1 2 41770 41771
0 41773 5 1 1 41772
0 41774 7 3 2 67811 95317
0 41775 7 1 2 66258 99007
0 41776 7 1 2 101456 41775
0 41777 7 1 2 98916 41776
0 41778 5 1 1 41777
0 41779 7 1 2 41773 41778
0 41780 5 1 1 41779
0 41781 7 1 2 63987 41780
0 41782 5 1 1 41781
0 41783 7 3 2 71742 93601
0 41784 5 1 1 101459
0 41785 7 1 2 63844 98615
0 41786 7 1 2 101460 41785
0 41787 7 1 2 98764 41786
0 41788 5 1 1 41787
0 41789 7 1 2 41782 41788
0 41790 5 1 1 41789
0 41791 7 1 2 62622 41790
0 41792 5 1 1 41791
0 41793 7 1 2 68229 80394
0 41794 5 1 1 41793
0 41795 7 2 2 61390 100118
0 41796 7 2 2 97652 101462
0 41797 7 1 2 63393 92518
0 41798 5 1 1 41797
0 41799 7 1 2 101464 41798
0 41800 7 1 2 41794 41799
0 41801 5 1 1 41800
0 41802 7 1 2 41792 41801
0 41803 5 1 1 41802
0 41804 7 1 2 63621 41803
0 41805 5 1 1 41804
0 41806 7 1 2 64385 100497
0 41807 7 3 2 83730 41806
0 41808 7 1 2 91344 87299
0 41809 7 1 2 101466 41808
0 41810 5 1 1 41809
0 41811 7 1 2 41805 41810
0 41812 5 1 1 41811
0 41813 7 1 2 62189 41812
0 41814 5 1 1 41813
0 41815 7 1 2 85129 98580
0 41816 7 1 2 97677 41815
0 41817 7 1 2 101164 41816
0 41818 5 1 1 41817
0 41819 7 1 2 41814 41818
0 41820 5 1 1 41819
0 41821 7 1 2 92541 41820
0 41822 5 1 1 41821
0 41823 7 1 2 67035 77306
0 41824 5 2 1 41823
0 41825 7 1 2 76217 100966
0 41826 5 2 1 41825
0 41827 7 1 2 62190 101471
0 41828 5 1 1 41827
0 41829 7 1 2 101469 41828
0 41830 5 1 1 41829
0 41831 7 1 2 75965 41830
0 41832 5 1 1 41831
0 41833 7 1 2 86634 82489
0 41834 5 1 1 41833
0 41835 7 1 2 41832 41834
0 41836 5 1 1 41835
0 41837 7 1 2 100073 41836
0 41838 5 1 1 41837
0 41839 7 1 2 94069 98613
0 41840 7 1 2 94217 41839
0 41841 5 1 1 41840
0 41842 7 1 2 41838 41841
0 41843 5 1 1 41842
0 41844 7 1 2 99414 41843
0 41845 5 1 1 41844
0 41846 7 1 2 97422 98728
0 41847 7 1 2 98204 41846
0 41848 5 1 1 41847
0 41849 7 3 2 63622 92176
0 41850 5 1 1 101473
0 41851 7 1 2 41784 41850
0 41852 5 1 1 41851
0 41853 7 1 2 90614 41852
0 41854 5 1 1 41853
0 41855 7 1 2 90954 93697
0 41856 5 1 1 41855
0 41857 7 1 2 41854 41856
0 41858 5 1 1 41857
0 41859 7 1 2 64291 71353
0 41860 7 1 2 41858 41859
0 41861 5 1 1 41860
0 41862 7 1 2 41848 41861
0 41863 5 1 1 41862
0 41864 7 1 2 71868 41863
0 41865 5 1 1 41864
0 41866 7 1 2 90615 100142
0 41867 7 1 2 101467 41866
0 41868 5 1 1 41867
0 41869 7 1 2 41865 41868
0 41870 5 1 1 41869
0 41871 7 1 2 62191 41870
0 41872 5 1 1 41871
0 41873 7 1 2 91345 74292
0 41874 7 1 2 101468 41873
0 41875 5 1 1 41874
0 41876 7 1 2 41872 41875
0 41877 5 1 1 41876
0 41878 7 1 2 82671 41877
0 41879 5 1 1 41878
0 41880 7 1 2 41845 41879
0 41881 5 1 1 41880
0 41882 7 1 2 65200 41881
0 41883 5 1 1 41882
0 41884 7 1 2 66535 41883
0 41885 7 1 2 41822 41884
0 41886 5 1 1 41885
0 41887 7 2 2 62192 79514
0 41888 5 2 1 101476
0 41889 7 1 2 90927 101478
0 41890 5 1 1 41889
0 41891 7 1 2 83681 74229
0 41892 5 2 1 41891
0 41893 7 1 2 41890 101480
0 41894 5 1 1 41893
0 41895 7 1 2 71989 41894
0 41896 5 1 1 41895
0 41897 7 1 2 89601 79304
0 41898 5 1 1 41897
0 41899 7 1 2 41896 41898
0 41900 5 1 1 41899
0 41901 7 1 2 65513 41900
0 41902 5 1 1 41901
0 41903 7 2 2 98975 101229
0 41904 5 1 1 101482
0 41905 7 1 2 81312 4169
0 41906 5 1 1 41905
0 41907 7 1 2 5048 41906
0 41908 7 1 2 96314 41907
0 41909 5 1 1 41908
0 41910 7 1 2 41904 41909
0 41911 5 1 1 41910
0 41912 7 1 2 83783 41911
0 41913 5 1 1 41912
0 41914 7 1 2 41902 41913
0 41915 5 1 1 41914
0 41916 7 1 2 93602 41915
0 41917 5 1 1 41916
0 41918 7 1 2 71597 97854
0 41919 5 1 1 41918
0 41920 7 2 2 62623 77915
0 41921 7 1 2 101484 98274
0 41922 5 1 1 41921
0 41923 7 1 2 41919 41922
0 41924 5 1 1 41923
0 41925 7 1 2 65201 41924
0 41926 5 1 1 41925
0 41927 7 1 2 80678 94061
0 41928 7 1 2 98944 41927
0 41929 5 1 1 41928
0 41930 7 1 2 41926 41929
0 41931 5 2 1 41930
0 41932 7 1 2 92177 101486
0 41933 5 1 1 41932
0 41934 7 1 2 41917 41933
0 41935 5 1 1 41934
0 41936 7 1 2 90616 41935
0 41937 5 1 1 41936
0 41938 7 1 2 98358 101487
0 41939 5 1 1 41938
0 41940 7 1 2 41937 41939
0 41941 5 1 1 41940
0 41942 7 1 2 63623 41941
0 41943 5 1 1 41942
0 41944 7 1 2 89634 98271
0 41945 5 1 1 41944
0 41946 7 1 2 79719 82490
0 41947 5 1 1 41946
0 41948 7 1 2 98353 41947
0 41949 5 1 1 41948
0 41950 7 1 2 81778 41949
0 41951 5 1 1 41950
0 41952 7 1 2 41945 41951
0 41953 5 1 1 41952
0 41954 7 1 2 100154 41953
0 41955 5 1 1 41954
0 41956 7 1 2 101424 98275
0 41957 5 1 1 41956
0 41958 7 1 2 75579 91332
0 41959 7 1 2 87958 41958
0 41960 5 1 1 41959
0 41961 7 1 2 41957 41960
0 41962 5 1 1 41961
0 41963 7 1 2 71869 100162
0 41964 7 1 2 41962 41963
0 41965 5 1 1 41964
0 41966 7 1 2 41955 41965
0 41967 5 1 1 41966
0 41968 7 1 2 65202 41967
0 41969 5 1 1 41968
0 41970 7 1 2 75734 83619
0 41971 5 1 1 41970
0 41972 7 1 2 99187 41971
0 41973 5 1 1 41972
0 41974 7 1 2 79611 81745
0 41975 7 1 2 100163 41974
0 41976 7 1 2 41973 41975
0 41977 5 1 1 41976
0 41978 7 1 2 41969 41977
0 41979 7 1 2 41943 41978
0 41980 5 1 1 41979
0 41981 7 1 2 64292 41980
0 41982 5 1 1 41981
0 41983 7 1 2 74230 101483
0 41984 5 1 1 41983
0 41985 7 1 2 67036 90928
0 41986 5 1 1 41985
0 41987 7 1 2 101481 41986
0 41988 5 1 1 41987
0 41989 7 1 2 65514 93358
0 41990 7 1 2 41988 41989
0 41991 5 1 1 41990
0 41992 7 1 2 41984 41991
0 41993 5 1 1 41992
0 41994 7 1 2 97461 99628
0 41995 7 1 2 98511 41994
0 41996 7 1 2 41993 41995
0 41997 5 1 1 41996
0 41998 7 1 2 65846 89726
0 41999 7 1 2 76624 41998
0 42000 7 1 2 94505 99189
0 42001 7 1 2 98861 42000
0 42002 7 1 2 41999 42001
0 42003 5 1 1 42002
0 42004 7 1 2 61646 42003
0 42005 7 1 2 41997 42004
0 42006 7 1 2 41982 42005
0 42007 5 1 1 42006
0 42008 7 1 2 64560 42007
0 42009 7 1 2 41886 42008
0 42010 5 1 1 42009
0 42011 7 1 2 77624 81598
0 42012 5 1 1 42011
0 42013 7 1 2 101119 42012
0 42014 5 1 1 42013
0 42015 7 1 2 70127 76181
0 42016 7 1 2 42014 42015
0 42017 5 1 1 42016
0 42018 7 1 2 91144 96527
0 42019 7 1 2 97185 42018
0 42020 5 1 1 42019
0 42021 7 1 2 42017 42020
0 42022 5 1 1 42021
0 42023 7 1 2 93603 42022
0 42024 5 1 1 42023
0 42025 7 1 2 76058 75200
0 42026 7 1 2 83550 42025
0 42027 7 1 2 79869 101474
0 42028 7 1 2 42026 42027
0 42029 5 1 1 42028
0 42030 7 1 2 42024 42029
0 42031 5 1 1 42030
0 42032 7 1 2 62193 42031
0 42033 5 1 1 42032
0 42034 7 1 2 77925 93155
0 42035 7 1 2 93661 42034
0 42036 7 1 2 97032 42035
0 42037 5 1 1 42036
0 42038 7 1 2 42033 42037
0 42039 5 1 1 42038
0 42040 7 2 2 64293 100736
0 42041 7 1 2 99097 101488
0 42042 7 1 2 42039 42041
0 42043 5 1 1 42042
0 42044 7 1 2 42010 42043
0 42045 5 1 1 42044
0 42046 7 1 2 69617 42045
0 42047 5 1 1 42046
0 42048 7 1 2 61313 42047
0 42049 7 1 2 41760 42048
0 42050 5 1 1 42049
0 42051 7 1 2 64386 89939
0 42052 7 1 2 91193 97370
0 42053 7 1 2 42051 42052
0 42054 7 1 2 100981 42053
0 42055 5 1 1 42054
0 42056 7 1 2 77578 94343
0 42057 7 1 2 97000 100184
0 42058 7 1 2 42056 42057
0 42059 5 1 1 42058
0 42060 7 1 2 42055 42059
0 42061 5 1 1 42060
0 42062 7 1 2 68465 42061
0 42063 5 1 1 42062
0 42064 7 1 2 66536 78796
0 42065 7 1 2 100143 42064
0 42066 7 1 2 92275 98442
0 42067 7 1 2 42065 42066
0 42068 5 1 1 42067
0 42069 7 1 2 42063 42068
0 42070 5 1 1 42069
0 42071 7 1 2 65203 95427
0 42072 7 1 2 42070 42071
0 42073 5 1 1 42072
0 42074 7 1 2 83559 93698
0 42075 7 1 2 90014 42074
0 42076 7 2 2 77131 79544
0 42077 7 1 2 99179 101490
0 42078 7 1 2 42075 42077
0 42079 5 1 1 42078
0 42080 7 1 2 42073 42079
0 42081 5 1 1 42080
0 42082 7 1 2 93808 42081
0 42083 5 1 1 42082
0 42084 7 2 2 93912 99453
0 42085 7 1 2 77307 90542
0 42086 7 3 2 101492 42085
0 42087 7 1 2 80679 100104
0 42088 7 1 2 101494 42087
0 42089 5 1 1 42088
0 42090 7 1 2 42083 42089
0 42091 5 1 1 42090
0 42092 7 1 2 68037 42091
0 42093 5 1 1 42092
0 42094 7 2 2 90721 98512
0 42095 7 1 2 65515 99182
0 42096 5 1 1 42095
0 42097 7 1 2 95589 42096
0 42098 5 1 1 42097
0 42099 7 1 2 101497 42098
0 42100 5 1 1 42099
0 42101 7 1 2 91346 93913
0 42102 7 1 2 99004 42101
0 42103 5 1 1 42102
0 42104 7 1 2 42100 42103
0 42105 5 1 1 42104
0 42106 7 1 2 67037 42105
0 42107 5 1 1 42106
0 42108 7 1 2 82493 100967
0 42109 5 1 1 42108
0 42110 7 3 2 90982 100123
0 42111 7 1 2 75966 93914
0 42112 7 1 2 101499 42111
0 42113 7 1 2 42109 42112
0 42114 5 1 1 42113
0 42115 7 1 2 42107 42114
0 42116 5 1 1 42115
0 42117 7 1 2 87071 42116
0 42118 5 1 1 42117
0 42119 7 1 2 61391 88269
0 42120 7 1 2 101495 42119
0 42121 5 1 1 42120
0 42122 7 1 2 42118 42121
0 42123 5 1 1 42122
0 42124 7 1 2 61647 42123
0 42125 5 1 1 42124
0 42126 7 1 2 92195 101491
0 42127 7 1 2 101496 42126
0 42128 5 1 1 42127
0 42129 7 1 2 42125 42128
0 42130 5 1 1 42129
0 42131 7 1 2 83819 42130
0 42132 5 1 1 42131
0 42133 7 1 2 42093 42132
0 42134 5 1 1 42133
0 42135 7 1 2 68230 42134
0 42136 5 1 1 42135
0 42137 7 1 2 76182 95534
0 42138 5 1 1 42137
0 42139 7 1 2 76059 76897
0 42140 7 1 2 85971 42139
0 42141 5 1 1 42140
0 42142 7 1 2 42138 42141
0 42143 5 1 1 42142
0 42144 7 1 2 101498 42143
0 42145 5 1 1 42144
0 42146 7 1 2 70753 76060
0 42147 7 1 2 89903 42146
0 42148 5 1 1 42147
0 42149 7 1 2 71870 95079
0 42150 5 1 1 42149
0 42151 7 1 2 42148 42150
0 42152 5 1 1 42151
0 42153 7 1 2 100634 97678
0 42154 7 1 2 42152 42153
0 42155 5 1 1 42154
0 42156 7 1 2 42145 42155
0 42157 5 1 1 42156
0 42158 7 1 2 69618 42157
0 42159 5 1 1 42158
0 42160 7 1 2 79757 93062
0 42161 7 1 2 99090 42160
0 42162 7 2 2 66259 77259
0 42163 5 1 1 101502
0 42164 7 2 2 99579 98180
0 42165 7 1 2 94344 101504
0 42166 7 1 2 101503 42165
0 42167 7 1 2 42161 42166
0 42168 5 1 1 42167
0 42169 7 1 2 42159 42168
0 42170 5 1 1 42169
0 42171 7 1 2 63624 42170
0 42172 5 1 1 42171
0 42173 7 1 2 87072 88069
0 42174 5 1 1 42173
0 42175 7 1 2 83594 98791
0 42176 5 1 1 42175
0 42177 7 1 2 42174 42176
0 42178 5 1 1 42177
0 42179 7 1 2 80384 99204
0 42180 7 1 2 101493 42179
0 42181 7 1 2 42178 42180
0 42182 5 1 1 42181
0 42183 7 1 2 42172 42182
0 42184 5 1 1 42183
0 42185 7 1 2 97878 42184
0 42186 5 1 1 42185
0 42187 7 1 2 66147 42186
0 42188 7 1 2 42136 42187
0 42189 5 1 1 42188
0 42190 7 1 2 72640 42189
0 42191 7 1 2 42050 42190
0 42192 5 1 1 42191
0 42193 7 1 2 41656 42192
0 42194 7 1 2 41050 42193
0 42195 7 1 2 39065 42194
0 42196 7 1 2 37575 42195
0 42197 5 1 1 42196
0 42198 7 1 2 100224 42197
0 42199 5 1 1 42198
0 42200 7 1 2 35481 42199
0 42201 7 1 2 31475 42200
0 42202 7 3 2 83764 77364
0 42203 5 7 1 101506
0 42204 7 2 2 62624 90359
0 42205 5 1 1 101516
0 42206 7 1 2 92417 101317
0 42207 5 1 1 42206
0 42208 7 1 2 42205 42207
0 42209 5 2 1 42208
0 42210 7 1 2 75056 101518
0 42211 5 1 1 42210
0 42212 7 1 2 75016 87535
0 42213 5 1 1 42212
0 42214 7 1 2 42211 42213
0 42215 5 1 1 42214
0 42216 7 1 2 63845 42215
0 42217 5 1 1 42216
0 42218 7 1 2 73717 86006
0 42219 7 1 2 90361 42218
0 42220 5 1 1 42219
0 42221 7 1 2 42217 42220
0 42222 5 1 1 42221
0 42223 7 1 2 99652 42222
0 42224 5 1 1 42223
0 42225 7 2 2 82243 94456
0 42226 7 1 2 75188 98995
0 42227 7 1 2 101520 42226
0 42228 5 1 1 42227
0 42229 7 1 2 42224 42228
0 42230 5 1 1 42229
0 42231 7 1 2 66260 42230
0 42232 5 1 1 42231
0 42233 7 1 2 93750 95385
0 42234 7 1 2 101521 42233
0 42235 5 1 1 42234
0 42236 7 1 2 42232 42235
0 42237 5 1 1 42236
0 42238 7 1 2 92901 42237
0 42239 5 1 1 42238
0 42240 7 3 2 69416 98731
0 42241 7 1 2 96791 101522
0 42242 5 1 1 42241
0 42243 7 1 2 88984 9555
0 42244 5 8 1 42243
0 42245 7 2 2 69417 101318
0 42246 7 1 2 100792 101533
0 42247 5 1 1 42246
0 42248 7 1 2 72571 99483
0 42249 5 1 1 42248
0 42250 7 1 2 42247 42249
0 42251 5 1 1 42250
0 42252 7 1 2 101525 42251
0 42253 5 1 1 42252
0 42254 7 1 2 81212 87171
0 42255 7 1 2 101523 42254
0 42256 5 1 1 42255
0 42257 7 1 2 42253 42256
0 42258 5 1 1 42257
0 42259 7 1 2 63846 42258
0 42260 5 1 1 42259
0 42261 7 1 2 42242 42260
0 42262 5 1 1 42261
0 42263 7 1 2 66769 42262
0 42264 5 1 1 42263
0 42265 7 1 2 76850 90906
0 42266 7 1 2 98088 42265
0 42267 7 1 2 85195 42266
0 42268 5 1 1 42267
0 42269 7 1 2 42264 42268
0 42270 5 1 1 42269
0 42271 7 1 2 68038 42270
0 42272 5 1 1 42271
0 42273 7 3 2 82381 80117
0 42274 7 1 2 66261 79860
0 42275 7 1 2 88734 42274
0 42276 7 1 2 101535 42275
0 42277 5 1 1 42276
0 42278 7 1 2 42272 42277
0 42279 5 1 1 42278
0 42280 7 1 2 65516 42279
0 42281 5 1 1 42280
0 42282 7 6 2 83372 72734
0 42283 5 1 1 101538
0 42284 7 1 2 100902 42283
0 42285 5 7 1 42284
0 42286 7 3 2 70432 101544
0 42287 7 2 2 69827 81828
0 42288 7 1 2 84437 91810
0 42289 7 1 2 101554 42288
0 42290 7 1 2 101551 42289
0 42291 5 1 1 42290
0 42292 7 1 2 42281 42291
0 42293 5 1 1 42292
0 42294 7 1 2 70128 42293
0 42295 5 1 1 42294
0 42296 7 1 2 66262 89338
0 42297 7 1 2 89766 42296
0 42298 7 1 2 92307 42297
0 42299 5 1 1 42298
0 42300 7 1 2 42295 42299
0 42301 5 1 1 42300
0 42302 7 1 2 68466 42301
0 42303 5 1 1 42302
0 42304 7 1 2 89806 13451
0 42305 5 3 1 42304
0 42306 7 2 2 81829 92290
0 42307 7 3 2 73700 86044
0 42308 7 1 2 98732 101561
0 42309 7 1 2 101559 42308
0 42310 7 1 2 101556 42309
0 42311 5 1 1 42310
0 42312 7 1 2 42303 42311
0 42313 5 1 1 42312
0 42314 7 1 2 67878 42313
0 42315 5 1 1 42314
0 42316 7 1 2 66263 97397
0 42317 7 1 2 86544 42316
0 42318 7 2 2 63847 84058
0 42319 7 1 2 91827 101564
0 42320 7 1 2 42317 42319
0 42321 5 1 1 42320
0 42322 7 1 2 42315 42321
0 42323 5 1 1 42322
0 42324 7 1 2 61648 42323
0 42325 5 1 1 42324
0 42326 7 1 2 42239 42325
0 42327 5 1 1 42326
0 42328 7 1 2 64781 42327
0 42329 5 1 1 42328
0 42330 7 1 2 89822 99998
0 42331 5 1 1 42330
0 42332 7 1 2 42331 101360
0 42333 5 1 1 42332
0 42334 7 1 2 67507 42333
0 42335 5 1 1 42334
0 42336 7 1 2 70954 82288
0 42337 7 1 2 98129 42336
0 42338 5 2 1 42337
0 42339 7 1 2 42335 101566
0 42340 5 2 1 42339
0 42341 7 1 2 80711 101568
0 42342 5 1 1 42341
0 42343 7 4 2 72839 90445
0 42344 7 1 2 99484 101570
0 42345 5 1 1 42344
0 42346 7 1 2 67508 72840
0 42347 5 5 1 42346
0 42348 7 1 2 85288 99999
0 42349 7 1 2 101574 42348
0 42350 5 1 1 42349
0 42351 7 1 2 42345 42350
0 42352 5 1 1 42351
0 42353 7 1 2 91705 42352
0 42354 5 1 1 42353
0 42355 7 1 2 42342 42354
0 42356 5 1 1 42355
0 42357 7 1 2 67879 42356
0 42358 5 1 1 42357
0 42359 7 1 2 63625 91282
0 42360 7 2 2 101545 42359
0 42361 7 1 2 93761 101579
0 42362 5 1 1 42361
0 42363 7 1 2 42358 42362
0 42364 5 1 1 42363
0 42365 7 1 2 80989 42364
0 42366 5 1 1 42365
0 42367 7 1 2 101580 99470
0 42368 5 1 1 42367
0 42369 7 1 2 42366 42368
0 42370 5 1 1 42369
0 42371 7 1 2 100225 42370
0 42372 5 1 1 42371
0 42373 7 1 2 80990 98381
0 42374 7 1 2 86539 42373
0 42375 7 1 2 101569 42374
0 42376 5 1 1 42375
0 42377 7 1 2 42372 42376
0 42378 5 1 1 42377
0 42379 7 1 2 68231 42378
0 42380 5 1 1 42379
0 42381 7 3 2 64561 101539
0 42382 7 3 2 92196 98495
0 42383 7 1 2 101581 101584
0 42384 5 1 1 42383
0 42385 7 4 2 61392 76562
0 42386 7 2 2 100896 101587
0 42387 7 1 2 93056 101591
0 42388 5 1 1 42387
0 42389 7 1 2 42384 42388
0 42390 5 1 1 42389
0 42391 7 1 2 78715 42390
0 42392 5 1 1 42391
0 42393 7 2 2 66537 97398
0 42394 7 2 2 78716 101593
0 42395 5 1 1 101595
0 42396 7 1 2 67880 95880
0 42397 5 1 1 42396
0 42398 7 1 2 42395 42397
0 42399 5 1 1 42398
0 42400 7 1 2 82289 42399
0 42401 5 1 1 42400
0 42402 7 1 2 76563 99580
0 42403 7 1 2 89877 42402
0 42404 5 1 1 42403
0 42405 7 1 2 42401 42404
0 42406 5 1 1 42405
0 42407 7 1 2 98300 42406
0 42408 5 1 1 42407
0 42409 7 1 2 95875 101582
0 42410 5 1 1 42409
0 42411 7 1 2 83820 82005
0 42412 7 1 2 101540 42411
0 42413 5 1 1 42412
0 42414 7 2 2 64970 94023
0 42415 7 1 2 84232 81658
0 42416 7 1 2 101597 42415
0 42417 5 1 1 42416
0 42418 7 1 2 42413 42417
0 42419 5 1 1 42418
0 42420 7 1 2 66538 42419
0 42421 5 1 1 42420
0 42422 7 1 2 42410 42421
0 42423 5 1 1 42422
0 42424 7 1 2 67881 42423
0 42425 5 1 1 42424
0 42426 7 1 2 101583 101596
0 42427 5 1 1 42426
0 42428 7 1 2 42425 42427
0 42429 7 1 2 42408 42428
0 42430 5 1 1 42429
0 42431 7 1 2 66264 42430
0 42432 5 1 1 42431
0 42433 7 1 2 42392 42432
0 42434 5 1 1 42433
0 42435 7 1 2 83432 42434
0 42436 5 1 1 42435
0 42437 7 1 2 69619 42436
0 42438 7 1 2 42380 42437
0 42439 5 1 1 42438
0 42440 7 3 2 79244 74507
0 42441 5 10 1 101599
0 42442 7 1 2 67725 101602
0 42443 5 1 1 42442
0 42444 7 1 2 84669 86736
0 42445 5 1 1 42444
0 42446 7 1 2 42443 42445
0 42447 5 3 1 42446
0 42448 7 1 2 99653 101612
0 42449 5 1 1 42448
0 42450 7 2 2 63032 69030
0 42451 7 2 2 88735 101615
0 42452 5 2 1 101617
0 42453 7 1 2 42449 101619
0 42454 5 1 1 42453
0 42455 7 1 2 66265 42454
0 42456 5 1 1 42455
0 42457 7 1 2 72572 100549
0 42458 5 1 1 42457
0 42459 7 1 2 42456 42458
0 42460 5 1 1 42459
0 42461 7 1 2 66770 101526
0 42462 5 1 1 42461
0 42463 7 1 2 96762 42462
0 42464 5 3 1 42463
0 42465 7 1 2 76183 101621
0 42466 5 1 1 42465
0 42467 7 2 2 69828 82382
0 42468 7 1 2 80991 101624
0 42469 5 1 1 42468
0 42470 7 1 2 42466 42469
0 42471 5 1 1 42470
0 42472 7 1 2 42460 42471
0 42473 5 1 1 42472
0 42474 7 2 2 83834 72573
0 42475 7 1 2 90668 101625
0 42476 7 1 2 101626 42475
0 42477 5 1 1 42476
0 42478 7 1 2 42473 42477
0 42479 5 1 1 42478
0 42480 7 1 2 80712 42479
0 42481 5 1 1 42480
0 42482 7 3 2 62625 75532
0 42483 5 2 1 101628
0 42484 7 3 2 67509 75547
0 42485 5 1 1 101633
0 42486 7 1 2 101631 42485
0 42487 5 2 1 42486
0 42488 7 1 2 69031 101636
0 42489 5 1 1 42488
0 42490 7 2 2 73582 79240
0 42491 5 2 1 101638
0 42492 7 1 2 42489 101640
0 42493 5 2 1 42492
0 42494 7 1 2 71064 101642
0 42495 5 1 1 42494
0 42496 7 1 2 71006 101637
0 42497 5 1 1 42496
0 42498 7 1 2 42495 42497
0 42499 5 1 1 42498
0 42500 7 1 2 100000 42499
0 42501 5 1 1 42500
0 42502 7 1 2 84106 99485
0 42503 5 1 1 42502
0 42504 7 1 2 42501 42503
0 42505 5 1 1 42504
0 42506 7 1 2 70129 99106
0 42507 7 1 2 91828 42506
0 42508 7 1 2 42505 42507
0 42509 5 1 1 42508
0 42510 7 1 2 64782 42509
0 42511 7 1 2 42481 42510
0 42512 5 1 1 42511
0 42513 7 1 2 74548 42512
0 42514 7 1 2 42439 42513
0 42515 5 1 1 42514
0 42516 7 1 2 90037 92072
0 42517 5 1 1 42516
0 42518 7 1 2 79861 79551
0 42519 5 1 1 42518
0 42520 7 1 2 42517 42519
0 42521 5 1 1 42520
0 42522 7 1 2 63626 42521
0 42523 5 1 1 42522
0 42524 7 1 2 83631 90109
0 42525 5 1 1 42524
0 42526 7 1 2 42523 42525
0 42527 5 1 1 42526
0 42528 7 3 2 92347 100288
0 42529 7 1 2 42527 101644
0 42530 5 1 1 42529
0 42531 7 1 2 78479 98996
0 42532 7 1 2 94457 42531
0 42533 7 1 2 101565 42532
0 42534 5 1 1 42533
0 42535 7 1 2 42530 42534
0 42536 5 1 1 42535
0 42537 7 1 2 76184 42536
0 42538 5 1 1 42537
0 42539 7 2 2 83260 92968
0 42540 5 1 1 101647
0 42541 7 1 2 75548 101648
0 42542 5 1 1 42541
0 42543 7 1 2 91112 28290
0 42544 5 6 1 42543
0 42545 7 2 2 79375 101649
0 42546 7 1 2 92554 101655
0 42547 5 1 1 42546
0 42548 7 1 2 42542 42547
0 42549 5 1 1 42548
0 42550 7 1 2 69032 42549
0 42551 5 1 1 42550
0 42552 7 3 2 79376 92555
0 42553 5 1 1 101657
0 42554 7 1 2 70955 101658
0 42555 5 1 1 42554
0 42556 7 2 2 67882 85898
0 42557 5 1 1 101660
0 42558 7 1 2 64783 88858
0 42559 7 1 2 101661 42558
0 42560 5 1 1 42559
0 42561 7 1 2 42555 42560
0 42562 5 1 1 42561
0 42563 7 1 2 67510 42562
0 42564 5 1 1 42563
0 42565 7 1 2 67726 84766
0 42566 5 2 1 42565
0 42567 7 1 2 101600 101662
0 42568 5 1 1 42567
0 42569 7 1 2 42568 101659
0 42570 5 1 1 42569
0 42571 7 1 2 83261 93003
0 42572 7 1 2 101603 42571
0 42573 5 1 1 42572
0 42574 7 1 2 42570 42573
0 42575 7 1 2 42564 42574
0 42576 7 1 2 42551 42575
0 42577 5 1 1 42576
0 42578 7 1 2 66539 42577
0 42579 5 1 1 42578
0 42580 7 2 2 84897 94499
0 42581 5 1 1 101664
0 42582 7 1 2 100903 101601
0 42583 7 1 2 101665 42582
0 42584 5 1 1 42583
0 42585 7 5 2 69620 99107
0 42586 7 1 2 83821 101666
0 42587 7 1 2 42584 42586
0 42588 5 1 1 42587
0 42589 7 1 2 42579 42588
0 42590 5 1 1 42589
0 42591 7 1 2 73995 86540
0 42592 7 1 2 42590 42591
0 42593 5 1 1 42592
0 42594 7 1 2 42538 42593
0 42595 5 1 1 42594
0 42596 7 1 2 66266 42595
0 42597 5 1 1 42596
0 42598 7 3 2 67883 92197
0 42599 7 2 2 100388 101671
0 42600 7 2 2 63197 73996
0 42601 7 1 2 83213 95992
0 42602 7 1 2 101676 42601
0 42603 7 1 2 101674 42602
0 42604 5 1 1 42603
0 42605 7 1 2 42597 42604
0 42606 5 1 1 42605
0 42607 7 1 2 83142 42606
0 42608 5 1 1 42607
0 42609 7 1 2 67884 91307
0 42610 5 1 1 42609
0 42611 7 2 2 87345 92556
0 42612 5 1 1 101678
0 42613 7 1 2 42610 42612
0 42614 5 1 1 42613
0 42615 7 1 2 42614 98721
0 42616 5 1 1 42615
0 42617 7 1 2 88975 98474
0 42618 7 1 2 101588 42617
0 42619 5 1 1 42618
0 42620 7 1 2 42616 42619
0 42621 5 1 1 42620
0 42622 7 1 2 101546 42621
0 42623 5 1 1 42622
0 42624 7 2 2 72641 85289
0 42625 7 1 2 101555 101585
0 42626 7 1 2 101680 42625
0 42627 5 1 1 42626
0 42628 7 1 2 42623 42627
0 42629 5 1 1 42628
0 42630 7 1 2 64562 42629
0 42631 5 1 1 42630
0 42632 7 1 2 89823 101527
0 42633 5 1 1 42632
0 42634 7 1 2 88927 81213
0 42635 5 1 1 42634
0 42636 7 1 2 42633 42635
0 42637 5 1 1 42636
0 42638 7 1 2 67511 42637
0 42639 5 1 1 42638
0 42640 7 1 2 90411 96688
0 42641 5 1 1 42640
0 42642 7 1 2 42639 42641
0 42643 5 1 1 42642
0 42644 7 1 2 87263 100202
0 42645 7 1 2 42643 42644
0 42646 5 1 1 42645
0 42647 7 1 2 42631 42646
0 42648 5 1 1 42647
0 42649 7 1 2 76898 96372
0 42650 7 1 2 42648 42649
0 42651 5 1 1 42650
0 42652 7 1 2 42608 42651
0 42653 7 1 2 42515 42652
0 42654 7 1 2 42329 42653
0 42655 5 1 1 42654
0 42656 7 1 2 96401 42655
0 42657 5 1 1 42656
0 42658 7 3 2 63033 93128
0 42659 5 2 1 101682
0 42660 7 1 2 101190 101683
0 42661 5 1 1 42660
0 42662 7 1 2 96148 101645
0 42663 5 1 1 42662
0 42664 7 1 2 42661 42663
0 42665 5 1 1 42664
0 42666 7 1 2 74710 82471
0 42667 7 1 2 42665 42666
0 42668 5 1 1 42667
0 42669 7 1 2 93418 100635
0 42670 5 1 1 42669
0 42671 7 1 2 76975 96930
0 42672 5 1 1 42671
0 42673 7 1 2 42670 42672
0 42674 5 1 1 42673
0 42675 7 1 2 101547 98382
0 42676 7 1 2 42674 42675
0 42677 5 1 1 42676
0 42678 7 1 2 42668 42677
0 42679 5 1 1 42678
0 42680 7 1 2 81937 42679
0 42681 5 1 1 42680
0 42682 7 1 2 68467 76976
0 42683 5 1 1 42682
0 42684 7 1 2 63627 89770
0 42685 5 1 1 42684
0 42686 7 1 2 42683 42685
0 42687 5 4 1 42686
0 42688 7 1 2 91322 98383
0 42689 7 1 2 96787 42688
0 42690 7 1 2 101687 42689
0 42691 5 1 1 42690
0 42692 7 1 2 42681 42691
0 42693 5 1 1 42692
0 42694 7 1 2 66267 42693
0 42695 5 1 1 42694
0 42696 7 1 2 76296 80631
0 42697 7 1 2 98594 42696
0 42698 7 2 2 64387 99275
0 42699 7 1 2 101247 101691
0 42700 7 1 2 42697 42699
0 42701 5 1 1 42700
0 42702 7 1 2 42695 42701
0 42703 5 1 1 42702
0 42704 7 1 2 63394 42703
0 42705 5 1 1 42704
0 42706 7 1 2 66028 101675
0 42707 5 1 1 42706
0 42708 7 7 2 66540 63034
0 42709 7 3 2 96853 101693
0 42710 5 1 1 101700
0 42711 7 1 2 64563 101701
0 42712 5 1 1 42711
0 42713 7 1 2 90268 101634
0 42714 5 1 1 42713
0 42715 7 1 2 61649 101656
0 42716 5 1 1 42715
0 42717 7 1 2 42714 42716
0 42718 5 1 1 42717
0 42719 7 1 2 69033 42718
0 42720 5 1 1 42719
0 42721 7 1 2 91506 101604
0 42722 5 1 1 42721
0 42723 7 1 2 84898 101663
0 42724 5 2 1 42723
0 42725 7 1 2 83961 101703
0 42726 5 1 1 42725
0 42727 7 1 2 90553 92597
0 42728 5 1 1 42727
0 42729 7 1 2 42726 42728
0 42730 7 1 2 42722 42729
0 42731 7 1 2 42720 42730
0 42732 5 1 1 42731
0 42733 7 1 2 67885 42732
0 42734 5 1 1 42733
0 42735 7 1 2 42712 42734
0 42736 5 1 1 42735
0 42737 7 1 2 66268 42736
0 42738 5 1 1 42737
0 42739 7 1 2 42707 42738
0 42740 5 1 1 42739
0 42741 7 1 2 101688 42740
0 42742 5 1 1 42741
0 42743 7 1 2 68468 74549
0 42744 7 3 2 79467 42743
0 42745 7 1 2 91876 101646
0 42746 7 1 2 101705 42745
0 42747 5 1 1 42746
0 42748 7 1 2 42742 42747
0 42749 5 1 1 42748
0 42750 7 1 2 66771 42749
0 42751 5 1 1 42750
0 42752 7 1 2 77949 84438
0 42753 7 1 2 93452 42752
0 42754 7 2 2 70956 100217
0 42755 7 1 2 100054 101708
0 42756 7 1 2 42753 42755
0 42757 5 1 1 42756
0 42758 7 1 2 42751 42757
0 42759 5 1 1 42758
0 42760 7 1 2 96832 42759
0 42761 5 1 1 42760
0 42762 7 1 2 42705 42761
0 42763 5 1 1 42762
0 42764 7 1 2 63198 42763
0 42765 5 1 1 42764
0 42766 7 2 2 98733 99581
0 42767 7 2 2 72073 101710
0 42768 7 1 2 87703 101706
0 42769 5 1 1 42768
0 42770 7 1 2 78243 100061
0 42771 7 1 2 88262 42770
0 42772 5 1 1 42771
0 42773 7 1 2 42769 42772
0 42774 5 1 1 42773
0 42775 7 1 2 101712 42774
0 42776 5 1 1 42775
0 42777 7 1 2 87211 86879
0 42778 5 1 1 42777
0 42779 7 1 2 75597 84149
0 42780 5 1 1 42779
0 42781 7 1 2 42778 42780
0 42782 5 1 1 42781
0 42783 7 1 2 61650 42782
0 42784 5 1 1 42783
0 42785 7 3 2 66772 86933
0 42786 7 2 2 68232 101714
0 42787 5 1 1 101717
0 42788 7 1 2 91593 42787
0 42789 5 1 1 42788
0 42790 7 2 2 66541 42789
0 42791 5 1 1 101719
0 42792 7 1 2 81878 101720
0 42793 5 1 1 42792
0 42794 7 1 2 42784 42793
0 42795 5 1 1 42794
0 42796 7 1 2 67886 42795
0 42797 5 1 1 42796
0 42798 7 2 2 94718 99409
0 42799 7 2 2 82746 101721
0 42800 5 1 1 101723
0 42801 7 1 2 67727 101724
0 42802 5 1 1 42801
0 42803 7 1 2 42797 42802
0 42804 5 1 1 42803
0 42805 7 1 2 66269 42804
0 42806 5 1 1 42805
0 42807 7 2 2 101589 99678
0 42808 7 1 2 67728 101725
0 42809 5 1 1 42808
0 42810 7 1 2 42806 42809
0 42811 5 1 1 42810
0 42812 7 1 2 98301 42811
0 42813 5 1 1 42812
0 42814 7 1 2 77205 93004
0 42815 7 1 2 97914 42814
0 42816 5 1 1 42815
0 42817 7 1 2 42800 42816
0 42818 5 1 1 42817
0 42819 7 1 2 101605 42818
0 42820 5 1 1 42819
0 42821 7 1 2 70957 100523
0 42822 5 1 1 42821
0 42823 7 1 2 89347 42822
0 42824 7 1 2 100525 42823
0 42825 5 1 1 42824
0 42826 7 1 2 90907 93005
0 42827 5 1 1 42826
0 42828 7 1 2 100530 42827
0 42829 5 1 1 42828
0 42830 7 1 2 81374 75585
0 42831 7 1 2 42829 42830
0 42832 5 1 1 42831
0 42833 7 1 2 42825 42832
0 42834 5 1 1 42833
0 42835 7 1 2 69034 42834
0 42836 5 1 1 42835
0 42837 7 1 2 86309 93006
0 42838 5 1 1 42837
0 42839 7 1 2 99610 42838
0 42840 5 1 1 42839
0 42841 7 2 2 80246 42840
0 42842 7 1 2 84217 101727
0 42843 5 1 1 42842
0 42844 7 1 2 66542 42843
0 42845 7 1 2 42836 42844
0 42846 5 1 1 42845
0 42847 7 1 2 75686 84150
0 42848 5 1 1 42847
0 42849 7 3 2 84126 86033
0 42850 5 1 1 101729
0 42851 7 1 2 42848 42850
0 42852 5 1 1 42851
0 42853 7 1 2 101606 42852
0 42854 5 1 1 42853
0 42855 7 2 2 69035 84151
0 42856 7 1 2 90078 101732
0 42857 5 1 1 42856
0 42858 7 1 2 42581 101730
0 42859 5 1 1 42858
0 42860 7 1 2 42857 42859
0 42861 7 1 2 42854 42860
0 42862 5 1 1 42861
0 42863 7 1 2 67887 42862
0 42864 5 1 1 42863
0 42865 7 1 2 83388 99593
0 42866 7 1 2 94799 42865
0 42867 5 1 1 42866
0 42868 7 1 2 61651 42867
0 42869 7 1 2 42864 42868
0 42870 5 1 1 42869
0 42871 7 1 2 42846 42870
0 42872 5 1 1 42871
0 42873 7 1 2 42820 42872
0 42874 5 1 1 42873
0 42875 7 1 2 66270 42874
0 42876 5 1 1 42875
0 42877 7 1 2 101607 101726
0 42878 5 1 1 42877
0 42879 7 1 2 15651 42791
0 42880 5 1 1 42879
0 42881 7 1 2 72574 42880
0 42882 5 1 1 42881
0 42883 7 1 2 84218 93218
0 42884 5 1 1 42883
0 42885 7 1 2 42882 42884
0 42886 5 1 1 42885
0 42887 7 1 2 100550 42886
0 42888 5 1 1 42887
0 42889 7 1 2 42878 42888
0 42890 7 1 2 42876 42889
0 42891 7 1 2 42813 42890
0 42892 5 1 1 42891
0 42893 7 1 2 101689 42892
0 42894 5 1 1 42893
0 42895 7 1 2 42776 42894
0 42896 5 1 1 42895
0 42897 7 1 2 96195 42896
0 42898 5 1 1 42897
0 42899 7 1 2 42765 42898
0 42900 5 1 1 42899
0 42901 7 1 2 69829 42900
0 42902 5 1 1 42901
0 42903 7 2 2 66543 88369
0 42904 5 1 1 101734
0 42905 7 1 2 81879 101735
0 42906 5 1 1 42905
0 42907 7 1 2 101172 42906
0 42908 5 1 1 42907
0 42909 7 1 2 67888 42908
0 42910 5 1 1 42909
0 42911 7 2 2 89000 101694
0 42912 7 1 2 78780 101736
0 42913 5 1 1 42912
0 42914 7 1 2 42910 42913
0 42915 5 1 1 42914
0 42916 7 1 2 66271 42915
0 42917 5 1 1 42916
0 42918 7 1 2 80992 78781
0 42919 7 1 2 100551 42918
0 42920 5 1 1 42919
0 42921 7 1 2 42917 42920
0 42922 5 1 1 42921
0 42923 7 1 2 98302 42922
0 42924 5 1 1 42923
0 42925 7 1 2 71131 84000
0 42926 5 1 1 42925
0 42927 7 1 2 79377 91454
0 42928 5 1 1 42927
0 42929 7 1 2 42926 42928
0 42930 5 1 1 42929
0 42931 7 1 2 67512 42930
0 42932 5 1 1 42931
0 42933 7 1 2 89241 80060
0 42934 5 1 1 42933
0 42935 7 1 2 42932 42934
0 42936 5 1 1 42935
0 42937 7 1 2 67889 42936
0 42938 5 1 1 42937
0 42939 7 1 2 68039 101616
0 42940 7 1 2 92130 42939
0 42941 5 1 1 42940
0 42942 7 1 2 61652 42941
0 42943 7 1 2 42938 42942
0 42944 5 1 1 42943
0 42945 7 1 2 80427 99594
0 42946 5 1 1 42945
0 42947 7 1 2 42540 42946
0 42948 5 1 1 42947
0 42949 7 1 2 62886 42948
0 42950 5 1 1 42949
0 42951 7 1 2 83234 100779
0 42952 5 1 1 42951
0 42953 7 1 2 64784 100607
0 42954 5 1 1 42953
0 42955 7 1 2 42952 42954
0 42956 5 1 1 42955
0 42957 7 1 2 66029 42956
0 42958 5 1 1 42957
0 42959 7 1 2 42950 42958
0 42960 5 1 1 42959
0 42961 7 1 2 69036 42960
0 42962 5 1 1 42961
0 42963 7 1 2 81521 101728
0 42964 5 1 1 42963
0 42965 7 1 2 66544 42964
0 42966 7 1 2 42962 42965
0 42967 5 1 1 42966
0 42968 7 1 2 66272 42967
0 42969 7 1 2 42944 42968
0 42970 5 1 1 42969
0 42971 7 1 2 67890 83264
0 42972 5 1 1 42971
0 42973 7 1 2 95255 99410
0 42974 5 1 1 42973
0 42975 7 1 2 42972 42974
0 42976 5 1 1 42975
0 42977 7 1 2 66273 42976
0 42978 5 1 1 42977
0 42979 7 1 2 98475 100041
0 42980 5 1 1 42979
0 42981 7 1 2 42978 42980
0 42982 5 1 1 42981
0 42983 7 1 2 101608 42982
0 42984 5 1 1 42983
0 42985 7 1 2 89092 42904
0 42986 5 1 1 42985
0 42987 7 1 2 72575 42986
0 42988 5 1 1 42987
0 42989 7 1 2 81673 91164
0 42990 5 1 1 42989
0 42991 7 1 2 42988 42990
0 42992 5 1 1 42991
0 42993 7 1 2 100552 42992
0 42994 5 1 1 42993
0 42995 7 1 2 42984 42994
0 42996 7 1 2 42970 42995
0 42997 7 1 2 42924 42996
0 42998 5 1 1 42997
0 42999 7 1 2 101690 42998
0 43000 5 1 1 42999
0 43001 7 1 2 76185 101713
0 43002 7 1 2 101707 43001
0 43003 5 1 1 43002
0 43004 7 1 2 43000 43003
0 43005 5 1 1 43004
0 43006 7 1 2 83143 43005
0 43007 5 1 1 43006
0 43008 7 1 2 86310 74892
0 43009 7 1 2 93244 43008
0 43010 7 1 2 101711 43009
0 43011 7 1 2 92908 43010
0 43012 5 1 1 43011
0 43013 7 1 2 43007 43012
0 43014 5 1 1 43013
0 43015 7 1 2 96451 43014
0 43016 5 1 1 43015
0 43017 7 1 2 42902 43016
0 43018 5 1 1 43017
0 43019 7 1 2 62440 43018
0 43020 5 1 1 43019
0 43021 7 1 2 67038 43020
0 43022 7 1 2 42657 43021
0 43023 5 1 1 43022
0 43024 7 1 2 85683 85694
0 43025 5 1 1 43024
0 43026 7 1 2 74550 82198
0 43027 5 1 1 43026
0 43028 7 1 2 43025 43027
0 43029 5 1 1 43028
0 43030 7 1 2 72718 101667
0 43031 5 1 1 43030
0 43032 7 1 2 100082 43031
0 43033 5 1 1 43032
0 43034 7 1 2 66274 43033
0 43035 5 1 1 43034
0 43036 7 2 2 92198 98852
0 43037 5 3 1 101738
0 43038 7 1 2 43035 101740
0 43039 5 1 1 43038
0 43040 7 1 2 66030 43039
0 43041 5 1 1 43040
0 43042 7 2 2 66275 80794
0 43043 7 1 2 101709 101743
0 43044 5 1 1 43043
0 43045 7 1 2 43041 43044
0 43046 5 1 1 43045
0 43047 7 1 2 69037 43046
0 43048 5 2 1 43047
0 43049 7 1 2 101744 101402
0 43050 5 1 1 43049
0 43051 7 1 2 101745 43050
0 43052 5 1 1 43051
0 43053 7 1 2 90197 43052
0 43054 5 1 1 43053
0 43055 7 1 2 94419 100904
0 43056 5 3 1 43055
0 43057 7 1 2 81938 101747
0 43058 5 1 1 43057
0 43059 7 1 2 43058 101242
0 43060 5 1 1 43059
0 43061 7 1 2 98562 43060
0 43062 5 1 1 43061
0 43063 7 1 2 43054 43062
0 43064 5 1 1 43063
0 43065 7 1 2 64971 43064
0 43066 5 1 1 43065
0 43067 7 1 2 71695 90669
0 43068 7 1 2 101571 43067
0 43069 7 1 2 96806 43068
0 43070 5 1 1 43069
0 43071 7 1 2 43066 43070
0 43072 5 1 1 43071
0 43073 7 1 2 43029 43072
0 43074 5 1 1 43073
0 43075 7 2 2 83144 74664
0 43076 7 1 2 79058 101750
0 43077 5 1 1 43076
0 43078 7 2 2 74869 86530
0 43079 7 1 2 83145 101752
0 43080 7 1 2 101748 43079
0 43081 5 1 1 43080
0 43082 7 1 2 43077 43081
0 43083 5 1 1 43082
0 43084 7 2 2 64785 101438
0 43085 7 1 2 43083 101754
0 43086 5 1 1 43085
0 43087 7 2 2 76253 74441
0 43088 5 2 1 101756
0 43089 7 1 2 77950 84760
0 43090 5 1 1 43089
0 43091 7 1 2 101758 43090
0 43092 5 1 1 43091
0 43093 7 1 2 79214 100561
0 43094 7 1 2 92620 43093
0 43095 7 1 2 43092 43094
0 43096 5 1 1 43095
0 43097 7 1 2 43086 43096
0 43098 5 1 1 43097
0 43099 7 1 2 69830 43098
0 43100 5 1 1 43099
0 43101 7 1 2 43074 43100
0 43102 5 1 1 43101
0 43103 7 1 2 69245 43102
0 43104 5 1 1 43103
0 43105 7 1 2 79112 20302
0 43106 5 1 1 43105
0 43107 7 3 2 4705 43106
0 43108 7 1 2 101439 101760
0 43109 5 1 1 43108
0 43110 7 1 2 88976 100562
0 43111 7 1 2 83867 43110
0 43112 5 1 1 43111
0 43113 7 1 2 43109 43112
0 43114 5 1 1 43113
0 43115 7 1 2 101753 43114
0 43116 5 1 1 43115
0 43117 7 1 2 61904 101528
0 43118 5 1 1 43117
0 43119 7 1 2 17744 43118
0 43120 5 2 1 43119
0 43121 7 1 2 76186 101763
0 43122 5 1 1 43121
0 43123 7 1 2 96019 43122
0 43124 5 1 1 43123
0 43125 7 1 2 67891 43124
0 43126 5 1 1 43125
0 43127 7 1 2 64972 101679
0 43128 5 1 1 43127
0 43129 7 1 2 43126 43128
0 43130 5 1 1 43129
0 43131 7 1 2 66276 43130
0 43132 5 1 1 43131
0 43133 7 2 2 85645 91811
0 43134 7 1 2 98503 101765
0 43135 5 1 1 43134
0 43136 7 1 2 43132 43135
0 43137 5 1 1 43136
0 43138 7 1 2 90784 43137
0 43139 5 1 1 43138
0 43140 7 1 2 43116 43139
0 43141 5 1 1 43140
0 43142 7 1 2 93063 43141
0 43143 5 1 1 43142
0 43144 7 2 2 63199 87481
0 43145 7 2 2 90617 101767
0 43146 7 1 2 80513 76433
0 43147 7 1 2 96910 43146
0 43148 7 1 2 101769 43147
0 43149 5 1 1 43148
0 43150 7 1 2 43143 43149
0 43151 5 1 1 43150
0 43152 7 1 2 72642 43151
0 43153 5 1 1 43152
0 43154 7 1 2 61393 83293
0 43155 7 1 2 91587 43154
0 43156 7 3 2 63035 64175
0 43157 7 2 2 90962 101771
0 43158 7 1 2 97510 101774
0 43159 7 1 2 43155 43158
0 43160 5 1 1 43159
0 43161 7 1 2 70130 43160
0 43162 7 1 2 43153 43161
0 43163 7 1 2 43104 43162
0 43164 5 1 1 43163
0 43165 7 1 2 96854 99383
0 43166 5 1 1 43165
0 43167 7 1 2 69621 101548
0 43168 7 1 2 101440 43167
0 43169 5 1 1 43168
0 43170 7 1 2 43166 43169
0 43171 5 1 1 43170
0 43172 7 1 2 76804 43171
0 43173 5 1 1 43172
0 43174 7 1 2 81939 101549
0 43175 5 1 1 43174
0 43176 7 1 2 101243 43175
0 43177 5 3 1 43176
0 43178 7 1 2 89982 101410
0 43179 7 1 2 101776 43178
0 43180 5 1 1 43179
0 43181 7 1 2 43173 43180
0 43182 5 1 1 43181
0 43183 7 1 2 68233 100226
0 43184 7 1 2 43182 43183
0 43185 5 1 1 43184
0 43186 7 3 2 72643 85764
0 43187 7 1 2 101779 100219
0 43188 5 1 1 43187
0 43189 7 1 2 101746 43188
0 43190 5 1 1 43189
0 43191 7 1 2 87256 43190
0 43192 5 1 1 43191
0 43193 7 1 2 66277 98500
0 43194 5 1 1 43193
0 43195 7 1 2 91812 98504
0 43196 5 1 1 43195
0 43197 7 1 2 43194 43196
0 43198 5 1 1 43197
0 43199 7 1 2 101777 43198
0 43200 5 1 1 43199
0 43201 7 1 2 43192 43200
0 43202 5 1 1 43201
0 43203 7 1 2 63395 76805
0 43204 7 1 2 43202 43203
0 43205 5 1 1 43204
0 43206 7 1 2 43185 43205
0 43207 5 1 1 43206
0 43208 7 1 2 96926 43207
0 43209 5 1 1 43208
0 43210 7 1 2 88486 81382
0 43211 7 2 2 61394 78519
0 43212 7 1 2 101775 101782
0 43213 7 1 2 43210 43212
0 43214 5 1 1 43213
0 43215 7 1 2 65204 43214
0 43216 7 1 2 43209 43215
0 43217 5 1 1 43216
0 43218 7 1 2 43164 43217
0 43219 5 1 1 43218
0 43220 7 1 2 64564 43219
0 43221 5 1 1 43220
0 43222 7 1 2 78962 101629
0 43223 5 1 1 43222
0 43224 7 1 2 66031 83772
0 43225 5 1 1 43224
0 43226 7 1 2 67513 43225
0 43227 7 1 2 88370 43226
0 43228 5 1 1 43227
0 43229 7 1 2 43223 43228
0 43230 5 1 1 43229
0 43231 7 1 2 69038 43230
0 43232 5 1 1 43231
0 43233 7 1 2 66032 88371
0 43234 5 1 1 43233
0 43235 7 1 2 78902 13862
0 43236 5 2 1 43235
0 43237 7 1 2 67729 101784
0 43238 5 1 1 43237
0 43239 7 1 2 43234 43238
0 43240 5 1 1 43239
0 43241 7 1 2 79241 43240
0 43242 5 1 1 43241
0 43243 7 1 2 43232 43242
0 43244 5 1 1 43243
0 43245 7 1 2 66545 43244
0 43246 5 1 1 43245
0 43247 7 1 2 89087 101613
0 43248 5 1 1 43247
0 43249 7 1 2 43246 43248
0 43250 5 1 1 43249
0 43251 7 1 2 95656 43250
0 43252 5 1 1 43251
0 43253 7 1 2 63628 78971
0 43254 7 1 2 75017 43253
0 43255 7 1 2 95482 43254
0 43256 5 1 1 43255
0 43257 7 1 2 43252 43256
0 43258 5 1 1 43257
0 43259 7 1 2 101529 43258
0 43260 5 1 1 43259
0 43261 7 1 2 74628 90462
0 43262 5 1 1 43261
0 43263 7 1 2 73855 101562
0 43264 5 1 1 43263
0 43265 7 1 2 43262 43264
0 43266 5 1 1 43265
0 43267 7 1 2 62626 43266
0 43268 5 1 1 43267
0 43269 7 3 2 90324 101319
0 43270 7 1 2 79780 101786
0 43271 5 1 1 43270
0 43272 7 1 2 43268 43271
0 43273 5 1 1 43272
0 43274 7 1 2 76102 81429
0 43275 5 1 1 43274
0 43276 7 1 2 64786 43275
0 43277 7 1 2 30223 43276
0 43278 7 1 2 43273 43277
0 43279 5 1 1 43278
0 43280 7 1 2 67514 100987
0 43281 5 1 1 43280
0 43282 7 4 2 72576 71677
0 43283 5 2 1 101789
0 43284 7 1 2 43281 101793
0 43285 5 5 1 43284
0 43286 7 2 2 99862 101795
0 43287 7 1 2 77206 91829
0 43288 7 1 2 101800 43287
0 43289 5 1 1 43288
0 43290 7 1 2 43279 43289
0 43291 7 1 2 43260 43290
0 43292 5 1 1 43291
0 43293 7 1 2 73031 43292
0 43294 5 1 1 43293
0 43295 7 2 2 88235 101796
0 43296 5 1 1 101802
0 43297 7 2 2 86380 101320
0 43298 5 1 1 101804
0 43299 7 3 2 62627 74753
0 43300 5 1 1 101806
0 43301 7 1 2 43298 43300
0 43302 5 2 1 43301
0 43303 7 1 2 86978 101809
0 43304 5 1 1 43303
0 43305 7 1 2 43296 43304
0 43306 5 1 1 43305
0 43307 7 1 2 91968 100227
0 43308 7 1 2 43306 43307
0 43309 5 1 1 43308
0 43310 7 1 2 43294 43309
0 43311 5 1 1 43310
0 43312 7 1 2 90670 100636
0 43313 7 1 2 43311 43312
0 43314 5 1 1 43313
0 43315 7 1 2 74908 74056
0 43316 5 4 1 43315
0 43317 7 5 2 67730 76597
0 43318 5 1 1 101815
0 43319 7 1 2 88469 99384
0 43320 5 1 1 43319
0 43321 7 1 2 88255 80672
0 43322 7 1 2 92631 43321
0 43323 5 1 1 43322
0 43324 7 1 2 43320 43323
0 43325 5 1 1 43324
0 43326 7 1 2 101816 43325
0 43327 5 1 1 43326
0 43328 7 2 2 80993 100803
0 43329 7 2 2 64176 101820
0 43330 7 1 2 62887 91362
0 43331 7 1 2 97973 43330
0 43332 7 1 2 101822 43331
0 43333 5 1 1 43332
0 43334 7 1 2 43327 43333
0 43335 5 1 1 43334
0 43336 7 1 2 87309 43335
0 43337 5 1 1 43336
0 43338 7 1 2 91255 101803
0 43339 5 1 1 43338
0 43340 7 1 2 64787 92909
0 43341 7 1 2 101810 43340
0 43342 5 1 1 43341
0 43343 7 1 2 43339 43342
0 43344 5 1 1 43343
0 43345 7 1 2 90671 96452
0 43346 7 1 2 43344 43345
0 43347 5 1 1 43346
0 43348 7 1 2 43337 43347
0 43349 5 1 1 43348
0 43350 7 1 2 101811 43349
0 43351 5 1 1 43350
0 43352 7 2 2 73032 92632
0 43353 7 1 2 62628 100321
0 43354 5 1 1 43353
0 43355 7 1 2 63629 101787
0 43356 5 1 1 43355
0 43357 7 1 2 43354 43356
0 43358 5 1 1 43357
0 43359 7 1 2 64973 92910
0 43360 7 1 2 43358 43359
0 43361 5 1 1 43360
0 43362 7 1 2 81011 101751
0 43363 7 1 2 101614 43362
0 43364 5 1 1 43363
0 43365 7 1 2 43361 43364
0 43366 5 1 1 43365
0 43367 7 1 2 64788 43366
0 43368 5 1 1 43367
0 43369 7 1 2 81599 87264
0 43370 7 1 2 101801 43369
0 43371 5 1 1 43370
0 43372 7 1 2 43368 43371
0 43373 5 1 1 43372
0 43374 7 1 2 101824 43373
0 43375 5 1 1 43374
0 43376 7 1 2 43351 43375
0 43377 5 1 1 43376
0 43378 7 1 2 70131 43377
0 43379 5 1 1 43378
0 43380 7 1 2 69418 43379
0 43381 7 1 2 43314 43380
0 43382 5 1 1 43381
0 43383 7 1 2 43221 43382
0 43384 5 1 1 43383
0 43385 7 1 2 62194 43384
0 43386 5 1 1 43385
0 43387 7 1 2 97315 43386
0 43388 7 1 2 43023 43387
0 43389 5 1 1 43388
0 43390 7 1 2 75255 92348
0 43391 7 1 2 90832 43390
0 43392 5 1 1 43391
0 43393 7 1 2 65517 85765
0 43394 7 1 2 95982 43393
0 43395 5 1 1 43394
0 43396 7 1 2 43392 43395
0 43397 5 1 1 43396
0 43398 7 1 2 64565 43397
0 43399 5 1 1 43398
0 43400 7 1 2 87895 100944
0 43401 7 1 2 97693 43400
0 43402 5 1 1 43401
0 43403 7 1 2 43399 43402
0 43404 5 1 1 43403
0 43405 7 1 2 64177 43404
0 43406 5 1 1 43405
0 43407 7 1 2 62629 88430
0 43408 5 1 1 43407
0 43409 7 1 2 16654 43408
0 43410 5 1 1 43409
0 43411 7 2 2 67039 74086
0 43412 7 1 2 79938 101826
0 43413 7 1 2 43410 43412
0 43414 5 1 1 43413
0 43415 7 1 2 43406 43414
0 43416 5 1 1 43415
0 43417 7 1 2 67299 43416
0 43418 5 1 1 43417
0 43419 7 1 2 82608 86796
0 43420 7 1 2 96795 43419
0 43421 5 1 1 43420
0 43422 7 1 2 43418 43421
0 43423 5 1 1 43422
0 43424 7 1 2 68708 43423
0 43425 5 1 1 43424
0 43426 7 1 2 73869 100452
0 43427 5 2 1 43426
0 43428 7 1 2 76187 82244
0 43429 7 1 2 77453 43428
0 43430 7 1 2 101828 43429
0 43431 5 1 1 43430
0 43432 7 1 2 43425 43431
0 43433 5 1 1 43432
0 43434 7 1 2 67892 43433
0 43435 5 1 1 43434
0 43436 7 1 2 79245 100905
0 43437 5 1 1 43436
0 43438 7 1 2 68709 89001
0 43439 7 1 2 79939 43438
0 43440 7 2 2 43437 43439
0 43441 7 1 2 79959 101695
0 43442 7 1 2 101830 43441
0 43443 5 1 1 43442
0 43444 7 1 2 43435 43443
0 43445 5 1 1 43444
0 43446 7 1 2 66278 43445
0 43447 5 1 1 43446
0 43448 7 1 2 79960 101672
0 43449 7 1 2 101831 43448
0 43450 5 1 1 43449
0 43451 7 1 2 43447 43450
0 43452 5 1 1 43451
0 43453 7 1 2 83146 43452
0 43454 5 1 1 43453
0 43455 7 6 2 82672 98089
0 43456 7 3 2 69831 75549
0 43457 7 1 2 81189 101838
0 43458 5 1 1 43457
0 43459 7 7 2 66033 72719
0 43460 7 1 2 71871 77092
0 43461 7 1 2 101841 43460
0 43462 5 2 1 43461
0 43463 7 1 2 43458 101848
0 43464 5 1 1 43463
0 43465 7 1 2 101832 43464
0 43466 5 1 1 43465
0 43467 7 1 2 9684 85936
0 43468 5 1 1 43467
0 43469 7 1 2 101842 43468
0 43470 5 1 1 43469
0 43471 7 1 2 70958 79781
0 43472 7 1 2 86119 43471
0 43473 5 1 1 43472
0 43474 7 1 2 43470 43473
0 43475 5 1 1 43474
0 43476 7 1 2 64974 43475
0 43477 5 1 1 43476
0 43478 7 1 2 71678 93334
0 43479 5 2 1 43478
0 43480 7 1 2 73164 75814
0 43481 5 1 1 43480
0 43482 7 1 2 101850 43481
0 43483 5 1 1 43482
0 43484 7 1 2 74824 71441
0 43485 7 1 2 43483 43484
0 43486 5 1 1 43485
0 43487 7 1 2 43477 43486
0 43488 5 1 1 43487
0 43489 7 1 2 68234 100620
0 43490 7 1 2 43488 43489
0 43491 5 1 1 43490
0 43492 7 1 2 43466 43491
0 43493 5 1 1 43492
0 43494 7 1 2 66546 43493
0 43495 5 1 1 43494
0 43496 7 1 2 74241 81190
0 43497 5 1 1 43496
0 43498 7 1 2 101849 43497
0 43499 5 2 1 43498
0 43500 7 1 2 90198 101852
0 43501 5 1 1 43500
0 43502 7 1 2 77579 77935
0 43503 7 1 2 76434 43502
0 43504 7 1 2 81427 43503
0 43505 5 1 1 43504
0 43506 7 1 2 43501 43505
0 43507 5 1 1 43506
0 43508 7 1 2 99023 43507
0 43509 5 1 1 43508
0 43510 7 1 2 43495 43509
0 43511 5 1 1 43510
0 43512 7 1 2 67893 43511
0 43513 5 1 1 43512
0 43514 7 1 2 91877 98389
0 43515 7 1 2 101853 43514
0 43516 5 1 1 43515
0 43517 7 1 2 43513 43516
0 43518 5 1 1 43517
0 43519 7 1 2 69039 43518
0 43520 5 1 1 43519
0 43521 7 4 2 66279 82673
0 43522 7 1 2 75422 101854
0 43523 5 1 1 43522
0 43524 7 1 2 81830 75815
0 43525 7 1 2 91813 43524
0 43526 5 1 1 43525
0 43527 7 1 2 43523 43526
0 43528 5 1 1 43527
0 43529 7 1 2 66547 43528
0 43530 5 1 1 43529
0 43531 7 1 2 91294 97574
0 43532 5 1 1 43531
0 43533 7 1 2 43530 43532
0 43534 5 1 1 43533
0 43535 7 1 2 67894 43534
0 43536 5 1 1 43535
0 43537 7 3 2 66280 76564
0 43538 7 1 2 89920 92557
0 43539 7 1 2 101858 43538
0 43540 5 1 1 43539
0 43541 7 1 2 43536 43540
0 43542 5 1 1 43541
0 43543 7 1 2 88931 43542
0 43544 5 1 1 43543
0 43545 7 1 2 85646 78717
0 43546 7 4 2 61395 61905
0 43547 5 1 1 101861
0 43548 7 1 2 93574 101862
0 43549 7 1 2 43545 43548
0 43550 5 1 1 43549
0 43551 7 1 2 43544 43550
0 43552 5 1 1 43551
0 43553 7 1 2 64178 43552
0 43554 5 1 1 43553
0 43555 7 1 2 82633 95851
0 43556 7 1 2 101441 43555
0 43557 5 1 1 43556
0 43558 7 1 2 43554 43557
0 43559 5 1 1 43558
0 43560 7 1 2 67515 43559
0 43561 5 1 1 43560
0 43562 7 2 2 81214 74249
0 43563 7 1 2 84191 101435
0 43564 7 1 2 101865 43563
0 43565 5 1 1 43564
0 43566 7 1 2 43561 43565
0 43567 5 1 1 43566
0 43568 7 1 2 74825 43567
0 43569 5 1 1 43568
0 43570 7 1 2 43520 43569
0 43571 5 1 1 43570
0 43572 7 1 2 64566 43571
0 43573 5 1 1 43572
0 43574 7 3 2 64975 98303
0 43575 7 1 2 94544 101867
0 43576 5 1 1 43575
0 43577 7 3 2 69832 82634
0 43578 5 1 1 101870
0 43579 7 1 2 72644 101871
0 43580 5 1 1 43579
0 43581 7 1 2 43576 43580
0 43582 5 1 1 43581
0 43583 7 1 2 62888 43582
0 43584 5 1 1 43583
0 43585 7 1 2 83491 101598
0 43586 5 1 1 43585
0 43587 7 1 2 43584 43586
0 43588 5 1 1 43587
0 43589 7 1 2 68469 43588
0 43590 5 1 1 43589
0 43591 7 1 2 75827 77485
0 43592 5 1 1 43591
0 43593 7 1 2 43590 43592
0 43594 5 1 1 43593
0 43595 7 1 2 68710 43594
0 43596 5 1 1 43595
0 43597 7 1 2 88414 89384
0 43598 7 1 2 101868 43597
0 43599 5 1 1 43598
0 43600 7 1 2 43596 43599
0 43601 5 1 1 43600
0 43602 7 4 2 91878 98476
0 43603 5 1 1 101873
0 43604 7 1 2 86873 101874
0 43605 7 1 2 43601 43604
0 43606 5 1 1 43605
0 43607 7 1 2 43573 43606
0 43608 5 1 1 43607
0 43609 7 1 2 65518 43608
0 43610 5 1 1 43609
0 43611 7 1 2 43454 43610
0 43612 5 1 1 43611
0 43613 7 1 2 69246 43612
0 43614 5 1 1 43613
0 43615 7 1 2 90925 101855
0 43616 5 1 1 43615
0 43617 7 1 2 82424 100621
0 43618 7 1 2 99139 43617
0 43619 5 1 1 43618
0 43620 7 1 2 43616 43619
0 43621 5 1 1 43620
0 43622 7 1 2 66548 43621
0 43623 5 1 1 43622
0 43624 7 1 2 90592 83784
0 43625 5 1 1 43624
0 43626 7 1 2 97851 43625
0 43627 5 1 1 43626
0 43628 7 1 2 99024 43627
0 43629 5 1 1 43628
0 43630 7 1 2 43623 43629
0 43631 5 1 1 43630
0 43632 7 1 2 67300 43631
0 43633 5 1 1 43632
0 43634 7 1 2 66281 71496
0 43635 7 1 2 76188 43634
0 43636 7 1 2 89693 43635
0 43637 5 1 1 43636
0 43638 7 1 2 43633 43637
0 43639 5 1 1 43638
0 43640 7 1 2 67895 43639
0 43641 5 1 1 43640
0 43642 7 1 2 93762 95524
0 43643 7 1 2 97849 43642
0 43644 5 1 1 43643
0 43645 7 1 2 43641 43644
0 43646 5 1 1 43645
0 43647 7 1 2 88381 93064
0 43648 7 1 2 43646 43647
0 43649 5 1 1 43648
0 43650 7 1 2 96021 98842
0 43651 7 3 2 69419 74629
0 43652 7 2 2 66282 98700
0 43653 7 1 2 101877 101880
0 43654 7 1 2 43650 43653
0 43655 5 1 1 43654
0 43656 7 1 2 43649 43655
0 43657 5 1 1 43656
0 43658 7 1 2 71102 43657
0 43659 5 1 1 43658
0 43660 7 2 2 64567 100133
0 43661 7 1 2 74375 101807
0 43662 5 1 1 43661
0 43663 7 1 2 84322 74406
0 43664 7 1 2 86898 43663
0 43665 5 1 1 43664
0 43666 7 1 2 43662 43665
0 43667 5 1 1 43666
0 43668 7 1 2 101882 43667
0 43669 5 1 1 43668
0 43670 7 2 2 74604 73655
0 43671 7 1 2 101684 101884
0 43672 5 1 1 43671
0 43673 7 1 2 43669 43672
0 43674 5 1 1 43673
0 43675 7 1 2 66283 43674
0 43676 5 1 1 43675
0 43677 7 3 2 93129 93751
0 43678 5 2 1 101886
0 43679 7 1 2 101885 101887
0 43680 5 1 1 43679
0 43681 7 1 2 43676 43680
0 43682 5 1 1 43681
0 43683 7 1 2 83694 43682
0 43684 5 1 1 43683
0 43685 7 1 2 81601 92973
0 43686 7 1 2 101135 43685
0 43687 7 1 2 79215 43686
0 43688 5 1 1 43687
0 43689 7 1 2 43684 43688
0 43690 5 1 1 43689
0 43691 7 1 2 69833 43690
0 43692 5 1 1 43691
0 43693 7 3 2 67731 94024
0 43694 7 1 2 92015 101891
0 43695 5 1 1 43694
0 43696 7 1 2 81100 101541
0 43697 5 1 1 43696
0 43698 7 1 2 43695 43697
0 43699 5 1 1 43698
0 43700 7 1 2 82747 43699
0 43701 5 1 1 43700
0 43702 7 1 2 79246 94420
0 43703 5 1 1 43702
0 43704 7 1 2 89005 43703
0 43705 5 1 1 43704
0 43706 7 1 2 43701 43705
0 43707 5 1 1 43706
0 43708 7 1 2 63630 43707
0 43709 5 1 1 43708
0 43710 7 2 2 64568 91308
0 43711 7 1 2 62195 94416
0 43712 7 1 2 101894 43711
0 43713 5 1 1 43712
0 43714 7 1 2 43709 43713
0 43715 5 1 1 43714
0 43716 7 1 2 67896 43715
0 43717 5 1 1 43716
0 43718 7 2 2 74376 72720
0 43719 5 1 1 101896
0 43720 7 1 2 72577 43719
0 43721 5 2 1 43720
0 43722 7 1 2 83373 93930
0 43723 7 2 2 101898 43722
0 43724 7 2 2 96439 101900
0 43725 7 1 2 101594 101902
0 43726 5 1 1 43725
0 43727 7 1 2 74442 101895
0 43728 5 1 1 43727
0 43729 7 1 2 73165 87346
0 43730 7 1 2 101239 43729
0 43731 5 1 1 43730
0 43732 7 1 2 43728 43731
0 43733 5 1 1 43732
0 43734 7 1 2 67897 43733
0 43735 5 1 1 43734
0 43736 7 1 2 82290 98701
0 43737 7 1 2 84287 43736
0 43738 5 1 1 43737
0 43739 7 1 2 43735 43738
0 43740 5 1 1 43739
0 43741 7 1 2 98304 43740
0 43742 5 1 1 43741
0 43743 7 1 2 43726 43742
0 43744 7 1 2 43717 43743
0 43745 5 1 1 43744
0 43746 7 1 2 66284 43745
0 43747 5 1 1 43746
0 43748 7 1 2 101586 101903
0 43749 5 1 1 43748
0 43750 7 1 2 64569 98488
0 43751 7 1 2 101592 43750
0 43752 5 1 1 43751
0 43753 7 1 2 43749 43752
0 43754 7 1 2 43747 43753
0 43755 5 1 1 43754
0 43756 7 1 2 70433 96453
0 43757 7 1 2 43755 43756
0 43758 5 1 1 43757
0 43759 7 1 2 43692 43758
0 43760 5 1 1 43759
0 43761 7 1 2 73033 43760
0 43762 5 1 1 43761
0 43763 7 1 2 43659 43762
0 43764 7 1 2 43614 43763
0 43765 5 1 1 43764
0 43766 7 1 2 70132 43765
0 43767 5 1 1 43766
0 43768 7 1 2 68470 74591
0 43769 5 2 1 43768
0 43770 7 1 2 74826 99871
0 43771 5 1 1 43770
0 43772 7 1 2 101904 43771
0 43773 5 3 1 43772
0 43774 7 1 2 101843 101906
0 43775 5 1 1 43774
0 43776 7 1 2 75816 74592
0 43777 5 1 1 43776
0 43778 7 1 2 86423 43777
0 43779 5 3 1 43778
0 43780 7 1 2 91108 101909
0 43781 5 1 1 43780
0 43782 7 1 2 43775 43781
0 43783 5 1 1 43782
0 43784 7 1 2 69040 43783
0 43785 5 1 1 43784
0 43786 7 1 2 101780 101910
0 43787 5 1 1 43786
0 43788 7 1 2 43785 43787
0 43789 5 1 1 43788
0 43790 7 4 2 64570 101442
0 43791 7 1 2 101622 101912
0 43792 5 1 1 43791
0 43793 7 2 2 76189 90672
0 43794 7 1 2 81701 82006
0 43795 7 1 2 101916 43794
0 43796 5 1 1 43795
0 43797 7 1 2 43792 43796
0 43798 5 1 1 43797
0 43799 7 1 2 43789 43798
0 43800 5 1 1 43799
0 43801 7 1 2 100409 101907
0 43802 5 1 1 43801
0 43803 7 1 2 79981 101911
0 43804 5 1 1 43803
0 43805 7 1 2 43802 43804
0 43806 5 1 1 43805
0 43807 7 1 2 67516 43806
0 43808 5 1 1 43807
0 43809 7 1 2 89031 78217
0 43810 5 1 1 43809
0 43811 7 1 2 63631 86797
0 43812 5 1 1 43811
0 43813 7 1 2 43810 43812
0 43814 5 1 1 43813
0 43815 7 1 2 67040 43814
0 43816 5 1 1 43815
0 43817 7 1 2 75116 86487
0 43818 5 1 1 43817
0 43819 7 1 2 67301 74665
0 43820 5 3 1 43819
0 43821 7 1 2 101918 98753
0 43822 5 2 1 43821
0 43823 7 1 2 101790 101921
0 43824 5 1 1 43823
0 43825 7 1 2 43818 43824
0 43826 7 1 2 43816 43825
0 43827 5 1 1 43826
0 43828 7 1 2 68711 43827
0 43829 5 1 1 43828
0 43830 7 2 2 75817 90342
0 43831 7 1 2 62630 85998
0 43832 7 1 2 101923 43831
0 43833 5 1 1 43832
0 43834 7 1 2 43829 43833
0 43835 7 1 2 43808 43834
0 43836 5 1 1 43835
0 43837 7 5 2 100001 100598
0 43838 7 1 2 101623 101925
0 43839 7 1 2 43836 43838
0 43840 5 1 1 43839
0 43841 7 1 2 43800 43840
0 43842 5 1 1 43841
0 43843 7 1 2 100637 43842
0 43844 5 1 1 43843
0 43845 7 1 2 43767 43844
0 43846 5 1 1 43845
0 43847 7 1 2 69622 43846
0 43848 5 1 1 43847
0 43849 7 1 2 80718 77675
0 43850 5 4 1 43849
0 43851 7 1 2 101635 101930
0 43852 5 1 1 43851
0 43853 7 1 2 78044 89197
0 43854 5 1 1 43853
0 43855 7 1 2 43852 43854
0 43856 5 1 1 43855
0 43857 7 1 2 69041 43856
0 43858 5 1 1 43857
0 43859 7 1 2 101639 101931
0 43860 5 1 1 43859
0 43861 7 1 2 43858 43860
0 43862 5 1 1 43861
0 43863 7 1 2 67302 43862
0 43864 5 1 1 43863
0 43865 7 1 2 68471 84703
0 43866 7 1 2 79623 43865
0 43867 5 1 1 43866
0 43868 7 1 2 43864 43867
0 43869 5 1 1 43868
0 43870 7 1 2 90075 43869
0 43871 5 1 1 43870
0 43872 7 1 2 77175 79266
0 43873 7 1 2 93466 43872
0 43874 5 1 1 43873
0 43875 7 1 2 43871 43874
0 43876 5 1 1 43875
0 43877 7 1 2 65519 43876
0 43878 5 1 1 43877
0 43879 7 3 2 78077 75256
0 43880 7 2 2 101797 101934
0 43881 7 1 2 87279 101937
0 43882 5 1 1 43881
0 43883 7 1 2 43878 43882
0 43884 5 1 1 43883
0 43885 7 1 2 69420 43884
0 43886 5 1 1 43885
0 43887 7 1 2 88407 89712
0 43888 7 1 2 101552 43887
0 43889 5 1 1 43888
0 43890 7 1 2 43886 43889
0 43891 5 1 1 43890
0 43892 7 1 2 68712 43891
0 43893 5 1 1 43892
0 43894 7 2 2 76579 79940
0 43895 7 1 2 101188 101939
0 43896 5 1 1 43895
0 43897 7 1 2 100323 98789
0 43898 5 1 1 43897
0 43899 7 1 2 43896 43898
0 43900 5 1 1 43899
0 43901 7 1 2 66549 43900
0 43902 5 1 1 43901
0 43903 7 1 2 76061 86657
0 43904 7 1 2 101940 43903
0 43905 5 1 1 43904
0 43906 7 1 2 43902 43905
0 43907 5 1 1 43906
0 43908 7 1 2 62889 43907
0 43909 5 1 1 43908
0 43910 7 1 2 70959 92318
0 43911 7 1 2 101935 43910
0 43912 5 1 1 43911
0 43913 7 1 2 43909 43912
0 43914 5 1 1 43913
0 43915 7 1 2 69421 43914
0 43916 5 1 1 43915
0 43917 7 2 2 83822 88591
0 43918 7 1 2 85766 90084
0 43919 7 1 2 101941 43918
0 43920 5 1 1 43919
0 43921 7 1 2 43916 43920
0 43922 5 1 1 43921
0 43923 7 1 2 64179 43922
0 43924 5 1 1 43923
0 43925 7 2 2 10137 101632
0 43926 5 1 1 101943
0 43927 7 1 2 82343 43926
0 43928 5 1 1 43927
0 43929 7 1 2 83835 73583
0 43930 7 1 2 88891 43929
0 43931 5 1 1 43930
0 43932 7 1 2 43928 43931
0 43933 5 1 1 43932
0 43934 7 1 2 69042 43933
0 43935 5 1 1 43934
0 43936 7 1 2 81101 84896
0 43937 5 1 1 43936
0 43938 7 1 2 43935 43937
0 43939 5 1 1 43938
0 43940 7 1 2 101936 43939
0 43941 5 1 1 43940
0 43942 7 1 2 43924 43941
0 43943 5 1 1 43942
0 43944 7 1 2 72944 43943
0 43945 5 1 1 43944
0 43946 7 1 2 43893 43945
0 43947 5 1 1 43946
0 43948 7 1 2 90673 43947
0 43949 5 1 1 43948
0 43950 7 1 2 75550 98748
0 43951 5 1 1 43950
0 43952 7 1 2 101851 43951
0 43953 5 1 1 43952
0 43954 7 1 2 99654 43953
0 43955 5 1 1 43954
0 43956 7 1 2 88736 98997
0 43957 5 1 1 43956
0 43958 7 1 2 43955 43957
0 43959 5 1 1 43958
0 43960 7 1 2 66285 43959
0 43961 5 1 1 43960
0 43962 7 1 2 93335 100553
0 43963 5 1 1 43962
0 43964 7 1 2 43961 43963
0 43965 5 1 1 43964
0 43966 7 1 2 64976 90540
0 43967 7 1 2 43965 43966
0 43968 5 1 1 43967
0 43969 7 1 2 89236 101926
0 43970 5 1 1 43969
0 43971 7 1 2 101844 101913
0 43972 5 1 1 43971
0 43973 7 1 2 43970 43972
0 43974 5 1 1 43973
0 43975 7 1 2 62196 81359
0 43976 7 1 2 43974 43975
0 43977 5 1 1 43976
0 43978 7 1 2 43968 43977
0 43979 5 1 1 43978
0 43980 7 1 2 69043 43979
0 43981 5 1 1 43980
0 43982 7 1 2 83214 75236
0 43983 7 1 2 81012 43982
0 43984 5 1 1 43983
0 43985 7 1 2 75818 88682
0 43986 7 1 2 90076 43985
0 43987 5 1 1 43986
0 43988 7 1 2 43984 43987
0 43989 5 1 1 43988
0 43990 7 1 2 86311 92974
0 43991 7 1 2 43989 43990
0 43992 5 1 1 43991
0 43993 7 1 2 43981 43992
0 43994 5 1 1 43993
0 43995 7 1 2 74593 43994
0 43996 5 1 1 43995
0 43997 7 1 2 77905 78045
0 43998 7 1 2 89598 79941
0 43999 7 1 2 43997 43998
0 44000 5 1 1 43999
0 44001 7 1 2 90085 92286
0 44002 7 1 2 101550 44001
0 44003 5 1 1 44002
0 44004 7 1 2 44000 44003
0 44005 5 1 1 44004
0 44006 7 1 2 66550 44005
0 44007 5 1 1 44006
0 44008 7 1 2 86584 91820
0 44009 7 1 2 98131 44008
0 44010 5 1 1 44009
0 44011 7 1 2 44007 44010
0 44012 5 1 1 44011
0 44013 7 8 2 64571 93809
0 44014 7 1 2 63632 101945
0 44015 7 1 2 44012 44014
0 44016 5 1 1 44015
0 44017 7 1 2 43996 44016
0 44018 7 1 2 43949 44017
0 44019 5 1 1 44018
0 44020 7 1 2 83147 44019
0 44021 5 1 1 44020
0 44022 7 2 2 72578 77768
0 44023 5 1 1 101953
0 44024 7 1 2 86079 44023
0 44025 5 1 1 44024
0 44026 7 1 2 62197 44025
0 44027 5 1 1 44026
0 44028 7 1 2 82199 74988
0 44029 5 1 1 44028
0 44030 7 1 2 44027 44029
0 44031 5 1 1 44030
0 44032 7 1 2 78555 44031
0 44033 5 1 1 44032
0 44034 7 1 2 94982 101954
0 44035 5 1 1 44034
0 44036 7 1 2 44033 44035
0 44037 5 1 1 44036
0 44038 7 1 2 62631 44037
0 44039 5 1 1 44038
0 44040 7 2 2 79982 94983
0 44041 5 1 1 101955
0 44042 7 1 2 76652 101956
0 44043 5 1 1 44042
0 44044 7 1 2 44039 44043
0 44045 5 2 1 44044
0 44046 7 1 2 99655 101957
0 44047 5 1 1 44046
0 44048 7 3 2 65205 82245
0 44049 7 1 2 68472 101542
0 44050 5 1 1 44049
0 44051 7 4 2 67041 72645
0 44052 5 1 1 101962
0 44053 7 1 2 67517 101963
0 44054 5 1 1 44053
0 44055 7 1 2 44050 44054
0 44056 5 1 1 44055
0 44057 7 2 2 101959 44056
0 44058 7 1 2 98761 101966
0 44059 5 1 1 44058
0 44060 7 1 2 44047 44059
0 44061 5 1 1 44060
0 44062 7 1 2 66286 44061
0 44063 5 1 1 44062
0 44064 7 2 2 62441 93752
0 44065 7 1 2 101967 101968
0 44066 5 1 1 44065
0 44067 7 1 2 44063 44066
0 44068 5 1 1 44067
0 44069 7 1 2 74551 44068
0 44070 5 1 1 44069
0 44071 7 1 2 85826 77563
0 44072 5 1 1 44071
0 44073 7 1 2 87609 44072
0 44074 5 1 1 44073
0 44075 7 1 2 62198 44074
0 44076 5 1 1 44075
0 44077 7 1 2 84704 78575
0 44078 5 2 1 44077
0 44079 7 1 2 77398 91701
0 44080 5 1 1 44079
0 44081 7 1 2 101970 44080
0 44082 7 1 2 44076 44081
0 44083 5 1 1 44082
0 44084 7 1 2 86798 44083
0 44085 5 1 1 44084
0 44086 7 2 2 78556 76598
0 44087 7 1 2 77801 74407
0 44088 7 1 2 101972 44087
0 44089 5 1 1 44088
0 44090 7 1 2 44085 44089
0 44091 5 1 1 44090
0 44092 7 1 2 99656 44091
0 44093 5 1 1 44092
0 44094 7 1 2 948 87188
0 44095 5 1 1 44094
0 44096 7 1 2 72579 44095
0 44097 5 1 1 44096
0 44098 7 1 2 491 44097
0 44099 5 2 1 44098
0 44100 7 2 2 90166 101974
0 44101 7 1 2 98762 101976
0 44102 5 1 1 44101
0 44103 7 1 2 44093 44102
0 44104 5 1 1 44103
0 44105 7 1 2 66287 44104
0 44106 5 1 1 44105
0 44107 7 1 2 101969 101977
0 44108 5 1 1 44107
0 44109 7 1 2 44106 44108
0 44110 5 1 1 44109
0 44111 7 1 2 68713 44110
0 44112 5 1 1 44111
0 44113 7 1 2 84965 44052
0 44114 5 1 1 44113
0 44115 7 1 2 67518 44114
0 44116 5 1 1 44115
0 44117 7 1 2 68473 94496
0 44118 5 1 1 44117
0 44119 7 1 2 44116 44118
0 44120 5 1 1 44119
0 44121 7 1 2 76966 44120
0 44122 5 1 1 44121
0 44123 7 1 2 79823 85054
0 44124 7 1 2 93966 44123
0 44125 5 1 1 44124
0 44126 7 1 2 44122 44125
0 44127 5 1 1 44126
0 44128 7 1 2 69834 44127
0 44129 5 1 1 44128
0 44130 7 1 2 101557 101975
0 44131 5 1 1 44130
0 44132 7 1 2 44129 44131
0 44133 5 1 1 44132
0 44134 7 1 2 101946 44133
0 44135 5 1 1 44134
0 44136 7 3 2 69835 94025
0 44137 7 1 2 67042 76977
0 44138 5 1 1 44137
0 44139 7 1 2 85684 95355
0 44140 5 1 1 44139
0 44141 7 1 2 44138 44140
0 44142 5 2 1 44141
0 44143 7 1 2 101978 101981
0 44144 5 1 1 44143
0 44145 7 1 2 74458 79493
0 44146 7 1 2 86905 44145
0 44147 5 1 1 44146
0 44148 7 1 2 44144 44147
0 44149 5 1 1 44148
0 44150 7 1 2 67732 44149
0 44151 5 1 1 44150
0 44152 7 1 2 95457 101973
0 44153 5 1 1 44152
0 44154 7 1 2 44151 44153
0 44155 5 1 1 44154
0 44156 7 1 2 100203 44155
0 44157 5 1 1 44156
0 44158 7 1 2 44135 44157
0 44159 5 1 1 44158
0 44160 7 1 2 67303 44159
0 44161 5 1 1 44160
0 44162 7 1 2 74827 101960
0 44163 7 1 2 99847 44162
0 44164 5 1 1 44163
0 44165 7 1 2 80300 93484
0 44166 7 1 2 101370 44165
0 44167 5 1 1 44166
0 44168 7 1 2 44164 44167
0 44169 5 1 1 44168
0 44170 7 1 2 63633 44169
0 44171 5 1 1 44170
0 44172 7 2 2 70434 93810
0 44173 7 1 2 67304 100070
0 44174 7 1 2 87598 44173
0 44175 7 1 2 101983 44174
0 44176 5 1 1 44175
0 44177 7 1 2 44171 44176
0 44178 5 1 1 44177
0 44179 7 1 2 101609 44178
0 44180 5 1 1 44179
0 44181 7 1 2 75819 100189
0 44182 5 1 1 44181
0 44183 7 3 2 66288 73166
0 44184 7 1 2 69422 93575
0 44185 7 1 2 101985 44184
0 44186 5 1 1 44185
0 44187 7 1 2 44182 44186
0 44188 5 1 1 44187
0 44189 7 1 2 78608 44188
0 44190 5 1 1 44189
0 44191 7 1 2 78557 83396
0 44192 7 1 2 92975 44191
0 44193 5 1 1 44192
0 44194 7 1 2 44190 44193
0 44195 5 1 1 44194
0 44196 7 1 2 74419 44195
0 44197 5 1 1 44196
0 44198 7 1 2 67043 79031
0 44199 5 1 1 44198
0 44200 7 1 2 86816 74870
0 44201 5 1 1 44200
0 44202 7 1 2 44199 44201
0 44203 5 2 1 44202
0 44204 7 1 2 100190 101988
0 44205 5 1 1 44204
0 44206 7 1 2 74377 74828
0 44207 5 1 1 44206
0 44208 7 1 2 74057 44207
0 44209 5 1 1 44208
0 44210 7 1 2 76868 99657
0 44211 7 1 2 100793 44210
0 44212 7 1 2 44209 44211
0 44213 5 1 1 44212
0 44214 7 1 2 44205 44213
0 44215 5 1 1 44214
0 44216 7 1 2 76781 44215
0 44217 5 1 1 44216
0 44218 7 1 2 44197 44217
0 44219 5 1 1 44218
0 44220 7 1 2 98305 44219
0 44221 5 1 1 44220
0 44222 7 1 2 86312 90674
0 44223 7 1 2 88710 44222
0 44224 7 1 2 92349 98282
0 44225 7 1 2 44223 44224
0 44226 5 1 1 44225
0 44227 7 1 2 44221 44226
0 44228 7 1 2 44180 44227
0 44229 7 1 2 44161 44228
0 44230 7 1 2 44112 44229
0 44231 7 1 2 44070 44230
0 44232 5 1 1 44231
0 44233 7 1 2 92911 44232
0 44234 5 1 1 44233
0 44235 7 1 2 101833 101982
0 44236 5 1 1 44235
0 44237 7 2 2 76899 91814
0 44238 7 1 2 81831 73923
0 44239 7 2 2 101990 44238
0 44240 5 1 1 101992
0 44241 7 1 2 44236 44240
0 44242 5 1 1 44241
0 44243 7 1 2 67305 44242
0 44244 5 1 1 44243
0 44245 7 1 2 94978 101834
0 44246 7 1 2 74557 44245
0 44247 5 1 1 44246
0 44248 7 1 2 44244 44247
0 44249 5 1 1 44248
0 44250 7 1 2 100897 44249
0 44251 5 1 1 44250
0 44252 7 1 2 87545 101991
0 44253 5 1 1 44252
0 44254 7 1 2 65206 101835
0 44255 7 1 2 101908 44254
0 44256 5 1 1 44255
0 44257 7 1 2 44253 44256
0 44258 5 1 1 44257
0 44259 7 1 2 94417 44258
0 44260 5 1 1 44259
0 44261 7 1 2 44251 44260
0 44262 5 1 1 44261
0 44263 7 1 2 69836 44262
0 44264 5 1 1 44263
0 44265 7 1 2 74420 94987
0 44266 5 1 1 44265
0 44267 7 1 2 76782 101989
0 44268 5 1 1 44267
0 44269 7 1 2 44266 44268
0 44270 5 1 1 44269
0 44271 7 1 2 101836 44270
0 44272 5 1 1 44271
0 44273 7 1 2 79880 101993
0 44274 5 1 1 44273
0 44275 7 1 2 44272 44274
0 44276 5 1 1 44275
0 44277 7 1 2 95870 44276
0 44278 5 1 1 44277
0 44279 7 2 2 61396 81560
0 44280 7 1 2 75967 80093
0 44281 7 1 2 101994 44280
0 44282 5 1 1 44281
0 44283 7 1 2 70435 72721
0 44284 7 1 2 101856 44283
0 44285 7 1 2 75390 44284
0 44286 5 1 1 44285
0 44287 7 1 2 44282 44286
0 44288 5 1 1 44287
0 44289 7 1 2 83273 44288
0 44290 5 1 1 44289
0 44291 7 1 2 44278 44290
0 44292 7 1 2 44264 44291
0 44293 5 1 1 44292
0 44294 7 1 2 64572 44293
0 44295 5 1 1 44294
0 44296 7 1 2 71065 101519
0 44297 5 1 1 44296
0 44298 7 1 2 76900 71442
0 44299 7 1 2 101798 44298
0 44300 5 1 1 44299
0 44301 7 1 2 44297 44300
0 44302 5 1 1 44301
0 44303 7 1 2 81832 98603
0 44304 7 1 2 88693 44303
0 44305 7 1 2 44302 44304
0 44306 5 1 1 44305
0 44307 7 1 2 44295 44306
0 44308 5 1 1 44307
0 44309 7 1 2 99108 44308
0 44310 5 1 1 44309
0 44311 7 1 2 44234 44310
0 44312 7 1 2 44021 44311
0 44313 5 1 1 44312
0 44314 7 1 2 92118 44313
0 44315 5 1 1 44314
0 44316 7 1 2 43848 44315
0 44317 5 1 1 44316
0 44318 7 1 2 96968 44317
0 44319 5 1 1 44318
0 44320 7 1 2 87408 92045
0 44321 5 1 1 44320
0 44322 7 1 2 32742 44321
0 44323 5 1 1 44322
0 44324 7 1 2 78078 86392
0 44325 7 2 2 101857 44324
0 44326 5 1 1 101996
0 44327 7 1 2 90343 99526
0 44328 7 1 2 91830 44327
0 44329 5 1 1 44328
0 44330 7 1 2 44326 44329
0 44331 5 1 1 44330
0 44332 7 1 2 44323 44331
0 44333 5 1 1 44332
0 44334 7 1 2 78680 90244
0 44335 5 1 1 44334
0 44336 7 1 2 69837 85827
0 44337 7 1 2 79267 44336
0 44338 5 1 1 44337
0 44339 7 1 2 44335 44338
0 44340 5 1 1 44339
0 44341 7 1 2 83148 44340
0 44342 5 1 1 44341
0 44343 7 1 2 83316 89210
0 44344 5 1 1 44343
0 44345 7 1 2 44342 44344
0 44346 5 1 1 44345
0 44347 7 1 2 64789 44346
0 44348 5 1 1 44347
0 44349 7 1 2 87610 86328
0 44350 5 3 1 44349
0 44351 7 1 2 68235 101998
0 44352 5 1 1 44351
0 44353 7 1 2 7802 44352
0 44354 5 1 1 44353
0 44355 7 1 2 62890 87076
0 44356 7 1 2 44354 44355
0 44357 5 1 1 44356
0 44358 7 1 2 44348 44357
0 44359 5 1 1 44358
0 44360 7 1 2 90344 44359
0 44361 5 1 1 44360
0 44362 7 2 2 78079 89983
0 44363 7 1 2 87409 81388
0 44364 5 1 1 44363
0 44365 7 2 2 68236 78480
0 44366 7 1 2 61653 102003
0 44367 5 1 1 44366
0 44368 7 1 2 44364 44367
0 44369 5 1 1 44368
0 44370 7 1 2 66773 44369
0 44371 5 1 1 44370
0 44372 7 2 2 83342 74242
0 44373 5 1 1 102005
0 44374 7 1 2 85647 102006
0 44375 5 1 1 44374
0 44376 7 1 2 44371 44375
0 44377 5 1 1 44376
0 44378 7 1 2 102001 44377
0 44379 5 1 1 44378
0 44380 7 1 2 44361 44379
0 44381 5 1 1 44380
0 44382 7 1 2 68040 44381
0 44383 5 1 1 44382
0 44384 7 3 2 75820 95463
0 44385 5 1 1 102007
0 44386 7 2 2 90345 102008
0 44387 7 1 2 102010 98032
0 44388 5 1 1 44387
0 44389 7 1 2 44383 44388
0 44390 5 1 1 44389
0 44391 7 1 2 61397 44390
0 44392 5 1 1 44391
0 44393 7 1 2 44333 44392
0 44394 5 1 1 44393
0 44395 7 1 2 69423 44394
0 44396 5 1 1 44395
0 44397 7 2 2 65520 71784
0 44398 7 1 2 91764 102012
0 44399 5 1 1 44398
0 44400 7 1 2 67306 83696
0 44401 5 1 1 44400
0 44402 7 1 2 44399 44401
0 44403 5 1 1 44402
0 44404 7 1 2 78080 82787
0 44405 7 1 2 99486 44404
0 44406 7 1 2 44403 44405
0 44407 5 1 1 44406
0 44408 7 1 2 44396 44407
0 44409 5 1 1 44408
0 44410 7 1 2 67519 44409
0 44411 5 1 1 44410
0 44412 7 2 2 61654 89454
0 44413 5 1 1 102014
0 44414 7 2 2 69838 84127
0 44415 7 1 2 77207 102016
0 44416 5 1 1 44415
0 44417 7 1 2 44413 44416
0 44418 5 5 1 44417
0 44419 7 1 2 94979 102018
0 44420 5 2 1 44419
0 44421 7 1 2 91984 92050
0 44422 5 1 1 44421
0 44423 7 1 2 102023 44422
0 44424 5 1 1 44423
0 44425 7 1 2 90346 44424
0 44426 5 2 1 44425
0 44427 7 4 2 75257 83595
0 44428 7 1 2 83294 93256
0 44429 7 1 2 102027 44428
0 44430 5 1 1 44429
0 44431 7 1 2 102025 44430
0 44432 5 1 1 44431
0 44433 7 1 2 80144 99487
0 44434 7 1 2 44432 44433
0 44435 5 1 1 44434
0 44436 7 1 2 44411 44435
0 44437 5 1 1 44436
0 44438 7 1 2 98306 44437
0 44439 5 1 1 44438
0 44440 7 1 2 62442 101829
0 44441 5 1 1 44440
0 44442 7 1 2 74378 90383
0 44443 5 1 1 44442
0 44444 7 1 2 44441 44443
0 44445 5 1 1 44444
0 44446 7 1 2 62632 44445
0 44447 5 1 1 44446
0 44448 7 3 2 67520 71171
0 44449 7 2 2 82200 102031
0 44450 5 1 1 102034
0 44451 7 1 2 70436 102035
0 44452 5 1 1 44451
0 44453 7 1 2 44447 44452
0 44454 5 1 1 44453
0 44455 7 1 2 88196 44454
0 44456 5 1 1 44455
0 44457 7 1 2 90347 93270
0 44458 7 1 2 67044 74715
0 44459 5 1 1 44458
0 44460 7 1 2 101845 44459
0 44461 7 1 2 44457 44460
0 44462 5 1 1 44461
0 44463 7 1 2 44456 44462
0 44464 5 1 1 44463
0 44465 7 1 2 83149 44464
0 44466 5 1 1 44465
0 44467 7 1 2 86979 72722
0 44468 5 1 1 44467
0 44469 7 1 2 69623 90082
0 44470 5 1 1 44469
0 44471 7 1 2 44468 44470
0 44472 5 1 1 44471
0 44473 7 1 2 66034 44472
0 44474 5 1 1 44473
0 44475 7 1 2 67521 95599
0 44476 5 1 1 44475
0 44477 7 1 2 44474 44476
0 44478 5 1 1 44477
0 44479 7 1 2 69044 44478
0 44480 5 1 1 44479
0 44481 7 1 2 28995 44480
0 44482 5 1 1 44481
0 44483 7 1 2 83569 102013
0 44484 7 1 2 44482 44483
0 44485 5 1 1 44484
0 44486 7 1 2 44466 44485
0 44487 5 1 1 44486
0 44488 7 1 2 69839 44487
0 44489 5 1 1 44488
0 44490 7 1 2 81940 90348
0 44491 5 1 1 44490
0 44492 7 1 2 44491 41451
0 44493 5 1 1 44492
0 44494 7 1 2 101897 44493
0 44495 5 1 1 44494
0 44496 7 1 2 61655 76824
0 44497 7 1 2 88129 44496
0 44498 5 1 1 44497
0 44499 7 1 2 44495 44498
0 44500 5 1 1 44499
0 44501 7 1 2 81215 101536
0 44502 7 1 2 44500 44501
0 44503 5 1 1 44502
0 44504 7 1 2 44489 44503
0 44505 5 1 1 44504
0 44506 7 1 2 70133 44505
0 44507 5 1 1 44506
0 44508 7 1 2 80863 80748
0 44509 7 1 2 90349 44508
0 44510 7 1 2 101846 44509
0 44511 7 1 2 102019 44510
0 44512 5 1 1 44511
0 44513 7 1 2 44507 44512
0 44514 5 1 1 44513
0 44515 7 1 2 99488 44514
0 44516 5 1 1 44515
0 44517 7 1 2 96055 101808
0 44518 5 1 1 44517
0 44519 7 1 2 7192 44385
0 44520 5 1 1 44519
0 44521 7 2 2 71172 86381
0 44522 7 1 2 44520 102036
0 44523 5 1 1 44522
0 44524 7 1 2 44518 44523
0 44525 5 1 1 44524
0 44526 7 1 2 67307 44525
0 44527 5 1 1 44526
0 44528 7 2 2 65207 74630
0 44529 7 1 2 87172 102038
0 44530 5 1 1 44529
0 44531 7 1 2 85192 93239
0 44532 5 1 1 44531
0 44533 7 1 2 44530 44532
0 44534 5 1 1 44533
0 44535 7 1 2 66774 44534
0 44536 5 1 1 44535
0 44537 7 1 2 68237 85880
0 44538 7 1 2 97898 44537
0 44539 5 1 1 44538
0 44540 7 1 2 44536 44539
0 44541 5 1 1 44540
0 44542 7 1 2 101284 44541
0 44543 5 1 1 44542
0 44544 7 1 2 44527 44543
0 44545 5 1 1 44544
0 44546 7 1 2 100622 44545
0 44547 5 1 1 44546
0 44548 7 1 2 85144 100623
0 44549 5 1 1 44548
0 44550 7 1 2 93082 98090
0 44551 5 1 1 44550
0 44552 7 1 2 44549 44551
0 44553 5 1 1 44552
0 44554 7 1 2 101517 44553
0 44555 5 1 1 44554
0 44556 7 1 2 100624 102009
0 44557 5 1 1 44556
0 44558 7 1 2 66289 88773
0 44559 7 1 2 91985 44558
0 44560 5 1 1 44559
0 44561 7 1 2 44557 44560
0 44562 5 1 1 44561
0 44563 7 1 2 65521 102032
0 44564 7 1 2 44562 44563
0 44565 5 1 1 44564
0 44566 7 1 2 44555 44565
0 44567 5 1 1 44566
0 44568 7 1 2 62443 44567
0 44569 5 1 1 44568
0 44570 7 1 2 44547 44569
0 44571 5 1 1 44570
0 44572 7 1 2 61656 44571
0 44573 5 1 1 44572
0 44574 7 1 2 73731 101630
0 44575 5 1 1 44574
0 44576 7 1 2 71173 98749
0 44577 5 1 1 44576
0 44578 7 1 2 44575 44577
0 44579 5 1 1 44578
0 44580 7 1 2 90350 44579
0 44581 5 1 1 44580
0 44582 7 1 2 84019 79831
0 44583 7 1 2 88617 44582
0 44584 5 1 1 44583
0 44585 7 1 2 44581 44584
0 44586 5 1 1 44585
0 44587 7 1 2 90048 99527
0 44588 7 1 2 44586 44587
0 44589 5 1 1 44588
0 44590 7 1 2 44573 44589
0 44591 5 1 1 44590
0 44592 7 1 2 64790 44591
0 44593 5 1 1 44592
0 44594 7 1 2 86393 101837
0 44595 5 1 1 44594
0 44596 7 1 2 61398 97818
0 44597 7 1 2 95613 44596
0 44598 5 1 1 44597
0 44599 7 1 2 44595 44598
0 44600 5 1 1 44599
0 44601 7 1 2 78081 44600
0 44602 5 1 1 44601
0 44603 7 1 2 100625 102011
0 44604 5 1 1 44603
0 44605 7 1 2 44602 44604
0 44606 5 1 1 44605
0 44607 7 1 2 91530 94026
0 44608 7 1 2 44606 44607
0 44609 5 1 1 44608
0 44610 7 1 2 44593 44609
0 44611 5 1 1 44610
0 44612 7 1 2 64977 44611
0 44613 5 1 1 44612
0 44614 7 2 2 65208 101924
0 44615 7 1 2 81848 102040
0 44616 5 1 1 44615
0 44617 7 1 2 88446 89171
0 44618 5 1 1 44617
0 44619 7 1 2 44616 44618
0 44620 5 1 1 44619
0 44621 7 1 2 100626 44620
0 44622 5 1 1 44621
0 44623 7 1 2 61657 101997
0 44624 5 1 1 44623
0 44625 7 1 2 44622 44624
0 44626 5 1 1 44625
0 44627 7 1 2 64791 44626
0 44628 5 1 1 44627
0 44629 7 1 2 88333 92199
0 44630 7 1 2 102041 44629
0 44631 5 1 1 44630
0 44632 7 1 2 44628 44631
0 44633 5 1 1 44632
0 44634 7 1 2 66775 44633
0 44635 5 1 1 44634
0 44636 7 2 2 61399 80994
0 44637 5 1 1 102042
0 44638 7 1 2 83596 85104
0 44639 7 1 2 93257 44638
0 44640 7 1 2 102043 44639
0 44641 5 1 1 44640
0 44642 7 1 2 44635 44641
0 44643 5 1 1 44642
0 44644 7 1 2 67733 101979
0 44645 7 1 2 44643 44644
0 44646 5 1 1 44645
0 44647 7 1 2 44613 44646
0 44648 5 1 1 44647
0 44649 7 1 2 69424 44648
0 44650 5 1 1 44649
0 44651 7 1 2 44516 44650
0 44652 7 1 2 44439 44651
0 44653 5 1 1 44652
0 44654 7 1 2 94786 99220
0 44655 7 1 2 44653 44654
0 44656 5 1 1 44655
0 44657 7 1 2 72074 95346
0 44658 5 1 1 44657
0 44659 7 3 2 74955 94027
0 44660 5 2 1 102044
0 44661 7 1 2 102045 101932
0 44662 5 1 1 44661
0 44663 7 1 2 44658 44662
0 44664 5 1 1 44663
0 44665 7 1 2 96879 44664
0 44666 5 1 1 44665
0 44667 7 1 2 89177 87696
0 44668 5 1 1 44667
0 44669 7 1 2 44666 44668
0 44670 5 1 1 44669
0 44671 7 1 2 64978 44670
0 44672 5 1 1 44671
0 44673 7 1 2 62199 88081
0 44674 5 1 1 44673
0 44675 7 1 2 83433 44674
0 44676 5 1 1 44675
0 44677 7 1 2 94883 44676
0 44678 5 1 1 44677
0 44679 7 1 2 72075 44678
0 44680 5 1 1 44679
0 44681 7 2 2 74010 87212
0 44682 7 1 2 74605 78046
0 44683 7 1 2 102049 44682
0 44684 5 1 1 44683
0 44685 7 1 2 44680 44684
0 44686 5 1 1 44685
0 44687 7 1 2 61906 44686
0 44688 5 1 1 44687
0 44689 7 1 2 81460 89178
0 44690 5 1 1 44689
0 44691 7 1 2 44688 44690
0 44692 5 1 1 44691
0 44693 7 1 2 92025 44692
0 44694 5 1 1 44693
0 44695 7 1 2 44672 44694
0 44696 5 1 1 44695
0 44697 7 1 2 69624 44696
0 44698 5 1 1 44697
0 44699 7 2 2 83295 79136
0 44700 7 2 2 65209 77580
0 44701 7 1 2 74443 102053
0 44702 5 2 1 44701
0 44703 7 1 2 70134 88082
0 44704 5 1 1 44703
0 44705 7 1 2 67045 81062
0 44706 7 1 2 44704 44705
0 44707 5 1 1 44706
0 44708 7 1 2 102055 44707
0 44709 5 1 1 44708
0 44710 7 1 2 63396 44709
0 44711 5 1 1 44710
0 44712 7 1 2 94884 44711
0 44713 5 1 1 44712
0 44714 7 1 2 72076 44713
0 44715 5 1 1 44714
0 44716 7 1 2 72580 102050
0 44717 7 1 2 101933 44716
0 44718 5 1 1 44717
0 44719 7 1 2 44715 44718
0 44720 5 1 1 44719
0 44721 7 1 2 102051 44720
0 44722 5 1 1 44721
0 44723 7 1 2 98307 102054
0 44724 7 1 2 102020 44723
0 44725 5 1 1 44724
0 44726 7 1 2 88352 83343
0 44727 7 1 2 89214 44726
0 44728 7 1 2 98976 44727
0 44729 5 1 1 44728
0 44730 7 1 2 44725 44729
0 44731 5 1 1 44730
0 44732 7 1 2 74379 44731
0 44733 5 1 1 44732
0 44734 7 1 2 83068 81941
0 44735 7 1 2 88829 44734
0 44736 7 1 2 96156 44735
0 44737 5 1 1 44736
0 44738 7 1 2 44733 44737
0 44739 5 1 1 44738
0 44740 7 1 2 62891 44739
0 44741 5 1 1 44740
0 44742 7 1 2 44722 44741
0 44743 7 1 2 44698 44742
0 44744 5 1 1 44743
0 44745 7 1 2 94615 44744
0 44746 5 1 1 44745
0 44747 7 1 2 94130 94726
0 44748 7 1 2 95894 44747
0 44749 7 1 2 95347 44748
0 44750 5 1 1 44749
0 44751 7 1 2 44746 44750
0 44752 5 1 1 44751
0 44753 7 1 2 63200 44752
0 44754 5 1 1 44753
0 44755 7 1 2 82084 99301
0 44756 5 1 1 44755
0 44757 7 2 2 83397 86096
0 44758 7 1 2 93915 102057
0 44759 5 1 1 44758
0 44760 7 1 2 44756 44759
0 44761 5 1 1 44760
0 44762 7 1 2 62200 44761
0 44763 5 1 1 44762
0 44764 7 1 2 75098 94376
0 44765 7 1 2 82085 44764
0 44766 5 1 1 44765
0 44767 7 1 2 44763 44766
0 44768 5 1 1 44767
0 44769 7 1 2 83150 44768
0 44770 5 1 1 44769
0 44771 7 1 2 81687 94406
0 44772 7 1 2 99241 44771
0 44773 5 1 1 44772
0 44774 7 1 2 44770 44773
0 44775 5 1 1 44774
0 44776 7 1 2 76062 94131
0 44777 7 1 2 44775 44776
0 44778 5 1 1 44777
0 44779 7 1 2 44754 44778
0 44780 5 1 1 44779
0 44781 7 1 2 65522 44780
0 44782 5 1 1 44781
0 44783 7 1 2 86980 87310
0 44784 5 1 1 44783
0 44785 7 1 2 61907 89254
0 44786 5 1 1 44785
0 44787 7 1 2 44784 44786
0 44788 5 2 1 44787
0 44789 7 1 2 94028 102059
0 44790 5 1 1 44789
0 44791 7 1 2 83344 79242
0 44792 7 1 2 97296 44791
0 44793 5 1 1 44792
0 44794 7 1 2 44790 44793
0 44795 5 1 1 44794
0 44796 7 1 2 67734 44795
0 44797 5 1 1 44796
0 44798 7 1 2 82585 92728
0 44799 7 1 2 100360 44798
0 44800 5 1 1 44799
0 44801 7 1 2 44797 44800
0 44802 5 1 1 44801
0 44803 7 1 2 63634 44802
0 44804 5 1 1 44803
0 44805 7 1 2 87173 94794
0 44806 7 1 2 97484 44805
0 44807 5 1 1 44806
0 44808 7 1 2 73167 98308
0 44809 7 1 2 102060 44808
0 44810 5 1 1 44809
0 44811 7 1 2 44807 44810
0 44812 7 1 2 44804 44811
0 44813 5 1 1 44812
0 44814 7 1 2 62444 44813
0 44815 5 1 1 44814
0 44816 7 1 2 64792 76851
0 44817 7 1 2 82251 74250
0 44818 7 1 2 44816 44817
0 44819 7 1 2 88618 44818
0 44820 5 1 1 44819
0 44821 7 1 2 44815 44820
0 44822 5 1 1 44821
0 44823 7 1 2 78733 44822
0 44824 5 1 1 44823
0 44825 7 1 2 75821 101892
0 44826 5 1 1 44825
0 44827 7 1 2 77478 100410
0 44828 5 1 1 44827
0 44829 7 1 2 44826 44828
0 44830 5 1 1 44829
0 44831 7 1 2 79592 44830
0 44832 7 1 2 102021 44831
0 44833 5 1 1 44832
0 44834 7 1 2 44824 44833
0 44835 5 1 1 44834
0 44836 7 1 2 95156 97435
0 44837 7 1 2 44835 44836
0 44838 5 1 1 44837
0 44839 7 1 2 68714 44838
0 44840 7 1 2 44782 44839
0 44841 5 1 1 44840
0 44842 7 2 2 83151 98309
0 44843 7 1 2 85828 81148
0 44844 7 1 2 102061 44843
0 44845 5 1 1 44844
0 44846 7 1 2 89455 94980
0 44847 7 1 2 100424 44846
0 44848 5 1 1 44847
0 44849 7 1 2 44845 44848
0 44850 5 1 1 44849
0 44851 7 1 2 61658 44850
0 44852 5 1 1 44851
0 44853 7 1 2 100411 101999
0 44854 5 1 1 44853
0 44855 7 1 2 44041 44854
0 44856 5 2 1 44855
0 44857 7 1 2 85426 83533
0 44858 7 1 2 102063 44857
0 44859 5 1 1 44858
0 44860 7 1 2 44852 44859
0 44861 5 1 1 44860
0 44862 7 1 2 67522 44861
0 44863 5 1 1 44862
0 44864 7 1 2 83597 88977
0 44865 7 1 2 82915 44864
0 44866 5 1 1 44865
0 44867 7 1 2 102024 44866
0 44868 5 1 1 44867
0 44869 7 1 2 101791 44868
0 44870 5 1 1 44869
0 44871 7 1 2 44863 44870
0 44872 5 1 1 44871
0 44873 7 1 2 90351 44872
0 44874 5 1 1 44873
0 44875 7 1 2 101643 102002
0 44876 5 1 1 44875
0 44877 7 1 2 70135 101922
0 44878 5 1 1 44877
0 44879 7 1 2 1273 2298
0 44880 5 1 1 44879
0 44881 7 1 2 62201 86397
0 44882 7 1 2 44880 44881
0 44883 5 1 1 44882
0 44884 7 1 2 44878 44883
0 44885 5 1 1 44884
0 44886 7 1 2 92604 44885
0 44887 5 1 1 44886
0 44888 7 1 2 44876 44887
0 44889 5 1 1 44888
0 44890 7 1 2 88986 44889
0 44891 5 1 1 44890
0 44892 7 1 2 85039 101938
0 44893 5 1 1 44892
0 44894 7 1 2 44891 44893
0 44895 5 1 1 44894
0 44896 7 1 2 86981 44895
0 44897 5 1 1 44896
0 44898 7 1 2 82058 80492
0 44899 7 1 2 90155 44898
0 44900 7 1 2 101799 44899
0 44901 5 1 1 44900
0 44902 7 1 2 44897 44901
0 44903 7 1 2 44874 44902
0 44904 5 1 1 44903
0 44905 7 1 2 95105 44904
0 44906 5 1 1 44905
0 44907 7 1 2 88288 88523
0 44908 7 2 2 79137 91283
0 44909 7 1 2 95377 96162
0 44910 7 1 2 102065 44909
0 44911 7 1 2 44907 44910
0 44912 5 1 1 44911
0 44913 7 1 2 63848 44912
0 44914 7 1 2 44906 44913
0 44915 5 1 1 44914
0 44916 7 1 2 93811 44915
0 44917 7 1 2 44841 44916
0 44918 5 1 1 44917
0 44919 7 1 2 84305 76404
0 44920 5 1 1 44919
0 44921 7 1 2 82201 84662
0 44922 5 1 1 44921
0 44923 7 1 2 44920 44922
0 44924 5 1 1 44923
0 44925 7 1 2 62633 44924
0 44926 5 1 1 44925
0 44927 7 1 2 44926 44450
0 44928 5 2 1 44927
0 44929 7 1 2 78893 102067
0 44930 5 1 1 44929
0 44931 7 3 2 67308 71679
0 44932 7 1 2 93730 102069
0 44933 5 1 1 44932
0 44934 7 1 2 91165 79832
0 44935 5 1 1 44934
0 44936 7 1 2 44933 44935
0 44937 5 1 1 44936
0 44938 7 1 2 62202 44937
0 44939 5 1 1 44938
0 44940 7 1 2 10596 102047
0 44941 5 1 1 44940
0 44942 7 1 2 88869 44941
0 44943 5 1 1 44942
0 44944 7 1 2 44939 44943
0 44945 7 1 2 44930 44944
0 44946 5 1 1 44945
0 44947 7 1 2 65523 44946
0 44948 5 1 1 44947
0 44949 7 1 2 93337 97071
0 44950 5 1 1 44949
0 44951 7 1 2 71116 101785
0 44952 5 1 1 44951
0 44953 7 1 2 69045 89059
0 44954 5 1 1 44953
0 44955 7 1 2 44952 44954
0 44956 5 1 1 44955
0 44957 7 1 2 67523 44956
0 44958 5 1 1 44957
0 44959 7 1 2 89065 85843
0 44960 5 1 1 44959
0 44961 7 1 2 44958 44960
0 44962 5 1 1 44961
0 44963 7 1 2 75822 44962
0 44964 5 1 1 44963
0 44965 7 1 2 44950 44964
0 44966 5 1 1 44965
0 44967 7 1 2 77549 44966
0 44968 5 1 1 44967
0 44969 7 1 2 44948 44968
0 44970 5 1 1 44969
0 44971 7 1 2 66551 44970
0 44972 5 1 1 44971
0 44973 7 1 2 62445 98541
0 44974 5 1 1 44973
0 44975 7 1 2 101919 44974
0 44976 5 4 1 44975
0 44977 7 1 2 102072 102033
0 44978 5 1 1 44977
0 44979 7 2 2 74380 85034
0 44980 5 1 1 102076
0 44981 7 1 2 84663 102077
0 44982 5 1 1 44981
0 44983 7 2 2 62446 74754
0 44984 5 1 1 102078
0 44985 7 1 2 68474 102079
0 44986 5 1 1 44985
0 44987 7 1 2 44982 44986
0 44988 5 1 1 44987
0 44989 7 1 2 62634 44988
0 44990 5 1 1 44989
0 44991 7 1 2 44978 44990
0 44992 5 1 1 44991
0 44993 7 1 2 89088 44992
0 44994 5 1 1 44993
0 44995 7 1 2 44972 44994
0 44996 5 1 1 44995
0 44997 7 1 2 69425 44996
0 44998 5 1 1 44997
0 44999 7 1 2 81880 95780
0 45000 5 1 1 44999
0 45001 7 1 2 101173 45000
0 45002 5 1 1 45001
0 45003 7 1 2 102073 45002
0 45004 5 1 1 45003
0 45005 7 1 2 98754 44980
0 45006 5 4 1 45005
0 45007 7 1 2 73168 98261
0 45008 7 1 2 102080 45007
0 45009 5 1 1 45008
0 45010 7 1 2 45004 45009
0 45011 5 1 1 45010
0 45012 7 1 2 98310 45011
0 45013 5 1 1 45012
0 45014 7 1 2 72723 102081
0 45015 7 1 2 98250 45014
0 45016 5 1 1 45015
0 45017 7 1 2 45013 45016
0 45018 7 1 2 44998 45017
0 45019 5 1 1 45018
0 45020 7 1 2 84487 45019
0 45021 5 1 1 45020
0 45022 7 1 2 90079 101560
0 45023 5 1 1 45022
0 45024 7 1 2 88719 101847
0 45025 5 1 1 45024
0 45026 7 1 2 45023 45025
0 45027 5 1 1 45026
0 45028 7 1 2 69046 45027
0 45029 5 1 1 45028
0 45030 7 1 2 80213 75598
0 45031 7 1 2 89863 45030
0 45032 5 1 1 45031
0 45033 7 1 2 45029 45032
0 45034 5 1 1 45033
0 45035 7 1 2 102082 45034
0 45036 5 1 1 45035
0 45037 7 4 2 82748 84082
0 45038 7 1 2 72077 102084
0 45039 7 1 2 76390 45038
0 45040 5 1 1 45039
0 45041 7 1 2 88720 98311
0 45042 5 1 1 45041
0 45043 7 1 2 94029 102085
0 45044 5 1 1 45043
0 45045 7 1 2 45042 45044
0 45046 5 1 1 45045
0 45047 7 1 2 67735 102074
0 45048 7 1 2 45046 45047
0 45049 5 1 1 45048
0 45050 7 1 2 45040 45049
0 45051 7 1 2 45036 45050
0 45052 5 1 1 45051
0 45053 7 1 2 87386 45052
0 45054 5 1 1 45053
0 45055 7 1 2 65210 45054
0 45056 7 1 2 45021 45055
0 45057 5 1 1 45056
0 45058 7 3 2 90618 93916
0 45059 7 1 2 78166 95068
0 45060 5 1 1 45059
0 45061 7 1 2 44984 45060
0 45062 5 1 1 45061
0 45063 7 1 2 74393 45062
0 45064 5 1 1 45063
0 45065 7 1 2 76825 101805
0 45066 5 1 1 45065
0 45067 7 1 2 45064 45066
0 45068 5 1 1 45067
0 45069 7 1 2 86143 45068
0 45070 5 1 1 45069
0 45071 7 1 2 83632 79961
0 45072 7 1 2 101788 45071
0 45073 5 1 1 45072
0 45074 7 1 2 45070 45073
0 45075 5 1 1 45074
0 45076 7 1 2 76190 45075
0 45077 5 1 1 45076
0 45078 7 1 2 77802 84083
0 45079 7 1 2 95809 45078
0 45080 7 1 2 99073 45079
0 45081 5 1 1 45080
0 45082 7 1 2 79962 82298
0 45083 7 1 2 99863 45082
0 45084 5 1 1 45083
0 45085 7 1 2 45081 45084
0 45086 5 1 1 45085
0 45087 7 1 2 98312 45086
0 45088 5 1 1 45087
0 45089 7 2 2 72078 86064
0 45090 5 1 1 102091
0 45091 7 1 2 94030 95617
0 45092 5 1 1 45091
0 45093 7 1 2 45090 45092
0 45094 5 2 1 45093
0 45095 7 2 2 79138 83398
0 45096 7 1 2 80995 102095
0 45097 7 1 2 102093 45096
0 45098 5 1 1 45097
0 45099 7 1 2 45088 45098
0 45100 7 1 2 45077 45099
0 45101 5 1 1 45100
0 45102 7 1 2 83152 45101
0 45103 5 1 1 45102
0 45104 7 2 2 75423 101162
0 45105 5 1 1 102097
0 45106 7 1 2 74381 86982
0 45107 5 1 1 45106
0 45108 7 1 2 23766 45107
0 45109 5 1 1 45108
0 45110 7 1 2 62447 85268
0 45111 7 1 2 45109 45110
0 45112 5 1 1 45111
0 45113 7 1 2 45105 45112
0 45114 5 1 1 45113
0 45115 7 1 2 85844 45114
0 45116 5 1 1 45115
0 45117 7 1 2 64180 90352
0 45118 7 1 2 87184 92296
0 45119 7 1 2 45117 45118
0 45120 5 1 1 45119
0 45121 7 1 2 45116 45120
0 45122 5 1 1 45121
0 45123 7 1 2 88706 45122
0 45124 5 1 1 45123
0 45125 7 1 2 66035 83823
0 45126 7 2 2 99074 45125
0 45127 7 1 2 80170 99060
0 45128 7 1 2 102099 45127
0 45129 5 1 1 45128
0 45130 7 1 2 45124 45129
0 45131 5 1 1 45130
0 45132 7 1 2 64979 45131
0 45133 5 1 1 45132
0 45134 7 2 2 85130 71443
0 45135 7 4 2 61659 80171
0 45136 5 1 1 102103
0 45137 7 1 2 102101 102104
0 45138 7 1 2 102100 45137
0 45139 5 1 1 45138
0 45140 7 1 2 45133 45139
0 45141 5 1 1 45140
0 45142 7 1 2 62635 45141
0 45143 5 1 1 45142
0 45144 7 1 2 89889 102098
0 45145 5 1 1 45144
0 45146 7 1 2 81942 87185
0 45147 5 1 1 45146
0 45148 7 1 2 10307 45147
0 45149 5 1 1 45148
0 45150 7 1 2 81833 77550
0 45151 7 1 2 89428 45150
0 45152 7 1 2 45149 45151
0 45153 5 1 1 45152
0 45154 7 1 2 45145 45153
0 45155 5 1 1 45154
0 45156 7 1 2 67524 45155
0 45157 5 1 1 45156
0 45158 7 1 2 71785 74711
0 45159 5 1 1 45158
0 45160 7 1 2 5360 45159
0 45161 5 2 1 45160
0 45162 7 1 2 89890 95684
0 45163 7 1 2 102107 45162
0 45164 5 1 1 45163
0 45165 7 1 2 45157 45164
0 45166 5 1 1 45165
0 45167 7 1 2 98313 45166
0 45168 5 1 1 45167
0 45169 7 1 2 84001 86246
0 45170 7 1 2 99085 45169
0 45171 5 1 1 45170
0 45172 7 1 2 84802 96089
0 45173 7 1 2 88878 45172
0 45174 7 1 2 97489 45173
0 45175 5 1 1 45174
0 45176 7 1 2 45171 45175
0 45177 5 1 1 45176
0 45178 7 1 2 71174 45177
0 45179 5 1 1 45178
0 45180 7 1 2 79083 90389
0 45181 7 1 2 81334 45180
0 45182 7 1 2 102108 45181
0 45183 5 1 1 45182
0 45184 7 1 2 45179 45183
0 45185 5 1 1 45184
0 45186 7 1 2 67525 45185
0 45187 5 1 1 45186
0 45188 7 2 2 79139 81849
0 45189 5 1 1 102109
0 45190 7 1 2 10222 45189
0 45191 5 1 1 45190
0 45192 7 1 2 88934 93931
0 45193 7 1 2 95659 45192
0 45194 7 1 2 62448 84375
0 45195 7 1 2 101899 45194
0 45196 7 1 2 45193 45195
0 45197 5 1 1 45196
0 45198 7 1 2 78303 102048
0 45199 5 1 1 45198
0 45200 7 1 2 89015 84197
0 45201 7 1 2 45199 45200
0 45202 5 1 1 45201
0 45203 7 1 2 45197 45202
0 45204 5 1 1 45203
0 45205 7 1 2 45191 45204
0 45206 5 1 1 45205
0 45207 7 1 2 88781 90010
0 45208 7 1 2 87186 100228
0 45209 7 1 2 98242 45208
0 45210 7 1 2 45207 45209
0 45211 5 1 1 45210
0 45212 7 1 2 70136 45211
0 45213 7 1 2 45206 45212
0 45214 7 1 2 45187 45213
0 45215 7 1 2 45168 45214
0 45216 7 1 2 45143 45215
0 45217 7 1 2 45103 45216
0 45218 5 1 1 45217
0 45219 7 1 2 102088 45218
0 45220 7 1 2 45057 45219
0 45221 5 1 1 45220
0 45222 7 1 2 81102 78481
0 45223 7 1 2 86799 97223
0 45224 7 1 2 45222 45223
0 45225 5 1 1 45224
0 45226 7 1 2 86920 92055
0 45227 7 2 2 79545 82903
0 45228 7 1 2 95460 102111
0 45229 7 1 2 45226 45228
0 45230 5 1 1 45229
0 45231 7 1 2 45225 45230
0 45232 5 1 1 45231
0 45233 7 1 2 99255 99918
0 45234 7 1 2 45232 45233
0 45235 5 1 1 45234
0 45236 7 1 2 45221 45235
0 45237 5 1 1 45236
0 45238 7 1 2 68715 45237
0 45239 5 1 1 45238
0 45240 7 1 2 95073 102056
0 45241 5 1 1 45240
0 45242 7 1 2 69840 45241
0 45243 5 1 1 45242
0 45244 7 1 2 101971 45243
0 45245 5 1 1 45244
0 45246 7 1 2 84020 45245
0 45247 5 1 1 45246
0 45248 7 3 2 78082 80301
0 45249 7 1 2 94259 102113
0 45250 5 1 1 45249
0 45251 7 1 2 45247 45250
0 45252 5 1 1 45251
0 45253 7 1 2 64181 45252
0 45254 5 1 1 45253
0 45255 7 2 2 74631 78609
0 45256 7 1 2 102070 102116
0 45257 5 1 1 45256
0 45258 7 1 2 62449 72724
0 45259 7 1 2 85767 45258
0 45260 7 1 2 89811 45259
0 45261 5 1 1 45260
0 45262 7 1 2 45257 45261
0 45263 5 1 1 45262
0 45264 7 1 2 74606 45263
0 45265 5 1 1 45264
0 45266 7 1 2 45254 45265
0 45267 5 1 1 45266
0 45268 7 1 2 68716 45267
0 45269 5 1 1 45268
0 45270 7 1 2 78558 102068
0 45271 5 1 1 45270
0 45272 7 1 2 82064 102046
0 45273 5 1 1 45272
0 45274 7 1 2 45271 45273
0 45275 5 1 1 45274
0 45276 7 1 2 74572 45275
0 45277 5 1 1 45276
0 45278 7 1 2 82072 101980
0 45279 5 1 1 45278
0 45280 7 1 2 64980 84306
0 45281 7 1 2 88054 45280
0 45282 5 1 1 45281
0 45283 7 1 2 45279 45282
0 45284 5 1 1 45283
0 45285 7 1 2 76978 45284
0 45286 5 1 1 45285
0 45287 7 1 2 78610 84021
0 45288 7 1 2 89101 45287
0 45289 5 1 1 45288
0 45290 7 1 2 72581 90899
0 45291 7 1 2 102071 45290
0 45292 5 1 1 45291
0 45293 7 1 2 45289 45292
0 45294 5 1 1 45293
0 45295 7 1 2 62203 45294
0 45296 5 1 1 45295
0 45297 7 1 2 45286 45296
0 45298 7 1 2 45277 45297
0 45299 7 1 2 45269 45298
0 45300 5 1 1 45299
0 45301 7 1 2 90269 45300
0 45302 5 1 1 45301
0 45303 7 1 2 86424 101905
0 45304 5 1 1 45303
0 45305 7 1 2 67736 83975
0 45306 5 1 1 45305
0 45307 7 1 2 14315 92624
0 45308 5 2 1 45307
0 45309 7 1 2 45306 102118
0 45310 7 1 2 45304 45309
0 45311 5 1 1 45310
0 45312 7 1 2 75237 91767
0 45313 7 1 2 97290 45312
0 45314 5 1 1 45313
0 45315 7 1 2 90245 93667
0 45316 7 1 2 74594 45315
0 45317 5 1 1 45316
0 45318 7 1 2 45314 45317
0 45319 7 1 2 45311 45318
0 45320 5 1 1 45319
0 45321 7 1 2 65211 45320
0 45322 5 1 1 45321
0 45323 7 1 2 75968 81569
0 45324 7 1 2 90510 45323
0 45325 5 1 1 45324
0 45326 7 1 2 45322 45325
0 45327 5 1 1 45326
0 45328 7 1 2 69841 45327
0 45329 5 1 1 45328
0 45330 7 1 2 73034 102114
0 45331 7 1 2 102119 45330
0 45332 5 1 1 45331
0 45333 7 1 2 45329 45332
0 45334 5 1 1 45333
0 45335 7 1 2 98314 45334
0 45336 5 1 1 45335
0 45337 7 1 2 94418 102000
0 45338 5 1 1 45337
0 45339 7 1 2 94984 95871
0 45340 5 1 1 45339
0 45341 7 1 2 45338 45340
0 45342 5 1 1 45341
0 45343 7 1 2 90225 45342
0 45344 5 1 1 45343
0 45345 7 1 2 90270 101958
0 45346 5 1 1 45345
0 45347 7 1 2 45344 45346
0 45348 5 1 1 45347
0 45349 7 1 2 74552 45348
0 45350 5 1 1 45349
0 45351 7 1 2 101558 101901
0 45352 5 1 1 45351
0 45353 7 1 2 89544 91157
0 45354 5 1 1 45353
0 45355 7 1 2 72725 74041
0 45356 7 1 2 86918 45355
0 45357 5 1 1 45356
0 45358 7 1 2 45354 45357
0 45359 5 1 1 45358
0 45360 7 1 2 69047 45359
0 45361 5 1 1 45360
0 45362 7 1 2 90123 85484
0 45363 5 1 1 45362
0 45364 7 1 2 72646 75823
0 45365 7 1 2 76967 45364
0 45366 5 1 1 45365
0 45367 7 1 2 45363 45366
0 45368 5 1 1 45367
0 45369 7 1 2 67526 45368
0 45370 5 1 1 45369
0 45371 7 1 2 45361 45370
0 45372 5 1 1 45371
0 45373 7 1 2 69842 45372
0 45374 5 1 1 45373
0 45375 7 1 2 45352 45374
0 45376 5 1 1 45375
0 45377 7 1 2 67309 45376
0 45378 5 1 1 45377
0 45379 7 1 2 71497 102115
0 45380 7 1 2 101543 45379
0 45381 5 1 1 45380
0 45382 7 1 2 45378 45381
0 45383 5 1 1 45382
0 45384 7 1 2 83962 45383
0 45385 5 1 1 45384
0 45386 7 1 2 45350 45385
0 45387 7 1 2 45336 45386
0 45388 7 1 2 45302 45387
0 45389 5 1 1 45388
0 45390 7 1 2 102089 45389
0 45391 5 1 1 45390
0 45392 7 2 2 79268 99166
0 45393 7 2 2 82078 96062
0 45394 7 1 2 102120 102122
0 45395 5 1 1 45394
0 45396 7 2 2 82904 95143
0 45397 7 1 2 95555 102124
0 45398 5 1 1 45397
0 45399 7 1 2 45395 45398
0 45400 5 1 1 45399
0 45401 7 1 2 93967 45400
0 45402 5 1 1 45401
0 45403 7 1 2 74382 90223
0 45404 7 1 2 86382 45403
0 45405 7 1 2 95382 45404
0 45406 7 1 2 101869 45405
0 45407 5 1 1 45406
0 45408 7 1 2 45402 45407
0 45409 5 1 1 45408
0 45410 7 1 2 70137 45409
0 45411 5 1 1 45410
0 45412 7 2 2 78611 82813
0 45413 7 1 2 93065 99795
0 45414 7 1 2 98315 45413
0 45415 7 1 2 102126 45414
0 45416 7 1 2 102083 45415
0 45417 5 1 1 45416
0 45418 7 1 2 45411 45417
0 45419 5 1 1 45418
0 45420 7 1 2 62892 45419
0 45421 5 1 1 45420
0 45422 7 1 2 87619 102094
0 45423 5 1 1 45422
0 45424 7 1 2 85623 101920
0 45425 5 1 1 45424
0 45426 7 1 2 101893 45425
0 45427 5 1 1 45426
0 45428 7 1 2 74666 73672
0 45429 5 1 1 45428
0 45430 7 1 2 45427 45429
0 45431 5 1 1 45430
0 45432 7 1 2 78612 45431
0 45433 5 1 1 45432
0 45434 7 1 2 45423 45433
0 45435 5 1 1 45434
0 45436 7 1 2 95096 45435
0 45437 5 1 1 45436
0 45438 7 2 2 64182 79269
0 45439 7 1 2 84452 102128
0 45440 7 2 2 65524 82079
0 45441 7 1 2 99473 102130
0 45442 7 1 2 45439 45441
0 45443 5 1 1 45442
0 45444 7 1 2 68717 45443
0 45445 7 1 2 45437 45444
0 45446 7 1 2 45421 45445
0 45447 5 1 1 45446
0 45448 7 1 2 90353 102064
0 45449 5 1 1 45448
0 45450 7 2 2 82202 89812
0 45451 5 1 1 102132
0 45452 7 1 2 100988 102133
0 45453 5 1 1 45452
0 45454 7 1 2 45449 45453
0 45455 5 1 1 45454
0 45456 7 1 2 67527 45455
0 45457 5 1 1 45456
0 45458 7 1 2 90354 94985
0 45459 5 1 1 45458
0 45460 7 1 2 45451 45459
0 45461 5 1 1 45460
0 45462 7 1 2 101792 45461
0 45463 5 1 1 45462
0 45464 7 1 2 45457 45463
0 45465 5 1 1 45464
0 45466 7 1 2 95097 45465
0 45467 5 1 1 45466
0 45468 7 1 2 86617 81861
0 45469 7 1 2 84754 94727
0 45470 7 1 2 45468 45469
0 45471 5 1 1 45470
0 45472 7 1 2 63849 45471
0 45473 7 1 2 45467 45472
0 45474 5 1 1 45473
0 45475 7 1 2 93812 45474
0 45476 7 1 2 45447 45475
0 45477 5 1 1 45476
0 45478 7 1 2 45391 45477
0 45479 5 1 1 45478
0 45480 7 1 2 90199 45479
0 45481 5 1 1 45480
0 45482 7 2 2 77581 84488
0 45483 7 1 2 81103 102134
0 45484 5 1 1 45483
0 45485 7 1 2 88950 89550
0 45486 7 1 2 90460 45485
0 45487 5 1 1 45486
0 45488 7 1 2 45484 45487
0 45489 5 1 1 45488
0 45490 7 1 2 84198 45489
0 45491 5 1 1 45490
0 45492 7 1 2 80302 96601
0 45493 7 1 2 93209 45492
0 45494 5 1 1 45493
0 45495 7 1 2 45491 45494
0 45496 5 1 1 45495
0 45497 7 1 2 69625 45496
0 45498 5 1 1 45497
0 45499 7 2 2 70437 101530
0 45500 7 1 2 76826 102136
0 45501 5 1 1 45500
0 45502 7 1 2 76783 89620
0 45503 5 1 1 45502
0 45504 7 1 2 45501 45503
0 45505 5 1 1 45504
0 45506 7 1 2 61908 45505
0 45507 5 1 1 45506
0 45508 7 1 2 74712 102102
0 45509 5 1 1 45508
0 45510 7 1 2 45507 45509
0 45511 5 1 1 45510
0 45512 7 1 2 91786 94651
0 45513 7 1 2 45511 45512
0 45514 5 1 1 45513
0 45515 7 1 2 45498 45514
0 45516 5 1 1 45515
0 45517 7 1 2 102090 45516
0 45518 5 1 1 45517
0 45519 7 2 2 82517 92854
0 45520 5 1 1 102138
0 45521 7 3 2 82080 88130
0 45522 7 1 2 87563 94377
0 45523 7 1 2 99025 45522
0 45524 7 1 2 102140 45523
0 45525 7 1 2 102139 45524
0 45526 5 1 1 45525
0 45527 7 1 2 45518 45526
0 45528 5 1 1 45527
0 45529 7 1 2 70138 45528
0 45530 5 1 1 45529
0 45531 7 2 2 91284 93917
0 45532 7 2 2 80655 90619
0 45533 7 1 2 102143 102145
0 45534 7 1 2 102075 45533
0 45535 7 1 2 102022 45534
0 45536 5 1 1 45535
0 45537 7 1 2 45530 45536
0 45538 5 1 1 45537
0 45539 7 1 2 68718 45538
0 45540 5 1 1 45539
0 45541 7 1 2 87052 96049
0 45542 7 1 2 102137 45541
0 45543 5 1 1 45542
0 45544 7 1 2 102026 45543
0 45545 5 1 1 45544
0 45546 7 1 2 82353 93918
0 45547 7 1 2 102146 45546
0 45548 7 1 2 45545 45547
0 45549 5 1 1 45548
0 45550 7 1 2 45540 45549
0 45551 5 1 1 45550
0 45552 7 1 2 72647 45551
0 45553 5 1 1 45552
0 45554 7 1 2 79084 100627
0 45555 7 1 2 86460 45554
0 45556 7 1 2 99214 45555
0 45557 5 1 1 45556
0 45558 7 2 2 92224 98161
0 45559 5 1 1 102147
0 45560 7 2 2 63397 80509
0 45561 7 1 2 94616 102149
0 45562 5 1 1 45561
0 45563 7 1 2 45559 45562
0 45564 5 1 1 45563
0 45565 7 1 2 86983 93813
0 45566 7 1 2 45564 45565
0 45567 5 1 1 45566
0 45568 7 1 2 45557 45567
0 45569 5 1 1 45568
0 45570 7 1 2 72079 45569
0 45571 5 1 1 45570
0 45572 7 1 2 94689 96347
0 45573 5 1 1 45572
0 45574 7 3 2 64981 96063
0 45575 7 2 2 95428 102151
0 45576 7 1 2 92499 102154
0 45577 5 1 1 45576
0 45578 7 1 2 45573 45577
0 45579 5 1 1 45578
0 45580 7 1 2 72648 99098
0 45581 7 1 2 45579 45580
0 45582 5 1 1 45581
0 45583 7 1 2 45571 45582
0 45584 5 1 1 45583
0 45585 7 1 2 76919 45584
0 45586 5 1 1 45585
0 45587 7 1 2 64388 89869
0 45588 7 2 2 66290 90011
0 45589 7 1 2 102066 102156
0 45590 7 1 2 101505 45589
0 45591 7 1 2 45587 45590
0 45592 5 1 1 45591
0 45593 7 1 2 45586 45592
0 45594 5 1 1 45593
0 45595 7 1 2 75837 45594
0 45596 5 1 1 45595
0 45597 7 1 2 45553 45596
0 45598 7 1 2 45481 45597
0 45599 7 1 2 45239 45598
0 45600 7 1 2 44918 45599
0 45601 7 1 2 44656 45600
0 45602 5 1 1 45601
0 45603 7 1 2 93871 45602
0 45604 5 1 1 45603
0 45605 7 1 2 81943 85398
0 45606 5 1 1 45605
0 45607 7 2 2 61660 72793
0 45608 7 1 2 76947 78809
0 45609 7 1 2 102158 45608
0 45610 5 1 1 45609
0 45611 7 1 2 45606 45610
0 45612 5 1 1 45611
0 45613 7 1 2 62636 45612
0 45614 5 1 1 45613
0 45615 7 2 2 64793 98316
0 45616 7 1 2 61661 102160
0 45617 5 1 1 45616
0 45618 7 1 2 84767 95600
0 45619 5 1 1 45618
0 45620 7 1 2 87015 17210
0 45621 5 3 1 45620
0 45622 7 1 2 71175 102162
0 45623 5 1 1 45622
0 45624 7 1 2 45619 45623
0 45625 7 1 2 45617 45624
0 45626 5 1 1 45625
0 45627 7 1 2 92418 45626
0 45628 5 1 1 45627
0 45629 7 1 2 45614 45628
0 45630 5 1 1 45629
0 45631 7 1 2 71066 45630
0 45632 5 1 1 45631
0 45633 7 1 2 92037 92419
0 45634 7 1 2 100989 45633
0 45635 5 1 1 45634
0 45636 7 1 2 45632 45635
0 45637 5 1 1 45636
0 45638 7 1 2 93872 99723
0 45639 7 1 2 45637 45638
0 45640 5 1 1 45639
0 45641 7 1 2 71067 101650
0 45642 5 1 1 45641
0 45643 7 1 2 75599 101839
0 45644 5 1 1 45643
0 45645 7 1 2 45642 45644
0 45646 5 1 1 45645
0 45647 7 1 2 81944 45646
0 45648 5 1 1 45647
0 45649 7 1 2 100229 101651
0 45650 5 1 1 45649
0 45651 7 1 2 89026 45650
0 45652 5 1 1 45651
0 45653 7 1 2 86984 45652
0 45654 5 1 1 45653
0 45655 7 1 2 45648 45654
0 45656 5 1 1 45655
0 45657 7 1 2 69048 45656
0 45658 5 1 1 45657
0 45659 7 2 2 69626 71481
0 45660 7 1 2 66552 102165
0 45661 5 1 1 45660
0 45662 7 1 2 92040 45661
0 45663 5 1 1 45662
0 45664 7 1 2 101610 45663
0 45665 5 1 1 45664
0 45666 7 1 2 92051 101704
0 45667 5 1 1 45666
0 45668 7 1 2 87896 91582
0 45669 5 1 1 45668
0 45670 7 1 2 66776 75677
0 45671 7 1 2 91231 45670
0 45672 5 1 1 45671
0 45673 7 1 2 45669 45672
0 45674 5 1 1 45673
0 45675 7 1 2 66036 45674
0 45676 5 1 1 45675
0 45677 7 1 2 45667 45676
0 45678 7 1 2 45665 45677
0 45679 7 1 2 45658 45678
0 45680 5 1 1 45679
0 45681 7 1 2 76901 91373
0 45682 7 1 2 99740 45681
0 45683 7 1 2 45680 45682
0 45684 5 1 1 45683
0 45685 7 1 2 45640 45684
0 45686 5 1 1 45685
0 45687 7 1 2 64294 45686
0 45688 5 1 1 45687
0 45689 7 1 2 92052 101681
0 45690 5 1 1 45689
0 45691 7 1 2 89436 101572
0 45692 5 1 1 45691
0 45693 7 1 2 91073 45692
0 45694 5 1 1 45693
0 45695 7 1 2 86985 45694
0 45696 5 1 1 45695
0 45697 7 1 2 45690 45696
0 45698 5 1 1 45697
0 45699 7 2 2 99965 97462
0 45700 7 1 2 79537 97788
0 45701 7 1 2 102167 45700
0 45702 7 1 2 45698 45701
0 45703 5 1 1 45702
0 45704 7 1 2 45688 45703
0 45705 5 1 1 45704
0 45706 7 1 2 69247 45705
0 45707 5 1 1 45706
0 45708 7 1 2 82649 100701
0 45709 5 1 1 45708
0 45710 7 2 2 81945 100823
0 45711 5 2 1 102169
0 45712 7 1 2 45709 102171
0 45713 5 2 1 45712
0 45714 7 1 2 72188 102173
0 45715 5 1 1 45714
0 45716 7 1 2 101778 100806
0 45717 5 1 1 45716
0 45718 7 1 2 45715 45717
0 45719 5 1 1 45718
0 45720 7 1 2 77037 45719
0 45721 5 1 1 45720
0 45722 7 1 2 91879 95560
0 45723 7 1 2 96752 45722
0 45724 7 1 2 101573 45723
0 45725 5 1 1 45724
0 45726 7 1 2 45721 45725
0 45727 5 1 1 45726
0 45728 7 1 2 70438 97993
0 45729 7 1 2 45727 45728
0 45730 5 1 1 45729
0 45731 7 2 2 88131 88169
0 45732 7 1 2 90450 102175
0 45733 7 1 2 100429 45732
0 45734 5 1 1 45733
0 45735 7 1 2 45730 45734
0 45736 5 1 1 45735
0 45737 7 1 2 66148 45736
0 45738 5 1 1 45737
0 45739 7 1 2 72189 93604
0 45740 5 1 1 45739
0 45741 7 1 2 85845 93641
0 45742 5 1 1 45741
0 45743 7 1 2 45740 45742
0 45744 5 1 1 45743
0 45745 7 1 2 91521 93708
0 45746 7 1 2 100729 45745
0 45747 7 1 2 45744 45746
0 45748 5 1 1 45747
0 45749 7 1 2 45738 45748
0 45750 5 1 1 45749
0 45751 7 1 2 100230 45750
0 45752 5 1 1 45751
0 45753 7 2 2 72855 92053
0 45754 7 1 2 99329 102177
0 45755 5 1 1 45754
0 45756 7 1 2 67737 76565
0 45757 7 1 2 97490 45756
0 45758 7 1 2 98527 45757
0 45759 5 1 1 45758
0 45760 7 1 2 45755 45759
0 45761 5 1 1 45760
0 45762 7 1 2 72190 45761
0 45763 5 1 1 45762
0 45764 7 1 2 74632 96969
0 45765 7 1 2 71103 45764
0 45766 5 1 1 45765
0 45767 7 1 2 75258 95495
0 45768 7 1 2 100494 45767
0 45769 5 1 1 45768
0 45770 7 1 2 45766 45769
0 45771 5 1 1 45770
0 45772 7 1 2 81946 45771
0 45773 5 1 1 45772
0 45774 7 1 2 45763 45773
0 45775 5 1 1 45774
0 45776 7 1 2 82940 100363
0 45777 7 1 2 45775 45776
0 45778 5 1 1 45777
0 45779 7 1 2 45752 45778
0 45780 7 1 2 45707 45779
0 45781 5 1 1 45780
0 45782 7 1 2 45781 98461
0 45783 5 1 1 45782
0 45784 7 2 2 83424 93149
0 45785 7 1 2 75424 98108
0 45786 7 1 2 102179 45785
0 45787 5 1 1 45786
0 45788 7 1 2 89578 924
0 45789 5 2 1 45788
0 45790 7 1 2 96420 98394
0 45791 7 1 2 102181 45790
0 45792 5 1 1 45791
0 45793 7 1 2 45787 45792
0 45794 5 1 1 45793
0 45795 7 1 2 67812 45794
0 45796 5 1 1 45795
0 45797 7 1 2 62979 84084
0 45798 7 1 2 93195 98496
0 45799 7 1 2 45797 45798
0 45800 7 1 2 96773 45799
0 45801 5 1 1 45800
0 45802 7 1 2 45796 45801
0 45803 5 1 1 45802
0 45804 7 1 2 66149 45803
0 45805 5 1 1 45804
0 45806 7 2 2 91831 91867
0 45807 7 2 2 61314 82635
0 45808 7 1 2 93150 102185
0 45809 7 1 2 102183 45808
0 45810 5 1 1 45809
0 45811 7 1 2 45805 45810
0 45812 5 1 1 45811
0 45813 7 1 2 95318 45812
0 45814 5 1 1 45813
0 45815 7 1 2 100231 98109
0 45816 7 1 2 101045 100740
0 45817 7 1 2 45815 45816
0 45818 5 1 1 45817
0 45819 7 1 2 45814 45818
0 45820 5 1 1 45819
0 45821 7 1 2 61662 45820
0 45822 5 1 1 45821
0 45823 7 6 2 67813 64573
0 45824 7 1 2 67738 102187
0 45825 7 1 2 100111 45824
0 45826 5 1 1 45825
0 45827 7 1 2 93130 98451
0 45828 5 1 1 45827
0 45829 7 1 2 45826 45828
0 45830 5 1 1 45829
0 45831 7 1 2 88043 45830
0 45832 5 1 1 45831
0 45833 7 1 2 74473 82081
0 45834 7 1 2 100611 45833
0 45835 5 1 1 45834
0 45836 7 1 2 45832 45835
0 45837 5 1 1 45836
0 45838 7 1 2 66150 45837
0 45839 5 1 1 45838
0 45840 7 1 2 82905 91868
0 45841 7 1 2 99558 45840
0 45842 5 1 1 45841
0 45843 7 1 2 45839 45842
0 45844 5 1 1 45843
0 45845 7 1 2 92902 95319
0 45846 7 1 2 45844 45845
0 45847 5 1 1 45846
0 45848 7 1 2 45822 45847
0 45849 5 1 1 45848
0 45850 7 1 2 66291 45849
0 45851 5 1 1 45850
0 45852 7 2 2 82082 93699
0 45853 7 1 2 100106 102193
0 45854 5 1 1 45853
0 45855 7 1 2 101685 36554
0 45856 5 4 1 45855
0 45857 7 1 2 88044 102195
0 45858 5 1 1 45857
0 45859 7 1 2 45854 45858
0 45860 5 1 1 45859
0 45861 7 1 2 92912 45860
0 45862 5 1 1 45861
0 45863 7 1 2 83699 92855
0 45864 7 1 2 102180 45863
0 45865 5 1 1 45864
0 45866 7 1 2 45862 45865
0 45867 5 1 1 45866
0 45868 7 1 2 101457 45867
0 45869 5 1 1 45868
0 45870 7 11 2 99796 98116
0 45871 7 1 2 74444 92809
0 45872 7 1 2 89838 45871
0 45873 7 1 2 102199 45872
0 45874 5 1 1 45873
0 45875 7 1 2 45869 45874
0 45876 5 1 1 45875
0 45877 7 1 2 90999 45876
0 45878 5 1 1 45877
0 45879 7 1 2 45851 45878
0 45880 5 1 1 45879
0 45881 7 1 2 64794 45880
0 45882 5 1 1 45881
0 45883 7 1 2 71471 82923
0 45884 7 4 2 61315 91880
0 45885 7 1 2 102210 98166
0 45886 7 1 2 45883 45885
0 45887 5 1 1 45886
0 45888 7 1 2 91309 93814
0 45889 5 1 1 45888
0 45890 7 1 2 92200 98390
0 45891 5 1 1 45890
0 45892 7 1 2 45889 45891
0 45893 5 4 1 45892
0 45894 7 1 2 67814 102214
0 45895 5 1 1 45894
0 45896 7 1 2 101859 98455
0 45897 5 1 1 45896
0 45898 7 1 2 45895 45897
0 45899 5 1 1 45898
0 45900 7 1 2 66151 45899
0 45901 5 1 1 45900
0 45902 7 1 2 93071 93692
0 45903 5 1 1 45902
0 45904 7 1 2 45901 45903
0 45905 5 1 1 45904
0 45906 7 1 2 95320 102182
0 45907 7 1 2 45905 45906
0 45908 5 1 1 45907
0 45909 7 1 2 45887 45908
0 45910 5 1 1 45909
0 45911 7 1 2 96104 45910
0 45912 5 1 1 45911
0 45913 7 1 2 45882 45912
0 45914 5 1 1 45913
0 45915 7 1 2 70139 45914
0 45916 5 1 1 45915
0 45917 7 1 2 87365 101046
0 45918 5 1 1 45917
0 45919 7 1 2 69627 101458
0 45920 7 1 2 100631 45919
0 45921 5 1 1 45920
0 45922 7 1 2 45918 45921
0 45923 5 1 1 45922
0 45924 7 1 2 68475 45923
0 45925 5 1 1 45924
0 45926 7 1 2 63635 79971
0 45927 7 1 2 82096 45926
0 45928 7 1 2 100711 45927
0 45929 5 1 1 45928
0 45930 7 1 2 45925 45929
0 45931 5 1 1 45930
0 45932 7 1 2 98415 45931
0 45933 5 1 1 45932
0 45934 7 1 2 87901 97316
0 45935 5 1 1 45934
0 45936 7 1 2 38306 45935
0 45937 5 1 1 45936
0 45938 7 1 2 45937 100571
0 45939 5 1 1 45938
0 45940 7 2 2 96970 99114
0 45941 7 1 2 82591 102218
0 45942 5 1 1 45941
0 45943 7 1 2 45939 45942
0 45944 5 1 1 45943
0 45945 7 1 2 90200 45944
0 45946 5 1 1 45945
0 45947 7 1 2 68719 93873
0 45948 7 2 2 69628 91881
0 45949 7 1 2 98556 102220
0 45950 7 1 2 45947 45949
0 45951 7 1 2 99081 45950
0 45952 5 1 1 45951
0 45953 7 1 2 45946 45952
0 45954 7 1 2 45933 45953
0 45955 5 1 1 45954
0 45956 7 1 2 93131 45955
0 45957 5 1 1 45956
0 45958 7 1 2 92913 93815
0 45959 5 1 1 45958
0 45960 7 2 2 99026 98384
0 45961 7 2 2 82674 102222
0 45962 5 1 1 102224
0 45963 7 1 2 45959 45962
0 45964 5 1 1 45963
0 45965 7 1 2 83307 93047
0 45966 7 2 2 45964 45965
0 45967 7 1 2 87902 97994
0 45968 7 1 2 102226 45967
0 45969 5 1 1 45968
0 45970 7 1 2 45957 45969
0 45971 5 1 1 45970
0 45972 7 1 2 78613 45971
0 45973 5 1 1 45972
0 45974 7 1 2 62450 45973
0 45975 7 1 2 45916 45974
0 45976 5 1 1 45975
0 45977 7 6 2 64295 65212
0 45978 7 2 2 74893 102228
0 45979 7 1 2 96950 102234
0 45980 5 2 1 45979
0 45981 7 2 2 95348 98187
0 45982 7 1 2 66152 102238
0 45983 5 1 1 45982
0 45984 7 1 2 102236 45983
0 45985 5 1 1 45984
0 45986 7 1 2 100572 45985
0 45987 5 1 1 45986
0 45988 7 2 2 78115 98181
0 45989 7 1 2 98074 102240
0 45990 5 1 1 45989
0 45991 7 1 2 88179 102235
0 45992 5 1 1 45991
0 45993 7 1 2 45990 45992
0 45994 5 1 1 45993
0 45995 7 1 2 61316 45994
0 45996 5 1 1 45995
0 45997 7 1 2 78153 99973
0 45998 7 1 2 101298 45997
0 45999 5 1 1 45998
0 46000 7 1 2 45996 45999
0 46001 5 1 1 46000
0 46002 7 1 2 84411 46001
0 46003 5 1 1 46002
0 46004 7 1 2 45987 46003
0 46005 5 1 1 46004
0 46006 7 1 2 90201 46005
0 46007 5 1 1 46006
0 46008 7 1 2 102241 99376
0 46009 5 1 1 46008
0 46010 7 1 2 102237 46009
0 46011 5 1 1 46010
0 46012 7 1 2 87366 46011
0 46013 5 1 1 46012
0 46014 7 5 2 66553 67815
0 46015 7 2 2 102242 97635
0 46016 7 1 2 88303 102247
0 46017 7 1 2 88824 46016
0 46018 5 1 1 46017
0 46019 7 1 2 46013 46018
0 46020 5 1 1 46019
0 46021 7 1 2 98416 46020
0 46022 5 1 1 46021
0 46023 7 1 2 81947 95349
0 46024 5 1 1 46023
0 46025 7 1 2 74338 88645
0 46026 5 1 1 46025
0 46027 7 1 2 46024 46026
0 46028 5 1 1 46027
0 46029 7 1 2 91256 99256
0 46030 7 1 2 99430 46029
0 46031 7 1 2 46028 46030
0 46032 5 1 1 46031
0 46033 7 1 2 46022 46032
0 46034 7 1 2 46007 46033
0 46035 5 1 1 46034
0 46036 7 1 2 93132 46035
0 46037 5 1 1 46036
0 46038 7 1 2 102227 102239
0 46039 5 1 1 46038
0 46040 7 1 2 46037 46039
0 46041 5 1 1 46040
0 46042 7 1 2 69843 46041
0 46043 5 1 1 46042
0 46044 7 1 2 92856 96557
0 46045 5 1 1 46044
0 46046 7 1 2 99411 100939
0 46047 5 1 1 46046
0 46048 7 1 2 46045 46047
0 46049 5 1 1 46048
0 46050 7 1 2 82387 15605
0 46051 5 1 1 46050
0 46052 7 1 2 5495 43547
0 46053 7 1 2 46051 46052
0 46054 7 1 2 46049 46053
0 46055 5 1 1 46054
0 46056 7 1 2 87704 93816
0 46057 7 1 2 96470 46056
0 46058 5 1 1 46057
0 46059 7 1 2 61663 93753
0 46060 7 1 2 85328 46059
0 46061 7 1 2 96105 46060
0 46062 5 1 1 46061
0 46063 7 2 2 63036 75687
0 46064 7 1 2 81779 91882
0 46065 7 1 2 91852 46064
0 46066 7 1 2 102249 46065
0 46067 5 1 1 46066
0 46068 7 1 2 46062 46067
0 46069 7 1 2 46058 46068
0 46070 7 1 2 46055 46069
0 46071 5 1 1 46070
0 46072 7 1 2 67816 46071
0 46073 5 1 1 46072
0 46074 7 2 2 90675 97605
0 46075 7 1 2 91257 96106
0 46076 7 1 2 102251 46075
0 46077 5 1 1 46076
0 46078 7 1 2 46073 46077
0 46079 5 1 1 46078
0 46080 7 1 2 66153 46079
0 46081 5 1 1 46080
0 46082 7 2 2 95901 102211
0 46083 5 1 1 102253
0 46084 7 1 2 82749 98724
0 46085 7 1 2 102254 46084
0 46086 5 1 1 46085
0 46087 7 1 2 46081 46086
0 46088 5 2 1 46087
0 46089 7 1 2 78083 77093
0 46090 7 1 2 98182 46089
0 46091 7 1 2 102255 46090
0 46092 5 1 1 46091
0 46093 7 1 2 67310 46092
0 46094 7 1 2 46043 46093
0 46095 5 1 1 46094
0 46096 7 1 2 65525 46095
0 46097 7 1 2 45976 46096
0 46098 5 1 1 46097
0 46099 7 1 2 78633 86329
0 46100 5 6 1 46099
0 46101 7 1 2 101812 102257
0 46102 7 1 2 102256 46101
0 46103 5 1 1 46102
0 46104 7 1 2 96558 99211
0 46105 5 1 1 46104
0 46106 7 1 2 46083 46105
0 46107 5 1 1 46106
0 46108 7 3 2 64982 80574
0 46109 7 1 2 61909 102263
0 46110 5 1 1 46109
0 46111 7 1 2 9889 46110
0 46112 5 3 1 46111
0 46113 7 1 2 46107 102266
0 46114 5 1 1 46113
0 46115 7 3 2 91374 93133
0 46116 7 1 2 83506 87133
0 46117 7 1 2 102269 46116
0 46118 5 1 1 46117
0 46119 7 1 2 46114 46118
0 46120 5 1 1 46119
0 46121 7 1 2 74829 102184
0 46122 7 1 2 46120 46121
0 46123 5 1 1 46122
0 46124 7 1 2 46103 46123
0 46125 5 1 1 46124
0 46126 7 1 2 69136 46125
0 46127 5 1 1 46126
0 46128 7 1 2 61664 98395
0 46129 5 1 1 46128
0 46130 7 1 2 90202 101696
0 46131 5 1 1 46130
0 46132 7 1 2 46129 46131
0 46133 5 1 1 46132
0 46134 7 1 2 61400 46133
0 46135 5 1 1 46134
0 46136 7 1 2 61665 98412
0 46137 5 1 1 46136
0 46138 7 1 2 46135 46137
0 46139 5 1 1 46138
0 46140 7 2 2 64795 46139
0 46141 7 1 2 87620 102272
0 46142 5 1 1 46141
0 46143 7 1 2 90940 102215
0 46144 5 1 1 46143
0 46145 7 1 2 46142 46144
0 46146 5 1 1 46145
0 46147 7 1 2 91901 100750
0 46148 7 1 2 46146 46147
0 46149 5 1 1 46148
0 46150 7 1 2 46127 46149
0 46151 5 1 1 46150
0 46152 7 1 2 70439 46151
0 46153 5 1 1 46152
0 46154 7 2 2 81797 78681
0 46155 5 2 1 102274
0 46156 7 3 2 83598 81901
0 46157 5 1 1 102278
0 46158 7 1 2 102276 46157
0 46159 5 10 1 46158
0 46160 7 2 2 97789 102281
0 46161 7 1 2 92645 102291
0 46162 5 1 1 46161
0 46163 7 3 2 79085 78419
0 46164 7 1 2 98528 102293
0 46165 5 1 1 46164
0 46166 7 1 2 46162 46165
0 46167 5 1 1 46166
0 46168 7 1 2 100761 46167
0 46169 5 1 1 46168
0 46170 7 1 2 93874 101875
0 46171 7 1 2 102292 46170
0 46172 5 1 1 46171
0 46173 7 1 2 46169 46172
0 46174 5 1 1 46173
0 46175 7 1 2 93134 46174
0 46176 5 1 1 46175
0 46177 7 1 2 64983 96465
0 46178 7 1 2 99385 46177
0 46179 7 1 2 101033 46178
0 46180 5 1 1 46179
0 46181 7 1 2 46176 46180
0 46182 5 1 1 46181
0 46183 7 1 2 101813 46182
0 46184 5 1 1 46183
0 46185 7 3 2 64389 100002
0 46186 7 3 2 80996 100841
0 46187 7 1 2 98042 102299
0 46188 5 1 1 46187
0 46189 7 1 2 70440 102200
0 46190 5 1 1 46189
0 46191 7 1 2 46188 46190
0 46192 5 2 1 46191
0 46193 7 1 2 61317 102302
0 46194 5 1 1 46193
0 46195 7 1 2 101105 100590
0 46196 5 1 1 46195
0 46197 7 1 2 46194 46196
0 46198 5 1 1 46197
0 46199 7 1 2 97169 46198
0 46200 5 1 1 46199
0 46201 7 6 2 67046 69137
0 46202 7 1 2 91702 102304
0 46203 7 1 2 99864 46202
0 46204 7 1 2 100603 46203
0 46205 5 1 1 46204
0 46206 7 1 2 46200 46205
0 46207 5 1 1 46206
0 46208 7 1 2 102296 46207
0 46209 5 1 1 46208
0 46210 7 1 2 100511 36292
0 46211 5 2 1 46210
0 46212 7 1 2 97170 102310
0 46213 5 1 1 46212
0 46214 7 1 2 99377 99884
0 46215 5 1 1 46214
0 46216 7 1 2 46213 46215
0 46217 5 1 1 46216
0 46218 7 1 2 100689 46217
0 46219 5 1 1 46218
0 46220 7 1 2 96413 102188
0 46221 7 1 2 99167 46220
0 46222 7 3 2 76902 79140
0 46223 7 1 2 102312 97782
0 46224 7 1 2 46221 46223
0 46225 5 1 1 46224
0 46226 7 1 2 46219 46225
0 46227 5 1 1 46226
0 46228 7 1 2 100674 46227
0 46229 5 1 1 46228
0 46230 7 4 2 81348 82906
0 46231 7 1 2 93167 102315
0 46232 5 1 1 46231
0 46233 7 1 2 92935 96931
0 46234 5 1 1 46233
0 46235 7 1 2 46232 46234
0 46236 5 1 1 46235
0 46237 7 1 2 46236 100508
0 46238 5 1 1 46237
0 46239 7 1 2 101014 102141
0 46240 7 1 2 95350 46239
0 46241 5 1 1 46240
0 46242 7 1 2 46238 46241
0 46243 5 1 1 46242
0 46244 7 1 2 67739 46243
0 46245 5 1 1 46244
0 46246 7 1 2 92646 99168
0 46247 7 1 2 93253 46246
0 46248 7 1 2 97161 46247
0 46249 5 1 1 46248
0 46250 7 1 2 46245 46249
0 46251 5 1 1 46250
0 46252 7 1 2 99386 46251
0 46253 5 1 1 46252
0 46254 7 1 2 102313 102121
0 46255 7 1 2 100800 101331
0 46256 7 1 2 46254 46255
0 46257 5 1 1 46256
0 46258 7 1 2 46253 46257
0 46259 7 1 2 46229 46258
0 46260 7 1 2 46209 46259
0 46261 5 1 1 46260
0 46262 7 1 2 73035 46261
0 46263 5 1 1 46262
0 46264 7 1 2 46184 46263
0 46265 5 1 1 46264
0 46266 7 1 2 83153 46265
0 46267 5 1 1 46266
0 46268 7 3 2 69138 93135
0 46269 7 2 2 92838 102319
0 46270 7 1 2 102178 102322
0 46271 5 1 1 46270
0 46272 7 1 2 61910 80795
0 46273 7 1 2 80514 46272
0 46274 7 1 2 100836 46273
0 46275 5 1 1 46274
0 46276 7 1 2 46271 46275
0 46277 5 1 1 46276
0 46278 7 1 2 70140 46277
0 46279 5 1 1 46278
0 46280 7 1 2 100232 98584
0 46281 7 1 2 101245 100648
0 46282 7 1 2 46280 46281
0 46283 5 1 1 46282
0 46284 7 1 2 46279 46283
0 46285 5 1 1 46284
0 46286 7 1 2 98458 46285
0 46287 5 1 1 46286
0 46288 7 1 2 46267 46287
0 46289 7 1 2 46153 46288
0 46290 7 1 2 46098 46289
0 46291 5 1 1 46290
0 46292 7 1 2 72191 46291
0 46293 5 1 1 46292
0 46294 7 1 2 45783 46293
0 46295 7 1 2 45604 46294
0 46296 7 1 2 44319 46295
0 46297 7 1 2 43389 46296
0 46298 5 1 1 46297
0 46299 7 1 2 101509 46298
0 46300 5 1 1 46299
0 46301 7 3 2 68041 93817
0 46302 7 1 2 84827 94546
0 46303 5 1 1 46302
0 46304 7 1 2 75486 87513
0 46305 5 1 1 46304
0 46306 7 1 2 46303 46305
0 46307 5 1 1 46306
0 46308 7 1 2 96971 46307
0 46309 5 1 1 46308
0 46310 7 3 2 65526 80575
0 46311 7 1 2 89287 76214
0 46312 7 1 2 101056 46311
0 46313 7 1 2 102327 46312
0 46314 5 1 1 46313
0 46315 7 1 2 46309 46314
0 46316 5 1 1 46315
0 46317 7 1 2 76526 46316
0 46318 5 1 1 46317
0 46319 7 1 2 79046 101418
0 46320 5 1 1 46319
0 46321 7 1 2 72794 46320
0 46322 5 1 1 46321
0 46323 7 2 2 76903 84687
0 46324 5 1 1 102330
0 46325 7 1 2 70754 102331
0 46326 5 1 1 46325
0 46327 7 1 2 46322 46326
0 46328 5 1 1 46327
0 46329 7 1 2 96972 46328
0 46330 5 1 1 46329
0 46331 7 1 2 72795 97025
0 46332 5 1 1 46331
0 46333 7 1 2 71743 84688
0 46334 5 1 1 46333
0 46335 7 1 2 46332 46334
0 46336 5 1 1 46335
0 46337 7 1 2 80576 97317
0 46338 7 1 2 46336 46337
0 46339 5 1 1 46338
0 46340 7 1 2 46330 46339
0 46341 5 1 1 46340
0 46342 7 1 2 94547 46341
0 46343 5 1 1 46342
0 46344 7 1 2 46318 46343
0 46345 5 1 1 46344
0 46346 7 1 2 68720 46345
0 46347 5 1 1 46346
0 46348 7 2 2 62980 84424
0 46349 7 1 2 93950 102229
0 46350 7 1 2 102332 46349
0 46351 7 1 2 96376 46350
0 46352 5 1 1 46351
0 46353 7 1 2 46347 46352
0 46354 5 1 1 46353
0 46355 7 1 2 69248 46354
0 46356 5 1 1 46355
0 46357 7 2 2 80577 93875
0 46358 7 1 2 67311 90922
0 46359 5 1 1 46358
0 46360 7 1 2 97952 46359
0 46361 5 1 1 46360
0 46362 7 1 2 86888 46361
0 46363 5 1 1 46362
0 46364 7 1 2 89984 76435
0 46365 7 1 2 84891 46364
0 46366 5 1 1 46365
0 46367 7 1 2 46363 46366
0 46368 5 1 1 46367
0 46369 7 1 2 68476 46368
0 46370 5 1 1 46369
0 46371 7 1 2 93986 19406
0 46372 5 1 1 46371
0 46373 7 1 2 101563 46372
0 46374 5 1 1 46373
0 46375 7 1 2 46370 46374
0 46376 5 1 1 46375
0 46377 7 1 2 102334 46376
0 46378 5 1 1 46377
0 46379 7 1 2 86889 95083
0 46380 5 1 1 46379
0 46381 7 1 2 88830 94587
0 46382 5 1 1 46381
0 46383 7 1 2 46380 46382
0 46384 5 1 1 46383
0 46385 7 1 2 70441 46384
0 46386 5 1 1 46385
0 46387 7 1 2 76405 96343
0 46388 5 1 1 46387
0 46389 7 1 2 62451 87157
0 46390 5 2 1 46389
0 46391 7 2 2 65527 102336
0 46392 7 1 2 63636 102338
0 46393 5 1 1 46392
0 46394 7 1 2 46388 46393
0 46395 5 1 1 46394
0 46396 7 1 2 65847 46395
0 46397 5 1 1 46396
0 46398 7 1 2 71264 101757
0 46399 5 1 1 46398
0 46400 7 1 2 46397 46399
0 46401 5 1 1 46400
0 46402 7 1 2 63850 46401
0 46403 5 1 1 46402
0 46404 7 1 2 72390 75457
0 46405 7 1 2 95476 46404
0 46406 5 1 1 46405
0 46407 7 1 2 46403 46406
0 46408 5 1 1 46407
0 46409 7 1 2 77382 46408
0 46410 5 1 1 46409
0 46411 7 1 2 46386 46410
0 46412 5 1 1 46411
0 46413 7 1 2 66777 93876
0 46414 7 1 2 46412 46413
0 46415 5 1 1 46414
0 46416 7 1 2 46378 46415
0 46417 5 1 1 46416
0 46418 7 1 2 94378 46417
0 46419 5 1 1 46418
0 46420 7 1 2 46356 46419
0 46421 5 1 1 46420
0 46422 7 1 2 68238 46421
0 46423 5 1 1 46422
0 46424 7 1 2 67528 101455
0 46425 5 1 1 46424
0 46426 7 1 2 93617 46425
0 46427 5 2 1 46426
0 46428 7 1 2 74087 102340
0 46429 5 1 1 46428
0 46430 7 1 2 72796 97361
0 46431 5 1 1 46430
0 46432 7 1 2 46429 46431
0 46433 5 1 1 46432
0 46434 7 1 2 99556 46433
0 46435 5 1 1 46434
0 46436 7 1 2 80014 92178
0 46437 5 1 1 46436
0 46438 7 1 2 93638 46437
0 46439 5 2 1 46438
0 46440 7 1 2 72797 102342
0 46441 5 1 1 46440
0 46442 7 1 2 75656 92179
0 46443 5 1 1 46442
0 46444 7 1 2 46441 46443
0 46445 5 1 1 46444
0 46446 7 1 2 81055 72856
0 46447 7 1 2 46445 46446
0 46448 5 1 1 46447
0 46449 7 1 2 46435 46448
0 46450 5 1 1 46449
0 46451 7 1 2 66154 46450
0 46452 5 1 1 46451
0 46453 7 1 2 74088 95490
0 46454 5 1 1 46453
0 46455 7 1 2 90106 84755
0 46456 5 1 1 46455
0 46457 7 1 2 46454 46456
0 46458 5 1 1 46457
0 46459 7 1 2 67047 46458
0 46460 5 1 1 46459
0 46461 7 1 2 90549 100200
0 46462 5 1 1 46461
0 46463 7 1 2 46460 46462
0 46464 5 1 1 46463
0 46465 7 1 2 99260 46464
0 46466 5 1 1 46465
0 46467 7 1 2 46452 46466
0 46468 5 1 1 46467
0 46469 7 1 2 69139 46468
0 46470 5 1 1 46469
0 46471 7 1 2 78661 101817
0 46472 5 1 1 46471
0 46473 7 1 2 65528 15913
0 46474 5 1 1 46473
0 46475 7 1 2 68477 84693
0 46476 7 1 2 46474 46475
0 46477 5 1 1 46476
0 46478 7 1 2 46472 46477
0 46479 5 1 1 46478
0 46480 7 1 2 70755 46479
0 46481 5 1 1 46480
0 46482 7 1 2 72493 94438
0 46483 5 2 1 46482
0 46484 7 1 2 84756 102344
0 46485 5 1 1 46484
0 46486 7 1 2 46481 46485
0 46487 5 1 1 46486
0 46488 7 1 2 96973 100638
0 46489 7 1 2 46487 46488
0 46490 5 1 1 46489
0 46491 7 1 2 46470 46490
0 46492 5 1 1 46491
0 46493 7 1 2 83154 46492
0 46494 5 1 1 46493
0 46495 7 1 2 5514 101759
0 46496 5 1 1 46495
0 46497 7 1 2 62204 46496
0 46498 5 1 1 46497
0 46499 7 1 2 67048 75458
0 46500 7 1 2 71760 46499
0 46501 5 1 1 46500
0 46502 7 1 2 46498 46501
0 46503 5 1 1 46502
0 46504 7 1 2 99420 46503
0 46505 5 1 1 46504
0 46506 7 1 2 96649 99288
0 46507 5 1 1 46506
0 46508 7 1 2 75166 76511
0 46509 5 1 1 46508
0 46510 7 1 2 46507 46509
0 46511 5 1 1 46510
0 46512 7 1 2 93513 46511
0 46513 5 1 1 46512
0 46514 7 1 2 46505 46513
0 46515 5 1 1 46514
0 46516 7 1 2 69140 46515
0 46517 5 1 1 46516
0 46518 7 1 2 99872 99432
0 46519 7 1 2 76506 46518
0 46520 5 1 1 46519
0 46521 7 1 2 46517 46520
0 46522 5 1 1 46521
0 46523 7 1 2 70141 46522
0 46524 5 1 1 46523
0 46525 7 1 2 66155 102343
0 46526 5 1 1 46525
0 46527 7 1 2 92961 93627
0 46528 5 1 1 46527
0 46529 7 1 2 46526 46528
0 46530 5 1 1 46529
0 46531 7 1 2 72798 46530
0 46532 5 1 1 46531
0 46533 7 1 2 75657 93514
0 46534 5 1 1 46533
0 46535 7 1 2 46532 46534
0 46536 5 1 1 46535
0 46537 7 1 2 96246 97790
0 46538 7 1 2 46536 46537
0 46539 5 1 1 46538
0 46540 7 1 2 46524 46539
0 46541 5 1 1 46540
0 46542 7 1 2 82750 46541
0 46543 5 1 1 46542
0 46544 7 1 2 46494 46543
0 46545 5 1 1 46544
0 46546 7 1 2 73036 46545
0 46547 5 1 1 46546
0 46548 7 1 2 79593 96344
0 46549 5 1 1 46548
0 46550 7 1 2 70142 102339
0 46551 5 1 1 46550
0 46552 7 1 2 46549 46551
0 46553 5 1 1 46552
0 46554 7 1 2 63851 46553
0 46555 5 1 1 46554
0 46556 7 1 2 87154 91097
0 46557 5 1 1 46556
0 46558 7 1 2 72923 95477
0 46559 5 1 1 46558
0 46560 7 1 2 46557 46559
0 46561 5 1 1 46560
0 46562 7 1 2 70143 46561
0 46563 5 1 1 46562
0 46564 7 1 2 46555 46563
0 46565 5 1 1 46564
0 46566 7 1 2 67049 46565
0 46567 5 1 1 46566
0 46568 7 1 2 75122 46567
0 46569 5 1 1 46568
0 46570 7 1 2 87155 91438
0 46571 5 1 1 46570
0 46572 7 1 2 68721 12784
0 46573 5 1 1 46572
0 46574 7 1 2 92516 46573
0 46575 5 1 1 46574
0 46576 7 1 2 74383 46575
0 46577 7 1 2 46571 46576
0 46578 5 1 1 46577
0 46579 7 1 2 65848 78738
0 46580 7 1 2 46578 46579
0 46581 7 1 2 46569 46580
0 46582 5 1 1 46581
0 46583 7 1 2 77335 75922
0 46584 7 1 2 86007 46583
0 46585 7 1 2 95159 46584
0 46586 5 1 1 46585
0 46587 7 1 2 91439 93429
0 46588 7 1 2 95351 46587
0 46589 5 1 1 46588
0 46590 7 1 2 46586 46589
0 46591 7 1 2 46582 46590
0 46592 5 1 1 46591
0 46593 7 1 2 98567 46592
0 46594 5 1 1 46593
0 46595 7 1 2 75437 596
0 46596 5 1 1 46595
0 46597 7 1 2 70144 74089
0 46598 7 1 2 46596 46597
0 46599 5 1 1 46598
0 46600 7 1 2 65213 95758
0 46601 5 1 1 46600
0 46602 7 1 2 9064 46601
0 46603 7 1 2 46599 46602
0 46604 5 1 1 46603
0 46605 7 1 2 65529 46604
0 46606 5 1 1 46605
0 46607 7 1 2 74090 78116
0 46608 7 1 2 93456 46607
0 46609 5 1 1 46608
0 46610 7 1 2 46606 46609
0 46611 5 1 1 46610
0 46612 7 1 2 67050 46611
0 46613 5 1 1 46612
0 46614 7 1 2 75969 81065
0 46615 5 1 1 46614
0 46616 7 1 2 46613 46615
0 46617 5 1 1 46616
0 46618 7 1 2 87841 96974
0 46619 7 1 2 46617 46618
0 46620 5 1 1 46619
0 46621 7 1 2 46594 46620
0 46622 5 1 1 46621
0 46623 7 1 2 83155 46622
0 46624 5 1 1 46623
0 46625 7 1 2 46547 46624
0 46626 7 1 2 46423 46625
0 46627 5 1 1 46626
0 46628 7 1 2 102324 46627
0 46629 5 1 1 46628
0 46630 7 1 2 96650 99448
0 46631 5 1 1 46630
0 46632 7 1 2 76507 98064
0 46633 5 1 1 46632
0 46634 7 2 2 91347 100498
0 46635 5 1 1 102346
0 46636 7 1 2 46633 46635
0 46637 5 1 1 46636
0 46638 7 1 2 67051 46637
0 46639 5 1 1 46638
0 46640 7 1 2 46631 46639
0 46641 5 1 1 46640
0 46642 7 1 2 70145 46641
0 46643 5 1 1 46642
0 46644 7 1 2 98043 98712
0 46645 7 1 2 99190 46644
0 46646 5 1 1 46645
0 46647 7 1 2 97690 46646
0 46648 5 1 1 46647
0 46649 7 1 2 76527 46648
0 46650 5 1 1 46649
0 46651 7 2 2 86890 93293
0 46652 5 1 1 102348
0 46653 7 1 2 102349 98018
0 46654 5 1 1 46653
0 46655 7 1 2 46650 46654
0 46656 5 1 1 46655
0 46657 7 1 2 77038 46656
0 46658 5 1 1 46657
0 46659 7 1 2 46643 46658
0 46660 5 1 1 46659
0 46661 7 1 2 87791 46660
0 46662 5 1 1 46661
0 46663 7 2 2 62637 79035
0 46664 5 1 1 102350
0 46665 7 1 2 67052 102351
0 46666 5 1 1 46665
0 46667 7 1 2 71756 79515
0 46668 7 1 2 80578 46667
0 46669 5 1 1 46668
0 46670 7 1 2 46666 46669
0 46671 5 1 1 46670
0 46672 7 1 2 98019 46671
0 46673 5 1 1 46672
0 46674 7 3 2 91348 102230
0 46675 7 1 2 83743 87959
0 46676 5 1 1 46675
0 46677 7 1 2 102352 46676
0 46678 5 1 1 46677
0 46679 7 1 2 46673 46678
0 46680 5 1 1 46679
0 46681 7 1 2 72799 46680
0 46682 5 1 1 46681
0 46683 7 1 2 94578 98020
0 46684 5 1 1 46683
0 46685 7 1 2 102231 97371
0 46686 7 1 2 99162 46685
0 46687 5 1 1 46686
0 46688 7 1 2 46684 46687
0 46689 5 1 1 46688
0 46690 7 1 2 70442 46689
0 46691 5 1 1 46690
0 46692 7 1 2 46682 46691
0 46693 5 1 1 46692
0 46694 7 1 2 87733 46693
0 46695 5 1 1 46694
0 46696 7 1 2 46662 46695
0 46697 5 1 1 46696
0 46698 7 1 2 62452 46697
0 46699 5 1 1 46698
0 46700 7 1 2 76948 84922
0 46701 5 1 1 46700
0 46702 7 1 2 13842 46701
0 46703 5 1 1 46702
0 46704 7 1 2 87734 46703
0 46705 5 1 1 46704
0 46706 7 1 2 66156 100639
0 46707 7 1 2 76512 46706
0 46708 5 1 1 46707
0 46709 7 1 2 46705 46708
0 46710 5 1 1 46709
0 46711 7 1 2 67312 46710
0 46712 5 1 1 46711
0 46713 7 2 2 61318 70146
0 46714 7 1 2 64390 102355
0 46715 7 1 2 101192 46714
0 46716 5 1 1 46715
0 46717 7 1 2 46712 46716
0 46718 5 1 1 46717
0 46719 7 1 2 62205 46718
0 46720 5 1 1 46719
0 46721 7 1 2 73779 87963
0 46722 5 2 1 46721
0 46723 7 1 2 76508 87792
0 46724 5 1 1 46723
0 46725 7 1 2 102357 46724
0 46726 5 1 1 46725
0 46727 7 1 2 72857 79581
0 46728 7 1 2 46726 46727
0 46729 5 1 1 46728
0 46730 7 1 2 46720 46729
0 46731 5 1 1 46730
0 46732 7 1 2 98021 46731
0 46733 5 1 1 46732
0 46734 7 1 2 46699 46733
0 46735 5 1 1 46734
0 46736 7 1 2 63852 46735
0 46737 5 1 1 46736
0 46738 7 1 2 76923 84831
0 46739 5 1 1 46738
0 46740 7 1 2 97679 46739
0 46741 5 1 1 46740
0 46742 7 2 2 91869 93031
0 46743 7 4 2 69141 65214
0 46744 7 1 2 86561 102361
0 46745 7 1 2 102359 46744
0 46746 5 1 1 46745
0 46747 7 1 2 46741 46746
0 46748 5 1 1 46747
0 46749 7 1 2 62206 46748
0 46750 5 1 1 46749
0 46751 7 1 2 99198 100182
0 46752 5 1 1 46751
0 46753 7 1 2 46750 46752
0 46754 5 1 1 46753
0 46755 7 1 2 76528 46754
0 46756 5 1 1 46755
0 46757 7 2 2 102232 101500
0 46758 5 1 1 102365
0 46759 7 1 2 80579 95321
0 46760 7 1 2 102360 46759
0 46761 5 1 1 46760
0 46762 7 1 2 46758 46761
0 46763 5 1 1 46762
0 46764 7 1 2 83731 84923
0 46765 7 1 2 46763 46764
0 46766 5 1 1 46765
0 46767 7 1 2 46756 46766
0 46768 5 1 1 46767
0 46769 7 1 2 87793 46768
0 46770 5 1 1 46769
0 46771 7 1 2 77383 94588
0 46772 5 1 1 46771
0 46773 7 2 2 64183 80580
0 46774 7 1 2 86008 85259
0 46775 7 1 2 102367 46774
0 46776 5 1 1 46775
0 46777 7 1 2 46772 46776
0 46778 5 1 1 46777
0 46779 7 1 2 98022 46778
0 46780 5 1 1 46779
0 46781 7 1 2 92331 102366
0 46782 5 1 1 46781
0 46783 7 1 2 46780 46782
0 46784 5 1 1 46783
0 46785 7 1 2 70443 46784
0 46786 5 1 1 46785
0 46787 7 1 2 80757 102347
0 46788 5 1 1 46787
0 46789 7 1 2 68722 91149
0 46790 7 1 2 98023 46789
0 46791 5 1 1 46790
0 46792 7 1 2 46788 46791
0 46793 5 1 1 46792
0 46794 7 1 2 64184 78018
0 46795 7 1 2 46793 46794
0 46796 5 1 1 46795
0 46797 7 1 2 46786 46796
0 46798 5 1 1 46797
0 46799 7 1 2 87735 46798
0 46800 5 1 1 46799
0 46801 7 1 2 46770 46800
0 46802 7 1 2 46737 46801
0 46803 5 1 1 46802
0 46804 7 1 2 63637 46803
0 46805 5 1 1 46804
0 46806 7 4 2 61319 93628
0 46807 5 1 1 102369
0 46808 7 1 2 92294 102370
0 46809 5 1 1 46808
0 46810 7 1 2 74144 87878
0 46811 5 1 1 46810
0 46812 7 1 2 46809 46811
0 46813 5 1 1 46812
0 46814 7 1 2 70147 46813
0 46815 5 1 1 46814
0 46816 7 1 2 96316 102371
0 46817 5 1 1 46816
0 46818 7 1 2 46815 46817
0 46819 5 1 1 46818
0 46820 7 2 2 93576 97463
0 46821 7 1 2 97791 102373
0 46822 7 1 2 46819 46821
0 46823 5 1 1 46822
0 46824 7 1 2 65215 101389
0 46825 5 1 1 46824
0 46826 7 4 2 66292 91870
0 46827 7 1 2 78200 94760
0 46828 7 1 2 102375 46827
0 46829 5 1 1 46828
0 46830 7 1 2 46825 46829
0 46831 5 1 1 46830
0 46832 7 1 2 71872 87736
0 46833 7 1 2 46831 46832
0 46834 5 1 1 46833
0 46835 7 1 2 92839 97995
0 46836 7 1 2 73037 46835
0 46837 7 1 2 88450 93579
0 46838 7 1 2 46836 46837
0 46839 5 1 1 46838
0 46840 7 1 2 46834 46839
0 46841 5 1 1 46840
0 46842 7 1 2 71354 46841
0 46843 5 1 1 46842
0 46844 7 1 2 82971 93635
0 46845 7 2 2 62638 90620
0 46846 7 1 2 99297 102379
0 46847 7 1 2 46844 46846
0 46848 5 1 1 46847
0 46849 7 1 2 46843 46848
0 46850 7 1 2 46823 46849
0 46851 5 1 1 46850
0 46852 7 1 2 72800 46851
0 46853 5 1 1 46852
0 46854 7 4 2 98197 99623
0 46855 7 1 2 79017 102381
0 46856 5 1 1 46855
0 46857 7 1 2 88357 94761
0 46858 7 1 2 93743 46857
0 46859 5 1 1 46858
0 46860 7 1 2 46856 46859
0 46861 5 1 1 46860
0 46862 7 1 2 86551 46861
0 46863 5 1 1 46862
0 46864 7 1 2 46853 46863
0 46865 5 1 1 46864
0 46866 7 1 2 62207 46865
0 46867 5 1 1 46866
0 46868 7 1 2 74384 99155
0 46869 7 1 2 76509 46868
0 46870 5 1 1 46869
0 46871 7 2 2 88032 99694
0 46872 5 1 1 102385
0 46873 7 1 2 87794 96651
0 46874 5 1 1 46873
0 46875 7 1 2 46872 46874
0 46876 5 1 1 46875
0 46877 7 1 2 99257 99775
0 46878 7 1 2 46876 46877
0 46879 5 1 1 46878
0 46880 7 1 2 46870 46879
0 46881 5 1 1 46880
0 46882 7 1 2 76986 46881
0 46883 5 1 1 46882
0 46884 7 3 2 80680 94379
0 46885 7 3 2 90880 99582
0 46886 7 1 2 73967 91375
0 46887 7 1 2 96257 46886
0 46888 7 1 2 102390 46887
0 46889 7 1 2 102387 46888
0 46890 5 1 1 46889
0 46891 7 1 2 46883 46890
0 46892 7 1 2 46867 46891
0 46893 7 1 2 46805 46892
0 46894 5 1 1 46893
0 46895 7 1 2 63398 46894
0 46896 5 1 1 46895
0 46897 7 1 2 86661 94566
0 46898 5 1 1 46897
0 46899 7 1 2 63638 102328
0 46900 5 1 1 46899
0 46901 7 1 2 46898 46900
0 46902 5 1 1 46901
0 46903 7 1 2 70756 46902
0 46904 5 1 1 46903
0 46905 7 1 2 78095 77753
0 46906 5 1 1 46905
0 46907 7 1 2 46904 46906
0 46908 5 1 1 46907
0 46909 7 1 2 63853 46908
0 46910 5 1 1 46909
0 46911 7 1 2 68723 75099
0 46912 7 1 2 80681 46911
0 46913 5 1 1 46912
0 46914 7 1 2 46910 46913
0 46915 5 1 1 46914
0 46916 7 1 2 62453 46915
0 46917 5 1 1 46916
0 46918 7 1 2 91683 93942
0 46919 5 1 1 46918
0 46920 7 1 2 75861 92744
0 46921 5 1 1 46920
0 46922 7 1 2 46919 46921
0 46923 5 1 1 46922
0 46924 7 1 2 78084 46923
0 46925 5 1 1 46924
0 46926 7 1 2 75204 101485
0 46927 5 1 1 46926
0 46928 7 2 2 73038 71744
0 46929 5 1 1 102393
0 46930 7 1 2 77854 89940
0 46931 5 1 1 46930
0 46932 7 1 2 46929 46931
0 46933 7 1 2 46927 46932
0 46934 5 1 1 46933
0 46935 7 1 2 62208 46934
0 46936 5 1 1 46935
0 46937 7 1 2 97835 46936
0 46938 5 1 1 46937
0 46939 7 1 2 94945 46938
0 46940 5 1 1 46939
0 46941 7 1 2 46925 46940
0 46942 7 1 2 46917 46941
0 46943 5 1 1 46942
0 46944 7 1 2 98887 46943
0 46945 5 1 1 46944
0 46946 7 1 2 62209 88419
0 46947 5 1 1 46946
0 46948 7 1 2 89320 91150
0 46949 5 1 1 46948
0 46950 7 1 2 46947 46949
0 46951 5 1 1 46950
0 46952 7 1 2 63639 46951
0 46953 5 1 1 46952
0 46954 7 1 2 77056 80015
0 46955 5 1 1 46954
0 46956 7 1 2 46953 46955
0 46957 5 1 1 46956
0 46958 7 1 2 97740 46957
0 46959 5 1 1 46958
0 46960 7 1 2 46945 46959
0 46961 5 1 1 46960
0 46962 7 1 2 72801 46961
0 46963 5 1 1 46962
0 46964 7 1 2 74091 93342
0 46965 5 1 1 46964
0 46966 7 1 2 94291 46965
0 46967 5 2 1 46966
0 46968 7 1 2 98937 102395
0 46969 5 1 1 46968
0 46970 7 1 2 67313 99952
0 46971 5 1 1 46970
0 46972 7 1 2 46969 46971
0 46973 5 1 1 46972
0 46974 7 1 2 76904 46973
0 46975 5 1 1 46974
0 46976 7 3 2 87842 97719
0 46977 5 1 1 102397
0 46978 7 2 2 65216 95132
0 46979 5 1 1 102400
0 46980 7 3 2 77676 46979
0 46981 5 1 1 102402
0 46982 7 1 2 102403 46324
0 46983 5 1 1 46982
0 46984 7 1 2 102398 46983
0 46985 5 1 1 46984
0 46986 7 1 2 66157 74092
0 46987 7 1 2 80581 46986
0 46988 7 1 2 98585 46987
0 46989 5 1 1 46988
0 46990 7 1 2 46985 46989
0 46991 5 1 1 46990
0 46992 7 1 2 62454 46991
0 46993 5 1 1 46992
0 46994 7 1 2 46975 46993
0 46995 5 1 1 46994
0 46996 7 1 2 63854 46995
0 46997 5 1 1 46996
0 46998 7 4 2 99282 99906
0 46999 7 1 2 79036 102405
0 47000 5 1 1 46999
0 47001 7 1 2 79876 102399
0 47002 5 1 1 47001
0 47003 7 2 2 66158 77155
0 47004 7 1 2 74093 94380
0 47005 7 1 2 102409 47004
0 47006 5 1 1 47005
0 47007 7 1 2 47002 47006
0 47008 5 1 1 47007
0 47009 7 1 2 75970 47008
0 47010 5 1 1 47009
0 47011 7 1 2 93951 98888
0 47012 7 1 2 94585 47011
0 47013 5 1 1 47012
0 47014 7 1 2 47010 47013
0 47015 5 1 1 47014
0 47016 7 1 2 84949 47015
0 47017 5 1 1 47016
0 47018 7 1 2 47000 47017
0 47019 7 1 2 46997 47018
0 47020 5 1 1 47019
0 47021 7 1 2 63640 47020
0 47022 5 1 1 47021
0 47023 7 2 2 76987 73222
0 47024 5 1 1 102411
0 47025 7 1 2 102406 102412
0 47026 5 1 1 47025
0 47027 7 1 2 47022 47026
0 47028 7 1 2 46963 47027
0 47029 5 1 1 47028
0 47030 7 1 2 63399 47029
0 47031 5 1 1 47030
0 47032 7 1 2 95283 99919
0 47033 7 2 2 94156 47032
0 47034 7 1 2 73718 85193
0 47035 7 1 2 102410 47034
0 47036 7 1 2 102413 47035
0 47037 5 1 1 47036
0 47038 7 1 2 47031 47037
0 47039 5 1 1 47038
0 47040 7 1 2 90722 47039
0 47041 5 1 1 47040
0 47042 7 1 2 77162 84721
0 47043 7 1 2 92984 102388
0 47044 7 1 2 47042 47043
0 47045 5 1 1 47044
0 47046 7 1 2 47041 47045
0 47047 7 1 2 46896 47046
0 47048 5 1 1 47047
0 47049 7 1 2 61911 47048
0 47050 5 1 1 47049
0 47051 7 1 2 88227 93377
0 47052 7 2 2 62893 91871
0 47053 7 1 2 102415 98486
0 47054 7 1 2 47051 47053
0 47055 7 1 2 102389 47054
0 47056 5 1 1 47055
0 47057 7 1 2 66159 90470
0 47058 7 1 2 100971 47057
0 47059 7 1 2 90723 102414
0 47060 7 1 2 47058 47059
0 47061 5 1 1 47060
0 47062 7 1 2 47056 47061
0 47063 7 1 2 47050 47062
0 47064 5 1 1 47063
0 47065 7 1 2 63201 47064
0 47066 5 1 1 47065
0 47067 7 1 2 46629 47066
0 47068 5 1 1 47067
0 47069 7 1 2 64984 47068
0 47070 5 1 1 47069
0 47071 7 1 2 79047 84832
0 47072 5 2 1 47071
0 47073 7 1 2 101825 102417
0 47074 5 1 1 47073
0 47075 7 1 2 64391 77855
0 47076 7 1 2 79006 47075
0 47077 7 1 2 102380 47076
0 47078 5 1 1 47077
0 47079 7 1 2 47074 47078
0 47080 5 1 1 47079
0 47081 7 1 2 75838 47080
0 47082 5 1 1 47081
0 47083 7 1 2 85269 74293
0 47084 5 1 1 47083
0 47085 7 1 2 76806 79782
0 47086 5 1 1 47085
0 47087 7 1 2 47084 47086
0 47088 5 1 1 47087
0 47089 7 1 2 71544 47088
0 47090 5 1 1 47089
0 47091 7 1 2 62639 74667
0 47092 7 1 2 92737 47091
0 47093 5 1 1 47092
0 47094 7 1 2 47090 47093
0 47095 5 1 1 47094
0 47096 7 1 2 62210 47095
0 47097 5 1 1 47096
0 47098 7 2 2 65849 76807
0 47099 7 1 2 90464 102419
0 47100 5 1 1 47099
0 47101 7 1 2 47097 47100
0 47102 5 1 1 47101
0 47103 7 1 2 65217 47102
0 47104 5 1 1 47103
0 47105 7 2 2 71786 78797
0 47106 7 1 2 76905 101177
0 47107 7 1 2 102421 47106
0 47108 5 1 1 47107
0 47109 7 1 2 47104 47108
0 47110 5 1 1 47109
0 47111 7 1 2 92633 47110
0 47112 5 1 1 47111
0 47113 7 1 2 47082 47112
0 47114 5 1 1 47113
0 47115 7 1 2 63400 47114
0 47116 5 1 1 47115
0 47117 7 2 2 67898 97775
0 47118 7 1 2 81602 102423
0 47119 7 1 2 97197 47118
0 47120 7 1 2 102418 47119
0 47121 5 1 1 47120
0 47122 7 1 2 47116 47121
0 47123 5 1 1 47122
0 47124 7 1 2 63202 47123
0 47125 5 1 1 47124
0 47126 7 2 2 73039 92711
0 47127 7 1 2 102425 99460
0 47128 5 1 1 47127
0 47129 7 1 2 84199 91588
0 47130 5 1 1 47129
0 47131 7 1 2 98607 47130
0 47132 5 1 1 47131
0 47133 7 1 2 90621 97423
0 47134 7 1 2 47132 47133
0 47135 5 1 1 47134
0 47136 7 1 2 47128 47135
0 47137 5 1 1 47136
0 47138 7 1 2 61912 47137
0 47139 5 1 1 47138
0 47140 7 1 2 76237 87097
0 47141 7 1 2 92634 47140
0 47142 7 1 2 74595 47141
0 47143 5 1 1 47142
0 47144 7 1 2 47139 47143
0 47145 5 1 1 47144
0 47146 7 1 2 63203 47145
0 47147 5 1 1 47146
0 47148 7 1 2 67053 74421
0 47149 5 1 1 47148
0 47150 7 1 2 18637 47149
0 47151 5 1 1 47150
0 47152 7 1 2 90491 87843
0 47153 7 1 2 93818 47152
0 47154 7 1 2 47151 47153
0 47155 5 1 1 47154
0 47156 7 1 2 47147 47155
0 47157 5 1 1 47156
0 47158 7 1 2 65218 47157
0 47159 5 1 1 47158
0 47160 7 2 2 73079 95126
0 47161 7 1 2 82636 102427
0 47162 7 1 2 101412 47161
0 47163 5 1 1 47162
0 47164 7 1 2 47159 47163
0 47165 5 1 1 47164
0 47166 7 1 2 71355 47165
0 47167 5 1 1 47166
0 47168 7 1 2 74339 84828
0 47169 5 1 1 47168
0 47170 7 1 2 78401 95352
0 47171 5 1 1 47170
0 47172 7 1 2 47169 47171
0 47173 5 1 1 47172
0 47174 7 1 2 73040 47173
0 47175 5 1 1 47174
0 47176 7 1 2 77039 102345
0 47177 5 1 1 47176
0 47178 7 1 2 76906 94070
0 47179 5 1 1 47178
0 47180 7 1 2 47177 47179
0 47181 5 1 1 47180
0 47182 7 1 2 88514 47181
0 47183 5 1 1 47182
0 47184 7 1 2 47175 47183
0 47185 5 1 1 47184
0 47186 7 1 2 96095 99415
0 47187 7 1 2 47185 47186
0 47188 5 1 1 47187
0 47189 7 1 2 47167 47188
0 47190 7 1 2 47125 47189
0 47191 5 1 1 47190
0 47192 7 1 2 72802 47191
0 47193 5 1 1 47192
0 47194 7 2 2 73041 84689
0 47195 7 1 2 98563 102429
0 47196 5 1 1 47195
0 47197 7 1 2 90040 93819
0 47198 7 1 2 96374 47197
0 47199 5 1 1 47198
0 47200 7 1 2 47196 47199
0 47201 5 1 1 47200
0 47202 7 1 2 68478 47201
0 47203 5 1 1 47202
0 47204 7 2 2 82675 90676
0 47205 7 1 2 95693 101178
0 47206 7 1 2 102431 47205
0 47207 5 1 1 47206
0 47208 7 1 2 47203 47207
0 47209 5 1 1 47208
0 47210 7 1 2 87844 47209
0 47211 5 1 1 47210
0 47212 7 1 2 84892 85972
0 47213 5 1 1 47212
0 47214 7 1 2 71873 80525
0 47215 5 1 1 47214
0 47216 7 1 2 74850 73491
0 47217 7 1 2 47215 47216
0 47218 5 1 1 47217
0 47219 7 2 2 47213 47218
0 47220 5 1 1 102433
0 47221 7 2 2 100364 98110
0 47222 7 1 2 85175 102435
0 47223 7 1 2 47220 47222
0 47224 5 1 1 47223
0 47225 7 1 2 47211 47224
0 47226 5 1 1 47225
0 47227 7 1 2 62211 47226
0 47228 5 1 1 47227
0 47229 7 2 2 80229 98497
0 47230 7 1 2 72426 96833
0 47231 7 1 2 102437 47230
0 47232 5 1 1 47231
0 47233 7 1 2 31793 47232
0 47234 5 1 1 47233
0 47235 7 1 2 61401 47234
0 47236 5 1 1 47235
0 47237 7 1 2 78380 96681
0 47238 7 1 2 98553 47237
0 47239 5 1 1 47238
0 47240 7 1 2 47236 47239
0 47241 5 1 1 47240
0 47242 7 1 2 67529 47241
0 47243 5 1 1 47242
0 47244 7 1 2 87859 101863
0 47245 7 1 2 98548 47244
0 47246 5 1 1 47245
0 47247 7 1 2 47243 47246
0 47248 5 1 1 47247
0 47249 7 1 2 73042 47248
0 47250 5 1 1 47249
0 47251 7 1 2 92259 102436
0 47252 7 1 2 102396 47251
0 47253 5 1 1 47252
0 47254 7 1 2 47250 47253
0 47255 5 1 1 47254
0 47256 7 1 2 75100 47255
0 47257 5 1 1 47256
0 47258 7 1 2 47228 47257
0 47259 5 1 1 47258
0 47260 7 1 2 65530 47259
0 47261 5 1 1 47260
0 47262 7 1 2 92857 95038
0 47263 5 1 1 47262
0 47264 7 2 2 91832 100334
0 47265 5 1 1 102439
0 47266 7 1 2 66778 102440
0 47267 5 1 1 47266
0 47268 7 1 2 47263 47267
0 47269 5 1 1 47268
0 47270 7 1 2 66293 47269
0 47271 5 1 1 47270
0 47272 7 1 2 80953 98498
0 47273 7 1 2 101995 47272
0 47274 5 1 1 47273
0 47275 7 1 2 47271 47274
0 47276 5 1 1 47275
0 47277 7 1 2 90889 47276
0 47278 5 1 1 47277
0 47279 7 1 2 75487 90442
0 47280 7 1 2 101413 47279
0 47281 5 1 1 47280
0 47282 7 1 2 47278 47281
0 47283 5 1 1 47282
0 47284 7 1 2 99344 47283
0 47285 5 1 1 47284
0 47286 7 1 2 47261 47285
0 47287 5 1 1 47286
0 47288 7 1 2 65219 47287
0 47289 5 1 1 47288
0 47290 7 1 2 36364 47265
0 47291 5 2 1 47290
0 47292 7 1 2 66294 102441
0 47293 5 1 1 47292
0 47294 7 1 2 47293 36421
0 47295 5 1 1 47294
0 47296 7 1 2 47295 102430
0 47297 5 1 1 47296
0 47298 7 1 2 94071 101414
0 47299 5 1 1 47298
0 47300 7 1 2 47297 47299
0 47301 5 1 1 47300
0 47302 7 1 2 66779 47301
0 47303 5 1 1 47302
0 47304 7 2 2 92858 98091
0 47305 7 1 2 90443 102443
0 47306 7 1 2 102426 47305
0 47307 5 1 1 47306
0 47308 7 1 2 47303 47307
0 47309 5 1 1 47308
0 47310 7 1 2 102428 47309
0 47311 5 1 1 47310
0 47312 7 1 2 92647 47311
0 47313 7 1 2 47289 47312
0 47314 7 1 2 47193 47313
0 47315 5 1 1 47314
0 47316 7 1 2 74094 85973
0 47317 5 1 1 47316
0 47318 7 1 2 91562 47317
0 47319 5 1 1 47318
0 47320 7 1 2 75167 47319
0 47321 5 1 1 47320
0 47322 7 1 2 47321 38366
0 47323 5 1 1 47322
0 47324 7 3 2 91497 102325
0 47325 7 1 2 47323 102445
0 47326 5 1 1 47325
0 47327 7 1 2 87903 102446
0 47328 5 1 1 47327
0 47329 7 1 2 76540 102444
0 47330 5 1 1 47329
0 47331 7 1 2 47328 47330
0 47332 5 1 1 47331
0 47333 7 1 2 71356 47332
0 47334 5 1 1 47333
0 47335 7 1 2 74042 102422
0 47336 7 1 2 102326 47335
0 47337 5 1 1 47336
0 47338 7 1 2 47334 47337
0 47339 5 1 1 47338
0 47340 7 1 2 72803 47339
0 47341 5 1 1 47340
0 47342 7 1 2 75193 102447
0 47343 7 1 2 102337 47342
0 47344 5 1 1 47343
0 47345 7 1 2 47341 47344
0 47346 5 1 1 47345
0 47347 7 1 2 65850 47346
0 47348 5 1 1 47347
0 47349 7 1 2 47326 47348
0 47350 5 1 1 47349
0 47351 7 1 2 68239 47350
0 47352 5 1 1 47351
0 47353 7 1 2 77754 95770
0 47354 5 1 1 47353
0 47355 7 1 2 47354 102434
0 47356 5 1 1 47355
0 47357 7 1 2 76391 47356
0 47358 5 1 1 47357
0 47359 7 1 2 93344 97900
0 47360 5 1 1 47359
0 47361 7 1 2 47358 47360
0 47362 5 1 1 47361
0 47363 7 1 2 61913 47362
0 47364 5 1 1 47363
0 47365 7 1 2 72351 86045
0 47366 7 1 2 95233 47365
0 47367 5 1 1 47366
0 47368 7 1 2 47364 47367
0 47369 5 1 1 47368
0 47370 7 1 2 102432 47369
0 47371 5 1 1 47370
0 47372 7 1 2 47352 47371
0 47373 5 1 1 47372
0 47374 7 1 2 95304 47373
0 47375 5 1 1 47374
0 47376 7 1 2 92659 47375
0 47377 5 1 1 47376
0 47378 7 2 2 69142 69844
0 47379 7 1 2 96953 102448
0 47380 7 1 2 47377 47379
0 47381 7 1 2 47315 47380
0 47382 5 1 1 47381
0 47383 7 1 2 64574 47382
0 47384 7 1 2 47070 47383
0 47385 5 1 1 47384
0 47386 7 2 2 73043 93642
0 47387 7 1 2 99946 102450
0 47388 5 1 1 47387
0 47389 7 1 2 62212 73997
0 47390 7 1 2 91744 97424
0 47391 7 1 2 47389 47390
0 47392 5 1 1 47391
0 47393 7 1 2 47388 47392
0 47394 5 1 1 47393
0 47395 7 1 2 90677 47394
0 47396 5 1 1 47395
0 47397 7 1 2 75037 98595
0 47398 7 1 2 97401 47397
0 47399 7 1 2 98917 47398
0 47400 5 1 1 47399
0 47401 7 1 2 47396 47400
0 47402 5 1 1 47401
0 47403 7 1 2 66160 47402
0 47404 5 1 1 47403
0 47405 7 1 2 63855 99439
0 47406 7 1 2 98055 47405
0 47407 7 1 2 98918 47406
0 47408 5 1 1 47407
0 47409 7 1 2 47404 47408
0 47410 5 1 1 47409
0 47411 7 1 2 94876 47410
0 47412 5 1 1 47411
0 47413 7 1 2 99949 102451
0 47414 5 1 1 47413
0 47415 7 2 2 79963 98843
0 47416 7 1 2 102452 98639
0 47417 5 1 1 47416
0 47418 7 1 2 47414 47417
0 47419 5 1 1 47418
0 47420 7 1 2 90678 47419
0 47421 5 1 1 47420
0 47422 7 2 2 79964 90644
0 47423 7 2 2 87649 98919
0 47424 7 1 2 102454 102456
0 47425 5 1 1 47424
0 47426 7 1 2 47421 47425
0 47427 5 1 1 47426
0 47428 7 1 2 66161 47427
0 47429 5 1 1 47428
0 47430 7 2 2 98075 99440
0 47431 7 1 2 102457 102458
0 47432 5 1 1 47431
0 47433 7 1 2 47429 47432
0 47434 5 1 1 47433
0 47435 7 1 2 94946 47434
0 47436 5 1 1 47435
0 47437 7 1 2 47412 47436
0 47438 5 1 1 47437
0 47439 7 1 2 64985 47438
0 47440 5 1 1 47439
0 47441 7 1 2 79483 102329
0 47442 5 1 1 47441
0 47443 7 1 2 67054 77617
0 47444 7 1 2 90107 47443
0 47445 5 1 1 47444
0 47446 7 1 2 47442 47445
0 47447 5 1 1 47446
0 47448 7 1 2 68724 47447
0 47449 5 1 1 47448
0 47450 7 1 2 72945 80665
0 47451 5 1 1 47450
0 47452 7 1 2 47449 47451
0 47453 5 1 1 47452
0 47454 7 1 2 68479 47453
0 47455 5 1 1 47454
0 47456 7 1 2 75101 80775
0 47457 7 1 2 102420 47456
0 47458 5 1 1 47457
0 47459 7 1 2 47455 47458
0 47460 5 2 1 47459
0 47461 7 1 2 62640 102460
0 47462 5 1 1 47461
0 47463 7 1 2 82976 77359
0 47464 7 1 2 90330 47463
0 47465 5 1 1 47464
0 47466 7 1 2 47462 47465
0 47467 5 1 1 47466
0 47468 7 1 2 92180 47467
0 47469 5 1 1 47468
0 47470 7 1 2 81017 100144
0 47471 7 1 2 102453 47470
0 47472 5 2 1 47471
0 47473 7 1 2 47469 102462
0 47474 5 1 1 47473
0 47475 7 1 2 90679 47474
0 47476 5 1 1 47475
0 47477 7 1 2 63641 98844
0 47478 7 2 2 81018 47477
0 47479 7 1 2 102455 102464
0 47480 5 2 1 47479
0 47481 7 1 2 47476 102466
0 47482 5 1 1 47481
0 47483 7 1 2 66162 47482
0 47484 5 1 1 47483
0 47485 7 1 2 102459 102465
0 47486 5 2 1 47485
0 47487 7 1 2 47484 102468
0 47488 5 1 1 47487
0 47489 7 1 2 88951 47488
0 47490 5 1 1 47489
0 47491 7 1 2 47440 47490
0 47492 5 1 1 47491
0 47493 7 1 2 66780 47492
0 47494 5 1 1 47493
0 47495 7 1 2 93643 102461
0 47496 5 1 1 47495
0 47497 7 1 2 102463 47496
0 47498 5 1 1 47497
0 47499 7 1 2 90680 47498
0 47500 5 1 1 47499
0 47501 7 1 2 102467 47500
0 47502 5 1 1 47501
0 47503 7 1 2 66163 47502
0 47504 5 1 1 47503
0 47505 7 1 2 102469 47504
0 47506 5 1 1 47505
0 47507 7 1 2 92009 47506
0 47508 5 1 1 47507
0 47509 7 1 2 47494 47508
0 47510 5 1 1 47509
0 47511 7 1 2 68042 47510
0 47512 5 1 1 47511
0 47513 7 1 2 66164 84866
0 47514 7 1 2 92827 97425
0 47515 7 1 2 47513 47514
0 47516 7 1 2 93820 101677
0 47517 7 1 2 47515 47516
0 47518 7 1 2 90454 47517
0 47519 5 1 1 47518
0 47520 7 1 2 47512 47519
0 47521 5 1 1 47520
0 47522 7 1 2 69143 47521
0 47523 5 1 1 47522
0 47524 7 1 2 102267 98799
0 47525 5 1 1 47524
0 47526 7 3 2 63988 97741
0 47527 7 1 2 71068 90228
0 47528 7 1 2 102470 47527
0 47529 5 1 1 47528
0 47530 7 1 2 47525 47529
0 47531 5 1 1 47530
0 47532 7 1 2 90724 47531
0 47533 5 1 1 47532
0 47534 7 2 2 63989 77336
0 47535 5 1 1 102473
0 47536 7 1 2 102474 99534
0 47537 7 3 2 64296 64986
0 47538 7 4 2 69249 102475
0 47539 7 1 2 102478 98875
0 47540 7 1 2 47536 47539
0 47541 5 1 1 47540
0 47542 7 1 2 65851 80582
0 47543 7 1 2 100233 98024
0 47544 7 1 2 47542 47543
0 47545 7 1 2 93021 99535
0 47546 5 2 1 47545
0 47547 7 1 2 87764 102482
0 47548 5 2 1 47547
0 47549 7 1 2 66781 77049
0 47550 7 1 2 102483 47549
0 47551 5 1 1 47550
0 47552 7 1 2 102484 47551
0 47553 7 1 2 47544 47552
0 47554 5 1 1 47553
0 47555 7 1 2 47541 47554
0 47556 7 1 2 47533 47555
0 47557 5 1 1 47556
0 47558 7 1 2 89653 47557
0 47559 5 1 1 47558
0 47560 7 2 2 90481 99048
0 47561 7 1 2 76827 83682
0 47562 7 1 2 95043 47561
0 47563 7 1 2 99995 47562
0 47564 7 1 2 102486 47563
0 47565 5 1 1 47564
0 47566 7 1 2 47559 47565
0 47567 5 1 1 47566
0 47568 7 1 2 74553 47567
0 47569 5 1 1 47568
0 47570 7 1 2 74145 94012
0 47571 7 1 2 100853 47570
0 47572 5 1 1 47571
0 47573 7 1 2 98596 98219
0 47574 7 1 2 99773 47573
0 47575 5 1 1 47574
0 47576 7 1 2 47572 47575
0 47577 5 1 1 47576
0 47578 7 1 2 83156 47577
0 47579 5 1 1 47578
0 47580 7 2 2 70757 101264
0 47581 7 1 2 88562 94787
0 47582 7 1 2 90413 47581
0 47583 7 1 2 102488 47582
0 47584 5 1 1 47583
0 47585 7 1 2 47579 47584
0 47586 5 1 1 47585
0 47587 7 1 2 65220 47586
0 47588 5 1 1 47587
0 47589 7 1 2 83069 79582
0 47590 7 1 2 93022 47589
0 47591 7 1 2 94145 47590
0 47592 7 1 2 91031 47591
0 47593 5 1 1 47592
0 47594 7 1 2 47588 47593
0 47595 5 1 1 47594
0 47596 7 1 2 68480 47595
0 47597 5 1 1 47596
0 47598 7 1 2 78085 70997
0 47599 7 1 2 96834 47598
0 47600 7 1 2 80359 47599
0 47601 7 1 2 91032 47600
0 47602 5 1 1 47601
0 47603 7 1 2 47597 47602
0 47604 5 1 1 47603
0 47605 7 1 2 68043 47604
0 47606 5 1 1 47605
0 47607 7 1 2 68875 72946
0 47608 7 1 2 86280 47607
0 47609 5 1 1 47608
0 47610 7 1 2 47024 47609
0 47611 5 1 1 47610
0 47612 7 1 2 82383 93700
0 47613 7 1 2 102487 47612
0 47614 7 1 2 47611 47613
0 47615 5 1 1 47614
0 47616 7 1 2 47606 47615
0 47617 5 1 1 47616
0 47618 7 1 2 102476 47617
0 47619 5 1 1 47618
0 47620 7 1 2 47569 47619
0 47621 7 1 2 47523 47620
0 47622 5 1 1 47621
0 47623 7 1 2 71176 47622
0 47624 5 1 1 47623
0 47625 7 2 2 68240 98477
0 47626 7 1 2 65531 97063
0 47627 5 1 1 47626
0 47628 7 1 2 91417 94002
0 47629 5 1 1 47628
0 47630 7 1 2 47627 47629
0 47631 5 1 1 47630
0 47632 7 1 2 67530 47631
0 47633 5 1 1 47632
0 47634 7 1 2 72377 97061
0 47635 5 1 1 47634
0 47636 7 1 2 47633 47635
0 47637 5 1 1 47636
0 47638 7 1 2 64185 47637
0 47639 5 1 1 47638
0 47640 7 1 2 76719 86011
0 47641 5 1 1 47640
0 47642 7 1 2 47639 47641
0 47643 5 2 1 47642
0 47644 7 1 2 78086 102492
0 47645 5 1 1 47644
0 47646 7 1 2 87150 102394
0 47647 5 1 1 47646
0 47648 7 1 2 75292 87974
0 47649 7 1 2 84705 47648
0 47650 5 1 1 47649
0 47651 7 1 2 47647 47650
0 47652 5 2 1 47651
0 47653 7 1 2 94947 102494
0 47654 5 1 1 47653
0 47655 7 1 2 47645 47654
0 47656 5 1 1 47655
0 47657 7 1 2 98568 47656
0 47658 5 1 1 47657
0 47659 7 1 2 65221 2767
0 47660 5 1 1 47659
0 47661 7 1 2 70148 99466
0 47662 5 1 1 47661
0 47663 7 2 2 47660 47662
0 47664 5 1 1 102496
0 47665 7 1 2 62641 102497
0 47666 5 1 1 47665
0 47667 7 1 2 88420 98642
0 47668 5 1 1 47667
0 47669 7 1 2 47666 47668
0 47670 5 1 1 47669
0 47671 7 1 2 95292 101001
0 47672 7 1 2 47670 47671
0 47673 5 1 1 47672
0 47674 7 1 2 47658 47673
0 47675 5 1 1 47674
0 47676 7 1 2 64987 47675
0 47677 5 1 1 47676
0 47678 7 1 2 86294 101356
0 47679 5 1 1 47678
0 47680 7 1 2 62894 47679
0 47681 5 1 1 47680
0 47682 7 1 2 62455 85601
0 47683 5 1 1 47682
0 47684 7 1 2 64186 91654
0 47685 7 1 2 47683 47684
0 47686 5 1 1 47685
0 47687 7 1 2 47681 47686
0 47688 5 1 1 47687
0 47689 7 1 2 68725 47688
0 47690 5 1 1 47689
0 47691 7 1 2 73492 87509
0 47692 5 1 1 47691
0 47693 7 1 2 87910 47692
0 47694 5 2 1 47693
0 47695 7 1 2 80477 102498
0 47696 5 1 1 47695
0 47697 7 1 2 47690 47696
0 47698 5 1 1 47697
0 47699 7 1 2 65532 47698
0 47700 5 1 1 47699
0 47701 7 1 2 67531 77873
0 47702 5 1 1 47701
0 47703 7 1 2 67740 77777
0 47704 7 1 2 85780 47703
0 47705 5 1 1 47704
0 47706 7 1 2 47702 47705
0 47707 5 1 1 47706
0 47708 7 1 2 67314 47707
0 47709 5 1 1 47708
0 47710 7 1 2 77874 82889
0 47711 5 1 1 47710
0 47712 7 1 2 47709 47711
0 47713 5 1 1 47712
0 47714 7 1 2 77951 47713
0 47715 5 1 1 47714
0 47716 7 1 2 47700 47715
0 47717 5 1 1 47716
0 47718 7 1 2 78614 93877
0 47719 7 1 2 99302 47718
0 47720 7 1 2 47717 47719
0 47721 5 1 1 47720
0 47722 7 1 2 47677 47721
0 47723 5 1 1 47722
0 47724 7 1 2 62213 47723
0 47725 5 1 1 47724
0 47726 7 2 2 102305 99421
0 47727 7 1 2 87621 102495
0 47728 5 1 1 47727
0 47729 7 2 2 65222 102493
0 47730 5 1 1 102502
0 47731 7 1 2 83522 102503
0 47732 5 1 1 47731
0 47733 7 1 2 47728 47732
0 47734 5 1 1 47733
0 47735 7 1 2 102500 47734
0 47736 5 1 1 47735
0 47737 7 1 2 47725 47736
0 47738 5 1 1 47737
0 47739 7 1 2 66782 47738
0 47740 5 1 1 47739
0 47741 7 1 2 73080 100932
0 47742 5 1 1 47741
0 47743 7 1 2 70444 87040
0 47744 7 1 2 85334 47743
0 47745 5 1 1 47744
0 47746 7 1 2 47742 47745
0 47747 5 2 1 47746
0 47748 7 1 2 86166 99303
0 47749 7 1 2 102335 47748
0 47750 7 1 2 102504 47749
0 47751 5 1 1 47750
0 47752 7 1 2 47740 47751
0 47753 5 1 1 47752
0 47754 7 1 2 102490 47753
0 47755 5 1 1 47754
0 47756 7 1 2 17766 36204
0 47757 5 2 1 47756
0 47758 7 1 2 70445 102506
0 47759 5 1 1 47758
0 47760 7 1 2 75311 47759
0 47761 5 1 1 47760
0 47762 7 2 2 97653 99036
0 47763 7 2 2 78682 102508
0 47764 7 1 2 47761 102510
0 47765 5 1 1 47764
0 47766 7 1 2 97318 102268
0 47767 7 1 2 102505 47766
0 47768 5 2 1 47767
0 47769 7 1 2 47765 102512
0 47770 5 1 1 47769
0 47771 7 1 2 71874 98111
0 47772 7 1 2 96911 47771
0 47773 7 1 2 47770 47772
0 47774 5 1 1 47773
0 47775 7 1 2 47755 47774
0 47776 5 1 1 47775
0 47777 7 1 2 66295 47776
0 47778 5 1 1 47777
0 47779 7 1 2 63642 47730
0 47780 5 1 1 47779
0 47781 7 1 2 91563 38668
0 47782 5 2 1 47781
0 47783 7 1 2 65533 102514
0 47784 5 1 1 47783
0 47785 7 1 2 71990 72710
0 47786 7 2 2 72890 47785
0 47787 5 1 1 102516
0 47788 7 1 2 47784 47787
0 47789 5 1 1 47788
0 47790 7 1 2 84503 47789
0 47791 5 1 1 47790
0 47792 7 1 2 88421 93410
0 47793 5 1 1 47792
0 47794 7 1 2 47791 47793
0 47795 5 1 1 47794
0 47796 7 1 2 65852 47795
0 47797 5 1 1 47796
0 47798 7 1 2 74131 101417
0 47799 5 2 1 47798
0 47800 7 1 2 92424 102518
0 47801 5 1 1 47800
0 47802 7 1 2 73044 47801
0 47803 5 1 1 47802
0 47804 7 1 2 68481 47803
0 47805 7 1 2 47797 47804
0 47806 5 1 1 47805
0 47807 7 1 2 98668 47806
0 47808 7 1 2 47780 47807
0 47809 5 1 1 47808
0 47810 7 1 2 71875 85607
0 47811 5 1 1 47810
0 47812 7 1 2 76472 47811
0 47813 5 1 1 47812
0 47814 7 1 2 65534 47813
0 47815 5 1 1 47814
0 47816 7 1 2 78433 91929
0 47817 5 1 1 47816
0 47818 7 1 2 70446 92507
0 47819 7 1 2 47817 47818
0 47820 5 1 1 47819
0 47821 7 1 2 78132 98655
0 47822 7 1 2 47820 47821
0 47823 7 1 2 47815 47822
0 47824 5 1 1 47823
0 47825 7 1 2 47809 47824
0 47826 5 1 1 47825
0 47827 7 1 2 64392 47826
0 47828 5 1 1 47827
0 47829 7 1 2 84504 96414
0 47830 7 1 2 99248 47829
0 47831 7 1 2 101275 47830
0 47832 5 1 1 47831
0 47833 7 1 2 47828 47832
0 47834 5 1 1 47833
0 47835 7 1 2 67055 47834
0 47836 5 1 1 47835
0 47837 7 1 2 73951 89781
0 47838 5 1 1 47837
0 47839 7 1 2 97021 47838
0 47840 5 1 1 47839
0 47841 7 1 2 73045 47840
0 47842 5 1 1 47841
0 47843 7 1 2 85817 83189
0 47844 5 1 1 47843
0 47845 7 1 2 47842 47844
0 47846 5 1 1 47845
0 47847 7 1 2 68482 47846
0 47848 5 1 1 47847
0 47849 7 1 2 82501 82890
0 47850 7 1 2 86354 47849
0 47851 5 1 1 47850
0 47852 7 1 2 47848 47851
0 47853 5 1 1 47852
0 47854 7 1 2 64187 47853
0 47855 5 1 1 47854
0 47856 7 1 2 69049 101421
0 47857 5 1 1 47856
0 47858 7 1 2 88358 93294
0 47859 5 1 1 47858
0 47860 7 1 2 47857 47859
0 47861 5 1 1 47860
0 47862 7 1 2 73837 47861
0 47863 5 1 1 47862
0 47864 7 1 2 47855 47863
0 47865 5 1 1 47864
0 47866 7 1 2 65223 102382
0 47867 7 1 2 47865 47866
0 47868 5 1 1 47867
0 47869 7 1 2 47836 47868
0 47870 5 1 1 47869
0 47871 7 1 2 78718 47870
0 47872 5 1 1 47871
0 47873 7 2 2 78615 98980
0 47874 7 1 2 88495 102520
0 47875 5 1 1 47874
0 47876 7 2 2 88760 102479
0 47877 7 1 2 62642 99359
0 47878 7 1 2 102522 47877
0 47879 5 1 1 47878
0 47880 7 1 2 47875 47879
0 47881 5 1 1 47880
0 47882 7 1 2 66165 47881
0 47883 5 1 1 47882
0 47884 7 2 2 62643 92962
0 47885 7 1 2 71876 102524
0 47886 7 1 2 102523 47885
0 47887 5 1 1 47886
0 47888 7 1 2 47883 47887
0 47889 5 1 1 47888
0 47890 7 1 2 94964 47889
0 47891 5 1 1 47890
0 47892 7 1 2 79299 94381
0 47893 7 1 2 99091 47892
0 47894 7 3 2 63990 83708
0 47895 7 1 2 77604 71004
0 47896 7 1 2 102526 47895
0 47897 7 1 2 47893 47896
0 47898 5 1 1 47897
0 47899 7 1 2 47891 47898
0 47900 5 1 1 47899
0 47901 7 1 2 63643 98369
0 47902 7 1 2 47900 47901
0 47903 5 1 1 47902
0 47904 7 1 2 64188 102515
0 47905 5 1 1 47904
0 47906 7 1 2 86013 47905
0 47907 5 1 1 47906
0 47908 7 1 2 96542 97636
0 47909 7 1 2 47907 47908
0 47910 5 1 1 47909
0 47911 7 1 2 85359 75330
0 47912 7 1 2 99441 47911
0 47913 7 1 2 95293 47912
0 47914 5 1 1 47913
0 47915 7 1 2 47910 47914
0 47916 5 1 1 47915
0 47917 7 1 2 65853 47916
0 47918 5 1 1 47917
0 47919 7 1 2 79833 98889
0 47920 7 1 2 91566 47919
0 47921 5 1 1 47920
0 47922 7 1 2 47918 47921
0 47923 5 1 1 47922
0 47924 7 1 2 90725 47923
0 47925 5 1 1 47924
0 47926 7 2 2 84544 96883
0 47927 5 1 1 102529
0 47928 7 1 2 71132 79699
0 47929 7 1 2 85931 87795
0 47930 7 1 2 47928 47929
0 47931 5 1 1 47930
0 47932 7 1 2 47927 47931
0 47933 5 1 1 47932
0 47934 7 1 2 97680 47933
0 47935 5 1 1 47934
0 47936 7 1 2 62456 87080
0 47937 5 1 1 47936
0 47938 7 1 2 72924 93390
0 47939 5 1 1 47938
0 47940 7 1 2 47937 47939
0 47941 5 1 1 47940
0 47942 7 1 2 68483 99263
0 47943 7 1 2 47941 47942
0 47944 5 1 1 47943
0 47945 7 1 2 47935 47944
0 47946 5 1 1 47945
0 47947 7 1 2 68726 47946
0 47948 5 1 1 47947
0 47949 7 1 2 98190 102499
0 47950 5 1 1 47949
0 47951 7 1 2 47950 41205
0 47952 5 1 1 47951
0 47953 7 1 2 102530 47952
0 47954 5 1 1 47953
0 47955 7 1 2 47948 47954
0 47956 7 1 2 47925 47955
0 47957 5 1 1 47956
0 47958 7 1 2 65535 47957
0 47959 5 1 1 47958
0 47960 7 1 2 94382 94686
0 47961 7 1 2 102517 47960
0 47962 7 1 2 92478 47961
0 47963 5 1 1 47962
0 47964 7 1 2 47959 47963
0 47965 5 1 1 47964
0 47966 7 1 2 65224 78719
0 47967 7 1 2 47965 47966
0 47968 5 1 1 47967
0 47969 7 1 2 47903 47968
0 47970 5 1 1 47969
0 47971 7 1 2 62214 47970
0 47972 5 1 1 47971
0 47973 7 1 2 47872 47972
0 47974 5 1 1 47973
0 47975 7 1 2 83157 47974
0 47976 5 1 1 47975
0 47977 7 1 2 85335 85431
0 47978 5 1 1 47977
0 47979 7 1 2 102519 47978
0 47980 5 1 1 47979
0 47981 7 1 2 63644 47980
0 47982 5 1 1 47981
0 47983 7 1 2 68484 90818
0 47984 7 1 2 94965 47983
0 47985 5 1 1 47984
0 47986 7 1 2 47982 47985
0 47987 5 1 1 47986
0 47988 7 1 2 98981 47987
0 47989 5 1 1 47988
0 47990 7 1 2 95452 99158
0 47991 7 1 2 100345 47990
0 47992 5 1 1 47991
0 47993 7 1 2 47989 47992
0 47994 5 1 1 47993
0 47995 7 1 2 64988 47994
0 47996 5 1 1 47995
0 47997 7 2 2 84592 73952
0 47998 7 1 2 79834 102531
0 47999 7 1 2 102521 47998
0 48000 5 1 1 47999
0 48001 7 1 2 47996 48000
0 48002 5 1 1 48001
0 48003 7 1 2 62215 48002
0 48004 5 1 1 48003
0 48005 7 2 2 64393 100712
0 48006 7 3 2 71357 80682
0 48007 7 1 2 89761 102535
0 48008 5 1 1 48007
0 48009 7 2 2 73493 81501
0 48010 5 1 1 102538
0 48011 7 1 2 85336 102539
0 48012 5 1 1 48011
0 48013 7 1 2 48008 48012
0 48014 5 1 1 48013
0 48015 7 1 2 63645 48014
0 48016 5 1 1 48015
0 48017 7 2 2 70447 100474
0 48018 5 1 1 102540
0 48019 7 1 2 87604 102541
0 48020 5 1 1 48019
0 48021 7 1 2 48016 48020
0 48022 5 1 1 48021
0 48023 7 1 2 102533 48022
0 48024 5 1 1 48023
0 48025 7 1 2 48004 48024
0 48026 5 1 1 48025
0 48027 7 1 2 73046 48026
0 48028 5 1 1 48027
0 48029 7 1 2 77094 95075
0 48030 5 1 1 48029
0 48031 7 1 2 78629 78389
0 48032 5 1 1 48031
0 48033 7 1 2 48030 48032
0 48034 5 1 1 48033
0 48035 7 1 2 93411 48034
0 48036 5 1 1 48035
0 48037 7 1 2 79720 93412
0 48038 5 1 1 48037
0 48039 7 1 2 62216 92342
0 48040 7 1 2 91440 48039
0 48041 5 1 1 48040
0 48042 7 1 2 48038 48041
0 48043 5 1 1 48042
0 48044 7 1 2 87622 48043
0 48045 5 1 1 48044
0 48046 7 1 2 78630 96305
0 48047 7 1 2 92390 48046
0 48048 5 1 1 48047
0 48049 7 1 2 48045 48048
0 48050 7 1 2 48036 48049
0 48051 5 1 1 48050
0 48052 7 1 2 98982 48051
0 48053 5 1 1 48052
0 48054 7 1 2 64989 85829
0 48055 7 1 2 95294 48054
0 48056 7 1 2 99218 48055
0 48057 5 1 1 48056
0 48058 7 1 2 48053 48057
0 48059 5 1 1 48058
0 48060 7 1 2 65854 48059
0 48061 5 1 1 48060
0 48062 7 1 2 79032 85159
0 48063 5 1 1 48062
0 48064 7 1 2 88422 79516
0 48065 5 1 1 48064
0 48066 7 1 2 48065 46664
0 48067 5 1 1 48066
0 48068 7 1 2 63646 48067
0 48069 5 1 1 48068
0 48070 7 1 2 48063 48069
0 48071 5 1 1 48070
0 48072 7 1 2 73742 98439
0 48073 7 1 2 102480 48072
0 48074 7 1 2 48071 48073
0 48075 5 1 1 48074
0 48076 7 1 2 48061 48075
0 48077 7 1 2 48028 48076
0 48078 5 1 1 48077
0 48079 7 1 2 66166 48078
0 48080 5 1 1 48079
0 48081 7 1 2 84293 93605
0 48082 7 1 2 86817 48081
0 48083 5 1 1 48082
0 48084 7 1 2 73047 100346
0 48085 5 1 1 48084
0 48086 7 1 2 47664 48085
0 48087 5 1 1 48086
0 48088 7 1 2 69250 101023
0 48089 7 1 2 48087 48088
0 48090 5 1 1 48089
0 48091 7 1 2 48083 48090
0 48092 5 1 1 48091
0 48093 7 1 2 62644 48092
0 48094 5 1 1 48093
0 48095 7 1 2 76473 101461
0 48096 5 1 1 48095
0 48097 7 1 2 77106 101475
0 48098 5 1 1 48097
0 48099 7 1 2 48096 48098
0 48100 5 1 1 48099
0 48101 7 1 2 65225 48100
0 48102 5 1 1 48101
0 48103 7 1 2 76907 96682
0 48104 7 1 2 99357 48103
0 48105 5 1 1 48104
0 48106 7 1 2 48102 48105
0 48107 5 1 1 48106
0 48108 7 1 2 63991 48107
0 48109 5 1 1 48108
0 48110 7 1 2 70758 96683
0 48111 7 1 2 99318 48110
0 48112 7 1 2 88423 48111
0 48113 5 1 1 48112
0 48114 7 1 2 48109 48113
0 48115 7 1 2 48094 48114
0 48116 5 1 1 48115
0 48117 7 1 2 62895 48116
0 48118 5 1 1 48117
0 48119 7 1 2 62981 77952
0 48120 7 1 2 95305 48119
0 48121 7 1 2 100999 48120
0 48122 5 1 1 48121
0 48123 7 1 2 48118 48122
0 48124 5 1 1 48123
0 48125 7 1 2 62217 48124
0 48126 5 1 1 48125
0 48127 7 1 2 87442 84829
0 48128 7 1 2 100150 48127
0 48129 5 1 1 48128
0 48130 7 1 2 48126 48129
0 48131 5 1 1 48130
0 48132 7 1 2 64990 97720
0 48133 7 1 2 48131 48132
0 48134 5 1 1 48133
0 48135 7 1 2 48080 48134
0 48136 5 1 1 48135
0 48137 7 1 2 98417 48136
0 48138 5 1 1 48137
0 48139 7 1 2 95284 95306
0 48140 7 2 2 100234 48139
0 48141 7 1 2 73924 93878
0 48142 7 1 2 102542 48141
0 48143 5 1 1 48142
0 48144 7 1 2 70149 96454
0 48145 7 2 2 99159 48144
0 48146 7 1 2 63856 84425
0 48147 7 1 2 95447 48146
0 48148 7 1 2 102544 48147
0 48149 5 1 1 48148
0 48150 7 1 2 48143 48149
0 48151 5 1 1 48150
0 48152 7 1 2 67315 48151
0 48153 5 1 1 48152
0 48154 7 1 2 71498 84426
0 48155 7 1 2 95448 48154
0 48156 7 1 2 102545 48155
0 48157 5 1 1 48156
0 48158 7 1 2 48153 48157
0 48159 5 1 1 48158
0 48160 7 1 2 102491 48159
0 48161 5 1 1 48160
0 48162 7 1 2 98481 99094
0 48163 7 1 2 102543 48162
0 48164 5 1 1 48163
0 48165 7 1 2 48161 48164
0 48166 5 1 1 48165
0 48167 7 1 2 66296 48166
0 48168 5 1 1 48167
0 48169 7 1 2 78133 91000
0 48170 7 1 2 100235 48169
0 48171 7 1 2 98983 48170
0 48172 7 1 2 98462 48171
0 48173 5 1 1 48172
0 48174 7 1 2 48168 48173
0 48175 5 1 1 48174
0 48176 7 1 2 62218 48175
0 48177 5 1 1 48176
0 48178 7 1 2 67817 98484
0 48179 5 1 1 48178
0 48180 7 1 2 87546 100377
0 48181 5 1 1 48180
0 48182 7 1 2 48179 48181
0 48183 5 1 1 48182
0 48184 7 1 2 66167 48183
0 48185 5 1 1 48184
0 48186 7 1 2 88515 99077
0 48187 7 1 2 98856 48186
0 48188 5 1 1 48187
0 48189 7 1 2 48185 48188
0 48190 5 1 1 48189
0 48191 7 1 2 95285 97380
0 48192 7 1 2 92685 48191
0 48193 7 1 2 48190 48192
0 48194 5 1 1 48193
0 48195 7 1 2 48177 48194
0 48196 5 1 1 48195
0 48197 7 1 2 73130 48196
0 48198 5 1 1 48197
0 48199 7 1 2 75312 48018
0 48200 5 1 1 48199
0 48201 7 1 2 102511 48200
0 48202 5 1 1 48201
0 48203 7 1 2 102513 48202
0 48204 5 1 1 48203
0 48205 7 1 2 98463 48204
0 48206 5 1 1 48205
0 48207 7 1 2 81309 85105
0 48208 7 1 2 92859 48207
0 48209 7 1 2 77564 95569
0 48210 7 1 2 98529 48209
0 48211 7 1 2 48208 48210
0 48212 5 1 1 48211
0 48213 7 1 2 48206 48212
0 48214 5 1 1 48213
0 48215 7 1 2 100365 48214
0 48216 5 1 1 48215
0 48217 7 1 2 69426 48216
0 48218 7 1 2 48198 48217
0 48219 7 1 2 48138 48218
0 48220 7 1 2 47976 48219
0 48221 7 1 2 47778 48220
0 48222 7 1 2 47624 48221
0 48223 5 1 1 48222
0 48224 7 1 2 102163 48223
0 48225 7 1 2 47385 48224
0 48226 5 1 1 48225
0 48227 7 1 2 84064 99008
0 48228 7 1 2 99867 48227
0 48229 5 1 1 48228
0 48230 7 1 2 91806 102150
0 48231 5 1 1 48230
0 48232 7 1 2 64991 98456
0 48233 5 1 1 48232
0 48234 7 1 2 48231 48233
0 48235 5 1 1 48234
0 48236 7 1 2 66168 48235
0 48237 5 1 1 48236
0 48238 7 2 2 68044 81286
0 48239 7 1 2 102546 99901
0 48240 5 1 1 48239
0 48241 7 1 2 48237 48240
0 48242 5 2 1 48241
0 48243 7 1 2 79689 100258
0 48244 5 2 1 48243
0 48245 7 1 2 69427 102550
0 48246 7 1 2 102548 48245
0 48247 5 1 1 48246
0 48248 7 1 2 48229 48247
0 48249 5 1 1 48248
0 48250 7 1 2 66037 48249
0 48251 5 1 1 48250
0 48252 7 1 2 81702 92860
0 48253 7 1 2 93879 48252
0 48254 7 1 2 95961 48253
0 48255 5 1 1 48254
0 48256 7 1 2 48251 48255
0 48257 5 1 1 48256
0 48258 7 1 2 64796 48257
0 48259 5 1 1 48258
0 48260 7 3 2 93880 94451
0 48261 7 1 2 76007 99679
0 48262 7 1 2 102552 48261
0 48263 5 1 1 48262
0 48264 7 1 2 48259 48263
0 48265 5 1 1 48264
0 48266 7 1 2 61666 48265
0 48267 5 1 1 48266
0 48268 7 1 2 81389 101737
0 48269 7 1 2 102553 48268
0 48270 5 1 1 48269
0 48271 7 1 2 48267 48270
0 48272 5 1 1 48271
0 48273 7 1 2 66297 48272
0 48274 5 1 1 48273
0 48275 7 1 2 81390 99489
0 48276 7 1 2 94452 48275
0 48277 7 1 2 100604 48276
0 48278 5 1 1 48277
0 48279 7 1 2 48274 48278
0 48280 5 1 1 48279
0 48281 7 1 2 86552 48280
0 48282 5 1 1 48281
0 48283 7 2 2 64797 94676
0 48284 7 1 2 85383 102555
0 48285 5 1 1 48284
0 48286 7 1 2 78223 93394
0 48287 5 2 1 48286
0 48288 7 2 2 69629 102557
0 48289 7 1 2 66554 102559
0 48290 5 1 1 48289
0 48291 7 1 2 48285 48290
0 48292 5 1 1 48291
0 48293 7 1 2 99782 48292
0 48294 5 1 1 48293
0 48295 7 1 2 67818 91001
0 48296 7 3 2 90868 48295
0 48297 7 1 2 93284 102561
0 48298 5 1 1 48297
0 48299 7 1 2 48294 48298
0 48300 5 1 1 48299
0 48301 7 1 2 70759 48300
0 48302 5 1 1 48301
0 48303 7 2 2 69630 98317
0 48304 7 1 2 66555 102564
0 48305 5 1 1 48304
0 48306 7 1 2 45136 48305
0 48307 5 2 1 48306
0 48308 7 1 2 72467 102562
0 48309 7 1 2 102566 48308
0 48310 5 1 1 48309
0 48311 7 1 2 48302 48310
0 48312 5 1 1 48311
0 48313 7 1 2 62896 48312
0 48314 5 1 1 48313
0 48315 7 1 2 73612 90554
0 48316 7 3 2 102551 48315
0 48317 7 1 2 102568 101380
0 48318 5 1 1 48317
0 48319 7 1 2 48314 48318
0 48320 5 1 1 48319
0 48321 7 1 2 62645 48320
0 48322 5 1 1 48321
0 48323 7 2 2 72279 79546
0 48324 7 1 2 89366 84562
0 48325 7 1 2 102571 48324
0 48326 7 1 2 99783 48325
0 48327 5 1 1 48326
0 48328 7 1 2 48322 48327
0 48329 5 2 1 48328
0 48330 7 1 2 81420 92861
0 48331 5 1 1 48330
0 48332 7 1 2 63037 102547
0 48333 5 1 1 48332
0 48334 7 1 2 48331 48333
0 48335 5 1 1 48334
0 48336 7 1 2 102573 48335
0 48337 5 1 1 48336
0 48338 7 1 2 90271 93392
0 48339 5 1 1 48338
0 48340 7 1 2 82858 102560
0 48341 5 1 1 48340
0 48342 7 1 2 48339 48341
0 48343 5 1 1 48342
0 48344 7 1 2 70760 48343
0 48345 5 1 1 48344
0 48346 7 1 2 70448 98259
0 48347 5 1 1 48346
0 48348 7 1 2 48345 48347
0 48349 5 1 1 48348
0 48350 7 1 2 62897 48349
0 48351 5 1 1 48350
0 48352 7 1 2 66556 102569
0 48353 5 1 1 48352
0 48354 7 1 2 48351 48353
0 48355 5 1 1 48354
0 48356 7 1 2 62646 48355
0 48357 5 1 1 48356
0 48358 7 3 2 88901 89268
0 48359 7 1 2 73631 102575
0 48360 5 1 1 48359
0 48361 7 1 2 48357 48360
0 48362 5 1 1 48361
0 48363 7 1 2 92479 48362
0 48364 5 1 1 48363
0 48365 7 2 2 89269 99793
0 48366 7 1 2 100882 102578
0 48367 5 1 1 48366
0 48368 7 2 2 80328 93739
0 48369 7 2 2 62982 64189
0 48370 7 1 2 66557 102582
0 48371 7 1 2 102580 48370
0 48372 5 1 1 48371
0 48373 7 1 2 48367 48372
0 48374 5 1 1 48373
0 48375 7 1 2 66169 48374
0 48376 5 1 1 48375
0 48377 7 1 2 92944 100480
0 48378 7 1 2 102581 48377
0 48379 5 1 1 48378
0 48380 7 1 2 48376 48379
0 48381 5 1 1 48380
0 48382 7 1 2 75373 93821
0 48383 7 1 2 48381 48382
0 48384 5 1 1 48383
0 48385 7 1 2 48364 48384
0 48386 5 2 1 48385
0 48387 7 1 2 95820 102584
0 48388 5 1 1 48387
0 48389 7 1 2 71358 91250
0 48390 5 1 1 48389
0 48391 7 1 2 62647 94163
0 48392 5 1 1 48391
0 48393 7 1 2 48390 48392
0 48394 5 1 1 48393
0 48395 7 1 2 70449 48394
0 48396 5 1 1 48395
0 48397 7 4 2 65536 77968
0 48398 5 1 1 102586
0 48399 7 1 2 89311 102587
0 48400 5 2 1 48399
0 48401 7 1 2 48396 102590
0 48402 5 1 1 48401
0 48403 7 1 2 102004 99049
0 48404 7 1 2 48402 48403
0 48405 5 1 1 48404
0 48406 7 1 2 64190 78384
0 48407 5 1 1 48406
0 48408 7 1 2 62648 72755
0 48409 7 1 2 48407 48408
0 48410 5 1 1 48409
0 48411 7 1 2 12967 48410
0 48412 5 1 1 48411
0 48413 7 1 2 66038 48412
0 48414 5 1 1 48413
0 48415 7 1 2 91719 48414
0 48416 5 1 1 48415
0 48417 7 1 2 81421 79547
0 48418 7 1 2 92480 48417
0 48419 7 1 2 48416 48418
0 48420 5 1 1 48419
0 48421 7 1 2 48405 48420
0 48422 5 1 1 48421
0 48423 7 1 2 64575 48422
0 48424 5 1 1 48423
0 48425 7 2 2 72649 76515
0 48426 7 2 2 92481 102592
0 48427 7 1 2 83633 85018
0 48428 7 1 2 102594 48427
0 48429 5 1 1 48428
0 48430 7 1 2 48424 48429
0 48431 5 1 1 48430
0 48432 7 1 2 76191 48431
0 48433 5 1 1 48432
0 48434 7 4 2 66298 63992
0 48435 7 2 2 69428 102596
0 48436 7 1 2 100883 102600
0 48437 5 1 1 48436
0 48438 7 1 2 61402 88440
0 48439 7 1 2 102558 48438
0 48440 5 1 1 48439
0 48441 7 1 2 48437 48440
0 48442 5 1 1 48441
0 48443 7 1 2 81948 48442
0 48444 5 1 1 48443
0 48445 7 1 2 91135 100003
0 48446 5 1 1 48445
0 48447 7 1 2 90115 99490
0 48448 5 1 1 48447
0 48449 7 1 2 48446 48448
0 48450 5 1 1 48449
0 48451 7 1 2 102556 48450
0 48452 5 1 1 48451
0 48453 7 1 2 48444 48452
0 48454 5 2 1 48453
0 48455 7 1 2 62649 102602
0 48456 5 1 1 48455
0 48457 7 2 2 73632 100042
0 48458 5 1 1 102604
0 48459 7 1 2 48456 48458
0 48460 5 1 1 48459
0 48461 7 1 2 102549 48460
0 48462 5 1 1 48461
0 48463 7 1 2 72468 94517
0 48464 5 1 1 48463
0 48465 7 2 2 70960 73525
0 48466 5 1 1 102606
0 48467 7 1 2 48464 48466
0 48468 5 1 1 48467
0 48469 7 1 2 91924 99050
0 48470 7 1 2 48468 48469
0 48471 5 1 1 48470
0 48472 7 1 2 93881 101443
0 48473 5 2 1 48472
0 48474 7 1 2 92648 101451
0 48475 5 1 1 48474
0 48476 7 1 2 102608 48475
0 48477 5 4 1 48476
0 48478 7 4 2 71359 86706
0 48479 5 1 1 102614
0 48480 7 1 2 74691 48479
0 48481 5 2 1 48480
0 48482 7 2 2 70450 102618
0 48483 5 1 1 102620
0 48484 7 1 2 81422 102621
0 48485 7 1 2 102610 48484
0 48486 5 1 1 48485
0 48487 7 1 2 48471 48486
0 48488 5 1 1 48487
0 48489 7 1 2 64798 48488
0 48490 5 1 1 48489
0 48491 7 1 2 102609 41267
0 48492 5 1 1 48491
0 48493 7 1 2 92915 98232
0 48494 7 1 2 48492 48493
0 48495 5 1 1 48494
0 48496 7 1 2 48490 48495
0 48497 5 1 1 48496
0 48498 7 1 2 64576 48497
0 48499 5 1 1 48498
0 48500 7 1 2 48462 48499
0 48501 5 1 1 48500
0 48502 7 1 2 62898 48501
0 48503 5 1 1 48502
0 48504 7 1 2 48433 48503
0 48505 7 1 2 48388 48504
0 48506 7 1 2 48337 48505
0 48507 7 1 2 48282 48506
0 48508 5 1 1 48507
0 48509 7 1 2 75839 48508
0 48510 5 1 1 48509
0 48511 7 1 2 92558 95197
0 48512 5 1 1 48511
0 48513 7 1 2 45520 48512
0 48514 5 1 1 48513
0 48515 7 1 2 102574 48514
0 48516 5 1 1 48515
0 48517 7 1 2 63204 95198
0 48518 5 1 1 48517
0 48519 7 1 2 25801 48518
0 48520 5 3 1 48519
0 48521 7 1 2 102585 102622
0 48522 5 1 1 48521
0 48523 7 1 2 62899 102603
0 48524 5 1 1 48523
0 48525 7 1 2 99027 102570
0 48526 5 1 1 48525
0 48527 7 1 2 48524 48526
0 48528 5 1 1 48527
0 48529 7 1 2 62650 48528
0 48530 5 1 1 48529
0 48531 7 1 2 62900 102605
0 48532 5 1 1 48531
0 48533 7 1 2 48530 48532
0 48534 5 1 1 48533
0 48535 7 1 2 99291 99776
0 48536 5 1 1 48535
0 48537 7 1 2 81659 93577
0 48538 7 1 2 98339 48537
0 48539 5 1 1 48538
0 48540 7 1 2 48536 48539
0 48541 5 1 1 48540
0 48542 7 1 2 66170 48541
0 48543 5 1 1 48542
0 48544 7 1 2 80037 91872
0 48545 7 1 2 102186 48544
0 48546 5 1 1 48545
0 48547 7 1 2 48543 48546
0 48548 5 1 1 48547
0 48549 7 1 2 48534 48548
0 48550 5 1 1 48549
0 48551 7 1 2 48522 48550
0 48552 7 1 2 48516 48551
0 48553 5 1 1 48552
0 48554 7 1 2 101531 48553
0 48555 5 1 1 48554
0 48556 7 1 2 66558 102623
0 48557 5 1 1 48556
0 48558 7 1 2 74340 90536
0 48559 5 1 1 48558
0 48560 7 1 2 48557 48559
0 48561 5 2 1 48560
0 48562 7 1 2 99051 102625
0 48563 5 1 1 48562
0 48564 7 2 2 75784 92894
0 48565 7 1 2 92482 102627
0 48566 5 1 1 48565
0 48567 7 1 2 48563 48566
0 48568 5 1 1 48567
0 48569 7 3 2 64577 48568
0 48570 7 1 2 88952 101343
0 48571 5 1 1 48570
0 48572 7 1 2 91246 95792
0 48573 5 7 1 48572
0 48574 7 1 2 88978 102632
0 48575 5 1 1 48574
0 48576 7 1 2 88953 94508
0 48577 5 1 1 48576
0 48578 7 1 2 48575 48577
0 48579 5 1 1 48578
0 48580 7 1 2 63993 48579
0 48581 5 1 1 48580
0 48582 7 1 2 48571 48581
0 48583 5 1 1 48582
0 48584 7 1 2 102629 48583
0 48585 5 1 1 48584
0 48586 7 1 2 69429 102595
0 48587 5 1 1 48586
0 48588 7 1 2 89564 99052
0 48589 5 1 1 48588
0 48590 7 1 2 48587 48589
0 48591 5 1 1 48590
0 48592 7 1 2 102626 48591
0 48593 5 1 1 48592
0 48594 7 1 2 89565 92483
0 48595 5 1 1 48594
0 48596 7 2 2 92649 100299
0 48597 7 1 2 102593 102639
0 48598 5 1 1 48597
0 48599 7 1 2 48595 48598
0 48600 5 1 1 48599
0 48601 7 1 2 102628 48600
0 48602 5 1 1 48601
0 48603 7 1 2 48593 48602
0 48604 5 1 1 48603
0 48605 7 1 2 63994 48604
0 48606 5 1 1 48605
0 48607 7 1 2 102630 102633
0 48608 5 1 1 48607
0 48609 7 1 2 48606 48608
0 48610 5 1 1 48609
0 48611 7 1 2 62651 88979
0 48612 7 1 2 48610 48611
0 48613 5 1 1 48612
0 48614 7 1 2 48585 48613
0 48615 5 1 1 48614
0 48616 7 1 2 64799 48615
0 48617 5 1 1 48616
0 48618 7 1 2 61667 102624
0 48619 5 1 1 48618
0 48620 7 1 2 88879 75785
0 48621 5 1 1 48620
0 48622 7 1 2 48619 48621
0 48623 5 1 1 48622
0 48624 7 1 2 92484 48623
0 48625 5 1 1 48624
0 48626 7 1 2 66783 96796
0 48627 7 1 2 99053 48626
0 48628 5 1 1 48627
0 48629 7 1 2 48625 48628
0 48630 5 1 1 48629
0 48631 7 1 2 88954 78011
0 48632 5 1 1 48631
0 48633 7 2 2 72582 78450
0 48634 5 1 1 102641
0 48635 7 1 2 77828 48634
0 48636 5 1 1 48635
0 48637 7 1 2 88980 48636
0 48638 5 1 1 48637
0 48639 7 1 2 48632 48638
0 48640 5 1 1 48639
0 48641 7 1 2 73344 48640
0 48642 5 1 1 48641
0 48643 7 1 2 65855 88959
0 48644 5 1 1 48643
0 48645 7 1 2 81330 77789
0 48646 5 1 1 48645
0 48647 7 1 2 48644 48646
0 48648 5 1 1 48647
0 48649 7 1 2 71360 48648
0 48650 5 1 1 48649
0 48651 7 1 2 62652 90488
0 48652 7 1 2 82174 48651
0 48653 5 1 1 48652
0 48654 7 1 2 48650 48653
0 48655 5 1 1 48654
0 48656 7 1 2 64191 48655
0 48657 5 1 1 48656
0 48658 7 1 2 48642 48657
0 48659 5 1 1 48658
0 48660 7 1 2 79378 48659
0 48661 7 1 2 48630 48660
0 48662 5 1 1 48661
0 48663 7 1 2 48617 48662
0 48664 5 1 1 48663
0 48665 7 1 2 70451 48664
0 48666 5 1 1 48665
0 48667 7 1 2 82552 89762
0 48668 7 1 2 102607 48667
0 48669 7 1 2 102631 48668
0 48670 5 1 1 48669
0 48671 7 1 2 48666 48670
0 48672 7 1 2 48555 48671
0 48673 7 1 2 48510 48672
0 48674 5 1 1 48673
0 48675 7 1 2 65226 48674
0 48676 5 1 1 48675
0 48677 7 1 2 102579 100477
0 48678 5 1 1 48677
0 48679 7 2 2 84412 99741
0 48680 7 1 2 89522 102643
0 48681 5 1 1 48680
0 48682 7 1 2 48678 48681
0 48683 5 1 1 48682
0 48684 7 1 2 63995 48683
0 48685 5 1 1 48684
0 48686 7 1 2 102634 102644
0 48687 5 1 1 48686
0 48688 7 1 2 48685 48687
0 48689 5 1 1 48688
0 48690 7 1 2 66171 48689
0 48691 5 1 1 48690
0 48692 7 1 2 84386 71598
0 48693 5 1 1 48692
0 48694 7 1 2 95793 48693
0 48695 5 1 1 48694
0 48696 7 4 2 64800 94719
0 48697 7 1 2 92963 102645
0 48698 7 1 2 48695 48697
0 48699 5 1 1 48698
0 48700 7 1 2 48691 48699
0 48701 5 1 1 48700
0 48702 7 1 2 62653 48701
0 48703 5 1 1 48702
0 48704 7 3 2 93882 94720
0 48705 7 2 2 81073 102649
0 48706 7 1 2 102635 102652
0 48707 5 1 1 48706
0 48708 7 1 2 48703 48707
0 48709 5 1 1 48708
0 48710 7 1 2 70452 48709
0 48711 5 1 1 48710
0 48712 7 3 2 73081 89501
0 48713 5 1 1 102654
0 48714 7 1 2 62654 102653
0 48715 7 1 2 102655 48714
0 48716 5 1 1 48715
0 48717 7 1 2 48711 48716
0 48718 5 1 1 48717
0 48719 7 1 2 93822 48718
0 48720 5 1 1 48719
0 48721 7 1 2 78451 87326
0 48722 5 1 1 48721
0 48723 7 1 2 14352 48722
0 48724 5 1 1 48723
0 48725 7 1 2 66039 48724
0 48726 5 1 1 48725
0 48727 7 1 2 75551 98256
0 48728 5 1 1 48727
0 48729 7 1 2 48726 48728
0 48730 5 1 1 48729
0 48731 7 1 2 69050 48730
0 48732 5 1 1 48731
0 48733 7 3 2 73584 90272
0 48734 5 1 1 102657
0 48735 7 1 2 64192 102658
0 48736 5 1 1 48735
0 48737 7 1 2 100892 48736
0 48738 5 2 1 48737
0 48739 7 1 2 65856 102660
0 48740 5 1 1 48739
0 48741 7 1 2 48732 48740
0 48742 5 1 1 48741
0 48743 7 1 2 73345 48742
0 48744 5 1 1 48743
0 48745 7 1 2 102576 102615
0 48746 5 1 1 48745
0 48747 7 1 2 48744 48746
0 48748 5 1 1 48747
0 48749 7 1 2 70453 48748
0 48750 5 1 1 48749
0 48751 7 1 2 12419 87335
0 48752 5 4 1 48751
0 48753 7 1 2 73082 93234
0 48754 7 1 2 102662 48753
0 48755 5 1 1 48754
0 48756 7 1 2 48750 48755
0 48757 5 1 1 48756
0 48758 7 1 2 92485 48757
0 48759 5 1 1 48758
0 48760 7 1 2 48720 48759
0 48761 5 1 1 48760
0 48762 7 1 2 90203 48761
0 48763 5 1 1 48762
0 48764 7 1 2 100878 99731
0 48765 5 1 1 48764
0 48766 7 1 2 90497 90947
0 48767 5 1 1 48766
0 48768 7 1 2 48765 48767
0 48769 5 1 1 48768
0 48770 7 1 2 63996 48769
0 48771 5 1 1 48770
0 48772 7 3 2 62983 99753
0 48773 5 1 1 102666
0 48774 7 1 2 86707 102667
0 48775 5 1 1 48774
0 48776 7 1 2 48771 48775
0 48777 5 1 1 48776
0 48778 7 1 2 66172 48777
0 48779 5 1 1 48778
0 48780 7 1 2 69051 80180
0 48781 5 1 1 48780
0 48782 7 1 2 77843 48781
0 48783 5 1 1 48782
0 48784 7 1 2 91376 102189
0 48785 7 1 2 48783 48784
0 48786 5 1 1 48785
0 48787 7 1 2 48779 48786
0 48788 5 1 1 48787
0 48789 7 1 2 62655 48788
0 48790 5 1 1 48789
0 48791 7 1 2 63997 86708
0 48792 7 1 2 99784 48791
0 48793 5 1 1 48792
0 48794 7 1 2 48790 48793
0 48795 5 1 1 48794
0 48796 7 1 2 70454 48795
0 48797 5 1 1 48796
0 48798 7 1 2 72480 73106
0 48799 5 2 1 48798
0 48800 7 1 2 84368 102669
0 48801 5 1 1 48800
0 48802 7 1 2 72413 94672
0 48803 5 1 1 48802
0 48804 7 1 2 48801 48803
0 48805 5 1 1 48804
0 48806 7 1 2 99785 48805
0 48807 5 1 1 48806
0 48808 7 1 2 62901 91136
0 48809 5 1 1 48808
0 48810 7 1 2 14151 48809
0 48811 5 1 1 48810
0 48812 7 1 2 102563 48811
0 48813 5 1 1 48812
0 48814 7 1 2 48807 48813
0 48815 5 1 1 48814
0 48816 7 1 2 62656 48815
0 48817 5 1 1 48816
0 48818 7 1 2 72192 78381
0 48819 5 2 1 48818
0 48820 7 1 2 65857 84369
0 48821 5 1 1 48820
0 48822 7 1 2 102671 48821
0 48823 5 1 1 48822
0 48824 7 1 2 73613 99786
0 48825 7 1 2 48823 48824
0 48826 5 1 1 48825
0 48827 7 1 2 48817 48826
0 48828 5 1 1 48827
0 48829 7 1 2 86986 48828
0 48830 5 1 1 48829
0 48831 7 1 2 65537 98734
0 48832 7 1 2 93426 48831
0 48833 7 1 2 101088 48832
0 48834 5 1 1 48833
0 48835 7 1 2 48830 48834
0 48836 7 1 2 48797 48835
0 48837 5 1 1 48836
0 48838 7 1 2 96038 48837
0 48839 5 1 1 48838
0 48840 7 1 2 73346 87499
0 48841 7 1 2 102221 48840
0 48842 7 1 2 102554 48841
0 48843 5 1 1 48842
0 48844 7 1 2 48839 48843
0 48845 5 1 1 48844
0 48846 7 1 2 98396 48845
0 48847 5 1 1 48846
0 48848 7 1 2 66173 99983
0 48849 5 1 1 48848
0 48850 7 1 2 68241 81660
0 48851 7 2 2 99902 48850
0 48852 5 1 1 102673
0 48853 7 1 2 48849 48852
0 48854 5 1 1 48853
0 48855 7 6 2 64801 87482
0 48856 5 2 1 102675
0 48857 7 2 2 63998 72469
0 48858 5 1 1 102683
0 48859 7 1 2 62657 102670
0 48860 5 1 1 48859
0 48861 7 1 2 48858 48860
0 48862 5 6 1 48861
0 48863 7 1 2 102676 102685
0 48864 5 1 1 48863
0 48865 7 2 2 70455 99393
0 48866 5 1 1 102691
0 48867 7 1 2 73347 102692
0 48868 5 1 1 48867
0 48869 7 1 2 48864 48868
0 48870 5 1 1 48869
0 48871 7 1 2 72650 48870
0 48872 5 1 1 48871
0 48873 7 1 2 102591 48483
0 48874 5 1 1 48873
0 48875 7 1 2 96039 48874
0 48876 5 1 1 48875
0 48877 7 1 2 91129 101256
0 48878 5 1 1 48877
0 48879 7 1 2 80796 87236
0 48880 7 1 2 83723 48879
0 48881 5 1 1 48880
0 48882 7 1 2 48878 48881
0 48883 5 1 1 48882
0 48884 7 1 2 70456 48883
0 48885 5 1 1 48884
0 48886 7 1 2 48876 48885
0 48887 7 1 2 48872 48886
0 48888 5 1 1 48887
0 48889 7 1 2 99491 48888
0 48890 5 1 1 48889
0 48891 7 1 2 96040 98318
0 48892 5 1 1 48891
0 48893 7 1 2 61668 100921
0 48894 5 1 1 48893
0 48895 7 1 2 48892 48894
0 48896 5 2 1 48895
0 48897 7 1 2 65858 102693
0 48898 5 1 1 48897
0 48899 7 1 2 86987 84638
0 48900 5 1 1 48899
0 48901 7 1 2 48898 48900
0 48902 5 1 1 48901
0 48903 7 1 2 70457 48902
0 48904 5 1 1 48903
0 48905 7 1 2 91133 102159
0 48906 5 1 1 48905
0 48907 7 1 2 48904 48906
0 48908 5 1 1 48907
0 48909 7 1 2 48908 100050
0 48910 5 1 1 48909
0 48911 7 1 2 48890 48910
0 48912 5 1 1 48911
0 48913 7 1 2 48854 48912
0 48914 5 1 1 48913
0 48915 7 1 2 64992 48914
0 48916 7 1 2 48847 48915
0 48917 7 1 2 48763 48916
0 48918 5 1 1 48917
0 48919 7 1 2 78810 102611
0 48920 5 1 1 48919
0 48921 7 1 2 101337 101385
0 48922 5 1 1 48921
0 48923 7 1 2 48920 48922
0 48924 5 1 1 48923
0 48925 7 1 2 65859 48924
0 48926 5 1 1 48925
0 48927 7 1 2 64802 99468
0 48928 5 2 1 48927
0 48929 7 1 2 92486 96475
0 48930 5 1 1 48929
0 48931 7 1 2 102695 48930
0 48932 5 1 1 48931
0 48933 7 1 2 85409 48932
0 48934 5 1 1 48933
0 48935 7 1 2 71133 88256
0 48936 7 1 2 102612 48935
0 48937 5 1 1 48936
0 48938 7 1 2 48934 48937
0 48939 7 1 2 48926 48938
0 48940 5 1 1 48939
0 48941 7 1 2 64578 48940
0 48942 5 1 1 48941
0 48943 7 1 2 62984 43603
0 48944 5 1 1 48943
0 48945 7 1 2 67819 100758
0 48946 5 1 1 48945
0 48947 7 3 2 48944 48946
0 48948 7 1 2 66174 102697
0 48949 5 1 1 48948
0 48950 7 1 2 102243 98857
0 48951 5 1 1 48950
0 48952 7 1 2 48949 48951
0 48953 5 2 1 48952
0 48954 7 1 2 102161 102700
0 48955 5 1 1 48954
0 48956 7 3 2 69631 92650
0 48957 7 1 2 84768 102702
0 48958 7 1 2 99387 48957
0 48959 5 1 1 48958
0 48960 7 1 2 48955 48959
0 48961 5 1 1 48960
0 48962 7 1 2 99717 48961
0 48963 5 1 1 48962
0 48964 7 1 2 48942 48963
0 48965 5 1 1 48964
0 48966 7 1 2 83158 73348
0 48967 7 1 2 48965 48966
0 48968 5 1 1 48967
0 48969 7 2 2 64579 86709
0 48970 7 1 2 87025 91661
0 48971 7 1 2 102705 48970
0 48972 7 1 2 102613 48971
0 48973 5 1 1 48972
0 48974 7 1 2 48968 48973
0 48975 5 1 1 48974
0 48976 7 1 2 70458 48975
0 48977 5 1 1 48976
0 48978 7 1 2 91945 92487
0 48979 5 1 1 48978
0 48980 7 1 2 102696 48979
0 48981 5 1 1 48980
0 48982 7 2 2 64193 88382
0 48983 7 1 2 75374 102707
0 48984 7 1 2 99478 48983
0 48985 7 1 2 48981 48984
0 48986 5 1 1 48985
0 48987 7 1 2 69845 48986
0 48988 7 1 2 48977 48987
0 48989 5 1 1 48988
0 48990 7 1 2 88714 48989
0 48991 7 1 2 48918 48990
0 48992 5 1 1 48991
0 48993 7 1 2 48676 48992
0 48994 5 1 1 48993
0 48995 7 1 2 94383 48994
0 48996 5 1 1 48995
0 48997 7 1 2 1458 28482
0 48998 5 1 1 48997
0 48999 7 1 2 62902 48998
0 49000 5 1 1 48999
0 49001 7 2 2 65538 94453
0 49002 7 1 2 69846 102709
0 49003 5 1 1 49002
0 49004 7 1 2 49000 49003
0 49005 5 1 1 49004
0 49006 7 1 2 75786 49005
0 49007 5 1 1 49006
0 49008 7 1 2 75678 73838
0 49009 7 1 2 77136 49008
0 49010 5 1 1 49009
0 49011 7 1 2 49007 49010
0 49012 5 1 1 49011
0 49013 7 1 2 63999 49012
0 49014 5 1 1 49013
0 49015 7 1 2 65227 19239
0 49016 5 1 1 49015
0 49017 7 1 2 2306 94509
0 49018 5 1 1 49017
0 49019 7 1 2 49016 49018
0 49020 5 2 1 49019
0 49021 7 1 2 83869 102711
0 49022 5 1 1 49021
0 49023 7 1 2 49014 49022
0 49024 5 1 1 49023
0 49025 7 1 2 99595 49024
0 49026 5 1 1 49025
0 49027 7 1 2 64000 78336
0 49028 5 2 1 49027
0 49029 7 1 2 80543 102713
0 49030 5 1 1 49029
0 49031 7 2 2 65228 49030
0 49032 5 1 1 102715
0 49033 7 2 2 74495 100879
0 49034 5 1 1 102717
0 49035 7 1 2 65229 77991
0 49036 5 1 1 49035
0 49037 7 1 2 49034 49036
0 49038 5 2 1 49037
0 49039 7 1 2 62903 102719
0 49040 5 1 1 49039
0 49041 7 1 2 49032 49040
0 49042 5 1 1 49041
0 49043 7 1 2 69430 83523
0 49044 7 1 2 98048 49043
0 49045 7 1 2 49042 49044
0 49046 5 1 1 49045
0 49047 7 1 2 49026 49046
0 49048 5 1 1 49047
0 49049 7 1 2 62658 49048
0 49050 5 1 1 49049
0 49051 7 1 2 99596 102712
0 49052 5 1 1 49051
0 49053 7 1 2 99676 101100
0 49054 5 1 1 49053
0 49055 7 1 2 49052 49054
0 49056 5 1 1 49055
0 49057 7 1 2 64001 49056
0 49058 5 1 1 49057
0 49059 7 1 2 95172 99658
0 49060 5 1 1 49059
0 49061 7 1 2 80549 99597
0 49062 5 1 1 49061
0 49063 7 1 2 49060 49062
0 49064 5 1 1 49063
0 49065 7 1 2 62904 49064
0 49066 5 1 1 49065
0 49067 7 2 2 64580 99063
0 49068 5 1 1 102721
0 49069 7 1 2 70761 102722
0 49070 5 1 1 49069
0 49071 7 1 2 49066 49070
0 49072 5 1 1 49071
0 49073 7 1 2 65230 49072
0 49074 5 1 1 49073
0 49075 7 1 2 49058 49074
0 49076 5 1 1 49075
0 49077 7 1 2 83870 49076
0 49078 5 1 1 49077
0 49079 7 1 2 49050 49078
0 49080 5 1 1 49079
0 49081 7 1 2 64803 49080
0 49082 5 1 1 49081
0 49083 7 1 2 99659 100412
0 49084 5 2 1 49083
0 49085 7 1 2 102723 100282
0 49086 5 1 1 49085
0 49087 7 1 2 65860 49086
0 49088 5 1 1 49087
0 49089 7 1 2 78452 101618
0 49090 5 1 1 49089
0 49091 7 1 2 49088 49090
0 49092 5 1 1 49091
0 49093 7 1 2 73349 49092
0 49094 5 1 1 49093
0 49095 7 1 2 63038 76277
0 49096 7 1 2 102706 49095
0 49097 5 1 1 49096
0 49098 7 1 2 49094 49097
0 49099 5 1 1 49098
0 49100 7 1 2 68485 49099
0 49101 5 1 1 49100
0 49102 7 1 2 87021 82446
0 49103 7 1 2 99629 49102
0 49104 5 1 1 49103
0 49105 7 1 2 49101 49104
0 49106 5 1 1 49105
0 49107 7 1 2 102294 49106
0 49108 5 1 1 49107
0 49109 7 2 2 67899 96907
0 49110 5 1 1 102725
0 49111 7 1 2 100283 49110
0 49112 5 1 1 49111
0 49113 7 1 2 72858 49112
0 49114 5 1 1 49113
0 49115 7 1 2 78317 99660
0 49116 5 1 1 49115
0 49117 7 1 2 101620 49116
0 49118 5 1 1 49117
0 49119 7 1 2 86065 49118
0 49120 5 1 1 49119
0 49121 7 1 2 49114 49120
0 49122 5 1 1 49121
0 49123 7 1 2 97171 49122
0 49124 5 1 1 49123
0 49125 7 1 2 49108 49124
0 49126 7 1 2 49082 49125
0 49127 5 1 1 49126
0 49128 7 1 2 77260 49127
0 49129 5 1 1 49128
0 49130 7 1 2 99842 102720
0 49131 5 1 1 49130
0 49132 7 1 2 97165 102718
0 49133 5 1 1 49132
0 49134 7 1 2 49131 49133
0 49135 5 1 1 49134
0 49136 7 1 2 62905 49135
0 49137 5 1 1 49136
0 49138 7 1 2 99843 102716
0 49139 5 1 1 49138
0 49140 7 1 2 49137 49139
0 49141 5 1 1 49140
0 49142 7 1 2 62659 49141
0 49143 5 1 1 49142
0 49144 7 2 2 84266 96159
0 49145 5 1 1 102727
0 49146 7 1 2 84370 86507
0 49147 5 1 1 49146
0 49148 7 1 2 5248 49147
0 49149 5 1 1 49148
0 49150 7 1 2 81149 49149
0 49151 5 1 1 49150
0 49152 7 1 2 49145 49151
0 49153 5 1 1 49152
0 49154 7 1 2 80713 49153
0 49155 5 1 1 49154
0 49156 7 1 2 67056 78337
0 49157 5 2 1 49156
0 49158 7 1 2 102729 30192
0 49159 5 1 1 49158
0 49160 7 1 2 4573 97172
0 49161 7 1 2 49159 49160
0 49162 5 1 1 49161
0 49163 7 1 2 49155 49162
0 49164 7 1 2 49143 49163
0 49165 5 1 1 49164
0 49166 7 2 2 69431 49165
0 49167 7 1 2 100668 102731
0 49168 5 1 1 49167
0 49169 7 1 2 49129 49168
0 49170 5 1 1 49169
0 49171 7 1 2 61403 49170
0 49172 5 1 1 49171
0 49173 7 2 2 64993 99830
0 49174 7 1 2 67057 93719
0 49175 5 1 1 49174
0 49176 7 1 2 85949 97265
0 49177 5 1 1 49176
0 49178 7 1 2 73350 49177
0 49179 5 1 1 49178
0 49180 7 1 2 74483 49179
0 49181 5 1 1 49180
0 49182 7 1 2 65539 49181
0 49183 5 1 1 49182
0 49184 7 1 2 76254 91716
0 49185 5 1 1 49184
0 49186 7 1 2 72873 49185
0 49187 5 1 1 49186
0 49188 7 1 2 75552 49187
0 49189 5 1 1 49188
0 49190 7 1 2 90069 49189
0 49191 7 1 2 49183 49190
0 49192 5 1 1 49191
0 49193 7 1 2 68486 49192
0 49194 5 1 1 49193
0 49195 7 1 2 49175 49194
0 49196 5 1 1 49195
0 49197 7 1 2 102733 49196
0 49198 5 1 1 49197
0 49199 7 3 2 69847 80489
0 49200 7 1 2 86513 94132
0 49201 5 1 1 49200
0 49202 7 1 2 85464 49201
0 49203 5 1 1 49202
0 49204 7 2 2 102735 49203
0 49205 7 1 2 98049 102738
0 49206 5 1 1 49205
0 49207 7 1 2 49198 49206
0 49208 5 1 1 49207
0 49209 7 1 2 61404 49208
0 49210 5 1 1 49209
0 49211 7 3 2 62219 93763
0 49212 7 1 2 102740 102739
0 49213 5 1 1 49212
0 49214 7 1 2 65231 49213
0 49215 7 1 2 49210 49214
0 49216 5 1 1 49215
0 49217 7 1 2 100107 102736
0 49218 5 1 1 49217
0 49219 7 1 2 74341 102734
0 49220 5 1 1 49219
0 49221 7 1 2 49218 49220
0 49222 5 1 1 49221
0 49223 7 1 2 61405 49222
0 49224 5 1 1 49223
0 49225 7 2 2 82788 74474
0 49226 7 1 2 101881 102743
0 49227 5 1 1 49226
0 49228 7 1 2 49224 49227
0 49229 5 1 1 49228
0 49230 7 1 2 72193 49229
0 49231 5 1 1 49230
0 49232 7 2 2 66040 93823
0 49233 7 1 2 80102 83871
0 49234 7 1 2 102745 49233
0 49235 5 1 1 49234
0 49236 7 1 2 49231 49235
0 49237 5 1 1 49236
0 49238 7 1 2 76720 49237
0 49239 5 1 1 49238
0 49240 7 1 2 75168 93824
0 49241 7 1 2 96508 49240
0 49242 7 1 2 95714 49241
0 49243 5 1 1 49242
0 49244 7 1 2 70150 49243
0 49245 7 1 2 49239 49244
0 49246 5 1 1 49245
0 49247 7 1 2 69432 49246
0 49248 7 1 2 49216 49247
0 49249 5 1 1 49248
0 49250 7 2 2 79379 90622
0 49251 7 1 2 89732 91627
0 49252 5 1 1 49251
0 49253 7 1 2 74496 101027
0 49254 5 1 1 49253
0 49255 7 1 2 75293 76721
0 49256 5 1 1 49255
0 49257 7 1 2 2321 49256
0 49258 5 1 1 49257
0 49259 7 1 2 62906 49258
0 49260 5 1 1 49259
0 49261 7 1 2 76959 49260
0 49262 7 1 2 49254 49261
0 49263 5 1 1 49262
0 49264 7 1 2 62660 49263
0 49265 5 1 1 49264
0 49266 7 1 2 49252 49265
0 49267 5 1 1 49266
0 49268 7 1 2 75787 49267
0 49269 5 1 1 49268
0 49270 7 1 2 70459 94999
0 49271 5 1 1 49270
0 49272 7 1 2 75735 96247
0 49273 5 1 1 49272
0 49274 7 1 2 49271 49273
0 49275 5 1 1 49274
0 49276 7 1 2 84670 49275
0 49277 5 1 1 49276
0 49278 7 1 2 85149 101227
0 49279 5 2 1 49278
0 49280 7 1 2 102749 100310
0 49281 5 2 1 49280
0 49282 7 1 2 62907 102750
0 49283 5 1 1 49282
0 49284 7 1 2 70151 49283
0 49285 7 1 2 102751 49284
0 49286 5 1 1 49285
0 49287 7 1 2 49277 49286
0 49288 7 1 2 49269 49287
0 49289 5 1 1 49288
0 49290 7 1 2 69848 49289
0 49291 5 1 1 49290
0 49292 7 1 2 96848 97139
0 49293 5 1 1 49292
0 49294 7 1 2 49291 49293
0 49295 5 1 1 49294
0 49296 7 1 2 102747 49295
0 49297 5 1 1 49296
0 49298 7 1 2 49249 49297
0 49299 5 1 1 49298
0 49300 7 1 2 76192 49299
0 49301 5 1 1 49300
0 49302 7 1 2 100755 102732
0 49303 5 1 1 49302
0 49304 7 1 2 81150 93726
0 49305 5 1 1 49304
0 49306 7 1 2 4576 49305
0 49307 5 1 1 49306
0 49308 7 1 2 100766 49307
0 49309 5 1 1 49308
0 49310 7 3 2 100608 99205
0 49311 7 1 2 81151 95173
0 49312 5 1 1 49311
0 49313 7 1 2 91821 96160
0 49314 5 1 1 49313
0 49315 7 1 2 49312 49314
0 49316 5 1 1 49315
0 49317 7 1 2 102753 49316
0 49318 5 1 1 49317
0 49319 7 1 2 49309 49318
0 49320 5 1 1 49319
0 49321 7 1 2 94948 49320
0 49322 5 1 1 49321
0 49323 7 1 2 49303 49322
0 49324 7 1 2 49301 49323
0 49325 7 1 2 49172 49324
0 49326 5 1 1 49325
0 49327 7 1 2 83159 49326
0 49328 5 1 1 49327
0 49329 7 9 2 64581 90623
0 49330 5 1 1 102756
0 49331 7 1 2 70460 101964
0 49332 5 3 1 49331
0 49333 7 1 2 36067 102765
0 49334 5 1 1 49333
0 49335 7 1 2 87623 49334
0 49336 5 1 1 49335
0 49337 7 1 2 85401 2249
0 49338 5 1 1 49337
0 49339 7 1 2 67058 49338
0 49340 5 1 1 49339
0 49341 7 1 2 62908 102619
0 49342 5 2 1 49341
0 49343 7 1 2 77969 77277
0 49344 5 1 1 49343
0 49345 7 1 2 102768 49344
0 49346 5 1 1 49345
0 49347 7 1 2 78420 49346
0 49348 5 1 1 49347
0 49349 7 1 2 49340 49348
0 49350 5 1 1 49349
0 49351 7 1 2 69849 49350
0 49352 5 1 1 49351
0 49353 7 1 2 75375 97140
0 49354 5 1 1 49353
0 49355 7 3 2 77384 80303
0 49356 7 1 2 72651 102770
0 49357 5 2 1 49356
0 49358 7 1 2 72652 76722
0 49359 7 1 2 86323 49358
0 49360 5 1 1 49359
0 49361 7 1 2 68487 49360
0 49362 7 1 2 102773 49361
0 49363 7 1 2 49354 49362
0 49364 7 1 2 49352 49363
0 49365 5 1 1 49364
0 49366 7 1 2 77340 18647
0 49367 5 1 1 49366
0 49368 7 1 2 62661 49367
0 49369 5 2 1 49368
0 49370 7 1 2 65232 86508
0 49371 5 1 1 49370
0 49372 7 1 2 102775 49371
0 49373 5 1 1 49372
0 49374 7 1 2 72653 49373
0 49375 5 1 1 49374
0 49376 7 1 2 77341 26290
0 49377 5 1 1 49376
0 49378 7 1 2 74989 49377
0 49379 5 1 1 49378
0 49380 7 1 2 76960 11844
0 49381 5 1 1 49380
0 49382 7 1 2 72726 49381
0 49383 5 1 1 49382
0 49384 7 1 2 74735 74501
0 49385 5 1 1 49384
0 49386 7 1 2 76961 49385
0 49387 5 1 1 49386
0 49388 7 1 2 71599 49387
0 49389 5 1 1 49388
0 49390 7 1 2 49383 49389
0 49391 7 1 2 49379 49390
0 49392 7 1 2 49375 49391
0 49393 5 1 1 49392
0 49394 7 1 2 77095 49393
0 49395 5 1 1 49394
0 49396 7 1 2 86367 102039
0 49397 5 1 1 49396
0 49398 7 1 2 63647 49397
0 49399 7 1 2 49395 49398
0 49400 5 1 1 49399
0 49401 7 1 2 49365 49400
0 49402 5 1 1 49401
0 49403 7 1 2 49336 49402
0 49404 5 1 1 49403
0 49405 7 1 2 69632 49404
0 49406 5 1 1 49405
0 49407 7 1 2 74206 78019
0 49408 7 1 2 82040 93241
0 49409 7 1 2 49407 49408
0 49410 5 1 1 49409
0 49411 7 1 2 49406 49410
0 49412 5 1 1 49411
0 49413 7 1 2 61669 49412
0 49414 5 1 1 49413
0 49415 7 1 2 69850 88451
0 49416 7 1 2 97058 49415
0 49417 7 1 2 96849 49416
0 49418 5 1 1 49417
0 49419 7 1 2 49414 49418
0 49420 5 1 1 49419
0 49421 7 1 2 102757 49420
0 49422 5 1 1 49421
0 49423 7 1 2 95353 100092
0 49424 5 1 1 49423
0 49425 7 1 2 81030 75123
0 49426 5 1 1 49425
0 49427 7 1 2 78739 100573
0 49428 7 1 2 49426 49427
0 49429 5 1 1 49428
0 49430 7 1 2 49424 49429
0 49431 5 1 1 49430
0 49432 7 1 2 69851 49431
0 49433 5 1 1 49432
0 49434 7 3 2 83599 77411
0 49435 7 2 2 61406 79270
0 49436 7 2 2 63039 102780
0 49437 7 1 2 102777 102782
0 49438 5 1 1 49437
0 49439 7 1 2 49433 49438
0 49440 5 1 1 49439
0 49441 7 1 2 72194 49440
0 49442 5 1 1 49441
0 49443 7 1 2 87611 89579
0 49444 5 1 1 49443
0 49445 7 1 2 101050 49444
0 49446 5 1 1 49445
0 49447 7 1 2 89580 27091
0 49448 5 1 1 49447
0 49449 7 1 2 83215 49448
0 49450 5 1 1 49449
0 49451 7 1 2 49446 49450
0 49452 5 1 1 49451
0 49453 7 1 2 100574 49452
0 49454 5 1 1 49453
0 49455 7 1 2 71177 89576
0 49456 5 1 1 49455
0 49457 7 1 2 98291 49456
0 49458 5 1 1 49457
0 49459 7 1 2 89581 100168
0 49460 5 1 1 49459
0 49461 7 1 2 73351 100093
0 49462 7 1 2 49460 49461
0 49463 7 1 2 49458 49462
0 49464 5 1 1 49463
0 49465 7 1 2 49454 49464
0 49466 7 1 2 49442 49465
0 49467 5 1 1 49466
0 49468 7 1 2 65861 49467
0 49469 5 1 1 49468
0 49470 7 2 2 63648 75294
0 49471 7 1 2 71680 96782
0 49472 7 1 2 102784 49471
0 49473 7 1 2 102783 49472
0 49474 5 1 1 49473
0 49475 7 1 2 49469 49474
0 49476 5 1 1 49475
0 49477 7 1 2 65540 49476
0 49478 5 1 1 49477
0 49479 7 1 2 63649 101159
0 49480 5 1 1 49479
0 49481 7 1 2 90750 49480
0 49482 5 1 1 49481
0 49483 7 1 2 100575 49482
0 49484 5 1 1 49483
0 49485 7 1 2 90751 19754
0 49486 5 1 1 49485
0 49487 7 1 2 100094 49486
0 49488 5 1 1 49487
0 49489 7 1 2 49484 49488
0 49490 5 1 1 49489
0 49491 7 1 2 62220 49490
0 49492 5 1 1 49491
0 49493 7 1 2 4674 93768
0 49494 5 1 1 49493
0 49495 7 1 2 89277 90635
0 49496 5 1 1 49495
0 49497 7 2 2 49494 49496
0 49498 7 2 2 70461 102786
0 49499 7 1 2 78096 102788
0 49500 5 1 1 49499
0 49501 7 1 2 49492 49500
0 49502 5 1 1 49501
0 49503 7 1 2 64994 49502
0 49504 5 1 1 49503
0 49505 7 1 2 81056 77399
0 49506 7 1 2 102789 49505
0 49507 5 1 1 49506
0 49508 7 1 2 49504 49507
0 49509 5 1 1 49508
0 49510 7 1 2 78338 49509
0 49511 5 1 1 49510
0 49512 7 1 2 72654 101269
0 49513 7 1 2 100089 49512
0 49514 5 1 1 49513
0 49515 7 2 2 70462 79517
0 49516 5 1 1 102790
0 49517 7 1 2 100095 102791
0 49518 5 1 1 49517
0 49519 7 2 2 62909 100096
0 49520 5 1 1 102792
0 49521 7 2 2 71361 93825
0 49522 7 1 2 89270 102794
0 49523 5 1 1 49522
0 49524 7 1 2 49520 49523
0 49525 5 1 1 49524
0 49526 7 1 2 80550 49525
0 49527 5 1 1 49526
0 49528 7 1 2 49518 49527
0 49529 7 1 2 49514 49528
0 49530 5 1 1 49529
0 49531 7 1 2 80714 77096
0 49532 7 1 2 49530 49531
0 49533 5 1 1 49532
0 49534 7 1 2 49511 49533
0 49535 7 1 2 49478 49534
0 49536 5 1 1 49535
0 49537 7 1 2 69433 49536
0 49538 5 1 1 49537
0 49539 7 1 2 49422 49538
0 49540 5 1 1 49539
0 49541 7 1 2 90204 49540
0 49542 5 1 1 49541
0 49543 7 1 2 3946 38233
0 49544 5 1 1 49543
0 49545 7 1 2 76723 49544
0 49546 5 1 1 49545
0 49547 7 1 2 89502 101270
0 49548 5 1 1 49547
0 49549 7 1 2 85465 96230
0 49550 7 1 2 49548 49549
0 49551 5 1 1 49550
0 49552 7 1 2 65233 49551
0 49553 5 1 1 49552
0 49554 7 1 2 49546 49553
0 49555 5 1 1 49554
0 49556 7 1 2 81949 49555
0 49557 5 1 1 49556
0 49558 7 2 2 71362 94280
0 49559 5 1 1 102796
0 49560 7 1 2 94271 49559
0 49561 5 1 1 49560
0 49562 7 1 2 65234 49561
0 49563 5 1 1 49562
0 49564 7 1 2 84671 78318
0 49565 5 1 1 49564
0 49566 7 1 2 85950 49565
0 49567 5 3 1 49566
0 49568 7 1 2 94431 102798
0 49569 5 1 1 49568
0 49570 7 1 2 72195 91151
0 49571 5 1 1 49570
0 49572 7 1 2 49569 49571
0 49573 7 1 2 49563 49572
0 49574 5 1 1 49573
0 49575 7 1 2 86988 49574
0 49576 5 1 1 49575
0 49577 7 1 2 63650 49576
0 49578 7 1 2 49557 49577
0 49579 5 1 1 49578
0 49580 7 2 2 87367 78339
0 49581 7 2 2 79612 102801
0 49582 5 1 1 102803
0 49583 7 1 2 68488 49582
0 49584 5 1 1 49583
0 49585 7 1 2 64995 49584
0 49586 7 1 2 49579 49585
0 49587 5 1 1 49586
0 49588 7 2 2 72196 87368
0 49589 5 1 1 102805
0 49590 7 1 2 81057 97445
0 49591 7 1 2 102806 49590
0 49592 5 1 1 49591
0 49593 7 1 2 62221 49592
0 49594 7 1 2 49587 49593
0 49595 5 1 1 49594
0 49596 7 1 2 81950 94802
0 49597 5 1 1 49596
0 49598 7 1 2 86989 94949
0 49599 5 1 1 49598
0 49600 7 1 2 49597 49599
0 49601 5 1 1 49600
0 49602 7 1 2 72197 49601
0 49603 5 1 1 49602
0 49604 7 1 2 78117 93275
0 49605 5 1 1 49604
0 49606 7 1 2 49603 49605
0 49607 5 1 1 49606
0 49608 7 1 2 76724 49607
0 49609 5 1 1 49608
0 49610 7 1 2 81058 78340
0 49611 7 1 2 99176 49610
0 49612 5 1 1 49611
0 49613 7 1 2 49609 49612
0 49614 5 1 1 49613
0 49615 7 1 2 69852 49614
0 49616 5 1 1 49615
0 49617 7 1 2 77412 102804
0 49618 5 1 1 49617
0 49619 7 1 2 67059 49618
0 49620 7 1 2 49616 49619
0 49621 5 1 1 49620
0 49622 7 1 2 49595 49621
0 49623 5 1 1 49622
0 49624 7 1 2 78421 86662
0 49625 7 1 2 87387 49624
0 49626 7 1 2 100478 49625
0 49627 5 1 1 49626
0 49628 7 1 2 49623 49627
0 49629 5 1 1 49628
0 49630 7 1 2 69434 49629
0 49631 5 1 1 49630
0 49632 7 1 2 75862 77137
0 49633 7 1 2 95971 100174
0 49634 7 1 2 49632 49633
0 49635 5 1 1 49634
0 49636 7 1 2 49631 49635
0 49637 5 1 1 49636
0 49638 7 1 2 98418 49637
0 49639 5 1 1 49638
0 49640 7 1 2 64394 49639
0 49641 7 1 2 72583 87073
0 49642 7 1 2 84167 49641
0 49643 5 1 1 49642
0 49644 7 1 2 77132 86046
0 49645 7 1 2 75376 49644
0 49646 7 1 2 98236 49645
0 49647 5 1 1 49646
0 49648 7 1 2 49643 49647
0 49649 5 1 1 49648
0 49650 7 1 2 62222 49649
0 49651 5 1 1 49650
0 49652 7 1 2 74642 78829
0 49653 5 2 1 49652
0 49654 7 1 2 65541 41064
0 49655 5 1 1 49654
0 49656 7 1 2 84672 72859
0 49657 5 1 1 49656
0 49658 7 1 2 49655 49657
0 49659 5 1 1 49658
0 49660 7 1 2 65235 49659
0 49661 5 1 1 49660
0 49662 7 1 2 81033 77351
0 49663 5 1 1 49662
0 49664 7 1 2 49661 49663
0 49665 5 1 1 49664
0 49666 7 1 2 68489 49665
0 49667 5 1 1 49666
0 49668 7 1 2 102807 49667
0 49669 5 1 1 49668
0 49670 7 1 2 69633 49669
0 49671 5 1 1 49670
0 49672 7 1 2 49651 49671
0 49673 5 1 1 49672
0 49674 7 1 2 66559 49673
0 49675 5 1 1 49674
0 49676 7 1 2 87022 94458
0 49677 5 1 1 49676
0 49678 7 1 2 72584 98280
0 49679 5 1 1 49678
0 49680 7 1 2 102769 49679
0 49681 5 1 1 49680
0 49682 7 1 2 65542 49681
0 49683 5 1 1 49682
0 49684 7 1 2 94447 94432
0 49685 5 1 1 49684
0 49686 7 1 2 102766 49685
0 49687 7 1 2 49683 49686
0 49688 5 1 1 49687
0 49689 7 1 2 65236 49688
0 49690 5 1 1 49689
0 49691 7 1 2 49677 49690
0 49692 5 1 1 49691
0 49693 7 1 2 68490 49692
0 49694 5 1 1 49693
0 49695 7 1 2 49694 102808
0 49696 5 1 1 49695
0 49697 7 1 2 86990 49696
0 49698 5 1 1 49697
0 49699 7 1 2 69853 49698
0 49700 7 1 2 49675 49699
0 49701 5 1 1 49700
0 49702 7 2 2 82676 99492
0 49703 7 4 2 98402 102809
0 49704 7 1 2 80551 96041
0 49705 5 1 1 49704
0 49706 7 1 2 88236 79518
0 49707 5 1 1 49706
0 49708 7 1 2 49705 49707
0 49709 5 1 1 49708
0 49710 7 1 2 65237 49709
0 49711 5 1 1 49710
0 49712 7 1 2 87990 102672
0 49713 5 1 1 49712
0 49714 7 1 2 86991 49713
0 49715 5 1 1 49714
0 49716 7 1 2 86690 49715
0 49717 5 1 1 49716
0 49718 7 1 2 71363 96042
0 49719 7 1 2 49717 49718
0 49720 5 1 1 49719
0 49721 7 1 2 81951 86911
0 49722 5 1 1 49721
0 49723 7 1 2 70961 95685
0 49724 5 1 1 49723
0 49725 7 1 2 49722 49724
0 49726 5 1 1 49725
0 49727 7 1 2 69052 73352
0 49728 7 1 2 49726 49727
0 49729 5 1 1 49728
0 49730 7 1 2 49720 49729
0 49731 5 1 1 49730
0 49732 7 1 2 65543 49731
0 49733 5 1 1 49732
0 49734 7 1 2 49711 49733
0 49735 5 1 1 49734
0 49736 7 1 2 75788 49735
0 49737 5 1 1 49736
0 49738 7 1 2 79271 91554
0 49739 5 1 1 49738
0 49740 7 2 2 70152 87369
0 49741 7 1 2 75169 102815
0 49742 5 1 1 49741
0 49743 7 1 2 49739 49742
0 49744 5 1 1 49743
0 49745 7 1 2 70463 49744
0 49746 5 1 1 49745
0 49747 7 1 2 102776 47535
0 49748 5 1 1 49747
0 49749 7 1 2 81952 49748
0 49750 5 1 1 49749
0 49751 7 4 2 86992 73936
0 49752 5 1 1 102817
0 49753 7 1 2 65238 102818
0 49754 5 1 1 49753
0 49755 7 1 2 49750 49754
0 49756 5 1 1 49755
0 49757 7 1 2 75789 49756
0 49758 5 1 1 49757
0 49759 7 1 2 49746 49758
0 49760 5 1 1 49759
0 49761 7 1 2 72655 49760
0 49762 5 1 1 49761
0 49763 7 1 2 102752 102816
0 49764 5 1 1 49763
0 49765 7 1 2 64996 49764
0 49766 7 1 2 49762 49765
0 49767 7 1 2 49737 49766
0 49768 5 1 1 49767
0 49769 7 1 2 102811 49768
0 49770 7 1 2 49701 49769
0 49771 5 1 1 49770
0 49772 7 6 2 75002 77533
0 49773 7 1 2 101668 102821
0 49774 5 1 1 49773
0 49775 7 1 2 100078 100413
0 49776 5 1 1 49775
0 49777 7 1 2 49774 49776
0 49778 5 1 1 49777
0 49779 7 1 2 61407 49778
0 49780 5 1 1 49779
0 49781 7 1 2 99028 99412
0 49782 7 1 2 102822 49781
0 49783 5 1 1 49782
0 49784 7 1 2 49780 49783
0 49785 5 1 1 49784
0 49786 7 1 2 69435 49785
0 49787 5 1 1 49786
0 49788 7 3 2 63040 99206
0 49789 7 6 2 79380 102827
0 49790 7 1 2 72656 102830
0 49791 5 1 1 49790
0 49792 7 1 2 49787 49791
0 49793 5 1 1 49792
0 49794 7 1 2 65862 49793
0 49795 5 1 1 49794
0 49796 7 1 2 102642 102831
0 49797 5 1 1 49796
0 49798 7 1 2 49795 49797
0 49799 5 1 1 49798
0 49800 7 1 2 76908 49799
0 49801 5 1 1 49800
0 49802 7 1 2 77337 99276
0 49803 7 2 2 101772 49802
0 49804 7 1 2 73856 102663
0 49805 7 1 2 102836 49804
0 49806 5 1 1 49805
0 49807 7 1 2 49801 49806
0 49808 5 1 1 49807
0 49809 7 1 2 73353 49808
0 49810 5 1 1 49809
0 49811 7 1 2 76278 102832
0 49812 7 1 2 97144 49811
0 49813 5 1 1 49812
0 49814 7 1 2 49810 49813
0 49815 5 1 1 49814
0 49816 7 1 2 90205 49815
0 49817 5 1 1 49816
0 49818 7 4 2 69436 98419
0 49819 7 1 2 93279 94513
0 49820 5 1 1 49819
0 49821 7 1 2 81953 102823
0 49822 5 1 1 49821
0 49823 7 1 2 98319 102677
0 49824 5 1 1 49823
0 49825 7 1 2 49822 49824
0 49826 5 1 1 49825
0 49827 7 1 2 91152 49826
0 49828 5 1 1 49827
0 49829 7 1 2 49820 49828
0 49830 5 1 1 49829
0 49831 7 1 2 102838 49830
0 49832 5 1 1 49831
0 49833 7 3 2 87370 102812
0 49834 7 1 2 70153 102710
0 49835 5 1 1 49834
0 49836 7 1 2 94969 49835
0 49837 5 1 1 49836
0 49838 7 1 2 102842 49837
0 49839 5 1 1 49838
0 49840 7 1 2 49832 49839
0 49841 5 1 1 49840
0 49842 7 1 2 73354 49841
0 49843 5 1 1 49842
0 49844 7 1 2 85830 92152
0 49845 7 1 2 102813 49844
0 49846 7 1 2 102616 49845
0 49847 5 1 1 49846
0 49848 7 1 2 64997 49847
0 49849 7 1 2 49843 49848
0 49850 7 1 2 49817 49849
0 49851 5 1 1 49850
0 49852 7 1 2 78894 100519
0 49853 5 1 1 49852
0 49854 7 1 2 42553 49853
0 49855 5 1 1 49854
0 49856 7 1 2 61670 49855
0 49857 5 1 1 49856
0 49858 7 1 2 101697 99975
0 49859 5 1 1 49858
0 49860 7 1 2 49857 49859
0 49861 5 1 1 49860
0 49862 7 1 2 61408 49861
0 49863 5 1 1 49862
0 49864 7 2 2 66299 87483
0 49865 7 1 2 94826 99831
0 49866 7 1 2 102845 49865
0 49867 5 1 1 49866
0 49868 7 1 2 49863 49867
0 49869 5 1 1 49868
0 49870 7 1 2 102062 49869
0 49871 5 1 1 49870
0 49872 7 1 2 71178 88197
0 49873 5 1 1 49872
0 49874 7 1 2 77261 95828
0 49875 5 1 1 49874
0 49876 7 1 2 49873 49875
0 49877 5 1 1 49876
0 49878 7 2 2 83160 102758
0 49879 7 1 2 49877 102847
0 49880 5 1 1 49879
0 49881 7 1 2 49871 49880
0 49882 5 1 1 49881
0 49883 7 1 2 65863 49882
0 49884 5 1 1 49883
0 49885 7 1 2 70762 96476
0 49886 5 1 1 49885
0 49887 7 1 2 17705 49886
0 49888 5 1 1 49887
0 49889 7 1 2 72585 102848
0 49890 7 1 2 49888 49889
0 49891 5 1 1 49890
0 49892 7 1 2 49884 49891
0 49893 5 1 1 49892
0 49894 7 1 2 76909 49893
0 49895 5 1 1 49894
0 49896 7 3 2 83161 91946
0 49897 7 2 2 70962 102849
0 49898 7 1 2 87500 102837
0 49899 7 1 2 102852 49898
0 49900 5 1 1 49899
0 49901 7 1 2 49895 49900
0 49902 5 1 1 49901
0 49903 7 1 2 73355 49902
0 49904 5 1 1 49903
0 49905 7 1 2 101770 102617
0 49906 7 1 2 99681 49905
0 49907 5 1 1 49906
0 49908 7 1 2 69854 49907
0 49909 7 1 2 49904 49908
0 49910 5 1 1 49909
0 49911 7 1 2 74385 49910
0 49912 7 1 2 49851 49911
0 49913 5 1 1 49912
0 49914 7 1 2 49771 49913
0 49915 7 1 2 49640 49914
0 49916 7 1 2 49542 49915
0 49917 7 1 2 49328 49916
0 49918 5 1 1 49917
0 49919 7 2 2 70464 90636
0 49920 7 1 2 63205 101329
0 49921 5 1 1 49920
0 49922 7 1 2 95231 49921
0 49923 5 1 1 49922
0 49924 7 1 2 71600 49923
0 49925 5 1 1 49924
0 49926 7 1 2 92091 101201
0 49927 5 1 1 49926
0 49928 7 1 2 73267 92438
0 49929 5 1 1 49928
0 49930 7 2 2 906 49929
0 49931 7 1 2 78937 102856
0 49932 5 1 1 49931
0 49933 7 1 2 49927 49932
0 49934 7 1 2 49925 49933
0 49935 5 1 1 49934
0 49936 7 1 2 66560 49935
0 49937 5 1 1 49936
0 49938 7 1 2 71601 101321
0 49939 5 1 1 49938
0 49940 7 1 2 72434 49939
0 49941 5 1 1 49940
0 49942 7 1 2 89089 49941
0 49943 5 1 1 49942
0 49944 7 1 2 49937 49943
0 49945 5 1 1 49944
0 49946 7 1 2 69437 49945
0 49947 5 1 1 49946
0 49948 7 1 2 96899 100427
0 49949 5 1 1 49948
0 49950 7 1 2 49947 49949
0 49951 5 1 1 49950
0 49952 7 1 2 90681 49951
0 49953 5 1 1 49952
0 49954 7 1 2 78938 85591
0 49955 5 1 1 49954
0 49956 7 1 2 78895 95715
0 49957 5 1 1 49956
0 49958 7 1 2 66561 49957
0 49959 7 1 2 49955 49958
0 49960 5 1 1 49959
0 49961 7 1 2 61671 27399
0 49962 5 1 1 49961
0 49963 7 1 2 64582 90692
0 49964 7 1 2 49962 49963
0 49965 7 1 2 49960 49964
0 49966 5 1 1 49965
0 49967 7 1 2 49953 49966
0 49968 5 1 1 49967
0 49969 7 1 2 102854 49968
0 49970 5 1 1 49969
0 49971 7 1 2 66562 89068
0 49972 5 1 1 49971
0 49973 7 1 2 4290 49972
0 49974 5 1 1 49973
0 49975 7 3 2 87218 100289
0 49976 7 1 2 102601 102858
0 49977 7 1 2 49974 49976
0 49978 5 1 1 49977
0 49979 7 1 2 49970 49978
0 49980 5 1 1 49979
0 49981 7 1 2 68491 49980
0 49982 5 1 1 49981
0 49983 7 2 2 89523 101947
0 49984 5 1 1 102861
0 49985 7 1 2 81269 84696
0 49986 7 1 2 102862 49985
0 49987 5 1 1 49986
0 49988 7 1 2 49982 49987
0 49989 5 1 1 49988
0 49990 7 1 2 84489 49989
0 49991 5 1 1 49990
0 49992 7 1 2 71364 86807
0 49993 5 1 1 49992
0 49994 7 1 2 94779 49993
0 49995 5 2 1 49994
0 49996 7 1 2 99661 102863
0 49997 5 1 1 49996
0 49998 7 1 2 63041 96900
0 49999 5 1 1 49998
0 50000 7 1 2 49997 49999
0 50001 5 1 1 50000
0 50002 7 1 2 87347 50001
0 50003 5 1 1 50002
0 50004 7 1 2 82384 99109
0 50005 7 1 2 96901 50004
0 50006 5 1 1 50005
0 50007 7 1 2 50003 50006
0 50008 5 1 1 50007
0 50009 7 1 2 66300 50008
0 50010 5 1 1 50009
0 50011 7 1 2 93057 101766
0 50012 7 1 2 85592 50011
0 50013 5 1 1 50012
0 50014 7 1 2 50010 50013
0 50015 5 1 1 50014
0 50016 7 1 2 70465 50015
0 50017 5 1 1 50016
0 50018 7 1 2 93068 102859
0 50019 7 1 2 101235 50018
0 50020 5 1 1 50019
0 50021 7 1 2 50017 50020
0 50022 5 1 1 50021
0 50023 7 1 2 78963 50022
0 50024 5 1 1 50023
0 50025 7 1 2 84094 102864
0 50026 5 1 1 50025
0 50027 7 1 2 81492 85593
0 50028 5 1 1 50027
0 50029 7 1 2 50026 50028
0 50030 5 1 1 50029
0 50031 7 1 2 90682 50030
0 50032 5 1 1 50031
0 50033 7 1 2 78972 90693
0 50034 7 1 2 96902 50033
0 50035 5 1 1 50034
0 50036 7 1 2 50032 50035
0 50037 5 1 1 50036
0 50038 7 1 2 102855 50037
0 50039 5 1 1 50038
0 50040 7 1 2 67900 89671
0 50041 7 1 2 80153 50040
0 50042 7 1 2 87219 101524
0 50043 7 1 2 50041 50042
0 50044 5 1 1 50043
0 50045 7 1 2 50039 50044
0 50046 5 1 1 50045
0 50047 7 1 2 87705 50046
0 50048 5 1 1 50047
0 50049 7 1 2 50024 50048
0 50050 5 1 1 50049
0 50051 7 1 2 75057 50050
0 50052 5 1 1 50051
0 50053 7 1 2 67060 50052
0 50054 7 1 2 49991 50053
0 50055 5 1 1 50054
0 50056 7 1 2 8473 49752
0 50057 5 1 1 50056
0 50058 7 1 2 72657 50057
0 50059 5 1 1 50058
0 50060 7 2 2 71745 81954
0 50061 5 1 1 102865
0 50062 7 1 2 50059 50061
0 50063 5 1 1 50062
0 50064 7 2 2 64583 50063
0 50065 7 1 2 98387 102867
0 50066 5 1 1 50065
0 50067 7 1 2 20230 95689
0 50068 5 1 1 50067
0 50069 7 1 2 64194 50068
0 50070 5 1 1 50069
0 50071 7 1 2 78453 102105
0 50072 5 1 1 50071
0 50073 7 1 2 50070 50072
0 50074 5 1 1 50073
0 50075 7 1 2 99662 50074
0 50076 5 1 1 50075
0 50077 7 1 2 230 101722
0 50078 5 1 1 50077
0 50079 7 1 2 50076 50078
0 50080 5 1 1 50079
0 50081 7 1 2 70466 50080
0 50082 5 1 1 50081
0 50083 7 2 2 86800 99663
0 50084 5 1 1 102869
0 50085 7 1 2 50084 100284
0 50086 5 1 1 50085
0 50087 7 1 2 102819 50086
0 50088 5 1 1 50087
0 50089 7 1 2 50082 50088
0 50090 5 1 1 50089
0 50091 7 1 2 91258 50090
0 50092 5 1 1 50091
0 50093 7 1 2 50066 50092
0 50094 5 1 1 50093
0 50095 7 1 2 66301 50094
0 50096 5 1 1 50095
0 50097 7 2 2 84413 101948
0 50098 7 1 2 101101 102871
0 50099 5 1 1 50098
0 50100 7 1 2 87336 48734
0 50101 5 1 1 50100
0 50102 7 1 2 64195 50101
0 50103 5 2 1 50102
0 50104 7 1 2 87337 29917
0 50105 5 2 1 50104
0 50106 7 1 2 27343 102875
0 50107 5 1 1 50106
0 50108 7 1 2 102873 50107
0 50109 5 1 1 50108
0 50110 7 1 2 70467 50109
0 50111 5 1 1 50110
0 50112 7 1 2 87338 14893
0 50113 5 1 1 50112
0 50114 7 1 2 79395 50113
0 50115 5 1 1 50114
0 50116 7 1 2 50111 50115
0 50117 5 1 1 50116
0 50118 7 1 2 90683 50117
0 50119 5 1 1 50118
0 50120 7 1 2 50099 50119
0 50121 5 1 1 50120
0 50122 7 1 2 90206 50121
0 50123 5 1 1 50122
0 50124 7 1 2 98559 102868
0 50125 5 1 1 50124
0 50126 7 2 2 70468 98320
0 50127 7 2 2 91259 100204
0 50128 7 1 2 102877 102879
0 50129 5 1 1 50128
0 50130 7 1 2 64584 80552
0 50131 7 1 2 98564 50130
0 50132 5 1 1 50131
0 50133 7 1 2 50129 50132
0 50134 5 1 1 50133
0 50135 7 1 2 96043 50134
0 50136 5 1 1 50135
0 50137 7 1 2 50125 50136
0 50138 7 1 2 50123 50137
0 50139 7 1 2 50096 50138
0 50140 5 1 1 50139
0 50141 7 1 2 71365 50140
0 50142 5 1 1 50141
0 50143 7 1 2 87220 92362
0 50144 5 2 1 50143
0 50145 7 1 2 70963 95940
0 50146 5 1 1 50145
0 50147 7 1 2 76602 50146
0 50148 5 1 1 50147
0 50149 7 2 2 64804 50148
0 50150 7 1 2 61672 102883
0 50151 5 1 1 50150
0 50152 7 1 2 102881 50151
0 50153 5 1 1 50152
0 50154 7 1 2 99664 50153
0 50155 5 1 1 50154
0 50156 7 1 2 91755 101698
0 50157 5 1 1 50156
0 50158 7 1 2 50155 50157
0 50159 5 1 1 50158
0 50160 7 1 2 91260 50159
0 50161 5 1 1 50160
0 50162 7 1 2 87501 87697
0 50163 7 1 2 101378 50162
0 50164 5 1 1 50163
0 50165 7 1 2 50161 50164
0 50166 5 1 1 50165
0 50167 7 1 2 66302 50166
0 50168 5 1 1 50167
0 50169 7 2 2 81955 99524
0 50170 5 1 1 102885
0 50171 7 1 2 98557 102886
0 50172 5 1 1 50171
0 50173 7 1 2 50168 50172
0 50174 5 1 1 50173
0 50175 7 1 2 73356 50174
0 50176 5 1 1 50175
0 50177 7 2 2 100275 98397
0 50178 5 1 1 102887
0 50179 7 3 2 67901 69053
0 50180 7 2 2 91647 102889
0 50181 5 1 1 102892
0 50182 7 1 2 91261 102893
0 50183 5 1 1 50182
0 50184 7 1 2 50178 50183
0 50185 5 1 1 50184
0 50186 7 1 2 62910 50185
0 50187 5 1 1 50186
0 50188 7 1 2 86313 86457
0 50189 7 1 2 102438 50188
0 50190 5 1 1 50189
0 50191 7 1 2 50187 50190
0 50192 5 1 1 50191
0 50193 7 1 2 86993 50192
0 50194 5 1 1 50193
0 50195 7 1 2 90560 102888
0 50196 5 1 1 50195
0 50197 7 1 2 50194 50196
0 50198 5 1 1 50197
0 50199 7 1 2 66303 50198
0 50200 5 1 1 50199
0 50201 7 1 2 100546 50181
0 50202 5 1 1 50201
0 50203 7 1 2 66304 50202
0 50204 5 1 1 50203
0 50205 7 1 2 50204 100544
0 50206 5 1 1 50205
0 50207 7 1 2 84414 50206
0 50208 5 1 1 50207
0 50209 7 1 2 67902 99029
0 50210 7 1 2 92282 50209
0 50211 5 1 1 50210
0 50212 7 1 2 50208 50211
0 50213 5 1 1 50212
0 50214 7 1 2 75553 50213
0 50215 5 1 1 50214
0 50216 7 1 2 73780 90684
0 50217 7 1 2 102659 50216
0 50218 5 1 1 50217
0 50219 7 1 2 64196 101669
0 50220 5 1 1 50219
0 50221 7 1 2 100083 50220
0 50222 5 1 1 50221
0 50223 7 1 2 66305 50222
0 50224 5 1 1 50223
0 50225 7 1 2 101741 50224
0 50226 5 1 1 50225
0 50227 7 1 2 64585 87984
0 50228 7 1 2 50226 50227
0 50229 5 1 1 50228
0 50230 7 1 2 50218 50229
0 50231 7 1 2 50215 50230
0 50232 5 1 1 50231
0 50233 7 1 2 90207 50232
0 50234 5 1 1 50233
0 50235 7 2 2 64586 78341
0 50236 7 1 2 98565 102894
0 50237 5 1 1 50236
0 50238 7 5 2 70763 98321
0 50239 7 1 2 102880 102896
0 50240 5 1 1 50239
0 50241 7 1 2 50237 50240
0 50242 5 1 1 50241
0 50243 7 1 2 96044 50242
0 50244 5 1 1 50243
0 50245 7 1 2 90563 102681
0 50246 5 1 1 50245
0 50247 7 1 2 100276 98560
0 50248 7 1 2 50246 50247
0 50249 5 1 1 50248
0 50250 7 1 2 50244 50249
0 50251 7 1 2 50234 50250
0 50252 7 1 2 50200 50251
0 50253 5 1 1 50252
0 50254 7 1 2 84608 50253
0 50255 5 1 1 50254
0 50256 7 1 2 82121 102884
0 50257 5 1 1 50256
0 50258 7 1 2 34927 50257
0 50259 5 1 1 50258
0 50260 7 1 2 91363 102597
0 50261 7 1 2 90208 50260
0 50262 7 1 2 50259 50261
0 50263 5 1 1 50262
0 50264 7 1 2 50255 50263
0 50265 7 1 2 50176 50264
0 50266 7 1 2 50142 50265
0 50267 5 1 1 50266
0 50268 7 1 2 77413 50267
0 50269 5 1 1 50268
0 50270 7 1 2 101917 102737
0 50271 5 1 1 50270
0 50272 7 1 2 83524 101755
0 50273 5 1 1 50272
0 50274 7 1 2 50271 50273
0 50275 5 1 1 50274
0 50276 7 1 2 71366 19235
0 50277 5 1 1 50276
0 50278 7 1 2 84609 85308
0 50279 5 1 1 50278
0 50280 7 1 2 86557 50279
0 50281 7 1 2 50277 50280
0 50282 5 1 1 50281
0 50283 7 1 2 50275 50282
0 50284 5 1 1 50283
0 50285 7 1 2 78482 84168
0 50286 7 1 2 76352 50285
0 50287 7 1 2 99388 50286
0 50288 5 1 1 50287
0 50289 7 1 2 50284 50288
0 50290 5 1 1 50289
0 50291 7 1 2 64587 50290
0 50292 5 1 1 50291
0 50293 7 1 2 77844 100419
0 50294 5 1 1 50293
0 50295 7 1 2 71367 50294
0 50296 5 1 1 50295
0 50297 7 1 2 62911 102897
0 50298 5 1 1 50297
0 50299 7 1 2 50296 50298
0 50300 5 1 1 50299
0 50301 7 1 2 70469 50300
0 50302 5 1 1 50301
0 50303 7 1 2 86496 100420
0 50304 5 1 1 50303
0 50305 7 1 2 87952 50304
0 50306 5 1 1 50305
0 50307 7 1 2 50302 50306
0 50308 5 1 1 50307
0 50309 7 1 2 101876 102096
0 50310 7 1 2 50308 50309
0 50311 5 1 1 50310
0 50312 7 1 2 50292 50311
0 50313 5 1 1 50312
0 50314 7 1 2 83162 50313
0 50315 5 1 1 50314
0 50316 7 1 2 76008 74927
0 50317 7 1 2 79928 99598
0 50318 7 1 2 50316 50317
0 50319 5 1 1 50318
0 50320 7 1 2 69855 84085
0 50321 7 1 2 99630 50320
0 50322 7 1 2 101425 50321
0 50323 5 1 1 50322
0 50324 7 1 2 50319 50323
0 50325 5 1 1 50324
0 50326 7 1 2 66563 50325
0 50327 5 1 1 50326
0 50328 7 1 2 80632 82291
0 50329 7 1 2 92559 50328
0 50330 7 1 2 84267 50329
0 50331 5 1 1 50330
0 50332 7 1 2 50327 50331
0 50333 5 1 1 50332
0 50334 7 1 2 94694 50333
0 50335 5 1 1 50334
0 50336 7 1 2 81956 89429
0 50337 7 1 2 98489 50336
0 50338 7 1 2 101426 50337
0 50339 5 1 1 50338
0 50340 7 1 2 50335 50339
0 50341 5 1 1 50340
0 50342 7 1 2 66306 50341
0 50343 5 1 1 50342
0 50344 7 1 2 74942 93754
0 50345 7 1 2 102142 50344
0 50346 7 1 2 92107 50345
0 50347 5 1 1 50346
0 50348 7 1 2 50343 50347
0 50349 5 1 1 50348
0 50350 7 1 2 72198 50349
0 50351 5 1 1 50350
0 50352 7 1 2 62223 50351
0 50353 7 1 2 50315 50352
0 50354 7 1 2 50269 50353
0 50355 5 1 1 50354
0 50356 7 1 2 65239 50355
0 50357 7 1 2 50055 50356
0 50358 5 1 1 50357
0 50359 7 1 2 101322 99892
0 50360 5 1 1 50359
0 50361 7 2 2 84128 71069
0 50362 7 1 2 100277 102901
0 50363 5 1 1 50362
0 50364 7 1 2 50360 50363
0 50365 5 1 1 50364
0 50366 7 1 2 68045 50365
0 50367 5 1 1 50366
0 50368 7 1 2 64805 101764
0 50369 5 1 1 50368
0 50370 7 1 2 68242 79105
0 50371 5 1 1 50370
0 50372 7 1 2 50369 50371
0 50373 5 2 1 50372
0 50374 7 1 2 63206 100278
0 50375 7 1 2 102903 50374
0 50376 5 1 1 50375
0 50377 7 1 2 50367 50376
0 50378 5 1 1 50377
0 50379 7 1 2 71602 50378
0 50380 5 1 1 50379
0 50381 7 2 2 69054 78483
0 50382 7 1 2 102086 102905
0 50383 5 1 1 50382
0 50384 7 1 2 78896 101532
0 50385 5 1 1 50384
0 50386 7 1 2 78939 95855
0 50387 5 1 1 50386
0 50388 7 1 2 50385 50387
0 50389 5 1 1 50388
0 50390 7 1 2 61914 50389
0 50391 5 1 1 50390
0 50392 7 1 2 81391 76676
0 50393 5 2 1 50392
0 50394 7 1 2 84129 96658
0 50395 5 1 1 50394
0 50396 7 1 2 102907 50395
0 50397 7 1 2 50391 50396
0 50398 5 1 1 50397
0 50399 7 1 2 64588 50398
0 50400 5 1 1 50399
0 50401 7 1 2 50383 50400
0 50402 5 1 1 50401
0 50403 7 1 2 73223 50402
0 50404 5 1 1 50403
0 50405 7 1 2 61673 50404
0 50406 7 1 2 50380 50405
0 50407 5 1 1 50406
0 50408 7 1 2 97187 101323
0 50409 5 1 1 50408
0 50410 7 1 2 68046 95227
0 50411 7 1 2 87311 50410
0 50412 5 1 1 50411
0 50413 7 1 2 50409 50412
0 50414 5 1 1 50413
0 50415 7 1 2 64806 50414
0 50416 5 1 1 50415
0 50417 7 1 2 95675 97364
0 50418 5 1 1 50417
0 50419 7 1 2 50416 50418
0 50420 5 1 1 50419
0 50421 7 1 2 71603 50420
0 50422 5 1 1 50421
0 50423 7 1 2 101761 102857
0 50424 5 1 1 50423
0 50425 7 2 2 74975 80172
0 50426 7 1 2 90493 102909
0 50427 5 1 1 50426
0 50428 7 1 2 50424 50427
0 50429 5 1 1 50428
0 50430 7 1 2 68047 50429
0 50431 5 1 1 50430
0 50432 7 1 2 76677 90796
0 50433 7 1 2 102910 50432
0 50434 5 1 1 50433
0 50435 7 1 2 50431 50434
0 50436 7 1 2 50422 50435
0 50437 5 1 1 50436
0 50438 7 1 2 69438 50437
0 50439 5 1 1 50438
0 50440 7 1 2 87312 101324
0 50441 5 1 1 50440
0 50442 7 1 2 72658 88987
0 50443 5 1 1 50442
0 50444 7 1 2 50441 50443
0 50445 5 1 1 50444
0 50446 7 1 2 71604 50445
0 50447 5 1 1 50446
0 50448 7 1 2 73224 96017
0 50449 5 1 1 50448
0 50450 7 1 2 50447 50449
0 50451 5 1 1 50450
0 50452 7 1 2 81493 50451
0 50453 5 1 1 50452
0 50454 7 1 2 66564 50453
0 50455 7 1 2 50439 50454
0 50456 5 1 1 50455
0 50457 7 1 2 66307 50456
0 50458 7 1 2 50407 50457
0 50459 5 1 1 50458
0 50460 7 1 2 93769 50459
0 50461 5 1 1 50460
0 50462 7 1 2 68048 102904
0 50463 5 1 1 50462
0 50464 7 1 2 78484 92265
0 50465 5 1 1 50464
0 50466 7 1 2 50463 50465
0 50467 5 1 1 50466
0 50468 7 1 2 66565 50467
0 50469 5 1 1 50468
0 50470 7 1 2 83389 87259
0 50471 5 1 1 50470
0 50472 7 1 2 50469 50471
0 50473 5 1 1 50472
0 50474 7 1 2 96903 50473
0 50475 5 1 1 50474
0 50476 7 1 2 90694 50475
0 50477 5 1 1 50476
0 50478 7 1 2 70470 50477
0 50479 7 1 2 50461 50478
0 50480 5 1 1 50479
0 50481 7 1 2 76193 99893
0 50482 5 1 1 50481
0 50483 7 1 2 90521 50482
0 50484 5 1 1 50483
0 50485 7 1 2 62912 50484
0 50486 5 1 1 50485
0 50487 7 1 2 91903 101762
0 50488 5 1 1 50487
0 50489 7 1 2 50486 50488
0 50490 5 1 1 50489
0 50491 7 1 2 102598 102860
0 50492 7 1 2 50490 50491
0 50493 5 1 1 50492
0 50494 7 1 2 50480 50493
0 50495 5 1 1 50494
0 50496 7 1 2 75170 50495
0 50497 5 1 1 50496
0 50498 7 1 2 95471 99389
0 50499 5 1 1 50498
0 50500 7 1 2 97224 101444
0 50501 5 1 1 50500
0 50502 7 1 2 50499 50501
0 50503 5 1 1 50502
0 50504 7 1 2 82175 97195
0 50505 7 1 2 84387 50504
0 50506 7 1 2 50503 50505
0 50507 5 1 1 50506
0 50508 7 1 2 50497 50507
0 50509 5 1 1 50508
0 50510 7 1 2 70154 50509
0 50511 5 1 1 50510
0 50512 7 1 2 69251 50511
0 50513 7 1 2 50358 50512
0 50514 5 1 1 50513
0 50515 7 1 2 49918 50514
0 50516 5 1 1 50515
0 50517 7 1 2 96951 50516
0 50518 5 1 1 50517
0 50519 7 1 2 98322 100090
0 50520 5 1 1 50519
0 50521 7 1 2 71179 100097
0 50522 5 1 1 50521
0 50523 7 1 2 50520 50522
0 50524 5 1 1 50523
0 50525 7 1 2 69439 50524
0 50526 5 1 1 50525
0 50527 7 1 2 84673 102833
0 50528 5 1 1 50527
0 50529 7 1 2 50526 50528
0 50530 5 1 1 50529
0 50531 7 1 2 62662 50530
0 50532 5 1 1 50531
0 50533 7 1 2 102828 100925
0 50534 5 1 1 50533
0 50535 7 1 2 50532 50534
0 50536 5 1 1 50535
0 50537 7 1 2 90209 50536
0 50538 5 1 1 50537
0 50539 7 1 2 102694 102839
0 50540 5 1 1 50539
0 50541 7 1 2 66566 84664
0 50542 5 1 1 50541
0 50543 7 1 2 102843 50542
0 50544 5 1 1 50543
0 50545 7 1 2 50540 50544
0 50546 5 1 1 50545
0 50547 7 1 2 62663 50546
0 50548 5 1 1 50547
0 50549 7 1 2 72804 93219
0 50550 5 1 1 50549
0 50551 7 1 2 23616 50550
0 50552 5 1 1 50551
0 50553 7 1 2 102814 50552
0 50554 5 1 1 50553
0 50555 7 1 2 64998 50554
0 50556 7 1 2 50548 50555
0 50557 7 1 2 50538 50556
0 50558 5 1 1 50557
0 50559 7 2 2 69440 98323
0 50560 7 1 2 93826 102911
0 50561 5 1 1 50560
0 50562 7 1 2 49330 50561
0 50563 5 1 1 50562
0 50564 7 1 2 91947 50563
0 50565 5 1 1 50564
0 50566 7 2 2 100079 100628
0 50567 5 1 1 102913
0 50568 7 1 2 102912 102914
0 50569 5 1 1 50568
0 50570 7 1 2 50565 50569
0 50571 5 1 1 50570
0 50572 7 1 2 87026 50571
0 50573 5 1 1 50572
0 50574 7 2 2 90624 100279
0 50575 7 1 2 102850 102915
0 50576 5 1 1 50575
0 50577 7 1 2 50573 50576
0 50578 5 1 1 50577
0 50579 7 1 2 62664 50578
0 50580 5 1 1 50579
0 50581 7 2 2 72805 102759
0 50582 7 1 2 102917 102853
0 50583 5 1 1 50582
0 50584 7 1 2 69856 50583
0 50585 7 1 2 50580 50584
0 50586 5 1 1 50585
0 50587 7 1 2 86509 50586
0 50588 7 1 2 50558 50587
0 50589 5 1 1 50588
0 50590 7 1 2 91720 97022
0 50591 5 1 1 50590
0 50592 7 1 2 50591 102793
0 50593 5 1 1 50592
0 50594 7 1 2 100576 102686
0 50595 5 1 1 50594
0 50596 7 1 2 50593 50595
0 50597 5 1 1 50596
0 50598 7 1 2 72080 50597
0 50599 5 1 1 50598
0 50600 7 1 2 100098 100974
0 50601 5 1 1 50600
0 50602 7 1 2 50599 50601
0 50603 5 1 1 50602
0 50604 7 1 2 69441 50603
0 50605 5 1 1 50604
0 50606 7 1 2 80385 102834
0 50607 5 1 1 50606
0 50608 7 1 2 50605 50607
0 50609 5 1 1 50608
0 50610 7 1 2 90210 50609
0 50611 5 1 1 50610
0 50612 7 1 2 87484 99464
0 50613 5 2 1 50612
0 50614 7 1 2 48866 102919
0 50615 5 1 1 50614
0 50616 7 1 2 71368 50615
0 50617 5 1 1 50616
0 50618 7 1 2 73083 81957
0 50619 5 1 1 50618
0 50620 7 1 2 34181 50619
0 50621 5 1 1 50620
0 50622 7 1 2 73357 50621
0 50623 5 1 1 50622
0 50624 7 1 2 50617 50623
0 50625 5 1 1 50624
0 50626 7 1 2 72081 50625
0 50627 5 1 1 50626
0 50628 7 1 2 93384 97905
0 50629 5 1 1 50628
0 50630 7 1 2 50627 50629
0 50631 5 1 1 50630
0 50632 7 1 2 102840 50631
0 50633 5 1 1 50632
0 50634 7 2 2 86034 90625
0 50635 7 1 2 92093 102921
0 50636 7 1 2 101225 50635
0 50637 5 1 1 50636
0 50638 7 1 2 50633 50637
0 50639 7 1 2 50611 50638
0 50640 5 1 1 50639
0 50641 7 1 2 64999 50640
0 50642 5 1 1 50641
0 50643 7 1 2 73626 102760
0 50644 5 1 1 50643
0 50645 7 1 2 86314 100775
0 50646 7 1 2 102687 50645
0 50647 5 1 1 50646
0 50648 7 1 2 50644 50647
0 50649 5 2 1 50648
0 50650 7 1 2 91948 102923
0 50651 5 1 1 50650
0 50652 7 2 2 72082 102688
0 50653 7 1 2 84095 99115
0 50654 7 1 2 102925 50653
0 50655 5 1 1 50654
0 50656 7 1 2 50651 50655
0 50657 5 1 1 50656
0 50658 7 1 2 87313 50657
0 50659 5 1 1 50658
0 50660 7 1 2 50642 50659
0 50661 7 1 2 50589 50660
0 50662 5 1 1 50661
0 50663 7 1 2 65240 50662
0 50664 5 1 1 50663
0 50665 7 1 2 71070 91323
0 50666 7 1 2 99832 50665
0 50667 7 1 2 79562 102810
0 50668 7 1 2 50666 50667
0 50669 5 1 1 50668
0 50670 7 1 2 50664 50669
0 50671 5 1 1 50670
0 50672 7 1 2 63651 50671
0 50673 5 1 1 50672
0 50674 7 1 2 78224 95402
0 50675 5 2 1 50674
0 50676 7 1 2 100300 102927
0 50677 5 1 1 50676
0 50678 7 4 2 89733 77957
0 50679 7 1 2 102761 102929
0 50680 5 1 1 50679
0 50681 7 1 2 50677 50680
0 50682 5 1 1 50681
0 50683 7 1 2 73225 50682
0 50684 5 1 1 50683
0 50685 7 3 2 71369 100737
0 50686 7 1 2 94133 102933
0 50687 7 1 2 99337 50686
0 50688 5 1 1 50687
0 50689 7 1 2 50684 50688
0 50690 5 1 1 50689
0 50691 7 1 2 88198 50690
0 50692 5 1 1 50691
0 50693 7 1 2 102926 100767
0 50694 5 1 1 50693
0 50695 7 1 2 94154 101452
0 50696 5 1 1 50695
0 50697 7 1 2 50694 50696
0 50698 5 2 1 50697
0 50699 7 1 2 64807 102936
0 50700 5 1 1 50699
0 50701 7 1 2 50692 50700
0 50702 5 1 1 50701
0 50703 7 1 2 87314 50702
0 50704 5 1 1 50703
0 50705 7 1 2 62665 102870
0 50706 5 1 1 50705
0 50707 7 1 2 49068 50706
0 50708 5 1 1 50707
0 50709 7 1 2 89271 50708
0 50710 5 1 1 50709
0 50711 7 1 2 84415 99699
0 50712 7 1 2 102930 50711
0 50713 5 1 1 50712
0 50714 7 1 2 50710 50713
0 50715 5 1 1 50714
0 50716 7 1 2 90211 50715
0 50717 5 1 1 50716
0 50718 7 1 2 88935 98779
0 50719 7 1 2 99177 50718
0 50720 5 1 1 50719
0 50721 7 1 2 86994 102931
0 50722 5 1 1 50721
0 50723 7 1 2 86488 92762
0 50724 5 1 1 50723
0 50725 7 1 2 50722 50724
0 50726 5 1 1 50725
0 50727 7 1 2 69442 98398
0 50728 7 1 2 50726 50727
0 50729 5 1 1 50728
0 50730 7 1 2 50720 50729
0 50731 7 1 2 50717 50730
0 50732 5 1 1 50731
0 50733 7 1 2 61409 50732
0 50734 5 1 1 50733
0 50735 7 1 2 88108 101537
0 50736 5 1 1 50735
0 50737 7 1 2 82385 89069
0 50738 5 1 1 50737
0 50739 7 1 2 81476 90557
0 50740 5 1 1 50739
0 50741 7 1 2 50738 50740
0 50742 5 1 1 50741
0 50743 7 1 2 86801 50742
0 50744 5 1 1 50743
0 50745 7 1 2 50736 50744
0 50746 5 1 1 50745
0 50747 7 1 2 61674 50746
0 50748 5 1 1 50747
0 50749 7 1 2 90021 89870
0 50750 7 1 2 91457 50749
0 50751 5 1 1 50750
0 50752 7 1 2 50748 50751
0 50753 5 1 1 50752
0 50754 7 1 2 100256 50753
0 50755 5 1 1 50754
0 50756 7 1 2 50734 50755
0 50757 5 1 1 50756
0 50758 7 1 2 73226 50757
0 50759 5 1 1 50758
0 50760 7 1 2 91221 102934
0 50761 7 1 2 102216 50760
0 50762 5 1 1 50761
0 50763 7 1 2 50759 50762
0 50764 5 1 1 50763
0 50765 7 1 2 65000 50764
0 50766 5 1 1 50765
0 50767 7 1 2 50704 50766
0 50768 5 1 1 50767
0 50769 7 1 2 78118 50768
0 50770 5 1 1 50769
0 50771 7 1 2 50673 50770
0 50772 5 1 1 50771
0 50773 7 1 2 62224 50772
0 50774 5 1 1 50773
0 50775 7 1 2 69634 72727
0 50776 7 1 2 90212 50775
0 50777 5 1 1 50776
0 50778 7 1 2 61915 101305
0 50779 5 1 1 50778
0 50780 7 1 2 50777 50779
0 50781 5 1 1 50780
0 50782 7 1 2 64589 50781
0 50783 5 1 1 50782
0 50784 7 1 2 92305 101733
0 50785 5 1 1 50784
0 50786 7 1 2 61675 50785
0 50787 7 1 2 50783 50786
0 50788 5 1 1 50787
0 50789 7 1 2 72728 88721
0 50790 5 1 1 50789
0 50791 7 1 2 100414 102087
0 50792 5 1 1 50791
0 50793 7 1 2 50790 50792
0 50794 5 1 1 50793
0 50795 7 1 2 69635 50794
0 50796 5 1 1 50795
0 50797 7 1 2 80173 90908
0 50798 7 1 2 90213 50797
0 50799 5 1 1 50798
0 50800 7 1 2 66567 50799
0 50801 7 1 2 50796 50800
0 50802 5 1 1 50801
0 50803 7 1 2 89577 50802
0 50804 7 1 2 50788 50803
0 50805 5 1 1 50804
0 50806 7 1 2 82754 78941
0 50807 5 1 1 50806
0 50808 7 1 2 82388 81481
0 50809 5 1 1 50808
0 50810 7 1 2 61676 50809
0 50811 7 1 2 50807 50810
0 50812 5 1 1 50811
0 50813 7 1 2 81477 87698
0 50814 5 1 1 50813
0 50815 7 1 2 50812 50814
0 50816 5 1 1 50815
0 50817 7 1 2 88045 100280
0 50818 7 1 2 50816 50817
0 50819 5 1 1 50818
0 50820 7 1 2 50805 50819
0 50821 5 1 1 50820
0 50822 7 1 2 65241 50821
0 50823 5 1 1 50822
0 50824 7 1 2 72659 75171
0 50825 7 1 2 92874 96722
0 50826 7 1 2 50824 50825
0 50827 5 1 1 50826
0 50828 7 1 2 50823 50827
0 50829 5 1 1 50828
0 50830 7 1 2 63042 50829
0 50831 5 1 1 50830
0 50832 7 1 2 93350 94795
0 50833 5 1 1 50832
0 50834 7 1 2 86934 98324
0 50835 7 1 2 91310 50834
0 50836 5 1 1 50835
0 50837 7 1 2 50833 50836
0 50838 5 1 1 50837
0 50839 7 2 2 83400 50838
0 50840 7 1 2 98050 102938
0 50841 5 1 1 50840
0 50842 7 1 2 50831 50841
0 50843 5 1 1 50842
0 50844 7 1 2 61410 50843
0 50845 5 1 1 50844
0 50846 7 1 2 101325 99599
0 50847 5 1 1 50846
0 50848 7 1 2 74502 99665
0 50849 5 1 1 50848
0 50850 7 1 2 50847 50849
0 50851 5 1 1 50850
0 50852 7 1 2 88715 50851
0 50853 5 1 1 50852
0 50854 7 1 2 72735 99600
0 50855 5 1 1 50854
0 50856 7 1 2 50855 102724
0 50857 5 1 1 50856
0 50858 7 1 2 96248 50857
0 50859 5 1 1 50858
0 50860 7 1 2 50853 50859
0 50861 5 1 1 50860
0 50862 7 1 2 82789 50861
0 50863 5 1 1 50862
0 50864 7 1 2 83637 100335
0 50865 7 1 2 101326 50864
0 50866 5 1 1 50865
0 50867 7 1 2 50863 50866
0 50868 5 1 1 50867
0 50869 7 1 2 61411 50868
0 50870 5 1 1 50869
0 50871 7 1 2 83216 86658
0 50872 5 1 1 50871
0 50873 7 1 2 89204 76869
0 50874 5 1 1 50873
0 50875 7 1 2 50872 50874
0 50876 5 1 1 50875
0 50877 7 1 2 62225 50876
0 50878 5 1 1 50877
0 50879 7 1 2 66041 78087
0 50880 7 1 2 78798 50879
0 50881 5 1 1 50880
0 50882 7 1 2 50878 50881
0 50883 5 1 1 50882
0 50884 7 1 2 69055 50883
0 50885 5 1 1 50884
0 50886 7 1 2 78048 86047
0 50887 5 1 1 50886
0 50888 7 1 2 50885 50887
0 50889 5 1 1 50888
0 50890 7 1 2 82795 93764
0 50891 7 1 2 50889 50890
0 50892 5 1 1 50891
0 50893 7 1 2 50870 50892
0 50894 5 1 1 50893
0 50895 7 1 2 76194 50894
0 50896 5 1 1 50895
0 50897 7 1 2 72729 102754
0 50898 5 1 1 50897
0 50899 7 1 2 100415 100768
0 50900 5 1 1 50899
0 50901 7 1 2 50898 50900
0 50902 5 1 1 50901
0 50903 7 1 2 50902 99844
0 50904 5 1 1 50903
0 50905 7 1 2 79086 94285
0 50906 7 1 2 102916 50905
0 50907 5 1 1 50906
0 50908 7 1 2 50904 50907
0 50909 5 1 1 50908
0 50910 7 1 2 65242 50909
0 50911 5 1 1 50910
0 50912 7 1 2 50896 50911
0 50913 5 1 1 50912
0 50914 7 1 2 83163 50913
0 50915 5 1 1 50914
0 50916 7 1 2 101534 102273
0 50917 5 1 1 50916
0 50918 7 1 2 72660 102748
0 50919 7 1 2 91311 50918
0 50920 5 1 1 50919
0 50921 7 1 2 50917 50920
0 50922 5 1 1 50921
0 50923 7 1 2 65001 50922
0 50924 5 1 1 50923
0 50925 7 1 2 94695 96157
0 50926 7 1 2 102755 50925
0 50927 5 1 1 50926
0 50928 7 1 2 50924 50927
0 50929 5 1 1 50928
0 50930 7 1 2 95000 50929
0 50931 5 1 1 50930
0 50932 7 1 2 102939 102741
0 50933 5 1 1 50932
0 50934 7 1 2 50931 50933
0 50935 7 1 2 50915 50934
0 50936 7 1 2 50845 50935
0 50937 5 1 1 50936
0 50938 7 1 2 70471 50937
0 50939 5 1 1 50938
0 50940 7 1 2 79087 91312
0 50941 5 1 1 50940
0 50942 7 1 2 69857 102851
0 50943 5 1 1 50942
0 50944 7 1 2 50941 50943
0 50945 5 1 1 50944
0 50946 7 1 2 70964 50945
0 50947 5 1 1 50946
0 50948 7 1 2 89348 91995
0 50949 5 1 1 50948
0 50950 7 1 2 50947 50949
0 50951 5 1 1 50950
0 50952 7 1 2 64197 50951
0 50953 5 1 1 50952
0 50954 7 1 2 95832 96695
0 50955 5 1 1 50954
0 50956 7 1 2 50953 50955
0 50957 5 1 1 50956
0 50958 7 1 2 62913 50957
0 50959 5 1 1 50958
0 50960 7 1 2 78817 92875
0 50961 5 1 1 50960
0 50962 7 1 2 50959 50961
0 50963 5 1 1 50962
0 50964 7 1 2 62666 96249
0 50965 7 1 2 102762 50964
0 50966 7 1 2 50963 50965
0 50967 5 1 1 50966
0 50968 7 1 2 50939 50967
0 50969 5 1 1 50968
0 50970 7 1 2 71605 50969
0 50971 5 1 1 50970
0 50972 7 1 2 93827 96477
0 50973 5 1 1 50972
0 50974 7 1 2 50567 50973
0 50975 5 1 1 50974
0 50976 7 1 2 87315 50975
0 50977 5 1 1 50976
0 50978 7 1 2 79088 102217
0 50979 5 1 1 50978
0 50980 7 1 2 50977 50979
0 50981 5 1 1 50980
0 50982 7 1 2 88716 50981
0 50983 5 1 1 50982
0 50984 7 1 2 79186 100762
0 50985 5 1 1 50984
0 50986 7 1 2 99390 97502
0 50987 5 1 1 50986
0 50988 7 1 2 50985 50987
0 50989 5 1 1 50988
0 50990 7 1 2 92712 50989
0 50991 5 1 1 50990
0 50992 7 2 2 100236 100577
0 50993 5 1 1 102940
0 50994 7 1 2 101590 99851
0 50995 5 1 1 50994
0 50996 7 1 2 50993 50995
0 50997 5 1 1 50996
0 50998 7 1 2 94917 50997
0 50999 5 1 1 50998
0 51000 7 1 2 61412 102442
0 51001 5 1 1 51000
0 51002 7 1 2 93083 102742
0 51003 5 1 1 51002
0 51004 7 1 2 51001 51003
0 51005 5 1 1 51004
0 51006 7 1 2 81958 100237
0 51007 5 1 1 51006
0 51008 7 1 2 92041 51007
0 51009 5 1 1 51008
0 51010 7 1 2 51005 51009
0 51011 5 1 1 51010
0 51012 7 1 2 50999 51011
0 51013 7 1 2 50991 51012
0 51014 5 1 1 51013
0 51015 7 1 2 65243 51014
0 51016 5 1 1 51015
0 51017 7 1 2 50983 51016
0 51018 5 1 1 51017
0 51019 7 1 2 85088 102935
0 51020 7 1 2 51018 51019
0 51021 5 1 1 51020
0 51022 7 1 2 98403 100124
0 51023 7 1 2 82360 51022
0 51024 7 1 2 96723 96984
0 51025 7 1 2 51023 51024
0 51026 5 1 1 51025
0 51027 7 1 2 51021 51026
0 51028 5 1 1 51027
0 51029 7 1 2 72199 51028
0 51030 5 1 1 51029
0 51031 7 2 2 93828 102058
0 51032 7 1 2 102928 102942
0 51033 5 1 1 51032
0 51034 7 1 2 83657 90626
0 51035 7 1 2 102932 51034
0 51036 5 1 1 51035
0 51037 7 1 2 51033 51036
0 51038 5 1 1 51037
0 51039 7 1 2 73227 51038
0 51040 5 1 1 51039
0 51041 7 1 2 72470 95411
0 51042 7 1 2 102943 51041
0 51043 5 1 1 51042
0 51044 7 1 2 51040 51043
0 51045 5 1 1 51044
0 51046 7 1 2 76195 51045
0 51047 5 1 1 51046
0 51048 7 1 2 97173 102937
0 51049 5 1 1 51048
0 51050 7 1 2 51047 51049
0 51051 5 1 1 51050
0 51052 7 1 2 83164 51051
0 51053 5 1 1 51052
0 51054 7 1 2 89279 102924
0 51055 5 1 1 51054
0 51056 7 1 2 79882 91611
0 51057 5 1 1 51056
0 51058 7 1 2 82065 102689
0 51059 5 1 1 51058
0 51060 7 1 2 51057 51059
0 51061 5 1 1 51060
0 51062 7 1 2 72083 51061
0 51063 5 1 1 51062
0 51064 7 1 2 102785 99925
0 51065 5 1 1 51064
0 51066 7 1 2 51063 51065
0 51067 5 1 1 51066
0 51068 7 1 2 90273 90627
0 51069 7 1 2 51067 51068
0 51070 5 1 1 51069
0 51071 7 1 2 51055 51070
0 51072 5 1 1 51071
0 51073 7 1 2 90214 51072
0 51074 5 1 1 51073
0 51075 7 1 2 81959 87624
0 51076 5 1 1 51075
0 51077 7 1 2 80633 99823
0 51078 5 1 1 51077
0 51079 7 1 2 51076 51078
0 51080 5 1 1 51079
0 51081 7 1 2 102690 51080
0 51082 5 1 1 51081
0 51083 7 1 2 73101 87485
0 51084 7 1 2 102778 51083
0 51085 5 1 1 51084
0 51086 7 1 2 51082 51085
0 51087 5 1 1 51086
0 51088 7 1 2 72084 51087
0 51089 5 1 1 51088
0 51090 7 1 2 71746 93385
0 51091 7 1 2 102779 51090
0 51092 5 1 1 51091
0 51093 7 1 2 51089 51092
0 51094 5 1 1 51093
0 51095 7 1 2 102841 51094
0 51096 5 1 1 51095
0 51097 7 1 2 87625 80386
0 51098 7 1 2 102844 51097
0 51099 5 1 1 51098
0 51100 7 1 2 51096 51099
0 51101 7 1 2 51074 51100
0 51102 7 1 2 51053 51101
0 51103 5 1 1 51102
0 51104 7 1 2 67061 51103
0 51105 5 1 1 51104
0 51106 7 1 2 51030 51105
0 51107 7 1 2 50971 51106
0 51108 7 1 2 50774 51107
0 51109 5 1 1 51108
0 51110 7 1 2 69252 51109
0 51111 5 1 1 51110
0 51112 7 1 2 96954 51111
0 51113 5 1 1 51112
0 51114 7 1 2 64297 92660
0 51115 7 1 2 51113 51114
0 51116 7 1 2 50518 51115
0 51117 5 1 1 51116
0 51118 7 1 2 48996 51117
0 51119 5 1 1 51118
0 51120 7 1 2 74851 51119
0 51121 5 1 1 51120
0 51122 7 1 2 70472 94533
0 51123 5 1 1 51122
0 51124 7 1 2 84039 51123
0 51125 5 2 1 51124
0 51126 7 2 2 70155 102944
0 51127 7 2 2 92731 102946
0 51128 7 1 2 98622 102948
0 51129 5 1 1 51128
0 51130 7 2 2 92936 99742
0 51131 7 1 2 84388 93496
0 51132 5 1 1 51131
0 51133 7 1 2 6730 102730
0 51134 7 1 2 51132 51133
0 51135 5 1 1 51134
0 51136 7 1 2 102950 51135
0 51137 5 1 1 51136
0 51138 7 1 2 51129 51137
0 51139 5 1 1 51138
0 51140 7 1 2 61320 51139
0 51141 5 1 1 51140
0 51142 7 1 2 102949 100383
0 51143 5 1 1 51142
0 51144 7 1 2 51141 51143
0 51145 5 1 1 51144
0 51146 7 1 2 93829 51145
0 51147 5 1 1 51146
0 51148 7 1 2 85665 92897
0 51149 5 1 1 51148
0 51150 7 1 2 82460 93309
0 51151 5 1 1 51150
0 51152 7 1 2 51149 51151
0 51153 5 1 1 51152
0 51154 7 1 2 62914 93670
0 51155 5 1 1 51154
0 51156 7 1 2 84323 83366
0 51157 5 1 1 51156
0 51158 7 1 2 51155 51157
0 51159 5 5 1 51158
0 51160 7 1 2 51153 102952
0 51161 5 1 1 51160
0 51162 7 1 2 73131 90448
0 51163 5 1 1 51162
0 51164 7 2 2 85728 85903
0 51165 5 2 1 102957
0 51166 7 1 2 86102 102959
0 51167 5 4 1 51166
0 51168 7 1 2 74743 12613
0 51169 5 2 1 51168
0 51170 7 1 2 102961 102965
0 51171 5 1 1 51170
0 51172 7 1 2 51163 51171
0 51173 7 1 2 51161 51172
0 51174 5 1 1 51173
0 51175 7 1 2 91033 51174
0 51176 5 1 1 51175
0 51177 7 1 2 51147 51176
0 51178 5 1 1 51177
0 51179 7 1 2 64298 51178
0 51180 5 1 1 51179
0 51181 7 1 2 68876 96714
0 51182 5 1 1 51181
0 51183 7 1 2 96708 51182
0 51184 5 1 1 51183
0 51185 7 1 2 99601 51184
0 51186 5 1 1 51185
0 51187 7 1 2 69056 99666
0 51188 7 1 2 100963 51187
0 51189 5 1 1 51188
0 51190 7 1 2 72200 99602
0 51191 7 1 2 96718 51190
0 51192 5 1 1 51191
0 51193 7 1 2 51189 51192
0 51194 5 1 1 51193
0 51195 7 1 2 67741 51194
0 51196 5 1 1 51195
0 51197 7 1 2 51186 51196
0 51198 5 1 1 51197
0 51199 7 1 2 66308 51198
0 51200 5 1 1 51199
0 51201 7 1 2 91247 101211
0 51202 5 1 1 51201
0 51203 7 1 2 76949 51202
0 51204 5 1 1 51203
0 51205 7 1 2 96716 51204
0 51206 5 1 1 51205
0 51207 7 1 2 100554 51206
0 51208 5 1 1 51207
0 51209 7 1 2 51200 51208
0 51210 5 1 1 51209
0 51211 7 1 2 67532 51210
0 51212 5 1 1 51211
0 51213 7 2 2 92866 93548
0 51214 5 1 1 102967
0 51215 7 1 2 84389 72471
0 51216 5 1 1 51215
0 51217 7 1 2 51214 51216
0 51218 5 1 1 51217
0 51219 7 1 2 77926 101949
0 51220 7 1 2 51218 51219
0 51221 5 1 1 51220
0 51222 7 1 2 51212 51221
0 51223 5 1 1 51222
0 51224 7 1 2 67062 51223
0 51225 5 1 1 51224
0 51226 7 1 2 85846 100205
0 51227 5 1 1 51226
0 51228 7 1 2 49984 51227
0 51229 5 1 1 51228
0 51230 7 1 2 94056 96472
0 51231 7 1 2 51229 51230
0 51232 5 1 1 51231
0 51233 7 1 2 51225 51232
0 51234 5 1 1 51233
0 51235 7 1 2 78485 51234
0 51236 5 1 1 51235
0 51237 7 1 2 75308 99583
0 51238 7 1 2 89228 51237
0 51239 5 1 1 51238
0 51240 7 1 2 99667 102953
0 51241 5 1 1 51240
0 51242 7 1 2 64198 100305
0 51243 5 1 1 51242
0 51244 7 1 2 51241 51243
0 51245 5 1 1 51244
0 51246 7 1 2 78486 78830
0 51247 7 1 2 51245 51246
0 51248 5 1 1 51247
0 51249 7 1 2 51239 51248
0 51250 5 1 1 51249
0 51251 7 1 2 66309 51250
0 51252 5 1 1 51251
0 51253 7 1 2 78786 101248
0 51254 7 1 2 100565 51253
0 51255 5 1 1 51254
0 51256 7 1 2 51252 51255
0 51257 5 1 1 51256
0 51258 7 1 2 73132 51257
0 51259 5 1 1 51258
0 51260 7 1 2 72925 102968
0 51261 5 2 1 51260
0 51262 7 1 2 67742 92402
0 51263 5 2 1 51262
0 51264 7 1 2 102971 41070
0 51265 5 1 1 51264
0 51266 7 1 2 65864 51265
0 51267 5 1 1 51266
0 51268 7 1 2 5867 75900
0 51269 7 1 2 92405 51268
0 51270 5 1 1 51269
0 51271 7 1 2 51267 51270
0 51272 5 1 1 51271
0 51273 7 1 2 69057 51272
0 51274 5 1 1 51273
0 51275 7 1 2 73585 85738
0 51276 7 1 2 95858 51275
0 51277 5 1 1 51276
0 51278 7 1 2 51274 51277
0 51279 5 1 1 51278
0 51280 7 1 2 70473 51279
0 51281 5 1 1 51280
0 51282 7 1 2 102969 51281
0 51283 5 1 1 51282
0 51284 7 1 2 83641 101296
0 51285 7 1 2 51283 51284
0 51286 5 1 1 51285
0 51287 7 1 2 51259 51286
0 51288 7 1 2 51236 51287
0 51289 5 1 1 51288
0 51290 7 1 2 97319 51289
0 51291 5 1 1 51290
0 51292 7 1 2 51180 51291
0 51293 5 1 1 51292
0 51294 7 1 2 69253 51293
0 51295 5 1 1 51294
0 51296 7 2 2 82086 102945
0 51297 7 1 2 98340 102973
0 51298 5 1 1 51297
0 51299 7 1 2 74132 89951
0 51300 5 1 1 51299
0 51301 7 1 2 90446 51300
0 51302 5 1 1 51301
0 51303 7 1 2 65865 1218
0 51304 7 1 2 51302 51303
0 51305 5 1 1 51304
0 51306 7 1 2 70764 84691
0 51307 7 1 2 89590 51306
0 51308 5 1 1 51307
0 51309 7 1 2 51305 51308
0 51310 5 1 1 51309
0 51311 7 1 2 84905 51310
0 51312 5 1 1 51311
0 51313 7 1 2 70474 51312
0 51314 5 1 1 51313
0 51315 7 1 2 100873 51314
0 51316 5 1 1 51315
0 51317 7 1 2 102316 98623
0 51318 7 1 2 51316 51317
0 51319 5 1 1 51318
0 51320 7 1 2 51298 51319
0 51321 5 1 1 51320
0 51322 7 1 2 66175 51321
0 51323 5 1 1 51322
0 51324 7 1 2 67063 92964
0 51325 7 1 2 102974 51324
0 51326 5 1 1 51325
0 51327 7 1 2 51323 51326
0 51328 5 1 1 51327
0 51329 7 1 2 69144 51328
0 51330 5 1 1 51329
0 51331 7 1 2 78342 95133
0 51332 5 2 1 51331
0 51333 7 1 2 132 102975
0 51334 5 2 1 51333
0 51335 7 1 2 97721 99765
0 51336 7 1 2 86097 51335
0 51337 7 1 2 102977 51336
0 51338 5 1 1 51337
0 51339 7 1 2 51330 51338
0 51340 5 1 1 51339
0 51341 7 1 2 93830 51340
0 51342 5 1 1 51341
0 51343 7 4 2 66042 80583
0 51344 7 1 2 102979 101223
0 51345 5 1 1 51344
0 51346 7 1 2 78831 101194
0 51347 5 1 1 51346
0 51348 7 1 2 51345 51347
0 51349 5 1 1 51348
0 51350 7 1 2 69058 51349
0 51351 5 1 1 51350
0 51352 7 2 2 64199 86202
0 51353 5 2 1 102983
0 51354 7 1 2 80662 102984
0 51355 5 1 1 51354
0 51356 7 1 2 51351 51355
0 51357 5 1 1 51356
0 51358 7 1 2 98669 51357
0 51359 5 1 1 51358
0 51360 7 2 2 79690 100355
0 51361 5 1 1 102987
0 51362 7 1 2 65544 51361
0 51363 5 1 1 51362
0 51364 7 1 2 85373 51363
0 51365 5 1 1 51364
0 51366 7 1 2 65244 98656
0 51367 7 1 2 51365 51366
0 51368 5 1 1 51367
0 51369 7 1 2 51359 51368
0 51370 5 1 1 51369
0 51371 7 1 2 79646 51370
0 51372 5 1 1 51371
0 51373 7 2 2 100353 102985
0 51374 5 5 1 102989
0 51375 7 1 2 82684 101148
0 51376 7 1 2 90086 51375
0 51377 7 1 2 102991 51376
0 51378 7 1 2 92488 51377
0 51379 5 1 1 51378
0 51380 7 1 2 51372 51379
0 51381 5 1 1 51380
0 51382 7 1 2 73494 51381
0 51383 5 1 1 51382
0 51384 7 1 2 65545 78360
0 51385 5 1 1 51384
0 51386 7 1 2 74728 51385
0 51387 5 1 1 51386
0 51388 7 1 2 102958 51387
0 51389 5 1 1 51388
0 51390 7 1 2 87506 102744
0 51391 5 1 1 51390
0 51392 7 1 2 51389 51391
0 51393 5 1 1 51392
0 51394 7 1 2 98670 51393
0 51395 5 1 1 51394
0 51396 7 1 2 84347 93310
0 51397 5 1 1 51396
0 51398 7 1 2 86935 90087
0 51399 7 1 2 102895 51398
0 51400 5 1 1 51399
0 51401 7 1 2 51397 51400
0 51402 5 1 1 51401
0 51403 7 1 2 98657 51402
0 51404 5 1 1 51403
0 51405 7 1 2 51395 51404
0 51406 5 1 1 51405
0 51407 7 1 2 71370 51406
0 51408 5 1 1 51407
0 51409 7 1 2 62915 98658
0 51410 7 1 2 102962 51409
0 51411 5 1 1 51410
0 51412 7 1 2 51408 51411
0 51413 7 1 2 51383 51412
0 51414 7 1 2 51342 51413
0 51415 5 1 1 51414
0 51416 7 1 2 64395 51415
0 51417 5 1 1 51416
0 51418 7 1 2 92489 102963
0 51419 5 1 1 51418
0 51420 7 1 2 102317 97585
0 51421 7 1 2 99683 51420
0 51422 5 1 1 51421
0 51423 7 1 2 51419 51422
0 51424 5 1 1 51423
0 51425 7 1 2 64396 51424
0 51426 5 1 1 51425
0 51427 7 3 2 92810 93831
0 51428 7 2 2 92937 102996
0 51429 7 1 2 99966 97586
0 51430 7 1 2 102999 51429
0 51431 5 1 1 51430
0 51432 7 1 2 51426 51431
0 51433 5 1 1 51432
0 51434 7 1 2 71371 51433
0 51435 5 1 1 51434
0 51436 7 2 2 90881 87873
0 51437 7 2 2 92840 98051
0 51438 7 1 2 83642 103003
0 51439 7 1 2 103001 51438
0 51440 5 1 1 51439
0 51441 7 1 2 78683 72230
0 51442 7 1 2 96064 51441
0 51443 7 1 2 99054 51442
0 51444 5 1 1 51443
0 51445 7 1 2 51440 51444
0 51446 5 1 1 51445
0 51447 7 1 2 64590 51446
0 51448 5 1 1 51447
0 51449 7 1 2 51435 51448
0 51450 5 1 1 51449
0 51451 7 1 2 70765 51450
0 51452 5 1 1 51451
0 51453 7 1 2 84577 99378
0 51454 7 1 2 103000 51453
0 51455 5 1 1 51454
0 51456 7 1 2 51452 51455
0 51457 5 1 1 51456
0 51458 7 1 2 65546 51457
0 51459 5 1 1 51458
0 51460 7 1 2 62226 97191
0 51461 5 1 1 51460
0 51462 7 1 2 87134 97179
0 51463 7 1 2 85575 51462
0 51464 5 1 1 51463
0 51465 7 1 2 51461 51464
0 51466 5 1 1 51465
0 51467 7 1 2 99099 51466
0 51468 5 1 1 51467
0 51469 7 1 2 1184 79703
0 51470 5 6 1 51469
0 51471 7 1 2 69254 78201
0 51472 7 2 2 103005 51471
0 51473 7 1 2 86144 102424
0 51474 7 1 2 103011 51473
0 51475 5 1 1 51474
0 51476 7 1 2 51468 51475
0 51477 5 1 1 51476
0 51478 7 1 2 92664 51477
0 51479 5 1 1 51478
0 51480 7 1 2 69145 51479
0 51481 7 1 2 51459 51480
0 51482 5 1 1 51481
0 51483 7 1 2 67064 41695
0 51484 5 3 1 51483
0 51485 7 1 2 93606 103013
0 51486 5 1 1 51485
0 51487 7 1 2 98624 98592
0 51488 5 1 1 51487
0 51489 7 1 2 51486 51488
0 51490 5 1 1 51489
0 51491 7 1 2 102318 51490
0 51492 5 1 1 51491
0 51493 7 1 2 62227 86514
0 51494 5 3 1 51493
0 51495 7 2 2 69255 99743
0 51496 7 1 2 92938 103019
0 51497 7 1 2 103016 51496
0 51498 5 1 1 51497
0 51499 7 1 2 51492 51498
0 51500 5 1 1 51499
0 51501 7 1 2 61321 51500
0 51502 5 1 1 51501
0 51503 7 1 2 79665 102125
0 51504 7 1 2 100384 51503
0 51505 5 1 1 51504
0 51506 7 1 2 51502 51505
0 51507 5 1 1 51506
0 51508 7 1 2 99100 51507
0 51509 5 1 1 51508
0 51510 7 1 2 67065 2323
0 51511 5 3 1 51510
0 51512 7 1 2 83662 103021
0 51513 5 1 1 51512
0 51514 7 1 2 102960 51513
0 51515 5 1 1 51514
0 51516 7 1 2 91358 51515
0 51517 5 1 1 51516
0 51518 7 1 2 64299 51517
0 51519 7 1 2 51509 51518
0 51520 5 1 1 51519
0 51521 7 1 2 72661 51520
0 51522 7 1 2 51482 51521
0 51523 5 1 1 51522
0 51524 7 1 2 51417 51523
0 51525 7 1 2 51295 51524
0 51526 5 1 1 51525
0 51527 7 1 2 76196 51526
0 51528 5 1 1 51527
0 51529 7 2 2 87826 102190
0 51530 7 1 2 93583 103024
0 51531 5 1 1 51530
0 51532 7 1 2 62916 99732
0 51533 5 1 1 51532
0 51534 7 1 2 48773 51533
0 51535 5 1 1 51534
0 51536 7 1 2 64397 72662
0 51537 7 1 2 51535 51536
0 51538 5 1 1 51537
0 51539 7 1 2 51531 51538
0 51540 5 1 1 51539
0 51541 7 1 2 64002 51540
0 51542 5 1 1 51541
0 51543 7 2 2 66310 88383
0 51544 7 1 2 72806 93607
0 51545 7 1 2 103026 51544
0 51546 5 1 1 51545
0 51547 7 1 2 51542 51546
0 51548 5 1 1 51547
0 51549 7 1 2 100675 51548
0 51550 5 1 1 51549
0 51551 7 2 2 64591 99277
0 51552 7 1 2 72085 103028
0 51553 5 2 1 51552
0 51554 7 1 2 89307 103030
0 51555 5 1 1 51554
0 51556 7 4 2 62917 100004
0 51557 5 1 1 103032
0 51558 7 1 2 99519 51557
0 51559 5 2 1 51558
0 51560 7 1 2 64398 100591
0 51561 7 2 2 103036 51560
0 51562 7 1 2 51555 103038
0 51563 5 1 1 51562
0 51564 7 1 2 99584 103025
0 51565 7 1 2 100784 51564
0 51566 5 1 1 51565
0 51567 7 1 2 51563 51566
0 51568 7 1 2 51550 51567
0 51569 5 1 1 51568
0 51570 7 1 2 70766 51569
0 51571 5 1 1 51570
0 51572 7 1 2 96486 99033
0 51573 5 1 1 51572
0 51574 7 1 2 93136 100752
0 51575 5 1 1 51574
0 51576 7 1 2 51573 51575
0 51577 5 1 1 51576
0 51578 7 1 2 93554 51577
0 51579 5 1 1 51578
0 51580 7 1 2 86893 102714
0 51581 5 2 1 51580
0 51582 7 1 2 92811 103040
0 51583 7 1 2 101445 51582
0 51584 5 1 1 51583
0 51585 7 1 2 51579 51584
0 51586 5 1 1 51585
0 51587 7 1 2 67820 51586
0 51588 5 1 1 51587
0 51589 7 1 2 84563 92181
0 51590 5 1 1 51589
0 51591 7 1 2 93639 51590
0 51592 5 1 1 51591
0 51593 7 1 2 99754 51592
0 51594 5 1 1 51593
0 51595 7 2 2 91648 100366
0 51596 5 1 1 103042
0 51597 7 1 2 97587 103043
0 51598 5 1 1 51597
0 51599 7 1 2 51594 51598
0 51600 5 1 1 51599
0 51601 7 1 2 100676 51600
0 51602 5 1 1 51601
0 51603 7 1 2 70767 103039
0 51604 5 1 1 51603
0 51605 7 1 2 96232 97588
0 51606 7 1 2 101436 51605
0 51607 5 1 1 51606
0 51608 7 1 2 51604 51607
0 51609 7 1 2 51602 51608
0 51610 5 1 1 51609
0 51611 7 1 2 72663 51610
0 51612 5 1 1 51611
0 51613 7 2 2 90696 100941
0 51614 5 3 1 103044
0 51615 7 1 2 93555 103045
0 51616 5 1 1 51615
0 51617 7 1 2 51612 51616
0 51618 7 1 2 51588 51617
0 51619 5 1 1 51618
0 51620 7 1 2 62667 51619
0 51621 5 1 1 51620
0 51622 7 1 2 51571 51621
0 51623 5 1 1 51622
0 51624 7 1 2 102279 51623
0 51625 5 1 1 51624
0 51626 7 1 2 44637 42163
0 51627 5 3 1 51626
0 51628 7 1 2 62985 93058
0 51629 5 2 1 51628
0 51630 7 1 2 99700 97589
0 51631 5 1 1 51630
0 51632 7 1 2 103052 51631
0 51633 5 1 1 51632
0 51634 7 1 2 103049 51633
0 51635 5 1 1 51634
0 51636 7 1 2 99611 36328
0 51637 5 1 1 51636
0 51638 7 1 2 32860 36529
0 51639 7 1 2 100586 51638
0 51640 7 1 2 51637 51639
0 51641 5 1 1 51640
0 51642 7 1 2 51635 51641
0 51643 5 2 1 51642
0 51644 7 1 2 89294 103054
0 51645 5 1 1 51644
0 51646 7 2 2 72086 88902
0 51647 7 1 2 61413 100592
0 51648 5 1 1 51647
0 51649 7 1 2 90948 100677
0 51650 5 1 1 51649
0 51651 7 1 2 51648 51650
0 51652 5 1 1 51651
0 51653 7 1 2 103056 51652
0 51654 5 1 1 51653
0 51655 7 1 2 51645 51654
0 51656 5 1 1 51655
0 51657 7 1 2 93629 51656
0 51658 5 1 1 51657
0 51659 7 1 2 92812 99585
0 51660 5 1 1 51659
0 51661 7 1 2 101686 51660
0 51662 5 2 1 51661
0 51663 7 1 2 103058 103050
0 51664 5 1 1 51663
0 51665 7 2 2 92813 93584
0 51666 5 1 1 103060
0 51667 7 1 2 100669 103061
0 51668 5 1 1 51667
0 51669 7 1 2 100223 100690
0 51670 5 2 1 51669
0 51671 7 1 2 51668 103062
0 51672 7 1 2 51664 51671
0 51673 5 1 1 51672
0 51674 7 1 2 67821 51673
0 51675 5 1 1 51674
0 51676 7 1 2 51675 103046
0 51677 5 1 1 51676
0 51678 7 1 2 93556 51677
0 51679 5 1 1 51678
0 51680 7 1 2 72664 93630
0 51681 7 1 2 103055 51680
0 51682 5 1 1 51681
0 51683 7 1 2 51679 51682
0 51684 5 1 1 51683
0 51685 7 1 2 62668 51684
0 51686 5 1 1 51685
0 51687 7 1 2 51658 51686
0 51688 5 1 1 51687
0 51689 7 1 2 78832 51688
0 51690 5 1 1 51689
0 51691 7 1 2 102196 103051
0 51692 5 1 1 51691
0 51693 7 3 2 66311 80942
0 51694 7 1 2 92560 92814
0 51695 7 1 2 103064 51694
0 51696 5 1 1 51695
0 51697 7 1 2 103063 51696
0 51698 7 1 2 51692 51697
0 51699 5 1 1 51698
0 51700 7 1 2 67822 51699
0 51701 5 1 1 51700
0 51702 7 1 2 103047 51701
0 51703 5 1 1 51702
0 51704 7 2 2 67533 80584
0 51705 7 1 2 100864 103067
0 51706 7 1 2 51703 51705
0 51707 5 1 1 51706
0 51708 7 1 2 51690 51707
0 51709 5 1 1 51708
0 51710 7 1 2 79089 51709
0 51711 5 1 1 51710
0 51712 7 1 2 65547 51711
0 51713 7 1 2 51625 51712
0 51714 5 1 1 51713
0 51715 7 3 2 61677 64399
0 51716 7 1 2 70965 98112
0 51717 7 1 2 103069 51716
0 51718 7 1 2 91615 51717
0 51719 5 1 1 51718
0 51720 7 2 2 87985 94488
0 51721 5 1 1 103072
0 51722 7 2 2 80997 100134
0 51723 7 1 2 5263 103074
0 51724 7 1 2 51721 51723
0 51725 5 1 1 51724
0 51726 7 1 2 51719 51725
0 51727 5 1 1 51726
0 51728 7 1 2 66312 51727
0 51729 5 1 1 51728
0 51730 7 1 2 91616 95545
0 51731 7 1 2 100753 51730
0 51732 5 1 1 51731
0 51733 7 1 2 51729 51732
0 51734 5 1 1 51733
0 51735 7 1 2 67534 51734
0 51736 5 1 1 51735
0 51737 7 1 2 67743 100395
0 51738 5 1 1 51737
0 51739 7 1 2 100438 51738
0 51740 5 1 1 51739
0 51741 7 1 2 64400 51740
0 51742 7 1 2 100763 51741
0 51743 5 1 1 51742
0 51744 7 1 2 51736 51743
0 51745 5 1 1 51744
0 51746 7 1 2 102280 51745
0 51747 5 1 1 51746
0 51748 7 2 2 70966 7277
0 51749 5 1 1 103076
0 51750 7 1 2 51749 100439
0 51751 5 2 1 51750
0 51752 7 1 2 64401 102275
0 51753 7 1 2 100764 51752
0 51754 7 1 2 103078 51753
0 51755 5 1 1 51754
0 51756 7 1 2 51747 51755
0 51757 5 1 1 51756
0 51758 7 1 2 69443 51757
0 51759 5 1 1 51758
0 51760 7 5 2 64402 102282
0 51761 7 1 2 85769 101453
0 51762 7 1 2 103080 51761
0 51763 5 1 1 51762
0 51764 7 1 2 102283 100432
0 51765 5 1 1 51764
0 51766 7 1 2 89122 81152
0 51767 7 1 2 82477 51766
0 51768 5 1 1 51767
0 51769 7 1 2 51765 51768
0 51770 5 1 1 51769
0 51771 7 1 2 69256 101446
0 51772 7 1 2 51770 51771
0 51773 5 1 1 51772
0 51774 7 1 2 51763 51773
0 51775 5 1 1 51774
0 51776 7 1 2 64592 51775
0 51777 5 1 1 51776
0 51778 7 1 2 67823 51777
0 51779 7 1 2 51759 51778
0 51780 5 1 1 51779
0 51781 7 1 2 85770 101914
0 51782 5 1 1 51781
0 51783 7 1 2 101927 103079
0 51784 5 1 1 51783
0 51785 7 1 2 51782 51784
0 51786 5 1 1 51785
0 51787 7 1 2 103081 51786
0 51788 5 1 1 51787
0 51789 7 1 2 62986 51788
0 51790 5 1 1 51789
0 51791 7 1 2 64200 51790
0 51792 7 1 2 51780 51791
0 51793 5 1 1 51792
0 51794 7 1 2 89946 102668
0 51795 5 1 1 51794
0 51796 7 3 2 66043 86842
0 51797 7 1 2 99733 103085
0 51798 5 1 1 51797
0 51799 7 1 2 51795 51798
0 51800 5 1 1 51799
0 51801 7 1 2 103082 51800
0 51802 5 1 1 51801
0 51803 7 1 2 81131 99755
0 51804 7 1 2 95736 51803
0 51805 7 1 2 99854 51804
0 51806 5 1 1 51805
0 51807 7 1 2 51802 51806
0 51808 5 1 1 51807
0 51809 7 1 2 100678 51808
0 51810 5 1 1 51809
0 51811 7 1 2 89947 99493
0 51812 5 1 1 51811
0 51813 7 1 2 100005 103086
0 51814 5 1 1 51813
0 51815 7 1 2 51812 51814
0 51816 5 1 1 51815
0 51817 7 1 2 100593 103083
0 51818 7 1 2 51816 51817
0 51819 5 1 1 51818
0 51820 7 1 2 91364 93689
0 51821 7 1 2 92125 51820
0 51822 7 1 2 95737 102781
0 51823 7 1 2 51821 51822
0 51824 5 1 1 51823
0 51825 7 1 2 70475 51824
0 51826 7 1 2 51819 51825
0 51827 7 1 2 51810 51826
0 51828 7 1 2 51793 51827
0 51829 5 1 1 51828
0 51830 7 1 2 66176 51829
0 51831 7 1 2 51714 51830
0 51832 5 1 1 51831
0 51833 7 1 2 83429 91887
0 51834 7 1 2 66044 72354
0 51835 5 1 1 51834
0 51836 7 1 2 97181 51835
0 51837 7 1 2 51833 51836
0 51838 7 1 2 99268 51837
0 51839 5 1 1 51838
0 51840 7 1 2 72352 93644
0 51841 5 1 1 51840
0 51842 7 1 2 75368 93608
0 51843 5 1 1 51842
0 51844 7 2 2 51841 51843
0 51845 5 1 1 103088
0 51846 7 1 2 92997 97454
0 51847 5 1 1 51846
0 51848 7 1 2 103089 51847
0 51849 5 1 1 51848
0 51850 7 1 2 66045 51849
0 51851 5 1 1 51850
0 51852 7 1 2 91109 102341
0 51853 5 1 1 51852
0 51854 7 1 2 51851 51853
0 51855 5 1 1 51854
0 51856 7 1 2 101447 51855
0 51857 5 1 1 51856
0 51858 7 1 2 91113 29471
0 51859 5 2 1 51858
0 51860 7 1 2 90645 100441
0 51861 7 1 2 103090 51860
0 51862 5 1 1 51861
0 51863 7 1 2 64593 51862
0 51864 7 1 2 51857 51863
0 51865 5 1 1 51864
0 51866 7 1 2 86828 101944
0 51867 5 2 1 51866
0 51868 7 1 2 64403 103092
0 51869 7 1 2 102698 51868
0 51870 5 1 1 51869
0 51871 7 1 2 101821 101406
0 51872 5 1 1 51871
0 51873 7 1 2 69444 51872
0 51874 7 1 2 51870 51873
0 51875 5 1 1 51874
0 51876 7 1 2 102284 51875
0 51877 7 1 2 51865 51876
0 51878 5 1 1 51877
0 51879 7 1 2 51839 51878
0 51880 5 1 1 51879
0 51881 7 1 2 66177 51880
0 51882 5 1 1 51881
0 51883 7 1 2 101915 103091
0 51884 5 1 1 51883
0 51885 7 1 2 101928 103093
0 51886 5 1 1 51885
0 51887 7 1 2 51884 51886
0 51888 5 1 1 51887
0 51889 7 1 2 92965 103084
0 51890 7 1 2 51888 51889
0 51891 5 1 1 51890
0 51892 7 1 2 51882 51891
0 51893 5 1 1 51892
0 51894 7 1 2 70476 51893
0 51895 5 1 1 51894
0 51896 7 1 2 87774 97359
0 51897 5 1 1 51896
0 51898 7 1 2 87941 93883
0 51899 5 1 1 51898
0 51900 7 1 2 51897 51899
0 51901 5 1 1 51900
0 51902 7 1 2 101448 51901
0 51903 5 1 1 51902
0 51904 7 1 2 87942 101383
0 51905 5 1 1 51904
0 51906 7 1 2 51903 51905
0 51907 5 1 1 51906
0 51908 7 1 2 66046 51907
0 51909 5 1 1 51908
0 51910 7 1 2 99541 97479
0 51911 7 1 2 101449 51910
0 51912 5 1 1 51911
0 51913 7 1 2 51909 51912
0 51914 5 1 1 51913
0 51915 7 1 2 64594 51914
0 51916 5 1 1 51915
0 51917 7 1 2 93050 97558
0 51918 7 1 2 101335 51917
0 51919 5 1 1 51918
0 51920 7 1 2 64404 84741
0 51921 7 1 2 102701 51920
0 51922 5 1 1 51921
0 51923 7 1 2 51919 51922
0 51924 5 1 1 51923
0 51925 7 1 2 69445 51924
0 51926 5 1 1 51925
0 51927 7 1 2 51916 51926
0 51928 5 1 1 51927
0 51929 7 1 2 80585 97201
0 51930 7 1 2 51928 51929
0 51931 5 1 1 51930
0 51932 7 1 2 51895 51931
0 51933 5 1 1 51932
0 51934 7 1 2 69059 51933
0 51935 5 1 1 51934
0 51936 7 2 2 89002 101673
0 51937 7 2 2 67744 73656
0 51938 5 2 1 103096
0 51939 7 1 2 48398 103098
0 51940 5 1 1 51939
0 51941 7 1 2 64201 51940
0 51942 5 1 1 51941
0 51943 7 1 2 72665 86558
0 51944 7 1 2 86510 51943
0 51945 5 1 1 51944
0 51946 7 2 2 51942 51945
0 51947 5 1 1 103100
0 51948 7 1 2 87221 101575
0 51949 5 1 1 51948
0 51950 7 1 2 103101 51949
0 51951 5 1 1 51950
0 51952 7 1 2 103094 51951
0 51953 5 1 1 51952
0 51954 7 1 2 71372 99603
0 51955 5 1 1 51954
0 51956 7 1 2 85758 99668
0 51957 5 1 1 51956
0 51958 7 1 2 51955 51957
0 51959 5 1 1 51958
0 51960 7 1 2 70768 51959
0 51961 5 1 1 51960
0 51962 7 1 2 92407 99669
0 51963 5 1 1 51962
0 51964 7 1 2 51961 51963
0 51965 5 1 1 51964
0 51966 7 1 2 64202 51965
0 51967 5 1 1 51966
0 51968 7 2 2 76279 99670
0 51969 5 1 1 103102
0 51970 7 1 2 64003 99604
0 51971 5 1 1 51970
0 51972 7 1 2 51969 51971
0 51973 5 1 1 51972
0 51974 7 1 2 74189 51973
0 51975 5 1 1 51974
0 51976 7 1 2 65548 51975
0 51977 7 1 2 51967 51976
0 51978 5 1 1 51977
0 51979 7 1 2 99671 103077
0 51980 5 1 1 51979
0 51981 7 1 2 85771 99605
0 51982 5 1 1 51981
0 51983 7 1 2 51980 51982
0 51984 5 1 1 51983
0 51985 7 1 2 64203 51984
0 51986 5 1 1 51985
0 51987 7 1 2 92969 101352
0 51988 5 1 1 51987
0 51989 7 1 2 100307 51988
0 51990 5 1 1 51989
0 51991 7 1 2 73495 51990
0 51992 5 1 1 51991
0 51993 7 1 2 70477 51992
0 51994 7 1 2 51986 51993
0 51995 5 1 1 51994
0 51996 7 1 2 80998 51995
0 51997 7 1 2 51978 51996
0 51998 5 1 1 51997
0 51999 7 1 2 67903 92689
0 52000 5 1 1 51999
0 52001 7 1 2 100308 36840
0 52002 5 1 1 52001
0 52003 7 1 2 80999 52002
0 52004 5 1 1 52003
0 52005 7 1 2 52000 52004
0 52006 5 1 1 52005
0 52007 7 1 2 73084 52006
0 52008 5 1 1 52007
0 52009 7 1 2 82122 98478
0 52010 7 1 2 96873 52009
0 52011 5 1 1 52010
0 52012 7 1 2 52008 52011
0 52013 5 1 1 52012
0 52014 7 1 2 101576 52013
0 52015 5 1 1 52014
0 52016 7 1 2 77262 93059
0 52017 7 1 2 51947 52016
0 52018 5 1 1 52017
0 52019 7 1 2 52015 52018
0 52020 7 1 2 51998 52019
0 52021 5 1 1 52020
0 52022 7 1 2 66313 52021
0 52023 5 1 1 52022
0 52024 7 1 2 51953 52023
0 52025 5 1 1 52024
0 52026 7 1 2 102285 52025
0 52027 5 1 1 52026
0 52028 7 1 2 78720 92583
0 52029 7 1 2 92976 99398
0 52030 7 1 2 52028 52029
0 52031 7 1 2 102980 52030
0 52032 5 1 1 52031
0 52033 7 1 2 52027 52032
0 52034 5 1 1 52033
0 52035 7 1 2 99261 52034
0 52036 5 1 1 52035
0 52037 7 1 2 51935 52036
0 52038 7 1 2 51832 52037
0 52039 5 1 1 52038
0 52040 7 1 2 69146 52039
0 52041 5 1 1 52040
0 52042 7 3 2 70478 80539
0 52043 5 1 1 103104
0 52044 7 1 2 84040 52043
0 52045 5 2 1 52044
0 52046 7 1 2 102286 103107
0 52047 5 1 1 52046
0 52048 7 1 2 85283 102824
0 52049 7 1 2 97204 52048
0 52050 5 1 1 52049
0 52051 7 1 2 52047 52050
0 52052 5 1 1 52051
0 52053 7 1 2 98424 52052
0 52054 5 1 1 52053
0 52055 7 1 2 86781 87416
0 52056 5 1 1 52055
0 52057 7 3 2 70769 95412
0 52058 5 1 1 103109
0 52059 7 1 2 94897 103110
0 52060 5 1 1 52059
0 52061 7 1 2 52056 52060
0 52062 5 1 1 52061
0 52063 7 1 2 70479 52062
0 52064 5 1 1 52063
0 52065 7 1 2 7194 100421
0 52066 5 1 1 52065
0 52067 7 1 2 65866 52066
0 52068 5 1 1 52067
0 52069 7 2 2 87049 52068
0 52070 5 1 1 103112
0 52071 7 2 2 84645 103113
0 52072 5 1 1 103114
0 52073 7 1 2 86848 103115
0 52074 5 3 1 52073
0 52075 7 1 2 102295 103116
0 52076 5 1 1 52075
0 52077 7 1 2 94898 95134
0 52078 5 1 1 52077
0 52079 7 1 2 102277 52078
0 52080 5 1 1 52079
0 52081 7 1 2 78343 52080
0 52082 5 2 1 52081
0 52083 7 1 2 52076 103119
0 52084 7 1 2 52064 52083
0 52085 5 1 1 52084
0 52086 7 1 2 99767 52085
0 52087 5 1 1 52086
0 52088 7 1 2 52054 52087
0 52089 5 1 1 52088
0 52090 7 1 2 99724 52089
0 52091 5 1 1 52090
0 52092 7 1 2 96277 102028
0 52093 5 1 1 52092
0 52094 7 1 2 72711 102898
0 52095 5 1 1 52094
0 52096 7 1 2 96218 52095
0 52097 5 1 1 52096
0 52098 7 1 2 65549 52097
0 52099 5 1 1 52098
0 52100 7 1 2 75364 86715
0 52101 5 1 1 52100
0 52102 7 1 2 72874 52101
0 52103 7 1 2 52099 52102
0 52104 5 1 1 52103
0 52105 7 1 2 87417 52104
0 52106 5 1 1 52105
0 52107 7 1 2 52093 52106
0 52108 5 1 1 52107
0 52109 7 1 2 91377 103020
0 52110 7 1 2 52108 52109
0 52111 5 1 1 52110
0 52112 7 1 2 52091 52111
0 52113 5 1 1 52112
0 52114 7 1 2 100679 52113
0 52115 5 1 1 52114
0 52116 7 1 2 100006 100990
0 52117 5 1 1 52116
0 52118 7 1 2 84674 99494
0 52119 5 1 1 52118
0 52120 7 1 2 52117 52119
0 52121 5 1 1 52120
0 52122 7 1 2 70770 52121
0 52123 5 1 1 52122
0 52124 7 1 2 52123 103031
0 52125 5 1 1 52124
0 52126 7 1 2 64004 52125
0 52127 5 1 1 52126
0 52128 7 1 2 79396 99495
0 52129 5 1 1 52128
0 52130 7 1 2 52127 52129
0 52131 5 1 1 52130
0 52132 7 1 2 62669 52131
0 52133 5 1 1 52132
0 52134 7 1 2 74190 99496
0 52135 7 1 2 79571 52134
0 52136 5 1 1 52135
0 52137 7 1 2 52133 52136
0 52138 5 2 1 52137
0 52139 7 1 2 94899 103121
0 52140 5 1 1 52139
0 52141 7 1 2 100007 102287
0 52142 5 1 1 52141
0 52143 7 1 2 67745 78684
0 52144 7 1 2 83179 52143
0 52145 7 1 2 98174 52144
0 52146 5 1 1 52145
0 52147 7 1 2 52142 52146
0 52148 5 1 1 52147
0 52149 7 1 2 72201 52148
0 52150 5 1 1 52149
0 52151 7 1 2 99520 35349
0 52152 5 1 1 52151
0 52153 7 1 2 102288 52152
0 52154 5 1 1 52153
0 52155 7 1 2 70480 52154
0 52156 7 1 2 52150 52155
0 52157 7 1 2 52140 52156
0 52158 5 1 1 52157
0 52159 7 1 2 89123 99497
0 52160 5 1 1 52159
0 52161 7 1 2 92291 100721
0 52162 5 1 1 52161
0 52163 7 1 2 52160 52162
0 52164 5 1 1 52163
0 52165 7 1 2 71545 52164
0 52166 5 1 1 52165
0 52167 7 1 2 97575 100861
0 52168 5 1 1 52167
0 52169 7 1 2 52166 52168
0 52170 5 1 1 52169
0 52171 7 1 2 64204 52170
0 52172 5 1 1 52171
0 52173 7 1 2 72391 99498
0 52174 7 1 2 100456 52173
0 52175 5 1 1 52174
0 52176 7 1 2 98325 100056
0 52177 5 1 1 52176
0 52178 7 1 2 52175 52177
0 52179 7 1 2 52172 52178
0 52180 5 1 1 52179
0 52181 7 1 2 87418 52180
0 52182 5 1 1 52181
0 52183 7 1 2 86315 79141
0 52184 7 1 2 97776 52183
0 52185 7 1 2 85198 52184
0 52186 5 1 1 52185
0 52187 7 1 2 65550 52186
0 52188 7 1 2 52182 52187
0 52189 5 1 1 52188
0 52190 7 1 2 100650 52189
0 52191 7 1 2 52158 52190
0 52192 5 1 1 52191
0 52193 7 1 2 65551 52072
0 52194 5 1 1 52193
0 52195 7 1 2 72472 90422
0 52196 5 3 1 52195
0 52197 7 1 2 72202 93497
0 52198 5 2 1 52197
0 52199 7 1 2 103123 103126
0 52200 7 1 2 52194 52199
0 52201 5 2 1 52200
0 52202 7 1 2 87419 103128
0 52203 5 1 1 52202
0 52204 7 1 2 71763 82041
0 52205 5 1 1 52204
0 52206 7 1 2 103120 52205
0 52207 7 1 2 52203 52206
0 52208 5 1 1 52207
0 52209 7 1 2 100008 52208
0 52210 5 1 1 52209
0 52211 7 1 2 79627 103037
0 52212 5 1 1 52211
0 52213 7 1 2 62228 99499
0 52214 5 1 1 52213
0 52215 7 1 2 52212 52214
0 52216 5 1 1 52215
0 52217 7 1 2 94900 52216
0 52218 5 1 1 52217
0 52219 7 1 2 90755 99528
0 52220 7 1 2 5273 52219
0 52221 5 1 1 52220
0 52222 7 1 2 52218 52221
0 52223 5 1 1 52222
0 52224 7 1 2 72666 52223
0 52225 5 1 1 52224
0 52226 7 1 2 77138 96755
0 52227 5 1 1 52226
0 52228 7 1 2 90038 80061
0 52229 5 1 1 52228
0 52230 7 1 2 52227 52229
0 52231 5 1 1 52230
0 52232 7 1 2 62918 52231
0 52233 5 1 1 52232
0 52234 7 2 2 21577 100906
0 52235 5 1 1 103130
0 52236 7 1 2 65552 52235
0 52237 5 1 1 52236
0 52238 7 1 2 78218 85078
0 52239 5 2 1 52238
0 52240 7 1 2 52237 103132
0 52241 5 1 1 52240
0 52242 7 1 2 87420 52241
0 52243 5 1 1 52242
0 52244 7 1 2 52233 52243
0 52245 5 1 1 52244
0 52246 7 1 2 99500 52245
0 52247 5 1 1 52246
0 52248 7 1 2 52225 52247
0 52249 7 1 2 52210 52248
0 52250 5 1 1 52249
0 52251 7 1 2 87737 100662
0 52252 7 1 2 52250 52251
0 52253 5 1 1 52252
0 52254 7 1 2 52192 52253
0 52255 7 1 2 52115 52254
0 52256 5 1 1 52255
0 52257 7 1 2 64300 52256
0 52258 5 1 1 52257
0 52259 7 8 2 97996 100599
0 52260 7 1 2 78799 103134
0 52261 7 1 2 100991 52260
0 52262 5 1 1 52261
0 52263 7 3 2 64301 98113
0 52264 7 1 2 72586 82310
0 52265 7 1 2 93175 52264
0 52266 7 1 2 103142 52265
0 52267 5 1 1 52266
0 52268 7 1 2 52262 52267
0 52269 5 1 1 52268
0 52270 7 1 2 69446 52269
0 52271 5 1 1 52270
0 52272 7 1 2 102191 102306
0 52273 7 1 2 100680 52272
0 52274 7 1 2 100557 52273
0 52275 5 1 1 52274
0 52276 7 1 2 66314 52275
0 52277 7 1 2 52271 52276
0 52278 5 1 1 52277
0 52279 7 1 2 77263 101367
0 52280 5 1 1 52279
0 52281 7 1 2 83940 92561
0 52282 5 1 1 52281
0 52283 7 1 2 52280 52282
0 52284 5 2 1 52283
0 52285 7 1 2 91800 98224
0 52286 7 1 2 103145 52285
0 52287 5 1 1 52286
0 52288 7 1 2 66568 89003
0 52289 7 1 2 97997 98070
0 52290 7 1 2 52288 52289
0 52291 7 1 2 100558 52290
0 52292 5 1 1 52291
0 52293 7 1 2 61414 52292
0 52294 7 1 2 52287 52293
0 52295 5 1 1 52294
0 52296 7 1 2 87421 52295
0 52297 7 1 2 52278 52296
0 52298 5 1 1 52297
0 52299 7 2 2 98210 98625
0 52300 7 1 2 81360 103147
0 52301 7 1 2 101929 52300
0 52302 7 1 2 102954 52301
0 52303 5 1 1 52302
0 52304 7 1 2 52298 52303
0 52305 5 1 1 52304
0 52306 7 1 2 69257 52305
0 52307 5 1 1 52306
0 52308 7 3 2 95286 96859
0 52309 7 1 2 102289 103149
0 52310 7 1 2 102699 52309
0 52311 5 1 1 52310
0 52312 7 1 2 66178 52311
0 52313 7 1 2 52307 52312
0 52314 5 1 1 52313
0 52315 7 4 2 82703 98725
0 52316 7 1 2 103152 103150
0 52317 5 1 1 52316
0 52318 7 1 2 99701 97346
0 52319 5 1 1 52318
0 52320 7 1 2 103053 52319
0 52321 5 1 1 52320
0 52322 7 1 2 77264 52321
0 52323 5 1 1 52322
0 52324 7 1 2 62987 81000
0 52325 7 1 2 101368 52324
0 52326 5 1 1 52325
0 52327 7 1 2 52323 52326
0 52328 5 1 1 52327
0 52329 7 1 2 72766 95453
0 52330 7 1 2 52328 52329
0 52331 5 1 1 52330
0 52332 7 1 2 52317 52331
0 52333 5 1 1 52332
0 52334 7 1 2 87422 52333
0 52335 5 1 1 52334
0 52336 7 1 2 94901 102300
0 52337 7 1 2 103151 52336
0 52338 5 1 1 52337
0 52339 7 1 2 52335 52338
0 52340 5 1 1 52339
0 52341 7 1 2 66315 52340
0 52342 5 1 1 52341
0 52343 7 1 2 67824 103146
0 52344 5 1 1 52343
0 52345 7 1 2 99744 100600
0 52346 5 1 1 52345
0 52347 7 1 2 52344 52346
0 52348 5 1 1 52347
0 52349 7 1 2 92573 95449
0 52350 7 1 2 100718 52349
0 52351 7 1 2 95892 52350
0 52352 7 1 2 52348 52351
0 52353 5 1 1 52352
0 52354 7 1 2 61322 52353
0 52355 7 1 2 52342 52354
0 52356 5 1 1 52355
0 52357 7 1 2 73133 52356
0 52358 7 1 2 52314 52357
0 52359 5 1 1 52358
0 52360 7 1 2 52258 52359
0 52361 7 1 2 52041 52360
0 52362 7 1 2 51528 52361
0 52363 5 1 1 52362
0 52364 7 1 2 83165 52363
0 52365 5 1 1 52364
0 52366 7 1 2 103108 100074
0 52367 5 1 1 52366
0 52368 7 1 2 52058 100294
0 52369 5 3 1 52368
0 52370 7 1 2 65553 103156
0 52371 5 2 1 52370
0 52372 7 1 2 70481 103117
0 52373 5 1 1 52372
0 52374 7 1 2 103159 52373
0 52375 5 2 1 52374
0 52376 7 1 2 98984 103161
0 52377 5 1 1 52376
0 52378 7 1 2 52367 52377
0 52379 5 1 1 52378
0 52380 7 1 2 66179 52379
0 52381 5 1 1 52380
0 52382 7 1 2 86489 92182
0 52383 5 1 1 52382
0 52384 7 1 2 93618 52383
0 52385 5 1 1 52384
0 52386 7 1 2 70771 52385
0 52387 5 1 1 52386
0 52388 7 1 2 92183 103105
0 52389 5 1 1 52388
0 52390 7 1 2 52387 52389
0 52391 5 1 1 52390
0 52392 7 1 2 97722 52391
0 52393 5 1 1 52392
0 52394 7 1 2 52381 52393
0 52395 5 1 1 52394
0 52396 7 1 2 96171 52395
0 52397 5 1 1 52396
0 52398 7 1 2 65554 96336
0 52399 5 1 1 52398
0 52400 7 1 2 84390 86843
0 52401 5 1 1 52400
0 52402 7 1 2 83719 94134
0 52403 5 1 1 52402
0 52404 7 1 2 70482 52403
0 52405 7 1 2 52401 52404
0 52406 5 1 1 52405
0 52407 7 1 2 93048 102248
0 52408 7 1 2 52406 52407
0 52409 7 1 2 52399 52408
0 52410 5 1 1 52409
0 52411 7 1 2 52397 52410
0 52412 5 1 1 52411
0 52413 7 1 2 93832 52412
0 52414 5 1 1 52413
0 52415 7 1 2 75554 102876
0 52416 5 1 1 52415
0 52417 7 1 2 102874 52416
0 52418 5 2 1 52417
0 52419 7 1 2 62670 103163
0 52420 5 1 1 52419
0 52421 7 1 2 74990 92626
0 52422 5 1 1 52421
0 52423 7 1 2 52420 52422
0 52424 5 1 1 52423
0 52425 7 1 2 70772 52424
0 52426 5 1 1 52425
0 52427 7 1 2 92606 52426
0 52428 5 1 1 52427
0 52429 7 1 2 64005 52428
0 52430 5 1 1 52429
0 52431 7 1 2 92629 52430
0 52432 5 1 1 52431
0 52433 7 1 2 52432 98065
0 52434 5 1 1 52433
0 52435 7 1 2 82123 87237
0 52436 5 1 1 52435
0 52437 7 1 2 87339 52436
0 52438 5 2 1 52437
0 52439 7 1 2 97681 103165
0 52440 5 1 1 52439
0 52441 7 1 2 83963 74526
0 52442 5 1 1 52441
0 52443 7 1 2 88627 93672
0 52444 5 1 1 52443
0 52445 7 1 2 52442 52444
0 52446 5 1 1 52445
0 52447 7 1 2 62919 52446
0 52448 5 1 1 52447
0 52449 7 1 2 79381 80072
0 52450 7 1 2 88640 52449
0 52451 5 1 1 52450
0 52452 7 1 2 52448 52451
0 52453 5 1 1 52452
0 52454 7 1 2 65867 52453
0 52455 5 1 1 52454
0 52456 7 1 2 77286 79706
0 52457 5 1 1 52456
0 52458 7 1 2 91507 52457
0 52459 5 1 1 52458
0 52460 7 1 2 79700 98257
0 52461 5 1 1 52460
0 52462 7 1 2 35151 52461
0 52463 5 1 1 52462
0 52464 7 1 2 98326 52463
0 52465 5 1 1 52464
0 52466 7 1 2 52459 52465
0 52467 7 1 2 52455 52466
0 52468 5 1 1 52467
0 52469 7 1 2 52468 98025
0 52470 5 1 1 52469
0 52471 7 1 2 52440 52470
0 52472 5 1 1 52471
0 52473 7 1 2 70483 52472
0 52474 5 1 1 52473
0 52475 7 1 2 52434 52474
0 52476 5 1 1 52475
0 52477 7 1 2 66180 52476
0 52478 5 1 1 52477
0 52479 7 2 2 91014 99125
0 52480 7 1 2 103166 103167
0 52481 5 1 1 52480
0 52482 7 1 2 52478 52481
0 52483 5 1 1 52482
0 52484 7 1 2 69258 52483
0 52485 5 1 1 52484
0 52486 7 1 2 76280 98044
0 52487 7 1 2 92490 52486
0 52488 5 1 1 52487
0 52489 7 1 2 98662 52488
0 52490 5 1 1 52489
0 52491 7 1 2 78344 52490
0 52492 5 1 1 52491
0 52493 7 1 2 71373 85847
0 52494 5 3 1 52493
0 52495 7 1 2 73496 102992
0 52496 5 1 1 52495
0 52497 7 1 2 103169 52496
0 52498 5 3 1 52497
0 52499 7 1 2 70484 103172
0 52500 7 1 2 98671 52499
0 52501 5 1 1 52500
0 52502 7 1 2 52492 52501
0 52503 5 1 1 52502
0 52504 7 1 2 90274 52503
0 52505 5 1 1 52504
0 52506 7 3 2 99618 99221
0 52507 7 2 2 100128 103175
0 52508 5 1 1 103178
0 52509 7 2 2 97013 98672
0 52510 5 1 1 103180
0 52511 7 1 2 102664 103181
0 52512 5 1 1 52511
0 52513 7 1 2 52508 52512
0 52514 5 1 1 52513
0 52515 7 1 2 72667 52514
0 52516 5 1 1 52515
0 52517 7 2 2 65555 101396
0 52518 7 1 2 95287 102577
0 52519 7 1 2 103182 52518
0 52520 5 1 1 52519
0 52521 7 1 2 52516 52520
0 52522 7 1 2 52505 52521
0 52523 5 1 1 52522
0 52524 7 1 2 64405 52523
0 52525 5 1 1 52524
0 52526 7 1 2 52485 52525
0 52527 7 1 2 52414 52526
0 52528 5 1 1 52527
0 52529 7 1 2 90215 52528
0 52530 5 1 1 52529
0 52531 7 3 2 97405 101312
0 52532 7 1 2 70485 76393
0 52533 5 1 1 52532
0 52534 7 1 2 100874 52533
0 52535 5 1 1 52534
0 52536 7 1 2 96045 52535
0 52537 5 1 1 52536
0 52538 7 1 2 75533 90561
0 52539 5 1 1 52538
0 52540 7 1 2 78811 88641
0 52541 5 1 1 52540
0 52542 7 1 2 52539 52541
0 52543 5 1 1 52542
0 52544 7 1 2 64205 52543
0 52545 5 1 1 52544
0 52546 7 1 2 86995 73586
0 52547 5 2 1 52546
0 52548 7 1 2 66569 101280
0 52549 5 1 1 52548
0 52550 7 1 2 103187 52549
0 52551 5 1 1 52550
0 52552 7 1 2 69060 52551
0 52553 5 1 1 52552
0 52554 7 1 2 66047 82650
0 52555 5 1 1 52554
0 52556 7 1 2 52553 52555
0 52557 5 1 1 52556
0 52558 7 1 2 70773 52557
0 52559 5 1 1 52558
0 52560 7 1 2 52545 52559
0 52561 5 1 1 52560
0 52562 7 1 2 67535 52561
0 52563 5 1 1 52562
0 52564 7 1 2 86996 79407
0 52565 7 1 2 28299 52564
0 52566 5 1 1 52565
0 52567 7 1 2 52563 52566
0 52568 5 1 1 52567
0 52569 7 1 2 70486 52568
0 52570 5 1 1 52569
0 52571 7 1 2 52537 52570
0 52572 5 1 1 52571
0 52573 7 1 2 87796 52572
0 52574 5 1 1 52573
0 52575 7 2 2 73085 74991
0 52576 5 1 1 103189
0 52577 7 2 2 88470 92945
0 52578 5 1 1 103191
0 52579 7 1 2 103190 103192
0 52580 5 1 1 52579
0 52581 7 3 2 87687 92119
0 52582 7 1 2 62920 103193
0 52583 5 1 1 52582
0 52584 7 1 2 52578 52583
0 52585 5 1 1 52584
0 52586 7 1 2 71374 52585
0 52587 5 1 1 52586
0 52588 7 2 2 80734 87114
0 52589 5 1 1 103196
0 52590 7 1 2 87797 103197
0 52591 5 1 1 52590
0 52592 7 1 2 52587 52591
0 52593 5 1 1 52592
0 52594 7 1 2 70774 52593
0 52595 5 1 1 52594
0 52596 7 1 2 69259 94835
0 52597 7 1 2 102527 52596
0 52598 5 1 1 52597
0 52599 7 1 2 52595 52598
0 52600 5 1 1 52599
0 52601 7 1 2 65556 52600
0 52602 5 1 1 52601
0 52603 7 5 2 70487 87798
0 52604 7 2 2 73497 102678
0 52605 7 1 2 75747 103203
0 52606 5 1 1 52605
0 52607 7 1 2 99436 52606
0 52608 5 1 1 52607
0 52609 7 1 2 103198 52608
0 52610 5 1 1 52609
0 52611 7 1 2 52602 52610
0 52612 5 1 1 52611
0 52613 7 1 2 72668 52612
0 52614 5 1 1 52613
0 52615 7 1 2 52580 52614
0 52616 7 1 2 52574 52615
0 52617 5 1 1 52616
0 52618 7 1 2 103184 52617
0 52619 5 1 1 52618
0 52620 7 1 2 94738 98404
0 52621 7 1 2 97436 98631
0 52622 7 1 2 52620 52621
0 52623 7 1 2 98906 52622
0 52624 5 1 1 52623
0 52625 7 1 2 52619 52624
0 52626 5 1 1 52625
0 52627 7 1 2 99501 52626
0 52628 5 1 1 52627
0 52629 7 2 2 69447 96046
0 52630 7 1 2 66316 103205
0 52631 5 1 1 52630
0 52632 7 1 2 34833 52631
0 52633 5 1 1 52632
0 52634 7 1 2 94518 52633
0 52635 5 1 1 52634
0 52636 7 1 2 92201 100926
0 52637 5 1 1 52636
0 52638 7 1 2 86997 76281
0 52639 5 1 1 52638
0 52640 7 2 2 52589 52639
0 52641 5 1 1 103207
0 52642 7 1 2 71375 97059
0 52643 5 1 1 52642
0 52644 7 1 2 103208 52643
0 52645 5 1 1 52644
0 52646 7 1 2 100009 52645
0 52647 5 1 1 52646
0 52648 7 1 2 52637 52647
0 52649 7 1 2 52635 52648
0 52650 5 1 1 52649
0 52651 7 1 2 70775 52650
0 52652 5 1 1 52651
0 52653 7 2 2 72087 100010
0 52654 7 1 2 103209 52641
0 52655 5 1 1 52654
0 52656 7 1 2 52652 52655
0 52657 5 1 1 52656
0 52658 7 1 2 65557 52657
0 52659 5 1 1 52658
0 52660 7 2 2 70488 100011
0 52661 7 1 2 81960 103118
0 52662 5 1 1 52661
0 52663 7 1 2 86998 103173
0 52664 5 1 1 52663
0 52665 7 1 2 52662 52664
0 52666 5 1 1 52665
0 52667 7 1 2 103211 52666
0 52668 5 1 1 52667
0 52669 7 1 2 52659 52668
0 52670 5 1 1 52669
0 52671 7 1 2 98890 52670
0 52672 5 1 1 52671
0 52673 7 1 2 99395 49589
0 52674 5 2 1 52673
0 52675 7 1 2 70489 103213
0 52676 5 1 1 52675
0 52677 7 1 2 102882 52676
0 52678 5 1 1 52677
0 52679 7 1 2 100012 52678
0 52680 5 1 1 52679
0 52681 7 1 2 50170 52680
0 52682 5 1 1 52681
0 52683 7 1 2 97742 52682
0 52684 5 1 1 52683
0 52685 7 1 2 52672 52684
0 52686 5 1 1 52685
0 52687 7 1 2 99984 52686
0 52688 5 1 1 52687
0 52689 7 5 2 98549 99069
0 52690 7 1 2 72203 103199
0 52691 5 1 1 52690
0 52692 7 1 2 46807 52691
0 52693 5 1 1 52692
0 52694 7 1 2 100013 52693
0 52695 5 1 1 52694
0 52696 7 1 2 87738 101359
0 52697 5 1 1 52696
0 52698 7 1 2 52695 52697
0 52699 5 1 1 52698
0 52700 7 1 2 103215 52699
0 52701 5 1 1 52700
0 52702 7 1 2 75600 90797
0 52703 7 1 2 95649 52702
0 52704 7 1 2 91047 101332
0 52705 7 1 2 99632 52704
0 52706 7 1 2 52703 52705
0 52707 5 1 1 52706
0 52708 7 1 2 52701 52707
0 52709 5 1 1 52708
0 52710 7 1 2 87371 52709
0 52711 5 1 1 52710
0 52712 7 1 2 80554 103216
0 52713 5 1 1 52712
0 52714 7 1 2 95676 97565
0 52715 7 1 2 73134 52714
0 52716 7 1 2 100992 52715
0 52717 5 1 1 52716
0 52718 7 1 2 52713 52717
0 52719 5 1 1 52718
0 52720 7 1 2 87799 52719
0 52721 5 1 1 52720
0 52722 7 1 2 94384 102674
0 52723 7 1 2 103162 52722
0 52724 5 1 1 52723
0 52725 7 1 2 52721 52724
0 52726 5 1 1 52725
0 52727 7 1 2 81961 52726
0 52728 5 1 1 52727
0 52729 7 1 2 87800 102955
0 52730 5 1 1 52729
0 52731 7 2 2 64206 87739
0 52732 5 1 1 103220
0 52733 7 1 2 52730 52732
0 52734 5 1 1 52733
0 52735 7 1 2 73135 52734
0 52736 5 1 1 52735
0 52737 7 1 2 73498 101327
0 52738 5 1 1 52737
0 52739 7 1 2 64207 85449
0 52740 5 1 1 52739
0 52741 7 1 2 103170 52740
0 52742 7 1 2 52738 52741
0 52743 5 1 1 52742
0 52744 7 1 2 70490 52743
0 52745 5 1 1 52744
0 52746 7 1 2 62671 73781
0 52747 5 1 1 52746
0 52748 7 1 2 74193 52747
0 52749 7 1 2 78364 52748
0 52750 5 1 1 52749
0 52751 7 1 2 93295 52750
0 52752 5 1 1 52751
0 52753 7 1 2 52745 52752
0 52754 5 1 1 52753
0 52755 7 1 2 87740 52754
0 52756 5 1 1 52755
0 52757 7 1 2 52736 52756
0 52758 5 1 1 52757
0 52759 7 1 2 103185 52758
0 52760 5 1 1 52759
0 52761 7 1 2 84458 95546
0 52762 7 1 2 99037 52761
0 52763 7 1 2 98167 52762
0 52764 5 1 1 52763
0 52765 7 1 2 52760 52764
0 52766 5 1 1 52765
0 52767 7 1 2 86999 52766
0 52768 5 1 1 52767
0 52769 7 1 2 52728 52768
0 52770 5 1 1 52769
0 52771 7 1 2 100014 52770
0 52772 5 1 1 52771
0 52773 7 1 2 52711 52772
0 52774 7 1 2 52688 52773
0 52775 7 1 2 52628 52774
0 52776 7 1 2 52530 52775
0 52777 5 1 1 52776
0 52778 7 1 2 102258 52777
0 52779 5 1 1 52778
0 52780 7 5 2 94385 99756
0 52781 7 1 2 94521 103222
0 52782 5 1 1 52781
0 52783 7 3 2 69260 70967
0 52784 7 1 2 95643 99725
0 52785 7 1 2 103227 52784
0 52786 5 1 1 52785
0 52787 7 1 2 52782 52786
0 52788 5 1 1 52787
0 52789 7 1 2 73086 52788
0 52790 5 1 1 52789
0 52791 7 9 2 93919 99726
0 52792 7 1 2 103230 103106
0 52793 5 1 1 52792
0 52794 7 1 2 52790 52793
0 52795 5 1 1 52794
0 52796 7 1 2 67825 52795
0 52797 5 1 1 52796
0 52798 7 1 2 70491 100807
0 52799 5 1 1 52798
0 52800 7 1 2 51596 52799
0 52801 5 1 1 52800
0 52802 7 1 2 97654 52801
0 52803 5 1 1 52802
0 52804 7 1 2 52797 52803
0 52805 5 1 1 52804
0 52806 7 1 2 81962 52805
0 52807 5 1 1 52806
0 52808 7 1 2 78345 93609
0 52809 5 1 1 52808
0 52810 7 1 2 92184 95660
0 52811 5 1 1 52810
0 52812 7 1 2 52809 52811
0 52813 5 1 1 52812
0 52814 7 1 2 99207 97512
0 52815 7 1 2 52813 52814
0 52816 5 1 1 52815
0 52817 7 1 2 52807 52816
0 52818 5 1 1 52817
0 52819 7 1 2 61323 52818
0 52820 5 1 1 52819
0 52821 7 1 2 100702 102679
0 52822 5 1 1 52821
0 52823 7 1 2 100367 103206
0 52824 5 1 1 52823
0 52825 7 1 2 52822 52824
0 52826 5 1 1 52825
0 52827 7 1 2 67826 52826
0 52828 5 1 1 52827
0 52829 7 1 2 66317 97606
0 52830 7 1 2 100178 52829
0 52831 5 1 1 52830
0 52832 7 1 2 52828 52831
0 52833 5 1 1 52832
0 52834 7 1 2 71376 52833
0 52835 5 1 1 52834
0 52836 7 2 2 79382 91883
0 52837 7 1 2 103002 103239
0 52838 5 1 1 52837
0 52839 7 1 2 52835 52838
0 52840 5 1 1 52839
0 52841 7 1 2 70776 52840
0 52842 5 1 1 52841
0 52843 7 2 2 87000 100808
0 52844 7 1 2 101107 103241
0 52845 5 1 1 52844
0 52846 7 1 2 52842 52845
0 52847 5 1 1 52846
0 52848 7 1 2 72669 52847
0 52849 5 1 1 52848
0 52850 7 1 2 102682 36063
0 52851 5 1 1 52850
0 52852 7 1 2 100691 52851
0 52853 5 1 1 52852
0 52854 7 2 2 92815 96047
0 52855 7 1 2 102599 103243
0 52856 5 1 1 52855
0 52857 7 1 2 52853 52856
0 52858 5 1 1 52857
0 52859 7 1 2 62672 52858
0 52860 5 1 1 52859
0 52861 7 1 2 90869 96113
0 52862 7 1 2 99404 52861
0 52863 5 1 1 52862
0 52864 7 1 2 52860 52863
0 52865 5 1 1 52864
0 52866 7 1 2 78346 52865
0 52867 5 1 1 52866
0 52868 7 1 2 66318 103244
0 52869 5 1 1 52868
0 52870 7 1 2 102172 52869
0 52871 5 1 1 52870
0 52872 7 1 2 75651 52871
0 52873 5 1 1 52872
0 52874 7 1 2 52867 52873
0 52875 5 1 1 52874
0 52876 7 1 2 67827 52875
0 52877 5 1 1 52876
0 52878 7 1 2 84307 93636
0 52879 7 1 2 103240 52878
0 52880 5 1 1 52879
0 52881 7 1 2 52877 52880
0 52882 7 1 2 52849 52881
0 52883 5 1 1 52882
0 52884 7 1 2 69147 52883
0 52885 5 1 1 52884
0 52886 7 1 2 102583 99407
0 52887 7 1 2 101141 52886
0 52888 5 1 1 52887
0 52889 7 1 2 65558 52888
0 52890 7 1 2 52885 52889
0 52891 5 1 1 52890
0 52892 7 1 2 73953 102164
0 52893 5 1 1 52892
0 52894 7 1 2 17837 52893
0 52895 5 1 1 52894
0 52896 7 1 2 73499 52895
0 52897 5 1 1 52896
0 52898 7 3 2 65868 101652
0 52899 5 1 1 103245
0 52900 7 2 2 95866 52899
0 52901 5 1 1 103248
0 52902 7 1 2 81963 52901
0 52903 5 1 1 52902
0 52904 7 1 2 52897 52903
0 52905 5 1 1 52904
0 52906 7 1 2 64208 52905
0 52907 5 1 1 52906
0 52908 7 1 2 81964 103087
0 52909 5 1 1 52908
0 52910 7 1 2 52907 52909
0 52911 5 1 1 52910
0 52912 7 1 2 100692 52911
0 52913 5 1 1 52912
0 52914 7 1 2 90564 93404
0 52915 5 1 1 52914
0 52916 7 2 2 93137 99989
0 52917 7 1 2 52915 103250
0 52918 5 1 1 52917
0 52919 7 1 2 81965 97329
0 52920 5 1 1 52919
0 52921 7 1 2 61678 97238
0 52922 5 1 1 52921
0 52923 7 1 2 52920 52922
0 52924 5 1 1 52923
0 52925 7 1 2 100809 52924
0 52926 5 1 1 52925
0 52927 7 1 2 52918 52926
0 52928 5 1 1 52927
0 52929 7 1 2 66048 52928
0 52930 5 1 1 52929
0 52931 7 1 2 87410 91194
0 52932 5 1 1 52931
0 52933 7 1 2 61679 94660
0 52934 5 1 1 52933
0 52935 7 1 2 52932 52934
0 52936 5 1 1 52935
0 52937 7 1 2 100693 52936
0 52938 5 1 1 52937
0 52939 7 1 2 85885 87845
0 52940 7 1 2 103065 52939
0 52941 5 1 1 52940
0 52942 7 1 2 52938 52941
0 52943 5 1 1 52942
0 52944 7 1 2 70968 52943
0 52945 5 1 1 52944
0 52946 7 1 2 100694 103204
0 52947 5 1 1 52946
0 52948 7 1 2 86844 102174
0 52949 5 1 1 52948
0 52950 7 1 2 52947 52949
0 52951 7 1 2 52945 52950
0 52952 7 1 2 52930 52951
0 52953 5 1 1 52952
0 52954 7 1 2 69061 52953
0 52955 5 1 1 52954
0 52956 7 1 2 97343 35908
0 52957 5 1 1 52956
0 52958 7 1 2 64209 52957
0 52959 5 1 1 52958
0 52960 7 1 2 62673 96828
0 52961 5 1 1 52960
0 52962 7 1 2 52959 52961
0 52963 5 1 1 52962
0 52964 7 1 2 87001 52963
0 52965 5 1 1 52964
0 52966 7 1 2 23376 100435
0 52967 5 1 1 52966
0 52968 7 1 2 95602 52967
0 52969 5 1 1 52968
0 52970 7 1 2 85546 102680
0 52971 5 1 1 52970
0 52972 7 1 2 99437 52971
0 52973 5 1 1 52972
0 52974 7 1 2 72670 52973
0 52975 5 1 1 52974
0 52976 7 1 2 52969 52975
0 52977 7 1 2 52965 52976
0 52978 5 1 1 52977
0 52979 7 1 2 100810 52978
0 52980 5 1 1 52979
0 52981 7 1 2 52955 52980
0 52982 7 1 2 52913 52981
0 52983 5 1 1 52982
0 52984 7 1 2 97998 52983
0 52985 5 1 1 52984
0 52986 7 1 2 88170 94617
0 52987 7 1 2 103214 52986
0 52988 5 1 1 52987
0 52989 7 1 2 70492 52988
0 52990 7 1 2 52985 52989
0 52991 5 1 1 52990
0 52992 7 1 2 66181 52991
0 52993 7 1 2 52891 52992
0 52994 5 1 1 52993
0 52995 7 1 2 52820 52994
0 52996 5 1 1 52995
0 52997 7 1 2 102259 52996
0 52998 5 1 1 52997
0 52999 7 5 2 94386 97576
0 53000 7 1 2 95380 103252
0 53001 5 1 1 53000
0 53002 7 1 2 94775 99278
0 53003 7 1 2 98158 53002
0 53004 5 1 1 53003
0 53005 7 1 2 53001 53004
0 53006 5 1 1 53005
0 53007 7 1 2 62674 53006
0 53008 5 1 1 53007
0 53009 7 2 2 94618 99990
0 53010 5 1 1 103257
0 53011 7 1 2 76229 103258
0 53012 5 1 1 53011
0 53013 7 1 2 71027 87502
0 53014 7 1 2 103253 53013
0 53015 5 1 1 53014
0 53016 7 1 2 53012 53015
0 53017 5 1 1 53016
0 53018 7 1 2 66049 53017
0 53019 5 1 1 53018
0 53020 7 1 2 53008 53019
0 53021 5 1 1 53020
0 53022 7 1 2 69062 53021
0 53023 5 1 1 53022
0 53024 7 1 2 72473 103231
0 53025 5 1 1 53024
0 53026 7 1 2 65559 76287
0 53027 5 1 1 53026
0 53028 7 1 2 70969 86559
0 53029 7 1 2 103223 53028
0 53030 7 1 2 53027 53029
0 53031 5 1 1 53030
0 53032 7 1 2 53025 53031
0 53033 5 1 1 53032
0 53034 7 1 2 67066 53033
0 53035 5 1 1 53034
0 53036 7 1 2 53023 53035
0 53037 5 1 1 53036
0 53038 7 1 2 65245 53037
0 53039 5 1 1 53038
0 53040 7 2 2 84059 103254
0 53041 7 1 2 84593 91214
0 53042 7 1 2 103259 53041
0 53043 5 1 1 53042
0 53044 7 1 2 53039 53043
0 53045 5 1 1 53044
0 53046 7 1 2 69858 53045
0 53047 5 1 1 53046
0 53048 7 2 2 94407 97777
0 53049 7 1 2 73587 103261
0 53050 5 1 1 53049
0 53051 7 2 2 85759 73228
0 53052 7 1 2 103232 103263
0 53053 5 1 1 53052
0 53054 7 1 2 53050 53053
0 53055 5 1 1 53054
0 53056 7 1 2 69063 53055
0 53057 5 1 1 53056
0 53058 7 1 2 84989 103224
0 53059 5 1 1 53058
0 53060 7 1 2 53010 53059
0 53061 5 1 1 53060
0 53062 7 1 2 62229 53061
0 53063 5 1 1 53062
0 53064 7 1 2 53057 53063
0 53065 5 1 1 53064
0 53066 7 1 2 70493 53065
0 53067 5 1 1 53066
0 53068 7 1 2 92219 93585
0 53069 7 1 2 100030 53068
0 53070 7 1 2 86114 53069
0 53071 5 1 1 53070
0 53072 7 1 2 53067 53071
0 53073 5 1 1 53072
0 53074 7 1 2 78559 53073
0 53075 5 1 1 53074
0 53076 7 1 2 88384 103255
0 53077 5 1 1 53076
0 53078 7 1 2 99727 99314
0 53079 7 1 2 103246 53078
0 53080 5 1 1 53079
0 53081 7 1 2 53077 53080
0 53082 5 1 1 53081
0 53083 7 1 2 62675 53082
0 53084 5 1 1 53083
0 53085 7 1 2 103027 99321
0 53086 5 1 1 53085
0 53087 7 1 2 53084 53086
0 53088 5 1 1 53087
0 53089 7 1 2 78616 53088
0 53090 5 1 1 53089
0 53091 7 1 2 93920 98647
0 53092 7 1 2 100125 53091
0 53093 7 1 2 89215 53092
0 53094 5 1 1 53093
0 53095 7 1 2 53090 53094
0 53096 5 1 1 53095
0 53097 7 1 2 65560 53096
0 53098 5 1 1 53097
0 53099 7 1 2 65561 75555
0 53100 7 1 2 103262 53099
0 53101 5 1 1 53100
0 53102 7 1 2 73614 103233
0 53103 7 1 2 100538 53102
0 53104 5 1 1 53103
0 53105 7 1 2 53101 53104
0 53106 5 1 1 53105
0 53107 7 1 2 78560 53106
0 53108 5 1 1 53107
0 53109 7 1 2 84022 103234
0 53110 5 1 1 53109
0 53111 7 1 2 94408 101986
0 53112 5 1 1 53111
0 53113 7 1 2 53110 53112
0 53114 5 1 1 53113
0 53115 7 1 2 78631 53114
0 53116 5 1 1 53115
0 53117 7 1 2 53108 53116
0 53118 5 1 1 53117
0 53119 7 1 2 70777 53118
0 53120 5 1 1 53119
0 53121 7 3 2 70494 84990
0 53122 7 1 2 101961 103256
0 53123 7 1 2 103265 53122
0 53124 5 1 1 53123
0 53125 7 1 2 53120 53124
0 53126 7 1 2 53098 53125
0 53127 5 1 1 53126
0 53128 7 1 2 64210 53127
0 53129 5 1 1 53128
0 53130 7 1 2 53075 53129
0 53131 7 1 2 53047 53130
0 53132 5 1 1 53131
0 53133 7 1 2 87002 53132
0 53134 5 1 1 53133
0 53135 7 2 2 73743 91749
0 53136 5 1 1 103268
0 53137 7 1 2 76962 96711
0 53138 5 2 1 53137
0 53139 7 1 2 67067 103270
0 53140 5 1 1 53139
0 53141 7 1 2 53136 53140
0 53142 5 2 1 53141
0 53143 7 1 2 69859 103272
0 53144 5 1 1 53143
0 53145 7 1 2 102774 53144
0 53146 5 1 1 53145
0 53147 7 1 2 73500 53146
0 53148 5 1 1 53147
0 53149 7 1 2 73744 89813
0 53150 7 1 2 97385 53149
0 53151 5 1 1 53150
0 53152 7 1 2 53148 53151
0 53153 5 1 1 53152
0 53154 7 1 2 103225 53153
0 53155 5 1 1 53154
0 53156 7 1 2 66319 102771
0 53157 7 1 2 98838 53156
0 53158 5 1 1 53157
0 53159 7 1 2 78561 80387
0 53160 5 2 1 53159
0 53161 7 1 2 76725 87162
0 53162 5 1 1 53161
0 53163 7 1 2 103274 53162
0 53164 5 4 1 53163
0 53165 7 1 2 91393 100833
0 53166 7 1 2 103276 53165
0 53167 5 1 1 53166
0 53168 7 1 2 53158 53167
0 53169 5 1 1 53168
0 53170 7 1 2 98327 53169
0 53171 5 1 1 53170
0 53172 7 1 2 93676 103277
0 53173 5 1 1 53172
0 53174 7 1 2 85881 86416
0 53175 7 1 2 73136 53174
0 53176 5 1 1 53175
0 53177 7 1 2 53173 53176
0 53178 5 1 1 53177
0 53179 7 1 2 103235 53178
0 53180 5 1 1 53179
0 53181 7 1 2 86335 103260
0 53182 5 1 1 53181
0 53183 7 1 2 53180 53182
0 53184 5 1 1 53183
0 53185 7 1 2 67746 53184
0 53186 5 1 1 53185
0 53187 7 1 2 53171 53186
0 53188 7 1 2 53155 53187
0 53189 5 1 1 53188
0 53190 7 1 2 81966 53189
0 53191 5 1 1 53190
0 53192 7 1 2 53134 53191
0 53193 5 1 1 53192
0 53194 7 1 2 93884 53193
0 53195 5 1 1 53194
0 53196 7 1 2 72088 102170
0 53197 5 1 1 53196
0 53198 7 1 2 70495 103242
0 53199 5 1 1 53198
0 53200 7 1 2 53197 53199
0 53201 5 1 1 53200
0 53202 7 1 2 67068 53201
0 53203 5 1 1 53202
0 53204 7 2 2 72587 100703
0 53205 5 1 1 103280
0 53206 7 1 2 36967 36673
0 53207 5 1 1 53206
0 53208 7 1 2 72204 53207
0 53209 5 1 1 53208
0 53210 7 1 2 53205 53209
0 53211 5 1 1 53210
0 53212 7 1 2 67536 53211
0 53213 5 1 1 53212
0 53214 7 1 2 84665 100695
0 53215 5 2 1 53214
0 53216 7 1 2 53213 103282
0 53217 5 1 1 53216
0 53218 7 1 2 68877 53217
0 53219 5 1 1 53218
0 53220 7 1 2 72733 100696
0 53221 5 1 1 53220
0 53222 7 1 2 53219 53221
0 53223 5 1 1 53222
0 53224 7 1 2 72474 53223
0 53225 5 1 1 53224
0 53226 7 1 2 96205 100811
0 53227 5 1 1 53226
0 53228 7 1 2 97102 100824
0 53229 5 1 1 53228
0 53230 7 1 2 53227 53229
0 53231 5 1 1 53230
0 53232 7 1 2 65869 53231
0 53233 5 1 1 53232
0 53234 7 1 2 97117 100697
0 53235 5 1 1 53234
0 53236 7 1 2 82447 101692
0 53237 5 1 1 53236
0 53238 7 1 2 97270 100812
0 53239 5 1 1 53238
0 53240 7 1 2 53237 53239
0 53241 5 1 1 53240
0 53242 7 1 2 98328 53241
0 53243 5 1 1 53242
0 53244 7 1 2 75295 100794
0 53245 7 1 2 96804 53244
0 53246 5 1 1 53245
0 53247 7 1 2 53243 53246
0 53248 7 1 2 53235 53247
0 53249 7 1 2 53233 53248
0 53250 5 1 1 53249
0 53251 7 1 2 65562 53250
0 53252 5 1 1 53251
0 53253 7 1 2 53225 53252
0 53254 5 1 1 53253
0 53255 7 1 2 87372 53254
0 53256 5 1 1 53255
0 53257 7 1 2 53203 53256
0 53258 5 1 1 53257
0 53259 7 1 2 78617 53258
0 53260 5 1 1 53259
0 53261 7 1 2 79628 100698
0 53262 5 1 1 53261
0 53263 7 1 2 62230 100704
0 53264 5 1 1 53263
0 53265 7 1 2 53262 53264
0 53266 5 1 1 53265
0 53267 7 1 2 62921 53266
0 53268 5 1 1 53267
0 53269 7 2 2 73358 100813
0 53270 5 1 1 103284
0 53271 7 1 2 71747 103285
0 53272 5 1 1 53271
0 53273 7 1 2 53268 53272
0 53274 5 1 1 53273
0 53275 7 1 2 87003 53274
0 53276 5 1 1 53275
0 53277 7 1 2 76282 100825
0 53278 5 1 1 53277
0 53279 7 1 2 53270 53278
0 53280 5 1 1 53279
0 53281 7 1 2 102866 53280
0 53282 5 1 1 53281
0 53283 7 1 2 53276 53282
0 53284 5 1 1 53283
0 53285 7 1 2 72671 53284
0 53286 5 1 1 53285
0 53287 7 1 2 36631 51666
0 53288 5 1 1 53287
0 53289 7 2 2 87373 53288
0 53290 7 1 2 86553 103286
0 53291 5 1 1 53290
0 53292 7 1 2 97001 100705
0 53293 5 1 1 53292
0 53294 7 1 2 53291 53293
0 53295 5 1 1 53294
0 53296 7 1 2 78347 53295
0 53297 5 1 1 53296
0 53298 7 1 2 92202 97162
0 53299 5 1 1 53298
0 53300 7 1 2 77953 75736
0 53301 7 1 2 103287 53300
0 53302 5 1 1 53301
0 53303 7 1 2 53299 53302
0 53304 5 1 1 53303
0 53305 7 1 2 70970 53304
0 53306 5 1 1 53305
0 53307 7 1 2 53297 53306
0 53308 7 1 2 53286 53307
0 53309 5 1 1 53308
0 53310 7 1 2 78562 53309
0 53311 5 1 1 53310
0 53312 7 1 2 53260 53311
0 53313 5 1 1 53312
0 53314 7 1 2 96975 53313
0 53315 5 1 1 53314
0 53316 7 1 2 66320 101153
0 53317 5 1 1 53316
0 53318 7 1 2 103283 53317
0 53319 5 1 1 53318
0 53320 7 1 2 87374 53319
0 53321 5 1 1 53320
0 53322 7 1 2 92203 95669
0 53323 7 1 2 96642 53322
0 53324 5 1 1 53323
0 53325 7 1 2 53321 53324
0 53326 5 1 1 53325
0 53327 7 1 2 80586 53326
0 53328 5 1 1 53327
0 53329 7 1 2 85729 87860
0 53330 7 1 2 99208 53329
0 53331 7 1 2 90415 53330
0 53332 5 1 1 53331
0 53333 7 1 2 53328 53332
0 53334 5 1 1 53333
0 53335 7 1 2 67537 53334
0 53336 5 1 1 53335
0 53337 7 3 2 87375 80587
0 53338 7 1 2 75910 103251
0 53339 7 1 2 103288 53338
0 53340 5 1 1 53339
0 53341 7 1 2 53336 53340
0 53342 5 1 1 53341
0 53343 7 1 2 76726 53342
0 53344 5 1 1 53343
0 53345 7 1 2 79758 90246
0 53346 7 1 2 100826 53345
0 53347 7 1 2 97281 53346
0 53348 5 1 1 53347
0 53349 7 1 2 53344 53348
0 53350 5 1 1 53349
0 53351 7 1 2 92651 102449
0 53352 7 1 2 53350 53351
0 53353 5 1 1 53352
0 53354 7 1 2 53315 53353
0 53355 7 1 2 53195 53354
0 53356 7 1 2 52998 53355
0 53357 5 1 1 53356
0 53358 7 1 2 98399 53357
0 53359 5 1 1 53358
0 53360 7 3 2 89734 86439
0 53361 7 1 2 62231 103291
0 53362 5 1 1 53361
0 53363 7 2 2 70778 102956
0 53364 7 1 2 73615 103294
0 53365 5 1 1 53364
0 53366 7 1 2 53362 53365
0 53367 5 2 1 53366
0 53368 7 1 2 87801 103296
0 53369 5 1 1 53368
0 53370 7 2 2 70496 103157
0 53371 5 1 1 103298
0 53372 7 1 2 87741 103299
0 53373 5 1 1 53372
0 53374 7 1 2 53369 53373
0 53375 5 1 1 53374
0 53376 7 1 2 78563 53375
0 53377 5 1 1 53376
0 53378 7 1 2 76231 19511
0 53379 5 1 1 53378
0 53380 7 1 2 67747 53379
0 53381 5 1 1 53380
0 53382 7 1 2 72926 72378
0 53383 7 1 2 100880 53382
0 53384 5 1 1 53383
0 53385 7 2 2 53381 53384
0 53386 5 1 1 103300
0 53387 7 1 2 67069 80555
0 53388 5 2 1 53387
0 53389 7 1 2 103301 103302
0 53390 5 2 1 53389
0 53391 7 1 2 87802 103304
0 53392 5 1 1 53391
0 53393 7 1 2 87742 103129
0 53394 5 1 1 53393
0 53395 7 1 2 53392 53394
0 53396 5 1 1 53395
0 53397 7 1 2 78618 53396
0 53398 5 1 1 53397
0 53399 7 1 2 53377 53398
0 53400 5 1 1 53399
0 53401 7 1 2 90275 53400
0 53402 5 1 1 53401
0 53403 7 1 2 75901 100930
0 53404 5 3 1 53403
0 53405 7 1 2 96219 103306
0 53406 5 2 1 53405
0 53407 7 1 2 87803 103309
0 53408 5 1 1 53407
0 53409 7 1 2 89952 96664
0 53410 7 1 2 103131 53409
0 53411 5 1 1 53410
0 53412 7 1 2 87743 53411
0 53413 5 1 1 53412
0 53414 7 1 2 53408 53413
0 53415 5 1 1 53414
0 53416 7 1 2 65563 53415
0 53417 5 1 1 53416
0 53418 7 1 2 71022 87775
0 53419 5 1 1 53418
0 53420 7 1 2 29757 53419
0 53421 5 1 1 53420
0 53422 7 1 2 69064 53421
0 53423 5 1 1 53422
0 53424 7 3 2 66050 93026
0 53425 7 1 2 72712 103311
0 53426 5 1 1 53425
0 53427 7 1 2 53423 53426
0 53428 5 1 1 53427
0 53429 7 1 2 72475 53428
0 53430 5 1 1 53429
0 53431 7 1 2 53417 53430
0 53432 5 1 1 53431
0 53433 7 1 2 78619 53432
0 53434 5 1 1 53433
0 53435 7 1 2 87765 7914
0 53436 5 1 1 53435
0 53437 7 1 2 72672 53436
0 53438 5 1 1 53437
0 53439 7 1 2 89640 87804
0 53440 5 1 1 53439
0 53441 7 1 2 53438 53440
0 53442 5 1 1 53441
0 53443 7 1 2 62676 53442
0 53444 5 1 1 53443
0 53445 7 1 2 87744 92403
0 53446 5 1 1 53445
0 53447 7 1 2 87745 94489
0 53448 5 1 1 53447
0 53449 7 1 2 103228 102528
0 53450 5 1 1 53449
0 53451 7 1 2 53448 53450
0 53452 5 1 1 53451
0 53453 7 1 2 64211 53452
0 53454 5 1 1 53453
0 53455 7 1 2 53446 53454
0 53456 7 1 2 53444 53455
0 53457 5 1 1 53456
0 53458 7 1 2 70779 53457
0 53459 5 1 1 53458
0 53460 7 1 2 87805 93235
0 53461 5 1 1 53460
0 53462 7 1 2 53459 53461
0 53463 5 1 1 53462
0 53464 7 1 2 86291 53463
0 53465 5 1 1 53464
0 53466 7 1 2 53434 53465
0 53467 5 1 1 53466
0 53468 7 1 2 83964 53467
0 53469 5 1 1 53468
0 53470 7 1 2 53402 53469
0 53471 5 1 1 53470
0 53472 7 1 2 99145 53471
0 53473 5 1 1 53472
0 53474 7 2 2 82998 92946
0 53475 7 1 2 70497 97516
0 53476 5 3 1 53475
0 53477 7 1 2 65564 103310
0 53478 5 2 1 53477
0 53479 7 1 2 103316 103319
0 53480 5 1 1 53479
0 53481 7 1 2 78620 53480
0 53482 5 1 1 53481
0 53483 7 1 2 62922 86554
0 53484 5 1 1 53483
0 53485 7 1 2 67070 53484
0 53486 5 1 1 53485
0 53487 7 1 2 78348 53486
0 53488 5 1 1 53487
0 53489 7 1 2 72807 74209
0 53490 5 1 1 53489
0 53491 7 1 2 75240 85163
0 53492 5 1 1 53491
0 53493 7 1 2 72673 53492
0 53494 5 1 1 53493
0 53495 7 1 2 53490 53494
0 53496 7 1 2 53488 53495
0 53497 5 1 1 53496
0 53498 7 1 2 78564 53497
0 53499 5 1 1 53498
0 53500 7 1 2 53482 53499
0 53501 5 1 1 53500
0 53502 7 1 2 103314 53501
0 53503 5 1 1 53502
0 53504 7 2 2 84885 102825
0 53505 7 3 2 73359 103321
0 53506 5 1 1 103323
0 53507 7 1 2 86292 103324
0 53508 5 1 1 53507
0 53509 7 2 2 65246 53386
0 53510 7 1 2 69860 103326
0 53511 5 1 1 53510
0 53512 7 1 2 53508 53511
0 53513 5 1 1 53512
0 53514 7 2 2 69636 53513
0 53515 7 1 2 100935 103328
0 53516 5 1 1 53515
0 53517 7 1 2 53503 53516
0 53518 5 1 1 53517
0 53519 7 1 2 93921 53518
0 53520 5 1 1 53519
0 53521 7 3 2 97637 102646
0 53522 7 1 2 77097 94526
0 53523 5 1 1 53522
0 53524 7 1 2 6607 53523
0 53525 5 1 1 53524
0 53526 7 1 2 65565 53525
0 53527 5 1 1 53526
0 53528 7 1 2 77098 83879
0 53529 5 1 1 53528
0 53530 7 1 2 53527 53529
0 53531 5 1 1 53530
0 53532 7 1 2 103330 53531
0 53533 5 1 1 53532
0 53534 7 1 2 11824 53371
0 53535 5 1 1 53534
0 53536 7 3 2 96172 97723
0 53537 7 1 2 65002 103333
0 53538 7 1 2 53535 53537
0 53539 5 1 1 53538
0 53540 7 1 2 53533 53539
0 53541 5 1 1 53540
0 53542 7 1 2 70156 53541
0 53543 5 1 1 53542
0 53544 7 1 2 65566 52070
0 53545 5 1 1 53544
0 53546 7 1 2 103124 53545
0 53547 5 1 1 53546
0 53548 7 1 2 103334 53547
0 53549 5 1 1 53548
0 53550 7 1 2 78225 35751
0 53551 5 2 1 53550
0 53552 7 1 2 71377 103336
0 53553 5 2 1 53552
0 53554 7 1 2 64212 84991
0 53555 5 2 1 53554
0 53556 7 1 2 89953 94500
0 53557 7 1 2 103340 53556
0 53558 5 1 1 53557
0 53559 7 1 2 70498 53558
0 53560 5 1 1 53559
0 53561 7 1 2 103338 53560
0 53562 5 1 1 53561
0 53563 7 1 2 103331 53562
0 53564 5 1 1 53563
0 53565 7 1 2 61324 86316
0 53566 7 1 2 80247 99797
0 53567 7 1 2 53565 53566
0 53568 5 1 1 53567
0 53569 7 1 2 53564 53568
0 53570 5 1 1 53569
0 53571 7 1 2 67071 53570
0 53572 5 1 1 53571
0 53573 7 1 2 90434 103332
0 53574 5 1 1 53573
0 53575 7 1 2 91324 78782
0 53576 7 1 2 97724 53575
0 53577 7 1 2 101878 53576
0 53578 5 1 1 53577
0 53579 7 1 2 53574 53578
0 53580 5 1 1 53579
0 53581 7 1 2 70780 53580
0 53582 5 1 1 53581
0 53583 7 1 2 53572 53582
0 53584 7 1 2 53549 53583
0 53585 5 1 1 53584
0 53586 7 1 2 78621 53585
0 53587 5 1 1 53586
0 53588 7 1 2 53543 53587
0 53589 5 1 1 53588
0 53590 7 1 2 64406 53589
0 53591 5 1 1 53590
0 53592 7 2 2 64407 82097
0 53593 7 1 2 96724 99960
0 53594 7 1 2 103342 53593
0 53595 5 1 1 53594
0 53596 7 1 2 91999 100743
0 53597 7 1 2 97240 53596
0 53598 5 1 1 53597
0 53599 7 1 2 53595 53598
0 53600 5 1 1 53599
0 53601 7 1 2 70499 53600
0 53602 5 1 1 53601
0 53603 7 2 2 97725 103070
0 53604 7 1 2 102127 103344
0 53605 7 1 2 100709 53604
0 53606 5 1 1 53605
0 53607 7 1 2 53602 53606
0 53608 5 1 1 53607
0 53609 7 1 2 72205 53608
0 53610 5 1 1 53609
0 53611 7 1 2 53591 53610
0 53612 7 1 2 53520 53611
0 53613 5 1 1 53612
0 53614 7 1 2 93833 53613
0 53615 5 1 1 53614
0 53616 7 1 2 53473 53615
0 53617 5 1 1 53616
0 53618 7 1 2 62988 53617
0 53619 5 1 1 53618
0 53620 7 1 2 95098 103327
0 53621 5 1 1 53620
0 53622 7 1 2 5616 96712
0 53623 5 3 1 53622
0 53624 7 1 2 73501 103346
0 53625 5 1 1 53624
0 53626 7 1 2 78226 23928
0 53627 5 1 1 53626
0 53628 7 1 2 62923 53627
0 53629 5 1 1 53628
0 53630 7 1 2 64213 103266
0 53631 5 1 1 53630
0 53632 7 1 2 53629 53631
0 53633 7 1 2 103339 53632
0 53634 5 1 1 53633
0 53635 7 1 2 65247 53634
0 53636 5 1 1 53635
0 53637 7 1 2 53625 53636
0 53638 5 1 1 53637
0 53639 7 1 2 82704 94858
0 53640 7 1 2 53638 53639
0 53641 5 1 1 53640
0 53642 7 1 2 53621 53641
0 53643 5 1 1 53642
0 53644 7 1 2 69861 53643
0 53645 5 1 1 53644
0 53646 7 1 2 95099 103325
0 53647 5 1 1 53646
0 53648 7 2 2 79272 94409
0 53649 7 1 2 94961 103349
0 53650 5 1 1 53649
0 53651 7 1 2 53647 53650
0 53652 5 1 1 53651
0 53653 7 1 2 70500 53652
0 53654 5 1 1 53653
0 53655 7 1 2 64808 103350
0 53656 7 1 2 102656 53655
0 53657 5 1 1 53656
0 53658 7 1 2 53654 53657
0 53659 5 1 1 53658
0 53660 7 1 2 78565 53659
0 53661 5 1 1 53660
0 53662 7 1 2 53645 53661
0 53663 5 1 1 53662
0 53664 7 1 2 61325 53663
0 53665 5 1 1 53664
0 53666 7 1 2 72206 97241
0 53667 5 1 1 53666
0 53668 7 1 2 27200 53667
0 53669 5 1 1 53668
0 53670 7 1 2 68878 53669
0 53671 5 1 1 53670
0 53672 7 1 2 80797 88471
0 53673 7 1 2 89554 53672
0 53674 5 1 1 53673
0 53675 7 1 2 53671 53674
0 53676 5 1 1 53675
0 53677 7 1 2 103068 53676
0 53678 5 1 1 53677
0 53679 7 1 2 90140 96107
0 53680 7 1 2 102981 53679
0 53681 5 1 1 53680
0 53682 7 1 2 53678 53681
0 53683 5 1 1 53682
0 53684 7 1 2 97638 97446
0 53685 7 1 2 53683 53684
0 53686 5 1 1 53685
0 53687 7 1 2 53665 53686
0 53688 5 1 1 53687
0 53689 7 1 2 93834 53688
0 53690 5 1 1 53689
0 53691 7 1 2 70971 86326
0 53692 5 1 1 53691
0 53693 7 1 2 78634 53692
0 53694 5 1 1 53693
0 53695 7 1 2 85295 53694
0 53696 5 1 1 53695
0 53697 7 1 2 71378 77530
0 53698 5 1 1 53697
0 53699 7 1 2 96665 53698
0 53700 5 1 1 53699
0 53701 7 1 2 100186 53700
0 53702 5 1 1 53701
0 53703 7 1 2 53696 53702
0 53704 5 1 1 53703
0 53705 7 1 2 70501 53704
0 53706 5 1 1 53705
0 53707 7 1 2 88146 92323
0 53708 7 1 2 102982 53707
0 53709 5 1 1 53708
0 53710 7 1 2 53706 53709
0 53711 5 1 1 53710
0 53712 7 1 2 83965 53711
0 53713 5 1 1 53712
0 53714 7 1 2 90363 87507
0 53715 5 1 1 53714
0 53716 7 2 2 76580 77322
0 53717 7 1 2 84184 83853
0 53718 7 1 2 103351 53717
0 53719 5 1 1 53718
0 53720 7 1 2 53715 53719
0 53721 5 1 1 53720
0 53722 7 1 2 62924 53721
0 53723 5 1 1 53722
0 53724 7 1 2 90423 80588
0 53725 5 1 1 53724
0 53726 7 1 2 77667 86243
0 53727 5 1 1 53726
0 53728 7 1 2 53725 53727
0 53729 5 1 1 53728
0 53730 7 1 2 88147 100915
0 53731 7 1 2 53729 53730
0 53732 5 1 1 53731
0 53733 7 1 2 53723 53732
0 53734 7 1 2 53713 53733
0 53735 5 1 1 53734
0 53736 7 1 2 87746 53735
0 53737 5 1 1 53736
0 53738 7 1 2 90555 83979
0 53739 5 1 1 53738
0 53740 7 1 2 83966 89524
0 53741 5 1 1 53740
0 53742 7 1 2 53739 53741
0 53743 5 1 1 53742
0 53744 7 2 2 97447 97547
0 53745 7 1 2 80589 103353
0 53746 7 1 2 53743 53745
0 53747 5 1 1 53746
0 53748 7 1 2 53737 53747
0 53749 5 1 1 53748
0 53750 7 1 2 99258 53749
0 53751 5 1 1 53750
0 53752 7 1 2 53690 53751
0 53753 5 1 1 53752
0 53754 7 1 2 67828 53753
0 53755 5 1 1 53754
0 53756 7 2 2 85497 91508
0 53757 5 1 1 103355
0 53758 7 1 2 103356 98938
0 53759 5 1 1 53758
0 53760 7 1 2 61680 89445
0 53761 5 1 1 53760
0 53762 7 1 2 15693 53761
0 53763 5 1 1 53762
0 53764 7 1 2 87934 99907
0 53765 7 1 2 53763 53764
0 53766 5 1 1 53765
0 53767 7 1 2 53759 53766
0 53768 5 1 1 53767
0 53769 7 1 2 65248 53768
0 53770 5 1 1 53769
0 53771 7 1 2 81674 89537
0 53772 5 1 1 53771
0 53773 7 1 2 53757 53772
0 53774 5 1 1 53773
0 53775 7 1 2 77668 98891
0 53776 7 1 2 53774 53775
0 53777 5 1 1 53776
0 53778 7 1 2 53770 53777
0 53779 5 1 1 53778
0 53780 7 1 2 65870 53779
0 53781 5 1 1 53780
0 53782 7 2 2 100640 97726
0 53783 7 1 2 75902 103357
0 53784 7 1 2 101282 53783
0 53785 5 1 1 53784
0 53786 7 1 2 53781 53785
0 53787 5 1 1 53786
0 53788 7 1 2 65567 53787
0 53789 5 1 1 53788
0 53790 7 1 2 95562 98927
0 53791 5 1 1 53790
0 53792 7 1 2 66570 93248
0 53793 5 1 1 53792
0 53794 7 1 2 12523 53793
0 53795 5 1 1 53794
0 53796 7 1 2 79505 97616
0 53797 7 1 2 53795 53796
0 53798 5 1 1 53797
0 53799 7 1 2 53791 53798
0 53800 5 1 1 53799
0 53801 7 1 2 76950 53800
0 53802 5 1 1 53801
0 53803 7 1 2 53789 53802
0 53804 5 1 1 53803
0 53805 7 1 2 69065 53804
0 53806 5 1 1 53805
0 53807 7 1 2 100048 101292
0 53808 5 1 1 53807
0 53809 7 1 2 67072 100044
0 53810 5 1 1 53809
0 53811 7 1 2 53808 53810
0 53812 5 1 1 53811
0 53813 7 1 2 70502 53812
0 53814 5 1 1 53813
0 53815 7 3 2 96436 97727
0 53816 7 1 2 71546 100559
0 53817 5 1 1 53816
0 53818 7 1 2 64214 100433
0 53819 5 1 1 53818
0 53820 7 1 2 53817 53819
0 53821 5 1 1 53820
0 53822 7 1 2 103359 53821
0 53823 5 1 1 53822
0 53824 7 1 2 53814 53823
0 53825 5 1 1 53824
0 53826 7 1 2 83967 53825
0 53827 5 1 1 53826
0 53828 7 1 2 85384 79701
0 53829 7 1 2 103247 53828
0 53830 5 1 1 53829
0 53831 7 1 2 103303 53830
0 53832 5 1 1 53831
0 53833 7 1 2 97743 53832
0 53834 5 1 1 53833
0 53835 7 1 2 90124 98892
0 53836 7 1 2 92375 53835
0 53837 5 1 1 53836
0 53838 7 1 2 53834 53837
0 53839 5 1 1 53838
0 53840 7 1 2 90276 53839
0 53841 5 1 1 53840
0 53842 7 1 2 53827 53841
0 53843 5 1 1 53842
0 53844 7 1 2 65249 53843
0 53845 5 1 1 53844
0 53846 7 2 2 79563 98142
0 53847 7 1 2 66182 81881
0 53848 7 1 2 82705 96065
0 53849 7 1 2 53847 53848
0 53850 7 1 2 103362 53849
0 53851 5 1 1 53850
0 53852 7 1 2 53845 53851
0 53853 7 1 2 53806 53852
0 53854 5 1 1 53853
0 53855 7 1 2 69862 53854
0 53856 5 1 1 53855
0 53857 7 1 2 87935 93922
0 53858 7 2 2 93571 53857
0 53859 5 1 1 103364
0 53860 7 1 2 98939 100910
0 53861 5 1 1 53860
0 53862 7 1 2 88026 98912
0 53863 5 1 1 53862
0 53864 7 1 2 34702 53863
0 53865 5 1 1 53864
0 53866 7 1 2 72674 53865
0 53867 5 1 1 53866
0 53868 7 1 2 53861 53867
0 53869 7 1 2 53859 53868
0 53870 5 1 1 53869
0 53871 7 1 2 83968 53870
0 53872 5 1 1 53871
0 53873 7 1 2 64006 103295
0 53874 5 1 1 53873
0 53875 7 1 2 74479 53874
0 53876 5 1 1 53875
0 53877 7 1 2 92947 95565
0 53878 7 1 2 53876 53877
0 53879 5 1 1 53878
0 53880 7 1 2 53872 53879
0 53881 5 1 1 53880
0 53882 7 1 2 70503 53881
0 53883 5 1 1 53882
0 53884 7 1 2 84177 92948
0 53885 7 1 2 94682 97974
0 53886 7 1 2 53884 53885
0 53887 5 1 1 53886
0 53888 7 1 2 53883 53887
0 53889 5 1 1 53888
0 53890 7 1 2 78566 53889
0 53891 5 1 1 53890
0 53892 7 1 2 53856 53891
0 53893 5 1 1 53892
0 53894 7 1 2 90726 53893
0 53895 5 1 1 53894
0 53896 7 1 2 53755 53895
0 53897 7 1 2 53619 53896
0 53898 5 1 1 53897
0 53899 7 1 2 90216 53898
0 53900 5 1 1 53899
0 53901 7 1 2 79704 97099
0 53902 5 1 1 53901
0 53903 7 1 2 87747 53902
0 53904 5 1 1 53903
0 53905 7 1 2 100985 53904
0 53906 5 1 1 53905
0 53907 7 1 2 65871 102485
0 53908 7 1 2 53906 53907
0 53909 5 1 1 53908
0 53910 7 1 2 87748 97118
0 53911 5 1 1 53910
0 53912 7 2 2 72280 72251
0 53913 7 1 2 87806 95372
0 53914 7 1 2 103366 53913
0 53915 5 1 1 53914
0 53916 7 1 2 53911 53915
0 53917 7 1 2 53909 53916
0 53918 5 1 1 53917
0 53919 7 1 2 65568 53918
0 53920 5 1 1 53919
0 53921 7 1 2 87749 84748
0 53922 5 1 1 53921
0 53923 7 1 2 90444 103312
0 53924 5 1 1 53923
0 53925 7 1 2 53922 53924
0 53926 5 1 1 53925
0 53927 7 1 2 72476 53926
0 53928 5 1 1 53927
0 53929 7 1 2 53920 53928
0 53930 5 1 1 53929
0 53931 7 1 2 87376 53930
0 53932 5 1 1 53931
0 53933 7 1 2 80556 103194
0 53934 5 1 1 53933
0 53935 7 1 2 93220 103221
0 53936 5 1 1 53935
0 53937 7 1 2 53934 53936
0 53938 5 1 1 53937
0 53939 7 1 2 67073 53938
0 53940 5 1 1 53939
0 53941 7 1 2 53932 53940
0 53942 5 1 1 53941
0 53943 7 1 2 100015 53942
0 53944 5 1 1 53943
0 53945 7 3 2 87377 99502
0 53946 7 1 2 84391 98946
0 53947 5 3 1 53946
0 53948 7 1 2 1064 103307
0 53949 5 1 1 53948
0 53950 7 1 2 65569 53949
0 53951 5 1 1 53950
0 53952 7 1 2 103371 53951
0 53953 5 1 1 53952
0 53954 7 1 2 87807 53953
0 53955 5 1 1 53954
0 53956 7 1 2 74928 98329
0 53957 5 1 1 53956
0 53958 7 1 2 103133 53957
0 53959 5 1 1 53958
0 53960 7 1 2 87750 53959
0 53961 5 1 1 53960
0 53962 7 1 2 74736 88020
0 53963 5 1 1 53962
0 53964 7 1 2 67074 103200
0 53965 5 1 1 53964
0 53966 7 1 2 53963 53965
0 53967 5 1 1 53966
0 53968 7 1 2 87004 53967
0 53969 5 1 1 53968
0 53970 7 1 2 53961 53969
0 53971 7 1 2 53955 53970
0 53972 5 1 1 53971
0 53973 7 1 2 103368 53972
0 53974 5 1 1 53973
0 53975 7 1 2 53944 53974
0 53976 5 1 1 53975
0 53977 7 1 2 78622 53976
0 53978 5 1 1 53977
0 53979 7 1 2 102270 102802
0 53980 5 1 1 53979
0 53981 7 1 2 78361 103369
0 53982 5 1 1 53981
0 53983 7 2 2 66321 91649
0 53984 5 1 1 103374
0 53985 7 1 2 62925 102567
0 53986 5 1 1 53985
0 53987 7 1 2 70972 102106
0 53988 5 1 1 53987
0 53989 7 1 2 92142 103188
0 53990 5 1 1 53989
0 53991 7 1 2 64215 53990
0 53992 5 1 1 53991
0 53993 7 1 2 53988 53992
0 53994 7 1 2 53986 53993
0 53995 5 1 1 53994
0 53996 7 1 2 103375 53995
0 53997 5 1 1 53996
0 53998 7 1 2 53982 53997
0 53999 5 1 1 53998
0 54000 7 1 2 87808 53999
0 54001 5 1 1 54000
0 54002 7 1 2 53980 54001
0 54003 5 1 1 54002
0 54004 7 1 2 62677 54003
0 54005 5 1 1 54004
0 54006 7 1 2 91394 87820
0 54007 7 1 2 93280 101987
0 54008 7 1 2 54006 54007
0 54009 5 1 1 54008
0 54010 7 1 2 54005 54009
0 54011 5 1 1 54010
0 54012 7 1 2 64007 54011
0 54013 5 1 1 54012
0 54014 7 2 2 87688 97778
0 54015 7 1 2 79458 96415
0 54016 7 1 2 103376 54015
0 54017 5 1 1 54016
0 54018 7 1 2 87751 79397
0 54019 7 1 2 103370 54018
0 54020 5 1 1 54019
0 54021 7 1 2 54017 54020
0 54022 7 1 2 54013 54021
0 54023 5 1 1 54022
0 54024 7 1 2 70504 54023
0 54025 5 1 1 54024
0 54026 7 1 2 86490 103033
0 54027 5 1 1 54026
0 54028 7 1 2 78349 99503
0 54029 5 1 1 54028
0 54030 7 1 2 54027 54029
0 54031 5 1 1 54030
0 54032 7 1 2 103195 54031
0 54033 5 1 1 54032
0 54034 7 1 2 96207 102212
0 54035 5 1 1 54034
0 54036 7 1 2 54033 54035
0 54037 5 1 1 54036
0 54038 7 1 2 62232 54037
0 54039 5 1 1 54038
0 54040 7 1 2 54025 54039
0 54041 5 1 1 54040
0 54042 7 1 2 78567 54041
0 54043 5 1 1 54042
0 54044 7 1 2 53978 54043
0 54045 5 1 1 54044
0 54046 7 1 2 103217 54045
0 54047 5 1 1 54046
0 54048 7 1 2 87005 103347
0 54049 5 1 1 54048
0 54050 7 1 2 81967 103271
0 54051 5 1 1 54050
0 54052 7 1 2 54049 54051
0 54053 5 1 1 54052
0 54054 7 1 2 67075 54053
0 54055 5 1 1 54054
0 54056 7 1 2 81968 103269
0 54057 5 1 1 54056
0 54058 7 1 2 54055 54057
0 54059 5 1 1 54058
0 54060 7 1 2 73502 54059
0 54061 5 1 1 54060
0 54062 7 1 2 66051 93281
0 54063 5 1 1 54062
0 54064 7 1 2 10383 54063
0 54065 5 1 1 54064
0 54066 7 1 2 67748 54065
0 54067 5 1 1 54066
0 54068 7 1 2 79691 94930
0 54069 5 1 1 54068
0 54070 7 1 2 87006 54069
0 54071 5 1 1 54070
0 54072 7 1 2 54067 54071
0 54073 5 1 1 54072
0 54074 7 1 2 70505 54073
0 54075 5 1 1 54074
0 54076 7 2 2 73782 73169
0 54077 5 1 1 103378
0 54078 7 1 2 94479 54077
0 54079 5 1 1 54078
0 54080 7 1 2 87007 54079
0 54081 5 1 1 54080
0 54082 7 1 2 54075 54081
0 54083 5 1 1 54082
0 54084 7 1 2 78833 54083
0 54085 5 1 1 54084
0 54086 7 1 2 54061 54085
0 54087 5 1 1 54086
0 54088 7 1 2 98893 54087
0 54089 5 1 1 54088
0 54090 7 1 2 103372 103320
0 54091 5 1 1 54090
0 54092 7 1 2 87378 54091
0 54093 5 1 1 54092
0 54094 7 1 2 70506 99445
0 54095 5 1 1 54094
0 54096 7 1 2 54093 54095
0 54097 5 1 1 54096
0 54098 7 1 2 103358 54097
0 54099 5 1 1 54098
0 54100 7 1 2 54089 54099
0 54101 5 1 1 54100
0 54102 7 1 2 69863 54101
0 54103 5 1 1 54102
0 54104 7 1 2 81969 100911
0 54105 5 1 1 54104
0 54106 7 1 2 61681 94962
0 54107 5 1 1 54106
0 54108 7 1 2 54105 54107
0 54109 5 1 1 54108
0 54110 7 1 2 98940 54109
0 54111 5 1 1 54110
0 54112 7 1 2 87379 103365
0 54113 5 1 1 54112
0 54114 7 1 2 54111 54113
0 54115 5 1 1 54114
0 54116 7 1 2 70507 54115
0 54117 5 1 1 54116
0 54118 7 1 2 87380 77970
0 54119 7 1 2 102471 54118
0 54120 5 1 1 54119
0 54121 7 1 2 81403 100031
0 54122 7 1 2 103343 54121
0 54123 5 1 1 54122
0 54124 7 1 2 54120 54123
0 54125 5 1 1 54124
0 54126 7 1 2 70508 54125
0 54127 5 1 1 54126
0 54128 7 1 2 73087 98894
0 54129 5 1 1 54128
0 54130 7 1 2 29800 54129
0 54131 5 1 1 54130
0 54132 7 3 2 87008 75238
0 54133 7 1 2 54131 103380
0 54134 5 1 1 54133
0 54135 7 1 2 54127 54134
0 54136 5 1 1 54135
0 54137 7 1 2 72675 54136
0 54138 5 1 1 54137
0 54139 7 1 2 78350 97744
0 54140 5 1 1 54139
0 54141 7 1 2 95288 95647
0 54142 7 1 2 87821 54141
0 54143 5 1 1 54142
0 54144 7 1 2 54140 54143
0 54145 5 1 1 54144
0 54146 7 1 2 97002 54145
0 54147 5 1 1 54146
0 54148 7 1 2 54138 54147
0 54149 7 1 2 54117 54148
0 54150 5 1 1 54149
0 54151 7 1 2 78568 54150
0 54152 5 1 1 54151
0 54153 7 1 2 54103 54152
0 54154 5 1 1 54153
0 54155 7 1 2 99504 54154
0 54156 5 1 1 54155
0 54157 7 1 2 81974 77677
0 54158 5 1 1 54157
0 54159 7 1 2 86244 54158
0 54160 5 1 1 54159
0 54161 7 1 2 12804 54160
0 54162 5 1 1 54161
0 54163 7 1 2 76727 103289
0 54164 7 1 2 54162 54163
0 54165 5 1 1 54164
0 54166 7 1 2 85365 93282
0 54167 7 1 2 103352 54166
0 54168 5 1 1 54167
0 54169 7 1 2 54165 54168
0 54170 5 1 1 54169
0 54171 7 2 2 69864 54170
0 54172 7 1 2 98895 103383
0 54173 5 1 1 54172
0 54174 7 1 2 78569 103297
0 54175 5 1 1 54174
0 54176 7 1 2 78623 103305
0 54177 5 1 1 54176
0 54178 7 1 2 54175 54177
0 54179 5 1 1 54178
0 54180 7 1 2 87009 54179
0 54181 5 1 1 54180
0 54182 7 1 2 66571 103329
0 54183 5 1 1 54182
0 54184 7 1 2 54181 54183
0 54185 5 1 1 54184
0 54186 7 1 2 97745 54185
0 54187 5 1 1 54186
0 54188 7 1 2 54173 54187
0 54189 5 1 1 54188
0 54190 7 1 2 100016 54189
0 54191 5 1 1 54190
0 54192 7 1 2 54156 54191
0 54193 5 1 1 54192
0 54194 7 1 2 99985 54193
0 54195 5 1 1 54194
0 54196 7 1 2 381 84929
0 54197 5 2 1 54196
0 54198 7 1 2 67538 103385
0 54199 5 1 1 54198
0 54200 7 1 2 100454 103341
0 54201 5 1 1 54200
0 54202 7 1 2 70509 54201
0 54203 5 1 1 54202
0 54204 7 1 2 54199 54203
0 54205 5 1 1 54204
0 54206 7 1 2 65250 54205
0 54207 5 1 1 54206
0 54208 7 1 2 76353 85432
0 54209 5 1 1 54208
0 54210 7 1 2 54207 54209
0 54211 5 1 1 54210
0 54212 7 1 2 77400 54211
0 54213 5 1 1 54212
0 54214 7 1 2 77099 102947
0 54215 5 1 1 54214
0 54216 7 1 2 54213 54215
0 54217 5 1 1 54216
0 54218 7 1 2 87010 54217
0 54219 5 1 1 54218
0 54220 7 1 2 73503 103273
0 54221 5 1 1 54220
0 54222 7 1 2 74095 80663
0 54223 5 1 1 54222
0 54224 7 1 2 54221 54223
0 54225 5 1 1 54224
0 54226 7 1 2 69865 54225
0 54227 5 1 1 54226
0 54228 7 1 2 94501 100907
0 54229 5 1 1 54228
0 54230 7 1 2 102772 54229
0 54231 5 1 1 54230
0 54232 7 1 2 54227 54231
0 54233 5 1 1 54232
0 54234 7 1 2 81970 54233
0 54235 5 1 1 54234
0 54236 7 1 2 54219 54235
0 54237 5 1 1 54236
0 54238 7 1 2 99505 54237
0 54239 5 1 1 54238
0 54240 7 1 2 100017 103384
0 54241 5 1 1 54240
0 54242 7 1 2 54239 54241
0 54243 5 1 1 54242
0 54244 7 1 2 87752 54243
0 54245 5 1 1 54244
0 54246 7 1 2 85848 100018
0 54247 5 1 1 54246
0 54248 7 1 2 61415 89566
0 54249 5 1 1 54248
0 54250 7 1 2 54247 54249
0 54251 5 1 1 54250
0 54252 7 1 2 103354 103290
0 54253 7 1 2 54251 54252
0 54254 5 1 1 54253
0 54255 7 1 2 54245 54254
0 54256 5 1 1 54255
0 54257 7 1 2 103186 54256
0 54258 5 1 1 54257
0 54259 7 1 2 87809 103278
0 54260 5 1 1 54259
0 54261 7 3 2 61326 97381
0 54262 7 1 2 88452 103387
0 54263 5 1 1 54262
0 54264 7 1 2 54260 54263
0 54265 5 1 1 54264
0 54266 7 1 2 62678 54265
0 54267 5 1 1 54266
0 54268 7 1 2 103275 48010
0 54269 5 1 1 54268
0 54270 7 1 2 87753 54269
0 54271 5 1 1 54270
0 54272 7 1 2 54267 54271
0 54273 5 1 1 54272
0 54274 7 1 2 99506 54273
0 54275 5 1 1 54274
0 54276 7 1 2 103034 103388
0 54277 7 1 2 102536 54276
0 54278 5 1 1 54277
0 54279 7 1 2 54275 54278
0 54280 5 1 1 54279
0 54281 7 1 2 87381 54280
0 54282 5 1 1 54281
0 54283 7 1 2 78570 100801
0 54284 7 1 2 103381 54283
0 54285 5 1 1 54284
0 54286 7 1 2 54282 54285
0 54287 5 1 1 54286
0 54288 7 1 2 103218 54287
0 54289 5 1 1 54288
0 54290 7 1 2 81971 89782
0 54291 5 1 1 54290
0 54292 7 1 2 102920 54291
0 54293 5 1 1 54292
0 54294 7 1 2 91815 102356
0 54295 7 1 2 100842 54294
0 54296 7 1 2 102148 54295
0 54297 7 1 2 54293 54296
0 54298 5 1 1 54297
0 54299 7 1 2 54289 54298
0 54300 5 1 1 54299
0 54301 7 1 2 72676 54300
0 54302 5 1 1 54301
0 54303 7 1 2 81972 78219
0 54304 7 1 2 100187 54303
0 54305 5 1 1 54304
0 54306 7 1 2 90247 99824
0 54307 7 1 2 103337 54306
0 54308 5 1 1 54307
0 54309 7 1 2 54305 54308
0 54310 5 1 1 54309
0 54311 7 1 2 66784 99619
0 54312 7 1 2 95432 54311
0 54313 7 1 2 98726 54312
0 54314 7 1 2 54310 54313
0 54315 5 1 1 54314
0 54316 7 1 2 99926 103210
0 54317 5 1 1 54316
0 54318 7 1 2 61416 84060
0 54319 7 1 2 102117 54318
0 54320 5 1 1 54319
0 54321 7 1 2 54317 54320
0 54322 5 1 1 54321
0 54323 7 1 2 87754 54322
0 54324 5 1 1 54323
0 54325 7 1 2 91002 87827
0 54326 7 1 2 90851 54325
0 54327 7 1 2 85199 54326
0 54328 5 1 1 54327
0 54329 7 1 2 54324 54328
0 54330 5 1 1 54329
0 54331 7 1 2 87382 103219
0 54332 7 1 2 54330 54331
0 54333 5 1 1 54332
0 54334 7 1 2 54315 54333
0 54335 5 1 1 54334
0 54336 7 1 2 71379 54335
0 54337 5 1 1 54336
0 54338 7 1 2 54302 54337
0 54339 7 1 2 54258 54338
0 54340 7 1 2 54195 54339
0 54341 7 1 2 54047 54340
0 54342 7 1 2 53900 54341
0 54343 7 1 2 53359 54342
0 54344 7 1 2 52779 54343
0 54345 7 1 2 52365 54344
0 54346 5 1 1 54345
0 54347 7 1 2 101814 54346
0 54348 5 1 1 54347
0 54349 7 1 2 94191 101064
0 54350 5 1 1 54349
0 54351 7 1 2 65872 95300
0 54352 5 1 1 54351
0 54353 7 1 2 84906 54352
0 54354 5 1 1 54353
0 54355 7 1 2 101950 54354
0 54356 5 1 1 54355
0 54357 7 1 2 68879 102799
0 54358 5 1 1 54357
0 54359 7 1 2 71656 101278
0 54360 5 1 1 54359
0 54361 7 1 2 54358 54360
0 54362 5 1 1 54361
0 54363 7 1 2 62679 54362
0 54364 5 1 1 54363
0 54365 7 1 2 64008 102800
0 54366 5 1 1 54365
0 54367 7 1 2 84324 96869
0 54368 5 1 1 54367
0 54369 7 1 2 78366 54368
0 54370 7 1 2 54366 54369
0 54371 5 1 1 54370
0 54372 7 1 2 67539 54371
0 54373 5 1 1 54372
0 54374 7 1 2 54364 54373
0 54375 5 2 1 54374
0 54376 7 1 2 100206 103390
0 54377 5 1 1 54376
0 54378 7 1 2 54356 54377
0 54379 5 1 1 54378
0 54380 7 1 2 78989 54379
0 54381 5 1 1 54380
0 54382 7 1 2 1222 102972
0 54383 5 1 1 54382
0 54384 7 1 2 69066 54383
0 54385 5 2 1 54384
0 54386 7 1 2 89848 40426
0 54387 5 2 1 54386
0 54388 7 1 2 64216 103394
0 54389 5 2 1 54388
0 54390 7 2 2 103392 103396
0 54391 5 1 1 103398
0 54392 7 1 2 65873 54391
0 54393 5 1 1 54392
0 54394 7 2 2 85498 82898
0 54395 7 1 2 72427 103400
0 54396 5 1 1 54395
0 54397 7 1 2 54393 54396
0 54398 5 1 1 54397
0 54399 7 1 2 89404 100563
0 54400 7 1 2 54398 54399
0 54401 5 1 1 54400
0 54402 7 1 2 54381 54401
0 54403 5 1 1 54402
0 54404 7 1 2 69261 54403
0 54405 5 1 1 54404
0 54406 7 1 2 102250 102906
0 54407 5 1 1 54406
0 54408 7 1 2 85925 98385
0 54409 5 1 1 54408
0 54410 7 1 2 54407 54409
0 54411 5 1 1 54410
0 54412 7 1 2 61417 54411
0 54413 5 1 1 54412
0 54414 7 1 2 85926 98409
0 54415 5 1 1 54414
0 54416 7 1 2 54413 54415
0 54417 5 1 1 54416
0 54418 7 1 2 76735 54417
0 54419 5 1 1 54418
0 54420 7 1 2 92587 97503
0 54421 7 1 2 100776 54420
0 54422 5 1 1 54421
0 54423 7 1 2 54419 54422
0 54424 5 1 1 54423
0 54425 7 1 2 93138 54424
0 54426 5 1 1 54425
0 54427 7 1 2 54405 54426
0 54428 5 1 1 54427
0 54429 7 1 2 67829 54428
0 54430 5 1 1 54429
0 54431 7 1 2 94534 101951
0 54432 5 1 1 54431
0 54433 7 2 2 84233 90685
0 54434 7 1 2 95218 103402
0 54435 5 1 1 54434
0 54436 7 1 2 54432 54435
0 54437 5 1 1 54436
0 54438 7 2 2 102152 54437
0 54439 7 1 2 97340 103404
0 54440 5 1 1 54439
0 54441 7 1 2 54430 54440
0 54442 5 1 1 54441
0 54443 7 1 2 66183 54442
0 54444 5 1 1 54443
0 54445 7 1 2 103405 98506
0 54446 5 1 1 54445
0 54447 7 2 2 90727 93139
0 54448 7 1 2 102993 103406
0 54449 5 1 1 54448
0 54450 7 1 2 67830 102997
0 54451 7 1 2 91251 54450
0 54452 5 1 1 54451
0 54453 7 1 2 54449 54452
0 54454 5 1 1 54453
0 54455 7 1 2 78990 54454
0 54456 5 1 1 54455
0 54457 7 2 2 87846 93060
0 54458 5 1 1 103408
0 54459 7 1 2 75534 103409
0 54460 5 1 1 54459
0 54461 7 1 2 92257 100119
0 54462 5 1 1 54461
0 54463 7 1 2 54460 54462
0 54464 5 1 1 54463
0 54465 7 1 2 66322 54464
0 54466 5 1 1 54465
0 54467 7 1 2 77824 101888
0 54468 5 1 1 54467
0 54469 7 1 2 54466 54468
0 54470 5 1 1 54469
0 54471 7 1 2 100481 97504
0 54472 7 1 2 54470 54471
0 54473 5 1 1 54472
0 54474 7 1 2 54456 54473
0 54475 5 1 1 54474
0 54476 7 1 2 66184 54475
0 54477 5 1 1 54476
0 54478 7 1 2 97084 97408
0 54479 7 1 2 102994 54478
0 54480 5 1 1 54479
0 54481 7 1 2 54477 54480
0 54482 5 1 1 54481
0 54483 7 1 2 73504 54482
0 54484 5 1 1 54483
0 54485 7 1 2 54446 54484
0 54486 7 1 2 54444 54485
0 54487 5 1 1 54486
0 54488 7 1 2 70510 54487
0 54489 5 1 1 54488
0 54490 7 2 2 92816 98713
0 54491 5 1 1 103410
0 54492 7 4 2 96114 99702
0 54493 5 2 1 103412
0 54494 7 1 2 54491 103416
0 54495 5 1 1 54494
0 54496 7 1 2 61418 54495
0 54497 5 1 1 54496
0 54498 7 1 2 64009 100804
0 54499 7 1 2 99614 54498
0 54500 5 1 1 54499
0 54501 7 1 2 54497 54500
0 54502 5 1 1 54501
0 54503 7 1 2 78991 54502
0 54504 5 1 1 54503
0 54505 7 1 2 66323 103059
0 54506 5 1 1 54505
0 54507 7 1 2 101889 54506
0 54508 5 2 1 54507
0 54509 7 1 2 82007 87115
0 54510 7 1 2 103418 54509
0 54511 5 1 1 54510
0 54512 7 1 2 54504 54511
0 54513 5 1 1 54512
0 54514 7 1 2 72089 54513
0 54515 5 1 1 54514
0 54516 7 1 2 99586 97505
0 54517 5 1 1 54516
0 54518 7 2 2 78851 99833
0 54519 5 1 1 103420
0 54520 7 1 2 54517 54519
0 54521 5 1 1 54520
0 54522 7 1 2 64595 86727
0 54523 7 1 2 54521 54522
0 54524 5 1 1 54523
0 54525 7 1 2 89641 73969
0 54526 5 1 1 54525
0 54527 7 1 2 84325 89295
0 54528 5 1 1 54527
0 54529 7 1 2 54526 54528
0 54530 5 1 1 54529
0 54531 7 1 2 67904 83903
0 54532 7 1 2 54530 54531
0 54533 5 1 1 54532
0 54534 7 1 2 54524 54533
0 54535 5 1 1 54534
0 54536 7 1 2 69262 54535
0 54537 5 1 1 54536
0 54538 7 1 2 86728 98405
0 54539 7 1 2 96550 54538
0 54540 5 1 1 54539
0 54541 7 1 2 66324 54540
0 54542 7 1 2 54537 54541
0 54543 5 1 1 54542
0 54544 7 1 2 67905 86729
0 54545 7 1 2 96505 54544
0 54546 5 1 1 54545
0 54547 7 1 2 82023 103413
0 54548 5 1 1 54547
0 54549 7 1 2 61419 54548
0 54550 7 1 2 54546 54549
0 54551 5 1 1 54550
0 54552 7 1 2 70781 54551
0 54553 7 1 2 54543 54552
0 54554 5 1 1 54553
0 54555 7 1 2 54515 54554
0 54556 5 1 1 54555
0 54557 7 1 2 62680 54556
0 54558 5 1 1 54557
0 54559 7 1 2 54458 103417
0 54560 5 1 1 54559
0 54561 7 1 2 61420 54560
0 54562 5 1 1 54561
0 54563 7 1 2 66325 87847
0 54564 7 1 2 100526 54563
0 54565 5 1 1 54564
0 54566 7 1 2 54562 54565
0 54567 5 1 1 54566
0 54568 7 1 2 78992 54567
0 54569 5 1 1 54568
0 54570 7 1 2 95012 103419
0 54571 5 1 1 54570
0 54572 7 1 2 54569 54571
0 54573 5 1 1 54572
0 54574 7 1 2 72090 54573
0 54575 5 1 1 54574
0 54576 7 1 2 91816 92035
0 54577 7 1 2 103414 54576
0 54578 5 1 1 54577
0 54579 7 1 2 54575 54578
0 54580 5 1 1 54579
0 54581 7 1 2 64010 54580
0 54582 5 1 1 54581
0 54583 7 1 2 54558 54582
0 54584 5 1 1 54583
0 54585 7 1 2 67831 54584
0 54586 5 1 1 54585
0 54587 7 1 2 88442 101773
0 54588 5 1 1 54587
0 54589 7 1 2 76283 102726
0 54590 5 1 1 54589
0 54591 7 1 2 54588 54590
0 54592 5 1 1 54591
0 54593 7 1 2 66326 54592
0 54594 5 1 1 54593
0 54595 7 1 2 75645 100555
0 54596 5 1 1 54595
0 54597 7 1 2 54594 54596
0 54598 5 1 1 54597
0 54599 7 2 2 102153 54598
0 54600 7 1 2 97341 103422
0 54601 5 1 1 54600
0 54602 7 1 2 54586 54601
0 54603 5 1 1 54602
0 54604 7 1 2 66185 54603
0 54605 5 1 1 54604
0 54606 7 1 2 98507 103423
0 54607 5 1 1 54606
0 54608 7 1 2 54605 54607
0 54609 5 1 1 54608
0 54610 7 1 2 65570 54609
0 54611 5 1 1 54610
0 54612 7 2 2 82008 82814
0 54613 7 1 2 97147 103424
0 54614 5 1 1 54613
0 54615 7 1 2 96349 97247
0 54616 5 1 1 54615
0 54617 7 1 2 54614 54616
0 54618 5 1 1 54617
0 54619 7 1 2 65571 54618
0 54620 5 1 1 54619
0 54621 7 1 2 92239 96501
0 54622 5 1 1 54621
0 54623 7 1 2 54620 54622
0 54624 5 1 1 54623
0 54625 7 1 2 67832 54624
0 54626 5 1 1 54625
0 54627 7 1 2 96920 99745
0 54628 7 1 2 98134 54627
0 54629 5 1 1 54628
0 54630 7 1 2 54626 54629
0 54631 5 1 1 54630
0 54632 7 1 2 99101 54631
0 54633 5 1 1 54632
0 54634 7 2 2 71380 83924
0 54635 7 1 2 65572 93631
0 54636 7 2 2 103426 54635
0 54637 7 1 2 90646 103428
0 54638 5 1 1 54637
0 54639 7 1 2 93610 103427
0 54640 5 1 1 54639
0 54641 7 1 2 89288 99306
0 54642 7 1 2 96077 54641
0 54643 5 1 1 54642
0 54644 7 1 2 54640 54643
0 54645 5 1 1 54644
0 54646 7 1 2 73088 54645
0 54647 5 1 1 54646
0 54648 7 1 2 69637 92830
0 54649 7 1 2 98444 103006
0 54650 7 1 2 54648 54649
0 54651 5 1 1 54650
0 54652 7 1 2 54647 54651
0 54653 5 1 1 54652
0 54654 7 1 2 90686 54653
0 54655 5 1 1 54654
0 54656 7 1 2 54638 54655
0 54657 7 1 2 54633 54656
0 54658 5 1 1 54657
0 54659 7 1 2 66186 54658
0 54660 5 1 1 54659
0 54661 7 1 2 92461 103429
0 54662 5 1 1 54661
0 54663 7 1 2 73089 102123
0 54664 7 1 2 98508 54663
0 54665 7 1 2 99102 54664
0 54666 5 1 1 54665
0 54667 7 1 2 54662 54666
0 54668 7 1 2 54660 54667
0 54669 5 1 1 54668
0 54670 7 1 2 72677 54669
0 54671 5 1 1 54670
0 54672 7 1 2 54611 54671
0 54673 7 1 2 54489 54672
0 54674 5 1 1 54673
0 54675 7 1 2 80590 54674
0 54676 5 1 1 54675
0 54677 7 1 2 66327 102197
0 54678 5 1 1 54677
0 54679 7 1 2 101890 54678
0 54680 5 1 1 54679
0 54681 7 1 2 72207 54680
0 54682 5 1 1 54681
0 54683 7 1 2 67906 103281
0 54684 5 1 1 54683
0 54685 7 1 2 54682 54684
0 54686 5 1 1 54685
0 54687 7 1 2 71265 54686
0 54688 5 1 1 54687
0 54689 7 1 2 64408 72588
0 54690 7 1 2 101376 54689
0 54691 5 1 1 54690
0 54692 7 1 2 54688 54691
0 54693 5 1 1 54692
0 54694 7 1 2 96867 54693
0 54695 5 1 1 54694
0 54696 7 1 2 76581 93632
0 54697 7 1 2 102918 54696
0 54698 5 1 1 54697
0 54699 7 1 2 54695 54698
0 54700 5 1 1 54699
0 54701 7 1 2 86066 54700
0 54702 5 1 1 54701
0 54703 7 1 2 90628 87943
0 54704 5 1 1 54703
0 54705 7 1 2 83762 103229
0 54706 7 1 2 92977 54705
0 54707 5 1 1 54706
0 54708 7 1 2 54704 54707
0 54709 5 1 1 54708
0 54710 7 1 2 64596 54709
0 54711 5 1 1 54710
0 54712 7 3 2 93140 93835
0 54713 7 1 2 64217 75668
0 54714 7 1 2 103430 54713
0 54715 5 1 1 54714
0 54716 7 1 2 85477 102890
0 54717 7 1 2 100814 54716
0 54718 5 1 1 54717
0 54719 7 1 2 54715 54718
0 54720 5 1 1 54719
0 54721 7 1 2 70973 54720
0 54722 5 1 1 54721
0 54723 7 1 2 90637 41096
0 54724 5 1 1 54723
0 54725 7 1 2 88033 101374
0 54726 7 1 2 54724 54725
0 54727 5 1 1 54726
0 54728 7 1 2 54722 54727
0 54729 5 1 1 54728
0 54730 7 1 2 67749 54729
0 54731 5 1 1 54730
0 54732 7 1 2 54711 54731
0 54733 5 1 1 54732
0 54734 7 1 2 77040 54733
0 54735 5 1 1 54734
0 54736 7 1 2 85344 103171
0 54737 5 2 1 54736
0 54738 7 1 2 102763 103433
0 54739 5 1 1 54738
0 54740 7 1 2 87986 94331
0 54741 5 1 1 54740
0 54742 7 1 2 96660 54741
0 54743 5 1 1 54742
0 54744 7 1 2 100301 54743
0 54745 5 1 1 54744
0 54746 7 1 2 54739 54745
0 54747 5 1 1 54746
0 54748 7 1 2 64409 77669
0 54749 7 1 2 54747 54748
0 54750 5 1 1 54749
0 54751 7 1 2 100795 99635
0 54752 7 2 2 96766 54751
0 54753 7 1 2 64218 103435
0 54754 5 1 1 54753
0 54755 7 1 2 72208 85478
0 54756 5 1 1 54755
0 54757 7 1 2 69067 77755
0 54758 5 1 1 54757
0 54759 7 1 2 54756 54758
0 54760 5 1 1 54759
0 54761 7 1 2 103431 54760
0 54762 5 1 1 54761
0 54763 7 1 2 54754 54762
0 54764 5 1 1 54763
0 54765 7 1 2 94806 54764
0 54766 5 1 1 54765
0 54767 7 3 2 62233 79300
0 54768 5 1 1 103437
0 54769 7 1 2 103415 103438
0 54770 5 1 1 54769
0 54771 7 2 2 92817 99636
0 54772 5 1 1 103440
0 54773 7 1 2 75903 77670
0 54774 7 1 2 103441 54773
0 54775 5 1 1 54774
0 54776 7 1 2 54770 54775
0 54777 5 1 1 54776
0 54778 7 1 2 66328 54777
0 54779 5 1 1 54778
0 54780 7 1 2 100520 103439
0 54781 5 1 1 54780
0 54782 7 1 2 95923 100336
0 54783 5 1 1 54782
0 54784 7 1 2 54781 54783
0 54785 5 1 1 54784
0 54786 7 1 2 100368 54785
0 54787 5 1 1 54786
0 54788 7 1 2 54779 54787
0 54789 5 1 1 54788
0 54790 7 1 2 98330 54789
0 54791 5 1 1 54790
0 54792 7 1 2 54766 54791
0 54793 7 1 2 54750 54792
0 54794 7 1 2 54735 54793
0 54795 5 1 1 54794
0 54796 7 1 2 70511 54795
0 54797 5 1 1 54796
0 54798 7 1 2 54702 54797
0 54799 5 1 1 54798
0 54800 7 1 2 82790 54799
0 54801 5 1 1 54800
0 54802 7 1 2 84733 102998
0 54803 5 1 1 54802
0 54804 7 1 2 85899 100120
0 54805 5 1 1 54804
0 54806 7 1 2 54772 54805
0 54807 5 1 1 54806
0 54808 7 1 2 61421 54807
0 54809 5 1 1 54808
0 54810 7 1 2 42557 99612
0 54811 5 1 1 54810
0 54812 7 1 2 66329 93023
0 54813 7 1 2 54811 54812
0 54814 5 1 1 54813
0 54815 7 1 2 54809 54814
0 54816 5 1 1 54815
0 54817 7 1 2 67540 54816
0 54818 5 1 1 54817
0 54819 7 1 2 89859 101463
0 54820 5 1 1 54819
0 54821 7 1 2 54818 54820
0 54822 5 1 1 54821
0 54823 7 1 2 69068 54822
0 54824 5 1 1 54823
0 54825 7 1 2 54803 54824
0 54826 5 1 1 54825
0 54827 7 1 2 67750 54826
0 54828 5 1 1 54827
0 54829 7 1 2 79659 92818
0 54830 7 1 2 102746 54829
0 54831 5 1 1 54830
0 54832 7 1 2 54828 54831
0 54833 5 2 1 54832
0 54834 7 1 2 79945 87135
0 54835 7 1 2 103442 54834
0 54836 5 1 1 54835
0 54837 7 1 2 54801 54836
0 54838 5 1 1 54837
0 54839 7 1 2 61916 54838
0 54840 5 1 1 54839
0 54841 7 1 2 78985 76728
0 54842 7 1 2 102260 54841
0 54843 7 1 2 103443 54842
0 54844 5 1 1 54843
0 54845 7 1 2 54840 54844
0 54846 5 1 1 54845
0 54847 7 1 2 67833 54846
0 54848 5 1 1 54847
0 54849 7 2 2 67907 64410
0 54850 7 2 2 86145 92686
0 54851 5 1 1 103446
0 54852 7 1 2 101195 103447
0 54853 5 1 1 54852
0 54854 7 1 2 75688 79459
0 54855 7 1 2 102261 54854
0 54856 5 1 1 54855
0 54857 7 1 2 62926 86103
0 54858 5 1 1 54857
0 54859 7 1 2 61917 102964
0 54860 7 1 2 54858 54859
0 54861 5 1 1 54860
0 54862 7 1 2 54856 54861
0 54863 5 1 1 54862
0 54864 7 1 2 84247 54863
0 54865 5 1 1 54864
0 54866 7 1 2 54853 54865
0 54867 5 1 1 54866
0 54868 7 1 2 69069 54867
0 54869 5 1 1 54868
0 54870 7 1 2 67076 102986
0 54871 5 1 1 54870
0 54872 7 1 2 80591 97945
0 54873 7 1 2 54871 54872
0 54874 5 1 1 54873
0 54875 7 1 2 54869 54874
0 54876 5 1 1 54875
0 54877 7 1 2 73505 54876
0 54878 5 1 1 54877
0 54879 7 1 2 43318 52576
0 54880 5 1 1 54879
0 54881 7 1 2 77041 54880
0 54882 5 1 1 54881
0 54883 7 1 2 76736 77671
0 54884 7 1 2 101818 54883
0 54885 5 1 1 54884
0 54886 7 1 2 54882 54885
0 54887 5 1 1 54886
0 54888 7 1 2 83911 54887
0 54889 5 1 1 54888
0 54890 7 1 2 54878 54889
0 54891 5 1 1 54890
0 54892 7 2 2 103444 54891
0 54893 7 1 2 90949 103448
0 54894 5 1 1 54893
0 54895 7 1 2 54848 54894
0 54896 5 1 1 54895
0 54897 7 1 2 66187 54896
0 54898 5 1 1 54897
0 54899 7 1 2 103449 100316
0 54900 5 1 1 54899
0 54901 7 1 2 69148 54900
0 54902 7 1 2 54898 54901
0 54903 7 1 2 54676 54902
0 54904 5 1 1 54903
0 54905 7 2 2 77912 86500
0 54906 5 1 1 103450
0 54907 7 1 2 86475 54906
0 54908 5 1 1 54907
0 54909 7 1 2 72209 54908
0 54910 5 1 1 54909
0 54911 7 1 2 96670 100422
0 54912 5 1 1 54911
0 54913 7 1 2 65874 54912
0 54914 5 1 1 54913
0 54915 7 1 2 87050 54914
0 54916 5 1 1 54915
0 54917 7 1 2 65573 54916
0 54918 5 1 1 54917
0 54919 7 1 2 54910 54918
0 54920 5 1 1 54919
0 54921 7 1 2 83904 54920
0 54922 5 1 1 54921
0 54923 7 1 2 65574 103174
0 54924 5 1 1 54923
0 54925 7 1 2 72233 54924
0 54926 5 1 1 54925
0 54927 7 1 2 83912 54926
0 54928 5 1 1 54927
0 54929 7 1 2 54922 54928
0 54930 5 1 1 54929
0 54931 7 1 2 70157 54930
0 54932 5 1 1 54931
0 54933 7 1 2 77050 103125
0 54934 5 1 1 54933
0 54935 7 1 2 83925 4645
0 54936 7 1 2 54934 54935
0 54937 5 1 1 54936
0 54938 7 1 2 54932 54937
0 54939 5 1 1 54938
0 54940 7 1 2 63043 54939
0 54941 5 1 1 54940
0 54942 7 1 2 63044 83926
0 54943 7 1 2 103022 54942
0 54944 5 1 1 54943
0 54945 7 1 2 82009 99762
0 54946 7 1 2 103103 54945
0 54947 5 1 1 54946
0 54948 7 1 2 54944 54947
0 54949 5 1 1 54948
0 54950 7 1 2 65251 54949
0 54951 5 1 1 54950
0 54952 7 1 2 100521 103017
0 54953 5 1 1 54952
0 54954 7 1 2 64597 100337
0 54955 5 1 1 54954
0 54956 7 1 2 54953 54955
0 54957 5 1 1 54956
0 54958 7 1 2 61918 86098
0 54959 7 1 2 54957 54958
0 54960 5 1 1 54959
0 54961 7 1 2 54951 54960
0 54962 5 1 1 54961
0 54963 7 1 2 72678 54962
0 54964 5 1 1 54963
0 54965 7 1 2 88318 78202
0 54966 5 1 1 54965
0 54967 7 1 2 81135 54966
0 54968 5 1 1 54967
0 54969 7 1 2 71381 54968
0 54970 5 1 1 54969
0 54971 7 1 2 73506 91252
0 54972 5 1 1 54971
0 54973 7 1 2 84907 54972
0 54974 5 1 1 54973
0 54975 7 1 2 65575 54974
0 54976 5 1 1 54975
0 54977 7 1 2 54976 103373
0 54978 5 1 1 54977
0 54979 7 1 2 70158 54978
0 54980 5 1 1 54979
0 54981 7 2 2 54970 54980
0 54982 5 1 1 103452
0 54983 7 1 2 99672 97506
0 54984 7 1 2 54982 54983
0 54985 5 1 1 54984
0 54986 7 1 2 54964 54985
0 54987 7 1 2 54941 54986
0 54988 5 1 1 54987
0 54989 7 1 2 61422 54988
0 54990 5 1 1 54989
0 54991 7 1 2 82010 98771
0 54992 7 1 2 46981 54991
0 54993 5 1 1 54992
0 54994 7 1 2 71382 79556
0 54995 5 1 1 54994
0 54996 7 1 2 77678 54995
0 54997 5 1 1 54996
0 54998 7 1 2 61423 103421
0 54999 7 1 2 54997 54998
0 55000 5 1 1 54999
0 55001 7 1 2 54993 55000
0 55002 5 1 1 55001
0 55003 7 1 2 69448 55002
0 55004 5 1 1 55003
0 55005 7 2 2 71383 86336
0 55006 7 1 2 86936 99507
0 55007 7 1 2 98406 55006
0 55008 7 1 2 103454 55007
0 55009 5 1 1 55008
0 55010 7 1 2 55004 55009
0 55011 5 1 1 55010
0 55012 7 1 2 78351 55011
0 55013 5 1 1 55012
0 55014 7 1 2 70159 103018
0 55015 5 1 1 55014
0 55016 7 1 2 55015 101419
0 55017 5 1 1 55016
0 55018 7 1 2 84371 55017
0 55019 5 1 1 55018
0 55020 7 1 2 103453 55019
0 55021 5 1 1 55020
0 55022 7 1 2 92732 98410
0 55023 7 1 2 55021 55022
0 55024 5 1 1 55023
0 55025 7 1 2 55013 55024
0 55026 7 1 2 54990 55025
0 55027 5 1 1 55026
0 55028 7 1 2 99768 55027
0 55029 5 1 1 55028
0 55030 7 2 2 76951 103322
0 55031 5 1 1 103456
0 55032 7 1 2 84666 91153
0 55033 5 1 1 55032
0 55034 7 1 2 55031 55033
0 55035 5 1 1 55034
0 55036 7 1 2 64011 55035
0 55037 5 1 1 55036
0 55038 7 1 2 79043 100993
0 55039 5 1 1 55038
0 55040 7 1 2 55037 55039
0 55041 5 1 1 55040
0 55042 7 1 2 62681 55041
0 55043 5 1 1 55042
0 55044 7 3 2 62234 77338
0 55045 5 1 1 103458
0 55046 7 1 2 72713 100957
0 55047 5 1 1 55046
0 55048 7 1 2 55045 55047
0 55049 5 1 1 55048
0 55050 7 1 2 86802 55049
0 55051 5 1 1 55050
0 55052 7 1 2 72210 94807
0 55053 5 1 1 55052
0 55054 7 1 2 2133 54768
0 55055 7 1 2 55053 55054
0 55056 5 1 1 55055
0 55057 7 1 2 70512 55056
0 55058 5 1 1 55057
0 55059 7 1 2 55051 55058
0 55060 7 1 2 55043 55059
0 55061 5 1 1 55060
0 55062 7 1 2 93885 103425
0 55063 7 1 2 55061 55062
0 55064 5 1 1 55063
0 55065 7 3 2 82932 102333
0 55066 7 1 2 85576 103461
0 55067 5 1 1 55066
0 55068 7 1 2 75425 82815
0 55069 7 1 2 99868 55068
0 55070 5 1 1 55069
0 55071 7 1 2 55067 55070
0 55072 5 1 1 55071
0 55073 7 1 2 65576 55072
0 55074 5 1 1 55073
0 55075 7 1 2 67077 103462
0 55076 5 1 1 55075
0 55077 7 1 2 55074 55076
0 55078 5 1 1 55077
0 55079 7 1 2 70160 55078
0 55080 5 1 1 55079
0 55081 7 1 2 84427 102951
0 55082 7 1 2 103014 55081
0 55083 5 1 1 55082
0 55084 7 1 2 55080 55083
0 55085 5 1 1 55084
0 55086 7 1 2 94135 55085
0 55087 5 1 1 55086
0 55088 7 1 2 76910 94559
0 55089 5 1 1 55088
0 55090 7 1 2 102404 55089
0 55091 5 1 1 55090
0 55092 7 1 2 70782 55091
0 55093 5 1 1 55092
0 55094 7 1 2 72901 93299
0 55095 5 2 1 55094
0 55096 7 1 2 89525 78203
0 55097 7 1 2 103464 55096
0 55098 5 1 1 55097
0 55099 7 1 2 55093 55098
0 55100 5 1 1 55099
0 55101 7 1 2 103463 55100
0 55102 5 1 1 55101
0 55103 7 1 2 55087 55102
0 55104 7 1 2 55064 55103
0 55105 5 1 1 55104
0 55106 7 1 2 93836 55105
0 55107 5 1 1 55106
0 55108 7 1 2 89157 86285
0 55109 5 1 1 55108
0 55110 7 1 2 83918 55109
0 55111 5 1 1 55110
0 55112 7 1 2 62682 55111
0 55113 5 1 1 55112
0 55114 7 1 2 89401 83919
0 55115 5 1 1 55114
0 55116 7 1 2 73558 55115
0 55117 5 1 1 55116
0 55118 7 1 2 55113 55117
0 55119 5 1 1 55118
0 55120 7 1 2 73229 55119
0 55121 5 1 1 55120
0 55122 7 1 2 86880 96015
0 55123 5 1 1 55122
0 55124 7 1 2 83905 101510
0 55125 5 1 1 55124
0 55126 7 1 2 55123 55125
0 55127 5 1 1 55126
0 55128 7 1 2 92350 55127
0 55129 5 1 1 55128
0 55130 7 1 2 55121 55129
0 55131 5 1 1 55130
0 55132 7 1 2 64219 55131
0 55133 5 1 1 55132
0 55134 7 1 2 74160 83989
0 55135 5 1 1 55134
0 55136 7 1 2 55133 55135
0 55137 5 1 1 55136
0 55138 7 1 2 76952 55137
0 55139 5 1 1 55138
0 55140 7 1 2 72752 86481
0 55141 5 1 1 55140
0 55142 7 1 2 79039 55141
0 55143 5 1 1 55142
0 55144 7 1 2 83913 55143
0 55145 5 1 1 55144
0 55146 7 1 2 79810 86286
0 55147 7 1 2 79055 55146
0 55148 5 1 1 55147
0 55149 7 1 2 55145 55148
0 55150 5 1 1 55149
0 55151 7 1 2 62683 55150
0 55152 5 1 1 55151
0 55153 7 3 2 67541 101511
0 55154 5 3 1 103466
0 55155 7 1 2 76255 103467
0 55156 7 1 2 89424 55155
0 55157 5 1 1 55156
0 55158 7 1 2 55152 55157
0 55159 5 1 1 55158
0 55160 7 1 2 75556 55159
0 55161 5 1 1 55160
0 55162 7 1 2 87997 100539
0 55163 5 1 1 55162
0 55164 7 1 2 101641 101794
0 55165 5 1 1 55164
0 55166 7 1 2 101512 55165
0 55167 5 1 1 55166
0 55168 7 1 2 73273 55167
0 55169 7 1 2 55163 55168
0 55170 5 1 1 55169
0 55171 7 1 2 65577 55170
0 55172 5 1 1 55171
0 55173 7 1 2 72739 55172
0 55174 5 1 1 55173
0 55175 7 1 2 89425 55174
0 55176 5 1 1 55175
0 55177 7 1 2 86287 102264
0 55178 5 1 1 55177
0 55179 7 1 2 54851 55178
0 55180 5 1 1 55179
0 55181 7 1 2 102966 55180
0 55182 5 1 1 55181
0 55183 7 1 2 55176 55182
0 55184 7 1 2 55161 55183
0 55185 7 1 2 55139 55184
0 55186 5 1 1 55185
0 55187 7 1 2 91034 55186
0 55188 5 1 1 55187
0 55189 7 1 2 55107 55188
0 55190 5 1 1 55189
0 55191 7 1 2 69263 55190
0 55192 5 1 1 55191
0 55193 7 1 2 64302 55192
0 55194 7 1 2 55029 55193
0 55195 5 1 1 55194
0 55196 7 1 2 76197 55195
0 55197 7 1 2 54904 55196
0 55198 5 1 1 55197
0 55199 7 1 2 74508 100908
0 55200 5 1 1 55199
0 55201 7 1 2 70783 55200
0 55202 5 1 1 55201
0 55203 7 1 2 72679 86845
0 55204 5 1 1 55203
0 55205 7 1 2 94511 55204
0 55206 7 1 2 55202 55205
0 55207 5 1 1 55206
0 55208 7 1 2 68880 55207
0 55209 5 1 1 55208
0 55210 7 1 2 64012 101781
0 55211 5 1 1 55210
0 55212 7 1 2 103393 55211
0 55213 5 1 1 55212
0 55214 7 1 2 65875 55213
0 55215 5 1 1 55214
0 55216 7 1 2 103308 55215
0 55217 7 1 2 55209 55216
0 55218 5 2 1 55217
0 55219 7 1 2 65578 103472
0 55220 5 1 1 55219
0 55221 7 1 2 103317 55220
0 55222 5 1 1 55221
0 55223 7 1 2 70161 55222
0 55224 5 1 1 55223
0 55225 7 1 2 76953 96274
0 55226 5 1 1 55225
0 55227 7 1 2 55224 55226
0 55228 5 2 1 55227
0 55229 7 1 2 98530 103474
0 55230 5 1 1 55229
0 55231 7 2 2 76954 96976
0 55232 5 1 1 103476
0 55233 7 1 2 100324 101025
0 55234 7 1 2 99909 55233
0 55235 5 1 1 55234
0 55236 7 1 2 55232 55235
0 55237 5 1 1 55236
0 55238 7 1 2 62235 55237
0 55239 5 1 1 55238
0 55240 7 1 2 70513 101294
0 55241 7 2 2 103473 55240
0 55242 7 1 2 99379 103478
0 55243 5 1 1 55242
0 55244 7 1 2 55239 55243
0 55245 7 1 2 55230 55244
0 55246 5 1 1 55245
0 55247 7 1 2 100815 55246
0 55248 5 1 1 55247
0 55249 7 2 2 73745 84248
0 55250 5 2 1 103480
0 55251 7 1 2 90070 103482
0 55252 5 1 1 55251
0 55253 7 1 2 73507 55252
0 55254 5 1 1 55253
0 55255 7 3 2 73090 94522
0 55256 5 1 1 103484
0 55257 7 1 2 94411 55256
0 55258 5 3 1 55257
0 55259 7 1 2 67078 103487
0 55260 5 1 1 55259
0 55261 7 1 2 55254 55260
0 55262 5 1 1 55261
0 55263 7 1 2 55262 103226
0 55264 5 1 1 55263
0 55265 7 2 2 96364 103469
0 55266 5 10 1 103490
0 55267 7 1 2 100994 103492
0 55268 5 1 1 55267
0 55269 7 1 2 62684 101507
0 55270 5 1 1 55269
0 55271 7 3 2 85552 55270
0 55272 5 1 1 103502
0 55273 7 2 2 66052 103503
0 55274 7 1 2 74096 103505
0 55275 5 1 1 55274
0 55276 7 1 2 55268 55275
0 55277 5 1 1 55276
0 55278 7 1 2 65579 55277
0 55279 5 1 1 55278
0 55280 7 1 2 72740 55279
0 55281 5 1 1 55280
0 55282 7 1 2 55281 103236
0 55283 5 1 1 55282
0 55284 7 1 2 55264 55283
0 55285 5 1 1 55284
0 55286 7 1 2 70162 55285
0 55287 5 1 1 55286
0 55288 7 1 2 87503 94387
0 55289 7 2 2 94957 55288
0 55290 7 1 2 66330 103507
0 55291 5 1 1 55290
0 55292 7 1 2 80557 103237
0 55293 5 1 1 55292
0 55294 7 1 2 55291 55293
0 55295 5 1 1 55294
0 55296 7 1 2 80592 55295
0 55297 5 1 1 55296
0 55298 7 1 2 73360 103238
0 55299 7 1 2 103457 55298
0 55300 5 1 1 55299
0 55301 7 1 2 55297 55300
0 55302 7 1 2 55287 55301
0 55303 5 1 1 55302
0 55304 7 1 2 93886 55303
0 55305 5 1 1 55304
0 55306 7 1 2 64220 84953
0 55307 5 1 1 55306
0 55308 7 1 2 85954 55307
0 55309 5 1 1 55308
0 55310 7 1 2 70514 55309
0 55311 5 2 1 55310
0 55312 7 2 2 74140 75737
0 55313 5 2 1 103511
0 55314 7 1 2 103509 103513
0 55315 5 1 1 55314
0 55316 7 1 2 70974 55315
0 55317 5 1 1 55316
0 55318 7 1 2 55317 46652
0 55319 5 1 1 55318
0 55320 7 1 2 97320 55319
0 55321 5 1 1 55320
0 55322 7 1 2 100503 55321
0 55323 5 1 1 55322
0 55324 7 1 2 67079 55323
0 55325 5 1 1 55324
0 55326 7 1 2 86212 100509
0 55327 5 1 1 55326
0 55328 7 1 2 72860 88113
0 55329 5 1 1 55328
0 55330 7 1 2 67751 103481
0 55331 5 1 1 55330
0 55332 7 1 2 55329 55331
0 55333 5 3 1 55332
0 55334 7 1 2 97321 103515
0 55335 5 1 1 55334
0 55336 7 1 2 55327 55335
0 55337 5 1 1 55336
0 55338 7 1 2 73508 55337
0 55339 5 1 1 55338
0 55340 7 1 2 101034 100265
0 55341 5 1 1 55340
0 55342 7 1 2 55339 55341
0 55343 7 1 2 55325 55342
0 55344 5 1 1 55343
0 55345 7 1 2 70163 55344
0 55346 5 1 1 55345
0 55347 7 1 2 103477 103111
0 55348 5 1 1 55347
0 55349 7 1 2 96977 102401
0 55350 5 1 1 55349
0 55351 7 2 2 90882 99967
0 55352 7 1 2 76911 95182
0 55353 7 1 2 103518 55352
0 55354 5 1 1 55353
0 55355 7 1 2 55350 55354
0 55356 5 1 1 55355
0 55357 7 1 2 78352 55356
0 55358 5 1 1 55357
0 55359 7 1 2 55348 55358
0 55360 7 1 2 55346 55359
0 55361 5 1 1 55360
0 55362 7 1 2 100699 55361
0 55363 5 1 1 55362
0 55364 7 1 2 55305 55363
0 55365 7 1 2 55248 55364
0 55366 5 1 1 55365
0 55367 7 1 2 100681 55366
0 55368 5 1 1 55367
0 55369 7 1 2 102201 103475
0 55370 5 1 1 55369
0 55371 7 1 2 103479 103153
0 55372 5 1 1 55371
0 55373 7 2 2 70515 102233
0 55374 7 1 2 103520 100663
0 55375 5 1 1 55374
0 55376 7 1 2 90530 98147
0 55377 7 1 2 103363 55376
0 55378 5 1 1 55377
0 55379 7 1 2 55375 55378
0 55380 5 1 1 55379
0 55381 7 1 2 62236 55380
0 55382 5 1 1 55381
0 55383 7 1 2 55372 55382
0 55384 7 1 2 55370 55383
0 55385 5 1 1 55384
0 55386 7 1 2 99508 55385
0 55387 5 1 1 55386
0 55388 7 1 2 65580 55272
0 55389 5 1 1 55388
0 55390 7 2 2 49516 55389
0 55391 7 1 2 102202 103522
0 55392 5 1 1 55391
0 55393 7 1 2 81001 92970
0 55394 7 1 2 97999 55393
0 55395 7 1 2 99941 55394
0 55396 5 1 1 55395
0 55397 7 1 2 55392 55396
0 55398 5 1 1 55397
0 55399 7 1 2 90451 55398
0 55400 5 1 1 55399
0 55401 7 1 2 92420 101513
0 55402 5 1 1 55401
0 55403 7 1 2 90250 55402
0 55404 5 1 1 55403
0 55405 7 1 2 102203 55404
0 55406 5 1 1 55405
0 55407 7 1 2 67542 98143
0 55408 7 1 2 80683 55407
0 55409 7 1 2 103154 55408
0 55410 5 1 1 55409
0 55411 7 1 2 55406 55410
0 55412 5 1 1 55411
0 55413 7 1 2 100995 55412
0 55414 5 1 1 55413
0 55415 7 1 2 80558 102204
0 55416 5 1 1 55415
0 55417 7 1 2 101819 103135
0 55418 7 1 2 103506 55417
0 55419 5 1 1 55418
0 55420 7 1 2 55416 55419
0 55421 5 1 1 55420
0 55422 7 1 2 80593 55421
0 55423 5 1 1 55422
0 55424 7 1 2 55414 55423
0 55425 7 1 2 55400 55424
0 55426 5 1 1 55425
0 55427 7 1 2 100019 55426
0 55428 5 1 1 55427
0 55429 7 1 2 55387 55428
0 55430 5 1 1 55429
0 55431 7 1 2 87810 55430
0 55432 5 1 1 55431
0 55433 7 1 2 100020 100260
0 55434 5 1 1 55433
0 55435 7 1 2 95637 99509
0 55436 5 1 1 55435
0 55437 7 1 2 55434 55436
0 55438 5 1 1 55437
0 55439 7 1 2 66053 55438
0 55440 5 1 1 55439
0 55441 7 1 2 101567 55440
0 55442 5 1 1 55441
0 55443 7 1 2 97792 103155
0 55444 5 1 1 55443
0 55445 7 2 2 98156 100664
0 55446 5 1 1 103524
0 55447 7 1 2 55444 55446
0 55448 5 1 1 55447
0 55449 7 1 2 55442 55448
0 55450 5 1 1 55449
0 55451 7 1 2 65581 102507
0 55452 5 1 1 55451
0 55453 7 1 2 103510 55452
0 55454 5 1 1 55453
0 55455 7 1 2 70975 55454
0 55456 5 1 1 55455
0 55457 7 2 2 92326 97014
0 55458 5 1 1 103526
0 55459 7 1 2 55456 55458
0 55460 5 1 1 55459
0 55461 7 1 2 100021 55460
0 55462 5 1 1 55461
0 55463 7 1 2 99510 103485
0 55464 5 1 1 55463
0 55465 7 1 2 55462 55464
0 55466 5 1 1 55465
0 55467 7 1 2 103136 55466
0 55468 5 1 1 55467
0 55469 7 1 2 101361 53984
0 55470 5 1 1 55469
0 55471 7 1 2 102205 55470
0 55472 5 1 1 55471
0 55473 7 1 2 55468 55472
0 55474 5 1 1 55473
0 55475 7 1 2 67080 55474
0 55476 5 1 1 55475
0 55477 7 1 2 55450 55476
0 55478 5 1 1 55477
0 55479 7 1 2 70164 55478
0 55480 5 1 1 55479
0 55481 7 1 2 103516 103137
0 55482 5 1 1 55481
0 55483 7 1 2 86750 102206
0 55484 5 1 1 55483
0 55485 7 1 2 55482 55484
0 55486 5 1 1 55485
0 55487 7 1 2 100022 55486
0 55488 5 1 1 55487
0 55489 7 1 2 73665 18493
0 55490 5 1 1 55489
0 55491 7 1 2 99511 102207
0 55492 7 1 2 55490 55491
0 55493 5 1 1 55492
0 55494 7 1 2 55488 55493
0 55495 5 1 1 55494
0 55496 7 1 2 70165 55495
0 55497 5 1 1 55496
0 55498 7 1 2 62237 103348
0 55499 5 1 1 55498
0 55500 7 1 2 72861 94971
0 55501 5 1 1 55500
0 55502 7 1 2 55499 55501
0 55503 5 1 1 55502
0 55504 7 1 2 99512 103138
0 55505 7 1 2 55503 55504
0 55506 5 1 1 55505
0 55507 7 1 2 55497 55506
0 55508 5 1 1 55507
0 55509 7 1 2 73509 55508
0 55510 5 1 1 55509
0 55511 7 1 2 75646 102208
0 55512 5 1 1 55511
0 55513 7 1 2 100849 55512
0 55514 5 1 1 55513
0 55515 7 1 2 62927 55514
0 55516 5 1 1 55515
0 55517 7 1 2 77992 102209
0 55518 5 1 1 55517
0 55519 7 1 2 55518 100850
0 55520 5 1 1 55519
0 55521 7 1 2 71384 55520
0 55522 5 1 1 55521
0 55523 7 1 2 101333 100846
0 55524 7 1 2 102129 55523
0 55525 5 1 1 55524
0 55526 7 1 2 55522 55525
0 55527 7 1 2 55516 55526
0 55528 5 1 1 55527
0 55529 7 1 2 99513 55528
0 55530 5 1 1 55529
0 55531 7 2 2 90983 99030
0 55532 7 1 2 95157 103528
0 55533 7 1 2 103158 55532
0 55534 5 1 1 55533
0 55535 7 1 2 55530 55534
0 55536 5 1 1 55535
0 55537 7 1 2 70516 55536
0 55538 5 1 1 55537
0 55539 7 1 2 66331 96908
0 55540 5 1 1 55539
0 55541 7 1 2 101362 55540
0 55542 5 1 1 55541
0 55543 7 1 2 100665 98636
0 55544 7 1 2 55542 55543
0 55545 5 1 1 55544
0 55546 7 1 2 55538 55545
0 55547 5 1 1 55546
0 55548 7 1 2 65252 55547
0 55549 5 1 1 55548
0 55550 7 1 2 55510 55549
0 55551 7 1 2 55480 55550
0 55552 5 1 1 55551
0 55553 7 1 2 87755 55552
0 55554 5 1 1 55553
0 55555 7 1 2 55432 55554
0 55556 7 1 2 55368 55555
0 55557 5 1 1 55556
0 55558 7 1 2 79187 55557
0 55559 5 1 1 55558
0 55560 7 1 2 65582 95995
0 55561 5 1 1 55560
0 55562 7 1 2 62238 55561
0 55563 5 1 1 55562
0 55564 7 1 2 96758 55563
0 55565 5 1 1 55564
0 55566 7 1 2 78283 96381
0 55567 5 1 1 55566
0 55568 7 1 2 87167 95243
0 55569 5 1 1 55568
0 55570 7 1 2 80081 83354
0 55571 5 1 1 55570
0 55572 7 1 2 55569 55571
0 55573 5 1 1 55572
0 55574 7 1 2 65583 55573
0 55575 5 1 1 55574
0 55576 7 1 2 55567 55575
0 55577 7 1 2 55565 55576
0 55578 5 1 1 55577
0 55579 7 2 2 101309 55578
0 55580 7 1 2 96952 103530
0 55581 5 1 1 55580
0 55582 7 1 2 70517 87127
0 55583 5 1 1 55582
0 55584 7 1 2 92870 55583
0 55585 5 1 1 55584
0 55586 7 1 2 64221 55585
0 55587 5 1 1 55586
0 55588 7 1 2 85349 101271
0 55589 5 1 1 55588
0 55590 7 1 2 55587 55589
0 55591 5 1 1 55590
0 55592 7 1 2 78284 55591
0 55593 5 1 1 55592
0 55594 7 1 2 76603 5422
0 55595 5 1 1 55594
0 55596 7 1 2 73510 55595
0 55597 5 1 1 55596
0 55598 7 1 2 27912 55597
0 55599 5 1 1 55598
0 55600 7 1 2 83355 55599
0 55601 5 1 1 55600
0 55602 7 1 2 55593 55601
0 55603 5 1 1 55602
0 55604 7 2 2 102362 55603
0 55605 7 1 2 100466 103532
0 55606 5 1 1 55605
0 55607 7 1 2 55581 55606
0 55608 5 1 1 55607
0 55609 7 1 2 70976 55608
0 55610 5 1 1 55609
0 55611 7 2 2 98828 103148
0 55612 7 2 2 78624 103534
0 55613 7 1 2 86900 103536
0 55614 5 1 1 55613
0 55615 7 2 2 79106 98531
0 55616 7 1 2 79666 103538
0 55617 5 1 1 55616
0 55618 7 2 2 65253 97322
0 55619 7 1 2 97202 101827
0 55620 5 1 1 55619
0 55621 7 1 2 75309 86230
0 55622 5 1 1 55621
0 55623 7 1 2 55620 55622
0 55624 5 1 1 55623
0 55625 7 1 2 61919 55624
0 55626 5 1 1 55625
0 55627 7 1 2 76256 85927
0 55628 7 1 2 95496 55627
0 55629 5 1 1 55628
0 55630 7 1 2 55626 55629
0 55631 5 1 1 55630
0 55632 7 1 2 103540 55631
0 55633 5 1 1 55632
0 55634 7 1 2 55617 55633
0 55635 5 1 1 55634
0 55636 7 1 2 66054 55635
0 55637 5 1 1 55636
0 55638 7 1 2 55614 55637
0 55639 5 1 1 55638
0 55640 7 1 2 73511 55639
0 55641 5 1 1 55640
0 55642 7 1 2 91215 103539
0 55643 5 1 1 55642
0 55644 7 1 2 74133 83356
0 55645 5 2 1 55644
0 55646 7 1 2 7522 103542
0 55647 5 1 1 55646
0 55648 7 1 2 80286 103541
0 55649 7 1 2 55647 55648
0 55650 5 1 1 55649
0 55651 7 1 2 55643 55650
0 55652 5 1 1 55651
0 55653 7 1 2 65584 55652
0 55654 5 1 1 55653
0 55655 7 1 2 74161 100495
0 55656 7 1 2 99825 103097
0 55657 7 1 2 55655 55656
0 55658 5 1 1 55657
0 55659 7 1 2 55654 55658
0 55660 5 1 1 55659
0 55661 7 1 2 71385 55660
0 55662 5 1 1 55661
0 55663 7 1 2 92392 96978
0 55664 5 1 1 55663
0 55665 7 1 2 77042 97323
0 55666 7 1 2 100261 55665
0 55667 5 1 1 55666
0 55668 7 1 2 55664 55667
0 55669 5 1 1 55668
0 55670 7 1 2 73657 55669
0 55671 5 1 1 55670
0 55672 7 2 2 73361 99330
0 55673 7 1 2 65585 103459
0 55674 7 1 2 103544 55673
0 55675 5 1 1 55674
0 55676 7 1 2 55671 55675
0 55677 5 1 1 55676
0 55678 7 1 2 78285 55677
0 55679 5 1 1 55678
0 55680 7 1 2 55662 55679
0 55681 7 1 2 55641 55680
0 55682 7 1 2 55610 55681
0 55683 5 1 1 55682
0 55684 7 1 2 99728 55683
0 55685 5 1 1 55684
0 55686 7 1 2 66055 102728
0 55687 5 2 1 55686
0 55688 7 3 2 64809 77686
0 55689 7 1 2 84178 103548
0 55690 5 1 1 55689
0 55691 7 1 2 103546 55690
0 55692 5 1 1 55691
0 55693 7 1 2 61920 55692
0 55694 5 1 1 55693
0 55695 7 3 2 76026 77459
0 55696 7 1 2 69866 103551
0 55697 5 2 1 55696
0 55698 7 1 2 77100 77954
0 55699 5 1 1 55698
0 55700 7 1 2 103554 55699
0 55701 5 2 1 55700
0 55702 7 1 2 78269 103556
0 55703 5 1 1 55702
0 55704 7 1 2 55694 55703
0 55705 5 1 1 55704
0 55706 7 1 2 73512 55705
0 55707 5 1 1 55706
0 55708 7 2 2 76852 78270
0 55709 5 1 1 103558
0 55710 7 1 2 74097 103559
0 55711 5 1 1 55710
0 55712 7 1 2 74251 82402
0 55713 5 1 1 55712
0 55714 7 1 2 55711 55713
0 55715 5 1 1 55714
0 55716 7 1 2 70518 55715
0 55717 5 1 1 55716
0 55718 7 1 2 95008 103543
0 55719 5 1 1 55718
0 55720 7 1 2 71712 55719
0 55721 5 1 1 55720
0 55722 7 1 2 71266 73588
0 55723 5 2 1 55722
0 55724 7 1 2 73783 79107
0 55725 7 1 2 103560 55724
0 55726 5 1 1 55725
0 55727 7 1 2 55721 55726
0 55728 5 1 1 55727
0 55729 7 1 2 65586 55728
0 55730 5 1 1 55729
0 55731 7 1 2 55717 55730
0 55732 5 2 1 55731
0 55733 7 1 2 62239 103562
0 55734 5 1 1 55733
0 55735 7 1 2 55707 55734
0 55736 5 1 1 55735
0 55737 7 1 2 99787 102363
0 55738 7 1 2 55736 55737
0 55739 5 1 1 55738
0 55740 7 1 2 55685 55739
0 55741 5 1 1 55740
0 55742 7 1 2 64411 55741
0 55743 5 1 1 55742
0 55744 7 1 2 5578 1587
0 55745 5 2 1 55744
0 55746 7 1 2 79188 99333
0 55747 5 1 1 55746
0 55748 7 1 2 98532 98934
0 55749 5 1 1 55748
0 55750 7 1 2 55747 55749
0 55751 5 1 1 55750
0 55752 7 1 2 70166 55751
0 55753 5 1 1 55752
0 55754 7 1 2 75488 92652
0 55755 7 1 2 101149 55754
0 55756 7 1 2 86592 55755
0 55757 5 1 1 55756
0 55758 7 1 2 55753 55757
0 55759 5 1 1 55758
0 55760 7 1 2 103564 55759
0 55761 5 1 1 55760
0 55762 7 1 2 102029 102509
0 55763 5 1 1 55762
0 55764 7 1 2 61921 102290
0 55765 5 1 1 55764
0 55766 7 1 2 78271 102262
0 55767 5 1 1 55766
0 55768 7 1 2 55765 55767
0 55769 5 1 1 55768
0 55770 7 1 2 92653 98045
0 55771 7 1 2 55769 55770
0 55772 5 1 1 55771
0 55773 7 1 2 55763 55772
0 55774 5 1 1 55773
0 55775 7 1 2 77907 55774
0 55776 5 1 1 55775
0 55777 7 1 2 55761 55776
0 55778 5 1 1 55777
0 55779 7 1 2 64412 55778
0 55780 5 1 1 55779
0 55781 7 1 2 80594 99126
0 55782 7 1 2 79189 55781
0 55783 7 1 2 98425 55782
0 55784 5 1 1 55783
0 55785 7 1 2 55780 55784
0 55786 5 1 1 55785
0 55787 7 1 2 99729 55786
0 55788 5 1 1 55787
0 55789 7 1 2 97298 102307
0 55790 7 2 2 100238 55789
0 55791 7 1 2 92654 103566
0 55792 5 1 1 55791
0 55793 7 1 2 70167 79190
0 55794 7 1 2 102311 55793
0 55795 5 1 1 55794
0 55796 7 1 2 55792 55795
0 55797 5 1 1 55796
0 55798 7 1 2 71267 55797
0 55799 5 1 1 55798
0 55800 7 1 2 103455 103535
0 55801 5 1 1 55800
0 55802 7 1 2 55799 55801
0 55803 5 1 1 55802
0 55804 7 1 2 65876 55803
0 55805 5 1 1 55804
0 55806 7 1 2 92521 103537
0 55807 5 1 1 55806
0 55808 7 1 2 55805 55807
0 55809 5 1 1 55808
0 55810 7 1 2 55809 100716
0 55811 5 1 1 55810
0 55812 7 1 2 55788 55811
0 55813 5 1 1 55812
0 55814 7 1 2 72211 55813
0 55815 5 1 1 55814
0 55816 7 2 2 75489 80304
0 55817 7 1 2 87917 103568
0 55818 5 1 1 55817
0 55819 7 1 2 100239 101183
0 55820 5 1 1 55819
0 55821 7 1 2 55818 55820
0 55822 5 1 1 55821
0 55823 7 1 2 66056 55822
0 55824 5 1 1 55823
0 55825 7 2 2 76853 73616
0 55826 7 1 2 85909 103570
0 55827 5 1 1 55826
0 55828 7 1 2 55824 55827
0 55829 5 1 1 55828
0 55830 7 1 2 69070 55829
0 55831 5 1 1 55830
0 55832 7 1 2 72680 103007
0 55833 5 2 1 55832
0 55834 7 1 2 103397 103572
0 55835 5 1 1 55834
0 55836 7 1 2 103569 55835
0 55837 5 1 1 55836
0 55838 7 1 2 55831 55837
0 55839 5 1 1 55838
0 55840 7 1 2 65877 55839
0 55841 5 2 1 55840
0 55842 7 1 2 86412 89645
0 55843 5 1 1 55842
0 55844 7 1 2 101354 55843
0 55845 5 1 1 55844
0 55846 7 1 2 70519 55845
0 55847 5 1 1 55846
0 55848 7 1 2 89746 93395
0 55849 5 1 1 55848
0 55850 7 1 2 62928 55849
0 55851 5 1 1 55850
0 55852 7 1 2 62685 296
0 55853 7 1 2 95174 55852
0 55854 7 1 2 12171 55853
0 55855 5 1 1 55854
0 55856 7 1 2 55851 55855
0 55857 7 1 2 55847 55856
0 55858 5 1 1 55857
0 55859 7 1 2 70784 55858
0 55860 5 1 1 55859
0 55861 7 1 2 84578 86491
0 55862 5 2 1 55861
0 55863 7 1 2 55860 103576
0 55864 5 1 1 55863
0 55865 7 1 2 81235 55864
0 55866 5 1 1 55865
0 55867 7 1 2 103574 55866
0 55868 5 1 1 55867
0 55869 7 1 2 69638 55868
0 55870 5 1 1 55869
0 55871 7 1 2 95795 95980
0 55872 5 1 1 55871
0 55873 7 1 2 89783 55872
0 55874 5 1 1 55873
0 55875 7 1 2 94433 95716
0 55876 5 1 1 55875
0 55877 7 1 2 73666 48713
0 55878 5 1 1 55877
0 55879 7 1 2 71386 55878
0 55880 5 1 1 55879
0 55881 7 1 2 55876 55880
0 55882 7 1 2 55874 55881
0 55883 5 1 1 55882
0 55884 7 1 2 85985 55883
0 55885 5 1 1 55884
0 55886 7 1 2 55870 55885
0 55887 5 1 1 55886
0 55888 7 1 2 65254 55887
0 55889 5 1 1 55888
0 55890 7 1 2 79159 55709
0 55891 5 3 1 55890
0 55892 7 1 2 76499 103578
0 55893 5 1 1 55892
0 55894 7 2 2 83345 80352
0 55895 5 1 1 103581
0 55896 7 1 2 95009 55895
0 55897 5 1 1 55896
0 55898 7 1 2 84548 55897
0 55899 5 1 1 55898
0 55900 7 1 2 55893 55899
0 55901 5 1 1 55900
0 55902 7 1 2 62686 55901
0 55903 5 1 1 55902
0 55904 7 1 2 76502 103579
0 55905 5 1 1 55904
0 55906 7 1 2 55903 55905
0 55907 5 1 1 55906
0 55908 7 1 2 65587 77672
0 55909 7 2 2 55907 55908
0 55910 5 1 1 103583
0 55911 7 1 2 55889 55910
0 55912 5 1 1 55911
0 55913 7 1 2 97324 100816
0 55914 7 1 2 55912 55913
0 55915 5 1 1 55914
0 55916 7 1 2 55815 55915
0 55917 7 1 2 55743 55916
0 55918 5 1 1 55917
0 55919 7 1 2 100682 55918
0 55920 5 1 1 55919
0 55921 7 2 2 98117 103345
0 55922 7 1 2 73513 103585
0 55923 5 1 1 55922
0 55924 7 2 2 89672 102391
0 55925 7 1 2 87828 97641
0 55926 7 1 2 103587 55925
0 55927 5 1 1 55926
0 55928 7 1 2 55923 55927
0 55929 5 1 1 55928
0 55930 7 1 2 70168 55929
0 55931 5 1 1 55930
0 55932 7 1 2 95289 100641
0 55933 7 1 2 100632 55932
0 55934 7 1 2 103588 55933
0 55935 5 1 1 55934
0 55936 7 1 2 55931 55935
0 55937 5 1 1 55936
0 55938 7 1 2 70785 55937
0 55939 5 1 1 55938
0 55940 7 1 2 71387 78204
0 55941 7 1 2 103586 55940
0 55942 5 1 1 55941
0 55943 7 1 2 55939 55942
0 55944 5 1 1 55943
0 55945 7 1 2 65003 55944
0 55946 5 1 1 55945
0 55947 7 2 2 79301 97552
0 55948 7 1 2 68049 99195
0 55949 7 1 2 97347 55948
0 55950 7 1 2 98287 55949
0 55951 7 1 2 103589 55950
0 55952 5 1 1 55951
0 55953 7 1 2 55946 55952
0 55954 5 1 1 55953
0 55955 7 1 2 66785 55954
0 55956 5 1 1 55955
0 55957 7 2 2 93007 99369
0 55958 7 1 2 69071 98162
0 55959 7 1 2 90519 55958
0 55960 7 1 2 103591 55959
0 55961 7 1 2 103590 55960
0 55962 5 1 1 55961
0 55963 7 1 2 65588 55962
0 55964 7 1 2 55956 55963
0 55965 5 1 1 55964
0 55966 7 1 2 87756 100262
0 55967 5 1 1 55966
0 55968 7 2 2 87811 103493
0 55969 5 1 1 103593
0 55970 7 1 2 72808 103594
0 55971 5 1 1 55970
0 55972 7 1 2 55967 55971
0 55973 5 1 1 55972
0 55974 7 1 2 77043 55973
0 55975 5 1 1 55974
0 55976 7 2 2 99968 103012
0 55977 5 1 1 103595
0 55978 7 1 2 72809 103596
0 55979 5 1 1 55978
0 55980 7 1 2 55975 55979
0 55981 5 1 1 55980
0 55982 7 1 2 103139 55981
0 55983 5 1 1 55982
0 55984 7 1 2 92542 99798
0 55985 7 1 2 87770 55984
0 55986 7 1 2 98127 55985
0 55987 5 1 1 55986
0 55988 7 1 2 55983 55987
0 55989 5 1 1 55988
0 55990 7 1 2 78852 55989
0 55991 5 1 1 55990
0 55992 7 1 2 70520 55991
0 55993 5 1 1 55992
0 55994 7 1 2 69639 55993
0 55995 7 1 2 55965 55994
0 55996 5 1 1 55995
0 55997 7 1 2 55969 97545
0 55998 5 1 1 55997
0 55999 7 1 2 77044 55998
0 56000 5 1 1 55999
0 56001 7 1 2 55977 56000
0 56002 5 1 1 56001
0 56003 7 1 2 64222 56002
0 56004 5 1 1 56003
0 56005 7 1 2 65255 90848
0 56006 7 1 2 102386 56005
0 56007 5 1 1 56006
0 56008 7 1 2 56004 56007
0 56009 5 1 1 56008
0 56010 7 1 2 70521 56009
0 56011 5 1 1 56010
0 56012 7 1 2 87879 102588
0 56013 7 1 2 102368 56012
0 56014 5 1 1 56013
0 56015 7 1 2 56011 56014
0 56016 5 1 1 56015
0 56017 7 1 2 79151 103140
0 56018 7 1 2 56016 56017
0 56019 5 1 1 56018
0 56020 7 1 2 55996 56019
0 56021 5 1 1 56020
0 56022 7 1 2 66057 56021
0 56023 5 1 1 56022
0 56024 7 1 2 86383 101514
0 56025 5 1 1 56024
0 56026 7 1 2 99709 56025
0 56027 5 1 1 56026
0 56028 7 1 2 77045 56027
0 56029 5 1 1 56028
0 56030 7 1 2 67543 102684
0 56031 5 1 1 56030
0 56032 7 1 2 99710 56031
0 56033 5 1 1 56032
0 56034 7 1 2 77673 56033
0 56035 5 1 1 56034
0 56036 7 1 2 56029 56035
0 56037 5 1 1 56036
0 56038 7 2 2 71180 87812
0 56039 7 1 2 79152 103597
0 56040 7 1 2 56037 56039
0 56041 5 1 1 56040
0 56042 7 1 2 78286 103527
0 56043 5 1 1 56042
0 56044 7 1 2 73514 86901
0 56045 5 1 1 56044
0 56046 7 1 2 103514 56045
0 56047 5 1 1 56046
0 56048 7 1 2 83357 56047
0 56049 5 1 1 56048
0 56050 7 1 2 56043 56049
0 56051 5 1 1 56050
0 56052 7 1 2 95307 99283
0 56053 7 1 2 56051 56052
0 56054 5 1 1 56053
0 56055 7 1 2 56041 56054
0 56056 5 1 1 56055
0 56057 7 1 2 103141 56056
0 56058 5 1 1 56057
0 56059 7 1 2 100666 103531
0 56060 5 1 1 56059
0 56061 7 1 2 102301 103533
0 56062 5 1 1 56061
0 56063 7 1 2 56060 56062
0 56064 5 1 1 56063
0 56065 7 1 2 87757 56064
0 56066 5 1 1 56065
0 56067 7 1 2 67544 76599
0 56068 5 2 1 56067
0 56069 7 1 2 64223 72936
0 56070 5 1 1 56069
0 56071 7 1 2 103599 56070
0 56072 5 1 1 56071
0 56073 7 1 2 83358 56072
0 56074 5 1 1 56073
0 56075 7 1 2 78287 102037
0 56076 5 1 1 56075
0 56077 7 1 2 56074 56076
0 56078 5 1 1 56077
0 56079 7 1 2 77360 56078
0 56080 5 1 1 56079
0 56081 7 1 2 79153 1753
0 56082 7 1 2 101577 56081
0 56083 5 1 1 56082
0 56084 7 2 2 71181 79108
0 56085 5 1 1 103601
0 56086 7 1 2 62687 103602
0 56087 5 1 1 56086
0 56088 7 1 2 56083 56087
0 56089 5 1 1 56088
0 56090 7 1 2 73137 56089
0 56091 5 1 1 56090
0 56092 7 1 2 89292 86465
0 56093 7 1 2 96756 56092
0 56094 5 1 1 56093
0 56095 7 1 2 56091 56094
0 56096 7 1 2 56080 56095
0 56097 5 1 1 56096
0 56098 7 1 2 80595 56097
0 56099 5 1 1 56098
0 56100 7 1 2 69072 79154
0 56101 5 1 1 56100
0 56102 7 1 2 56085 56101
0 56103 5 1 1 56102
0 56104 7 1 2 72893 103460
0 56105 7 1 2 56103 56104
0 56106 5 1 1 56105
0 56107 7 1 2 56099 56106
0 56108 5 1 1 56107
0 56109 7 1 2 97325 103075
0 56110 7 1 2 56108 56109
0 56111 5 1 1 56110
0 56112 7 1 2 56066 56111
0 56113 5 1 1 56112
0 56114 7 1 2 70977 56113
0 56115 5 1 1 56114
0 56116 7 1 2 56058 56115
0 56117 7 1 2 56023 56116
0 56118 5 1 1 56117
0 56119 7 1 2 100023 56118
0 56120 5 1 1 56119
0 56121 7 1 2 99521 37006
0 56122 5 2 1 56121
0 56123 7 1 2 103523 103603
0 56124 5 1 1 56123
0 56125 7 1 2 103451 103029
0 56126 5 1 1 56125
0 56127 7 1 2 56124 56126
0 56128 5 1 1 56127
0 56129 7 1 2 66058 56128
0 56130 5 1 1 56129
0 56131 7 1 2 103494 103035
0 56132 5 1 1 56131
0 56133 7 1 2 77361 99993
0 56134 5 1 1 56133
0 56135 7 1 2 56132 56134
0 56136 5 1 1 56135
0 56137 7 1 2 84023 56136
0 56138 5 1 1 56137
0 56139 7 1 2 56130 56138
0 56140 5 1 1 56139
0 56141 7 1 2 69073 56140
0 56142 5 1 1 56141
0 56143 7 1 2 64224 100024
0 56144 7 1 2 101653 56143
0 56145 5 1 1 56144
0 56146 7 1 2 101363 56145
0 56147 5 1 1 56146
0 56148 7 1 2 103495 56147
0 56149 5 1 1 56148
0 56150 7 1 2 79686 99514
0 56151 7 1 2 103395 56150
0 56152 5 1 1 56151
0 56153 7 1 2 56149 56152
0 56154 5 1 1 56153
0 56155 7 1 2 65589 56154
0 56156 5 1 1 56155
0 56157 7 1 2 56142 56156
0 56158 5 1 1 56157
0 56159 7 1 2 97746 56158
0 56160 5 1 1 56159
0 56161 7 1 2 102323 103517
0 56162 5 1 1 56161
0 56163 7 1 2 96416 97728
0 56164 7 1 2 102899 56163
0 56165 5 1 1 56164
0 56166 7 1 2 66188 83467
0 56167 7 1 2 99266 56166
0 56168 5 1 1 56167
0 56169 7 1 2 56165 56168
0 56170 5 1 1 56169
0 56171 7 1 2 65590 56170
0 56172 5 1 1 56171
0 56173 7 3 2 70522 100035
0 56174 5 1 1 103605
0 56175 7 1 2 64225 103606
0 56176 5 1 1 56175
0 56177 7 1 2 56172 56176
0 56178 5 1 1 56177
0 56179 7 1 2 99515 56178
0 56180 5 1 1 56179
0 56181 7 1 2 56162 56180
0 56182 5 1 1 56181
0 56183 7 1 2 73515 56182
0 56184 5 1 1 56183
0 56185 7 1 2 84911 100997
0 56186 5 1 1 56185
0 56187 7 1 2 70523 56186
0 56188 5 1 1 56187
0 56189 7 1 2 103160 56188
0 56190 5 2 1 56189
0 56191 7 1 2 100025 103608
0 56192 5 1 1 56191
0 56193 7 1 2 99516 103488
0 56194 5 1 1 56193
0 56195 7 1 2 56192 56194
0 56196 5 1 1 56195
0 56197 7 1 2 100036 56196
0 56198 5 1 1 56197
0 56199 7 1 2 56184 56198
0 56200 7 1 2 56160 56199
0 56201 5 1 1 56200
0 56202 7 1 2 70169 56201
0 56203 5 1 1 56202
0 56204 7 1 2 91003 103508
0 56205 5 1 1 56204
0 56206 7 1 2 80559 100026
0 56207 5 1 1 56206
0 56208 7 1 2 33831 56207
0 56209 5 1 1 56208
0 56210 7 1 2 97747 56209
0 56211 5 1 1 56210
0 56212 7 1 2 56205 56211
0 56213 5 1 1 56212
0 56214 7 1 2 80596 56213
0 56215 5 1 1 56214
0 56216 7 1 2 76955 97748
0 56217 7 1 2 103122 56216
0 56218 5 1 1 56217
0 56219 7 1 2 56215 56218
0 56220 7 1 2 56203 56219
0 56221 5 1 1 56220
0 56222 7 1 2 79191 56221
0 56223 5 1 1 56222
0 56224 7 1 2 76999 103549
0 56225 5 1 1 56224
0 56226 7 1 2 56225 29519
0 56227 5 2 1 56226
0 56228 7 1 2 99517 103610
0 56229 5 1 1 56228
0 56230 7 1 2 73954 103580
0 56231 5 1 1 56230
0 56232 7 1 2 66059 83359
0 56233 5 1 1 56232
0 56234 7 1 2 56231 56233
0 56235 5 1 1 56234
0 56236 7 1 2 103212 56235
0 56237 5 1 1 56236
0 56238 7 1 2 56229 56237
0 56239 5 1 1 56238
0 56240 7 1 2 64226 56239
0 56241 5 1 1 56240
0 56242 7 1 2 69074 98092
0 56243 7 1 2 84185 56242
0 56244 7 1 2 101196 56243
0 56245 5 1 1 56244
0 56246 7 1 2 56241 56245
0 56247 5 1 1 56246
0 56248 7 1 2 62240 56247
0 56249 5 1 1 56248
0 56250 7 1 2 80103 84203
0 56251 7 1 2 100240 56250
0 56252 7 1 2 103604 56251
0 56253 5 1 1 56252
0 56254 7 1 2 56249 56253
0 56255 5 1 1 56254
0 56256 7 1 2 73516 56255
0 56257 5 1 1 56256
0 56258 7 1 2 95010 44373
0 56259 5 1 1 56258
0 56260 7 1 2 71388 56259
0 56261 5 1 1 56260
0 56262 7 1 2 79090 75613
0 56263 5 1 1 56262
0 56264 7 1 2 56261 56263
0 56265 5 1 1 56264
0 56266 7 1 2 65591 56265
0 56267 5 1 1 56266
0 56268 7 1 2 71268 103611
0 56269 5 1 1 56268
0 56270 7 1 2 69640 75689
0 56271 7 1 2 80317 56270
0 56272 5 1 1 56271
0 56273 7 1 2 56269 56272
0 56274 7 1 2 56267 56273
0 56275 5 1 1 56274
0 56276 7 1 2 70978 56275
0 56277 5 1 1 56276
0 56278 7 1 2 90298 101715
0 56279 5 1 1 56278
0 56280 7 1 2 79160 34301
0 56281 5 1 1 56280
0 56282 7 1 2 97015 56281
0 56283 5 1 1 56282
0 56284 7 1 2 56279 56283
0 56285 7 1 2 56277 56284
0 56286 5 1 1 56285
0 56287 7 1 2 64227 56286
0 56288 5 1 1 56287
0 56289 7 1 2 83346 101840
0 56290 5 1 1 56289
0 56291 7 1 2 7432 56290
0 56292 5 1 1 56291
0 56293 7 1 2 73091 56292
0 56294 5 1 1 56293
0 56295 7 1 2 79155 74720
0 56296 5 1 1 56295
0 56297 7 1 2 56294 56296
0 56298 5 1 1 56297
0 56299 7 1 2 71389 56298
0 56300 5 1 1 56299
0 56301 7 1 2 87991 91730
0 56302 5 1 1 56301
0 56303 7 1 2 76600 56302
0 56304 5 1 1 56303
0 56305 7 1 2 73527 56304
0 56306 5 1 1 56305
0 56307 7 1 2 78288 56306
0 56308 5 1 1 56307
0 56309 7 1 2 56300 56308
0 56310 7 1 2 56288 56309
0 56311 5 1 1 56310
0 56312 7 1 2 100027 56311
0 56313 5 1 1 56312
0 56314 7 1 2 99518 103563
0 56315 5 1 1 56314
0 56316 7 1 2 56313 56315
0 56317 5 1 1 56316
0 56318 7 1 2 62241 56317
0 56319 5 1 1 56318
0 56320 7 1 2 56257 56319
0 56321 5 1 1 56320
0 56322 7 1 2 56321 99921
0 56323 5 1 1 56322
0 56324 7 1 2 56223 56323
0 56325 5 1 1 56324
0 56326 7 1 2 100594 56325
0 56327 5 1 1 56326
0 56328 7 1 2 100756 98341
0 56329 7 1 2 101489 56328
0 56330 5 1 1 56329
0 56331 7 1 2 78434 100654
0 56332 7 1 2 102303 56331
0 56333 5 1 1 56332
0 56334 7 1 2 56330 56333
0 56335 5 1 1 56334
0 56336 7 1 2 70170 56335
0 56337 5 1 1 56336
0 56338 7 1 2 63207 87675
0 56339 7 1 2 103521 56338
0 56340 7 1 2 103529 56339
0 56341 5 1 1 56340
0 56342 7 1 2 56337 56341
0 56343 5 1 1 56342
0 56344 7 1 2 87813 56343
0 56345 5 1 1 56344
0 56346 7 2 2 71269 81715
0 56347 7 1 2 99923 103612
0 56348 5 1 1 56347
0 56349 7 1 2 97729 97437
0 56350 7 1 2 80597 56349
0 56351 5 1 1 56350
0 56352 7 1 2 56348 56351
0 56353 5 1 1 56352
0 56354 7 1 2 100028 56353
0 56355 5 1 1 56354
0 56356 7 1 2 82891 86281
0 56357 7 1 2 100837 56356
0 56358 5 1 1 56357
0 56359 7 1 2 56355 56358
0 56360 5 1 1 56359
0 56361 7 1 2 100595 56360
0 56362 5 1 1 56361
0 56363 7 1 2 68881 77385
0 56364 7 1 2 81522 56363
0 56365 7 2 2 61327 76729
0 56366 7 1 2 91888 102320
0 56367 7 1 2 103614 56366
0 56368 7 1 2 56364 56367
0 56369 5 1 1 56368
0 56370 7 1 2 56362 56369
0 56371 7 1 2 56345 56370
0 56372 5 1 1 56371
0 56373 7 1 2 79192 56372
0 56374 5 1 1 56373
0 56375 7 1 2 78272 102265
0 56376 5 1 1 56375
0 56377 7 1 2 75426 94902
0 56378 5 1 1 56377
0 56379 7 1 2 56376 56378
0 56380 5 1 1 56379
0 56381 7 1 2 97793 100605
0 56382 7 1 2 56380 56381
0 56383 5 1 1 56382
0 56384 7 1 2 61328 82011
0 56385 7 1 2 83600 56384
0 56386 7 1 2 103525 56385
0 56387 5 1 1 56386
0 56388 7 1 2 56383 56387
0 56389 5 1 1 56388
0 56390 7 1 2 102297 56389
0 56391 5 1 1 56390
0 56392 7 1 2 67752 83785
0 56393 7 1 2 93755 56392
0 56394 7 1 2 97255 99826
0 56395 7 1 2 101143 56394
0 56396 7 1 2 56393 56395
0 56397 5 1 1 56396
0 56398 7 1 2 56391 56397
0 56399 5 1 1 56398
0 56400 7 1 2 103565 56399
0 56401 5 1 1 56400
0 56402 7 1 2 102298 100596
0 56403 5 1 1 56402
0 56404 7 2 2 98479 102244
0 56405 7 1 2 92819 99991
0 56406 7 1 2 103616 56405
0 56407 5 1 1 56406
0 56408 7 1 2 56403 56407
0 56409 5 1 1 56408
0 56410 7 1 2 66189 56409
0 56411 5 1 1 56410
0 56412 7 1 2 102271 103617
0 56413 5 1 1 56412
0 56414 7 1 2 56411 56413
0 56415 5 1 1 56414
0 56416 7 1 2 103567 56415
0 56417 5 1 1 56416
0 56418 7 1 2 93141 99065
0 56419 7 1 2 102030 56418
0 56420 7 1 2 100656 103143
0 56421 7 1 2 56419 56420
0 56422 5 1 1 56421
0 56423 7 1 2 56417 56422
0 56424 5 1 1 56423
0 56425 7 1 2 77908 56424
0 56426 5 1 1 56425
0 56427 7 1 2 56401 56426
0 56428 7 1 2 56374 56427
0 56429 5 1 1 56428
0 56430 7 1 2 72212 56429
0 56431 5 1 1 56430
0 56432 7 1 2 77502 87758
0 56433 5 1 1 56432
0 56434 7 1 2 94136 99428
0 56435 5 1 1 56434
0 56436 7 1 2 56433 56435
0 56437 5 1 1 56436
0 56438 7 1 2 65592 56437
0 56439 5 1 1 56438
0 56440 7 1 2 72884 103201
0 56441 5 1 1 56440
0 56442 7 1 2 56439 56441
0 56443 5 1 1 56442
0 56444 7 1 2 71390 56443
0 56445 5 1 1 56444
0 56446 7 1 2 95797 103202
0 56447 5 1 1 56446
0 56448 7 1 2 56447 102358
0 56449 5 1 1 56448
0 56450 7 1 2 73517 56449
0 56451 5 1 1 56450
0 56452 7 1 2 77955 87771
0 56453 5 1 1 56452
0 56454 7 1 2 89503 98252
0 56455 5 1 1 56454
0 56456 7 1 2 73528 56455
0 56457 5 1 1 56456
0 56458 7 1 2 87814 56457
0 56459 5 1 1 56458
0 56460 7 1 2 56453 56459
0 56461 7 1 2 56451 56460
0 56462 7 1 2 56445 56461
0 56463 5 1 1 56462
0 56464 7 1 2 85986 56463
0 56465 5 1 1 56464
0 56466 7 1 2 72681 98253
0 56467 5 1 1 56466
0 56468 7 1 2 76601 103401
0 56469 5 1 1 56468
0 56470 7 1 2 74737 94042
0 56471 5 1 1 56470
0 56472 7 1 2 56469 56471
0 56473 7 1 2 56467 56472
0 56474 5 1 1 56473
0 56475 7 1 2 70786 56474
0 56476 5 1 1 56475
0 56477 7 1 2 103577 56476
0 56478 5 1 1 56477
0 56479 7 1 2 81236 56478
0 56480 5 1 1 56479
0 56481 7 1 2 103575 56480
0 56482 5 1 1 56481
0 56483 7 1 2 87815 56482
0 56484 5 1 1 56483
0 56485 7 1 2 87759 103557
0 56486 5 1 1 56485
0 56487 7 1 2 88009 97917
0 56488 7 1 2 100898 56487
0 56489 5 1 1 56488
0 56490 7 1 2 56486 56489
0 56491 5 1 1 56490
0 56492 7 1 2 66786 56491
0 56493 5 1 1 56492
0 56494 7 1 2 61922 103389
0 56495 7 1 2 103552 56494
0 56496 5 1 1 56495
0 56497 7 1 2 56493 56496
0 56498 5 1 1 56497
0 56499 7 1 2 73518 56498
0 56500 5 1 1 56499
0 56501 7 1 2 81237 87760
0 56502 7 1 2 103489 56501
0 56503 5 1 1 56502
0 56504 7 1 2 56500 56503
0 56505 7 1 2 56484 56504
0 56506 5 1 1 56505
0 56507 7 1 2 69641 56506
0 56508 5 1 1 56507
0 56509 7 1 2 56465 56508
0 56510 5 1 1 56509
0 56511 7 1 2 65256 56510
0 56512 5 1 1 56511
0 56513 7 1 2 87816 103584
0 56514 5 1 1 56513
0 56515 7 1 2 56512 56514
0 56516 5 1 1 56515
0 56517 7 1 2 98000 103095
0 56518 7 1 2 56516 56517
0 56519 5 1 1 56518
0 56520 7 1 2 56431 56519
0 56521 7 1 2 56327 56520
0 56522 7 1 2 56120 56521
0 56523 7 1 2 55920 56522
0 56524 7 1 2 55559 56523
0 56525 7 1 2 55198 56524
0 56526 5 1 1 56525
0 56527 7 1 2 54350 56526
0 56528 5 1 1 56527
0 56529 7 1 2 90791 94552
0 56530 5 1 1 56529
0 56531 7 1 2 66332 100085
0 56532 5 1 1 56531
0 56533 7 1 2 101742 56532
0 56534 5 1 1 56533
0 56535 7 1 2 71391 56534
0 56536 5 1 1 56535
0 56537 7 1 2 69642 98714
0 56538 7 1 2 100782 56537
0 56539 5 1 1 56538
0 56540 7 1 2 56536 56539
0 56541 5 1 1 56540
0 56542 7 1 2 65878 56541
0 56543 5 1 1 56542
0 56544 7 1 2 85479 82899
0 56545 7 1 2 100220 56544
0 56546 5 1 1 56545
0 56547 7 1 2 56543 56546
0 56548 5 1 1 56547
0 56549 7 1 2 64598 56548
0 56550 5 1 1 56549
0 56551 7 1 2 84416 103403
0 56552 7 1 2 103504 56551
0 56553 5 1 1 56552
0 56554 7 1 2 56550 56553
0 56555 5 1 1 56554
0 56556 7 1 2 69264 56555
0 56557 5 1 1 56556
0 56558 7 1 2 91662 99116
0 56559 5 1 1 56558
0 56560 7 1 2 70787 100578
0 56561 5 1 1 56560
0 56562 7 1 2 56559 56561
0 56563 5 1 1 56562
0 56564 7 1 2 97482 56563
0 56565 5 1 1 56564
0 56566 7 1 2 56557 56565
0 56567 5 1 1 56566
0 56568 7 1 2 100241 56567
0 56569 5 1 1 56568
0 56570 7 1 2 102922 103071
0 56571 7 1 2 97334 56570
0 56572 5 1 1 56571
0 56573 7 1 2 56569 56572
0 56574 5 1 1 56573
0 56575 7 1 2 92655 56574
0 56576 5 1 1 56575
0 56577 7 2 2 84417 93837
0 56578 7 1 2 77017 103618
0 56579 5 1 1 56578
0 56580 7 1 2 102223 97335
0 56581 5 1 1 56580
0 56582 7 1 2 56579 56581
0 56583 5 1 1 56582
0 56584 7 1 2 64599 56583
0 56585 5 1 1 56584
0 56586 7 1 2 89022 90687
0 56587 7 1 2 100917 56586
0 56588 5 1 1 56587
0 56589 7 1 2 56585 56588
0 56590 5 1 1 56589
0 56591 7 1 2 64413 92661
0 56592 7 1 2 56590 56591
0 56593 5 1 1 56592
0 56594 7 1 2 56576 56593
0 56595 5 1 1 56594
0 56596 7 1 2 93952 96955
0 56597 7 1 2 56595 56596
0 56598 5 1 1 56597
0 56599 7 2 2 79142 90849
0 56600 7 1 2 70524 99422
0 56601 7 1 2 103620 56600
0 56602 5 1 1 56601
0 56603 7 2 2 79091 87817
0 56604 7 1 2 85456 99370
0 56605 7 1 2 103622 56604
0 56606 5 1 1 56605
0 56607 7 1 2 56602 56606
0 56608 5 1 1 56607
0 56609 7 1 2 66787 56608
0 56610 5 1 1 56609
0 56611 7 2 2 71270 99371
0 56612 7 2 2 92120 103624
0 56613 7 1 2 88148 98829
0 56614 7 1 2 103626 56613
0 56615 5 1 1 56614
0 56616 7 1 2 56610 56615
0 56617 5 1 1 56616
0 56618 7 1 2 66572 56617
0 56619 5 1 1 56618
0 56620 7 1 2 83317 99910
0 56621 7 1 2 103627 56620
0 56622 5 1 1 56621
0 56623 7 1 2 56619 56622
0 56624 5 1 1 56623
0 56625 7 1 2 101371 56624
0 56626 5 1 1 56625
0 56627 7 2 2 101883 98095
0 56628 7 1 2 89571 92828
0 56629 7 1 2 101258 56628
0 56630 7 1 2 103628 56629
0 56631 5 1 1 56630
0 56632 7 1 2 56626 56631
0 56633 7 1 2 56598 56632
0 56634 5 1 1 56633
0 56635 7 1 2 66060 56634
0 56636 5 1 1 56635
0 56637 7 1 2 71457 95953
0 56638 5 3 1 56637
0 56639 7 1 2 82292 103630
0 56640 7 1 2 92491 56639
0 56641 5 1 1 56640
0 56642 7 2 2 77825 100242
0 56643 7 1 2 62929 103633
0 56644 7 1 2 102640 56643
0 56645 5 1 1 56644
0 56646 7 1 2 56641 56645
0 56647 5 1 1 56646
0 56648 7 1 2 64414 56647
0 56649 5 1 1 56648
0 56650 7 1 2 92841 97348
0 56651 7 1 2 103411 56650
0 56652 7 1 2 103634 56651
0 56653 5 1 1 56652
0 56654 7 1 2 56649 56653
0 56655 5 1 1 56654
0 56656 7 1 2 89272 56655
0 56657 5 1 1 56656
0 56658 7 1 2 75557 92842
0 56659 7 2 2 102245 56658
0 56660 7 1 2 100243 100136
0 56661 7 1 2 103635 56660
0 56662 7 1 2 103496 56661
0 56663 5 1 1 56662
0 56664 7 1 2 56657 56663
0 56665 5 1 1 56664
0 56666 7 1 2 70525 56665
0 56667 5 1 1 56666
0 56668 7 1 2 69265 80329
0 56669 7 1 2 74497 56668
0 56670 7 1 2 100244 100780
0 56671 7 1 2 56669 56670
0 56672 7 1 2 103636 56671
0 56673 5 1 1 56672
0 56674 7 1 2 56667 56673
0 56675 5 1 1 56674
0 56676 7 1 2 62242 56675
0 56677 5 1 1 56676
0 56678 7 1 2 56636 56677
0 56679 5 1 1 56678
0 56680 7 1 2 69075 56679
0 56681 5 1 1 56680
0 56682 7 1 2 71071 84982
0 56683 5 1 1 56682
0 56684 7 1 2 85503 94904
0 56685 5 1 1 56684
0 56686 7 1 2 56683 56685
0 56687 5 1 1 56686
0 56688 7 1 2 65593 56687
0 56689 5 1 1 56688
0 56690 7 1 2 71444 103267
0 56691 5 1 1 56690
0 56692 7 1 2 56689 56691
0 56693 5 1 1 56692
0 56694 7 1 2 64228 56693
0 56695 5 1 1 56694
0 56696 7 1 2 73706 93381
0 56697 5 1 1 56696
0 56698 7 1 2 72481 91079
0 56699 5 1 1 56698
0 56700 7 1 2 71072 56699
0 56701 5 1 1 56700
0 56702 7 1 2 56697 56701
0 56703 7 1 2 56695 56702
0 56704 5 1 1 56703
0 56705 7 1 2 99055 102647
0 56706 7 1 2 56704 56705
0 56707 5 1 1 56706
0 56708 7 3 2 76566 84186
0 56709 7 1 2 92376 103637
0 56710 5 1 1 56709
0 56711 7 2 2 83534 76591
0 56712 7 1 2 97508 103640
0 56713 5 1 1 56712
0 56714 7 1 2 56710 56713
0 56715 5 1 1 56714
0 56716 7 1 2 64229 92492
0 56717 7 1 2 56715 56716
0 56718 5 1 1 56717
0 56719 7 1 2 56707 56718
0 56720 5 1 1 56719
0 56721 7 1 2 64415 56720
0 56722 5 1 1 56721
0 56723 7 1 2 90277 85309
0 56724 5 1 1 56723
0 56725 7 1 2 77993 87327
0 56726 5 1 1 56725
0 56727 7 1 2 56724 56726
0 56728 5 1 1 56727
0 56729 7 1 2 71392 56728
0 56730 5 1 1 56729
0 56731 7 1 2 88376 100927
0 56732 5 1 1 56731
0 56733 7 1 2 56730 56732
0 56734 5 1 1 56733
0 56735 7 1 2 65594 103445
0 56736 7 2 2 56734 56735
0 56737 7 1 2 100317 103642
0 56738 5 1 1 56737
0 56739 7 1 2 90950 103643
0 56740 5 1 1 56739
0 56741 7 1 2 70526 103249
0 56742 5 1 1 56741
0 56743 7 1 2 92412 35903
0 56744 5 1 1 56743
0 56745 7 1 2 64230 56744
0 56746 7 1 2 56742 56745
0 56747 5 1 1 56746
0 56748 7 1 2 35916 56747
0 56749 5 1 1 56748
0 56750 7 1 2 100579 56749
0 56751 5 1 1 56750
0 56752 7 1 2 93296 100099
0 56753 7 1 2 85310 56752
0 56754 5 1 1 56753
0 56755 7 1 2 56751 56754
0 56756 5 1 1 56755
0 56757 7 1 2 69449 56756
0 56758 5 1 1 56757
0 56759 7 1 2 102835 103486
0 56760 5 1 1 56759
0 56761 7 1 2 64416 56760
0 56762 7 1 2 56758 56761
0 56763 5 1 1 56762
0 56764 7 1 2 86384 102661
0 56765 5 1 1 56764
0 56766 7 1 2 74741 100160
0 56767 5 1 1 56766
0 56768 7 1 2 56765 56767
0 56769 5 1 1 56768
0 56770 7 1 2 101515 56769
0 56771 5 1 1 56770
0 56772 7 1 2 102665 100542
0 56773 5 1 1 56772
0 56774 7 1 2 83367 87328
0 56775 5 1 1 56774
0 56776 7 1 2 56773 56775
0 56777 5 1 1 56776
0 56778 7 1 2 73138 56777
0 56779 5 1 1 56778
0 56780 7 1 2 72414 98263
0 56781 5 1 1 56780
0 56782 7 1 2 56781 102970
0 56783 5 1 1 56782
0 56784 7 1 2 83969 56783
0 56785 5 1 1 56784
0 56786 7 1 2 56779 56785
0 56787 7 1 2 56771 56786
0 56788 5 1 1 56787
0 56789 7 1 2 90688 56788
0 56790 5 1 1 56789
0 56791 7 1 2 72902 92871
0 56792 5 1 1 56791
0 56793 7 1 2 94137 56792
0 56794 5 1 1 56793
0 56795 7 1 2 73529 56794
0 56796 5 1 1 56795
0 56797 7 1 2 102872 56796
0 56798 5 1 1 56797
0 56799 7 1 2 69266 56798
0 56800 7 1 2 56790 56799
0 56801 5 1 1 56800
0 56802 7 1 2 67834 56801
0 56803 7 1 2 56763 56802
0 56804 5 1 1 56803
0 56805 7 1 2 56740 56804
0 56806 5 1 1 56805
0 56807 7 1 2 66190 56806
0 56808 5 1 1 56807
0 56809 7 1 2 56738 56808
0 56810 5 1 1 56809
0 56811 7 1 2 100245 56810
0 56812 5 1 1 56811
0 56813 7 1 2 56722 56812
0 56814 5 1 1 56813
0 56815 7 1 2 62243 56814
0 56816 5 1 1 56815
0 56817 7 1 2 61682 84239
0 56818 5 1 1 56817
0 56819 7 1 2 4402 56818
0 56820 5 1 1 56819
0 56821 7 1 2 103553 56820
0 56822 5 1 1 56821
0 56823 7 3 2 93953 100246
0 56824 7 1 2 90278 102995
0 56825 5 1 1 56824
0 56826 7 1 2 83970 96689
0 56827 5 1 1 56826
0 56828 7 1 2 56825 56827
0 56829 5 1 1 56828
0 56830 7 1 2 103644 56829
0 56831 5 1 1 56830
0 56832 7 1 2 56822 56831
0 56833 5 1 1 56832
0 56834 7 1 2 92493 56833
0 56835 5 1 1 56834
0 56836 7 1 2 81153 103386
0 56837 5 1 1 56836
0 56838 7 1 2 103547 56837
0 56839 5 1 1 56838
0 56840 7 1 2 102650 56839
0 56841 5 1 1 56840
0 56842 7 1 2 87689 98626
0 56843 7 1 2 102112 56842
0 56844 7 1 2 86748 56843
0 56845 5 1 1 56844
0 56846 7 1 2 56841 56845
0 56847 5 1 1 56846
0 56848 7 1 2 66788 56847
0 56849 5 1 1 56848
0 56850 7 1 2 80305 97439
0 56851 5 1 1 56850
0 56852 7 1 2 103555 56851
0 56853 5 1 1 56852
0 56854 7 1 2 67753 56853
0 56855 5 1 1 56854
0 56856 7 1 2 77101 96704
0 56857 5 1 1 56856
0 56858 7 1 2 56855 56857
0 56859 5 1 1 56858
0 56860 7 1 2 95920 102703
0 56861 7 1 2 56859 56860
0 56862 5 1 1 56861
0 56863 7 1 2 56849 56862
0 56864 5 1 1 56863
0 56865 7 1 2 93838 56864
0 56866 5 1 1 56865
0 56867 7 1 2 56835 56866
0 56868 5 1 1 56867
0 56869 7 1 2 64417 56868
0 56870 5 1 1 56869
0 56871 7 1 2 87238 101699
0 56872 5 1 1 56871
0 56873 7 1 2 99110 102565
0 56874 5 1 1 56873
0 56875 7 1 2 56872 56874
0 56876 5 1 1 56875
0 56877 7 1 2 67754 56876
0 56878 5 1 1 56877
0 56879 7 1 2 42710 56878
0 56880 5 1 1 56879
0 56881 7 1 2 70788 56880
0 56882 5 1 1 56881
0 56883 7 1 2 95790 100080
0 56884 5 1 1 56883
0 56885 7 1 2 56882 56884
0 56886 5 1 1 56885
0 56887 7 1 2 66333 56886
0 56888 5 1 1 56887
0 56889 7 1 2 101739 102636
0 56890 5 1 1 56889
0 56891 7 1 2 56888 56890
0 56892 5 1 1 56891
0 56893 7 1 2 92656 92820
0 56894 7 1 2 103645 56893
0 56895 7 1 2 56892 56894
0 56896 5 1 1 56895
0 56897 7 1 2 56870 56896
0 56898 5 1 1 56897
0 56899 7 1 2 73519 56898
0 56900 5 1 1 56899
0 56901 7 1 2 91195 87818
0 56902 7 1 2 91498 56901
0 56903 7 1 2 103625 56902
0 56904 5 1 1 56903
0 56905 7 1 2 77756 93515
0 56906 5 1 1 56905
0 56907 7 1 2 33613 56906
0 56908 5 1 1 56907
0 56909 7 1 2 81132 85106
0 56910 7 1 2 56908 56909
0 56911 5 1 1 56910
0 56912 7 1 2 56904 56911
0 56913 5 1 1 56912
0 56914 7 1 2 100191 56913
0 56915 5 1 1 56914
0 56916 7 1 2 85730 78273
0 56917 7 1 2 85457 56916
0 56918 7 1 2 92674 56917
0 56919 5 1 1 56918
0 56920 7 1 2 56915 56919
0 56921 5 1 1 56920
0 56922 7 1 2 65004 56921
0 56923 5 1 1 56922
0 56924 7 1 2 75427 95624
0 56925 5 1 1 56924
0 56926 7 1 2 20830 56925
0 56927 5 1 1 56926
0 56928 7 1 2 71468 92657
0 56929 7 1 2 93839 56928
0 56930 7 1 2 97245 56929
0 56931 7 1 2 56927 56930
0 56932 5 1 1 56931
0 56933 7 1 2 56923 56932
0 56934 5 1 1 56933
0 56935 7 1 2 66573 56934
0 56936 5 1 1 56935
0 56937 7 1 2 96612 101184
0 56938 5 1 1 56937
0 56939 7 1 2 71393 96108
0 56940 7 1 2 103646 56939
0 56941 5 1 1 56940
0 56942 7 1 2 56938 56941
0 56943 5 1 1 56942
0 56944 7 1 2 93840 56943
0 56945 5 1 1 56944
0 56946 7 1 2 75712 98071
0 56947 7 1 2 97491 56946
0 56948 7 1 2 100820 56947
0 56949 5 1 1 56948
0 56950 7 1 2 56945 56949
0 56951 5 1 1 56950
0 56952 7 1 2 87177 92658
0 56953 7 1 2 56951 56952
0 56954 5 1 1 56953
0 56955 7 1 2 56936 56954
0 56956 5 1 1 56955
0 56957 7 1 2 72213 56956
0 56958 5 1 1 56957
0 56959 7 1 2 69149 56958
0 56960 7 1 2 56900 56959
0 56961 7 1 2 56816 56960
0 56962 7 1 2 56681 56961
0 56963 5 1 1 56962
0 56964 7 1 2 77706 103008
0 56965 5 1 1 56964
0 56966 7 1 2 75616 56965
0 56967 5 1 1 56966
0 56968 7 1 2 70527 56967
0 56969 5 1 1 56968
0 56970 7 1 2 62244 76793
0 56971 5 1 1 56970
0 56972 7 1 2 56969 56971
0 56973 5 1 1 56972
0 56974 7 1 2 70789 56973
0 56975 5 1 1 56974
0 56976 7 1 2 65879 77632
0 56977 5 1 1 56976
0 56978 7 1 2 6198 56977
0 56979 5 1 1 56978
0 56980 7 1 2 77707 56979
0 56981 5 1 1 56980
0 56982 7 1 2 56975 56981
0 56983 5 1 1 56982
0 56984 7 1 2 70979 56983
0 56985 5 1 1 56984
0 56986 7 1 2 71096 325
0 56987 5 3 1 56986
0 56988 7 1 2 73589 85160
0 56989 7 1 2 103647 56988
0 56990 5 1 1 56989
0 56991 7 1 2 56985 56990
0 56992 5 1 1 56991
0 56993 7 1 2 64231 56992
0 56994 5 1 1 56993
0 56995 7 1 2 71073 103264
0 56996 5 1 1 56995
0 56997 7 1 2 89829 86200
0 56998 5 1 1 56997
0 56999 7 1 2 56996 56998
0 57000 5 1 1 56999
0 57001 7 1 2 69076 57000
0 57002 5 1 1 57001
0 57003 7 1 2 72214 100247
0 57004 5 1 1 57003
0 57005 7 1 2 95058 57004
0 57006 5 1 1 57005
0 57007 7 1 2 62245 57006
0 57008 5 1 1 57007
0 57009 7 1 2 57002 57008
0 57010 5 1 1 57009
0 57011 7 1 2 70528 57010
0 57012 5 1 1 57011
0 57013 7 1 2 56994 57012
0 57014 5 1 1 57013
0 57015 7 1 2 90279 57014
0 57016 5 1 1 57015
0 57017 7 1 2 100248 100062
0 57018 7 1 2 96278 57017
0 57019 5 1 1 57018
0 57020 7 1 2 57016 57019
0 57021 5 1 1 57020
0 57022 7 1 2 91035 57021
0 57023 5 1 1 57022
0 57024 7 1 2 87286 75614
0 57025 5 1 1 57024
0 57026 7 1 2 77708 103015
0 57027 5 1 1 57026
0 57028 7 1 2 57025 57027
0 57029 5 1 1 57028
0 57030 7 1 2 72682 57029
0 57031 5 1 1 57030
0 57032 7 1 2 78353 74166
0 57033 5 1 1 57032
0 57034 7 1 2 908 100295
0 57035 5 1 1 57034
0 57036 7 1 2 103648 57035
0 57037 5 1 1 57036
0 57038 7 1 2 11699 57037
0 57039 5 1 1 57038
0 57040 7 1 2 70529 57039
0 57041 5 1 1 57040
0 57042 7 1 2 57033 57041
0 57043 7 1 2 57031 57042
0 57044 5 1 1 57043
0 57045 7 1 2 103315 99293
0 57046 7 1 2 57044 57045
0 57047 5 1 1 57046
0 57048 7 1 2 6623 53506
0 57049 5 1 1 57048
0 57050 7 1 2 70530 57049
0 57051 5 1 1 57050
0 57052 7 1 2 70790 102092
0 57053 5 1 1 57052
0 57054 7 1 2 57051 57053
0 57055 5 1 1 57054
0 57056 7 2 2 69450 102941
0 57057 7 1 2 93887 103650
0 57058 7 1 2 57055 57057
0 57059 5 1 1 57058
0 57060 7 1 2 57047 57059
0 57061 7 1 2 57023 57060
0 57062 5 1 1 57061
0 57063 7 1 2 69267 57062
0 57064 5 1 1 57063
0 57065 7 1 2 79629 94138
0 57066 5 1 1 57065
0 57067 7 1 2 102976 57066
0 57068 5 1 1 57067
0 57069 7 1 2 103651 57068
0 57070 5 1 1 57069
0 57071 7 1 2 62930 103638
0 57072 5 1 1 57071
0 57073 7 1 2 71074 87329
0 57074 5 1 1 57073
0 57075 7 1 2 57072 57074
0 57076 5 1 1 57075
0 57077 7 1 2 79630 57076
0 57078 5 1 1 57077
0 57079 7 1 2 74167 87330
0 57080 5 1 1 57079
0 57081 7 1 2 57078 57080
0 57082 5 1 1 57081
0 57083 7 1 2 72683 57082
0 57084 5 1 1 57083
0 57085 7 1 2 71075 90280
0 57086 5 1 1 57085
0 57087 7 1 2 71445 87331
0 57088 5 1 1 57087
0 57089 7 1 2 57086 57088
0 57090 5 1 1 57089
0 57091 7 1 2 84675 103023
0 57092 5 1 1 57091
0 57093 7 1 2 73857 96345
0 57094 5 1 1 57093
0 57095 7 1 2 57092 57094
0 57096 5 1 1 57095
0 57097 7 1 2 57090 57096
0 57098 5 1 1 57097
0 57099 7 1 2 103639 102978
0 57100 5 1 1 57099
0 57101 7 1 2 71748 103641
0 57102 7 1 2 103057 57101
0 57103 5 1 1 57102
0 57104 7 1 2 57100 57103
0 57105 7 1 2 57098 57104
0 57106 7 1 2 57084 57105
0 57107 5 1 1 57106
0 57108 7 1 2 90629 57107
0 57109 5 1 1 57108
0 57110 7 1 2 57070 57109
0 57111 5 1 1 57110
0 57112 7 1 2 99769 57111
0 57113 5 1 1 57112
0 57114 7 1 2 64303 57113
0 57115 7 1 2 57064 57114
0 57116 5 1 1 57115
0 57117 7 1 2 65257 57116
0 57118 7 1 2 56963 57117
0 57119 5 1 1 57118
0 57120 7 1 2 88889 98687
0 57121 5 1 1 57120
0 57122 7 3 2 92843 97566
0 57123 7 1 2 75558 78800
0 57124 7 1 2 103652 57123
0 57125 5 1 1 57124
0 57126 7 1 2 57121 57125
0 57127 5 1 1 57126
0 57128 7 1 2 69451 57127
0 57129 5 1 1 57128
0 57130 7 1 2 64304 88737
0 57131 7 1 2 84281 57130
0 57132 7 1 2 99294 57131
0 57133 5 1 1 57132
0 57134 7 1 2 57129 57133
0 57135 5 1 1 57134
0 57136 7 1 2 70531 57135
0 57137 5 1 1 57136
0 57138 7 1 2 72767 100515
0 57139 7 1 2 101372 57138
0 57140 5 1 1 57139
0 57141 7 1 2 57137 57140
0 57142 5 1 1 57141
0 57143 7 1 2 84418 57142
0 57144 5 1 1 57143
0 57145 7 1 2 89033 94638
0 57146 7 1 2 99056 57145
0 57147 5 1 1 57146
0 57148 7 1 2 88738 97567
0 57149 7 1 2 100747 57148
0 57150 5 1 1 57149
0 57151 7 1 2 57147 57150
0 57152 5 1 1 57151
0 57153 7 1 2 101167 57152
0 57154 5 1 1 57153
0 57155 7 1 2 69077 57154
0 57156 7 1 2 57144 57155
0 57157 5 1 1 57156
0 57158 7 1 2 94639 101654
0 57159 7 2 2 99848 57158
0 57160 7 1 2 62989 103655
0 57161 5 1 1 57160
0 57162 7 1 2 64600 99132
0 57163 5 1 1 57162
0 57164 7 1 2 57161 57163
0 57165 5 1 1 57164
0 57166 7 1 2 62688 57165
0 57167 5 1 1 57166
0 57168 7 3 2 99196 97590
0 57169 7 1 2 95279 97577
0 57170 7 1 2 103657 57169
0 57171 5 1 1 57170
0 57172 7 1 2 57167 57171
0 57173 5 1 1 57172
0 57174 7 1 2 66191 57173
0 57175 5 1 1 57174
0 57176 7 1 2 103656 102525
0 57177 5 1 1 57176
0 57178 7 1 2 57175 57177
0 57179 5 1 1 57178
0 57180 7 1 2 89273 57179
0 57181 5 1 1 57180
0 57182 7 1 2 90281 72862
0 57183 7 1 2 100540 57182
0 57184 7 1 2 103653 57183
0 57185 5 1 1 57184
0 57186 7 1 2 64232 57185
0 57187 7 1 2 57181 57186
0 57188 5 1 1 57187
0 57189 7 1 2 57157 57188
0 57190 5 1 1 57189
0 57191 7 2 2 92844 99111
0 57192 7 2 2 95429 103660
0 57193 7 1 2 77936 90883
0 57194 7 1 2 79548 57193
0 57195 7 1 2 103662 57194
0 57196 5 1 1 57195
0 57197 7 1 2 57190 57196
0 57198 5 1 1 57197
0 57199 7 1 2 68882 57198
0 57200 5 1 1 57199
0 57201 7 2 2 82706 101267
0 57202 7 1 2 94244 103600
0 57203 5 1 1 57202
0 57204 7 1 2 62931 57203
0 57205 5 1 1 57204
0 57206 7 1 2 67545 102878
0 57207 5 1 1 57206
0 57208 7 1 2 57205 57207
0 57209 5 1 1 57208
0 57210 7 1 2 103664 57209
0 57211 5 1 1 57210
0 57212 7 1 2 90781 99229
0 57213 7 1 2 94031 57212
0 57214 5 1 1 57213
0 57215 7 1 2 70532 101611
0 57216 7 1 2 103665 57215
0 57217 5 1 1 57216
0 57218 7 1 2 57214 57217
0 57219 5 1 1 57218
0 57220 7 1 2 67755 57219
0 57221 5 1 1 57220
0 57222 7 1 2 57211 57221
0 57223 5 1 1 57222
0 57224 7 1 2 66334 57223
0 57225 5 1 1 57224
0 57226 7 1 2 62689 101702
0 57227 5 1 1 57226
0 57228 7 1 2 94032 101670
0 57229 5 1 1 57228
0 57230 7 1 2 57227 57229
0 57231 5 1 1 57230
0 57232 7 1 2 74929 98738
0 57233 7 1 2 57231 57232
0 57234 5 1 1 57233
0 57235 7 1 2 57225 57234
0 57236 5 1 1 57235
0 57237 7 1 2 69452 57236
0 57238 5 1 1 57237
0 57239 7 1 2 87332 98081
0 57240 7 1 2 101553 57239
0 57241 5 1 1 57240
0 57242 7 1 2 57238 57241
0 57243 5 1 1 57242
0 57244 7 1 2 64013 57243
0 57245 5 1 1 57244
0 57246 7 1 2 97655 99703
0 57247 5 1 1 57246
0 57248 7 1 2 69150 87518
0 57249 7 1 2 102392 57248
0 57250 5 1 1 57249
0 57251 7 1 2 57247 57250
0 57252 5 1 1 57251
0 57253 7 1 2 66335 57252
0 57254 5 1 1 57253
0 57255 7 1 2 99673 98739
0 57256 5 1 1 57255
0 57257 7 1 2 57254 57256
0 57258 5 1 1 57257
0 57259 7 1 2 89274 72863
0 57260 7 1 2 57258 57259
0 57261 5 1 1 57260
0 57262 7 1 2 57245 57261
0 57263 5 1 1 57262
0 57264 7 1 2 66192 57263
0 57265 5 1 1 57264
0 57266 7 1 2 67835 102787
0 57267 5 1 1 57266
0 57268 7 1 2 64810 102252
0 57269 5 1 1 57268
0 57270 7 1 2 57267 57269
0 57271 5 1 1 57270
0 57272 7 1 2 74503 57271
0 57273 5 1 1 57272
0 57274 7 1 2 79243 91382
0 57275 7 1 2 100569 57274
0 57276 5 1 1 57275
0 57277 7 1 2 57273 57276
0 57278 5 1 1 57277
0 57279 7 1 2 65595 72252
0 57280 7 1 2 57278 57279
0 57281 5 1 1 57280
0 57282 7 1 2 81798 91383
0 57283 7 1 2 101984 57282
0 57284 5 1 1 57283
0 57285 7 1 2 57281 57284
0 57286 5 1 1 57285
0 57287 7 1 2 69453 97730
0 57288 7 1 2 57286 57287
0 57289 5 1 1 57288
0 57290 7 1 2 57265 57289
0 57291 7 1 2 57200 57290
0 57292 5 1 1 57291
0 57293 7 1 2 65880 57292
0 57294 5 1 1 57293
0 57295 7 2 2 65596 98688
0 57296 5 1 1 103666
0 57297 7 1 2 66193 99133
0 57298 5 1 1 57297
0 57299 7 1 2 57296 57298
0 57300 5 1 1 57299
0 57301 7 1 2 85849 57300
0 57302 5 1 1 57301
0 57303 7 2 2 100290 102308
0 57304 7 1 2 84024 92845
0 57305 7 1 2 97591 57304
0 57306 7 1 2 103668 57305
0 57307 5 1 1 57306
0 57308 7 1 2 57302 57307
0 57309 5 1 1 57308
0 57310 7 1 2 90282 57309
0 57311 5 1 1 57310
0 57312 7 1 2 69078 99372
0 57313 7 1 2 84051 57312
0 57314 7 1 2 103663 57313
0 57315 5 1 1 57314
0 57316 7 1 2 57311 57315
0 57317 5 1 1 57316
0 57318 7 1 2 103009 57317
0 57319 5 1 1 57318
0 57320 7 1 2 69454 94739
0 57321 7 1 2 96742 57320
0 57322 7 1 2 93888 57321
0 57323 5 1 1 57322
0 57324 7 1 2 87411 102192
0 57325 7 1 2 97639 57324
0 57326 7 1 2 91663 57325
0 57327 5 1 1 57326
0 57328 7 1 2 57323 57327
0 57329 5 1 1 57328
0 57330 7 1 2 64233 57329
0 57331 5 1 1 57330
0 57332 7 1 2 102648 103545
0 57333 5 1 1 57332
0 57334 7 1 2 57331 57333
0 57335 5 1 1 57334
0 57336 7 1 2 93841 57335
0 57337 5 1 1 57336
0 57338 7 1 2 64014 103164
0 57339 5 1 1 57338
0 57340 7 1 2 61683 100928
0 57341 5 1 1 57340
0 57342 7 1 2 57339 57341
0 57343 5 1 1 57342
0 57344 7 1 2 62690 57343
0 57345 5 1 1 57344
0 57346 7 1 2 72810 96743
0 57347 7 1 2 85666 57346
0 57348 5 1 1 57347
0 57349 7 1 2 57345 57348
0 57350 5 1 1 57349
0 57351 7 1 2 103654 57350
0 57352 5 1 1 57351
0 57353 7 1 2 57337 57352
0 57354 5 1 1 57353
0 57355 7 1 2 65597 57354
0 57356 5 1 1 57355
0 57357 7 1 2 83789 97592
0 57358 7 1 2 95652 103661
0 57359 7 1 2 57357 57358
0 57360 5 1 1 57359
0 57361 7 1 2 57356 57360
0 57362 5 1 1 57361
0 57363 7 1 2 67081 57362
0 57364 5 1 1 57363
0 57365 7 1 2 57319 57364
0 57366 5 1 1 57365
0 57367 7 1 2 70791 57366
0 57368 5 1 1 57367
0 57369 7 1 2 94139 103619
0 57370 5 1 1 57369
0 57371 7 1 2 80248 100291
0 57372 7 1 2 102846 57371
0 57373 5 1 1 57372
0 57374 7 1 2 57370 57373
0 57375 5 1 1 57374
0 57376 7 1 2 93740 95183
0 57377 7 1 2 103519 57376
0 57378 7 1 2 57375 57377
0 57379 5 1 1 57378
0 57380 7 1 2 69268 57379
0 57381 7 1 2 57368 57380
0 57382 7 1 2 57294 57381
0 57383 5 1 1 57382
0 57384 7 2 2 96979 100100
0 57385 5 1 1 103670
0 57386 7 1 2 61684 95543
0 57387 7 1 2 102704 57386
0 57388 7 1 2 99849 57387
0 57389 5 1 1 57388
0 57390 7 1 2 57385 57389
0 57391 5 1 1 57390
0 57392 7 1 2 78354 57391
0 57393 5 1 1 57392
0 57394 7 1 2 73092 95413
0 57395 5 1 1 57394
0 57396 7 1 2 101018 57395
0 57397 5 1 1 57396
0 57398 7 1 2 97326 57397
0 57399 5 1 1 57398
0 57400 7 1 2 100504 57399
0 57401 5 1 1 57400
0 57402 7 1 2 100580 57401
0 57403 5 1 1 57402
0 57404 7 1 2 57393 57403
0 57405 5 1 1 57404
0 57406 7 1 2 69455 57405
0 57407 5 1 1 57406
0 57408 7 1 2 98663 52510
0 57409 5 1 1 57408
0 57410 7 1 2 100889 57409
0 57411 5 1 1 57410
0 57412 7 1 2 57407 57411
0 57413 5 1 1 57412
0 57414 7 1 2 67082 57413
0 57415 5 1 1 57414
0 57416 7 2 2 84908 36219
0 57417 5 1 1 103672
0 57418 7 1 2 102219 100065
0 57419 7 1 2 57417 57418
0 57420 5 1 1 57419
0 57421 7 1 2 64418 57420
0 57422 7 1 2 57415 57421
0 57423 5 1 1 57422
0 57424 7 1 2 100249 57423
0 57425 7 1 2 57383 57424
0 57426 5 1 1 57425
0 57427 7 1 2 103399 103573
0 57428 5 1 1 57427
0 57429 7 1 2 65881 57428
0 57430 5 1 1 57429
0 57431 7 1 2 94421 95873
0 57432 5 1 1 57431
0 57433 7 1 2 70792 86233
0 57434 7 1 2 57432 57433
0 57435 5 1 1 57434
0 57436 7 1 2 57430 57435
0 57437 5 1 1 57436
0 57438 7 1 2 65598 57437
0 57439 5 1 1 57438
0 57440 7 1 2 103318 57439
0 57441 5 1 1 57440
0 57442 7 1 2 71076 57441
0 57443 5 1 1 57442
0 57444 7 1 2 65599 103391
0 57445 5 1 1 57444
0 57446 7 1 2 67083 103292
0 57447 5 1 1 57446
0 57448 7 1 2 72741 57447
0 57449 7 1 2 57445 57448
0 57450 5 1 1 57449
0 57451 7 1 2 71446 57450
0 57452 5 1 1 57451
0 57453 7 1 2 57443 57452
0 57454 5 1 1 57453
0 57455 7 1 2 99746 97520
0 57456 7 1 2 57454 57455
0 57457 5 1 1 57456
0 57458 7 1 2 75559 101508
0 57459 5 1 1 57458
0 57460 7 1 2 65600 57459
0 57461 7 1 2 103073 57460
0 57462 5 1 1 57461
0 57463 7 1 2 40586 57462
0 57464 5 1 1 57463
0 57465 7 1 2 67546 57464
0 57466 5 1 1 57465
0 57467 7 1 2 66061 77971
0 57468 7 1 2 89743 57467
0 57469 5 1 1 57468
0 57470 7 1 2 57466 57469
0 57471 5 1 1 57470
0 57472 7 1 2 71077 57471
0 57473 5 1 1 57472
0 57474 7 1 2 82637 96812
0 57475 5 1 1 57474
0 57476 7 1 2 57473 57475
0 57477 5 1 1 57476
0 57478 7 1 2 69079 57477
0 57479 5 1 1 57478
0 57480 7 1 2 101866 103468
0 57481 5 1 1 57480
0 57482 7 1 2 77691 101965
0 57483 5 1 1 57482
0 57484 7 1 2 57481 57483
0 57485 5 1 1 57484
0 57486 7 1 2 62932 57485
0 57487 5 1 1 57486
0 57488 7 1 2 73784 76854
0 57489 7 1 2 85922 57488
0 57490 5 1 1 57489
0 57491 7 1 2 57487 57490
0 57492 5 1 1 57491
0 57493 7 1 2 65601 57492
0 57494 5 1 1 57493
0 57495 7 1 2 57479 57494
0 57496 5 1 1 57495
0 57497 7 1 2 69456 99057
0 57498 7 1 2 57496 57497
0 57499 5 1 1 57498
0 57500 7 1 2 57457 57499
0 57501 5 1 1 57500
0 57502 7 1 2 69269 57501
0 57503 5 1 1 57502
0 57504 7 1 2 71104 103465
0 57505 5 1 1 57504
0 57506 7 1 2 85385 77709
0 57507 5 1 1 57506
0 57508 7 1 2 57505 57507
0 57509 5 1 1 57508
0 57510 7 1 2 66062 57509
0 57511 5 1 1 57510
0 57512 7 1 2 79660 95951
0 57513 5 1 1 57512
0 57514 7 1 2 57511 57513
0 57515 5 1 1 57514
0 57516 7 1 2 65882 57515
0 57517 5 1 1 57516
0 57518 7 1 2 71078 24364
0 57519 5 1 1 57518
0 57520 7 1 2 89884 94140
0 57521 5 1 1 57520
0 57522 7 1 2 57519 57521
0 57523 5 1 1 57522
0 57524 7 1 2 65602 57523
0 57525 5 1 1 57524
0 57526 7 1 2 94110 95954
0 57527 5 1 1 57526
0 57528 7 1 2 67084 103631
0 57529 7 1 2 57527 57528
0 57530 5 1 1 57529
0 57531 7 1 2 57525 57530
0 57532 7 1 2 57517 57531
0 57533 5 1 1 57532
0 57534 7 1 2 100302 57533
0 57535 5 1 1 57534
0 57536 7 1 2 71394 71482
0 57537 5 1 1 57536
0 57538 7 1 2 75634 57537
0 57539 5 1 1 57538
0 57540 7 1 2 72589 57539
0 57541 5 1 1 57540
0 57542 7 1 2 89023 98331
0 57543 5 1 1 57542
0 57544 7 1 2 57541 57543
0 57545 5 2 1 57544
0 57546 7 1 2 65603 103674
0 57547 5 1 1 57546
0 57548 7 1 2 67085 77007
0 57549 5 1 1 57548
0 57550 7 1 2 57547 57549
0 57551 5 1 1 57550
0 57552 7 1 2 102764 57551
0 57553 5 1 1 57552
0 57554 7 1 2 57535 57553
0 57555 5 1 1 57554
0 57556 7 1 2 99770 57555
0 57557 5 1 1 57556
0 57558 7 1 2 57503 57557
0 57559 5 1 1 57558
0 57560 7 1 2 64305 57559
0 57561 5 1 1 57560
0 57562 7 1 2 77505 71461
0 57563 5 1 1 57562
0 57564 7 1 2 102826 97430
0 57565 5 1 1 57564
0 57566 7 1 2 57563 57565
0 57567 5 1 1 57566
0 57568 7 1 2 65883 57567
0 57569 5 1 1 57568
0 57570 7 1 2 89882 95948
0 57571 5 1 1 57570
0 57572 7 1 2 84107 78382
0 57573 5 1 1 57572
0 57574 7 1 2 57571 57573
0 57575 7 1 2 57569 57574
0 57576 5 1 1 57575
0 57577 7 1 2 103432 57576
0 57578 5 1 1 57577
0 57579 7 1 2 72684 10532
0 57580 7 1 2 100250 57579
0 57581 7 1 2 103436 57580
0 57582 5 1 1 57581
0 57583 7 1 2 57578 57582
0 57584 5 1 1 57583
0 57585 7 1 2 66194 57584
0 57586 5 1 1 57585
0 57587 7 1 2 92220 97599
0 57588 7 1 2 103675 57587
0 57589 5 1 1 57588
0 57590 7 1 2 57586 57589
0 57591 5 1 1 57590
0 57592 7 1 2 70533 57591
0 57593 5 1 1 57592
0 57594 7 1 2 72811 90689
0 57595 7 1 2 99038 57594
0 57596 7 1 2 86115 98705
0 57597 7 1 2 57595 57596
0 57598 5 1 1 57597
0 57599 7 1 2 57593 57598
0 57600 5 1 1 57599
0 57601 7 1 2 100713 57600
0 57602 5 1 1 57601
0 57603 7 1 2 57561 57602
0 57604 5 1 1 57603
0 57605 7 1 2 89275 57604
0 57606 5 1 1 57605
0 57607 7 1 2 91248 87992
0 57608 5 1 1 57607
0 57609 7 2 2 91384 99969
0 57610 7 1 2 69457 79549
0 57611 7 1 2 103676 57610
0 57612 7 1 2 57608 57611
0 57613 5 1 1 57612
0 57614 7 1 2 102767 103483
0 57615 5 1 1 57614
0 57616 7 1 2 64811 102651
0 57617 7 1 2 57615 57616
0 57618 5 1 1 57617
0 57619 7 1 2 57613 57618
0 57620 5 1 1 57619
0 57621 7 1 2 69151 57620
0 57622 5 1 1 57621
0 57623 7 1 2 103335 99311
0 57624 7 1 2 102637 57623
0 57625 5 1 1 57624
0 57626 7 1 2 57622 57625
0 57627 5 1 1 57626
0 57628 7 1 2 71447 57627
0 57629 5 1 1 57628
0 57630 7 1 2 67756 94932
0 57631 5 1 1 57630
0 57632 7 1 2 76336 80544
0 57633 5 1 1 57632
0 57634 7 1 2 57631 57633
0 57635 5 1 1 57634
0 57636 7 1 2 96980 57635
0 57637 5 1 1 57636
0 57638 7 1 2 84326 78355
0 57639 7 1 2 99334 57638
0 57640 5 1 1 57639
0 57641 7 1 2 57637 57640
0 57642 5 1 1 57641
0 57643 7 1 2 79092 95921
0 57644 7 1 2 57642 57643
0 57645 5 1 1 57644
0 57646 7 1 2 57629 57645
0 57647 5 1 1 57646
0 57648 7 1 2 64419 57647
0 57649 5 1 1 57648
0 57650 7 1 2 71079 102638
0 57651 5 1 1 57650
0 57652 7 1 2 77692 100899
0 57653 5 1 1 57652
0 57654 7 1 2 57651 57653
0 57655 5 1 1 57654
0 57656 7 1 2 96167 101035
0 57657 7 1 2 57655 57656
0 57658 5 1 1 57657
0 57659 7 1 2 57649 57658
0 57660 5 1 1 57659
0 57661 7 1 2 93842 57660
0 57662 5 1 1 57661
0 57663 7 1 2 91509 92494
0 57664 5 1 1 57663
0 57665 7 1 2 91385 83310
0 57666 7 1 2 98772 57665
0 57667 5 1 1 57666
0 57668 7 1 2 57664 57667
0 57669 5 1 1 57668
0 57670 7 1 2 100448 57669
0 57671 5 1 1 57670
0 57672 7 1 2 101092 103677
0 57673 7 1 2 100777 57672
0 57674 5 1 1 57673
0 57675 7 1 2 57671 57674
0 57676 5 1 1 57675
0 57677 7 1 2 97426 57676
0 57678 5 1 1 57677
0 57679 7 1 2 102572 103592
0 57680 7 2 2 64234 92821
0 57681 7 1 2 101259 103678
0 57682 7 1 2 57679 57681
0 57683 5 1 1 57682
0 57684 7 1 2 57678 57683
0 57685 5 1 1 57684
0 57686 7 1 2 69152 57685
0 57687 5 1 1 57686
0 57688 7 2 2 93142 103671
0 57689 7 1 2 103680 101215
0 57690 5 1 1 57689
0 57691 7 1 2 57687 57690
0 57692 5 1 1 57691
0 57693 7 1 2 100251 57692
0 57694 5 1 1 57693
0 57695 7 1 2 99880 101400
0 57696 5 1 1 57695
0 57697 7 1 2 76330 95450
0 57698 7 1 2 91349 57697
0 57699 5 1 1 57698
0 57700 7 1 2 57696 57699
0 57701 5 1 1 57700
0 57702 7 1 2 61329 57701
0 57703 5 1 1 57702
0 57704 7 1 2 90125 97882
0 57705 5 1 1 57704
0 57706 7 1 2 57703 57705
0 57707 5 1 1 57706
0 57708 7 1 2 71483 57707
0 57709 5 1 1 57708
0 57710 7 3 2 92495 102309
0 57711 7 1 2 95955 102988
0 57712 5 1 1 57711
0 57713 7 1 2 103632 57712
0 57714 7 1 2 103682 57713
0 57715 5 1 1 57714
0 57716 7 1 2 57709 57715
0 57717 5 1 1 57716
0 57718 7 1 2 83971 57717
0 57719 5 1 1 57718
0 57720 7 1 2 89230 73955
0 57721 5 1 1 57720
0 57722 7 1 2 66063 71080
0 57723 5 1 1 57722
0 57724 7 1 2 57721 57723
0 57725 5 1 1 57724
0 57726 7 1 2 64235 57725
0 57727 5 1 1 57726
0 57728 7 1 2 66064 77699
0 57729 5 1 1 57728
0 57730 7 1 2 77695 95956
0 57731 5 1 1 57730
0 57732 7 1 2 69080 57731
0 57733 5 1 1 57732
0 57734 7 1 2 57729 57733
0 57735 7 1 2 57727 57734
0 57736 5 1 1 57735
0 57737 7 1 2 90316 103683
0 57738 7 1 2 57736 57737
0 57739 5 1 1 57738
0 57740 7 1 2 57719 57739
0 57741 5 1 1 57740
0 57742 7 1 2 70534 57741
0 57743 5 1 1 57742
0 57744 7 1 2 20740 102990
0 57745 5 1 1 57744
0 57746 7 1 2 65604 96690
0 57747 7 1 2 100252 57746
0 57748 7 1 2 103179 57747
0 57749 7 1 2 57745 57748
0 57750 5 1 1 57749
0 57751 7 1 2 57743 57750
0 57752 5 1 1 57751
0 57753 7 1 2 64420 57752
0 57754 5 1 1 57753
0 57755 7 1 2 98332 103667
0 57756 5 1 1 57755
0 57757 7 1 2 70980 97794
0 57758 7 1 2 102891 57757
0 57759 7 1 2 102168 57758
0 57760 5 1 1 57759
0 57761 7 1 2 57756 57760
0 57762 5 1 1 57761
0 57763 7 1 2 87897 92822
0 57764 7 1 2 91523 57763
0 57765 7 1 2 57762 57764
0 57766 5 1 1 57765
0 57767 7 1 2 57754 57766
0 57768 7 1 2 57694 57767
0 57769 7 1 2 57662 57768
0 57770 5 1 1 57769
0 57771 7 1 2 73520 57770
0 57772 5 1 1 57771
0 57773 7 1 2 103609 98896
0 57774 5 1 1 57773
0 57775 7 1 2 80560 97749
0 57776 5 1 1 57775
0 57777 7 1 2 57774 57776
0 57778 5 1 1 57777
0 57779 7 1 2 71448 57778
0 57780 5 1 1 57779
0 57781 7 1 2 89735 97750
0 57782 5 1 1 57781
0 57783 7 1 2 95175 98897
0 57784 7 1 2 102797 57783
0 57785 5 1 1 57784
0 57786 7 1 2 57782 57785
0 57787 5 1 1 57786
0 57788 7 1 2 71081 86440
0 57789 7 1 2 57787 57788
0 57790 5 1 1 57789
0 57791 7 1 2 57780 57790
0 57792 5 1 1 57791
0 57793 7 1 2 67086 57792
0 57794 5 1 1 57793
0 57795 7 1 2 69081 95957
0 57796 5 1 1 57795
0 57797 7 1 2 72215 103649
0 57798 7 2 2 57796 57797
0 57799 5 1 1 103685
0 57800 7 1 2 71182 89231
0 57801 5 1 1 57800
0 57802 7 1 2 57799 57801
0 57803 5 1 1 57802
0 57804 7 1 2 103497 57803
0 57805 5 1 1 57804
0 57806 7 1 2 85920 85360
0 57807 7 1 2 88017 57806
0 57808 5 1 1 57807
0 57809 7 1 2 57805 57808
0 57810 5 1 1 57809
0 57811 7 1 2 103360 57810
0 57812 5 1 1 57811
0 57813 7 1 2 57794 57812
0 57814 5 1 1 57813
0 57815 7 1 2 90283 57814
0 57816 5 1 1 57815
0 57817 7 1 2 68883 102589
0 57818 5 1 1 57817
0 57819 7 1 2 1032 57818
0 57820 5 1 1 57819
0 57821 7 1 2 97751 57820
0 57822 5 1 1 57821
0 57823 7 1 2 64015 103607
0 57824 5 1 1 57823
0 57825 7 1 2 57822 57824
0 57826 5 1 1 57825
0 57827 7 1 2 71484 57826
0 57828 5 1 1 57827
0 57829 7 2 2 99039 102481
0 57830 7 1 2 86501 100485
0 57831 7 1 2 103687 57830
0 57832 5 1 1 57831
0 57833 7 1 2 57828 57832
0 57834 5 1 1 57833
0 57835 7 1 2 66065 57834
0 57836 5 1 1 57835
0 57837 7 1 2 96726 99298
0 57838 5 1 1 57837
0 57839 7 1 2 56174 57838
0 57840 5 1 1 57839
0 57841 7 1 2 70981 89027
0 57842 5 1 1 57841
0 57843 7 1 2 88892 71082
0 57844 5 1 1 57843
0 57845 7 1 2 78640 57844
0 57846 5 1 1 57845
0 57847 7 1 2 57842 57846
0 57848 7 1 2 57840 57847
0 57849 5 1 1 57848
0 57850 7 2 2 76794 97617
0 57851 7 1 2 75560 103689
0 57852 7 1 2 103498 57851
0 57853 5 1 1 57852
0 57854 7 1 2 57849 57853
0 57855 7 1 2 57836 57854
0 57856 5 1 1 57855
0 57857 7 1 2 69082 57856
0 57858 5 1 1 57857
0 57859 7 1 2 91080 103099
0 57860 5 1 1 57859
0 57861 7 1 2 100037 57860
0 57862 5 1 1 57861
0 57863 7 1 2 65884 85739
0 57864 7 1 2 103561 57863
0 57865 5 1 1 57864
0 57866 7 1 2 103470 57865
0 57867 5 1 1 57866
0 57868 7 1 2 103361 57867
0 57869 5 1 1 57868
0 57870 7 1 2 57862 57869
0 57871 5 1 1 57870
0 57872 7 1 2 71083 57871
0 57873 5 1 1 57872
0 57874 7 1 2 73590 103491
0 57875 5 1 1 57874
0 57876 7 1 2 73559 101477
0 57877 5 1 1 57876
0 57878 7 1 2 103690 57877
0 57879 7 1 2 57875 57878
0 57880 5 1 1 57879
0 57881 7 1 2 57873 57880
0 57882 5 1 1 57881
0 57883 7 1 2 64236 57882
0 57884 5 1 1 57883
0 57885 7 1 2 72864 71485
0 57886 5 1 1 57885
0 57887 7 2 2 71084 84025
0 57888 7 1 2 103499 103691
0 57889 5 1 1 57888
0 57890 7 1 2 57886 57889
0 57891 5 1 1 57890
0 57892 7 1 2 97752 57891
0 57893 5 1 1 57892
0 57894 7 1 2 57884 57893
0 57895 7 1 2 57858 57894
0 57896 5 1 1 57895
0 57897 7 1 2 83972 57896
0 57898 5 1 1 57897
0 57899 7 1 2 57816 57898
0 57900 5 1 1 57899
0 57901 7 1 2 90728 57900
0 57902 5 1 1 57901
0 57903 7 1 2 93756 97242
0 57904 5 1 1 57903
0 57905 7 1 2 82999 100112
0 57906 7 1 2 103066 57905
0 57907 5 1 1 57906
0 57908 7 1 2 57904 57907
0 57909 5 1 1 57908
0 57910 7 1 2 100516 57909
0 57911 5 1 1 57910
0 57912 7 1 2 101155 103377
0 57913 5 1 1 57912
0 57914 7 1 2 57913 41336
0 57915 5 1 1 57914
0 57916 7 1 2 102198 57915
0 57917 5 1 1 57916
0 57918 7 2 2 100113 101078
0 57919 7 1 2 102213 101012
0 57920 7 1 2 103693 57919
0 57921 5 1 1 57920
0 57922 7 1 2 57917 57921
0 57923 7 1 2 57911 57922
0 57924 5 1 1 57923
0 57925 7 1 2 71271 57924
0 57926 5 1 1 57925
0 57927 7 1 2 93297 103681
0 57928 5 1 1 57927
0 57929 7 1 2 57926 57928
0 57930 5 1 1 57929
0 57931 7 1 2 65885 57930
0 57932 5 1 1 57931
0 57933 7 1 2 82707 95566
0 57934 7 1 2 101254 57933
0 57935 5 1 1 57934
0 57936 7 1 2 57932 57935
0 57937 5 1 1 57936
0 57938 7 1 2 100253 57937
0 57939 5 1 1 57938
0 57940 7 1 2 95383 102166
0 57941 5 1 1 57940
0 57942 7 1 2 96581 102155
0 57943 5 1 1 57942
0 57944 7 1 2 57941 57943
0 57945 5 1 1 57944
0 57946 7 1 2 93889 57945
0 57947 5 1 1 57946
0 57948 7 1 2 71395 93440
0 57949 7 1 2 97327 57948
0 57950 7 1 2 97243 57949
0 57951 5 1 1 57950
0 57952 7 1 2 57947 57951
0 57953 5 1 1 57952
0 57954 7 1 2 67087 57953
0 57955 5 1 1 57954
0 57956 7 1 2 97142 97731
0 57957 7 3 2 82816 82397
0 57958 7 1 2 97533 103695
0 57959 7 1 2 57956 57958
0 57960 5 1 1 57959
0 57961 7 1 2 57955 57960
0 57962 5 1 1 57961
0 57963 7 1 2 93843 57962
0 57964 5 1 1 57963
0 57965 7 1 2 99230 99475
0 57966 5 1 1 57965
0 57967 7 1 2 71396 84419
0 57968 7 1 2 92966 57967
0 57969 7 1 2 100207 98513
0 57970 7 1 2 57968 57969
0 57971 5 1 1 57970
0 57972 7 1 2 57966 57971
0 57973 5 1 1 57972
0 57974 7 1 2 101872 57973
0 57975 5 1 1 57974
0 57976 7 3 2 68884 82176
0 57977 7 1 2 91643 99212
0 57978 7 1 2 103698 57977
0 57979 7 1 2 103694 57978
0 57980 5 1 1 57979
0 57981 7 1 2 57975 57980
0 57982 7 1 2 57964 57981
0 57983 5 1 1 57982
0 57984 7 1 2 70535 57983
0 57985 5 1 1 57984
0 57986 7 1 2 101273 99817
0 57987 7 1 2 77758 57986
0 57988 5 1 1 57987
0 57989 7 1 2 82454 103699
0 57990 5 1 1 57989
0 57991 7 1 2 43578 57990
0 57992 5 1 1 57991
0 57993 7 1 2 87333 97618
0 57994 7 1 2 57992 57993
0 57995 5 1 1 57994
0 57996 7 1 2 57988 57995
0 57997 5 1 1 57996
0 57998 7 1 2 70536 57997
0 57999 5 1 1 57998
0 58000 7 1 2 64812 76567
0 58001 7 1 2 88149 58000
0 58002 7 1 2 102321 103613
0 58003 7 1 2 58001 58002
0 58004 5 1 1 58003
0 58005 7 1 2 57999 58004
0 58006 5 1 1 58005
0 58007 7 1 2 90729 58006
0 58008 5 1 1 58007
0 58009 7 1 2 97233 98052
0 58010 7 1 2 101860 101070
0 58011 7 1 2 58009 58010
0 58012 5 1 1 58011
0 58013 7 1 2 78520 96551
0 58014 5 1 1 58013
0 58015 7 1 2 78487 97256
0 58016 5 1 1 58015
0 58017 7 1 2 58014 58016
0 58018 5 1 1 58017
0 58019 7 1 2 102795 101079
0 58020 7 1 2 58018 58019
0 58021 5 1 1 58020
0 58022 7 1 2 58012 58021
0 58023 5 1 1 58022
0 58024 7 1 2 103615 58023
0 58025 5 1 1 58024
0 58026 7 1 2 58008 58025
0 58027 7 1 2 57985 58026
0 58028 7 1 2 57939 58027
0 58029 5 1 1 58028
0 58030 7 1 2 72216 58029
0 58031 5 1 1 58030
0 58032 7 1 2 64237 103500
0 58033 5 1 1 58032
0 58034 7 1 2 75748 100487
0 58035 5 1 1 58034
0 58036 7 1 2 72590 87960
0 58037 7 1 2 58035 58036
0 58038 5 1 1 58037
0 58039 7 1 2 58033 58038
0 58040 5 1 1 58039
0 58041 7 1 2 101036 58040
0 58042 5 1 1 58041
0 58043 7 1 2 72865 96981
0 58044 5 1 1 58043
0 58045 7 1 2 58042 58044
0 58046 5 1 1 58045
0 58047 7 1 2 71449 58046
0 58048 5 1 1 58047
0 58049 7 1 2 81225 93305
0 58050 5 1 1 58049
0 58051 7 1 2 101037 58050
0 58052 5 1 1 58051
0 58053 7 1 2 76529 101041
0 58054 5 1 1 58053
0 58055 7 1 2 58052 58054
0 58056 5 1 1 58055
0 58057 7 1 2 71085 58056
0 58058 5 1 1 58057
0 58059 7 1 2 72903 97023
0 58060 5 1 1 58059
0 58061 7 1 2 58060 99916
0 58062 5 1 1 58061
0 58063 7 1 2 96982 101219
0 58064 5 1 1 58063
0 58065 7 1 2 58062 58064
0 58066 5 1 1 58065
0 58067 7 1 2 97431 58066
0 58068 5 1 1 58067
0 58069 7 1 2 71547 101578
0 58070 5 1 1 58069
0 58071 7 1 2 103471 58070
0 58072 5 1 1 58071
0 58073 7 1 2 71450 101038
0 58074 7 1 2 58072 58073
0 58075 5 1 1 58074
0 58076 7 1 2 58068 58075
0 58077 5 1 1 58076
0 58078 7 1 2 70982 58077
0 58079 5 1 1 58078
0 58080 7 1 2 58058 58079
0 58081 7 1 2 58048 58080
0 58082 5 1 1 58081
0 58083 7 1 2 69270 58082
0 58084 5 1 1 58083
0 58085 7 1 2 89437 75296
0 58086 5 1 1 58085
0 58087 7 1 2 17910 58086
0 58088 5 1 1 58087
0 58089 7 1 2 70537 58088
0 58090 5 1 1 58089
0 58091 7 1 2 94923 26670
0 58092 5 1 1 58091
0 58093 7 1 2 73093 58092
0 58094 5 1 1 58093
0 58095 7 1 2 58090 58094
0 58096 5 1 1 58095
0 58097 7 1 2 58096 102501
0 58098 5 1 1 58097
0 58099 7 1 2 71451 101749
0 58100 5 1 1 58099
0 58101 7 1 2 4492 58100
0 58102 5 1 1 58101
0 58103 7 1 2 99373 98586
0 58104 5 1 1 58103
0 58105 7 1 2 62990 95167
0 58106 7 1 2 96727 58105
0 58107 5 1 1 58106
0 58108 7 1 2 58104 58107
0 58109 5 1 1 58108
0 58110 7 1 2 61330 58109
0 58111 5 1 1 58110
0 58112 7 1 2 87928 99307
0 58113 5 1 1 58112
0 58114 7 1 2 93619 58113
0 58115 5 1 1 58114
0 58116 7 1 2 99970 97795
0 58117 7 1 2 58115 58116
0 58118 5 1 1 58117
0 58119 7 1 2 58111 58118
0 58120 5 1 1 58119
0 58121 7 1 2 58102 58120
0 58122 5 1 1 58121
0 58123 7 1 2 58098 58122
0 58124 7 1 2 58084 58123
0 58125 5 1 1 58124
0 58126 7 1 2 101952 58125
0 58127 5 1 1 58126
0 58128 7 1 2 76530 103692
0 58129 5 1 1 58128
0 58130 7 1 2 67757 84109
0 58131 5 1 1 58130
0 58132 7 1 2 58129 58131
0 58133 5 1 1 58132
0 58134 7 1 2 71397 58133
0 58135 5 1 1 58134
0 58136 7 1 2 70538 103673
0 58137 5 1 1 58136
0 58138 7 1 2 71398 84924
0 58139 5 1 1 58138
0 58140 7 1 2 65605 100296
0 58141 7 1 2 58139 58140
0 58142 5 1 1 58141
0 58143 7 1 2 71452 58142
0 58144 7 1 2 58137 58143
0 58145 5 1 1 58144
0 58146 7 1 2 58135 58145
0 58147 5 1 1 58146
0 58148 7 1 2 99264 58147
0 58149 5 1 1 58148
0 58150 7 1 2 71453 80561
0 58151 5 1 1 58150
0 58152 7 1 2 71086 103293
0 58153 5 1 1 58152
0 58154 7 1 2 58151 58153
0 58155 5 1 1 58154
0 58156 7 1 2 99156 58155
0 58157 5 1 1 58156
0 58158 7 1 2 58149 58157
0 58159 5 1 1 58158
0 58160 7 1 2 67088 58159
0 58161 5 1 1 58160
0 58162 7 1 2 103501 98709
0 58163 5 1 1 58162
0 58164 7 1 2 89572 99737
0 58165 7 1 2 97568 58164
0 58166 5 1 1 58165
0 58167 7 1 2 58163 58166
0 58168 5 1 1 58167
0 58169 7 1 2 103598 58168
0 58170 5 1 1 58169
0 58171 7 1 2 103512 99232
0 58172 5 1 1 58171
0 58173 7 1 2 58170 58172
0 58174 5 1 1 58173
0 58175 7 1 2 89232 58174
0 58176 5 1 1 58175
0 58177 7 1 2 103010 103686
0 58178 5 1 1 58177
0 58179 7 1 2 93303 95952
0 58180 5 1 1 58179
0 58181 7 1 2 58178 58180
0 58182 5 1 1 58181
0 58183 7 1 2 100949 58182
0 58184 5 1 1 58183
0 58185 7 1 2 103313 103379
0 58186 5 1 1 58185
0 58187 7 1 2 67758 88024
0 58188 5 1 1 58187
0 58189 7 1 2 58186 58188
0 58190 5 1 1 58189
0 58191 7 1 2 71454 58190
0 58192 5 1 1 58191
0 58193 7 1 2 71087 97548
0 58194 7 1 2 102900 58193
0 58195 5 1 1 58194
0 58196 7 1 2 58192 58195
0 58197 5 1 1 58196
0 58198 7 1 2 99449 58197
0 58199 5 1 1 58198
0 58200 7 1 2 58184 58199
0 58201 7 1 2 58176 58200
0 58202 7 1 2 58161 58201
0 58203 5 1 1 58202
0 58204 7 1 2 69458 58203
0 58205 5 1 1 58204
0 58206 7 1 2 73094 72231
0 58207 7 1 2 95508 58206
0 58208 7 1 2 89233 58207
0 58209 7 1 2 99058 58208
0 58210 5 1 1 58209
0 58211 7 1 2 58205 58210
0 58212 7 1 2 58127 58211
0 58213 5 1 1 58212
0 58214 7 1 2 84420 58213
0 58215 5 1 1 58214
0 58216 7 1 2 58031 58215
0 58217 7 1 2 57902 58216
0 58218 7 1 2 57772 58217
0 58219 7 1 2 57606 58218
0 58220 7 1 2 57426 58219
0 58221 5 1 1 58220
0 58222 7 1 2 70171 58221
0 58223 5 1 1 58222
0 58224 7 1 2 57119 58223
0 58225 5 1 1 58224
0 58226 7 1 2 56530 58225
0 58227 5 1 1 58226
0 58228 7 1 2 56528 58227
0 58229 7 1 2 54348 58228
0 58230 7 1 2 51121 58229
0 58231 7 1 2 62246 12491
0 58232 5 1 1 58231
0 58233 7 1 2 71877 58232
0 58234 5 1 1 58233
0 58235 7 1 2 71620 84296
0 58236 7 1 2 86268 58235
0 58237 5 1 1 58236
0 58238 7 1 2 58234 58237
0 58239 5 1 1 58238
0 58240 7 1 2 77000 58239
0 58241 5 1 1 58240
0 58242 7 1 2 89704 94157
0 58243 5 1 1 58242
0 58244 7 1 2 58241 58243
0 58245 5 1 1 58244
0 58246 7 1 2 65005 58245
0 58247 5 1 1 58246
0 58248 7 1 2 71878 72404
0 58249 5 1 1 58248
0 58250 7 1 2 70793 76634
0 58251 5 1 1 58250
0 58252 7 1 2 58249 58251
0 58253 5 1 1 58252
0 58254 7 1 2 71455 58253
0 58255 5 1 1 58254
0 58256 7 1 2 58247 58255
0 58257 5 1 1 58256
0 58258 7 1 2 97682 58257
0 58259 5 1 1 58258
0 58260 7 1 2 89075 92617
0 58261 5 1 1 58260
0 58262 7 1 2 79702 85978
0 58263 5 1 1 58262
0 58264 7 1 2 58261 58263
0 58265 5 2 1 58264
0 58266 7 1 2 71879 99134
0 58267 7 1 2 103701 58266
0 58268 5 1 1 58267
0 58269 7 1 2 58259 58268
0 58270 5 1 1 58269
0 58271 7 1 2 63652 58270
0 58272 5 1 1 58271
0 58273 7 3 2 91350 99807
0 58274 7 1 2 71606 90545
0 58275 5 1 1 58274
0 58276 7 1 2 71272 75428
0 58277 7 1 2 94339 58276
0 58278 5 1 1 58277
0 58279 7 1 2 58275 58278
0 58280 5 1 1 58279
0 58281 7 1 2 68492 58280
0 58282 5 1 1 58281
0 58283 7 1 2 65606 89705
0 58284 7 1 2 73888 58283
0 58285 5 1 1 58284
0 58286 7 1 2 58282 58285
0 58287 5 1 1 58286
0 58288 7 1 2 103703 58287
0 58289 5 1 1 58288
0 58290 7 1 2 58272 58289
0 58291 5 1 1 58290
0 58292 7 1 2 63401 58291
0 58293 5 1 1 58292
0 58294 7 1 2 70794 100170
0 58295 5 1 1 58294
0 58296 7 1 2 71880 100180
0 58297 5 1 1 58296
0 58298 7 1 2 58295 58297
0 58299 5 2 1 58298
0 58300 7 1 2 99808 99935
0 58301 7 1 2 103706 58300
0 58302 5 1 1 58301
0 58303 7 1 2 58293 58302
0 58304 5 1 1 58303
0 58305 7 1 2 64813 58304
0 58306 5 1 1 58305
0 58307 7 1 2 89460 99251
0 58308 5 1 1 58307
0 58309 7 1 2 68243 100172
0 58310 5 1 1 58309
0 58311 7 1 2 96894 99246
0 58312 5 1 1 58311
0 58313 7 1 2 58310 58312
0 58314 5 1 1 58313
0 58315 7 1 2 70795 58314
0 58316 5 1 1 58315
0 58317 7 1 2 89490 99243
0 58318 5 1 1 58317
0 58319 7 1 2 76218 72398
0 58320 5 1 1 58319
0 58321 7 1 2 62247 58320
0 58322 5 1 1 58321
0 58323 7 1 2 101470 58322
0 58324 5 1 1 58323
0 58325 7 1 2 90937 58324
0 58326 5 1 1 58325
0 58327 7 1 2 58318 58326
0 58328 7 1 2 58316 58327
0 58329 5 1 1 58328
0 58330 7 1 2 66789 58329
0 58331 5 1 1 58330
0 58332 7 1 2 58308 58331
0 58333 5 1 1 58332
0 58334 7 3 2 64306 79093
0 58335 7 1 2 91351 103708
0 58336 7 1 2 58333 58335
0 58337 5 1 1 58336
0 58338 7 1 2 58306 58337
0 58339 5 1 1 58338
0 58340 7 1 2 70172 58339
0 58341 5 1 1 58340
0 58342 7 1 2 68244 90892
0 58343 5 1 1 58342
0 58344 7 1 2 94839 58343
0 58345 5 1 1 58344
0 58346 7 1 2 70796 58345
0 58347 5 1 1 58346
0 58348 7 1 2 65607 82143
0 58349 7 1 2 101472 58348
0 58350 5 1 1 58349
0 58351 7 1 2 58347 58350
0 58352 5 1 1 58351
0 58353 7 1 2 62248 58352
0 58354 5 1 1 58353
0 58355 7 1 2 71607 98605
0 58356 5 1 1 58355
0 58357 7 1 2 58354 58356
0 58358 5 1 1 58357
0 58359 7 1 2 79193 58358
0 58360 5 1 1 58359
0 58361 7 1 2 81461 103550
0 58362 7 1 2 77649 58361
0 58363 5 1 1 58362
0 58364 7 1 2 58360 58363
0 58365 5 1 1 58364
0 58366 7 1 2 102353 58365
0 58367 5 1 1 58366
0 58368 7 1 2 58341 58367
0 58369 5 1 1 58368
0 58370 7 1 2 63208 58369
0 58371 5 1 1 58370
0 58372 7 1 2 74011 103279
0 58373 5 1 1 58372
0 58374 7 1 2 77133 77414
0 58375 5 1 1 58374
0 58376 7 1 2 71608 82066
0 58377 5 1 1 58376
0 58378 7 1 2 58375 58377
0 58379 5 1 1 58378
0 58380 7 1 2 65608 58379
0 58381 5 1 1 58380
0 58382 7 1 2 58373 58381
0 58383 5 1 1 58382
0 58384 7 1 2 68727 58383
0 58385 5 1 1 58384
0 58386 7 1 2 92087 98960
0 58387 5 1 1 58386
0 58388 7 1 2 58385 58387
0 58389 5 1 1 58388
0 58390 7 1 2 62249 58389
0 58391 5 1 1 58390
0 58392 7 1 2 74894 81502
0 58393 5 1 1 58392
0 58394 7 1 2 71881 87626
0 58395 5 1 1 58394
0 58396 7 1 2 58393 58395
0 58397 5 1 1 58396
0 58398 7 1 2 72402 58397
0 58399 5 1 1 58398
0 58400 7 1 2 58391 58399
0 58401 5 1 1 58400
0 58402 7 1 2 63402 58401
0 58403 5 1 1 58402
0 58404 7 2 2 77687 90896
0 58405 7 1 2 88677 103711
0 58406 5 1 1 58405
0 58407 7 1 2 58403 58406
0 58408 5 1 1 58407
0 58409 7 1 2 69643 58408
0 58410 5 1 1 58409
0 58411 7 1 2 88482 74294
0 58412 7 1 2 97199 58411
0 58413 5 1 1 58412
0 58414 7 1 2 58410 58413
0 58415 5 1 1 58414
0 58416 7 1 2 61923 58415
0 58417 5 1 1 58416
0 58418 7 2 2 77308 95234
0 58419 7 1 2 84130 99927
0 58420 7 1 2 103713 58419
0 58421 5 1 1 58420
0 58422 7 1 2 58417 58421
0 58423 5 1 1 58422
0 58424 7 1 2 101314 58423
0 58425 5 1 1 58424
0 58426 7 1 2 61685 58425
0 58427 7 1 2 58371 58426
0 58428 5 1 1 58427
0 58429 7 1 2 78662 99319
0 58430 7 1 2 98445 58429
0 58431 7 1 2 98719 58430
0 58432 5 1 1 58431
0 58433 7 2 2 72399 21595
0 58434 5 1 1 103715
0 58435 7 1 2 61924 58434
0 58436 5 1 1 58435
0 58437 7 1 2 75866 80388
0 58438 5 1 1 58437
0 58439 7 1 2 58436 58438
0 58440 5 1 1 58439
0 58441 7 1 2 63653 58440
0 58442 5 1 1 58441
0 58443 7 1 2 74162 98961
0 58444 5 1 1 58443
0 58445 7 1 2 58442 58444
0 58446 5 1 1 58445
0 58447 7 1 2 88180 102477
0 58448 7 1 2 58446 58447
0 58449 5 1 1 58448
0 58450 7 1 2 58432 58449
0 58451 5 1 1 58450
0 58452 7 1 2 70173 58451
0 58453 5 1 1 58452
0 58454 7 1 2 82491 97175
0 58455 7 1 2 97683 58454
0 58456 5 1 1 58455
0 58457 7 1 2 58453 58456
0 58458 5 1 1 58457
0 58459 7 1 2 71882 58458
0 58460 5 1 1 58459
0 58461 7 1 2 75038 96362
0 58462 5 1 1 58461
0 58463 7 1 2 96916 58462
0 58464 5 1 1 58463
0 58465 7 1 2 81503 58464
0 58466 5 1 1 58465
0 58467 7 1 2 73362 75039
0 58468 7 1 2 99928 58467
0 58469 5 1 1 58468
0 58470 7 1 2 58466 58469
0 58471 5 1 1 58470
0 58472 7 1 2 94665 98876
0 58473 7 1 2 58471 58472
0 58474 5 1 1 58473
0 58475 7 1 2 58460 58474
0 58476 5 1 1 58475
0 58477 7 1 2 63403 58476
0 58478 5 1 1 58477
0 58479 7 3 2 100126 99066
0 58480 7 1 2 99355 103717
0 58481 7 1 2 103712 58480
0 58482 5 1 1 58481
0 58483 7 1 2 58478 58482
0 58484 5 1 1 58483
0 58485 7 1 2 69644 58484
0 58486 5 1 1 58485
0 58487 7 2 2 95168 101864
0 58488 7 2 2 80686 103720
0 58489 7 1 2 81383 99454
0 58490 7 1 2 103722 58489
0 58491 5 1 1 58490
0 58492 7 1 2 58486 58491
0 58493 5 1 1 58492
0 58494 7 1 2 63209 58493
0 58495 5 1 1 58494
0 58496 7 1 2 93156 100771
0 58497 7 1 2 102017 58496
0 58498 7 1 2 103723 58497
0 58499 5 1 1 58498
0 58500 7 1 2 66574 58499
0 58501 7 1 2 58495 58500
0 58502 5 1 1 58501
0 58503 7 1 2 64601 58502
0 58504 7 1 2 58428 58503
0 58505 5 1 1 58504
0 58506 7 1 2 75979 93971
0 58507 5 1 1 58506
0 58508 7 2 2 77447 58507
0 58509 7 1 2 88568 95837
0 58510 7 1 2 103724 58509
0 58511 5 1 1 58510
0 58512 7 1 2 76828 75863
0 58513 7 1 2 95236 58512
0 58514 7 1 2 95839 58513
0 58515 5 1 1 58514
0 58516 7 1 2 58511 58515
0 58517 5 1 1 58516
0 58518 7 1 2 66790 58517
0 58519 5 1 1 58518
0 58520 7 1 2 80306 95271
0 58521 7 1 2 101428 58520
0 58522 5 1 1 58521
0 58523 7 1 2 58519 58522
0 58524 5 1 1 58523
0 58525 7 2 2 68050 64307
0 58526 7 1 2 92205 103726
0 58527 7 1 2 92917 58526
0 58528 7 1 2 58524 58527
0 58529 5 1 1 58528
0 58530 7 1 2 58505 58529
0 58531 5 1 1 58530
0 58532 7 1 2 69271 58531
0 58533 5 1 1 58532
0 58534 7 1 2 89941 95154
0 58535 7 1 2 88457 58534
0 58536 7 1 2 90088 91352
0 58537 7 1 2 95902 100972
0 58538 7 1 2 58536 58537
0 58539 7 1 2 58535 58538
0 58540 5 1 1 58539
0 58541 7 1 2 58533 58540
0 58542 5 1 1 58541
0 58543 7 1 2 66195 58542
0 58544 5 1 1 58543
0 58545 7 1 2 99536 102376
0 58546 7 1 2 100058 58545
0 58547 5 1 1 58546
0 58548 7 1 2 18134 58547
0 58549 5 1 1 58548
0 58550 7 1 2 62250 58549
0 58551 5 1 1 58550
0 58552 7 1 2 67908 99971
0 58553 7 1 2 99191 58552
0 58554 7 1 2 99642 58553
0 58555 5 1 1 58554
0 58556 7 1 2 58551 58555
0 58557 5 1 1 58556
0 58558 7 1 2 83166 58557
0 58559 5 1 1 58558
0 58560 7 1 2 79783 84594
0 58561 5 1 1 58560
0 58562 7 1 2 82952 79631
0 58563 5 1 1 58562
0 58564 7 1 2 58561 58563
0 58565 5 1 1 58564
0 58566 7 1 2 84803 58565
0 58567 7 1 2 92675 58566
0 58568 5 1 1 58567
0 58569 7 1 2 58559 58568
0 58570 5 1 1 58569
0 58571 7 1 2 79143 58570
0 58572 5 1 1 58571
0 58573 7 2 2 79942 93705
0 58574 7 1 2 88472 89461
0 58575 7 1 2 103728 58574
0 58576 5 1 1 58575
0 58577 7 1 2 58572 58576
0 58578 5 1 1 58577
0 58579 7 1 2 70174 58578
0 58580 5 1 1 58579
0 58581 7 2 2 90782 87168
0 58582 7 1 2 75490 103730
0 58583 5 1 1 58582
0 58584 7 1 2 79194 94934
0 58585 5 1 1 58584
0 58586 7 1 2 58583 58585
0 58587 5 1 1 58586
0 58588 7 1 2 92676 58587
0 58589 5 1 1 58588
0 58590 7 2 2 103623 97467
0 58591 7 1 2 70998 99947
0 58592 7 1 2 103732 58591
0 58593 5 1 1 58592
0 58594 7 1 2 58589 58593
0 58595 5 1 1 58594
0 58596 7 1 2 94877 58595
0 58597 5 1 1 58596
0 58598 7 1 2 67089 103731
0 58599 5 1 1 58598
0 58600 7 1 2 71749 103621
0 58601 5 1 1 58600
0 58602 7 1 2 58599 58601
0 58603 5 1 1 58602
0 58604 7 1 2 63404 58603
0 58605 5 1 1 58604
0 58606 7 1 2 79094 88678
0 58607 7 1 2 79632 58606
0 58608 5 1 1 58607
0 58609 7 1 2 58605 58608
0 58610 5 1 1 58609
0 58611 7 1 2 92677 58610
0 58612 5 1 1 58611
0 58613 7 1 2 62691 103733
0 58614 7 1 2 99950 58613
0 58615 5 1 1 58614
0 58616 7 1 2 58612 58615
0 58617 5 1 1 58616
0 58618 7 1 2 66791 58617
0 58619 5 1 1 58618
0 58620 7 1 2 90160 93196
0 58621 7 1 2 97906 58620
0 58622 7 1 2 93528 58621
0 58623 5 1 1 58622
0 58624 7 1 2 58619 58623
0 58625 5 1 1 58624
0 58626 7 1 2 94950 58625
0 58627 5 1 1 58626
0 58628 7 1 2 58597 58627
0 58629 7 1 2 58580 58628
0 58630 5 1 1 58629
0 58631 7 1 2 69153 58630
0 58632 5 1 1 58631
0 58633 7 1 2 70539 81392
0 58634 7 1 2 102383 58633
0 58635 5 1 1 58634
0 58636 7 2 2 66196 100796
0 58637 7 1 2 63405 99169
0 58638 7 1 2 103734 58637
0 58639 7 2 2 76784 92121
0 58640 7 1 2 102416 103736
0 58641 7 1 2 58638 58640
0 58642 5 1 1 58641
0 58643 7 1 2 58635 58642
0 58644 5 1 1 58643
0 58645 7 1 2 65258 58644
0 58646 5 1 1 58645
0 58647 7 1 2 67836 73839
0 58648 7 1 2 102314 58647
0 58649 7 1 2 103735 100745
0 58650 7 1 2 58648 58649
0 58651 5 1 1 58650
0 58652 7 1 2 58646 58651
0 58653 5 1 1 58652
0 58654 7 1 2 67090 58653
0 58655 5 1 1 58654
0 58656 7 1 2 100748 103658
0 58657 7 1 2 103737 58656
0 58658 7 1 2 94878 58657
0 58659 5 1 1 58658
0 58660 7 1 2 58655 58659
0 58661 5 1 1 58660
0 58662 7 1 2 61925 58661
0 58663 5 1 1 58662
0 58664 7 2 2 76956 79095
0 58665 7 1 2 81462 98577
0 58666 7 1 2 103738 58665
0 58667 7 1 2 101465 58666
0 58668 5 1 1 58667
0 58669 7 1 2 58663 58668
0 58670 5 1 1 58669
0 58671 7 1 2 73268 58670
0 58672 5 1 1 58671
0 58673 7 2 2 79195 97016
0 58674 5 1 1 103740
0 58675 7 1 2 62251 103741
0 58676 5 1 1 58675
0 58677 7 1 2 89784 99859
0 58678 5 1 1 58677
0 58679 7 1 2 58676 58678
0 58680 5 1 1 58679
0 58681 7 1 2 83551 58680
0 58682 5 1 1 58681
0 58683 7 1 2 85315 103739
0 58684 5 1 1 58683
0 58685 7 1 2 78274 98903
0 58686 5 1 1 58685
0 58687 7 1 2 58674 58686
0 58688 5 1 1 58687
0 58689 7 1 2 94879 58688
0 58690 5 1 1 58689
0 58691 7 1 2 58684 58690
0 58692 7 1 2 58682 58691
0 58693 5 1 1 58692
0 58694 7 1 2 100164 58693
0 58695 5 1 1 58694
0 58696 7 1 2 83360 95818
0 58697 5 1 1 58696
0 58698 7 1 2 79109 89211
0 58699 5 1 1 58698
0 58700 7 1 2 58697 58699
0 58701 5 1 1 58700
0 58702 7 1 2 73139 58701
0 58703 5 1 1 58702
0 58704 7 1 2 68885 82751
0 58705 7 1 2 100148 58704
0 58706 5 1 1 58705
0 58707 7 1 2 58703 58706
0 58708 5 1 1 58707
0 58709 7 2 2 69272 58708
0 58710 7 1 2 62692 90730
0 58711 7 1 2 103742 58710
0 58712 5 1 1 58711
0 58713 7 1 2 58695 58712
0 58714 5 1 1 58713
0 58715 7 1 2 61331 58714
0 58716 5 1 1 58715
0 58717 7 1 2 103743 99457
0 58718 5 1 1 58717
0 58719 7 1 2 66792 96437
0 58720 7 1 2 78734 58719
0 58721 7 1 2 87953 58720
0 58722 7 1 2 91036 58721
0 58723 5 1 1 58722
0 58724 7 1 2 75438 32038
0 58725 5 1 1 58724
0 58726 7 1 2 76957 100121
0 58727 7 1 2 99350 58726
0 58728 7 1 2 58725 58727
0 58729 5 1 1 58728
0 58730 7 1 2 58723 58729
0 58731 5 1 1 58730
0 58732 7 1 2 81393 58731
0 58733 5 1 1 58732
0 58734 7 1 2 58718 58733
0 58735 7 1 2 58716 58734
0 58736 5 1 1 58735
0 58737 7 1 2 64308 58736
0 58738 5 1 1 58737
0 58739 7 1 2 58672 58738
0 58740 7 1 2 58632 58739
0 58741 5 1 1 58740
0 58742 7 1 2 63210 58741
0 58743 5 1 1 58742
0 58744 7 3 2 97796 102377
0 58745 7 1 2 76222 103744
0 58746 5 1 1 58745
0 58747 7 1 2 34651 58746
0 58748 5 1 1 58747
0 58749 7 1 2 78571 58748
0 58750 5 1 1 58749
0 58751 7 1 2 89407 94762
0 58752 7 1 2 81019 58751
0 58753 7 1 2 102378 58752
0 58754 5 1 1 58753
0 58755 7 1 2 58750 58754
0 58756 5 1 1 58755
0 58757 7 1 2 62252 58756
0 58758 5 1 1 58757
0 58759 7 1 2 76785 91703
0 58760 7 2 2 98082 58759
0 58761 5 1 1 103747
0 58762 7 1 2 71548 103748
0 58763 5 1 1 58762
0 58764 7 1 2 58758 58763
0 58765 5 1 1 58764
0 58766 7 1 2 99547 58765
0 58767 5 1 1 58766
0 58768 7 1 2 86067 97541
0 58769 5 1 1 58768
0 58770 7 1 2 67091 99550
0 58771 5 1 1 58770
0 58772 7 1 2 58769 58771
0 58773 5 1 1 58772
0 58774 7 1 2 98026 58773
0 58775 5 1 1 58774
0 58776 7 2 2 99458 99896
0 58777 7 1 2 64309 103749
0 58778 5 1 1 58777
0 58779 7 1 2 58775 58778
0 58780 5 1 1 58779
0 58781 7 1 2 87627 58780
0 58782 5 1 1 58781
0 58783 7 2 2 76786 102364
0 58784 7 1 2 98076 103751
0 58785 5 1 1 58784
0 58786 7 1 2 80307 101310
0 58787 7 1 2 91353 58786
0 58788 5 2 1 58787
0 58789 7 1 2 58785 103753
0 58790 5 1 1 58789
0 58791 7 1 2 93181 58790
0 58792 5 1 1 58791
0 58793 7 3 2 65259 99809
0 58794 7 1 2 88171 98998
0 58795 7 1 2 97017 58794
0 58796 7 1 2 103755 58795
0 58797 5 1 1 58796
0 58798 7 1 2 58792 58797
0 58799 5 1 1 58798
0 58800 7 1 2 87761 58799
0 58801 5 1 1 58800
0 58802 7 1 2 58782 58801
0 58803 7 1 2 58767 58802
0 58804 5 1 1 58803
0 58805 7 1 2 63406 58804
0 58806 5 1 1 58805
0 58807 7 1 2 93648 102372
0 58808 5 1 1 58807
0 58809 7 1 2 93027 94228
0 58810 5 1 1 58809
0 58811 7 1 2 58808 58810
0 58812 5 1 1 58811
0 58813 7 1 2 70175 58812
0 58814 5 1 1 58813
0 58815 7 1 2 65260 99537
0 58816 7 1 2 99643 58815
0 58817 5 1 1 58816
0 58818 7 1 2 58814 58817
0 58819 5 1 1 58818
0 58820 7 1 2 62253 58819
0 58821 5 1 1 58820
0 58822 7 1 2 93168 98578
0 58823 7 1 2 102537 58822
0 58824 5 1 1 58823
0 58825 7 1 2 58821 58824
0 58826 5 1 1 58825
0 58827 7 1 2 98027 58826
0 58828 5 1 1 58827
0 58829 7 1 2 78735 97018
0 58830 7 1 2 102384 58829
0 58831 5 1 1 58830
0 58832 7 1 2 58828 58831
0 58833 5 1 1 58832
0 58834 7 1 2 88955 58833
0 58835 5 1 1 58834
0 58836 7 1 2 90823 99953
0 58837 5 1 1 58836
0 58838 7 1 2 90455 100045
0 58839 5 1 1 58838
0 58840 7 1 2 58837 58839
0 58841 5 1 1 58840
0 58842 7 1 2 65609 58841
0 58843 5 1 1 58842
0 58844 7 1 2 99978 99837
0 58845 7 1 2 90824 58844
0 58846 5 1 1 58845
0 58847 7 1 2 58843 58846
0 58848 5 1 1 58847
0 58849 7 1 2 63407 58848
0 58850 5 1 1 58849
0 58851 7 1 2 68245 90089
0 58852 7 1 2 98898 58851
0 58853 7 1 2 97157 58852
0 58854 5 1 1 58853
0 58855 7 1 2 58850 58854
0 58856 5 1 1 58855
0 58857 7 1 2 90731 58856
0 58858 5 1 1 58857
0 58859 7 1 2 58835 58858
0 58860 7 1 2 58806 58859
0 58861 5 1 1 58860
0 58862 7 1 2 69645 84469
0 58863 7 1 2 58861 58862
0 58864 5 1 1 58863
0 58865 7 1 2 58743 58864
0 58866 5 1 1 58865
0 58867 7 1 2 61686 58866
0 58868 5 1 1 58867
0 58869 7 1 2 90825 103168
0 58870 5 1 1 58869
0 58871 7 1 2 103752 102374
0 58872 5 1 1 58871
0 58873 7 1 2 103754 58872
0 58874 5 1 1 58873
0 58875 7 1 2 62254 58874
0 58876 5 1 1 58875
0 58877 7 1 2 87628 101390
0 58878 5 1 1 58877
0 58879 7 1 2 58761 58878
0 58880 7 1 2 58876 58879
0 58881 5 1 1 58880
0 58882 7 1 2 66197 58881
0 58883 5 1 1 58882
0 58884 7 1 2 58870 58883
0 58885 5 1 1 58884
0 58886 7 1 2 71549 58885
0 58887 5 1 1 58886
0 58888 7 1 2 76215 103756
0 58889 7 1 2 102489 58888
0 58890 5 1 1 58889
0 58891 7 1 2 58887 58890
0 58892 5 1 1 58891
0 58893 7 1 2 69273 58892
0 58894 5 1 1 58893
0 58895 7 2 2 91354 84545
0 58896 7 1 2 64421 99810
0 58897 7 1 2 80817 58896
0 58898 7 1 2 103758 58897
0 58899 5 1 1 58898
0 58900 7 1 2 58894 58899
0 58901 5 1 1 58900
0 58902 7 1 2 62693 58901
0 58903 5 1 1 58902
0 58904 7 1 2 73102 103757
0 58905 7 1 2 103759 58904
0 58906 5 1 1 58905
0 58907 7 1 2 101394 30727
0 58908 5 1 1 58907
0 58909 7 1 2 61332 58908
0 58910 5 1 1 58909
0 58911 7 1 2 86068 97883
0 58912 5 1 1 58911
0 58913 7 1 2 58910 58912
0 58914 5 1 1 58913
0 58915 7 1 2 78572 93182
0 58916 7 1 2 58914 58915
0 58917 5 1 1 58916
0 58918 7 1 2 58906 58917
0 58919 5 1 1 58918
0 58920 7 1 2 64422 58919
0 58921 5 1 1 58920
0 58922 7 1 2 58903 58921
0 58923 5 1 1 58922
0 58924 7 1 2 63408 58923
0 58925 5 1 1 58924
0 58926 7 1 2 74386 98710
0 58927 5 1 1 58926
0 58928 7 1 2 75172 103745
0 58929 5 1 1 58928
0 58930 7 1 2 58927 58929
0 58931 5 1 1 58930
0 58932 7 1 2 61333 58931
0 58933 5 1 1 58932
0 58934 7 1 2 84117 97884
0 58935 5 1 1 58934
0 58936 7 1 2 58933 58935
0 58937 5 1 1 58936
0 58938 7 1 2 97148 58937
0 58939 5 1 1 58938
0 58940 7 1 2 72394 99170
0 58941 7 1 2 97784 58940
0 58942 5 1 1 58941
0 58943 7 1 2 58939 58942
0 58944 5 1 1 58943
0 58945 7 1 2 70176 88956
0 58946 7 1 2 58944 58945
0 58947 5 1 1 58946
0 58948 7 1 2 58925 58947
0 58949 5 1 1 58948
0 58950 7 1 2 77208 81478
0 58951 7 1 2 58949 58950
0 58952 5 1 1 58951
0 58953 7 1 2 58868 58952
0 58954 5 1 1 58953
0 58955 7 1 2 64602 58954
0 58956 5 1 1 58955
0 58957 7 2 2 76009 75738
0 58958 7 1 2 99882 103760
0 58959 5 1 1 58958
0 58960 7 1 2 75355 92574
0 58961 7 1 2 101217 58960
0 58962 7 1 2 99184 58961
0 58963 5 1 1 58962
0 58964 7 1 2 58959 58963
0 58965 5 1 1 58964
0 58966 7 1 2 65261 58965
0 58967 5 1 1 58966
0 58968 7 1 2 83601 76010
0 58969 7 1 2 98028 58968
0 58970 7 1 2 97158 58969
0 58971 5 1 1 58970
0 58972 7 1 2 58967 58971
0 58973 5 1 1 58972
0 58974 7 1 2 61334 58973
0 58975 5 1 1 58974
0 58976 7 1 2 98211 103761
0 58977 7 1 2 92451 58976
0 58978 7 1 2 95001 58977
0 58979 5 1 1 58978
0 58980 7 1 2 58975 58979
0 58981 5 1 1 58980
0 58982 7 1 2 68246 58981
0 58983 5 1 1 58982
0 58984 7 1 2 78685 80749
0 58985 5 1 1 58984
0 58986 7 1 2 88835 75356
0 58987 5 1 1 58986
0 58988 7 1 2 58985 58987
0 58989 5 1 1 58988
0 58990 7 1 2 67092 58989
0 58991 5 1 1 58990
0 58992 7 1 2 81363 95268
0 58993 5 1 1 58992
0 58994 7 1 2 58991 58993
0 58995 5 1 1 58994
0 58996 7 1 2 71399 87100
0 58997 7 1 2 98673 58996
0 58998 7 1 2 58995 58997
0 58999 5 1 1 58998
0 59000 7 1 2 58983 58999
0 59001 5 1 1 59000
0 59002 7 1 2 66793 59001
0 59003 5 1 1 59002
0 59004 7 1 2 77115 94593
0 59005 7 1 2 91666 59004
0 59006 7 1 2 95840 59005
0 59007 7 1 2 98703 59006
0 59008 5 1 1 59007
0 59009 7 1 2 59003 59008
0 59010 5 1 1 59009
0 59011 7 1 2 70540 59010
0 59012 5 1 1 59011
0 59013 7 1 2 78736 87257
0 59014 5 1 1 59013
0 59015 7 1 2 87605 76678
0 59016 5 1 1 59015
0 59017 7 1 2 59014 59016
0 59018 5 1 1 59017
0 59019 7 1 2 68247 59018
0 59020 5 1 1 59019
0 59021 7 1 2 87606 90174
0 59022 5 1 1 59021
0 59023 7 1 2 59020 59022
0 59024 5 1 1 59023
0 59025 7 1 2 62933 59024
0 59026 5 1 1 59025
0 59027 7 1 2 76011 95466
0 59028 5 1 1 59027
0 59029 7 1 2 59026 59028
0 59030 5 1 1 59029
0 59031 7 1 2 64814 59030
0 59032 5 1 1 59031
0 59033 7 1 2 78737 78721
0 59034 7 1 2 101718 59033
0 59035 5 1 1 59034
0 59036 7 1 2 59032 59035
0 59037 5 1 1 59036
0 59038 7 1 2 97019 98659
0 59039 7 1 2 59037 59038
0 59040 5 1 1 59039
0 59041 7 1 2 59012 59040
0 59042 5 1 1 59041
0 59043 7 1 2 66575 59042
0 59044 5 1 1 59043
0 59045 7 1 2 61335 75739
0 59046 7 2 2 92562 98616
0 59047 7 1 2 91542 102176
0 59048 7 1 2 103762 59047
0 59049 7 1 2 59045 59048
0 59050 7 1 2 90826 59049
0 59051 5 1 1 59050
0 59052 7 1 2 59044 59051
0 59053 5 1 1 59052
0 59054 7 1 2 93143 59053
0 59055 5 1 1 59054
0 59056 7 1 2 58956 59055
0 59057 5 1 1 59056
0 59058 7 1 2 73048 59057
0 59059 5 1 1 59058
0 59060 7 1 2 64603 95881
0 59061 5 1 1 59060
0 59062 7 1 2 82609 87265
0 59063 5 1 1 59062
0 59064 7 1 2 59061 59063
0 59065 5 1 1 59064
0 59066 7 1 2 89898 59065
0 59067 5 1 1 59066
0 59068 7 2 2 76787 84439
0 59069 7 1 2 94816 103764
0 59070 5 1 1 59069
0 59071 7 1 2 59067 59070
0 59072 5 1 1 59071
0 59073 7 1 2 97753 59072
0 59074 5 1 1 59073
0 59075 7 1 2 96352 98706
0 59076 7 1 2 99981 59075
0 59077 7 1 2 93979 59076
0 59078 5 1 1 59077
0 59079 7 1 2 59074 59078
0 59080 5 1 1 59079
0 59081 7 1 2 63409 59080
0 59082 5 1 1 59081
0 59083 7 1 2 96696 103765
0 59084 5 1 1 59083
0 59085 7 1 2 73617 83560
0 59086 7 1 2 95238 59085
0 59087 7 1 2 77018 59086
0 59088 5 1 1 59087
0 59089 7 1 2 59084 59088
0 59090 5 1 1 59089
0 59091 7 1 2 96835 97732
0 59092 7 1 2 59090 59091
0 59093 5 1 1 59092
0 59094 7 1 2 59082 59093
0 59095 5 1 1 59094
0 59096 7 1 2 70797 59095
0 59097 5 1 1 59096
0 59098 7 1 2 95003 97619
0 59099 5 2 1 59098
0 59100 7 2 2 81874 93197
0 59101 7 1 2 83167 97797
0 59102 7 1 2 103768 59101
0 59103 5 1 1 59102
0 59104 7 1 2 103766 59103
0 59105 5 1 1 59104
0 59106 7 1 2 71991 59105
0 59107 5 1 1 59106
0 59108 7 1 2 98183 103769
0 59109 7 1 2 97857 59108
0 59110 5 1 1 59109
0 59111 7 1 2 59107 59110
0 59112 5 1 1 59111
0 59113 7 1 2 68886 59112
0 59114 5 1 1 59113
0 59115 7 1 2 75931 97007
0 59116 5 1 1 59115
0 59117 7 1 2 87316 98899
0 59118 7 1 2 59116 59117
0 59119 5 1 1 59118
0 59120 7 1 2 59114 59119
0 59121 5 1 1 59120
0 59122 7 1 2 65886 59121
0 59123 5 1 1 59122
0 59124 7 1 2 79226 86578
0 59125 7 1 2 103688 59124
0 59126 5 1 1 59125
0 59127 7 1 2 59123 59126
0 59128 5 1 1 59127
0 59129 7 1 2 81104 59128
0 59130 5 1 1 59129
0 59131 7 1 2 59097 59130
0 59132 5 1 1 59131
0 59133 7 1 2 62255 59132
0 59134 5 1 1 59133
0 59135 7 1 2 83168 98810
0 59136 5 1 1 59135
0 59137 7 1 2 70541 81463
0 59138 7 1 2 100046 59137
0 59139 5 1 1 59138
0 59140 7 1 2 59136 59139
0 59141 5 1 1 59140
0 59142 7 1 2 69867 59141
0 59143 5 1 1 59142
0 59144 7 1 2 103767 59143
0 59145 5 1 1 59144
0 59146 7 1 2 67093 59145
0 59147 5 1 1 59146
0 59148 7 1 2 103702 97757
0 59149 5 1 1 59148
0 59150 7 1 2 59147 59149
0 59151 5 1 1 59150
0 59152 7 1 2 62457 59151
0 59153 5 1 1 59152
0 59154 7 2 2 73521 97918
0 59155 7 2 2 94388 103770
0 59156 7 1 2 98830 98226
0 59157 7 1 2 103772 59156
0 59158 5 1 1 59157
0 59159 7 1 2 59153 59158
0 59160 5 1 1 59159
0 59161 7 1 2 91908 59160
0 59162 5 1 1 59161
0 59163 7 1 2 59134 59162
0 59164 5 1 1 59163
0 59165 7 1 2 63654 59164
0 59166 5 1 1 59165
0 59167 7 1 2 98811 97807
0 59168 5 1 1 59167
0 59169 7 1 2 98800 98822
0 59170 5 1 1 59169
0 59171 7 1 2 71273 97754
0 59172 7 1 2 94340 59171
0 59173 5 1 1 59172
0 59174 7 1 2 59170 59173
0 59175 5 1 1 59174
0 59176 7 1 2 84804 59175
0 59177 5 1 1 59176
0 59178 7 1 2 59168 59177
0 59179 5 1 1 59178
0 59180 7 1 2 69868 59179
0 59181 5 1 1 59180
0 59182 7 1 2 62256 87650
0 59183 7 1 2 99569 59182
0 59184 7 1 2 103771 59183
0 59185 5 1 1 59184
0 59186 7 1 2 59181 59185
0 59187 5 1 1 59186
0 59188 7 1 2 61926 59187
0 59189 5 1 1 59188
0 59190 7 2 2 69869 98812
0 59191 7 1 2 85131 82479
0 59192 7 1 2 103774 59191
0 59193 5 1 1 59192
0 59194 7 1 2 59189 59193
0 59195 5 1 1 59194
0 59196 7 1 2 68493 59195
0 59197 5 1 1 59196
0 59198 7 1 2 83070 80375
0 59199 5 1 1 59198
0 59200 7 1 2 65610 92612
0 59201 5 1 1 59200
0 59202 7 1 2 59199 59201
0 59203 5 1 1 59202
0 59204 7 1 2 69870 102407
0 59205 7 1 2 59203 59204
0 59206 5 1 1 59205
0 59207 7 1 2 59197 59206
0 59208 5 1 1 59207
0 59209 7 1 2 81105 59208
0 59210 5 1 1 59209
0 59211 7 1 2 59166 59210
0 59212 5 1 1 59211
0 59213 7 1 2 70177 59212
0 59214 5 1 1 59213
0 59215 7 1 2 86680 98948
0 59216 5 1 1 59215
0 59217 7 1 2 97620 98355
0 59218 5 1 1 59217
0 59219 7 1 2 59216 59218
0 59220 5 1 1 59219
0 59221 7 1 2 69871 59220
0 59222 5 1 1 59221
0 59223 7 1 2 75246 83461
0 59224 7 1 2 103773 59223
0 59225 5 1 1 59224
0 59226 7 1 2 59222 59225
0 59227 5 1 1 59226
0 59228 7 1 2 61927 59227
0 59229 5 1 1 59228
0 59230 7 1 2 77693 97621
0 59231 7 1 2 77650 59230
0 59232 5 1 1 59231
0 59233 7 1 2 59229 59232
0 59234 5 1 1 59233
0 59235 7 1 2 63410 59234
0 59236 5 1 1 59235
0 59237 7 1 2 87592 94893
0 59238 7 1 2 97622 59237
0 59239 7 1 2 90893 59238
0 59240 5 1 1 59239
0 59241 7 1 2 59236 59240
0 59242 5 1 1 59241
0 59243 7 1 2 65262 81106
0 59244 7 1 2 59242 59243
0 59245 5 1 1 59244
0 59246 7 1 2 64815 59245
0 59247 7 1 2 59214 59246
0 59248 5 1 1 59247
0 59249 7 1 2 81850 92505
0 59250 5 1 1 59249
0 59251 7 1 2 14558 59250
0 59252 5 1 1 59251
0 59253 7 1 2 61928 59252
0 59254 5 1 1 59253
0 59255 7 1 2 78521 83425
0 59256 7 1 2 91604 59255
0 59257 5 1 1 59256
0 59258 7 1 2 59254 59257
0 59259 5 1 1 59258
0 59260 7 1 2 67094 59259
0 59261 5 1 1 59260
0 59262 7 1 2 89959 76436
0 59263 5 1 1 59262
0 59264 7 1 2 88539 92231
0 59265 5 1 1 59264
0 59266 7 1 2 59263 59265
0 59267 5 1 1 59266
0 59268 7 1 2 99962 59267
0 59269 5 1 1 59268
0 59270 7 1 2 59261 59269
0 59271 5 1 1 59270
0 59272 7 1 2 63211 59271
0 59273 5 1 1 59272
0 59274 7 1 2 89485 84476
0 59275 7 1 2 91605 59274
0 59276 5 1 1 59275
0 59277 7 1 2 59273 59276
0 59278 5 1 1 59277
0 59279 7 1 2 92221 98163
0 59280 7 1 2 59278 59279
0 59281 5 1 1 59280
0 59282 7 1 2 68887 94389
0 59283 7 1 2 95461 59282
0 59284 7 1 2 101133 59283
0 59285 5 1 1 59284
0 59286 7 1 2 87874 100499
0 59287 7 1 2 90484 59286
0 59288 7 1 2 82926 59287
0 59289 5 1 1 59288
0 59290 7 1 2 59285 59289
0 59291 5 1 1 59290
0 59292 7 1 2 69872 98648
0 59293 7 1 2 59291 59292
0 59294 5 1 1 59293
0 59295 7 1 2 59281 59294
0 59296 5 1 1 59295
0 59297 7 1 2 70542 59296
0 59298 5 1 1 59297
0 59299 7 1 2 91313 98987
0 59300 5 1 1 59299
0 59301 7 1 2 79920 92921
0 59302 7 1 2 92713 59301
0 59303 5 1 1 59302
0 59304 7 1 2 59300 59303
0 59305 5 1 1 59304
0 59306 7 1 2 65006 59305
0 59307 5 1 1 59306
0 59308 7 1 2 82012 79921
0 59309 7 1 2 99402 59308
0 59310 5 1 1 59309
0 59311 7 1 2 59307 59310
0 59312 5 1 1 59311
0 59313 7 1 2 63857 59312
0 59314 5 1 1 59313
0 59315 7 2 2 73363 95882
0 59316 7 1 2 75971 92714
0 59317 7 1 2 103776 59316
0 59318 5 1 1 59317
0 59319 7 1 2 59314 59318
0 59320 5 1 1 59319
0 59321 7 1 2 94390 100724
0 59322 7 1 2 59320 59321
0 59323 5 1 1 59322
0 59324 7 1 2 59298 59323
0 59325 5 1 1 59324
0 59326 7 1 2 66198 59325
0 59327 5 1 1 59326
0 59328 7 1 2 90217 103707
0 59329 5 1 1 59328
0 59330 7 1 2 83169 95332
0 59331 7 1 2 99252 59330
0 59332 5 1 1 59331
0 59333 7 1 2 71750 85023
0 59334 7 1 2 90051 101179
0 59335 7 1 2 59333 59334
0 59336 5 1 1 59335
0 59337 7 1 2 59332 59336
0 59338 7 1 2 59329 59337
0 59339 5 1 1 59338
0 59340 7 1 2 61687 59339
0 59341 5 1 1 59340
0 59342 7 1 2 67316 93955
0 59343 5 1 1 59342
0 59344 7 1 2 82494 103716
0 59345 5 1 1 59344
0 59346 7 1 2 71883 74387
0 59347 7 1 2 59345 59346
0 59348 5 1 1 59347
0 59349 7 1 2 59343 59348
0 59350 5 1 1 59349
0 59351 7 1 2 61929 59350
0 59352 5 1 1 59351
0 59353 7 1 2 71751 103714
0 59354 5 1 1 59353
0 59355 7 1 2 59352 59354
0 59356 5 1 1 59355
0 59357 7 1 2 93479 59356
0 59358 5 1 1 59357
0 59359 7 1 2 59341 59358
0 59360 5 1 1 59359
0 59361 7 1 2 65007 59360
0 59362 5 1 1 59361
0 59363 7 1 2 87651 83525
0 59364 7 1 2 73627 59363
0 59365 7 1 2 90057 59364
0 59366 5 1 1 59365
0 59367 7 1 2 59362 59366
0 59368 5 1 1 59367
0 59369 7 1 2 64604 59368
0 59370 5 1 1 59369
0 59371 7 1 2 70798 98649
0 59372 7 1 2 75716 59371
0 59373 7 1 2 84288 59372
0 59374 7 1 2 103725 59373
0 59375 5 1 1 59374
0 59376 7 1 2 59370 59375
0 59377 5 1 1 59376
0 59378 7 1 2 69274 59377
0 59379 5 1 1 59378
0 59380 7 1 2 75259 78703
0 59381 7 1 2 77625 59380
0 59382 7 1 2 82916 100741
0 59383 7 1 2 59381 59382
0 59384 5 1 1 59383
0 59385 7 1 2 59379 59384
0 59386 5 1 1 59385
0 59387 7 1 2 97733 59386
0 59388 5 1 1 59387
0 59389 7 1 2 59327 59388
0 59390 5 1 1 59389
0 59391 7 1 2 70178 59390
0 59392 5 1 1 59391
0 59393 7 1 2 68728 98806
0 59394 5 1 1 59393
0 59395 7 1 2 63858 32204
0 59396 5 1 1 59395
0 59397 7 1 2 95876 59396
0 59398 7 1 2 59394 59397
0 59399 5 1 1 59398
0 59400 7 1 2 77209 80854
0 59401 7 1 2 103775 59400
0 59402 5 1 1 59401
0 59403 7 1 2 59399 59402
0 59404 5 1 1 59403
0 59405 7 1 2 65611 59404
0 59406 5 1 1 59405
0 59407 7 1 2 80308 94391
0 59408 7 2 2 91606 59407
0 59409 7 1 2 66199 91334
0 59410 7 1 2 103778 59409
0 59411 5 1 1 59410
0 59412 7 1 2 59406 59411
0 59413 5 1 1 59412
0 59414 7 1 2 63411 59413
0 59415 5 1 1 59414
0 59416 7 1 2 81780 83300
0 59417 7 1 2 103779 59416
0 59418 5 1 1 59417
0 59419 7 1 2 59415 59418
0 59420 5 1 1 59419
0 59421 7 1 2 75173 59420
0 59422 5 1 1 59421
0 59423 7 1 2 71752 88793
0 59424 5 1 1 59423
0 59425 7 1 2 27683 59424
0 59426 5 1 1 59425
0 59427 7 1 2 102472 59426
0 59428 5 1 1 59427
0 59429 7 1 2 98804 46977
0 59430 5 1 1 59429
0 59431 7 1 2 92715 59430
0 59432 5 1 1 59431
0 59433 7 1 2 59428 59432
0 59434 5 1 1 59433
0 59435 7 1 2 71884 59434
0 59436 5 1 1 59435
0 59437 7 1 2 98787 102408
0 59438 5 1 1 59437
0 59439 7 1 2 59436 59438
0 59440 5 1 1 59439
0 59441 7 1 2 95883 59440
0 59442 5 1 1 59441
0 59443 7 1 2 66200 88281
0 59444 7 1 2 100032 59443
0 59445 7 1 2 91965 96912
0 59446 7 1 2 59444 59445
0 59447 7 1 2 98904 59446
0 59448 5 1 1 59447
0 59449 7 1 2 59442 59448
0 59450 7 1 2 59422 59449
0 59451 5 1 1 59450
0 59452 7 1 2 91285 59451
0 59453 5 1 1 59452
0 59454 7 1 2 69646 59453
0 59455 7 1 2 59392 59454
0 59456 5 1 1 59455
0 59457 7 1 2 90732 59456
0 59458 7 1 2 59248 59457
0 59459 5 1 1 59458
0 59460 7 1 2 88957 94434
0 59461 5 1 1 59460
0 59462 7 1 2 84867 80309
0 59463 5 1 1 59462
0 59464 7 1 2 59461 59463
0 59465 5 1 1 59464
0 59466 7 1 2 75790 59465
0 59467 5 1 1 59466
0 59468 7 1 2 97921 101430
0 59469 5 1 1 59468
0 59470 7 1 2 59467 59469
0 59471 5 1 1 59470
0 59472 7 1 2 76198 59471
0 59473 5 1 1 59472
0 59474 7 1 2 81287 80634
0 59475 7 1 2 72866 89599
0 59476 7 1 2 59474 59475
0 59477 5 1 1 59476
0 59478 7 1 2 59473 59477
0 59479 5 1 1 59478
0 59480 7 1 2 69647 59479
0 59481 5 1 1 59480
0 59482 7 1 2 77265 79144
0 59483 7 1 2 86448 59482
0 59484 7 1 2 92716 59483
0 59485 5 1 1 59484
0 59486 7 1 2 59481 59485
0 59487 5 1 1 59486
0 59488 7 1 2 61930 59487
0 59489 5 1 1 59488
0 59490 7 1 2 75791 81394
0 59491 5 1 1 59490
0 59492 7 1 2 79096 89491
0 59493 5 1 1 59492
0 59494 7 1 2 59491 59493
0 59495 5 1 1 59494
0 59496 7 1 2 86449 92922
0 59497 7 1 2 59495 59496
0 59498 5 1 1 59497
0 59499 7 1 2 59489 59498
0 59500 5 1 1 59499
0 59501 7 1 2 68729 59500
0 59502 5 1 1 59501
0 59503 7 1 2 61931 87525
0 59504 5 1 1 59503
0 59505 7 1 2 102908 59504
0 59506 5 1 1 59505
0 59507 7 1 2 61688 59506
0 59508 5 1 1 59507
0 59509 7 1 2 84131 96645
0 59510 5 1 1 59509
0 59511 7 1 2 59508 59510
0 59512 5 1 1 59511
0 59513 7 1 2 98988 59512
0 59514 5 1 1 59513
0 59515 7 1 2 84535 92038
0 59516 5 1 1 59515
0 59517 7 1 2 92717 95024
0 59518 5 1 1 59517
0 59519 7 1 2 59516 59518
0 59520 5 1 1 59519
0 59521 7 1 2 79922 59520
0 59522 5 1 1 59521
0 59523 7 1 2 59514 59522
0 59524 5 1 1 59523
0 59525 7 1 2 63859 59524
0 59526 5 1 1 59525
0 59527 7 1 2 92046 94909
0 59528 5 1 1 59527
0 59529 7 1 2 61932 94895
0 59530 5 1 1 59529
0 59531 7 1 2 81395 75840
0 59532 5 1 1 59531
0 59533 7 1 2 89493 59532
0 59534 7 1 2 59530 59533
0 59535 5 1 1 59534
0 59536 7 1 2 63212 59535
0 59537 5 1 1 59536
0 59538 7 1 2 59528 59537
0 59539 5 2 1 59538
0 59540 7 1 2 86769 72894
0 59541 7 1 2 103780 59540
0 59542 5 1 1 59541
0 59543 7 1 2 59526 59542
0 59544 7 1 2 59502 59543
0 59545 5 1 1 59544
0 59546 7 1 2 100725 59545
0 59547 5 1 1 59546
0 59548 7 1 2 80287 86579
0 59549 7 1 2 90943 59548
0 59550 7 1 2 96676 59549
0 59551 5 1 1 59550
0 59552 7 1 2 81865 96509
0 59553 7 1 2 92721 59552
0 59554 5 1 1 59553
0 59555 7 1 2 59551 59554
0 59556 5 1 1 59555
0 59557 7 1 2 62934 59556
0 59558 5 1 1 59557
0 59559 7 1 2 88642 100733
0 59560 7 1 2 103781 59559
0 59561 5 1 1 59560
0 59562 7 1 2 59558 59561
0 59563 5 1 1 59562
0 59564 7 1 2 85715 59563
0 59565 5 1 1 59564
0 59566 7 1 2 59547 59565
0 59567 5 1 1 59566
0 59568 7 1 2 98029 59567
0 59569 5 1 1 59568
0 59570 7 2 2 86461 94921
0 59571 7 1 2 83744 103782
0 59572 5 1 1 59571
0 59573 7 1 2 81703 71757
0 59574 7 1 2 91996 59573
0 59575 5 1 1 59574
0 59576 7 1 2 59572 59575
0 59577 5 1 1 59576
0 59578 7 1 2 66794 59577
0 59579 5 1 1 59578
0 59580 7 1 2 81781 82177
0 59581 5 1 1 59580
0 59582 7 1 2 65612 89624
0 59583 5 1 1 59582
0 59584 7 1 2 59581 59583
0 59585 5 1 1 59584
0 59586 7 1 2 61689 59585
0 59587 5 1 1 59586
0 59588 7 1 2 76788 93480
0 59589 5 1 1 59588
0 59590 7 1 2 59587 59589
0 59591 5 1 1 59590
0 59592 7 1 2 86035 59591
0 59593 5 1 1 59592
0 59594 7 1 2 59579 59593
0 59595 5 1 1 59594
0 59596 7 1 2 68494 59595
0 59597 5 1 1 59596
0 59598 7 1 2 95664 102131
0 59599 7 1 2 96124 59598
0 59600 5 1 1 59599
0 59601 7 1 2 59597 59600
0 59602 5 1 1 59601
0 59603 7 1 2 67095 59602
0 59604 5 1 1 59603
0 59605 7 1 2 95583 103700
0 59606 5 1 1 59605
0 59607 7 1 2 10838 59606
0 59608 5 1 1 59607
0 59609 7 1 2 61933 59608
0 59610 5 1 1 59609
0 59611 7 1 2 76012 75828
0 59612 5 1 1 59611
0 59613 7 1 2 59610 59612
0 59614 5 1 1 59613
0 59615 7 1 2 68248 59614
0 59616 5 1 1 59615
0 59617 7 1 2 76679 95993
0 59618 7 1 2 82980 59617
0 59619 5 1 1 59618
0 59620 7 1 2 59616 59619
0 59621 5 1 1 59620
0 59622 7 1 2 61690 59621
0 59623 5 1 1 59622
0 59624 7 1 2 81782 97214
0 59625 5 1 1 59624
0 59626 7 1 2 59623 59625
0 59627 5 1 1 59626
0 59628 7 1 2 93741 59627
0 59629 5 1 1 59628
0 59630 7 1 2 59604 59629
0 59631 5 1 1 59630
0 59632 7 1 2 69648 59631
0 59633 5 1 1 59632
0 59634 7 1 2 74388 79519
0 59635 5 1 1 59634
0 59636 7 1 2 68495 76027
0 59637 5 1 1 59636
0 59638 7 1 2 33001 59637
0 59639 5 1 1 59638
0 59640 7 1 2 63412 59639
0 59641 7 1 2 59635 59640
0 59642 5 1 1 59641
0 59643 7 1 2 68249 99289
0 59644 5 1 1 59643
0 59645 7 1 2 59642 59644
0 59646 5 1 1 59645
0 59647 7 1 2 83836 79156
0 59648 7 1 2 59646 59647
0 59649 5 1 1 59648
0 59650 7 1 2 59633 59649
0 59651 5 1 1 59650
0 59652 7 1 2 71992 59651
0 59653 5 1 1 59652
0 59654 7 1 2 95063 26343
0 59655 5 1 1 59654
0 59656 7 1 2 82013 59655
0 59657 5 1 1 59656
0 59658 7 1 2 97212 59657
0 59659 5 1 1 59658
0 59660 7 1 2 64605 59659
0 59661 5 1 1 59660
0 59662 7 1 2 82024 99888
0 59663 5 1 1 59662
0 59664 7 1 2 59661 59663
0 59665 5 1 1 59664
0 59666 7 1 2 71885 59665
0 59667 5 1 1 59666
0 59668 7 2 2 84440 96284
0 59669 7 1 2 102902 103784
0 59670 5 1 1 59669
0 59671 7 1 2 59667 59670
0 59672 5 1 1 59671
0 59673 7 1 2 73364 59672
0 59674 5 1 1 59673
0 59675 7 1 2 88051 101731
0 59676 7 1 2 94288 59675
0 59677 5 1 1 59676
0 59678 7 1 2 59674 59677
0 59679 5 1 1 59678
0 59680 7 1 2 76199 59679
0 59681 5 1 1 59680
0 59682 7 1 2 77266 103785
0 59683 5 1 1 59682
0 59684 7 1 2 83840 15353
0 59685 5 1 1 59684
0 59686 7 1 2 91637 59685
0 59687 5 1 1 59686
0 59688 7 1 2 59683 59687
0 59689 5 1 1 59688
0 59690 7 1 2 73365 59689
0 59691 5 1 1 59690
0 59692 7 1 2 83837 74281
0 59693 7 1 2 94289 59692
0 59694 5 1 1 59693
0 59695 7 1 2 59691 59694
0 59696 5 1 1 59695
0 59697 7 1 2 95896 59696
0 59698 5 1 1 59697
0 59699 7 1 2 83634 73701
0 59700 5 1 1 59699
0 59701 7 1 2 83920 59700
0 59702 5 1 1 59701
0 59703 7 1 2 81002 59702
0 59704 5 1 1 59703
0 59705 7 1 2 82933 94817
0 59706 5 1 1 59705
0 59707 7 1 2 59704 59706
0 59708 5 1 1 59707
0 59709 7 1 2 63413 84719
0 59710 7 1 2 88055 59709
0 59711 7 1 2 59708 59710
0 59712 5 1 1 59711
0 59713 7 1 2 59698 59712
0 59714 7 1 2 59681 59713
0 59715 5 1 1 59714
0 59716 7 1 2 70543 59715
0 59717 5 1 1 59716
0 59718 7 1 2 103783 101286
0 59719 5 1 1 59718
0 59720 7 2 2 76789 98971
0 59721 7 1 2 73170 96397
0 59722 7 1 2 103786 59721
0 59723 5 1 1 59722
0 59724 7 1 2 59719 59723
0 59725 5 1 1 59724
0 59726 7 1 2 66795 59725
0 59727 5 1 1 59726
0 59728 7 1 2 81107 85461
0 59729 7 2 2 84490 59728
0 59730 5 1 1 103788
0 59731 7 1 2 74871 103789
0 59732 5 1 1 59731
0 59733 7 1 2 59727 59732
0 59734 5 1 1 59733
0 59735 7 1 2 67096 59734
0 59736 5 1 1 59735
0 59737 7 1 2 75601 89551
0 59738 7 1 2 103787 59737
0 59739 5 1 1 59738
0 59740 7 1 2 59730 59739
0 59741 5 1 1 59740
0 59742 7 1 2 88516 59741
0 59743 5 1 1 59742
0 59744 7 1 2 59736 59743
0 59745 5 1 1 59744
0 59746 7 1 2 69649 59745
0 59747 5 1 1 59746
0 59748 7 1 2 83745 82398
0 59749 7 1 2 91658 59748
0 59750 7 1 2 99129 59749
0 59751 5 1 1 59750
0 59752 7 1 2 59747 59751
0 59753 7 1 2 59717 59752
0 59754 7 1 2 59653 59753
0 59755 5 1 1 59754
0 59756 7 1 2 97684 59755
0 59757 5 1 1 59756
0 59758 7 1 2 59569 59757
0 59759 5 1 1 59758
0 59760 7 1 2 70179 59759
0 59761 5 1 1 59760
0 59762 7 1 2 61691 99890
0 59763 5 1 1 59762
0 59764 7 1 2 61934 95841
0 59765 5 1 1 59764
0 59766 7 1 2 62935 93373
0 59767 5 1 1 59766
0 59768 7 1 2 59765 59767
0 59769 5 1 1 59768
0 59770 7 1 2 90284 59769
0 59771 5 1 1 59770
0 59772 7 1 2 59763 59771
0 59773 5 1 1 59772
0 59774 7 1 2 76490 59773
0 59775 5 1 1 59774
0 59776 7 1 2 84152 87551
0 59777 7 1 2 88052 59776
0 59778 5 1 1 59777
0 59779 7 1 2 59775 59778
0 59780 5 1 1 59779
0 59781 7 1 2 95609 59780
0 59782 5 1 1 59781
0 59783 7 1 2 68250 16991
0 59784 5 1 1 59783
0 59785 7 1 2 63414 92042
0 59786 5 1 1 59785
0 59787 7 1 2 86777 59786
0 59788 7 1 2 59784 59787
0 59789 5 1 1 59788
0 59790 7 1 2 63860 98751
0 59791 5 1 1 59790
0 59792 7 1 2 85673 59791
0 59793 5 1 1 59792
0 59794 7 1 2 65887 102015
0 59795 7 1 2 59793 59794
0 59796 5 1 1 59795
0 59797 7 1 2 59789 59796
0 59798 5 1 1 59797
0 59799 7 1 2 64606 59798
0 59800 5 1 1 59799
0 59801 7 1 2 85015 90870
0 59802 7 1 2 79328 59801
0 59803 7 1 2 76491 59802
0 59804 5 1 1 59803
0 59805 7 1 2 59800 59804
0 59806 5 1 1 59805
0 59807 7 1 2 63213 59806
0 59808 5 1 1 59807
0 59809 7 1 2 59782 59808
0 59810 5 1 1 59809
0 59811 7 1 2 70544 59810
0 59812 5 1 1 59811
0 59813 7 1 2 83251 86681
0 59814 5 1 1 59813
0 59815 7 1 2 6849 82215
0 59816 5 1 1 59815
0 59817 7 1 2 65888 59816
0 59818 5 1 1 59817
0 59819 7 1 2 71993 74389
0 59820 7 1 2 33253 59819
0 59821 5 1 1 59820
0 59822 7 1 2 59818 59821
0 59823 5 1 1 59822
0 59824 7 1 2 64607 59823
0 59825 7 1 2 95025 59824
0 59826 5 1 1 59825
0 59827 7 1 2 59814 59826
0 59828 5 1 1 59827
0 59829 7 1 2 65613 59828
0 59830 5 1 1 59829
0 59831 7 1 2 79145 90543
0 59832 5 1 1 59831
0 59833 7 1 2 91196 83184
0 59834 7 1 2 97291 59833
0 59835 5 1 1 59834
0 59836 7 1 2 59832 59835
0 59837 5 1 1 59836
0 59838 7 1 2 66796 59837
0 59839 5 1 1 59838
0 59840 7 1 2 82403 97950
0 59841 5 1 1 59840
0 59842 7 1 2 59839 59841
0 59843 5 1 1 59842
0 59844 7 1 2 101942 59843
0 59845 5 1 1 59844
0 59846 7 1 2 59830 59845
0 59847 5 1 1 59846
0 59848 7 1 2 63415 59847
0 59849 5 1 1 59848
0 59850 7 1 2 86682 91768
0 59851 5 1 1 59850
0 59852 7 1 2 74408 91200
0 59853 7 1 2 91461 59852
0 59854 5 1 1 59853
0 59855 7 1 2 59851 59854
0 59856 5 1 1 59855
0 59857 7 1 2 81783 71088
0 59858 7 1 2 59856 59857
0 59859 5 1 1 59858
0 59860 7 1 2 59849 59859
0 59861 7 1 2 59812 59860
0 59862 5 1 1 59861
0 59863 7 1 2 97685 59862
0 59864 5 1 1 59863
0 59865 7 1 2 103777 98609
0 59866 5 1 1 59865
0 59867 7 1 2 89125 80310
0 59868 5 1 1 59867
0 59869 7 1 2 86580 96333
0 59870 5 1 1 59869
0 59871 7 1 2 59868 59870
0 59872 5 1 1 59871
0 59873 7 1 2 61935 59872
0 59874 5 1 1 59873
0 59875 7 1 2 74554 90499
0 59876 5 1 1 59875
0 59877 7 1 2 59874 59876
0 59878 5 1 1 59877
0 59879 7 1 2 79914 59878
0 59880 5 1 1 59879
0 59881 7 1 2 70545 80611
0 59882 7 1 2 102135 59881
0 59883 5 1 1 59882
0 59884 7 1 2 59880 59883
0 59885 5 1 1 59884
0 59886 7 1 2 61692 75174
0 59887 7 1 2 59885 59886
0 59888 5 1 1 59887
0 59889 7 1 2 59866 59888
0 59890 5 1 1 59889
0 59891 7 1 2 69650 59890
0 59892 5 1 1 59891
0 59893 7 1 2 84820 80656
0 59894 7 1 2 102052 59893
0 59895 7 1 2 95418 59894
0 59896 5 1 1 59895
0 59897 7 1 2 59892 59896
0 59898 5 1 1 59897
0 59899 7 1 2 90690 100727
0 59900 7 1 2 59898 59899
0 59901 5 1 1 59900
0 59902 7 1 2 59864 59901
0 59903 5 1 1 59902
0 59904 7 1 2 65263 59903
0 59905 5 1 1 59904
0 59906 7 1 2 75175 102820
0 59907 5 1 1 59906
0 59908 7 1 2 86618 95823
0 59909 5 1 1 59908
0 59910 7 1 2 59907 59909
0 59911 5 1 1 59910
0 59912 7 1 2 103746 59911
0 59913 5 1 1 59912
0 59914 7 1 2 63655 86394
0 59915 7 1 2 94740 59914
0 59916 7 1 2 92206 59915
0 59917 5 1 1 59916
0 59918 7 1 2 59913 59917
0 59919 5 1 1 59918
0 59920 7 1 2 71706 59919
0 59921 5 1 1 59920
0 59922 7 2 2 85685 98221
0 59923 7 1 2 99446 99811
0 59924 7 1 2 103790 59923
0 59925 5 1 1 59924
0 59926 7 1 2 59921 59925
0 59927 5 1 1 59926
0 59928 7 1 2 61936 59927
0 59929 5 1 1 59928
0 59930 7 1 2 103709 103791
0 59931 5 1 1 59930
0 59932 7 1 2 76829 86231
0 59933 7 1 2 98191 59932
0 59934 5 1 1 59933
0 59935 7 1 2 59931 59934
0 59936 5 1 1 59935
0 59937 7 1 2 88524 59936
0 59938 5 1 1 59937
0 59939 7 1 2 59929 59938
0 59940 5 1 1 59939
0 59941 7 1 2 63416 59940
0 59942 5 1 1 59941
0 59943 7 1 2 82059 81851
0 59944 7 1 2 85686 59943
0 59945 7 1 2 103710 99937
0 59946 7 1 2 59944 59945
0 59947 5 1 1 59946
0 59948 7 1 2 59942 59947
0 59949 5 1 1 59948
0 59950 7 1 2 83824 59949
0 59951 5 1 1 59950
0 59952 7 1 2 74976 91873
0 59953 7 1 2 89867 59952
0 59954 7 1 2 99174 59953
0 59955 7 1 2 89221 59954
0 59956 5 1 1 59955
0 59957 7 1 2 91712 103696
0 59958 5 1 1 59957
0 59959 7 1 2 83838 89456
0 59960 5 1 1 59959
0 59961 7 1 2 59958 59960
0 59962 5 1 1 59961
0 59963 7 1 2 68496 98342
0 59964 7 1 2 99146 59963
0 59965 7 1 2 59962 59964
0 59966 5 1 1 59965
0 59967 7 1 2 59956 59966
0 59968 5 1 1 59967
0 59969 7 1 2 74586 59968
0 59970 5 1 1 59969
0 59971 7 1 2 6347 25950
0 59972 5 1 1 59971
0 59973 7 1 2 91818 98440
0 59974 7 1 2 103697 103763
0 59975 7 1 2 59973 59974
0 59976 7 1 2 59972 59975
0 59977 5 1 1 59976
0 59978 7 1 2 59970 59977
0 59979 7 1 2 59951 59978
0 59980 5 1 1 59979
0 59981 7 1 2 70180 59980
0 59982 5 1 1 59981
0 59983 7 1 2 87383 84200
0 59984 7 1 2 103704 59983
0 59985 5 1 1 59984
0 59986 7 1 2 91884 99171
0 59987 7 1 2 83021 59986
0 59988 7 1 2 100843 59987
0 59989 5 1 1 59988
0 59990 7 1 2 59985 59989
0 59991 5 1 1 59990
0 59992 7 1 2 62458 59991
0 59993 5 1 1 59992
0 59994 7 1 2 99172 97919
0 59995 7 1 2 103382 97468
0 59996 7 1 2 59994 59995
0 59997 5 1 1 59996
0 59998 7 1 2 59993 59997
0 59999 5 1 1 59998
0 60000 7 1 2 63214 59999
0 60001 5 1 1 60000
0 60002 7 1 2 97492 103727
0 60003 7 2 2 67097 98492
0 60004 7 1 2 102829 103792
0 60005 7 1 2 60002 60004
0 60006 5 1 1 60005
0 60007 7 1 2 60001 60006
0 60008 5 1 1 60007
0 60009 7 1 2 61937 60008
0 60010 5 1 1 60009
0 60011 7 1 2 101783 99865
0 60012 7 1 2 103144 103793
0 60013 7 1 2 60011 60012
0 60014 5 1 1 60013
0 60015 7 1 2 60010 60014
0 60016 5 1 1 60015
0 60017 7 1 2 81704 79007
0 60018 7 1 2 60016 60017
0 60019 5 1 1 60018
0 60020 7 1 2 59982 60019
0 60021 5 1 1 60020
0 60022 7 1 2 73522 60021
0 60023 5 1 1 60022
0 60024 7 1 2 59905 60023
0 60025 7 1 2 59761 60024
0 60026 5 1 1 60025
0 60027 7 1 2 64423 60026
0 60028 5 1 1 60027
0 60029 7 1 2 92733 95360
0 60030 7 1 2 101108 60029
0 60031 7 1 2 77156 80684
0 60032 7 1 2 102225 60031
0 60033 7 1 2 60030 60032
0 60034 5 1 1 60033
0 60035 7 1 2 60028 60034
0 60036 5 1 1 60035
0 60037 7 1 2 61336 60036
0 60038 5 1 1 60037
0 60039 7 1 2 91874 92748
0 60040 7 1 2 101043 98136
0 60041 7 1 2 60039 60040
0 60042 5 1 1 60041
0 60043 7 1 2 70546 99222
0 60044 7 1 2 103718 60043
0 60045 7 1 2 90910 60044
0 60046 5 1 1 60045
0 60047 7 1 2 60042 60046
0 60048 5 1 1 60047
0 60049 7 1 2 64608 60048
0 60050 5 1 1 60049
0 60051 7 1 2 85657 79231
0 60052 7 1 2 91833 97569
0 60053 7 1 2 98137 60052
0 60054 7 1 2 60051 60053
0 60055 5 1 1 60054
0 60056 7 1 2 60050 60055
0 60057 5 1 1 60056
0 60058 7 1 2 70181 60057
0 60059 5 1 1 60058
0 60060 7 1 2 88073 95734
0 60061 5 1 1 60060
0 60062 7 1 2 88936 77645
0 60063 5 1 1 60062
0 60064 7 1 2 60061 60063
0 60065 5 1 1 60064
0 60066 7 1 2 97819 102354
0 60067 7 1 2 60065 60066
0 60068 5 1 1 60067
0 60069 7 1 2 60059 60068
0 60070 5 1 1 60069
0 60071 7 1 2 61693 60070
0 60072 5 1 1 60071
0 60073 7 1 2 83552 89991
0 60074 5 1 1 60073
0 60075 7 1 2 8475 60074
0 60076 5 1 1 60075
0 60077 7 1 2 91725 60076
0 60078 5 1 1 60077
0 60079 7 1 2 76765 79538
0 60080 7 1 2 87660 60079
0 60081 5 1 1 60080
0 60082 7 1 2 60078 60081
0 60083 5 1 1 60082
0 60084 7 1 2 90803 97686
0 60085 7 1 2 60083 60084
0 60086 5 1 1 60085
0 60087 7 1 2 60072 60086
0 60088 5 1 1 60087
0 60089 7 1 2 64816 60088
0 60090 5 1 1 60089
0 60091 7 1 2 88815 96320
0 60092 5 1 1 60091
0 60093 7 1 2 89331 90788
0 60094 5 1 1 60093
0 60095 7 1 2 60092 60094
0 60096 5 1 1 60095
0 60097 7 1 2 99747 60096
0 60098 5 1 1 60097
0 60099 7 2 2 63861 82941
0 60100 7 1 2 77267 99092
0 60101 7 1 2 89217 60100
0 60102 7 1 2 103794 60101
0 60103 5 1 1 60102
0 60104 7 1 2 60098 60103
0 60105 5 1 1 60104
0 60106 7 1 2 90630 60105
0 60107 5 1 1 60106
0 60108 7 1 2 87567 98452
0 60109 7 1 2 102157 103795
0 60110 7 1 2 60108 60109
0 60111 5 1 1 60110
0 60112 7 1 2 60107 60111
0 60113 5 1 1 60112
0 60114 7 1 2 62257 85107
0 60115 7 1 2 94741 60114
0 60116 7 1 2 60113 60115
0 60117 5 1 1 60116
0 60118 7 1 2 60090 60117
0 60119 5 1 1 60118
0 60120 7 1 2 69873 60119
0 60121 5 1 1 60120
0 60122 7 1 2 79460 92903
0 60123 5 1 1 60122
0 60124 7 1 2 92269 60123
0 60125 5 1 1 60124
0 60126 7 1 2 86818 60125
0 60127 5 1 1 60126
0 60128 7 1 2 61694 86341
0 60129 5 1 1 60128
0 60130 7 1 2 79232 86462
0 60131 5 1 1 60130
0 60132 7 1 2 60129 60131
0 60133 5 1 1 60132
0 60134 7 1 2 78964 60133
0 60135 5 1 1 60134
0 60136 7 1 2 80841 82924
0 60137 5 1 1 60136
0 60138 7 1 2 19867 60137
0 60139 5 1 1 60138
0 60140 7 1 2 99976 60139
0 60141 5 1 1 60140
0 60142 7 1 2 60135 60141
0 60143 5 1 1 60142
0 60144 7 1 2 82472 60143
0 60145 5 1 1 60144
0 60146 7 1 2 60127 60145
0 60147 5 1 1 60146
0 60148 7 1 2 77102 101391
0 60149 7 1 2 60147 60148
0 60150 5 1 1 60149
0 60151 7 1 2 60121 60150
0 60152 5 1 1 60151
0 60153 7 1 2 93633 60152
0 60154 5 1 1 60153
0 60155 7 1 2 82144 86086
0 60156 5 1 1 60155
0 60157 7 1 2 78625 90938
0 60158 5 1 1 60157
0 60159 7 1 2 60156 60158
0 60160 5 2 1 60159
0 60161 7 1 2 88199 103796
0 60162 5 1 1 60161
0 60163 7 2 2 63215 88424
0 60164 7 1 2 102110 103798
0 60165 5 1 1 60164
0 60166 7 1 2 60162 60165
0 60167 5 1 1 60166
0 60168 7 1 2 61938 60167
0 60169 5 1 1 60168
0 60170 7 1 2 78522 81396
0 60171 7 1 2 103799 60170
0 60172 5 1 1 60171
0 60173 7 1 2 60169 60172
0 60174 5 1 1 60173
0 60175 7 1 2 75792 99566
0 60176 7 1 2 90733 60175
0 60177 7 1 2 60174 60176
0 60178 5 1 1 60177
0 60179 7 1 2 61337 60178
0 60180 7 1 2 60154 60179
0 60181 5 1 1 60180
0 60182 7 1 2 82685 100719
0 60183 7 1 2 91589 60182
0 60184 7 1 2 98168 60183
0 60185 5 1 1 60184
0 60186 7 1 2 88403 92057
0 60187 5 1 1 60186
0 60188 7 1 2 83574 60187
0 60189 5 1 1 60188
0 60190 7 1 2 77323 94392
0 60191 7 1 2 90734 60190
0 60192 7 1 2 60189 60191
0 60193 5 1 1 60192
0 60194 7 1 2 60185 60193
0 60195 5 1 1 60194
0 60196 7 1 2 76912 60195
0 60197 5 1 1 60196
0 60198 7 1 2 77157 88172
0 60199 7 1 2 102144 60198
0 60200 7 1 2 98482 60199
0 60201 5 1 1 60200
0 60202 7 1 2 60197 60201
0 60203 5 1 1 60202
0 60204 7 1 2 66797 60203
0 60205 5 1 1 60204
0 60206 7 1 2 99567 103719
0 60207 7 1 2 100658 60206
0 60208 7 1 2 88425 60207
0 60209 5 1 1 60208
0 60210 7 1 2 60205 60209
0 60211 5 1 1 60210
0 60212 7 1 2 64817 60211
0 60213 5 1 1 60212
0 60214 7 1 2 89113 96241
0 60215 5 1 1 60214
0 60216 7 1 2 79613 87098
0 60217 7 1 2 90963 98650
0 60218 7 1 2 60216 60217
0 60219 5 1 1 60218
0 60220 7 1 2 60215 60219
0 60221 5 1 1 60220
0 60222 7 1 2 76541 98878
0 60223 7 1 2 60221 60222
0 60224 5 1 1 60223
0 60225 7 1 2 60213 60224
0 60226 5 1 1 60225
0 60227 7 1 2 69874 60226
0 60228 5 1 1 60227
0 60229 7 1 2 94742 102194
0 60230 7 1 2 101501 60229
0 60231 7 1 2 76924 90182
0 60232 5 1 1 60231
0 60233 7 1 2 88426 90218
0 60234 7 1 2 60232 60233
0 60235 7 1 2 60230 60234
0 60236 5 1 1 60235
0 60237 7 1 2 60228 60236
0 60238 5 1 1 60237
0 60239 7 1 2 61695 60238
0 60240 5 1 1 60239
0 60241 7 1 2 86036 81479
0 60242 7 1 2 93701 98637
0 60243 7 1 2 60241 60242
0 60244 7 1 2 92207 60243
0 60245 7 1 2 103797 60244
0 60246 5 1 1 60245
0 60247 7 1 2 66201 60246
0 60248 7 1 2 60240 60247
0 60249 5 1 1 60248
0 60250 7 1 2 71400 60249
0 60251 7 1 2 60181 60250
0 60252 5 1 1 60251
0 60253 7 1 2 60038 60252
0 60254 7 1 2 59459 60253
0 60255 7 1 2 59059 60254
0 60256 7 1 2 58544 60255
0 60257 5 1 1 60256
0 60258 7 1 2 72685 60257
0 60259 5 1 1 60258
0 60260 7 1 2 65614 97403
0 60261 5 1 1 60260
0 60262 7 1 2 90735 97428
0 60263 7 1 2 97411 60262
0 60264 5 1 1 60263
0 60265 7 1 2 60261 60264
0 60266 5 1 1 60265
0 60267 7 1 2 62258 60266
0 60268 5 1 1 60267
0 60269 7 1 2 93205 97764
0 60270 5 1 1 60269
0 60271 7 1 2 92635 99308
0 60272 7 1 2 101339 60271
0 60273 5 1 1 60272
0 60274 7 1 2 60270 60273
0 60275 5 1 1 60274
0 60276 7 1 2 86297 60275
0 60277 5 1 1 60276
0 60278 7 1 2 93144 102246
0 60279 7 1 2 98759 60278
0 60280 5 1 1 60279
0 60281 7 1 2 103048 60280
0 60282 5 1 1 60281
0 60283 7 1 2 103041 60282
0 60284 5 1 1 60283
0 60285 7 1 2 72281 99674
0 60286 7 1 2 97593 60285
0 60287 7 1 2 101823 60286
0 60288 5 1 1 60287
0 60289 7 1 2 83825 78356
0 60290 7 1 2 92636 97596
0 60291 7 1 2 60289 60290
0 60292 5 1 1 60291
0 60293 7 1 2 60288 60292
0 60294 5 1 1 60293
0 60295 7 1 2 64016 60294
0 60296 5 1 1 60295
0 60297 7 2 2 92823 100583
0 60298 7 1 2 90691 96744
0 60299 7 1 2 84925 60298
0 60300 7 1 2 103800 60299
0 60301 5 1 1 60300
0 60302 7 1 2 60296 60301
0 60303 7 1 2 60284 60302
0 60304 5 1 1 60303
0 60305 7 1 2 69651 60304
0 60306 5 1 1 60305
0 60307 7 1 2 60277 60306
0 60308 5 1 1 60307
0 60309 7 1 2 62694 60308
0 60310 5 1 1 60309
0 60311 7 1 2 78903 38169
0 60312 5 1 1 60311
0 60313 7 1 2 87412 60312
0 60314 5 1 1 60313
0 60315 7 1 2 70983 89090
0 60316 5 1 1 60315
0 60317 7 1 2 60314 60316
0 60318 5 2 1 60317
0 60319 7 1 2 103407 103802
0 60320 5 1 1 60319
0 60321 7 1 2 80249 97594
0 60322 7 1 2 99471 60321
0 60323 7 1 2 103679 60322
0 60324 5 1 1 60323
0 60325 7 1 2 60320 60324
0 60326 5 1 1 60325
0 60327 7 1 2 73230 60326
0 60328 5 1 1 60327
0 60329 7 1 2 60310 60328
0 60330 5 1 1 60329
0 60331 7 1 2 82638 80311
0 60332 7 1 2 60330 60331
0 60333 5 1 1 60332
0 60334 7 1 2 60268 60333
0 60335 5 1 1 60334
0 60336 7 1 2 66202 60335
0 60337 5 1 1 60336
0 60338 7 1 2 93539 101627
0 60339 5 1 1 60338
0 60340 7 1 2 65615 84914
0 60341 5 1 1 60340
0 60342 7 1 2 103127 60341
0 60343 5 1 1 60342
0 60344 7 1 2 82344 60343
0 60345 5 1 1 60344
0 60346 7 1 2 60339 60345
0 60347 5 1 1 60346
0 60348 7 1 2 69652 60347
0 60349 5 1 1 60348
0 60350 7 1 2 97393 102532
0 60351 5 1 1 60350
0 60352 7 1 2 60349 60351
0 60353 5 1 1 60352
0 60354 7 1 2 62259 60353
0 60355 5 1 1 60354
0 60356 7 1 2 71401 103803
0 60357 5 1 1 60356
0 60358 7 1 2 73366 92532
0 60359 5 1 1 60358
0 60360 7 1 2 60357 60359
0 60361 5 1 1 60360
0 60362 7 1 2 70799 60361
0 60363 5 1 1 60362
0 60364 7 1 2 72091 87116
0 60365 7 1 2 80673 60364
0 60366 5 1 1 60365
0 60367 7 1 2 60363 60366
0 60368 5 1 1 60367
0 60369 7 1 2 100443 60368
0 60370 5 1 1 60369
0 60371 7 1 2 60355 60370
0 60372 5 1 1 60371
0 60373 7 1 2 97409 97382
0 60374 7 1 2 60372 60373
0 60375 5 1 1 60374
0 60376 7 1 2 60337 60375
0 60377 5 1 1 60376
0 60378 7 1 2 69154 60377
0 60379 5 1 1 60378
0 60380 7 2 2 62991 100942
0 60381 7 1 2 72591 103804
0 60382 5 1 1 60381
0 60383 7 1 2 72592 82345
0 60384 5 1 1 60383
0 60385 7 1 2 81118 60384
0 60386 5 1 1 60385
0 60387 7 1 2 86737 97480
0 60388 7 1 2 60386 60387
0 60389 5 1 1 60388
0 60390 7 1 2 60382 60389
0 60391 5 1 1 60390
0 60392 7 1 2 76745 60391
0 60393 5 1 1 60392
0 60394 7 1 2 82311 100584
0 60395 7 1 2 97561 60394
0 60396 5 1 1 60395
0 60397 7 1 2 60393 60396
0 60398 5 1 1 60397
0 60399 7 1 2 103004 100829
0 60400 7 1 2 60398 60399
0 60401 5 1 1 60400
0 60402 7 1 2 90951 83709
0 60403 7 1 2 95547 60402
0 60404 7 1 2 103669 60403
0 60405 5 1 1 60404
0 60406 7 1 2 72593 92998
0 60407 7 1 2 95169 99620
0 60408 7 1 2 100114 60407
0 60409 7 1 2 60406 60408
0 60410 5 1 1 60409
0 60411 7 1 2 60405 60410
0 60412 5 1 1 60411
0 60413 7 1 2 81108 60412
0 60414 5 1 1 60413
0 60415 7 1 2 320 35730
0 60416 5 1 1 60415
0 60417 7 1 2 92185 60416
0 60418 5 1 1 60417
0 60419 7 1 2 72769 101307
0 60420 5 1 1 60419
0 60421 7 1 2 93611 60420
0 60422 5 1 1 60421
0 60423 7 1 2 60418 60422
0 60424 5 1 1 60423
0 60425 7 1 2 90631 94640
0 60426 7 1 2 100947 60425
0 60427 7 1 2 60424 60426
0 60428 5 1 1 60427
0 60429 7 1 2 60414 60428
0 60430 5 1 1 60429
0 60431 7 1 2 70800 60430
0 60432 5 1 1 60431
0 60433 7 1 2 72594 51845
0 60434 5 1 1 60433
0 60435 7 1 2 74992 97362
0 60436 5 1 1 60435
0 60437 7 1 2 60434 60436
0 60438 5 1 1 60437
0 60439 7 1 2 81109 60438
0 60440 5 1 1 60439
0 60441 7 1 2 86742 92440
0 60442 7 1 2 103805 60441
0 60443 5 1 1 60442
0 60444 7 1 2 60440 60443
0 60445 5 1 1 60444
0 60446 7 1 2 103176 60445
0 60447 5 1 1 60446
0 60448 7 1 2 60432 60447
0 60449 7 1 2 60401 60448
0 60450 5 1 1 60449
0 60451 7 1 2 70547 60450
0 60452 5 1 1 60451
0 60453 7 1 2 81110 97330
0 60454 5 1 1 60453
0 60455 7 1 2 89673 91650
0 60456 7 1 2 93399 60455
0 60457 5 1 1 60456
0 60458 7 1 2 60454 60457
0 60459 5 1 1 60458
0 60460 7 1 2 100075 60459
0 60461 5 1 1 60460
0 60462 7 1 2 79273 98001
0 60463 7 1 2 87944 60462
0 60464 7 1 2 91935 60463
0 60465 5 1 1 60464
0 60466 7 1 2 60461 60465
0 60467 5 1 1 60466
0 60468 7 1 2 72595 60467
0 60469 5 1 1 60468
0 60470 7 1 2 70801 102534
0 60471 5 1 1 60470
0 60472 7 1 2 71550 100076
0 60473 5 1 1 60472
0 60474 7 1 2 60471 60473
0 60475 5 1 1 60474
0 60476 7 1 2 60475 100868
0 60477 5 1 1 60476
0 60478 7 1 2 82708 93157
0 60479 7 1 2 94643 60478
0 60480 5 1 1 60479
0 60481 7 1 2 60477 60480
0 60482 5 1 1 60481
0 60483 7 1 2 72092 60482
0 60484 5 1 1 60483
0 60485 7 1 2 60469 60484
0 60486 5 1 1 60485
0 60487 7 1 2 70548 60486
0 60488 5 1 1 60487
0 60489 7 1 2 1303 92016
0 60490 5 1 1 60489
0 60491 7 1 2 83841 60490
0 60492 5 1 1 60491
0 60493 7 1 2 62260 60492
0 60494 5 2 1 60493
0 60495 7 1 2 93572 100869
0 60496 5 1 1 60495
0 60497 7 1 2 103806 60496
0 60498 5 1 1 60497
0 60499 7 1 2 60498 98571
0 60500 5 1 1 60499
0 60501 7 1 2 60488 60500
0 60502 5 1 1 60501
0 60503 7 1 2 97522 60502
0 60504 5 1 1 60503
0 60505 7 1 2 92103 102708
0 60506 5 1 1 60505
0 60507 7 2 2 80674 90871
0 60508 5 1 1 103808
0 60509 7 1 2 60506 60508
0 60510 5 1 1 60509
0 60511 7 1 2 93612 60510
0 60512 5 1 1 60511
0 60513 7 1 2 87486 103801
0 60514 7 1 2 94043 60513
0 60515 5 1 1 60514
0 60516 7 1 2 60512 60515
0 60517 5 1 1 60516
0 60518 7 1 2 70802 60517
0 60519 5 1 1 60518
0 60520 7 1 2 81111 93236
0 60521 5 1 1 60520
0 60522 7 1 2 103807 60521
0 60523 5 1 1 60522
0 60524 7 1 2 92186 60523
0 60525 5 1 1 60524
0 60526 7 1 2 60519 60525
0 60527 5 1 1 60526
0 60528 7 1 2 103177 60527
0 60529 5 1 1 60528
0 60530 7 1 2 100786 60529
0 60531 5 1 1 60530
0 60532 7 1 2 65616 60531
0 60533 5 1 1 60532
0 60534 7 1 2 60504 60533
0 60535 7 1 2 60452 60534
0 60536 5 1 1 60535
0 60537 7 1 2 79196 60536
0 60538 5 1 1 60537
0 60539 7 1 2 67759 93645
0 60540 5 1 1 60539
0 60541 7 1 2 93620 60540
0 60542 5 1 1 60541
0 60543 7 1 2 103582 60542
0 60544 5 1 1 60543
0 60545 7 1 2 90884 97559
0 60546 7 1 2 99840 60545
0 60547 5 1 1 60546
0 60548 7 1 2 60544 60547
0 60549 5 1 1 60548
0 60550 7 1 2 73140 60549
0 60551 5 1 1 60550
0 60552 7 1 2 70549 36249
0 60553 5 1 1 60552
0 60554 7 1 2 62992 95548
0 60555 7 1 2 79157 60554
0 60556 7 1 2 1722 60555
0 60557 7 1 2 60553 60556
0 60558 5 1 1 60557
0 60559 7 1 2 60551 60558
0 60560 5 1 1 60559
0 60561 7 1 2 90632 60560
0 60562 5 1 1 60561
0 60563 7 2 2 91110 83361
0 60564 5 1 1 103810
0 60565 7 1 2 81216 101716
0 60566 5 1 1 60565
0 60567 7 1 2 60564 60566
0 60568 5 1 1 60567
0 60569 7 1 2 99708 98359
0 60570 7 1 2 60568 60569
0 60571 5 1 1 60570
0 60572 7 1 2 60562 60571
0 60573 5 1 1 60572
0 60574 7 1 2 68051 60573
0 60575 5 1 1 60574
0 60576 7 1 2 78897 70999
0 60577 7 2 2 73141 60576
0 60578 7 1 2 87898 100155
0 60579 7 1 2 103812 60578
0 60580 5 1 1 60579
0 60581 7 1 2 60575 60580
0 60582 5 1 1 60581
0 60583 7 1 2 61338 60582
0 60584 5 1 1 60583
0 60585 7 1 2 78853 80237
0 60586 5 1 1 60585
0 60587 7 1 2 68052 103811
0 60588 5 1 1 60587
0 60589 7 1 2 60586 60588
0 60590 5 1 1 60589
0 60591 7 1 2 103750 60590
0 60592 5 1 1 60591
0 60593 7 1 2 60584 60592
0 60594 5 1 1 60593
0 60595 7 1 2 64238 60594
0 60596 5 1 1 60595
0 60597 7 1 2 75626 96684
0 60598 7 1 2 103813 60597
0 60599 7 1 2 91037 60598
0 60600 5 1 1 60599
0 60601 7 1 2 60596 60600
0 60602 5 1 1 60601
0 60603 7 1 2 64310 82124
0 60604 7 1 2 60602 60603
0 60605 5 1 1 60604
0 60606 7 1 2 60538 60605
0 60607 7 1 2 60379 60606
0 60608 5 1 1 60607
0 60609 7 1 2 73049 60608
0 60610 5 1 1 60609
0 60611 7 1 2 86274 97927
0 60612 5 1 1 60611
0 60613 7 1 2 97388 60612
0 60614 5 1 1 60613
0 60615 7 1 2 86269 97698
0 60616 5 1 1 60615
0 60617 7 1 2 60614 60616
0 60618 5 1 1 60617
0 60619 7 1 2 66066 60618
0 60620 5 1 1 60619
0 60621 7 1 2 86622 100954
0 60622 5 1 1 60621
0 60623 7 1 2 81112 60622
0 60624 5 1 1 60623
0 60625 7 1 2 86623 94574
0 60626 5 1 1 60625
0 60627 7 1 2 82346 60626
0 60628 5 1 1 60627
0 60629 7 1 2 60624 60628
0 60630 5 1 1 60629
0 60631 7 1 2 63862 60630
0 60632 5 1 1 60631
0 60633 7 2 2 71402 77826
0 60634 7 1 2 84518 101768
0 60635 7 1 2 103814 60634
0 60636 5 1 1 60635
0 60637 7 1 2 60632 60636
0 60638 7 1 2 60620 60637
0 60639 5 1 1 60638
0 60640 7 1 2 70550 60639
0 60641 5 1 1 60640
0 60642 7 1 2 81113 97892
0 60643 5 1 1 60642
0 60644 7 1 2 86270 92017
0 60645 5 1 1 60644
0 60646 7 1 2 60643 60645
0 60647 5 1 1 60646
0 60648 7 1 2 73095 60647
0 60649 5 1 1 60648
0 60650 7 1 2 60641 60649
0 60651 5 1 1 60650
0 60652 7 1 2 79197 60651
0 60653 5 1 1 60652
0 60654 7 1 2 84840 86271
0 60655 7 1 2 7632 60654
0 60656 5 1 1 60655
0 60657 7 1 2 65889 101127
0 60658 5 1 1 60657
0 60659 7 1 2 60656 60658
0 60660 5 1 1 60659
0 60661 7 1 2 83362 60660
0 60662 5 1 1 60661
0 60663 7 1 2 72477 94580
0 60664 7 1 2 96152 60663
0 60665 5 1 1 60664
0 60666 7 1 2 60662 60665
0 60667 5 1 1 60666
0 60668 7 1 2 82347 60667
0 60669 5 1 1 60668
0 60670 7 1 2 60653 60669
0 60671 5 1 1 60670
0 60672 7 1 2 98660 60671
0 60673 5 1 1 60672
0 60674 7 1 2 66067 103809
0 60675 5 1 1 60674
0 60676 7 1 2 70984 93319
0 60677 5 1 1 60676
0 60678 7 1 2 60675 60677
0 60679 5 2 1 60678
0 60680 7 1 2 68730 103816
0 60681 5 1 1 60680
0 60682 7 1 2 91209 96059
0 60683 5 1 1 60682
0 60684 7 1 2 60681 60683
0 60685 5 1 1 60684
0 60686 7 1 2 62936 60685
0 60687 5 1 1 60686
0 60688 7 1 2 82348 94581
0 60689 5 1 1 60688
0 60690 7 1 2 60687 60689
0 60691 5 1 1 60690
0 60692 7 1 2 69653 60691
0 60693 5 1 1 60692
0 60694 7 2 2 80943 80827
0 60695 7 1 2 79915 79461
0 60696 7 1 2 103818 60695
0 60697 5 1 1 60696
0 60698 7 1 2 60693 60697
0 60699 5 1 1 60698
0 60700 7 1 2 65617 60699
0 60701 5 1 1 60700
0 60702 7 1 2 71994 72415
0 60703 7 1 2 101169 60702
0 60704 5 1 1 60703
0 60705 7 1 2 60701 60704
0 60706 5 1 1 60705
0 60707 7 1 2 62261 60706
0 60708 5 1 1 60707
0 60709 7 1 2 86937 86635
0 60710 7 1 2 103817 60709
0 60711 5 1 1 60710
0 60712 7 1 2 60708 60711
0 60713 5 1 1 60712
0 60714 7 1 2 64239 60713
0 60715 5 1 1 60714
0 60716 7 1 2 86069 91684
0 60717 5 1 1 60716
0 60718 7 1 2 60717 97948
0 60719 5 1 1 60718
0 60720 7 1 2 80118 91773
0 60721 7 1 2 60719 60720
0 60722 5 1 1 60721
0 60723 7 1 2 60715 60722
0 60724 5 1 1 60723
0 60725 7 1 2 65890 60724
0 60726 5 1 1 60725
0 60727 7 1 2 79721 93386
0 60728 7 1 2 100919 60727
0 60729 5 1 1 60728
0 60730 7 1 2 60726 60729
0 60731 5 1 1 60730
0 60732 7 1 2 78854 60731
0 60733 5 1 1 60732
0 60734 7 1 2 81013 86520
0 60735 7 1 2 101879 60734
0 60736 5 1 1 60735
0 60737 7 1 2 74134 81114
0 60738 5 1 1 60737
0 60739 7 1 2 37299 60738
0 60740 5 1 1 60739
0 60741 7 1 2 77605 103571
0 60742 7 1 2 60740 60741
0 60743 5 1 1 60742
0 60744 7 1 2 60736 60743
0 60745 5 1 1 60744
0 60746 7 1 2 61939 60745
0 60747 5 1 1 60746
0 60748 7 1 2 80830 87118
0 60749 7 2 2 69875 73858
0 60750 7 1 2 93427 103820
0 60751 7 1 2 60748 60750
0 60752 5 1 1 60751
0 60753 7 1 2 60747 60752
0 60754 5 1 1 60753
0 60755 7 1 2 64818 60754
0 60756 5 1 1 60755
0 60757 7 1 2 76592 89819
0 60758 5 1 1 60757
0 60759 7 1 2 90395 80735
0 60760 7 1 2 103821 60759
0 60761 5 1 1 60760
0 60762 7 1 2 60758 60761
0 60763 5 1 1 60762
0 60764 7 1 2 79383 76680
0 60765 7 1 2 60763 60764
0 60766 5 1 1 60765
0 60767 7 1 2 60756 60766
0 60768 5 1 1 60767
0 60769 7 1 2 62459 60768
0 60770 5 1 1 60769
0 60771 7 1 2 78523 80119
0 60772 7 1 2 90756 60771
0 60773 7 1 2 95248 60772
0 60774 5 1 1 60773
0 60775 7 1 2 60770 60774
0 60776 5 1 1 60775
0 60777 7 1 2 62262 60776
0 60778 5 1 1 60777
0 60779 7 1 2 88343 76625
0 60780 5 1 1 60779
0 60781 7 1 2 62263 86178
0 60782 7 1 2 83851 60781
0 60783 5 1 1 60782
0 60784 7 1 2 60780 60783
0 60785 5 1 1 60784
0 60786 7 1 2 72596 60785
0 60787 5 1 1 60786
0 60788 7 1 2 78031 90248
0 60789 7 1 2 73692 60788
0 60790 7 1 2 93259 60789
0 60791 5 1 1 60790
0 60792 7 1 2 60787 60791
0 60793 5 1 1 60792
0 60794 7 1 2 70551 60793
0 60795 5 1 1 60794
0 60796 7 1 2 75518 87676
0 60797 7 1 2 89557 60796
0 60798 7 1 2 89896 60797
0 60799 5 1 1 60798
0 60800 7 1 2 60795 60799
0 60801 5 1 1 60800
0 60802 7 1 2 79198 60801
0 60803 5 1 1 60802
0 60804 7 1 2 86636 88058
0 60805 7 1 2 92923 60804
0 60806 7 1 2 76753 60805
0 60807 5 1 1 60806
0 60808 7 1 2 60803 60807
0 60809 7 1 2 60778 60808
0 60810 5 1 1 60809
0 60811 7 1 2 70803 60810
0 60812 5 1 1 60811
0 60813 7 1 2 90551 103815
0 60814 5 1 1 60813
0 60815 7 1 2 92383 103819
0 60816 5 1 1 60815
0 60817 7 1 2 60814 60816
0 60818 5 1 1 60817
0 60819 7 1 2 86037 75310
0 60820 7 1 2 85863 60819
0 60821 7 1 2 60818 60820
0 60822 5 1 1 60821
0 60823 7 1 2 60812 60822
0 60824 7 1 2 60733 60823
0 60825 5 1 1 60824
0 60826 7 1 2 98674 60825
0 60827 5 1 1 60826
0 60828 7 1 2 60673 60827
0 60829 5 1 1 60828
0 60830 7 1 2 64424 60829
0 60831 5 1 1 60830
0 60832 7 1 2 79722 73231
0 60833 5 2 1 60832
0 60834 7 1 2 62264 101341
0 60835 5 1 1 60834
0 60836 7 1 2 103822 60835
0 60837 5 1 1 60836
0 60838 7 1 2 81115 97799
0 60839 7 1 2 60837 60838
0 60840 5 1 1 60839
0 60841 7 1 2 79723 78763
0 60842 7 1 2 97227 60841
0 60843 5 1 1 60842
0 60844 7 1 2 75972 73702
0 60845 7 1 2 73746 60844
0 60846 7 1 2 80378 60845
0 60847 5 1 1 60846
0 60848 7 1 2 60843 60847
0 60849 5 1 1 60848
0 60850 7 1 2 71609 60849
0 60851 5 1 1 60850
0 60852 7 1 2 62265 91443
0 60853 5 1 1 60852
0 60854 7 1 2 62266 94149
0 60855 5 1 1 60854
0 60856 7 1 2 67098 94294
0 60857 5 1 1 60856
0 60858 7 1 2 72093 60857
0 60859 7 1 2 60855 60858
0 60860 5 1 1 60859
0 60861 7 1 2 62267 94202
0 60862 5 1 1 60861
0 60863 7 1 2 72217 103823
0 60864 7 1 2 60862 60863
0 60865 5 1 1 60864
0 60866 7 1 2 60860 60865
0 60867 5 1 1 60866
0 60868 7 1 2 60853 60867
0 60869 5 1 1 60868
0 60870 7 1 2 79199 60869
0 60871 5 1 1 60870
0 60872 7 1 2 9943 75635
0 60873 5 1 1 60872
0 60874 7 1 2 80502 77158
0 60875 7 1 2 81075 60874
0 60876 7 1 2 60873 60875
0 60877 5 1 1 60876
0 60878 7 1 2 60871 60877
0 60879 5 1 1 60878
0 60880 7 1 2 68053 60879
0 60881 5 1 1 60880
0 60882 7 1 2 60851 60881
0 60883 5 1 1 60882
0 60884 7 1 2 82125 91038
0 60885 7 1 2 60883 60884
0 60886 5 1 1 60885
0 60887 7 1 2 60840 60886
0 60888 5 1 1 60887
0 60889 7 1 2 93923 60888
0 60890 5 1 1 60889
0 60891 7 1 2 66336 69654
0 60892 7 1 2 75535 60891
0 60893 7 1 2 92310 60892
0 60894 7 1 2 97942 101261
0 60895 7 1 2 60893 60894
0 60896 5 1 1 60895
0 60897 7 1 2 73591 97687
0 60898 5 1 1 60897
0 60899 7 1 2 66337 72094
0 60900 7 1 2 79506 60899
0 60901 7 1 2 103659 60900
0 60902 5 1 1 60901
0 60903 7 1 2 60898 60902
0 60904 5 1 1 60903
0 60905 7 1 2 89430 88132
0 60906 7 1 2 60904 60905
0 60907 5 1 1 60906
0 60908 7 1 2 60896 60907
0 60909 5 1 1 60908
0 60910 7 1 2 66203 60909
0 60911 5 1 1 60910
0 60912 7 1 2 73592 84428
0 60913 7 1 2 94641 60912
0 60914 7 1 2 80515 60913
0 60915 7 1 2 90736 60914
0 60916 5 1 1 60915
0 60917 7 1 2 60911 60916
0 60918 5 1 1 60917
0 60919 7 1 2 69275 60918
0 60920 5 1 1 60919
0 60921 7 1 2 65618 97472
0 60922 5 1 1 60921
0 60923 7 1 2 70552 29663
0 60924 5 1 1 60923
0 60925 7 1 2 84240 60924
0 60926 7 1 2 60922 60925
0 60927 5 1 1 60926
0 60928 7 1 2 84236 86420
0 60929 5 1 1 60928
0 60930 7 1 2 60929 97494
0 60931 5 1 1 60930
0 60932 7 1 2 92678 60931
0 60933 5 1 1 60932
0 60934 7 2 2 66204 98093
0 60935 7 1 2 100138 103824
0 60936 7 1 2 103629 60935
0 60937 5 1 1 60936
0 60938 7 1 2 60933 60937
0 60939 7 1 2 60927 60938
0 60940 5 1 1 60939
0 60941 7 1 2 66068 60940
0 60942 5 1 1 60941
0 60943 7 1 2 72485 93011
0 60944 7 1 2 96078 103825
0 60945 7 1 2 60943 60944
0 60946 5 1 1 60945
0 60947 7 1 2 69459 83770
0 60948 7 1 2 96921 60947
0 60949 7 1 2 103729 60948
0 60950 5 1 1 60949
0 60951 7 1 2 60946 60950
0 60952 7 1 2 60942 60951
0 60953 5 1 1 60952
0 60954 7 1 2 69155 60953
0 60955 5 1 1 60954
0 60956 7 2 2 78855 95567
0 60957 7 1 2 101265 103826
0 60958 5 1 1 60957
0 60959 7 1 2 60955 60958
0 60960 5 1 1 60959
0 60961 7 1 2 69083 60960
0 60962 5 1 1 60961
0 60963 7 1 2 60920 60962
0 60964 5 1 1 60963
0 60965 7 1 2 62268 60964
0 60966 5 1 1 60965
0 60967 7 1 2 71403 87762
0 60968 5 1 1 60967
0 60969 7 1 2 64017 98865
0 60970 5 1 1 60969
0 60971 7 1 2 60968 60970
0 60972 5 1 1 60971
0 60973 7 1 2 98030 60972
0 60974 5 1 1 60973
0 60975 7 1 2 33028 60974
0 60976 5 1 1 60975
0 60977 7 1 2 67099 60976
0 60978 5 1 1 60977
0 60979 7 1 2 65891 93924
0 60980 7 1 2 99236 60979
0 60981 5 1 1 60980
0 60982 7 1 2 60978 60981
0 60983 5 1 1 60982
0 60984 7 1 2 70553 60983
0 60985 5 1 1 60984
0 60986 7 1 2 99835 99932
0 60987 5 1 1 60986
0 60988 7 1 2 60985 60987
0 60989 5 1 1 60988
0 60990 7 1 2 74993 60989
0 60991 5 1 1 60990
0 60992 7 1 2 71404 100038
0 60993 5 1 1 60992
0 60994 7 1 2 97755 101479
0 60995 5 1 1 60994
0 60996 7 1 2 60993 60995
0 60997 5 1 1 60996
0 60998 7 1 2 70554 60997
0 60999 5 1 1 60998
0 61000 7 1 2 76616 93925
0 61001 7 1 2 98850 61000
0 61002 5 1 1 61001
0 61003 7 1 2 60999 61002
0 61004 5 1 1 61003
0 61005 7 1 2 74994 61004
0 61006 5 1 1 61005
0 61007 7 1 2 86385 97623
0 61008 7 1 2 72309 61007
0 61009 5 1 1 61008
0 61010 7 1 2 61006 61009
0 61011 5 1 1 61010
0 61012 7 1 2 90737 61011
0 61013 5 1 1 61012
0 61014 7 1 2 70555 95295
0 61015 7 1 2 103367 61014
0 61016 7 1 2 99933 61015
0 61017 5 1 1 61016
0 61018 7 1 2 61013 61017
0 61019 7 1 2 60991 61018
0 61020 5 1 1 61019
0 61021 7 1 2 83906 61020
0 61022 5 1 1 61021
0 61023 7 1 2 97027 99040
0 61024 7 1 2 101392 61023
0 61025 7 1 2 103434 61024
0 61026 5 1 1 61025
0 61027 7 1 2 61022 61026
0 61028 7 1 2 60966 61027
0 61029 5 1 1 61028
0 61030 7 1 2 73050 61029
0 61031 5 1 1 61030
0 61032 7 1 2 84241 100033
0 61033 7 1 2 93535 61032
0 61034 5 1 1 61033
0 61035 7 1 2 88903 74252
0 61036 7 1 2 96924 61035
0 61037 7 1 2 98661 61036
0 61038 5 1 1 61037
0 61039 7 1 2 61034 61038
0 61040 5 1 1 61039
0 61041 7 1 2 85254 61040
0 61042 5 1 1 61041
0 61043 7 1 2 77001 73747
0 61044 7 1 2 95430 61043
0 61045 7 1 2 97229 61044
0 61046 7 1 2 93529 61045
0 61047 5 1 1 61046
0 61048 7 1 2 61042 61047
0 61049 5 1 1 61048
0 61050 7 1 2 68731 61049
0 61051 5 1 1 61050
0 61052 7 1 2 86619 84308
0 61053 5 1 1 61052
0 61054 7 1 2 83468 82892
0 61055 5 1 1 61054
0 61056 7 1 2 61053 61055
0 61057 5 1 1 61056
0 61058 7 1 2 83907 61057
0 61059 5 1 1 61058
0 61060 7 2 2 84061 97230
0 61061 7 1 2 71274 74163
0 61062 7 1 2 103828 61061
0 61063 5 1 1 61062
0 61064 7 1 2 61059 61063
0 61065 5 1 1 61064
0 61066 7 1 2 92496 98184
0 61067 7 1 2 61065 61066
0 61068 5 1 1 61067
0 61069 7 1 2 61051 61068
0 61070 5 1 1 61069
0 61071 7 1 2 70804 61070
0 61072 5 1 1 61071
0 61073 7 1 2 76437 84579
0 61074 7 1 2 103829 61073
0 61075 5 1 1 61074
0 61076 7 1 2 84339 93378
0 61077 5 1 1 61076
0 61078 7 1 2 6486 61077
0 61079 5 1 1 61078
0 61080 7 1 2 79801 97960
0 61081 7 1 2 61079 61080
0 61082 5 1 1 61081
0 61083 7 1 2 61075 61082
0 61084 5 1 1 61083
0 61085 7 1 2 62269 98675
0 61086 7 1 2 61084 61085
0 61087 5 1 1 61086
0 61088 7 1 2 65619 61087
0 61089 7 1 2 61072 61088
0 61090 5 1 1 61089
0 61091 7 2 2 79384 103705
0 61092 7 1 2 88282 103830
0 61093 5 1 1 61092
0 61094 7 1 2 68732 79647
0 61095 7 1 2 100844 98717
0 61096 7 1 2 61094 61095
0 61097 5 1 1 61096
0 61098 7 1 2 61093 61097
0 61099 5 1 1 61098
0 61100 7 1 2 61339 61099
0 61101 5 1 1 61100
0 61102 7 1 2 73816 99815
0 61103 7 1 2 98213 61102
0 61104 7 1 2 90738 61103
0 61105 5 1 1 61104
0 61106 7 1 2 61101 61105
0 61107 5 1 1 61106
0 61108 7 1 2 67317 61107
0 61109 5 1 1 61108
0 61110 7 1 2 61340 90821
0 61111 7 1 2 103721 99455
0 61112 7 1 2 61110 61111
0 61113 5 1 1 61112
0 61114 7 1 2 61109 61113
0 61115 5 1 1 61114
0 61116 7 1 2 71183 61115
0 61117 5 1 1 61116
0 61118 7 2 2 99041 103831
0 61119 7 1 2 71275 75228
0 61120 7 1 2 103832 61119
0 61121 5 1 1 61120
0 61122 7 1 2 65892 61121
0 61123 7 1 2 61117 61122
0 61124 5 1 1 61123
0 61125 7 1 2 83927 89795
0 61126 5 1 1 61125
0 61127 7 1 2 63863 97931
0 61128 5 1 1 61127
0 61129 7 1 2 61126 61128
0 61130 5 1 1 61129
0 61131 7 1 2 74995 61130
0 61132 5 1 1 61131
0 61133 7 1 2 72597 83635
0 61134 7 1 2 97958 61133
0 61135 5 1 1 61134
0 61136 7 1 2 61132 61135
0 61137 5 1 1 61136
0 61138 7 1 2 103684 61137
0 61139 5 1 1 61138
0 61140 7 1 2 83928 97963
0 61141 5 1 1 61140
0 61142 7 1 2 83914 94325
0 61143 5 1 1 61142
0 61144 7 1 2 61141 61143
0 61145 5 1 1 61144
0 61146 7 1 2 72598 99695
0 61147 7 1 2 97688 61146
0 61148 7 1 2 61145 61147
0 61149 5 1 1 61148
0 61150 7 1 2 70805 61149
0 61151 7 1 2 61139 61150
0 61152 5 1 1 61151
0 61153 7 1 2 61124 61152
0 61154 5 1 1 61153
0 61155 7 1 2 83929 98665
0 61156 5 1 1 61155
0 61157 7 1 2 70556 61156
0 61158 7 1 2 61154 61157
0 61159 5 1 1 61158
0 61160 7 1 2 61090 61159
0 61161 5 1 1 61160
0 61162 7 1 2 74484 97285
0 61163 5 1 1 61162
0 61164 7 1 2 103833 61163
0 61165 5 1 1 61164
0 61166 7 1 2 66798 92452
0 61167 5 1 1 61166
0 61168 7 1 2 29501 61167
0 61169 5 1 1 61168
0 61170 7 1 2 71276 73748
0 61171 7 1 2 98214 61170
0 61172 7 1 2 91734 61171
0 61173 7 1 2 61169 61172
0 61174 5 1 1 61173
0 61175 7 1 2 61165 61174
0 61176 5 1 1 61175
0 61177 7 1 2 70557 61176
0 61178 5 1 1 61177
0 61179 7 1 2 88415 92588
0 61180 7 1 2 98215 61179
0 61181 7 1 2 103183 61180
0 61182 5 1 1 61181
0 61183 7 1 2 61178 61182
0 61184 5 1 1 61183
0 61185 7 1 2 71995 61184
0 61186 5 1 1 61185
0 61187 7 1 2 83620 97282
0 61188 5 1 1 61187
0 61189 7 1 2 79870 76626
0 61190 7 1 2 85946 61189
0 61191 5 1 1 61190
0 61192 7 1 2 61188 61191
0 61193 5 1 1 61192
0 61194 7 1 2 83908 98676
0 61195 7 1 2 61193 61194
0 61196 5 1 1 61195
0 61197 7 1 2 61186 61196
0 61198 7 1 2 61161 61197
0 61199 5 1 1 61198
0 61200 7 1 2 64425 61199
0 61201 5 1 1 61200
0 61202 7 1 2 74475 95478
0 61203 5 1 1 61202
0 61204 7 1 2 71184 86637
0 61205 5 1 1 61204
0 61206 7 1 2 61203 61205
0 61207 5 1 1 61206
0 61208 7 1 2 71610 61207
0 61209 5 1 1 61208
0 61210 7 1 2 6261 75006
0 61211 5 1 1 61210
0 61212 7 1 2 73232 61211
0 61213 5 1 1 61212
0 61214 7 1 2 62937 76835
0 61215 7 1 2 100396 61214
0 61216 5 1 1 61215
0 61217 7 1 2 67100 61216
0 61218 7 1 2 61213 61217
0 61219 5 1 1 61218
0 61220 7 1 2 73269 89728
0 61221 5 1 1 61220
0 61222 7 1 2 62270 61221
0 61223 7 1 2 97864 61222
0 61224 5 1 1 61223
0 61225 7 1 2 61219 61224
0 61226 5 1 1 61225
0 61227 7 1 2 61209 61226
0 61228 5 1 1 61227
0 61229 7 1 2 91039 103827
0 61230 7 1 2 61228 61229
0 61231 5 1 1 61230
0 61232 7 1 2 61201 61231
0 61233 7 1 2 61031 61232
0 61234 5 1 1 61233
0 61235 7 1 2 76200 61234
0 61236 5 1 1 61235
0 61237 7 1 2 60890 61236
0 61238 7 1 2 60831 61237
0 61239 7 1 2 60610 61238
0 61240 5 1 1 61239
0 61241 7 1 2 94880 61240
0 61242 5 1 1 61241
0 61243 7 1 2 60259 61242
0 61244 7 1 2 58230 61243
0 61245 7 1 2 48226 61244
0 61246 7 1 2 46300 61245
0 61247 7 1 2 42201 61246
0 61248 7 1 2 29347 61247
0 61249 7 1 2 18439 61248
0 61250 7 1 2 14226 61249
3 129999 5 0 1 61250
