1 0 0 2 0
2 16 1 0
2 17 1 0
1 1 0 2 0
2 18 1 1
2 19 1 1
1 2 0 2 0
2 20 1 2
2 21 1 2
1 3 0 2 0
2 22 1 3
2 23 1 3
1 4 0 2 0
2 24 1 4
2 25 1 4
1 5 0 2 0
2 46 1 5
2 58 1 5
1 6 0 2 0
2 74 1 6
2 90 1 6
1 7 0 2 0
2 106 1 7
2 122 1 7
1 8 0 2 0
2 138 1 8
2 154 1 8
1 9 0 2 0
2 157 1 9
2 158 1 9
1 10 0 2 0
2 159 1 10
2 160 1 10
1 11 0 2 0
2 161 1 11
2 162 1 11
1 12 0 2 0
2 163 1 12
2 164 1 12
1 13 0 2 0
2 165 1 13
2 166 1 13
1 14 0 2 0
2 167 1 14
2 168 1 14
1 15 0 2 0
2 169 1 15
2 170 1 15
2 171 1 42
2 172 1 42
2 173 1 43
2 174 1 43
2 175 1 43
2 176 1 48
2 177 1 48
2 178 1 50
2 179 1 50
2 180 1 51
2 181 1 51
2 182 1 60
2 183 1 60
2 184 1 62
2 185 1 62
2 186 1 63
2 187 1 63
2 188 1 67
2 189 1 67
2 190 1 68
2 191 1 68
2 192 1 76
2 193 1 76
2 194 1 78
2 195 1 78
2 196 1 79
2 197 1 79
2 198 1 83
2 199 1 83
2 200 1 84
2 201 1 84
2 202 1 92
2 203 1 92
2 204 1 94
2 205 1 94
2 206 1 95
2 207 1 95
2 208 1 99
2 209 1 99
2 210 1 100
2 211 1 100
2 212 1 108
2 213 1 108
2 214 1 110
2 215 1 110
2 216 1 111
2 217 1 111
2 218 1 115
2 219 1 115
2 220 1 116
2 221 1 116
2 222 1 124
2 223 1 124
2 224 1 126
2 225 1 126
2 226 1 127
2 227 1 127
2 228 1 131
2 229 1 131
2 230 1 132
2 231 1 132
2 232 1 140
2 233 1 140
2 234 1 142
2 235 1 142
2 236 1 143
2 237 1 143
2 238 1 147
2 239 1 147
2 240 1 148
2 241 1 148
0 26 5 1 1 16
0 27 5 1 1 18
0 28 5 1 1 20
0 29 5 1 1 22
0 30 5 1 1 24
0 31 5 1 1 46
0 32 5 1 1 74
0 33 5 1 1 106
0 34 5 1 1 138
0 35 5 1 1 157
0 36 5 1 1 159
0 37 5 1 1 161
0 38 5 1 1 163
0 39 5 1 1 165
0 40 5 1 1 167
0 41 5 1 1 169
0 42 7 2 2 17 154
0 43 5 3 1 171
0 44 7 1 2 26 34
0 45 5 1 1 44
3 291 7 0 2 173 45
0 47 7 1 2 27 35
0 48 5 2 1 47
0 49 7 1 2 19 158
0 50 5 2 1 49
0 51 7 2 2 176 178
0 52 5 1 1 180
0 53 7 1 2 172 52
0 54 5 1 1 53
0 55 7 1 2 174 181
0 56 5 1 1 55
0 57 7 1 2 54 56
3 292 5 0 1 57
0 59 7 1 2 28 36
0 60 5 2 1 59
0 61 7 1 2 21 160
0 62 5 2 1 61
0 63 7 2 2 182 184
0 64 5 1 1 186
0 65 7 1 2 175 179
0 66 5 1 1 65
0 67 7 2 2 177 66
0 68 5 2 1 188
0 69 7 1 2 64 189
0 70 5 1 1 69
0 71 7 1 2 187 190
0 72 5 1 1 71
0 73 7 1 2 70 72
3 293 5 0 1 73
0 75 7 1 2 29 37
0 76 5 2 1 75
0 77 7 1 2 23 162
0 78 5 2 1 77
0 79 7 2 2 192 194
0 80 5 1 1 196
0 81 7 1 2 185 191
0 82 5 1 1 81
0 83 7 2 2 183 82
0 84 5 2 1 198
0 85 7 1 2 80 199
0 86 5 1 1 85
0 87 7 1 2 197 200
0 88 5 1 1 87
0 89 7 1 2 86 88
3 294 5 0 1 89
0 91 7 1 2 30 38
0 92 5 2 1 91
0 93 7 1 2 25 164
0 94 5 2 1 93
0 95 7 2 2 202 204
0 96 5 1 1 206
0 97 7 1 2 195 201
0 98 5 1 1 97
0 99 7 2 2 193 98
0 100 5 2 1 208
0 101 7 1 2 96 209
0 102 5 1 1 101
0 103 7 1 2 207 210
0 104 5 1 1 103
0 105 7 1 2 102 104
3 295 5 0 1 105
0 107 7 1 2 31 39
0 108 5 2 1 107
0 109 7 1 2 58 166
0 110 5 2 1 109
0 111 7 2 2 212 214
0 112 5 1 1 216
0 113 7 1 2 205 211
0 114 5 1 1 113
0 115 7 2 2 203 114
0 116 5 2 1 218
0 117 7 1 2 112 219
0 118 5 1 1 117
0 119 7 1 2 217 220
0 120 5 1 1 119
0 121 7 1 2 118 120
3 296 5 0 1 121
0 123 7 1 2 32 40
0 124 5 2 1 123
0 125 7 1 2 90 168
0 126 5 2 1 125
0 127 7 2 2 222 224
0 128 5 1 1 226
0 129 7 1 2 215 221
0 130 5 1 1 129
0 131 7 2 2 213 130
0 132 5 2 1 228
0 133 7 1 2 128 229
0 134 5 1 1 133
0 135 7 1 2 227 230
0 136 5 1 1 135
0 137 7 1 2 134 136
3 297 5 0 1 137
0 139 7 1 2 122 170
0 140 5 2 1 139
0 141 7 1 2 33 41
0 142 5 2 1 141
0 143 7 2 2 232 234
0 144 5 1 1 236
0 145 7 1 2 225 231
0 146 5 1 1 145
0 147 7 2 2 223 146
0 148 5 2 1 238
0 149 7 1 2 237 240
0 150 5 1 1 149
0 151 7 1 2 144 239
0 152 5 1 1 151
0 153 7 1 2 150 152
3 298 5 0 1 153
0 155 7 1 2 233 241
0 156 5 1 1 155
3 299 7 0 2 235 156
