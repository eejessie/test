1 0 0 1 0
1 1 0 2 0
2 14 1 1
2 15 1 1
1 2 0 3 0
2 125 1 2
2 126 1 2
2 127 1 2
1 3 0 4 0
2 128 1 3
2 129 1 3
2 130 1 3
2 131 1 3
1 4 0 2 0
2 132 1 4
2 133 1 4
1 5 0 2 0
2 134 1 5
2 135 1 5
1 6 0 2 0
2 136 1 6
2 137 1 6
1 7 0 2 0
2 138 1 7
2 139 1 7
1 8 0 2 0
2 140 1 8
2 141 1 8
1 9 0 0 0
1 10 0 0 0
1 11 0 2 0
2 142 1 11
2 143 1 11
1 12 0 2 0
2 144 1 12
2 145 1 12
1 13 0 3 0
2 146 1 13
2 147 1 13
2 148 1 13
2 149 1 18
2 150 1 18
2 151 1 18
2 152 1 19
2 153 1 19
2 154 1 19
2 155 1 27
2 156 1 27
2 157 1 37
2 158 1 37
2 159 1 37
2 160 1 39
2 161 1 39
2 162 1 43
2 163 1 43
2 164 1 48
2 165 1 48
2 166 1 48
2 167 1 51
2 168 1 51
2 169 1 51
2 170 1 52
2 171 1 52
2 172 1 57
2 173 1 57
2 174 1 58
2 175 1 58
2 176 1 59
2 177 1 59
2 178 1 59
2 179 1 65
2 180 1 65
2 181 1 70
2 182 1 70
2 183 1 72
2 184 1 72
2 185 1 72
2 186 1 72
2 187 1 73
2 188 1 73
2 189 1 86
2 190 1 86
2 191 1 87
2 192 1 87
2 193 1 88
2 194 1 88
2 195 1 92
2 196 1 92
0 16 5 1 1 0
0 17 5 1 1 14
0 18 5 3 1 125
0 19 5 3 1 128
0 20 5 1 1 132
0 21 5 1 1 134
0 22 5 1 1 136
0 23 5 1 1 138
0 24 5 1 1 140
0 25 5 1 1 142
0 26 5 1 1 144
0 27 5 2 1 146
0 28 7 1 2 133 141
0 29 5 1 1 28
0 30 7 1 2 16 29
0 31 5 1 1 30
0 32 7 1 2 20 24
0 33 5 1 1 32
0 34 7 1 2 17 21
0 35 5 1 1 34
0 36 7 1 2 33 35
0 37 7 3 2 31 36
0 38 5 1 1 157
0 39 7 2 2 139 26
0 40 5 1 1 160
0 41 7 1 2 147 161
0 42 5 1 1 41
0 43 7 2 2 23 145
0 44 5 1 1 162
0 45 7 1 2 155 163
0 46 5 1 1 45
0 47 7 1 2 42 46
0 48 5 3 1 47
0 49 7 1 2 129 164
0 50 5 1 1 49
0 51 7 3 2 40 44
0 52 7 2 2 152 156
0 53 5 1 1 170
0 54 7 1 2 167 171
0 55 5 1 1 54
0 56 7 1 2 50 55
0 57 5 2 1 56
0 58 7 2 2 22 143
0 59 5 3 1 174
0 60 7 1 2 149 175
0 61 7 1 2 172 60
0 62 5 1 1 61
0 63 7 1 2 153 165
0 64 5 1 1 63
0 65 7 2 2 130 148
0 66 5 1 1 179
0 67 7 1 2 168 180
0 68 5 1 1 67
0 69 7 1 2 64 68
0 70 5 2 1 69
0 71 7 1 2 137 25
0 72 5 4 1 71
0 73 7 2 2 183 176
0 74 5 1 1 187
0 75 7 1 2 126 74
0 76 5 1 1 75
0 77 7 1 2 150 184
0 78 5 1 1 77
0 79 7 1 2 76 78
0 80 7 1 2 181 79
0 81 5 1 1 80
0 82 7 1 2 62 81
0 83 5 1 1 82
0 84 7 1 2 158 83
0 85 5 1 1 84
0 86 7 2 2 15 135
0 87 5 2 1 189
0 88 7 2 2 127 190
0 89 5 1 1 193
0 90 7 1 2 182 194
0 91 5 1 1 90
0 92 7 2 2 151 191
0 93 5 1 1 195
0 94 7 1 2 196 38
0 95 7 1 2 173 94
0 96 5 1 1 95
0 97 7 1 2 91 96
0 98 5 1 1 97
0 99 7 1 2 188 98
0 100 5 1 1 99
0 101 7 1 2 177 66
0 102 5 1 1 101
0 103 7 1 2 185 53
0 104 5 1 1 103
0 105 7 1 2 169 104
0 106 7 1 2 102 105
0 107 5 1 1 106
0 108 7 1 2 154 186
0 109 5 1 1 108
0 110 7 1 2 131 178
0 111 5 1 1 110
0 112 7 1 2 109 111
0 113 7 1 2 166 112
0 114 5 1 1 113
0 115 7 1 2 107 114
0 116 5 1 1 115
0 117 7 1 2 192 159
0 118 5 1 1 117
0 119 7 1 2 89 93
0 120 7 1 2 118 119
0 121 7 1 2 116 120
0 122 5 1 1 121
0 123 7 1 2 100 122
0 124 7 1 2 85 123
3 699 5 0 1 124
