1 0 0 2 0
2 49 1 0
2 744 1 0
1 1 0 2 0
2 745 1 1
2 746 1 1
1 2 0 2 0
2 747 1 2
2 748 1 2
1 3 0 2 0
2 749 1 3
2 750 1 3
1 4 0 2 0
2 751 1 4
2 752 1 4
1 5 0 2 0
2 753 1 5
2 754 1 5
1 6 0 2 0
2 755 1 6
2 756 1 6
1 7 0 2 0
2 757 1 7
2 758 1 7
1 8 0 2 0
2 759 1 8
2 760 1 8
1 9 0 2 0
2 761 1 9
2 762 1 9
1 10 0 2 0
2 763 1 10
2 764 1 10
1 11 0 2 0
2 765 1 11
2 766 1 11
1 12 0 2 0
2 767 1 12
2 768 1 12
1 13 0 2 0
2 769 1 13
2 770 1 13
1 14 0 2 0
2 771 1 14
2 772 1 14
1 15 0 2 0
2 773 1 15
2 774 1 15
1 16 0 2 0
2 775 1 16
2 776 1 16
1 17 0 2 0
2 777 1 17
2 778 1 17
1 18 0 2 0
2 779 1 18
2 780 1 18
1 19 0 2 0
2 781 1 19
2 782 1 19
1 20 0 2 0
2 783 1 20
2 784 1 20
1 21 0 2 0
2 785 1 21
2 786 1 21
1 22 0 2 0
2 787 1 22
2 788 1 22
1 23 0 2 0
2 789 1 23
2 790 1 23
1 24 0 2 0
2 791 1 24
2 792 1 24
1 25 0 2 0
2 793 1 25
2 794 1 25
1 26 0 2 0
2 795 1 26
2 796 1 26
1 27 0 2 0
2 797 1 27
2 798 1 27
1 28 0 2 0
2 799 1 28
2 800 1 28
1 29 0 2 0
2 801 1 29
2 802 1 29
1 30 0 2 0
2 803 1 30
2 804 1 30
1 31 0 2 0
2 805 1 31
2 806 1 31
1 32 0 2 0
2 807 1 32
2 808 1 32
1 33 0 2 0
2 809 1 33
2 810 1 33
1 34 0 2 0
2 811 1 34
2 812 1 34
1 35 0 2 0
2 813 1 35
2 814 1 35
1 36 0 2 0
2 815 1 36
2 816 1 36
1 37 0 2 0
2 817 1 37
2 818 1 37
1 38 0 2 0
2 819 1 38
2 820 1 38
1 39 0 2 0
2 821 1 39
2 822 1 39
1 40 0 2 0
2 823 1 40
2 824 1 40
1 41 0 2 0
2 825 1 41
2 826 1 41
1 42 0 2 0
2 827 1 42
2 828 1 42
1 43 0 2 0
2 829 1 43
2 830 1 43
1 44 0 2 0
2 831 1 44
2 832 1 44
1 45 0 2 0
2 833 1 45
2 834 1 45
1 46 0 2 0
2 835 1 46
2 836 1 46
1 47 0 2 0
2 837 1 47
2 838 1 47
1 48 0 2 0
2 839 1 48
2 840 1 48
2 841 1 69
2 842 1 69
2 843 1 70
2 844 1 70
2 845 1 71
2 846 1 71
2 847 1 72
2 848 1 72
2 849 1 73
2 850 1 73
2 851 1 74
2 852 1 74
2 853 1 75
2 854 1 75
2 855 1 76
2 856 1 76
2 857 1 77
2 858 1 77
2 859 1 78
2 860 1 78
2 861 1 79
2 862 1 79
2 863 1 80
2 864 1 80
2 865 1 81
2 866 1 81
2 867 1 100
2 868 1 100
2 869 1 102
2 870 1 102
2 871 1 104
2 872 1 104
2 873 1 106
2 874 1 106
2 875 1 107
2 876 1 107
2 877 1 108
2 878 1 108
2 879 1 108
2 880 1 111
2 881 1 111
2 882 1 112
2 883 1 112
2 884 1 115
2 885 1 115
2 886 1 118
2 887 1 118
2 888 1 120
2 889 1 120
2 890 1 123
2 891 1 123
2 892 1 126
2 893 1 126
2 894 1 128
2 895 1 128
2 896 1 131
2 897 1 131
2 898 1 134
2 899 1 134
2 900 1 136
2 901 1 136
2 902 1 139
2 903 1 139
2 904 1 142
2 905 1 142
2 906 1 144
2 907 1 144
2 908 1 147
2 909 1 147
2 910 1 150
2 911 1 150
2 912 1 152
2 913 1 152
2 914 1 155
2 915 1 155
2 916 1 158
2 917 1 158
2 918 1 160
2 919 1 160
2 920 1 163
2 921 1 163
2 922 1 166
2 923 1 166
2 924 1 168
2 925 1 168
2 926 1 171
2 927 1 171
2 928 1 174
2 929 1 174
2 930 1 176
2 931 1 176
2 932 1 179
2 933 1 179
2 934 1 182
2 935 1 182
2 936 1 184
2 937 1 184
2 938 1 187
2 939 1 187
2 940 1 190
2 941 1 190
2 942 1 192
2 943 1 192
2 944 1 195
2 945 1 195
2 946 1 198
2 947 1 198
2 948 1 200
2 949 1 200
2 950 1 203
2 951 1 203
2 952 1 206
2 953 1 206
2 954 1 208
2 955 1 208
2 956 1 211
2 957 1 211
2 958 1 214
2 959 1 214
2 960 1 216
2 961 1 216
2 962 1 219
2 963 1 219
2 964 1 221
2 965 1 221
2 966 1 222
2 967 1 222
2 968 1 223
2 969 1 223
2 970 1 224
2 971 1 224
2 972 1 225
2 973 1 225
2 974 1 231
2 975 1 231
2 976 1 234
2 977 1 234
2 978 1 234
2 979 1 235
2 980 1 235
2 981 1 241
2 982 1 241
2 983 1 244
2 984 1 244
2 985 1 244
2 986 1 244
2 987 1 246
2 988 1 246
2 989 1 246
2 990 1 247
2 991 1 247
2 992 1 253
2 993 1 253
2 994 1 256
2 995 1 256
2 996 1 256
2 997 1 256
2 998 1 258
2 999 1 258
2 1000 1 258
2 1001 1 259
2 1002 1 259
2 1003 1 265
2 1004 1 265
2 1005 1 268
2 1006 1 268
2 1007 1 268
2 1008 1 268
2 1009 1 269
2 1010 1 269
2 1011 1 275
2 1012 1 275
2 1013 1 278
2 1014 1 278
2 1015 1 278
2 1016 1 278
2 1017 1 280
2 1018 1 280
2 1019 1 280
2 1020 1 280
2 1021 1 281
2 1022 1 281
2 1023 1 287
2 1024 1 287
2 1025 1 290
2 1026 1 290
2 1027 1 290
2 1028 1 290
2 1029 1 292
2 1030 1 292
2 1031 1 292
2 1032 1 292
2 1033 1 293
2 1034 1 293
2 1035 1 299
2 1036 1 299
2 1037 1 302
2 1038 1 302
2 1039 1 302
2 1040 1 302
2 1041 1 304
2 1042 1 304
2 1043 1 304
2 1044 1 304
2 1045 1 305
2 1046 1 305
2 1047 1 311
2 1048 1 311
2 1049 1 314
2 1050 1 314
2 1051 1 314
2 1052 1 314
2 1053 1 316
2 1054 1 316
2 1055 1 316
2 1056 1 317
2 1057 1 317
2 1058 1 323
2 1059 1 323
2 1060 1 326
2 1061 1 326
2 1062 1 326
2 1063 1 328
2 1064 1 328
2 1065 1 328
2 1066 1 328
2 1067 1 329
2 1068 1 329
2 1069 1 335
2 1070 1 335
2 1071 1 338
2 1072 1 338
2 1073 1 338
2 1074 1 340
2 1075 1 340
2 1076 1 340
2 1077 1 341
2 1078 1 341
2 1079 1 347
2 1080 1 347
2 1081 1 350
2 1082 1 350
2 1083 1 350
2 1084 1 352
2 1085 1 352
2 1086 1 352
2 1087 1 353
2 1088 1 353
2 1089 1 359
2 1090 1 359
2 1091 1 362
2 1092 1 362
2 1093 1 362
2 1094 1 364
2 1095 1 364
2 1096 1 364
2 1097 1 365
2 1098 1 365
2 1099 1 371
2 1100 1 371
2 1101 1 374
2 1102 1 374
2 1103 1 374
2 1104 1 376
2 1105 1 376
2 1106 1 376
2 1107 1 377
2 1108 1 377
2 1109 1 383
2 1110 1 383
2 1111 1 386
2 1112 1 386
2 1113 1 386
2 1114 1 388
2 1115 1 388
2 1116 1 388
2 1117 1 389
2 1118 1 389
2 1119 1 395
2 1120 1 395
2 1121 1 398
2 1122 1 398
2 1123 1 400
2 1124 1 400
2 1125 1 403
2 1126 1 403
2 1127 1 407
2 1128 1 407
2 1129 1 409
2 1130 1 409
2 1131 1 410
2 1132 1 410
2 1133 1 413
2 1134 1 413
2 1135 1 414
2 1136 1 414
2 1137 1 417
2 1138 1 417
2 1139 1 418
2 1140 1 418
2 1141 1 421
2 1142 1 421
2 1143 1 422
2 1144 1 422
2 1145 1 425
2 1146 1 425
2 1147 1 426
2 1148 1 426
2 1149 1 429
2 1150 1 429
2 1151 1 430
2 1152 1 430
2 1153 1 433
2 1154 1 433
2 1155 1 435
2 1156 1 435
2 1157 1 437
2 1158 1 437
2 1159 1 439
2 1160 1 439
2 1161 1 441
2 1162 1 441
2 1163 1 444
2 1164 1 444
2 1165 1 448
2 1166 1 448
2 1167 1 453
2 1168 1 453
2 1169 1 453
2 1170 1 453
2 1171 1 456
2 1172 1 456
2 1173 1 462
2 1174 1 462
2 1175 1 464
2 1176 1 464
2 1177 1 464
2 1178 1 467
2 1179 1 467
2 1180 1 471
2 1181 1 471
2 1182 1 475
2 1183 1 475
2 1184 1 475
2 1185 1 476
2 1186 1 476
2 1187 1 481
2 1188 1 481
2 1189 1 481
2 1190 1 487
2 1191 1 487
2 1192 1 488
2 1193 1 488
2 1194 1 491
2 1195 1 491
2 1196 1 496
2 1197 1 496
2 1198 1 502
2 1199 1 502
2 1200 1 508
2 1201 1 508
2 1202 1 513
2 1203 1 513
2 1204 1 514
2 1205 1 514
2 1206 1 517
2 1207 1 517
2 1208 1 518
2 1209 1 518
2 1210 1 521
2 1211 1 521
2 1212 1 521
2 1213 1 522
2 1214 1 522
2 1215 1 525
2 1216 1 525
2 1217 1 525
2 1218 1 526
2 1219 1 526
2 1220 1 533
2 1221 1 533
2 1222 1 533
2 1223 1 534
2 1224 1 534
2 1225 1 539
2 1226 1 539
2 1227 1 539
2 1228 1 540
2 1229 1 540
2 1230 1 545
2 1231 1 545
2 1232 1 545
2 1233 1 546
2 1234 1 546
2 1235 1 553
2 1236 1 553
2 1237 1 556
2 1238 1 556
2 1239 1 591
2 1240 1 591
2 1241 1 591
2 1242 1 595
2 1243 1 595
2 1244 1 595
2 1245 1 599
2 1246 1 599
2 1247 1 600
2 1248 1 600
2 1249 1 603
2 1250 1 603
2 1251 1 604
2 1252 1 604
2 1253 1 607
2 1254 1 607
2 1255 1 608
2 1256 1 608
2 1257 1 611
2 1258 1 611
2 1259 1 613
2 1260 1 613
2 1261 1 615
2 1262 1 615
2 1263 1 616
2 1264 1 616
2 1265 1 619
2 1266 1 619
2 1267 1 621
2 1268 1 621
2 1269 1 623
2 1270 1 623
2 1271 1 626
2 1272 1 626
2 1273 1 630
2 1274 1 630
2 1275 1 635
2 1276 1 635
2 1277 1 639
2 1278 1 639
2 1279 1 640
2 1280 1 640
2 1281 1 643
2 1282 1 643
2 1283 1 644
2 1284 1 644
2 1285 1 733
2 1286 1 733
0 50 5 1 1 49
0 51 5 1 1 745
0 52 5 1 1 747
0 53 5 1 1 749
0 54 5 1 1 751
0 55 5 1 1 753
0 56 5 1 1 755
0 57 5 1 1 757
0 58 5 1 1 759
0 59 5 1 1 761
0 60 5 1 1 763
0 61 5 1 1 765
0 62 5 1 1 767
0 63 5 1 1 769
0 64 5 1 1 771
0 65 5 1 1 773
0 66 5 1 1 775
0 67 5 1 1 777
0 68 5 1 1 779
0 69 5 2 1 781
0 70 5 2 1 783
0 71 5 2 1 785
0 72 5 2 1 787
0 73 5 2 1 789
0 74 5 2 1 791
0 75 5 2 1 793
0 76 5 2 1 795
0 77 5 2 1 797
0 78 5 2 1 799
0 79 5 2 1 801
0 80 5 2 1 803
0 81 5 2 1 805
0 82 5 1 1 807
0 83 5 1 1 809
0 84 5 1 1 811
0 85 5 1 1 813
0 86 5 1 1 815
0 87 5 1 1 817
0 88 5 1 1 819
0 89 5 1 1 821
0 90 5 1 1 823
0 91 5 1 1 825
0 92 5 1 1 827
0 93 5 1 1 829
0 94 5 1 1 831
0 95 5 1 1 833
0 96 5 1 1 835
0 97 5 1 1 837
0 98 5 1 1 839
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 748 780
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 746 778
0 106 5 2 1 105
0 107 7 2 2 744 776
0 108 5 3 1 875
0 109 7 1 2 873 877
0 110 5 1 1 109
0 111 7 2 2 871 110
0 112 5 2 1 880
0 113 7 1 2 869 882
0 114 5 1 1 113
0 115 7 2 2 867 114
0 116 5 1 1 884
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 750 885
0 120 5 2 1 119
0 121 7 1 2 841 888
0 122 5 1 1 121
0 123 7 2 2 886 122
0 124 5 1 1 890
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 752 891
0 128 5 2 1 127
0 129 7 1 2 843 894
0 130 5 1 1 129
0 131 7 2 2 892 130
0 132 5 1 1 896
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 754 897
0 136 5 2 1 135
0 137 7 1 2 845 900
0 138 5 1 1 137
0 139 7 2 2 898 138
0 140 5 1 1 902
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 756 903
0 144 5 2 1 143
0 145 7 1 2 847 906
0 146 5 1 1 145
0 147 7 2 2 904 146
0 148 5 1 1 908
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 758 909
0 152 5 2 1 151
0 153 7 1 2 849 912
0 154 5 1 1 153
0 155 7 2 2 910 154
0 156 5 1 1 914
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 760 915
0 160 5 2 1 159
0 161 7 1 2 851 918
0 162 5 1 1 161
0 163 7 2 2 916 162
0 164 5 1 1 920
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 762 921
0 168 5 2 1 167
0 169 7 1 2 853 924
0 170 5 1 1 169
0 171 7 2 2 922 170
0 172 5 1 1 926
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 764 927
0 176 5 2 1 175
0 177 7 1 2 855 930
0 178 5 1 1 177
0 179 7 2 2 928 178
0 180 5 1 1 932
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 766 933
0 184 5 2 1 183
0 185 7 1 2 857 936
0 186 5 1 1 185
0 187 7 2 2 934 186
0 188 5 1 1 938
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 768 939
0 192 5 2 1 191
0 193 7 1 2 859 942
0 194 5 1 1 193
0 195 7 2 2 940 194
0 196 5 1 1 944
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 770 945
0 200 5 2 1 199
0 201 7 1 2 861 948
0 202 5 1 1 201
0 203 7 2 2 946 202
0 204 5 1 1 950
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 772 951
0 208 5 2 1 207
0 209 7 1 2 863 954
0 210 5 1 1 209
0 211 7 2 2 952 210
0 212 5 1 1 956
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 774 957
0 216 5 2 1 215
0 217 7 1 2 865 960
0 218 5 1 1 217
0 219 7 2 2 958 218
0 220 5 1 1 962
0 221 7 2 2 840 220
0 222 5 2 1 964
0 223 7 2 2 98 963
0 224 5 2 1 968
0 225 7 2 2 959 961
0 226 5 1 1 972
0 227 7 1 2 806 226
0 228 5 1 1 227
0 229 7 1 2 866 973
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 974
0 233 7 1 2 838 975
0 234 5 3 1 233
0 235 7 2 2 953 955
0 236 5 1 1 979
0 237 7 1 2 804 980
0 238 5 1 1 237
0 239 7 1 2 864 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 981
0 243 7 1 2 836 242
0 244 5 4 1 243
0 245 7 1 2 96 982
0 246 5 3 1 245
0 247 7 2 2 947 949
0 248 5 1 1 990
0 249 7 1 2 802 991
0 250 5 1 1 249
0 251 7 1 2 862 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 992
0 255 7 1 2 834 254
0 256 5 4 1 255
0 257 7 1 2 95 993
0 258 5 3 1 257
0 259 7 2 2 941 943
0 260 5 1 1 1001
0 261 7 1 2 800 1002
0 262 5 1 1 261
0 263 7 1 2 860 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 1003
0 267 7 1 2 832 266
0 268 5 4 1 267
0 269 7 2 2 935 937
0 270 5 1 1 1009
0 271 7 1 2 798 1010
0 272 5 1 1 271
0 273 7 1 2 858 270
0 274 5 1 1 273
0 275 7 2 2 272 274
0 276 5 1 1 1011
0 277 7 1 2 830 276
0 278 5 4 1 277
0 279 7 1 2 93 1012
0 280 5 4 1 279
0 281 7 2 2 929 931
0 282 5 1 1 1021
0 283 7 1 2 796 1022
0 284 5 1 1 283
0 285 7 1 2 856 282
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 1023
0 289 7 1 2 828 288
0 290 5 4 1 289
0 291 7 1 2 92 1024
0 292 5 4 1 291
0 293 7 2 2 923 925
0 294 5 1 1 1033
0 295 7 1 2 794 1034
0 296 5 1 1 295
0 297 7 1 2 854 294
0 298 5 1 1 297
0 299 7 2 2 296 298
0 300 5 1 1 1035
0 301 7 1 2 91 1036
0 302 5 4 1 301
0 303 7 1 2 826 300
0 304 5 4 1 303
0 305 7 2 2 917 919
0 306 5 1 1 1045
0 307 7 1 2 792 1046
0 308 5 1 1 307
0 309 7 1 2 852 306
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 1047
0 313 7 1 2 824 312
0 314 5 4 1 313
0 315 7 1 2 90 1048
0 316 5 3 1 315
0 317 7 2 2 911 913
0 318 5 1 1 1056
0 319 7 1 2 790 1057
0 320 5 1 1 319
0 321 7 1 2 850 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1058
0 325 7 1 2 89 1059
0 326 5 3 1 325
0 327 7 1 2 822 324
0 328 5 4 1 327
0 329 7 2 2 905 907
0 330 5 1 1 1067
0 331 7 1 2 788 1068
0 332 5 1 1 331
0 333 7 1 2 848 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1069
0 337 7 1 2 88 1070
0 338 5 3 1 337
0 339 7 1 2 820 336
0 340 5 3 1 339
0 341 7 2 2 899 901
0 342 5 1 1 1077
0 343 7 1 2 786 1078
0 344 5 1 1 343
0 345 7 1 2 846 342
0 346 5 1 1 345
0 347 7 2 2 344 346
0 348 5 1 1 1079
0 349 7 1 2 87 1080
0 350 5 3 1 349
0 351 7 1 2 818 348
0 352 5 3 1 351
0 353 7 2 2 893 895
0 354 5 1 1 1087
0 355 7 1 2 784 1088
0 356 5 1 1 355
0 357 7 1 2 844 354
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 1089
0 361 7 1 2 86 1090
0 362 5 3 1 361
0 363 7 1 2 816 360
0 364 5 3 1 363
0 365 7 2 2 887 889
0 366 5 1 1 1097
0 367 7 1 2 782 1098
0 368 5 1 1 367
0 369 7 1 2 842 366
0 370 5 1 1 369
0 371 7 2 2 368 370
0 372 5 1 1 1099
0 373 7 1 2 85 1100
0 374 5 3 1 373
0 375 7 1 2 814 372
0 376 5 3 1 375
0 377 7 2 2 868 870
0 378 5 1 1 1107
0 379 7 1 2 881 378
0 380 5 1 1 379
0 381 7 1 2 883 1108
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 1109
0 385 7 1 2 84 384
0 386 5 3 1 385
0 387 7 1 2 812 1110
0 388 5 3 1 387
0 389 7 2 2 872 874
0 390 5 1 1 1117
0 391 7 1 2 876 390
0 392 5 1 1 391
0 393 7 1 2 878 1118
0 394 5 1 1 393
0 395 7 2 2 392 394
0 396 5 1 1 1119
0 397 7 1 2 83 396
0 398 5 2 1 397
0 399 7 1 2 810 1120
0 400 5 2 1 399
0 401 7 1 2 50 66
0 402 5 1 1 401
0 403 7 2 2 879 402
0 404 5 1 1 1125
0 405 7 1 2 808 404
0 406 5 1 1 405
0 407 7 2 2 1123 406
0 408 5 1 1 1127
0 409 7 2 2 1121 408
0 410 5 2 1 1129
0 411 7 1 2 1114 1131
0 412 5 1 1 411
0 413 7 2 2 1111 412
0 414 5 2 1 1133
0 415 7 1 2 1104 1135
0 416 5 1 1 415
0 417 7 2 2 1101 416
0 418 5 2 1 1137
0 419 7 1 2 1094 1139
0 420 5 1 1 419
0 421 7 2 2 1091 420
0 422 5 2 1 1141
0 423 7 1 2 1084 1143
0 424 5 1 1 423
0 425 7 2 2 1081 424
0 426 5 2 1 1145
0 427 7 1 2 1074 1147
0 428 5 1 1 427
0 429 7 2 2 1071 428
0 430 5 2 1 1149
0 431 7 1 2 1063 1151
0 432 5 1 1 431
0 433 7 2 2 1060 432
0 434 5 1 1 1153
0 435 7 2 2 1053 1154
0 436 5 1 1 1155
0 437 7 2 2 1049 436
0 438 5 1 1 1157
0 439 7 2 2 1041 1158
0 440 5 1 1 1159
0 441 7 2 2 1037 440
0 442 5 1 1 1161
0 443 7 1 2 1029 1162
0 444 5 2 1 443
0 445 7 1 2 1025 1163
0 446 5 1 1 445
0 447 7 1 2 1017 446
0 448 5 2 1 447
0 449 7 1 2 1013 1165
0 450 7 1 2 1005 449
0 451 5 1 1 450
0 452 7 1 2 94 1004
0 453 5 4 1 452
0 454 7 1 2 451 1167
0 455 7 1 2 998 454
0 456 5 2 1 455
0 457 7 1 2 994 1171
0 458 5 1 1 457
0 459 7 1 2 987 458
0 460 5 1 1 459
0 461 7 1 2 983 460
0 462 5 2 1 461
0 463 7 1 2 97 232
0 464 5 3 1 463
0 465 7 1 2 1173 1175
0 466 5 1 1 465
0 467 7 2 2 976 466
0 468 5 1 1 1178
0 469 7 1 2 970 468
0 470 5 1 1 469
0 471 7 2 2 966 470
0 472 5 1 1 1180
0 473 7 1 2 969 1179
0 474 5 1 1 473
0 475 7 3 2 1176 977
0 476 5 2 1 1182
0 477 7 1 2 984 1185
0 478 5 1 1 477
0 479 7 1 2 1174 1183
0 480 5 1 1 479
0 481 7 3 2 985 988
0 482 5 1 1 1187
0 483 7 1 2 1172 1188
0 484 5 1 1 483
0 485 7 1 2 995 484
0 486 5 1 1 485
0 487 7 2 2 996 999
0 488 5 2 1 1190
0 489 7 1 2 1006 1192
0 490 5 1 1 489
0 491 7 2 2 1007 1168
0 492 7 1 2 1166 1194
0 493 5 1 1 492
0 494 7 1 2 1014 493
0 495 5 1 1 494
0 496 7 2 2 1015 1018
0 497 7 1 2 1164 1196
0 498 5 1 1 497
0 499 7 1 2 1026 498
0 500 5 1 1 499
0 501 7 1 2 1027 1030
0 502 5 2 1 501
0 503 7 1 2 442 1198
0 504 5 1 1 503
0 505 7 1 2 1038 1160
0 506 5 1 1 505
0 507 7 1 2 1039 1042
0 508 5 2 1 507
0 509 7 1 2 438 1200
0 510 5 1 1 509
0 511 7 1 2 1050 1156
0 512 5 1 1 511
0 513 7 2 2 1051 1054
0 514 5 2 1 1202
0 515 7 1 2 434 1204
0 516 5 1 1 515
0 517 7 2 2 1061 1064
0 518 5 2 1 1206
0 519 7 1 2 1152 1207
0 520 5 1 1 519
0 521 7 3 2 1072 1075
0 522 5 2 1 1210
0 523 7 1 2 1146 1211
0 524 5 1 1 523
0 525 7 3 2 1082 1085
0 526 5 2 1 1215
0 527 7 1 2 1142 1216
0 528 5 1 1 527
0 529 7 1 2 1144 1218
0 530 5 1 1 529
0 531 7 1 2 528 530
0 532 5 1 1 531
0 533 7 3 2 1092 1095
0 534 5 2 1 1220
0 535 7 1 2 1138 1223
0 536 5 1 1 535
0 537 7 1 2 1140 1221
0 538 5 1 1 537
0 539 7 3 2 1102 1105
0 540 5 2 1 1225
0 541 7 1 2 1136 1226
0 542 5 1 1 541
0 543 7 1 2 1134 1228
0 544 5 1 1 543
0 545 7 3 2 1112 1115
0 546 5 2 1 1230
0 547 7 1 2 1130 1233
0 548 5 1 1 547
0 549 7 1 2 1132 1231
0 550 5 1 1 549
0 551 7 1 2 82 1126
0 552 5 1 1 551
0 553 7 2 2 1122 552
0 554 5 1 1 1235
0 555 7 1 2 1128 1236
0 556 5 2 1 555
0 557 7 1 2 550 1237
0 558 7 1 2 548 557
0 559 7 1 2 544 558
0 560 7 1 2 542 559
0 561 7 1 2 538 560
0 562 7 1 2 536 561
0 563 7 1 2 532 562
0 564 5 1 1 563
0 565 7 1 2 1148 1213
0 566 5 1 1 565
0 567 7 1 2 564 566
0 568 7 1 2 524 567
0 569 5 1 1 568
0 570 7 1 2 1150 1208
0 571 5 1 1 570
0 572 7 1 2 569 571
0 573 7 1 2 520 572
0 574 5 1 1 573
0 575 7 1 2 516 574
0 576 7 1 2 512 575
0 577 5 1 1 576
0 578 7 1 2 510 577
0 579 7 1 2 506 578
0 580 5 1 1 579
0 581 7 1 2 504 580
0 582 7 1 2 500 581
0 583 7 1 2 495 582
0 584 7 1 2 490 583
0 585 7 1 2 486 584
0 586 7 1 2 480 585
0 587 7 1 2 478 586
0 588 7 1 2 474 587
0 589 7 1 2 1181 588
0 590 5 1 1 589
0 591 7 3 2 1124 554
0 592 5 1 1 1239
0 593 7 1 2 1116 1240
0 594 5 1 1 593
0 595 7 3 2 1113 594
0 596 5 1 1 1242
0 597 7 1 2 1103 1243
0 598 5 1 1 597
0 599 7 2 2 1106 598
0 600 5 2 1 1245
0 601 7 1 2 1093 1247
0 602 5 1 1 601
0 603 7 2 2 1096 602
0 604 5 2 1 1249
0 605 7 1 2 1083 1251
0 606 5 1 1 605
0 607 7 2 2 1086 606
0 608 5 2 1 1253
0 609 7 1 2 1073 1255
0 610 5 1 1 609
0 611 7 2 2 1076 610
0 612 5 1 1 1257
0 613 7 2 2 1062 612
0 614 5 1 1 1259
0 615 7 2 2 1065 614
0 616 5 2 1 1261
0 617 7 1 2 1055 1263
0 618 5 1 1 617
0 619 7 2 2 1052 618
0 620 5 1 1 1265
0 621 7 2 2 1040 620
0 622 5 1 1 1267
0 623 7 2 2 1043 622
0 624 5 1 1 1269
0 625 7 1 2 1028 1270
0 626 5 2 1 625
0 627 7 1 2 1031 1271
0 628 5 1 1 627
0 629 7 1 2 1016 628
0 630 5 2 1 629
0 631 7 1 2 1019 1273
0 632 5 1 1 631
0 633 7 1 2 1008 632
0 634 5 1 1 633
0 635 7 2 2 1169 634
0 636 5 1 1 1275
0 637 7 1 2 1000 1276
0 638 5 1 1 637
0 639 7 2 2 997 638
0 640 5 2 1 1277
0 641 7 1 2 989 1279
0 642 5 1 1 641
0 643 7 2 2 986 642
0 644 5 2 1 1281
0 645 7 1 2 1184 1283
0 646 5 1 1 645
0 647 7 1 2 1186 1282
0 648 5 1 1 647
0 649 7 1 2 646 648
0 650 5 1 1 649
0 651 7 1 2 1191 636
0 652 5 1 1 651
0 653 7 1 2 1170 1193
0 654 5 1 1 653
0 655 7 1 2 1195 1274
0 656 5 1 1 655
0 657 7 1 2 1020 656
0 658 5 1 1 657
0 659 7 1 2 1197 1272
0 660 5 1 1 659
0 661 7 1 2 1032 660
0 662 5 1 1 661
0 663 7 1 2 1199 624
0 664 5 1 1 663
0 665 7 1 2 1044 1268
0 666 5 1 1 665
0 667 7 1 2 1201 1266
0 668 5 1 1 667
0 669 7 1 2 1203 1262
0 670 5 1 1 669
0 671 7 1 2 1066 1260
0 672 5 1 1 671
0 673 7 1 2 1209 1258
0 674 5 1 1 673
0 675 7 1 2 1212 1254
0 676 5 1 1 675
0 677 7 1 2 1219 1250
0 678 5 1 1 677
0 679 7 1 2 1217 1252
0 680 5 1 1 679
0 681 7 1 2 1222 1248
0 682 5 1 1 681
0 683 7 1 2 1224 1246
0 684 5 1 1 683
0 685 7 1 2 1227 1244
0 686 5 1 1 685
0 687 7 1 2 1229 596
0 688 5 1 1 687
0 689 7 1 2 1234 1241
0 690 5 1 1 689
0 691 7 1 2 1232 592
0 692 5 1 1 691
0 693 7 1 2 1238 692
0 694 7 1 2 690 693
0 695 7 1 2 688 694
0 696 7 1 2 686 695
0 697 7 1 2 684 696
0 698 7 1 2 682 697
0 699 7 1 2 680 698
0 700 7 1 2 678 699
0 701 5 1 1 700
0 702 7 1 2 1214 1256
0 703 5 1 1 702
0 704 7 1 2 701 703
0 705 7 1 2 676 704
0 706 5 1 1 705
0 707 7 1 2 674 706
0 708 7 1 2 672 707
0 709 5 1 1 708
0 710 7 1 2 1205 1264
0 711 5 1 1 710
0 712 7 1 2 709 711
0 713 7 1 2 670 712
0 714 5 1 1 713
0 715 7 1 2 668 714
0 716 7 1 2 666 715
0 717 5 1 1 716
0 718 7 1 2 664 717
0 719 7 1 2 662 718
0 720 7 1 2 658 719
0 721 7 1 2 654 720
0 722 7 1 2 652 721
0 723 7 1 2 971 722
0 724 7 1 2 482 1280
0 725 5 1 1 724
0 726 7 1 2 1189 1278
0 727 5 1 1 726
0 728 7 1 2 725 727
0 729 7 1 2 723 728
0 730 7 1 2 650 729
0 731 7 1 2 1177 1284
0 732 5 1 1 731
0 733 7 2 2 978 732
0 734 5 1 1 1285
0 735 7 1 2 965 734
0 736 5 1 1 735
0 737 7 1 2 967 1286
0 738 5 1 1 737
0 739 7 1 2 736 738
0 740 7 1 2 730 739
0 741 7 1 2 472 740
0 742 5 1 1 741
0 743 7 1 2 590 742
3 3499 5 0 1 743
