1 0 0 2 0
2 49 1 0
2 717 1 0
1 1 0 2 0
2 718 1 1
2 719 1 1
1 2 0 2 0
2 720 1 2
2 721 1 2
1 3 0 2 0
2 722 1 3
2 723 1 3
1 4 0 2 0
2 724 1 4
2 725 1 4
1 5 0 2 0
2 726 1 5
2 727 1 5
1 6 0 2 0
2 728 1 6
2 729 1 6
1 7 0 2 0
2 730 1 7
2 731 1 7
1 8 0 2 0
2 732 1 8
2 733 1 8
1 9 0 2 0
2 734 1 9
2 735 1 9
1 10 0 2 0
2 736 1 10
2 737 1 10
1 11 0 2 0
2 738 1 11
2 739 1 11
1 12 0 2 0
2 740 1 12
2 741 1 12
1 13 0 2 0
2 742 1 13
2 743 1 13
1 14 0 2 0
2 744 1 14
2 745 1 14
1 15 0 2 0
2 746 1 15
2 747 1 15
1 16 0 2 0
2 748 1 16
2 749 1 16
1 17 0 2 0
2 750 1 17
2 751 1 17
1 18 0 2 0
2 752 1 18
2 753 1 18
1 19 0 2 0
2 754 1 19
2 755 1 19
1 20 0 2 0
2 756 1 20
2 757 1 20
1 21 0 2 0
2 758 1 21
2 759 1 21
1 22 0 2 0
2 760 1 22
2 761 1 22
1 23 0 2 0
2 762 1 23
2 763 1 23
1 24 0 2 0
2 764 1 24
2 765 1 24
1 25 0 2 0
2 766 1 25
2 767 1 25
1 26 0 2 0
2 768 1 26
2 769 1 26
1 27 0 2 0
2 770 1 27
2 771 1 27
1 28 0 2 0
2 772 1 28
2 773 1 28
1 29 0 2 0
2 774 1 29
2 775 1 29
1 30 0 2 0
2 776 1 30
2 777 1 30
1 31 0 2 0
2 778 1 31
2 779 1 31
1 32 0 2 0
2 780 1 32
2 781 1 32
1 33 0 2 0
2 782 1 33
2 783 1 33
1 34 0 2 0
2 784 1 34
2 785 1 34
1 35 0 2 0
2 786 1 35
2 787 1 35
1 36 0 2 0
2 788 1 36
2 789 1 36
1 37 0 2 0
2 790 1 37
2 791 1 37
1 38 0 2 0
2 792 1 38
2 793 1 38
1 39 0 2 0
2 794 1 39
2 795 1 39
1 40 0 2 0
2 796 1 40
2 797 1 40
1 41 0 2 0
2 798 1 41
2 799 1 41
1 42 0 2 0
2 800 1 42
2 801 1 42
1 43 0 2 0
2 802 1 43
2 803 1 43
1 44 0 2 0
2 804 1 44
2 805 1 44
1 45 0 2 0
2 806 1 45
2 807 1 45
1 46 0 2 0
2 808 1 46
2 809 1 46
1 47 0 2 0
2 810 1 47
2 811 1 47
1 48 0 2 0
2 812 1 48
2 813 1 48
2 814 1 69
2 815 1 69
2 816 1 70
2 817 1 70
2 818 1 71
2 819 1 71
2 820 1 72
2 821 1 72
2 822 1 73
2 823 1 73
2 824 1 74
2 825 1 74
2 826 1 75
2 827 1 75
2 828 1 76
2 829 1 76
2 830 1 77
2 831 1 77
2 832 1 78
2 833 1 78
2 834 1 79
2 835 1 79
2 836 1 80
2 837 1 80
2 838 1 81
2 839 1 81
2 840 1 100
2 841 1 100
2 842 1 102
2 843 1 102
2 844 1 104
2 845 1 104
2 846 1 106
2 847 1 106
2 848 1 107
2 849 1 107
2 850 1 108
2 851 1 108
2 852 1 108
2 853 1 111
2 854 1 111
2 855 1 112
2 856 1 112
2 857 1 115
2 858 1 115
2 859 1 118
2 860 1 118
2 861 1 120
2 862 1 120
2 863 1 123
2 864 1 123
2 865 1 126
2 866 1 126
2 867 1 128
2 868 1 128
2 869 1 131
2 870 1 131
2 871 1 134
2 872 1 134
2 873 1 136
2 874 1 136
2 875 1 139
2 876 1 139
2 877 1 142
2 878 1 142
2 879 1 144
2 880 1 144
2 881 1 147
2 882 1 147
2 883 1 150
2 884 1 150
2 885 1 152
2 886 1 152
2 887 1 155
2 888 1 155
2 889 1 158
2 890 1 158
2 891 1 160
2 892 1 160
2 893 1 163
2 894 1 163
2 895 1 166
2 896 1 166
2 897 1 168
2 898 1 168
2 899 1 171
2 900 1 171
2 901 1 174
2 902 1 174
2 903 1 176
2 904 1 176
2 905 1 179
2 906 1 179
2 907 1 182
2 908 1 182
2 909 1 184
2 910 1 184
2 911 1 187
2 912 1 187
2 913 1 190
2 914 1 190
2 915 1 192
2 916 1 192
2 917 1 195
2 918 1 195
2 919 1 198
2 920 1 198
2 921 1 200
2 922 1 200
2 923 1 203
2 924 1 203
2 925 1 206
2 926 1 206
2 927 1 208
2 928 1 208
2 929 1 211
2 930 1 211
2 931 1 214
2 932 1 214
2 933 1 216
2 934 1 216
2 935 1 219
2 936 1 219
2 937 1 221
2 938 1 221
2 939 1 222
2 940 1 222
2 941 1 223
2 942 1 223
2 943 1 224
2 944 1 224
2 945 1 225
2 946 1 225
2 947 1 231
2 948 1 231
2 949 1 234
2 950 1 234
2 951 1 234
2 952 1 235
2 953 1 235
2 954 1 241
2 955 1 241
2 956 1 244
2 957 1 244
2 958 1 244
2 959 1 244
2 960 1 246
2 961 1 246
2 962 1 246
2 963 1 247
2 964 1 247
2 965 1 253
2 966 1 253
2 967 1 256
2 968 1 256
2 969 1 256
2 970 1 256
2 971 1 258
2 972 1 258
2 973 1 258
2 974 1 259
2 975 1 259
2 976 1 265
2 977 1 265
2 978 1 268
2 979 1 268
2 980 1 268
2 981 1 268
2 982 1 270
2 983 1 270
2 984 1 270
2 985 1 271
2 986 1 271
2 987 1 277
2 988 1 277
2 989 1 280
2 990 1 280
2 991 1 280
2 992 1 280
2 993 1 281
2 994 1 281
2 995 1 287
2 996 1 287
2 997 1 290
2 998 1 290
2 999 1 290
2 1000 1 290
2 1001 1 292
2 1002 1 292
2 1003 1 292
2 1004 1 292
2 1005 1 293
2 1006 1 293
2 1007 1 299
2 1008 1 299
2 1009 1 302
2 1010 1 302
2 1011 1 302
2 1012 1 302
2 1013 1 304
2 1014 1 304
2 1015 1 304
2 1016 1 305
2 1017 1 305
2 1018 1 311
2 1019 1 311
2 1020 1 314
2 1021 1 314
2 1022 1 314
2 1023 1 316
2 1024 1 316
2 1025 1 316
2 1026 1 317
2 1027 1 317
2 1028 1 323
2 1029 1 323
2 1030 1 326
2 1031 1 326
2 1032 1 326
2 1033 1 326
2 1034 1 328
2 1035 1 328
2 1036 1 328
2 1037 1 329
2 1038 1 329
2 1039 1 335
2 1040 1 335
2 1041 1 338
2 1042 1 338
2 1043 1 338
2 1044 1 338
2 1045 1 340
2 1046 1 340
2 1047 1 340
2 1048 1 341
2 1049 1 341
2 1050 1 347
2 1051 1 347
2 1052 1 350
2 1053 1 350
2 1054 1 350
2 1055 1 350
2 1056 1 350
2 1057 1 352
2 1058 1 352
2 1059 1 352
2 1060 1 352
2 1061 1 353
2 1062 1 353
2 1063 1 359
2 1064 1 359
2 1065 1 361
2 1066 1 361
2 1067 1 361
2 1068 1 362
2 1069 1 362
2 1070 1 363
2 1071 1 363
2 1072 1 363
2 1073 1 364
2 1074 1 364
2 1075 1 365
2 1076 1 365
2 1077 1 371
2 1078 1 371
2 1079 1 374
2 1080 1 374
2 1081 1 374
2 1082 1 376
2 1083 1 376
2 1084 1 376
2 1085 1 377
2 1086 1 377
2 1087 1 383
2 1088 1 383
2 1089 1 386
2 1090 1 386
2 1091 1 386
2 1092 1 386
2 1093 1 388
2 1094 1 388
2 1095 1 388
2 1096 1 389
2 1097 1 389
2 1098 1 395
2 1099 1 395
2 1100 1 398
2 1101 1 398
2 1102 1 400
2 1103 1 400
2 1104 1 403
2 1105 1 403
2 1106 1 409
2 1107 1 409
2 1108 1 410
2 1109 1 410
2 1110 1 413
2 1111 1 413
2 1112 1 413
2 1113 1 417
2 1114 1 417
2 1115 1 418
2 1116 1 418
2 1117 1 424
2 1118 1 424
2 1119 1 428
2 1120 1 428
2 1121 1 429
2 1122 1 429
2 1123 1 432
2 1124 1 432
2 1125 1 433
2 1126 1 433
2 1127 1 436
2 1128 1 436
2 1129 1 439
2 1130 1 439
2 1131 1 443
2 1132 1 443
2 1133 1 448
2 1134 1 448
2 1135 1 448
2 1136 1 448
2 1137 1 451
2 1138 1 451
2 1139 1 455
2 1140 1 455
2 1141 1 461
2 1142 1 461
2 1143 1 463
2 1144 1 463
2 1145 1 463
2 1146 1 466
2 1147 1 466
2 1148 1 470
2 1149 1 470
2 1150 1 474
2 1151 1 474
2 1152 1 474
2 1153 1 475
2 1154 1 475
2 1155 1 480
2 1156 1 480
2 1157 1 480
2 1158 1 486
2 1159 1 486
2 1160 1 486
2 1161 1 492
2 1162 1 492
2 1163 1 493
2 1164 1 493
2 1165 1 496
2 1166 1 496
2 1167 1 501
2 1168 1 501
2 1169 1 507
2 1170 1 507
2 1171 1 507
2 1172 1 508
2 1173 1 508
2 1174 1 513
2 1175 1 513
2 1176 1 514
2 1177 1 514
2 1178 1 519
2 1179 1 519
2 1180 1 519
2 1181 1 520
2 1182 1 520
2 1183 1 533
2 1184 1 533
2 1185 1 533
2 1186 1 534
2 1187 1 534
2 1188 1 538
2 1189 1 538
2 1190 1 540
2 1191 1 540
2 1192 1 544
2 1193 1 544
2 1194 1 565
2 1195 1 565
2 1196 1 566
2 1197 1 566
2 1198 1 584
2 1199 1 584
2 1200 1 587
2 1201 1 587
2 1202 1 588
2 1203 1 588
2 1204 1 598
2 1205 1 598
2 1206 1 600
2 1207 1 600
2 1208 1 601
2 1209 1 601
2 1210 1 604
2 1211 1 604
2 1212 1 605
2 1213 1 605
2 1214 1 608
2 1215 1 608
2 1216 1 611
2 1217 1 611
2 1218 1 616
2 1219 1 616
2 1220 1 620
2 1221 1 620
2 1222 1 621
2 1223 1 621
2 1224 1 624
2 1225 1 624
2 1226 1 625
2 1227 1 625
2 1228 1 628
2 1229 1 628
2 1230 1 629
2 1231 1 629
2 1232 1 706
2 1233 1 706
0 50 5 1 1 49
0 51 5 1 1 718
0 52 5 1 1 720
0 53 5 1 1 722
0 54 5 1 1 724
0 55 5 1 1 726
0 56 5 1 1 728
0 57 5 1 1 730
0 58 5 1 1 732
0 59 5 1 1 734
0 60 5 1 1 736
0 61 5 1 1 738
0 62 5 1 1 740
0 63 5 1 1 742
0 64 5 1 1 744
0 65 5 1 1 746
0 66 5 1 1 748
0 67 5 1 1 750
0 68 5 1 1 752
0 69 5 2 1 754
0 70 5 2 1 756
0 71 5 2 1 758
0 72 5 2 1 760
0 73 5 2 1 762
0 74 5 2 1 764
0 75 5 2 1 766
0 76 5 2 1 768
0 77 5 2 1 770
0 78 5 2 1 772
0 79 5 2 1 774
0 80 5 2 1 776
0 81 5 2 1 778
0 82 5 1 1 780
0 83 5 1 1 782
0 84 5 1 1 784
0 85 5 1 1 786
0 86 5 1 1 788
0 87 5 1 1 790
0 88 5 1 1 792
0 89 5 1 1 794
0 90 5 1 1 796
0 91 5 1 1 798
0 92 5 1 1 800
0 93 5 1 1 802
0 94 5 1 1 804
0 95 5 1 1 806
0 96 5 1 1 808
0 97 5 1 1 810
0 98 5 1 1 812
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 721 753
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 719 751
0 106 5 2 1 105
0 107 7 2 2 717 749
0 108 5 3 1 848
0 109 7 1 2 846 850
0 110 5 1 1 109
0 111 7 2 2 844 110
0 112 5 2 1 853
0 113 7 1 2 842 855
0 114 5 1 1 113
0 115 7 2 2 840 114
0 116 5 1 1 857
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 723 858
0 120 5 2 1 119
0 121 7 1 2 814 861
0 122 5 1 1 121
0 123 7 2 2 859 122
0 124 5 1 1 863
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 725 864
0 128 5 2 1 127
0 129 7 1 2 816 867
0 130 5 1 1 129
0 131 7 2 2 865 130
0 132 5 1 1 869
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 727 870
0 136 5 2 1 135
0 137 7 1 2 818 873
0 138 5 1 1 137
0 139 7 2 2 871 138
0 140 5 1 1 875
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 729 876
0 144 5 2 1 143
0 145 7 1 2 820 879
0 146 5 1 1 145
0 147 7 2 2 877 146
0 148 5 1 1 881
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 731 882
0 152 5 2 1 151
0 153 7 1 2 822 885
0 154 5 1 1 153
0 155 7 2 2 883 154
0 156 5 1 1 887
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 733 888
0 160 5 2 1 159
0 161 7 1 2 824 891
0 162 5 1 1 161
0 163 7 2 2 889 162
0 164 5 1 1 893
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 735 894
0 168 5 2 1 167
0 169 7 1 2 826 897
0 170 5 1 1 169
0 171 7 2 2 895 170
0 172 5 1 1 899
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 737 900
0 176 5 2 1 175
0 177 7 1 2 828 903
0 178 5 1 1 177
0 179 7 2 2 901 178
0 180 5 1 1 905
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 739 906
0 184 5 2 1 183
0 185 7 1 2 830 909
0 186 5 1 1 185
0 187 7 2 2 907 186
0 188 5 1 1 911
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 741 912
0 192 5 2 1 191
0 193 7 1 2 832 915
0 194 5 1 1 193
0 195 7 2 2 913 194
0 196 5 1 1 917
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 743 918
0 200 5 2 1 199
0 201 7 1 2 834 921
0 202 5 1 1 201
0 203 7 2 2 919 202
0 204 5 1 1 923
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 745 924
0 208 5 2 1 207
0 209 7 1 2 836 927
0 210 5 1 1 209
0 211 7 2 2 925 210
0 212 5 1 1 929
0 213 7 1 2 65 212
0 214 5 2 1 213
0 215 7 1 2 747 930
0 216 5 2 1 215
0 217 7 1 2 838 933
0 218 5 1 1 217
0 219 7 2 2 931 218
0 220 5 1 1 935
0 221 7 2 2 813 220
0 222 5 2 1 937
0 223 7 2 2 98 936
0 224 5 2 1 941
0 225 7 2 2 932 934
0 226 5 1 1 945
0 227 7 1 2 779 226
0 228 5 1 1 227
0 229 7 1 2 839 946
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 947
0 233 7 1 2 811 948
0 234 5 3 1 233
0 235 7 2 2 926 928
0 236 5 1 1 952
0 237 7 1 2 777 953
0 238 5 1 1 237
0 239 7 1 2 837 236
0 240 5 1 1 239
0 241 7 2 2 238 240
0 242 5 1 1 954
0 243 7 1 2 809 242
0 244 5 4 1 243
0 245 7 1 2 96 955
0 246 5 3 1 245
0 247 7 2 2 920 922
0 248 5 1 1 963
0 249 7 1 2 775 964
0 250 5 1 1 249
0 251 7 1 2 835 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 1 1 965
0 255 7 1 2 807 254
0 256 5 4 1 255
0 257 7 1 2 95 966
0 258 5 3 1 257
0 259 7 2 2 914 916
0 260 5 1 1 974
0 261 7 1 2 773 975
0 262 5 1 1 261
0 263 7 1 2 833 260
0 264 5 1 1 263
0 265 7 2 2 262 264
0 266 5 1 1 976
0 267 7 1 2 805 266
0 268 5 4 1 267
0 269 7 1 2 94 977
0 270 5 3 1 269
0 271 7 2 2 908 910
0 272 5 1 1 985
0 273 7 1 2 771 986
0 274 5 1 1 273
0 275 7 1 2 831 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 1 1 987
0 279 7 1 2 803 278
0 280 5 4 1 279
0 281 7 2 2 902 904
0 282 5 1 1 993
0 283 7 1 2 769 994
0 284 5 1 1 283
0 285 7 1 2 829 282
0 286 5 1 1 285
0 287 7 2 2 284 286
0 288 5 1 1 995
0 289 7 1 2 801 288
0 290 5 4 1 289
0 291 7 1 2 92 996
0 292 5 4 1 291
0 293 7 2 2 896 898
0 294 5 1 1 1005
0 295 7 1 2 767 1006
0 296 5 1 1 295
0 297 7 1 2 827 294
0 298 5 1 1 297
0 299 7 2 2 296 298
0 300 5 1 1 1007
0 301 7 1 2 799 300
0 302 5 4 1 301
0 303 7 1 2 91 1008
0 304 5 3 1 303
0 305 7 2 2 890 892
0 306 5 1 1 1016
0 307 7 1 2 765 1017
0 308 5 1 1 307
0 309 7 1 2 825 306
0 310 5 1 1 309
0 311 7 2 2 308 310
0 312 5 1 1 1018
0 313 7 1 2 797 312
0 314 5 3 1 313
0 315 7 1 2 90 1019
0 316 5 3 1 315
0 317 7 2 2 884 886
0 318 5 1 1 1026
0 319 7 1 2 763 1027
0 320 5 1 1 319
0 321 7 1 2 823 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1028
0 325 7 1 2 795 324
0 326 5 4 1 325
0 327 7 1 2 89 1029
0 328 5 3 1 327
0 329 7 2 2 878 880
0 330 5 1 1 1037
0 331 7 1 2 761 1038
0 332 5 1 1 331
0 333 7 1 2 821 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1039
0 337 7 1 2 793 336
0 338 5 4 1 337
0 339 7 1 2 88 1040
0 340 5 3 1 339
0 341 7 2 2 872 874
0 342 5 1 1 1048
0 343 7 1 2 759 1049
0 344 5 1 1 343
0 345 7 1 2 819 342
0 346 5 1 1 345
0 347 7 2 2 344 346
0 348 5 1 1 1050
0 349 7 1 2 87 1051
0 350 5 5 1 349
0 351 7 1 2 791 348
0 352 5 4 1 351
0 353 7 2 2 866 868
0 354 5 1 1 1061
0 355 7 1 2 757 1062
0 356 5 1 1 355
0 357 7 1 2 817 354
0 358 5 1 1 357
0 359 7 2 2 356 358
0 360 5 1 1 1063
0 361 7 3 2 789 360
0 362 5 2 1 1065
0 363 7 3 2 86 1064
0 364 5 2 1 1070
0 365 7 2 2 860 862
0 366 5 1 1 1075
0 367 7 1 2 755 1076
0 368 5 1 1 367
0 369 7 1 2 815 366
0 370 5 1 1 369
0 371 7 2 2 368 370
0 372 5 1 1 1077
0 373 7 1 2 787 372
0 374 5 3 1 373
0 375 7 1 2 85 1078
0 376 5 3 1 375
0 377 7 2 2 841 843
0 378 5 1 1 1085
0 379 7 1 2 854 378
0 380 5 1 1 379
0 381 7 1 2 856 1086
0 382 5 1 1 381
0 383 7 2 2 380 382
0 384 5 1 1 1087
0 385 7 1 2 84 384
0 386 5 4 1 385
0 387 7 1 2 785 1088
0 388 5 3 1 387
0 389 7 2 2 845 847
0 390 5 1 1 1096
0 391 7 1 2 849 390
0 392 5 1 1 391
0 393 7 1 2 851 1097
0 394 5 1 1 393
0 395 7 2 2 392 394
0 396 5 1 1 1098
0 397 7 1 2 83 396
0 398 5 2 1 397
0 399 7 1 2 783 1099
0 400 5 2 1 399
0 401 7 1 2 50 66
0 402 5 1 1 401
0 403 7 2 2 852 402
0 404 5 1 1 1104
0 405 7 1 2 781 404
0 406 5 1 1 405
0 407 7 1 2 1102 406
0 408 5 1 1 407
0 409 7 2 2 1100 408
0 410 5 2 1 1106
0 411 7 1 2 1093 1108
0 412 5 1 1 411
0 413 7 3 2 1089 412
0 414 5 1 1 1110
0 415 7 1 2 1082 1111
0 416 5 1 1 415
0 417 7 2 2 1079 416
0 418 5 2 1 1113
0 419 7 1 2 1073 1115
0 420 5 1 1 419
0 421 7 1 2 1068 420
0 422 7 1 2 1057 421
0 423 5 1 1 422
0 424 7 2 2 1052 423
0 425 5 1 1 1117
0 426 7 1 2 1045 1118
0 427 5 1 1 426
0 428 7 2 2 1041 427
0 429 5 2 1 1119
0 430 7 1 2 1034 1121
0 431 5 1 1 430
0 432 7 2 2 1030 431
0 433 5 2 1 1123
0 434 7 1 2 1023 1125
0 435 5 1 1 434
0 436 7 2 2 1020 435
0 437 5 1 1 1127
0 438 7 1 2 1013 437
0 439 5 2 1 438
0 440 7 1 2 1009 1129
0 441 5 1 1 440
0 442 7 1 2 1001 441
0 443 5 2 1 442
0 444 7 1 2 997 1131
0 445 7 1 2 989 444
0 446 5 1 1 445
0 447 7 1 2 93 988
0 448 5 4 1 447
0 449 7 1 2 446 1133
0 450 7 1 2 982 449
0 451 5 2 1 450
0 452 7 1 2 978 1137
0 453 5 1 1 452
0 454 7 1 2 971 453
0 455 5 2 1 454
0 456 7 1 2 967 1139
0 457 5 1 1 456
0 458 7 1 2 960 457
0 459 5 1 1 458
0 460 7 1 2 956 459
0 461 5 2 1 460
0 462 7 1 2 97 232
0 463 5 3 1 462
0 464 7 1 2 1141 1143
0 465 5 1 1 464
0 466 7 2 2 949 465
0 467 5 1 1 1146
0 468 7 1 2 943 467
0 469 5 1 1 468
0 470 7 2 2 939 469
0 471 5 1 1 1148
0 472 7 1 2 942 1147
0 473 5 1 1 472
0 474 7 3 2 1144 950
0 475 5 2 1 1150
0 476 7 1 2 957 1153
0 477 5 1 1 476
0 478 7 1 2 1142 1151
0 479 5 1 1 478
0 480 7 3 2 958 961
0 481 5 1 1 1155
0 482 7 1 2 1140 1156
0 483 5 1 1 482
0 484 7 1 2 968 483
0 485 5 1 1 484
0 486 7 3 2 969 972
0 487 5 1 1 1158
0 488 7 1 2 1138 1159
0 489 5 1 1 488
0 490 7 1 2 979 489
0 491 5 1 1 490
0 492 7 2 2 980 983
0 493 5 2 1 1161
0 494 7 1 2 990 1163
0 495 5 1 1 494
0 496 7 2 2 991 1134
0 497 7 1 2 1132 1165
0 498 5 1 1 497
0 499 7 1 2 998 498
0 500 5 1 1 499
0 501 7 2 2 999 1002
0 502 5 1 1 1167
0 503 7 1 2 1130 1168
0 504 5 1 1 503
0 505 7 1 2 1010 504
0 506 5 1 1 505
0 507 7 3 2 1021 1024
0 508 5 2 1 1169
0 509 7 1 2 1124 1170
0 510 5 1 1 509
0 511 7 1 2 1126 1172
0 512 5 1 1 511
0 513 7 2 2 1031 1035
0 514 5 2 1 1174
0 515 7 1 2 1122 1176
0 516 5 1 1 515
0 517 7 1 2 1120 1175
0 518 5 1 1 517
0 519 7 3 2 1042 1046
0 520 5 2 1 1178
0 521 7 1 2 1053 1181
0 522 5 1 1 521
0 523 7 1 2 425 1179
0 524 5 1 1 523
0 525 7 1 2 1054 1058
0 526 5 1 1 525
0 527 7 1 2 1071 1114
0 528 5 1 1 527
0 529 7 1 2 526 528
0 530 5 1 1 529
0 531 7 1 2 1066 1116
0 532 5 1 1 531
0 533 7 3 2 1080 1083
0 534 5 2 1 1183
0 535 7 1 2 1112 1184
0 536 5 1 1 535
0 537 7 1 2 1090 1094
0 538 5 2 1 537
0 539 7 1 2 1107 1188
0 540 5 2 1 539
0 541 7 1 2 82 1105
0 542 5 1 1 541
0 543 7 1 2 1101 542
0 544 5 2 1 543
0 545 7 1 2 1189 1192
0 546 5 1 1 545
0 547 7 1 2 1109 546
0 548 5 1 1 547
0 549 7 1 2 1190 548
0 550 5 1 1 549
0 551 7 1 2 414 1186
0 552 5 1 1 551
0 553 7 1 2 550 552
0 554 7 1 2 536 553
0 555 5 1 1 554
0 556 7 1 2 532 555
0 557 7 1 2 530 556
0 558 7 1 2 524 557
0 559 7 1 2 522 558
0 560 7 1 2 518 559
0 561 7 1 2 516 560
0 562 7 1 2 512 561
0 563 7 1 2 510 562
0 564 5 1 1 563
0 565 7 2 2 1011 1014
0 566 5 2 1 1194
0 567 7 1 2 1128 1196
0 568 5 1 1 567
0 569 7 1 2 564 568
0 570 7 1 2 506 569
0 571 7 1 2 500 570
0 572 7 1 2 495 571
0 573 7 1 2 491 572
0 574 7 1 2 485 573
0 575 7 1 2 479 574
0 576 7 1 2 477 575
0 577 7 1 2 473 576
0 578 7 1 2 1149 577
0 579 5 1 1 578
0 580 7 1 2 1095 1103
0 581 7 1 2 1193 580
0 582 5 1 1 581
0 583 7 1 2 1091 582
0 584 5 2 1 583
0 585 7 1 2 1081 1198
0 586 5 1 1 585
0 587 7 2 2 1084 586
0 588 5 2 1 1200
0 589 7 1 2 1069 1202
0 590 5 1 1 589
0 591 7 1 2 1074 590
0 592 7 1 2 1055 591
0 593 5 1 1 592
0 594 7 1 2 1059 593
0 595 7 1 2 1043 594
0 596 5 1 1 595
0 597 7 1 2 1047 596
0 598 7 2 2 1036 597
0 599 5 1 1 1204
0 600 7 2 2 1032 599
0 601 5 2 1 1206
0 602 7 1 2 1025 1208
0 603 5 1 1 602
0 604 7 2 2 1022 603
0 605 5 2 1 1210
0 606 7 1 2 1015 1212
0 607 5 1 1 606
0 608 7 2 2 1012 607
0 609 5 1 1 1214
0 610 7 1 2 1000 1215
0 611 5 2 1 610
0 612 7 1 2 1003 1216
0 613 5 1 1 612
0 614 7 1 2 992 613
0 615 5 1 1 614
0 616 7 2 2 1135 615
0 617 5 1 1 1218
0 618 7 1 2 984 1219
0 619 5 1 1 618
0 620 7 2 2 981 619
0 621 5 2 1 1220
0 622 7 1 2 973 1222
0 623 5 1 1 622
0 624 7 2 2 970 623
0 625 5 2 1 1224
0 626 7 1 2 962 1226
0 627 5 1 1 626
0 628 7 2 2 959 627
0 629 5 2 1 1228
0 630 7 1 2 1152 1230
0 631 5 1 1 630
0 632 7 1 2 1154 1229
0 633 5 1 1 632
0 634 7 1 2 631 633
0 635 5 1 1 634
0 636 7 1 2 1160 1221
0 637 5 1 1 636
0 638 7 1 2 487 1223
0 639 5 1 1 638
0 640 7 1 2 1162 617
0 641 5 1 1 640
0 642 7 1 2 1136 1164
0 643 5 1 1 642
0 644 7 1 2 1166 1217
0 645 5 1 1 644
0 646 7 1 2 1004 645
0 647 5 1 1 646
0 648 7 1 2 502 609
0 649 5 1 1 648
0 650 7 1 2 1195 1213
0 651 5 1 1 650
0 652 7 1 2 1197 1211
0 653 5 1 1 652
0 654 7 1 2 651 653
0 655 5 1 1 654
0 656 7 1 2 1171 1209
0 657 5 1 1 656
0 658 7 1 2 1173 1207
0 659 5 1 1 658
0 660 7 1 2 1044 1177
0 661 5 1 1 660
0 662 7 1 2 1033 1205
0 663 5 1 1 662
0 664 7 1 2 1056 1180
0 665 5 1 1 664
0 666 7 1 2 1067 1201
0 667 5 1 1 666
0 668 7 1 2 665 667
0 669 5 1 1 668
0 670 7 1 2 1060 1182
0 671 5 1 1 670
0 672 7 1 2 1072 1203
0 673 5 1 1 672
0 674 7 1 2 1092 1187
0 675 5 1 1 674
0 676 7 1 2 1185 1199
0 677 5 1 1 676
0 678 7 1 2 1191 677
0 679 7 1 2 675 678
0 680 5 1 1 679
0 681 7 1 2 673 680
0 682 7 1 2 671 681
0 683 7 1 2 669 682
0 684 7 1 2 663 683
0 685 7 1 2 661 684
0 686 7 1 2 659 685
0 687 7 1 2 657 686
0 688 5 1 1 687
0 689 7 1 2 655 688
0 690 7 1 2 649 689
0 691 7 1 2 647 690
0 692 7 1 2 643 691
0 693 7 1 2 641 692
0 694 7 1 2 639 693
0 695 7 1 2 637 694
0 696 7 1 2 944 695
0 697 7 1 2 481 1227
0 698 5 1 1 697
0 699 7 1 2 1157 1225
0 700 5 1 1 699
0 701 7 1 2 698 700
0 702 7 1 2 696 701
0 703 7 1 2 635 702
0 704 7 1 2 1145 1231
0 705 5 1 1 704
0 706 7 2 2 951 705
0 707 5 1 1 1232
0 708 7 1 2 938 707
0 709 5 1 1 708
0 710 7 1 2 940 1233
0 711 5 1 1 710
0 712 7 1 2 709 711
0 713 7 1 2 703 712
0 714 7 1 2 471 713
0 715 5 1 1 714
0 716 7 1 2 579 715
3 3499 5 0 1 716
