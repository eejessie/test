1 0 0 3 0
2 49 1 0
2 1829 1 0
2 1830 1 0
1 1 0 3 0
2 1831 1 1
2 1832 1 1
2 1833 1 1
1 2 0 3 0
2 1834 1 2
2 1835 1 2
2 1836 1 2
1 3 0 3 0
2 1837 1 3
2 1838 1 3
2 1839 1 3
1 4 0 3 0
2 1840 1 4
2 1841 1 4
2 1842 1 4
1 5 0 3 0
2 1843 1 5
2 1844 1 5
2 1845 1 5
1 6 0 3 0
2 1846 1 6
2 1847 1 6
2 1848 1 6
1 7 0 3 0
2 1849 1 7
2 1850 1 7
2 1851 1 7
1 8 0 3 0
2 1852 1 8
2 1853 1 8
2 1854 1 8
1 9 0 3 0
2 1855 1 9
2 1856 1 9
2 1857 1 9
1 10 0 3 0
2 1858 1 10
2 1859 1 10
2 1860 1 10
1 11 0 3 0
2 1861 1 11
2 1862 1 11
2 1863 1 11
1 12 0 3 0
2 1864 1 12
2 1865 1 12
2 1866 1 12
1 13 0 3 0
2 1867 1 13
2 1868 1 13
2 1869 1 13
1 14 0 3 0
2 1870 1 14
2 1871 1 14
2 1872 1 14
1 15 0 3 0
2 1873 1 15
2 1874 1 15
2 1875 1 15
1 16 0 3 0
2 1876 1 16
2 1877 1 16
2 1878 1 16
1 17 0 3 0
2 1879 1 17
2 1880 1 17
2 1881 1 17
1 18 0 3 0
2 1882 1 18
2 1883 1 18
2 1884 1 18
1 19 0 3 0
2 1885 1 19
2 1886 1 19
2 1887 1 19
1 20 0 3 0
2 1888 1 20
2 1889 1 20
2 1890 1 20
1 21 0 3 0
2 1891 1 21
2 1892 1 21
2 1893 1 21
1 22 0 3 0
2 1894 1 22
2 1895 1 22
2 1896 1 22
1 23 0 3 0
2 1897 1 23
2 1898 1 23
2 1899 1 23
1 24 0 3 0
2 1900 1 24
2 1901 1 24
2 1902 1 24
1 25 0 3 0
2 1903 1 25
2 1904 1 25
2 1905 1 25
1 26 0 3 0
2 1906 1 26
2 1907 1 26
2 1908 1 26
1 27 0 3 0
2 1909 1 27
2 1910 1 27
2 1911 1 27
1 28 0 3 0
2 1912 1 28
2 1913 1 28
2 1914 1 28
1 29 0 3 0
2 1915 1 29
2 1916 1 29
2 1917 1 29
1 30 0 3 0
2 1918 1 30
2 1919 1 30
2 1920 1 30
1 31 0 3 0
2 1921 1 31
2 1922 1 31
2 1923 1 31
1 32 0 3 0
2 1924 1 32
2 1925 1 32
2 1926 1 32
1 33 0 3 0
2 1927 1 33
2 1928 1 33
2 1929 1 33
1 34 0 3 0
2 1930 1 34
2 1931 1 34
2 1932 1 34
1 35 0 3 0
2 1933 1 35
2 1934 1 35
2 1935 1 35
1 36 0 3 0
2 1936 1 36
2 1937 1 36
2 1938 1 36
1 37 0 3 0
2 1939 1 37
2 1940 1 37
2 1941 1 37
1 38 0 3 0
2 1942 1 38
2 1943 1 38
2 1944 1 38
1 39 0 3 0
2 1945 1 39
2 1946 1 39
2 1947 1 39
1 40 0 3 0
2 1948 1 40
2 1949 1 40
2 1950 1 40
1 41 0 3 0
2 1951 1 41
2 1952 1 41
2 1953 1 41
1 42 0 3 0
2 1954 1 42
2 1955 1 42
2 1956 1 42
1 43 0 3 0
2 1957 1 43
2 1958 1 43
2 1959 1 43
1 44 0 3 0
2 1960 1 44
2 1961 1 44
2 1962 1 44
1 45 0 4 0
2 1963 1 45
2 1964 1 45
2 1965 1 45
2 1966 1 45
1 46 0 3 0
2 1967 1 46
2 1968 1 46
2 1969 1 46
1 47 0 4 0
2 1970 1 47
2 1971 1 47
2 1972 1 47
2 1973 1 47
1 48 0 4 0
2 1974 1 48
2 1975 1 48
2 1976 1 48
2 1977 1 48
2 1978 1 50
2 1979 1 50
2 1980 1 51
2 1981 1 51
2 1982 1 51
2 1983 1 52
2 1984 1 52
2 1985 1 52
2 1986 1 53
2 1987 1 53
2 1988 1 53
2 1989 1 54
2 1990 1 54
2 1991 1 54
2 1992 1 55
2 1993 1 55
2 1994 1 55
2 1995 1 56
2 1996 1 56
2 1997 1 56
2 1998 1 57
2 1999 1 57
2 2000 1 57
2 2001 1 58
2 2002 1 58
2 2003 1 58
2 2004 1 59
2 2005 1 59
2 2006 1 59
2 2007 1 60
2 2008 1 60
2 2009 1 60
2 2010 1 61
2 2011 1 61
2 2012 1 61
2 2013 1 62
2 2014 1 62
2 2015 1 62
2 2016 1 63
2 2017 1 63
2 2018 1 63
2 2019 1 64
2 2020 1 64
2 2021 1 64
2 2022 1 65
2 2023 1 65
2 2024 1 65
2 2025 1 66
2 2026 1 66
2 2027 1 66
2 2028 1 67
2 2029 1 67
2 2030 1 67
2 2031 1 68
2 2032 1 68
2 2033 1 68
2 2034 1 69
2 2035 1 69
2 2036 1 69
2 2037 1 69
2 2038 1 70
2 2039 1 70
2 2040 1 70
2 2041 1 70
2 2042 1 71
2 2043 1 71
2 2044 1 71
2 2045 1 71
2 2046 1 72
2 2047 1 72
2 2048 1 72
2 2049 1 72
2 2050 1 73
2 2051 1 73
2 2052 1 73
2 2053 1 73
2 2054 1 74
2 2055 1 74
2 2056 1 74
2 2057 1 74
2 2058 1 75
2 2059 1 75
2 2060 1 75
2 2061 1 75
2 2062 1 76
2 2063 1 76
2 2064 1 76
2 2065 1 76
2 2066 1 77
2 2067 1 77
2 2068 1 77
2 2069 1 77
2 2070 1 78
2 2071 1 78
2 2072 1 78
2 2073 1 78
2 2074 1 79
2 2075 1 79
2 2076 1 79
2 2077 1 79
2 2078 1 80
2 2079 1 80
2 2080 1 80
2 2081 1 80
2 2082 1 81
2 2083 1 81
2 2084 1 81
2 2085 1 81
2 2086 1 82
2 2087 1 82
2 2088 1 82
2 2089 1 83
2 2090 1 83
2 2091 1 83
2 2092 1 84
2 2093 1 84
2 2094 1 84
2 2095 1 85
2 2096 1 85
2 2097 1 85
2 2098 1 86
2 2099 1 86
2 2100 1 86
2 2101 1 87
2 2102 1 87
2 2103 1 87
2 2104 1 88
2 2105 1 88
2 2106 1 88
2 2107 1 89
2 2108 1 89
2 2109 1 89
2 2110 1 90
2 2111 1 90
2 2112 1 90
2 2113 1 91
2 2114 1 91
2 2115 1 91
2 2116 1 92
2 2117 1 92
2 2118 1 92
2 2119 1 93
2 2120 1 93
2 2121 1 93
2 2122 1 94
2 2123 1 94
2 2124 1 94
2 2125 1 95
2 2126 1 95
2 2127 1 95
2 2128 1 95
2 2129 1 96
2 2130 1 96
2 2131 1 96
2 2132 1 97
2 2133 1 97
2 2134 1 98
2 2135 1 98
2 2136 1 99
2 2137 1 99
2 2138 1 101
2 2139 1 101
2 2140 1 107
2 2141 1 107
2 2142 1 109
2 2143 1 109
2 2144 1 113
2 2145 1 113
2 2146 1 113
2 2147 1 117
2 2148 1 117
2 2149 1 118
2 2150 1 118
2 2151 1 122
2 2152 1 122
2 2153 1 125
2 2154 1 125
2 2155 1 128
2 2156 1 128
2 2157 1 130
2 2158 1 130
2 2159 1 131
2 2160 1 131
2 2161 1 136
2 2162 1 136
2 2163 1 139
2 2164 1 139
2 2165 1 140
2 2166 1 140
2 2167 1 143
2 2168 1 143
2 2169 1 146
2 2170 1 146
2 2171 1 148
2 2172 1 148
2 2173 1 149
2 2174 1 149
2 2175 1 154
2 2176 1 154
2 2177 1 157
2 2178 1 157
2 2179 1 162
2 2180 1 162
2 2181 1 162
2 2182 1 168
2 2183 1 168
2 2184 1 168
2 2185 1 170
2 2186 1 170
2 2187 1 173
2 2188 1 173
2 2189 1 176
2 2190 1 176
2 2191 1 178
2 2192 1 178
2 2193 1 179
2 2194 1 179
2 2195 1 184
2 2196 1 184
2 2197 1 187
2 2198 1 187
2 2199 1 188
2 2200 1 188
2 2201 1 191
2 2202 1 191
2 2203 1 194
2 2204 1 194
2 2205 1 196
2 2206 1 196
2 2207 1 197
2 2208 1 197
2 2209 1 202
2 2210 1 202
2 2211 1 205
2 2212 1 205
2 2213 1 210
2 2214 1 210
2 2215 1 210
2 2216 1 216
2 2217 1 216
2 2218 1 216
2 2219 1 218
2 2220 1 218
2 2221 1 221
2 2222 1 221
2 2223 1 224
2 2224 1 224
2 2225 1 226
2 2226 1 226
2 2227 1 227
2 2228 1 227
2 2229 1 232
2 2230 1 232
2 2231 1 235
2 2232 1 235
2 2233 1 236
2 2234 1 236
2 2235 1 239
2 2236 1 239
2 2237 1 242
2 2238 1 242
2 2239 1 244
2 2240 1 244
2 2241 1 245
2 2242 1 245
2 2243 1 250
2 2244 1 250
2 2245 1 253
2 2246 1 253
2 2247 1 258
2 2248 1 258
2 2249 1 258
2 2250 1 264
2 2251 1 264
2 2252 1 264
2 2253 1 266
2 2254 1 266
2 2255 1 269
2 2256 1 269
2 2257 1 272
2 2258 1 272
2 2259 1 274
2 2260 1 274
2 2261 1 275
2 2262 1 275
2 2263 1 280
2 2264 1 280
2 2265 1 283
2 2266 1 283
2 2267 1 284
2 2268 1 284
2 2269 1 287
2 2270 1 287
2 2271 1 290
2 2272 1 290
2 2273 1 292
2 2274 1 292
2 2275 1 293
2 2276 1 293
2 2277 1 298
2 2278 1 298
2 2279 1 301
2 2280 1 301
2 2281 1 306
2 2282 1 306
2 2283 1 306
2 2284 1 312
2 2285 1 312
2 2286 1 312
2 2287 1 314
2 2288 1 314
2 2289 1 317
2 2290 1 317
2 2291 1 320
2 2292 1 320
2 2293 1 322
2 2294 1 322
2 2295 1 323
2 2296 1 323
2 2297 1 328
2 2298 1 328
2 2299 1 331
2 2300 1 331
2 2301 1 332
2 2302 1 332
2 2303 1 335
2 2304 1 335
2 2305 1 338
2 2306 1 338
2 2307 1 340
2 2308 1 340
2 2309 1 341
2 2310 1 341
2 2311 1 346
2 2312 1 346
2 2313 1 349
2 2314 1 349
2 2315 1 354
2 2316 1 354
2 2317 1 354
2 2318 1 360
2 2319 1 360
2 2320 1 360
2 2321 1 362
2 2322 1 362
2 2323 1 365
2 2324 1 365
2 2325 1 368
2 2326 1 368
2 2327 1 370
2 2328 1 370
2 2329 1 371
2 2330 1 371
2 2331 1 376
2 2332 1 376
2 2333 1 379
2 2334 1 379
2 2335 1 380
2 2336 1 380
2 2337 1 383
2 2338 1 383
2 2339 1 386
2 2340 1 386
2 2341 1 388
2 2342 1 388
2 2343 1 389
2 2344 1 389
2 2345 1 394
2 2346 1 394
2 2347 1 397
2 2348 1 397
2 2349 1 402
2 2350 1 402
2 2351 1 402
2 2352 1 408
2 2353 1 408
2 2354 1 408
2 2355 1 410
2 2356 1 410
2 2357 1 413
2 2358 1 413
2 2359 1 416
2 2360 1 416
2 2361 1 418
2 2362 1 418
2 2363 1 419
2 2364 1 419
2 2365 1 424
2 2366 1 424
2 2367 1 427
2 2368 1 427
2 2369 1 428
2 2370 1 428
2 2371 1 431
2 2372 1 431
2 2373 1 434
2 2374 1 434
2 2375 1 436
2 2376 1 436
2 2377 1 437
2 2378 1 437
2 2379 1 442
2 2380 1 442
2 2381 1 445
2 2382 1 445
2 2383 1 450
2 2384 1 450
2 2385 1 450
2 2386 1 456
2 2387 1 456
2 2388 1 456
2 2389 1 458
2 2390 1 458
2 2391 1 461
2 2392 1 461
2 2393 1 464
2 2394 1 464
2 2395 1 466
2 2396 1 466
2 2397 1 467
2 2398 1 467
2 2399 1 472
2 2400 1 472
2 2401 1 475
2 2402 1 475
2 2403 1 476
2 2404 1 476
2 2405 1 479
2 2406 1 479
2 2407 1 482
2 2408 1 482
2 2409 1 484
2 2410 1 484
2 2411 1 485
2 2412 1 485
2 2413 1 490
2 2414 1 490
2 2415 1 493
2 2416 1 493
2 2417 1 498
2 2418 1 498
2 2419 1 498
2 2420 1 504
2 2421 1 504
2 2422 1 504
2 2423 1 506
2 2424 1 506
2 2425 1 509
2 2426 1 509
2 2427 1 512
2 2428 1 512
2 2429 1 514
2 2430 1 514
2 2431 1 515
2 2432 1 515
2 2433 1 520
2 2434 1 520
2 2435 1 523
2 2436 1 523
2 2437 1 524
2 2438 1 524
2 2439 1 527
2 2440 1 527
2 2441 1 530
2 2442 1 530
2 2443 1 532
2 2444 1 532
2 2445 1 533
2 2446 1 533
2 2447 1 538
2 2448 1 538
2 2449 1 541
2 2450 1 541
2 2451 1 546
2 2452 1 546
2 2453 1 546
2 2454 1 552
2 2455 1 552
2 2456 1 552
2 2457 1 554
2 2458 1 554
2 2459 1 557
2 2460 1 557
2 2461 1 560
2 2462 1 560
2 2463 1 562
2 2464 1 562
2 2465 1 563
2 2466 1 563
2 2467 1 568
2 2468 1 568
2 2469 1 571
2 2470 1 571
2 2471 1 572
2 2472 1 572
2 2473 1 575
2 2474 1 575
2 2475 1 578
2 2476 1 578
2 2477 1 580
2 2478 1 580
2 2479 1 581
2 2480 1 581
2 2481 1 586
2 2482 1 586
2 2483 1 589
2 2484 1 589
2 2485 1 594
2 2486 1 594
2 2487 1 594
2 2488 1 600
2 2489 1 600
2 2490 1 600
2 2491 1 602
2 2492 1 602
2 2493 1 605
2 2494 1 605
2 2495 1 608
2 2496 1 608
2 2497 1 610
2 2498 1 610
2 2499 1 611
2 2500 1 611
2 2501 1 616
2 2502 1 616
2 2503 1 619
2 2504 1 619
2 2505 1 620
2 2506 1 620
2 2507 1 623
2 2508 1 623
2 2509 1 626
2 2510 1 626
2 2511 1 628
2 2512 1 628
2 2513 1 629
2 2514 1 629
2 2515 1 634
2 2516 1 634
2 2517 1 637
2 2518 1 637
2 2519 1 642
2 2520 1 642
2 2521 1 642
2 2522 1 648
2 2523 1 648
2 2524 1 648
2 2525 1 650
2 2526 1 650
2 2527 1 653
2 2528 1 653
2 2529 1 656
2 2530 1 656
2 2531 1 658
2 2532 1 658
2 2533 1 659
2 2534 1 659
2 2535 1 664
2 2536 1 664
2 2537 1 667
2 2538 1 667
2 2539 1 668
2 2540 1 668
2 2541 1 671
2 2542 1 671
2 2543 1 674
2 2544 1 674
2 2545 1 676
2 2546 1 676
2 2547 1 677
2 2548 1 677
2 2549 1 682
2 2550 1 682
2 2551 1 685
2 2552 1 685
2 2553 1 690
2 2554 1 690
2 2555 1 690
2 2556 1 696
2 2557 1 696
2 2558 1 696
2 2559 1 698
2 2560 1 698
2 2561 1 701
2 2562 1 701
2 2563 1 704
2 2564 1 704
2 2565 1 706
2 2566 1 706
2 2567 1 707
2 2568 1 707
2 2569 1 712
2 2570 1 712
2 2571 1 715
2 2572 1 715
2 2573 1 716
2 2574 1 716
2 2575 1 719
2 2576 1 719
2 2577 1 722
2 2578 1 722
2 2579 1 724
2 2580 1 724
2 2581 1 725
2 2582 1 725
2 2583 1 730
2 2584 1 730
2 2585 1 733
2 2586 1 733
2 2587 1 738
2 2588 1 738
2 2589 1 738
2 2590 1 744
2 2591 1 744
2 2592 1 744
2 2593 1 746
2 2594 1 746
2 2595 1 749
2 2596 1 749
2 2597 1 752
2 2598 1 752
2 2599 1 754
2 2600 1 754
2 2601 1 755
2 2602 1 755
2 2603 1 760
2 2604 1 760
2 2605 1 763
2 2606 1 763
2 2607 1 764
2 2608 1 764
2 2609 1 767
2 2610 1 767
2 2611 1 770
2 2612 1 770
2 2613 1 772
2 2614 1 772
2 2615 1 773
2 2616 1 773
2 2617 1 778
2 2618 1 778
2 2619 1 781
2 2620 1 781
2 2621 1 786
2 2622 1 786
2 2623 1 786
2 2624 1 792
2 2625 1 792
2 2626 1 792
2 2627 1 794
2 2628 1 794
2 2629 1 797
2 2630 1 797
2 2631 1 800
2 2632 1 800
2 2633 1 802
2 2634 1 802
2 2635 1 803
2 2636 1 803
2 2637 1 808
2 2638 1 808
2 2639 1 811
2 2640 1 811
2 2641 1 812
2 2642 1 812
2 2643 1 815
2 2644 1 815
2 2645 1 818
2 2646 1 818
2 2647 1 820
2 2648 1 820
2 2649 1 821
2 2650 1 821
2 2651 1 826
2 2652 1 826
2 2653 1 829
2 2654 1 829
2 2655 1 834
2 2656 1 834
2 2657 1 834
2 2658 1 840
2 2659 1 840
2 2660 1 840
2 2661 1 842
2 2662 1 842
2 2663 1 845
2 2664 1 845
2 2665 1 848
2 2666 1 848
2 2667 1 850
2 2668 1 850
2 2669 1 851
2 2670 1 851
2 2671 1 856
2 2672 1 856
2 2673 1 859
2 2674 1 859
2 2675 1 860
2 2676 1 860
2 2677 1 863
2 2678 1 863
2 2679 1 866
2 2680 1 866
2 2681 1 868
2 2682 1 868
2 2683 1 869
2 2684 1 869
2 2685 1 874
2 2686 1 874
2 2687 1 877
2 2688 1 877
2 2689 1 882
2 2690 1 882
2 2691 1 882
2 2692 1 888
2 2693 1 888
2 2694 1 888
2 2695 1 890
2 2696 1 890
2 2697 1 893
2 2698 1 893
2 2699 1 896
2 2700 1 896
2 2701 1 898
2 2702 1 898
2 2703 1 899
2 2704 1 899
2 2705 1 904
2 2706 1 904
2 2707 1 907
2 2708 1 907
2 2709 1 908
2 2710 1 908
2 2711 1 911
2 2712 1 911
2 2713 1 914
2 2714 1 914
2 2715 1 916
2 2716 1 916
2 2717 1 917
2 2718 1 917
2 2719 1 922
2 2720 1 922
2 2721 1 925
2 2722 1 925
2 2723 1 930
2 2724 1 930
2 2725 1 930
2 2726 1 936
2 2727 1 936
2 2728 1 936
2 2729 1 938
2 2730 1 938
2 2731 1 941
2 2732 1 941
2 2733 1 944
2 2734 1 944
2 2735 1 946
2 2736 1 946
2 2737 1 947
2 2738 1 947
2 2739 1 952
2 2740 1 952
2 2741 1 955
2 2742 1 955
2 2743 1 956
2 2744 1 956
2 2745 1 959
2 2746 1 959
2 2747 1 962
2 2748 1 962
2 2749 1 964
2 2750 1 964
2 2751 1 965
2 2752 1 965
2 2753 1 970
2 2754 1 970
2 2755 1 973
2 2756 1 973
2 2757 1 978
2 2758 1 978
2 2759 1 978
2 2760 1 984
2 2761 1 984
2 2762 1 984
2 2763 1 986
2 2764 1 986
2 2765 1 989
2 2766 1 989
2 2767 1 992
2 2768 1 992
2 2769 1 994
2 2770 1 994
2 2771 1 995
2 2772 1 995
2 2773 1 1000
2 2774 1 1000
2 2775 1 1003
2 2776 1 1003
2 2777 1 1004
2 2778 1 1004
2 2779 1 1007
2 2780 1 1007
2 2781 1 1010
2 2782 1 1010
2 2783 1 1012
2 2784 1 1012
2 2785 1 1013
2 2786 1 1013
2 2787 1 1018
2 2788 1 1018
2 2789 1 1021
2 2790 1 1021
2 2791 1 1026
2 2792 1 1026
2 2793 1 1026
2 2794 1 1032
2 2795 1 1032
2 2796 1 1032
2 2797 1 1034
2 2798 1 1034
2 2799 1 1037
2 2800 1 1037
2 2801 1 1040
2 2802 1 1040
2 2803 1 1042
2 2804 1 1042
2 2805 1 1043
2 2806 1 1043
2 2807 1 1048
2 2808 1 1048
2 2809 1 1051
2 2810 1 1051
2 2811 1 1052
2 2812 1 1052
2 2813 1 1055
2 2814 1 1055
2 2815 1 1058
2 2816 1 1058
2 2817 1 1060
2 2818 1 1060
2 2819 1 1061
2 2820 1 1061
2 2821 1 1066
2 2822 1 1066
2 2823 1 1069
2 2824 1 1069
2 2825 1 1074
2 2826 1 1074
2 2827 1 1074
2 2828 1 1080
2 2829 1 1080
2 2830 1 1080
2 2831 1 1082
2 2832 1 1082
2 2833 1 1085
2 2834 1 1085
2 2835 1 1088
2 2836 1 1088
2 2837 1 1090
2 2838 1 1090
2 2839 1 1091
2 2840 1 1091
2 2841 1 1096
2 2842 1 1096
2 2843 1 1099
2 2844 1 1099
2 2845 1 1100
2 2846 1 1100
2 2847 1 1103
2 2848 1 1103
2 2849 1 1106
2 2850 1 1106
2 2851 1 1108
2 2852 1 1108
2 2853 1 1109
2 2854 1 1109
2 2855 1 1114
2 2856 1 1114
2 2857 1 1117
2 2858 1 1117
2 2859 1 1122
2 2860 1 1122
2 2861 1 1122
2 2862 1 1128
2 2863 1 1128
2 2864 1 1128
2 2865 1 1130
2 2866 1 1130
2 2867 1 1133
2 2868 1 1133
2 2869 1 1136
2 2870 1 1136
2 2871 1 1138
2 2872 1 1138
2 2873 1 1139
2 2874 1 1139
2 2875 1 1144
2 2876 1 1144
2 2877 1 1147
2 2878 1 1147
2 2879 1 1148
2 2880 1 1148
2 2881 1 1151
2 2882 1 1151
2 2883 1 1154
2 2884 1 1154
2 2885 1 1156
2 2886 1 1156
2 2887 1 1162
2 2888 1 1162
2 2889 1 1165
2 2890 1 1165
2 2891 1 1170
2 2892 1 1170
2 2893 1 1171
2 2894 1 1171
2 2895 1 1175
2 2896 1 1175
2 2897 1 1176
2 2898 1 1176
2 2899 1 1180
2 2900 1 1180
2 2901 1 1183
2 2902 1 1183
2 2903 1 1198
2 2904 1 1198
2 2905 1 1201
2 2906 1 1201
2 2907 1 1203
2 2908 1 1203
2 2909 1 1205
2 2910 1 1205
2 2911 1 1207
2 2912 1 1207
2 2913 1 1208
2 2914 1 1208
2 2915 1 1209
2 2916 1 1209
2 2917 1 1209
2 2918 1 1212
2 2919 1 1212
2 2920 1 1213
2 2921 1 1213
2 2922 1 1216
2 2923 1 1216
2 2924 1 1219
2 2925 1 1219
2 2926 1 1221
2 2927 1 1221
2 2928 1 1224
2 2929 1 1224
2 2930 1 1227
2 2931 1 1227
2 2932 1 1229
2 2933 1 1229
2 2934 1 1232
2 2935 1 1232
2 2936 1 1235
2 2937 1 1235
2 2938 1 1237
2 2939 1 1237
2 2940 1 1240
2 2941 1 1240
2 2942 1 1243
2 2943 1 1243
2 2944 1 1245
2 2945 1 1245
2 2946 1 1248
2 2947 1 1248
2 2948 1 1251
2 2949 1 1251
2 2950 1 1253
2 2951 1 1253
2 2952 1 1256
2 2953 1 1256
2 2954 1 1259
2 2955 1 1259
2 2956 1 1261
2 2957 1 1261
2 2958 1 1264
2 2959 1 1264
2 2960 1 1267
2 2961 1 1267
2 2962 1 1269
2 2963 1 1269
2 2964 1 1272
2 2965 1 1272
2 2966 1 1275
2 2967 1 1275
2 2968 1 1277
2 2969 1 1277
2 2970 1 1280
2 2971 1 1280
2 2972 1 1283
2 2973 1 1283
2 2974 1 1285
2 2975 1 1285
2 2976 1 1288
2 2977 1 1288
2 2978 1 1291
2 2979 1 1291
2 2980 1 1293
2 2981 1 1293
2 2982 1 1296
2 2983 1 1296
2 2984 1 1299
2 2985 1 1299
2 2986 1 1301
2 2987 1 1301
2 2988 1 1304
2 2989 1 1304
2 2990 1 1307
2 2991 1 1307
2 2992 1 1309
2 2993 1 1309
2 2994 1 1312
2 2995 1 1312
2 2996 1 1315
2 2997 1 1315
2 2998 1 1317
2 2999 1 1317
2 3000 1 1318
2 3001 1 1318
2 3002 1 1324
2 3003 1 1324
2 3004 1 1327
2 3005 1 1327
2 3006 1 1327
2 3007 1 1330
2 3008 1 1330
2 3009 1 1333
2 3010 1 1333
2 3011 1 1333
2 3012 1 1335
2 3013 1 1335
2 3014 1 1335
2 3015 1 1335
2 3016 1 1336
2 3017 1 1336
2 3018 1 1342
2 3019 1 1342
2 3020 1 1345
2 3021 1 1345
2 3022 1 1345
2 3023 1 1347
2 3024 1 1347
2 3025 1 1347
2 3026 1 1347
2 3027 1 1348
2 3028 1 1348
2 3029 1 1354
2 3030 1 1354
2 3031 1 1357
2 3032 1 1357
2 3033 1 1357
2 3034 1 1359
2 3035 1 1359
2 3036 1 1359
2 3037 1 1359
2 3038 1 1359
2 3039 1 1360
2 3040 1 1360
2 3041 1 1366
2 3042 1 1366
2 3043 1 1369
2 3044 1 1369
2 3045 1 1369
2 3046 1 1371
2 3047 1 1371
2 3048 1 1371
2 3049 1 1371
2 3050 1 1371
2 3051 1 1372
2 3052 1 1372
2 3053 1 1378
2 3054 1 1378
2 3055 1 1381
2 3056 1 1381
2 3057 1 1381
2 3058 1 1381
2 3059 1 1382
2 3060 1 1382
2 3061 1 1388
2 3062 1 1388
2 3063 1 1391
2 3064 1 1391
2 3065 1 1391
2 3066 1 1393
2 3067 1 1393
2 3068 1 1393
2 3069 1 1393
2 3070 1 1394
2 3071 1 1394
2 3072 1 1400
2 3073 1 1400
2 3074 1 1403
2 3075 1 1403
2 3076 1 1403
2 3077 1 1403
2 3078 1 1405
2 3079 1 1405
2 3080 1 1405
2 3081 1 1406
2 3082 1 1406
2 3083 1 1412
2 3084 1 1412
2 3085 1 1415
2 3086 1 1415
2 3087 1 1415
2 3088 1 1415
2 3089 1 1417
2 3090 1 1417
2 3091 1 1417
2 3092 1 1418
2 3093 1 1418
2 3094 1 1424
2 3095 1 1424
2 3096 1 1427
2 3097 1 1427
2 3098 1 1427
2 3099 1 1427
2 3100 1 1429
2 3101 1 1429
2 3102 1 1429
2 3103 1 1429
2 3104 1 1430
2 3105 1 1430
2 3106 1 1436
2 3107 1 1436
2 3108 1 1439
2 3109 1 1439
2 3110 1 1439
2 3111 1 1439
2 3112 1 1439
2 3113 1 1441
2 3114 1 1441
2 3115 1 1441
2 3116 1 1441
2 3117 1 1442
2 3118 1 1442
2 3119 1 1448
2 3120 1 1448
2 3121 1 1451
2 3122 1 1451
2 3123 1 1451
2 3124 1 1451
2 3125 1 1453
2 3126 1 1453
2 3127 1 1453
2 3128 1 1454
2 3129 1 1454
2 3130 1 1460
2 3131 1 1460
2 3132 1 1463
2 3133 1 1463
2 3134 1 1463
2 3135 1 1463
2 3136 1 1465
2 3137 1 1465
2 3138 1 1465
2 3139 1 1466
2 3140 1 1466
2 3141 1 1472
2 3142 1 1472
2 3143 1 1475
2 3144 1 1475
2 3145 1 1476
2 3146 1 1476
2 3147 1 1482
2 3148 1 1482
2 3149 1 1486
2 3150 1 1486
2 3151 1 1490
2 3152 1 1490
2 3153 1 1494
2 3154 1 1494
2 3155 1 1496
2 3156 1 1496
2 3157 1 1501
2 3158 1 1501
2 3159 1 1501
2 3160 1 1503
2 3161 1 1503
2 3162 1 1504
2 3163 1 1504
2 3164 1 1507
2 3165 1 1507
2 3166 1 1508
2 3167 1 1508
2 3168 1 1511
2 3169 1 1511
2 3170 1 1514
2 3171 1 1514
2 3172 1 1520
2 3173 1 1520
2 3174 1 1523
2 3175 1 1523
2 3176 1 1524
2 3177 1 1524
2 3178 1 1527
2 3179 1 1527
2 3180 1 1527
2 3181 1 1531
2 3182 1 1531
2 3183 1 1531
2 3184 1 1533
2 3185 1 1533
2 3186 1 1539
2 3187 1 1539
2 3188 1 1541
2 3189 1 1541
2 3190 1 1541
2 3191 1 1542
2 3192 1 1542
2 3193 1 1545
2 3194 1 1545
2 3195 1 1545
2 3196 1 1546
2 3197 1 1546
2 3198 1 1548
2 3199 1 1548
2 3200 1 1548
2 3201 1 1548
2 3202 1 1549
2 3203 1 1549
2 3204 1 1553
2 3205 1 1553
2 3206 1 1556
2 3207 1 1556
2 3208 1 1557
2 3209 1 1557
2 3210 1 1560
2 3211 1 1560
2 3212 1 1561
2 3213 1 1561
2 3214 1 1564
2 3215 1 1564
2 3216 1 1564
2 3217 1 1572
2 3218 1 1572
2 3219 1 1574
2 3220 1 1574
2 3221 1 1579
2 3222 1 1579
2 3223 1 1579
2 3224 1 1581
2 3225 1 1581
2 3226 1 1582
2 3227 1 1582
2 3228 1 1585
2 3229 1 1585
2 3230 1 1585
2 3231 1 1586
2 3232 1 1586
2 3233 1 1591
2 3234 1 1591
2 3235 1 1592
2 3236 1 1592
2 3237 1 1597
2 3238 1 1597
2 3239 1 1598
2 3240 1 1598
2 3241 1 1604
2 3242 1 1604
2 3243 1 1611
2 3244 1 1611
2 3245 1 1611
2 3246 1 1612
2 3247 1 1612
2 3248 1 1617
2 3249 1 1617
2 3250 1 1617
2 3251 1 1618
2 3252 1 1618
2 3253 1 1623
2 3254 1 1623
2 3255 1 1623
2 3256 1 1624
2 3257 1 1624
2 3258 1 1629
2 3259 1 1629
2 3260 1 1635
2 3261 1 1635
2 3262 1 1638
2 3263 1 1638
2 3264 1 1638
2 3265 1 1639
2 3266 1 1639
2 3267 1 1642
2 3268 1 1642
2 3269 1 1642
2 3270 1 1643
2 3271 1 1643
2 3272 1 1649
2 3273 1 1649
2 3274 1 1649
2 3275 1 1652
2 3276 1 1652
2 3277 1 1684
2 3278 1 1684
2 3279 1 1687
2 3280 1 1687
2 3281 1 1688
2 3282 1 1688
2 3283 1 1691
2 3284 1 1691
2 3285 1 1692
2 3286 1 1692
2 3287 1 1695
2 3288 1 1695
2 3289 1 1695
2 3290 1 1702
2 3291 1 1702
2 3292 1 1705
2 3293 1 1705
2 3294 1 1706
2 3295 1 1706
2 3296 1 1709
2 3297 1 1709
2 3298 1 1710
2 3299 1 1710
2 3300 1 1713
2 3301 1 1713
2 3302 1 1714
2 3303 1 1714
2 3304 1 1724
2 3305 1 1724
2 3306 1 1726
2 3307 1 1726
2 3308 1 1727
2 3309 1 1727
2 3310 1 1730
2 3311 1 1730
0 50 5 2 1 49
0 51 5 3 1 1831
0 52 5 3 1 1834
0 53 5 3 1 1837
0 54 5 3 1 1840
0 55 5 3 1 1843
0 56 5 3 1 1846
0 57 5 3 1 1849
0 58 5 3 1 1852
0 59 5 3 1 1855
0 60 5 3 1 1858
0 61 5 3 1 1861
0 62 5 3 1 1864
0 63 5 3 1 1867
0 64 5 3 1 1870
0 65 5 3 1 1873
0 66 5 3 1 1876
0 67 5 3 1 1879
0 68 5 3 1 1882
0 69 5 4 1 1885
0 70 5 4 1 1888
0 71 5 4 1 1891
0 72 5 4 1 1894
0 73 5 4 1 1897
0 74 5 4 1 1900
0 75 5 4 1 1903
0 76 5 4 1 1906
0 77 5 4 1 1909
0 78 5 4 1 1912
0 79 5 4 1 1915
0 80 5 4 1 1918
0 81 5 4 1 1921
0 82 5 3 1 1924
0 83 5 3 1 1927
0 84 5 3 1 1930
0 85 5 3 1 1933
0 86 5 3 1 1936
0 87 5 3 1 1939
0 88 5 3 1 1942
0 89 5 3 1 1945
0 90 5 3 1 1948
0 91 5 3 1 1951
0 92 5 3 1 1954
0 93 5 3 1 1957
0 94 5 3 1 1960
0 95 5 4 1 1963
0 96 5 3 1 1967
0 97 5 2 1 1970
0 98 5 2 1 1974
0 99 7 2 2 2129 2132
0 100 5 1 1 2136
0 101 7 2 2 2130 1975
0 102 5 1 1 2138
0 103 7 1 2 100 2139
0 104 5 1 1 103
0 105 7 1 2 1968 2134
0 106 5 1 1 105
0 107 7 2 2 104 106
0 108 5 1 1 2140
0 109 7 2 2 2125 2141
0 110 5 1 1 2142
0 111 7 1 2 1971 2143
0 112 5 1 1 111
0 113 7 3 2 1976 2137
0 114 5 1 1 2144
0 115 7 1 2 1964 2145
0 116 5 1 1 115
0 117 7 2 2 112 116
0 118 5 2 1 2147
0 119 7 1 2 1972 102
0 120 7 1 2 110 119
0 121 5 1 1 120
0 122 7 2 2 114 121
0 123 5 1 1 2151
0 124 7 1 2 2126 123
0 125 5 2 1 124
0 126 7 1 2 1965 2152
0 127 5 1 1 126
0 128 7 2 2 2153 127
0 129 5 1 1 2155
0 130 7 2 2 2122 2156
0 131 5 2 1 2157
0 132 7 1 2 108 2154
0 133 5 1 1 132
0 134 7 1 2 2127 2146
0 135 5 1 1 134
0 136 7 2 2 133 135
0 137 5 1 1 2161
0 138 7 1 2 2159 137
0 139 5 2 1 138
0 140 7 2 2 2148 2163
0 141 5 1 1 2165
0 142 7 1 2 2123 141
0 143 5 2 1 142
0 144 7 1 2 1961 2166
0 145 5 1 1 144
0 146 7 2 2 2167 145
0 147 5 1 1 2169
0 148 7 2 2 2119 2170
0 149 5 2 1 2171
0 150 7 1 2 129 2168
0 151 5 1 1 150
0 152 7 1 2 2149 2158
0 153 5 1 1 152
0 154 7 2 2 151 153
0 155 5 1 1 2175
0 156 7 1 2 2173 155
0 157 5 2 1 156
0 158 7 1 2 2150 2160
0 159 5 1 1 158
0 160 7 1 2 2162 159
0 161 5 1 1 160
0 162 7 3 2 2164 161
0 163 5 1 1 2179
0 164 7 1 2 2174 2180
0 165 5 1 1 164
0 166 7 1 2 2176 165
0 167 5 1 1 166
0 168 7 3 2 2177 167
0 169 5 1 1 2182
0 170 7 2 2 2178 163
0 171 5 1 1 2185
0 172 7 1 2 2120 171
0 173 5 2 1 172
0 174 7 1 2 1958 2186
0 175 5 1 1 174
0 176 7 2 2 2187 175
0 177 5 1 1 2189
0 178 7 2 2 2116 2190
0 179 5 2 1 2191
0 180 7 1 2 147 2188
0 181 5 1 1 180
0 182 7 1 2 2172 2181
0 183 5 1 1 182
0 184 7 2 2 181 183
0 185 5 1 1 2195
0 186 7 1 2 2193 185
0 187 5 2 1 186
0 188 7 2 2 169 2197
0 189 5 1 1 2199
0 190 7 1 2 2117 189
0 191 5 2 1 190
0 192 7 1 2 1955 2200
0 193 5 1 1 192
0 194 7 2 2 2201 193
0 195 5 1 1 2203
0 196 7 2 2 2113 2204
0 197 5 2 1 2205
0 198 7 1 2 177 2202
0 199 5 1 1 198
0 200 7 1 2 2183 2192
0 201 5 1 1 200
0 202 7 2 2 199 201
0 203 5 1 1 2209
0 204 7 1 2 2207 203
0 205 5 2 1 204
0 206 7 1 2 2184 2194
0 207 5 1 1 206
0 208 7 1 2 2196 207
0 209 5 1 1 208
0 210 7 3 2 2198 209
0 211 5 1 1 2213
0 212 7 1 2 2208 2214
0 213 5 1 1 212
0 214 7 1 2 2210 213
0 215 5 1 1 214
0 216 7 3 2 2211 215
0 217 5 1 1 2216
0 218 7 2 2 2212 211
0 219 5 1 1 2219
0 220 7 1 2 2114 219
0 221 5 2 1 220
0 222 7 1 2 1952 2220
0 223 5 1 1 222
0 224 7 2 2 2221 223
0 225 5 1 1 2223
0 226 7 2 2 2110 2224
0 227 5 2 1 2225
0 228 7 1 2 195 2222
0 229 5 1 1 228
0 230 7 1 2 2206 2215
0 231 5 1 1 230
0 232 7 2 2 229 231
0 233 5 1 1 2229
0 234 7 1 2 2227 233
0 235 5 2 1 234
0 236 7 2 2 217 2231
0 237 5 1 1 2233
0 238 7 1 2 2111 237
0 239 5 2 1 238
0 240 7 1 2 1949 2234
0 241 5 1 1 240
0 242 7 2 2 2235 241
0 243 5 1 1 2237
0 244 7 2 2 2107 2238
0 245 5 2 1 2239
0 246 7 1 2 225 2236
0 247 5 1 1 246
0 248 7 1 2 2217 2226
0 249 5 1 1 248
0 250 7 2 2 247 249
0 251 5 1 1 2243
0 252 7 1 2 2241 251
0 253 5 2 1 252
0 254 7 1 2 2218 2228
0 255 5 1 1 254
0 256 7 1 2 2230 255
0 257 5 1 1 256
0 258 7 3 2 2232 257
0 259 5 1 1 2247
0 260 7 1 2 2242 2248
0 261 5 1 1 260
0 262 7 1 2 2244 261
0 263 5 1 1 262
0 264 7 3 2 2245 263
0 265 5 1 1 2250
0 266 7 2 2 2246 259
0 267 5 1 1 2253
0 268 7 1 2 2108 267
0 269 5 2 1 268
0 270 7 1 2 1946 2254
0 271 5 1 1 270
0 272 7 2 2 2255 271
0 273 5 1 1 2257
0 274 7 2 2 2104 2258
0 275 5 2 1 2259
0 276 7 1 2 243 2256
0 277 5 1 1 276
0 278 7 1 2 2240 2249
0 279 5 1 1 278
0 280 7 2 2 277 279
0 281 5 1 1 2263
0 282 7 1 2 2261 281
0 283 5 2 1 282
0 284 7 2 2 265 2265
0 285 5 1 1 2267
0 286 7 1 2 2105 285
0 287 5 2 1 286
0 288 7 1 2 1943 2268
0 289 5 1 1 288
0 290 7 2 2 2269 289
0 291 5 1 1 2271
0 292 7 2 2 2101 2272
0 293 5 2 1 2273
0 294 7 1 2 273 2270
0 295 5 1 1 294
0 296 7 1 2 2251 2260
0 297 5 1 1 296
0 298 7 2 2 295 297
0 299 5 1 1 2277
0 300 7 1 2 2275 299
0 301 5 2 1 300
0 302 7 1 2 2252 2262
0 303 5 1 1 302
0 304 7 1 2 2264 303
0 305 5 1 1 304
0 306 7 3 2 2266 305
0 307 5 1 1 2281
0 308 7 1 2 2276 2282
0 309 5 1 1 308
0 310 7 1 2 2278 309
0 311 5 1 1 310
0 312 7 3 2 2279 311
0 313 5 1 1 2284
0 314 7 2 2 2280 307
0 315 5 1 1 2287
0 316 7 1 2 2102 315
0 317 5 2 1 316
0 318 7 1 2 1940 2288
0 319 5 1 1 318
0 320 7 2 2 2289 319
0 321 5 1 1 2291
0 322 7 2 2 2098 2292
0 323 5 2 1 2293
0 324 7 1 2 291 2290
0 325 5 1 1 324
0 326 7 1 2 2274 2283
0 327 5 1 1 326
0 328 7 2 2 325 327
0 329 5 1 1 2297
0 330 7 1 2 2295 329
0 331 5 2 1 330
0 332 7 2 2 313 2299
0 333 5 1 1 2301
0 334 7 1 2 2099 333
0 335 5 2 1 334
0 336 7 1 2 1937 2302
0 337 5 1 1 336
0 338 7 2 2 2303 337
0 339 5 1 1 2305
0 340 7 2 2 2095 2306
0 341 5 2 1 2307
0 342 7 1 2 321 2304
0 343 5 1 1 342
0 344 7 1 2 2285 2294
0 345 5 1 1 344
0 346 7 2 2 343 345
0 347 5 1 1 2311
0 348 7 1 2 2309 347
0 349 5 2 1 348
0 350 7 1 2 2286 2296
0 351 5 1 1 350
0 352 7 1 2 2298 351
0 353 5 1 1 352
0 354 7 3 2 2300 353
0 355 5 1 1 2315
0 356 7 1 2 2310 2316
0 357 5 1 1 356
0 358 7 1 2 2312 357
0 359 5 1 1 358
0 360 7 3 2 2313 359
0 361 5 1 1 2318
0 362 7 2 2 2314 355
0 363 5 1 1 2321
0 364 7 1 2 2096 363
0 365 5 2 1 364
0 366 7 1 2 1934 2322
0 367 5 1 1 366
0 368 7 2 2 2323 367
0 369 5 1 1 2325
0 370 7 2 2 2092 2326
0 371 5 2 1 2327
0 372 7 1 2 339 2324
0 373 5 1 1 372
0 374 7 1 2 2308 2317
0 375 5 1 1 374
0 376 7 2 2 373 375
0 377 5 1 1 2331
0 378 7 1 2 2329 377
0 379 5 2 1 378
0 380 7 2 2 361 2333
0 381 5 1 1 2335
0 382 7 1 2 2093 381
0 383 5 2 1 382
0 384 7 1 2 1931 2336
0 385 5 1 1 384
0 386 7 2 2 2337 385
0 387 5 1 1 2339
0 388 7 2 2 2089 2340
0 389 5 2 1 2341
0 390 7 1 2 369 2338
0 391 5 1 1 390
0 392 7 1 2 2319 2328
0 393 5 1 1 392
0 394 7 2 2 391 393
0 395 5 1 1 2345
0 396 7 1 2 2343 395
0 397 5 2 1 396
0 398 7 1 2 2320 2330
0 399 5 1 1 398
0 400 7 1 2 2332 399
0 401 5 1 1 400
0 402 7 3 2 2334 401
0 403 5 1 1 2349
0 404 7 1 2 2344 2350
0 405 5 1 1 404
0 406 7 1 2 2346 405
0 407 5 1 1 406
0 408 7 3 2 2347 407
0 409 5 1 1 2352
0 410 7 2 2 2348 403
0 411 5 1 1 2355
0 412 7 1 2 2090 411
0 413 5 2 1 412
0 414 7 1 2 1928 2356
0 415 5 1 1 414
0 416 7 2 2 2357 415
0 417 5 1 1 2359
0 418 7 2 2 2086 2360
0 419 5 2 1 2361
0 420 7 1 2 387 2358
0 421 5 1 1 420
0 422 7 1 2 2342 2351
0 423 5 1 1 422
0 424 7 2 2 421 423
0 425 5 1 1 2365
0 426 7 1 2 2363 425
0 427 5 2 1 426
0 428 7 2 2 409 2367
0 429 5 1 1 2369
0 430 7 1 2 2087 429
0 431 5 2 1 430
0 432 7 1 2 1925 2370
0 433 5 1 1 432
0 434 7 2 2 2371 433
0 435 5 1 1 2373
0 436 7 2 2 2082 2374
0 437 5 2 1 2375
0 438 7 1 2 417 2372
0 439 5 1 1 438
0 440 7 1 2 2353 2362
0 441 5 1 1 440
0 442 7 2 2 439 441
0 443 5 1 1 2379
0 444 7 1 2 2377 443
0 445 5 2 1 444
0 446 7 1 2 2354 2364
0 447 5 1 1 446
0 448 7 1 2 2366 447
0 449 5 1 1 448
0 450 7 3 2 2368 449
0 451 5 1 1 2383
0 452 7 1 2 2378 2384
0 453 5 1 1 452
0 454 7 1 2 2380 453
0 455 5 1 1 454
0 456 7 3 2 2381 455
0 457 5 1 1 2386
0 458 7 2 2 2382 451
0 459 5 1 1 2389
0 460 7 1 2 2083 459
0 461 5 2 1 460
0 462 7 1 2 1922 2390
0 463 5 1 1 462
0 464 7 2 2 2391 463
0 465 5 1 1 2393
0 466 7 2 2 2078 2394
0 467 5 2 1 2395
0 468 7 1 2 435 2392
0 469 5 1 1 468
0 470 7 1 2 2376 2385
0 471 5 1 1 470
0 472 7 2 2 469 471
0 473 5 1 1 2399
0 474 7 1 2 2397 473
0 475 5 2 1 474
0 476 7 2 2 457 2401
0 477 5 1 1 2403
0 478 7 1 2 2079 477
0 479 5 2 1 478
0 480 7 1 2 1919 2404
0 481 5 1 1 480
0 482 7 2 2 2405 481
0 483 5 1 1 2407
0 484 7 2 2 2074 2408
0 485 5 2 1 2409
0 486 7 1 2 465 2406
0 487 5 1 1 486
0 488 7 1 2 2387 2396
0 489 5 1 1 488
0 490 7 2 2 487 489
0 491 5 1 1 2413
0 492 7 1 2 2411 491
0 493 5 2 1 492
0 494 7 1 2 2388 2398
0 495 5 1 1 494
0 496 7 1 2 2400 495
0 497 5 1 1 496
0 498 7 3 2 2402 497
0 499 5 1 1 2417
0 500 7 1 2 2412 2418
0 501 5 1 1 500
0 502 7 1 2 2414 501
0 503 5 1 1 502
0 504 7 3 2 2415 503
0 505 5 1 1 2420
0 506 7 2 2 2416 499
0 507 5 1 1 2423
0 508 7 1 2 2075 507
0 509 5 2 1 508
0 510 7 1 2 1916 2424
0 511 5 1 1 510
0 512 7 2 2 2425 511
0 513 5 1 1 2427
0 514 7 2 2 2070 2428
0 515 5 2 1 2429
0 516 7 1 2 483 2426
0 517 5 1 1 516
0 518 7 1 2 2410 2419
0 519 5 1 1 518
0 520 7 2 2 517 519
0 521 5 1 1 2433
0 522 7 1 2 2431 521
0 523 5 2 1 522
0 524 7 2 2 505 2435
0 525 5 1 1 2437
0 526 7 1 2 2071 525
0 527 5 2 1 526
0 528 7 1 2 1913 2438
0 529 5 1 1 528
0 530 7 2 2 2439 529
0 531 5 1 1 2441
0 532 7 2 2 2066 2442
0 533 5 2 1 2443
0 534 7 1 2 513 2440
0 535 5 1 1 534
0 536 7 1 2 2421 2430
0 537 5 1 1 536
0 538 7 2 2 535 537
0 539 5 1 1 2447
0 540 7 1 2 2445 539
0 541 5 2 1 540
0 542 7 1 2 2422 2432
0 543 5 1 1 542
0 544 7 1 2 2434 543
0 545 5 1 1 544
0 546 7 3 2 2436 545
0 547 5 1 1 2451
0 548 7 1 2 2446 2452
0 549 5 1 1 548
0 550 7 1 2 2448 549
0 551 5 1 1 550
0 552 7 3 2 2449 551
0 553 5 1 1 2454
0 554 7 2 2 2450 547
0 555 5 1 1 2457
0 556 7 1 2 2067 555
0 557 5 2 1 556
0 558 7 1 2 1910 2458
0 559 5 1 1 558
0 560 7 2 2 2459 559
0 561 5 1 1 2461
0 562 7 2 2 2062 2462
0 563 5 2 1 2463
0 564 7 1 2 531 2460
0 565 5 1 1 564
0 566 7 1 2 2444 2453
0 567 5 1 1 566
0 568 7 2 2 565 567
0 569 5 1 1 2467
0 570 7 1 2 2465 569
0 571 5 2 1 570
0 572 7 2 2 553 2469
0 573 5 1 1 2471
0 574 7 1 2 2063 573
0 575 5 2 1 574
0 576 7 1 2 1907 2472
0 577 5 1 1 576
0 578 7 2 2 2473 577
0 579 5 1 1 2475
0 580 7 2 2 2058 2476
0 581 5 2 1 2477
0 582 7 1 2 561 2474
0 583 5 1 1 582
0 584 7 1 2 2455 2464
0 585 5 1 1 584
0 586 7 2 2 583 585
0 587 5 1 1 2481
0 588 7 1 2 2479 587
0 589 5 2 1 588
0 590 7 1 2 2456 2466
0 591 5 1 1 590
0 592 7 1 2 2468 591
0 593 5 1 1 592
0 594 7 3 2 2470 593
0 595 5 1 1 2485
0 596 7 1 2 2480 2486
0 597 5 1 1 596
0 598 7 1 2 2482 597
0 599 5 1 1 598
0 600 7 3 2 2483 599
0 601 5 1 1 2488
0 602 7 2 2 2484 595
0 603 5 1 1 2491
0 604 7 1 2 2059 603
0 605 5 2 1 604
0 606 7 1 2 1904 2492
0 607 5 1 1 606
0 608 7 2 2 2493 607
0 609 5 1 1 2495
0 610 7 2 2 2054 2496
0 611 5 2 1 2497
0 612 7 1 2 579 2494
0 613 5 1 1 612
0 614 7 1 2 2478 2487
0 615 5 1 1 614
0 616 7 2 2 613 615
0 617 5 1 1 2501
0 618 7 1 2 2499 617
0 619 5 2 1 618
0 620 7 2 2 601 2503
0 621 5 1 1 2505
0 622 7 1 2 2055 621
0 623 5 2 1 622
0 624 7 1 2 1901 2506
0 625 5 1 1 624
0 626 7 2 2 2507 625
0 627 5 1 1 2509
0 628 7 2 2 2050 2510
0 629 5 2 1 2511
0 630 7 1 2 609 2508
0 631 5 1 1 630
0 632 7 1 2 2489 2498
0 633 5 1 1 632
0 634 7 2 2 631 633
0 635 5 1 1 2515
0 636 7 1 2 2513 635
0 637 5 2 1 636
0 638 7 1 2 2490 2500
0 639 5 1 1 638
0 640 7 1 2 2502 639
0 641 5 1 1 640
0 642 7 3 2 2504 641
0 643 5 1 1 2519
0 644 7 1 2 2514 2520
0 645 5 1 1 644
0 646 7 1 2 2516 645
0 647 5 1 1 646
0 648 7 3 2 2517 647
0 649 5 1 1 2522
0 650 7 2 2 2518 643
0 651 5 1 1 2525
0 652 7 1 2 2051 651
0 653 5 2 1 652
0 654 7 1 2 1898 2526
0 655 5 1 1 654
0 656 7 2 2 2527 655
0 657 5 1 1 2529
0 658 7 2 2 2046 2530
0 659 5 2 1 2531
0 660 7 1 2 627 2528
0 661 5 1 1 660
0 662 7 1 2 2512 2521
0 663 5 1 1 662
0 664 7 2 2 661 663
0 665 5 1 1 2535
0 666 7 1 2 2533 665
0 667 5 2 1 666
0 668 7 2 2 649 2537
0 669 5 1 1 2539
0 670 7 1 2 2047 669
0 671 5 2 1 670
0 672 7 1 2 1895 2540
0 673 5 1 1 672
0 674 7 2 2 2541 673
0 675 5 1 1 2543
0 676 7 2 2 2042 2544
0 677 5 2 1 2545
0 678 7 1 2 657 2542
0 679 5 1 1 678
0 680 7 1 2 2523 2532
0 681 5 1 1 680
0 682 7 2 2 679 681
0 683 5 1 1 2549
0 684 7 1 2 2547 683
0 685 5 2 1 684
0 686 7 1 2 2524 2534
0 687 5 1 1 686
0 688 7 1 2 2536 687
0 689 5 1 1 688
0 690 7 3 2 2538 689
0 691 5 1 1 2553
0 692 7 1 2 2548 2554
0 693 5 1 1 692
0 694 7 1 2 2550 693
0 695 5 1 1 694
0 696 7 3 2 2551 695
0 697 5 1 1 2556
0 698 7 2 2 2552 691
0 699 5 1 1 2559
0 700 7 1 2 2043 699
0 701 5 2 1 700
0 702 7 1 2 1892 2560
0 703 5 1 1 702
0 704 7 2 2 2561 703
0 705 5 1 1 2563
0 706 7 2 2 2038 2564
0 707 5 2 1 2565
0 708 7 1 2 675 2562
0 709 5 1 1 708
0 710 7 1 2 2546 2555
0 711 5 1 1 710
0 712 7 2 2 709 711
0 713 5 1 1 2569
0 714 7 1 2 2567 713
0 715 5 2 1 714
0 716 7 2 2 697 2571
0 717 5 1 1 2573
0 718 7 1 2 2039 717
0 719 5 2 1 718
0 720 7 1 2 1889 2574
0 721 5 1 1 720
0 722 7 2 2 2575 721
0 723 5 1 1 2577
0 724 7 2 2 2034 2578
0 725 5 2 1 2579
0 726 7 1 2 705 2576
0 727 5 1 1 726
0 728 7 1 2 2557 2566
0 729 5 1 1 728
0 730 7 2 2 727 729
0 731 5 1 1 2583
0 732 7 1 2 2581 731
0 733 5 2 1 732
0 734 7 1 2 2558 2568
0 735 5 1 1 734
0 736 7 1 2 2570 735
0 737 5 1 1 736
0 738 7 3 2 2572 737
0 739 5 1 1 2587
0 740 7 1 2 2582 2588
0 741 5 1 1 740
0 742 7 1 2 2584 741
0 743 5 1 1 742
0 744 7 3 2 2585 743
0 745 5 1 1 2590
0 746 7 2 2 2586 739
0 747 5 1 1 2593
0 748 7 1 2 2035 747
0 749 5 2 1 748
0 750 7 1 2 1886 2594
0 751 5 1 1 750
0 752 7 2 2 2595 751
0 753 5 1 1 2597
0 754 7 2 2 2031 2598
0 755 5 2 1 2599
0 756 7 1 2 723 2596
0 757 5 1 1 756
0 758 7 1 2 2580 2589
0 759 5 1 1 758
0 760 7 2 2 757 759
0 761 5 1 1 2603
0 762 7 1 2 2601 761
0 763 5 2 1 762
0 764 7 2 2 745 2605
0 765 5 1 1 2607
0 766 7 1 2 2032 765
0 767 5 2 1 766
0 768 7 1 2 1883 2608
0 769 5 1 1 768
0 770 7 2 2 2609 769
0 771 5 1 1 2611
0 772 7 2 2 2028 2612
0 773 5 2 1 2613
0 774 7 1 2 753 2610
0 775 5 1 1 774
0 776 7 1 2 2591 2600
0 777 5 1 1 776
0 778 7 2 2 775 777
0 779 5 1 1 2617
0 780 7 1 2 2615 779
0 781 5 2 1 780
0 782 7 1 2 2592 2602
0 783 5 1 1 782
0 784 7 1 2 2604 783
0 785 5 1 1 784
0 786 7 3 2 2606 785
0 787 5 1 1 2621
0 788 7 1 2 2616 2622
0 789 5 1 1 788
0 790 7 1 2 2618 789
0 791 5 1 1 790
0 792 7 3 2 2619 791
0 793 5 1 1 2624
0 794 7 2 2 2620 787
0 795 5 1 1 2627
0 796 7 1 2 2029 795
0 797 5 2 1 796
0 798 7 1 2 1880 2628
0 799 5 1 1 798
0 800 7 2 2 2629 799
0 801 5 1 1 2631
0 802 7 2 2 2025 2632
0 803 5 2 1 2633
0 804 7 1 2 771 2630
0 805 5 1 1 804
0 806 7 1 2 2614 2623
0 807 5 1 1 806
0 808 7 2 2 805 807
0 809 5 1 1 2637
0 810 7 1 2 2635 809
0 811 5 2 1 810
0 812 7 2 2 793 2639
0 813 5 1 1 2641
0 814 7 1 2 2026 813
0 815 5 2 1 814
0 816 7 1 2 1877 2642
0 817 5 1 1 816
0 818 7 2 2 2643 817
0 819 5 1 1 2645
0 820 7 2 2 2022 2646
0 821 5 2 1 2647
0 822 7 1 2 801 2644
0 823 5 1 1 822
0 824 7 1 2 2625 2634
0 825 5 1 1 824
0 826 7 2 2 823 825
0 827 5 1 1 2651
0 828 7 1 2 2649 827
0 829 5 2 1 828
0 830 7 1 2 2626 2636
0 831 5 1 1 830
0 832 7 1 2 2638 831
0 833 5 1 1 832
0 834 7 3 2 2640 833
0 835 5 1 1 2655
0 836 7 1 2 2650 2656
0 837 5 1 1 836
0 838 7 1 2 2652 837
0 839 5 1 1 838
0 840 7 3 2 2653 839
0 841 5 1 1 2658
0 842 7 2 2 2654 835
0 843 5 1 1 2661
0 844 7 1 2 2023 843
0 845 5 2 1 844
0 846 7 1 2 1874 2662
0 847 5 1 1 846
0 848 7 2 2 2663 847
0 849 5 1 1 2665
0 850 7 2 2 2019 2666
0 851 5 2 1 2667
0 852 7 1 2 819 2664
0 853 5 1 1 852
0 854 7 1 2 2648 2657
0 855 5 1 1 854
0 856 7 2 2 853 855
0 857 5 1 1 2671
0 858 7 1 2 2669 857
0 859 5 2 1 858
0 860 7 2 2 841 2673
0 861 5 1 1 2675
0 862 7 1 2 2020 861
0 863 5 2 1 862
0 864 7 1 2 1871 2676
0 865 5 1 1 864
0 866 7 2 2 2677 865
0 867 5 1 1 2679
0 868 7 2 2 2016 2680
0 869 5 2 1 2681
0 870 7 1 2 849 2678
0 871 5 1 1 870
0 872 7 1 2 2659 2668
0 873 5 1 1 872
0 874 7 2 2 871 873
0 875 5 1 1 2685
0 876 7 1 2 2683 875
0 877 5 2 1 876
0 878 7 1 2 2660 2670
0 879 5 1 1 878
0 880 7 1 2 2672 879
0 881 5 1 1 880
0 882 7 3 2 2674 881
0 883 5 1 1 2689
0 884 7 1 2 2684 2690
0 885 5 1 1 884
0 886 7 1 2 2686 885
0 887 5 1 1 886
0 888 7 3 2 2687 887
0 889 5 1 1 2692
0 890 7 2 2 2688 883
0 891 5 1 1 2695
0 892 7 1 2 2017 891
0 893 5 2 1 892
0 894 7 1 2 1868 2696
0 895 5 1 1 894
0 896 7 2 2 2697 895
0 897 5 1 1 2699
0 898 7 2 2 2013 2700
0 899 5 2 1 2701
0 900 7 1 2 867 2698
0 901 5 1 1 900
0 902 7 1 2 2682 2691
0 903 5 1 1 902
0 904 7 2 2 901 903
0 905 5 1 1 2705
0 906 7 1 2 2703 905
0 907 5 2 1 906
0 908 7 2 2 889 2707
0 909 5 1 1 2709
0 910 7 1 2 2014 909
0 911 5 2 1 910
0 912 7 1 2 1865 2710
0 913 5 1 1 912
0 914 7 2 2 2711 913
0 915 5 1 1 2713
0 916 7 2 2 2010 2714
0 917 5 2 1 2715
0 918 7 1 2 897 2712
0 919 5 1 1 918
0 920 7 1 2 2693 2702
0 921 5 1 1 920
0 922 7 2 2 919 921
0 923 5 1 1 2719
0 924 7 1 2 2717 923
0 925 5 2 1 924
0 926 7 1 2 2694 2704
0 927 5 1 1 926
0 928 7 1 2 2706 927
0 929 5 1 1 928
0 930 7 3 2 2708 929
0 931 5 1 1 2723
0 932 7 1 2 2718 2724
0 933 5 1 1 932
0 934 7 1 2 2720 933
0 935 5 1 1 934
0 936 7 3 2 2721 935
0 937 5 1 1 2726
0 938 7 2 2 2722 931
0 939 5 1 1 2729
0 940 7 1 2 2011 939
0 941 5 2 1 940
0 942 7 1 2 1862 2730
0 943 5 1 1 942
0 944 7 2 2 2731 943
0 945 5 1 1 2733
0 946 7 2 2 2007 2734
0 947 5 2 1 2735
0 948 7 1 2 915 2732
0 949 5 1 1 948
0 950 7 1 2 2716 2725
0 951 5 1 1 950
0 952 7 2 2 949 951
0 953 5 1 1 2739
0 954 7 1 2 2737 953
0 955 5 2 1 954
0 956 7 2 2 937 2741
0 957 5 1 1 2743
0 958 7 1 2 2008 957
0 959 5 2 1 958
0 960 7 1 2 1859 2744
0 961 5 1 1 960
0 962 7 2 2 2745 961
0 963 5 1 1 2747
0 964 7 2 2 2004 2748
0 965 5 2 1 2749
0 966 7 1 2 945 2746
0 967 5 1 1 966
0 968 7 1 2 2727 2736
0 969 5 1 1 968
0 970 7 2 2 967 969
0 971 5 1 1 2753
0 972 7 1 2 2751 971
0 973 5 2 1 972
0 974 7 1 2 2728 2738
0 975 5 1 1 974
0 976 7 1 2 2740 975
0 977 5 1 1 976
0 978 7 3 2 2742 977
0 979 5 1 1 2757
0 980 7 1 2 2752 2758
0 981 5 1 1 980
0 982 7 1 2 2754 981
0 983 5 1 1 982
0 984 7 3 2 2755 983
0 985 5 1 1 2760
0 986 7 2 2 2756 979
0 987 5 1 1 2763
0 988 7 1 2 2005 987
0 989 5 2 1 988
0 990 7 1 2 1856 2764
0 991 5 1 1 990
0 992 7 2 2 2765 991
0 993 5 1 1 2767
0 994 7 2 2 2001 2768
0 995 5 2 1 2769
0 996 7 1 2 963 2766
0 997 5 1 1 996
0 998 7 1 2 2750 2759
0 999 5 1 1 998
0 1000 7 2 2 997 999
0 1001 5 1 1 2773
0 1002 7 1 2 2771 1001
0 1003 5 2 1 1002
0 1004 7 2 2 985 2775
0 1005 5 1 1 2777
0 1006 7 1 2 2002 1005
0 1007 5 2 1 1006
0 1008 7 1 2 1853 2778
0 1009 5 1 1 1008
0 1010 7 2 2 2779 1009
0 1011 5 1 1 2781
0 1012 7 2 2 1998 2782
0 1013 5 2 1 2783
0 1014 7 1 2 993 2780
0 1015 5 1 1 1014
0 1016 7 1 2 2761 2770
0 1017 5 1 1 1016
0 1018 7 2 2 1015 1017
0 1019 5 1 1 2787
0 1020 7 1 2 2785 1019
0 1021 5 2 1 1020
0 1022 7 1 2 2762 2772
0 1023 5 1 1 1022
0 1024 7 1 2 2774 1023
0 1025 5 1 1 1024
0 1026 7 3 2 2776 1025
0 1027 5 1 1 2791
0 1028 7 1 2 2786 2792
0 1029 5 1 1 1028
0 1030 7 1 2 2788 1029
0 1031 5 1 1 1030
0 1032 7 3 2 2789 1031
0 1033 5 1 1 2794
0 1034 7 2 2 2790 1027
0 1035 5 1 1 2797
0 1036 7 1 2 1999 1035
0 1037 5 2 1 1036
0 1038 7 1 2 1850 2798
0 1039 5 1 1 1038
0 1040 7 2 2 2799 1039
0 1041 5 1 1 2801
0 1042 7 2 2 1995 2802
0 1043 5 2 1 2803
0 1044 7 1 2 1011 2800
0 1045 5 1 1 1044
0 1046 7 1 2 2784 2793
0 1047 5 1 1 1046
0 1048 7 2 2 1045 1047
0 1049 5 1 1 2807
0 1050 7 1 2 2805 1049
0 1051 5 2 1 1050
0 1052 7 2 2 1033 2809
0 1053 5 1 1 2811
0 1054 7 1 2 1996 1053
0 1055 5 2 1 1054
0 1056 7 1 2 1847 2812
0 1057 5 1 1 1056
0 1058 7 2 2 2813 1057
0 1059 5 1 1 2815
0 1060 7 2 2 1992 2816
0 1061 5 2 1 2817
0 1062 7 1 2 1041 2814
0 1063 5 1 1 1062
0 1064 7 1 2 2795 2804
0 1065 5 1 1 1064
0 1066 7 2 2 1063 1065
0 1067 5 1 1 2821
0 1068 7 1 2 2819 1067
0 1069 5 2 1 1068
0 1070 7 1 2 2796 2806
0 1071 5 1 1 1070
0 1072 7 1 2 2808 1071
0 1073 5 1 1 1072
0 1074 7 3 2 2810 1073
0 1075 5 1 1 2825
0 1076 7 1 2 2820 2826
0 1077 5 1 1 1076
0 1078 7 1 2 2822 1077
0 1079 5 1 1 1078
0 1080 7 3 2 2823 1079
0 1081 5 1 1 2828
0 1082 7 2 2 2824 1075
0 1083 5 1 1 2831
0 1084 7 1 2 1993 1083
0 1085 5 2 1 1084
0 1086 7 1 2 1844 2832
0 1087 5 1 1 1086
0 1088 7 2 2 2833 1087
0 1089 5 1 1 2835
0 1090 7 2 2 1989 2836
0 1091 5 2 1 2837
0 1092 7 1 2 1059 2834
0 1093 5 1 1 1092
0 1094 7 1 2 2818 2827
0 1095 5 1 1 1094
0 1096 7 2 2 1093 1095
0 1097 5 1 1 2841
0 1098 7 1 2 2839 1097
0 1099 5 2 1 1098
0 1100 7 2 2 1081 2843
0 1101 5 1 1 2845
0 1102 7 1 2 1990 1101
0 1103 5 2 1 1102
0 1104 7 1 2 1841 2846
0 1105 5 1 1 1104
0 1106 7 2 2 2847 1105
0 1107 5 1 1 2849
0 1108 7 2 2 1986 2850
0 1109 5 2 1 2851
0 1110 7 1 2 1089 2848
0 1111 5 1 1 1110
0 1112 7 1 2 2829 2838
0 1113 5 1 1 1112
0 1114 7 2 2 1111 1113
0 1115 5 1 1 2855
0 1116 7 1 2 2853 1115
0 1117 5 2 1 1116
0 1118 7 1 2 2830 2840
0 1119 5 1 1 1118
0 1120 7 1 2 2842 1119
0 1121 5 1 1 1120
0 1122 7 3 2 2844 1121
0 1123 5 1 1 2859
0 1124 7 1 2 2854 2860
0 1125 5 1 1 1124
0 1126 7 1 2 2856 1125
0 1127 5 1 1 1126
0 1128 7 3 2 2857 1127
0 1129 5 1 1 2862
0 1130 7 2 2 2858 1123
0 1131 5 1 1 2865
0 1132 7 1 2 1987 1131
0 1133 5 2 1 1132
0 1134 7 1 2 1838 2866
0 1135 5 1 1 1134
0 1136 7 2 2 2867 1135
0 1137 5 1 1 2869
0 1138 7 2 2 1983 2870
0 1139 5 2 1 2871
0 1140 7 1 2 1107 2868
0 1141 5 1 1 1140
0 1142 7 1 2 2852 2861
0 1143 5 1 1 1142
0 1144 7 2 2 1141 1143
0 1145 5 1 1 2875
0 1146 7 1 2 2873 1145
0 1147 5 2 1 1146
0 1148 7 2 2 1129 2877
0 1149 5 1 1 2879
0 1150 7 1 2 1984 1149
0 1151 5 2 1 1150
0 1152 7 1 2 1835 2880
0 1153 5 1 1 1152
0 1154 7 2 2 2881 1153
0 1155 5 1 1 2883
0 1156 7 2 2 1980 2884
0 1157 5 1 1 2885
0 1158 7 1 2 1137 2882
0 1159 5 1 1 1158
0 1160 7 1 2 2863 2872
0 1161 5 1 1 1160
0 1162 7 2 2 1159 1161
0 1163 5 1 1 2887
0 1164 7 1 2 1157 1163
0 1165 5 2 1 1164
0 1166 7 1 2 2864 2874
0 1167 5 1 1 1166
0 1168 7 1 2 2876 1167
0 1169 5 1 1 1168
0 1170 7 2 2 2878 1169
0 1171 5 2 1 2891
0 1172 7 1 2 2889 2893
0 1173 5 1 1 1172
0 1174 7 1 2 1981 1173
0 1175 5 2 1 1174
0 1176 7 2 2 2888 2894
0 1177 5 1 1 2897
0 1178 7 1 2 1832 2898
0 1179 5 1 1 1178
0 1180 7 2 2 2895 1179
0 1181 5 1 1 2899
0 1182 7 1 2 1155 2896
0 1183 5 2 1 1182
0 1184 7 1 2 2886 2892
0 1185 5 1 1 1184
0 1186 7 1 2 2901 1185
0 1187 7 1 2 1181 1186
0 1188 5 1 1 1187
0 1189 7 1 2 2890 1177
0 1190 5 1 1 1189
0 1191 7 1 2 2902 1190
0 1192 5 1 1 1191
0 1193 7 1 2 1829 1192
0 1194 5 1 1 1193
0 1195 7 1 2 1978 2900
0 1196 5 1 1 1195
0 1197 7 1 2 1194 1196
0 1198 7 2 2 1188 1197
0 1199 5 1 1 2903
0 1200 7 1 2 1985 2033
0 1201 5 2 1 1200
0 1202 7 1 2 1836 1884
0 1203 5 2 1 1202
0 1204 7 1 2 1982 2030
0 1205 5 2 1 1204
0 1206 7 1 2 1833 1881
0 1207 5 2 1 1206
0 1208 7 2 2 1830 1878
0 1209 5 3 1 2913
0 1210 7 1 2 2911 2915
0 1211 5 1 1 1210
0 1212 7 2 2 2909 1211
0 1213 5 2 1 2918
0 1214 7 1 2 2907 2920
0 1215 5 1 1 1214
0 1216 7 2 2 2905 1215
0 1217 5 1 1 2922
0 1218 7 1 2 1988 1217
0 1219 5 2 1 1218
0 1220 7 1 2 1839 2923
0 1221 5 2 1 1220
0 1222 7 1 2 2036 2926
0 1223 5 1 1 1222
0 1224 7 2 2 2924 1223
0 1225 5 1 1 2928
0 1226 7 1 2 1991 1225
0 1227 5 2 1 1226
0 1228 7 1 2 1842 2929
0 1229 5 2 1 1228
0 1230 7 1 2 2040 2932
0 1231 5 1 1 1230
0 1232 7 2 2 2930 1231
0 1233 5 1 1 2934
0 1234 7 1 2 1994 1233
0 1235 5 2 1 1234
0 1236 7 1 2 1845 2935
0 1237 5 2 1 1236
0 1238 7 1 2 2044 2938
0 1239 5 1 1 1238
0 1240 7 2 2 2936 1239
0 1241 5 1 1 2940
0 1242 7 1 2 1997 1241
0 1243 5 2 1 1242
0 1244 7 1 2 1848 2941
0 1245 5 2 1 1244
0 1246 7 1 2 2048 2944
0 1247 5 1 1 1246
0 1248 7 2 2 2942 1247
0 1249 5 1 1 2946
0 1250 7 1 2 2000 1249
0 1251 5 2 1 1250
0 1252 7 1 2 1851 2947
0 1253 5 2 1 1252
0 1254 7 1 2 2052 2950
0 1255 5 1 1 1254
0 1256 7 2 2 2948 1255
0 1257 5 1 1 2952
0 1258 7 1 2 2003 1257
0 1259 5 2 1 1258
0 1260 7 1 2 1854 2953
0 1261 5 2 1 1260
0 1262 7 1 2 2056 2956
0 1263 5 1 1 1262
0 1264 7 2 2 2954 1263
0 1265 5 1 1 2958
0 1266 7 1 2 2006 1265
0 1267 5 2 1 1266
0 1268 7 1 2 1857 2959
0 1269 5 2 1 1268
0 1270 7 1 2 2060 2962
0 1271 5 1 1 1270
0 1272 7 2 2 2960 1271
0 1273 5 1 1 2964
0 1274 7 1 2 2009 1273
0 1275 5 2 1 1274
0 1276 7 1 2 1860 2965
0 1277 5 2 1 1276
0 1278 7 1 2 2064 2968
0 1279 5 1 1 1278
0 1280 7 2 2 2966 1279
0 1281 5 1 1 2970
0 1282 7 1 2 2012 1281
0 1283 5 2 1 1282
0 1284 7 1 2 1863 2971
0 1285 5 2 1 1284
0 1286 7 1 2 2068 2974
0 1287 5 1 1 1286
0 1288 7 2 2 2972 1287
0 1289 5 1 1 2976
0 1290 7 1 2 2015 1289
0 1291 5 2 1 1290
0 1292 7 1 2 1866 2977
0 1293 5 2 1 1292
0 1294 7 1 2 2072 2980
0 1295 5 1 1 1294
0 1296 7 2 2 2978 1295
0 1297 5 1 1 2982
0 1298 7 1 2 2018 1297
0 1299 5 2 1 1298
0 1300 7 1 2 1869 2983
0 1301 5 2 1 1300
0 1302 7 1 2 2076 2986
0 1303 5 1 1 1302
0 1304 7 2 2 2984 1303
0 1305 5 1 1 2988
0 1306 7 1 2 2021 1305
0 1307 5 2 1 1306
0 1308 7 1 2 1872 2989
0 1309 5 2 1 1308
0 1310 7 1 2 2080 2992
0 1311 5 1 1 1310
0 1312 7 2 2 2990 1311
0 1313 5 1 1 2994
0 1314 7 1 2 2024 1313
0 1315 5 2 1 1314
0 1316 7 1 2 1875 2995
0 1317 5 2 1 1316
0 1318 7 2 2 2996 2998
0 1319 5 1 1 3000
0 1320 7 1 2 1923 3001
0 1321 5 1 1 1320
0 1322 7 1 2 2084 1319
0 1323 5 1 1 1322
0 1324 7 2 2 1321 1323
0 1325 5 1 1 3002
0 1326 7 1 2 1973 1325
0 1327 5 3 1 1326
0 1328 7 1 2 2085 2999
0 1329 5 1 1 1328
0 1330 7 2 2 2997 1329
0 1331 5 1 1 3007
0 1332 7 1 2 2135 3008
0 1333 5 3 1 1332
0 1334 7 1 2 2133 3003
0 1335 5 4 1 1334
0 1336 7 2 2 2991 2993
0 1337 5 1 1 3016
0 1338 7 1 2 1920 3017
0 1339 5 1 1 1338
0 1340 7 1 2 2081 1337
0 1341 5 1 1 1340
0 1342 7 2 2 1339 1341
0 1343 5 1 1 3018
0 1344 7 1 2 1969 1343
0 1345 5 3 1 1344
0 1346 7 1 2 2131 3019
0 1347 5 4 1 1346
0 1348 7 2 2 2985 2987
0 1349 5 1 1 3027
0 1350 7 1 2 1917 3028
0 1351 5 1 1 1350
0 1352 7 1 2 2077 1349
0 1353 5 1 1 1352
0 1354 7 2 2 1351 1353
0 1355 5 1 1 3029
0 1356 7 1 2 1966 1355
0 1357 5 3 1 1356
0 1358 7 1 2 2128 3030
0 1359 5 5 1 1358
0 1360 7 2 2 2979 2981
0 1361 5 1 1 3039
0 1362 7 1 2 1914 3040
0 1363 5 1 1 1362
0 1364 7 1 2 2073 1361
0 1365 5 1 1 1364
0 1366 7 2 2 1363 1365
0 1367 5 1 1 3041
0 1368 7 1 2 1962 1367
0 1369 5 3 1 1368
0 1370 7 1 2 2124 3042
0 1371 5 5 1 1370
0 1372 7 2 2 2973 2975
0 1373 5 1 1 3051
0 1374 7 1 2 1911 3052
0 1375 5 1 1 1374
0 1376 7 1 2 2069 1373
0 1377 5 1 1 1376
0 1378 7 2 2 1375 1377
0 1379 5 1 1 3053
0 1380 7 1 2 1959 1379
0 1381 5 4 1 1380
0 1382 7 2 2 2961 2963
0 1383 5 1 1 3059
0 1384 7 1 2 1905 3060
0 1385 5 1 1 1384
0 1386 7 1 2 2061 1383
0 1387 5 1 1 1386
0 1388 7 2 2 1385 1387
0 1389 5 1 1 3061
0 1390 7 1 2 1953 1389
0 1391 5 3 1 1390
0 1392 7 1 2 2115 3062
0 1393 5 4 1 1392
0 1394 7 2 2 2955 2957
0 1395 5 1 1 3070
0 1396 7 1 2 1902 3071
0 1397 5 1 1 1396
0 1398 7 1 2 2057 1395
0 1399 5 1 1 1398
0 1400 7 2 2 1397 1399
0 1401 5 1 1 3072
0 1402 7 1 2 2112 3073
0 1403 5 4 1 1402
0 1404 7 1 2 1950 1401
0 1405 5 3 1 1404
0 1406 7 2 2 2949 2951
0 1407 5 1 1 3081
0 1408 7 1 2 1899 3082
0 1409 5 1 1 1408
0 1410 7 1 2 2053 1407
0 1411 5 1 1 1410
0 1412 7 2 2 1409 1411
0 1413 5 1 1 3083
0 1414 7 1 2 2109 3084
0 1415 5 4 1 1414
0 1416 7 1 2 1947 1413
0 1417 5 3 1 1416
0 1418 7 2 2 2943 2945
0 1419 5 1 1 3092
0 1420 7 1 2 1896 3093
0 1421 5 1 1 1420
0 1422 7 1 2 2049 1419
0 1423 5 1 1 1422
0 1424 7 2 2 1421 1423
0 1425 5 1 1 3094
0 1426 7 1 2 2106 3095
0 1427 5 4 1 1426
0 1428 7 1 2 1944 1425
0 1429 5 4 1 1428
0 1430 7 2 2 2937 2939
0 1431 5 1 1 3104
0 1432 7 1 2 1893 3105
0 1433 5 1 1 1432
0 1434 7 1 2 2045 1431
0 1435 5 1 1 1434
0 1436 7 2 2 1433 1435
0 1437 5 1 1 3106
0 1438 7 1 2 2103 3107
0 1439 5 5 1 1438
0 1440 7 1 2 1941 1437
0 1441 5 4 1 1440
0 1442 7 2 2 2931 2933
0 1443 5 1 1 3117
0 1444 7 1 2 1890 3118
0 1445 5 1 1 1444
0 1446 7 1 2 2041 1443
0 1447 5 1 1 1446
0 1448 7 2 2 1445 1447
0 1449 5 1 1 3119
0 1450 7 1 2 2100 3120
0 1451 5 4 1 1450
0 1452 7 1 2 1938 1449
0 1453 5 3 1 1452
0 1454 7 2 2 2925 2927
0 1455 5 1 1 3128
0 1456 7 1 2 1887 3129
0 1457 5 1 1 1456
0 1458 7 1 2 2037 1455
0 1459 5 1 1 1458
0 1460 7 2 2 1457 1459
0 1461 5 1 1 3130
0 1462 7 1 2 2097 3131
0 1463 5 4 1 1462
0 1464 7 1 2 1935 1461
0 1465 5 3 1 1464
0 1466 7 2 2 2906 2908
0 1467 5 1 1 3139
0 1468 7 1 2 2919 1467
0 1469 5 1 1 1468
0 1470 7 1 2 2921 3140
0 1471 5 1 1 1470
0 1472 7 2 2 1469 1471
0 1473 5 1 1 3141
0 1474 7 1 2 1932 3142
0 1475 5 2 1 1474
0 1476 7 2 2 2910 2912
0 1477 5 1 1 3145
0 1478 7 1 2 2914 1477
0 1479 5 1 1 1478
0 1480 7 1 2 2916 3146
0 1481 5 1 1 1480
0 1482 7 2 2 1479 1481
0 1483 5 1 1 3147
0 1484 7 1 2 1929 3148
0 1485 5 1 1 1484
0 1486 7 2 2 3143 1485
0 1487 5 1 1 3149
0 1488 7 1 2 1979 2027
0 1489 5 1 1 1488
0 1490 7 2 2 2917 1489
0 1491 5 1 1 3151
0 1492 7 1 2 1926 1491
0 1493 5 1 1 1492
0 1494 7 2 2 3150 1493
0 1495 5 1 1 3153
0 1496 7 2 2 2091 1483
0 1497 5 1 1 3155
0 1498 7 1 2 3144 3156
0 1499 5 1 1 1498
0 1500 7 1 2 2094 1473
0 1501 5 3 1 1500
0 1502 7 1 2 1499 3157
0 1503 7 2 2 1495 1502
0 1504 5 2 1 3160
0 1505 7 1 2 3136 3162
0 1506 5 1 1 1505
0 1507 7 2 2 3132 1506
0 1508 5 2 1 3164
0 1509 7 1 2 3125 3166
0 1510 5 1 1 1509
0 1511 7 2 2 3121 1510
0 1512 5 1 1 3168
0 1513 7 1 2 3113 1512
0 1514 5 2 1 1513
0 1515 7 1 2 3108 3170
0 1516 5 1 1 1515
0 1517 7 1 2 3100 1516
0 1518 5 1 1 1517
0 1519 7 1 2 3096 1518
0 1520 5 2 1 1519
0 1521 7 1 2 3089 3172
0 1522 5 1 1 1521
0 1523 7 2 2 3085 1522
0 1524 5 2 1 3174
0 1525 7 1 2 3078 3176
0 1526 5 1 1 1525
0 1527 7 3 2 3074 1526
0 1528 5 1 1 3178
0 1529 7 1 2 3066 3179
0 1530 5 1 1 1529
0 1531 7 3 2 3063 1530
0 1532 5 1 1 3181
0 1533 7 2 2 2967 2969
0 1534 5 1 1 3184
0 1535 7 1 2 1908 3185
0 1536 5 1 1 1535
0 1537 7 1 2 2065 1534
0 1538 5 1 1 1537
0 1539 7 2 2 1536 1538
0 1540 5 1 1 3186
0 1541 7 3 2 1956 1540
0 1542 5 2 1 3188
0 1543 7 1 2 3182 3191
0 1544 5 1 1 1543
0 1545 7 3 2 2118 3187
0 1546 5 2 1 3193
0 1547 7 1 2 2121 3054
0 1548 5 4 1 1547
0 1549 7 2 2 3196 3198
0 1550 7 1 2 1544 3202
0 1551 5 1 1 1550
0 1552 7 1 2 3055 1551
0 1553 5 2 1 1552
0 1554 7 1 2 3046 3204
0 1555 5 1 1 1554
0 1556 7 2 2 3043 1555
0 1557 5 2 1 3206
0 1558 7 1 2 3034 3208
0 1559 5 1 1 1558
0 1560 7 2 2 3031 1559
0 1561 5 2 1 3210
0 1562 7 1 2 3023 3212
0 1563 5 1 1 1562
0 1564 7 3 2 3020 1563
0 1565 5 1 1 3214
0 1566 7 1 2 3012 1565
0 1567 5 1 1 1566
0 1568 7 1 2 3009 1567
0 1569 5 1 1 1568
0 1570 7 1 2 3004 1569
0 1571 5 1 1 1570
0 1572 7 2 2 1977 1331
0 1573 5 1 1 3217
0 1574 7 2 2 3010 3013
0 1575 7 1 2 3005 3215
0 1576 5 1 1 1575
0 1577 7 1 2 3219 1576
0 1578 5 1 1 1577
0 1579 7 3 2 1573 1578
0 1580 5 1 1 3221
0 1581 7 2 2 3014 3006
0 1582 5 2 1 3224
0 1583 7 1 2 3216 3226
0 1584 5 1 1 1583
0 1585 7 3 2 3021 3024
0 1586 5 2 1 3228
0 1587 7 1 2 3211 3231
0 1588 5 1 1 1587
0 1589 7 1 2 3213 3229
0 1590 5 1 1 1589
0 1591 7 2 2 3032 3035
0 1592 5 2 1 3233
0 1593 7 1 2 3207 3235
0 1594 5 1 1 1593
0 1595 7 1 2 3209 3234
0 1596 5 1 1 1595
0 1597 7 2 2 3044 3047
0 1598 5 2 1 3237
0 1599 7 1 2 3056 3239
0 1600 5 1 1 1599
0 1601 7 1 2 3205 3238
0 1602 5 1 1 1601
0 1603 7 1 2 3057 3199
0 1604 5 2 1 1603
0 1605 7 1 2 1532 3189
0 1606 5 1 1 1605
0 1607 7 1 2 3241 1606
0 1608 5 1 1 1607
0 1609 7 1 2 3194 3183
0 1610 5 1 1 1609
0 1611 7 3 2 3064 3067
0 1612 5 2 1 3243
0 1613 7 1 2 1528 3244
0 1614 5 1 1 1613
0 1615 7 1 2 3180 3246
0 1616 5 1 1 1615
0 1617 7 3 2 3075 3079
0 1618 5 2 1 3248
0 1619 7 1 2 3175 3251
0 1620 5 1 1 1619
0 1621 7 1 2 3177 3249
0 1622 5 1 1 1621
0 1623 7 3 2 3086 3090
0 1624 5 2 1 3253
0 1625 7 1 2 3173 3254
0 1626 5 1 1 1625
0 1627 7 1 2 3097 3256
0 1628 5 1 1 1627
0 1629 7 2 2 3098 3101
0 1630 7 1 2 3171 3258
0 1631 5 1 1 1630
0 1632 7 1 2 3109 1631
0 1633 5 1 1 1632
0 1634 7 1 2 3110 3114
0 1635 5 2 1 1634
0 1636 7 1 2 3169 3260
0 1637 5 1 1 1636
0 1638 7 3 2 3122 3126
0 1639 5 2 1 3262
0 1640 7 1 2 3165 3263
0 1641 5 1 1 1640
0 1642 7 3 2 3133 3137
0 1643 5 2 1 3267
0 1644 7 1 2 3163 3268
0 1645 5 1 1 1644
0 1646 7 1 2 2088 3152
0 1647 5 1 1 1646
0 1648 7 1 2 1497 1647
0 1649 7 3 2 3158 1648
0 1650 5 1 1 3272
0 1651 7 1 2 3154 3273
0 1652 5 2 1 1651
0 1653 7 1 2 3161 3270
0 1654 5 1 1 1653
0 1655 7 1 2 3275 1654
0 1656 7 1 2 1645 1655
0 1657 5 1 1 1656
0 1658 7 1 2 3167 3265
0 1659 5 1 1 1658
0 1660 7 1 2 1657 1659
0 1661 7 1 2 1641 1660
0 1662 5 1 1 1661
0 1663 7 1 2 1637 1662
0 1664 7 1 2 1633 1663
0 1665 7 1 2 1628 1664
0 1666 7 1 2 1626 1665
0 1667 7 1 2 1622 1666
0 1668 7 1 2 1620 1667
0 1669 7 1 2 1616 1668
0 1670 7 1 2 1614 1669
0 1671 5 1 1 1670
0 1672 7 1 2 1610 1671
0 1673 7 1 2 1608 1672
0 1674 7 1 2 1602 1673
0 1675 7 1 2 1600 1674
0 1676 7 1 2 1596 1675
0 1677 7 1 2 1594 1676
0 1678 7 1 2 1590 1677
0 1679 7 1 2 1588 1678
0 1680 7 1 2 1584 1679
0 1681 7 1 2 3222 1680
0 1682 7 1 2 1571 1681
0 1683 5 1 1 1682
0 1684 7 2 2 3099 3111
0 1685 7 1 2 1487 3159
0 1686 5 1 1 1685
0 1687 7 2 2 1650 1686
0 1688 5 2 1 3279
0 1689 7 1 2 3134 3281
0 1690 5 1 1 1689
0 1691 7 2 2 3138 1690
0 1692 5 2 1 3283
0 1693 7 1 2 3123 3285
0 1694 5 1 1 1693
0 1695 7 3 2 3127 1694
0 1696 5 1 1 3287
0 1697 7 1 2 3115 3288
0 1698 5 1 1 1697
0 1699 7 1 2 3277 1698
0 1700 5 1 1 1699
0 1701 7 1 2 3102 1700
0 1702 5 2 1 1701
0 1703 7 1 2 3087 3290
0 1704 5 1 1 1703
0 1705 7 2 2 3091 1704
0 1706 5 2 1 3292
0 1707 7 1 2 3076 3294
0 1708 5 1 1 1707
0 1709 7 2 2 3080 1708
0 1710 5 2 1 3296
0 1711 7 1 2 3068 3298
0 1712 5 1 1 1711
0 1713 7 2 2 3065 1712
0 1714 5 2 1 3300
0 1715 7 1 2 3197 3302
0 1716 5 1 1 1715
0 1717 7 1 2 3192 1716
0 1718 7 1 2 3058 1717
0 1719 5 1 1 1718
0 1720 7 1 2 3200 1719
0 1721 7 1 2 3048 1720
0 1722 5 1 1 1721
0 1723 7 1 2 3045 1722
0 1724 7 2 2 3033 1723
0 1725 5 1 1 3304
0 1726 7 2 2 3036 1725
0 1727 5 2 1 3306
0 1728 7 1 2 3022 3308
0 1729 5 1 1 1728
0 1730 7 2 2 3025 1729
0 1731 5 1 1 3310
0 1732 7 1 2 3227 3311
0 1733 5 1 1 1732
0 1734 7 1 2 3225 1731
0 1735 5 1 1 1734
0 1736 7 1 2 3218 3015
0 1737 5 1 1 1736
0 1738 7 1 2 3232 3309
0 1739 5 1 1 1738
0 1740 7 1 2 3230 3307
0 1741 5 1 1 1740
0 1742 7 1 2 1739 1741
0 1743 5 1 1 1742
0 1744 7 1 2 3037 3305
0 1745 5 1 1 1744
0 1746 7 1 2 3049 3236
0 1747 5 1 1 1746
0 1748 7 1 2 3201 3240
0 1749 5 1 1 1748
0 1750 7 1 2 3195 3301
0 1751 5 1 1 1750
0 1752 7 1 2 3242 1751
0 1753 5 1 1 1752
0 1754 7 1 2 3190 3303
0 1755 5 1 1 1754
0 1756 7 1 2 3247 3297
0 1757 5 1 1 1756
0 1758 7 1 2 3245 3299
0 1759 5 1 1 1758
0 1760 7 1 2 3252 3293
0 1761 5 1 1 1760
0 1762 7 1 2 3250 3295
0 1763 5 1 1 1762
0 1764 7 1 2 3103 3257
0 1765 5 1 1 1764
0 1766 7 1 2 3255 3291
0 1767 5 1 1 1766
0 1768 7 1 2 3112 1696
0 1769 5 1 1 1768
0 1770 7 1 2 3259 1769
0 1771 5 1 1 1770
0 1772 7 1 2 3116 1771
0 1773 5 1 1 1772
0 1774 7 1 2 3261 3289
0 1775 5 1 1 1774
0 1776 7 1 2 3264 3284
0 1777 5 1 1 1776
0 1778 7 1 2 3269 3282
0 1779 5 1 1 1778
0 1780 7 1 2 3271 3280
0 1781 5 1 1 1780
0 1782 7 1 2 3276 1781
0 1783 7 1 2 1779 1782
0 1784 5 1 1 1783
0 1785 7 1 2 3266 3286
0 1786 5 1 1 1785
0 1787 7 1 2 1784 1786
0 1788 7 1 2 1777 1787
0 1789 5 1 1 1788
0 1790 7 1 2 1775 1789
0 1791 7 1 2 1773 1790
0 1792 7 1 2 1767 1791
0 1793 7 1 2 1765 1792
0 1794 7 1 2 1763 1793
0 1795 7 1 2 1761 1794
0 1796 7 1 2 1759 1795
0 1797 7 1 2 1757 1796
0 1798 5 1 1 1797
0 1799 7 1 2 1755 1798
0 1800 7 1 2 1753 1799
0 1801 7 1 2 1749 1800
0 1802 7 1 2 1747 1801
0 1803 7 1 2 1745 1802
0 1804 7 1 2 3011 1803
0 1805 7 1 2 1743 1804
0 1806 7 1 2 1737 1805
0 1807 7 1 2 1735 1806
0 1808 7 1 2 1733 1807
0 1809 7 1 2 1580 1808
0 1810 5 1 1 1809
0 1811 7 1 2 1683 1810
0 1812 7 1 2 2904 1811
0 1813 5 1 1 1812
0 1814 7 1 2 3135 3274
0 1815 7 1 2 3124 1814
0 1816 7 1 2 3278 1815
0 1817 7 1 2 3088 1816
0 1818 7 1 2 3077 1817
0 1819 7 1 2 3069 1818
0 1820 7 1 2 3203 1819
0 1821 7 1 2 3050 1820
0 1822 7 1 2 3038 1821
0 1823 7 1 2 3026 1822
0 1824 7 1 2 3220 1823
0 1825 7 1 2 3223 1824
0 1826 5 1 1 1825
0 1827 7 1 2 1199 1826
0 1828 5 1 1 1827
3 9999 7 0 2 1813 1828
