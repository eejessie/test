1 0 0 2 0
2 8 1 0
2 9 1 0
1 1 0 2 0
2 10 1 1
2 11 1 1
1 2 0 2 0
2 12 1 2
2 25 1 2
1 3 0 2 0
2 37 1 3
2 52 1 3
1 4 0 2 0
2 68 1 4
2 71 1 4
1 5 0 2 0
2 72 1 5
2 73 1 5
1 6 0 2 0
2 74 1 6
2 75 1 6
1 7 0 2 0
2 76 1 7
2 77 1 7
2 78 1 19
2 79 1 19
2 80 1 21
2 81 1 21
2 82 1 22
2 83 1 22
2 84 1 22
2 85 1 27
2 86 1 27
2 87 1 29
2 88 1 29
2 89 1 30
2 90 1 30
2 91 1 40
2 92 1 40
2 93 1 43
2 94 1 43
2 95 1 45
2 96 1 45
2 97 1 46
2 98 1 46
2 99 1 55
2 100 1 55
2 101 1 56
2 102 1 56
2 103 1 58
2 104 1 58
2 105 1 60
2 106 1 60
2 107 1 61
2 108 1 61
0 13 5 1 1 8
0 14 5 1 1 10
0 15 5 1 1 12
0 16 5 1 1 37
0 17 5 1 1 68
0 18 5 1 1 72
0 19 5 2 1 74
0 20 5 1 1 76
0 21 7 2 2 9 71
0 22 5 3 1 80
0 23 7 1 2 13 17
0 24 5 1 1 23
3 195 7 0 2 82 24
0 26 7 1 2 11 73
0 27 5 2 1 26
0 28 7 1 2 14 18
0 29 5 2 1 28
0 30 7 2 2 85 87
0 31 5 1 1 89
0 32 7 1 2 81 31
0 33 5 1 1 32
0 34 7 1 2 83 90
0 35 5 1 1 34
0 36 7 1 2 33 35
3 196 5 0 1 36
0 38 7 1 2 84 86
0 39 5 1 1 38
0 40 7 2 2 88 39
0 41 5 1 1 91
0 42 7 1 2 25 92
0 43 5 2 1 42
0 44 7 1 2 15 41
0 45 5 2 1 44
0 46 7 2 2 93 95
0 47 5 1 1 97
0 48 7 1 2 75 98
0 49 5 1 1 48
0 50 7 1 2 78 47
0 51 5 1 1 50
3 197 7 0 2 49 51
0 53 7 1 2 79 94
0 54 5 1 1 53
0 55 7 2 2 96 54
0 56 5 2 1 99
0 57 7 1 2 16 20
0 58 5 2 1 57
0 59 7 1 2 52 77
0 60 5 2 1 59
0 61 7 2 2 103 105
0 62 5 1 1 107
0 63 7 1 2 100 62
0 64 5 1 1 63
0 65 7 1 2 101 108
0 66 5 1 1 65
0 67 7 1 2 64 66
3 198 5 0 1 67
0 69 7 1 2 102 106
0 70 5 1 1 69
3 199 7 0 2 104 70
