1 0 0 8 0
2 32 1 0
2 2181 1 0
2 2182 1 0
2 2183 1 0
2 2184 1 0
2 2185 1 0
2 2186 1 0
2 2187 1 0
1 1 0 8 0
2 2188 1 1
2 2189 1 1
2 2190 1 1
2 2191 1 1
2 2192 1 1
2 2193 1 1
2 2194 1 1
2 2195 1 1
1 2 0 8 0
2 2196 1 2
2 2197 1 2
2 2198 1 2
2 2199 1 2
2 2200 1 2
2 2201 1 2
2 2202 1 2
2 2203 1 2
1 3 0 9 0
2 2204 1 3
2 2205 1 3
2 2206 1 3
2 2207 1 3
2 2208 1 3
2 2209 1 3
2 2210 1 3
2 2211 1 3
2 2212 1 3
1 4 0 8 0
2 2213 1 4
2 2214 1 4
2 2215 1 4
2 2216 1 4
2 2217 1 4
2 2218 1 4
2 2219 1 4
2 2220 1 4
1 5 0 9 0
2 2221 1 5
2 2222 1 5
2 2223 1 5
2 2224 1 5
2 2225 1 5
2 2226 1 5
2 2227 1 5
2 2228 1 5
2 2229 1 5
1 6 0 8 0
2 2230 1 6
2 2231 1 6
2 2232 1 6
2 2233 1 6
2 2234 1 6
2 2235 1 6
2 2236 1 6
2 2237 1 6
1 7 0 8 0
2 2238 1 7
2 2239 1 7
2 2240 1 7
2 2241 1 7
2 2242 1 7
2 2243 1 7
2 2244 1 7
2 2245 1 7
1 8 0 8 0
2 2246 1 8
2 2247 1 8
2 2248 1 8
2 2249 1 8
2 2250 1 8
2 2251 1 8
2 2252 1 8
2 2253 1 8
1 9 0 8 0
2 2254 1 9
2 2255 1 9
2 2256 1 9
2 2257 1 9
2 2258 1 9
2 2259 1 9
2 2260 1 9
2 2261 1 9
1 10 0 9 0
2 2262 1 10
2 2263 1 10
2 2264 1 10
2 2265 1 10
2 2266 1 10
2 2267 1 10
2 2268 1 10
2 2269 1 10
2 2270 1 10
1 11 0 8 0
2 2271 1 11
2 2272 1 11
2 2273 1 11
2 2274 1 11
2 2275 1 11
2 2276 1 11
2 2277 1 11
2 2278 1 11
1 12 0 8 0
2 2279 1 12
2 2280 1 12
2 2281 1 12
2 2282 1 12
2 2283 1 12
2 2284 1 12
2 2285 1 12
2 2286 1 12
1 13 0 8 0
2 2287 1 13
2 2288 1 13
2 2289 1 13
2 2290 1 13
2 2291 1 13
2 2292 1 13
2 2293 1 13
2 2294 1 13
1 14 0 8 0
2 2295 1 14
2 2296 1 14
2 2297 1 14
2 2298 1 14
2 2299 1 14
2 2300 1 14
2 2301 1 14
2 2302 1 14
1 15 0 8 0
2 2303 1 15
2 2304 1 15
2 2305 1 15
2 2306 1 15
2 2307 1 15
2 2308 1 15
2 2309 1 15
2 2310 1 15
1 16 0 2 0
2 2311 1 16
2 2312 1 16
1 17 0 2 0
2 2313 1 17
2 2314 1 17
1 18 0 2 0
2 2315 1 18
2 2316 1 18
1 19 0 2 0
2 2317 1 19
2 2318 1 19
1 20 0 2 0
2 2319 1 20
2 2320 1 20
1 21 0 2 0
2 2321 1 21
2 2322 1 21
1 22 0 2 0
2 2323 1 22
2 2324 1 22
1 23 0 2 0
2 2325 1 23
2 2326 1 23
1 24 0 2 0
2 2327 1 24
2 2328 1 24
1 25 0 2 0
2 2329 1 25
2 2330 1 25
1 26 0 2 0
2 2331 1 26
2 2332 1 26
1 27 0 2 0
2 2333 1 27
2 2334 1 27
1 28 0 2 0
2 2335 1 28
2 2336 1 28
1 29 0 2 0
2 2337 1 29
2 2338 1 29
1 30 0 2 0
2 2339 1 30
2 2340 1 30
1 31 0 2 0
2 2341 1 31
2 2342 1 31
2 2343 1 49
2 2344 1 49
2 2345 1 51
2 2346 1 51
2 2347 1 52
2 2348 1 52
2 2349 1 53
2 2350 1 53
2 2351 1 55
2 2352 1 55
2 2353 1 58
2 2354 1 58
2 2355 1 61
2 2356 1 61
2 2357 1 64
2 2358 1 64
2 2359 1 65
2 2360 1 65
2 2361 1 67
2 2362 1 67
2 2363 1 69
2 2364 1 69
2 2365 1 75
2 2366 1 75
2 2367 1 78
2 2368 1 78
2 2369 1 78
2 2370 1 81
2 2371 1 81
2 2372 1 82
2 2373 1 82
2 2374 1 83
2 2375 1 83
2 2376 1 85
2 2377 1 85
2 2378 1 88
2 2379 1 88
2 2380 1 89
2 2381 1 89
2 2382 1 93
2 2383 1 93
2 2384 1 96
2 2385 1 96
2 2386 1 97
2 2387 1 97
2 2388 1 101
2 2389 1 101
2 2390 1 104
2 2391 1 104
2 2392 1 105
2 2393 1 105
2 2394 1 109
2 2395 1 109
2 2396 1 112
2 2397 1 112
2 2398 1 113
2 2399 1 113
2 2400 1 115
2 2401 1 115
2 2402 1 118
2 2403 1 118
2 2404 1 119
2 2405 1 119
2 2406 1 123
2 2407 1 123
2 2408 1 126
2 2409 1 126
2 2410 1 127
2 2411 1 127
2 2412 1 131
2 2413 1 131
2 2414 1 134
2 2415 1 134
2 2416 1 135
2 2417 1 135
2 2418 1 139
2 2419 1 139
2 2420 1 142
2 2421 1 142
2 2422 1 143
2 2423 1 143
2 2424 1 147
2 2425 1 147
2 2426 1 150
2 2427 1 150
2 2428 1 151
2 2429 1 151
2 2430 1 155
2 2431 1 155
2 2432 1 158
2 2433 1 158
2 2434 1 159
2 2435 1 159
2 2436 1 163
2 2437 1 163
2 2438 1 166
2 2439 1 166
2 2440 1 167
2 2441 1 167
2 2442 1 171
2 2443 1 171
2 2444 1 174
2 2445 1 174
2 2446 1 175
2 2447 1 175
2 2448 1 177
2 2449 1 177
2 2450 1 179
2 2451 1 179
2 2452 1 181
2 2453 1 181
2 2454 1 182
2 2455 1 182
2 2456 1 183
2 2457 1 183
2 2458 1 184
2 2459 1 184
2 2460 1 186
2 2461 1 186
2 2462 1 187
2 2463 1 187
2 2464 1 191
2 2465 1 191
2 2466 1 194
2 2467 1 194
2 2468 1 195
2 2469 1 195
2 2470 1 199
2 2471 1 199
2 2472 1 202
2 2473 1 202
2 2474 1 203
2 2475 1 203
2 2476 1 207
2 2477 1 207
2 2478 1 210
2 2479 1 210
2 2480 1 211
2 2481 1 211
2 2482 1 215
2 2483 1 215
2 2484 1 218
2 2485 1 218
2 2486 1 219
2 2487 1 219
2 2488 1 223
2 2489 1 223
2 2490 1 226
2 2491 1 226
2 2492 1 227
2 2493 1 227
2 2494 1 231
2 2495 1 231
2 2496 1 234
2 2497 1 234
2 2498 1 235
2 2499 1 235
2 2500 1 239
2 2501 1 239
2 2502 1 242
2 2503 1 242
2 2504 1 243
2 2505 1 243
2 2506 1 245
2 2507 1 245
2 2508 1 248
2 2509 1 248
2 2510 1 251
2 2511 1 251
2 2512 1 255
2 2513 1 255
2 2514 1 258
2 2515 1 258
2 2516 1 259
2 2517 1 259
2 2518 1 263
2 2519 1 263
2 2520 1 266
2 2521 1 266
2 2522 1 267
2 2523 1 267
2 2524 1 269
2 2525 1 269
2 2526 1 272
2 2527 1 272
2 2528 1 273
2 2529 1 273
2 2530 1 275
2 2531 1 275
2 2532 1 281
2 2533 1 281
2 2534 1 284
2 2535 1 284
2 2536 1 287
2 2537 1 287
2 2538 1 290
2 2539 1 290
2 2540 1 293
2 2541 1 293
2 2542 1 297
2 2543 1 297
2 2544 1 300
2 2545 1 300
2 2546 1 301
2 2547 1 301
2 2548 1 305
2 2549 1 305
2 2550 1 308
2 2551 1 308
2 2552 1 309
2 2553 1 309
2 2554 1 311
2 2555 1 311
2 2556 1 314
2 2557 1 314
2 2558 1 317
2 2559 1 317
2 2560 1 321
2 2561 1 321
2 2562 1 324
2 2563 1 324
2 2564 1 325
2 2565 1 325
2 2566 1 329
2 2567 1 329
2 2568 1 332
2 2569 1 332
2 2570 1 333
2 2571 1 333
2 2572 1 337
2 2573 1 337
2 2574 1 340
2 2575 1 340
2 2576 1 341
2 2577 1 341
2 2578 1 345
2 2579 1 345
2 2580 1 348
2 2581 1 348
2 2582 1 349
2 2583 1 349
2 2584 1 353
2 2585 1 353
2 2586 1 356
2 2587 1 356
2 2588 1 357
2 2589 1 357
2 2590 1 359
2 2591 1 359
2 2592 1 362
2 2593 1 362
2 2594 1 363
2 2595 1 363
2 2596 1 367
2 2597 1 367
2 2598 1 370
2 2599 1 370
2 2600 1 371
2 2601 1 371
2 2602 1 373
2 2603 1 373
2 2604 1 375
2 2605 1 375
2 2606 1 378
2 2607 1 378
2 2608 1 379
2 2609 1 379
2 2610 1 381
2 2611 1 381
2 2612 1 383
2 2613 1 383
2 2614 1 385
2 2615 1 385
2 2616 1 387
2 2617 1 387
2 2618 1 388
2 2619 1 388
2 2620 1 389
2 2621 1 389
2 2622 1 390
2 2623 1 390
2 2624 1 391
2 2625 1 391
2 2626 1 392
2 2627 1 392
2 2628 1 393
2 2629 1 393
2 2630 1 394
2 2631 1 394
2 2632 1 396
2 2633 1 396
2 2634 1 399
2 2635 1 399
2 2636 1 403
2 2637 1 403
2 2638 1 406
2 2639 1 406
2 2640 1 409
2 2641 1 409
2 2642 1 413
2 2643 1 413
2 2644 1 416
2 2645 1 416
2 2646 1 417
2 2647 1 417
2 2648 1 420
2 2649 1 420
2 2650 1 421
2 2651 1 421
2 2652 1 425
2 2653 1 425
2 2654 1 428
2 2655 1 428
2 2656 1 429
2 2657 1 429
2 2658 1 433
2 2659 1 433
2 2660 1 436
2 2661 1 436
2 2662 1 437
2 2663 1 437
2 2664 1 441
2 2665 1 441
2 2666 1 444
2 2667 1 444
2 2668 1 447
2 2669 1 447
2 2670 1 451
2 2671 1 451
2 2672 1 454
2 2673 1 454
2 2674 1 457
2 2675 1 457
2 2676 1 461
2 2677 1 461
2 2678 1 464
2 2679 1 464
2 2680 1 465
2 2681 1 465
2 2682 1 467
2 2683 1 467
2 2684 1 470
2 2685 1 470
2 2686 1 471
2 2687 1 471
2 2688 1 475
2 2689 1 475
2 2690 1 478
2 2691 1 478
2 2692 1 479
2 2693 1 479
2 2694 1 483
2 2695 1 483
2 2696 1 486
2 2697 1 486
2 2698 1 487
2 2699 1 487
2 2700 1 491
2 2701 1 491
2 2702 1 494
2 2703 1 494
2 2704 1 495
2 2705 1 495
2 2706 1 499
2 2707 1 499
2 2708 1 502
2 2709 1 502
2 2710 1 503
2 2711 1 503
2 2712 1 507
2 2713 1 507
2 2714 1 510
2 2715 1 510
2 2716 1 511
2 2717 1 511
2 2718 1 513
2 2719 1 513
2 2720 1 519
2 2721 1 519
2 2722 1 522
2 2723 1 522
2 2724 1 525
2 2725 1 525
2 2726 1 528
2 2727 1 528
2 2728 1 531
2 2729 1 531
2 2730 1 535
2 2731 1 535
2 2732 1 538
2 2733 1 538
2 2734 1 539
2 2735 1 539
2 2736 1 543
2 2737 1 543
2 2738 1 546
2 2739 1 546
2 2740 1 547
2 2741 1 547
2 2742 1 551
2 2743 1 551
2 2744 1 554
2 2745 1 554
2 2746 1 555
2 2747 1 555
2 2748 1 559
2 2749 1 559
2 2750 1 562
2 2751 1 562
2 2752 1 563
2 2753 1 563
2 2754 1 567
2 2755 1 567
2 2756 1 570
2 2757 1 570
2 2758 1 571
2 2759 1 571
2 2760 1 575
2 2761 1 575
2 2762 1 578
2 2763 1 578
2 2764 1 579
2 2765 1 579
2 2766 1 583
2 2767 1 583
2 2768 1 586
2 2769 1 586
2 2770 1 587
2 2771 1 587
2 2772 1 589
2 2773 1 589
2 2774 1 592
2 2775 1 592
2 2776 1 595
2 2777 1 595
2 2778 1 599
2 2779 1 599
2 2780 1 602
2 2781 1 602
2 2782 1 603
2 2783 1 603
2 2784 1 607
2 2785 1 607
2 2786 1 610
2 2787 1 610
2 2788 1 611
2 2789 1 611
2 2790 1 615
2 2791 1 615
2 2792 1 618
2 2793 1 618
2 2794 1 619
2 2795 1 619
2 2796 1 623
2 2797 1 623
2 2798 1 626
2 2799 1 626
2 2800 1 627
2 2801 1 627
2 2802 1 633
2 2803 1 633
2 2804 1 636
2 2805 1 636
2 2806 1 637
2 2807 1 637
2 2808 1 641
2 2809 1 641
2 2810 1 644
2 2811 1 644
2 2812 1 645
2 2813 1 645
2 2814 1 649
2 2815 1 649
2 2816 1 652
2 2817 1 652
2 2818 1 653
2 2819 1 653
2 2820 1 657
2 2821 1 657
2 2822 1 660
2 2823 1 660
2 2824 1 661
2 2825 1 661
2 2826 1 663
2 2827 1 663
2 2828 1 666
2 2829 1 666
2 2830 1 669
2 2831 1 669
2 2832 1 673
2 2833 1 673
2 2834 1 676
2 2835 1 676
2 2836 1 677
2 2837 1 677
2 2838 1 681
2 2839 1 681
2 2840 1 684
2 2841 1 684
2 2842 1 687
2 2843 1 687
2 2844 1 689
2 2845 1 689
2 2846 1 691
2 2847 1 691
2 2848 1 693
2 2849 1 693
2 2850 1 695
2 2851 1 695
2 2852 1 697
2 2853 1 697
2 2854 1 699
2 2855 1 699
2 2856 1 700
2 2857 1 700
2 2858 1 701
2 2859 1 701
2 2860 1 701
2 2861 1 704
2 2862 1 704
2 2863 1 707
2 2864 1 707
2 2865 1 715
2 2866 1 715
2 2867 1 718
2 2868 1 718
2 2869 1 719
2 2870 1 719
2 2871 1 723
2 2872 1 723
2 2873 1 726
2 2874 1 726
2 2875 1 729
2 2876 1 729
2 2877 1 729
2 2878 1 730
2 2879 1 730
2 2880 1 731
2 2881 1 731
2 2882 1 733
2 2883 1 733
2 2884 1 735
2 2885 1 735
2 2886 1 736
2 2887 1 736
2 2888 1 738
2 2889 1 738
2 2890 1 739
2 2891 1 739
2 2892 1 743
2 2893 1 743
2 2894 1 746
2 2895 1 746
2 2896 1 747
2 2897 1 747
2 2898 1 751
2 2899 1 751
2 2900 1 754
2 2901 1 754
2 2902 1 755
2 2903 1 755
2 2904 1 759
2 2905 1 759
2 2906 1 762
2 2907 1 762
2 2908 1 763
2 2909 1 763
2 2910 1 767
2 2911 1 767
2 2912 1 770
2 2913 1 770
2 2914 1 771
2 2915 1 771
2 2916 1 775
2 2917 1 775
2 2918 1 778
2 2919 1 778
2 2920 1 779
2 2921 1 779
2 2922 1 783
2 2923 1 783
2 2924 1 786
2 2925 1 786
2 2926 1 787
2 2927 1 787
2 2928 1 791
2 2929 1 791
2 2930 1 794
2 2931 1 794
2 2932 1 795
2 2933 1 795
2 2934 1 799
2 2935 1 799
2 2936 1 802
2 2937 1 802
2 2938 1 803
2 2939 1 803
2 2940 1 807
2 2941 1 807
2 2942 1 810
2 2943 1 810
2 2944 1 811
2 2945 1 811
2 2946 1 815
2 2947 1 815
2 2948 1 818
2 2949 1 818
2 2950 1 819
2 2951 1 819
2 2952 1 823
2 2953 1 823
2 2954 1 826
2 2955 1 826
2 2956 1 827
2 2957 1 827
2 2958 1 827
2 2959 1 828
2 2960 1 828
2 2961 1 829
2 2962 1 829
2 2963 1 831
2 2964 1 831
2 2965 1 834
2 2966 1 834
2 2967 1 835
2 2968 1 835
2 2969 1 835
2 2970 1 836
2 2971 1 836
2 2972 1 838
2 2973 1 838
2 2974 1 838
2 2975 1 838
2 2976 1 838
2 2977 1 840
2 2978 1 840
2 2979 1 840
2 2980 1 840
2 2981 1 840
2 2982 1 843
2 2983 1 843
2 2984 1 843
2 2985 1 844
2 2986 1 844
2 2987 1 846
2 2988 1 846
2 2989 1 846
2 2990 1 849
2 2991 1 849
2 2992 1 849
2 2993 1 849
2 2994 1 850
2 2995 1 850
2 2996 1 850
2 2997 1 852
2 2998 1 852
2 2999 1 852
2 3000 1 855
2 3001 1 855
2 3002 1 855
2 3003 1 855
2 3004 1 856
2 3005 1 856
2 3006 1 856
2 3007 1 858
2 3008 1 858
2 3009 1 858
2 3010 1 861
2 3011 1 861
2 3012 1 861
2 3013 1 861
2 3014 1 862
2 3015 1 862
2 3016 1 862
2 3017 1 864
2 3018 1 864
2 3019 1 864
2 3020 1 867
2 3021 1 867
2 3022 1 867
2 3023 1 867
2 3024 1 868
2 3025 1 868
2 3026 1 868
2 3027 1 870
2 3028 1 870
2 3029 1 870
2 3030 1 873
2 3031 1 873
2 3032 1 873
2 3033 1 873
2 3034 1 874
2 3035 1 874
2 3036 1 874
2 3037 1 876
2 3038 1 876
2 3039 1 876
2 3040 1 879
2 3041 1 879
2 3042 1 879
2 3043 1 879
2 3044 1 880
2 3045 1 880
2 3046 1 880
2 3047 1 882
2 3048 1 882
2 3049 1 882
2 3050 1 884
2 3051 1 884
2 3052 1 884
2 3053 1 887
2 3054 1 887
2 3055 1 887
2 3056 1 887
2 3057 1 888
2 3058 1 888
2 3059 1 888
2 3060 1 890
2 3061 1 890
2 3062 1 890
2 3063 1 893
2 3064 1 893
2 3065 1 893
2 3066 1 893
2 3067 1 894
2 3068 1 894
2 3069 1 894
2 3070 1 896
2 3071 1 896
2 3072 1 896
2 3073 1 898
2 3074 1 898
2 3075 1 898
2 3076 1 901
2 3077 1 901
2 3078 1 901
2 3079 1 901
2 3080 1 902
2 3081 1 902
2 3082 1 902
2 3083 1 904
2 3084 1 904
2 3085 1 904
2 3086 1 907
2 3087 1 907
2 3088 1 907
2 3089 1 907
2 3090 1 908
2 3091 1 908
2 3092 1 908
2 3093 1 910
2 3094 1 910
2 3095 1 910
2 3096 1 913
2 3097 1 913
2 3098 1 913
2 3099 1 913
2 3100 1 914
2 3101 1 914
2 3102 1 914
2 3103 1 916
2 3104 1 916
2 3105 1 916
2 3106 1 919
2 3107 1 919
2 3108 1 919
2 3109 1 920
2 3110 1 920
2 3111 1 920
2 3112 1 922
2 3113 1 922
2 3114 1 922
2 3115 1 924
2 3116 1 924
2 3117 1 924
2 3118 1 925
2 3119 1 925
2 3120 1 927
2 3121 1 927
2 3122 1 927
2 3123 1 927
2 3124 1 928
2 3125 1 928
2 3126 1 930
2 3127 1 930
2 3128 1 930
2 3129 1 932
2 3130 1 932
2 3131 1 932
2 3132 1 933
2 3133 1 933
2 3134 1 933
2 3135 1 934
2 3136 1 934
2 3137 1 934
2 3138 1 935
2 3139 1 935
2 3140 1 936
2 3141 1 936
2 3142 1 936
2 3143 1 939
2 3144 1 939
2 3145 1 940
2 3146 1 940
2 3147 1 943
2 3148 1 943
2 3149 1 944
2 3150 1 944
2 3151 1 946
2 3152 1 946
2 3153 1 946
2 3154 1 949
2 3155 1 949
2 3156 1 950
2 3157 1 950
2 3158 1 952
2 3159 1 952
2 3160 1 952
2 3161 1 955
2 3162 1 955
2 3163 1 956
2 3164 1 956
2 3165 1 958
2 3166 1 958
2 3167 1 958
2 3168 1 961
2 3169 1 961
2 3170 1 962
2 3171 1 962
2 3172 1 965
2 3173 1 965
2 3174 1 966
2 3175 1 966
2 3176 1 968
2 3177 1 968
2 3178 1 968
2 3179 1 971
2 3180 1 971
2 3181 1 972
2 3182 1 972
2 3183 1 975
2 3184 1 975
2 3185 1 976
2 3186 1 976
2 3187 1 978
2 3188 1 978
2 3189 1 978
2 3190 1 981
2 3191 1 981
2 3192 1 982
2 3193 1 982
2 3194 1 984
2 3195 1 984
2 3196 1 984
2 3197 1 987
2 3198 1 987
2 3199 1 988
2 3200 1 988
2 3201 1 990
2 3202 1 990
2 3203 1 990
2 3204 1 993
2 3205 1 993
2 3206 1 994
2 3207 1 994
2 3208 1 996
2 3209 1 996
2 3210 1 996
2 3211 1 999
2 3212 1 999
2 3213 1 1000
2 3214 1 1000
2 3215 1 1002
2 3216 1 1002
2 3217 1 1002
2 3218 1 1005
2 3219 1 1005
2 3220 1 1006
2 3221 1 1006
2 3222 1 1008
2 3223 1 1008
2 3224 1 1008
2 3225 1 1011
2 3226 1 1011
2 3227 1 1011
2 3228 1 1011
2 3229 1 1012
2 3230 1 1012
2 3231 1 1015
2 3232 1 1015
2 3233 1 1015
2 3234 1 1017
2 3235 1 1017
2 3236 1 1017
2 3237 1 1018
2 3238 1 1018
2 3239 1 1023
2 3240 1 1023
2 3241 1 1023
2 3242 1 1024
2 3243 1 1024
2 3244 1 1026
2 3245 1 1026
2 3246 1 1027
2 3247 1 1027
2 3248 1 1027
2 3249 1 1028
2 3250 1 1028
2 3251 1 1033
2 3252 1 1033
2 3253 1 1033
2 3254 1 1034
2 3255 1 1034
2 3256 1 1035
2 3257 1 1035
2 3258 1 1035
2 3259 1 1036
2 3260 1 1036
2 3261 1 1041
2 3262 1 1041
2 3263 1 1044
2 3264 1 1044
2 3265 1 1045
2 3266 1 1045
2 3267 1 1045
2 3268 1 1046
2 3269 1 1046
2 3270 1 1051
2 3271 1 1051
2 3272 1 1051
2 3273 1 1052
2 3274 1 1052
2 3275 1 1054
2 3276 1 1054
2 3277 1 1055
2 3278 1 1055
2 3279 1 1055
2 3280 1 1056
2 3281 1 1056
2 3282 1 1061
2 3283 1 1061
2 3284 1 1061
2 3285 1 1062
2 3286 1 1062
2 3287 1 1064
2 3288 1 1064
2 3289 1 1065
2 3290 1 1065
2 3291 1 1065
2 3292 1 1066
2 3293 1 1066
2 3294 1 1071
2 3295 1 1071
2 3296 1 1071
2 3297 1 1072
2 3298 1 1072
2 3299 1 1074
2 3300 1 1074
2 3301 1 1075
2 3302 1 1075
2 3303 1 1075
2 3304 1 1076
2 3305 1 1076
2 3306 1 1081
2 3307 1 1081
2 3308 1 1081
2 3309 1 1082
2 3310 1 1082
2 3311 1 1084
2 3312 1 1084
2 3313 1 1085
2 3314 1 1085
2 3315 1 1085
2 3316 1 1086
2 3317 1 1086
2 3318 1 1091
2 3319 1 1091
2 3320 1 1091
2 3321 1 1092
2 3322 1 1092
2 3323 1 1094
2 3324 1 1094
2 3325 1 1095
2 3326 1 1095
2 3327 1 1095
2 3328 1 1096
2 3329 1 1096
2 3330 1 1101
2 3331 1 1101
2 3332 1 1101
2 3333 1 1102
2 3334 1 1102
2 3335 1 1104
2 3336 1 1104
2 3337 1 1105
2 3338 1 1105
2 3339 1 1105
2 3340 1 1106
2 3341 1 1106
2 3342 1 1111
2 3343 1 1111
2 3344 1 1111
2 3345 1 1112
2 3346 1 1112
2 3347 1 1114
2 3348 1 1114
2 3349 1 1115
2 3350 1 1115
2 3351 1 1115
2 3352 1 1116
2 3353 1 1116
2 3354 1 1121
2 3355 1 1121
2 3356 1 1121
2 3357 1 1122
2 3358 1 1122
2 3359 1 1124
2 3360 1 1124
2 3361 1 1125
2 3362 1 1125
2 3363 1 1125
2 3364 1 1126
2 3365 1 1126
2 3366 1 1131
2 3367 1 1131
2 3368 1 1131
2 3369 1 1132
2 3370 1 1132
2 3371 1 1134
2 3372 1 1134
2 3373 1 1135
2 3374 1 1135
2 3375 1 1135
2 3376 1 1136
2 3377 1 1136
2 3378 1 1141
2 3379 1 1141
2 3380 1 1141
2 3381 1 1142
2 3382 1 1142
2 3383 1 1144
2 3384 1 1144
2 3385 1 1145
2 3386 1 1145
2 3387 1 1145
2 3388 1 1146
2 3389 1 1146
2 3390 1 1151
2 3391 1 1151
2 3392 1 1151
2 3393 1 1152
2 3394 1 1152
2 3395 1 1154
2 3396 1 1154
2 3397 1 1155
2 3398 1 1155
2 3399 1 1155
2 3400 1 1156
2 3401 1 1156
2 3402 1 1161
2 3403 1 1161
2 3404 1 1162
2 3405 1 1162
2 3406 1 1164
2 3407 1 1164
2 3408 1 1165
2 3409 1 1165
2 3410 1 1165
2 3411 1 1166
2 3412 1 1166
2 3413 1 1166
2 3414 1 1167
2 3415 1 1167
2 3416 1 1167
2 3417 1 1168
2 3418 1 1168
2 3419 1 1169
2 3420 1 1169
2 3421 1 1170
2 3422 1 1170
2 3423 1 1173
2 3424 1 1173
2 3425 1 1176
2 3426 1 1176
2 3427 1 1177
2 3428 1 1177
2 3429 1 1181
2 3430 1 1181
2 3431 1 1184
2 3432 1 1184
2 3433 1 1185
2 3434 1 1185
2 3435 1 1189
2 3436 1 1189
2 3437 1 1192
2 3438 1 1192
2 3439 1 1193
2 3440 1 1193
2 3441 1 1197
2 3442 1 1197
2 3443 1 1200
2 3444 1 1200
2 3445 1 1201
2 3446 1 1201
2 3447 1 1205
2 3448 1 1205
2 3449 1 1208
2 3450 1 1208
2 3451 1 1209
2 3452 1 1209
2 3453 1 1213
2 3454 1 1213
2 3455 1 1216
2 3456 1 1216
2 3457 1 1217
2 3458 1 1217
2 3459 1 1221
2 3460 1 1221
2 3461 1 1224
2 3462 1 1224
2 3463 1 1225
2 3464 1 1225
2 3465 1 1229
2 3466 1 1229
2 3467 1 1232
2 3468 1 1232
2 3469 1 1233
2 3470 1 1233
2 3471 1 1237
2 3472 1 1237
2 3473 1 1240
2 3474 1 1240
2 3475 1 1241
2 3476 1 1241
2 3477 1 1245
2 3478 1 1245
2 3479 1 1248
2 3480 1 1248
2 3481 1 1249
2 3482 1 1249
2 3483 1 1253
2 3484 1 1253
2 3485 1 1256
2 3486 1 1256
2 3487 1 1257
2 3488 1 1257
2 3489 1 1261
2 3490 1 1261
2 3491 1 1264
2 3492 1 1264
2 3493 1 1265
2 3494 1 1265
2 3495 1 1269
2 3496 1 1269
2 3497 1 1272
2 3498 1 1272
2 3499 1 1273
2 3500 1 1273
2 3501 1 1277
2 3502 1 1277
2 3503 1 1280
2 3504 1 1280
2 3505 1 1281
2 3506 1 1281
2 3507 1 1287
2 3508 1 1287
2 3509 1 1290
2 3510 1 1290
2 3511 1 1292
2 3512 1 1292
2 3513 1 1296
2 3514 1 1296
2 3515 1 1298
2 3516 1 1298
2 3517 1 1300
2 3518 1 1300
2 3519 1 1302
2 3520 1 1302
2 3521 1 1304
2 3522 1 1304
2 3523 1 1306
2 3524 1 1306
2 3525 1 1308
2 3526 1 1308
2 3527 1 1310
2 3528 1 1310
2 3529 1 1312
2 3530 1 1312
2 3531 1 1314
2 3532 1 1314
2 3533 1 1316
2 3534 1 1316
2 3535 1 1318
2 3536 1 1318
2 3537 1 1320
2 3538 1 1320
2 3539 1 1323
2 3540 1 1323
2 3541 1 1327
2 3542 1 1327
2 3543 1 1328
2 3544 1 1328
2 3545 1 1330
2 3546 1 1330
2 3547 1 1331
2 3548 1 1331
2 3549 1 1335
2 3550 1 1335
2 3551 1 1338
2 3552 1 1338
2 3553 1 1339
2 3554 1 1339
2 3555 1 1343
2 3556 1 1343
2 3557 1 1346
2 3558 1 1346
2 3559 1 1347
2 3560 1 1347
2 3561 1 1351
2 3562 1 1351
2 3563 1 1354
2 3564 1 1354
2 3565 1 1355
2 3566 1 1355
2 3567 1 1359
2 3568 1 1359
2 3569 1 1362
2 3570 1 1362
2 3571 1 1363
2 3572 1 1363
2 3573 1 1367
2 3574 1 1367
2 3575 1 1370
2 3576 1 1370
2 3577 1 1371
2 3578 1 1371
2 3579 1 1375
2 3580 1 1375
2 3581 1 1378
2 3582 1 1378
2 3583 1 1379
2 3584 1 1379
2 3585 1 1383
2 3586 1 1383
2 3587 1 1386
2 3588 1 1386
2 3589 1 1387
2 3590 1 1387
2 3591 1 1391
2 3592 1 1391
2 3593 1 1394
2 3594 1 1394
2 3595 1 1395
2 3596 1 1395
2 3597 1 1399
2 3598 1 1399
2 3599 1 1402
2 3600 1 1402
2 3601 1 1403
2 3602 1 1403
2 3603 1 1407
2 3604 1 1407
2 3605 1 1410
2 3606 1 1410
2 3607 1 1411
2 3608 1 1411
2 3609 1 1415
2 3610 1 1415
2 3611 1 1418
2 3612 1 1418
2 3613 1 1419
2 3614 1 1419
2 3615 1 1423
2 3616 1 1423
2 3617 1 1425
2 3618 1 1425
2 3619 1 1426
2 3620 1 1426
2 3621 1 1429
2 3622 1 1429
2 3623 1 1429
2 3624 1 1429
2 3625 1 1429
2 3626 1 1435
2 3627 1 1435
2 3628 1 1438
2 3629 1 1438
2 3630 1 1438
2 3631 1 1439
2 3632 1 1439
2 3633 1 1447
2 3634 1 1447
2 3635 1 1447
2 3636 1 1448
2 3637 1 1448
2 3638 1 1451
2 3639 1 1451
2 3640 1 1459
2 3641 1 1459
2 3642 1 1459
2 3643 1 1460
2 3644 1 1460
2 3645 1 1463
2 3646 1 1463
2 3647 1 1471
2 3648 1 1471
2 3649 1 1471
2 3650 1 1472
2 3651 1 1472
2 3652 1 1475
2 3653 1 1475
2 3654 1 1483
2 3655 1 1483
2 3656 1 1483
2 3657 1 1484
2 3658 1 1484
2 3659 1 1487
2 3660 1 1487
2 3661 1 1495
2 3662 1 1495
2 3663 1 1495
2 3664 1 1496
2 3665 1 1496
2 3666 1 1499
2 3667 1 1499
2 3668 1 1507
2 3669 1 1507
2 3670 1 1507
2 3671 1 1508
2 3672 1 1508
2 3673 1 1511
2 3674 1 1511
2 3675 1 1519
2 3676 1 1519
2 3677 1 1520
2 3678 1 1520
2 3679 1 1523
2 3680 1 1523
2 3681 1 1531
2 3682 1 1531
2 3683 1 1531
2 3684 1 1532
2 3685 1 1532
2 3686 1 1535
2 3687 1 1535
2 3688 1 1543
2 3689 1 1543
2 3690 1 1544
2 3691 1 1544
2 3692 1 1547
2 3693 1 1547
2 3694 1 1559
2 3695 1 1559
2 3696 1 1559
2 3697 1 1560
2 3698 1 1560
2 3699 1 1563
2 3700 1 1563
2 3701 1 1564
2 3702 1 1564
2 3703 1 1567
2 3704 1 1567
2 3705 1 1567
2 3706 1 1571
2 3707 1 1571
2 3708 1 1575
2 3709 1 1575
2 3710 1 1575
2 3711 1 1579
2 3712 1 1579
2 3713 1 1581
2 3714 1 1581
2 3715 1 1589
2 3716 1 1589
2 3717 1 1590
2 3718 1 1590
2 3719 1 1593
2 3720 1 1593
2 3721 1 1596
2 3722 1 1596
2 3723 1 1601
2 3724 1 1601
2 3725 1 1605
2 3726 1 1605
2 3727 1 1613
2 3728 1 1613
2 3729 1 1621
2 3730 1 1621
2 3731 1 1629
2 3732 1 1629
2 3733 1 1640
2 3734 1 1640
2 3735 1 1698
2 3736 1 1698
2 3737 1 1699
2 3738 1 1699
2 3739 1 1700
2 3740 1 1700
2 3741 1 1703
2 3742 1 1703
2 3743 1 1704
2 3744 1 1704
2 3745 1 1707
2 3746 1 1707
2 3747 1 1708
2 3748 1 1708
2 3749 1 1711
2 3750 1 1711
2 3751 1 1712
2 3752 1 1712
2 3753 1 1715
2 3754 1 1715
2 3755 1 1716
2 3756 1 1716
2 3757 1 1719
2 3758 1 1719
2 3759 1 1720
2 3760 1 1720
2 3761 1 1723
2 3762 1 1723
2 3763 1 1724
2 3764 1 1724
2 3765 1 1727
2 3766 1 1727
2 3767 1 1728
2 3768 1 1728
2 3769 1 1731
2 3770 1 1731
2 3771 1 1732
2 3772 1 1732
2 3773 1 1735
2 3774 1 1735
2 3775 1 1736
2 3776 1 1736
2 3777 1 1739
2 3778 1 1739
2 3779 1 1740
2 3780 1 1740
2 3781 1 1743
2 3782 1 1743
2 3783 1 1744
2 3784 1 1744
2 3785 1 1747
2 3786 1 1747
2 3787 1 1748
2 3788 1 1748
2 3789 1 1751
2 3790 1 1751
2 3791 1 1751
2 3792 1 1752
2 3793 1 1752
2 3794 1 1752
2 3795 1 1755
2 3796 1 1755
2 3797 1 1755
2 3798 1 1756
2 3799 1 1756
2 3800 1 1763
2 3801 1 1763
2 3802 1 1763
2 3803 1 1764
2 3804 1 1764
2 3805 1 1769
2 3806 1 1769
2 3807 1 1769
2 3808 1 1770
2 3809 1 1770
2 3810 1 1772
2 3811 1 1772
2 3812 1 1777
2 3813 1 1777
2 3814 1 1777
2 3815 1 1778
2 3816 1 1778
2 3817 1 1783
2 3818 1 1783
2 3819 1 1783
2 3820 1 1784
2 3821 1 1784
2 3822 1 1786
2 3823 1 1786
2 3824 1 1791
2 3825 1 1791
2 3826 1 1791
2 3827 1 1792
2 3828 1 1792
2 3829 1 1794
2 3830 1 1794
2 3831 1 1799
2 3832 1 1799
2 3833 1 1799
2 3834 1 1800
2 3835 1 1800
2 3836 1 1802
2 3837 1 1802
2 3838 1 1807
2 3839 1 1807
2 3840 1 1807
2 3841 1 1808
2 3842 1 1808
2 3843 1 1810
2 3844 1 1810
2 3845 1 1815
2 3846 1 1815
2 3847 1 1815
2 3848 1 1816
2 3849 1 1816
2 3850 1 1818
2 3851 1 1818
2 3852 1 1823
2 3853 1 1823
2 3854 1 1823
2 3855 1 1824
2 3856 1 1824
2 3857 1 1826
2 3858 1 1826
2 3859 1 1831
2 3860 1 1831
2 3861 1 1831
2 3862 1 1832
2 3863 1 1832
2 3864 1 1834
2 3865 1 1834
2 3866 1 1837
2 3867 1 1837
2 3868 1 1837
2 3869 1 1840
2 3870 1 1840
2 3871 1 1841
2 3872 1 1841
2 3873 1 1842
2 3874 1 1842
2 3875 1 1845
2 3876 1 1845
2 3877 1 1848
2 3878 1 1848
2 3879 1 1849
2 3880 1 1849
2 3881 1 1853
2 3882 1 1853
2 3883 1 1856
2 3884 1 1856
2 3885 1 1857
2 3886 1 1857
2 3887 1 1861
2 3888 1 1861
2 3889 1 1864
2 3890 1 1864
2 3891 1 1865
2 3892 1 1865
2 3893 1 1869
2 3894 1 1869
2 3895 1 1872
2 3896 1 1872
2 3897 1 1873
2 3898 1 1873
2 3899 1 1877
2 3900 1 1877
2 3901 1 1880
2 3902 1 1880
2 3903 1 1881
2 3904 1 1881
2 3905 1 1885
2 3906 1 1885
2 3907 1 1888
2 3908 1 1888
2 3909 1 1889
2 3910 1 1889
2 3911 1 1893
2 3912 1 1893
2 3913 1 1896
2 3914 1 1896
2 3915 1 1897
2 3916 1 1897
2 3917 1 1901
2 3918 1 1901
2 3919 1 1904
2 3920 1 1904
2 3921 1 1905
2 3922 1 1905
2 3923 1 1909
2 3924 1 1909
2 3925 1 1912
2 3926 1 1912
2 3927 1 1913
2 3928 1 1913
2 3929 1 1919
2 3930 1 1919
2 3931 1 1919
2 3932 1 1920
2 3933 1 1920
2 3934 1 1922
2 3935 1 1922
2 3936 1 1925
2 3937 1 1925
2 3938 1 1928
2 3939 1 1928
2 3940 1 1931
2 3941 1 1931
2 3942 1 1937
2 3943 1 1937
2 3944 1 1945
2 3945 1 1945
2 3946 1 1951
2 3947 1 1951
2 3948 1 1955
2 3949 1 1955
2 3950 1 1963
2 3951 1 1963
2 3952 1 1967
2 3953 1 1967
2 3954 1 1975
2 3955 1 1975
2 3956 1 1979
2 3957 1 1979
2 3958 1 1987
2 3959 1 1987
2 3960 1 1997
2 3961 1 1997
2 3962 1 2014
2 3963 1 2014
2 3964 1 2026
2 3965 1 2026
2 3966 1 2038
2 3967 1 2038
2 3968 1 2061
2 3969 1 2061
2 3970 1 2067
2 3971 1 2067
2 3972 1 2067
2 3973 1 2068
2 3974 1 2068
2 3975 1 2070
2 3976 1 2070
2 3977 1 2073
2 3978 1 2073
2 3979 1 2076
2 3980 1 2076
2 3981 1 2079
2 3982 1 2079
2 3983 1 2086
2 3984 1 2086
2 3985 1 2092
2 3986 1 2092
2 3987 1 2092
2 3988 1 2093
2 3989 1 2093
2 3990 1 2095
2 3991 1 2095
2 3992 1 2098
2 3993 1 2098
2 3994 1 2101
2 3995 1 2101
2 3996 1 2104
2 3997 1 2104
2 3998 1 2113
2 3999 1 2113
2 4000 1 2119
2 4001 1 2119
2 4002 1 2122
2 4003 1 2122
2 4004 1 2125
2 4005 1 2125
2 4006 1 2128
2 4007 1 2128
2 4008 1 2131
2 4009 1 2131
2 4010 1 2140
2 4011 1 2140
2 4012 1 2146
2 4013 1 2146
2 4014 1 2155
2 4015 1 2155
2 4016 1 2156
2 4017 1 2156
2 4018 1 2162
2 4019 1 2162
0 33 5 1 1 2311
0 34 5 1 1 2313
0 35 5 1 1 2315
0 36 5 1 1 2317
0 37 5 1 1 2319
0 38 5 1 1 2321
0 39 5 1 1 2323
0 40 5 1 1 2325
0 41 5 1 1 2327
0 42 5 1 1 2329
0 43 5 1 1 2331
0 44 5 1 1 2333
0 45 5 1 1 2335
0 46 5 1 1 2337
0 47 5 1 1 2339
0 48 5 1 1 2341
0 49 7 2 2 2238 2303
0 50 5 1 1 2343
0 51 7 2 2 2230 2295
0 52 5 2 1 2345
0 53 7 2 2 2221 2304
0 54 5 1 1 2349
0 55 7 2 2 2239 2287
0 56 5 1 1 2351
0 57 7 1 2 2350 2352
0 58 5 2 1 57
0 59 7 1 2 54 56
0 60 5 1 1 59
0 61 7 2 2 2353 60
0 62 5 1 1 2355
0 63 7 1 2 2346 2356
0 64 5 2 1 63
0 65 7 2 2 2354 2357
0 66 5 1 1 2359
0 67 7 2 2 2231 2305
0 68 5 1 1 2361
0 69 7 2 2 2240 2296
0 70 5 1 1 2363
0 71 7 1 2 68 2364
0 72 5 1 1 71
0 73 7 1 2 2362 70
0 74 5 1 1 73
0 75 7 2 2 72 74
0 76 5 1 1 2365
0 77 7 1 2 66 76
0 78 5 3 1 77
0 79 7 1 2 2347 2367
0 80 5 1 1 79
0 81 7 2 2 2344 80
0 82 5 2 1 2370
0 83 7 2 2 2213 2306
0 84 5 1 1 2374
0 85 7 2 2 2241 2279
0 86 5 1 1 2376
0 87 7 1 2 2375 2377
0 88 5 2 1 87
0 89 7 2 2 2232 2288
0 90 5 1 1 2380
0 91 7 1 2 84 86
0 92 5 1 1 91
0 93 7 2 2 2378 92
0 94 5 1 1 2382
0 95 7 1 2 2381 2383
0 96 5 2 1 95
0 97 7 2 2 2379 2384
0 98 5 1 1 2386
0 99 7 1 2 2348 62
0 100 5 1 1 99
0 101 7 2 2 2358 100
0 102 5 1 1 2388
0 103 7 1 2 98 2389
0 104 5 2 1 103
0 105 7 2 2 2222 2297
0 106 5 1 1 2392
0 107 7 1 2 90 94
0 108 5 1 1 107
0 109 7 2 2 2385 108
0 110 5 1 1 2394
0 111 7 1 2 2393 2395
0 112 5 2 1 111
0 113 7 2 2 2204 2307
0 114 5 1 1 2398
0 115 7 2 2 2242 2271
0 116 5 1 1 2400
0 117 7 1 2 2399 2401
0 118 5 2 1 117
0 119 7 2 2 2233 2280
0 120 5 1 1 2404
0 121 7 1 2 114 116
0 122 5 1 1 121
0 123 7 2 2 2402 122
0 124 5 1 1 2406
0 125 7 1 2 2405 2407
0 126 5 2 1 125
0 127 7 2 2 2403 2408
0 128 5 1 1 2410
0 129 7 1 2 106 110
0 130 5 1 1 129
0 131 7 2 2 2396 130
0 132 5 1 1 2412
0 133 7 1 2 128 2413
0 134 5 2 1 133
0 135 7 2 2 2397 2414
0 136 5 1 1 2416
0 137 7 1 2 2387 102
0 138 5 1 1 137
0 139 7 2 2 2390 138
0 140 5 1 1 2418
0 141 7 1 2 136 2419
0 142 5 2 1 141
0 143 7 2 2 2391 2420
0 144 5 1 1 2422
0 145 7 1 2 2360 2366
0 146 5 1 1 145
0 147 7 2 2 2368 146
0 148 5 1 1 2424
0 149 7 1 2 144 2425
0 150 5 2 1 149
0 151 7 2 2 2214 2298
0 152 5 1 1 2428
0 153 7 1 2 120 124
0 154 5 1 1 153
0 155 7 2 2 2409 154
0 156 5 1 1 2430
0 157 7 1 2 2429 2431
0 158 5 2 1 157
0 159 7 2 2 2223 2289
0 160 5 1 1 2434
0 161 7 1 2 152 156
0 162 5 1 1 161
0 163 7 2 2 2432 162
0 164 5 1 1 2436
0 165 7 1 2 2435 2437
0 166 5 2 1 165
0 167 7 2 2 2433 2438
0 168 5 1 1 2440
0 169 7 1 2 2411 132
0 170 5 1 1 169
0 171 7 2 2 2415 170
0 172 5 1 1 2442
0 173 7 1 2 168 2443
0 174 5 2 1 173
0 175 7 2 2 2196 2308
0 176 5 1 1 2446
0 177 7 2 2 2243 2246
0 178 5 1 1 2448
0 179 7 2 2 2234 2254
0 180 5 1 1 2450
0 181 7 2 2 2449 2451
0 182 5 2 1 2452
0 183 7 2 2 2262 2453
0 184 5 2 1 2456
0 185 7 1 2 2447 2457
0 186 5 2 1 185
0 187 7 2 2 2244 2263
0 188 5 1 1 2462
0 189 7 1 2 176 2458
0 190 5 1 1 189
0 191 7 2 2 2460 190
0 192 5 1 1 2464
0 193 7 1 2 2463 2465
0 194 5 2 1 193
0 195 7 2 2 2461 2466
0 196 5 1 1 2468
0 197 7 1 2 160 164
0 198 5 1 1 197
0 199 7 2 2 2439 198
0 200 5 1 1 2470
0 201 7 1 2 196 2471
0 202 5 2 1 201
0 203 7 2 2 2224 2281
0 204 5 1 1 2474
0 205 7 1 2 188 192
0 206 5 1 1 205
0 207 7 2 2 2467 206
0 208 5 1 1 2476
0 209 7 1 2 2475 2477
0 210 5 2 1 209
0 211 7 2 2 2235 2272
0 212 5 1 1 2480
0 213 7 1 2 204 208
0 214 5 1 1 213
0 215 7 2 2 2478 214
0 216 5 1 1 2482
0 217 7 1 2 2481 2483
0 218 5 2 1 217
0 219 7 2 2 2479 2484
0 220 5 1 1 2486
0 221 7 1 2 2469 200
0 222 5 1 1 221
0 223 7 2 2 2472 222
0 224 5 1 1 2488
0 225 7 1 2 220 2489
0 226 5 2 1 225
0 227 7 2 2 2473 2490
0 228 5 1 1 2492
0 229 7 1 2 2441 172
0 230 5 1 1 229
0 231 7 2 2 2444 230
0 232 5 1 1 2494
0 233 7 1 2 228 2495
0 234 5 2 1 233
0 235 7 2 2 2445 2496
0 236 5 1 1 2498
0 237 7 1 2 2417 140
0 238 5 1 1 237
0 239 7 2 2 2421 238
0 240 5 1 1 2500
0 241 7 1 2 236 2501
0 242 5 2 1 241
0 243 7 2 2 2205 2299
0 244 5 1 1 2504
0 245 7 2 2 2215 2290
0 246 5 1 1 2506
0 247 7 1 2 2505 2507
0 248 5 2 1 247
0 249 7 1 2 212 216
0 250 5 1 1 249
0 251 7 2 2 2485 250
0 252 5 1 1 2510
0 253 7 1 2 244 246
0 254 5 1 1 253
0 255 7 2 2 2508 254
0 256 5 1 1 2512
0 257 7 1 2 2511 2513
0 258 5 2 1 257
0 259 7 2 2 2509 2514
0 260 5 1 1 2516
0 261 7 1 2 2487 224
0 262 5 1 1 261
0 263 7 2 2 2491 262
0 264 5 1 1 2518
0 265 7 1 2 260 2519
0 266 5 2 1 265
0 267 7 2 2 2225 2273
0 268 5 1 1 2522
0 269 7 2 2 2197 2300
0 270 5 1 1 2524
0 271 7 1 2 2523 2525
0 272 5 2 1 271
0 273 7 2 2 2188 2309
0 274 5 1 1 2528
0 275 7 2 2 2216 2282
0 276 5 1 1 2530
0 277 7 1 2 2236 2264
0 278 5 1 1 277
0 279 7 1 2 2454 278
0 280 5 1 1 279
0 281 7 2 2 2459 280
0 282 5 1 1 2532
0 283 7 1 2 2531 2533
0 284 5 2 1 283
0 285 7 1 2 276 282
0 286 5 1 1 285
0 287 7 2 2 2534 286
0 288 5 1 1 2536
0 289 7 1 2 2529 2537
0 290 5 2 1 289
0 291 7 1 2 274 288
0 292 5 1 1 291
0 293 7 2 2 2538 292
0 294 5 1 1 2540
0 295 7 1 2 268 270
0 296 5 1 1 295
0 297 7 2 2 2526 296
0 298 5 1 1 2542
0 299 7 1 2 2541 2543
0 300 5 2 1 299
0 301 7 2 2 2527 2544
0 302 5 1 1 2546
0 303 7 1 2 252 256
0 304 5 1 1 303
0 305 7 2 2 2515 304
0 306 5 1 1 2548
0 307 7 1 2 302 2549
0 308 5 2 1 307
0 309 7 2 2 2245 2255
0 310 5 1 1 2552
0 311 7 2 2 2206 2291
0 312 5 1 1 2554
0 313 7 1 2 2553 2555
0 314 5 2 1 313
0 315 7 1 2 294 298
0 316 5 1 1 315
0 317 7 2 2 2545 316
0 318 5 1 1 2558
0 319 7 1 2 310 312
0 320 5 1 1 319
0 321 7 2 2 2556 320
0 322 5 1 1 2560
0 323 7 1 2 2559 2561
0 324 5 2 1 323
0 325 7 2 2 2557 2562
0 326 5 1 1 2564
0 327 7 1 2 2547 306
0 328 5 1 1 327
0 329 7 2 2 2550 328
0 330 5 1 1 2566
0 331 7 1 2 326 2567
0 332 5 2 1 331
0 333 7 2 2 2551 2568
0 334 5 1 1 2570
0 335 7 1 2 2517 264
0 336 5 1 1 335
0 337 7 2 2 2520 336
0 338 5 1 1 2572
0 339 7 1 2 334 2573
0 340 5 2 1 339
0 341 7 2 2 2521 2574
0 342 5 1 1 2576
0 343 7 1 2 2493 232
0 344 5 1 1 343
0 345 7 2 2 2497 344
0 346 5 1 1 2578
0 347 7 1 2 342 2579
0 348 5 2 1 347
0 349 7 2 2 2535 2539
0 350 5 1 1 2582
0 351 7 1 2 2565 330
0 352 5 1 1 351
0 353 7 2 2 2569 352
0 354 5 1 1 2584
0 355 7 1 2 350 2585
0 356 5 2 1 355
0 357 7 2 2 2226 2265
0 358 5 1 1 2588
0 359 7 2 2 2217 2274
0 360 5 1 1 2590
0 361 7 1 2 2589 2591
0 362 5 2 1 361
0 363 7 2 2 2189 2301
0 364 5 1 1 2594
0 365 7 1 2 358 360
0 366 5 1 1 365
0 367 7 2 2 2592 366
0 368 5 1 1 2596
0 369 7 1 2 2595 2597
0 370 5 2 1 369
0 371 7 2 2 2593 2598
0 372 5 1 1 2600
0 373 7 2 2 2198 2292
0 374 5 1 1 2602
0 375 7 2 2 32 2310
0 376 5 1 1 2604
0 377 7 1 2 2603 2605
0 378 5 2 1 377
0 379 7 2 2 2207 2283
0 380 5 1 1 2608
0 381 7 2 2 2218 2256
0 382 5 1 1 2610
0 383 7 2 2 2181 2275
0 384 5 1 1 2612
0 385 7 2 2 2199 2257
0 386 5 1 1 2614
0 387 7 2 2 2613 2615
0 388 5 2 1 2616
0 389 7 2 2 2208 2617
0 390 5 2 1 2620
0 391 7 2 2 2611 2621
0 392 5 2 1 2624
0 393 7 2 2 2227 2625
0 394 5 2 1 2628
0 395 7 1 2 2609 2629
0 396 5 2 1 395
0 397 7 1 2 380 2630
0 398 5 1 1 397
0 399 7 2 2 2632 398
0 400 5 1 1 2634
0 401 7 1 2 178 180
0 402 5 1 1 401
0 403 7 2 2 2455 402
0 404 5 1 1 2636
0 405 7 1 2 2635 2637
0 406 5 2 1 405
0 407 7 1 2 400 404
0 408 5 1 1 407
0 409 7 2 2 2638 408
0 410 5 1 1 2640
0 411 7 1 2 374 376
0 412 5 1 1 411
0 413 7 2 2 2606 412
0 414 5 1 1 2642
0 415 7 1 2 2641 2643
0 416 5 2 1 415
0 417 7 2 2 2607 2644
0 418 5 1 1 2646
0 419 7 1 2 372 418
0 420 5 2 1 419
0 421 7 2 2 2633 2639
0 422 5 1 1 2650
0 423 7 1 2 2601 2647
0 424 5 1 1 423
0 425 7 2 2 2648 424
0 426 5 1 1 2652
0 427 7 1 2 422 2653
0 428 5 2 1 427
0 429 7 2 2 2649 2654
0 430 5 1 1 2656
0 431 7 1 2 2583 354
0 432 5 1 1 431
0 433 7 2 2 2586 432
0 434 5 1 1 2658
0 435 7 1 2 430 2659
0 436 5 2 1 435
0 437 7 2 2 2587 2660
0 438 5 1 1 2662
0 439 7 1 2 2571 338
0 440 5 1 1 439
0 441 7 2 2 2575 440
0 442 5 1 1 2664
0 443 7 1 2 438 2665
0 444 5 2 1 443
0 445 7 1 2 318 322
0 446 5 1 1 445
0 447 7 2 2 2563 446
0 448 5 1 1 2668
0 449 7 1 2 2651 426
0 450 5 1 1 449
0 451 7 2 2 2655 450
0 452 5 1 1 2670
0 453 7 1 2 2669 2671
0 454 5 2 1 453
0 455 7 1 2 364 368
0 456 5 1 1 455
0 457 7 2 2 2599 456
0 458 5 1 1 2674
0 459 7 1 2 410 414
0 460 5 1 1 459
0 461 7 2 2 2645 460
0 462 5 1 1 2676
0 463 7 1 2 2675 2677
0 464 5 2 1 463
0 465 7 2 2 2209 2276
0 466 5 1 1 2680
0 467 7 2 2 2200 2284
0 468 5 1 1 2682
0 469 7 1 2 2681 2683
0 470 5 2 1 469
0 471 7 2 2 2190 2293
0 472 5 1 1 2686
0 473 7 1 2 466 468
0 474 5 1 1 473
0 475 7 2 2 2684 474
0 476 5 1 1 2688
0 477 7 1 2 2687 2689
0 478 5 2 1 477
0 479 7 2 2 2685 2690
0 480 5 1 1 2692
0 481 7 1 2 458 462
0 482 5 1 1 481
0 483 7 2 2 2678 482
0 484 5 1 1 2694
0 485 7 1 2 480 2695
0 486 5 2 1 485
0 487 7 2 2 2679 2696
0 488 5 1 1 2698
0 489 7 1 2 448 452
0 490 5 1 1 489
0 491 7 2 2 2672 490
0 492 5 1 1 2700
0 493 7 1 2 488 2701
0 494 5 2 1 493
0 495 7 2 2 2673 2702
0 496 5 1 1 2704
0 497 7 1 2 2657 434
0 498 5 1 1 497
0 499 7 2 2 2661 498
0 500 5 1 1 2706
0 501 7 1 2 496 2707
0 502 5 2 1 501
0 503 7 2 2 2182 2302
0 504 5 1 1 2710
0 505 7 1 2 472 476
0 506 5 1 1 505
0 507 7 2 2 2691 506
0 508 5 1 1 2712
0 509 7 1 2 2711 2713
0 510 5 2 1 509
0 511 7 2 2 2237 2247
0 512 5 1 1 2716
0 513 7 2 2 2219 2266
0 514 5 1 1 2718
0 515 7 1 2 2228 2258
0 516 5 1 1 515
0 517 7 1 2 2626 516
0 518 5 1 1 517
0 519 7 2 2 2631 518
0 520 5 1 1 2720
0 521 7 1 2 2719 2721
0 522 5 2 1 521
0 523 7 1 2 514 520
0 524 5 1 1 523
0 525 7 2 2 2722 524
0 526 5 1 1 2724
0 527 7 1 2 2717 2725
0 528 5 2 1 527
0 529 7 1 2 512 526
0 530 5 1 1 529
0 531 7 2 2 2726 530
0 532 5 1 1 2728
0 533 7 1 2 504 508
0 534 5 1 1 533
0 535 7 2 2 2714 534
0 536 5 1 1 2730
0 537 7 1 2 2729 2731
0 538 5 2 1 537
0 539 7 2 2 2715 2732
0 540 5 1 1 2734
0 541 7 1 2 2693 484
0 542 5 1 1 541
0 543 7 2 2 2697 542
0 544 5 1 1 2736
0 545 7 1 2 540 2737
0 546 5 2 1 545
0 547 7 2 2 2723 2727
0 548 5 1 1 2740
0 549 7 1 2 2735 544
0 550 5 1 1 549
0 551 7 2 2 2738 550
0 552 5 1 1 2742
0 553 7 1 2 548 2743
0 554 5 2 1 553
0 555 7 2 2 2739 2744
0 556 5 1 1 2746
0 557 7 1 2 2699 492
0 558 5 1 1 557
0 559 7 2 2 2703 558
0 560 5 1 1 2748
0 561 7 1 2 556 2749
0 562 5 2 1 561
0 563 7 2 2 2210 2267
0 564 5 1 1 2752
0 565 7 1 2 382 2622
0 566 5 1 1 565
0 567 7 2 2 2627 566
0 568 5 1 1 2754
0 569 7 1 2 2753 2755
0 570 5 2 1 569
0 571 7 2 2 2229 2248
0 572 5 1 1 2758
0 573 7 1 2 564 568
0 574 5 1 1 573
0 575 7 2 2 2756 574
0 576 5 1 1 2760
0 577 7 1 2 2759 2761
0 578 5 2 1 577
0 579 7 2 2 2757 2762
0 580 5 1 1 2764
0 581 7 1 2 532 536
0 582 5 1 1 581
0 583 7 2 2 2733 582
0 584 5 1 1 2766
0 585 7 1 2 580 2767
0 586 5 2 1 585
0 587 7 2 2 2201 2277
0 588 5 1 1 2770
0 589 7 2 2 2183 2294
0 590 5 1 1 2772
0 591 7 1 2 2771 2773
0 592 5 2 1 591
0 593 7 1 2 572 576
0 594 5 1 1 593
0 595 7 2 2 2763 594
0 596 5 1 1 2776
0 597 7 1 2 588 590
0 598 5 1 1 597
0 599 7 2 2 2774 598
0 600 5 1 1 2778
0 601 7 1 2 2777 2779
0 602 5 2 1 601
0 603 7 2 2 2775 2780
0 604 5 1 1 2782
0 605 7 1 2 2765 584
0 606 5 1 1 605
0 607 7 2 2 2768 606
0 608 5 1 1 2784
0 609 7 1 2 604 2785
0 610 5 2 1 609
0 611 7 2 2 2769 2786
0 612 5 1 1 2788
0 613 7 1 2 2741 552
0 614 5 1 1 613
0 615 7 2 2 2745 614
0 616 5 1 1 2790
0 617 7 1 2 612 2791
0 618 5 2 1 617
0 619 7 2 2 2191 2285
0 620 5 1 1 2794
0 621 7 1 2 596 600
0 622 5 1 1 621
0 623 7 2 2 2781 622
0 624 5 1 1 2796
0 625 7 1 2 2795 2797
0 626 5 2 1 625
0 627 7 2 2 2202 2268
0 628 5 1 1 2800
0 629 7 1 2 2211 2259
0 630 5 1 1 629
0 631 7 1 2 2618 630
0 632 5 1 1 631
0 633 7 2 2 2623 632
0 634 5 1 1 2802
0 635 7 1 2 2801 2803
0 636 5 2 1 635
0 637 7 2 2 2220 2249
0 638 5 1 1 2806
0 639 7 1 2 628 634
0 640 5 1 1 639
0 641 7 2 2 2804 640
0 642 5 1 1 2808
0 643 7 1 2 2807 2809
0 644 5 2 1 643
0 645 7 2 2 2805 2810
0 646 5 1 1 2812
0 647 7 1 2 620 624
0 648 5 1 1 647
0 649 7 2 2 2798 648
0 650 5 1 1 2814
0 651 7 1 2 646 2815
0 652 5 2 1 651
0 653 7 2 2 2799 2816
0 654 5 1 1 2818
0 655 7 1 2 2783 608
0 656 5 1 1 655
0 657 7 2 2 2787 656
0 658 5 1 1 2820
0 659 7 1 2 654 2821
0 660 5 2 1 659
0 661 7 2 2 2184 2286
0 662 5 1 1 2824
0 663 7 2 2 2192 2278
0 664 5 1 1 2826
0 665 7 1 2 2825 2827
0 666 5 2 1 665
0 667 7 1 2 638 642
0 668 5 1 1 667
0 669 7 2 2 2811 668
0 670 5 1 1 2830
0 671 7 1 2 662 664
0 672 5 1 1 671
0 673 7 2 2 2828 672
0 674 5 1 1 2832
0 675 7 1 2 2831 2833
0 676 5 2 1 675
0 677 7 2 2 2829 2834
0 678 5 1 1 2836
0 679 7 1 2 2813 650
0 680 5 1 1 679
0 681 7 2 2 2817 680
0 682 5 1 1 2838
0 683 7 1 2 678 2839
0 684 5 2 1 683
0 685 7 1 2 670 674
0 686 5 1 1 685
0 687 7 2 2 2835 686
0 688 5 1 1 2842
0 689 7 2 2 2193 2269
0 690 5 1 1 2844
0 691 7 2 2 2212 2250
0 692 5 1 1 2846
0 693 7 2 2 2845 2847
0 694 5 1 1 2848
0 695 7 2 2 2194 2260
0 696 5 1 1 2850
0 697 7 2 2 2185 2270
0 698 5 1 1 2852
0 699 7 2 2 2851 2853
0 700 5 2 1 2854
0 701 7 3 2 694 2856
0 702 5 1 1 2858
0 703 7 1 2 2843 702
0 704 5 2 1 703
0 705 7 1 2 384 386
0 706 5 1 1 705
0 707 7 2 2 2619 706
0 708 5 1 1 2863
0 709 7 1 2 690 692
0 710 5 1 1 709
0 711 7 1 2 2859 710
0 712 5 1 1 711
0 713 7 1 2 2849 2855
0 714 5 1 1 713
0 715 7 2 2 712 714
0 716 5 1 1 2865
0 717 7 1 2 2864 716
0 718 5 2 1 717
0 719 7 2 2 2203 2251
0 720 5 1 1 2869
0 721 7 1 2 696 698
0 722 5 1 1 721
0 723 7 2 2 2857 722
0 724 5 1 1 2871
0 725 7 1 2 2870 2872
0 726 5 2 1 725
0 727 7 1 2 720 724
0 728 5 1 1 727
0 729 7 3 2 2873 728
0 730 5 2 1 2875
0 731 7 2 2 2186 2261
0 732 5 1 1 2880
0 733 7 2 2 2195 2252
0 734 5 1 1 2882
0 735 7 2 2 2881 2883
0 736 5 2 1 2884
0 737 7 1 2 2876 2885
0 738 5 2 1 737
0 739 7 2 2 2874 2888
0 740 5 1 1 2890
0 741 7 1 2 708 2866
0 742 5 1 1 741
0 743 7 2 2 2867 742
0 744 5 1 1 2892
0 745 7 1 2 740 2893
0 746 5 2 1 745
0 747 7 2 2 2868 2894
0 748 5 1 1 2896
0 749 7 1 2 688 2860
0 750 5 1 1 749
0 751 7 2 2 2861 750
0 752 5 1 1 2898
0 753 7 1 2 748 2899
0 754 5 2 1 753
0 755 7 2 2 2862 2900
0 756 5 1 1 2902
0 757 7 1 2 2837 682
0 758 5 1 1 757
0 759 7 2 2 2840 758
0 760 5 1 1 2904
0 761 7 1 2 756 2905
0 762 5 2 1 761
0 763 7 2 2 2841 2906
0 764 5 1 1 2908
0 765 7 1 2 2819 658
0 766 5 1 1 765
0 767 7 2 2 2822 766
0 768 5 1 1 2910
0 769 7 1 2 764 2911
0 770 5 2 1 769
0 771 7 2 2 2823 2912
0 772 5 1 1 2914
0 773 7 1 2 2789 616
0 774 5 1 1 773
0 775 7 2 2 2792 774
0 776 5 1 1 2916
0 777 7 1 2 772 2917
0 778 5 2 1 777
0 779 7 2 2 2793 2918
0 780 5 1 1 2920
0 781 7 1 2 2747 560
0 782 5 1 1 781
0 783 7 2 2 2750 782
0 784 5 1 1 2922
0 785 7 1 2 780 2923
0 786 5 2 1 785
0 787 7 2 2 2751 2924
0 788 5 1 1 2926
0 789 7 1 2 2705 500
0 790 5 1 1 789
0 791 7 2 2 2708 790
0 792 5 1 1 2928
0 793 7 1 2 788 2929
0 794 5 2 1 793
0 795 7 2 2 2709 2930
0 796 5 1 1 2932
0 797 7 1 2 2663 442
0 798 5 1 1 797
0 799 7 2 2 2666 798
0 800 5 1 1 2934
0 801 7 1 2 796 2935
0 802 5 2 1 801
0 803 7 2 2 2667 2936
0 804 5 1 1 2938
0 805 7 1 2 2577 346
0 806 5 1 1 805
0 807 7 2 2 2580 806
0 808 5 1 1 2940
0 809 7 1 2 804 2941
0 810 5 2 1 809
0 811 7 2 2 2581 2942
0 812 5 1 1 2944
0 813 7 1 2 2499 240
0 814 5 1 1 813
0 815 7 2 2 2502 814
0 816 5 1 1 2946
0 817 7 1 2 812 2947
0 818 5 2 1 817
0 819 7 2 2 2503 2948
0 820 5 1 1 2950
0 821 7 1 2 2423 148
0 822 5 1 1 821
0 823 7 2 2 2426 822
0 824 5 1 1 2952
0 825 7 1 2 820 2953
0 826 5 2 1 825
0 827 7 3 2 2427 2954
0 828 5 2 1 2956
0 829 7 2 2 50 2369
0 830 5 1 1 2961
0 831 7 2 2 2372 830
0 832 5 1 1 2963
0 833 7 1 2 2959 2964
0 834 5 2 1 833
0 835 7 3 2 2373 2965
0 836 5 2 1 2967
0 837 7 1 2 48 2970
0 838 5 5 1 837
0 839 7 1 2 2342 2968
0 840 5 5 1 839
0 841 7 1 2 2957 832
0 842 5 1 1 841
0 843 7 3 2 2966 842
0 844 5 2 1 2982
0 845 7 1 2 2340 2985
0 846 5 3 1 845
0 847 7 1 2 2951 824
0 848 5 1 1 847
0 849 7 4 2 2955 848
0 850 5 3 1 2990
0 851 7 1 2 2338 2994
0 852 5 3 1 851
0 853 7 1 2 2945 816
0 854 5 1 1 853
0 855 7 4 2 2949 854
0 856 5 3 1 3000
0 857 7 1 2 2336 3004
0 858 5 3 1 857
0 859 7 1 2 2939 808
0 860 5 1 1 859
0 861 7 4 2 2943 860
0 862 5 3 1 3010
0 863 7 1 2 2334 3014
0 864 5 3 1 863
0 865 7 1 2 2933 800
0 866 5 1 1 865
0 867 7 4 2 2937 866
0 868 5 3 1 3020
0 869 7 1 2 2332 3024
0 870 5 3 1 869
0 871 7 1 2 2927 792
0 872 5 1 1 871
0 873 7 4 2 2931 872
0 874 5 3 1 3030
0 875 7 1 2 2330 3034
0 876 5 3 1 875
0 877 7 1 2 2921 784
0 878 5 1 1 877
0 879 7 4 2 2925 878
0 880 5 3 1 3040
0 881 7 1 2 2328 3044
0 882 5 3 1 881
0 883 7 1 2 41 3041
0 884 5 3 1 883
0 885 7 1 2 2915 776
0 886 5 1 1 885
0 887 7 4 2 2919 886
0 888 5 3 1 3053
0 889 7 1 2 2326 3057
0 890 5 3 1 889
0 891 7 1 2 2909 768
0 892 5 1 1 891
0 893 7 4 2 2913 892
0 894 5 3 1 3063
0 895 7 1 2 2324 3067
0 896 5 3 1 895
0 897 7 1 2 39 3064
0 898 5 3 1 897
0 899 7 1 2 2903 760
0 900 5 1 1 899
0 901 7 4 2 2907 900
0 902 5 3 1 3076
0 903 7 1 2 2322 3080
0 904 5 3 1 903
0 905 7 1 2 2897 752
0 906 5 1 1 905
0 907 7 4 2 2901 906
0 908 5 3 1 3086
0 909 7 1 2 2320 3090
0 910 5 3 1 909
0 911 7 1 2 2891 744
0 912 5 1 1 911
0 913 7 4 2 2895 912
0 914 5 3 1 3096
0 915 7 1 2 2318 3100
0 916 5 3 1 915
0 917 7 1 2 2878 2886
0 918 5 1 1 917
0 919 7 3 2 2889 918
0 920 5 3 1 3106
0 921 7 1 2 2316 3109
0 922 5 3 1 921
0 923 7 1 2 35 3107
0 924 5 3 1 923
0 925 7 2 2 732 734
0 926 5 1 1 3118
0 927 7 4 2 2887 926
0 928 5 2 1 3120
0 929 7 1 2 2314 3124
0 930 5 3 1 929
0 931 7 1 2 34 3121
0 932 5 3 1 931
0 933 7 3 2 2187 2253
0 934 5 3 1 3132
0 935 7 2 2 33 3133
0 936 5 3 1 3138
0 937 7 1 2 3129 3140
0 938 5 1 1 937
0 939 7 2 2 3126 938
0 940 5 2 1 3143
0 941 7 1 2 3115 3145
0 942 5 1 1 941
0 943 7 2 2 3112 942
0 944 5 2 1 3147
0 945 7 1 2 36 3097
0 946 5 3 1 945
0 947 7 1 2 3149 3151
0 948 5 1 1 947
0 949 7 2 2 3103 948
0 950 5 2 1 3154
0 951 7 1 2 37 3087
0 952 5 3 1 951
0 953 7 1 2 3156 3158
0 954 5 1 1 953
0 955 7 2 2 3093 954
0 956 5 2 1 3161
0 957 7 1 2 38 3077
0 958 5 3 1 957
0 959 7 1 2 3163 3165
0 960 5 1 1 959
0 961 7 2 2 3083 960
0 962 5 2 1 3168
0 963 7 1 2 3073 3170
0 964 5 1 1 963
0 965 7 2 2 3070 964
0 966 5 2 1 3172
0 967 7 1 2 40 3054
0 968 5 3 1 967
0 969 7 1 2 3174 3176
0 970 5 1 1 969
0 971 7 2 2 3060 970
0 972 5 2 1 3179
0 973 7 1 2 3050 3181
0 974 5 1 1 973
0 975 7 2 2 3047 974
0 976 5 2 1 3183
0 977 7 1 2 42 3031
0 978 5 3 1 977
0 979 7 1 2 3185 3187
0 980 5 1 1 979
0 981 7 2 2 3037 980
0 982 5 2 1 3190
0 983 7 1 2 43 3021
0 984 5 3 1 983
0 985 7 1 2 3192 3194
0 986 5 1 1 985
0 987 7 2 2 3027 986
0 988 5 2 1 3197
0 989 7 1 2 44 3011
0 990 5 3 1 989
0 991 7 1 2 3199 3201
0 992 5 1 1 991
0 993 7 2 2 3017 992
0 994 5 2 1 3204
0 995 7 1 2 45 3001
0 996 5 3 1 995
0 997 7 1 2 3206 3208
0 998 5 1 1 997
0 999 7 2 2 3007 998
0 1000 5 2 1 3211
0 1001 7 1 2 46 2991
0 1002 5 3 1 1001
0 1003 7 1 2 3213 3215
0 1004 5 1 1 1003
0 1005 7 2 2 2997 1004
0 1006 5 2 1 3218
0 1007 7 1 2 47 2983
0 1008 5 3 1 1007
0 1009 7 1 2 3220 3222
0 1010 5 1 1 1009
0 1011 7 4 2 2987 1010
0 1012 5 2 1 3225
0 1013 7 1 2 2977 3226
0 1014 5 1 1 1013
0 1015 7 3 2 2972 1014
0 1016 5 1 1 3231
0 1017 7 3 2 2988 3223
0 1018 5 2 1 3234
0 1019 7 1 2 3219 3237
0 1020 5 1 1 1019
0 1021 7 1 2 3221 3235
0 1022 5 1 1 1021
0 1023 7 3 2 1020 1022
0 1024 5 2 1 3239
0 1025 7 1 2 1016 3240
0 1026 5 2 1 1025
0 1027 7 3 2 2998 3216
0 1028 5 2 1 3246
0 1029 7 1 2 3212 3249
0 1030 5 1 1 1029
0 1031 7 1 2 3214 3247
0 1032 5 1 1 1031
0 1033 7 3 2 1030 1032
0 1034 5 2 1 3251
0 1035 7 3 2 2973 2978
0 1036 5 2 1 3256
0 1037 7 1 2 3229 3257
0 1038 5 1 1 1037
0 1039 7 1 2 3227 3259
0 1040 5 1 1 1039
0 1041 7 2 2 1038 1040
0 1042 5 1 1 3261
0 1043 7 1 2 3252 3262
0 1044 5 2 1 1043
0 1045 7 3 2 3008 3209
0 1046 5 2 1 3265
0 1047 7 1 2 3205 3268
0 1048 5 1 1 1047
0 1049 7 1 2 3207 3266
0 1050 5 1 1 1049
0 1051 7 3 2 1048 1050
0 1052 5 2 1 3270
0 1053 7 1 2 3241 3271
0 1054 5 2 1 1053
0 1055 7 3 2 3018 3202
0 1056 5 2 1 3277
0 1057 7 1 2 3198 3280
0 1058 5 1 1 1057
0 1059 7 1 2 3200 3278
0 1060 5 1 1 1059
0 1061 7 3 2 1058 1060
0 1062 5 2 1 3282
0 1063 7 1 2 3253 3283
0 1064 5 2 1 1063
0 1065 7 3 2 3028 3195
0 1066 5 2 1 3289
0 1067 7 1 2 3191 3292
0 1068 5 1 1 1067
0 1069 7 1 2 3193 3290
0 1070 5 1 1 1069
0 1071 7 3 2 1068 1070
0 1072 5 2 1 3294
0 1073 7 1 2 3272 3295
0 1074 5 2 1 1073
0 1075 7 3 2 3038 3188
0 1076 5 2 1 3301
0 1077 7 1 2 3184 3304
0 1078 5 1 1 1077
0 1079 7 1 2 3186 3302
0 1080 5 1 1 1079
0 1081 7 3 2 1078 1080
0 1082 5 2 1 3306
0 1083 7 1 2 3284 3307
0 1084 5 2 1 1083
0 1085 7 3 2 3048 3051
0 1086 5 2 1 3313
0 1087 7 1 2 3182 3314
0 1088 5 1 1 1087
0 1089 7 1 2 3180 3316
0 1090 5 1 1 1089
0 1091 7 3 2 1088 1090
0 1092 5 2 1 3318
0 1093 7 1 2 3296 3319
0 1094 5 2 1 1093
0 1095 7 3 2 3061 3177
0 1096 5 2 1 3325
0 1097 7 1 2 3173 3328
0 1098 5 1 1 1097
0 1099 7 1 2 3175 3326
0 1100 5 1 1 1099
0 1101 7 3 2 1098 1100
0 1102 5 2 1 3330
0 1103 7 1 2 3308 3331
0 1104 5 2 1 1103
0 1105 7 3 2 3071 3074
0 1106 5 2 1 3337
0 1107 7 1 2 3171 3338
0 1108 5 1 1 1107
0 1109 7 1 2 3169 3340
0 1110 5 1 1 1109
0 1111 7 3 2 1108 1110
0 1112 5 2 1 3342
0 1113 7 1 2 3320 3343
0 1114 5 2 1 1113
0 1115 7 3 2 3084 3166
0 1116 5 2 1 3349
0 1117 7 1 2 3162 3352
0 1118 5 1 1 1117
0 1119 7 1 2 3164 3350
0 1120 5 1 1 1119
0 1121 7 3 2 1118 1120
0 1122 5 2 1 3354
0 1123 7 1 2 3332 3355
0 1124 5 2 1 1123
0 1125 7 3 2 3094 3159
0 1126 5 2 1 3361
0 1127 7 1 2 3155 3364
0 1128 5 1 1 1127
0 1129 7 1 2 3157 3362
0 1130 5 1 1 1129
0 1131 7 3 2 1128 1130
0 1132 5 2 1 3366
0 1133 7 1 2 3344 3367
0 1134 5 2 1 1133
0 1135 7 3 2 3104 3152
0 1136 5 2 1 3373
0 1137 7 1 2 3148 3376
0 1138 5 1 1 1137
0 1139 7 1 2 3150 3374
0 1140 5 1 1 1139
0 1141 7 3 2 1138 1140
0 1142 5 2 1 3378
0 1143 7 1 2 3356 3379
0 1144 5 2 1 1143
0 1145 7 3 2 3113 3116
0 1146 5 2 1 3385
0 1147 7 1 2 3146 3386
0 1148 5 1 1 1147
0 1149 7 1 2 3144 3388
0 1150 5 1 1 1149
0 1151 7 3 2 1148 1150
0 1152 5 2 1 3390
0 1153 7 1 2 3368 3391
0 1154 5 2 1 1153
0 1155 7 3 2 3127 3130
0 1156 5 2 1 3397
0 1157 7 1 2 3141 3398
0 1158 5 1 1 1157
0 1159 7 1 2 3139 3400
0 1160 5 1 1 1159
0 1161 7 2 2 1158 1160
0 1162 5 2 1 3402
0 1163 7 1 2 3380 3403
0 1164 5 2 1 1163
0 1165 7 3 2 2312 3135
0 1166 5 3 1 3408
0 1167 7 3 2 3142 3411
0 1168 5 2 1 3414
0 1169 7 2 2 3392 3417
0 1170 5 2 1 3419
0 1171 7 1 2 3381 3404
0 1172 5 1 1 1171
0 1173 7 2 2 3406 1172
0 1174 5 1 1 3423
0 1175 7 1 2 3420 3424
0 1176 5 2 1 1175
0 1177 7 2 2 3407 3425
0 1178 5 1 1 3427
0 1179 7 1 2 3369 3393
0 1180 5 1 1 1179
0 1181 7 2 2 3395 1180
0 1182 5 1 1 3429
0 1183 7 1 2 1178 3430
0 1184 5 2 1 1183
0 1185 7 2 2 3396 3431
0 1186 5 1 1 3433
0 1187 7 1 2 3357 3382
0 1188 5 1 1 1187
0 1189 7 2 2 3383 1188
0 1190 5 1 1 3435
0 1191 7 1 2 1186 3436
0 1192 5 2 1 1191
0 1193 7 2 2 3384 3437
0 1194 5 1 1 3439
0 1195 7 1 2 3345 3370
0 1196 5 1 1 1195
0 1197 7 2 2 3371 1196
0 1198 5 1 1 3441
0 1199 7 1 2 1194 3442
0 1200 5 2 1 1199
0 1201 7 2 2 3372 3443
0 1202 5 1 1 3445
0 1203 7 1 2 3333 3358
0 1204 5 1 1 1203
0 1205 7 2 2 3359 1204
0 1206 5 1 1 3447
0 1207 7 1 2 1202 3448
0 1208 5 2 1 1207
0 1209 7 2 2 3360 3449
0 1210 5 1 1 3451
0 1211 7 1 2 3321 3346
0 1212 5 1 1 1211
0 1213 7 2 2 3347 1212
0 1214 5 1 1 3453
0 1215 7 1 2 1210 3454
0 1216 5 2 1 1215
0 1217 7 2 2 3348 3455
0 1218 5 1 1 3457
0 1219 7 1 2 3309 3334
0 1220 5 1 1 1219
0 1221 7 2 2 3335 1220
0 1222 5 1 1 3459
0 1223 7 1 2 1218 3460
0 1224 5 2 1 1223
0 1225 7 2 2 3336 3461
0 1226 5 1 1 3463
0 1227 7 1 2 3297 3322
0 1228 5 1 1 1227
0 1229 7 2 2 3323 1228
0 1230 5 1 1 3465
0 1231 7 1 2 1226 3466
0 1232 5 2 1 1231
0 1233 7 2 2 3324 3467
0 1234 5 1 1 3469
0 1235 7 1 2 3285 3310
0 1236 5 1 1 1235
0 1237 7 2 2 3311 1236
0 1238 5 1 1 3471
0 1239 7 1 2 1234 3472
0 1240 5 2 1 1239
0 1241 7 2 2 3312 3473
0 1242 5 1 1 3475
0 1243 7 1 2 3273 3298
0 1244 5 1 1 1243
0 1245 7 2 2 3299 1244
0 1246 5 1 1 3477
0 1247 7 1 2 1242 3478
0 1248 5 2 1 1247
0 1249 7 2 2 3300 3479
0 1250 5 1 1 3481
0 1251 7 1 2 3254 3286
0 1252 5 1 1 1251
0 1253 7 2 2 3287 1252
0 1254 5 1 1 3483
0 1255 7 1 2 1250 3484
0 1256 5 2 1 1255
0 1257 7 2 2 3288 3485
0 1258 5 1 1 3487
0 1259 7 1 2 3242 3274
0 1260 5 1 1 1259
0 1261 7 2 2 3275 1260
0 1262 5 1 1 3489
0 1263 7 1 2 1258 3490
0 1264 5 2 1 1263
0 1265 7 2 2 3276 3491
0 1266 5 1 1 3493
0 1267 7 1 2 3255 1042
0 1268 5 1 1 1267
0 1269 7 2 2 3263 1268
0 1270 5 1 1 3495
0 1271 7 1 2 1266 3496
0 1272 5 2 1 1271
0 1273 7 2 2 3264 3497
0 1274 5 1 1 3499
0 1275 7 1 2 3232 3243
0 1276 5 1 1 1275
0 1277 7 2 2 3244 1276
0 1278 5 1 1 3501
0 1279 7 1 2 1274 3502
0 1280 5 2 1 1279
0 1281 7 2 2 3245 3503
0 1282 5 1 1 3505
0 1283 7 1 2 2974 3228
0 1284 5 1 1 1283
0 1285 7 1 2 2979 3230
0 1286 5 1 1 1285
0 1287 7 2 2 1284 1286
0 1288 5 1 1 3507
0 1289 7 1 2 1282 3508
0 1290 5 2 1 1289
0 1291 7 1 2 3506 1288
0 1292 5 2 1 1291
0 1293 7 1 2 3509 3511
0 1294 5 1 1 1293
0 1295 7 1 2 2371 2960
0 1296 5 2 1 1295
0 1297 7 1 2 2984 2992
0 1298 5 2 1 1297
0 1299 7 1 2 2993 3002
0 1300 5 2 1 1299
0 1301 7 1 2 3003 3012
0 1302 5 2 1 1301
0 1303 7 1 2 3013 3022
0 1304 5 2 1 1303
0 1305 7 1 2 3023 3032
0 1306 5 2 1 1305
0 1307 7 1 2 3033 3042
0 1308 5 2 1 1307
0 1309 7 1 2 3043 3055
0 1310 5 2 1 1309
0 1311 7 1 2 3056 3065
0 1312 5 2 1 1311
0 1313 7 1 2 3066 3078
0 1314 5 2 1 1313
0 1315 7 1 2 3079 3088
0 1316 5 2 1 1315
0 1317 7 1 2 3089 3098
0 1318 5 2 1 1317
0 1319 7 1 2 3099 3108
0 1320 5 2 1 1319
0 1321 7 1 2 3101 3110
0 1322 5 1 1 1321
0 1323 7 2 2 3537 1322
0 1324 5 1 1 3539
0 1325 7 1 2 2879 3136
0 1326 5 1 1 1325
0 1327 7 2 2 3122 1326
0 1328 5 2 1 3541
0 1329 7 1 2 3540 3542
0 1330 5 2 1 1329
0 1331 7 2 2 3538 3545
0 1332 5 1 1 3547
0 1333 7 1 2 3091 3102
0 1334 5 1 1 1333
0 1335 7 2 2 3535 1334
0 1336 5 1 1 3549
0 1337 7 1 2 1332 3550
0 1338 5 2 1 1337
0 1339 7 2 2 3536 3551
0 1340 5 1 1 3553
0 1341 7 1 2 3081 3092
0 1342 5 1 1 1341
0 1343 7 2 2 3533 1342
0 1344 5 1 1 3555
0 1345 7 1 2 1340 3556
0 1346 5 2 1 1345
0 1347 7 2 2 3534 3557
0 1348 5 1 1 3559
0 1349 7 1 2 3068 3082
0 1350 5 1 1 1349
0 1351 7 2 2 3531 1350
0 1352 5 1 1 3561
0 1353 7 1 2 1348 3562
0 1354 5 2 1 1353
0 1355 7 2 2 3532 3563
0 1356 5 1 1 3565
0 1357 7 1 2 3058 3069
0 1358 5 1 1 1357
0 1359 7 2 2 3529 1358
0 1360 5 1 1 3567
0 1361 7 1 2 1356 3568
0 1362 5 2 1 1361
0 1363 7 2 2 3530 3569
0 1364 5 1 1 3571
0 1365 7 1 2 3045 3059
0 1366 5 1 1 1365
0 1367 7 2 2 3527 1366
0 1368 5 1 1 3573
0 1369 7 1 2 1364 3574
0 1370 5 2 1 1369
0 1371 7 2 2 3528 3575
0 1372 5 1 1 3577
0 1373 7 1 2 3035 3046
0 1374 5 1 1 1373
0 1375 7 2 2 3525 1374
0 1376 5 1 1 3579
0 1377 7 1 2 1372 3580
0 1378 5 2 1 1377
0 1379 7 2 2 3526 3581
0 1380 5 1 1 3583
0 1381 7 1 2 3025 3036
0 1382 5 1 1 1381
0 1383 7 2 2 3523 1382
0 1384 5 1 1 3585
0 1385 7 1 2 1380 3586
0 1386 5 2 1 1385
0 1387 7 2 2 3524 3587
0 1388 5 1 1 3589
0 1389 7 1 2 3015 3026
0 1390 5 1 1 1389
0 1391 7 2 2 3521 1390
0 1392 5 1 1 3591
0 1393 7 1 2 1388 3592
0 1394 5 2 1 1393
0 1395 7 2 2 3522 3593
0 1396 5 1 1 3595
0 1397 7 1 2 3005 3016
0 1398 5 1 1 1397
0 1399 7 2 2 3519 1398
0 1400 5 1 1 3597
0 1401 7 1 2 1396 3598
0 1402 5 2 1 1401
0 1403 7 2 2 3520 3599
0 1404 5 1 1 3601
0 1405 7 1 2 2995 3006
0 1406 5 1 1 1405
0 1407 7 2 2 3517 1406
0 1408 5 1 1 3603
0 1409 7 1 2 1404 3604
0 1410 5 2 1 1409
0 1411 7 2 2 3518 3605
0 1412 5 1 1 3607
0 1413 7 1 2 2986 2996
0 1414 5 1 1 1413
0 1415 7 2 2 3515 1414
0 1416 5 1 1 3609
0 1417 7 1 2 1412 3610
0 1418 5 2 1 1417
0 1419 7 2 2 3516 3611
0 1420 5 1 1 3613
0 1421 7 1 2 2958 2962
0 1422 5 1 1 1421
0 1423 7 2 2 3513 1422
0 1424 5 1 1 3615
0 1425 7 2 2 1420 3616
0 1426 5 2 1 3617
0 1427 7 1 2 2971 3618
0 1428 5 1 1 1427
0 1429 7 5 2 3514 1428
0 1430 5 1 1 3621
0 1431 7 1 2 1294 1430
0 1432 5 1 1 1431
0 1433 7 1 2 3500 1278
0 1434 5 1 1 1433
0 1435 7 2 2 3504 1434
0 1436 5 1 1 3626
0 1437 7 1 2 2969 3619
0 1438 5 3 1 1437
0 1439 7 2 2 3622 3628
0 1440 5 1 1 3631
0 1441 7 1 2 3627 1440
0 1442 5 1 1 1441
0 1443 7 1 2 1436 3632
0 1444 5 1 1 1443
0 1445 7 1 2 3614 1424
0 1446 5 1 1 1445
0 1447 7 3 2 3620 1446
0 1448 5 2 1 3633
0 1449 7 1 2 3494 1270
0 1450 5 1 1 1449
0 1451 7 2 2 3498 1450
0 1452 5 1 1 3638
0 1453 7 1 2 3634 1452
0 1454 5 1 1 1453
0 1455 7 1 2 3636 3639
0 1456 5 1 1 1455
0 1457 7 1 2 3608 1416
0 1458 5 1 1 1457
0 1459 7 3 2 3612 1458
0 1460 5 2 1 3640
0 1461 7 1 2 3488 1262
0 1462 5 1 1 1461
0 1463 7 2 2 3492 1462
0 1464 5 1 1 3645
0 1465 7 1 2 3641 1464
0 1466 5 1 1 1465
0 1467 7 1 2 3643 3646
0 1468 5 1 1 1467
0 1469 7 1 2 3602 1408
0 1470 5 1 1 1469
0 1471 7 3 2 3606 1470
0 1472 5 2 1 3647
0 1473 7 1 2 3482 1254
0 1474 5 1 1 1473
0 1475 7 2 2 3486 1474
0 1476 5 1 1 3652
0 1477 7 1 2 3648 1476
0 1478 5 1 1 1477
0 1479 7 1 2 3650 3653
0 1480 5 1 1 1479
0 1481 7 1 2 3596 1400
0 1482 5 1 1 1481
0 1483 7 3 2 3600 1482
0 1484 5 2 1 3654
0 1485 7 1 2 3476 1246
0 1486 5 1 1 1485
0 1487 7 2 2 3480 1486
0 1488 5 1 1 3659
0 1489 7 1 2 3655 1488
0 1490 5 1 1 1489
0 1491 7 1 2 3657 3660
0 1492 5 1 1 1491
0 1493 7 1 2 3590 1392
0 1494 5 1 1 1493
0 1495 7 3 2 3594 1494
0 1496 5 2 1 3661
0 1497 7 1 2 3470 1238
0 1498 5 1 1 1497
0 1499 7 2 2 3474 1498
0 1500 5 1 1 3666
0 1501 7 1 2 3662 1500
0 1502 5 1 1 1501
0 1503 7 1 2 3664 3667
0 1504 5 1 1 1503
0 1505 7 1 2 3584 1384
0 1506 5 1 1 1505
0 1507 7 3 2 3588 1506
0 1508 5 2 1 3668
0 1509 7 1 2 3464 1230
0 1510 5 1 1 1509
0 1511 7 2 2 3468 1510
0 1512 5 1 1 3673
0 1513 7 1 2 3669 1512
0 1514 5 1 1 1513
0 1515 7 1 2 3671 3674
0 1516 5 1 1 1515
0 1517 7 1 2 3578 1376
0 1518 5 1 1 1517
0 1519 7 2 2 3582 1518
0 1520 5 2 1 3675
0 1521 7 1 2 3458 1222
0 1522 5 1 1 1521
0 1523 7 2 2 3462 1522
0 1524 5 1 1 3679
0 1525 7 1 2 3676 1524
0 1526 5 1 1 1525
0 1527 7 1 2 3677 3680
0 1528 5 1 1 1527
0 1529 7 1 2 3572 1368
0 1530 5 1 1 1529
0 1531 7 3 2 3576 1530
0 1532 5 2 1 3681
0 1533 7 1 2 3452 1214
0 1534 5 1 1 1533
0 1535 7 2 2 3456 1534
0 1536 5 1 1 3686
0 1537 7 1 2 3682 1536
0 1538 5 1 1 1537
0 1539 7 1 2 3684 3687
0 1540 5 1 1 1539
0 1541 7 1 2 3566 1360
0 1542 5 1 1 1541
0 1543 7 2 2 3570 1542
0 1544 5 2 1 3688
0 1545 7 1 2 3446 1206
0 1546 5 1 1 1545
0 1547 7 2 2 3450 1546
0 1548 5 1 1 3692
0 1549 7 1 2 3689 1548
0 1550 5 1 1 1549
0 1551 7 1 2 3690 3693
0 1552 5 1 1 1551
0 1553 7 1 2 3440 1198
0 1554 5 1 1 1553
0 1555 7 1 2 3444 1554
0 1556 5 1 1 1555
0 1557 7 1 2 3560 1352
0 1558 5 1 1 1557
0 1559 7 3 2 3564 1558
0 1560 5 2 1 3694
0 1561 7 1 2 3554 1344
0 1562 5 1 1 1561
0 1563 7 2 2 3558 1562
0 1564 5 2 1 3699
0 1565 7 1 2 3548 1336
0 1566 5 1 1 1565
0 1567 7 3 2 3552 1566
0 1568 5 1 1 3703
0 1569 7 1 2 3428 1182
0 1570 5 1 1 1569
0 1571 7 2 2 3432 1570
0 1572 5 1 1 3706
0 1573 7 1 2 1324 3543
0 1574 5 1 1 1573
0 1575 7 3 2 3546 1574
0 1576 5 1 1 3708
0 1577 7 1 2 3421 1174
0 1578 5 1 1 1577
0 1579 7 2 2 3426 1578
0 1580 5 1 1 3711
0 1581 7 2 2 3123 3134
0 1582 5 1 1 3713
0 1583 7 1 2 2877 3714
0 1584 5 1 1 1583
0 1585 7 1 2 3111 3125
0 1586 5 1 1 1585
0 1587 7 1 2 3544 1586
0 1588 5 1 1 1587
0 1589 7 2 2 1584 1588
0 1590 5 2 1 3715
0 1591 7 1 2 3119 3137
0 1592 5 1 1 1591
0 1593 7 2 2 1582 1592
0 1594 5 1 1 3719
0 1595 7 1 2 3401 3409
0 1596 5 2 1 1595
0 1597 7 1 2 3720 3721
0 1598 5 1 1 1597
0 1599 7 1 2 3405 3412
0 1600 5 1 1 1599
0 1601 7 2 2 1598 1600
0 1602 5 1 1 3723
0 1603 7 1 2 3394 3415
0 1604 5 1 1 1603
0 1605 7 2 2 3422 1604
0 1606 5 1 1 3725
0 1607 7 1 2 3724 3726
0 1608 5 1 1 1607
0 1609 7 1 2 3717 1608
0 1610 5 1 1 1609
0 1611 7 1 2 1602 1606
0 1612 5 1 1 1611
0 1613 7 2 2 1610 1612
0 1614 5 1 1 3727
0 1615 7 1 2 3712 3728
0 1616 5 1 1 1615
0 1617 7 1 2 3709 1616
0 1618 5 1 1 1617
0 1619 7 1 2 1580 1614
0 1620 5 1 1 1619
0 1621 7 2 2 1618 1620
0 1622 5 1 1 3729
0 1623 7 1 2 3707 3730
0 1624 5 1 1 1623
0 1625 7 1 2 3704 1624
0 1626 5 1 1 1625
0 1627 7 1 2 1572 1622
0 1628 5 1 1 1627
0 1629 7 2 2 1626 1628
0 1630 5 1 1 3731
0 1631 7 1 2 3701 3732
0 1632 5 1 1 1631
0 1633 7 1 2 3434 1190
0 1634 5 1 1 1633
0 1635 7 1 2 3700 1630
0 1636 5 1 1 1635
0 1637 7 1 2 3438 1636
0 1638 7 1 2 1634 1637
0 1639 5 1 1 1638
0 1640 7 2 2 1632 1639
0 1641 5 1 1 3733
0 1642 7 1 2 3697 1641
0 1643 5 1 1 1642
0 1644 7 1 2 1556 1643
0 1645 5 1 1 1644
0 1646 7 1 2 3695 3734
0 1647 5 1 1 1646
0 1648 7 1 2 1645 1647
0 1649 5 1 1 1648
0 1650 7 1 2 1552 1649
0 1651 5 1 1 1650
0 1652 7 1 2 1550 1651
0 1653 5 1 1 1652
0 1654 7 1 2 1540 1653
0 1655 5 1 1 1654
0 1656 7 1 2 1538 1655
0 1657 5 1 1 1656
0 1658 7 1 2 1528 1657
0 1659 5 1 1 1658
0 1660 7 1 2 1526 1659
0 1661 5 1 1 1660
0 1662 7 1 2 1516 1661
0 1663 5 1 1 1662
0 1664 7 1 2 1514 1663
0 1665 5 1 1 1664
0 1666 7 1 2 1504 1665
0 1667 5 1 1 1666
0 1668 7 1 2 1502 1667
0 1669 5 1 1 1668
0 1670 7 1 2 1492 1669
0 1671 5 1 1 1670
0 1672 7 1 2 1490 1671
0 1673 5 1 1 1672
0 1674 7 1 2 1480 1673
0 1675 5 1 1 1674
0 1676 7 1 2 1478 1675
0 1677 5 1 1 1676
0 1678 7 1 2 1468 1677
0 1679 5 1 1 1678
0 1680 7 1 2 1466 1679
0 1681 5 1 1 1680
0 1682 7 1 2 1456 1681
0 1683 5 1 1 1682
0 1684 7 1 2 1454 1683
0 1685 7 1 2 1444 1684
0 1686 5 1 1 1685
0 1687 7 1 2 1442 1686
0 1688 5 1 1 1687
0 1689 7 1 2 1432 1688
0 1690 5 1 1 1689
0 1691 7 1 2 3512 3623
0 1692 5 1 1 1691
0 1693 7 1 2 3233 3510
0 1694 7 1 2 1692 1693
0 1695 7 1 2 1690 1694
0 1696 5 1 1 1695
0 1697 7 1 2 3131 3410
0 1698 5 2 1 1697
0 1699 7 2 2 3128 3735
0 1700 5 2 1 3737
0 1701 7 1 2 3117 3739
0 1702 5 1 1 1701
0 1703 7 2 2 3114 1702
0 1704 5 2 1 3741
0 1705 7 1 2 3153 3743
0 1706 5 1 1 1705
0 1707 7 2 2 3105 1706
0 1708 5 2 1 3745
0 1709 7 1 2 3160 3747
0 1710 5 1 1 1709
0 1711 7 2 2 3095 1710
0 1712 5 2 1 3749
0 1713 7 1 2 3167 3751
0 1714 5 1 1 1713
0 1715 7 2 2 3085 1714
0 1716 5 2 1 3753
0 1717 7 1 2 3075 3755
0 1718 5 1 1 1717
0 1719 7 2 2 3072 1718
0 1720 5 2 1 3757
0 1721 7 1 2 3178 3759
0 1722 5 1 1 1721
0 1723 7 2 2 3062 1722
0 1724 5 2 1 3761
0 1725 7 1 2 3052 3763
0 1726 5 1 1 1725
0 1727 7 2 2 3049 1726
0 1728 5 2 1 3765
0 1729 7 1 2 3189 3767
0 1730 5 1 1 1729
0 1731 7 2 2 3039 1730
0 1732 5 2 1 3769
0 1733 7 1 2 3196 3771
0 1734 5 1 1 1733
0 1735 7 2 2 3029 1734
0 1736 5 2 1 3773
0 1737 7 1 2 3203 3775
0 1738 5 1 1 1737
0 1739 7 2 2 3019 1738
0 1740 5 2 1 3777
0 1741 7 1 2 3210 3779
0 1742 5 1 1 1741
0 1743 7 2 2 3009 1742
0 1744 5 2 1 3781
0 1745 7 1 2 3217 3783
0 1746 5 1 1 1745
0 1747 7 2 2 2999 1746
0 1748 5 2 1 3785
0 1749 7 1 2 3224 3787
0 1750 5 1 1 1749
0 1751 7 3 2 2989 1750
0 1752 5 3 1 3789
0 1753 7 1 2 2975 3792
0 1754 5 1 1 1753
0 1755 7 3 2 2980 1754
0 1756 5 2 1 3795
0 1757 7 1 2 1696 3798
0 1758 5 1 1 1757
0 1759 7 1 2 3279 3776
0 1760 5 1 1 1759
0 1761 7 1 2 3281 3774
0 1762 5 1 1 1761
0 1763 7 3 2 1760 1762
0 1764 5 2 1 3800
0 1765 7 1 2 3303 3768
0 1766 5 1 1 1765
0 1767 7 1 2 3305 3766
0 1768 5 1 1 1767
0 1769 7 3 2 1766 1768
0 1770 5 2 1 3805
0 1771 7 1 2 3803 3808
0 1772 5 2 1 1771
0 1773 7 1 2 3291 3772
0 1774 5 1 1 1773
0 1775 7 1 2 3293 3770
0 1776 5 1 1 1775
0 1777 7 3 2 1774 1776
0 1778 5 2 1 3812
0 1779 7 1 2 3315 3764
0 1780 5 1 1 1779
0 1781 7 1 2 3317 3762
0 1782 5 1 1 1781
0 1783 7 3 2 1780 1782
0 1784 5 2 1 3817
0 1785 7 1 2 3815 3820
0 1786 5 2 1 1785
0 1787 7 1 2 3327 3760
0 1788 5 1 1 1787
0 1789 7 1 2 3329 3758
0 1790 5 1 1 1789
0 1791 7 3 2 1788 1790
0 1792 5 2 1 3824
0 1793 7 1 2 3809 3827
0 1794 5 2 1 1793
0 1795 7 1 2 3339 3756
0 1796 5 1 1 1795
0 1797 7 1 2 3341 3754
0 1798 5 1 1 1797
0 1799 7 3 2 1796 1798
0 1800 5 2 1 3831
0 1801 7 1 2 3821 3834
0 1802 5 2 1 1801
0 1803 7 1 2 3351 3752
0 1804 5 1 1 1803
0 1805 7 1 2 3353 3750
0 1806 5 1 1 1805
0 1807 7 3 2 1804 1806
0 1808 5 2 1 3838
0 1809 7 1 2 3828 3841
0 1810 5 2 1 1809
0 1811 7 1 2 3363 3748
0 1812 5 1 1 1811
0 1813 7 1 2 3365 3746
0 1814 5 1 1 1813
0 1815 7 3 2 1812 1814
0 1816 5 2 1 3845
0 1817 7 1 2 3835 3848
0 1818 5 2 1 1817
0 1819 7 1 2 3375 3744
0 1820 5 1 1 1819
0 1821 7 1 2 3377 3742
0 1822 5 1 1 1821
0 1823 7 3 2 1820 1822
0 1824 5 2 1 3852
0 1825 7 1 2 3842 3855
0 1826 5 2 1 1825
0 1827 7 1 2 3387 3740
0 1828 5 1 1 1827
0 1829 7 1 2 3389 3738
0 1830 5 1 1 1829
0 1831 7 3 2 1828 1830
0 1832 5 2 1 3859
0 1833 7 1 2 3849 3862
0 1834 5 2 1 1833
0 1835 7 1 2 3399 3413
0 1836 5 1 1 1835
0 1837 7 3 2 3722 1836
0 1838 5 1 1 3866
0 1839 7 1 2 3856 3867
0 1840 5 2 1 1839
0 1841 7 2 2 3418 3863
0 1842 5 2 1 3871
0 1843 7 1 2 3853 1838
0 1844 5 1 1 1843
0 1845 7 2 2 3869 1844
0 1846 5 1 1 3875
0 1847 7 1 2 3872 3876
0 1848 5 2 1 1847
0 1849 7 2 2 3870 3877
0 1850 5 1 1 3879
0 1851 7 1 2 3846 3860
0 1852 5 1 1 1851
0 1853 7 2 2 3864 1852
0 1854 5 1 1 3881
0 1855 7 1 2 1850 3882
0 1856 5 2 1 1855
0 1857 7 2 2 3865 3883
0 1858 5 1 1 3885
0 1859 7 1 2 3839 3854
0 1860 5 1 1 1859
0 1861 7 2 2 3857 1860
0 1862 5 1 1 3887
0 1863 7 1 2 1858 3888
0 1864 5 2 1 1863
0 1865 7 2 2 3858 3889
0 1866 5 1 1 3891
0 1867 7 1 2 3832 3847
0 1868 5 1 1 1867
0 1869 7 2 2 3850 1868
0 1870 5 1 1 3893
0 1871 7 1 2 1866 3894
0 1872 5 2 1 1871
0 1873 7 2 2 3851 3895
0 1874 5 1 1 3897
0 1875 7 1 2 3825 3840
0 1876 5 1 1 1875
0 1877 7 2 2 3843 1876
0 1878 5 1 1 3899
0 1879 7 1 2 1874 3900
0 1880 5 2 1 1879
0 1881 7 2 2 3844 3901
0 1882 5 1 1 3903
0 1883 7 1 2 3818 3833
0 1884 5 1 1 1883
0 1885 7 2 2 3836 1884
0 1886 5 1 1 3905
0 1887 7 1 2 1882 3906
0 1888 5 2 1 1887
0 1889 7 2 2 3837 3907
0 1890 5 1 1 3909
0 1891 7 1 2 3806 3826
0 1892 5 1 1 1891
0 1893 7 2 2 3829 1892
0 1894 5 1 1 3911
0 1895 7 1 2 1890 3912
0 1896 5 2 1 1895
0 1897 7 2 2 3830 3913
0 1898 5 1 1 3915
0 1899 7 1 2 3813 3819
0 1900 5 1 1 1899
0 1901 7 2 2 3822 1900
0 1902 5 1 1 3917
0 1903 7 1 2 1898 3918
0 1904 5 2 1 1903
0 1905 7 2 2 3823 3919
0 1906 5 1 1 3921
0 1907 7 1 2 3801 3807
0 1908 5 1 1 1907
0 1909 7 2 2 3810 1908
0 1910 5 1 1 3923
0 1911 7 1 2 1906 3924
0 1912 5 2 1 1911
0 1913 7 2 2 3811 3925
0 1914 5 1 1 3927
0 1915 7 1 2 3267 3780
0 1916 5 1 1 1915
0 1917 7 1 2 3269 3778
0 1918 5 1 1 1917
0 1919 7 3 2 1916 1918
0 1920 5 2 1 3929
0 1921 7 1 2 3932 3816
0 1922 5 2 1 1921
0 1923 7 1 2 3930 3814
0 1924 5 1 1 1923
0 1925 7 2 2 3934 1924
0 1926 5 1 1 3936
0 1927 7 1 2 1914 3937
0 1928 5 2 1 1927
0 1929 7 1 2 3928 1926
0 1930 5 1 1 1929
0 1931 7 2 2 3938 1930
0 1932 5 1 1 3940
0 1933 7 1 2 3658 3941
0 1934 5 1 1 1933
0 1935 7 1 2 3922 1910
0 1936 5 1 1 1935
0 1937 7 2 2 3926 1936
0 1938 5 1 1 3942
0 1939 7 1 2 3663 1938
0 1940 5 1 1 1939
0 1941 7 1 2 3665 3943
0 1942 5 1 1 1941
0 1943 7 1 2 3916 1902
0 1944 5 1 1 1943
0 1945 7 2 2 3920 1944
0 1946 5 1 1 3944
0 1947 7 1 2 3670 1946
0 1948 5 1 1 1947
0 1949 7 1 2 3910 1894
0 1950 5 1 1 1949
0 1951 7 2 2 3914 1950
0 1952 5 1 1 3946
0 1953 7 1 2 3904 1886
0 1954 5 1 1 1953
0 1955 7 2 2 3908 1954
0 1956 5 1 1 3948
0 1957 7 1 2 3685 3949
0 1958 5 1 1 1957
0 1959 7 1 2 3683 1956
0 1960 5 1 1 1959
0 1961 7 1 2 3898 1878
0 1962 5 1 1 1961
0 1963 7 2 2 3902 1962
0 1964 5 1 1 3950
0 1965 7 1 2 3892 1870
0 1966 5 1 1 1965
0 1967 7 2 2 3896 1966
0 1968 5 1 1 3952
0 1969 7 1 2 3698 3953
0 1970 5 1 1 1969
0 1971 7 1 2 3696 1968
0 1972 5 1 1 1971
0 1973 7 1 2 3886 1862
0 1974 5 1 1 1973
0 1975 7 2 2 3890 1974
0 1976 5 1 1 3954
0 1977 7 1 2 3880 1854
0 1978 5 1 1 1977
0 1979 7 2 2 3884 1978
0 1980 5 1 1 3956
0 1981 7 1 2 1568 3957
0 1982 5 1 1 1981
0 1983 7 1 2 3705 1980
0 1984 5 1 1 1983
0 1985 7 1 2 3873 1846
0 1986 5 1 1 1985
0 1987 7 2 2 3878 1986
0 1988 5 1 1 3958
0 1989 7 1 2 1576 3959
0 1990 5 1 1 1989
0 1991 7 1 2 3710 1988
0 1992 5 1 1 1991
0 1993 7 1 2 3416 3861
0 1994 5 1 1 1993
0 1995 7 1 2 1594 3868
0 1996 5 1 1 1995
0 1997 7 2 2 3736 1996
0 1998 5 1 1 3960
0 1999 7 1 2 3718 3961
0 2000 5 1 1 1999
0 2001 7 1 2 3874 2000
0 2002 7 1 2 1994 2001
0 2003 5 1 1 2002
0 2004 7 1 2 3716 1998
0 2005 5 1 1 2004
0 2006 7 1 2 2003 2005
0 2007 5 1 1 2006
0 2008 7 1 2 1992 2007
0 2009 5 1 1 2008
0 2010 7 1 2 1990 2009
0 2011 5 1 1 2010
0 2012 7 1 2 1984 2011
0 2013 5 1 1 2012
0 2014 7 2 2 1982 2013
0 2015 5 1 1 3962
0 2016 7 1 2 3955 2015
0 2017 5 1 1 2016
0 2018 7 1 2 1976 3963
0 2019 5 1 1 2018
0 2020 7 1 2 3702 2019
0 2021 5 1 1 2020
0 2022 7 1 2 2017 2021
0 2023 5 1 1 2022
0 2024 7 1 2 1972 2023
0 2025 5 1 1 2024
0 2026 7 2 2 1970 2025
0 2027 5 1 1 3964
0 2028 7 1 2 3951 2027
0 2029 5 1 1 2028
0 2030 7 1 2 1964 3965
0 2031 5 1 1 2030
0 2032 7 1 2 3691 2031
0 2033 5 1 1 2032
0 2034 7 1 2 2029 2033
0 2035 5 1 1 2034
0 2036 7 1 2 1960 2035
0 2037 5 1 1 2036
0 2038 7 2 2 1958 2037
0 2039 5 1 1 3966
0 2040 7 1 2 1952 3967
0 2041 5 1 1 2040
0 2042 7 1 2 3678 2041
0 2043 5 1 1 2042
0 2044 7 1 2 3947 2039
0 2045 5 1 1 2044
0 2046 7 1 2 3672 3945
0 2047 5 1 1 2046
0 2048 7 1 2 2045 2047
0 2049 7 1 2 2043 2048
0 2050 5 1 1 2049
0 2051 7 1 2 1948 2050
0 2052 5 1 1 2051
0 2053 7 1 2 1942 2052
0 2054 5 1 1 2053
0 2055 7 1 2 1940 2054
0 2056 5 1 1 2055
0 2057 7 1 2 1934 2056
0 2058 5 1 1 2057
0 2059 7 1 2 3656 1932
0 2060 5 1 1 2059
0 2061 7 2 2 3935 3939
0 2062 5 1 1 3968
0 2063 7 1 2 3248 3784
0 2064 5 1 1 2063
0 2065 7 1 2 3250 3782
0 2066 5 1 1 2065
0 2067 7 3 2 2064 2066
0 2068 5 2 1 3970
0 2069 7 1 2 3973 3804
0 2070 5 2 1 2069
0 2071 7 1 2 3971 3802
0 2072 5 1 1 2071
0 2073 7 2 2 3975 2072
0 2074 5 1 1 3977
0 2075 7 1 2 2062 3978
0 2076 5 2 1 2075
0 2077 7 1 2 3969 2074
0 2078 5 1 1 2077
0 2079 7 2 2 3979 2078
0 2080 5 1 1 3981
0 2081 7 1 2 3649 2080
0 2082 5 1 1 2081
0 2083 7 1 2 2060 2082
0 2084 7 1 2 2058 2083
0 2085 5 1 1 2084
0 2086 7 2 2 3976 3980
0 2087 5 1 1 3983
0 2088 7 1 2 3236 3788
0 2089 5 1 1 2088
0 2090 7 1 2 3238 3786
0 2091 5 1 1 2090
0 2092 7 3 2 2089 2091
0 2093 5 2 1 3985
0 2094 7 1 2 3933 3988
0 2095 5 2 1 2094
0 2096 7 1 2 3931 3986
0 2097 5 1 1 2096
0 2098 7 2 2 3990 2097
0 2099 5 1 1 3992
0 2100 7 1 2 2087 3993
0 2101 5 2 1 2100
0 2102 7 1 2 3984 2099
0 2103 5 1 1 2102
0 2104 7 2 2 3994 2103
0 2105 5 1 1 3996
0 2106 7 1 2 3644 3997
0 2107 5 1 1 2106
0 2108 7 1 2 3651 3982
0 2109 5 1 1 2108
0 2110 7 1 2 2107 2109
0 2111 7 1 2 2085 2110
0 2112 5 1 1 2111
0 2113 7 2 2 3991 3995
0 2114 5 1 1 3998
0 2115 7 1 2 3258 3793
0 2116 5 1 1 2115
0 2117 7 1 2 3260 3790
0 2118 5 1 1 2117
0 2119 7 2 2 2116 2118
0 2120 5 1 1 4000
0 2121 7 1 2 2120 3974
0 2122 5 2 1 2121
0 2123 7 1 2 4001 3972
0 2124 5 1 1 2123
0 2125 7 2 2 4002 2124
0 2126 5 1 1 4004
0 2127 7 1 2 2114 4005
0 2128 5 2 1 2127
0 2129 7 1 2 3999 2126
0 2130 5 1 1 2129
0 2131 7 2 2 4006 2130
0 2132 5 1 1 4008
0 2133 7 1 2 3635 2132
0 2134 5 1 1 2133
0 2135 7 1 2 3642 2105
0 2136 5 1 1 2135
0 2137 7 1 2 2134 2136
0 2138 7 1 2 2112 2137
0 2139 5 1 1 2138
0 2140 7 2 2 4003 4007
0 2141 5 1 1 4010
0 2142 7 1 2 3796 3987
0 2143 5 1 1 2142
0 2144 7 1 2 3799 3989
0 2145 5 1 1 2144
0 2146 7 2 2 2143 2145
0 2147 5 1 1 4012
0 2148 7 1 2 2141 4013
0 2149 5 1 1 2148
0 2150 7 1 2 2976 3791
0 2151 5 1 1 2150
0 2152 7 1 2 2981 3794
0 2153 5 1 1 2152
0 2154 7 1 2 2151 2153
0 2155 5 2 1 2154
0 2156 7 2 2 2149 4014
0 2157 5 1 1 4016
0 2158 7 1 2 3624 2157
0 2159 5 1 1 2158
0 2160 7 1 2 3637 4009
0 2161 5 1 1 2160
0 2162 7 2 2 4011 2147
0 2163 5 1 1 4018
0 2164 7 1 2 3629 4015
0 2165 5 1 1 2164
0 2166 7 1 2 2163 2165
0 2167 5 1 1 2166
0 2168 7 1 2 2161 2167
0 2169 7 1 2 2159 2168
0 2170 7 1 2 2139 2169
0 2171 5 1 1 2170
0 2172 7 1 2 3630 4019
0 2173 5 1 1 2172
0 2174 7 1 2 3625 2173
0 2175 5 1 1 2174
0 2176 7 1 2 4017 2175
0 2177 5 1 1 2176
0 2178 7 1 2 3797 2177
0 2179 7 1 2 2171 2178
0 2180 5 1 1 2179
3 4299 7 0 2 1758 2180
