1 0 0 8 0
2 32 1 0
2 1972 1 0
2 1973 1 0
2 1974 1 0
2 1975 1 0
2 1976 1 0
2 1977 1 0
2 1978 1 0
1 1 0 8 0
2 1979 1 1
2 1980 1 1
2 1981 1 1
2 1982 1 1
2 1983 1 1
2 1984 1 1
2 1985 1 1
2 1986 1 1
1 2 0 8 0
2 1987 1 2
2 1988 1 2
2 1989 1 2
2 1990 1 2
2 1991 1 2
2 1992 1 2
2 1993 1 2
2 1994 1 2
1 3 0 9 0
2 1995 1 3
2 1996 1 3
2 1997 1 3
2 1998 1 3
2 1999 1 3
2 2000 1 3
2 2001 1 3
2 2002 1 3
2 2003 1 3
1 4 0 8 0
2 2004 1 4
2 2005 1 4
2 2006 1 4
2 2007 1 4
2 2008 1 4
2 2009 1 4
2 2010 1 4
2 2011 1 4
1 5 0 9 0
2 2012 1 5
2 2013 1 5
2 2014 1 5
2 2015 1 5
2 2016 1 5
2 2017 1 5
2 2018 1 5
2 2019 1 5
2 2020 1 5
1 6 0 8 0
2 2021 1 6
2 2022 1 6
2 2023 1 6
2 2024 1 6
2 2025 1 6
2 2026 1 6
2 2027 1 6
2 2028 1 6
1 7 0 8 0
2 2029 1 7
2 2030 1 7
2 2031 1 7
2 2032 1 7
2 2033 1 7
2 2034 1 7
2 2035 1 7
2 2036 1 7
1 8 0 8 0
2 2037 1 8
2 2038 1 8
2 2039 1 8
2 2040 1 8
2 2041 1 8
2 2042 1 8
2 2043 1 8
2 2044 1 8
1 9 0 8 0
2 2045 1 9
2 2046 1 9
2 2047 1 9
2 2048 1 9
2 2049 1 9
2 2050 1 9
2 2051 1 9
2 2052 1 9
1 10 0 9 0
2 2053 1 10
2 2054 1 10
2 2055 1 10
2 2056 1 10
2 2057 1 10
2 2058 1 10
2 2059 1 10
2 2060 1 10
2 2061 1 10
1 11 0 8 0
2 2062 1 11
2 2063 1 11
2 2064 1 11
2 2065 1 11
2 2066 1 11
2 2067 1 11
2 2068 1 11
2 2069 1 11
1 12 0 8 0
2 2070 1 12
2 2071 1 12
2 2072 1 12
2 2073 1 12
2 2074 1 12
2 2075 1 12
2 2076 1 12
2 2077 1 12
1 13 0 8 0
2 2078 1 13
2 2079 1 13
2 2080 1 13
2 2081 1 13
2 2082 1 13
2 2083 1 13
2 2084 1 13
2 2085 1 13
1 14 0 8 0
2 2086 1 14
2 2087 1 14
2 2088 1 14
2 2089 1 14
2 2090 1 14
2 2091 1 14
2 2092 1 14
2 2093 1 14
1 15 0 8 0
2 2094 1 15
2 2095 1 15
2 2096 1 15
2 2097 1 15
2 2098 1 15
2 2099 1 15
2 2100 1 15
2 2101 1 15
1 16 0 2 0
2 2102 1 16
2 2103 1 16
1 17 0 2 0
2 2104 1 17
2 2105 1 17
1 18 0 2 0
2 2106 1 18
2 2107 1 18
1 19 0 2 0
2 2108 1 19
2 2109 1 19
1 20 0 2 0
2 2110 1 20
2 2111 1 20
1 21 0 2 0
2 2112 1 21
2 2113 1 21
1 22 0 2 0
2 2114 1 22
2 2115 1 22
1 23 0 2 0
2 2116 1 23
2 2117 1 23
1 24 0 2 0
2 2118 1 24
2 2119 1 24
1 25 0 2 0
2 2120 1 25
2 2121 1 25
1 26 0 2 0
2 2122 1 26
2 2123 1 26
1 27 0 2 0
2 2124 1 27
2 2125 1 27
1 28 0 2 0
2 2126 1 28
2 2127 1 28
1 29 0 2 0
2 2128 1 29
2 2129 1 29
1 30 0 2 0
2 2130 1 30
2 2131 1 30
1 31 0 2 0
2 2132 1 31
2 2133 1 31
2 2134 1 49
2 2135 1 49
2 2136 1 51
2 2137 1 51
2 2138 1 52
2 2139 1 52
2 2140 1 53
2 2141 1 53
2 2142 1 55
2 2143 1 55
2 2144 1 58
2 2145 1 58
2 2146 1 61
2 2147 1 61
2 2148 1 64
2 2149 1 64
2 2150 1 65
2 2151 1 65
2 2152 1 67
2 2153 1 67
2 2154 1 69
2 2155 1 69
2 2156 1 75
2 2157 1 75
2 2158 1 78
2 2159 1 78
2 2160 1 78
2 2161 1 82
2 2162 1 82
2 2163 1 83
2 2164 1 83
2 2165 1 85
2 2166 1 85
2 2167 1 88
2 2168 1 88
2 2169 1 89
2 2170 1 89
2 2171 1 93
2 2172 1 93
2 2173 1 96
2 2174 1 96
2 2175 1 97
2 2176 1 97
2 2177 1 101
2 2178 1 101
2 2179 1 104
2 2180 1 104
2 2181 1 105
2 2182 1 105
2 2183 1 109
2 2184 1 109
2 2185 1 112
2 2186 1 112
2 2187 1 113
2 2188 1 113
2 2189 1 115
2 2190 1 115
2 2191 1 118
2 2192 1 118
2 2193 1 119
2 2194 1 119
2 2195 1 123
2 2196 1 123
2 2197 1 126
2 2198 1 126
2 2199 1 127
2 2200 1 127
2 2201 1 131
2 2202 1 131
2 2203 1 134
2 2204 1 134
2 2205 1 135
2 2206 1 135
2 2207 1 139
2 2208 1 139
2 2209 1 142
2 2210 1 142
2 2211 1 143
2 2212 1 143
2 2213 1 147
2 2214 1 147
2 2215 1 150
2 2216 1 150
2 2217 1 151
2 2218 1 151
2 2219 1 155
2 2220 1 155
2 2221 1 158
2 2222 1 158
2 2223 1 159
2 2224 1 159
2 2225 1 163
2 2226 1 163
2 2227 1 166
2 2228 1 166
2 2229 1 167
2 2230 1 167
2 2231 1 171
2 2232 1 171
2 2233 1 174
2 2234 1 174
2 2235 1 175
2 2236 1 175
2 2237 1 177
2 2238 1 177
2 2239 1 179
2 2240 1 179
2 2241 1 181
2 2242 1 181
2 2243 1 182
2 2244 1 182
2 2245 1 183
2 2246 1 183
2 2247 1 184
2 2248 1 184
2 2249 1 186
2 2250 1 186
2 2251 1 187
2 2252 1 187
2 2253 1 191
2 2254 1 191
2 2255 1 194
2 2256 1 194
2 2257 1 195
2 2258 1 195
2 2259 1 199
2 2260 1 199
2 2261 1 202
2 2262 1 202
2 2263 1 203
2 2264 1 203
2 2265 1 207
2 2266 1 207
2 2267 1 210
2 2268 1 210
2 2269 1 211
2 2270 1 211
2 2271 1 215
2 2272 1 215
2 2273 1 218
2 2274 1 218
2 2275 1 219
2 2276 1 219
2 2277 1 223
2 2278 1 223
2 2279 1 226
2 2280 1 226
2 2281 1 227
2 2282 1 227
2 2283 1 231
2 2284 1 231
2 2285 1 234
2 2286 1 234
2 2287 1 235
2 2288 1 235
2 2289 1 239
2 2290 1 239
2 2291 1 242
2 2292 1 242
2 2293 1 243
2 2294 1 243
2 2295 1 245
2 2296 1 245
2 2297 1 248
2 2298 1 248
2 2299 1 251
2 2300 1 251
2 2301 1 255
2 2302 1 255
2 2303 1 258
2 2304 1 258
2 2305 1 259
2 2306 1 259
2 2307 1 263
2 2308 1 263
2 2309 1 266
2 2310 1 266
2 2311 1 267
2 2312 1 267
2 2313 1 269
2 2314 1 269
2 2315 1 272
2 2316 1 272
2 2317 1 273
2 2318 1 273
2 2319 1 275
2 2320 1 275
2 2321 1 281
2 2322 1 281
2 2323 1 284
2 2324 1 284
2 2325 1 287
2 2326 1 287
2 2327 1 290
2 2328 1 290
2 2329 1 293
2 2330 1 293
2 2331 1 297
2 2332 1 297
2 2333 1 300
2 2334 1 300
2 2335 1 301
2 2336 1 301
2 2337 1 305
2 2338 1 305
2 2339 1 308
2 2340 1 308
2 2341 1 309
2 2342 1 309
2 2343 1 311
2 2344 1 311
2 2345 1 314
2 2346 1 314
2 2347 1 317
2 2348 1 317
2 2349 1 321
2 2350 1 321
2 2351 1 324
2 2352 1 324
2 2353 1 325
2 2354 1 325
2 2355 1 329
2 2356 1 329
2 2357 1 332
2 2358 1 332
2 2359 1 333
2 2360 1 333
2 2361 1 337
2 2362 1 337
2 2363 1 340
2 2364 1 340
2 2365 1 341
2 2366 1 341
2 2367 1 345
2 2368 1 345
2 2369 1 348
2 2370 1 348
2 2371 1 349
2 2372 1 349
2 2373 1 353
2 2374 1 353
2 2375 1 356
2 2376 1 356
2 2377 1 357
2 2378 1 357
2 2379 1 359
2 2380 1 359
2 2381 1 362
2 2382 1 362
2 2383 1 363
2 2384 1 363
2 2385 1 367
2 2386 1 367
2 2387 1 370
2 2388 1 370
2 2389 1 371
2 2390 1 371
2 2391 1 373
2 2392 1 373
2 2393 1 375
2 2394 1 375
2 2395 1 378
2 2396 1 378
2 2397 1 379
2 2398 1 379
2 2399 1 381
2 2400 1 381
2 2401 1 383
2 2402 1 383
2 2403 1 385
2 2404 1 385
2 2405 1 387
2 2406 1 387
2 2407 1 388
2 2408 1 388
2 2409 1 389
2 2410 1 389
2 2411 1 390
2 2412 1 390
2 2413 1 391
2 2414 1 391
2 2415 1 392
2 2416 1 392
2 2417 1 393
2 2418 1 393
2 2419 1 394
2 2420 1 394
2 2421 1 396
2 2422 1 396
2 2423 1 399
2 2424 1 399
2 2425 1 403
2 2426 1 403
2 2427 1 406
2 2428 1 406
2 2429 1 409
2 2430 1 409
2 2431 1 413
2 2432 1 413
2 2433 1 416
2 2434 1 416
2 2435 1 417
2 2436 1 417
2 2437 1 420
2 2438 1 420
2 2439 1 421
2 2440 1 421
2 2441 1 425
2 2442 1 425
2 2443 1 428
2 2444 1 428
2 2445 1 429
2 2446 1 429
2 2447 1 433
2 2448 1 433
2 2449 1 436
2 2450 1 436
2 2451 1 437
2 2452 1 437
2 2453 1 441
2 2454 1 441
2 2455 1 444
2 2456 1 444
2 2457 1 447
2 2458 1 447
2 2459 1 451
2 2460 1 451
2 2461 1 454
2 2462 1 454
2 2463 1 457
2 2464 1 457
2 2465 1 461
2 2466 1 461
2 2467 1 464
2 2468 1 464
2 2469 1 465
2 2470 1 465
2 2471 1 467
2 2472 1 467
2 2473 1 470
2 2474 1 470
2 2475 1 471
2 2476 1 471
2 2477 1 475
2 2478 1 475
2 2479 1 478
2 2480 1 478
2 2481 1 479
2 2482 1 479
2 2483 1 483
2 2484 1 483
2 2485 1 486
2 2486 1 486
2 2487 1 487
2 2488 1 487
2 2489 1 491
2 2490 1 491
2 2491 1 494
2 2492 1 494
2 2493 1 495
2 2494 1 495
2 2495 1 499
2 2496 1 499
2 2497 1 502
2 2498 1 502
2 2499 1 503
2 2500 1 503
2 2501 1 507
2 2502 1 507
2 2503 1 510
2 2504 1 510
2 2505 1 511
2 2506 1 511
2 2507 1 513
2 2508 1 513
2 2509 1 519
2 2510 1 519
2 2511 1 522
2 2512 1 522
2 2513 1 525
2 2514 1 525
2 2515 1 528
2 2516 1 528
2 2517 1 531
2 2518 1 531
2 2519 1 535
2 2520 1 535
2 2521 1 538
2 2522 1 538
2 2523 1 539
2 2524 1 539
2 2525 1 543
2 2526 1 543
2 2527 1 546
2 2528 1 546
2 2529 1 547
2 2530 1 547
2 2531 1 551
2 2532 1 551
2 2533 1 554
2 2534 1 554
2 2535 1 555
2 2536 1 555
2 2537 1 559
2 2538 1 559
2 2539 1 562
2 2540 1 562
2 2541 1 563
2 2542 1 563
2 2543 1 567
2 2544 1 567
2 2545 1 570
2 2546 1 570
2 2547 1 571
2 2548 1 571
2 2549 1 575
2 2550 1 575
2 2551 1 578
2 2552 1 578
2 2553 1 579
2 2554 1 579
2 2555 1 583
2 2556 1 583
2 2557 1 586
2 2558 1 586
2 2559 1 587
2 2560 1 587
2 2561 1 589
2 2562 1 589
2 2563 1 592
2 2564 1 592
2 2565 1 595
2 2566 1 595
2 2567 1 599
2 2568 1 599
2 2569 1 602
2 2570 1 602
2 2571 1 603
2 2572 1 603
2 2573 1 607
2 2574 1 607
2 2575 1 610
2 2576 1 610
2 2577 1 611
2 2578 1 611
2 2579 1 615
2 2580 1 615
2 2581 1 618
2 2582 1 618
2 2583 1 619
2 2584 1 619
2 2585 1 623
2 2586 1 623
2 2587 1 626
2 2588 1 626
2 2589 1 627
2 2590 1 627
2 2591 1 633
2 2592 1 633
2 2593 1 636
2 2594 1 636
2 2595 1 637
2 2596 1 637
2 2597 1 641
2 2598 1 641
2 2599 1 644
2 2600 1 644
2 2601 1 645
2 2602 1 645
2 2603 1 649
2 2604 1 649
2 2605 1 652
2 2606 1 652
2 2607 1 653
2 2608 1 653
2 2609 1 657
2 2610 1 657
2 2611 1 660
2 2612 1 660
2 2613 1 661
2 2614 1 661
2 2615 1 663
2 2616 1 663
2 2617 1 666
2 2618 1 666
2 2619 1 669
2 2620 1 669
2 2621 1 673
2 2622 1 673
2 2623 1 676
2 2624 1 676
2 2625 1 677
2 2626 1 677
2 2627 1 681
2 2628 1 681
2 2629 1 684
2 2630 1 684
2 2631 1 687
2 2632 1 687
2 2633 1 689
2 2634 1 689
2 2635 1 691
2 2636 1 691
2 2637 1 693
2 2638 1 693
2 2639 1 695
2 2640 1 695
2 2641 1 697
2 2642 1 697
2 2643 1 699
2 2644 1 699
2 2645 1 700
2 2646 1 700
2 2647 1 701
2 2648 1 701
2 2649 1 701
2 2650 1 704
2 2651 1 704
2 2652 1 707
2 2653 1 707
2 2654 1 715
2 2655 1 715
2 2656 1 718
2 2657 1 718
2 2658 1 719
2 2659 1 719
2 2660 1 723
2 2661 1 723
2 2662 1 726
2 2663 1 726
2 2664 1 729
2 2665 1 729
2 2666 1 731
2 2667 1 731
2 2668 1 733
2 2669 1 733
2 2670 1 735
2 2671 1 735
2 2672 1 736
2 2673 1 736
2 2674 1 738
2 2675 1 738
2 2676 1 739
2 2677 1 739
2 2678 1 743
2 2679 1 743
2 2680 1 746
2 2681 1 746
2 2682 1 747
2 2683 1 747
2 2684 1 751
2 2685 1 751
2 2686 1 754
2 2687 1 754
2 2688 1 755
2 2689 1 755
2 2690 1 759
2 2691 1 759
2 2692 1 762
2 2693 1 762
2 2694 1 763
2 2695 1 763
2 2696 1 767
2 2697 1 767
2 2698 1 770
2 2699 1 770
2 2700 1 771
2 2701 1 771
2 2702 1 775
2 2703 1 775
2 2704 1 778
2 2705 1 778
2 2706 1 779
2 2707 1 779
2 2708 1 783
2 2709 1 783
2 2710 1 786
2 2711 1 786
2 2712 1 787
2 2713 1 787
2 2714 1 791
2 2715 1 791
2 2716 1 794
2 2717 1 794
2 2718 1 795
2 2719 1 795
2 2720 1 799
2 2721 1 799
2 2722 1 802
2 2723 1 802
2 2724 1 803
2 2725 1 803
2 2726 1 807
2 2727 1 807
2 2728 1 810
2 2729 1 810
2 2730 1 811
2 2731 1 811
2 2732 1 815
2 2733 1 815
2 2734 1 818
2 2735 1 818
2 2736 1 819
2 2737 1 819
2 2738 1 823
2 2739 1 823
2 2740 1 826
2 2741 1 826
2 2742 1 827
2 2743 1 827
2 2744 1 831
2 2745 1 831
2 2746 1 834
2 2747 1 834
2 2748 1 835
2 2749 1 835
2 2750 1 835
2 2751 1 835
2 2752 1 836
2 2753 1 836
2 2754 1 836
2 2755 1 837
2 2756 1 837
2 2757 1 837
2 2758 1 838
2 2759 1 838
2 2760 1 838
2 2761 1 839
2 2762 1 839
2 2763 1 839
2 2764 1 840
2 2765 1 840
2 2766 1 840
2 2767 1 843
2 2768 1 843
2 2769 1 843
2 2770 1 843
2 2771 1 844
2 2772 1 844
2 2773 1 844
2 2774 1 846
2 2775 1 846
2 2776 1 846
2 2777 1 848
2 2778 1 848
2 2779 1 848
2 2780 1 851
2 2781 1 851
2 2782 1 851
2 2783 1 851
2 2784 1 852
2 2785 1 852
2 2786 1 852
2 2787 1 854
2 2788 1 854
2 2789 1 854
2 2790 1 856
2 2791 1 856
2 2792 1 856
2 2793 1 859
2 2794 1 859
2 2795 1 859
2 2796 1 859
2 2797 1 860
2 2798 1 860
2 2799 1 860
2 2800 1 862
2 2801 1 862
2 2802 1 862
2 2803 1 864
2 2804 1 864
2 2805 1 864
2 2806 1 867
2 2807 1 867
2 2808 1 867
2 2809 1 867
2 2810 1 868
2 2811 1 868
2 2812 1 868
2 2813 1 870
2 2814 1 870
2 2815 1 870
2 2816 1 872
2 2817 1 872
2 2818 1 872
2 2819 1 875
2 2820 1 875
2 2821 1 875
2 2822 1 875
2 2823 1 876
2 2824 1 876
2 2825 1 876
2 2826 1 878
2 2827 1 878
2 2828 1 878
2 2829 1 880
2 2830 1 880
2 2831 1 880
2 2832 1 883
2 2833 1 883
2 2834 1 883
2 2835 1 883
2 2836 1 884
2 2837 1 884
2 2838 1 884
2 2839 1 886
2 2840 1 886
2 2841 1 886
2 2842 1 888
2 2843 1 888
2 2844 1 888
2 2845 1 891
2 2846 1 891
2 2847 1 891
2 2848 1 891
2 2849 1 892
2 2850 1 892
2 2851 1 892
2 2852 1 894
2 2853 1 894
2 2854 1 894
2 2855 1 896
2 2856 1 896
2 2857 1 896
2 2858 1 899
2 2859 1 899
2 2860 1 899
2 2861 1 899
2 2862 1 900
2 2863 1 900
2 2864 1 900
2 2865 1 902
2 2866 1 902
2 2867 1 902
2 2868 1 904
2 2869 1 904
2 2870 1 904
2 2871 1 907
2 2872 1 907
2 2873 1 907
2 2874 1 907
2 2875 1 908
2 2876 1 908
2 2877 1 908
2 2878 1 910
2 2879 1 910
2 2880 1 910
2 2881 1 912
2 2882 1 912
2 2883 1 912
2 2884 1 915
2 2885 1 915
2 2886 1 915
2 2887 1 915
2 2888 1 916
2 2889 1 916
2 2890 1 916
2 2891 1 918
2 2892 1 918
2 2893 1 918
2 2894 1 920
2 2895 1 920
2 2896 1 920
2 2897 1 923
2 2898 1 923
2 2899 1 923
2 2900 1 923
2 2901 1 924
2 2902 1 924
2 2903 1 924
2 2904 1 926
2 2905 1 926
2 2906 1 926
2 2907 1 928
2 2908 1 928
2 2909 1 928
2 2910 1 931
2 2911 1 931
2 2912 1 931
2 2913 1 931
2 2914 1 932
2 2915 1 932
2 2916 1 932
2 2917 1 934
2 2918 1 934
2 2919 1 934
2 2920 1 936
2 2921 1 936
2 2922 1 936
2 2923 1 939
2 2924 1 939
2 2925 1 940
2 2926 1 940
2 2927 1 940
2 2928 1 942
2 2929 1 942
2 2930 1 942
2 2931 1 944
2 2932 1 944
2 2933 1 944
2 2934 1 947
2 2935 1 947
2 2936 1 947
2 2937 1 947
2 2938 1 948
2 2939 1 948
2 2940 1 948
2 2941 1 950
2 2942 1 950
2 2943 1 950
2 2944 1 952
2 2945 1 952
2 2946 1 952
2 2947 1 952
2 2948 1 953
2 2949 1 953
2 2950 1 953
2 2951 1 954
2 2952 1 954
2 2953 1 955
2 2954 1 955
2 2955 1 956
2 2956 1 956
2 2957 1 956
2 2958 1 956
2 2959 1 959
2 2960 1 959
2 2961 1 960
2 2962 1 960
2 2963 1 963
2 2964 1 963
2 2965 1 964
2 2966 1 964
2 2967 1 967
2 2968 1 967
2 2969 1 968
2 2970 1 968
2 2971 1 971
2 2972 1 971
2 2973 1 972
2 2974 1 972
2 2975 1 975
2 2976 1 975
2 2977 1 976
2 2978 1 976
2 2979 1 979
2 2980 1 979
2 2981 1 980
2 2982 1 980
2 2983 1 983
2 2984 1 983
2 2985 1 984
2 2986 1 984
2 2987 1 987
2 2988 1 987
2 2989 1 988
2 2990 1 988
2 2991 1 991
2 2992 1 991
2 2993 1 992
2 2994 1 992
2 2995 1 995
2 2996 1 995
2 2997 1 996
2 2998 1 996
2 2999 1 999
2 3000 1 999
2 3001 1 1000
2 3002 1 1000
2 3003 1 1003
2 3004 1 1003
2 3005 1 1004
2 3006 1 1004
2 3007 1 1007
2 3008 1 1007
2 3009 1 1008
2 3010 1 1008
2 3011 1 1011
2 3012 1 1011
2 3013 1 1011
2 3014 1 1011
2 3015 1 1012
2 3016 1 1012
2 3017 1 1014
2 3018 1 1014
2 3019 1 1015
2 3020 1 1015
2 3021 1 1017
2 3022 1 1017
2 3023 1 1017
2 3024 1 1018
2 3025 1 1018
2 3026 1 1023
2 3027 1 1023
2 3028 1 1023
2 3029 1 1024
2 3030 1 1024
2 3031 1 1026
2 3032 1 1026
2 3033 1 1027
2 3034 1 1027
2 3035 1 1027
2 3036 1 1028
2 3037 1 1028
2 3038 1 1033
2 3039 1 1033
2 3040 1 1035
2 3041 1 1035
2 3042 1 1035
2 3043 1 1036
2 3044 1 1036
2 3045 1 1041
2 3046 1 1041
2 3047 1 1041
2 3048 1 1042
2 3049 1 1042
2 3050 1 1044
2 3051 1 1044
2 3052 1 1045
2 3053 1 1045
2 3054 1 1045
2 3055 1 1046
2 3056 1 1046
2 3057 1 1051
2 3058 1 1051
2 3059 1 1051
2 3060 1 1052
2 3061 1 1052
2 3062 1 1054
2 3063 1 1054
2 3064 1 1055
2 3065 1 1055
2 3066 1 1055
2 3067 1 1056
2 3068 1 1056
2 3069 1 1061
2 3070 1 1061
2 3071 1 1061
2 3072 1 1062
2 3073 1 1062
2 3074 1 1064
2 3075 1 1064
2 3076 1 1065
2 3077 1 1065
2 3078 1 1065
2 3079 1 1066
2 3080 1 1066
2 3081 1 1071
2 3082 1 1071
2 3083 1 1071
2 3084 1 1072
2 3085 1 1072
2 3086 1 1074
2 3087 1 1074
2 3088 1 1075
2 3089 1 1075
2 3090 1 1075
2 3091 1 1076
2 3092 1 1076
2 3093 1 1081
2 3094 1 1081
2 3095 1 1081
2 3096 1 1082
2 3097 1 1082
2 3098 1 1084
2 3099 1 1084
2 3100 1 1085
2 3101 1 1085
2 3102 1 1085
2 3103 1 1086
2 3104 1 1086
2 3105 1 1091
2 3106 1 1091
2 3107 1 1091
2 3108 1 1092
2 3109 1 1092
2 3110 1 1094
2 3111 1 1094
2 3112 1 1095
2 3113 1 1095
2 3114 1 1095
2 3115 1 1096
2 3116 1 1096
2 3117 1 1101
2 3118 1 1101
2 3119 1 1101
2 3120 1 1102
2 3121 1 1102
2 3122 1 1104
2 3123 1 1104
2 3124 1 1105
2 3125 1 1105
2 3126 1 1105
2 3127 1 1106
2 3128 1 1106
2 3129 1 1111
2 3130 1 1111
2 3131 1 1111
2 3132 1 1112
2 3133 1 1112
2 3134 1 1114
2 3135 1 1114
2 3136 1 1115
2 3137 1 1115
2 3138 1 1115
2 3139 1 1116
2 3140 1 1116
2 3141 1 1121
2 3142 1 1121
2 3143 1 1121
2 3144 1 1122
2 3145 1 1122
2 3146 1 1124
2 3147 1 1124
2 3148 1 1125
2 3149 1 1125
2 3150 1 1125
2 3151 1 1126
2 3152 1 1126
2 3153 1 1131
2 3154 1 1131
2 3155 1 1131
2 3156 1 1132
2 3157 1 1132
2 3158 1 1134
2 3159 1 1134
2 3160 1 1135
2 3161 1 1135
2 3162 1 1135
2 3163 1 1136
2 3164 1 1136
2 3165 1 1141
2 3166 1 1141
2 3167 1 1141
2 3168 1 1142
2 3169 1 1142
2 3170 1 1144
2 3171 1 1144
2 3172 1 1145
2 3173 1 1145
2 3174 1 1145
2 3175 1 1146
2 3176 1 1146
2 3177 1 1151
2 3178 1 1151
2 3179 1 1151
2 3180 1 1152
2 3181 1 1152
2 3182 1 1154
2 3183 1 1154
2 3184 1 1155
2 3185 1 1155
2 3186 1 1156
2 3187 1 1156
2 3188 1 1161
2 3189 1 1161
2 3190 1 1164
2 3191 1 1164
2 3192 1 1165
2 3193 1 1165
2 3194 1 1166
2 3195 1 1166
2 3196 1 1167
2 3197 1 1167
2 3198 1 1167
2 3199 1 1168
2 3200 1 1168
2 3201 1 1169
2 3202 1 1169
2 3203 1 1170
2 3204 1 1170
2 3205 1 1173
2 3206 1 1173
2 3207 1 1176
2 3208 1 1176
2 3209 1 1177
2 3210 1 1177
2 3211 1 1181
2 3212 1 1181
2 3213 1 1184
2 3214 1 1184
2 3215 1 1185
2 3216 1 1185
2 3217 1 1189
2 3218 1 1189
2 3219 1 1192
2 3220 1 1192
2 3221 1 1193
2 3222 1 1193
2 3223 1 1197
2 3224 1 1197
2 3225 1 1200
2 3226 1 1200
2 3227 1 1201
2 3228 1 1201
2 3229 1 1205
2 3230 1 1205
2 3231 1 1208
2 3232 1 1208
2 3233 1 1209
2 3234 1 1209
2 3235 1 1213
2 3236 1 1213
2 3237 1 1216
2 3238 1 1216
2 3239 1 1217
2 3240 1 1217
2 3241 1 1221
2 3242 1 1221
2 3243 1 1224
2 3244 1 1224
2 3245 1 1225
2 3246 1 1225
2 3247 1 1229
2 3248 1 1229
2 3249 1 1232
2 3250 1 1232
2 3251 1 1233
2 3252 1 1233
2 3253 1 1237
2 3254 1 1237
2 3255 1 1240
2 3256 1 1240
2 3257 1 1241
2 3258 1 1241
2 3259 1 1245
2 3260 1 1245
2 3261 1 1248
2 3262 1 1248
2 3263 1 1249
2 3264 1 1249
2 3265 1 1253
2 3266 1 1253
2 3267 1 1256
2 3268 1 1256
2 3269 1 1257
2 3270 1 1257
2 3271 1 1261
2 3272 1 1261
2 3273 1 1264
2 3274 1 1264
2 3275 1 1265
2 3276 1 1265
2 3277 1 1269
2 3278 1 1269
2 3279 1 1272
2 3280 1 1272
2 3281 1 1273
2 3282 1 1273
2 3283 1 1277
2 3284 1 1277
2 3285 1 1280
2 3286 1 1280
2 3287 1 1281
2 3288 1 1281
2 3289 1 1287
2 3290 1 1287
2 3291 1 1290
2 3292 1 1290
2 3293 1 1293
2 3294 1 1293
2 3295 1 1299
2 3296 1 1299
2 3297 1 1307
2 3298 1 1307
2 3299 1 1315
2 3300 1 1315
2 3301 1 1323
2 3302 1 1323
2 3303 1 1331
2 3304 1 1331
2 3305 1 1339
2 3306 1 1339
2 3307 1 1347
2 3308 1 1347
2 3309 1 1355
2 3310 1 1355
2 3311 1 1363
2 3312 1 1363
2 3313 1 1371
2 3314 1 1371
2 3315 1 1379
2 3316 1 1379
2 3317 1 1387
2 3318 1 1387
2 3319 1 1391
2 3320 1 1391
2 3321 1 1395
2 3322 1 1395
2 3323 1 1397
2 3324 1 1397
2 3325 1 1398
2 3326 1 1398
2 3327 1 1400
2 3328 1 1400
2 3329 1 1405
2 3330 1 1405
2 3331 1 1414
2 3332 1 1414
2 3333 1 1426
2 3334 1 1426
2 3335 1 1484
2 3336 1 1484
2 3337 1 1485
2 3338 1 1485
2 3339 1 1488
2 3340 1 1488
2 3341 1 1489
2 3342 1 1489
2 3343 1 1492
2 3344 1 1492
2 3345 1 1493
2 3346 1 1493
2 3347 1 1496
2 3348 1 1496
2 3349 1 1497
2 3350 1 1497
2 3351 1 1500
2 3352 1 1500
2 3353 1 1501
2 3354 1 1501
2 3355 1 1504
2 3356 1 1504
2 3357 1 1505
2 3358 1 1505
2 3359 1 1508
2 3360 1 1508
2 3361 1 1509
2 3362 1 1509
2 3363 1 1512
2 3364 1 1512
2 3365 1 1513
2 3366 1 1513
2 3367 1 1516
2 3368 1 1516
2 3369 1 1517
2 3370 1 1517
2 3371 1 1520
2 3372 1 1520
2 3373 1 1521
2 3374 1 1521
2 3375 1 1524
2 3376 1 1524
2 3377 1 1525
2 3378 1 1525
2 3379 1 1528
2 3380 1 1528
2 3381 1 1529
2 3382 1 1529
2 3383 1 1532
2 3384 1 1532
2 3385 1 1533
2 3386 1 1533
2 3387 1 1536
2 3388 1 1536
2 3389 1 1536
2 3390 1 1537
2 3391 1 1537
2 3392 1 1537
2 3393 1 1540
2 3394 1 1540
2 3395 1 1540
2 3396 1 1541
2 3397 1 1541
2 3398 1 1551
2 3399 1 1551
2 3400 1 1551
2 3401 1 1552
2 3402 1 1552
2 3403 1 1554
2 3404 1 1554
2 3405 1 1559
2 3406 1 1559
2 3407 1 1565
2 3408 1 1565
2 3409 1 1565
2 3410 1 1566
2 3411 1 1566
2 3412 1 1568
2 3413 1 1568
2 3414 1 1573
2 3415 1 1573
2 3416 1 1573
2 3417 1 1574
2 3418 1 1574
2 3419 1 1576
2 3420 1 1576
2 3421 1 1581
2 3422 1 1581
2 3423 1 1581
2 3424 1 1582
2 3425 1 1582
2 3426 1 1584
2 3427 1 1584
2 3428 1 1589
2 3429 1 1589
2 3430 1 1589
2 3431 1 1590
2 3432 1 1590
2 3433 1 1592
2 3434 1 1592
2 3435 1 1597
2 3436 1 1597
2 3437 1 1597
2 3438 1 1598
2 3439 1 1598
2 3440 1 1600
2 3441 1 1600
2 3442 1 1605
2 3443 1 1605
2 3444 1 1605
2 3445 1 1606
2 3446 1 1606
2 3447 1 1608
2 3448 1 1608
2 3449 1 1613
2 3450 1 1613
2 3451 1 1613
2 3452 1 1614
2 3453 1 1614
2 3454 1 1616
2 3455 1 1616
2 3456 1 1621
2 3457 1 1621
2 3458 1 1621
2 3459 1 1622
2 3460 1 1622
2 3461 1 1624
2 3462 1 1624
2 3463 1 1629
2 3464 1 1629
2 3465 1 1629
2 3466 1 1630
2 3467 1 1630
2 3468 1 1632
2 3469 1 1632
2 3470 1 1637
2 3471 1 1637
2 3472 1 1637
2 3473 1 1638
2 3474 1 1638
2 3475 1 1640
2 3476 1 1640
2 3477 1 1645
2 3478 1 1645
2 3479 1 1645
2 3480 1 1646
2 3481 1 1646
2 3482 1 1648
2 3483 1 1648
2 3484 1 1653
2 3485 1 1653
2 3486 1 1653
2 3487 1 1654
2 3488 1 1654
2 3489 1 1656
2 3490 1 1656
2 3491 1 1659
2 3492 1 1659
2 3493 1 1662
2 3494 1 1662
2 3495 1 1663
2 3496 1 1663
2 3497 1 1664
2 3498 1 1664
2 3499 1 1667
2 3500 1 1667
2 3501 1 1670
2 3502 1 1670
2 3503 1 1671
2 3504 1 1671
2 3505 1 1675
2 3506 1 1675
2 3507 1 1678
2 3508 1 1678
2 3509 1 1679
2 3510 1 1679
2 3511 1 1683
2 3512 1 1683
2 3513 1 1686
2 3514 1 1686
2 3515 1 1687
2 3516 1 1687
2 3517 1 1691
2 3518 1 1691
2 3519 1 1694
2 3520 1 1694
2 3521 1 1695
2 3522 1 1695
2 3523 1 1699
2 3524 1 1699
2 3525 1 1702
2 3526 1 1702
2 3527 1 1703
2 3528 1 1703
2 3529 1 1707
2 3530 1 1707
2 3531 1 1710
2 3532 1 1710
2 3533 1 1711
2 3534 1 1711
2 3535 1 1715
2 3536 1 1715
2 3537 1 1718
2 3538 1 1718
2 3539 1 1719
2 3540 1 1719
2 3541 1 1723
2 3542 1 1723
2 3543 1 1726
2 3544 1 1726
2 3545 1 1727
2 3546 1 1727
2 3547 1 1731
2 3548 1 1731
2 3549 1 1734
2 3550 1 1734
2 3551 1 1735
2 3552 1 1735
2 3553 1 1739
2 3554 1 1739
2 3555 1 1742
2 3556 1 1742
2 3557 1 1743
2 3558 1 1743
2 3559 1 1747
2 3560 1 1747
2 3561 1 1750
2 3562 1 1750
2 3563 1 1751
2 3564 1 1751
2 3565 1 1755
2 3566 1 1755
2 3567 1 1758
2 3568 1 1758
2 3569 1 1759
2 3570 1 1759
2 3571 1 1763
2 3572 1 1763
2 3573 1 1766
2 3574 1 1766
2 3575 1 1767
2 3576 1 1767
2 3577 1 1771
2 3578 1 1771
2 3579 1 1774
2 3580 1 1774
2 3581 1 1775
2 3582 1 1775
2 3583 1 1781
2 3584 1 1781
2 3585 1 1784
2 3586 1 1784
2 3587 1 1786
2 3588 1 1786
2 3589 1 1793
2 3590 1 1793
2 3591 1 1799
2 3592 1 1799
2 3593 1 1807
2 3594 1 1807
2 3595 1 1815
2 3596 1 1815
2 3597 1 1823
2 3598 1 1823
2 3599 1 1831
2 3600 1 1831
2 3601 1 1839
2 3602 1 1839
2 3603 1 1847
2 3604 1 1847
2 3605 1 1855
2 3606 1 1855
2 3607 1 1863
2 3608 1 1863
2 3609 1 1871
2 3610 1 1871
2 3611 1 1879
2 3612 1 1879
2 3613 1 1883
2 3614 1 1883
2 3615 1 1897
2 3616 1 1897
2 3617 1 1909
2 3618 1 1909
0 33 5 1 1 2102
0 34 5 1 1 2104
0 35 5 1 1 2106
0 36 5 1 1 2108
0 37 5 1 1 2110
0 38 5 1 1 2112
0 39 5 1 1 2114
0 40 5 1 1 2116
0 41 5 1 1 2118
0 42 5 1 1 2120
0 43 5 1 1 2122
0 44 5 1 1 2124
0 45 5 1 1 2126
0 46 5 1 1 2128
0 47 5 1 1 2130
0 48 5 1 1 2132
0 49 7 2 2 2029 2094
0 50 5 1 1 2134
0 51 7 2 2 2021 2086
0 52 5 2 1 2136
0 53 7 2 2 2012 2095
0 54 5 1 1 2140
0 55 7 2 2 2030 2078
0 56 5 1 1 2142
0 57 7 1 2 2141 2143
0 58 5 2 1 57
0 59 7 1 2 54 56
0 60 5 1 1 59
0 61 7 2 2 2144 60
0 62 5 1 1 2146
0 63 7 1 2 2137 2147
0 64 5 2 1 63
0 65 7 2 2 2145 2148
0 66 5 1 1 2150
0 67 7 2 2 2022 2096
0 68 5 1 1 2152
0 69 7 2 2 2031 2087
0 70 5 1 1 2154
0 71 7 1 2 68 2155
0 72 5 1 1 71
0 73 7 1 2 2153 70
0 74 5 1 1 73
0 75 7 2 2 72 74
0 76 5 1 1 2156
0 77 7 1 2 66 76
0 78 5 3 1 77
0 79 7 1 2 2138 2158
0 80 5 1 1 79
0 81 7 1 2 2135 80
0 82 5 2 1 81
0 83 7 2 2 2004 2097
0 84 5 1 1 2163
0 85 7 2 2 2032 2070
0 86 5 1 1 2165
0 87 7 1 2 2164 2166
0 88 5 2 1 87
0 89 7 2 2 2023 2079
0 90 5 1 1 2169
0 91 7 1 2 84 86
0 92 5 1 1 91
0 93 7 2 2 2167 92
0 94 5 1 1 2171
0 95 7 1 2 2170 2172
0 96 5 2 1 95
0 97 7 2 2 2168 2173
0 98 5 1 1 2175
0 99 7 1 2 2139 62
0 100 5 1 1 99
0 101 7 2 2 2149 100
0 102 5 1 1 2177
0 103 7 1 2 98 2178
0 104 5 2 1 103
0 105 7 2 2 2013 2088
0 106 5 1 1 2181
0 107 7 1 2 90 94
0 108 5 1 1 107
0 109 7 2 2 2174 108
0 110 5 1 1 2183
0 111 7 1 2 2182 2184
0 112 5 2 1 111
0 113 7 2 2 1995 2098
0 114 5 1 1 2187
0 115 7 2 2 2033 2062
0 116 5 1 1 2189
0 117 7 1 2 2188 2190
0 118 5 2 1 117
0 119 7 2 2 2024 2071
0 120 5 1 1 2193
0 121 7 1 2 114 116
0 122 5 1 1 121
0 123 7 2 2 2191 122
0 124 5 1 1 2195
0 125 7 1 2 2194 2196
0 126 5 2 1 125
0 127 7 2 2 2192 2197
0 128 5 1 1 2199
0 129 7 1 2 106 110
0 130 5 1 1 129
0 131 7 2 2 2185 130
0 132 5 1 1 2201
0 133 7 1 2 128 2202
0 134 5 2 1 133
0 135 7 2 2 2186 2203
0 136 5 1 1 2205
0 137 7 1 2 2176 102
0 138 5 1 1 137
0 139 7 2 2 2179 138
0 140 5 1 1 2207
0 141 7 1 2 136 2208
0 142 5 2 1 141
0 143 7 2 2 2180 2209
0 144 5 1 1 2211
0 145 7 1 2 2151 2157
0 146 5 1 1 145
0 147 7 2 2 2159 146
0 148 5 1 1 2213
0 149 7 1 2 144 2214
0 150 5 2 1 149
0 151 7 2 2 2005 2089
0 152 5 1 1 2217
0 153 7 1 2 120 124
0 154 5 1 1 153
0 155 7 2 2 2198 154
0 156 5 1 1 2219
0 157 7 1 2 2218 2220
0 158 5 2 1 157
0 159 7 2 2 2014 2080
0 160 5 1 1 2223
0 161 7 1 2 152 156
0 162 5 1 1 161
0 163 7 2 2 2221 162
0 164 5 1 1 2225
0 165 7 1 2 2224 2226
0 166 5 2 1 165
0 167 7 2 2 2222 2227
0 168 5 1 1 2229
0 169 7 1 2 2200 132
0 170 5 1 1 169
0 171 7 2 2 2204 170
0 172 5 1 1 2231
0 173 7 1 2 168 2232
0 174 5 2 1 173
0 175 7 2 2 1987 2099
0 176 5 1 1 2235
0 177 7 2 2 2034 2037
0 178 5 1 1 2237
0 179 7 2 2 2025 2045
0 180 5 1 1 2239
0 181 7 2 2 2238 2240
0 182 5 2 1 2241
0 183 7 2 2 2053 2242
0 184 5 2 1 2245
0 185 7 1 2 2236 2246
0 186 5 2 1 185
0 187 7 2 2 2035 2054
0 188 5 1 1 2251
0 189 7 1 2 176 2247
0 190 5 1 1 189
0 191 7 2 2 2249 190
0 192 5 1 1 2253
0 193 7 1 2 2252 2254
0 194 5 2 1 193
0 195 7 2 2 2250 2255
0 196 5 1 1 2257
0 197 7 1 2 160 164
0 198 5 1 1 197
0 199 7 2 2 2228 198
0 200 5 1 1 2259
0 201 7 1 2 196 2260
0 202 5 2 1 201
0 203 7 2 2 2015 2072
0 204 5 1 1 2263
0 205 7 1 2 188 192
0 206 5 1 1 205
0 207 7 2 2 2256 206
0 208 5 1 1 2265
0 209 7 1 2 2264 2266
0 210 5 2 1 209
0 211 7 2 2 2026 2063
0 212 5 1 1 2269
0 213 7 1 2 204 208
0 214 5 1 1 213
0 215 7 2 2 2267 214
0 216 5 1 1 2271
0 217 7 1 2 2270 2272
0 218 5 2 1 217
0 219 7 2 2 2268 2273
0 220 5 1 1 2275
0 221 7 1 2 2258 200
0 222 5 1 1 221
0 223 7 2 2 2261 222
0 224 5 1 1 2277
0 225 7 1 2 220 2278
0 226 5 2 1 225
0 227 7 2 2 2262 2279
0 228 5 1 1 2281
0 229 7 1 2 2230 172
0 230 5 1 1 229
0 231 7 2 2 2233 230
0 232 5 1 1 2283
0 233 7 1 2 228 2284
0 234 5 2 1 233
0 235 7 2 2 2234 2285
0 236 5 1 1 2287
0 237 7 1 2 2206 140
0 238 5 1 1 237
0 239 7 2 2 2210 238
0 240 5 1 1 2289
0 241 7 1 2 236 2290
0 242 5 2 1 241
0 243 7 2 2 1996 2090
0 244 5 1 1 2293
0 245 7 2 2 2006 2081
0 246 5 1 1 2295
0 247 7 1 2 2294 2296
0 248 5 2 1 247
0 249 7 1 2 212 216
0 250 5 1 1 249
0 251 7 2 2 2274 250
0 252 5 1 1 2299
0 253 7 1 2 244 246
0 254 5 1 1 253
0 255 7 2 2 2297 254
0 256 5 1 1 2301
0 257 7 1 2 2300 2302
0 258 5 2 1 257
0 259 7 2 2 2298 2303
0 260 5 1 1 2305
0 261 7 1 2 2276 224
0 262 5 1 1 261
0 263 7 2 2 2280 262
0 264 5 1 1 2307
0 265 7 1 2 260 2308
0 266 5 2 1 265
0 267 7 2 2 2016 2064
0 268 5 1 1 2311
0 269 7 2 2 1988 2091
0 270 5 1 1 2313
0 271 7 1 2 2312 2314
0 272 5 2 1 271
0 273 7 2 2 1979 2100
0 274 5 1 1 2317
0 275 7 2 2 2007 2073
0 276 5 1 1 2319
0 277 7 1 2 2027 2055
0 278 5 1 1 277
0 279 7 1 2 2243 278
0 280 5 1 1 279
0 281 7 2 2 2248 280
0 282 5 1 1 2321
0 283 7 1 2 2320 2322
0 284 5 2 1 283
0 285 7 1 2 276 282
0 286 5 1 1 285
0 287 7 2 2 2323 286
0 288 5 1 1 2325
0 289 7 1 2 2318 2326
0 290 5 2 1 289
0 291 7 1 2 274 288
0 292 5 1 1 291
0 293 7 2 2 2327 292
0 294 5 1 1 2329
0 295 7 1 2 268 270
0 296 5 1 1 295
0 297 7 2 2 2315 296
0 298 5 1 1 2331
0 299 7 1 2 2330 2332
0 300 5 2 1 299
0 301 7 2 2 2316 2333
0 302 5 1 1 2335
0 303 7 1 2 252 256
0 304 5 1 1 303
0 305 7 2 2 2304 304
0 306 5 1 1 2337
0 307 7 1 2 302 2338
0 308 5 2 1 307
0 309 7 2 2 2036 2046
0 310 5 1 1 2341
0 311 7 2 2 1997 2082
0 312 5 1 1 2343
0 313 7 1 2 2342 2344
0 314 5 2 1 313
0 315 7 1 2 294 298
0 316 5 1 1 315
0 317 7 2 2 2334 316
0 318 5 1 1 2347
0 319 7 1 2 310 312
0 320 5 1 1 319
0 321 7 2 2 2345 320
0 322 5 1 1 2349
0 323 7 1 2 2348 2350
0 324 5 2 1 323
0 325 7 2 2 2346 2351
0 326 5 1 1 2353
0 327 7 1 2 2336 306
0 328 5 1 1 327
0 329 7 2 2 2339 328
0 330 5 1 1 2355
0 331 7 1 2 326 2356
0 332 5 2 1 331
0 333 7 2 2 2340 2357
0 334 5 1 1 2359
0 335 7 1 2 2306 264
0 336 5 1 1 335
0 337 7 2 2 2309 336
0 338 5 1 1 2361
0 339 7 1 2 334 2362
0 340 5 2 1 339
0 341 7 2 2 2310 2363
0 342 5 1 1 2365
0 343 7 1 2 2282 232
0 344 5 1 1 343
0 345 7 2 2 2286 344
0 346 5 1 1 2367
0 347 7 1 2 342 2368
0 348 5 2 1 347
0 349 7 2 2 2324 2328
0 350 5 1 1 2371
0 351 7 1 2 2354 330
0 352 5 1 1 351
0 353 7 2 2 2358 352
0 354 5 1 1 2373
0 355 7 1 2 350 2374
0 356 5 2 1 355
0 357 7 2 2 2017 2056
0 358 5 1 1 2377
0 359 7 2 2 2008 2065
0 360 5 1 1 2379
0 361 7 1 2 2378 2380
0 362 5 2 1 361
0 363 7 2 2 1980 2092
0 364 5 1 1 2383
0 365 7 1 2 358 360
0 366 5 1 1 365
0 367 7 2 2 2381 366
0 368 5 1 1 2385
0 369 7 1 2 2384 2386
0 370 5 2 1 369
0 371 7 2 2 2382 2387
0 372 5 1 1 2389
0 373 7 2 2 1989 2083
0 374 5 1 1 2391
0 375 7 2 2 32 2101
0 376 5 1 1 2393
0 377 7 1 2 2392 2394
0 378 5 2 1 377
0 379 7 2 2 1998 2074
0 380 5 1 1 2397
0 381 7 2 2 2009 2047
0 382 5 1 1 2399
0 383 7 2 2 1972 2066
0 384 5 1 1 2401
0 385 7 2 2 1990 2048
0 386 5 1 1 2403
0 387 7 2 2 2402 2404
0 388 5 2 1 2405
0 389 7 2 2 1999 2406
0 390 5 2 1 2409
0 391 7 2 2 2400 2410
0 392 5 2 1 2413
0 393 7 2 2 2018 2414
0 394 5 2 1 2417
0 395 7 1 2 2398 2418
0 396 5 2 1 395
0 397 7 1 2 380 2419
0 398 5 1 1 397
0 399 7 2 2 2421 398
0 400 5 1 1 2423
0 401 7 1 2 178 180
0 402 5 1 1 401
0 403 7 2 2 2244 402
0 404 5 1 1 2425
0 405 7 1 2 2424 2426
0 406 5 2 1 405
0 407 7 1 2 400 404
0 408 5 1 1 407
0 409 7 2 2 2427 408
0 410 5 1 1 2429
0 411 7 1 2 374 376
0 412 5 1 1 411
0 413 7 2 2 2395 412
0 414 5 1 1 2431
0 415 7 1 2 2430 2432
0 416 5 2 1 415
0 417 7 2 2 2396 2433
0 418 5 1 1 2435
0 419 7 1 2 372 418
0 420 5 2 1 419
0 421 7 2 2 2422 2428
0 422 5 1 1 2439
0 423 7 1 2 2390 2436
0 424 5 1 1 423
0 425 7 2 2 2437 424
0 426 5 1 1 2441
0 427 7 1 2 422 2442
0 428 5 2 1 427
0 429 7 2 2 2438 2443
0 430 5 1 1 2445
0 431 7 1 2 2372 354
0 432 5 1 1 431
0 433 7 2 2 2375 432
0 434 5 1 1 2447
0 435 7 1 2 430 2448
0 436 5 2 1 435
0 437 7 2 2 2376 2449
0 438 5 1 1 2451
0 439 7 1 2 2360 338
0 440 5 1 1 439
0 441 7 2 2 2364 440
0 442 5 1 1 2453
0 443 7 1 2 438 2454
0 444 5 2 1 443
0 445 7 1 2 318 322
0 446 5 1 1 445
0 447 7 2 2 2352 446
0 448 5 1 1 2457
0 449 7 1 2 2440 426
0 450 5 1 1 449
0 451 7 2 2 2444 450
0 452 5 1 1 2459
0 453 7 1 2 2458 2460
0 454 5 2 1 453
0 455 7 1 2 364 368
0 456 5 1 1 455
0 457 7 2 2 2388 456
0 458 5 1 1 2463
0 459 7 1 2 410 414
0 460 5 1 1 459
0 461 7 2 2 2434 460
0 462 5 1 1 2465
0 463 7 1 2 2464 2466
0 464 5 2 1 463
0 465 7 2 2 2000 2067
0 466 5 1 1 2469
0 467 7 2 2 1991 2075
0 468 5 1 1 2471
0 469 7 1 2 2470 2472
0 470 5 2 1 469
0 471 7 2 2 1981 2084
0 472 5 1 1 2475
0 473 7 1 2 466 468
0 474 5 1 1 473
0 475 7 2 2 2473 474
0 476 5 1 1 2477
0 477 7 1 2 2476 2478
0 478 5 2 1 477
0 479 7 2 2 2474 2479
0 480 5 1 1 2481
0 481 7 1 2 458 462
0 482 5 1 1 481
0 483 7 2 2 2467 482
0 484 5 1 1 2483
0 485 7 1 2 480 2484
0 486 5 2 1 485
0 487 7 2 2 2468 2485
0 488 5 1 1 2487
0 489 7 1 2 448 452
0 490 5 1 1 489
0 491 7 2 2 2461 490
0 492 5 1 1 2489
0 493 7 1 2 488 2490
0 494 5 2 1 493
0 495 7 2 2 2462 2491
0 496 5 1 1 2493
0 497 7 1 2 2446 434
0 498 5 1 1 497
0 499 7 2 2 2450 498
0 500 5 1 1 2495
0 501 7 1 2 496 2496
0 502 5 2 1 501
0 503 7 2 2 1973 2093
0 504 5 1 1 2499
0 505 7 1 2 472 476
0 506 5 1 1 505
0 507 7 2 2 2480 506
0 508 5 1 1 2501
0 509 7 1 2 2500 2502
0 510 5 2 1 509
0 511 7 2 2 2028 2038
0 512 5 1 1 2505
0 513 7 2 2 2010 2057
0 514 5 1 1 2507
0 515 7 1 2 2019 2049
0 516 5 1 1 515
0 517 7 1 2 2415 516
0 518 5 1 1 517
0 519 7 2 2 2420 518
0 520 5 1 1 2509
0 521 7 1 2 2508 2510
0 522 5 2 1 521
0 523 7 1 2 514 520
0 524 5 1 1 523
0 525 7 2 2 2511 524
0 526 5 1 1 2513
0 527 7 1 2 2506 2514
0 528 5 2 1 527
0 529 7 1 2 512 526
0 530 5 1 1 529
0 531 7 2 2 2515 530
0 532 5 1 1 2517
0 533 7 1 2 504 508
0 534 5 1 1 533
0 535 7 2 2 2503 534
0 536 5 1 1 2519
0 537 7 1 2 2518 2520
0 538 5 2 1 537
0 539 7 2 2 2504 2521
0 540 5 1 1 2523
0 541 7 1 2 2482 484
0 542 5 1 1 541
0 543 7 2 2 2486 542
0 544 5 1 1 2525
0 545 7 1 2 540 2526
0 546 5 2 1 545
0 547 7 2 2 2512 2516
0 548 5 1 1 2529
0 549 7 1 2 2524 544
0 550 5 1 1 549
0 551 7 2 2 2527 550
0 552 5 1 1 2531
0 553 7 1 2 548 2532
0 554 5 2 1 553
0 555 7 2 2 2528 2533
0 556 5 1 1 2535
0 557 7 1 2 2488 492
0 558 5 1 1 557
0 559 7 2 2 2492 558
0 560 5 1 1 2537
0 561 7 1 2 556 2538
0 562 5 2 1 561
0 563 7 2 2 2001 2058
0 564 5 1 1 2541
0 565 7 1 2 382 2411
0 566 5 1 1 565
0 567 7 2 2 2416 566
0 568 5 1 1 2543
0 569 7 1 2 2542 2544
0 570 5 2 1 569
0 571 7 2 2 2020 2039
0 572 5 1 1 2547
0 573 7 1 2 564 568
0 574 5 1 1 573
0 575 7 2 2 2545 574
0 576 5 1 1 2549
0 577 7 1 2 2548 2550
0 578 5 2 1 577
0 579 7 2 2 2546 2551
0 580 5 1 1 2553
0 581 7 1 2 532 536
0 582 5 1 1 581
0 583 7 2 2 2522 582
0 584 5 1 1 2555
0 585 7 1 2 580 2556
0 586 5 2 1 585
0 587 7 2 2 1992 2068
0 588 5 1 1 2559
0 589 7 2 2 1974 2085
0 590 5 1 1 2561
0 591 7 1 2 2560 2562
0 592 5 2 1 591
0 593 7 1 2 572 576
0 594 5 1 1 593
0 595 7 2 2 2552 594
0 596 5 1 1 2565
0 597 7 1 2 588 590
0 598 5 1 1 597
0 599 7 2 2 2563 598
0 600 5 1 1 2567
0 601 7 1 2 2566 2568
0 602 5 2 1 601
0 603 7 2 2 2564 2569
0 604 5 1 1 2571
0 605 7 1 2 2554 584
0 606 5 1 1 605
0 607 7 2 2 2557 606
0 608 5 1 1 2573
0 609 7 1 2 604 2574
0 610 5 2 1 609
0 611 7 2 2 2558 2575
0 612 5 1 1 2577
0 613 7 1 2 2530 552
0 614 5 1 1 613
0 615 7 2 2 2534 614
0 616 5 1 1 2579
0 617 7 1 2 612 2580
0 618 5 2 1 617
0 619 7 2 2 1982 2076
0 620 5 1 1 2583
0 621 7 1 2 596 600
0 622 5 1 1 621
0 623 7 2 2 2570 622
0 624 5 1 1 2585
0 625 7 1 2 2584 2586
0 626 5 2 1 625
0 627 7 2 2 1993 2059
0 628 5 1 1 2589
0 629 7 1 2 2002 2050
0 630 5 1 1 629
0 631 7 1 2 2407 630
0 632 5 1 1 631
0 633 7 2 2 2412 632
0 634 5 1 1 2591
0 635 7 1 2 2590 2592
0 636 5 2 1 635
0 637 7 2 2 2011 2040
0 638 5 1 1 2595
0 639 7 1 2 628 634
0 640 5 1 1 639
0 641 7 2 2 2593 640
0 642 5 1 1 2597
0 643 7 1 2 2596 2598
0 644 5 2 1 643
0 645 7 2 2 2594 2599
0 646 5 1 1 2601
0 647 7 1 2 620 624
0 648 5 1 1 647
0 649 7 2 2 2587 648
0 650 5 1 1 2603
0 651 7 1 2 646 2604
0 652 5 2 1 651
0 653 7 2 2 2588 2605
0 654 5 1 1 2607
0 655 7 1 2 2572 608
0 656 5 1 1 655
0 657 7 2 2 2576 656
0 658 5 1 1 2609
0 659 7 1 2 654 2610
0 660 5 2 1 659
0 661 7 2 2 1975 2077
0 662 5 1 1 2613
0 663 7 2 2 1983 2069
0 664 5 1 1 2615
0 665 7 1 2 2614 2616
0 666 5 2 1 665
0 667 7 1 2 638 642
0 668 5 1 1 667
0 669 7 2 2 2600 668
0 670 5 1 1 2619
0 671 7 1 2 662 664
0 672 5 1 1 671
0 673 7 2 2 2617 672
0 674 5 1 1 2621
0 675 7 1 2 2620 2622
0 676 5 2 1 675
0 677 7 2 2 2618 2623
0 678 5 1 1 2625
0 679 7 1 2 2602 650
0 680 5 1 1 679
0 681 7 2 2 2606 680
0 682 5 1 1 2627
0 683 7 1 2 678 2628
0 684 5 2 1 683
0 685 7 1 2 670 674
0 686 5 1 1 685
0 687 7 2 2 2624 686
0 688 5 1 1 2631
0 689 7 2 2 1984 2060
0 690 5 1 1 2633
0 691 7 2 2 2003 2041
0 692 5 1 1 2635
0 693 7 2 2 2634 2636
0 694 5 1 1 2637
0 695 7 2 2 1985 2051
0 696 5 1 1 2639
0 697 7 2 2 1976 2061
0 698 5 1 1 2641
0 699 7 2 2 2640 2642
0 700 5 2 1 2643
0 701 7 3 2 694 2645
0 702 5 1 1 2647
0 703 7 1 2 2632 702
0 704 5 2 1 703
0 705 7 1 2 384 386
0 706 5 1 1 705
0 707 7 2 2 2408 706
0 708 5 1 1 2652
0 709 7 1 2 690 692
0 710 5 1 1 709
0 711 7 1 2 2648 710
0 712 5 1 1 711
0 713 7 1 2 2638 2644
0 714 5 1 1 713
0 715 7 2 2 712 714
0 716 5 1 1 2654
0 717 7 1 2 2653 716
0 718 5 2 1 717
0 719 7 2 2 1994 2042
0 720 5 1 1 2658
0 721 7 1 2 696 698
0 722 5 1 1 721
0 723 7 2 2 2646 722
0 724 5 1 1 2660
0 725 7 1 2 2659 2661
0 726 5 2 1 725
0 727 7 1 2 720 724
0 728 5 1 1 727
0 729 7 2 2 2662 728
0 730 5 1 1 2664
0 731 7 2 2 1977 2052
0 732 5 1 1 2666
0 733 7 2 2 1986 2043
0 734 5 1 1 2668
0 735 7 2 2 2667 2669
0 736 5 2 1 2670
0 737 7 1 2 2665 2671
0 738 5 2 1 737
0 739 7 2 2 2663 2674
0 740 5 1 1 2676
0 741 7 1 2 708 2655
0 742 5 1 1 741
0 743 7 2 2 2656 742
0 744 5 1 1 2678
0 745 7 1 2 740 2679
0 746 5 2 1 745
0 747 7 2 2 2657 2680
0 748 5 1 1 2682
0 749 7 1 2 688 2649
0 750 5 1 1 749
0 751 7 2 2 2650 750
0 752 5 1 1 2684
0 753 7 1 2 748 2685
0 754 5 2 1 753
0 755 7 2 2 2651 2686
0 756 5 1 1 2688
0 757 7 1 2 2626 682
0 758 5 1 1 757
0 759 7 2 2 2629 758
0 760 5 1 1 2690
0 761 7 1 2 756 2691
0 762 5 2 1 761
0 763 7 2 2 2630 2692
0 764 5 1 1 2694
0 765 7 1 2 2608 658
0 766 5 1 1 765
0 767 7 2 2 2611 766
0 768 5 1 1 2696
0 769 7 1 2 764 2697
0 770 5 2 1 769
0 771 7 2 2 2612 2698
0 772 5 1 1 2700
0 773 7 1 2 2578 616
0 774 5 1 1 773
0 775 7 2 2 2581 774
0 776 5 1 1 2702
0 777 7 1 2 772 2703
0 778 5 2 1 777
0 779 7 2 2 2582 2704
0 780 5 1 1 2706
0 781 7 1 2 2536 560
0 782 5 1 1 781
0 783 7 2 2 2539 782
0 784 5 1 1 2708
0 785 7 1 2 780 2709
0 786 5 2 1 785
0 787 7 2 2 2540 2710
0 788 5 1 1 2712
0 789 7 1 2 2494 500
0 790 5 1 1 789
0 791 7 2 2 2497 790
0 792 5 1 1 2714
0 793 7 1 2 788 2715
0 794 5 2 1 793
0 795 7 2 2 2498 2716
0 796 5 1 1 2718
0 797 7 1 2 2452 442
0 798 5 1 1 797
0 799 7 2 2 2455 798
0 800 5 1 1 2720
0 801 7 1 2 796 2721
0 802 5 2 1 801
0 803 7 2 2 2456 2722
0 804 5 1 1 2724
0 805 7 1 2 2366 346
0 806 5 1 1 805
0 807 7 2 2 2369 806
0 808 5 1 1 2726
0 809 7 1 2 804 2727
0 810 5 2 1 809
0 811 7 2 2 2370 2728
0 812 5 1 1 2730
0 813 7 1 2 2288 240
0 814 5 1 1 813
0 815 7 2 2 2291 814
0 816 5 1 1 2732
0 817 7 1 2 812 2733
0 818 5 2 1 817
0 819 7 2 2 2292 2734
0 820 5 1 1 2736
0 821 7 1 2 2212 148
0 822 5 1 1 821
0 823 7 2 2 2215 822
0 824 5 1 1 2738
0 825 7 1 2 820 2739
0 826 5 2 1 825
0 827 7 2 2 2216 2740
0 828 5 1 1 2742
0 829 7 1 2 50 2160
0 830 5 1 1 829
0 831 7 2 2 2161 830
0 832 5 1 1 2744
0 833 7 1 2 828 2745
0 834 5 2 1 833
0 835 7 4 2 2162 2746
0 836 5 3 1 2748
0 837 7 3 2 48 2752
0 838 5 3 1 2755
0 839 7 3 2 2133 2749
0 840 5 3 1 2761
0 841 7 1 2 2743 832
0 842 5 1 1 841
0 843 7 4 2 2747 842
0 844 5 3 1 2767
0 845 7 1 2 2131 2771
0 846 5 3 1 845
0 847 7 1 2 47 2768
0 848 5 3 1 847
0 849 7 1 2 2737 824
0 850 5 1 1 849
0 851 7 4 2 2741 850
0 852 5 3 1 2780
0 853 7 1 2 2129 2784
0 854 5 3 1 853
0 855 7 1 2 46 2781
0 856 5 3 1 855
0 857 7 1 2 2731 816
0 858 5 1 1 857
0 859 7 4 2 2735 858
0 860 5 3 1 2793
0 861 7 1 2 2127 2797
0 862 5 3 1 861
0 863 7 1 2 45 2794
0 864 5 3 1 863
0 865 7 1 2 2725 808
0 866 5 1 1 865
0 867 7 4 2 2729 866
0 868 5 3 1 2806
0 869 7 1 2 2125 2810
0 870 5 3 1 869
0 871 7 1 2 44 2807
0 872 5 3 1 871
0 873 7 1 2 2719 800
0 874 5 1 1 873
0 875 7 4 2 2723 874
0 876 5 3 1 2819
0 877 7 1 2 2123 2823
0 878 5 3 1 877
0 879 7 1 2 43 2820
0 880 5 3 1 879
0 881 7 1 2 2713 792
0 882 5 1 1 881
0 883 7 4 2 2717 882
0 884 5 3 1 2832
0 885 7 1 2 2121 2836
0 886 5 3 1 885
0 887 7 1 2 42 2833
0 888 5 3 1 887
0 889 7 1 2 2707 784
0 890 5 1 1 889
0 891 7 4 2 2711 890
0 892 5 3 1 2845
0 893 7 1 2 2119 2849
0 894 5 3 1 893
0 895 7 1 2 41 2846
0 896 5 3 1 895
0 897 7 1 2 2701 776
0 898 5 1 1 897
0 899 7 4 2 2705 898
0 900 5 3 1 2858
0 901 7 1 2 2117 2862
0 902 5 3 1 901
0 903 7 1 2 40 2859
0 904 5 3 1 903
0 905 7 1 2 2695 768
0 906 5 1 1 905
0 907 7 4 2 2699 906
0 908 5 3 1 2871
0 909 7 1 2 2115 2875
0 910 5 3 1 909
0 911 7 1 2 39 2872
0 912 5 3 1 911
0 913 7 1 2 2689 760
0 914 5 1 1 913
0 915 7 4 2 2693 914
0 916 5 3 1 2884
0 917 7 1 2 2113 2888
0 918 5 3 1 917
0 919 7 1 2 38 2885
0 920 5 3 1 919
0 921 7 1 2 2683 752
0 922 5 1 1 921
0 923 7 4 2 2687 922
0 924 5 3 1 2897
0 925 7 1 2 2111 2901
0 926 5 3 1 925
0 927 7 1 2 37 2898
0 928 5 3 1 927
0 929 7 1 2 2677 744
0 930 5 1 1 929
0 931 7 4 2 2681 930
0 932 5 3 1 2910
0 933 7 1 2 2109 2914
0 934 5 3 1 933
0 935 7 1 2 36 2911
0 936 5 3 1 935
0 937 7 1 2 730 2672
0 938 5 1 1 937
0 939 7 2 2 2675 938
0 940 5 3 1 2923
0 941 7 1 2 2107 2925
0 942 5 3 1 941
0 943 7 1 2 35 2924
0 944 5 3 1 943
0 945 7 1 2 732 734
0 946 5 1 1 945
0 947 7 4 2 2673 946
0 948 5 3 1 2934
0 949 7 1 2 2105 2938
0 950 5 3 1 949
0 951 7 1 2 34 2935
0 952 5 4 1 951
0 953 7 3 2 1978 2044
0 954 5 2 1 2948
0 955 7 2 2 33 2949
0 956 5 4 1 2953
0 957 7 1 2 2944 2955
0 958 5 1 1 957
0 959 7 2 2 2941 958
0 960 5 2 1 2959
0 961 7 1 2 2931 2961
0 962 5 1 1 961
0 963 7 2 2 2928 962
0 964 5 2 1 2963
0 965 7 1 2 2920 2965
0 966 5 1 1 965
0 967 7 2 2 2917 966
0 968 5 2 1 2967
0 969 7 1 2 2907 2969
0 970 5 1 1 969
0 971 7 2 2 2904 970
0 972 5 2 1 2971
0 973 7 1 2 2894 2973
0 974 5 1 1 973
0 975 7 2 2 2891 974
0 976 5 2 1 2975
0 977 7 1 2 2881 2977
0 978 5 1 1 977
0 979 7 2 2 2878 978
0 980 5 2 1 2979
0 981 7 1 2 2868 2981
0 982 5 1 1 981
0 983 7 2 2 2865 982
0 984 5 2 1 2983
0 985 7 1 2 2855 2985
0 986 5 1 1 985
0 987 7 2 2 2852 986
0 988 5 2 1 2987
0 989 7 1 2 2842 2989
0 990 5 1 1 989
0 991 7 2 2 2839 990
0 992 5 2 1 2991
0 993 7 1 2 2829 2993
0 994 5 1 1 993
0 995 7 2 2 2826 994
0 996 5 2 1 2995
0 997 7 1 2 2816 2997
0 998 5 1 1 997
0 999 7 2 2 2813 998
0 1000 5 2 1 2999
0 1001 7 1 2 2803 3001
0 1002 5 1 1 1001
0 1003 7 2 2 2800 1002
0 1004 5 2 1 3003
0 1005 7 1 2 2790 3005
0 1006 5 1 1 1005
0 1007 7 2 2 2787 1006
0 1008 5 2 1 3007
0 1009 7 1 2 2777 3009
0 1010 5 1 1 1009
0 1011 7 4 2 2774 1010
0 1012 5 2 1 3011
0 1013 7 1 2 2764 3012
0 1014 5 2 1 1013
0 1015 7 2 2 2758 3017
0 1016 5 1 1 3019
0 1017 7 3 2 2775 2778
0 1018 5 2 1 3021
0 1019 7 1 2 3010 3022
0 1020 5 1 1 1019
0 1021 7 1 2 3008 3024
0 1022 5 1 1 1021
0 1023 7 3 2 1020 1022
0 1024 5 2 1 3026
0 1025 7 1 2 1016 3027
0 1026 5 2 1 1025
0 1027 7 3 2 2759 2765
0 1028 5 2 1 3033
0 1029 7 1 2 3015 3034
0 1030 5 1 1 1029
0 1031 7 1 2 3013 3036
0 1032 5 1 1 1031
0 1033 7 2 2 1030 1032
0 1034 5 1 1 3038
0 1035 7 3 2 2788 2791
0 1036 5 2 1 3040
0 1037 7 1 2 3004 3041
0 1038 5 1 1 1037
0 1039 7 1 2 3006 3043
0 1040 5 1 1 1039
0 1041 7 3 2 1038 1040
0 1042 5 2 1 3045
0 1043 7 1 2 3039 3048
0 1044 5 2 1 1043
0 1045 7 3 2 2801 2804
0 1046 5 2 1 3052
0 1047 7 1 2 3000 3053
0 1048 5 1 1 1047
0 1049 7 1 2 3002 3055
0 1050 5 1 1 1049
0 1051 7 3 2 1048 1050
0 1052 5 2 1 3057
0 1053 7 1 2 3028 3060
0 1054 5 2 1 1053
0 1055 7 3 2 2814 2817
0 1056 5 2 1 3064
0 1057 7 1 2 2996 3065
0 1058 5 1 1 1057
0 1059 7 1 2 2998 3067
0 1060 5 1 1 1059
0 1061 7 3 2 1058 1060
0 1062 5 2 1 3069
0 1063 7 1 2 3049 3072
0 1064 5 2 1 1063
0 1065 7 3 2 2827 2830
0 1066 5 2 1 3076
0 1067 7 1 2 2992 3077
0 1068 5 1 1 1067
0 1069 7 1 2 2994 3079
0 1070 5 1 1 1069
0 1071 7 3 2 1068 1070
0 1072 5 2 1 3081
0 1073 7 1 2 3061 3084
0 1074 5 2 1 1073
0 1075 7 3 2 2840 2843
0 1076 5 2 1 3088
0 1077 7 1 2 2988 3089
0 1078 5 1 1 1077
0 1079 7 1 2 2990 3091
0 1080 5 1 1 1079
0 1081 7 3 2 1078 1080
0 1082 5 2 1 3093
0 1083 7 1 2 3073 3096
0 1084 5 2 1 1083
0 1085 7 3 2 2853 2856
0 1086 5 2 1 3100
0 1087 7 1 2 2984 3101
0 1088 5 1 1 1087
0 1089 7 1 2 2986 3103
0 1090 5 1 1 1089
0 1091 7 3 2 1088 1090
0 1092 5 2 1 3105
0 1093 7 1 2 3085 3108
0 1094 5 2 1 1093
0 1095 7 3 2 2866 2869
0 1096 5 2 1 3112
0 1097 7 1 2 2980 3113
0 1098 5 1 1 1097
0 1099 7 1 2 2982 3115
0 1100 5 1 1 1099
0 1101 7 3 2 1098 1100
0 1102 5 2 1 3117
0 1103 7 1 2 3097 3120
0 1104 5 2 1 1103
0 1105 7 3 2 2879 2882
0 1106 5 2 1 3124
0 1107 7 1 2 2976 3125
0 1108 5 1 1 1107
0 1109 7 1 2 2978 3127
0 1110 5 1 1 1109
0 1111 7 3 2 1108 1110
0 1112 5 2 1 3129
0 1113 7 1 2 3109 3132
0 1114 5 2 1 1113
0 1115 7 3 2 2892 2895
0 1116 5 2 1 3136
0 1117 7 1 2 2972 3137
0 1118 5 1 1 1117
0 1119 7 1 2 2974 3139
0 1120 5 1 1 1119
0 1121 7 3 2 1118 1120
0 1122 5 2 1 3141
0 1123 7 1 2 3121 3144
0 1124 5 2 1 1123
0 1125 7 3 2 2905 2908
0 1126 5 2 1 3148
0 1127 7 1 2 2968 3149
0 1128 5 1 1 1127
0 1129 7 1 2 2970 3151
0 1130 5 1 1 1129
0 1131 7 3 2 1128 1130
0 1132 5 2 1 3153
0 1133 7 1 2 3133 3156
0 1134 5 2 1 1133
0 1135 7 3 2 2918 2921
0 1136 5 2 1 3160
0 1137 7 1 2 2964 3161
0 1138 5 1 1 1137
0 1139 7 1 2 2966 3163
0 1140 5 1 1 1139
0 1141 7 3 2 1138 1140
0 1142 5 2 1 3165
0 1143 7 1 2 3145 3168
0 1144 5 2 1 1143
0 1145 7 3 2 2929 2932
0 1146 5 2 1 3172
0 1147 7 1 2 2960 3173
0 1148 5 1 1 1147
0 1149 7 1 2 2962 3175
0 1150 5 1 1 1149
0 1151 7 3 2 1148 1150
0 1152 5 2 1 3177
0 1153 7 1 2 3157 3180
0 1154 5 2 1 1153
0 1155 7 2 2 2942 2945
0 1156 5 2 1 3184
0 1157 7 1 2 2954 3185
0 1158 5 1 1 1157
0 1159 7 1 2 2956 3186
0 1160 5 1 1 1159
0 1161 7 2 2 1158 1160
0 1162 5 1 1 3188
0 1163 7 1 2 3169 1162
0 1164 5 2 1 1163
0 1165 7 2 2 2103 2951
0 1166 5 2 1 3192
0 1167 7 3 2 2957 3194
0 1168 5 2 1 3196
0 1169 7 2 2 3181 3199
0 1170 5 2 1 3201
0 1171 7 1 2 3166 3189
0 1172 5 1 1 1171
0 1173 7 2 2 3190 1172
0 1174 5 1 1 3205
0 1175 7 1 2 3202 3206
0 1176 5 2 1 1175
0 1177 7 2 2 3191 3207
0 1178 5 1 1 3209
0 1179 7 1 2 3154 3178
0 1180 5 1 1 1179
0 1181 7 2 2 3182 1180
0 1182 5 1 1 3211
0 1183 7 1 2 1178 3212
0 1184 5 2 1 1183
0 1185 7 2 2 3183 3213
0 1186 5 1 1 3215
0 1187 7 1 2 3142 3167
0 1188 5 1 1 1187
0 1189 7 2 2 3170 1188
0 1190 5 1 1 3217
0 1191 7 1 2 1186 3218
0 1192 5 2 1 1191
0 1193 7 2 2 3171 3219
0 1194 5 1 1 3221
0 1195 7 1 2 3130 3155
0 1196 5 1 1 1195
0 1197 7 2 2 3158 1196
0 1198 5 1 1 3223
0 1199 7 1 2 1194 3224
0 1200 5 2 1 1199
0 1201 7 2 2 3159 3225
0 1202 5 1 1 3227
0 1203 7 1 2 3118 3143
0 1204 5 1 1 1203
0 1205 7 2 2 3146 1204
0 1206 5 1 1 3229
0 1207 7 1 2 1202 3230
0 1208 5 2 1 1207
0 1209 7 2 2 3147 3231
0 1210 5 1 1 3233
0 1211 7 1 2 3106 3131
0 1212 5 1 1 1211
0 1213 7 2 2 3134 1212
0 1214 5 1 1 3235
0 1215 7 1 2 1210 3236
0 1216 5 2 1 1215
0 1217 7 2 2 3135 3237
0 1218 5 1 1 3239
0 1219 7 1 2 3094 3119
0 1220 5 1 1 1219
0 1221 7 2 2 3122 1220
0 1222 5 1 1 3241
0 1223 7 1 2 1218 3242
0 1224 5 2 1 1223
0 1225 7 2 2 3123 3243
0 1226 5 1 1 3245
0 1227 7 1 2 3082 3107
0 1228 5 1 1 1227
0 1229 7 2 2 3110 1228
0 1230 5 1 1 3247
0 1231 7 1 2 1226 3248
0 1232 5 2 1 1231
0 1233 7 2 2 3111 3249
0 1234 5 1 1 3251
0 1235 7 1 2 3070 3095
0 1236 5 1 1 1235
0 1237 7 2 2 3098 1236
0 1238 5 1 1 3253
0 1239 7 1 2 1234 3254
0 1240 5 2 1 1239
0 1241 7 2 2 3099 3255
0 1242 5 1 1 3257
0 1243 7 1 2 3058 3083
0 1244 5 1 1 1243
0 1245 7 2 2 3086 1244
0 1246 5 1 1 3259
0 1247 7 1 2 1242 3260
0 1248 5 2 1 1247
0 1249 7 2 2 3087 3261
0 1250 5 1 1 3263
0 1251 7 1 2 3046 3071
0 1252 5 1 1 1251
0 1253 7 2 2 3074 1252
0 1254 5 1 1 3265
0 1255 7 1 2 1250 3266
0 1256 5 2 1 1255
0 1257 7 2 2 3075 3267
0 1258 5 1 1 3269
0 1259 7 1 2 3029 3059
0 1260 5 1 1 1259
0 1261 7 2 2 3062 1260
0 1262 5 1 1 3271
0 1263 7 1 2 1258 3272
0 1264 5 2 1 1263
0 1265 7 2 2 3063 3273
0 1266 5 1 1 3275
0 1267 7 1 2 1034 3047
0 1268 5 1 1 1267
0 1269 7 2 2 3050 1268
0 1270 5 1 1 3277
0 1271 7 1 2 1266 3278
0 1272 5 2 1 1271
0 1273 7 2 2 3051 3279
0 1274 5 1 1 3281
0 1275 7 1 2 3020 3030
0 1276 5 1 1 1275
0 1277 7 2 2 3031 1276
0 1278 5 1 1 3283
0 1279 7 1 2 1274 3284
0 1280 5 2 1 1279
0 1281 7 2 2 3032 3285
0 1282 5 1 1 3287
0 1283 7 1 2 2762 3016
0 1284 5 1 1 1283
0 1285 7 1 2 2756 3014
0 1286 5 1 1 1285
0 1287 7 2 2 1284 1286
0 1288 5 1 1 3289
0 1289 7 1 2 1282 1288
0 1290 5 2 1 1289
0 1291 7 1 2 3288 3290
0 1292 5 1 1 1291
0 1293 7 2 2 3291 1292
0 1294 5 1 1 3293
0 1295 7 1 2 2753 1294
0 1296 5 1 1 1295
0 1297 7 1 2 3282 1278
0 1298 5 1 1 1297
0 1299 7 2 2 3286 1298
0 1300 5 1 1 3295
0 1301 7 1 2 2772 3296
0 1302 5 1 1 1301
0 1303 7 1 2 2769 1300
0 1304 5 1 1 1303
0 1305 7 1 2 3276 1270
0 1306 5 1 1 1305
0 1307 7 2 2 3280 1306
0 1308 5 1 1 3297
0 1309 7 1 2 2785 3298
0 1310 5 1 1 1309
0 1311 7 1 2 2782 1308
0 1312 5 1 1 1311
0 1313 7 1 2 3270 1262
0 1314 5 1 1 1313
0 1315 7 2 2 3274 1314
0 1316 5 1 1 3299
0 1317 7 1 2 2798 3300
0 1318 5 1 1 1317
0 1319 7 1 2 2795 1316
0 1320 5 1 1 1319
0 1321 7 1 2 3264 1254
0 1322 5 1 1 1321
0 1323 7 2 2 3268 1322
0 1324 5 1 1 3301
0 1325 7 1 2 2811 3302
0 1326 5 1 1 1325
0 1327 7 1 2 2808 1324
0 1328 5 1 1 1327
0 1329 7 1 2 3258 1246
0 1330 5 1 1 1329
0 1331 7 2 2 3262 1330
0 1332 5 1 1 3303
0 1333 7 1 2 2824 3304
0 1334 5 1 1 1333
0 1335 7 1 2 2821 1332
0 1336 5 1 1 1335
0 1337 7 1 2 3252 1238
0 1338 5 1 1 1337
0 1339 7 2 2 3256 1338
0 1340 5 1 1 3305
0 1341 7 1 2 2837 3306
0 1342 5 1 1 1341
0 1343 7 1 2 2834 1340
0 1344 5 1 1 1343
0 1345 7 1 2 3246 1230
0 1346 5 1 1 1345
0 1347 7 2 2 3250 1346
0 1348 5 1 1 3307
0 1349 7 1 2 2850 3308
0 1350 5 1 1 1349
0 1351 7 1 2 2847 1348
0 1352 5 1 1 1351
0 1353 7 1 2 3240 1222
0 1354 5 1 1 1353
0 1355 7 2 2 3244 1354
0 1356 5 1 1 3309
0 1357 7 1 2 2863 3310
0 1358 5 1 1 1357
0 1359 7 1 2 2860 1356
0 1360 5 1 1 1359
0 1361 7 1 2 3234 1214
0 1362 5 1 1 1361
0 1363 7 2 2 3238 1362
0 1364 5 1 1 3311
0 1365 7 1 2 2876 3312
0 1366 5 1 1 1365
0 1367 7 1 2 2873 1364
0 1368 5 1 1 1367
0 1369 7 1 2 3228 1206
0 1370 5 1 1 1369
0 1371 7 2 2 3232 1370
0 1372 5 1 1 3313
0 1373 7 1 2 2889 3314
0 1374 5 1 1 1373
0 1375 7 1 2 2886 1372
0 1376 5 1 1 1375
0 1377 7 1 2 3222 1198
0 1378 5 1 1 1377
0 1379 7 2 2 3226 1378
0 1380 5 1 1 3315
0 1381 7 1 2 2902 3316
0 1382 5 1 1 1381
0 1383 7 1 2 2899 1380
0 1384 5 1 1 1383
0 1385 7 1 2 3210 1182
0 1386 5 1 1 1385
0 1387 7 2 2 3214 1386
0 1388 5 1 1 3317
0 1389 7 1 2 3203 1174
0 1390 5 1 1 1389
0 1391 7 2 2 3208 1390
0 1392 5 1 1 3319
0 1393 7 1 2 2939 3320
0 1394 5 1 1 1393
0 1395 7 2 2 2943 3195
0 1396 5 1 1 3321
0 1397 7 2 2 2946 3322
0 1398 5 2 1 3323
0 1399 7 1 2 2952 3325
0 1400 5 2 1 1399
0 1401 7 1 2 3179 3197
0 1402 5 1 1 1401
0 1403 7 1 2 2950 2958
0 1404 7 1 2 3324 1403
0 1405 5 2 1 1404
0 1406 7 1 2 3204 3329
0 1407 7 1 2 1402 1406
0 1408 5 1 1 1407
0 1409 7 1 2 3327 1408
0 1410 7 1 2 1394 1409
0 1411 5 1 1 1410
0 1412 7 1 2 2936 1392
0 1413 5 1 1 1412
0 1414 7 2 2 1411 1413
0 1415 5 1 1 3331
0 1416 7 1 2 1388 1415
0 1417 5 1 1 1416
0 1418 7 1 2 2926 1417
0 1419 5 1 1 1418
0 1420 7 1 2 3318 3332
0 1421 5 1 1 1420
0 1422 7 1 2 1419 1421
0 1423 5 1 1 1422
0 1424 7 1 2 3216 1190
0 1425 5 1 1 1424
0 1426 7 2 2 3220 1425
0 1427 5 1 1 3333
0 1428 7 1 2 2912 1427
0 1429 5 1 1 1428
0 1430 7 1 2 1423 1429
0 1431 5 1 1 1430
0 1432 7 1 2 2915 3334
0 1433 5 1 1 1432
0 1434 7 1 2 1431 1433
0 1435 5 1 1 1434
0 1436 7 1 2 1384 1435
0 1437 5 1 1 1436
0 1438 7 1 2 1382 1437
0 1439 5 1 1 1438
0 1440 7 1 2 1376 1439
0 1441 5 1 1 1440
0 1442 7 1 2 1374 1441
0 1443 5 1 1 1442
0 1444 7 1 2 1368 1443
0 1445 5 1 1 1444
0 1446 7 1 2 1366 1445
0 1447 5 1 1 1446
0 1448 7 1 2 1360 1447
0 1449 5 1 1 1448
0 1450 7 1 2 1358 1449
0 1451 5 1 1 1450
0 1452 7 1 2 1352 1451
0 1453 5 1 1 1452
0 1454 7 1 2 1350 1453
0 1455 5 1 1 1454
0 1456 7 1 2 1344 1455
0 1457 5 1 1 1456
0 1458 7 1 2 1342 1457
0 1459 5 1 1 1458
0 1460 7 1 2 1336 1459
0 1461 5 1 1 1460
0 1462 7 1 2 1334 1461
0 1463 5 1 1 1462
0 1464 7 1 2 1328 1463
0 1465 5 1 1 1464
0 1466 7 1 2 1326 1465
0 1467 5 1 1 1466
0 1468 7 1 2 1320 1467
0 1469 5 1 1 1468
0 1470 7 1 2 1318 1469
0 1471 5 1 1 1470
0 1472 7 1 2 1312 1471
0 1473 5 1 1 1472
0 1474 7 1 2 1310 1473
0 1475 5 1 1 1474
0 1476 7 1 2 1304 1475
0 1477 5 1 1 1476
0 1478 7 1 2 1302 1477
0 1479 5 1 1 1478
0 1480 7 1 2 1296 1479
0 1481 5 1 1 1480
0 1482 7 1 2 2750 3294
0 1483 5 1 1 1482
0 1484 7 2 2 2947 1396
0 1485 5 2 1 3335
0 1486 7 1 2 2930 3337
0 1487 5 1 1 1486
0 1488 7 2 2 2933 1487
0 1489 5 2 1 3339
0 1490 7 1 2 2919 3341
0 1491 5 1 1 1490
0 1492 7 2 2 2922 1491
0 1493 5 2 1 3343
0 1494 7 1 2 2906 3345
0 1495 5 1 1 1494
0 1496 7 2 2 2909 1495
0 1497 5 2 1 3347
0 1498 7 1 2 2893 3349
0 1499 5 1 1 1498
0 1500 7 2 2 2896 1499
0 1501 5 2 1 3351
0 1502 7 1 2 2880 3353
0 1503 5 1 1 1502
0 1504 7 2 2 2883 1503
0 1505 5 2 1 3355
0 1506 7 1 2 2867 3357
0 1507 5 1 1 1506
0 1508 7 2 2 2870 1507
0 1509 5 2 1 3359
0 1510 7 1 2 2854 3361
0 1511 5 1 1 1510
0 1512 7 2 2 2857 1511
0 1513 5 2 1 3363
0 1514 7 1 2 2841 3365
0 1515 5 1 1 1514
0 1516 7 2 2 2844 1515
0 1517 5 2 1 3367
0 1518 7 1 2 2828 3369
0 1519 5 1 1 1518
0 1520 7 2 2 2831 1519
0 1521 5 2 1 3371
0 1522 7 1 2 2815 3373
0 1523 5 1 1 1522
0 1524 7 2 2 2818 1523
0 1525 5 2 1 3375
0 1526 7 1 2 2802 3377
0 1527 5 1 1 1526
0 1528 7 2 2 2805 1527
0 1529 5 2 1 3379
0 1530 7 1 2 2789 3381
0 1531 5 1 1 1530
0 1532 7 2 2 2792 1531
0 1533 5 2 1 3383
0 1534 7 1 2 2776 3385
0 1535 5 1 1 1534
0 1536 7 3 2 2779 1535
0 1537 5 3 1 3387
0 1538 7 1 2 2766 3390
0 1539 5 1 1 1538
0 1540 7 3 2 2760 1539
0 1541 5 2 1 3393
0 1542 7 1 2 3018 3394
0 1543 7 1 2 3292 1542
0 1544 7 1 2 1483 1543
0 1545 7 1 2 1481 1544
0 1546 5 1 1 1545
0 1547 7 1 2 3025 3384
0 1548 5 1 1 1547
0 1549 7 1 2 3023 3386
0 1550 5 1 1 1549
0 1551 7 3 2 1548 1550
0 1552 5 2 1 3398
0 1553 7 1 2 3395 3399
0 1554 5 2 1 1553
0 1555 7 1 2 3037 3388
0 1556 5 1 1 1555
0 1557 7 1 2 3035 3391
0 1558 5 1 1 1557
0 1559 7 2 2 1556 1558
0 1560 5 1 1 3405
0 1561 7 1 2 3044 3380
0 1562 5 1 1 1561
0 1563 7 1 2 3042 3382
0 1564 5 1 1 1563
0 1565 7 3 2 1562 1564
0 1566 5 2 1 3407
0 1567 7 1 2 3406 3408
0 1568 5 2 1 1567
0 1569 7 1 2 3056 3376
0 1570 5 1 1 1569
0 1571 7 1 2 3054 3378
0 1572 5 1 1 1571
0 1573 7 3 2 1570 1572
0 1574 5 2 1 3414
0 1575 7 1 2 3400 3415
0 1576 5 2 1 1575
0 1577 7 1 2 3068 3372
0 1578 5 1 1 1577
0 1579 7 1 2 3066 3374
0 1580 5 1 1 1579
0 1581 7 3 2 1578 1580
0 1582 5 2 1 3421
0 1583 7 1 2 3409 3422
0 1584 5 2 1 1583
0 1585 7 1 2 3080 3368
0 1586 5 1 1 1585
0 1587 7 1 2 3078 3370
0 1588 5 1 1 1587
0 1589 7 3 2 1586 1588
0 1590 5 2 1 3428
0 1591 7 1 2 3416 3429
0 1592 5 2 1 1591
0 1593 7 1 2 3092 3364
0 1594 5 1 1 1593
0 1595 7 1 2 3090 3366
0 1596 5 1 1 1595
0 1597 7 3 2 1594 1596
0 1598 5 2 1 3435
0 1599 7 1 2 3423 3436
0 1600 5 2 1 1599
0 1601 7 1 2 3104 3360
0 1602 5 1 1 1601
0 1603 7 1 2 3102 3362
0 1604 5 1 1 1603
0 1605 7 3 2 1602 1604
0 1606 5 2 1 3442
0 1607 7 1 2 3430 3443
0 1608 5 2 1 1607
0 1609 7 1 2 3116 3356
0 1610 5 1 1 1609
0 1611 7 1 2 3114 3358
0 1612 5 1 1 1611
0 1613 7 3 2 1610 1612
0 1614 5 2 1 3449
0 1615 7 1 2 3437 3450
0 1616 5 2 1 1615
0 1617 7 1 2 3128 3352
0 1618 5 1 1 1617
0 1619 7 1 2 3126 3354
0 1620 5 1 1 1619
0 1621 7 3 2 1618 1620
0 1622 5 2 1 3456
0 1623 7 1 2 3444 3457
0 1624 5 2 1 1623
0 1625 7 1 2 3140 3348
0 1626 5 1 1 1625
0 1627 7 1 2 3138 3350
0 1628 5 1 1 1627
0 1629 7 3 2 1626 1628
0 1630 5 2 1 3463
0 1631 7 1 2 3451 3464
0 1632 5 2 1 1631
0 1633 7 1 2 3152 3344
0 1634 5 1 1 1633
0 1635 7 1 2 3150 3346
0 1636 5 1 1 1635
0 1637 7 3 2 1634 1636
0 1638 5 2 1 3470
0 1639 7 1 2 3458 3471
0 1640 5 2 1 1639
0 1641 7 1 2 3164 3340
0 1642 5 1 1 1641
0 1643 7 1 2 3162 3342
0 1644 5 1 1 1643
0 1645 7 3 2 1642 1644
0 1646 5 2 1 3477
0 1647 7 1 2 3465 3478
0 1648 5 2 1 1647
0 1649 7 1 2 3176 3336
0 1650 5 1 1 1649
0 1651 7 1 2 3174 3338
0 1652 5 1 1 1651
0 1653 7 3 2 1650 1652
0 1654 5 2 1 3484
0 1655 7 1 2 3472 3485
0 1656 5 2 1 1655
0 1657 7 1 2 3187 3193
0 1658 5 1 1 1657
0 1659 7 2 2 3326 1658
0 1660 5 1 1 3491
0 1661 7 1 2 3479 3492
0 1662 5 2 1 1661
0 1663 7 2 2 3200 3486
0 1664 5 2 1 3495
0 1665 7 1 2 3480 1660
0 1666 5 1 1 1665
0 1667 7 2 2 3493 1666
0 1668 5 1 1 3499
0 1669 7 1 2 3496 3500
0 1670 5 2 1 1669
0 1671 7 2 2 3494 3501
0 1672 5 1 1 3503
0 1673 7 1 2 3473 3487
0 1674 5 1 1 1673
0 1675 7 2 2 3489 1674
0 1676 5 1 1 3505
0 1677 7 1 2 1672 3506
0 1678 5 2 1 1677
0 1679 7 2 2 3490 3507
0 1680 5 1 1 3509
0 1681 7 1 2 3466 3481
0 1682 5 1 1 1681
0 1683 7 2 2 3482 1682
0 1684 5 1 1 3511
0 1685 7 1 2 1680 3512
0 1686 5 2 1 1685
0 1687 7 2 2 3483 3513
0 1688 5 1 1 3515
0 1689 7 1 2 3459 3474
0 1690 5 1 1 1689
0 1691 7 2 2 3475 1690
0 1692 5 1 1 3517
0 1693 7 1 2 1688 3518
0 1694 5 2 1 1693
0 1695 7 2 2 3476 3519
0 1696 5 1 1 3521
0 1697 7 1 2 3452 3467
0 1698 5 1 1 1697
0 1699 7 2 2 3468 1698
0 1700 5 1 1 3523
0 1701 7 1 2 1696 3524
0 1702 5 2 1 1701
0 1703 7 2 2 3469 3525
0 1704 5 1 1 3527
0 1705 7 1 2 3445 3460
0 1706 5 1 1 1705
0 1707 7 2 2 3461 1706
0 1708 5 1 1 3529
0 1709 7 1 2 1704 3530
0 1710 5 2 1 1709
0 1711 7 2 2 3462 3531
0 1712 5 1 1 3533
0 1713 7 1 2 3438 3453
0 1714 5 1 1 1713
0 1715 7 2 2 3454 1714
0 1716 5 1 1 3535
0 1717 7 1 2 1712 3536
0 1718 5 2 1 1717
0 1719 7 2 2 3455 3537
0 1720 5 1 1 3539
0 1721 7 1 2 3431 3446
0 1722 5 1 1 1721
0 1723 7 2 2 3447 1722
0 1724 5 1 1 3541
0 1725 7 1 2 1720 3542
0 1726 5 2 1 1725
0 1727 7 2 2 3448 3543
0 1728 5 1 1 3545
0 1729 7 1 2 3424 3439
0 1730 5 1 1 1729
0 1731 7 2 2 3440 1730
0 1732 5 1 1 3547
0 1733 7 1 2 1728 3548
0 1734 5 2 1 1733
0 1735 7 2 2 3441 3549
0 1736 5 1 1 3551
0 1737 7 1 2 3417 3432
0 1738 5 1 1 1737
0 1739 7 2 2 3433 1738
0 1740 5 1 1 3553
0 1741 7 1 2 1736 3554
0 1742 5 2 1 1741
0 1743 7 2 2 3434 3555
0 1744 5 1 1 3557
0 1745 7 1 2 3410 3425
0 1746 5 1 1 1745
0 1747 7 2 2 3426 1746
0 1748 5 1 1 3559
0 1749 7 1 2 1744 3560
0 1750 5 2 1 1749
0 1751 7 2 2 3427 3561
0 1752 5 1 1 3563
0 1753 7 1 2 3401 3418
0 1754 5 1 1 1753
0 1755 7 2 2 3419 1754
0 1756 5 1 1 3565
0 1757 7 1 2 1752 3566
0 1758 5 2 1 1757
0 1759 7 2 2 3420 3567
0 1760 5 1 1 3569
0 1761 7 1 2 1560 3411
0 1762 5 1 1 1761
0 1763 7 2 2 3412 1762
0 1764 5 1 1 3571
0 1765 7 1 2 1760 3572
0 1766 5 2 1 1765
0 1767 7 2 2 3413 3573
0 1768 5 1 1 3575
0 1769 7 1 2 3396 3402
0 1770 5 1 1 1769
0 1771 7 2 2 3403 1770
0 1772 5 1 1 3577
0 1773 7 1 2 1768 3578
0 1774 5 2 1 1773
0 1775 7 2 2 3404 3579
0 1776 5 1 1 3581
0 1777 7 1 2 2757 3392
0 1778 5 1 1 1777
0 1779 7 1 2 2763 3389
0 1780 5 1 1 1779
0 1781 7 2 2 1778 1780
0 1782 5 1 1 3583
0 1783 7 1 2 1776 1782
0 1784 5 2 1 1783
0 1785 7 1 2 3582 3584
0 1786 5 2 1 1785
0 1787 7 1 2 3585 3587
0 1788 5 1 1 1787
0 1789 7 1 2 2754 1788
0 1790 5 1 1 1789
0 1791 7 1 2 3576 1772
0 1792 5 1 1 1791
0 1793 7 2 2 3580 1792
0 1794 5 1 1 3589
0 1795 7 1 2 2773 3590
0 1796 5 1 1 1795
0 1797 7 1 2 3570 1764
0 1798 5 1 1 1797
0 1799 7 2 2 3574 1798
0 1800 5 1 1 3591
0 1801 7 1 2 2783 1800
0 1802 5 1 1 1801
0 1803 7 1 2 2786 3592
0 1804 5 1 1 1803
0 1805 7 1 2 3564 1756
0 1806 5 1 1 1805
0 1807 7 2 2 3568 1806
0 1808 5 1 1 3593
0 1809 7 1 2 2796 1808
0 1810 5 1 1 1809
0 1811 7 1 2 2799 3594
0 1812 5 1 1 1811
0 1813 7 1 2 3558 1748
0 1814 5 1 1 1813
0 1815 7 2 2 3562 1814
0 1816 5 1 1 3595
0 1817 7 1 2 2809 1816
0 1818 5 1 1 1817
0 1819 7 1 2 2812 3596
0 1820 5 1 1 1819
0 1821 7 1 2 3552 1740
0 1822 5 1 1 1821
0 1823 7 2 2 3556 1822
0 1824 5 1 1 3597
0 1825 7 1 2 2822 1824
0 1826 5 1 1 1825
0 1827 7 1 2 2825 3598
0 1828 5 1 1 1827
0 1829 7 1 2 3546 1732
0 1830 5 1 1 1829
0 1831 7 2 2 3550 1830
0 1832 5 1 1 3599
0 1833 7 1 2 2838 3600
0 1834 5 1 1 1833
0 1835 7 1 2 2835 1832
0 1836 5 1 1 1835
0 1837 7 1 2 3540 1724
0 1838 5 1 1 1837
0 1839 7 2 2 3544 1838
0 1840 5 1 1 3601
0 1841 7 1 2 2851 3602
0 1842 5 1 1 1841
0 1843 7 1 2 2848 1840
0 1844 5 1 1 1843
0 1845 7 1 2 3534 1716
0 1846 5 1 1 1845
0 1847 7 2 2 3538 1846
0 1848 5 1 1 3603
0 1849 7 1 2 2864 3604
0 1850 5 1 1 1849
0 1851 7 1 2 2861 1848
0 1852 5 1 1 1851
0 1853 7 1 2 3528 1708
0 1854 5 1 1 1853
0 1855 7 2 2 3532 1854
0 1856 5 1 1 3605
0 1857 7 1 2 2877 3606
0 1858 5 1 1 1857
0 1859 7 1 2 2874 1856
0 1860 5 1 1 1859
0 1861 7 1 2 3522 1700
0 1862 5 1 1 1861
0 1863 7 2 2 3526 1862
0 1864 5 1 1 3607
0 1865 7 1 2 2890 3608
0 1866 5 1 1 1865
0 1867 7 1 2 2887 1864
0 1868 5 1 1 1867
0 1869 7 1 2 3516 1692
0 1870 5 1 1 1869
0 1871 7 2 2 3520 1870
0 1872 5 1 1 3609
0 1873 7 1 2 2903 3610
0 1874 5 1 1 1873
0 1875 7 1 2 2900 1872
0 1876 5 1 1 1875
0 1877 7 1 2 3504 1676
0 1878 5 1 1 1877
0 1879 7 2 2 3508 1878
0 1880 5 1 1 3611
0 1881 7 1 2 3497 1668
0 1882 5 1 1 1881
0 1883 7 2 2 3502 1882
0 1884 5 1 1 3613
0 1885 7 1 2 2940 3614
0 1886 5 1 1 1885
0 1887 7 1 2 3198 3488
0 1888 5 1 1 1887
0 1889 7 1 2 3330 3498
0 1890 7 1 2 1888 1889
0 1891 5 1 1 1890
0 1892 7 1 2 3328 1891
0 1893 7 1 2 1886 1892
0 1894 5 1 1 1893
0 1895 7 1 2 2937 1884
0 1896 5 1 1 1895
0 1897 7 2 2 1894 1896
0 1898 5 1 1 3615
0 1899 7 1 2 1880 1898
0 1900 5 1 1 1899
0 1901 7 1 2 2927 1900
0 1902 5 1 1 1901
0 1903 7 1 2 3612 3616
0 1904 5 1 1 1903
0 1905 7 1 2 1902 1904
0 1906 5 1 1 1905
0 1907 7 1 2 3510 1684
0 1908 5 1 1 1907
0 1909 7 2 2 3514 1908
0 1910 5 1 1 3617
0 1911 7 1 2 2913 1910
0 1912 5 1 1 1911
0 1913 7 1 2 1906 1912
0 1914 5 1 1 1913
0 1915 7 1 2 2916 3618
0 1916 5 1 1 1915
0 1917 7 1 2 1914 1916
0 1918 5 1 1 1917
0 1919 7 1 2 1876 1918
0 1920 5 1 1 1919
0 1921 7 1 2 1874 1920
0 1922 5 1 1 1921
0 1923 7 1 2 1868 1922
0 1924 5 1 1 1923
0 1925 7 1 2 1866 1924
0 1926 5 1 1 1925
0 1927 7 1 2 1860 1926
0 1928 5 1 1 1927
0 1929 7 1 2 1858 1928
0 1930 5 1 1 1929
0 1931 7 1 2 1852 1930
0 1932 5 1 1 1931
0 1933 7 1 2 1850 1932
0 1934 5 1 1 1933
0 1935 7 1 2 1844 1934
0 1936 5 1 1 1935
0 1937 7 1 2 1842 1936
0 1938 5 1 1 1937
0 1939 7 1 2 1836 1938
0 1940 5 1 1 1939
0 1941 7 1 2 1834 1940
0 1942 7 1 2 1828 1941
0 1943 5 1 1 1942
0 1944 7 1 2 1826 1943
0 1945 5 1 1 1944
0 1946 7 1 2 1820 1945
0 1947 5 1 1 1946
0 1948 7 1 2 1818 1947
0 1949 5 1 1 1948
0 1950 7 1 2 1812 1949
0 1951 5 1 1 1950
0 1952 7 1 2 1810 1951
0 1953 5 1 1 1952
0 1954 7 1 2 1804 1953
0 1955 5 1 1 1954
0 1956 7 1 2 1802 1955
0 1957 5 1 1 1956
0 1958 7 1 2 1796 1957
0 1959 5 1 1 1958
0 1960 7 1 2 2770 1794
0 1961 5 1 1 1960
0 1962 7 1 2 1959 1961
0 1963 7 1 2 1790 1962
0 1964 5 1 1 1963
0 1965 7 1 2 2751 3588
0 1966 5 1 1 1965
0 1967 7 1 2 3397 3586
0 1968 7 1 2 1966 1967
0 1969 7 1 2 1964 1968
0 1970 5 1 1 1969
0 1971 7 1 2 1546 1970
3 4299 5 0 1 1971
