1 0 0 3 0
2 13 1 0
2 14 1 0
2 15 1 0
1 1 0 2 0
2 16 1 1
2 17 1 1
1 2 0 2 0
2 18 1 2
2 19 1 2
1 3 0 2 0
2 44 1 3
2 64 1 3
1 4 0 2 0
2 83 1 4
2 103 1 4
1 5 0 2 0
2 126 1 5
2 147 1 5
1 6 0 2 0
2 154 1 6
2 155 1 6
1 7 0 2 0
2 156 1 7
2 157 1 7
1 8 0 2 0
2 158 1 8
2 159 1 8
1 9 0 2 0
2 160 1 9
2 161 1 9
1 10 0 2 0
2 162 1 10
2 163 1 10
1 11 0 2 0
2 164 1 11
2 165 1 11
1 12 0 2 0
2 166 1 12
2 167 1 12
2 168 1 20
2 169 1 20
2 170 1 34
2 171 1 34
2 172 1 34
2 173 1 36
2 174 1 36
2 175 1 36
2 176 1 37
2 177 1 37
2 178 1 48
2 179 1 48
2 180 1 48
2 181 1 50
2 182 1 50
2 183 1 50
2 184 1 50
2 185 1 52
2 186 1 52
2 187 1 52
2 188 1 53
2 189 1 53
2 190 1 60
2 191 1 60
2 192 1 66
2 193 1 66
2 194 1 66
2 195 1 66
2 196 1 70
2 197 1 70
2 198 1 70
2 199 1 71
2 200 1 71
2 201 1 72
2 202 1 72
2 203 1 84
2 204 1 84
2 205 1 89
2 206 1 89
2 207 1 91
2 208 1 91
2 209 1 91
2 210 1 91
2 211 1 93
2 212 1 93
2 213 1 93
2 214 1 93
2 215 1 94
2 216 1 94
2 217 1 100
2 218 1 100
2 219 1 105
2 220 1 105
2 221 1 105
2 222 1 106
2 223 1 106
2 224 1 107
2 225 1 107
2 226 1 107
2 227 1 108
2 228 1 108
2 229 1 108
2 230 1 116
2 231 1 116
2 232 1 116
2 233 1 121
2 234 1 121
2 235 1 128
2 236 1 128
2 237 1 130
2 238 1 130
2 239 1 131
2 240 1 131
2 241 1 131
0 20 5 2 1 13
0 21 5 1 1 16
0 22 5 1 1 18
0 23 5 1 1 44
0 24 5 1 1 83
0 25 5 1 1 126
0 26 5 1 1 154
0 27 5 1 1 156
0 28 5 1 1 158
0 29 5 1 1 160
0 30 5 1 1 162
0 31 5 1 1 164
0 32 5 1 1 166
0 33 7 1 2 155 167
0 34 5 3 1 33
0 35 7 1 2 26 32
0 36 5 3 1 35
0 37 7 2 2 170 173
0 38 5 1 1 176
0 39 7 1 2 14 38
0 40 5 1 1 39
0 41 7 1 2 168 177
0 42 5 1 1 41
0 43 7 1 2 40 42
3 593 5 0 1 43
0 45 7 1 2 15 174
0 46 5 1 1 45
0 47 7 1 2 171 46
0 48 5 3 1 47
0 49 7 1 2 17 157
0 50 5 4 1 49
0 51 7 1 2 21 27
0 52 5 3 1 51
0 53 7 2 2 181 185
0 54 5 1 1 188
0 55 7 1 2 178 54
0 56 5 1 1 55
0 57 7 1 2 169 172
0 58 5 1 1 57
0 59 7 1 2 175 58
0 60 5 2 1 59
0 61 7 1 2 189 190
0 62 5 1 1 61
0 63 7 1 2 56 62
3 594 5 0 1 63
0 65 7 1 2 19 159
0 66 5 4 1 65
0 67 7 1 2 182 191
0 68 5 1 1 67
0 69 7 1 2 22 28
0 70 5 3 1 69
0 71 7 2 2 186 196
0 72 7 2 2 68 199
0 73 5 1 1 201
0 74 7 1 2 192 202
0 75 5 1 1 74
0 76 7 1 2 179 187
0 77 5 1 1 76
0 78 7 1 2 193 197
0 79 5 1 1 78
0 80 7 1 2 183 79
0 81 7 1 2 77 80
0 82 5 1 1 81
3 595 7 0 2 75 82
0 84 7 2 2 180 200
0 85 5 1 1 203
0 86 7 1 2 184 194
0 87 5 1 1 86
0 88 7 1 2 198 87
0 89 5 2 1 88
0 90 7 1 2 64 161
0 91 5 4 1 90
0 92 7 1 2 23 29
0 93 5 4 1 92
0 94 7 2 2 207 211
0 95 5 1 1 215
0 96 7 1 2 205 95
0 97 7 1 2 85 96
0 98 5 1 1 97
0 99 7 1 2 195 73
0 100 5 2 1 99
0 101 7 1 2 216 217
0 102 5 1 1 101
3 596 7 0 2 98 102
0 104 7 1 2 103 163
0 105 5 3 1 104
0 106 7 2 2 24 30
0 107 5 3 1 222
0 108 7 3 2 219 224
0 109 5 1 1 227
0 110 7 1 2 206 208
0 111 5 1 1 110
0 112 7 1 2 212 111
0 113 5 1 1 112
0 114 7 1 2 204 213
0 115 5 1 1 114
0 116 7 3 2 113 115
0 117 5 1 1 230
0 118 7 1 2 109 117
0 119 5 1 1 118
0 120 7 1 2 214 218
0 121 5 2 1 120
0 122 7 1 2 209 228
0 123 7 1 2 233 122
0 124 5 1 1 123
0 125 7 1 2 119 124
3 597 5 0 1 125
0 127 7 1 2 147 165
0 128 5 2 1 127
0 129 7 1 2 25 31
0 130 5 2 1 129
0 131 7 3 2 235 237
0 132 5 1 1 239
0 133 7 1 2 210 220
0 134 7 1 2 240 133
0 135 7 1 2 234 134
0 136 5 1 1 135
0 137 7 1 2 229 231
0 138 5 1 1 137
0 139 7 1 2 223 132
0 140 5 1 1 139
0 141 7 1 2 225 241
0 142 5 1 1 141
0 143 7 1 2 140 142
0 144 7 1 2 138 143
0 145 5 1 1 144
0 146 7 1 2 136 145
3 598 5 0 1 146
0 148 7 1 2 221 232
0 149 5 1 1 148
0 150 7 1 2 226 238
0 151 7 1 2 149 150
0 152 5 1 1 151
0 153 7 1 2 236 152
3 599 5 0 1 153
