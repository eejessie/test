1 0 0 3 0
2 21 1 0
2 22 1 0
2 23 1 0
1 1 0 2 0
2 24 1 1
2 25 1 1
1 2 0 2 0
2 26 1 2
2 27 1 2
1 3 0 2 0
2 28 1 3
2 29 1 3
1 4 0 2 0
2 30 1 4
2 31 1 4
1 5 0 2 0
2 64 1 5
2 84 1 5
1 6 0 2 0
2 102 1 6
2 124 1 6
1 7 0 2 0
2 142 1 7
2 165 1 7
1 8 0 2 0
2 191 1 8
2 214 1 8
1 9 0 2 0
2 233 1 9
2 271 1 9
1 10 0 2 0
2 274 1 10
2 275 1 10
1 11 0 2 0
2 276 1 11
2 277 1 11
1 12 0 2 0
2 278 1 12
2 279 1 12
1 13 0 2 0
2 280 1 13
2 281 1 13
1 14 0 2 0
2 282 1 14
2 283 1 14
1 15 0 2 0
2 284 1 15
2 285 1 15
1 16 0 2 0
2 286 1 16
2 287 1 16
1 17 0 2 0
2 288 1 17
2 289 1 17
1 18 0 2 0
2 290 1 18
2 291 1 18
1 19 0 2 0
2 292 1 19
2 293 1 19
1 20 0 2 0
2 294 1 20
2 295 1 20
2 296 1 32
2 297 1 32
2 298 1 54
2 299 1 54
2 300 1 54
2 301 1 56
2 302 1 56
2 303 1 56
2 304 1 57
2 305 1 57
2 306 1 68
2 307 1 68
2 308 1 70
2 309 1 70
2 310 1 70
2 311 1 70
2 312 1 71
2 313 1 71
2 314 1 72
2 315 1 72
2 316 1 72
2 317 1 73
2 318 1 73
2 319 1 80
2 320 1 80
2 321 1 80
2 322 1 86
2 323 1 86
2 324 1 86
2 325 1 86
2 326 1 88
2 327 1 88
2 328 1 88
2 329 1 89
2 330 1 89
2 331 1 93
2 332 1 93
2 333 1 97
2 334 1 97
2 335 1 98
2 336 1 98
2 337 1 104
2 338 1 104
2 339 1 104
2 340 1 104
2 341 1 106
2 342 1 106
2 343 1 106
2 344 1 109
2 345 1 109
2 346 1 109
2 347 1 114
2 348 1 114
2 349 1 117
2 350 1 117
2 351 1 117
2 352 1 117
2 353 1 120
2 354 1 120
2 355 1 126
2 356 1 126
2 357 1 126
2 358 1 126
2 359 1 126
2 360 1 126
2 361 1 128
2 362 1 128
2 363 1 129
2 364 1 129
2 365 1 129
2 366 1 130
2 367 1 130
2 368 1 144
2 369 1 144
2 370 1 144
2 371 1 144
2 372 1 146
2 373 1 146
2 374 1 146
2 375 1 146
2 376 1 147
2 377 1 147
2 378 1 149
2 379 1 149
2 380 1 154
2 381 1 154
2 382 1 154
2 383 1 161
2 384 1 161
2 385 1 167
2 386 1 167
2 387 1 167
2 388 1 167
2 389 1 169
2 390 1 169
2 391 1 169
2 392 1 171
2 393 1 171
2 394 1 175
2 395 1 175
2 396 1 180
2 397 1 180
2 398 1 180
2 399 1 181
2 400 1 181
2 401 1 193
2 402 1 193
2 403 1 193
2 404 1 195
2 405 1 195
2 406 1 195
2 407 1 195
2 408 1 195
2 409 1 195
2 410 1 201
2 411 1 201
2 412 1 202
2 413 1 202
2 414 1 208
2 415 1 208
2 416 1 209
2 417 1 209
2 418 1 218
2 419 1 218
2 420 1 220
2 421 1 220
2 422 1 220
2 423 1 222
2 424 1 222
2 425 1 222
2 426 1 223
2 427 1 223
2 428 1 226
2 429 1 226
2 430 1 235
2 431 1 235
2 432 1 237
2 433 1 237
2 434 1 238
2 435 1 238
2 436 1 244
2 437 1 244
0 32 5 2 1 21
0 33 5 1 1 24
0 34 5 1 1 26
0 35 5 1 1 28
0 36 5 1 1 30
0 37 5 1 1 64
0 38 5 1 1 102
0 39 5 1 1 142
0 40 5 1 1 191
0 41 5 1 1 233
0 42 5 1 1 274
0 43 5 1 1 276
0 44 5 1 1 278
0 45 5 1 1 280
0 46 5 1 1 282
0 47 5 1 1 284
0 48 5 1 1 286
0 49 5 1 1 288
0 50 5 1 1 290
0 51 5 1 1 292
0 52 5 1 1 294
0 53 7 1 2 275 295
0 54 5 3 1 53
0 55 7 1 2 42 52
0 56 5 3 1 55
0 57 7 2 2 298 301
0 58 5 1 1 304
0 59 7 1 2 22 58
0 60 5 1 1 59
0 61 7 1 2 296 305
0 62 5 1 1 61
0 63 7 1 2 60 62
3 589 5 0 1 63
0 65 7 1 2 23 302
0 66 5 1 1 65
0 67 7 1 2 299 66
0 68 5 2 1 67
0 69 7 1 2 25 277
0 70 5 4 1 69
0 71 7 2 2 33 43
0 72 5 3 1 312
0 73 7 2 2 308 314
0 74 5 1 1 317
0 75 7 1 2 306 74
0 76 5 1 1 75
0 77 7 1 2 297 300
0 78 5 1 1 77
0 79 7 1 2 303 78
0 80 5 3 1 79
0 81 7 1 2 318 319
0 82 5 1 1 81
0 83 7 1 2 76 82
3 590 5 0 1 83
0 85 7 1 2 27 279
0 86 5 4 1 85
0 87 7 1 2 34 44
0 88 5 3 1 87
0 89 7 2 2 322 326
0 90 5 1 1 329
0 91 7 1 2 309 320
0 92 5 1 1 91
0 93 7 2 2 315 92
0 94 5 1 1 331
0 95 7 1 2 330 332
0 96 5 1 1 95
0 97 7 2 2 307 316
0 98 5 2 1 333
0 99 7 1 2 310 90
0 100 7 1 2 335 99
0 101 5 1 1 100
3 591 7 0 2 96 101
0 103 7 1 2 29 281
0 104 5 4 1 103
0 105 7 1 2 35 45
0 106 5 3 1 105
0 107 7 1 2 337 341
0 108 5 1 1 107
0 109 7 3 2 311 323
0 110 5 1 1 344
0 111 7 1 2 336 345
0 112 5 1 1 111
0 113 7 1 2 327 112
0 114 5 2 1 113
0 115 7 1 2 108 347
0 116 5 1 1 115
0 117 7 4 2 328 342
0 118 7 1 2 324 94
0 119 5 1 1 118
0 120 7 2 2 349 119
0 121 5 1 1 353
0 122 7 1 2 338 354
0 123 5 1 1 122
3 592 7 0 2 116 123
0 125 7 1 2 36 46
0 126 5 6 1 125
0 127 7 1 2 31 283
0 128 5 2 1 127
0 129 7 3 2 339 361
0 130 7 2 2 121 363
0 131 5 1 1 366
0 132 7 1 2 355 367
0 133 5 1 1 132
0 134 7 1 2 340 348
0 135 5 1 1 134
0 136 7 1 2 356 362
0 137 5 1 1 136
0 138 7 1 2 343 137
0 139 7 1 2 135 138
0 140 5 1 1 139
0 141 7 1 2 133 140
3 593 5 0 1 141
0 143 7 1 2 84 285
0 144 5 4 1 143
0 145 7 1 2 37 47
0 146 5 4 1 145
0 147 7 2 2 368 372
0 148 5 1 1 376
0 149 7 2 2 357 131
0 150 5 1 1 378
0 151 7 1 2 377 379
0 152 5 1 1 151
0 153 7 1 2 350 358
0 154 7 3 2 334 153
0 155 5 1 1 380
0 156 7 1 2 110 351
0 157 5 1 1 156
0 158 7 1 2 364 157
0 159 5 1 1 158
0 160 7 1 2 359 159
0 161 5 2 1 160
0 162 7 1 2 148 383
0 163 7 1 2 155 162
0 164 5 1 1 163
3 594 7 0 2 152 164
0 166 7 1 2 124 287
0 167 5 4 1 166
0 168 7 1 2 38 48
0 169 5 3 1 168
0 170 7 1 2 385 389
0 171 5 2 1 170
0 172 7 1 2 369 384
0 173 5 1 1 172
0 174 7 1 2 373 173
0 175 5 2 1 174
0 176 7 1 2 392 394
0 177 5 1 1 176
0 178 7 1 2 370 150
0 179 5 1 1 178
0 180 7 3 2 374 390
0 181 7 2 2 179 396
0 182 5 1 1 399
0 183 7 1 2 386 400
0 184 5 1 1 183
0 185 7 1 2 177 184
0 186 5 1 1 185
0 187 7 1 2 375 393
0 188 7 1 2 381 187
0 189 5 1 1 188
0 190 7 1 2 186 189
3 595 5 0 1 190
0 192 7 1 2 165 289
0 193 5 3 1 192
0 194 7 1 2 39 49
0 195 5 6 1 194
0 196 7 1 2 401 404
0 197 5 1 1 196
0 198 7 1 2 387 395
0 199 5 1 1 198
0 200 7 1 2 391 199
0 201 5 2 1 200
0 202 7 2 2 382 397
0 203 5 1 1 412
0 204 7 1 2 410 203
0 205 5 1 1 204
0 206 7 1 2 197 205
0 207 5 1 1 206
0 208 7 2 2 388 402
0 209 7 2 2 182 414
0 210 5 1 1 416
0 211 7 1 2 405 417
0 212 5 1 1 211
0 213 7 1 2 207 212
3 596 5 0 1 213
0 215 7 1 2 403 411
0 216 5 1 1 215
0 217 7 1 2 406 216
0 218 5 2 1 217
0 219 7 1 2 214 291
0 220 5 3 1 219
0 221 7 1 2 40 50
0 222 5 3 1 221
0 223 7 2 2 420 423
0 224 5 1 1 426
0 225 7 1 2 407 413
0 226 5 2 1 225
0 227 7 1 2 224 428
0 228 7 1 2 418 227
0 229 5 1 1 228
0 230 7 1 2 408 427
0 231 7 1 2 210 230
0 232 5 1 1 231
3 597 7 0 2 229 232
0 234 7 1 2 271 293
0 235 5 2 1 234
0 236 7 1 2 41 51
0 237 5 2 1 236
0 238 7 2 2 430 432
0 239 5 1 1 434
0 240 7 1 2 421 429
0 241 7 1 2 419 240
0 242 5 1 1 241
0 243 7 1 2 424 242
0 244 5 2 1 243
0 245 7 1 2 239 436
0 246 5 1 1 245
0 247 7 1 2 321 346
0 248 5 1 1 247
0 249 7 1 2 313 325
0 250 5 1 1 249
0 251 7 1 2 352 250
0 252 7 1 2 248 251
0 253 5 1 1 252
0 254 7 1 2 365 253
0 255 5 1 1 254
0 256 7 1 2 360 255
0 257 5 1 1 256
0 258 7 1 2 371 257
0 259 5 1 1 258
0 260 7 1 2 398 259
0 261 5 1 1 260
0 262 7 1 2 415 261
0 263 5 1 1 262
0 264 7 1 2 409 263
0 265 5 1 1 264
0 266 7 1 2 422 265
0 267 5 1 1 266
0 268 7 1 2 425 435
0 269 7 1 2 267 268
0 270 5 1 1 269
3 598 7 0 2 246 270
0 272 7 1 2 431 437
0 273 5 1 1 272
3 599 7 0 2 433 273
