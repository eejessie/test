1 0 0 291 0
2 25 1 0
2 26 1 0
2 47734 1 0
2 47735 1 0
2 47736 1 0
2 47737 1 0
2 47738 1 0
2 47739 1 0
2 47740 1 0
2 47741 1 0
2 47742 1 0
2 47743 1 0
2 47744 1 0
2 47745 1 0
2 47746 1 0
2 47747 1 0
2 47748 1 0
2 47749 1 0
2 47750 1 0
2 47751 1 0
2 47752 1 0
2 47753 1 0
2 47754 1 0
2 47755 1 0
2 47756 1 0
2 47757 1 0
2 47758 1 0
2 47759 1 0
2 47760 1 0
2 47761 1 0
2 47762 1 0
2 47763 1 0
2 47764 1 0
2 47765 1 0
2 47766 1 0
2 47767 1 0
2 47768 1 0
2 47769 1 0
2 47770 1 0
2 47771 1 0
2 47772 1 0
2 47773 1 0
2 47774 1 0
2 47775 1 0
2 47776 1 0
2 47777 1 0
2 47778 1 0
2 47779 1 0
2 47780 1 0
2 47781 1 0
2 47782 1 0
2 47783 1 0
2 47784 1 0
2 47785 1 0
2 47786 1 0
2 47787 1 0
2 47788 1 0
2 47789 1 0
2 47790 1 0
2 47791 1 0
2 47792 1 0
2 47793 1 0
2 47794 1 0
2 47795 1 0
2 47796 1 0
2 47797 1 0
2 47798 1 0
2 47799 1 0
2 47800 1 0
2 47801 1 0
2 47802 1 0
2 47803 1 0
2 47804 1 0
2 47805 1 0
2 47806 1 0
2 47807 1 0
2 47808 1 0
2 47809 1 0
2 47810 1 0
2 47811 1 0
2 47812 1 0
2 47813 1 0
2 47814 1 0
2 47815 1 0
2 47816 1 0
2 47817 1 0
2 47818 1 0
2 47819 1 0
2 47820 1 0
2 47821 1 0
2 47822 1 0
2 47823 1 0
2 47824 1 0
2 47825 1 0
2 47826 1 0
2 47827 1 0
2 47828 1 0
2 47829 1 0
2 47830 1 0
2 47831 1 0
2 47832 1 0
2 47833 1 0
2 47834 1 0
2 47835 1 0
2 47836 1 0
2 47837 1 0
2 47838 1 0
2 47839 1 0
2 47840 1 0
2 47841 1 0
2 47842 1 0
2 47843 1 0
2 47844 1 0
2 47845 1 0
2 47846 1 0
2 47847 1 0
2 47848 1 0
2 47849 1 0
2 47850 1 0
2 47851 1 0
2 47852 1 0
2 47853 1 0
2 47854 1 0
2 47855 1 0
2 47856 1 0
2 47857 1 0
2 47858 1 0
2 47859 1 0
2 47860 1 0
2 47861 1 0
2 47862 1 0
2 47863 1 0
2 47864 1 0
2 47865 1 0
2 47866 1 0
2 47867 1 0
2 47868 1 0
2 47869 1 0
2 47870 1 0
2 47871 1 0
2 47872 1 0
2 47873 1 0
2 47874 1 0
2 47875 1 0
2 47876 1 0
2 47877 1 0
2 47878 1 0
2 47879 1 0
2 47880 1 0
2 47881 1 0
2 47882 1 0
2 47883 1 0
2 47884 1 0
2 47885 1 0
2 47886 1 0
2 47887 1 0
2 47888 1 0
2 47889 1 0
2 47890 1 0
2 47891 1 0
2 47892 1 0
2 47893 1 0
2 47894 1 0
2 47895 1 0
2 47896 1 0
2 47897 1 0
2 47898 1 0
2 47899 1 0
2 47900 1 0
2 47901 1 0
2 47902 1 0
2 47903 1 0
2 47904 1 0
2 47905 1 0
2 47906 1 0
2 47907 1 0
2 47908 1 0
2 47909 1 0
2 47910 1 0
2 47911 1 0
2 47912 1 0
2 47913 1 0
2 47914 1 0
2 47915 1 0
2 47916 1 0
2 47917 1 0
2 47918 1 0
2 47919 1 0
2 47920 1 0
2 47921 1 0
2 47922 1 0
2 47923 1 0
2 47924 1 0
2 47925 1 0
2 47926 1 0
2 47927 1 0
2 47928 1 0
2 47929 1 0
2 47930 1 0
2 47931 1 0
2 47932 1 0
2 47933 1 0
2 47934 1 0
2 47935 1 0
2 47936 1 0
2 47937 1 0
2 47938 1 0
2 47939 1 0
2 47940 1 0
2 47941 1 0
2 47942 1 0
2 47943 1 0
2 47944 1 0
2 47945 1 0
2 47946 1 0
2 47947 1 0
2 47948 1 0
2 47949 1 0
2 47950 1 0
2 47951 1 0
2 47952 1 0
2 47953 1 0
2 47954 1 0
2 47955 1 0
2 47956 1 0
2 47957 1 0
2 47958 1 0
2 47959 1 0
2 47960 1 0
2 47961 1 0
2 47962 1 0
2 47963 1 0
2 47964 1 0
2 47965 1 0
2 47966 1 0
2 47967 1 0
2 47968 1 0
2 47969 1 0
2 47970 1 0
2 47971 1 0
2 47972 1 0
2 47973 1 0
2 47974 1 0
2 47975 1 0
2 47976 1 0
2 47977 1 0
2 47978 1 0
2 47979 1 0
2 47980 1 0
2 47981 1 0
2 47982 1 0
2 47983 1 0
2 47984 1 0
2 47985 1 0
2 47986 1 0
2 47987 1 0
2 47988 1 0
2 47989 1 0
2 47990 1 0
2 47991 1 0
2 47992 1 0
2 47993 1 0
2 47994 1 0
2 47995 1 0
2 47996 1 0
2 47997 1 0
2 47998 1 0
2 47999 1 0
2 48000 1 0
2 48001 1 0
2 48002 1 0
2 48003 1 0
2 48004 1 0
2 48005 1 0
2 48006 1 0
2 48007 1 0
2 48008 1 0
2 48009 1 0
2 48010 1 0
2 48011 1 0
2 48012 1 0
2 48013 1 0
2 48014 1 0
2 48015 1 0
2 48016 1 0
2 48017 1 0
2 48018 1 0
2 48019 1 0
2 48020 1 0
2 48021 1 0
2 48022 1 0
1 1 0 255 0
2 48023 1 1
2 48024 1 1
2 48025 1 1
2 48026 1 1
2 48027 1 1
2 48028 1 1
2 48029 1 1
2 48030 1 1
2 48031 1 1
2 48032 1 1
2 48033 1 1
2 48034 1 1
2 48035 1 1
2 48036 1 1
2 48037 1 1
2 48038 1 1
2 48039 1 1
2 48040 1 1
2 48041 1 1
2 48042 1 1
2 48043 1 1
2 48044 1 1
2 48045 1 1
2 48046 1 1
2 48047 1 1
2 48048 1 1
2 48049 1 1
2 48050 1 1
2 48051 1 1
2 48052 1 1
2 48053 1 1
2 48054 1 1
2 48055 1 1
2 48056 1 1
2 48057 1 1
2 48058 1 1
2 48059 1 1
2 48060 1 1
2 48061 1 1
2 48062 1 1
2 48063 1 1
2 48064 1 1
2 48065 1 1
2 48066 1 1
2 48067 1 1
2 48068 1 1
2 48069 1 1
2 48070 1 1
2 48071 1 1
2 48072 1 1
2 48073 1 1
2 48074 1 1
2 48075 1 1
2 48076 1 1
2 48077 1 1
2 48078 1 1
2 48079 1 1
2 48080 1 1
2 48081 1 1
2 48082 1 1
2 48083 1 1
2 48084 1 1
2 48085 1 1
2 48086 1 1
2 48087 1 1
2 48088 1 1
2 48089 1 1
2 48090 1 1
2 48091 1 1
2 48092 1 1
2 48093 1 1
2 48094 1 1
2 48095 1 1
2 48096 1 1
2 48097 1 1
2 48098 1 1
2 48099 1 1
2 48100 1 1
2 48101 1 1
2 48102 1 1
2 48103 1 1
2 48104 1 1
2 48105 1 1
2 48106 1 1
2 48107 1 1
2 48108 1 1
2 48109 1 1
2 48110 1 1
2 48111 1 1
2 48112 1 1
2 48113 1 1
2 48114 1 1
2 48115 1 1
2 48116 1 1
2 48117 1 1
2 48118 1 1
2 48119 1 1
2 48120 1 1
2 48121 1 1
2 48122 1 1
2 48123 1 1
2 48124 1 1
2 48125 1 1
2 48126 1 1
2 48127 1 1
2 48128 1 1
2 48129 1 1
2 48130 1 1
2 48131 1 1
2 48132 1 1
2 48133 1 1
2 48134 1 1
2 48135 1 1
2 48136 1 1
2 48137 1 1
2 48138 1 1
2 48139 1 1
2 48140 1 1
2 48141 1 1
2 48142 1 1
2 48143 1 1
2 48144 1 1
2 48145 1 1
2 48146 1 1
2 48147 1 1
2 48148 1 1
2 48149 1 1
2 48150 1 1
2 48151 1 1
2 48152 1 1
2 48153 1 1
2 48154 1 1
2 48155 1 1
2 48156 1 1
2 48157 1 1
2 48158 1 1
2 48159 1 1
2 48160 1 1
2 48161 1 1
2 48162 1 1
2 48163 1 1
2 48164 1 1
2 48165 1 1
2 48166 1 1
2 48167 1 1
2 48168 1 1
2 48169 1 1
2 48170 1 1
2 48171 1 1
2 48172 1 1
2 48173 1 1
2 48174 1 1
2 48175 1 1
2 48176 1 1
2 48177 1 1
2 48178 1 1
2 48179 1 1
2 48180 1 1
2 48181 1 1
2 48182 1 1
2 48183 1 1
2 48184 1 1
2 48185 1 1
2 48186 1 1
2 48187 1 1
2 48188 1 1
2 48189 1 1
2 48190 1 1
2 48191 1 1
2 48192 1 1
2 48193 1 1
2 48194 1 1
2 48195 1 1
2 48196 1 1
2 48197 1 1
2 48198 1 1
2 48199 1 1
2 48200 1 1
2 48201 1 1
2 48202 1 1
2 48203 1 1
2 48204 1 1
2 48205 1 1
2 48206 1 1
2 48207 1 1
2 48208 1 1
2 48209 1 1
2 48210 1 1
2 48211 1 1
2 48212 1 1
2 48213 1 1
2 48214 1 1
2 48215 1 1
2 48216 1 1
2 48217 1 1
2 48218 1 1
2 48219 1 1
2 48220 1 1
2 48221 1 1
2 48222 1 1
2 48223 1 1
2 48224 1 1
2 48225 1 1
2 48226 1 1
2 48227 1 1
2 48228 1 1
2 48229 1 1
2 48230 1 1
2 48231 1 1
2 48232 1 1
2 48233 1 1
2 48234 1 1
2 48235 1 1
2 48236 1 1
2 48237 1 1
2 48238 1 1
2 48239 1 1
2 48240 1 1
2 48241 1 1
2 48242 1 1
2 48243 1 1
2 48244 1 1
2 48245 1 1
2 48246 1 1
2 48247 1 1
2 48248 1 1
2 48249 1 1
2 48250 1 1
2 48251 1 1
2 48252 1 1
2 48253 1 1
2 48254 1 1
2 48255 1 1
2 48256 1 1
2 48257 1 1
2 48258 1 1
2 48259 1 1
2 48260 1 1
2 48261 1 1
2 48262 1 1
2 48263 1 1
2 48264 1 1
2 48265 1 1
2 48266 1 1
2 48267 1 1
2 48268 1 1
2 48269 1 1
2 48270 1 1
2 48271 1 1
2 48272 1 1
2 48273 1 1
2 48274 1 1
2 48275 1 1
2 48276 1 1
2 48277 1 1
1 2 0 175 0
2 48278 1 2
2 48279 1 2
2 48280 1 2
2 48281 1 2
2 48282 1 2
2 48283 1 2
2 48284 1 2
2 48285 1 2
2 48286 1 2
2 48287 1 2
2 48288 1 2
2 48289 1 2
2 48290 1 2
2 48291 1 2
2 48292 1 2
2 48293 1 2
2 48294 1 2
2 48295 1 2
2 48296 1 2
2 48297 1 2
2 48298 1 2
2 48299 1 2
2 48300 1 2
2 48301 1 2
2 48302 1 2
2 48303 1 2
2 48304 1 2
2 48305 1 2
2 48306 1 2
2 48307 1 2
2 48308 1 2
2 48309 1 2
2 48310 1 2
2 48311 1 2
2 48312 1 2
2 48313 1 2
2 48314 1 2
2 48315 1 2
2 48316 1 2
2 48317 1 2
2 48318 1 2
2 48319 1 2
2 48320 1 2
2 48321 1 2
2 48322 1 2
2 48323 1 2
2 48324 1 2
2 48325 1 2
2 48326 1 2
2 48327 1 2
2 48328 1 2
2 48329 1 2
2 48330 1 2
2 48331 1 2
2 48332 1 2
2 48333 1 2
2 48334 1 2
2 48335 1 2
2 48336 1 2
2 48337 1 2
2 48338 1 2
2 48339 1 2
2 48340 1 2
2 48341 1 2
2 48342 1 2
2 48343 1 2
2 48344 1 2
2 48345 1 2
2 48346 1 2
2 48347 1 2
2 48348 1 2
2 48349 1 2
2 48350 1 2
2 48351 1 2
2 48352 1 2
2 48353 1 2
2 48354 1 2
2 48355 1 2
2 48356 1 2
2 48357 1 2
2 48358 1 2
2 48359 1 2
2 48360 1 2
2 48361 1 2
2 48362 1 2
2 48363 1 2
2 48364 1 2
2 48365 1 2
2 48366 1 2
2 48367 1 2
2 48368 1 2
2 48369 1 2
2 48370 1 2
2 48371 1 2
2 48372 1 2
2 48373 1 2
2 48374 1 2
2 48375 1 2
2 48376 1 2
2 48377 1 2
2 48378 1 2
2 48379 1 2
2 48380 1 2
2 48381 1 2
2 48382 1 2
2 48383 1 2
2 48384 1 2
2 48385 1 2
2 48386 1 2
2 48387 1 2
2 48388 1 2
2 48389 1 2
2 48390 1 2
2 48391 1 2
2 48392 1 2
2 48393 1 2
2 48394 1 2
2 48395 1 2
2 48396 1 2
2 48397 1 2
2 48398 1 2
2 48399 1 2
2 48400 1 2
2 48401 1 2
2 48402 1 2
2 48403 1 2
2 48404 1 2
2 48405 1 2
2 48406 1 2
2 48407 1 2
2 48408 1 2
2 48409 1 2
2 48410 1 2
2 48411 1 2
2 48412 1 2
2 48413 1 2
2 48414 1 2
2 48415 1 2
2 48416 1 2
2 48417 1 2
2 48418 1 2
2 48419 1 2
2 48420 1 2
2 48421 1 2
2 48422 1 2
2 48423 1 2
2 48424 1 2
2 48425 1 2
2 48426 1 2
2 48427 1 2
2 48428 1 2
2 48429 1 2
2 48430 1 2
2 48431 1 2
2 48432 1 2
2 48433 1 2
2 48434 1 2
2 48435 1 2
2 48436 1 2
2 48437 1 2
2 48438 1 2
2 48439 1 2
2 48440 1 2
2 48441 1 2
2 48442 1 2
2 48443 1 2
2 48444 1 2
2 48445 1 2
2 48446 1 2
2 48447 1 2
2 48448 1 2
2 48449 1 2
2 48450 1 2
2 48451 1 2
2 48452 1 2
1 3 0 114 0
2 48453 1 3
2 48454 1 3
2 48455 1 3
2 48456 1 3
2 48457 1 3
2 48458 1 3
2 48459 1 3
2 48460 1 3
2 48461 1 3
2 48462 1 3
2 48463 1 3
2 48464 1 3
2 48465 1 3
2 48466 1 3
2 48467 1 3
2 48468 1 3
2 48469 1 3
2 48470 1 3
2 48471 1 3
2 48472 1 3
2 48473 1 3
2 48474 1 3
2 48475 1 3
2 48476 1 3
2 48477 1 3
2 48478 1 3
2 48479 1 3
2 48480 1 3
2 48481 1 3
2 48482 1 3
2 48483 1 3
2 48484 1 3
2 48485 1 3
2 48486 1 3
2 48487 1 3
2 48488 1 3
2 48489 1 3
2 48490 1 3
2 48491 1 3
2 48492 1 3
2 48493 1 3
2 48494 1 3
2 48495 1 3
2 48496 1 3
2 48497 1 3
2 48498 1 3
2 48499 1 3
2 48500 1 3
2 48501 1 3
2 48502 1 3
2 48503 1 3
2 48504 1 3
2 48505 1 3
2 48506 1 3
2 48507 1 3
2 48508 1 3
2 48509 1 3
2 48510 1 3
2 48511 1 3
2 48512 1 3
2 48513 1 3
2 48514 1 3
2 48515 1 3
2 48516 1 3
2 48517 1 3
2 48518 1 3
2 48519 1 3
2 48520 1 3
2 48521 1 3
2 48522 1 3
2 48523 1 3
2 48524 1 3
2 48525 1 3
2 48526 1 3
2 48527 1 3
2 48528 1 3
2 48529 1 3
2 48530 1 3
2 48531 1 3
2 48532 1 3
2 48533 1 3
2 48534 1 3
2 48535 1 3
2 48536 1 3
2 48537 1 3
2 48538 1 3
2 48539 1 3
2 48540 1 3
2 48541 1 3
2 48542 1 3
2 48543 1 3
2 48544 1 3
2 48545 1 3
2 48546 1 3
2 48547 1 3
2 48548 1 3
2 48549 1 3
2 48550 1 3
2 48551 1 3
2 48552 1 3
2 48553 1 3
2 48554 1 3
2 48555 1 3
2 48556 1 3
2 48557 1 3
2 48558 1 3
2 48559 1 3
2 48560 1 3
2 48561 1 3
2 48562 1 3
2 48563 1 3
2 48564 1 3
2 48565 1 3
2 48566 1 3
1 4 0 111 0
2 48567 1 4
2 48568 1 4
2 48569 1 4
2 48570 1 4
2 48571 1 4
2 48572 1 4
2 48573 1 4
2 48574 1 4
2 48575 1 4
2 48576 1 4
2 48577 1 4
2 48578 1 4
2 48579 1 4
2 48580 1 4
2 48581 1 4
2 48582 1 4
2 48583 1 4
2 48584 1 4
2 48585 1 4
2 48586 1 4
2 48587 1 4
2 48588 1 4
2 48589 1 4
2 48590 1 4
2 48591 1 4
2 48592 1 4
2 48593 1 4
2 48594 1 4
2 48595 1 4
2 48596 1 4
2 48597 1 4
2 48598 1 4
2 48599 1 4
2 48600 1 4
2 48601 1 4
2 48602 1 4
2 48603 1 4
2 48604 1 4
2 48605 1 4
2 48606 1 4
2 48607 1 4
2 48608 1 4
2 48609 1 4
2 48610 1 4
2 48611 1 4
2 48612 1 4
2 48613 1 4
2 48614 1 4
2 48615 1 4
2 48616 1 4
2 48617 1 4
2 48618 1 4
2 48619 1 4
2 48620 1 4
2 48621 1 4
2 48622 1 4
2 48623 1 4
2 48624 1 4
2 48625 1 4
2 48626 1 4
2 48627 1 4
2 48628 1 4
2 48629 1 4
2 48630 1 4
2 48631 1 4
2 48632 1 4
2 48633 1 4
2 48634 1 4
2 48635 1 4
2 48636 1 4
2 48637 1 4
2 48638 1 4
2 48639 1 4
2 48640 1 4
2 48641 1 4
2 48642 1 4
2 48643 1 4
2 48644 1 4
2 48645 1 4
2 48646 1 4
2 48647 1 4
2 48648 1 4
2 48649 1 4
2 48650 1 4
2 48651 1 4
2 48652 1 4
2 48653 1 4
2 48654 1 4
2 48655 1 4
2 48656 1 4
2 48657 1 4
2 48658 1 4
2 48659 1 4
2 48660 1 4
2 48661 1 4
2 48662 1 4
2 48663 1 4
2 48664 1 4
2 48665 1 4
2 48666 1 4
2 48667 1 4
2 48668 1 4
2 48669 1 4
2 48670 1 4
2 48671 1 4
2 48672 1 4
2 48673 1 4
2 48674 1 4
2 48675 1 4
2 48676 1 4
2 48677 1 4
1 5 0 158 0
2 48678 1 5
2 48679 1 5
2 48680 1 5
2 48681 1 5
2 48682 1 5
2 48683 1 5
2 48684 1 5
2 48685 1 5
2 48686 1 5
2 48687 1 5
2 48688 1 5
2 48689 1 5
2 48690 1 5
2 48691 1 5
2 48692 1 5
2 48693 1 5
2 48694 1 5
2 48695 1 5
2 48696 1 5
2 48697 1 5
2 48698 1 5
2 48699 1 5
2 48700 1 5
2 48701 1 5
2 48702 1 5
2 48703 1 5
2 48704 1 5
2 48705 1 5
2 48706 1 5
2 48707 1 5
2 48708 1 5
2 48709 1 5
2 48710 1 5
2 48711 1 5
2 48712 1 5
2 48713 1 5
2 48714 1 5
2 48715 1 5
2 48716 1 5
2 48717 1 5
2 48718 1 5
2 48719 1 5
2 48720 1 5
2 48721 1 5
2 48722 1 5
2 48723 1 5
2 48724 1 5
2 48725 1 5
2 48726 1 5
2 48727 1 5
2 48728 1 5
2 48729 1 5
2 48730 1 5
2 48731 1 5
2 48732 1 5
2 48733 1 5
2 48734 1 5
2 48735 1 5
2 48736 1 5
2 48737 1 5
2 48738 1 5
2 48739 1 5
2 48740 1 5
2 48741 1 5
2 48742 1 5
2 48743 1 5
2 48744 1 5
2 48745 1 5
2 48746 1 5
2 48747 1 5
2 48748 1 5
2 48749 1 5
2 48750 1 5
2 48751 1 5
2 48752 1 5
2 48753 1 5
2 48754 1 5
2 48755 1 5
2 48756 1 5
2 48757 1 5
2 48758 1 5
2 48759 1 5
2 48760 1 5
2 48761 1 5
2 48762 1 5
2 48763 1 5
2 48764 1 5
2 48765 1 5
2 48766 1 5
2 48767 1 5
2 48768 1 5
2 48769 1 5
2 48770 1 5
2 48771 1 5
2 48772 1 5
2 48773 1 5
2 48774 1 5
2 48775 1 5
2 48776 1 5
2 48777 1 5
2 48778 1 5
2 48779 1 5
2 48780 1 5
2 48781 1 5
2 48782 1 5
2 48783 1 5
2 48784 1 5
2 48785 1 5
2 48786 1 5
2 48787 1 5
2 48788 1 5
2 48789 1 5
2 48790 1 5
2 48791 1 5
2 48792 1 5
2 48793 1 5
2 48794 1 5
2 48795 1 5
2 48796 1 5
2 48797 1 5
2 48798 1 5
2 48799 1 5
2 48800 1 5
2 48801 1 5
2 48802 1 5
2 48803 1 5
2 48804 1 5
2 48805 1 5
2 48806 1 5
2 48807 1 5
2 48808 1 5
2 48809 1 5
2 48810 1 5
2 48811 1 5
2 48812 1 5
2 48813 1 5
2 48814 1 5
2 48815 1 5
2 48816 1 5
2 48817 1 5
2 48818 1 5
2 48819 1 5
2 48820 1 5
2 48821 1 5
2 48822 1 5
2 48823 1 5
2 48824 1 5
2 48825 1 5
2 48826 1 5
2 48827 1 5
2 48828 1 5
2 48829 1 5
2 48830 1 5
2 48831 1 5
2 48832 1 5
2 48833 1 5
2 48834 1 5
2 48835 1 5
1 6 0 147 0
2 48836 1 6
2 48837 1 6
2 48838 1 6
2 48839 1 6
2 48840 1 6
2 48841 1 6
2 48842 1 6
2 48843 1 6
2 48844 1 6
2 48845 1 6
2 48846 1 6
2 48847 1 6
2 48848 1 6
2 48849 1 6
2 48850 1 6
2 48851 1 6
2 48852 1 6
2 48853 1 6
2 48854 1 6
2 48855 1 6
2 48856 1 6
2 48857 1 6
2 48858 1 6
2 48859 1 6
2 48860 1 6
2 48861 1 6
2 48862 1 6
2 48863 1 6
2 48864 1 6
2 48865 1 6
2 48866 1 6
2 48867 1 6
2 48868 1 6
2 48869 1 6
2 48870 1 6
2 48871 1 6
2 48872 1 6
2 48873 1 6
2 48874 1 6
2 48875 1 6
2 48876 1 6
2 48877 1 6
2 48878 1 6
2 48879 1 6
2 48880 1 6
2 48881 1 6
2 48882 1 6
2 48883 1 6
2 48884 1 6
2 48885 1 6
2 48886 1 6
2 48887 1 6
2 48888 1 6
2 48889 1 6
2 48890 1 6
2 48891 1 6
2 48892 1 6
2 48893 1 6
2 48894 1 6
2 48895 1 6
2 48896 1 6
2 48897 1 6
2 48898 1 6
2 48899 1 6
2 48900 1 6
2 48901 1 6
2 48902 1 6
2 48903 1 6
2 48904 1 6
2 48905 1 6
2 48906 1 6
2 48907 1 6
2 48908 1 6
2 48909 1 6
2 48910 1 6
2 48911 1 6
2 48912 1 6
2 48913 1 6
2 48914 1 6
2 48915 1 6
2 48916 1 6
2 48917 1 6
2 48918 1 6
2 48919 1 6
2 48920 1 6
2 48921 1 6
2 48922 1 6
2 48923 1 6
2 48924 1 6
2 48925 1 6
2 48926 1 6
2 48927 1 6
2 48928 1 6
2 48929 1 6
2 48930 1 6
2 48931 1 6
2 48932 1 6
2 48933 1 6
2 48934 1 6
2 48935 1 6
2 48936 1 6
2 48937 1 6
2 48938 1 6
2 48939 1 6
2 48940 1 6
2 48941 1 6
2 48942 1 6
2 48943 1 6
2 48944 1 6
2 48945 1 6
2 48946 1 6
2 48947 1 6
2 48948 1 6
2 48949 1 6
2 48950 1 6
2 48951 1 6
2 48952 1 6
2 48953 1 6
2 48954 1 6
2 48955 1 6
2 48956 1 6
2 48957 1 6
2 48958 1 6
2 48959 1 6
2 48960 1 6
2 48961 1 6
2 48962 1 6
2 48963 1 6
2 48964 1 6
2 48965 1 6
2 48966 1 6
2 48967 1 6
2 48968 1 6
2 48969 1 6
2 48970 1 6
2 48971 1 6
2 48972 1 6
2 48973 1 6
2 48974 1 6
2 48975 1 6
2 48976 1 6
2 48977 1 6
2 48978 1 6
2 48979 1 6
2 48980 1 6
2 48981 1 6
2 48982 1 6
1 7 0 99 0
2 48983 1 7
2 48984 1 7
2 48985 1 7
2 48986 1 7
2 48987 1 7
2 48988 1 7
2 48989 1 7
2 48990 1 7
2 48991 1 7
2 48992 1 7
2 48993 1 7
2 48994 1 7
2 48995 1 7
2 48996 1 7
2 48997 1 7
2 48998 1 7
2 48999 1 7
2 49000 1 7
2 49001 1 7
2 49002 1 7
2 49003 1 7
2 49004 1 7
2 49005 1 7
2 49006 1 7
2 49007 1 7
2 49008 1 7
2 49009 1 7
2 49010 1 7
2 49011 1 7
2 49012 1 7
2 49013 1 7
2 49014 1 7
2 49015 1 7
2 49016 1 7
2 49017 1 7
2 49018 1 7
2 49019 1 7
2 49020 1 7
2 49021 1 7
2 49022 1 7
2 49023 1 7
2 49024 1 7
2 49025 1 7
2 49026 1 7
2 49027 1 7
2 49028 1 7
2 49029 1 7
2 49030 1 7
2 49031 1 7
2 49032 1 7
2 49033 1 7
2 49034 1 7
2 49035 1 7
2 49036 1 7
2 49037 1 7
2 49038 1 7
2 49039 1 7
2 49040 1 7
2 49041 1 7
2 49042 1 7
2 49043 1 7
2 49044 1 7
2 49045 1 7
2 49046 1 7
2 49047 1 7
2 49048 1 7
2 49049 1 7
2 49050 1 7
2 49051 1 7
2 49052 1 7
2 49053 1 7
2 49054 1 7
2 49055 1 7
2 49056 1 7
2 49057 1 7
2 49058 1 7
2 49059 1 7
2 49060 1 7
2 49061 1 7
2 49062 1 7
2 49063 1 7
2 49064 1 7
2 49065 1 7
2 49066 1 7
2 49067 1 7
2 49068 1 7
2 49069 1 7
2 49070 1 7
2 49071 1 7
2 49072 1 7
2 49073 1 7
2 49074 1 7
2 49075 1 7
2 49076 1 7
2 49077 1 7
2 49078 1 7
2 49079 1 7
2 49080 1 7
2 49081 1 7
1 8 0 57 0
2 49082 1 8
2 49083 1 8
2 49084 1 8
2 49085 1 8
2 49086 1 8
2 49087 1 8
2 49088 1 8
2 49089 1 8
2 49090 1 8
2 49091 1 8
2 49092 1 8
2 49093 1 8
2 49094 1 8
2 49095 1 8
2 49096 1 8
2 49097 1 8
2 49098 1 8
2 49099 1 8
2 49100 1 8
2 49101 1 8
2 49102 1 8
2 49103 1 8
2 49104 1 8
2 49105 1 8
2 49106 1 8
2 49107 1 8
2 49108 1 8
2 49109 1 8
2 49110 1 8
2 49111 1 8
2 49112 1 8
2 49113 1 8
2 49114 1 8
2 49115 1 8
2 49116 1 8
2 49117 1 8
2 49118 1 8
2 49119 1 8
2 49120 1 8
2 49121 1 8
2 49122 1 8
2 49123 1 8
2 49124 1 8
2 49125 1 8
2 49126 1 8
2 49127 1 8
2 49128 1 8
2 49129 1 8
2 49130 1 8
2 49131 1 8
2 49132 1 8
2 49133 1 8
2 49134 1 8
2 49135 1 8
2 49136 1 8
2 49137 1 8
2 49138 1 8
1 9 0 121 0
2 49139 1 9
2 49140 1 9
2 49141 1 9
2 49142 1 9
2 49143 1 9
2 49144 1 9
2 49145 1 9
2 49146 1 9
2 49147 1 9
2 49148 1 9
2 49149 1 9
2 49150 1 9
2 49151 1 9
2 49152 1 9
2 49153 1 9
2 49154 1 9
2 49155 1 9
2 49156 1 9
2 49157 1 9
2 49158 1 9
2 49159 1 9
2 49160 1 9
2 49161 1 9
2 49162 1 9
2 49163 1 9
2 49164 1 9
2 49165 1 9
2 49166 1 9
2 49167 1 9
2 49168 1 9
2 49169 1 9
2 49170 1 9
2 49171 1 9
2 49172 1 9
2 49173 1 9
2 49174 1 9
2 49175 1 9
2 49176 1 9
2 49177 1 9
2 49178 1 9
2 49179 1 9
2 49180 1 9
2 49181 1 9
2 49182 1 9
2 49183 1 9
2 49184 1 9
2 49185 1 9
2 49186 1 9
2 49187 1 9
2 49188 1 9
2 49189 1 9
2 49190 1 9
2 49191 1 9
2 49192 1 9
2 49193 1 9
2 49194 1 9
2 49195 1 9
2 49196 1 9
2 49197 1 9
2 49198 1 9
2 49199 1 9
2 49200 1 9
2 49201 1 9
2 49202 1 9
2 49203 1 9
2 49204 1 9
2 49205 1 9
2 49206 1 9
2 49207 1 9
2 49208 1 9
2 49209 1 9
2 49210 1 9
2 49211 1 9
2 49212 1 9
2 49213 1 9
2 49214 1 9
2 49215 1 9
2 49216 1 9
2 49217 1 9
2 49218 1 9
2 49219 1 9
2 49220 1 9
2 49221 1 9
2 49222 1 9
2 49223 1 9
2 49224 1 9
2 49225 1 9
2 49226 1 9
2 49227 1 9
2 49228 1 9
2 49229 1 9
2 49230 1 9
2 49231 1 9
2 49232 1 9
2 49233 1 9
2 49234 1 9
2 49235 1 9
2 49236 1 9
2 49237 1 9
2 49238 1 9
2 49239 1 9
2 49240 1 9
2 49241 1 9
2 49242 1 9
2 49243 1 9
2 49244 1 9
2 49245 1 9
2 49246 1 9
2 49247 1 9
2 49248 1 9
2 49249 1 9
2 49250 1 9
2 49251 1 9
2 49252 1 9
2 49253 1 9
2 49254 1 9
2 49255 1 9
2 49256 1 9
2 49257 1 9
2 49258 1 9
2 49259 1 9
1 10 0 124 0
2 49260 1 10
2 49261 1 10
2 49262 1 10
2 49263 1 10
2 49264 1 10
2 49265 1 10
2 49266 1 10
2 49267 1 10
2 49268 1 10
2 49269 1 10
2 49270 1 10
2 49271 1 10
2 49272 1 10
2 49273 1 10
2 49274 1 10
2 49275 1 10
2 49276 1 10
2 49277 1 10
2 49278 1 10
2 49279 1 10
2 49280 1 10
2 49281 1 10
2 49282 1 10
2 49283 1 10
2 49284 1 10
2 49285 1 10
2 49286 1 10
2 49287 1 10
2 49288 1 10
2 49289 1 10
2 49290 1 10
2 49291 1 10
2 49292 1 10
2 49293 1 10
2 49294 1 10
2 49295 1 10
2 49296 1 10
2 49297 1 10
2 49298 1 10
2 49299 1 10
2 49300 1 10
2 49301 1 10
2 49302 1 10
2 49303 1 10
2 49304 1 10
2 49305 1 10
2 49306 1 10
2 49307 1 10
2 49308 1 10
2 49309 1 10
2 49310 1 10
2 49311 1 10
2 49312 1 10
2 49313 1 10
2 49314 1 10
2 49315 1 10
2 49316 1 10
2 49317 1 10
2 49318 1 10
2 49319 1 10
2 49320 1 10
2 49321 1 10
2 49322 1 10
2 49323 1 10
2 49324 1 10
2 49325 1 10
2 49326 1 10
2 49327 1 10
2 49328 1 10
2 49329 1 10
2 49330 1 10
2 49331 1 10
2 49332 1 10
2 49333 1 10
2 49334 1 10
2 49335 1 10
2 49336 1 10
2 49337 1 10
2 49338 1 10
2 49339 1 10
2 49340 1 10
2 49341 1 10
2 49342 1 10
2 49343 1 10
2 49344 1 10
2 49345 1 10
2 49346 1 10
2 49347 1 10
2 49348 1 10
2 49349 1 10
2 49350 1 10
2 49351 1 10
2 49352 1 10
2 49353 1 10
2 49354 1 10
2 49355 1 10
2 49356 1 10
2 49357 1 10
2 49358 1 10
2 49359 1 10
2 49360 1 10
2 49361 1 10
2 49362 1 10
2 49363 1 10
2 49364 1 10
2 49365 1 10
2 49366 1 10
2 49367 1 10
2 49368 1 10
2 49369 1 10
2 49370 1 10
2 49371 1 10
2 49372 1 10
2 49373 1 10
2 49374 1 10
2 49375 1 10
2 49376 1 10
2 49377 1 10
2 49378 1 10
2 49379 1 10
2 49380 1 10
2 49381 1 10
2 49382 1 10
2 49383 1 10
1 11 0 122 0
2 49384 1 11
2 49385 1 11
2 49386 1 11
2 49387 1 11
2 49388 1 11
2 49389 1 11
2 49390 1 11
2 49391 1 11
2 49392 1 11
2 49393 1 11
2 49394 1 11
2 49395 1 11
2 49396 1 11
2 49397 1 11
2 49398 1 11
2 49399 1 11
2 49400 1 11
2 49401 1 11
2 49402 1 11
2 49403 1 11
2 49404 1 11
2 49405 1 11
2 49406 1 11
2 49407 1 11
2 49408 1 11
2 49409 1 11
2 49410 1 11
2 49411 1 11
2 49412 1 11
2 49413 1 11
2 49414 1 11
2 49415 1 11
2 49416 1 11
2 49417 1 11
2 49418 1 11
2 49419 1 11
2 49420 1 11
2 49421 1 11
2 49422 1 11
2 49423 1 11
2 49424 1 11
2 49425 1 11
2 49426 1 11
2 49427 1 11
2 49428 1 11
2 49429 1 11
2 49430 1 11
2 49431 1 11
2 49432 1 11
2 49433 1 11
2 49434 1 11
2 49435 1 11
2 49436 1 11
2 49437 1 11
2 49438 1 11
2 49439 1 11
2 49440 1 11
2 49441 1 11
2 49442 1 11
2 49443 1 11
2 49444 1 11
2 49445 1 11
2 49446 1 11
2 49447 1 11
2 49448 1 11
2 49449 1 11
2 49450 1 11
2 49451 1 11
2 49452 1 11
2 49453 1 11
2 49454 1 11
2 49455 1 11
2 49456 1 11
2 49457 1 11
2 49458 1 11
2 49459 1 11
2 49460 1 11
2 49461 1 11
2 49462 1 11
2 49463 1 11
2 49464 1 11
2 49465 1 11
2 49466 1 11
2 49467 1 11
2 49468 1 11
2 49469 1 11
2 49470 1 11
2 49471 1 11
2 49472 1 11
2 49473 1 11
2 49474 1 11
2 49475 1 11
2 49476 1 11
2 49477 1 11
2 49478 1 11
2 49479 1 11
2 49480 1 11
2 49481 1 11
2 49482 1 11
2 49483 1 11
2 49484 1 11
2 49485 1 11
2 49486 1 11
2 49487 1 11
2 49488 1 11
2 49489 1 11
2 49490 1 11
2 49491 1 11
2 49492 1 11
2 49493 1 11
2 49494 1 11
2 49495 1 11
2 49496 1 11
2 49497 1 11
2 49498 1 11
2 49499 1 11
2 49500 1 11
2 49501 1 11
2 49502 1 11
2 49503 1 11
2 49504 1 11
2 49505 1 11
1 12 0 140 0
2 49506 1 12
2 49507 1 12
2 49508 1 12
2 49509 1 12
2 49510 1 12
2 49511 1 12
2 49512 1 12
2 49513 1 12
2 49514 1 12
2 49515 1 12
2 49516 1 12
2 49517 1 12
2 49518 1 12
2 49519 1 12
2 49520 1 12
2 49521 1 12
2 49522 1 12
2 49523 1 12
2 49524 1 12
2 49525 1 12
2 49526 1 12
2 49527 1 12
2 49528 1 12
2 49529 1 12
2 49530 1 12
2 49531 1 12
2 49532 1 12
2 49533 1 12
2 49534 1 12
2 49535 1 12
2 49536 1 12
2 49537 1 12
2 49538 1 12
2 49539 1 12
2 49540 1 12
2 49541 1 12
2 49542 1 12
2 49543 1 12
2 49544 1 12
2 49545 1 12
2 49546 1 12
2 49547 1 12
2 49548 1 12
2 49549 1 12
2 49550 1 12
2 49551 1 12
2 49552 1 12
2 49553 1 12
2 49554 1 12
2 49555 1 12
2 49556 1 12
2 49557 1 12
2 49558 1 12
2 49559 1 12
2 49560 1 12
2 49561 1 12
2 49562 1 12
2 49563 1 12
2 49564 1 12
2 49565 1 12
2 49566 1 12
2 49567 1 12
2 49568 1 12
2 49569 1 12
2 49570 1 12
2 49571 1 12
2 49572 1 12
2 49573 1 12
2 49574 1 12
2 49575 1 12
2 49576 1 12
2 49577 1 12
2 49578 1 12
2 49579 1 12
2 49580 1 12
2 49581 1 12
2 49582 1 12
2 49583 1 12
2 49584 1 12
2 49585 1 12
2 49586 1 12
2 49587 1 12
2 49588 1 12
2 49589 1 12
2 49590 1 12
2 49591 1 12
2 49592 1 12
2 49593 1 12
2 49594 1 12
2 49595 1 12
2 49596 1 12
2 49597 1 12
2 49598 1 12
2 49599 1 12
2 49600 1 12
2 49601 1 12
2 49602 1 12
2 49603 1 12
2 49604 1 12
2 49605 1 12
2 49606 1 12
2 49607 1 12
2 49608 1 12
2 49609 1 12
2 49610 1 12
2 49611 1 12
2 49612 1 12
2 49613 1 12
2 49614 1 12
2 49615 1 12
2 49616 1 12
2 49617 1 12
2 49618 1 12
2 49619 1 12
2 49620 1 12
2 49621 1 12
2 49622 1 12
2 49623 1 12
2 49624 1 12
2 49625 1 12
2 49626 1 12
2 49627 1 12
2 49628 1 12
2 49629 1 12
2 49630 1 12
2 49631 1 12
2 49632 1 12
2 49633 1 12
2 49634 1 12
2 49635 1 12
2 49636 1 12
2 49637 1 12
2 49638 1 12
2 49639 1 12
2 49640 1 12
2 49641 1 12
2 49642 1 12
2 49643 1 12
2 49644 1 12
2 49645 1 12
1 13 0 183 0
2 49646 1 13
2 49647 1 13
2 49648 1 13
2 49649 1 13
2 49650 1 13
2 49651 1 13
2 49652 1 13
2 49653 1 13
2 49654 1 13
2 49655 1 13
2 49656 1 13
2 49657 1 13
2 49658 1 13
2 49659 1 13
2 49660 1 13
2 49661 1 13
2 49662 1 13
2 49663 1 13
2 49664 1 13
2 49665 1 13
2 49666 1 13
2 49667 1 13
2 49668 1 13
2 49669 1 13
2 49670 1 13
2 49671 1 13
2 49672 1 13
2 49673 1 13
2 49674 1 13
2 49675 1 13
2 49676 1 13
2 49677 1 13
2 49678 1 13
2 49679 1 13
2 49680 1 13
2 49681 1 13
2 49682 1 13
2 49683 1 13
2 49684 1 13
2 49685 1 13
2 49686 1 13
2 49687 1 13
2 49688 1 13
2 49689 1 13
2 49690 1 13
2 49691 1 13
2 49692 1 13
2 49693 1 13
2 49694 1 13
2 49695 1 13
2 49696 1 13
2 49697 1 13
2 49698 1 13
2 49699 1 13
2 49700 1 13
2 49701 1 13
2 49702 1 13
2 49703 1 13
2 49704 1 13
2 49705 1 13
2 49706 1 13
2 49707 1 13
2 49708 1 13
2 49709 1 13
2 49710 1 13
2 49711 1 13
2 49712 1 13
2 49713 1 13
2 49714 1 13
2 49715 1 13
2 49716 1 13
2 49717 1 13
2 49718 1 13
2 49719 1 13
2 49720 1 13
2 49721 1 13
2 49722 1 13
2 49723 1 13
2 49724 1 13
2 49725 1 13
2 49726 1 13
2 49727 1 13
2 49728 1 13
2 49729 1 13
2 49730 1 13
2 49731 1 13
2 49732 1 13
2 49733 1 13
2 49734 1 13
2 49735 1 13
2 49736 1 13
2 49737 1 13
2 49738 1 13
2 49739 1 13
2 49740 1 13
2 49741 1 13
2 49742 1 13
2 49743 1 13
2 49744 1 13
2 49745 1 13
2 49746 1 13
2 49747 1 13
2 49748 1 13
2 49749 1 13
2 49750 1 13
2 49751 1 13
2 49752 1 13
2 49753 1 13
2 49754 1 13
2 49755 1 13
2 49756 1 13
2 49757 1 13
2 49758 1 13
2 49759 1 13
2 49760 1 13
2 49761 1 13
2 49762 1 13
2 49763 1 13
2 49764 1 13
2 49765 1 13
2 49766 1 13
2 49767 1 13
2 49768 1 13
2 49769 1 13
2 49770 1 13
2 49771 1 13
2 49772 1 13
2 49773 1 13
2 49774 1 13
2 49775 1 13
2 49776 1 13
2 49777 1 13
2 49778 1 13
2 49779 1 13
2 49780 1 13
2 49781 1 13
2 49782 1 13
2 49783 1 13
2 49784 1 13
2 49785 1 13
2 49786 1 13
2 49787 1 13
2 49788 1 13
2 49789 1 13
2 49790 1 13
2 49791 1 13
2 49792 1 13
2 49793 1 13
2 49794 1 13
2 49795 1 13
2 49796 1 13
2 49797 1 13
2 49798 1 13
2 49799 1 13
2 49800 1 13
2 49801 1 13
2 49802 1 13
2 49803 1 13
2 49804 1 13
2 49805 1 13
2 49806 1 13
2 49807 1 13
2 49808 1 13
2 49809 1 13
2 49810 1 13
2 49811 1 13
2 49812 1 13
2 49813 1 13
2 49814 1 13
2 49815 1 13
2 49816 1 13
2 49817 1 13
2 49818 1 13
2 49819 1 13
2 49820 1 13
2 49821 1 13
2 49822 1 13
2 49823 1 13
2 49824 1 13
2 49825 1 13
2 49826 1 13
2 49827 1 13
2 49828 1 13
1 14 0 162 0
2 49829 1 14
2 49830 1 14
2 49831 1 14
2 49832 1 14
2 49833 1 14
2 49834 1 14
2 49835 1 14
2 49836 1 14
2 49837 1 14
2 49838 1 14
2 49839 1 14
2 49840 1 14
2 49841 1 14
2 49842 1 14
2 49843 1 14
2 49844 1 14
2 49845 1 14
2 49846 1 14
2 49847 1 14
2 49848 1 14
2 49849 1 14
2 49850 1 14
2 49851 1 14
2 49852 1 14
2 49853 1 14
2 49854 1 14
2 49855 1 14
2 49856 1 14
2 49857 1 14
2 49858 1 14
2 49859 1 14
2 49860 1 14
2 49861 1 14
2 49862 1 14
2 49863 1 14
2 49864 1 14
2 49865 1 14
2 49866 1 14
2 49867 1 14
2 49868 1 14
2 49869 1 14
2 49870 1 14
2 49871 1 14
2 49872 1 14
2 49873 1 14
2 49874 1 14
2 49875 1 14
2 49876 1 14
2 49877 1 14
2 49878 1 14
2 49879 1 14
2 49880 1 14
2 49881 1 14
2 49882 1 14
2 49883 1 14
2 49884 1 14
2 49885 1 14
2 49886 1 14
2 49887 1 14
2 49888 1 14
2 49889 1 14
2 49890 1 14
2 49891 1 14
2 49892 1 14
2 49893 1 14
2 49894 1 14
2 49895 1 14
2 49896 1 14
2 49897 1 14
2 49898 1 14
2 49899 1 14
2 49900 1 14
2 49901 1 14
2 49902 1 14
2 49903 1 14
2 49904 1 14
2 49905 1 14
2 49906 1 14
2 49907 1 14
2 49908 1 14
2 49909 1 14
2 49910 1 14
2 49911 1 14
2 49912 1 14
2 49913 1 14
2 49914 1 14
2 49915 1 14
2 49916 1 14
2 49917 1 14
2 49918 1 14
2 49919 1 14
2 49920 1 14
2 49921 1 14
2 49922 1 14
2 49923 1 14
2 49924 1 14
2 49925 1 14
2 49926 1 14
2 49927 1 14
2 49928 1 14
2 49929 1 14
2 49930 1 14
2 49931 1 14
2 49932 1 14
2 49933 1 14
2 49934 1 14
2 49935 1 14
2 49936 1 14
2 49937 1 14
2 49938 1 14
2 49939 1 14
2 49940 1 14
2 49941 1 14
2 49942 1 14
2 49943 1 14
2 49944 1 14
2 49945 1 14
2 49946 1 14
2 49947 1 14
2 49948 1 14
2 49949 1 14
2 49950 1 14
2 49951 1 14
2 49952 1 14
2 49953 1 14
2 49954 1 14
2 49955 1 14
2 49956 1 14
2 49957 1 14
2 49958 1 14
2 49959 1 14
2 49960 1 14
2 49961 1 14
2 49962 1 14
2 49963 1 14
2 49964 1 14
2 49965 1 14
2 49966 1 14
2 49967 1 14
2 49968 1 14
2 49969 1 14
2 49970 1 14
2 49971 1 14
2 49972 1 14
2 49973 1 14
2 49974 1 14
2 49975 1 14
2 49976 1 14
2 49977 1 14
2 49978 1 14
2 49979 1 14
2 49980 1 14
2 49981 1 14
2 49982 1 14
2 49983 1 14
2 49984 1 14
2 49985 1 14
2 49986 1 14
2 49987 1 14
2 49988 1 14
2 49989 1 14
2 49990 1 14
1 15 0 84 0
2 49991 1 15
2 49992 1 15
2 49993 1 15
2 49994 1 15
2 49995 1 15
2 49996 1 15
2 49997 1 15
2 49998 1 15
2 49999 1 15
2 50000 1 15
2 50001 1 15
2 50002 1 15
2 50003 1 15
2 50004 1 15
2 50005 1 15
2 50006 1 15
2 50007 1 15
2 50008 1 15
2 50009 1 15
2 50010 1 15
2 50011 1 15
2 50012 1 15
2 50013 1 15
2 50014 1 15
2 50015 1 15
2 50016 1 15
2 50017 1 15
2 50018 1 15
2 50019 1 15
2 50020 1 15
2 50021 1 15
2 50022 1 15
2 50023 1 15
2 50024 1 15
2 50025 1 15
2 50026 1 15
2 50027 1 15
2 50028 1 15
2 50029 1 15
2 50030 1 15
2 50031 1 15
2 50032 1 15
2 50033 1 15
2 50034 1 15
2 50035 1 15
2 50036 1 15
2 50037 1 15
2 50038 1 15
2 50039 1 15
2 50040 1 15
2 50041 1 15
2 50042 1 15
2 50043 1 15
2 50044 1 15
2 50045 1 15
2 50046 1 15
2 50047 1 15
2 50048 1 15
2 50049 1 15
2 50050 1 15
2 50051 1 15
2 50052 1 15
2 50053 1 15
2 50054 1 15
2 50055 1 15
2 50056 1 15
2 50057 1 15
2 50058 1 15
2 50059 1 15
2 50060 1 15
2 50061 1 15
2 50062 1 15
2 50063 1 15
2 50064 1 15
2 50065 1 15
2 50066 1 15
2 50067 1 15
2 50068 1 15
2 50069 1 15
2 50070 1 15
2 50071 1 15
2 50072 1 15
2 50073 1 15
2 50074 1 15
1 16 0 41 0
2 50075 1 16
2 50076 1 16
2 50077 1 16
2 50078 1 16
2 50079 1 16
2 50080 1 16
2 50081 1 16
2 50082 1 16
2 50083 1 16
2 50084 1 16
2 50085 1 16
2 50086 1 16
2 50087 1 16
2 50088 1 16
2 50089 1 16
2 50090 1 16
2 50091 1 16
2 50092 1 16
2 50093 1 16
2 50094 1 16
2 50095 1 16
2 50096 1 16
2 50097 1 16
2 50098 1 16
2 50099 1 16
2 50100 1 16
2 50101 1 16
2 50102 1 16
2 50103 1 16
2 50104 1 16
2 50105 1 16
2 50106 1 16
2 50107 1 16
2 50108 1 16
2 50109 1 16
2 50110 1 16
2 50111 1 16
2 50112 1 16
2 50113 1 16
2 50114 1 16
2 50115 1 16
1 17 0 204 0
2 50116 1 17
2 50117 1 17
2 50118 1 17
2 50119 1 17
2 50120 1 17
2 50121 1 17
2 50122 1 17
2 50123 1 17
2 50124 1 17
2 50125 1 17
2 50126 1 17
2 50127 1 17
2 50128 1 17
2 50129 1 17
2 50130 1 17
2 50131 1 17
2 50132 1 17
2 50133 1 17
2 50134 1 17
2 50135 1 17
2 50136 1 17
2 50137 1 17
2 50138 1 17
2 50139 1 17
2 50140 1 17
2 50141 1 17
2 50142 1 17
2 50143 1 17
2 50144 1 17
2 50145 1 17
2 50146 1 17
2 50147 1 17
2 50148 1 17
2 50149 1 17
2 50150 1 17
2 50151 1 17
2 50152 1 17
2 50153 1 17
2 50154 1 17
2 50155 1 17
2 50156 1 17
2 50157 1 17
2 50158 1 17
2 50159 1 17
2 50160 1 17
2 50161 1 17
2 50162 1 17
2 50163 1 17
2 50164 1 17
2 50165 1 17
2 50166 1 17
2 50167 1 17
2 50168 1 17
2 50169 1 17
2 50170 1 17
2 50171 1 17
2 50172 1 17
2 50173 1 17
2 50174 1 17
2 50175 1 17
2 50176 1 17
2 50177 1 17
2 50178 1 17
2 50179 1 17
2 50180 1 17
2 50181 1 17
2 50182 1 17
2 50183 1 17
2 50184 1 17
2 50185 1 17
2 50186 1 17
2 50187 1 17
2 50188 1 17
2 50189 1 17
2 50190 1 17
2 50191 1 17
2 50192 1 17
2 50193 1 17
2 50194 1 17
2 50195 1 17
2 50196 1 17
2 50197 1 17
2 50198 1 17
2 50199 1 17
2 50200 1 17
2 50201 1 17
2 50202 1 17
2 50203 1 17
2 50204 1 17
2 50205 1 17
2 50206 1 17
2 50207 1 17
2 50208 1 17
2 50209 1 17
2 50210 1 17
2 50211 1 17
2 50212 1 17
2 50213 1 17
2 50214 1 17
2 50215 1 17
2 50216 1 17
2 50217 1 17
2 50218 1 17
2 50219 1 17
2 50220 1 17
2 50221 1 17
2 50222 1 17
2 50223 1 17
2 50224 1 17
2 50225 1 17
2 50226 1 17
2 50227 1 17
2 50228 1 17
2 50229 1 17
2 50230 1 17
2 50231 1 17
2 50232 1 17
2 50233 1 17
2 50234 1 17
2 50235 1 17
2 50236 1 17
2 50237 1 17
2 50238 1 17
2 50239 1 17
2 50240 1 17
2 50241 1 17
2 50242 1 17
2 50243 1 17
2 50244 1 17
2 50245 1 17
2 50246 1 17
2 50247 1 17
2 50248 1 17
2 50249 1 17
2 50250 1 17
2 50251 1 17
2 50252 1 17
2 50253 1 17
2 50254 1 17
2 50255 1 17
2 50256 1 17
2 50257 1 17
2 50258 1 17
2 50259 1 17
2 50260 1 17
2 50261 1 17
2 50262 1 17
2 50263 1 17
2 50264 1 17
2 50265 1 17
2 50266 1 17
2 50267 1 17
2 50268 1 17
2 50269 1 17
2 50270 1 17
2 50271 1 17
2 50272 1 17
2 50273 1 17
2 50274 1 17
2 50275 1 17
2 50276 1 17
2 50277 1 17
2 50278 1 17
2 50279 1 17
2 50280 1 17
2 50281 1 17
2 50282 1 17
2 50283 1 17
2 50284 1 17
2 50285 1 17
2 50286 1 17
2 50287 1 17
2 50288 1 17
2 50289 1 17
2 50290 1 17
2 50291 1 17
2 50292 1 17
2 50293 1 17
2 50294 1 17
2 50295 1 17
2 50296 1 17
2 50297 1 17
2 50298 1 17
2 50299 1 17
2 50300 1 17
2 50301 1 17
2 50302 1 17
2 50303 1 17
2 50304 1 17
2 50305 1 17
2 50306 1 17
2 50307 1 17
2 50308 1 17
2 50309 1 17
2 50310 1 17
2 50311 1 17
2 50312 1 17
2 50313 1 17
2 50314 1 17
2 50315 1 17
2 50316 1 17
2 50317 1 17
2 50318 1 17
2 50319 1 17
1 18 0 257 0
2 50320 1 18
2 50321 1 18
2 50322 1 18
2 50323 1 18
2 50324 1 18
2 50325 1 18
2 50326 1 18
2 50327 1 18
2 50328 1 18
2 50329 1 18
2 50330 1 18
2 50331 1 18
2 50332 1 18
2 50333 1 18
2 50334 1 18
2 50335 1 18
2 50336 1 18
2 50337 1 18
2 50338 1 18
2 50339 1 18
2 50340 1 18
2 50341 1 18
2 50342 1 18
2 50343 1 18
2 50344 1 18
2 50345 1 18
2 50346 1 18
2 50347 1 18
2 50348 1 18
2 50349 1 18
2 50350 1 18
2 50351 1 18
2 50352 1 18
2 50353 1 18
2 50354 1 18
2 50355 1 18
2 50356 1 18
2 50357 1 18
2 50358 1 18
2 50359 1 18
2 50360 1 18
2 50361 1 18
2 50362 1 18
2 50363 1 18
2 50364 1 18
2 50365 1 18
2 50366 1 18
2 50367 1 18
2 50368 1 18
2 50369 1 18
2 50370 1 18
2 50371 1 18
2 50372 1 18
2 50373 1 18
2 50374 1 18
2 50375 1 18
2 50376 1 18
2 50377 1 18
2 50378 1 18
2 50379 1 18
2 50380 1 18
2 50381 1 18
2 50382 1 18
2 50383 1 18
2 50384 1 18
2 50385 1 18
2 50386 1 18
2 50387 1 18
2 50388 1 18
2 50389 1 18
2 50390 1 18
2 50391 1 18
2 50392 1 18
2 50393 1 18
2 50394 1 18
2 50395 1 18
2 50396 1 18
2 50397 1 18
2 50398 1 18
2 50399 1 18
2 50400 1 18
2 50401 1 18
2 50402 1 18
2 50403 1 18
2 50404 1 18
2 50405 1 18
2 50406 1 18
2 50407 1 18
2 50408 1 18
2 50409 1 18
2 50410 1 18
2 50411 1 18
2 50412 1 18
2 50413 1 18
2 50414 1 18
2 50415 1 18
2 50416 1 18
2 50417 1 18
2 50418 1 18
2 50419 1 18
2 50420 1 18
2 50421 1 18
2 50422 1 18
2 50423 1 18
2 50424 1 18
2 50425 1 18
2 50426 1 18
2 50427 1 18
2 50428 1 18
2 50429 1 18
2 50430 1 18
2 50431 1 18
2 50432 1 18
2 50433 1 18
2 50434 1 18
2 50435 1 18
2 50436 1 18
2 50437 1 18
2 50438 1 18
2 50439 1 18
2 50440 1 18
2 50441 1 18
2 50442 1 18
2 50443 1 18
2 50444 1 18
2 50445 1 18
2 50446 1 18
2 50447 1 18
2 50448 1 18
2 50449 1 18
2 50450 1 18
2 50451 1 18
2 50452 1 18
2 50453 1 18
2 50454 1 18
2 50455 1 18
2 50456 1 18
2 50457 1 18
2 50458 1 18
2 50459 1 18
2 50460 1 18
2 50461 1 18
2 50462 1 18
2 50463 1 18
2 50464 1 18
2 50465 1 18
2 50466 1 18
2 50467 1 18
2 50468 1 18
2 50469 1 18
2 50470 1 18
2 50471 1 18
2 50472 1 18
2 50473 1 18
2 50474 1 18
2 50475 1 18
2 50476 1 18
2 50477 1 18
2 50478 1 18
2 50479 1 18
2 50480 1 18
2 50481 1 18
2 50482 1 18
2 50483 1 18
2 50484 1 18
2 50485 1 18
2 50486 1 18
2 50487 1 18
2 50488 1 18
2 50489 1 18
2 50490 1 18
2 50491 1 18
2 50492 1 18
2 50493 1 18
2 50494 1 18
2 50495 1 18
2 50496 1 18
2 50497 1 18
2 50498 1 18
2 50499 1 18
2 50500 1 18
2 50501 1 18
2 50502 1 18
2 50503 1 18
2 50504 1 18
2 50505 1 18
2 50506 1 18
2 50507 1 18
2 50508 1 18
2 50509 1 18
2 50510 1 18
2 50511 1 18
2 50512 1 18
2 50513 1 18
2 50514 1 18
2 50515 1 18
2 50516 1 18
2 50517 1 18
2 50518 1 18
2 50519 1 18
2 50520 1 18
2 50521 1 18
2 50522 1 18
2 50523 1 18
2 50524 1 18
2 50525 1 18
2 50526 1 18
2 50527 1 18
2 50528 1 18
2 50529 1 18
2 50530 1 18
2 50531 1 18
2 50532 1 18
2 50533 1 18
2 50534 1 18
2 50535 1 18
2 50536 1 18
2 50537 1 18
2 50538 1 18
2 50539 1 18
2 50540 1 18
2 50541 1 18
2 50542 1 18
2 50543 1 18
2 50544 1 18
2 50545 1 18
2 50546 1 18
2 50547 1 18
2 50548 1 18
2 50549 1 18
2 50550 1 18
2 50551 1 18
2 50552 1 18
2 50553 1 18
2 50554 1 18
2 50555 1 18
2 50556 1 18
2 50557 1 18
2 50558 1 18
2 50559 1 18
2 50560 1 18
2 50561 1 18
2 50562 1 18
2 50563 1 18
2 50564 1 18
2 50565 1 18
2 50566 1 18
2 50567 1 18
2 50568 1 18
2 50569 1 18
2 50570 1 18
2 50571 1 18
2 50572 1 18
2 50573 1 18
2 50574 1 18
2 50575 1 18
2 50576 1 18
1 19 0 310 0
2 50577 1 19
2 50578 1 19
2 50579 1 19
2 50580 1 19
2 50581 1 19
2 50582 1 19
2 50583 1 19
2 50584 1 19
2 50585 1 19
2 50586 1 19
2 50587 1 19
2 50588 1 19
2 50589 1 19
2 50590 1 19
2 50591 1 19
2 50592 1 19
2 50593 1 19
2 50594 1 19
2 50595 1 19
2 50596 1 19
2 50597 1 19
2 50598 1 19
2 50599 1 19
2 50600 1 19
2 50601 1 19
2 50602 1 19
2 50603 1 19
2 50604 1 19
2 50605 1 19
2 50606 1 19
2 50607 1 19
2 50608 1 19
2 50609 1 19
2 50610 1 19
2 50611 1 19
2 50612 1 19
2 50613 1 19
2 50614 1 19
2 50615 1 19
2 50616 1 19
2 50617 1 19
2 50618 1 19
2 50619 1 19
2 50620 1 19
2 50621 1 19
2 50622 1 19
2 50623 1 19
2 50624 1 19
2 50625 1 19
2 50626 1 19
2 50627 1 19
2 50628 1 19
2 50629 1 19
2 50630 1 19
2 50631 1 19
2 50632 1 19
2 50633 1 19
2 50634 1 19
2 50635 1 19
2 50636 1 19
2 50637 1 19
2 50638 1 19
2 50639 1 19
2 50640 1 19
2 50641 1 19
2 50642 1 19
2 50643 1 19
2 50644 1 19
2 50645 1 19
2 50646 1 19
2 50647 1 19
2 50648 1 19
2 50649 1 19
2 50650 1 19
2 50651 1 19
2 50652 1 19
2 50653 1 19
2 50654 1 19
2 50655 1 19
2 50656 1 19
2 50657 1 19
2 50658 1 19
2 50659 1 19
2 50660 1 19
2 50661 1 19
2 50662 1 19
2 50663 1 19
2 50664 1 19
2 50665 1 19
2 50666 1 19
2 50667 1 19
2 50668 1 19
2 50669 1 19
2 50670 1 19
2 50671 1 19
2 50672 1 19
2 50673 1 19
2 50674 1 19
2 50675 1 19
2 50676 1 19
2 50677 1 19
2 50678 1 19
2 50679 1 19
2 50680 1 19
2 50681 1 19
2 50682 1 19
2 50683 1 19
2 50684 1 19
2 50685 1 19
2 50686 1 19
2 50687 1 19
2 50688 1 19
2 50689 1 19
2 50690 1 19
2 50691 1 19
2 50692 1 19
2 50693 1 19
2 50694 1 19
2 50695 1 19
2 50696 1 19
2 50697 1 19
2 50698 1 19
2 50699 1 19
2 50700 1 19
2 50701 1 19
2 50702 1 19
2 50703 1 19
2 50704 1 19
2 50705 1 19
2 50706 1 19
2 50707 1 19
2 50708 1 19
2 50709 1 19
2 50710 1 19
2 50711 1 19
2 50712 1 19
2 50713 1 19
2 50714 1 19
2 50715 1 19
2 50716 1 19
2 50717 1 19
2 50718 1 19
2 50719 1 19
2 50720 1 19
2 50721 1 19
2 50722 1 19
2 50723 1 19
2 50724 1 19
2 50725 1 19
2 50726 1 19
2 50727 1 19
2 50728 1 19
2 50729 1 19
2 50730 1 19
2 50731 1 19
2 50732 1 19
2 50733 1 19
2 50734 1 19
2 50735 1 19
2 50736 1 19
2 50737 1 19
2 50738 1 19
2 50739 1 19
2 50740 1 19
2 50741 1 19
2 50742 1 19
2 50743 1 19
2 50744 1 19
2 50745 1 19
2 50746 1 19
2 50747 1 19
2 50748 1 19
2 50749 1 19
2 50750 1 19
2 50751 1 19
2 50752 1 19
2 50753 1 19
2 50754 1 19
2 50755 1 19
2 50756 1 19
2 50757 1 19
2 50758 1 19
2 50759 1 19
2 50760 1 19
2 50761 1 19
2 50762 1 19
2 50763 1 19
2 50764 1 19
2 50765 1 19
2 50766 1 19
2 50767 1 19
2 50768 1 19
2 50769 1 19
2 50770 1 19
2 50771 1 19
2 50772 1 19
2 50773 1 19
2 50774 1 19
2 50775 1 19
2 50776 1 19
2 50777 1 19
2 50778 1 19
2 50779 1 19
2 50780 1 19
2 50781 1 19
2 50782 1 19
2 50783 1 19
2 50784 1 19
2 50785 1 19
2 50786 1 19
2 50787 1 19
2 50788 1 19
2 50789 1 19
2 50790 1 19
2 50791 1 19
2 50792 1 19
2 50793 1 19
2 50794 1 19
2 50795 1 19
2 50796 1 19
2 50797 1 19
2 50798 1 19
2 50799 1 19
2 50800 1 19
2 50801 1 19
2 50802 1 19
2 50803 1 19
2 50804 1 19
2 50805 1 19
2 50806 1 19
2 50807 1 19
2 50808 1 19
2 50809 1 19
2 50810 1 19
2 50811 1 19
2 50812 1 19
2 50813 1 19
2 50814 1 19
2 50815 1 19
2 50816 1 19
2 50817 1 19
2 50818 1 19
2 50819 1 19
2 50820 1 19
2 50821 1 19
2 50822 1 19
2 50823 1 19
2 50824 1 19
2 50825 1 19
2 50826 1 19
2 50827 1 19
2 50828 1 19
2 50829 1 19
2 50830 1 19
2 50831 1 19
2 50832 1 19
2 50833 1 19
2 50834 1 19
2 50835 1 19
2 50836 1 19
2 50837 1 19
2 50838 1 19
2 50839 1 19
2 50840 1 19
2 50841 1 19
2 50842 1 19
2 50843 1 19
2 50844 1 19
2 50845 1 19
2 50846 1 19
2 50847 1 19
2 50848 1 19
2 50849 1 19
2 50850 1 19
2 50851 1 19
2 50852 1 19
2 50853 1 19
2 50854 1 19
2 50855 1 19
2 50856 1 19
2 50857 1 19
2 50858 1 19
2 50859 1 19
2 50860 1 19
2 50861 1 19
2 50862 1 19
2 50863 1 19
2 50864 1 19
2 50865 1 19
2 50866 1 19
2 50867 1 19
2 50868 1 19
2 50869 1 19
2 50870 1 19
2 50871 1 19
2 50872 1 19
2 50873 1 19
2 50874 1 19
2 50875 1 19
2 50876 1 19
2 50877 1 19
2 50878 1 19
2 50879 1 19
2 50880 1 19
2 50881 1 19
2 50882 1 19
2 50883 1 19
2 50884 1 19
2 50885 1 19
2 50886 1 19
1 20 0 309 0
2 50887 1 20
2 50888 1 20
2 50889 1 20
2 50890 1 20
2 50891 1 20
2 50892 1 20
2 50893 1 20
2 50894 1 20
2 50895 1 20
2 50896 1 20
2 50897 1 20
2 50898 1 20
2 50899 1 20
2 50900 1 20
2 50901 1 20
2 50902 1 20
2 50903 1 20
2 50904 1 20
2 50905 1 20
2 50906 1 20
2 50907 1 20
2 50908 1 20
2 50909 1 20
2 50910 1 20
2 50911 1 20
2 50912 1 20
2 50913 1 20
2 50914 1 20
2 50915 1 20
2 50916 1 20
2 50917 1 20
2 50918 1 20
2 50919 1 20
2 50920 1 20
2 50921 1 20
2 50922 1 20
2 50923 1 20
2 50924 1 20
2 50925 1 20
2 50926 1 20
2 50927 1 20
2 50928 1 20
2 50929 1 20
2 50930 1 20
2 50931 1 20
2 50932 1 20
2 50933 1 20
2 50934 1 20
2 50935 1 20
2 50936 1 20
2 50937 1 20
2 50938 1 20
2 50939 1 20
2 50940 1 20
2 50941 1 20
2 50942 1 20
2 50943 1 20
2 50944 1 20
2 50945 1 20
2 50946 1 20
2 50947 1 20
2 50948 1 20
2 50949 1 20
2 50950 1 20
2 50951 1 20
2 50952 1 20
2 50953 1 20
2 50954 1 20
2 50955 1 20
2 50956 1 20
2 50957 1 20
2 50958 1 20
2 50959 1 20
2 50960 1 20
2 50961 1 20
2 50962 1 20
2 50963 1 20
2 50964 1 20
2 50965 1 20
2 50966 1 20
2 50967 1 20
2 50968 1 20
2 50969 1 20
2 50970 1 20
2 50971 1 20
2 50972 1 20
2 50973 1 20
2 50974 1 20
2 50975 1 20
2 50976 1 20
2 50977 1 20
2 50978 1 20
2 50979 1 20
2 50980 1 20
2 50981 1 20
2 50982 1 20
2 50983 1 20
2 50984 1 20
2 50985 1 20
2 50986 1 20
2 50987 1 20
2 50988 1 20
2 50989 1 20
2 50990 1 20
2 50991 1 20
2 50992 1 20
2 50993 1 20
2 50994 1 20
2 50995 1 20
2 50996 1 20
2 50997 1 20
2 50998 1 20
2 50999 1 20
2 51000 1 20
2 51001 1 20
2 51002 1 20
2 51003 1 20
2 51004 1 20
2 51005 1 20
2 51006 1 20
2 51007 1 20
2 51008 1 20
2 51009 1 20
2 51010 1 20
2 51011 1 20
2 51012 1 20
2 51013 1 20
2 51014 1 20
2 51015 1 20
2 51016 1 20
2 51017 1 20
2 51018 1 20
2 51019 1 20
2 51020 1 20
2 51021 1 20
2 51022 1 20
2 51023 1 20
2 51024 1 20
2 51025 1 20
2 51026 1 20
2 51027 1 20
2 51028 1 20
2 51029 1 20
2 51030 1 20
2 51031 1 20
2 51032 1 20
2 51033 1 20
2 51034 1 20
2 51035 1 20
2 51036 1 20
2 51037 1 20
2 51038 1 20
2 51039 1 20
2 51040 1 20
2 51041 1 20
2 51042 1 20
2 51043 1 20
2 51044 1 20
2 51045 1 20
2 51046 1 20
2 51047 1 20
2 51048 1 20
2 51049 1 20
2 51050 1 20
2 51051 1 20
2 51052 1 20
2 51053 1 20
2 51054 1 20
2 51055 1 20
2 51056 1 20
2 51057 1 20
2 51058 1 20
2 51059 1 20
2 51060 1 20
2 51061 1 20
2 51062 1 20
2 51063 1 20
2 51064 1 20
2 51065 1 20
2 51066 1 20
2 51067 1 20
2 51068 1 20
2 51069 1 20
2 51070 1 20
2 51071 1 20
2 51072 1 20
2 51073 1 20
2 51074 1 20
2 51075 1 20
2 51076 1 20
2 51077 1 20
2 51078 1 20
2 51079 1 20
2 51080 1 20
2 51081 1 20
2 51082 1 20
2 51083 1 20
2 51084 1 20
2 51085 1 20
2 51086 1 20
2 51087 1 20
2 51088 1 20
2 51089 1 20
2 51090 1 20
2 51091 1 20
2 51092 1 20
2 51093 1 20
2 51094 1 20
2 51095 1 20
2 51096 1 20
2 51097 1 20
2 51098 1 20
2 51099 1 20
2 51100 1 20
2 51101 1 20
2 51102 1 20
2 51103 1 20
2 51104 1 20
2 51105 1 20
2 51106 1 20
2 51107 1 20
2 51108 1 20
2 51109 1 20
2 51110 1 20
2 51111 1 20
2 51112 1 20
2 51113 1 20
2 51114 1 20
2 51115 1 20
2 51116 1 20
2 51117 1 20
2 51118 1 20
2 51119 1 20
2 51120 1 20
2 51121 1 20
2 51122 1 20
2 51123 1 20
2 51124 1 20
2 51125 1 20
2 51126 1 20
2 51127 1 20
2 51128 1 20
2 51129 1 20
2 51130 1 20
2 51131 1 20
2 51132 1 20
2 51133 1 20
2 51134 1 20
2 51135 1 20
2 51136 1 20
2 51137 1 20
2 51138 1 20
2 51139 1 20
2 51140 1 20
2 51141 1 20
2 51142 1 20
2 51143 1 20
2 51144 1 20
2 51145 1 20
2 51146 1 20
2 51147 1 20
2 51148 1 20
2 51149 1 20
2 51150 1 20
2 51151 1 20
2 51152 1 20
2 51153 1 20
2 51154 1 20
2 51155 1 20
2 51156 1 20
2 51157 1 20
2 51158 1 20
2 51159 1 20
2 51160 1 20
2 51161 1 20
2 51162 1 20
2 51163 1 20
2 51164 1 20
2 51165 1 20
2 51166 1 20
2 51167 1 20
2 51168 1 20
2 51169 1 20
2 51170 1 20
2 51171 1 20
2 51172 1 20
2 51173 1 20
2 51174 1 20
2 51175 1 20
2 51176 1 20
2 51177 1 20
2 51178 1 20
2 51179 1 20
2 51180 1 20
2 51181 1 20
2 51182 1 20
2 51183 1 20
2 51184 1 20
2 51185 1 20
2 51186 1 20
2 51187 1 20
2 51188 1 20
2 51189 1 20
2 51190 1 20
2 51191 1 20
2 51192 1 20
2 51193 1 20
2 51194 1 20
2 51195 1 20
1 21 0 283 0
2 51196 1 21
2 51197 1 21
2 51198 1 21
2 51199 1 21
2 51200 1 21
2 51201 1 21
2 51202 1 21
2 51203 1 21
2 51204 1 21
2 51205 1 21
2 51206 1 21
2 51207 1 21
2 51208 1 21
2 51209 1 21
2 51210 1 21
2 51211 1 21
2 51212 1 21
2 51213 1 21
2 51214 1 21
2 51215 1 21
2 51216 1 21
2 51217 1 21
2 51218 1 21
2 51219 1 21
2 51220 1 21
2 51221 1 21
2 51222 1 21
2 51223 1 21
2 51224 1 21
2 51225 1 21
2 51226 1 21
2 51227 1 21
2 51228 1 21
2 51229 1 21
2 51230 1 21
2 51231 1 21
2 51232 1 21
2 51233 1 21
2 51234 1 21
2 51235 1 21
2 51236 1 21
2 51237 1 21
2 51238 1 21
2 51239 1 21
2 51240 1 21
2 51241 1 21
2 51242 1 21
2 51243 1 21
2 51244 1 21
2 51245 1 21
2 51246 1 21
2 51247 1 21
2 51248 1 21
2 51249 1 21
2 51250 1 21
2 51251 1 21
2 51252 1 21
2 51253 1 21
2 51254 1 21
2 51255 1 21
2 51256 1 21
2 51257 1 21
2 51258 1 21
2 51259 1 21
2 51260 1 21
2 51261 1 21
2 51262 1 21
2 51263 1 21
2 51264 1 21
2 51265 1 21
2 51266 1 21
2 51267 1 21
2 51268 1 21
2 51269 1 21
2 51270 1 21
2 51271 1 21
2 51272 1 21
2 51273 1 21
2 51274 1 21
2 51275 1 21
2 51276 1 21
2 51277 1 21
2 51278 1 21
2 51279 1 21
2 51280 1 21
2 51281 1 21
2 51282 1 21
2 51283 1 21
2 51284 1 21
2 51285 1 21
2 51286 1 21
2 51287 1 21
2 51288 1 21
2 51289 1 21
2 51290 1 21
2 51291 1 21
2 51292 1 21
2 51293 1 21
2 51294 1 21
2 51295 1 21
2 51296 1 21
2 51297 1 21
2 51298 1 21
2 51299 1 21
2 51300 1 21
2 51301 1 21
2 51302 1 21
2 51303 1 21
2 51304 1 21
2 51305 1 21
2 51306 1 21
2 51307 1 21
2 51308 1 21
2 51309 1 21
2 51310 1 21
2 51311 1 21
2 51312 1 21
2 51313 1 21
2 51314 1 21
2 51315 1 21
2 51316 1 21
2 51317 1 21
2 51318 1 21
2 51319 1 21
2 51320 1 21
2 51321 1 21
2 51322 1 21
2 51323 1 21
2 51324 1 21
2 51325 1 21
2 51326 1 21
2 51327 1 21
2 51328 1 21
2 51329 1 21
2 51330 1 21
2 51331 1 21
2 51332 1 21
2 51333 1 21
2 51334 1 21
2 51335 1 21
2 51336 1 21
2 51337 1 21
2 51338 1 21
2 51339 1 21
2 51340 1 21
2 51341 1 21
2 51342 1 21
2 51343 1 21
2 51344 1 21
2 51345 1 21
2 51346 1 21
2 51347 1 21
2 51348 1 21
2 51349 1 21
2 51350 1 21
2 51351 1 21
2 51352 1 21
2 51353 1 21
2 51354 1 21
2 51355 1 21
2 51356 1 21
2 51357 1 21
2 51358 1 21
2 51359 1 21
2 51360 1 21
2 51361 1 21
2 51362 1 21
2 51363 1 21
2 51364 1 21
2 51365 1 21
2 51366 1 21
2 51367 1 21
2 51368 1 21
2 51369 1 21
2 51370 1 21
2 51371 1 21
2 51372 1 21
2 51373 1 21
2 51374 1 21
2 51375 1 21
2 51376 1 21
2 51377 1 21
2 51378 1 21
2 51379 1 21
2 51380 1 21
2 51381 1 21
2 51382 1 21
2 51383 1 21
2 51384 1 21
2 51385 1 21
2 51386 1 21
2 51387 1 21
2 51388 1 21
2 51389 1 21
2 51390 1 21
2 51391 1 21
2 51392 1 21
2 51393 1 21
2 51394 1 21
2 51395 1 21
2 51396 1 21
2 51397 1 21
2 51398 1 21
2 51399 1 21
2 51400 1 21
2 51401 1 21
2 51402 1 21
2 51403 1 21
2 51404 1 21
2 51405 1 21
2 51406 1 21
2 51407 1 21
2 51408 1 21
2 51409 1 21
2 51410 1 21
2 51411 1 21
2 51412 1 21
2 51413 1 21
2 51414 1 21
2 51415 1 21
2 51416 1 21
2 51417 1 21
2 51418 1 21
2 51419 1 21
2 51420 1 21
2 51421 1 21
2 51422 1 21
2 51423 1 21
2 51424 1 21
2 51425 1 21
2 51426 1 21
2 51427 1 21
2 51428 1 21
2 51429 1 21
2 51430 1 21
2 51431 1 21
2 51432 1 21
2 51433 1 21
2 51434 1 21
2 51435 1 21
2 51436 1 21
2 51437 1 21
2 51438 1 21
2 51439 1 21
2 51440 1 21
2 51441 1 21
2 51442 1 21
2 51443 1 21
2 51444 1 21
2 51445 1 21
2 51446 1 21
2 51447 1 21
2 51448 1 21
2 51449 1 21
2 51450 1 21
2 51451 1 21
2 51452 1 21
2 51453 1 21
2 51454 1 21
2 51455 1 21
2 51456 1 21
2 51457 1 21
2 51458 1 21
2 51459 1 21
2 51460 1 21
2 51461 1 21
2 51462 1 21
2 51463 1 21
2 51464 1 21
2 51465 1 21
2 51466 1 21
2 51467 1 21
2 51468 1 21
2 51469 1 21
2 51470 1 21
2 51471 1 21
2 51472 1 21
2 51473 1 21
2 51474 1 21
2 51475 1 21
2 51476 1 21
2 51477 1 21
2 51478 1 21
1 22 0 203 0
2 51479 1 22
2 51480 1 22
2 51481 1 22
2 51482 1 22
2 51483 1 22
2 51484 1 22
2 51485 1 22
2 51486 1 22
2 51487 1 22
2 51488 1 22
2 51489 1 22
2 51490 1 22
2 51491 1 22
2 51492 1 22
2 51493 1 22
2 51494 1 22
2 51495 1 22
2 51496 1 22
2 51497 1 22
2 51498 1 22
2 51499 1 22
2 51500 1 22
2 51501 1 22
2 51502 1 22
2 51503 1 22
2 51504 1 22
2 51505 1 22
2 51506 1 22
2 51507 1 22
2 51508 1 22
2 51509 1 22
2 51510 1 22
2 51511 1 22
2 51512 1 22
2 51513 1 22
2 51514 1 22
2 51515 1 22
2 51516 1 22
2 51517 1 22
2 51518 1 22
2 51519 1 22
2 51520 1 22
2 51521 1 22
2 51522 1 22
2 51523 1 22
2 51524 1 22
2 51525 1 22
2 51526 1 22
2 51527 1 22
2 51528 1 22
2 51529 1 22
2 51530 1 22
2 51531 1 22
2 51532 1 22
2 51533 1 22
2 51534 1 22
2 51535 1 22
2 51536 1 22
2 51537 1 22
2 51538 1 22
2 51539 1 22
2 51540 1 22
2 51541 1 22
2 51542 1 22
2 51543 1 22
2 51544 1 22
2 51545 1 22
2 51546 1 22
2 51547 1 22
2 51548 1 22
2 51549 1 22
2 51550 1 22
2 51551 1 22
2 51552 1 22
2 51553 1 22
2 51554 1 22
2 51555 1 22
2 51556 1 22
2 51557 1 22
2 51558 1 22
2 51559 1 22
2 51560 1 22
2 51561 1 22
2 51562 1 22
2 51563 1 22
2 51564 1 22
2 51565 1 22
2 51566 1 22
2 51567 1 22
2 51568 1 22
2 51569 1 22
2 51570 1 22
2 51571 1 22
2 51572 1 22
2 51573 1 22
2 51574 1 22
2 51575 1 22
2 51576 1 22
2 51577 1 22
2 51578 1 22
2 51579 1 22
2 51580 1 22
2 51581 1 22
2 51582 1 22
2 51583 1 22
2 51584 1 22
2 51585 1 22
2 51586 1 22
2 51587 1 22
2 51588 1 22
2 51589 1 22
2 51590 1 22
2 51591 1 22
2 51592 1 22
2 51593 1 22
2 51594 1 22
2 51595 1 22
2 51596 1 22
2 51597 1 22
2 51598 1 22
2 51599 1 22
2 51600 1 22
2 51601 1 22
2 51602 1 22
2 51603 1 22
2 51604 1 22
2 51605 1 22
2 51606 1 22
2 51607 1 22
2 51608 1 22
2 51609 1 22
2 51610 1 22
2 51611 1 22
2 51612 1 22
2 51613 1 22
2 51614 1 22
2 51615 1 22
2 51616 1 22
2 51617 1 22
2 51618 1 22
2 51619 1 22
2 51620 1 22
2 51621 1 22
2 51622 1 22
2 51623 1 22
2 51624 1 22
2 51625 1 22
2 51626 1 22
2 51627 1 22
2 51628 1 22
2 51629 1 22
2 51630 1 22
2 51631 1 22
2 51632 1 22
2 51633 1 22
2 51634 1 22
2 51635 1 22
2 51636 1 22
2 51637 1 22
2 51638 1 22
2 51639 1 22
2 51640 1 22
2 51641 1 22
2 51642 1 22
2 51643 1 22
2 51644 1 22
2 51645 1 22
2 51646 1 22
2 51647 1 22
2 51648 1 22
2 51649 1 22
2 51650 1 22
2 51651 1 22
2 51652 1 22
2 51653 1 22
2 51654 1 22
2 51655 1 22
2 51656 1 22
2 51657 1 22
2 51658 1 22
2 51659 1 22
2 51660 1 22
2 51661 1 22
2 51662 1 22
2 51663 1 22
2 51664 1 22
2 51665 1 22
2 51666 1 22
2 51667 1 22
2 51668 1 22
2 51669 1 22
2 51670 1 22
2 51671 1 22
2 51672 1 22
2 51673 1 22
2 51674 1 22
2 51675 1 22
2 51676 1 22
2 51677 1 22
2 51678 1 22
2 51679 1 22
2 51680 1 22
2 51681 1 22
1 23 0 147 0
2 51682 1 23
2 51683 1 23
2 51684 1 23
2 51685 1 23
2 51686 1 23
2 51687 1 23
2 51688 1 23
2 51689 1 23
2 51690 1 23
2 51691 1 23
2 51692 1 23
2 51693 1 23
2 51694 1 23
2 51695 1 23
2 51696 1 23
2 51697 1 23
2 51698 1 23
2 51699 1 23
2 51700 1 23
2 51701 1 23
2 51702 1 23
2 51703 1 23
2 51704 1 23
2 51705 1 23
2 51706 1 23
2 51707 1 23
2 51708 1 23
2 51709 1 23
2 51710 1 23
2 51711 1 23
2 51712 1 23
2 51713 1 23
2 51714 1 23
2 51715 1 23
2 51716 1 23
2 51717 1 23
2 51718 1 23
2 51719 1 23
2 51720 1 23
2 51721 1 23
2 51722 1 23
2 51723 1 23
2 51724 1 23
2 51725 1 23
2 51726 1 23
2 51727 1 23
2 51728 1 23
2 51729 1 23
2 51730 1 23
2 51731 1 23
2 51732 1 23
2 51733 1 23
2 51734 1 23
2 51735 1 23
2 51736 1 23
2 51737 1 23
2 51738 1 23
2 51739 1 23
2 51740 1 23
2 51741 1 23
2 51742 1 23
2 51743 1 23
2 51744 1 23
2 51745 1 23
2 51746 1 23
2 51747 1 23
2 51748 1 23
2 51749 1 23
2 51750 1 23
2 51751 1 23
2 51752 1 23
2 51753 1 23
2 51754 1 23
2 51755 1 23
2 51756 1 23
2 51757 1 23
2 51758 1 23
2 51759 1 23
2 51760 1 23
2 51761 1 23
2 51762 1 23
2 51763 1 23
2 51764 1 23
2 51765 1 23
2 51766 1 23
2 51767 1 23
2 51768 1 23
2 51769 1 23
2 51770 1 23
2 51771 1 23
2 51772 1 23
2 51773 1 23
2 51774 1 23
2 51775 1 23
2 51776 1 23
2 51777 1 23
2 51778 1 23
2 51779 1 23
2 51780 1 23
2 51781 1 23
2 51782 1 23
2 51783 1 23
2 51784 1 23
2 51785 1 23
2 51786 1 23
2 51787 1 23
2 51788 1 23
2 51789 1 23
2 51790 1 23
2 51791 1 23
2 51792 1 23
2 51793 1 23
2 51794 1 23
2 51795 1 23
2 51796 1 23
2 51797 1 23
2 51798 1 23
2 51799 1 23
2 51800 1 23
2 51801 1 23
2 51802 1 23
2 51803 1 23
2 51804 1 23
2 51805 1 23
2 51806 1 23
2 51807 1 23
2 51808 1 23
2 51809 1 23
2 51810 1 23
2 51811 1 23
2 51812 1 23
2 51813 1 23
2 51814 1 23
2 51815 1 23
2 51816 1 23
2 51817 1 23
2 51818 1 23
2 51819 1 23
2 51820 1 23
2 51821 1 23
2 51822 1 23
2 51823 1 23
2 51824 1 23
2 51825 1 23
2 51826 1 23
2 51827 1 23
2 51828 1 23
1 24 0 2 0
2 51829 1 24
2 51830 1 24
2 51831 1 27
2 51832 1 27
2 51833 1 27
2 51834 1 27
2 51835 1 27
2 51836 1 27
2 51837 1 27
2 51838 1 27
2 51839 1 27
2 51840 1 27
2 51841 1 27
2 51842 1 27
2 51843 1 27
2 51844 1 27
2 51845 1 27
2 51846 1 27
2 51847 1 27
2 51848 1 27
2 51849 1 27
2 51850 1 27
2 51851 1 27
2 51852 1 27
2 51853 1 27
2 51854 1 27
2 51855 1 27
2 51856 1 27
2 51857 1 27
2 51858 1 27
2 51859 1 27
2 51860 1 27
2 51861 1 27
2 51862 1 27
2 51863 1 27
2 51864 1 27
2 51865 1 27
2 51866 1 27
2 51867 1 27
2 51868 1 27
2 51869 1 27
2 51870 1 27
2 51871 1 27
2 51872 1 27
2 51873 1 27
2 51874 1 27
2 51875 1 27
2 51876 1 27
2 51877 1 27
2 51878 1 27
2 51879 1 27
2 51880 1 27
2 51881 1 27
2 51882 1 27
2 51883 1 27
2 51884 1 27
2 51885 1 27
2 51886 1 27
2 51887 1 27
2 51888 1 27
2 51889 1 27
2 51890 1 27
2 51891 1 27
2 51892 1 27
2 51893 1 27
2 51894 1 27
2 51895 1 27
2 51896 1 27
2 51897 1 27
2 51898 1 27
2 51899 1 27
2 51900 1 27
2 51901 1 27
2 51902 1 27
2 51903 1 27
2 51904 1 27
2 51905 1 27
2 51906 1 27
2 51907 1 27
2 51908 1 27
2 51909 1 27
2 51910 1 27
2 51911 1 27
2 51912 1 27
2 51913 1 27
2 51914 1 27
2 51915 1 27
2 51916 1 27
2 51917 1 27
2 51918 1 27
2 51919 1 27
2 51920 1 27
2 51921 1 27
2 51922 1 27
2 51923 1 27
2 51924 1 27
2 51925 1 27
2 51926 1 27
2 51927 1 27
2 51928 1 27
2 51929 1 27
2 51930 1 27
2 51931 1 27
2 51932 1 27
2 51933 1 27
2 51934 1 27
2 51935 1 27
2 51936 1 27
2 51937 1 27
2 51938 1 27
2 51939 1 27
2 51940 1 27
2 51941 1 27
2 51942 1 27
2 51943 1 27
2 51944 1 27
2 51945 1 27
2 51946 1 27
2 51947 1 27
2 51948 1 27
2 51949 1 27
2 51950 1 27
2 51951 1 27
2 51952 1 27
2 51953 1 27
2 51954 1 27
2 51955 1 27
2 51956 1 27
2 51957 1 27
2 51958 1 27
2 51959 1 27
2 51960 1 27
2 51961 1 27
2 51962 1 27
2 51963 1 27
2 51964 1 27
2 51965 1 27
2 51966 1 27
2 51967 1 27
2 51968 1 27
2 51969 1 27
2 51970 1 27
2 51971 1 27
2 51972 1 27
2 51973 1 27
2 51974 1 27
2 51975 1 27
2 51976 1 27
2 51977 1 27
2 51978 1 27
2 51979 1 27
2 51980 1 27
2 51981 1 27
2 51982 1 27
2 51983 1 27
2 51984 1 27
2 51985 1 27
2 51986 1 27
2 51987 1 27
2 51988 1 27
2 51989 1 27
2 51990 1 27
2 51991 1 27
2 51992 1 27
2 51993 1 27
2 51994 1 27
2 51995 1 27
2 51996 1 27
2 51997 1 27
2 51998 1 27
2 51999 1 27
2 52000 1 27
2 52001 1 27
2 52002 1 27
2 52003 1 27
2 52004 1 27
2 52005 1 27
2 52006 1 27
2 52007 1 27
2 52008 1 27
2 52009 1 27
2 52010 1 27
2 52011 1 27
2 52012 1 27
2 52013 1 27
2 52014 1 27
2 52015 1 27
2 52016 1 27
2 52017 1 27
2 52018 1 27
2 52019 1 27
2 52020 1 27
2 52021 1 27
2 52022 1 27
2 52023 1 27
2 52024 1 27
2 52025 1 27
2 52026 1 27
2 52027 1 27
2 52028 1 27
2 52029 1 27
2 52030 1 27
2 52031 1 27
2 52032 1 27
2 52033 1 27
2 52034 1 27
2 52035 1 27
2 52036 1 27
2 52037 1 27
2 52038 1 27
2 52039 1 27
2 52040 1 27
2 52041 1 27
2 52042 1 27
2 52043 1 27
2 52044 1 27
2 52045 1 28
2 52046 1 28
2 52047 1 28
2 52048 1 28
2 52049 1 28
2 52050 1 28
2 52051 1 28
2 52052 1 28
2 52053 1 28
2 52054 1 28
2 52055 1 28
2 52056 1 28
2 52057 1 28
2 52058 1 28
2 52059 1 28
2 52060 1 28
2 52061 1 28
2 52062 1 28
2 52063 1 28
2 52064 1 28
2 52065 1 28
2 52066 1 28
2 52067 1 28
2 52068 1 28
2 52069 1 28
2 52070 1 28
2 52071 1 28
2 52072 1 28
2 52073 1 28
2 52074 1 28
2 52075 1 28
2 52076 1 28
2 52077 1 28
2 52078 1 28
2 52079 1 28
2 52080 1 28
2 52081 1 28
2 52082 1 28
2 52083 1 28
2 52084 1 28
2 52085 1 28
2 52086 1 28
2 52087 1 28
2 52088 1 28
2 52089 1 28
2 52090 1 28
2 52091 1 28
2 52092 1 28
2 52093 1 28
2 52094 1 28
2 52095 1 28
2 52096 1 28
2 52097 1 28
2 52098 1 28
2 52099 1 28
2 52100 1 28
2 52101 1 28
2 52102 1 28
2 52103 1 28
2 52104 1 28
2 52105 1 28
2 52106 1 28
2 52107 1 28
2 52108 1 28
2 52109 1 28
2 52110 1 28
2 52111 1 28
2 52112 1 28
2 52113 1 28
2 52114 1 28
2 52115 1 28
2 52116 1 28
2 52117 1 28
2 52118 1 28
2 52119 1 28
2 52120 1 28
2 52121 1 28
2 52122 1 28
2 52123 1 28
2 52124 1 28
2 52125 1 28
2 52126 1 28
2 52127 1 28
2 52128 1 28
2 52129 1 28
2 52130 1 28
2 52131 1 28
2 52132 1 28
2 52133 1 28
2 52134 1 28
2 52135 1 28
2 52136 1 28
2 52137 1 28
2 52138 1 28
2 52139 1 28
2 52140 1 28
2 52141 1 28
2 52142 1 28
2 52143 1 28
2 52144 1 28
2 52145 1 28
2 52146 1 28
2 52147 1 28
2 52148 1 28
2 52149 1 28
2 52150 1 28
2 52151 1 28
2 52152 1 28
2 52153 1 28
2 52154 1 28
2 52155 1 28
2 52156 1 28
2 52157 1 28
2 52158 1 28
2 52159 1 28
2 52160 1 28
2 52161 1 28
2 52162 1 28
2 52163 1 28
2 52164 1 28
2 52165 1 28
2 52166 1 28
2 52167 1 28
2 52168 1 28
2 52169 1 28
2 52170 1 28
2 52171 1 28
2 52172 1 28
2 52173 1 28
2 52174 1 28
2 52175 1 28
2 52176 1 28
2 52177 1 28
2 52178 1 28
2 52179 1 28
2 52180 1 28
2 52181 1 28
2 52182 1 28
2 52183 1 28
2 52184 1 28
2 52185 1 28
2 52186 1 28
2 52187 1 28
2 52188 1 28
2 52189 1 28
2 52190 1 28
2 52191 1 28
2 52192 1 28
2 52193 1 28
2 52194 1 28
2 52195 1 28
2 52196 1 28
2 52197 1 28
2 52198 1 28
2 52199 1 28
2 52200 1 28
2 52201 1 28
2 52202 1 28
2 52203 1 28
2 52204 1 28
2 52205 1 28
2 52206 1 28
2 52207 1 28
2 52208 1 28
2 52209 1 28
2 52210 1 28
2 52211 1 28
2 52212 1 29
2 52213 1 29
2 52214 1 29
2 52215 1 29
2 52216 1 29
2 52217 1 29
2 52218 1 29
2 52219 1 29
2 52220 1 29
2 52221 1 29
2 52222 1 29
2 52223 1 29
2 52224 1 29
2 52225 1 29
2 52226 1 29
2 52227 1 29
2 52228 1 29
2 52229 1 29
2 52230 1 29
2 52231 1 29
2 52232 1 29
2 52233 1 29
2 52234 1 29
2 52235 1 29
2 52236 1 29
2 52237 1 29
2 52238 1 29
2 52239 1 29
2 52240 1 29
2 52241 1 29
2 52242 1 29
2 52243 1 29
2 52244 1 29
2 52245 1 29
2 52246 1 29
2 52247 1 29
2 52248 1 29
2 52249 1 29
2 52250 1 29
2 52251 1 29
2 52252 1 29
2 52253 1 29
2 52254 1 29
2 52255 1 29
2 52256 1 29
2 52257 1 29
2 52258 1 29
2 52259 1 29
2 52260 1 29
2 52261 1 29
2 52262 1 29
2 52263 1 29
2 52264 1 29
2 52265 1 29
2 52266 1 29
2 52267 1 29
2 52268 1 29
2 52269 1 29
2 52270 1 29
2 52271 1 29
2 52272 1 29
2 52273 1 29
2 52274 1 29
2 52275 1 29
2 52276 1 29
2 52277 1 29
2 52278 1 29
2 52279 1 29
2 52280 1 29
2 52281 1 29
2 52282 1 29
2 52283 1 29
2 52284 1 29
2 52285 1 29
2 52286 1 29
2 52287 1 29
2 52288 1 29
2 52289 1 29
2 52290 1 29
2 52291 1 29
2 52292 1 29
2 52293 1 29
2 52294 1 29
2 52295 1 29
2 52296 1 29
2 52297 1 29
2 52298 1 29
2 52299 1 29
2 52300 1 29
2 52301 1 29
2 52302 1 29
2 52303 1 29
2 52304 1 29
2 52305 1 29
2 52306 1 29
2 52307 1 29
2 52308 1 29
2 52309 1 29
2 52310 1 29
2 52311 1 29
2 52312 1 29
2 52313 1 29
2 52314 1 29
2 52315 1 29
2 52316 1 29
2 52317 1 29
2 52318 1 29
2 52319 1 29
2 52320 1 29
2 52321 1 29
2 52322 1 29
2 52323 1 29
2 52324 1 29
2 52325 1 29
2 52326 1 29
2 52327 1 29
2 52328 1 29
2 52329 1 29
2 52330 1 29
2 52331 1 29
2 52332 1 29
2 52333 1 29
2 52334 1 29
2 52335 1 29
2 52336 1 29
2 52337 1 29
2 52338 1 29
2 52339 1 29
2 52340 1 29
2 52341 1 29
2 52342 1 29
2 52343 1 29
2 52344 1 29
2 52345 1 29
2 52346 1 29
2 52347 1 29
2 52348 1 29
2 52349 1 29
2 52350 1 29
2 52351 1 29
2 52352 1 29
2 52353 1 29
2 52354 1 29
2 52355 1 29
2 52356 1 29
2 52357 1 29
2 52358 1 29
2 52359 1 29
2 52360 1 30
2 52361 1 30
2 52362 1 30
2 52363 1 30
2 52364 1 30
2 52365 1 30
2 52366 1 30
2 52367 1 30
2 52368 1 30
2 52369 1 30
2 52370 1 30
2 52371 1 30
2 52372 1 30
2 52373 1 30
2 52374 1 30
2 52375 1 30
2 52376 1 30
2 52377 1 30
2 52378 1 30
2 52379 1 30
2 52380 1 30
2 52381 1 30
2 52382 1 30
2 52383 1 30
2 52384 1 30
2 52385 1 30
2 52386 1 30
2 52387 1 30
2 52388 1 30
2 52389 1 30
2 52390 1 30
2 52391 1 30
2 52392 1 30
2 52393 1 30
2 52394 1 30
2 52395 1 30
2 52396 1 30
2 52397 1 30
2 52398 1 30
2 52399 1 30
2 52400 1 30
2 52401 1 30
2 52402 1 30
2 52403 1 30
2 52404 1 30
2 52405 1 30
2 52406 1 30
2 52407 1 30
2 52408 1 30
2 52409 1 30
2 52410 1 30
2 52411 1 30
2 52412 1 30
2 52413 1 30
2 52414 1 30
2 52415 1 30
2 52416 1 30
2 52417 1 30
2 52418 1 30
2 52419 1 30
2 52420 1 30
2 52421 1 30
2 52422 1 30
2 52423 1 30
2 52424 1 30
2 52425 1 30
2 52426 1 30
2 52427 1 30
2 52428 1 30
2 52429 1 30
2 52430 1 30
2 52431 1 30
2 52432 1 30
2 52433 1 30
2 52434 1 30
2 52435 1 30
2 52436 1 30
2 52437 1 30
2 52438 1 30
2 52439 1 30
2 52440 1 30
2 52441 1 30
2 52442 1 30
2 52443 1 30
2 52444 1 30
2 52445 1 30
2 52446 1 30
2 52447 1 30
2 52448 1 30
2 52449 1 30
2 52450 1 30
2 52451 1 30
2 52452 1 30
2 52453 1 30
2 52454 1 30
2 52455 1 30
2 52456 1 30
2 52457 1 30
2 52458 1 30
2 52459 1 30
2 52460 1 30
2 52461 1 30
2 52462 1 30
2 52463 1 30
2 52464 1 30
2 52465 1 30
2 52466 1 30
2 52467 1 30
2 52468 1 30
2 52469 1 30
2 52470 1 31
2 52471 1 31
2 52472 1 31
2 52473 1 31
2 52474 1 31
2 52475 1 31
2 52476 1 31
2 52477 1 31
2 52478 1 31
2 52479 1 31
2 52480 1 31
2 52481 1 31
2 52482 1 31
2 52483 1 31
2 52484 1 31
2 52485 1 31
2 52486 1 31
2 52487 1 31
2 52488 1 31
2 52489 1 31
2 52490 1 31
2 52491 1 31
2 52492 1 31
2 52493 1 31
2 52494 1 31
2 52495 1 31
2 52496 1 31
2 52497 1 31
2 52498 1 31
2 52499 1 31
2 52500 1 31
2 52501 1 31
2 52502 1 31
2 52503 1 31
2 52504 1 31
2 52505 1 31
2 52506 1 31
2 52507 1 31
2 52508 1 31
2 52509 1 31
2 52510 1 31
2 52511 1 31
2 52512 1 31
2 52513 1 31
2 52514 1 31
2 52515 1 31
2 52516 1 31
2 52517 1 31
2 52518 1 31
2 52519 1 31
2 52520 1 31
2 52521 1 31
2 52522 1 31
2 52523 1 31
2 52524 1 31
2 52525 1 31
2 52526 1 31
2 52527 1 31
2 52528 1 31
2 52529 1 31
2 52530 1 31
2 52531 1 31
2 52532 1 31
2 52533 1 31
2 52534 1 31
2 52535 1 31
2 52536 1 31
2 52537 1 31
2 52538 1 31
2 52539 1 31
2 52540 1 31
2 52541 1 31
2 52542 1 31
2 52543 1 31
2 52544 1 31
2 52545 1 31
2 52546 1 31
2 52547 1 31
2 52548 1 31
2 52549 1 31
2 52550 1 31
2 52551 1 31
2 52552 1 31
2 52553 1 31
2 52554 1 31
2 52555 1 31
2 52556 1 31
2 52557 1 31
2 52558 1 31
2 52559 1 31
2 52560 1 31
2 52561 1 31
2 52562 1 31
2 52563 1 31
2 52564 1 31
2 52565 1 31
2 52566 1 31
2 52567 1 31
2 52568 1 31
2 52569 1 31
2 52570 1 31
2 52571 1 31
2 52572 1 31
2 52573 1 31
2 52574 1 31
2 52575 1 31
2 52576 1 31
2 52577 1 31
2 52578 1 31
2 52579 1 31
2 52580 1 31
2 52581 1 31
2 52582 1 31
2 52583 1 31
2 52584 1 31
2 52585 1 31
2 52586 1 32
2 52587 1 32
2 52588 1 32
2 52589 1 32
2 52590 1 32
2 52591 1 32
2 52592 1 32
2 52593 1 32
2 52594 1 32
2 52595 1 32
2 52596 1 32
2 52597 1 32
2 52598 1 32
2 52599 1 32
2 52600 1 32
2 52601 1 32
2 52602 1 32
2 52603 1 32
2 52604 1 32
2 52605 1 32
2 52606 1 32
2 52607 1 32
2 52608 1 32
2 52609 1 32
2 52610 1 32
2 52611 1 32
2 52612 1 32
2 52613 1 32
2 52614 1 32
2 52615 1 32
2 52616 1 32
2 52617 1 32
2 52618 1 32
2 52619 1 32
2 52620 1 32
2 52621 1 32
2 52622 1 32
2 52623 1 32
2 52624 1 32
2 52625 1 32
2 52626 1 32
2 52627 1 32
2 52628 1 32
2 52629 1 32
2 52630 1 32
2 52631 1 32
2 52632 1 32
2 52633 1 32
2 52634 1 32
2 52635 1 32
2 52636 1 32
2 52637 1 32
2 52638 1 32
2 52639 1 32
2 52640 1 32
2 52641 1 32
2 52642 1 32
2 52643 1 32
2 52644 1 32
2 52645 1 32
2 52646 1 32
2 52647 1 32
2 52648 1 32
2 52649 1 32
2 52650 1 32
2 52651 1 32
2 52652 1 32
2 52653 1 32
2 52654 1 32
2 52655 1 32
2 52656 1 32
2 52657 1 32
2 52658 1 32
2 52659 1 32
2 52660 1 32
2 52661 1 32
2 52662 1 32
2 52663 1 32
2 52664 1 32
2 52665 1 32
2 52666 1 32
2 52667 1 32
2 52668 1 32
2 52669 1 32
2 52670 1 32
2 52671 1 32
2 52672 1 32
2 52673 1 32
2 52674 1 32
2 52675 1 32
2 52676 1 32
2 52677 1 32
2 52678 1 32
2 52679 1 32
2 52680 1 32
2 52681 1 32
2 52682 1 32
2 52683 1 32
2 52684 1 32
2 52685 1 32
2 52686 1 32
2 52687 1 32
2 52688 1 32
2 52689 1 32
2 52690 1 32
2 52691 1 32
2 52692 1 32
2 52693 1 32
2 52694 1 32
2 52695 1 32
2 52696 1 32
2 52697 1 32
2 52698 1 32
2 52699 1 32
2 52700 1 32
2 52701 1 32
2 52702 1 32
2 52703 1 32
2 52704 1 32
2 52705 1 32
2 52706 1 32
2 52707 1 32
2 52708 1 32
2 52709 1 32
2 52710 1 32
2 52711 1 32
2 52712 1 32
2 52713 1 32
2 52714 1 32
2 52715 1 32
2 52716 1 32
2 52717 1 32
2 52718 1 32
2 52719 1 32
2 52720 1 32
2 52721 1 32
2 52722 1 32
2 52723 1 32
2 52724 1 32
2 52725 1 32
2 52726 1 32
2 52727 1 32
2 52728 1 32
2 52729 1 32
2 52730 1 32
2 52731 1 32
2 52732 1 32
2 52733 1 32
2 52734 1 32
2 52735 1 32
2 52736 1 32
2 52737 1 32
2 52738 1 32
2 52739 1 32
2 52740 1 32
2 52741 1 33
2 52742 1 33
2 52743 1 33
2 52744 1 33
2 52745 1 33
2 52746 1 33
2 52747 1 33
2 52748 1 33
2 52749 1 33
2 52750 1 33
2 52751 1 33
2 52752 1 33
2 52753 1 33
2 52754 1 33
2 52755 1 33
2 52756 1 33
2 52757 1 33
2 52758 1 33
2 52759 1 33
2 52760 1 33
2 52761 1 33
2 52762 1 33
2 52763 1 33
2 52764 1 33
2 52765 1 33
2 52766 1 33
2 52767 1 33
2 52768 1 33
2 52769 1 33
2 52770 1 33
2 52771 1 33
2 52772 1 33
2 52773 1 33
2 52774 1 33
2 52775 1 33
2 52776 1 33
2 52777 1 33
2 52778 1 33
2 52779 1 33
2 52780 1 33
2 52781 1 33
2 52782 1 33
2 52783 1 33
2 52784 1 33
2 52785 1 33
2 52786 1 33
2 52787 1 33
2 52788 1 33
2 52789 1 33
2 52790 1 33
2 52791 1 33
2 52792 1 33
2 52793 1 33
2 52794 1 33
2 52795 1 33
2 52796 1 33
2 52797 1 33
2 52798 1 33
2 52799 1 33
2 52800 1 33
2 52801 1 33
2 52802 1 33
2 52803 1 33
2 52804 1 33
2 52805 1 33
2 52806 1 33
2 52807 1 33
2 52808 1 33
2 52809 1 33
2 52810 1 33
2 52811 1 33
2 52812 1 33
2 52813 1 33
2 52814 1 33
2 52815 1 33
2 52816 1 33
2 52817 1 33
2 52818 1 33
2 52819 1 33
2 52820 1 33
2 52821 1 33
2 52822 1 33
2 52823 1 33
2 52824 1 33
2 52825 1 33
2 52826 1 33
2 52827 1 33
2 52828 1 33
2 52829 1 33
2 52830 1 33
2 52831 1 33
2 52832 1 33
2 52833 1 33
2 52834 1 33
2 52835 1 33
2 52836 1 33
2 52837 1 33
2 52838 1 33
2 52839 1 33
2 52840 1 33
2 52841 1 33
2 52842 1 33
2 52843 1 33
2 52844 1 33
2 52845 1 33
2 52846 1 33
2 52847 1 33
2 52848 1 33
2 52849 1 33
2 52850 1 33
2 52851 1 33
2 52852 1 33
2 52853 1 34
2 52854 1 34
2 52855 1 34
2 52856 1 34
2 52857 1 34
2 52858 1 34
2 52859 1 34
2 52860 1 34
2 52861 1 34
2 52862 1 34
2 52863 1 34
2 52864 1 34
2 52865 1 34
2 52866 1 34
2 52867 1 34
2 52868 1 34
2 52869 1 34
2 52870 1 35
2 52871 1 35
2 52872 1 35
2 52873 1 35
2 52874 1 35
2 52875 1 35
2 52876 1 35
2 52877 1 35
2 52878 1 35
2 52879 1 35
2 52880 1 35
2 52881 1 35
2 52882 1 35
2 52883 1 35
2 52884 1 35
2 52885 1 35
2 52886 1 35
2 52887 1 35
2 52888 1 35
2 52889 1 35
2 52890 1 35
2 52891 1 35
2 52892 1 35
2 52893 1 35
2 52894 1 35
2 52895 1 35
2 52896 1 35
2 52897 1 35
2 52898 1 35
2 52899 1 35
2 52900 1 35
2 52901 1 35
2 52902 1 35
2 52903 1 35
2 52904 1 35
2 52905 1 35
2 52906 1 35
2 52907 1 35
2 52908 1 35
2 52909 1 35
2 52910 1 35
2 52911 1 35
2 52912 1 36
2 52913 1 36
2 52914 1 36
2 52915 1 36
2 52916 1 36
2 52917 1 36
2 52918 1 36
2 52919 1 36
2 52920 1 36
2 52921 1 36
2 52922 1 36
2 52923 1 36
2 52924 1 36
2 52925 1 36
2 52926 1 36
2 52927 1 36
2 52928 1 36
2 52929 1 36
2 52930 1 36
2 52931 1 36
2 52932 1 36
2 52933 1 36
2 52934 1 36
2 52935 1 36
2 52936 1 36
2 52937 1 36
2 52938 1 36
2 52939 1 36
2 52940 1 36
2 52941 1 36
2 52942 1 36
2 52943 1 36
2 52944 1 36
2 52945 1 36
2 52946 1 36
2 52947 1 36
2 52948 1 36
2 52949 1 36
2 52950 1 36
2 52951 1 36
2 52952 1 36
2 52953 1 36
2 52954 1 36
2 52955 1 36
2 52956 1 36
2 52957 1 36
2 52958 1 36
2 52959 1 36
2 52960 1 36
2 52961 1 36
2 52962 1 36
2 52963 1 36
2 52964 1 36
2 52965 1 36
2 52966 1 36
2 52967 1 36
2 52968 1 36
2 52969 1 36
2 52970 1 36
2 52971 1 36
2 52972 1 36
2 52973 1 36
2 52974 1 36
2 52975 1 36
2 52976 1 36
2 52977 1 36
2 52978 1 36
2 52979 1 36
2 52980 1 36
2 52981 1 36
2 52982 1 36
2 52983 1 36
2 52984 1 36
2 52985 1 36
2 52986 1 36
2 52987 1 36
2 52988 1 36
2 52989 1 36
2 52990 1 36
2 52991 1 36
2 52992 1 36
2 52993 1 36
2 52994 1 36
2 52995 1 36
2 52996 1 36
2 52997 1 36
2 52998 1 36
2 52999 1 36
2 53000 1 36
2 53001 1 36
2 53002 1 36
2 53003 1 36
2 53004 1 36
2 53005 1 36
2 53006 1 36
2 53007 1 36
2 53008 1 36
2 53009 1 36
2 53010 1 36
2 53011 1 36
2 53012 1 36
2 53013 1 36
2 53014 1 36
2 53015 1 36
2 53016 1 36
2 53017 1 36
2 53018 1 36
2 53019 1 36
2 53020 1 36
2 53021 1 36
2 53022 1 36
2 53023 1 36
2 53024 1 36
2 53025 1 36
2 53026 1 36
2 53027 1 36
2 53028 1 36
2 53029 1 36
2 53030 1 36
2 53031 1 36
2 53032 1 37
2 53033 1 37
2 53034 1 37
2 53035 1 37
2 53036 1 37
2 53037 1 37
2 53038 1 37
2 53039 1 37
2 53040 1 37
2 53041 1 37
2 53042 1 37
2 53043 1 37
2 53044 1 37
2 53045 1 37
2 53046 1 37
2 53047 1 37
2 53048 1 37
2 53049 1 37
2 53050 1 37
2 53051 1 37
2 53052 1 37
2 53053 1 37
2 53054 1 37
2 53055 1 37
2 53056 1 37
2 53057 1 37
2 53058 1 37
2 53059 1 37
2 53060 1 37
2 53061 1 37
2 53062 1 37
2 53063 1 37
2 53064 1 37
2 53065 1 37
2 53066 1 37
2 53067 1 37
2 53068 1 37
2 53069 1 37
2 53070 1 37
2 53071 1 37
2 53072 1 37
2 53073 1 37
2 53074 1 37
2 53075 1 37
2 53076 1 37
2 53077 1 37
2 53078 1 37
2 53079 1 37
2 53080 1 37
2 53081 1 37
2 53082 1 37
2 53083 1 37
2 53084 1 37
2 53085 1 37
2 53086 1 37
2 53087 1 37
2 53088 1 37
2 53089 1 37
2 53090 1 37
2 53091 1 37
2 53092 1 37
2 53093 1 37
2 53094 1 37
2 53095 1 37
2 53096 1 37
2 53097 1 37
2 53098 1 37
2 53099 1 37
2 53100 1 37
2 53101 1 37
2 53102 1 37
2 53103 1 37
2 53104 1 37
2 53105 1 37
2 53106 1 37
2 53107 1 37
2 53108 1 37
2 53109 1 37
2 53110 1 37
2 53111 1 37
2 53112 1 37
2 53113 1 37
2 53114 1 37
2 53115 1 37
2 53116 1 37
2 53117 1 37
2 53118 1 37
2 53119 1 37
2 53120 1 37
2 53121 1 37
2 53122 1 37
2 53123 1 37
2 53124 1 37
2 53125 1 37
2 53126 1 37
2 53127 1 37
2 53128 1 37
2 53129 1 37
2 53130 1 37
2 53131 1 37
2 53132 1 37
2 53133 1 37
2 53134 1 37
2 53135 1 37
2 53136 1 37
2 53137 1 37
2 53138 1 37
2 53139 1 37
2 53140 1 37
2 53141 1 38
2 53142 1 38
2 53143 1 38
2 53144 1 38
2 53145 1 38
2 53146 1 38
2 53147 1 38
2 53148 1 38
2 53149 1 38
2 53150 1 38
2 53151 1 38
2 53152 1 38
2 53153 1 38
2 53154 1 38
2 53155 1 38
2 53156 1 38
2 53157 1 38
2 53158 1 38
2 53159 1 38
2 53160 1 38
2 53161 1 38
2 53162 1 38
2 53163 1 38
2 53164 1 38
2 53165 1 38
2 53166 1 38
2 53167 1 38
2 53168 1 38
2 53169 1 38
2 53170 1 38
2 53171 1 38
2 53172 1 38
2 53173 1 38
2 53174 1 38
2 53175 1 38
2 53176 1 38
2 53177 1 38
2 53178 1 38
2 53179 1 38
2 53180 1 38
2 53181 1 38
2 53182 1 38
2 53183 1 38
2 53184 1 38
2 53185 1 38
2 53186 1 38
2 53187 1 38
2 53188 1 38
2 53189 1 38
2 53190 1 38
2 53191 1 38
2 53192 1 38
2 53193 1 38
2 53194 1 38
2 53195 1 38
2 53196 1 38
2 53197 1 38
2 53198 1 38
2 53199 1 38
2 53200 1 38
2 53201 1 38
2 53202 1 38
2 53203 1 38
2 53204 1 38
2 53205 1 38
2 53206 1 38
2 53207 1 38
2 53208 1 38
2 53209 1 38
2 53210 1 38
2 53211 1 38
2 53212 1 38
2 53213 1 38
2 53214 1 38
2 53215 1 38
2 53216 1 38
2 53217 1 38
2 53218 1 38
2 53219 1 38
2 53220 1 38
2 53221 1 38
2 53222 1 38
2 53223 1 38
2 53224 1 38
2 53225 1 38
2 53226 1 38
2 53227 1 38
2 53228 1 38
2 53229 1 38
2 53230 1 38
2 53231 1 38
2 53232 1 38
2 53233 1 38
2 53234 1 38
2 53235 1 38
2 53236 1 38
2 53237 1 38
2 53238 1 38
2 53239 1 38
2 53240 1 38
2 53241 1 38
2 53242 1 38
2 53243 1 38
2 53244 1 38
2 53245 1 38
2 53246 1 38
2 53247 1 38
2 53248 1 38
2 53249 1 38
2 53250 1 38
2 53251 1 38
2 53252 1 38
2 53253 1 38
2 53254 1 38
2 53255 1 38
2 53256 1 38
2 53257 1 38
2 53258 1 39
2 53259 1 39
2 53260 1 39
2 53261 1 39
2 53262 1 39
2 53263 1 39
2 53264 1 39
2 53265 1 39
2 53266 1 39
2 53267 1 39
2 53268 1 39
2 53269 1 39
2 53270 1 39
2 53271 1 39
2 53272 1 39
2 53273 1 39
2 53274 1 39
2 53275 1 39
2 53276 1 39
2 53277 1 39
2 53278 1 39
2 53279 1 39
2 53280 1 39
2 53281 1 39
2 53282 1 39
2 53283 1 39
2 53284 1 39
2 53285 1 39
2 53286 1 39
2 53287 1 39
2 53288 1 39
2 53289 1 39
2 53290 1 39
2 53291 1 39
2 53292 1 39
2 53293 1 39
2 53294 1 39
2 53295 1 39
2 53296 1 39
2 53297 1 39
2 53298 1 39
2 53299 1 39
2 53300 1 39
2 53301 1 39
2 53302 1 39
2 53303 1 39
2 53304 1 39
2 53305 1 39
2 53306 1 39
2 53307 1 39
2 53308 1 39
2 53309 1 39
2 53310 1 39
2 53311 1 39
2 53312 1 39
2 53313 1 39
2 53314 1 39
2 53315 1 39
2 53316 1 39
2 53317 1 39
2 53318 1 39
2 53319 1 39
2 53320 1 39
2 53321 1 39
2 53322 1 39
2 53323 1 39
2 53324 1 39
2 53325 1 39
2 53326 1 39
2 53327 1 39
2 53328 1 39
2 53329 1 39
2 53330 1 39
2 53331 1 39
2 53332 1 39
2 53333 1 39
2 53334 1 39
2 53335 1 39
2 53336 1 39
2 53337 1 39
2 53338 1 39
2 53339 1 39
2 53340 1 39
2 53341 1 39
2 53342 1 39
2 53343 1 39
2 53344 1 39
2 53345 1 39
2 53346 1 39
2 53347 1 39
2 53348 1 39
2 53349 1 39
2 53350 1 39
2 53351 1 39
2 53352 1 39
2 53353 1 39
2 53354 1 39
2 53355 1 39
2 53356 1 39
2 53357 1 39
2 53358 1 39
2 53359 1 39
2 53360 1 39
2 53361 1 39
2 53362 1 39
2 53363 1 39
2 53364 1 39
2 53365 1 39
2 53366 1 39
2 53367 1 39
2 53368 1 39
2 53369 1 39
2 53370 1 39
2 53371 1 39
2 53372 1 39
2 53373 1 39
2 53374 1 39
2 53375 1 39
2 53376 1 39
2 53377 1 39
2 53378 1 39
2 53379 1 39
2 53380 1 39
2 53381 1 39
2 53382 1 39
2 53383 1 39
2 53384 1 39
2 53385 1 39
2 53386 1 39
2 53387 1 39
2 53388 1 39
2 53389 1 39
2 53390 1 39
2 53391 1 39
2 53392 1 39
2 53393 1 39
2 53394 1 39
2 53395 1 39
2 53396 1 39
2 53397 1 39
2 53398 1 39
2 53399 1 39
2 53400 1 39
2 53401 1 39
2 53402 1 39
2 53403 1 40
2 53404 1 40
2 53405 1 40
2 53406 1 40
2 53407 1 40
2 53408 1 40
2 53409 1 40
2 53410 1 40
2 53411 1 40
2 53412 1 40
2 53413 1 40
2 53414 1 40
2 53415 1 40
2 53416 1 40
2 53417 1 40
2 53418 1 40
2 53419 1 40
2 53420 1 40
2 53421 1 40
2 53422 1 40
2 53423 1 40
2 53424 1 40
2 53425 1 40
2 53426 1 40
2 53427 1 40
2 53428 1 40
2 53429 1 40
2 53430 1 40
2 53431 1 40
2 53432 1 40
2 53433 1 40
2 53434 1 40
2 53435 1 40
2 53436 1 40
2 53437 1 40
2 53438 1 40
2 53439 1 40
2 53440 1 40
2 53441 1 40
2 53442 1 40
2 53443 1 40
2 53444 1 40
2 53445 1 40
2 53446 1 40
2 53447 1 40
2 53448 1 40
2 53449 1 40
2 53450 1 40
2 53451 1 40
2 53452 1 40
2 53453 1 40
2 53454 1 40
2 53455 1 40
2 53456 1 40
2 53457 1 40
2 53458 1 40
2 53459 1 40
2 53460 1 40
2 53461 1 40
2 53462 1 40
2 53463 1 40
2 53464 1 40
2 53465 1 40
2 53466 1 40
2 53467 1 40
2 53468 1 40
2 53469 1 40
2 53470 1 40
2 53471 1 40
2 53472 1 40
2 53473 1 40
2 53474 1 40
2 53475 1 40
2 53476 1 40
2 53477 1 40
2 53478 1 40
2 53479 1 40
2 53480 1 40
2 53481 1 40
2 53482 1 40
2 53483 1 40
2 53484 1 40
2 53485 1 40
2 53486 1 40
2 53487 1 40
2 53488 1 40
2 53489 1 40
2 53490 1 40
2 53491 1 40
2 53492 1 40
2 53493 1 40
2 53494 1 40
2 53495 1 40
2 53496 1 40
2 53497 1 40
2 53498 1 40
2 53499 1 40
2 53500 1 40
2 53501 1 40
2 53502 1 40
2 53503 1 40
2 53504 1 40
2 53505 1 40
2 53506 1 40
2 53507 1 40
2 53508 1 40
2 53509 1 40
2 53510 1 40
2 53511 1 40
2 53512 1 40
2 53513 1 40
2 53514 1 40
2 53515 1 40
2 53516 1 40
2 53517 1 40
2 53518 1 40
2 53519 1 40
2 53520 1 40
2 53521 1 40
2 53522 1 40
2 53523 1 40
2 53524 1 40
2 53525 1 40
2 53526 1 40
2 53527 1 40
2 53528 1 40
2 53529 1 40
2 53530 1 40
2 53531 1 40
2 53532 1 40
2 53533 1 40
2 53534 1 40
2 53535 1 40
2 53536 1 40
2 53537 1 40
2 53538 1 40
2 53539 1 40
2 53540 1 40
2 53541 1 40
2 53542 1 40
2 53543 1 40
2 53544 1 40
2 53545 1 40
2 53546 1 40
2 53547 1 40
2 53548 1 40
2 53549 1 40
2 53550 1 40
2 53551 1 40
2 53552 1 40
2 53553 1 40
2 53554 1 40
2 53555 1 40
2 53556 1 40
2 53557 1 40
2 53558 1 40
2 53559 1 40
2 53560 1 40
2 53561 1 40
2 53562 1 40
2 53563 1 40
2 53564 1 40
2 53565 1 40
2 53566 1 40
2 53567 1 40
2 53568 1 40
2 53569 1 40
2 53570 1 40
2 53571 1 40
2 53572 1 40
2 53573 1 40
2 53574 1 40
2 53575 1 40
2 53576 1 40
2 53577 1 40
2 53578 1 40
2 53579 1 40
2 53580 1 40
2 53581 1 40
2 53582 1 40
2 53583 1 40
2 53584 1 40
2 53585 1 40
2 53586 1 40
2 53587 1 40
2 53588 1 40
2 53589 1 40
2 53590 1 40
2 53591 1 40
2 53592 1 40
2 53593 1 40
2 53594 1 40
2 53595 1 40
2 53596 1 40
2 53597 1 40
2 53598 1 40
2 53599 1 40
2 53600 1 40
2 53601 1 40
2 53602 1 40
2 53603 1 40
2 53604 1 40
2 53605 1 40
2 53606 1 40
2 53607 1 40
2 53608 1 40
2 53609 1 41
2 53610 1 41
2 53611 1 41
2 53612 1 41
2 53613 1 41
2 53614 1 41
2 53615 1 41
2 53616 1 41
2 53617 1 41
2 53618 1 41
2 53619 1 41
2 53620 1 41
2 53621 1 41
2 53622 1 41
2 53623 1 41
2 53624 1 41
2 53625 1 41
2 53626 1 41
2 53627 1 41
2 53628 1 41
2 53629 1 41
2 53630 1 41
2 53631 1 41
2 53632 1 41
2 53633 1 41
2 53634 1 41
2 53635 1 41
2 53636 1 41
2 53637 1 41
2 53638 1 41
2 53639 1 41
2 53640 1 41
2 53641 1 41
2 53642 1 41
2 53643 1 41
2 53644 1 41
2 53645 1 41
2 53646 1 41
2 53647 1 41
2 53648 1 41
2 53649 1 41
2 53650 1 41
2 53651 1 41
2 53652 1 41
2 53653 1 41
2 53654 1 41
2 53655 1 41
2 53656 1 41
2 53657 1 41
2 53658 1 41
2 53659 1 41
2 53660 1 41
2 53661 1 41
2 53662 1 41
2 53663 1 41
2 53664 1 41
2 53665 1 41
2 53666 1 41
2 53667 1 41
2 53668 1 41
2 53669 1 41
2 53670 1 41
2 53671 1 41
2 53672 1 41
2 53673 1 41
2 53674 1 41
2 53675 1 41
2 53676 1 41
2 53677 1 41
2 53678 1 41
2 53679 1 41
2 53680 1 41
2 53681 1 41
2 53682 1 41
2 53683 1 41
2 53684 1 41
2 53685 1 41
2 53686 1 41
2 53687 1 41
2 53688 1 41
2 53689 1 41
2 53690 1 41
2 53691 1 41
2 53692 1 41
2 53693 1 41
2 53694 1 41
2 53695 1 41
2 53696 1 41
2 53697 1 41
2 53698 1 41
2 53699 1 41
2 53700 1 41
2 53701 1 41
2 53702 1 41
2 53703 1 41
2 53704 1 41
2 53705 1 41
2 53706 1 41
2 53707 1 41
2 53708 1 41
2 53709 1 41
2 53710 1 41
2 53711 1 41
2 53712 1 41
2 53713 1 41
2 53714 1 41
2 53715 1 41
2 53716 1 41
2 53717 1 41
2 53718 1 41
2 53719 1 41
2 53720 1 41
2 53721 1 41
2 53722 1 41
2 53723 1 41
2 53724 1 41
2 53725 1 41
2 53726 1 41
2 53727 1 41
2 53728 1 41
2 53729 1 41
2 53730 1 41
2 53731 1 41
2 53732 1 41
2 53733 1 41
2 53734 1 41
2 53735 1 41
2 53736 1 41
2 53737 1 41
2 53738 1 41
2 53739 1 41
2 53740 1 41
2 53741 1 41
2 53742 1 41
2 53743 1 41
2 53744 1 41
2 53745 1 41
2 53746 1 41
2 53747 1 41
2 53748 1 41
2 53749 1 41
2 53750 1 41
2 53751 1 41
2 53752 1 41
2 53753 1 41
2 53754 1 41
2 53755 1 41
2 53756 1 41
2 53757 1 41
2 53758 1 41
2 53759 1 41
2 53760 1 41
2 53761 1 41
2 53762 1 41
2 53763 1 41
2 53764 1 41
2 53765 1 42
2 53766 1 42
2 53767 1 42
2 53768 1 42
2 53769 1 42
2 53770 1 42
2 53771 1 42
2 53772 1 42
2 53773 1 42
2 53774 1 42
2 53775 1 42
2 53776 1 42
2 53777 1 42
2 53778 1 42
2 53779 1 42
2 53780 1 42
2 53781 1 42
2 53782 1 42
2 53783 1 42
2 53784 1 42
2 53785 1 42
2 53786 1 42
2 53787 1 42
2 53788 1 42
2 53789 1 42
2 53790 1 42
2 53791 1 42
2 53792 1 42
2 53793 1 42
2 53794 1 42
2 53795 1 42
2 53796 1 42
2 53797 1 42
2 53798 1 42
2 53799 1 42
2 53800 1 42
2 53801 1 42
2 53802 1 42
2 53803 1 42
2 53804 1 42
2 53805 1 42
2 53806 1 42
2 53807 1 42
2 53808 1 42
2 53809 1 42
2 53810 1 42
2 53811 1 42
2 53812 1 42
2 53813 1 42
2 53814 1 42
2 53815 1 42
2 53816 1 42
2 53817 1 42
2 53818 1 42
2 53819 1 42
2 53820 1 42
2 53821 1 42
2 53822 1 42
2 53823 1 42
2 53824 1 42
2 53825 1 42
2 53826 1 42
2 53827 1 42
2 53828 1 42
2 53829 1 42
2 53830 1 42
2 53831 1 42
2 53832 1 42
2 53833 1 42
2 53834 1 42
2 53835 1 42
2 53836 1 42
2 53837 1 42
2 53838 1 42
2 53839 1 42
2 53840 1 42
2 53841 1 42
2 53842 1 42
2 53843 1 42
2 53844 1 42
2 53845 1 42
2 53846 1 42
2 53847 1 42
2 53848 1 42
2 53849 1 42
2 53850 1 42
2 53851 1 43
2 53852 1 43
2 53853 1 43
2 53854 1 43
2 53855 1 43
2 53856 1 43
2 53857 1 43
2 53858 1 43
2 53859 1 43
2 53860 1 43
2 53861 1 43
2 53862 1 43
2 53863 1 43
2 53864 1 43
2 53865 1 43
2 53866 1 43
2 53867 1 43
2 53868 1 43
2 53869 1 43
2 53870 1 43
2 53871 1 43
2 53872 1 43
2 53873 1 43
2 53874 1 43
2 53875 1 43
2 53876 1 43
2 53877 1 43
2 53878 1 43
2 53879 1 43
2 53880 1 43
2 53881 1 43
2 53882 1 43
2 53883 1 43
2 53884 1 43
2 53885 1 43
2 53886 1 43
2 53887 1 43
2 53888 1 43
2 53889 1 43
2 53890 1 43
2 53891 1 43
2 53892 1 43
2 53893 1 43
2 53894 1 43
2 53895 1 43
2 53896 1 43
2 53897 1 43
2 53898 1 43
2 53899 1 43
2 53900 1 43
2 53901 1 43
2 53902 1 43
2 53903 1 43
2 53904 1 43
2 53905 1 43
2 53906 1 43
2 53907 1 43
2 53908 1 43
2 53909 1 43
2 53910 1 43
2 53911 1 43
2 53912 1 43
2 53913 1 43
2 53914 1 43
2 53915 1 43
2 53916 1 43
2 53917 1 44
2 53918 1 44
2 53919 1 44
2 53920 1 44
2 53921 1 44
2 53922 1 44
2 53923 1 44
2 53924 1 44
2 53925 1 44
2 53926 1 44
2 53927 1 44
2 53928 1 44
2 53929 1 44
2 53930 1 44
2 53931 1 44
2 53932 1 44
2 53933 1 44
2 53934 1 44
2 53935 1 44
2 53936 1 44
2 53937 1 44
2 53938 1 44
2 53939 1 44
2 53940 1 44
2 53941 1 44
2 53942 1 44
2 53943 1 44
2 53944 1 44
2 53945 1 44
2 53946 1 44
2 53947 1 44
2 53948 1 44
2 53949 1 44
2 53950 1 44
2 53951 1 44
2 53952 1 44
2 53953 1 44
2 53954 1 44
2 53955 1 44
2 53956 1 44
2 53957 1 44
2 53958 1 44
2 53959 1 44
2 53960 1 44
2 53961 1 44
2 53962 1 44
2 53963 1 44
2 53964 1 44
2 53965 1 44
2 53966 1 44
2 53967 1 44
2 53968 1 44
2 53969 1 44
2 53970 1 44
2 53971 1 44
2 53972 1 44
2 53973 1 44
2 53974 1 44
2 53975 1 44
2 53976 1 44
2 53977 1 44
2 53978 1 44
2 53979 1 44
2 53980 1 44
2 53981 1 44
2 53982 1 44
2 53983 1 44
2 53984 1 44
2 53985 1 44
2 53986 1 44
2 53987 1 44
2 53988 1 44
2 53989 1 44
2 53990 1 44
2 53991 1 44
2 53992 1 44
2 53993 1 44
2 53994 1 44
2 53995 1 44
2 53996 1 44
2 53997 1 44
2 53998 1 44
2 53999 1 44
2 54000 1 44
2 54001 1 44
2 54002 1 44
2 54003 1 44
2 54004 1 44
2 54005 1 44
2 54006 1 44
2 54007 1 44
2 54008 1 44
2 54009 1 44
2 54010 1 44
2 54011 1 44
2 54012 1 44
2 54013 1 44
2 54014 1 44
2 54015 1 44
2 54016 1 44
2 54017 1 44
2 54018 1 44
2 54019 1 44
2 54020 1 44
2 54021 1 44
2 54022 1 44
2 54023 1 44
2 54024 1 44
2 54025 1 44
2 54026 1 44
2 54027 1 44
2 54028 1 44
2 54029 1 44
2 54030 1 44
2 54031 1 44
2 54032 1 44
2 54033 1 44
2 54034 1 44
2 54035 1 44
2 54036 1 44
2 54037 1 44
2 54038 1 44
2 54039 1 44
2 54040 1 44
2 54041 1 44
2 54042 1 44
2 54043 1 44
2 54044 1 44
2 54045 1 44
2 54046 1 44
2 54047 1 44
2 54048 1 44
2 54049 1 44
2 54050 1 44
2 54051 1 44
2 54052 1 44
2 54053 1 44
2 54054 1 44
2 54055 1 44
2 54056 1 44
2 54057 1 44
2 54058 1 44
2 54059 1 44
2 54060 1 44
2 54061 1 44
2 54062 1 44
2 54063 1 44
2 54064 1 44
2 54065 1 44
2 54066 1 44
2 54067 1 44
2 54068 1 44
2 54069 1 44
2 54070 1 44
2 54071 1 44
2 54072 1 44
2 54073 1 44
2 54074 1 44
2 54075 1 44
2 54076 1 44
2 54077 1 44
2 54078 1 44
2 54079 1 44
2 54080 1 44
2 54081 1 44
2 54082 1 44
2 54083 1 44
2 54084 1 44
2 54085 1 44
2 54086 1 44
2 54087 1 44
2 54088 1 44
2 54089 1 44
2 54090 1 44
2 54091 1 44
2 54092 1 44
2 54093 1 44
2 54094 1 44
2 54095 1 44
2 54096 1 44
2 54097 1 44
2 54098 1 44
2 54099 1 44
2 54100 1 44
2 54101 1 44
2 54102 1 44
2 54103 1 44
2 54104 1 44
2 54105 1 44
2 54106 1 44
2 54107 1 44
2 54108 1 44
2 54109 1 44
2 54110 1 44
2 54111 1 44
2 54112 1 44
2 54113 1 44
2 54114 1 44
2 54115 1 44
2 54116 1 44
2 54117 1 45
2 54118 1 45
2 54119 1 45
2 54120 1 45
2 54121 1 45
2 54122 1 45
2 54123 1 45
2 54124 1 45
2 54125 1 45
2 54126 1 45
2 54127 1 45
2 54128 1 45
2 54129 1 45
2 54130 1 45
2 54131 1 45
2 54132 1 45
2 54133 1 45
2 54134 1 45
2 54135 1 45
2 54136 1 45
2 54137 1 45
2 54138 1 45
2 54139 1 45
2 54140 1 45
2 54141 1 45
2 54142 1 45
2 54143 1 45
2 54144 1 45
2 54145 1 45
2 54146 1 45
2 54147 1 45
2 54148 1 45
2 54149 1 45
2 54150 1 45
2 54151 1 45
2 54152 1 45
2 54153 1 45
2 54154 1 45
2 54155 1 45
2 54156 1 45
2 54157 1 45
2 54158 1 45
2 54159 1 45
2 54160 1 45
2 54161 1 45
2 54162 1 45
2 54163 1 45
2 54164 1 45
2 54165 1 45
2 54166 1 45
2 54167 1 45
2 54168 1 45
2 54169 1 45
2 54170 1 45
2 54171 1 45
2 54172 1 45
2 54173 1 45
2 54174 1 45
2 54175 1 45
2 54176 1 45
2 54177 1 45
2 54178 1 45
2 54179 1 45
2 54180 1 45
2 54181 1 45
2 54182 1 45
2 54183 1 45
2 54184 1 45
2 54185 1 45
2 54186 1 45
2 54187 1 45
2 54188 1 45
2 54189 1 45
2 54190 1 45
2 54191 1 45
2 54192 1 45
2 54193 1 45
2 54194 1 45
2 54195 1 45
2 54196 1 45
2 54197 1 45
2 54198 1 45
2 54199 1 45
2 54200 1 45
2 54201 1 45
2 54202 1 45
2 54203 1 45
2 54204 1 45
2 54205 1 45
2 54206 1 45
2 54207 1 45
2 54208 1 45
2 54209 1 45
2 54210 1 45
2 54211 1 45
2 54212 1 45
2 54213 1 45
2 54214 1 45
2 54215 1 45
2 54216 1 45
2 54217 1 45
2 54218 1 45
2 54219 1 45
2 54220 1 45
2 54221 1 45
2 54222 1 45
2 54223 1 45
2 54224 1 45
2 54225 1 45
2 54226 1 45
2 54227 1 45
2 54228 1 45
2 54229 1 45
2 54230 1 45
2 54231 1 45
2 54232 1 45
2 54233 1 45
2 54234 1 45
2 54235 1 45
2 54236 1 45
2 54237 1 45
2 54238 1 45
2 54239 1 45
2 54240 1 45
2 54241 1 45
2 54242 1 45
2 54243 1 45
2 54244 1 45
2 54245 1 45
2 54246 1 45
2 54247 1 45
2 54248 1 45
2 54249 1 45
2 54250 1 45
2 54251 1 45
2 54252 1 45
2 54253 1 45
2 54254 1 45
2 54255 1 45
2 54256 1 45
2 54257 1 45
2 54258 1 45
2 54259 1 45
2 54260 1 45
2 54261 1 45
2 54262 1 45
2 54263 1 45
2 54264 1 45
2 54265 1 45
2 54266 1 45
2 54267 1 45
2 54268 1 45
2 54269 1 45
2 54270 1 45
2 54271 1 45
2 54272 1 45
2 54273 1 45
2 54274 1 45
2 54275 1 45
2 54276 1 45
2 54277 1 45
2 54278 1 45
2 54279 1 45
2 54280 1 45
2 54281 1 45
2 54282 1 45
2 54283 1 45
2 54284 1 45
2 54285 1 45
2 54286 1 45
2 54287 1 45
2 54288 1 45
2 54289 1 45
2 54290 1 45
2 54291 1 45
2 54292 1 45
2 54293 1 45
2 54294 1 45
2 54295 1 45
2 54296 1 45
2 54297 1 45
2 54298 1 45
2 54299 1 45
2 54300 1 45
2 54301 1 45
2 54302 1 45
2 54303 1 45
2 54304 1 45
2 54305 1 45
2 54306 1 45
2 54307 1 45
2 54308 1 45
2 54309 1 45
2 54310 1 45
2 54311 1 45
2 54312 1 45
2 54313 1 45
2 54314 1 45
2 54315 1 45
2 54316 1 45
2 54317 1 45
2 54318 1 45
2 54319 1 45
2 54320 1 45
2 54321 1 45
2 54322 1 45
2 54323 1 45
2 54324 1 45
2 54325 1 45
2 54326 1 45
2 54327 1 45
2 54328 1 45
2 54329 1 45
2 54330 1 45
2 54331 1 45
2 54332 1 45
2 54333 1 45
2 54334 1 45
2 54335 1 45
2 54336 1 45
2 54337 1 45
2 54338 1 45
2 54339 1 45
2 54340 1 45
2 54341 1 45
2 54342 1 45
2 54343 1 45
2 54344 1 45
2 54345 1 45
2 54346 1 45
2 54347 1 45
2 54348 1 45
2 54349 1 45
2 54350 1 45
2 54351 1 45
2 54352 1 45
2 54353 1 45
2 54354 1 45
2 54355 1 45
2 54356 1 45
2 54357 1 45
2 54358 1 45
2 54359 1 45
2 54360 1 45
2 54361 1 45
2 54362 1 45
2 54363 1 45
2 54364 1 45
2 54365 1 45
2 54366 1 45
2 54367 1 45
2 54368 1 45
2 54369 1 45
2 54370 1 45
2 54371 1 45
2 54372 1 45
2 54373 1 45
2 54374 1 45
2 54375 1 45
2 54376 1 45
2 54377 1 45
2 54378 1 45
2 54379 1 45
2 54380 1 45
2 54381 1 45
2 54382 1 45
2 54383 1 45
2 54384 1 45
2 54385 1 45
2 54386 1 45
2 54387 1 45
2 54388 1 45
2 54389 1 45
2 54390 1 45
2 54391 1 45
2 54392 1 45
2 54393 1 45
2 54394 1 45
2 54395 1 45
2 54396 1 45
2 54397 1 45
2 54398 1 45
2 54399 1 45
2 54400 1 45
2 54401 1 45
2 54402 1 45
2 54403 1 45
2 54404 1 45
2 54405 1 45
2 54406 1 45
2 54407 1 45
2 54408 1 45
2 54409 1 45
2 54410 1 45
2 54411 1 45
2 54412 1 45
2 54413 1 45
2 54414 1 45
2 54415 1 45
2 54416 1 45
2 54417 1 45
2 54418 1 46
2 54419 1 46
2 54420 1 46
2 54421 1 46
2 54422 1 46
2 54423 1 46
2 54424 1 46
2 54425 1 46
2 54426 1 46
2 54427 1 46
2 54428 1 46
2 54429 1 46
2 54430 1 46
2 54431 1 46
2 54432 1 46
2 54433 1 46
2 54434 1 46
2 54435 1 46
2 54436 1 46
2 54437 1 46
2 54438 1 46
2 54439 1 46
2 54440 1 46
2 54441 1 46
2 54442 1 46
2 54443 1 46
2 54444 1 46
2 54445 1 46
2 54446 1 46
2 54447 1 46
2 54448 1 46
2 54449 1 46
2 54450 1 46
2 54451 1 46
2 54452 1 46
2 54453 1 46
2 54454 1 46
2 54455 1 46
2 54456 1 46
2 54457 1 46
2 54458 1 46
2 54459 1 46
2 54460 1 46
2 54461 1 46
2 54462 1 46
2 54463 1 46
2 54464 1 46
2 54465 1 46
2 54466 1 46
2 54467 1 46
2 54468 1 46
2 54469 1 46
2 54470 1 46
2 54471 1 46
2 54472 1 46
2 54473 1 46
2 54474 1 46
2 54475 1 46
2 54476 1 46
2 54477 1 46
2 54478 1 46
2 54479 1 46
2 54480 1 46
2 54481 1 46
2 54482 1 46
2 54483 1 46
2 54484 1 46
2 54485 1 46
2 54486 1 46
2 54487 1 46
2 54488 1 46
2 54489 1 46
2 54490 1 46
2 54491 1 46
2 54492 1 46
2 54493 1 46
2 54494 1 46
2 54495 1 46
2 54496 1 46
2 54497 1 46
2 54498 1 46
2 54499 1 46
2 54500 1 46
2 54501 1 46
2 54502 1 46
2 54503 1 46
2 54504 1 46
2 54505 1 46
2 54506 1 46
2 54507 1 46
2 54508 1 46
2 54509 1 46
2 54510 1 46
2 54511 1 46
2 54512 1 46
2 54513 1 46
2 54514 1 46
2 54515 1 46
2 54516 1 46
2 54517 1 46
2 54518 1 46
2 54519 1 46
2 54520 1 46
2 54521 1 46
2 54522 1 46
2 54523 1 46
2 54524 1 46
2 54525 1 46
2 54526 1 46
2 54527 1 46
2 54528 1 46
2 54529 1 46
2 54530 1 46
2 54531 1 46
2 54532 1 46
2 54533 1 46
2 54534 1 46
2 54535 1 46
2 54536 1 46
2 54537 1 46
2 54538 1 46
2 54539 1 46
2 54540 1 46
2 54541 1 46
2 54542 1 46
2 54543 1 46
2 54544 1 46
2 54545 1 46
2 54546 1 46
2 54547 1 46
2 54548 1 46
2 54549 1 46
2 54550 1 46
2 54551 1 46
2 54552 1 46
2 54553 1 46
2 54554 1 46
2 54555 1 46
2 54556 1 46
2 54557 1 46
2 54558 1 46
2 54559 1 46
2 54560 1 46
2 54561 1 46
2 54562 1 46
2 54563 1 46
2 54564 1 46
2 54565 1 46
2 54566 1 46
2 54567 1 46
2 54568 1 46
2 54569 1 46
2 54570 1 46
2 54571 1 46
2 54572 1 46
2 54573 1 46
2 54574 1 46
2 54575 1 46
2 54576 1 46
2 54577 1 46
2 54578 1 46
2 54579 1 46
2 54580 1 46
2 54581 1 46
2 54582 1 46
2 54583 1 46
2 54584 1 46
2 54585 1 46
2 54586 1 46
2 54587 1 46
2 54588 1 46
2 54589 1 46
2 54590 1 46
2 54591 1 46
2 54592 1 46
2 54593 1 46
2 54594 1 46
2 54595 1 46
2 54596 1 46
2 54597 1 46
2 54598 1 46
2 54599 1 46
2 54600 1 46
2 54601 1 46
2 54602 1 46
2 54603 1 46
2 54604 1 46
2 54605 1 46
2 54606 1 46
2 54607 1 46
2 54608 1 46
2 54609 1 46
2 54610 1 46
2 54611 1 46
2 54612 1 46
2 54613 1 46
2 54614 1 46
2 54615 1 46
2 54616 1 46
2 54617 1 46
2 54618 1 46
2 54619 1 46
2 54620 1 46
2 54621 1 46
2 54622 1 46
2 54623 1 46
2 54624 1 46
2 54625 1 46
2 54626 1 46
2 54627 1 46
2 54628 1 46
2 54629 1 46
2 54630 1 46
2 54631 1 46
2 54632 1 46
2 54633 1 46
2 54634 1 46
2 54635 1 46
2 54636 1 46
2 54637 1 46
2 54638 1 46
2 54639 1 46
2 54640 1 46
2 54641 1 46
2 54642 1 46
2 54643 1 46
2 54644 1 46
2 54645 1 46
2 54646 1 46
2 54647 1 46
2 54648 1 46
2 54649 1 46
2 54650 1 46
2 54651 1 46
2 54652 1 46
2 54653 1 46
2 54654 1 46
2 54655 1 46
2 54656 1 46
2 54657 1 46
2 54658 1 46
2 54659 1 46
2 54660 1 46
2 54661 1 46
2 54662 1 46
2 54663 1 46
2 54664 1 46
2 54665 1 46
2 54666 1 46
2 54667 1 46
2 54668 1 46
2 54669 1 46
2 54670 1 46
2 54671 1 46
2 54672 1 46
2 54673 1 46
2 54674 1 46
2 54675 1 46
2 54676 1 46
2 54677 1 46
2 54678 1 46
2 54679 1 46
2 54680 1 46
2 54681 1 46
2 54682 1 46
2 54683 1 46
2 54684 1 46
2 54685 1 46
2 54686 1 46
2 54687 1 46
2 54688 1 46
2 54689 1 46
2 54690 1 46
2 54691 1 46
2 54692 1 46
2 54693 1 46
2 54694 1 46
2 54695 1 46
2 54696 1 46
2 54697 1 46
2 54698 1 46
2 54699 1 46
2 54700 1 46
2 54701 1 46
2 54702 1 46
2 54703 1 46
2 54704 1 46
2 54705 1 46
2 54706 1 46
2 54707 1 46
2 54708 1 46
2 54709 1 46
2 54710 1 46
2 54711 1 46
2 54712 1 46
2 54713 1 46
2 54714 1 46
2 54715 1 46
2 54716 1 46
2 54717 1 46
2 54718 1 46
2 54719 1 46
2 54720 1 46
2 54721 1 46
2 54722 1 46
2 54723 1 46
2 54724 1 46
2 54725 1 46
2 54726 1 46
2 54727 1 46
2 54728 1 46
2 54729 1 46
2 54730 1 46
2 54731 1 46
2 54732 1 46
2 54733 1 46
2 54734 1 46
2 54735 1 46
2 54736 1 46
2 54737 1 46
2 54738 1 46
2 54739 1 46
2 54740 1 46
2 54741 1 46
2 54742 1 46
2 54743 1 46
2 54744 1 46
2 54745 1 46
2 54746 1 46
2 54747 1 46
2 54748 1 46
2 54749 1 46
2 54750 1 46
2 54751 1 46
2 54752 1 46
2 54753 1 46
2 54754 1 46
2 54755 1 46
2 54756 1 46
2 54757 1 46
2 54758 1 46
2 54759 1 46
2 54760 1 46
2 54761 1 46
2 54762 1 46
2 54763 1 46
2 54764 1 46
2 54765 1 46
2 54766 1 46
2 54767 1 46
2 54768 1 46
2 54769 1 46
2 54770 1 46
2 54771 1 46
2 54772 1 46
2 54773 1 46
2 54774 1 46
2 54775 1 46
2 54776 1 46
2 54777 1 46
2 54778 1 46
2 54779 1 46
2 54780 1 46
2 54781 1 46
2 54782 1 46
2 54783 1 46
2 54784 1 46
2 54785 1 46
2 54786 1 46
2 54787 1 46
2 54788 1 46
2 54789 1 46
2 54790 1 46
2 54791 1 46
2 54792 1 46
2 54793 1 46
2 54794 1 46
2 54795 1 46
2 54796 1 46
2 54797 1 46
2 54798 1 46
2 54799 1 46
2 54800 1 46
2 54801 1 46
2 54802 1 46
2 54803 1 46
2 54804 1 46
2 54805 1 46
2 54806 1 46
2 54807 1 46
2 54808 1 46
2 54809 1 46
2 54810 1 46
2 54811 1 47
2 54812 1 47
2 54813 1 47
2 54814 1 47
2 54815 1 47
2 54816 1 47
2 54817 1 47
2 54818 1 47
2 54819 1 47
2 54820 1 47
2 54821 1 47
2 54822 1 47
2 54823 1 47
2 54824 1 47
2 54825 1 47
2 54826 1 47
2 54827 1 47
2 54828 1 47
2 54829 1 47
2 54830 1 47
2 54831 1 47
2 54832 1 47
2 54833 1 47
2 54834 1 47
2 54835 1 47
2 54836 1 47
2 54837 1 47
2 54838 1 47
2 54839 1 47
2 54840 1 47
2 54841 1 47
2 54842 1 47
2 54843 1 47
2 54844 1 47
2 54845 1 47
2 54846 1 47
2 54847 1 47
2 54848 1 47
2 54849 1 47
2 54850 1 47
2 54851 1 47
2 54852 1 47
2 54853 1 47
2 54854 1 47
2 54855 1 47
2 54856 1 47
2 54857 1 47
2 54858 1 47
2 54859 1 47
2 54860 1 47
2 54861 1 47
2 54862 1 47
2 54863 1 47
2 54864 1 47
2 54865 1 47
2 54866 1 47
2 54867 1 47
2 54868 1 47
2 54869 1 47
2 54870 1 47
2 54871 1 47
2 54872 1 47
2 54873 1 47
2 54874 1 47
2 54875 1 47
2 54876 1 47
2 54877 1 47
2 54878 1 47
2 54879 1 47
2 54880 1 47
2 54881 1 47
2 54882 1 47
2 54883 1 47
2 54884 1 47
2 54885 1 47
2 54886 1 47
2 54887 1 47
2 54888 1 47
2 54889 1 47
2 54890 1 47
2 54891 1 47
2 54892 1 47
2 54893 1 47
2 54894 1 47
2 54895 1 47
2 54896 1 47
2 54897 1 47
2 54898 1 47
2 54899 1 47
2 54900 1 47
2 54901 1 47
2 54902 1 47
2 54903 1 47
2 54904 1 47
2 54905 1 47
2 54906 1 47
2 54907 1 47
2 54908 1 47
2 54909 1 47
2 54910 1 47
2 54911 1 47
2 54912 1 47
2 54913 1 47
2 54914 1 47
2 54915 1 47
2 54916 1 47
2 54917 1 47
2 54918 1 47
2 54919 1 47
2 54920 1 47
2 54921 1 47
2 54922 1 47
2 54923 1 47
2 54924 1 47
2 54925 1 47
2 54926 1 47
2 54927 1 47
2 54928 1 47
2 54929 1 47
2 54930 1 47
2 54931 1 47
2 54932 1 47
2 54933 1 47
2 54934 1 47
2 54935 1 47
2 54936 1 47
2 54937 1 47
2 54938 1 47
2 54939 1 47
2 54940 1 47
2 54941 1 47
2 54942 1 47
2 54943 1 47
2 54944 1 47
2 54945 1 47
2 54946 1 47
2 54947 1 47
2 54948 1 47
2 54949 1 47
2 54950 1 47
2 54951 1 47
2 54952 1 47
2 54953 1 47
2 54954 1 47
2 54955 1 47
2 54956 1 47
2 54957 1 47
2 54958 1 47
2 54959 1 47
2 54960 1 47
2 54961 1 47
2 54962 1 47
2 54963 1 47
2 54964 1 47
2 54965 1 47
2 54966 1 47
2 54967 1 47
2 54968 1 47
2 54969 1 47
2 54970 1 47
2 54971 1 47
2 54972 1 47
2 54973 1 47
2 54974 1 47
2 54975 1 47
2 54976 1 47
2 54977 1 47
2 54978 1 47
2 54979 1 47
2 54980 1 47
2 54981 1 47
2 54982 1 47
2 54983 1 47
2 54984 1 47
2 54985 1 47
2 54986 1 47
2 54987 1 47
2 54988 1 47
2 54989 1 47
2 54990 1 47
2 54991 1 47
2 54992 1 47
2 54993 1 47
2 54994 1 47
2 54995 1 47
2 54996 1 47
2 54997 1 47
2 54998 1 47
2 54999 1 47
2 55000 1 47
2 55001 1 47
2 55002 1 47
2 55003 1 47
2 55004 1 47
2 55005 1 47
2 55006 1 47
2 55007 1 47
2 55008 1 47
2 55009 1 47
2 55010 1 47
2 55011 1 47
2 55012 1 47
2 55013 1 47
2 55014 1 47
2 55015 1 47
2 55016 1 47
2 55017 1 47
2 55018 1 47
2 55019 1 47
2 55020 1 47
2 55021 1 47
2 55022 1 47
2 55023 1 47
2 55024 1 47
2 55025 1 47
2 55026 1 47
2 55027 1 47
2 55028 1 47
2 55029 1 47
2 55030 1 47
2 55031 1 47
2 55032 1 47
2 55033 1 47
2 55034 1 47
2 55035 1 47
2 55036 1 47
2 55037 1 47
2 55038 1 47
2 55039 1 47
2 55040 1 47
2 55041 1 47
2 55042 1 47
2 55043 1 47
2 55044 1 47
2 55045 1 47
2 55046 1 47
2 55047 1 47
2 55048 1 47
2 55049 1 47
2 55050 1 47
2 55051 1 47
2 55052 1 47
2 55053 1 47
2 55054 1 47
2 55055 1 47
2 55056 1 47
2 55057 1 47
2 55058 1 47
2 55059 1 47
2 55060 1 47
2 55061 1 47
2 55062 1 47
2 55063 1 47
2 55064 1 47
2 55065 1 47
2 55066 1 47
2 55067 1 47
2 55068 1 47
2 55069 1 47
2 55070 1 47
2 55071 1 47
2 55072 1 47
2 55073 1 47
2 55074 1 47
2 55075 1 47
2 55076 1 47
2 55077 1 47
2 55078 1 47
2 55079 1 47
2 55080 1 47
2 55081 1 47
2 55082 1 47
2 55083 1 47
2 55084 1 47
2 55085 1 47
2 55086 1 47
2 55087 1 47
2 55088 1 47
2 55089 1 47
2 55090 1 47
2 55091 1 47
2 55092 1 47
2 55093 1 47
2 55094 1 47
2 55095 1 47
2 55096 1 47
2 55097 1 47
2 55098 1 47
2 55099 1 47
2 55100 1 47
2 55101 1 47
2 55102 1 47
2 55103 1 47
2 55104 1 47
2 55105 1 47
2 55106 1 47
2 55107 1 47
2 55108 1 47
2 55109 1 47
2 55110 1 47
2 55111 1 47
2 55112 1 47
2 55113 1 47
2 55114 1 47
2 55115 1 47
2 55116 1 47
2 55117 1 47
2 55118 1 47
2 55119 1 47
2 55120 1 47
2 55121 1 47
2 55122 1 47
2 55123 1 47
2 55124 1 47
2 55125 1 47
2 55126 1 47
2 55127 1 47
2 55128 1 47
2 55129 1 47
2 55130 1 47
2 55131 1 47
2 55132 1 47
2 55133 1 47
2 55134 1 47
2 55135 1 47
2 55136 1 47
2 55137 1 47
2 55138 1 47
2 55139 1 47
2 55140 1 47
2 55141 1 47
2 55142 1 47
2 55143 1 47
2 55144 1 47
2 55145 1 47
2 55146 1 47
2 55147 1 47
2 55148 1 47
2 55149 1 47
2 55150 1 47
2 55151 1 47
2 55152 1 47
2 55153 1 47
2 55154 1 47
2 55155 1 47
2 55156 1 47
2 55157 1 47
2 55158 1 47
2 55159 1 47
2 55160 1 48
2 55161 1 48
2 55162 1 48
2 55163 1 48
2 55164 1 48
2 55165 1 48
2 55166 1 48
2 55167 1 48
2 55168 1 48
2 55169 1 48
2 55170 1 48
2 55171 1 48
2 55172 1 48
2 55173 1 48
2 55174 1 48
2 55175 1 48
2 55176 1 48
2 55177 1 48
2 55178 1 48
2 55179 1 48
2 55180 1 48
2 55181 1 48
2 55182 1 48
2 55183 1 48
2 55184 1 48
2 55185 1 48
2 55186 1 48
2 55187 1 48
2 55188 1 48
2 55189 1 48
2 55190 1 48
2 55191 1 48
2 55192 1 48
2 55193 1 48
2 55194 1 48
2 55195 1 48
2 55196 1 48
2 55197 1 48
2 55198 1 48
2 55199 1 48
2 55200 1 48
2 55201 1 48
2 55202 1 48
2 55203 1 48
2 55204 1 48
2 55205 1 48
2 55206 1 48
2 55207 1 48
2 55208 1 48
2 55209 1 48
2 55210 1 48
2 55211 1 48
2 55212 1 48
2 55213 1 48
2 55214 1 48
2 55215 1 48
2 55216 1 48
2 55217 1 48
2 55218 1 48
2 55219 1 48
2 55220 1 48
2 55221 1 48
2 55222 1 48
2 55223 1 48
2 55224 1 48
2 55225 1 48
2 55226 1 48
2 55227 1 48
2 55228 1 48
2 55229 1 48
2 55230 1 48
2 55231 1 48
2 55232 1 48
2 55233 1 48
2 55234 1 48
2 55235 1 48
2 55236 1 48
2 55237 1 48
2 55238 1 48
2 55239 1 48
2 55240 1 48
2 55241 1 48
2 55242 1 48
2 55243 1 48
2 55244 1 48
2 55245 1 48
2 55246 1 48
2 55247 1 48
2 55248 1 48
2 55249 1 48
2 55250 1 48
2 55251 1 48
2 55252 1 48
2 55253 1 48
2 55254 1 48
2 55255 1 48
2 55256 1 48
2 55257 1 48
2 55258 1 48
2 55259 1 48
2 55260 1 48
2 55261 1 48
2 55262 1 48
2 55263 1 48
2 55264 1 48
2 55265 1 48
2 55266 1 48
2 55267 1 48
2 55268 1 48
2 55269 1 48
2 55270 1 48
2 55271 1 48
2 55272 1 48
2 55273 1 48
2 55274 1 48
2 55275 1 48
2 55276 1 48
2 55277 1 48
2 55278 1 48
2 55279 1 48
2 55280 1 48
2 55281 1 48
2 55282 1 48
2 55283 1 48
2 55284 1 48
2 55285 1 48
2 55286 1 48
2 55287 1 48
2 55288 1 48
2 55289 1 48
2 55290 1 48
2 55291 1 48
2 55292 1 48
2 55293 1 48
2 55294 1 48
2 55295 1 48
2 55296 1 48
2 55297 1 48
2 55298 1 48
2 55299 1 48
2 55300 1 48
2 55301 1 48
2 55302 1 48
2 55303 1 48
2 55304 1 48
2 55305 1 48
2 55306 1 48
2 55307 1 48
2 55308 1 48
2 55309 1 48
2 55310 1 48
2 55311 1 48
2 55312 1 48
2 55313 1 48
2 55314 1 48
2 55315 1 48
2 55316 1 48
2 55317 1 48
2 55318 1 48
2 55319 1 48
2 55320 1 48
2 55321 1 48
2 55322 1 48
2 55323 1 48
2 55324 1 48
2 55325 1 48
2 55326 1 48
2 55327 1 48
2 55328 1 48
2 55329 1 48
2 55330 1 48
2 55331 1 48
2 55332 1 48
2 55333 1 48
2 55334 1 48
2 55335 1 48
2 55336 1 48
2 55337 1 48
2 55338 1 48
2 55339 1 48
2 55340 1 48
2 55341 1 48
2 55342 1 48
2 55343 1 48
2 55344 1 48
2 55345 1 48
2 55346 1 48
2 55347 1 48
2 55348 1 48
2 55349 1 48
2 55350 1 48
2 55351 1 48
2 55352 1 48
2 55353 1 48
2 55354 1 48
2 55355 1 48
2 55356 1 48
2 55357 1 48
2 55358 1 48
2 55359 1 48
2 55360 1 48
2 55361 1 48
2 55362 1 48
2 55363 1 48
2 55364 1 48
2 55365 1 48
2 55366 1 48
2 55367 1 48
2 55368 1 48
2 55369 1 48
2 55370 1 48
2 55371 1 48
2 55372 1 48
2 55373 1 48
2 55374 1 48
2 55375 1 48
2 55376 1 48
2 55377 1 48
2 55378 1 48
2 55379 1 48
2 55380 1 48
2 55381 1 48
2 55382 1 48
2 55383 1 48
2 55384 1 48
2 55385 1 48
2 55386 1 48
2 55387 1 48
2 55388 1 48
2 55389 1 48
2 55390 1 48
2 55391 1 48
2 55392 1 48
2 55393 1 48
2 55394 1 48
2 55395 1 48
2 55396 1 48
2 55397 1 48
2 55398 1 48
2 55399 1 48
2 55400 1 48
2 55401 1 48
2 55402 1 48
2 55403 1 48
2 55404 1 48
2 55405 1 48
2 55406 1 48
2 55407 1 48
2 55408 1 48
2 55409 1 48
2 55410 1 48
2 55411 1 48
2 55412 1 48
2 55413 1 48
2 55414 1 48
2 55415 1 48
2 55416 1 48
2 55417 1 48
2 55418 1 48
2 55419 1 48
2 55420 1 48
2 55421 1 48
2 55422 1 48
2 55423 1 48
2 55424 1 48
2 55425 1 48
2 55426 1 48
2 55427 1 48
2 55428 1 48
2 55429 1 48
2 55430 1 48
2 55431 1 48
2 55432 1 49
2 55433 1 49
2 55434 1 49
2 55435 1 49
2 55436 1 49
2 55437 1 49
2 55438 1 49
2 55439 1 49
2 55440 1 49
2 55441 1 49
2 55442 1 49
2 55443 1 49
2 55444 1 49
2 55445 1 49
2 55446 1 49
2 55447 1 49
2 55448 1 49
2 55449 1 49
2 55450 1 49
2 55451 1 49
2 55452 1 49
2 55453 1 49
2 55454 1 49
2 55455 1 49
2 55456 1 49
2 55457 1 49
2 55458 1 49
2 55459 1 49
2 55460 1 49
2 55461 1 49
2 55462 1 49
2 55463 1 49
2 55464 1 49
2 55465 1 49
2 55466 1 49
2 55467 1 49
2 55468 1 49
2 55469 1 49
2 55470 1 49
2 55471 1 49
2 55472 1 49
2 55473 1 49
2 55474 1 49
2 55475 1 49
2 55476 1 49
2 55477 1 49
2 55478 1 49
2 55479 1 49
2 55480 1 49
2 55481 1 49
2 55482 1 49
2 55483 1 49
2 55484 1 49
2 55485 1 49
2 55486 1 49
2 55487 1 49
2 55488 1 49
2 55489 1 49
2 55490 1 49
2 55491 1 49
2 55492 1 49
2 55493 1 49
2 55494 1 49
2 55495 1 49
2 55496 1 49
2 55497 1 49
2 55498 1 49
2 55499 1 49
2 55500 1 49
2 55501 1 49
2 55502 1 49
2 55503 1 49
2 55504 1 49
2 55505 1 49
2 55506 1 49
2 55507 1 49
2 55508 1 49
2 55509 1 49
2 55510 1 49
2 55511 1 49
2 55512 1 49
2 55513 1 49
2 55514 1 49
2 55515 1 49
2 55516 1 49
2 55517 1 49
2 55518 1 49
2 55519 1 49
2 55520 1 49
2 55521 1 49
2 55522 1 49
2 55523 1 49
2 55524 1 49
2 55525 1 49
2 55526 1 49
2 55527 1 49
2 55528 1 49
2 55529 1 49
2 55530 1 49
2 55531 1 49
2 55532 1 49
2 55533 1 49
2 55534 1 49
2 55535 1 49
2 55536 1 49
2 55537 1 49
2 55538 1 49
2 55539 1 49
2 55540 1 49
2 55541 1 49
2 55542 1 49
2 55543 1 49
2 55544 1 49
2 55545 1 49
2 55546 1 49
2 55547 1 49
2 55548 1 49
2 55549 1 49
2 55550 1 49
2 55551 1 49
2 55552 1 49
2 55553 1 49
2 55554 1 49
2 55555 1 49
2 55556 1 49
2 55557 1 49
2 55558 1 49
2 55559 1 49
2 55560 1 49
2 55561 1 49
2 55562 1 49
2 55563 1 49
2 55564 1 49
2 55565 1 49
2 55566 1 49
2 55567 1 49
2 55568 1 49
2 55569 1 49
2 55570 1 49
2 55571 1 49
2 55572 1 49
2 55573 1 49
2 55574 1 49
2 55575 1 49
2 55576 1 49
2 55577 1 49
2 55578 1 49
2 55579 1 49
2 55580 1 49
2 55581 1 49
2 55582 1 49
2 55583 1 49
2 55584 1 49
2 55585 1 49
2 55586 1 49
2 55587 1 49
2 55588 1 49
2 55589 1 49
2 55590 1 49
2 55591 1 49
2 55592 1 49
2 55593 1 50
2 55594 1 50
2 55595 1 50
2 55596 1 50
2 55597 1 50
2 55598 1 50
2 55599 1 50
2 55600 1 50
2 55601 1 50
2 55602 1 50
2 55603 1 50
2 55604 1 50
2 55605 1 50
2 55606 1 50
2 55607 1 50
2 55608 1 50
2 55609 1 50
2 55610 1 50
2 55611 1 50
2 55612 1 50
2 55613 1 50
2 55614 1 50
2 55615 1 50
2 55616 1 50
2 55617 1 50
2 55618 1 50
2 55619 1 50
2 55620 1 50
2 55621 1 50
2 55622 1 50
2 55623 1 50
2 55624 1 50
2 55625 1 50
2 55626 1 50
2 55627 1 50
2 55628 1 50
2 55629 1 50
2 55630 1 50
2 55631 1 50
2 55632 1 50
2 55633 1 50
2 55634 1 50
2 55635 1 50
2 55636 1 50
2 55637 1 50
2 55638 1 50
2 55639 1 50
2 55640 1 50
2 55641 1 50
2 55642 1 50
2 55643 1 50
2 55644 1 50
2 55645 1 50
2 55646 1 50
2 55647 1 50
2 55648 1 50
2 55649 1 50
2 55650 1 50
2 55651 1 50
2 55652 1 50
2 55653 1 50
2 55654 1 50
2 55655 1 50
2 55656 1 50
2 55657 1 50
2 55658 1 50
2 55659 1 50
2 55660 1 52
2 55661 1 52
2 55662 1 52
2 55663 1 52
2 55664 1 52
2 55665 1 52
2 55666 1 52
2 55667 1 52
2 55668 1 52
2 55669 1 52
2 55670 1 52
2 55671 1 52
2 55672 1 52
2 55673 1 52
2 55674 1 52
2 55675 1 52
2 55676 1 52
2 55677 1 52
2 55678 1 52
2 55679 1 52
2 55680 1 52
2 55681 1 52
2 55682 1 52
2 55683 1 52
2 55684 1 52
2 55685 1 52
2 55686 1 52
2 55687 1 52
2 55688 1 52
2 55689 1 52
2 55690 1 52
2 55691 1 52
2 55692 1 52
2 55693 1 52
2 55694 1 52
2 55695 1 52
2 55696 1 52
2 55697 1 52
2 55698 1 52
2 55699 1 52
2 55700 1 52
2 55701 1 52
2 55702 1 52
2 55703 1 52
2 55704 1 52
2 55705 1 52
2 55706 1 52
2 55707 1 52
2 55708 1 52
2 55709 1 52
2 55710 1 52
2 55711 1 52
2 55712 1 52
2 55713 1 52
2 55714 1 52
2 55715 1 52
2 55716 1 52
2 55717 1 52
2 55718 1 52
2 55719 1 52
2 55720 1 52
2 55721 1 53
2 55722 1 53
2 55723 1 53
2 55724 1 53
2 55725 1 53
2 55726 1 53
2 55727 1 53
2 55728 1 53
2 55729 1 53
2 55730 1 53
2 55731 1 53
2 55732 1 53
2 55733 1 53
2 55734 1 53
2 55735 1 53
2 55736 1 53
2 55737 1 53
2 55738 1 53
2 55739 1 53
2 55740 1 53
2 55741 1 53
2 55742 1 53
2 55743 1 53
2 55744 1 53
2 55745 1 53
2 55746 1 53
2 55747 1 53
2 55748 1 53
2 55749 1 53
2 55750 1 53
2 55751 1 53
2 55752 1 53
2 55753 1 53
2 55754 1 53
2 55755 1 53
2 55756 1 53
2 55757 1 53
2 55758 1 53
2 55759 1 53
2 55760 1 53
2 55761 1 53
2 55762 1 53
2 55763 1 53
2 55764 1 53
2 55765 1 53
2 55766 1 53
2 55767 1 53
2 55768 1 53
2 55769 1 53
2 55770 1 53
2 55771 1 53
2 55772 1 53
2 55773 1 53
2 55774 1 53
2 55775 1 53
2 55776 1 53
2 55777 1 53
2 55778 1 53
2 55779 1 53
2 55780 1 53
2 55781 1 53
2 55782 1 53
2 55783 1 53
2 55784 1 53
2 55785 1 53
2 55786 1 53
2 55787 1 53
2 55788 1 53
2 55789 1 53
2 55790 1 53
2 55791 1 53
2 55792 1 53
2 55793 1 53
2 55794 1 53
2 55795 1 53
2 55796 1 53
2 55797 1 53
2 55798 1 53
2 55799 1 53
2 55800 1 53
2 55801 1 53
2 55802 1 53
2 55803 1 53
2 55804 1 53
2 55805 1 53
2 55806 1 53
2 55807 1 53
2 55808 1 53
2 55809 1 53
2 55810 1 53
2 55811 1 53
2 55812 1 53
2 55813 1 53
2 55814 1 53
2 55815 1 53
2 55816 1 53
2 55817 1 53
2 55818 1 53
2 55819 1 53
2 55820 1 53
2 55821 1 53
2 55822 1 53
2 55823 1 53
2 55824 1 53
2 55825 1 53
2 55826 1 53
2 55827 1 53
2 55828 1 53
2 55829 1 53
2 55830 1 53
2 55831 1 53
2 55832 1 53
2 55833 1 53
2 55834 1 53
2 55835 1 53
2 55836 1 53
2 55837 1 54
2 55838 1 54
2 55839 1 54
2 55840 1 54
2 55841 1 54
2 55842 1 54
2 55843 1 54
2 55844 1 54
2 55845 1 54
2 55846 1 54
2 55847 1 54
2 55848 1 54
2 55849 1 54
2 55850 1 54
2 55851 1 54
2 55852 1 54
2 55853 1 54
2 55854 1 54
2 55855 1 54
2 55856 1 54
2 55857 1 54
2 55858 1 54
2 55859 1 54
2 55860 1 54
2 55861 1 54
2 55862 1 54
2 55863 1 54
2 55864 1 54
2 55865 1 54
2 55866 1 54
2 55867 1 54
2 55868 1 54
2 55869 1 54
2 55870 1 54
2 55871 1 54
2 55872 1 54
2 55873 1 54
2 55874 1 54
2 55875 1 54
2 55876 1 54
2 55877 1 54
2 55878 1 54
2 55879 1 54
2 55880 1 54
2 55881 1 54
2 55882 1 54
2 55883 1 54
2 55884 1 54
2 55885 1 54
2 55886 1 54
2 55887 1 54
2 55888 1 54
2 55889 1 54
2 55890 1 54
2 55891 1 54
2 55892 1 54
2 55893 1 54
2 55894 1 54
2 55895 1 54
2 55896 1 54
2 55897 1 54
2 55898 1 54
2 55899 1 54
2 55900 1 54
2 55901 1 54
2 55902 1 54
2 55903 1 54
2 55904 1 54
2 55905 1 54
2 55906 1 54
2 55907 1 54
2 55908 1 54
2 55909 1 54
2 55910 1 54
2 55911 1 54
2 55912 1 54
2 55913 1 54
2 55914 1 54
2 55915 1 54
2 55916 1 54
2 55917 1 54
2 55918 1 54
2 55919 1 54
2 55920 1 54
2 55921 1 54
2 55922 1 54
2 55923 1 54
2 55924 1 54
2 55925 1 54
2 55926 1 54
2 55927 1 54
2 55928 1 54
2 55929 1 54
2 55930 1 54
2 55931 1 54
2 55932 1 54
2 55933 1 54
2 55934 1 54
2 55935 1 54
2 55936 1 54
2 55937 1 54
2 55938 1 54
2 55939 1 54
2 55940 1 54
2 55941 1 54
2 55942 1 54
2 55943 1 54
2 55944 1 54
2 55945 1 54
2 55946 1 54
2 55947 1 54
2 55948 1 54
2 55949 1 54
2 55950 1 54
2 55951 1 54
2 55952 1 54
2 55953 1 54
2 55954 1 54
2 55955 1 54
2 55956 1 54
2 55957 1 54
2 55958 1 54
2 55959 1 54
2 55960 1 54
2 55961 1 54
2 55962 1 54
2 55963 1 54
2 55964 1 54
2 55965 1 54
2 55966 1 54
2 55967 1 54
2 55968 1 54
2 55969 1 54
2 55970 1 54
2 55971 1 54
2 55972 1 55
2 55973 1 55
2 55974 1 55
2 55975 1 55
2 55976 1 55
2 55977 1 55
2 55978 1 55
2 55979 1 55
2 55980 1 55
2 55981 1 55
2 55982 1 55
2 55983 1 55
2 55984 1 55
2 55985 1 55
2 55986 1 55
2 55987 1 55
2 55988 1 55
2 55989 1 55
2 55990 1 55
2 55991 1 55
2 55992 1 55
2 55993 1 55
2 55994 1 55
2 55995 1 55
2 55996 1 55
2 55997 1 55
2 55998 1 55
2 55999 1 55
2 56000 1 55
2 56001 1 55
2 56002 1 55
2 56003 1 55
2 56004 1 55
2 56005 1 55
2 56006 1 55
2 56007 1 55
2 56008 1 55
2 56009 1 55
2 56010 1 55
2 56011 1 55
2 56012 1 55
2 56013 1 55
2 56014 1 55
2 56015 1 55
2 56016 1 55
2 56017 1 55
2 56018 1 55
2 56019 1 55
2 56020 1 55
2 56021 1 55
2 56022 1 55
2 56023 1 55
2 56024 1 55
2 56025 1 55
2 56026 1 55
2 56027 1 55
2 56028 1 55
2 56029 1 55
2 56030 1 55
2 56031 1 55
2 56032 1 55
2 56033 1 55
2 56034 1 55
2 56035 1 55
2 56036 1 55
2 56037 1 55
2 56038 1 55
2 56039 1 55
2 56040 1 55
2 56041 1 55
2 56042 1 55
2 56043 1 55
2 56044 1 55
2 56045 1 55
2 56046 1 55
2 56047 1 55
2 56048 1 55
2 56049 1 55
2 56050 1 55
2 56051 1 55
2 56052 1 55
2 56053 1 55
2 56054 1 55
2 56055 1 55
2 56056 1 55
2 56057 1 55
2 56058 1 55
2 56059 1 55
2 56060 1 55
2 56061 1 55
2 56062 1 55
2 56063 1 55
2 56064 1 55
2 56065 1 55
2 56066 1 55
2 56067 1 55
2 56068 1 55
2 56069 1 55
2 56070 1 55
2 56071 1 55
2 56072 1 55
2 56073 1 55
2 56074 1 55
2 56075 1 55
2 56076 1 55
2 56077 1 55
2 56078 1 55
2 56079 1 55
2 56080 1 55
2 56081 1 55
2 56082 1 55
2 56083 1 55
2 56084 1 55
2 56085 1 55
2 56086 1 55
2 56087 1 55
2 56088 1 55
2 56089 1 55
2 56090 1 55
2 56091 1 55
2 56092 1 55
2 56093 1 55
2 56094 1 55
2 56095 1 55
2 56096 1 55
2 56097 1 55
2 56098 1 55
2 56099 1 55
2 56100 1 55
2 56101 1 55
2 56102 1 55
2 56103 1 55
2 56104 1 55
2 56105 1 55
2 56106 1 55
2 56107 1 55
2 56108 1 55
2 56109 1 55
2 56110 1 55
2 56111 1 55
2 56112 1 55
2 56113 1 55
2 56114 1 55
2 56115 1 55
2 56116 1 55
2 56117 1 55
2 56118 1 55
2 56119 1 55
2 56120 1 55
2 56121 1 55
2 56122 1 55
2 56123 1 55
2 56124 1 55
2 56125 1 55
2 56126 1 55
2 56127 1 55
2 56128 1 55
2 56129 1 55
2 56130 1 55
2 56131 1 55
2 56132 1 55
2 56133 1 55
2 56134 1 55
2 56135 1 55
2 56136 1 55
2 56137 1 55
2 56138 1 55
2 56139 1 55
2 56140 1 55
2 56141 1 55
2 56142 1 55
2 56143 1 55
2 56144 1 55
2 56145 1 55
2 56146 1 55
2 56147 1 55
2 56148 1 55
2 56149 1 55
2 56150 1 55
2 56151 1 55
2 56152 1 55
2 56153 1 55
2 56154 1 55
2 56155 1 55
2 56156 1 55
2 56157 1 55
2 56158 1 55
2 56159 1 55
2 56160 1 55
2 56161 1 55
2 56162 1 55
2 56163 1 55
2 56164 1 55
2 56165 1 55
2 56166 1 55
2 56167 1 55
2 56168 1 55
2 56169 1 55
2 56170 1 56
2 56171 1 56
2 56172 1 56
2 56173 1 56
2 56174 1 56
2 56175 1 56
2 56176 1 56
2 56177 1 56
2 56178 1 56
2 56179 1 56
2 56180 1 56
2 56181 1 56
2 56182 1 56
2 56183 1 56
2 56184 1 56
2 56185 1 56
2 56186 1 56
2 56187 1 56
2 56188 1 56
2 56189 1 56
2 56190 1 56
2 56191 1 56
2 56192 1 56
2 56193 1 56
2 56194 1 56
2 56195 1 56
2 56196 1 56
2 56197 1 56
2 56198 1 56
2 56199 1 56
2 56200 1 56
2 56201 1 56
2 56202 1 56
2 56203 1 56
2 56204 1 56
2 56205 1 56
2 56206 1 56
2 56207 1 56
2 56208 1 56
2 56209 1 56
2 56210 1 56
2 56211 1 56
2 56212 1 56
2 56213 1 56
2 56214 1 56
2 56215 1 56
2 56216 1 56
2 56217 1 56
2 56218 1 56
2 56219 1 56
2 56220 1 56
2 56221 1 56
2 56222 1 56
2 56223 1 56
2 56224 1 56
2 56225 1 56
2 56226 1 56
2 56227 1 56
2 56228 1 56
2 56229 1 56
2 56230 1 56
2 56231 1 56
2 56232 1 56
2 56233 1 56
2 56234 1 56
2 56235 1 56
2 56236 1 56
2 56237 1 56
2 56238 1 56
2 56239 1 56
2 56240 1 56
2 56241 1 56
2 56242 1 56
2 56243 1 56
2 56244 1 56
2 56245 1 56
2 56246 1 56
2 56247 1 56
2 56248 1 56
2 56249 1 56
2 56250 1 56
2 56251 1 56
2 56252 1 56
2 56253 1 56
2 56254 1 56
2 56255 1 56
2 56256 1 56
2 56257 1 56
2 56258 1 56
2 56259 1 56
2 56260 1 56
2 56261 1 56
2 56262 1 56
2 56263 1 56
2 56264 1 56
2 56265 1 56
2 56266 1 56
2 56267 1 56
2 56268 1 56
2 56269 1 57
2 56270 1 57
2 56271 1 57
2 56272 1 57
2 56273 1 57
2 56274 1 57
2 56275 1 57
2 56276 1 57
2 56277 1 57
2 56278 1 57
2 56279 1 57
2 56280 1 57
2 56281 1 57
2 56282 1 57
2 56283 1 57
2 56284 1 57
2 56285 1 57
2 56286 1 57
2 56287 1 57
2 56288 1 57
2 56289 1 57
2 56290 1 57
2 56291 1 57
2 56292 1 57
2 56293 1 57
2 56294 1 57
2 56295 1 57
2 56296 1 57
2 56297 1 57
2 56298 1 57
2 56299 1 57
2 56300 1 57
2 56301 1 57
2 56302 1 57
2 56303 1 57
2 56304 1 57
2 56305 1 57
2 56306 1 57
2 56307 1 57
2 56308 1 57
2 56309 1 57
2 56310 1 57
2 56311 1 57
2 56312 1 57
2 56313 1 57
2 56314 1 57
2 56315 1 57
2 56316 1 57
2 56317 1 57
2 56318 1 57
2 56319 1 57
2 56320 1 57
2 56321 1 57
2 56322 1 57
2 56323 1 57
2 56324 1 57
2 56325 1 57
2 56326 1 57
2 56327 1 57
2 56328 1 57
2 56329 1 57
2 56330 1 57
2 56331 1 57
2 56332 1 57
2 56333 1 57
2 56334 1 57
2 56335 1 57
2 56336 1 57
2 56337 1 57
2 56338 1 57
2 56339 1 57
2 56340 1 57
2 56341 1 57
2 56342 1 57
2 56343 1 57
2 56344 1 57
2 56345 1 57
2 56346 1 57
2 56347 1 57
2 56348 1 57
2 56349 1 57
2 56350 1 57
2 56351 1 57
2 56352 1 57
2 56353 1 57
2 56354 1 57
2 56355 1 57
2 56356 1 57
2 56357 1 57
2 56358 1 57
2 56359 1 57
2 56360 1 57
2 56361 1 57
2 56362 1 57
2 56363 1 57
2 56364 1 57
2 56365 1 57
2 56366 1 57
2 56367 1 57
2 56368 1 57
2 56369 1 57
2 56370 1 57
2 56371 1 57
2 56372 1 57
2 56373 1 57
2 56374 1 57
2 56375 1 57
2 56376 1 57
2 56377 1 57
2 56378 1 57
2 56379 1 57
2 56380 1 57
2 56381 1 57
2 56382 1 57
2 56383 1 57
2 56384 1 57
2 56385 1 57
2 56386 1 57
2 56387 1 57
2 56388 1 57
2 56389 1 57
2 56390 1 57
2 56391 1 57
2 56392 1 57
2 56393 1 57
2 56394 1 57
2 56395 1 57
2 56396 1 57
2 56397 1 57
2 56398 1 57
2 56399 1 57
2 56400 1 57
2 56401 1 57
2 56402 1 57
2 56403 1 57
2 56404 1 57
2 56405 1 57
2 56406 1 57
2 56407 1 57
2 56408 1 57
2 56409 1 57
2 56410 1 57
2 56411 1 57
2 56412 1 57
2 56413 1 57
2 56414 1 57
2 56415 1 57
2 56416 1 57
2 56417 1 57
2 56418 1 57
2 56419 1 57
2 56420 1 57
2 56421 1 57
2 56422 1 57
2 56423 1 57
2 56424 1 57
2 56425 1 57
2 56426 1 57
2 56427 1 57
2 56428 1 57
2 56429 1 57
2 56430 1 57
2 56431 1 58
2 56432 1 58
2 56433 1 58
2 56434 1 58
2 56435 1 58
2 56436 1 58
2 56437 1 58
2 56438 1 58
2 56439 1 58
2 56440 1 58
2 56441 1 58
2 56442 1 58
2 56443 1 58
2 56444 1 58
2 56445 1 58
2 56446 1 58
2 56447 1 58
2 56448 1 58
2 56449 1 58
2 56450 1 58
2 56451 1 58
2 56452 1 58
2 56453 1 58
2 56454 1 58
2 56455 1 58
2 56456 1 58
2 56457 1 58
2 56458 1 58
2 56459 1 58
2 56460 1 58
2 56461 1 58
2 56462 1 58
2 56463 1 58
2 56464 1 58
2 56465 1 58
2 56466 1 58
2 56467 1 58
2 56468 1 58
2 56469 1 58
2 56470 1 58
2 56471 1 58
2 56472 1 58
2 56473 1 58
2 56474 1 58
2 56475 1 58
2 56476 1 58
2 56477 1 58
2 56478 1 58
2 56479 1 58
2 56480 1 58
2 56481 1 58
2 56482 1 58
2 56483 1 58
2 56484 1 58
2 56485 1 58
2 56486 1 59
2 56487 1 59
2 56488 1 59
2 56489 1 59
2 56490 1 59
2 56491 1 59
2 56492 1 59
2 56493 1 59
2 56494 1 59
2 56495 1 59
2 56496 1 59
2 56497 1 59
2 56498 1 59
2 56499 1 59
2 56500 1 59
2 56501 1 59
2 56502 1 59
2 56503 1 59
2 56504 1 59
2 56505 1 59
2 56506 1 59
2 56507 1 59
2 56508 1 59
2 56509 1 59
2 56510 1 59
2 56511 1 59
2 56512 1 59
2 56513 1 59
2 56514 1 59
2 56515 1 59
2 56516 1 59
2 56517 1 59
2 56518 1 59
2 56519 1 59
2 56520 1 59
2 56521 1 59
2 56522 1 59
2 56523 1 59
2 56524 1 59
2 56525 1 59
2 56526 1 59
2 56527 1 59
2 56528 1 59
2 56529 1 59
2 56530 1 59
2 56531 1 59
2 56532 1 59
2 56533 1 59
2 56534 1 59
2 56535 1 59
2 56536 1 59
2 56537 1 59
2 56538 1 59
2 56539 1 59
2 56540 1 59
2 56541 1 59
2 56542 1 59
2 56543 1 59
2 56544 1 59
2 56545 1 59
2 56546 1 59
2 56547 1 59
2 56548 1 59
2 56549 1 59
2 56550 1 59
2 56551 1 59
2 56552 1 59
2 56553 1 59
2 56554 1 59
2 56555 1 59
2 56556 1 59
2 56557 1 59
2 56558 1 59
2 56559 1 59
2 56560 1 59
2 56561 1 59
2 56562 1 59
2 56563 1 59
2 56564 1 59
2 56565 1 59
2 56566 1 59
2 56567 1 59
2 56568 1 59
2 56569 1 59
2 56570 1 59
2 56571 1 59
2 56572 1 59
2 56573 1 59
2 56574 1 59
2 56575 1 59
2 56576 1 59
2 56577 1 59
2 56578 1 59
2 56579 1 59
2 56580 1 59
2 56581 1 59
2 56582 1 59
2 56583 1 59
2 56584 1 59
2 56585 1 59
2 56586 1 59
2 56587 1 59
2 56588 1 59
2 56589 1 59
2 56590 1 59
2 56591 1 59
2 56592 1 59
2 56593 1 59
2 56594 1 59
2 56595 1 59
2 56596 1 59
2 56597 1 59
2 56598 1 59
2 56599 1 59
2 56600 1 59
2 56601 1 60
2 56602 1 60
2 56603 1 60
2 56604 1 60
2 56605 1 60
2 56606 1 60
2 56607 1 60
2 56608 1 60
2 56609 1 60
2 56610 1 60
2 56611 1 60
2 56612 1 60
2 56613 1 60
2 56614 1 60
2 56615 1 60
2 56616 1 60
2 56617 1 60
2 56618 1 60
2 56619 1 60
2 56620 1 60
2 56621 1 60
2 56622 1 60
2 56623 1 60
2 56624 1 60
2 56625 1 60
2 56626 1 60
2 56627 1 60
2 56628 1 60
2 56629 1 60
2 56630 1 60
2 56631 1 60
2 56632 1 60
2 56633 1 60
2 56634 1 60
2 56635 1 60
2 56636 1 60
2 56637 1 60
2 56638 1 60
2 56639 1 60
2 56640 1 60
2 56641 1 60
2 56642 1 60
2 56643 1 60
2 56644 1 60
2 56645 1 60
2 56646 1 60
2 56647 1 60
2 56648 1 60
2 56649 1 60
2 56650 1 60
2 56651 1 60
2 56652 1 60
2 56653 1 60
2 56654 1 60
2 56655 1 60
2 56656 1 60
2 56657 1 60
2 56658 1 60
2 56659 1 60
2 56660 1 60
2 56661 1 60
2 56662 1 60
2 56663 1 60
2 56664 1 60
2 56665 1 60
2 56666 1 60
2 56667 1 60
2 56668 1 60
2 56669 1 61
2 56670 1 61
2 56671 1 61
2 56672 1 61
2 56673 1 61
2 56674 1 61
2 56675 1 61
2 56676 1 61
2 56677 1 61
2 56678 1 61
2 56679 1 61
2 56680 1 61
2 56681 1 61
2 56682 1 61
2 56683 1 61
2 56684 1 61
2 56685 1 61
2 56686 1 61
2 56687 1 61
2 56688 1 61
2 56689 1 61
2 56690 1 61
2 56691 1 61
2 56692 1 61
2 56693 1 61
2 56694 1 61
2 56695 1 61
2 56696 1 61
2 56697 1 61
2 56698 1 61
2 56699 1 61
2 56700 1 61
2 56701 1 61
2 56702 1 61
2 56703 1 61
2 56704 1 61
2 56705 1 61
2 56706 1 61
2 56707 1 61
2 56708 1 61
2 56709 1 61
2 56710 1 61
2 56711 1 61
2 56712 1 61
2 56713 1 61
2 56714 1 61
2 56715 1 61
2 56716 1 61
2 56717 1 61
2 56718 1 61
2 56719 1 61
2 56720 1 61
2 56721 1 61
2 56722 1 61
2 56723 1 61
2 56724 1 61
2 56725 1 61
2 56726 1 61
2 56727 1 61
2 56728 1 61
2 56729 1 61
2 56730 1 61
2 56731 1 61
2 56732 1 61
2 56733 1 61
2 56734 1 61
2 56735 1 61
2 56736 1 61
2 56737 1 61
2 56738 1 61
2 56739 1 61
2 56740 1 61
2 56741 1 61
2 56742 1 61
2 56743 1 61
2 56744 1 61
2 56745 1 61
2 56746 1 61
2 56747 1 61
2 56748 1 61
2 56749 1 61
2 56750 1 61
2 56751 1 61
2 56752 1 61
2 56753 1 61
2 56754 1 61
2 56755 1 61
2 56756 1 61
2 56757 1 61
2 56758 1 61
2 56759 1 61
2 56760 1 61
2 56761 1 61
2 56762 1 61
2 56763 1 61
2 56764 1 61
2 56765 1 61
2 56766 1 61
2 56767 1 61
2 56768 1 61
2 56769 1 61
2 56770 1 61
2 56771 1 61
2 56772 1 61
2 56773 1 61
2 56774 1 61
2 56775 1 61
2 56776 1 61
2 56777 1 61
2 56778 1 61
2 56779 1 61
2 56780 1 61
2 56781 1 61
2 56782 1 62
2 56783 1 62
2 56784 1 64
2 56785 1 64
2 56786 1 65
2 56787 1 65
2 56788 1 66
2 56789 1 66
2 56790 1 66
2 56791 1 66
2 56792 1 66
2 56793 1 66
2 56794 1 66
2 56795 1 66
2 56796 1 66
2 56797 1 66
2 56798 1 66
2 56799 1 66
2 56800 1 66
2 56801 1 66
2 56802 1 66
2 56803 1 66
2 56804 1 66
2 56805 1 66
2 56806 1 66
2 56807 1 66
2 56808 1 66
2 56809 1 66
2 56810 1 66
2 56811 1 66
2 56812 1 66
2 56813 1 66
2 56814 1 66
2 56815 1 66
2 56816 1 66
2 56817 1 66
2 56818 1 66
2 56819 1 66
2 56820 1 66
2 56821 1 66
2 56822 1 66
2 56823 1 66
2 56824 1 66
2 56825 1 66
2 56826 1 66
2 56827 1 66
2 56828 1 66
2 56829 1 66
2 56830 1 66
2 56831 1 66
2 56832 1 66
2 56833 1 66
2 56834 1 66
2 56835 1 66
2 56836 1 66
2 56837 1 66
2 56838 1 66
2 56839 1 66
2 56840 1 66
2 56841 1 66
2 56842 1 66
2 56843 1 66
2 56844 1 66
2 56845 1 66
2 56846 1 66
2 56847 1 66
2 56848 1 66
2 56849 1 66
2 56850 1 66
2 56851 1 66
2 56852 1 66
2 56853 1 66
2 56854 1 66
2 56855 1 66
2 56856 1 66
2 56857 1 66
2 56858 1 66
2 56859 1 66
2 56860 1 66
2 56861 1 66
2 56862 1 66
2 56863 1 66
2 56864 1 66
2 56865 1 66
2 56866 1 66
2 56867 1 66
2 56868 1 66
2 56869 1 66
2 56870 1 66
2 56871 1 66
2 56872 1 66
2 56873 1 66
2 56874 1 66
2 56875 1 66
2 56876 1 66
2 56877 1 66
2 56878 1 66
2 56879 1 66
2 56880 1 66
2 56881 1 66
2 56882 1 66
2 56883 1 66
2 56884 1 66
2 56885 1 66
2 56886 1 66
2 56887 1 66
2 56888 1 66
2 56889 1 66
2 56890 1 66
2 56891 1 66
2 56892 1 66
2 56893 1 66
2 56894 1 66
2 56895 1 66
2 56896 1 66
2 56897 1 66
2 56898 1 66
2 56899 1 66
2 56900 1 66
2 56901 1 66
2 56902 1 66
2 56903 1 66
2 56904 1 66
2 56905 1 66
2 56906 1 66
2 56907 1 66
2 56908 1 66
2 56909 1 66
2 56910 1 66
2 56911 1 66
2 56912 1 66
2 56913 1 66
2 56914 1 66
2 56915 1 66
2 56916 1 66
2 56917 1 66
2 56918 1 66
2 56919 1 66
2 56920 1 66
2 56921 1 66
2 56922 1 66
2 56923 1 66
2 56924 1 66
2 56925 1 66
2 56926 1 66
2 56927 1 66
2 56928 1 66
2 56929 1 66
2 56930 1 66
2 56931 1 66
2 56932 1 66
2 56933 1 66
2 56934 1 66
2 56935 1 66
2 56936 1 66
2 56937 1 66
2 56938 1 66
2 56939 1 66
2 56940 1 66
2 56941 1 66
2 56942 1 66
2 56943 1 66
2 56944 1 66
2 56945 1 66
2 56946 1 66
2 56947 1 66
2 56948 1 66
2 56949 1 66
2 56950 1 66
2 56951 1 66
2 56952 1 66
2 56953 1 66
2 56954 1 66
2 56955 1 66
2 56956 1 66
2 56957 1 66
2 56958 1 66
2 56959 1 66
2 56960 1 66
2 56961 1 66
2 56962 1 66
2 56963 1 66
2 56964 1 66
2 56965 1 66
2 56966 1 66
2 56967 1 66
2 56968 1 66
2 56969 1 66
2 56970 1 66
2 56971 1 67
2 56972 1 67
2 56973 1 67
2 56974 1 67
2 56975 1 67
2 56976 1 67
2 56977 1 67
2 56978 1 67
2 56979 1 67
2 56980 1 67
2 56981 1 67
2 56982 1 67
2 56983 1 67
2 56984 1 67
2 56985 1 67
2 56986 1 67
2 56987 1 67
2 56988 1 67
2 56989 1 67
2 56990 1 67
2 56991 1 67
2 56992 1 67
2 56993 1 67
2 56994 1 67
2 56995 1 67
2 56996 1 67
2 56997 1 67
2 56998 1 67
2 56999 1 67
2 57000 1 67
2 57001 1 67
2 57002 1 67
2 57003 1 67
2 57004 1 67
2 57005 1 67
2 57006 1 67
2 57007 1 67
2 57008 1 67
2 57009 1 67
2 57010 1 67
2 57011 1 67
2 57012 1 67
2 57013 1 67
2 57014 1 67
2 57015 1 67
2 57016 1 67
2 57017 1 67
2 57018 1 67
2 57019 1 67
2 57020 1 67
2 57021 1 67
2 57022 1 67
2 57023 1 67
2 57024 1 67
2 57025 1 67
2 57026 1 67
2 57027 1 67
2 57028 1 67
2 57029 1 67
2 57030 1 67
2 57031 1 67
2 57032 1 67
2 57033 1 67
2 57034 1 67
2 57035 1 67
2 57036 1 67
2 57037 1 67
2 57038 1 67
2 57039 1 67
2 57040 1 67
2 57041 1 67
2 57042 1 67
2 57043 1 67
2 57044 1 67
2 57045 1 67
2 57046 1 67
2 57047 1 67
2 57048 1 67
2 57049 1 67
2 57050 1 67
2 57051 1 67
2 57052 1 67
2 57053 1 67
2 57054 1 67
2 57055 1 67
2 57056 1 67
2 57057 1 67
2 57058 1 67
2 57059 1 67
2 57060 1 67
2 57061 1 67
2 57062 1 67
2 57063 1 67
2 57064 1 67
2 57065 1 67
2 57066 1 67
2 57067 1 67
2 57068 1 67
2 57069 1 67
2 57070 1 67
2 57071 1 67
2 57072 1 67
2 57073 1 67
2 57074 1 68
2 57075 1 68
2 57076 1 68
2 57077 1 68
2 57078 1 69
2 57079 1 69
2 57080 1 69
2 57081 1 69
2 57082 1 69
2 57083 1 69
2 57084 1 69
2 57085 1 69
2 57086 1 69
2 57087 1 69
2 57088 1 69
2 57089 1 69
2 57090 1 69
2 57091 1 69
2 57092 1 69
2 57093 1 69
2 57094 1 69
2 57095 1 69
2 57096 1 69
2 57097 1 69
2 57098 1 69
2 57099 1 69
2 57100 1 69
2 57101 1 69
2 57102 1 69
2 57103 1 69
2 57104 1 69
2 57105 1 69
2 57106 1 69
2 57107 1 69
2 57108 1 69
2 57109 1 69
2 57110 1 69
2 57111 1 69
2 57112 1 69
2 57113 1 69
2 57114 1 69
2 57115 1 70
2 57116 1 70
2 57117 1 70
2 57118 1 70
2 57119 1 70
2 57120 1 70
2 57121 1 70
2 57122 1 70
2 57123 1 70
2 57124 1 70
2 57125 1 70
2 57126 1 70
2 57127 1 70
2 57128 1 70
2 57129 1 70
2 57130 1 70
2 57131 1 70
2 57132 1 70
2 57133 1 70
2 57134 1 70
2 57135 1 70
2 57136 1 70
2 57137 1 70
2 57138 1 70
2 57139 1 70
2 57140 1 70
2 57141 1 70
2 57142 1 70
2 57143 1 70
2 57144 1 70
2 57145 1 70
2 57146 1 70
2 57147 1 70
2 57148 1 70
2 57149 1 70
2 57150 1 70
2 57151 1 70
2 57152 1 70
2 57153 1 70
2 57154 1 70
2 57155 1 70
2 57156 1 70
2 57157 1 70
2 57158 1 70
2 57159 1 70
2 57160 1 70
2 57161 1 70
2 57162 1 70
2 57163 1 70
2 57164 1 70
2 57165 1 70
2 57166 1 70
2 57167 1 70
2 57168 1 70
2 57169 1 70
2 57170 1 70
2 57171 1 70
2 57172 1 70
2 57173 1 70
2 57174 1 70
2 57175 1 70
2 57176 1 70
2 57177 1 70
2 57178 1 70
2 57179 1 70
2 57180 1 70
2 57181 1 70
2 57182 1 70
2 57183 1 70
2 57184 1 70
2 57185 1 70
2 57186 1 70
2 57187 1 70
2 57188 1 70
2 57189 1 70
2 57190 1 70
2 57191 1 70
2 57192 1 71
2 57193 1 71
2 57194 1 71
2 57195 1 71
2 57196 1 71
2 57197 1 71
2 57198 1 71
2 57199 1 71
2 57200 1 71
2 57201 1 71
2 57202 1 71
2 57203 1 71
2 57204 1 71
2 57205 1 71
2 57206 1 71
2 57207 1 71
2 57208 1 71
2 57209 1 71
2 57210 1 71
2 57211 1 71
2 57212 1 71
2 57213 1 71
2 57214 1 71
2 57215 1 71
2 57216 1 71
2 57217 1 71
2 57218 1 71
2 57219 1 71
2 57220 1 71
2 57221 1 71
2 57222 1 71
2 57223 1 71
2 57224 1 71
2 57225 1 71
2 57226 1 71
2 57227 1 71
2 57228 1 71
2 57229 1 71
2 57230 1 71
2 57231 1 71
2 57232 1 71
2 57233 1 71
2 57234 1 71
2 57235 1 71
2 57236 1 71
2 57237 1 71
2 57238 1 71
2 57239 1 71
2 57240 1 71
2 57241 1 71
2 57242 1 71
2 57243 1 71
2 57244 1 71
2 57245 1 71
2 57246 1 71
2 57247 1 71
2 57248 1 71
2 57249 1 71
2 57250 1 71
2 57251 1 71
2 57252 1 71
2 57253 1 71
2 57254 1 71
2 57255 1 71
2 57256 1 71
2 57257 1 71
2 57258 1 71
2 57259 1 71
2 57260 1 71
2 57261 1 71
2 57262 1 71
2 57263 1 71
2 57264 1 71
2 57265 1 71
2 57266 1 71
2 57267 1 71
2 57268 1 71
2 57269 1 71
2 57270 1 72
2 57271 1 72
2 57272 1 73
2 57273 1 73
2 57274 1 73
2 57275 1 73
2 57276 1 73
2 57277 1 73
2 57278 1 73
2 57279 1 73
2 57280 1 73
2 57281 1 73
2 57282 1 73
2 57283 1 73
2 57284 1 73
2 57285 1 73
2 57286 1 73
2 57287 1 73
2 57288 1 74
2 57289 1 74
2 57290 1 74
2 57291 1 81
2 57292 1 81
2 57293 1 81
2 57294 1 81
2 57295 1 81
2 57296 1 81
2 57297 1 81
2 57298 1 83
2 57299 1 83
2 57300 1 83
2 57301 1 83
2 57302 1 88
2 57303 1 88
2 57304 1 88
2 57305 1 88
2 57306 1 88
2 57307 1 88
2 57308 1 89
2 57309 1 89
2 57310 1 89
2 57311 1 89
2 57312 1 89
2 57313 1 89
2 57314 1 89
2 57315 1 89
2 57316 1 89
2 57317 1 89
2 57318 1 89
2 57319 1 89
2 57320 1 89
2 57321 1 89
2 57322 1 89
2 57323 1 89
2 57324 1 89
2 57325 1 89
2 57326 1 89
2 57327 1 89
2 57328 1 89
2 57329 1 89
2 57330 1 89
2 57331 1 89
2 57332 1 89
2 57333 1 89
2 57334 1 89
2 57335 1 89
2 57336 1 89
2 57337 1 89
2 57338 1 89
2 57339 1 89
2 57340 1 89
2 57341 1 89
2 57342 1 89
2 57343 1 89
2 57344 1 89
2 57345 1 89
2 57346 1 89
2 57347 1 89
2 57348 1 89
2 57349 1 90
2 57350 1 90
2 57351 1 90
2 57352 1 90
2 57353 1 91
2 57354 1 91
2 57355 1 91
2 57356 1 91
2 57357 1 91
2 57358 1 92
2 57359 1 92
2 57360 1 92
2 57361 1 92
2 57362 1 92
2 57363 1 92
2 57364 1 92
2 57365 1 92
2 57366 1 92
2 57367 1 92
2 57368 1 93
2 57369 1 93
2 57370 1 93
2 57371 1 93
2 57372 1 93
2 57373 1 93
2 57374 1 93
2 57375 1 93
2 57376 1 93
2 57377 1 93
2 57378 1 93
2 57379 1 93
2 57380 1 94
2 57381 1 94
2 57382 1 94
2 57383 1 94
2 57384 1 94
2 57385 1 94
2 57386 1 94
2 57387 1 94
2 57388 1 94
2 57389 1 94
2 57390 1 94
2 57391 1 94
2 57392 1 94
2 57393 1 94
2 57394 1 94
2 57395 1 94
2 57396 1 94
2 57397 1 94
2 57398 1 94
2 57399 1 94
2 57400 1 94
2 57401 1 94
2 57402 1 94
2 57403 1 94
2 57404 1 94
2 57405 1 94
2 57406 1 94
2 57407 1 94
2 57408 1 94
2 57409 1 94
2 57410 1 94
2 57411 1 94
2 57412 1 94
2 57413 1 94
2 57414 1 94
2 57415 1 94
2 57416 1 94
2 57417 1 94
2 57418 1 94
2 57419 1 94
2 57420 1 94
2 57421 1 94
2 57422 1 94
2 57423 1 94
2 57424 1 94
2 57425 1 94
2 57426 1 94
2 57427 1 94
2 57428 1 94
2 57429 1 94
2 57430 1 94
2 57431 1 94
2 57432 1 94
2 57433 1 94
2 57434 1 94
2 57435 1 94
2 57436 1 94
2 57437 1 94
2 57438 1 94
2 57439 1 94
2 57440 1 94
2 57441 1 94
2 57442 1 94
2 57443 1 94
2 57444 1 94
2 57445 1 94
2 57446 1 94
2 57447 1 94
2 57448 1 94
2 57449 1 94
2 57450 1 94
2 57451 1 94
2 57452 1 94
2 57453 1 94
2 57454 1 94
2 57455 1 94
2 57456 1 94
2 57457 1 94
2 57458 1 94
2 57459 1 94
2 57460 1 94
2 57461 1 94
2 57462 1 94
2 57463 1 94
2 57464 1 94
2 57465 1 94
2 57466 1 94
2 57467 1 94
2 57468 1 94
2 57469 1 94
2 57470 1 94
2 57471 1 94
2 57472 1 94
2 57473 1 94
2 57474 1 94
2 57475 1 94
2 57476 1 94
2 57477 1 94
2 57478 1 94
2 57479 1 94
2 57480 1 94
2 57481 1 94
2 57482 1 94
2 57483 1 94
2 57484 1 94
2 57485 1 94
2 57486 1 94
2 57487 1 94
2 57488 1 94
2 57489 1 94
2 57490 1 94
2 57491 1 94
2 57492 1 94
2 57493 1 94
2 57494 1 94
2 57495 1 94
2 57496 1 94
2 57497 1 94
2 57498 1 94
2 57499 1 94
2 57500 1 94
2 57501 1 94
2 57502 1 94
2 57503 1 94
2 57504 1 94
2 57505 1 94
2 57506 1 94
2 57507 1 94
2 57508 1 94
2 57509 1 94
2 57510 1 94
2 57511 1 94
2 57512 1 94
2 57513 1 94
2 57514 1 94
2 57515 1 94
2 57516 1 94
2 57517 1 94
2 57518 1 94
2 57519 1 94
2 57520 1 94
2 57521 1 94
2 57522 1 94
2 57523 1 94
2 57524 1 94
2 57525 1 94
2 57526 1 94
2 57527 1 94
2 57528 1 94
2 57529 1 94
2 57530 1 94
2 57531 1 94
2 57532 1 94
2 57533 1 94
2 57534 1 94
2 57535 1 94
2 57536 1 94
2 57537 1 94
2 57538 1 94
2 57539 1 94
2 57540 1 94
2 57541 1 94
2 57542 1 94
2 57543 1 94
2 57544 1 94
2 57545 1 94
2 57546 1 94
2 57547 1 94
2 57548 1 94
2 57549 1 94
2 57550 1 95
2 57551 1 95
2 57552 1 95
2 57553 1 95
2 57554 1 95
2 57555 1 95
2 57556 1 95
2 57557 1 95
2 57558 1 95
2 57559 1 95
2 57560 1 95
2 57561 1 95
2 57562 1 95
2 57563 1 95
2 57564 1 95
2 57565 1 95
2 57566 1 95
2 57567 1 95
2 57568 1 95
2 57569 1 95
2 57570 1 95
2 57571 1 95
2 57572 1 95
2 57573 1 95
2 57574 1 95
2 57575 1 95
2 57576 1 95
2 57577 1 95
2 57578 1 95
2 57579 1 95
2 57580 1 95
2 57581 1 95
2 57582 1 95
2 57583 1 95
2 57584 1 95
2 57585 1 95
2 57586 1 95
2 57587 1 95
2 57588 1 95
2 57589 1 95
2 57590 1 95
2 57591 1 95
2 57592 1 95
2 57593 1 95
2 57594 1 95
2 57595 1 95
2 57596 1 95
2 57597 1 95
2 57598 1 95
2 57599 1 95
2 57600 1 95
2 57601 1 95
2 57602 1 95
2 57603 1 95
2 57604 1 95
2 57605 1 95
2 57606 1 95
2 57607 1 95
2 57608 1 95
2 57609 1 95
2 57610 1 95
2 57611 1 95
2 57612 1 95
2 57613 1 95
2 57614 1 95
2 57615 1 95
2 57616 1 95
2 57617 1 95
2 57618 1 95
2 57619 1 95
2 57620 1 95
2 57621 1 95
2 57622 1 95
2 57623 1 95
2 57624 1 95
2 57625 1 95
2 57626 1 95
2 57627 1 95
2 57628 1 95
2 57629 1 95
2 57630 1 95
2 57631 1 95
2 57632 1 95
2 57633 1 95
2 57634 1 95
2 57635 1 95
2 57636 1 95
2 57637 1 95
2 57638 1 95
2 57639 1 95
2 57640 1 95
2 57641 1 95
2 57642 1 95
2 57643 1 95
2 57644 1 95
2 57645 1 95
2 57646 1 95
2 57647 1 95
2 57648 1 95
2 57649 1 95
2 57650 1 95
2 57651 1 95
2 57652 1 95
2 57653 1 95
2 57654 1 95
2 57655 1 95
2 57656 1 95
2 57657 1 95
2 57658 1 95
2 57659 1 95
2 57660 1 95
2 57661 1 95
2 57662 1 95
2 57663 1 95
2 57664 1 95
2 57665 1 95
2 57666 1 95
2 57667 1 95
2 57668 1 95
2 57669 1 95
2 57670 1 95
2 57671 1 95
2 57672 1 95
2 57673 1 95
2 57674 1 95
2 57675 1 95
2 57676 1 95
2 57677 1 95
2 57678 1 95
2 57679 1 95
2 57680 1 95
2 57681 1 95
2 57682 1 95
2 57683 1 95
2 57684 1 95
2 57685 1 95
2 57686 1 95
2 57687 1 95
2 57688 1 95
2 57689 1 95
2 57690 1 95
2 57691 1 95
2 57692 1 95
2 57693 1 95
2 57694 1 95
2 57695 1 95
2 57696 1 95
2 57697 1 95
2 57698 1 95
2 57699 1 95
2 57700 1 95
2 57701 1 95
2 57702 1 95
2 57703 1 95
2 57704 1 95
2 57705 1 95
2 57706 1 95
2 57707 1 95
2 57708 1 95
2 57709 1 95
2 57710 1 95
2 57711 1 95
2 57712 1 96
2 57713 1 96
2 57714 1 97
2 57715 1 97
2 57716 1 99
2 57717 1 99
2 57718 1 99
2 57719 1 99
2 57720 1 99
2 57721 1 99
2 57722 1 99
2 57723 1 99
2 57724 1 99
2 57725 1 99
2 57726 1 99
2 57727 1 99
2 57728 1 100
2 57729 1 100
2 57730 1 100
2 57731 1 100
2 57732 1 100
2 57733 1 100
2 57734 1 100
2 57735 1 100
2 57736 1 100
2 57737 1 100
2 57738 1 100
2 57739 1 100
2 57740 1 100
2 57741 1 100
2 57742 1 100
2 57743 1 100
2 57744 1 100
2 57745 1 100
2 57746 1 100
2 57747 1 100
2 57748 1 100
2 57749 1 100
2 57750 1 101
2 57751 1 101
2 57752 1 101
2 57753 1 101
2 57754 1 101
2 57755 1 101
2 57756 1 101
2 57757 1 101
2 57758 1 101
2 57759 1 101
2 57760 1 102
2 57761 1 102
2 57762 1 102
2 57763 1 102
2 57764 1 102
2 57765 1 102
2 57766 1 102
2 57767 1 102
2 57768 1 102
2 57769 1 102
2 57770 1 102
2 57771 1 102
2 57772 1 102
2 57773 1 102
2 57774 1 102
2 57775 1 102
2 57776 1 102
2 57777 1 103
2 57778 1 103
2 57779 1 103
2 57780 1 103
2 57781 1 103
2 57782 1 103
2 57783 1 103
2 57784 1 103
2 57785 1 103
2 57786 1 104
2 57787 1 104
2 57788 1 105
2 57789 1 105
2 57790 1 105
2 57791 1 105
2 57792 1 105
2 57793 1 105
2 57794 1 110
2 57795 1 110
2 57796 1 110
2 57797 1 110
2 57798 1 110
2 57799 1 110
2 57800 1 111
2 57801 1 111
2 57802 1 111
2 57803 1 111
2 57804 1 113
2 57805 1 113
2 57806 1 113
2 57807 1 113
2 57808 1 113
2 57809 1 114
2 57810 1 114
2 57811 1 114
2 57812 1 114
2 57813 1 114
2 57814 1 114
2 57815 1 114
2 57816 1 114
2 57817 1 114
2 57818 1 114
2 57819 1 114
2 57820 1 114
2 57821 1 114
2 57822 1 114
2 57823 1 114
2 57824 1 114
2 57825 1 114
2 57826 1 114
2 57827 1 114
2 57828 1 114
2 57829 1 114
2 57830 1 114
2 57831 1 114
2 57832 1 114
2 57833 1 114
2 57834 1 114
2 57835 1 114
2 57836 1 114
2 57837 1 114
2 57838 1 114
2 57839 1 115
2 57840 1 115
2 57841 1 115
2 57842 1 115
2 57843 1 115
2 57844 1 115
2 57845 1 115
2 57846 1 115
2 57847 1 116
2 57848 1 116
2 57849 1 116
2 57850 1 116
2 57851 1 116
2 57852 1 117
2 57853 1 117
2 57854 1 117
2 57855 1 126
2 57856 1 126
2 57857 1 126
2 57858 1 126
2 57859 1 126
2 57860 1 126
2 57861 1 126
2 57862 1 126
2 57863 1 126
2 57864 1 126
2 57865 1 126
2 57866 1 126
2 57867 1 126
2 57868 1 126
2 57869 1 126
2 57870 1 126
2 57871 1 126
2 57872 1 126
2 57873 1 126
2 57874 1 126
2 57875 1 126
2 57876 1 126
2 57877 1 126
2 57878 1 126
2 57879 1 126
2 57880 1 126
2 57881 1 126
2 57882 1 126
2 57883 1 126
2 57884 1 126
2 57885 1 126
2 57886 1 126
2 57887 1 126
2 57888 1 126
2 57889 1 126
2 57890 1 126
2 57891 1 126
2 57892 1 126
2 57893 1 126
2 57894 1 126
2 57895 1 126
2 57896 1 126
2 57897 1 126
2 57898 1 126
2 57899 1 126
2 57900 1 126
2 57901 1 126
2 57902 1 126
2 57903 1 126
2 57904 1 126
2 57905 1 126
2 57906 1 126
2 57907 1 126
2 57908 1 126
2 57909 1 126
2 57910 1 126
2 57911 1 126
2 57912 1 126
2 57913 1 126
2 57914 1 126
2 57915 1 126
2 57916 1 126
2 57917 1 126
2 57918 1 126
2 57919 1 126
2 57920 1 126
2 57921 1 126
2 57922 1 126
2 57923 1 126
2 57924 1 126
2 57925 1 126
2 57926 1 126
2 57927 1 126
2 57928 1 126
2 57929 1 126
2 57930 1 126
2 57931 1 126
2 57932 1 126
2 57933 1 126
2 57934 1 126
2 57935 1 126
2 57936 1 126
2 57937 1 126
2 57938 1 126
2 57939 1 126
2 57940 1 126
2 57941 1 126
2 57942 1 126
2 57943 1 126
2 57944 1 126
2 57945 1 126
2 57946 1 126
2 57947 1 126
2 57948 1 126
2 57949 1 126
2 57950 1 126
2 57951 1 126
2 57952 1 126
2 57953 1 126
2 57954 1 126
2 57955 1 126
2 57956 1 126
2 57957 1 126
2 57958 1 126
2 57959 1 126
2 57960 1 126
2 57961 1 126
2 57962 1 126
2 57963 1 126
2 57964 1 126
2 57965 1 126
2 57966 1 126
2 57967 1 126
2 57968 1 126
2 57969 1 127
2 57970 1 127
2 57971 1 127
2 57972 1 127
2 57973 1 127
2 57974 1 127
2 57975 1 127
2 57976 1 127
2 57977 1 127
2 57978 1 127
2 57979 1 127
2 57980 1 127
2 57981 1 127
2 57982 1 127
2 57983 1 127
2 57984 1 127
2 57985 1 127
2 57986 1 127
2 57987 1 127
2 57988 1 127
2 57989 1 127
2 57990 1 127
2 57991 1 127
2 57992 1 127
2 57993 1 127
2 57994 1 127
2 57995 1 127
2 57996 1 127
2 57997 1 127
2 57998 1 127
2 57999 1 127
2 58000 1 127
2 58001 1 127
2 58002 1 127
2 58003 1 127
2 58004 1 127
2 58005 1 127
2 58006 1 127
2 58007 1 127
2 58008 1 127
2 58009 1 127
2 58010 1 127
2 58011 1 127
2 58012 1 127
2 58013 1 127
2 58014 1 127
2 58015 1 127
2 58016 1 127
2 58017 1 127
2 58018 1 127
2 58019 1 127
2 58020 1 127
2 58021 1 127
2 58022 1 127
2 58023 1 127
2 58024 1 127
2 58025 1 127
2 58026 1 127
2 58027 1 127
2 58028 1 127
2 58029 1 127
2 58030 1 127
2 58031 1 127
2 58032 1 127
2 58033 1 127
2 58034 1 127
2 58035 1 127
2 58036 1 127
2 58037 1 127
2 58038 1 127
2 58039 1 127
2 58040 1 127
2 58041 1 127
2 58042 1 127
2 58043 1 127
2 58044 1 127
2 58045 1 127
2 58046 1 127
2 58047 1 127
2 58048 1 127
2 58049 1 127
2 58050 1 127
2 58051 1 127
2 58052 1 127
2 58053 1 127
2 58054 1 127
2 58055 1 127
2 58056 1 127
2 58057 1 127
2 58058 1 127
2 58059 1 127
2 58060 1 127
2 58061 1 127
2 58062 1 127
2 58063 1 127
2 58064 1 127
2 58065 1 127
2 58066 1 127
2 58067 1 128
2 58068 1 128
2 58069 1 128
2 58070 1 128
2 58071 1 128
2 58072 1 128
2 58073 1 128
2 58074 1 128
2 58075 1 128
2 58076 1 129
2 58077 1 129
2 58078 1 129
2 58079 1 129
2 58080 1 129
2 58081 1 129
2 58082 1 129
2 58083 1 129
2 58084 1 129
2 58085 1 129
2 58086 1 129
2 58087 1 129
2 58088 1 129
2 58089 1 129
2 58090 1 129
2 58091 1 129
2 58092 1 129
2 58093 1 129
2 58094 1 129
2 58095 1 129
2 58096 1 129
2 58097 1 129
2 58098 1 129
2 58099 1 129
2 58100 1 129
2 58101 1 129
2 58102 1 129
2 58103 1 129
2 58104 1 129
2 58105 1 129
2 58106 1 129
2 58107 1 129
2 58108 1 129
2 58109 1 129
2 58110 1 129
2 58111 1 129
2 58112 1 129
2 58113 1 129
2 58114 1 129
2 58115 1 129
2 58116 1 129
2 58117 1 129
2 58118 1 129
2 58119 1 129
2 58120 1 129
2 58121 1 129
2 58122 1 129
2 58123 1 129
2 58124 1 129
2 58125 1 129
2 58126 1 129
2 58127 1 129
2 58128 1 129
2 58129 1 130
2 58130 1 130
2 58131 1 130
2 58132 1 130
2 58133 1 130
2 58134 1 130
2 58135 1 130
2 58136 1 130
2 58137 1 130
2 58138 1 130
2 58139 1 130
2 58140 1 131
2 58141 1 131
2 58142 1 131
2 58143 1 132
2 58144 1 132
2 58145 1 132
2 58146 1 132
2 58147 1 132
2 58148 1 132
2 58149 1 132
2 58150 1 132
2 58151 1 132
2 58152 1 134
2 58153 1 134
2 58154 1 135
2 58155 1 135
2 58156 1 135
2 58157 1 135
2 58158 1 137
2 58159 1 137
2 58160 1 137
2 58161 1 137
2 58162 1 137
2 58163 1 138
2 58164 1 138
2 58165 1 138
2 58166 1 138
2 58167 1 138
2 58168 1 138
2 58169 1 138
2 58170 1 138
2 58171 1 138
2 58172 1 138
2 58173 1 138
2 58174 1 138
2 58175 1 138
2 58176 1 138
2 58177 1 138
2 58178 1 139
2 58179 1 139
2 58180 1 139
2 58181 1 139
2 58182 1 139
2 58183 1 139
2 58184 1 139
2 58185 1 140
2 58186 1 140
2 58187 1 140
2 58188 1 140
2 58189 1 140
2 58190 1 141
2 58191 1 141
2 58192 1 143
2 58193 1 143
2 58194 1 143
2 58195 1 146
2 58196 1 146
2 58197 1 146
2 58198 1 146
2 58199 1 146
2 58200 1 146
2 58201 1 146
2 58202 1 146
2 58203 1 146
2 58204 1 146
2 58205 1 146
2 58206 1 146
2 58207 1 146
2 58208 1 147
2 58209 1 147
2 58210 1 147
2 58211 1 147
2 58212 1 147
2 58213 1 147
2 58214 1 147
2 58215 1 147
2 58216 1 147
2 58217 1 147
2 58218 1 148
2 58219 1 148
2 58220 1 149
2 58221 1 149
2 58222 1 149
2 58223 1 150
2 58224 1 150
2 58225 1 150
2 58226 1 150
2 58227 1 150
2 58228 1 150
2 58229 1 150
2 58230 1 150
2 58231 1 150
2 58232 1 150
2 58233 1 151
2 58234 1 151
2 58235 1 151
2 58236 1 151
2 58237 1 151
2 58238 1 151
2 58239 1 151
2 58240 1 151
2 58241 1 151
2 58242 1 151
2 58243 1 151
2 58244 1 151
2 58245 1 151
2 58246 1 151
2 58247 1 151
2 58248 1 151
2 58249 1 151
2 58250 1 151
2 58251 1 151
2 58252 1 151
2 58253 1 151
2 58254 1 151
2 58255 1 151
2 58256 1 151
2 58257 1 151
2 58258 1 151
2 58259 1 151
2 58260 1 151
2 58261 1 151
2 58262 1 152
2 58263 1 152
2 58264 1 152
2 58265 1 152
2 58266 1 152
2 58267 1 152
2 58268 1 152
2 58269 1 152
2 58270 1 152
2 58271 1 152
2 58272 1 152
2 58273 1 152
2 58274 1 153
2 58275 1 153
2 58276 1 153
2 58277 1 153
2 58278 1 153
2 58279 1 153
2 58280 1 162
2 58281 1 162
2 58282 1 162
2 58283 1 162
2 58284 1 162
2 58285 1 162
2 58286 1 162
2 58287 1 162
2 58288 1 162
2 58289 1 162
2 58290 1 163
2 58291 1 163
2 58292 1 163
2 58293 1 163
2 58294 1 163
2 58295 1 163
2 58296 1 164
2 58297 1 164
2 58298 1 164
2 58299 1 165
2 58300 1 165
2 58301 1 165
2 58302 1 165
2 58303 1 165
2 58304 1 165
2 58305 1 165
2 58306 1 165
2 58307 1 165
2 58308 1 165
2 58309 1 165
2 58310 1 165
2 58311 1 165
2 58312 1 165
2 58313 1 165
2 58314 1 165
2 58315 1 165
2 58316 1 165
2 58317 1 166
2 58318 1 166
2 58319 1 166
2 58320 1 166
2 58321 1 166
2 58322 1 166
2 58323 1 166
2 58324 1 167
2 58325 1 167
2 58326 1 167
2 58327 1 167
2 58328 1 167
2 58329 1 167
2 58330 1 167
2 58331 1 168
2 58332 1 168
2 58333 1 168
2 58334 1 168
2 58335 1 169
2 58336 1 169
2 58337 1 170
2 58338 1 170
2 58339 1 170
2 58340 1 170
2 58341 1 170
2 58342 1 174
2 58343 1 174
2 58344 1 175
2 58345 1 175
2 58346 1 175
2 58347 1 175
2 58348 1 175
2 58349 1 175
2 58350 1 175
2 58351 1 182
2 58352 1 182
2 58353 1 182
2 58354 1 182
2 58355 1 182
2 58356 1 182
2 58357 1 182
2 58358 1 182
2 58359 1 182
2 58360 1 182
2 58361 1 182
2 58362 1 182
2 58363 1 182
2 58364 1 182
2 58365 1 182
2 58366 1 182
2 58367 1 182
2 58368 1 182
2 58369 1 182
2 58370 1 182
2 58371 1 182
2 58372 1 182
2 58373 1 182
2 58374 1 182
2 58375 1 182
2 58376 1 182
2 58377 1 182
2 58378 1 182
2 58379 1 182
2 58380 1 182
2 58381 1 182
2 58382 1 182
2 58383 1 182
2 58384 1 182
2 58385 1 182
2 58386 1 182
2 58387 1 182
2 58388 1 182
2 58389 1 182
2 58390 1 182
2 58391 1 182
2 58392 1 182
2 58393 1 182
2 58394 1 182
2 58395 1 182
2 58396 1 182
2 58397 1 182
2 58398 1 182
2 58399 1 182
2 58400 1 182
2 58401 1 182
2 58402 1 182
2 58403 1 182
2 58404 1 182
2 58405 1 182
2 58406 1 182
2 58407 1 182
2 58408 1 182
2 58409 1 182
2 58410 1 182
2 58411 1 182
2 58412 1 182
2 58413 1 182
2 58414 1 183
2 58415 1 183
2 58416 1 183
2 58417 1 183
2 58418 1 183
2 58419 1 183
2 58420 1 183
2 58421 1 183
2 58422 1 183
2 58423 1 183
2 58424 1 183
2 58425 1 183
2 58426 1 183
2 58427 1 183
2 58428 1 183
2 58429 1 183
2 58430 1 183
2 58431 1 183
2 58432 1 183
2 58433 1 183
2 58434 1 183
2 58435 1 183
2 58436 1 183
2 58437 1 183
2 58438 1 183
2 58439 1 183
2 58440 1 183
2 58441 1 183
2 58442 1 183
2 58443 1 183
2 58444 1 183
2 58445 1 183
2 58446 1 183
2 58447 1 183
2 58448 1 183
2 58449 1 183
2 58450 1 183
2 58451 1 183
2 58452 1 183
2 58453 1 183
2 58454 1 183
2 58455 1 183
2 58456 1 183
2 58457 1 183
2 58458 1 183
2 58459 1 183
2 58460 1 183
2 58461 1 183
2 58462 1 183
2 58463 1 183
2 58464 1 183
2 58465 1 183
2 58466 1 183
2 58467 1 183
2 58468 1 183
2 58469 1 183
2 58470 1 184
2 58471 1 184
2 58472 1 184
2 58473 1 184
2 58474 1 184
2 58475 1 184
2 58476 1 184
2 58477 1 184
2 58478 1 184
2 58479 1 184
2 58480 1 184
2 58481 1 184
2 58482 1 184
2 58483 1 184
2 58484 1 185
2 58485 1 185
2 58486 1 185
2 58487 1 185
2 58488 1 186
2 58489 1 186
2 58490 1 186
2 58491 1 186
2 58492 1 186
2 58493 1 186
2 58494 1 186
2 58495 1 188
2 58496 1 188
2 58497 1 189
2 58498 1 189
2 58499 1 190
2 58500 1 190
2 58501 1 194
2 58502 1 194
2 58503 1 195
2 58504 1 195
2 58505 1 195
2 58506 1 195
2 58507 1 195
2 58508 1 195
2 58509 1 195
2 58510 1 196
2 58511 1 196
2 58512 1 197
2 58513 1 197
2 58514 1 205
2 58515 1 205
2 58516 1 205
2 58517 1 205
2 58518 1 205
2 58519 1 205
2 58520 1 205
2 58521 1 205
2 58522 1 205
2 58523 1 206
2 58524 1 206
2 58525 1 206
2 58526 1 206
2 58527 1 206
2 58528 1 206
2 58529 1 206
2 58530 1 206
2 58531 1 206
2 58532 1 206
2 58533 1 206
2 58534 1 206
2 58535 1 206
2 58536 1 206
2 58537 1 206
2 58538 1 206
2 58539 1 206
2 58540 1 206
2 58541 1 206
2 58542 1 206
2 58543 1 206
2 58544 1 206
2 58545 1 206
2 58546 1 206
2 58547 1 206
2 58548 1 206
2 58549 1 206
2 58550 1 207
2 58551 1 207
2 58552 1 207
2 58553 1 207
2 58554 1 207
2 58555 1 207
2 58556 1 207
2 58557 1 207
2 58558 1 208
2 58559 1 208
2 58560 1 208
2 58561 1 208
2 58562 1 208
2 58563 1 208
2 58564 1 208
2 58565 1 208
2 58566 1 209
2 58567 1 209
2 58568 1 209
2 58569 1 209
2 58570 1 209
2 58571 1 209
2 58572 1 209
2 58573 1 209
2 58574 1 209
2 58575 1 210
2 58576 1 210
2 58577 1 210
2 58578 1 210
2 58579 1 210
2 58580 1 210
2 58581 1 210
2 58582 1 210
2 58583 1 210
2 58584 1 210
2 58585 1 210
2 58586 1 211
2 58587 1 211
2 58588 1 211
2 58589 1 211
2 58590 1 219
2 58591 1 219
2 58592 1 220
2 58593 1 220
2 58594 1 220
2 58595 1 220
2 58596 1 220
2 58597 1 220
2 58598 1 220
2 58599 1 220
2 58600 1 220
2 58601 1 220
2 58602 1 220
2 58603 1 220
2 58604 1 220
2 58605 1 220
2 58606 1 220
2 58607 1 220
2 58608 1 220
2 58609 1 220
2 58610 1 220
2 58611 1 220
2 58612 1 220
2 58613 1 220
2 58614 1 220
2 58615 1 220
2 58616 1 220
2 58617 1 220
2 58618 1 220
2 58619 1 220
2 58620 1 220
2 58621 1 220
2 58622 1 220
2 58623 1 220
2 58624 1 220
2 58625 1 220
2 58626 1 220
2 58627 1 220
2 58628 1 220
2 58629 1 220
2 58630 1 220
2 58631 1 220
2 58632 1 220
2 58633 1 224
2 58634 1 224
2 58635 1 227
2 58636 1 227
2 58637 1 227
2 58638 1 227
2 58639 1 227
2 58640 1 227
2 58641 1 227
2 58642 1 227
2 58643 1 227
2 58644 1 228
2 58645 1 228
2 58646 1 228
2 58647 1 228
2 58648 1 228
2 58649 1 231
2 58650 1 231
2 58651 1 231
2 58652 1 231
2 58653 1 231
2 58654 1 231
2 58655 1 231
2 58656 1 231
2 58657 1 231
2 58658 1 231
2 58659 1 231
2 58660 1 231
2 58661 1 231
2 58662 1 231
2 58663 1 231
2 58664 1 231
2 58665 1 231
2 58666 1 231
2 58667 1 231
2 58668 1 231
2 58669 1 231
2 58670 1 231
2 58671 1 231
2 58672 1 231
2 58673 1 231
2 58674 1 231
2 58675 1 231
2 58676 1 231
2 58677 1 231
2 58678 1 231
2 58679 1 231
2 58680 1 231
2 58681 1 231
2 58682 1 231
2 58683 1 231
2 58684 1 231
2 58685 1 231
2 58686 1 231
2 58687 1 231
2 58688 1 231
2 58689 1 231
2 58690 1 231
2 58691 1 231
2 58692 1 231
2 58693 1 231
2 58694 1 231
2 58695 1 231
2 58696 1 231
2 58697 1 231
2 58698 1 231
2 58699 1 231
2 58700 1 231
2 58701 1 231
2 58702 1 231
2 58703 1 232
2 58704 1 232
2 58705 1 232
2 58706 1 232
2 58707 1 232
2 58708 1 232
2 58709 1 232
2 58710 1 232
2 58711 1 232
2 58712 1 232
2 58713 1 232
2 58714 1 232
2 58715 1 232
2 58716 1 232
2 58717 1 232
2 58718 1 232
2 58719 1 232
2 58720 1 232
2 58721 1 232
2 58722 1 232
2 58723 1 232
2 58724 1 249
2 58725 1 249
2 58726 1 249
2 58727 1 249
2 58728 1 249
2 58729 1 249
2 58730 1 249
2 58731 1 249
2 58732 1 249
2 58733 1 249
2 58734 1 249
2 58735 1 250
2 58736 1 250
2 58737 1 250
2 58738 1 250
2 58739 1 250
2 58740 1 250
2 58741 1 250
2 58742 1 250
2 58743 1 250
2 58744 1 250
2 58745 1 250
2 58746 1 250
2 58747 1 250
2 58748 1 250
2 58749 1 250
2 58750 1 250
2 58751 1 250
2 58752 1 250
2 58753 1 250
2 58754 1 250
2 58755 1 250
2 58756 1 250
2 58757 1 250
2 58758 1 250
2 58759 1 250
2 58760 1 250
2 58761 1 250
2 58762 1 250
2 58763 1 250
2 58764 1 250
2 58765 1 250
2 58766 1 250
2 58767 1 250
2 58768 1 250
2 58769 1 250
2 58770 1 250
2 58771 1 250
2 58772 1 250
2 58773 1 250
2 58774 1 250
2 58775 1 250
2 58776 1 250
2 58777 1 250
2 58778 1 250
2 58779 1 250
2 58780 1 250
2 58781 1 250
2 58782 1 250
2 58783 1 250
2 58784 1 250
2 58785 1 250
2 58786 1 250
2 58787 1 250
2 58788 1 250
2 58789 1 250
2 58790 1 250
2 58791 1 250
2 58792 1 251
2 58793 1 251
2 58794 1 251
2 58795 1 251
2 58796 1 251
2 58797 1 253
2 58798 1 253
2 58799 1 253
2 58800 1 253
2 58801 1 253
2 58802 1 253
2 58803 1 253
2 58804 1 253
2 58805 1 253
2 58806 1 253
2 58807 1 253
2 58808 1 254
2 58809 1 254
2 58810 1 254
2 58811 1 254
2 58812 1 255
2 58813 1 255
2 58814 1 255
2 58815 1 255
2 58816 1 255
2 58817 1 255
2 58818 1 255
2 58819 1 255
2 58820 1 255
2 58821 1 255
2 58822 1 255
2 58823 1 255
2 58824 1 256
2 58825 1 256
2 58826 1 256
2 58827 1 257
2 58828 1 257
2 58829 1 257
2 58830 1 258
2 58831 1 258
2 58832 1 258
2 58833 1 258
2 58834 1 258
2 58835 1 258
2 58836 1 258
2 58837 1 258
2 58838 1 258
2 58839 1 258
2 58840 1 258
2 58841 1 258
2 58842 1 258
2 58843 1 258
2 58844 1 258
2 58845 1 258
2 58846 1 259
2 58847 1 259
2 58848 1 259
2 58849 1 259
2 58850 1 259
2 58851 1 259
2 58852 1 259
2 58853 1 259
2 58854 1 259
2 58855 1 259
2 58856 1 259
2 58857 1 259
2 58858 1 259
2 58859 1 259
2 58860 1 259
2 58861 1 259
2 58862 1 259
2 58863 1 259
2 58864 1 259
2 58865 1 259
2 58866 1 259
2 58867 1 259
2 58868 1 259
2 58869 1 259
2 58870 1 259
2 58871 1 259
2 58872 1 259
2 58873 1 259
2 58874 1 259
2 58875 1 259
2 58876 1 259
2 58877 1 259
2 58878 1 259
2 58879 1 259
2 58880 1 259
2 58881 1 259
2 58882 1 259
2 58883 1 259
2 58884 1 260
2 58885 1 260
2 58886 1 260
2 58887 1 260
2 58888 1 260
2 58889 1 260
2 58890 1 260
2 58891 1 260
2 58892 1 260
2 58893 1 260
2 58894 1 260
2 58895 1 260
2 58896 1 260
2 58897 1 260
2 58898 1 262
2 58899 1 262
2 58900 1 262
2 58901 1 262
2 58902 1 262
2 58903 1 262
2 58904 1 263
2 58905 1 263
2 58906 1 263
2 58907 1 271
2 58908 1 271
2 58909 1 271
2 58910 1 271
2 58911 1 272
2 58912 1 272
2 58913 1 273
2 58914 1 273
2 58915 1 273
2 58916 1 273
2 58917 1 273
2 58918 1 274
2 58919 1 274
2 58920 1 274
2 58921 1 275
2 58922 1 275
2 58923 1 275
2 58924 1 275
2 58925 1 275
2 58926 1 275
2 58927 1 275
2 58928 1 275
2 58929 1 275
2 58930 1 275
2 58931 1 276
2 58932 1 276
2 58933 1 276
2 58934 1 276
2 58935 1 276
2 58936 1 276
2 58937 1 276
2 58938 1 276
2 58939 1 276
2 58940 1 276
2 58941 1 276
2 58942 1 276
2 58943 1 276
2 58944 1 276
2 58945 1 276
2 58946 1 276
2 58947 1 276
2 58948 1 276
2 58949 1 276
2 58950 1 276
2 58951 1 278
2 58952 1 278
2 58953 1 279
2 58954 1 279
2 58955 1 279
2 58956 1 279
2 58957 1 279
2 58958 1 280
2 58959 1 280
2 58960 1 280
2 58961 1 280
2 58962 1 280
2 58963 1 280
2 58964 1 280
2 58965 1 280
2 58966 1 280
2 58967 1 280
2 58968 1 280
2 58969 1 280
2 58970 1 280
2 58971 1 280
2 58972 1 280
2 58973 1 280
2 58974 1 280
2 58975 1 280
2 58976 1 280
2 58977 1 280
2 58978 1 280
2 58979 1 280
2 58980 1 280
2 58981 1 280
2 58982 1 280
2 58983 1 280
2 58984 1 280
2 58985 1 280
2 58986 1 280
2 58987 1 280
2 58988 1 280
2 58989 1 280
2 58990 1 280
2 58991 1 280
2 58992 1 280
2 58993 1 280
2 58994 1 280
2 58995 1 282
2 58996 1 282
2 58997 1 289
2 58998 1 289
2 58999 1 289
2 59000 1 289
2 59001 1 289
2 59002 1 289
2 59003 1 289
2 59004 1 289
2 59005 1 289
2 59006 1 289
2 59007 1 289
2 59008 1 289
2 59009 1 290
2 59010 1 290
2 59011 1 290
2 59012 1 290
2 59013 1 290
2 59014 1 290
2 59015 1 290
2 59016 1 291
2 59017 1 291
2 59018 1 291
2 59019 1 291
2 59020 1 291
2 59021 1 291
2 59022 1 291
2 59023 1 291
2 59024 1 291
2 59025 1 291
2 59026 1 291
2 59027 1 292
2 59028 1 292
2 59029 1 292
2 59030 1 292
2 59031 1 293
2 59032 1 293
2 59033 1 293
2 59034 1 293
2 59035 1 293
2 59036 1 293
2 59037 1 293
2 59038 1 293
2 59039 1 293
2 59040 1 294
2 59041 1 294
2 59042 1 294
2 59043 1 294
2 59044 1 294
2 59045 1 294
2 59046 1 295
2 59047 1 295
2 59048 1 295
2 59049 1 295
2 59050 1 296
2 59051 1 296
2 59052 1 296
2 59053 1 296
2 59054 1 296
2 59055 1 296
2 59056 1 297
2 59057 1 297
2 59058 1 298
2 59059 1 298
2 59060 1 298
2 59061 1 298
2 59062 1 298
2 59063 1 298
2 59064 1 298
2 59065 1 298
2 59066 1 298
2 59067 1 298
2 59068 1 303
2 59069 1 303
2 59070 1 303
2 59071 1 304
2 59072 1 304
2 59073 1 304
2 59074 1 304
2 59075 1 305
2 59076 1 305
2 59077 1 305
2 59078 1 305
2 59079 1 305
2 59080 1 305
2 59081 1 305
2 59082 1 305
2 59083 1 306
2 59084 1 306
2 59085 1 306
2 59086 1 306
2 59087 1 306
2 59088 1 306
2 59089 1 307
2 59090 1 307
2 59091 1 307
2 59092 1 308
2 59093 1 308
2 59094 1 308
2 59095 1 309
2 59096 1 309
2 59097 1 309
2 59098 1 309
2 59099 1 309
2 59100 1 309
2 59101 1 309
2 59102 1 309
2 59103 1 309
2 59104 1 309
2 59105 1 309
2 59106 1 309
2 59107 1 309
2 59108 1 309
2 59109 1 309
2 59110 1 309
2 59111 1 309
2 59112 1 309
2 59113 1 309
2 59114 1 313
2 59115 1 313
2 59116 1 313
2 59117 1 313
2 59118 1 313
2 59119 1 314
2 59120 1 314
2 59121 1 314
2 59122 1 314
2 59123 1 314
2 59124 1 314
2 59125 1 314
2 59126 1 314
2 59127 1 314
2 59128 1 314
2 59129 1 314
2 59130 1 314
2 59131 1 314
2 59132 1 314
2 59133 1 314
2 59134 1 314
2 59135 1 314
2 59136 1 314
2 59137 1 314
2 59138 1 314
2 59139 1 314
2 59140 1 314
2 59141 1 314
2 59142 1 314
2 59143 1 314
2 59144 1 314
2 59145 1 314
2 59146 1 314
2 59147 1 314
2 59148 1 314
2 59149 1 314
2 59150 1 314
2 59151 1 314
2 59152 1 314
2 59153 1 314
2 59154 1 314
2 59155 1 314
2 59156 1 314
2 59157 1 314
2 59158 1 314
2 59159 1 314
2 59160 1 315
2 59161 1 315
2 59162 1 315
2 59163 1 315
2 59164 1 315
2 59165 1 315
2 59166 1 315
2 59167 1 315
2 59168 1 316
2 59169 1 316
2 59170 1 316
2 59171 1 324
2 59172 1 324
2 59173 1 324
2 59174 1 324
2 59175 1 324
2 59176 1 324
2 59177 1 325
2 59178 1 325
2 59179 1 325
2 59180 1 325
2 59181 1 325
2 59182 1 325
2 59183 1 325
2 59184 1 325
2 59185 1 325
2 59186 1 325
2 59187 1 325
2 59188 1 325
2 59189 1 325
2 59190 1 325
2 59191 1 326
2 59192 1 326
2 59193 1 326
2 59194 1 326
2 59195 1 326
2 59196 1 326
2 59197 1 326
2 59198 1 326
2 59199 1 326
2 59200 1 327
2 59201 1 327
2 59202 1 327
2 59203 1 327
2 59204 1 327
2 59205 1 327
2 59206 1 327
2 59207 1 327
2 59208 1 327
2 59209 1 327
2 59210 1 327
2 59211 1 327
2 59212 1 327
2 59213 1 327
2 59214 1 327
2 59215 1 327
2 59216 1 327
2 59217 1 327
2 59218 1 327
2 59219 1 327
2 59220 1 327
2 59221 1 327
2 59222 1 327
2 59223 1 327
2 59224 1 327
2 59225 1 327
2 59226 1 327
2 59227 1 327
2 59228 1 327
2 59229 1 327
2 59230 1 327
2 59231 1 327
2 59232 1 327
2 59233 1 327
2 59234 1 327
2 59235 1 327
2 59236 1 327
2 59237 1 327
2 59238 1 327
2 59239 1 331
2 59240 1 331
2 59241 1 331
2 59242 1 332
2 59243 1 332
2 59244 1 335
2 59245 1 335
2 59246 1 338
2 59247 1 338
2 59248 1 338
2 59249 1 338
2 59250 1 338
2 59251 1 338
2 59252 1 338
2 59253 1 338
2 59254 1 338
2 59255 1 338
2 59256 1 338
2 59257 1 338
2 59258 1 338
2 59259 1 338
2 59260 1 338
2 59261 1 338
2 59262 1 338
2 59263 1 338
2 59264 1 338
2 59265 1 338
2 59266 1 338
2 59267 1 338
2 59268 1 338
2 59269 1 338
2 59270 1 338
2 59271 1 338
2 59272 1 338
2 59273 1 338
2 59274 1 339
2 59275 1 339
2 59276 1 340
2 59277 1 340
2 59278 1 341
2 59279 1 341
2 59280 1 341
2 59281 1 342
2 59282 1 342
2 59283 1 342
2 59284 1 352
2 59285 1 352
2 59286 1 352
2 59287 1 352
2 59288 1 352
2 59289 1 352
2 59290 1 353
2 59291 1 353
2 59292 1 353
2 59293 1 353
2 59294 1 353
2 59295 1 353
2 59296 1 354
2 59297 1 354
2 59298 1 354
2 59299 1 354
2 59300 1 354
2 59301 1 354
2 59302 1 354
2 59303 1 354
2 59304 1 355
2 59305 1 355
2 59306 1 355
2 59307 1 355
2 59308 1 355
2 59309 1 355
2 59310 1 356
2 59311 1 356
2 59312 1 356
2 59313 1 356
2 59314 1 356
2 59315 1 356
2 59316 1 356
2 59317 1 356
2 59318 1 357
2 59319 1 357
2 59320 1 357
2 59321 1 357
2 59322 1 357
2 59323 1 357
2 59324 1 357
2 59325 1 357
2 59326 1 357
2 59327 1 366
2 59328 1 366
2 59329 1 366
2 59330 1 366
2 59331 1 367
2 59332 1 367
2 59333 1 367
2 59334 1 368
2 59335 1 368
2 59336 1 368
2 59337 1 368
2 59338 1 368
2 59339 1 368
2 59340 1 369
2 59341 1 369
2 59342 1 369
2 59343 1 375
2 59344 1 375
2 59345 1 378
2 59346 1 378
2 59347 1 379
2 59348 1 379
2 59349 1 379
2 59350 1 379
2 59351 1 379
2 59352 1 379
2 59353 1 379
2 59354 1 379
2 59355 1 379
2 59356 1 379
2 59357 1 379
2 59358 1 379
2 59359 1 379
2 59360 1 379
2 59361 1 380
2 59362 1 380
2 59363 1 381
2 59364 1 381
2 59365 1 381
2 59366 1 381
2 59367 1 381
2 59368 1 381
2 59369 1 381
2 59370 1 381
2 59371 1 381
2 59372 1 381
2 59373 1 381
2 59374 1 381
2 59375 1 381
2 59376 1 381
2 59377 1 381
2 59378 1 381
2 59379 1 382
2 59380 1 382
2 59381 1 382
2 59382 1 383
2 59383 1 383
2 59384 1 391
2 59385 1 391
2 59386 1 392
2 59387 1 392
2 59388 1 392
2 59389 1 392
2 59390 1 397
2 59391 1 397
2 59392 1 397
2 59393 1 397
2 59394 1 398
2 59395 1 398
2 59396 1 399
2 59397 1 399
2 59398 1 399
2 59399 1 399
2 59400 1 408
2 59401 1 408
2 59402 1 408
2 59403 1 408
2 59404 1 408
2 59405 1 409
2 59406 1 409
2 59407 1 409
2 59408 1 409
2 59409 1 409
2 59410 1 409
2 59411 1 409
2 59412 1 409
2 59413 1 409
2 59414 1 410
2 59415 1 410
2 59416 1 412
2 59417 1 412
2 59418 1 413
2 59419 1 413
2 59420 1 413
2 59421 1 413
2 59422 1 414
2 59423 1 414
2 59424 1 414
2 59425 1 414
2 59426 1 414
2 59427 1 414
2 59428 1 414
2 59429 1 414
2 59430 1 414
2 59431 1 414
2 59432 1 414
2 59433 1 414
2 59434 1 414
2 59435 1 414
2 59436 1 414
2 59437 1 414
2 59438 1 415
2 59439 1 415
2 59440 1 415
2 59441 1 416
2 59442 1 416
2 59443 1 416
2 59444 1 416
2 59445 1 416
2 59446 1 416
2 59447 1 417
2 59448 1 417
2 59449 1 417
2 59450 1 417
2 59451 1 418
2 59452 1 418
2 59453 1 418
2 59454 1 418
2 59455 1 418
2 59456 1 418
2 59457 1 418
2 59458 1 419
2 59459 1 419
2 59460 1 419
2 59461 1 419
2 59462 1 419
2 59463 1 419
2 59464 1 419
2 59465 1 420
2 59466 1 420
2 59467 1 423
2 59468 1 423
2 59469 1 426
2 59470 1 426
2 59471 1 426
2 59472 1 426
2 59473 1 426
2 59474 1 426
2 59475 1 426
2 59476 1 426
2 59477 1 426
2 59478 1 426
2 59479 1 426
2 59480 1 426
2 59481 1 426
2 59482 1 427
2 59483 1 427
2 59484 1 427
2 59485 1 427
2 59486 1 427
2 59487 1 427
2 59488 1 432
2 59489 1 432
2 59490 1 432
2 59491 1 432
2 59492 1 452
2 59493 1 452
2 59494 1 452
2 59495 1 452
2 59496 1 452
2 59497 1 452
2 59498 1 452
2 59499 1 452
2 59500 1 452
2 59501 1 452
2 59502 1 452
2 59503 1 452
2 59504 1 452
2 59505 1 452
2 59506 1 453
2 59507 1 453
2 59508 1 453
2 59509 1 453
2 59510 1 454
2 59511 1 454
2 59512 1 454
2 59513 1 454
2 59514 1 455
2 59515 1 455
2 59516 1 455
2 59517 1 455
2 59518 1 457
2 59519 1 457
2 59520 1 457
2 59521 1 457
2 59522 1 457
2 59523 1 460
2 59524 1 460
2 59525 1 460
2 59526 1 460
2 59527 1 460
2 59528 1 460
2 59529 1 460
2 59530 1 460
2 59531 1 463
2 59532 1 463
2 59533 1 463
2 59534 1 464
2 59535 1 464
2 59536 1 470
2 59537 1 470
2 59538 1 484
2 59539 1 484
2 59540 1 484
2 59541 1 484
2 59542 1 484
2 59543 1 484
2 59544 1 484
2 59545 1 484
2 59546 1 484
2 59547 1 484
2 59548 1 484
2 59549 1 484
2 59550 1 484
2 59551 1 484
2 59552 1 484
2 59553 1 484
2 59554 1 485
2 59555 1 485
2 59556 1 485
2 59557 1 485
2 59558 1 485
2 59559 1 485
2 59560 1 485
2 59561 1 485
2 59562 1 487
2 59563 1 487
2 59564 1 487
2 59565 1 487
2 59566 1 487
2 59567 1 487
2 59568 1 487
2 59569 1 487
2 59570 1 487
2 59571 1 487
2 59572 1 487
2 59573 1 488
2 59574 1 488
2 59575 1 488
2 59576 1 488
2 59577 1 488
2 59578 1 502
2 59579 1 502
2 59580 1 502
2 59581 1 502
2 59582 1 502
2 59583 1 502
2 59584 1 502
2 59585 1 505
2 59586 1 505
2 59587 1 505
2 59588 1 505
2 59589 1 505
2 59590 1 505
2 59591 1 505
2 59592 1 505
2 59593 1 506
2 59594 1 506
2 59595 1 521
2 59596 1 521
2 59597 1 521
2 59598 1 522
2 59599 1 522
2 59600 1 522
2 59601 1 522
2 59602 1 522
2 59603 1 529
2 59604 1 529
2 59605 1 529
2 59606 1 529
2 59607 1 529
2 59608 1 529
2 59609 1 529
2 59610 1 529
2 59611 1 529
2 59612 1 529
2 59613 1 529
2 59614 1 529
2 59615 1 529
2 59616 1 529
2 59617 1 529
2 59618 1 529
2 59619 1 529
2 59620 1 529
2 59621 1 529
2 59622 1 529
2 59623 1 529
2 59624 1 529
2 59625 1 529
2 59626 1 529
2 59627 1 530
2 59628 1 530
2 59629 1 530
2 59630 1 530
2 59631 1 530
2 59632 1 530
2 59633 1 530
2 59634 1 530
2 59635 1 530
2 59636 1 530
2 59637 1 530
2 59638 1 530
2 59639 1 530
2 59640 1 530
2 59641 1 530
2 59642 1 530
2 59643 1 530
2 59644 1 530
2 59645 1 531
2 59646 1 531
2 59647 1 531
2 59648 1 531
2 59649 1 531
2 59650 1 531
2 59651 1 531
2 59652 1 531
2 59653 1 531
2 59654 1 531
2 59655 1 531
2 59656 1 531
2 59657 1 531
2 59658 1 531
2 59659 1 531
2 59660 1 531
2 59661 1 531
2 59662 1 531
2 59663 1 531
2 59664 1 531
2 59665 1 531
2 59666 1 531
2 59667 1 532
2 59668 1 532
2 59669 1 532
2 59670 1 532
2 59671 1 532
2 59672 1 532
2 59673 1 532
2 59674 1 532
2 59675 1 532
2 59676 1 532
2 59677 1 532
2 59678 1 532
2 59679 1 532
2 59680 1 532
2 59681 1 532
2 59682 1 532
2 59683 1 532
2 59684 1 532
2 59685 1 532
2 59686 1 532
2 59687 1 532
2 59688 1 532
2 59689 1 532
2 59690 1 534
2 59691 1 534
2 59692 1 534
2 59693 1 534
2 59694 1 534
2 59695 1 535
2 59696 1 535
2 59697 1 535
2 59698 1 535
2 59699 1 535
2 59700 1 536
2 59701 1 536
2 59702 1 536
2 59703 1 536
2 59704 1 536
2 59705 1 536
2 59706 1 537
2 59707 1 537
2 59708 1 537
2 59709 1 537
2 59710 1 537
2 59711 1 537
2 59712 1 537
2 59713 1 537
2 59714 1 538
2 59715 1 538
2 59716 1 539
2 59717 1 539
2 59718 1 539
2 59719 1 539
2 59720 1 539
2 59721 1 539
2 59722 1 539
2 59723 1 539
2 59724 1 539
2 59725 1 539
2 59726 1 540
2 59727 1 540
2 59728 1 540
2 59729 1 540
2 59730 1 540
2 59731 1 540
2 59732 1 540
2 59733 1 540
2 59734 1 557
2 59735 1 557
2 59736 1 557
2 59737 1 557
2 59738 1 557
2 59739 1 557
2 59740 1 557
2 59741 1 557
2 59742 1 557
2 59743 1 557
2 59744 1 557
2 59745 1 557
2 59746 1 557
2 59747 1 558
2 59748 1 558
2 59749 1 558
2 59750 1 558
2 59751 1 558
2 59752 1 558
2 59753 1 558
2 59754 1 558
2 59755 1 558
2 59756 1 559
2 59757 1 559
2 59758 1 559
2 59759 1 559
2 59760 1 559
2 59761 1 559
2 59762 1 559
2 59763 1 560
2 59764 1 560
2 59765 1 560
2 59766 1 560
2 59767 1 560
2 59768 1 560
2 59769 1 560
2 59770 1 560
2 59771 1 560
2 59772 1 561
2 59773 1 561
2 59774 1 561
2 59775 1 561
2 59776 1 561
2 59777 1 561
2 59778 1 561
2 59779 1 561
2 59780 1 561
2 59781 1 561
2 59782 1 561
2 59783 1 562
2 59784 1 562
2 59785 1 562
2 59786 1 562
2 59787 1 564
2 59788 1 564
2 59789 1 564
2 59790 1 564
2 59791 1 565
2 59792 1 565
2 59793 1 565
2 59794 1 565
2 59795 1 565
2 59796 1 567
2 59797 1 567
2 59798 1 567
2 59799 1 567
2 59800 1 567
2 59801 1 567
2 59802 1 568
2 59803 1 568
2 59804 1 568
2 59805 1 568
2 59806 1 568
2 59807 1 568
2 59808 1 568
2 59809 1 568
2 59810 1 568
2 59811 1 569
2 59812 1 569
2 59813 1 570
2 59814 1 570
2 59815 1 570
2 59816 1 570
2 59817 1 570
2 59818 1 570
2 59819 1 570
2 59820 1 571
2 59821 1 571
2 59822 1 572
2 59823 1 572
2 59824 1 572
2 59825 1 573
2 59826 1 573
2 59827 1 573
2 59828 1 573
2 59829 1 573
2 59830 1 573
2 59831 1 578
2 59832 1 578
2 59833 1 586
2 59834 1 586
2 59835 1 586
2 59836 1 586
2 59837 1 586
2 59838 1 587
2 59839 1 587
2 59840 1 587
2 59841 1 587
2 59842 1 587
2 59843 1 587
2 59844 1 587
2 59845 1 587
2 59846 1 587
2 59847 1 587
2 59848 1 587
2 59849 1 587
2 59850 1 587
2 59851 1 587
2 59852 1 587
2 59853 1 587
2 59854 1 587
2 59855 1 587
2 59856 1 587
2 59857 1 587
2 59858 1 587
2 59859 1 587
2 59860 1 587
2 59861 1 587
2 59862 1 587
2 59863 1 587
2 59864 1 587
2 59865 1 587
2 59866 1 587
2 59867 1 587
2 59868 1 587
2 59869 1 587
2 59870 1 587
2 59871 1 588
2 59872 1 588
2 59873 1 588
2 59874 1 588
2 59875 1 588
2 59876 1 588
2 59877 1 588
2 59878 1 588
2 59879 1 588
2 59880 1 588
2 59881 1 588
2 59882 1 588
2 59883 1 588
2 59884 1 588
2 59885 1 588
2 59886 1 588
2 59887 1 588
2 59888 1 588
2 59889 1 588
2 59890 1 588
2 59891 1 589
2 59892 1 589
2 59893 1 589
2 59894 1 589
2 59895 1 590
2 59896 1 590
2 59897 1 590
2 59898 1 590
2 59899 1 590
2 59900 1 590
2 59901 1 590
2 59902 1 590
2 59903 1 590
2 59904 1 590
2 59905 1 590
2 59906 1 591
2 59907 1 591
2 59908 1 591
2 59909 1 591
2 59910 1 602
2 59911 1 602
2 59912 1 602
2 59913 1 602
2 59914 1 602
2 59915 1 602
2 59916 1 602
2 59917 1 602
2 59918 1 602
2 59919 1 602
2 59920 1 602
2 59921 1 602
2 59922 1 602
2 59923 1 602
2 59924 1 602
2 59925 1 602
2 59926 1 604
2 59927 1 604
2 59928 1 604
2 59929 1 604
2 59930 1 604
2 59931 1 604
2 59932 1 604
2 59933 1 604
2 59934 1 604
2 59935 1 604
2 59936 1 604
2 59937 1 604
2 59938 1 604
2 59939 1 604
2 59940 1 604
2 59941 1 604
2 59942 1 604
2 59943 1 604
2 59944 1 604
2 59945 1 604
2 59946 1 604
2 59947 1 604
2 59948 1 604
2 59949 1 604
2 59950 1 604
2 59951 1 604
2 59952 1 604
2 59953 1 604
2 59954 1 604
2 59955 1 605
2 59956 1 605
2 59957 1 605
2 59958 1 605
2 59959 1 605
2 59960 1 605
2 59961 1 605
2 59962 1 605
2 59963 1 605
2 59964 1 605
2 59965 1 605
2 59966 1 605
2 59967 1 605
2 59968 1 605
2 59969 1 605
2 59970 1 605
2 59971 1 605
2 59972 1 605
2 59973 1 605
2 59974 1 605
2 59975 1 605
2 59976 1 605
2 59977 1 605
2 59978 1 605
2 59979 1 605
2 59980 1 605
2 59981 1 605
2 59982 1 605
2 59983 1 605
2 59984 1 605
2 59985 1 605
2 59986 1 605
2 59987 1 605
2 59988 1 605
2 59989 1 605
2 59990 1 605
2 59991 1 605
2 59992 1 605
2 59993 1 605
2 59994 1 605
2 59995 1 605
2 59996 1 605
2 59997 1 605
2 59998 1 605
2 59999 1 605
2 60000 1 605
2 60001 1 605
2 60002 1 605
2 60003 1 605
2 60004 1 606
2 60005 1 606
2 60006 1 606
2 60007 1 606
2 60008 1 607
2 60009 1 607
2 60010 1 607
2 60011 1 607
2 60012 1 607
2 60013 1 607
2 60014 1 607
2 60015 1 607
2 60016 1 607
2 60017 1 607
2 60018 1 607
2 60019 1 607
2 60020 1 607
2 60021 1 607
2 60022 1 607
2 60023 1 608
2 60024 1 608
2 60025 1 608
2 60026 1 608
2 60027 1 609
2 60028 1 609
2 60029 1 609
2 60030 1 609
2 60031 1 609
2 60032 1 609
2 60033 1 610
2 60034 1 610
2 60035 1 610
2 60036 1 610
2 60037 1 610
2 60038 1 617
2 60039 1 617
2 60040 1 618
2 60041 1 618
2 60042 1 619
2 60043 1 619
2 60044 1 619
2 60045 1 619
2 60046 1 619
2 60047 1 619
2 60048 1 619
2 60049 1 619
2 60050 1 619
2 60051 1 624
2 60052 1 624
2 60053 1 624
2 60054 1 624
2 60055 1 624
2 60056 1 624
2 60057 1 624
2 60058 1 624
2 60059 1 624
2 60060 1 624
2 60061 1 624
2 60062 1 625
2 60063 1 625
2 60064 1 625
2 60065 1 626
2 60066 1 626
2 60067 1 626
2 60068 1 629
2 60069 1 629
2 60070 1 629
2 60071 1 633
2 60072 1 633
2 60073 1 633
2 60074 1 633
2 60075 1 633
2 60076 1 633
2 60077 1 633
2 60078 1 633
2 60079 1 633
2 60080 1 633
2 60081 1 633
2 60082 1 633
2 60083 1 634
2 60084 1 634
2 60085 1 634
2 60086 1 634
2 60087 1 634
2 60088 1 634
2 60089 1 635
2 60090 1 635
2 60091 1 635
2 60092 1 637
2 60093 1 637
2 60094 1 641
2 60095 1 641
2 60096 1 641
2 60097 1 641
2 60098 1 641
2 60099 1 641
2 60100 1 641
2 60101 1 642
2 60102 1 642
2 60103 1 643
2 60104 1 643
2 60105 1 643
2 60106 1 643
2 60107 1 644
2 60108 1 644
2 60109 1 645
2 60110 1 645
2 60111 1 646
2 60112 1 646
2 60113 1 646
2 60114 1 646
2 60115 1 646
2 60116 1 646
2 60117 1 646
2 60118 1 646
2 60119 1 646
2 60120 1 646
2 60121 1 646
2 60122 1 646
2 60123 1 646
2 60124 1 646
2 60125 1 646
2 60126 1 646
2 60127 1 646
2 60128 1 647
2 60129 1 647
2 60130 1 647
2 60131 1 647
2 60132 1 647
2 60133 1 647
2 60134 1 647
2 60135 1 647
2 60136 1 647
2 60137 1 648
2 60138 1 648
2 60139 1 649
2 60140 1 649
2 60141 1 649
2 60142 1 649
2 60143 1 649
2 60144 1 649
2 60145 1 649
2 60146 1 649
2 60147 1 649
2 60148 1 649
2 60149 1 649
2 60150 1 649
2 60151 1 649
2 60152 1 649
2 60153 1 649
2 60154 1 649
2 60155 1 649
2 60156 1 649
2 60157 1 649
2 60158 1 649
2 60159 1 650
2 60160 1 650
2 60161 1 650
2 60162 1 666
2 60163 1 666
2 60164 1 666
2 60165 1 666
2 60166 1 666
2 60167 1 666
2 60168 1 666
2 60169 1 668
2 60170 1 668
2 60171 1 668
2 60172 1 671
2 60173 1 671
2 60174 1 672
2 60175 1 672
2 60176 1 673
2 60177 1 673
2 60178 1 673
2 60179 1 674
2 60180 1 674
2 60181 1 674
2 60182 1 674
2 60183 1 674
2 60184 1 674
2 60185 1 674
2 60186 1 674
2 60187 1 674
2 60188 1 674
2 60189 1 674
2 60190 1 674
2 60191 1 674
2 60192 1 674
2 60193 1 674
2 60194 1 674
2 60195 1 674
2 60196 1 674
2 60197 1 674
2 60198 1 674
2 60199 1 674
2 60200 1 674
2 60201 1 674
2 60202 1 674
2 60203 1 674
2 60204 1 674
2 60205 1 674
2 60206 1 674
2 60207 1 674
2 60208 1 674
2 60209 1 674
2 60210 1 674
2 60211 1 674
2 60212 1 674
2 60213 1 674
2 60214 1 674
2 60215 1 674
2 60216 1 674
2 60217 1 674
2 60218 1 674
2 60219 1 674
2 60220 1 674
2 60221 1 674
2 60222 1 674
2 60223 1 674
2 60224 1 674
2 60225 1 674
2 60226 1 674
2 60227 1 674
2 60228 1 674
2 60229 1 675
2 60230 1 675
2 60231 1 675
2 60232 1 675
2 60233 1 675
2 60234 1 675
2 60235 1 675
2 60236 1 675
2 60237 1 675
2 60238 1 675
2 60239 1 675
2 60240 1 675
2 60241 1 675
2 60242 1 675
2 60243 1 675
2 60244 1 675
2 60245 1 675
2 60246 1 675
2 60247 1 675
2 60248 1 675
2 60249 1 675
2 60250 1 675
2 60251 1 675
2 60252 1 675
2 60253 1 675
2 60254 1 675
2 60255 1 675
2 60256 1 675
2 60257 1 675
2 60258 1 676
2 60259 1 676
2 60260 1 676
2 60261 1 676
2 60262 1 676
2 60263 1 676
2 60264 1 676
2 60265 1 676
2 60266 1 676
2 60267 1 676
2 60268 1 676
2 60269 1 676
2 60270 1 676
2 60271 1 676
2 60272 1 676
2 60273 1 676
2 60274 1 676
2 60275 1 677
2 60276 1 677
2 60277 1 677
2 60278 1 677
2 60279 1 677
2 60280 1 677
2 60281 1 677
2 60282 1 677
2 60283 1 677
2 60284 1 677
2 60285 1 677
2 60286 1 677
2 60287 1 677
2 60288 1 677
2 60289 1 677
2 60290 1 677
2 60291 1 677
2 60292 1 677
2 60293 1 677
2 60294 1 677
2 60295 1 677
2 60296 1 677
2 60297 1 677
2 60298 1 677
2 60299 1 677
2 60300 1 677
2 60301 1 677
2 60302 1 677
2 60303 1 677
2 60304 1 677
2 60305 1 677
2 60306 1 677
2 60307 1 677
2 60308 1 677
2 60309 1 677
2 60310 1 677
2 60311 1 677
2 60312 1 677
2 60313 1 677
2 60314 1 677
2 60315 1 677
2 60316 1 677
2 60317 1 677
2 60318 1 678
2 60319 1 678
2 60320 1 678
2 60321 1 678
2 60322 1 678
2 60323 1 678
2 60324 1 678
2 60325 1 678
2 60326 1 678
2 60327 1 678
2 60328 1 678
2 60329 1 679
2 60330 1 679
2 60331 1 679
2 60332 1 679
2 60333 1 679
2 60334 1 679
2 60335 1 679
2 60336 1 679
2 60337 1 679
2 60338 1 679
2 60339 1 679
2 60340 1 679
2 60341 1 679
2 60342 1 679
2 60343 1 679
2 60344 1 679
2 60345 1 680
2 60346 1 680
2 60347 1 680
2 60348 1 680
2 60349 1 680
2 60350 1 680
2 60351 1 680
2 60352 1 680
2 60353 1 681
2 60354 1 681
2 60355 1 681
2 60356 1 681
2 60357 1 681
2 60358 1 681
2 60359 1 681
2 60360 1 681
2 60361 1 681
2 60362 1 683
2 60363 1 683
2 60364 1 683
2 60365 1 684
2 60366 1 684
2 60367 1 686
2 60368 1 686
2 60369 1 688
2 60370 1 688
2 60371 1 688
2 60372 1 688
2 60373 1 688
2 60374 1 688
2 60375 1 688
2 60376 1 688
2 60377 1 688
2 60378 1 688
2 60379 1 688
2 60380 1 688
2 60381 1 688
2 60382 1 688
2 60383 1 688
2 60384 1 688
2 60385 1 688
2 60386 1 688
2 60387 1 688
2 60388 1 688
2 60389 1 688
2 60390 1 688
2 60391 1 688
2 60392 1 688
2 60393 1 688
2 60394 1 688
2 60395 1 688
2 60396 1 688
2 60397 1 688
2 60398 1 688
2 60399 1 688
2 60400 1 688
2 60401 1 688
2 60402 1 688
2 60403 1 688
2 60404 1 688
2 60405 1 689
2 60406 1 689
2 60407 1 689
2 60408 1 689
2 60409 1 689
2 60410 1 689
2 60411 1 689
2 60412 1 689
2 60413 1 689
2 60414 1 689
2 60415 1 689
2 60416 1 689
2 60417 1 689
2 60418 1 689
2 60419 1 689
2 60420 1 689
2 60421 1 689
2 60422 1 689
2 60423 1 689
2 60424 1 689
2 60425 1 689
2 60426 1 689
2 60427 1 689
2 60428 1 689
2 60429 1 689
2 60430 1 689
2 60431 1 689
2 60432 1 689
2 60433 1 690
2 60434 1 690
2 60435 1 691
2 60436 1 691
2 60437 1 691
2 60438 1 693
2 60439 1 693
2 60440 1 693
2 60441 1 693
2 60442 1 693
2 60443 1 693
2 60444 1 698
2 60445 1 698
2 60446 1 698
2 60447 1 698
2 60448 1 698
2 60449 1 698
2 60450 1 699
2 60451 1 699
2 60452 1 699
2 60453 1 699
2 60454 1 699
2 60455 1 703
2 60456 1 703
2 60457 1 703
2 60458 1 703
2 60459 1 703
2 60460 1 703
2 60461 1 703
2 60462 1 703
2 60463 1 704
2 60464 1 704
2 60465 1 704
2 60466 1 711
2 60467 1 711
2 60468 1 711
2 60469 1 711
2 60470 1 711
2 60471 1 711
2 60472 1 711
2 60473 1 711
2 60474 1 711
2 60475 1 711
2 60476 1 711
2 60477 1 711
2 60478 1 711
2 60479 1 711
2 60480 1 711
2 60481 1 711
2 60482 1 711
2 60483 1 711
2 60484 1 713
2 60485 1 713
2 60486 1 713
2 60487 1 713
2 60488 1 713
2 60489 1 714
2 60490 1 714
2 60491 1 714
2 60492 1 714
2 60493 1 714
2 60494 1 714
2 60495 1 716
2 60496 1 716
2 60497 1 716
2 60498 1 716
2 60499 1 716
2 60500 1 717
2 60501 1 717
2 60502 1 718
2 60503 1 718
2 60504 1 718
2 60505 1 718
2 60506 1 723
2 60507 1 723
2 60508 1 729
2 60509 1 729
2 60510 1 732
2 60511 1 732
2 60512 1 732
2 60513 1 732
2 60514 1 732
2 60515 1 732
2 60516 1 732
2 60517 1 732
2 60518 1 733
2 60519 1 733
2 60520 1 733
2 60521 1 733
2 60522 1 733
2 60523 1 734
2 60524 1 734
2 60525 1 734
2 60526 1 734
2 60527 1 734
2 60528 1 734
2 60529 1 734
2 60530 1 734
2 60531 1 734
2 60532 1 734
2 60533 1 734
2 60534 1 734
2 60535 1 734
2 60536 1 734
2 60537 1 734
2 60538 1 734
2 60539 1 734
2 60540 1 734
2 60541 1 734
2 60542 1 734
2 60543 1 734
2 60544 1 734
2 60545 1 734
2 60546 1 734
2 60547 1 734
2 60548 1 734
2 60549 1 734
2 60550 1 734
2 60551 1 734
2 60552 1 734
2 60553 1 734
2 60554 1 734
2 60555 1 734
2 60556 1 734
2 60557 1 734
2 60558 1 734
2 60559 1 734
2 60560 1 734
2 60561 1 734
2 60562 1 734
2 60563 1 734
2 60564 1 735
2 60565 1 735
2 60566 1 735
2 60567 1 735
2 60568 1 735
2 60569 1 735
2 60570 1 735
2 60571 1 735
2 60572 1 735
2 60573 1 735
2 60574 1 735
2 60575 1 735
2 60576 1 735
2 60577 1 735
2 60578 1 735
2 60579 1 736
2 60580 1 736
2 60581 1 736
2 60582 1 737
2 60583 1 737
2 60584 1 737
2 60585 1 737
2 60586 1 738
2 60587 1 738
2 60588 1 746
2 60589 1 746
2 60590 1 746
2 60591 1 747
2 60592 1 747
2 60593 1 748
2 60594 1 748
2 60595 1 748
2 60596 1 748
2 60597 1 748
2 60598 1 748
2 60599 1 748
2 60600 1 748
2 60601 1 748
2 60602 1 748
2 60603 1 748
2 60604 1 748
2 60605 1 749
2 60606 1 749
2 60607 1 749
2 60608 1 750
2 60609 1 750
2 60610 1 750
2 60611 1 750
2 60612 1 751
2 60613 1 751
2 60614 1 751
2 60615 1 751
2 60616 1 751
2 60617 1 751
2 60618 1 751
2 60619 1 752
2 60620 1 752
2 60621 1 752
2 60622 1 752
2 60623 1 752
2 60624 1 752
2 60625 1 752
2 60626 1 753
2 60627 1 753
2 60628 1 753
2 60629 1 753
2 60630 1 753
2 60631 1 753
2 60632 1 753
2 60633 1 753
2 60634 1 753
2 60635 1 753
2 60636 1 753
2 60637 1 753
2 60638 1 753
2 60639 1 754
2 60640 1 754
2 60641 1 754
2 60642 1 754
2 60643 1 754
2 60644 1 754
2 60645 1 754
2 60646 1 754
2 60647 1 754
2 60648 1 754
2 60649 1 755
2 60650 1 755
2 60651 1 755
2 60652 1 755
2 60653 1 755
2 60654 1 755
2 60655 1 755
2 60656 1 755
2 60657 1 755
2 60658 1 755
2 60659 1 755
2 60660 1 756
2 60661 1 756
2 60662 1 756
2 60663 1 757
2 60664 1 757
2 60665 1 757
2 60666 1 757
2 60667 1 757
2 60668 1 757
2 60669 1 757
2 60670 1 757
2 60671 1 761
2 60672 1 761
2 60673 1 763
2 60674 1 763
2 60675 1 763
2 60676 1 766
2 60677 1 766
2 60678 1 766
2 60679 1 766
2 60680 1 766
2 60681 1 766
2 60682 1 766
2 60683 1 766
2 60684 1 766
2 60685 1 766
2 60686 1 766
2 60687 1 766
2 60688 1 767
2 60689 1 767
2 60690 1 767
2 60691 1 767
2 60692 1 767
2 60693 1 767
2 60694 1 767
2 60695 1 767
2 60696 1 767
2 60697 1 767
2 60698 1 767
2 60699 1 767
2 60700 1 767
2 60701 1 767
2 60702 1 767
2 60703 1 767
2 60704 1 767
2 60705 1 767
2 60706 1 767
2 60707 1 767
2 60708 1 767
2 60709 1 767
2 60710 1 768
2 60711 1 768
2 60712 1 768
2 60713 1 768
2 60714 1 769
2 60715 1 769
2 60716 1 769
2 60717 1 769
2 60718 1 769
2 60719 1 769
2 60720 1 771
2 60721 1 771
2 60722 1 771
2 60723 1 771
2 60724 1 771
2 60725 1 771
2 60726 1 771
2 60727 1 771
2 60728 1 771
2 60729 1 771
2 60730 1 771
2 60731 1 771
2 60732 1 771
2 60733 1 771
2 60734 1 772
2 60735 1 772
2 60736 1 772
2 60737 1 772
2 60738 1 773
2 60739 1 773
2 60740 1 774
2 60741 1 774
2 60742 1 774
2 60743 1 774
2 60744 1 774
2 60745 1 774
2 60746 1 774
2 60747 1 774
2 60748 1 774
2 60749 1 774
2 60750 1 774
2 60751 1 775
2 60752 1 775
2 60753 1 775
2 60754 1 775
2 60755 1 775
2 60756 1 775
2 60757 1 775
2 60758 1 775
2 60759 1 775
2 60760 1 775
2 60761 1 775
2 60762 1 776
2 60763 1 776
2 60764 1 777
2 60765 1 777
2 60766 1 777
2 60767 1 777
2 60768 1 778
2 60769 1 778
2 60770 1 778
2 60771 1 778
2 60772 1 778
2 60773 1 778
2 60774 1 778
2 60775 1 779
2 60776 1 779
2 60777 1 780
2 60778 1 780
2 60779 1 781
2 60780 1 781
2 60781 1 781
2 60782 1 781
2 60783 1 781
2 60784 1 781
2 60785 1 781
2 60786 1 781
2 60787 1 782
2 60788 1 782
2 60789 1 783
2 60790 1 783
2 60791 1 784
2 60792 1 784
2 60793 1 788
2 60794 1 788
2 60795 1 788
2 60796 1 788
2 60797 1 788
2 60798 1 789
2 60799 1 789
2 60800 1 789
2 60801 1 789
2 60802 1 790
2 60803 1 790
2 60804 1 790
2 60805 1 790
2 60806 1 790
2 60807 1 793
2 60808 1 793
2 60809 1 793
2 60810 1 793
2 60811 1 793
2 60812 1 793
2 60813 1 794
2 60814 1 794
2 60815 1 795
2 60816 1 795
2 60817 1 795
2 60818 1 795
2 60819 1 795
2 60820 1 795
2 60821 1 796
2 60822 1 796
2 60823 1 796
2 60824 1 796
2 60825 1 796
2 60826 1 800
2 60827 1 800
2 60828 1 805
2 60829 1 805
2 60830 1 805
2 60831 1 806
2 60832 1 806
2 60833 1 811
2 60834 1 811
2 60835 1 811
2 60836 1 811
2 60837 1 811
2 60838 1 811
2 60839 1 811
2 60840 1 811
2 60841 1 811
2 60842 1 812
2 60843 1 812
2 60844 1 812
2 60845 1 812
2 60846 1 812
2 60847 1 812
2 60848 1 812
2 60849 1 812
2 60850 1 812
2 60851 1 812
2 60852 1 812
2 60853 1 812
2 60854 1 812
2 60855 1 812
2 60856 1 812
2 60857 1 812
2 60858 1 812
2 60859 1 812
2 60860 1 812
2 60861 1 812
2 60862 1 812
2 60863 1 812
2 60864 1 812
2 60865 1 812
2 60866 1 813
2 60867 1 813
2 60868 1 814
2 60869 1 814
2 60870 1 815
2 60871 1 815
2 60872 1 815
2 60873 1 816
2 60874 1 816
2 60875 1 816
2 60876 1 816
2 60877 1 817
2 60878 1 817
2 60879 1 817
2 60880 1 818
2 60881 1 818
2 60882 1 819
2 60883 1 819
2 60884 1 819
2 60885 1 819
2 60886 1 819
2 60887 1 820
2 60888 1 820
2 60889 1 820
2 60890 1 821
2 60891 1 821
2 60892 1 822
2 60893 1 822
2 60894 1 824
2 60895 1 824
2 60896 1 831
2 60897 1 831
2 60898 1 832
2 60899 1 832
2 60900 1 832
2 60901 1 832
2 60902 1 832
2 60903 1 832
2 60904 1 833
2 60905 1 833
2 60906 1 833
2 60907 1 833
2 60908 1 833
2 60909 1 833
2 60910 1 833
2 60911 1 833
2 60912 1 833
2 60913 1 833
2 60914 1 833
2 60915 1 833
2 60916 1 833
2 60917 1 833
2 60918 1 833
2 60919 1 833
2 60920 1 833
2 60921 1 833
2 60922 1 833
2 60923 1 833
2 60924 1 833
2 60925 1 833
2 60926 1 833
2 60927 1 833
2 60928 1 833
2 60929 1 833
2 60930 1 833
2 60931 1 833
2 60932 1 833
2 60933 1 833
2 60934 1 833
2 60935 1 833
2 60936 1 833
2 60937 1 833
2 60938 1 833
2 60939 1 834
2 60940 1 834
2 60941 1 834
2 60942 1 834
2 60943 1 834
2 60944 1 834
2 60945 1 834
2 60946 1 834
2 60947 1 834
2 60948 1 834
2 60949 1 834
2 60950 1 835
2 60951 1 835
2 60952 1 835
2 60953 1 835
2 60954 1 835
2 60955 1 836
2 60956 1 836
2 60957 1 837
2 60958 1 837
2 60959 1 837
2 60960 1 837
2 60961 1 837
2 60962 1 838
2 60963 1 838
2 60964 1 841
2 60965 1 841
2 60966 1 841
2 60967 1 841
2 60968 1 841
2 60969 1 841
2 60970 1 841
2 60971 1 841
2 60972 1 841
2 60973 1 841
2 60974 1 841
2 60975 1 841
2 60976 1 841
2 60977 1 841
2 60978 1 842
2 60979 1 842
2 60980 1 842
2 60981 1 842
2 60982 1 842
2 60983 1 842
2 60984 1 842
2 60985 1 842
2 60986 1 842
2 60987 1 842
2 60988 1 842
2 60989 1 842
2 60990 1 842
2 60991 1 842
2 60992 1 843
2 60993 1 843
2 60994 1 844
2 60995 1 844
2 60996 1 849
2 60997 1 849
2 60998 1 849
2 60999 1 849
2 61000 1 849
2 61001 1 849
2 61002 1 849
2 61003 1 849
2 61004 1 850
2 61005 1 850
2 61006 1 850
2 61007 1 864
2 61008 1 864
2 61009 1 864
2 61010 1 864
2 61011 1 864
2 61012 1 864
2 61013 1 864
2 61014 1 864
2 61015 1 864
2 61016 1 864
2 61017 1 864
2 61018 1 864
2 61019 1 864
2 61020 1 864
2 61021 1 864
2 61022 1 864
2 61023 1 864
2 61024 1 864
2 61025 1 864
2 61026 1 864
2 61027 1 864
2 61028 1 865
2 61029 1 865
2 61030 1 865
2 61031 1 865
2 61032 1 874
2 61033 1 874
2 61034 1 875
2 61035 1 875
2 61036 1 878
2 61037 1 878
2 61038 1 899
2 61039 1 899
2 61040 1 899
2 61041 1 900
2 61042 1 900
2 61043 1 900
2 61044 1 900
2 61045 1 900
2 61046 1 900
2 61047 1 900
2 61048 1 900
2 61049 1 900
2 61050 1 901
2 61051 1 901
2 61052 1 901
2 61053 1 901
2 61054 1 901
2 61055 1 901
2 61056 1 901
2 61057 1 901
2 61058 1 901
2 61059 1 902
2 61060 1 902
2 61061 1 902
2 61062 1 902
2 61063 1 902
2 61064 1 902
2 61065 1 902
2 61066 1 902
2 61067 1 902
2 61068 1 903
2 61069 1 903
2 61070 1 903
2 61071 1 903
2 61072 1 903
2 61073 1 903
2 61074 1 903
2 61075 1 903
2 61076 1 903
2 61077 1 904
2 61078 1 904
2 61079 1 905
2 61080 1 905
2 61081 1 905
2 61082 1 905
2 61083 1 905
2 61084 1 908
2 61085 1 908
2 61086 1 908
2 61087 1 908
2 61088 1 908
2 61089 1 908
2 61090 1 908
2 61091 1 908
2 61092 1 908
2 61093 1 908
2 61094 1 908
2 61095 1 908
2 61096 1 908
2 61097 1 911
2 61098 1 911
2 61099 1 911
2 61100 1 911
2 61101 1 911
2 61102 1 911
2 61103 1 911
2 61104 1 911
2 61105 1 919
2 61106 1 919
2 61107 1 919
2 61108 1 919
2 61109 1 919
2 61110 1 919
2 61111 1 919
2 61112 1 920
2 61113 1 920
2 61114 1 920
2 61115 1 920
2 61116 1 920
2 61117 1 920
2 61118 1 920
2 61119 1 920
2 61120 1 920
2 61121 1 920
2 61122 1 920
2 61123 1 920
2 61124 1 920
2 61125 1 920
2 61126 1 920
2 61127 1 920
2 61128 1 921
2 61129 1 921
2 61130 1 921
2 61131 1 921
2 61132 1 921
2 61133 1 922
2 61134 1 922
2 61135 1 922
2 61136 1 922
2 61137 1 922
2 61138 1 922
2 61139 1 922
2 61140 1 922
2 61141 1 922
2 61142 1 922
2 61143 1 922
2 61144 1 922
2 61145 1 922
2 61146 1 923
2 61147 1 923
2 61148 1 924
2 61149 1 924
2 61150 1 925
2 61151 1 925
2 61152 1 931
2 61153 1 931
2 61154 1 933
2 61155 1 933
2 61156 1 949
2 61157 1 949
2 61158 1 949
2 61159 1 949
2 61160 1 949
2 61161 1 950
2 61162 1 950
2 61163 1 950
2 61164 1 950
2 61165 1 951
2 61166 1 951
2 61167 1 952
2 61168 1 952
2 61169 1 955
2 61170 1 955
2 61171 1 957
2 61172 1 957
2 61173 1 970
2 61174 1 970
2 61175 1 970
2 61176 1 970
2 61177 1 971
2 61178 1 971
2 61179 1 971
2 61180 1 971
2 61181 1 971
2 61182 1 971
2 61183 1 971
2 61184 1 971
2 61185 1 971
2 61186 1 971
2 61187 1 971
2 61188 1 971
2 61189 1 971
2 61190 1 971
2 61191 1 971
2 61192 1 971
2 61193 1 971
2 61194 1 971
2 61195 1 972
2 61196 1 972
2 61197 1 972
2 61198 1 973
2 61199 1 973
2 61200 1 974
2 61201 1 974
2 61202 1 974
2 61203 1 974
2 61204 1 974
2 61205 1 979
2 61206 1 979
2 61207 1 979
2 61208 1 979
2 61209 1 991
2 61210 1 991
2 61211 1 991
2 61212 1 992
2 61213 1 992
2 61214 1 992
2 61215 1 992
2 61216 1 992
2 61217 1 993
2 61218 1 993
2 61219 1 993
2 61220 1 993
2 61221 1 993
2 61222 1 993
2 61223 1 993
2 61224 1 993
2 61225 1 994
2 61226 1 994
2 61227 1 994
2 61228 1 994
2 61229 1 994
2 61230 1 994
2 61231 1 995
2 61232 1 995
2 61233 1 995
2 61234 1 995
2 61235 1 997
2 61236 1 997
2 61237 1 998
2 61238 1 998
2 61239 1 998
2 61240 1 998
2 61241 1 999
2 61242 1 999
2 61243 1 999
2 61244 1 1003
2 61245 1 1003
2 61246 1 1003
2 61247 1 1003
2 61248 1 1003
2 61249 1 1003
2 61250 1 1003
2 61251 1 1003
2 61252 1 1003
2 61253 1 1004
2 61254 1 1004
2 61255 1 1005
2 61256 1 1005
2 61257 1 1005
2 61258 1 1005
2 61259 1 1006
2 61260 1 1006
2 61261 1 1006
2 61262 1 1006
2 61263 1 1006
2 61264 1 1006
2 61265 1 1006
2 61266 1 1009
2 61267 1 1009
2 61268 1 1009
2 61269 1 1009
2 61270 1 1009
2 61271 1 1009
2 61272 1 1009
2 61273 1 1009
2 61274 1 1009
2 61275 1 1010
2 61276 1 1010
2 61277 1 1010
2 61278 1 1010
2 61279 1 1015
2 61280 1 1015
2 61281 1 1015
2 61282 1 1016
2 61283 1 1016
2 61284 1 1016
2 61285 1 1017
2 61286 1 1017
2 61287 1 1019
2 61288 1 1019
2 61289 1 1020
2 61290 1 1020
2 61291 1 1020
2 61292 1 1020
2 61293 1 1020
2 61294 1 1021
2 61295 1 1021
2 61296 1 1021
2 61297 1 1021
2 61298 1 1021
2 61299 1 1021
2 61300 1 1021
2 61301 1 1022
2 61302 1 1022
2 61303 1 1022
2 61304 1 1022
2 61305 1 1022
2 61306 1 1022
2 61307 1 1022
2 61308 1 1022
2 61309 1 1022
2 61310 1 1031
2 61311 1 1031
2 61312 1 1031
2 61313 1 1031
2 61314 1 1032
2 61315 1 1032
2 61316 1 1032
2 61317 1 1033
2 61318 1 1033
2 61319 1 1033
2 61320 1 1033
2 61321 1 1033
2 61322 1 1033
2 61323 1 1033
2 61324 1 1034
2 61325 1 1034
2 61326 1 1034
2 61327 1 1034
2 61328 1 1034
2 61329 1 1034
2 61330 1 1034
2 61331 1 1034
2 61332 1 1034
2 61333 1 1034
2 61334 1 1034
2 61335 1 1034
2 61336 1 1034
2 61337 1 1034
2 61338 1 1034
2 61339 1 1034
2 61340 1 1034
2 61341 1 1034
2 61342 1 1034
2 61343 1 1034
2 61344 1 1034
2 61345 1 1034
2 61346 1 1034
2 61347 1 1034
2 61348 1 1034
2 61349 1 1034
2 61350 1 1034
2 61351 1 1034
2 61352 1 1034
2 61353 1 1034
2 61354 1 1034
2 61355 1 1034
2 61356 1 1034
2 61357 1 1034
2 61358 1 1035
2 61359 1 1035
2 61360 1 1035
2 61361 1 1035
2 61362 1 1036
2 61363 1 1036
2 61364 1 1036
2 61365 1 1036
2 61366 1 1036
2 61367 1 1036
2 61368 1 1036
2 61369 1 1036
2 61370 1 1038
2 61371 1 1038
2 61372 1 1051
2 61373 1 1051
2 61374 1 1052
2 61375 1 1052
2 61376 1 1052
2 61377 1 1053
2 61378 1 1053
2 61379 1 1054
2 61380 1 1054
2 61381 1 1058
2 61382 1 1058
2 61383 1 1063
2 61384 1 1063
2 61385 1 1074
2 61386 1 1074
2 61387 1 1074
2 61388 1 1074
2 61389 1 1074
2 61390 1 1074
2 61391 1 1074
2 61392 1 1074
2 61393 1 1074
2 61394 1 1074
2 61395 1 1075
2 61396 1 1075
2 61397 1 1075
2 61398 1 1075
2 61399 1 1075
2 61400 1 1076
2 61401 1 1076
2 61402 1 1076
2 61403 1 1076
2 61404 1 1076
2 61405 1 1076
2 61406 1 1076
2 61407 1 1079
2 61408 1 1079
2 61409 1 1084
2 61410 1 1084
2 61411 1 1087
2 61412 1 1087
2 61413 1 1087
2 61414 1 1087
2 61415 1 1088
2 61416 1 1088
2 61417 1 1088
2 61418 1 1089
2 61419 1 1089
2 61420 1 1089
2 61421 1 1089
2 61422 1 1090
2 61423 1 1090
2 61424 1 1095
2 61425 1 1095
2 61426 1 1125
2 61427 1 1125
2 61428 1 1127
2 61429 1 1127
2 61430 1 1127
2 61431 1 1128
2 61432 1 1128
2 61433 1 1133
2 61434 1 1133
2 61435 1 1133
2 61436 1 1133
2 61437 1 1133
2 61438 1 1133
2 61439 1 1133
2 61440 1 1133
2 61441 1 1133
2 61442 1 1134
2 61443 1 1134
2 61444 1 1134
2 61445 1 1134
2 61446 1 1135
2 61447 1 1135
2 61448 1 1135
2 61449 1 1135
2 61450 1 1149
2 61451 1 1149
2 61452 1 1149
2 61453 1 1149
2 61454 1 1149
2 61455 1 1149
2 61456 1 1149
2 61457 1 1149
2 61458 1 1149
2 61459 1 1149
2 61460 1 1151
2 61461 1 1151
2 61462 1 1154
2 61463 1 1154
2 61464 1 1154
2 61465 1 1155
2 61466 1 1155
2 61467 1 1155
2 61468 1 1155
2 61469 1 1155
2 61470 1 1155
2 61471 1 1155
2 61472 1 1155
2 61473 1 1155
2 61474 1 1155
2 61475 1 1155
2 61476 1 1155
2 61477 1 1158
2 61478 1 1158
2 61479 1 1158
2 61480 1 1158
2 61481 1 1158
2 61482 1 1158
2 61483 1 1158
2 61484 1 1159
2 61485 1 1159
2 61486 1 1159
2 61487 1 1160
2 61488 1 1160
2 61489 1 1160
2 61490 1 1160
2 61491 1 1161
2 61492 1 1161
2 61493 1 1168
2 61494 1 1168
2 61495 1 1168
2 61496 1 1168
2 61497 1 1168
2 61498 1 1168
2 61499 1 1168
2 61500 1 1168
2 61501 1 1168
2 61502 1 1168
2 61503 1 1168
2 61504 1 1168
2 61505 1 1168
2 61506 1 1169
2 61507 1 1169
2 61508 1 1169
2 61509 1 1169
2 61510 1 1169
2 61511 1 1169
2 61512 1 1170
2 61513 1 1170
2 61514 1 1170
2 61515 1 1170
2 61516 1 1170
2 61517 1 1170
2 61518 1 1170
2 61519 1 1170
2 61520 1 1170
2 61521 1 1170
2 61522 1 1170
2 61523 1 1170
2 61524 1 1170
2 61525 1 1170
2 61526 1 1170
2 61527 1 1170
2 61528 1 1170
2 61529 1 1170
2 61530 1 1170
2 61531 1 1170
2 61532 1 1170
2 61533 1 1170
2 61534 1 1170
2 61535 1 1171
2 61536 1 1171
2 61537 1 1171
2 61538 1 1171
2 61539 1 1171
2 61540 1 1171
2 61541 1 1171
2 61542 1 1171
2 61543 1 1171
2 61544 1 1171
2 61545 1 1171
2 61546 1 1171
2 61547 1 1171
2 61548 1 1171
2 61549 1 1171
2 61550 1 1171
2 61551 1 1171
2 61552 1 1171
2 61553 1 1171
2 61554 1 1171
2 61555 1 1171
2 61556 1 1171
2 61557 1 1171
2 61558 1 1171
2 61559 1 1171
2 61560 1 1171
2 61561 1 1171
2 61562 1 1171
2 61563 1 1171
2 61564 1 1171
2 61565 1 1171
2 61566 1 1171
2 61567 1 1171
2 61568 1 1171
2 61569 1 1171
2 61570 1 1171
2 61571 1 1171
2 61572 1 1171
2 61573 1 1171
2 61574 1 1171
2 61575 1 1171
2 61576 1 1171
2 61577 1 1171
2 61578 1 1171
2 61579 1 1171
2 61580 1 1171
2 61581 1 1171
2 61582 1 1171
2 61583 1 1171
2 61584 1 1171
2 61585 1 1171
2 61586 1 1171
2 61587 1 1171
2 61588 1 1171
2 61589 1 1172
2 61590 1 1172
2 61591 1 1172
2 61592 1 1172
2 61593 1 1172
2 61594 1 1172
2 61595 1 1173
2 61596 1 1173
2 61597 1 1174
2 61598 1 1174
2 61599 1 1175
2 61600 1 1175
2 61601 1 1180
2 61602 1 1180
2 61603 1 1180
2 61604 1 1180
2 61605 1 1181
2 61606 1 1181
2 61607 1 1181
2 61608 1 1181
2 61609 1 1181
2 61610 1 1181
2 61611 1 1181
2 61612 1 1182
2 61613 1 1182
2 61614 1 1183
2 61615 1 1183
2 61616 1 1183
2 61617 1 1194
2 61618 1 1194
2 61619 1 1195
2 61620 1 1195
2 61621 1 1195
2 61622 1 1195
2 61623 1 1196
2 61624 1 1196
2 61625 1 1196
2 61626 1 1196
2 61627 1 1196
2 61628 1 1196
2 61629 1 1196
2 61630 1 1196
2 61631 1 1196
2 61632 1 1196
2 61633 1 1197
2 61634 1 1197
2 61635 1 1197
2 61636 1 1197
2 61637 1 1197
2 61638 1 1199
2 61639 1 1199
2 61640 1 1199
2 61641 1 1199
2 61642 1 1211
2 61643 1 1211
2 61644 1 1217
2 61645 1 1217
2 61646 1 1217
2 61647 1 1217
2 61648 1 1218
2 61649 1 1218
2 61650 1 1218
2 61651 1 1219
2 61652 1 1219
2 61653 1 1219
2 61654 1 1219
2 61655 1 1219
2 61656 1 1219
2 61657 1 1219
2 61658 1 1219
2 61659 1 1219
2 61660 1 1219
2 61661 1 1219
2 61662 1 1219
2 61663 1 1219
2 61664 1 1219
2 61665 1 1220
2 61666 1 1220
2 61667 1 1220
2 61668 1 1220
2 61669 1 1220
2 61670 1 1222
2 61671 1 1222
2 61672 1 1222
2 61673 1 1222
2 61674 1 1222
2 61675 1 1224
2 61676 1 1224
2 61677 1 1224
2 61678 1 1225
2 61679 1 1225
2 61680 1 1226
2 61681 1 1226
2 61682 1 1226
2 61683 1 1226
2 61684 1 1237
2 61685 1 1237
2 61686 1 1238
2 61687 1 1238
2 61688 1 1239
2 61689 1 1239
2 61690 1 1243
2 61691 1 1243
2 61692 1 1243
2 61693 1 1243
2 61694 1 1243
2 61695 1 1243
2 61696 1 1244
2 61697 1 1244
2 61698 1 1244
2 61699 1 1244
2 61700 1 1244
2 61701 1 1244
2 61702 1 1244
2 61703 1 1244
2 61704 1 1244
2 61705 1 1244
2 61706 1 1244
2 61707 1 1244
2 61708 1 1244
2 61709 1 1244
2 61710 1 1244
2 61711 1 1247
2 61712 1 1247
2 61713 1 1247
2 61714 1 1247
2 61715 1 1247
2 61716 1 1247
2 61717 1 1247
2 61718 1 1247
2 61719 1 1247
2 61720 1 1247
2 61721 1 1247
2 61722 1 1248
2 61723 1 1248
2 61724 1 1248
2 61725 1 1249
2 61726 1 1249
2 61727 1 1249
2 61728 1 1249
2 61729 1 1250
2 61730 1 1250
2 61731 1 1250
2 61732 1 1250
2 61733 1 1256
2 61734 1 1256
2 61735 1 1256
2 61736 1 1256
2 61737 1 1256
2 61738 1 1256
2 61739 1 1256
2 61740 1 1256
2 61741 1 1256
2 61742 1 1256
2 61743 1 1256
2 61744 1 1256
2 61745 1 1256
2 61746 1 1256
2 61747 1 1256
2 61748 1 1256
2 61749 1 1256
2 61750 1 1256
2 61751 1 1256
2 61752 1 1256
2 61753 1 1256
2 61754 1 1256
2 61755 1 1256
2 61756 1 1256
2 61757 1 1256
2 61758 1 1256
2 61759 1 1256
2 61760 1 1256
2 61761 1 1256
2 61762 1 1256
2 61763 1 1256
2 61764 1 1256
2 61765 1 1257
2 61766 1 1257
2 61767 1 1257
2 61768 1 1257
2 61769 1 1257
2 61770 1 1257
2 61771 1 1257
2 61772 1 1257
2 61773 1 1257
2 61774 1 1257
2 61775 1 1257
2 61776 1 1257
2 61777 1 1258
2 61778 1 1258
2 61779 1 1258
2 61780 1 1258
2 61781 1 1258
2 61782 1 1259
2 61783 1 1259
2 61784 1 1259
2 61785 1 1259
2 61786 1 1260
2 61787 1 1260
2 61788 1 1261
2 61789 1 1261
2 61790 1 1261
2 61791 1 1261
2 61792 1 1261
2 61793 1 1261
2 61794 1 1261
2 61795 1 1261
2 61796 1 1261
2 61797 1 1261
2 61798 1 1261
2 61799 1 1266
2 61800 1 1266
2 61801 1 1266
2 61802 1 1266
2 61803 1 1266
2 61804 1 1266
2 61805 1 1267
2 61806 1 1267
2 61807 1 1267
2 61808 1 1267
2 61809 1 1271
2 61810 1 1271
2 61811 1 1280
2 61812 1 1280
2 61813 1 1280
2 61814 1 1282
2 61815 1 1282
2 61816 1 1282
2 61817 1 1282
2 61818 1 1282
2 61819 1 1282
2 61820 1 1282
2 61821 1 1282
2 61822 1 1282
2 61823 1 1282
2 61824 1 1282
2 61825 1 1282
2 61826 1 1283
2 61827 1 1283
2 61828 1 1283
2 61829 1 1283
2 61830 1 1283
2 61831 1 1283
2 61832 1 1283
2 61833 1 1285
2 61834 1 1285
2 61835 1 1285
2 61836 1 1285
2 61837 1 1285
2 61838 1 1285
2 61839 1 1285
2 61840 1 1285
2 61841 1 1285
2 61842 1 1285
2 61843 1 1285
2 61844 1 1285
2 61845 1 1299
2 61846 1 1299
2 61847 1 1300
2 61848 1 1300
2 61849 1 1300
2 61850 1 1300
2 61851 1 1300
2 61852 1 1300
2 61853 1 1302
2 61854 1 1302
2 61855 1 1305
2 61856 1 1305
2 61857 1 1305
2 61858 1 1305
2 61859 1 1305
2 61860 1 1305
2 61861 1 1305
2 61862 1 1305
2 61863 1 1306
2 61864 1 1306
2 61865 1 1306
2 61866 1 1306
2 61867 1 1306
2 61868 1 1306
2 61869 1 1306
2 61870 1 1306
2 61871 1 1317
2 61872 1 1317
2 61873 1 1318
2 61874 1 1318
2 61875 1 1318
2 61876 1 1318
2 61877 1 1319
2 61878 1 1319
2 61879 1 1320
2 61880 1 1320
2 61881 1 1320
2 61882 1 1323
2 61883 1 1323
2 61884 1 1323
2 61885 1 1323
2 61886 1 1323
2 61887 1 1323
2 61888 1 1323
2 61889 1 1323
2 61890 1 1323
2 61891 1 1323
2 61892 1 1323
2 61893 1 1323
2 61894 1 1323
2 61895 1 1323
2 61896 1 1323
2 61897 1 1323
2 61898 1 1323
2 61899 1 1323
2 61900 1 1323
2 61901 1 1323
2 61902 1 1323
2 61903 1 1323
2 61904 1 1323
2 61905 1 1323
2 61906 1 1323
2 61907 1 1323
2 61908 1 1323
2 61909 1 1323
2 61910 1 1323
2 61911 1 1323
2 61912 1 1323
2 61913 1 1323
2 61914 1 1323
2 61915 1 1323
2 61916 1 1323
2 61917 1 1323
2 61918 1 1324
2 61919 1 1324
2 61920 1 1324
2 61921 1 1324
2 61922 1 1324
2 61923 1 1324
2 61924 1 1324
2 61925 1 1324
2 61926 1 1325
2 61927 1 1325
2 61928 1 1325
2 61929 1 1326
2 61930 1 1326
2 61931 1 1329
2 61932 1 1329
2 61933 1 1329
2 61934 1 1329
2 61935 1 1329
2 61936 1 1329
2 61937 1 1329
2 61938 1 1329
2 61939 1 1329
2 61940 1 1329
2 61941 1 1329
2 61942 1 1330
2 61943 1 1330
2 61944 1 1330
2 61945 1 1345
2 61946 1 1345
2 61947 1 1345
2 61948 1 1345
2 61949 1 1345
2 61950 1 1345
2 61951 1 1345
2 61952 1 1346
2 61953 1 1346
2 61954 1 1346
2 61955 1 1347
2 61956 1 1347
2 61957 1 1347
2 61958 1 1347
2 61959 1 1347
2 61960 1 1347
2 61961 1 1347
2 61962 1 1348
2 61963 1 1348
2 61964 1 1348
2 61965 1 1349
2 61966 1 1349
2 61967 1 1354
2 61968 1 1354
2 61969 1 1354
2 61970 1 1355
2 61971 1 1355
2 61972 1 1355
2 61973 1 1355
2 61974 1 1355
2 61975 1 1355
2 61976 1 1355
2 61977 1 1355
2 61978 1 1355
2 61979 1 1355
2 61980 1 1355
2 61981 1 1355
2 61982 1 1355
2 61983 1 1355
2 61984 1 1355
2 61985 1 1356
2 61986 1 1356
2 61987 1 1357
2 61988 1 1357
2 61989 1 1357
2 61990 1 1357
2 61991 1 1357
2 61992 1 1357
2 61993 1 1360
2 61994 1 1360
2 61995 1 1360
2 61996 1 1360
2 61997 1 1360
2 61998 1 1363
2 61999 1 1363
2 62000 1 1364
2 62001 1 1364
2 62002 1 1372
2 62003 1 1372
2 62004 1 1372
2 62005 1 1372
2 62006 1 1372
2 62007 1 1372
2 62008 1 1372
2 62009 1 1372
2 62010 1 1372
2 62011 1 1372
2 62012 1 1372
2 62013 1 1374
2 62014 1 1374
2 62015 1 1374
2 62016 1 1376
2 62017 1 1376
2 62018 1 1377
2 62019 1 1377
2 62020 1 1377
2 62021 1 1377
2 62022 1 1379
2 62023 1 1379
2 62024 1 1389
2 62025 1 1389
2 62026 1 1389
2 62027 1 1389
2 62028 1 1390
2 62029 1 1390
2 62030 1 1390
2 62031 1 1391
2 62032 1 1391
2 62033 1 1391
2 62034 1 1391
2 62035 1 1391
2 62036 1 1392
2 62037 1 1392
2 62038 1 1392
2 62039 1 1392
2 62040 1 1392
2 62041 1 1392
2 62042 1 1392
2 62043 1 1392
2 62044 1 1392
2 62045 1 1397
2 62046 1 1397
2 62047 1 1397
2 62048 1 1397
2 62049 1 1397
2 62050 1 1398
2 62051 1 1398
2 62052 1 1398
2 62053 1 1398
2 62054 1 1398
2 62055 1 1398
2 62056 1 1398
2 62057 1 1398
2 62058 1 1398
2 62059 1 1398
2 62060 1 1398
2 62061 1 1398
2 62062 1 1398
2 62063 1 1398
2 62064 1 1398
2 62065 1 1398
2 62066 1 1398
2 62067 1 1398
2 62068 1 1399
2 62069 1 1399
2 62070 1 1399
2 62071 1 1399
2 62072 1 1399
2 62073 1 1399
2 62074 1 1399
2 62075 1 1400
2 62076 1 1400
2 62077 1 1400
2 62078 1 1400
2 62079 1 1400
2 62080 1 1400
2 62081 1 1401
2 62082 1 1401
2 62083 1 1401
2 62084 1 1401
2 62085 1 1401
2 62086 1 1401
2 62087 1 1402
2 62088 1 1402
2 62089 1 1402
2 62090 1 1402
2 62091 1 1402
2 62092 1 1402
2 62093 1 1409
2 62094 1 1409
2 62095 1 1409
2 62096 1 1409
2 62097 1 1409
2 62098 1 1409
2 62099 1 1409
2 62100 1 1410
2 62101 1 1410
2 62102 1 1410
2 62103 1 1410
2 62104 1 1410
2 62105 1 1411
2 62106 1 1411
2 62107 1 1411
2 62108 1 1411
2 62109 1 1411
2 62110 1 1411
2 62111 1 1412
2 62112 1 1412
2 62113 1 1412
2 62114 1 1412
2 62115 1 1412
2 62116 1 1412
2 62117 1 1412
2 62118 1 1412
2 62119 1 1412
2 62120 1 1413
2 62121 1 1413
2 62122 1 1413
2 62123 1 1413
2 62124 1 1413
2 62125 1 1413
2 62126 1 1413
2 62127 1 1413
2 62128 1 1413
2 62129 1 1413
2 62130 1 1413
2 62131 1 1413
2 62132 1 1413
2 62133 1 1422
2 62134 1 1422
2 62135 1 1422
2 62136 1 1422
2 62137 1 1422
2 62138 1 1422
2 62139 1 1422
2 62140 1 1422
2 62141 1 1422
2 62142 1 1422
2 62143 1 1423
2 62144 1 1423
2 62145 1 1425
2 62146 1 1425
2 62147 1 1427
2 62148 1 1427
2 62149 1 1427
2 62150 1 1427
2 62151 1 1427
2 62152 1 1427
2 62153 1 1428
2 62154 1 1428
2 62155 1 1428
2 62156 1 1428
2 62157 1 1428
2 62158 1 1428
2 62159 1 1428
2 62160 1 1428
2 62161 1 1428
2 62162 1 1428
2 62163 1 1428
2 62164 1 1428
2 62165 1 1428
2 62166 1 1429
2 62167 1 1429
2 62168 1 1429
2 62169 1 1429
2 62170 1 1429
2 62171 1 1429
2 62172 1 1429
2 62173 1 1429
2 62174 1 1429
2 62175 1 1429
2 62176 1 1429
2 62177 1 1429
2 62178 1 1429
2 62179 1 1429
2 62180 1 1429
2 62181 1 1430
2 62182 1 1430
2 62183 1 1430
2 62184 1 1431
2 62185 1 1431
2 62186 1 1442
2 62187 1 1442
2 62188 1 1442
2 62189 1 1442
2 62190 1 1442
2 62191 1 1442
2 62192 1 1442
2 62193 1 1442
2 62194 1 1442
2 62195 1 1442
2 62196 1 1442
2 62197 1 1443
2 62198 1 1443
2 62199 1 1443
2 62200 1 1443
2 62201 1 1443
2 62202 1 1444
2 62203 1 1444
2 62204 1 1444
2 62205 1 1446
2 62206 1 1446
2 62207 1 1446
2 62208 1 1446
2 62209 1 1446
2 62210 1 1446
2 62211 1 1446
2 62212 1 1446
2 62213 1 1446
2 62214 1 1446
2 62215 1 1446
2 62216 1 1447
2 62217 1 1447
2 62218 1 1457
2 62219 1 1457
2 62220 1 1457
2 62221 1 1458
2 62222 1 1458
2 62223 1 1458
2 62224 1 1460
2 62225 1 1460
2 62226 1 1461
2 62227 1 1461
2 62228 1 1461
2 62229 1 1462
2 62230 1 1462
2 62231 1 1463
2 62232 1 1463
2 62233 1 1463
2 62234 1 1467
2 62235 1 1467
2 62236 1 1467
2 62237 1 1468
2 62238 1 1468
2 62239 1 1470
2 62240 1 1470
2 62241 1 1470
2 62242 1 1470
2 62243 1 1470
2 62244 1 1472
2 62245 1 1472
2 62246 1 1483
2 62247 1 1483
2 62248 1 1483
2 62249 1 1483
2 62250 1 1483
2 62251 1 1483
2 62252 1 1484
2 62253 1 1484
2 62254 1 1485
2 62255 1 1485
2 62256 1 1485
2 62257 1 1485
2 62258 1 1485
2 62259 1 1485
2 62260 1 1485
2 62261 1 1485
2 62262 1 1485
2 62263 1 1485
2 62264 1 1487
2 62265 1 1487
2 62266 1 1487
2 62267 1 1487
2 62268 1 1488
2 62269 1 1488
2 62270 1 1488
2 62271 1 1488
2 62272 1 1488
2 62273 1 1488
2 62274 1 1488
2 62275 1 1490
2 62276 1 1490
2 62277 1 1497
2 62278 1 1497
2 62279 1 1497
2 62280 1 1497
2 62281 1 1497
2 62282 1 1497
2 62283 1 1497
2 62284 1 1498
2 62285 1 1498
2 62286 1 1498
2 62287 1 1504
2 62288 1 1504
2 62289 1 1505
2 62290 1 1505
2 62291 1 1505
2 62292 1 1512
2 62293 1 1512
2 62294 1 1512
2 62295 1 1514
2 62296 1 1514
2 62297 1 1514
2 62298 1 1514
2 62299 1 1516
2 62300 1 1516
2 62301 1 1516
2 62302 1 1516
2 62303 1 1516
2 62304 1 1516
2 62305 1 1516
2 62306 1 1516
2 62307 1 1516
2 62308 1 1516
2 62309 1 1516
2 62310 1 1516
2 62311 1 1516
2 62312 1 1520
2 62313 1 1520
2 62314 1 1520
2 62315 1 1523
2 62316 1 1523
2 62317 1 1523
2 62318 1 1523
2 62319 1 1523
2 62320 1 1523
2 62321 1 1523
2 62322 1 1523
2 62323 1 1523
2 62324 1 1523
2 62325 1 1523
2 62326 1 1523
2 62327 1 1523
2 62328 1 1523
2 62329 1 1523
2 62330 1 1523
2 62331 1 1523
2 62332 1 1523
2 62333 1 1524
2 62334 1 1524
2 62335 1 1524
2 62336 1 1524
2 62337 1 1524
2 62338 1 1524
2 62339 1 1524
2 62340 1 1524
2 62341 1 1524
2 62342 1 1524
2 62343 1 1525
2 62344 1 1525
2 62345 1 1525
2 62346 1 1526
2 62347 1 1526
2 62348 1 1526
2 62349 1 1528
2 62350 1 1528
2 62351 1 1545
2 62352 1 1545
2 62353 1 1545
2 62354 1 1545
2 62355 1 1545
2 62356 1 1545
2 62357 1 1545
2 62358 1 1545
2 62359 1 1545
2 62360 1 1545
2 62361 1 1545
2 62362 1 1545
2 62363 1 1545
2 62364 1 1545
2 62365 1 1546
2 62366 1 1546
2 62367 1 1546
2 62368 1 1546
2 62369 1 1546
2 62370 1 1546
2 62371 1 1546
2 62372 1 1546
2 62373 1 1546
2 62374 1 1546
2 62375 1 1546
2 62376 1 1546
2 62377 1 1547
2 62378 1 1547
2 62379 1 1547
2 62380 1 1547
2 62381 1 1547
2 62382 1 1548
2 62383 1 1548
2 62384 1 1548
2 62385 1 1548
2 62386 1 1568
2 62387 1 1568
2 62388 1 1570
2 62389 1 1570
2 62390 1 1570
2 62391 1 1570
2 62392 1 1570
2 62393 1 1571
2 62394 1 1571
2 62395 1 1571
2 62396 1 1571
2 62397 1 1571
2 62398 1 1571
2 62399 1 1571
2 62400 1 1571
2 62401 1 1571
2 62402 1 1571
2 62403 1 1571
2 62404 1 1571
2 62405 1 1571
2 62406 1 1571
2 62407 1 1571
2 62408 1 1571
2 62409 1 1571
2 62410 1 1571
2 62411 1 1571
2 62412 1 1571
2 62413 1 1571
2 62414 1 1571
2 62415 1 1571
2 62416 1 1571
2 62417 1 1571
2 62418 1 1571
2 62419 1 1572
2 62420 1 1572
2 62421 1 1572
2 62422 1 1572
2 62423 1 1591
2 62424 1 1591
2 62425 1 1591
2 62426 1 1591
2 62427 1 1591
2 62428 1 1591
2 62429 1 1591
2 62430 1 1591
2 62431 1 1592
2 62432 1 1592
2 62433 1 1592
2 62434 1 1592
2 62435 1 1592
2 62436 1 1592
2 62437 1 1592
2 62438 1 1592
2 62439 1 1592
2 62440 1 1592
2 62441 1 1592
2 62442 1 1593
2 62443 1 1593
2 62444 1 1593
2 62445 1 1593
2 62446 1 1593
2 62447 1 1593
2 62448 1 1593
2 62449 1 1594
2 62450 1 1594
2 62451 1 1595
2 62452 1 1595
2 62453 1 1595
2 62454 1 1595
2 62455 1 1595
2 62456 1 1595
2 62457 1 1595
2 62458 1 1595
2 62459 1 1595
2 62460 1 1598
2 62461 1 1598
2 62462 1 1598
2 62463 1 1599
2 62464 1 1599
2 62465 1 1600
2 62466 1 1600
2 62467 1 1600
2 62468 1 1600
2 62469 1 1601
2 62470 1 1601
2 62471 1 1601
2 62472 1 1601
2 62473 1 1601
2 62474 1 1601
2 62475 1 1601
2 62476 1 1601
2 62477 1 1601
2 62478 1 1601
2 62479 1 1601
2 62480 1 1601
2 62481 1 1601
2 62482 1 1601
2 62483 1 1601
2 62484 1 1601
2 62485 1 1601
2 62486 1 1601
2 62487 1 1601
2 62488 1 1601
2 62489 1 1601
2 62490 1 1601
2 62491 1 1601
2 62492 1 1601
2 62493 1 1601
2 62494 1 1601
2 62495 1 1601
2 62496 1 1601
2 62497 1 1601
2 62498 1 1601
2 62499 1 1601
2 62500 1 1601
2 62501 1 1601
2 62502 1 1601
2 62503 1 1601
2 62504 1 1601
2 62505 1 1601
2 62506 1 1601
2 62507 1 1601
2 62508 1 1601
2 62509 1 1601
2 62510 1 1601
2 62511 1 1601
2 62512 1 1601
2 62513 1 1602
2 62514 1 1602
2 62515 1 1602
2 62516 1 1602
2 62517 1 1602
2 62518 1 1602
2 62519 1 1602
2 62520 1 1602
2 62521 1 1602
2 62522 1 1602
2 62523 1 1602
2 62524 1 1602
2 62525 1 1602
2 62526 1 1602
2 62527 1 1602
2 62528 1 1602
2 62529 1 1602
2 62530 1 1602
2 62531 1 1602
2 62532 1 1602
2 62533 1 1602
2 62534 1 1602
2 62535 1 1602
2 62536 1 1602
2 62537 1 1602
2 62538 1 1602
2 62539 1 1602
2 62540 1 1602
2 62541 1 1602
2 62542 1 1602
2 62543 1 1602
2 62544 1 1602
2 62545 1 1602
2 62546 1 1602
2 62547 1 1602
2 62548 1 1602
2 62549 1 1602
2 62550 1 1602
2 62551 1 1602
2 62552 1 1602
2 62553 1 1602
2 62554 1 1602
2 62555 1 1602
2 62556 1 1602
2 62557 1 1602
2 62558 1 1602
2 62559 1 1602
2 62560 1 1602
2 62561 1 1602
2 62562 1 1602
2 62563 1 1602
2 62564 1 1602
2 62565 1 1602
2 62566 1 1602
2 62567 1 1602
2 62568 1 1602
2 62569 1 1602
2 62570 1 1602
2 62571 1 1602
2 62572 1 1602
2 62573 1 1602
2 62574 1 1602
2 62575 1 1602
2 62576 1 1602
2 62577 1 1602
2 62578 1 1602
2 62579 1 1602
2 62580 1 1602
2 62581 1 1602
2 62582 1 1602
2 62583 1 1602
2 62584 1 1602
2 62585 1 1602
2 62586 1 1602
2 62587 1 1602
2 62588 1 1602
2 62589 1 1602
2 62590 1 1602
2 62591 1 1602
2 62592 1 1603
2 62593 1 1603
2 62594 1 1603
2 62595 1 1603
2 62596 1 1603
2 62597 1 1603
2 62598 1 1603
2 62599 1 1603
2 62600 1 1604
2 62601 1 1604
2 62602 1 1605
2 62603 1 1605
2 62604 1 1605
2 62605 1 1605
2 62606 1 1605
2 62607 1 1605
2 62608 1 1605
2 62609 1 1605
2 62610 1 1605
2 62611 1 1605
2 62612 1 1605
2 62613 1 1605
2 62614 1 1605
2 62615 1 1606
2 62616 1 1606
2 62617 1 1606
2 62618 1 1615
2 62619 1 1615
2 62620 1 1617
2 62621 1 1617
2 62622 1 1618
2 62623 1 1618
2 62624 1 1627
2 62625 1 1627
2 62626 1 1630
2 62627 1 1630
2 62628 1 1630
2 62629 1 1630
2 62630 1 1630
2 62631 1 1630
2 62632 1 1630
2 62633 1 1630
2 62634 1 1630
2 62635 1 1630
2 62636 1 1630
2 62637 1 1630
2 62638 1 1630
2 62639 1 1630
2 62640 1 1630
2 62641 1 1630
2 62642 1 1630
2 62643 1 1630
2 62644 1 1630
2 62645 1 1630
2 62646 1 1638
2 62647 1 1638
2 62648 1 1638
2 62649 1 1638
2 62650 1 1638
2 62651 1 1638
2 62652 1 1638
2 62653 1 1639
2 62654 1 1639
2 62655 1 1639
2 62656 1 1640
2 62657 1 1640
2 62658 1 1641
2 62659 1 1641
2 62660 1 1641
2 62661 1 1641
2 62662 1 1642
2 62663 1 1642
2 62664 1 1643
2 62665 1 1643
2 62666 1 1643
2 62667 1 1643
2 62668 1 1644
2 62669 1 1644
2 62670 1 1646
2 62671 1 1646
2 62672 1 1657
2 62673 1 1657
2 62674 1 1657
2 62675 1 1657
2 62676 1 1657
2 62677 1 1657
2 62678 1 1657
2 62679 1 1657
2 62680 1 1657
2 62681 1 1657
2 62682 1 1657
2 62683 1 1657
2 62684 1 1657
2 62685 1 1657
2 62686 1 1657
2 62687 1 1657
2 62688 1 1657
2 62689 1 1657
2 62690 1 1657
2 62691 1 1658
2 62692 1 1658
2 62693 1 1659
2 62694 1 1659
2 62695 1 1659
2 62696 1 1660
2 62697 1 1660
2 62698 1 1665
2 62699 1 1665
2 62700 1 1673
2 62701 1 1673
2 62702 1 1673
2 62703 1 1673
2 62704 1 1673
2 62705 1 1673
2 62706 1 1673
2 62707 1 1673
2 62708 1 1673
2 62709 1 1673
2 62710 1 1673
2 62711 1 1673
2 62712 1 1673
2 62713 1 1673
2 62714 1 1673
2 62715 1 1673
2 62716 1 1673
2 62717 1 1673
2 62718 1 1673
2 62719 1 1673
2 62720 1 1673
2 62721 1 1673
2 62722 1 1673
2 62723 1 1673
2 62724 1 1673
2 62725 1 1673
2 62726 1 1673
2 62727 1 1673
2 62728 1 1673
2 62729 1 1673
2 62730 1 1673
2 62731 1 1673
2 62732 1 1673
2 62733 1 1673
2 62734 1 1673
2 62735 1 1673
2 62736 1 1673
2 62737 1 1673
2 62738 1 1673
2 62739 1 1674
2 62740 1 1674
2 62741 1 1674
2 62742 1 1674
2 62743 1 1674
2 62744 1 1674
2 62745 1 1674
2 62746 1 1674
2 62747 1 1675
2 62748 1 1675
2 62749 1 1676
2 62750 1 1676
2 62751 1 1678
2 62752 1 1678
2 62753 1 1678
2 62754 1 1678
2 62755 1 1678
2 62756 1 1678
2 62757 1 1678
2 62758 1 1678
2 62759 1 1678
2 62760 1 1678
2 62761 1 1678
2 62762 1 1680
2 62763 1 1680
2 62764 1 1685
2 62765 1 1685
2 62766 1 1685
2 62767 1 1685
2 62768 1 1685
2 62769 1 1687
2 62770 1 1687
2 62771 1 1687
2 62772 1 1687
2 62773 1 1688
2 62774 1 1688
2 62775 1 1688
2 62776 1 1688
2 62777 1 1688
2 62778 1 1688
2 62779 1 1688
2 62780 1 1688
2 62781 1 1688
2 62782 1 1688
2 62783 1 1688
2 62784 1 1690
2 62785 1 1690
2 62786 1 1701
2 62787 1 1701
2 62788 1 1701
2 62789 1 1701
2 62790 1 1702
2 62791 1 1702
2 62792 1 1702
2 62793 1 1702
2 62794 1 1705
2 62795 1 1705
2 62796 1 1705
2 62797 1 1706
2 62798 1 1706
2 62799 1 1706
2 62800 1 1706
2 62801 1 1706
2 62802 1 1706
2 62803 1 1706
2 62804 1 1706
2 62805 1 1706
2 62806 1 1706
2 62807 1 1706
2 62808 1 1706
2 62809 1 1711
2 62810 1 1711
2 62811 1 1712
2 62812 1 1712
2 62813 1 1713
2 62814 1 1713
2 62815 1 1713
2 62816 1 1713
2 62817 1 1715
2 62818 1 1715
2 62819 1 1716
2 62820 1 1716
2 62821 1 1724
2 62822 1 1724
2 62823 1 1724
2 62824 1 1724
2 62825 1 1724
2 62826 1 1724
2 62827 1 1724
2 62828 1 1724
2 62829 1 1724
2 62830 1 1724
2 62831 1 1724
2 62832 1 1725
2 62833 1 1725
2 62834 1 1725
2 62835 1 1725
2 62836 1 1726
2 62837 1 1726
2 62838 1 1727
2 62839 1 1727
2 62840 1 1727
2 62841 1 1727
2 62842 1 1727
2 62843 1 1727
2 62844 1 1727
2 62845 1 1727
2 62846 1 1727
2 62847 1 1727
2 62848 1 1738
2 62849 1 1738
2 62850 1 1738
2 62851 1 1738
2 62852 1 1738
2 62853 1 1741
2 62854 1 1741
2 62855 1 1741
2 62856 1 1741
2 62857 1 1741
2 62858 1 1742
2 62859 1 1742
2 62860 1 1743
2 62861 1 1743
2 62862 1 1750
2 62863 1 1750
2 62864 1 1750
2 62865 1 1750
2 62866 1 1750
2 62867 1 1751
2 62868 1 1751
2 62869 1 1751
2 62870 1 1758
2 62871 1 1758
2 62872 1 1759
2 62873 1 1759
2 62874 1 1761
2 62875 1 1761
2 62876 1 1763
2 62877 1 1763
2 62878 1 1763
2 62879 1 1763
2 62880 1 1763
2 62881 1 1763
2 62882 1 1779
2 62883 1 1779
2 62884 1 1779
2 62885 1 1779
2 62886 1 1779
2 62887 1 1779
2 62888 1 1779
2 62889 1 1779
2 62890 1 1779
2 62891 1 1779
2 62892 1 1779
2 62893 1 1779
2 62894 1 1779
2 62895 1 1779
2 62896 1 1779
2 62897 1 1779
2 62898 1 1779
2 62899 1 1779
2 62900 1 1779
2 62901 1 1779
2 62902 1 1779
2 62903 1 1779
2 62904 1 1779
2 62905 1 1779
2 62906 1 1779
2 62907 1 1779
2 62908 1 1779
2 62909 1 1779
2 62910 1 1779
2 62911 1 1779
2 62912 1 1779
2 62913 1 1779
2 62914 1 1779
2 62915 1 1779
2 62916 1 1779
2 62917 1 1779
2 62918 1 1779
2 62919 1 1779
2 62920 1 1779
2 62921 1 1779
2 62922 1 1779
2 62923 1 1779
2 62924 1 1779
2 62925 1 1779
2 62926 1 1779
2 62927 1 1779
2 62928 1 1779
2 62929 1 1779
2 62930 1 1779
2 62931 1 1779
2 62932 1 1779
2 62933 1 1779
2 62934 1 1779
2 62935 1 1779
2 62936 1 1779
2 62937 1 1779
2 62938 1 1779
2 62939 1 1780
2 62940 1 1780
2 62941 1 1780
2 62942 1 1780
2 62943 1 1780
2 62944 1 1780
2 62945 1 1780
2 62946 1 1780
2 62947 1 1780
2 62948 1 1780
2 62949 1 1780
2 62950 1 1780
2 62951 1 1780
2 62952 1 1780
2 62953 1 1780
2 62954 1 1780
2 62955 1 1780
2 62956 1 1780
2 62957 1 1780
2 62958 1 1780
2 62959 1 1780
2 62960 1 1780
2 62961 1 1780
2 62962 1 1780
2 62963 1 1780
2 62964 1 1780
2 62965 1 1780
2 62966 1 1780
2 62967 1 1780
2 62968 1 1780
2 62969 1 1780
2 62970 1 1780
2 62971 1 1780
2 62972 1 1780
2 62973 1 1780
2 62974 1 1780
2 62975 1 1780
2 62976 1 1780
2 62977 1 1780
2 62978 1 1780
2 62979 1 1780
2 62980 1 1780
2 62981 1 1780
2 62982 1 1780
2 62983 1 1780
2 62984 1 1780
2 62985 1 1780
2 62986 1 1780
2 62987 1 1780
2 62988 1 1780
2 62989 1 1780
2 62990 1 1780
2 62991 1 1780
2 62992 1 1780
2 62993 1 1780
2 62994 1 1780
2 62995 1 1780
2 62996 1 1780
2 62997 1 1780
2 62998 1 1781
2 62999 1 1781
2 63000 1 1781
2 63001 1 1782
2 63002 1 1782
2 63003 1 1783
2 63004 1 1783
2 63005 1 1783
2 63006 1 1783
2 63007 1 1784
2 63008 1 1784
2 63009 1 1784
2 63010 1 1784
2 63011 1 1784
2 63012 1 1784
2 63013 1 1784
2 63014 1 1784
2 63015 1 1784
2 63016 1 1784
2 63017 1 1784
2 63018 1 1784
2 63019 1 1784
2 63020 1 1784
2 63021 1 1784
2 63022 1 1786
2 63023 1 1786
2 63024 1 1786
2 63025 1 1786
2 63026 1 1787
2 63027 1 1787
2 63028 1 1788
2 63029 1 1788
2 63030 1 1788
2 63031 1 1788
2 63032 1 1788
2 63033 1 1788
2 63034 1 1790
2 63035 1 1790
2 63036 1 1790
2 63037 1 1790
2 63038 1 1790
2 63039 1 1791
2 63040 1 1791
2 63041 1 1797
2 63042 1 1797
2 63043 1 1797
2 63044 1 1802
2 63045 1 1802
2 63046 1 1812
2 63047 1 1812
2 63048 1 1812
2 63049 1 1817
2 63050 1 1817
2 63051 1 1817
2 63052 1 1818
2 63053 1 1818
2 63054 1 1818
2 63055 1 1818
2 63056 1 1819
2 63057 1 1819
2 63058 1 1827
2 63059 1 1827
2 63060 1 1827
2 63061 1 1827
2 63062 1 1827
2 63063 1 1827
2 63064 1 1827
2 63065 1 1828
2 63066 1 1828
2 63067 1 1828
2 63068 1 1828
2 63069 1 1828
2 63070 1 1828
2 63071 1 1828
2 63072 1 1828
2 63073 1 1828
2 63074 1 1828
2 63075 1 1828
2 63076 1 1828
2 63077 1 1828
2 63078 1 1828
2 63079 1 1828
2 63080 1 1828
2 63081 1 1828
2 63082 1 1828
2 63083 1 1828
2 63084 1 1828
2 63085 1 1828
2 63086 1 1828
2 63087 1 1828
2 63088 1 1828
2 63089 1 1828
2 63090 1 1828
2 63091 1 1828
2 63092 1 1828
2 63093 1 1829
2 63094 1 1829
2 63095 1 1829
2 63096 1 1833
2 63097 1 1833
2 63098 1 1835
2 63099 1 1835
2 63100 1 1836
2 63101 1 1836
2 63102 1 1836
2 63103 1 1838
2 63104 1 1838
2 63105 1 1838
2 63106 1 1839
2 63107 1 1839
2 63108 1 1839
2 63109 1 1839
2 63110 1 1839
2 63111 1 1851
2 63112 1 1851
2 63113 1 1851
2 63114 1 1851
2 63115 1 1851
2 63116 1 1853
2 63117 1 1853
2 63118 1 1854
2 63119 1 1854
2 63120 1 1854
2 63121 1 1854
2 63122 1 1854
2 63123 1 1854
2 63124 1 1854
2 63125 1 1855
2 63126 1 1855
2 63127 1 1855
2 63128 1 1856
2 63129 1 1856
2 63130 1 1856
2 63131 1 1856
2 63132 1 1856
2 63133 1 1856
2 63134 1 1856
2 63135 1 1857
2 63136 1 1857
2 63137 1 1857
2 63138 1 1857
2 63139 1 1857
2 63140 1 1857
2 63141 1 1858
2 63142 1 1858
2 63143 1 1858
2 63144 1 1858
2 63145 1 1859
2 63146 1 1859
2 63147 1 1859
2 63148 1 1860
2 63149 1 1860
2 63150 1 1865
2 63151 1 1865
2 63152 1 1865
2 63153 1 1865
2 63154 1 1866
2 63155 1 1866
2 63156 1 1866
2 63157 1 1866
2 63158 1 1871
2 63159 1 1871
2 63160 1 1873
2 63161 1 1873
2 63162 1 1873
2 63163 1 1873
2 63164 1 1873
2 63165 1 1873
2 63166 1 1873
2 63167 1 1873
2 63168 1 1880
2 63169 1 1880
2 63170 1 1880
2 63171 1 1880
2 63172 1 1880
2 63173 1 1880
2 63174 1 1880
2 63175 1 1880
2 63176 1 1880
2 63177 1 1880
2 63178 1 1880
2 63179 1 1880
2 63180 1 1880
2 63181 1 1880
2 63182 1 1880
2 63183 1 1880
2 63184 1 1880
2 63185 1 1880
2 63186 1 1881
2 63187 1 1881
2 63188 1 1881
2 63189 1 1884
2 63190 1 1884
2 63191 1 1884
2 63192 1 1884
2 63193 1 1884
2 63194 1 1885
2 63195 1 1885
2 63196 1 1887
2 63197 1 1887
2 63198 1 1892
2 63199 1 1892
2 63200 1 1892
2 63201 1 1892
2 63202 1 1892
2 63203 1 1892
2 63204 1 1892
2 63205 1 1892
2 63206 1 1892
2 63207 1 1892
2 63208 1 1892
2 63209 1 1892
2 63210 1 1892
2 63211 1 1892
2 63212 1 1892
2 63213 1 1892
2 63214 1 1893
2 63215 1 1893
2 63216 1 1893
2 63217 1 1893
2 63218 1 1894
2 63219 1 1894
2 63220 1 1894
2 63221 1 1894
2 63222 1 1894
2 63223 1 1894
2 63224 1 1894
2 63225 1 1894
2 63226 1 1894
2 63227 1 1894
2 63228 1 1895
2 63229 1 1895
2 63230 1 1895
2 63231 1 1895
2 63232 1 1895
2 63233 1 1896
2 63234 1 1896
2 63235 1 1897
2 63236 1 1897
2 63237 1 1904
2 63238 1 1904
2 63239 1 1904
2 63240 1 1904
2 63241 1 1906
2 63242 1 1906
2 63243 1 1906
2 63244 1 1906
2 63245 1 1906
2 63246 1 1906
2 63247 1 1906
2 63248 1 1906
2 63249 1 1906
2 63250 1 1906
2 63251 1 1906
2 63252 1 1906
2 63253 1 1906
2 63254 1 1906
2 63255 1 1907
2 63256 1 1907
2 63257 1 1907
2 63258 1 1908
2 63259 1 1908
2 63260 1 1908
2 63261 1 1908
2 63262 1 1927
2 63263 1 1927
2 63264 1 1927
2 63265 1 1929
2 63266 1 1929
2 63267 1 1929
2 63268 1 1929
2 63269 1 1929
2 63270 1 1930
2 63271 1 1930
2 63272 1 1930
2 63273 1 1931
2 63274 1 1931
2 63275 1 1932
2 63276 1 1932
2 63277 1 1933
2 63278 1 1933
2 63279 1 1933
2 63280 1 1933
2 63281 1 1933
2 63282 1 1933
2 63283 1 1933
2 63284 1 1933
2 63285 1 1933
2 63286 1 1933
2 63287 1 1933
2 63288 1 1933
2 63289 1 1933
2 63290 1 1933
2 63291 1 1935
2 63292 1 1935
2 63293 1 1935
2 63294 1 1939
2 63295 1 1939
2 63296 1 1939
2 63297 1 1939
2 63298 1 1940
2 63299 1 1940
2 63300 1 1940
2 63301 1 1940
2 63302 1 1940
2 63303 1 1940
2 63304 1 1940
2 63305 1 1940
2 63306 1 1940
2 63307 1 1940
2 63308 1 1940
2 63309 1 1940
2 63310 1 1940
2 63311 1 1940
2 63312 1 1940
2 63313 1 1940
2 63314 1 1940
2 63315 1 1940
2 63316 1 1940
2 63317 1 1940
2 63318 1 1942
2 63319 1 1942
2 63320 1 1944
2 63321 1 1944
2 63322 1 1952
2 63323 1 1952
2 63324 1 1953
2 63325 1 1953
2 63326 1 1953
2 63327 1 1953
2 63328 1 1953
2 63329 1 1954
2 63330 1 1954
2 63331 1 1954
2 63332 1 1955
2 63333 1 1955
2 63334 1 1956
2 63335 1 1956
2 63336 1 1956
2 63337 1 1971
2 63338 1 1971
2 63339 1 1972
2 63340 1 1972
2 63341 1 1972
2 63342 1 1972
2 63343 1 1972
2 63344 1 1972
2 63345 1 1972
2 63346 1 1972
2 63347 1 1972
2 63348 1 1972
2 63349 1 1980
2 63350 1 1980
2 63351 1 1980
2 63352 1 1980
2 63353 1 1982
2 63354 1 1982
2 63355 1 1982
2 63356 1 1989
2 63357 1 1989
2 63358 1 1989
2 63359 1 1989
2 63360 1 1989
2 63361 1 1990
2 63362 1 1990
2 63363 1 2000
2 63364 1 2000
2 63365 1 2000
2 63366 1 2001
2 63367 1 2001
2 63368 1 2001
2 63369 1 2002
2 63370 1 2002
2 63371 1 2003
2 63372 1 2003
2 63373 1 2004
2 63374 1 2004
2 63375 1 2009
2 63376 1 2009
2 63377 1 2009
2 63378 1 2009
2 63379 1 2009
2 63380 1 2010
2 63381 1 2010
2 63382 1 2028
2 63383 1 2028
2 63384 1 2028
2 63385 1 2029
2 63386 1 2029
2 63387 1 2030
2 63388 1 2030
2 63389 1 2030
2 63390 1 2030
2 63391 1 2032
2 63392 1 2032
2 63393 1 2038
2 63394 1 2038
2 63395 1 2040
2 63396 1 2040
2 63397 1 2040
2 63398 1 2049
2 63399 1 2049
2 63400 1 2049
2 63401 1 2049
2 63402 1 2049
2 63403 1 2049
2 63404 1 2049
2 63405 1 2049
2 63406 1 2049
2 63407 1 2049
2 63408 1 2050
2 63409 1 2050
2 63410 1 2050
2 63411 1 2050
2 63412 1 2051
2 63413 1 2051
2 63414 1 2052
2 63415 1 2052
2 63416 1 2059
2 63417 1 2059
2 63418 1 2059
2 63419 1 2059
2 63420 1 2059
2 63421 1 2059
2 63422 1 2059
2 63423 1 2059
2 63424 1 2059
2 63425 1 2059
2 63426 1 2060
2 63427 1 2060
2 63428 1 2060
2 63429 1 2060
2 63430 1 2061
2 63431 1 2061
2 63432 1 2061
2 63433 1 2061
2 63434 1 2061
2 63435 1 2061
2 63436 1 2061
2 63437 1 2061
2 63438 1 2061
2 63439 1 2061
2 63440 1 2061
2 63441 1 2061
2 63442 1 2061
2 63443 1 2061
2 63444 1 2061
2 63445 1 2061
2 63446 1 2061
2 63447 1 2061
2 63448 1 2061
2 63449 1 2061
2 63450 1 2061
2 63451 1 2061
2 63452 1 2061
2 63453 1 2061
2 63454 1 2061
2 63455 1 2061
2 63456 1 2061
2 63457 1 2061
2 63458 1 2061
2 63459 1 2061
2 63460 1 2061
2 63461 1 2061
2 63462 1 2061
2 63463 1 2061
2 63464 1 2062
2 63465 1 2062
2 63466 1 2062
2 63467 1 2062
2 63468 1 2062
2 63469 1 2062
2 63470 1 2062
2 63471 1 2062
2 63472 1 2062
2 63473 1 2062
2 63474 1 2062
2 63475 1 2063
2 63476 1 2063
2 63477 1 2064
2 63478 1 2064
2 63479 1 2064
2 63480 1 2066
2 63481 1 2066
2 63482 1 2066
2 63483 1 2073
2 63484 1 2073
2 63485 1 2073
2 63486 1 2073
2 63487 1 2073
2 63488 1 2073
2 63489 1 2073
2 63490 1 2073
2 63491 1 2073
2 63492 1 2075
2 63493 1 2075
2 63494 1 2075
2 63495 1 2076
2 63496 1 2076
2 63497 1 2076
2 63498 1 2077
2 63499 1 2077
2 63500 1 2077
2 63501 1 2084
2 63502 1 2084
2 63503 1 2084
2 63504 1 2084
2 63505 1 2084
2 63506 1 2084
2 63507 1 2084
2 63508 1 2084
2 63509 1 2084
2 63510 1 2084
2 63511 1 2084
2 63512 1 2084
2 63513 1 2084
2 63514 1 2084
2 63515 1 2084
2 63516 1 2084
2 63517 1 2084
2 63518 1 2084
2 63519 1 2084
2 63520 1 2084
2 63521 1 2084
2 63522 1 2084
2 63523 1 2084
2 63524 1 2084
2 63525 1 2084
2 63526 1 2084
2 63527 1 2084
2 63528 1 2084
2 63529 1 2084
2 63530 1 2084
2 63531 1 2084
2 63532 1 2084
2 63533 1 2084
2 63534 1 2084
2 63535 1 2084
2 63536 1 2084
2 63537 1 2084
2 63538 1 2084
2 63539 1 2084
2 63540 1 2084
2 63541 1 2084
2 63542 1 2085
2 63543 1 2085
2 63544 1 2085
2 63545 1 2085
2 63546 1 2085
2 63547 1 2085
2 63548 1 2085
2 63549 1 2085
2 63550 1 2085
2 63551 1 2085
2 63552 1 2085
2 63553 1 2086
2 63554 1 2086
2 63555 1 2086
2 63556 1 2086
2 63557 1 2086
2 63558 1 2086
2 63559 1 2086
2 63560 1 2086
2 63561 1 2087
2 63562 1 2087
2 63563 1 2087
2 63564 1 2090
2 63565 1 2090
2 63566 1 2090
2 63567 1 2090
2 63568 1 2090
2 63569 1 2090
2 63570 1 2090
2 63571 1 2090
2 63572 1 2090
2 63573 1 2090
2 63574 1 2090
2 63575 1 2090
2 63576 1 2090
2 63577 1 2092
2 63578 1 2092
2 63579 1 2092
2 63580 1 2092
2 63581 1 2092
2 63582 1 2092
2 63583 1 2092
2 63584 1 2094
2 63585 1 2094
2 63586 1 2094
2 63587 1 2094
2 63588 1 2094
2 63589 1 2096
2 63590 1 2096
2 63591 1 2096
2 63592 1 2108
2 63593 1 2108
2 63594 1 2108
2 63595 1 2108
2 63596 1 2108
2 63597 1 2108
2 63598 1 2108
2 63599 1 2108
2 63600 1 2117
2 63601 1 2117
2 63602 1 2117
2 63603 1 2117
2 63604 1 2117
2 63605 1 2117
2 63606 1 2117
2 63607 1 2117
2 63608 1 2117
2 63609 1 2117
2 63610 1 2117
2 63611 1 2117
2 63612 1 2117
2 63613 1 2117
2 63614 1 2117
2 63615 1 2117
2 63616 1 2117
2 63617 1 2117
2 63618 1 2117
2 63619 1 2117
2 63620 1 2117
2 63621 1 2117
2 63622 1 2118
2 63623 1 2118
2 63624 1 2118
2 63625 1 2118
2 63626 1 2118
2 63627 1 2118
2 63628 1 2118
2 63629 1 2118
2 63630 1 2118
2 63631 1 2118
2 63632 1 2118
2 63633 1 2118
2 63634 1 2119
2 63635 1 2119
2 63636 1 2119
2 63637 1 2119
2 63638 1 2119
2 63639 1 2119
2 63640 1 2119
2 63641 1 2119
2 63642 1 2119
2 63643 1 2119
2 63644 1 2119
2 63645 1 2119
2 63646 1 2119
2 63647 1 2119
2 63648 1 2119
2 63649 1 2122
2 63650 1 2122
2 63651 1 2122
2 63652 1 2123
2 63653 1 2123
2 63654 1 2123
2 63655 1 2123
2 63656 1 2123
2 63657 1 2123
2 63658 1 2123
2 63659 1 2123
2 63660 1 2123
2 63661 1 2123
2 63662 1 2123
2 63663 1 2123
2 63664 1 2123
2 63665 1 2123
2 63666 1 2123
2 63667 1 2123
2 63668 1 2124
2 63669 1 2124
2 63670 1 2124
2 63671 1 2125
2 63672 1 2125
2 63673 1 2125
2 63674 1 2125
2 63675 1 2125
2 63676 1 2125
2 63677 1 2125
2 63678 1 2126
2 63679 1 2126
2 63680 1 2126
2 63681 1 2127
2 63682 1 2127
2 63683 1 2127
2 63684 1 2127
2 63685 1 2128
2 63686 1 2128
2 63687 1 2128
2 63688 1 2130
2 63689 1 2130
2 63690 1 2130
2 63691 1 2141
2 63692 1 2141
2 63693 1 2141
2 63694 1 2141
2 63695 1 2141
2 63696 1 2141
2 63697 1 2142
2 63698 1 2142
2 63699 1 2149
2 63700 1 2149
2 63701 1 2149
2 63702 1 2149
2 63703 1 2149
2 63704 1 2149
2 63705 1 2149
2 63706 1 2149
2 63707 1 2152
2 63708 1 2152
2 63709 1 2157
2 63710 1 2157
2 63711 1 2158
2 63712 1 2158
2 63713 1 2158
2 63714 1 2182
2 63715 1 2182
2 63716 1 2182
2 63717 1 2182
2 63718 1 2182
2 63719 1 2182
2 63720 1 2182
2 63721 1 2182
2 63722 1 2182
2 63723 1 2182
2 63724 1 2182
2 63725 1 2182
2 63726 1 2182
2 63727 1 2182
2 63728 1 2182
2 63729 1 2182
2 63730 1 2182
2 63731 1 2182
2 63732 1 2182
2 63733 1 2182
2 63734 1 2182
2 63735 1 2182
2 63736 1 2182
2 63737 1 2182
2 63738 1 2182
2 63739 1 2182
2 63740 1 2182
2 63741 1 2182
2 63742 1 2182
2 63743 1 2182
2 63744 1 2182
2 63745 1 2182
2 63746 1 2182
2 63747 1 2183
2 63748 1 2183
2 63749 1 2183
2 63750 1 2183
2 63751 1 2183
2 63752 1 2183
2 63753 1 2184
2 63754 1 2184
2 63755 1 2185
2 63756 1 2185
2 63757 1 2185
2 63758 1 2185
2 63759 1 2185
2 63760 1 2185
2 63761 1 2185
2 63762 1 2185
2 63763 1 2185
2 63764 1 2185
2 63765 1 2185
2 63766 1 2185
2 63767 1 2186
2 63768 1 2186
2 63769 1 2186
2 63770 1 2186
2 63771 1 2186
2 63772 1 2186
2 63773 1 2187
2 63774 1 2187
2 63775 1 2187
2 63776 1 2197
2 63777 1 2197
2 63778 1 2197
2 63779 1 2197
2 63780 1 2197
2 63781 1 2197
2 63782 1 2197
2 63783 1 2197
2 63784 1 2197
2 63785 1 2197
2 63786 1 2197
2 63787 1 2197
2 63788 1 2197
2 63789 1 2197
2 63790 1 2197
2 63791 1 2197
2 63792 1 2197
2 63793 1 2197
2 63794 1 2198
2 63795 1 2198
2 63796 1 2198
2 63797 1 2198
2 63798 1 2198
2 63799 1 2199
2 63800 1 2199
2 63801 1 2199
2 63802 1 2199
2 63803 1 2200
2 63804 1 2200
2 63805 1 2200
2 63806 1 2200
2 63807 1 2200
2 63808 1 2200
2 63809 1 2200
2 63810 1 2200
2 63811 1 2207
2 63812 1 2207
2 63813 1 2207
2 63814 1 2207
2 63815 1 2207
2 63816 1 2207
2 63817 1 2207
2 63818 1 2207
2 63819 1 2207
2 63820 1 2207
2 63821 1 2207
2 63822 1 2207
2 63823 1 2207
2 63824 1 2207
2 63825 1 2207
2 63826 1 2207
2 63827 1 2207
2 63828 1 2207
2 63829 1 2207
2 63830 1 2207
2 63831 1 2207
2 63832 1 2207
2 63833 1 2207
2 63834 1 2207
2 63835 1 2207
2 63836 1 2207
2 63837 1 2207
2 63838 1 2207
2 63839 1 2207
2 63840 1 2207
2 63841 1 2207
2 63842 1 2207
2 63843 1 2207
2 63844 1 2207
2 63845 1 2208
2 63846 1 2208
2 63847 1 2208
2 63848 1 2208
2 63849 1 2208
2 63850 1 2208
2 63851 1 2209
2 63852 1 2209
2 63853 1 2209
2 63854 1 2216
2 63855 1 2216
2 63856 1 2216
2 63857 1 2216
2 63858 1 2216
2 63859 1 2227
2 63860 1 2227
2 63861 1 2227
2 63862 1 2227
2 63863 1 2227
2 63864 1 2227
2 63865 1 2232
2 63866 1 2232
2 63867 1 2232
2 63868 1 2233
2 63869 1 2233
2 63870 1 2238
2 63871 1 2238
2 63872 1 2238
2 63873 1 2241
2 63874 1 2241
2 63875 1 2241
2 63876 1 2241
2 63877 1 2241
2 63878 1 2241
2 63879 1 2243
2 63880 1 2243
2 63881 1 2244
2 63882 1 2244
2 63883 1 2244
2 63884 1 2244
2 63885 1 2244
2 63886 1 2244
2 63887 1 2244
2 63888 1 2244
2 63889 1 2244
2 63890 1 2244
2 63891 1 2244
2 63892 1 2245
2 63893 1 2245
2 63894 1 2245
2 63895 1 2247
2 63896 1 2247
2 63897 1 2248
2 63898 1 2248
2 63899 1 2257
2 63900 1 2257
2 63901 1 2260
2 63902 1 2260
2 63903 1 2260
2 63904 1 2269
2 63905 1 2269
2 63906 1 2269
2 63907 1 2270
2 63908 1 2270
2 63909 1 2270
2 63910 1 2270
2 63911 1 2271
2 63912 1 2271
2 63913 1 2272
2 63914 1 2272
2 63915 1 2272
2 63916 1 2272
2 63917 1 2272
2 63918 1 2272
2 63919 1 2274
2 63920 1 2274
2 63921 1 2274
2 63922 1 2275
2 63923 1 2275
2 63924 1 2276
2 63925 1 2276
2 63926 1 2276
2 63927 1 2290
2 63928 1 2290
2 63929 1 2290
2 63930 1 2290
2 63931 1 2291
2 63932 1 2291
2 63933 1 2291
2 63934 1 2291
2 63935 1 2291
2 63936 1 2291
2 63937 1 2291
2 63938 1 2291
2 63939 1 2291
2 63940 1 2291
2 63941 1 2291
2 63942 1 2291
2 63943 1 2291
2 63944 1 2291
2 63945 1 2291
2 63946 1 2291
2 63947 1 2291
2 63948 1 2291
2 63949 1 2291
2 63950 1 2291
2 63951 1 2298
2 63952 1 2298
2 63953 1 2298
2 63954 1 2298
2 63955 1 2298
2 63956 1 2299
2 63957 1 2299
2 63958 1 2299
2 63959 1 2301
2 63960 1 2301
2 63961 1 2301
2 63962 1 2306
2 63963 1 2306
2 63964 1 2306
2 63965 1 2306
2 63966 1 2306
2 63967 1 2306
2 63968 1 2306
2 63969 1 2306
2 63970 1 2306
2 63971 1 2307
2 63972 1 2307
2 63973 1 2307
2 63974 1 2307
2 63975 1 2307
2 63976 1 2308
2 63977 1 2308
2 63978 1 2308
2 63979 1 2308
2 63980 1 2308
2 63981 1 2308
2 63982 1 2308
2 63983 1 2308
2 63984 1 2308
2 63985 1 2308
2 63986 1 2309
2 63987 1 2309
2 63988 1 2309
2 63989 1 2309
2 63990 1 2314
2 63991 1 2314
2 63992 1 2314
2 63993 1 2314
2 63994 1 2314
2 63995 1 2314
2 63996 1 2314
2 63997 1 2314
2 63998 1 2314
2 63999 1 2314
2 64000 1 2314
2 64001 1 2314
2 64002 1 2314
2 64003 1 2314
2 64004 1 2314
2 64005 1 2314
2 64006 1 2314
2 64007 1 2314
2 64008 1 2314
2 64009 1 2314
2 64010 1 2314
2 64011 1 2314
2 64012 1 2315
2 64013 1 2315
2 64014 1 2315
2 64015 1 2315
2 64016 1 2315
2 64017 1 2315
2 64018 1 2315
2 64019 1 2315
2 64020 1 2315
2 64021 1 2315
2 64022 1 2316
2 64023 1 2316
2 64024 1 2316
2 64025 1 2317
2 64026 1 2317
2 64027 1 2317
2 64028 1 2317
2 64029 1 2319
2 64030 1 2319
2 64031 1 2319
2 64032 1 2331
2 64033 1 2331
2 64034 1 2331
2 64035 1 2331
2 64036 1 2332
2 64037 1 2332
2 64038 1 2333
2 64039 1 2333
2 64040 1 2335
2 64041 1 2335
2 64042 1 2336
2 64043 1 2336
2 64044 1 2341
2 64045 1 2341
2 64046 1 2342
2 64047 1 2342
2 64048 1 2342
2 64049 1 2342
2 64050 1 2342
2 64051 1 2342
2 64052 1 2342
2 64053 1 2342
2 64054 1 2344
2 64055 1 2344
2 64056 1 2344
2 64057 1 2345
2 64058 1 2345
2 64059 1 2346
2 64060 1 2346
2 64061 1 2346
2 64062 1 2346
2 64063 1 2346
2 64064 1 2355
2 64065 1 2355
2 64066 1 2356
2 64067 1 2356
2 64068 1 2363
2 64069 1 2363
2 64070 1 2363
2 64071 1 2363
2 64072 1 2363
2 64073 1 2363
2 64074 1 2363
2 64075 1 2363
2 64076 1 2363
2 64077 1 2363
2 64078 1 2364
2 64079 1 2364
2 64080 1 2364
2 64081 1 2365
2 64082 1 2365
2 64083 1 2368
2 64084 1 2368
2 64085 1 2368
2 64086 1 2368
2 64087 1 2376
2 64088 1 2376
2 64089 1 2376
2 64090 1 2386
2 64091 1 2386
2 64092 1 2388
2 64093 1 2388
2 64094 1 2388
2 64095 1 2405
2 64096 1 2405
2 64097 1 2406
2 64098 1 2406
2 64099 1 2406
2 64100 1 2406
2 64101 1 2406
2 64102 1 2410
2 64103 1 2410
2 64104 1 2411
2 64105 1 2411
2 64106 1 2411
2 64107 1 2411
2 64108 1 2412
2 64109 1 2412
2 64110 1 2414
2 64111 1 2414
2 64112 1 2421
2 64113 1 2421
2 64114 1 2421
2 64115 1 2421
2 64116 1 2434
2 64117 1 2434
2 64118 1 2434
2 64119 1 2434
2 64120 1 2434
2 64121 1 2434
2 64122 1 2434
2 64123 1 2434
2 64124 1 2434
2 64125 1 2434
2 64126 1 2434
2 64127 1 2435
2 64128 1 2435
2 64129 1 2435
2 64130 1 2435
2 64131 1 2435
2 64132 1 2435
2 64133 1 2435
2 64134 1 2435
2 64135 1 2435
2 64136 1 2435
2 64137 1 2435
2 64138 1 2435
2 64139 1 2435
2 64140 1 2435
2 64141 1 2435
2 64142 1 2435
2 64143 1 2435
2 64144 1 2435
2 64145 1 2435
2 64146 1 2435
2 64147 1 2435
2 64148 1 2435
2 64149 1 2435
2 64150 1 2435
2 64151 1 2435
2 64152 1 2435
2 64153 1 2436
2 64154 1 2436
2 64155 1 2436
2 64156 1 2436
2 64157 1 2436
2 64158 1 2436
2 64159 1 2437
2 64160 1 2437
2 64161 1 2437
2 64162 1 2437
2 64163 1 2439
2 64164 1 2439
2 64165 1 2439
2 64166 1 2440
2 64167 1 2440
2 64168 1 2445
2 64169 1 2445
2 64170 1 2445
2 64171 1 2445
2 64172 1 2445
2 64173 1 2445
2 64174 1 2445
2 64175 1 2445
2 64176 1 2445
2 64177 1 2445
2 64178 1 2445
2 64179 1 2453
2 64180 1 2453
2 64181 1 2453
2 64182 1 2461
2 64183 1 2461
2 64184 1 2462
2 64185 1 2462
2 64186 1 2462
2 64187 1 2462
2 64188 1 2471
2 64189 1 2471
2 64190 1 2471
2 64191 1 2471
2 64192 1 2471
2 64193 1 2471
2 64194 1 2471
2 64195 1 2471
2 64196 1 2471
2 64197 1 2471
2 64198 1 2471
2 64199 1 2471
2 64200 1 2471
2 64201 1 2471
2 64202 1 2471
2 64203 1 2471
2 64204 1 2472
2 64205 1 2472
2 64206 1 2473
2 64207 1 2473
2 64208 1 2473
2 64209 1 2473
2 64210 1 2473
2 64211 1 2474
2 64212 1 2474
2 64213 1 2474
2 64214 1 2474
2 64215 1 2474
2 64216 1 2474
2 64217 1 2474
2 64218 1 2474
2 64219 1 2474
2 64220 1 2474
2 64221 1 2474
2 64222 1 2474
2 64223 1 2474
2 64224 1 2474
2 64225 1 2475
2 64226 1 2475
2 64227 1 2476
2 64228 1 2476
2 64229 1 2476
2 64230 1 2487
2 64231 1 2487
2 64232 1 2487
2 64233 1 2487
2 64234 1 2487
2 64235 1 2487
2 64236 1 2487
2 64237 1 2487
2 64238 1 2487
2 64239 1 2487
2 64240 1 2487
2 64241 1 2487
2 64242 1 2487
2 64243 1 2487
2 64244 1 2489
2 64245 1 2489
2 64246 1 2489
2 64247 1 2489
2 64248 1 2491
2 64249 1 2491
2 64250 1 2498
2 64251 1 2498
2 64252 1 2498
2 64253 1 2499
2 64254 1 2499
2 64255 1 2499
2 64256 1 2499
2 64257 1 2499
2 64258 1 2507
2 64259 1 2507
2 64260 1 2507
2 64261 1 2507
2 64262 1 2508
2 64263 1 2508
2 64264 1 2518
2 64265 1 2518
2 64266 1 2518
2 64267 1 2518
2 64268 1 2518
2 64269 1 2518
2 64270 1 2518
2 64271 1 2518
2 64272 1 2520
2 64273 1 2520
2 64274 1 2520
2 64275 1 2520
2 64276 1 2520
2 64277 1 2520
2 64278 1 2520
2 64279 1 2520
2 64280 1 2521
2 64281 1 2521
2 64282 1 2521
2 64283 1 2522
2 64284 1 2522
2 64285 1 2522
2 64286 1 2522
2 64287 1 2522
2 64288 1 2522
2 64289 1 2522
2 64290 1 2522
2 64291 1 2522
2 64292 1 2522
2 64293 1 2522
2 64294 1 2522
2 64295 1 2523
2 64296 1 2523
2 64297 1 2523
2 64298 1 2523
2 64299 1 2525
2 64300 1 2525
2 64301 1 2525
2 64302 1 2532
2 64303 1 2532
2 64304 1 2533
2 64305 1 2533
2 64306 1 2533
2 64307 1 2533
2 64308 1 2534
2 64309 1 2534
2 64310 1 2541
2 64311 1 2541
2 64312 1 2541
2 64313 1 2541
2 64314 1 2543
2 64315 1 2543
2 64316 1 2543
2 64317 1 2543
2 64318 1 2543
2 64319 1 2543
2 64320 1 2543
2 64321 1 2545
2 64322 1 2545
2 64323 1 2545
2 64324 1 2545
2 64325 1 2545
2 64326 1 2545
2 64327 1 2545
2 64328 1 2545
2 64329 1 2545
2 64330 1 2545
2 64331 1 2545
2 64332 1 2545
2 64333 1 2545
2 64334 1 2545
2 64335 1 2545
2 64336 1 2545
2 64337 1 2547
2 64338 1 2547
2 64339 1 2547
2 64340 1 2549
2 64341 1 2549
2 64342 1 2549
2 64343 1 2555
2 64344 1 2555
2 64345 1 2555
2 64346 1 2555
2 64347 1 2555
2 64348 1 2555
2 64349 1 2555
2 64350 1 2555
2 64351 1 2555
2 64352 1 2555
2 64353 1 2555
2 64354 1 2556
2 64355 1 2556
2 64356 1 2556
2 64357 1 2556
2 64358 1 2563
2 64359 1 2563
2 64360 1 2565
2 64361 1 2565
2 64362 1 2567
2 64363 1 2567
2 64364 1 2567
2 64365 1 2567
2 64366 1 2567
2 64367 1 2567
2 64368 1 2576
2 64369 1 2576
2 64370 1 2576
2 64371 1 2576
2 64372 1 2576
2 64373 1 2576
2 64374 1 2576
2 64375 1 2577
2 64376 1 2577
2 64377 1 2577
2 64378 1 2577
2 64379 1 2577
2 64380 1 2577
2 64381 1 2577
2 64382 1 2577
2 64383 1 2577
2 64384 1 2577
2 64385 1 2577
2 64386 1 2577
2 64387 1 2577
2 64388 1 2577
2 64389 1 2577
2 64390 1 2577
2 64391 1 2577
2 64392 1 2578
2 64393 1 2578
2 64394 1 2581
2 64395 1 2581
2 64396 1 2581
2 64397 1 2583
2 64398 1 2583
2 64399 1 2586
2 64400 1 2586
2 64401 1 2588
2 64402 1 2588
2 64403 1 2589
2 64404 1 2589
2 64405 1 2599
2 64406 1 2599
2 64407 1 2599
2 64408 1 2599
2 64409 1 2599
2 64410 1 2599
2 64411 1 2600
2 64412 1 2600
2 64413 1 2602
2 64414 1 2602
2 64415 1 2602
2 64416 1 2602
2 64417 1 2602
2 64418 1 2602
2 64419 1 2602
2 64420 1 2604
2 64421 1 2604
2 64422 1 2613
2 64423 1 2613
2 64424 1 2613
2 64425 1 2617
2 64426 1 2617
2 64427 1 2619
2 64428 1 2619
2 64429 1 2621
2 64430 1 2621
2 64431 1 2621
2 64432 1 2621
2 64433 1 2621
2 64434 1 2622
2 64435 1 2622
2 64436 1 2622
2 64437 1 2622
2 64438 1 2622
2 64439 1 2622
2 64440 1 2623
2 64441 1 2623
2 64442 1 2634
2 64443 1 2634
2 64444 1 2634
2 64445 1 2634
2 64446 1 2634
2 64447 1 2634
2 64448 1 2634
2 64449 1 2634
2 64450 1 2634
2 64451 1 2634
2 64452 1 2634
2 64453 1 2634
2 64454 1 2634
2 64455 1 2634
2 64456 1 2635
2 64457 1 2635
2 64458 1 2635
2 64459 1 2647
2 64460 1 2647
2 64461 1 2647
2 64462 1 2647
2 64463 1 2647
2 64464 1 2647
2 64465 1 2647
2 64466 1 2647
2 64467 1 2648
2 64468 1 2648
2 64469 1 2648
2 64470 1 2648
2 64471 1 2648
2 64472 1 2648
2 64473 1 2648
2 64474 1 2648
2 64475 1 2648
2 64476 1 2649
2 64477 1 2649
2 64478 1 2649
2 64479 1 2649
2 64480 1 2649
2 64481 1 2649
2 64482 1 2649
2 64483 1 2658
2 64484 1 2658
2 64485 1 2659
2 64486 1 2659
2 64487 1 2659
2 64488 1 2659
2 64489 1 2659
2 64490 1 2659
2 64491 1 2661
2 64492 1 2661
2 64493 1 2661
2 64494 1 2661
2 64495 1 2662
2 64496 1 2662
2 64497 1 2671
2 64498 1 2671
2 64499 1 2671
2 64500 1 2671
2 64501 1 2671
2 64502 1 2671
2 64503 1 2671
2 64504 1 2671
2 64505 1 2671
2 64506 1 2671
2 64507 1 2671
2 64508 1 2671
2 64509 1 2671
2 64510 1 2671
2 64511 1 2671
2 64512 1 2671
2 64513 1 2672
2 64514 1 2672
2 64515 1 2681
2 64516 1 2681
2 64517 1 2681
2 64518 1 2681
2 64519 1 2681
2 64520 1 2681
2 64521 1 2682
2 64522 1 2682
2 64523 1 2682
2 64524 1 2682
2 64525 1 2702
2 64526 1 2702
2 64527 1 2703
2 64528 1 2703
2 64529 1 2725
2 64530 1 2725
2 64531 1 2725
2 64532 1 2738
2 64533 1 2738
2 64534 1 2746
2 64535 1 2746
2 64536 1 2746
2 64537 1 2746
2 64538 1 2746
2 64539 1 2746
2 64540 1 2746
2 64541 1 2746
2 64542 1 2746
2 64543 1 2747
2 64544 1 2747
2 64545 1 2747
2 64546 1 2748
2 64547 1 2748
2 64548 1 2749
2 64549 1 2749
2 64550 1 2749
2 64551 1 2749
2 64552 1 2757
2 64553 1 2757
2 64554 1 2757
2 64555 1 2762
2 64556 1 2762
2 64557 1 2765
2 64558 1 2765
2 64559 1 2765
2 64560 1 2765
2 64561 1 2766
2 64562 1 2766
2 64563 1 2766
2 64564 1 2766
2 64565 1 2766
2 64566 1 2766
2 64567 1 2767
2 64568 1 2767
2 64569 1 2767
2 64570 1 2767
2 64571 1 2767
2 64572 1 2767
2 64573 1 2767
2 64574 1 2767
2 64575 1 2767
2 64576 1 2767
2 64577 1 2768
2 64578 1 2768
2 64579 1 2768
2 64580 1 2768
2 64581 1 2782
2 64582 1 2782
2 64583 1 2782
2 64584 1 2782
2 64585 1 2782
2 64586 1 2782
2 64587 1 2782
2 64588 1 2782
2 64589 1 2782
2 64590 1 2782
2 64591 1 2782
2 64592 1 2782
2 64593 1 2782
2 64594 1 2782
2 64595 1 2782
2 64596 1 2782
2 64597 1 2782
2 64598 1 2782
2 64599 1 2782
2 64600 1 2782
2 64601 1 2783
2 64602 1 2783
2 64603 1 2783
2 64604 1 2783
2 64605 1 2783
2 64606 1 2783
2 64607 1 2783
2 64608 1 2783
2 64609 1 2784
2 64610 1 2784
2 64611 1 2784
2 64612 1 2786
2 64613 1 2786
2 64614 1 2786
2 64615 1 2786
2 64616 1 2786
2 64617 1 2789
2 64618 1 2789
2 64619 1 2789
2 64620 1 2789
2 64621 1 2789
2 64622 1 2789
2 64623 1 2803
2 64624 1 2803
2 64625 1 2803
2 64626 1 2803
2 64627 1 2803
2 64628 1 2803
2 64629 1 2810
2 64630 1 2810
2 64631 1 2815
2 64632 1 2815
2 64633 1 2818
2 64634 1 2818
2 64635 1 2818
2 64636 1 2818
2 64637 1 2818
2 64638 1 2818
2 64639 1 2818
2 64640 1 2818
2 64641 1 2818
2 64642 1 2818
2 64643 1 2818
2 64644 1 2818
2 64645 1 2818
2 64646 1 2820
2 64647 1 2820
2 64648 1 2826
2 64649 1 2826
2 64650 1 2826
2 64651 1 2826
2 64652 1 2826
2 64653 1 2826
2 64654 1 2826
2 64655 1 2826
2 64656 1 2826
2 64657 1 2826
2 64658 1 2826
2 64659 1 2844
2 64660 1 2844
2 64661 1 2844
2 64662 1 2844
2 64663 1 2844
2 64664 1 2844
2 64665 1 2845
2 64666 1 2845
2 64667 1 2845
2 64668 1 2845
2 64669 1 2845
2 64670 1 2845
2 64671 1 2847
2 64672 1 2847
2 64673 1 2855
2 64674 1 2855
2 64675 1 2863
2 64676 1 2863
2 64677 1 2865
2 64678 1 2865
2 64679 1 2865
2 64680 1 2865
2 64681 1 2875
2 64682 1 2875
2 64683 1 2875
2 64684 1 2875
2 64685 1 2876
2 64686 1 2876
2 64687 1 2876
2 64688 1 2876
2 64689 1 2877
2 64690 1 2877
2 64691 1 2889
2 64692 1 2889
2 64693 1 2889
2 64694 1 2889
2 64695 1 2895
2 64696 1 2895
2 64697 1 2895
2 64698 1 2895
2 64699 1 2895
2 64700 1 2895
2 64701 1 2895
2 64702 1 2895
2 64703 1 2895
2 64704 1 2895
2 64705 1 2895
2 64706 1 2895
2 64707 1 2895
2 64708 1 2895
2 64709 1 2895
2 64710 1 2895
2 64711 1 2895
2 64712 1 2895
2 64713 1 2895
2 64714 1 2896
2 64715 1 2896
2 64716 1 2897
2 64717 1 2897
2 64718 1 2897
2 64719 1 2898
2 64720 1 2898
2 64721 1 2917
2 64722 1 2917
2 64723 1 2917
2 64724 1 2917
2 64725 1 2918
2 64726 1 2918
2 64727 1 2918
2 64728 1 2919
2 64729 1 2919
2 64730 1 2919
2 64731 1 2920
2 64732 1 2920
2 64733 1 2920
2 64734 1 2927
2 64735 1 2927
2 64736 1 2927
2 64737 1 2927
2 64738 1 2927
2 64739 1 2927
2 64740 1 2927
2 64741 1 2927
2 64742 1 2928
2 64743 1 2928
2 64744 1 2933
2 64745 1 2933
2 64746 1 2933
2 64747 1 2934
2 64748 1 2934
2 64749 1 2934
2 64750 1 2934
2 64751 1 2937
2 64752 1 2937
2 64753 1 2937
2 64754 1 2937
2 64755 1 2937
2 64756 1 2937
2 64757 1 2937
2 64758 1 2937
2 64759 1 2937
2 64760 1 2937
2 64761 1 2958
2 64762 1 2958
2 64763 1 2958
2 64764 1 2958
2 64765 1 2958
2 64766 1 2959
2 64767 1 2959
2 64768 1 2959
2 64769 1 2959
2 64770 1 2959
2 64771 1 2959
2 64772 1 2966
2 64773 1 2966
2 64774 1 2969
2 64775 1 2969
2 64776 1 2969
2 64777 1 2978
2 64778 1 2978
2 64779 1 2978
2 64780 1 2978
2 64781 1 2978
2 64782 1 2978
2 64783 1 2978
2 64784 1 2978
2 64785 1 2978
2 64786 1 2978
2 64787 1 2978
2 64788 1 2978
2 64789 1 2978
2 64790 1 2978
2 64791 1 2978
2 64792 1 2978
2 64793 1 2979
2 64794 1 2979
2 64795 1 2980
2 64796 1 2980
2 64797 1 2980
2 64798 1 2985
2 64799 1 2985
2 64800 1 2986
2 64801 1 2986
2 64802 1 2986
2 64803 1 2986
2 64804 1 2986
2 64805 1 2986
2 64806 1 2986
2 64807 1 2986
2 64808 1 2986
2 64809 1 2986
2 64810 1 2986
2 64811 1 2986
2 64812 1 2986
2 64813 1 2986
2 64814 1 2986
2 64815 1 2999
2 64816 1 2999
2 64817 1 2999
2 64818 1 2999
2 64819 1 2999
2 64820 1 2999
2 64821 1 2999
2 64822 1 2999
2 64823 1 3000
2 64824 1 3000
2 64825 1 3000
2 64826 1 3000
2 64827 1 3000
2 64828 1 3001
2 64829 1 3001
2 64830 1 3001
2 64831 1 3001
2 64832 1 3009
2 64833 1 3009
2 64834 1 3010
2 64835 1 3010
2 64836 1 3010
2 64837 1 3011
2 64838 1 3011
2 64839 1 3013
2 64840 1 3013
2 64841 1 3013
2 64842 1 3014
2 64843 1 3014
2 64844 1 3016
2 64845 1 3016
2 64846 1 3016
2 64847 1 3017
2 64848 1 3017
2 64849 1 3018
2 64850 1 3018
2 64851 1 3018
2 64852 1 3019
2 64853 1 3019
2 64854 1 3020
2 64855 1 3020
2 64856 1 3020
2 64857 1 3020
2 64858 1 3020
2 64859 1 3032
2 64860 1 3032
2 64861 1 3032
2 64862 1 3032
2 64863 1 3032
2 64864 1 3059
2 64865 1 3059
2 64866 1 3059
2 64867 1 3059
2 64868 1 3059
2 64869 1 3059
2 64870 1 3059
2 64871 1 3059
2 64872 1 3059
2 64873 1 3059
2 64874 1 3059
2 64875 1 3060
2 64876 1 3060
2 64877 1 3060
2 64878 1 3061
2 64879 1 3061
2 64880 1 3061
2 64881 1 3061
2 64882 1 3061
2 64883 1 3061
2 64884 1 3062
2 64885 1 3062
2 64886 1 3062
2 64887 1 3062
2 64888 1 3065
2 64889 1 3065
2 64890 1 3065
2 64891 1 3068
2 64892 1 3068
2 64893 1 3068
2 64894 1 3068
2 64895 1 3068
2 64896 1 3068
2 64897 1 3068
2 64898 1 3080
2 64899 1 3080
2 64900 1 3080
2 64901 1 3080
2 64902 1 3080
2 64903 1 3081
2 64904 1 3081
2 64905 1 3081
2 64906 1 3081
2 64907 1 3081
2 64908 1 3081
2 64909 1 3081
2 64910 1 3082
2 64911 1 3082
2 64912 1 3087
2 64913 1 3087
2 64914 1 3090
2 64915 1 3090
2 64916 1 3090
2 64917 1 3090
2 64918 1 3090
2 64919 1 3090
2 64920 1 3090
2 64921 1 3090
2 64922 1 3090
2 64923 1 3091
2 64924 1 3091
2 64925 1 3091
2 64926 1 3091
2 64927 1 3092
2 64928 1 3092
2 64929 1 3092
2 64930 1 3093
2 64931 1 3093
2 64932 1 3093
2 64933 1 3094
2 64934 1 3094
2 64935 1 3106
2 64936 1 3106
2 64937 1 3106
2 64938 1 3106
2 64939 1 3106
2 64940 1 3107
2 64941 1 3107
2 64942 1 3108
2 64943 1 3108
2 64944 1 3108
2 64945 1 3108
2 64946 1 3108
2 64947 1 3108
2 64948 1 3112
2 64949 1 3112
2 64950 1 3112
2 64951 1 3112
2 64952 1 3113
2 64953 1 3113
2 64954 1 3113
2 64955 1 3113
2 64956 1 3113
2 64957 1 3115
2 64958 1 3115
2 64959 1 3115
2 64960 1 3115
2 64961 1 3118
2 64962 1 3118
2 64963 1 3118
2 64964 1 3118
2 64965 1 3119
2 64966 1 3119
2 64967 1 3119
2 64968 1 3120
2 64969 1 3120
2 64970 1 3120
2 64971 1 3121
2 64972 1 3121
2 64973 1 3121
2 64974 1 3121
2 64975 1 3121
2 64976 1 3121
2 64977 1 3122
2 64978 1 3122
2 64979 1 3133
2 64980 1 3133
2 64981 1 3149
2 64982 1 3149
2 64983 1 3149
2 64984 1 3149
2 64985 1 3149
2 64986 1 3151
2 64987 1 3151
2 64988 1 3151
2 64989 1 3151
2 64990 1 3153
2 64991 1 3153
2 64992 1 3153
2 64993 1 3153
2 64994 1 3157
2 64995 1 3157
2 64996 1 3158
2 64997 1 3158
2 64998 1 3163
2 64999 1 3163
2 65000 1 3163
2 65001 1 3163
2 65002 1 3163
2 65003 1 3163
2 65004 1 3163
2 65005 1 3163
2 65006 1 3163
2 65007 1 3163
2 65008 1 3163
2 65009 1 3163
2 65010 1 3163
2 65011 1 3163
2 65012 1 3163
2 65013 1 3163
2 65014 1 3164
2 65015 1 3164
2 65016 1 3164
2 65017 1 3164
2 65018 1 3164
2 65019 1 3164
2 65020 1 3164
2 65021 1 3165
2 65022 1 3165
2 65023 1 3166
2 65024 1 3166
2 65025 1 3169
2 65026 1 3169
2 65027 1 3169
2 65028 1 3169
2 65029 1 3169
2 65030 1 3169
2 65031 1 3169
2 65032 1 3170
2 65033 1 3170
2 65034 1 3172
2 65035 1 3172
2 65036 1 3179
2 65037 1 3179
2 65038 1 3179
2 65039 1 3180
2 65040 1 3180
2 65041 1 3181
2 65042 1 3181
2 65043 1 3181
2 65044 1 3181
2 65045 1 3181
2 65046 1 3181
2 65047 1 3182
2 65048 1 3182
2 65049 1 3183
2 65050 1 3183
2 65051 1 3183
2 65052 1 3187
2 65053 1 3187
2 65054 1 3187
2 65055 1 3187
2 65056 1 3187
2 65057 1 3187
2 65058 1 3187
2 65059 1 3187
2 65060 1 3187
2 65061 1 3188
2 65062 1 3188
2 65063 1 3189
2 65064 1 3189
2 65065 1 3189
2 65066 1 3189
2 65067 1 3189
2 65068 1 3189
2 65069 1 3189
2 65070 1 3189
2 65071 1 3189
2 65072 1 3189
2 65073 1 3189
2 65074 1 3189
2 65075 1 3189
2 65076 1 3190
2 65077 1 3190
2 65078 1 3190
2 65079 1 3190
2 65080 1 3197
2 65081 1 3197
2 65082 1 3209
2 65083 1 3209
2 65084 1 3210
2 65085 1 3210
2 65086 1 3211
2 65087 1 3211
2 65088 1 3211
2 65089 1 3211
2 65090 1 3215
2 65091 1 3215
2 65092 1 3215
2 65093 1 3218
2 65094 1 3218
2 65095 1 3218
2 65096 1 3218
2 65097 1 3218
2 65098 1 3218
2 65099 1 3218
2 65100 1 3219
2 65101 1 3219
2 65102 1 3220
2 65103 1 3220
2 65104 1 3226
2 65105 1 3226
2 65106 1 3226
2 65107 1 3227
2 65108 1 3227
2 65109 1 3230
2 65110 1 3230
2 65111 1 3230
2 65112 1 3230
2 65113 1 3232
2 65114 1 3232
2 65115 1 3232
2 65116 1 3232
2 65117 1 3232
2 65118 1 3232
2 65119 1 3232
2 65120 1 3232
2 65121 1 3232
2 65122 1 3232
2 65123 1 3232
2 65124 1 3232
2 65125 1 3232
2 65126 1 3232
2 65127 1 3233
2 65128 1 3233
2 65129 1 3233
2 65130 1 3233
2 65131 1 3233
2 65132 1 3247
2 65133 1 3247
2 65134 1 3250
2 65135 1 3250
2 65136 1 3250
2 65137 1 3250
2 65138 1 3250
2 65139 1 3252
2 65140 1 3252
2 65141 1 3256
2 65142 1 3256
2 65143 1 3256
2 65144 1 3257
2 65145 1 3257
2 65146 1 3257
2 65147 1 3257
2 65148 1 3257
2 65149 1 3257
2 65150 1 3257
2 65151 1 3257
2 65152 1 3258
2 65153 1 3258
2 65154 1 3269
2 65155 1 3269
2 65156 1 3276
2 65157 1 3276
2 65158 1 3276
2 65159 1 3276
2 65160 1 3276
2 65161 1 3276
2 65162 1 3276
2 65163 1 3277
2 65164 1 3277
2 65165 1 3277
2 65166 1 3278
2 65167 1 3278
2 65168 1 3278
2 65169 1 3278
2 65170 1 3278
2 65171 1 3278
2 65172 1 3279
2 65173 1 3279
2 65174 1 3279
2 65175 1 3285
2 65176 1 3285
2 65177 1 3287
2 65178 1 3287
2 65179 1 3288
2 65180 1 3288
2 65181 1 3289
2 65182 1 3289
2 65183 1 3289
2 65184 1 3289
2 65185 1 3289
2 65186 1 3289
2 65187 1 3290
2 65188 1 3290
2 65189 1 3290
2 65190 1 3295
2 65191 1 3295
2 65192 1 3296
2 65193 1 3296
2 65194 1 3296
2 65195 1 3306
2 65196 1 3306
2 65197 1 3306
2 65198 1 3307
2 65199 1 3307
2 65200 1 3307
2 65201 1 3307
2 65202 1 3307
2 65203 1 3307
2 65204 1 3307
2 65205 1 3307
2 65206 1 3307
2 65207 1 3307
2 65208 1 3307
2 65209 1 3307
2 65210 1 3307
2 65211 1 3307
2 65212 1 3307
2 65213 1 3309
2 65214 1 3309
2 65215 1 3314
2 65216 1 3314
2 65217 1 3314
2 65218 1 3314
2 65219 1 3314
2 65220 1 3314
2 65221 1 3314
2 65222 1 3314
2 65223 1 3314
2 65224 1 3315
2 65225 1 3315
2 65226 1 3316
2 65227 1 3316
2 65228 1 3316
2 65229 1 3316
2 65230 1 3316
2 65231 1 3316
2 65232 1 3316
2 65233 1 3317
2 65234 1 3317
2 65235 1 3317
2 65236 1 3317
2 65237 1 3317
2 65238 1 3318
2 65239 1 3318
2 65240 1 3322
2 65241 1 3322
2 65242 1 3322
2 65243 1 3322
2 65244 1 3322
2 65245 1 3322
2 65246 1 3322
2 65247 1 3322
2 65248 1 3322
2 65249 1 3322
2 65250 1 3322
2 65251 1 3322
2 65252 1 3322
2 65253 1 3322
2 65254 1 3323
2 65255 1 3323
2 65256 1 3323
2 65257 1 3323
2 65258 1 3323
2 65259 1 3324
2 65260 1 3324
2 65261 1 3324
2 65262 1 3326
2 65263 1 3326
2 65264 1 3326
2 65265 1 3329
2 65266 1 3329
2 65267 1 3332
2 65268 1 3332
2 65269 1 3348
2 65270 1 3348
2 65271 1 3348
2 65272 1 3348
2 65273 1 3348
2 65274 1 3354
2 65275 1 3354
2 65276 1 3354
2 65277 1 3354
2 65278 1 3354
2 65279 1 3354
2 65280 1 3354
2 65281 1 3354
2 65282 1 3365
2 65283 1 3365
2 65284 1 3369
2 65285 1 3369
2 65286 1 3378
2 65287 1 3378
2 65288 1 3378
2 65289 1 3380
2 65290 1 3380
2 65291 1 3380
2 65292 1 3386
2 65293 1 3386
2 65294 1 3386
2 65295 1 3386
2 65296 1 3386
2 65297 1 3386
2 65298 1 3386
2 65299 1 3386
2 65300 1 3387
2 65301 1 3387
2 65302 1 3387
2 65303 1 3389
2 65304 1 3389
2 65305 1 3389
2 65306 1 3392
2 65307 1 3392
2 65308 1 3411
2 65309 1 3411
2 65310 1 3412
2 65311 1 3412
2 65312 1 3415
2 65313 1 3415
2 65314 1 3415
2 65315 1 3415
2 65316 1 3423
2 65317 1 3423
2 65318 1 3423
2 65319 1 3423
2 65320 1 3423
2 65321 1 3423
2 65322 1 3424
2 65323 1 3424
2 65324 1 3428
2 65325 1 3428
2 65326 1 3428
2 65327 1 3438
2 65328 1 3438
2 65329 1 3438
2 65330 1 3438
2 65331 1 3438
2 65332 1 3439
2 65333 1 3439
2 65334 1 3447
2 65335 1 3447
2 65336 1 3447
2 65337 1 3447
2 65338 1 3447
2 65339 1 3447
2 65340 1 3447
2 65341 1 3447
2 65342 1 3447
2 65343 1 3447
2 65344 1 3447
2 65345 1 3447
2 65346 1 3447
2 65347 1 3447
2 65348 1 3448
2 65349 1 3448
2 65350 1 3448
2 65351 1 3448
2 65352 1 3448
2 65353 1 3448
2 65354 1 3448
2 65355 1 3449
2 65356 1 3449
2 65357 1 3449
2 65358 1 3449
2 65359 1 3450
2 65360 1 3450
2 65361 1 3450
2 65362 1 3450
2 65363 1 3450
2 65364 1 3450
2 65365 1 3452
2 65366 1 3452
2 65367 1 3452
2 65368 1 3457
2 65369 1 3457
2 65370 1 3457
2 65371 1 3458
2 65372 1 3458
2 65373 1 3458
2 65374 1 3458
2 65375 1 3458
2 65376 1 3458
2 65377 1 3458
2 65378 1 3458
2 65379 1 3458
2 65380 1 3458
2 65381 1 3459
2 65382 1 3459
2 65383 1 3459
2 65384 1 3460
2 65385 1 3460
2 65386 1 3487
2 65387 1 3487
2 65388 1 3490
2 65389 1 3490
2 65390 1 3490
2 65391 1 3491
2 65392 1 3491
2 65393 1 3492
2 65394 1 3492
2 65395 1 3492
2 65396 1 3493
2 65397 1 3493
2 65398 1 3495
2 65399 1 3495
2 65400 1 3499
2 65401 1 3499
2 65402 1 3499
2 65403 1 3499
2 65404 1 3500
2 65405 1 3500
2 65406 1 3500
2 65407 1 3502
2 65408 1 3502
2 65409 1 3519
2 65410 1 3519
2 65411 1 3520
2 65412 1 3520
2 65413 1 3521
2 65414 1 3521
2 65415 1 3529
2 65416 1 3529
2 65417 1 3529
2 65418 1 3530
2 65419 1 3530
2 65420 1 3530
2 65421 1 3531
2 65422 1 3531
2 65423 1 3539
2 65424 1 3539
2 65425 1 3539
2 65426 1 3539
2 65427 1 3539
2 65428 1 3540
2 65429 1 3540
2 65430 1 3540
2 65431 1 3541
2 65432 1 3541
2 65433 1 3541
2 65434 1 3541
2 65435 1 3543
2 65436 1 3543
2 65437 1 3543
2 65438 1 3543
2 65439 1 3543
2 65440 1 3543
2 65441 1 3545
2 65442 1 3545
2 65443 1 3549
2 65444 1 3549
2 65445 1 3549
2 65446 1 3549
2 65447 1 3549
2 65448 1 3550
2 65449 1 3550
2 65450 1 3550
2 65451 1 3552
2 65452 1 3552
2 65453 1 3552
2 65454 1 3552
2 65455 1 3552
2 65456 1 3560
2 65457 1 3560
2 65458 1 3561
2 65459 1 3561
2 65460 1 3564
2 65461 1 3564
2 65462 1 3565
2 65463 1 3565
2 65464 1 3565
2 65465 1 3565
2 65466 1 3581
2 65467 1 3581
2 65468 1 3581
2 65469 1 3581
2 65470 1 3581
2 65471 1 3583
2 65472 1 3583
2 65473 1 3583
2 65474 1 3583
2 65475 1 3583
2 65476 1 3583
2 65477 1 3583
2 65478 1 3583
2 65479 1 3583
2 65480 1 3583
2 65481 1 3584
2 65482 1 3584
2 65483 1 3585
2 65484 1 3585
2 65485 1 3594
2 65486 1 3594
2 65487 1 3602
2 65488 1 3602
2 65489 1 3604
2 65490 1 3604
2 65491 1 3604
2 65492 1 3604
2 65493 1 3605
2 65494 1 3605
2 65495 1 3605
2 65496 1 3612
2 65497 1 3612
2 65498 1 3613
2 65499 1 3613
2 65500 1 3618
2 65501 1 3618
2 65502 1 3620
2 65503 1 3620
2 65504 1 3641
2 65505 1 3641
2 65506 1 3641
2 65507 1 3641
2 65508 1 3641
2 65509 1 3641
2 65510 1 3656
2 65511 1 3656
2 65512 1 3662
2 65513 1 3662
2 65514 1 3662
2 65515 1 3665
2 65516 1 3665
2 65517 1 3665
2 65518 1 3666
2 65519 1 3666
2 65520 1 3666
2 65521 1 3666
2 65522 1 3666
2 65523 1 3666
2 65524 1 3666
2 65525 1 3676
2 65526 1 3676
2 65527 1 3676
2 65528 1 3676
2 65529 1 3676
2 65530 1 3676
2 65531 1 3676
2 65532 1 3676
2 65533 1 3676
2 65534 1 3677
2 65535 1 3677
2 65536 1 3680
2 65537 1 3680
2 65538 1 3680
2 65539 1 3680
2 65540 1 3680
2 65541 1 3680
2 65542 1 3680
2 65543 1 3680
2 65544 1 3680
2 65545 1 3680
2 65546 1 3680
2 65547 1 3680
2 65548 1 3707
2 65549 1 3707
2 65550 1 3707
2 65551 1 3711
2 65552 1 3711
2 65553 1 3711
2 65554 1 3711
2 65555 1 3712
2 65556 1 3712
2 65557 1 3712
2 65558 1 3751
2 65559 1 3751
2 65560 1 3751
2 65561 1 3751
2 65562 1 3751
2 65563 1 3754
2 65564 1 3754
2 65565 1 3755
2 65566 1 3755
2 65567 1 3782
2 65568 1 3782
2 65569 1 3791
2 65570 1 3791
2 65571 1 3795
2 65572 1 3795
2 65573 1 3795
2 65574 1 3795
2 65575 1 3795
2 65576 1 3796
2 65577 1 3796
2 65578 1 3803
2 65579 1 3803
2 65580 1 3804
2 65581 1 3804
2 65582 1 3805
2 65583 1 3805
2 65584 1 3805
2 65585 1 3805
2 65586 1 3805
2 65587 1 3805
2 65588 1 3805
2 65589 1 3818
2 65590 1 3818
2 65591 1 3822
2 65592 1 3822
2 65593 1 3822
2 65594 1 3822
2 65595 1 3823
2 65596 1 3823
2 65597 1 3823
2 65598 1 3823
2 65599 1 3826
2 65600 1 3826
2 65601 1 3827
2 65602 1 3827
2 65603 1 3828
2 65604 1 3828
2 65605 1 3828
2 65606 1 3829
2 65607 1 3829
2 65608 1 3829
2 65609 1 3841
2 65610 1 3841
2 65611 1 3841
2 65612 1 3841
2 65613 1 3841
2 65614 1 3841
2 65615 1 3858
2 65616 1 3858
2 65617 1 3858
2 65618 1 3858
2 65619 1 3858
2 65620 1 3858
2 65621 1 3858
2 65622 1 3858
2 65623 1 3858
2 65624 1 3858
2 65625 1 3858
2 65626 1 3858
2 65627 1 3858
2 65628 1 3858
2 65629 1 3858
2 65630 1 3858
2 65631 1 3858
2 65632 1 3858
2 65633 1 3860
2 65634 1 3860
2 65635 1 3884
2 65636 1 3884
2 65637 1 3884
2 65638 1 3886
2 65639 1 3886
2 65640 1 3886
2 65641 1 3892
2 65642 1 3892
2 65643 1 3896
2 65644 1 3896
2 65645 1 3925
2 65646 1 3925
2 65647 1 3935
2 65648 1 3935
2 65649 1 3935
2 65650 1 3935
2 65651 1 3936
2 65652 1 3936
2 65653 1 3947
2 65654 1 3947
2 65655 1 3959
2 65656 1 3959
2 65657 1 3990
2 65658 1 3990
2 65659 1 3990
2 65660 1 3990
2 65661 1 4015
2 65662 1 4015
2 65663 1 4015
2 65664 1 4015
2 65665 1 4030
2 65666 1 4030
2 65667 1 4034
2 65668 1 4034
2 65669 1 4034
2 65670 1 4034
2 65671 1 4034
2 65672 1 4034
2 65673 1 4034
2 65674 1 4034
2 65675 1 4035
2 65676 1 4035
2 65677 1 4035
2 65678 1 4035
2 65679 1 4035
2 65680 1 4035
2 65681 1 4035
2 65682 1 4035
2 65683 1 4046
2 65684 1 4046
2 65685 1 4046
2 65686 1 4046
2 65687 1 4061
2 65688 1 4061
2 65689 1 4061
2 65690 1 4061
2 65691 1 4063
2 65692 1 4063
2 65693 1 4093
2 65694 1 4093
2 65695 1 4093
2 65696 1 4093
2 65697 1 4093
2 65698 1 4093
2 65699 1 4093
2 65700 1 4093
2 65701 1 4093
2 65702 1 4093
2 65703 1 4093
2 65704 1 4093
2 65705 1 4093
2 65706 1 4093
2 65707 1 4117
2 65708 1 4117
2 65709 1 4117
2 65710 1 4137
2 65711 1 4137
2 65712 1 4137
2 65713 1 4137
2 65714 1 4137
2 65715 1 4137
2 65716 1 4137
2 65717 1 4137
2 65718 1 4137
2 65719 1 4137
2 65720 1 4137
2 65721 1 4137
2 65722 1 4137
2 65723 1 4137
2 65724 1 4137
2 65725 1 4137
2 65726 1 4137
2 65727 1 4137
2 65728 1 4137
2 65729 1 4137
2 65730 1 4137
2 65731 1 4137
2 65732 1 4137
2 65733 1 4137
2 65734 1 4137
2 65735 1 4137
2 65736 1 4137
2 65737 1 4137
2 65738 1 4137
2 65739 1 4137
2 65740 1 4137
2 65741 1 4137
2 65742 1 4137
2 65743 1 4137
2 65744 1 4137
2 65745 1 4137
2 65746 1 4138
2 65747 1 4138
2 65748 1 4138
2 65749 1 4138
2 65750 1 4142
2 65751 1 4142
2 65752 1 4148
2 65753 1 4148
2 65754 1 4149
2 65755 1 4149
2 65756 1 4151
2 65757 1 4151
2 65758 1 4152
2 65759 1 4152
2 65760 1 4152
2 65761 1 4154
2 65762 1 4154
2 65763 1 4160
2 65764 1 4160
2 65765 1 4171
2 65766 1 4171
2 65767 1 4171
2 65768 1 4171
2 65769 1 4171
2 65770 1 4171
2 65771 1 4171
2 65772 1 4171
2 65773 1 4171
2 65774 1 4171
2 65775 1 4171
2 65776 1 4171
2 65777 1 4180
2 65778 1 4180
2 65779 1 4181
2 65780 1 4181
2 65781 1 4181
2 65782 1 4183
2 65783 1 4183
2 65784 1 4183
2 65785 1 4183
2 65786 1 4183
2 65787 1 4183
2 65788 1 4183
2 65789 1 4193
2 65790 1 4193
2 65791 1 4193
2 65792 1 4214
2 65793 1 4214
2 65794 1 4218
2 65795 1 4218
2 65796 1 4218
2 65797 1 4218
2 65798 1 4219
2 65799 1 4219
2 65800 1 4219
2 65801 1 4219
2 65802 1 4219
2 65803 1 4219
2 65804 1 4219
2 65805 1 4219
2 65806 1 4219
2 65807 1 4219
2 65808 1 4219
2 65809 1 4219
2 65810 1 4219
2 65811 1 4225
2 65812 1 4225
2 65813 1 4239
2 65814 1 4239
2 65815 1 4239
2 65816 1 4239
2 65817 1 4239
2 65818 1 4239
2 65819 1 4239
2 65820 1 4242
2 65821 1 4242
2 65822 1 4242
2 65823 1 4242
2 65824 1 4243
2 65825 1 4243
2 65826 1 4243
2 65827 1 4243
2 65828 1 4243
2 65829 1 4243
2 65830 1 4243
2 65831 1 4244
2 65832 1 4244
2 65833 1 4244
2 65834 1 4245
2 65835 1 4245
2 65836 1 4245
2 65837 1 4245
2 65838 1 4245
2 65839 1 4245
2 65840 1 4245
2 65841 1 4245
2 65842 1 4246
2 65843 1 4246
2 65844 1 4259
2 65845 1 4259
2 65846 1 4259
2 65847 1 4260
2 65848 1 4260
2 65849 1 4261
2 65850 1 4261
2 65851 1 4262
2 65852 1 4262
2 65853 1 4262
2 65854 1 4262
2 65855 1 4262
2 65856 1 4262
2 65857 1 4266
2 65858 1 4266
2 65859 1 4276
2 65860 1 4276
2 65861 1 4276
2 65862 1 4279
2 65863 1 4279
2 65864 1 4280
2 65865 1 4280
2 65866 1 4280
2 65867 1 4281
2 65868 1 4281
2 65869 1 4282
2 65870 1 4282
2 65871 1 4282
2 65872 1 4282
2 65873 1 4282
2 65874 1 4287
2 65875 1 4287
2 65876 1 4300
2 65877 1 4300
2 65878 1 4301
2 65879 1 4301
2 65880 1 4301
2 65881 1 4302
2 65882 1 4302
2 65883 1 4303
2 65884 1 4303
2 65885 1 4303
2 65886 1 4303
2 65887 1 4303
2 65888 1 4303
2 65889 1 4303
2 65890 1 4303
2 65891 1 4310
2 65892 1 4310
2 65893 1 4310
2 65894 1 4310
2 65895 1 4310
2 65896 1 4310
2 65897 1 4310
2 65898 1 4310
2 65899 1 4311
2 65900 1 4311
2 65901 1 4311
2 65902 1 4316
2 65903 1 4316
2 65904 1 4316
2 65905 1 4316
2 65906 1 4325
2 65907 1 4325
2 65908 1 4325
2 65909 1 4325
2 65910 1 4325
2 65911 1 4325
2 65912 1 4325
2 65913 1 4325
2 65914 1 4326
2 65915 1 4326
2 65916 1 4326
2 65917 1 4326
2 65918 1 4326
2 65919 1 4326
2 65920 1 4327
2 65921 1 4327
2 65922 1 4329
2 65923 1 4329
2 65924 1 4330
2 65925 1 4330
2 65926 1 4330
2 65927 1 4330
2 65928 1 4330
2 65929 1 4331
2 65930 1 4331
2 65931 1 4331
2 65932 1 4331
2 65933 1 4332
2 65934 1 4332
2 65935 1 4332
2 65936 1 4332
2 65937 1 4355
2 65938 1 4355
2 65939 1 4355
2 65940 1 4355
2 65941 1 4355
2 65942 1 4356
2 65943 1 4356
2 65944 1 4356
2 65945 1 4357
2 65946 1 4357
2 65947 1 4363
2 65948 1 4363
2 65949 1 4363
2 65950 1 4363
2 65951 1 4363
2 65952 1 4365
2 65953 1 4365
2 65954 1 4387
2 65955 1 4387
2 65956 1 4390
2 65957 1 4390
2 65958 1 4390
2 65959 1 4390
2 65960 1 4390
2 65961 1 4390
2 65962 1 4390
2 65963 1 4390
2 65964 1 4390
2 65965 1 4390
2 65966 1 4390
2 65967 1 4390
2 65968 1 4390
2 65969 1 4390
2 65970 1 4390
2 65971 1 4390
2 65972 1 4390
2 65973 1 4390
2 65974 1 4390
2 65975 1 4390
2 65976 1 4390
2 65977 1 4390
2 65978 1 4390
2 65979 1 4390
2 65980 1 4390
2 65981 1 4390
2 65982 1 4390
2 65983 1 4390
2 65984 1 4390
2 65985 1 4390
2 65986 1 4390
2 65987 1 4390
2 65988 1 4390
2 65989 1 4390
2 65990 1 4390
2 65991 1 4390
2 65992 1 4390
2 65993 1 4390
2 65994 1 4390
2 65995 1 4390
2 65996 1 4390
2 65997 1 4390
2 65998 1 4390
2 65999 1 4390
2 66000 1 4391
2 66001 1 4391
2 66002 1 4392
2 66003 1 4392
2 66004 1 4392
2 66005 1 4392
2 66006 1 4392
2 66007 1 4393
2 66008 1 4393
2 66009 1 4393
2 66010 1 4393
2 66011 1 4393
2 66012 1 4394
2 66013 1 4394
2 66014 1 4394
2 66015 1 4404
2 66016 1 4404
2 66017 1 4416
2 66018 1 4416
2 66019 1 4418
2 66020 1 4418
2 66021 1 4418
2 66022 1 4426
2 66023 1 4426
2 66024 1 4426
2 66025 1 4426
2 66026 1 4426
2 66027 1 4426
2 66028 1 4426
2 66029 1 4426
2 66030 1 4426
2 66031 1 4426
2 66032 1 4426
2 66033 1 4426
2 66034 1 4426
2 66035 1 4427
2 66036 1 4427
2 66037 1 4428
2 66038 1 4428
2 66039 1 4428
2 66040 1 4428
2 66041 1 4428
2 66042 1 4430
2 66043 1 4430
2 66044 1 4430
2 66045 1 4430
2 66046 1 4430
2 66047 1 4430
2 66048 1 4430
2 66049 1 4430
2 66050 1 4430
2 66051 1 4430
2 66052 1 4430
2 66053 1 4430
2 66054 1 4430
2 66055 1 4430
2 66056 1 4431
2 66057 1 4431
2 66058 1 4431
2 66059 1 4431
2 66060 1 4431
2 66061 1 4432
2 66062 1 4432
2 66063 1 4432
2 66064 1 4432
2 66065 1 4432
2 66066 1 4432
2 66067 1 4432
2 66068 1 4432
2 66069 1 4432
2 66070 1 4432
2 66071 1 4432
2 66072 1 4432
2 66073 1 4432
2 66074 1 4432
2 66075 1 4432
2 66076 1 4432
2 66077 1 4432
2 66078 1 4432
2 66079 1 4432
2 66080 1 4432
2 66081 1 4432
2 66082 1 4432
2 66083 1 4432
2 66084 1 4432
2 66085 1 4432
2 66086 1 4432
2 66087 1 4432
2 66088 1 4432
2 66089 1 4432
2 66090 1 4432
2 66091 1 4432
2 66092 1 4432
2 66093 1 4432
2 66094 1 4432
2 66095 1 4432
2 66096 1 4432
2 66097 1 4432
2 66098 1 4432
2 66099 1 4432
2 66100 1 4432
2 66101 1 4432
2 66102 1 4432
2 66103 1 4432
2 66104 1 4432
2 66105 1 4432
2 66106 1 4432
2 66107 1 4432
2 66108 1 4432
2 66109 1 4432
2 66110 1 4433
2 66111 1 4433
2 66112 1 4433
2 66113 1 4433
2 66114 1 4433
2 66115 1 4433
2 66116 1 4433
2 66117 1 4434
2 66118 1 4434
2 66119 1 4437
2 66120 1 4437
2 66121 1 4437
2 66122 1 4437
2 66123 1 4437
2 66124 1 4437
2 66125 1 4439
2 66126 1 4439
2 66127 1 4444
2 66128 1 4444
2 66129 1 4445
2 66130 1 4445
2 66131 1 4447
2 66132 1 4447
2 66133 1 4458
2 66134 1 4458
2 66135 1 4471
2 66136 1 4471
2 66137 1 4472
2 66138 1 4472
2 66139 1 4474
2 66140 1 4474
2 66141 1 4476
2 66142 1 4476
2 66143 1 4491
2 66144 1 4491
2 66145 1 4495
2 66146 1 4495
2 66147 1 4506
2 66148 1 4506
2 66149 1 4508
2 66150 1 4508
2 66151 1 4508
2 66152 1 4521
2 66153 1 4521
2 66154 1 4521
2 66155 1 4521
2 66156 1 4521
2 66157 1 4521
2 66158 1 4521
2 66159 1 4521
2 66160 1 4522
2 66161 1 4522
2 66162 1 4523
2 66163 1 4523
2 66164 1 4524
2 66165 1 4524
2 66166 1 4528
2 66167 1 4528
2 66168 1 4528
2 66169 1 4528
2 66170 1 4529
2 66171 1 4529
2 66172 1 4529
2 66173 1 4536
2 66174 1 4536
2 66175 1 4536
2 66176 1 4536
2 66177 1 4536
2 66178 1 4538
2 66179 1 4538
2 66180 1 4547
2 66181 1 4547
2 66182 1 4549
2 66183 1 4549
2 66184 1 4565
2 66185 1 4565
2 66186 1 4566
2 66187 1 4566
2 66188 1 4591
2 66189 1 4591
2 66190 1 4591
2 66191 1 4591
2 66192 1 4591
2 66193 1 4591
2 66194 1 4592
2 66195 1 4592
2 66196 1 4593
2 66197 1 4593
2 66198 1 4593
2 66199 1 4593
2 66200 1 4594
2 66201 1 4594
2 66202 1 4594
2 66203 1 4594
2 66204 1 4594
2 66205 1 4594
2 66206 1 4594
2 66207 1 4594
2 66208 1 4595
2 66209 1 4595
2 66210 1 4614
2 66211 1 4614
2 66212 1 4614
2 66213 1 4626
2 66214 1 4626
2 66215 1 4626
2 66216 1 4626
2 66217 1 4626
2 66218 1 4626
2 66219 1 4626
2 66220 1 4626
2 66221 1 4626
2 66222 1 4635
2 66223 1 4635
2 66224 1 4635
2 66225 1 4637
2 66226 1 4637
2 66227 1 4638
2 66228 1 4638
2 66229 1 4640
2 66230 1 4640
2 66231 1 4649
2 66232 1 4649
2 66233 1 4649
2 66234 1 4649
2 66235 1 4649
2 66236 1 4649
2 66237 1 4649
2 66238 1 4650
2 66239 1 4650
2 66240 1 4651
2 66241 1 4651
2 66242 1 4663
2 66243 1 4663
2 66244 1 4663
2 66245 1 4663
2 66246 1 4663
2 66247 1 4663
2 66248 1 4663
2 66249 1 4663
2 66250 1 4663
2 66251 1 4663
2 66252 1 4663
2 66253 1 4663
2 66254 1 4663
2 66255 1 4663
2 66256 1 4663
2 66257 1 4663
2 66258 1 4663
2 66259 1 4665
2 66260 1 4665
2 66261 1 4665
2 66262 1 4668
2 66263 1 4668
2 66264 1 4669
2 66265 1 4669
2 66266 1 4669
2 66267 1 4669
2 66268 1 4669
2 66269 1 4677
2 66270 1 4677
2 66271 1 4677
2 66272 1 4677
2 66273 1 4677
2 66274 1 4677
2 66275 1 4677
2 66276 1 4677
2 66277 1 4677
2 66278 1 4677
2 66279 1 4677
2 66280 1 4677
2 66281 1 4677
2 66282 1 4677
2 66283 1 4677
2 66284 1 4678
2 66285 1 4678
2 66286 1 4678
2 66287 1 4679
2 66288 1 4679
2 66289 1 4679
2 66290 1 4679
2 66291 1 4679
2 66292 1 4679
2 66293 1 4679
2 66294 1 4679
2 66295 1 4679
2 66296 1 4679
2 66297 1 4679
2 66298 1 4679
2 66299 1 4679
2 66300 1 4679
2 66301 1 4679
2 66302 1 4679
2 66303 1 4680
2 66304 1 4680
2 66305 1 4680
2 66306 1 4680
2 66307 1 4680
2 66308 1 4680
2 66309 1 4680
2 66310 1 4680
2 66311 1 4680
2 66312 1 4680
2 66313 1 4680
2 66314 1 4680
2 66315 1 4680
2 66316 1 4681
2 66317 1 4681
2 66318 1 4681
2 66319 1 4681
2 66320 1 4696
2 66321 1 4696
2 66322 1 4697
2 66323 1 4697
2 66324 1 4697
2 66325 1 4697
2 66326 1 4710
2 66327 1 4710
2 66328 1 4710
2 66329 1 4710
2 66330 1 4710
2 66331 1 4711
2 66332 1 4711
2 66333 1 4712
2 66334 1 4712
2 66335 1 4732
2 66336 1 4732
2 66337 1 4732
2 66338 1 4732
2 66339 1 4732
2 66340 1 4733
2 66341 1 4733
2 66342 1 4741
2 66343 1 4741
2 66344 1 4741
2 66345 1 4744
2 66346 1 4744
2 66347 1 4744
2 66348 1 4744
2 66349 1 4744
2 66350 1 4744
2 66351 1 4744
2 66352 1 4744
2 66353 1 4744
2 66354 1 4744
2 66355 1 4745
2 66356 1 4745
2 66357 1 4745
2 66358 1 4745
2 66359 1 4746
2 66360 1 4746
2 66361 1 4759
2 66362 1 4759
2 66363 1 4772
2 66364 1 4772
2 66365 1 4772
2 66366 1 4772
2 66367 1 4772
2 66368 1 4799
2 66369 1 4799
2 66370 1 4799
2 66371 1 4799
2 66372 1 4799
2 66373 1 4799
2 66374 1 4799
2 66375 1 4799
2 66376 1 4799
2 66377 1 4799
2 66378 1 4799
2 66379 1 4799
2 66380 1 4799
2 66381 1 4800
2 66382 1 4800
2 66383 1 4801
2 66384 1 4801
2 66385 1 4803
2 66386 1 4803
2 66387 1 4803
2 66388 1 4804
2 66389 1 4804
2 66390 1 4806
2 66391 1 4806
2 66392 1 4806
2 66393 1 4806
2 66394 1 4806
2 66395 1 4806
2 66396 1 4806
2 66397 1 4806
2 66398 1 4806
2 66399 1 4806
2 66400 1 4806
2 66401 1 4806
2 66402 1 4807
2 66403 1 4807
2 66404 1 4807
2 66405 1 4807
2 66406 1 4807
2 66407 1 4809
2 66408 1 4809
2 66409 1 4809
2 66410 1 4809
2 66411 1 4809
2 66412 1 4809
2 66413 1 4809
2 66414 1 4809
2 66415 1 4809
2 66416 1 4809
2 66417 1 4809
2 66418 1 4809
2 66419 1 4809
2 66420 1 4809
2 66421 1 4809
2 66422 1 4809
2 66423 1 4809
2 66424 1 4809
2 66425 1 4809
2 66426 1 4809
2 66427 1 4809
2 66428 1 4810
2 66429 1 4810
2 66430 1 4810
2 66431 1 4810
2 66432 1 4810
2 66433 1 4810
2 66434 1 4811
2 66435 1 4811
2 66436 1 4811
2 66437 1 4811
2 66438 1 4811
2 66439 1 4811
2 66440 1 4811
2 66441 1 4811
2 66442 1 4812
2 66443 1 4812
2 66444 1 4812
2 66445 1 4812
2 66446 1 4812
2 66447 1 4812
2 66448 1 4812
2 66449 1 4812
2 66450 1 4812
2 66451 1 4812
2 66452 1 4814
2 66453 1 4814
2 66454 1 4816
2 66455 1 4816
2 66456 1 4819
2 66457 1 4819
2 66458 1 4819
2 66459 1 4819
2 66460 1 4819
2 66461 1 4819
2 66462 1 4819
2 66463 1 4819
2 66464 1 4819
2 66465 1 4819
2 66466 1 4819
2 66467 1 4819
2 66468 1 4819
2 66469 1 4819
2 66470 1 4819
2 66471 1 4819
2 66472 1 4819
2 66473 1 4819
2 66474 1 4819
2 66475 1 4819
2 66476 1 4819
2 66477 1 4819
2 66478 1 4819
2 66479 1 4819
2 66480 1 4819
2 66481 1 4819
2 66482 1 4820
2 66483 1 4820
2 66484 1 4821
2 66485 1 4821
2 66486 1 4821
2 66487 1 4821
2 66488 1 4832
2 66489 1 4832
2 66490 1 4832
2 66491 1 4832
2 66492 1 4832
2 66493 1 4832
2 66494 1 4833
2 66495 1 4833
2 66496 1 4833
2 66497 1 4833
2 66498 1 4833
2 66499 1 4833
2 66500 1 4833
2 66501 1 4833
2 66502 1 4834
2 66503 1 4834
2 66504 1 4846
2 66505 1 4846
2 66506 1 4846
2 66507 1 4846
2 66508 1 4846
2 66509 1 4847
2 66510 1 4847
2 66511 1 4847
2 66512 1 4847
2 66513 1 4848
2 66514 1 4848
2 66515 1 4848
2 66516 1 4848
2 66517 1 4848
2 66518 1 4848
2 66519 1 4848
2 66520 1 4848
2 66521 1 4848
2 66522 1 4848
2 66523 1 4850
2 66524 1 4850
2 66525 1 4851
2 66526 1 4851
2 66527 1 4851
2 66528 1 4851
2 66529 1 4851
2 66530 1 4852
2 66531 1 4852
2 66532 1 4859
2 66533 1 4859
2 66534 1 4859
2 66535 1 4859
2 66536 1 4859
2 66537 1 4859
2 66538 1 4860
2 66539 1 4860
2 66540 1 4860
2 66541 1 4867
2 66542 1 4867
2 66543 1 4867
2 66544 1 4868
2 66545 1 4868
2 66546 1 4869
2 66547 1 4869
2 66548 1 4877
2 66549 1 4877
2 66550 1 4877
2 66551 1 4877
2 66552 1 4877
2 66553 1 4877
2 66554 1 4878
2 66555 1 4878
2 66556 1 4879
2 66557 1 4879
2 66558 1 4880
2 66559 1 4880
2 66560 1 4881
2 66561 1 4881
2 66562 1 4881
2 66563 1 4886
2 66564 1 4886
2 66565 1 4907
2 66566 1 4907
2 66567 1 4908
2 66568 1 4908
2 66569 1 4908
2 66570 1 4908
2 66571 1 4908
2 66572 1 4916
2 66573 1 4916
2 66574 1 4924
2 66575 1 4924
2 66576 1 4924
2 66577 1 4924
2 66578 1 4924
2 66579 1 4924
2 66580 1 4924
2 66581 1 4924
2 66582 1 4924
2 66583 1 4924
2 66584 1 4924
2 66585 1 4924
2 66586 1 4924
2 66587 1 4931
2 66588 1 4931
2 66589 1 4932
2 66590 1 4932
2 66591 1 4932
2 66592 1 4932
2 66593 1 4932
2 66594 1 4932
2 66595 1 4932
2 66596 1 4932
2 66597 1 4932
2 66598 1 4932
2 66599 1 4932
2 66600 1 4932
2 66601 1 4932
2 66602 1 4932
2 66603 1 4932
2 66604 1 4932
2 66605 1 4932
2 66606 1 4932
2 66607 1 4932
2 66608 1 4932
2 66609 1 4932
2 66610 1 4932
2 66611 1 4932
2 66612 1 4932
2 66613 1 4932
2 66614 1 4932
2 66615 1 4932
2 66616 1 4932
2 66617 1 4943
2 66618 1 4943
2 66619 1 4943
2 66620 1 4944
2 66621 1 4944
2 66622 1 4947
2 66623 1 4947
2 66624 1 4947
2 66625 1 4948
2 66626 1 4948
2 66627 1 4948
2 66628 1 4949
2 66629 1 4949
2 66630 1 4949
2 66631 1 4949
2 66632 1 4949
2 66633 1 4949
2 66634 1 4949
2 66635 1 4949
2 66636 1 4949
2 66637 1 4950
2 66638 1 4950
2 66639 1 4950
2 66640 1 4950
2 66641 1 4950
2 66642 1 4950
2 66643 1 4950
2 66644 1 4950
2 66645 1 4951
2 66646 1 4951
2 66647 1 4951
2 66648 1 4951
2 66649 1 4951
2 66650 1 4951
2 66651 1 4951
2 66652 1 4951
2 66653 1 4951
2 66654 1 4951
2 66655 1 4951
2 66656 1 4951
2 66657 1 4951
2 66658 1 4951
2 66659 1 4951
2 66660 1 4951
2 66661 1 4951
2 66662 1 4951
2 66663 1 4951
2 66664 1 4951
2 66665 1 4951
2 66666 1 4951
2 66667 1 4951
2 66668 1 4951
2 66669 1 4951
2 66670 1 4951
2 66671 1 4951
2 66672 1 4951
2 66673 1 4951
2 66674 1 4963
2 66675 1 4963
2 66676 1 4964
2 66677 1 4964
2 66678 1 4964
2 66679 1 4964
2 66680 1 4964
2 66681 1 4964
2 66682 1 4972
2 66683 1 4972
2 66684 1 4972
2 66685 1 4972
2 66686 1 4974
2 66687 1 4974
2 66688 1 4974
2 66689 1 4974
2 66690 1 4974
2 66691 1 4976
2 66692 1 4976
2 66693 1 4976
2 66694 1 4978
2 66695 1 4978
2 66696 1 4982
2 66697 1 4982
2 66698 1 4982
2 66699 1 4982
2 66700 1 4982
2 66701 1 4982
2 66702 1 4982
2 66703 1 4982
2 66704 1 4982
2 66705 1 4982
2 66706 1 4982
2 66707 1 4982
2 66708 1 4982
2 66709 1 4983
2 66710 1 4983
2 66711 1 4983
2 66712 1 4983
2 66713 1 4983
2 66714 1 4986
2 66715 1 4986
2 66716 1 4986
2 66717 1 4987
2 66718 1 4987
2 66719 1 5000
2 66720 1 5000
2 66721 1 5000
2 66722 1 5000
2 66723 1 5000
2 66724 1 5000
2 66725 1 5001
2 66726 1 5001
2 66727 1 5009
2 66728 1 5009
2 66729 1 5009
2 66730 1 5016
2 66731 1 5016
2 66732 1 5016
2 66733 1 5016
2 66734 1 5016
2 66735 1 5016
2 66736 1 5016
2 66737 1 5016
2 66738 1 5016
2 66739 1 5016
2 66740 1 5016
2 66741 1 5016
2 66742 1 5016
2 66743 1 5016
2 66744 1 5022
2 66745 1 5022
2 66746 1 5022
2 66747 1 5022
2 66748 1 5023
2 66749 1 5023
2 66750 1 5027
2 66751 1 5027
2 66752 1 5027
2 66753 1 5027
2 66754 1 5027
2 66755 1 5027
2 66756 1 5027
2 66757 1 5027
2 66758 1 5027
2 66759 1 5027
2 66760 1 5027
2 66761 1 5027
2 66762 1 5027
2 66763 1 5027
2 66764 1 5027
2 66765 1 5027
2 66766 1 5027
2 66767 1 5027
2 66768 1 5027
2 66769 1 5027
2 66770 1 5029
2 66771 1 5029
2 66772 1 5029
2 66773 1 5029
2 66774 1 5029
2 66775 1 5037
2 66776 1 5037
2 66777 1 5039
2 66778 1 5039
2 66779 1 5039
2 66780 1 5039
2 66781 1 5039
2 66782 1 5046
2 66783 1 5046
2 66784 1 5046
2 66785 1 5046
2 66786 1 5046
2 66787 1 5064
2 66788 1 5064
2 66789 1 5065
2 66790 1 5065
2 66791 1 5074
2 66792 1 5074
2 66793 1 5077
2 66794 1 5077
2 66795 1 5078
2 66796 1 5078
2 66797 1 5078
2 66798 1 5078
2 66799 1 5078
2 66800 1 5078
2 66801 1 5078
2 66802 1 5079
2 66803 1 5079
2 66804 1 5079
2 66805 1 5079
2 66806 1 5080
2 66807 1 5080
2 66808 1 5080
2 66809 1 5082
2 66810 1 5082
2 66811 1 5083
2 66812 1 5083
2 66813 1 5083
2 66814 1 5083
2 66815 1 5083
2 66816 1 5083
2 66817 1 5083
2 66818 1 5083
2 66819 1 5083
2 66820 1 5083
2 66821 1 5083
2 66822 1 5084
2 66823 1 5084
2 66824 1 5084
2 66825 1 5084
2 66826 1 5100
2 66827 1 5100
2 66828 1 5100
2 66829 1 5104
2 66830 1 5104
2 66831 1 5108
2 66832 1 5108
2 66833 1 5125
2 66834 1 5125
2 66835 1 5140
2 66836 1 5140
2 66837 1 5140
2 66838 1 5141
2 66839 1 5141
2 66840 1 5141
2 66841 1 5147
2 66842 1 5147
2 66843 1 5147
2 66844 1 5147
2 66845 1 5148
2 66846 1 5148
2 66847 1 5148
2 66848 1 5151
2 66849 1 5151
2 66850 1 5154
2 66851 1 5154
2 66852 1 5154
2 66853 1 5154
2 66854 1 5155
2 66855 1 5155
2 66856 1 5163
2 66857 1 5163
2 66858 1 5165
2 66859 1 5165
2 66860 1 5165
2 66861 1 5165
2 66862 1 5165
2 66863 1 5165
2 66864 1 5166
2 66865 1 5166
2 66866 1 5166
2 66867 1 5166
2 66868 1 5167
2 66869 1 5167
2 66870 1 5168
2 66871 1 5168
2 66872 1 5168
2 66873 1 5186
2 66874 1 5186
2 66875 1 5188
2 66876 1 5188
2 66877 1 5188
2 66878 1 5188
2 66879 1 5189
2 66880 1 5189
2 66881 1 5202
2 66882 1 5202
2 66883 1 5202
2 66884 1 5202
2 66885 1 5202
2 66886 1 5202
2 66887 1 5202
2 66888 1 5202
2 66889 1 5202
2 66890 1 5202
2 66891 1 5202
2 66892 1 5202
2 66893 1 5203
2 66894 1 5203
2 66895 1 5203
2 66896 1 5204
2 66897 1 5204
2 66898 1 5204
2 66899 1 5204
2 66900 1 5204
2 66901 1 5204
2 66902 1 5204
2 66903 1 5204
2 66904 1 5205
2 66905 1 5205
2 66906 1 5205
2 66907 1 5205
2 66908 1 5206
2 66909 1 5206
2 66910 1 5213
2 66911 1 5213
2 66912 1 5213
2 66913 1 5216
2 66914 1 5216
2 66915 1 5216
2 66916 1 5232
2 66917 1 5232
2 66918 1 5232
2 66919 1 5232
2 66920 1 5232
2 66921 1 5236
2 66922 1 5236
2 66923 1 5245
2 66924 1 5245
2 66925 1 5246
2 66926 1 5246
2 66927 1 5247
2 66928 1 5247
2 66929 1 5247
2 66930 1 5247
2 66931 1 5249
2 66932 1 5249
2 66933 1 5256
2 66934 1 5256
2 66935 1 5256
2 66936 1 5257
2 66937 1 5257
2 66938 1 5264
2 66939 1 5264
2 66940 1 5267
2 66941 1 5267
2 66942 1 5306
2 66943 1 5306
2 66944 1 5307
2 66945 1 5307
2 66946 1 5316
2 66947 1 5316
2 66948 1 5331
2 66949 1 5331
2 66950 1 5333
2 66951 1 5333
2 66952 1 5358
2 66953 1 5358
2 66954 1 5364
2 66955 1 5364
2 66956 1 5364
2 66957 1 5364
2 66958 1 5364
2 66959 1 5364
2 66960 1 5364
2 66961 1 5364
2 66962 1 5364
2 66963 1 5364
2 66964 1 5364
2 66965 1 5364
2 66966 1 5364
2 66967 1 5364
2 66968 1 5365
2 66969 1 5365
2 66970 1 5373
2 66971 1 5373
2 66972 1 5373
2 66973 1 5373
2 66974 1 5373
2 66975 1 5373
2 66976 1 5373
2 66977 1 5373
2 66978 1 5376
2 66979 1 5376
2 66980 1 5376
2 66981 1 5376
2 66982 1 5376
2 66983 1 5376
2 66984 1 5376
2 66985 1 5376
2 66986 1 5376
2 66987 1 5376
2 66988 1 5386
2 66989 1 5386
2 66990 1 5386
2 66991 1 5386
2 66992 1 5386
2 66993 1 5386
2 66994 1 5395
2 66995 1 5395
2 66996 1 5397
2 66997 1 5397
2 66998 1 5397
2 66999 1 5397
2 67000 1 5397
2 67001 1 5397
2 67002 1 5397
2 67003 1 5399
2 67004 1 5399
2 67005 1 5406
2 67006 1 5406
2 67007 1 5406
2 67008 1 5406
2 67009 1 5406
2 67010 1 5406
2 67011 1 5406
2 67012 1 5406
2 67013 1 5406
2 67014 1 5406
2 67015 1 5406
2 67016 1 5406
2 67017 1 5406
2 67018 1 5406
2 67019 1 5407
2 67020 1 5407
2 67021 1 5407
2 67022 1 5414
2 67023 1 5414
2 67024 1 5414
2 67025 1 5417
2 67026 1 5417
2 67027 1 5417
2 67028 1 5417
2 67029 1 5417
2 67030 1 5417
2 67031 1 5417
2 67032 1 5417
2 67033 1 5417
2 67034 1 5419
2 67035 1 5419
2 67036 1 5420
2 67037 1 5420
2 67038 1 5420
2 67039 1 5420
2 67040 1 5420
2 67041 1 5421
2 67042 1 5421
2 67043 1 5428
2 67044 1 5428
2 67045 1 5435
2 67046 1 5435
2 67047 1 5435
2 67048 1 5435
2 67049 1 5435
2 67050 1 5435
2 67051 1 5436
2 67052 1 5436
2 67053 1 5450
2 67054 1 5450
2 67055 1 5450
2 67056 1 5450
2 67057 1 5450
2 67058 1 5451
2 67059 1 5451
2 67060 1 5451
2 67061 1 5451
2 67062 1 5452
2 67063 1 5452
2 67064 1 5452
2 67065 1 5452
2 67066 1 5452
2 67067 1 5452
2 67068 1 5452
2 67069 1 5460
2 67070 1 5460
2 67071 1 5460
2 67072 1 5464
2 67073 1 5464
2 67074 1 5472
2 67075 1 5472
2 67076 1 5473
2 67077 1 5473
2 67078 1 5473
2 67079 1 5474
2 67080 1 5474
2 67081 1 5482
2 67082 1 5482
2 67083 1 5490
2 67084 1 5490
2 67085 1 5490
2 67086 1 5490
2 67087 1 5491
2 67088 1 5491
2 67089 1 5499
2 67090 1 5499
2 67091 1 5499
2 67092 1 5499
2 67093 1 5506
2 67094 1 5506
2 67095 1 5506
2 67096 1 5506
2 67097 1 5506
2 67098 1 5506
2 67099 1 5507
2 67100 1 5507
2 67101 1 5507
2 67102 1 5527
2 67103 1 5527
2 67104 1 5527
2 67105 1 5530
2 67106 1 5530
2 67107 1 5531
2 67108 1 5531
2 67109 1 5531
2 67110 1 5531
2 67111 1 5531
2 67112 1 5532
2 67113 1 5532
2 67114 1 5532
2 67115 1 5532
2 67116 1 5532
2 67117 1 5532
2 67118 1 5532
2 67119 1 5532
2 67120 1 5532
2 67121 1 5532
2 67122 1 5532
2 67123 1 5532
2 67124 1 5532
2 67125 1 5532
2 67126 1 5532
2 67127 1 5532
2 67128 1 5532
2 67129 1 5532
2 67130 1 5533
2 67131 1 5533
2 67132 1 5533
2 67133 1 5533
2 67134 1 5533
2 67135 1 5533
2 67136 1 5533
2 67137 1 5533
2 67138 1 5545
2 67139 1 5545
2 67140 1 5545
2 67141 1 5545
2 67142 1 5547
2 67143 1 5547
2 67144 1 5555
2 67145 1 5555
2 67146 1 5555
2 67147 1 5556
2 67148 1 5556
2 67149 1 5559
2 67150 1 5559
2 67151 1 5559
2 67152 1 5559
2 67153 1 5572
2 67154 1 5572
2 67155 1 5572
2 67156 1 5573
2 67157 1 5573
2 67158 1 5599
2 67159 1 5599
2 67160 1 5599
2 67161 1 5599
2 67162 1 5599
2 67163 1 5599
2 67164 1 5599
2 67165 1 5600
2 67166 1 5600
2 67167 1 5604
2 67168 1 5604
2 67169 1 5608
2 67170 1 5608
2 67171 1 5624
2 67172 1 5624
2 67173 1 5624
2 67174 1 5624
2 67175 1 5624
2 67176 1 5624
2 67177 1 5624
2 67178 1 5624
2 67179 1 5624
2 67180 1 5624
2 67181 1 5624
2 67182 1 5624
2 67183 1 5624
2 67184 1 5624
2 67185 1 5624
2 67186 1 5624
2 67187 1 5624
2 67188 1 5624
2 67189 1 5624
2 67190 1 5624
2 67191 1 5624
2 67192 1 5625
2 67193 1 5625
2 67194 1 5626
2 67195 1 5626
2 67196 1 5646
2 67197 1 5646
2 67198 1 5646
2 67199 1 5646
2 67200 1 5646
2 67201 1 5646
2 67202 1 5646
2 67203 1 5646
2 67204 1 5646
2 67205 1 5646
2 67206 1 5647
2 67207 1 5647
2 67208 1 5647
2 67209 1 5647
2 67210 1 5647
2 67211 1 5647
2 67212 1 5647
2 67213 1 5647
2 67214 1 5647
2 67215 1 5647
2 67216 1 5647
2 67217 1 5647
2 67218 1 5647
2 67219 1 5647
2 67220 1 5647
2 67221 1 5647
2 67222 1 5647
2 67223 1 5647
2 67224 1 5647
2 67225 1 5647
2 67226 1 5647
2 67227 1 5647
2 67228 1 5647
2 67229 1 5647
2 67230 1 5647
2 67231 1 5647
2 67232 1 5647
2 67233 1 5647
2 67234 1 5648
2 67235 1 5648
2 67236 1 5648
2 67237 1 5648
2 67238 1 5648
2 67239 1 5648
2 67240 1 5648
2 67241 1 5649
2 67242 1 5649
2 67243 1 5650
2 67244 1 5650
2 67245 1 5658
2 67246 1 5658
2 67247 1 5686
2 67248 1 5686
2 67249 1 5694
2 67250 1 5694
2 67251 1 5695
2 67252 1 5695
2 67253 1 5695
2 67254 1 5695
2 67255 1 5695
2 67256 1 5695
2 67257 1 5695
2 67258 1 5703
2 67259 1 5703
2 67260 1 5704
2 67261 1 5704
2 67262 1 5704
2 67263 1 5704
2 67264 1 5712
2 67265 1 5712
2 67266 1 5712
2 67267 1 5720
2 67268 1 5720
2 67269 1 5730
2 67270 1 5730
2 67271 1 5733
2 67272 1 5733
2 67273 1 5745
2 67274 1 5745
2 67275 1 5745
2 67276 1 5745
2 67277 1 5746
2 67278 1 5746
2 67279 1 5746
2 67280 1 5753
2 67281 1 5753
2 67282 1 5755
2 67283 1 5755
2 67284 1 5755
2 67285 1 5756
2 67286 1 5756
2 67287 1 5756
2 67288 1 5756
2 67289 1 5764
2 67290 1 5764
2 67291 1 5772
2 67292 1 5772
2 67293 1 5772
2 67294 1 5772
2 67295 1 5779
2 67296 1 5779
2 67297 1 5779
2 67298 1 5779
2 67299 1 5779
2 67300 1 5779
2 67301 1 5779
2 67302 1 5780
2 67303 1 5780
2 67304 1 5780
2 67305 1 5791
2 67306 1 5791
2 67307 1 5791
2 67308 1 5791
2 67309 1 5794
2 67310 1 5794
2 67311 1 5821
2 67312 1 5821
2 67313 1 5821
2 67314 1 5829
2 67315 1 5829
2 67316 1 5863
2 67317 1 5863
2 67318 1 5874
2 67319 1 5874
2 67320 1 5874
2 67321 1 5882
2 67322 1 5882
2 67323 1 5901
2 67324 1 5901
2 67325 1 5901
2 67326 1 5901
2 67327 1 5901
2 67328 1 5901
2 67329 1 5901
2 67330 1 5901
2 67331 1 5901
2 67332 1 5901
2 67333 1 5901
2 67334 1 5901
2 67335 1 5901
2 67336 1 5901
2 67337 1 5901
2 67338 1 5901
2 67339 1 5901
2 67340 1 5902
2 67341 1 5902
2 67342 1 5902
2 67343 1 5902
2 67344 1 5902
2 67345 1 5903
2 67346 1 5903
2 67347 1 5903
2 67348 1 5903
2 67349 1 5903
2 67350 1 5903
2 67351 1 5904
2 67352 1 5904
2 67353 1 5910
2 67354 1 5910
2 67355 1 5926
2 67356 1 5926
2 67357 1 5939
2 67358 1 5939
2 67359 1 5940
2 67360 1 5940
2 67361 1 5952
2 67362 1 5952
2 67363 1 5955
2 67364 1 5955
2 67365 1 5955
2 67366 1 5956
2 67367 1 5956
2 67368 1 5957
2 67369 1 5957
2 67370 1 5957
2 67371 1 5976
2 67372 1 5976
2 67373 1 5976
2 67374 1 5977
2 67375 1 5977
2 67376 1 5987
2 67377 1 5987
2 67378 1 5988
2 67379 1 5988
2 67380 1 5999
2 67381 1 5999
2 67382 1 5999
2 67383 1 6005
2 67384 1 6005
2 67385 1 6007
2 67386 1 6007
2 67387 1 6027
2 67388 1 6027
2 67389 1 6028
2 67390 1 6028
2 67391 1 6037
2 67392 1 6037
2 67393 1 6060
2 67394 1 6060
2 67395 1 6060
2 67396 1 6060
2 67397 1 6060
2 67398 1 6060
2 67399 1 6060
2 67400 1 6060
2 67401 1 6060
2 67402 1 6060
2 67403 1 6060
2 67404 1 6060
2 67405 1 6060
2 67406 1 6060
2 67407 1 6060
2 67408 1 6060
2 67409 1 6060
2 67410 1 6060
2 67411 1 6060
2 67412 1 6060
2 67413 1 6060
2 67414 1 6076
2 67415 1 6076
2 67416 1 6079
2 67417 1 6079
2 67418 1 6079
2 67419 1 6079
2 67420 1 6079
2 67421 1 6079
2 67422 1 6079
2 67423 1 6106
2 67424 1 6106
2 67425 1 6106
2 67426 1 6106
2 67427 1 6127
2 67428 1 6127
2 67429 1 6128
2 67430 1 6128
2 67431 1 6128
2 67432 1 6137
2 67433 1 6137
2 67434 1 6141
2 67435 1 6141
2 67436 1 6156
2 67437 1 6156
2 67438 1 6156
2 67439 1 6156
2 67440 1 6165
2 67441 1 6165
2 67442 1 6165
2 67443 1 6165
2 67444 1 6165
2 67445 1 6165
2 67446 1 6165
2 67447 1 6183
2 67448 1 6183
2 67449 1 6183
2 67450 1 6185
2 67451 1 6185
2 67452 1 6186
2 67453 1 6186
2 67454 1 6197
2 67455 1 6197
2 67456 1 6216
2 67457 1 6216
2 67458 1 6216
2 67459 1 6218
2 67460 1 6218
2 67461 1 6246
2 67462 1 6246
2 67463 1 6246
2 67464 1 6267
2 67465 1 6267
2 67466 1 6268
2 67467 1 6268
2 67468 1 6270
2 67469 1 6270
2 67470 1 6291
2 67471 1 6291
2 67472 1 6291
2 67473 1 6291
2 67474 1 6299
2 67475 1 6299
2 67476 1 6299
2 67477 1 6299
2 67478 1 6299
2 67479 1 6299
2 67480 1 6306
2 67481 1 6306
2 67482 1 6307
2 67483 1 6307
2 67484 1 6354
2 67485 1 6354
2 67486 1 6357
2 67487 1 6357
2 67488 1 6357
2 67489 1 6366
2 67490 1 6366
2 67491 1 6366
2 67492 1 6367
2 67493 1 6367
2 67494 1 6367
2 67495 1 6368
2 67496 1 6368
2 67497 1 6368
2 67498 1 6375
2 67499 1 6375
2 67500 1 6376
2 67501 1 6376
2 67502 1 6376
2 67503 1 6378
2 67504 1 6378
2 67505 1 6386
2 67506 1 6386
2 67507 1 6387
2 67508 1 6387
2 67509 1 6388
2 67510 1 6388
2 67511 1 6388
2 67512 1 6388
2 67513 1 6388
2 67514 1 6388
2 67515 1 6389
2 67516 1 6389
2 67517 1 6392
2 67518 1 6392
2 67519 1 6392
2 67520 1 6392
2 67521 1 6392
2 67522 1 6422
2 67523 1 6422
2 67524 1 6422
2 67525 1 6422
2 67526 1 6422
2 67527 1 6422
2 67528 1 6422
2 67529 1 6422
2 67530 1 6422
2 67531 1 6422
2 67532 1 6422
2 67533 1 6422
2 67534 1 6422
2 67535 1 6422
2 67536 1 6422
2 67537 1 6423
2 67538 1 6423
2 67539 1 6423
2 67540 1 6437
2 67541 1 6437
2 67542 1 6437
2 67543 1 6437
2 67544 1 6437
2 67545 1 6437
2 67546 1 6437
2 67547 1 6439
2 67548 1 6439
2 67549 1 6444
2 67550 1 6444
2 67551 1 6444
2 67552 1 6444
2 67553 1 6444
2 67554 1 6444
2 67555 1 6444
2 67556 1 6444
2 67557 1 6444
2 67558 1 6444
2 67559 1 6445
2 67560 1 6445
2 67561 1 6445
2 67562 1 6445
2 67563 1 6446
2 67564 1 6446
2 67565 1 6458
2 67566 1 6458
2 67567 1 6458
2 67568 1 6458
2 67569 1 6458
2 67570 1 6458
2 67571 1 6458
2 67572 1 6458
2 67573 1 6458
2 67574 1 6461
2 67575 1 6461
2 67576 1 6482
2 67577 1 6482
2 67578 1 6485
2 67579 1 6485
2 67580 1 6485
2 67581 1 6485
2 67582 1 6485
2 67583 1 6485
2 67584 1 6485
2 67585 1 6485
2 67586 1 6507
2 67587 1 6507
2 67588 1 6507
2 67589 1 6521
2 67590 1 6521
2 67591 1 6524
2 67592 1 6524
2 67593 1 6535
2 67594 1 6535
2 67595 1 6535
2 67596 1 6535
2 67597 1 6545
2 67598 1 6545
2 67599 1 6552
2 67600 1 6552
2 67601 1 6575
2 67602 1 6575
2 67603 1 6577
2 67604 1 6577
2 67605 1 6579
2 67606 1 6579
2 67607 1 6579
2 67608 1 6585
2 67609 1 6585
2 67610 1 6585
2 67611 1 6585
2 67612 1 6585
2 67613 1 6585
2 67614 1 6585
2 67615 1 6585
2 67616 1 6585
2 67617 1 6585
2 67618 1 6585
2 67619 1 6586
2 67620 1 6586
2 67621 1 6586
2 67622 1 6587
2 67623 1 6587
2 67624 1 6597
2 67625 1 6597
2 67626 1 6618
2 67627 1 6618
2 67628 1 6619
2 67629 1 6619
2 67630 1 6632
2 67631 1 6632
2 67632 1 6632
2 67633 1 6632
2 67634 1 6632
2 67635 1 6632
2 67636 1 6632
2 67637 1 6633
2 67638 1 6633
2 67639 1 6646
2 67640 1 6646
2 67641 1 6646
2 67642 1 6649
2 67643 1 6649
2 67644 1 6649
2 67645 1 6649
2 67646 1 6649
2 67647 1 6649
2 67648 1 6650
2 67649 1 6650
2 67650 1 6670
2 67651 1 6670
2 67652 1 6670
2 67653 1 6670
2 67654 1 6670
2 67655 1 6670
2 67656 1 6670
2 67657 1 6670
2 67658 1 6670
2 67659 1 6670
2 67660 1 6682
2 67661 1 6682
2 67662 1 6682
2 67663 1 6695
2 67664 1 6695
2 67665 1 6723
2 67666 1 6723
2 67667 1 6723
2 67668 1 6744
2 67669 1 6744
2 67670 1 6757
2 67671 1 6757
2 67672 1 6779
2 67673 1 6779
2 67674 1 6779
2 67675 1 6779
2 67676 1 6779
2 67677 1 6779
2 67678 1 6779
2 67679 1 6779
2 67680 1 6779
2 67681 1 6779
2 67682 1 6779
2 67683 1 6779
2 67684 1 6779
2 67685 1 6779
2 67686 1 6779
2 67687 1 6779
2 67688 1 6780
2 67689 1 6780
2 67690 1 6780
2 67691 1 6780
2 67692 1 6781
2 67693 1 6781
2 67694 1 6781
2 67695 1 6781
2 67696 1 6781
2 67697 1 6781
2 67698 1 6781
2 67699 1 6781
2 67700 1 6782
2 67701 1 6782
2 67702 1 6812
2 67703 1 6812
2 67704 1 6813
2 67705 1 6813
2 67706 1 6821
2 67707 1 6821
2 67708 1 6853
2 67709 1 6853
2 67710 1 6854
2 67711 1 6854
2 67712 1 6854
2 67713 1 6855
2 67714 1 6855
2 67715 1 6864
2 67716 1 6864
2 67717 1 6864
2 67718 1 6864
2 67719 1 6864
2 67720 1 6864
2 67721 1 6868
2 67722 1 6868
2 67723 1 6879
2 67724 1 6879
2 67725 1 6879
2 67726 1 6880
2 67727 1 6880
2 67728 1 6881
2 67729 1 6881
2 67730 1 6881
2 67731 1 6881
2 67732 1 6881
2 67733 1 6881
2 67734 1 6882
2 67735 1 6882
2 67736 1 6882
2 67737 1 6884
2 67738 1 6884
2 67739 1 6887
2 67740 1 6887
2 67741 1 6917
2 67742 1 6917
2 67743 1 6917
2 67744 1 6925
2 67745 1 6925
2 67746 1 6947
2 67747 1 6947
2 67748 1 6948
2 67749 1 6948
2 67750 1 6948
2 67751 1 6948
2 67752 1 6948
2 67753 1 6948
2 67754 1 6948
2 67755 1 6948
2 67756 1 6948
2 67757 1 6948
2 67758 1 6948
2 67759 1 6949
2 67760 1 6949
2 67761 1 6949
2 67762 1 6949
2 67763 1 6949
2 67764 1 6949
2 67765 1 6949
2 67766 1 6949
2 67767 1 6949
2 67768 1 6949
2 67769 1 6949
2 67770 1 6949
2 67771 1 6949
2 67772 1 6949
2 67773 1 6949
2 67774 1 6949
2 67775 1 6949
2 67776 1 6949
2 67777 1 6949
2 67778 1 6949
2 67779 1 6949
2 67780 1 6949
2 67781 1 6949
2 67782 1 6949
2 67783 1 6949
2 67784 1 6949
2 67785 1 6949
2 67786 1 6949
2 67787 1 6949
2 67788 1 6949
2 67789 1 6949
2 67790 1 6949
2 67791 1 6949
2 67792 1 6949
2 67793 1 6949
2 67794 1 6949
2 67795 1 6950
2 67796 1 6950
2 67797 1 6950
2 67798 1 6950
2 67799 1 6950
2 67800 1 6950
2 67801 1 6950
2 67802 1 6950
2 67803 1 6950
2 67804 1 6952
2 67805 1 6952
2 67806 1 6955
2 67807 1 6955
2 67808 1 6955
2 67809 1 6955
2 67810 1 6955
2 67811 1 6955
2 67812 1 6955
2 67813 1 6955
2 67814 1 6955
2 67815 1 6955
2 67816 1 6958
2 67817 1 6958
2 67818 1 6958
2 67819 1 6960
2 67820 1 6960
2 67821 1 6961
2 67822 1 6961
2 67823 1 6961
2 67824 1 6961
2 67825 1 6961
2 67826 1 6961
2 67827 1 6961
2 67828 1 6961
2 67829 1 6961
2 67830 1 6961
2 67831 1 6961
2 67832 1 6961
2 67833 1 6961
2 67834 1 6961
2 67835 1 6961
2 67836 1 6969
2 67837 1 6969
2 67838 1 6969
2 67839 1 6969
2 67840 1 6969
2 67841 1 6969
2 67842 1 6969
2 67843 1 6970
2 67844 1 6970
2 67845 1 6970
2 67846 1 6971
2 67847 1 6971
2 67848 1 6971
2 67849 1 6971
2 67850 1 6971
2 67851 1 6972
2 67852 1 6972
2 67853 1 6972
2 67854 1 6972
2 67855 1 6972
2 67856 1 6972
2 67857 1 6972
2 67858 1 6972
2 67859 1 6972
2 67860 1 6972
2 67861 1 6972
2 67862 1 6972
2 67863 1 6972
2 67864 1 6972
2 67865 1 6972
2 67866 1 6972
2 67867 1 6972
2 67868 1 6972
2 67869 1 6972
2 67870 1 6972
2 67871 1 6973
2 67872 1 6973
2 67873 1 6973
2 67874 1 6973
2 67875 1 6973
2 67876 1 6973
2 67877 1 6974
2 67878 1 6974
2 67879 1 6975
2 67880 1 6975
2 67881 1 6975
2 67882 1 6975
2 67883 1 6975
2 67884 1 6975
2 67885 1 6975
2 67886 1 6975
2 67887 1 6975
2 67888 1 6975
2 67889 1 6975
2 67890 1 6975
2 67891 1 6975
2 67892 1 6978
2 67893 1 6978
2 67894 1 6978
2 67895 1 6978
2 67896 1 6991
2 67897 1 6991
2 67898 1 6991
2 67899 1 6991
2 67900 1 6991
2 67901 1 6991
2 67902 1 6991
2 67903 1 6991
2 67904 1 6991
2 67905 1 6992
2 67906 1 6992
2 67907 1 6992
2 67908 1 6992
2 67909 1 6992
2 67910 1 6992
2 67911 1 6992
2 67912 1 6992
2 67913 1 6992
2 67914 1 6992
2 67915 1 6992
2 67916 1 6992
2 67917 1 6992
2 67918 1 6992
2 67919 1 6992
2 67920 1 6992
2 67921 1 6992
2 67922 1 6992
2 67923 1 6992
2 67924 1 6992
2 67925 1 6992
2 67926 1 6992
2 67927 1 6992
2 67928 1 6992
2 67929 1 6992
2 67930 1 6992
2 67931 1 6992
2 67932 1 6992
2 67933 1 6992
2 67934 1 6992
2 67935 1 6992
2 67936 1 6992
2 67937 1 6992
2 67938 1 6992
2 67939 1 6992
2 67940 1 6992
2 67941 1 6992
2 67942 1 6992
2 67943 1 6992
2 67944 1 6992
2 67945 1 6992
2 67946 1 6992
2 67947 1 6992
2 67948 1 6992
2 67949 1 6992
2 67950 1 6992
2 67951 1 6992
2 67952 1 6992
2 67953 1 6992
2 67954 1 6992
2 67955 1 6992
2 67956 1 6992
2 67957 1 7001
2 67958 1 7001
2 67959 1 7007
2 67960 1 7007
2 67961 1 7007
2 67962 1 7007
2 67963 1 7007
2 67964 1 7007
2 67965 1 7009
2 67966 1 7009
2 67967 1 7009
2 67968 1 7009
2 67969 1 7010
2 67970 1 7010
2 67971 1 7011
2 67972 1 7011
2 67973 1 7023
2 67974 1 7023
2 67975 1 7023
2 67976 1 7028
2 67977 1 7028
2 67978 1 7029
2 67979 1 7029
2 67980 1 7029
2 67981 1 7029
2 67982 1 7030
2 67983 1 7030
2 67984 1 7030
2 67985 1 7031
2 67986 1 7031
2 67987 1 7031
2 67988 1 7031
2 67989 1 7031
2 67990 1 7032
2 67991 1 7032
2 67992 1 7032
2 67993 1 7032
2 67994 1 7032
2 67995 1 7032
2 67996 1 7041
2 67997 1 7041
2 67998 1 7043
2 67999 1 7043
2 68000 1 7043
2 68001 1 7043
2 68002 1 7044
2 68003 1 7044
2 68004 1 7055
2 68005 1 7055
2 68006 1 7057
2 68007 1 7057
2 68008 1 7058
2 68009 1 7058
2 68010 1 7059
2 68011 1 7059
2 68012 1 7060
2 68013 1 7060
2 68014 1 7079
2 68015 1 7079
2 68016 1 7079
2 68017 1 7079
2 68018 1 7080
2 68019 1 7080
2 68020 1 7080
2 68021 1 7080
2 68022 1 7080
2 68023 1 7081
2 68024 1 7081
2 68025 1 7094
2 68026 1 7094
2 68027 1 7096
2 68028 1 7096
2 68029 1 7097
2 68030 1 7097
2 68031 1 7097
2 68032 1 7098
2 68033 1 7098
2 68034 1 7098
2 68035 1 7098
2 68036 1 7106
2 68037 1 7106
2 68038 1 7109
2 68039 1 7109
2 68040 1 7109
2 68041 1 7109
2 68042 1 7112
2 68043 1 7112
2 68044 1 7129
2 68045 1 7129
2 68046 1 7130
2 68047 1 7130
2 68048 1 7134
2 68049 1 7134
2 68050 1 7136
2 68051 1 7136
2 68052 1 7149
2 68053 1 7149
2 68054 1 7161
2 68055 1 7161
2 68056 1 7162
2 68057 1 7162
2 68058 1 7162
2 68059 1 7162
2 68060 1 7163
2 68061 1 7163
2 68062 1 7171
2 68063 1 7171
2 68064 1 7171
2 68065 1 7171
2 68066 1 7171
2 68067 1 7172
2 68068 1 7172
2 68069 1 7172
2 68070 1 7172
2 68071 1 7172
2 68072 1 7173
2 68073 1 7173
2 68074 1 7177
2 68075 1 7177
2 68076 1 7177
2 68077 1 7177
2 68078 1 7177
2 68079 1 7177
2 68080 1 7177
2 68081 1 7185
2 68082 1 7185
2 68083 1 7185
2 68084 1 7185
2 68085 1 7185
2 68086 1 7192
2 68087 1 7192
2 68088 1 7205
2 68089 1 7205
2 68090 1 7221
2 68091 1 7221
2 68092 1 7221
2 68093 1 7221
2 68094 1 7241
2 68095 1 7241
2 68096 1 7241
2 68097 1 7241
2 68098 1 7241
2 68099 1 7241
2 68100 1 7249
2 68101 1 7249
2 68102 1 7249
2 68103 1 7250
2 68104 1 7250
2 68105 1 7250
2 68106 1 7252
2 68107 1 7252
2 68108 1 7254
2 68109 1 7254
2 68110 1 7257
2 68111 1 7257
2 68112 1 7257
2 68113 1 7257
2 68114 1 7257
2 68115 1 7258
2 68116 1 7258
2 68117 1 7258
2 68118 1 7258
2 68119 1 7258
2 68120 1 7258
2 68121 1 7258
2 68122 1 7258
2 68123 1 7259
2 68124 1 7259
2 68125 1 7259
2 68126 1 7259
2 68127 1 7261
2 68128 1 7261
2 68129 1 7277
2 68130 1 7277
2 68131 1 7277
2 68132 1 7290
2 68133 1 7290
2 68134 1 7290
2 68135 1 7291
2 68136 1 7291
2 68137 1 7291
2 68138 1 7291
2 68139 1 7291
2 68140 1 7291
2 68141 1 7291
2 68142 1 7291
2 68143 1 7291
2 68144 1 7291
2 68145 1 7291
2 68146 1 7296
2 68147 1 7296
2 68148 1 7296
2 68149 1 7297
2 68150 1 7297
2 68151 1 7305
2 68152 1 7305
2 68153 1 7306
2 68154 1 7306
2 68155 1 7306
2 68156 1 7306
2 68157 1 7308
2 68158 1 7308
2 68159 1 7309
2 68160 1 7309
2 68161 1 7316
2 68162 1 7316
2 68163 1 7317
2 68164 1 7317
2 68165 1 7317
2 68166 1 7317
2 68167 1 7345
2 68168 1 7345
2 68169 1 7346
2 68170 1 7346
2 68171 1 7346
2 68172 1 7358
2 68173 1 7358
2 68174 1 7364
2 68175 1 7364
2 68176 1 7364
2 68177 1 7364
2 68178 1 7364
2 68179 1 7364
2 68180 1 7364
2 68181 1 7364
2 68182 1 7364
2 68183 1 7366
2 68184 1 7366
2 68185 1 7366
2 68186 1 7366
2 68187 1 7366
2 68188 1 7366
2 68189 1 7366
2 68190 1 7366
2 68191 1 7366
2 68192 1 7366
2 68193 1 7366
2 68194 1 7366
2 68195 1 7366
2 68196 1 7366
2 68197 1 7366
2 68198 1 7366
2 68199 1 7368
2 68200 1 7368
2 68201 1 7373
2 68202 1 7373
2 68203 1 7395
2 68204 1 7395
2 68205 1 7395
2 68206 1 7395
2 68207 1 7395
2 68208 1 7395
2 68209 1 7395
2 68210 1 7395
2 68211 1 7395
2 68212 1 7395
2 68213 1 7395
2 68214 1 7396
2 68215 1 7396
2 68216 1 7396
2 68217 1 7396
2 68218 1 7396
2 68219 1 7396
2 68220 1 7396
2 68221 1 7396
2 68222 1 7396
2 68223 1 7396
2 68224 1 7396
2 68225 1 7397
2 68226 1 7397
2 68227 1 7397
2 68228 1 7397
2 68229 1 7397
2 68230 1 7397
2 68231 1 7397
2 68232 1 7397
2 68233 1 7397
2 68234 1 7397
2 68235 1 7397
2 68236 1 7397
2 68237 1 7397
2 68238 1 7397
2 68239 1 7397
2 68240 1 7397
2 68241 1 7397
2 68242 1 7397
2 68243 1 7397
2 68244 1 7397
2 68245 1 7397
2 68246 1 7397
2 68247 1 7397
2 68248 1 7397
2 68249 1 7397
2 68250 1 7397
2 68251 1 7397
2 68252 1 7397
2 68253 1 7397
2 68254 1 7397
2 68255 1 7397
2 68256 1 7397
2 68257 1 7397
2 68258 1 7397
2 68259 1 7397
2 68260 1 7397
2 68261 1 7397
2 68262 1 7397
2 68263 1 7397
2 68264 1 7397
2 68265 1 7397
2 68266 1 7397
2 68267 1 7397
2 68268 1 7397
2 68269 1 7397
2 68270 1 7397
2 68271 1 7397
2 68272 1 7397
2 68273 1 7397
2 68274 1 7398
2 68275 1 7398
2 68276 1 7398
2 68277 1 7399
2 68278 1 7399
2 68279 1 7399
2 68280 1 7399
2 68281 1 7403
2 68282 1 7403
2 68283 1 7404
2 68284 1 7404
2 68285 1 7404
2 68286 1 7404
2 68287 1 7408
2 68288 1 7408
2 68289 1 7409
2 68290 1 7409
2 68291 1 7409
2 68292 1 7409
2 68293 1 7409
2 68294 1 7409
2 68295 1 7409
2 68296 1 7409
2 68297 1 7409
2 68298 1 7410
2 68299 1 7410
2 68300 1 7413
2 68301 1 7413
2 68302 1 7419
2 68303 1 7419
2 68304 1 7419
2 68305 1 7419
2 68306 1 7419
2 68307 1 7419
2 68308 1 7419
2 68309 1 7419
2 68310 1 7419
2 68311 1 7419
2 68312 1 7419
2 68313 1 7419
2 68314 1 7419
2 68315 1 7419
2 68316 1 7419
2 68317 1 7427
2 68318 1 7427
2 68319 1 7427
2 68320 1 7427
2 68321 1 7427
2 68322 1 7427
2 68323 1 7427
2 68324 1 7427
2 68325 1 7428
2 68326 1 7428
2 68327 1 7428
2 68328 1 7436
2 68329 1 7436
2 68330 1 7436
2 68331 1 7436
2 68332 1 7436
2 68333 1 7436
2 68334 1 7436
2 68335 1 7437
2 68336 1 7437
2 68337 1 7437
2 68338 1 7444
2 68339 1 7444
2 68340 1 7444
2 68341 1 7444
2 68342 1 7444
2 68343 1 7444
2 68344 1 7444
2 68345 1 7444
2 68346 1 7444
2 68347 1 7444
2 68348 1 7444
2 68349 1 7444
2 68350 1 7444
2 68351 1 7444
2 68352 1 7445
2 68353 1 7445
2 68354 1 7453
2 68355 1 7453
2 68356 1 7453
2 68357 1 7453
2 68358 1 7453
2 68359 1 7453
2 68360 1 7474
2 68361 1 7474
2 68362 1 7475
2 68363 1 7475
2 68364 1 7475
2 68365 1 7475
2 68366 1 7475
2 68367 1 7477
2 68368 1 7477
2 68369 1 7477
2 68370 1 7477
2 68371 1 7478
2 68372 1 7478
2 68373 1 7479
2 68374 1 7479
2 68375 1 7509
2 68376 1 7509
2 68377 1 7509
2 68378 1 7509
2 68379 1 7509
2 68380 1 7509
2 68381 1 7509
2 68382 1 7509
2 68383 1 7509
2 68384 1 7509
2 68385 1 7509
2 68386 1 7509
2 68387 1 7509
2 68388 1 7509
2 68389 1 7509
2 68390 1 7509
2 68391 1 7509
2 68392 1 7509
2 68393 1 7509
2 68394 1 7509
2 68395 1 7509
2 68396 1 7509
2 68397 1 7509
2 68398 1 7509
2 68399 1 7509
2 68400 1 7509
2 68401 1 7509
2 68402 1 7509
2 68403 1 7509
2 68404 1 7509
2 68405 1 7509
2 68406 1 7509
2 68407 1 7509
2 68408 1 7509
2 68409 1 7510
2 68410 1 7510
2 68411 1 7511
2 68412 1 7511
2 68413 1 7511
2 68414 1 7515
2 68415 1 7515
2 68416 1 7520
2 68417 1 7520
2 68418 1 7527
2 68419 1 7527
2 68420 1 7536
2 68421 1 7536
2 68422 1 7537
2 68423 1 7537
2 68424 1 7538
2 68425 1 7538
2 68426 1 7539
2 68427 1 7539
2 68428 1 7539
2 68429 1 7539
2 68430 1 7539
2 68431 1 7539
2 68432 1 7552
2 68433 1 7552
2 68434 1 7553
2 68435 1 7553
2 68436 1 7553
2 68437 1 7553
2 68438 1 7554
2 68439 1 7554
2 68440 1 7554
2 68441 1 7554
2 68442 1 7563
2 68443 1 7563
2 68444 1 7563
2 68445 1 7563
2 68446 1 7579
2 68447 1 7579
2 68448 1 7579
2 68449 1 7579
2 68450 1 7579
2 68451 1 7579
2 68452 1 7579
2 68453 1 7579
2 68454 1 7579
2 68455 1 7579
2 68456 1 7579
2 68457 1 7579
2 68458 1 7579
2 68459 1 7579
2 68460 1 7579
2 68461 1 7579
2 68462 1 7579
2 68463 1 7579
2 68464 1 7579
2 68465 1 7579
2 68466 1 7579
2 68467 1 7579
2 68468 1 7579
2 68469 1 7579
2 68470 1 7579
2 68471 1 7579
2 68472 1 7580
2 68473 1 7580
2 68474 1 7580
2 68475 1 7581
2 68476 1 7581
2 68477 1 7581
2 68478 1 7581
2 68479 1 7581
2 68480 1 7581
2 68481 1 7581
2 68482 1 7582
2 68483 1 7582
2 68484 1 7582
2 68485 1 7584
2 68486 1 7584
2 68487 1 7585
2 68488 1 7585
2 68489 1 7585
2 68490 1 7585
2 68491 1 7586
2 68492 1 7586
2 68493 1 7586
2 68494 1 7586
2 68495 1 7586
2 68496 1 7586
2 68497 1 7586
2 68498 1 7586
2 68499 1 7586
2 68500 1 7586
2 68501 1 7586
2 68502 1 7586
2 68503 1 7586
2 68504 1 7586
2 68505 1 7586
2 68506 1 7587
2 68507 1 7587
2 68508 1 7588
2 68509 1 7588
2 68510 1 7588
2 68511 1 7588
2 68512 1 7588
2 68513 1 7588
2 68514 1 7588
2 68515 1 7589
2 68516 1 7589
2 68517 1 7597
2 68518 1 7597
2 68519 1 7597
2 68520 1 7597
2 68521 1 7597
2 68522 1 7597
2 68523 1 7597
2 68524 1 7597
2 68525 1 7597
2 68526 1 7597
2 68527 1 7597
2 68528 1 7597
2 68529 1 7597
2 68530 1 7597
2 68531 1 7597
2 68532 1 7598
2 68533 1 7598
2 68534 1 7598
2 68535 1 7599
2 68536 1 7599
2 68537 1 7614
2 68538 1 7614
2 68539 1 7615
2 68540 1 7615
2 68541 1 7628
2 68542 1 7628
2 68543 1 7628
2 68544 1 7628
2 68545 1 7628
2 68546 1 7628
2 68547 1 7628
2 68548 1 7628
2 68549 1 7628
2 68550 1 7628
2 68551 1 7628
2 68552 1 7628
2 68553 1 7628
2 68554 1 7629
2 68555 1 7629
2 68556 1 7629
2 68557 1 7629
2 68558 1 7631
2 68559 1 7631
2 68560 1 7635
2 68561 1 7635
2 68562 1 7642
2 68563 1 7642
2 68564 1 7643
2 68565 1 7643
2 68566 1 7643
2 68567 1 7643
2 68568 1 7644
2 68569 1 7644
2 68570 1 7644
2 68571 1 7644
2 68572 1 7644
2 68573 1 7644
2 68574 1 7644
2 68575 1 7644
2 68576 1 7644
2 68577 1 7644
2 68578 1 7644
2 68579 1 7644
2 68580 1 7644
2 68581 1 7644
2 68582 1 7644
2 68583 1 7644
2 68584 1 7644
2 68585 1 7644
2 68586 1 7644
2 68587 1 7644
2 68588 1 7644
2 68589 1 7644
2 68590 1 7644
2 68591 1 7644
2 68592 1 7644
2 68593 1 7644
2 68594 1 7644
2 68595 1 7644
2 68596 1 7644
2 68597 1 7644
2 68598 1 7644
2 68599 1 7644
2 68600 1 7645
2 68601 1 7645
2 68602 1 7645
2 68603 1 7645
2 68604 1 7645
2 68605 1 7645
2 68606 1 7645
2 68607 1 7645
2 68608 1 7645
2 68609 1 7645
2 68610 1 7646
2 68611 1 7646
2 68612 1 7646
2 68613 1 7646
2 68614 1 7646
2 68615 1 7646
2 68616 1 7646
2 68617 1 7646
2 68618 1 7647
2 68619 1 7647
2 68620 1 7647
2 68621 1 7647
2 68622 1 7654
2 68623 1 7654
2 68624 1 7654
2 68625 1 7655
2 68626 1 7655
2 68627 1 7662
2 68628 1 7662
2 68629 1 7662
2 68630 1 7662
2 68631 1 7662
2 68632 1 7663
2 68633 1 7663
2 68634 1 7672
2 68635 1 7672
2 68636 1 7674
2 68637 1 7674
2 68638 1 7674
2 68639 1 7688
2 68640 1 7688
2 68641 1 7688
2 68642 1 7688
2 68643 1 7688
2 68644 1 7689
2 68645 1 7689
2 68646 1 7690
2 68647 1 7690
2 68648 1 7708
2 68649 1 7708
2 68650 1 7711
2 68651 1 7711
2 68652 1 7719
2 68653 1 7719
2 68654 1 7719
2 68655 1 7719
2 68656 1 7726
2 68657 1 7726
2 68658 1 7726
2 68659 1 7726
2 68660 1 7726
2 68661 1 7726
2 68662 1 7726
2 68663 1 7726
2 68664 1 7726
2 68665 1 7726
2 68666 1 7726
2 68667 1 7726
2 68668 1 7726
2 68669 1 7726
2 68670 1 7726
2 68671 1 7727
2 68672 1 7727
2 68673 1 7729
2 68674 1 7729
2 68675 1 7734
2 68676 1 7734
2 68677 1 7735
2 68678 1 7735
2 68679 1 7735
2 68680 1 7735
2 68681 1 7736
2 68682 1 7736
2 68683 1 7736
2 68684 1 7736
2 68685 1 7736
2 68686 1 7740
2 68687 1 7740
2 68688 1 7740
2 68689 1 7740
2 68690 1 7740
2 68691 1 7740
2 68692 1 7740
2 68693 1 7740
2 68694 1 7740
2 68695 1 7740
2 68696 1 7740
2 68697 1 7740
2 68698 1 7740
2 68699 1 7740
2 68700 1 7740
2 68701 1 7740
2 68702 1 7740
2 68703 1 7740
2 68704 1 7740
2 68705 1 7740
2 68706 1 7740
2 68707 1 7742
2 68708 1 7742
2 68709 1 7742
2 68710 1 7742
2 68711 1 7742
2 68712 1 7755
2 68713 1 7755
2 68714 1 7755
2 68715 1 7755
2 68716 1 7755
2 68717 1 7755
2 68718 1 7755
2 68719 1 7755
2 68720 1 7756
2 68721 1 7756
2 68722 1 7756
2 68723 1 7758
2 68724 1 7758
2 68725 1 7758
2 68726 1 7761
2 68727 1 7761
2 68728 1 7773
2 68729 1 7773
2 68730 1 7773
2 68731 1 7773
2 68732 1 7774
2 68733 1 7774
2 68734 1 7775
2 68735 1 7775
2 68736 1 7775
2 68737 1 7777
2 68738 1 7777
2 68739 1 7777
2 68740 1 7778
2 68741 1 7778
2 68742 1 7778
2 68743 1 7786
2 68744 1 7786
2 68745 1 7786
2 68746 1 7786
2 68747 1 7786
2 68748 1 7786
2 68749 1 7786
2 68750 1 7786
2 68751 1 7786
2 68752 1 7786
2 68753 1 7786
2 68754 1 7786
2 68755 1 7786
2 68756 1 7786
2 68757 1 7788
2 68758 1 7788
2 68759 1 7788
2 68760 1 7789
2 68761 1 7789
2 68762 1 7789
2 68763 1 7789
2 68764 1 7789
2 68765 1 7792
2 68766 1 7792
2 68767 1 7792
2 68768 1 7792
2 68769 1 7792
2 68770 1 7792
2 68771 1 7792
2 68772 1 7792
2 68773 1 7792
2 68774 1 7792
2 68775 1 7792
2 68776 1 7792
2 68777 1 7793
2 68778 1 7793
2 68779 1 7794
2 68780 1 7794
2 68781 1 7794
2 68782 1 7810
2 68783 1 7810
2 68784 1 7810
2 68785 1 7811
2 68786 1 7811
2 68787 1 7812
2 68788 1 7812
2 68789 1 7818
2 68790 1 7818
2 68791 1 7818
2 68792 1 7819
2 68793 1 7819
2 68794 1 7819
2 68795 1 7819
2 68796 1 7819
2 68797 1 7826
2 68798 1 7826
2 68799 1 7826
2 68800 1 7826
2 68801 1 7826
2 68802 1 7826
2 68803 1 7826
2 68804 1 7826
2 68805 1 7826
2 68806 1 7826
2 68807 1 7826
2 68808 1 7826
2 68809 1 7826
2 68810 1 7826
2 68811 1 7826
2 68812 1 7826
2 68813 1 7826
2 68814 1 7826
2 68815 1 7827
2 68816 1 7827
2 68817 1 7827
2 68818 1 7828
2 68819 1 7828
2 68820 1 7828
2 68821 1 7828
2 68822 1 7828
2 68823 1 7828
2 68824 1 7828
2 68825 1 7828
2 68826 1 7828
2 68827 1 7828
2 68828 1 7828
2 68829 1 7828
2 68830 1 7828
2 68831 1 7828
2 68832 1 7828
2 68833 1 7828
2 68834 1 7828
2 68835 1 7828
2 68836 1 7828
2 68837 1 7829
2 68838 1 7829
2 68839 1 7829
2 68840 1 7829
2 68841 1 7830
2 68842 1 7830
2 68843 1 7830
2 68844 1 7830
2 68845 1 7830
2 68846 1 7831
2 68847 1 7831
2 68848 1 7832
2 68849 1 7832
2 68850 1 7832
2 68851 1 7833
2 68852 1 7833
2 68853 1 7846
2 68854 1 7846
2 68855 1 7846
2 68856 1 7847
2 68857 1 7847
2 68858 1 7847
2 68859 1 7847
2 68860 1 7847
2 68861 1 7847
2 68862 1 7847
2 68863 1 7847
2 68864 1 7848
2 68865 1 7848
2 68866 1 7850
2 68867 1 7850
2 68868 1 7850
2 68869 1 7856
2 68870 1 7856
2 68871 1 7856
2 68872 1 7856
2 68873 1 7856
2 68874 1 7856
2 68875 1 7856
2 68876 1 7856
2 68877 1 7856
2 68878 1 7856
2 68879 1 7856
2 68880 1 7856
2 68881 1 7856
2 68882 1 7856
2 68883 1 7856
2 68884 1 7857
2 68885 1 7857
2 68886 1 7857
2 68887 1 7857
2 68888 1 7857
2 68889 1 7865
2 68890 1 7865
2 68891 1 7865
2 68892 1 7865
2 68893 1 7865
2 68894 1 7865
2 68895 1 7865
2 68896 1 7865
2 68897 1 7865
2 68898 1 7865
2 68899 1 7865
2 68900 1 7865
2 68901 1 7865
2 68902 1 7865
2 68903 1 7865
2 68904 1 7865
2 68905 1 7865
2 68906 1 7865
2 68907 1 7865
2 68908 1 7866
2 68909 1 7866
2 68910 1 7879
2 68911 1 7879
2 68912 1 7880
2 68913 1 7880
2 68914 1 7886
2 68915 1 7886
2 68916 1 7886
2 68917 1 7886
2 68918 1 7886
2 68919 1 7886
2 68920 1 7886
2 68921 1 7886
2 68922 1 7886
2 68923 1 7886
2 68924 1 7886
2 68925 1 7886
2 68926 1 7886
2 68927 1 7886
2 68928 1 7886
2 68929 1 7886
2 68930 1 7886
2 68931 1 7886
2 68932 1 7886
2 68933 1 7886
2 68934 1 7886
2 68935 1 7886
2 68936 1 7886
2 68937 1 7886
2 68938 1 7886
2 68939 1 7886
2 68940 1 7888
2 68941 1 7888
2 68942 1 7888
2 68943 1 7893
2 68944 1 7893
2 68945 1 7893
2 68946 1 7893
2 68947 1 7893
2 68948 1 7893
2 68949 1 7902
2 68950 1 7902
2 68951 1 7902
2 68952 1 7902
2 68953 1 7902
2 68954 1 7902
2 68955 1 7902
2 68956 1 7902
2 68957 1 7903
2 68958 1 7903
2 68959 1 7903
2 68960 1 7903
2 68961 1 7903
2 68962 1 7903
2 68963 1 7903
2 68964 1 7903
2 68965 1 7903
2 68966 1 7904
2 68967 1 7904
2 68968 1 7904
2 68969 1 7905
2 68970 1 7905
2 68971 1 7908
2 68972 1 7908
2 68973 1 7908
2 68974 1 7908
2 68975 1 7908
2 68976 1 7908
2 68977 1 7908
2 68978 1 7908
2 68979 1 7908
2 68980 1 7908
2 68981 1 7908
2 68982 1 7909
2 68983 1 7909
2 68984 1 7909
2 68985 1 7909
2 68986 1 7909
2 68987 1 7909
2 68988 1 7910
2 68989 1 7910
2 68990 1 7912
2 68991 1 7912
2 68992 1 7912
2 68993 1 7913
2 68994 1 7913
2 68995 1 7913
2 68996 1 7913
2 68997 1 7913
2 68998 1 7913
2 68999 1 7914
2 69000 1 7914
2 69001 1 7914
2 69002 1 7914
2 69003 1 7914
2 69004 1 7926
2 69005 1 7926
2 69006 1 7926
2 69007 1 7930
2 69008 1 7930
2 69009 1 7930
2 69010 1 7932
2 69011 1 7932
2 69012 1 7946
2 69013 1 7946
2 69014 1 7946
2 69015 1 7946
2 69016 1 7946
2 69017 1 7946
2 69018 1 7946
2 69019 1 7946
2 69020 1 7949
2 69021 1 7949
2 69022 1 7949
2 69023 1 7949
2 69024 1 7949
2 69025 1 7949
2 69026 1 7949
2 69027 1 7949
2 69028 1 7949
2 69029 1 7949
2 69030 1 7949
2 69031 1 7950
2 69032 1 7950
2 69033 1 7950
2 69034 1 7950
2 69035 1 7958
2 69036 1 7958
2 69037 1 7959
2 69038 1 7959
2 69039 1 7959
2 69040 1 7959
2 69041 1 7962
2 69042 1 7962
2 69043 1 7962
2 69044 1 7962
2 69045 1 7962
2 69046 1 7962
2 69047 1 7962
2 69048 1 7970
2 69049 1 7970
2 69050 1 7970
2 69051 1 7970
2 69052 1 7970
2 69053 1 7971
2 69054 1 7971
2 69055 1 7971
2 69056 1 7972
2 69057 1 7972
2 69058 1 7972
2 69059 1 7975
2 69060 1 7975
2 69061 1 7976
2 69062 1 7976
2 69063 1 7978
2 69064 1 7978
2 69065 1 7993
2 69066 1 7993
2 69067 1 7993
2 69068 1 7993
2 69069 1 7994
2 69070 1 7994
2 69071 1 7994
2 69072 1 7996
2 69073 1 7996
2 69074 1 7996
2 69075 1 7996
2 69076 1 7996
2 69077 1 7996
2 69078 1 7996
2 69079 1 7996
2 69080 1 7996
2 69081 1 7996
2 69082 1 7996
2 69083 1 7996
2 69084 1 7996
2 69085 1 7996
2 69086 1 7996
2 69087 1 7996
2 69088 1 7996
2 69089 1 7996
2 69090 1 7996
2 69091 1 7996
2 69092 1 7996
2 69093 1 7996
2 69094 1 7996
2 69095 1 8000
2 69096 1 8000
2 69097 1 8012
2 69098 1 8012
2 69099 1 8012
2 69100 1 8012
2 69101 1 8012
2 69102 1 8012
2 69103 1 8012
2 69104 1 8012
2 69105 1 8012
2 69106 1 8014
2 69107 1 8014
2 69108 1 8014
2 69109 1 8014
2 69110 1 8014
2 69111 1 8014
2 69112 1 8015
2 69113 1 8015
2 69114 1 8015
2 69115 1 8015
2 69116 1 8022
2 69117 1 8022
2 69118 1 8022
2 69119 1 8022
2 69120 1 8023
2 69121 1 8023
2 69122 1 8024
2 69123 1 8024
2 69124 1 8024
2 69125 1 8024
2 69126 1 8024
2 69127 1 8024
2 69128 1 8025
2 69129 1 8025
2 69130 1 8027
2 69131 1 8027
2 69132 1 8031
2 69133 1 8031
2 69134 1 8039
2 69135 1 8039
2 69136 1 8059
2 69137 1 8059
2 69138 1 8067
2 69139 1 8067
2 69140 1 8067
2 69141 1 8067
2 69142 1 8067
2 69143 1 8067
2 69144 1 8068
2 69145 1 8068
2 69146 1 8068
2 69147 1 8068
2 69148 1 8068
2 69149 1 8068
2 69150 1 8068
2 69151 1 8068
2 69152 1 8069
2 69153 1 8069
2 69154 1 8076
2 69155 1 8076
2 69156 1 8076
2 69157 1 8076
2 69158 1 8077
2 69159 1 8077
2 69160 1 8077
2 69161 1 8079
2 69162 1 8079
2 69163 1 8081
2 69164 1 8081
2 69165 1 8090
2 69166 1 8090
2 69167 1 8090
2 69168 1 8090
2 69169 1 8090
2 69170 1 8090
2 69171 1 8091
2 69172 1 8091
2 69173 1 8091
2 69174 1 8091
2 69175 1 8091
2 69176 1 8091
2 69177 1 8091
2 69178 1 8091
2 69179 1 8092
2 69180 1 8092
2 69181 1 8092
2 69182 1 8092
2 69183 1 8095
2 69184 1 8095
2 69185 1 8095
2 69186 1 8095
2 69187 1 8095
2 69188 1 8095
2 69189 1 8095
2 69190 1 8097
2 69191 1 8097
2 69192 1 8097
2 69193 1 8098
2 69194 1 8098
2 69195 1 8099
2 69196 1 8099
2 69197 1 8099
2 69198 1 8104
2 69199 1 8104
2 69200 1 8104
2 69201 1 8104
2 69202 1 8104
2 69203 1 8104
2 69204 1 8107
2 69205 1 8107
2 69206 1 8107
2 69207 1 8107
2 69208 1 8107
2 69209 1 8108
2 69210 1 8108
2 69211 1 8109
2 69212 1 8109
2 69213 1 8109
2 69214 1 8109
2 69215 1 8109
2 69216 1 8109
2 69217 1 8118
2 69218 1 8118
2 69219 1 8118
2 69220 1 8121
2 69221 1 8121
2 69222 1 8128
2 69223 1 8128
2 69224 1 8136
2 69225 1 8136
2 69226 1 8147
2 69227 1 8147
2 69228 1 8147
2 69229 1 8148
2 69230 1 8148
2 69231 1 8149
2 69232 1 8149
2 69233 1 8152
2 69234 1 8152
2 69235 1 8152
2 69236 1 8163
2 69237 1 8163
2 69238 1 8163
2 69239 1 8164
2 69240 1 8164
2 69241 1 8164
2 69242 1 8164
2 69243 1 8164
2 69244 1 8164
2 69245 1 8164
2 69246 1 8165
2 69247 1 8165
2 69248 1 8169
2 69249 1 8169
2 69250 1 8170
2 69251 1 8170
2 69252 1 8170
2 69253 1 8172
2 69254 1 8172
2 69255 1 8172
2 69256 1 8172
2 69257 1 8179
2 69258 1 8179
2 69259 1 8201
2 69260 1 8201
2 69261 1 8201
2 69262 1 8201
2 69263 1 8201
2 69264 1 8201
2 69265 1 8201
2 69266 1 8201
2 69267 1 8201
2 69268 1 8201
2 69269 1 8201
2 69270 1 8202
2 69271 1 8202
2 69272 1 8202
2 69273 1 8202
2 69274 1 8202
2 69275 1 8202
2 69276 1 8202
2 69277 1 8202
2 69278 1 8204
2 69279 1 8204
2 69280 1 8229
2 69281 1 8229
2 69282 1 8230
2 69283 1 8230
2 69284 1 8243
2 69285 1 8243
2 69286 1 8243
2 69287 1 8243
2 69288 1 8243
2 69289 1 8243
2 69290 1 8243
2 69291 1 8243
2 69292 1 8244
2 69293 1 8244
2 69294 1 8244
2 69295 1 8244
2 69296 1 8245
2 69297 1 8245
2 69298 1 8252
2 69299 1 8252
2 69300 1 8252
2 69301 1 8252
2 69302 1 8252
2 69303 1 8252
2 69304 1 8252
2 69305 1 8253
2 69306 1 8253
2 69307 1 8253
2 69308 1 8253
2 69309 1 8253
2 69310 1 8253
2 69311 1 8253
2 69312 1 8253
2 69313 1 8253
2 69314 1 8253
2 69315 1 8254
2 69316 1 8254
2 69317 1 8254
2 69318 1 8255
2 69319 1 8255
2 69320 1 8255
2 69321 1 8255
2 69322 1 8255
2 69323 1 8257
2 69324 1 8257
2 69325 1 8257
2 69326 1 8257
2 69327 1 8264
2 69328 1 8264
2 69329 1 8265
2 69330 1 8265
2 69331 1 8266
2 69332 1 8266
2 69333 1 8266
2 69334 1 8266
2 69335 1 8266
2 69336 1 8266
2 69337 1 8269
2 69338 1 8269
2 69339 1 8270
2 69340 1 8270
2 69341 1 8270
2 69342 1 8273
2 69343 1 8273
2 69344 1 8273
2 69345 1 8273
2 69346 1 8273
2 69347 1 8273
2 69348 1 8273
2 69349 1 8273
2 69350 1 8273
2 69351 1 8273
2 69352 1 8273
2 69353 1 8273
2 69354 1 8273
2 69355 1 8273
2 69356 1 8273
2 69357 1 8273
2 69358 1 8273
2 69359 1 8274
2 69360 1 8274
2 69361 1 8274
2 69362 1 8289
2 69363 1 8289
2 69364 1 8289
2 69365 1 8289
2 69366 1 8289
2 69367 1 8289
2 69368 1 8296
2 69369 1 8296
2 69370 1 8314
2 69371 1 8314
2 69372 1 8314
2 69373 1 8315
2 69374 1 8315
2 69375 1 8326
2 69376 1 8326
2 69377 1 8326
2 69378 1 8326
2 69379 1 8326
2 69380 1 8326
2 69381 1 8326
2 69382 1 8327
2 69383 1 8327
2 69384 1 8328
2 69385 1 8328
2 69386 1 8328
2 69387 1 8330
2 69388 1 8330
2 69389 1 8330
2 69390 1 8345
2 69391 1 8345
2 69392 1 8346
2 69393 1 8346
2 69394 1 8346
2 69395 1 8346
2 69396 1 8346
2 69397 1 8347
2 69398 1 8347
2 69399 1 8350
2 69400 1 8350
2 69401 1 8350
2 69402 1 8358
2 69403 1 8358
2 69404 1 8367
2 69405 1 8367
2 69406 1 8367
2 69407 1 8367
2 69408 1 8367
2 69409 1 8367
2 69410 1 8367
2 69411 1 8367
2 69412 1 8367
2 69413 1 8368
2 69414 1 8368
2 69415 1 8368
2 69416 1 8368
2 69417 1 8368
2 69418 1 8369
2 69419 1 8369
2 69420 1 8369
2 69421 1 8369
2 69422 1 8369
2 69423 1 8377
2 69424 1 8377
2 69425 1 8377
2 69426 1 8377
2 69427 1 8377
2 69428 1 8377
2 69429 1 8377
2 69430 1 8377
2 69431 1 8378
2 69432 1 8378
2 69433 1 8378
2 69434 1 8378
2 69435 1 8378
2 69436 1 8382
2 69437 1 8382
2 69438 1 8382
2 69439 1 8383
2 69440 1 8383
2 69441 1 8383
2 69442 1 8393
2 69443 1 8393
2 69444 1 8393
2 69445 1 8393
2 69446 1 8393
2 69447 1 8393
2 69448 1 8393
2 69449 1 8403
2 69450 1 8403
2 69451 1 8411
2 69452 1 8411
2 69453 1 8411
2 69454 1 8411
2 69455 1 8411
2 69456 1 8411
2 69457 1 8411
2 69458 1 8418
2 69459 1 8418
2 69460 1 8418
2 69461 1 8418
2 69462 1 8418
2 69463 1 8418
2 69464 1 8418
2 69465 1 8418
2 69466 1 8418
2 69467 1 8418
2 69468 1 8418
2 69469 1 8418
2 69470 1 8419
2 69471 1 8419
2 69472 1 8419
2 69473 1 8427
2 69474 1 8427
2 69475 1 8434
2 69476 1 8434
2 69477 1 8434
2 69478 1 8434
2 69479 1 8434
2 69480 1 8435
2 69481 1 8435
2 69482 1 8448
2 69483 1 8448
2 69484 1 8449
2 69485 1 8449
2 69486 1 8449
2 69487 1 8449
2 69488 1 8453
2 69489 1 8453
2 69490 1 8469
2 69491 1 8469
2 69492 1 8473
2 69493 1 8473
2 69494 1 8475
2 69495 1 8475
2 69496 1 8484
2 69497 1 8484
2 69498 1 8484
2 69499 1 8484
2 69500 1 8484
2 69501 1 8485
2 69502 1 8485
2 69503 1 8512
2 69504 1 8512
2 69505 1 8512
2 69506 1 8512
2 69507 1 8522
2 69508 1 8522
2 69509 1 8525
2 69510 1 8525
2 69511 1 8525
2 69512 1 8525
2 69513 1 8525
2 69514 1 8528
2 69515 1 8528
2 69516 1 8529
2 69517 1 8529
2 69518 1 8529
2 69519 1 8529
2 69520 1 8529
2 69521 1 8529
2 69522 1 8529
2 69523 1 8529
2 69524 1 8529
2 69525 1 8529
2 69526 1 8529
2 69527 1 8529
2 69528 1 8529
2 69529 1 8529
2 69530 1 8529
2 69531 1 8529
2 69532 1 8529
2 69533 1 8529
2 69534 1 8529
2 69535 1 8529
2 69536 1 8529
2 69537 1 8529
2 69538 1 8529
2 69539 1 8529
2 69540 1 8529
2 69541 1 8529
2 69542 1 8529
2 69543 1 8529
2 69544 1 8529
2 69545 1 8529
2 69546 1 8529
2 69547 1 8529
2 69548 1 8529
2 69549 1 8530
2 69550 1 8530
2 69551 1 8530
2 69552 1 8530
2 69553 1 8530
2 69554 1 8530
2 69555 1 8530
2 69556 1 8530
2 69557 1 8530
2 69558 1 8530
2 69559 1 8530
2 69560 1 8530
2 69561 1 8530
2 69562 1 8530
2 69563 1 8530
2 69564 1 8530
2 69565 1 8530
2 69566 1 8530
2 69567 1 8530
2 69568 1 8530
2 69569 1 8530
2 69570 1 8530
2 69571 1 8530
2 69572 1 8530
2 69573 1 8530
2 69574 1 8530
2 69575 1 8530
2 69576 1 8530
2 69577 1 8530
2 69578 1 8530
2 69579 1 8530
2 69580 1 8531
2 69581 1 8531
2 69582 1 8543
2 69583 1 8543
2 69584 1 8543
2 69585 1 8543
2 69586 1 8543
2 69587 1 8543
2 69588 1 8564
2 69589 1 8564
2 69590 1 8565
2 69591 1 8565
2 69592 1 8573
2 69593 1 8573
2 69594 1 8573
2 69595 1 8573
2 69596 1 8573
2 69597 1 8573
2 69598 1 8573
2 69599 1 8573
2 69600 1 8573
2 69601 1 8573
2 69602 1 8575
2 69603 1 8575
2 69604 1 8575
2 69605 1 8575
2 69606 1 8575
2 69607 1 8577
2 69608 1 8577
2 69609 1 8582
2 69610 1 8582
2 69611 1 8582
2 69612 1 8582
2 69613 1 8582
2 69614 1 8582
2 69615 1 8582
2 69616 1 8582
2 69617 1 8582
2 69618 1 8582
2 69619 1 8582
2 69620 1 8582
2 69621 1 8582
2 69622 1 8582
2 69623 1 8582
2 69624 1 8582
2 69625 1 8582
2 69626 1 8582
2 69627 1 8582
2 69628 1 8582
2 69629 1 8582
2 69630 1 8582
2 69631 1 8582
2 69632 1 8582
2 69633 1 8582
2 69634 1 8582
2 69635 1 8582
2 69636 1 8582
2 69637 1 8582
2 69638 1 8582
2 69639 1 8582
2 69640 1 8583
2 69641 1 8583
2 69642 1 8583
2 69643 1 8583
2 69644 1 8583
2 69645 1 8583
2 69646 1 8583
2 69647 1 8583
2 69648 1 8583
2 69649 1 8583
2 69650 1 8583
2 69651 1 8583
2 69652 1 8583
2 69653 1 8583
2 69654 1 8583
2 69655 1 8583
2 69656 1 8583
2 69657 1 8584
2 69658 1 8584
2 69659 1 8585
2 69660 1 8585
2 69661 1 8594
2 69662 1 8594
2 69663 1 8594
2 69664 1 8594
2 69665 1 8595
2 69666 1 8595
2 69667 1 8595
2 69668 1 8595
2 69669 1 8596
2 69670 1 8596
2 69671 1 8596
2 69672 1 8613
2 69673 1 8613
2 69674 1 8614
2 69675 1 8614
2 69676 1 8614
2 69677 1 8616
2 69678 1 8616
2 69679 1 8625
2 69680 1 8625
2 69681 1 8633
2 69682 1 8633
2 69683 1 8634
2 69684 1 8634
2 69685 1 8634
2 69686 1 8635
2 69687 1 8635
2 69688 1 8635
2 69689 1 8640
2 69690 1 8640
2 69691 1 8660
2 69692 1 8660
2 69693 1 8660
2 69694 1 8660
2 69695 1 8660
2 69696 1 8660
2 69697 1 8660
2 69698 1 8660
2 69699 1 8661
2 69700 1 8661
2 69701 1 8663
2 69702 1 8663
2 69703 1 8663
2 69704 1 8663
2 69705 1 8663
2 69706 1 8665
2 69707 1 8665
2 69708 1 8666
2 69709 1 8666
2 69710 1 8666
2 69711 1 8666
2 69712 1 8666
2 69713 1 8666
2 69714 1 8666
2 69715 1 8667
2 69716 1 8667
2 69717 1 8673
2 69718 1 8673
2 69719 1 8680
2 69720 1 8680
2 69721 1 8680
2 69722 1 8680
2 69723 1 8680
2 69724 1 8681
2 69725 1 8681
2 69726 1 8694
2 69727 1 8694
2 69728 1 8707
2 69729 1 8707
2 69730 1 8725
2 69731 1 8725
2 69732 1 8725
2 69733 1 8725
2 69734 1 8734
2 69735 1 8734
2 69736 1 8735
2 69737 1 8735
2 69738 1 8739
2 69739 1 8739
2 69740 1 8743
2 69741 1 8743
2 69742 1 8743
2 69743 1 8743
2 69744 1 8755
2 69745 1 8755
2 69746 1 8755
2 69747 1 8755
2 69748 1 8756
2 69749 1 8756
2 69750 1 8756
2 69751 1 8779
2 69752 1 8779
2 69753 1 8779
2 69754 1 8780
2 69755 1 8780
2 69756 1 8780
2 69757 1 8780
2 69758 1 8781
2 69759 1 8781
2 69760 1 8782
2 69761 1 8782
2 69762 1 8802
2 69763 1 8802
2 69764 1 8802
2 69765 1 8802
2 69766 1 8802
2 69767 1 8803
2 69768 1 8803
2 69769 1 8803
2 69770 1 8804
2 69771 1 8804
2 69772 1 8810
2 69773 1 8810
2 69774 1 8810
2 69775 1 8813
2 69776 1 8813
2 69777 1 8815
2 69778 1 8815
2 69779 1 8823
2 69780 1 8823
2 69781 1 8840
2 69782 1 8840
2 69783 1 8840
2 69784 1 8851
2 69785 1 8851
2 69786 1 8851
2 69787 1 8851
2 69788 1 8851
2 69789 1 8851
2 69790 1 8851
2 69791 1 8851
2 69792 1 8851
2 69793 1 8851
2 69794 1 8851
2 69795 1 8851
2 69796 1 8851
2 69797 1 8851
2 69798 1 8851
2 69799 1 8851
2 69800 1 8851
2 69801 1 8851
2 69802 1 8851
2 69803 1 8851
2 69804 1 8851
2 69805 1 8851
2 69806 1 8851
2 69807 1 8851
2 69808 1 8851
2 69809 1 8851
2 69810 1 8851
2 69811 1 8851
2 69812 1 8860
2 69813 1 8860
2 69814 1 8860
2 69815 1 8860
2 69816 1 8860
2 69817 1 8862
2 69818 1 8862
2 69819 1 8866
2 69820 1 8866
2 69821 1 8866
2 69822 1 8867
2 69823 1 8867
2 69824 1 8867
2 69825 1 8867
2 69826 1 8867
2 69827 1 8869
2 69828 1 8869
2 69829 1 8870
2 69830 1 8870
2 69831 1 8870
2 69832 1 8871
2 69833 1 8871
2 69834 1 8888
2 69835 1 8888
2 69836 1 8892
2 69837 1 8892
2 69838 1 8915
2 69839 1 8915
2 69840 1 8915
2 69841 1 8915
2 69842 1 8916
2 69843 1 8916
2 69844 1 8916
2 69845 1 8918
2 69846 1 8918
2 69847 1 8918
2 69848 1 8918
2 69849 1 8924
2 69850 1 8924
2 69851 1 8933
2 69852 1 8933
2 69853 1 8933
2 69854 1 8934
2 69855 1 8934
2 69856 1 8935
2 69857 1 8935
2 69858 1 8939
2 69859 1 8939
2 69860 1 8939
2 69861 1 8939
2 69862 1 8939
2 69863 1 8939
2 69864 1 8940
2 69865 1 8940
2 69866 1 8949
2 69867 1 8949
2 69868 1 8950
2 69869 1 8950
2 69870 1 8951
2 69871 1 8951
2 69872 1 8951
2 69873 1 8951
2 69874 1 8951
2 69875 1 8952
2 69876 1 8952
2 69877 1 8952
2 69878 1 8952
2 69879 1 8952
2 69880 1 8952
2 69881 1 8952
2 69882 1 8952
2 69883 1 8952
2 69884 1 8952
2 69885 1 8952
2 69886 1 8952
2 69887 1 8952
2 69888 1 8952
2 69889 1 8952
2 69890 1 8952
2 69891 1 8952
2 69892 1 8953
2 69893 1 8953
2 69894 1 8961
2 69895 1 8961
2 69896 1 8961
2 69897 1 8961
2 69898 1 8964
2 69899 1 8964
2 69900 1 8964
2 69901 1 8964
2 69902 1 8964
2 69903 1 8965
2 69904 1 8965
2 69905 1 8967
2 69906 1 8967
2 69907 1 8967
2 69908 1 8967
2 69909 1 8967
2 69910 1 8967
2 69911 1 8967
2 69912 1 8967
2 69913 1 8967
2 69914 1 8967
2 69915 1 8967
2 69916 1 8968
2 69917 1 8968
2 69918 1 8973
2 69919 1 8973
2 69920 1 8973
2 69921 1 8981
2 69922 1 8981
2 69923 1 8981
2 69924 1 8993
2 69925 1 8993
2 69926 1 8993
2 69927 1 8993
2 69928 1 9000
2 69929 1 9000
2 69930 1 9000
2 69931 1 9000
2 69932 1 9000
2 69933 1 9000
2 69934 1 9000
2 69935 1 9008
2 69936 1 9008
2 69937 1 9009
2 69938 1 9009
2 69939 1 9009
2 69940 1 9009
2 69941 1 9009
2 69942 1 9009
2 69943 1 9009
2 69944 1 9009
2 69945 1 9009
2 69946 1 9009
2 69947 1 9009
2 69948 1 9010
2 69949 1 9010
2 69950 1 9030
2 69951 1 9030
2 69952 1 9030
2 69953 1 9030
2 69954 1 9030
2 69955 1 9030
2 69956 1 9031
2 69957 1 9031
2 69958 1 9032
2 69959 1 9032
2 69960 1 9032
2 69961 1 9048
2 69962 1 9048
2 69963 1 9048
2 69964 1 9048
2 69965 1 9048
2 69966 1 9048
2 69967 1 9048
2 69968 1 9048
2 69969 1 9048
2 69970 1 9052
2 69971 1 9052
2 69972 1 9052
2 69973 1 9059
2 69974 1 9059
2 69975 1 9077
2 69976 1 9077
2 69977 1 9077
2 69978 1 9077
2 69979 1 9077
2 69980 1 9077
2 69981 1 9078
2 69982 1 9078
2 69983 1 9078
2 69984 1 9078
2 69985 1 9080
2 69986 1 9080
2 69987 1 9080
2 69988 1 9080
2 69989 1 9080
2 69990 1 9080
2 69991 1 9080
2 69992 1 9080
2 69993 1 9081
2 69994 1 9081
2 69995 1 9081
2 69996 1 9081
2 69997 1 9081
2 69998 1 9099
2 69999 1 9099
2 70000 1 9099
2 70001 1 9107
2 70002 1 9107
2 70003 1 9107
2 70004 1 9107
2 70005 1 9108
2 70006 1 9108
2 70007 1 9109
2 70008 1 9109
2 70009 1 9109
2 70010 1 9109
2 70011 1 9109
2 70012 1 9110
2 70013 1 9110
2 70014 1 9110
2 70015 1 9110
2 70016 1 9110
2 70017 1 9110
2 70018 1 9110
2 70019 1 9110
2 70020 1 9110
2 70021 1 9110
2 70022 1 9110
2 70023 1 9110
2 70024 1 9115
2 70025 1 9115
2 70026 1 9115
2 70027 1 9115
2 70028 1 9115
2 70029 1 9115
2 70030 1 9115
2 70031 1 9115
2 70032 1 9116
2 70033 1 9116
2 70034 1 9116
2 70035 1 9116
2 70036 1 9117
2 70037 1 9117
2 70038 1 9120
2 70039 1 9120
2 70040 1 9137
2 70041 1 9137
2 70042 1 9137
2 70043 1 9138
2 70044 1 9138
2 70045 1 9138
2 70046 1 9138
2 70047 1 9139
2 70048 1 9139
2 70049 1 9139
2 70050 1 9139
2 70051 1 9139
2 70052 1 9139
2 70053 1 9140
2 70054 1 9140
2 70055 1 9151
2 70056 1 9151
2 70057 1 9151
2 70058 1 9152
2 70059 1 9152
2 70060 1 9153
2 70061 1 9153
2 70062 1 9153
2 70063 1 9153
2 70064 1 9153
2 70065 1 9153
2 70066 1 9154
2 70067 1 9154
2 70068 1 9154
2 70069 1 9154
2 70070 1 9154
2 70071 1 9154
2 70072 1 9154
2 70073 1 9154
2 70074 1 9158
2 70075 1 9158
2 70076 1 9158
2 70077 1 9159
2 70078 1 9159
2 70079 1 9159
2 70080 1 9160
2 70081 1 9160
2 70082 1 9173
2 70083 1 9173
2 70084 1 9173
2 70085 1 9173
2 70086 1 9173
2 70087 1 9173
2 70088 1 9173
2 70089 1 9173
2 70090 1 9173
2 70091 1 9173
2 70092 1 9173
2 70093 1 9173
2 70094 1 9175
2 70095 1 9175
2 70096 1 9183
2 70097 1 9183
2 70098 1 9183
2 70099 1 9184
2 70100 1 9184
2 70101 1 9201
2 70102 1 9201
2 70103 1 9201
2 70104 1 9201
2 70105 1 9201
2 70106 1 9201
2 70107 1 9201
2 70108 1 9201
2 70109 1 9202
2 70110 1 9202
2 70111 1 9202
2 70112 1 9203
2 70113 1 9203
2 70114 1 9203
2 70115 1 9204
2 70116 1 9204
2 70117 1 9205
2 70118 1 9205
2 70119 1 9205
2 70120 1 9205
2 70121 1 9205
2 70122 1 9206
2 70123 1 9206
2 70124 1 9206
2 70125 1 9206
2 70126 1 9206
2 70127 1 9206
2 70128 1 9206
2 70129 1 9206
2 70130 1 9206
2 70131 1 9206
2 70132 1 9206
2 70133 1 9206
2 70134 1 9206
2 70135 1 9206
2 70136 1 9206
2 70137 1 9206
2 70138 1 9206
2 70139 1 9206
2 70140 1 9209
2 70141 1 9209
2 70142 1 9209
2 70143 1 9209
2 70144 1 9209
2 70145 1 9209
2 70146 1 9209
2 70147 1 9209
2 70148 1 9209
2 70149 1 9209
2 70150 1 9209
2 70151 1 9209
2 70152 1 9209
2 70153 1 9209
2 70154 1 9209
2 70155 1 9209
2 70156 1 9209
2 70157 1 9210
2 70158 1 9210
2 70159 1 9210
2 70160 1 9211
2 70161 1 9211
2 70162 1 9211
2 70163 1 9211
2 70164 1 9211
2 70165 1 9211
2 70166 1 9211
2 70167 1 9211
2 70168 1 9211
2 70169 1 9211
2 70170 1 9211
2 70171 1 9211
2 70172 1 9211
2 70173 1 9211
2 70174 1 9211
2 70175 1 9211
2 70176 1 9211
2 70177 1 9211
2 70178 1 9211
2 70179 1 9212
2 70180 1 9212
2 70181 1 9212
2 70182 1 9212
2 70183 1 9212
2 70184 1 9213
2 70185 1 9213
2 70186 1 9214
2 70187 1 9214
2 70188 1 9215
2 70189 1 9215
2 70190 1 9217
2 70191 1 9217
2 70192 1 9218
2 70193 1 9218
2 70194 1 9219
2 70195 1 9219
2 70196 1 9220
2 70197 1 9220
2 70198 1 9221
2 70199 1 9221
2 70200 1 9221
2 70201 1 9222
2 70202 1 9222
2 70203 1 9222
2 70204 1 9222
2 70205 1 9222
2 70206 1 9222
2 70207 1 9222
2 70208 1 9223
2 70209 1 9223
2 70210 1 9223
2 70211 1 9223
2 70212 1 9224
2 70213 1 9224
2 70214 1 9224
2 70215 1 9224
2 70216 1 9224
2 70217 1 9224
2 70218 1 9224
2 70219 1 9224
2 70220 1 9224
2 70221 1 9224
2 70222 1 9224
2 70223 1 9225
2 70224 1 9225
2 70225 1 9228
2 70226 1 9228
2 70227 1 9237
2 70228 1 9237
2 70229 1 9237
2 70230 1 9241
2 70231 1 9241
2 70232 1 9244
2 70233 1 9244
2 70234 1 9244
2 70235 1 9244
2 70236 1 9244
2 70237 1 9244
2 70238 1 9245
2 70239 1 9245
2 70240 1 9245
2 70241 1 9245
2 70242 1 9245
2 70243 1 9245
2 70244 1 9245
2 70245 1 9245
2 70246 1 9245
2 70247 1 9245
2 70248 1 9245
2 70249 1 9245
2 70250 1 9245
2 70251 1 9245
2 70252 1 9245
2 70253 1 9245
2 70254 1 9245
2 70255 1 9245
2 70256 1 9245
2 70257 1 9245
2 70258 1 9245
2 70259 1 9245
2 70260 1 9246
2 70261 1 9246
2 70262 1 9246
2 70263 1 9247
2 70264 1 9247
2 70265 1 9248
2 70266 1 9248
2 70267 1 9249
2 70268 1 9249
2 70269 1 9252
2 70270 1 9252
2 70271 1 9257
2 70272 1 9257
2 70273 1 9258
2 70274 1 9258
2 70275 1 9259
2 70276 1 9259
2 70277 1 9263
2 70278 1 9263
2 70279 1 9263
2 70280 1 9263
2 70281 1 9264
2 70282 1 9264
2 70283 1 9264
2 70284 1 9265
2 70285 1 9265
2 70286 1 9275
2 70287 1 9275
2 70288 1 9275
2 70289 1 9281
2 70290 1 9281
2 70291 1 9281
2 70292 1 9281
2 70293 1 9281
2 70294 1 9281
2 70295 1 9281
2 70296 1 9288
2 70297 1 9288
2 70298 1 9288
2 70299 1 9288
2 70300 1 9288
2 70301 1 9289
2 70302 1 9289
2 70303 1 9291
2 70304 1 9291
2 70305 1 9294
2 70306 1 9294
2 70307 1 9294
2 70308 1 9309
2 70309 1 9309
2 70310 1 9310
2 70311 1 9310
2 70312 1 9315
2 70313 1 9315
2 70314 1 9315
2 70315 1 9320
2 70316 1 9320
2 70317 1 9320
2 70318 1 9329
2 70319 1 9329
2 70320 1 9329
2 70321 1 9334
2 70322 1 9334
2 70323 1 9335
2 70324 1 9335
2 70325 1 9335
2 70326 1 9335
2 70327 1 9335
2 70328 1 9335
2 70329 1 9335
2 70330 1 9335
2 70331 1 9335
2 70332 1 9335
2 70333 1 9336
2 70334 1 9336
2 70335 1 9336
2 70336 1 9336
2 70337 1 9336
2 70338 1 9337
2 70339 1 9337
2 70340 1 9337
2 70341 1 9338
2 70342 1 9338
2 70343 1 9346
2 70344 1 9346
2 70345 1 9349
2 70346 1 9349
2 70347 1 9349
2 70348 1 9349
2 70349 1 9357
2 70350 1 9357
2 70351 1 9377
2 70352 1 9377
2 70353 1 9378
2 70354 1 9378
2 70355 1 9378
2 70356 1 9387
2 70357 1 9387
2 70358 1 9399
2 70359 1 9399
2 70360 1 9399
2 70361 1 9399
2 70362 1 9399
2 70363 1 9399
2 70364 1 9399
2 70365 1 9400
2 70366 1 9400
2 70367 1 9400
2 70368 1 9400
2 70369 1 9400
2 70370 1 9400
2 70371 1 9400
2 70372 1 9400
2 70373 1 9400
2 70374 1 9400
2 70375 1 9400
2 70376 1 9400
2 70377 1 9400
2 70378 1 9400
2 70379 1 9400
2 70380 1 9400
2 70381 1 9400
2 70382 1 9400
2 70383 1 9400
2 70384 1 9400
2 70385 1 9401
2 70386 1 9401
2 70387 1 9401
2 70388 1 9402
2 70389 1 9402
2 70390 1 9402
2 70391 1 9402
2 70392 1 9402
2 70393 1 9402
2 70394 1 9402
2 70395 1 9402
2 70396 1 9402
2 70397 1 9402
2 70398 1 9402
2 70399 1 9402
2 70400 1 9402
2 70401 1 9402
2 70402 1 9402
2 70403 1 9402
2 70404 1 9402
2 70405 1 9402
2 70406 1 9402
2 70407 1 9404
2 70408 1 9404
2 70409 1 9405
2 70410 1 9405
2 70411 1 9405
2 70412 1 9405
2 70413 1 9405
2 70414 1 9405
2 70415 1 9405
2 70416 1 9405
2 70417 1 9405
2 70418 1 9405
2 70419 1 9405
2 70420 1 9405
2 70421 1 9405
2 70422 1 9405
2 70423 1 9406
2 70424 1 9406
2 70425 1 9406
2 70426 1 9407
2 70427 1 9407
2 70428 1 9407
2 70429 1 9419
2 70430 1 9419
2 70431 1 9422
2 70432 1 9422
2 70433 1 9422
2 70434 1 9422
2 70435 1 9422
2 70436 1 9422
2 70437 1 9422
2 70438 1 9422
2 70439 1 9422
2 70440 1 9424
2 70441 1 9424
2 70442 1 9424
2 70443 1 9424
2 70444 1 9424
2 70445 1 9424
2 70446 1 9424
2 70447 1 9424
2 70448 1 9424
2 70449 1 9424
2 70450 1 9424
2 70451 1 9424
2 70452 1 9424
2 70453 1 9424
2 70454 1 9426
2 70455 1 9426
2 70456 1 9426
2 70457 1 9428
2 70458 1 9428
2 70459 1 9428
2 70460 1 9428
2 70461 1 9429
2 70462 1 9429
2 70463 1 9429
2 70464 1 9429
2 70465 1 9429
2 70466 1 9431
2 70467 1 9431
2 70468 1 9431
2 70469 1 9431
2 70470 1 9431
2 70471 1 9431
2 70472 1 9431
2 70473 1 9432
2 70474 1 9432
2 70475 1 9436
2 70476 1 9436
2 70477 1 9436
2 70478 1 9436
2 70479 1 9436
2 70480 1 9449
2 70481 1 9449
2 70482 1 9449
2 70483 1 9449
2 70484 1 9449
2 70485 1 9449
2 70486 1 9449
2 70487 1 9449
2 70488 1 9451
2 70489 1 9451
2 70490 1 9459
2 70491 1 9459
2 70492 1 9459
2 70493 1 9460
2 70494 1 9460
2 70495 1 9460
2 70496 1 9460
2 70497 1 9460
2 70498 1 9461
2 70499 1 9461
2 70500 1 9461
2 70501 1 9461
2 70502 1 9461
2 70503 1 9462
2 70504 1 9462
2 70505 1 9462
2 70506 1 9462
2 70507 1 9463
2 70508 1 9463
2 70509 1 9463
2 70510 1 9474
2 70511 1 9474
2 70512 1 9474
2 70513 1 9474
2 70514 1 9477
2 70515 1 9477
2 70516 1 9478
2 70517 1 9478
2 70518 1 9486
2 70519 1 9486
2 70520 1 9486
2 70521 1 9490
2 70522 1 9490
2 70523 1 9490
2 70524 1 9506
2 70525 1 9506
2 70526 1 9507
2 70527 1 9507
2 70528 1 9507
2 70529 1 9509
2 70530 1 9509
2 70531 1 9520
2 70532 1 9520
2 70533 1 9520
2 70534 1 9520
2 70535 1 9520
2 70536 1 9521
2 70537 1 9521
2 70538 1 9528
2 70539 1 9528
2 70540 1 9528
2 70541 1 9528
2 70542 1 9530
2 70543 1 9530
2 70544 1 9530
2 70545 1 9531
2 70546 1 9531
2 70547 1 9538
2 70548 1 9538
2 70549 1 9541
2 70550 1 9541
2 70551 1 9548
2 70552 1 9548
2 70553 1 9548
2 70554 1 9548
2 70555 1 9556
2 70556 1 9556
2 70557 1 9556
2 70558 1 9556
2 70559 1 9556
2 70560 1 9565
2 70561 1 9565
2 70562 1 9565
2 70563 1 9565
2 70564 1 9566
2 70565 1 9566
2 70566 1 9566
2 70567 1 9566
2 70568 1 9570
2 70569 1 9570
2 70570 1 9570
2 70571 1 9570
2 70572 1 9573
2 70573 1 9573
2 70574 1 9576
2 70575 1 9576
2 70576 1 9580
2 70577 1 9580
2 70578 1 9580
2 70579 1 9580
2 70580 1 9580
2 70581 1 9583
2 70582 1 9583
2 70583 1 9585
2 70584 1 9585
2 70585 1 9585
2 70586 1 9586
2 70587 1 9586
2 70588 1 9586
2 70589 1 9586
2 70590 1 9586
2 70591 1 9586
2 70592 1 9586
2 70593 1 9586
2 70594 1 9586
2 70595 1 9586
2 70596 1 9586
2 70597 1 9586
2 70598 1 9586
2 70599 1 9588
2 70600 1 9588
2 70601 1 9588
2 70602 1 9588
2 70603 1 9588
2 70604 1 9588
2 70605 1 9588
2 70606 1 9588
2 70607 1 9588
2 70608 1 9588
2 70609 1 9588
2 70610 1 9588
2 70611 1 9588
2 70612 1 9588
2 70613 1 9588
2 70614 1 9591
2 70615 1 9591
2 70616 1 9591
2 70617 1 9591
2 70618 1 9610
2 70619 1 9610
2 70620 1 9610
2 70621 1 9610
2 70622 1 9611
2 70623 1 9611
2 70624 1 9611
2 70625 1 9613
2 70626 1 9613
2 70627 1 9613
2 70628 1 9614
2 70629 1 9614
2 70630 1 9627
2 70631 1 9627
2 70632 1 9627
2 70633 1 9627
2 70634 1 9627
2 70635 1 9630
2 70636 1 9630
2 70637 1 9630
2 70638 1 9630
2 70639 1 9630
2 70640 1 9630
2 70641 1 9630
2 70642 1 9630
2 70643 1 9630
2 70644 1 9630
2 70645 1 9630
2 70646 1 9630
2 70647 1 9630
2 70648 1 9630
2 70649 1 9630
2 70650 1 9631
2 70651 1 9631
2 70652 1 9631
2 70653 1 9631
2 70654 1 9631
2 70655 1 9632
2 70656 1 9632
2 70657 1 9632
2 70658 1 9655
2 70659 1 9655
2 70660 1 9655
2 70661 1 9655
2 70662 1 9655
2 70663 1 9655
2 70664 1 9655
2 70665 1 9656
2 70666 1 9656
2 70667 1 9656
2 70668 1 9656
2 70669 1 9656
2 70670 1 9656
2 70671 1 9656
2 70672 1 9656
2 70673 1 9656
2 70674 1 9656
2 70675 1 9657
2 70676 1 9657
2 70677 1 9657
2 70678 1 9657
2 70679 1 9657
2 70680 1 9657
2 70681 1 9657
2 70682 1 9657
2 70683 1 9657
2 70684 1 9657
2 70685 1 9657
2 70686 1 9657
2 70687 1 9657
2 70688 1 9658
2 70689 1 9658
2 70690 1 9658
2 70691 1 9659
2 70692 1 9659
2 70693 1 9659
2 70694 1 9659
2 70695 1 9659
2 70696 1 9659
2 70697 1 9660
2 70698 1 9660
2 70699 1 9661
2 70700 1 9661
2 70701 1 9661
2 70702 1 9661
2 70703 1 9667
2 70704 1 9667
2 70705 1 9667
2 70706 1 9668
2 70707 1 9668
2 70708 1 9680
2 70709 1 9680
2 70710 1 9681
2 70711 1 9681
2 70712 1 9684
2 70713 1 9684
2 70714 1 9689
2 70715 1 9689
2 70716 1 9690
2 70717 1 9690
2 70718 1 9690
2 70719 1 9690
2 70720 1 9690
2 70721 1 9690
2 70722 1 9690
2 70723 1 9690
2 70724 1 9690
2 70725 1 9690
2 70726 1 9690
2 70727 1 9690
2 70728 1 9690
2 70729 1 9690
2 70730 1 9691
2 70731 1 9691
2 70732 1 9698
2 70733 1 9698
2 70734 1 9698
2 70735 1 9698
2 70736 1 9698
2 70737 1 9698
2 70738 1 9698
2 70739 1 9698
2 70740 1 9698
2 70741 1 9698
2 70742 1 9698
2 70743 1 9698
2 70744 1 9698
2 70745 1 9699
2 70746 1 9699
2 70747 1 9700
2 70748 1 9700
2 70749 1 9700
2 70750 1 9700
2 70751 1 9700
2 70752 1 9700
2 70753 1 9701
2 70754 1 9701
2 70755 1 9701
2 70756 1 9701
2 70757 1 9705
2 70758 1 9705
2 70759 1 9705
2 70760 1 9705
2 70761 1 9706
2 70762 1 9706
2 70763 1 9724
2 70764 1 9724
2 70765 1 9725
2 70766 1 9725
2 70767 1 9725
2 70768 1 9725
2 70769 1 9725
2 70770 1 9725
2 70771 1 9727
2 70772 1 9727
2 70773 1 9727
2 70774 1 9730
2 70775 1 9730
2 70776 1 9730
2 70777 1 9730
2 70778 1 9730
2 70779 1 9730
2 70780 1 9730
2 70781 1 9730
2 70782 1 9730
2 70783 1 9731
2 70784 1 9731
2 70785 1 9731
2 70786 1 9731
2 70787 1 9731
2 70788 1 9732
2 70789 1 9732
2 70790 1 9733
2 70791 1 9733
2 70792 1 9733
2 70793 1 9733
2 70794 1 9733
2 70795 1 9734
2 70796 1 9734
2 70797 1 9740
2 70798 1 9740
2 70799 1 9740
2 70800 1 9741
2 70801 1 9741
2 70802 1 9741
2 70803 1 9741
2 70804 1 9741
2 70805 1 9741
2 70806 1 9741
2 70807 1 9744
2 70808 1 9744
2 70809 1 9744
2 70810 1 9744
2 70811 1 9744
2 70812 1 9744
2 70813 1 9744
2 70814 1 9754
2 70815 1 9754
2 70816 1 9754
2 70817 1 9754
2 70818 1 9754
2 70819 1 9754
2 70820 1 9754
2 70821 1 9756
2 70822 1 9756
2 70823 1 9756
2 70824 1 9757
2 70825 1 9757
2 70826 1 9757
2 70827 1 9757
2 70828 1 9758
2 70829 1 9758
2 70830 1 9759
2 70831 1 9759
2 70832 1 9760
2 70833 1 9760
2 70834 1 9779
2 70835 1 9779
2 70836 1 9779
2 70837 1 9779
2 70838 1 9780
2 70839 1 9780
2 70840 1 9780
2 70841 1 9780
2 70842 1 9780
2 70843 1 9782
2 70844 1 9782
2 70845 1 9786
2 70846 1 9786
2 70847 1 9787
2 70848 1 9787
2 70849 1 9787
2 70850 1 9788
2 70851 1 9788
2 70852 1 9788
2 70853 1 9788
2 70854 1 9790
2 70855 1 9790
2 70856 1 9790
2 70857 1 9805
2 70858 1 9805
2 70859 1 9805
2 70860 1 9805
2 70861 1 9805
2 70862 1 9805
2 70863 1 9805
2 70864 1 9805
2 70865 1 9805
2 70866 1 9805
2 70867 1 9826
2 70868 1 9826
2 70869 1 9826
2 70870 1 9826
2 70871 1 9827
2 70872 1 9827
2 70873 1 9827
2 70874 1 9829
2 70875 1 9829
2 70876 1 9829
2 70877 1 9829
2 70878 1 9832
2 70879 1 9832
2 70880 1 9846
2 70881 1 9846
2 70882 1 9847
2 70883 1 9847
2 70884 1 9850
2 70885 1 9850
2 70886 1 9850
2 70887 1 9850
2 70888 1 9850
2 70889 1 9850
2 70890 1 9850
2 70891 1 9850
2 70892 1 9850
2 70893 1 9850
2 70894 1 9851
2 70895 1 9851
2 70896 1 9853
2 70897 1 9853
2 70898 1 9855
2 70899 1 9855
2 70900 1 9856
2 70901 1 9856
2 70902 1 9856
2 70903 1 9856
2 70904 1 9858
2 70905 1 9858
2 70906 1 9859
2 70907 1 9859
2 70908 1 9859
2 70909 1 9859
2 70910 1 9863
2 70911 1 9863
2 70912 1 9867
2 70913 1 9867
2 70914 1 9867
2 70915 1 9868
2 70916 1 9868
2 70917 1 9870
2 70918 1 9870
2 70919 1 9870
2 70920 1 9884
2 70921 1 9884
2 70922 1 9887
2 70923 1 9887
2 70924 1 9890
2 70925 1 9890
2 70926 1 9892
2 70927 1 9892
2 70928 1 9918
2 70929 1 9918
2 70930 1 9925
2 70931 1 9925
2 70932 1 9925
2 70933 1 9926
2 70934 1 9926
2 70935 1 9926
2 70936 1 9927
2 70937 1 9927
2 70938 1 9927
2 70939 1 9927
2 70940 1 9927
2 70941 1 9927
2 70942 1 9929
2 70943 1 9929
2 70944 1 9929
2 70945 1 9929
2 70946 1 9929
2 70947 1 9929
2 70948 1 9929
2 70949 1 9930
2 70950 1 9930
2 70951 1 9930
2 70952 1 9939
2 70953 1 9939
2 70954 1 9939
2 70955 1 9939
2 70956 1 9939
2 70957 1 9939
2 70958 1 9939
2 70959 1 9945
2 70960 1 9945
2 70961 1 9946
2 70962 1 9946
2 70963 1 9953
2 70964 1 9953
2 70965 1 9954
2 70966 1 9954
2 70967 1 9959
2 70968 1 9959
2 70969 1 9961
2 70970 1 9961
2 70971 1 9966
2 70972 1 9966
2 70973 1 9968
2 70974 1 9968
2 70975 1 9969
2 70976 1 9969
2 70977 1 9971
2 70978 1 9971
2 70979 1 9973
2 70980 1 9973
2 70981 1 9974
2 70982 1 9974
2 70983 1 9974
2 70984 1 9982
2 70985 1 9982
2 70986 1 9983
2 70987 1 9983
2 70988 1 9983
2 70989 1 9983
2 70990 1 9985
2 70991 1 9985
2 70992 1 9985
2 70993 1 9985
2 70994 1 9986
2 70995 1 9986
2 70996 1 9997
2 70997 1 9997
2 70998 1 9997
2 70999 1 9997
2 71000 1 9997
2 71001 1 9997
2 71002 1 9997
2 71003 1 9998
2 71004 1 9998
2 71005 1 9998
2 71006 1 9998
2 71007 1 9998
2 71008 1 9998
2 71009 1 9998
2 71010 1 10005
2 71011 1 10005
2 71012 1 10005
2 71013 1 10005
2 71014 1 10005
2 71015 1 10005
2 71016 1 10005
2 71017 1 10005
2 71018 1 10005
2 71019 1 10005
2 71020 1 10006
2 71021 1 10006
2 71022 1 10006
2 71023 1 10007
2 71024 1 10007
2 71025 1 10008
2 71026 1 10008
2 71027 1 10020
2 71028 1 10020
2 71029 1 10020
2 71030 1 10021
2 71031 1 10021
2 71032 1 10021
2 71033 1 10021
2 71034 1 10028
2 71035 1 10028
2 71036 1 10029
2 71037 1 10029
2 71038 1 10029
2 71039 1 10031
2 71040 1 10031
2 71041 1 10039
2 71042 1 10039
2 71043 1 10040
2 71044 1 10040
2 71045 1 10040
2 71046 1 10040
2 71047 1 10040
2 71048 1 10041
2 71049 1 10041
2 71050 1 10042
2 71051 1 10042
2 71052 1 10042
2 71053 1 10069
2 71054 1 10069
2 71055 1 10069
2 71056 1 10070
2 71057 1 10070
2 71058 1 10070
2 71059 1 10070
2 71060 1 10070
2 71061 1 10073
2 71062 1 10073
2 71063 1 10073
2 71064 1 10073
2 71065 1 10073
2 71066 1 10073
2 71067 1 10073
2 71068 1 10075
2 71069 1 10075
2 71070 1 10081
2 71071 1 10081
2 71072 1 10081
2 71073 1 10089
2 71074 1 10089
2 71075 1 10089
2 71076 1 10089
2 71077 1 10089
2 71078 1 10089
2 71079 1 10089
2 71080 1 10089
2 71081 1 10089
2 71082 1 10089
2 71083 1 10089
2 71084 1 10089
2 71085 1 10090
2 71086 1 10090
2 71087 1 10091
2 71088 1 10091
2 71089 1 10091
2 71090 1 10091
2 71091 1 10091
2 71092 1 10091
2 71093 1 10091
2 71094 1 10091
2 71095 1 10091
2 71096 1 10092
2 71097 1 10092
2 71098 1 10095
2 71099 1 10095
2 71100 1 10103
2 71101 1 10103
2 71102 1 10105
2 71103 1 10105
2 71104 1 10109
2 71105 1 10109
2 71106 1 10115
2 71107 1 10115
2 71108 1 10116
2 71109 1 10116
2 71110 1 10116
2 71111 1 10116
2 71112 1 10116
2 71113 1 10116
2 71114 1 10116
2 71115 1 10116
2 71116 1 10116
2 71117 1 10117
2 71118 1 10117
2 71119 1 10117
2 71120 1 10117
2 71121 1 10118
2 71122 1 10118
2 71123 1 10118
2 71124 1 10118
2 71125 1 10119
2 71126 1 10119
2 71127 1 10120
2 71128 1 10120
2 71129 1 10144
2 71130 1 10144
2 71131 1 10144
2 71132 1 10146
2 71133 1 10146
2 71134 1 10146
2 71135 1 10146
2 71136 1 10147
2 71137 1 10147
2 71138 1 10156
2 71139 1 10156
2 71140 1 10156
2 71141 1 10156
2 71142 1 10156
2 71143 1 10158
2 71144 1 10158
2 71145 1 10158
2 71146 1 10159
2 71147 1 10159
2 71148 1 10159
2 71149 1 10159
2 71150 1 10159
2 71151 1 10159
2 71152 1 10159
2 71153 1 10159
2 71154 1 10159
2 71155 1 10159
2 71156 1 10159
2 71157 1 10159
2 71158 1 10159
2 71159 1 10159
2 71160 1 10159
2 71161 1 10159
2 71162 1 10159
2 71163 1 10159
2 71164 1 10160
2 71165 1 10160
2 71166 1 10160
2 71167 1 10160
2 71168 1 10160
2 71169 1 10161
2 71170 1 10161
2 71171 1 10161
2 71172 1 10169
2 71173 1 10169
2 71174 1 10169
2 71175 1 10169
2 71176 1 10169
2 71177 1 10169
2 71178 1 10169
2 71179 1 10174
2 71180 1 10174
2 71181 1 10174
2 71182 1 10176
2 71183 1 10176
2 71184 1 10189
2 71185 1 10189
2 71186 1 10189
2 71187 1 10189
2 71188 1 10189
2 71189 1 10189
2 71190 1 10189
2 71191 1 10189
2 71192 1 10189
2 71193 1 10189
2 71194 1 10189
2 71195 1 10191
2 71196 1 10191
2 71197 1 10191
2 71198 1 10198
2 71199 1 10198
2 71200 1 10198
2 71201 1 10198
2 71202 1 10198
2 71203 1 10198
2 71204 1 10200
2 71205 1 10200
2 71206 1 10201
2 71207 1 10201
2 71208 1 10201
2 71209 1 10201
2 71210 1 10201
2 71211 1 10202
2 71212 1 10202
2 71213 1 10214
2 71214 1 10214
2 71215 1 10214
2 71216 1 10214
2 71217 1 10215
2 71218 1 10215
2 71219 1 10222
2 71220 1 10222
2 71221 1 10222
2 71222 1 10222
2 71223 1 10222
2 71224 1 10222
2 71225 1 10222
2 71226 1 10224
2 71227 1 10224
2 71228 1 10224
2 71229 1 10224
2 71230 1 10224
2 71231 1 10225
2 71232 1 10225
2 71233 1 10232
2 71234 1 10232
2 71235 1 10232
2 71236 1 10232
2 71237 1 10232
2 71238 1 10233
2 71239 1 10233
2 71240 1 10235
2 71241 1 10235
2 71242 1 10235
2 71243 1 10235
2 71244 1 10242
2 71245 1 10242
2 71246 1 10242
2 71247 1 10242
2 71248 1 10243
2 71249 1 10243
2 71250 1 10243
2 71251 1 10244
2 71252 1 10244
2 71253 1 10245
2 71254 1 10245
2 71255 1 10245
2 71256 1 10245
2 71257 1 10245
2 71258 1 10245
2 71259 1 10245
2 71260 1 10254
2 71261 1 10254
2 71262 1 10254
2 71263 1 10255
2 71264 1 10255
2 71265 1 10255
2 71266 1 10256
2 71267 1 10256
2 71268 1 10257
2 71269 1 10257
2 71270 1 10269
2 71271 1 10269
2 71272 1 10271
2 71273 1 10271
2 71274 1 10274
2 71275 1 10274
2 71276 1 10274
2 71277 1 10274
2 71278 1 10276
2 71279 1 10276
2 71280 1 10277
2 71281 1 10277
2 71282 1 10278
2 71283 1 10278
2 71284 1 10278
2 71285 1 10278
2 71286 1 10278
2 71287 1 10280
2 71288 1 10280
2 71289 1 10280
2 71290 1 10281
2 71291 1 10281
2 71292 1 10281
2 71293 1 10281
2 71294 1 10289
2 71295 1 10289
2 71296 1 10289
2 71297 1 10303
2 71298 1 10303
2 71299 1 10316
2 71300 1 10316
2 71301 1 10316
2 71302 1 10317
2 71303 1 10317
2 71304 1 10317
2 71305 1 10318
2 71306 1 10318
2 71307 1 10318
2 71308 1 10318
2 71309 1 10318
2 71310 1 10326
2 71311 1 10326
2 71312 1 10326
2 71313 1 10326
2 71314 1 10327
2 71315 1 10327
2 71316 1 10327
2 71317 1 10329
2 71318 1 10329
2 71319 1 10329
2 71320 1 10336
2 71321 1 10336
2 71322 1 10336
2 71323 1 10336
2 71324 1 10337
2 71325 1 10337
2 71326 1 10337
2 71327 1 10337
2 71328 1 10353
2 71329 1 10353
2 71330 1 10353
2 71331 1 10353
2 71332 1 10353
2 71333 1 10353
2 71334 1 10353
2 71335 1 10353
2 71336 1 10353
2 71337 1 10353
2 71338 1 10353
2 71339 1 10353
2 71340 1 10353
2 71341 1 10353
2 71342 1 10353
2 71343 1 10353
2 71344 1 10354
2 71345 1 10354
2 71346 1 10355
2 71347 1 10355
2 71348 1 10355
2 71349 1 10355
2 71350 1 10356
2 71351 1 10356
2 71352 1 10356
2 71353 1 10357
2 71354 1 10357
2 71355 1 10357
2 71356 1 10357
2 71357 1 10361
2 71358 1 10361
2 71359 1 10361
2 71360 1 10361
2 71361 1 10361
2 71362 1 10365
2 71363 1 10365
2 71364 1 10365
2 71365 1 10365
2 71366 1 10366
2 71367 1 10366
2 71368 1 10366
2 71369 1 10366
2 71370 1 10366
2 71371 1 10366
2 71372 1 10367
2 71373 1 10367
2 71374 1 10368
2 71375 1 10368
2 71376 1 10368
2 71377 1 10374
2 71378 1 10374
2 71379 1 10386
2 71380 1 10386
2 71381 1 10387
2 71382 1 10387
2 71383 1 10387
2 71384 1 10387
2 71385 1 10387
2 71386 1 10387
2 71387 1 10387
2 71388 1 10387
2 71389 1 10395
2 71390 1 10395
2 71391 1 10398
2 71392 1 10398
2 71393 1 10398
2 71394 1 10398
2 71395 1 10398
2 71396 1 10399
2 71397 1 10399
2 71398 1 10401
2 71399 1 10401
2 71400 1 10401
2 71401 1 10402
2 71402 1 10402
2 71403 1 10402
2 71404 1 10402
2 71405 1 10402
2 71406 1 10402
2 71407 1 10402
2 71408 1 10402
2 71409 1 10402
2 71410 1 10402
2 71411 1 10403
2 71412 1 10403
2 71413 1 10406
2 71414 1 10406
2 71415 1 10409
2 71416 1 10409
2 71417 1 10409
2 71418 1 10409
2 71419 1 10409
2 71420 1 10409
2 71421 1 10409
2 71422 1 10409
2 71423 1 10409
2 71424 1 10409
2 71425 1 10409
2 71426 1 10423
2 71427 1 10423
2 71428 1 10424
2 71429 1 10424
2 71430 1 10424
2 71431 1 10424
2 71432 1 10424
2 71433 1 10429
2 71434 1 10429
2 71435 1 10429
2 71436 1 10438
2 71437 1 10438
2 71438 1 10438
2 71439 1 10455
2 71440 1 10455
2 71441 1 10455
2 71442 1 10456
2 71443 1 10456
2 71444 1 10456
2 71445 1 10458
2 71446 1 10458
2 71447 1 10463
2 71448 1 10463
2 71449 1 10463
2 71450 1 10473
2 71451 1 10473
2 71452 1 10489
2 71453 1 10489
2 71454 1 10508
2 71455 1 10508
2 71456 1 10508
2 71457 1 10508
2 71458 1 10508
2 71459 1 10508
2 71460 1 10508
2 71461 1 10508
2 71462 1 10508
2 71463 1 10508
2 71464 1 10508
2 71465 1 10509
2 71466 1 10509
2 71467 1 10510
2 71468 1 10510
2 71469 1 10510
2 71470 1 10517
2 71471 1 10517
2 71472 1 10528
2 71473 1 10528
2 71474 1 10528
2 71475 1 10528
2 71476 1 10528
2 71477 1 10531
2 71478 1 10531
2 71479 1 10532
2 71480 1 10532
2 71481 1 10532
2 71482 1 10535
2 71483 1 10535
2 71484 1 10539
2 71485 1 10539
2 71486 1 10539
2 71487 1 10539
2 71488 1 10551
2 71489 1 10551
2 71490 1 10551
2 71491 1 10559
2 71492 1 10559
2 71493 1 10559
2 71494 1 10559
2 71495 1 10559
2 71496 1 10559
2 71497 1 10559
2 71498 1 10560
2 71499 1 10560
2 71500 1 10564
2 71501 1 10564
2 71502 1 10567
2 71503 1 10567
2 71504 1 10585
2 71505 1 10585
2 71506 1 10585
2 71507 1 10585
2 71508 1 10585
2 71509 1 10585
2 71510 1 10585
2 71511 1 10585
2 71512 1 10585
2 71513 1 10585
2 71514 1 10585
2 71515 1 10585
2 71516 1 10585
2 71517 1 10585
2 71518 1 10585
2 71519 1 10585
2 71520 1 10585
2 71521 1 10585
2 71522 1 10585
2 71523 1 10586
2 71524 1 10586
2 71525 1 10586
2 71526 1 10586
2 71527 1 10587
2 71528 1 10587
2 71529 1 10588
2 71530 1 10588
2 71531 1 10588
2 71532 1 10588
2 71533 1 10588
2 71534 1 10588
2 71535 1 10588
2 71536 1 10588
2 71537 1 10589
2 71538 1 10589
2 71539 1 10589
2 71540 1 10589
2 71541 1 10590
2 71542 1 10590
2 71543 1 10592
2 71544 1 10592
2 71545 1 10592
2 71546 1 10601
2 71547 1 10601
2 71548 1 10602
2 71549 1 10602
2 71550 1 10603
2 71551 1 10603
2 71552 1 10603
2 71553 1 10609
2 71554 1 10609
2 71555 1 10613
2 71556 1 10613
2 71557 1 10613
2 71558 1 10614
2 71559 1 10614
2 71560 1 10615
2 71561 1 10615
2 71562 1 10615
2 71563 1 10615
2 71564 1 10615
2 71565 1 10615
2 71566 1 10626
2 71567 1 10626
2 71568 1 10627
2 71569 1 10627
2 71570 1 10628
2 71571 1 10628
2 71572 1 10628
2 71573 1 10628
2 71574 1 10628
2 71575 1 10628
2 71576 1 10629
2 71577 1 10629
2 71578 1 10637
2 71579 1 10637
2 71580 1 10638
2 71581 1 10638
2 71582 1 10639
2 71583 1 10639
2 71584 1 10639
2 71585 1 10642
2 71586 1 10642
2 71587 1 10642
2 71588 1 10642
2 71589 1 10654
2 71590 1 10654
2 71591 1 10664
2 71592 1 10664
2 71593 1 10664
2 71594 1 10673
2 71595 1 10673
2 71596 1 10673
2 71597 1 10674
2 71598 1 10674
2 71599 1 10681
2 71600 1 10681
2 71601 1 10694
2 71602 1 10694
2 71603 1 10694
2 71604 1 10694
2 71605 1 10722
2 71606 1 10722
2 71607 1 10722
2 71608 1 10723
2 71609 1 10723
2 71610 1 10723
2 71611 1 10724
2 71612 1 10724
2 71613 1 10725
2 71614 1 10725
2 71615 1 10750
2 71616 1 10750
2 71617 1 10770
2 71618 1 10770
2 71619 1 10771
2 71620 1 10771
2 71621 1 10771
2 71622 1 10771
2 71623 1 10771
2 71624 1 10772
2 71625 1 10772
2 71626 1 10772
2 71627 1 10772
2 71628 1 10772
2 71629 1 10773
2 71630 1 10773
2 71631 1 10774
2 71632 1 10774
2 71633 1 10789
2 71634 1 10789
2 71635 1 10789
2 71636 1 10814
2 71637 1 10814
2 71638 1 10814
2 71639 1 10836
2 71640 1 10836
2 71641 1 10838
2 71642 1 10838
2 71643 1 10841
2 71644 1 10841
2 71645 1 10870
2 71646 1 10870
2 71647 1 10876
2 71648 1 10876
2 71649 1 10876
2 71650 1 10884
2 71651 1 10884
2 71652 1 10886
2 71653 1 10886
2 71654 1 10886
2 71655 1 10886
2 71656 1 10886
2 71657 1 10886
2 71658 1 10916
2 71659 1 10916
2 71660 1 10916
2 71661 1 10918
2 71662 1 10918
2 71663 1 10928
2 71664 1 10928
2 71665 1 10928
2 71666 1 10939
2 71667 1 10939
2 71668 1 10939
2 71669 1 10940
2 71670 1 10940
2 71671 1 10940
2 71672 1 10940
2 71673 1 10940
2 71674 1 10940
2 71675 1 10940
2 71676 1 10940
2 71677 1 10940
2 71678 1 10940
2 71679 1 10948
2 71680 1 10948
2 71681 1 10952
2 71682 1 10952
2 71683 1 10954
2 71684 1 10954
2 71685 1 10981
2 71686 1 10981
2 71687 1 10981
2 71688 1 10990
2 71689 1 10990
2 71690 1 11008
2 71691 1 11008
2 71692 1 11008
2 71693 1 11008
2 71694 1 11016
2 71695 1 11016
2 71696 1 11016
2 71697 1 11016
2 71698 1 11016
2 71699 1 11017
2 71700 1 11017
2 71701 1 11017
2 71702 1 11030
2 71703 1 11030
2 71704 1 11030
2 71705 1 11030
2 71706 1 11040
2 71707 1 11040
2 71708 1 11049
2 71709 1 11049
2 71710 1 11049
2 71711 1 11049
2 71712 1 11050
2 71713 1 11050
2 71714 1 11051
2 71715 1 11051
2 71716 1 11051
2 71717 1 11051
2 71718 1 11052
2 71719 1 11052
2 71720 1 11060
2 71721 1 11060
2 71722 1 11060
2 71723 1 11060
2 71724 1 11077
2 71725 1 11077
2 71726 1 11098
2 71727 1 11098
2 71728 1 11105
2 71729 1 11105
2 71730 1 11112
2 71731 1 11112
2 71732 1 11112
2 71733 1 11112
2 71734 1 11112
2 71735 1 11114
2 71736 1 11114
2 71737 1 11120
2 71738 1 11120
2 71739 1 11120
2 71740 1 11121
2 71741 1 11121
2 71742 1 11121
2 71743 1 11123
2 71744 1 11123
2 71745 1 11123
2 71746 1 11123
2 71747 1 11123
2 71748 1 11123
2 71749 1 11123
2 71750 1 11125
2 71751 1 11125
2 71752 1 11125
2 71753 1 11126
2 71754 1 11126
2 71755 1 11133
2 71756 1 11133
2 71757 1 11133
2 71758 1 11133
2 71759 1 11133
2 71760 1 11133
2 71761 1 11133
2 71762 1 11133
2 71763 1 11133
2 71764 1 11133
2 71765 1 11133
2 71766 1 11133
2 71767 1 11133
2 71768 1 11133
2 71769 1 11133
2 71770 1 11133
2 71771 1 11133
2 71772 1 11133
2 71773 1 11133
2 71774 1 11133
2 71775 1 11135
2 71776 1 11135
2 71777 1 11136
2 71778 1 11136
2 71779 1 11136
2 71780 1 11140
2 71781 1 11140
2 71782 1 11140
2 71783 1 11144
2 71784 1 11144
2 71785 1 11145
2 71786 1 11145
2 71787 1 11145
2 71788 1 11145
2 71789 1 11145
2 71790 1 11145
2 71791 1 11146
2 71792 1 11146
2 71793 1 11147
2 71794 1 11147
2 71795 1 11147
2 71796 1 11149
2 71797 1 11149
2 71798 1 11157
2 71799 1 11157
2 71800 1 11157
2 71801 1 11157
2 71802 1 11157
2 71803 1 11157
2 71804 1 11157
2 71805 1 11158
2 71806 1 11158
2 71807 1 11158
2 71808 1 11159
2 71809 1 11159
2 71810 1 11167
2 71811 1 11167
2 71812 1 11167
2 71813 1 11195
2 71814 1 11195
2 71815 1 11195
2 71816 1 11195
2 71817 1 11198
2 71818 1 11198
2 71819 1 11228
2 71820 1 11228
2 71821 1 11228
2 71822 1 11228
2 71823 1 11228
2 71824 1 11228
2 71825 1 11228
2 71826 1 11254
2 71827 1 11254
2 71828 1 11254
2 71829 1 11254
2 71830 1 11254
2 71831 1 11255
2 71832 1 11255
2 71833 1 11255
2 71834 1 11255
2 71835 1 11255
2 71836 1 11264
2 71837 1 11264
2 71838 1 11270
2 71839 1 11270
2 71840 1 11270
2 71841 1 11271
2 71842 1 11271
2 71843 1 11271
2 71844 1 11271
2 71845 1 11271
2 71846 1 11271
2 71847 1 11271
2 71848 1 11272
2 71849 1 11272
2 71850 1 11272
2 71851 1 11272
2 71852 1 11272
2 71853 1 11272
2 71854 1 11273
2 71855 1 11273
2 71856 1 11273
2 71857 1 11273
2 71858 1 11273
2 71859 1 11273
2 71860 1 11305
2 71861 1 11305
2 71862 1 11318
2 71863 1 11318
2 71864 1 11319
2 71865 1 11319
2 71866 1 11332
2 71867 1 11332
2 71868 1 11332
2 71869 1 11332
2 71870 1 11332
2 71871 1 11356
2 71872 1 11356
2 71873 1 11356
2 71874 1 11365
2 71875 1 11365
2 71876 1 11365
2 71877 1 11365
2 71878 1 11365
2 71879 1 11365
2 71880 1 11365
2 71881 1 11365
2 71882 1 11365
2 71883 1 11365
2 71884 1 11365
2 71885 1 11365
2 71886 1 11365
2 71887 1 11366
2 71888 1 11366
2 71889 1 11368
2 71890 1 11368
2 71891 1 11368
2 71892 1 11368
2 71893 1 11379
2 71894 1 11379
2 71895 1 11379
2 71896 1 11379
2 71897 1 11381
2 71898 1 11381
2 71899 1 11381
2 71900 1 11381
2 71901 1 11382
2 71902 1 11382
2 71903 1 11396
2 71904 1 11396
2 71905 1 11397
2 71906 1 11397
2 71907 1 11398
2 71908 1 11398
2 71909 1 11409
2 71910 1 11409
2 71911 1 11410
2 71912 1 11410
2 71913 1 11422
2 71914 1 11422
2 71915 1 11422
2 71916 1 11422
2 71917 1 11422
2 71918 1 11422
2 71919 1 11428
2 71920 1 11428
2 71921 1 11428
2 71922 1 11428
2 71923 1 11428
2 71924 1 11431
2 71925 1 11431
2 71926 1 11447
2 71927 1 11447
2 71928 1 11447
2 71929 1 11450
2 71930 1 11450
2 71931 1 11451
2 71932 1 11451
2 71933 1 11451
2 71934 1 11451
2 71935 1 11451
2 71936 1 11459
2 71937 1 11459
2 71938 1 11460
2 71939 1 11460
2 71940 1 11489
2 71941 1 11489
2 71942 1 11500
2 71943 1 11500
2 71944 1 11500
2 71945 1 11531
2 71946 1 11531
2 71947 1 11547
2 71948 1 11547
2 71949 1 11547
2 71950 1 11547
2 71951 1 11547
2 71952 1 11547
2 71953 1 11548
2 71954 1 11548
2 71955 1 11549
2 71956 1 11549
2 71957 1 11550
2 71958 1 11550
2 71959 1 11550
2 71960 1 11550
2 71961 1 11556
2 71962 1 11556
2 71963 1 11556
2 71964 1 11562
2 71965 1 11562
2 71966 1 11583
2 71967 1 11583
2 71968 1 11583
2 71969 1 11583
2 71970 1 11584
2 71971 1 11584
2 71972 1 11607
2 71973 1 11607
2 71974 1 11610
2 71975 1 11610
2 71976 1 11610
2 71977 1 11611
2 71978 1 11611
2 71979 1 11611
2 71980 1 11611
2 71981 1 11611
2 71982 1 11611
2 71983 1 11611
2 71984 1 11616
2 71985 1 11616
2 71986 1 11621
2 71987 1 11621
2 71988 1 11621
2 71989 1 11622
2 71990 1 11622
2 71991 1 11655
2 71992 1 11655
2 71993 1 11655
2 71994 1 11660
2 71995 1 11660
2 71996 1 11693
2 71997 1 11693
2 71998 1 11693
2 71999 1 11693
2 72000 1 11694
2 72001 1 11694
2 72002 1 11702
2 72003 1 11702
2 72004 1 11702
2 72005 1 11709
2 72006 1 11709
2 72007 1 11710
2 72008 1 11710
2 72009 1 11718
2 72010 1 11718
2 72011 1 11718
2 72012 1 11718
2 72013 1 11719
2 72014 1 11719
2 72015 1 11719
2 72016 1 11720
2 72017 1 11720
2 72018 1 11722
2 72019 1 11722
2 72020 1 11737
2 72021 1 11737
2 72022 1 11745
2 72023 1 11745
2 72024 1 11745
2 72025 1 11784
2 72026 1 11784
2 72027 1 11786
2 72028 1 11786
2 72029 1 11803
2 72030 1 11803
2 72031 1 11803
2 72032 1 11803
2 72033 1 11806
2 72034 1 11806
2 72035 1 11810
2 72036 1 11810
2 72037 1 11810
2 72038 1 11818
2 72039 1 11818
2 72040 1 11828
2 72041 1 11828
2 72042 1 11850
2 72043 1 11850
2 72044 1 11850
2 72045 1 11877
2 72046 1 11877
2 72047 1 11877
2 72048 1 11878
2 72049 1 11878
2 72050 1 11910
2 72051 1 11910
2 72052 1 11910
2 72053 1 11910
2 72054 1 11910
2 72055 1 11910
2 72056 1 11910
2 72057 1 11918
2 72058 1 11918
2 72059 1 11918
2 72060 1 11920
2 72061 1 11920
2 72062 1 11920
2 72063 1 11920
2 72064 1 11920
2 72065 1 11920
2 72066 1 11920
2 72067 1 11920
2 72068 1 11920
2 72069 1 11920
2 72070 1 11921
2 72071 1 11921
2 72072 1 11937
2 72073 1 11937
2 72074 1 11985
2 72075 1 11985
2 72076 1 11988
2 72077 1 11988
2 72078 1 11988
2 72079 1 11990
2 72080 1 11990
2 72081 1 11992
2 72082 1 11992
2 72083 1 12005
2 72084 1 12005
2 72085 1 12005
2 72086 1 12006
2 72087 1 12006
2 72088 1 12008
2 72089 1 12008
2 72090 1 12011
2 72091 1 12011
2 72092 1 12019
2 72093 1 12019
2 72094 1 12019
2 72095 1 12019
2 72096 1 12021
2 72097 1 12021
2 72098 1 12021
2 72099 1 12043
2 72100 1 12043
2 72101 1 12045
2 72102 1 12045
2 72103 1 12053
2 72104 1 12053
2 72105 1 12053
2 72106 1 12053
2 72107 1 12053
2 72108 1 12053
2 72109 1 12053
2 72110 1 12054
2 72111 1 12054
2 72112 1 12058
2 72113 1 12058
2 72114 1 12058
2 72115 1 12059
2 72116 1 12059
2 72117 1 12083
2 72118 1 12083
2 72119 1 12084
2 72120 1 12084
2 72121 1 12085
2 72122 1 12085
2 72123 1 12087
2 72124 1 12087
2 72125 1 12090
2 72126 1 12090
2 72127 1 12095
2 72128 1 12095
2 72129 1 12117
2 72130 1 12117
2 72131 1 12117
2 72132 1 12123
2 72133 1 12123
2 72134 1 12123
2 72135 1 12123
2 72136 1 12123
2 72137 1 12123
2 72138 1 12123
2 72139 1 12123
2 72140 1 12130
2 72141 1 12130
2 72142 1 12130
2 72143 1 12130
2 72144 1 12130
2 72145 1 12131
2 72146 1 12131
2 72147 1 12132
2 72148 1 12132
2 72149 1 12132
2 72150 1 12132
2 72151 1 12133
2 72152 1 12133
2 72153 1 12148
2 72154 1 12148
2 72155 1 12149
2 72156 1 12149
2 72157 1 12149
2 72158 1 12150
2 72159 1 12150
2 72160 1 12155
2 72161 1 12155
2 72162 1 12156
2 72163 1 12156
2 72164 1 12161
2 72165 1 12161
2 72166 1 12174
2 72167 1 12174
2 72168 1 12175
2 72169 1 12175
2 72170 1 12175
2 72171 1 12175
2 72172 1 12175
2 72173 1 12175
2 72174 1 12176
2 72175 1 12176
2 72176 1 12176
2 72177 1 12181
2 72178 1 12181
2 72179 1 12189
2 72180 1 12189
2 72181 1 12189
2 72182 1 12189
2 72183 1 12192
2 72184 1 12192
2 72185 1 12192
2 72186 1 12192
2 72187 1 12194
2 72188 1 12194
2 72189 1 12203
2 72190 1 12203
2 72191 1 12203
2 72192 1 12203
2 72193 1 12204
2 72194 1 12204
2 72195 1 12205
2 72196 1 12205
2 72197 1 12205
2 72198 1 12206
2 72199 1 12206
2 72200 1 12208
2 72201 1 12208
2 72202 1 12209
2 72203 1 12209
2 72204 1 12209
2 72205 1 12209
2 72206 1 12211
2 72207 1 12211
2 72208 1 12211
2 72209 1 12211
2 72210 1 12212
2 72211 1 12212
2 72212 1 12214
2 72213 1 12214
2 72214 1 12215
2 72215 1 12215
2 72216 1 12215
2 72217 1 12229
2 72218 1 12229
2 72219 1 12229
2 72220 1 12229
2 72221 1 12229
2 72222 1 12229
2 72223 1 12229
2 72224 1 12229
2 72225 1 12229
2 72226 1 12230
2 72227 1 12230
2 72228 1 12232
2 72229 1 12232
2 72230 1 12232
2 72231 1 12247
2 72232 1 12247
2 72233 1 12247
2 72234 1 12275
2 72235 1 12275
2 72236 1 12289
2 72237 1 12289
2 72238 1 12289
2 72239 1 12289
2 72240 1 12289
2 72241 1 12289
2 72242 1 12289
2 72243 1 12298
2 72244 1 12298
2 72245 1 12299
2 72246 1 12299
2 72247 1 12302
2 72248 1 12302
2 72249 1 12302
2 72250 1 12315
2 72251 1 12315
2 72252 1 12316
2 72253 1 12316
2 72254 1 12319
2 72255 1 12319
2 72256 1 12338
2 72257 1 12338
2 72258 1 12339
2 72259 1 12339
2 72260 1 12347
2 72261 1 12347
2 72262 1 12349
2 72263 1 12349
2 72264 1 12372
2 72265 1 12372
2 72266 1 12372
2 72267 1 12372
2 72268 1 12373
2 72269 1 12373
2 72270 1 12373
2 72271 1 12376
2 72272 1 12376
2 72273 1 12377
2 72274 1 12377
2 72275 1 12385
2 72276 1 12385
2 72277 1 12385
2 72278 1 12385
2 72279 1 12385
2 72280 1 12385
2 72281 1 12385
2 72282 1 12385
2 72283 1 12385
2 72284 1 12385
2 72285 1 12394
2 72286 1 12394
2 72287 1 12394
2 72288 1 12394
2 72289 1 12394
2 72290 1 12394
2 72291 1 12394
2 72292 1 12394
2 72293 1 12394
2 72294 1 12394
2 72295 1 12394
2 72296 1 12395
2 72297 1 12395
2 72298 1 12395
2 72299 1 12409
2 72300 1 12409
2 72301 1 12409
2 72302 1 12409
2 72303 1 12409
2 72304 1 12409
2 72305 1 12411
2 72306 1 12411
2 72307 1 12411
2 72308 1 12411
2 72309 1 12411
2 72310 1 12411
2 72311 1 12412
2 72312 1 12412
2 72313 1 12412
2 72314 1 12412
2 72315 1 12412
2 72316 1 12412
2 72317 1 12412
2 72318 1 12412
2 72319 1 12412
2 72320 1 12412
2 72321 1 12412
2 72322 1 12412
2 72323 1 12412
2 72324 1 12412
2 72325 1 12412
2 72326 1 12412
2 72327 1 12412
2 72328 1 12412
2 72329 1 12413
2 72330 1 12413
2 72331 1 12414
2 72332 1 12414
2 72333 1 12414
2 72334 1 12415
2 72335 1 12415
2 72336 1 12428
2 72337 1 12428
2 72338 1 12428
2 72339 1 12428
2 72340 1 12428
2 72341 1 12430
2 72342 1 12430
2 72343 1 12447
2 72344 1 12447
2 72345 1 12447
2 72346 1 12447
2 72347 1 12467
2 72348 1 12467
2 72349 1 12467
2 72350 1 12481
2 72351 1 12481
2 72352 1 12481
2 72353 1 12481
2 72354 1 12481
2 72355 1 12481
2 72356 1 12482
2 72357 1 12482
2 72358 1 12482
2 72359 1 12482
2 72360 1 12482
2 72361 1 12482
2 72362 1 12482
2 72363 1 12483
2 72364 1 12483
2 72365 1 12483
2 72366 1 12502
2 72367 1 12502
2 72368 1 12503
2 72369 1 12503
2 72370 1 12503
2 72371 1 12503
2 72372 1 12504
2 72373 1 12504
2 72374 1 12513
2 72375 1 12513
2 72376 1 12513
2 72377 1 12526
2 72378 1 12526
2 72379 1 12526
2 72380 1 12526
2 72381 1 12532
2 72382 1 12532
2 72383 1 12540
2 72384 1 12540
2 72385 1 12540
2 72386 1 12541
2 72387 1 12541
2 72388 1 12541
2 72389 1 12541
2 72390 1 12541
2 72391 1 12544
2 72392 1 12544
2 72393 1 12563
2 72394 1 12563
2 72395 1 12563
2 72396 1 12564
2 72397 1 12564
2 72398 1 12568
2 72399 1 12568
2 72400 1 12569
2 72401 1 12569
2 72402 1 12577
2 72403 1 12577
2 72404 1 12587
2 72405 1 12587
2 72406 1 12587
2 72407 1 12587
2 72408 1 12587
2 72409 1 12587
2 72410 1 12587
2 72411 1 12587
2 72412 1 12587
2 72413 1 12587
2 72414 1 12597
2 72415 1 12597
2 72416 1 12597
2 72417 1 12598
2 72418 1 12598
2 72419 1 12605
2 72420 1 12605
2 72421 1 12605
2 72422 1 12605
2 72423 1 12645
2 72424 1 12645
2 72425 1 12645
2 72426 1 12646
2 72427 1 12646
2 72428 1 12658
2 72429 1 12658
2 72430 1 12658
2 72431 1 12665
2 72432 1 12665
2 72433 1 12716
2 72434 1 12716
2 72435 1 12717
2 72436 1 12717
2 72437 1 12717
2 72438 1 12754
2 72439 1 12754
2 72440 1 12754
2 72441 1 12754
2 72442 1 12754
2 72443 1 12754
2 72444 1 12754
2 72445 1 12754
2 72446 1 12755
2 72447 1 12755
2 72448 1 12755
2 72449 1 12755
2 72450 1 12756
2 72451 1 12756
2 72452 1 12758
2 72453 1 12758
2 72454 1 12759
2 72455 1 12759
2 72456 1 12760
2 72457 1 12760
2 72458 1 12760
2 72459 1 12783
2 72460 1 12783
2 72461 1 12784
2 72462 1 12784
2 72463 1 12807
2 72464 1 12807
2 72465 1 12814
2 72466 1 12814
2 72467 1 12814
2 72468 1 12827
2 72469 1 12827
2 72470 1 12829
2 72471 1 12829
2 72472 1 12829
2 72473 1 12829
2 72474 1 12833
2 72475 1 12833
2 72476 1 12838
2 72477 1 12838
2 72478 1 12838
2 72479 1 12846
2 72480 1 12846
2 72481 1 12846
2 72482 1 12846
2 72483 1 12846
2 72484 1 12880
2 72485 1 12880
2 72486 1 12880
2 72487 1 12880
2 72488 1 12880
2 72489 1 12880
2 72490 1 12884
2 72491 1 12884
2 72492 1 12894
2 72493 1 12894
2 72494 1 12904
2 72495 1 12904
2 72496 1 12904
2 72497 1 12905
2 72498 1 12905
2 72499 1 12923
2 72500 1 12923
2 72501 1 12936
2 72502 1 12936
2 72503 1 12937
2 72504 1 12937
2 72505 1 12946
2 72506 1 12946
2 72507 1 12957
2 72508 1 12957
2 72509 1 12957
2 72510 1 12959
2 72511 1 12959
2 72512 1 12959
2 72513 1 12970
2 72514 1 12970
2 72515 1 12972
2 72516 1 12972
2 72517 1 12973
2 72518 1 12973
2 72519 1 12984
2 72520 1 12984
2 72521 1 13015
2 72522 1 13015
2 72523 1 13015
2 72524 1 13027
2 72525 1 13027
2 72526 1 13028
2 72527 1 13028
2 72528 1 13028
2 72529 1 13028
2 72530 1 13028
2 72531 1 13028
2 72532 1 13029
2 72533 1 13029
2 72534 1 13049
2 72535 1 13049
2 72536 1 13049
2 72537 1 13049
2 72538 1 13049
2 72539 1 13049
2 72540 1 13070
2 72541 1 13070
2 72542 1 13073
2 72543 1 13073
2 72544 1 13073
2 72545 1 13081
2 72546 1 13081
2 72547 1 13081
2 72548 1 13100
2 72549 1 13100
2 72550 1 13108
2 72551 1 13108
2 72552 1 13109
2 72553 1 13109
2 72554 1 13109
2 72555 1 13118
2 72556 1 13118
2 72557 1 13139
2 72558 1 13139
2 72559 1 13149
2 72560 1 13149
2 72561 1 13153
2 72562 1 13153
2 72563 1 13153
2 72564 1 13153
2 72565 1 13154
2 72566 1 13154
2 72567 1 13154
2 72568 1 13156
2 72569 1 13156
2 72570 1 13178
2 72571 1 13178
2 72572 1 13178
2 72573 1 13178
2 72574 1 13178
2 72575 1 13178
2 72576 1 13178
2 72577 1 13179
2 72578 1 13179
2 72579 1 13179
2 72580 1 13179
2 72581 1 13199
2 72582 1 13199
2 72583 1 13200
2 72584 1 13200
2 72585 1 13232
2 72586 1 13232
2 72587 1 13232
2 72588 1 13248
2 72589 1 13248
2 72590 1 13248
2 72591 1 13255
2 72592 1 13255
2 72593 1 13255
2 72594 1 13255
2 72595 1 13255
2 72596 1 13255
2 72597 1 13255
2 72598 1 13255
2 72599 1 13255
2 72600 1 13255
2 72601 1 13255
2 72602 1 13255
2 72603 1 13255
2 72604 1 13270
2 72605 1 13270
2 72606 1 13279
2 72607 1 13279
2 72608 1 13279
2 72609 1 13280
2 72610 1 13280
2 72611 1 13303
2 72612 1 13303
2 72613 1 13308
2 72614 1 13308
2 72615 1 13309
2 72616 1 13309
2 72617 1 13309
2 72618 1 13309
2 72619 1 13310
2 72620 1 13310
2 72621 1 13322
2 72622 1 13322
2 72623 1 13322
2 72624 1 13337
2 72625 1 13337
2 72626 1 13342
2 72627 1 13342
2 72628 1 13343
2 72629 1 13343
2 72630 1 13344
2 72631 1 13344
2 72632 1 13344
2 72633 1 13344
2 72634 1 13345
2 72635 1 13345
2 72636 1 13355
2 72637 1 13355
2 72638 1 13355
2 72639 1 13366
2 72640 1 13366
2 72641 1 13369
2 72642 1 13369
2 72643 1 13389
2 72644 1 13389
2 72645 1 13389
2 72646 1 13394
2 72647 1 13394
2 72648 1 13394
2 72649 1 13394
2 72650 1 13394
2 72651 1 13394
2 72652 1 13394
2 72653 1 13395
2 72654 1 13395
2 72655 1 13396
2 72656 1 13396
2 72657 1 13397
2 72658 1 13397
2 72659 1 13401
2 72660 1 13401
2 72661 1 13409
2 72662 1 13409
2 72663 1 13410
2 72664 1 13410
2 72665 1 13411
2 72666 1 13411
2 72667 1 13412
2 72668 1 13412
2 72669 1 13418
2 72670 1 13418
2 72671 1 13422
2 72672 1 13422
2 72673 1 13428
2 72674 1 13428
2 72675 1 13431
2 72676 1 13431
2 72677 1 13431
2 72678 1 13432
2 72679 1 13432
2 72680 1 13432
2 72681 1 13432
2 72682 1 13432
2 72683 1 13435
2 72684 1 13435
2 72685 1 13435
2 72686 1 13435
2 72687 1 13436
2 72688 1 13436
2 72689 1 13460
2 72690 1 13460
2 72691 1 13460
2 72692 1 13460
2 72693 1 13460
2 72694 1 13461
2 72695 1 13461
2 72696 1 13462
2 72697 1 13462
2 72698 1 13462
2 72699 1 13469
2 72700 1 13469
2 72701 1 13470
2 72702 1 13470
2 72703 1 13470
2 72704 1 13471
2 72705 1 13471
2 72706 1 13471
2 72707 1 13471
2 72708 1 13471
2 72709 1 13471
2 72710 1 13471
2 72711 1 13471
2 72712 1 13471
2 72713 1 13471
2 72714 1 13471
2 72715 1 13471
2 72716 1 13471
2 72717 1 13471
2 72718 1 13471
2 72719 1 13471
2 72720 1 13471
2 72721 1 13471
2 72722 1 13471
2 72723 1 13472
2 72724 1 13472
2 72725 1 13472
2 72726 1 13473
2 72727 1 13473
2 72728 1 13473
2 72729 1 13486
2 72730 1 13486
2 72731 1 13486
2 72732 1 13486
2 72733 1 13488
2 72734 1 13488
2 72735 1 13490
2 72736 1 13490
2 72737 1 13491
2 72738 1 13491
2 72739 1 13491
2 72740 1 13493
2 72741 1 13493
2 72742 1 13505
2 72743 1 13505
2 72744 1 13532
2 72745 1 13532
2 72746 1 13536
2 72747 1 13536
2 72748 1 13543
2 72749 1 13543
2 72750 1 13569
2 72751 1 13569
2 72752 1 13570
2 72753 1 13570
2 72754 1 13570
2 72755 1 13570
2 72756 1 13572
2 72757 1 13572
2 72758 1 13572
2 72759 1 13572
2 72760 1 13572
2 72761 1 13577
2 72762 1 13577
2 72763 1 13590
2 72764 1 13590
2 72765 1 13590
2 72766 1 13590
2 72767 1 13590
2 72768 1 13590
2 72769 1 13592
2 72770 1 13592
2 72771 1 13594
2 72772 1 13594
2 72773 1 13597
2 72774 1 13597
2 72775 1 13611
2 72776 1 13611
2 72777 1 13644
2 72778 1 13644
2 72779 1 13645
2 72780 1 13645
2 72781 1 13645
2 72782 1 13645
2 72783 1 13645
2 72784 1 13645
2 72785 1 13646
2 72786 1 13646
2 72787 1 13647
2 72788 1 13647
2 72789 1 13650
2 72790 1 13650
2 72791 1 13650
2 72792 1 13650
2 72793 1 13650
2 72794 1 13650
2 72795 1 13650
2 72796 1 13651
2 72797 1 13651
2 72798 1 13651
2 72799 1 13654
2 72800 1 13654
2 72801 1 13654
2 72802 1 13658
2 72803 1 13658
2 72804 1 13700
2 72805 1 13700
2 72806 1 13725
2 72807 1 13725
2 72808 1 13726
2 72809 1 13726
2 72810 1 13726
2 72811 1 13726
2 72812 1 13726
2 72813 1 13726
2 72814 1 13726
2 72815 1 13738
2 72816 1 13738
2 72817 1 13741
2 72818 1 13741
2 72819 1 13762
2 72820 1 13762
2 72821 1 13762
2 72822 1 13762
2 72823 1 13762
2 72824 1 13762
2 72825 1 13788
2 72826 1 13788
2 72827 1 13789
2 72828 1 13789
2 72829 1 13798
2 72830 1 13798
2 72831 1 13820
2 72832 1 13820
2 72833 1 13834
2 72834 1 13834
2 72835 1 13835
2 72836 1 13835
2 72837 1 13836
2 72838 1 13836
2 72839 1 13864
2 72840 1 13864
2 72841 1 13864
2 72842 1 13864
2 72843 1 13864
2 72844 1 13869
2 72845 1 13869
2 72846 1 13898
2 72847 1 13898
2 72848 1 13898
2 72849 1 13905
2 72850 1 13905
2 72851 1 13922
2 72852 1 13922
2 72853 1 13922
2 72854 1 13922
2 72855 1 13922
2 72856 1 13923
2 72857 1 13923
2 72858 1 13923
2 72859 1 13924
2 72860 1 13924
2 72861 1 13939
2 72862 1 13939
2 72863 1 13960
2 72864 1 13960
2 72865 1 13974
2 72866 1 13974
2 72867 1 13975
2 72868 1 13975
2 72869 1 13986
2 72870 1 13986
2 72871 1 13986
2 72872 1 13986
2 72873 1 14007
2 72874 1 14007
2 72875 1 14007
2 72876 1 14007
2 72877 1 14009
2 72878 1 14009
2 72879 1 14023
2 72880 1 14023
2 72881 1 14041
2 72882 1 14041
2 72883 1 14041
2 72884 1 14041
2 72885 1 14041
2 72886 1 14049
2 72887 1 14049
2 72888 1 14049
2 72889 1 14049
2 72890 1 14049
2 72891 1 14057
2 72892 1 14057
2 72893 1 14057
2 72894 1 14057
2 72895 1 14057
2 72896 1 14058
2 72897 1 14058
2 72898 1 14078
2 72899 1 14078
2 72900 1 14109
2 72901 1 14109
2 72902 1 14109
2 72903 1 14109
2 72904 1 14109
2 72905 1 14109
2 72906 1 14110
2 72907 1 14110
2 72908 1 14111
2 72909 1 14111
2 72910 1 14115
2 72911 1 14115
2 72912 1 14115
2 72913 1 14125
2 72914 1 14125
2 72915 1 14154
2 72916 1 14154
2 72917 1 14160
2 72918 1 14160
2 72919 1 14168
2 72920 1 14168
2 72921 1 14172
2 72922 1 14172
2 72923 1 14172
2 72924 1 14174
2 72925 1 14174
2 72926 1 14177
2 72927 1 14177
2 72928 1 14177
2 72929 1 14177
2 72930 1 14177
2 72931 1 14177
2 72932 1 14177
2 72933 1 14177
2 72934 1 14178
2 72935 1 14178
2 72936 1 14194
2 72937 1 14194
2 72938 1 14200
2 72939 1 14200
2 72940 1 14200
2 72941 1 14200
2 72942 1 14201
2 72943 1 14201
2 72944 1 14201
2 72945 1 14201
2 72946 1 14202
2 72947 1 14202
2 72948 1 14202
2 72949 1 14220
2 72950 1 14220
2 72951 1 14221
2 72952 1 14221
2 72953 1 14228
2 72954 1 14228
2 72955 1 14232
2 72956 1 14232
2 72957 1 14232
2 72958 1 14240
2 72959 1 14240
2 72960 1 14240
2 72961 1 14240
2 72962 1 14241
2 72963 1 14241
2 72964 1 14244
2 72965 1 14244
2 72966 1 14244
2 72967 1 14244
2 72968 1 14244
2 72969 1 14245
2 72970 1 14245
2 72971 1 14247
2 72972 1 14247
2 72973 1 14266
2 72974 1 14266
2 72975 1 14266
2 72976 1 14266
2 72977 1 14266
2 72978 1 14266
2 72979 1 14267
2 72980 1 14267
2 72981 1 14268
2 72982 1 14268
2 72983 1 14268
2 72984 1 14279
2 72985 1 14279
2 72986 1 14279
2 72987 1 14279
2 72988 1 14279
2 72989 1 14279
2 72990 1 14279
2 72991 1 14281
2 72992 1 14281
2 72993 1 14281
2 72994 1 14294
2 72995 1 14294
2 72996 1 14294
2 72997 1 14294
2 72998 1 14294
2 72999 1 14294
2 73000 1 14294
2 73001 1 14294
2 73002 1 14294
2 73003 1 14294
2 73004 1 14294
2 73005 1 14296
2 73006 1 14296
2 73007 1 14298
2 73008 1 14298
2 73009 1 14299
2 73010 1 14299
2 73011 1 14303
2 73012 1 14303
2 73013 1 14304
2 73014 1 14304
2 73015 1 14329
2 73016 1 14329
2 73017 1 14329
2 73018 1 14329
2 73019 1 14329
2 73020 1 14329
2 73021 1 14329
2 73022 1 14329
2 73023 1 14329
2 73024 1 14329
2 73025 1 14330
2 73026 1 14330
2 73027 1 14331
2 73028 1 14331
2 73029 1 14337
2 73030 1 14337
2 73031 1 14338
2 73032 1 14338
2 73033 1 14338
2 73034 1 14345
2 73035 1 14345
2 73036 1 14345
2 73037 1 14345
2 73038 1 14345
2 73039 1 14345
2 73040 1 14345
2 73041 1 14345
2 73042 1 14345
2 73043 1 14345
2 73044 1 14345
2 73045 1 14345
2 73046 1 14345
2 73047 1 14350
2 73048 1 14350
2 73049 1 14368
2 73050 1 14368
2 73051 1 14377
2 73052 1 14377
2 73053 1 14377
2 73054 1 14377
2 73055 1 14378
2 73056 1 14378
2 73057 1 14378
2 73058 1 14379
2 73059 1 14379
2 73060 1 14379
2 73061 1 14386
2 73062 1 14386
2 73063 1 14386
2 73064 1 14398
2 73065 1 14398
2 73066 1 14398
2 73067 1 14398
2 73068 1 14398
2 73069 1 14399
2 73070 1 14399
2 73071 1 14401
2 73072 1 14401
2 73073 1 14402
2 73074 1 14402
2 73075 1 14404
2 73076 1 14404
2 73077 1 14404
2 73078 1 14404
2 73079 1 14404
2 73080 1 14404
2 73081 1 14404
2 73082 1 14404
2 73083 1 14404
2 73084 1 14405
2 73085 1 14405
2 73086 1 14407
2 73087 1 14407
2 73088 1 14415
2 73089 1 14415
2 73090 1 14415
2 73091 1 14415
2 73092 1 14415
2 73093 1 14415
2 73094 1 14417
2 73095 1 14417
2 73096 1 14418
2 73097 1 14418
2 73098 1 14418
2 73099 1 14418
2 73100 1 14420
2 73101 1 14420
2 73102 1 14421
2 73103 1 14421
2 73104 1 14423
2 73105 1 14423
2 73106 1 14434
2 73107 1 14434
2 73108 1 14448
2 73109 1 14448
2 73110 1 14448
2 73111 1 14448
2 73112 1 14448
2 73113 1 14448
2 73114 1 14450
2 73115 1 14450
2 73116 1 14451
2 73117 1 14451
2 73118 1 14457
2 73119 1 14457
2 73120 1 14457
2 73121 1 14457
2 73122 1 14457
2 73123 1 14457
2 73124 1 14458
2 73125 1 14458
2 73126 1 14467
2 73127 1 14467
2 73128 1 14467
2 73129 1 14467
2 73130 1 14467
2 73131 1 14468
2 73132 1 14468
2 73133 1 14475
2 73134 1 14475
2 73135 1 14475
2 73136 1 14475
2 73137 1 14476
2 73138 1 14476
2 73139 1 14476
2 73140 1 14481
2 73141 1 14481
2 73142 1 14491
2 73143 1 14491
2 73144 1 14515
2 73145 1 14515
2 73146 1 14516
2 73147 1 14516
2 73148 1 14518
2 73149 1 14518
2 73150 1 14519
2 73151 1 14519
2 73152 1 14529
2 73153 1 14529
2 73154 1 14529
2 73155 1 14529
2 73156 1 14529
2 73157 1 14529
2 73158 1 14533
2 73159 1 14533
2 73160 1 14533
2 73161 1 14533
2 73162 1 14533
2 73163 1 14533
2 73164 1 14540
2 73165 1 14540
2 73166 1 14540
2 73167 1 14541
2 73168 1 14541
2 73169 1 14548
2 73170 1 14548
2 73171 1 14566
2 73172 1 14566
2 73173 1 14566
2 73174 1 14566
2 73175 1 14566
2 73176 1 14578
2 73177 1 14578
2 73178 1 14584
2 73179 1 14584
2 73180 1 14585
2 73181 1 14585
2 73182 1 14585
2 73183 1 14586
2 73184 1 14586
2 73185 1 14592
2 73186 1 14592
2 73187 1 14593
2 73188 1 14593
2 73189 1 14593
2 73190 1 14611
2 73191 1 14611
2 73192 1 14611
2 73193 1 14613
2 73194 1 14613
2 73195 1 14614
2 73196 1 14614
2 73197 1 14617
2 73198 1 14617
2 73199 1 14617
2 73200 1 14617
2 73201 1 14617
2 73202 1 14617
2 73203 1 14617
2 73204 1 14617
2 73205 1 14617
2 73206 1 14617
2 73207 1 14617
2 73208 1 14618
2 73209 1 14618
2 73210 1 14626
2 73211 1 14626
2 73212 1 14626
2 73213 1 14628
2 73214 1 14628
2 73215 1 14628
2 73216 1 14630
2 73217 1 14630
2 73218 1 14630
2 73219 1 14631
2 73220 1 14631
2 73221 1 14646
2 73222 1 14646
2 73223 1 14646
2 73224 1 14646
2 73225 1 14646
2 73226 1 14646
2 73227 1 14647
2 73228 1 14647
2 73229 1 14652
2 73230 1 14652
2 73231 1 14652
2 73232 1 14652
2 73233 1 14663
2 73234 1 14663
2 73235 1 14663
2 73236 1 14663
2 73237 1 14684
2 73238 1 14684
2 73239 1 14688
2 73240 1 14688
2 73241 1 14697
2 73242 1 14697
2 73243 1 14707
2 73244 1 14707
2 73245 1 14709
2 73246 1 14709
2 73247 1 14709
2 73248 1 14709
2 73249 1 14709
2 73250 1 14709
2 73251 1 14709
2 73252 1 14709
2 73253 1 14709
2 73254 1 14709
2 73255 1 14709
2 73256 1 14709
2 73257 1 14709
2 73258 1 14711
2 73259 1 14711
2 73260 1 14711
2 73261 1 14728
2 73262 1 14728
2 73263 1 14737
2 73264 1 14737
2 73265 1 14737
2 73266 1 14737
2 73267 1 14737
2 73268 1 14737
2 73269 1 14745
2 73270 1 14745
2 73271 1 14745
2 73272 1 14746
2 73273 1 14746
2 73274 1 14746
2 73275 1 14746
2 73276 1 14746
2 73277 1 14749
2 73278 1 14749
2 73279 1 14771
2 73280 1 14771
2 73281 1 14771
2 73282 1 14774
2 73283 1 14774
2 73284 1 14774
2 73285 1 14790
2 73286 1 14790
2 73287 1 14804
2 73288 1 14804
2 73289 1 14804
2 73290 1 14804
2 73291 1 14804
2 73292 1 14804
2 73293 1 14805
2 73294 1 14805
2 73295 1 14805
2 73296 1 14808
2 73297 1 14808
2 73298 1 14808
2 73299 1 14809
2 73300 1 14809
2 73301 1 14823
2 73302 1 14823
2 73303 1 14823
2 73304 1 14823
2 73305 1 14823
2 73306 1 14823
2 73307 1 14823
2 73308 1 14823
2 73309 1 14824
2 73310 1 14824
2 73311 1 14824
2 73312 1 14825
2 73313 1 14825
2 73314 1 14825
2 73315 1 14825
2 73316 1 14834
2 73317 1 14834
2 73318 1 14834
2 73319 1 14834
2 73320 1 14834
2 73321 1 14834
2 73322 1 14834
2 73323 1 14834
2 73324 1 14834
2 73325 1 14835
2 73326 1 14835
2 73327 1 14835
2 73328 1 14839
2 73329 1 14839
2 73330 1 14841
2 73331 1 14841
2 73332 1 14842
2 73333 1 14842
2 73334 1 14861
2 73335 1 14861
2 73336 1 14871
2 73337 1 14871
2 73338 1 14871
2 73339 1 14871
2 73340 1 14872
2 73341 1 14872
2 73342 1 14872
2 73343 1 14872
2 73344 1 14874
2 73345 1 14874
2 73346 1 14874
2 73347 1 14874
2 73348 1 14877
2 73349 1 14877
2 73350 1 14884
2 73351 1 14884
2 73352 1 14884
2 73353 1 14891
2 73354 1 14891
2 73355 1 14891
2 73356 1 14891
2 73357 1 14891
2 73358 1 14893
2 73359 1 14893
2 73360 1 14893
2 73361 1 14893
2 73362 1 14893
2 73363 1 14893
2 73364 1 14893
2 73365 1 14894
2 73366 1 14894
2 73367 1 14905
2 73368 1 14905
2 73369 1 14905
2 73370 1 14905
2 73371 1 14905
2 73372 1 14905
2 73373 1 14905
2 73374 1 14905
2 73375 1 14905
2 73376 1 14905
2 73377 1 14908
2 73378 1 14908
2 73379 1 14918
2 73380 1 14918
2 73381 1 14918
2 73382 1 14918
2 73383 1 14918
2 73384 1 14918
2 73385 1 14918
2 73386 1 14918
2 73387 1 14918
2 73388 1 14919
2 73389 1 14919
2 73390 1 14920
2 73391 1 14920
2 73392 1 14920
2 73393 1 14920
2 73394 1 14931
2 73395 1 14931
2 73396 1 14931
2 73397 1 14934
2 73398 1 14934
2 73399 1 14943
2 73400 1 14943
2 73401 1 14943
2 73402 1 14951
2 73403 1 14951
2 73404 1 14951
2 73405 1 14951
2 73406 1 14951
2 73407 1 14952
2 73408 1 14952
2 73409 1 14977
2 73410 1 14977
2 73411 1 14977
2 73412 1 14977
2 73413 1 14977
2 73414 1 14977
2 73415 1 14977
2 73416 1 14979
2 73417 1 14979
2 73418 1 14979
2 73419 1 14980
2 73420 1 14980
2 73421 1 14997
2 73422 1 14997
2 73423 1 14998
2 73424 1 14998
2 73425 1 14998
2 73426 1 14998
2 73427 1 14998
2 73428 1 14998
2 73429 1 14998
2 73430 1 14998
2 73431 1 14998
2 73432 1 14998
2 73433 1 14999
2 73434 1 14999
2 73435 1 14999
2 73436 1 15011
2 73437 1 15011
2 73438 1 15011
2 73439 1 15011
2 73440 1 15011
2 73441 1 15011
2 73442 1 15011
2 73443 1 15011
2 73444 1 15011
2 73445 1 15011
2 73446 1 15012
2 73447 1 15012
2 73448 1 15018
2 73449 1 15018
2 73450 1 15020
2 73451 1 15020
2 73452 1 15020
2 73453 1 15033
2 73454 1 15033
2 73455 1 15033
2 73456 1 15047
2 73457 1 15047
2 73458 1 15048
2 73459 1 15048
2 73460 1 15048
2 73461 1 15070
2 73462 1 15070
2 73463 1 15070
2 73464 1 15074
2 73465 1 15074
2 73466 1 15074
2 73467 1 15075
2 73468 1 15075
2 73469 1 15075
2 73470 1 15083
2 73471 1 15083
2 73472 1 15083
2 73473 1 15089
2 73474 1 15089
2 73475 1 15099
2 73476 1 15099
2 73477 1 15099
2 73478 1 15099
2 73479 1 15100
2 73480 1 15100
2 73481 1 15100
2 73482 1 15100
2 73483 1 15100
2 73484 1 15100
2 73485 1 15101
2 73486 1 15101
2 73487 1 15103
2 73488 1 15103
2 73489 1 15103
2 73490 1 15106
2 73491 1 15106
2 73492 1 15106
2 73493 1 15106
2 73494 1 15106
2 73495 1 15106
2 73496 1 15107
2 73497 1 15107
2 73498 1 15109
2 73499 1 15109
2 73500 1 15109
2 73501 1 15110
2 73502 1 15110
2 73503 1 15110
2 73504 1 15122
2 73505 1 15122
2 73506 1 15122
2 73507 1 15135
2 73508 1 15135
2 73509 1 15146
2 73510 1 15146
2 73511 1 15147
2 73512 1 15147
2 73513 1 15156
2 73514 1 15156
2 73515 1 15156
2 73516 1 15156
2 73517 1 15156
2 73518 1 15156
2 73519 1 15157
2 73520 1 15157
2 73521 1 15157
2 73522 1 15157
2 73523 1 15157
2 73524 1 15157
2 73525 1 15157
2 73526 1 15157
2 73527 1 15157
2 73528 1 15157
2 73529 1 15157
2 73530 1 15157
2 73531 1 15157
2 73532 1 15157
2 73533 1 15157
2 73534 1 15157
2 73535 1 15158
2 73536 1 15158
2 73537 1 15170
2 73538 1 15170
2 73539 1 15178
2 73540 1 15178
2 73541 1 15178
2 73542 1 15178
2 73543 1 15179
2 73544 1 15179
2 73545 1 15179
2 73546 1 15187
2 73547 1 15187
2 73548 1 15187
2 73549 1 15187
2 73550 1 15198
2 73551 1 15198
2 73552 1 15198
2 73553 1 15198
2 73554 1 15198
2 73555 1 15198
2 73556 1 15200
2 73557 1 15200
2 73558 1 15202
2 73559 1 15202
2 73560 1 15207
2 73561 1 15207
2 73562 1 15207
2 73563 1 15207
2 73564 1 15207
2 73565 1 15207
2 73566 1 15207
2 73567 1 15215
2 73568 1 15215
2 73569 1 15215
2 73570 1 15215
2 73571 1 15215
2 73572 1 15215
2 73573 1 15215
2 73574 1 15215
2 73575 1 15215
2 73576 1 15215
2 73577 1 15217
2 73578 1 15217
2 73579 1 15231
2 73580 1 15231
2 73581 1 15233
2 73582 1 15233
2 73583 1 15234
2 73584 1 15234
2 73585 1 15235
2 73586 1 15235
2 73587 1 15244
2 73588 1 15244
2 73589 1 15262
2 73590 1 15262
2 73591 1 15272
2 73592 1 15272
2 73593 1 15272
2 73594 1 15272
2 73595 1 15273
2 73596 1 15273
2 73597 1 15295
2 73598 1 15295
2 73599 1 15295
2 73600 1 15309
2 73601 1 15309
2 73602 1 15309
2 73603 1 15309
2 73604 1 15310
2 73605 1 15310
2 73606 1 15311
2 73607 1 15311
2 73608 1 15311
2 73609 1 15318
2 73610 1 15318
2 73611 1 15318
2 73612 1 15340
2 73613 1 15340
2 73614 1 15340
2 73615 1 15340
2 73616 1 15341
2 73617 1 15341
2 73618 1 15359
2 73619 1 15359
2 73620 1 15366
2 73621 1 15366
2 73622 1 15367
2 73623 1 15367
2 73624 1 15367
2 73625 1 15375
2 73626 1 15375
2 73627 1 15376
2 73628 1 15376
2 73629 1 15377
2 73630 1 15377
2 73631 1 15383
2 73632 1 15383
2 73633 1 15383
2 73634 1 15383
2 73635 1 15383
2 73636 1 15384
2 73637 1 15384
2 73638 1 15402
2 73639 1 15402
2 73640 1 15405
2 73641 1 15405
2 73642 1 15405
2 73643 1 15405
2 73644 1 15405
2 73645 1 15405
2 73646 1 15405
2 73647 1 15412
2 73648 1 15412
2 73649 1 15412
2 73650 1 15412
2 73651 1 15412
2 73652 1 15412
2 73653 1 15412
2 73654 1 15413
2 73655 1 15413
2 73656 1 15413
2 73657 1 15413
2 73658 1 15413
2 73659 1 15413
2 73660 1 15414
2 73661 1 15414
2 73662 1 15415
2 73663 1 15415
2 73664 1 15423
2 73665 1 15423
2 73666 1 15439
2 73667 1 15439
2 73668 1 15442
2 73669 1 15442
2 73670 1 15442
2 73671 1 15455
2 73672 1 15455
2 73673 1 15457
2 73674 1 15457
2 73675 1 15457
2 73676 1 15457
2 73677 1 15457
2 73678 1 15457
2 73679 1 15457
2 73680 1 15457
2 73681 1 15458
2 73682 1 15458
2 73683 1 15465
2 73684 1 15465
2 73685 1 15474
2 73686 1 15474
2 73687 1 15475
2 73688 1 15475
2 73689 1 15485
2 73690 1 15485
2 73691 1 15508
2 73692 1 15508
2 73693 1 15508
2 73694 1 15514
2 73695 1 15514
2 73696 1 15515
2 73697 1 15515
2 73698 1 15515
2 73699 1 15515
2 73700 1 15530
2 73701 1 15530
2 73702 1 15532
2 73703 1 15532
2 73704 1 15532
2 73705 1 15532
2 73706 1 15532
2 73707 1 15532
2 73708 1 15532
2 73709 1 15532
2 73710 1 15535
2 73711 1 15535
2 73712 1 15535
2 73713 1 15535
2 73714 1 15535
2 73715 1 15535
2 73716 1 15535
2 73717 1 15535
2 73718 1 15539
2 73719 1 15539
2 73720 1 15546
2 73721 1 15546
2 73722 1 15551
2 73723 1 15551
2 73724 1 15551
2 73725 1 15551
2 73726 1 15552
2 73727 1 15552
2 73728 1 15552
2 73729 1 15552
2 73730 1 15552
2 73731 1 15552
2 73732 1 15552
2 73733 1 15573
2 73734 1 15573
2 73735 1 15575
2 73736 1 15575
2 73737 1 15575
2 73738 1 15575
2 73739 1 15575
2 73740 1 15575
2 73741 1 15576
2 73742 1 15576
2 73743 1 15576
2 73744 1 15576
2 73745 1 15577
2 73746 1 15577
2 73747 1 15577
2 73748 1 15577
2 73749 1 15577
2 73750 1 15577
2 73751 1 15578
2 73752 1 15578
2 73753 1 15581
2 73754 1 15581
2 73755 1 15582
2 73756 1 15582
2 73757 1 15582
2 73758 1 15582
2 73759 1 15585
2 73760 1 15585
2 73761 1 15596
2 73762 1 15596
2 73763 1 15596
2 73764 1 15596
2 73765 1 15597
2 73766 1 15597
2 73767 1 15608
2 73768 1 15608
2 73769 1 15608
2 73770 1 15608
2 73771 1 15608
2 73772 1 15608
2 73773 1 15608
2 73774 1 15609
2 73775 1 15609
2 73776 1 15613
2 73777 1 15613
2 73778 1 15613
2 73779 1 15619
2 73780 1 15619
2 73781 1 15619
2 73782 1 15619
2 73783 1 15620
2 73784 1 15620
2 73785 1 15645
2 73786 1 15645
2 73787 1 15655
2 73788 1 15655
2 73789 1 15657
2 73790 1 15657
2 73791 1 15658
2 73792 1 15658
2 73793 1 15658
2 73794 1 15661
2 73795 1 15661
2 73796 1 15661
2 73797 1 15668
2 73798 1 15668
2 73799 1 15668
2 73800 1 15668
2 73801 1 15682
2 73802 1 15682
2 73803 1 15682
2 73804 1 15682
2 73805 1 15683
2 73806 1 15683
2 73807 1 15684
2 73808 1 15684
2 73809 1 15692
2 73810 1 15692
2 73811 1 15692
2 73812 1 15695
2 73813 1 15695
2 73814 1 15703
2 73815 1 15703
2 73816 1 15706
2 73817 1 15706
2 73818 1 15706
2 73819 1 15706
2 73820 1 15706
2 73821 1 15706
2 73822 1 15706
2 73823 1 15706
2 73824 1 15706
2 73825 1 15706
2 73826 1 15706
2 73827 1 15706
2 73828 1 15706
2 73829 1 15708
2 73830 1 15708
2 73831 1 15708
2 73832 1 15711
2 73833 1 15711
2 73834 1 15723
2 73835 1 15723
2 73836 1 15724
2 73837 1 15724
2 73838 1 15724
2 73839 1 15724
2 73840 1 15724
2 73841 1 15724
2 73842 1 15724
2 73843 1 15724
2 73844 1 15736
2 73845 1 15736
2 73846 1 15765
2 73847 1 15765
2 73848 1 15778
2 73849 1 15778
2 73850 1 15778
2 73851 1 15783
2 73852 1 15783
2 73853 1 15783
2 73854 1 15788
2 73855 1 15788
2 73856 1 15796
2 73857 1 15796
2 73858 1 15796
2 73859 1 15796
2 73860 1 15796
2 73861 1 15796
2 73862 1 15797
2 73863 1 15797
2 73864 1 15800
2 73865 1 15800
2 73866 1 15803
2 73867 1 15803
2 73868 1 15806
2 73869 1 15806
2 73870 1 15806
2 73871 1 15806
2 73872 1 15825
2 73873 1 15825
2 73874 1 15839
2 73875 1 15839
2 73876 1 15839
2 73877 1 15840
2 73878 1 15840
2 73879 1 15845
2 73880 1 15845
2 73881 1 15857
2 73882 1 15857
2 73883 1 15857
2 73884 1 15858
2 73885 1 15858
2 73886 1 15876
2 73887 1 15876
2 73888 1 15876
2 73889 1 15878
2 73890 1 15878
2 73891 1 15878
2 73892 1 15886
2 73893 1 15886
2 73894 1 15886
2 73895 1 15886
2 73896 1 15888
2 73897 1 15888
2 73898 1 15896
2 73899 1 15896
2 73900 1 15913
2 73901 1 15913
2 73902 1 15914
2 73903 1 15914
2 73904 1 15914
2 73905 1 15934
2 73906 1 15934
2 73907 1 15949
2 73908 1 15949
2 73909 1 15950
2 73910 1 15950
2 73911 1 15984
2 73912 1 15984
2 73913 1 15984
2 73914 1 15984
2 73915 1 15984
2 73916 1 15985
2 73917 1 15985
2 73918 1 15985
2 73919 1 15985
2 73920 1 15985
2 73921 1 15986
2 73922 1 15986
2 73923 1 16008
2 73924 1 16008
2 73925 1 16008
2 73926 1 16009
2 73927 1 16009
2 73928 1 16024
2 73929 1 16024
2 73930 1 16048
2 73931 1 16048
2 73932 1 16051
2 73933 1 16051
2 73934 1 16051
2 73935 1 16058
2 73936 1 16058
2 73937 1 16083
2 73938 1 16083
2 73939 1 16134
2 73940 1 16134
2 73941 1 16146
2 73942 1 16146
2 73943 1 16148
2 73944 1 16148
2 73945 1 16153
2 73946 1 16153
2 73947 1 16153
2 73948 1 16153
2 73949 1 16153
2 73950 1 16153
2 73951 1 16155
2 73952 1 16155
2 73953 1 16160
2 73954 1 16160
2 73955 1 16177
2 73956 1 16177
2 73957 1 16180
2 73958 1 16180
2 73959 1 16189
2 73960 1 16189
2 73961 1 16190
2 73962 1 16190
2 73963 1 16208
2 73964 1 16208
2 73965 1 16208
2 73966 1 16208
2 73967 1 16233
2 73968 1 16233
2 73969 1 16233
2 73970 1 16250
2 73971 1 16250
2 73972 1 16256
2 73973 1 16256
2 73974 1 16256
2 73975 1 16259
2 73976 1 16259
2 73977 1 16277
2 73978 1 16277
2 73979 1 16286
2 73980 1 16286
2 73981 1 16310
2 73982 1 16310
2 73983 1 16368
2 73984 1 16368
2 73985 1 16371
2 73986 1 16371
2 73987 1 16371
2 73988 1 16371
2 73989 1 16382
2 73990 1 16382
2 73991 1 16382
2 73992 1 16383
2 73993 1 16383
2 73994 1 16384
2 73995 1 16384
2 73996 1 16385
2 73997 1 16385
2 73998 1 16385
2 73999 1 16385
2 74000 1 16400
2 74001 1 16400
2 74002 1 16400
2 74003 1 16400
2 74004 1 16401
2 74005 1 16401
2 74006 1 16417
2 74007 1 16417
2 74008 1 16444
2 74009 1 16444
2 74010 1 16445
2 74011 1 16445
2 74012 1 16445
2 74013 1 16446
2 74014 1 16446
2 74015 1 16446
2 74016 1 16446
2 74017 1 16446
2 74018 1 16448
2 74019 1 16448
2 74020 1 16450
2 74021 1 16450
2 74022 1 16451
2 74023 1 16451
2 74024 1 16451
2 74025 1 16456
2 74026 1 16456
2 74027 1 16457
2 74028 1 16457
2 74029 1 16458
2 74030 1 16458
2 74031 1 16460
2 74032 1 16460
2 74033 1 16469
2 74034 1 16469
2 74035 1 16470
2 74036 1 16470
2 74037 1 16471
2 74038 1 16471
2 74039 1 16471
2 74040 1 16473
2 74041 1 16473
2 74042 1 16473
2 74043 1 16476
2 74044 1 16476
2 74045 1 16477
2 74046 1 16477
2 74047 1 16487
2 74048 1 16487
2 74049 1 16487
2 74050 1 16487
2 74051 1 16489
2 74052 1 16489
2 74053 1 16490
2 74054 1 16490
2 74055 1 16491
2 74056 1 16491
2 74057 1 16492
2 74058 1 16492
2 74059 1 16528
2 74060 1 16528
2 74061 1 16532
2 74062 1 16532
2 74063 1 16538
2 74064 1 16538
2 74065 1 16539
2 74066 1 16539
2 74067 1 16546
2 74068 1 16546
2 74069 1 16548
2 74070 1 16548
2 74071 1 16557
2 74072 1 16557
2 74073 1 16557
2 74074 1 16558
2 74075 1 16558
2 74076 1 16558
2 74077 1 16558
2 74078 1 16558
2 74079 1 16559
2 74080 1 16559
2 74081 1 16560
2 74082 1 16560
2 74083 1 16571
2 74084 1 16571
2 74085 1 16572
2 74086 1 16572
2 74087 1 16572
2 74088 1 16572
2 74089 1 16589
2 74090 1 16589
2 74091 1 16604
2 74092 1 16604
2 74093 1 16625
2 74094 1 16625
2 74095 1 16628
2 74096 1 16628
2 74097 1 16633
2 74098 1 16633
2 74099 1 16651
2 74100 1 16651
2 74101 1 16665
2 74102 1 16665
2 74103 1 16666
2 74104 1 16666
2 74105 1 16676
2 74106 1 16676
2 74107 1 16692
2 74108 1 16692
2 74109 1 16694
2 74110 1 16694
2 74111 1 16702
2 74112 1 16702
2 74113 1 16705
2 74114 1 16705
2 74115 1 16736
2 74116 1 16736
2 74117 1 16736
2 74118 1 16771
2 74119 1 16771
2 74120 1 16771
2 74121 1 16779
2 74122 1 16779
2 74123 1 16793
2 74124 1 16793
2 74125 1 16793
2 74126 1 16794
2 74127 1 16794
2 74128 1 16794
2 74129 1 16794
2 74130 1 16821
2 74131 1 16821
2 74132 1 16830
2 74133 1 16830
2 74134 1 16853
2 74135 1 16853
2 74136 1 16853
2 74137 1 16862
2 74138 1 16862
2 74139 1 16866
2 74140 1 16866
2 74141 1 16869
2 74142 1 16869
2 74143 1 16869
2 74144 1 16876
2 74145 1 16876
2 74146 1 16877
2 74147 1 16877
2 74148 1 16888
2 74149 1 16888
2 74150 1 16905
2 74151 1 16905
2 74152 1 16906
2 74153 1 16906
2 74154 1 16919
2 74155 1 16919
2 74156 1 16941
2 74157 1 16941
2 74158 1 16942
2 74159 1 16942
2 74160 1 16942
2 74161 1 16942
2 74162 1 16944
2 74163 1 16944
2 74164 1 16952
2 74165 1 16952
2 74166 1 17000
2 74167 1 17000
2 74168 1 17034
2 74169 1 17034
2 74170 1 17050
2 74171 1 17050
2 74172 1 17064
2 74173 1 17064
2 74174 1 17075
2 74175 1 17075
2 74176 1 17077
2 74177 1 17077
2 74178 1 17090
2 74179 1 17090
2 74180 1 17090
2 74181 1 17144
2 74182 1 17144
2 74183 1 17144
2 74184 1 17144
2 74185 1 17147
2 74186 1 17147
2 74187 1 17147
2 74188 1 17186
2 74189 1 17186
2 74190 1 17186
2 74191 1 17186
2 74192 1 17186
2 74193 1 17187
2 74194 1 17187
2 74195 1 17192
2 74196 1 17192
2 74197 1 17193
2 74198 1 17193
2 74199 1 17193
2 74200 1 17193
2 74201 1 17193
2 74202 1 17196
2 74203 1 17196
2 74204 1 17223
2 74205 1 17223
2 74206 1 17223
2 74207 1 17241
2 74208 1 17241
2 74209 1 17262
2 74210 1 17262
2 74211 1 17270
2 74212 1 17270
2 74213 1 17274
2 74214 1 17274
2 74215 1 17284
2 74216 1 17284
2 74217 1 17288
2 74218 1 17288
2 74219 1 17304
2 74220 1 17304
2 74221 1 17308
2 74222 1 17308
2 74223 1 17309
2 74224 1 17309
2 74225 1 17314
2 74226 1 17314
2 74227 1 17314
2 74228 1 17348
2 74229 1 17348
2 74230 1 17352
2 74231 1 17352
2 74232 1 17353
2 74233 1 17353
2 74234 1 17353
2 74235 1 17353
2 74236 1 17359
2 74237 1 17359
2 74238 1 17360
2 74239 1 17360
2 74240 1 17368
2 74241 1 17368
2 74242 1 17368
2 74243 1 17368
2 74244 1 17368
2 74245 1 17368
2 74246 1 17370
2 74247 1 17370
2 74248 1 17376
2 74249 1 17376
2 74250 1 17376
2 74251 1 17376
2 74252 1 17380
2 74253 1 17380
2 74254 1 17381
2 74255 1 17381
2 74256 1 17387
2 74257 1 17387
2 74258 1 17498
2 74259 1 17498
2 74260 1 17521
2 74261 1 17521
2 74262 1 17534
2 74263 1 17534
2 74264 1 17534
2 74265 1 17534
2 74266 1 17574
2 74267 1 17574
2 74268 1 17574
2 74269 1 17574
2 74270 1 17574
2 74271 1 17574
2 74272 1 17617
2 74273 1 17617
2 74274 1 17643
2 74275 1 17643
2 74276 1 17656
2 74277 1 17656
2 74278 1 17656
2 74279 1 17738
2 74280 1 17738
2 74281 1 17739
2 74282 1 17739
2 74283 1 17755
2 74284 1 17755
2 74285 1 17755
2 74286 1 17755
2 74287 1 17755
2 74288 1 17755
2 74289 1 17755
2 74290 1 17755
2 74291 1 17755
2 74292 1 17755
2 74293 1 17755
2 74294 1 17755
2 74295 1 17755
2 74296 1 17755
2 74297 1 17755
2 74298 1 17755
2 74299 1 17755
2 74300 1 17755
2 74301 1 17755
2 74302 1 17755
2 74303 1 17757
2 74304 1 17757
2 74305 1 17779
2 74306 1 17779
2 74307 1 17838
2 74308 1 17838
2 74309 1 17838
2 74310 1 17838
2 74311 1 17839
2 74312 1 17839
2 74313 1 17848
2 74314 1 17848
2 74315 1 17895
2 74316 1 17895
2 74317 1 17895
2 74318 1 17899
2 74319 1 17899
2 74320 1 17900
2 74321 1 17900
2 74322 1 17911
2 74323 1 17911
2 74324 1 17916
2 74325 1 17916
2 74326 1 17940
2 74327 1 17940
2 74328 1 17951
2 74329 1 17951
2 74330 1 17993
2 74331 1 17993
2 74332 1 18011
2 74333 1 18011
2 74334 1 18050
2 74335 1 18050
2 74336 1 18050
2 74337 1 18050
2 74338 1 18050
2 74339 1 18050
2 74340 1 18052
2 74341 1 18052
2 74342 1 18065
2 74343 1 18065
2 74344 1 18069
2 74345 1 18069
2 74346 1 18070
2 74347 1 18070
2 74348 1 18070
2 74349 1 18070
2 74350 1 18077
2 74351 1 18077
2 74352 1 18078
2 74353 1 18078
2 74354 1 18082
2 74355 1 18082
2 74356 1 18083
2 74357 1 18083
2 74358 1 18083
2 74359 1 18083
2 74360 1 18083
2 74361 1 18084
2 74362 1 18084
2 74363 1 18110
2 74364 1 18110
2 74365 1 18130
2 74366 1 18130
2 74367 1 18137
2 74368 1 18137
2 74369 1 18137
2 74370 1 18145
2 74371 1 18145
2 74372 1 18146
2 74373 1 18146
2 74374 1 18154
2 74375 1 18154
2 74376 1 18154
2 74377 1 18166
2 74378 1 18166
2 74379 1 18232
2 74380 1 18232
2 74381 1 18232
2 74382 1 18232
2 74383 1 18235
2 74384 1 18235
2 74385 1 18242
2 74386 1 18242
2 74387 1 18253
2 74388 1 18253
2 74389 1 18255
2 74390 1 18255
2 74391 1 18338
2 74392 1 18338
2 74393 1 18338
2 74394 1 18347
2 74395 1 18347
2 74396 1 18347
2 74397 1 18350
2 74398 1 18350
2 74399 1 18350
2 74400 1 18350
2 74401 1 18359
2 74402 1 18359
2 74403 1 18359
2 74404 1 18361
2 74405 1 18361
2 74406 1 18362
2 74407 1 18362
2 74408 1 18390
2 74409 1 18390
2 74410 1 18392
2 74411 1 18392
2 74412 1 18400
2 74413 1 18400
2 74414 1 18400
2 74415 1 18400
2 74416 1 18400
2 74417 1 18400
2 74418 1 18420
2 74419 1 18420
2 74420 1 18428
2 74421 1 18428
2 74422 1 18428
2 74423 1 18463
2 74424 1 18463
2 74425 1 18463
2 74426 1 18463
2 74427 1 18463
2 74428 1 18493
2 74429 1 18493
2 74430 1 18515
2 74431 1 18515
2 74432 1 18515
2 74433 1 18515
2 74434 1 18515
2 74435 1 18515
2 74436 1 18540
2 74437 1 18540
2 74438 1 18540
2 74439 1 18567
2 74440 1 18567
2 74441 1 18567
2 74442 1 18583
2 74443 1 18583
2 74444 1 18612
2 74445 1 18612
2 74446 1 18612
2 74447 1 18636
2 74448 1 18636
2 74449 1 18650
2 74450 1 18650
2 74451 1 18650
2 74452 1 18658
2 74453 1 18658
2 74454 1 18658
2 74455 1 18659
2 74456 1 18659
2 74457 1 18666
2 74458 1 18666
2 74459 1 18666
2 74460 1 18666
2 74461 1 18666
2 74462 1 18682
2 74463 1 18682
2 74464 1 18687
2 74465 1 18687
2 74466 1 18699
2 74467 1 18699
2 74468 1 18699
2 74469 1 18699
2 74470 1 18707
2 74471 1 18707
2 74472 1 18708
2 74473 1 18708
2 74474 1 18709
2 74475 1 18709
2 74476 1 18711
2 74477 1 18711
2 74478 1 18719
2 74479 1 18719
2 74480 1 18728
2 74481 1 18728
2 74482 1 18728
2 74483 1 18729
2 74484 1 18729
2 74485 1 18739
2 74486 1 18739
2 74487 1 18753
2 74488 1 18753
2 74489 1 18754
2 74490 1 18754
2 74491 1 18754
2 74492 1 18781
2 74493 1 18781
2 74494 1 18781
2 74495 1 18815
2 74496 1 18815
2 74497 1 18823
2 74498 1 18823
2 74499 1 18831
2 74500 1 18831
2 74501 1 18890
2 74502 1 18890
2 74503 1 18895
2 74504 1 18895
2 74505 1 18896
2 74506 1 18896
2 74507 1 18916
2 74508 1 18916
2 74509 1 18917
2 74510 1 18917
2 74511 1 18918
2 74512 1 18918
2 74513 1 18918
2 74514 1 18925
2 74515 1 18925
2 74516 1 18925
2 74517 1 18953
2 74518 1 18953
2 74519 1 18953
2 74520 1 18957
2 74521 1 18957
2 74522 1 18964
2 74523 1 18964
2 74524 1 18990
2 74525 1 18990
2 74526 1 18990
2 74527 1 18990
2 74528 1 19005
2 74529 1 19005
2 74530 1 19005
2 74531 1 19009
2 74532 1 19009
2 74533 1 19022
2 74534 1 19022
2 74535 1 19023
2 74536 1 19023
2 74537 1 19029
2 74538 1 19029
2 74539 1 19049
2 74540 1 19049
2 74541 1 19062
2 74542 1 19062
2 74543 1 19113
2 74544 1 19113
2 74545 1 19115
2 74546 1 19115
2 74547 1 19115
2 74548 1 19115
2 74549 1 19146
2 74550 1 19146
2 74551 1 19148
2 74552 1 19148
2 74553 1 19178
2 74554 1 19178
2 74555 1 19187
2 74556 1 19187
2 74557 1 19189
2 74558 1 19189
2 74559 1 19223
2 74560 1 19223
2 74561 1 19256
2 74562 1 19256
2 74563 1 19256
2 74564 1 19259
2 74565 1 19259
2 74566 1 19263
2 74567 1 19263
2 74568 1 19263
2 74569 1 19263
2 74570 1 19264
2 74571 1 19264
2 74572 1 19264
2 74573 1 19269
2 74574 1 19269
2 74575 1 19270
2 74576 1 19270
2 74577 1 19271
2 74578 1 19271
2 74579 1 19273
2 74580 1 19273
2 74581 1 19273
2 74582 1 19273
2 74583 1 19273
2 74584 1 19273
2 74585 1 19273
2 74586 1 19273
2 74587 1 19281
2 74588 1 19281
2 74589 1 19284
2 74590 1 19284
2 74591 1 19284
2 74592 1 19299
2 74593 1 19299
2 74594 1 19302
2 74595 1 19302
2 74596 1 19315
2 74597 1 19315
2 74598 1 19316
2 74599 1 19316
2 74600 1 19316
2 74601 1 19335
2 74602 1 19335
2 74603 1 19336
2 74604 1 19336
2 74605 1 19338
2 74606 1 19338
2 74607 1 19341
2 74608 1 19341
2 74609 1 19351
2 74610 1 19351
2 74611 1 19351
2 74612 1 19351
2 74613 1 19366
2 74614 1 19366
2 74615 1 19366
2 74616 1 19367
2 74617 1 19367
2 74618 1 19407
2 74619 1 19407
2 74620 1 19446
2 74621 1 19446
2 74622 1 19460
2 74623 1 19460
2 74624 1 19481
2 74625 1 19481
2 74626 1 19545
2 74627 1 19545
2 74628 1 19545
2 74629 1 19569
2 74630 1 19569
2 74631 1 19589
2 74632 1 19589
2 74633 1 19590
2 74634 1 19590
2 74635 1 19590
2 74636 1 19590
2 74637 1 19590
2 74638 1 19590
2 74639 1 19626
2 74640 1 19626
2 74641 1 19644
2 74642 1 19644
2 74643 1 19644
2 74644 1 19756
2 74645 1 19756
2 74646 1 19777
2 74647 1 19777
2 74648 1 19813
2 74649 1 19813
2 74650 1 19834
2 74651 1 19834
2 74652 1 19868
2 74653 1 19868
2 74654 1 19885
2 74655 1 19885
2 74656 1 19899
2 74657 1 19899
2 74658 1 19933
2 74659 1 19933
2 74660 1 19933
2 74661 1 19933
2 74662 1 19933
2 74663 1 20002
2 74664 1 20002
2 74665 1 20002
2 74666 1 20027
2 74667 1 20027
2 74668 1 20055
2 74669 1 20055
2 74670 1 20063
2 74671 1 20063
2 74672 1 20063
2 74673 1 20075
2 74674 1 20075
2 74675 1 20102
2 74676 1 20102
2 74677 1 20110
2 74678 1 20110
2 74679 1 20120
2 74680 1 20120
2 74681 1 20128
2 74682 1 20128
2 74683 1 20132
2 74684 1 20132
2 74685 1 20132
2 74686 1 20153
2 74687 1 20153
2 74688 1 20186
2 74689 1 20186
2 74690 1 20186
2 74691 1 20210
2 74692 1 20210
2 74693 1 20227
2 74694 1 20227
2 74695 1 20234
2 74696 1 20234
2 74697 1 20253
2 74698 1 20253
2 74699 1 20265
2 74700 1 20265
2 74701 1 20265
2 74702 1 20272
2 74703 1 20272
2 74704 1 20311
2 74705 1 20311
2 74706 1 20323
2 74707 1 20323
2 74708 1 20331
2 74709 1 20331
2 74710 1 20334
2 74711 1 20334
2 74712 1 20364
2 74713 1 20364
2 74714 1 20367
2 74715 1 20367
2 74716 1 20367
2 74717 1 20367
2 74718 1 20369
2 74719 1 20369
2 74720 1 20369
2 74721 1 20374
2 74722 1 20374
2 74723 1 20378
2 74724 1 20378
2 74725 1 20379
2 74726 1 20379
2 74727 1 20391
2 74728 1 20391
2 74729 1 20435
2 74730 1 20435
2 74731 1 20438
2 74732 1 20438
2 74733 1 20439
2 74734 1 20439
2 74735 1 20446
2 74736 1 20446
2 74737 1 20447
2 74738 1 20447
2 74739 1 20475
2 74740 1 20475
2 74741 1 20508
2 74742 1 20508
2 74743 1 20533
2 74744 1 20533
2 74745 1 20584
2 74746 1 20584
2 74747 1 20587
2 74748 1 20587
2 74749 1 20599
2 74750 1 20599
2 74751 1 20604
2 74752 1 20604
2 74753 1 20604
2 74754 1 20604
2 74755 1 20604
2 74756 1 20604
2 74757 1 20607
2 74758 1 20607
2 74759 1 20607
2 74760 1 20607
2 74761 1 20608
2 74762 1 20608
2 74763 1 20609
2 74764 1 20609
2 74765 1 20617
2 74766 1 20617
2 74767 1 20618
2 74768 1 20618
2 74769 1 20618
2 74770 1 20618
2 74771 1 20655
2 74772 1 20655
2 74773 1 20661
2 74774 1 20661
2 74775 1 20676
2 74776 1 20676
2 74777 1 20677
2 74778 1 20677
2 74779 1 20677
2 74780 1 20687
2 74781 1 20687
2 74782 1 20703
2 74783 1 20703
2 74784 1 20705
2 74785 1 20705
2 74786 1 20722
2 74787 1 20722
2 74788 1 20730
2 74789 1 20730
2 74790 1 20739
2 74791 1 20739
2 74792 1 20739
2 74793 1 20740
2 74794 1 20740
2 74795 1 20744
2 74796 1 20744
2 74797 1 20749
2 74798 1 20749
2 74799 1 20749
2 74800 1 20813
2 74801 1 20813
2 74802 1 20813
2 74803 1 20817
2 74804 1 20817
2 74805 1 20819
2 74806 1 20819
2 74807 1 20822
2 74808 1 20822
2 74809 1 20828
2 74810 1 20828
2 74811 1 20851
2 74812 1 20851
2 74813 1 20873
2 74814 1 20873
2 74815 1 20874
2 74816 1 20874
2 74817 1 20906
2 74818 1 20906
2 74819 1 20909
2 74820 1 20909
2 74821 1 20909
2 74822 1 20909
2 74823 1 20936
2 74824 1 20936
2 74825 1 20944
2 74826 1 20944
2 74827 1 20950
2 74828 1 20950
2 74829 1 20967
2 74830 1 20967
2 74831 1 20967
2 74832 1 20967
2 74833 1 20967
2 74834 1 20967
2 74835 1 20967
2 74836 1 20967
2 74837 1 20967
2 74838 1 20967
2 74839 1 20968
2 74840 1 20968
2 74841 1 20968
2 74842 1 20968
2 74843 1 20982
2 74844 1 20982
2 74845 1 20987
2 74846 1 20987
2 74847 1 20987
2 74848 1 20990
2 74849 1 20990
2 74850 1 20991
2 74851 1 20991
2 74852 1 20995
2 74853 1 20995
2 74854 1 21025
2 74855 1 21025
2 74856 1 21026
2 74857 1 21026
2 74858 1 21035
2 74859 1 21035
2 74860 1 21035
2 74861 1 21036
2 74862 1 21036
2 74863 1 21045
2 74864 1 21045
2 74865 1 21076
2 74866 1 21076
2 74867 1 21104
2 74868 1 21104
2 74869 1 21105
2 74870 1 21105
2 74871 1 21108
2 74872 1 21108
2 74873 1 21108
2 74874 1 21108
2 74875 1 21114
2 74876 1 21114
2 74877 1 21117
2 74878 1 21117
2 74879 1 21118
2 74880 1 21118
2 74881 1 21129
2 74882 1 21129
2 74883 1 21138
2 74884 1 21138
2 74885 1 21139
2 74886 1 21139
2 74887 1 21139
2 74888 1 21139
2 74889 1 21139
2 74890 1 21139
2 74891 1 21141
2 74892 1 21141
2 74893 1 21153
2 74894 1 21153
2 74895 1 21156
2 74896 1 21156
2 74897 1 21156
2 74898 1 21157
2 74899 1 21157
2 74900 1 21160
2 74901 1 21160
2 74902 1 21161
2 74903 1 21161
2 74904 1 21161
2 74905 1 21169
2 74906 1 21169
2 74907 1 21170
2 74908 1 21170
2 74909 1 21170
2 74910 1 21176
2 74911 1 21176
2 74912 1 21179
2 74913 1 21179
2 74914 1 21183
2 74915 1 21183
2 74916 1 21184
2 74917 1 21184
2 74918 1 21184
2 74919 1 21184
2 74920 1 21184
2 74921 1 21184
2 74922 1 21195
2 74923 1 21195
2 74924 1 21223
2 74925 1 21223
2 74926 1 21223
2 74927 1 21231
2 74928 1 21231
2 74929 1 21238
2 74930 1 21238
2 74931 1 21249
2 74932 1 21249
2 74933 1 21251
2 74934 1 21251
2 74935 1 21251
2 74936 1 21252
2 74937 1 21252
2 74938 1 21256
2 74939 1 21256
2 74940 1 21256
2 74941 1 21266
2 74942 1 21266
2 74943 1 21266
2 74944 1 21273
2 74945 1 21273
2 74946 1 21273
2 74947 1 21280
2 74948 1 21280
2 74949 1 21292
2 74950 1 21292
2 74951 1 21295
2 74952 1 21295
2 74953 1 21298
2 74954 1 21298
2 74955 1 21301
2 74956 1 21301
2 74957 1 21302
2 74958 1 21302
2 74959 1 21305
2 74960 1 21305
2 74961 1 21308
2 74962 1 21308
2 74963 1 21308
2 74964 1 21309
2 74965 1 21309
2 74966 1 21309
2 74967 1 21309
2 74968 1 21354
2 74969 1 21354
2 74970 1 21355
2 74971 1 21355
2 74972 1 21355
2 74973 1 21355
2 74974 1 21357
2 74975 1 21357
2 74976 1 21362
2 74977 1 21362
2 74978 1 21372
2 74979 1 21372
2 74980 1 21375
2 74981 1 21375
2 74982 1 21376
2 74983 1 21376
2 74984 1 21388
2 74985 1 21388
2 74986 1 21401
2 74987 1 21401
2 74988 1 21403
2 74989 1 21403
2 74990 1 21415
2 74991 1 21415
2 74992 1 21415
2 74993 1 21416
2 74994 1 21416
2 74995 1 21416
2 74996 1 21416
2 74997 1 21448
2 74998 1 21448
2 74999 1 21452
2 75000 1 21452
2 75001 1 21470
2 75002 1 21470
2 75003 1 21470
2 75004 1 21470
2 75005 1 21470
2 75006 1 21482
2 75007 1 21482
2 75008 1 21496
2 75009 1 21496
2 75010 1 21508
2 75011 1 21508
2 75012 1 21543
2 75013 1 21543
2 75014 1 21543
2 75015 1 21557
2 75016 1 21557
2 75017 1 21570
2 75018 1 21570
2 75019 1 21570
2 75020 1 21571
2 75021 1 21571
2 75022 1 21571
2 75023 1 21572
2 75024 1 21572
2 75025 1 21584
2 75026 1 21584
2 75027 1 21588
2 75028 1 21588
2 75029 1 21625
2 75030 1 21625
2 75031 1 21653
2 75032 1 21653
2 75033 1 21672
2 75034 1 21672
2 75035 1 21672
2 75036 1 21681
2 75037 1 21681
2 75038 1 21682
2 75039 1 21682
2 75040 1 21682
2 75041 1 21682
2 75042 1 21682
2 75043 1 21709
2 75044 1 21709
2 75045 1 21712
2 75046 1 21712
2 75047 1 21714
2 75048 1 21714
2 75049 1 21725
2 75050 1 21725
2 75051 1 21725
2 75052 1 21770
2 75053 1 21770
2 75054 1 21801
2 75055 1 21801
2 75056 1 21826
2 75057 1 21826
2 75058 1 21826
2 75059 1 21826
2 75060 1 21827
2 75061 1 21827
2 75062 1 21827
2 75063 1 21828
2 75064 1 21828
2 75065 1 21828
2 75066 1 21828
2 75067 1 21829
2 75068 1 21829
2 75069 1 21832
2 75070 1 21832
2 75071 1 21832
2 75072 1 21860
2 75073 1 21860
2 75074 1 21880
2 75075 1 21880
2 75076 1 21896
2 75077 1 21896
2 75078 1 21910
2 75079 1 21910
2 75080 1 21926
2 75081 1 21926
2 75082 1 21935
2 75083 1 21935
2 75084 1 21935
2 75085 1 21935
2 75086 1 21979
2 75087 1 21979
2 75088 1 21998
2 75089 1 21998
2 75090 1 21999
2 75091 1 21999
2 75092 1 22000
2 75093 1 22000
2 75094 1 22000
2 75095 1 22000
2 75096 1 22000
2 75097 1 22000
2 75098 1 22000
2 75099 1 22002
2 75100 1 22002
2 75101 1 22002
2 75102 1 22002
2 75103 1 22002
2 75104 1 22041
2 75105 1 22041
2 75106 1 22041
2 75107 1 22041
2 75108 1 22041
2 75109 1 22041
2 75110 1 22041
2 75111 1 22041
2 75112 1 22041
2 75113 1 22041
2 75114 1 22041
2 75115 1 22041
2 75116 1 22042
2 75117 1 22042
2 75118 1 22043
2 75119 1 22043
2 75120 1 22093
2 75121 1 22093
2 75122 1 22093
2 75123 1 22093
2 75124 1 22093
2 75125 1 22093
2 75126 1 22094
2 75127 1 22094
2 75128 1 22095
2 75129 1 22095
2 75130 1 22126
2 75131 1 22126
2 75132 1 22126
2 75133 1 22137
2 75134 1 22137
2 75135 1 22137
2 75136 1 22140
2 75137 1 22140
2 75138 1 22153
2 75139 1 22153
2 75140 1 22153
2 75141 1 22153
2 75142 1 22157
2 75143 1 22157
2 75144 1 22158
2 75145 1 22158
2 75146 1 22158
2 75147 1 22166
2 75148 1 22166
2 75149 1 22182
2 75150 1 22182
2 75151 1 22209
2 75152 1 22209
2 75153 1 22247
2 75154 1 22247
2 75155 1 22247
2 75156 1 22247
2 75157 1 22247
2 75158 1 22247
2 75159 1 22248
2 75160 1 22248
2 75161 1 22256
2 75162 1 22256
2 75163 1 22274
2 75164 1 22274
2 75165 1 22277
2 75166 1 22277
2 75167 1 22277
2 75168 1 22277
2 75169 1 22279
2 75170 1 22279
2 75171 1 22279
2 75172 1 22279
2 75173 1 22298
2 75174 1 22298
2 75175 1 22310
2 75176 1 22310
2 75177 1 22332
2 75178 1 22332
2 75179 1 22354
2 75180 1 22354
2 75181 1 22354
2 75182 1 22354
2 75183 1 22354
2 75184 1 22354
2 75185 1 22355
2 75186 1 22355
2 75187 1 22365
2 75188 1 22365
2 75189 1 22377
2 75190 1 22377
2 75191 1 22378
2 75192 1 22378
2 75193 1 22384
2 75194 1 22384
2 75195 1 22385
2 75196 1 22385
2 75197 1 22400
2 75198 1 22400
2 75199 1 22400
2 75200 1 22400
2 75201 1 22400
2 75202 1 22400
2 75203 1 22456
2 75204 1 22456
2 75205 1 22458
2 75206 1 22458
2 75207 1 22459
2 75208 1 22459
2 75209 1 22460
2 75210 1 22460
2 75211 1 22460
2 75212 1 22460
2 75213 1 22460
2 75214 1 22460
2 75215 1 22460
2 75216 1 22461
2 75217 1 22461
2 75218 1 22469
2 75219 1 22469
2 75220 1 22475
2 75221 1 22475
2 75222 1 22483
2 75223 1 22483
2 75224 1 22488
2 75225 1 22488
2 75226 1 22488
2 75227 1 22488
2 75228 1 22488
2 75229 1 22488
2 75230 1 22488
2 75231 1 22488
2 75232 1 22488
2 75233 1 22489
2 75234 1 22489
2 75235 1 22489
2 75236 1 22490
2 75237 1 22490
2 75238 1 22490
2 75239 1 22490
2 75240 1 22490
2 75241 1 22490
2 75242 1 22490
2 75243 1 22490
2 75244 1 22490
2 75245 1 22490
2 75246 1 22490
2 75247 1 22491
2 75248 1 22491
2 75249 1 22491
2 75250 1 22491
2 75251 1 22491
2 75252 1 22491
2 75253 1 22491
2 75254 1 22491
2 75255 1 22491
2 75256 1 22493
2 75257 1 22493
2 75258 1 22493
2 75259 1 22493
2 75260 1 22493
2 75261 1 22493
2 75262 1 22493
2 75263 1 22494
2 75264 1 22494
2 75265 1 22496
2 75266 1 22496
2 75267 1 22498
2 75268 1 22498
2 75269 1 22498
2 75270 1 22498
2 75271 1 22499
2 75272 1 22499
2 75273 1 22499
2 75274 1 22499
2 75275 1 22499
2 75276 1 22499
2 75277 1 22499
2 75278 1 22499
2 75279 1 22499
2 75280 1 22499
2 75281 1 22499
2 75282 1 22499
2 75283 1 22499
2 75284 1 22499
2 75285 1 22499
2 75286 1 22499
2 75287 1 22499
2 75288 1 22499
2 75289 1 22499
2 75290 1 22499
2 75291 1 22499
2 75292 1 22499
2 75293 1 22499
2 75294 1 22499
2 75295 1 22499
2 75296 1 22499
2 75297 1 22500
2 75298 1 22500
2 75299 1 22506
2 75300 1 22506
2 75301 1 22506
2 75302 1 22506
2 75303 1 22506
2 75304 1 22508
2 75305 1 22508
2 75306 1 22508
2 75307 1 22509
2 75308 1 22509
2 75309 1 22509
2 75310 1 22509
2 75311 1 22516
2 75312 1 22516
2 75313 1 22516
2 75314 1 22524
2 75315 1 22524
2 75316 1 22524
2 75317 1 22525
2 75318 1 22525
2 75319 1 22530
2 75320 1 22530
2 75321 1 22534
2 75322 1 22534
2 75323 1 22536
2 75324 1 22536
2 75325 1 22546
2 75326 1 22546
2 75327 1 22548
2 75328 1 22548
2 75329 1 22555
2 75330 1 22555
2 75331 1 22555
2 75332 1 22555
2 75333 1 22555
2 75334 1 22556
2 75335 1 22556
2 75336 1 22556
2 75337 1 22556
2 75338 1 22557
2 75339 1 22557
2 75340 1 22557
2 75341 1 22557
2 75342 1 22566
2 75343 1 22566
2 75344 1 22566
2 75345 1 22566
2 75346 1 22566
2 75347 1 22566
2 75348 1 22566
2 75349 1 22577
2 75350 1 22577
2 75351 1 22577
2 75352 1 22577
2 75353 1 22577
2 75354 1 22577
2 75355 1 22577
2 75356 1 22577
2 75357 1 22586
2 75358 1 22586
2 75359 1 22586
2 75360 1 22586
2 75361 1 22586
2 75362 1 22586
2 75363 1 22587
2 75364 1 22587
2 75365 1 22587
2 75366 1 22589
2 75367 1 22589
2 75368 1 22593
2 75369 1 22593
2 75370 1 22593
2 75371 1 22608
2 75372 1 22608
2 75373 1 22616
2 75374 1 22616
2 75375 1 22616
2 75376 1 22616
2 75377 1 22638
2 75378 1 22638
2 75379 1 22650
2 75380 1 22650
2 75381 1 22650
2 75382 1 22650
2 75383 1 22651
2 75384 1 22651
2 75385 1 22651
2 75386 1 22651
2 75387 1 22651
2 75388 1 22654
2 75389 1 22654
2 75390 1 22655
2 75391 1 22655
2 75392 1 22655
2 75393 1 22688
2 75394 1 22688
2 75395 1 22689
2 75396 1 22689
2 75397 1 22689
2 75398 1 22690
2 75399 1 22690
2 75400 1 22690
2 75401 1 22707
2 75402 1 22707
2 75403 1 22710
2 75404 1 22710
2 75405 1 22714
2 75406 1 22714
2 75407 1 22714
2 75408 1 22714
2 75409 1 22714
2 75410 1 22717
2 75411 1 22717
2 75412 1 22717
2 75413 1 22718
2 75414 1 22718
2 75415 1 22718
2 75416 1 22718
2 75417 1 22718
2 75418 1 22728
2 75419 1 22728
2 75420 1 22743
2 75421 1 22743
2 75422 1 22755
2 75423 1 22755
2 75424 1 22755
2 75425 1 22755
2 75426 1 22755
2 75427 1 22755
2 75428 1 22755
2 75429 1 22757
2 75430 1 22757
2 75431 1 22764
2 75432 1 22764
2 75433 1 22764
2 75434 1 22764
2 75435 1 22764
2 75436 1 22764
2 75437 1 22764
2 75438 1 22764
2 75439 1 22764
2 75440 1 22764
2 75441 1 22764
2 75442 1 22764
2 75443 1 22764
2 75444 1 22764
2 75445 1 22764
2 75446 1 22765
2 75447 1 22765
2 75448 1 22765
2 75449 1 22765
2 75450 1 22765
2 75451 1 22766
2 75452 1 22766
2 75453 1 22768
2 75454 1 22768
2 75455 1 22778
2 75456 1 22778
2 75457 1 22795
2 75458 1 22795
2 75459 1 22796
2 75460 1 22796
2 75461 1 22796
2 75462 1 22810
2 75463 1 22810
2 75464 1 22829
2 75465 1 22829
2 75466 1 22829
2 75467 1 22829
2 75468 1 22829
2 75469 1 22829
2 75470 1 22833
2 75471 1 22833
2 75472 1 22843
2 75473 1 22843
2 75474 1 22871
2 75475 1 22871
2 75476 1 22877
2 75477 1 22877
2 75478 1 22877
2 75479 1 22877
2 75480 1 22877
2 75481 1 22881
2 75482 1 22881
2 75483 1 22881
2 75484 1 22881
2 75485 1 22881
2 75486 1 22881
2 75487 1 22881
2 75488 1 22881
2 75489 1 22881
2 75490 1 22881
2 75491 1 22881
2 75492 1 22881
2 75493 1 22883
2 75494 1 22883
2 75495 1 22883
2 75496 1 22883
2 75497 1 22890
2 75498 1 22890
2 75499 1 22890
2 75500 1 22890
2 75501 1 22890
2 75502 1 22890
2 75503 1 22890
2 75504 1 22890
2 75505 1 22890
2 75506 1 22891
2 75507 1 22891
2 75508 1 22891
2 75509 1 22891
2 75510 1 22891
2 75511 1 22891
2 75512 1 22891
2 75513 1 22892
2 75514 1 22892
2 75515 1 22892
2 75516 1 22892
2 75517 1 22892
2 75518 1 22892
2 75519 1 22892
2 75520 1 22892
2 75521 1 22892
2 75522 1 22893
2 75523 1 22893
2 75524 1 22893
2 75525 1 22893
2 75526 1 22893
2 75527 1 22894
2 75528 1 22894
2 75529 1 22897
2 75530 1 22897
2 75531 1 22912
2 75532 1 22912
2 75533 1 22912
2 75534 1 22912
2 75535 1 22912
2 75536 1 22924
2 75537 1 22924
2 75538 1 22931
2 75539 1 22931
2 75540 1 22969
2 75541 1 22969
2 75542 1 22969
2 75543 1 22969
2 75544 1 22969
2 75545 1 22969
2 75546 1 22970
2 75547 1 22970
2 75548 1 22970
2 75549 1 22970
2 75550 1 22972
2 75551 1 22972
2 75552 1 22975
2 75553 1 22975
2 75554 1 22975
2 75555 1 23000
2 75556 1 23000
2 75557 1 23000
2 75558 1 23015
2 75559 1 23015
2 75560 1 23045
2 75561 1 23045
2 75562 1 23045
2 75563 1 23045
2 75564 1 23047
2 75565 1 23047
2 75566 1 23050
2 75567 1 23050
2 75568 1 23050
2 75569 1 23051
2 75570 1 23051
2 75571 1 23052
2 75572 1 23052
2 75573 1 23052
2 75574 1 23065
2 75575 1 23065
2 75576 1 23080
2 75577 1 23080
2 75578 1 23087
2 75579 1 23087
2 75580 1 23095
2 75581 1 23095
2 75582 1 23095
2 75583 1 23095
2 75584 1 23095
2 75585 1 23103
2 75586 1 23103
2 75587 1 23107
2 75588 1 23107
2 75589 1 23110
2 75590 1 23110
2 75591 1 23111
2 75592 1 23111
2 75593 1 23111
2 75594 1 23133
2 75595 1 23133
2 75596 1 23134
2 75597 1 23134
2 75598 1 23135
2 75599 1 23135
2 75600 1 23137
2 75601 1 23137
2 75602 1 23137
2 75603 1 23143
2 75604 1 23143
2 75605 1 23161
2 75606 1 23161
2 75607 1 23164
2 75608 1 23164
2 75609 1 23170
2 75610 1 23170
2 75611 1 23176
2 75612 1 23176
2 75613 1 23190
2 75614 1 23190
2 75615 1 23194
2 75616 1 23194
2 75617 1 23194
2 75618 1 23194
2 75619 1 23194
2 75620 1 23205
2 75621 1 23205
2 75622 1 23206
2 75623 1 23206
2 75624 1 23206
2 75625 1 23206
2 75626 1 23206
2 75627 1 23207
2 75628 1 23207
2 75629 1 23207
2 75630 1 23207
2 75631 1 23229
2 75632 1 23229
2 75633 1 23229
2 75634 1 23238
2 75635 1 23238
2 75636 1 23238
2 75637 1 23238
2 75638 1 23242
2 75639 1 23242
2 75640 1 23243
2 75641 1 23243
2 75642 1 23243
2 75643 1 23243
2 75644 1 23259
2 75645 1 23259
2 75646 1 23259
2 75647 1 23259
2 75648 1 23260
2 75649 1 23260
2 75650 1 23268
2 75651 1 23268
2 75652 1 23272
2 75653 1 23272
2 75654 1 23272
2 75655 1 23272
2 75656 1 23272
2 75657 1 23284
2 75658 1 23284
2 75659 1 23284
2 75660 1 23284
2 75661 1 23288
2 75662 1 23288
2 75663 1 23319
2 75664 1 23319
2 75665 1 23328
2 75666 1 23328
2 75667 1 23337
2 75668 1 23337
2 75669 1 23337
2 75670 1 23337
2 75671 1 23337
2 75672 1 23337
2 75673 1 23337
2 75674 1 23339
2 75675 1 23339
2 75676 1 23339
2 75677 1 23346
2 75678 1 23346
2 75679 1 23346
2 75680 1 23346
2 75681 1 23346
2 75682 1 23346
2 75683 1 23346
2 75684 1 23346
2 75685 1 23346
2 75686 1 23346
2 75687 1 23354
2 75688 1 23354
2 75689 1 23355
2 75690 1 23355
2 75691 1 23357
2 75692 1 23357
2 75693 1 23361
2 75694 1 23361
2 75695 1 23361
2 75696 1 23361
2 75697 1 23361
2 75698 1 23364
2 75699 1 23364
2 75700 1 23364
2 75701 1 23365
2 75702 1 23365
2 75703 1 23365
2 75704 1 23373
2 75705 1 23373
2 75706 1 23376
2 75707 1 23376
2 75708 1 23377
2 75709 1 23377
2 75710 1 23378
2 75711 1 23378
2 75712 1 23405
2 75713 1 23405
2 75714 1 23406
2 75715 1 23406
2 75716 1 23408
2 75717 1 23408
2 75718 1 23416
2 75719 1 23416
2 75720 1 23416
2 75721 1 23416
2 75722 1 23416
2 75723 1 23416
2 75724 1 23424
2 75725 1 23424
2 75726 1 23426
2 75727 1 23426
2 75728 1 23426
2 75729 1 23436
2 75730 1 23436
2 75731 1 23436
2 75732 1 23437
2 75733 1 23437
2 75734 1 23448
2 75735 1 23448
2 75736 1 23452
2 75737 1 23452
2 75738 1 23452
2 75739 1 23453
2 75740 1 23453
2 75741 1 23464
2 75742 1 23464
2 75743 1 23464
2 75744 1 23479
2 75745 1 23479
2 75746 1 23479
2 75747 1 23479
2 75748 1 23481
2 75749 1 23481
2 75750 1 23503
2 75751 1 23503
2 75752 1 23506
2 75753 1 23506
2 75754 1 23507
2 75755 1 23507
2 75756 1 23507
2 75757 1 23507
2 75758 1 23507
2 75759 1 23507
2 75760 1 23507
2 75761 1 23507
2 75762 1 23507
2 75763 1 23507
2 75764 1 23507
2 75765 1 23507
2 75766 1 23509
2 75767 1 23509
2 75768 1 23509
2 75769 1 23516
2 75770 1 23516
2 75771 1 23516
2 75772 1 23517
2 75773 1 23517
2 75774 1 23517
2 75775 1 23517
2 75776 1 23517
2 75777 1 23517
2 75778 1 23520
2 75779 1 23520
2 75780 1 23533
2 75781 1 23533
2 75782 1 23533
2 75783 1 23533
2 75784 1 23559
2 75785 1 23559
2 75786 1 23559
2 75787 1 23559
2 75788 1 23559
2 75789 1 23579
2 75790 1 23579
2 75791 1 23579
2 75792 1 23579
2 75793 1 23581
2 75794 1 23581
2 75795 1 23597
2 75796 1 23597
2 75797 1 23599
2 75798 1 23599
2 75799 1 23600
2 75800 1 23600
2 75801 1 23602
2 75802 1 23602
2 75803 1 23602
2 75804 1 23602
2 75805 1 23603
2 75806 1 23603
2 75807 1 23610
2 75808 1 23610
2 75809 1 23610
2 75810 1 23610
2 75811 1 23610
2 75812 1 23610
2 75813 1 23610
2 75814 1 23610
2 75815 1 23610
2 75816 1 23610
2 75817 1 23610
2 75818 1 23612
2 75819 1 23612
2 75820 1 23613
2 75821 1 23613
2 75822 1 23613
2 75823 1 23613
2 75824 1 23613
2 75825 1 23614
2 75826 1 23614
2 75827 1 23614
2 75828 1 23614
2 75829 1 23614
2 75830 1 23621
2 75831 1 23621
2 75832 1 23621
2 75833 1 23621
2 75834 1 23621
2 75835 1 23634
2 75836 1 23634
2 75837 1 23634
2 75838 1 23634
2 75839 1 23634
2 75840 1 23647
2 75841 1 23647
2 75842 1 23650
2 75843 1 23650
2 75844 1 23653
2 75845 1 23653
2 75846 1 23656
2 75847 1 23656
2 75848 1 23659
2 75849 1 23659
2 75850 1 23659
2 75851 1 23659
2 75852 1 23661
2 75853 1 23661
2 75854 1 23661
2 75855 1 23661
2 75856 1 23662
2 75857 1 23662
2 75858 1 23662
2 75859 1 23663
2 75860 1 23663
2 75861 1 23665
2 75862 1 23665
2 75863 1 23673
2 75864 1 23673
2 75865 1 23673
2 75866 1 23673
2 75867 1 23688
2 75868 1 23688
2 75869 1 23688
2 75870 1 23691
2 75871 1 23691
2 75872 1 23694
2 75873 1 23694
2 75874 1 23694
2 75875 1 23694
2 75876 1 23695
2 75877 1 23695
2 75878 1 23697
2 75879 1 23697
2 75880 1 23697
2 75881 1 23697
2 75882 1 23697
2 75883 1 23714
2 75884 1 23714
2 75885 1 23715
2 75886 1 23715
2 75887 1 23715
2 75888 1 23715
2 75889 1 23718
2 75890 1 23718
2 75891 1 23719
2 75892 1 23719
2 75893 1 23720
2 75894 1 23720
2 75895 1 23727
2 75896 1 23727
2 75897 1 23727
2 75898 1 23727
2 75899 1 23727
2 75900 1 23727
2 75901 1 23727
2 75902 1 23727
2 75903 1 23727
2 75904 1 23727
2 75905 1 23727
2 75906 1 23727
2 75907 1 23727
2 75908 1 23727
2 75909 1 23727
2 75910 1 23728
2 75911 1 23728
2 75912 1 23728
2 75913 1 23733
2 75914 1 23733
2 75915 1 23733
2 75916 1 23736
2 75917 1 23736
2 75918 1 23751
2 75919 1 23751
2 75920 1 23751
2 75921 1 23753
2 75922 1 23753
2 75923 1 23753
2 75924 1 23753
2 75925 1 23754
2 75926 1 23754
2 75927 1 23754
2 75928 1 23756
2 75929 1 23756
2 75930 1 23757
2 75931 1 23757
2 75932 1 23757
2 75933 1 23758
2 75934 1 23758
2 75935 1 23765
2 75936 1 23765
2 75937 1 23768
2 75938 1 23768
2 75939 1 23768
2 75940 1 23768
2 75941 1 23768
2 75942 1 23768
2 75943 1 23768
2 75944 1 23768
2 75945 1 23768
2 75946 1 23769
2 75947 1 23769
2 75948 1 23769
2 75949 1 23769
2 75950 1 23770
2 75951 1 23770
2 75952 1 23771
2 75953 1 23771
2 75954 1 23771
2 75955 1 23778
2 75956 1 23778
2 75957 1 23779
2 75958 1 23779
2 75959 1 23781
2 75960 1 23781
2 75961 1 23781
2 75962 1 23781
2 75963 1 23781
2 75964 1 23781
2 75965 1 23781
2 75966 1 23781
2 75967 1 23781
2 75968 1 23781
2 75969 1 23785
2 75970 1 23785
2 75971 1 23785
2 75972 1 23785
2 75973 1 23786
2 75974 1 23786
2 75975 1 23798
2 75976 1 23798
2 75977 1 23799
2 75978 1 23799
2 75979 1 23800
2 75980 1 23800
2 75981 1 23800
2 75982 1 23807
2 75983 1 23807
2 75984 1 23807
2 75985 1 23808
2 75986 1 23808
2 75987 1 23819
2 75988 1 23819
2 75989 1 23819
2 75990 1 23822
2 75991 1 23822
2 75992 1 23822
2 75993 1 23823
2 75994 1 23823
2 75995 1 23824
2 75996 1 23824
2 75997 1 23824
2 75998 1 23837
2 75999 1 23837
2 76000 1 23837
2 76001 1 23837
2 76002 1 23837
2 76003 1 23838
2 76004 1 23838
2 76005 1 23838
2 76006 1 23838
2 76007 1 23838
2 76008 1 23838
2 76009 1 23838
2 76010 1 23838
2 76011 1 23858
2 76012 1 23858
2 76013 1 23858
2 76014 1 23861
2 76015 1 23861
2 76016 1 23861
2 76017 1 23880
2 76018 1 23880
2 76019 1 23881
2 76020 1 23881
2 76021 1 23892
2 76022 1 23892
2 76023 1 23892
2 76024 1 23897
2 76025 1 23897
2 76026 1 23903
2 76027 1 23903
2 76028 1 23920
2 76029 1 23920
2 76030 1 23920
2 76031 1 23921
2 76032 1 23921
2 76033 1 23922
2 76034 1 23922
2 76035 1 23923
2 76036 1 23923
2 76037 1 23938
2 76038 1 23938
2 76039 1 23948
2 76040 1 23948
2 76041 1 23949
2 76042 1 23949
2 76043 1 23954
2 76044 1 23954
2 76045 1 23973
2 76046 1 23973
2 76047 1 23975
2 76048 1 23975
2 76049 1 23975
2 76050 1 23975
2 76051 1 23976
2 76052 1 23976
2 76053 1 23976
2 76054 1 23976
2 76055 1 23976
2 76056 1 23976
2 76057 1 23978
2 76058 1 23978
2 76059 1 23990
2 76060 1 23990
2 76061 1 23990
2 76062 1 23991
2 76063 1 23991
2 76064 1 23992
2 76065 1 23992
2 76066 1 23993
2 76067 1 23993
2 76068 1 23993
2 76069 1 23996
2 76070 1 23996
2 76071 1 24004
2 76072 1 24004
2 76073 1 24004
2 76074 1 24007
2 76075 1 24007
2 76076 1 24019
2 76077 1 24019
2 76078 1 24019
2 76079 1 24026
2 76080 1 24026
2 76081 1 24026
2 76082 1 24026
2 76083 1 24029
2 76084 1 24029
2 76085 1 24029
2 76086 1 24037
2 76087 1 24037
2 76088 1 24038
2 76089 1 24038
2 76090 1 24039
2 76091 1 24039
2 76092 1 24045
2 76093 1 24045
2 76094 1 24080
2 76095 1 24080
2 76096 1 24080
2 76097 1 24080
2 76098 1 24080
2 76099 1 24080
2 76100 1 24080
2 76101 1 24084
2 76102 1 24084
2 76103 1 24098
2 76104 1 24098
2 76105 1 24102
2 76106 1 24102
2 76107 1 24109
2 76108 1 24109
2 76109 1 24109
2 76110 1 24113
2 76111 1 24113
2 76112 1 24121
2 76113 1 24121
2 76114 1 24121
2 76115 1 24121
2 76116 1 24125
2 76117 1 24125
2 76118 1 24146
2 76119 1 24146
2 76120 1 24152
2 76121 1 24152
2 76122 1 24152
2 76123 1 24156
2 76124 1 24156
2 76125 1 24159
2 76126 1 24159
2 76127 1 24172
2 76128 1 24172
2 76129 1 24174
2 76130 1 24174
2 76131 1 24183
2 76132 1 24183
2 76133 1 24185
2 76134 1 24185
2 76135 1 24185
2 76136 1 24187
2 76137 1 24187
2 76138 1 24187
2 76139 1 24187
2 76140 1 24187
2 76141 1 24189
2 76142 1 24189
2 76143 1 24189
2 76144 1 24199
2 76145 1 24199
2 76146 1 24199
2 76147 1 24200
2 76148 1 24200
2 76149 1 24201
2 76150 1 24201
2 76151 1 24201
2 76152 1 24201
2 76153 1 24208
2 76154 1 24208
2 76155 1 24222
2 76156 1 24222
2 76157 1 24222
2 76158 1 24231
2 76159 1 24231
2 76160 1 24241
2 76161 1 24241
2 76162 1 24241
2 76163 1 24241
2 76164 1 24241
2 76165 1 24241
2 76166 1 24242
2 76167 1 24242
2 76168 1 24243
2 76169 1 24243
2 76170 1 24244
2 76171 1 24244
2 76172 1 24244
2 76173 1 24245
2 76174 1 24245
2 76175 1 24252
2 76176 1 24252
2 76177 1 24252
2 76178 1 24261
2 76179 1 24261
2 76180 1 24271
2 76181 1 24271
2 76182 1 24271
2 76183 1 24271
2 76184 1 24290
2 76185 1 24290
2 76186 1 24291
2 76187 1 24291
2 76188 1 24303
2 76189 1 24303
2 76190 1 24313
2 76191 1 24313
2 76192 1 24321
2 76193 1 24321
2 76194 1 24323
2 76195 1 24323
2 76196 1 24326
2 76197 1 24326
2 76198 1 24326
2 76199 1 24326
2 76200 1 24333
2 76201 1 24333
2 76202 1 24344
2 76203 1 24344
2 76204 1 24344
2 76205 1 24344
2 76206 1 24344
2 76207 1 24344
2 76208 1 24345
2 76209 1 24345
2 76210 1 24345
2 76211 1 24357
2 76212 1 24357
2 76213 1 24357
2 76214 1 24357
2 76215 1 24357
2 76216 1 24357
2 76217 1 24369
2 76218 1 24369
2 76219 1 24369
2 76220 1 24370
2 76221 1 24370
2 76222 1 24378
2 76223 1 24378
2 76224 1 24378
2 76225 1 24378
2 76226 1 24378
2 76227 1 24378
2 76228 1 24378
2 76229 1 24378
2 76230 1 24392
2 76231 1 24392
2 76232 1 24407
2 76233 1 24407
2 76234 1 24416
2 76235 1 24416
2 76236 1 24416
2 76237 1 24416
2 76238 1 24416
2 76239 1 24427
2 76240 1 24427
2 76241 1 24433
2 76242 1 24433
2 76243 1 24434
2 76244 1 24434
2 76245 1 24448
2 76246 1 24448
2 76247 1 24451
2 76248 1 24451
2 76249 1 24460
2 76250 1 24460
2 76251 1 24485
2 76252 1 24485
2 76253 1 24485
2 76254 1 24485
2 76255 1 24486
2 76256 1 24486
2 76257 1 24487
2 76258 1 24487
2 76259 1 24489
2 76260 1 24489
2 76261 1 24490
2 76262 1 24490
2 76263 1 24497
2 76264 1 24497
2 76265 1 24497
2 76266 1 24514
2 76267 1 24514
2 76268 1 24514
2 76269 1 24516
2 76270 1 24516
2 76271 1 24529
2 76272 1 24529
2 76273 1 24529
2 76274 1 24530
2 76275 1 24530
2 76276 1 24553
2 76277 1 24553
2 76278 1 24561
2 76279 1 24561
2 76280 1 24561
2 76281 1 24568
2 76282 1 24568
2 76283 1 24579
2 76284 1 24579
2 76285 1 24581
2 76286 1 24581
2 76287 1 24597
2 76288 1 24597
2 76289 1 24601
2 76290 1 24601
2 76291 1 24601
2 76292 1 24602
2 76293 1 24602
2 76294 1 24602
2 76295 1 24602
2 76296 1 24604
2 76297 1 24604
2 76298 1 24607
2 76299 1 24607
2 76300 1 24614
2 76301 1 24614
2 76302 1 24614
2 76303 1 24622
2 76304 1 24622
2 76305 1 24632
2 76306 1 24632
2 76307 1 24644
2 76308 1 24644
2 76309 1 24662
2 76310 1 24662
2 76311 1 24676
2 76312 1 24676
2 76313 1 24680
2 76314 1 24680
2 76315 1 24695
2 76316 1 24695
2 76317 1 24695
2 76318 1 24695
2 76319 1 24696
2 76320 1 24696
2 76321 1 24703
2 76322 1 24703
2 76323 1 24703
2 76324 1 24703
2 76325 1 24714
2 76326 1 24714
2 76327 1 24714
2 76328 1 24714
2 76329 1 24714
2 76330 1 24714
2 76331 1 24716
2 76332 1 24716
2 76333 1 24718
2 76334 1 24718
2 76335 1 24726
2 76336 1 24726
2 76337 1 24743
2 76338 1 24743
2 76339 1 24744
2 76340 1 24744
2 76341 1 24744
2 76342 1 24744
2 76343 1 24744
2 76344 1 24787
2 76345 1 24787
2 76346 1 24787
2 76347 1 24787
2 76348 1 24787
2 76349 1 24787
2 76350 1 24789
2 76351 1 24789
2 76352 1 24789
2 76353 1 24789
2 76354 1 24801
2 76355 1 24801
2 76356 1 24812
2 76357 1 24812
2 76358 1 24815
2 76359 1 24815
2 76360 1 24823
2 76361 1 24823
2 76362 1 24827
2 76363 1 24827
2 76364 1 24827
2 76365 1 24841
2 76366 1 24841
2 76367 1 24841
2 76368 1 24842
2 76369 1 24842
2 76370 1 24842
2 76371 1 24842
2 76372 1 24844
2 76373 1 24844
2 76374 1 24846
2 76375 1 24846
2 76376 1 24855
2 76377 1 24855
2 76378 1 24856
2 76379 1 24856
2 76380 1 24864
2 76381 1 24864
2 76382 1 24864
2 76383 1 24864
2 76384 1 24873
2 76385 1 24873
2 76386 1 24878
2 76387 1 24878
2 76388 1 24879
2 76389 1 24879
2 76390 1 24879
2 76391 1 24879
2 76392 1 24879
2 76393 1 24879
2 76394 1 24879
2 76395 1 24889
2 76396 1 24889
2 76397 1 24902
2 76398 1 24902
2 76399 1 24910
2 76400 1 24910
2 76401 1 24910
2 76402 1 24910
2 76403 1 24910
2 76404 1 24910
2 76405 1 24940
2 76406 1 24940
2 76407 1 24944
2 76408 1 24944
2 76409 1 24947
2 76410 1 24947
2 76411 1 24954
2 76412 1 24954
2 76413 1 24954
2 76414 1 24958
2 76415 1 24958
2 76416 1 24958
2 76417 1 24958
2 76418 1 24958
2 76419 1 24958
2 76420 1 24959
2 76421 1 24959
2 76422 1 24974
2 76423 1 24974
2 76424 1 24977
2 76425 1 24977
2 76426 1 24977
2 76427 1 24984
2 76428 1 24984
2 76429 1 24984
2 76430 1 24984
2 76431 1 24984
2 76432 1 24985
2 76433 1 24985
2 76434 1 24985
2 76435 1 24985
2 76436 1 25002
2 76437 1 25002
2 76438 1 25006
2 76439 1 25006
2 76440 1 25015
2 76441 1 25015
2 76442 1 25026
2 76443 1 25026
2 76444 1 25026
2 76445 1 25028
2 76446 1 25028
2 76447 1 25028
2 76448 1 25032
2 76449 1 25032
2 76450 1 25032
2 76451 1 25038
2 76452 1 25038
2 76453 1 25038
2 76454 1 25038
2 76455 1 25039
2 76456 1 25039
2 76457 1 25054
2 76458 1 25054
2 76459 1 25054
2 76460 1 25055
2 76461 1 25055
2 76462 1 25056
2 76463 1 25056
2 76464 1 25057
2 76465 1 25057
2 76466 1 25061
2 76467 1 25061
2 76468 1 25061
2 76469 1 25074
2 76470 1 25074
2 76471 1 25074
2 76472 1 25083
2 76473 1 25083
2 76474 1 25083
2 76475 1 25099
2 76476 1 25099
2 76477 1 25109
2 76478 1 25109
2 76479 1 25110
2 76480 1 25110
2 76481 1 25112
2 76482 1 25112
2 76483 1 25122
2 76484 1 25122
2 76485 1 25125
2 76486 1 25125
2 76487 1 25127
2 76488 1 25127
2 76489 1 25128
2 76490 1 25128
2 76491 1 25130
2 76492 1 25130
2 76493 1 25136
2 76494 1 25136
2 76495 1 25137
2 76496 1 25137
2 76497 1 25141
2 76498 1 25141
2 76499 1 25144
2 76500 1 25144
2 76501 1 25161
2 76502 1 25161
2 76503 1 25161
2 76504 1 25161
2 76505 1 25178
2 76506 1 25178
2 76507 1 25185
2 76508 1 25185
2 76509 1 25189
2 76510 1 25189
2 76511 1 25198
2 76512 1 25198
2 76513 1 25198
2 76514 1 25198
2 76515 1 25238
2 76516 1 25238
2 76517 1 25239
2 76518 1 25239
2 76519 1 25257
2 76520 1 25257
2 76521 1 25259
2 76522 1 25259
2 76523 1 25259
2 76524 1 25259
2 76525 1 25261
2 76526 1 25261
2 76527 1 25266
2 76528 1 25266
2 76529 1 25266
2 76530 1 25268
2 76531 1 25268
2 76532 1 25268
2 76533 1 25281
2 76534 1 25281
2 76535 1 25281
2 76536 1 25281
2 76537 1 25282
2 76538 1 25282
2 76539 1 25291
2 76540 1 25291
2 76541 1 25291
2 76542 1 25291
2 76543 1 25303
2 76544 1 25303
2 76545 1 25306
2 76546 1 25306
2 76547 1 25308
2 76548 1 25308
2 76549 1 25309
2 76550 1 25309
2 76551 1 25309
2 76552 1 25314
2 76553 1 25314
2 76554 1 25314
2 76555 1 25314
2 76556 1 25325
2 76557 1 25325
2 76558 1 25327
2 76559 1 25327
2 76560 1 25327
2 76561 1 25327
2 76562 1 25327
2 76563 1 25327
2 76564 1 25327
2 76565 1 25327
2 76566 1 25328
2 76567 1 25328
2 76568 1 25328
2 76569 1 25328
2 76570 1 25328
2 76571 1 25331
2 76572 1 25331
2 76573 1 25337
2 76574 1 25337
2 76575 1 25337
2 76576 1 25337
2 76577 1 25337
2 76578 1 25337
2 76579 1 25345
2 76580 1 25345
2 76581 1 25345
2 76582 1 25352
2 76583 1 25352
2 76584 1 25352
2 76585 1 25352
2 76586 1 25352
2 76587 1 25360
2 76588 1 25360
2 76589 1 25360
2 76590 1 25360
2 76591 1 25364
2 76592 1 25364
2 76593 1 25381
2 76594 1 25381
2 76595 1 25383
2 76596 1 25383
2 76597 1 25388
2 76598 1 25388
2 76599 1 25389
2 76600 1 25389
2 76601 1 25389
2 76602 1 25400
2 76603 1 25400
2 76604 1 25401
2 76605 1 25401
2 76606 1 25423
2 76607 1 25423
2 76608 1 25427
2 76609 1 25427
2 76610 1 25451
2 76611 1 25451
2 76612 1 25458
2 76613 1 25458
2 76614 1 25458
2 76615 1 25458
2 76616 1 25458
2 76617 1 25458
2 76618 1 25458
2 76619 1 25458
2 76620 1 25458
2 76621 1 25458
2 76622 1 25460
2 76623 1 25460
2 76624 1 25469
2 76625 1 25469
2 76626 1 25517
2 76627 1 25517
2 76628 1 25517
2 76629 1 25528
2 76630 1 25528
2 76631 1 25536
2 76632 1 25536
2 76633 1 25543
2 76634 1 25543
2 76635 1 25543
2 76636 1 25546
2 76637 1 25546
2 76638 1 25546
2 76639 1 25550
2 76640 1 25550
2 76641 1 25553
2 76642 1 25553
2 76643 1 25553
2 76644 1 25553
2 76645 1 25553
2 76646 1 25554
2 76647 1 25554
2 76648 1 25554
2 76649 1 25555
2 76650 1 25555
2 76651 1 25555
2 76652 1 25556
2 76653 1 25556
2 76654 1 25570
2 76655 1 25570
2 76656 1 25599
2 76657 1 25599
2 76658 1 25599
2 76659 1 25599
2 76660 1 25599
2 76661 1 25599
2 76662 1 25601
2 76663 1 25601
2 76664 1 25602
2 76665 1 25602
2 76666 1 25602
2 76667 1 25603
2 76668 1 25603
2 76669 1 25603
2 76670 1 25603
2 76671 1 25604
2 76672 1 25604
2 76673 1 25608
2 76674 1 25608
2 76675 1 25608
2 76676 1 25609
2 76677 1 25609
2 76678 1 25609
2 76679 1 25610
2 76680 1 25610
2 76681 1 25615
2 76682 1 25615
2 76683 1 25616
2 76684 1 25616
2 76685 1 25625
2 76686 1 25625
2 76687 1 25625
2 76688 1 25625
2 76689 1 25625
2 76690 1 25626
2 76691 1 25626
2 76692 1 25626
2 76693 1 25633
2 76694 1 25633
2 76695 1 25633
2 76696 1 25633
2 76697 1 25633
2 76698 1 25633
2 76699 1 25634
2 76700 1 25634
2 76701 1 25635
2 76702 1 25635
2 76703 1 25636
2 76704 1 25636
2 76705 1 25636
2 76706 1 25636
2 76707 1 25636
2 76708 1 25636
2 76709 1 25636
2 76710 1 25643
2 76711 1 25643
2 76712 1 25644
2 76713 1 25644
2 76714 1 25644
2 76715 1 25654
2 76716 1 25654
2 76717 1 25657
2 76718 1 25657
2 76719 1 25657
2 76720 1 25657
2 76721 1 25667
2 76722 1 25667
2 76723 1 25670
2 76724 1 25670
2 76725 1 25673
2 76726 1 25673
2 76727 1 25673
2 76728 1 25675
2 76729 1 25675
2 76730 1 25675
2 76731 1 25679
2 76732 1 25679
2 76733 1 25679
2 76734 1 25687
2 76735 1 25687
2 76736 1 25687
2 76737 1 25689
2 76738 1 25689
2 76739 1 25698
2 76740 1 25698
2 76741 1 25698
2 76742 1 25698
2 76743 1 25699
2 76744 1 25699
2 76745 1 25699
2 76746 1 25699
2 76747 1 25700
2 76748 1 25700
2 76749 1 25702
2 76750 1 25702
2 76751 1 25711
2 76752 1 25711
2 76753 1 25711
2 76754 1 25713
2 76755 1 25713
2 76756 1 25716
2 76757 1 25716
2 76758 1 25721
2 76759 1 25721
2 76760 1 25721
2 76761 1 25721
2 76762 1 25725
2 76763 1 25725
2 76764 1 25725
2 76765 1 25725
2 76766 1 25740
2 76767 1 25740
2 76768 1 25743
2 76769 1 25743
2 76770 1 25749
2 76771 1 25749
2 76772 1 25752
2 76773 1 25752
2 76774 1 25753
2 76775 1 25753
2 76776 1 25753
2 76777 1 25753
2 76778 1 25765
2 76779 1 25765
2 76780 1 25765
2 76781 1 25765
2 76782 1 25768
2 76783 1 25768
2 76784 1 25770
2 76785 1 25770
2 76786 1 25770
2 76787 1 25775
2 76788 1 25775
2 76789 1 25781
2 76790 1 25781
2 76791 1 25788
2 76792 1 25788
2 76793 1 25796
2 76794 1 25796
2 76795 1 25797
2 76796 1 25797
2 76797 1 25798
2 76798 1 25798
2 76799 1 25800
2 76800 1 25800
2 76801 1 25800
2 76802 1 25801
2 76803 1 25801
2 76804 1 25802
2 76805 1 25802
2 76806 1 25810
2 76807 1 25810
2 76808 1 25810
2 76809 1 25810
2 76810 1 25825
2 76811 1 25825
2 76812 1 25825
2 76813 1 25857
2 76814 1 25857
2 76815 1 25857
2 76816 1 25857
2 76817 1 25877
2 76818 1 25877
2 76819 1 25877
2 76820 1 25903
2 76821 1 25903
2 76822 1 25911
2 76823 1 25911
2 76824 1 25934
2 76825 1 25934
2 76826 1 25946
2 76827 1 25946
2 76828 1 25950
2 76829 1 25950
2 76830 1 25950
2 76831 1 25951
2 76832 1 25951
2 76833 1 25965
2 76834 1 25965
2 76835 1 25980
2 76836 1 25980
2 76837 1 25982
2 76838 1 25982
2 76839 1 25990
2 76840 1 25990
2 76841 1 25992
2 76842 1 25992
2 76843 1 25994
2 76844 1 25994
2 76845 1 25999
2 76846 1 25999
2 76847 1 25999
2 76848 1 25999
2 76849 1 26006
2 76850 1 26006
2 76851 1 26006
2 76852 1 26006
2 76853 1 26007
2 76854 1 26007
2 76855 1 26007
2 76856 1 26007
2 76857 1 26007
2 76858 1 26007
2 76859 1 26007
2 76860 1 26007
2 76861 1 26015
2 76862 1 26015
2 76863 1 26015
2 76864 1 26015
2 76865 1 26020
2 76866 1 26020
2 76867 1 26023
2 76868 1 26023
2 76869 1 26043
2 76870 1 26043
2 76871 1 26050
2 76872 1 26050
2 76873 1 26051
2 76874 1 26051
2 76875 1 26067
2 76876 1 26067
2 76877 1 26076
2 76878 1 26076
2 76879 1 26077
2 76880 1 26077
2 76881 1 26077
2 76882 1 26102
2 76883 1 26102
2 76884 1 26103
2 76885 1 26103
2 76886 1 26104
2 76887 1 26104
2 76888 1 26105
2 76889 1 26105
2 76890 1 26125
2 76891 1 26125
2 76892 1 26125
2 76893 1 26126
2 76894 1 26126
2 76895 1 26139
2 76896 1 26139
2 76897 1 26139
2 76898 1 26139
2 76899 1 26139
2 76900 1 26151
2 76901 1 26151
2 76902 1 26151
2 76903 1 26151
2 76904 1 26153
2 76905 1 26153
2 76906 1 26154
2 76907 1 26154
2 76908 1 26182
2 76909 1 26182
2 76910 1 26189
2 76911 1 26189
2 76912 1 26189
2 76913 1 26189
2 76914 1 26189
2 76915 1 26189
2 76916 1 26189
2 76917 1 26202
2 76918 1 26202
2 76919 1 26207
2 76920 1 26207
2 76921 1 26232
2 76922 1 26232
2 76923 1 26233
2 76924 1 26233
2 76925 1 26233
2 76926 1 26233
2 76927 1 26268
2 76928 1 26268
2 76929 1 26268
2 76930 1 26268
2 76931 1 26268
2 76932 1 26298
2 76933 1 26298
2 76934 1 26300
2 76935 1 26300
2 76936 1 26301
2 76937 1 26301
2 76938 1 26301
2 76939 1 26306
2 76940 1 26306
2 76941 1 26321
2 76942 1 26321
2 76943 1 26322
2 76944 1 26322
2 76945 1 26333
2 76946 1 26333
2 76947 1 26348
2 76948 1 26348
2 76949 1 26368
2 76950 1 26368
2 76951 1 26368
2 76952 1 26368
2 76953 1 26377
2 76954 1 26377
2 76955 1 26377
2 76956 1 26378
2 76957 1 26378
2 76958 1 26380
2 76959 1 26380
2 76960 1 26380
2 76961 1 26380
2 76962 1 26415
2 76963 1 26415
2 76964 1 26415
2 76965 1 26433
2 76966 1 26433
2 76967 1 26433
2 76968 1 26433
2 76969 1 26433
2 76970 1 26434
2 76971 1 26434
2 76972 1 26438
2 76973 1 26438
2 76974 1 26438
2 76975 1 26439
2 76976 1 26439
2 76977 1 26439
2 76978 1 26449
2 76979 1 26449
2 76980 1 26449
2 76981 1 26500
2 76982 1 26500
2 76983 1 26511
2 76984 1 26511
2 76985 1 26515
2 76986 1 26515
2 76987 1 26558
2 76988 1 26558
2 76989 1 26567
2 76990 1 26567
2 76991 1 26569
2 76992 1 26569
2 76993 1 26588
2 76994 1 26588
2 76995 1 26588
2 76996 1 26588
2 76997 1 26598
2 76998 1 26598
2 76999 1 26620
2 77000 1 26620
2 77001 1 26621
2 77002 1 26621
2 77003 1 26621
2 77004 1 26641
2 77005 1 26641
2 77006 1 26643
2 77007 1 26643
2 77008 1 26643
2 77009 1 26659
2 77010 1 26659
2 77011 1 26689
2 77012 1 26689
2 77013 1 26700
2 77014 1 26700
2 77015 1 26717
2 77016 1 26717
2 77017 1 26722
2 77018 1 26722
2 77019 1 26734
2 77020 1 26734
2 77021 1 26741
2 77022 1 26741
2 77023 1 26746
2 77024 1 26746
2 77025 1 26746
2 77026 1 26753
2 77027 1 26753
2 77028 1 26810
2 77029 1 26810
2 77030 1 26812
2 77031 1 26812
2 77032 1 26817
2 77033 1 26817
2 77034 1 26861
2 77035 1 26861
2 77036 1 26870
2 77037 1 26870
2 77038 1 26870
2 77039 1 26870
2 77040 1 26876
2 77041 1 26876
2 77042 1 26899
2 77043 1 26899
2 77044 1 26900
2 77045 1 26900
2 77046 1 26906
2 77047 1 26906
2 77048 1 26915
2 77049 1 26915
2 77050 1 26917
2 77051 1 26917
2 77052 1 26929
2 77053 1 26929
2 77054 1 26944
2 77055 1 26944
2 77056 1 26963
2 77057 1 26963
2 77058 1 26963
2 77059 1 26965
2 77060 1 26965
2 77061 1 26977
2 77062 1 26977
2 77063 1 26984
2 77064 1 26984
2 77065 1 27002
2 77066 1 27002
2 77067 1 27007
2 77068 1 27007
2 77069 1 27007
2 77070 1 27024
2 77071 1 27024
2 77072 1 27076
2 77073 1 27076
2 77074 1 27078
2 77075 1 27078
2 77076 1 27082
2 77077 1 27082
2 77078 1 27085
2 77079 1 27085
2 77080 1 27085
2 77081 1 27086
2 77082 1 27086
2 77083 1 27088
2 77084 1 27088
2 77085 1 27095
2 77086 1 27095
2 77087 1 27107
2 77088 1 27107
2 77089 1 27112
2 77090 1 27112
2 77091 1 27118
2 77092 1 27118
2 77093 1 27129
2 77094 1 27129
2 77095 1 27130
2 77096 1 27130
2 77097 1 27160
2 77098 1 27160
2 77099 1 27161
2 77100 1 27161
2 77101 1 27231
2 77102 1 27231
2 77103 1 27231
2 77104 1 27232
2 77105 1 27232
2 77106 1 27243
2 77107 1 27243
2 77108 1 27244
2 77109 1 27244
2 77110 1 27244
2 77111 1 27244
2 77112 1 27247
2 77113 1 27247
2 77114 1 27248
2 77115 1 27248
2 77116 1 27260
2 77117 1 27260
2 77118 1 27263
2 77119 1 27263
2 77120 1 27274
2 77121 1 27274
2 77122 1 27275
2 77123 1 27275
2 77124 1 27281
2 77125 1 27281
2 77126 1 27281
2 77127 1 27281
2 77128 1 27281
2 77129 1 27281
2 77130 1 27281
2 77131 1 27281
2 77132 1 27281
2 77133 1 27281
2 77134 1 27304
2 77135 1 27304
2 77136 1 27327
2 77137 1 27327
2 77138 1 27329
2 77139 1 27329
2 77140 1 27332
2 77141 1 27332
2 77142 1 27340
2 77143 1 27340
2 77144 1 27362
2 77145 1 27362
2 77146 1 27388
2 77147 1 27388
2 77148 1 27399
2 77149 1 27399
2 77150 1 27407
2 77151 1 27407
2 77152 1 27414
2 77153 1 27414
2 77154 1 27414
2 77155 1 27433
2 77156 1 27433
2 77157 1 27434
2 77158 1 27434
2 77159 1 27437
2 77160 1 27437
2 77161 1 27460
2 77162 1 27460
2 77163 1 27461
2 77164 1 27461
2 77165 1 27470
2 77166 1 27470
2 77167 1 27470
2 77168 1 27471
2 77169 1 27471
2 77170 1 27471
2 77171 1 27471
2 77172 1 27471
2 77173 1 27475
2 77174 1 27475
2 77175 1 27483
2 77176 1 27483
2 77177 1 27488
2 77178 1 27488
2 77179 1 27502
2 77180 1 27502
2 77181 1 27507
2 77182 1 27507
2 77183 1 27515
2 77184 1 27515
2 77185 1 27520
2 77186 1 27520
2 77187 1 27523
2 77188 1 27523
2 77189 1 27527
2 77190 1 27527
2 77191 1 27546
2 77192 1 27546
2 77193 1 27546
2 77194 1 27551
2 77195 1 27551
2 77196 1 27571
2 77197 1 27571
2 77198 1 27572
2 77199 1 27572
2 77200 1 27573
2 77201 1 27573
2 77202 1 27592
2 77203 1 27592
2 77204 1 27601
2 77205 1 27601
2 77206 1 27605
2 77207 1 27605
2 77208 1 27631
2 77209 1 27631
2 77210 1 27631
2 77211 1 27659
2 77212 1 27659
2 77213 1 27668
2 77214 1 27668
2 77215 1 27671
2 77216 1 27671
2 77217 1 27685
2 77218 1 27685
2 77219 1 27700
2 77220 1 27700
2 77221 1 27710
2 77222 1 27710
2 77223 1 27710
2 77224 1 27710
2 77225 1 27710
2 77226 1 27711
2 77227 1 27711
2 77228 1 27728
2 77229 1 27728
2 77230 1 27729
2 77231 1 27729
2 77232 1 27730
2 77233 1 27730
2 77234 1 27744
2 77235 1 27744
2 77236 1 27744
2 77237 1 27745
2 77238 1 27745
2 77239 1 27745
2 77240 1 27757
2 77241 1 27757
2 77242 1 27770
2 77243 1 27770
2 77244 1 27770
2 77245 1 27773
2 77246 1 27773
2 77247 1 27773
2 77248 1 27773
2 77249 1 27777
2 77250 1 27777
2 77251 1 27777
2 77252 1 27807
2 77253 1 27807
2 77254 1 27823
2 77255 1 27823
2 77256 1 27825
2 77257 1 27825
2 77258 1 27836
2 77259 1 27836
2 77260 1 27836
2 77261 1 27837
2 77262 1 27837
2 77263 1 27837
2 77264 1 27837
2 77265 1 27837
2 77266 1 27839
2 77267 1 27839
2 77268 1 27846
2 77269 1 27846
2 77270 1 27852
2 77271 1 27852
2 77272 1 27862
2 77273 1 27862
2 77274 1 27868
2 77275 1 27868
2 77276 1 27884
2 77277 1 27884
2 77278 1 27884
2 77279 1 27885
2 77280 1 27885
2 77281 1 27885
2 77282 1 27894
2 77283 1 27894
2 77284 1 27911
2 77285 1 27911
2 77286 1 27927
2 77287 1 27927
2 77288 1 27929
2 77289 1 27929
2 77290 1 27943
2 77291 1 27943
2 77292 1 27943
2 77293 1 27943
2 77294 1 27943
2 77295 1 27943
2 77296 1 27946
2 77297 1 27946
2 77298 1 27948
2 77299 1 27948
2 77300 1 27956
2 77301 1 27956
2 77302 1 27962
2 77303 1 27962
2 77304 1 27982
2 77305 1 27982
2 77306 1 27989
2 77307 1 27989
2 77308 1 27989
2 77309 1 27990
2 77310 1 27990
2 77311 1 27993
2 77312 1 27993
2 77313 1 27996
2 77314 1 27996
2 77315 1 27998
2 77316 1 27998
2 77317 1 28011
2 77318 1 28011
2 77319 1 28011
2 77320 1 28014
2 77321 1 28014
2 77322 1 28014
2 77323 1 28014
2 77324 1 28014
2 77325 1 28014
2 77326 1 28015
2 77327 1 28015
2 77328 1 28021
2 77329 1 28021
2 77330 1 28021
2 77331 1 28048
2 77332 1 28048
2 77333 1 28050
2 77334 1 28050
2 77335 1 28050
2 77336 1 28055
2 77337 1 28055
2 77338 1 28086
2 77339 1 28086
2 77340 1 28092
2 77341 1 28092
2 77342 1 28092
2 77343 1 28092
2 77344 1 28102
2 77345 1 28102
2 77346 1 28130
2 77347 1 28130
2 77348 1 28155
2 77349 1 28155
2 77350 1 28168
2 77351 1 28168
2 77352 1 28168
2 77353 1 28168
2 77354 1 28168
2 77355 1 28197
2 77356 1 28197
2 77357 1 28197
2 77358 1 28197
2 77359 1 28200
2 77360 1 28200
2 77361 1 28200
2 77362 1 28201
2 77363 1 28201
2 77364 1 28201
2 77365 1 28201
2 77366 1 28201
2 77367 1 28209
2 77368 1 28209
2 77369 1 28226
2 77370 1 28226
2 77371 1 28236
2 77372 1 28236
2 77373 1 28266
2 77374 1 28266
2 77375 1 28277
2 77376 1 28277
2 77377 1 28277
2 77378 1 28277
2 77379 1 28280
2 77380 1 28280
2 77381 1 28280
2 77382 1 28280
2 77383 1 28280
2 77384 1 28280
2 77385 1 28288
2 77386 1 28288
2 77387 1 28288
2 77388 1 28301
2 77389 1 28301
2 77390 1 28301
2 77391 1 28301
2 77392 1 28301
2 77393 1 28313
2 77394 1 28313
2 77395 1 28319
2 77396 1 28319
2 77397 1 28348
2 77398 1 28348
2 77399 1 28350
2 77400 1 28350
2 77401 1 28368
2 77402 1 28368
2 77403 1 28375
2 77404 1 28375
2 77405 1 28382
2 77406 1 28382
2 77407 1 28382
2 77408 1 28384
2 77409 1 28384
2 77410 1 28389
2 77411 1 28389
2 77412 1 28393
2 77413 1 28393
2 77414 1 28411
2 77415 1 28411
2 77416 1 28432
2 77417 1 28432
2 77418 1 28439
2 77419 1 28439
2 77420 1 28449
2 77421 1 28449
2 77422 1 28451
2 77423 1 28451
2 77424 1 28455
2 77425 1 28455
2 77426 1 28460
2 77427 1 28460
2 77428 1 28476
2 77429 1 28476
2 77430 1 28482
2 77431 1 28482
2 77432 1 28497
2 77433 1 28497
2 77434 1 28498
2 77435 1 28498
2 77436 1 28498
2 77437 1 28512
2 77438 1 28512
2 77439 1 28513
2 77440 1 28513
2 77441 1 28514
2 77442 1 28514
2 77443 1 28519
2 77444 1 28519
2 77445 1 28532
2 77446 1 28532
2 77447 1 28554
2 77448 1 28554
2 77449 1 28558
2 77450 1 28558
2 77451 1 28560
2 77452 1 28560
2 77453 1 28560
2 77454 1 28561
2 77455 1 28561
2 77456 1 28563
2 77457 1 28563
2 77458 1 28563
2 77459 1 28583
2 77460 1 28583
2 77461 1 28585
2 77462 1 28585
2 77463 1 28617
2 77464 1 28617
2 77465 1 28617
2 77466 1 28622
2 77467 1 28622
2 77468 1 28627
2 77469 1 28627
2 77470 1 28630
2 77471 1 28630
2 77472 1 28641
2 77473 1 28641
2 77474 1 28642
2 77475 1 28642
2 77476 1 28648
2 77477 1 28648
2 77478 1 28648
2 77479 1 28665
2 77480 1 28665
2 77481 1 28687
2 77482 1 28687
2 77483 1 28690
2 77484 1 28690
2 77485 1 28690
2 77486 1 28699
2 77487 1 28699
2 77488 1 28718
2 77489 1 28718
2 77490 1 28724
2 77491 1 28724
2 77492 1 28733
2 77493 1 28733
2 77494 1 28734
2 77495 1 28734
2 77496 1 28734
2 77497 1 28734
2 77498 1 28744
2 77499 1 28744
2 77500 1 28764
2 77501 1 28764
2 77502 1 28764
2 77503 1 28776
2 77504 1 28776
2 77505 1 28779
2 77506 1 28779
2 77507 1 28783
2 77508 1 28783
2 77509 1 28783
2 77510 1 28783
2 77511 1 28783
2 77512 1 28785
2 77513 1 28785
2 77514 1 28787
2 77515 1 28787
2 77516 1 28788
2 77517 1 28788
2 77518 1 28789
2 77519 1 28789
2 77520 1 28796
2 77521 1 28796
2 77522 1 28796
2 77523 1 28826
2 77524 1 28826
2 77525 1 28830
2 77526 1 28830
2 77527 1 28838
2 77528 1 28838
2 77529 1 28855
2 77530 1 28855
2 77531 1 28861
2 77532 1 28861
2 77533 1 28861
2 77534 1 28862
2 77535 1 28862
2 77536 1 28863
2 77537 1 28863
2 77538 1 28863
2 77539 1 28863
2 77540 1 28863
2 77541 1 28876
2 77542 1 28876
2 77543 1 28884
2 77544 1 28884
2 77545 1 28896
2 77546 1 28896
2 77547 1 28900
2 77548 1 28900
2 77549 1 28912
2 77550 1 28912
2 77551 1 28914
2 77552 1 28914
2 77553 1 28927
2 77554 1 28927
2 77555 1 28934
2 77556 1 28934
2 77557 1 28946
2 77558 1 28946
2 77559 1 28956
2 77560 1 28956
2 77561 1 28957
2 77562 1 28957
2 77563 1 28960
2 77564 1 28960
2 77565 1 28978
2 77566 1 28978
2 77567 1 28987
2 77568 1 28987
2 77569 1 28988
2 77570 1 28988
2 77571 1 29038
2 77572 1 29038
2 77573 1 29038
2 77574 1 29040
2 77575 1 29040
2 77576 1 29051
2 77577 1 29051
2 77578 1 29085
2 77579 1 29085
2 77580 1 29085
2 77581 1 29166
2 77582 1 29166
2 77583 1 29166
2 77584 1 29208
2 77585 1 29208
2 77586 1 29244
2 77587 1 29244
2 77588 1 29246
2 77589 1 29246
2 77590 1 29265
2 77591 1 29265
2 77592 1 29265
2 77593 1 29265
2 77594 1 29272
2 77595 1 29272
2 77596 1 29296
2 77597 1 29296
2 77598 1 29346
2 77599 1 29346
2 77600 1 29355
2 77601 1 29355
2 77602 1 29368
2 77603 1 29368
2 77604 1 29384
2 77605 1 29384
2 77606 1 29416
2 77607 1 29416
2 77608 1 29418
2 77609 1 29418
2 77610 1 29440
2 77611 1 29440
2 77612 1 29453
2 77613 1 29453
2 77614 1 29526
2 77615 1 29526
2 77616 1 29527
2 77617 1 29527
2 77618 1 29540
2 77619 1 29540
2 77620 1 29600
2 77621 1 29600
2 77622 1 29601
2 77623 1 29601
2 77624 1 29622
2 77625 1 29622
2 77626 1 29622
2 77627 1 29622
2 77628 1 29653
2 77629 1 29653
2 77630 1 29657
2 77631 1 29657
2 77632 1 29662
2 77633 1 29662
2 77634 1 29692
2 77635 1 29692
2 77636 1 29750
2 77637 1 29750
2 77638 1 29750
2 77639 1 29759
2 77640 1 29759
2 77641 1 29778
2 77642 1 29778
2 77643 1 29784
2 77644 1 29784
2 77645 1 29788
2 77646 1 29788
2 77647 1 29833
2 77648 1 29833
2 77649 1 29833
2 77650 1 29834
2 77651 1 29834
2 77652 1 29834
2 77653 1 29881
2 77654 1 29881
2 77655 1 29897
2 77656 1 29897
2 77657 1 29900
2 77658 1 29900
2 77659 1 29948
2 77660 1 29948
2 77661 1 29960
2 77662 1 29960
2 77663 1 29961
2 77664 1 29961
2 77665 1 29965
2 77666 1 29965
2 77667 1 29999
2 77668 1 29999
2 77669 1 30007
2 77670 1 30007
2 77671 1 30033
2 77672 1 30033
2 77673 1 30046
2 77674 1 30046
2 77675 1 30048
2 77676 1 30048
2 77677 1 30100
2 77678 1 30100
2 77679 1 30100
2 77680 1 30100
2 77681 1 30111
2 77682 1 30111
2 77683 1 30111
2 77684 1 30124
2 77685 1 30124
2 77686 1 30145
2 77687 1 30145
2 77688 1 30164
2 77689 1 30164
2 77690 1 30167
2 77691 1 30167
2 77692 1 30167
2 77693 1 30181
2 77694 1 30181
2 77695 1 30191
2 77696 1 30191
2 77697 1 30192
2 77698 1 30192
2 77699 1 30192
2 77700 1 30192
2 77701 1 30206
2 77702 1 30206
2 77703 1 30238
2 77704 1 30238
2 77705 1 30259
2 77706 1 30259
2 77707 1 30263
2 77708 1 30263
2 77709 1 30297
2 77710 1 30297
2 77711 1 30300
2 77712 1 30300
2 77713 1 30342
2 77714 1 30342
2 77715 1 30451
2 77716 1 30451
2 77717 1 30463
2 77718 1 30463
2 77719 1 30464
2 77720 1 30464
2 77721 1 30468
2 77722 1 30468
2 77723 1 30468
2 77724 1 30492
2 77725 1 30492
2 77726 1 30492
2 77727 1 30492
2 77728 1 30535
2 77729 1 30535
2 77730 1 30547
2 77731 1 30547
2 77732 1 30547
2 77733 1 30547
2 77734 1 30547
2 77735 1 30550
2 77736 1 30550
2 77737 1 30550
2 77738 1 30550
2 77739 1 30550
2 77740 1 30550
2 77741 1 30550
2 77742 1 30550
2 77743 1 30551
2 77744 1 30551
2 77745 1 30569
2 77746 1 30569
2 77747 1 30571
2 77748 1 30571
2 77749 1 30592
2 77750 1 30592
2 77751 1 30593
2 77752 1 30593
2 77753 1 30599
2 77754 1 30599
2 77755 1 30602
2 77756 1 30602
2 77757 1 30612
2 77758 1 30612
2 77759 1 30629
2 77760 1 30629
2 77761 1 30675
2 77762 1 30675
2 77763 1 30683
2 77764 1 30683
2 77765 1 30688
2 77766 1 30688
2 77767 1 30700
2 77768 1 30700
2 77769 1 30732
2 77770 1 30732
2 77771 1 30732
2 77772 1 30732
2 77773 1 30732
2 77774 1 30773
2 77775 1 30773
2 77776 1 30791
2 77777 1 30791
2 77778 1 30797
2 77779 1 30797
2 77780 1 30805
2 77781 1 30805
2 77782 1 30805
2 77783 1 30805
2 77784 1 30807
2 77785 1 30807
2 77786 1 30856
2 77787 1 30856
2 77788 1 30856
2 77789 1 30858
2 77790 1 30858
2 77791 1 30860
2 77792 1 30860
2 77793 1 30899
2 77794 1 30899
2 77795 1 30900
2 77796 1 30900
2 77797 1 30916
2 77798 1 30916
2 77799 1 30917
2 77800 1 30917
2 77801 1 30942
2 77802 1 30942
2 77803 1 30952
2 77804 1 30952
2 77805 1 30974
2 77806 1 30974
2 77807 1 30975
2 77808 1 30975
2 77809 1 30987
2 77810 1 30987
2 77811 1 30988
2 77812 1 30988
2 77813 1 30994
2 77814 1 30994
2 77815 1 30997
2 77816 1 30997
2 77817 1 31029
2 77818 1 31029
2 77819 1 31048
2 77820 1 31048
2 77821 1 31097
2 77822 1 31097
2 77823 1 31131
2 77824 1 31131
2 77825 1 31139
2 77826 1 31139
2 77827 1 31213
2 77828 1 31213
2 77829 1 31227
2 77830 1 31227
2 77831 1 31248
2 77832 1 31248
2 77833 1 31265
2 77834 1 31265
2 77835 1 31317
2 77836 1 31317
2 77837 1 31332
2 77838 1 31332
2 77839 1 31380
2 77840 1 31380
2 77841 1 31384
2 77842 1 31384
2 77843 1 31386
2 77844 1 31386
2 77845 1 31393
2 77846 1 31393
2 77847 1 31405
2 77848 1 31405
2 77849 1 31405
2 77850 1 31405
2 77851 1 31406
2 77852 1 31406
2 77853 1 31407
2 77854 1 31407
2 77855 1 31408
2 77856 1 31408
2 77857 1 31429
2 77858 1 31429
2 77859 1 31432
2 77860 1 31432
2 77861 1 31433
2 77862 1 31433
2 77863 1 31442
2 77864 1 31442
2 77865 1 31476
2 77866 1 31476
2 77867 1 31476
2 77868 1 31484
2 77869 1 31484
2 77870 1 31508
2 77871 1 31508
2 77872 1 31510
2 77873 1 31510
2 77874 1 31525
2 77875 1 31525
2 77876 1 31525
2 77877 1 31540
2 77878 1 31540
2 77879 1 31562
2 77880 1 31562
2 77881 1 31661
2 77882 1 31661
2 77883 1 31664
2 77884 1 31664
2 77885 1 31664
2 77886 1 31664
2 77887 1 31666
2 77888 1 31666
2 77889 1 31666
2 77890 1 31714
2 77891 1 31714
2 77892 1 31717
2 77893 1 31717
2 77894 1 31726
2 77895 1 31726
2 77896 1 31780
2 77897 1 31780
2 77898 1 31822
2 77899 1 31822
2 77900 1 31824
2 77901 1 31824
2 77902 1 31845
2 77903 1 31845
2 77904 1 31854
2 77905 1 31854
2 77906 1 31908
2 77907 1 31908
2 77908 1 31909
2 77909 1 31909
2 77910 1 31910
2 77911 1 31910
2 77912 1 31916
2 77913 1 31916
2 77914 1 31929
2 77915 1 31929
2 77916 1 31930
2 77917 1 31930
2 77918 1 31930
2 77919 1 31955
2 77920 1 31955
2 77921 1 31972
2 77922 1 31972
2 77923 1 32010
2 77924 1 32010
2 77925 1 32021
2 77926 1 32021
2 77927 1 32026
2 77928 1 32026
2 77929 1 32026
2 77930 1 32027
2 77931 1 32027
2 77932 1 32066
2 77933 1 32066
2 77934 1 32066
2 77935 1 32075
2 77936 1 32075
2 77937 1 32094
2 77938 1 32094
2 77939 1 32094
2 77940 1 32135
2 77941 1 32135
2 77942 1 32135
2 77943 1 32194
2 77944 1 32194
2 77945 1 32204
2 77946 1 32204
2 77947 1 32353
2 77948 1 32353
2 77949 1 32353
2 77950 1 32353
2 77951 1 32373
2 77952 1 32373
2 77953 1 32380
2 77954 1 32380
2 77955 1 32436
2 77956 1 32436
2 77957 1 32485
2 77958 1 32485
2 77959 1 32485
2 77960 1 32485
2 77961 1 32485
2 77962 1 32499
2 77963 1 32499
2 77964 1 32499
2 77965 1 32506
2 77966 1 32506
2 77967 1 32506
2 77968 1 32506
2 77969 1 32507
2 77970 1 32507
2 77971 1 32517
2 77972 1 32517
2 77973 1 32519
2 77974 1 32519
2 77975 1 32548
2 77976 1 32548
2 77977 1 32548
2 77978 1 32548
2 77979 1 32548
2 77980 1 32548
2 77981 1 32548
2 77982 1 32548
2 77983 1 32549
2 77984 1 32549
2 77985 1 32549
2 77986 1 32550
2 77987 1 32550
2 77988 1 32550
2 77989 1 32559
2 77990 1 32559
2 77991 1 32563
2 77992 1 32563
2 77993 1 32644
2 77994 1 32644
2 77995 1 32645
2 77996 1 32645
2 77997 1 32660
2 77998 1 32660
2 77999 1 32673
2 78000 1 32673
2 78001 1 32680
2 78002 1 32680
2 78003 1 32690
2 78004 1 32690
2 78005 1 32690
2 78006 1 32690
2 78007 1 32701
2 78008 1 32701
2 78009 1 32736
2 78010 1 32736
2 78011 1 32736
2 78012 1 32738
2 78013 1 32738
2 78014 1 32770
2 78015 1 32770
2 78016 1 32775
2 78017 1 32775
2 78018 1 32775
2 78019 1 32775
2 78020 1 32790
2 78021 1 32790
2 78022 1 32790
2 78023 1 32791
2 78024 1 32791
2 78025 1 32791
2 78026 1 32804
2 78027 1 32804
2 78028 1 32817
2 78029 1 32817
2 78030 1 32839
2 78031 1 32839
2 78032 1 32852
2 78033 1 32852
2 78034 1 32852
2 78035 1 32879
2 78036 1 32879
2 78037 1 32879
2 78038 1 32879
2 78039 1 32881
2 78040 1 32881
2 78041 1 32994
2 78042 1 32994
2 78043 1 32995
2 78044 1 32995
2 78045 1 33017
2 78046 1 33017
2 78047 1 33027
2 78048 1 33027
2 78049 1 33088
2 78050 1 33088
2 78051 1 33088
2 78052 1 33089
2 78053 1 33089
2 78054 1 33089
2 78055 1 33113
2 78056 1 33113
2 78057 1 33113
2 78058 1 33132
2 78059 1 33132
2 78060 1 33132
2 78061 1 33133
2 78062 1 33133
2 78063 1 33156
2 78064 1 33156
2 78065 1 33159
2 78066 1 33159
2 78067 1 33160
2 78068 1 33160
2 78069 1 33223
2 78070 1 33223
2 78071 1 33260
2 78072 1 33260
2 78073 1 33306
2 78074 1 33306
2 78075 1 33307
2 78076 1 33307
2 78077 1 33354
2 78078 1 33354
2 78079 1 33409
2 78080 1 33409
2 78081 1 33483
2 78082 1 33483
2 78083 1 33491
2 78084 1 33491
2 78085 1 33491
2 78086 1 33549
2 78087 1 33549
2 78088 1 33558
2 78089 1 33558
2 78090 1 33564
2 78091 1 33564
2 78092 1 33596
2 78093 1 33596
2 78094 1 33597
2 78095 1 33597
2 78096 1 33629
2 78097 1 33629
2 78098 1 33629
2 78099 1 33630
2 78100 1 33630
2 78101 1 33630
2 78102 1 33655
2 78103 1 33655
2 78104 1 33656
2 78105 1 33656
2 78106 1 33656
2 78107 1 33666
2 78108 1 33666
2 78109 1 33714
2 78110 1 33714
2 78111 1 33881
2 78112 1 33881
2 78113 1 33892
2 78114 1 33892
2 78115 1 33897
2 78116 1 33897
2 78117 1 33916
2 78118 1 33916
2 78119 1 33916
2 78120 1 33964
2 78121 1 33964
2 78122 1 33980
2 78123 1 33980
2 78124 1 33991
2 78125 1 33991
2 78126 1 34020
2 78127 1 34020
2 78128 1 34021
2 78129 1 34021
2 78130 1 34033
2 78131 1 34033
2 78132 1 34074
2 78133 1 34074
2 78134 1 34075
2 78135 1 34075
2 78136 1 34075
2 78137 1 34095
2 78138 1 34095
2 78139 1 34103
2 78140 1 34103
2 78141 1 34104
2 78142 1 34104
2 78143 1 34114
2 78144 1 34114
2 78145 1 34114
2 78146 1 34118
2 78147 1 34118
2 78148 1 34118
2 78149 1 34118
2 78150 1 34118
2 78151 1 34127
2 78152 1 34127
2 78153 1 34141
2 78154 1 34141
2 78155 1 34160
2 78156 1 34160
2 78157 1 34208
2 78158 1 34208
2 78159 1 34209
2 78160 1 34209
2 78161 1 34209
2 78162 1 34209
2 78163 1 34217
2 78164 1 34217
2 78165 1 34255
2 78166 1 34255
2 78167 1 34262
2 78168 1 34262
2 78169 1 34319
2 78170 1 34319
2 78171 1 34351
2 78172 1 34351
2 78173 1 34363
2 78174 1 34363
2 78175 1 34364
2 78176 1 34364
2 78177 1 34384
2 78178 1 34384
2 78179 1 34423
2 78180 1 34423
2 78181 1 34426
2 78182 1 34426
2 78183 1 34451
2 78184 1 34451
2 78185 1 34529
2 78186 1 34529
2 78187 1 34538
2 78188 1 34538
2 78189 1 34541
2 78190 1 34541
2 78191 1 34566
2 78192 1 34566
2 78193 1 34566
2 78194 1 34573
2 78195 1 34573
2 78196 1 34698
2 78197 1 34698
2 78198 1 34714
2 78199 1 34714
2 78200 1 34778
2 78201 1 34778
2 78202 1 34872
2 78203 1 34872
2 78204 1 34905
2 78205 1 34905
2 78206 1 34921
2 78207 1 34921
2 78208 1 34922
2 78209 1 34922
2 78210 1 34982
2 78211 1 34982
2 78212 1 35000
2 78213 1 35000
2 78214 1 35017
2 78215 1 35017
2 78216 1 35037
2 78217 1 35037
2 78218 1 35039
2 78219 1 35039
2 78220 1 35059
2 78221 1 35059
2 78222 1 35105
2 78223 1 35105
2 78224 1 35124
2 78225 1 35124
2 78226 1 35125
2 78227 1 35125
2 78228 1 35128
2 78229 1 35128
2 78230 1 35137
2 78231 1 35137
2 78232 1 35141
2 78233 1 35141
2 78234 1 35143
2 78235 1 35143
2 78236 1 35154
2 78237 1 35154
2 78238 1 35159
2 78239 1 35159
2 78240 1 35159
2 78241 1 35160
2 78242 1 35160
2 78243 1 35160
2 78244 1 35160
2 78245 1 35166
2 78246 1 35166
2 78247 1 35208
2 78248 1 35208
2 78249 1 35208
2 78250 1 35209
2 78251 1 35209
2 78252 1 35210
2 78253 1 35210
2 78254 1 35225
2 78255 1 35225
2 78256 1 35226
2 78257 1 35226
2 78258 1 35289
2 78259 1 35289
2 78260 1 35319
2 78261 1 35319
2 78262 1 35319
2 78263 1 35319
2 78264 1 35321
2 78265 1 35321
2 78266 1 35322
2 78267 1 35322
2 78268 1 35341
2 78269 1 35341
2 78270 1 35345
2 78271 1 35345
2 78272 1 35381
2 78273 1 35381
2 78274 1 35446
2 78275 1 35446
2 78276 1 35480
2 78277 1 35480
2 78278 1 35593
2 78279 1 35593
2 78280 1 35603
2 78281 1 35603
2 78282 1 35671
2 78283 1 35671
2 78284 1 35671
2 78285 1 35671
2 78286 1 35675
2 78287 1 35675
2 78288 1 35677
2 78289 1 35677
2 78290 1 35700
2 78291 1 35700
2 78292 1 35700
2 78293 1 35715
2 78294 1 35715
2 78295 1 35722
2 78296 1 35722
2 78297 1 35727
2 78298 1 35727
2 78299 1 35791
2 78300 1 35791
2 78301 1 35791
2 78302 1 35866
2 78303 1 35866
2 78304 1 35882
2 78305 1 35882
2 78306 1 35882
2 78307 1 35883
2 78308 1 35883
2 78309 1 35908
2 78310 1 35908
2 78311 1 35908
2 78312 1 35908
2 78313 1 35917
2 78314 1 35917
2 78315 1 35937
2 78316 1 35937
2 78317 1 35943
2 78318 1 35943
2 78319 1 35943
2 78320 1 35943
2 78321 1 35950
2 78322 1 35950
2 78323 1 35969
2 78324 1 35969
2 78325 1 35970
2 78326 1 35970
2 78327 1 35981
2 78328 1 35981
2 78329 1 35986
2 78330 1 35986
2 78331 1 35988
2 78332 1 35988
2 78333 1 35989
2 78334 1 35989
2 78335 1 35989
2 78336 1 36001
2 78337 1 36001
2 78338 1 36002
2 78339 1 36002
2 78340 1 36004
2 78341 1 36004
2 78342 1 36021
2 78343 1 36021
2 78344 1 36023
2 78345 1 36023
2 78346 1 36053
2 78347 1 36053
2 78348 1 36053
2 78349 1 36053
2 78350 1 36058
2 78351 1 36058
2 78352 1 36059
2 78353 1 36059
2 78354 1 36072
2 78355 1 36072
2 78356 1 36072
2 78357 1 36072
2 78358 1 36072
2 78359 1 36093
2 78360 1 36093
2 78361 1 36143
2 78362 1 36143
2 78363 1 36196
2 78364 1 36196
2 78365 1 36196
2 78366 1 36196
2 78367 1 36196
2 78368 1 36228
2 78369 1 36228
2 78370 1 36279
2 78371 1 36279
2 78372 1 36280
2 78373 1 36280
2 78374 1 36280
2 78375 1 36296
2 78376 1 36296
2 78377 1 36302
2 78378 1 36302
2 78379 1 36307
2 78380 1 36307
2 78381 1 36317
2 78382 1 36317
2 78383 1 36329
2 78384 1 36329
2 78385 1 36376
2 78386 1 36376
2 78387 1 36407
2 78388 1 36407
2 78389 1 36413
2 78390 1 36413
2 78391 1 36414
2 78392 1 36414
2 78393 1 36414
2 78394 1 36424
2 78395 1 36424
2 78396 1 36448
2 78397 1 36448
2 78398 1 36485
2 78399 1 36485
2 78400 1 36485
2 78401 1 36489
2 78402 1 36489
2 78403 1 36584
2 78404 1 36584
2 78405 1 36606
2 78406 1 36606
2 78407 1 36608
2 78408 1 36608
2 78409 1 36612
2 78410 1 36612
2 78411 1 36689
2 78412 1 36689
2 78413 1 36696
2 78414 1 36696
2 78415 1 36732
2 78416 1 36732
2 78417 1 36739
2 78418 1 36739
2 78419 1 36741
2 78420 1 36741
2 78421 1 36777
2 78422 1 36777
2 78423 1 36828
2 78424 1 36828
2 78425 1 36880
2 78426 1 36880
2 78427 1 36887
2 78428 1 36887
2 78429 1 36887
2 78430 1 36887
2 78431 1 36888
2 78432 1 36888
2 78433 1 36888
2 78434 1 36931
2 78435 1 36931
2 78436 1 36937
2 78437 1 36937
2 78438 1 36944
2 78439 1 36944
2 78440 1 36965
2 78441 1 36965
2 78442 1 36966
2 78443 1 36966
2 78444 1 36967
2 78445 1 36967
2 78446 1 36967
2 78447 1 37002
2 78448 1 37002
2 78449 1 37090
2 78450 1 37090
2 78451 1 37102
2 78452 1 37102
2 78453 1 37105
2 78454 1 37105
2 78455 1 37163
2 78456 1 37163
2 78457 1 37180
2 78458 1 37180
2 78459 1 37209
2 78460 1 37209
2 78461 1 37269
2 78462 1 37269
2 78463 1 37318
2 78464 1 37318
2 78465 1 37319
2 78466 1 37319
2 78467 1 37324
2 78468 1 37324
2 78469 1 37356
2 78470 1 37356
2 78471 1 37387
2 78472 1 37387
2 78473 1 37530
2 78474 1 37530
2 78475 1 37581
2 78476 1 37581
2 78477 1 37581
2 78478 1 37597
2 78479 1 37597
2 78480 1 37604
2 78481 1 37604
2 78482 1 37605
2 78483 1 37605
2 78484 1 37607
2 78485 1 37607
2 78486 1 37608
2 78487 1 37608
2 78488 1 37615
2 78489 1 37615
2 78490 1 37615
2 78491 1 37615
2 78492 1 37615
2 78493 1 37615
2 78494 1 37615
2 78495 1 37632
2 78496 1 37632
2 78497 1 37633
2 78498 1 37633
2 78499 1 37633
2 78500 1 37653
2 78501 1 37653
2 78502 1 37666
2 78503 1 37666
2 78504 1 37666
2 78505 1 37666
2 78506 1 37672
2 78507 1 37672
2 78508 1 37683
2 78509 1 37683
2 78510 1 37684
2 78511 1 37684
2 78512 1 37688
2 78513 1 37688
2 78514 1 37688
2 78515 1 37688
2 78516 1 37692
2 78517 1 37692
2 78518 1 37698
2 78519 1 37698
2 78520 1 37706
2 78521 1 37706
2 78522 1 37707
2 78523 1 37707
2 78524 1 37708
2 78525 1 37708
2 78526 1 37709
2 78527 1 37709
2 78528 1 37712
2 78529 1 37712
2 78530 1 37715
2 78531 1 37715
2 78532 1 37740
2 78533 1 37740
2 78534 1 37753
2 78535 1 37753
2 78536 1 37775
2 78537 1 37775
2 78538 1 37778
2 78539 1 37778
2 78540 1 37782
2 78541 1 37782
2 78542 1 37798
2 78543 1 37798
2 78544 1 37798
2 78545 1 37808
2 78546 1 37808
2 78547 1 37809
2 78548 1 37809
2 78549 1 37809
2 78550 1 37839
2 78551 1 37839
2 78552 1 37840
2 78553 1 37840
2 78554 1 37844
2 78555 1 37844
2 78556 1 37844
2 78557 1 37846
2 78558 1 37846
2 78559 1 37846
2 78560 1 37854
2 78561 1 37854
2 78562 1 37854
2 78563 1 37867
2 78564 1 37867
2 78565 1 37912
2 78566 1 37912
2 78567 1 37912
2 78568 1 37914
2 78569 1 37914
2 78570 1 37914
2 78571 1 37918
2 78572 1 37918
2 78573 1 37918
2 78574 1 37918
2 78575 1 37918
2 78576 1 37919
2 78577 1 37919
2 78578 1 37940
2 78579 1 37940
2 78580 1 37940
2 78581 1 37940
2 78582 1 37941
2 78583 1 37941
2 78584 1 37941
2 78585 1 37942
2 78586 1 37942
2 78587 1 37965
2 78588 1 37965
2 78589 1 37967
2 78590 1 37967
2 78591 1 37979
2 78592 1 37979
2 78593 1 37995
2 78594 1 37995
2 78595 1 38009
2 78596 1 38009
2 78597 1 38009
2 78598 1 38009
2 78599 1 38009
2 78600 1 38009
2 78601 1 38009
2 78602 1 38009
2 78603 1 38009
2 78604 1 38009
2 78605 1 38062
2 78606 1 38062
2 78607 1 38075
2 78608 1 38075
2 78609 1 38081
2 78610 1 38081
2 78611 1 38086
2 78612 1 38086
2 78613 1 38096
2 78614 1 38096
2 78615 1 38096
2 78616 1 38098
2 78617 1 38098
2 78618 1 38110
2 78619 1 38110
2 78620 1 38137
2 78621 1 38137
2 78622 1 38156
2 78623 1 38156
2 78624 1 38156
2 78625 1 38158
2 78626 1 38158
2 78627 1 38160
2 78628 1 38160
2 78629 1 38169
2 78630 1 38169
2 78631 1 38221
2 78632 1 38221
2 78633 1 38221
2 78634 1 38268
2 78635 1 38268
2 78636 1 38305
2 78637 1 38305
2 78638 1 38365
2 78639 1 38365
2 78640 1 38382
2 78641 1 38382
2 78642 1 38382
2 78643 1 38382
2 78644 1 38383
2 78645 1 38383
2 78646 1 38385
2 78647 1 38385
2 78648 1 38386
2 78649 1 38386
2 78650 1 38386
2 78651 1 38386
2 78652 1 38399
2 78653 1 38399
2 78654 1 38427
2 78655 1 38427
2 78656 1 38427
2 78657 1 38498
2 78658 1 38498
2 78659 1 38516
2 78660 1 38516
2 78661 1 38531
2 78662 1 38531
2 78663 1 38540
2 78664 1 38540
2 78665 1 38549
2 78666 1 38549
2 78667 1 38549
2 78668 1 38549
2 78669 1 38549
2 78670 1 38549
2 78671 1 38549
2 78672 1 38569
2 78673 1 38569
2 78674 1 38617
2 78675 1 38617
2 78676 1 38620
2 78677 1 38620
2 78678 1 38624
2 78679 1 38624
2 78680 1 38650
2 78681 1 38650
2 78682 1 38670
2 78683 1 38670
2 78684 1 38676
2 78685 1 38676
2 78686 1 38676
2 78687 1 38691
2 78688 1 38691
2 78689 1 38705
2 78690 1 38705
2 78691 1 38712
2 78692 1 38712
2 78693 1 38712
2 78694 1 38712
2 78695 1 38756
2 78696 1 38756
2 78697 1 38767
2 78698 1 38767
2 78699 1 38768
2 78700 1 38768
2 78701 1 38852
2 78702 1 38852
2 78703 1 38866
2 78704 1 38866
2 78705 1 38890
2 78706 1 38890
2 78707 1 38898
2 78708 1 38898
2 78709 1 38898
2 78710 1 38900
2 78711 1 38900
2 78712 1 38900
2 78713 1 38903
2 78714 1 38903
2 78715 1 38974
2 78716 1 38974
2 78717 1 38975
2 78718 1 38975
2 78719 1 38975
2 78720 1 39008
2 78721 1 39008
2 78722 1 39012
2 78723 1 39012
2 78724 1 39086
2 78725 1 39086
2 78726 1 39087
2 78727 1 39087
2 78728 1 39099
2 78729 1 39099
2 78730 1 39108
2 78731 1 39108
2 78732 1 39108
2 78733 1 39108
2 78734 1 39120
2 78735 1 39120
2 78736 1 39132
2 78737 1 39132
2 78738 1 39132
2 78739 1 39132
2 78740 1 39132
2 78741 1 39132
2 78742 1 39132
2 78743 1 39132
2 78744 1 39132
2 78745 1 39133
2 78746 1 39133
2 78747 1 39140
2 78748 1 39140
2 78749 1 39140
2 78750 1 39140
2 78751 1 39140
2 78752 1 39140
2 78753 1 39140
2 78754 1 39141
2 78755 1 39141
2 78756 1 39170
2 78757 1 39170
2 78758 1 39170
2 78759 1 39171
2 78760 1 39171
2 78761 1 39171
2 78762 1 39189
2 78763 1 39189
2 78764 1 39189
2 78765 1 39189
2 78766 1 39231
2 78767 1 39231
2 78768 1 39246
2 78769 1 39246
2 78770 1 39254
2 78771 1 39254
2 78772 1 39257
2 78773 1 39257
2 78774 1 39257
2 78775 1 39257
2 78776 1 39257
2 78777 1 39262
2 78778 1 39262
2 78779 1 39299
2 78780 1 39299
2 78781 1 39357
2 78782 1 39357
2 78783 1 39360
2 78784 1 39360
2 78785 1 39363
2 78786 1 39363
2 78787 1 39406
2 78788 1 39406
2 78789 1 39439
2 78790 1 39439
2 78791 1 39449
2 78792 1 39449
2 78793 1 39506
2 78794 1 39506
2 78795 1 39523
2 78796 1 39523
2 78797 1 39618
2 78798 1 39618
2 78799 1 39621
2 78800 1 39621
2 78801 1 39624
2 78802 1 39624
2 78803 1 39637
2 78804 1 39637
2 78805 1 39640
2 78806 1 39640
2 78807 1 39683
2 78808 1 39683
2 78809 1 39696
2 78810 1 39696
2 78811 1 39750
2 78812 1 39750
2 78813 1 39765
2 78814 1 39765
2 78815 1 39765
2 78816 1 39828
2 78817 1 39828
2 78818 1 39829
2 78819 1 39829
2 78820 1 39847
2 78821 1 39847
2 78822 1 39879
2 78823 1 39879
2 78824 1 39941
2 78825 1 39941
2 78826 1 39941
2 78827 1 39941
2 78828 1 39941
2 78829 1 39941
2 78830 1 39942
2 78831 1 39942
2 78832 1 39943
2 78833 1 39943
2 78834 1 39943
2 78835 1 39948
2 78836 1 39948
2 78837 1 39976
2 78838 1 39976
2 78839 1 39983
2 78840 1 39983
2 78841 1 39991
2 78842 1 39991
2 78843 1 40001
2 78844 1 40001
2 78845 1 40008
2 78846 1 40008
2 78847 1 40011
2 78848 1 40011
2 78849 1 40025
2 78850 1 40025
2 78851 1 40067
2 78852 1 40067
2 78853 1 40067
2 78854 1 40103
2 78855 1 40103
2 78856 1 40103
2 78857 1 40103
2 78858 1 40107
2 78859 1 40107
2 78860 1 40107
2 78861 1 40180
2 78862 1 40180
2 78863 1 40180
2 78864 1 40180
2 78865 1 40193
2 78866 1 40193
2 78867 1 40193
2 78868 1 40193
2 78869 1 40193
2 78870 1 40193
2 78871 1 40193
2 78872 1 40193
2 78873 1 40263
2 78874 1 40263
2 78875 1 40263
2 78876 1 40263
2 78877 1 40263
2 78878 1 40263
2 78879 1 40263
2 78880 1 40264
2 78881 1 40264
2 78882 1 40267
2 78883 1 40267
2 78884 1 40278
2 78885 1 40278
2 78886 1 40278
2 78887 1 40328
2 78888 1 40328
2 78889 1 40344
2 78890 1 40344
2 78891 1 40433
2 78892 1 40433
2 78893 1 40470
2 78894 1 40470
2 78895 1 40482
2 78896 1 40482
2 78897 1 40482
2 78898 1 40482
2 78899 1 40482
2 78900 1 40482
2 78901 1 40482
2 78902 1 40482
2 78903 1 40484
2 78904 1 40484
2 78905 1 40488
2 78906 1 40488
2 78907 1 40488
2 78908 1 40492
2 78909 1 40492
2 78910 1 40492
2 78911 1 40492
2 78912 1 40492
2 78913 1 40494
2 78914 1 40494
2 78915 1 40494
2 78916 1 40499
2 78917 1 40499
2 78918 1 40507
2 78919 1 40507
2 78920 1 40508
2 78921 1 40508
2 78922 1 40508
2 78923 1 40510
2 78924 1 40510
2 78925 1 40511
2 78926 1 40511
2 78927 1 40512
2 78928 1 40512
2 78929 1 40516
2 78930 1 40516
2 78931 1 40527
2 78932 1 40527
2 78933 1 40539
2 78934 1 40539
2 78935 1 40546
2 78936 1 40546
2 78937 1 40546
2 78938 1 40546
2 78939 1 40547
2 78940 1 40547
2 78941 1 40613
2 78942 1 40613
2 78943 1 40614
2 78944 1 40614
2 78945 1 40614
2 78946 1 40727
2 78947 1 40727
2 78948 1 40727
2 78949 1 40727
2 78950 1 40746
2 78951 1 40746
2 78952 1 40746
2 78953 1 40746
2 78954 1 40746
2 78955 1 40763
2 78956 1 40763
2 78957 1 40771
2 78958 1 40771
2 78959 1 40810
2 78960 1 40810
2 78961 1 40815
2 78962 1 40815
2 78963 1 40829
2 78964 1 40829
2 78965 1 40829
2 78966 1 40829
2 78967 1 40850
2 78968 1 40850
2 78969 1 40850
2 78970 1 40850
2 78971 1 40850
2 78972 1 40851
2 78973 1 40851
2 78974 1 40851
2 78975 1 40863
2 78976 1 40863
2 78977 1 40875
2 78978 1 40875
2 78979 1 40875
2 78980 1 40889
2 78981 1 40889
2 78982 1 40890
2 78983 1 40890
2 78984 1 40891
2 78985 1 40891
2 78986 1 40891
2 78987 1 40894
2 78988 1 40894
2 78989 1 40894
2 78990 1 40894
2 78991 1 40895
2 78992 1 40895
2 78993 1 40895
2 78994 1 40897
2 78995 1 40897
2 78996 1 40897
2 78997 1 40916
2 78998 1 40916
2 78999 1 40924
2 79000 1 40924
2 79001 1 40926
2 79002 1 40926
2 79003 1 40939
2 79004 1 40939
2 79005 1 40939
2 79006 1 40956
2 79007 1 40956
2 79008 1 40959
2 79009 1 40959
2 79010 1 40968
2 79011 1 40968
2 79012 1 40969
2 79013 1 40969
2 79014 1 40969
2 79015 1 40972
2 79016 1 40972
2 79017 1 40976
2 79018 1 40976
2 79019 1 40988
2 79020 1 40988
2 79021 1 40996
2 79022 1 40996
2 79023 1 41002
2 79024 1 41002
2 79025 1 41009
2 79026 1 41009
2 79027 1 41009
2 79028 1 41016
2 79029 1 41016
2 79030 1 41016
2 79031 1 41016
2 79032 1 41016
2 79033 1 41018
2 79034 1 41018
2 79035 1 41040
2 79036 1 41040
2 79037 1 41048
2 79038 1 41048
2 79039 1 41049
2 79040 1 41049
2 79041 1 41053
2 79042 1 41053
2 79043 1 41067
2 79044 1 41067
2 79045 1 41067
2 79046 1 41121
2 79047 1 41121
2 79048 1 41122
2 79049 1 41122
2 79050 1 41122
2 79051 1 41125
2 79052 1 41125
2 79053 1 41139
2 79054 1 41139
2 79055 1 41164
2 79056 1 41164
2 79057 1 41170
2 79058 1 41170
2 79059 1 41184
2 79060 1 41184
2 79061 1 41198
2 79062 1 41198
2 79063 1 41199
2 79064 1 41199
2 79065 1 41201
2 79066 1 41201
2 79067 1 41202
2 79068 1 41202
2 79069 1 41235
2 79070 1 41235
2 79071 1 41240
2 79072 1 41240
2 79073 1 41241
2 79074 1 41241
2 79075 1 41248
2 79076 1 41248
2 79077 1 41253
2 79078 1 41253
2 79079 1 41255
2 79080 1 41255
2 79081 1 41255
2 79082 1 41283
2 79083 1 41283
2 79084 1 41283
2 79085 1 41283
2 79086 1 41283
2 79087 1 41284
2 79088 1 41284
2 79089 1 41284
2 79090 1 41294
2 79091 1 41294
2 79092 1 41297
2 79093 1 41297
2 79094 1 41297
2 79095 1 41297
2 79096 1 41297
2 79097 1 41297
2 79098 1 41297
2 79099 1 41297
2 79100 1 41297
2 79101 1 41311
2 79102 1 41311
2 79103 1 41319
2 79104 1 41319
2 79105 1 41321
2 79106 1 41321
2 79107 1 41321
2 79108 1 41343
2 79109 1 41343
2 79110 1 41344
2 79111 1 41344
2 79112 1 41347
2 79113 1 41347
2 79114 1 41348
2 79115 1 41348
2 79116 1 41349
2 79117 1 41349
2 79118 1 41349
2 79119 1 41356
2 79120 1 41356
2 79121 1 41369
2 79122 1 41369
2 79123 1 41369
2 79124 1 41384
2 79125 1 41384
2 79126 1 41391
2 79127 1 41391
2 79128 1 41404
2 79129 1 41404
2 79130 1 41416
2 79131 1 41416
2 79132 1 41425
2 79133 1 41425
2 79134 1 41435
2 79135 1 41435
2 79136 1 41446
2 79137 1 41446
2 79138 1 41452
2 79139 1 41452
2 79140 1 41455
2 79141 1 41455
2 79142 1 41455
2 79143 1 41467
2 79144 1 41467
2 79145 1 41475
2 79146 1 41475
2 79147 1 41502
2 79148 1 41502
2 79149 1 41506
2 79150 1 41506
2 79151 1 41506
2 79152 1 41510
2 79153 1 41510
2 79154 1 41511
2 79155 1 41511
2 79156 1 41544
2 79157 1 41544
2 79158 1 41570
2 79159 1 41570
2 79160 1 41573
2 79161 1 41573
2 79162 1 41593
2 79163 1 41593
2 79164 1 41596
2 79165 1 41596
2 79166 1 41603
2 79167 1 41603
2 79168 1 41603
2 79169 1 41604
2 79170 1 41604
2 79171 1 41617
2 79172 1 41617
2 79173 1 41617
2 79174 1 41620
2 79175 1 41620
2 79176 1 41629
2 79177 1 41629
2 79178 1 41632
2 79179 1 41632
2 79180 1 41681
2 79181 1 41681
2 79182 1 41681
2 79183 1 41688
2 79184 1 41688
2 79185 1 41696
2 79186 1 41696
2 79187 1 41736
2 79188 1 41736
2 79189 1 41749
2 79190 1 41749
2 79191 1 41769
2 79192 1 41769
2 79193 1 41829
2 79194 1 41829
2 79195 1 41878
2 79196 1 41878
2 79197 1 41899
2 79198 1 41899
2 79199 1 41916
2 79200 1 41916
2 79201 1 41918
2 79202 1 41918
2 79203 1 41918
2 79204 1 42001
2 79205 1 42001
2 79206 1 42050
2 79207 1 42050
2 79208 1 42146
2 79209 1 42146
2 79210 1 42174
2 79211 1 42174
2 79212 1 42183
2 79213 1 42183
2 79214 1 42193
2 79215 1 42193
2 79216 1 42193
2 79217 1 42237
2 79218 1 42237
2 79219 1 42238
2 79220 1 42238
2 79221 1 42239
2 79222 1 42239
2 79223 1 42250
2 79224 1 42250
2 79225 1 42250
2 79226 1 42250
2 79227 1 42250
2 79228 1 42250
2 79229 1 42274
2 79230 1 42274
2 79231 1 42342
2 79232 1 42342
2 79233 1 42343
2 79234 1 42343
2 79235 1 42347
2 79236 1 42347
2 79237 1 42350
2 79238 1 42350
2 79239 1 42351
2 79240 1 42351
2 79241 1 42357
2 79242 1 42357
2 79243 1 42357
2 79244 1 42358
2 79245 1 42358
2 79246 1 42360
2 79247 1 42360
2 79248 1 42360
2 79249 1 42361
2 79250 1 42361
2 79251 1 42369
2 79252 1 42369
2 79253 1 42369
2 79254 1 42370
2 79255 1 42370
2 79256 1 42376
2 79257 1 42376
2 79258 1 42399
2 79259 1 42399
2 79260 1 42409
2 79261 1 42409
2 79262 1 42422
2 79263 1 42422
2 79264 1 42428
2 79265 1 42428
2 79266 1 42429
2 79267 1 42429
2 79268 1 42451
2 79269 1 42451
2 79270 1 42454
2 79271 1 42454
2 79272 1 42559
2 79273 1 42559
2 79274 1 42559
2 79275 1 42559
2 79276 1 42559
2 79277 1 42606
2 79278 1 42606
2 79279 1 42606
2 79280 1 42694
2 79281 1 42694
2 79282 1 42695
2 79283 1 42695
2 79284 1 42715
2 79285 1 42715
2 79286 1 42730
2 79287 1 42730
2 79288 1 42734
2 79289 1 42734
2 79290 1 42741
2 79291 1 42741
2 79292 1 42745
2 79293 1 42745
2 79294 1 42758
2 79295 1 42758
2 79296 1 42766
2 79297 1 42766
2 79298 1 42767
2 79299 1 42767
2 79300 1 42767
2 79301 1 42795
2 79302 1 42795
2 79303 1 42795
2 79304 1 42798
2 79305 1 42798
2 79306 1 42799
2 79307 1 42799
2 79308 1 42815
2 79309 1 42815
2 79310 1 42815
2 79311 1 42816
2 79312 1 42816
2 79313 1 42819
2 79314 1 42819
2 79315 1 42826
2 79316 1 42826
2 79317 1 42826
2 79318 1 42826
2 79319 1 42826
2 79320 1 42830
2 79321 1 42830
2 79322 1 42838
2 79323 1 42838
2 79324 1 42849
2 79325 1 42849
2 79326 1 42850
2 79327 1 42850
2 79328 1 42890
2 79329 1 42890
2 79330 1 42911
2 79331 1 42911
2 79332 1 42919
2 79333 1 42919
2 79334 1 42920
2 79335 1 42920
2 79336 1 42930
2 79337 1 42930
2 79338 1 42946
2 79339 1 42946
2 79340 1 42971
2 79341 1 42971
2 79342 1 42977
2 79343 1 42977
2 79344 1 42999
2 79345 1 42999
2 79346 1 43004
2 79347 1 43004
2 79348 1 43011
2 79349 1 43011
2 79350 1 43013
2 79351 1 43013
2 79352 1 43020
2 79353 1 43020
2 79354 1 43028
2 79355 1 43028
2 79356 1 43028
2 79357 1 43029
2 79358 1 43029
2 79359 1 43035
2 79360 1 43035
2 79361 1 43042
2 79362 1 43042
2 79363 1 43053
2 79364 1 43053
2 79365 1 43060
2 79366 1 43060
2 79367 1 43063
2 79368 1 43063
2 79369 1 43073
2 79370 1 43073
2 79371 1 43099
2 79372 1 43099
2 79373 1 43107
2 79374 1 43107
2 79375 1 43107
2 79376 1 43137
2 79377 1 43137
2 79378 1 43146
2 79379 1 43146
2 79380 1 43146
2 79381 1 43146
2 79382 1 43207
2 79383 1 43207
2 79384 1 43207
2 79385 1 43207
2 79386 1 43207
2 79387 1 43207
2 79388 1 43207
2 79389 1 43207
2 79390 1 43207
2 79391 1 43207
2 79392 1 43207
2 79393 1 43209
2 79394 1 43209
2 79395 1 43217
2 79396 1 43217
2 79397 1 43239
2 79398 1 43239
2 79399 1 43239
2 79400 1 43248
2 79401 1 43248
2 79402 1 43248
2 79403 1 43248
2 79404 1 43250
2 79405 1 43250
2 79406 1 43277
2 79407 1 43277
2 79408 1 43283
2 79409 1 43283
2 79410 1 43302
2 79411 1 43302
2 79412 1 43302
2 79413 1 43302
2 79414 1 43308
2 79415 1 43308
2 79416 1 43313
2 79417 1 43313
2 79418 1 43313
2 79419 1 43321
2 79420 1 43321
2 79421 1 43323
2 79422 1 43323
2 79423 1 43324
2 79424 1 43324
2 79425 1 43325
2 79426 1 43325
2 79427 1 43325
2 79428 1 43326
2 79429 1 43326
2 79430 1 43339
2 79431 1 43339
2 79432 1 43367
2 79433 1 43367
2 79434 1 43405
2 79435 1 43405
2 79436 1 43430
2 79437 1 43430
2 79438 1 43451
2 79439 1 43451
2 79440 1 43451
2 79441 1 43464
2 79442 1 43464
2 79443 1 43478
2 79444 1 43478
2 79445 1 43493
2 79446 1 43493
2 79447 1 43493
2 79448 1 43496
2 79449 1 43496
2 79450 1 43496
2 79451 1 43498
2 79452 1 43498
2 79453 1 43524
2 79454 1 43524
2 79455 1 43532
2 79456 1 43532
2 79457 1 43536
2 79458 1 43536
2 79459 1 43540
2 79460 1 43540
2 79461 1 43551
2 79462 1 43551
2 79463 1 43573
2 79464 1 43573
2 79465 1 43574
2 79466 1 43574
2 79467 1 43577
2 79468 1 43577
2 79469 1 43582
2 79470 1 43582
2 79471 1 43582
2 79472 1 43583
2 79473 1 43583
2 79474 1 43584
2 79475 1 43584
2 79476 1 43599
2 79477 1 43599
2 79478 1 43599
2 79479 1 43599
2 79480 1 43602
2 79481 1 43602
2 79482 1 43607
2 79483 1 43607
2 79484 1 43611
2 79485 1 43611
2 79486 1 43611
2 79487 1 43613
2 79488 1 43613
2 79489 1 43617
2 79490 1 43617
2 79491 1 43628
2 79492 1 43628
2 79493 1 43655
2 79494 1 43655
2 79495 1 43701
2 79496 1 43701
2 79497 1 43708
2 79498 1 43708
2 79499 1 43711
2 79500 1 43711
2 79501 1 43728
2 79502 1 43728
2 79503 1 43758
2 79504 1 43758
2 79505 1 43769
2 79506 1 43769
2 79507 1 43799
2 79508 1 43799
2 79509 1 43803
2 79510 1 43803
2 79511 1 43822
2 79512 1 43822
2 79513 1 43869
2 79514 1 43869
2 79515 1 43878
2 79516 1 43878
2 79517 1 43976
2 79518 1 43976
2 79519 1 43986
2 79520 1 43986
2 79521 1 44007
2 79522 1 44007
2 79523 1 44021
2 79524 1 44021
2 79525 1 44021
2 79526 1 44021
2 79527 1 44053
2 79528 1 44053
2 79529 1 44099
2 79530 1 44099
2 79531 1 44105
2 79532 1 44105
2 79533 1 44114
2 79534 1 44114
2 79535 1 44156
2 79536 1 44156
2 79537 1 44156
2 79538 1 44246
2 79539 1 44246
2 79540 1 44304
2 79541 1 44304
2 79542 1 44331
2 79543 1 44331
2 79544 1 44332
2 79545 1 44332
2 79546 1 44332
2 79547 1 44334
2 79548 1 44334
2 79549 1 44358
2 79550 1 44358
2 79551 1 44358
2 79552 1 44358
2 79553 1 44358
2 79554 1 44378
2 79555 1 44378
2 79556 1 44404
2 79557 1 44404
2 79558 1 44435
2 79559 1 44435
2 79560 1 44438
2 79561 1 44438
2 79562 1 44443
2 79563 1 44443
2 79564 1 44445
2 79565 1 44445
2 79566 1 44445
2 79567 1 44474
2 79568 1 44474
2 79569 1 44474
2 79570 1 44475
2 79571 1 44475
2 79572 1 44549
2 79573 1 44549
2 79574 1 44613
2 79575 1 44613
2 79576 1 44631
2 79577 1 44631
2 79578 1 44719
2 79579 1 44719
2 79580 1 44719
2 79581 1 44739
2 79582 1 44739
2 79583 1 44741
2 79584 1 44741
2 79585 1 44750
2 79586 1 44750
2 79587 1 44750
2 79588 1 44750
2 79589 1 44750
2 79590 1 44770
2 79591 1 44770
2 79592 1 44829
2 79593 1 44829
2 79594 1 44866
2 79595 1 44866
2 79596 1 44866
2 79597 1 44866
2 79598 1 44866
2 79599 1 44866
2 79600 1 44871
2 79601 1 44871
2 79602 1 44872
2 79603 1 44872
2 79604 1 44884
2 79605 1 44884
2 79606 1 44885
2 79607 1 44885
2 79608 1 44951
2 79609 1 44951
2 79610 1 44955
2 79611 1 44955
2 79612 1 44968
2 79613 1 44968
2 79614 1 44973
2 79615 1 44973
2 79616 1 44974
2 79617 1 44974
2 79618 1 44988
2 79619 1 44988
2 79620 1 45007
2 79621 1 45007
2 79622 1 45009
2 79623 1 45009
2 79624 1 45032
2 79625 1 45032
2 79626 1 45033
2 79627 1 45033
2 79628 1 45201
2 79629 1 45201
2 79630 1 45261
2 79631 1 45261
2 79632 1 45274
2 79633 1 45274
2 79634 1 45282
2 79635 1 45282
2 79636 1 45321
2 79637 1 45321
2 79638 1 45325
2 79639 1 45325
2 79640 1 45349
2 79641 1 45349
2 79642 1 45368
2 79643 1 45368
2 79644 1 45373
2 79645 1 45373
2 79646 1 45388
2 79647 1 45388
2 79648 1 45400
2 79649 1 45400
2 79650 1 45404
2 79651 1 45404
2 79652 1 45426
2 79653 1 45426
2 79654 1 45426
2 79655 1 45427
2 79656 1 45427
2 79657 1 45434
2 79658 1 45434
2 79659 1 45464
2 79660 1 45464
2 79661 1 45473
2 79662 1 45473
2 79663 1 45476
2 79664 1 45476
2 79665 1 45522
2 79666 1 45522
2 79667 1 45523
2 79668 1 45523
2 79669 1 45546
2 79670 1 45546
2 79671 1 45586
2 79672 1 45586
2 79673 1 45592
2 79674 1 45592
2 79675 1 45635
2 79676 1 45635
2 79677 1 45684
2 79678 1 45684
2 79679 1 45684
2 79680 1 45716
2 79681 1 45716
2 79682 1 45727
2 79683 1 45727
2 79684 1 45728
2 79685 1 45728
2 79686 1 45750
2 79687 1 45750
2 79688 1 45874
2 79689 1 45874
2 79690 1 45880
2 79691 1 45880
2 79692 1 45925
2 79693 1 45925
2 79694 1 45953
2 79695 1 45953
2 79696 1 45953
2 79697 1 45954
2 79698 1 45954
2 79699 1 45957
2 79700 1 45957
2 79701 1 45961
2 79702 1 45961
2 79703 1 45968
2 79704 1 45968
2 79705 1 45987
2 79706 1 45987
2 79707 1 45988
2 79708 1 45988
2 79709 1 45989
2 79710 1 45989
2 79711 1 46023
2 79712 1 46023
2 79713 1 46166
2 79714 1 46166
2 79715 1 46166
2 79716 1 46166
2 79717 1 46166
2 79718 1 46166
2 79719 1 46166
2 79720 1 46207
2 79721 1 46207
2 79722 1 46275
2 79723 1 46275
2 79724 1 46290
2 79725 1 46290
2 79726 1 46290
2 79727 1 46290
2 79728 1 46290
2 79729 1 46291
2 79730 1 46291
2 79731 1 46291
2 79732 1 46293
2 79733 1 46293
2 79734 1 46310
2 79735 1 46310
2 79736 1 46310
2 79737 1 46334
2 79738 1 46334
2 79739 1 46355
2 79740 1 46355
2 79741 1 46355
2 79742 1 46355
2 79743 1 46435
2 79744 1 46435
2 79745 1 46467
2 79746 1 46467
2 79747 1 46468
2 79748 1 46468
2 79749 1 46534
2 79750 1 46534
2 79751 1 46534
2 79752 1 46564
2 79753 1 46564
2 79754 1 46596
2 79755 1 46596
2 79756 1 46597
2 79757 1 46597
2 79758 1 46600
2 79759 1 46600
2 79760 1 46611
2 79761 1 46611
2 79762 1 46613
2 79763 1 46613
2 79764 1 46613
2 79765 1 46618
2 79766 1 46618
2 79767 1 46621
2 79768 1 46621
2 79769 1 46621
2 79770 1 46621
2 79771 1 46645
2 79772 1 46645
2 79773 1 46764
2 79774 1 46764
2 79775 1 46900
2 79776 1 46900
2 79777 1 46901
2 79778 1 46901
2 79779 1 46911
2 79780 1 46911
2 79781 1 46911
2 79782 1 46926
2 79783 1 46926
2 79784 1 46935
2 79785 1 46935
2 79786 1 46937
2 79787 1 46937
2 79788 1 46937
2 79789 1 46937
2 79790 1 46987
2 79791 1 46987
2 79792 1 46990
2 79793 1 46990
2 79794 1 46990
2 79795 1 47011
2 79796 1 47011
2 79797 1 47192
2 79798 1 47192
2 79799 1 47297
2 79800 1 47297
2 79801 1 47401
2 79802 1 47401
2 79803 1 47401
2 79804 1 47401
2 79805 1 47474
2 79806 1 47474
2 79807 1 47476
2 79808 1 47476
2 79809 1 47532
2 79810 1 47532
2 79811 1 47681
2 79812 1 47681
0 27 5 214 1 25
0 28 5 167 1 48023
0 29 5 148 1 48278
0 30 5 110 1 48453
0 31 5 116 1 48567
0 32 5 155 1 48678
0 33 5 112 1 48836
0 34 5 17 1 48983
0 35 5 42 1 49082
0 36 5 120 1 49139
0 37 5 109 1 49260
0 38 5 117 1 49384
0 39 5 145 1 49506
0 40 5 206 1 49646
0 41 5 156 1 49829
0 42 5 86 1 49991
0 43 5 66 1 50075
0 44 5 200 1 50116
0 45 5 301 1 50320
0 46 5 393 1 50577
0 47 5 349 1 50887
0 48 5 272 1 51196
0 49 5 161 1 51479
0 50 5 67 1 51682
0 51 5 1 1 51829
0 52 7 61 2 52870 50076
0 53 5 116 1 55660
0 54 7 135 2 52212 53032
0 55 5 198 1 55837
0 56 7 99 2 52360 53141
0 57 5 162 1 56170
0 58 7 55 2 52470 53258
0 59 5 115 1 56431
0 60 7 68 2 52045 52912
0 61 5 113 1 56601
0 62 7 2 2 56486 56669
0 63 5 1 1 56782
0 64 7 2 2 56269 56783
0 65 5 2 1 56784
0 66 7 183 2 48454 49385
0 67 5 103 1 56788
0 68 7 4 2 56432 56971
0 69 5 37 1 57074
0 70 7 77 2 48024 49140
0 71 5 78 1 57115
0 72 7 2 2 50321 57192
0 73 5 16 1 57270
0 74 7 3 2 54418 57272
0 75 7 1 2 57078 57288
0 76 5 1 1 75
0 77 7 1 2 56786 76
0 78 5 1 1 77
0 79 7 1 2 26 78
0 80 5 1 1 79
0 81 7 7 2 54117 56487
0 82 7 1 2 56270 57291
0 83 5 4 1 82
0 84 7 1 2 80 57298
0 85 5 1 1 84
0 86 7 1 2 55972 85
0 87 5 1 1 86
0 88 7 6 2 48568 56271
0 89 5 41 1 57302
0 90 7 4 2 49507 56272
0 91 5 5 1 57349
0 92 7 10 2 57308 57353
0 93 5 12 1 57358
0 94 7 170 2 48279 49261
0 95 5 162 1 57380
0 96 7 2 2 57381 57079
0 97 5 2 1 57712
0 98 7 1 2 57359 57714
0 99 5 12 1 98
0 100 7 22 2 47734 54419
0 101 5 10 1 57728
0 102 7 17 2 49141 54118
0 103 5 9 1 57760
0 104 7 2 2 48025 57761
0 105 5 6 1 57786
0 106 7 1 2 57750 57788
0 107 5 1 1 106
0 108 7 1 2 57716 107
0 109 5 1 1 108
0 110 7 6 2 57382 56273
0 111 5 4 1 57794
0 112 7 1 2 57800 57075
0 113 5 5 1 112
0 114 7 30 2 47735 54119
0 115 5 8 1 57809
0 116 7 5 2 54420 57116
0 117 5 3 1 57847
0 118 7 1 2 57810 57848
0 119 7 1 2 57804 118
0 120 5 1 1 119
0 121 7 1 2 109 120
0 122 7 1 2 87 121
0 123 5 1 1 122
0 124 7 1 2 55721 123
0 125 5 1 1 124
0 126 7 114 2 48569 49508
0 127 5 98 1 57855
0 128 7 9 2 52586 57969
0 129 5 53 1 58067
0 130 7 11 2 49142 53851
0 131 5 3 1 58129
0 132 7 9 2 49083 49262
0 133 5 1 1 58143
0 134 7 2 2 58130 58144
0 135 5 4 1 58152
0 136 7 1 2 53142 58154
0 137 5 5 1 136
0 138 7 15 2 48280 54120
0 139 5 7 1 58163
0 140 7 5 2 47736 58164
0 141 5 2 1 58185
0 142 7 1 2 52361 58190
0 143 5 3 1 142
0 144 7 1 2 56488 58192
0 145 5 1 1 144
0 146 7 13 2 48026 54421
0 147 5 10 1 58195
0 148 7 2 2 56489 58196
0 149 5 3 1 58218
0 150 7 10 2 48281 48455
0 151 7 29 2 48027 54121
0 152 5 12 1 58233
0 153 7 6 2 54422 58234
0 154 7 1 2 58223 58274
0 155 5 1 1 154
0 156 7 1 2 58220 155
0 157 7 1 2 145 156
0 158 5 1 1 157
0 159 7 1 2 58158 158
0 160 5 1 1 159
0 161 7 1 2 58068 160
0 162 7 10 2 49084 58131
0 163 5 6 1 58280
0 164 7 3 2 53033 58290
0 165 5 18 1 58296
0 166 7 7 2 52213 50322
0 167 5 7 1 58317
0 168 7 4 2 54423 58324
0 169 5 2 1 58331
0 170 7 5 2 48028 57080
0 171 5 1 1 58337
0 172 7 1 2 58332 58338
0 173 5 1 1 172
0 174 7 2 2 52214 57839
0 175 5 7 1 58342
0 176 7 1 2 58344 57368
0 177 5 1 1 176
0 178 7 1 2 173 177
0 179 5 1 1 178
0 180 7 1 2 58299 179
0 181 5 1 1 180
0 182 7 63 2 49085 53852
0 183 5 56 1 58351
0 184 7 14 2 49143 49263
0 185 5 4 1 58470
0 186 7 7 2 49386 58471
0 187 7 1 2 58352 58488
0 188 5 2 1 187
0 189 7 2 2 53259 58495
0 190 5 2 1 58497
0 191 7 1 2 52471 58498
0 192 5 1 1 191
0 193 7 1 2 52362 58178
0 194 5 2 1 193
0 195 7 7 2 47737 48456
0 196 7 2 2 58165 58503
0 197 5 2 1 58510
0 198 7 1 2 58208 58512
0 199 5 1 1 198
0 200 7 1 2 58501 199
0 201 7 1 2 192 200
0 202 5 1 1 201
0 203 7 1 2 181 202
0 204 7 1 2 161 203
0 205 7 9 2 48457 55973
0 206 5 27 1 58514
0 207 7 8 2 49387 55974
0 208 5 8 1 58550
0 209 7 9 2 58523 58558
0 210 5 11 1 58566
0 211 7 4 2 58575 56670
0 212 5 1 1 58586
0 213 7 1 2 54122 58587
0 214 5 1 1 213
0 215 7 1 2 58496 214
0 216 5 1 1 215
0 217 7 1 2 56490 216
0 218 5 1 1 217
0 219 7 2 2 52913 58414
0 220 5 41 1 58590
0 221 7 1 2 47738 58235
0 222 5 1 1 221
0 223 7 1 2 50578 222
0 224 5 2 1 223
0 225 7 1 2 57717 58633
0 226 5 1 1 225
0 227 7 9 2 48029 56274
0 228 5 5 1 58635
0 229 7 1 2 56491 58636
0 230 5 1 1 229
0 231 7 54 2 54123 54424
0 232 5 21 1 58649
0 233 7 1 2 57081 58650
0 234 5 1 1 233
0 235 7 1 2 230 234
0 236 5 1 1 235
0 237 7 1 2 55975 236
0 238 5 1 1 237
0 239 7 1 2 226 238
0 240 5 1 1 239
0 241 7 1 2 58592 240
0 242 5 1 1 241
0 243 7 1 2 218 242
0 244 7 1 2 204 243
0 245 7 1 2 125 244
0 246 5 1 1 245
0 247 7 1 2 52741 246
0 248 5 1 1 247
0 249 7 11 2 48679 56492
0 250 5 57 1 58724
0 251 7 5 2 50323 58735
0 252 5 1 1 58792
0 253 7 11 2 49647 50579
0 254 5 4 1 58797
0 255 7 12 2 52914 53034
0 256 5 3 1 58812
0 257 7 3 2 50077 58813
0 258 7 16 2 51831 52871
0 259 5 38 1 58830
0 260 7 14 2 52046 52215
0 261 5 1 1 58884
0 262 7 6 2 58831 58885
0 263 7 3 2 58827 58898
0 264 7 1 2 58798 58904
0 265 7 1 2 58793 264
0 266 5 1 1 265
0 267 7 1 2 248 266
0 268 5 1 1 267
0 269 7 1 2 54811 268
0 270 5 1 1 269
0 271 7 4 2 49648 56275
0 272 5 2 1 58907
0 273 7 5 2 54425 56671
0 274 5 3 1 58913
0 275 7 10 2 56972 57801
0 276 5 20 1 58921
0 277 7 1 2 56493 58931
0 278 5 2 1 277
0 279 7 5 2 53403 58069
0 280 5 37 1 58953
0 281 7 1 2 58951 58954
0 282 5 2 1 281
0 283 7 1 2 58914 58995
0 284 5 1 1 283
0 285 7 1 2 58911 284
0 286 5 1 1 285
0 287 7 1 2 52742 286
0 288 5 1 1 287
0 289 7 12 2 52743 49649
0 290 5 7 1 58997
0 291 7 11 2 53404 50580
0 292 5 4 1 59016
0 293 7 9 2 50888 59017
0 294 7 6 2 49388 56494
0 295 7 4 2 48458 59040
0 296 5 6 1 59046
0 297 7 2 2 59050 58070
0 298 5 10 1 59056
0 299 7 1 2 59031 59058
0 300 5 1 1 299
0 301 7 1 2 59009 300
0 302 5 1 1 301
0 303 7 3 2 52915 57550
0 304 5 4 1 59068
0 305 7 8 2 48030 55976
0 306 5 6 1 59075
0 307 7 3 2 57551 59083
0 308 5 3 1 59089
0 309 7 19 2 59071 59092
0 310 5 1 1 59095
0 311 7 1 2 302 59096
0 312 5 1 1 311
0 313 7 5 2 53405 58076
0 314 7 41 2 50581 50889
0 315 5 8 1 59119
0 316 7 3 2 56276 59120
0 317 7 1 2 59114 59168
0 318 5 1 1 317
0 319 7 1 2 312 318
0 320 7 1 2 288 319
0 321 5 1 1 320
0 322 7 1 2 54124 321
0 323 5 1 1 322
0 324 7 6 2 52363 57552
0 325 5 14 1 59171
0 326 7 9 2 53143 59172
0 327 5 39 1 59191
0 328 7 1 2 59200 57117
0 329 5 1 1 328
0 330 7 1 2 58567 329
0 331 5 3 1 330
0 332 7 2 2 58077 59032
0 333 5 1 1 59242
0 334 7 1 2 59010 333
0 335 5 2 1 334
0 336 7 1 2 59239 59244
0 337 5 1 1 336
0 338 7 28 2 57383 57118
0 339 5 2 1 59246
0 340 7 2 2 48459 59247
0 341 7 3 2 49389 59276
0 342 7 3 2 50890 56495
0 343 7 1 2 59018 59281
0 344 7 1 2 59278 343
0 345 5 1 1 344
0 346 7 1 2 337 345
0 347 7 1 2 323 346
0 348 5 1 1 347
0 349 7 1 2 47739 348
0 350 5 1 1 349
0 351 7 1 2 59051 58955
0 352 5 6 1 351
0 353 7 6 2 49144 55977
0 354 5 8 1 59290
0 355 7 6 2 59296 59084
0 356 5 8 1 59304
0 357 7 9 2 52744 54426
0 358 5 1 1 59318
0 359 7 1 2 59310 59319
0 360 7 1 2 59284 359
0 361 5 1 1 360
0 362 7 1 2 350 361
0 363 5 1 1 362
0 364 7 1 2 55722 363
0 365 5 1 1 364
0 366 7 4 2 48031 58472
0 367 5 3 1 59327
0 368 7 6 2 47740 49264
0 369 5 3 1 59334
0 370 7 1 2 58262 59340
0 371 5 1 1 370
0 372 7 1 2 58593 371
0 373 5 1 1 372
0 374 7 1 2 59331 373
0 375 5 2 1 374
0 376 7 1 2 59343 59320
0 377 5 1 1 376
0 378 7 2 2 57119 58145
0 379 7 14 2 53406 50891
0 380 5 2 1 59347
0 381 7 16 2 54125 50582
0 382 5 3 1 59363
0 383 7 2 2 53853 59364
0 384 7 1 2 59348 59382
0 385 7 1 2 59345 384
0 386 5 1 1 385
0 387 7 1 2 377 386
0 388 5 1 1 387
0 389 7 1 2 56789 388
0 390 5 1 1 389
0 391 7 2 2 47741 58594
0 392 5 4 1 59384
0 393 7 1 2 57193 59386
0 394 5 1 1 393
0 395 7 1 2 59321 394
0 396 5 1 1 395
0 397 7 4 2 53854 50583
0 398 7 2 2 50892 59390
0 399 7 4 2 49145 53407
0 400 7 1 2 49086 58236
0 401 7 1 2 59396 400
0 402 7 1 2 59394 401
0 403 5 1 1 402
0 404 7 1 2 396 403
0 405 5 1 1 404
0 406 7 1 2 56790 405
0 407 5 1 1 406
0 408 7 5 2 58353 57762
0 409 5 9 1 59400
0 410 7 2 2 56973 59405
0 411 5 1 1 59414
0 412 7 2 2 54126 58595
0 413 5 4 1 59416
0 414 7 16 2 49087 49146
0 415 5 3 1 59422
0 416 7 6 2 47742 53855
0 417 5 4 1 59441
0 418 7 7 2 59423 59442
0 419 5 7 1 59451
0 420 7 2 2 59418 59458
0 421 5 1 1 59465
0 422 7 1 2 48032 421
0 423 5 2 1 422
0 424 7 1 2 59415 59467
0 425 5 1 1 424
0 426 7 13 2 54427 56277
0 427 5 6 1 59469
0 428 7 1 2 52745 59470
0 429 7 1 2 425 428
0 430 5 1 1 429
0 431 7 1 2 50324 58291
0 432 5 4 1 431
0 433 7 1 2 48033 59488
0 434 5 1 1 433
0 435 7 1 2 59419 434
0 436 5 1 1 435
0 437 7 1 2 56791 59033
0 438 7 1 2 436 437
0 439 5 1 1 438
0 440 7 1 2 430 439
0 441 5 1 1 440
0 442 7 1 2 49265 441
0 443 5 1 1 442
0 444 7 1 2 407 443
0 445 5 1 1 444
0 446 7 1 2 48282 445
0 447 5 1 1 446
0 448 7 1 2 390 447
0 449 5 1 1 448
0 450 7 1 2 56496 449
0 451 5 1 1 450
0 452 7 14 2 53856 54127
0 453 5 4 1 59492
0 454 7 4 2 49088 59493
0 455 5 4 1 59510
0 456 7 1 2 50584 59514
0 457 5 5 1 456
0 458 7 1 2 55978 59518
0 459 5 1 1 458
0 460 7 8 2 49266 53857
0 461 5 1 1 59523
0 462 7 1 2 48283 49089
0 463 7 3 2 59524 462
0 464 5 2 1 59531
0 465 7 1 2 459 59534
0 466 5 1 1 465
0 467 7 1 2 57120 466
0 468 5 1 1 467
0 469 7 1 2 50585 58263
0 470 5 2 1 469
0 471 7 1 2 59201 59536
0 472 5 1 1 471
0 473 7 1 2 468 472
0 474 5 1 1 473
0 475 7 1 2 49650 474
0 476 5 1 1 475
0 477 7 1 2 58197 58078
0 478 7 1 2 59291 477
0 479 5 1 1 478
0 480 7 1 2 476 479
0 481 5 1 1 480
0 482 7 1 2 52746 481
0 483 5 1 1 482
0 484 7 16 2 47743 48034
0 485 5 8 1 59538
0 486 7 1 2 50325 59554
0 487 5 11 1 486
0 488 7 5 2 54428 59562
0 489 7 1 2 59573 59285
0 490 5 1 1 489
0 491 7 1 2 49651 58637
0 492 5 1 1 491
0 493 7 1 2 490 492
0 494 5 1 1 493
0 495 7 1 2 52747 494
0 496 5 1 1 495
0 497 7 1 2 58638 59243
0 498 5 1 1 497
0 499 7 1 2 496 498
0 500 5 1 1 499
0 501 7 1 2 55838 58292
0 502 5 7 1 501
0 503 7 1 2 500 59578
0 504 5 1 1 503
0 505 7 8 2 47744 55979
0 506 5 2 1 59585
0 507 7 1 2 58264 59593
0 508 5 1 1 507
0 509 7 1 2 58958 59322
0 510 7 1 2 508 509
0 511 5 1 1 510
0 512 7 1 2 50326 58568
0 513 5 1 1 512
0 514 7 1 2 59202 59245
0 515 7 1 2 513 514
0 516 5 1 1 515
0 517 7 1 2 511 516
0 518 5 1 1 517
0 519 7 1 2 58596 518
0 520 5 1 1 519
0 521 7 3 2 48035 53408
0 522 7 5 2 54128 59121
0 523 7 1 2 59595 59598
0 524 5 1 1 523
0 525 7 1 2 358 524
0 526 5 1 1 525
0 527 7 1 2 59203 526
0 528 5 1 1 527
0 529 7 24 2 49267 54129
0 530 5 18 1 59603
0 531 7 22 2 53035 50327
0 532 5 23 1 59645
0 533 7 1 2 48284 59667
0 534 5 5 1 533
0 535 7 5 2 59627 59690
0 536 5 6 1 59695
0 537 7 8 2 48036 53858
0 538 5 2 1 59706
0 539 7 10 2 59424 59707
0 540 5 8 1 59716
0 541 7 1 2 59717 59034
0 542 7 1 2 59700 541
0 543 5 1 1 542
0 544 7 1 2 528 543
0 545 5 1 1 544
0 546 7 1 2 58079 545
0 547 5 1 1 546
0 548 7 1 2 520 547
0 549 7 1 2 504 548
0 550 7 1 2 483 549
0 551 7 1 2 451 550
0 552 7 1 2 365 551
0 553 7 1 2 270 552
0 554 5 1 1 553
0 555 7 1 2 53917 554
0 556 5 1 1 555
0 557 7 13 2 53036 50117
0 558 5 9 1 59734
0 559 7 7 2 52216 59735
0 560 5 9 1 59756
0 561 7 11 2 52916 55661
0 562 5 4 1 59772
0 563 7 1 2 55980 59783
0 564 5 4 1 563
0 565 7 5 2 57553 59787
0 566 5 1 1 59791
0 567 7 6 2 51832 57554
0 568 5 9 1 59796
0 569 7 2 2 59802 59072
0 570 7 7 2 52917 50078
0 571 5 2 1 59813
0 572 7 3 2 58832 59814
0 573 5 6 1 59822
0 574 7 1 2 59811 59825
0 575 5 1 1 574
0 576 7 1 2 50118 575
0 577 5 1 1 576
0 578 7 2 2 566 577
0 579 5 1 1 59831
0 580 7 1 2 52047 579
0 581 5 1 1 580
0 582 7 1 2 59763 581
0 583 5 1 1 582
0 584 7 1 2 50893 583
0 585 5 1 1 584
0 586 7 5 2 49147 55723
0 587 5 33 1 59833
0 588 7 20 2 50119 50894
0 589 5 4 1 59871
0 590 7 11 2 51833 50895
0 591 5 4 1 59895
0 592 7 1 2 50586 59757
0 593 5 1 1 592
0 594 7 1 2 59906 593
0 595 5 1 1 594
0 596 7 1 2 52048 595
0 597 5 1 1 596
0 598 7 1 2 59891 597
0 599 5 1 1 598
0 600 7 1 2 50328 599
0 601 5 1 1 600
0 602 7 16 2 50896 57555
0 603 5 1 1 59910
0 604 7 29 2 51834 50120
0 605 5 49 1 59926
0 606 7 4 2 49268 59955
0 607 5 15 1 60004
0 608 7 4 2 48285 59956
0 609 5 6 1 60023
0 610 7 5 2 60008 60027
0 611 5 1 1 60033
0 612 7 1 2 59911 60034
0 613 5 1 1 612
0 614 7 1 2 601 613
0 615 5 1 1 614
0 616 7 1 2 59838 615
0 617 5 2 1 616
0 618 7 2 2 49269 59784
0 619 5 9 1 60040
0 620 7 1 2 51835 60042
0 621 5 1 1 620
0 622 7 1 2 48286 621
0 623 5 1 1 622
0 624 7 11 2 49270 53918
0 625 5 3 1 60051
0 626 7 3 2 49148 59539
0 627 5 1 1 60065
0 628 7 1 2 60052 60066
0 629 5 3 1 628
0 630 7 1 2 623 60068
0 631 5 1 1 630
0 632 7 1 2 53037 57194
0 633 5 12 1 632
0 634 7 6 2 48037 49271
0 635 5 3 1 60083
0 636 7 1 2 50121 60089
0 637 5 2 1 636
0 638 7 1 2 60071 60092
0 639 7 1 2 631 638
0 640 5 1 1 639
0 641 7 7 2 53038 50079
0 642 5 2 1 60094
0 643 7 4 2 52217 60095
0 644 5 2 1 60103
0 645 7 2 2 52918 60104
0 646 7 17 2 51836 52049
0 647 5 9 1 60111
0 648 7 2 2 53919 60128
0 649 5 20 1 60137
0 650 7 3 2 52872 50587
0 651 7 1 2 60139 60159
0 652 7 1 2 60109 651
0 653 5 1 1 652
0 654 7 1 2 54812 653
0 655 5 1 1 654
0 656 7 1 2 50329 655
0 657 7 1 2 640 656
0 658 5 1 1 657
0 659 7 1 2 60038 658
0 660 7 1 2 585 659
0 661 5 1 1 660
0 662 7 1 2 53409 661
0 663 5 1 1 662
0 664 7 1 2 58725 663
0 665 5 1 1 664
0 666 7 7 2 52873 52919
0 667 5 1 1 60162
0 668 7 3 2 50080 60163
0 669 5 1 1 60169
0 670 7 1 2 54130 669
0 671 5 2 1 670
0 672 7 2 2 52050 60172
0 673 5 3 1 60174
0 674 7 50 2 50122 50330
0 675 5 29 1 60179
0 676 7 17 2 52051 50123
0 677 5 43 1 60258
0 678 7 11 2 54131 60275
0 679 5 16 1 60318
0 680 7 8 2 47745 49149
0 681 5 9 1 60345
0 682 7 1 2 60329 60353
0 683 5 3 1 682
0 684 7 2 2 60229 60362
0 685 5 1 1 60365
0 686 7 2 2 60176 60366
0 687 5 1 1 60367
0 688 7 36 2 53920 54132
0 689 5 28 1 60369
0 690 7 2 2 52218 60405
0 691 5 3 1 60433
0 692 7 1 2 53039 60434
0 693 5 6 1 692
0 694 7 1 2 60368 60438
0 695 5 1 1 694
0 696 7 1 2 57556 695
0 697 5 1 1 696
0 698 7 6 2 52052 55839
0 699 5 5 1 60444
0 700 7 1 2 60330 59823
0 701 5 1 1 700
0 702 7 1 2 50331 60259
0 703 5 8 1 702
0 704 7 3 2 701 60455
0 705 5 1 1 60463
0 706 7 1 2 60450 60464
0 707 7 1 2 697 706
0 708 5 1 1 707
0 709 7 1 2 50897 708
0 710 5 1 1 709
0 711 7 18 2 52219 52920
0 712 5 1 1 60466
0 713 7 5 2 53040 60467
0 714 7 6 2 50081 50332
0 715 5 1 1 60489
0 716 7 5 2 52874 60490
0 717 5 2 1 60495
0 718 7 4 2 60484 60496
0 719 5 1 1 60502
0 720 7 1 2 50124 60503
0 721 5 1 1 720
0 722 7 1 2 54813 721
0 723 5 2 1 722
0 724 7 1 2 50588 60506
0 725 5 1 1 724
0 726 7 1 2 49652 725
0 727 7 1 2 60039 726
0 728 7 1 2 710 727
0 729 5 2 1 728
0 730 7 1 2 665 60508
0 731 5 1 1 730
0 732 7 8 2 53144 53260
0 733 7 5 2 52472 60510
0 734 7 41 2 50333 50589
0 735 5 15 1 60523
0 736 7 3 2 54814 60564
0 737 5 4 1 60579
0 738 7 2 2 52364 60582
0 739 5 1 1 60586
0 740 7 1 2 60518 60587
0 741 5 1 1 740
0 742 7 1 2 731 741
0 743 5 1 1 742
0 744 7 1 2 48837 743
0 745 5 1 1 744
0 746 7 3 2 49653 56171
0 747 7 2 2 56433 60588
0 748 7 12 2 51837 52220
0 749 5 3 1 60593
0 750 7 4 2 59736 60594
0 751 5 7 1 60608
0 752 7 7 2 50334 57557
0 753 5 13 1 60619
0 754 7 10 2 51838 55662
0 755 5 11 1 60639
0 756 7 3 2 53921 60649
0 757 5 8 1 60660
0 758 7 1 2 55981 60661
0 759 5 1 1 758
0 760 7 1 2 60620 759
0 761 5 2 1 760
0 762 7 1 2 60612 60671
0 763 5 3 1 762
0 764 7 1 2 57195 60673
0 765 5 1 1 764
0 766 7 12 2 50082 50125
0 767 5 22 1 60676
0 768 7 4 2 52875 60677
0 769 5 6 1 60710
0 770 7 1 2 54133 60714
0 771 5 14 1 770
0 772 7 4 2 51839 60720
0 773 5 2 1 60734
0 774 7 11 2 54134 56672
0 775 5 11 1 60740
0 776 7 2 2 50126 60751
0 777 5 4 1 60762
0 778 7 7 2 52053 52876
0 779 5 2 1 60768
0 780 7 2 2 59815 60769
0 781 5 8 1 60777
0 782 7 2 2 60764 60779
0 783 5 2 1 60787
0 784 7 2 2 60738 60788
0 785 5 1 1 60791
0 786 7 1 2 55840 785
0 787 5 1 1 786
0 788 7 5 2 52054 60180
0 789 5 4 1 60793
0 790 7 5 2 55663 60794
0 791 5 1 1 60802
0 792 7 1 2 52921 60803
0 793 5 6 1 792
0 794 7 2 2 60181 55664
0 795 5 6 1 60813
0 796 7 5 2 51840 56602
0 797 5 1 1 60821
0 798 7 1 2 60822 60721
0 799 5 1 1 798
0 800 7 2 2 60815 799
0 801 5 1 1 60826
0 802 7 1 2 57558 801
0 803 5 1 1 802
0 804 7 1 2 60807 803
0 805 7 3 2 787 804
0 806 5 2 1 60828
0 807 7 1 2 765 60829
0 808 5 1 1 807
0 809 7 1 2 54429 808
0 810 5 1 1 809
0 811 7 9 2 53922 55724
0 812 5 24 1 60833
0 813 7 2 2 52922 60842
0 814 5 2 1 60866
0 815 7 3 2 52055 60843
0 816 5 4 1 60870
0 817 7 3 2 60868 60873
0 818 5 2 1 60877
0 819 7 5 2 49272 56673
0 820 5 3 1 60882
0 821 7 2 2 60024 60883
0 822 5 2 1 60890
0 823 7 1 2 60878 60891
0 824 5 2 1 823
0 825 7 1 2 59365 60894
0 826 5 1 1 825
0 827 7 1 2 810 826
0 828 5 1 1 827
0 829 7 1 2 60591 828
0 830 5 1 1 829
0 831 7 2 2 50590 59628
0 832 5 6 1 60896
0 833 7 35 2 47746 49090
0 834 5 11 1 60904
0 835 7 5 2 57121 60905
0 836 5 2 1 60950
0 837 7 5 2 53859 60951
0 838 5 2 1 60957
0 839 7 1 2 60898 60958
0 840 5 1 1 839
0 841 7 14 2 47747 58354
0 842 5 14 1 60964
0 843 7 2 2 57196 60978
0 844 5 2 1 60992
0 845 7 1 2 50335 60993
0 846 5 1 1 845
0 847 7 1 2 49273 846
0 848 5 1 1 847
0 849 7 8 2 54135 57122
0 850 5 3 1 60996
0 851 7 1 2 59341 59515
0 852 5 1 1 851
0 853 7 1 2 56674 852
0 854 5 1 1 853
0 855 7 1 2 61004 854
0 856 7 1 2 848 855
0 857 5 1 1 856
0 858 7 1 2 54430 857
0 859 5 1 1 858
0 860 7 1 2 840 859
0 861 5 1 1 860
0 862 7 1 2 48287 861
0 863 5 1 1 862
0 864 7 21 2 49274 54431
0 865 5 4 1 61007
0 866 7 1 2 59406 59468
0 867 5 1 1 866
0 868 7 1 2 61008 867
0 869 5 1 1 868
0 870 7 1 2 863 869
0 871 5 1 1 870
0 872 7 1 2 57082 871
0 873 5 1 1 872
0 874 7 2 2 627 60752
0 875 5 2 1 61032
0 876 7 1 2 57369 61034
0 877 5 1 1 876
0 878 7 2 2 57083 57811
0 879 7 1 2 58915 61036
0 880 5 1 1 879
0 881 7 1 2 877 880
0 882 5 1 1 881
0 883 7 1 2 55982 882
0 884 5 1 1 883
0 885 7 1 2 57718 58916
0 886 5 1 1 885
0 887 7 1 2 47748 58996
0 888 5 1 1 887
0 889 7 1 2 886 888
0 890 7 1 2 884 889
0 891 5 1 1 890
0 892 7 1 2 55725 891
0 893 5 1 1 892
0 894 7 1 2 58591 60445
0 895 5 1 1 894
0 896 7 1 2 59286 895
0 897 5 1 1 896
0 898 7 1 2 48288 58300
0 899 5 3 1 898
0 900 7 9 2 51841 52923
0 901 5 9 1 61041
0 902 7 9 2 54136 55983
0 903 5 9 1 61059
0 904 7 2 2 50591 61068
0 905 5 5 1 61077
0 906 7 1 2 61050 61079
0 907 5 1 1 906
0 908 7 13 2 53860 59425
0 909 5 1 1 61084
0 910 7 1 2 53041 57840
0 911 5 8 1 910
0 912 7 1 2 61085 61097
0 913 5 1 1 912
0 914 7 1 2 907 913
0 915 7 1 2 61038 914
0 916 5 1 1 915
0 917 7 1 2 48038 916
0 918 5 1 1 917
0 919 7 7 2 48289 59604
0 920 5 16 1 61105
0 921 7 5 2 50336 55841
0 922 5 13 1 61128
0 923 7 2 2 54432 61133
0 924 5 2 1 61146
0 925 7 2 2 61112 61148
0 926 7 1 2 48290 61098
0 927 5 1 1 926
0 928 7 1 2 47749 60899
0 929 5 1 1 928
0 930 7 1 2 927 929
0 931 5 2 1 930
0 932 7 1 2 58597 61152
0 933 5 2 1 932
0 934 7 1 2 61150 61154
0 935 7 1 2 918 934
0 936 5 1 1 935
0 937 7 1 2 57370 936
0 938 5 1 1 937
0 939 7 1 2 897 938
0 940 7 1 2 893 939
0 941 7 1 2 873 940
0 942 5 1 1 941
0 943 7 1 2 52748 942
0 944 5 1 1 943
0 945 7 1 2 830 944
0 946 5 1 1 945
0 947 7 1 2 54815 946
0 948 5 1 1 947
0 949 7 5 2 47750 56278
0 950 5 4 1 61156
0 951 7 2 2 55984 61157
0 952 5 2 1 61165
0 953 7 1 2 52924 61167
0 954 5 1 1 953
0 955 7 2 2 58355 59563
0 956 5 1 1 61169
0 957 7 2 2 59085 59594
0 958 5 1 1 61171
0 959 7 1 2 56279 958
0 960 5 1 1 959
0 961 7 1 2 956 960
0 962 5 1 1 961
0 963 7 1 2 954 962
0 964 5 1 1 963
0 965 7 1 2 58265 964
0 966 5 1 1 965
0 967 7 1 2 59204 58598
0 968 7 1 2 966 967
0 969 5 1 1 968
0 970 7 4 2 48039 55726
0 971 5 18 1 61173
0 972 7 3 2 59839 61177
0 973 5 2 1 61195
0 974 7 5 2 54137 59205
0 975 5 1 1 61200
0 976 7 1 2 47751 61201
0 977 5 1 1 976
0 978 7 1 2 58569 977
0 979 5 4 1 978
0 980 7 1 2 61198 61205
0 981 5 1 1 980
0 982 7 1 2 56280 59803
0 983 7 1 2 59093 982
0 984 5 1 1 983
0 985 7 1 2 52587 984
0 986 7 1 2 981 985
0 987 7 1 2 969 986
0 988 5 1 1 987
0 989 7 1 2 49654 988
0 990 5 1 1 989
0 991 7 3 2 49655 56497
0 992 5 5 1 61209
0 993 7 8 2 58736 61212
0 994 5 6 1 61217
0 995 7 4 2 56792 58959
0 996 5 1 1 61231
0 997 7 2 2 61218 996
0 998 5 4 1 61235
0 999 7 3 2 56281 58960
0 1000 5 1 1 61241
0 1001 7 1 2 1000 59696
0 1002 5 1 1 1001
0 1003 7 9 2 52925 60112
0 1004 5 2 1 61244
0 1005 7 4 2 55665 61245
0 1006 5 7 1 61255
0 1007 7 1 2 1002 61259
0 1008 5 1 1 1007
0 1009 7 9 2 54138 57384
0 1010 5 4 1 61266
0 1011 7 1 2 1008 61275
0 1012 5 1 1 1011
0 1013 7 1 2 59287 1012
0 1014 5 1 1 1013
0 1015 7 3 2 59840 59387
0 1016 5 3 1 61279
0 1017 7 2 2 48040 61282
0 1018 5 1 1 61285
0 1019 7 2 2 59459 1018
0 1020 5 5 1 61287
0 1021 7 7 2 52221 59646
0 1022 5 9 1 61294
0 1023 7 1 2 61301 59288
0 1024 5 1 1 1023
0 1025 7 1 2 57795 57292
0 1026 5 1 1 1025
0 1027 7 1 2 1024 1026
0 1028 5 1 1 1027
0 1029 7 1 2 61289 1028
0 1030 5 1 1 1029
0 1031 7 4 2 48680 56282
0 1032 5 3 1 61310
0 1033 7 7 2 49509 57303
0 1034 5 34 1 61317
0 1035 7 4 2 61314 61324
0 1036 5 8 1 61358
0 1037 7 1 2 55985 61362
0 1038 5 2 1 1037
0 1039 7 1 2 1030 61370
0 1040 7 1 2 1014 1039
0 1041 5 1 1 1040
0 1042 7 1 2 54433 1041
0 1043 5 1 1 1042
0 1044 7 1 2 61236 1043
0 1045 7 1 2 990 1044
0 1046 5 1 1 1045
0 1047 7 1 2 52749 1046
0 1048 5 1 1 1047
0 1049 7 1 2 56283 58301
0 1050 5 1 1 1049
0 1051 7 2 2 52365 58155
0 1052 5 3 1 61372
0 1053 7 2 2 53145 61373
0 1054 5 2 1 61377
0 1055 7 1 2 48291 61379
0 1056 5 1 1 1055
0 1057 7 1 2 1050 1056
0 1058 5 2 1 1057
0 1059 7 1 2 59564 61381
0 1060 5 1 1 1059
0 1061 7 1 2 56284 59344
0 1062 5 1 1 1061
0 1063 7 2 2 48292 60072
0 1064 5 1 1 61383
0 1065 7 1 2 49390 61384
0 1066 5 1 1 1065
0 1067 7 1 2 1062 1066
0 1068 7 1 2 1060 1067
0 1069 5 1 1 1068
0 1070 7 1 2 58080 1069
0 1071 5 1 1 1070
0 1072 7 1 2 58081 61206
0 1073 5 1 1 1072
0 1074 7 10 2 47752 48293
0 1075 5 5 1 61385
0 1076 7 7 2 48460 49275
0 1077 5 1 1 61400
0 1078 7 1 2 54139 61401
0 1079 7 2 2 59041 1078
0 1080 5 1 1 61407
0 1081 7 1 2 61386 61408
0 1082 5 1 1 1081
0 1083 7 1 2 1073 1082
0 1084 5 2 1 1083
0 1085 7 1 2 61199 61409
0 1086 5 1 1 1085
0 1087 7 4 2 47753 49391
0 1088 5 3 1 61411
0 1089 7 4 2 48041 59605
0 1090 5 2 1 61418
0 1091 7 1 2 61415 61422
0 1092 5 1 1 1091
0 1093 7 1 2 58082 1092
0 1094 5 1 1 1093
0 1095 7 2 2 47754 58083
0 1096 5 1 1 61424
0 1097 7 1 2 59042 61419
0 1098 5 1 1 1097
0 1099 7 1 2 1096 1098
0 1100 5 1 1 1099
0 1101 7 1 2 48461 1100
0 1102 5 1 1 1101
0 1103 7 1 2 1094 1102
0 1104 5 1 1 1103
0 1105 7 1 2 58599 1104
0 1106 5 1 1 1105
0 1107 7 1 2 58084 60073
0 1108 5 1 1 1107
0 1109 7 1 2 59043 58473
0 1110 7 1 2 61170 1109
0 1111 5 1 1 1110
0 1112 7 1 2 1108 1111
0 1113 5 1 1 1112
0 1114 7 1 2 48462 1113
0 1115 5 1 1 1114
0 1116 7 1 2 1106 1115
0 1117 5 1 1 1116
0 1118 7 1 2 48294 1117
0 1119 5 1 1 1118
0 1120 7 1 2 1086 1119
0 1121 7 1 2 1071 1120
0 1122 5 1 1 1121
0 1123 7 1 2 59035 1122
0 1124 5 1 1 1123
0 1125 7 2 2 55986 58908
0 1126 5 1 1 61426
0 1127 7 3 2 54816 59059
0 1128 5 2 1 61428
0 1129 7 1 2 1126 61431
0 1130 5 1 1 1129
0 1131 7 1 2 52750 1130
0 1132 5 1 1 1131
0 1133 7 9 2 52588 49656
0 1134 5 4 1 61433
0 1135 7 4 2 54817 61434
0 1136 7 1 2 56434 61446
0 1137 5 1 1 1136
0 1138 7 1 2 1132 1137
0 1139 5 1 1 1138
0 1140 7 1 2 60565 1139
0 1141 5 1 1 1140
0 1142 7 1 2 55160 1141
0 1143 7 1 2 1124 1142
0 1144 7 1 2 1048 1143
0 1145 7 1 2 948 1144
0 1146 7 1 2 745 1145
0 1147 7 1 2 556 1146
0 1148 5 1 1 1147
0 1149 7 10 2 57559 60035
0 1150 7 1 2 52056 59841
0 1151 5 2 1 1150
0 1152 7 1 2 59842 60170
0 1153 5 1 1 1152
0 1154 7 3 2 61460 1153
0 1155 5 12 1 61462
0 1156 7 1 2 61450 61465
0 1157 5 1 1 1156
0 1158 7 7 2 48042 60346
0 1159 5 3 1 61477
0 1160 7 4 2 50127 61484
0 1161 5 2 1 61487
0 1162 7 1 2 55842 61488
0 1163 5 1 1 1162
0 1164 7 1 2 1157 1163
0 1165 5 1 1 1164
0 1166 7 1 2 50592 1165
0 1167 5 1 1 1166
0 1168 7 13 2 51842 50593
0 1169 5 6 1 61493
0 1170 7 23 2 52926 50128
0 1171 5 54 1 61512
0 1172 7 6 2 52057 53042
0 1173 5 2 1 61589
0 1174 7 2 2 61513 61590
0 1175 5 2 1 61597
0 1176 7 1 2 61506 61599
0 1177 5 1 1 1176
0 1178 7 1 2 55666 1177
0 1179 5 1 1 1178
0 1180 7 4 2 51843 57197
0 1181 5 7 1 61601
0 1182 7 2 2 53923 61605
0 1183 5 3 1 61612
0 1184 7 1 2 60884 61613
0 1185 5 1 1 1184
0 1186 7 1 2 50594 1185
0 1187 5 1 1 1186
0 1188 7 1 2 1179 1187
0 1189 5 1 1 1188
0 1190 7 1 2 52222 1189
0 1191 5 1 1 1190
0 1192 7 1 2 60140 60043
0 1193 5 1 1 1192
0 1194 7 2 2 52058 58814
0 1195 5 4 1 61617
0 1196 7 10 2 51844 53043
0 1197 5 5 1 61623
0 1198 7 1 2 60276 61633
0 1199 5 4 1 1198
0 1200 7 1 2 59843 61638
0 1201 5 1 1 1200
0 1202 7 1 2 61619 1201
0 1203 7 1 2 1193 1202
0 1204 5 1 1 1203
0 1205 7 1 2 50595 1204
0 1206 5 1 1 1205
0 1207 7 1 2 1191 1206
0 1208 5 1 1 1207
0 1209 7 1 2 50337 1208
0 1210 5 1 1 1209
0 1211 7 2 2 1167 1210
0 1212 5 1 1 61642
0 1213 7 1 2 56498 61643
0 1214 5 1 1 1213
0 1215 7 1 2 48838 1214
0 1216 5 1 1 1215
0 1217 7 4 2 54434 61535
0 1218 5 3 1 61644
0 1219 7 14 2 53861 53924
0 1220 5 5 1 61651
0 1221 7 1 2 52927 61665
0 1222 5 5 1 1221
0 1223 7 1 2 58846 61670
0 1224 5 3 1 1223
0 1225 7 2 2 52928 60939
0 1226 5 4 1 61678
0 1227 7 1 2 60688 61680
0 1228 5 1 1 1227
0 1229 7 1 2 61675 1228
0 1230 5 1 1 1229
0 1231 7 1 2 55987 1230
0 1232 5 1 1 1231
0 1233 7 1 2 61648 1232
0 1234 5 1 1 1233
0 1235 7 1 2 48043 1234
0 1236 5 1 1 1235
0 1237 7 2 2 51845 55843
0 1238 5 2 1 61684
0 1239 7 2 2 55667 61685
0 1240 5 1 1 61688
0 1241 7 1 2 56285 1240
0 1242 5 1 1 1241
0 1243 7 6 2 52059 61514
0 1244 5 15 1 61690
0 1245 7 1 2 59177 61696
0 1246 5 1 1 1245
0 1247 7 11 2 49276 61387
0 1248 5 3 1 61711
0 1249 7 4 2 58356 59957
0 1250 5 4 1 61725
0 1251 7 1 2 59292 61726
0 1252 5 1 1 1251
0 1253 7 1 2 61722 1252
0 1254 7 1 2 1246 1253
0 1255 7 1 2 1242 1254
0 1256 7 32 2 49150 53925
0 1257 5 12 1 61733
0 1258 7 5 2 52223 61765
0 1259 5 4 1 61777
0 1260 7 2 2 53044 61778
0 1261 5 11 1 61786
0 1262 7 1 2 61787 60979
0 1263 5 1 1 1262
0 1264 7 1 2 54435 1263
0 1265 5 1 1 1264
0 1266 7 6 2 47755 61734
0 1267 5 4 1 61799
0 1268 7 1 2 55988 61800
0 1269 5 1 1 1268
0 1270 7 1 2 57560 1269
0 1271 5 2 1 1270
0 1272 7 1 2 55727 61809
0 1273 5 1 1 1272
0 1274 7 1 2 1265 1273
0 1275 7 1 2 1255 1274
0 1276 7 1 2 1236 1275
0 1277 5 1 1 1276
0 1278 7 1 2 58726 1277
0 1279 5 1 1 1278
0 1280 7 3 2 56793 56675
0 1281 5 1 1 61811
0 1282 7 12 2 53926 56676
0 1283 5 7 1 61814
0 1284 7 1 2 57198 61826
0 1285 5 12 1 1284
0 1286 7 1 2 59471 61833
0 1287 5 1 1 1286
0 1288 7 1 2 1281 1287
0 1289 5 1 1 1288
0 1290 7 1 2 53862 1289
0 1291 5 1 1 1290
0 1292 7 1 2 56794 61815
0 1293 5 1 1 1292
0 1294 7 1 2 1291 1293
0 1295 5 1 1 1294
0 1296 7 1 2 49091 1295
0 1297 5 1 1 1296
0 1298 7 1 2 52060 61666
0 1299 5 2 1 1298
0 1300 7 6 2 61671 61845
0 1301 5 1 1 61847
0 1302 7 2 2 56677 61848
0 1303 7 1 2 48463 61853
0 1304 5 1 1 1303
0 1305 7 8 2 48044 61735
0 1306 5 8 1 61855
0 1307 7 1 2 54436 61856
0 1308 5 1 1 1307
0 1309 7 1 2 1304 1308
0 1310 5 1 1 1309
0 1311 7 1 2 49392 1310
0 1312 5 1 1 1311
0 1313 7 1 2 1297 1312
0 1314 5 1 1 1313
0 1315 7 1 2 47756 1314
0 1316 5 1 1 1315
0 1317 7 2 2 59426 61652
0 1318 5 4 1 61871
0 1319 7 2 2 50596 61873
0 1320 5 3 1 61877
0 1321 7 1 2 48464 61879
0 1322 5 1 1 1321
0 1323 7 36 2 53927 54437
0 1324 5 8 1 61882
0 1325 7 3 2 52366 61918
0 1326 5 2 1 61926
0 1327 7 1 2 59834 61929
0 1328 5 1 1 1327
0 1329 7 11 2 53928 58357
0 1330 5 3 1 61931
0 1331 7 1 2 48465 61932
0 1332 5 1 1 1331
0 1333 7 1 2 1328 1332
0 1334 5 1 1 1333
0 1335 7 1 2 48045 1334
0 1336 5 1 1 1335
0 1337 7 1 2 1322 1336
0 1338 5 1 1 1337
0 1339 7 1 2 49393 1338
0 1340 5 1 1 1339
0 1341 7 1 2 1316 1340
0 1342 5 1 1 1341
0 1343 7 1 2 55989 1342
0 1344 5 1 1 1343
0 1345 7 7 2 49277 58224
0 1346 7 3 2 48046 61536
0 1347 5 7 1 61952
0 1348 7 3 2 61766 60980
0 1349 5 2 1 61962
0 1350 7 1 2 61955 61963
0 1351 5 1 1 1350
0 1352 7 1 2 61945 1351
0 1353 5 1 1 1352
0 1354 7 3 2 58415 56603
0 1355 5 15 1 61967
0 1356 7 2 2 50129 61968
0 1357 5 6 1 61985
0 1358 7 1 2 47757 61987
0 1359 5 1 1 1358
0 1360 7 5 2 61767 61956
0 1361 7 1 2 60844 61196
0 1362 7 1 2 61993 1361
0 1363 7 2 2 1359 1362
0 1364 5 2 1 61998
0 1365 7 1 2 49394 59178
0 1366 7 1 2 62000 1365
0 1367 5 1 1 1366
0 1368 7 1 2 1353 1367
0 1369 5 1 1 1368
0 1370 7 1 2 54438 1369
0 1371 5 1 1 1370
0 1372 7 11 2 49278 49395
0 1373 5 1 1 62002
0 1374 7 3 2 48466 62003
0 1375 5 1 1 62013
0 1376 7 2 2 48295 60650
0 1377 5 4 1 62016
0 1378 7 1 2 62014 62017
0 1379 5 2 1 1378
0 1380 7 1 2 1371 62022
0 1381 7 1 2 1344 1380
0 1382 5 1 1 1381
0 1383 7 1 2 58085 1382
0 1384 5 1 1 1383
0 1385 7 1 2 1279 1384
0 1386 5 1 1 1385
0 1387 7 1 2 54140 1386
0 1388 5 1 1 1387
0 1389 7 4 2 49396 57385
0 1390 5 3 1 62024
0 1391 7 5 2 53146 57561
0 1392 5 9 1 62031
0 1393 7 1 2 61736 62036
0 1394 5 1 1 1393
0 1395 7 1 2 58559 1394
0 1396 5 1 1 1395
0 1397 7 5 2 52061 58416
0 1398 5 18 1 62045
0 1399 7 7 2 47758 55728
0 1400 5 6 1 62068
0 1401 7 6 2 62046 62075
0 1402 5 6 1 62081
0 1403 7 1 2 1396 62087
0 1404 5 1 1 1403
0 1405 7 1 2 62028 1404
0 1406 5 1 1 1405
0 1407 7 1 2 54439 1406
0 1408 5 1 1 1407
0 1409 7 7 2 52062 50083
0 1410 5 5 1 62093
0 1411 7 6 2 58833 62094
0 1412 5 9 1 62105
0 1413 7 13 2 48296 53929
0 1414 5 1 1 62120
0 1415 7 1 2 62121 58489
0 1416 7 1 2 62111 1415
0 1417 5 1 1 1416
0 1418 7 1 2 1408 1417
0 1419 5 1 1 1418
0 1420 7 1 2 48467 1419
0 1421 5 1 1 1420
0 1422 7 10 2 49397 54440
0 1423 5 2 1 62133
0 1424 7 1 2 58515 62134
0 1425 5 2 1 1424
0 1426 7 1 2 51846 58417
0 1427 5 6 1 1426
0 1428 7 13 2 55729 62147
0 1429 5 15 1 62153
0 1430 7 3 2 54441 62154
0 1431 5 2 1 62181
0 1432 7 1 2 58932 62182
0 1433 5 1 1 1432
0 1434 7 1 2 62023 1433
0 1435 5 1 1 1434
0 1436 7 1 2 48047 1435
0 1437 5 1 1 1436
0 1438 7 1 2 62145 1437
0 1439 5 1 1 1438
0 1440 7 1 2 61537 1439
0 1441 5 1 1 1440
0 1442 7 11 2 49398 53930
0 1443 5 5 1 62186
0 1444 7 3 2 49279 62187
0 1445 5 1 1 62202
0 1446 7 11 2 48297 49151
0 1447 5 2 1 62205
0 1448 7 1 2 54442 62206
0 1449 7 1 2 62203 1448
0 1450 7 1 2 62088 1449
0 1451 5 1 1 1450
0 1452 7 1 2 1441 1451
0 1453 7 1 2 1421 1452
0 1454 5 1 1 1453
0 1455 7 1 2 58086 1454
0 1456 5 1 1 1455
0 1457 7 3 2 50084 57562
0 1458 5 3 1 62218
0 1459 7 1 2 52877 57563
0 1460 5 2 1 1459
0 1461 7 3 2 62221 62224
0 1462 5 2 1 62226
0 1463 7 3 2 59094 62227
0 1464 5 1 1 62231
0 1465 7 1 2 47759 62232
0 1466 5 1 1 1465
0 1467 7 3 2 50085 60770
0 1468 5 2 1 62234
0 1469 7 1 2 57386 62237
0 1470 5 5 1 1469
0 1471 7 1 2 1466 62239
0 1472 5 2 1 1471
0 1473 7 1 2 61737 62244
0 1474 5 1 1 1473
0 1475 7 1 2 56172 58209
0 1476 5 1 1 1475
0 1477 7 1 2 62112 1476
0 1478 5 1 1 1477
0 1479 7 1 2 62184 1478
0 1480 5 1 1 1479
0 1481 7 1 2 61788 1480
0 1482 5 1 1 1481
0 1483 7 6 2 54443 59206
0 1484 5 2 1 62246
0 1485 7 10 2 48048 49092
0 1486 5 1 1 62254
0 1487 7 4 2 59443 62255
0 1488 5 7 1 62264
0 1489 7 1 2 59179 62265
0 1490 5 2 1 1489
0 1491 7 1 2 62252 62275
0 1492 7 1 2 1482 1491
0 1493 7 1 2 1474 1492
0 1494 5 1 1 1493
0 1495 7 1 2 58727 1494
0 1496 5 1 1 1495
0 1497 7 7 2 49399 53863
0 1498 7 3 2 49093 62277
0 1499 5 1 1 62284
0 1500 7 1 2 58703 1499
0 1501 5 1 1 1500
0 1502 7 1 2 47760 1501
0 1503 5 1 1 1502
0 1504 7 2 2 54444 55730
0 1505 5 3 1 62287
0 1506 7 1 2 53147 62289
0 1507 5 1 1 1506
0 1508 7 1 2 54141 1507
0 1509 5 1 1 1508
0 1510 7 1 2 1503 1509
0 1511 5 1 1 1510
0 1512 7 3 2 48468 58087
0 1513 7 1 2 49280 61538
0 1514 5 4 1 1513
0 1515 7 1 2 53045 61768
0 1516 5 13 1 1515
0 1517 7 1 2 48049 62299
0 1518 5 1 1 1517
0 1519 7 1 2 62295 1518
0 1520 5 3 1 1519
0 1521 7 1 2 48298 62312
0 1522 5 1 1 1521
0 1523 7 18 2 48050 53931
0 1524 5 10 1 62315
0 1525 7 3 2 62316 58474
0 1526 5 3 1 62343
0 1527 7 1 2 1522 62346
0 1528 5 2 1 1527
0 1529 7 1 2 62292 62349
0 1530 5 1 1 1529
0 1531 7 1 2 58728 61697
0 1532 5 1 1 1531
0 1533 7 1 2 1530 1532
0 1534 5 1 1 1533
0 1535 7 1 2 1511 1534
0 1536 5 1 1 1535
0 1537 7 1 2 59207 60651
0 1538 5 1 1 1537
0 1539 7 1 2 62185 1538
0 1540 5 1 1 1539
0 1541 7 1 2 48051 1540
0 1542 5 1 1 1541
0 1543 7 1 2 59180 60965
0 1544 5 1 1 1543
0 1545 7 14 2 53148 50597
0 1546 5 12 1 62351
0 1547 7 5 2 52367 62352
0 1548 5 4 1 62377
0 1549 7 1 2 55990 62382
0 1550 5 1 1 1549
0 1551 7 1 2 1544 1550
0 1552 7 1 2 1542 1551
0 1553 5 1 1 1552
0 1554 7 1 2 58729 61539
0 1555 7 1 2 1553 1554
0 1556 5 1 1 1555
0 1557 7 1 2 1536 1556
0 1558 7 1 2 1496 1557
0 1559 7 1 2 1456 1558
0 1560 7 1 2 1388 1559
0 1561 5 1 1 1560
0 1562 7 1 2 53410 1561
0 1563 5 1 1 1562
0 1564 7 1 2 1216 1563
0 1565 5 1 1 1564
0 1566 7 1 2 54818 1565
0 1567 5 1 1 1566
0 1568 7 2 2 59872 59311
0 1569 5 1 1 62386
0 1570 7 5 2 55844 57199
0 1571 5 26 1 62388
0 1572 7 4 2 53411 53932
0 1573 7 1 2 62393 62419
0 1574 5 1 1 1573
0 1575 7 1 2 1569 1574
0 1576 5 1 1 1575
0 1577 7 1 2 56286 1576
0 1578 5 1 1 1577
0 1579 7 1 2 59248 62420
0 1580 5 1 1 1579
0 1581 7 1 2 1578 1580
0 1582 5 1 1 1581
0 1583 7 1 2 48681 1582
0 1584 5 1 1 1583
0 1585 7 1 2 58909 62387
0 1586 5 1 1 1585
0 1587 7 1 2 1584 1586
0 1588 5 1 1 1587
0 1589 7 1 2 54142 1588
0 1590 5 1 1 1589
0 1591 7 8 2 52224 57200
0 1592 5 11 1 62423
0 1593 7 7 2 60074 62431
0 1594 5 2 1 62442
0 1595 7 9 2 55991 62443
0 1596 5 1 1 62451
0 1597 7 1 2 56287 62452
0 1598 5 3 1 1597
0 1599 7 2 2 56974 62460
0 1600 5 4 1 62463
0 1601 7 44 2 52589 53412
0 1602 5 79 1 62469
0 1603 7 8 2 50898 62513
0 1604 5 2 1 62592
0 1605 7 13 2 53933 50338
0 1606 5 3 1 62602
0 1607 7 1 2 62593 62603
0 1608 7 1 2 62465 1607
0 1609 5 1 1 1608
0 1610 7 1 2 1590 1609
0 1611 5 1 1 1610
0 1612 7 1 2 54445 1611
0 1613 5 1 1 1612
0 1614 7 1 2 55992 61834
0 1615 5 2 1 1614
0 1616 7 1 2 57564 62618
0 1617 5 2 1 1616
0 1618 7 2 2 56795 62620
0 1619 5 1 1 62622
0 1620 7 1 2 50598 62594
0 1621 7 1 2 62623 1620
0 1622 5 1 1 1621
0 1623 7 1 2 1613 1622
0 1624 5 1 1 1623
0 1625 7 1 2 47761 1624
0 1626 5 1 1 1625
0 1627 7 2 2 50599 58237
0 1628 7 1 2 61738 62624
0 1629 5 1 1 1628
0 1630 7 20 2 50339 54446
0 1631 5 1 1 62626
0 1632 7 1 2 56678 62627
0 1633 5 1 1 1632
0 1634 7 1 2 1629 1633
0 1635 5 1 1 1634
0 1636 7 1 2 58933 1635
0 1637 5 1 1 1636
0 1638 7 7 2 49400 50600
0 1639 7 3 2 48469 62646
0 1640 7 2 2 48299 61540
0 1641 5 4 1 62656
0 1642 7 2 2 62296 62658
0 1643 5 4 1 62662
0 1644 7 2 2 59086 62663
0 1645 5 1 1 62668
0 1646 7 2 2 54143 1645
0 1647 7 1 2 62653 62670
0 1648 5 1 1 1647
0 1649 7 1 2 1637 1648
0 1650 5 1 1 1649
0 1651 7 1 2 62595 1650
0 1652 5 1 1 1651
0 1653 7 1 2 1626 1652
0 1654 5 1 1 1653
0 1655 7 1 2 56499 1654
0 1656 5 1 1 1655
0 1657 7 19 2 49657 50899
0 1658 5 2 1 62672
0 1659 7 3 2 53934 62394
0 1660 5 2 1 62693
0 1661 7 1 2 59305 62696
0 1662 5 1 1 1661
0 1663 7 1 2 54144 1662
0 1664 5 1 1 1663
0 1665 7 2 2 62032 62619
0 1666 5 1 1 62698
0 1667 7 1 2 47762 1666
0 1668 5 1 1 1667
0 1669 7 1 2 1664 1668
0 1670 5 1 1 1669
0 1671 7 1 2 50601 1670
0 1672 5 1 1 1671
0 1673 7 39 2 47763 53935
0 1674 5 8 1 62700
0 1675 7 2 2 52063 62739
0 1676 5 2 1 62747
0 1677 7 1 2 52929 62748
0 1678 5 11 1 1677
0 1679 7 1 2 62751 62628
0 1680 5 2 1 1679
0 1681 7 1 2 1672 62762
0 1682 5 1 1 1681
0 1683 7 1 2 62673 1682
0 1684 5 1 1 1683
0 1685 7 5 2 49658 59122
0 1686 5 1 1 62764
0 1687 7 4 2 49401 53413
0 1688 7 11 2 53936 58651
0 1689 5 1 1 62773
0 1690 7 2 2 62774 59249
0 1691 7 1 2 62769 62784
0 1692 5 1 1 1691
0 1693 7 1 2 1686 1692
0 1694 5 1 1 1693
0 1695 7 1 2 58504 1694
0 1696 5 1 1 1695
0 1697 7 1 2 1684 1696
0 1698 5 1 1 1697
0 1699 7 1 2 58088 1698
0 1700 5 1 1 1699
0 1701 7 4 2 49152 60053
0 1702 5 4 1 62786
0 1703 7 1 2 48300 62300
0 1704 5 1 1 1703
0 1705 7 3 2 62790 1704
0 1706 5 12 1 62794
0 1707 7 1 2 56173 62795
0 1708 5 1 1 1707
0 1709 7 1 2 47764 1708
0 1710 5 1 1 1709
0 1711 7 2 2 58238 61789
0 1712 5 2 1 62809
0 1713 7 4 2 61541 59565
0 1714 5 1 1 62813
0 1715 7 2 2 55993 62814
0 1716 5 2 1 62817
0 1717 7 1 2 62811 62819
0 1718 7 1 2 1710 1717
0 1719 5 1 1 1718
0 1720 7 1 2 50602 1719
0 1721 5 1 1 1720
0 1722 7 1 2 62763 1721
0 1723 5 1 1 1722
0 1724 7 11 2 48682 57856
0 1725 5 4 1 62821
0 1726 7 2 2 52751 62832
0 1727 5 10 1 62836
0 1728 7 1 2 50900 62838
0 1729 7 1 2 1723 1728
0 1730 5 1 1 1729
0 1731 7 1 2 1700 1730
0 1732 7 1 2 1656 1731
0 1733 5 1 1 1732
0 1734 7 1 2 55731 1733
0 1735 5 1 1 1734
0 1736 7 1 2 48839 58704
0 1737 5 1 1 1736
0 1738 7 5 2 50603 60277
0 1739 7 1 2 56796 62848
0 1740 5 1 1 1739
0 1741 7 5 2 54447 58358
0 1742 5 2 1 62853
0 1743 7 2 2 50130 56288
0 1744 7 1 2 62854 62860
0 1745 5 1 1 1744
0 1746 7 1 2 1740 1745
0 1747 5 1 1 1746
0 1748 7 1 2 61060 1747
0 1749 5 1 1 1748
0 1750 7 5 2 48052 50340
0 1751 7 3 2 54448 58934
0 1752 7 1 2 62862 62867
0 1753 5 1 1 1752
0 1754 7 1 2 1749 1753
0 1755 5 1 1 1754
0 1756 7 1 2 49153 1755
0 1757 5 1 1 1756
0 1758 7 2 2 57387 59366
0 1759 5 2 1 62870
0 1760 7 1 2 50604 62333
0 1761 5 2 1 1760
0 1762 7 1 2 59379 1631
0 1763 5 6 1 1762
0 1764 7 1 2 55994 62876
0 1765 7 1 2 62874 1764
0 1766 5 1 1 1765
0 1767 7 1 2 62872 1766
0 1768 5 1 1 1767
0 1769 7 1 2 56797 1768
0 1770 5 1 1 1769
0 1771 7 1 2 1757 1770
0 1772 5 1 1 1771
0 1773 7 1 2 56500 1772
0 1774 5 1 1 1773
0 1775 7 1 2 1737 1774
0 1776 5 1 1 1775
0 1777 7 1 2 62514 1776
0 1778 5 1 1 1777
0 1779 7 57 2 48683 49659
0 1780 5 59 1 62882
0 1781 7 3 2 62515 57857
0 1782 5 2 1 62998
0 1783 7 4 2 62939 63001
0 1784 5 15 1 63003
0 1785 7 1 2 52752 63004
0 1786 5 4 1 1785
0 1787 7 2 2 52930 62334
0 1788 5 6 1 63026
0 1789 7 1 2 60319 63028
0 1790 5 5 1 1789
0 1791 7 2 2 56174 63034
0 1792 7 1 2 50605 63039
0 1793 5 1 1 1792
0 1794 7 1 2 55995 58705
0 1795 7 1 2 1793 1794
0 1796 5 1 1 1795
0 1797 7 3 2 56975 975
0 1798 5 1 1 63041
0 1799 7 1 2 50606 1798
0 1800 5 1 1 1799
0 1801 7 1 2 56175 57201
0 1802 5 2 1 1801
0 1803 7 1 2 62629 63044
0 1804 5 1 1 1803
0 1805 7 1 2 1800 1804
0 1806 7 1 2 1796 1805
0 1807 5 1 1 1806
0 1808 7 1 2 63022 1807
0 1809 5 1 1 1808
0 1810 7 1 2 58193 62849
0 1811 5 1 1 1810
0 1812 7 3 2 58198 59958
0 1813 5 1 1 63046
0 1814 7 1 2 50341 63047
0 1815 5 1 1 1814
0 1816 7 1 2 1811 1815
0 1817 5 3 1 1816
0 1818 7 4 2 49094 49510
0 1819 7 2 2 48684 63052
0 1820 7 1 2 62004 58132
0 1821 7 1 2 63056 1820
0 1822 5 1 1 1821
0 1823 7 1 2 52753 1822
0 1824 5 1 1 1823
0 1825 7 1 2 63049 1824
0 1826 5 1 1 1825
0 1827 7 7 2 52754 62940
0 1828 5 28 1 63058
0 1829 7 3 2 56501 63065
0 1830 5 1 1 63093
0 1831 7 1 2 58706 63094
0 1832 5 1 1 1831
0 1833 7 2 2 48301 55732
0 1834 5 1 1 63096
0 1835 7 2 2 49281 63097
0 1836 5 3 1 63098
0 1837 7 1 2 57123 63099
0 1838 5 3 1 1837
0 1839 7 5 2 48840 54145
0 1840 7 1 2 54449 63106
0 1841 7 1 2 63103 1840
0 1842 5 1 1 1841
0 1843 7 1 2 1832 1842
0 1844 7 1 2 1826 1843
0 1845 7 1 2 1809 1844
0 1846 7 1 2 1778 1845
0 1847 5 1 1 1846
0 1848 7 1 2 50901 1847
0 1849 5 1 1 1848
0 1850 7 1 2 55845 62335
0 1851 5 5 1 1850
0 1852 7 1 2 57812 63111
0 1853 5 2 1 1852
0 1854 7 7 2 52064 57565
0 1855 5 3 1 63118
0 1856 7 7 2 50131 57566
0 1857 5 6 1 63128
0 1858 7 4 2 55996 63135
0 1859 7 3 2 63125 63141
0 1860 5 2 1 63145
0 1861 7 1 2 63116 63148
0 1862 5 1 1 1861
0 1863 7 1 2 50607 1862
0 1864 5 1 1 1863
0 1865 7 4 2 54450 59959
0 1866 5 4 1 63150
0 1867 7 1 2 50342 63151
0 1868 5 1 1 1867
0 1869 7 1 2 1864 1868
0 1870 5 1 1 1869
0 1871 7 2 2 50902 63023
0 1872 5 1 1 63158
0 1873 7 8 2 62516 56798
0 1874 7 1 2 63160 59282
0 1875 5 1 1 1874
0 1876 7 1 2 1872 1875
0 1877 5 1 1 1876
0 1878 7 1 2 1870 1877
0 1879 5 1 1 1878
0 1880 7 18 2 50132 54146
0 1881 5 3 1 63168
0 1882 7 1 2 59076 63169
0 1883 5 1 1 1882
0 1884 7 5 2 50343 57388
0 1885 5 2 1 63189
0 1886 7 1 2 59960 63190
0 1887 5 2 1 1886
0 1888 7 1 2 1883 63196
0 1889 5 1 1 1888
0 1890 7 1 2 62596 1889
0 1891 5 1 1 1890
0 1892 7 16 2 48685 53414
0 1893 5 4 1 63198
0 1894 7 10 2 53937 55997
0 1895 5 5 1 63218
0 1896 7 2 2 54147 63219
0 1897 5 2 1 63233
0 1898 7 1 2 63199 63234
0 1899 5 1 1 1898
0 1900 7 1 2 1891 1899
0 1901 5 1 1 1900
0 1902 7 1 2 54451 1901
0 1903 5 1 1 1902
0 1904 7 4 2 53938 59367
0 1905 5 1 1 63237
0 1906 7 14 2 48053 48302
0 1907 5 3 1 63241
0 1908 7 4 2 63242 59335
0 1909 5 1 1 63258
0 1910 7 1 2 63259 62597
0 1911 7 1 2 63238 1910
0 1912 5 1 1 1911
0 1913 7 1 2 1903 1912
0 1914 5 1 1 1913
0 1915 7 1 2 56502 1914
0 1916 5 1 1 1915
0 1917 7 1 2 50608 63159
0 1918 5 1 1 1917
0 1919 7 1 2 1916 1918
0 1920 5 1 1 1919
0 1921 7 1 2 56289 1920
0 1922 5 1 1 1921
0 1923 7 1 2 1879 1922
0 1924 5 1 1 1923
0 1925 7 1 2 58600 1924
0 1926 5 1 1 1925
0 1927 7 3 2 48054 61225
0 1928 5 1 1 63262
0 1929 7 5 2 53939 56290
0 1930 5 3 1 63265
0 1931 7 2 2 61161 63270
0 1932 5 2 1 63273
0 1933 7 14 2 48303 54452
0 1934 5 1 1 63277
0 1935 7 3 2 50344 63278
0 1936 7 1 2 63275 63291
0 1937 7 1 2 63263 1936
0 1938 5 1 1 1937
0 1939 7 4 2 57970 59052
0 1940 5 20 1 63294
0 1941 7 1 2 62517 63298
0 1942 5 2 1 1941
0 1943 7 1 2 63059 63318
0 1944 5 2 1 1943
0 1945 7 1 2 58345 62850
0 1946 7 1 2 63320 1945
0 1947 5 1 1 1946
0 1948 7 1 2 1938 1947
0 1949 5 1 1 1948
0 1950 7 1 2 50903 1949
0 1951 5 1 1 1950
0 1952 7 2 2 48055 48686
0 1953 7 5 2 53415 54148
0 1954 7 3 2 61883 63324
0 1955 7 2 2 56503 63329
0 1956 7 3 2 56291 63332
0 1957 7 1 2 63322 63334
0 1958 5 1 1 1957
0 1959 7 1 2 1951 1958
0 1960 5 1 1 1959
0 1961 7 1 2 58302 1960
0 1962 5 1 1 1961
0 1963 7 1 2 57971 58513
0 1964 5 1 1 1963
0 1965 7 1 2 61226 1964
0 1966 5 1 1 1965
0 1967 7 1 2 63060 1966
0 1968 5 1 1 1967
0 1969 7 1 2 62851 1968
0 1970 5 1 1 1969
0 1971 7 2 2 59961 61227
0 1972 7 10 2 48470 54453
0 1973 7 1 2 63339 62863
0 1974 7 1 2 63337 1973
0 1975 5 1 1 1974
0 1976 7 1 2 1970 1975
0 1977 5 1 1 1976
0 1978 7 1 2 50904 1977
0 1979 5 1 1 1978
0 1980 7 4 2 48304 48687
0 1981 5 1 1 63349
0 1982 7 3 2 48056 63350
0 1983 7 1 2 63333 63353
0 1984 5 1 1 1983
0 1985 7 1 2 1979 1984
0 1986 5 1 1 1985
0 1987 7 1 2 58159 1986
0 1988 5 1 1 1987
0 1989 7 5 2 48057 48471
0 1990 7 2 2 63356 63351
0 1991 7 1 2 63330 63361
0 1992 5 1 1 1991
0 1993 7 1 2 48570 62598
0 1994 7 1 2 63050 1993
0 1995 5 1 1 1994
0 1996 7 1 2 1992 1995
0 1997 5 1 1 1996
0 1998 7 1 2 58499 1997
0 1999 5 1 1 1998
0 2000 7 3 2 49095 58475
0 2001 7 3 2 49511 53864
0 2002 7 2 2 49402 63366
0 2003 7 2 2 63363 63369
0 2004 5 2 1 63371
0 2005 7 1 2 52590 63373
0 2006 5 1 1 2005
0 2007 7 1 2 62674 63051
0 2008 5 1 1 2007
0 2009 7 5 2 48305 48571
0 2010 7 2 2 63375 63357
0 2011 7 1 2 63331 63380
0 2012 5 1 1 2011
0 2013 7 1 2 2008 2012
0 2014 5 1 1 2013
0 2015 7 1 2 2006 2014
0 2016 5 1 1 2015
0 2017 7 1 2 51197 2016
0 2018 7 1 2 1999 2017
0 2019 7 1 2 1988 2018
0 2020 7 1 2 1962 2019
0 2021 7 1 2 1926 2020
0 2022 7 1 2 1849 2021
0 2023 7 1 2 1735 2022
0 2024 7 1 2 1567 2023
0 2025 5 1 1 2024
0 2026 7 1 2 1148 2025
0 2027 5 1 1 2026
0 2028 7 3 2 52878 50345
0 2029 5 2 1 63382
0 2030 7 4 2 60096 63383
0 2031 5 1 1 63387
0 2032 7 2 2 50133 63388
0 2033 5 1 1 63391
0 2034 7 1 2 48306 2033
0 2035 5 1 1 2034
0 2036 7 1 2 53046 60735
0 2037 5 1 1 2036
0 2038 7 2 2 60816 2037
0 2039 5 1 1 63393
0 2040 7 3 2 2035 2039
0 2041 7 1 2 50905 63395
0 2042 5 1 1 2041
0 2043 7 1 2 53416 60845
0 2044 5 1 1 2043
0 2045 7 1 2 2042 2044
0 2046 5 1 1 2045
0 2047 7 1 2 48841 2046
0 2048 5 1 1 2047
0 2049 7 10 2 49660 54149
0 2050 5 4 1 63398
0 2051 7 2 2 52591 63399
0 2052 7 2 2 54819 60846
0 2053 7 1 2 63412 63414
0 2054 5 1 1 2053
0 2055 7 1 2 2048 2054
0 2056 5 1 1 2055
0 2057 7 1 2 50609 2056
0 2058 5 1 1 2057
0 2059 7 10 2 48842 53417
0 2060 5 4 1 63416
0 2061 7 34 2 54454 54820
0 2062 5 11 1 63430
0 2063 7 2 2 63431 61435
0 2064 5 3 1 63475
0 2065 7 1 2 63426 63477
0 2066 5 3 1 2065
0 2067 7 1 2 60674 63480
0 2068 5 1 1 2067
0 2069 7 1 2 2058 2068
0 2070 5 1 1 2069
0 2071 7 1 2 55161 2070
0 2072 5 1 1 2071
0 2073 7 9 2 48843 51198
0 2074 5 1 1 63483
0 2075 7 3 2 54821 63484
0 2076 7 3 2 59606 60025
0 2077 5 3 1 63495
0 2078 7 1 2 63492 63498
0 2079 5 1 1 2078
0 2080 7 1 2 2072 2079
0 2081 5 1 1 2080
0 2082 7 1 2 57202 2081
0 2083 5 1 1 2082
0 2084 7 41 2 54455 50906
0 2085 5 11 1 63501
0 2086 7 8 2 54150 63502
0 2087 5 3 1 63553
0 2088 7 1 2 63485 63554
0 2089 5 1 1 2088
0 2090 7 13 2 49661 54822
0 2091 5 1 1 63564
0 2092 7 7 2 52592 54456
0 2093 5 1 1 63577
0 2094 7 5 2 56604 58834
0 2095 5 1 1 63584
0 2096 7 3 2 53940 60524
0 2097 7 1 2 60105 63589
0 2098 7 1 2 63585 2097
0 2099 5 1 1 2098
0 2100 7 1 2 2093 2099
0 2101 5 1 1 2100
0 2102 7 1 2 63565 2101
0 2103 5 1 1 2102
0 2104 7 1 2 48844 60509
0 2105 5 1 1 2104
0 2106 7 1 2 2103 2105
0 2107 5 1 1 2106
0 2108 7 8 2 53149 55162
0 2109 5 1 1 63592
0 2110 7 1 2 52368 63593
0 2111 7 1 2 2107 2110
0 2112 5 1 1 2111
0 2113 7 1 2 2089 2112
0 2114 5 1 1 2113
0 2115 7 1 2 57972 2114
0 2116 5 1 1 2115
0 2117 7 22 2 50134 50610
0 2118 5 12 1 63600
0 2119 7 15 2 50346 50907
0 2120 5 1 1 63634
0 2121 7 1 2 63601 63635
0 2122 5 3 1 2121
0 2123 7 16 2 53418 50347
0 2124 5 3 1 63652
0 2125 7 7 2 53419 50135
0 2126 5 3 1 63671
0 2127 7 4 2 50348 59123
0 2128 5 3 1 63681
0 2129 7 1 2 63678 63685
0 2130 5 3 1 2129
0 2131 7 1 2 55668 63688
0 2132 5 1 1 2131
0 2133 7 1 2 63668 2132
0 2134 5 1 1 2133
0 2135 7 1 2 51847 2134
0 2136 5 1 1 2135
0 2137 7 1 2 63649 2136
0 2138 5 1 1 2137
0 2139 7 1 2 56605 2138
0 2140 5 1 1 2139
0 2141 7 6 2 53420 60182
0 2142 5 2 1 63691
0 2143 7 1 2 55669 63692
0 2144 5 1 1 2143
0 2145 7 1 2 2140 2144
0 2146 5 1 1 2145
0 2147 7 1 2 57567 2146
0 2148 5 1 1 2147
0 2149 7 8 2 50908 56606
0 2150 5 1 1 63699
0 2151 7 1 2 63602 63700
0 2152 5 2 1 2151
0 2153 7 1 2 63669 63707
0 2154 5 1 1 2153
0 2155 7 1 2 51848 2154
0 2156 5 1 1 2155
0 2157 7 2 2 56679 60652
0 2158 5 3 1 63709
0 2159 7 1 2 63689 63711
0 2160 5 1 1 2159
0 2161 7 1 2 2160 63650
0 2162 7 1 2 2156 2161
0 2163 5 1 1 2162
0 2164 7 1 2 55846 2163
0 2165 5 1 1 2164
0 2166 7 1 2 62941 60583
0 2167 5 1 1 2166
0 2168 7 1 2 60230 60780
0 2169 5 1 1 2168
0 2170 7 1 2 55847 2169
0 2171 5 1 1 2170
0 2172 7 1 2 60808 2171
0 2173 5 1 1 2172
0 2174 7 1 2 53421 2173
0 2175 5 1 1 2174
0 2176 7 1 2 2167 2175
0 2177 7 1 2 2165 2176
0 2178 7 1 2 2148 2177
0 2179 5 1 1 2178
0 2180 7 1 2 55163 2179
0 2181 5 1 1 2180
0 2182 7 33 2 54823 51199
0 2183 5 6 1 63714
0 2184 7 2 2 54457 63142
0 2185 7 12 2 51849 50349
0 2186 5 6 1 63755
0 2187 7 3 2 63767 60765
0 2188 7 1 2 60626 63773
0 2189 7 1 2 63753 2188
0 2190 5 1 1 2189
0 2191 7 1 2 63715 2190
0 2192 5 1 1 2191
0 2193 7 1 2 2181 2192
0 2194 5 1 1 2193
0 2195 7 1 2 48845 2194
0 2196 5 1 1 2195
0 2197 7 18 2 50611 55164
0 2198 7 5 2 53422 63776
0 2199 5 4 1 63794
0 2200 7 8 2 54824 55670
0 2201 7 1 2 51200 63803
0 2202 5 1 1 2201
0 2203 7 1 2 63799 2202
0 2204 5 1 1 2203
0 2205 7 1 2 48846 2204
0 2206 5 1 1 2205
0 2207 7 34 2 54825 55165
0 2208 5 6 1 63811
0 2209 7 3 2 50612 63812
0 2210 7 1 2 63413 63851
0 2211 5 1 1 2210
0 2212 7 1 2 2206 2211
0 2213 5 1 1 2212
0 2214 7 1 2 60892 2213
0 2215 5 1 1 2214
0 2216 7 5 2 55166 63432
0 2217 7 1 2 63854 61436
0 2218 7 1 2 60831 2217
0 2219 5 1 1 2218
0 2220 7 1 2 2215 2219
0 2221 7 1 2 2196 2220
0 2222 7 1 2 2116 2221
0 2223 7 1 2 2083 2222
0 2224 5 1 1 2223
0 2225 7 1 2 61325 2224
0 2226 5 1 1 2225
0 2227 7 6 2 54458 60370
0 2228 5 1 1 63859
0 2229 7 1 2 47765 63860
0 2230 5 1 1 2229
0 2231 7 1 2 50909 2230
0 2232 5 3 1 2231
0 2233 7 2 2 55733 63865
0 2234 5 1 1 63868
0 2235 7 1 2 53941 61153
0 2236 5 1 1 2235
0 2237 7 1 2 58707 2236
0 2238 5 3 1 2237
0 2239 7 1 2 57084 63870
0 2240 5 1 1 2239
0 2241 7 6 2 53942 56504
0 2242 5 1 1 63873
0 2243 7 2 2 50350 62740
0 2244 5 11 1 63879
0 2245 7 3 2 57389 63881
0 2246 5 1 1 63892
0 2247 7 2 2 54459 63893
0 2248 5 2 1 63895
0 2249 7 1 2 2242 63897
0 2250 5 1 1 2249
0 2251 7 1 2 56292 2250
0 2252 5 1 1 2251
0 2253 7 1 2 2240 2252
0 2254 5 1 1 2253
0 2255 7 1 2 56680 2254
0 2256 5 1 1 2255
0 2257 7 2 2 47766 62395
0 2258 5 1 1 63899
0 2259 7 1 2 2258 60406
0 2260 5 3 1 2259
0 2261 7 1 2 54460 63901
0 2262 5 1 1 2261
0 2263 7 1 2 61061 62444
0 2264 5 1 1 2263
0 2265 7 1 2 2262 2264
0 2266 5 1 1 2265
0 2267 7 1 2 57085 2266
0 2268 5 1 1 2267
0 2269 7 3 2 59607 62122
0 2270 5 4 1 63904
0 2271 7 2 2 48307 60371
0 2272 5 6 1 63911
0 2273 7 1 2 53047 63913
0 2274 5 3 1 2273
0 2275 7 2 2 60407 61395
0 2276 5 3 1 63922
0 2277 7 1 2 57124 63924
0 2278 7 1 2 63919 2277
0 2279 5 1 1 2278
0 2280 7 1 2 63907 2279
0 2281 5 1 1 2280
0 2282 7 1 2 59472 2281
0 2283 5 1 1 2282
0 2284 7 1 2 57299 2283
0 2285 7 1 2 2268 2284
0 2286 7 1 2 2256 2285
0 2287 5 1 1 2286
0 2288 7 1 2 63869 2287
0 2289 5 1 1 2288
0 2290 7 4 2 50136 58418
0 2291 5 20 1 63927
0 2292 7 1 2 58652 59097
0 2293 5 1 1 2292
0 2294 7 1 2 63 2293
0 2295 5 1 1 2294
0 2296 7 1 2 47767 2295
0 2297 5 1 1 2296
0 2298 7 5 2 48058 62207
0 2299 5 3 1 63951
0 2300 7 1 2 61009 63952
0 2301 5 3 1 2300
0 2302 7 1 2 2297 63959
0 2303 5 1 1 2302
0 2304 7 1 2 56293 2303
0 2305 5 1 1 2304
0 2306 7 9 2 48308 59336
0 2307 5 5 1 63962
0 2308 7 10 2 49154 54461
0 2309 5 4 1 63976
0 2310 7 1 2 63971 63986
0 2311 5 1 1 2310
0 2312 7 1 2 48059 2311
0 2313 5 1 1 2312
0 2314 7 22 2 54462 55998
0 2315 5 10 1 63990
0 2316 7 3 2 48309 58476
0 2317 5 4 1 64022
0 2318 7 1 2 58708 64025
0 2319 5 3 1 2318
0 2320 7 1 2 47768 64029
0 2321 5 1 1 2320
0 2322 7 1 2 64012 2321
0 2323 7 1 2 2313 2322
0 2324 5 1 1 2323
0 2325 7 1 2 57086 2324
0 2326 5 1 1 2325
0 2327 7 1 2 2305 2326
0 2328 5 1 1 2327
0 2329 7 1 2 63931 2328
0 2330 5 1 1 2329
0 2331 7 4 2 49512 55999
0 2332 5 2 1 64032
0 2333 7 2 2 48572 56000
0 2334 5 1 1 64038
0 2335 7 2 2 64036 2334
0 2336 5 2 1 64040
0 2337 7 1 2 64041 63960
0 2338 5 1 1 2337
0 2339 7 1 2 54151 2338
0 2340 5 1 1 2339
0 2341 7 2 2 50351 61942
0 2342 5 8 1 64044
0 2343 7 1 2 47769 64046
0 2344 5 3 1 2343
0 2345 7 2 2 60408 64054
0 2346 5 5 1 64057
0 2347 7 1 2 50613 64058
0 2348 5 1 1 2347
0 2349 7 1 2 56505 2348
0 2350 5 1 1 2349
0 2351 7 1 2 2340 2350
0 2352 5 1 1 2351
0 2353 7 1 2 56294 2352
0 2354 5 1 1 2353
0 2355 7 2 2 64013 61113
0 2356 7 2 2 54463 64047
0 2357 7 1 2 59962 64066
0 2358 5 1 1 2357
0 2359 7 1 2 64064 2358
0 2360 5 1 1 2359
0 2361 7 1 2 57087 2360
0 2362 5 1 1 2361
0 2363 7 10 2 54152 58359
0 2364 7 3 2 62701 64068
0 2365 5 2 1 64078
0 2366 7 1 2 59473 64079
0 2367 5 1 1 2366
0 2368 7 4 2 54153 57088
0 2369 5 1 1 64083
0 2370 7 1 2 61727 64084
0 2371 5 1 1 2370
0 2372 7 1 2 2367 2371
0 2373 5 1 1 2372
0 2374 7 1 2 56001 2373
0 2375 5 1 1 2374
0 2376 7 3 2 64048 59963
0 2377 7 1 2 54464 57796
0 2378 7 1 2 64087 2377
0 2379 5 1 1 2378
0 2380 7 1 2 57300 2379
0 2381 7 1 2 2375 2380
0 2382 7 1 2 2362 2381
0 2383 5 1 1 2382
0 2384 7 1 2 56681 2383
0 2385 5 1 1 2384
0 2386 7 2 2 57568 57789
0 2387 5 1 1 64090
0 2388 7 3 2 61069 64091
0 2389 5 1 1 64092
0 2390 7 1 2 54465 2389
0 2391 5 1 1 2390
0 2392 7 1 2 59098 64059
0 2393 5 1 1 2392
0 2394 7 1 2 2391 2393
0 2395 5 1 1 2394
0 2396 7 1 2 57089 2395
0 2397 5 1 1 2396
0 2398 7 1 2 2385 2397
0 2399 7 1 2 2354 2398
0 2400 7 1 2 2330 2399
0 2401 7 1 2 2289 2400
0 2402 5 1 1 2401
0 2403 7 1 2 54826 2402
0 2404 5 1 1 2403
0 2405 7 2 2 56506 58576
0 2406 5 5 1 64095
0 2407 7 1 2 57125 57719
0 2408 5 1 1 2407
0 2409 7 1 2 64097 2408
0 2410 5 2 1 2409
0 2411 7 4 2 54827 59964
0 2412 5 2 1 64104
0 2413 7 1 2 60372 62855
0 2414 5 2 1 2413
0 2415 7 1 2 64108 64110
0 2416 7 1 2 2234 2415
0 2417 5 1 1 2416
0 2418 7 1 2 64102 2417
0 2419 5 1 1 2418
0 2420 7 1 2 50910 1689
0 2421 5 4 1 2420
0 2422 7 1 2 56682 64112
0 2423 7 1 2 64096 2422
0 2424 5 1 1 2423
0 2425 7 1 2 2419 2424
0 2426 7 1 2 2404 2425
0 2427 5 1 1 2426
0 2428 7 1 2 58998 2427
0 2429 5 1 1 2428
0 2430 7 1 2 55432 2429
0 2431 7 1 2 2226 2430
0 2432 7 1 2 2027 2431
0 2433 5 1 1 2432
0 2434 7 11 2 55167 62518
0 2435 7 26 2 54154 54828
0 2436 5 6 1 64127
0 2437 7 4 2 48060 64128
0 2438 5 1 1 64159
0 2439 7 3 2 49155 49513
0 2440 5 2 1 64163
0 2441 7 1 2 2438 64166
0 2442 5 1 1 2441
0 2443 7 1 2 62702 2442
0 2444 5 1 1 2443
0 2445 7 11 2 49514 54155
0 2446 5 1 1 64168
0 2447 7 1 2 48061 64169
0 2448 5 1 1 2447
0 2449 7 1 2 2444 2448
0 2450 5 1 1 2449
0 2451 7 1 2 49282 2450
0 2452 5 1 1 2451
0 2453 7 3 2 48062 64164
0 2454 5 1 1 64179
0 2455 7 1 2 60373 64180
0 2456 5 1 1 2455
0 2457 7 1 2 2452 2456
0 2458 5 1 1 2457
0 2459 7 1 2 48310 2458
0 2460 5 1 1 2459
0 2461 7 2 2 61739 61420
0 2462 5 4 1 64182
0 2463 7 1 2 50911 64184
0 2464 5 1 1 2463
0 2465 7 1 2 49515 2464
0 2466 5 1 1 2465
0 2467 7 1 2 2460 2466
0 2468 5 1 1 2467
0 2469 7 1 2 54466 2468
0 2470 5 1 1 2469
0 2471 7 16 2 49516 54829
0 2472 5 2 1 64188
0 2473 7 5 2 50352 61769
0 2474 5 14 1 64206
0 2475 7 2 2 48063 64211
0 2476 5 3 1 64225
0 2477 7 1 2 47770 64226
0 2478 5 1 1 2477
0 2479 7 1 2 59297 2478
0 2480 5 1 1 2479
0 2481 7 1 2 64189 2480
0 2482 5 1 1 2481
0 2483 7 1 2 2470 2482
0 2484 5 1 1 2483
0 2485 7 1 2 48573 2484
0 2486 5 1 1 2485
0 2487 7 14 2 49517 54467
0 2488 5 1 1 64230
0 2489 7 4 2 53943 64129
0 2490 5 1 1 64244
0 2491 7 2 2 64231 64245
0 2492 7 1 2 63260 64248
0 2493 5 1 1 2492
0 2494 7 1 2 2486 2493
0 2495 5 1 1 2494
0 2496 7 1 2 56799 2495
0 2497 5 1 1 2496
0 2498 7 3 2 48574 49283
0 2499 7 5 2 48311 59540
0 2500 7 1 2 64250 64253
0 2501 7 1 2 64249 2500
0 2502 5 1 1 2501
0 2503 7 1 2 2497 2502
0 2504 5 1 1 2503
0 2505 7 1 2 64116 2504
0 2506 5 1 1 2505
0 2507 7 4 2 48575 49156
0 2508 7 2 2 49518 56800
0 2509 5 1 1 64262
0 2510 7 1 2 64258 64263
0 2511 5 1 1 2510
0 2512 7 1 2 49284 63855
0 2513 5 1 1 2512
0 2514 7 1 2 2511 2513
0 2515 5 1 1 2514
0 2516 7 1 2 48312 2515
0 2517 5 1 1 2516
0 2518 7 8 2 48472 48576
0 2519 5 1 1 64264
0 2520 7 8 2 49403 49519
0 2521 5 3 1 64272
0 2522 7 12 2 64265 64273
0 2523 5 4 1 64283
0 2524 7 1 2 50614 58484
0 2525 5 3 1 2524
0 2526 7 1 2 64284 64299
0 2527 5 1 1 2526
0 2528 7 1 2 2517 2527
0 2529 5 1 1 2528
0 2530 7 1 2 54156 2529
0 2531 5 1 1 2530
0 2532 7 2 2 49285 64274
0 2533 7 4 2 48473 49157
0 2534 7 2 2 63376 64304
0 2535 7 1 2 64302 64308
0 2536 5 1 1 2535
0 2537 7 1 2 2531 2536
0 2538 5 1 1 2537
0 2539 7 1 2 53944 2538
0 2540 5 1 1 2539
0 2541 7 4 2 49286 49520
0 2542 5 1 1 64310
0 2543 7 7 2 64311 63377
0 2544 5 1 1 64314
0 2545 7 16 2 49404 54157
0 2546 5 1 1 64321
0 2547 7 3 2 48474 64322
0 2548 5 1 1 64337
0 2549 7 3 2 64315 64338
0 2550 5 1 1 64340
0 2551 7 1 2 2540 2550
0 2552 5 1 1 2551
0 2553 7 1 2 48064 2552
0 2554 5 1 1 2553
0 2555 7 11 2 48577 56801
0 2556 5 4 1 64343
0 2557 7 1 2 64190 64344
0 2558 5 1 1 2557
0 2559 7 1 2 2554 2558
0 2560 5 1 1 2559
0 2561 7 1 2 47771 2560
0 2562 5 1 1 2561
0 2563 7 2 2 56002 64212
0 2564 5 1 1 64358
0 2565 7 2 2 57569 2564
0 2566 5 1 1 64360
0 2567 7 6 2 49405 57858
0 2568 5 1 1 64362
0 2569 7 1 2 64363 63340
0 2570 7 1 2 2566 2569
0 2571 5 1 1 2570
0 2572 7 1 2 2562 2571
0 2573 5 1 1 2572
0 2574 7 1 2 63066 2573
0 2575 5 1 1 2574
0 2576 7 7 2 48847 62519
0 2577 5 17 1 64368
0 2578 7 2 2 63067 63299
0 2579 5 1 1 64392
0 2580 7 1 2 64375 2579
0 2581 5 3 1 2580
0 2582 7 1 2 61770 61295
0 2583 5 2 1 2582
0 2584 7 1 2 55168 64397
0 2585 5 1 1 2584
0 2586 7 2 2 58166 62787
0 2587 5 1 1 64399
0 2588 7 2 2 49158 60374
0 2589 5 2 1 64401
0 2590 7 1 2 64361 64403
0 2591 5 1 1 2590
0 2592 7 1 2 54468 59804
0 2593 7 1 2 2591 2592
0 2594 5 1 1 2593
0 2595 7 1 2 2587 2594
0 2596 5 1 1 2595
0 2597 7 1 2 48065 2596
0 2598 5 1 1 2597
0 2599 7 6 2 54469 57390
0 2600 5 2 1 64405
0 2601 7 1 2 52931 62741
0 2602 5 7 1 2601
0 2603 7 1 2 64406 64413
0 2604 5 2 1 2603
0 2605 7 1 2 2598 64420
0 2606 5 1 1 2605
0 2607 7 1 2 54830 2606
0 2608 5 1 1 2607
0 2609 7 1 2 2585 2608
0 2610 5 1 1 2609
0 2611 7 1 2 64394 2610
0 2612 5 1 1 2611
0 2613 7 3 2 49159 58653
0 2614 5 1 1 64422
0 2615 7 1 2 57090 64369
0 2616 5 1 1 2615
0 2617 7 2 2 63068 64285
0 2618 5 1 1 64425
0 2619 7 2 2 2616 2618
0 2620 5 1 1 64427
0 2621 7 5 2 48313 54831
0 2622 7 6 2 49287 55169
0 2623 7 2 2 64429 64434
0 2624 5 1 1 64440
0 2625 7 1 2 64441 63321
0 2626 5 1 1 2625
0 2627 7 1 2 64428 2626
0 2628 5 1 1 2627
0 2629 7 1 2 64423 2628
0 2630 5 1 1 2629
0 2631 7 1 2 63813 63069
0 2632 7 1 2 57091 2631
0 2633 5 1 1 2632
0 2634 7 14 2 54832 57859
0 2635 5 3 1 64442
0 2636 7 1 2 55170 64443
0 2637 7 1 2 63161 2636
0 2638 5 1 1 2637
0 2639 7 1 2 2633 2638
0 2640 5 1 1 2639
0 2641 7 1 2 56003 2640
0 2642 5 1 1 2641
0 2643 7 1 2 2630 2642
0 2644 5 1 1 2643
0 2645 7 1 2 62749 2644
0 2646 5 1 1 2645
0 2647 7 8 2 50615 57570
0 2648 5 9 1 64459
0 2649 7 7 2 64467 63136
0 2650 7 1 2 58239 64476
0 2651 5 1 1 2650
0 2652 7 1 2 50912 2651
0 2653 5 1 1 2652
0 2654 7 1 2 47772 2653
0 2655 5 1 1 2654
0 2656 7 1 2 61884 59293
0 2657 5 1 1 2656
0 2658 7 2 2 57126 62703
0 2659 5 6 1 64483
0 2660 7 1 2 50616 64485
0 2661 5 4 1 2660
0 2662 7 2 2 56004 64491
0 2663 5 1 1 64495
0 2664 7 1 2 60627 64496
0 2665 5 1 1 2664
0 2666 7 1 2 2657 2665
0 2667 7 1 2 2655 2666
0 2668 5 1 1 2667
0 2669 7 1 2 64370 2668
0 2670 5 1 1 2669
0 2671 7 16 2 47773 54833
0 2672 5 2 1 64497
0 2673 7 1 2 64213 64498
0 2674 5 1 1 2673
0 2675 7 1 2 58654 62797
0 2676 5 1 1 2675
0 2677 7 1 2 2674 2676
0 2678 5 1 1 2677
0 2679 7 1 2 48066 2678
0 2680 5 1 1 2679
0 2681 7 6 2 54834 56005
0 2682 5 4 1 64515
0 2683 7 1 2 61885 63963
0 2684 5 1 1 2683
0 2685 7 1 2 64521 2684
0 2686 5 1 1 2685
0 2687 7 1 2 49160 2686
0 2688 5 1 1 2687
0 2689 7 1 2 63464 2688
0 2690 7 1 2 2680 2689
0 2691 5 1 1 2690
0 2692 7 1 2 55171 63070
0 2693 7 1 2 2691 2692
0 2694 5 1 1 2693
0 2695 7 1 2 2670 2694
0 2696 5 1 1 2695
0 2697 7 1 2 57092 2696
0 2698 5 1 1 2697
0 2699 7 1 2 2646 2698
0 2700 7 1 2 2612 2699
0 2701 7 1 2 2575 2700
0 2702 7 2 2 55172 58639
0 2703 5 2 1 64525
0 2704 7 1 2 63024 64526
0 2705 5 1 1 2704
0 2706 7 1 2 57813 64395
0 2707 5 1 1 2706
0 2708 7 1 2 2705 2707
0 2709 5 1 1 2708
0 2710 7 1 2 54470 2709
0 2711 5 1 1 2710
0 2712 7 1 2 48848 59566
0 2713 7 1 2 61363 2712
0 2714 5 1 1 2713
0 2715 7 1 2 2711 2714
0 2716 5 1 1 2715
0 2717 7 1 2 54835 2716
0 2718 5 1 1 2717
0 2719 7 1 2 58199 2620
0 2720 5 1 1 2719
0 2721 7 1 2 2718 2720
0 2722 5 1 1 2721
0 2723 7 1 2 56006 2722
0 2724 5 1 1 2723
0 2725 7 3 2 64430 59608
0 2726 5 1 1 64529
0 2727 7 1 2 2726 58221
0 2728 5 1 1 2727
0 2729 7 1 2 63071 2728
0 2730 5 1 1 2729
0 2731 7 1 2 62520 64130
0 2732 7 1 2 64316 2731
0 2733 5 1 1 2732
0 2734 7 1 2 2730 2733
0 2735 5 1 1 2734
0 2736 7 1 2 55173 2735
0 2737 5 1 1 2736
0 2738 7 2 2 62521 57293
0 2739 5 1 1 64532
0 2740 7 1 2 48849 64533
0 2741 5 1 1 2740
0 2742 7 1 2 2737 2741
0 2743 5 1 1 2742
0 2744 7 1 2 47774 2743
0 2745 5 1 1 2744
0 2746 7 9 2 48067 57391
0 2747 5 3 1 64534
0 2748 7 2 2 58709 64543
0 2749 5 4 1 64546
0 2750 7 1 2 55174 64548
0 2751 7 1 2 63095 2750
0 2752 5 1 1 2751
0 2753 7 1 2 2745 2752
0 2754 5 1 1 2753
0 2755 7 1 2 56295 2754
0 2756 5 1 1 2755
0 2757 7 3 2 47775 63072
0 2758 7 1 2 64341 64552
0 2759 5 1 1 2758
0 2760 7 1 2 48068 64396
0 2761 5 1 1 2760
0 2762 7 2 2 57814 63162
0 2763 7 1 2 64444 64555
0 2764 5 1 1 2763
0 2765 7 4 2 48850 56507
0 2766 5 6 1 64557
0 2767 7 10 2 49521 49662
0 2768 5 4 1 64567
0 2769 7 1 2 64345 64568
0 2770 5 1 1 2769
0 2771 7 1 2 64561 2770
0 2772 5 1 1 2771
0 2773 7 1 2 57392 59574
0 2774 7 1 2 2772 2773
0 2775 5 1 1 2774
0 2776 7 1 2 2764 2775
0 2777 7 1 2 2761 2776
0 2778 5 1 1 2777
0 2779 7 1 2 55175 2778
0 2780 5 1 1 2779
0 2781 7 1 2 2759 2780
0 2782 7 20 2 54471 55176
0 2783 5 8 1 64581
0 2784 7 3 2 49663 64582
0 2785 5 1 1 64609
0 2786 7 5 2 48688 54158
0 2787 7 1 2 64610 64612
0 2788 5 1 1 2787
0 2789 7 6 2 55177 62883
0 2790 5 1 1 64617
0 2791 7 1 2 58200 64618
0 2792 5 1 1 2791
0 2793 7 1 2 54159 64371
0 2794 5 1 1 2793
0 2795 7 1 2 2792 2794
0 2796 5 1 1 2795
0 2797 7 1 2 47776 2796
0 2798 5 1 1 2797
0 2799 7 1 2 2788 2798
0 2800 5 1 1 2799
0 2801 7 1 2 57393 2800
0 2802 5 1 1 2801
0 2803 7 6 2 54160 63814
0 2804 7 1 2 64553 64623
0 2805 5 1 1 2804
0 2806 7 1 2 2802 2805
0 2807 5 1 1 2806
0 2808 7 1 2 57093 2807
0 2809 5 1 1 2808
0 2810 7 2 2 49406 61010
0 2811 5 1 1 64629
0 2812 7 1 2 55178 64630
0 2813 5 1 1 2812
0 2814 7 1 2 2091 2813
0 2815 5 2 1 2814
0 2816 7 1 2 48475 64631
0 2817 5 1 1 2816
0 2818 7 13 2 49407 54836
0 2819 5 1 1 64633
0 2820 7 2 2 49664 64634
0 2821 5 1 1 64646
0 2822 7 1 2 2817 2821
0 2823 5 1 1 2822
0 2824 7 1 2 48314 2823
0 2825 5 1 1 2824
0 2826 7 11 2 49288 54837
0 2827 5 1 1 64648
0 2828 7 1 2 64649 58910
0 2829 5 1 1 2828
0 2830 7 1 2 2825 2829
0 2831 5 1 1 2830
0 2832 7 1 2 62839 59567
0 2833 7 1 2 2831 2832
0 2834 5 1 1 2833
0 2835 7 1 2 2809 2834
0 2836 7 1 2 2781 2835
0 2837 7 1 2 2756 2836
0 2838 7 1 2 2724 2837
0 2839 5 1 1 2838
0 2840 7 1 2 61542 2839
0 2841 5 1 1 2840
0 2842 7 1 2 61740 64042
0 2843 5 1 1 2842
0 2844 7 6 2 49161 54838
0 2845 5 6 1 64659
0 2846 7 1 2 61886 64660
0 2847 5 2 1 2846
0 2848 7 1 2 2843 64671
0 2849 5 1 1 2848
0 2850 7 1 2 47777 2849
0 2851 5 1 1 2850
0 2852 7 1 2 57394 64499
0 2853 5 1 1 2852
0 2854 7 1 2 52473 64167
0 2855 5 2 1 2854
0 2856 7 1 2 56007 64414
0 2857 7 1 2 64673 2856
0 2858 5 1 1 2857
0 2859 7 1 2 2853 2858
0 2860 5 1 1 2859
0 2861 7 1 2 48069 2860
0 2862 5 1 1 2861
0 2863 7 2 2 56008 63433
0 2864 5 1 1 64675
0 2865 7 4 2 56508 57395
0 2866 5 1 1 64677
0 2867 7 1 2 2864 2866
0 2868 7 1 2 2862 2867
0 2869 7 1 2 2851 2868
0 2870 5 1 1 2869
0 2871 7 1 2 55179 2870
0 2872 5 1 1 2871
0 2873 7 1 2 53261 64665
0 2874 5 1 1 2873
0 2875 7 4 2 55180 56009
0 2876 5 4 1 64681
0 2877 7 2 2 63279 64251
0 2878 5 1 1 64689
0 2879 7 1 2 64685 2878
0 2880 5 1 1 2879
0 2881 7 1 2 62704 2880
0 2882 5 1 1 2881
0 2883 7 1 2 64601 2882
0 2884 5 1 1 2883
0 2885 7 1 2 2874 2884
0 2886 5 1 1 2885
0 2887 7 1 2 64445 61790
0 2888 5 1 1 2887
0 2889 7 4 2 48315 64312
0 2890 5 1 1 64691
0 2891 7 1 2 49162 64692
0 2892 5 1 1 2891
0 2893 7 1 2 51201 2892
0 2894 5 1 1 2893
0 2895 7 19 2 53945 54839
0 2896 5 2 1 64695
0 2897 7 3 2 47778 64696
0 2898 5 2 1 64716
0 2899 7 1 2 52474 64719
0 2900 5 1 1 2899
0 2901 7 1 2 54472 2900
0 2902 7 1 2 2894 2901
0 2903 5 1 1 2902
0 2904 7 1 2 2888 2903
0 2905 7 1 2 2886 2904
0 2906 5 1 1 2905
0 2907 7 1 2 48070 2906
0 2908 5 1 1 2907
0 2909 7 1 2 62705 64165
0 2910 7 1 2 64690 2909
0 2911 5 1 1 2910
0 2912 7 1 2 2908 2911
0 2913 7 1 2 2872 2912
0 2914 5 1 1 2913
0 2915 7 1 2 54161 2914
0 2916 5 1 1 2915
0 2917 7 4 2 55181 56509
0 2918 5 3 1 64721
0 2919 7 3 2 57396 61741
0 2920 5 3 1 64728
0 2921 7 1 2 61791 57729
0 2922 5 1 1 2921
0 2923 7 1 2 64731 2922
0 2924 5 1 1 2923
0 2925 7 1 2 64722 2924
0 2926 5 1 1 2925
0 2927 7 8 2 47779 57860
0 2928 5 2 1 64734
0 2929 7 1 2 64742 64602
0 2930 5 1 1 2929
0 2931 7 1 2 62798 2930
0 2932 5 1 1 2931
0 2933 7 3 2 48578 64232
0 2934 5 4 1 64744
0 2935 7 1 2 64415 64745
0 2936 5 1 1 2935
0 2937 7 10 2 55182 57397
0 2938 7 1 2 61801 64751
0 2939 5 1 1 2938
0 2940 7 1 2 64747 2939
0 2941 5 1 1 2940
0 2942 7 1 2 48071 2941
0 2943 5 1 1 2942
0 2944 7 1 2 2936 2943
0 2945 7 1 2 2932 2944
0 2946 5 1 1 2945
0 2947 7 1 2 54840 2946
0 2948 5 1 1 2947
0 2949 7 1 2 2926 2948
0 2950 7 1 2 2916 2949
0 2951 5 1 1 2950
0 2952 7 1 2 63073 2951
0 2953 5 1 1 2952
0 2954 7 1 2 56435 64666
0 2955 5 1 1 2954
0 2956 7 1 2 48851 2955
0 2957 5 1 1 2956
0 2958 7 5 2 48072 57861
0 2959 7 6 2 49163 64761
0 2960 7 1 2 64624 64766
0 2961 5 1 1 2960
0 2962 7 1 2 2957 2961
0 2963 5 1 1 2962
0 2964 7 1 2 56010 2963
0 2965 5 1 1 2964
0 2966 7 2 2 57862 64435
0 2967 5 1 1 64772
0 2968 7 1 2 64431 64773
0 2969 5 3 1 2968
0 2970 7 1 2 64562 64774
0 2971 5 1 1 2970
0 2972 7 1 2 57127 2971
0 2973 5 1 1 2972
0 2974 7 1 2 2965 2973
0 2975 5 1 1 2974
0 2976 7 1 2 53946 2975
0 2977 5 1 1 2976
0 2978 7 16 2 54162 55183
0 2979 5 2 1 64777
0 2980 7 3 2 48073 64778
0 2981 5 1 1 64795
0 2982 7 1 2 57863 64796
0 2983 5 1 1 2982
0 2984 7 1 2 52755 2983
0 2985 5 2 1 2984
0 2986 7 15 2 54841 57398
0 2987 5 1 1 64800
0 2988 7 1 2 64798 64801
0 2989 5 1 1 2988
0 2990 7 1 2 64558 58240
0 2991 5 1 1 2990
0 2992 7 1 2 2989 2991
0 2993 7 1 2 2977 2992
0 2994 5 1 1 2993
0 2995 7 1 2 47780 2994
0 2996 5 1 1 2995
0 2997 7 1 2 48852 62752
0 2998 5 1 1 2997
0 2999 7 8 2 49522 55184
0 3000 7 5 2 48579 64815
0 3001 5 4 1 64823
0 3002 7 1 2 62799 64824
0 3003 5 1 1 3002
0 3004 7 1 2 2998 3003
0 3005 5 1 1 3004
0 3006 7 1 2 54842 3005
0 3007 5 1 1 3006
0 3008 7 1 2 64446 64682
0 3009 5 2 1 3008
0 3010 7 3 2 48853 49289
0 3011 7 2 2 48316 64834
0 3012 5 1 1 64837
0 3013 7 3 2 57864 63815
0 3014 5 2 1 64839
0 3015 7 1 2 3012 64842
0 3016 5 3 1 3015
0 3017 7 2 2 62706 56683
0 3018 5 3 1 64847
0 3019 7 2 2 57203 64849
0 3020 5 5 1 64852
0 3021 7 1 2 64844 64854
0 3022 5 1 1 3021
0 3023 7 1 2 64832 3022
0 3024 5 1 1 3023
0 3025 7 1 2 54163 3024
0 3026 5 1 1 3025
0 3027 7 1 2 64563 3026
0 3028 7 1 2 3007 3027
0 3029 5 1 1 3028
0 3030 7 1 2 54473 3029
0 3031 5 1 1 3030
0 3032 7 5 2 48854 54843
0 3033 5 1 1 64859
0 3034 7 1 2 64860 62810
0 3035 5 1 1 3034
0 3036 7 1 2 3031 3035
0 3037 7 1 2 2996 3036
0 3038 5 1 1 3037
0 3039 7 1 2 62522 3038
0 3040 5 1 1 3039
0 3041 7 1 2 48855 61210
0 3042 7 1 2 59312 3041
0 3043 5 1 1 3042
0 3044 7 1 2 3040 3043
0 3045 7 1 2 2953 3044
0 3046 5 1 1 3045
0 3047 7 1 2 56296 3046
0 3048 5 1 1 3047
0 3049 7 1 2 2841 3048
0 3050 7 1 2 2701 3049
0 3051 7 1 2 2506 3050
0 3052 5 1 1 3051
0 3053 7 1 2 55734 3052
0 3054 5 1 1 3053
0 3055 7 1 2 62253 64714
0 3056 5 1 1 3055
0 3057 7 1 2 55185 3056
0 3058 5 1 1 3057
0 3059 7 11 2 48476 54164
0 3060 5 3 1 64864
0 3061 7 6 2 48317 62005
0 3062 7 4 2 64865 64878
0 3063 5 1 1 64884
0 3064 7 1 2 51202 3063
0 3065 5 3 1 3064
0 3066 7 1 2 47781 64888
0 3067 5 1 1 3066
0 3068 7 7 2 54165 58935
0 3069 5 1 1 64891
0 3070 7 1 2 64892 61887
0 3071 5 1 1 3070
0 3072 7 1 2 3067 3071
0 3073 5 1 1 3072
0 3074 7 1 2 54844 3073
0 3075 5 1 1 3074
0 3076 7 1 2 3058 3075
0 3077 5 1 1 3076
0 3078 7 1 2 48074 3077
0 3079 5 1 1 3078
0 3080 7 5 2 48477 64635
0 3081 5 7 1 64898
0 3082 7 2 2 60375 64899
0 3083 5 1 1 64910
0 3084 7 1 2 61712 64911
0 3085 5 1 1 3084
0 3086 7 1 2 61919 63972
0 3087 5 2 1 3086
0 3088 7 1 2 56297 64912
0 3089 5 1 1 3088
0 3090 7 9 2 47782 56802
0 3091 5 4 1 64914
0 3092 7 3 2 61011 62123
0 3093 5 3 1 64927
0 3094 7 2 2 64153 64930
0 3095 5 1 1 64933
0 3096 7 1 2 64923 64934
0 3097 7 1 2 3089 3096
0 3098 5 1 1 3097
0 3099 7 1 2 55186 3098
0 3100 5 1 1 3099
0 3101 7 1 2 3085 3100
0 3102 7 1 2 3079 3101
0 3103 5 1 1 3102
0 3104 7 1 2 58360 3103
0 3105 5 1 1 3104
0 3106 7 5 2 54845 60278
0 3107 5 2 1 64935
0 3108 7 6 2 63341 64879
0 3109 5 1 1 64942
0 3110 7 1 2 64936 64943
0 3111 5 1 1 3110
0 3112 7 4 2 48318 60054
0 3113 5 5 1 64948
0 3114 7 1 2 58710 64952
0 3115 5 4 1 3114
0 3116 7 1 2 56298 64957
0 3117 5 1 1 3116
0 3118 7 4 2 48478 62188
0 3119 5 3 1 64961
0 3120 7 3 2 58167 61012
0 3121 5 6 1 64968
0 3122 7 2 2 64965 64971
0 3123 5 1 1 64977
0 3124 7 1 2 3117 64978
0 3125 5 1 1 3124
0 3126 7 1 2 48075 3125
0 3127 5 1 1 3126
0 3128 7 1 2 2228 2246
0 3129 5 1 1 3128
0 3130 7 1 2 56299 3129
0 3131 5 1 1 3130
0 3132 7 1 2 50913 63908
0 3133 5 2 1 3132
0 3134 7 1 2 54474 64979
0 3135 5 1 1 3134
0 3136 7 1 2 56803 63882
0 3137 5 1 1 3136
0 3138 7 1 2 3135 3137
0 3139 7 1 2 3131 3138
0 3140 7 1 2 3127 3139
0 3141 5 1 1 3140
0 3142 7 1 2 55187 3141
0 3143 5 1 1 3142
0 3144 7 1 2 3111 3143
0 3145 7 1 2 3105 3144
0 3146 5 1 1 3145
0 3147 7 1 2 49164 3146
0 3148 5 1 1 3147
0 3149 7 5 2 47783 58655
0 3150 5 1 1 64981
0 3151 7 4 2 49096 60279
0 3152 5 1 1 64986
0 3153 7 4 2 53865 64987
0 3154 5 1 1 64990
0 3155 7 1 2 64982 64991
0 3156 5 1 1 3155
0 3157 7 2 2 64940 3156
0 3158 5 2 1 64994
0 3159 7 1 2 56976 64995
0 3160 5 1 1 3159
0 3161 7 1 2 49165 3160
0 3162 5 1 1 3161
0 3163 7 16 2 52065 50353
0 3164 5 7 1 64998
0 3165 7 2 2 56977 59482
0 3166 5 2 1 65021
0 3167 7 1 2 65014 65023
0 3168 5 1 1 3167
0 3169 7 7 2 58361 57815
0 3170 5 2 1 65025
0 3171 7 1 2 58640 65026
0 3172 5 2 1 3171
0 3173 7 1 2 65034 63465
0 3174 7 1 2 3168 3173
0 3175 7 1 2 3162 3174
0 3176 5 1 1 3175
0 3177 7 1 2 55188 3176
0 3178 5 1 1 3177
0 3179 7 3 2 64866 62135
0 3180 5 2 1 65036
0 3181 7 6 2 53866 54846
0 3182 5 2 1 65041
0 3183 7 3 2 59427 65042
0 3184 5 1 1 65049
0 3185 7 1 2 65037 65050
0 3186 5 1 1 3185
0 3187 7 9 2 48076 54847
0 3188 5 2 1 65052
0 3189 7 13 2 54475 56804
0 3190 5 4 1 65063
0 3191 7 1 2 65064 61086
0 3192 5 1 1 3191
0 3193 7 1 2 51203 3192
0 3194 5 1 1 3193
0 3195 7 1 2 65053 3194
0 3196 5 1 1 3195
0 3197 7 2 2 56300 411
0 3198 7 1 2 55189 65080
0 3199 5 1 1 3198
0 3200 7 1 2 3196 3199
0 3201 5 1 1 3200
0 3202 7 1 2 59965 3201
0 3203 5 1 1 3202
0 3204 7 1 2 3186 3203
0 3205 7 1 2 3178 3204
0 3206 5 1 1 3205
0 3207 7 1 2 56011 3206
0 3208 5 1 1 3207
0 3209 7 2 2 64535 59966
0 3210 7 2 2 64636 63342
0 3211 5 4 1 65084
0 3212 7 1 2 65082 65085
0 3213 5 1 1 3212
0 3214 7 1 2 60260 63756
0 3215 5 3 1 3214
0 3216 7 1 2 54848 65090
0 3217 5 1 1 3216
0 3218 7 7 2 48077 59967
0 3219 5 2 1 65093
0 3220 7 2 2 65094 61202
0 3221 5 1 1 65102
0 3222 7 1 2 3217 3221
0 3223 5 1 1 3222
0 3224 7 1 2 54476 3223
0 3225 5 1 1 3224
0 3226 7 3 2 50617 60331
0 3227 5 2 1 65104
0 3228 7 1 2 58936 65107
0 3229 5 1 1 3228
0 3230 7 4 2 54849 59208
0 3231 5 1 1 65109
0 3232 7 14 2 62006 58225
0 3233 5 5 1 65113
0 3234 7 1 2 3231 65127
0 3235 7 1 2 3229 3234
0 3236 7 1 2 3225 3235
0 3237 5 1 1 3236
0 3238 7 1 2 55190 3237
0 3239 5 1 1 3238
0 3240 7 1 2 3213 3239
0 3241 7 1 2 3208 3240
0 3242 7 1 2 3148 3241
0 3243 5 1 1 3242
0 3244 7 1 2 63074 3243
0 3245 5 1 1 3244
0 3246 7 1 2 48856 59209
0 3247 5 2 1 3246
0 3248 7 1 2 48857 56012
0 3249 5 1 1 3248
0 3250 7 5 2 48319 55191
0 3251 5 1 1 65134
0 3252 7 2 2 61402 65135
0 3253 7 1 2 64637 65139
0 3254 5 1 1 3253
0 3255 7 1 2 52756 3254
0 3256 5 3 1 3255
0 3257 7 8 2 53867 60906
0 3258 5 2 1 65144
0 3259 7 1 2 65141 65145
0 3260 5 1 1 3259
0 3261 7 1 2 3249 3260
0 3262 5 1 1 3261
0 3263 7 1 2 54166 3262
0 3264 5 1 1 3263
0 3265 7 1 2 65132 3264
0 3266 5 1 1 3265
0 3267 7 1 2 54477 3266
0 3268 5 1 1 3267
0 3269 7 2 2 56013 63266
0 3270 7 1 2 48858 65154
0 3271 5 1 1 3270
0 3272 7 1 2 3268 3271
0 3273 5 1 1 3272
0 3274 7 1 2 56684 3273
0 3275 5 1 1 3274
0 3276 7 7 2 54850 61888
0 3277 7 3 2 59494 65156
0 3278 7 6 2 49166 49408
0 3279 7 3 2 49097 65166
0 3280 7 1 2 65140 65172
0 3281 7 1 2 65163 3280
0 3282 5 1 1 3281
0 3283 7 1 2 52757 3282
0 3284 5 1 1 3283
0 3285 7 2 2 62317 59428
0 3286 5 1 1 65175
0 3287 7 2 2 59495 65176
0 3288 5 2 1 65177
0 3289 7 6 2 47784 63932
0 3290 5 3 1 65181
0 3291 7 1 2 62336 65187
0 3292 5 1 1 3291
0 3293 7 1 2 49167 3292
0 3294 5 1 1 3293
0 3295 7 2 2 53150 60409
0 3296 5 3 1 65190
0 3297 7 1 2 52369 65191
0 3298 7 1 2 3294 3297
0 3299 5 1 1 3298
0 3300 7 1 2 54478 3299
0 3301 5 1 1 3300
0 3302 7 1 2 65179 3301
0 3303 5 1 1 3302
0 3304 7 1 2 56014 3303
0 3305 5 1 1 3304
0 3306 7 3 2 50354 62337
0 3307 5 15 1 65195
0 3308 7 1 2 65198 61087
0 3309 5 2 1 3308
0 3310 7 1 2 63154 65213
0 3311 5 1 1 3310
0 3312 7 1 2 59210 3311
0 3313 5 1 1 3312
0 3314 7 9 2 53048 50618
0 3315 5 2 1 65215
0 3316 7 7 2 52225 65216
0 3317 5 5 1 65226
0 3318 7 2 2 64999 65227
0 3319 5 1 1 65238
0 3320 7 1 2 54851 3319
0 3321 5 1 1 3320
0 3322 7 14 2 53868 54479
0 3323 5 5 1 65240
0 3324 7 3 2 49098 65241
0 3325 7 1 2 64402 65259
0 3326 5 3 1 3325
0 3327 7 1 2 51204 65262
0 3328 7 1 2 53151 58711
0 3329 5 2 1 3328
0 3330 7 1 2 57399 65265
0 3331 5 1 1 3330
0 3332 7 2 2 48479 62037
0 3333 5 1 1 65267
0 3334 7 1 2 3331 3333
0 3335 7 1 2 3327 3334
0 3336 7 1 2 3321 3335
0 3337 7 1 2 3313 3336
0 3338 7 1 2 3305 3337
0 3339 5 1 1 3338
0 3340 7 1 2 3284 3339
0 3341 5 1 1 3340
0 3342 7 1 2 3275 3341
0 3343 5 1 1 3342
0 3344 7 1 2 62523 3343
0 3345 5 1 1 3344
0 3346 7 1 2 47785 61382
0 3347 5 1 1 3346
0 3348 7 5 2 49168 56301
0 3349 5 1 1 65269
0 3350 7 1 2 56015 65270
0 3351 5 1 1 3350
0 3352 7 1 2 3347 3351
0 3353 5 1 1 3352
0 3354 7 8 2 48859 49665
0 3355 5 1 1 65274
0 3356 7 1 2 48078 65275
0 3357 7 1 2 3353 3356
0 3358 5 1 1 3357
0 3359 7 1 2 3345 3358
0 3360 7 1 2 3245 3359
0 3361 5 1 1 3360
0 3362 7 1 2 56510 3361
0 3363 5 1 1 3362
0 3364 7 1 2 65196 65188
0 3365 5 2 1 3364
0 3366 7 1 2 49169 65282
0 3367 5 1 1 3366
0 3368 7 1 2 60332 3367
0 3369 5 2 1 3368
0 3370 7 1 2 54480 65284
0 3371 5 1 1 3370
0 3372 7 1 2 3371 65180
0 3373 5 1 1 3372
0 3374 7 1 2 64638 3373
0 3375 5 1 1 3374
0 3376 7 1 2 54481 65283
0 3377 5 1 1 3376
0 3378 7 3 2 58362 62318
0 3379 5 1 1 65286
0 3380 7 3 2 54167 65287
0 3381 5 1 1 65289
0 3382 7 1 2 3377 3381
0 3383 5 1 1 3382
0 3384 7 1 2 49170 3383
0 3385 5 1 1 3384
0 3386 7 8 2 53152 50137
0 3387 5 3 1 65292
0 3388 7 1 2 54482 65300
0 3389 5 3 1 3388
0 3390 7 1 2 52066 65303
0 3391 5 1 1 3390
0 3392 7 2 2 50138 61494
0 3393 5 1 1 65306
0 3394 7 1 2 3393 65266
0 3395 7 1 2 3391 3394
0 3396 5 1 1 3395
0 3397 7 1 2 3385 3396
0 3398 5 1 1 3397
0 3399 7 1 2 54852 3398
0 3400 5 1 1 3399
0 3401 7 1 2 65167 64996
0 3402 5 1 1 3401
0 3403 7 1 2 3400 3402
0 3404 5 1 1 3403
0 3405 7 1 2 48480 3404
0 3406 5 1 1 3405
0 3407 7 1 2 3375 3406
0 3408 5 1 1 3407
0 3409 7 1 2 56016 3408
0 3410 5 1 1 3409
0 3411 7 2 2 50619 59726
0 3412 5 2 1 65308
0 3413 7 1 2 56302 65310
0 3414 5 1 1 3413
0 3415 7 4 2 53869 58656
0 3416 5 1 1 65312
0 3417 7 1 2 59429 65313
0 3418 5 1 1 3417
0 3419 7 1 2 3414 3418
0 3420 5 1 1 3419
0 3421 7 1 2 57400 3420
0 3422 5 1 1 3421
0 3423 7 6 2 49409 63358
0 3424 5 2 1 65316
0 3425 7 1 2 56303 58657
0 3426 5 1 1 3425
0 3427 7 1 2 65322 3426
0 3428 5 3 1 3427
0 3429 7 1 2 61088 65324
0 3430 5 1 1 3429
0 3431 7 1 2 65076 3430
0 3432 7 1 2 3422 3431
0 3433 5 1 1 3432
0 3434 7 1 2 59968 3433
0 3435 5 1 1 3434
0 3436 7 1 2 57401 65081
0 3437 5 1 1 3436
0 3438 7 5 2 48481 49099
0 3439 7 2 2 62278 65327
0 3440 7 1 2 57763 65332
0 3441 5 1 1 3440
0 3442 7 1 2 3437 3441
0 3443 7 1 2 3435 3442
0 3444 5 1 1 3443
0 3445 7 1 2 54853 3444
0 3446 5 1 1 3445
0 3447 7 14 2 52932 50355
0 3448 5 7 1 65334
0 3449 7 4 2 52067 65335
0 3450 5 6 1 65355
0 3451 7 1 2 56805 65359
0 3452 5 3 1 3451
0 3453 7 1 2 65365 65035
0 3454 5 1 1 3453
0 3455 7 1 2 54854 3454
0 3456 5 1 1 3455
0 3457 7 3 2 50356 58419
0 3458 5 10 1 65368
0 3459 7 3 2 49171 65371
0 3460 5 2 1 65381
0 3461 7 1 2 56806 65382
0 3462 5 1 1 3461
0 3463 7 1 2 50914 3462
0 3464 5 1 1 3463
0 3465 7 1 2 48079 65027
0 3466 5 1 1 3465
0 3467 7 1 2 56176 3466
0 3468 5 1 1 3467
0 3469 7 1 2 65348 59892
0 3470 5 1 1 3469
0 3471 7 1 2 52068 3470
0 3472 5 1 1 3471
0 3473 7 1 2 57402 3472
0 3474 7 1 2 3468 3473
0 3475 7 1 2 3464 3474
0 3476 5 1 1 3475
0 3477 7 1 2 3456 3476
0 3478 5 1 1 3477
0 3479 7 1 2 54483 3478
0 3480 5 1 1 3479
0 3481 7 1 2 65038 65083
0 3482 5 1 1 3481
0 3483 7 1 2 3480 3482
0 3484 7 1 2 3446 3483
0 3485 7 1 2 3410 3484
0 3486 5 1 1 3485
0 3487 7 2 2 55192 3486
0 3488 5 1 1 65386
0 3489 7 1 2 50620 65032
0 3490 5 3 1 3489
0 3491 7 2 2 57403 60280
0 3492 5 3 1 65391
0 3493 7 2 2 58644 63271
0 3494 5 1 1 65396
0 3495 7 2 2 65393 65397
0 3496 5 1 1 65398
0 3497 7 1 2 65388 3496
0 3498 5 1 1 3497
0 3499 7 4 2 48080 58363
0 3500 5 3 1 65400
0 3501 7 1 2 65401 62775
0 3502 5 2 1 3501
0 3503 7 1 2 3498 65407
0 3504 5 1 1 3503
0 3505 7 1 2 49172 3504
0 3506 5 1 1 3505
0 3507 7 1 2 59969 62247
0 3508 5 1 1 3507
0 3509 7 1 2 58922 3508
0 3510 5 1 1 3509
0 3511 7 1 2 48081 3510
0 3512 5 1 1 3511
0 3513 7 1 2 65077 3069
0 3514 7 1 2 3512 3513
0 3515 7 1 2 3506 3514
0 3516 5 1 1 3515
0 3517 7 1 2 54855 3516
0 3518 5 1 1 3517
0 3519 7 2 2 58241 59970
0 3520 5 2 1 65409
0 3521 7 2 2 50621 65411
0 3522 5 1 1 65413
0 3523 7 1 2 60281 65383
0 3524 5 1 1 3523
0 3525 7 1 2 65414 3524
0 3526 5 1 1 3525
0 3527 7 1 2 56304 3526
0 3528 5 1 1 3527
0 3529 7 3 2 50357 65100
0 3530 5 3 1 65415
0 3531 7 2 2 59430 65242
0 3532 7 1 2 65418 65421
0 3533 5 1 1 3532
0 3534 7 1 2 56978 3533
0 3535 7 1 2 3528 3534
0 3536 5 1 1 3535
0 3537 7 1 2 54856 3536
0 3538 5 1 1 3537
0 3539 7 5 2 49173 61653
0 3540 5 3 1 65423
0 3541 7 4 2 49100 49410
0 3542 5 1 1 65431
0 3543 7 6 2 48482 65432
0 3544 5 1 1 65435
0 3545 7 2 2 65424 65436
0 3546 5 1 1 65441
0 3547 7 1 2 58242 65442
0 3548 5 1 1 3547
0 3549 7 5 2 52933 60183
0 3550 5 3 1 65443
0 3551 7 1 2 60113 65444
0 3552 5 5 1 3551
0 3553 7 1 2 55193 65451
0 3554 5 1 1 3553
0 3555 7 1 2 3548 3554
0 3556 7 1 2 3538 3555
0 3557 5 1 1 3556
0 3558 7 1 2 56017 3557
0 3559 5 1 1 3558
0 3560 7 2 2 49174 65199
0 3561 5 2 1 65456
0 3562 7 1 2 65114 65457
0 3563 5 1 1 3562
0 3564 7 2 2 49175 59971
0 3565 5 4 1 65460
0 3566 7 1 2 59555 65462
0 3567 5 1 1 3566
0 3568 7 1 2 54484 3567
0 3569 7 1 2 64893 3568
0 3570 5 1 1 3569
0 3571 7 1 2 3563 3570
0 3572 5 1 1 3571
0 3573 7 1 2 58364 3572
0 3574 5 1 1 3573
0 3575 7 1 2 51205 62146
0 3576 5 1 1 3575
0 3577 7 1 2 65285 3576
0 3578 5 1 1 3577
0 3579 7 1 2 65452 64944
0 3580 5 1 1 3579
0 3581 7 5 2 52370 50622
0 3582 5 1 1 65466
0 3583 7 10 2 53153 50915
0 3584 5 2 1 65471
0 3585 7 2 2 65467 65472
0 3586 7 1 2 57571 65483
0 3587 5 1 1 3586
0 3588 7 1 2 55194 3587
0 3589 5 1 1 3588
0 3590 7 1 2 3580 3589
0 3591 7 1 2 3578 3590
0 3592 7 1 2 3574 3591
0 3593 7 1 2 3559 3592
0 3594 7 2 2 3518 3593
0 3595 5 1 1 65485
0 3596 7 1 2 57865 3595
0 3597 5 1 1 3596
0 3598 7 1 2 3488 3597
0 3599 5 1 1 3598
0 3600 7 1 2 63075 3599
0 3601 5 1 1 3600
0 3602 7 2 2 54168 63300
0 3603 5 1 1 65487
0 3604 7 4 2 55195 56305
0 3605 5 3 1 65489
0 3606 7 1 2 47786 65490
0 3607 5 1 1 3606
0 3608 7 1 2 3603 3607
0 3609 5 1 1 3608
0 3610 7 1 2 54857 3609
0 3611 5 1 1 3610
0 3612 7 2 2 56807 64735
0 3613 5 2 1 65496
0 3614 7 1 2 3611 65498
0 3615 5 1 1 3614
0 3616 7 1 2 63076 3615
0 3617 5 1 1 3616
0 3618 7 2 2 54858 63107
0 3619 5 1 1 65500
0 3620 7 2 2 48860 49411
0 3621 5 1 1 65502
0 3622 7 1 2 64843 3621
0 3623 5 1 1 3622
0 3624 7 1 2 48483 3623
0 3625 5 1 1 3624
0 3626 7 1 2 63816 64364
0 3627 5 1 1 3626
0 3628 7 1 2 64564 3627
0 3629 7 1 2 3625 3628
0 3630 5 1 1 3629
0 3631 7 1 2 47787 3630
0 3632 5 1 1 3631
0 3633 7 1 2 3619 3632
0 3634 5 1 1 3633
0 3635 7 1 2 62524 3634
0 3636 5 1 1 3635
0 3637 7 1 2 3617 3636
0 3638 5 1 1 3637
0 3639 7 1 2 58201 3638
0 3640 5 1 1 3639
0 3641 7 6 2 54859 62525
0 3642 7 1 2 63108 61412
0 3643 7 1 2 65504 3642
0 3644 5 1 1 3643
0 3645 7 1 2 3640 3644
0 3646 5 1 1 3645
0 3647 7 1 2 56018 3646
0 3648 5 1 1 3647
0 3649 7 1 2 47788 64549
0 3650 5 1 1 3649
0 3651 7 1 2 1934 3650
0 3652 5 1 1 3651
0 3653 7 1 2 56511 3652
0 3654 5 1 1 3653
0 3655 7 1 2 64536 64131
0 3656 5 2 1 3655
0 3657 7 1 2 3654 65510
0 3658 5 1 1 3657
0 3659 7 1 2 56306 3658
0 3660 5 1 1 3659
0 3661 7 1 2 64154 64924
0 3662 5 3 1 3661
0 3663 7 1 2 56512 65512
0 3664 5 1 1 3663
0 3665 7 3 2 64639 64867
0 3666 5 7 1 65515
0 3667 7 1 2 64743 65518
0 3668 7 1 2 3664 3667
0 3669 5 1 1 3668
0 3670 7 1 2 48082 3669
0 3671 5 1 1 3670
0 3672 7 1 2 3660 3671
0 3673 5 1 1 3672
0 3674 7 1 2 55196 3673
0 3675 5 1 1 3674
0 3676 7 9 2 54860 56307
0 3677 5 2 1 65525
0 3678 7 1 2 65526 58346
0 3679 5 1 1 3678
0 3680 7 12 2 54169 56808
0 3681 7 1 2 65536 63243
0 3682 5 1 1 3681
0 3683 7 1 2 3679 3682
0 3684 5 1 1 3683
0 3685 7 1 2 49523 64252
0 3686 7 1 2 3684 3685
0 3687 5 1 1 3686
0 3688 7 1 2 49290 64583
0 3689 5 1 1 3688
0 3690 7 1 2 49524 64640
0 3691 5 1 1 3690
0 3692 7 1 2 3689 3691
0 3693 5 1 1 3692
0 3694 7 1 2 48580 3693
0 3695 5 1 1 3694
0 3696 7 1 2 61013 64816
0 3697 5 1 1 3696
0 3698 7 1 2 3695 3697
0 3699 5 1 1 3698
0 3700 7 1 2 58194 3699
0 3701 5 1 1 3700
0 3702 7 1 2 3687 3701
0 3703 7 1 2 3675 3702
0 3704 5 1 1 3703
0 3705 7 1 2 63077 3704
0 3706 5 1 1 3705
0 3707 7 3 2 54861 58937
0 3708 5 1 1 65548
0 3709 7 1 2 65549 64799
0 3710 5 1 1 3709
0 3711 7 4 2 48083 55197
0 3712 5 3 1 65551
0 3713 7 1 2 64650 64868
0 3714 5 1 1 3713
0 3715 7 1 2 65555 3714
0 3716 5 1 1 3715
0 3717 7 1 2 47789 3716
0 3718 5 1 1 3717
0 3719 7 1 2 58243 57720
0 3720 5 1 1 3719
0 3721 7 1 2 3718 3720
0 3722 5 1 1 3721
0 3723 7 1 2 48861 3722
0 3724 5 1 1 3723
0 3725 7 1 2 3710 3724
0 3726 5 1 1 3725
0 3727 7 1 2 62526 3726
0 3728 5 1 1 3727
0 3729 7 1 2 62007 64611
0 3730 5 1 1 3729
0 3731 7 1 2 3033 3730
0 3732 5 1 1 3731
0 3733 7 1 2 58186 62293
0 3734 5 1 1 3733
0 3735 7 1 2 58737 3734
0 3736 5 1 1 3735
0 3737 7 1 2 3732 3736
0 3738 5 1 1 3737
0 3739 7 1 2 62840 58511
0 3740 5 1 1 3739
0 3741 7 1 2 64565 3740
0 3742 5 1 1 3741
0 3743 7 1 2 3742 64632
0 3744 5 1 1 3743
0 3745 7 1 2 3738 3744
0 3746 7 1 2 3728 3745
0 3747 7 1 2 3706 3746
0 3748 7 1 2 3648 3747
0 3749 5 1 1 3748
0 3750 7 1 2 58420 61515
0 3751 5 5 1 3750
0 3752 7 1 2 3749 65558
0 3753 5 1 1 3752
0 3754 7 2 2 48484 65503
0 3755 5 2 1 65563
0 3756 7 1 2 64566 57204
0 3757 5 1 1 3756
0 3758 7 1 2 56513 65142
0 3759 5 1 1 3758
0 3760 7 1 2 3759 64775
0 3761 5 1 1 3760
0 3762 7 1 2 3757 3761
0 3763 5 1 1 3762
0 3764 7 1 2 65565 3763
0 3765 5 1 1 3764
0 3766 7 1 2 63900 3765
0 3767 5 1 1 3766
0 3768 7 1 2 48862 65110
0 3769 5 1 1 3768
0 3770 7 1 2 57128 64845
0 3771 5 1 1 3770
0 3772 7 1 2 3771 64833
0 3773 5 1 1 3772
0 3774 7 1 2 61158 3773
0 3775 5 1 1 3774
0 3776 7 1 2 3769 3775
0 3777 7 1 2 3767 3776
0 3778 5 1 1 3777
0 3779 7 1 2 62527 3778
0 3780 5 1 1 3779
0 3781 7 1 2 63845 2544
0 3782 5 2 1 3781
0 3783 7 1 2 57129 65567
0 3784 5 1 1 3783
0 3785 7 1 2 56019 63817
0 3786 5 1 1 3785
0 3787 7 1 2 3784 3786
0 3788 5 1 1 3787
0 3789 7 1 2 56308 3788
0 3790 5 1 1 3789
0 3791 7 2 2 64295 2624
0 3792 5 1 1 65569
0 3793 7 1 2 57130 3792
0 3794 5 1 1 3793
0 3795 7 5 2 49412 64266
0 3796 7 2 2 64033 65571
0 3797 5 1 1 65576
0 3798 7 1 2 3794 3797
0 3799 7 1 2 3790 3798
0 3800 5 1 1 3799
0 3801 7 1 2 47790 3800
0 3802 5 1 1 3801
0 3803 7 2 2 57866 65527
0 3804 5 2 1 65578
0 3805 7 7 2 48320 64651
0 3806 5 1 1 65582
0 3807 7 1 2 63301 65583
0 3808 5 1 1 3807
0 3809 7 1 2 65580 3808
0 3810 7 1 2 3802 3809
0 3811 5 1 1 3810
0 3812 7 1 2 63078 3811
0 3813 5 1 1 3812
0 3814 7 1 2 3780 3813
0 3815 5 1 1 3814
0 3816 7 1 2 54485 3815
0 3817 5 1 1 3816
0 3818 7 2 2 62528 58577
0 3819 5 1 1 65589
0 3820 7 1 2 64559 65590
0 3821 5 1 1 3820
0 3822 7 4 2 57973 58952
0 3823 5 4 1 65591
0 3824 7 1 2 47791 65595
0 3825 5 1 1 3824
0 3826 7 2 2 54862 57094
0 3827 5 2 1 65599
0 3828 7 3 2 47792 56514
0 3829 7 3 2 56309 57131
0 3830 5 1 1 65606
0 3831 7 1 2 65603 65607
0 3832 5 1 1 3831
0 3833 7 1 2 65601 3832
0 3834 5 1 1 3833
0 3835 7 1 2 56020 3834
0 3836 5 1 1 3835
0 3837 7 1 2 3825 3836
0 3838 5 1 1 3837
0 3839 7 1 2 63079 3838
0 3840 5 1 1 3839
0 3841 7 6 2 47793 48863
0 3842 5 1 1 65609
0 3843 7 1 2 54863 65577
0 3844 5 1 1 3843
0 3845 7 1 2 3842 3844
0 3846 5 1 1 3845
0 3847 7 1 2 62529 3846
0 3848 5 1 1 3847
0 3849 7 1 2 3840 3848
0 3850 5 1 1 3849
0 3851 7 1 2 55198 3850
0 3852 5 1 1 3851
0 3853 7 1 2 3821 3852
0 3854 7 1 2 3817 3853
0 3855 5 1 1 3854
0 3856 7 1 2 64049 3855
0 3857 5 1 1 3856
0 3858 7 18 2 48689 48864
0 3859 5 1 1 65615
0 3860 7 2 2 65115 60952
0 3861 5 1 1 65633
0 3862 7 1 2 53870 65634
0 3863 7 1 2 62841 3862
0 3864 5 1 1 3863
0 3865 7 1 2 3859 3864
0 3866 5 1 1 3865
0 3867 7 1 2 49666 3866
0 3868 5 1 1 3867
0 3869 7 1 2 51480 3868
0 3870 7 1 2 3857 3869
0 3871 7 1 2 3753 3870
0 3872 7 1 2 3601 3871
0 3873 7 1 2 3363 3872
0 3874 7 1 2 57974 65486
0 3875 5 1 1 3874
0 3876 7 1 2 48865 3875
0 3877 5 1 1 3876
0 3878 7 1 2 57867 65387
0 3879 5 1 1 3878
0 3880 7 1 2 3877 3879
0 3881 5 1 1 3880
0 3882 7 1 2 62530 3881
0 3883 5 1 1 3882
0 3884 7 3 2 56809 61014
0 3885 5 1 1 65635
0 3886 7 3 2 55199 65636
0 3887 5 1 1 65638
0 3888 7 1 2 57868 65639
0 3889 5 1 1 3888
0 3890 7 1 2 48866 65528
0 3891 5 1 1 3890
0 3892 7 2 2 3889 3891
0 3893 5 1 1 65641
0 3894 7 1 2 48321 3893
0 3895 5 1 1 3894
0 3896 7 2 2 49291 64861
0 3897 5 1 1 65643
0 3898 7 1 2 56310 65644
0 3899 5 1 1 3898
0 3900 7 1 2 3895 3899
0 3901 5 1 1 3900
0 3902 7 1 2 48084 3901
0 3903 5 1 1 3902
0 3904 7 1 2 65065 64825
0 3905 5 1 1 3904
0 3906 7 1 2 3897 3905
0 3907 5 1 1 3906
0 3908 7 1 2 48322 3907
0 3909 5 1 1 3908
0 3910 7 1 2 65642 3909
0 3911 5 1 1 3910
0 3912 7 1 2 47794 3911
0 3913 5 1 1 3912
0 3914 7 1 2 56311 64846
0 3915 5 1 1 3914
0 3916 7 1 2 65566 64776
0 3917 7 1 2 3915 3916
0 3918 5 1 1 3917
0 3919 7 1 2 54486 3918
0 3920 5 1 1 3919
0 3921 7 1 2 3913 3920
0 3922 5 1 1 3921
0 3923 7 1 2 48085 3922
0 3924 5 1 1 3923
0 3925 7 2 2 55200 58938
0 3926 5 1 1 65645
0 3927 7 1 2 57869 65646
0 3928 5 1 1 3927
0 3929 7 1 2 48867 63991
0 3930 5 1 1 3929
0 3931 7 1 2 3928 3930
0 3932 5 1 1 3931
0 3933 7 1 2 54864 3932
0 3934 5 1 1 3933
0 3935 7 4 2 48485 48868
0 3936 7 2 2 62025 65647
0 3937 5 1 1 65651
0 3938 7 1 2 3934 3937
0 3939 7 1 2 3924 3938
0 3940 5 1 1 3939
0 3941 7 1 2 54170 3940
0 3942 5 1 1 3941
0 3943 7 1 2 3903 3942
0 3944 5 1 1 3943
0 3945 7 1 2 53947 3944
0 3946 5 1 1 3945
0 3947 7 2 2 64817 64346
0 3948 5 1 1 65653
0 3949 7 1 2 48869 61015
0 3950 5 1 1 3949
0 3951 7 1 2 3948 3950
0 3952 5 1 1 3951
0 3953 7 1 2 48323 3952
0 3954 5 1 1 3953
0 3955 7 1 2 48870 62136
0 3956 5 1 1 3955
0 3957 7 1 2 48871 54487
0 3958 5 1 1 3957
0 3959 7 2 2 49413 64436
0 3960 5 1 1 65655
0 3961 7 1 2 57870 65656
0 3962 5 1 1 3961
0 3963 7 1 2 3958 3962
0 3964 5 1 1 3963
0 3965 7 1 2 48486 3964
0 3966 5 1 1 3965
0 3967 7 1 2 3956 3966
0 3968 7 1 2 3954 3967
0 3969 5 1 1 3968
0 3970 7 1 2 64500 3969
0 3971 5 1 1 3970
0 3972 7 1 2 3946 3971
0 3973 5 1 1 3972
0 3974 7 1 2 62531 3973
0 3975 5 1 1 3974
0 3976 7 1 2 56021 65579
0 3977 5 1 1 3976
0 3978 7 1 2 48324 65640
0 3979 5 1 1 3978
0 3980 7 1 2 3977 3979
0 3981 5 1 1 3980
0 3982 7 1 2 48086 3981
0 3983 5 1 1 3982
0 3984 7 1 2 56312 65568
0 3985 5 1 1 3984
0 3986 7 1 2 65570 3985
0 3987 5 1 1 3986
0 3988 7 1 2 54488 3987
0 3989 5 1 1 3988
0 3990 7 4 2 49414 55201
0 3991 5 1 1 65657
0 3992 7 1 2 63343 65658
0 3993 5 1 1 3992
0 3994 7 1 2 49292 64447
0 3995 5 1 1 3994
0 3996 7 1 2 3993 3995
0 3997 5 1 1 3996
0 3998 7 1 2 48325 3997
0 3999 5 1 1 3998
0 4000 7 1 2 65581 3887
0 4001 7 1 2 3999 4000
0 4002 5 1 1 4001
0 4003 7 1 2 47795 4002
0 4004 5 1 1 4003
0 4005 7 1 2 3989 4004
0 4006 5 1 1 4005
0 4007 7 1 2 48087 4006
0 4008 5 1 1 4007
0 4009 7 1 2 56022 64746
0 4010 5 1 1 4009
0 4011 7 1 2 3926 4010
0 4012 5 1 1 4011
0 4013 7 1 2 54865 4012
0 4014 5 1 1 4013
0 4015 7 4 2 64365 61946
0 4016 5 1 1 65661
0 4017 7 1 2 4014 4016
0 4018 7 1 2 4008 4017
0 4019 5 1 1 4018
0 4020 7 1 2 54171 4019
0 4021 5 1 1 4020
0 4022 7 1 2 3983 4021
0 4023 5 1 1 4022
0 4024 7 1 2 53948 4023
0 4025 5 1 1 4024
0 4026 7 1 2 51206 3885
0 4027 5 1 1 4026
0 4028 7 1 2 54866 4027
0 4029 5 1 1 4028
0 4030 7 2 2 64652 56810
0 4031 5 1 1 65665
0 4032 7 1 2 64603 4031
0 4033 5 1 1 4032
0 4034 7 8 2 53949 58244
0 4035 5 8 1 65667
0 4036 7 1 2 4033 65668
0 4037 5 1 1 4036
0 4038 7 1 2 4029 4037
0 4039 5 1 1 4038
0 4040 7 1 2 47796 4039
0 4041 5 1 1 4040
0 4042 7 1 2 64527 65086
0 4043 5 1 1 4042
0 4044 7 1 2 54172 4043
0 4045 5 1 1 4044
0 4046 7 4 2 48088 61016
0 4047 5 1 1 65683
0 4048 7 1 2 55202 65684
0 4049 5 1 1 4048
0 4050 7 1 2 4045 4049
0 4051 5 1 1 4050
0 4052 7 1 2 53950 4051
0 4053 5 1 1 4052
0 4054 7 1 2 4041 4053
0 4055 5 1 1 4054
0 4056 7 1 2 48326 4055
0 4057 5 1 1 4056
0 4058 7 1 2 64246 65637
0 4059 5 1 1 4058
0 4060 7 1 2 58245 61889
0 4061 5 4 1 4060
0 4062 7 1 2 50916 65687
0 4063 5 2 1 4062
0 4064 7 1 2 47797 65691
0 4065 5 1 1 4064
0 4066 7 1 2 56313 65669
0 4067 5 1 1 4066
0 4068 7 1 2 4065 4067
0 4069 5 1 1 4068
0 4070 7 1 2 49293 4069
0 4071 5 1 1 4070
0 4072 7 1 2 48089 59474
0 4073 5 1 1 4072
0 4074 7 1 2 64155 4073
0 4075 5 1 1 4074
0 4076 7 1 2 53951 4075
0 4077 5 1 1 4076
0 4078 7 1 2 4071 4077
0 4079 5 1 1 4078
0 4080 7 1 2 55203 4079
0 4081 5 1 1 4080
0 4082 7 1 2 4059 4081
0 4083 7 1 2 4057 4082
0 4084 5 1 1 4083
0 4085 7 1 2 56515 4084
0 4086 5 1 1 4085
0 4087 7 1 2 64748 3960
0 4088 5 1 1 4087
0 4089 7 1 2 48487 4088
0 4090 5 1 1 4089
0 4091 7 1 2 54489 64366
0 4092 5 1 1 4091
0 4093 7 14 2 55204 56811
0 4094 5 1 1 65693
0 4095 7 1 2 57871 61017
0 4096 5 1 1 4095
0 4097 7 1 2 4094 4096
0 4098 5 1 1 4097
0 4099 7 1 2 48327 4098
0 4100 5 1 1 4099
0 4101 7 1 2 4092 4100
0 4102 7 1 2 4090 4101
0 4103 5 1 1 4102
0 4104 7 1 2 64501 4103
0 4105 5 1 1 4104
0 4106 7 1 2 4086 4105
0 4107 7 1 2 4025 4106
0 4108 5 1 1 4107
0 4109 7 1 2 63080 4108
0 4110 5 1 1 4109
0 4111 7 1 2 65610 61427
0 4112 5 1 1 4111
0 4113 7 1 2 65143 58202
0 4114 5 1 1 4113
0 4115 7 1 2 65133 4114
0 4116 5 1 1 4115
0 4117 7 3 2 53952 62532
0 4118 7 1 2 54173 65707
0 4119 7 1 2 4116 4118
0 4120 5 1 1 4119
0 4121 7 1 2 4112 4120
0 4122 5 1 1 4121
0 4123 7 1 2 56516 4122
0 4124 5 1 1 4123
0 4125 7 1 2 4110 4124
0 4126 7 1 2 3975 4125
0 4127 5 1 1 4126
0 4128 7 1 2 58601 4127
0 4129 5 1 1 4128
0 4130 7 1 2 3883 4129
0 4131 7 1 2 3873 4130
0 4132 7 1 2 3054 4131
0 4133 5 1 1 4132
0 4134 7 1 2 49830 4133
0 4135 7 1 2 2433 4134
0 4136 5 1 1 4135
0 4137 7 36 2 53609 55433
0 4138 5 4 1 65710
0 4139 7 1 2 58658 63146
0 4140 5 1 1 4139
0 4141 7 1 2 60410 60009
0 4142 5 2 1 4141
0 4143 7 1 2 48090 65750
0 4144 5 1 1 4143
0 4145 7 1 2 59629 4144
0 4146 5 1 1 4145
0 4147 7 1 2 54490 4146
0 4148 5 2 1 4147
0 4149 7 2 2 54491 65200
0 4150 5 1 1 65754
0 4151 7 2 2 49294 60376
0 4152 5 3 1 65756
0 4153 7 1 2 48091 60900
0 4154 5 2 1 4153
0 4155 7 1 2 65758 65761
0 4156 5 1 1 4155
0 4157 7 1 2 47798 4156
0 4158 5 1 1 4157
0 4159 7 1 2 4150 4158
0 4160 5 2 1 4159
0 4161 7 1 2 48328 65763
0 4162 5 1 1 4161
0 4163 7 1 2 65752 4162
0 4164 5 1 1 4163
0 4165 7 1 2 61089 4164
0 4166 5 1 1 4165
0 4167 7 1 2 4140 4166
0 4168 5 1 1 4167
0 4169 7 1 2 57095 4168
0 4170 5 1 1 4169
0 4171 7 12 2 50623 60184
0 4172 7 1 2 60446 65765
0 4173 5 1 1 4172
0 4174 7 1 2 63302 4173
0 4175 5 1 1 4174
0 4176 7 1 2 4170 4175
0 4177 5 1 1 4176
0 4178 7 1 2 54867 4177
0 4179 5 1 1 4178
0 4180 7 2 2 59609 58281
0 4181 5 3 1 65777
0 4182 7 1 2 47799 58303
0 4183 5 7 1 4182
0 4184 7 1 2 58485 65782
0 4185 5 1 1 4184
0 4186 7 1 2 54492 4185
0 4187 5 1 1 4186
0 4188 7 1 2 65779 4187
0 4189 5 1 1 4188
0 4190 7 1 2 53953 4189
0 4191 5 1 1 4190
0 4192 7 1 2 49295 58659
0 4193 5 3 1 4192
0 4194 7 1 2 61920 58156
0 4195 5 1 1 4194
0 4196 7 1 2 47800 4195
0 4197 5 1 1 4196
0 4198 7 1 2 59668 61880
0 4199 5 1 1 4198
0 4200 7 1 2 59630 63987
0 4201 5 1 1 4200
0 4202 7 1 2 53954 4201
0 4203 5 1 1 4202
0 4204 7 1 2 4199 4203
0 4205 7 1 2 4197 4204
0 4206 5 1 1 4205
0 4207 7 1 2 48329 4206
0 4208 5 1 1 4207
0 4209 7 1 2 65789 4208
0 4210 7 1 2 4191 4209
0 4211 5 1 1 4210
0 4212 7 1 2 48092 4211
0 4213 5 1 1 4212
0 4214 7 2 2 59631 57751
0 4215 5 1 1 65792
0 4216 7 1 2 48330 4215
0 4217 5 1 1 4216
0 4218 7 4 2 54174 59972
0 4219 5 13 1 65794
0 4220 7 1 2 59342 65798
0 4221 5 1 1 4220
0 4222 7 1 2 54493 4221
0 4223 5 1 1 4222
0 4224 7 1 2 4217 4223
0 4225 5 2 1 4224
0 4226 7 1 2 61090 65811
0 4227 5 1 1 4226
0 4228 7 1 2 64296 64972
0 4229 7 1 2 4227 4228
0 4230 7 1 2 4213 4229
0 4231 5 1 1 4230
0 4232 7 1 2 63303 4231
0 4233 5 1 1 4232
0 4234 7 1 2 4179 4233
0 4235 5 1 1 4234
0 4236 7 1 2 55205 4235
0 4237 5 1 1 4236
0 4238 7 1 2 53049 58343
0 4239 5 7 1 4238
0 4240 7 1 2 64937 65813
0 4241 5 1 1 4240
0 4242 7 4 2 48093 62707
0 4243 5 7 1 65820
0 4244 7 3 2 65799 65824
0 4245 5 8 1 65831
0 4246 7 2 2 57404 65834
0 4247 7 1 2 54494 65842
0 4248 5 1 1 4247
0 4249 7 1 2 4241 4248
0 4250 5 1 1 4249
0 4251 7 1 2 58365 4250
0 4252 5 1 1 4251
0 4253 7 1 2 56023 64247
0 4254 5 1 1 4253
0 4255 7 1 2 4252 4254
0 4256 5 1 1 4255
0 4257 7 1 2 49176 4256
0 4258 5 1 1 4257
0 4259 7 3 2 47801 60377
0 4260 5 2 1 65844
0 4261 7 2 2 50624 65847
0 4262 5 6 1 65849
0 4263 7 1 2 56024 65851
0 4264 5 1 1 4263
0 4265 7 1 2 54175 64468
0 4266 5 2 1 4265
0 4267 7 1 2 65394 65857
0 4268 7 1 2 4264 4267
0 4269 5 1 1 4268
0 4270 7 1 2 54868 4269
0 4271 5 1 1 4270
0 4272 7 1 2 4258 4271
0 4273 5 1 1 4272
0 4274 7 1 2 56517 4273
0 4275 5 1 1 4274
0 4276 7 3 2 49101 59250
0 4277 7 1 2 65164 65859
0 4278 5 1 1 4277
0 4279 7 2 2 58366 65461
0 4280 5 3 1 65862
0 4281 7 2 2 50625 60411
0 4282 5 5 1 65867
0 4283 7 1 2 65864 65868
0 4284 5 1 1 4283
0 4285 7 1 2 48094 4284
0 4286 5 1 1 4285
0 4287 7 2 2 57572 59407
0 4288 5 1 1 65874
0 4289 7 1 2 64014 61070
0 4290 7 1 2 65875 4289
0 4291 7 1 2 4286 4290
0 4292 5 1 1 4291
0 4293 7 1 2 57872 4292
0 4294 5 1 1 4293
0 4295 7 1 2 4278 4294
0 4296 7 1 2 4275 4295
0 4297 5 1 1 4296
0 4298 7 1 2 55206 4297
0 4299 5 1 1 4298
0 4300 7 2 2 54176 59586
0 4301 5 3 1 65876
0 4302 7 2 2 57573 65878
0 4303 5 8 1 65881
0 4304 7 1 2 64992 65883
0 4305 5 1 1 4304
0 4306 7 1 2 63909 4305
0 4307 5 1 1 4306
0 4308 7 1 2 49177 4307
0 4309 5 1 1 4308
0 4310 7 8 2 49296 62124
0 4311 5 3 1 65891
0 4312 7 1 2 57816 65892
0 4313 5 1 1 4312
0 4314 7 1 2 4309 4313
0 4315 5 1 1 4314
0 4316 7 4 2 48581 54495
0 4317 5 1 1 65902
0 4318 7 1 2 64191 65903
0 4319 7 1 2 4315 4318
0 4320 5 1 1 4319
0 4321 7 1 2 4299 4320
0 4322 5 1 1 4321
0 4323 7 1 2 56314 4322
0 4324 5 1 1 4323
0 4325 7 8 2 53955 57764
0 4326 5 6 1 65906
0 4327 7 2 2 58203 65907
0 4328 5 1 1 65920
0 4329 7 2 2 59532 65921
0 4330 5 5 1 65922
0 4331 7 4 2 52226 60981
0 4332 5 4 1 65929
0 4333 7 1 2 48095 65933
0 4334 5 1 1 4333
0 4335 7 1 2 59516 4334
0 4336 5 1 1 4335
0 4337 7 1 2 53956 4336
0 4338 5 1 1 4337
0 4339 7 1 2 65146 58325
0 4340 5 1 1 4339
0 4341 7 1 2 4338 4340
0 4342 5 1 1 4341
0 4343 7 1 2 49297 4342
0 4344 5 1 1 4343
0 4345 7 1 2 58367 60026
0 4346 5 1 1 4345
0 4347 7 1 2 61921 4346
0 4348 5 1 1 4347
0 4349 7 1 2 54177 4348
0 4350 5 1 1 4349
0 4351 7 1 2 4344 4350
0 4352 5 1 1 4351
0 4353 7 1 2 49178 4352
0 4354 5 1 1 4353
0 4355 7 5 2 50358 59737
0 4356 5 3 1 65937
0 4357 7 2 2 54496 65942
0 4358 5 1 1 65945
0 4359 7 1 2 65762 4358
0 4360 5 1 1 4359
0 4361 7 1 2 48331 4360
0 4362 5 1 1 4361
0 4363 7 5 2 54497 60282
0 4364 5 1 1 65947
0 4365 7 2 2 62319 61388
0 4366 5 1 1 65952
0 4367 7 1 2 4364 4366
0 4368 5 1 1 4367
0 4369 7 1 2 58304 4368
0 4370 5 1 1 4369
0 4371 7 1 2 53050 62742
0 4372 5 1 1 4371
0 4373 7 1 2 58660 4372
0 4374 5 1 1 4373
0 4375 7 1 2 4370 4374
0 4376 7 1 2 4362 4375
0 4377 7 1 2 4354 4376
0 4378 5 1 1 4377
0 4379 7 1 2 54869 4378
0 4380 5 1 1 4379
0 4381 7 1 2 65924 4380
0 4382 5 1 1 4381
0 4383 7 1 2 64286 4382
0 4384 5 1 1 4383
0 4385 7 1 2 4324 4384
0 4386 7 1 2 4237 4385
0 4387 5 2 1 4386
0 4388 7 1 2 65711 65954
0 4389 5 1 1 4388
0 4390 7 44 2 55207 51481
0 4391 5 2 1 65956
0 4392 7 5 2 57873 65957
0 4393 5 5 1 66002
0 4394 7 3 2 48096 62038
0 4395 7 1 2 64105 66012
0 4396 5 1 1 4395
0 4397 7 1 2 49415 65948
0 4398 7 1 2 65884 4397
0 4399 5 1 1 4398
0 4400 7 1 2 4396 4399
0 4401 5 1 1 4400
0 4402 7 1 2 58368 4401
0 4403 5 1 1 4402
0 4404 7 2 2 63861 62026
0 4405 5 1 1 66015
0 4406 7 1 2 4403 4405
0 4407 5 1 1 4406
0 4408 7 1 2 49179 4407
0 4409 5 1 1 4408
0 4410 7 1 2 62027 63866
0 4411 5 1 1 4410
0 4412 7 1 2 4409 4411
0 4413 5 1 1 4412
0 4414 7 1 2 48488 4413
0 4415 5 1 1 4414
0 4416 7 2 2 58369 60084
0 4417 5 1 1 66017
0 4418 7 3 2 62208 66018
0 4419 7 1 2 64641 59973
0 4420 7 1 2 66019 4419
0 4421 5 1 1 4420
0 4422 7 1 2 4415 4421
0 4423 5 1 1 4422
0 4424 7 1 2 66003 4423
0 4425 5 1 1 4424
0 4426 7 13 2 52371 53051
0 4427 5 2 1 66022
0 4428 7 5 2 52227 53154
0 4429 5 1 1 66037
0 4430 7 14 2 66023 66038
0 4431 5 5 1 66042
0 4432 7 49 2 51207 55434
0 4433 5 7 1 66061
0 4434 7 2 2 63636 66062
0 4435 7 1 2 66056 66117
0 4436 5 1 1 4435
0 4437 7 6 2 54870 56518
0 4438 5 1 1 66119
0 4439 7 2 2 65201 66120
0 4440 5 1 1 66125
0 4441 7 1 2 3154 60412
0 4442 5 1 1 4441
0 4443 7 1 2 49180 4442
0 4444 5 2 1 4443
0 4445 7 2 2 65848 66127
0 4446 5 1 1 66129
0 4447 7 2 2 55208 4446
0 4448 5 1 1 66131
0 4449 7 1 2 4440 4448
0 4450 5 1 1 4449
0 4451 7 1 2 57405 4450
0 4452 5 1 1 4451
0 4453 7 1 2 64456 4452
0 4454 5 1 1 4453
0 4455 7 1 2 49416 4454
0 4456 5 1 1 4455
0 4457 7 1 2 54871 65015
0 4458 5 2 1 4457
0 4459 7 1 2 56436 66133
0 4460 5 1 1 4459
0 4461 7 1 2 55209 4460
0 4462 5 1 1 4461
0 4463 7 1 2 56519 65051
0 4464 7 1 2 65670 4463
0 4465 5 1 1 4464
0 4466 7 1 2 4462 4465
0 4467 7 1 2 4456 4466
0 4468 5 1 1 4467
0 4469 7 1 2 65268 4468
0 4470 5 1 1 4469
0 4471 7 2 2 62338 58293
0 4472 5 2 1 66135
0 4473 7 1 2 47802 66137
0 4474 5 2 1 4473
0 4475 7 1 2 64227 66139
0 4476 5 2 1 4475
0 4477 7 1 2 65529 66141
0 4478 5 1 1 4477
0 4479 7 1 2 59452 64085
0 4480 5 1 1 4479
0 4481 7 1 2 57360 4480
0 4482 5 1 1 4481
0 4483 7 1 2 60283 4482
0 4484 5 1 1 4483
0 4485 7 1 2 65602 57301
0 4486 7 1 2 4484 4485
0 4487 7 1 2 4478 4486
0 4488 5 1 1 4487
0 4489 7 1 2 55210 4488
0 4490 5 1 1 4489
0 4491 7 2 2 53957 59489
0 4492 5 1 1 66143
0 4493 7 1 2 48097 66144
0 4494 5 1 1 4493
0 4495 7 2 2 59408 4494
0 4496 5 1 1 66145
0 4497 7 1 2 61326 66146
0 4498 5 1 1 4497
0 4499 7 1 2 54872 63304
0 4500 7 1 2 4498 4499
0 4501 5 1 1 4500
0 4502 7 1 2 4490 4501
0 4503 5 1 1 4502
0 4504 7 1 2 56025 4503
0 4505 5 1 1 4504
0 4506 7 2 2 55211 65016
0 4507 5 1 1 66147
0 4508 7 3 2 59496 62189
0 4509 7 1 2 65860 66149
0 4510 5 1 1 4509
0 4511 7 1 2 4507 4510
0 4512 5 1 1 4511
0 4513 7 1 2 54873 4512
0 4514 5 1 1 4513
0 4515 7 1 2 59211 66132
0 4516 5 1 1 4515
0 4517 7 1 2 4514 4516
0 4518 5 1 1 4517
0 4519 7 1 2 56520 4518
0 4520 5 1 1 4519
0 4521 7 8 2 49102 54178
0 4522 5 2 1 66152
0 4523 7 2 2 65425 66153
0 4524 5 2 1 66162
0 4525 7 1 2 57975 59460
0 4526 7 1 2 66164 4525
0 4527 5 1 1 4526
0 4528 7 4 2 51208 57976
0 4529 5 3 1 66166
0 4530 7 1 2 65202 66170
0 4531 7 1 2 59212 4530
0 4532 7 1 2 4527 4531
0 4533 5 1 1 4532
0 4534 7 1 2 64323 64752
0 4535 5 1 1 4534
0 4536 7 5 2 48098 59431
0 4537 5 1 1 66173
0 4538 7 2 2 48582 63367
0 4539 7 1 2 60378 66178
0 4540 7 1 2 66174 4539
0 4541 5 1 1 4540
0 4542 7 1 2 4535 4541
0 4543 7 1 2 4533 4542
0 4544 5 1 1 4543
0 4545 7 1 2 54874 4544
0 4546 5 1 1 4545
0 4547 7 2 2 52475 65061
0 4548 7 1 2 53262 66180
0 4549 5 2 1 4548
0 4550 7 1 2 49417 64753
0 4551 7 1 2 66182 4550
0 4552 5 1 1 4551
0 4553 7 1 2 64828 4552
0 4554 7 1 2 4546 4553
0 4555 7 1 2 4520 4554
0 4556 7 1 2 4505 4555
0 4557 7 1 2 4470 4556
0 4558 5 1 1 4557
0 4559 7 1 2 51482 4558
0 4560 5 1 1 4559
0 4561 7 1 2 4436 4560
0 4562 5 1 1 4561
0 4563 7 1 2 54498 4562
0 4564 5 1 1 4563
0 4565 7 2 2 58157 61039
0 4566 5 2 1 66184
0 4567 7 1 2 47803 66186
0 4568 5 1 1 4567
0 4569 7 1 2 64026 4568
0 4570 5 1 1 4569
0 4571 7 1 2 53958 4570
0 4572 5 1 1 4571
0 4573 7 1 2 61114 4572
0 4574 5 1 1 4573
0 4575 7 1 2 56315 4574
0 4576 5 1 1 4575
0 4577 7 1 2 64966 3184
0 4578 5 1 1 4577
0 4579 7 1 2 47804 4578
0 4580 5 1 1 4579
0 4581 7 1 2 64697 59490
0 4582 5 1 1 4581
0 4583 7 1 2 56812 61782
0 4584 5 1 1 4583
0 4585 7 1 2 4582 4584
0 4586 7 1 2 4580 4585
0 4587 7 1 2 4576 4586
0 4588 5 1 1 4587
0 4589 7 1 2 48099 4588
0 4590 5 1 1 4589
0 4591 7 6 2 48100 56813
0 4592 5 2 1 66188
0 4593 7 4 2 50917 56979
0 4594 5 8 1 66196
0 4595 7 2 2 65271 60966
0 4596 5 1 1 66208
0 4597 7 1 2 66197 4596
0 4598 5 1 1 4597
0 4599 7 1 2 48332 4598
0 4600 5 1 1 4599
0 4601 7 1 2 66194 4600
0 4602 5 1 1 4601
0 4603 7 1 2 59669 4602
0 4604 5 1 1 4603
0 4605 7 1 2 64132 58305
0 4606 5 1 1 4605
0 4607 7 1 2 65534 4606
0 4608 7 1 2 59632 59461
0 4609 5 1 1 4608
0 4610 7 1 2 56814 4609
0 4611 5 1 1 4610
0 4612 7 1 2 1414 60010
0 4613 5 1 1 4612
0 4614 7 3 2 56316 57765
0 4615 5 1 1 66210
0 4616 7 1 2 58370 66211
0 4617 7 1 2 4613 4616
0 4618 5 1 1 4617
0 4619 7 1 2 4611 4618
0 4620 7 1 2 4607 4619
0 4621 7 1 2 4604 4620
0 4622 7 1 2 4590 4621
0 4623 5 1 1 4622
0 4624 7 1 2 65958 4623
0 4625 5 1 1 4624
0 4626 7 9 2 50918 66063
0 4627 7 1 2 58712 66213
0 4628 5 1 1 4627
0 4629 7 1 2 4625 4628
0 4630 5 1 1 4629
0 4631 7 1 2 56521 4630
0 4632 5 1 1 4631
0 4633 7 1 2 57874 65017
0 4634 5 1 1 4633
0 4635 7 3 2 49103 61742
0 4636 5 1 1 66222
0 4637 7 2 2 59708 66223
0 4638 5 2 1 66225
0 4639 7 1 2 52372 66227
0 4640 5 2 1 4639
0 4641 7 1 2 59670 66229
0 4642 5 1 1 4641
0 4643 7 1 2 59610 66138
0 4644 5 1 1 4643
0 4645 7 1 2 4642 4644
0 4646 5 1 1 4645
0 4647 7 1 2 49418 4646
0 4648 5 1 1 4647
0 4649 7 7 2 48489 53959
0 4650 5 2 1 66231
0 4651 7 2 2 48101 66232
0 4652 5 1 1 66240
0 4653 7 1 2 59401 66241
0 4654 5 1 1 4653
0 4655 7 1 2 4648 4654
0 4656 5 1 1 4655
0 4657 7 1 2 54875 4656
0 4658 5 1 1 4657
0 4659 7 1 2 4634 4658
0 4660 5 1 1 4659
0 4661 7 1 2 65959 4660
0 4662 5 1 1 4661
0 4663 7 17 2 53960 50626
0 4664 5 1 1 66242
0 4665 7 3 2 66214 66243
0 4666 5 1 1 66259
0 4667 7 1 2 54179 66260
0 4668 5 2 1 4667
0 4669 7 5 2 54876 65960
0 4670 7 1 2 62279 59346
0 4671 7 1 2 66264 4670
0 4672 5 1 1 4671
0 4673 7 1 2 66262 4672
0 4674 5 1 1 4673
0 4675 7 1 2 47805 4674
0 4676 5 1 1 4675
0 4677 7 15 2 50627 51209
0 4678 5 3 1 66269
0 4679 7 16 2 50919 55435
0 4680 7 13 2 66270 66287
0 4681 5 4 1 66303
0 4682 7 1 2 56177 66128
0 4683 5 1 1 4682
0 4684 7 1 2 66304 4683
0 4685 5 1 1 4684
0 4686 7 1 2 4676 4685
0 4687 7 1 2 4662 4686
0 4688 5 1 1 4687
0 4689 7 1 2 48333 4688
0 4690 5 1 1 4689
0 4691 7 1 2 60413 65865
0 4692 5 1 1 4691
0 4693 7 1 2 48102 4692
0 4694 5 1 1 4693
0 4695 7 1 2 59409 4694
0 4696 5 2 1 4695
0 4697 7 4 2 48490 54877
0 4698 7 1 2 66320 66322
0 4699 5 1 1 4698
0 4700 7 1 2 57977 4699
0 4701 5 1 1 4700
0 4702 7 1 2 65961 4701
0 4703 5 1 1 4702
0 4704 7 1 2 60456 66305
0 4705 5 1 1 4704
0 4706 7 1 2 4703 4705
0 4707 5 1 1 4706
0 4708 7 1 2 62039 4707
0 4709 5 1 1 4708
0 4710 7 5 2 48583 64170
0 4711 5 2 1 66326
0 4712 7 2 2 59497 64698
0 4713 5 1 1 66333
0 4714 7 1 2 65173 66334
0 4715 5 1 1 4714
0 4716 7 1 2 57978 4715
0 4717 5 1 1 4716
0 4718 7 1 2 48103 4717
0 4719 5 1 1 4718
0 4720 7 1 2 66331 4719
0 4721 5 1 1 4720
0 4722 7 1 2 65962 4721
0 4723 5 1 1 4722
0 4724 7 1 2 53155 66130
0 4725 5 1 1 4724
0 4726 7 1 2 66306 4725
0 4727 5 1 1 4726
0 4728 7 1 2 4723 4727
0 4729 5 1 1 4728
0 4730 7 1 2 49298 4729
0 4731 5 1 1 4730
0 4732 7 5 2 54180 61654
0 4733 7 2 2 63364 66335
0 4734 5 1 1 66340
0 4735 7 1 2 66265 66341
0 4736 5 1 1 4735
0 4737 7 1 2 66316 4736
0 4738 5 1 1 4737
0 4739 7 1 2 48104 4738
0 4740 5 1 1 4739
0 4741 7 3 2 64324 65963
0 4742 7 1 2 64653 66342
0 4743 5 1 1 4742
0 4744 7 10 2 53156 50359
0 4745 5 4 1 66345
0 4746 7 2 2 59738 66346
0 4747 5 1 1 66359
0 4748 7 1 2 66307 4747
0 4749 5 1 1 4748
0 4750 7 1 2 66007 4749
0 4751 7 1 2 4743 4750
0 4752 7 1 2 4740 4751
0 4753 5 1 1 4752
0 4754 7 1 2 48491 4753
0 4755 5 1 1 4754
0 4756 7 1 2 59402 66308
0 4757 5 1 1 4756
0 4758 7 1 2 53961 66004
0 4759 5 2 1 4758
0 4760 7 1 2 4757 66361
0 4761 5 1 1 4760
0 4762 7 1 2 48105 4761
0 4763 5 1 1 4762
0 4764 7 1 2 66008 66263
0 4765 5 1 1 4764
0 4766 7 1 2 61091 4765
0 4767 5 1 1 4766
0 4768 7 1 2 4763 4767
0 4769 5 1 1 4768
0 4770 7 1 2 47806 4769
0 4771 5 1 1 4770
0 4772 7 5 2 51483 57875
0 4773 7 1 2 50920 64228
0 4774 5 1 1 4773
0 4775 7 1 2 66363 4774
0 4776 5 1 1 4775
0 4777 7 1 2 65746 4776
0 4778 5 1 1 4777
0 4779 7 1 2 55212 4778
0 4780 5 1 1 4779
0 4781 7 1 2 4771 4780
0 4782 7 1 2 4755 4781
0 4783 7 1 2 4731 4782
0 4784 7 1 2 4709 4783
0 4785 7 1 2 4690 4784
0 4786 7 1 2 4632 4785
0 4787 7 1 2 4564 4786
0 4788 5 1 1 4787
0 4789 7 1 2 48690 4788
0 4790 5 1 1 4789
0 4791 7 1 2 4425 4790
0 4792 5 1 1 4791
0 4793 7 1 2 49667 4792
0 4794 5 1 1 4793
0 4795 7 1 2 4389 4794
0 4796 5 1 1 4795
0 4797 7 1 2 48872 4796
0 4798 5 1 1 4797
0 4799 7 13 2 49668 54499
0 4800 5 2 1 66368
0 4801 7 2 2 65964 66369
0 4802 5 1 1 66383
0 4803 7 3 2 64835 63352
0 4804 7 2 2 66384 66385
0 4805 5 1 1 66388
0 4806 7 12 2 48873 51484
0 4807 7 5 2 64619 66390
0 4808 5 1 1 66402
0 4809 7 21 2 55213 55436
0 4810 7 6 2 53610 66407
0 4811 5 8 1 66428
0 4812 7 10 2 51485 56815
0 4813 7 1 2 48874 66442
0 4814 5 2 1 4813
0 4815 7 1 2 66434 66452
0 4816 5 2 1 4815
0 4817 7 1 2 62884 66454
0 4818 5 1 1 4817
0 4819 7 26 2 53611 55214
0 4820 5 2 1 66456
0 4821 7 4 2 55437 66457
0 4822 7 1 2 48875 66484
0 4823 5 1 1 4822
0 4824 7 1 2 4818 4823
0 4825 5 1 1 4824
0 4826 7 1 2 63992 4825
0 4827 5 1 1 4826
0 4828 7 1 2 4808 4827
0 4829 5 1 1 4828
0 4830 7 1 2 54878 4829
0 4831 5 1 1 4830
0 4832 7 6 2 53612 63081
0 4833 7 8 2 55438 66488
0 4834 7 2 2 65116 66494
0 4835 5 1 1 66502
0 4836 7 1 2 55215 66503
0 4837 5 1 1 4836
0 4838 7 1 2 4831 4837
0 4839 5 1 1 4838
0 4840 7 1 2 48106 4839
0 4841 5 1 1 4840
0 4842 7 1 2 4805 4841
0 4843 5 1 1 4842
0 4844 7 1 2 49181 4843
0 4845 5 1 1 4844
0 4846 7 5 2 48691 54879
0 4847 5 4 1 66504
0 4848 7 10 2 54500 51486
0 4849 7 1 2 64836 66513
0 4850 7 2 2 66505 4849
0 4851 7 5 2 49419 49669
0 4852 7 2 2 58226 66525
0 4853 7 1 2 66523 66530
0 4854 5 1 1 4853
0 4855 7 1 2 4845 4854
0 4856 5 1 1 4855
0 4857 7 1 2 53962 4856
0 4858 5 1 1 4857
0 4859 7 6 2 55439 56816
0 4860 7 3 2 63818 66489
0 4861 7 1 2 66532 66538
0 4862 5 1 1 4861
0 4863 7 1 2 4858 4862
0 4864 5 1 1 4863
0 4865 7 1 2 47807 4864
0 4866 5 1 1 4865
0 4867 7 3 2 65276 65965
0 4868 7 2 2 48692 54501
0 4869 7 2 2 66541 66544
0 4870 5 1 1 66546
0 4871 7 1 2 54880 66547
0 4872 5 1 1 4871
0 4873 7 1 2 4866 4872
0 4874 5 1 1 4873
0 4875 7 1 2 56522 4874
0 4876 5 1 1 4875
0 4877 7 6 2 49525 53613
0 4878 7 2 2 48584 55440
0 4879 7 2 2 66548 66554
0 4880 5 2 1 66556
0 4881 7 3 2 63819 66557
0 4882 5 1 1 66560
0 4883 7 1 2 49420 61302
0 4884 5 1 1 4883
0 4885 7 1 2 61115 4884
0 4886 5 2 1 4885
0 4887 7 1 2 57132 66563
0 4888 5 1 1 4887
0 4889 7 1 2 58551 60628
0 4890 5 1 1 4889
0 4891 7 1 2 4888 4890
0 4892 5 1 1 4891
0 4893 7 1 2 53963 4892
0 4894 5 1 1 4893
0 4895 7 1 2 58552 60741
0 4896 5 1 1 4895
0 4897 7 1 2 4894 4896
0 4898 5 1 1 4897
0 4899 7 1 2 47808 4898
0 4900 5 1 1 4899
0 4901 7 1 2 64880 56685
0 4902 5 1 1 4901
0 4903 7 1 2 4900 4902
0 4904 5 1 1 4903
0 4905 7 1 2 48492 4904
0 4906 5 1 1 4905
0 4907 7 2 2 60055 64325
0 4908 7 5 2 63244 60347
0 4909 5 1 1 66567
0 4910 7 1 2 66565 66568
0 4911 5 1 1 4910
0 4912 7 1 2 4906 4911
0 4913 5 1 1 4912
0 4914 7 1 2 54502 4913
0 4915 5 1 1 4914
0 4916 7 2 2 63359 62209
0 4917 5 1 1 66572
0 4918 7 1 2 66566 66573
0 4919 5 1 1 4918
0 4920 7 1 2 4915 4919
0 4921 5 1 1 4920
0 4922 7 1 2 66561 4921
0 4923 5 1 1 4922
0 4924 7 13 2 53614 53964
0 4925 5 1 1 66574
0 4926 7 1 2 54881 66575
0 4927 5 1 1 4926
0 4928 7 1 2 50139 65877
0 4929 5 1 1 4928
0 4930 7 1 2 63194 4929
0 4931 5 2 1 4930
0 4932 7 28 2 50921 51210
0 4933 5 1 1 66589
0 4934 7 1 2 59475 66590
0 4935 7 1 2 66587 4934
0 4936 5 1 1 4935
0 4937 7 1 2 4927 4936
0 4938 5 1 1 4937
0 4939 7 1 2 59192 65879
0 4940 5 1 1 4939
0 4941 7 1 2 4938 4940
0 4942 5 1 1 4941
0 4943 7 3 2 49421 50360
0 4944 7 2 2 63344 66617
0 4945 7 1 2 66591 66620
0 4946 5 1 1 4945
0 4947 7 3 2 53615 63434
0 4948 5 3 1 66622
0 4949 7 9 2 50628 66592
0 4950 7 8 2 49422 58516
0 4951 5 29 1 66637
0 4952 7 1 2 66628 66638
0 4953 5 1 1 4952
0 4954 7 1 2 66625 4953
0 4955 5 1 1 4954
0 4956 7 1 2 63883 4955
0 4957 5 1 1 4956
0 4958 7 1 2 4946 4957
0 4959 7 1 2 4942 4958
0 4960 5 1 1 4959
0 4961 7 1 2 55441 4960
0 4962 5 1 1 4961
0 4963 7 2 2 57406 64915
0 4964 7 6 2 51487 63820
0 4965 7 1 2 63862 66676
0 4966 7 1 2 66674 4965
0 4967 5 1 1 4966
0 4968 7 1 2 4962 4967
0 4969 5 1 1 4968
0 4970 7 1 2 56686 4969
0 4971 5 1 1 4970
0 4972 7 4 2 49423 50922
0 4973 5 1 1 66682
0 4974 7 5 2 48493 50629
0 4975 5 1 1 66686
0 4976 7 3 2 66683 66687
0 4977 5 1 1 66691
0 4978 7 2 2 51211 66692
0 4979 5 1 1 66694
0 4980 7 1 2 59099 66695
0 4981 5 1 1 4980
0 4982 7 13 2 53965 56817
0 4983 7 5 2 51212 63637
0 4984 7 1 2 66696 66709
0 4985 5 1 1 4984
0 4986 7 3 2 50923 57205
0 4987 5 2 1 66714
0 4988 7 1 2 53616 62396
0 4989 7 1 2 66717 4988
0 4990 7 1 2 64980 4989
0 4991 5 1 1 4990
0 4992 7 1 2 4985 4991
0 4993 5 1 1 4992
0 4994 7 1 2 54503 4993
0 4995 5 1 1 4994
0 4996 7 1 2 4981 4995
0 4997 5 1 1 4996
0 4998 7 1 2 47809 4997
0 4999 5 1 1 4998
0 5000 7 6 2 50361 66593
0 5001 7 2 2 57407 66719
0 5002 5 1 1 66725
0 5003 7 1 2 53617 60997
0 5004 5 1 1 5003
0 5005 7 1 2 5002 5004
0 5006 5 1 1 5005
0 5007 7 1 2 57730 5006
0 5008 5 1 1 5007
0 5009 7 3 2 59368 66594
0 5010 7 1 2 59251 66727
0 5011 5 1 1 5010
0 5012 7 1 2 5008 5011
0 5013 5 1 1 5012
0 5014 7 1 2 53966 5013
0 5015 5 1 1 5014
0 5016 7 14 2 53618 54181
0 5017 5 1 1 66730
0 5018 7 1 2 57133 66720
0 5019 5 1 1 5018
0 5020 7 1 2 5017 5019
0 5021 5 1 1 5020
0 5022 7 4 2 54504 62708
0 5023 5 2 1 66744
0 5024 7 1 2 56026 66745
0 5025 7 1 2 5021 5024
0 5026 5 1 1 5025
0 5027 7 20 2 53619 54882
0 5028 7 1 2 50362 62389
0 5029 5 5 1 5028
0 5030 7 1 2 66750 66770
0 5031 5 1 1 5030
0 5032 7 1 2 5026 5031
0 5033 7 1 2 5015 5032
0 5034 5 1 1 5033
0 5035 7 1 2 56317 5034
0 5036 5 1 1 5035
0 5037 7 2 2 57134 66751
0 5038 5 1 1 66775
0 5039 7 5 2 66595 66244
0 5040 7 1 2 56818 66777
0 5041 5 1 1 5040
0 5042 7 1 2 5038 5041
0 5043 5 1 1 5042
0 5044 7 1 2 56027 5043
0 5045 5 1 1 5044
0 5046 7 5 2 57135 56819
0 5047 7 1 2 66778 66782
0 5048 5 1 1 5047
0 5049 7 1 2 64477 66752
0 5050 5 1 1 5049
0 5051 7 1 2 5048 5050
0 5052 7 1 2 5045 5051
0 5053 5 1 1 5052
0 5054 7 1 2 54182 5053
0 5055 5 1 1 5054
0 5056 7 1 2 57408 66776
0 5057 5 1 1 5056
0 5058 7 1 2 5055 5057
0 5059 7 1 2 5036 5058
0 5060 7 1 2 4999 5059
0 5061 5 1 1 5060
0 5062 7 1 2 55442 5061
0 5063 5 1 1 5062
0 5064 7 2 2 64869 65168
0 5065 7 2 2 61018 66787
0 5066 7 1 2 63245 66266
0 5067 7 1 2 66789 5066
0 5068 5 1 1 5067
0 5069 7 1 2 5063 5068
0 5070 7 1 2 4971 5069
0 5071 5 1 1 5070
0 5072 7 1 2 56523 5071
0 5073 5 1 1 5072
0 5074 7 2 2 57876 59369
0 5075 5 1 1 66791
0 5076 7 1 2 66596 66792
0 5077 5 2 1 5076
0 5078 7 7 2 51213 57877
0 5079 7 4 2 47810 50630
0 5080 7 3 2 50924 66802
0 5081 7 1 2 66795 66806
0 5082 5 2 1 5081
0 5083 7 11 2 53620 54505
0 5084 7 4 2 55216 66811
0 5085 5 1 1 66822
0 5086 7 1 2 66809 5085
0 5087 5 1 1 5086
0 5088 7 1 2 48107 5087
0 5089 5 1 1 5088
0 5090 7 1 2 66793 5089
0 5091 5 1 1 5090
0 5092 7 1 2 56028 5091
0 5093 5 1 1 5092
0 5094 7 1 2 57409 65325
0 5095 5 1 1 5094
0 5096 7 1 2 65039 5095
0 5097 5 1 1 5096
0 5098 7 1 2 54883 5097
0 5099 5 1 1 5098
0 5100 7 3 2 49299 63435
0 5101 7 1 2 63246 66826
0 5102 5 1 1 5101
0 5103 7 1 2 64793 5102
0 5104 5 2 1 5103
0 5105 7 1 2 56318 66829
0 5106 5 1 1 5105
0 5107 7 1 2 64437 58168
0 5108 5 2 1 5107
0 5109 7 1 2 63436 66189
0 5110 5 1 1 5109
0 5111 7 1 2 66831 5110
0 5112 7 1 2 5106 5111
0 5113 5 1 1 5112
0 5114 7 1 2 47811 5113
0 5115 5 1 1 5114
0 5116 7 1 2 5099 5115
0 5117 5 1 1 5116
0 5118 7 1 2 53621 5117
0 5119 5 1 1 5118
0 5120 7 1 2 5093 5119
0 5121 5 1 1 5120
0 5122 7 1 2 61543 5121
0 5123 5 1 1 5122
0 5124 7 1 2 57410 61802
0 5125 5 2 1 5124
0 5126 7 1 2 50925 66833
0 5127 5 1 1 5126
0 5128 7 1 2 65317 5127
0 5129 5 1 1 5128
0 5130 7 1 2 64686 5129
0 5131 5 1 1 5130
0 5132 7 1 2 54506 5131
0 5133 5 1 1 5132
0 5134 7 1 2 56029 64900
0 5135 5 1 1 5134
0 5136 7 1 2 64604 5135
0 5137 5 1 1 5136
0 5138 7 1 2 64855 5137
0 5139 5 1 1 5138
0 5140 7 3 2 64881 66323
0 5141 5 3 1 66835
0 5142 7 1 2 5139 66838
0 5143 7 1 2 5133 5142
0 5144 5 1 1 5143
0 5145 7 1 2 54183 5144
0 5146 5 1 1 5145
0 5147 7 4 2 47812 55217
0 5148 7 3 2 64537 61743
0 5149 5 1 1 66845
0 5150 7 1 2 50926 5149
0 5151 5 2 1 5150
0 5152 7 1 2 66841 66848
0 5153 5 1 1 5152
0 5154 7 4 2 48334 61744
0 5155 5 2 1 66850
0 5156 7 1 2 65666 66851
0 5157 5 1 1 5156
0 5158 7 1 2 5153 5157
0 5159 7 1 2 5146 5158
0 5160 5 1 1 5159
0 5161 7 1 2 53622 5160
0 5162 5 1 1 5161
0 5163 7 2 2 65552 64214
0 5164 5 1 1 66856
0 5165 7 6 2 48335 61019
0 5166 5 4 1 66858
0 5167 7 2 2 49182 64699
0 5168 7 3 2 66859 66868
0 5169 5 1 1 66870
0 5170 7 1 2 5164 5169
0 5171 5 1 1 5170
0 5172 7 1 2 47813 5171
0 5173 5 1 1 5172
0 5174 7 1 2 64605 5173
0 5175 5 1 1 5174
0 5176 7 1 2 53623 5175
0 5177 5 1 1 5176
0 5178 7 1 2 5177 66810
0 5179 5 1 1 5178
0 5180 7 1 2 56319 5179
0 5181 5 1 1 5180
0 5182 7 1 2 56320 64160
0 5183 5 1 1 5182
0 5184 7 1 2 51214 5183
0 5185 5 1 1 5184
0 5186 7 2 2 66812 5185
0 5187 5 1 1 66873
0 5188 7 4 2 59124 66796
0 5189 5 2 1 66875
0 5190 7 1 2 58246 66458
0 5191 5 1 1 5190
0 5192 7 1 2 66879 5191
0 5193 5 1 1 5192
0 5194 7 1 2 47814 5193
0 5195 5 1 1 5194
0 5196 7 1 2 5187 5195
0 5197 5 1 1 5196
0 5198 7 1 2 62800 5197
0 5199 5 1 1 5198
0 5200 7 1 2 58578 66459
0 5201 5 1 1 5200
0 5202 7 12 2 50363 51215
0 5203 5 3 1 66881
0 5204 7 8 2 48585 50927
0 5205 5 4 1 66896
0 5206 7 2 2 64233 66897
0 5207 7 1 2 66882 66908
0 5208 5 1 1 5207
0 5209 7 1 2 5201 5208
0 5210 5 1 1 5209
0 5211 7 1 2 62753 5210
0 5212 5 1 1 5211
0 5213 7 3 2 54184 64762
0 5214 7 1 2 66629 66910
0 5215 5 1 1 5214
0 5216 7 3 2 64916 63437
0 5217 5 1 1 66913
0 5218 7 1 2 53624 66914
0 5219 5 1 1 5218
0 5220 7 1 2 5215 5219
0 5221 5 1 1 5220
0 5222 7 1 2 61792 5221
0 5223 5 1 1 5222
0 5224 7 1 2 5212 5223
0 5225 7 1 2 5199 5224
0 5226 7 1 2 5181 5225
0 5227 7 1 2 5162 5226
0 5228 7 1 2 5123 5227
0 5229 5 1 1 5228
0 5230 7 1 2 55443 5229
0 5231 5 1 1 5230
0 5232 7 5 2 63821 66364
0 5233 5 1 1 66916
0 5234 7 1 2 54507 63220
0 5235 5 1 1 5234
0 5236 7 2 2 47815 64478
0 5237 5 1 1 66921
0 5238 7 1 2 54185 66922
0 5239 5 1 1 5238
0 5240 7 1 2 5235 5239
0 5241 5 1 1 5240
0 5242 7 1 2 56687 5241
0 5243 5 1 1 5242
0 5244 7 1 2 59100 65852
0 5245 5 2 1 5244
0 5246 7 2 2 56030 58661
0 5247 5 4 1 66925
0 5248 7 1 2 58247 63977
0 5249 5 2 1 5248
0 5250 7 1 2 66927 66931
0 5251 7 1 2 66923 5250
0 5252 7 1 2 5243 5251
0 5253 5 1 1 5252
0 5254 7 1 2 56321 5253
0 5255 5 1 1 5254
0 5256 7 3 2 47816 60742
0 5257 5 2 1 66933
0 5258 7 1 2 65850 66936
0 5259 5 1 1 5258
0 5260 7 1 2 56820 5259
0 5261 5 1 1 5260
0 5262 7 1 2 64928 66934
0 5263 5 1 1 5262
0 5264 7 2 2 57136 63280
0 5265 5 1 1 66938
0 5266 7 1 2 59611 66939
0 5267 5 2 1 5266
0 5268 7 1 2 5263 66940
0 5269 7 1 2 5261 5268
0 5270 7 1 2 5255 5269
0 5271 5 1 1 5270
0 5272 7 1 2 66917 5271
0 5273 5 1 1 5272
0 5274 7 1 2 5231 5273
0 5275 7 1 2 5073 5274
0 5276 5 1 1 5275
0 5277 7 1 2 48876 5276
0 5278 5 1 1 5277
0 5279 7 1 2 4923 5278
0 5280 5 1 1 5279
0 5281 7 1 2 62533 5280
0 5282 5 1 1 5281
0 5283 7 1 2 64779 66183
0 5284 5 1 1 5283
0 5285 7 1 2 64457 5284
0 5286 5 1 1 5285
0 5287 7 1 2 61803 5286
0 5288 5 1 1 5287
0 5289 7 1 2 56524 64797
0 5290 7 1 2 64416 5289
0 5291 5 1 1 5290
0 5292 7 1 2 5288 5291
0 5293 5 1 1 5292
0 5294 7 1 2 57411 5293
0 5295 5 1 1 5294
0 5296 7 1 2 64829 5295
0 5297 5 1 1 5296
0 5298 7 1 2 54508 5297
0 5299 5 1 1 5298
0 5300 7 1 2 64736 66857
0 5301 5 1 1 5300
0 5302 7 1 2 5299 5301
0 5303 5 1 1 5302
0 5304 7 1 2 66490 5303
0 5305 5 1 1 5304
0 5306 7 2 2 47817 65616
0 5307 7 2 2 62675 66271
0 5308 5 1 1 66944
0 5309 7 1 2 66942 66945
0 5310 5 1 1 5309
0 5311 7 1 2 5305 5310
0 5312 5 1 1 5311
0 5313 7 1 2 55444 5312
0 5314 5 1 1 5313
0 5315 7 1 2 48108 64030
0 5316 5 2 1 5315
0 5317 7 1 2 2614 66946
0 5318 5 1 1 5317
0 5319 7 1 2 55218 5318
0 5320 5 1 1 5319
0 5321 7 1 2 64749 5320
0 5322 5 1 1 5321
0 5323 7 1 2 64502 5322
0 5324 5 1 1 5323
0 5325 7 1 2 56031 66935
0 5326 5 1 1 5325
0 5327 7 1 2 64027 5326
0 5328 5 1 1 5327
0 5329 7 1 2 55219 5328
0 5330 5 1 1 5329
0 5331 7 2 2 57137 57817
0 5332 5 1 1 66948
0 5333 7 2 2 64654 63281
0 5334 7 1 2 66949 66950
0 5335 5 1 1 5334
0 5336 7 1 2 5330 5335
0 5337 5 1 1 5336
0 5338 7 1 2 56525 5337
0 5339 5 1 1 5338
0 5340 7 1 2 5324 5339
0 5341 5 1 1 5340
0 5342 7 1 2 53967 5341
0 5343 5 1 1 5342
0 5344 7 1 2 56526 59101
0 5345 5 1 1 5344
0 5346 7 1 2 62397 63438
0 5347 5 1 1 5346
0 5348 7 1 2 58222 5347
0 5349 7 1 2 5345 5348
0 5350 5 1 1 5349
0 5351 7 1 2 64780 5350
0 5352 5 1 1 5351
0 5353 7 1 2 5343 5352
0 5354 5 1 1 5353
0 5355 7 1 2 48693 5354
0 5356 5 1 1 5355
0 5357 7 1 2 53968 59541
0 5358 7 2 2 64023 5357
0 5359 5 1 1 66952
0 5360 7 1 2 64840 66953
0 5361 5 1 1 5360
0 5362 7 1 2 5356 5361
0 5363 5 1 1 5362
0 5364 7 14 2 49670 51488
0 5365 5 2 1 66954
0 5366 7 1 2 48877 66955
0 5367 7 1 2 5363 5366
0 5368 5 1 1 5367
0 5369 7 1 2 5314 5368
0 5370 5 1 1 5369
0 5371 7 1 2 56322 5370
0 5372 5 1 1 5371
0 5373 7 8 2 49424 58505
0 5374 7 1 2 65712 66970
0 5375 5 1 1 5374
0 5376 7 10 2 48694 66956
0 5377 5 1 1 66978
0 5378 7 1 2 54509 66979
0 5379 5 1 1 5378
0 5380 7 1 2 5375 5379
0 5381 5 1 1 5380
0 5382 7 1 2 56527 5381
0 5383 5 1 1 5382
0 5384 7 1 2 64737 65713
0 5385 5 1 1 5384
0 5386 7 6 2 51489 58089
0 5387 7 1 2 56821 66370
0 5388 7 1 2 66988 5387
0 5389 5 1 1 5388
0 5390 7 1 2 5385 5389
0 5391 7 1 2 5383 5390
0 5392 5 1 1 5391
0 5393 7 1 2 48878 5392
0 5394 5 1 1 5393
0 5395 7 2 2 63305 65714
0 5396 5 1 1 66994
0 5397 7 7 2 47818 48695
0 5398 5 1 1 66996
0 5399 7 2 2 49671 66997
0 5400 7 1 2 66995 67003
0 5401 5 1 1 5400
0 5402 7 1 2 5394 5401
0 5403 5 1 1 5402
0 5404 7 1 2 58248 5403
0 5405 5 1 1 5404
0 5406 7 14 2 54510 55445
0 5407 7 3 2 53625 67005
0 5408 7 1 2 64393 67019
0 5409 5 1 1 5408
0 5410 7 1 2 5405 5409
0 5411 5 1 1 5410
0 5412 7 1 2 55220 5411
0 5413 5 1 1 5412
0 5414 7 3 2 62885 65611
0 5415 7 1 2 66309 67022
0 5416 5 1 1 5415
0 5417 7 9 2 49672 65617
0 5418 7 1 2 66514 67025
0 5419 5 2 1 5418
0 5420 7 5 2 48109 48879
0 5421 7 2 2 66980 67036
0 5422 5 1 1 67041
0 5423 7 1 2 54186 67042
0 5424 5 1 1 5423
0 5425 7 1 2 56528 66495
0 5426 5 1 1 5425
0 5427 7 1 2 5424 5426
0 5428 5 2 1 5427
0 5429 7 1 2 47819 67043
0 5430 5 1 1 5429
0 5431 7 1 2 67034 5430
0 5432 5 1 1 5431
0 5433 7 1 2 55221 5432
0 5434 5 1 1 5433
0 5435 7 6 2 53626 58662
0 5436 7 2 2 55446 67045
0 5437 5 1 1 67051
0 5438 7 1 2 63082 64763
0 5439 7 1 2 67052 5438
0 5440 5 1 1 5439
0 5441 7 1 2 5434 5440
0 5442 5 1 1 5441
0 5443 7 1 2 65530 5442
0 5444 5 1 1 5443
0 5445 7 1 2 5416 5444
0 5446 7 1 2 5413 5445
0 5447 5 1 1 5446
0 5448 7 1 2 62801 5447
0 5449 5 1 1 5448
0 5450 7 5 2 54884 56822
0 5451 7 4 2 55447 63083
0 5452 7 7 2 48586 66549
0 5453 7 1 2 64729 67062
0 5454 7 1 2 67058 5453
0 5455 5 1 1 5454
0 5456 7 1 2 4870 5455
0 5457 5 1 1 5456
0 5458 7 1 2 67053 5457
0 5459 5 1 1 5458
0 5460 7 3 2 48110 65715
0 5461 5 1 1 67069
0 5462 7 1 2 64133 67070
0 5463 5 1 1 5462
0 5464 7 2 2 47820 66391
0 5465 5 1 1 67072
0 5466 7 1 2 54511 67073
0 5467 5 1 1 5466
0 5468 7 1 2 5463 5467
0 5469 5 1 1 5468
0 5470 7 1 2 56323 5469
0 5471 5 1 1 5470
0 5472 7 2 2 64134 65716
0 5473 7 3 2 47821 58204
0 5474 5 2 1 67076
0 5475 7 1 2 67074 67077
0 5476 5 1 1 5475
0 5477 7 1 2 5476 66453
0 5478 7 1 2 5471 5477
0 5479 5 1 1 5478
0 5480 7 1 2 55222 5479
0 5481 5 1 1 5480
0 5482 7 2 2 64503 66515
0 5483 7 1 2 63109 66190
0 5484 7 1 2 67081 5483
0 5485 5 1 1 5484
0 5486 7 1 2 5481 5485
0 5487 5 1 1 5486
0 5488 7 1 2 56529 5487
0 5489 5 1 1 5488
0 5490 7 4 2 54885 57731
0 5491 7 2 2 66533 66460
0 5492 5 1 1 67087
0 5493 7 1 2 57878 66392
0 5494 5 1 1 5493
0 5495 7 1 2 5492 5494
0 5496 5 1 1 5495
0 5497 7 1 2 58249 5496
0 5498 5 1 1 5497
0 5499 7 4 2 55448 66550
0 5500 7 1 2 64347 67089
0 5501 5 1 1 5500
0 5502 7 1 2 5498 5501
0 5503 5 1 1 5502
0 5504 7 1 2 67083 5503
0 5505 5 1 1 5504
0 5506 7 6 2 50928 59370
0 5507 7 3 2 48111 66064
0 5508 5 1 1 67099
0 5509 7 1 2 67093 67100
0 5510 5 1 1 5509
0 5511 7 1 2 66009 5510
0 5512 5 1 1 5511
0 5513 7 1 2 48880 5512
0 5514 5 1 1 5513
0 5515 7 1 2 5505 5514
0 5516 7 1 2 5489 5515
0 5517 5 1 1 5516
0 5518 7 1 2 62886 5517
0 5519 5 1 1 5518
0 5520 7 1 2 57979 2981
0 5521 5 1 1 5520
0 5522 7 1 2 48881 67006
0 5523 7 1 2 66753 5522
0 5524 7 1 2 64917 5523
0 5525 7 1 2 5521 5524
0 5526 5 1 1 5525
0 5527 7 3 2 48112 57294
0 5528 5 1 1 67102
0 5529 7 1 2 56178 57752
0 5530 5 2 1 5529
0 5531 7 5 2 55449 63822
0 5532 7 18 2 48882 53627
0 5533 5 8 1 67112
0 5534 7 1 2 67107 67113
0 5535 7 1 2 67105 5534
0 5536 7 1 2 67103 5535
0 5537 5 1 1 5536
0 5538 7 1 2 5526 5537
0 5539 7 1 2 5519 5538
0 5540 5 1 1 5539
0 5541 7 1 2 61793 5540
0 5542 5 1 1 5541
0 5543 7 1 2 5459 5542
0 5544 7 1 2 5449 5543
0 5545 7 4 2 55223 66393
0 5546 5 1 1 67138
0 5547 7 2 2 57412 65717
0 5548 5 1 1 67142
0 5549 7 1 2 64192 67143
0 5550 5 1 1 5549
0 5551 7 1 2 5546 5550
0 5552 5 1 1 5551
0 5553 7 1 2 59575 5552
0 5554 5 1 1 5553
0 5555 7 3 2 55450 66731
0 5556 7 2 2 47822 49526
0 5557 7 1 2 67144 67147
0 5558 5 1 1 5557
0 5559 7 4 2 51490 57413
0 5560 7 1 2 67149 67037
0 5561 5 1 1 5560
0 5562 7 1 2 5558 5561
0 5563 5 1 1 5562
0 5564 7 1 2 55224 5563
0 5565 5 1 1 5564
0 5566 7 1 2 5554 5565
0 5567 5 1 1 5566
0 5568 7 1 2 62887 5567
0 5569 5 1 1 5568
0 5570 7 1 2 47823 66830
0 5571 5 1 1 5570
0 5572 7 3 2 58663 64802
0 5573 5 2 1 67153
0 5574 7 1 2 5571 67156
0 5575 5 1 1 5574
0 5576 7 1 2 48883 67090
0 5577 7 1 2 5575 5576
0 5578 5 1 1 5577
0 5579 7 1 2 5569 5578
0 5580 5 1 1 5579
0 5581 7 1 2 48587 5580
0 5582 5 1 1 5581
0 5583 7 1 2 64547 67079
0 5584 5 1 1 5583
0 5585 7 1 2 49527 5584
0 5586 5 1 1 5585
0 5587 7 1 2 64504 61267
0 5588 5 1 1 5587
0 5589 7 1 2 5586 5588
0 5590 5 1 1 5589
0 5591 7 1 2 66403 5590
0 5592 5 1 1 5591
0 5593 7 1 2 5582 5592
0 5594 5 1 1 5593
0 5595 7 1 2 56324 5594
0 5596 5 1 1 5595
0 5597 7 1 2 57371 66539
0 5598 5 1 1 5597
0 5599 7 7 2 48696 65277
0 5600 5 2 1 67158
0 5601 7 1 2 67159 66630
0 5602 5 1 1 5601
0 5603 7 1 2 5598 5602
0 5604 5 2 1 5603
0 5605 7 1 2 59568 67167
0 5606 5 1 1 5605
0 5607 7 1 2 48113 63306
0 5608 5 2 1 5607
0 5609 7 1 2 54886 61037
0 5610 5 1 1 5609
0 5611 7 1 2 67169 5610
0 5612 5 1 1 5611
0 5613 7 1 2 64584 66491
0 5614 7 1 2 5612 5613
0 5615 5 1 1 5614
0 5616 7 1 2 5606 5615
0 5617 5 1 1 5616
0 5618 7 1 2 55451 5617
0 5619 5 1 1 5618
0 5620 7 1 2 47824 65488
0 5621 5 1 1 5620
0 5622 7 1 2 64528 5621
0 5623 5 1 1 5622
0 5624 7 21 2 54887 51491
0 5625 7 2 2 67171 66371
0 5626 5 2 1 67192
0 5627 7 1 2 65618 67193
0 5628 7 1 2 5623 5627
0 5629 5 1 1 5628
0 5630 7 1 2 5619 5629
0 5631 5 1 1 5630
0 5632 7 1 2 56032 5631
0 5633 5 1 1 5632
0 5634 7 1 2 64234 65054
0 5635 5 1 1 5634
0 5636 7 1 2 66832 5635
0 5637 5 1 1 5636
0 5638 7 1 2 47825 5637
0 5639 5 1 1 5638
0 5640 7 1 2 64550 64193
0 5641 5 1 1 5640
0 5642 7 1 2 5639 5641
0 5643 5 1 1 5642
0 5644 7 1 2 64348 5643
0 5645 5 1 1 5644
0 5646 7 10 2 52476 56980
0 5647 5 28 1 67196
0 5648 7 7 2 49528 67206
0 5649 5 2 1 67234
0 5650 7 2 2 64754 67235
0 5651 7 1 2 57818 67243
0 5652 5 1 1 5651
0 5653 7 1 2 5645 5652
0 5654 5 1 1 5653
0 5655 7 1 2 66496 5654
0 5656 5 1 1 5655
0 5657 7 1 2 63282 60085
0 5658 5 2 1 5657
0 5659 7 1 2 64156 67245
0 5660 5 1 1 5659
0 5661 7 1 2 47826 5660
0 5662 5 1 1 5661
0 5663 7 1 2 64973 5662
0 5664 5 1 1 5663
0 5665 7 1 2 57096 5664
0 5666 5 1 1 5665
0 5667 7 1 2 67170 5666
0 5668 5 1 1 5667
0 5669 7 1 2 48697 5668
0 5670 5 1 1 5669
0 5671 7 1 2 59576 65662
0 5672 5 1 1 5671
0 5673 7 1 2 5670 5672
0 5674 5 1 1 5673
0 5675 7 1 2 66542 5674
0 5676 5 1 1 5675
0 5677 7 1 2 5656 5676
0 5678 7 1 2 5633 5677
0 5679 7 1 2 5596 5678
0 5680 5 1 1 5679
0 5681 7 1 2 61544 5680
0 5682 5 1 1 5681
0 5683 7 1 2 61311 67091
0 5684 5 1 1 5683
0 5685 7 1 2 52593 2509
0 5686 5 2 1 5685
0 5687 7 1 2 48884 67172
0 5688 7 1 2 67247 5687
0 5689 5 1 1 5688
0 5690 7 1 2 5684 5689
0 5691 5 1 1 5690
0 5692 7 1 2 48588 5691
0 5693 5 1 1 5692
0 5694 7 2 2 53263 56981
0 5695 5 7 1 67249
0 5696 7 1 2 65619 67173
0 5697 7 1 2 67251 5696
0 5698 5 1 1 5697
0 5699 7 1 2 5693 5698
0 5700 5 1 1 5699
0 5701 7 1 2 49673 5700
0 5702 5 1 1 5701
0 5703 7 2 2 48885 49529
0 5704 7 4 2 48589 67258
0 5705 7 1 2 56325 65718
0 5706 7 1 2 67260 5705
0 5707 5 1 1 5706
0 5708 7 1 2 5702 5707
0 5709 5 1 1 5708
0 5710 7 1 2 56033 5709
0 5711 5 1 1 5710
0 5712 7 3 2 54888 67059
0 5713 7 1 2 57721 66813
0 5714 7 1 2 67264 5713
0 5715 5 1 1 5714
0 5716 7 1 2 5711 5715
0 5717 5 1 1 5716
0 5718 7 1 2 55225 5717
0 5719 5 1 1 5718
0 5720 7 2 2 63503 66065
0 5721 7 1 2 50364 67026
0 5722 7 1 2 67267 5721
0 5723 5 1 1 5722
0 5724 7 1 2 5719 5723
0 5725 5 1 1 5724
0 5726 7 1 2 62754 5725
0 5727 5 1 1 5726
0 5728 7 1 2 5682 5727
0 5729 7 1 2 5544 5728
0 5730 7 2 2 56034 63084
0 5731 5 1 1 67269
0 5732 7 1 2 48114 66754
0 5733 7 2 2 67270 5732
0 5734 7 1 2 67007 67271
0 5735 5 1 1 5734
0 5736 7 1 2 65062 66864
0 5737 5 1 1 5736
0 5738 7 1 2 65278 66989
0 5739 7 1 2 5737 5738
0 5740 5 1 1 5739
0 5741 7 1 2 5735 5740
0 5742 5 1 1 5741
0 5743 7 1 2 56823 5742
0 5744 5 1 1 5743
0 5745 7 4 2 48115 55452
0 5746 7 3 2 66492 67273
0 5747 7 1 2 64317 67277
0 5748 5 1 1 5747
0 5749 7 1 2 5744 5748
0 5750 5 1 1 5749
0 5751 7 1 2 55226 5750
0 5752 5 1 1 5751
0 5753 7 2 2 48116 49674
0 5754 7 1 2 64034 67280
0 5755 7 3 2 48590 65620
0 5756 7 4 2 54512 67174
0 5757 7 1 2 67282 67285
0 5758 7 1 2 5754 5757
0 5759 5 1 1 5758
0 5760 7 1 2 5752 5759
0 5761 5 1 1 5760
0 5762 7 1 2 49183 5761
0 5763 5 1 1 5762
0 5764 7 2 2 48591 64569
0 5765 7 1 2 48336 67289
0 5766 7 1 2 66524 5765
0 5767 5 1 1 5766
0 5768 7 1 2 5763 5767
0 5769 5 1 1 5768
0 5770 7 1 2 53969 5769
0 5771 5 1 1 5770
0 5772 7 4 2 55453 57879
0 5773 7 1 2 66540 67291
0 5774 5 1 1 5773
0 5775 7 1 2 5771 5774
0 5776 5 1 1 5775
0 5777 7 1 2 47827 5776
0 5778 5 1 1 5777
0 5779 7 7 2 53970 57138
0 5780 5 3 1 67295
0 5781 7 1 2 54513 64738
0 5782 5 1 1 5781
0 5783 7 1 2 63846 5782
0 5784 5 1 1 5783
0 5785 7 1 2 67296 5784
0 5786 5 1 1 5785
0 5787 7 1 2 64458 5786
0 5788 5 1 1 5787
0 5789 7 1 2 49300 5788
0 5790 5 1 1 5789
0 5791 7 4 2 54514 56530
0 5792 5 1 1 67305
0 5793 7 1 2 55227 67306
0 5794 5 2 1 5793
0 5795 7 1 2 5790 67309
0 5796 5 1 1 5795
0 5797 7 1 2 56824 5796
0 5798 5 1 1 5797
0 5799 7 1 2 62344 66121
0 5800 5 1 1 5799
0 5801 7 1 2 64750 5800
0 5802 5 1 1 5801
0 5803 7 1 2 55228 5802
0 5804 5 1 1 5803
0 5805 7 1 2 5798 5804
0 5806 5 1 1 5805
0 5807 7 1 2 48337 5806
0 5808 5 1 1 5807
0 5809 7 1 2 56531 64438
0 5810 5 1 1 5809
0 5811 7 1 2 48117 64448
0 5812 5 1 1 5811
0 5813 7 1 2 5810 5812
0 5814 5 1 1 5813
0 5815 7 1 2 56825 5814
0 5816 5 1 1 5815
0 5817 7 1 2 2967 5816
0 5818 5 1 1 5817
0 5819 7 1 2 54515 5818
0 5820 5 1 1 5819
0 5821 7 3 2 48592 64194
0 5822 7 1 2 56035 67311
0 5823 5 1 1 5822
0 5824 7 1 2 67310 5823
0 5825 5 1 1 5824
0 5826 7 1 2 56826 5825
0 5827 5 1 1 5826
0 5828 7 1 2 57880 64585
0 5829 5 2 1 5828
0 5830 7 1 2 5827 67314
0 5831 5 1 1 5830
0 5832 7 1 2 64856 5831
0 5833 5 1 1 5832
0 5834 7 1 2 5820 5833
0 5835 7 1 2 5808 5834
0 5836 5 1 1 5835
0 5837 7 1 2 66497 5836
0 5838 5 1 1 5837
0 5839 7 1 2 64505 58339
0 5840 5 1 1 5839
0 5841 7 1 2 63295 5840
0 5842 5 1 1 5841
0 5843 7 1 2 66404 5842
0 5844 5 1 1 5843
0 5845 7 1 2 54889 64857
0 5846 7 1 2 66389 5845
0 5847 5 1 1 5846
0 5848 7 1 2 5844 5847
0 5849 7 1 2 5838 5848
0 5850 5 1 1 5849
0 5851 7 1 2 54187 5850
0 5852 5 1 1 5851
0 5853 7 1 2 5778 5852
0 5854 7 1 2 5729 5853
0 5855 7 1 2 5372 5854
0 5856 7 1 2 5282 5855
0 5857 7 1 2 4876 5856
0 5858 5 1 1 5857
0 5859 7 1 2 55735 5858
0 5860 5 1 1 5859
0 5861 7 1 2 62280 62776
0 5862 7 1 2 65861 5861
0 5863 5 2 1 5862
0 5864 7 1 2 58371 65764
0 5865 5 1 1 5864
0 5866 7 1 2 4047 5865
0 5867 5 1 1 5866
0 5868 7 1 2 49184 5867
0 5869 5 1 1 5868
0 5870 7 1 2 65753 5869
0 5871 5 1 1 5870
0 5872 7 1 2 48338 5871
0 5873 5 1 1 5872
0 5874 7 3 2 53971 59671
0 5875 7 1 2 909 59633
0 5876 5 1 1 5875
0 5877 7 1 2 67318 5876
0 5878 5 1 1 5877
0 5879 7 1 2 59444 63365
0 5880 5 1 1 5879
0 5881 7 1 2 5878 5880
0 5882 5 2 1 5881
0 5883 7 1 2 48118 67321
0 5884 5 1 1 5883
0 5885 7 1 2 5884 65780
0 5886 5 1 1 5885
0 5887 7 1 2 54516 5886
0 5888 5 1 1 5887
0 5889 7 1 2 5873 5888
0 5890 5 1 1 5889
0 5891 7 1 2 49425 5890
0 5892 5 1 1 5891
0 5893 7 1 2 65925 5892
0 5894 5 1 1 5893
0 5895 7 1 2 48494 5894
0 5896 5 1 1 5895
0 5897 7 1 2 67316 5896
0 5898 5 1 1 5897
0 5899 7 1 2 5898 66562
0 5900 5 1 1 5899
0 5901 7 17 2 49530 50929
0 5902 5 5 1 67323
0 5903 7 6 2 48593 67324
0 5904 7 2 2 66883 67345
0 5905 5 1 1 67351
0 5906 7 1 2 67352 66057
0 5907 5 1 1 5906
0 5908 7 1 2 55229 65835
0 5909 5 1 1 5908
0 5910 7 2 2 58250 65893
0 5911 5 1 1 67353
0 5912 7 1 2 64941 5911
0 5913 5 1 1 5912
0 5914 7 1 2 56827 5913
0 5915 5 1 1 5914
0 5916 7 1 2 5909 5915
0 5917 5 1 1 5916
0 5918 7 1 2 58372 5917
0 5919 5 1 1 5918
0 5920 7 1 2 3083 5919
0 5921 5 1 1 5920
0 5922 7 1 2 49185 5921
0 5923 5 1 1 5922
0 5924 7 1 2 55230 66142
0 5925 5 1 1 5924
0 5926 7 2 2 57766 60967
0 5927 5 1 1 67355
0 5928 7 1 2 56326 64938
0 5929 7 1 2 67356 5928
0 5930 5 1 1 5929
0 5931 7 1 2 60798 67054
0 5932 5 1 1 5931
0 5933 7 1 2 65493 5932
0 5934 7 1 2 5930 5933
0 5935 7 1 2 5925 5934
0 5936 5 1 1 5935
0 5937 7 1 2 56036 5936
0 5938 5 1 1 5937
0 5939 7 2 2 63137 60629
0 5940 7 2 2 59805 67357
0 5941 7 1 2 56828 67359
0 5942 5 1 1 5941
0 5943 7 1 2 51216 5942
0 5944 5 1 1 5943
0 5945 7 1 2 54890 5944
0 5946 5 1 1 5945
0 5947 7 1 2 57414 66148
0 5948 5 1 1 5947
0 5949 7 1 2 65584 58282
0 5950 5 1 1 5949
0 5951 7 1 2 51217 5950
0 5952 5 2 1 5951
0 5953 7 1 2 48119 67361
0 5954 5 1 1 5953
0 5955 7 3 2 57841 65384
0 5956 5 2 1 67363
0 5957 7 3 2 64655 62125
0 5958 5 1 1 67368
0 5959 7 1 2 67366 67369
0 5960 5 1 1 5959
0 5961 7 1 2 5954 5960
0 5962 5 1 1 5961
0 5963 7 1 2 56327 5962
0 5964 5 1 1 5963
0 5965 7 1 2 5948 5964
0 5966 7 1 2 5946 5965
0 5967 7 1 2 5938 5966
0 5968 7 1 2 5923 5967
0 5969 5 1 1 5968
0 5970 7 1 2 53628 5969
0 5971 5 1 1 5970
0 5972 7 1 2 5907 5971
0 5973 5 1 1 5972
0 5974 7 1 2 54517 5973
0 5975 5 1 1 5974
0 5976 7 3 2 48120 64305
0 5977 7 2 2 62285 67371
0 5978 7 1 2 66755 67374
0 5979 5 1 1 5978
0 5980 7 1 2 5979 66794
0 5981 5 1 1 5980
0 5982 7 1 2 47828 5981
0 5983 5 1 1 5982
0 5984 7 1 2 65372 66876
0 5985 5 1 1 5984
0 5986 7 1 2 65556 64903
0 5987 5 2 1 5986
0 5988 7 2 2 58373 66732
0 5989 7 1 2 67376 67378
0 5990 5 1 1 5989
0 5991 7 1 2 5985 5990
0 5992 5 1 1 5991
0 5993 7 1 2 49186 5992
0 5994 5 1 1 5993
0 5995 7 1 2 5983 5994
0 5996 5 1 1 5995
0 5997 7 1 2 56037 5996
0 5998 5 1 1 5997
0 5999 7 3 2 56829 59252
0 6000 5 1 1 67380
0 6001 7 1 2 51218 6000
0 6002 5 1 1 6001
0 6003 7 1 2 66756 6002
0 6004 5 1 1 6003
0 6005 7 2 2 54188 64259
0 6006 5 1 1 67383
0 6007 7 2 2 53871 63053
0 6008 7 1 2 66631 67385
0 6009 7 1 2 67384 6008
0 6010 5 1 1 6009
0 6011 7 1 2 53629 65318
0 6012 7 1 2 64803 6011
0 6013 5 1 1 6012
0 6014 7 1 2 6010 6013
0 6015 5 1 1 6014
0 6016 7 1 2 47829 6015
0 6017 5 1 1 6016
0 6018 7 1 2 6004 6017
0 6019 7 1 2 5998 6018
0 6020 5 1 1 6019
0 6021 7 1 2 53972 6020
0 6022 5 1 1 6021
0 6023 7 1 2 56982 59697
0 6024 5 1 1 6023
0 6025 7 1 2 65491 6024
0 6026 5 1 1 6025
0 6027 7 2 2 47830 58227
0 6028 7 2 2 65433 58133
0 6029 7 1 2 67387 67389
0 6030 5 1 1 6029
0 6031 7 1 2 51219 6030
0 6032 5 1 1 6031
0 6033 7 1 2 59672 6032
0 6034 5 1 1 6033
0 6035 7 1 2 48121 64889
0 6036 5 1 1 6035
0 6037 7 2 2 64326 59525
0 6038 5 1 1 67391
0 6039 7 1 2 65328 60348
0 6040 7 1 2 67392 6039
0 6041 5 1 1 6040
0 6042 7 1 2 3251 6041
0 6043 7 1 2 6036 6042
0 6044 7 1 2 6034 6043
0 6045 5 1 1 6044
0 6046 7 1 2 54891 6045
0 6047 5 1 1 6046
0 6048 7 1 2 6026 6047
0 6049 5 1 1 6048
0 6050 7 1 2 53630 6049
0 6051 5 1 1 6050
0 6052 7 1 2 66461 66321
0 6053 5 1 1 6052
0 6054 7 1 2 60457 66877
0 6055 5 1 1 6054
0 6056 7 1 2 6053 6055
0 6057 5 1 1 6056
0 6058 7 1 2 59213 6057
0 6059 5 1 1 6058
0 6060 7 21 2 58570 56983
0 6061 5 1 1 67393
0 6062 7 1 2 59718 65814
0 6063 5 1 1 6062
0 6064 7 1 2 67394 6063
0 6065 5 1 1 6064
0 6066 7 1 2 66878 6065
0 6067 5 1 1 6066
0 6068 7 1 2 6059 6067
0 6069 7 1 2 6051 6068
0 6070 7 1 2 6022 6069
0 6071 7 1 2 5975 6070
0 6072 5 1 1 6071
0 6073 7 1 2 55454 6072
0 6074 5 1 1 6073
0 6075 7 1 2 61378 61040
0 6076 5 2 1 6075
0 6077 7 1 2 65719 67414
0 6078 5 1 1 6077
0 6079 7 7 2 54518 65966
0 6080 7 1 2 65117 58283
0 6081 7 1 2 67416 6080
0 6082 5 1 1 6081
0 6083 7 1 2 6078 6082
0 6084 5 1 1 6083
0 6085 7 1 2 47831 6084
0 6086 5 1 1 6085
0 6087 7 1 2 49187 65720
0 6088 7 1 2 59214 6087
0 6089 5 1 1 6088
0 6090 7 1 2 6086 6089
0 6091 5 1 1 6090
0 6092 7 1 2 65203 6091
0 6093 5 1 1 6092
0 6094 7 1 2 56038 65091
0 6095 5 1 1 6094
0 6096 7 1 2 52934 6095
0 6097 5 1 1 6096
0 6098 7 1 2 53052 65930
0 6099 5 1 1 6098
0 6100 7 1 2 6097 6099
0 6101 5 1 1 6100
0 6102 7 1 2 65105 6101
0 6103 5 1 1 6102
0 6104 7 1 2 65721 6103
0 6105 5 1 1 6104
0 6106 7 4 2 57415 57767
0 6107 5 1 1 67423
0 6108 7 1 2 58374 62190
0 6109 7 1 2 67417 6108
0 6110 7 1 2 67424 6109
0 6111 5 1 1 6110
0 6112 7 1 2 6105 6111
0 6113 5 1 1 6112
0 6114 7 1 2 48495 6113
0 6115 5 1 1 6114
0 6116 7 1 2 58160 63925
0 6117 5 1 1 6116
0 6118 7 1 2 62040 59537
0 6119 5 1 1 6118
0 6120 7 1 2 58553 65349
0 6121 5 1 1 6120
0 6122 7 1 2 6121 66928
0 6123 7 1 2 6119 6122
0 6124 7 1 2 6117 6123
0 6125 7 1 2 58297 65688
0 6126 5 1 1 6125
0 6127 7 2 2 50631 58179
0 6128 5 3 1 67427
0 6129 7 1 2 53973 67429
0 6130 5 1 1 6129
0 6131 7 1 2 58210 61416
0 6132 7 1 2 6130 6131
0 6133 5 1 1 6132
0 6134 7 1 2 6126 6133
0 6135 5 1 1 6134
0 6136 7 1 2 54189 61051
0 6137 5 2 1 6136
0 6138 7 1 2 52228 58560
0 6139 7 1 2 67432 6138
0 6140 5 1 1 6139
0 6141 7 2 2 50632 58561
0 6142 5 1 1 67434
0 6143 7 1 2 60284 6142
0 6144 7 1 2 6140 6143
0 6145 5 1 1 6144
0 6146 7 1 2 6135 6145
0 6147 7 1 2 6124 6146
0 6148 5 1 1 6147
0 6149 7 1 2 65722 6148
0 6150 5 1 1 6149
0 6151 7 1 2 6115 6150
0 6152 7 1 2 6093 6151
0 6153 5 1 1 6152
0 6154 7 1 2 54892 6153
0 6155 5 1 1 6154
0 6156 7 4 2 54190 66576
0 6157 5 1 1 67436
0 6158 7 1 2 66721 65863
0 6159 5 1 1 6158
0 6160 7 1 2 6157 6159
0 6161 5 1 1 6160
0 6162 7 1 2 56039 6161
0 6163 5 1 1 6162
0 6164 7 1 2 50140 61042
0 6165 5 7 1 6164
0 6166 7 1 2 67440 66726
0 6167 5 1 1 6166
0 6168 7 1 2 61745 67379
0 6169 5 1 1 6168
0 6170 7 1 2 6167 6169
0 6171 7 1 2 6163 6170
0 6172 5 1 1 6171
0 6173 7 1 2 48122 6172
0 6174 5 1 1 6173
0 6175 7 1 2 56040 63170
0 6176 7 1 2 66597 6175
0 6177 7 1 2 58284 6176
0 6178 5 1 1 6177
0 6179 7 1 2 6174 6178
0 6180 5 1 1 6179
0 6181 7 1 2 54519 6180
0 6182 5 1 1 6181
0 6183 7 3 2 58146 59445
0 6184 5 1 1 67447
0 6185 7 2 2 62210 67448
0 6186 7 2 2 60320 67450
0 6187 7 1 2 66632 67452
0 6188 5 1 1 6187
0 6189 7 1 2 6182 6188
0 6190 5 1 1 6189
0 6191 7 1 2 56328 6190
0 6192 5 1 1 6191
0 6193 7 1 2 51220 65926
0 6194 5 1 1 6193
0 6195 7 1 2 53631 6194
0 6196 5 1 1 6195
0 6197 7 2 2 56830 66598
0 6198 7 1 2 57574 67364
0 6199 5 1 1 6198
0 6200 7 1 2 56041 60285
0 6201 7 1 2 6199 6200
0 6202 5 1 1 6201
0 6203 7 1 2 63235 5927
0 6204 5 1 1 6203
0 6205 7 1 2 48123 6204
0 6206 5 1 1 6205
0 6207 7 1 2 47832 66163
0 6208 5 1 1 6207
0 6209 7 1 2 61276 6208
0 6210 7 1 2 6206 6209
0 6211 7 1 2 6202 6210
0 6212 5 1 1 6211
0 6213 7 1 2 50633 6212
0 6214 5 1 1 6213
0 6215 7 1 2 48124 67441
0 6216 5 3 1 6215
0 6217 7 1 2 55848 67456
0 6218 5 2 1 6217
0 6219 7 1 2 62630 67459
0 6220 5 1 1 6219
0 6221 7 1 2 6214 6220
0 6222 5 1 1 6221
0 6223 7 1 2 67454 6222
0 6224 5 1 1 6223
0 6225 7 1 2 6196 6224
0 6226 7 1 2 6192 6225
0 6227 5 1 1 6226
0 6228 7 1 2 55455 6227
0 6229 5 1 1 6228
0 6230 7 1 2 6155 6229
0 6231 5 1 1 6230
0 6232 7 1 2 56532 6231
0 6233 5 1 1 6232
0 6234 7 1 2 58641 63221
0 6235 5 1 1 6234
0 6236 7 1 2 61168 65832
0 6237 5 1 1 6236
0 6238 7 1 2 58375 59215
0 6239 7 1 2 6237 6238
0 6240 5 1 1 6239
0 6241 7 1 2 6235 6240
0 6242 5 1 1 6241
0 6243 7 1 2 49188 6242
0 6244 5 1 1 6243
0 6245 7 1 2 59647 58886
0 6246 5 3 1 6245
0 6247 7 1 2 56831 67461
0 6248 5 1 1 6247
0 6249 7 1 2 59087 61116
0 6250 5 1 1 6249
0 6251 7 1 2 57575 63880
0 6252 5 1 1 6251
0 6253 7 1 2 56329 6252
0 6254 7 1 2 6250 6253
0 6255 5 1 1 6254
0 6256 7 1 2 6248 6255
0 6257 7 1 2 6244 6256
0 6258 5 1 1 6257
0 6259 7 1 2 54520 6258
0 6260 5 1 1 6259
0 6261 7 1 2 63247 63267
0 6262 5 1 1 6261
0 6263 7 1 2 56984 6262
0 6264 5 1 1 6263
0 6265 7 1 2 58306 6264
0 6266 5 1 1 6265
0 6267 7 2 2 52229 62339
0 6268 5 2 1 67464
0 6269 7 1 2 56330 61374
0 6270 7 2 2 58161 6269
0 6271 7 1 2 67466 67468
0 6272 5 1 1 6271
0 6273 7 1 2 6266 6272
0 6274 5 1 1 6273
0 6275 7 1 2 54191 6274
0 6276 5 1 1 6275
0 6277 7 1 2 6260 6276
0 6278 5 1 1 6277
0 6279 7 1 2 66918 6278
0 6280 5 1 1 6279
0 6281 7 1 2 48125 67145
0 6282 5 1 1 6281
0 6283 7 1 2 66010 6282
0 6284 5 1 1 6283
0 6285 7 1 2 64804 6284
0 6286 5 1 1 6285
0 6287 7 1 2 66435 6286
0 6288 5 1 1 6287
0 6289 7 1 2 56331 6288
0 6290 5 1 1 6289
0 6291 7 4 2 54893 66733
0 6292 5 1 1 67470
0 6293 7 1 2 56832 67471
0 6294 5 1 1 6293
0 6295 7 1 2 5905 6294
0 6296 5 1 1 6295
0 6297 7 1 2 48126 6296
0 6298 5 1 1 6297
0 6299 7 6 2 49301 53632
0 6300 7 1 2 65136 67474
0 6301 5 1 1 6300
0 6302 7 1 2 6298 6301
0 6303 5 1 1 6302
0 6304 7 1 2 55456 6303
0 6305 5 1 1 6304
0 6306 7 2 2 65694 67175
0 6307 5 2 1 67480
0 6308 7 1 2 57881 67481
0 6309 5 1 1 6308
0 6310 7 1 2 6305 6309
0 6311 7 1 2 6290 6310
0 6312 5 1 1 6311
0 6313 7 1 2 54521 6312
0 6314 5 1 1 6313
0 6315 7 1 2 65118 67075
0 6316 5 1 1 6315
0 6317 7 1 2 67286 66327
0 6318 5 1 1 6317
0 6319 7 1 2 5461 6318
0 6320 5 1 1 6319
0 6321 7 1 2 56332 6320
0 6322 5 1 1 6321
0 6323 7 1 2 6322 5437
0 6324 5 1 1 6323
0 6325 7 1 2 55231 6324
0 6326 5 1 1 6325
0 6327 7 1 2 66310 66911
0 6328 5 1 1 6327
0 6329 7 1 2 6326 6328
0 6330 5 1 1 6329
0 6331 7 1 2 56042 6330
0 6332 5 1 1 6331
0 6333 7 1 2 6316 6332
0 6334 7 1 2 6314 6333
0 6335 5 1 1 6334
0 6336 7 1 2 67442 6335
0 6337 5 1 1 6336
0 6338 7 1 2 6280 6337
0 6339 7 1 2 6233 6338
0 6340 7 1 2 6074 6339
0 6341 5 1 1 6340
0 6342 7 1 2 48886 6341
0 6343 5 1 1 6342
0 6344 7 1 2 5900 6343
0 6345 5 1 1 6344
0 6346 7 1 2 62534 6345
0 6347 5 1 1 6346
0 6348 7 1 2 65531 66981
0 6349 5 1 1 6348
0 6350 7 1 2 5396 6349
0 6351 5 1 1 6350
0 6352 7 1 2 60286 6351
0 6353 5 1 1 6352
0 6354 7 2 2 56833 58090
0 6355 5 1 1 67484
0 6356 7 1 2 58738 6355
0 6357 5 3 1 6356
0 6358 7 1 2 51492 62320
0 6359 7 1 2 63400 6358
0 6360 7 1 2 67486 6359
0 6361 5 1 1 6360
0 6362 7 1 2 6353 6361
0 6363 5 1 1 6362
0 6364 7 1 2 48887 6363
0 6365 5 1 1 6364
0 6366 7 3 2 55457 62888
0 6367 7 3 2 53633 67489
0 6368 7 3 2 63307 60287
0 6369 7 1 2 67492 67495
0 6370 5 1 1 6369
0 6371 7 1 2 6365 6370
0 6372 5 1 1 6371
0 6373 7 1 2 47833 6372
0 6374 5 1 1 6373
0 6375 7 2 2 53974 57097
0 6376 5 3 1 67498
0 6377 7 1 2 171 67500
0 6378 5 2 1 6377
0 6379 7 1 2 67060 67472
0 6380 7 1 2 67503 6379
0 6381 5 1 1 6380
0 6382 7 1 2 6374 6381
0 6383 5 1 1 6382
0 6384 7 1 2 55232 6383
0 6385 5 1 1 6384
0 6386 7 2 2 49531 60288
0 6387 7 2 2 48496 48698
0 6388 7 6 2 66526 67507
0 6389 7 2 2 66394 67509
0 6390 7 1 2 67505 67515
0 6391 5 1 1 6390
0 6392 7 5 2 53975 51493
0 6393 7 1 2 67027 67517
0 6394 5 1 1 6393
0 6395 7 1 2 5422 6394
0 6396 5 1 1 6395
0 6397 7 1 2 67252 6396
0 6398 5 1 1 6397
0 6399 7 1 2 67274 66577
0 6400 7 1 2 57350 6399
0 6401 7 1 2 64554 6400
0 6402 5 1 1 6401
0 6403 7 1 2 6398 6402
0 6404 5 1 1 6403
0 6405 7 1 2 48594 6404
0 6406 5 1 1 6405
0 6407 7 1 2 6391 6406
0 6408 5 1 1 6407
0 6409 7 1 2 64135 6408
0 6410 5 1 1 6409
0 6411 7 1 2 6385 6410
0 6412 5 1 1 6411
0 6413 7 1 2 54522 6412
0 6414 5 1 1 6413
0 6415 7 1 2 55458 62321
0 6416 7 1 2 67168 6415
0 6417 5 1 1 6416
0 6418 7 1 2 6414 6417
0 6419 5 1 1 6418
0 6420 7 1 2 56043 6419
0 6421 5 1 1 6420
0 6422 7 15 2 50141 51221
0 6423 5 3 1 67522
0 6424 7 1 2 48127 50930
0 6425 7 1 2 67523 6424
0 6426 5 1 1 6425
0 6427 7 1 2 4925 6426
0 6428 5 1 1 6427
0 6429 7 1 2 63993 6428
0 6430 5 1 1 6429
0 6431 7 1 2 63261 66779
0 6432 5 1 1 6431
0 6433 7 1 2 6430 6432
0 6434 5 1 1 6433
0 6435 7 1 2 54192 6434
0 6436 5 1 1 6435
0 6437 7 7 2 47834 53634
0 6438 7 1 2 64939 67540
0 6439 5 2 1 6438
0 6440 7 1 2 6436 67547
0 6441 5 1 1 6440
0 6442 7 1 2 56333 6441
0 6443 5 1 1 6442
0 6444 7 10 2 54193 51222
0 6445 7 4 2 50931 56834
0 6446 7 2 2 67559 66803
0 6447 5 1 1 67563
0 6448 7 1 2 67549 67564
0 6449 5 1 1 6448
0 6450 7 1 2 66626 6449
0 6451 5 1 1 6450
0 6452 7 1 2 63112 6451
0 6453 5 1 1 6452
0 6454 7 1 2 67548 4979
0 6455 5 1 1 6454
0 6456 7 1 2 57416 6455
0 6457 5 1 1 6456
0 6458 7 9 2 54194 63439
0 6459 7 1 2 67541 67565
0 6460 5 1 1 6459
0 6461 7 2 2 56044 65319
0 6462 7 1 2 66780 67574
0 6463 5 1 1 6462
0 6464 7 1 2 6460 6463
0 6465 7 1 2 6457 6464
0 6466 7 1 2 6453 6465
0 6467 7 1 2 6443 6466
0 6468 5 1 1 6467
0 6469 7 1 2 56533 6468
0 6470 5 1 1 6469
0 6471 7 1 2 64764 66781
0 6472 5 1 1 6471
0 6473 7 1 2 50142 65557
0 6474 5 1 1 6473
0 6475 7 1 2 47835 6474
0 6476 7 1 2 66874 6475
0 6477 5 1 1 6476
0 6478 7 1 2 6472 6477
0 6479 5 1 1 6478
0 6480 7 1 2 56045 6479
0 6481 5 1 1 6480
0 6482 7 2 2 60289 66971
0 6483 5 1 1 67576
0 6484 7 1 2 57842 62340
0 6485 5 8 1 6484
0 6486 7 1 2 59476 67578
0 6487 5 1 1 6486
0 6488 7 1 2 6483 6487
0 6489 5 1 1 6488
0 6490 7 1 2 57417 6489
0 6491 5 1 1 6490
0 6492 7 1 2 65537 57732
0 6493 5 1 1 6492
0 6494 7 1 2 51223 6493
0 6495 7 1 2 6491 6494
0 6496 5 1 1 6495
0 6497 7 1 2 66757 6496
0 6498 5 1 1 6497
0 6499 7 1 2 64739 66728
0 6500 5 1 1 6499
0 6501 7 1 2 65066 66758
0 6502 5 1 1 6501
0 6503 7 1 2 6500 6502
0 6504 5 1 1 6503
0 6505 7 1 2 63113 6504
0 6506 5 1 1 6505
0 6507 7 3 2 55233 60290
0 6508 7 1 2 66734 67586
0 6509 5 1 1 6508
0 6510 7 1 2 66880 6509
0 6511 5 1 1 6510
0 6512 7 1 2 59216 6511
0 6513 5 1 1 6512
0 6514 7 1 2 6506 6513
0 6515 7 1 2 6498 6514
0 6516 7 1 2 6481 6515
0 6517 7 1 2 6470 6516
0 6518 5 1 1 6517
0 6519 7 1 2 55459 6518
0 6520 5 1 1 6519
0 6521 7 2 2 56046 57733
0 6522 5 1 1 67589
0 6523 7 1 2 61117 6522
0 6524 5 2 1 6523
0 6525 7 1 2 3494 67591
0 6526 5 1 1 6525
0 6527 7 1 2 65538 60291
0 6528 5 1 1 6527
0 6529 7 1 2 6526 6528
0 6530 5 1 1 6529
0 6531 7 1 2 66919 6530
0 6532 5 1 1 6531
0 6533 7 1 2 67287 66912
0 6534 5 1 1 6533
0 6535 7 4 2 55460 56047
0 6536 7 1 2 53635 67593
0 6537 5 1 1 6536
0 6538 7 1 2 6534 6537
0 6539 5 1 1 6538
0 6540 7 1 2 56334 6539
0 6541 5 1 1 6540
0 6542 7 1 2 64449 67150
0 6543 5 1 1 6542
0 6544 7 1 2 65747 6543
0 6545 5 2 1 6544
0 6546 7 1 2 58275 67597
0 6547 5 1 1 6546
0 6548 7 1 2 6541 6547
0 6549 5 1 1 6548
0 6550 7 1 2 55234 6549
0 6551 5 1 1 6550
0 6552 7 2 2 62631 66599
0 6553 7 1 2 65596 67599
0 6554 5 1 1 6553
0 6555 7 1 2 64516 66735
0 6556 7 1 2 58340 6555
0 6557 5 1 1 6556
0 6558 7 1 2 6554 6557
0 6559 5 1 1 6558
0 6560 7 1 2 55461 6559
0 6561 5 1 1 6560
0 6562 7 1 2 58219 66677
0 6563 7 1 2 64885 6562
0 6564 5 1 1 6563
0 6565 7 1 2 6561 6564
0 6566 7 1 2 6551 6565
0 6567 5 1 1 6566
0 6568 7 1 2 59974 6567
0 6569 5 1 1 6568
0 6570 7 1 2 6532 6569
0 6571 7 1 2 6520 6570
0 6572 5 1 1 6571
0 6573 7 1 2 48888 6572
0 6574 5 1 1 6573
0 6575 7 2 2 58251 62709
0 6576 5 1 1 67601
0 6577 7 2 2 63155 6576
0 6578 5 1 1 67603
0 6579 7 3 2 57418 6578
0 6580 5 1 1 67605
0 6581 7 1 2 60321 63994
0 6582 5 1 1 6581
0 6583 7 1 2 6580 6582
0 6584 5 1 1 6583
0 6585 7 11 2 54894 55462
0 6586 7 3 2 67608 66462
0 6587 5 2 1 67619
0 6588 7 1 2 64287 67620
0 6589 7 1 2 6584 6588
0 6590 5 1 1 6589
0 6591 7 1 2 6574 6590
0 6592 5 1 1 6591
0 6593 7 1 2 62535 6592
0 6594 5 1 1 6593
0 6595 7 1 2 67160 67600
0 6596 5 1 1 6595
0 6597 7 2 2 64367 64870
0 6598 5 1 1 67624
0 6599 7 1 2 67625 67272
0 6600 5 1 1 6599
0 6601 7 1 2 6596 6600
0 6602 5 1 1 6601
0 6603 7 1 2 55463 6602
0 6604 5 1 1 6603
0 6605 7 1 2 59217 67044
0 6606 5 1 1 6605
0 6607 7 1 2 4835 6606
0 6608 5 1 1 6607
0 6609 7 1 2 54895 6608
0 6610 5 1 1 6609
0 6611 7 1 2 54195 67278
0 6612 7 1 2 65597 6611
0 6613 5 1 1 6612
0 6614 7 1 2 6610 6613
0 6615 5 1 1 6614
0 6616 7 1 2 54523 6615
0 6617 5 1 1 6616
0 6618 7 2 2 56048 67487
0 6619 7 2 2 49675 67176
0 6620 7 1 2 67626 67628
0 6621 5 1 1 6620
0 6622 7 1 2 66982 67104
0 6623 5 1 1 6622
0 6624 7 1 2 66558 6623
0 6625 5 1 1 6624
0 6626 7 1 2 58579 6625
0 6627 5 1 1 6626
0 6628 7 1 2 6621 6627
0 6629 5 1 1 6628
0 6630 7 1 2 48889 6629
0 6631 5 1 1 6630
0 6632 7 7 2 57882 62889
0 6633 5 2 1 67630
0 6634 7 1 2 65723 67631
0 6635 7 1 2 58580 6634
0 6636 5 1 1 6635
0 6637 7 1 2 6631 6636
0 6638 7 1 2 6617 6637
0 6639 5 1 1 6638
0 6640 7 1 2 55235 6639
0 6641 5 1 1 6640
0 6642 7 1 2 6604 6641
0 6643 5 1 1 6642
0 6644 7 1 2 59975 6643
0 6645 5 1 1 6644
0 6646 7 3 2 67063 67265
0 6647 7 1 2 49426 67639
0 6648 5 1 1 6647
0 6649 7 6 2 53636 67609
0 6650 5 2 1 67642
0 6651 7 1 2 67643 67261
0 6652 5 1 1 6651
0 6653 7 1 2 62822 67644
0 6654 5 1 1 6653
0 6655 7 1 2 49427 58091
0 6656 7 1 2 67139 6655
0 6657 5 1 1 6656
0 6658 7 1 2 6654 6657
0 6659 5 1 1 6658
0 6660 7 1 2 49676 6659
0 6661 5 1 1 6660
0 6662 7 1 2 6652 6661
0 6663 5 1 1 6662
0 6664 7 1 2 48497 6663
0 6665 5 1 1 6664
0 6666 7 1 2 6648 6665
0 6667 5 1 1 6666
0 6668 7 1 2 67579 6667
0 6669 5 1 1 6668
0 6670 7 10 2 49677 53976
0 6671 5 1 1 67650
0 6672 7 1 2 66395 67651
0 6673 7 1 2 58730 6672
0 6674 7 1 2 67377 6673
0 6675 5 1 1 6674
0 6676 7 1 2 6669 6675
0 6677 5 1 1 6676
0 6678 7 1 2 54524 6677
0 6679 5 1 1 6678
0 6680 7 1 2 67640 67577
0 6681 5 1 1 6680
0 6682 7 3 2 51494 60292
0 6683 7 1 2 65612 67660
0 6684 5 1 1 6683
0 6685 7 1 2 67648 6684
0 6686 5 1 1 6685
0 6687 7 1 2 56534 6686
0 6688 5 1 1 6687
0 6689 7 1 2 65501 67661
0 6690 5 1 1 6689
0 6691 7 1 2 6688 6690
0 6692 5 1 1 6691
0 6693 7 1 2 62890 6692
0 6694 5 1 1 6693
0 6695 7 2 2 55464 56535
0 6696 7 1 2 53637 64862
0 6697 7 1 2 67663 6696
0 6698 5 1 1 6697
0 6699 7 1 2 6694 6698
0 6700 5 1 1 6699
0 6701 7 1 2 56335 6700
0 6702 5 1 1 6701
0 6703 7 1 2 59053 64720
0 6704 5 1 1 6703
0 6705 7 1 2 58341 6704
0 6706 5 1 1 6705
0 6707 7 1 2 59044 66233
0 6708 5 1 1 6707
0 6709 7 1 2 6706 6708
0 6710 5 1 1 6709
0 6711 7 1 2 67061 66736
0 6712 7 1 2 6710 6711
0 6713 5 1 1 6712
0 6714 7 1 2 6702 6713
0 6715 5 1 1 6714
0 6716 7 1 2 55236 6715
0 6717 5 1 1 6716
0 6718 7 1 2 6681 6717
0 6719 7 1 2 6679 6718
0 6720 5 1 1 6719
0 6721 7 1 2 57419 6720
0 6722 5 1 1 6721
0 6723 7 3 2 47836 64781
0 6724 5 1 1 67665
0 6725 7 1 2 56536 67666
0 6726 5 1 1 6725
0 6727 7 1 2 53977 67312
0 6728 5 1 1 6727
0 6729 7 1 2 6726 6728
0 6730 5 1 1 6729
0 6731 7 1 2 66516 6730
0 6732 5 1 1 6731
0 6733 7 1 2 6732 66317
0 6734 5 1 1 6733
0 6735 7 1 2 67028 6734
0 6736 5 1 1 6735
0 6737 7 1 2 60322 64826
0 6738 7 1 2 66498 6737
0 6739 5 1 1 6738
0 6740 7 1 2 6736 6739
0 6741 5 1 1 6740
0 6742 7 1 2 59218 6741
0 6743 5 1 1 6742
0 6744 7 2 2 47837 62891
0 6745 7 1 2 67140 67668
0 6746 7 1 2 67496 6745
0 6747 5 1 1 6746
0 6748 7 1 2 6743 6747
0 6749 7 1 2 64426 66623
0 6750 5 1 1 6749
0 6751 7 1 2 66729 67023
0 6752 5 1 1 6751
0 6753 7 1 2 6750 6752
0 6754 5 1 1 6753
0 6755 7 1 2 55465 6754
0 6756 5 1 1 6755
0 6757 7 2 2 47838 66737
0 6758 7 1 2 67266 67670
0 6759 5 1 1 6758
0 6760 7 1 2 6759 67035
0 6761 5 1 1 6760
0 6762 7 1 2 56336 64723
0 6763 7 1 2 6761 6762
0 6764 5 1 1 6763
0 6765 7 1 2 6756 6764
0 6766 5 1 1 6765
0 6767 7 1 2 63114 6766
0 6768 5 1 1 6767
0 6769 7 1 2 57883 64983
0 6770 5 1 1 6769
0 6771 7 1 2 64725 6770
0 6772 5 1 1 6771
0 6773 7 1 2 56835 6772
0 6774 5 1 1 6773
0 6775 7 1 2 64830 6774
0 6776 5 1 1 6775
0 6777 7 1 2 66499 6776
0 6778 5 1 1 6777
0 6779 7 16 2 49678 55237
0 6780 5 4 1 67672
0 6781 7 8 2 54196 51495
0 6782 7 2 2 67673 67692
0 6783 5 1 1 67700
0 6784 7 1 2 65621 67701
0 6785 7 1 2 67504 6784
0 6786 5 1 1 6785
0 6787 7 1 2 6778 6786
0 6788 5 1 1 6787
0 6789 7 1 2 54896 6788
0 6790 5 1 1 6789
0 6791 7 1 2 6768 6790
0 6792 7 1 2 6748 6791
0 6793 7 1 2 6722 6792
0 6794 7 1 2 6645 6793
0 6795 7 1 2 6594 6794
0 6796 7 1 2 6421 6795
0 6797 5 1 1 6796
0 6798 7 1 2 58602 6797
0 6799 5 1 1 6798
0 6800 7 1 2 63308 64755
0 6801 5 1 1 6800
0 6802 7 1 2 57098 64756
0 6803 5 1 1 6802
0 6804 7 1 2 6598 6803
0 6805 5 1 1 6804
0 6806 7 1 2 65055 6805
0 6807 5 1 1 6806
0 6808 7 1 2 6801 6807
0 6809 5 1 1 6808
0 6810 7 1 2 66493 6809
0 6811 5 1 1 6810
0 6812 7 2 2 62676 66884
0 6813 5 2 1 67702
0 6814 7 1 2 48128 65622
0 6815 7 1 2 67703 6814
0 6816 5 1 1 6815
0 6817 7 1 2 6811 6816
0 6818 5 1 1 6817
0 6819 7 1 2 55466 6818
0 6820 5 1 1 6819
0 6821 7 2 2 57884 61106
0 6822 5 1 1 67706
0 6823 7 1 2 64726 6822
0 6824 5 1 1 6823
0 6825 7 1 2 65056 6824
0 6826 5 1 1 6825
0 6827 7 1 2 64831 6826
0 6828 5 1 1 6827
0 6829 7 1 2 6828 66500
0 6830 5 1 1 6829
0 6831 7 1 2 2987 5528
0 6832 5 1 1 6831
0 6833 7 1 2 66405 6832
0 6834 5 1 1 6833
0 6835 7 1 2 6830 6834
0 6836 5 1 1 6835
0 6837 7 1 2 56337 6836
0 6838 5 1 1 6837
0 6839 7 1 2 57420 58252
0 6840 7 1 2 67488 6839
0 6841 5 1 1 6840
0 6842 7 1 2 48699 65600
0 6843 5 1 1 6842
0 6844 7 1 2 6841 6843
0 6845 5 1 1 6844
0 6846 7 1 2 66543 6845
0 6847 5 1 1 6846
0 6848 7 1 2 6838 6847
0 6849 7 1 2 6820 6848
0 6850 5 1 1 6849
0 6851 7 1 2 54525 6850
0 6852 5 1 1 6851
0 6853 7 2 2 52069 56985
0 6854 5 3 1 67708
0 6855 7 2 2 67710 66200
0 6856 7 1 2 67713 66983
0 6857 5 1 1 6856
0 6858 7 1 2 66534 67046
0 6859 5 1 1 6858
0 6860 7 1 2 6857 6859
0 6861 5 1 1 6860
0 6862 7 1 2 56537 6861
0 6863 5 1 1 6862
0 6864 7 6 2 54197 67008
0 6865 7 1 2 67064 67715
0 6866 5 1 1 6865
0 6867 7 1 2 56836 65057
0 6868 5 2 1 6867
0 6869 7 1 2 62833 67721
0 6870 5 1 1 6869
0 6871 7 1 2 49679 66990
0 6872 7 1 2 6870 6871
0 6873 5 1 1 6872
0 6874 7 1 2 6866 6873
0 6875 7 1 2 6863 6874
0 6876 5 1 1 6875
0 6877 7 1 2 48890 6876
0 6878 5 1 1 6877
0 6879 7 3 2 50365 57980
0 6880 5 2 1 67723
0 6881 7 6 2 50932 57981
0 6882 5 3 1 67728
0 6883 7 1 2 56538 67734
0 6884 7 2 2 67726 6883
0 6885 7 1 2 67737 67279
0 6886 5 1 1 6885
0 6887 7 2 2 64136 66517
0 6888 7 1 2 67161 67739
0 6889 5 1 1 6888
0 6890 7 1 2 6886 6889
0 6891 5 1 1 6890
0 6892 7 1 2 56338 6891
0 6893 5 1 1 6892
0 6894 7 1 2 58664 67493
0 6895 7 1 2 63309 6894
0 6896 5 1 1 6895
0 6897 7 1 2 6893 6896
0 6898 7 1 2 6878 6897
0 6899 5 1 1 6898
0 6900 7 1 2 55238 6899
0 6901 5 1 1 6900
0 6902 7 1 2 62625 66215
0 6903 7 1 2 67029 6902
0 6904 5 1 1 6903
0 6905 7 1 2 6901 6904
0 6906 5 1 1 6905
0 6907 7 1 2 56049 6906
0 6908 5 1 1 6907
0 6909 7 1 2 57421 67641
0 6910 5 1 1 6909
0 6911 7 1 2 56539 66406
0 6912 5 1 1 6911
0 6913 7 1 2 6910 6912
0 6914 5 1 1 6913
0 6915 7 1 2 56837 6914
0 6916 5 1 1 6915
0 6917 7 3 2 64570 65967
0 6918 7 1 2 67283 67741
0 6919 5 1 1 6918
0 6920 7 1 2 6916 6919
0 6921 5 1 1 6920
0 6922 7 1 2 54198 6921
0 6923 5 1 1 6922
0 6924 7 1 2 64560 61312
0 6925 7 2 2 49680 64782
0 6926 5 1 1 67744
0 6927 7 1 2 67151 67745
0 6928 7 1 2 6924 6927
0 6929 5 1 1 6928
0 6930 7 1 2 6923 6929
0 6931 7 1 2 6908 6930
0 6932 7 1 2 6852 6931
0 6933 5 1 1 6932
0 6934 7 1 2 6933 67443
0 6935 5 1 1 6934
0 6936 7 1 2 67494 65955
0 6937 5 1 1 6936
0 6938 7 1 2 6935 6937
0 6939 7 1 2 6799 6938
0 6940 7 1 2 6347 6939
0 6941 7 1 2 5860 6940
0 6942 7 1 2 4798 6941
0 6943 7 1 2 4136 6942
0 6944 5 1 1 6943
0 6945 7 1 2 55593 6944
0 6946 5 1 1 6945
0 6947 7 2 2 50933 58713
0 6948 5 11 1 67746
0 6949 7 36 2 49831 51496
0 6950 5 9 1 67759
0 6951 7 1 2 5548 67795
0 6952 5 2 1 6951
0 6953 7 1 2 64372 67804
0 6954 5 1 1 6953
0 6955 7 10 2 53423 51224
0 6956 5 1 1 67806
0 6957 7 1 2 48700 67807
0 6958 5 3 1 6957
0 6959 7 1 2 59011 67816
0 6960 5 2 1 6959
0 6961 7 15 2 49832 55467
0 6962 7 1 2 57422 67821
0 6963 7 1 2 67819 6962
0 6964 5 1 1 6963
0 6965 7 1 2 6954 6964
0 6966 5 1 1 6965
0 6967 7 1 2 56339 6966
0 6968 5 1 1 6967
0 6969 7 7 2 52758 49833
0 6970 5 3 1 67836
0 6971 7 5 2 67130 67843
0 6972 5 20 1 67846
0 6973 7 6 2 49681 67851
0 6974 5 2 1 67871
0 6975 7 13 2 49834 51225
0 6976 5 1 1 67879
0 6977 7 1 2 53424 67880
0 6978 5 4 1 6977
0 6979 7 1 2 67131 67892
0 6980 5 1 1 6979
0 6981 7 1 2 48701 6980
0 6982 5 1 1 6981
0 6983 7 1 2 67877 6982
0 6984 5 1 1 6983
0 6985 7 1 2 66535 6984
0 6986 5 1 1 6985
0 6987 7 1 2 6968 6986
0 6988 5 1 1 6987
0 6989 7 1 2 55594 6988
0 6990 5 1 1 6989
0 6991 7 9 2 49835 55239
0 6992 7 52 2 55468 51683
0 6993 7 1 2 67896 67905
0 6994 7 1 2 67162 6993
0 6995 5 1 1 6994
0 6996 7 1 2 6990 6995
0 6997 5 1 1 6996
0 6998 7 1 2 56540 6997
0 6999 5 1 1 6998
0 7000 7 1 2 49682 58092
0 7001 5 2 1 7000
0 7002 7 1 2 65494 67957
0 7003 5 1 1 7002
0 7004 7 1 2 52759 58961
0 7005 7 1 2 7003 7004
0 7006 5 1 1 7005
0 7007 7 6 2 52594 48891
0 7008 5 1 1 67959
0 7009 7 4 2 48702 49532
0 7010 5 2 1 67965
0 7011 7 2 2 53425 67966
0 7012 7 1 2 48595 67971
0 7013 5 1 1 7012
0 7014 7 1 2 7008 7013
0 7015 5 1 1 7014
0 7016 7 1 2 51226 7015
0 7017 5 1 1 7016
0 7018 7 1 2 49836 7017
0 7019 7 1 2 7006 7018
0 7020 5 1 1 7019
0 7021 7 1 2 63061 64376
0 7022 5 1 1 7021
0 7023 7 3 2 57982 64377
0 7024 5 1 1 67973
0 7025 7 1 2 65492 7024
0 7026 7 1 2 7022 7025
0 7027 5 1 1 7026
0 7028 7 2 2 53426 57983
0 7029 5 4 1 67976
0 7030 7 3 2 58093 67978
0 7031 5 5 1 67982
0 7032 7 6 2 62536 67983
0 7033 7 1 2 48892 67990
0 7034 5 1 1 7033
0 7035 7 1 2 53638 7034
0 7036 7 1 2 7027 7035
0 7037 5 1 1 7036
0 7038 7 1 2 55595 7037
0 7039 7 1 2 7020 7038
0 7040 5 1 1 7039
0 7041 7 2 2 58939 58094
0 7042 5 1 1 67996
0 7043 7 4 2 51684 67897
0 7044 7 2 2 65279 67998
0 7045 7 1 2 67997 68002
0 7046 5 1 1 7045
0 7047 7 1 2 7040 7046
0 7048 5 1 1 7047
0 7049 7 1 2 55469 7048
0 7050 5 1 1 7049
0 7051 7 1 2 6999 7050
0 7052 5 1 1 7051
0 7053 7 1 2 67748 7052
0 7054 5 1 1 7053
0 7055 7 2 2 53872 61794
0 7056 5 1 1 68004
0 7057 7 2 2 53157 59634
0 7058 5 2 1 68006
0 7059 7 2 2 52373 68007
0 7060 5 2 1 68010
0 7061 7 1 2 58095 68012
0 7062 5 1 1 7061
0 7063 7 1 2 1080 7062
0 7064 5 1 1 7063
0 7065 7 1 2 48129 7064
0 7066 5 1 1 7065
0 7067 7 1 2 64656 57372
0 7068 5 1 1 7067
0 7069 7 1 2 7066 7068
0 7070 5 1 1 7069
0 7071 7 1 2 48339 7070
0 7072 5 1 1 7071
0 7073 7 1 2 61364 60086
0 7074 5 1 1 7073
0 7075 7 1 2 7072 7074
0 7076 5 1 1 7075
0 7077 7 1 2 61746 7076
0 7078 5 1 1 7077
0 7079 7 4 2 54199 56340
0 7080 5 5 1 68014
0 7081 7 2 2 58096 68015
0 7082 7 1 2 48130 68023
0 7083 5 1 1 7082
0 7084 7 1 2 61432 7083
0 7085 7 1 2 7078 7084
0 7086 5 1 1 7085
0 7087 7 1 2 68005 7086
0 7088 5 1 1 7087
0 7089 7 1 2 53873 56050
0 7090 7 1 2 68024 7089
0 7091 5 1 1 7090
0 7092 7 1 2 56541 57797
0 7093 5 1 1 7092
0 7094 7 2 2 63296 7093
0 7095 7 1 2 52595 68025
0 7096 5 2 1 7095
0 7097 7 3 2 50366 59714
0 7098 5 4 1 68029
0 7099 7 1 2 54897 68032
0 7100 7 1 2 68027 7099
0 7101 5 1 1 7100
0 7102 7 1 2 7091 7101
0 7103 5 1 1 7102
0 7104 7 1 2 61545 7103
0 7105 5 1 1 7104
0 7106 7 2 2 58739 7042
0 7107 5 1 1 68036
0 7108 7 1 2 61667 56607
0 7109 5 4 1 7108
0 7110 7 1 2 7107 68038
0 7111 5 1 1 7110
0 7112 7 2 2 56341 62802
0 7113 5 1 1 68042
0 7114 7 1 2 56542 68043
0 7115 5 1 1 7114
0 7116 7 1 2 59057 7115
0 7117 5 1 1 7116
0 7118 7 1 2 64161 7117
0 7119 5 1 1 7118
0 7120 7 1 2 7111 7119
0 7121 7 1 2 7105 7120
0 7122 7 1 2 7088 7121
0 7123 5 1 1 7122
0 7124 7 1 2 54526 7123
0 7125 5 1 1 7124
0 7126 7 1 2 57423 59060
0 7127 5 1 1 7126
0 7128 7 1 2 61359 7127
0 7129 5 2 1 7128
0 7130 7 2 2 64207 61957
0 7131 5 1 1 68046
0 7132 7 1 2 68044 7131
0 7133 5 1 1 7132
0 7134 7 2 2 56051 59061
0 7135 5 1 1 68048
0 7136 7 2 2 60743 61849
0 7137 5 1 1 68050
0 7138 7 1 2 68049 68051
0 7139 5 1 1 7138
0 7140 7 1 2 61371 7139
0 7141 7 1 2 7133 7140
0 7142 5 1 1 7141
0 7143 7 1 2 54898 7142
0 7144 5 1 1 7143
0 7145 7 1 2 7125 7144
0 7146 5 1 1 7145
0 7147 7 1 2 58847 7146
0 7148 5 1 1 7147
0 7149 7 2 2 60744 60968
0 7150 5 1 1 68052
0 7151 7 1 2 63268 68053
0 7152 5 1 1 7151
0 7153 7 1 2 65366 7152
0 7154 5 1 1 7153
0 7155 7 1 2 54899 7154
0 7156 5 1 1 7155
0 7157 7 1 2 52596 7156
0 7158 5 1 1 7157
0 7159 7 1 2 54527 7158
0 7160 5 1 1 7159
0 7161 7 2 2 58506 62256
0 7162 7 4 2 53874 64700
0 7163 5 2 1 68056
0 7164 7 1 2 65169 68057
0 7165 7 1 2 68054 7164
0 7166 5 1 1 7165
0 7167 7 1 2 7160 7166
0 7168 5 1 1 7167
0 7169 7 1 2 56052 7168
0 7170 5 1 1 7169
0 7171 7 5 2 60907 61655
0 7172 5 5 1 68062
0 7173 7 2 2 60753 68067
0 7174 5 1 1 68072
0 7175 7 1 2 66836 7174
0 7176 5 1 1 7175
0 7177 7 7 2 48131 60908
0 7178 5 1 1 68074
0 7179 7 1 2 65908 68075
0 7180 5 1 1 7179
0 7181 7 1 2 50934 7180
0 7182 5 1 1 7181
0 7183 7 1 2 56838 7182
0 7184 5 1 1 7183
0 7185 7 5 2 53978 60909
0 7186 5 1 1 68081
0 7187 7 1 2 57777 7186
0 7188 5 1 1 7187
0 7189 7 1 2 48132 7188
0 7190 5 1 1 7189
0 7191 7 1 2 59432 62710
0 7192 5 2 1 7191
0 7193 7 1 2 7190 68086
0 7194 5 1 1 7193
0 7195 7 1 2 65532 7194
0 7196 5 1 1 7195
0 7197 7 1 2 7184 7196
0 7198 5 1 1 7197
0 7199 7 1 2 57424 7198
0 7200 5 1 1 7199
0 7201 7 1 2 60910 61816
0 7202 5 1 1 7201
0 7203 7 1 2 61005 7202
0 7204 5 1 1 7203
0 7205 7 2 2 54900 7204
0 7206 5 1 1 68088
0 7207 7 1 2 56839 68089
0 7208 5 1 1 7207
0 7209 7 1 2 48703 63045
0 7210 5 1 1 7209
0 7211 7 1 2 7208 7210
0 7212 7 1 2 7200 7211
0 7213 5 1 1 7212
0 7214 7 1 2 54528 7213
0 7215 5 1 1 7214
0 7216 7 1 2 7176 7215
0 7217 7 1 2 7170 7216
0 7218 5 1 1 7217
0 7219 7 1 2 56543 7218
0 7220 5 1 1 7219
0 7221 7 4 2 64469 59073
0 7222 5 1 1 68090
0 7223 7 1 2 54200 68091
0 7224 5 1 1 7223
0 7225 7 1 2 66947 7224
0 7226 5 1 1 7225
0 7227 7 1 2 54901 7226
0 7228 5 1 1 7227
0 7229 7 1 2 64667 66865
0 7230 5 1 1 7229
0 7231 7 1 2 48133 7230
0 7232 5 1 1 7231
0 7233 7 1 2 64407 61681
0 7234 5 1 1 7233
0 7235 7 1 2 64157 7234
0 7236 7 1 2 7232 7235
0 7237 5 1 1 7236
0 7238 7 1 2 56342 7237
0 7239 5 1 1 7238
0 7240 7 1 2 60940 56608
0 7241 5 6 1 7240
0 7242 7 1 2 65067 68094
0 7243 5 1 1 7242
0 7244 7 1 2 7239 7243
0 7245 7 1 2 7228 7244
0 7246 5 1 1 7245
0 7247 7 1 2 58097 7246
0 7248 5 1 1 7247
0 7249 7 3 2 49104 59542
0 7250 5 3 1 68100
0 7251 7 1 2 63978 68101
0 7252 5 2 1 7251
0 7253 7 1 2 50935 68106
0 7254 5 2 1 7253
0 7255 7 1 2 61365 68108
0 7256 5 1 1 7255
0 7257 7 5 2 52070 60941
0 7258 5 8 1 68110
0 7259 7 4 2 61682 68115
0 7260 5 1 1 68123
0 7261 7 2 2 60745 68124
0 7262 5 1 1 68127
0 7263 7 1 2 61429 68128
0 7264 5 1 1 7263
0 7265 7 1 2 7256 7264
0 7266 5 1 1 7265
0 7267 7 1 2 56053 7266
0 7268 5 1 1 7267
0 7269 7 1 2 48704 68095
0 7270 5 1 1 7269
0 7271 7 1 2 65550 60746
0 7272 5 1 1 7271
0 7273 7 1 2 7270 7272
0 7274 5 1 1 7273
0 7275 7 1 2 54529 7274
0 7276 5 1 1 7275
0 7277 7 3 2 54902 57273
0 7278 5 1 1 68129
0 7279 7 1 2 65119 68130
0 7280 5 1 1 7279
0 7281 7 1 2 7276 7280
0 7282 5 1 1 7281
0 7283 7 1 2 56544 7282
0 7284 5 1 1 7283
0 7285 7 1 2 7268 7284
0 7286 7 1 2 7248 7285
0 7287 5 1 1 7286
0 7288 7 1 2 60689 7287
0 7289 5 1 1 7288
0 7290 7 3 2 50143 60942
0 7291 5 11 1 68132
0 7292 7 1 2 65047 66929
0 7293 5 1 1 7292
0 7294 7 1 2 61366 7293
0 7295 5 1 1 7294
0 7296 7 3 2 48340 59526
0 7297 5 2 1 68146
0 7298 7 1 2 61430 68147
0 7299 5 1 1 7298
0 7300 7 1 2 7295 7299
0 7301 5 1 1 7300
0 7302 7 1 2 56688 7301
0 7303 5 1 1 7302
0 7304 7 1 2 57425 59498
0 7305 5 2 1 7304
0 7306 7 4 2 49189 59077
0 7307 5 1 1 68153
0 7308 7 2 2 60630 68154
0 7309 5 2 1 68157
0 7310 7 1 2 62222 68158
0 7311 5 1 1 7310
0 7312 7 1 2 68151 7311
0 7313 5 1 1 7312
0 7314 7 1 2 57373 7313
0 7315 5 1 1 7314
0 7316 7 2 2 53053 59506
0 7317 5 4 1 68161
0 7318 7 1 2 62424 68162
0 7319 5 1 1 7318
0 7320 7 1 2 59062 7319
0 7321 5 1 1 7320
0 7322 7 1 2 7315 7321
0 7323 5 1 1 7322
0 7324 7 1 2 63440 7323
0 7325 5 1 1 7324
0 7326 7 1 2 7303 7325
0 7327 5 1 1 7326
0 7328 7 1 2 68135 7327
0 7329 5 1 1 7328
0 7330 7 1 2 60911 61890
0 7331 5 1 1 7330
0 7332 7 1 2 50936 7331
0 7333 5 1 1 7332
0 7334 7 1 2 54201 7333
0 7335 5 1 1 7334
0 7336 7 1 2 56689 66718
0 7337 7 1 2 67749 7336
0 7338 5 1 1 7337
0 7339 7 1 2 7335 7338
0 7340 5 1 1 7339
0 7341 7 1 2 56343 7340
0 7342 5 1 1 7341
0 7343 7 1 2 54530 65360
0 7344 5 1 1 7343
0 7345 7 2 2 65426 68076
0 7346 5 3 1 68167
0 7347 7 1 2 7344 68169
0 7348 5 1 1 7347
0 7349 7 1 2 54903 7348
0 7350 5 1 1 7349
0 7351 7 1 2 65078 7350
0 7352 7 1 2 7342 7351
0 7353 5 1 1 7352
0 7354 7 1 2 56054 58098
0 7355 7 1 2 7353 7354
0 7356 5 1 1 7355
0 7357 7 1 2 57139 58940
0 7358 5 2 1 7357
0 7359 7 1 2 7206 68172
0 7360 5 1 1 7359
0 7361 7 1 2 54531 58099
0 7362 7 1 2 7360 7361
0 7363 5 1 1 7362
0 7364 7 9 2 48596 48705
0 7365 5 1 1 68174
0 7366 7 16 2 49533 68175
0 7367 5 1 1 68183
0 7368 7 2 2 59219 58100
0 7369 7 1 2 65048 66932
0 7370 5 1 1 7369
0 7371 7 1 2 68082 7370
0 7372 5 1 1 7371
0 7373 7 2 2 50634 60754
0 7374 5 1 1 68201
0 7375 7 1 2 54904 7374
0 7376 5 1 1 7375
0 7377 7 1 2 7372 7376
0 7378 5 1 1 7377
0 7379 7 1 2 68199 7378
0 7380 5 1 1 7379
0 7381 7 1 2 7367 7380
0 7382 7 1 2 7363 7381
0 7383 7 1 2 7356 7382
0 7384 7 1 2 7329 7383
0 7385 7 1 2 7289 7384
0 7386 7 1 2 7220 7385
0 7387 7 1 2 7148 7386
0 7388 5 1 1 7387
0 7389 7 1 2 55470 68003
0 7390 7 1 2 7388 7389
0 7391 5 1 1 7390
0 7392 7 1 2 7054 7391
0 7393 7 1 2 6946 7392
0 7394 5 1 1 7393
0 7395 7 11 2 52853 53765
0 7396 5 11 1 68203
0 7397 7 49 2 48984 49992
0 7398 5 3 1 68225
0 7399 7 4 2 68214 68274
0 7400 5 1 1 68277
0 7401 7 1 2 7394 68278
0 7402 5 1 1 7401
0 7403 7 2 2 65157 66957
0 7404 5 4 1 68281
0 7405 7 1 2 66318 68283
0 7406 5 1 1 7405
0 7407 7 1 2 52760 7406
0 7408 5 2 1 7407
0 7409 7 9 2 54202 50937
0 7410 7 2 2 56840 68289
0 7411 7 1 2 66842 68298
0 7412 5 1 1 7411
0 7413 7 2 2 51227 64701
0 7414 5 1 1 68300
0 7415 7 1 2 58101 68301
0 7416 5 1 1 7415
0 7417 7 1 2 7412 7416
0 7418 5 1 1 7417
0 7419 7 15 2 53427 54532
0 7420 7 1 2 51497 68302
0 7421 7 1 2 7418 7420
0 7422 5 1 1 7421
0 7423 7 1 2 68287 7422
0 7424 5 1 1 7423
0 7425 7 1 2 55596 7424
0 7426 5 1 1 7425
0 7427 7 8 2 63007 67906
0 7428 5 3 1 68317
0 7429 7 1 2 64702 66843
0 7430 7 1 2 68318 7429
0 7431 5 1 1 7430
0 7432 7 1 2 7426 7431
0 7433 5 1 1 7432
0 7434 7 1 2 53639 7433
0 7435 5 1 1 7434
0 7436 7 7 2 63777 66288
0 7437 5 3 1 68328
0 7438 7 1 2 64717 67760
0 7439 5 1 1 7438
0 7440 7 1 2 68335 7439
0 7441 5 1 1 7440
0 7442 7 1 2 56841 7441
0 7443 5 1 1 7442
0 7444 7 14 2 49837 53979
0 7445 7 2 2 65968 68338
0 7446 5 1 1 68352
0 7447 7 1 2 54203 68353
0 7448 5 1 1 7447
0 7449 7 1 2 7443 7448
0 7450 5 1 1 7449
0 7451 7 1 2 62537 7450
0 7452 5 1 1 7451
0 7453 7 6 2 54204 66066
0 7454 5 1 1 68354
0 7455 7 1 2 67482 7454
0 7456 5 1 1 7455
0 7457 7 1 2 47839 7456
0 7458 5 1 1 7457
0 7459 7 1 2 66267 66697
0 7460 5 1 1 7459
0 7461 7 1 2 7458 7460
0 7462 5 1 1 7461
0 7463 7 1 2 54533 7462
0 7464 5 1 1 7463
0 7465 7 1 2 67796 7464
0 7466 5 1 1 7465
0 7467 7 1 2 62892 7466
0 7468 5 1 1 7467
0 7469 7 1 2 7452 7468
0 7470 5 1 1 7469
0 7471 7 1 2 57885 7470
0 7472 5 1 1 7471
0 7473 7 1 2 67510 68329
0 7474 5 2 1 7473
0 7475 7 5 2 50938 66408
0 7476 7 1 2 62654 68362
0 7477 5 4 1 7476
0 7478 7 2 2 53428 66409
0 7479 5 2 1 68371
0 7480 7 1 2 62893 66443
0 7481 5 1 1 7480
0 7482 7 1 2 68373 7481
0 7483 5 1 1 7482
0 7484 7 1 2 64506 7483
0 7485 5 1 1 7484
0 7486 7 1 2 64783 66984
0 7487 5 1 1 7486
0 7488 7 1 2 7485 7487
0 7489 5 1 1 7488
0 7490 7 1 2 53980 7489
0 7491 5 1 1 7490
0 7492 7 1 2 68367 7491
0 7493 5 1 1 7492
0 7494 7 1 2 49838 7493
0 7495 5 1 1 7494
0 7496 7 1 2 68360 7495
0 7497 7 1 2 7472 7496
0 7498 5 1 1 7497
0 7499 7 1 2 51685 7498
0 7500 5 1 1 7499
0 7501 7 1 2 7435 7500
0 7502 5 1 1 7501
0 7503 7 1 2 58376 7502
0 7504 5 1 1 7503
0 7505 7 1 2 66319 67194
0 7506 5 1 1 7505
0 7507 7 1 2 52761 7506
0 7508 5 1 1 7507
0 7509 7 34 2 50939 55240
0 7510 5 2 1 68375
0 7511 7 3 2 56842 68376
0 7512 5 1 1 68411
0 7513 7 1 2 62711 68412
0 7514 5 1 1 7513
0 7515 7 2 2 51228 58102
0 7516 7 1 2 54905 68414
0 7517 5 1 1 7516
0 7518 7 1 2 7514 7517
0 7519 5 1 1 7518
0 7520 7 2 2 66518 7519
0 7521 7 1 2 53429 68416
0 7522 5 1 1 7521
0 7523 7 1 2 7508 7522
0 7524 5 1 1 7523
0 7525 7 1 2 55597 7524
0 7526 5 1 1 7525
0 7527 7 2 2 59976 63008
0 7528 7 1 2 63823 67907
0 7529 7 1 2 68418 7528
0 7530 5 1 1 7529
0 7531 7 1 2 7526 7530
0 7532 5 1 1 7531
0 7533 7 1 2 53640 7532
0 7534 5 1 1 7533
0 7535 7 1 2 62894 66365
0 7536 5 2 1 7535
0 7537 7 2 2 68420 68368
0 7538 5 2 1 68422
0 7539 7 6 2 51498 67991
0 7540 5 1 1 68426
0 7541 7 1 2 56843 68427
0 7542 5 1 1 7541
0 7543 7 1 2 68374 7542
0 7544 5 1 1 7543
0 7545 7 1 2 64106 7544
0 7546 5 1 1 7545
0 7547 7 1 2 68423 7546
0 7548 5 1 1 7547
0 7549 7 1 2 49839 7548
0 7550 5 1 1 7549
0 7551 7 1 2 58799 66289
0 7552 5 2 1 7551
0 7553 7 4 2 50635 66290
0 7554 5 4 1 68434
0 7555 7 1 2 67195 68438
0 7556 5 1 1 7555
0 7557 7 1 2 48706 7556
0 7558 5 1 1 7557
0 7559 7 1 2 68432 7558
0 7560 5 1 1 7559
0 7561 7 1 2 65695 7560
0 7562 5 1 1 7561
0 7563 7 4 2 61891 66067
0 7564 7 1 2 67669 68442
0 7565 5 1 1 7564
0 7566 7 1 2 7562 7565
0 7567 5 1 1 7566
0 7568 7 1 2 57886 7567
0 7569 5 1 1 7568
0 7570 7 1 2 68361 7569
0 7571 7 1 2 7550 7570
0 7572 5 1 1 7571
0 7573 7 1 2 51686 7572
0 7574 5 1 1 7573
0 7575 7 1 2 7534 7574
0 7576 5 1 1 7575
0 7577 7 1 2 54205 7576
0 7578 5 1 1 7577
0 7579 7 26 2 51499 55598
0 7580 7 3 2 54906 68446
0 7581 7 7 2 53641 50367
0 7582 7 3 2 53430 68475
0 7583 7 1 2 68472 68482
0 7584 5 2 1 7583
0 7585 7 4 2 53642 62942
0 7586 5 15 1 68487
0 7587 7 2 2 63002 68488
0 7588 5 7 1 68506
0 7589 7 2 2 50940 68508
0 7590 7 1 2 53981 67908
0 7591 7 1 2 68515 7590
0 7592 5 1 1 7591
0 7593 7 1 2 68485 7592
0 7594 5 1 1 7593
0 7595 7 1 2 65696 7594
0 7596 5 1 1 7595
0 7597 7 15 2 51229 55599
0 7598 7 3 2 66291 68517
0 7599 7 2 2 52762 66578
0 7600 7 1 2 68532 68535
0 7601 5 1 1 7600
0 7602 7 1 2 7596 7601
0 7603 5 1 1 7602
0 7604 7 1 2 50636 7603
0 7605 5 1 1 7604
0 7606 7 1 2 64586 68419
0 7607 5 1 1 7606
0 7608 7 1 2 62823 67652
0 7609 5 1 1 7608
0 7610 7 1 2 7607 7609
0 7611 5 1 1 7610
0 7612 7 1 2 67761 7611
0 7613 5 1 1 7612
0 7614 7 2 2 63566 66068
0 7615 5 2 1 68537
0 7616 7 1 2 62824 68538
0 7617 5 1 1 7616
0 7618 7 1 2 7613 7617
0 7619 5 1 1 7618
0 7620 7 1 2 51687 7619
0 7621 5 1 1 7620
0 7622 7 1 2 7605 7621
0 7623 7 1 2 7578 7622
0 7624 7 1 2 7504 7623
0 7625 5 1 1 7624
0 7626 7 1 2 57140 7625
0 7627 5 1 1 7626
0 7628 7 13 2 53643 55600
0 7629 7 4 2 51500 63441
0 7630 7 1 2 63401 68554
0 7631 5 2 1 7630
0 7632 7 1 2 4666 68558
0 7633 5 1 1 7632
0 7634 7 1 2 52763 7633
0 7635 5 2 1 7634
0 7636 7 1 2 63325 68417
0 7637 5 1 1 7636
0 7638 7 1 2 68560 7637
0 7639 5 1 1 7638
0 7640 7 1 2 68541 7639
0 7641 5 1 1 7640
0 7642 7 2 2 49840 65969
0 7643 5 4 1 68562
0 7644 7 32 2 49683 51230
0 7645 5 10 1 68568
0 7646 7 8 2 54206 55471
0 7647 7 4 2 53982 68610
0 7648 7 1 2 68569 68618
0 7649 5 1 1 7648
0 7650 7 1 2 68564 7649
0 7651 5 1 1 7650
0 7652 7 1 2 47840 7651
0 7653 5 1 1 7652
0 7654 7 3 2 64137 65970
0 7655 7 2 2 48498 66527
0 7656 7 1 2 68622 68625
0 7657 5 1 1 7656
0 7658 7 1 2 7653 7657
0 7659 5 1 1 7658
0 7660 7 1 2 54534 7659
0 7661 5 1 1 7660
0 7662 7 5 2 49684 67762
0 7663 5 2 1 68627
0 7664 7 1 2 68632 68369
0 7665 5 1 1 7664
0 7666 7 1 2 53983 7665
0 7667 5 1 1 7666
0 7668 7 1 2 7661 7667
0 7669 5 1 1 7668
0 7670 7 1 2 48707 7669
0 7671 5 1 1 7670
0 7672 7 2 2 66698 68435
0 7673 5 1 1 68634
0 7674 7 3 2 47841 67763
0 7675 5 1 1 68636
0 7676 7 1 2 54535 68637
0 7677 5 1 1 7676
0 7678 7 1 2 7673 7677
0 7679 5 1 1 7678
0 7680 7 1 2 67674 7679
0 7681 5 1 1 7680
0 7682 7 1 2 7671 7681
0 7683 5 1 1 7682
0 7684 7 1 2 57887 7683
0 7685 5 1 1 7684
0 7686 7 1 2 68491 68635
0 7687 5 1 1 7686
0 7688 7 5 2 49841 54536
0 7689 7 2 2 66958 66998
0 7690 5 2 1 68644
0 7691 7 1 2 68639 68645
0 7692 5 1 1 7691
0 7693 7 1 2 7687 7692
0 7694 5 1 1 7693
0 7695 7 1 2 55241 7694
0 7696 5 1 1 7695
0 7697 7 1 2 7685 7696
0 7698 5 1 1 7697
0 7699 7 1 2 51688 7698
0 7700 5 1 1 7699
0 7701 7 1 2 7641 7700
0 7702 5 1 1 7701
0 7703 7 1 2 58377 7702
0 7704 5 1 1 7703
0 7705 7 1 2 64625 64962
0 7706 7 1 2 68184 7705
0 7707 5 1 1 7706
0 7708 7 2 2 55242 63884
0 7709 5 1 1 68648
0 7710 7 1 2 64904 7709
0 7711 5 2 1 7710
0 7712 7 1 2 49842 58103
0 7713 7 1 2 68650 7712
0 7714 5 1 1 7713
0 7715 7 1 2 7707 7714
0 7716 5 1 1 7715
0 7717 7 1 2 51689 7716
0 7718 5 1 1 7717
0 7719 7 4 2 55601 64138
0 7720 7 1 2 68652 68536
0 7721 5 1 1 7720
0 7722 7 1 2 7718 7721
0 7723 5 1 1 7722
0 7724 7 1 2 54537 7723
0 7725 5 1 1 7724
0 7726 7 15 2 52764 55243
0 7727 5 2 1 68656
0 7728 7 1 2 68657 68542
0 7729 5 2 1 7728
0 7730 7 1 2 7725 68673
0 7731 5 1 1 7730
0 7732 7 1 2 49685 7731
0 7733 5 1 1 7732
0 7734 7 2 2 49534 49843
0 7735 7 4 2 68176 68675
0 7736 7 5 2 54538 51690
0 7737 7 1 2 68677 68681
0 7738 7 1 2 68651 7737
0 7739 5 1 1 7738
0 7740 7 21 2 54539 51231
0 7741 5 1 1 68686
0 7742 7 5 2 60379 68687
0 7743 5 1 1 68707
0 7744 7 1 2 54907 7743
0 7745 5 1 1 7744
0 7746 7 1 2 4933 68543
0 7747 7 1 2 59115 7746
0 7748 7 1 2 7745 7747
0 7749 5 1 1 7748
0 7750 7 1 2 7739 7749
0 7751 7 1 2 7733 7750
0 7752 5 1 1 7751
0 7753 7 1 2 51501 7752
0 7754 5 1 1 7753
0 7755 7 8 2 53644 50637
0 7756 7 3 2 52765 68712
0 7757 7 1 2 68720 68533
0 7758 5 3 1 7757
0 7759 7 1 2 49844 68424
0 7760 5 1 1 7759
0 7761 7 2 2 56844 63778
0 7762 7 1 2 66292 68726
0 7763 7 1 2 63009 7762
0 7764 5 1 1 7763
0 7765 7 1 2 7760 7764
0 7766 5 1 1 7765
0 7767 7 1 2 51691 7766
0 7768 5 1 1 7767
0 7769 7 1 2 68723 7768
0 7770 5 1 1 7769
0 7771 7 1 2 54207 7770
0 7772 5 1 1 7771
0 7773 7 4 2 49686 66069
0 7774 5 2 1 68728
0 7775 7 3 2 62825 68729
0 7776 5 1 1 68734
0 7777 7 3 2 63010 67693
0 7778 5 3 1 68737
0 7779 7 1 2 49845 65333
0 7780 7 1 2 68738 7779
0 7781 5 1 1 7780
0 7782 7 1 2 7776 7781
0 7783 5 1 1 7782
0 7784 7 1 2 51692 7783
0 7785 5 1 1 7784
0 7786 7 14 2 53431 53645
0 7787 5 1 1 68743
0 7788 7 3 2 56845 68744
0 7789 7 5 2 60525 68447
0 7790 7 1 2 68757 68760
0 7791 5 1 1 7790
0 7792 7 12 2 49687 49846
0 7793 5 2 1 68765
0 7794 7 3 2 68777 68509
0 7795 7 1 2 64069 67909
0 7796 7 1 2 68779 7795
0 7797 5 1 1 7796
0 7798 7 1 2 7791 7797
0 7799 5 1 1 7798
0 7800 7 1 2 55244 7799
0 7801 5 1 1 7800
0 7802 7 1 2 7785 7801
0 7803 5 1 1 7802
0 7804 7 1 2 54908 7803
0 7805 5 1 1 7804
0 7806 7 1 2 7772 7805
0 7807 5 1 1 7806
0 7808 7 1 2 59977 7807
0 7809 5 1 1 7808
0 7810 7 3 2 56846 68570
0 7811 5 2 1 68782
0 7812 7 2 2 63442 66463
0 7813 5 1 1 68787
0 7814 7 1 2 68785 7813
0 7815 5 1 1 7814
0 7816 7 1 2 48708 7815
0 7817 5 1 1 7816
0 7818 7 3 2 66464 66372
0 7819 5 5 1 68789
0 7820 7 1 2 54909 68790
0 7821 5 1 1 7820
0 7822 7 1 2 7817 7821
0 7823 5 1 1 7822
0 7824 7 1 2 57888 7823
0 7825 5 1 1 7824
0 7826 7 18 2 53432 49847
0 7827 5 3 1 68797
0 7828 7 19 2 49688 53646
0 7829 5 4 1 68818
0 7830 7 5 2 48709 68819
0 7831 5 2 1 68841
0 7832 7 3 2 68815 68846
0 7833 5 2 1 68848
0 7834 7 1 2 63856 68851
0 7835 5 1 1 7834
0 7836 7 1 2 7825 7835
0 7837 5 1 1 7836
0 7838 7 1 2 67910 7837
0 7839 5 1 1 7838
0 7840 7 1 2 7809 7839
0 7841 7 1 2 7754 7840
0 7842 7 1 2 7704 7841
0 7843 5 1 1 7842
0 7844 7 1 2 56690 7843
0 7845 5 1 1 7844
0 7846 7 3 2 53647 51502
0 7847 7 8 2 55602 68853
0 7848 7 2 2 60912 56691
0 7849 7 1 2 53875 68864
0 7850 5 3 1 7849
0 7851 7 1 2 60755 67302
0 7852 7 1 2 68866 7851
0 7853 5 1 1 7852
0 7854 7 1 2 67560 7853
0 7855 5 1 1 7854
0 7856 7 15 2 50368 54910
0 7857 7 5 2 50144 68869
0 7858 5 1 1 68884
0 7859 7 1 2 60959 68885
0 7860 5 1 1 7859
0 7861 7 1 2 7855 7860
0 7862 5 1 1 7861
0 7863 7 1 2 68856 7862
0 7864 5 1 1 7863
0 7865 7 19 2 51693 67822
0 7866 5 2 1 68889
0 7867 7 1 2 59543 65909
0 7868 5 1 1 7867
0 7869 7 1 2 50941 7868
0 7870 5 1 1 7869
0 7871 7 1 2 68890 7870
0 7872 5 1 1 7871
0 7873 7 1 2 7864 7872
0 7874 5 1 1 7873
0 7875 7 1 2 54540 7874
0 7876 5 1 1 7875
0 7877 7 1 2 56692 64107
0 7878 5 1 1 7877
0 7879 7 2 2 48134 64661
0 7880 5 2 1 68910
0 7881 7 1 2 65367 68912
0 7882 7 1 2 7878 7881
0 7883 5 1 1 7882
0 7884 7 1 2 68891 7883
0 7885 5 1 1 7884
0 7886 7 26 2 50638 54911
0 7887 5 1 1 68914
0 7888 7 3 2 61656 68290
0 7889 7 1 2 66175 68940
0 7890 5 1 1 7889
0 7891 7 1 2 7887 7890
0 7892 5 1 1 7891
0 7893 7 6 2 55603 56847
0 7894 7 1 2 68854 68943
0 7895 7 1 2 7892 7894
0 7896 5 1 1 7895
0 7897 7 1 2 7885 7896
0 7898 7 1 2 7876 7897
0 7899 5 1 1 7898
0 7900 7 1 2 51232 7899
0 7901 5 1 1 7900
0 7902 7 8 2 49848 54208
0 7903 7 9 2 55245 51694
0 7904 7 3 2 54912 68957
0 7905 7 2 2 66444 68966
0 7906 7 1 2 68949 68969
0 7907 5 1 1 7906
0 7908 7 11 2 53648 50942
0 7909 7 6 2 55604 68971
0 7910 7 2 2 66445 68982
0 7911 5 1 1 68988
0 7912 7 3 2 49849 53876
0 7913 7 6 2 49105 68990
0 7914 7 5 2 51695 68611
0 7915 7 1 2 68993 68999
0 7916 5 1 1 7915
0 7917 7 1 2 7911 7916
0 7918 5 1 1 7917
0 7919 7 1 2 47842 51233
0 7920 7 1 2 7918 7919
0 7921 5 1 1 7920
0 7922 7 1 2 7907 7921
0 7923 5 1 1 7922
0 7924 7 1 2 61835 7923
0 7925 5 1 1 7924
0 7926 7 3 2 57141 59978
0 7927 5 1 1 69004
0 7928 7 1 2 60756 7927
0 7929 5 1 1 7928
0 7930 7 3 2 54913 58378
0 7931 5 1 1 69007
0 7932 7 2 2 56848 69008
0 7933 5 1 1 69010
0 7934 7 1 2 51503 67999
0 7935 7 1 2 69011 7934
0 7936 7 1 2 7929 7935
0 7937 5 1 1 7936
0 7938 7 1 2 7925 7937
0 7939 5 1 1 7938
0 7940 7 1 2 54541 7939
0 7941 5 1 1 7940
0 7942 7 1 2 7901 7941
0 7943 5 1 1 7942
0 7944 7 1 2 58962 7943
0 7945 5 1 1 7944
0 7946 7 8 2 55605 68745
0 7947 7 1 2 69012 68291
0 7948 5 1 1 7947
0 7949 7 11 2 49850 51696
0 7950 7 4 2 49689 69020
0 7951 5 1 1 69031
0 7952 7 1 2 54914 69032
0 7953 5 1 1 7952
0 7954 7 1 2 7948 7953
0 7955 5 1 1 7954
0 7956 7 1 2 58104 7955
0 7957 5 1 1 7956
0 7958 7 2 2 54209 55606
0 7959 7 4 2 53649 58999
0 7960 7 1 2 69035 69037
0 7961 5 1 1 7960
0 7962 7 7 2 54915 51697
0 7963 7 1 2 68678 69041
0 7964 5 1 1 7963
0 7965 7 1 2 7961 7964
0 7966 7 1 2 7957 7965
0 7967 5 1 1 7966
0 7968 7 1 2 65971 7967
0 7969 5 1 1 7968
0 7970 7 5 2 51698 57889
0 7971 7 3 2 67490 69048
0 7972 7 3 2 51234 63443
0 7973 7 1 2 69053 69056
0 7974 5 1 1 7973
0 7975 7 2 2 66814 68448
0 7976 7 2 2 52766 63824
0 7977 7 1 2 69059 69061
0 7978 5 2 1 7977
0 7979 7 1 2 67550 69054
0 7980 5 1 1 7979
0 7981 7 1 2 69063 7980
0 7982 5 1 1 7981
0 7983 7 1 2 56849 7982
0 7984 5 1 1 7983
0 7985 7 1 2 7974 7984
0 7986 7 1 2 7969 7985
0 7987 7 1 2 7945 7986
0 7988 7 1 2 7845 7987
0 7989 7 1 2 7627 7988
0 7990 5 1 1 7989
0 7991 7 1 2 68226 7990
0 7992 5 1 1 7991
0 7993 7 4 2 54210 51699
0 7994 7 3 2 48985 69065
0 7995 5 1 1 69069
0 7996 7 23 2 48986 51700
0 7997 5 1 1 69072
0 7998 7 1 2 63933 69073
0 7999 5 1 1 7998
0 8000 7 2 2 49106 68758
0 8001 7 1 2 55607 68941
0 8002 7 1 2 69095 8001
0 8003 5 1 1 8002
0 8004 7 1 2 7999 8003
0 8005 5 1 1 8004
0 8006 7 1 2 47843 8005
0 8007 5 1 1 8006
0 8008 7 1 2 7995 8007
0 8009 5 1 1 8008
0 8010 7 1 2 51504 8009
0 8011 5 1 1 8010
0 8012 7 9 2 49851 54916
0 8013 5 1 1 69097
0 8014 7 6 2 67911 69098
0 8015 5 4 1 69106
0 8016 7 1 2 53433 69107
0 8017 5 1 1 8016
0 8018 7 1 2 8011 8017
0 8019 5 1 1 8018
0 8020 7 1 2 48710 8019
0 8021 5 1 1 8020
0 8022 7 4 2 51505 51701
0 8023 7 2 2 48987 69116
0 8024 7 6 2 47844 49690
0 8025 5 2 1 69122
0 8026 7 1 2 65519 69128
0 8027 5 2 1 8026
0 8028 7 1 2 63934 69130
0 8029 5 1 1 8028
0 8030 7 1 2 63408 8029
0 8031 5 2 1 8030
0 8032 7 1 2 69120 69132
0 8033 5 1 1 8032
0 8034 7 1 2 8021 8033
0 8035 5 1 1 8034
0 8036 7 1 2 57890 8035
0 8037 5 1 1 8036
0 8038 7 1 2 54211 68492
0 8039 5 2 1 8038
0 8040 7 1 2 47845 68493
0 8041 5 1 1 8040
0 8042 7 1 2 64139 63163
0 8043 5 1 1 8042
0 8044 7 1 2 8041 8043
0 8045 5 1 1 8044
0 8046 7 1 2 63935 8045
0 8047 5 1 1 8046
0 8048 7 1 2 69134 8047
0 8049 5 1 1 8048
0 8050 7 1 2 51506 8049
0 8051 5 1 1 8050
0 8052 7 1 2 67649 8051
0 8053 5 1 1 8052
0 8054 7 1 2 69074 8053
0 8055 5 1 1 8054
0 8056 7 1 2 49993 8055
0 8057 7 1 2 8037 8056
0 8058 5 1 1 8057
0 8059 7 2 2 47846 65329
0 8060 7 1 2 66150 68449
0 8061 7 1 2 69136 8060
0 8062 5 1 1 8061
0 8063 7 1 2 69112 8062
0 8064 5 1 1 8063
0 8065 7 1 2 48988 8064
0 8066 5 1 1 8065
0 8067 7 6 2 55472 55608
0 8068 7 8 2 52854 49852
0 8069 7 2 2 69138 69144
0 8070 7 1 2 69133 69152
0 8071 5 1 1 8070
0 8072 7 1 2 8066 8071
0 8073 5 1 1 8072
0 8074 7 1 2 68185 8073
0 8075 5 1 1 8074
0 8076 7 4 2 54212 63936
0 8077 5 3 1 69154
0 8078 7 1 2 55609 67610
0 8079 7 2 2 66528 8078
0 8080 7 1 2 62294 69145
0 8081 7 2 2 69161 8080
0 8082 7 1 2 69155 69163
0 8083 5 1 1 8082
0 8084 7 1 2 53766 8083
0 8085 7 1 2 8075 8084
0 8086 5 1 1 8085
0 8087 7 1 2 55246 8086
0 8088 7 1 2 8058 8087
0 8089 5 1 1 8088
0 8090 7 6 2 49994 51702
0 8091 7 8 2 48989 51507
0 8092 7 4 2 69171 68510
0 8093 7 1 2 69165 69179
0 8094 5 1 1 8093
0 8095 7 7 2 53767 55473
0 8096 5 1 1 69183
0 8097 7 3 2 52855 68766
0 8098 7 2 2 69184 69190
0 8099 7 3 2 55610 69193
0 8100 5 1 1 69195
0 8101 7 1 2 62826 69196
0 8102 5 1 1 8101
0 8103 7 1 2 8094 8102
0 8104 5 6 1 8103
0 8105 7 1 2 67055 69198
0 8106 5 1 1 8105
0 8107 7 5 2 51235 68227
0 8108 7 2 2 58963 69204
0 8109 7 6 2 67912 69209
0 8110 5 1 1 69211
0 8111 7 1 2 64080 69212
0 8112 5 1 1 8111
0 8113 7 1 2 8106 8112
0 8114 7 1 2 8089 8113
0 8115 5 1 1 8114
0 8116 7 1 2 54542 8115
0 8117 5 1 1 8116
0 8118 7 3 2 50639 55611
0 8119 7 1 2 55247 69217
0 8120 7 1 2 68483 8119
0 8121 5 2 1 8120
0 8122 7 1 2 64070 69075
0 8123 5 1 1 8122
0 8124 7 1 2 69220 8123
0 8125 5 1 1 8124
0 8126 7 1 2 66446 8125
0 8127 5 1 1 8126
0 8128 7 2 2 64784 67913
0 8129 7 1 2 53434 68994
0 8130 7 1 2 69222 8129
0 8131 5 1 1 8130
0 8132 7 1 2 8127 8131
0 8133 5 1 1 8132
0 8134 7 1 2 48711 8133
0 8135 5 1 1 8134
0 8136 7 2 2 64871 62286
0 8137 7 1 2 66959 69224
0 8138 5 1 1 8137
0 8139 7 1 2 66110 8138
0 8140 5 1 1 8139
0 8141 7 1 2 69076 8140
0 8142 5 1 1 8141
0 8143 7 1 2 8135 8142
0 8144 5 1 1 8143
0 8145 7 1 2 57891 8144
0 8146 5 1 1 8145
0 8147 7 3 2 62538 66070
0 8148 5 2 1 69226
0 8149 7 2 2 66447 68494
0 8150 5 1 1 69231
0 8151 7 1 2 66436 8150
0 8152 5 3 1 8151
0 8153 7 1 2 59511 69233
0 8154 5 1 1 8153
0 8155 7 1 2 69229 8154
0 8156 5 1 1 8155
0 8157 7 1 2 69077 8156
0 8158 5 1 1 8157
0 8159 7 1 2 8146 8158
0 8160 5 1 1 8159
0 8161 7 1 2 54917 8160
0 8162 5 1 1 8161
0 8163 7 3 2 49853 62539
0 8164 5 7 1 69236
0 8165 7 2 2 57892 68495
0 8166 5 1 1 69246
0 8167 7 1 2 69239 8166
0 8168 5 1 1 8167
0 8169 7 2 2 51508 8168
0 8170 5 3 1 69248
0 8171 7 1 2 69250 68370
0 8172 5 4 1 8171
0 8173 7 1 2 69070 69253
0 8174 5 1 1 8173
0 8175 7 1 2 8162 8174
0 8176 5 1 1 8175
0 8177 7 1 2 49995 8176
0 8178 5 1 1 8177
0 8179 7 2 2 48990 65972
0 8180 5 1 1 69257
0 8181 7 1 2 55474 64071
0 8182 7 1 2 69191 8181
0 8183 5 1 1 8182
0 8184 7 1 2 8180 8183
0 8185 5 1 1 8184
0 8186 7 1 2 68944 8185
0 8187 5 1 1 8186
0 8188 7 1 2 48991 68995
0 8189 7 1 2 69223 8188
0 8190 5 1 1 8189
0 8191 7 1 2 8187 8190
0 8192 5 1 1 8191
0 8193 7 1 2 53768 64195
0 8194 7 1 2 68177 8193
0 8195 7 1 2 8192 8194
0 8196 5 1 1 8195
0 8197 7 1 2 8178 8196
0 8198 5 1 1 8197
0 8199 7 1 2 59979 8198
0 8200 5 1 1 8199
0 8201 7 11 2 51703 68228
0 8202 7 8 2 51236 58964
0 8203 7 1 2 66536 69270
0 8204 5 2 1 8203
0 8205 7 1 2 61933 69254
0 8206 5 1 1 8205
0 8207 7 1 2 69278 8206
0 8208 5 1 1 8207
0 8209 7 1 2 69259 8208
0 8210 5 1 1 8209
0 8211 7 1 2 8200 8210
0 8212 7 1 2 8117 8211
0 8213 5 1 1 8212
0 8214 7 1 2 56693 8213
0 8215 5 1 1 8214
0 8216 7 1 2 65539 69213
0 8217 5 1 1 8216
0 8218 7 1 2 55248 69199
0 8219 5 1 1 8218
0 8220 7 1 2 67009 69260
0 8221 7 1 2 69271 8220
0 8222 5 1 1 8221
0 8223 7 1 2 8219 8222
0 8224 5 1 1 8223
0 8225 7 1 2 54918 8224
0 8226 5 1 1 8225
0 8227 7 1 2 8217 8226
0 8228 7 1 2 8215 8227
0 8229 7 2 2 68950 68967
0 8230 5 2 1 69280
0 8231 7 1 2 68996 68968
0 8232 5 1 1 8231
0 8233 7 1 2 51237 68983
0 8234 5 1 1 8233
0 8235 7 1 2 8232 8234
0 8236 5 1 1 8235
0 8237 7 1 2 59980 8236
0 8238 5 1 1 8237
0 8239 7 1 2 69282 8238
0 8240 5 1 1 8239
0 8241 7 1 2 54543 8240
0 8242 5 1 1 8241
0 8243 7 8 2 53650 51238
0 8244 7 4 2 49107 55612
0 8245 7 2 2 69284 69292
0 8246 7 1 2 68942 69296
0 8247 5 1 1 8246
0 8248 7 1 2 8242 8247
0 8249 5 1 1 8248
0 8250 7 1 2 66960 8249
0 8251 5 1 1 8250
0 8252 7 7 2 55249 67914
0 8253 7 10 2 49854 50640
0 8254 7 3 2 50943 69305
0 8255 7 5 2 69298 69315
0 8256 7 1 2 58421 60185
0 8257 5 4 1 8256
0 8258 7 1 2 69318 69323
0 8259 5 1 1 8258
0 8260 7 1 2 8251 8259
0 8261 5 1 1 8260
0 8262 7 1 2 56850 8261
0 8263 5 1 1 8262
0 8264 7 2 2 67915 68951
0 8265 5 2 1 69327
0 8266 7 6 2 66759 68450
0 8267 7 1 2 60186 69331
0 8268 5 1 1 8267
0 8269 7 2 2 69329 8268
0 8270 5 3 1 69337
0 8271 7 1 2 58379 69339
0 8272 5 1 1 8271
0 8273 7 17 2 49855 67916
0 8274 5 3 1 69342
0 8275 7 1 2 60380 69343
0 8276 5 1 1 8275
0 8277 7 1 2 8272 8276
0 8278 5 1 1 8277
0 8279 7 1 2 57734 8278
0 8280 5 1 1 8279
0 8281 7 1 2 69113 8280
0 8282 5 1 1 8281
0 8283 7 1 2 68571 8282
0 8284 5 1 1 8283
0 8285 7 1 2 8263 8284
0 8286 5 1 1 8285
0 8287 7 1 2 57142 8286
0 8288 5 1 1 8287
0 8289 7 6 2 50944 68518
0 8290 7 1 2 67542 69362
0 8291 5 1 1 8290
0 8292 7 1 2 69283 8291
0 8293 5 1 1 8292
0 8294 7 1 2 63937 8293
0 8295 5 1 1 8294
0 8296 7 2 2 66738 69363
0 8297 5 1 1 69368
0 8298 7 1 2 8295 8297
0 8299 5 1 1 8298
0 8300 7 1 2 66519 8299
0 8301 5 1 1 8300
0 8302 7 1 2 51239 68892
0 8303 5 1 1 8302
0 8304 7 1 2 8301 8303
0 8305 5 1 1 8304
0 8306 7 1 2 49691 8305
0 8307 5 1 1 8306
0 8308 7 1 2 64088 69319
0 8309 5 1 1 8308
0 8310 7 1 2 8307 8309
0 8311 5 1 1 8310
0 8312 7 1 2 56851 8311
0 8313 5 1 1 8312
0 8314 7 3 2 68730 69021
0 8315 5 2 1 69370
0 8316 7 1 2 65028 61892
0 8317 5 1 1 8316
0 8318 7 1 2 64109 8317
0 8319 5 1 1 8318
0 8320 7 1 2 69371 8319
0 8321 5 1 1 8320
0 8322 7 1 2 8313 8321
0 8323 5 1 1 8322
0 8324 7 1 2 56694 8323
0 8325 5 1 1 8324
0 8326 7 7 2 68451 68713
0 8327 7 2 2 54919 69375
0 8328 5 3 1 69382
0 8329 7 1 2 69330 69384
0 8330 5 3 1 8329
0 8331 7 1 2 56852 69387
0 8332 5 1 1 8331
0 8333 7 1 2 63444 68893
0 8334 5 1 1 8333
0 8335 7 1 2 8332 8334
0 8336 5 1 1 8335
0 8337 7 1 2 68572 8336
0 8338 5 1 1 8337
0 8339 7 1 2 8325 8338
0 8340 7 1 2 8288 8339
0 8341 5 1 1 8340
0 8342 7 1 2 68186 8341
0 8343 5 1 1 8342
0 8344 7 1 2 57143 69324
0 8345 5 2 1 8344
0 8346 7 5 2 56695 64089
0 8347 5 2 1 69392
0 8348 7 1 2 69390 69397
0 8349 5 1 1 8348
0 8350 7 3 2 58105 68626
0 8351 7 1 2 69399 69320
0 8352 7 1 2 8349 8351
0 8353 5 1 1 8352
0 8354 7 1 2 8343 8353
0 8355 5 1 1 8354
0 8356 7 1 2 68215 8355
0 8357 5 1 1 8356
0 8358 7 2 2 69185 69146
0 8359 7 1 2 53435 7933
0 8360 5 1 1 8359
0 8361 7 1 2 59981 8360
0 8362 5 1 1 8361
0 8363 7 1 2 65520 8362
0 8364 5 1 1 8363
0 8365 7 1 2 69402 8364
0 8366 5 1 1 8365
0 8367 7 9 2 50945 51509
0 8368 7 5 2 49996 69404
0 8369 7 5 2 68746 69413
0 8370 7 1 2 65540 65182
0 8371 7 1 2 69418 8370
0 8372 5 1 1 8371
0 8373 7 1 2 8366 8372
0 8374 5 1 1 8373
0 8375 7 1 2 54544 8374
0 8376 5 1 1 8375
0 8377 7 8 2 54920 60526
0 8378 7 5 2 49997 51510
0 8379 7 1 2 69431 68759
0 8380 7 1 2 69423 8379
0 8381 5 1 1 8380
0 8382 7 3 2 49108 53769
0 8383 7 3 2 49692 53877
0 8384 7 1 2 69439 69147
0 8385 7 1 2 69436 8384
0 8386 7 1 2 68619 8385
0 8387 5 1 1 8386
0 8388 7 1 2 8381 8387
0 8389 7 1 2 8376 8388
0 8390 5 1 1 8389
0 8391 7 1 2 55613 8390
0 8392 5 1 1 8391
0 8393 7 7 2 53436 49998
0 8394 5 1 1 69442
0 8395 7 1 2 69443 69108
0 8396 7 1 2 64060 8395
0 8397 5 1 1 8396
0 8398 7 1 2 8392 8397
0 8399 5 1 1 8398
0 8400 7 1 2 55250 8399
0 8401 5 1 1 8400
0 8402 7 1 2 48499 53770
0 8403 7 2 2 69148 8402
0 8404 7 1 2 69449 69162
0 8405 7 1 2 64061 8404
0 8406 5 1 1 8405
0 8407 7 1 2 8401 8406
0 8408 5 1 1 8407
0 8409 7 1 2 62827 8408
0 8410 5 1 1 8409
0 8411 7 7 2 51511 68511
0 8412 7 1 2 56853 69451
0 8413 5 1 1 8412
0 8414 7 1 2 66437 8413
0 8415 5 1 1 8414
0 8416 7 1 2 49999 8415
0 8417 5 1 1 8416
0 8418 7 12 2 53771 55251
0 8419 7 3 2 68187 69458
0 8420 5 1 1 69470
0 8421 7 1 2 67823 69471
0 8422 5 1 1 8421
0 8423 7 1 2 8417 8422
0 8424 5 1 1 8423
0 8425 7 1 2 64062 8424
0 8426 5 1 1 8425
0 8427 7 2 2 58380 64918
0 8428 7 1 2 67418 69473
0 8429 5 1 1 8428
0 8430 7 1 2 66111 8429
0 8431 5 1 1 8430
0 8432 7 1 2 50000 8431
0 8433 5 1 1 8432
0 8434 7 5 2 50001 55252
0 8435 7 2 2 66448 69475
0 8436 7 1 2 64067 69480
0 8437 5 1 1 8436
0 8438 7 1 2 8433 8437
0 8439 5 1 1 8438
0 8440 7 1 2 58965 8439
0 8441 5 1 1 8440
0 8442 7 1 2 8426 8441
0 8443 5 1 1 8442
0 8444 7 1 2 54921 8443
0 8445 5 1 1 8444
0 8446 7 1 2 69255 69325
0 8447 5 1 1 8446
0 8448 7 2 2 54213 65183
0 8449 5 4 1 69482
0 8450 7 1 2 67010 69272
0 8451 7 1 2 69483 8450
0 8452 5 1 1 8451
0 8453 7 2 2 53984 59519
0 8454 5 1 1 69488
0 8455 7 1 2 57753 8454
0 8456 5 1 1 8455
0 8457 7 1 2 55253 69452
0 8458 7 1 2 8456 8457
0 8459 5 1 1 8458
0 8460 7 1 2 8452 8459
0 8461 7 1 2 8447 8460
0 8462 5 1 1 8461
0 8463 7 1 2 50002 8462
0 8464 5 1 1 8463
0 8465 7 1 2 8445 8464
0 8466 5 1 1 8465
0 8467 7 1 2 51704 8466
0 8468 5 1 1 8467
0 8469 7 2 2 58665 65184
0 8470 5 1 1 69490
0 8471 7 1 2 50946 8470
0 8472 5 1 1 8471
0 8473 7 2 2 53772 68452
0 8474 5 1 1 69492
0 8475 7 2 2 65697 69493
0 8476 5 1 1 69494
0 8477 7 1 2 68188 69495
0 8478 7 1 2 8472 8477
0 8479 5 1 1 8478
0 8480 7 1 2 8468 8479
0 8481 5 1 1 8480
0 8482 7 1 2 48992 8481
0 8483 5 1 1 8482
0 8484 7 5 2 53773 54545
0 8485 7 2 2 55254 69496
0 8486 5 1 1 69501
0 8487 7 1 2 50369 61729
0 8488 5 1 1 8487
0 8489 7 1 2 69502 8488
0 8490 7 1 2 69164 8489
0 8491 5 1 1 8490
0 8492 7 1 2 8483 8491
0 8493 7 1 2 8410 8492
0 8494 5 1 1 8493
0 8495 7 1 2 57144 8494
0 8496 5 1 1 8495
0 8497 7 1 2 8357 8496
0 8498 7 1 2 8228 8497
0 8499 5 1 1 8498
0 8500 7 1 2 48893 8499
0 8501 5 1 1 8500
0 8502 7 1 2 7992 8501
0 8503 5 1 1 8502
0 8504 7 1 2 56055 8503
0 8505 5 1 1 8504
0 8506 7 1 2 66336 69057
0 8507 5 1 1 8506
0 8508 7 1 2 68409 8507
0 8509 5 1 1 8508
0 8510 7 1 2 53437 8509
0 8511 5 1 1 8510
0 8512 7 4 2 51240 63504
0 8513 7 1 2 65541 69503
0 8514 5 1 1 8513
0 8515 7 1 2 8511 8514
0 8516 5 1 1 8515
0 8517 7 1 2 68544 8516
0 8518 5 1 1 8517
0 8519 7 1 2 63110 68339
0 8520 5 1 1 8519
0 8521 7 1 2 56854 65043
0 8522 5 2 1 8521
0 8523 7 1 2 6926 69507
0 8524 5 1 1 8523
0 8525 7 5 2 53985 64785
0 8526 5 1 1 69509
0 8527 7 1 2 53438 8526
0 8528 5 2 1 8527
0 8529 7 33 2 52767 53651
0 8530 5 31 1 69516
0 8531 7 2 2 54546 69549
0 8532 7 1 2 69514 69580
0 8533 7 1 2 8524 8532
0 8534 5 1 1 8533
0 8535 7 1 2 8520 8534
0 8536 5 1 1 8535
0 8537 7 1 2 51705 8536
0 8538 5 1 1 8537
0 8539 7 1 2 8518 8538
0 8540 5 1 1 8539
0 8541 7 1 2 51512 8540
0 8542 5 1 1 8541
0 8543 7 6 2 51241 69550
0 8544 7 1 2 56986 68060
0 8545 5 1 1 8544
0 8546 7 1 2 69582 8545
0 8547 5 1 1 8546
0 8548 7 1 2 67094 66699
0 8549 5 1 1 8548
0 8550 7 1 2 65044 66815
0 8551 5 1 1 8550
0 8552 7 1 2 8549 8551
0 8553 5 1 1 8552
0 8554 7 1 2 67675 8553
0 8555 5 1 1 8554
0 8556 7 1 2 8547 8555
0 8557 5 1 1 8556
0 8558 7 1 2 67917 8557
0 8559 5 1 1 8558
0 8560 7 1 2 8542 8559
0 8561 5 1 1 8560
0 8562 7 1 2 48993 8561
0 8563 5 1 1 8562
0 8564 7 2 2 59599 69299
0 8565 7 2 2 49856 67653
0 8566 7 1 2 65564 69590
0 8567 7 1 2 69588 8566
0 8568 5 1 1 8567
0 8569 7 1 2 8563 8568
0 8570 5 1 1 8569
0 8571 7 1 2 58848 8570
0 8572 5 1 1 8571
0 8573 7 10 2 51513 69551
0 8574 5 1 1 69592
0 8575 7 5 2 53986 55255
0 8576 7 1 2 65147 69602
0 8577 5 2 1 8576
0 8578 7 1 2 65521 69607
0 8579 5 1 1 8578
0 8580 7 1 2 49693 8579
0 8581 5 1 1 8580
0 8582 7 31 2 48894 49857
0 8583 5 17 1 69609
0 8584 7 2 2 64786 64703
0 8585 7 2 2 56855 60913
0 8586 5 1 1 69659
0 8587 7 1 2 69657 69660
0 8588 5 1 1 8587
0 8589 7 1 2 69640 8588
0 8590 7 1 2 8581 8589
0 8591 5 1 1 8590
0 8592 7 1 2 69593 8591
0 8593 5 1 1 8592
0 8594 7 4 2 50370 56987
0 8595 5 4 1 69661
0 8596 7 3 2 66201 69665
0 8597 7 1 2 66410 68820
0 8598 7 1 2 69669 8597
0 8599 5 1 1 8598
0 8600 7 1 2 8593 8599
0 8601 5 1 1 8600
0 8602 7 1 2 54547 8601
0 8603 5 1 1 8602
0 8604 7 1 2 59499 69610
0 8605 5 1 1 8604
0 8606 7 1 2 66373 69552
0 8607 7 1 2 67056 8606
0 8608 5 1 1 8607
0 8609 7 1 2 8605 8608
0 8610 5 1 1 8609
0 8611 7 1 2 51514 8610
0 8612 5 1 1 8611
0 8613 7 2 2 55475 67676
0 8614 7 3 2 48500 62281
0 8615 7 1 2 59600 69674
0 8616 5 2 1 8615
0 8617 7 1 2 66627 69677
0 8618 5 1 1 8617
0 8619 7 1 2 69672 8618
0 8620 5 1 1 8619
0 8621 7 1 2 8612 8620
0 8622 5 1 1 8621
0 8623 7 1 2 68136 8622
0 8624 5 1 1 8623
0 8625 7 2 2 55476 64140
0 8626 7 1 2 69583 69679
0 8627 5 1 1 8626
0 8628 7 1 2 8624 8627
0 8629 7 1 2 8603 8628
0 8630 5 1 1 8629
0 8631 7 1 2 51706 8630
0 8632 5 1 1 8631
0 8633 7 2 2 53439 64141
0 8634 5 3 1 69681
0 8635 7 3 2 53878 50947
0 8636 7 1 2 56856 69686
0 8637 5 1 1 8636
0 8638 7 1 2 69683 8637
0 8639 5 1 1 8638
0 8640 7 2 2 68453 68688
0 8641 7 1 2 53652 68083
0 8642 7 1 2 69689 8641
0 8643 7 1 2 8639 8642
0 8644 5 1 1 8643
0 8645 7 1 2 8632 8644
0 8646 5 1 1 8645
0 8647 7 1 2 48994 8646
0 8648 5 1 1 8647
0 8649 7 1 2 59500 65280
0 8650 7 1 2 67918 69306
0 8651 7 1 2 8649 8650
0 8652 7 1 2 68137 68413
0 8653 7 1 2 8651 8652
0 8654 5 1 1 8653
0 8655 7 1 2 8648 8654
0 8656 7 1 2 8572 8655
0 8657 5 1 1 8656
0 8658 7 1 2 58106 8657
0 8659 5 1 1 8658
0 8660 7 8 2 67259 68178
0 8661 5 2 1 69691
0 8662 7 1 2 52856 69699
0 8663 5 5 1 8662
0 8664 7 1 2 67177 68640
0 8665 5 2 1 8664
0 8666 7 7 2 50641 55477
0 8667 7 2 2 69708 69687
0 8668 7 1 2 68138 69715
0 8669 5 1 1 8668
0 8670 7 1 2 60914 68282
0 8671 5 1 1 8670
0 8672 7 1 2 8669 8671
0 8673 5 2 1 8672
0 8674 7 1 2 55256 69717
0 8675 5 1 1 8674
0 8676 7 1 2 69706 8675
0 8677 5 1 1 8676
0 8678 7 1 2 56857 8677
0 8679 5 1 1 8678
0 8680 7 5 2 54922 66071
0 8681 5 2 1 69719
0 8682 7 1 2 61668 60982
0 8683 5 1 1 8682
0 8684 7 1 2 67764 8683
0 8685 5 1 1 8684
0 8686 7 1 2 69724 8685
0 8687 5 1 1 8686
0 8688 7 1 2 49694 8687
0 8689 5 1 1 8688
0 8690 7 1 2 8679 8689
0 8691 5 1 1 8690
0 8692 7 1 2 62842 8691
0 8693 5 1 1 8692
0 8694 7 2 2 53879 68139
0 8695 5 1 1 69726
0 8696 7 1 2 49695 69727
0 8697 5 1 1 8696
0 8698 7 1 2 65087 8697
0 8699 5 1 1 8698
0 8700 7 1 2 51515 69692
0 8701 7 1 2 8699 8700
0 8702 5 1 1 8701
0 8703 7 1 2 8693 8702
0 8704 5 1 1 8703
0 8705 7 1 2 51707 8704
0 8706 5 1 1 8705
0 8707 7 2 2 52768 55614
0 8708 7 1 2 53880 66261
0 8709 5 1 1 8708
0 8710 7 1 2 67483 8709
0 8711 5 1 1 8710
0 8712 7 1 2 69728 8711
0 8713 5 1 1 8712
0 8714 7 1 2 63857 67919
0 8715 7 1 2 62843 8714
0 8716 5 1 1 8715
0 8717 7 1 2 8713 8716
0 8718 5 1 1 8717
0 8719 7 1 2 53653 8718
0 8720 5 1 1 8719
0 8721 7 1 2 51242 69716
0 8722 5 1 1 8721
0 8723 7 1 2 68284 8722
0 8724 5 1 1 8723
0 8725 7 4 2 55615 69517
0 8726 7 1 2 60915 69730
0 8727 7 1 2 8724 8726
0 8728 5 1 1 8727
0 8729 7 1 2 8720 8728
0 8730 7 1 2 8706 8729
0 8731 5 1 1 8730
0 8732 7 1 2 54214 8731
0 8733 5 1 1 8732
0 8734 7 2 2 52769 68476
0 8735 7 2 2 68534 69734
0 8736 5 1 1 69736
0 8737 7 1 2 56988 68133
0 8738 5 1 1 8737
0 8739 7 2 2 66202 8738
0 8740 7 1 2 62844 66485
0 8741 7 1 2 69738 8740
0 8742 5 1 1 8741
0 8743 7 4 2 53881 69603
0 8744 5 1 1 69740
0 8745 7 1 2 64905 8744
0 8746 5 1 1 8745
0 8747 7 1 2 60916 8746
0 8748 5 1 1 8747
0 8749 7 1 2 54923 64963
0 8750 5 1 1 8749
0 8751 7 1 2 53440 8750
0 8752 7 1 2 8748 8751
0 8753 5 1 1 8752
0 8754 7 1 2 53654 62834
0 8755 5 4 1 8754
0 8756 7 3 2 62845 69744
0 8757 5 1 1 69748
0 8758 7 1 2 69594 69749
0 8759 7 1 2 8753 8758
0 8760 5 1 1 8759
0 8761 7 1 2 8742 8760
0 8762 5 1 1 8761
0 8763 7 1 2 51708 8762
0 8764 5 1 1 8763
0 8765 7 1 2 8736 8764
0 8766 5 1 1 8765
0 8767 7 1 2 54548 8766
0 8768 5 1 1 8767
0 8769 7 1 2 63858 69675
0 8770 5 1 1 8769
0 8771 7 1 2 53655 8770
0 8772 5 1 1 8771
0 8773 7 1 2 62846 8772
0 8774 5 1 1 8773
0 8775 7 1 2 69700 8774
0 8776 5 1 1 8775
0 8777 7 1 2 51709 8776
0 8778 5 1 1 8777
0 8779 7 3 2 54924 55616
0 8780 7 4 2 54549 69751
0 8781 7 2 2 53656 53882
0 8782 7 2 2 52770 69758
0 8783 7 1 2 69754 69760
0 8784 5 1 1 8783
0 8785 7 1 2 8778 8784
0 8786 5 1 1 8785
0 8787 7 1 2 60381 8786
0 8788 5 1 1 8787
0 8789 7 1 2 68674 8788
0 8790 5 1 1 8789
0 8791 7 1 2 49696 8790
0 8792 5 1 1 8791
0 8793 7 1 2 64794 69508
0 8794 5 1 1 8793
0 8795 7 1 2 51710 69581
0 8796 7 1 2 8794 8795
0 8797 7 1 2 69750 8796
0 8798 5 1 1 8797
0 8799 7 1 2 51516 8798
0 8800 7 1 2 8792 8799
0 8801 5 1 1 8800
0 8802 7 5 2 50642 68377
0 8803 5 3 1 69762
0 8804 7 2 2 60382 69763
0 8805 5 1 1 69770
0 8806 7 1 2 68600 8805
0 8807 5 1 1 8806
0 8808 7 1 2 56858 8807
0 8809 5 1 1 8808
0 8810 7 3 2 53657 64587
0 8811 5 1 1 69772
0 8812 7 1 2 51243 67654
0 8813 5 2 1 8812
0 8814 7 1 2 8811 69775
0 8815 5 2 1 8814
0 8816 7 1 2 65045 69777
0 8817 5 1 1 8816
0 8818 7 1 2 8809 8817
0 8819 5 1 1 8818
0 8820 7 1 2 51711 62847
0 8821 7 1 2 8819 8820
0 8822 5 1 1 8821
0 8823 7 2 2 66245 68292
0 8824 7 1 2 69518 68519
0 8825 7 1 2 69779 8824
0 8826 5 1 1 8825
0 8827 7 1 2 55478 8826
0 8828 7 1 2 8822 8827
0 8829 5 1 1 8828
0 8830 7 1 2 58849 8829
0 8831 7 1 2 8801 8830
0 8832 5 1 1 8831
0 8833 7 1 2 8768 8832
0 8834 7 1 2 8733 8833
0 8835 5 1 1 8834
0 8836 7 1 2 48995 8835
0 8837 5 1 1 8836
0 8838 7 1 2 56859 69718
0 8839 5 1 1 8838
0 8840 7 3 2 53441 63445
0 8841 7 1 2 55479 69781
0 8842 5 1 1 8841
0 8843 7 1 2 8839 8842
0 8844 5 1 1 8843
0 8845 7 1 2 55257 8844
0 8846 5 1 1 8845
0 8847 7 1 2 68539 8846
0 8848 5 1 1 8847
0 8849 7 1 2 54215 8848
0 8850 5 1 1 8849
0 8851 7 28 2 53442 55258
0 8852 5 1 1 69784
0 8853 7 1 2 67011 69785
0 8854 7 1 2 69739 8853
0 8855 5 1 1 8854
0 8856 7 1 2 8850 8855
0 8857 5 1 1 8856
0 8858 7 1 2 69022 8857
0 8859 5 1 1 8858
0 8860 7 5 2 69405 68520
0 8861 7 1 2 67655 66816
0 8862 7 2 2 69812 8861
0 8863 5 1 1 69817
0 8864 7 1 2 69818 69474
0 8865 5 1 1 8864
0 8866 7 3 2 67920 68641
0 8867 5 5 1 69819
0 8868 7 1 2 69786 69820
0 8869 5 2 1 8868
0 8870 7 3 2 56860 65973
0 8871 7 2 2 60527 69013
0 8872 5 1 1 69832
0 8873 7 1 2 49858 63402
0 8874 7 1 2 68682 8873
0 8875 5 1 1 8874
0 8876 7 1 2 8872 8875
0 8877 5 1 1 8876
0 8878 7 1 2 69829 8877
0 8879 5 1 1 8878
0 8880 7 1 2 69373 8879
0 8881 5 1 1 8880
0 8882 7 1 2 53987 8881
0 8883 5 1 1 8882
0 8884 7 1 2 69827 8883
0 8885 5 1 1 8884
0 8886 7 1 2 65046 8885
0 8887 5 1 1 8886
0 8888 7 2 2 50948 68454
0 8889 7 1 2 67047 69834
0 8890 5 1 1 8889
0 8891 7 1 2 69359 8890
0 8892 5 2 1 8891
0 8893 7 1 2 68573 69836
0 8894 5 1 1 8893
0 8895 7 1 2 60383 69321
0 8896 5 1 1 8895
0 8897 7 1 2 8894 8896
0 8898 5 1 1 8897
0 8899 7 1 2 56861 8898
0 8900 5 1 1 8899
0 8901 7 1 2 8887 8900
0 8902 5 1 1 8901
0 8903 7 1 2 58850 8902
0 8904 5 1 1 8903
0 8905 7 1 2 8865 8904
0 8906 7 1 2 8859 8905
0 8907 7 1 2 8837 8906
0 8908 5 1 1 8907
0 8909 7 1 2 69701 8908
0 8910 5 1 1 8909
0 8911 7 1 2 8659 8910
0 8912 5 1 1 8911
0 8913 7 1 2 50003 8912
0 8914 5 1 1 8913
0 8915 7 4 2 68204 68945
0 8916 7 3 2 54550 69838
0 8917 5 1 1 69842
0 8918 7 4 2 50145 62076
0 8919 5 1 1 69845
0 8920 7 1 2 65369 69846
0 8921 5 1 1 8920
0 8922 7 1 2 69843 8921
0 8923 5 1 1 8922
0 8924 7 2 2 53988 69078
0 8925 5 1 1 69849
0 8926 7 1 2 51244 59446
0 8927 7 1 2 69850 8926
0 8928 5 1 1 8927
0 8929 7 1 2 8923 8928
0 8930 5 1 1 8929
0 8931 7 1 2 54925 8930
0 8932 5 1 1 8931
0 8933 7 3 2 55617 64588
0 8934 7 2 2 54216 68205
0 8935 7 2 2 69851 69854
0 8936 5 1 1 69856
0 8937 7 1 2 49109 69857
0 8938 5 1 1 8937
0 8939 7 6 2 48996 56862
0 8940 7 2 2 51245 51712
0 8941 7 1 2 58851 69864
0 8942 7 1 2 69858 8941
0 8943 5 1 1 8942
0 8944 7 1 2 8938 8943
0 8945 7 1 2 8932 8944
0 8946 5 1 1 8945
0 8947 7 1 2 55480 8946
0 8948 5 1 1 8947
0 8949 7 2 2 48997 63863
0 8950 7 2 2 56863 69866
0 8951 7 5 2 58422 62077
0 8952 5 17 1 69870
0 8953 7 2 2 51713 69875
0 8954 7 1 2 66678 69892
0 8955 7 1 2 69868 8954
0 8956 5 1 1 8955
0 8957 7 1 2 8948 8956
0 8958 5 1 1 8957
0 8959 7 1 2 49859 8958
0 8960 5 1 1 8959
0 8961 7 4 2 48998 51246
0 8962 7 1 2 69894 69109
0 8963 5 1 1 8962
0 8964 7 5 2 67824 69459
0 8965 7 2 2 52857 69898
0 8966 5 1 1 69903
0 8967 7 11 2 51247 51517
0 8968 7 2 2 69905 68972
0 8969 7 1 2 69916 69859
0 8970 5 1 1 8969
0 8971 7 1 2 8966 8970
0 8972 5 1 1 8971
0 8973 7 3 2 54551 55618
0 8974 7 1 2 47847 69918
0 8975 7 1 2 8972 8974
0 8976 5 1 1 8975
0 8977 7 1 2 8963 8976
0 8978 5 1 1 8977
0 8979 7 1 2 64050 8978
0 8980 5 1 1 8979
0 8981 7 3 2 51518 69860
0 8982 5 1 1 69921
0 8983 7 1 2 63555 69297
0 8984 7 1 2 69922 8983
0 8985 5 1 1 8984
0 8986 7 1 2 8980 8985
0 8987 7 1 2 8960 8986
0 8988 5 1 1 8987
0 8989 7 1 2 49697 8988
0 8990 5 1 1 8989
0 8991 7 1 2 67095 68894
0 8992 5 1 1 8991
0 8993 7 4 2 53774 53883
0 8994 7 1 2 68473 69924
0 8995 5 1 1 8994
0 8996 7 1 2 8992 8995
0 8997 5 1 1 8996
0 8998 7 1 2 48999 8997
0 8999 5 1 1 8998
0 9000 7 7 2 54926 58666
0 9001 7 1 2 69928 69925
0 9002 7 1 2 69153 9001
0 9003 5 1 1 9002
0 9004 7 1 2 8999 9003
0 9005 5 1 1 9004
0 9006 7 1 2 66700 9005
0 9007 5 1 1 9006
0 9008 7 2 2 63446 67921
0 9009 7 11 2 49860 53775
0 9010 7 2 2 49000 53884
0 9011 7 1 2 69937 69948
0 9012 7 1 2 69935 9011
0 9013 5 1 1 9012
0 9014 7 1 2 9007 9013
0 9015 5 1 1 9014
0 9016 7 1 2 58852 9015
0 9017 5 1 1 9016
0 9018 7 1 2 53776 63447
0 9019 5 1 1 9018
0 9020 7 1 2 69678 9019
0 9021 5 1 1 9020
0 9022 7 1 2 68140 9021
0 9023 5 1 1 9022
0 9024 7 1 2 69497 69670
0 9025 5 1 1 9024
0 9026 7 1 2 9023 9025
0 9027 5 1 1 9026
0 9028 7 1 2 69079 9027
0 9029 5 1 1 9028
0 9030 7 6 2 52858 55619
0 9031 7 2 2 65437 69950
0 9032 7 3 2 53777 60384
0 9033 7 1 2 67084 69958
0 9034 7 1 2 69956 9033
0 9035 5 1 1 9034
0 9036 7 1 2 9029 9035
0 9037 5 1 1 9036
0 9038 7 1 2 67825 9037
0 9039 5 1 1 9038
0 9040 7 1 2 9017 9039
0 9041 5 1 1 9040
0 9042 7 1 2 55259 9041
0 9043 5 1 1 9042
0 9044 7 1 2 8990 9043
0 9045 5 1 1 9044
0 9046 7 1 2 68189 9045
0 9047 5 1 1 9046
0 9048 7 9 2 59125 69080
0 9049 5 1 1 69961
0 9050 7 1 2 65185 69962
0 9051 5 1 1 9050
0 9052 7 3 2 47848 68206
0 9053 7 1 2 69755 69970
0 9054 5 1 1 9053
0 9055 7 1 2 9049 9054
0 9056 5 1 1 9055
0 9057 7 1 2 55736 9056
0 9058 5 1 1 9057
0 9059 7 2 2 63448 69951
0 9060 7 1 2 53885 69437
0 9061 7 1 2 69973 9060
0 9062 5 1 1 9061
0 9063 7 1 2 9058 9062
0 9064 5 1 1 9063
0 9065 7 1 2 53989 9064
0 9066 5 1 1 9065
0 9067 7 1 2 9051 9066
0 9068 5 1 1 9067
0 9069 7 1 2 67898 68612
0 9070 7 1 2 69400 9069
0 9071 7 1 2 9068 9070
0 9072 5 1 1 9071
0 9073 7 1 2 9047 9072
0 9074 5 1 1 9073
0 9075 7 1 2 48895 9074
0 9076 5 1 1 9075
0 9077 7 6 2 50949 55620
0 9078 7 4 2 68747 69975
0 9079 5 1 1 69981
0 9080 7 8 2 51714 69553
0 9081 7 5 2 62540 69985
0 9082 7 1 2 58667 69993
0 9083 5 1 1 9082
0 9084 7 1 2 9079 9083
0 9085 5 1 1 9084
0 9086 7 1 2 49001 9085
0 9087 5 1 1 9086
0 9088 7 1 2 64642 65648
0 9089 7 1 2 63200 66804
0 9090 7 1 2 68477 69293
0 9091 7 1 2 9089 9090
0 9092 7 1 2 9088 9091
0 9093 5 1 1 9092
0 9094 7 1 2 9087 9093
0 9095 5 1 1 9094
0 9096 7 1 2 55260 9095
0 9097 5 1 1 9096
0 9098 7 1 2 52859 67165
0 9099 5 3 1 9098
0 9100 7 1 2 65068 69998
0 9101 7 1 2 69369 9100
0 9102 5 1 1 9101
0 9103 7 1 2 9097 9102
0 9104 5 1 1 9103
0 9105 7 1 2 51519 9104
0 9106 5 1 1 9105
0 9107 7 4 2 62895 69611
0 9108 5 2 1 70001
0 9109 7 5 2 62943 69519
0 9110 5 12 1 70007
0 9111 7 1 2 49002 70012
0 9112 5 1 1 9111
0 9113 7 1 2 70005 9112
0 9114 5 1 1 9113
0 9115 7 8 2 51715 66072
0 9116 7 4 2 54927 60917
0 9117 5 2 1 70032
0 9118 7 1 2 56989 70036
0 9119 5 1 1 9118
0 9120 7 2 2 70024 9119
0 9121 7 1 2 9114 70038
0 9122 5 1 1 9121
0 9123 7 1 2 9106 9122
0 9124 5 1 1 9123
0 9125 7 1 2 50004 9124
0 9126 5 1 1 9125
0 9127 7 1 2 69374 8476
0 9128 5 1 1 9127
0 9129 7 1 2 70033 9128
0 9130 5 1 1 9129
0 9131 7 1 2 68783 69837
0 9132 5 1 1 9131
0 9133 7 1 2 9130 9132
0 9134 5 1 1 9133
0 9135 7 1 2 49003 9134
0 9136 5 1 1 9135
0 9137 7 3 2 52860 49698
0 9138 7 4 2 69938 70040
0 9139 7 6 2 55261 69139
0 9140 7 2 2 58668 70047
0 9141 7 1 2 70043 70053
0 9142 5 1 1 9141
0 9143 7 1 2 9136 9142
0 9144 5 1 1 9143
0 9145 7 1 2 65623 9144
0 9146 5 1 1 9145
0 9147 7 1 2 9126 9146
0 9148 5 1 1 9147
0 9149 7 1 2 57893 9148
0 9150 5 1 1 9149
0 9151 7 3 2 63085 68496
0 9152 5 2 1 70055
0 9153 7 6 2 69554 70056
0 9154 7 8 2 51716 70060
0 9155 5 1 1 70066
0 9156 7 1 2 58669 70067
0 9157 5 1 1 9156
0 9158 7 3 2 48712 50950
0 9159 5 3 1 70074
0 9160 7 2 2 53443 70077
0 9161 7 1 2 62647 68870
0 9162 7 1 2 69137 9161
0 9163 5 1 1 9162
0 9164 7 1 2 70080 9163
0 9165 5 1 1 9164
0 9166 7 1 2 3355 68545
0 9167 7 1 2 9165 9166
0 9168 5 1 1 9167
0 9169 7 1 2 9157 9168
0 9170 5 1 1 9169
0 9171 7 1 2 55262 9170
0 9172 5 1 1 9171
0 9173 7 12 2 51248 62541
0 9174 5 1 1 70082
0 9175 7 2 2 69976 70083
0 9176 7 1 2 65542 66817
0 9177 7 1 2 70094 9176
0 9178 5 1 1 9177
0 9179 7 1 2 9172 9178
0 9180 5 1 1 9179
0 9181 7 1 2 51520 9180
0 9182 5 1 1 9181
0 9183 7 3 2 64378 69240
0 9184 5 2 1 70096
0 9185 7 1 2 70099 70039
0 9186 5 1 1 9185
0 9187 7 1 2 9182 9186
0 9188 5 1 1 9187
0 9189 7 1 2 68229 9188
0 9190 5 1 1 9189
0 9191 7 1 2 9150 9190
0 9192 5 1 1 9191
0 9193 7 1 2 60690 9192
0 9194 5 1 1 9193
0 9195 7 1 2 9076 9194
0 9196 7 1 2 8914 9195
0 9197 7 1 2 8505 9196
0 9198 5 1 1 9197
0 9199 7 1 2 62398 9198
0 9200 5 1 1 9199
0 9201 7 8 2 52477 56179
0 9202 5 3 1 70101
0 9203 7 3 2 53264 57309
0 9204 5 2 1 70112
0 9205 7 5 2 70109 70115
0 9206 5 18 1 70117
0 9207 7 1 2 1212 70122
0 9208 5 1 1 9207
0 9209 7 17 2 52374 52478
0 9210 5 3 1 70140
0 9211 7 19 2 60511 70141
0 9212 5 5 1 70160
0 9213 7 2 2 50371 61805
0 9214 5 2 1 70184
0 9215 7 2 2 63995 70186
0 9216 5 1 1 70188
0 9217 7 2 2 54217 60869
0 9218 5 2 1 70190
0 9219 7 2 2 52071 70192
0 9220 5 2 1 70194
0 9221 7 3 2 57426 59982
0 9222 5 7 1 70198
0 9223 7 4 2 49190 61174
0 9224 5 11 1 70208
0 9225 7 2 2 70201 70212
0 9226 5 1 1 70223
0 9227 7 1 2 67358 9226
0 9228 7 2 2 70196 9227
0 9229 7 1 2 70189 70225
0 9230 5 1 1 9229
0 9231 7 1 2 70161 9230
0 9232 5 1 1 9231
0 9233 7 1 2 9208 9232
0 9234 5 1 1 9233
0 9235 7 1 2 62944 9234
0 9236 5 1 1 9235
0 9237 7 3 2 54218 59806
0 9238 5 1 1 70227
0 9239 7 1 2 56056 70228
0 9240 5 1 1 9239
0 9241 7 2 2 63228 9240
0 9242 7 1 2 61466 70230
0 9243 5 1 1 9242
0 9244 7 6 2 54219 61546
0 9245 5 22 1 70232
0 9246 7 3 2 53054 70238
0 9247 5 2 1 70260
0 9248 7 2 2 65350 59747
0 9249 5 2 1 70265
0 9250 7 1 2 52072 70267
0 9251 5 1 1 9250
0 9252 7 2 2 70263 9251
0 9253 7 1 2 60231 70269
0 9254 5 1 1 9253
0 9255 7 1 2 52230 9254
0 9256 5 1 1 9255
0 9257 7 2 2 52935 60771
0 9258 7 2 2 60491 70271
0 9259 5 2 1 70273
0 9260 7 1 2 59764 70275
0 9261 5 1 1 9260
0 9262 7 1 2 51850 9261
0 9263 5 4 1 9262
0 9264 7 3 2 50372 61827
0 9265 5 2 1 70281
0 9266 7 1 2 53055 70282
0 9267 5 1 1 9266
0 9268 7 1 2 61318 9267
0 9269 7 1 2 70277 9268
0 9270 7 1 2 9256 9269
0 9271 7 1 2 9243 9270
0 9272 5 1 1 9271
0 9273 7 1 2 50643 9272
0 9274 5 1 1 9273
0 9275 7 3 2 60435 63920
0 9276 7 1 2 70187 70286
0 9277 7 1 2 70197 9276
0 9278 5 1 1 9277
0 9279 7 1 2 61327 9278
0 9280 5 1 1 9279
0 9281 7 7 2 50644 63757
0 9282 7 1 2 57576 70289
0 9283 5 1 1 9282
0 9284 7 1 2 61319 9283
0 9285 5 1 1 9284
0 9286 7 1 2 70224 9285
0 9287 5 1 1 9286
0 9288 7 5 2 52879 60097
0 9289 7 2 2 58318 70296
0 9290 5 1 1 70301
0 9291 7 2 2 60261 70302
0 9292 5 1 1 70303
0 9293 7 1 2 52936 70304
0 9294 5 3 1 9293
0 9295 7 1 2 56545 70305
0 9296 7 1 2 9287 9295
0 9297 7 1 2 9280 9296
0 9298 7 1 2 9274 9297
0 9299 5 1 1 9298
0 9300 7 1 2 70097 9299
0 9301 5 1 1 9300
0 9302 7 1 2 9236 9301
0 9303 5 1 1 9302
0 9304 7 1 2 54928 69641
0 9305 7 1 2 9303 9304
0 9306 5 1 1 9305
0 9307 7 1 2 67750 70008
0 9308 5 1 1 9307
0 9309 7 2 2 58670 69642
0 9310 7 2 2 62542 70110
0 9311 5 1 1 70310
0 9312 7 1 2 70116 70311
0 9313 5 1 1 9312
0 9314 7 1 2 62945 9313
0 9315 5 3 1 9314
0 9316 7 1 2 69555 70312
0 9317 5 1 1 9316
0 9318 7 1 2 70308 9317
0 9319 5 1 1 9318
0 9320 7 3 2 50645 60114
0 9321 5 1 1 70315
0 9322 7 1 2 61134 9321
0 9323 5 1 1 9322
0 9324 7 1 2 50146 9323
0 9325 5 1 1 9324
0 9326 7 1 2 52073 64460
0 9327 5 1 1 9326
0 9328 7 1 2 54552 60451
0 9329 5 3 1 9328
0 9330 7 1 2 63758 70318
0 9331 5 1 1 9330
0 9332 7 1 2 9327 9331
0 9333 7 1 2 9325 9332
0 9334 5 2 1 9333
0 9335 7 10 2 49699 58740
0 9336 5 5 1 70323
0 9337 7 3 2 61360 70324
0 9338 5 2 1 70338
0 9339 7 1 2 53658 70339
0 9340 7 1 2 70321 9339
0 9341 5 1 1 9340
0 9342 7 1 2 9319 9341
0 9343 5 1 1 9342
0 9344 7 1 2 59844 9343
0 9345 5 1 1 9344
0 9346 7 2 2 57427 68714
0 9347 5 1 1 70343
0 9348 7 1 2 62126 60087
0 9349 5 4 1 9348
0 9350 7 1 2 54553 69241
0 9351 7 1 2 70345 9350
0 9352 5 1 1 9351
0 9353 7 1 2 9347 9352
0 9354 5 1 1 9353
0 9355 7 1 2 54220 9354
0 9356 5 1 1 9355
0 9357 7 2 2 56864 68715
0 9358 5 1 1 70349
0 9359 7 1 2 9356 9358
0 9360 5 1 1 9359
0 9361 7 1 2 52771 9360
0 9362 5 1 1 9361
0 9363 7 1 2 54554 62470
0 9364 7 1 2 66739 9363
0 9365 7 1 2 70346 9364
0 9366 5 1 1 9365
0 9367 7 1 2 9362 9366
0 9368 7 1 2 9345 9367
0 9369 5 1 1 9368
0 9370 7 1 2 50951 9369
0 9371 5 1 1 9370
0 9372 7 1 2 9308 9371
0 9373 7 1 2 9306 9372
0 9374 5 1 1 9373
0 9375 7 1 2 55481 9374
0 9376 5 1 1 9375
0 9377 7 2 2 65336 55671
0 9378 5 3 1 70351
0 9379 7 1 2 58326 70353
0 9380 5 1 1 9379
0 9381 7 1 2 53056 9380
0 9382 5 1 1 9381
0 9383 7 1 2 64470 9382
0 9384 5 1 1 9383
0 9385 7 1 2 52074 9384
0 9386 5 1 1 9385
0 9387 7 2 2 54221 59826
0 9388 5 1 1 70356
0 9389 7 1 2 59812 70357
0 9390 5 1 1 9389
0 9391 7 1 2 50646 9390
0 9392 5 1 1 9391
0 9393 7 1 2 9386 9392
0 9394 5 1 1 9393
0 9395 7 1 2 50147 9394
0 9396 5 1 1 9395
0 9397 7 1 2 50647 59792
0 9398 5 1 1 9397
0 9399 7 7 2 48341 56696
0 9400 5 20 1 70358
0 9401 7 3 2 49302 70359
0 9402 5 19 1 70385
0 9403 7 1 2 50648 70388
0 9404 5 2 1 9403
0 9405 7 14 2 52075 50649
0 9406 5 3 1 70409
0 9407 7 3 2 55672 60485
0 9408 5 1 1 70426
0 9409 7 1 2 70423 9408
0 9410 5 1 1 9409
0 9411 7 1 2 51851 9410
0 9412 5 1 1 9411
0 9413 7 1 2 70407 9412
0 9414 5 1 1 9413
0 9415 7 1 2 50373 9414
0 9416 5 1 1 9415
0 9417 7 1 2 9398 9416
0 9418 7 1 2 9396 9417
0 9419 5 2 1 9418
0 9420 7 1 2 67837 70429
0 9421 5 1 1 9420
0 9422 7 9 2 52231 56609
0 9423 5 1 1 70431
0 9424 7 14 2 50148 55673
0 9425 5 1 1 70440
0 9426 7 3 2 70432 70441
0 9427 5 1 1 70454
0 9428 7 4 2 55482 69643
0 9429 7 5 2 51852 54222
0 9430 5 1 1 70461
0 9431 7 7 2 53057 54555
0 9432 7 2 2 70462 70466
0 9433 5 1 1 70473
0 9434 7 1 2 70457 70474
0 9435 5 1 1 9434
0 9436 7 5 2 49861 50374
0 9437 5 1 1 70475
0 9438 7 1 2 52772 70476
0 9439 5 1 1 9438
0 9440 7 1 2 9435 9439
0 9441 5 1 1 9440
0 9442 7 1 2 70455 9441
0 9443 5 1 1 9442
0 9444 7 1 2 9421 9443
0 9445 5 1 1 9444
0 9446 7 1 2 62946 9445
0 9447 5 1 1 9446
0 9448 7 1 2 61442 63427
0 9449 5 8 1 9448
0 9450 7 1 2 53659 66968
0 9451 7 2 2 70480 9450
0 9452 7 1 2 59648 59773
0 9453 5 1 1 9452
0 9454 7 1 2 63622 9453
0 9455 5 1 1 9454
0 9456 7 1 2 51853 9455
0 9457 5 1 1 9456
0 9458 7 1 2 54556 60458
0 9459 5 3 1 9458
0 9460 7 5 2 50149 57206
0 9461 5 5 1 70493
0 9462 7 4 2 54223 70498
0 9463 5 3 1 70503
0 9464 7 1 2 50650 70507
0 9465 5 1 1 9464
0 9466 7 1 2 60041 9465
0 9467 5 1 1 9466
0 9468 7 1 2 70490 9467
0 9469 5 1 1 9468
0 9470 7 1 2 9457 9469
0 9471 5 1 1 9470
0 9472 7 1 2 52232 9471
0 9473 5 1 1 9472
0 9474 7 4 2 56610 70442
0 9475 5 1 1 70510
0 9476 7 1 2 59649 70511
0 9477 5 2 1 9476
0 9478 7 2 2 65018 59748
0 9479 5 1 1 70516
0 9480 7 1 2 55674 60011
0 9481 5 1 1 9480
0 9482 7 1 2 70517 9481
0 9483 5 1 1 9482
0 9484 7 1 2 52937 9483
0 9485 5 1 1 9484
0 9486 7 3 2 53058 60333
0 9487 5 1 1 70518
0 9488 7 1 2 51854 9479
0 9489 5 1 1 9488
0 9490 7 3 2 60232 9489
0 9491 5 1 1 70521
0 9492 7 1 2 9487 70522
0 9493 7 1 2 9485 9492
0 9494 5 1 1 9493
0 9495 7 1 2 50651 9494
0 9496 5 1 1 9495
0 9497 7 1 2 70514 9496
0 9498 7 1 2 9473 9497
0 9499 5 1 1 9498
0 9500 7 1 2 70488 9499
0 9501 5 1 1 9500
0 9502 7 1 2 9447 9501
0 9503 5 1 1 9502
0 9504 7 1 2 61328 9503
0 9505 5 1 1 9504
0 9506 7 2 2 49862 64379
0 9507 5 3 1 70524
0 9508 7 1 2 49700 65724
0 9509 5 2 1 9508
0 9510 7 1 2 70526 70529
0 9511 5 1 1 9510
0 9512 7 1 2 9511 70430
0 9513 5 1 1 9512
0 9514 7 1 2 61624 67716
0 9515 5 1 1 9514
0 9516 7 1 2 9437 9515
0 9517 5 1 1 9516
0 9518 7 1 2 64380 9517
0 9519 5 1 1 9518
0 9520 7 5 2 49701 50375
0 9521 5 2 1 70531
0 9522 7 1 2 70536 9433
0 9523 5 1 1 9522
0 9524 7 1 2 65725 9523
0 9525 5 1 1 9524
0 9526 7 1 2 9519 9525
0 9527 5 1 1 9526
0 9528 7 4 2 52880 50150
0 9529 5 1 1 70538
0 9530 7 3 2 62095 70539
0 9531 7 2 2 60468 70542
0 9532 7 1 2 9527 70545
0 9533 5 1 1 9532
0 9534 7 1 2 9513 9533
0 9535 5 1 1 9534
0 9536 7 1 2 56180 9535
0 9537 5 1 1 9536
0 9538 7 2 2 62947 58671
0 9539 7 1 2 70458 70547
0 9540 7 1 2 70347 9539
0 9541 5 2 1 9540
0 9542 7 1 2 9537 70549
0 9543 5 1 1 9542
0 9544 7 1 2 56437 9543
0 9545 5 1 1 9544
0 9546 7 1 2 50376 70489
0 9547 5 1 1 9546
0 9548 7 4 2 50377 62948
0 9549 7 1 2 67838 70551
0 9550 5 1 1 9549
0 9551 7 1 2 70550 9550
0 9552 7 1 2 9547 9551
0 9553 5 1 1 9552
0 9554 7 1 2 56181 9553
0 9555 5 1 1 9554
0 9556 7 5 2 69644 70098
0 9557 5 1 1 70555
0 9558 7 1 2 55483 58672
0 9559 7 1 2 70556 9558
0 9560 5 1 1 9559
0 9561 7 1 2 9555 9560
0 9562 5 1 1 9561
0 9563 7 1 2 57984 9562
0 9564 5 1 1 9563
0 9565 7 4 2 48896 68748
0 9566 5 4 1 70560
0 9567 7 1 2 49863 63062
0 9568 5 1 1 9567
0 9569 7 1 2 70564 9568
0 9570 5 4 1 9569
0 9571 7 1 2 61329 70568
0 9572 5 1 1 9571
0 9573 7 2 2 70162 70525
0 9574 5 1 1 70572
0 9575 7 1 2 9572 9574
0 9576 5 2 1 9575
0 9577 7 1 2 59845 70574
0 9578 7 1 2 70322 9577
0 9579 5 1 1 9578
0 9580 7 5 2 53444 67852
0 9581 5 1 1 70576
0 9582 7 1 2 58741 70577
0 9583 5 2 1 9582
0 9584 7 1 2 67844 70530
0 9585 5 3 1 9584
0 9586 7 13 2 52479 52597
0 9587 5 1 1 70586
0 9588 7 15 2 53265 70587
0 9589 7 1 2 70583 70599
0 9590 5 1 1 9589
0 9591 7 4 2 48713 52773
0 9592 7 1 2 65726 70614
0 9593 5 1 1 9592
0 9594 7 1 2 9590 9593
0 9595 7 1 2 70581 9594
0 9596 5 1 1 9595
0 9597 7 1 2 58714 9596
0 9598 5 1 1 9597
0 9599 7 1 2 9579 9598
0 9600 7 1 2 9564 9599
0 9601 7 1 2 9545 9600
0 9602 7 1 2 9505 9601
0 9603 5 1 1 9602
0 9604 7 1 2 50952 9603
0 9605 5 1 1 9604
0 9606 7 1 2 9376 9605
0 9607 5 1 1 9606
0 9608 7 1 2 69205 9607
0 9609 5 1 1 9608
0 9610 7 4 2 53158 66024
0 9611 5 3 1 70618
0 9612 7 1 2 49303 56344
0 9613 5 3 1 9612
0 9614 7 2 2 59483 70625
0 9615 5 1 1 70628
0 9616 7 1 2 52233 58645
0 9617 7 1 2 70629 9616
0 9618 5 1 1 9617
0 9619 7 1 2 70622 9618
0 9620 5 1 1 9619
0 9621 7 1 2 59927 9620
0 9622 5 1 1 9621
0 9623 7 1 2 66058 9622
0 9624 5 1 1 9623
0 9625 7 1 2 59846 9624
0 9626 5 1 1 9625
0 9627 7 5 2 52076 56182
0 9628 7 1 2 59793 70630
0 9629 5 1 1 9628
0 9630 7 15 2 59298 59090
0 9631 5 5 1 70635
0 9632 7 3 2 51855 58887
0 9633 5 1 1 70655
0 9634 7 1 2 70650 9633
0 9635 5 1 1 9634
0 9636 7 1 2 56183 9635
0 9637 5 1 1 9636
0 9638 7 1 2 60044 70631
0 9639 5 1 1 9638
0 9640 7 1 2 60160 60110
0 9641 5 1 1 9640
0 9642 7 1 2 9639 9641
0 9643 5 1 1 9642
0 9644 7 1 2 51856 9643
0 9645 5 1 1 9644
0 9646 7 1 2 9637 9645
0 9647 5 1 1 9646
0 9648 7 1 2 50151 9647
0 9649 5 1 1 9648
0 9650 7 1 2 9629 9649
0 9651 7 1 2 9626 9650
0 9652 5 1 1 9651
0 9653 7 1 2 50953 9652
0 9654 5 1 1 9653
0 9655 7 7 2 52375 65473
0 9656 5 10 1 70658
0 9657 7 13 2 53059 50954
0 9658 5 3 1 70675
0 9659 7 6 2 52234 50152
0 9660 5 2 1 70691
0 9661 7 4 2 70676 70692
0 9662 5 1 1 70699
0 9663 7 1 2 50378 70700
0 9664 5 1 1 9663
0 9665 7 1 2 56546 9664
0 9666 5 1 1 9665
0 9667 7 3 2 54224 60005
0 9668 5 2 1 70703
0 9669 7 1 2 70360 70704
0 9670 7 1 2 60879 9669
0 9671 5 1 1 9670
0 9672 7 1 2 9666 9671
0 9673 5 1 1 9672
0 9674 7 1 2 70665 9673
0 9675 5 1 1 9674
0 9676 7 1 2 50652 9675
0 9677 5 1 1 9676
0 9678 7 1 2 55675 63119
0 9679 5 1 1 9678
0 9680 7 2 2 56057 9679
0 9681 5 2 1 70708
0 9682 7 1 2 47849 60452
0 9683 5 1 1 9682
0 9684 7 2 2 70710 9683
0 9685 5 1 1 70712
0 9686 7 1 2 70239 70713
0 9687 5 1 1 9686
0 9688 7 1 2 54929 9687
0 9689 7 2 2 53990 61052
0 9690 5 14 1 70714
0 9691 7 2 2 57577 70716
0 9692 7 1 2 50379 70730
0 9693 5 1 1 9692
0 9694 7 1 2 60613 9693
0 9695 5 1 1 9694
0 9696 7 1 2 61178 9695
0 9697 5 1 1 9696
0 9698 7 13 2 61071 63229
0 9699 5 2 1 70732
0 9700 7 6 2 52077 55676
0 9701 5 4 1 70747
0 9702 7 1 2 70733 70748
0 9703 5 1 1 9702
0 9704 7 1 2 48342 59749
0 9705 5 4 1 9704
0 9706 7 2 2 50380 70757
0 9707 5 1 1 70761
0 9708 7 1 2 60062 70762
0 9709 5 1 1 9708
0 9710 7 1 2 9703 9709
0 9711 5 1 1 9710
0 9712 7 1 2 52938 9711
0 9713 5 1 1 9712
0 9714 7 1 2 9697 9713
0 9715 7 1 2 9688 9714
0 9716 5 1 1 9715
0 9717 7 1 2 56438 9716
0 9718 5 1 1 9717
0 9719 7 1 2 9677 9718
0 9720 5 1 1 9719
0 9721 7 1 2 53445 9720
0 9722 5 1 1 9721
0 9723 7 1 2 48343 70688
0 9724 5 2 1 9723
0 9725 7 6 2 53060 53159
0 9726 5 1 1 70765
0 9727 7 3 2 52376 70766
0 9728 5 1 1 70771
0 9729 7 1 2 54930 9728
0 9730 5 9 1 9729
0 9731 7 5 2 70763 70774
0 9732 7 2 2 61516 55677
0 9733 5 5 1 70788
0 9734 7 2 2 50153 59847
0 9735 5 1 1 70795
0 9736 7 1 2 59827 9735
0 9737 5 1 1 9736
0 9738 7 1 2 52078 9737
0 9739 5 1 1 9738
0 9740 7 3 2 70790 9739
0 9741 5 7 1 70797
0 9742 7 1 2 70783 70800
0 9743 5 1 1 9742
0 9744 7 7 2 50955 55849
0 9745 5 1 1 70807
0 9746 7 1 2 61606 63710
0 9747 5 1 1 9746
0 9748 7 1 2 70808 9747
0 9749 5 1 1 9748
0 9750 7 1 2 9743 9749
0 9751 5 1 1 9750
0 9752 7 1 2 50653 9751
0 9753 5 1 1 9752
0 9754 7 7 2 50956 56184
0 9755 5 1 1 70814
0 9756 7 3 2 51857 70389
0 9757 5 4 1 70821
0 9758 7 2 2 63230 63100
0 9759 5 2 1 70828
0 9760 7 2 2 70824 70830
0 9761 5 1 1 70832
0 9762 7 1 2 57428 60662
0 9763 5 1 1 9762
0 9764 7 1 2 57207 9763
0 9765 5 1 1 9764
0 9766 7 1 2 70833 9765
0 9767 5 1 1 9766
0 9768 7 1 2 70815 9767
0 9769 5 1 1 9768
0 9770 7 1 2 9753 9769
0 9771 5 1 1 9770
0 9772 7 1 2 50381 9771
0 9773 5 1 1 9772
0 9774 7 1 2 9722 9773
0 9775 7 1 2 9654 9774
0 9776 5 1 1 9775
0 9777 7 1 2 61213 9776
0 9778 5 1 1 9777
0 9779 7 4 2 52377 65293
0 9780 5 5 1 70834
0 9781 7 1 2 63389 70433
0 9782 5 2 1 9781
0 9783 7 1 2 70838 70843
0 9784 5 1 1 9783
0 9785 7 1 2 51858 9784
0 9786 5 2 1 9785
0 9787 7 3 2 59739 58319
0 9788 5 4 1 70847
0 9789 7 1 2 56345 70850
0 9790 5 3 1 9789
0 9791 7 1 2 61268 70499
0 9792 5 1 1 9791
0 9793 7 1 2 56185 9792
0 9794 5 1 1 9793
0 9795 7 1 2 61463 9794
0 9796 5 1 1 9795
0 9797 7 1 2 70854 9796
0 9798 5 1 1 9797
0 9799 7 1 2 70845 9798
0 9800 5 1 1 9799
0 9801 7 1 2 50654 9800
0 9802 5 1 1 9801
0 9803 7 1 2 54931 9802
0 9804 5 1 1 9803
0 9805 7 10 2 60766 57274
0 9806 5 1 1 70857
0 9807 7 1 2 60436 70858
0 9808 5 1 1 9807
0 9809 7 1 2 53061 9808
0 9810 5 1 1 9809
0 9811 7 1 2 50154 58320
0 9812 5 1 1 9811
0 9813 7 1 2 59477 9812
0 9814 7 1 2 9810 9813
0 9815 5 1 1 9814
0 9816 7 1 2 9804 9815
0 9817 5 1 1 9816
0 9818 7 1 2 50957 62240
0 9819 5 1 1 9818
0 9820 7 1 2 56186 70711
0 9821 5 1 1 9820
0 9822 7 1 2 9819 9821
0 9823 5 1 1 9822
0 9824 7 1 2 70240 9823
0 9825 5 1 1 9824
0 9826 7 4 2 52235 56187
0 9827 5 3 1 70867
0 9828 7 1 2 54932 70871
0 9829 5 4 1 9828
0 9830 7 1 2 70268 70874
0 9831 5 1 1 9830
0 9832 7 2 2 52378 58815
0 9833 7 1 2 66347 70878
0 9834 5 1 1 9833
0 9835 7 1 2 52236 59873
0 9836 5 1 1 9835
0 9837 7 1 2 9834 9836
0 9838 7 1 2 9831 9837
0 9839 5 1 1 9838
0 9840 7 1 2 61179 9839
0 9841 5 1 1 9840
0 9842 7 1 2 9825 9841
0 9843 5 1 1 9842
0 9844 7 1 2 51859 9843
0 9845 5 1 1 9844
0 9846 7 2 2 52237 59848
0 9847 5 2 1 70880
0 9848 7 1 2 48135 70882
0 9849 5 1 1 9848
0 9850 7 10 2 52379 50155
0 9851 5 2 1 70884
0 9852 7 1 2 66348 70885
0 9853 5 2 1 9852
0 9854 7 1 2 70689 70896
0 9855 5 2 1 9854
0 9856 7 4 2 52881 59816
0 9857 5 1 1 70900
0 9858 7 2 2 48344 9857
0 9859 5 4 1 70904
0 9860 7 1 2 70898 70906
0 9861 7 1 2 9849 9860
0 9862 5 1 1 9861
0 9863 7 2 2 57275 70500
0 9864 5 1 1 70910
0 9865 7 1 2 55737 70911
0 9866 5 1 1 9865
0 9867 7 3 2 60757 61863
0 9868 5 2 1 70912
0 9869 7 1 2 48345 60233
0 9870 5 3 1 9869
0 9871 7 1 2 70775 70917
0 9872 7 1 2 70913 9871
0 9873 7 1 2 9866 9872
0 9874 5 1 1 9873
0 9875 7 1 2 9862 9874
0 9876 7 1 2 9845 9875
0 9877 7 1 2 9817 9876
0 9878 5 1 1 9877
0 9879 7 1 2 53446 9878
0 9880 5 1 1 9879
0 9881 7 1 2 51860 70519
0 9882 5 1 1 9881
0 9883 7 1 2 60799 9882
0 9884 5 2 1 9883
0 9885 7 1 2 52238 70920
0 9886 5 1 1 9885
0 9887 7 2 2 60262 59650
0 9888 5 1 1 70922
0 9889 7 1 2 9886 9888
0 9890 5 2 1 9889
0 9891 7 1 2 59849 70924
0 9892 5 2 1 9891
0 9893 7 1 2 60621 60141
0 9894 5 1 1 9893
0 9895 7 1 2 60614 9894
0 9896 5 1 1 9895
0 9897 7 1 2 55678 9896
0 9898 5 1 1 9897
0 9899 7 1 2 67462 9898
0 9900 5 1 1 9899
0 9901 7 1 2 52939 9900
0 9902 5 1 1 9901
0 9903 7 1 2 60115 61296
0 9904 5 1 1 9903
0 9905 7 1 2 9902 9904
0 9906 7 1 2 70926 9905
0 9907 5 1 1 9906
0 9908 7 1 2 65484 9907
0 9909 5 1 1 9908
0 9910 7 1 2 9880 9909
0 9911 5 1 1 9910
0 9912 7 1 2 57985 9911
0 9913 5 1 1 9912
0 9914 7 1 2 49864 9913
0 9915 7 1 2 9778 9914
0 9916 5 1 1 9915
0 9917 7 1 2 53660 63567
0 9918 5 2 1 9917
0 9919 7 1 2 52598 69556
0 9920 7 1 2 70928 9919
0 9921 7 1 2 9916 9920
0 9922 5 1 1 9921
0 9923 7 1 2 64045 56990
0 9924 5 1 1 9923
0 9925 7 3 2 53062 56991
0 9926 5 3 1 70930
0 9927 7 6 2 52239 56992
0 9928 5 1 1 70936
0 9929 7 7 2 70933 9928
0 9930 5 3 1 70942
0 9931 7 1 2 63449 70943
0 9932 7 1 2 9924 9931
0 9933 5 1 1 9932
0 9934 7 1 2 52599 9933
0 9935 5 1 1 9934
0 9936 7 1 2 68821 9935
0 9937 5 1 1 9936
0 9938 7 1 2 62896 70118
0 9939 5 7 1 9938
0 9940 7 1 2 56697 63496
0 9941 5 1 1 9940
0 9942 7 1 2 50655 9941
0 9943 5 1 1 9942
0 9944 7 1 2 50656 60847
0 9945 5 2 1 9944
0 9946 7 2 2 60615 70959
0 9947 5 1 1 70961
0 9948 7 1 2 60672 70962
0 9949 5 1 1 9948
0 9950 7 1 2 57208 9949
0 9951 5 1 1 9950
0 9952 7 1 2 9943 9951
0 9953 7 2 2 60830 9952
0 9954 5 2 1 70963
0 9955 7 1 2 54933 70964
0 9956 5 1 1 9955
0 9957 7 1 2 70952 9956
0 9958 5 1 1 9957
0 9959 7 2 2 50156 61330
0 9960 5 1 1 70967
0 9961 7 2 2 60528 70968
0 9962 5 1 1 70969
0 9963 7 1 2 62425 70297
0 9964 7 1 2 70970 9963
0 9965 5 1 1 9964
0 9966 7 2 2 70179 9965
0 9967 7 1 2 9958 70971
0 9968 7 2 2 50382 60063
0 9969 5 2 1 70973
0 9970 7 1 2 59750 60500
0 9971 5 2 1 9970
0 9972 7 1 2 51861 70977
0 9973 5 2 1 9972
0 9974 7 3 2 70975 70979
0 9975 7 1 2 52240 70706
0 9976 5 1 1 9975
0 9977 7 1 2 70981 9976
0 9978 5 1 1 9977
0 9979 7 1 2 61331 9978
0 9980 5 1 1 9979
0 9981 7 1 2 63759 65217
0 9982 5 2 1 9981
0 9983 7 4 2 50657 55679
0 9984 7 1 2 54225 61634
0 9985 5 4 1 9984
0 9986 7 2 2 50157 70990
0 9987 7 1 2 70986 70994
0 9988 5 1 1 9987
0 9989 7 1 2 70984 9988
0 9990 5 1 1 9989
0 9991 7 1 2 52241 9990
0 9992 5 1 1 9991
0 9993 7 1 2 9980 9992
0 9994 5 1 1 9993
0 9995 7 1 2 57209 9994
0 9996 5 1 1 9995
0 9997 7 7 2 55850 56611
0 9998 5 7 1 70996
0 9999 7 1 2 60663 70636
0 10000 5 1 1 9999
0 10001 7 1 2 71003 10000
0 10002 5 1 1 10001
0 10003 7 1 2 50383 10002
0 10004 5 1 1 10003
0 10005 7 10 2 50158 55851
0 10006 5 3 1 71010
0 10007 7 2 2 61246 71011
0 10008 5 2 1 71023
0 10009 7 1 2 57210 63392
0 10010 5 1 1 10009
0 10011 7 1 2 71025 10010
0 10012 7 1 2 10004 10011
0 10013 5 1 1 10012
0 10014 7 1 2 50658 10013
0 10015 5 1 1 10014
0 10016 7 1 2 9996 10015
0 10017 5 1 1 10016
0 10018 7 1 2 50958 10017
0 10019 5 1 1 10018
0 10020 7 3 2 54226 60834
0 10021 5 4 1 71027
0 10022 7 1 2 53063 71030
0 10023 5 1 1 10022
0 10024 7 1 2 60792 10023
0 10025 5 1 1 10024
0 10026 7 1 2 50959 10025
0 10027 5 1 1 10026
0 10028 7 2 2 50659 60664
0 10029 7 3 2 59651 56612
0 10030 5 1 1 71036
0 10031 7 2 2 71034 71037
0 10032 5 1 1 71039
0 10033 7 1 2 10027 10032
0 10034 5 1 1 10033
0 10035 7 1 2 52242 10034
0 10036 5 1 1 10035
0 10037 7 1 2 53064 60789
0 10038 5 1 1 10037
0 10039 7 2 2 54557 60817
0 10040 5 5 1 71041
0 10041 7 2 2 51862 60887
0 10042 5 3 1 71048
0 10043 7 1 2 60722 71049
0 10044 5 1 1 10043
0 10045 7 1 2 71042 10044
0 10046 7 1 2 10038 10045
0 10047 5 1 1 10046
0 10048 7 1 2 50960 10047
0 10049 5 1 1 10048
0 10050 7 1 2 62897 10049
0 10051 7 1 2 10036 10050
0 10052 5 1 1 10051
0 10053 7 1 2 56346 62999
0 10054 5 1 1 10053
0 10055 7 1 2 10052 10054
0 10056 5 1 1 10055
0 10057 7 1 2 10019 10056
0 10058 7 1 2 9967 10057
0 10059 5 1 1 10058
0 10060 7 1 2 49865 10059
0 10061 5 1 1 10060
0 10062 7 1 2 9937 10061
0 10063 5 1 1 10062
0 10064 7 1 2 52774 10063
0 10065 5 1 1 10064
0 10066 7 1 2 60354 67114
0 10067 5 1 1 10066
0 10068 7 1 2 54227 60605
0 10069 5 3 1 10068
0 10070 7 5 2 50961 70123
0 10071 7 1 2 71053 71056
0 10072 5 1 1 10071
0 10073 7 7 2 53266 50384
0 10074 5 1 1 71061
0 10075 7 2 2 70142 71062
0 10076 5 1 1 71068
0 10077 7 1 2 66039 71069
0 10078 5 1 1 10077
0 10079 7 1 2 10072 10078
0 10080 5 1 1 10079
0 10081 7 3 2 53065 49866
0 10082 7 1 2 71070 70901
0 10083 7 1 2 10080 10082
0 10084 5 1 1 10083
0 10085 7 1 2 10067 10084
0 10086 5 1 1 10085
0 10087 7 1 2 50660 10086
0 10088 5 1 1 10087
0 10089 7 12 2 49867 50962
0 10090 7 2 2 53160 71073
0 10091 7 9 2 52243 52380
0 10092 7 2 2 56439 71087
0 10093 7 1 2 71085 71096
0 10094 5 1 1 10093
0 10095 7 2 2 59774 67115
0 10096 5 1 1 71098
0 10097 7 1 2 53066 71099
0 10098 5 1 1 10097
0 10099 7 1 2 10094 10098
0 10100 5 1 1 10099
0 10101 7 1 2 51863 10100
0 10102 5 1 1 10101
0 10103 7 2 2 49868 56440
0 10104 7 1 2 70816 71100
0 10105 5 2 1 10104
0 10106 7 1 2 52244 67116
0 10107 5 1 1 10106
0 10108 7 1 2 71102 10107
0 10109 5 2 1 10108
0 10110 7 1 2 54228 58824
0 10111 5 1 1 10110
0 10112 7 1 2 71104 10111
0 10113 5 1 1 10112
0 10114 7 1 2 48897 68716
0 10115 5 2 1 10114
0 10116 7 9 2 53267 50963
0 10117 5 4 1 71108
0 10118 7 4 2 70102 71109
0 10119 5 2 1 71121
0 10120 7 2 2 49869 71122
0 10121 7 1 2 60469 71127
0 10122 5 1 1 10121
0 10123 7 1 2 71106 10122
0 10124 7 1 2 10113 10123
0 10125 7 1 2 10102 10124
0 10126 5 1 1 10125
0 10127 7 1 2 52079 10126
0 10128 5 1 1 10127
0 10129 7 1 2 51864 71105
0 10130 5 1 1 10129
0 10131 7 1 2 48898 68478
0 10132 5 1 1 10131
0 10133 7 1 2 10130 10132
0 10134 5 1 1 10133
0 10135 7 1 2 52080 10134
0 10136 5 1 1 10135
0 10137 7 1 2 58321 69307
0 10138 7 1 2 71057 10137
0 10139 5 1 1 10138
0 10140 7 1 2 10136 10139
0 10141 5 1 1 10140
0 10142 7 1 2 60045 10141
0 10143 5 1 1 10142
0 10144 7 3 2 52245 59635
0 10145 5 1 1 71129
0 10146 7 4 2 59673 10145
0 10147 5 2 1 71132
0 10148 7 1 2 71136 71128
0 10149 5 1 1 10148
0 10150 7 1 2 10143 10149
0 10151 7 1 2 10128 10150
0 10152 7 1 2 10088 10151
0 10153 5 1 1 10152
0 10154 7 1 2 53447 10153
0 10155 5 1 1 10154
0 10156 7 5 2 59691 70991
0 10157 5 1 1 71138
0 10158 7 3 2 50964 67117
0 10159 7 18 2 52940 50661
0 10160 5 5 1 71146
0 10161 7 3 2 55680 71147
0 10162 7 1 2 71143 71169
0 10163 7 1 2 71139 10162
0 10164 5 1 1 10163
0 10165 7 1 2 10155 10164
0 10166 5 1 1 10165
0 10167 7 1 2 50159 10166
0 10168 5 1 1 10167
0 10169 7 7 2 52081 50965
0 10170 5 1 1 71172
0 10171 7 1 2 67132 70119
0 10172 5 1 1 10171
0 10173 7 1 2 67133 68816
0 10174 5 3 1 10173
0 10175 7 1 2 50662 71179
0 10176 7 2 2 10172 10175
0 10177 7 1 2 71173 71182
0 10178 5 1 1 10177
0 10179 7 1 2 70565 10178
0 10180 5 1 1 10179
0 10181 7 1 2 59775 10180
0 10182 5 1 1 10181
0 10183 7 1 2 71123 68798
0 10184 5 1 1 10183
0 10185 7 1 2 10182 10184
0 10186 5 1 1 10185
0 10187 7 1 2 51865 10186
0 10188 5 1 1 10187
0 10189 7 11 2 53161 70143
0 10190 7 1 2 53268 68799
0 10191 7 3 2 71184 10190
0 10192 7 1 2 66715 71195
0 10193 5 1 1 10192
0 10194 7 1 2 10188 10193
0 10195 5 1 1 10194
0 10196 7 1 2 50385 10195
0 10197 5 1 1 10196
0 10198 7 6 2 52381 52941
0 10199 5 1 1 71198
0 10200 7 2 2 60772 71199
0 10201 7 5 2 50086 50966
0 10202 7 2 2 53162 71206
0 10203 7 1 2 71211 71101
0 10204 7 1 2 71204 10203
0 10205 5 1 1 10204
0 10206 7 1 2 71107 10205
0 10207 5 1 1 10206
0 10208 7 1 2 53448 10207
0 10209 5 1 1 10208
0 10210 7 1 2 10197 10209
0 10211 5 1 1 10210
0 10212 7 1 2 57578 10211
0 10213 5 1 1 10212
0 10214 7 4 2 53269 50087
0 10215 7 2 2 60164 71213
0 10216 5 1 1 71217
0 10217 7 1 2 54934 10216
0 10218 5 1 1 10217
0 10219 7 1 2 65218 58888
0 10220 7 1 2 10218 10219
0 10221 5 1 1 10220
0 10222 7 7 2 52942 53270
0 10223 5 1 1 71219
0 10224 7 5 2 52882 71207
0 10225 5 2 1 71226
0 10226 7 1 2 71220 71227
0 10227 5 1 1 10226
0 10228 7 1 2 10221 10227
0 10229 5 1 1 10228
0 10230 7 1 2 51866 10229
0 10231 5 1 1 10230
0 10232 7 5 2 50663 56613
0 10233 5 2 1 71233
0 10234 7 1 2 49535 71238
0 10235 5 4 1 10234
0 10236 7 1 2 70809 71240
0 10237 5 1 1 10236
0 10238 7 1 2 10231 10237
0 10239 5 1 1 10238
0 10240 7 1 2 70103 10239
0 10241 5 1 1 10240
0 10242 7 4 2 55852 57310
0 10243 5 3 1 71244
0 10244 7 2 2 60355 59126
0 10245 7 7 2 52082 53271
0 10246 5 1 1 71253
0 10247 7 1 2 71251 71254
0 10248 7 1 2 71245 10247
0 10249 5 1 1 10248
0 10250 7 1 2 10241 10249
0 10251 5 1 1 10250
0 10252 7 1 2 49870 10251
0 10253 5 1 1 10252
0 10254 7 3 2 48899 53067
0 10255 7 3 2 52246 53661
0 10256 7 2 2 71260 71263
0 10257 5 2 1 71266
0 10258 7 1 2 61485 71267
0 10259 5 1 1 10258
0 10260 7 1 2 10253 10259
0 10261 5 1 1 10260
0 10262 7 1 2 50386 10261
0 10263 5 1 1 10262
0 10264 7 1 2 71103 10096
0 10265 5 1 1 10264
0 10266 7 1 2 70319 10265
0 10267 5 1 1 10266
0 10268 7 1 2 51867 60622
0 10269 5 2 1 10268
0 10270 7 1 2 54558 71270
0 10271 5 2 1 10270
0 10272 7 1 2 67118 71272
0 10273 5 1 1 10272
0 10274 7 4 2 52382 60187
0 10275 5 1 1 71274
0 10276 7 2 2 62353 71275
0 10277 5 2 1 71278
0 10278 7 5 2 52480 53068
0 10279 5 1 1 71282
0 10280 7 3 2 52247 53272
0 10281 7 4 2 71283 71287
0 10282 7 1 2 49871 71290
0 10283 7 1 2 71279 10282
0 10284 5 1 1 10283
0 10285 7 1 2 10273 10284
0 10286 5 1 1 10285
0 10287 7 1 2 52083 10286
0 10288 5 1 1 10287
0 10289 7 3 2 50160 67119
0 10290 7 1 2 71140 71294
0 10291 5 1 1 10290
0 10292 7 1 2 10288 10291
0 10293 5 1 1 10292
0 10294 7 1 2 59850 10293
0 10295 5 1 1 10294
0 10296 7 1 2 10267 10295
0 10297 7 1 2 10263 10296
0 10298 5 1 1 10297
0 10299 7 1 2 53449 10298
0 10300 5 1 1 10299
0 10301 7 1 2 71183 70925
0 10302 5 1 1 10301
0 10303 7 2 2 52248 60012
0 10304 5 1 1 71297
0 10305 7 1 2 70523 10304
0 10306 5 1 1 10305
0 10307 7 1 2 71196 10306
0 10308 5 1 1 10307
0 10309 7 1 2 10302 10308
0 10310 5 1 1 10309
0 10311 7 1 2 50967 59851
0 10312 7 1 2 10310 10311
0 10313 5 1 1 10312
0 10314 7 1 2 49702 59160
0 10315 5 1 1 10314
0 10316 7 3 2 52249 52600
0 10317 7 3 2 66025 71299
0 10318 7 5 2 49872 50161
0 10319 7 1 2 66349 71305
0 10320 7 1 2 71302 10319
0 10321 5 1 1 10320
0 10322 7 1 2 67134 10321
0 10323 5 1 1 10322
0 10324 7 1 2 57986 10323
0 10325 5 1 1 10324
0 10326 7 4 2 49873 70600
0 10327 5 3 1 71310
0 10328 7 1 2 67135 71314
0 10329 5 3 1 10328
0 10330 7 1 2 70855 71317
0 10331 5 1 1 10330
0 10332 7 1 2 10325 10331
0 10333 5 1 1 10332
0 10334 7 1 2 10315 10333
0 10335 5 1 1 10334
0 10336 7 4 2 53662 55853
0 10337 7 4 2 48900 50387
0 10338 5 1 1 71324
0 10339 7 1 2 52084 71325
0 10340 7 1 2 71320 10339
0 10341 7 1 2 71252 10340
0 10342 5 1 1 10341
0 10343 7 1 2 10335 10342
0 10344 7 1 2 10313 10343
0 10345 7 1 2 10300 10344
0 10346 7 1 2 10213 10345
0 10347 7 1 2 10168 10346
0 10348 7 1 2 10065 10347
0 10349 7 1 2 9922 10348
0 10350 5 1 1 10349
0 10351 7 1 2 68230 10350
0 10352 5 1 1 10351
0 10353 7 16 2 53663 50005
0 10354 5 2 1 71328
0 10355 7 4 2 49004 53450
0 10356 7 3 2 71329 71346
0 10357 7 4 2 64142 68689
0 10358 5 1 1 71353
0 10359 7 1 2 71350 71354
0 10360 5 1 1 10359
0 10361 7 5 2 61893 63716
0 10362 7 1 2 71351 71357
0 10363 5 1 1 10362
0 10364 7 1 2 49005 53778
0 10365 5 4 1 10364
0 10366 7 6 2 50162 59127
0 10367 5 2 1 71366
0 10368 7 3 2 53451 66885
0 10369 7 1 2 50006 71374
0 10370 7 1 2 71367 10369
0 10371 5 1 1 10370
0 10372 7 1 2 71362 10371
0 10373 5 1 1 10372
0 10374 7 2 2 49874 65613
0 10375 7 1 2 66783 71377
0 10376 7 1 2 10373 10375
0 10377 5 1 1 10376
0 10378 7 1 2 10363 10377
0 10379 5 1 1 10378
0 10380 7 1 2 58381 10379
0 10381 5 1 1 10380
0 10382 7 1 2 10360 10381
0 10383 5 1 1 10382
0 10384 7 1 2 57429 10383
0 10385 5 1 1 10384
0 10386 7 2 2 53452 69861
0 10387 7 8 2 54559 63717
0 10388 7 1 2 71330 71381
0 10389 7 1 2 71379 10388
0 10390 5 1 1 10389
0 10391 7 1 2 10385 10390
0 10392 5 1 1 10391
0 10393 7 1 2 58107 10392
0 10394 5 1 1 10393
0 10395 7 2 2 67030 68216
0 10396 5 1 1 71389
0 10397 7 1 2 68275 10396
0 10398 5 5 1 10397
0 10399 7 2 2 57894 71391
0 10400 5 1 1 71396
0 10401 7 3 2 49110 61657
0 10402 5 10 1 71398
0 10403 7 2 2 50664 71401
0 10404 5 1 1 71411
0 10405 7 1 2 57211 71412
0 10406 5 2 1 10405
0 10407 7 1 2 68299 71413
0 10408 5 1 1 10407
0 10409 7 11 2 50163 54560
0 10410 7 1 2 71415 68871
0 10411 7 1 2 60994 10410
0 10412 5 1 1 10411
0 10413 7 1 2 10408 10412
0 10414 5 1 1 10413
0 10415 7 1 2 57430 10414
0 10416 5 1 1 10415
0 10417 7 1 2 65543 68915
0 10418 5 1 1 10417
0 10419 7 1 2 10416 10418
0 10420 5 1 1 10419
0 10421 7 1 2 71397 10420
0 10422 5 1 1 10421
0 10423 7 2 2 50388 60356
0 10424 5 5 1 71426
0 10425 7 1 2 64035 68179
0 10426 7 1 2 71428 10425
0 10427 7 1 2 70226 10426
0 10428 5 1 1 10427
0 10429 7 3 2 48901 49006
0 10430 7 1 2 50007 71433
0 10431 7 1 2 10428 10430
0 10432 5 1 1 10431
0 10433 7 1 2 10422 10432
0 10434 5 1 1 10433
0 10435 7 1 2 53664 10434
0 10436 5 1 1 10435
0 10437 7 1 2 58322 70677
0 10438 5 3 1 10437
0 10439 7 1 2 57579 61332
0 10440 5 1 1 10439
0 10441 7 1 2 54935 10440
0 10442 5 1 1 10441
0 10443 7 1 2 63603 10442
0 10444 5 1 1 10443
0 10445 7 1 2 71436 10444
0 10446 5 1 1 10445
0 10447 7 1 2 51868 10446
0 10448 5 1 1 10447
0 10449 7 1 2 10448 9962
0 10450 5 1 1 10449
0 10451 7 1 2 61467 10450
0 10452 5 1 1 10451
0 10453 7 1 2 54936 67979
0 10454 5 1 1 10453
0 10455 7 3 2 59776 61591
0 10456 5 3 1 71439
0 10457 7 1 2 54561 71442
0 10458 5 2 1 10457
0 10459 7 1 2 71054 71445
0 10460 5 1 1 10459
0 10461 7 1 2 53069 61495
0 10462 5 1 1 10461
0 10463 7 3 2 60470 60773
0 10464 7 1 2 60492 71447
0 10465 5 1 1 10464
0 10466 7 1 2 10462 10465
0 10467 7 1 2 10460 10466
0 10468 5 1 1 10467
0 10469 7 1 2 50164 10468
0 10470 5 1 1 10469
0 10471 7 1 2 56614 61118
0 10472 5 1 1 10471
0 10473 7 2 2 49536 64039
0 10474 5 1 1 71450
0 10475 7 1 2 60631 71451
0 10476 7 1 2 10472 10475
0 10477 5 1 1 10476
0 10478 7 1 2 5792 10477
0 10479 5 1 1 10478
0 10480 7 1 2 49703 10479
0 10481 7 1 2 10470 10480
0 10482 5 1 1 10481
0 10483 7 1 2 10454 10482
0 10484 5 1 1 10483
0 10485 7 1 2 54937 70515
0 10486 5 1 1 10485
0 10487 7 1 2 52250 10486
0 10488 5 1 1 10487
0 10489 7 2 2 56698 63222
0 10490 5 1 1 71452
0 10491 7 1 2 60623 10490
0 10492 5 1 1 10491
0 10493 7 1 2 71004 10492
0 10494 7 1 2 70278 10493
0 10495 5 1 1 10494
0 10496 7 1 2 50665 10495
0 10497 5 1 1 10496
0 10498 7 1 2 10488 10497
0 10499 5 1 1 10498
0 10500 7 1 2 61333 10499
0 10501 5 1 1 10500
0 10502 7 1 2 10484 10501
0 10503 7 1 2 10452 10502
0 10504 5 1 1 10503
0 10505 7 1 2 52601 10504
0 10506 5 1 1 10505
0 10507 7 1 2 56547 62898
0 10508 5 11 1 10507
0 10509 7 2 2 53070 59874
0 10510 5 3 1 71465
0 10511 7 1 2 51869 62378
0 10512 5 1 1 10511
0 10513 7 1 2 71467 10512
0 10514 5 1 1 10513
0 10515 7 1 2 52251 10514
0 10516 5 1 1 10515
0 10517 7 2 2 50666 70776
0 10518 7 1 2 51870 71470
0 10519 5 1 1 10518
0 10520 7 1 2 10516 10519
0 10521 5 1 1 10520
0 10522 7 1 2 50389 10521
0 10523 5 1 1 10522
0 10524 7 1 2 70666 10523
0 10525 5 1 1 10524
0 10526 7 1 2 71454 10525
0 10527 5 1 1 10526
0 10528 7 5 2 50968 62949
0 10529 5 1 1 71472
0 10530 7 1 2 53453 57580
0 10531 5 2 1 10530
0 10532 7 3 2 52602 57581
0 10533 5 1 1 71479
0 10534 7 1 2 71477 10533
0 10535 5 2 1 10534
0 10536 7 1 2 61496 71482
0 10537 5 1 1 10536
0 10538 7 1 2 61507 59765
0 10539 5 4 1 10538
0 10540 7 1 2 71484 70817
0 10541 5 1 1 10540
0 10542 7 1 2 10537 10541
0 10543 5 1 1 10542
0 10544 7 1 2 50390 10543
0 10545 5 1 1 10544
0 10546 7 1 2 10529 10545
0 10547 5 1 1 10546
0 10548 7 1 2 57987 10547
0 10549 5 1 1 10548
0 10550 7 1 2 48902 70313
0 10551 5 3 1 10550
0 10552 7 1 2 70202 71488
0 10553 5 1 1 10552
0 10554 7 1 2 10549 10553
0 10555 7 1 2 10527 10554
0 10556 5 1 1 10555
0 10557 7 1 2 70213 10556
0 10558 5 1 1 10557
0 10559 7 7 2 50667 57212
0 10560 5 2 1 71491
0 10561 7 1 2 56188 71455
0 10562 5 1 1 10561
0 10563 7 1 2 67984 10562
0 10564 5 2 1 10563
0 10565 7 1 2 55854 71500
0 10566 5 1 1 10565
0 10567 7 2 2 59912 70953
0 10568 5 1 1 71502
0 10569 7 1 2 10566 10568
0 10570 5 1 1 10569
0 10571 7 1 2 71492 10570
0 10572 5 1 1 10571
0 10573 7 1 2 56615 71489
0 10574 5 1 1 10573
0 10575 7 1 2 10572 10574
0 10576 5 1 1 10575
0 10577 7 1 2 60848 10576
0 10578 5 1 1 10577
0 10579 7 1 2 57988 70875
0 10580 5 1 1 10579
0 10581 7 1 2 70667 10580
0 10582 5 1 1 10581
0 10583 7 1 2 62950 10582
0 10584 5 1 1 10583
0 10585 7 19 2 52603 56441
0 10586 5 4 1 71504
0 10587 7 2 2 48903 71523
0 10588 5 8 1 71527
0 10589 7 4 2 53454 58742
0 10590 5 2 1 71537
0 10591 7 1 2 71528 71541
0 10592 5 3 1 10591
0 10593 7 1 2 52252 71543
0 10594 5 1 1 10593
0 10595 7 1 2 71125 10594
0 10596 7 1 2 10584 10595
0 10597 5 1 1 10596
0 10598 7 1 2 65759 10597
0 10599 5 1 1 10598
0 10600 7 1 2 50391 64486
0 10601 5 2 1 10600
0 10602 7 2 2 53071 60414
0 10603 5 3 1 71548
0 10604 7 1 2 54562 71550
0 10605 7 1 2 71546 10604
0 10606 5 1 1 10605
0 10607 7 1 2 71490 10606
0 10608 5 1 1 10607
0 10609 7 2 2 64450 62899
0 10610 5 1 1 71553
0 10611 7 1 2 52775 10610
0 10612 5 1 1 10611
0 10613 7 3 2 50969 56442
0 10614 7 2 2 50165 60529
0 10615 5 6 1 71558
0 10616 7 1 2 49704 71560
0 10617 5 1 1 10616
0 10618 7 1 2 71555 10617
0 10619 5 1 1 10618
0 10620 7 1 2 10612 10619
0 10621 7 1 2 10608 10620
0 10622 7 1 2 10599 10621
0 10623 7 1 2 10578 10622
0 10624 7 1 2 10558 10623
0 10625 7 1 2 10506 10624
0 10626 7 2 2 53455 60530
0 10627 5 2 1 71566
0 10628 7 6 2 52253 66026
0 10629 7 2 2 53163 59875
0 10630 5 1 1 71576
0 10631 7 1 2 71570 71577
0 10632 5 1 1 10631
0 10633 7 1 2 71568 10632
0 10634 5 1 1 10633
0 10635 7 1 2 51871 10634
0 10636 5 1 1 10635
0 10637 7 2 2 65474 66027
0 10638 5 2 1 71578
0 10639 7 3 2 53072 53456
0 10640 5 1 1 71582
0 10641 7 1 2 70668 10640
0 10642 5 4 1 10641
0 10643 7 1 2 52254 71585
0 10644 5 1 1 10643
0 10645 7 1 2 71580 10644
0 10646 5 1 1 10645
0 10647 7 1 2 60188 10646
0 10648 5 1 1 10647
0 10649 7 1 2 10636 10648
0 10650 5 1 1 10649
0 10651 7 1 2 55681 10650
0 10652 5 1 1 10651
0 10653 7 1 2 71478 70669
0 10654 5 2 1 10653
0 10655 7 1 2 48346 70670
0 10656 5 1 1 10655
0 10657 7 1 2 53073 10656
0 10658 5 1 1 10657
0 10659 7 1 2 54229 10658
0 10660 5 1 1 10659
0 10661 7 1 2 71589 10660
0 10662 5 1 1 10661
0 10663 7 1 2 65475 71088
0 10664 5 3 1 10663
0 10665 7 1 2 10662 71591
0 10666 5 1 1 10665
0 10667 7 1 2 50668 10666
0 10668 5 1 1 10667
0 10669 7 1 2 10652 10668
0 10670 5 1 1 10669
0 10671 7 1 2 56616 10670
0 10672 5 1 1 10671
0 10673 7 3 2 53457 63604
0 10674 5 2 1 71594
0 10675 7 1 2 59652 70659
0 10676 5 1 1 10675
0 10677 7 1 2 71597 10676
0 10678 5 1 1 10677
0 10679 7 1 2 52255 10678
0 10680 5 1 1 10679
0 10681 7 2 2 50669 71586
0 10682 7 1 2 50166 71599
0 10683 5 1 1 10682
0 10684 7 1 2 10680 10683
0 10685 5 1 1 10684
0 10686 7 1 2 51872 10685
0 10687 5 1 1 10686
0 10688 7 1 2 50670 63693
0 10689 5 1 1 10688
0 10690 7 1 2 10687 10689
0 10691 5 1 1 10690
0 10692 7 1 2 61468 10691
0 10693 5 1 1 10692
0 10694 7 4 2 52256 50970
0 10695 5 1 1 71601
0 10696 7 1 2 53458 71602
0 10697 5 1 1 10696
0 10698 7 1 2 65800 70619
0 10699 5 1 1 10698
0 10700 7 1 2 49705 10699
0 10701 5 1 1 10700
0 10702 7 1 2 50971 10701
0 10703 5 1 1 10702
0 10704 7 1 2 63697 71581
0 10705 5 1 1 10704
0 10706 7 1 2 52257 10705
0 10707 5 1 1 10706
0 10708 7 1 2 65801 70918
0 10709 7 1 2 71587 10708
0 10710 5 1 1 10709
0 10711 7 1 2 10707 10710
0 10712 7 1 2 10703 10711
0 10713 5 1 1 10712
0 10714 7 1 2 50671 10713
0 10715 5 1 1 10714
0 10716 7 1 2 10697 10715
0 10717 7 1 2 10693 10716
0 10718 7 1 2 10672 10717
0 10719 5 1 1 10718
0 10720 7 1 2 57989 10719
0 10721 5 1 1 10720
0 10722 7 3 2 52383 50392
0 10723 5 3 1 71605
0 10724 7 2 2 62354 71606
0 10725 5 2 1 71611
0 10726 7 1 2 9662 71613
0 10727 5 1 1 10726
0 10728 7 1 2 51873 10727
0 10729 5 1 1 10728
0 10730 7 1 2 60189 70784
0 10731 5 1 1 10730
0 10732 7 1 2 10729 10731
0 10733 5 1 1 10732
0 10734 7 1 2 55682 10733
0 10735 5 1 1 10734
0 10736 7 1 2 59636 70876
0 10737 5 1 1 10736
0 10738 7 1 2 50393 70620
0 10739 5 1 1 10738
0 10740 7 1 2 10695 10739
0 10741 7 1 2 10737 10740
0 10742 5 1 1 10741
0 10743 7 1 2 50672 10742
0 10744 5 1 1 10743
0 10745 7 1 2 10735 10744
0 10746 5 1 1 10745
0 10747 7 1 2 56617 10746
0 10748 5 1 1 10747
0 10749 7 1 2 62355 70886
0 10750 5 2 1 10749
0 10751 7 1 2 50394 70678
0 10752 5 1 1 10751
0 10753 7 1 2 71615 10752
0 10754 5 1 1 10753
0 10755 7 1 2 52258 10754
0 10756 5 1 1 10755
0 10757 7 1 2 50167 71471
0 10758 5 1 1 10757
0 10759 7 1 2 10756 10758
0 10760 5 1 1 10759
0 10761 7 1 2 51874 10760
0 10762 5 1 1 10761
0 10763 7 1 2 10762 71280
0 10764 5 1 1 10763
0 10765 7 1 2 61469 10764
0 10766 5 1 1 10765
0 10767 7 1 2 65802 70785
0 10768 5 1 1 10767
0 10769 7 1 2 52259 70899
0 10770 5 2 1 10769
0 10771 7 5 2 53164 60190
0 10772 5 5 1 71619
0 10773 7 2 2 66028 71620
0 10774 5 2 1 71629
0 10775 7 1 2 71617 71631
0 10776 7 1 2 10768 10775
0 10777 5 1 1 10776
0 10778 7 1 2 50673 10777
0 10779 5 1 1 10778
0 10780 7 1 2 71592 10779
0 10781 7 1 2 10766 10780
0 10782 7 1 2 10748 10781
0 10783 5 1 1 10782
0 10784 7 1 2 61214 10783
0 10785 5 1 1 10784
0 10786 7 1 2 10721 10785
0 10787 7 1 2 10625 10786
0 10788 5 1 1 10787
0 10789 7 3 2 49007 49875
0 10790 7 1 2 50008 71633
0 10791 7 1 2 10788 10790
0 10792 5 1 1 10791
0 10793 7 1 2 10436 10792
0 10794 5 1 1 10793
0 10795 7 1 2 51249 10794
0 10796 5 1 1 10795
0 10797 7 1 2 10394 10796
0 10798 7 1 2 10352 10797
0 10799 5 1 1 10798
0 10800 7 1 2 51521 10799
0 10801 5 1 1 10800
0 10802 7 1 2 9609 10801
0 10803 5 1 1 10802
0 10804 7 1 2 55621 10803
0 10805 5 1 1 10804
0 10806 7 1 2 54230 68989
0 10807 5 1 1 10806
0 10808 7 1 2 61894 69344
0 10809 5 1 1 10808
0 10810 7 1 2 10807 10809
0 10811 5 1 1 10810
0 10812 7 1 2 57431 10811
0 10813 5 1 1 10812
0 10814 7 3 2 56865 63505
0 10815 5 1 1 71636
0 10816 7 1 2 66579 68455
0 10817 7 1 2 71637 10816
0 10818 5 1 1 10817
0 10819 7 1 2 69114 10818
0 10820 5 1 1 10819
0 10821 7 1 2 54231 10820
0 10822 5 1 1 10821
0 10823 7 1 2 10813 10822
0 10824 5 1 1 10823
0 10825 7 1 2 47850 10824
0 10826 5 1 1 10825
0 10827 7 1 2 66860 69340
0 10828 5 1 1 10827
0 10829 7 1 2 66701 68895
0 10830 5 1 1 10829
0 10831 7 1 2 10828 10830
0 10832 7 1 2 10826 10831
0 10833 5 1 1 10832
0 10834 7 1 2 51250 10833
0 10835 5 1 1 10834
0 10836 7 2 2 66268 68683
0 10837 7 1 2 49876 62008
0 10838 7 2 2 58228 10837
0 10839 7 1 2 71639 71641
0 10840 5 1 1 10839
0 10841 7 2 2 10835 10840
0 10842 5 1 1 71643
0 10843 7 1 2 51251 69110
0 10844 5 1 1 10843
0 10845 7 1 2 66580 69364
0 10846 5 1 1 10845
0 10847 7 1 2 47851 69281
0 10848 5 1 1 10847
0 10849 7 1 2 10846 10848
0 10850 5 1 1 10849
0 10851 7 1 2 49428 51522
0 10852 7 1 2 63345 10851
0 10853 7 1 2 10850 10852
0 10854 5 1 1 10853
0 10855 7 1 2 10844 10854
0 10856 5 1 1 10855
0 10857 7 1 2 56058 10856
0 10858 5 1 1 10857
0 10859 7 1 2 71644 10858
0 10860 5 1 1 10859
0 10861 7 1 2 58966 10860
0 10862 5 1 1 10861
0 10863 7 1 2 54563 69737
0 10864 5 1 1 10863
0 10865 7 1 2 57432 68355
0 10866 5 1 1 10865
0 10867 7 1 2 67797 10866
0 10868 5 1 1 10867
0 10869 7 1 2 57433 67765
0 10870 5 2 1 10869
0 10871 7 1 2 57754 71645
0 10872 5 1 1 10871
0 10873 7 1 2 53991 10872
0 10874 7 1 2 10868 10873
0 10875 5 1 1 10874
0 10876 7 3 2 49877 66520
0 10877 5 1 1 71647
0 10878 7 1 2 54232 71648
0 10879 5 1 1 10878
0 10880 7 1 2 10875 10879
0 10881 5 1 1 10880
0 10882 7 1 2 63011 10881
0 10883 5 1 1 10882
0 10884 7 2 2 55484 68708
0 10885 5 1 1 71650
0 10886 7 6 2 49878 57434
0 10887 7 1 2 47852 71652
0 10888 7 1 2 71651 10887
0 10889 5 1 1 10888
0 10890 7 1 2 10883 10889
0 10891 5 1 1 10890
0 10892 7 1 2 54938 10891
0 10893 5 1 1 10892
0 10894 7 1 2 53992 68735
0 10895 5 1 1 10894
0 10896 7 1 2 10893 10895
0 10897 5 1 1 10896
0 10898 7 1 2 56866 10897
0 10899 5 1 1 10898
0 10900 7 1 2 47853 3095
0 10901 5 1 1 10900
0 10902 7 1 2 64974 10901
0 10903 5 1 1 10902
0 10904 7 1 2 66073 10903
0 10905 5 1 1 10904
0 10906 7 1 2 10877 10905
0 10907 5 1 1 10906
0 10908 7 1 2 67632 10907
0 10909 5 1 1 10908
0 10910 7 1 2 10899 10909
0 10911 5 1 1 10910
0 10912 7 1 2 51717 10911
0 10913 5 1 1 10912
0 10914 7 1 2 10864 10913
0 10915 7 1 2 10862 10914
0 10916 7 3 2 69308 68363
0 10917 5 1 1 71658
0 10918 7 2 2 67178 68952
0 10919 5 1 1 71661
0 10920 7 1 2 10919 68336
0 10921 5 1 1 10920
0 10922 7 1 2 63012 10921
0 10923 5 1 1 10922
0 10924 7 1 2 10917 10923
0 10925 5 1 1 10924
0 10926 7 1 2 56867 10925
0 10927 5 1 1 10926
0 10928 7 3 2 54939 66411
0 10929 7 1 2 63326 71663
0 10930 5 1 1 10929
0 10931 7 1 2 68421 10930
0 10932 5 1 1 10931
0 10933 7 1 2 49879 10932
0 10934 5 1 1 10933
0 10935 7 1 2 10927 10934
0 10936 5 1 1 10935
0 10937 7 1 2 53993 10936
0 10938 5 1 1 10937
0 10939 7 3 2 64349 67967
0 10940 7 10 2 51523 67677
0 10941 7 1 2 71669 69929
0 10942 7 1 2 71666 10941
0 10943 5 1 1 10942
0 10944 7 1 2 10938 10943
0 10945 5 1 1 10944
0 10946 7 1 2 47854 10945
0 10947 5 1 1 10946
0 10948 7 2 2 64620 67518
0 10949 5 1 1 71679
0 10950 7 1 2 68642 71680
0 10951 5 1 1 10950
0 10952 7 2 2 62900 69720
0 10953 5 1 1 71681
0 10954 7 2 2 53994 64589
0 10955 5 1 1 71683
0 10956 7 1 2 63409 10955
0 10957 5 1 1 10956
0 10958 7 1 2 48714 10957
0 10959 5 1 1 10958
0 10960 7 1 2 66374 69604
0 10961 5 1 1 10960
0 10962 7 1 2 10959 10961
0 10963 5 1 1 10962
0 10964 7 1 2 67766 10963
0 10965 5 1 1 10964
0 10966 7 1 2 10953 10965
0 10967 5 1 1 10966
0 10968 7 1 2 57895 10967
0 10969 5 1 1 10968
0 10970 7 1 2 10951 10969
0 10971 7 1 2 10947 10970
0 10972 5 1 1 10971
0 10973 7 1 2 51718 10972
0 10974 5 1 1 10973
0 10975 7 1 2 69000 68516
0 10976 5 1 1 10975
0 10977 7 1 2 68486 10976
0 10978 5 1 1 10977
0 10979 7 1 2 65698 10978
0 10980 5 1 1 10979
0 10981 7 3 2 52776 66293
0 10982 5 1 1 71685
0 10983 7 1 2 66740 68521
0 10984 7 1 2 71686 10983
0 10985 5 1 1 10984
0 10986 7 1 2 10980 10985
0 10987 5 1 1 10986
0 10988 7 1 2 50674 10987
0 10989 5 1 1 10988
0 10990 7 2 2 66991 69058
0 10991 7 1 2 63327 71688
0 10992 5 1 1 10991
0 10993 7 1 2 68561 10992
0 10994 5 1 1 10993
0 10995 7 1 2 55622 10994
0 10996 5 1 1 10995
0 10997 7 1 2 68319 69658
0 10998 5 1 1 10997
0 10999 7 1 2 10996 10998
0 11000 5 1 1 10999
0 11001 7 1 2 67543 11000
0 11002 5 1 1 11001
0 11003 7 1 2 10989 11002
0 11004 7 1 2 10974 11003
0 11005 5 1 1 11004
0 11006 7 1 2 56059 11005
0 11007 5 1 1 11006
0 11008 7 4 2 52777 57435
0 11009 7 1 2 55623 67694
0 11010 7 1 2 71690 11009
0 11011 5 1 1 11010
0 11012 7 1 2 68325 11011
0 11013 5 1 1 11012
0 11014 7 1 2 61895 11013
0 11015 5 1 1 11014
0 11016 7 5 2 52778 54233
0 11017 7 3 2 56868 68456
0 11018 7 1 2 71694 71699
0 11019 5 1 1 11018
0 11020 7 1 2 11015 11019
0 11021 5 1 1 11020
0 11022 7 1 2 47855 11021
0 11023 5 1 1 11022
0 11024 7 1 2 64958 68320
0 11025 5 1 1 11024
0 11026 7 1 2 11023 11025
0 11027 5 1 1 11026
0 11028 7 1 2 54940 11027
0 11029 5 1 1 11028
0 11030 7 4 2 59349 68457
0 11031 7 1 2 63894 71702
0 11032 5 1 1 11031
0 11033 7 1 2 68326 11032
0 11034 5 1 1 11033
0 11035 7 1 2 65069 11034
0 11036 5 1 1 11035
0 11037 7 1 2 50972 59116
0 11038 5 1 1 11037
0 11039 7 1 2 59012 11038
0 11040 5 2 1 11039
0 11041 7 1 2 53995 68458
0 11042 7 1 2 71706 11041
0 11043 5 1 1 11042
0 11044 7 1 2 11036 11043
0 11045 7 1 2 11029 11044
0 11046 5 1 1 11045
0 11047 7 1 2 53665 11046
0 11048 5 1 1 11047
0 11049 7 4 2 55485 68800
0 11050 5 2 1 71708
0 11051 7 4 2 48715 57436
0 11052 7 2 2 49706 71714
0 11053 7 1 2 51524 64451
0 11054 7 1 2 71718 11053
0 11055 5 1 1 11054
0 11056 7 1 2 71712 11055
0 11057 5 1 1 11056
0 11058 7 1 2 56869 11057
0 11059 5 1 1 11058
0 11060 7 4 2 53459 67611
0 11061 5 1 1 71720
0 11062 7 1 2 68740 11061
0 11063 5 1 1 11062
0 11064 7 1 2 62712 11063
0 11065 5 1 1 11064
0 11066 7 1 2 55486 69682
0 11067 5 1 1 11066
0 11068 7 1 2 11065 11067
0 11069 5 1 1 11068
0 11070 7 1 2 49880 11069
0 11071 5 1 1 11070
0 11072 7 1 2 11059 11071
0 11073 5 1 1 11072
0 11074 7 1 2 54564 11073
0 11075 5 1 1 11074
0 11076 7 1 2 47856 68739
0 11077 5 2 1 11076
0 11078 7 1 2 53996 71721
0 11079 5 1 1 11078
0 11080 7 1 2 71724 11079
0 11081 5 1 1 11080
0 11082 7 1 2 71653 11081
0 11083 5 1 1 11082
0 11084 7 1 2 11075 11083
0 11085 5 1 1 11084
0 11086 7 1 2 51719 11085
0 11087 5 1 1 11086
0 11088 7 1 2 11048 11087
0 11089 5 1 1 11088
0 11090 7 1 2 55263 11089
0 11091 5 1 1 11090
0 11092 7 1 2 11007 11091
0 11093 7 1 2 10915 11092
0 11094 5 1 1 11093
0 11095 7 1 2 56699 11094
0 11096 5 1 1 11095
0 11097 7 1 2 67594 68690
0 11098 5 2 1 11097
0 11099 7 1 2 65974 66837
0 11100 5 1 1 11099
0 11101 7 1 2 71726 11100
0 11102 5 1 1 11101
0 11103 7 1 2 69023 11102
0 11104 5 1 1 11103
0 11105 7 2 2 63718 68459
0 11106 7 1 2 70344 71728
0 11107 5 1 1 11106
0 11108 7 1 2 11104 11107
0 11109 5 1 1 11108
0 11110 7 1 2 57145 11109
0 11111 5 1 1 11110
0 11112 7 5 2 49304 49881
0 11113 7 1 2 63283 71730
0 11114 7 2 2 70025 11113
0 11115 5 1 1 71735
0 11116 7 1 2 11111 11115
0 11117 5 1 1 11116
0 11118 7 1 2 58967 11117
0 11119 5 1 1 11118
0 11120 7 3 2 67922 68574
0 11121 7 3 2 62828 71737
0 11122 5 1 1 71740
0 11123 7 7 2 51525 68378
0 11124 5 1 1 71743
0 11125 7 3 2 69014 71744
0 11126 5 2 1 71750
0 11127 7 1 2 56870 71751
0 11128 5 1 1 11127
0 11129 7 1 2 11122 11128
0 11130 5 1 1 11129
0 11131 7 1 2 59102 11130
0 11132 5 1 1 11131
0 11133 7 20 2 53460 55487
0 11134 5 1 1 71755
0 11135 7 2 2 67899 71756
0 11136 5 3 1 71775
0 11137 7 1 2 56871 67767
0 11138 5 1 1 11137
0 11139 7 1 2 66438 11138
0 11140 5 3 1 11139
0 11141 7 1 2 63013 71780
0 11142 5 1 1 11141
0 11143 7 1 2 71777 11142
0 11144 5 2 1 11143
0 11145 7 6 2 47857 57437
0 11146 7 2 2 57146 71785
0 11147 5 3 1 71791
0 11148 7 1 2 50973 71793
0 11149 5 2 1 11148
0 11150 7 1 2 51720 71796
0 11151 7 1 2 71783 11150
0 11152 5 1 1 11151
0 11153 7 1 2 11132 11152
0 11154 5 1 1 11153
0 11155 7 1 2 54565 11154
0 11156 5 1 1 11155
0 11157 7 7 2 49305 63248
0 11158 7 3 2 49191 71798
0 11159 7 2 2 67633 71805
0 11160 7 1 2 71808 68970
0 11161 5 1 1 11160
0 11162 7 1 2 11156 11161
0 11163 7 1 2 11119 11162
0 11164 5 1 1 11163
0 11165 7 1 2 53997 11164
0 11166 5 1 1 11165
0 11167 7 3 2 65585 57849
0 11168 5 1 1 71810
0 11169 7 1 2 49707 71811
0 11170 5 1 1 11169
0 11171 7 1 2 53666 11170
0 11172 5 1 1 11171
0 11173 7 1 2 66074 11172
0 11174 5 1 1 11173
0 11175 7 1 2 66961 69099
0 11176 7 1 2 59103 11175
0 11177 5 1 1 11176
0 11178 7 1 2 11174 11177
0 11179 5 1 1 11178
0 11180 7 1 2 56872 11179
0 11181 5 1 1 11180
0 11182 7 1 2 67108 68822
0 11183 7 1 2 62453 11182
0 11184 5 1 1 11183
0 11185 7 1 2 11181 11184
0 11186 5 1 1 11185
0 11187 7 1 2 51721 11186
0 11188 5 1 1 11187
0 11189 7 1 2 11188 71753
0 11190 5 1 1 11189
0 11191 7 1 2 58108 11190
0 11192 5 1 1 11191
0 11193 7 1 2 53461 11168
0 11194 5 1 1 11193
0 11195 7 4 2 56873 70026
0 11196 7 1 2 69745 71813
0 11197 5 1 1 11196
0 11198 7 2 2 68658 68460
0 11199 7 1 2 53667 71817
0 11200 5 1 1 11199
0 11201 7 1 2 11197 11200
0 11202 5 1 1 11201
0 11203 7 1 2 11194 11202
0 11204 5 1 1 11203
0 11205 7 1 2 68190 71781
0 11206 5 1 1 11205
0 11207 7 1 2 71778 11206
0 11208 5 1 1 11207
0 11209 7 1 2 62454 69042
0 11210 7 1 2 11208 11209
0 11211 5 1 1 11210
0 11212 7 1 2 11204 11211
0 11213 7 1 2 11192 11212
0 11214 7 1 2 11166 11213
0 11215 5 1 1 11214
0 11216 7 1 2 54234 11215
0 11217 5 1 1 11216
0 11218 7 1 2 62421 71689
0 11219 5 1 1 11218
0 11220 7 1 2 68288 11219
0 11221 5 1 1 11220
0 11222 7 1 2 68546 11221
0 11223 5 1 1 11222
0 11224 7 1 2 68439 68285
0 11225 5 1 1 11224
0 11226 7 1 2 69746 11225
0 11227 5 1 1 11226
0 11228 7 7 2 53998 63450
0 11229 7 1 2 67768 71819
0 11230 5 1 1 11229
0 11231 7 1 2 68433 11230
0 11232 5 1 1 11231
0 11233 7 1 2 58109 11232
0 11234 5 1 1 11233
0 11235 7 1 2 11227 11234
0 11236 5 1 1 11235
0 11237 7 1 2 65699 11236
0 11238 5 1 1 11237
0 11239 7 1 2 62829 68628
0 11240 5 1 1 11239
0 11241 7 1 2 11238 11240
0 11242 5 1 1 11241
0 11243 7 1 2 51722 11242
0 11244 5 1 1 11243
0 11245 7 1 2 11223 11244
0 11246 5 1 1 11245
0 11247 7 1 2 59104 11246
0 11248 5 1 1 11247
0 11249 7 1 2 53999 69140
0 11250 7 1 2 69504 11249
0 11251 7 1 2 69735 11250
0 11252 5 1 1 11251
0 11253 7 1 2 11248 11252
0 11254 7 5 2 54566 66075
0 11255 5 5 1 71826
0 11256 7 1 2 66362 71831
0 11257 5 1 1 11256
0 11258 7 1 2 59253 11257
0 11259 5 1 1 11258
0 11260 7 1 2 5233 11259
0 11261 5 1 1 11260
0 11262 7 1 2 62543 11261
0 11263 5 1 1 11262
0 11264 7 2 2 67292 68691
0 11265 5 1 1 71836
0 11266 7 1 2 11265 10949
0 11267 5 1 1 11266
0 11268 7 1 2 59254 11267
0 11269 5 1 1 11268
0 11270 7 3 2 51526 62901
0 11271 7 7 2 49537 54000
0 11272 5 6 1 71841
0 11273 7 6 2 54567 71842
0 11274 7 1 2 48597 71854
0 11275 5 1 1 11274
0 11276 7 1 2 63847 11275
0 11277 5 1 1 11276
0 11278 7 1 2 71838 11277
0 11279 5 1 1 11278
0 11280 7 1 2 11269 11279
0 11281 7 1 2 11263 11280
0 11282 5 1 1 11281
0 11283 7 1 2 49882 11282
0 11284 5 1 1 11283
0 11285 7 1 2 71827 71809
0 11286 5 1 1 11285
0 11287 7 1 2 11284 11286
0 11288 5 1 1 11287
0 11289 7 1 2 51723 11288
0 11290 5 1 1 11289
0 11291 7 1 2 59255 71703
0 11292 5 1 1 11291
0 11293 7 1 2 54001 68321
0 11294 5 1 1 11293
0 11295 7 1 2 11292 11294
0 11296 5 1 1 11295
0 11297 7 1 2 53668 11296
0 11298 5 1 1 11297
0 11299 7 1 2 62422 68896
0 11300 5 1 1 11299
0 11301 7 1 2 11298 11300
0 11302 5 1 1 11301
0 11303 7 1 2 64590 11302
0 11304 5 1 1 11303
0 11305 7 2 2 63466 68857
0 11306 7 1 2 66849 71860
0 11307 7 1 2 69273 11306
0 11308 5 1 1 11307
0 11309 7 1 2 11304 11308
0 11310 5 1 1 11309
0 11311 7 1 2 56874 11310
0 11312 5 1 1 11311
0 11313 7 1 2 11290 11312
0 11314 7 1 2 11253 11313
0 11315 5 1 1 11314
0 11316 7 1 2 47858 11315
0 11317 5 1 1 11316
0 11318 7 2 2 59105 68461
0 11319 7 2 2 56875 68973
0 11320 7 1 2 71862 71864
0 11321 5 1 1 11320
0 11322 7 1 2 69115 11321
0 11323 5 1 1 11322
0 11324 7 1 2 58968 11323
0 11325 5 1 1 11324
0 11326 7 1 2 67923 71554
0 11327 5 1 1 11326
0 11328 7 1 2 11325 11327
0 11329 5 1 1 11328
0 11330 7 1 2 51252 11329
0 11331 5 1 1 11330
0 11332 7 5 2 54941 69520
0 11333 7 1 2 68946 71866
0 11334 5 1 1 11333
0 11335 7 1 2 63014 69024
0 11336 7 1 2 62455 11335
0 11337 5 1 1 11336
0 11338 7 1 2 11334 11337
0 11339 5 1 1 11338
0 11340 7 1 2 65975 11339
0 11341 5 1 1 11340
0 11342 7 1 2 11331 11341
0 11343 5 1 1 11342
0 11344 7 1 2 65853 11343
0 11345 5 1 1 11344
0 11346 7 1 2 59256 69043
0 11347 7 1 2 71784 11346
0 11348 5 1 1 11347
0 11349 7 1 2 11345 11348
0 11350 7 1 2 11317 11349
0 11351 7 1 2 11217 11350
0 11352 7 1 2 11096 11351
0 11353 5 1 1 11352
0 11354 7 1 2 68231 11353
0 11355 5 1 1 11354
0 11356 7 3 2 49429 67508
0 11357 7 1 2 71871 71752
0 11358 5 1 1 11357
0 11359 7 1 2 49008 70027
0 11360 5 1 1 11359
0 11361 7 1 2 11358 11360
0 11362 5 1 1 11361
0 11363 7 1 2 57438 11362
0 11364 5 1 1 11363
0 11365 7 13 2 51527 62544
0 11366 7 2 2 71874 69862
0 11367 5 1 1 71887
0 11368 7 4 2 48716 68801
0 11369 7 1 2 66412 71889
0 11370 5 1 1 11369
0 11371 7 1 2 11367 11370
0 11372 5 1 1 11371
0 11373 7 1 2 69044 11372
0 11374 5 1 1 11373
0 11375 7 1 2 11364 11374
0 11376 5 1 1 11375
0 11377 7 1 2 57896 11376
0 11378 5 1 1 11377
0 11379 7 4 2 55264 66760
0 11380 5 1 1 71893
0 11381 7 4 2 62545 57439
0 11382 7 2 2 51253 71897
0 11383 5 1 1 71901
0 11384 7 1 2 11380 11383
0 11385 5 1 1 11384
0 11386 7 1 2 55488 11385
0 11387 5 1 1 11386
0 11388 7 1 2 54942 69232
0 11389 5 1 1 11388
0 11390 7 1 2 11387 11389
0 11391 5 1 1 11390
0 11392 7 1 2 69081 11391
0 11393 5 1 1 11392
0 11394 7 1 2 11378 11393
0 11395 5 1 1 11394
0 11396 7 2 2 58266 61806
0 11397 5 2 1 71903
0 11398 7 2 2 54568 71905
0 11399 7 1 2 11395 71907
0 11400 5 1 1 11399
0 11401 7 1 2 65845 68512
0 11402 5 1 1 11401
0 11403 7 1 2 65586 61232
0 11404 5 1 1 11403
0 11405 7 1 2 11402 11404
0 11406 5 1 1 11405
0 11407 7 1 2 56700 11406
0 11408 5 1 1 11407
0 11409 7 2 2 54943 58969
0 11410 7 2 2 56876 62713
0 11411 5 1 1 71911
0 11412 7 1 2 71909 71912
0 11413 5 1 1 11412
0 11414 7 1 2 68507 11413
0 11415 5 1 1 11414
0 11416 7 1 2 57440 11415
0 11417 5 1 1 11416
0 11418 7 1 2 11408 11417
0 11419 5 1 1 11418
0 11420 7 1 2 69172 11419
0 11421 5 1 1 11420
0 11422 7 6 2 49009 53669
0 11423 5 1 1 71913
0 11424 7 1 2 57897 71890
0 11425 5 1 1 11424
0 11426 7 1 2 11423 11425
0 11427 5 1 1 11426
0 11428 7 5 2 55489 11427
0 11429 7 1 2 56993 70348
0 11430 5 1 1 11429
0 11431 7 2 2 56994 57843
0 11432 5 1 1 71924
0 11433 7 1 2 49192 11432
0 11434 7 1 2 11430 11433
0 11435 5 1 1 11434
0 11436 7 1 2 62714 67714
0 11437 5 1 1 11436
0 11438 7 1 2 65323 11437
0 11439 7 1 2 11435 11438
0 11440 5 1 1 11439
0 11441 7 1 2 71919 11440
0 11442 5 1 1 11441
0 11443 7 1 2 11421 11442
0 11444 5 1 1 11443
0 11445 7 1 2 55265 11444
0 11446 5 1 1 11445
0 11447 7 3 2 47859 67519
0 11448 7 1 2 63005 8013
0 11449 5 1 1 11448
0 11450 7 2 2 50974 6107
0 11451 5 5 1 71929
0 11452 7 1 2 66191 71931
0 11453 7 1 2 11449 11452
0 11454 5 1 1 11453
0 11455 7 1 2 67637 11454
0 11456 5 1 1 11455
0 11457 7 1 2 71926 11456
0 11458 5 1 1 11457
0 11459 7 2 2 60385 66076
0 11460 7 2 2 54944 66675
0 11461 7 1 2 71936 71938
0 11462 5 1 1 11461
0 11463 7 1 2 69251 11462
0 11464 5 1 1 11463
0 11465 7 1 2 56701 11464
0 11466 5 1 1 11465
0 11467 7 1 2 61269 66784
0 11468 5 1 1 11467
0 11469 7 1 2 58956 11468
0 11470 5 1 1 11469
0 11471 7 1 2 54002 68638
0 11472 5 1 1 11471
0 11473 7 1 2 69725 11472
0 11474 5 1 1 11473
0 11475 7 1 2 11470 11474
0 11476 5 1 1 11475
0 11477 7 1 2 11466 11476
0 11478 7 1 2 11458 11477
0 11479 5 1 1 11478
0 11480 7 1 2 49010 11479
0 11481 5 1 1 11480
0 11482 7 1 2 11446 11481
0 11483 5 1 1 11482
0 11484 7 1 2 54569 11483
0 11485 5 1 1 11484
0 11486 7 1 2 47860 65553
0 11487 5 1 1 11486
0 11488 7 1 2 64906 11487
0 11489 5 2 1 11488
0 11490 7 1 2 69453 71940
0 11491 5 1 1 11490
0 11492 7 1 2 67622 11491
0 11493 5 1 1 11492
0 11494 7 1 2 57441 11493
0 11495 5 1 1 11494
0 11496 7 1 2 11495 69279
0 11497 5 1 1 11496
0 11498 7 1 2 64215 11497
0 11499 5 1 1 11498
0 11500 7 3 2 55490 67551
0 11501 7 1 2 65058 71942
0 11502 5 1 1 11501
0 11503 7 1 2 71646 11502
0 11504 5 1 1 11503
0 11505 7 1 2 47861 11504
0 11506 5 1 1 11505
0 11507 7 1 2 64024 68623
0 11508 5 1 1 11507
0 11509 7 1 2 66112 11508
0 11510 5 1 1 11509
0 11511 7 1 2 63360 62191
0 11512 7 1 2 11510 11511
0 11513 5 1 1 11512
0 11514 7 1 2 11506 11513
0 11515 5 1 1 11514
0 11516 7 1 2 58970 11515
0 11517 5 1 1 11516
0 11518 7 1 2 57442 68425
0 11519 5 1 1 11518
0 11520 7 1 2 66679 68513
0 11521 5 1 1 11520
0 11522 7 1 2 11519 11521
0 11523 5 1 1 11522
0 11524 7 1 2 47862 11523
0 11525 5 1 1 11524
0 11526 7 1 2 11517 11525
0 11527 7 1 2 11499 11526
0 11528 5 1 1 11527
0 11529 7 1 2 49011 11528
0 11530 5 1 1 11529
0 11531 7 2 2 57898 71715
0 11532 7 1 2 64216 68802
0 11533 7 1 2 67109 11532
0 11534 7 1 2 71945 11533
0 11535 5 1 1 11534
0 11536 7 1 2 11530 11535
0 11537 7 1 2 11485 11536
0 11538 5 1 1 11537
0 11539 7 1 2 51724 11538
0 11540 5 1 1 11539
0 11541 7 1 2 11400 11540
0 11542 5 1 1 11541
0 11543 7 1 2 50009 11542
0 11544 5 1 1 11543
0 11545 7 1 2 49708 10842
0 11546 5 1 1 11545
0 11547 7 6 2 48347 61403
0 11548 5 2 1 71947
0 11549 7 2 2 62777 71948
0 11550 7 4 2 47863 66077
0 11551 5 1 1 71957
0 11552 7 1 2 64643 69025
0 11553 7 1 2 71958 11552
0 11554 7 1 2 71955 11553
0 11555 5 1 1 11554
0 11556 7 3 2 66294 66246
0 11557 5 1 1 71961
0 11558 7 1 2 68559 11557
0 11559 5 1 1 11558
0 11560 7 1 2 47864 11559
0 11561 5 1 1 11560
0 11562 7 2 2 59371 66295
0 11563 5 1 1 71964
0 11564 7 1 2 11561 11563
0 11565 5 1 1 11564
0 11566 7 1 2 68000 11565
0 11567 5 1 1 11566
0 11568 7 1 2 11567 8863
0 11569 5 1 1 11568
0 11570 7 1 2 56877 11569
0 11571 5 1 1 11570
0 11572 7 1 2 68575 69111
0 11573 5 1 1 11572
0 11574 7 1 2 11571 11573
0 11575 5 1 1 11574
0 11576 7 1 2 56060 11575
0 11577 5 1 1 11576
0 11578 7 1 2 11555 11577
0 11579 7 1 2 11546 11578
0 11580 5 1 1 11579
0 11581 7 1 2 68191 11580
0 11582 5 1 1 11581
0 11583 7 4 2 49306 50675
0 11584 7 2 2 68379 71966
0 11585 5 1 1 71970
0 11586 7 1 2 59612 71382
0 11587 5 1 1 11586
0 11588 7 1 2 69767 11587
0 11589 5 1 1 11588
0 11590 7 1 2 48348 11589
0 11591 5 1 1 11590
0 11592 7 1 2 11585 11591
0 11593 5 1 1 11592
0 11594 7 1 2 62715 11593
0 11595 5 1 1 11594
0 11596 7 1 2 64683 67096
0 11597 5 1 1 11596
0 11598 7 1 2 11595 11597
0 11599 5 1 1 11598
0 11600 7 1 2 68897 69401
0 11601 7 1 2 11599 11600
0 11602 5 1 1 11601
0 11603 7 1 2 11582 11602
0 11604 5 1 1 11603
0 11605 7 1 2 56702 11604
0 11606 5 1 1 11605
0 11607 7 2 2 66805 68380
0 11608 7 1 2 59106 71972
0 11609 5 1 1 11608
0 11610 7 3 2 54945 59257
0 11611 7 7 2 54235 68692
0 11612 7 1 2 71974 71977
0 11613 5 1 1 11612
0 11614 7 1 2 11609 11613
0 11615 5 1 1 11614
0 11616 7 2 2 68898 11615
0 11617 7 1 2 67511 71984
0 11618 5 1 1 11617
0 11619 7 1 2 63164 71985
0 11620 5 1 1 11619
0 11621 7 3 2 65910 71799
0 11622 5 2 1 71986
0 11623 7 1 2 64925 71989
0 11624 5 1 1 11623
0 11625 7 1 2 68916 11624
0 11626 5 1 1 11625
0 11627 7 1 2 5359 66924
0 11628 5 1 1 11627
0 11629 7 1 2 67561 11628
0 11630 5 1 1 11629
0 11631 7 1 2 11626 11630
0 11632 5 1 1 11631
0 11633 7 1 2 68858 11632
0 11634 5 1 1 11633
0 11635 7 1 2 61896 59107
0 11636 5 1 1 11635
0 11637 7 1 2 56995 11636
0 11638 5 1 1 11637
0 11639 7 1 2 54236 11638
0 11640 5 1 1 11639
0 11641 7 1 2 2490 63961
0 11642 5 1 1 11641
0 11643 7 1 2 47865 11642
0 11644 5 1 1 11643
0 11645 7 1 2 63467 11644
0 11646 7 1 2 11640 11645
0 11647 5 1 1 11646
0 11648 7 1 2 68899 11647
0 11649 5 1 1 11648
0 11650 7 1 2 11634 11649
0 11651 5 1 1 11650
0 11652 7 1 2 51254 11651
0 11653 5 1 1 11652
0 11654 7 1 2 64538 57768
0 11655 5 3 1 11654
0 11656 7 1 2 62445 67590
0 11657 5 1 1 11656
0 11658 7 1 2 71991 11657
0 11659 5 1 1 11658
0 11660 7 2 2 67179 68958
0 11661 7 1 2 56878 68340
0 11662 7 1 2 71994 11661
0 11663 7 1 2 11659 11662
0 11664 5 1 1 11663
0 11665 7 1 2 11653 11664
0 11666 5 1 1 11665
0 11667 7 1 2 62902 11666
0 11668 5 1 1 11667
0 11669 7 1 2 11620 11668
0 11670 5 1 1 11669
0 11671 7 1 2 57899 11670
0 11672 5 1 1 11671
0 11673 7 1 2 11618 11672
0 11674 7 1 2 11606 11673
0 11675 7 1 2 11544 11674
0 11676 5 1 1 11675
0 11677 7 1 2 68217 11676
0 11678 5 1 1 11677
0 11679 7 1 2 65088 63410
0 11680 5 1 1 11679
0 11681 7 1 2 62716 11680
0 11682 5 1 1 11681
0 11683 7 1 2 66381 11682
0 11684 5 1 1 11683
0 11685 7 1 2 55266 11684
0 11686 5 1 1 11685
0 11687 7 1 2 63403 67057
0 11688 5 1 1 11687
0 11689 7 1 2 11686 11688
0 11690 5 1 1 11689
0 11691 7 1 2 69952 11690
0 11692 5 1 1 11691
0 11693 7 4 2 49012 54946
0 11694 7 2 2 68959 71996
0 11695 5 1 1 72000
0 11696 7 1 2 54237 72001
0 11697 5 1 1 11696
0 11698 7 1 2 11692 11697
0 11699 5 1 1 11698
0 11700 7 1 2 67826 11699
0 11701 5 1 1 11700
0 11702 7 3 2 55267 68462
0 11703 7 1 2 72002 69869
0 11704 5 1 1 11703
0 11705 7 1 2 11701 11704
0 11706 5 1 1 11705
0 11707 7 1 2 48717 11706
0 11708 5 1 1 11707
0 11709 7 2 2 56879 69149
0 11710 7 2 2 69123 72005
0 11711 7 1 2 70048 71820
0 11712 7 1 2 72007 11711
0 11713 5 1 1 11712
0 11714 7 1 2 11708 11713
0 11715 5 1 1 11714
0 11716 7 1 2 57900 11715
0 11717 5 1 1 11716
0 11718 7 4 2 55268 55624
0 11719 7 3 2 67612 72009
0 11720 7 2 2 49883 72013
0 11721 7 1 2 47866 52861
0 11722 7 2 2 67512 11721
0 11723 7 1 2 61897 72018
0 11724 7 1 2 72016 11723
0 11725 5 1 1 11724
0 11726 7 1 2 53779 11725
0 11727 7 1 2 11717 11726
0 11728 5 1 1 11727
0 11729 7 1 2 64507 69082
0 11730 5 1 1 11729
0 11731 7 1 2 64613 69982
0 11732 5 1 1 11731
0 11733 7 1 2 11730 11732
0 11734 5 1 1 11733
0 11735 7 1 2 65070 11734
0 11736 5 1 1 11735
0 11737 7 2 2 51725 62546
0 11738 7 1 2 49013 57819
0 11739 7 1 2 72020 11738
0 11740 5 1 1 11739
0 11741 7 1 2 11736 11740
0 11742 5 1 1 11741
0 11743 7 1 2 54003 11742
0 11744 5 1 1 11743
0 11745 7 3 2 49014 54570
0 11746 7 1 2 72022 72021
0 11747 5 1 1 11746
0 11748 7 1 2 11744 11747
0 11749 5 1 1 11748
0 11750 7 1 2 51528 11749
0 11751 5 1 1 11750
0 11752 7 1 2 66506 68803
0 11753 7 1 2 69001 11752
0 11754 5 1 1 11753
0 11755 7 1 2 11751 11754
0 11756 5 1 1 11755
0 11757 7 1 2 57901 11756
0 11758 5 1 1 11757
0 11759 7 1 2 65505 65071
0 11760 5 1 1 11759
0 11761 7 1 2 69135 11760
0 11762 5 1 1 11761
0 11763 7 1 2 62717 11762
0 11764 5 1 1 11763
0 11765 7 1 2 54571 68497
0 11766 5 1 1 11765
0 11767 7 1 2 51529 11766
0 11768 7 1 2 11764 11767
0 11769 5 1 1 11768
0 11770 7 1 2 55491 6292
0 11771 7 1 2 6447 11770
0 11772 5 1 1 11771
0 11773 7 1 2 69083 11772
0 11774 7 1 2 11769 11773
0 11775 5 1 1 11774
0 11776 7 1 2 11758 11775
0 11777 5 1 1 11776
0 11778 7 1 2 55269 11777
0 11779 5 1 1 11778
0 11780 7 1 2 10885 7675
0 11781 5 1 1 11780
0 11782 7 1 2 58971 11781
0 11783 5 1 1 11782
0 11784 7 2 2 62830 69124
0 11785 5 1 1 72025
0 11786 7 2 2 54947 68514
0 11787 7 1 2 65544 72027
0 11788 5 1 1 11787
0 11789 7 1 2 11785 11788
0 11790 5 1 1 11789
0 11791 7 1 2 51530 11790
0 11792 5 1 1 11791
0 11793 7 1 2 11783 11792
0 11794 5 1 1 11793
0 11795 7 1 2 69084 11794
0 11796 5 1 1 11795
0 11797 7 1 2 50010 11796
0 11798 7 1 2 11779 11797
0 11799 5 1 1 11798
0 11800 7 1 2 57147 11799
0 11801 7 1 2 11728 11800
0 11802 5 1 1 11801
0 11803 7 4 2 49015 55625
0 11804 7 1 2 66449 72029
0 11805 5 1 1 11804
0 11806 7 2 2 65072 69953
0 11807 5 1 1 72033
0 11808 7 1 2 11807 8925
0 11809 5 1 1 11808
0 11810 7 3 2 47867 49884
0 11811 7 1 2 68613 72035
0 11812 7 1 2 11809 11811
0 11813 5 1 1 11812
0 11814 7 1 2 11805 11813
0 11815 5 1 1 11814
0 11816 7 1 2 55270 11815
0 11817 5 1 1 11816
0 11818 7 2 2 55492 68341
0 11819 7 1 2 52862 58507
0 11820 7 1 2 66529 69036
0 11821 7 1 2 11819 11820
0 11822 7 1 2 72038 11821
0 11823 5 1 1 11822
0 11824 7 1 2 11817 11823
0 11825 5 1 1 11824
0 11826 7 1 2 54948 11825
0 11827 5 1 1 11826
0 11828 7 2 2 67012 72010
0 11829 7 1 2 68342 70041
0 11830 7 1 2 72040 11829
0 11831 5 1 1 11830
0 11832 7 1 2 11827 11831
0 11833 5 1 1 11832
0 11834 7 1 2 48718 11833
0 11835 5 1 1 11834
0 11836 7 1 2 54949 72008
0 11837 7 1 2 70054 11836
0 11838 5 1 1 11837
0 11839 7 1 2 11835 11838
0 11840 5 1 1 11839
0 11841 7 1 2 57902 11840
0 11842 5 1 1 11841
0 11843 7 1 2 58673 72019
0 11844 7 1 2 72017 11843
0 11845 5 1 1 11844
0 11846 7 1 2 53780 11845
0 11847 7 1 2 11842 11846
0 11848 5 1 1 11847
0 11849 7 1 2 64606 6671
0 11850 5 3 1 11849
0 11851 7 1 2 64919 67695
0 11852 7 1 2 72042 11851
0 11853 5 1 1 11852
0 11854 7 1 2 66113 11853
0 11855 5 1 1 11854
0 11856 7 1 2 57903 11855
0 11857 5 1 1 11856
0 11858 7 1 2 65846 69234
0 11859 5 1 1 11858
0 11860 7 1 2 64556 67419
0 11861 5 1 1 11860
0 11862 7 1 2 69230 11861
0 11863 7 1 2 11859 11862
0 11864 7 1 2 11857 11863
0 11865 5 1 1 11864
0 11866 7 1 2 54950 11865
0 11867 5 1 1 11866
0 11868 7 1 2 69454 71684
0 11869 5 1 1 11868
0 11870 7 1 2 63885 69256
0 11871 5 1 1 11870
0 11872 7 1 2 11869 11871
0 11873 7 1 2 11867 11872
0 11874 5 1 1 11873
0 11875 7 1 2 69085 11874
0 11876 5 1 1 11875
0 11877 7 3 2 53670 56880
0 11878 7 2 2 72045 68761
0 11879 5 1 1 72048
0 11880 7 1 2 69787 72049
0 11881 5 1 1 11880
0 11882 7 1 2 71779 8982
0 11883 5 1 1 11882
0 11884 7 1 2 62718 69066
0 11885 7 1 2 11883 11884
0 11886 5 1 1 11885
0 11887 7 1 2 11881 11886
0 11888 5 1 1 11887
0 11889 7 1 2 48719 67313
0 11890 7 1 2 11888 11889
0 11891 5 1 1 11890
0 11892 7 1 2 50011 11891
0 11893 7 1 2 11876 11892
0 11894 5 1 1 11893
0 11895 7 1 2 56703 11894
0 11896 7 1 2 11848 11895
0 11897 5 1 1 11896
0 11898 7 1 2 11802 11897
0 11899 5 1 1 11898
0 11900 7 1 2 56061 11899
0 11901 5 1 1 11900
0 11902 7 1 2 67613 69192
0 11903 5 1 1 11902
0 11904 7 1 2 57443 69258
0 11905 5 1 1 11904
0 11906 7 1 2 11903 11905
0 11907 5 1 1 11906
0 11908 7 1 2 68947 11907
0 11909 5 1 1 11908
0 11910 7 7 2 51726 66413
0 11911 7 1 2 49885 71997
0 11912 7 1 2 72050 11911
0 11913 5 1 1 11912
0 11914 7 1 2 11909 11913
0 11915 5 1 1 11914
0 11916 7 1 2 71908 11915
0 11917 5 1 1 11916
0 11918 7 3 2 49016 68960
0 11919 5 1 1 72057
0 11920 7 10 2 55626 70042
0 11921 5 2 1 72060
0 11922 7 1 2 56881 72061
0 11923 5 1 1 11922
0 11924 7 1 2 11919 11923
0 11925 5 1 1 11924
0 11926 7 1 2 71932 11925
0 11927 5 1 1 11926
0 11928 7 1 2 64787 72062
0 11929 5 1 1 11928
0 11930 7 1 2 11927 11929
0 11931 5 1 1 11930
0 11932 7 1 2 48136 11931
0 11933 5 1 1 11932
0 11934 7 1 2 64805 69954
0 11935 5 1 1 11934
0 11936 7 1 2 7997 11935
0 11937 5 2 1 11936
0 11938 7 1 2 56882 72072
0 11939 5 1 1 11938
0 11940 7 1 2 57769 72063
0 11941 5 1 1 11940
0 11942 7 1 2 11939 11941
0 11943 5 1 1 11942
0 11944 7 1 2 55271 11943
0 11945 5 1 1 11944
0 11946 7 1 2 11933 11945
0 11947 5 1 1 11946
0 11948 7 1 2 62719 11947
0 11949 5 1 1 11948
0 11950 7 1 2 57444 72064
0 11951 5 1 1 11950
0 11952 7 1 2 61812 72073
0 11953 5 1 1 11952
0 11954 7 1 2 11951 11953
0 11955 5 1 1 11954
0 11956 7 1 2 55272 11955
0 11957 5 1 1 11956
0 11958 7 1 2 11949 11957
0 11959 5 1 1 11958
0 11960 7 1 2 54572 11959
0 11961 5 1 1 11960
0 11962 7 1 2 63905 66785
0 11963 5 1 1 11962
0 11964 7 1 2 69129 11963
0 11965 5 1 1 11964
0 11966 7 1 2 63825 69955
0 11967 7 1 2 11965 11966
0 11968 5 1 1 11967
0 11969 7 1 2 72065 71941
0 11970 5 1 1 11969
0 11971 7 1 2 11695 11970
0 11972 5 1 1 11971
0 11973 7 1 2 57445 64217
0 11974 7 1 2 11972 11973
0 11975 5 1 1 11974
0 11976 7 1 2 11968 11975
0 11977 7 1 2 11961 11976
0 11978 5 1 1 11977
0 11979 7 1 2 67827 11978
0 11980 5 1 1 11979
0 11981 7 1 2 11917 11980
0 11982 5 1 1 11981
0 11983 7 1 2 68192 11982
0 11984 5 1 1 11983
0 11985 7 2 2 54573 64417
0 11986 5 1 1 72074
0 11987 7 1 2 50676 65914
0 11988 5 3 1 11987
0 11989 7 1 2 48137 72076
0 11990 5 2 1 11989
0 11991 7 1 2 11986 72079
0 11992 5 2 1 11991
0 11993 7 1 2 58110 69150
0 11994 7 1 2 64647 61947
0 11995 7 1 2 70049 11994
0 11996 7 1 2 11993 11995
0 11997 7 1 2 72081 11996
0 11998 5 1 1 11997
0 11999 7 1 2 11984 11998
0 12000 5 1 1 11999
0 12001 7 1 2 53781 12000
0 12002 5 1 1 12001
0 12003 7 1 2 69261 69235
0 12004 5 1 1 12003
0 12005 7 3 2 69173 69166
0 12006 5 2 1 72083
0 12007 7 1 2 72086 8100
0 12008 5 2 1 12007
0 12009 7 1 2 48720 72088
0 12010 5 1 1 12009
0 12011 7 2 2 66962 68232
0 12012 7 1 2 51727 72090
0 12013 5 1 1 12012
0 12014 7 1 2 12010 12013
0 12015 5 1 1 12014
0 12016 7 1 2 56883 12015
0 12017 5 1 1 12016
0 12018 7 1 2 8394 71363
0 12019 5 4 1 12018
0 12020 7 1 2 48721 67900
0 12021 7 3 2 72092 12020
0 12022 7 1 2 67924 72096
0 12023 5 1 1 12022
0 12024 7 1 2 12017 12023
0 12025 5 1 1 12024
0 12026 7 1 2 57904 12025
0 12027 5 1 1 12026
0 12028 7 1 2 12004 12027
0 12029 5 1 1 12028
0 12030 7 1 2 54574 12029
0 12031 5 1 1 12030
0 12032 7 1 2 47868 69214
0 12033 5 1 1 12032
0 12034 7 1 2 12031 12033
0 12035 5 1 1 12034
0 12036 7 1 2 64143 12035
0 12037 5 1 1 12036
0 12038 7 1 2 67722 6724
0 12039 5 1 1 12038
0 12040 7 1 2 69200 12039
0 12041 5 1 1 12040
0 12042 7 1 2 68974 69444
0 12043 5 2 1 12042
0 12044 7 1 2 71364 72099
0 12045 5 2 1 12044
0 12046 7 1 2 72003 71667
0 12047 7 1 2 72101 12046
0 12048 5 1 1 12047
0 12049 7 1 2 8110 12048
0 12050 5 1 1 12049
0 12051 7 1 2 59577 12050
0 12052 5 1 1 12051
0 12053 7 7 2 49017 71331
0 12054 5 2 1 72103
0 12055 7 1 2 72093 68679
0 12056 5 1 1 12055
0 12057 7 1 2 72110 12056
0 12058 5 3 1 12057
0 12059 7 2 2 55493 72112
0 12060 7 1 2 65059 68961
0 12061 7 1 2 72115 12060
0 12062 5 1 1 12061
0 12063 7 1 2 12052 12062
0 12064 7 1 2 12041 12063
0 12065 5 1 1 12064
0 12066 7 1 2 57446 12065
0 12067 5 1 1 12066
0 12068 7 1 2 12037 12067
0 12069 5 1 1 12068
0 12070 7 1 2 61547 12069
0 12071 5 1 1 12070
0 12072 7 1 2 12002 12071
0 12073 7 1 2 11901 12072
0 12074 7 1 2 11678 12073
0 12075 5 1 1 12074
0 12076 7 1 2 48904 12075
0 12077 5 1 1 12076
0 12078 7 1 2 11355 12077
0 12079 5 1 1 12078
0 12080 7 1 2 55738 12079
0 12081 5 1 1 12080
0 12082 7 1 2 67958 8757
0 12083 5 2 1 12082
0 12084 7 2 2 69595 72117
0 12085 7 2 2 69863 72119
0 12086 5 1 1 72121
0 12087 7 2 2 53886 51255
0 12088 7 1 2 65330 72123
0 12089 7 1 2 64882 12088
0 12090 5 2 1 12089
0 12091 7 1 2 8852 72125
0 12092 5 1 1 12091
0 12093 7 1 2 69702 12092
0 12094 5 1 1 12093
0 12095 7 2 2 58382 68576
0 12096 5 1 1 72127
0 12097 7 1 2 58111 72128
0 12098 7 1 2 65652 12097
0 12099 5 1 1 12098
0 12100 7 1 2 12094 12099
0 12101 5 1 1 12100
0 12102 7 1 2 49886 12101
0 12103 5 1 1 12102
0 12104 7 1 2 66482 72126
0 12105 5 1 1 12104
0 12106 7 1 2 49018 63025
0 12107 7 1 2 12105 12106
0 12108 5 1 1 12107
0 12109 7 1 2 12103 12108
0 12110 5 1 1 12109
0 12111 7 1 2 55494 12110
0 12112 5 1 1 12111
0 12113 7 1 2 12086 12112
0 12114 5 1 1 12113
0 12115 7 1 2 50012 12114
0 12116 5 1 1 12115
0 12117 7 3 2 51256 67992
0 12118 7 1 2 65438 68148
0 12119 7 1 2 72129 12118
0 12120 5 1 1 12119
0 12121 7 1 2 8420 12120
0 12122 5 1 1 12121
0 12123 7 8 2 48905 55495
0 12124 7 1 2 71634 72132
0 12125 7 1 2 12122 12124
0 12126 5 1 1 12125
0 12127 7 1 2 51728 12126
0 12128 7 1 2 12116 12127
0 12129 5 1 1 12128
0 12130 7 5 2 52779 71332
0 12131 5 2 1 72140
0 12132 7 4 2 53887 65976
0 12133 7 2 2 49019 49111
0 12134 7 1 2 57447 72151
0 12135 7 1 2 72147 12134
0 12136 7 1 2 72141 12135
0 12137 5 1 1 12136
0 12138 7 1 2 64571 69186
0 12139 7 1 2 67284 12138
0 12140 7 1 2 72006 12139
0 12141 5 1 1 12140
0 12142 7 1 2 55627 12141
0 12143 7 1 2 12137 12142
0 12144 5 1 1 12143
0 12145 7 1 2 54951 12144
0 12146 7 1 2 12129 12145
0 12147 5 1 1 12146
0 12148 7 2 2 69986 72118
0 12149 7 3 2 53888 55273
0 12150 7 2 2 49112 72155
0 12151 5 1 1 72158
0 12152 7 1 2 49020 72159
0 12153 7 1 2 72153 12152
0 12154 5 1 1 12153
0 12155 7 2 2 57448 69788
0 12156 5 2 1 72160
0 12157 7 1 2 72162 12096
0 12158 5 1 1 12157
0 12159 7 1 2 69703 12158
0 12160 5 1 1 12159
0 12161 7 2 2 49021 68415
0 12162 7 1 2 58383 72164
0 12163 5 1 1 12162
0 12164 7 1 2 12160 12163
0 12165 5 1 1 12164
0 12166 7 1 2 68975 68948
0 12167 7 1 2 12165 12166
0 12168 5 1 1 12167
0 12169 7 1 2 12154 12168
0 12170 5 1 1 12169
0 12171 7 1 2 50013 12170
0 12172 5 1 1 12171
0 12173 7 1 2 57449 69460
0 12174 5 2 1 12173
0 12175 7 6 2 51257 62677
0 12176 7 3 2 49113 69759
0 12177 7 1 2 72168 72174
0 12178 5 1 1 12177
0 12179 7 1 2 72166 12178
0 12180 5 1 1 12179
0 12181 7 2 2 56884 69693
0 12182 7 1 2 72030 72177
0 12183 7 1 2 12180 12182
0 12184 5 1 1 12183
0 12185 7 1 2 12172 12184
0 12186 5 1 1 12185
0 12187 7 1 2 51531 12186
0 12188 5 1 1 12187
0 12189 7 4 2 48906 52863
0 12190 7 1 2 66555 72179
0 12191 7 1 2 63057 12190
0 12192 7 4 2 49709 69939
0 12193 5 1 1 72183
0 12194 7 2 2 55628 72156
0 12195 7 1 2 72184 72187
0 12196 7 1 2 12191 12195
0 12197 5 1 1 12196
0 12198 7 1 2 12188 12197
0 12199 7 1 2 12147 12198
0 12200 5 1 1 12199
0 12201 7 1 2 56704 12200
0 12202 5 1 1 12201
0 12203 7 4 2 52780 51532
0 12204 5 2 1 72189
0 12205 7 3 2 55629 72190
0 12206 7 2 2 71914 72195
0 12207 7 1 2 69476 72198
0 12208 5 2 1 12207
0 12209 7 4 2 50014 69557
0 12210 5 1 1 72202
0 12211 7 4 2 49022 72203
0 12212 5 2 1 72206
0 12213 7 1 2 68276 69645
0 12214 5 2 1 12213
0 12215 7 3 2 68218 72212
0 12216 7 1 2 63015 72214
0 12217 5 1 1 12216
0 12218 7 1 2 72210 12217
0 12219 5 1 1 12218
0 12220 7 1 2 71814 12219
0 12221 5 1 1 12220
0 12222 7 1 2 72200 12221
0 12223 5 1 1 12222
0 12224 7 1 2 71975 12223
0 12225 5 1 1 12224
0 12226 7 1 2 62903 72215
0 12227 5 1 1 12226
0 12228 7 1 2 12227 72211
0 12229 5 9 1 12228
0 12230 7 2 2 57905 72217
0 12231 5 1 1 72226
0 12232 7 3 2 62547 68233
0 12233 5 1 1 72228
0 12234 7 1 2 69558 72229
0 12235 5 1 1 12234
0 12236 7 1 2 12231 12235
0 12237 5 1 1 12236
0 12238 7 1 2 70028 71800
0 12239 7 1 2 12237 12238
0 12240 5 1 1 12239
0 12241 7 1 2 12225 12240
0 12242 7 1 2 12202 12241
0 12243 5 1 1 12242
0 12244 7 1 2 54238 12243
0 12245 5 1 1 12244
0 12246 7 1 2 64806 66963
0 12247 5 3 1 12246
0 12248 7 1 2 11134 72231
0 12249 5 1 1 12248
0 12250 7 1 2 69704 12249
0 12251 5 1 1 12250
0 12252 7 1 2 57450 71998
0 12253 7 1 2 66992 12252
0 12254 5 1 1 12253
0 12255 7 1 2 12251 12254
0 12256 5 1 1 12255
0 12257 7 1 2 49887 12256
0 12258 5 1 1 12257
0 12259 7 1 2 63086 67598
0 12260 5 1 1 12259
0 12261 7 1 2 64838 67180
0 12262 5 1 1 12261
0 12263 7 1 2 66559 12262
0 12264 5 1 1 12263
0 12265 7 1 2 62548 12264
0 12266 5 1 1 12265
0 12267 7 1 2 12260 12266
0 12268 5 1 1 12267
0 12269 7 1 2 49023 12268
0 12270 5 1 1 12269
0 12271 7 1 2 12258 12270
0 12272 5 1 1 12271
0 12273 7 1 2 65700 12272
0 12274 5 1 1 12273
0 12275 7 2 2 57906 70061
0 12276 5 1 1 72234
0 12277 7 1 2 49888 64373
0 12278 5 1 1 12277
0 12279 7 1 2 12276 12278
0 12280 5 1 1 12279
0 12281 7 1 2 69174 12280
0 12282 5 1 1 12281
0 12283 7 1 2 12274 12282
0 12284 5 1 1 12283
0 12285 7 1 2 50015 12284
0 12286 5 1 1 12285
0 12287 7 1 2 8096 72232
0 12288 5 1 1 12287
0 12289 7 7 2 48722 49889
0 12290 7 1 2 72236 71434
0 12291 7 1 2 65654 12290
0 12292 7 1 2 12288 12291
0 12293 5 1 1 12292
0 12294 7 1 2 12286 12293
0 12295 5 1 1 12294
0 12296 7 1 2 51729 12295
0 12297 5 1 1 12296
0 12298 7 2 2 52781 50016
0 12299 7 2 2 71915 72243
0 12300 7 1 2 66710 72245
0 12301 5 1 1 12300
0 12302 7 3 2 68207 69612
0 12303 7 1 2 64807 65701
0 12304 7 1 2 72247 12303
0 12305 7 1 2 63016 12304
0 12306 5 1 1 12305
0 12307 7 1 2 12301 12306
0 12308 5 1 1 12307
0 12309 7 1 2 69141 12308
0 12310 5 1 1 12309
0 12311 7 1 2 12297 12310
0 12312 5 1 1 12311
0 12313 7 1 2 61970 12312
0 12314 5 1 1 12313
0 12315 7 2 2 69477 69994
0 12316 5 2 1 72250
0 12317 7 1 2 53782 67166
0 12318 5 1 1 12317
0 12319 7 2 2 68522 12318
0 12320 7 1 2 72254 71865
0 12321 5 1 1 12320
0 12322 7 1 2 72252 12321
0 12323 5 1 1 12322
0 12324 7 1 2 57907 12323
0 12325 5 1 1 12324
0 12326 7 1 2 72046 70095
0 12327 5 1 1 12326
0 12328 7 1 2 68962 70062
0 12329 5 1 1 12328
0 12330 7 1 2 12327 12329
0 12331 5 1 1 12330
0 12332 7 1 2 50017 12331
0 12333 5 1 1 12332
0 12334 7 1 2 12325 12333
0 12335 5 1 1 12334
0 12336 7 1 2 49024 12335
0 12337 5 1 1 12336
0 12338 7 2 2 49710 71333
0 12339 5 2 1 72256
0 12340 7 1 2 69365 72257
0 12341 7 1 2 72178 12340
0 12342 5 1 1 12341
0 12343 7 1 2 12337 12342
0 12344 5 1 1 12343
0 12345 7 1 2 51533 12344
0 12346 5 1 1 12345
0 12347 7 2 2 53783 68680
0 12348 5 1 1 72260
0 12349 7 2 2 49711 72180
0 12350 7 1 2 70050 72262
0 12351 7 1 2 72261 12350
0 12352 5 1 1 12351
0 12353 7 1 2 12346 12352
0 12354 5 1 1 12353
0 12355 7 1 2 57451 12354
0 12356 5 1 1 12355
0 12357 7 1 2 64901 72104
0 12358 7 1 2 71818 12357
0 12359 5 1 1 12358
0 12360 7 1 2 12356 12359
0 12361 7 1 2 12314 12360
0 12362 7 1 2 12245 12361
0 12363 5 1 1 12362
0 12364 7 1 2 54575 12363
0 12365 5 1 1 12364
0 12366 7 1 2 64907 12151
0 12367 5 1 1 12366
0 12368 7 1 2 57148 12367
0 12369 5 1 1 12368
0 12370 7 1 2 65522 12369
0 12371 5 1 1 12370
0 12372 7 4 2 72084 70063
0 12373 5 3 1 72264
0 12374 7 1 2 48907 72089
0 12375 5 1 1 12374
0 12376 7 2 2 67769 69262
0 12377 5 2 1 72271
0 12378 7 1 2 12375 72273
0 12379 5 1 1 12378
0 12380 7 1 2 48723 12379
0 12381 5 1 1 12380
0 12382 7 1 2 69987 72091
0 12383 5 1 1 12382
0 12384 7 1 2 12381 12383
0 12385 5 10 1 12384
0 12386 7 1 2 57908 72275
0 12387 5 1 1 12386
0 12388 7 1 2 72268 12387
0 12389 5 1 1 12388
0 12390 7 1 2 12371 12389
0 12391 5 1 1 12390
0 12392 7 1 2 12233 10400
0 12393 5 1 1 12392
0 12394 7 11 2 55630 69906
0 12395 7 3 2 68976 72285
0 12396 7 1 2 67375 72296
0 12397 7 1 2 12393 12396
0 12398 5 1 1 12397
0 12399 7 1 2 71344 12348
0 12400 5 1 1 12399
0 12401 7 1 2 48908 12400
0 12402 5 1 1 12401
0 12403 7 1 2 50018 68780
0 12404 5 1 1 12403
0 12405 7 1 2 12402 12404
0 12406 5 1 1 12405
0 12407 7 1 2 49025 12406
0 12408 5 1 1 12407
0 12409 7 6 2 49890 50019
0 12410 5 1 1 72299
0 12411 7 6 2 65624 72300
0 12412 7 18 2 49538 53462
0 12413 5 2 1 72311
0 12414 7 3 2 48598 72312
0 12415 5 2 1 72331
0 12416 7 1 2 72305 72332
0 12417 5 1 1 12416
0 12418 7 1 2 12408 12417
0 12419 5 1 1 12418
0 12420 7 1 2 68131 69300
0 12421 7 1 2 12419 12420
0 12422 5 1 1 12421
0 12423 7 1 2 12398 12422
0 12424 7 1 2 12391 12423
0 12425 5 1 1 12424
0 12426 7 1 2 57452 12425
0 12427 5 1 1 12426
0 12428 7 5 2 56885 66078
0 12429 5 1 1 72336
0 12430 7 2 2 69559 72337
0 12431 5 1 1 72341
0 12432 7 1 2 51730 72342
0 12433 5 1 1 12432
0 12434 7 1 2 71754 12433
0 12435 5 1 1 12434
0 12436 7 1 2 58112 12435
0 12437 5 1 1 12436
0 12438 7 1 2 53671 62837
0 12439 5 1 1 12438
0 12440 7 1 2 56886 71738
0 12441 7 1 2 12439 12440
0 12442 5 1 1 12441
0 12443 7 1 2 12437 12442
0 12444 5 1 1 12443
0 12445 7 1 2 50020 12444
0 12446 5 1 1 12445
0 12447 7 4 2 64288 69613
0 12448 7 1 2 62904 70029
0 12449 7 1 2 72343 12448
0 12450 5 1 1 12449
0 12451 7 1 2 12446 12450
0 12452 5 1 1 12451
0 12453 7 1 2 49026 12452
0 12454 5 1 1 12453
0 12455 7 1 2 64289 71739
0 12456 7 1 2 72306 12455
0 12457 5 1 1 12456
0 12458 7 1 2 12454 12457
0 12459 5 1 1 12458
0 12460 7 1 2 54239 12459
0 12461 5 1 1 12460
0 12462 7 1 2 12427 12461
0 12463 7 1 2 12365 12462
0 12464 5 1 1 12463
0 12465 7 1 2 59983 12464
0 12466 5 1 1 12465
0 12467 7 3 2 65572 67325
0 12468 7 1 2 69709 72347
0 12469 5 1 1 12468
0 12470 7 1 2 64662 66972
0 12471 5 1 1 12470
0 12472 7 1 2 57990 12471
0 12473 5 1 1 12472
0 12474 7 1 2 58253 69596
0 12475 7 1 2 12473 12474
0 12476 5 1 1 12475
0 12477 7 1 2 12469 12476
0 12478 5 1 1 12477
0 12479 7 1 2 55274 12478
0 12480 5 1 1 12479
0 12481 7 6 2 48909 67770
0 12482 5 7 1 72350
0 12483 7 3 2 57276 61607
0 12484 7 1 2 67013 69584
0 12485 7 1 2 72363 12484
0 12486 5 1 1 12485
0 12487 7 1 2 72356 12486
0 12488 7 1 2 12480 12487
0 12489 5 1 1 12488
0 12490 7 1 2 50021 12489
0 12491 5 1 1 12490
0 12492 7 1 2 68330 72344
0 12493 5 1 1 12492
0 12494 7 1 2 12491 12493
0 12495 5 1 1 12494
0 12496 7 1 2 57453 12495
0 12497 5 1 1 12496
0 12498 7 1 2 56887 69597
0 12499 5 1 1 12498
0 12500 7 1 2 66439 12499
0 12501 5 1 1 12500
0 12502 7 2 2 54952 64171
0 12503 7 4 2 47869 48599
0 12504 7 2 2 50022 54576
0 12505 7 1 2 72368 72372
0 12506 7 1 2 72366 12505
0 12507 7 1 2 12501 12506
0 12508 5 1 1 12507
0 12509 7 1 2 12497 12508
0 12510 5 1 1 12509
0 12511 7 1 2 51731 12510
0 12512 5 1 1 12511
0 12513 7 3 2 61107 61478
0 12514 5 1 1 72374
0 12515 7 1 2 56996 12514
0 12516 5 1 1 12515
0 12517 7 1 2 71334 68917
0 12518 7 1 2 72286 12517
0 12519 7 1 2 12516 12518
0 12520 5 1 1 12519
0 12521 7 1 2 12512 12520
0 12522 5 1 1 12521
0 12523 7 1 2 49027 12522
0 12524 5 1 1 12523
0 12525 7 1 2 59128 69167
0 12526 5 4 1 12525
0 12527 7 1 2 57149 68653
0 12528 7 1 2 69971 12527
0 12529 5 1 1 12528
0 12530 7 1 2 72377 12529
0 12531 5 1 1 12530
0 12532 7 2 2 66414 72345
0 12533 7 1 2 57454 72381
0 12534 7 1 2 12531 12533
0 12535 5 1 1 12534
0 12536 7 1 2 12524 12535
0 12537 5 1 1 12536
0 12538 7 1 2 62549 12537
0 12539 5 1 1 12538
0 12540 7 3 2 49307 53463
0 12541 7 5 2 48349 72383
0 12542 7 1 2 66465 69977
0 12543 7 1 2 72386 12542
0 12544 5 2 1 12543
0 12545 7 1 2 69614 69045
0 12546 5 1 1 12545
0 12547 7 1 2 72391 12546
0 12548 5 1 1 12547
0 12549 7 1 2 66450 12548
0 12550 5 1 1 12549
0 12551 7 1 2 64318 69585
0 12552 5 1 1 12551
0 12553 7 1 2 63826 71180
0 12554 5 1 1 12553
0 12555 7 1 2 12552 12554
0 12556 5 1 1 12555
0 12557 7 1 2 67925 12556
0 12558 5 1 1 12557
0 12559 7 1 2 12550 12558
0 12560 5 1 1 12559
0 12561 7 1 2 54577 12560
0 12562 5 1 1 12561
0 12563 7 3 2 68717 68523
0 12564 5 2 1 72393
0 12565 7 1 2 65702 69988
0 12566 5 1 1 12565
0 12567 7 1 2 72396 12566
0 12568 5 2 1 12567
0 12569 7 2 2 51534 71976
0 12570 7 1 2 57909 72400
0 12571 7 1 2 72398 12570
0 12572 5 1 1 12571
0 12573 7 1 2 12562 12572
0 12574 5 1 1 12573
0 12575 7 1 2 47870 12574
0 12576 5 1 1 12575
0 12577 7 2 2 48350 67771
0 12578 5 1 1 72402
0 12579 7 1 2 51732 64439
0 12580 7 1 2 67038 12579
0 12581 7 1 2 72403 12580
0 12582 5 1 1 12581
0 12583 7 1 2 12576 12582
0 12584 5 1 1 12583
0 12585 7 1 2 54240 12584
0 12586 5 1 1 12585
0 12587 7 10 2 52782 55496
0 12588 7 1 2 66272 72404
0 12589 5 1 1 12588
0 12590 7 1 2 59397 67420
0 12591 7 1 2 66192 12590
0 12592 5 1 1 12591
0 12593 7 1 2 12589 12592
0 12594 5 1 1 12593
0 12595 7 1 2 68547 12594
0 12596 5 1 1 12595
0 12597 7 3 2 55497 69989
0 12598 5 2 1 72414
0 12599 7 1 2 72415 68727
0 12600 5 1 1 12599
0 12601 7 1 2 12596 12600
0 12602 5 1 1 12601
0 12603 7 1 2 50975 12602
0 12604 5 1 1 12603
0 12605 7 4 2 57150 71828
0 12606 5 1 1 72419
0 12607 7 1 2 69560 72420
0 12608 5 1 1 12607
0 12609 7 1 2 72357 12608
0 12610 5 1 1 12609
0 12611 7 1 2 69049 12610
0 12612 5 1 1 12611
0 12613 7 1 2 12604 12612
0 12614 5 1 1 12613
0 12615 7 1 2 57455 12614
0 12616 5 1 1 12615
0 12617 7 1 2 64644 66688
0 12618 7 1 2 67065 12617
0 12619 7 1 2 72287 12618
0 12620 5 1 1 12619
0 12621 7 1 2 12616 12620
0 12622 7 1 2 12586 12621
0 12623 5 1 1 12622
0 12624 7 1 2 68234 12623
0 12625 5 1 1 12624
0 12626 7 1 2 12539 12625
0 12627 7 1 2 56888 68001
0 12628 5 1 1 12627
0 12629 7 1 2 72397 12628
0 12630 5 1 1 12629
0 12631 7 1 2 72375 12630
0 12632 5 1 1 12631
0 12633 7 1 2 56889 72394
0 12634 5 1 1 12633
0 12635 7 1 2 12632 12634
0 12636 5 1 1 12635
0 12637 7 1 2 67181 12636
0 12638 5 1 1 12637
0 12639 7 1 2 71736 72364
0 12640 5 1 1 12639
0 12641 7 1 2 12638 12640
0 12642 5 1 1 12641
0 12643 7 1 2 57910 12642
0 12644 5 1 1 12643
0 12645 7 3 2 55275 59129
0 12646 7 2 2 67926 72423
0 12647 7 1 2 71642 72426
0 12648 5 1 1 12647
0 12649 7 1 2 12644 12648
0 12650 5 1 1 12649
0 12651 7 1 2 68219 12650
0 12652 5 1 1 12651
0 12653 7 1 2 52864 57911
0 12654 7 1 2 69940 69142
0 12655 7 1 2 12653 12654
0 12656 5 1 1 12655
0 12657 7 1 2 72087 12656
0 12658 5 3 1 12657
0 12659 7 1 2 48138 64757
0 12660 5 1 1 12659
0 12661 7 1 2 5217 12660
0 12662 5 1 1 12661
0 12663 7 1 2 72428 12662
0 12664 5 1 1 12663
0 12665 7 2 2 61413 59258
0 12666 7 1 2 72014 69450
0 12667 7 1 2 72431 12666
0 12668 5 1 1 12667
0 12669 7 1 2 12664 12668
0 12670 5 1 1 12669
0 12671 7 1 2 54241 12670
0 12672 5 1 1 12671
0 12673 7 1 2 50023 64319
0 12674 7 1 2 69121 12673
0 12675 5 1 1 12674
0 12676 7 1 2 12672 12675
0 12677 7 1 2 12652 12676
0 12678 5 1 1 12677
0 12679 7 1 2 48910 12678
0 12680 5 1 1 12679
0 12681 7 1 2 58254 67772
0 12682 5 1 1 12681
0 12683 7 1 2 55498 66693
0 12684 5 1 1 12683
0 12685 7 1 2 12682 12684
0 12686 5 1 1 12685
0 12687 7 1 2 55276 12686
0 12688 5 1 1 12687
0 12689 7 1 2 64645 65977
0 12690 7 1 2 67372 12689
0 12691 5 1 1 12690
0 12692 7 1 2 71832 12691
0 12693 5 1 1 12692
0 12694 7 1 2 57820 12693
0 12695 5 1 1 12694
0 12696 7 1 2 67798 12606
0 12697 7 1 2 12695 12696
0 12698 5 1 1 12697
0 12699 7 1 2 57912 12698
0 12700 5 1 1 12699
0 12701 7 1 2 12688 12700
0 12702 5 1 1 12701
0 12703 7 1 2 57456 12702
0 12704 5 1 1 12703
0 12705 7 1 2 64144 57735
0 12706 7 1 2 71782 12705
0 12707 5 1 1 12706
0 12708 7 1 2 12704 12707
0 12709 5 1 1 12708
0 12710 7 1 2 69263 12709
0 12711 5 1 1 12710
0 12712 7 1 2 12680 12711
0 12713 5 1 1 12712
0 12714 7 1 2 49712 12713
0 12715 5 1 1 12714
0 12716 7 2 2 55499 72036
0 12717 7 3 2 54242 69046
0 12718 7 1 2 72094 72435
0 12719 7 1 2 72433 12718
0 12720 5 1 1 12719
0 12721 7 1 2 57457 71700
0 12722 7 1 2 72102 12721
0 12723 7 1 2 72365 12722
0 12724 5 1 1 12723
0 12725 7 1 2 12720 12724
0 12726 5 1 1 12725
0 12727 7 1 2 64591 67262
0 12728 7 1 2 12726 12727
0 12729 5 1 1 12728
0 12730 7 1 2 12715 12729
0 12731 5 1 1 12730
0 12732 7 1 2 48724 12731
0 12733 5 1 1 12732
0 12734 7 1 2 64886 69274
0 12735 5 1 1 12734
0 12736 7 1 2 61425 69789
0 12737 5 1 1 12736
0 12738 7 1 2 12735 12737
0 12739 5 1 1 12738
0 12740 7 1 2 50976 12739
0 12741 5 1 1 12740
0 12742 7 1 2 68659 69131
0 12743 5 1 1 12742
0 12744 7 1 2 12741 12743
0 12745 5 1 1 12744
0 12746 7 1 2 68548 12745
0 12747 5 1 1 12746
0 12748 7 1 2 71939 72154
0 12749 5 1 1 12748
0 12750 7 1 2 12747 12749
0 12751 5 1 1 12750
0 12752 7 1 2 51535 12751
0 12753 5 1 1 12752
0 12754 7 8 2 49539 51258
0 12755 7 4 2 48600 72438
0 12756 5 2 1 72446
0 12757 7 1 2 64145 72447
0 12758 5 2 1 12757
0 12759 7 2 2 56890 66797
0 12760 5 3 1 72454
0 12761 7 1 2 57458 71894
0 12762 5 1 1 12761
0 12763 7 1 2 72456 12762
0 12764 5 1 1 12763
0 12765 7 1 2 47871 12764
0 12766 5 1 1 12765
0 12767 7 1 2 72452 12766
0 12768 5 1 1 12767
0 12769 7 1 2 63087 12768
0 12770 5 1 1 12769
0 12771 7 1 2 54953 72161
0 12772 5 1 1 12771
0 12773 7 1 2 72457 12772
0 12774 5 1 1 12773
0 12775 7 1 2 47872 12774
0 12776 5 1 1 12775
0 12777 7 1 2 12776 72453
0 12778 5 1 1 12777
0 12779 7 1 2 49891 12778
0 12780 5 1 1 12779
0 12781 7 1 2 65513 69586
0 12782 5 1 1 12781
0 12783 7 2 2 57459 72369
0 12784 7 2 2 64196 66466
0 12785 5 1 1 72461
0 12786 7 1 2 72459 72462
0 12787 5 1 1 12786
0 12788 7 1 2 12782 12787
0 12789 5 1 1 12788
0 12790 7 1 2 62550 12789
0 12791 5 1 1 12790
0 12792 7 1 2 12780 12791
0 12793 7 1 2 12770 12792
0 12794 5 1 1 12793
0 12795 7 1 2 67927 12794
0 12796 5 1 1 12795
0 12797 7 1 2 12753 12796
0 12798 5 1 1 12797
0 12799 7 1 2 50024 12798
0 12800 5 1 1 12799
0 12801 7 1 2 64808 69461
0 12802 5 1 1 12801
0 12803 7 1 2 68786 12802
0 12804 5 1 1 12803
0 12805 7 1 2 47873 12804
0 12806 5 1 1 12805
0 12807 7 2 2 49713 67552
0 12808 7 1 2 54954 72463
0 12809 5 1 1 12808
0 12810 7 1 2 12806 12809
0 12811 5 1 1 12810
0 12812 7 1 2 68900 12811
0 12813 5 1 1 12812
0 12814 7 3 2 51259 68463
0 12815 7 1 2 67475 68293
0 12816 7 1 2 66531 12815
0 12817 7 1 2 72465 12816
0 12818 5 1 1 12817
0 12819 7 1 2 12813 12818
0 12820 5 1 1 12819
0 12821 7 1 2 69694 12820
0 12822 5 1 1 12821
0 12823 7 1 2 12800 12822
0 12824 5 1 1 12823
0 12825 7 1 2 49028 12824
0 12826 5 1 1 12825
0 12827 7 2 2 50025 69865
0 12828 5 1 1 72468
0 12829 7 4 2 53784 55631
0 12830 7 1 2 52865 49308
0 12831 7 1 2 64432 12830
0 12832 7 1 2 72470 12831
0 12833 5 2 1 12832
0 12834 7 1 2 12828 72474
0 12835 5 1 1 12834
0 12836 7 1 2 72434 12835
0 12837 5 1 1 12836
0 12838 7 3 2 50977 71335
0 12839 7 1 2 61108 72476
0 12840 7 1 2 72288 12839
0 12841 5 1 1 12840
0 12842 7 1 2 12837 12841
0 12843 5 1 1 12842
0 12844 7 1 2 56891 12843
0 12845 5 1 1 12844
0 12846 7 5 2 50026 54243
0 12847 7 1 2 63719 72479
0 12848 7 1 2 69345 12847
0 12849 5 1 1 12848
0 12850 7 1 2 12845 12849
0 12851 5 1 1 12850
0 12852 7 1 2 49714 12851
0 12853 5 1 1 12852
0 12854 7 1 2 69445 69100
0 12855 7 1 2 61713 12854
0 12856 7 1 2 69301 12855
0 12857 5 1 1 12856
0 12858 7 1 2 12853 12857
0 12859 5 1 1 12858
0 12860 7 1 2 69695 12859
0 12861 5 1 1 12860
0 12862 7 1 2 12826 12861
0 12863 5 1 1 12862
0 12864 7 1 2 56705 12863
0 12865 5 1 1 12864
0 12866 7 1 2 12733 12865
0 12867 7 1 2 12626 12866
0 12868 5 1 1 12867
0 12869 7 1 2 63938 12868
0 12870 5 1 1 12869
0 12871 7 1 2 57991 69608
0 12872 5 1 1 12871
0 12873 7 1 2 65516 12872
0 12874 5 1 1 12873
0 12875 7 1 2 67315 69646
0 12876 7 1 2 12874 12875
0 12877 5 1 1 12876
0 12878 7 1 2 69990 12877
0 12879 5 1 1 12878
0 12880 7 6 2 47874 60191
0 12881 5 1 1 72484
0 12882 7 1 2 54955 12881
0 12883 5 1 1 12882
0 12884 7 2 2 66818 68524
0 12885 7 1 2 66203 72490
0 12886 7 1 2 12883 12885
0 12887 5 1 1 12886
0 12888 7 1 2 12879 12887
0 12889 5 1 1 12888
0 12890 7 1 2 51536 12889
0 12891 5 1 1 12890
0 12892 7 1 2 72051 72348
0 12893 5 1 1 12892
0 12894 7 2 2 53889 72289
0 12895 7 1 2 67437 70034
0 12896 7 1 2 72492 12895
0 12897 5 1 1 12896
0 12898 7 1 2 12893 12897
0 12899 5 1 1 12898
0 12900 7 1 2 50677 12899
0 12901 5 1 1 12900
0 12902 7 1 2 64626 67066
0 12903 5 1 1 12902
0 12904 7 3 2 54004 51260
0 12905 7 2 2 69561 72494
0 12906 5 1 1 72497
0 12907 7 1 2 65260 72498
0 12908 5 1 1 12907
0 12909 7 1 2 12903 12908
0 12910 5 1 1 12909
0 12911 7 1 2 67928 12910
0 12912 5 1 1 12911
0 12913 7 1 2 12901 12912
0 12914 7 1 2 12891 12913
0 12915 5 1 1 12914
0 12916 7 1 2 57460 12915
0 12917 5 1 1 12916
0 12918 7 1 2 70350 71729
0 12919 5 1 1 12918
0 12920 7 1 2 64290 68331
0 12921 5 1 1 12920
0 12922 7 1 2 72358 12921
0 12923 5 2 1 12922
0 12924 7 1 2 68063 72499
0 12925 5 1 1 12924
0 12926 7 1 2 12925 12431
0 12927 5 1 1 12926
0 12928 7 1 2 69067 12927
0 12929 5 1 1 12928
0 12930 7 1 2 12919 12929
0 12931 7 1 2 12917 12930
0 12932 5 1 1 12931
0 12933 7 1 2 50027 12932
0 12934 5 1 1 12933
0 12935 7 1 2 57582 68068
0 12936 5 2 1 12935
0 12937 7 2 2 60632 72501
0 12938 7 1 2 72346 72427
0 12939 7 1 2 72503 12938
0 12940 5 1 1 12939
0 12941 7 1 2 12934 12940
0 12942 5 1 1 12941
0 12943 7 1 2 49029 12942
0 12944 5 1 1 12943
0 12945 7 1 2 72378 72475
0 12946 5 2 1 12945
0 12947 7 1 2 72505 72504
0 12948 7 1 2 64081 72379
0 12949 5 1 1 12948
0 12950 7 1 2 12949 72382
0 12951 7 1 2 12947 12950
0 12952 5 1 1 12951
0 12953 7 1 2 12944 12952
0 12954 5 1 1 12953
0 12955 7 1 2 56706 12954
0 12956 5 1 1 12955
0 12957 7 3 2 54005 66079
0 12958 7 1 2 53785 69647
0 12959 5 3 1 12958
0 12960 7 1 2 72507 72510
0 12961 7 1 2 60960 12960
0 12962 5 1 1 12961
0 12963 7 1 2 51537 72204
0 12964 5 1 1 12963
0 12965 7 1 2 12962 12964
0 12966 5 1 1 12965
0 12967 7 1 2 49030 12966
0 12968 5 1 1 12967
0 12969 7 1 2 47875 67101
0 12970 7 2 2 48911 68343
0 12971 5 1 1 72513
0 12972 7 2 2 50028 53890
0 12973 7 2 2 59433 72515
0 12974 7 1 2 72514 72517
0 12975 7 1 2 12969 12974
0 12976 5 1 1 12975
0 12977 7 1 2 12968 12976
0 12978 5 1 1 12977
0 12979 7 1 2 69050 12978
0 12980 5 1 1 12979
0 12981 7 1 2 48912 72429
0 12982 5 1 1 12981
0 12983 7 1 2 72274 12982
0 12984 5 2 1 12983
0 12985 7 1 2 55277 57277
0 12986 7 1 2 72519 12985
0 12987 5 1 1 12986
0 12988 7 1 2 12980 12987
0 12989 5 1 1 12988
0 12990 7 1 2 56892 12989
0 12991 5 1 1 12990
0 12992 7 1 2 57913 72052
0 12993 5 1 1 12992
0 12994 7 1 2 60192 72290
0 12995 7 1 2 60995 12994
0 12996 5 1 1 12995
0 12997 7 1 2 12993 12996
0 12998 5 1 1 12997
0 12999 7 1 2 72105 12998
0 13000 5 1 1 12999
0 13001 7 1 2 12991 13000
0 13002 5 1 1 13001
0 13003 7 1 2 57461 13002
0 13004 5 1 1 13003
0 13005 7 1 2 51261 3546
0 13006 5 1 1 13005
0 13007 7 1 2 66366 13006
0 13008 5 1 1 13007
0 13009 7 1 2 65351 66080
0 13010 5 1 1 13009
0 13011 7 1 2 13008 13010
0 13012 5 1 1 13011
0 13013 7 1 2 69562 13012
0 13014 5 1 1 13013
0 13015 7 3 2 48601 63054
0 13016 7 1 2 65427 66429
0 13017 7 1 2 72521 13016
0 13018 5 1 1 13017
0 13019 7 1 2 13014 13018
0 13020 5 1 1 13019
0 13021 7 1 2 69264 13020
0 13022 5 1 1 13021
0 13023 7 1 2 13004 13022
0 13024 5 1 1 13023
0 13025 7 1 2 54578 13024
0 13026 5 1 1 13025
0 13027 7 2 2 56893 66741
0 13028 7 6 2 50678 51538
0 13029 7 2 2 68525 72526
0 13030 7 1 2 72524 72532
0 13031 5 1 1 13030
0 13032 7 1 2 48602 65331
0 13033 7 1 2 63370 13032
0 13034 7 1 2 71927 13033
0 13035 5 1 1 13034
0 13036 7 1 2 66114 13035
0 13037 5 1 1 13036
0 13038 7 1 2 57462 13037
0 13039 5 1 1 13038
0 13040 7 1 2 65352 66005
0 13041 5 1 1 13040
0 13042 7 1 2 68356 71399
0 13043 5 1 1 13042
0 13044 7 1 2 13041 13043
0 13045 7 1 2 13039 13044
0 13046 5 1 1 13045
0 13047 7 1 2 69563 13046
0 13048 5 1 1 13047
0 13049 7 6 2 54006 57463
0 13050 7 1 2 60969 72534
0 13051 5 1 1 13050
0 13052 7 1 2 56997 13051
0 13053 5 1 1 13052
0 13054 7 1 2 66467 67293
0 13055 7 1 2 13053 13054
0 13056 5 1 1 13055
0 13057 7 1 2 72359 13056
0 13058 7 1 2 13048 13057
0 13059 5 1 1 13058
0 13060 7 1 2 51733 13059
0 13061 5 1 1 13060
0 13062 7 1 2 13031 13061
0 13063 5 1 1 13062
0 13064 7 1 2 68235 13063
0 13065 5 1 1 13064
0 13066 7 1 2 13026 13065
0 13067 5 1 1 13066
0 13068 7 1 2 54956 13067
0 13069 5 1 1 13068
0 13070 7 2 2 68464 69285
0 13071 7 1 2 57914 63468
0 13072 5 1 1 13071
0 13073 7 3 2 50978 57464
0 13074 7 1 2 65545 72542
0 13075 7 1 2 71414 13074
0 13076 5 1 1 13075
0 13077 7 1 2 13072 13076
0 13078 5 1 1 13077
0 13079 7 1 2 72540 13078
0 13080 5 1 1 13079
0 13081 7 3 2 54244 65978
0 13082 7 1 2 64320 72545
0 13083 5 1 1 13082
0 13084 7 1 2 56894 71959
0 13085 5 1 1 13084
0 13086 7 1 2 13083 13085
0 13087 5 1 1 13086
0 13088 7 1 2 61934 13087
0 13089 5 1 1 13088
0 13090 7 1 2 66328 67421
0 13091 5 1 1 13090
0 13092 7 1 2 12429 13091
0 13093 5 1 1 13092
0 13094 7 1 2 57465 13093
0 13095 5 1 1 13094
0 13096 7 1 2 66011 71833
0 13097 5 1 1 13096
0 13098 7 1 2 56895 13097
0 13099 5 1 1 13098
0 13100 7 2 2 57915 66081
0 13101 5 1 1 72548
0 13102 7 1 2 13099 13101
0 13103 7 1 2 13095 13102
0 13104 7 1 2 13089 13103
0 13105 5 1 1 13104
0 13106 7 1 2 69564 13105
0 13107 5 1 1 13106
0 13108 7 2 2 51262 56998
0 13109 5 3 1 72550
0 13110 7 1 2 67773 72552
0 13111 5 1 1 13110
0 13112 7 1 2 66440 13111
0 13113 5 1 1 13112
0 13114 7 1 2 48913 13113
0 13115 5 1 1 13114
0 13116 7 1 2 57466 72500
0 13117 5 1 1 13116
0 13118 7 2 2 56896 65727
0 13119 5 1 1 72555
0 13120 7 1 2 64827 72556
0 13121 5 1 1 13120
0 13122 7 1 2 72360 13121
0 13123 5 1 1 13122
0 13124 7 1 2 54579 13123
0 13125 5 1 1 13124
0 13126 7 1 2 13117 13125
0 13127 5 1 1 13126
0 13128 7 1 2 54245 13127
0 13129 5 1 1 13128
0 13130 7 1 2 13115 13129
0 13131 7 1 2 13107 13130
0 13132 5 1 1 13131
0 13133 7 1 2 51734 13132
0 13134 5 1 1 13133
0 13135 7 1 2 13080 13134
0 13136 5 1 1 13135
0 13137 7 1 2 68236 13136
0 13138 5 1 1 13137
0 13139 7 2 2 48914 68220
0 13140 7 1 2 64342 72557
0 13141 7 1 2 69322 13140
0 13142 5 1 1 13141
0 13143 7 1 2 13138 13142
0 13144 7 1 2 13069 13143
0 13145 7 1 2 12956 13144
0 13146 5 1 1 13145
0 13147 7 1 2 62551 13146
0 13148 5 1 1 13147
0 13149 7 2 2 61935 69790
0 13150 5 1 1 72559
0 13151 7 1 2 48139 72560
0 13152 5 1 1 13151
0 13153 7 4 2 52085 59928
0 13154 5 3 1 72561
0 13155 7 1 2 68577 72565
0 13156 5 2 1 13155
0 13157 7 1 2 13152 72568
0 13158 5 1 1 13157
0 13159 7 1 2 69705 13158
0 13160 5 1 1 13159
0 13161 7 1 2 72566 72165
0 13162 5 1 1 13161
0 13163 7 1 2 13160 13162
0 13164 5 1 1 13163
0 13165 7 1 2 49892 13164
0 13166 5 1 1 13165
0 13167 7 1 2 48915 66171
0 13168 5 1 1 13167
0 13169 7 1 2 62471 13168
0 13170 5 1 1 13169
0 13171 7 1 2 49031 13170
0 13172 7 1 2 51263 72567
0 13173 5 1 1 13172
0 13174 7 1 2 65402 66581
0 13175 5 1 1 13174
0 13176 7 1 2 13173 13175
0 13177 5 1 1 13176
0 13178 7 7 2 51264 62951
0 13179 5 4 1 72570
0 13180 7 1 2 57916 72577
0 13181 5 1 1 13180
0 13182 7 1 2 52783 2790
0 13183 7 1 2 13181 13182
0 13184 5 1 1 13183
0 13185 7 1 2 13177 13184
0 13186 7 1 2 13171 13185
0 13187 5 1 1 13186
0 13188 7 1 2 13166 13187
0 13189 5 1 1 13188
0 13190 7 1 2 55500 13189
0 13191 5 1 1 13190
0 13192 7 1 2 65288 72122
0 13193 5 1 1 13192
0 13194 7 1 2 13191 13193
0 13195 5 1 1 13194
0 13196 7 1 2 54580 13195
0 13197 5 1 1 13196
0 13198 7 1 2 58423 60263
0 13199 5 2 1 13198
0 13200 7 2 2 55278 72581
0 13201 5 1 1 72583
0 13202 7 1 2 49032 72584
0 13203 7 1 2 72120 13202
0 13204 5 1 1 13203
0 13205 7 1 2 13197 13204
0 13206 5 1 1 13205
0 13207 7 1 2 50029 13206
0 13208 5 1 1 13207
0 13209 7 1 2 48140 69438
0 13210 7 1 2 69741 13209
0 13211 5 1 1 13210
0 13212 7 1 2 72569 13211
0 13213 5 1 1 13212
0 13214 7 1 2 67828 72023
0 13215 7 1 2 69696 13214
0 13216 7 1 2 13213 13215
0 13217 5 1 1 13216
0 13218 7 1 2 13208 13217
0 13219 5 1 1 13218
0 13220 7 1 2 71933 13219
0 13221 5 1 1 13220
0 13222 7 1 2 64461 68069
0 13223 5 1 1 13222
0 13224 7 1 2 57917 13223
0 13225 5 1 1 13224
0 13226 7 1 2 68064 71812
0 13227 5 1 1 13226
0 13228 7 1 2 13225 13227
0 13229 5 1 1 13228
0 13230 7 1 2 56897 13229
0 13231 5 1 1 13230
0 13232 7 3 2 54246 10404
0 13233 5 1 1 72585
0 13234 7 1 2 7222 13233
0 13235 5 1 1 13234
0 13236 7 1 2 64452 13235
0 13237 5 1 1 13236
0 13238 7 1 2 13231 13237
0 13239 5 1 1 13238
0 13240 7 1 2 72218 13239
0 13241 5 1 1 13240
0 13242 7 1 2 70057 72207
0 13243 5 1 1 13242
0 13244 7 1 2 13241 13243
0 13245 5 1 1 13244
0 13246 7 1 2 51265 13245
0 13247 5 1 1 13246
0 13248 7 3 2 48916 68804
0 13249 7 1 2 68237 72588
0 13250 5 1 1 13249
0 13251 7 1 2 13247 13250
0 13252 5 1 1 13251
0 13253 7 1 2 55501 13252
0 13254 5 1 1 13253
0 13255 7 13 2 51539 68238
0 13256 7 1 2 66198 65858
0 13257 5 1 1 13256
0 13258 7 1 2 72235 13257
0 13259 5 1 1 13258
0 13260 7 1 2 70006 13259
0 13261 5 1 1 13260
0 13262 7 1 2 72591 13261
0 13263 5 1 1 13262
0 13264 7 1 2 13254 13263
0 13265 7 1 2 13221 13264
0 13266 5 1 1 13265
0 13267 7 1 2 51735 13266
0 13268 5 1 1 13267
0 13269 7 1 2 61898 58285
0 13270 5 2 1 13269
0 13271 7 1 2 50679 68070
0 13272 5 1 1 13271
0 13273 7 1 2 57467 13272
0 13274 5 1 1 13273
0 13275 7 1 2 72604 13274
0 13276 5 1 1 13275
0 13277 7 1 2 56898 13276
0 13278 5 1 1 13277
0 13279 7 3 2 52943 60531
0 13280 5 2 1 72606
0 13281 7 1 2 55279 72609
0 13282 5 1 1 13281
0 13283 7 1 2 13278 13282
0 13284 5 1 1 13283
0 13285 7 1 2 54957 13284
0 13286 5 1 1 13285
0 13287 7 1 2 57468 72586
0 13288 5 1 1 13287
0 13289 7 1 2 56999 13288
0 13290 5 1 1 13289
0 13291 7 1 2 55280 13290
0 13292 5 1 1 13291
0 13293 7 1 2 13286 13292
0 13294 5 1 1 13293
0 13295 7 1 2 62905 72520
0 13296 5 1 1 13295
0 13297 7 1 2 48917 72272
0 13298 5 1 1 13297
0 13299 7 1 2 13296 13298
0 13300 5 1 1 13299
0 13301 7 1 2 13294 13300
0 13302 5 1 1 13301
0 13303 7 2 2 62322 65243
0 13304 7 1 2 65439 72611
0 13305 5 1 1 13304
0 13306 7 1 2 13201 13305
0 13307 5 1 1 13306
0 13308 7 2 2 65625 68208
0 13309 7 4 2 68767 72613
0 13310 7 2 2 69143 72615
0 13311 5 1 1 72619
0 13312 7 1 2 57918 71934
0 13313 7 1 2 72620 13312
0 13314 7 1 2 13307 13313
0 13315 5 1 1 13314
0 13316 7 1 2 13302 13315
0 13317 7 1 2 13268 13316
0 13318 7 1 2 13148 13317
0 13319 7 1 2 12870 13318
0 13320 7 1 2 12466 13319
0 13321 7 1 2 12081 13320
0 13322 7 3 2 57992 57361
0 13323 5 1 1 72621
0 13324 7 1 2 63774 71551
0 13325 7 1 2 57213 70707
0 13326 5 1 1 13325
0 13327 7 1 2 56707 60006
0 13328 5 1 1 13327
0 13329 7 1 2 55683 13328
0 13330 5 1 1 13329
0 13331 7 1 2 13326 13330
0 13332 7 1 2 13324 13331
0 13333 5 1 1 13332
0 13334 7 1 2 52260 13333
0 13335 5 1 1 13334
0 13336 7 1 2 50395 59852
0 13337 5 2 1 13336
0 13338 7 1 2 70791 72624
0 13339 5 1 1 13338
0 13340 7 1 2 52086 13339
0 13341 5 1 1 13340
0 13342 7 2 2 70354 13341
0 13343 5 2 1 72626
0 13344 7 4 2 51875 72628
0 13345 5 2 1 72630
0 13346 7 1 2 70214 70995
0 13347 5 1 1 13346
0 13348 7 1 2 60781 57278
0 13349 7 1 2 63775 13348
0 13350 5 1 1 13349
0 13351 7 1 2 53074 13350
0 13352 5 1 1 13351
0 13353 7 1 2 13347 13352
0 13354 7 1 2 72634 13353
0 13355 7 3 2 13335 13354
0 13356 7 1 2 13323 72636
0 13357 5 1 1 13356
0 13358 7 1 2 61334 13357
0 13359 5 1 1 13358
0 13360 7 1 2 49715 13359
0 13361 5 1 1 13360
0 13362 7 1 2 58972 72477
0 13363 7 1 2 13361 13362
0 13364 5 1 1 13363
0 13365 7 1 2 53786 69697
0 13366 5 2 1 13365
0 13367 7 1 2 72100 72639
0 13368 5 1 1 13367
0 13369 7 2 2 57151 61948
0 13370 7 1 2 64327 72641
0 13371 7 1 2 13368 13370
0 13372 5 1 1 13371
0 13373 7 1 2 13364 13372
0 13374 5 1 1 13373
0 13375 7 1 2 54581 13374
0 13376 5 1 1 13375
0 13377 7 1 2 71707 72502
0 13378 5 1 1 13377
0 13379 7 1 2 69125 71695
0 13380 5 1 1 13379
0 13381 7 1 2 13378 13380
0 13382 5 1 1 13381
0 13383 7 1 2 71336 13382
0 13384 5 1 1 13383
0 13385 7 1 2 13376 13384
0 13386 5 1 1 13385
0 13387 7 1 2 51540 13386
0 13388 5 1 1 13387
0 13389 7 3 2 50030 55502
0 13390 7 1 2 54582 72637
0 13391 5 1 1 13390
0 13392 7 1 2 71058 13391
0 13393 5 1 1 13392
0 13394 7 7 2 52261 50680
0 13395 7 2 2 59653 72646
0 13396 5 2 1 72653
0 13397 7 2 2 72654 70801
0 13398 5 1 1 72657
0 13399 7 1 2 70124 72658
0 13400 5 1 1 13399
0 13401 7 2 2 60293 59828
0 13402 5 1 1 72659
0 13403 7 1 2 59853 60142
0 13404 5 1 1 13403
0 13405 7 1 2 72660 13404
0 13406 5 1 1 13405
0 13407 7 1 2 57583 13406
0 13408 5 1 1 13407
0 13409 7 2 2 55855 64487
0 13410 5 2 1 72661
0 13411 7 2 2 54583 9475
0 13412 5 2 1 72665
0 13413 7 1 2 72663 72666
0 13414 7 1 2 13408 13413
0 13415 5 1 1 13414
0 13416 7 1 2 50396 13415
0 13417 5 1 1 13416
0 13418 7 2 2 52262 60046
0 13419 7 1 2 72562 72669
0 13420 5 1 1 13419
0 13421 7 1 2 60616 70424
0 13422 5 2 1 13421
0 13423 7 1 2 59854 72671
0 13424 5 1 1 13423
0 13425 7 1 2 13420 13424
0 13426 7 1 2 50681 60047
0 13427 5 1 1 13426
0 13428 7 2 2 54958 13427
0 13429 5 1 1 72673
0 13430 7 1 2 48141 71164
0 13431 5 3 1 13430
0 13432 7 5 2 52263 58816
0 13433 5 1 1 72678
0 13434 7 1 2 54584 13433
0 13435 5 4 1 13434
0 13436 7 2 2 72675 72683
0 13437 5 1 1 72687
0 13438 7 1 2 50168 72688
0 13439 5 1 1 13438
0 13440 7 1 2 60028 71446
0 13441 5 1 1 13440
0 13442 7 1 2 13439 13441
0 13443 7 1 2 72674 13442
0 13444 7 1 2 13425 13443
0 13445 7 1 2 13417 13444
0 13446 5 1 1 13445
0 13447 7 1 2 70163 13446
0 13448 5 1 1 13447
0 13449 7 1 2 13400 13448
0 13450 7 1 2 13393 13449
0 13451 5 1 1 13450
0 13452 7 1 2 62472 13451
0 13453 5 1 1 13452
0 13454 7 1 2 59794 60143
0 13455 5 1 1 13454
0 13456 7 1 2 71005 13455
0 13457 5 1 1 13456
0 13458 7 1 2 50397 13457
0 13459 5 1 1 13458
0 13460 7 5 2 52264 52883
0 13461 7 2 2 51876 72689
0 13462 7 3 2 59740 59817
0 13463 5 1 1 72696
0 13464 7 1 2 72694 72697
0 13465 5 1 1 13464
0 13466 7 1 2 13459 13465
0 13467 7 1 2 70927 13466
0 13468 5 1 1 13467
0 13469 7 2 2 49716 71524
0 13470 5 3 1 72699
0 13471 7 19 2 58743 72701
0 13472 5 3 1 72704
0 13473 7 3 2 56189 72705
0 13474 5 1 1 72726
0 13475 7 1 2 58973 13474
0 13476 5 1 1 13475
0 13477 7 1 2 59130 13476
0 13478 7 1 2 13468 13477
0 13479 5 1 1 13478
0 13480 7 1 2 13453 13479
0 13481 5 1 1 13480
0 13482 7 1 2 69648 13481
0 13483 5 1 1 13482
0 13484 7 1 2 62952 60334
0 13485 5 1 1 13484
0 13486 7 4 2 65000 59131
0 13487 5 1 1 72729
0 13488 7 2 2 13485 13487
0 13489 5 1 1 72733
0 13490 7 2 2 59929 59132
0 13491 5 3 1 72735
0 13492 7 1 2 52087 62953
0 13493 5 2 1 13492
0 13494 7 1 2 72737 72740
0 13495 5 1 1 13494
0 13496 7 1 2 55684 13495
0 13497 5 1 1 13496
0 13498 7 1 2 72734 13497
0 13499 5 1 1 13498
0 13500 7 1 2 52265 13499
0 13501 5 1 1 13500
0 13502 7 1 2 51877 13489
0 13503 5 1 1 13502
0 13504 7 1 2 63651 13503
0 13505 5 2 1 13504
0 13506 7 1 2 55685 72742
0 13507 5 1 1 13506
0 13508 7 1 2 13501 13507
0 13509 5 1 1 13508
0 13510 7 1 2 52944 13509
0 13511 5 1 1 13510
0 13512 7 1 2 67465 70552
0 13513 5 1 1 13512
0 13514 7 1 2 13511 13513
0 13515 5 1 1 13514
0 13516 7 1 2 53075 13515
0 13517 5 1 1 13516
0 13518 7 1 2 59741 72730
0 13519 5 1 1 13518
0 13520 7 1 2 62954 9491
0 13521 5 1 1 13520
0 13522 7 1 2 59133 70921
0 13523 5 1 1 13522
0 13524 7 1 2 13521 13523
0 13525 5 1 1 13524
0 13526 7 1 2 52266 13525
0 13527 5 1 1 13526
0 13528 7 1 2 13519 13527
0 13529 5 1 1 13528
0 13530 7 1 2 59855 13529
0 13531 5 1 1 13530
0 13532 7 2 2 50398 61625
0 13533 5 1 1 72744
0 13534 7 1 2 54585 13533
0 13535 5 1 1 13534
0 13536 7 2 2 52088 13535
0 13537 5 1 1 72746
0 13538 7 1 2 65943 13537
0 13539 5 1 1 13538
0 13540 7 1 2 59856 13539
0 13541 5 1 1 13540
0 13542 7 1 2 50682 60357
0 13543 5 2 1 13542
0 13544 7 1 2 48142 72748
0 13545 5 1 1 13544
0 13546 7 1 2 50169 58335
0 13547 7 1 2 13545 13546
0 13548 5 1 1 13547
0 13549 7 1 2 54959 67430
0 13550 7 1 2 13548 13549
0 13551 7 1 2 13541 13550
0 13552 5 1 1 13551
0 13553 7 1 2 62955 13552
0 13554 5 1 1 13553
0 13555 7 1 2 52267 72743
0 13556 5 1 1 13555
0 13557 7 1 2 62956 70491
0 13558 5 1 1 13557
0 13559 7 1 2 13556 13558
0 13560 5 1 1 13559
0 13561 7 1 2 60048 13560
0 13562 5 1 1 13561
0 13563 7 1 2 13554 13562
0 13564 7 1 2 13531 13563
0 13565 7 1 2 13517 13564
0 13566 5 1 1 13565
0 13567 7 1 2 61335 13566
0 13568 5 1 1 13567
0 13569 7 2 2 50088 50683
0 13570 7 4 2 52884 53076
0 13571 5 1 1 72752
0 13572 7 5 2 52268 72753
0 13573 5 1 1 72756
0 13574 7 1 2 72750 72757
0 13575 5 1 1 13574
0 13576 7 1 2 54960 13575
0 13577 5 2 1 13576
0 13578 7 1 2 52089 72761
0 13579 5 1 1 13578
0 13580 7 1 2 71231 13579
0 13581 5 1 1 13580
0 13582 7 1 2 70717 13581
0 13583 5 1 1 13582
0 13584 7 1 2 57584 64488
0 13585 5 1 1 13584
0 13586 7 1 2 62664 13585
0 13587 5 1 1 13586
0 13588 7 1 2 50979 13587
0 13589 5 1 1 13588
0 13590 7 6 2 50684 55856
0 13591 5 1 1 72763
0 13592 7 2 2 61691 72764
0 13593 5 1 1 72769
0 13594 7 2 2 50980 60116
0 13595 5 1 1 72771
0 13596 7 1 2 61517 65228
0 13597 5 2 1 13596
0 13598 7 1 2 13595 72773
0 13599 5 1 1 13598
0 13600 7 1 2 55686 13599
0 13601 5 1 1 13600
0 13602 7 1 2 13593 13601
0 13603 7 1 2 13589 13602
0 13604 7 1 2 13583 13603
0 13605 5 1 1 13604
0 13606 7 1 2 50399 13605
0 13607 5 1 1 13606
0 13608 7 1 2 50170 70822
0 13609 5 1 1 13608
0 13610 7 1 2 70651 13609
0 13611 5 2 1 13610
0 13612 7 1 2 55687 72775
0 13613 5 1 1 13612
0 13614 7 1 2 63129 59306
0 13615 5 1 1 13614
0 13616 7 1 2 54586 13615
0 13617 7 1 2 13613 13616
0 13618 5 1 1 13617
0 13619 7 1 2 50981 13618
0 13620 5 1 1 13619
0 13621 7 1 2 13607 13620
0 13622 5 1 1 13621
0 13623 7 1 2 70954 13622
0 13624 5 1 1 13623
0 13625 7 1 2 61180 70718
0 13626 5 1 1 13625
0 13627 7 1 2 61548 62113
0 13628 7 1 2 13626 13627
0 13629 5 1 1 13628
0 13630 7 1 2 57585 13629
0 13631 5 1 1 13630
0 13632 7 1 2 56062 70792
0 13633 5 1 1 13632
0 13634 7 1 2 52090 13633
0 13635 5 1 1 13634
0 13636 7 1 2 55857 61807
0 13637 5 1 1 13636
0 13638 7 1 2 54587 13637
0 13639 7 1 2 13635 13638
0 13640 7 1 2 13631 13639
0 13641 5 1 1 13640
0 13642 7 1 2 50400 13641
0 13643 5 1 1 13642
0 13644 7 2 2 50171 61256
0 13645 5 6 1 72777
0 13646 7 2 2 54588 72779
0 13647 5 2 1 72785
0 13648 7 1 2 57586 72787
0 13649 5 1 1 13648
0 13650 7 7 2 65101 65463
0 13651 7 3 2 55858 55688
0 13652 5 1 1 72796
0 13653 7 1 2 54589 13652
0 13654 5 3 1 13653
0 13655 7 1 2 72789 72799
0 13656 5 1 1 13655
0 13657 7 1 2 56618 59758
0 13658 5 2 1 13657
0 13659 7 1 2 54961 72802
0 13660 7 1 2 13656 13659
0 13661 7 1 2 13649 13660
0 13662 7 1 2 13643 13661
0 13663 5 1 1 13662
0 13664 7 1 2 70164 13663
0 13665 5 1 1 13664
0 13666 7 1 2 70165 9947
0 13667 5 1 1 13666
0 13668 7 1 2 60036 71503
0 13669 5 1 1 13668
0 13670 7 1 2 13667 13669
0 13671 5 1 1 13670
0 13672 7 1 2 57214 13671
0 13673 5 1 1 13672
0 13674 7 1 2 70314 13673
0 13675 7 1 2 13665 13674
0 13676 7 1 2 13624 13675
0 13677 7 1 2 13568 13676
0 13678 5 1 1 13677
0 13679 7 1 2 69521 13678
0 13680 5 1 1 13679
0 13681 7 1 2 13483 13680
0 13682 5 1 1 13681
0 13683 7 1 2 72643 13682
0 13684 5 1 1 13683
0 13685 7 1 2 13388 13684
0 13686 5 1 1 13685
0 13687 7 1 2 55632 13686
0 13688 5 1 1 13687
0 13689 7 1 2 61320 72638
0 13690 5 1 1 13689
0 13691 7 1 2 68768 13690
0 13692 5 1 1 13691
0 13693 7 1 2 65120 59372
0 13694 7 1 2 70013 13693
0 13695 5 1 1 13694
0 13696 7 1 2 13692 13695
0 13697 5 1 1 13696
0 13698 7 1 2 50982 13697
0 13699 5 1 1 13698
0 13700 7 2 2 67136 68849
0 13701 5 1 1 72804
0 13702 7 1 2 57993 65040
0 13703 5 1 1 13702
0 13704 7 1 2 13701 13703
0 13705 5 1 1 13704
0 13706 7 1 2 61336 70965
0 13707 5 1 1 13706
0 13708 7 1 2 67163 70120
0 13709 7 1 2 13398 13708
0 13710 7 1 2 13707 13709
0 13711 5 1 1 13710
0 13712 7 1 2 69237 13711
0 13713 5 1 1 13712
0 13714 7 1 2 13705 13713
0 13715 7 1 2 13699 13714
0 13716 5 1 1 13715
0 13717 7 1 2 50031 13716
0 13718 5 1 1 13717
0 13719 7 1 2 57919 69498
0 13720 5 1 1 13719
0 13721 7 1 2 57469 62765
0 13722 5 1 1 13721
0 13723 7 1 2 13720 13722
0 13724 5 1 1 13723
0 13725 7 2 2 48725 49430
0 13726 7 7 2 65649 72806
0 13727 7 1 2 68953 72808
0 13728 7 1 2 13724 13727
0 13729 5 1 1 13728
0 13730 7 1 2 13718 13729
0 13731 5 1 1 13730
0 13732 7 1 2 67929 13731
0 13733 5 1 1 13732
0 13734 7 1 2 13688 13733
0 13735 5 1 1 13734
0 13736 7 1 2 49033 13735
0 13737 5 1 1 13736
0 13738 7 2 2 72480 72809
0 13739 7 1 2 58800 69346
0 13740 5 1 1 13739
0 13741 7 2 2 68749 68465
0 13742 7 1 2 64765 63979
0 13743 7 1 2 72817 13742
0 13744 5 1 1 13743
0 13745 7 1 2 13740 13744
0 13746 5 1 1 13745
0 13747 7 1 2 72543 13746
0 13748 5 1 1 13747
0 13749 7 1 2 69821 72333
0 13750 5 1 1 13749
0 13751 7 1 2 13748 13750
0 13752 5 1 1 13751
0 13753 7 1 2 72815 13752
0 13754 5 1 1 13753
0 13755 7 1 2 56899 72587
0 13756 5 1 1 13755
0 13757 7 1 2 58071 13756
0 13758 5 1 1 13757
0 13759 7 1 2 52784 13758
0 13760 5 1 1 13759
0 13761 7 1 2 48726 70121
0 13762 5 6 1 13761
0 13763 7 1 2 72819 70966
0 13764 5 1 1 13763
0 13765 7 1 2 52269 71040
0 13766 5 1 1 13765
0 13767 7 1 2 48727 13766
0 13768 5 1 1 13767
0 13769 7 1 2 61337 13768
0 13770 5 1 1 13769
0 13771 7 1 2 70972 13770
0 13772 7 1 2 13764 13771
0 13773 5 1 1 13772
0 13774 7 1 2 49717 13773
0 13775 5 1 1 13774
0 13776 7 1 2 13760 13775
0 13777 5 1 1 13776
0 13778 7 1 2 72106 68466
0 13779 7 1 2 13777 13778
0 13780 5 1 1 13779
0 13781 7 1 2 69117 72227
0 13782 5 1 1 13781
0 13783 7 1 2 13311 13782
0 13784 5 1 1 13783
0 13785 7 1 2 56900 57279
0 13786 7 1 2 13784 13785
0 13787 5 1 1 13786
0 13788 7 2 2 71928 69731
0 13789 7 2 2 48143 49034
0 13790 7 1 2 72827 72518
0 13791 7 1 2 72825 13790
0 13792 5 1 1 13791
0 13793 7 1 2 13787 13792
0 13794 5 1 1 13793
0 13795 7 1 2 54590 13794
0 13796 5 1 1 13795
0 13797 7 1 2 71337 71567
0 13798 5 2 1 13797
0 13799 7 1 2 72829 72640
0 13800 5 1 1 13799
0 13801 7 1 2 71701 13800
0 13802 5 1 1 13801
0 13803 7 1 2 67263 69941
0 13804 5 1 1 13803
0 13805 7 1 2 72258 13804
0 13806 5 1 1 13805
0 13807 7 1 2 48728 13806
0 13808 5 1 1 13807
0 13809 7 1 2 50032 71181
0 13810 5 1 1 13809
0 13811 7 1 2 13808 13810
0 13812 5 1 1 13811
0 13813 7 1 2 67930 68065
0 13814 7 1 2 13812 13813
0 13815 5 1 1 13814
0 13816 7 1 2 13802 13815
0 13817 5 1 1 13816
0 13818 7 1 2 49035 13817
0 13819 5 1 1 13818
0 13820 7 2 2 47876 69347
0 13821 5 1 1 72831
0 13822 7 1 2 61936 72832
0 13823 5 1 1 13822
0 13824 7 1 2 11879 13823
0 13825 5 1 1 13824
0 13826 7 1 2 69446 69698
0 13827 7 1 2 13825 13826
0 13828 5 1 1 13827
0 13829 7 1 2 13819 13828
0 13830 7 1 2 13796 13829
0 13831 5 1 1 13830
0 13832 7 1 2 57470 13831
0 13833 5 1 1 13832
0 13834 7 2 2 68239 68823
0 13835 5 2 1 72833
0 13836 7 2 2 69615 72095
0 13837 5 1 1 72837
0 13838 7 1 2 57920 72838
0 13839 5 1 1 13838
0 13840 7 1 2 72835 13839
0 13841 5 1 1 13840
0 13842 7 1 2 48729 13841
0 13843 5 1 1 13842
0 13844 7 1 2 68778 72208
0 13845 5 1 1 13844
0 13846 7 1 2 13843 13845
0 13847 5 1 1 13846
0 13848 7 1 2 57000 64411
0 13849 7 1 2 72605 13848
0 13850 5 1 1 13849
0 13851 7 1 2 67931 13850
0 13852 7 1 2 13847 13851
0 13853 5 1 1 13852
0 13854 7 1 2 13833 13853
0 13855 7 1 2 13780 13854
0 13856 5 1 1 13855
0 13857 7 1 2 54962 13856
0 13858 5 1 1 13857
0 13859 7 1 2 13754 13858
0 13860 7 1 2 13737 13859
0 13861 5 1 1 13860
0 13862 7 1 2 55281 13861
0 13863 5 1 1 13862
0 13864 7 5 2 50172 62632
0 13865 5 1 1 72839
0 13866 7 1 2 58384 63239
0 13867 5 1 1 13866
0 13868 7 1 2 13865 13867
0 13869 5 2 1 13868
0 13870 7 1 2 64740 72844
0 13871 5 1 1 13870
0 13872 7 1 2 61899 59117
0 13873 5 1 1 13872
0 13874 7 1 2 13871 13873
0 13875 5 1 1 13874
0 13876 7 1 2 51266 13875
0 13877 5 1 1 13876
0 13878 7 1 2 61900 59000
0 13879 5 1 1 13878
0 13880 7 1 2 13877 13879
0 13881 5 1 1 13880
0 13882 7 1 2 54963 13881
0 13883 5 1 1 13882
0 13884 7 1 2 72450 13150
0 13885 5 1 1 13884
0 13886 7 1 2 71638 13885
0 13887 5 1 1 13886
0 13888 7 1 2 13883 13887
0 13889 5 1 1 13888
0 13890 7 1 2 51541 13889
0 13891 5 1 1 13890
0 13892 7 1 2 66273 71687
0 13893 5 1 1 13892
0 13894 7 1 2 13891 13893
0 13895 5 1 1 13894
0 13896 7 1 2 55633 13895
0 13897 5 1 1 13896
0 13898 7 3 2 63088 67932
0 13899 7 1 2 64627 72846
0 13900 5 1 1 13899
0 13901 7 1 2 13897 13900
0 13902 5 1 1 13901
0 13903 7 1 2 53672 13902
0 13904 5 1 1 13903
0 13905 7 2 2 60386 67182
0 13906 7 1 2 57921 60970
0 13907 7 1 2 72849 13906
0 13908 5 1 1 13907
0 13909 7 1 2 68440 13908
0 13910 5 1 1 13909
0 13911 7 1 2 65703 13910
0 13912 5 1 1 13911
0 13913 7 1 2 53891 68443
0 13914 7 1 2 72522 13913
0 13915 5 1 1 13914
0 13916 7 1 2 13912 13915
0 13917 5 1 1 13916
0 13918 7 1 2 70014 13917
0 13919 5 1 1 13918
0 13920 7 1 2 64628 71709
0 13921 5 1 1 13920
0 13922 7 5 2 51542 70064
0 13923 5 3 1 72851
0 13924 7 2 2 65523 64607
0 13925 5 1 1 72859
0 13926 7 1 2 57994 72860
0 13927 5 1 1 13926
0 13928 7 1 2 72852 13927
0 13929 5 1 1 13928
0 13930 7 1 2 13921 13929
0 13931 7 1 2 13919 13930
0 13932 5 1 1 13931
0 13933 7 1 2 51736 13932
0 13934 5 1 1 13933
0 13935 7 1 2 13904 13934
0 13936 5 1 1 13935
0 13937 7 1 2 50033 13936
0 13938 5 1 1 13937
0 13939 7 2 2 69026 69680
0 13940 5 1 1 72861
0 13941 7 1 2 53787 72862
0 13942 5 1 1 13941
0 13943 7 1 2 53788 69919
0 13944 5 1 1 13943
0 13945 7 1 2 47877 68769
0 13946 7 1 2 72436 13945
0 13947 5 1 1 13946
0 13948 7 1 2 13944 13947
0 13949 5 1 1 13948
0 13950 7 1 2 61937 66451
0 13951 7 1 2 13949 13950
0 13952 5 1 1 13951
0 13953 7 1 2 13942 13952
0 13954 5 1 1 13953
0 13955 7 1 2 55282 13954
0 13956 5 1 1 13955
0 13957 7 1 2 64508 72845
0 13958 5 1 1 13957
0 13959 7 1 2 10815 13958
0 13960 5 2 1 13959
0 13961 7 1 2 68859 72863
0 13962 5 1 1 13961
0 13963 7 1 2 61901 67933
0 13964 7 1 2 68997 13963
0 13965 5 1 1 13964
0 13966 7 1 2 13962 13965
0 13967 5 1 1 13966
0 13968 7 1 2 68578 13967
0 13969 5 1 1 13968
0 13970 7 1 2 13956 13969
0 13971 5 1 1 13970
0 13972 7 1 2 57922 13971
0 13973 5 1 1 13972
0 13974 7 2 2 62766 72053
0 13975 7 2 2 49893 56901
0 13976 7 1 2 72865 72867
0 13977 5 1 1 13976
0 13978 7 1 2 13973 13977
0 13979 5 1 1 13978
0 13980 7 1 2 65626 13979
0 13981 5 1 1 13980
0 13982 7 1 2 13938 13981
0 13983 5 1 1 13982
0 13984 7 1 2 49036 13983
0 13985 5 1 1 13984
0 13986 7 4 2 71338 69907
0 13987 7 1 2 72869 72864
0 13988 5 1 1 13987
0 13989 7 1 2 13925 69403
0 13990 5 1 1 13989
0 13991 7 1 2 13988 13990
0 13992 5 1 1 13991
0 13993 7 1 2 55634 13992
0 13994 5 1 1 13993
0 13995 7 1 2 64920 68624
0 13996 5 1 1 13995
0 13997 7 1 2 71834 13996
0 13998 5 1 1 13997
0 13999 7 1 2 58385 68344
0 14000 7 1 2 69168 13999
0 14001 7 1 2 13998 14000
0 14002 5 1 1 14001
0 14003 7 1 2 13994 14002
0 14004 5 1 1 14003
0 14005 7 1 2 49718 14004
0 14006 5 1 1 14005
0 14007 7 4 2 55635 69406
0 14008 7 1 2 48501 72873
0 14009 7 2 2 49431 61902
0 14010 5 1 1 72877
0 14011 7 1 2 72175 72878
0 14012 7 1 2 14008 14011
0 14013 5 1 1 14012
0 14014 7 1 2 13940 14013
0 14015 5 1 1 14014
0 14016 7 1 2 50034 69791
0 14017 7 1 2 14015 14016
0 14018 5 1 1 14017
0 14019 7 1 2 14006 14018
0 14020 5 1 1 14019
0 14021 7 1 2 57923 14020
0 14022 5 1 1 14021
0 14023 7 2 2 61658 64509
0 14024 5 1 1 72879
0 14025 7 1 2 69294 69855
0 14026 7 1 2 72880 14025
0 14027 5 1 1 14026
0 14028 7 1 2 72380 14027
0 14029 5 1 1 14028
0 14030 7 1 2 72868 69673
0 14031 7 1 2 14029 14030
0 14032 5 1 1 14031
0 14033 7 1 2 14022 14032
0 14034 5 1 1 14033
0 14035 7 1 2 65627 14034
0 14036 5 1 1 14035
0 14037 7 1 2 13985 14036
0 14038 5 1 1 14037
0 14039 7 1 2 57471 14038
0 14040 5 1 1 14039
0 14041 7 5 2 49719 65979
0 14042 5 1 1 72881
0 14043 7 1 2 66311 68066
0 14044 5 1 1 14043
0 14045 7 1 2 14042 14044
0 14046 5 1 1 14045
0 14047 7 1 2 52785 14046
0 14048 5 1 1 14047
0 14049 7 5 2 55283 59350
0 14050 5 1 1 72886
0 14051 7 1 2 66993 72887
0 14052 5 1 1 14051
0 14053 7 1 2 14048 14052
0 14054 5 1 1 14053
0 14055 7 1 2 68549 14054
0 14056 5 1 1 14055
0 14057 7 5 2 47878 61659
0 14058 5 2 1 72891
0 14059 7 1 2 72523 72892
0 14060 7 1 2 72853 14059
0 14061 5 1 1 14060
0 14062 7 1 2 71400 71973
0 14063 5 1 1 14062
0 14064 7 1 2 72451 14063
0 14065 5 1 1 14064
0 14066 7 1 2 66537 70015
0 14067 7 1 2 14065 14066
0 14068 5 1 1 14067
0 14069 7 1 2 14061 14068
0 14070 5 1 1 14069
0 14071 7 1 2 51737 14070
0 14072 5 1 1 14071
0 14073 7 1 2 14056 14072
0 14074 5 1 1 14073
0 14075 7 1 2 54247 14074
0 14076 5 1 1 14075
0 14077 7 1 2 52786 64592
0 14078 5 2 1 14077
0 14079 7 1 2 50685 72448
0 14080 5 1 1 14079
0 14081 7 1 2 72898 14080
0 14082 5 1 1 14081
0 14083 7 1 2 56902 69332
0 14084 7 1 2 14082 14083
0 14085 5 1 1 14084
0 14086 7 1 2 14076 14085
0 14087 5 1 1 14086
0 14088 7 1 2 68240 14087
0 14089 5 1 1 14088
0 14090 7 1 2 66798 69388
0 14091 5 1 1 14090
0 14092 7 1 2 61938 72037
0 14093 7 1 2 69589 14092
0 14094 5 1 1 14093
0 14095 7 1 2 14091 14094
0 14096 5 1 1 14095
0 14097 7 1 2 67513 72558
0 14098 7 1 2 14096 14097
0 14099 5 1 1 14098
0 14100 7 1 2 14089 14099
0 14101 7 1 2 14040 14100
0 14102 5 1 1 14101
0 14103 7 1 2 56708 14102
0 14104 5 1 1 14103
0 14105 7 1 2 13863 14104
0 14106 7 1 2 13321 14105
0 14107 7 1 2 10805 14106
0 14108 7 1 2 9200 14107
0 14109 7 6 2 49894 68279
0 14110 7 2 2 50173 59373
0 14111 5 2 1 72906
0 14112 7 1 2 50401 72776
0 14113 5 1 1 14112
0 14114 7 1 2 61626 70434
0 14115 5 3 1 14114
0 14116 7 1 2 14113 72910
0 14117 5 1 1 14116
0 14118 7 1 2 54591 14117
0 14119 5 1 1 14118
0 14120 7 1 2 72908 14119
0 14121 5 1 1 14120
0 14122 7 1 2 61447 14121
0 14123 5 1 1 14122
0 14124 7 1 2 56190 59913
0 14125 5 2 1 14124
0 14126 7 1 2 70786 70290
0 14127 5 1 1 14126
0 14128 7 1 2 72913 14127
0 14129 5 1 1 14128
0 14130 7 1 2 50174 14129
0 14131 5 1 1 14130
0 14132 7 1 2 60532 70810
0 14133 5 1 1 14132
0 14134 7 1 2 53464 71485
0 14135 5 1 1 14134
0 14136 7 1 2 14133 14135
0 14137 7 1 2 14131 14136
0 14138 5 1 1 14137
0 14139 7 1 2 48918 14138
0 14140 5 1 1 14139
0 14141 7 1 2 54592 71020
0 14142 5 1 1 14141
0 14143 7 1 2 50686 9430
0 14144 5 1 1 14143
0 14145 7 1 2 61448 14144
0 14146 7 1 2 14142 14145
0 14147 5 1 1 14146
0 14148 7 1 2 14140 14147
0 14149 5 1 1 14148
0 14150 7 1 2 57215 14149
0 14151 5 1 1 14150
0 14152 7 1 2 63760 71590
0 14153 5 1 1 14152
0 14154 7 2 2 70679 72647
0 14155 5 1 1 72915
0 14156 7 1 2 53465 63761
0 14157 5 1 1 14156
0 14158 7 1 2 14155 14157
0 14159 5 1 1 14158
0 14160 7 2 2 56619 14159
0 14161 5 1 1 72917
0 14162 7 1 2 59027 14161
0 14163 7 1 2 14153 14162
0 14164 5 1 1 14163
0 14165 7 1 2 50175 14164
0 14166 5 1 1 14165
0 14167 7 1 2 60758 70365
0 14168 7 2 2 71055 14167
0 14169 7 1 2 72919 71588
0 14170 5 1 1 14169
0 14171 7 1 2 51878 70366
0 14172 5 3 1 14171
0 14173 7 1 2 54248 72921
0 14174 5 2 1 14173
0 14175 7 1 2 72924 71579
0 14176 5 1 1 14175
0 14177 7 8 2 52945 58889
0 14178 5 2 1 72926
0 14179 7 1 2 63653 72927
0 14180 5 1 1 14179
0 14181 7 1 2 14176 14180
0 14182 7 1 2 14170 14181
0 14183 7 1 2 14166 14182
0 14184 5 1 1 14183
0 14185 7 1 2 48919 14184
0 14186 5 1 1 14185
0 14187 7 1 2 14151 14186
0 14188 7 1 2 14123 14187
0 14189 5 1 1 14188
0 14190 7 1 2 57995 14189
0 14191 5 1 1 14190
0 14192 7 1 2 64146 60589
0 14193 5 1 1 14192
0 14194 7 2 2 71012 71326
0 14195 5 1 1 72936
0 14196 7 1 2 14193 14195
0 14197 5 1 1 14196
0 14198 7 1 2 61497 14197
0 14199 5 1 1 14198
0 14200 7 4 2 48920 50983
0 14201 5 4 1 72938
0 14202 7 3 2 56191 70467
0 14203 5 1 1 72946
0 14204 7 1 2 63568 72947
0 14205 5 1 1 14204
0 14206 7 1 2 72942 14205
0 14207 5 1 1 14206
0 14208 7 1 2 52270 14207
0 14209 5 1 1 14208
0 14210 7 1 2 48921 70680
0 14211 5 1 1 14210
0 14212 7 1 2 14209 14211
0 14213 5 1 1 14212
0 14214 7 1 2 50176 14213
0 14215 5 1 1 14214
0 14216 7 1 2 14199 14215
0 14217 5 1 1 14216
0 14218 7 1 2 57216 14217
0 14219 5 1 1 14218
0 14220 7 2 2 51879 71416
0 14221 7 2 2 56192 63569
0 14222 7 1 2 72949 72951
0 14223 5 1 1 14222
0 14224 7 1 2 72943 14223
0 14225 5 1 1 14224
0 14226 7 1 2 70390 14225
0 14227 5 1 1 14226
0 14228 7 2 2 54593 63570
0 14229 7 1 2 56193 72953
0 14230 7 1 2 70637 14229
0 14231 5 1 1 14230
0 14232 7 3 2 48922 50177
0 14233 7 1 2 59896 72955
0 14234 5 1 1 14233
0 14235 7 1 2 14231 14234
0 14236 7 1 2 14227 14235
0 14237 5 1 1 14236
0 14238 7 1 2 50402 14237
0 14239 5 1 1 14238
0 14240 7 4 2 51880 48923
0 14241 7 2 2 50984 70638
0 14242 7 1 2 72958 72962
0 14243 5 1 1 14242
0 14244 7 5 2 51881 54594
0 14245 7 2 2 58890 72964
0 14246 7 1 2 58817 72969
0 14247 5 2 1 14246
0 14248 7 1 2 72909 72971
0 14249 5 1 1 14248
0 14250 7 1 2 72952 14249
0 14251 5 1 1 14250
0 14252 7 1 2 14243 14251
0 14253 7 1 2 14239 14252
0 14254 7 1 2 14219 14253
0 14255 5 1 1 14254
0 14256 7 1 2 58744 14255
0 14257 5 1 1 14256
0 14258 7 1 2 53466 70777
0 14259 5 1 1 14258
0 14260 7 1 2 63762 71600
0 14261 5 1 1 14260
0 14262 7 1 2 14259 14261
0 14263 5 1 1 14262
0 14264 7 1 2 52271 14263
0 14265 5 1 1 14264
0 14266 7 6 2 51882 52384
0 14267 7 2 2 53165 60533
0 14268 5 3 1 72979
0 14269 7 1 2 72973 72980
0 14270 5 1 1 14269
0 14271 7 1 2 49720 14270
0 14272 5 1 1 14271
0 14273 7 1 2 70681 14272
0 14274 5 1 1 14273
0 14275 7 1 2 14265 14274
0 14276 5 1 1 14275
0 14277 7 1 2 50178 14276
0 14278 5 1 1 14277
0 14279 7 7 2 50687 56194
0 14280 5 1 1 72984
0 14281 7 3 2 51883 53467
0 14282 5 1 1 72991
0 14283 7 1 2 14282 71437
0 14284 5 1 1 14283
0 14285 7 1 2 72985 14284
0 14286 5 1 1 14285
0 14287 7 1 2 14278 14286
0 14288 5 1 1 14287
0 14289 7 1 2 57217 14288
0 14290 5 1 1 14289
0 14291 7 1 2 72918 70835
0 14292 5 1 1 14291
0 14293 7 1 2 54249 61253
0 14294 5 11 1 14293
0 14295 7 1 2 57587 72994
0 14296 5 2 1 14295
0 14297 7 1 2 51884 70734
0 14298 5 2 1 14297
0 14299 7 2 2 65361 73007
0 14300 5 1 1 73009
0 14301 7 1 2 73005 73010
0 14302 5 1 1 14301
0 14303 7 2 2 50985 14302
0 14304 5 2 1 73011
0 14305 7 1 2 56620 71141
0 14306 5 1 1 14305
0 14307 7 1 2 61303 14306
0 14308 5 1 1 14307
0 14309 7 1 2 56195 14308
0 14310 5 1 1 14309
0 14311 7 1 2 70836 71273
0 14312 5 1 1 14311
0 14313 7 1 2 14310 14312
0 14314 7 1 2 73013 14313
0 14315 5 1 1 14314
0 14316 7 1 2 53468 14315
0 14317 5 1 1 14316
0 14318 7 1 2 14292 14317
0 14319 7 1 2 14290 14318
0 14320 5 1 1 14319
0 14321 7 1 2 48924 14320
0 14322 5 1 1 14321
0 14323 7 1 2 14257 14322
0 14324 7 1 2 14191 14323
0 14325 5 1 1 14324
0 14326 7 1 2 55284 14325
0 14327 5 1 1 14326
0 14328 7 1 2 54595 65448
0 14329 5 10 1 14328
0 14330 7 2 2 53077 73015
0 14331 7 2 2 52272 73025
0 14332 5 1 1 73027
0 14333 7 1 2 71561 14332
0 14334 5 1 1 14333
0 14335 7 1 2 52091 14334
0 14336 5 1 1 14335
0 14337 7 2 2 61518 60534
0 14338 5 3 1 73029
0 14339 7 1 2 14336 73031
0 14340 5 1 1 14339
0 14341 7 1 2 51885 14340
0 14342 5 1 1 14341
0 14343 7 1 2 51886 61338
0 14344 5 1 1 14343
0 14345 7 13 2 60759 9864
0 14346 5 1 1 73034
0 14347 7 1 2 50688 73035
0 14348 5 1 1 14347
0 14349 7 1 2 14344 14348
0 14350 5 2 1 14349
0 14351 7 1 2 57588 73047
0 14352 5 1 1 14351
0 14353 7 1 2 61339 70241
0 14354 5 1 1 14353
0 14355 7 1 2 52092 61340
0 14356 5 1 1 14355
0 14357 7 1 2 65233 14356
0 14358 5 1 1 14357
0 14359 7 1 2 70719 14358
0 14360 5 1 1 14359
0 14361 7 1 2 14354 14360
0 14362 7 1 2 14352 14361
0 14363 7 1 2 14342 14362
0 14364 5 1 1 14363
0 14365 7 1 2 54964 14364
0 14366 5 1 1 14365
0 14367 7 1 2 63506 70463
0 14368 5 2 1 14367
0 14369 7 1 2 14366 73049
0 14370 5 1 1 14369
0 14371 7 1 2 63486 14370
0 14372 5 1 1 14371
0 14373 7 1 2 14327 14372
0 14374 5 1 1 14373
0 14375 7 1 2 72900 14374
0 14376 5 1 1 14375
0 14377 7 4 2 68241 69649
0 14378 7 3 2 55859 63720
0 14379 5 3 1 73055
0 14380 7 1 2 55285 71501
0 14381 5 1 1 14380
0 14382 7 1 2 73058 14381
0 14383 5 1 1 14382
0 14384 7 1 2 73016 14383
0 14385 5 1 1 14384
0 14386 7 3 2 55286 70955
0 14387 7 1 2 55860 73061
0 14388 5 1 1 14387
0 14389 7 1 2 63747 14388
0 14390 5 1 1 14389
0 14391 7 1 2 65766 14390
0 14392 5 1 1 14391
0 14393 7 1 2 14385 14392
0 14394 5 1 1 14393
0 14395 7 1 2 52093 14394
0 14396 5 1 1 14395
0 14397 7 1 2 54965 73032
0 14398 5 5 1 14397
0 14399 7 2 2 67751 73064
0 14400 7 1 2 51267 73069
0 14401 5 2 1 14400
0 14402 7 2 2 55861 73065
0 14403 5 1 1 73073
0 14404 7 9 2 50179 63638
0 14405 5 2 1 73075
0 14406 7 1 2 14403 73084
0 14407 5 2 1 14406
0 14408 7 1 2 73086 73062
0 14409 5 1 1 14408
0 14410 7 1 2 73071 14409
0 14411 7 1 2 14396 14410
0 14412 5 1 1 14411
0 14413 7 1 2 51887 14412
0 14414 5 1 1 14413
0 14415 7 6 2 55287 55862
0 14416 7 1 2 73088 70166
0 14417 5 2 1 14416
0 14418 7 4 2 50986 70410
0 14419 5 1 1 73096
0 14420 7 2 2 49721 14419
0 14421 5 2 1 73100
0 14422 7 1 2 48730 73101
0 14423 5 2 1 14422
0 14424 7 1 2 73089 73104
0 14425 5 1 1 14424
0 14426 7 1 2 63748 14425
0 14427 5 1 1 14426
0 14428 7 1 2 61341 14427
0 14429 5 1 1 14428
0 14430 7 1 2 73094 14429
0 14431 5 1 1 14430
0 14432 7 1 2 70242 14431
0 14433 5 1 1 14432
0 14434 7 2 2 65337 68381
0 14435 7 1 2 52094 70956
0 14436 5 1 1 14435
0 14437 7 1 2 61342 72765
0 14438 5 1 1 14437
0 14439 7 1 2 14436 14438
0 14440 5 1 1 14439
0 14441 7 1 2 73106 14440
0 14442 5 1 1 14441
0 14443 7 1 2 14433 14442
0 14444 7 1 2 14414 14443
0 14445 5 1 1 14444
0 14446 7 1 2 52787 14445
0 14447 5 1 1 14446
0 14448 7 6 2 50403 55288
0 14449 7 1 2 57218 72736
0 14450 5 2 1 14449
0 14451 7 2 2 62957 72790
0 14452 5 1 1 73116
0 14453 7 1 2 73114 14452
0 14454 5 1 1 14453
0 14455 7 1 2 73108 14454
0 14456 5 1 1 14455
0 14457 7 6 2 51888 51268
0 14458 5 2 1 73118
0 14459 7 1 2 54966 73119
0 14460 5 1 1 14459
0 14461 7 1 2 14456 14460
0 14462 5 1 1 14461
0 14463 7 1 2 61343 14462
0 14464 5 1 1 14463
0 14465 7 1 2 68382 70957
0 14466 5 1 1 14465
0 14467 7 5 2 50689 63721
0 14468 5 2 1 73126
0 14469 7 1 2 52095 73127
0 14470 5 1 1 14469
0 14471 7 1 2 14466 14470
0 14472 5 1 1 14471
0 14473 7 1 2 70243 14472
0 14474 5 1 1 14473
0 14475 7 4 2 63594 70144
0 14476 7 3 2 53273 73133
0 14477 5 1 1 73137
0 14478 7 1 2 73138 72791
0 14479 5 1 1 14478
0 14480 7 1 2 63722 71148
0 14481 5 2 1 14480
0 14482 7 1 2 14479 73140
0 14483 5 1 1 14482
0 14484 7 1 2 50404 14483
0 14485 5 1 1 14484
0 14486 7 1 2 14474 14485
0 14487 7 1 2 14464 14486
0 14488 5 1 1 14487
0 14489 7 1 2 52788 14488
0 14490 5 1 1 14489
0 14491 7 2 2 66600 70340
0 14492 7 1 2 60117 73017
0 14493 7 1 2 73142 14492
0 14494 5 1 1 14493
0 14495 7 1 2 14490 14494
0 14496 5 1 1 14495
0 14497 7 1 2 57589 14496
0 14498 5 1 1 14497
0 14499 7 1 2 61592 68660
0 14500 5 1 1 14499
0 14501 7 1 2 5308 14500
0 14502 5 1 1 14501
0 14503 7 1 2 52273 14502
0 14504 5 1 1 14503
0 14505 7 1 2 53078 72169
0 14506 5 1 1 14505
0 14507 7 1 2 68671 14506
0 14508 5 1 1 14507
0 14509 7 1 2 50690 14508
0 14510 5 1 1 14509
0 14511 7 1 2 14504 14510
0 14512 5 1 1 14511
0 14513 7 1 2 52604 14512
0 14514 5 1 1 14513
0 14515 7 2 2 55863 69792
0 14516 5 2 1 73144
0 14517 7 1 2 63749 73146
0 14518 5 2 1 14517
0 14519 7 2 2 52096 73148
0 14520 5 1 1 73150
0 14521 7 1 2 63800 14520
0 14522 5 1 1 14521
0 14523 7 1 2 52789 14522
0 14524 5 1 1 14523
0 14525 7 1 2 14514 14524
0 14526 5 1 1 14525
0 14527 7 1 2 61344 14526
0 14528 5 1 1 14527
0 14529 7 6 2 49722 66274
0 14530 5 1 1 73152
0 14531 7 1 2 70167 73153
0 14532 5 1 1 14531
0 14533 7 6 2 52097 52790
0 14534 7 1 2 73063 73158
0 14535 5 1 1 14534
0 14536 7 1 2 14532 14535
0 14537 5 1 1 14536
0 14538 7 1 2 59914 14537
0 14539 5 1 1 14538
0 14540 7 3 2 52098 70145
0 14541 7 2 2 55289 60512
0 14542 7 1 2 73164 73167
0 14543 5 1 1 14542
0 14544 7 1 2 73131 14543
0 14545 5 1 1 14544
0 14546 7 1 2 55864 14545
0 14547 5 1 1 14546
0 14548 7 2 2 50691 70146
0 14549 5 1 1 73169
0 14550 7 1 2 73168 73170
0 14551 5 1 1 14550
0 14552 7 1 2 14547 14551
0 14553 5 1 1 14552
0 14554 7 1 2 52791 14553
0 14555 5 1 1 14554
0 14556 7 1 2 14539 14555
0 14557 7 1 2 14528 14556
0 14558 5 1 1 14557
0 14559 7 1 2 70720 14558
0 14560 5 1 1 14559
0 14561 7 1 2 60617 13437
0 14562 5 1 1 14561
0 14563 7 1 2 50405 14562
0 14564 5 1 1 14563
0 14565 7 1 2 61519 70411
0 14566 5 5 1 14565
0 14567 7 1 2 14564 73171
0 14568 5 1 1 14567
0 14569 7 1 2 73143 14568
0 14570 5 1 1 14569
0 14571 7 1 2 14560 14570
0 14572 7 1 2 14498 14571
0 14573 7 1 2 14447 14572
0 14574 5 1 1 14573
0 14575 7 1 2 53673 14574
0 14576 5 1 1 14575
0 14577 7 1 2 60633 73008
0 14578 5 2 1 14577
0 14579 7 1 2 52946 73176
0 14580 5 1 1 14579
0 14581 7 1 2 59766 14580
0 14582 5 1 1 14581
0 14583 7 1 2 50692 14582
0 14584 5 2 1 14583
0 14585 7 3 2 50693 70244
0 14586 5 2 1 73180
0 14587 7 1 2 51889 73026
0 14588 5 1 1 14587
0 14589 7 1 2 73183 14588
0 14590 5 1 1 14589
0 14591 7 1 2 52274 14590
0 14592 5 2 1 14591
0 14593 7 3 2 51890 60193
0 14594 5 1 1 73187
0 14595 7 1 2 70264 14594
0 14596 5 1 1 14595
0 14597 7 1 2 50694 14596
0 14598 5 1 1 14597
0 14599 7 1 2 73185 14598
0 14600 5 1 1 14599
0 14601 7 1 2 52099 14600
0 14602 5 1 1 14601
0 14603 7 1 2 73178 14602
0 14604 5 1 1 14603
0 14605 7 1 2 54967 14604
0 14606 5 1 1 14605
0 14607 7 1 2 73050 14606
0 14608 5 1 1 14607
0 14609 7 1 2 14608 70125
0 14610 5 1 1 14609
0 14611 7 3 2 52100 70721
0 14612 5 1 1 73190
0 14613 7 2 2 70233 14612
0 14614 5 2 1 73193
0 14615 7 1 2 59807 73194
0 14616 5 1 1 14615
0 14617 7 11 2 53274 54968
0 14618 5 2 1 73197
0 14619 7 1 2 73198 71185
0 14620 7 1 2 14616 14619
0 14621 5 1 1 14620
0 14622 7 1 2 14610 14621
0 14623 5 1 1 14622
0 14624 7 1 2 51269 14623
0 14625 5 1 1 14624
0 14626 7 3 2 50695 56443
0 14627 5 1 1 73210
0 14628 7 3 2 56196 73211
0 14629 5 1 1 73213
0 14630 7 3 2 68383 73214
0 14631 7 2 2 57219 61451
0 14632 7 1 2 50406 73219
0 14633 5 1 1 14632
0 14634 7 1 2 72803 14633
0 14635 5 1 1 14634
0 14636 7 1 2 73216 14635
0 14637 5 1 1 14636
0 14638 7 1 2 14625 14637
0 14639 5 1 1 14638
0 14640 7 1 2 62958 14639
0 14641 5 1 1 14640
0 14642 7 1 2 63723 73048
0 14643 5 1 1 14642
0 14644 7 1 2 61520 71059
0 14645 5 1 1 14644
0 14646 7 6 2 52481 71221
0 14647 5 2 1 73221
0 14648 7 1 2 73227 72738
0 14649 5 1 1 14648
0 14650 7 1 2 52101 14649
0 14651 5 1 1 14650
0 14652 7 4 2 50987 59930
0 14653 5 1 1 73229
0 14654 7 1 2 73230 71149
0 14655 5 1 1 14654
0 14656 7 1 2 14651 14655
0 14657 5 1 1 14656
0 14658 7 1 2 56197 14657
0 14659 5 1 1 14658
0 14660 7 1 2 51891 70837
0 14661 5 1 1 14660
0 14662 7 1 2 54969 14661
0 14663 5 4 1 14662
0 14664 7 1 2 56444 73233
0 14665 5 1 1 14664
0 14666 7 1 2 70671 73115
0 14667 5 1 1 14666
0 14668 7 1 2 57996 14667
0 14669 5 1 1 14668
0 14670 7 1 2 14665 14669
0 14671 7 1 2 14659 14670
0 14672 5 1 1 14671
0 14673 7 1 2 50407 14672
0 14674 5 1 1 14673
0 14675 7 1 2 14645 14674
0 14676 5 1 1 14675
0 14677 7 1 2 55290 14676
0 14678 5 1 1 14677
0 14679 7 1 2 14643 14678
0 14680 5 1 1 14679
0 14681 7 1 2 57590 14680
0 14682 5 1 1 14681
0 14683 7 1 2 14477 73059
0 14684 5 2 1 14683
0 14685 7 1 2 73018 73237
0 14686 5 1 1 14685
0 14687 7 1 2 70126 73090
0 14688 5 2 1 14687
0 14689 7 1 2 63750 73239
0 14690 5 1 1 14689
0 14691 7 1 2 65767 14690
0 14692 5 1 1 14691
0 14693 7 1 2 14686 14692
0 14694 5 1 1 14693
0 14695 7 1 2 52102 14694
0 14696 5 1 1 14695
0 14697 7 2 2 55291 70127
0 14698 7 1 2 73241 73087
0 14699 5 1 1 14698
0 14700 7 1 2 73072 14699
0 14701 7 1 2 14696 14700
0 14702 5 1 1 14701
0 14703 7 1 2 51892 14702
0 14704 5 1 1 14703
0 14705 7 1 2 50696 73238
0 14706 5 1 1 14705
0 14707 7 2 2 51270 61345
0 14708 5 1 1 73243
0 14709 7 13 2 52385 55865
0 14710 5 1 1 73245
0 14711 7 3 2 60519 73246
0 14712 5 1 1 73258
0 14713 7 1 2 14708 14712
0 14714 5 1 1 14713
0 14715 7 1 2 54970 14714
0 14716 5 1 1 14715
0 14717 7 1 2 59915 73242
0 14718 5 1 1 14717
0 14719 7 1 2 14716 14718
0 14720 5 1 1 14719
0 14721 7 1 2 52103 14720
0 14722 5 1 1 14721
0 14723 7 1 2 14706 14722
0 14724 5 1 1 14723
0 14725 7 1 2 70722 14724
0 14726 5 1 1 14725
0 14727 7 1 2 60447 69764
0 14728 5 2 1 14727
0 14729 7 1 2 63751 73261
0 14730 5 1 1 14729
0 14731 7 1 2 61346 14730
0 14732 5 1 1 14731
0 14733 7 1 2 73095 14732
0 14734 5 1 1 14733
0 14735 7 1 2 70245 14734
0 14736 5 1 1 14735
0 14737 7 6 2 52104 52386
0 14738 5 1 1 73263
0 14739 7 1 2 53166 73264
0 14740 5 1 1 14739
0 14741 7 1 2 13591 14740
0 14742 5 1 1 14741
0 14743 7 1 2 57997 14742
0 14744 5 1 1 14743
0 14745 7 3 2 52105 52482
0 14746 7 5 2 53275 73269
0 14747 5 1 1 73272
0 14748 7 1 2 56198 65229
0 14749 5 2 1 14748
0 14750 7 1 2 14747 73277
0 14751 7 1 2 14744 14750
0 14752 5 1 1 14751
0 14753 7 1 2 73107 14752
0 14754 5 1 1 14753
0 14755 7 1 2 14736 14754
0 14756 7 1 2 14726 14755
0 14757 7 1 2 14704 14756
0 14758 7 1 2 14682 14757
0 14759 5 1 1 14758
0 14760 7 1 2 62473 14759
0 14761 5 1 1 14760
0 14762 7 1 2 14641 14761
0 14763 7 1 2 14576 14762
0 14764 5 1 1 14763
0 14765 7 1 2 73051 14764
0 14766 5 1 1 14765
0 14767 7 1 2 14376 14766
0 14768 5 1 1 14767
0 14769 7 1 2 55503 14768
0 14770 5 1 1 14769
0 14771 7 3 2 55866 62959
0 14772 5 1 1 73279
0 14773 7 1 2 55292 14772
0 14774 5 3 1 14773
0 14775 7 1 2 65768 73282
0 14776 5 1 1 14775
0 14777 7 1 2 51271 73028
0 14778 5 1 1 14777
0 14779 7 1 2 14776 14778
0 14780 5 1 1 14779
0 14781 7 1 2 53276 14780
0 14782 5 1 1 14781
0 14783 7 1 2 52792 73019
0 14784 5 1 1 14783
0 14785 7 1 2 14782 14784
0 14786 5 1 1 14785
0 14787 7 1 2 52106 14786
0 14788 5 1 1 14787
0 14789 7 1 2 59759 66722
0 14790 5 2 1 14789
0 14791 7 1 2 73066 73283
0 14792 5 1 1 14791
0 14793 7 1 2 60194 71473
0 14794 5 1 1 14793
0 14795 7 1 2 14792 14794
0 14796 5 1 1 14795
0 14797 7 1 2 53277 14796
0 14798 5 1 1 14797
0 14799 7 1 2 73285 14798
0 14800 7 1 2 14788 14799
0 14801 5 1 1 14800
0 14802 7 1 2 70104 14801
0 14803 5 1 1 14802
0 14804 7 6 2 52275 71583
0 14805 7 3 2 59876 66886
0 14806 7 1 2 73287 73293
0 14807 5 1 1 14806
0 14808 7 3 2 52387 60513
0 14809 5 2 1 73296
0 14810 7 1 2 58731 73299
0 14811 5 1 1 14810
0 14812 7 1 2 73020 73159
0 14813 5 1 1 14812
0 14814 7 1 2 73286 14813
0 14815 5 1 1 14814
0 14816 7 1 2 14811 14815
0 14817 5 1 1 14816
0 14818 7 1 2 14807 14817
0 14819 7 1 2 14803 14818
0 14820 5 1 1 14819
0 14821 7 1 2 49895 14820
0 14822 5 1 1 14821
0 14823 7 8 2 53674 63827
0 14824 5 3 1 73301
0 14825 7 4 2 52107 49723
0 14826 7 1 2 73302 73312
0 14827 7 1 2 73021 14826
0 14828 7 1 2 72820 14827
0 14829 5 1 1 14828
0 14830 7 1 2 14822 14829
0 14831 5 1 1 14830
0 14832 7 1 2 51893 14831
0 14833 5 1 1 14832
0 14834 7 9 2 69650 69565
0 14835 5 3 1 73316
0 14836 7 1 2 67960 70128
0 14837 5 1 1 14836
0 14838 7 1 2 73325 14837
0 14839 5 2 1 14838
0 14840 7 1 2 55293 63698
0 14841 5 2 1 14840
0 14842 7 2 2 52108 73330
0 14843 5 1 1 73332
0 14844 7 1 2 59028 14843
0 14845 5 1 1 14844
0 14846 7 1 2 51894 14845
0 14847 5 1 1 14846
0 14848 7 1 2 53469 60118
0 14849 5 1 1 14848
0 14850 7 1 2 63686 14849
0 14851 5 1 1 14850
0 14852 7 1 2 55867 14851
0 14853 5 1 1 14852
0 14854 7 1 2 14847 14853
0 14855 5 1 1 14854
0 14856 7 1 2 52947 14855
0 14857 5 1 1 14856
0 14858 7 1 2 51272 60264
0 14859 5 1 1 14858
0 14860 7 1 2 52109 71486
0 14861 5 2 1 14860
0 14862 7 1 2 63623 73334
0 14863 5 1 1 14862
0 14864 7 1 2 53470 14863
0 14865 5 1 1 14864
0 14866 7 1 2 14859 14865
0 14867 7 1 2 14857 14866
0 14868 5 1 1 14867
0 14869 7 1 2 73328 14868
0 14870 5 1 1 14869
0 14871 7 4 2 63571 66468
0 14872 5 4 1 73336
0 14873 7 1 2 67845 73340
0 14874 5 4 1 14873
0 14875 7 1 2 73344 70320
0 14876 5 1 1 14875
0 14877 7 2 2 51273 68805
0 14878 7 1 2 52110 73348
0 14879 5 1 1 14878
0 14880 7 1 2 14876 14879
0 14881 5 1 1 14880
0 14882 7 1 2 72821 14881
0 14883 5 1 1 14882
0 14884 7 3 2 50697 67881
0 14885 7 1 2 73259 73350
0 14886 5 1 1 14885
0 14887 7 1 2 14883 14886
0 14888 5 1 1 14887
0 14889 7 1 2 70723 14888
0 14890 5 1 1 14889
0 14891 7 5 2 53079 51274
0 14892 5 1 1 73353
0 14893 7 7 2 52276 73354
0 14894 5 2 1 73358
0 14895 7 1 2 70180 73365
0 14896 5 1 1 14895
0 14897 7 1 2 52111 14896
0 14898 5 1 1 14897
0 14899 7 1 2 66284 14898
0 14900 5 1 1 14899
0 14901 7 1 2 62960 14900
0 14902 5 1 1 14901
0 14903 7 1 2 62474 72766
0 14904 5 1 1 14903
0 14905 7 10 2 52112 51275
0 14906 5 1 1 73367
0 14907 7 1 2 59029 14906
0 14908 5 2 1 14907
0 14909 7 1 2 55868 73377
0 14910 5 1 1 14909
0 14911 7 1 2 66285 14910
0 14912 5 1 1 14911
0 14913 7 1 2 70129 14912
0 14914 5 1 1 14913
0 14915 7 1 2 14904 14914
0 14916 7 1 2 14902 14915
0 14917 5 1 1 14916
0 14918 7 9 2 52948 50988
0 14919 5 2 1 73379
0 14920 7 4 2 50408 73380
0 14921 5 1 1 73390
0 14922 7 1 2 49896 73391
0 14923 7 1 2 14917 14922
0 14924 5 1 1 14923
0 14925 7 1 2 14890 14924
0 14926 7 1 2 14870 14925
0 14927 7 1 2 14833 14926
0 14928 5 1 1 14927
0 14929 7 1 2 51543 14928
0 14930 5 1 1 14929
0 14931 7 3 2 52949 62961
0 14932 5 1 1 73394
0 14933 7 1 2 72741 14932
0 14934 5 2 1 14933
0 14935 7 1 2 66275 73397
0 14936 5 1 1 14935
0 14937 7 1 2 50989 64381
0 14938 5 1 1 14937
0 14939 7 1 2 14936 14938
0 14940 5 1 1 14939
0 14941 7 1 2 49897 14940
0 14942 5 1 1 14941
0 14943 7 3 2 54596 68384
0 14944 7 1 2 68824 73399
0 14945 5 1 1 14944
0 14946 7 1 2 14942 14945
0 14947 5 1 1 14946
0 14948 7 1 2 50409 14947
0 14949 5 1 1 14948
0 14950 7 1 2 70527 68792
0 14951 5 5 1 14950
0 14952 7 2 2 50990 73402
0 14953 7 1 2 61521 73407
0 14954 5 1 1 14953
0 14955 7 1 2 70724 73408
0 14956 5 1 1 14955
0 14957 7 1 2 61522 69309
0 14958 7 1 2 72571 14957
0 14959 5 1 1 14958
0 14960 7 1 2 14956 14959
0 14961 5 1 1 14960
0 14962 7 1 2 52113 14961
0 14963 5 1 1 14962
0 14964 7 1 2 14954 14963
0 14965 7 1 2 14949 14964
0 14966 5 1 1 14965
0 14967 7 1 2 61347 14966
0 14968 5 1 1 14967
0 14969 7 1 2 56199 73222
0 14970 5 1 1 14969
0 14971 7 1 2 66286 14970
0 14972 5 1 1 14971
0 14973 7 1 2 60144 14972
0 14974 5 1 1 14973
0 14975 7 1 2 61043 66276
0 14976 5 1 1 14975
0 14977 7 7 2 52114 53167
0 14978 5 1 1 73409
0 14979 7 3 2 53278 50180
0 14980 7 2 2 70147 73416
0 14981 7 1 2 73410 73419
0 14982 5 1 1 14981
0 14983 7 1 2 14976 14982
0 14984 7 1 2 14974 14983
0 14985 5 1 1 14984
0 14986 7 1 2 62962 14985
0 14987 5 1 1 14986
0 14988 7 1 2 61614 66277
0 14989 7 1 2 72622 14988
0 14990 5 1 1 14989
0 14991 7 1 2 14987 14990
0 14992 5 1 1 14991
0 14993 7 1 2 50991 14992
0 14994 5 1 1 14993
0 14995 7 1 2 72992 72822
0 14996 5 1 1 14995
0 14997 7 2 2 73270 71200
0 14998 7 10 2 53279 50698
0 14999 5 3 1 73423
0 15000 7 1 2 65294 73424
0 15001 7 1 2 73421 15000
0 15002 5 1 1 15001
0 15003 7 1 2 14996 15002
0 15004 5 1 1 15003
0 15005 7 1 2 51276 15004
0 15006 5 1 1 15005
0 15007 7 1 2 14994 15006
0 15008 5 1 1 15007
0 15009 7 1 2 49898 15008
0 15010 5 1 1 15009
0 15011 7 10 2 52950 53471
0 15012 5 2 1 73436
0 15013 7 1 2 72739 73446
0 15014 5 1 1 15013
0 15015 7 1 2 52115 15014
0 15016 5 1 1 15015
0 15017 7 1 2 52951 59134
0 15018 5 2 1 15017
0 15019 7 1 2 49724 73448
0 15020 5 3 1 15019
0 15021 7 1 2 59931 73450
0 15022 5 1 1 15021
0 15023 7 1 2 15016 15022
0 15024 5 1 1 15023
0 15025 7 1 2 50410 15024
0 15026 5 1 1 15025
0 15027 7 1 2 73124 15026
0 15028 5 1 1 15027
0 15029 7 1 2 73329 15028
0 15030 5 1 1 15029
0 15031 7 1 2 72792 73345
0 15032 5 1 1 15031
0 15033 7 3 2 52116 59019
0 15034 5 1 1 73453
0 15035 7 1 2 49193 15034
0 15036 5 1 1 15035
0 15037 7 1 2 49899 73231
0 15038 7 1 2 73378 15037
0 15039 7 1 2 15036 15038
0 15040 5 1 1 15039
0 15041 7 1 2 15032 15040
0 15042 5 1 1 15041
0 15043 7 1 2 72823 15042
0 15044 5 1 1 15043
0 15045 7 1 2 62963 71124
0 15046 5 1 1 15045
0 15047 7 2 2 61523 60119
0 15048 5 3 1 73456
0 15049 7 1 2 59351 73457
0 15050 5 1 1 15049
0 15051 7 1 2 14629 15050
0 15052 5 1 1 15051
0 15053 7 1 2 51277 57220
0 15054 7 1 2 15052 15053
0 15055 5 1 1 15054
0 15056 7 1 2 15046 15055
0 15057 5 1 1 15056
0 15058 7 1 2 49900 15057
0 15059 5 1 1 15058
0 15060 7 1 2 15044 15059
0 15061 5 1 1 15060
0 15062 7 1 2 50411 15061
0 15063 5 1 1 15062
0 15064 7 1 2 15030 15063
0 15065 7 1 2 15010 15064
0 15066 7 1 2 14968 15065
0 15067 5 1 1 15066
0 15068 7 1 2 51544 15067
0 15069 5 1 1 15068
0 15070 7 3 2 73022 72676
0 15071 7 1 2 51895 73461
0 15072 5 1 1 15071
0 15073 7 1 2 63624 15072
0 15074 5 3 1 15073
0 15075 7 3 2 51278 73464
0 15076 7 1 2 50992 70575
0 15077 7 1 2 73467 15076
0 15078 5 1 1 15077
0 15079 7 1 2 15069 15078
0 15080 5 1 1 15079
0 15081 7 1 2 57591 15080
0 15082 5 1 1 15081
0 15083 7 3 2 52605 67882
0 15084 5 1 1 73470
0 15085 7 1 2 50993 73454
0 15086 5 1 1 15085
0 15087 7 1 2 48925 15086
0 15088 5 1 1 15087
0 15089 7 2 2 49901 15088
0 15090 5 1 1 73473
0 15091 7 1 2 73341 15090
0 15092 5 1 1 15091
0 15093 7 1 2 55869 15092
0 15094 5 1 1 15093
0 15095 7 1 2 15084 15094
0 15096 5 1 1 15095
0 15097 7 1 2 70130 15096
0 15098 5 1 1 15097
0 15099 7 4 2 52606 53080
0 15100 7 6 2 52277 73475
0 15101 5 2 1 73479
0 15102 7 1 2 55294 73485
0 15103 5 3 1 15102
0 15104 7 1 2 70131 73487
0 15105 5 1 1 15104
0 15106 7 6 2 52278 52793
0 15107 7 2 2 53081 73490
0 15108 5 1 1 73496
0 15109 7 3 2 52607 51279
0 15110 5 3 1 73498
0 15111 7 1 2 15108 73501
0 15112 7 1 2 15105 15111
0 15113 5 1 1 15112
0 15114 7 1 2 49902 15113
0 15115 5 1 1 15114
0 15116 7 1 2 71268 15115
0 15117 5 1 1 15116
0 15118 7 1 2 73102 15117
0 15119 5 1 1 15118
0 15120 7 1 2 73488 73474
0 15121 5 1 1 15120
0 15122 7 3 2 49725 63828
0 15123 7 1 2 73480 73504
0 15124 5 1 1 15123
0 15125 7 1 2 2074 15124
0 15126 5 1 1 15125
0 15127 7 1 2 53675 15126
0 15128 5 1 1 15127
0 15129 7 1 2 15121 15128
0 15130 7 1 2 15119 15129
0 15131 7 1 2 15098 15130
0 15132 5 1 1 15131
0 15133 7 1 2 51545 15132
0 15134 5 1 1 15133
0 15135 7 2 2 51280 64382
0 15136 7 1 2 73165 73425
0 15137 7 1 2 71086 15136
0 15138 7 1 2 73507 15137
0 15139 5 1 1 15138
0 15140 7 1 2 15134 15139
0 15141 5 1 1 15140
0 15142 7 1 2 70246 15141
0 15143 5 1 1 15142
0 15144 7 1 2 55870 64383
0 15145 5 1 1 15144
0 15146 7 2 2 72578 15145
0 15147 5 2 1 73509
0 15148 7 1 2 51546 59932
0 15149 7 1 2 73511 15148
0 15150 5 1 1 15149
0 15151 7 1 2 63063 66601
0 15152 5 1 1 15151
0 15153 7 1 2 49903 15152
0 15154 7 1 2 15150 15153
0 15155 5 1 1 15154
0 15156 7 6 2 49726 55871
0 15157 7 16 2 50181 54971
0 15158 7 2 2 65980 73519
0 15159 7 1 2 51896 73535
0 15160 7 1 2 73513 15159
0 15161 5 1 1 15160
0 15162 7 1 2 63417 66602
0 15163 5 1 1 15162
0 15164 7 1 2 53676 15163
0 15165 7 1 2 15161 15164
0 15166 5 1 1 15165
0 15167 7 1 2 50412 15166
0 15168 7 1 2 15155 15167
0 15169 5 1 1 15168
0 15170 7 2 2 51547 72572
0 15171 7 1 2 60595 71071
0 15172 7 1 2 73537 15171
0 15173 5 1 1 15172
0 15174 7 1 2 15169 15173
0 15175 5 1 1 15174
0 15176 7 1 2 57221 15175
0 15177 5 1 1 15176
0 15178 7 4 2 49904 62964
0 15179 7 3 2 51548 55872
0 15180 5 1 1 73543
0 15181 7 1 2 73160 73381
0 15182 5 1 1 15181
0 15183 7 1 2 15180 15182
0 15184 5 1 1 15183
0 15185 7 1 2 73539 15184
0 15186 5 1 1 15185
0 15187 7 4 2 52117 73437
0 15188 7 1 2 73546 71144
0 15189 5 1 1 15188
0 15190 7 1 2 15186 15189
0 15191 5 1 1 15190
0 15192 7 1 2 67524 15191
0 15193 5 1 1 15192
0 15194 7 1 2 15177 15193
0 15195 5 1 1 15194
0 15196 7 1 2 50699 15195
0 15197 5 1 1 15196
0 15198 7 6 2 51897 51549
0 15199 7 1 2 49905 73512
0 15200 5 2 1 15199
0 15201 7 1 2 73514 69773
0 15202 5 2 1 15201
0 15203 7 1 2 73556 73558
0 15204 5 1 1 15203
0 15205 7 1 2 73550 15204
0 15206 5 1 1 15205
0 15207 7 7 2 51281 55873
0 15208 7 1 2 63064 73560
0 15209 5 1 1 15208
0 15210 7 1 2 51550 64384
0 15211 5 1 1 15210
0 15212 7 1 2 49906 15211
0 15213 7 1 2 15209 15212
0 15214 5 1 1 15213
0 15215 7 10 2 65416 65464
0 15216 5 1 1 73567
0 15217 7 2 2 48926 73288
0 15218 5 1 1 73577
0 15219 7 1 2 51282 73578
0 15220 5 1 1 15219
0 15221 7 1 2 53677 4802
0 15222 7 1 2 15220 15221
0 15223 5 1 1 15222
0 15224 7 1 2 73568 15223
0 15225 7 1 2 15214 15224
0 15226 5 1 1 15225
0 15227 7 1 2 15206 15226
0 15228 5 1 1 15227
0 15229 7 1 2 50994 15228
0 15230 5 1 1 15229
0 15231 7 2 2 61524 63763
0 15232 5 1 1 73579
0 15233 7 2 2 52118 73580
0 15234 5 2 1 73581
0 15235 7 2 2 49907 55874
0 15236 7 1 2 73538 73585
0 15237 7 1 2 73582 15236
0 15238 5 1 1 15237
0 15239 7 1 2 15230 15238
0 15240 7 1 2 15197 15239
0 15241 5 1 1 15240
0 15242 7 1 2 61348 15241
0 15243 5 1 1 15242
0 15244 7 2 2 55875 72793
0 15245 5 1 1 73587
0 15246 7 1 2 71165 15245
0 15247 5 1 1 15246
0 15248 7 1 2 66723 70573
0 15249 7 1 2 15247 15248
0 15250 5 1 1 15249
0 15251 7 1 2 15243 15250
0 15252 7 1 2 15143 15251
0 15253 7 1 2 15082 15252
0 15254 7 1 2 14930 15253
0 15255 5 1 1 15254
0 15256 7 1 2 68242 15255
0 15257 5 1 1 15256
0 15258 7 1 2 14770 15257
0 15259 5 1 1 15258
0 15260 7 1 2 55636 15259
0 15261 5 1 1 15260
0 15262 7 2 2 50995 73462
0 15263 5 1 1 73589
0 15264 7 1 2 49727 15263
0 15265 5 1 1 15264
0 15266 7 1 2 48927 15265
0 15267 5 1 1 15266
0 15268 7 1 2 63478 15267
0 15269 5 1 1 15268
0 15270 7 1 2 51898 15269
0 15271 5 1 1 15270
0 15272 7 4 2 48928 50700
0 15273 5 2 1 73591
0 15274 7 1 2 59877 73592
0 15275 5 1 1 15274
0 15276 7 1 2 15271 15275
0 15277 5 1 1 15276
0 15278 7 1 2 72901 15277
0 15279 5 1 1 15278
0 15280 7 1 2 51899 70009
0 15281 5 1 1 15280
0 15282 7 1 2 50996 70557
0 15283 7 1 2 73465 15282
0 15284 5 1 1 15283
0 15285 7 1 2 15281 15284
0 15286 5 1 1 15285
0 15287 7 1 2 68243 15286
0 15288 5 1 1 15287
0 15289 7 1 2 15279 15288
0 15290 5 1 1 15289
0 15291 7 1 2 55295 15290
0 15292 5 1 1 15291
0 15293 7 1 2 61437 68479
0 15294 5 1 1 15293
0 15295 7 3 2 61958 70725
0 15296 7 1 2 62965 70309
0 15297 7 1 2 73597 15296
0 15298 5 1 1 15297
0 15299 7 1 2 15294 15298
0 15300 5 1 1 15299
0 15301 7 1 2 50997 69206
0 15302 7 1 2 15300 15301
0 15303 5 1 1 15302
0 15304 7 1 2 15292 15303
0 15305 5 1 1 15304
0 15306 7 1 2 55504 15305
0 15307 5 1 1 15306
0 15308 7 1 2 70528 73342
0 15309 5 4 1 15308
0 15310 7 2 2 57222 60535
0 15311 5 3 1 73604
0 15312 7 1 2 73172 73606
0 15313 5 1 1 15312
0 15314 7 1 2 73600 15313
0 15315 5 1 1 15314
0 15316 7 1 2 67883 73117
0 15317 5 1 1 15316
0 15318 7 3 2 59933 66603
0 15319 7 1 2 49908 73609
0 15320 7 1 2 71493 15319
0 15321 5 1 1 15320
0 15322 7 1 2 15317 15321
0 15323 5 1 1 15322
0 15324 7 1 2 50413 15323
0 15325 5 1 1 15324
0 15326 7 1 2 15315 15325
0 15327 5 1 1 15326
0 15328 7 1 2 51551 15327
0 15329 5 1 1 15328
0 15330 7 1 2 66711 70569
0 15331 5 1 1 15330
0 15332 7 1 2 15329 15331
0 15333 5 1 1 15332
0 15334 7 1 2 68244 15333
0 15335 5 1 1 15334
0 15336 7 1 2 15307 15335
0 15337 5 1 1 15336
0 15338 7 1 2 55637 15337
0 15339 5 1 1 15338
0 15340 7 4 2 51900 49728
0 15341 7 2 2 73612 71635
0 15342 7 1 2 67934 69478
0 15343 7 1 2 73616 15342
0 15344 5 1 1 15343
0 15345 7 1 2 15339 15344
0 15346 5 1 1 15345
0 15347 7 1 2 57998 15346
0 15348 5 1 1 15347
0 15349 7 1 2 50035 73610
0 15350 7 1 2 70584 15349
0 15351 5 1 1 15350
0 15352 7 1 2 64704 66415
0 15353 7 1 2 72185 15352
0 15354 5 1 1 15353
0 15355 7 1 2 15351 15354
0 15356 5 1 1 15355
0 15357 7 1 2 50414 15356
0 15358 5 1 1 15357
0 15359 7 2 2 51901 68806
0 15360 7 1 2 69414 73618
0 15361 5 1 1 15360
0 15362 7 1 2 15358 15361
0 15363 5 1 1 15362
0 15364 7 1 2 49037 15363
0 15365 5 1 1 15364
0 15366 7 2 2 50415 67656
0 15367 7 3 2 52866 72301
0 15368 7 1 2 67110 73622
0 15369 7 1 2 73620 15368
0 15370 5 1 1 15369
0 15371 7 1 2 15365 15370
0 15372 5 1 1 15371
0 15373 7 1 2 58745 15372
0 15374 5 1 1 15373
0 15375 7 2 2 49909 71529
0 15376 5 2 1 73625
0 15377 7 2 2 63672 66887
0 15378 5 1 1 73629
0 15379 7 1 2 55505 15378
0 15380 5 1 1 15379
0 15381 7 1 2 73626 15380
0 15382 5 1 1 15381
0 15383 7 5 2 50182 66888
0 15384 5 2 1 73631
0 15385 7 1 2 63418 73632
0 15386 5 1 1 15385
0 15387 7 1 2 60387 72882
0 15388 5 1 1 15387
0 15389 7 1 2 15386 15388
0 15390 5 1 1 15389
0 15391 7 1 2 53678 15390
0 15392 5 1 1 15391
0 15393 7 1 2 15382 15392
0 15394 5 1 1 15393
0 15395 7 1 2 59897 68245
0 15396 7 1 2 15394 15395
0 15397 5 1 1 15396
0 15398 7 1 2 15374 15397
0 15399 5 1 1 15398
0 15400 7 1 2 57223 15399
0 15401 5 1 1 15400
0 15402 7 2 2 65728 69793
0 15403 7 1 2 65338 73638
0 15404 5 1 1 15403
0 15405 7 7 2 49910 69407
0 15406 7 1 2 50183 73640
0 15407 5 1 1 15406
0 15408 7 1 2 15404 15407
0 15409 5 1 1 15408
0 15410 7 1 2 71530 15409
0 15411 5 1 1 15410
0 15412 7 7 2 52608 52794
0 15413 7 6 2 56445 73647
0 15414 7 2 2 52952 55296
0 15415 7 2 2 55506 73660
0 15416 7 1 2 63654 73662
0 15417 7 1 2 73654 15416
0 15418 5 1 1 15417
0 15419 7 1 2 15411 15418
0 15420 5 1 1 15419
0 15421 7 1 2 50036 15420
0 15422 5 1 1 15421
0 15423 7 2 2 71074 69432
0 15424 7 1 2 63673 73664
0 15425 5 1 1 15424
0 15426 7 1 2 68480 72244
0 15427 5 1 1 15426
0 15428 7 1 2 64147 60265
0 15429 7 1 2 72186 15428
0 15430 5 1 1 15429
0 15431 7 1 2 15427 15430
0 15432 5 1 1 15431
0 15433 7 1 2 73663 15432
0 15434 5 1 1 15433
0 15435 7 1 2 15425 15434
0 15436 5 1 1 15435
0 15437 7 1 2 58746 15436
0 15438 5 1 1 15437
0 15439 7 2 2 50416 73438
0 15440 7 1 2 73666 69899
0 15441 5 1 1 15440
0 15442 7 3 2 50037 50184
0 15443 7 1 2 53679 69408
0 15444 7 1 2 73668 15443
0 15445 5 1 1 15444
0 15446 7 1 2 15441 15445
0 15447 5 1 1 15446
0 15448 7 1 2 48929 15447
0 15449 5 1 1 15448
0 15450 7 1 2 15438 15449
0 15451 7 1 2 15422 15450
0 15452 5 1 1 15451
0 15453 7 1 2 49038 15452
0 15454 5 1 1 15453
0 15455 7 2 2 50185 58747
0 15456 5 1 1 73671
0 15457 7 8 2 52119 54972
0 15458 7 2 2 63404 73673
0 15459 7 1 2 73672 73681
0 15460 5 1 1 15459
0 15461 7 1 2 48930 63655
0 15462 5 1 1 15461
0 15463 7 1 2 15460 15462
0 15464 5 1 1 15463
0 15465 7 2 2 55507 73623
0 15466 7 1 2 73661 73683
0 15467 7 1 2 15464 15466
0 15468 5 1 1 15467
0 15469 7 1 2 15454 15468
0 15470 7 1 2 15401 15469
0 15471 5 1 1 15470
0 15472 7 1 2 50701 15471
0 15473 5 1 1 15472
0 15474 7 2 2 55508 72794
0 15475 7 2 2 69566 71525
0 15476 5 1 1 73687
0 15477 7 1 2 73688 71542
0 15478 5 1 1 15477
0 15479 7 1 2 73052 15478
0 15480 5 1 1 15479
0 15481 7 1 2 68280 69616
0 15482 5 1 1 15481
0 15483 7 1 2 15480 15482
0 15484 5 1 1 15483
0 15485 7 2 2 68872 15484
0 15486 7 1 2 73685 73689
0 15487 5 1 1 15486
0 15488 7 1 2 49039 71456
0 15489 7 1 2 73665 15488
0 15490 7 1 2 73191 15489
0 15491 5 1 1 15490
0 15492 7 1 2 15487 15491
0 15493 5 1 1 15492
0 15494 7 1 2 51283 15493
0 15495 5 1 1 15494
0 15496 7 1 2 73076 73547
0 15497 5 1 1 15496
0 15498 7 1 2 48931 15497
0 15499 5 1 1 15498
0 15500 7 1 2 49911 15499
0 15501 5 1 1 15500
0 15502 7 1 2 73343 15501
0 15503 5 1 1 15502
0 15504 7 1 2 58748 15503
0 15505 5 1 1 15504
0 15506 7 1 2 53680 64608
0 15507 5 1 1 15506
0 15508 7 3 2 60795 73382
0 15509 5 1 1 73691
0 15510 7 1 2 15507 73692
0 15511 5 1 1 15510
0 15512 7 1 2 49729 15511
0 15513 5 1 1 15512
0 15514 7 2 2 67137 73627
0 15515 5 4 1 73694
0 15516 7 1 2 68837 73695
0 15517 5 1 1 15516
0 15518 7 1 2 15513 15517
0 15519 5 1 1 15518
0 15520 7 1 2 15505 15519
0 15521 5 1 1 15520
0 15522 7 1 2 68246 73551
0 15523 7 1 2 15521 15522
0 15524 5 1 1 15523
0 15525 7 1 2 15495 15524
0 15526 7 1 2 15473 15525
0 15527 5 1 1 15526
0 15528 7 1 2 55638 15527
0 15529 5 1 1 15528
0 15530 7 2 2 68770 69302
0 15531 5 1 1 73700
0 15532 7 8 2 68247 73701
0 15533 7 1 2 73702 72607
0 15534 5 1 1 15533
0 15535 7 8 2 69651 15476
0 15536 5 1 1 73710
0 15537 7 1 2 68248 15536
0 15538 5 1 1 15537
0 15539 7 2 2 72216 15538
0 15540 7 1 2 53472 73718
0 15541 5 1 1 15540
0 15542 7 1 2 58749 72246
0 15543 5 1 1 15542
0 15544 7 1 2 15541 15543
0 15545 5 1 1 15544
0 15546 7 2 2 55509 15545
0 15547 5 1 1 73720
0 15548 7 1 2 55297 70412
0 15549 7 1 2 73721 15548
0 15550 5 1 1 15549
0 15551 7 4 2 51284 71457
0 15552 7 7 2 51552 71075
0 15553 5 1 1 73726
0 15554 7 1 2 68249 73727
0 15555 7 1 2 73722 15554
0 15556 5 1 1 15555
0 15557 7 1 2 15550 15556
0 15558 5 1 1 15557
0 15559 7 1 2 55639 15558
0 15560 5 1 1 15559
0 15561 7 1 2 70413 73703
0 15562 5 1 1 15561
0 15563 7 1 2 15560 15562
0 15564 5 1 1 15563
0 15565 7 1 2 70247 15564
0 15566 5 1 1 15565
0 15567 7 1 2 15534 15566
0 15568 7 1 2 15529 15567
0 15569 7 1 2 15348 15568
0 15570 5 1 1 15569
0 15571 7 1 2 57592 15570
0 15572 5 1 1 15571
0 15573 7 2 2 51902 62475
0 15574 5 1 1 73733
0 15575 7 6 2 56446 73734
0 15576 5 4 1 73735
0 15577 7 6 2 50417 63779
0 15578 5 2 1 73745
0 15579 7 1 2 73736 73746
0 15580 5 1 1 15579
0 15581 7 2 2 51903 60536
0 15582 5 4 1 73753
0 15583 7 1 2 56548 73755
0 15584 5 1 1 15583
0 15585 7 2 2 57999 15584
0 15586 5 1 1 73759
0 15587 7 1 2 62552 15586
0 15588 5 1 1 15587
0 15589 7 1 2 63724 73280
0 15590 7 1 2 15588 15589
0 15591 5 1 1 15590
0 15592 7 1 2 15580 15591
0 15593 5 1 1 15592
0 15594 7 1 2 69652 15593
0 15595 5 1 1 15594
0 15596 7 4 2 51904 56447
0 15597 5 2 1 73761
0 15598 7 1 2 73747 73762
0 15599 5 1 1 15598
0 15600 7 1 2 73060 15599
0 15601 5 1 1 15600
0 15602 7 1 2 69522 15601
0 15603 5 1 1 15602
0 15604 7 1 2 15595 15603
0 15605 5 1 1 15604
0 15606 7 1 2 68250 15605
0 15607 5 1 1 15606
0 15608 7 7 2 54973 58000
0 15609 7 2 2 52609 73767
0 15610 5 1 1 73774
0 15611 7 1 2 66375 73775
0 15612 5 1 1 15611
0 15613 7 3 2 48932 58750
0 15614 7 1 2 70291 73776
0 15615 5 1 1 15614
0 15616 7 1 2 55298 15615
0 15617 7 1 2 15612 15616
0 15618 5 1 1 15617
0 15619 7 4 2 52279 54974
0 15620 7 2 2 71261 73779
0 15621 5 1 1 73783
0 15622 7 1 2 51285 15621
0 15623 5 1 1 15622
0 15624 7 1 2 72902 15623
0 15625 7 1 2 15618 15624
0 15626 5 1 1 15625
0 15627 7 1 2 15607 15626
0 15628 5 1 1 15627
0 15629 7 1 2 55510 15628
0 15630 5 1 1 15629
0 15631 7 1 2 73601 73760
0 15632 5 1 1 15631
0 15633 7 1 2 61297 73351
0 15634 7 1 2 73763 15633
0 15635 5 1 1 15634
0 15636 7 1 2 52610 73346
0 15637 5 1 1 15636
0 15638 7 1 2 15637 9581
0 15639 7 1 2 15635 15638
0 15640 7 1 2 15632 15639
0 15641 5 1 1 15640
0 15642 7 1 2 72592 15641
0 15643 5 1 1 15642
0 15644 7 1 2 57924 73756
0 15645 5 2 1 15644
0 15646 7 1 2 69479 72181
0 15647 7 1 2 71710 15646
0 15648 7 1 2 73785 15647
0 15649 5 1 1 15648
0 15650 7 1 2 15643 15649
0 15651 7 1 2 15630 15650
0 15652 5 1 1 15651
0 15653 7 1 2 55640 15652
0 15654 5 1 1 15653
0 15655 7 2 2 65729 68661
0 15656 5 1 1 73787
0 15657 7 2 2 67774 73359
0 15658 5 3 1 73789
0 15659 7 1 2 15656 73791
0 15660 5 1 1 15659
0 15661 7 3 2 62966 15660
0 15662 7 1 2 55641 73794
0 15663 5 1 1 15662
0 15664 7 1 2 15531 15663
0 15665 5 1 1 15664
0 15666 7 1 2 50038 15665
0 15667 5 1 1 15666
0 15668 7 4 2 48933 69942
0 15669 5 1 1 73797
0 15670 7 1 2 55642 73798
0 15671 7 1 2 68372 15670
0 15672 5 1 1 15671
0 15673 7 1 2 15667 15672
0 15674 5 1 1 15673
0 15675 7 1 2 49040 73786
0 15676 7 1 2 15674 15675
0 15677 5 1 1 15676
0 15678 7 1 2 15654 15677
0 15679 5 1 1 15678
0 15680 7 1 2 50186 15679
0 15681 5 1 1 15680
0 15682 7 4 2 51905 58751
0 15683 5 2 1 73801
0 15684 7 2 2 64148 73515
0 15685 5 1 1 73807
0 15686 7 1 2 73802 73808
0 15687 5 1 1 15686
0 15688 7 1 2 67729 71327
0 15689 5 1 1 15688
0 15690 7 1 2 15687 15689
0 15691 5 1 1 15690
0 15692 7 3 2 66416 72903
0 15693 7 1 2 15691 73809
0 15694 5 1 1 15693
0 15695 7 2 2 52611 51553
0 15696 5 1 1 73812
0 15697 7 1 2 52795 73360
0 15698 5 1 1 15697
0 15699 7 1 2 15696 15698
0 15700 5 1 1 15699
0 15701 7 1 2 61215 15700
0 15702 5 1 1 15701
0 15703 7 2 2 55876 69908
0 15704 7 1 2 58001 73814
0 15705 5 1 1 15704
0 15706 7 13 2 53280 53473
0 15707 5 1 1 73816
0 15708 7 3 2 52483 73817
0 15709 5 1 1 73829
0 15710 7 1 2 48934 15709
0 15711 5 2 1 15710
0 15712 7 1 2 52612 73361
0 15713 5 1 1 15712
0 15714 7 1 2 55511 15713
0 15715 5 1 1 15714
0 15716 7 1 2 73832 15715
0 15717 5 1 1 15716
0 15718 7 1 2 15705 15717
0 15719 7 1 2 15702 15718
0 15720 5 1 1 15719
0 15721 7 1 2 49912 15720
0 15722 5 1 1 15721
0 15723 7 2 2 55512 58002
0 15724 7 8 2 55299 62476
0 15725 7 1 2 52796 73836
0 15726 7 1 2 73834 15725
0 15727 5 1 1 15726
0 15728 7 1 2 53474 73561
0 15729 5 1 1 15728
0 15730 7 1 2 55513 15729
0 15731 5 1 1 15730
0 15732 7 1 2 48935 15731
0 15733 5 1 1 15732
0 15734 7 1 2 55300 67974
0 15735 5 1 1 15734
0 15736 7 2 2 70325 73362
0 15737 5 1 1 73844
0 15738 7 1 2 15735 15737
0 15739 7 1 2 15733 15738
0 15740 5 1 1 15739
0 15741 7 1 2 53681 72193
0 15742 7 1 2 15740 15741
0 15743 5 1 1 15742
0 15744 7 1 2 15727 15743
0 15745 7 1 2 15722 15744
0 15746 5 1 1 15745
0 15747 7 1 2 63639 68251
0 15748 7 1 2 15746 15747
0 15749 5 1 1 15748
0 15750 7 1 2 15694 15749
0 15751 5 1 1 15750
0 15752 7 1 2 69218 15751
0 15753 5 1 1 15752
0 15754 7 1 2 15681 15753
0 15755 5 1 1 15754
0 15756 7 1 2 57224 15755
0 15757 5 1 1 15756
0 15758 7 1 2 66376 68886
0 15759 7 1 2 70997 15758
0 15760 5 1 1 15759
0 15761 7 1 2 72944 15760
0 15762 5 1 1 15761
0 15763 7 1 2 51906 15762
0 15764 5 1 1 15763
0 15765 7 2 2 63171 68918
0 15766 7 1 2 73516 73846
0 15767 5 1 1 15766
0 15768 7 1 2 15764 15767
0 15769 5 1 1 15768
0 15770 7 1 2 58752 15769
0 15771 5 1 1 15770
0 15772 7 1 2 59352 72959
0 15773 5 1 1 15772
0 15774 7 1 2 15771 15773
0 15775 5 1 1 15774
0 15776 7 1 2 55301 15775
0 15777 5 1 1 15776
0 15778 7 3 2 51286 72995
0 15779 7 1 2 73848 73784
0 15780 5 1 1 15779
0 15781 7 1 2 15777 15780
0 15782 5 1 1 15781
0 15783 7 3 2 55514 72904
0 15784 7 1 2 15782 73851
0 15785 5 1 1 15784
0 15786 7 1 2 68385 73737
0 15787 5 1 1 15786
0 15788 7 2 2 54975 72996
0 15789 7 1 2 73562 73854
0 15790 7 1 2 72706 15789
0 15791 5 1 1 15790
0 15792 7 1 2 15787 15791
0 15793 5 1 1 15792
0 15794 7 1 2 72405 15793
0 15795 5 1 1 15794
0 15796 7 6 2 52484 50187
0 15797 7 2 2 73426 73856
0 15798 5 1 1 73862
0 15799 7 1 2 66893 15798
0 15800 5 2 1 15799
0 15801 7 1 2 51554 73864
0 15802 5 1 1 15801
0 15803 7 2 2 50188 66278
0 15804 7 1 2 52797 73866
0 15805 5 1 1 15804
0 15806 7 4 2 50418 56448
0 15807 5 1 1 73868
0 15808 7 1 2 51555 73869
0 15809 5 1 1 15808
0 15810 7 1 2 15805 15809
0 15811 5 1 1 15810
0 15812 7 1 2 55877 15811
0 15813 5 1 1 15812
0 15814 7 1 2 15802 15813
0 15815 5 1 1 15814
0 15816 7 1 2 56621 15815
0 15817 5 1 1 15816
0 15818 7 1 2 73857 71063
0 15819 5 1 1 15818
0 15820 7 1 2 55302 15819
0 15821 5 1 1 15820
0 15822 7 1 2 55878 15821
0 15823 5 1 1 15822
0 15824 7 1 2 73636 15823
0 15825 5 2 1 15824
0 15826 7 1 2 73552 73872
0 15827 5 1 1 15826
0 15828 7 1 2 15817 15827
0 15829 5 1 1 15828
0 15830 7 1 2 50998 15829
0 15831 5 1 1 15830
0 15832 7 1 2 72997 72191
0 15833 5 1 1 15832
0 15834 7 1 2 15831 15833
0 15835 5 1 1 15834
0 15836 7 1 2 62967 15835
0 15837 5 1 1 15836
0 15838 7 1 2 61304 63625
0 15839 5 3 1 15838
0 15840 7 2 2 52120 73874
0 15841 5 1 1 73877
0 15842 7 1 2 73383 73878
0 15843 5 1 1 15842
0 15844 7 1 2 56449 56622
0 15845 5 2 1 15844
0 15846 7 1 2 55879 73077
0 15847 5 1 1 15846
0 15848 7 1 2 73879 15847
0 15849 5 1 1 15848
0 15850 7 1 2 51907 15849
0 15851 5 1 1 15850
0 15852 7 1 2 15807 15851
0 15853 7 1 2 15843 15852
0 15854 5 1 1 15853
0 15855 7 1 2 51556 15854
0 15856 5 1 1 15855
0 15857 7 3 2 52280 52485
0 15858 7 2 2 53281 73881
0 15859 5 1 1 73884
0 15860 7 1 2 61598 66633
0 15861 7 1 2 73885 15860
0 15862 5 1 1 15861
0 15863 7 1 2 15856 15862
0 15864 5 1 1 15863
0 15865 7 1 2 64385 15864
0 15866 5 1 1 15865
0 15867 7 1 2 69909 71556
0 15868 7 1 2 14300 15867
0 15869 5 1 1 15868
0 15870 7 1 2 49913 15869
0 15871 7 1 2 15866 15870
0 15872 7 1 2 15837 15871
0 15873 5 1 1 15872
0 15874 7 1 2 73855 71544
0 15875 5 1 1 15874
0 15876 7 3 2 58753 56623
0 15877 5 1 1 73886
0 15878 7 3 2 59878 58801
0 15879 5 1 1 73889
0 15880 7 1 2 73887 73890
0 15881 5 1 1 15880
0 15882 7 1 2 15875 15881
0 15883 5 1 1 15882
0 15884 7 1 2 55515 15883
0 15885 5 1 1 15884
0 15886 7 4 2 48936 52953
0 15887 7 1 2 63605 71174
0 15888 7 2 2 73892 15887
0 15889 5 1 1 73896
0 15890 7 1 2 53475 73897
0 15891 5 1 1 15890
0 15892 7 1 2 15885 15891
0 15893 5 1 1 15892
0 15894 7 1 2 51287 15893
0 15895 5 1 1 15894
0 15896 7 2 2 63507 71670
0 15897 7 1 2 73569 73898
0 15898 5 1 1 15897
0 15899 7 1 2 15895 15898
0 15900 5 1 1 15899
0 15901 7 1 2 55880 15900
0 15902 5 1 1 15901
0 15903 7 1 2 58754 73505
0 15904 5 1 1 15903
0 15905 7 1 2 63428 15904
0 15906 5 1 1 15905
0 15907 7 1 2 72998 15906
0 15908 5 1 1 15907
0 15909 7 1 2 15889 15908
0 15910 5 1 1 15909
0 15911 7 1 2 51557 15910
0 15912 5 1 1 15911
0 15913 7 2 2 64386 1830
0 15914 7 3 2 51908 68386
0 15915 7 1 2 55516 73902
0 15916 7 1 2 73900 15915
0 15917 5 1 1 15916
0 15918 7 1 2 53682 15917
0 15919 7 1 2 15912 15918
0 15920 7 1 2 15902 15919
0 15921 5 1 1 15920
0 15922 7 1 2 15873 15921
0 15923 5 1 1 15922
0 15924 7 1 2 15795 15923
0 15925 5 1 1 15924
0 15926 7 1 2 68252 15925
0 15927 5 1 1 15926
0 15928 7 1 2 15785 15927
0 15929 5 1 1 15928
0 15930 7 1 2 55643 15929
0 15931 5 1 1 15930
0 15932 7 1 2 50039 73795
0 15933 5 1 1 15932
0 15934 7 2 2 63481 66417
0 15935 7 1 2 69943 73905
0 15936 5 1 1 15935
0 15937 7 1 2 15933 15936
0 15938 5 1 1 15937
0 15939 7 1 2 49041 15938
0 15940 5 1 1 15939
0 15941 7 1 2 73624 73906
0 15942 5 1 1 15941
0 15943 7 1 2 15940 15942
0 15944 5 1 1 15943
0 15945 7 1 2 55644 15944
0 15946 5 1 1 15945
0 15947 7 1 2 49730 50040
0 15948 7 1 2 67829 15947
0 15949 7 2 2 72058 15948
0 15950 5 2 1 73907
0 15951 7 1 2 15946 73909
0 15952 5 1 1 15951
0 15953 7 1 2 72999 15952
0 15954 5 1 1 15953
0 15955 7 1 2 70570 73570
0 15956 5 1 1 15955
0 15957 7 1 2 67775 72770
0 15958 5 1 1 15957
0 15959 7 1 2 15956 15958
0 15960 5 1 1 15959
0 15961 7 1 2 51288 15960
0 15962 5 1 1 15961
0 15963 7 1 2 73403 73553
0 15964 5 1 1 15963
0 15965 7 1 2 15962 15964
0 15966 5 1 1 15965
0 15967 7 1 2 68253 15966
0 15968 5 1 1 15967
0 15969 7 1 2 50419 73588
0 15970 5 1 1 15969
0 15971 7 1 2 73173 15970
0 15972 5 1 1 15971
0 15973 7 1 2 7400 9557
0 15974 5 1 1 15973
0 15975 7 1 2 55303 72213
0 15976 7 1 2 15974 15975
0 15977 7 1 2 15972 15976
0 15978 5 1 1 15977
0 15979 7 1 2 52613 68579
0 15980 7 1 2 72107 15979
0 15981 7 1 2 73571 15980
0 15982 5 1 1 15981
0 15983 7 1 2 60596 72024
0 15984 7 5 2 50041 51289
0 15985 7 5 2 53082 54250
0 15986 5 2 1 73916
0 15987 7 1 2 73911 73917
0 15988 7 1 2 15983 15987
0 15989 7 1 2 70058 15988
0 15990 5 1 1 15989
0 15991 7 1 2 15982 15990
0 15992 7 1 2 15978 15991
0 15993 5 1 1 15992
0 15994 7 1 2 55517 15993
0 15995 5 1 1 15994
0 15996 7 1 2 15968 15995
0 15997 5 1 1 15996
0 15998 7 1 2 69978 15997
0 15999 5 1 1 15998
0 16000 7 1 2 15954 15999
0 16001 5 1 1 16000
0 16002 7 1 2 58003 16001
0 16003 5 1 1 16002
0 16004 7 1 2 59898 73704
0 16005 5 1 1 16004
0 16006 7 1 2 73149 73719
0 16007 5 1 1 16006
0 16008 7 3 2 53476 63725
0 16009 5 2 1 73923
0 16010 7 1 2 68662 71321
0 16011 5 1 1 16010
0 16012 7 1 2 73926 16011
0 16013 5 1 1 16012
0 16014 7 1 2 58755 73053
0 16015 7 1 2 16013 16014
0 16016 5 1 1 16015
0 16017 7 1 2 16007 16016
0 16018 5 1 1 16017
0 16019 7 1 2 55518 16018
0 16020 5 1 1 16019
0 16021 7 1 2 73303 73517
0 16022 5 1 1 16021
0 16023 7 1 2 73557 16022
0 16024 5 2 1 16023
0 16025 7 1 2 58004 72593
0 16026 7 1 2 73928 16025
0 16027 5 1 1 16026
0 16028 7 1 2 16020 16027
0 16029 5 1 1 16028
0 16030 7 1 2 55645 16029
0 16031 5 1 1 16030
0 16032 7 1 2 55881 73705
0 16033 5 1 1 16032
0 16034 7 1 2 16031 16033
0 16035 5 1 1 16034
0 16036 7 1 2 73466 16035
0 16037 5 1 1 16036
0 16038 7 1 2 16005 16037
0 16039 7 1 2 16003 16038
0 16040 7 1 2 15931 16039
0 16041 7 1 2 15757 16040
0 16042 7 1 2 15572 16041
0 16043 5 1 1 16042
0 16044 7 1 2 57001 16043
0 16045 5 1 1 16044
0 16046 7 1 2 60624 59307
0 16047 5 1 1 16046
0 16048 7 2 2 63626 16047
0 16049 7 1 2 56624 70735
0 16050 5 1 1 16049
0 16051 7 3 2 50420 63130
0 16052 5 1 1 73932
0 16053 7 1 2 16050 16052
0 16054 5 1 1 16053
0 16055 7 1 2 51909 16054
0 16056 5 1 1 16055
0 16057 7 1 2 73930 16056
0 16058 5 2 1 16057
0 16059 7 1 2 61349 73935
0 16060 5 1 1 16059
0 16061 7 1 2 61350 71487
0 16062 5 1 1 16061
0 16063 7 1 2 54976 70985
0 16064 5 1 1 16063
0 16065 7 1 2 50189 70764
0 16066 7 1 2 16064 16065
0 16067 5 1 1 16066
0 16068 7 1 2 16062 16067
0 16069 5 1 1 16068
0 16070 7 1 2 57225 16069
0 16071 5 1 1 16070
0 16072 7 1 2 73014 16071
0 16073 7 1 2 16060 16072
0 16074 5 1 1 16073
0 16075 7 1 2 73706 16074
0 16076 5 1 1 16075
0 16077 7 1 2 16045 16076
0 16078 7 1 2 15261 16077
0 16079 5 1 1 16078
0 16080 7 1 2 58424 16079
0 16081 5 1 1 16080
0 16082 7 1 2 48731 49042
0 16083 7 2 2 51738 16082
0 16084 7 1 2 61305 73937
0 16085 5 1 1 16084
0 16086 7 1 2 52867 71898
0 16087 7 1 2 68654 16086
0 16088 5 1 1 16087
0 16089 7 1 2 16085 16088
0 16090 5 1 1 16089
0 16091 7 1 2 57152 16090
0 16092 5 1 1 16091
0 16093 7 1 2 59701 73938
0 16094 5 1 1 16093
0 16095 7 1 2 16092 16094
0 16096 5 1 1 16095
0 16097 7 1 2 54597 16096
0 16098 5 1 1 16097
0 16099 7 1 2 48732 72066
0 16100 7 1 2 66771 16099
0 16101 5 1 1 16100
0 16102 7 1 2 16098 16101
0 16103 5 1 1 16102
0 16104 7 1 2 54007 16103
0 16105 5 1 1 16104
0 16106 7 1 2 63996 69086
0 16107 5 1 1 16106
0 16108 7 1 2 72070 16107
0 16109 5 1 1 16108
0 16110 7 1 2 48733 60747
0 16111 7 1 2 16109 16110
0 16112 5 1 1 16111
0 16113 7 1 2 16105 16112
0 16114 5 1 1 16113
0 16115 7 1 2 53892 16114
0 16116 5 1 1 16115
0 16117 7 1 2 61020 69087
0 16118 5 1 1 16117
0 16119 7 1 2 72071 16118
0 16120 5 1 1 16119
0 16121 7 1 2 48351 16120
0 16122 5 1 1 16121
0 16123 7 1 2 49309 72067
0 16124 5 1 1 16123
0 16125 7 1 2 64705 69088
0 16126 5 1 1 16125
0 16127 7 1 2 16124 16126
0 16128 7 1 2 16122 16127
0 16129 5 1 1 16128
0 16130 7 1 2 56709 16129
0 16131 5 1 1 16130
0 16132 7 1 2 54598 72068
0 16133 5 1 1 16132
0 16134 7 2 2 49043 66772
0 16135 7 1 2 69047 73939
0 16136 5 1 1 16135
0 16137 7 1 2 16133 16136
0 16138 7 1 2 16131 16137
0 16139 5 1 1 16138
0 16140 7 1 2 48734 16139
0 16141 5 1 1 16140
0 16142 7 1 2 16116 16141
0 16143 5 1 1 16142
0 16144 7 1 2 55304 16143
0 16145 5 1 1 16144
0 16146 7 2 2 58267 65428
0 16147 5 1 1 73941
0 16148 7 2 2 61549 68033
0 16149 5 1 1 73943
0 16150 7 1 2 73942 16149
0 16151 5 1 1 16150
0 16152 7 1 2 58255 61747
0 16153 5 6 1 16152
0 16154 7 1 2 53083 73945
0 16155 5 2 1 16154
0 16156 7 1 2 48352 73951
0 16157 7 1 2 16151 16156
0 16158 5 1 1 16157
0 16159 7 1 2 64185 16158
0 16160 5 2 1 16159
0 16161 7 1 2 62906 69974
0 16162 7 1 2 73953 16161
0 16163 5 1 1 16162
0 16164 7 1 2 16145 16163
0 16165 5 1 1 16164
0 16166 7 1 2 67830 16165
0 16167 5 1 1 16166
0 16168 7 1 2 49044 58477
0 16169 7 1 2 63354 16168
0 16170 7 1 2 68058 72004
0 16171 7 1 2 16169 16170
0 16172 5 1 1 16171
0 16173 7 1 2 16167 16172
0 16174 5 1 1 16173
0 16175 7 1 2 57925 16174
0 16176 5 1 1 16175
0 16177 7 2 2 59501 61903
0 16178 5 1 1 73955
0 16179 7 1 2 59259 73956
0 16180 7 2 2 62907 69151
0 16181 7 1 2 73957 72015
0 16182 7 1 2 16179 16181
0 16183 5 1 1 16182
0 16184 7 1 2 53789 16183
0 16185 7 1 2 16176 16184
0 16186 5 1 1 16185
0 16187 7 1 2 61645 69089
0 16188 5 1 1 16187
0 16189 7 2 2 49194 62604
0 16190 5 2 1 73959
0 16191 7 1 2 63795 68550
0 16192 7 1 2 73960 16191
0 16193 5 1 1 16192
0 16194 7 1 2 16188 16193
0 16195 5 1 1 16194
0 16196 7 1 2 53893 16195
0 16197 5 1 1 16196
0 16198 7 1 2 54599 69071
0 16199 5 1 1 16198
0 16200 7 1 2 16197 16199
0 16201 5 1 1 16200
0 16202 7 1 2 67183 16201
0 16203 5 1 1 16202
0 16204 7 1 2 69828 16203
0 16205 5 1 1 16204
0 16206 7 1 2 48735 16205
0 16207 5 1 1 16206
0 16208 7 4 2 53894 61550
0 16209 5 1 1 73963
0 16210 7 1 2 73447 73964
0 16211 7 1 2 69515 16210
0 16212 5 1 1 16211
0 16213 7 1 2 63411 16212
0 16214 5 1 1 16213
0 16215 7 1 2 68555 16214
0 16216 5 1 1 16215
0 16217 7 1 2 61551 66082
0 16218 5 1 1 16217
0 16219 7 1 2 16216 16218
0 16220 5 1 1 16219
0 16221 7 1 2 69090 16220
0 16222 5 1 1 16221
0 16223 7 1 2 16207 16222
0 16224 5 1 1 16223
0 16225 7 1 2 57926 16224
0 16226 5 1 1 16225
0 16227 7 1 2 49195 69742
0 16228 5 1 1 16227
0 16229 7 1 2 53477 16228
0 16230 5 1 1 16229
0 16231 7 1 2 48736 16230
0 16232 5 1 1 16231
0 16233 7 3 2 49196 49731
0 16234 7 1 2 69743 73967
0 16235 5 1 1 16234
0 16236 7 1 2 53683 16235
0 16237 7 1 2 16232 16236
0 16238 5 1 1 16237
0 16239 7 1 2 68556 16238
0 16240 5 1 1 16239
0 16241 7 1 2 61748 59135
0 16242 7 1 2 66418 16241
0 16243 5 1 1 16242
0 16244 7 1 2 16240 16243
0 16245 5 1 1 16244
0 16246 7 1 2 54251 16245
0 16247 5 1 1 16246
0 16248 7 1 2 55519 69774
0 16249 5 1 1 16248
0 16250 7 2 2 67288 69440
0 16251 5 1 1 73970
0 16252 7 1 2 66115 16251
0 16253 5 1 1 16252
0 16254 7 1 2 48737 16253
0 16255 5 1 1 16254
0 16256 7 3 2 51558 68991
0 16257 5 1 1 73972
0 16258 7 1 2 63451 73973
0 16259 5 2 1 16258
0 16260 7 1 2 68732 73975
0 16261 7 1 2 16255 16260
0 16262 5 1 1 16261
0 16263 7 1 2 61552 16262
0 16264 5 1 1 16263
0 16265 7 1 2 16249 16264
0 16266 7 1 2 16247 16265
0 16267 5 1 1 16266
0 16268 7 1 2 69091 16267
0 16269 5 1 1 16268
0 16270 7 1 2 16226 16269
0 16271 5 1 1 16270
0 16272 7 1 2 48144 16271
0 16273 5 1 1 16272
0 16274 7 1 2 55305 61672
0 16275 7 1 2 71920 16274
0 16276 5 1 1 16275
0 16277 7 2 2 65429 70248
0 16278 5 1 1 73977
0 16279 7 1 2 16278 71999
0 16280 7 1 2 69455 16279
0 16281 5 1 1 16280
0 16282 7 1 2 16276 16281
0 16283 5 1 1 16282
0 16284 7 1 2 54600 16283
0 16285 5 1 1 16284
0 16286 7 2 2 55520 69895
0 16287 7 1 2 64218 73979
0 16288 7 1 2 58974 16287
0 16289 5 1 1 16288
0 16290 7 1 2 16285 16289
0 16291 5 1 1 16290
0 16292 7 1 2 51739 16291
0 16293 5 1 1 16292
0 16294 7 1 2 16273 16293
0 16295 5 1 1 16294
0 16296 7 1 2 49310 16295
0 16297 5 1 1 16296
0 16298 7 1 2 65244 70859
0 16299 5 1 1 16298
0 16300 7 1 2 50999 16299
0 16301 5 1 1 16300
0 16302 7 1 2 71921 16301
0 16303 5 1 1 16302
0 16304 7 1 2 68039 69180
0 16305 5 1 1 16304
0 16306 7 1 2 16303 16305
0 16307 5 1 1 16306
0 16308 7 1 2 55306 16307
0 16309 5 1 1 16308
0 16310 7 2 2 53895 66083
0 16311 5 1 1 73981
0 16312 7 1 2 64767 72850
0 16313 5 1 1 16312
0 16314 7 1 2 16311 16313
0 16315 5 1 1 16314
0 16316 7 1 2 54601 16315
0 16317 5 1 1 16316
0 16318 7 1 2 61854 68357
0 16319 5 1 1 16318
0 16320 7 1 2 16317 16319
0 16321 5 1 1 16320
0 16322 7 1 2 62553 16321
0 16323 5 1 1 16322
0 16324 7 1 2 53896 71837
0 16325 5 1 1 16324
0 16326 7 1 2 57850 67184
0 16327 7 1 2 68498 16326
0 16328 5 1 1 16327
0 16329 7 1 2 56710 66084
0 16330 7 1 2 66179 16329
0 16331 5 1 1 16330
0 16332 7 1 2 16328 16331
0 16333 5 1 1 16332
0 16334 7 1 2 54008 16333
0 16335 5 1 1 16334
0 16336 7 1 2 64768 66085
0 16337 5 1 1 16336
0 16338 7 1 2 16335 16337
0 16339 5 1 1 16338
0 16340 7 1 2 54252 16339
0 16341 5 1 1 16340
0 16342 7 1 2 16325 16341
0 16343 7 1 2 16323 16342
0 16344 5 1 1 16343
0 16345 7 1 2 49045 16344
0 16346 5 1 1 16345
0 16347 7 1 2 16309 16346
0 16348 5 1 1 16347
0 16349 7 1 2 51740 16348
0 16350 5 1 1 16349
0 16351 7 1 2 16297 16350
0 16352 5 1 1 16351
0 16353 7 1 2 48353 16352
0 16354 5 1 1 16353
0 16355 7 1 2 53897 65685
0 16356 5 1 1 16355
0 16357 7 1 2 51000 16356
0 16358 5 1 1 16357
0 16359 7 1 2 71922 16358
0 16360 5 1 1 16359
0 16361 7 1 2 59709 69181
0 16362 5 1 1 16361
0 16363 7 1 2 16360 16362
0 16364 5 1 1 16363
0 16365 7 1 2 64219 16364
0 16366 5 1 1 16365
0 16367 7 1 2 51001 16178
0 16368 5 2 1 16367
0 16369 7 1 2 60075 73983
0 16370 5 1 1 16369
0 16371 7 4 2 48145 64706
0 16372 5 1 1 73985
0 16373 7 1 2 64424 59527
0 16374 5 1 1 16373
0 16375 7 1 2 16372 16374
0 16376 7 1 2 16370 16375
0 16377 5 1 1 16376
0 16378 7 1 2 71923 16377
0 16379 5 1 1 16378
0 16380 7 1 2 49197 68163
0 16381 5 1 1 16380
0 16382 7 3 2 53898 60388
0 16383 5 2 1 73989
0 16384 7 2 2 50702 73992
0 16385 5 4 1 73994
0 16386 7 1 2 49311 61846
0 16387 5 1 1 16386
0 16388 7 1 2 73995 16387
0 16389 7 1 2 16381 16388
0 16390 5 1 1 16389
0 16391 7 1 2 69182 16390
0 16392 5 1 1 16391
0 16393 7 1 2 16379 16392
0 16394 7 1 2 16366 16393
0 16395 5 1 1 16394
0 16396 7 1 2 55307 16395
0 16397 5 1 1 16396
0 16398 7 1 2 53899 67634
0 16399 5 1 1 16398
0 16400 7 4 2 54009 58478
0 16401 5 2 1 74000
0 16402 7 1 2 58276 74001
0 16403 7 1 2 72028 16402
0 16404 5 1 1 16403
0 16405 7 1 2 16399 16404
0 16406 5 1 1 16405
0 16407 7 1 2 51559 16406
0 16408 5 1 1 16407
0 16409 7 1 2 54602 61698
0 16410 5 1 1 16409
0 16411 7 1 2 60885 61850
0 16412 5 1 1 16411
0 16413 7 1 2 16410 16412
0 16414 5 1 1 16413
0 16415 7 1 2 54253 16414
0 16416 5 1 1 16415
0 16417 7 2 2 53084 61994
0 16418 5 1 1 74006
0 16419 7 1 2 65245 16418
0 16420 5 1 1 16419
0 16421 7 1 2 16416 16420
0 16422 5 1 1 16421
0 16423 7 1 2 66086 16422
0 16424 5 1 1 16423
0 16425 7 1 2 16424 16257
0 16426 5 1 1 16425
0 16427 7 1 2 58975 16426
0 16428 5 1 1 16427
0 16429 7 1 2 16408 16428
0 16430 5 1 1 16429
0 16431 7 1 2 49046 16430
0 16432 5 1 1 16431
0 16433 7 1 2 16397 16432
0 16434 5 1 1 16433
0 16435 7 1 2 51741 16434
0 16436 5 1 1 16435
0 16437 7 1 2 50042 16436
0 16438 7 1 2 16354 16437
0 16439 5 1 1 16438
0 16440 7 1 2 58853 16439
0 16441 7 1 2 16186 16440
0 16442 5 1 1 16441
0 16443 7 1 2 49114 73965
0 16444 5 2 1 16443
0 16445 7 3 2 61771 74008
0 16446 5 5 1 74010
0 16447 7 1 2 47879 74013
0 16448 5 2 1 16447
0 16449 7 1 2 54010 59835
0 16450 5 2 1 16449
0 16451 7 3 2 74018 74020
0 16452 5 1 1 74022
0 16453 7 1 2 48146 16452
0 16454 5 1 1 16453
0 16455 7 1 2 54011 59453
0 16456 5 2 1 16455
0 16457 7 2 2 16454 74025
0 16458 5 2 1 74027
0 16459 7 1 2 69765 69328
0 16460 7 2 2 74029 16459
0 16461 7 1 2 71899 74031
0 16462 5 1 1 16461
0 16463 7 1 2 53684 61021
0 16464 7 1 2 72874 16463
0 16465 5 1 1 16464
0 16466 7 1 2 68908 16465
0 16467 5 1 1 16466
0 16468 7 1 2 48354 16467
0 16469 5 2 1 16468
0 16470 7 2 2 67935 71731
0 16471 5 3 1 74035
0 16472 7 1 2 74033 74037
0 16473 5 3 1 16472
0 16474 7 1 2 59984 74040
0 16475 5 1 1 16474
0 16476 7 2 2 47880 66582
0 16477 7 2 2 68919 68467
0 16478 7 1 2 74043 74045
0 16479 5 1 1 16478
0 16480 7 1 2 16475 16479
0 16481 5 1 1 16480
0 16482 7 1 2 54254 16481
0 16483 5 1 1 16482
0 16484 7 1 2 64657 69376
0 16485 5 1 1 16484
0 16486 7 1 2 69822 16485
0 16487 5 4 1 16486
0 16488 7 1 2 54012 74047
0 16489 5 2 1 16488
0 16490 7 2 2 66247 69333
0 16491 5 2 1 74053
0 16492 7 2 2 59337 69348
0 16493 5 1 1 74057
0 16494 7 1 2 74055 16493
0 16495 5 1 1 16494
0 16496 7 1 2 48355 16495
0 16497 5 1 1 16496
0 16498 7 1 2 74051 16497
0 16499 7 1 2 16483 16498
0 16500 5 1 1 16499
0 16501 7 1 2 48147 16500
0 16502 5 1 1 16501
0 16503 7 1 2 67671 74046
0 16504 5 1 1 16503
0 16505 7 1 2 69823 16504
0 16506 5 1 1 16505
0 16507 7 1 2 56063 16506
0 16508 5 1 1 16507
0 16509 7 1 2 62720 69349
0 16510 5 1 1 16509
0 16511 7 1 2 69385 16510
0 16512 5 1 1 16511
0 16513 7 1 2 57472 16512
0 16514 5 1 1 16513
0 16515 7 1 2 57736 69341
0 16516 5 1 1 16515
0 16517 7 1 2 16514 16516
0 16518 7 1 2 16508 16517
0 16519 7 1 2 16502 16518
0 16520 5 1 1 16519
0 16521 7 1 2 58603 16520
0 16522 5 1 1 16521
0 16523 7 1 2 65836 74041
0 16524 5 1 1 16523
0 16525 7 1 2 65815 69383
0 16526 5 1 1 16525
0 16527 7 1 2 69824 16526
0 16528 5 2 1 16527
0 16529 7 1 2 60294 74059
0 16530 5 1 1 16529
0 16531 7 1 2 69350 71786
0 16532 5 2 1 16531
0 16533 7 1 2 16530 74061
0 16534 7 1 2 16524 16533
0 16535 5 1 1 16534
0 16536 7 1 2 61092 16535
0 16537 5 1 1 16536
0 16538 7 2 2 74038 74056
0 16539 5 2 1 74063
0 16540 7 1 2 48356 74065
0 16541 5 1 1 16540
0 16542 7 1 2 74052 16541
0 16543 5 1 1 16542
0 16544 7 1 2 54255 16543
0 16545 5 1 1 16544
0 16546 7 2 2 67696 69219
0 16547 7 1 2 66761 74067
0 16548 5 2 1 16547
0 16549 7 1 2 60056 68901
0 16550 5 1 1 16549
0 16551 7 1 2 74069 16550
0 16552 5 1 1 16551
0 16553 7 1 2 48357 16552
0 16554 5 1 1 16553
0 16555 7 1 2 58674 69351
0 16556 5 1 1 16555
0 16557 7 3 2 54603 60234
0 16558 5 5 1 74071
0 16559 7 2 2 69334 74074
0 16560 7 2 2 60901 74079
0 16561 5 1 1 74081
0 16562 7 1 2 16556 16561
0 16563 7 1 2 16554 16562
0 16564 5 1 1 16563
0 16565 7 1 2 48148 16564
0 16566 5 1 1 16565
0 16567 7 1 2 16545 16566
0 16568 5 1 1 16567
0 16569 7 1 2 61053 16568
0 16570 5 1 1 16569
0 16571 7 2 2 54604 59674
0 16572 5 4 1 74083
0 16573 7 1 2 60266 74085
0 16574 5 1 1 16573
0 16575 7 1 2 48358 60902
0 16576 7 1 2 69352 16575
0 16577 7 1 2 16574 16576
0 16578 5 1 1 16577
0 16579 7 1 2 60088 66583
0 16580 7 1 2 74068 16579
0 16581 5 1 1 16580
0 16582 7 1 2 69360 16581
0 16583 5 1 1 16582
0 16584 7 1 2 54977 16583
0 16585 5 1 1 16584
0 16586 7 1 2 64433 69377
0 16587 5 1 1 16586
0 16588 7 1 2 69825 16587
0 16589 5 2 1 16588
0 16590 7 1 2 49312 60459
0 16591 5 1 1 16590
0 16592 7 1 2 65675 16591
0 16593 5 1 1 16592
0 16594 7 1 2 74089 16593
0 16595 5 1 1 16594
0 16596 7 1 2 16585 16595
0 16597 7 1 2 16578 16596
0 16598 7 1 2 16570 16597
0 16599 7 1 2 16537 16598
0 16600 7 1 2 16522 16599
0 16601 5 1 1 16600
0 16602 7 1 2 51290 16601
0 16603 5 1 1 16602
0 16604 7 2 2 57473 66742
0 16605 7 1 2 69835 74091
0 16606 5 1 1 16605
0 16607 7 1 2 68909 16606
0 16608 5 1 1 16607
0 16609 7 1 2 62721 16608
0 16610 5 1 1 16609
0 16611 7 1 2 69338 16610
0 16612 5 1 1 16611
0 16613 7 1 2 54605 16612
0 16614 5 1 1 16613
0 16615 7 1 2 69353 72535
0 16616 5 1 1 16615
0 16617 7 1 2 62722 69389
0 16618 5 1 1 16617
0 16619 7 1 2 74070 16618
0 16620 5 1 1 16619
0 16621 7 1 2 56064 16620
0 16622 5 1 1 16621
0 16623 7 1 2 16616 16622
0 16624 7 1 2 16614 16623
0 16625 5 2 1 16624
0 16626 7 1 2 56711 74093
0 16627 5 1 1 16626
0 16628 7 2 2 68468 68977
0 16629 5 1 1 74095
0 16630 7 1 2 59260 74096
0 16631 5 1 1 16630
0 16632 7 1 2 67936 68345
0 16633 5 2 1 16632
0 16634 7 1 2 16631 74097
0 16635 5 1 1 16634
0 16636 7 1 2 54606 16635
0 16637 5 1 1 16636
0 16638 7 1 2 62456 68902
0 16639 5 1 1 16638
0 16640 7 1 2 16637 16639
0 16641 5 1 1 16640
0 16642 7 1 2 54256 16641
0 16643 5 1 1 16642
0 16644 7 1 2 67544 68920
0 16645 7 1 2 71863 16644
0 16646 5 1 1 16645
0 16647 7 1 2 59261 69354
0 16648 5 1 1 16647
0 16649 7 1 2 57737 69355
0 16650 5 1 1 16649
0 16651 7 2 2 60389 69335
0 16652 7 1 2 50703 74099
0 16653 5 1 1 16652
0 16654 7 1 2 16650 16653
0 16655 5 1 1 16654
0 16656 7 1 2 62399 16655
0 16657 5 1 1 16656
0 16658 7 1 2 16648 16657
0 16659 7 1 2 16646 16658
0 16660 7 1 2 16643 16659
0 16661 7 1 2 16627 16660
0 16662 5 1 1 16661
0 16663 7 1 2 51291 16662
0 16664 5 1 1 16663
0 16665 7 2 2 62778 71995
0 16666 7 2 2 48359 71732
0 16667 7 1 2 60067 74103
0 16668 7 1 2 74101 16667
0 16669 5 1 1 16668
0 16670 7 1 2 16664 16669
0 16671 5 1 1 16670
0 16672 7 1 2 55739 16671
0 16673 5 1 1 16672
0 16674 7 1 2 59262 68998
0 16675 7 1 2 74102 16674
0 16676 5 2 1 16675
0 16677 7 1 2 16673 74105
0 16678 7 1 2 16603 16677
0 16679 5 1 1 16678
0 16680 7 1 2 62908 16679
0 16681 5 1 1 16680
0 16682 7 1 2 16462 16681
0 16683 5 1 1 16682
0 16684 7 1 2 57927 16683
0 16685 5 1 1 16684
0 16686 7 1 2 74032 71719
0 16687 5 1 1 16686
0 16688 7 1 2 16685 16687
0 16689 5 1 1 16688
0 16690 7 1 2 68221 16689
0 16691 5 1 1 16690
0 16692 7 2 2 72469 72828
0 16693 5 1 1 74107
0 16694 7 2 2 53790 54257
0 16695 7 1 2 73958 74109
0 16696 7 1 2 69756 16695
0 16697 5 1 1 16696
0 16698 7 1 2 16693 16697
0 16699 5 1 1 16698
0 16700 7 1 2 57474 16699
0 16701 5 1 1 16700
0 16702 7 2 2 54607 68254
0 16703 7 1 2 67553 74111
0 16704 5 1 1 16703
0 16705 7 2 2 54978 72097
0 16706 5 1 1 74113
0 16707 7 1 2 48149 74114
0 16708 5 1 1 16707
0 16709 7 1 2 16704 16708
0 16710 5 1 1 16709
0 16711 7 1 2 51742 16710
0 16712 5 1 1 16711
0 16713 7 1 2 16701 16712
0 16714 5 1 1 16713
0 16715 7 1 2 57928 16714
0 16716 5 1 1 16715
0 16717 7 1 2 64551 70084
0 16718 5 1 1 16717
0 16719 7 1 2 48150 71895
0 16720 5 1 1 16719
0 16721 7 1 2 16718 16720
0 16722 5 1 1 16721
0 16723 7 1 2 69265 16722
0 16724 5 1 1 16723
0 16725 7 1 2 16716 16724
0 16726 5 1 1 16725
0 16727 7 1 2 55521 16726
0 16728 5 1 1 16727
0 16729 7 1 2 67154 69266
0 16730 7 1 2 69456 16729
0 16731 5 1 1 16730
0 16732 7 1 2 16728 16731
0 16733 5 1 1 16732
0 16734 7 1 2 68141 16733
0 16735 5 1 1 16734
0 16736 7 3 2 49115 56065
0 16737 7 1 2 59544 74115
0 16738 5 1 1 16737
0 16739 7 1 2 57593 16738
0 16740 5 1 1 16739
0 16741 7 1 2 69275 16740
0 16742 5 1 1 16741
0 16743 7 1 2 73309 16742
0 16744 5 1 1 16743
0 16745 7 1 2 50043 16744
0 16746 5 1 1 16745
0 16747 7 1 2 69101 69472
0 16748 5 1 1 16747
0 16749 7 1 2 16746 16748
0 16750 5 1 1 16749
0 16751 7 1 2 49047 16750
0 16752 5 1 1 16751
0 16753 7 1 2 50044 64841
0 16754 7 1 2 71891 16753
0 16755 5 1 1 16754
0 16756 7 1 2 16752 16755
0 16757 5 1 1 16756
0 16758 7 1 2 61749 67937
0 16759 7 1 2 16757 16758
0 16760 5 1 1 16759
0 16761 7 1 2 16735 16760
0 16762 5 1 1 16761
0 16763 7 1 2 53900 16762
0 16764 5 1 1 16763
0 16765 7 1 2 64687 67157
0 16766 5 1 1 16765
0 16767 7 1 2 69201 16766
0 16768 5 1 1 16767
0 16769 7 1 2 61022 72098
0 16770 5 1 1 16769
0 16771 7 3 2 49116 72481
0 16772 7 1 2 47881 69896
0 16773 7 1 2 74118 16772
0 16774 5 1 1 16773
0 16775 7 1 2 16770 16774
0 16776 5 1 1 16775
0 16777 7 1 2 57929 16776
0 16778 5 1 1 16777
0 16779 7 2 2 54258 70085
0 16780 5 1 1 74121
0 16781 7 1 2 60918 74122
0 16782 5 1 1 16781
0 16783 7 1 2 49313 66823
0 16784 5 1 1 16783
0 16785 7 1 2 16782 16784
0 16786 5 1 1 16785
0 16787 7 1 2 68255 16786
0 16788 5 1 1 16787
0 16789 7 1 2 16778 16788
0 16790 5 1 1 16789
0 16791 7 1 2 48360 16790
0 16792 5 1 1 16791
0 16793 7 3 2 54259 58976
0 16794 7 4 2 47882 58147
0 16795 5 1 1 74126
0 16796 7 1 2 50704 16795
0 16797 5 1 1 16796
0 16798 7 1 2 69207 16797
0 16799 7 1 2 74123 16798
0 16800 5 1 1 16799
0 16801 7 1 2 16792 16800
0 16802 5 1 1 16801
0 16803 7 1 2 67938 16802
0 16804 5 1 1 16803
0 16805 7 1 2 16768 16804
0 16806 5 1 1 16805
0 16807 7 1 2 56712 16806
0 16808 5 1 1 16807
0 16809 7 1 2 56066 68109
0 16810 5 1 1 16809
0 16811 7 1 2 60919 66861
0 16812 5 1 1 16811
0 16813 7 1 2 7278 16812
0 16814 7 1 2 16810 16813
0 16815 5 1 1 16814
0 16816 7 1 2 72116 16815
0 16817 5 1 1 16816
0 16818 7 1 2 62400 60920
0 16819 5 1 1 16818
0 16820 7 1 2 50705 16819
0 16821 5 2 1 16820
0 16822 7 1 2 68256 69457
0 16823 7 1 2 74130 16822
0 16824 5 1 1 16823
0 16825 7 1 2 16817 16824
0 16826 5 1 1 16825
0 16827 7 1 2 51743 16826
0 16828 5 1 1 16827
0 16829 7 1 2 50706 60955
0 16830 5 2 1 16829
0 16831 7 1 2 69194 74132
0 16832 5 1 1 16831
0 16833 7 1 2 67595 70044
0 16834 5 1 1 16833
0 16835 7 1 2 71365 72830
0 16836 5 1 1 16835
0 16837 7 1 2 16836 72401
0 16838 5 1 1 16837
0 16839 7 1 2 16834 16838
0 16840 5 1 1 16839
0 16841 7 1 2 60921 16840
0 16842 5 1 1 16841
0 16843 7 1 2 16832 16842
0 16844 5 1 1 16843
0 16845 7 1 2 55646 68193
0 16846 7 1 2 16844 16845
0 16847 5 1 1 16846
0 16848 7 1 2 16828 16847
0 16849 5 1 1 16848
0 16850 7 1 2 55308 16849
0 16851 5 1 1 16850
0 16852 7 1 2 61119 68159
0 16853 5 3 1 16852
0 16854 7 1 2 69215 74134
0 16855 5 1 1 16854
0 16856 7 1 2 16851 16855
0 16857 7 1 2 16808 16856
0 16858 7 1 2 16764 16857
0 16859 5 1 1 16858
0 16860 7 1 2 60691 16859
0 16861 5 1 1 16860
0 16862 7 2 2 66871 68102
0 16863 5 1 1 74137
0 16864 7 1 2 72430 74138
0 16865 5 1 1 16864
0 16866 7 2 2 57930 72085
0 16867 7 1 2 61779 65219
0 16868 7 1 2 68103 16867
0 16869 5 3 1 16868
0 16870 7 1 2 74139 74141
0 16871 5 1 1 16870
0 16872 7 1 2 16865 16871
0 16873 5 1 1 16872
0 16874 7 1 2 54260 16873
0 16875 5 1 1 16874
0 16876 7 2 2 56067 71498
0 16877 5 2 1 74144
0 16878 7 1 2 59916 58918
0 16879 7 1 2 74146 16878
0 16880 5 1 1 16879
0 16881 7 1 2 74140 16880
0 16882 5 1 1 16881
0 16883 7 1 2 16875 16882
0 16884 5 1 1 16883
0 16885 7 1 2 55309 16884
0 16886 5 1 1 16885
0 16887 7 1 2 48151 68092
0 16888 5 2 1 16887
0 16889 7 1 2 48361 64300
0 16890 5 1 1 16889
0 16891 7 1 2 61028 16890
0 16892 7 1 2 74148 16891
0 16893 5 1 1 16892
0 16894 7 1 2 54261 16893
0 16895 5 1 1 16894
0 16896 7 1 2 51002 16895
0 16897 5 1 1 16896
0 16898 7 1 2 66087 16897
0 16899 5 1 1 16898
0 16900 7 1 2 57475 67740
0 16901 7 1 2 64769 16900
0 16902 5 1 1 16901
0 16903 7 1 2 67776 72655
0 16904 5 1 1 16903
0 16905 7 2 2 64408 66088
0 16906 5 2 1 74150
0 16907 7 1 2 16904 74152
0 16908 7 1 2 16902 16907
0 16909 7 1 2 16899 16908
0 16910 5 1 1 16909
0 16911 7 1 2 69267 16910
0 16912 5 1 1 16911
0 16913 7 1 2 16886 16912
0 16914 5 1 1 16913
0 16915 7 1 2 62554 16914
0 16916 5 1 1 16915
0 16917 7 1 2 51003 58211
0 16918 7 1 2 74147 16917
0 16919 5 2 1 16918
0 16920 7 1 2 57931 74154
0 16921 5 1 1 16920
0 16922 7 1 2 57932 74142
0 16923 5 1 1 16922
0 16924 7 1 2 16863 16923
0 16925 5 1 1 16924
0 16926 7 1 2 54262 16925
0 16927 5 1 1 16926
0 16928 7 1 2 16921 16927
0 16929 5 1 1 16928
0 16930 7 1 2 55310 16929
0 16931 5 1 1 16930
0 16932 7 1 2 64770 67155
0 16933 5 1 1 16932
0 16934 7 1 2 16931 16933
0 16935 5 1 1 16934
0 16936 7 1 2 48738 69197
0 16937 7 1 2 16935 16936
0 16938 5 1 1 16937
0 16939 7 1 2 61795 69216
0 16940 5 1 1 16939
0 16941 7 2 2 60634 62223
0 16942 7 4 2 56068 74156
0 16943 5 1 1 74158
0 16944 7 2 2 54979 74159
0 16945 7 1 2 61750 74162
0 16946 7 1 2 69202 16945
0 16947 5 1 1 16946
0 16948 7 1 2 16940 16947
0 16949 5 1 1 16948
0 16950 7 1 2 54608 16949
0 16951 5 1 1 16950
0 16952 7 2 2 59383 68364
0 16953 5 1 1 74164
0 16954 7 1 2 64730 74165
0 16955 5 1 1 16954
0 16956 7 1 2 69252 16955
0 16957 5 1 1 16956
0 16958 7 1 2 69268 16957
0 16959 5 1 1 16958
0 16960 7 1 2 16951 16959
0 16961 5 1 1 16960
0 16962 7 1 2 68116 16961
0 16963 5 1 1 16962
0 16964 7 1 2 54263 74108
0 16965 5 1 1 16964
0 16966 7 1 2 48739 72011
0 16967 7 1 2 70045 16966
0 16968 5 1 1 16967
0 16969 7 1 2 16965 16968
0 16970 5 1 1 16969
0 16971 7 1 2 67294 16970
0 16972 5 1 1 16971
0 16973 7 1 2 65981 68499
0 16974 7 1 2 69269 16973
0 16975 5 1 1 16974
0 16976 7 1 2 16972 16975
0 16977 5 1 1 16976
0 16978 7 1 2 68093 16977
0 16979 5 1 1 16978
0 16980 7 1 2 16963 16979
0 16981 7 1 2 16938 16980
0 16982 7 1 2 16916 16981
0 16983 7 1 2 64788 68117
0 16984 5 1 1 16983
0 16985 7 1 2 57738 62257
0 16986 7 1 2 74163 16985
0 16987 5 1 1 16986
0 16988 7 1 2 16984 16987
0 16989 5 1 1 16988
0 16990 7 1 2 69203 16989
0 16991 5 1 1 16990
0 16992 7 1 2 66926 68118
0 16993 5 1 1 16992
0 16994 7 1 2 47883 69009
0 16995 5 1 1 16994
0 16996 7 1 2 16993 16995
0 16997 5 1 1 16996
0 16998 7 1 2 72113 16997
0 16999 5 1 1 16998
0 17000 7 2 2 64254 72152
0 17001 7 1 2 59613 59136
0 17002 7 1 2 72516 17001
0 17003 7 1 2 74166 17002
0 17004 5 1 1 17003
0 17005 7 1 2 16999 17004
0 17006 5 1 1 17005
0 17007 7 1 2 55311 17006
0 17008 5 1 1 17007
0 17009 7 1 2 58212 68149
0 17010 5 1 1 17009
0 17011 7 1 2 60922 17010
0 17012 5 1 1 17011
0 17013 7 1 2 64015 17012
0 17014 5 1 1 17013
0 17015 7 1 2 69210 17014
0 17016 5 1 1 17015
0 17017 7 1 2 17008 17016
0 17018 5 1 1 17017
0 17019 7 1 2 55522 17018
0 17020 5 1 1 17019
0 17021 7 1 2 68257 69249
0 17022 5 1 1 17021
0 17023 7 1 2 17020 17022
0 17024 5 1 1 17023
0 17025 7 1 2 51744 17024
0 17026 5 1 1 17025
0 17027 7 1 2 16991 17026
0 17028 5 1 1 17027
0 17029 7 1 2 61553 17028
0 17030 5 1 1 17029
0 17031 7 1 2 68500 74143
0 17032 5 1 1 17031
0 17033 7 1 2 62211 66827
0 17034 7 2 2 48603 71843
0 17035 7 1 2 68077 74168
0 17036 7 1 2 17033 17035
0 17037 5 1 1 17036
0 17038 7 1 2 17032 17037
0 17039 5 1 1 17038
0 17040 7 1 2 54264 17039
0 17041 5 1 1 17040
0 17042 7 1 2 68501 74155
0 17043 5 1 1 17042
0 17044 7 1 2 17041 17043
0 17045 5 1 1 17044
0 17046 7 1 2 55312 17045
0 17047 5 1 1 17046
0 17048 7 1 2 57933 72656
0 17049 5 1 1 17048
0 17050 7 2 2 59328 67566
0 17051 5 1 1 74170
0 17052 7 1 2 48362 74171
0 17053 5 1 1 17052
0 17054 7 1 2 17049 17053
0 17055 5 1 1 17054
0 17056 7 1 2 68502 17055
0 17057 5 1 1 17056
0 17058 7 1 2 17047 17057
0 17059 5 1 1 17058
0 17060 7 1 2 72594 17059
0 17061 5 1 1 17060
0 17062 7 1 2 49198 64113
0 17063 5 1 1 17062
0 17064 7 2 2 47884 62258
0 17065 7 1 2 58675 74172
0 17066 5 1 1 17065
0 17067 7 1 2 66134 17066
0 17068 7 1 2 17063 17067
0 17069 5 1 1 17068
0 17070 7 1 2 56069 17069
0 17071 5 1 1 17070
0 17072 7 1 2 57476 67752
0 17073 5 1 1 17072
0 17074 7 1 2 60923 60390
0 17075 5 2 1 17074
0 17076 7 1 2 57594 74174
0 17077 5 2 1 17076
0 17078 7 1 2 63980 74176
0 17079 5 1 1 17078
0 17080 7 1 2 64158 17079
0 17081 5 1 1 17080
0 17082 7 1 2 48152 17081
0 17083 5 1 1 17082
0 17084 7 1 2 17073 17083
0 17085 7 1 2 17071 17084
0 17086 5 1 1 17085
0 17087 7 1 2 55313 72114
0 17088 7 1 2 17086 17087
0 17089 5 1 1 17088
0 17090 7 3 2 50707 57778
0 17091 5 1 1 74178
0 17092 7 1 2 57477 69208
0 17093 5 1 1 17092
0 17094 7 1 2 16706 17093
0 17095 5 1 1 17094
0 17096 7 1 2 57934 17095
0 17097 5 1 1 17096
0 17098 7 1 2 63829 72108
0 17099 5 1 1 17098
0 17100 7 1 2 17097 17099
0 17101 5 1 1 17100
0 17102 7 1 2 17091 17101
0 17103 5 1 1 17102
0 17104 7 1 2 51004 66930
0 17105 5 1 1 17104
0 17106 7 1 2 66799 68258
0 17107 7 1 2 17105 17106
0 17108 5 1 1 17107
0 17109 7 1 2 17103 17108
0 17110 7 1 2 17089 17109
0 17111 5 1 1 17110
0 17112 7 1 2 55523 17111
0 17113 5 1 1 17112
0 17114 7 1 2 17061 17113
0 17115 5 1 1 17114
0 17116 7 1 2 51745 17115
0 17117 5 1 1 17116
0 17118 7 1 2 17030 17117
0 17119 7 1 2 16982 17118
0 17120 7 1 2 16861 17119
0 17121 7 1 2 16691 17120
0 17122 7 1 2 16442 17121
0 17123 5 1 1 17122
0 17124 7 1 2 48937 17123
0 17125 5 1 1 17124
0 17126 7 1 2 63871 69055
0 17127 5 1 1 17126
0 17128 7 1 2 58977 74094
0 17129 5 1 1 17128
0 17130 7 1 2 17127 17129
0 17131 5 1 1 17130
0 17132 7 1 2 51292 17131
0 17133 5 1 1 17132
0 17134 7 1 2 63997 68322
0 17135 5 1 1 17134
0 17136 7 1 2 54980 72196
0 17137 7 1 2 64479 17136
0 17138 5 1 1 17137
0 17139 7 1 2 17135 17138
0 17140 5 1 1 17139
0 17141 7 1 2 57821 17140
0 17142 5 1 1 17141
0 17143 7 1 2 64412 64715
0 17144 5 4 1 17143
0 17145 7 1 2 74181 68323
0 17146 5 1 1 17145
0 17147 7 3 2 61904 67185
0 17148 7 1 2 56070 69729
0 17149 7 1 2 74185 17148
0 17150 5 1 1 17149
0 17151 7 1 2 17146 17150
0 17152 7 1 2 17142 17151
0 17153 5 1 1 17152
0 17154 7 1 2 53685 17153
0 17155 5 1 1 17154
0 17156 7 1 2 53478 57822
0 17157 7 1 2 67014 17156
0 17158 5 1 1 17157
0 17159 7 1 2 7540 17158
0 17160 5 1 1 17159
0 17161 7 1 2 56071 17160
0 17162 5 1 1 17161
0 17163 7 1 2 74182 71757
0 17164 5 1 1 17163
0 17165 7 1 2 71725 17164
0 17166 7 1 2 17162 17165
0 17167 5 1 1 17166
0 17168 7 1 2 69027 17167
0 17169 5 1 1 17168
0 17170 7 1 2 17155 17169
0 17171 5 1 1 17170
0 17172 7 1 2 55314 17171
0 17173 5 1 1 17172
0 17174 7 1 2 49914 69118
0 17175 7 1 2 63886 17174
0 17176 7 1 2 66951 17175
0 17177 7 1 2 63017 17176
0 17178 5 1 1 17177
0 17179 7 1 2 17173 17178
0 17180 7 1 2 17133 17179
0 17181 5 1 1 17180
0 17182 7 1 2 55740 17181
0 17183 5 1 1 17182
0 17184 7 1 2 64453 66469
0 17185 5 1 1 17184
0 17186 7 5 2 49314 51293
0 17187 7 2 2 48363 49915
0 17188 7 1 2 74188 74193
0 17189 5 1 1 17188
0 17190 7 1 2 17185 17189
0 17191 5 1 1 17190
0 17192 7 2 2 50421 65152
0 17193 5 5 1 74195
0 17194 7 1 2 17191 74197
0 17195 5 1 1 17194
0 17196 7 2 2 49916 68693
0 17197 5 1 1 74202
0 17198 7 1 2 64818 59601
0 17199 7 1 2 72460 17198
0 17200 5 1 1 17199
0 17201 7 1 2 17197 17200
0 17202 5 1 1 17201
0 17203 7 1 2 58386 17202
0 17204 5 1 1 17203
0 17205 7 1 2 49917 71978
0 17206 5 1 1 17205
0 17207 7 1 2 17204 17206
0 17208 5 1 1 17207
0 17209 7 1 2 54013 17208
0 17210 5 1 1 17209
0 17211 7 1 2 17195 17210
0 17212 5 1 1 17211
0 17213 7 1 2 55524 17212
0 17214 5 1 1 17213
0 17215 7 1 2 59985 66089
0 17216 5 1 1 17215
0 17217 7 1 2 67082 74169
0 17218 5 1 1 17217
0 17219 7 1 2 17216 17218
0 17220 5 1 1 17219
0 17221 7 1 2 49918 17220
0 17222 5 1 1 17221
0 17223 7 3 2 54609 66419
0 17224 7 1 2 67067 74204
0 17225 5 1 1 17224
0 17226 7 1 2 17222 17225
0 17227 5 1 1 17226
0 17228 7 1 2 64072 17227
0 17229 5 1 1 17228
0 17230 7 1 2 4882 17229
0 17231 5 1 1 17230
0 17232 7 1 2 56072 17231
0 17233 5 1 1 17232
0 17234 7 1 2 65373 67370
0 17235 5 1 1 17234
0 17236 7 1 2 51294 17235
0 17237 5 1 1 17236
0 17238 7 1 2 54610 17237
0 17239 5 1 1 17238
0 17240 7 1 2 58387 64789
0 17241 5 2 1 17240
0 17242 7 1 2 17239 74207
0 17243 5 1 1 17242
0 17244 7 1 2 57935 67777
0 17245 7 1 2 17243 17244
0 17246 5 1 1 17245
0 17247 7 1 2 17233 17246
0 17248 7 1 2 17214 17247
0 17249 5 1 1 17248
0 17250 7 1 2 62555 17249
0 17251 5 1 1 17250
0 17252 7 1 2 65374 65234
0 17253 7 1 2 69489 17252
0 17254 5 1 1 17253
0 17255 7 1 2 65148 59702
0 17256 5 1 1 17255
0 17257 7 1 2 61277 17256
0 17258 7 1 2 17254 17257
0 17259 5 1 1 17258
0 17260 7 1 2 66800 17259
0 17261 5 1 1 17260
0 17262 7 2 2 57478 60971
0 17263 7 1 2 69771 74209
0 17264 5 1 1 17263
0 17265 7 1 2 17261 17264
0 17266 5 1 1 17265
0 17267 7 1 2 68503 17266
0 17268 5 1 1 17267
0 17269 7 1 2 59654 65931
0 17270 5 2 1 17269
0 17271 7 1 2 54981 74211
0 17272 5 1 1 17271
0 17273 7 1 2 65261 61062
0 17274 5 2 1 17273
0 17275 7 1 2 17272 74213
0 17276 5 1 1 17275
0 17277 7 1 2 55315 68852
0 17278 7 1 2 17276 17277
0 17279 5 1 1 17278
0 17280 7 1 2 17268 17279
0 17281 5 1 1 17280
0 17282 7 1 2 55525 17281
0 17283 5 1 1 17282
0 17284 7 2 2 66964 72237
0 17285 7 1 2 58388 65885
0 17286 5 1 1 17285
0 17287 7 1 2 61120 17286
0 17288 5 2 1 17287
0 17289 7 1 2 64707 74217
0 17290 5 1 1 17289
0 17291 7 1 2 51295 17290
0 17292 5 1 1 17291
0 17293 7 1 2 54611 17292
0 17294 5 1 1 17293
0 17295 7 1 2 74208 17294
0 17296 5 1 1 17295
0 17297 7 1 2 74215 17296
0 17298 5 1 1 17297
0 17299 7 1 2 17283 17298
0 17300 7 1 2 17251 17299
0 17301 5 1 1 17300
0 17302 7 1 2 51746 17301
0 17303 5 1 1 17302
0 17304 7 2 2 47885 74183
0 17305 5 1 1 74219
0 17306 7 1 2 63469 74220
0 17307 5 1 1 17306
0 17308 7 2 2 51005 64929
0 17309 5 2 1 74221
0 17310 7 1 2 17307 74223
0 17311 5 1 1 17310
0 17312 7 1 2 54265 17311
0 17313 5 1 1 17312
0 17314 7 3 2 50708 56073
0 17315 7 1 2 64708 74225
0 17316 5 1 1 17315
0 17317 7 1 2 17313 17316
0 17318 5 1 1 17317
0 17319 7 1 2 69276 17318
0 17320 5 1 1 17319
0 17321 7 1 2 65812 69062
0 17322 5 1 1 17321
0 17323 7 1 2 17320 17322
0 17324 5 1 1 17323
0 17325 7 1 2 58389 17324
0 17326 5 1 1 17325
0 17327 7 1 2 66248 69277
0 17328 5 1 1 17327
0 17329 7 1 2 72899 17328
0 17330 5 1 1 17329
0 17331 7 1 2 61063 17330
0 17332 5 1 1 17331
0 17333 7 1 2 64758 59323
0 17334 5 1 1 17333
0 17335 7 1 2 17332 17334
0 17336 5 1 1 17335
0 17337 7 1 2 54982 17336
0 17338 5 1 1 17337
0 17339 7 1 2 17326 17338
0 17340 5 1 1 17339
0 17341 7 1 2 68860 17340
0 17342 5 1 1 17341
0 17343 7 1 2 17303 17342
0 17344 7 1 2 17183 17343
0 17345 5 1 1 17344
0 17346 7 1 2 56713 17345
0 17347 5 1 1 17346
0 17348 7 2 2 50422 59447
0 17349 5 1 1 74228
0 17350 7 1 2 55882 74229
0 17351 5 1 1 17350
0 17352 7 2 2 54014 62069
0 17353 5 4 1 74230
0 17354 7 1 2 73605 74232
0 17355 5 1 1 17354
0 17356 7 1 2 69051 72238
0 17357 7 1 2 17355 17356
0 17358 5 1 1 17357
0 17359 7 2 2 49117 53686
0 17360 7 2 2 52798 74236
0 17361 7 1 2 64484 68655
0 17362 7 1 2 74238 17361
0 17363 5 1 1 17362
0 17364 7 1 2 17358 17363
0 17365 5 1 1 17364
0 17366 7 1 2 55316 17365
0 17367 5 1 1 17366
0 17368 7 6 2 52799 68825
0 17369 5 1 1 74240
0 17370 7 2 2 69757 74241
0 17371 5 1 1 74246
0 17372 7 1 2 17367 17371
0 17373 5 1 1 17372
0 17374 7 1 2 51560 17373
0 17375 5 1 1 17374
0 17376 7 4 2 49732 68694
0 17377 5 1 1 74248
0 17378 7 1 2 62831 74249
0 17379 5 1 1 17378
0 17380 7 2 2 57226 74233
0 17381 5 2 1 74252
0 17382 7 1 2 54612 74254
0 17383 5 1 1 17382
0 17384 7 1 2 51006 17383
0 17385 5 1 1 17384
0 17386 7 1 2 66551 68180
0 17387 5 2 1 17386
0 17388 7 1 2 68817 74256
0 17389 5 1 1 17388
0 17390 7 1 2 55317 17389
0 17391 7 1 2 17385 17390
0 17392 5 1 1 17391
0 17393 7 1 2 17379 17392
0 17394 5 1 1 17393
0 17395 7 1 2 54266 17394
0 17396 5 1 1 17395
0 17397 7 1 2 50709 3286
0 17398 5 1 1 17397
0 17399 7 1 2 72124 17398
0 17400 7 1 2 72026 17399
0 17401 5 1 1 17400
0 17402 7 1 2 17396 17401
0 17403 5 1 1 17402
0 17404 7 1 2 67939 17403
0 17405 5 1 1 17404
0 17406 7 1 2 17375 17405
0 17407 5 1 1 17406
0 17408 7 1 2 56074 17407
0 17409 5 1 1 17408
0 17410 7 1 2 69052 74216
0 17411 5 1 1 17410
0 17412 7 1 2 17411 68724
0 17413 7 1 2 17409 17412
0 17414 5 1 1 17413
0 17415 7 1 2 17351 17414
0 17416 5 1 1 17415
0 17417 7 1 2 63926 74048
0 17418 5 1 1 17417
0 17419 7 1 2 58169 74066
0 17420 5 1 1 17419
0 17421 7 1 2 54613 74058
0 17422 5 1 1 17421
0 17423 7 1 2 17420 17422
0 17424 7 1 2 17418 17423
0 17425 5 1 1 17424
0 17426 7 1 2 51296 17425
0 17427 5 1 1 17426
0 17428 7 1 2 74034 74064
0 17429 5 1 1 17428
0 17430 7 1 2 51297 17429
0 17431 5 1 1 17430
0 17432 7 1 2 63964 68346
0 17433 7 1 2 71640 17432
0 17434 5 1 1 17433
0 17435 7 1 2 17431 17434
0 17436 5 1 1 17435
0 17437 7 1 2 54267 17436
0 17438 5 1 1 17437
0 17439 7 1 2 64510 69378
0 17440 5 1 1 17439
0 17441 7 1 2 74039 17440
0 17442 5 1 1 17441
0 17443 7 1 2 48364 17442
0 17444 5 1 1 17443
0 17445 7 1 2 47886 74049
0 17446 5 1 1 17445
0 17447 7 1 2 17444 17446
0 17448 5 1 1 17447
0 17449 7 1 2 51298 17448
0 17450 5 1 1 17449
0 17451 7 1 2 17438 17450
0 17452 5 1 1 17451
0 17453 7 1 2 57153 17452
0 17454 5 1 1 17453
0 17455 7 1 2 17427 17454
0 17456 5 1 1 17455
0 17457 7 1 2 55741 17456
0 17458 5 1 1 17457
0 17459 7 1 2 64063 74042
0 17460 5 1 1 17459
0 17461 7 1 2 63939 74060
0 17462 5 1 1 17461
0 17463 7 1 2 61080 74080
0 17464 5 1 1 17463
0 17465 7 1 2 58715 70203
0 17466 5 1 1 17465
0 17467 7 1 2 68903 17466
0 17468 5 1 1 17467
0 17469 7 1 2 17464 17468
0 17470 7 1 2 17462 17469
0 17471 7 1 2 17460 17470
0 17472 5 1 1 17471
0 17473 7 1 2 57154 17472
0 17474 5 1 1 17473
0 17475 7 1 2 69386 74098
0 17476 7 1 2 13821 17475
0 17477 5 1 1 17476
0 17478 7 1 2 59614 17477
0 17479 5 1 1 17478
0 17480 7 1 2 65946 69356
0 17481 5 1 1 17480
0 17482 7 1 2 61099 74054
0 17483 5 1 1 17482
0 17484 7 1 2 17481 17483
0 17485 7 1 2 17479 17484
0 17486 5 1 1 17485
0 17487 7 1 2 48365 17486
0 17488 5 1 1 17487
0 17489 7 1 2 61023 69357
0 17490 5 1 1 17489
0 17491 7 1 2 57823 74050
0 17492 5 1 1 17491
0 17493 7 1 2 17490 17492
0 17494 5 1 1 17493
0 17495 7 1 2 54015 17494
0 17496 5 1 1 17495
0 17497 7 1 2 51007 65790
0 17498 5 2 1 17497
0 17499 7 1 2 68904 74258
0 17500 5 1 1 17499
0 17501 7 1 2 17496 17500
0 17502 7 1 2 17488 17501
0 17503 7 1 2 17474 17502
0 17504 5 1 1 17503
0 17505 7 1 2 51299 17504
0 17506 5 1 1 17505
0 17507 7 1 2 74106 17506
0 17508 7 1 2 17458 17507
0 17509 5 1 1 17508
0 17510 7 1 2 58978 17509
0 17511 5 1 1 17510
0 17512 7 1 2 17416 17511
0 17513 7 1 2 67799 71727
0 17514 5 1 1 17513
0 17515 7 1 2 67635 17514
0 17516 5 1 1 17515
0 17517 7 1 2 16953 69707
0 17518 5 1 1 17517
0 17519 7 1 2 49315 17518
0 17520 5 1 1 17519
0 17521 7 2 2 73974 69930
0 17522 5 1 1 74260
0 17523 7 1 2 17520 17522
0 17524 5 1 1 17523
0 17525 7 1 2 63018 17524
0 17526 5 1 1 17525
0 17527 7 1 2 59502 67831
0 17528 7 1 2 71971 17527
0 17529 5 1 1 17528
0 17530 7 1 2 17526 17529
0 17531 5 1 1 17530
0 17532 7 1 2 48366 17531
0 17533 5 1 1 17532
0 17534 7 4 2 55526 68695
0 17535 7 1 2 62909 74262
0 17536 5 1 1 17535
0 17537 7 1 2 49316 62556
0 17538 7 1 2 74261 17537
0 17539 5 1 1 17538
0 17540 7 1 2 17536 17539
0 17541 5 1 1 17540
0 17542 7 1 2 57936 17541
0 17543 5 1 1 17542
0 17544 7 1 2 64614 71733
0 17545 7 1 2 73971 17544
0 17546 5 1 1 17545
0 17547 7 1 2 17543 17546
0 17548 7 1 2 17533 17547
0 17549 5 1 1 17548
0 17550 7 1 2 57155 17549
0 17551 5 1 1 17550
0 17552 7 1 2 17516 17551
0 17553 5 1 1 17552
0 17554 7 1 2 51747 17553
0 17555 5 1 1 17554
0 17556 7 1 2 68725 17555
0 17557 5 1 1 17556
0 17558 7 1 2 68142 17557
0 17559 5 1 1 17558
0 17560 7 1 2 53901 66430
0 17561 5 1 1 17560
0 17562 7 1 2 56075 71662
0 17563 5 1 1 17562
0 17564 7 1 2 17561 17563
0 17565 5 1 1 17564
0 17566 7 1 2 61147 17565
0 17567 5 1 1 17566
0 17568 7 1 2 49919 72148
0 17569 5 1 1 17568
0 17570 7 1 2 17567 17569
0 17571 5 1 1 17570
0 17572 7 1 2 54016 17571
0 17573 5 1 1 17572
0 17574 7 6 2 50710 60391
0 17575 5 1 1 74266
0 17576 7 1 2 68365 74267
0 17577 5 1 1 17576
0 17578 7 1 2 73976 17577
0 17579 5 1 1 17578
0 17580 7 1 2 57479 17579
0 17581 5 1 1 17580
0 17582 7 1 2 67623 17581
0 17583 7 1 2 17573 17582
0 17584 5 1 1 17583
0 17585 7 1 2 67993 17584
0 17586 5 1 1 17585
0 17587 7 1 2 65246 63405
0 17588 7 1 2 67520 17587
0 17589 7 1 2 71946 17588
0 17590 5 1 1 17589
0 17591 7 1 2 71713 17590
0 17592 5 1 1 17591
0 17593 7 1 2 54983 17592
0 17594 5 1 1 17593
0 17595 7 1 2 57480 59602
0 17596 5 1 1 17595
0 17597 7 1 2 53479 65247
0 17598 7 1 2 61306 17597
0 17599 5 1 1 17598
0 17600 7 1 2 17596 17599
0 17601 5 1 1 17600
0 17602 7 1 2 72039 17601
0 17603 5 1 1 17602
0 17604 7 1 2 17594 17603
0 17605 5 1 1 17604
0 17606 7 1 2 55318 17605
0 17607 5 1 1 17606
0 17608 7 1 2 65254 59698
0 17609 5 1 1 17608
0 17610 7 1 2 68736 17609
0 17611 5 1 1 17610
0 17612 7 1 2 17607 17611
0 17613 7 1 2 17586 17612
0 17614 5 1 1 17613
0 17615 7 1 2 57156 17614
0 17616 5 1 1 17615
0 17617 7 2 2 69794 69102
0 17618 5 1 1 74272
0 17619 7 1 2 62910 74189
0 17620 7 1 2 66329 17619
0 17621 5 1 1 17620
0 17622 7 1 2 17618 17621
0 17623 5 1 1 17622
0 17624 7 1 2 48367 17623
0 17625 5 1 1 17624
0 17626 7 1 2 59675 74273
0 17627 5 1 1 17626
0 17628 7 1 2 67636 68709
0 17629 5 1 1 17628
0 17630 7 1 2 17627 17629
0 17631 7 1 2 17625 17630
0 17632 5 1 1 17631
0 17633 7 1 2 55527 17632
0 17634 5 1 1 17633
0 17635 7 1 2 63906 71649
0 17636 5 1 1 17635
0 17637 7 1 2 61307 66486
0 17638 5 1 1 17637
0 17639 7 1 2 17636 17638
0 17640 5 1 1 17639
0 17641 7 1 2 54984 17640
0 17642 5 1 1 17641
0 17643 7 2 2 65982 68643
0 17644 5 1 1 74274
0 17645 7 1 2 17642 17644
0 17646 5 1 1 17645
0 17647 7 1 2 63019 17646
0 17648 5 1 1 17647
0 17649 7 1 2 17634 17648
0 17650 7 1 2 17616 17649
0 17651 5 1 1 17650
0 17652 7 1 2 51748 17651
0 17653 5 1 1 17652
0 17654 7 1 2 59703 59324
0 17655 5 1 1 17654
0 17656 7 3 2 59391 62605
0 17657 7 1 2 72387 74276
0 17658 5 1 1 17657
0 17659 7 1 2 55883 58716
0 17660 5 1 1 17659
0 17661 7 1 2 52800 17660
0 17662 7 1 2 73996 17661
0 17663 5 1 1 17662
0 17664 7 1 2 17658 17663
0 17665 5 1 1 17664
0 17666 7 1 2 57157 17665
0 17667 5 1 1 17666
0 17668 7 1 2 17655 17667
0 17669 5 1 1 17668
0 17670 7 1 2 73304 68469
0 17671 7 1 2 17669 17670
0 17672 5 1 1 17671
0 17673 7 1 2 17653 17672
0 17674 5 1 1 17673
0 17675 7 1 2 58854 17674
0 17676 5 1 1 17675
0 17677 7 1 2 17559 17676
0 17678 7 1 2 17512 17677
0 17679 7 1 2 65748 72233
0 17680 5 1 1 17679
0 17681 7 1 2 60924 69605
0 17682 7 1 2 17680 17681
0 17683 5 1 1 17682
0 17684 7 1 2 65587 67778
0 17685 5 1 1 17684
0 17686 7 1 2 68733 17685
0 17687 7 1 2 17683 17686
0 17688 5 1 1 17687
0 17689 7 1 2 57158 17688
0 17690 5 1 1 17689
0 17691 7 1 2 67779 68059
0 17692 5 1 1 17691
0 17693 7 1 2 66441 17692
0 17694 5 1 1 17693
0 17695 7 1 2 57481 17694
0 17696 5 1 1 17695
0 17697 7 1 2 69441 72508
0 17698 5 1 1 17697
0 17699 7 1 2 17698 68565
0 17700 7 1 2 17696 17699
0 17701 7 1 2 17690 17700
0 17702 5 1 1 17701
0 17703 7 1 2 54268 17702
0 17704 5 1 1 17703
0 17705 7 1 2 66470 74255
0 17706 5 1 1 17705
0 17707 7 1 2 68601 17706
0 17708 5 1 1 17707
0 17709 7 1 2 57482 17708
0 17710 5 1 1 17709
0 17711 7 1 2 73310 17710
0 17712 5 1 1 17711
0 17713 7 1 2 55528 17712
0 17714 5 1 1 17713
0 17715 7 1 2 17714 68633
0 17716 7 1 2 17704 17715
0 17717 5 1 1 17716
0 17718 7 1 2 54614 17717
0 17719 5 1 1 17718
0 17720 7 1 2 54985 67805
0 17721 5 1 1 17720
0 17722 7 1 2 57595 74253
0 17723 5 1 1 17722
0 17724 7 1 2 60635 67780
0 17725 7 1 2 17723 17724
0 17726 5 1 1 17725
0 17727 7 1 2 17721 17726
0 17728 5 1 1 17727
0 17729 7 1 2 55319 17728
0 17730 5 1 1 17729
0 17731 7 1 2 68540 17730
0 17732 7 1 2 17719 17731
0 17733 5 1 1 17732
0 17734 7 1 2 68194 17733
0 17735 5 1 1 17734
0 17736 7 1 2 57159 74177
0 17737 5 1 1 17736
0 17738 7 2 2 50423 74234
0 17739 5 2 1 74279
0 17740 7 1 2 57483 74281
0 17741 5 1 1 17740
0 17742 7 1 2 17737 17741
0 17743 5 1 1 17742
0 17744 7 1 2 54615 17743
0 17745 5 1 1 17744
0 17746 7 1 2 51008 17745
0 17747 5 1 1 17746
0 17748 7 1 2 64471 71776
0 17749 7 1 2 17747 17748
0 17750 5 1 1 17749
0 17751 7 1 2 17735 17750
0 17752 5 1 1 17751
0 17753 7 1 2 51749 17752
0 17754 5 1 1 17753
0 17755 7 20 2 53480 54986
0 17756 5 1 1 74283
0 17757 7 2 2 74284 72491
0 17758 5 1 1 74303
0 17759 7 1 2 51561 74304
0 17760 5 1 1 17759
0 17761 7 1 2 63284 65730
0 17762 5 1 1 17761
0 17763 7 1 2 67800 17762
0 17764 5 1 1 17763
0 17765 7 1 2 59676 17764
0 17766 5 1 1 17765
0 17767 7 1 2 67717 67476
0 17768 5 1 1 17767
0 17769 7 1 2 12578 17768
0 17770 7 1 2 17766 17769
0 17771 5 1 1 17770
0 17772 7 1 2 51750 67678
0 17773 7 1 2 17771 17772
0 17774 5 1 1 17773
0 17775 7 1 2 17760 17774
0 17776 5 1 1 17775
0 17777 7 1 2 55742 17776
0 17778 5 1 1 17777
0 17779 7 2 2 68826 72054
0 17780 7 1 2 58676 66176
0 17781 7 1 2 74305 17780
0 17782 5 1 1 17781
0 17783 7 1 2 17778 17782
0 17784 5 1 1 17783
0 17785 7 1 2 47887 17784
0 17786 5 1 1 17785
0 17787 7 1 2 63572 68992
0 17788 7 1 2 69119 17787
0 17789 7 1 2 64969 17788
0 17790 5 1 1 17789
0 17791 7 1 2 17786 17790
0 17792 5 1 1 17791
0 17793 7 1 2 54017 17792
0 17794 5 1 1 17793
0 17795 7 1 2 51009 57852
0 17796 5 1 1 17795
0 17797 7 1 2 59704 17796
0 17798 5 1 1 17797
0 17799 7 1 2 51010 61121
0 17800 5 1 1 17799
0 17801 7 1 2 54616 17800
0 17802 5 1 1 17801
0 17803 7 1 2 17798 17802
0 17804 5 1 1 17803
0 17805 7 1 2 74306 17804
0 17806 5 1 1 17805
0 17807 7 1 2 51300 66941
0 17808 5 1 1 17807
0 17809 7 1 2 54987 17808
0 17810 5 1 1 17809
0 17811 7 1 2 64684 60636
0 17812 5 1 1 17811
0 17813 7 1 2 17810 17812
0 17814 5 1 1 17813
0 17815 7 1 2 69033 17814
0 17816 5 1 1 17815
0 17817 7 1 2 69795 68984
0 17818 5 1 1 17817
0 17819 7 1 2 68771 68963
0 17820 7 1 2 71499 17819
0 17821 5 1 1 17820
0 17822 7 1 2 17758 17821
0 17823 5 1 1 17822
0 17824 7 1 2 61308 17823
0 17825 5 1 1 17824
0 17826 7 1 2 17818 17825
0 17827 7 1 2 17816 17826
0 17828 5 1 1 17827
0 17829 7 1 2 51562 17828
0 17830 5 1 1 17829
0 17831 7 1 2 17806 17830
0 17832 7 1 2 17794 17831
0 17833 5 1 1 17832
0 17834 7 1 2 58113 17833
0 17835 5 1 1 17834
0 17836 7 1 2 50711 65886
0 17837 5 1 1 17836
0 17838 7 4 2 47888 50424
0 17839 7 2 2 71417 74307
0 17840 5 1 1 74311
0 17841 7 1 2 17837 17840
0 17842 5 1 1 17841
0 17843 7 1 2 69336 17842
0 17844 5 1 1 17843
0 17845 7 1 2 47889 64959
0 17846 5 1 1 17845
0 17847 7 1 2 64016 17846
0 17848 5 2 1 17847
0 17849 7 1 2 67940 69747
0 17850 7 1 2 74313 17849
0 17851 5 1 1 17850
0 17852 7 1 2 17844 17851
0 17853 5 1 1 17852
0 17854 7 1 2 49733 17853
0 17855 5 1 1 17854
0 17856 7 1 2 74285 69060
0 17857 5 1 1 17856
0 17858 7 1 2 74062 17857
0 17859 5 1 1 17858
0 17860 7 1 2 54018 17859
0 17861 5 1 1 17860
0 17862 7 1 2 63285 68905
0 17863 5 1 1 17862
0 17864 7 1 2 17861 17863
0 17865 7 1 2 47890 74082
0 17866 5 1 1 17865
0 17867 7 1 2 61100 74090
0 17868 5 1 1 17867
0 17869 7 1 2 17866 17868
0 17870 7 1 2 17864 17869
0 17871 5 1 1 17870
0 17872 7 1 2 58114 17871
0 17873 5 1 1 17872
0 17874 7 1 2 55529 69979
0 17875 7 1 2 68721 17874
0 17876 5 1 1 17875
0 17877 7 1 2 17873 17876
0 17878 7 1 2 17855 17877
0 17879 5 1 1 17878
0 17880 7 1 2 51301 17879
0 17881 5 1 1 17880
0 17882 7 1 2 61714 67567
0 17883 7 1 2 67994 17882
0 17884 5 1 1 17883
0 17885 7 1 2 67638 17884
0 17886 5 1 1 17885
0 17887 7 1 2 69028 17886
0 17888 5 1 1 17887
0 17889 7 1 2 54019 74247
0 17890 5 1 1 17889
0 17891 7 1 2 17888 17890
0 17892 5 1 1 17891
0 17893 7 1 2 51563 17892
0 17894 5 1 1 17893
0 17895 7 3 2 53481 68347
0 17896 7 1 2 67718 74315
0 17897 5 1 1 17896
0 17898 7 1 2 66819 68620
0 17899 5 2 1 17898
0 17900 7 2 2 51564 59986
0 17901 7 1 2 49920 74320
0 17902 5 1 1 17901
0 17903 7 1 2 74318 17902
0 17904 5 1 1 17903
0 17905 7 1 2 63020 17904
0 17906 5 1 1 17905
0 17907 7 1 2 17897 17906
0 17908 5 1 1 17907
0 17909 7 1 2 56076 17908
0 17910 5 1 1 17909
0 17911 7 2 2 63021 67521
0 17912 5 1 1 74322
0 17913 7 1 2 68954 74323
0 17914 5 1 1 17913
0 17915 7 1 2 64931 17305
0 17916 5 2 1 17915
0 17917 7 1 2 55530 68781
0 17918 7 1 2 74324 17917
0 17919 5 1 1 17918
0 17920 7 1 2 17914 17919
0 17921 7 1 2 17910 17920
0 17922 5 1 1 17921
0 17923 7 1 2 51751 17922
0 17924 5 1 1 17923
0 17925 7 1 2 74100 71691
0 17926 5 1 1 17925
0 17927 7 1 2 64676 72826
0 17928 5 1 1 17927
0 17929 7 1 2 17926 17928
0 17930 7 1 2 17924 17929
0 17931 5 1 1 17930
0 17932 7 1 2 55320 17931
0 17933 5 1 1 17932
0 17934 7 1 2 17894 17933
0 17935 7 1 2 17881 17934
0 17936 5 1 1 17935
0 17937 7 1 2 61971 17936
0 17938 5 1 1 17937
0 17939 7 1 2 54988 62432
0 17940 5 2 1 17939
0 17941 7 1 2 60953 63998
0 17942 5 1 1 17941
0 17943 7 1 2 74326 17942
0 17944 5 1 1 17943
0 17945 7 1 2 68324 17944
0 17946 5 1 1 17945
0 17947 7 1 2 59637 63956
0 17948 5 1 1 17947
0 17949 7 1 2 59325 17948
0 17950 5 1 1 17949
0 17951 7 2 2 62212 62864
0 17952 5 1 1 74328
0 17953 7 1 2 59020 74127
0 17954 7 1 2 74329 17953
0 17955 5 1 1 17954
0 17956 7 1 2 17950 17955
0 17957 5 1 1 17956
0 17958 7 1 2 68474 17957
0 17959 5 1 1 17958
0 17960 7 1 2 17946 17959
0 17961 5 1 1 17960
0 17962 7 1 2 53687 17961
0 17963 5 1 1 17962
0 17964 7 1 2 49199 67078
0 17965 7 1 2 74116 17964
0 17966 5 1 1 17965
0 17967 7 1 2 74327 17966
0 17968 5 1 1 17967
0 17969 7 1 2 71758 17968
0 17970 5 1 1 17969
0 17971 7 1 2 74133 68428
0 17972 5 1 1 17971
0 17973 7 1 2 17970 17972
0 17974 5 1 1 17973
0 17975 7 1 2 69029 17974
0 17976 5 1 1 17975
0 17977 7 1 2 17963 17976
0 17978 5 1 1 17977
0 17979 7 1 2 55321 17978
0 17980 5 1 1 17979
0 17981 7 1 2 48368 71741
0 17982 5 1 1 17981
0 17983 7 1 2 69064 17982
0 17984 5 1 1 17983
0 17985 7 1 2 57160 17984
0 17986 5 1 1 17985
0 17987 7 1 2 63286 72197
0 17988 5 1 1 17987
0 17989 7 1 2 17988 68327
0 17990 5 1 1 17989
0 17991 7 1 2 53688 17990
0 17992 5 1 1 17991
0 17993 7 2 2 67941 68807
0 17994 5 1 1 74330
0 17995 7 1 2 17992 17994
0 17996 5 1 1 17995
0 17997 7 1 2 63830 17996
0 17998 5 1 1 17997
0 17999 7 1 2 17986 17998
0 18000 5 1 1 17999
0 18001 7 1 2 59677 18000
0 18002 5 1 1 18001
0 18003 7 1 2 59615 62433
0 18004 7 1 2 71742 18003
0 18005 5 1 1 18004
0 18006 7 1 2 18002 18005
0 18007 7 1 2 17980 18006
0 18008 5 1 1 18007
0 18009 7 1 2 60692 18008
0 18010 5 1 1 18009
0 18011 7 2 2 58390 66746
0 18012 5 1 1 74332
0 18013 7 1 2 61122 18012
0 18014 5 1 1 18013
0 18015 7 1 2 57161 18014
0 18016 5 1 1 18015
0 18017 7 1 2 50712 74235
0 18018 5 1 1 18017
0 18019 7 1 2 61270 18018
0 18020 5 1 1 18019
0 18021 7 1 2 18016 18020
0 18022 5 1 1 18021
0 18023 7 1 2 55322 18022
0 18024 5 1 1 18023
0 18025 7 1 2 66377 74282
0 18026 5 1 1 18025
0 18027 7 1 2 18024 18026
0 18028 5 1 1 18027
0 18029 7 1 2 54989 18028
0 18030 5 1 1 18029
0 18031 7 1 2 67688 18030
0 18032 5 1 1 18031
0 18033 7 1 2 51565 18032
0 18034 5 1 1 18033
0 18035 7 1 2 67015 66712
0 18036 5 1 1 18035
0 18037 7 1 2 18034 18036
0 18038 5 1 1 18037
0 18039 7 1 2 69732 18038
0 18040 5 1 1 18039
0 18041 7 1 2 18010 18040
0 18042 7 1 2 17938 18041
0 18043 7 1 2 17835 18042
0 18044 7 1 2 17754 18043
0 18045 7 1 2 17678 18044
0 18046 7 1 2 17347 18045
0 18047 5 1 1 18046
0 18048 7 1 2 68259 18047
0 18049 5 1 1 18048
0 18050 7 6 2 51302 70016
0 18051 7 1 2 55531 65854
0 18052 7 2 2 74334 18051
0 18053 5 1 1 74340
0 18054 7 1 2 47891 69598
0 18055 5 1 1 18054
0 18056 7 1 2 74319 18055
0 18057 5 1 1 18056
0 18058 7 1 2 64117 18057
0 18059 5 1 1 18058
0 18060 7 1 2 18053 18059
0 18061 5 1 1 18060
0 18062 7 1 2 50045 18061
0 18063 5 1 1 18062
0 18064 7 1 2 65855 68580
0 18065 5 2 1 18064
0 18066 7 1 2 64593 69959
0 18067 5 1 1 18066
0 18068 7 1 2 74342 18067
0 18069 5 2 1 18068
0 18070 7 4 2 65628 67832
0 18071 7 1 2 74344 74346
0 18072 5 1 1 18071
0 18073 7 1 2 18063 18072
0 18074 5 1 1 18073
0 18075 7 1 2 49048 18074
0 18076 5 1 1 18075
0 18077 7 2 2 53482 64594
0 18078 5 2 1 74350
0 18079 7 1 2 60392 74351
0 18080 5 1 1 18079
0 18081 7 1 2 74343 18080
0 18082 5 2 1 18081
0 18083 7 5 2 49921 65629
0 18084 7 2 2 72644 74356
0 18085 7 1 2 74354 74361
0 18086 5 1 1 18085
0 18087 7 1 2 18076 18086
0 18088 5 1 1 18087
0 18089 7 1 2 49118 18088
0 18090 5 1 1 18089
0 18091 7 1 2 17349 69599
0 18092 5 1 1 18091
0 18093 7 1 2 67020 73990
0 18094 5 1 1 18093
0 18095 7 1 2 18092 18094
0 18096 5 1 1 18095
0 18097 7 1 2 64118 18096
0 18098 5 1 1 18097
0 18099 7 1 2 50089 61922
0 18100 5 1 1 18099
0 18101 7 1 2 74341 18100
0 18102 5 1 1 18101
0 18103 7 1 2 18098 18102
0 18104 5 1 1 18103
0 18105 7 1 2 50046 18104
0 18106 5 1 1 18105
0 18107 7 1 2 53902 74345
0 18108 5 1 1 18107
0 18109 7 1 2 67657 68696
0 18110 5 2 1 18109
0 18111 7 1 2 18108 74363
0 18112 5 1 1 18111
0 18113 7 1 2 18112 74347
0 18114 5 1 1 18113
0 18115 7 1 2 18106 18114
0 18116 5 1 1 18115
0 18117 7 1 2 49049 18116
0 18118 5 1 1 18117
0 18119 7 1 2 53903 74355
0 18120 5 1 1 18119
0 18121 7 1 2 74364 18120
0 18122 5 1 1 18121
0 18123 7 1 2 18122 74362
0 18124 5 1 1 18123
0 18125 7 1 2 18118 18124
0 18126 7 1 2 18090 18125
0 18127 5 1 1 18126
0 18128 7 1 2 48153 18127
0 18129 5 1 1 18128
0 18130 7 2 2 50047 62557
0 18131 7 1 2 67719 67545
0 18132 5 1 1 18131
0 18133 7 1 2 8574 18132
0 18134 5 1 1 18133
0 18135 7 1 2 74365 18134
0 18136 5 1 1 18135
0 18137 7 3 2 65614 72239
0 18138 7 1 2 68614 69499
0 18139 7 1 2 74367 18138
0 18140 5 1 1 18139
0 18141 7 1 2 18136 18140
0 18142 5 1 1 18141
0 18143 7 1 2 49050 18142
0 18144 5 1 1 18143
0 18145 7 2 2 53483 72302
0 18146 7 2 2 66943 74370
0 18147 7 1 2 67720 74372
0 18148 5 1 1 18147
0 18149 7 1 2 18144 18148
0 18150 5 1 1 18149
0 18151 7 1 2 67587 18150
0 18152 5 1 1 18151
0 18153 7 1 2 57755 65676
0 18154 5 3 1 18153
0 18155 7 1 2 66090 74374
0 18156 7 1 2 72219 18155
0 18157 5 1 1 18156
0 18158 7 1 2 18152 18157
0 18159 5 1 1 18158
0 18160 7 1 2 58391 18159
0 18161 5 1 1 18160
0 18162 7 1 2 18129 18161
0 18163 5 1 1 18162
0 18164 7 1 2 49200 18163
0 18165 5 1 1 18164
0 18166 7 2 2 68697 70002
0 18167 7 1 2 68222 68615
0 18168 7 1 2 74377 18167
0 18169 5 1 1 18168
0 18170 7 1 2 67016 74335
0 18171 5 1 1 18170
0 18172 7 1 2 69567 69606
0 18173 7 1 2 71875 18172
0 18174 5 1 1 18173
0 18175 7 1 2 18171 18174
0 18176 5 1 1 18175
0 18177 7 1 2 54269 18176
0 18178 5 1 1 18177
0 18179 7 1 2 18178 72856
0 18180 5 1 1 18179
0 18181 7 1 2 68260 18180
0 18182 5 1 1 18181
0 18183 7 1 2 18169 18182
0 18184 5 1 1 18183
0 18185 7 1 2 55743 18184
0 18186 5 1 1 18185
0 18187 7 1 2 62911 60235
0 18188 5 1 1 18187
0 18189 7 1 2 54617 64119
0 18190 5 1 1 18189
0 18191 7 1 2 18188 18190
0 18192 5 1 1 18191
0 18193 7 1 2 69568 18192
0 18194 5 1 1 18193
0 18195 7 1 2 60236 69617
0 18196 5 1 1 18195
0 18197 7 1 2 18194 18196
0 18198 5 1 1 18197
0 18199 7 1 2 72595 18198
0 18200 5 1 1 18199
0 18201 7 1 2 18186 18200
0 18202 7 1 2 18165 18201
0 18203 5 1 1 18202
0 18204 7 1 2 54990 18203
0 18205 5 1 1 18204
0 18206 7 1 2 71659 71390
0 18207 5 1 1 18206
0 18208 7 1 2 70017 68332
0 18209 5 1 1 18208
0 18210 7 1 2 60835 57280
0 18211 5 1 1 18210
0 18212 7 1 2 59727 18211
0 18213 5 1 1 18212
0 18214 7 1 2 47892 18213
0 18215 5 1 1 18214
0 18216 7 1 2 65214 18215
0 18217 5 1 1 18216
0 18218 7 1 2 66521 70065
0 18219 7 1 2 18217 18218
0 18220 5 1 1 18219
0 18221 7 1 2 18209 18220
0 18222 5 1 1 18221
0 18223 7 1 2 68261 18222
0 18224 5 1 1 18223
0 18225 7 1 2 18207 18224
0 18226 7 1 2 18205 18225
0 18227 5 1 1 18226
0 18228 7 1 2 51752 18227
0 18229 5 1 1 18228
0 18230 7 1 2 72645 74378
0 18231 5 1 1 18230
0 18232 7 4 2 50048 54020
0 18233 7 1 2 65983 74379
0 18234 5 1 1 18233
0 18235 7 2 2 66091 68772
0 18236 7 1 2 54618 74383
0 18237 5 1 1 18236
0 18238 7 1 2 18234 18237
0 18239 5 1 1 18238
0 18240 7 1 2 48938 18239
0 18241 5 1 1 18240
0 18242 7 2 2 66092 66378
0 18243 5 1 1 74385
0 18244 7 1 2 7446 18243
0 18245 5 1 1 18244
0 18246 7 1 2 50049 18245
0 18247 5 1 1 18246
0 18248 7 1 2 18241 18247
0 18249 5 1 1 18248
0 18250 7 1 2 48740 18249
0 18251 5 1 1 18250
0 18252 7 1 2 65984 67658
0 18253 5 2 1 18252
0 18254 7 1 2 71835 74387
0 18255 5 2 1 18254
0 18256 7 1 2 72205 74389
0 18257 5 1 1 18256
0 18258 7 1 2 18251 18257
0 18259 5 1 1 18258
0 18260 7 1 2 49051 18259
0 18261 5 1 1 18260
0 18262 7 1 2 18231 18261
0 18263 5 1 1 18262
0 18264 7 1 2 51753 18263
0 18265 5 1 1 18264
0 18266 7 1 2 72614 70051
0 18267 7 1 2 69591 18266
0 18268 5 1 1 18267
0 18269 7 1 2 18265 18268
0 18270 5 1 1 18269
0 18271 7 1 2 54270 18270
0 18272 5 1 1 18271
0 18273 7 1 2 72276 68649
0 18274 5 1 1 18273
0 18275 7 1 2 51754 68444
0 18276 7 1 2 72220 18275
0 18277 5 1 1 18276
0 18278 7 1 2 18274 18277
0 18279 5 1 1 18278
0 18280 7 1 2 55744 18279
0 18281 5 1 1 18280
0 18282 7 1 2 72269 18281
0 18283 7 1 2 18272 18282
0 18284 5 1 1 18283
0 18285 7 1 2 54991 18284
0 18286 5 1 1 18285
0 18287 7 1 2 62558 71916
0 18288 5 1 1 18287
0 18289 7 1 2 63419 72240
0 18290 7 1 2 65769 18289
0 18291 5 1 1 18290
0 18292 7 1 2 18288 18291
0 18293 5 1 1 18292
0 18294 7 1 2 51303 18293
0 18295 5 1 1 18294
0 18296 7 1 2 66584 71347
0 18297 7 1 2 67667 18296
0 18298 5 1 1 18297
0 18299 7 1 2 18295 18298
0 18300 5 1 1 18299
0 18301 7 1 2 69980 18300
0 18302 5 1 1 18301
0 18303 7 1 2 49052 64984
0 18304 7 1 2 70068 18303
0 18305 5 1 1 18304
0 18306 7 1 2 18302 18305
0 18307 5 1 1 18306
0 18308 7 1 2 50050 18307
0 18309 5 1 1 18308
0 18310 7 1 2 72241 72471
0 18311 7 1 2 71435 18310
0 18312 5 1 1 18311
0 18313 7 1 2 18309 18312
0 18314 5 1 1 18313
0 18315 7 1 2 51566 55745
0 18316 7 1 2 18314 18315
0 18317 5 1 1 18316
0 18318 7 1 2 18286 18317
0 18319 5 1 1 18318
0 18320 7 1 2 56714 18319
0 18321 5 1 1 18320
0 18322 7 1 2 48154 70086
0 18323 5 1 1 18322
0 18324 7 1 2 58392 69796
0 18325 7 1 2 65837 18324
0 18326 5 1 1 18325
0 18327 7 1 2 18323 18326
0 18328 5 1 1 18327
0 18329 7 1 2 72478 18328
0 18330 5 1 1 18329
0 18331 7 1 2 63323 73799
0 18332 5 1 1 18331
0 18333 7 1 2 18330 18332
0 18334 5 1 1 18333
0 18335 7 1 2 49053 18334
0 18336 5 1 1 18335
0 18337 7 1 2 67039 66634
0 18338 7 3 2 50425 73669
0 18339 7 1 2 71892 74391
0 18340 7 1 2 18337 18339
0 18341 5 1 1 18340
0 18342 7 1 2 18336 18341
0 18343 5 1 1 18342
0 18344 7 1 2 51567 18343
0 18345 5 1 1 18344
0 18346 7 1 2 48155 65375
0 18347 5 3 1 18346
0 18348 7 1 2 71402 74394
0 18349 5 1 1 18348
0 18350 7 4 2 67614 72616
0 18351 5 1 1 74397
0 18352 7 1 2 55323 74398
0 18353 7 1 2 18349 18352
0 18354 5 1 1 18353
0 18355 7 1 2 18345 18354
0 18356 5 1 1 18355
0 18357 7 1 2 49201 18356
0 18358 5 1 1 18357
0 18359 7 3 2 49054 69419
0 18360 7 1 2 54619 74401
0 18361 5 2 1 18360
0 18362 7 2 2 73968 72248
0 18363 7 1 2 67275 66507
0 18364 7 1 2 74406 18363
0 18365 5 1 1 18364
0 18366 7 1 2 74404 18365
0 18367 5 1 1 18366
0 18368 7 1 2 47893 18367
0 18369 5 1 1 18368
0 18370 7 1 2 54021 74399
0 18371 5 1 1 18370
0 18372 7 1 2 57162 74402
0 18373 5 1 1 18372
0 18374 7 1 2 18371 18373
0 18375 5 1 1 18374
0 18376 7 1 2 54271 18375
0 18377 5 1 1 18376
0 18378 7 1 2 18369 18377
0 18379 5 1 1 18378
0 18380 7 1 2 55324 18379
0 18381 5 1 1 18380
0 18382 7 1 2 62723 68978
0 18383 7 1 2 72596 18382
0 18384 7 1 2 70087 18383
0 18385 5 1 1 18384
0 18386 7 1 2 18381 18385
0 18387 5 1 1 18386
0 18388 7 1 2 55746 18387
0 18389 5 1 1 18388
0 18390 7 2 2 68262 69917
0 18391 5 1 1 74408
0 18392 7 2 2 67615 69462
0 18393 7 1 2 49922 74410
0 18394 7 1 2 72263 18393
0 18395 5 1 1 18394
0 18396 7 1 2 18391 18395
0 18397 5 1 1 18396
0 18398 7 1 2 48741 18397
0 18399 5 1 1 18398
0 18400 7 6 2 67689 6956
0 18401 5 1 1 74412
0 18402 7 1 2 63670 71917
0 18403 7 1 2 69415 18402
0 18404 7 1 2 74413 18403
0 18405 5 1 1 18404
0 18406 7 1 2 18399 18405
0 18407 5 1 1 18406
0 18408 7 1 2 54620 18407
0 18409 5 1 1 18408
0 18410 7 1 2 18389 18409
0 18411 7 1 2 18358 18410
0 18412 5 1 1 18411
0 18413 7 1 2 55647 18412
0 18414 5 1 1 18413
0 18415 7 1 2 18321 18414
0 18416 7 1 2 18229 18415
0 18417 5 1 1 18416
0 18418 7 1 2 56077 18417
0 18419 5 1 1 18418
0 18420 7 2 2 60295 72221
0 18421 7 1 2 67554 74418
0 18422 5 1 1 18421
0 18423 7 1 2 72111 13837
0 18424 5 1 1 18423
0 18425 7 1 2 48742 18424
0 18426 5 1 1 18425
0 18427 7 1 2 18426 72836
0 18428 5 3 1 18427
0 18429 7 1 2 64595 67580
0 18430 7 1 2 74420 18429
0 18431 5 1 1 18430
0 18432 7 1 2 18422 18431
0 18433 5 1 1 18432
0 18434 7 1 2 57484 18433
0 18435 5 1 1 18434
0 18436 7 1 2 63048 67555
0 18437 7 1 2 72222 18436
0 18438 5 1 1 18437
0 18439 7 1 2 18435 18438
0 18440 5 1 1 18439
0 18441 7 1 2 55532 18440
0 18442 5 1 1 18441
0 18443 7 1 2 57596 67604
0 18444 5 1 1 18443
0 18445 7 1 2 64120 18444
0 18446 5 1 1 18445
0 18447 7 1 2 60296 67004
0 18448 5 1 1 18447
0 18449 7 1 2 18446 18448
0 18450 5 1 1 18449
0 18451 7 1 2 69569 18450
0 18452 5 1 1 18451
0 18453 7 1 2 60297 71378
0 18454 5 1 1 18453
0 18455 7 1 2 18452 18454
0 18456 5 1 1 18455
0 18457 7 1 2 72597 18456
0 18458 5 1 1 18457
0 18459 7 1 2 18442 18458
0 18460 5 1 1 18459
0 18461 7 1 2 54992 18460
0 18462 5 1 1 18461
0 18463 7 5 2 63287 58256
0 18464 5 1 1 74423
0 18465 7 1 2 49317 49734
0 18466 7 1 2 74321 18465
0 18467 7 1 2 74424 18466
0 18468 5 1 1 18467
0 18469 7 1 2 68441 18468
0 18470 5 1 1 18469
0 18471 7 1 2 55325 69570
0 18472 7 1 2 18470 18471
0 18473 5 1 1 18472
0 18474 7 1 2 49923 66396
0 18475 7 1 2 67606 18474
0 18476 5 1 1 18475
0 18477 7 1 2 18473 18476
0 18478 5 1 1 18477
0 18479 7 1 2 68263 18478
0 18480 5 1 1 18479
0 18481 7 1 2 67607 69600
0 18482 5 1 1 18481
0 18483 7 1 2 18482 68337
0 18484 5 1 1 18483
0 18485 7 1 2 50051 18484
0 18486 5 1 1 18485
0 18487 7 1 2 48939 71660
0 18488 5 1 1 18487
0 18489 7 1 2 18486 18488
0 18490 5 1 1 18489
0 18491 7 1 2 49055 18490
0 18492 5 1 1 18491
0 18493 7 2 2 48940 72303
0 18494 7 1 2 68333 74428
0 18495 5 1 1 18494
0 18496 7 1 2 18492 18495
0 18497 5 1 1 18496
0 18498 7 1 2 49735 18497
0 18499 5 1 1 18498
0 18500 7 1 2 63249 67422
0 18501 7 1 2 72209 18500
0 18502 7 1 2 70705 18501
0 18503 5 1 1 18502
0 18504 7 1 2 18499 18503
0 18505 5 1 1 18504
0 18506 7 1 2 48743 18505
0 18507 5 1 1 18506
0 18508 7 1 2 18480 18507
0 18509 7 1 2 18462 18508
0 18510 5 1 1 18509
0 18511 7 1 2 51755 18510
0 18512 5 1 1 18511
0 18513 7 1 2 67581 72277
0 18514 5 1 1 18513
0 18515 7 6 2 67942 74421
0 18516 7 1 2 62779 59545
0 18517 7 1 2 74430 18516
0 18518 5 1 1 18517
0 18519 7 1 2 18514 18518
0 18520 5 1 1 18519
0 18521 7 1 2 55326 18520
0 18522 5 1 1 18521
0 18523 7 1 2 57739 70030
0 18524 7 1 2 74419 18523
0 18525 5 1 1 18524
0 18526 7 1 2 18522 18525
0 18527 5 1 1 18526
0 18528 7 1 2 54993 18527
0 18529 5 1 1 18528
0 18530 7 1 2 58257 69797
0 18531 5 1 1 18530
0 18532 7 1 2 9174 18531
0 18533 5 1 1 18532
0 18534 7 1 2 59987 18533
0 18535 5 1 1 18534
0 18536 7 1 2 74352 18535
0 18537 5 1 1 18536
0 18538 7 1 2 68985 18537
0 18539 5 1 1 18538
0 18540 7 3 2 54621 70069
0 18541 7 1 2 60323 74436
0 18542 5 1 1 18541
0 18543 7 1 2 18539 18542
0 18544 5 1 1 18543
0 18545 7 1 2 50052 18544
0 18546 5 1 1 18545
0 18547 7 1 2 72472 74368
0 18548 5 1 1 18547
0 18549 7 1 2 18546 18548
0 18550 5 1 1 18549
0 18551 7 1 2 49056 18550
0 18552 5 1 1 18551
0 18553 7 1 2 65770 69366
0 18554 7 1 2 74373 18553
0 18555 5 1 1 18554
0 18556 7 1 2 18552 18555
0 18557 5 1 1 18556
0 18558 7 1 2 51568 18557
0 18559 5 1 1 18558
0 18560 7 1 2 18529 18559
0 18561 5 1 1 18560
0 18562 7 1 2 56078 18561
0 18563 5 1 1 18562
0 18564 7 1 2 68616 72617
0 18565 7 1 2 74325 18564
0 18566 5 1 1 18565
0 18567 7 3 2 53484 68979
0 18568 7 1 2 72598 74439
0 18569 7 1 2 64913 18568
0 18570 5 1 1 18569
0 18571 7 1 2 18566 18570
0 18572 5 1 1 18571
0 18573 7 1 2 48156 18572
0 18574 5 1 1 18573
0 18575 7 1 2 62724 74403
0 18576 5 1 1 18575
0 18577 7 1 2 18351 18576
0 18578 5 1 1 18577
0 18579 7 1 2 57485 18578
0 18580 5 1 1 18579
0 18581 7 1 2 59988 74400
0 18582 5 1 1 18581
0 18583 7 2 2 67546 71348
0 18584 7 1 2 69409 72482
0 18585 7 1 2 74442 18584
0 18586 5 1 1 18585
0 18587 7 1 2 18582 18586
0 18588 5 1 1 18587
0 18589 7 1 2 54622 18588
0 18590 5 1 1 18589
0 18591 7 1 2 18580 18590
0 18592 7 1 2 18574 18591
0 18593 5 1 1 18592
0 18594 7 1 2 55327 18593
0 18595 5 1 1 18594
0 18596 7 1 2 62559 60324
0 18597 7 1 2 74409 18596
0 18598 5 1 1 18597
0 18599 7 1 2 18595 18598
0 18600 5 1 1 18599
0 18601 7 1 2 55648 18600
0 18602 5 1 1 18601
0 18603 7 1 2 18563 18602
0 18604 7 1 2 18512 18603
0 18605 5 1 1 18604
0 18606 7 1 2 58604 18605
0 18607 5 1 1 18606
0 18608 7 1 2 65204 72854
0 18609 5 1 1 18608
0 18610 7 1 2 65458 60415
0 18611 5 1 1 18610
0 18612 7 3 2 66093 18611
0 18613 7 1 2 61715 70018
0 18614 7 1 2 74444 18613
0 18615 5 1 1 18614
0 18616 7 1 2 18609 18615
0 18617 5 1 1 18616
0 18618 7 1 2 50053 18617
0 18619 5 1 1 18618
0 18620 7 1 2 67024 74104
0 18621 7 1 2 74445 18620
0 18622 5 1 1 18621
0 18623 7 1 2 18619 18622
0 18624 5 1 1 18623
0 18625 7 1 2 49057 18624
0 18626 5 1 1 18625
0 18627 7 1 2 49736 71787
0 18628 7 1 2 72307 18627
0 18629 7 1 2 74446 18628
0 18630 5 1 1 18629
0 18631 7 1 2 18626 18630
0 18632 5 1 1 18631
0 18633 7 1 2 51756 18632
0 18634 5 1 1 18633
0 18635 7 1 2 63973 73946
0 18636 5 2 1 18635
0 18637 7 1 2 55328 74447
0 18638 7 1 2 72278 18637
0 18639 5 1 1 18638
0 18640 7 1 2 18634 18639
0 18641 5 1 1 18640
0 18642 7 1 2 54994 18641
0 18643 5 1 1 18642
0 18644 7 1 2 60349 70088
0 18645 5 1 1 18644
0 18646 7 1 2 18645 72163
0 18647 5 1 1 18646
0 18648 7 1 2 65205 18647
0 18649 5 1 1 18648
0 18650 7 3 2 51304 57824
0 18651 7 1 2 62560 60298
0 18652 7 1 2 74449 18651
0 18653 5 1 1 18652
0 18654 7 1 2 18649 18653
0 18655 5 1 1 18654
0 18656 7 1 2 68861 18655
0 18657 5 1 1 18656
0 18658 7 3 2 67943 70019
0 18659 7 2 2 63780 74452
0 18660 7 1 2 47894 74455
0 18661 5 1 1 18660
0 18662 7 1 2 18657 18661
0 18663 5 1 1 18662
0 18664 7 1 2 51011 18663
0 18665 5 1 1 18664
0 18666 7 5 2 51569 70070
0 18667 5 1 1 74457
0 18668 7 1 2 74458 71987
0 18669 5 1 1 18668
0 18670 7 1 2 18665 18669
0 18671 5 1 1 18670
0 18672 7 1 2 68264 18671
0 18673 5 1 1 18672
0 18674 7 1 2 68223 74369
0 18675 7 1 2 72866 18674
0 18676 5 1 1 18675
0 18677 7 1 2 18673 18676
0 18678 7 1 2 18643 18677
0 18679 5 1 1 18678
0 18680 7 1 2 55747 18679
0 18681 5 1 1 18680
0 18682 7 2 2 64809 74431
0 18683 5 1 1 74462
0 18684 7 1 2 69420 72031
0 18685 5 1 1 18684
0 18686 7 1 2 18683 18685
0 18687 5 2 1 18686
0 18688 7 1 2 57779 65825
0 18689 5 1 1 18688
0 18690 7 1 2 74464 18689
0 18691 5 1 1 18690
0 18692 7 1 2 62750 71935
0 18693 7 1 2 72279 18692
0 18694 5 1 1 18693
0 18695 7 1 2 18691 18694
0 18696 5 1 1 18695
0 18697 7 1 2 55329 18696
0 18698 5 1 1 18697
0 18699 7 4 2 47895 64149
0 18700 7 1 2 61857 72388
0 18701 7 1 2 74466 18700
0 18702 5 1 1 18701
0 18703 7 1 2 62600 18702
0 18704 5 1 1 18703
0 18705 7 1 2 68862 18704
0 18706 5 1 1 18705
0 18707 7 2 2 54995 74453
0 18708 7 2 2 54272 64858
0 18709 5 2 1 74472
0 18710 7 1 2 57597 74474
0 18711 5 2 1 18710
0 18712 7 1 2 74470 74476
0 18713 5 1 1 18712
0 18714 7 1 2 18706 18713
0 18715 5 1 1 18714
0 18716 7 1 2 51305 18715
0 18717 5 1 1 18716
0 18718 7 1 2 62725 2387
0 18719 5 2 1 18718
0 18720 7 1 2 64544 74478
0 18721 5 1 1 18720
0 18722 7 1 2 74459 18721
0 18723 5 1 1 18722
0 18724 7 1 2 18717 18723
0 18725 5 1 1 18724
0 18726 7 1 2 68265 18725
0 18727 5 1 1 18726
0 18728 7 3 2 63726 67944
0 18729 7 2 2 68224 74480
0 18730 7 1 2 70003 74483
0 18731 7 1 2 74477 18730
0 18732 5 1 1 18731
0 18733 7 1 2 18727 18732
0 18734 7 1 2 18698 18733
0 18735 5 1 1 18734
0 18736 7 1 2 55748 18735
0 18737 5 1 1 18736
0 18738 7 1 2 67164 71654
0 18739 7 2 2 74484 18738
0 18740 7 1 2 65453 74485
0 18741 5 1 1 18740
0 18742 7 1 2 65454 62599
0 18743 5 1 1 18742
0 18744 7 1 2 64709 63328
0 18745 7 1 2 66020 18744
0 18746 5 1 1 18745
0 18747 7 1 2 18743 18746
0 18748 5 1 1 18747
0 18749 7 1 2 72541 18748
0 18750 5 1 1 18749
0 18751 7 1 2 69571 71839
0 18752 5 1 1 18751
0 18753 7 2 2 72361 18752
0 18754 5 3 1 74487
0 18755 7 1 2 54996 74489
0 18756 5 1 1 18755
0 18757 7 1 2 59438 67457
0 18758 5 1 1 18757
0 18759 7 1 2 74490 18758
0 18760 5 1 1 18759
0 18761 7 1 2 67616 73583
0 18762 7 1 2 74336 18761
0 18763 5 1 1 18762
0 18764 7 1 2 18760 18763
0 18765 5 1 1 18764
0 18766 7 1 2 57486 18765
0 18767 5 1 1 18766
0 18768 7 1 2 18756 18767
0 18769 5 1 1 18768
0 18770 7 1 2 51757 18769
0 18771 5 1 1 18770
0 18772 7 1 2 18750 18771
0 18773 5 1 1 18772
0 18774 7 1 2 68266 18773
0 18775 5 1 1 18774
0 18776 7 1 2 18741 18775
0 18777 7 1 2 18737 18776
0 18778 5 1 1 18777
0 18779 7 1 2 54623 18778
0 18780 5 1 1 18779
0 18781 7 3 2 63573 67945
0 18782 7 1 2 57740 74492
0 18783 5 1 1 18782
0 18784 7 1 2 16629 18783
0 18785 5 1 1 18784
0 18786 7 1 2 48744 18785
0 18787 5 1 1 18786
0 18788 7 1 2 68827 72875
0 18789 5 1 1 18788
0 18790 7 1 2 67085 72416
0 18791 5 1 1 18790
0 18792 7 1 2 18789 18791
0 18793 7 1 2 18787 18792
0 18794 5 1 1 18793
0 18795 7 1 2 65206 18794
0 18796 5 1 1 18795
0 18797 7 1 2 63864 74471
0 18798 5 1 1 18797
0 18799 7 1 2 59546 68986
0 18800 7 1 2 71876 18799
0 18801 5 1 1 18800
0 18802 7 1 2 18798 18801
0 18803 7 1 2 18796 18802
0 18804 5 1 1 18803
0 18805 7 1 2 51306 18804
0 18806 5 1 1 18805
0 18807 7 1 2 64513 65689
0 18808 5 1 1 18807
0 18809 7 1 2 74460 18808
0 18810 5 1 1 18809
0 18811 7 1 2 18806 18810
0 18812 5 1 1 18811
0 18813 7 1 2 50054 18812
0 18814 5 1 1 18813
0 18815 7 2 2 61905 74493
0 18816 5 1 1 74495
0 18817 7 1 2 51307 74496
0 18818 5 1 1 18817
0 18819 7 1 2 8474 18818
0 18820 5 1 1 18819
0 18821 7 1 2 48157 18820
0 18822 5 1 1 18821
0 18823 7 2 2 58677 74494
0 18824 5 1 1 74497
0 18825 7 1 2 51308 74498
0 18826 5 1 1 18825
0 18827 7 1 2 18822 18826
0 18828 5 1 1 18827
0 18829 7 1 2 47896 18828
0 18830 5 1 1 18829
0 18831 7 2 2 61906 63406
0 18832 7 1 2 74481 74499
0 18833 5 1 1 18832
0 18834 7 1 2 18830 18833
0 18835 5 1 1 18834
0 18836 7 1 2 74357 18835
0 18837 5 1 1 18836
0 18838 7 1 2 18814 18837
0 18839 5 1 1 18838
0 18840 7 1 2 49058 18839
0 18841 5 1 1 18840
0 18842 7 1 2 67491 72249
0 18843 7 1 2 74467 18842
0 18844 5 1 1 18843
0 18845 7 1 2 74405 18844
0 18846 5 1 1 18845
0 18847 7 1 2 55649 18846
0 18848 5 1 1 18847
0 18849 7 1 2 72599 74468
0 18850 7 1 2 69995 18849
0 18851 5 1 1 18850
0 18852 7 1 2 18848 18851
0 18853 5 1 1 18852
0 18854 7 1 2 67588 18853
0 18855 5 1 1 18854
0 18856 7 1 2 65771 71704
0 18857 5 1 1 18856
0 18858 7 1 2 18816 18857
0 18859 5 1 1 18858
0 18860 7 1 2 48158 18859
0 18861 5 1 1 18860
0 18862 7 1 2 18824 18861
0 18863 5 1 1 18862
0 18864 7 1 2 47897 18863
0 18865 5 1 1 18864
0 18866 7 1 2 49737 60393
0 18867 7 1 2 69936 18866
0 18868 5 1 1 18867
0 18869 7 1 2 18865 18868
0 18870 5 1 1 18869
0 18871 7 1 2 51309 72308
0 18872 7 1 2 18870 18871
0 18873 5 1 1 18872
0 18874 7 1 2 18855 18873
0 18875 7 1 2 18841 18874
0 18876 5 1 1 18875
0 18877 7 1 2 59579 18876
0 18878 5 1 1 18877
0 18879 7 1 2 57844 4636
0 18880 5 1 1 18879
0 18881 7 1 2 48159 18880
0 18882 5 1 1 18881
0 18883 7 1 2 49119 57770
0 18884 5 1 1 18883
0 18885 7 1 2 18882 18884
0 18886 5 1 1 18885
0 18887 7 1 2 53904 18886
0 18888 5 1 1 18887
0 18889 7 1 2 65677 18888
0 18890 5 2 1 18889
0 18891 7 1 2 74486 74501
0 18892 5 1 1 18891
0 18893 7 1 2 48160 60394
0 18894 5 1 1 18893
0 18895 7 2 2 57598 18894
0 18896 5 2 1 74503
0 18897 7 1 2 51012 74504
0 18898 5 1 1 18897
0 18899 7 1 2 71861 18898
0 18900 5 1 1 18899
0 18901 7 1 2 72417 18900
0 18902 5 1 1 18901
0 18903 7 1 2 62561 18902
0 18904 5 1 1 18903
0 18905 7 1 2 64810 74454
0 18906 7 1 2 74502 18905
0 18907 5 1 1 18906
0 18908 7 1 2 18904 18907
0 18909 5 1 1 18908
0 18910 7 1 2 51310 18909
0 18911 5 1 1 18910
0 18912 7 1 2 65197 3152
0 18913 5 1 1 18912
0 18914 7 1 2 54997 18913
0 18915 5 1 1 18914
0 18916 7 2 2 64988 61389
0 18917 7 2 2 49318 59503
0 18918 5 3 1 74509
0 18919 7 1 2 74507 74510
0 18920 5 1 1 18919
0 18921 7 1 2 18915 18920
0 18922 5 1 1 18921
0 18923 7 1 2 49202 18922
0 18924 5 1 1 18923
0 18925 7 3 2 47898 65207
0 18926 5 1 1 74514
0 18927 7 1 2 57599 18926
0 18928 5 1 1 18927
0 18929 7 1 2 54998 18928
0 18930 5 1 1 18929
0 18931 7 1 2 18924 18930
0 18932 5 1 1 18931
0 18933 7 1 2 74461 18932
0 18934 5 1 1 18933
0 18935 7 1 2 18911 18934
0 18936 5 1 1 18935
0 18937 7 1 2 68267 18936
0 18938 5 1 1 18937
0 18939 7 1 2 18892 18938
0 18940 7 1 2 18878 18939
0 18941 7 1 2 18780 18940
0 18942 7 1 2 18681 18941
0 18943 7 1 2 74505 69983
0 18944 5 1 1 18943
0 18945 7 1 2 59439 59556
0 18946 5 1 1 18945
0 18947 7 1 2 57487 66337
0 18948 5 1 1 18947
0 18949 7 1 2 51013 18948
0 18950 5 1 1 18949
0 18951 7 1 2 18946 18950
0 18952 5 1 1 18951
0 18953 7 3 2 54999 61554
0 18954 5 1 1 74517
0 18955 7 1 2 48161 74518
0 18956 5 1 1 18955
0 18957 7 2 2 47899 58134
0 18958 5 1 1 74520
0 18959 7 1 2 57488 66154
0 18960 7 1 2 74521 18959
0 18961 5 1 1 18960
0 18962 7 1 2 18956 18961
0 18963 7 1 2 18952 18962
0 18964 5 2 1 18963
0 18965 7 1 2 69996 74522
0 18966 5 1 1 18965
0 18967 7 1 2 18944 18966
0 18968 5 1 1 18967
0 18969 7 1 2 51570 18968
0 18970 5 1 1 18969
0 18971 7 1 2 66743 71900
0 18972 7 1 2 73986 18971
0 18973 5 1 1 18972
0 18974 7 1 2 72805 18973
0 18975 5 1 1 18974
0 18976 7 1 2 67946 18975
0 18977 5 1 1 18976
0 18978 7 1 2 18970 18977
0 18979 5 1 1 18978
0 18980 7 1 2 50055 18979
0 18981 5 1 1 18980
0 18982 7 1 2 64863 63355
0 18983 7 1 2 74036 69960
0 18984 7 1 2 18982 18983
0 18985 5 1 1 18984
0 18986 7 1 2 18981 18985
0 18987 5 1 1 18986
0 18988 7 1 2 49059 18987
0 18989 5 1 1 18988
0 18990 7 4 2 47900 59434
0 18991 5 1 1 74524
0 18992 7 1 2 54273 59820
0 18993 5 1 1 18992
0 18994 7 1 2 18991 18993
0 18995 5 1 1 18994
0 18996 7 1 2 74465 18995
0 18997 5 1 1 18996
0 18998 7 1 2 71918 74119
0 18999 7 1 2 71705 18998
0 19000 5 1 1 18999
0 19001 7 1 2 18997 19000
0 19002 5 1 1 19001
0 19003 7 1 2 60299 19002
0 19004 5 1 1 19003
0 19005 7 3 2 53791 72069
0 19006 5 1 1 74528
0 19007 7 1 2 74523 74529
0 19008 5 1 1 19007
0 19009 7 2 2 63250 72384
0 19010 7 1 2 74380 72437
0 19011 7 1 2 74531 19010
0 19012 5 1 1 19011
0 19013 7 1 2 19008 19012
0 19014 5 1 1 19013
0 19015 7 1 2 74348 19014
0 19016 5 1 1 19015
0 19017 7 1 2 19004 19016
0 19018 7 1 2 18989 19017
0 19019 5 1 1 19018
0 19020 7 1 2 54624 19019
0 19021 5 1 1 19020
0 19022 7 2 2 52121 59448
0 19023 5 2 1 74533
0 19024 7 1 2 50190 74534
0 19025 5 1 1 19024
0 19026 7 1 2 59435 19025
0 19027 5 1 1 19026
0 19028 7 1 2 48162 70715
0 19029 5 2 1 19028
0 19030 7 1 2 67433 74537
0 19031 7 1 2 19027 19030
0 19032 5 1 1 19031
0 19033 7 1 2 69984 19032
0 19034 5 1 1 19033
0 19035 7 1 2 65506 60460
0 19036 7 1 2 69991 19035
0 19037 5 1 1 19036
0 19038 7 1 2 19034 19037
0 19039 5 1 1 19038
0 19040 7 1 2 57489 19039
0 19041 5 1 1 19040
0 19042 7 1 2 69523 69752
0 19043 5 1 1 19042
0 19044 7 1 2 19041 19043
0 19045 5 1 1 19044
0 19046 7 1 2 51571 19045
0 19047 5 1 1 19046
0 19048 7 1 2 59137 67947
0 19049 7 2 2 60461 19048
0 19050 7 1 2 70020 74539
0 19051 5 1 1 19050
0 19052 7 1 2 19047 19051
0 19053 5 1 1 19052
0 19054 7 1 2 50056 19053
0 19055 5 1 1 19054
0 19056 7 1 2 70004 74540
0 19057 5 1 1 19056
0 19058 7 1 2 19055 19057
0 19059 5 1 1 19058
0 19060 7 1 2 49060 19059
0 19061 5 1 1 19060
0 19062 7 2 2 67031 67833
0 19063 7 1 2 60462 74541
0 19064 7 1 2 72506 19063
0 19065 5 1 1 19064
0 19066 7 1 2 19061 19065
0 19067 7 1 2 19021 19066
0 19068 5 1 1 19067
0 19069 7 1 2 55330 19068
0 19070 5 1 1 19069
0 19071 7 1 2 50426 58140
0 19072 5 1 1 19071
0 19073 7 1 2 65894 68078
0 19074 5 1 1 19073
0 19075 7 1 2 51014 19074
0 19076 5 1 1 19075
0 19077 7 1 2 72280 19076
0 19078 5 1 1 19077
0 19079 7 1 2 58855 74463
0 19080 5 1 1 19079
0 19081 7 1 2 55650 69416
0 19082 7 1 2 74443 19081
0 19083 5 1 1 19082
0 19084 7 1 2 19080 19083
0 19085 5 1 1 19084
0 19086 7 1 2 60300 19085
0 19087 5 1 1 19086
0 19088 7 1 2 19078 19087
0 19089 5 1 1 19088
0 19090 7 1 2 55331 19089
0 19091 5 1 1 19090
0 19092 7 1 2 57490 72265
0 19093 5 1 1 19092
0 19094 7 1 2 19091 19093
0 19095 5 1 1 19094
0 19096 7 1 2 54625 19095
0 19097 5 1 1 19096
0 19098 7 1 2 55000 70071
0 19099 5 1 1 19098
0 19100 7 1 2 72392 19099
0 19101 5 1 1 19100
0 19102 7 1 2 67662 19101
0 19103 5 1 1 19102
0 19104 7 1 2 64811 68079
0 19105 7 1 2 70021 70031
0 19106 7 1 2 19104 19105
0 19107 5 1 1 19106
0 19108 7 1 2 19103 19107
0 19109 5 1 1 19108
0 19110 7 1 2 50057 19109
0 19111 5 1 1 19110
0 19112 7 1 2 64539 74482
0 19113 7 2 2 48745 60925
0 19114 5 1 1 74543
0 19115 7 4 2 48941 68773
0 19116 7 1 2 74544 74545
0 19117 7 1 2 19112 19116
0 19118 5 1 1 19117
0 19119 7 1 2 19111 19118
0 19120 5 1 1 19119
0 19121 7 1 2 49061 19120
0 19122 5 1 1 19121
0 19123 7 1 2 51758 58148
0 19124 7 1 2 64255 19123
0 19125 7 1 2 74429 19124
0 19126 7 1 2 71682 19125
0 19127 5 1 1 19126
0 19128 7 1 2 19122 19127
0 19129 7 1 2 19097 19128
0 19130 5 1 1 19129
0 19131 7 1 2 19072 19130
0 19132 5 1 1 19131
0 19133 7 1 2 19070 19132
0 19134 7 1 2 18942 19133
0 19135 7 1 2 18607 19134
0 19136 7 1 2 18419 19135
0 19137 5 1 1 19136
0 19138 7 1 2 56549 19137
0 19139 5 1 1 19138
0 19140 7 1 2 18049 19139
0 19141 7 1 2 17125 19140
0 19142 5 1 1 19141
0 19143 7 1 2 56347 19142
0 19144 5 1 1 19143
0 19145 7 1 2 16081 19144
0 19146 7 2 2 49319 59719
0 19147 5 1 1 74549
0 19148 7 2 2 49320 62050
0 19149 5 1 1 74551
0 19150 7 1 2 59728 58486
0 19151 7 1 2 19149 19150
0 19152 5 1 1 19151
0 19153 7 1 2 48369 19152
0 19154 5 1 1 19153
0 19155 7 1 2 19147 19154
0 19156 5 1 1 19155
0 19157 7 1 2 60195 72047
0 19158 7 1 2 72255 19157
0 19159 5 1 1 19158
0 19160 7 1 2 72253 19159
0 19161 5 1 1 19160
0 19162 7 1 2 49062 19161
0 19163 5 1 1 19162
0 19164 7 1 2 67120 68526
0 19165 7 1 2 67514 19164
0 19166 7 1 2 74392 19165
0 19167 5 1 1 19166
0 19168 7 1 2 19163 19167
0 19169 5 1 1 19168
0 19170 7 1 2 51572 19169
0 19171 5 1 1 19170
0 19172 7 1 2 72618 70052
0 19173 5 1 1 19172
0 19174 7 1 2 19171 19173
0 19175 5 1 1 19174
0 19176 7 1 2 19156 19175
0 19177 5 1 1 19176
0 19178 7 2 2 57491 68581
0 19179 7 1 2 74553 70915
0 19180 5 1 1 19179
0 19181 7 1 2 65704 74110
0 19182 5 1 1 19181
0 19183 7 1 2 19180 19182
0 19184 5 1 1 19183
0 19185 7 1 2 74358 19184
0 19186 5 1 1 19185
0 19187 7 2 2 63165 66471
0 19188 5 1 1 74555
0 19189 7 2 2 56715 74337
0 19190 5 1 1 74557
0 19191 7 1 2 57492 74558
0 19192 5 1 1 19191
0 19193 7 1 2 19188 19192
0 19194 5 1 1 19193
0 19195 7 1 2 54274 19194
0 19196 5 1 1 19195
0 19197 7 1 2 66846 74338
0 19198 5 1 1 19197
0 19199 7 1 2 19196 19198
0 19200 5 1 1 19199
0 19201 7 1 2 50058 19200
0 19202 5 1 1 19201
0 19203 7 1 2 19186 19202
0 19204 5 1 1 19203
0 19205 7 1 2 58393 19204
0 19206 5 1 1 19205
0 19207 7 1 2 62912 72511
0 19208 5 1 1 19207
0 19209 7 1 2 12210 19208
0 19210 5 1 1 19209
0 19211 7 1 2 59263 67556
0 19212 7 1 2 19210 19211
0 19213 5 1 1 19212
0 19214 7 1 2 19206 19213
0 19215 5 1 1 19214
0 19216 7 1 2 49063 19215
0 19217 5 1 1 19216
0 19218 7 1 2 59420 61874
0 19219 5 1 1 19218
0 19220 7 1 2 48163 19219
0 19221 5 1 1 19220
0 19222 7 1 2 59410 19221
0 19223 5 2 1 19222
0 19224 7 1 2 74554 74559
0 19225 5 1 1 19224
0 19226 7 1 2 69798 69225
0 19227 5 1 1 19226
0 19228 7 1 2 19225 19227
0 19229 5 1 1 19228
0 19230 7 1 2 72309 19229
0 19231 5 1 1 19230
0 19232 7 1 2 19217 19231
0 19233 5 1 1 19232
0 19234 7 1 2 55533 19233
0 19235 5 1 1 19234
0 19236 7 1 2 74120 69949
0 19237 7 1 2 72855 19236
0 19238 5 1 1 19237
0 19239 7 1 2 19235 19238
0 19240 5 1 1 19239
0 19241 7 1 2 51759 19240
0 19242 5 1 1 19241
0 19243 7 1 2 19177 19242
0 19244 5 1 1 19243
0 19245 7 1 2 47901 19244
0 19246 5 1 1 19245
0 19247 7 1 2 62562 67088
0 19248 5 1 1 19247
0 19249 7 1 2 72857 19248
0 19250 5 1 1 19249
0 19251 7 1 2 50059 19250
0 19252 5 1 1 19251
0 19253 7 1 2 69900 72810
0 19254 5 1 1 19253
0 19255 7 1 2 19252 19254
0 19256 5 3 1 19255
0 19257 7 1 2 49064 74561
0 19258 5 1 1 19257
0 19259 7 2 2 74371 72811
0 19260 7 1 2 66420 74564
0 19261 5 1 1 19260
0 19262 7 1 2 19258 19261
0 19263 5 4 1 19262
0 19264 7 3 2 53085 58425
0 19265 7 1 2 50427 74570
0 19266 5 1 1 19265
0 19267 7 1 2 74566 19266
0 19268 5 1 1 19267
0 19269 7 2 2 60057 71943
0 19270 7 2 2 48164 58605
0 19271 5 2 1 74575
0 19272 7 1 2 58294 74577
0 19273 5 8 1 19272
0 19274 7 1 2 74573 74579
0 19275 7 1 2 72223 19274
0 19276 5 1 1 19275
0 19277 7 1 2 19268 19276
0 19278 5 1 1 19277
0 19279 7 1 2 51760 19278
0 19280 5 1 1 19279
0 19281 7 2 2 56716 71349
0 19282 7 1 2 74381 74587
0 19283 5 1 1 19282
0 19284 7 3 2 48165 60196
0 19285 5 1 1 74589
0 19286 7 1 2 49203 74590
0 19287 7 1 2 71392 19286
0 19288 5 1 1 19287
0 19289 7 1 2 19283 19288
0 19290 5 1 1 19289
0 19291 7 1 2 56903 67477
0 19292 7 1 2 72291 19291
0 19293 7 1 2 19290 19292
0 19294 5 1 1 19293
0 19295 7 1 2 19280 19294
0 19296 5 1 1 19295
0 19297 7 1 2 48370 19296
0 19298 5 1 1 19297
0 19299 7 2 2 49321 65376
0 19300 5 1 1 74592
0 19301 7 1 2 61864 19300
0 19302 5 2 1 19301
0 19303 7 1 2 67948 74556
0 19304 5 1 1 19303
0 19305 7 1 2 18667 19304
0 19306 5 1 1 19305
0 19307 7 1 2 74594 19306
0 19308 5 1 1 19307
0 19309 7 1 2 67820 68863
0 19310 5 1 1 19309
0 19311 7 1 2 19308 19310
0 19312 5 1 1 19311
0 19313 7 1 2 50060 19312
0 19314 5 1 1 19313
0 19315 7 2 2 72055 74595
0 19316 7 3 2 73800 71872
0 19317 5 1 1 74598
0 19318 7 1 2 74596 74599
0 19319 5 1 1 19318
0 19320 7 1 2 19314 19319
0 19321 5 1 1 19320
0 19322 7 1 2 49065 19321
0 19323 5 1 1 19322
0 19324 7 1 2 72870 71380
0 19325 5 1 1 19324
0 19326 7 1 2 67032 69904
0 19327 5 1 1 19326
0 19328 7 1 2 19325 19327
0 19329 5 1 1 19328
0 19330 7 1 2 55651 19329
0 19331 5 1 1 19330
0 19332 7 1 2 69175 72251
0 19333 5 1 1 19332
0 19334 7 1 2 19331 19333
0 19335 5 2 1 19334
0 19336 7 2 2 57600 71403
0 19337 5 1 1 74603
0 19338 7 2 2 62446 19337
0 19339 7 1 2 54275 74605
0 19340 5 1 1 19339
0 19341 7 2 2 49120 62457
0 19342 7 1 2 61660 74607
0 19343 5 1 1 19342
0 19344 7 1 2 19340 19343
0 19345 5 1 1 19344
0 19346 7 1 2 74601 19345
0 19347 5 1 1 19346
0 19348 7 1 2 72224 71815
0 19349 5 1 1 19348
0 19350 7 1 2 72201 19349
0 19351 5 4 1 19350
0 19352 7 1 2 63768 74609
0 19353 5 1 1 19352
0 19354 7 1 2 74565 74597
0 19355 5 1 1 19354
0 19356 7 1 2 19353 19355
0 19357 7 1 2 19347 19356
0 19358 7 1 2 19323 19357
0 19359 7 1 2 19298 19358
0 19360 7 1 2 19246 19359
0 19361 5 1 1 19360
0 19362 7 1 2 54626 19361
0 19363 5 1 1 19362
0 19364 7 1 2 66639 74432
0 19365 5 1 1 19364
0 19366 7 3 2 59808 64472
0 19367 7 2 2 54022 74613
0 19368 7 1 2 72281 74616
0 19369 5 1 1 19368
0 19370 7 1 2 19365 19369
0 19371 5 1 1 19370
0 19372 7 1 2 55332 19371
0 19373 5 1 1 19372
0 19374 7 1 2 66702 69379
0 19375 5 1 1 19374
0 19376 7 1 2 69826 19375
0 19377 5 1 1 19376
0 19378 7 1 2 71393 19377
0 19379 5 1 1 19378
0 19380 7 1 2 74112 72847
0 19381 5 1 1 19380
0 19382 7 1 2 19379 19381
0 19383 5 1 1 19382
0 19384 7 1 2 74190 19383
0 19385 5 1 1 19384
0 19386 7 1 2 72270 19385
0 19387 5 1 1 19386
0 19388 7 1 2 48371 19387
0 19389 5 1 1 19388
0 19390 7 1 2 49322 70072
0 19391 5 1 1 19390
0 19392 7 1 2 68551 72495
0 19393 7 1 2 68303 19392
0 19394 7 1 2 64921 19393
0 19395 5 1 1 19394
0 19396 7 1 2 19391 19395
0 19397 5 1 1 19396
0 19398 7 1 2 72600 19397
0 19399 5 1 1 19398
0 19400 7 1 2 19389 19399
0 19401 7 1 2 19373 19400
0 19402 5 1 1 19401
0 19403 7 1 2 49204 19402
0 19404 5 1 1 19403
0 19405 7 1 2 56079 74567
0 19406 5 1 1 19405
0 19407 7 2 2 74151 72225
0 19408 5 1 1 74618
0 19409 7 1 2 19406 19408
0 19410 5 1 1 19409
0 19411 7 1 2 51761 62726
0 19412 7 1 2 19410 19411
0 19413 5 1 1 19412
0 19414 7 1 2 19404 19413
0 19415 5 1 1 19414
0 19416 7 1 2 48166 19415
0 19417 5 1 1 19416
0 19418 7 1 2 59587 74602
0 19419 5 1 1 19418
0 19420 7 1 2 51762 74568
0 19421 5 1 1 19420
0 19422 7 1 2 19419 19421
0 19423 5 1 1 19422
0 19424 7 1 2 54627 19423
0 19425 5 1 1 19424
0 19426 7 1 2 47902 74610
0 19427 5 1 1 19426
0 19428 7 1 2 19425 19427
0 19429 5 1 1 19428
0 19430 7 1 2 61699 19429
0 19431 5 1 1 19430
0 19432 7 1 2 61810 74569
0 19433 5 1 1 19432
0 19434 7 1 2 61804 74619
0 19435 5 1 1 19434
0 19436 7 1 2 19433 19435
0 19437 5 1 1 19436
0 19438 7 1 2 51763 19437
0 19439 5 1 1 19438
0 19440 7 1 2 19431 19439
0 19441 7 1 2 19417 19440
0 19442 5 1 1 19441
0 19443 7 1 2 54276 19442
0 19444 5 1 1 19443
0 19445 7 1 2 60197 68828
0 19446 7 2 2 69690 19445
0 19447 5 1 1 74620
0 19448 7 1 2 57493 74621
0 19449 5 1 1 19448
0 19450 7 1 2 51764 69901
0 19451 7 1 2 74617 19450
0 19452 5 1 1 19451
0 19453 7 1 2 19449 19452
0 19454 5 1 1 19453
0 19455 7 1 2 56717 19454
0 19456 5 1 1 19455
0 19457 7 1 2 69776 8486
0 19458 5 1 1 19457
0 19459 7 1 2 47903 19458
0 19460 5 2 1 19459
0 19461 7 1 2 74622 72167
0 19462 5 1 1 19461
0 19463 7 1 2 57163 19462
0 19464 5 1 1 19463
0 19465 7 1 2 17377 19464
0 19466 5 1 1 19465
0 19467 7 1 2 68906 19466
0 19468 5 1 1 19467
0 19469 7 1 2 19456 19468
0 19470 5 1 1 19469
0 19471 7 1 2 72812 19470
0 19472 5 1 1 19471
0 19473 7 1 2 51311 64945
0 19474 5 1 1 19473
0 19475 7 1 2 57164 73748
0 19476 5 1 1 19475
0 19477 7 1 2 19474 19476
0 19478 5 1 1 19477
0 19479 7 1 2 69015 19478
0 19480 5 1 1 19479
0 19481 7 2 2 62563 64759
0 19482 5 1 1 74624
0 19483 7 1 2 62913 56718
0 19484 5 1 1 19483
0 19485 7 1 2 19482 19484
0 19486 5 1 1 19485
0 19487 7 1 2 69572 19486
0 19488 5 1 1 19487
0 19489 7 1 2 56719 69618
0 19490 5 1 1 19489
0 19491 7 1 2 19488 19490
0 19492 5 1 1 19491
0 19493 7 1 2 68684 19492
0 19494 5 1 1 19493
0 19495 7 1 2 19480 19494
0 19496 5 1 1 19495
0 19497 7 1 2 54023 19496
0 19498 5 1 1 19497
0 19499 7 1 2 57165 74437
0 19500 5 1 1 19499
0 19501 7 1 2 62564 72399
0 19502 5 1 1 19501
0 19503 7 1 2 19500 19502
0 19504 7 1 2 19498 19503
0 19505 5 1 1 19504
0 19506 7 1 2 47904 19505
0 19507 5 1 1 19506
0 19508 7 1 2 57166 70073
0 19509 5 1 1 19508
0 19510 7 1 2 52614 2785
0 19511 5 1 1 19510
0 19512 7 1 2 69573 72043
0 19513 7 1 2 19511 19512
0 19514 5 1 1 19513
0 19515 7 1 2 12971 19514
0 19516 5 1 1 19515
0 19517 7 1 2 51765 19516
0 19518 5 1 1 19517
0 19519 7 1 2 67525 68552
0 19520 7 1 2 66621 19519
0 19521 5 1 1 19520
0 19522 7 1 2 19518 19521
0 19523 5 1 1 19522
0 19524 7 1 2 56720 19523
0 19525 5 1 1 19524
0 19526 7 1 2 19509 19525
0 19527 5 1 1 19526
0 19528 7 1 2 57494 19527
0 19529 5 1 1 19528
0 19530 7 1 2 69524 69852
0 19531 5 1 1 19530
0 19532 7 1 2 19529 19531
0 19533 7 1 2 19507 19532
0 19534 5 1 1 19533
0 19535 7 1 2 51573 19534
0 19536 5 1 1 19535
0 19537 7 1 2 64492 74339
0 19538 5 1 1 19537
0 19539 7 1 2 62565 66472
0 19540 7 1 2 61836 19539
0 19541 7 1 2 74614 19540
0 19542 5 1 1 19541
0 19543 7 1 2 19538 19542
0 19544 5 1 1 19543
0 19545 7 3 2 51766 56904
0 19546 7 1 2 55534 74626
0 19547 7 1 2 19544 19546
0 19548 5 1 1 19547
0 19549 7 1 2 19536 19548
0 19550 5 1 1 19549
0 19551 7 1 2 50061 19550
0 19552 5 1 1 19551
0 19553 7 1 2 19472 19552
0 19554 5 1 1 19553
0 19555 7 1 2 49066 19554
0 19556 5 1 1 19555
0 19557 7 1 2 48746 69778
0 19558 5 1 1 19557
0 19559 7 1 2 68793 12906
0 19560 7 1 2 19558 19559
0 19561 5 1 1 19560
0 19562 7 1 2 47905 19561
0 19563 5 1 1 19562
0 19564 7 1 2 19190 19563
0 19565 5 1 1 19564
0 19566 7 1 2 50062 19565
0 19567 5 1 1 19566
0 19568 7 1 2 56721 68582
0 19569 5 2 1 19568
0 19570 7 1 2 74623 74629
0 19571 5 1 1 19570
0 19572 7 1 2 74359 19571
0 19573 5 1 1 19572
0 19574 7 1 2 19567 19573
0 19575 5 1 1 19574
0 19576 7 1 2 49067 19575
0 19577 5 1 1 19576
0 19578 7 1 2 47906 67690
0 19579 7 1 2 72044 19578
0 19580 5 1 1 19579
0 19581 7 1 2 74630 19580
0 19582 5 1 1 19581
0 19583 7 1 2 72310 19582
0 19584 5 1 1 19583
0 19585 7 1 2 19577 19584
0 19586 5 1 1 19585
0 19587 7 1 2 74627 19586
0 19588 5 1 1 19587
0 19589 7 2 2 48167 72012
0 19590 7 6 2 48747 54024
0 19591 5 1 1 74633
0 19592 7 1 2 57741 74634
0 19593 7 1 2 74631 19592
0 19594 7 1 2 74407 19593
0 19595 5 1 1 19594
0 19596 7 1 2 19588 19595
0 19597 5 1 1 19596
0 19598 7 1 2 55535 19597
0 19599 5 1 1 19598
0 19600 7 1 2 62755 69833
0 19601 5 1 1 19600
0 19602 7 1 2 63981 65821
0 19603 7 1 2 69997 19602
0 19604 5 1 1 19603
0 19605 7 1 2 19601 19604
0 19606 5 1 1 19605
0 19607 7 1 2 55333 19606
0 19608 5 1 1 19607
0 19609 7 1 2 66786 72496
0 19610 7 1 2 69016 19609
0 19611 5 1 1 19610
0 19612 7 1 2 9155 19611
0 19613 5 1 1 19612
0 19614 7 1 2 57742 19613
0 19615 5 1 1 19614
0 19616 7 1 2 19608 19615
0 19617 5 1 1 19616
0 19618 7 1 2 72601 19617
0 19619 5 1 1 19618
0 19620 7 1 2 19599 19619
0 19621 5 1 1 19620
0 19622 7 1 2 56080 19621
0 19623 5 1 1 19622
0 19624 7 1 2 70046 72041
0 19625 5 1 1 19624
0 19626 7 2 2 69303 74316
0 19627 5 1 1 74639
0 19628 7 1 2 19447 19627
0 19629 5 1 1 19628
0 19630 7 1 2 50063 56905
0 19631 7 1 2 19629 19630
0 19632 5 1 1 19631
0 19633 7 1 2 19625 19632
0 19634 5 1 1 19633
0 19635 7 1 2 57495 19634
0 19636 5 1 1 19635
0 19637 7 1 2 66973 72373
0 19638 7 1 2 74640 19637
0 19639 5 1 1 19638
0 19640 7 1 2 19636 19639
0 19641 5 1 1 19640
0 19642 7 1 2 56722 19641
0 19643 5 1 1 19642
0 19644 7 3 2 51767 69447
0 19645 7 1 2 57851 74641
0 19646 5 1 1 19645
0 19647 7 1 2 19006 19646
0 19648 5 1 1 19647
0 19649 7 1 2 47907 19648
0 19650 5 1 1 19649
0 19651 7 1 2 59264 74642
0 19652 5 1 1 19651
0 19653 7 1 2 19650 19652
0 19654 5 1 1 19653
0 19655 7 1 2 56906 19654
0 19656 5 1 1 19655
0 19657 7 1 2 49738 69920
0 19658 7 1 2 65895 19657
0 19659 7 1 2 69972 19658
0 19660 5 1 1 19659
0 19661 7 1 2 19656 19660
0 19662 5 1 1 19661
0 19663 7 1 2 55334 19662
0 19664 5 1 1 19663
0 19665 7 1 2 69169 68784
0 19666 7 1 2 64493 19665
0 19667 5 1 1 19666
0 19668 7 1 2 19664 19667
0 19669 5 1 1 19668
0 19670 7 1 2 67834 19669
0 19671 5 1 1 19670
0 19672 7 1 2 19643 19671
0 19673 5 1 1 19672
0 19674 7 1 2 65630 19673
0 19675 5 1 1 19674
0 19676 7 1 2 19623 19675
0 19677 7 1 2 19556 19676
0 19678 7 1 2 19444 19677
0 19679 5 1 1 19678
0 19680 7 1 2 55749 19679
0 19681 5 1 1 19680
0 19682 7 1 2 64073 69601
0 19683 5 1 1 19682
0 19684 7 1 2 13119 19683
0 19685 5 1 1 19684
0 19686 7 1 2 64121 19685
0 19687 5 1 1 19686
0 19688 7 1 2 72858 19687
0 19689 5 1 1 19688
0 19690 7 1 2 51768 19689
0 19691 5 1 1 19690
0 19692 7 1 2 59504 72292
0 19693 7 1 2 69096 19692
0 19694 5 1 1 19693
0 19695 7 1 2 19691 19694
0 19696 5 1 1 19695
0 19697 7 1 2 50064 19696
0 19698 5 1 1 19697
0 19699 7 1 2 69304 74600
0 19700 5 1 1 19699
0 19701 7 1 2 19698 19700
0 19702 5 1 1 19701
0 19703 7 1 2 56081 19702
0 19704 5 1 1 19703
0 19705 7 1 2 47908 69068
0 19706 7 1 2 74562 19705
0 19707 5 1 1 19706
0 19708 7 1 2 19704 19707
0 19709 5 1 1 19708
0 19710 7 1 2 54628 19709
0 19711 5 1 1 19710
0 19712 7 1 2 70100 69481
0 19713 5 1 1 19712
0 19714 7 1 2 57496 74198
0 19715 7 1 2 74563 19714
0 19716 5 1 1 19715
0 19717 7 1 2 19713 19716
0 19718 5 1 1 19717
0 19719 7 1 2 51769 19718
0 19720 5 1 1 19719
0 19721 7 1 2 51574 74366
0 19722 7 1 2 72395 19721
0 19723 5 1 1 19722
0 19724 7 1 2 19720 19723
0 19725 7 1 2 19711 19724
0 19726 5 1 1 19725
0 19727 7 1 2 49068 19726
0 19728 5 1 1 19727
0 19729 7 1 2 57002 74214
0 19730 5 1 1 19729
0 19731 7 1 2 74530 19730
0 19732 5 1 1 19731
0 19733 7 1 2 58717 59535
0 19734 5 1 1 19733
0 19735 7 1 2 47909 19734
0 19736 5 1 1 19735
0 19737 7 1 2 64065 19736
0 19738 5 1 1 19737
0 19739 7 1 2 56907 74643
0 19740 7 1 2 19738 19739
0 19741 5 1 1 19740
0 19742 7 1 2 19732 19741
0 19743 5 1 1 19742
0 19744 7 1 2 55335 74349
0 19745 7 1 2 19743 19744
0 19746 5 1 1 19745
0 19747 7 1 2 59520 74611
0 19748 5 1 1 19747
0 19749 7 1 2 19746 19748
0 19750 7 1 2 19728 19749
0 19751 5 1 1 19750
0 19752 7 1 2 61700 19751
0 19753 5 1 1 19752
0 19754 7 1 2 68762 71352
0 19755 5 1 1 19754
0 19756 7 2 2 53905 66234
0 19757 7 1 2 65174 74644
0 19758 7 1 2 74433 19757
0 19759 5 1 1 19758
0 19760 7 1 2 19755 19759
0 19761 5 1 1 19760
0 19762 7 1 2 48168 19761
0 19763 5 1 1 19762
0 19764 7 1 2 59398 72109
0 19765 7 1 2 68763 19764
0 19766 5 1 1 19765
0 19767 7 1 2 19763 19766
0 19768 5 1 1 19767
0 19769 7 1 2 56082 19768
0 19770 5 1 1 19769
0 19771 7 1 2 64887 74434
0 19772 5 1 1 19771
0 19773 7 1 2 19770 19772
0 19774 5 1 1 19773
0 19775 7 1 2 47910 19774
0 19776 5 1 1 19775
0 19777 7 2 2 50713 68470
0 19778 7 1 2 63656 71339
0 19779 7 1 2 62401 19778
0 19780 7 1 2 74646 19779
0 19781 5 1 1 19780
0 19782 7 1 2 63166 71340
0 19783 5 1 1 19782
0 19784 7 1 2 19317 19783
0 19785 5 1 1 19784
0 19786 7 1 2 59313 69002
0 19787 7 1 2 19785 19786
0 19788 5 1 1 19787
0 19789 7 1 2 19781 19788
0 19790 5 1 1 19789
0 19791 7 1 2 58394 19790
0 19792 5 1 1 19791
0 19793 7 1 2 48748 12410
0 19794 7 1 2 72512 19793
0 19795 5 1 1 19794
0 19796 7 1 2 72259 19795
0 19797 5 1 1 19796
0 19798 7 1 2 49205 69003
0 19799 7 1 2 67575 19798
0 19800 7 1 2 19797 19799
0 19801 5 1 1 19800
0 19802 7 1 2 19792 19801
0 19803 5 1 1 19802
0 19804 7 1 2 59989 19803
0 19805 5 1 1 19804
0 19806 7 1 2 62566 66585
0 19807 7 1 2 59279 19806
0 19808 5 1 1 19807
0 19809 7 1 2 68850 19808
0 19810 5 1 1 19809
0 19811 7 1 2 50065 19810
0 19812 5 1 1 19811
0 19813 7 2 2 48749 58490
0 19814 7 1 2 63251 66235
0 19815 7 1 2 69944 19814
0 19816 7 1 2 74648 19815
0 19817 5 1 1 19816
0 19818 7 1 2 71345 19817
0 19819 5 1 1 19818
0 19820 7 1 2 48942 19819
0 19821 5 1 1 19820
0 19822 7 1 2 19812 19821
0 19823 5 1 1 19822
0 19824 7 1 2 67949 19823
0 19825 5 1 1 19824
0 19826 7 1 2 71341 72389
0 19827 7 1 2 68764 19826
0 19828 5 1 1 19827
0 19829 7 1 2 19825 19828
0 19830 7 1 2 19805 19829
0 19831 5 1 1 19830
0 19832 7 1 2 49069 19831
0 19833 5 1 1 19832
0 19834 7 2 2 52281 58426
0 19835 7 1 2 53086 74650
0 19836 5 1 1 19835
0 19837 7 1 2 56908 19836
0 19838 5 1 1 19837
0 19839 7 1 2 54025 72376
0 19840 5 1 1 19839
0 19841 7 1 2 19838 19840
0 19842 5 1 1 19841
0 19843 7 1 2 72282 19842
0 19844 5 1 1 19843
0 19845 7 1 2 65631 74382
0 19846 7 1 2 67381 19845
0 19847 5 1 1 19846
0 19848 7 1 2 611 72816
0 19849 7 1 2 74580 19848
0 19850 5 1 1 19849
0 19851 7 1 2 19847 19850
0 19852 5 1 1 19851
0 19853 7 1 2 74331 19852
0 19854 5 1 1 19853
0 19855 7 1 2 55336 19854
0 19856 7 1 2 19844 19855
0 19857 7 1 2 19833 19856
0 19858 7 1 2 19776 19857
0 19859 5 1 1 19858
0 19860 7 1 2 64400 69380
0 19861 5 1 1 19860
0 19862 7 1 2 59580 68907
0 19863 5 1 1 19862
0 19864 7 1 2 19861 19863
0 19865 5 1 1 19864
0 19866 7 1 2 47911 19865
0 19867 5 1 1 19866
0 19868 7 2 2 49206 49924
0 19869 7 1 2 67950 74652
0 19870 7 1 2 61939 19869
0 19871 5 1 1 19870
0 19872 7 1 2 19867 19871
0 19873 5 1 1 19872
0 19874 7 1 2 48169 19873
0 19875 5 1 1 19874
0 19876 7 1 2 59388 74604
0 19877 5 1 1 19876
0 19878 7 1 2 56083 69358
0 19879 7 1 2 19877 19878
0 19880 5 1 1 19879
0 19881 7 1 2 19875 19880
0 19882 5 1 1 19881
0 19883 7 1 2 71394 19882
0 19884 5 1 1 19883
0 19885 7 2 2 68268 72848
0 19886 5 1 1 74654
0 19887 7 1 2 62402 61728
0 19888 5 1 1 19887
0 19889 7 1 2 59809 70652
0 19890 5 1 1 19889
0 19891 7 1 2 19888 19890
0 19892 5 1 1 19891
0 19893 7 1 2 74655 19892
0 19894 5 1 1 19893
0 19895 7 1 2 19884 19894
0 19896 5 1 1 19895
0 19897 7 1 2 56909 19896
0 19898 5 1 1 19897
0 19899 7 2 2 58427 61129
0 19900 5 1 1 74656
0 19901 7 1 2 69381 19900
0 19902 5 1 1 19901
0 19903 7 1 2 72418 19902
0 19904 5 1 1 19903
0 19905 7 1 2 19904 72230
0 19906 5 1 1 19905
0 19907 7 1 2 51312 19906
0 19908 7 1 2 19898 19907
0 19909 5 1 1 19908
0 19910 7 1 2 19859 19909
0 19911 5 1 1 19910
0 19912 7 1 2 65389 72283
0 19913 5 1 1 19912
0 19914 7 1 2 66974 74435
0 19915 5 1 1 19914
0 19916 7 1 2 19913 19915
0 19917 5 1 1 19916
0 19918 7 1 2 57497 19917
0 19919 5 1 1 19918
0 19920 7 1 2 72483 72199
0 19921 5 1 1 19920
0 19922 7 1 2 65377 67017
0 19923 7 1 2 74628 19922
0 19924 7 1 2 74422 19923
0 19925 5 1 1 19924
0 19926 7 1 2 19921 19925
0 19927 7 1 2 19919 19926
0 19928 5 1 1 19927
0 19929 7 1 2 55337 19928
0 19930 5 1 1 19929
0 19931 7 1 2 64122 69992
0 19932 5 1 1 19931
0 19933 7 5 2 51313 56910
0 19934 5 1 1 74658
0 19935 7 1 2 74659 69017
0 19936 5 1 1 19935
0 19937 7 1 2 19932 19936
0 19938 5 1 1 19937
0 19939 7 1 2 58678 19938
0 19940 5 1 1 19939
0 19941 7 1 2 19940 69221
0 19942 5 1 1 19941
0 19943 7 1 2 51575 19942
0 19944 5 1 1 19943
0 19945 7 1 2 70022 71816
0 19946 5 1 1 19945
0 19947 7 1 2 19944 19946
0 19948 5 1 1 19947
0 19949 7 1 2 50066 19948
0 19950 5 1 1 19949
0 19951 7 1 2 72813 69372
0 19952 5 1 1 19951
0 19953 7 1 2 19950 19952
0 19954 5 1 1 19953
0 19955 7 1 2 49070 19954
0 19956 5 1 1 19955
0 19957 7 1 2 69170 74660
0 19958 5 1 1 19957
0 19959 7 1 2 8936 19958
0 19960 5 1 1 19959
0 19961 7 1 2 74542 19960
0 19962 5 1 1 19961
0 19963 7 1 2 19956 19962
0 19964 5 1 1 19963
0 19965 7 1 2 56084 19964
0 19966 5 1 1 19965
0 19967 7 1 2 61716 74647
0 19968 7 1 2 72176 19967
0 19969 5 1 1 19968
0 19970 7 1 2 69361 19969
0 19971 5 1 1 19970
0 19972 7 1 2 71395 19971
0 19973 5 1 1 19972
0 19974 7 1 2 19973 19886
0 19975 5 1 1 19974
0 19976 7 1 2 74661 19975
0 19977 5 1 1 19976
0 19978 7 1 2 72602 74438
0 19979 5 1 1 19978
0 19980 7 1 2 19977 19979
0 19981 5 1 1 19980
0 19982 7 1 2 54277 19981
0 19983 5 1 1 19982
0 19984 7 1 2 61723 62858
0 19985 5 1 1 19984
0 19986 7 1 2 72266 19985
0 19987 5 1 1 19986
0 19988 7 1 2 19983 19987
0 19989 7 1 2 19966 19988
0 19990 7 1 2 19930 19989
0 19991 5 1 1 19990
0 19992 7 1 2 61837 19991
0 19993 5 1 1 19992
0 19994 7 1 2 56085 74612
0 19995 5 1 1 19994
0 19996 7 1 2 65705 72284
0 19997 5 1 1 19996
0 19998 7 1 2 19995 19997
0 19999 5 1 1 19998
0 20000 7 1 2 60566 19999
0 20001 5 1 1 20000
0 20002 7 3 2 54278 74581
0 20003 5 1 1 74663
0 20004 7 1 2 59990 74664
0 20005 5 1 1 20004
0 20006 7 1 2 68170 20005
0 20007 5 1 1 20006
0 20008 7 1 2 56086 20007
0 20009 5 1 1 20008
0 20010 7 1 2 61865 71925
0 20011 5 1 1 20010
0 20012 7 1 2 70944 20011
0 20013 5 1 1 20012
0 20014 7 1 2 20009 20013
0 20015 5 1 1 20014
0 20016 7 1 2 72267 20015
0 20017 5 1 1 20016
0 20018 7 1 2 20001 20017
0 20019 7 1 2 19993 20018
0 20020 7 1 2 19911 20019
0 20021 7 1 2 19753 20020
0 20022 7 1 2 19681 20021
0 20023 7 1 2 19363 20022
0 20024 5 1 1 20023
0 20025 7 1 2 55001 20024
0 20026 5 1 1 20025
0 20027 7 2 2 49323 74173
0 20028 5 1 1 74666
0 20029 7 1 2 61923 20028
0 20030 5 1 1 20029
0 20031 7 1 2 53906 20030
0 20032 5 1 1 20031
0 20033 7 1 2 60926 59678
0 20034 5 1 1 20033
0 20035 7 1 2 50714 20034
0 20036 5 1 1 20035
0 20037 7 1 2 48170 20036
0 20038 5 1 1 20037
0 20039 7 1 2 59638 20038
0 20040 5 1 1 20039
0 20041 7 1 2 54026 20040
0 20042 5 1 1 20041
0 20043 7 1 2 20032 20042
0 20044 5 1 1 20043
0 20045 7 1 2 49207 20044
0 20046 5 1 1 20045
0 20047 7 1 2 58679 60101
0 20048 5 1 1 20047
0 20049 7 1 2 20046 20048
0 20050 5 1 1 20049
0 20051 7 1 2 48372 20050
0 20052 5 1 1 20051
0 20053 7 1 2 49324 62100
0 20054 5 1 1 20053
0 20055 7 2 2 50191 59715
0 20056 5 1 1 74668
0 20057 7 1 2 20056 68865
0 20058 5 1 1 20057
0 20059 7 1 2 20054 20058
0 20060 5 1 1 20059
0 20061 7 1 2 54279 20060
0 20062 5 1 1 20061
0 20063 7 3 2 49121 59528
0 20064 5 1 1 74670
0 20065 7 1 2 59547 74671
0 20066 5 1 1 20065
0 20067 7 1 2 20062 20066
0 20068 5 1 1 20067
0 20069 7 1 2 54629 20068
0 20070 5 1 1 20069
0 20071 7 1 2 20052 20070
0 20072 5 1 1 20071
0 20073 7 1 2 69839 20072
0 20074 5 1 1 20073
0 20075 7 2 2 49208 62127
0 20076 5 1 1 74673
0 20077 7 1 2 74511 20076
0 20078 5 1 1 20077
0 20079 7 1 2 69963 20078
0 20080 5 1 1 20079
0 20081 7 1 2 57771 69926
0 20082 7 1 2 72034 20081
0 20083 5 1 1 20082
0 20084 7 1 2 20080 20083
0 20085 5 1 1 20084
0 20086 7 1 2 68119 20085
0 20087 5 1 1 20086
0 20088 7 1 2 54280 66852
0 20089 5 1 1 20088
0 20090 7 1 2 57003 20089
0 20091 5 1 1 20090
0 20092 7 1 2 69964 20091
0 20093 5 1 1 20092
0 20094 7 1 2 20087 20093
0 20095 7 1 2 20074 20094
0 20096 5 1 1 20095
0 20097 7 1 2 55338 20096
0 20098 5 1 1 20097
0 20099 7 1 2 62051 69844
0 20100 5 1 1 20099
0 20101 7 1 2 50428 61181
0 20102 5 2 1 20101
0 20103 7 1 2 69965 74675
0 20104 5 1 1 20103
0 20105 7 1 2 20100 20104
0 20106 5 1 1 20105
0 20107 7 1 2 47912 20106
0 20108 5 1 1 20107
0 20109 7 1 2 54281 69966
0 20110 5 2 1 20109
0 20111 7 1 2 69500 69957
0 20112 5 1 1 20111
0 20113 7 1 2 74677 20112
0 20114 5 1 1 20113
0 20115 7 1 2 48171 20114
0 20116 5 1 1 20115
0 20117 7 1 2 49122 69967
0 20118 5 1 1 20117
0 20119 7 1 2 8917 20118
0 20120 5 2 1 20119
0 20121 7 1 2 68034 74679
0 20122 5 1 1 20121
0 20123 7 1 2 20116 20122
0 20124 7 1 2 20108 20123
0 20125 5 1 1 20124
0 20126 7 1 2 65137 20125
0 20127 5 1 1 20126
0 20128 7 2 2 49432 68698
0 20129 7 1 2 58229 74681
0 20130 5 1 1 20129
0 20131 7 1 2 69768 20130
0 20132 5 3 1 20131
0 20133 7 1 2 62101 74683
0 20134 5 1 1 20133
0 20135 7 1 2 62282 68699
0 20136 7 1 2 68055 20135
0 20137 5 1 1 20136
0 20138 7 1 2 20134 20137
0 20139 5 1 1 20138
0 20140 7 1 2 69092 20139
0 20141 5 1 1 20140
0 20142 7 1 2 55652 58230
0 20143 7 1 2 65659 68209
0 20144 7 1 2 20142 20143
0 20145 7 1 2 62089 20144
0 20146 5 1 1 20145
0 20147 7 1 2 20141 20146
0 20148 5 1 1 20147
0 20149 7 1 2 54282 20148
0 20150 5 1 1 20149
0 20151 7 1 2 65932 68030
0 20152 5 1 1 20151
0 20153 7 2 2 64596 69840
0 20154 7 1 2 20152 74686
0 20155 5 1 1 20154
0 20156 7 1 2 58856 69093
0 20157 7 1 2 68035 20156
0 20158 7 1 2 74684 20157
0 20159 5 1 1 20158
0 20160 7 1 2 20155 20159
0 20161 7 1 2 20150 20160
0 20162 5 1 1 20161
0 20163 7 1 2 49325 20162
0 20164 5 1 1 20163
0 20165 7 1 2 20127 20164
0 20166 5 1 1 20165
0 20167 7 1 2 61555 20166
0 20168 5 1 1 20167
0 20169 7 1 2 56911 65248
0 20170 7 1 2 68210 69295
0 20171 7 1 2 20169 20170
0 20172 5 1 1 20171
0 20173 7 1 2 74678 20172
0 20174 5 1 1 20173
0 20175 7 1 2 47913 20174
0 20176 5 1 1 20175
0 20177 7 1 2 54283 74680
0 20178 5 1 1 20177
0 20179 7 1 2 20176 20178
0 20180 5 1 1 20179
0 20181 7 1 2 65554 20180
0 20182 5 1 1 20181
0 20183 7 1 2 60927 68211
0 20184 7 1 2 74632 20183
0 20185 5 1 1 20184
0 20186 7 3 2 69897 68685
0 20187 5 1 1 74688
0 20188 7 1 2 53907 68120
0 20189 7 1 2 74689 20188
0 20190 5 1 1 20189
0 20191 7 1 2 20185 20190
0 20192 5 1 1 20191
0 20193 7 1 2 54284 20192
0 20194 5 1 1 20193
0 20195 7 1 2 62102 68212
0 20196 7 1 2 69853 20195
0 20197 5 1 1 20196
0 20198 7 1 2 20194 20197
0 20199 5 1 1 20198
0 20200 7 1 2 56912 20199
0 20201 5 1 1 20200
0 20202 7 1 2 67097 72059
0 20203 5 1 1 20202
0 20204 7 1 2 69968 72157
0 20205 5 1 1 20204
0 20206 7 1 2 68213 72188
0 20207 5 1 1 20206
0 20208 7 1 2 20187 20207
0 20209 5 1 1 20208
0 20210 7 2 2 56913 58258
0 20211 5 1 1 74691
0 20212 7 1 2 20209 74692
0 20213 5 1 1 20212
0 20214 7 1 2 20205 20213
0 20215 5 1 1 20214
0 20216 7 1 2 58857 20215
0 20217 5 1 1 20216
0 20218 7 1 2 20203 20217
0 20219 7 1 2 20201 20218
0 20220 5 1 1 20219
0 20221 7 1 2 49326 20220
0 20222 5 1 1 20221
0 20223 7 1 2 20182 20222
0 20224 5 1 1 20223
0 20225 7 1 2 61783 20224
0 20226 5 1 1 20225
0 20227 7 2 2 62128 58135
0 20228 5 1 1 74693
0 20229 7 1 2 61423 20228
0 20230 5 1 1 20229
0 20231 7 1 2 69969 20230
0 20232 5 1 1 20231
0 20233 7 1 2 54630 62434
0 20234 5 2 1 20233
0 20235 7 1 2 59710 74674
0 20236 5 1 1 20235
0 20237 7 1 2 74695 20236
0 20238 5 1 1 20237
0 20239 7 1 2 59679 20238
0 20240 5 1 1 20239
0 20241 7 1 2 59639 66854
0 20242 5 1 1 20241
0 20243 7 1 2 54631 20242
0 20244 5 1 1 20243
0 20245 7 1 2 20240 20244
0 20246 5 1 1 20245
0 20247 7 1 2 69841 20246
0 20248 5 1 1 20247
0 20249 7 1 2 20232 20248
0 20250 5 1 1 20249
0 20251 7 1 2 55339 20250
0 20252 5 1 1 20251
0 20253 7 2 2 64964 74690
0 20254 7 1 2 58268 461
0 20255 5 1 1 20254
0 20256 7 1 2 62213 20255
0 20257 7 1 2 74697 20256
0 20258 5 1 1 20257
0 20259 7 1 2 20252 20258
0 20260 5 1 1 20259
0 20261 7 1 2 58858 20260
0 20262 5 1 1 20261
0 20263 7 1 2 67425 74698
0 20264 5 1 1 20263
0 20265 7 3 2 56723 68125
0 20266 7 1 2 50192 60956
0 20267 5 1 1 20266
0 20268 7 1 2 74685 20267
0 20269 7 1 2 74699 20268
0 20270 5 1 1 20269
0 20271 7 1 2 56625 68134
0 20272 5 2 1 20271
0 20273 7 1 2 65138 59138
0 20274 7 1 2 74702 20273
0 20275 5 1 1 20274
0 20276 7 1 2 20270 20275
0 20277 5 1 1 20276
0 20278 7 1 2 69094 20277
0 20279 5 1 1 20278
0 20280 7 1 2 58859 61817
0 20281 7 1 2 74687 20280
0 20282 5 1 1 20281
0 20283 7 1 2 20279 20282
0 20284 5 1 1 20283
0 20285 7 1 2 68164 20284
0 20286 5 1 1 20285
0 20287 7 1 2 20264 20286
0 20288 7 1 2 20262 20287
0 20289 7 1 2 20226 20288
0 20290 7 1 2 20168 20289
0 20291 7 1 2 20098 20290
0 20292 5 1 1 20291
0 20293 7 1 2 49739 20292
0 20294 5 1 1 20293
0 20295 7 1 2 67382 69463
0 20296 7 1 2 69867 20295
0 20297 7 1 2 69893 20296
0 20298 5 1 1 20297
0 20299 7 1 2 20294 20298
0 20300 5 1 1 20299
0 20301 7 1 2 55536 20300
0 20302 5 1 1 20301
0 20303 7 1 2 58479 68471
0 20304 7 1 2 69927 20303
0 20305 7 1 2 74167 20304
0 20306 5 1 1 20305
0 20307 7 1 2 20302 20306
0 20308 5 1 1 20307
0 20309 7 1 2 74360 20308
0 20310 5 1 1 20309
0 20311 7 2 2 54632 61818
0 20312 5 1 1 74704
0 20313 7 1 2 64545 20312
0 20314 5 1 1 20313
0 20315 7 1 2 47914 20314
0 20316 5 1 1 20315
0 20317 7 1 2 2663 57853
0 20318 7 1 2 20316 20317
0 20319 5 1 1 20318
0 20320 7 1 2 54285 20319
0 20321 5 1 1 20320
0 20322 7 1 2 54633 62301
0 20323 5 2 1 20322
0 20324 7 1 2 59338 67297
0 20325 5 1 1 20324
0 20326 7 1 2 74706 20325
0 20327 5 1 1 20326
0 20328 7 1 2 48373 20327
0 20329 5 1 1 20328
0 20330 7 1 2 61024 61751
0 20331 5 2 1 20330
0 20332 7 1 2 20329 74708
0 20333 7 1 2 20321 20332
0 20334 5 2 1 20333
0 20335 7 1 2 74710 69830
0 20336 5 1 1 20335
0 20337 7 1 2 64398 66094
0 20338 5 1 1 20337
0 20339 7 1 2 57498 57825
0 20340 5 1 1 20339
0 20341 7 1 2 48172 63999
0 20342 5 1 1 20341
0 20343 7 1 2 20340 20342
0 20344 5 1 1 20343
0 20345 7 1 2 69831 20344
0 20346 5 1 1 20345
0 20347 7 1 2 5508 20346
0 20348 5 1 1 20347
0 20349 7 1 2 61556 20348
0 20350 5 1 1 20349
0 20351 7 1 2 20338 20350
0 20352 7 1 2 20336 20351
0 20353 5 1 1 20352
0 20354 7 1 2 48943 20353
0 20355 5 1 1 20354
0 20356 7 1 2 66431 65953
0 20357 7 1 2 66790 20356
0 20358 5 1 1 20357
0 20359 7 1 2 20355 20358
0 20360 5 1 1 20359
0 20361 7 1 2 62567 20360
0 20362 5 1 1 20361
0 20363 7 1 2 58269 61396
0 20364 5 2 1 20363
0 20365 7 1 2 62302 74712
0 20366 5 1 1 20365
0 20367 7 4 2 48173 58170
0 20368 5 1 1 74714
0 20369 7 3 2 61752 59339
0 20370 5 1 1 74718
0 20371 7 1 2 20368 20370
0 20372 7 1 2 20366 20371
0 20373 7 1 2 62820 20372
0 20374 5 2 1 20373
0 20375 7 1 2 67516 74721
0 20376 5 1 1 20375
0 20377 7 1 2 1714 71904
0 20378 5 2 1 20377
0 20379 7 2 2 73952 74723
0 20380 7 1 2 74725 72338
0 20381 5 1 1 20380
0 20382 7 1 2 67697 67040
0 20383 7 1 2 74719 20382
0 20384 5 1 1 20383
0 20385 7 1 2 20381 20384
0 20386 5 1 1 20385
0 20387 7 1 2 48374 20386
0 20388 5 1 1 20387
0 20389 7 1 2 62756 66455
0 20390 5 1 1 20389
0 20391 7 2 2 57167 61404
0 20392 7 1 2 62192 71944
0 20393 7 1 2 74727 20392
0 20394 5 1 1 20393
0 20395 7 1 2 20390 20394
0 20396 7 1 2 20388 20395
0 20397 5 1 1 20396
0 20398 7 1 2 62914 20397
0 20399 5 1 1 20398
0 20400 7 1 2 62757 66473
0 20401 5 1 1 20400
0 20402 7 1 2 48375 74726
0 20403 5 1 1 20402
0 20404 7 1 2 64186 20403
0 20405 5 1 1 20404
0 20406 7 1 2 74662 20405
0 20407 5 1 1 20406
0 20408 7 1 2 20401 20407
0 20409 5 1 1 20408
0 20410 7 1 2 72133 20409
0 20411 5 1 1 20410
0 20412 7 1 2 20399 20411
0 20413 5 1 1 20412
0 20414 7 1 2 54634 20413
0 20415 5 1 1 20414
0 20416 7 1 2 20376 20415
0 20417 7 1 2 20362 20416
0 20418 5 1 1 20417
0 20419 7 1 2 49071 20418
0 20420 5 1 1 20419
0 20421 7 1 2 63089 56724
0 20422 5 1 1 20421
0 20423 7 1 2 64123 60998
0 20424 5 1 1 20423
0 20425 7 1 2 20422 20424
0 20426 5 1 1 20425
0 20427 7 1 2 56087 20426
0 20428 5 1 1 20427
0 20429 7 1 2 57281 74625
0 20430 5 1 1 20429
0 20431 7 1 2 20428 20430
0 20432 5 1 1 20431
0 20433 7 1 2 20432 69923
0 20434 5 1 1 20433
0 20435 7 2 2 70386 72339
0 20436 5 1 1 74729
0 20437 7 1 2 57004 71992
0 20438 5 2 1 20437
0 20439 7 2 2 51576 63090
0 20440 7 1 2 74731 74733
0 20441 5 1 1 20440
0 20442 7 1 2 20436 20441
0 20443 5 1 1 20442
0 20444 7 1 2 49072 20443
0 20445 5 1 1 20444
0 20446 7 2 2 62568 56725
0 20447 7 2 2 69176 74735
0 20448 5 1 1 74737
0 20449 7 1 2 65632 71759
0 20450 7 1 2 59265 20449
0 20451 5 1 1 20450
0 20452 7 1 2 20448 20451
0 20453 5 1 1 20452
0 20454 7 1 2 65546 20453
0 20455 5 1 1 20454
0 20456 7 1 2 49073 71760
0 20457 5 1 1 20456
0 20458 7 1 2 20455 20457
0 20459 5 1 1 20458
0 20460 7 1 2 55340 20459
0 20461 5 1 1 20460
0 20462 7 1 2 67033 74730
0 20463 5 1 1 20462
0 20464 7 1 2 20461 20463
0 20465 7 1 2 20445 20464
0 20466 5 1 1 20465
0 20467 7 1 2 54635 20466
0 20468 5 1 1 20467
0 20469 7 1 2 20434 20468
0 20470 5 1 1 20469
0 20471 7 1 2 47915 20470
0 20472 5 1 1 20471
0 20473 7 1 2 73980 74736
0 20474 5 1 1 20473
0 20475 7 2 2 63091 69177
0 20476 5 1 1 74739
0 20477 7 1 2 69999 72421
0 20478 5 1 1 20477
0 20479 7 1 2 20476 20478
0 20480 5 1 1 20479
0 20481 7 1 2 56088 20480
0 20482 5 1 1 20481
0 20483 7 1 2 66386 74386
0 20484 5 1 1 20483
0 20485 7 1 2 57168 74734
0 20486 5 1 1 20485
0 20487 7 1 2 74153 20486
0 20488 5 1 1 20487
0 20489 7 1 2 49074 20488
0 20490 5 1 1 20489
0 20491 7 1 2 20484 20490
0 20492 7 1 2 20482 20491
0 20493 5 1 1 20492
0 20494 7 1 2 54286 20493
0 20495 5 1 1 20494
0 20496 7 1 2 56089 64597
0 20497 7 1 2 74738 20496
0 20498 5 1 1 20497
0 20499 7 1 2 20495 20498
0 20500 5 1 1 20499
0 20501 7 1 2 56914 20500
0 20502 5 1 1 20501
0 20503 7 1 2 20474 20502
0 20504 7 1 2 20472 20503
0 20505 5 1 1 20504
0 20506 7 1 2 54027 20505
0 20507 5 1 1 20506
0 20508 7 2 2 63965 64124
0 20509 5 1 1 74741
0 20510 7 1 2 5731 20509
0 20511 5 1 1 20510
0 20512 7 1 2 54287 20511
0 20513 5 1 1 20512
0 20514 7 1 2 54636 63092
0 20515 5 1 1 20514
0 20516 7 1 2 20513 20515
0 20517 5 1 1 20516
0 20518 7 1 2 51577 20517
0 20519 5 1 1 20518
0 20520 7 1 2 61109 71829
0 20521 5 1 1 20520
0 20522 7 1 2 20519 20521
0 20523 5 1 1 20522
0 20524 7 1 2 49075 20523
0 20525 5 1 1 20524
0 20526 7 1 2 66387 68617
0 20527 7 1 2 74250 20526
0 20528 5 1 1 20527
0 20529 7 1 2 20525 20528
0 20530 5 1 1 20529
0 20531 7 1 2 56726 20530
0 20532 5 1 1 20531
0 20533 7 2 2 64125 69178
0 20534 7 1 2 61135 74743
0 20535 5 1 1 20534
0 20536 7 1 2 57499 71960
0 20537 7 1 2 70000 20536
0 20538 5 1 1 20537
0 20539 7 1 2 20535 20538
0 20540 5 1 1 20539
0 20541 7 1 2 57169 20540
0 20542 5 1 1 20541
0 20543 7 1 2 59705 74744
0 20544 5 1 1 20543
0 20545 7 1 2 20542 20544
0 20546 5 1 1 20545
0 20547 7 1 2 54637 20546
0 20548 5 1 1 20547
0 20549 7 1 2 47916 74740
0 20550 7 1 2 62458 20549
0 20551 5 1 1 20550
0 20552 7 1 2 20548 20551
0 20553 7 1 2 20532 20552
0 20554 5 1 1 20553
0 20555 7 1 2 56915 20554
0 20556 5 1 1 20555
0 20557 7 1 2 73940 69227
0 20558 5 1 1 20557
0 20559 7 1 2 74205 74588
0 20560 5 1 1 20559
0 20561 7 1 2 20558 20560
0 20562 7 1 2 20556 20561
0 20563 7 1 2 20507 20562
0 20564 5 1 1 20563
0 20565 7 1 2 49925 20564
0 20566 5 1 1 20565
0 20567 7 1 2 20420 20566
0 20568 5 1 1 20567
0 20569 7 1 2 55750 20568
0 20570 5 1 1 20569
0 20571 7 1 2 65290 65650
0 20572 7 1 2 74649 20571
0 20573 5 1 1 20572
0 20574 7 1 2 52868 20573
0 20575 5 1 1 20574
0 20576 7 1 2 71761 20575
0 20577 5 1 1 20576
0 20578 7 1 2 50429 74007
0 20579 5 1 1 20578
0 20580 7 1 2 47917 20579
0 20581 5 1 1 20580
0 20582 7 1 2 61701 74199
0 20583 5 1 1 20582
0 20584 7 2 2 61866 20583
0 20585 5 1 1 74745
0 20586 7 1 2 61525 65001
0 20587 5 2 1 20586
0 20588 7 1 2 49327 74747
0 20589 5 1 1 20588
0 20590 7 1 2 74746 20589
0 20591 7 1 2 20581 20590
0 20592 5 1 1 20591
0 20593 7 1 2 71888 20592
0 20594 5 1 1 20593
0 20595 7 1 2 20577 20594
0 20596 5 1 1 20595
0 20597 7 1 2 74194 20596
0 20598 5 1 1 20597
0 20599 7 2 2 49209 67478
0 20600 7 1 2 68621 74749
0 20601 5 1 1 20600
0 20602 7 1 2 5465 20601
0 20603 5 1 1 20602
0 20604 7 6 2 58395 63252
0 20605 7 1 2 20603 74751
0 20606 5 1 1 20605
0 20607 7 4 2 47918 61557
0 20608 5 2 1 74757
0 20609 7 2 2 64208 74761
0 20610 5 1 1 74763
0 20611 7 1 2 53087 74764
0 20612 5 1 1 20611
0 20613 7 1 2 48376 20612
0 20614 5 1 1 20613
0 20615 7 1 2 59680 61965
0 20616 5 1 1 20615
0 20617 7 2 2 53088 71404
0 20618 5 4 1 74765
0 20619 7 1 2 71429 74767
0 20620 5 1 1 20619
0 20621 7 1 2 57780 60064
0 20622 5 1 1 20621
0 20623 7 1 2 47919 20622
0 20624 5 1 1 20623
0 20625 7 1 2 20620 20624
0 20626 7 1 2 20616 20625
0 20627 7 1 2 20614 20626
0 20628 5 1 1 20627
0 20629 7 1 2 48174 20628
0 20630 5 1 1 20629
0 20631 7 1 2 48377 61635
0 20632 5 1 1 20631
0 20633 7 1 2 61875 20632
0 20634 7 1 2 65783 20633
0 20635 5 1 1 20634
0 20636 7 1 2 54288 20635
0 20637 5 1 1 20636
0 20638 7 1 2 47920 62803
0 20639 5 1 1 20638
0 20640 7 1 2 57601 74196
0 20641 5 1 1 20640
0 20642 7 1 2 62665 20641
0 20643 5 1 1 20642
0 20644 7 1 2 20639 20643
0 20645 7 1 2 20637 20644
0 20646 7 1 2 20630 20645
0 20647 5 1 1 20646
0 20648 7 1 2 66397 20647
0 20649 5 1 1 20648
0 20650 7 1 2 20606 20649
0 20651 5 1 1 20650
0 20652 7 1 2 63167 20651
0 20653 5 1 1 20652
0 20654 7 1 2 59991 61972
0 20655 5 2 1 20654
0 20656 7 1 2 57227 59655
0 20657 7 1 2 74771 20656
0 20658 5 1 1 20657
0 20659 7 1 2 71762 20658
0 20660 5 1 1 20659
0 20661 7 2 2 56916 71877
0 20662 7 1 2 58298 74578
0 20663 5 1 1 20662
0 20664 7 1 2 54289 20663
0 20665 5 1 1 20664
0 20666 7 1 2 59332 20665
0 20667 5 1 1 20666
0 20668 7 1 2 59992 20667
0 20669 5 1 1 20668
0 20670 7 1 2 65186 56727
0 20671 5 1 1 20670
0 20672 7 1 2 68073 20671
0 20673 5 1 1 20672
0 20674 7 1 2 49328 20673
0 20675 5 1 1 20674
0 20676 7 2 2 60972 61858
0 20677 5 3 1 74775
0 20678 7 1 2 20675 74777
0 20679 7 1 2 20669 20678
0 20680 5 1 1 20679
0 20681 7 1 2 74773 20680
0 20682 5 1 1 20681
0 20683 7 1 2 20660 20682
0 20684 5 1 1 20683
0 20685 7 1 2 49926 20684
0 20686 5 1 1 20685
0 20687 7 2 2 57271 74772
0 20688 5 1 1 74780
0 20689 7 1 2 55884 74781
0 20690 5 1 1 20689
0 20691 7 1 2 66501 20690
0 20692 5 1 1 20691
0 20693 7 1 2 20686 20692
0 20694 7 1 2 20653 20693
0 20695 5 1 1 20694
0 20696 7 1 2 49076 20695
0 20697 5 1 1 20696
0 20698 7 1 2 20598 20697
0 20699 5 1 1 20698
0 20700 7 1 2 55341 20699
0 20701 5 1 1 20700
0 20702 7 1 2 64993 63029
0 20703 5 2 1 20702
0 20704 7 1 2 67303 74782
0 20705 5 2 1 20704
0 20706 7 1 2 65887 74784
0 20707 5 1 1 20706
0 20708 7 1 2 61964 74762
0 20709 7 1 2 67458 20708
0 20710 5 1 1 20709
0 20711 7 1 2 61271 20710
0 20712 5 1 1 20711
0 20713 7 1 2 20707 20712
0 20714 5 1 1 20713
0 20715 7 1 2 74384 72814
0 20716 7 1 2 20714 20715
0 20717 5 1 1 20716
0 20718 7 1 2 20701 20717
0 20719 5 1 1 20718
0 20720 7 1 2 54638 20719
0 20721 5 1 1 20720
0 20722 7 2 2 54290 62303
0 20723 7 1 2 47921 74786
0 20724 5 1 1 20723
0 20725 7 1 2 62791 20724
0 20726 5 1 1 20725
0 20727 7 1 2 62052 20726
0 20728 5 1 1 20727
0 20729 7 1 2 49329 60129
0 20730 5 2 1 20729
0 20731 7 1 2 62268 74788
0 20732 5 1 1 20731
0 20733 7 1 2 54291 20732
0 20734 5 1 1 20733
0 20735 7 1 2 4417 20734
0 20736 5 1 1 20735
0 20737 7 1 2 61558 20736
0 20738 5 1 1 20737
0 20739 7 3 2 61753 59616
0 20740 5 2 1 74790
0 20741 7 1 2 20738 74793
0 20742 7 1 2 20728 20741
0 20743 5 1 1 20742
0 20744 7 2 2 72340 20743
0 20745 5 1 1 74795
0 20746 7 1 2 62345 64074
0 20747 5 1 1 20746
0 20748 7 1 2 57005 20747
0 20749 5 3 1 20748
0 20750 7 1 2 66985 74797
0 20751 5 1 1 20750
0 20752 7 1 2 20745 20751
0 20753 5 1 1 20752
0 20754 7 1 2 69574 20753
0 20755 5 1 1 20754
0 20756 7 1 2 62915 74796
0 20757 5 1 1 20756
0 20758 7 1 2 72351 74798
0 20759 5 1 1 20758
0 20760 7 1 2 20757 20759
0 20761 7 1 2 20755 20760
0 20762 5 1 1 20761
0 20763 7 1 2 48378 20762
0 20764 5 1 1 20763
0 20765 7 1 2 69575 69228
0 20766 5 1 1 20765
0 20767 7 1 2 57170 74574
0 20768 5 1 1 20767
0 20769 7 1 2 61973 66986
0 20770 5 1 1 20769
0 20771 7 1 2 20768 20770
0 20772 5 1 1 20771
0 20773 7 1 2 69576 20772
0 20774 5 1 1 20773
0 20775 7 1 2 61974 72352
0 20776 5 1 1 20775
0 20777 7 1 2 62916 59329
0 20778 7 1 2 71937 20777
0 20779 5 1 1 20778
0 20780 7 1 2 20776 20779
0 20781 7 1 2 20774 20780
0 20782 5 1 1 20781
0 20783 7 1 2 47922 20782
0 20784 5 1 1 20783
0 20785 7 1 2 68047 74766
0 20786 5 1 1 20785
0 20787 7 1 2 67449 69577
0 20788 7 1 2 68358 20787
0 20789 5 1 1 20788
0 20790 7 1 2 62917 60928
0 20791 7 1 2 59617 20790
0 20792 7 1 2 73982 20791
0 20793 5 1 1 20792
0 20794 7 1 2 20789 20793
0 20795 5 1 1 20794
0 20796 7 1 2 61838 20795
0 20797 5 1 1 20796
0 20798 7 1 2 74488 20797
0 20799 5 1 1 20798
0 20800 7 1 2 20786 20799
0 20801 5 1 1 20800
0 20802 7 1 2 20784 20801
0 20803 5 1 1 20802
0 20804 7 1 2 56917 20803
0 20805 5 1 1 20804
0 20806 7 1 2 20766 20805
0 20807 7 1 2 20764 20806
0 20808 5 1 1 20807
0 20809 7 1 2 54639 20808
0 20810 5 1 1 20809
0 20811 7 1 2 61988 65888
0 20812 5 1 1 20811
0 20813 7 3 2 58396 56090
0 20814 5 1 1 74800
0 20815 7 1 2 65033 61072
0 20816 7 1 2 20814 20815
0 20817 5 2 1 20816
0 20818 7 1 2 61839 74803
0 20819 5 2 1 20818
0 20820 7 1 2 61101 67298
0 20821 5 1 1 20820
0 20822 7 2 2 59640 61867
0 20823 5 1 1 74807
0 20824 7 1 2 48379 20823
0 20825 5 1 1 20824
0 20826 7 1 2 20821 20825
0 20827 7 1 2 74805 20826
0 20828 7 2 2 20812 20827
0 20829 5 1 1 74809
0 20830 7 1 2 56918 20829
0 20831 5 1 1 20830
0 20832 7 1 2 51314 20831
0 20833 5 1 1 20832
0 20834 7 1 2 74491 20833
0 20835 5 1 1 20834
0 20836 7 1 2 66343 71949
0 20837 5 1 1 20836
0 20838 7 1 2 11551 20837
0 20839 5 1 1 20838
0 20840 7 1 2 62053 20839
0 20841 5 1 1 20840
0 20842 7 1 2 55537 74191
0 20843 5 1 1 20842
0 20844 7 1 2 20841 20843
0 20845 5 1 1 20844
0 20846 7 1 2 61559 20845
0 20847 5 1 1 20846
0 20848 7 1 2 50430 65404
0 20849 5 1 1 20848
0 20850 7 1 2 47923 20849
0 20851 5 2 1 20850
0 20852 7 1 2 58327 61620
0 20853 5 1 1 20852
0 20854 7 1 2 58180 20853
0 20855 7 1 2 74811 20854
0 20856 5 1 1 20855
0 20857 7 1 2 66095 20856
0 20858 5 1 1 20857
0 20859 7 1 2 62015 66853
0 20860 7 1 2 72546 20859
0 20861 5 1 1 20860
0 20862 7 1 2 20858 20861
0 20863 7 1 2 60130 66096
0 20864 5 1 1 20863
0 20865 7 1 2 65440 72149
0 20866 7 1 2 74715 20865
0 20867 5 1 1 20866
0 20868 7 1 2 20864 20867
0 20869 5 1 1 20868
0 20870 7 1 2 62304 20869
0 20871 5 1 1 20870
0 20872 7 1 2 60416 60029
0 20873 5 2 1 20872
0 20874 7 2 2 64306 62259
0 20875 7 1 2 62009 72150
0 20876 7 1 2 74815 20875
0 20877 5 1 1 20876
0 20878 7 1 2 66116 20877
0 20879 5 1 1 20878
0 20880 7 1 2 74813 20879
0 20881 5 1 1 20880
0 20882 7 1 2 20871 20881
0 20883 7 1 2 20862 20882
0 20884 7 1 2 20847 20883
0 20885 5 1 1 20884
0 20886 7 1 2 69578 20885
0 20887 5 1 1 20886
0 20888 7 1 2 72362 20887
0 20889 5 1 1 20888
0 20890 7 1 2 62569 20889
0 20891 5 1 1 20890
0 20892 7 1 2 20835 20891
0 20893 7 1 2 20810 20892
0 20894 5 1 1 20893
0 20895 7 1 2 49077 20894
0 20896 5 1 1 20895
0 20897 7 1 2 20721 20896
0 20898 7 1 2 20570 20897
0 20899 5 1 1 20898
0 20900 7 1 2 51770 20899
0 20901 5 1 1 20900
0 20902 7 1 2 55751 74722
0 20903 5 1 1 20902
0 20904 7 1 2 57006 20903
0 20905 7 1 2 74810 20904
0 20906 5 2 1 20905
0 20907 7 1 2 74456 74817
0 20908 5 1 1 20907
0 20909 7 4 2 53485 65985
0 20910 7 1 2 49123 74160
0 20911 5 1 1 20910
0 20912 7 1 2 68150 20911
0 20913 5 1 1 20912
0 20914 7 1 2 47924 20913
0 20915 5 1 1 20914
0 20916 7 1 2 48380 74593
0 20917 5 1 1 20916
0 20918 7 1 2 20915 20917
0 20919 5 1 1 20918
0 20920 7 1 2 58205 20919
0 20921 5 1 1 20920
0 20922 7 1 2 56919 74212
0 20923 5 1 1 20922
0 20924 7 1 2 20921 20923
0 20925 5 1 1 20924
0 20926 7 1 2 61560 20925
0 20927 5 1 1 20926
0 20928 7 1 2 55752 74713
0 20929 5 1 1 20928
0 20930 7 1 2 58347 62054
0 20931 5 1 1 20930
0 20932 7 1 2 20929 20931
0 20933 5 1 1 20932
0 20934 7 1 2 49330 20933
0 20935 5 1 1 20934
0 20936 7 2 2 58397 58187
0 20937 5 1 1 74823
0 20938 7 1 2 20935 20937
0 20939 5 1 1 20938
0 20940 7 1 2 54640 61754
0 20941 7 1 2 20939 20940
0 20942 5 1 1 20941
0 20943 7 1 2 49210 60715
0 20944 5 2 1 20943
0 20945 7 1 2 51910 74825
0 20946 5 1 1 20945
0 20947 7 1 2 65559 20946
0 20948 5 1 1 20947
0 20949 7 1 2 60849 20948
0 20950 5 2 1 20949
0 20951 7 1 2 64975 66195
0 20952 5 1 1 20951
0 20953 7 1 2 74827 20952
0 20954 5 1 1 20953
0 20955 7 1 2 60090 58323
0 20956 5 1 1 20955
0 20957 7 1 2 61627 70749
0 20958 5 1 1 20957
0 20959 7 1 2 20956 20958
0 20960 5 1 1 20959
0 20961 7 1 2 67428 20960
0 20962 5 1 1 20961
0 20963 7 1 2 56920 20962
0 20964 5 1 1 20963
0 20965 7 1 2 57007 18464
0 20966 5 1 1 20965
0 20967 7 10 2 50090 58835
0 20968 5 4 1 74829
0 20969 7 1 2 62305 74839
0 20970 7 1 2 20966 20969
0 20971 5 1 1 20970
0 20972 7 1 2 52615 20971
0 20973 7 1 2 20964 20972
0 20974 7 1 2 20954 20973
0 20975 7 1 2 20942 20974
0 20976 7 1 2 20927 20975
0 20977 5 1 1 20976
0 20978 7 1 2 74819 20977
0 20979 5 1 1 20978
0 20980 7 1 2 58718 72406
0 20981 5 1 1 20980
0 20982 7 2 2 53908 62323
0 20983 5 1 1 74843
0 20984 7 1 2 49211 74844
0 20985 5 1 1 20984
0 20986 7 1 2 50715 20985
0 20987 5 3 1 20986
0 20988 7 1 2 54292 74845
0 20989 5 1 1 20988
0 20990 7 2 2 63030 65949
0 20991 5 2 1 74848
0 20992 7 1 2 20989 74850
0 20993 5 1 1 20992
0 20994 7 1 2 58860 20993
0 20995 5 2 1 20994
0 20996 7 1 2 65249 56728
0 20997 5 1 1 20996
0 20998 7 1 2 60929 60999
0 20999 5 1 1 20998
0 21000 7 1 2 20997 20999
0 21001 5 1 1 21000
0 21002 7 1 2 54028 21001
0 21003 5 1 1 21002
0 21004 7 1 2 3416 21003
0 21005 7 1 2 74852 21004
0 21006 5 1 1 21005
0 21007 7 1 2 56091 21006
0 21008 5 1 1 21007
0 21009 7 1 2 61136 63982
0 21010 5 1 1 21009
0 21011 7 1 2 60930 64031
0 21012 5 1 1 21011
0 21013 7 1 2 21010 21012
0 21014 5 1 1 21013
0 21015 7 1 2 48175 21014
0 21016 5 1 1 21015
0 21017 7 1 2 58680 74525
0 21018 5 1 1 21017
0 21019 7 1 2 21016 21018
0 21020 5 1 1 21019
0 21021 7 1 2 60693 21020
0 21022 5 1 1 21021
0 21023 7 1 2 64000 74200
0 21024 5 1 1 21023
0 21025 7 2 2 54293 62155
0 21026 5 2 1 74854
0 21027 7 1 2 50716 74856
0 21028 5 1 1 21027
0 21029 7 1 2 57500 21028
0 21030 5 1 1 21029
0 21031 7 1 2 21024 21030
0 21032 5 1 1 21031
0 21033 7 1 2 61702 21032
0 21034 5 1 1 21033
0 21035 7 3 2 56729 58861
0 21036 7 2 2 61851 74858
0 21037 5 1 1 74861
0 21038 7 1 2 54294 74862
0 21039 5 1 1 21038
0 21040 7 1 2 74778 21039
0 21041 5 1 1 21040
0 21042 7 1 2 54641 21041
0 21043 5 1 1 21042
0 21044 7 1 2 58862 74846
0 21045 5 2 1 21044
0 21046 7 1 2 54642 715
0 21047 5 1 1 21046
0 21048 7 1 2 57008 21047
0 21049 7 1 2 63035 21048
0 21050 7 1 2 74863 21049
0 21051 5 1 1 21050
0 21052 7 1 2 70945 21051
0 21053 5 1 1 21052
0 21054 7 1 2 21043 21053
0 21055 7 1 2 21034 21054
0 21056 7 1 2 21022 21055
0 21057 7 1 2 21008 21056
0 21058 5 1 1 21057
0 21059 7 1 2 71878 21058
0 21060 5 1 1 21059
0 21061 7 1 2 20981 21060
0 21062 5 1 1 21061
0 21063 7 1 2 51315 21062
0 21064 5 1 1 21063
0 21065 7 1 2 20979 21064
0 21066 5 1 1 21065
0 21067 7 1 2 68553 21066
0 21068 5 1 1 21067
0 21069 7 1 2 20908 21068
0 21070 5 1 1 21069
0 21071 7 1 2 49078 21070
0 21072 5 1 1 21071
0 21073 7 1 2 67679 67951
0 21074 7 1 2 74818 21073
0 21075 5 1 1 21074
0 21076 7 2 2 58149 63694
0 21077 5 1 1 74865
0 21078 7 1 2 66569 72493
0 21079 7 1 2 74866 21078
0 21080 5 1 1 21079
0 21081 7 1 2 21075 21080
0 21082 5 1 1 21081
0 21083 7 1 2 73593 72242
0 21084 7 1 2 21082 21083
0 21085 5 1 1 21084
0 21086 7 1 2 21072 21085
0 21087 5 1 1 21086
0 21088 7 1 2 51015 21087
0 21089 5 1 1 21088
0 21090 7 1 2 52801 66965
0 21091 7 1 2 66474 72032
0 21092 7 1 2 21090 21091
0 21093 5 1 1 21092
0 21094 7 1 2 21089 21093
0 21095 7 1 2 20901 21094
0 21096 5 1 1 21095
0 21097 7 1 2 50067 21096
0 21098 5 1 1 21097
0 21099 7 1 2 20310 21098
0 21100 7 1 2 20026 21099
0 21101 5 1 1 21100
0 21102 7 1 2 56550 21101
0 21103 5 1 1 21102
0 21104 7 2 2 52954 62606
0 21105 5 2 1 74867
0 21106 7 1 2 70750 74868
0 21107 5 1 1 21106
0 21108 7 4 2 54295 55885
0 21109 7 1 2 50193 74871
0 21110 5 1 1 21109
0 21111 7 1 2 21107 21110
0 21112 5 1 1 21111
0 21113 7 1 2 51911 21112
0 21114 5 2 1 21113
0 21115 7 1 2 52122 63172
0 21116 5 1 1 21115
0 21117 7 2 2 62615 21116
0 21118 5 2 1 74877
0 21119 7 1 2 54296 60867
0 21120 5 1 1 21119
0 21121 7 1 2 74878 21120
0 21122 5 1 1 21121
0 21123 7 1 2 55886 21122
0 21124 5 1 1 21123
0 21125 7 1 2 74875 21124
0 21126 5 1 1 21125
0 21127 7 1 2 50717 21126
0 21128 5 1 1 21127
0 21129 7 2 2 54643 70274
0 21130 5 1 1 74881
0 21131 7 1 2 59760 74882
0 21132 5 1 1 21131
0 21133 7 1 2 21128 21132
0 21134 5 1 1 21133
0 21135 7 1 2 63574 21134
0 21136 5 1 1 21135
0 21137 7 1 2 51016 65678
0 21138 5 2 1 21137
0 21139 7 6 2 52955 63606
0 21140 5 1 1 74885
0 21141 7 2 2 55689 74886
0 21142 5 1 1 74891
0 21143 7 1 2 50431 74892
0 21144 5 1 1 21143
0 21145 7 1 2 74883 21144
0 21146 5 1 1 21145
0 21147 7 1 2 48944 21146
0 21148 5 1 1 21147
0 21149 7 1 2 21136 21148
0 21150 5 1 1 21149
0 21151 7 1 2 58756 21150
0 21152 5 1 1 21151
0 21153 7 2 2 53089 60850
0 21154 5 1 1 74893
0 21155 7 1 2 52282 74894
0 21156 5 3 1 21155
0 21157 7 2 2 60818 74895
0 21158 5 1 1 74898
0 21159 7 1 2 52956 21158
0 21160 5 2 1 21159
0 21161 7 3 2 70279 74900
0 21162 5 1 1 74902
0 21163 7 1 2 52283 70520
0 21164 5 1 1 21163
0 21165 7 1 2 74903 21164
0 21166 5 1 1 21165
0 21167 7 1 2 50718 21166
0 21168 5 1 1 21167
0 21169 7 2 2 51017 60417
0 21170 5 3 1 74905
0 21171 7 1 2 48176 74907
0 21172 5 1 1 21171
0 21173 7 1 2 60507 21172
0 21174 5 1 1 21173
0 21175 7 1 2 21168 21174
0 21176 5 2 1 21175
0 21177 7 1 2 63420 74910
0 21178 5 1 1 21177
0 21179 7 2 2 65019 70793
0 21180 5 1 1 74912
0 21181 7 1 2 51912 21180
0 21182 5 1 1 21181
0 21183 7 2 2 70284 21182
0 21184 5 6 1 74914
0 21185 7 1 2 56092 74915
0 21186 5 1 1 21185
0 21187 7 1 2 59139 21186
0 21188 5 1 1 21187
0 21189 7 1 2 65002 70701
0 21190 5 1 1 21189
0 21191 7 1 2 21188 21190
0 21192 5 1 1 21191
0 21193 7 1 2 48945 21192
0 21194 5 1 1 21193
0 21195 7 2 2 60177 70745
0 21196 7 1 2 54644 74922
0 21197 5 1 1 21196
0 21198 7 1 2 60567 61449
0 21199 5 1 1 21198
0 21200 7 1 2 63429 21199
0 21201 5 1 1 21200
0 21202 7 1 2 21197 21201
0 21203 5 1 1 21202
0 21204 7 1 2 60358 63482
0 21205 5 1 1 21204
0 21206 7 1 2 59899 73893
0 21207 7 1 2 72797 21206
0 21208 5 1 1 21207
0 21209 7 1 2 21205 21208
0 21210 5 1 1 21209
0 21211 7 1 2 60335 21210
0 21212 5 1 1 21211
0 21213 7 1 2 21203 21212
0 21214 7 1 2 21194 21213
0 21215 5 1 1 21214
0 21216 7 1 2 58005 21215
0 21217 5 1 1 21216
0 21218 7 1 2 21178 21217
0 21219 7 1 2 21152 21218
0 21220 5 1 1 21219
0 21221 7 1 2 55342 21220
0 21222 5 1 1 21221
0 21223 7 3 2 65465 60851
0 21224 5 1 1 74924
0 21225 7 1 2 60325 21224
0 21226 5 1 1 21225
0 21227 7 1 2 50719 21226
0 21228 5 1 1 21227
0 21229 7 1 2 55887 685
0 21230 5 1 1 21229
0 21231 7 2 2 65445 55690
0 21232 5 1 1 74927
0 21233 7 1 2 56093 21232
0 21234 5 1 1 21233
0 21235 7 1 2 60175 21234
0 21236 5 1 1 21235
0 21237 7 1 2 21230 21236
0 21238 7 2 2 21228 21237
0 21239 7 1 2 64454 74929
0 21240 5 1 1 21239
0 21241 7 1 2 63487 67753
0 21242 7 1 2 21240 21241
0 21243 5 1 1 21242
0 21244 7 1 2 21222 21243
0 21245 5 1 1 21244
0 21246 7 1 2 73852 21245
0 21247 5 1 1 21246
0 21248 7 1 2 49927 73901
0 21249 5 2 1 21248
0 21250 7 1 2 70566 74931
0 21251 5 3 1 21250
0 21252 7 2 2 50720 74916
0 21253 5 1 1 74936
0 21254 7 1 2 74933 74937
0 21255 5 1 1 21254
0 21256 7 3 2 58006 70571
0 21257 7 1 2 50432 74938
0 21258 5 1 1 21257
0 21259 7 1 2 21255 21258
0 21260 5 1 1 21259
0 21261 7 1 2 55888 21260
0 21262 5 1 1 21261
0 21263 7 1 2 50433 13402
0 21264 5 1 1 21263
0 21265 7 1 2 54645 21264
0 21266 5 3 1 21265
0 21267 7 1 2 74939 74941
0 21268 5 1 1 21267
0 21269 7 1 2 21262 21268
0 21270 5 1 1 21269
0 21271 7 1 2 66604 21270
0 21272 5 1 1 21271
0 21273 7 3 2 60471 72754
0 21274 5 1 1 74944
0 21275 7 1 2 60678 74945
0 21276 5 1 1 21275
0 21277 7 1 2 60568 21276
0 21278 5 1 1 21277
0 21279 7 1 2 52123 21278
0 21280 5 2 1 21279
0 21281 7 1 2 719 74947
0 21282 5 1 1 21281
0 21283 7 1 2 51913 21282
0 21284 5 1 1 21283
0 21285 7 1 2 59767 71166
0 21286 5 1 1 21285
0 21287 7 1 2 52124 21286
0 21288 5 1 1 21287
0 21289 7 1 2 63627 21288
0 21290 5 1 1 21289
0 21291 7 1 2 50434 21290
0 21292 5 2 1 21291
0 21293 7 1 2 21284 74949
0 21294 5 1 1 21293
0 21295 7 2 2 55343 21294
0 21296 7 1 2 53486 74951
0 21297 5 1 1 21296
0 21298 7 2 2 61526 60640
0 21299 5 1 1 74953
0 21300 7 1 2 56094 21299
0 21301 5 2 1 21300
0 21302 7 2 2 58681 73368
0 21303 5 1 1 74957
0 21304 7 1 2 63801 21303
0 21305 5 2 1 21304
0 21306 7 1 2 74955 74959
0 21307 5 1 1 21306
0 21308 7 3 2 50194 58682
0 21309 5 4 1 74961
0 21310 7 1 2 74964 70537
0 21311 5 1 1 21310
0 21312 7 1 2 55889 21311
0 21313 5 1 1 21312
0 21314 7 1 2 49740 74942
0 21315 5 1 1 21314
0 21316 7 1 2 21313 21315
0 21317 5 1 1 21316
0 21318 7 1 2 51316 21317
0 21319 5 1 1 21318
0 21320 7 1 2 21307 21319
0 21321 7 1 2 21297 21320
0 21322 5 1 1 21321
0 21323 7 1 2 51018 21322
0 21324 5 1 1 21323
0 21325 7 1 2 60504 73128
0 21326 5 1 1 21325
0 21327 7 1 2 50195 68663
0 21328 5 1 1 21327
0 21329 7 1 2 21326 21328
0 21330 5 1 1 21329
0 21331 7 1 2 51914 21330
0 21332 5 1 1 21331
0 21333 7 1 2 68664 70193
0 21334 5 1 1 21333
0 21335 7 1 2 21332 21334
0 21336 5 1 1 21335
0 21337 7 1 2 52125 21336
0 21338 5 1 1 21337
0 21339 7 1 2 68665 9216
0 21340 5 1 1 21339
0 21341 7 1 2 63804 73030
0 21342 7 1 2 73563 21341
0 21343 5 1 1 21342
0 21344 7 1 2 73927 21343
0 21345 7 1 2 21340 21344
0 21346 7 1 2 21338 21345
0 21347 7 1 2 21324 21346
0 21348 5 1 1 21347
0 21349 7 1 2 52616 21348
0 21350 5 1 1 21349
0 21351 7 1 2 52802 74952
0 21352 5 1 1 21351
0 21353 7 1 2 52803 63781
0 21354 5 2 1 21353
0 21355 7 4 2 52126 53487
0 21356 7 1 2 71979 74970
0 21357 5 2 1 21356
0 21358 7 1 2 74968 74974
0 21359 5 1 1 21358
0 21360 7 1 2 74956 21359
0 21361 5 1 1 21360
0 21362 7 2 2 63173 68700
0 21363 7 1 2 73289 74976
0 21364 5 1 1 21363
0 21365 7 1 2 21361 21364
0 21366 7 1 2 21352 21365
0 21367 5 1 1 21366
0 21368 7 1 2 51019 21367
0 21369 5 1 1 21368
0 21370 7 1 2 52804 63727
0 21371 5 1 1 21370
0 21372 7 2 2 67526 68921
0 21373 7 1 2 70427 74978
0 21374 5 1 1 21373
0 21375 7 2 2 51915 50091
0 21376 5 2 1 74980
0 21377 7 1 2 65220 63728
0 21378 7 1 2 74981 21377
0 21379 7 1 2 71448 21378
0 21380 5 1 1 21379
0 21381 7 1 2 21374 21380
0 21382 5 1 1 21381
0 21383 7 1 2 50435 21382
0 21384 5 1 1 21383
0 21385 7 1 2 68672 21384
0 21386 5 1 1 21385
0 21387 7 1 2 52127 74925
0 21388 5 2 1 21387
0 21389 7 1 2 64001 71547
0 21390 7 1 2 74984 21389
0 21391 5 1 1 21390
0 21392 7 1 2 53488 21391
0 21393 7 1 2 21386 21392
0 21394 5 1 1 21393
0 21395 7 1 2 21371 21394
0 21396 7 1 2 21369 21395
0 21397 7 1 2 21350 21396
0 21398 5 1 1 21397
0 21399 7 1 2 53689 21398
0 21400 5 1 1 21399
0 21401 7 2 2 61130 68922
0 21402 5 1 1 74986
0 21403 7 2 2 63174 63508
0 21404 5 1 1 74988
0 21405 7 1 2 21402 21404
0 21406 5 1 1 21405
0 21407 7 1 2 59824 21406
0 21408 5 1 1 21407
0 21409 7 1 2 55890 63556
0 21410 5 1 1 21409
0 21411 7 1 2 21408 21410
0 21412 5 1 1 21411
0 21413 7 1 2 52128 21412
0 21414 5 1 1 21413
0 21415 7 3 2 52617 74286
0 21416 5 4 1 74990
0 21417 7 1 2 60171 69424
0 21418 5 1 1 21417
0 21419 7 1 2 63561 21418
0 21420 5 1 1 21419
0 21421 7 1 2 71013 21420
0 21422 5 1 1 21421
0 21423 7 1 2 74993 21422
0 21424 7 1 2 21414 21423
0 21425 5 1 1 21424
0 21426 7 1 2 72573 21425
0 21427 5 1 1 21426
0 21428 7 1 2 59777 73875
0 21429 5 1 1 21428
0 21430 7 1 2 74948 21429
0 21431 5 1 1 21430
0 21432 7 1 2 51916 21431
0 21433 5 1 1 21432
0 21434 7 1 2 65235 74950
0 21435 7 1 2 21433 21434
0 21436 5 1 1 21435
0 21437 7 1 2 62477 68387
0 21438 7 1 2 21436 21437
0 21439 5 1 1 21438
0 21440 7 1 2 21427 21439
0 21441 5 1 1 21440
0 21442 7 1 2 52805 21441
0 21443 5 1 1 21442
0 21444 7 1 2 21400 21443
0 21445 5 1 1 21444
0 21446 7 1 2 58007 21445
0 21447 5 1 1 21446
0 21448 7 2 2 53489 69653
0 21449 5 1 1 74997
0 21450 7 1 2 55002 74930
0 21451 5 1 1 21450
0 21452 7 2 2 67754 21451
0 21453 7 1 2 74998 74999
0 21454 5 1 1 21453
0 21455 7 1 2 72916 68829
0 21456 7 1 2 74917 21455
0 21457 5 1 1 21456
0 21458 7 1 2 21454 21457
0 21459 5 1 1 21458
0 21460 7 1 2 58757 21459
0 21461 5 1 1 21460
0 21462 7 1 2 73711 75000
0 21463 5 1 1 21462
0 21464 7 1 2 21461 21463
0 21465 5 1 1 21464
0 21466 7 1 2 51317 21465
0 21467 5 1 1 21466
0 21468 7 1 2 69799 73712
0 21469 5 1 1 21468
0 21470 7 5 2 55344 58758
0 21471 7 1 2 69525 75001
0 21472 5 1 1 21471
0 21473 7 1 2 21469 21472
0 21474 5 1 1 21473
0 21475 7 1 2 74911 21474
0 21476 5 1 1 21475
0 21477 7 1 2 55538 21476
0 21478 7 1 2 21467 21477
0 21479 7 1 2 21447 21478
0 21480 5 1 1 21479
0 21481 7 1 2 55891 66167
0 21482 5 2 1 21481
0 21483 7 1 2 72723 75006
0 21484 5 1 1 21483
0 21485 7 1 2 48946 21484
0 21486 5 1 1 21485
0 21487 7 1 2 67847 21486
0 21488 5 1 1 21487
0 21489 7 1 2 74918 21488
0 21490 5 1 1 21489
0 21491 7 1 2 56450 73284
0 21492 5 1 1 21491
0 21493 7 1 2 73510 21492
0 21494 5 1 1 21493
0 21495 7 1 2 49928 21494
0 21496 5 2 1 21495
0 21497 7 1 2 71269 75008
0 21498 7 1 2 21490 21497
0 21499 5 1 1 21498
0 21500 7 1 2 50721 21499
0 21501 5 1 1 21500
0 21502 7 1 2 52129 73873
0 21503 5 1 1 21502
0 21504 7 1 2 66172 21503
0 21505 5 1 1 21504
0 21506 7 1 2 62968 21505
0 21507 5 1 1 21506
0 21508 7 2 2 51318 70736
0 21509 7 1 2 73273 75010
0 21510 5 1 1 21509
0 21511 7 1 2 21507 21510
0 21512 5 1 1 21511
0 21513 7 1 2 49929 21512
0 21514 5 1 1 21513
0 21515 7 1 2 58008 73404
0 21516 5 1 1 21515
0 21517 7 1 2 73586 73723
0 21518 5 1 1 21517
0 21519 7 1 2 21516 21518
0 21520 5 1 1 21519
0 21521 7 1 2 60418 21520
0 21522 5 1 1 21521
0 21523 7 1 2 21514 21522
0 21524 7 1 2 21501 21523
0 21525 5 1 1 21524
0 21526 7 1 2 51020 21525
0 21527 5 1 1 21526
0 21528 7 1 2 50722 21162
0 21529 5 1 1 21528
0 21530 7 1 2 21529 70306
0 21531 5 1 1 21530
0 21532 7 1 2 73602 21531
0 21533 5 1 1 21532
0 21534 7 1 2 70276 72749
0 21535 5 1 1 21534
0 21536 7 1 2 67527 73540
0 21537 7 1 2 21535 21536
0 21538 5 1 1 21537
0 21539 7 1 2 21533 21538
0 21540 5 1 1 21539
0 21541 7 1 2 58009 21540
0 21542 5 1 1 21541
0 21543 7 3 2 50723 58010
0 21544 7 1 2 73929 75012
0 21545 5 1 1 21544
0 21546 7 1 2 73559 75009
0 21547 5 1 1 21546
0 21548 7 1 2 59900 70902
0 21549 7 1 2 21547 21548
0 21550 5 1 1 21549
0 21551 7 1 2 21545 21550
0 21552 5 1 1 21551
0 21553 7 1 2 60336 21552
0 21554 5 1 1 21553
0 21555 7 1 2 56451 60145
0 21556 5 1 1 21555
0 21557 7 2 2 62969 60120
0 21558 5 1 1 75015
0 21559 7 1 2 21556 21558
0 21560 5 1 1 21559
0 21561 7 1 2 50724 60505
0 21562 7 1 2 21560 21561
0 21563 5 1 1 21562
0 21564 7 1 2 69619 72724
0 21565 7 1 2 21563 21564
0 21566 5 1 1 21565
0 21567 7 1 2 69587 21566
0 21568 5 1 1 21567
0 21569 7 1 2 57937 70851
0 21570 5 3 1 21569
0 21571 7 3 2 62970 67884
0 21572 5 2 1 75020
0 21573 7 1 2 75021 71170
0 21574 5 1 1 21573
0 21575 7 1 2 73405 71175
0 21576 5 1 1 21575
0 21577 7 1 2 21574 21576
0 21578 5 1 1 21577
0 21579 7 1 2 75017 21578
0 21580 5 1 1 21579
0 21581 7 1 2 51578 21580
0 21582 7 1 2 21568 21581
0 21583 7 1 2 58759 73347
0 21584 5 2 1 21583
0 21585 7 1 2 53490 73696
0 21586 5 1 1 21585
0 21587 7 1 2 75025 21586
0 21588 5 2 1 21587
0 21589 7 1 2 64017 75027
0 21590 5 1 1 21589
0 21591 7 1 2 53491 71531
0 21592 5 1 1 21591
0 21593 7 1 2 75007 21592
0 21594 5 1 1 21593
0 21595 7 1 2 73541 21594
0 21596 5 1 1 21595
0 21597 7 1 2 70567 75026
0 21598 7 1 2 21596 21597
0 21599 5 1 1 21598
0 21600 7 1 2 687 21599
0 21601 5 1 1 21600
0 21602 7 1 2 21590 21601
0 21603 7 1 2 21582 21602
0 21604 7 1 2 21554 21603
0 21605 7 1 2 21542 21604
0 21606 7 1 2 21527 21605
0 21607 5 1 1 21606
0 21608 7 1 2 21480 21607
0 21609 5 1 1 21608
0 21610 7 1 2 21272 21609
0 21611 5 1 1 21610
0 21612 7 1 2 68269 21611
0 21613 5 1 1 21612
0 21614 7 1 2 21247 21613
0 21615 5 1 1 21614
0 21616 7 1 2 55653 21615
0 21617 5 1 1 21616
0 21618 7 1 2 58011 67186
0 21619 7 1 2 72834 21618
0 21620 5 1 1 21619
0 21621 7 1 2 15547 21620
0 21622 5 1 1 21621
0 21623 7 1 2 55345 21622
0 21624 5 1 1 21623
0 21625 7 2 2 67781 68270
0 21626 7 1 2 67975 75029
0 21627 5 1 1 21626
0 21628 7 1 2 21624 21627
0 21629 5 1 1 21628
0 21630 7 1 2 55654 21629
0 21631 5 1 1 21630
0 21632 7 1 2 73910 21631
0 21633 5 1 1 21632
0 21634 7 1 2 60337 21633
0 21635 5 1 1 21634
0 21636 7 1 2 70326 69753
0 21637 7 1 2 74879 21636
0 21638 7 1 2 73810 21637
0 21639 5 1 1 21638
0 21640 7 1 2 21635 21639
0 21641 5 1 1 21640
0 21642 7 1 2 50725 21641
0 21643 5 1 1 21642
0 21644 7 1 2 52130 73690
0 21645 5 1 1 21644
0 21646 7 1 2 73054 74989
0 21647 7 1 2 67985 21646
0 21648 5 1 1 21647
0 21649 7 1 2 21645 21648
0 21650 5 1 1 21649
0 21651 7 1 2 55539 21650
0 21652 5 1 1 21651
0 21653 7 2 2 52131 70553
0 21654 7 1 2 58012 75031
0 21655 5 1 1 21654
0 21656 7 1 2 59879 71458
0 21657 5 1 1 21656
0 21658 7 1 2 21655 21657
0 21659 5 1 1 21658
0 21660 7 1 2 75030 21659
0 21661 5 1 1 21660
0 21662 7 1 2 21652 21661
0 21663 5 1 1 21662
0 21664 7 1 2 68527 21663
0 21665 5 1 1 21664
0 21666 7 1 2 21643 21665
0 21667 5 1 1 21666
0 21668 7 1 2 51917 21667
0 21669 5 1 1 21668
0 21670 7 1 2 58013 73908
0 21671 5 1 1 21670
0 21672 7 3 2 60267 60537
0 21673 5 1 1 75033
0 21674 7 1 2 66605 75034
0 21675 5 1 1 21674
0 21676 7 1 2 55540 21675
0 21677 5 1 1 21676
0 21678 7 1 2 74934 21677
0 21679 5 1 1 21678
0 21680 7 1 2 53492 67782
0 21681 5 2 1 21680
0 21682 7 5 2 60198 66097
0 21683 7 1 2 68830 75038
0 21684 5 1 1 21683
0 21685 7 1 2 75036 21684
0 21686 5 1 1 21685
0 21687 7 1 2 73097 21686
0 21688 5 1 1 21687
0 21689 7 1 2 73630 70459
0 21690 5 1 1 21689
0 21691 7 1 2 53690 71671
0 21692 5 1 1 21691
0 21693 7 1 2 21690 21692
0 21694 5 1 1 21693
0 21695 7 1 2 55003 21694
0 21696 5 1 1 21695
0 21697 7 1 2 21688 21696
0 21698 5 1 1 21697
0 21699 7 1 2 58760 21698
0 21700 5 1 1 21699
0 21701 7 1 2 70414 73728
0 21702 5 1 1 21701
0 21703 7 1 2 66762 75039
0 21704 5 1 1 21703
0 21705 7 1 2 21702 21704
0 21706 5 1 1 21705
0 21707 7 1 2 71532 21706
0 21708 5 1 1 21707
0 21709 7 2 2 55004 75040
0 21710 7 1 2 73655 75043
0 21711 5 1 1 21710
0 21712 7 2 2 72883 68294
0 21713 5 1 1 75045
0 21714 7 2 2 52132 53691
0 21715 7 1 2 66249 75047
0 21716 7 1 2 75046 21715
0 21717 5 1 1 21716
0 21718 7 1 2 21711 21717
0 21719 7 1 2 21708 21718
0 21720 7 1 2 21700 21719
0 21721 7 1 2 21679 21720
0 21722 5 1 1 21721
0 21723 7 1 2 50068 21722
0 21724 5 1 1 21723
0 21725 7 3 2 63488 67835
0 21726 7 1 2 53792 68887
0 21727 7 1 2 75049 21726
0 21728 5 1 1 21727
0 21729 7 1 2 21724 21728
0 21730 5 1 1 21729
0 21731 7 1 2 49079 21730
0 21732 5 1 1 21731
0 21733 7 1 2 48947 73103
0 21734 5 1 1 21733
0 21735 7 1 2 63479 21734
0 21736 5 1 1 21735
0 21737 7 1 2 72905 21736
0 21738 5 1 1 21737
0 21739 7 1 2 73098 70558
0 21740 5 1 1 21739
0 21741 7 1 2 70023 21740
0 21742 5 1 1 21741
0 21743 7 1 2 68271 21742
0 21744 5 1 1 21743
0 21745 7 1 2 21738 21744
0 21746 5 1 1 21745
0 21747 7 1 2 66421 21746
0 21748 5 1 1 21747
0 21749 7 1 2 60199 67885
0 21750 7 1 2 72603 21749
0 21751 7 1 2 73105 21750
0 21752 5 1 1 21751
0 21753 7 1 2 21748 21752
0 21754 5 1 1 21753
0 21755 7 1 2 58014 21754
0 21756 5 1 1 21755
0 21757 7 1 2 72304 72182
0 21758 7 1 2 75044 21757
0 21759 5 1 1 21758
0 21760 7 1 2 21756 21759
0 21761 7 1 2 21732 21760
0 21762 5 1 1 21761
0 21763 7 1 2 55655 21762
0 21764 5 1 1 21763
0 21765 7 1 2 21671 21764
0 21766 7 1 2 21669 21765
0 21767 5 1 1 21766
0 21768 7 1 2 57602 21767
0 21769 5 1 1 21768
0 21770 7 2 2 65106 73697
0 21771 5 1 1 75052
0 21772 7 1 2 68794 73628
0 21773 5 1 1 21772
0 21774 7 1 2 55892 21773
0 21775 5 1 1 21774
0 21776 7 1 2 67893 21775
0 21777 5 1 1 21776
0 21778 7 1 2 65003 21777
0 21779 5 1 1 21778
0 21780 7 1 2 21771 21779
0 21781 5 1 1 21780
0 21782 7 1 2 51918 21781
0 21783 5 1 1 21782
0 21784 7 1 2 68791 70848
0 21785 5 1 1 21784
0 21786 7 1 2 71533 70849
0 21787 5 1 1 21786
0 21788 7 1 2 53493 75011
0 21789 5 1 1 21788
0 21790 7 1 2 21787 21789
0 21791 5 1 1 21790
0 21792 7 1 2 49930 21791
0 21793 5 1 1 21792
0 21794 7 1 2 21785 21793
0 21795 7 1 2 21783 21794
0 21796 5 1 1 21795
0 21797 7 1 2 51579 21796
0 21798 5 1 1 21797
0 21799 7 1 2 66422 73713
0 21800 5 1 1 21799
0 21801 7 2 2 60597 73355
0 21802 5 1 1 75054
0 21803 7 1 2 75053 75055
0 21804 5 1 1 21803
0 21805 7 1 2 21800 21804
0 21806 5 1 1 21805
0 21807 7 1 2 53494 21806
0 21808 5 1 1 21807
0 21809 7 1 2 21798 21808
0 21810 5 1 1 21809
0 21811 7 1 2 51021 21810
0 21812 5 1 1 21811
0 21813 7 1 2 71322 69721
0 21814 5 1 1 21813
0 21815 7 1 2 75037 21814
0 21816 5 1 1 21815
0 21817 7 1 2 51919 21816
0 21818 5 1 1 21817
0 21819 7 1 2 52133 60538
0 21820 7 1 2 73639 21819
0 21821 5 1 1 21820
0 21822 7 1 2 21818 21821
0 21823 5 1 1 21822
0 21824 7 1 2 71534 21823
0 21825 5 1 1 21824
0 21826 7 4 2 52618 53282
0 21827 5 3 1 75056
0 21828 7 4 2 71284 75057
0 21829 7 2 2 73491 75063
0 21830 7 1 2 69722 75067
0 21831 5 1 1 21830
0 21832 7 3 2 48948 68855
0 21833 5 1 1 75069
0 21834 7 1 2 53495 75070
0 21835 5 1 1 21834
0 21836 7 1 2 21831 21835
0 21837 5 1 1 21836
0 21838 7 1 2 51920 21837
0 21839 5 1 1 21838
0 21840 7 1 2 66423 73656
0 21841 5 1 1 21840
0 21842 7 1 2 73792 21841
0 21843 5 1 1 21842
0 21844 7 1 2 63657 70415
0 21845 7 1 2 21843 21844
0 21846 5 1 1 21845
0 21847 7 1 2 21839 21846
0 21848 7 1 2 21825 21847
0 21849 5 1 1 21848
0 21850 7 1 2 50196 21849
0 21851 5 1 1 21850
0 21852 7 1 2 73151 69710
0 21853 7 1 2 73714 21852
0 21854 5 1 1 21853
0 21855 7 1 2 21851 21854
0 21856 7 1 2 21812 21855
0 21857 5 1 1 21856
0 21858 7 1 2 50069 21857
0 21859 5 1 1 21858
0 21860 7 2 2 66894 71598
0 21861 5 1 1 75072
0 21862 7 1 2 52134 21861
0 21863 5 1 1 21862
0 21864 7 1 2 71569 21863
0 21865 5 1 1 21864
0 21866 7 1 2 51921 21865
0 21867 5 1 1 21866
0 21868 7 1 2 73637 21867
0 21869 5 1 1 21868
0 21870 7 1 2 73729 21869
0 21871 5 1 1 21870
0 21872 7 1 2 73455 69723
0 21873 5 1 1 21872
0 21874 7 1 2 73554 71306
0 21875 5 1 1 21874
0 21876 7 1 2 21873 21875
0 21877 5 1 1 21876
0 21878 7 1 2 52806 21877
0 21879 5 1 1 21878
0 21880 7 2 2 73369 69711
0 21881 7 1 2 53496 75074
0 21882 5 1 1 21881
0 21883 7 1 2 59934 71672
0 21884 5 1 1 21883
0 21885 7 1 2 21882 21884
0 21886 5 1 1 21885
0 21887 7 1 2 66763 21886
0 21888 5 1 1 21887
0 21889 7 1 2 21879 21888
0 21890 7 1 2 21871 21889
0 21891 5 1 1 21890
0 21892 7 1 2 50070 21891
0 21893 5 1 1 21892
0 21894 7 1 2 66432 73161
0 21895 5 1 1 21894
0 21896 7 2 2 51319 59901
0 21897 7 1 2 60338 75076
0 21898 7 1 2 70585 21897
0 21899 5 1 1 21898
0 21900 7 1 2 21895 21899
0 21901 5 1 1 21900
0 21902 7 1 2 50071 21901
0 21903 5 1 1 21902
0 21904 7 1 2 69902 73682
0 21905 5 1 1 21904
0 21906 7 1 2 21903 21905
0 21907 5 1 1 21906
0 21908 7 1 2 50726 21907
0 21909 5 1 1 21908
0 21910 7 2 2 59935 63729
0 21911 5 1 1 75078
0 21912 7 1 2 70460 75079
0 21913 5 1 1 21912
0 21914 7 1 2 50436 60146
0 21915 7 1 2 73730 21914
0 21916 5 1 1 21915
0 21917 7 1 2 21913 21916
0 21918 5 1 1 21917
0 21919 7 1 2 69448 21918
0 21920 5 1 1 21919
0 21921 7 1 2 21909 21920
0 21922 5 1 1 21921
0 21923 7 1 2 55893 21922
0 21924 5 1 1 21923
0 21925 7 1 2 55005 21673
0 21926 5 2 1 21925
0 21927 7 1 2 69464 72134
0 21928 5 1 1 21927
0 21929 7 1 2 73564 69433
0 21930 5 1 1 21929
0 21931 7 1 2 21928 21930
0 21932 5 1 1 21931
0 21933 7 1 2 49931 21932
0 21934 5 1 1 21933
0 21935 7 4 2 50072 69526
0 21936 7 1 2 66424 75082
0 21937 5 1 1 21936
0 21938 7 1 2 21934 21937
0 21939 5 1 1 21938
0 21940 7 1 2 75080 21939
0 21941 5 1 1 21940
0 21942 7 1 2 21924 21941
0 21943 7 1 2 21893 21942
0 21944 5 1 1 21943
0 21945 7 1 2 58761 21944
0 21946 5 1 1 21945
0 21947 7 1 2 73333 68923
0 21948 5 1 1 21947
0 21949 7 1 2 68924 74971
0 21950 5 1 1 21949
0 21951 7 1 2 21911 21950
0 21952 5 1 1 21951
0 21953 7 1 2 55894 21952
0 21954 5 1 1 21953
0 21955 7 1 2 14050 21954
0 21956 7 1 2 21948 21955
0 21957 5 1 1 21956
0 21958 7 1 2 69945 72135
0 21959 7 1 2 21957 21958
0 21960 5 1 1 21959
0 21961 7 1 2 21946 21960
0 21962 7 1 2 21859 21961
0 21963 5 1 1 21962
0 21964 7 1 2 49080 21963
0 21965 5 1 1 21964
0 21966 7 1 2 50437 72956
0 21967 5 1 1 21966
0 21968 7 1 2 15685 21967
0 21969 5 1 1 21968
0 21970 7 1 2 70416 21969
0 21971 5 1 1 21970
0 21972 7 1 2 72945 21971
0 21973 5 1 1 21972
0 21974 7 1 2 58762 21973
0 21975 5 1 1 21974
0 21976 7 1 2 70737 70417
0 21977 5 1 1 21976
0 21978 7 1 2 55006 21977
0 21979 5 2 1 21978
0 21980 7 1 2 63421 75086
0 21981 5 1 1 21980
0 21982 7 1 2 21975 21981
0 21983 5 1 1 21982
0 21984 7 1 2 55346 21983
0 21985 5 1 1 21984
0 21986 7 1 2 63493 72672
0 21987 5 1 1 21986
0 21988 7 1 2 21985 21987
0 21989 5 1 1 21988
0 21990 7 1 2 73684 21989
0 21991 5 1 1 21990
0 21992 7 1 2 21965 21991
0 21993 5 1 1 21992
0 21994 7 1 2 55656 21993
0 21995 5 1 1 21994
0 21996 7 1 2 73707 75087
0 21997 5 1 1 21996
0 21998 7 2 2 48949 67808
0 21999 5 2 1 75088
0 22000 7 7 2 52619 55541
0 22001 7 1 2 73147 68602
0 22002 5 5 1 22001
0 22003 7 1 2 75092 75099
0 22004 5 1 1 22003
0 22005 7 1 2 75090 22004
0 22006 5 1 1 22005
0 22007 7 1 2 53692 22006
0 22008 5 1 1 22007
0 22009 7 1 2 55895 66425
0 22010 7 1 2 69242 22009
0 22011 5 1 1 22010
0 22012 7 1 2 75023 22011
0 22013 5 1 1 22012
0 22014 7 1 2 52807 22013
0 22015 5 1 1 22014
0 22016 7 1 2 22008 22015
0 22017 5 1 1 22016
0 22018 7 1 2 60147 22017
0 22019 5 1 1 22018
0 22020 7 1 2 66426 70559
0 22021 5 1 1 22020
0 22022 7 1 2 73793 22021
0 22023 5 1 1 22022
0 22024 7 1 2 61498 22023
0 22025 5 1 1 22024
0 22026 7 1 2 22019 22025
0 22027 5 1 1 22026
0 22028 7 1 2 50438 22027
0 22029 5 1 1 22028
0 22030 7 1 2 59742 66279
0 22031 7 1 2 70656 22030
0 22032 5 1 1 22031
0 22033 7 1 2 64374 22032
0 22034 5 1 1 22033
0 22035 7 1 2 49932 22034
0 22036 5 1 1 22035
0 22037 7 1 2 68795 22036
0 22038 5 1 1 22037
0 22039 7 1 2 51580 22038
0 22040 5 1 1 22039
0 22041 7 12 2 52620 55347
0 22042 5 2 1 75104
0 22043 7 2 2 75105 72563
0 22044 7 1 2 59021 75118
0 22045 5 1 1 22044
0 22046 7 1 2 73565 70548
0 22047 5 1 1 22046
0 22048 7 1 2 22045 22047
0 22049 5 1 1 22048
0 22050 7 1 2 69654 22049
0 22051 5 1 1 22050
0 22052 7 1 2 55348 68722
0 22053 7 1 2 72564 22052
0 22054 5 1 1 22053
0 22055 7 1 2 22051 22054
0 22056 5 1 1 22055
0 22057 7 1 2 55542 22056
0 22058 5 1 1 22057
0 22059 7 1 2 22040 22058
0 22060 7 1 2 22029 22059
0 22061 5 1 1 22060
0 22062 7 1 2 51022 22061
0 22063 5 1 1 22062
0 22064 7 1 2 59936 73796
0 22065 5 1 1 22064
0 22066 7 1 2 70738 73603
0 22067 5 1 1 22066
0 22068 7 1 2 75024 22067
0 22069 5 1 1 22068
0 22070 7 1 2 51581 22069
0 22071 5 1 1 22070
0 22072 7 1 2 55543 60200
0 22073 7 1 2 73056 22072
0 22074 7 1 2 70059 22073
0 22075 5 1 1 22074
0 22076 7 1 2 22071 22075
0 22077 5 1 1 22076
0 22078 7 1 2 70418 22077
0 22079 5 1 1 22078
0 22080 7 1 2 22065 22079
0 22081 7 1 2 22063 22080
0 22082 5 1 1 22081
0 22083 7 1 2 68272 22082
0 22084 5 1 1 22083
0 22085 7 1 2 60569 15841
0 22086 5 1 1 22085
0 22087 7 1 2 51023 22086
0 22088 5 1 1 22087
0 22089 7 1 2 63679 22088
0 22090 5 1 1 22089
0 22091 7 1 2 48950 22090
0 22092 5 1 1 22091
0 22093 7 6 2 49741 50197
0 22094 5 2 1 75120
0 22095 7 2 2 52621 75121
0 22096 7 1 2 63452 75128
0 22097 5 1 1 22096
0 22098 7 1 2 22092 22097
0 22099 5 1 1 22098
0 22100 7 1 2 51922 22099
0 22101 5 1 1 22100
0 22102 7 1 2 51024 72937
0 22103 5 1 1 22102
0 22104 7 1 2 22101 22103
0 22105 5 1 1 22104
0 22106 7 1 2 73811 22105
0 22107 5 1 1 22106
0 22108 7 1 2 22084 22107
0 22109 5 1 1 22108
0 22110 7 1 2 55657 22109
0 22111 5 1 1 22110
0 22112 7 1 2 73617 73670
0 22113 7 1 2 72056 22112
0 22114 5 1 1 22113
0 22115 7 1 2 22111 22114
0 22116 5 1 1 22115
0 22117 7 1 2 58015 22116
0 22118 5 1 1 22117
0 22119 7 1 2 21997 22118
0 22120 7 1 2 21995 22119
0 22121 7 1 2 21769 22120
0 22122 5 1 1 22121
0 22123 7 1 2 59857 22122
0 22124 5 1 1 22123
0 22125 7 1 2 50198 59557
0 22126 5 3 1 22125
0 22127 7 1 2 70191 75130
0 22128 5 1 1 22127
0 22129 7 1 2 67730 22128
0 22130 5 1 1 22129
0 22131 7 1 2 53497 74919
0 22132 5 1 1 22131
0 22133 7 1 2 22130 22132
0 22134 5 1 1 22133
0 22135 7 1 2 50727 22134
0 22136 5 1 1 22135
0 22137 7 3 2 58016 65679
0 22138 5 1 1 75133
0 22139 7 1 2 55691 73693
0 22140 5 2 1 22139
0 22141 7 1 2 49742 75136
0 22142 5 1 1 22141
0 22143 7 1 2 75134 22142
0 22144 5 1 1 22143
0 22145 7 1 2 59361 22144
0 22146 7 1 2 22136 22145
0 22147 5 1 1 22146
0 22148 7 1 2 48951 22147
0 22149 5 1 1 22148
0 22150 7 1 2 63476 75135
0 22151 5 1 1 22150
0 22152 7 1 2 55007 71562
0 22153 5 4 1 22152
0 22154 7 1 2 48952 75138
0 22155 5 1 1 22154
0 22156 7 1 2 52135 62607
0 22157 5 2 1 22156
0 22158 7 3 2 50092 63175
0 22159 7 1 2 60165 75144
0 22160 5 1 1 22159
0 22161 7 1 2 75142 22160
0 22162 5 1 1 22161
0 22163 7 1 2 51923 22162
0 22164 5 1 1 22163
0 22165 7 1 2 56626 62608
0 22166 5 2 1 22165
0 22167 7 1 2 22164 75147
0 22168 5 1 1 22167
0 22169 7 1 2 49743 68925
0 22170 7 1 2 22168 22169
0 22171 5 1 1 22170
0 22172 7 1 2 22155 22171
0 22173 5 1 1 22172
0 22174 7 1 2 58763 22173
0 22175 5 1 1 22174
0 22176 7 1 2 22151 22175
0 22177 7 1 2 22149 22176
0 22178 5 1 1 22177
0 22179 7 1 2 55349 22178
0 22180 5 1 1 22179
0 22181 7 1 2 54646 60465
0 22182 5 2 1 22181
0 22183 7 1 2 63494 75149
0 22184 5 1 1 22183
0 22185 7 1 2 22180 22184
0 22186 5 1 1 22185
0 22187 7 1 2 73853 22186
0 22188 5 1 1 22187
0 22189 7 1 2 64387 74920
0 22190 5 1 1 22189
0 22191 7 1 2 72579 22190
0 22192 5 1 1 22191
0 22193 7 1 2 49933 22192
0 22194 5 1 1 22193
0 22195 7 1 2 73337 74921
0 22196 5 1 1 22195
0 22197 7 1 2 22194 22196
0 22198 5 1 1 22197
0 22199 7 1 2 50728 22198
0 22200 5 1 1 22199
0 22201 7 1 2 705 75022
0 22202 5 1 1 22201
0 22203 7 1 2 22200 22202
0 22204 5 1 1 22203
0 22205 7 1 2 58017 22204
0 22206 5 1 1 22205
0 22207 7 1 2 60173 71545
0 22208 5 1 1 22207
0 22209 7 2 2 58018 60148
0 22210 5 1 1 75151
0 22211 7 1 2 51320 70352
0 22212 7 1 2 75152 22211
0 22213 5 1 1 22212
0 22214 7 1 2 22208 22213
0 22215 5 1 1 22214
0 22216 7 1 2 50729 22215
0 22217 5 1 1 22216
0 22218 7 1 2 60237 74985
0 22219 5 1 1 22218
0 22220 7 1 2 73724 22219
0 22221 5 1 1 22220
0 22222 7 1 2 73858 71218
0 22223 7 1 2 75032 22222
0 22224 5 1 1 22223
0 22225 7 1 2 22221 22224
0 22226 7 1 2 22217 22225
0 22227 5 1 1 22226
0 22228 7 1 2 49934 22227
0 22229 5 1 1 22228
0 22230 7 1 2 62971 73865
0 22231 5 1 1 22230
0 22232 7 1 2 51321 73870
0 22233 5 1 1 22232
0 22234 7 1 2 64388 63607
0 22235 5 1 1 22234
0 22236 7 1 2 22233 22235
0 22237 7 1 2 22231 22236
0 22238 5 1 1 22237
0 22239 7 1 2 49935 22238
0 22240 5 1 1 22239
0 22241 7 1 2 50730 71295
0 22242 5 1 1 22241
0 22243 7 1 2 22240 22242
0 22244 5 1 1 22243
0 22245 7 1 2 61486 22244
0 22246 5 1 1 22245
0 22247 7 6 2 52957 49744
0 22248 7 2 2 52885 75153
0 22249 7 1 2 50093 69510
0 22250 7 1 2 75159 22249
0 22251 5 1 1 22250
0 22252 7 1 2 10338 22251
0 22253 5 1 1 22252
0 22254 7 1 2 68718 22253
0 22255 5 1 1 22254
0 22256 7 2 2 48604 60809
0 22257 5 1 1 75161
0 22258 7 1 2 49540 75162
0 22259 5 1 1 22258
0 22260 7 1 2 73406 22259
0 22261 5 1 1 22260
0 22262 7 1 2 22255 22261
0 22263 7 1 2 22246 22262
0 22264 7 1 2 22229 22263
0 22265 5 1 1 22264
0 22266 7 1 2 51025 22265
0 22267 5 1 1 22266
0 22268 7 1 2 65680 75028
0 22269 5 1 1 22268
0 22270 7 1 2 51582 22269
0 22271 7 1 2 22267 22270
0 22272 7 1 2 22206 22271
0 22273 5 1 1 22272
0 22274 7 2 2 52622 53693
0 22275 7 1 2 64489 68583
0 22276 5 1 1 22275
0 22277 7 4 2 50094 60268
0 22278 5 1 1 75165
0 22279 7 4 2 60166 75166
0 22280 7 1 2 69800 75169
0 22281 5 1 1 22280
0 22282 7 1 2 22276 22281
0 22283 5 1 1 22282
0 22284 7 1 2 50439 22283
0 22285 5 1 1 22284
0 22286 7 1 2 60339 63796
0 22287 5 1 1 22286
0 22288 7 1 2 22285 22287
0 22289 5 1 1 22288
0 22290 7 1 2 75163 22289
0 22291 5 1 1 22290
0 22292 7 1 2 50731 66475
0 22293 5 1 1 22292
0 22294 7 1 2 74975 22293
0 22295 5 1 1 22294
0 22296 7 1 2 52808 22295
0 22297 5 1 1 22296
0 22298 7 2 2 52623 69655
0 22299 5 1 1 75173
0 22300 7 1 2 74960 75174
0 22301 5 1 1 22300
0 22302 7 1 2 68750 74958
0 22303 5 1 1 22302
0 22304 7 1 2 22301 22303
0 22305 7 1 2 22297 22304
0 22306 5 1 1 22305
0 22307 7 1 2 74926 22306
0 22308 5 1 1 22307
0 22309 7 1 2 65108 60810
0 22310 5 2 1 22309
0 22311 7 1 2 68666 69243
0 22312 7 1 2 75175 22311
0 22313 5 1 1 22312
0 22314 7 1 2 22308 22313
0 22315 7 1 2 22291 22314
0 22316 5 1 1 22315
0 22317 7 1 2 51026 22316
0 22318 5 1 1 22317
0 22319 7 1 2 65681 68667
0 22320 7 1 2 68489 22319
0 22321 5 1 1 22320
0 22322 7 1 2 22318 22321
0 22323 5 1 1 22322
0 22324 7 1 2 58019 22323
0 22325 5 1 1 22324
0 22326 7 1 2 73924 74943
0 22327 5 1 1 22326
0 22328 7 1 2 56730 60138
0 22329 5 1 1 22328
0 22330 7 1 2 68668 22329
0 22331 5 1 1 22330
0 22332 7 2 2 50095 66606
0 22333 7 1 2 60149 75160
0 22334 7 1 2 75177 22333
0 22335 5 1 1 22334
0 22336 7 1 2 22331 22335
0 22337 5 1 1 22336
0 22338 7 1 2 60539 22337
0 22339 5 1 1 22338
0 22340 7 1 2 52809 68388
0 22341 5 1 1 22340
0 22342 7 1 2 52136 73925
0 22343 5 1 1 22342
0 22344 7 1 2 74969 22343
0 22345 5 1 1 22344
0 22346 7 1 2 74954 22345
0 22347 5 1 1 22346
0 22348 7 1 2 22341 22347
0 22349 7 1 2 22339 22348
0 22350 7 1 2 22327 22349
0 22351 5 1 1 22350
0 22352 7 1 2 53694 22351
0 22353 5 1 1 22352
0 22354 7 6 2 52810 53498
0 22355 5 2 1 75179
0 22356 7 1 2 63730 75180
0 22357 7 1 2 75150 22356
0 22358 5 1 1 22357
0 22359 7 1 2 22353 22358
0 22360 5 1 1 22359
0 22361 7 1 2 58764 22360
0 22362 5 1 1 22361
0 22363 7 1 2 59778 63731
0 22364 5 1 1 22363
0 22365 7 2 2 52137 63797
0 22366 5 1 1 75187
0 22367 7 1 2 22364 22366
0 22368 5 1 1 22367
0 22369 7 1 2 51924 22368
0 22370 5 1 1 22369
0 22371 7 1 2 52958 75188
0 22372 5 1 1 22371
0 22373 7 1 2 22370 22372
0 22374 5 1 1 22373
0 22375 7 1 2 50440 22374
0 22376 5 1 1 22375
0 22377 7 2 2 50199 9388
0 22378 7 2 2 55008 73370
0 22379 5 1 1 75191
0 22380 7 1 2 63802 22379
0 22381 5 1 1 22380
0 22382 7 1 2 75189 22381
0 22383 5 1 1 22382
0 22384 7 2 2 53499 68389
0 22385 5 2 1 75193
0 22386 7 1 2 73132 75195
0 22387 7 1 2 22383 22386
0 22388 7 1 2 22376 22387
0 22389 5 1 1 22388
0 22390 7 1 2 73715 22389
0 22391 5 1 1 22390
0 22392 7 1 2 55544 22391
0 22393 7 1 2 22362 22392
0 22394 7 1 2 22325 22393
0 22395 5 1 1 22394
0 22396 7 1 2 22273 22395
0 22397 5 1 1 22396
0 22398 7 1 2 64490 74940
0 22399 5 1 1 22398
0 22400 7 6 2 50732 60150
0 22401 5 1 1 75197
0 22402 7 1 2 59779 75198
0 22403 7 1 2 74935 22402
0 22404 5 1 1 22403
0 22405 7 1 2 22399 22404
0 22406 5 1 1 22405
0 22407 7 1 2 66724 22406
0 22408 5 1 1 22407
0 22409 7 1 2 22397 22408
0 22410 5 1 1 22409
0 22411 7 1 2 68273 22410
0 22412 5 1 1 22411
0 22413 7 1 2 22188 22412
0 22414 5 1 1 22413
0 22415 7 1 2 55658 22414
0 22416 5 1 1 22415
0 22417 7 1 2 55009 22138
0 22418 7 1 2 21253 22417
0 22419 5 1 1 22418
0 22420 7 1 2 73708 22419
0 22421 5 1 1 22420
0 22422 7 1 2 22416 22421
0 22423 5 1 1 22422
0 22424 7 1 2 57603 22423
0 22425 5 1 1 22424
0 22426 7 1 2 57938 74904
0 22427 5 1 1 22426
0 22428 7 1 2 50733 22427
0 22429 5 1 1 22428
0 22430 7 1 2 60363 74923
0 22431 5 1 1 22430
0 22432 7 1 2 58020 22431
0 22433 5 1 1 22432
0 22434 7 1 2 55896 75176
0 22435 5 1 1 22434
0 22436 7 1 2 74884 22435
0 22437 7 1 2 22433 22436
0 22438 7 1 2 22429 22437
0 22439 5 1 1 22438
0 22440 7 1 2 73709 22439
0 22441 5 1 1 22440
0 22442 7 1 2 22425 22441
0 22443 7 1 2 22124 22442
0 22444 7 1 2 21617 22443
0 22445 5 1 1 22444
0 22446 7 1 2 57009 22445
0 22447 5 1 1 22446
0 22448 7 1 2 21103 22447
0 22449 7 1 2 19145 22448
0 22450 7 1 2 14108 22449
0 22451 7 1 2 7402 22450
0 22452 5 1 1 22451
0 22453 7 1 2 51830 22452
0 22454 5 1 1 22453
0 22455 7 1 2 63928 62078
0 22456 5 2 1 22455
0 22457 7 1 2 52138 60665
0 22458 5 2 1 22457
0 22459 7 2 2 75203 75205
0 22460 5 7 1 75207
0 22461 7 2 2 59656 75209
0 22462 5 1 1 75216
0 22463 7 1 2 52139 70978
0 22464 5 1 1 22463
0 22465 7 1 2 50200 70298
0 22466 5 1 1 22465
0 22467 7 1 2 70976 22466
0 22468 5 1 1 22467
0 22469 7 2 2 20064 22468
0 22470 5 1 1 75218
0 22471 7 1 2 22464 22470
0 22472 5 1 1 22471
0 22473 7 1 2 51925 22472
0 22474 5 1 1 22473
0 22475 7 2 2 74395 69158
0 22476 5 1 1 75220
0 22477 7 1 2 53090 75221
0 22478 5 1 1 22477
0 22479 7 1 2 60201 61182
0 22480 5 1 1 22479
0 22481 7 1 2 22478 22480
0 22482 7 1 2 22474 22481
0 22483 5 2 1 22482
0 22484 7 1 2 52284 75222
0 22485 5 1 1 22484
0 22486 7 1 2 22462 22485
0 22487 5 1 1 22486
0 22488 7 9 2 52486 49541
0 22489 5 3 1 75224
0 22490 7 11 2 48750 53283
0 22491 5 9 1 75236
0 22492 7 1 2 75233 75247
0 22493 5 7 1 22492
0 22494 7 2 2 59140 75154
0 22495 5 1 1 75263
0 22496 7 2 2 75256 75264
0 22497 5 1 1 75265
0 22498 7 4 2 61443 63214
0 22499 5 26 1 75267
0 22500 7 2 2 73768 75271
0 22501 5 1 1 75297
0 22502 7 1 2 22497 22501
0 22503 5 1 1 22502
0 22504 7 1 2 51583 22503
0 22505 5 1 1 22504
0 22506 7 5 2 52487 52959
0 22507 5 1 1 75299
0 22508 7 3 2 75058 75300
0 22509 7 4 2 59022 66296
0 22510 7 1 2 75304 75307
0 22511 5 1 1 22510
0 22512 7 1 2 22505 22511
0 22513 5 1 1 22512
0 22514 7 1 2 22487 22513
0 22515 5 1 1 22514
0 22516 7 3 2 48751 50734
0 22517 5 1 1 75311
0 22518 7 1 2 58428 70731
0 22519 5 1 1 22518
0 22520 7 1 2 59832 22519
0 22521 5 1 1 22520
0 22522 7 1 2 52140 22521
0 22523 5 1 1 22522
0 22524 7 3 2 59836 62148
0 22525 5 2 1 75314
0 22526 7 1 2 55897 75317
0 22527 5 1 1 22526
0 22528 7 1 2 56095 61283
0 22529 5 1 1 22528
0 22530 7 2 2 57604 22529
0 22531 7 1 2 50201 75319
0 22532 5 1 1 22531
0 22533 7 1 2 22527 22532
0 22534 7 2 2 22523 22533
0 22535 5 1 1 75321
0 22536 7 2 2 58683 22535
0 22537 5 1 1 75323
0 22538 7 1 2 22517 22537
0 22539 5 1 1 22538
0 22540 7 1 2 51027 22539
0 22541 5 1 1 22540
0 22542 7 1 2 62260 72893
0 22543 5 1 1 22542
0 22544 7 1 2 57605 22543
0 22545 5 1 1 22544
0 22546 7 2 2 56096 22545
0 22547 5 1 1 75325
0 22548 7 2 2 70075 22547
0 22549 5 1 1 75327
0 22550 7 1 2 75208 22549
0 22551 5 1 1 22550
0 22552 7 1 2 52960 65230
0 22553 5 1 1 22552
0 22554 7 1 2 55010 22553
0 22555 5 5 1 22554
0 22556 7 4 2 52624 51028
0 22557 5 4 1 75334
0 22558 7 1 2 50441 75338
0 22559 7 1 2 75329 22558
0 22560 7 1 2 22551 22559
0 22561 5 1 1 22560
0 22562 7 1 2 22541 22561
0 22563 5 1 1 22562
0 22564 7 1 2 53284 22563
0 22565 5 1 1 22564
0 22566 7 7 2 51926 49542
0 22567 7 1 2 62096 75342
0 22568 7 1 2 71368 22567
0 22569 7 1 2 72758 22568
0 22570 5 1 1 22569
0 22571 7 1 2 22565 22570
0 22572 5 1 1 22571
0 22573 7 1 2 52488 22572
0 22574 5 1 1 22573
0 22575 7 1 2 53091 72690
0 22576 7 1 2 75237 22575
0 22577 7 8 2 50096 59880
0 22578 5 1 1 75349
0 22579 7 1 2 70316 75350
0 22580 7 1 2 22576 22579
0 22581 5 1 1 22580
0 22582 7 1 2 22574 22581
0 22583 5 1 1 22582
0 22584 7 1 2 49745 22583
0 22585 5 1 1 22584
0 22586 7 6 2 49543 50735
0 22587 5 3 1 75357
0 22588 7 1 2 57606 59858
0 22589 5 2 1 22588
0 22590 7 1 2 48177 75366
0 22591 5 1 1 22590
0 22592 7 1 2 57501 59785
0 22593 5 3 1 22592
0 22594 7 1 2 51927 75368
0 22595 7 1 2 22591 22594
0 22596 5 1 1 22595
0 22597 7 1 2 70653 22596
0 22598 5 1 1 22597
0 22599 7 1 2 50202 22598
0 22600 5 1 1 22599
0 22601 7 1 2 53092 59859
0 22602 5 1 1 22601
0 22603 7 1 2 48178 22602
0 22604 5 1 1 22603
0 22605 7 1 2 72670 22604
0 22606 5 1 1 22605
0 22607 7 1 2 71443 22606
0 22608 7 2 2 22600 22607
0 22609 5 1 1 75371
0 22610 7 1 2 58684 22609
0 22611 5 1 1 22610
0 22612 7 1 2 75363 22611
0 22613 5 1 1 22612
0 22614 7 1 2 51029 22613
0 22615 5 1 1 22614
0 22616 7 4 2 49544 50442
0 22617 5 1 1 75373
0 22618 7 1 2 70204 75374
0 22619 5 1 1 22618
0 22620 7 1 2 57607 73598
0 22621 5 1 1 22620
0 22622 7 1 2 61686 22621
0 22623 5 1 1 22622
0 22624 7 1 2 58685 22623
0 22625 5 1 1 22624
0 22626 7 1 2 22619 22625
0 22627 5 1 1 22626
0 22628 7 1 2 51030 22627
0 22629 5 1 1 22628
0 22630 7 1 2 61044 68926
0 22631 7 1 2 75018 22630
0 22632 5 1 1 22631
0 22633 7 1 2 22629 22632
0 22634 5 1 1 22633
0 22635 7 1 2 58429 22634
0 22636 5 1 1 22635
0 22637 7 1 2 57608 65826
0 22638 5 2 1 22637
0 22639 7 1 2 62666 75377
0 22640 5 1 1 22639
0 22641 7 1 2 67326 22640
0 22642 5 1 1 22641
0 22643 7 1 2 60716 75206
0 22644 7 1 2 22642 22643
0 22645 5 1 1 22644
0 22646 7 1 2 50443 71117
0 22647 7 1 2 75330 22646
0 22648 7 1 2 22645 22647
0 22649 5 1 1 22648
0 22650 7 4 2 52489 73199
0 22651 5 5 1 75379
0 22652 7 1 2 71167 70852
0 22653 5 1 1 22652
0 22654 7 2 2 62324 55753
0 22655 5 3 1 75388
0 22656 7 1 2 22653 75390
0 22657 5 1 1 22656
0 22658 7 1 2 55011 22657
0 22659 5 1 1 22658
0 22660 7 1 2 58021 67755
0 22661 7 1 2 22659 22660
0 22662 5 1 1 22661
0 22663 7 1 2 75383 22662
0 22664 7 1 2 22649 22663
0 22665 7 1 2 22636 22664
0 22666 7 1 2 22615 22665
0 22667 5 1 1 22666
0 22668 7 1 2 75272 22667
0 22669 5 1 1 22668
0 22670 7 1 2 22585 22669
0 22671 5 1 1 22670
0 22672 7 1 2 51584 22671
0 22673 5 1 1 22672
0 22674 7 1 2 22515 22673
0 22675 5 1 1 22674
0 22676 7 1 2 51322 22675
0 22677 5 1 1 22676
0 22678 7 1 2 21140 9290
0 22679 5 1 1 22678
0 22680 7 1 2 52141 22679
0 22681 5 1 1 22680
0 22682 7 1 2 60723 71150
0 22683 5 1 1 22682
0 22684 7 1 2 22681 22683
0 22685 5 1 1 22684
0 22686 7 1 2 51928 22685
0 22687 5 1 1 22686
0 22688 7 2 2 48179 62156
0 22689 5 3 1 75393
0 22690 7 3 2 52961 65221
0 22691 5 1 1 75398
0 22692 7 1 2 65944 71168
0 22693 5 1 1 22692
0 22694 7 1 2 52285 22693
0 22695 5 1 1 22694
0 22696 7 1 2 22691 22695
0 22697 5 1 1 22696
0 22698 7 1 2 75395 22697
0 22699 5 1 1 22698
0 22700 7 1 2 63138 22476
0 22701 5 1 1 22700
0 22702 7 1 2 71151 22701
0 22703 5 1 1 22702
0 22704 7 1 2 22699 22703
0 22705 7 1 2 22687 22704
0 22706 5 1 1 22705
0 22707 7 2 2 53285 75273
0 22708 5 1 1 75401
0 22709 7 1 2 52490 75402
0 22710 5 2 1 22709
0 22711 7 1 2 49545 62478
0 22712 5 1 1 22711
0 22713 7 1 2 75403 22712
0 22714 5 5 1 22713
0 22715 7 1 2 22706 75405
0 22716 5 1 1 22715
0 22717 7 3 2 62149 75389
0 22718 5 5 1 75410
0 22719 7 1 2 61110 75411
0 22720 5 1 1 22719
0 22721 7 1 2 70588 72313
0 22722 7 1 2 22720 22721
0 22723 5 1 1 22722
0 22724 7 1 2 22716 22723
0 22725 5 1 1 22724
0 22726 7 1 2 51031 22725
0 22727 5 1 1 22726
0 22728 7 2 2 49546 60202
0 22729 5 1 1 75418
0 22730 7 1 2 55012 74872
0 22731 5 1 1 22730
0 22732 7 1 2 22729 22731
0 22733 5 1 1 22732
0 22734 7 1 2 51929 22733
0 22735 5 1 1 22734
0 22736 7 1 2 60625 64710
0 22737 5 1 1 22736
0 22738 7 1 2 22735 22737
0 22739 5 1 1 22738
0 22740 7 1 2 52491 22739
0 22741 5 1 1 22740
0 22742 7 1 2 53093 62609
0 22743 5 2 1 22742
0 22744 7 1 2 52286 60238
0 22745 7 1 2 70992 22744
0 22746 5 1 1 22745
0 22747 7 1 2 75420 22746
0 22748 5 1 1 22747
0 22749 7 1 2 73200 22748
0 22750 5 1 1 22749
0 22751 7 1 2 22741 22750
0 22752 5 1 1 22751
0 22753 7 1 2 50736 22752
0 22754 5 1 1 22753
0 22755 7 7 2 52492 55013
0 22756 5 1 1 75422
0 22757 7 2 2 54647 73417
0 22758 7 1 2 75423 75429
0 22759 5 1 1 22758
0 22760 7 1 2 22754 22759
0 22761 5 1 1 22760
0 22762 7 1 2 57228 22761
0 22763 5 1 1 22762
0 22764 7 15 2 53286 54648
0 22765 7 5 2 52493 75431
0 22766 5 2 1 75446
0 22767 7 1 2 54297 70825
0 22768 5 2 1 22767
0 22769 7 1 2 75447 75453
0 22770 5 1 1 22769
0 22771 7 1 2 51930 61298
0 22772 5 1 1 22771
0 22773 7 1 2 64473 22772
0 22774 5 1 1 22773
0 22775 7 1 2 56627 22774
0 22776 5 1 1 22775
0 22777 7 1 2 65236 22776
0 22778 5 2 1 22777
0 22779 7 1 2 50203 58022
0 22780 7 1 2 60570 22779
0 22781 7 1 2 75455 22780
0 22782 5 1 1 22781
0 22783 7 1 2 22770 22782
0 22784 5 1 1 22783
0 22785 7 1 2 55014 22784
0 22786 5 1 1 22785
0 22787 7 1 2 22763 22786
0 22788 5 1 1 22787
0 22789 7 1 2 58430 22788
0 22790 5 1 1 22789
0 22791 7 1 2 59380 21130
0 22792 5 1 1 22791
0 22793 7 1 2 61489 22792
0 22794 5 1 1 22793
0 22795 7 2 2 54298 55754
0 22796 5 3 1 75457
0 22797 7 1 2 60239 74179
0 22798 7 1 2 75459 22797
0 22799 5 1 1 22798
0 22800 7 1 2 75451 22799
0 22801 7 1 2 22794 22800
0 22802 5 1 1 22801
0 22803 7 1 2 55898 58023
0 22804 7 1 2 22802 22803
0 22805 5 1 1 22804
0 22806 7 1 2 58836 75145
0 22807 5 1 1 22806
0 22808 7 1 2 75143 22807
0 22809 5 1 1 22808
0 22810 7 2 2 58024 71152
0 22811 7 1 2 22809 75462
0 22812 5 1 1 22811
0 22813 7 1 2 60419 75448
0 22814 5 1 1 22813
0 22815 7 1 2 22812 22814
0 22816 5 1 1 22815
0 22817 7 1 2 57609 22816
0 22818 5 1 1 22817
0 22819 7 1 2 60364 65755
0 22820 5 1 1 22819
0 22821 7 1 2 56452 60571
0 22822 7 1 2 22820 22821
0 22823 5 1 1 22822
0 22824 7 1 2 22818 22823
0 22825 7 1 2 22805 22824
0 22826 5 1 1 22825
0 22827 7 1 2 55015 22826
0 22828 5 1 1 22827
0 22829 7 6 2 52494 50737
0 22830 7 1 2 75464 75419
0 22831 5 1 1 22830
0 22832 7 1 2 63764 66250
0 22833 5 2 1 22832
0 22834 7 1 2 75452 75470
0 22835 5 1 1 22834
0 22836 7 1 2 52142 73769
0 22837 7 1 2 22835 22836
0 22838 5 1 1 22837
0 22839 7 1 2 22831 22838
0 22840 5 1 1 22839
0 22841 7 1 2 75369 22840
0 22842 5 1 1 22841
0 22843 7 2 2 58891 73918
0 22844 5 1 1 75472
0 22845 7 1 2 59797 74880
0 22846 5 1 1 22845
0 22847 7 1 2 22844 22846
0 22848 5 1 1 22847
0 22849 7 1 2 75013 22848
0 22850 5 1 1 22849
0 22851 7 1 2 70205 75449
0 22852 5 1 1 22851
0 22853 7 1 2 22850 22852
0 22854 5 1 1 22853
0 22855 7 1 2 55016 22854
0 22856 5 1 1 22855
0 22857 7 1 2 75035 75225
0 22858 5 1 1 22857
0 22859 7 1 2 22856 22858
0 22860 5 1 1 22859
0 22861 7 1 2 59860 22860
0 22862 5 1 1 22861
0 22863 7 1 2 22842 22862
0 22864 7 1 2 22828 22863
0 22865 7 1 2 22790 22864
0 22866 5 1 1 22865
0 22867 7 1 2 62479 22866
0 22868 5 1 1 22867
0 22869 7 1 2 22727 22868
0 22870 5 1 1 22869
0 22871 7 2 2 65986 22870
0 22872 5 1 1 75474
0 22873 7 1 2 22677 22872
0 22874 5 1 1 22873
0 22875 7 1 2 57010 22874
0 22876 5 1 1 22875
0 22877 7 5 2 52495 48752
0 22878 5 1 1 75476
0 22879 7 1 2 63176 68304
0 22880 5 1 1 22879
0 22881 7 12 2 53287 49746
0 22882 5 1 1 75481
0 22883 7 4 2 50738 75482
0 22884 7 1 2 55899 75493
0 22885 5 1 1 22884
0 22886 7 1 2 22880 22885
0 22887 5 1 1 22886
0 22888 7 1 2 75477 22887
0 22889 5 1 1 22888
0 22890 7 9 2 52625 49547
0 22891 5 7 1 75497
0 22892 7 9 2 48605 53288
0 22893 5 5 1 75513
0 22894 7 2 2 50204 75514
0 22895 5 1 1 75527
0 22896 7 1 2 75506 22895
0 22897 5 2 1 22896
0 22898 7 1 2 56731 75529
0 22899 5 1 1 22898
0 22900 7 1 2 52626 63874
0 22901 5 1 1 22900
0 22902 7 1 2 22899 22901
0 22903 5 1 1 22902
0 22904 7 1 2 54299 22903
0 22905 5 1 1 22904
0 22906 7 1 2 67299 75498
0 22907 5 1 1 22906
0 22908 7 1 2 22905 22907
0 22909 5 1 1 22908
0 22910 7 1 2 56097 22909
0 22911 5 1 1 22910
0 22912 7 5 2 52627 54029
0 22913 5 1 1 75531
0 22914 7 1 2 57171 57295
0 22915 5 1 1 22914
0 22916 7 1 2 2890 22915
0 22917 5 1 1 22916
0 22918 7 1 2 75532 22917
0 22919 5 1 1 22918
0 22920 7 1 2 22911 22919
0 22921 5 1 1 22920
0 22922 7 1 2 47925 22921
0 22923 5 1 1 22922
0 22924 7 2 2 52628 56732
0 22925 7 1 2 64693 75536
0 22926 5 1 1 22925
0 22927 7 1 2 22923 22926
0 22928 5 1 1 22927
0 22929 7 1 2 55755 22928
0 22930 5 1 1 22929
0 22931 7 2 2 48180 63875
0 22932 5 1 1 75538
0 22933 7 1 2 49548 58286
0 22934 5 1 1 22933
0 22935 7 1 2 22932 22934
0 22936 5 1 1 22935
0 22937 7 1 2 52629 22936
0 22938 5 1 1 22937
0 22939 7 1 2 61093 75528
0 22940 5 1 1 22939
0 22941 7 1 2 22938 22940
0 22942 5 1 1 22941
0 22943 7 1 2 54300 22942
0 22944 5 1 1 22943
0 22945 7 1 2 52630 67386
0 22946 7 1 2 69005 22945
0 22947 5 1 1 22946
0 22948 7 1 2 22944 22947
0 22949 5 1 1 22948
0 22950 7 1 2 56098 22949
0 22951 5 1 1 22950
0 22952 7 1 2 64540 67444
0 22953 5 1 1 22952
0 22954 7 1 2 52496 22953
0 22955 5 1 1 22954
0 22956 7 1 2 49549 22955
0 22957 5 1 1 22956
0 22958 7 1 2 57296 74606
0 22959 5 1 1 22958
0 22960 7 1 2 22957 22959
0 22961 5 1 1 22960
0 22962 7 1 2 52631 22961
0 22963 5 1 1 22962
0 22964 7 1 2 22951 22963
0 22965 7 1 2 22930 22964
0 22966 5 1 1 22965
0 22967 7 1 2 54649 22966
0 22968 5 1 1 22967
0 22969 7 6 2 48606 52632
0 22970 7 4 2 49550 75540
0 22971 5 1 1 75546
0 22972 7 2 2 48607 73427
0 22973 5 1 1 75550
0 22974 7 1 2 22973 75507
0 22975 5 3 1 22974
0 22976 7 1 2 67453 75552
0 22977 5 1 1 22976
0 22978 7 1 2 22971 22977
0 22979 5 1 1 22978
0 22980 7 1 2 60240 22979
0 22981 5 1 1 22980
0 22982 7 1 2 55756 71988
0 22983 7 1 2 75553 22982
0 22984 5 1 1 22983
0 22985 7 1 2 22981 22984
0 22986 7 1 2 22968 22985
0 22987 5 1 1 22986
0 22988 7 1 2 56348 22987
0 22989 5 1 1 22988
0 22990 7 1 2 50739 59308
0 22991 5 1 1 22990
0 22992 7 1 2 49551 22991
0 22993 5 1 1 22992
0 22994 7 1 2 61000 66862
0 22995 5 1 1 22994
0 22996 7 1 2 22993 22995
0 22997 5 1 1 22996
0 22998 7 1 2 47926 22997
0 22999 5 1 1 22998
0 23000 7 3 2 54301 62403
0 23001 5 1 1 75555
0 23002 7 1 2 49552 75556
0 23003 5 1 1 23002
0 23004 7 1 2 22999 23003
0 23005 5 1 1 23004
0 23006 7 1 2 67207 23005
0 23007 5 1 1 23006
0 23008 7 1 2 64235 61001
0 23009 7 1 2 71788 23008
0 23010 5 1 1 23009
0 23011 7 1 2 23007 23010
0 23012 5 1 1 23011
0 23013 7 1 2 54030 23012
0 23014 5 1 1 23013
0 23015 7 2 2 56733 61081
0 23016 5 1 1 75558
0 23017 7 1 2 67236 75559
0 23018 5 1 1 23017
0 23019 7 1 2 23014 23018
0 23020 5 1 1 23019
0 23021 7 1 2 55757 23020
0 23022 5 1 1 23021
0 23023 7 1 2 49553 67445
0 23024 5 1 1 23023
0 23025 7 1 2 62856 74002
0 23026 5 1 1 23025
0 23027 7 1 2 23024 23026
0 23028 5 1 1 23027
0 23029 7 1 2 67208 23028
0 23030 5 1 1 23029
0 23031 7 1 2 58153 71855
0 23032 5 1 1 23031
0 23033 7 1 2 23030 23032
0 23034 5 1 1 23033
0 23035 7 1 2 48381 23034
0 23036 5 1 1 23035
0 23037 7 1 2 62297 65784
0 23038 5 1 1 23037
0 23039 7 1 2 67237 23038
0 23040 5 1 1 23039
0 23041 7 1 2 23036 23040
0 23042 5 1 1 23041
0 23043 7 1 2 48181 23042
0 23044 5 1 1 23043
0 23045 7 4 2 48608 49433
0 23046 5 1 1 75560
0 23047 7 2 2 63346 75561
0 23048 5 1 1 75564
0 23049 7 1 2 47927 59581
0 23050 5 3 1 23049
0 23051 7 2 2 59299 75566
0 23052 5 3 1 75569
0 23053 7 1 2 54031 75571
0 23054 5 1 1 23053
0 23055 7 1 2 64462 23054
0 23056 5 1 1 23055
0 23057 7 1 2 67238 23056
0 23058 5 1 1 23057
0 23059 7 1 2 23048 23058
0 23060 7 1 2 23044 23059
0 23061 5 1 1 23060
0 23062 7 1 2 54302 23061
0 23063 5 1 1 23062
0 23064 7 1 2 54650 67460
0 23065 5 2 1 23064
0 23066 7 1 2 61094 63223
0 23067 5 1 1 23066
0 23068 7 1 2 65899 23067
0 23069 7 1 2 75574 23068
0 23070 5 1 1 23069
0 23071 7 1 2 67239 23070
0 23072 5 1 1 23071
0 23073 7 1 2 23063 23072
0 23074 7 1 2 23022 23073
0 23075 5 1 1 23074
0 23076 7 1 2 52633 23075
0 23077 5 1 1 23076
0 23078 7 1 2 64002 75530
0 23079 5 1 1 23078
0 23080 7 2 2 54032 75554
0 23081 7 1 2 63966 75576
0 23082 5 1 1 23081
0 23083 7 1 2 23079 23082
0 23084 5 1 1 23083
0 23085 7 1 2 48182 23084
0 23086 5 1 1 23085
0 23087 7 2 2 54651 75533
0 23088 5 1 1 75578
0 23089 7 1 2 64043 75579
0 23090 5 1 1 23089
0 23091 7 1 2 23086 23090
0 23092 5 1 1 23091
0 23093 7 1 2 54303 23092
0 23094 5 1 1 23093
0 23095 7 5 2 54652 75499
0 23096 5 1 1 75580
0 23097 7 1 2 70199 75581
0 23098 5 1 1 23097
0 23099 7 1 2 23094 23098
0 23100 5 1 1 23099
0 23101 7 1 2 56349 23100
0 23102 5 1 1 23101
0 23103 7 2 2 67209 75500
0 23104 5 1 1 75585
0 23105 7 1 2 63152 75586
0 23106 5 1 1 23105
0 23107 7 2 2 64350 73428
0 23108 5 1 1 75587
0 23109 7 1 2 23108 23104
0 23110 5 2 1 23109
0 23111 7 3 2 56099 62325
0 23112 5 1 1 75591
0 23113 7 1 2 63117 23112
0 23114 5 1 1 23113
0 23115 7 1 2 75589 23114
0 23116 5 1 1 23115
0 23117 7 1 2 23106 23116
0 23118 7 1 2 23102 23117
0 23119 5 1 1 23118
0 23120 7 1 2 58606 23119
0 23121 5 1 1 23120
0 23122 7 1 2 48183 75572
0 23123 5 1 1 23122
0 23124 7 1 2 63149 23123
0 23125 5 1 1 23124
0 23126 7 1 2 54304 23125
0 23127 5 1 1 23126
0 23128 7 1 2 54305 75573
0 23129 5 1 1 23128
0 23130 7 1 2 66185 23129
0 23131 5 1 1 23130
0 23132 7 1 2 54033 23131
0 23133 5 2 1 23132
0 23134 7 2 2 64850 60760
0 23135 5 2 1 75596
0 23136 7 1 2 60420 75597
0 23137 5 3 1 23136
0 23138 7 1 2 56100 75600
0 23139 5 1 1 23138
0 23140 7 1 2 73947 23139
0 23141 5 1 1 23140
0 23142 7 1 2 55758 23141
0 23143 5 2 1 23142
0 23144 7 1 2 75594 75603
0 23145 7 1 2 23127 23144
0 23146 5 1 1 23145
0 23147 7 1 2 75588 23146
0 23148 5 1 1 23147
0 23149 7 1 2 23121 23148
0 23150 7 1 2 23077 23149
0 23151 7 1 2 22989 23150
0 23152 5 1 1 23151
0 23153 7 1 2 53500 23152
0 23154 5 1 1 23153
0 23155 7 1 2 22889 23154
0 23156 5 1 1 23155
0 23157 7 1 2 51032 23156
0 23158 5 1 1 23157
0 23159 7 1 2 56101 69393
0 23160 5 1 1 23159
0 23161 7 2 2 58398 61819
0 23162 5 1 1 75605
0 23163 7 1 2 62404 63940
0 23164 5 2 1 23163
0 23165 7 1 2 23162 75607
0 23166 5 1 1 23165
0 23167 7 1 2 57826 23166
0 23168 5 1 1 23167
0 23169 7 1 2 59193 7307
0 23170 5 2 1 23169
0 23171 7 1 2 60241 75609
0 23172 5 1 1 23171
0 23173 7 1 2 52497 23172
0 23174 7 1 2 23168 23173
0 23175 7 1 2 23160 23174
0 23176 7 2 2 75604 23175
0 23177 5 1 1 75611
0 23178 7 1 2 51033 23177
0 23179 5 1 1 23178
0 23180 7 1 2 22756 23179
0 23181 5 1 1 23180
0 23182 7 1 2 50740 23181
0 23183 5 1 1 23182
0 23184 7 1 2 52498 63557
0 23185 5 1 1 23184
0 23186 7 1 2 23183 23185
0 23187 5 1 1 23186
0 23188 7 1 2 53289 23187
0 23189 5 1 1 23188
0 23190 7 2 2 59141 75226
0 23191 5 1 1 75613
0 23192 7 1 2 56102 23191
0 23193 5 1 1 23192
0 23194 7 5 2 49554 59142
0 23195 5 1 1 75615
0 23196 7 1 2 75384 23195
0 23197 5 1 1 23196
0 23198 7 1 2 23193 23197
0 23199 5 1 1 23198
0 23200 7 1 2 23189 23199
0 23201 5 1 1 23200
0 23202 7 1 2 75274 23201
0 23203 5 1 1 23202
0 23204 7 1 2 63215 70333
0 23205 5 2 1 23204
0 23206 7 5 2 52388 54306
0 23207 5 4 1 75622
0 23208 7 1 2 51034 61772
0 23209 7 1 2 75623 23208
0 23210 7 1 2 75620 23209
0 23211 5 1 1 23210
0 23212 7 1 2 52389 62697
0 23213 7 1 2 23001 23212
0 23214 7 1 2 69484 23213
0 23215 7 1 2 55759 75601
0 23216 5 1 1 23215
0 23217 7 1 2 69398 23216
0 23218 7 1 2 23214 23217
0 23219 5 1 1 23218
0 23220 7 1 2 62480 64197
0 23221 7 1 2 23219 23220
0 23222 5 1 1 23221
0 23223 7 1 2 23211 23222
0 23224 5 1 1 23223
0 23225 7 1 2 54653 23224
0 23226 5 1 1 23225
0 23227 7 1 2 62481 64455
0 23228 5 1 1 23227
0 23229 7 3 2 52962 63201
0 23230 5 1 1 75631
0 23231 7 1 2 73520 75632
0 23232 5 1 1 23231
0 23233 7 1 2 67340 73208
0 23234 5 1 1 23233
0 23235 7 1 2 52499 18954
0 23236 7 1 2 23234 23235
0 23237 5 1 1 23236
0 23238 7 4 2 52634 52963
0 23239 5 1 1 75634
0 23240 7 1 2 73521 75635
0 23241 5 1 1 23240
0 23242 7 2 2 48753 71110
0 23243 5 4 1 75638
0 23244 7 1 2 23241 75640
0 23245 7 1 2 23237 23244
0 23246 5 1 1 23245
0 23247 7 1 2 49747 23246
0 23248 5 1 1 23247
0 23249 7 1 2 23232 23248
0 23250 5 1 1 23249
0 23251 7 1 2 55900 65468
0 23252 7 1 2 23250 23251
0 23253 5 1 1 23252
0 23254 7 1 2 23228 23253
0 23255 7 1 2 23226 23254
0 23256 5 1 1 23255
0 23257 7 1 2 53168 23256
0 23258 5 1 1 23257
0 23259 7 4 2 52500 64275
0 23260 5 2 1 75644
0 23261 7 1 2 62461 67197
0 23262 5 1 1 23261
0 23263 7 1 2 63941 23262
0 23264 5 1 1 23263
0 23265 7 1 2 61940 58588
0 23266 5 1 1 23265
0 23267 7 1 2 23264 23266
0 23268 5 2 1 23267
0 23269 7 1 2 57827 75650
0 23270 5 1 1 23269
0 23271 7 1 2 57802 67198
0 23272 5 5 1 23271
0 23273 7 1 2 69394 75652
0 23274 5 1 1 23273
0 23275 7 1 2 57311 23274
0 23276 7 1 2 23270 23275
0 23277 5 1 1 23276
0 23278 7 1 2 53290 23277
0 23279 5 1 1 23278
0 23280 7 1 2 75648 23279
0 23281 5 1 1 23280
0 23282 7 1 2 54654 23281
0 23283 5 1 1 23282
0 23284 7 4 2 56103 57099
0 23285 5 1 1 75657
0 23286 7 1 2 74560 75658
0 23287 5 1 1 23286
0 23288 7 2 2 50444 64098
0 23289 7 1 2 61995 75661
0 23290 5 1 1 23289
0 23291 7 1 2 57722 23290
0 23292 5 1 1 23291
0 23293 7 1 2 23287 23292
0 23294 5 1 1 23293
0 23295 7 1 2 47928 23294
0 23296 5 1 1 23295
0 23297 7 1 2 59512 66703
0 23298 5 1 1 23297
0 23299 7 1 2 64075 63876
0 23300 5 1 1 23299
0 23301 7 1 2 57362 23300
0 23302 7 1 2 23298 23301
0 23303 5 1 1 23302
0 23304 7 1 2 56734 23303
0 23305 5 1 1 23304
0 23306 7 1 2 64086 67300
0 23307 5 1 1 23306
0 23308 7 1 2 23305 23307
0 23309 5 1 1 23308
0 23310 7 1 2 56104 23309
0 23311 5 1 1 23310
0 23312 7 1 2 57723 20585
0 23313 5 1 1 23312
0 23314 7 1 2 65592 23313
0 23315 7 1 2 23311 23314
0 23316 7 1 2 23296 23315
0 23317 5 1 1 23316
0 23318 7 1 2 50741 23317
0 23319 5 2 1 23318
0 23320 7 1 2 71806 75432
0 23321 5 1 1 23320
0 23322 7 1 2 56551 74226
0 23323 5 1 1 23322
0 23324 7 1 2 23321 23323
0 23325 5 1 1 23324
0 23326 7 1 2 56350 23325
0 23327 5 1 1 23326
0 23328 7 2 2 67210 75433
0 23329 7 1 2 62405 75665
0 23330 5 1 1 23329
0 23331 7 1 2 23327 23330
0 23332 5 1 1 23331
0 23333 7 1 2 60242 23332
0 23334 5 1 1 23333
0 23335 7 1 2 50742 57724
0 23336 5 1 1 23335
0 23337 7 7 2 47929 53291
0 23338 5 1 1 75667
0 23339 7 3 2 54655 75653
0 23340 7 1 2 75668 75674
0 23341 5 1 1 23340
0 23342 7 1 2 23336 23341
0 23343 5 1 1 23342
0 23344 7 1 2 54034 23343
0 23345 5 1 1 23344
0 23346 7 10 2 53292 54307
0 23347 5 1 1 75677
0 23348 7 1 2 75678 75675
0 23349 5 1 1 23348
0 23350 7 1 2 23345 23349
0 23351 5 1 1 23350
0 23352 7 1 2 56735 23351
0 23353 5 1 1 23352
0 23354 7 2 2 48184 53293
0 23355 7 2 2 65911 75687
0 23356 5 1 1 75689
0 23357 7 2 2 54656 75690
0 23358 5 1 1 75691
0 23359 7 1 2 56105 75692
0 23360 5 1 1 23359
0 23361 7 5 2 50743 56552
0 23362 7 1 2 66773 75693
0 23363 5 1 1 23362
0 23364 7 3 2 49331 53294
0 23365 7 3 2 48382 75698
0 23366 7 1 2 62780 75701
0 23367 5 1 1 23366
0 23368 7 1 2 23363 23367
0 23369 7 1 2 23360 23368
0 23370 5 1 1 23369
0 23371 7 1 2 56351 23370
0 23372 5 1 1 23371
0 23373 7 2 2 61907 75679
0 23374 7 1 2 67211 75704
0 23375 5 1 1 23374
0 23376 7 2 2 23372 23375
0 23377 7 2 2 48383 71967
0 23378 5 2 1 75708
0 23379 7 1 2 57282 75709
0 23380 5 1 1 23379
0 23381 7 1 2 74227 74473
0 23382 5 1 1 23381
0 23383 7 1 2 23380 23382
0 23384 5 1 1 23383
0 23385 7 1 2 57100 23384
0 23386 5 1 1 23385
0 23387 7 1 2 75706 23386
0 23388 7 1 2 23353 23387
0 23389 5 1 1 23388
0 23390 7 1 2 55760 23389
0 23391 5 1 1 23390
0 23392 7 1 2 23334 23391
0 23393 7 1 2 75663 23392
0 23394 7 1 2 23283 23393
0 23395 5 1 1 23394
0 23396 7 1 2 74991 23395
0 23397 5 1 1 23396
0 23398 7 1 2 23258 23397
0 23399 7 1 2 23203 23398
0 23400 7 1 2 23158 23399
0 23401 5 1 1 23400
0 23402 7 1 2 51323 23401
0 23403 5 1 1 23402
0 23404 7 1 2 58399 60395
0 23405 5 2 1 23404
0 23406 7 2 2 57610 75712
0 23407 5 1 1 75714
0 23408 7 2 2 49212 64051
0 23409 5 1 1 75716
0 23410 7 1 2 48185 75717
0 23411 5 1 1 23410
0 23412 7 1 2 75715 23411
0 23413 5 1 1 23412
0 23414 7 1 2 50744 23413
0 23415 5 1 1 23414
0 23416 7 6 2 52501 54657
0 23417 5 1 1 75718
0 23418 7 1 2 63942 59374
0 23419 5 1 1 23418
0 23420 7 1 2 23417 23419
0 23421 5 1 1 23420
0 23422 7 1 2 56736 23421
0 23423 5 1 1 23422
0 23424 7 2 2 48502 52502
0 23425 5 1 1 75724
0 23426 7 3 2 47930 65311
0 23427 5 1 1 75726
0 23428 7 1 2 4317 75727
0 23429 5 1 1 23428
0 23430 7 1 2 23425 23429
0 23431 7 1 2 23423 23430
0 23432 7 1 2 23415 23431
0 23433 5 1 1 23432
0 23434 7 1 2 49434 23433
0 23435 5 1 1 23434
0 23436 7 3 2 49435 55761
0 23437 5 2 1 75729
0 23438 7 1 2 54035 74582
0 23439 5 1 1 23438
0 23440 7 1 2 52390 23439
0 23441 5 1 1 23440
0 23442 7 1 2 54308 23441
0 23443 5 1 1 23442
0 23444 7 1 2 75732 23443
0 23445 5 1 1 23444
0 23446 7 1 2 75719 23445
0 23447 5 1 1 23446
0 23448 7 2 2 59220 70860
0 23449 5 1 1 75734
0 23450 7 1 2 50745 75735
0 23451 5 1 1 23450
0 23452 7 3 2 52503 54036
0 23453 7 2 2 54658 60748
0 23454 5 1 1 75739
0 23455 7 1 2 75736 75740
0 23456 5 1 1 23455
0 23457 7 1 2 23451 23456
0 23458 5 1 1 23457
0 23459 7 1 2 62070 23458
0 23460 5 1 1 23459
0 23461 7 1 2 23447 23460
0 23462 7 1 2 23435 23461
0 23463 7 1 2 54309 74014
0 23464 5 3 1 23463
0 23465 7 1 2 59466 4492
0 23466 5 1 1 23465
0 23467 7 1 2 48186 23466
0 23468 5 1 1 23467
0 23469 7 1 2 75741 23468
0 23470 5 1 1 23469
0 23471 7 1 2 59181 23470
0 23472 5 1 1 23471
0 23473 7 1 2 71953 23472
0 23474 5 1 1 23473
0 23475 7 1 2 50746 23474
0 23476 5 1 1 23475
0 23477 7 1 2 65192 75720
0 23478 5 1 1 23477
0 23479 7 4 2 58646 3349
0 23480 7 1 2 56200 57790
0 23481 5 2 1 23480
0 23482 7 1 2 62727 75748
0 23483 5 1 1 23482
0 23484 7 1 2 75744 23483
0 23485 5 1 1 23484
0 23486 7 1 2 55762 23485
0 23487 5 1 1 23486
0 23488 7 1 2 54310 66226
0 23489 5 1 1 23488
0 23490 7 1 2 56352 20688
0 23491 5 1 1 23490
0 23492 7 1 2 23489 23491
0 23493 7 1 2 23487 23492
0 23494 5 1 1 23493
0 23495 7 1 2 50747 23494
0 23496 5 1 1 23495
0 23497 7 1 2 23478 23496
0 23498 5 1 1 23497
0 23499 7 1 2 56106 23498
0 23500 5 1 1 23499
0 23501 7 1 2 23476 23500
0 23502 7 1 2 23462 23501
0 23503 5 2 1 23502
0 23504 7 1 2 53295 75750
0 23505 5 1 1 23504
0 23506 7 2 2 75234 75522
0 23507 5 12 1 75752
0 23508 7 1 2 56201 75754
0 23509 5 3 1 23508
0 23510 7 1 2 55901 61280
0 23511 5 1 1 23510
0 23512 7 1 2 48187 23511
0 23513 5 1 1 23512
0 23514 7 1 2 59795 75567
0 23515 7 1 2 23513 23514
0 23516 5 3 1 23515
0 23517 7 6 2 53169 54311
0 23518 5 1 1 75772
0 23519 7 1 2 75773 75434
0 23520 7 2 2 75769 23519
0 23521 5 1 1 75778
0 23522 7 1 2 49555 71246
0 23523 5 1 1 23522
0 23524 7 1 2 23521 23523
0 23525 5 1 1 23524
0 23526 7 1 2 50205 23525
0 23527 5 1 1 23526
0 23528 7 1 2 75766 23527
0 23529 7 1 2 23505 23528
0 23530 5 1 1 23529
0 23531 7 1 2 51035 23530
0 23532 5 1 1 23531
0 23533 7 4 2 54659 56202
0 23534 5 1 1 75780
0 23535 7 1 2 52964 72907
0 23536 5 1 1 23535
0 23537 7 1 2 23534 23536
0 23538 5 1 1 23537
0 23539 7 1 2 75380 23538
0 23540 5 1 1 23539
0 23541 7 1 2 23532 23540
0 23542 5 1 1 23541
0 23543 7 1 2 53501 23542
0 23544 5 1 1 23543
0 23545 7 1 2 60592 70702
0 23546 5 1 1 23545
0 23547 7 1 2 23544 23546
0 23548 5 1 1 23547
0 23549 7 1 2 52635 23548
0 23550 5 1 1 23549
0 23551 7 1 2 63202 73882
0 23552 7 1 2 73297 23551
0 23553 7 1 2 71466 23552
0 23554 5 1 1 23553
0 23555 7 1 2 23550 23554
0 23556 5 1 1 23555
0 23557 7 1 2 55350 23556
0 23558 5 1 1 23557
0 23559 7 5 2 52391 49748
0 23560 7 1 2 73363 75784
0 23561 5 1 1 23560
0 23562 7 1 2 53502 75627
0 23563 5 1 1 23562
0 23564 7 1 2 58025 74414
0 23565 7 1 2 23563 23564
0 23566 5 1 1 23565
0 23567 7 1 2 23561 23566
0 23568 5 1 1 23567
0 23569 7 1 2 53170 23568
0 23570 5 1 1 23569
0 23571 7 1 2 64790 73830
0 23572 5 1 1 23571
0 23573 7 1 2 23570 23572
0 23574 5 1 1 23573
0 23575 7 1 2 55017 23574
0 23576 5 1 1 23575
0 23577 7 1 2 56553 14710
0 23578 5 1 1 23577
0 23579 7 4 2 58026 23578
0 23580 7 1 2 49749 75789
0 23581 5 2 1 23580
0 23582 7 1 2 72329 75793
0 23583 5 1 1 23582
0 23584 7 1 2 63595 23583
0 23585 5 1 1 23584
0 23586 7 1 2 49750 72439
0 23587 5 1 1 23586
0 23588 7 1 2 23585 23587
0 23589 5 1 1 23588
0 23590 7 1 2 75351 23589
0 23591 5 1 1 23590
0 23592 7 1 2 23576 23591
0 23593 5 1 1 23592
0 23594 7 1 2 50748 23593
0 23595 5 1 1 23594
0 23596 7 1 2 49436 72440
0 23597 5 2 1 23596
0 23598 7 1 2 73240 75795
0 23599 5 2 1 23598
0 23600 7 2 2 55018 75797
0 23601 5 1 1 75799
0 23602 7 4 2 53296 55351
0 23603 7 2 2 75352 75801
0 23604 7 1 2 64328 75805
0 23605 5 1 1 23604
0 23606 7 1 2 23601 23605
0 23607 5 1 1 23606
0 23608 7 1 2 54660 23607
0 23609 5 1 1 23608
0 23610 7 11 2 53094 71089
0 23611 5 1 1 75807
0 23612 7 2 2 48609 23611
0 23613 5 5 1 75818
0 23614 7 5 2 49556 68390
0 23615 7 1 2 60679 75825
0 23616 7 1 2 75820 23615
0 23617 5 1 1 23616
0 23618 7 1 2 53503 23617
0 23619 7 1 2 23609 23618
0 23620 5 1 1 23619
0 23621 7 5 2 52392 58027
0 23622 7 1 2 52504 75806
0 23623 5 1 1 23622
0 23624 7 1 2 63752 23623
0 23625 5 1 1 23624
0 23626 7 1 2 75830 23625
0 23627 5 1 1 23626
0 23628 7 1 2 75146 69505
0 23629 5 1 1 23628
0 23630 7 1 2 23627 23629
0 23631 5 1 1 23630
0 23632 7 1 2 55902 23631
0 23633 5 1 1 23632
0 23634 7 5 2 55019 56453
0 23635 7 1 2 51324 75835
0 23636 5 1 1 23635
0 23637 7 1 2 49751 23636
0 23638 7 1 2 23633 23637
0 23639 5 1 1 23638
0 23640 7 1 2 52965 23639
0 23641 7 1 2 23620 23640
0 23642 5 1 1 23641
0 23643 7 1 2 23595 23642
0 23644 5 1 1 23643
0 23645 7 1 2 52636 23644
0 23646 5 1 1 23645
0 23647 7 2 2 60472 66029
0 23648 5 1 1 75840
0 23649 7 1 2 62365 23648
0 23650 5 2 1 23649
0 23651 7 1 2 58028 75842
0 23652 5 1 1 23651
0 23653 7 2 2 73228 73278
0 23654 5 1 1 75844
0 23655 7 1 2 23652 75845
0 23656 5 2 1 23655
0 23657 7 1 2 63203 75846
0 23658 5 1 1 23657
0 23659 7 4 2 55903 70148
0 23660 5 1 1 75848
0 23661 7 4 2 53171 49752
0 23662 7 3 2 73429 75852
0 23663 5 2 1 75856
0 23664 7 1 2 75849 75857
0 23665 5 2 1 23664
0 23666 7 1 2 23658 75861
0 23667 5 1 1 23666
0 23668 7 1 2 63732 23667
0 23669 5 1 1 23668
0 23670 7 1 2 50749 75257
0 23671 7 1 2 75100 23670
0 23672 5 1 1 23671
0 23673 7 4 2 58686 60486
0 23674 7 1 2 49753 66168
0 23675 7 1 2 75863 23674
0 23676 5 1 1 23675
0 23677 7 1 2 23672 23676
0 23678 5 1 1 23677
0 23679 7 1 2 53172 23678
0 23680 5 1 1 23679
0 23681 7 1 2 55352 71291
0 23682 7 1 2 75633 23681
0 23683 5 1 1 23682
0 23684 7 1 2 23680 23683
0 23685 5 1 1 23684
0 23686 7 1 2 52393 23685
0 23687 5 1 1 23686
0 23688 7 3 2 60520 63204
0 23689 7 1 2 63782 75867
0 23690 5 1 1 23689
0 23691 7 2 2 62570 61216
0 23692 7 1 2 75864 75870
0 23693 5 1 1 23692
0 23694 7 4 2 52505 75483
0 23695 5 2 1 75872
0 23696 7 1 2 72330 75876
0 23697 5 5 1 23696
0 23698 7 1 2 75878 75312
0 23699 5 1 1 23698
0 23700 7 1 2 23693 23699
0 23701 5 1 1 23700
0 23702 7 1 2 51325 23701
0 23703 5 1 1 23702
0 23704 7 1 2 23690 23703
0 23705 7 1 2 23687 23704
0 23706 5 1 1 23705
0 23707 7 1 2 75353 23706
0 23708 5 1 1 23707
0 23709 7 1 2 23669 23708
0 23710 7 1 2 23646 23709
0 23711 5 1 1 23710
0 23712 7 1 2 52886 23711
0 23713 5 1 1 23712
0 23714 7 2 2 50097 55020
0 23715 7 4 2 51326 75275
0 23716 7 1 2 75885 75843
0 23717 5 1 1 23716
0 23718 7 2 2 60572 72684
0 23719 7 2 2 55353 75889
0 23720 7 2 2 62482 56203
0 23721 7 1 2 75891 75893
0 23722 5 1 1 23721
0 23723 7 1 2 23717 23722
0 23724 5 1 1 23723
0 23725 7 1 2 58029 23724
0 23726 5 1 1 23725
0 23727 7 15 2 56454 62483
0 23728 5 3 1 75895
0 23729 7 1 2 75892 75896
0 23730 5 1 1 23729
0 23731 7 1 2 75276 23654
0 23732 5 1 1 23731
0 23733 7 3 2 52966 49437
0 23734 7 1 2 62484 64236
0 23735 7 1 2 75913 23734
0 23736 5 2 1 23735
0 23737 7 1 2 75916 75862
0 23738 7 1 2 23732 23737
0 23739 5 1 1 23738
0 23740 7 1 2 51327 23739
0 23741 5 1 1 23740
0 23742 7 1 2 23730 23741
0 23743 7 1 2 23726 23742
0 23744 5 1 1 23743
0 23745 7 1 2 75883 23744
0 23746 5 1 1 23745
0 23747 7 1 2 23713 23746
0 23748 5 1 1 23747
0 23749 7 1 2 51931 23748
0 23750 5 1 1 23749
0 23751 7 3 2 67756 75331
0 23752 7 1 2 48754 70111
0 23753 5 4 1 23752
0 23754 7 3 2 49754 75921
0 23755 5 1 1 75925
0 23756 7 2 2 63216 23755
0 23757 5 3 1 75928
0 23758 7 2 2 53297 75930
0 23759 5 1 1 75933
0 23760 7 1 2 75918 75934
0 23761 5 1 1 23760
0 23762 7 1 2 52967 75821
0 23763 5 1 1 23762
0 23764 7 1 2 62366 23763
0 23765 5 2 1 23764
0 23766 7 1 2 75277 75935
0 23767 5 1 1 23766
0 23768 7 9 2 52506 53173
0 23769 5 4 1 75937
0 23770 7 2 2 75938 75785
0 23771 5 3 1 75950
0 23772 7 1 2 72767 75951
0 23773 5 1 1 23772
0 23774 7 1 2 23767 23773
0 23775 5 1 1 23774
0 23776 7 1 2 53298 23775
0 23777 5 1 1 23776
0 23778 7 2 2 52507 62356
0 23779 5 2 1 75955
0 23780 7 1 2 62367 22507
0 23781 5 10 1 23780
0 23782 7 1 2 75808 75959
0 23783 5 1 1 23782
0 23784 7 1 2 75957 23783
0 23785 5 4 1 23784
0 23786 7 2 2 75278 75969
0 23787 5 1 1 75973
0 23788 7 1 2 23787 75917
0 23789 7 1 2 23777 23788
0 23790 5 1 1 23789
0 23791 7 1 2 63805 23790
0 23792 5 1 1 23791
0 23793 7 1 2 23761 23792
0 23794 5 1 1 23793
0 23795 7 1 2 51328 23794
0 23796 5 1 1 23795
0 23797 7 1 2 75919 75886
0 23798 5 2 1 23797
0 23799 7 2 2 52887 71222
0 23800 7 3 2 50098 63453
0 23801 7 1 2 75977 75979
0 23802 5 1 1 23801
0 23803 7 1 2 67341 23802
0 23804 5 1 1 23803
0 23805 7 1 2 55904 23804
0 23806 5 1 1 23805
0 23807 7 3 2 50750 64150
0 23808 7 2 2 59861 75982
0 23809 7 1 2 53299 75985
0 23810 5 1 1 23809
0 23811 7 1 2 23806 23810
0 23812 5 1 1 23811
0 23813 7 1 2 73837 23812
0 23814 5 1 1 23813
0 23815 7 1 2 75975 23814
0 23816 5 1 1 23815
0 23817 7 1 2 57312 23816
0 23818 5 1 1 23817
0 23819 7 3 2 52637 73818
0 23820 7 1 2 66898 75987
0 23821 5 1 1 23820
0 23822 7 3 2 53300 62678
0 23823 5 2 1 75990
0 23824 7 3 2 52888 73439
0 23825 7 1 2 75980 75995
0 23826 5 1 1 23825
0 23827 7 1 2 75993 23826
0 23828 5 1 1 23827
0 23829 7 1 2 55905 23828
0 23830 5 1 1 23829
0 23831 7 1 2 53504 75986
0 23832 5 1 1 23831
0 23833 7 1 2 23830 23832
0 23834 5 1 1 23833
0 23835 7 1 2 52638 23834
0 23836 5 1 1 23835
0 23837 7 5 2 48755 73819
0 23838 5 8 1 75998
0 23839 7 1 2 70811 75999
0 23840 5 1 1 23839
0 23841 7 1 2 23836 23840
0 23842 5 1 1 23841
0 23843 7 1 2 70149 23842
0 23844 5 1 1 23843
0 23845 7 1 2 23821 23844
0 23846 5 1 1 23845
0 23847 7 1 2 63596 23846
0 23848 5 1 1 23847
0 23849 7 1 2 23818 23848
0 23850 7 1 2 23796 23849
0 23851 7 1 2 23750 23850
0 23852 5 1 1 23851
0 23853 7 1 2 52143 23852
0 23854 5 1 1 23853
0 23855 7 1 2 51036 73134
0 23856 5 1 1 23855
0 23857 7 1 2 73141 23856
0 23858 5 3 1 23857
0 23859 7 1 2 55906 76011
0 23860 5 1 1 23859
0 23861 7 3 2 63509 67557
0 23862 5 1 1 76014
0 23863 7 1 2 23860 23862
0 23864 5 1 1 23863
0 23865 7 1 2 75279 23864
0 23866 5 1 1 23865
0 23867 7 1 2 66899 73838
0 23868 5 1 1 23867
0 23869 7 1 2 70150 68584
0 23870 7 1 2 75920 23869
0 23871 5 1 1 23870
0 23872 7 1 2 23868 23871
0 23873 5 1 1 23872
0 23874 7 1 2 53174 23873
0 23875 5 1 1 23874
0 23876 7 1 2 23866 23875
0 23877 5 1 1 23876
0 23878 7 1 2 53301 23877
0 23879 5 1 1 23878
0 23880 7 2 2 55907 67327
0 23881 5 2 1 76017
0 23882 7 1 2 71223 75983
0 23883 5 1 1 23882
0 23884 7 1 2 76019 23883
0 23885 5 1 1 23884
0 23886 7 1 2 73839 23885
0 23887 5 1 1 23886
0 23888 7 1 2 75976 23887
0 23889 5 1 1 23888
0 23890 7 1 2 57313 23889
0 23891 5 1 1 23890
0 23892 7 3 2 52639 70151
0 23893 7 1 2 73440 75774
0 23894 7 1 2 63852 23893
0 23895 7 1 2 76021 23894
0 23896 5 1 1 23895
0 23897 7 2 2 23891 23896
0 23898 7 1 2 23879 76024
0 23899 5 1 1 23898
0 23900 7 1 2 62166 23899
0 23901 5 1 1 23900
0 23902 7 1 2 56204 64018
0 23903 5 2 1 23902
0 23904 7 1 2 72774 76026
0 23905 5 1 1 23904
0 23906 7 1 2 55021 23905
0 23907 5 1 1 23906
0 23908 7 1 2 52968 63558
0 23909 5 1 1 23908
0 23910 7 1 2 23907 23909
0 23911 5 1 1 23910
0 23912 7 1 2 75280 23911
0 23913 5 1 1 23912
0 23914 7 1 2 63559 75129
0 23915 5 1 1 23914
0 23916 7 1 2 23913 23915
0 23917 5 1 1 23916
0 23918 7 1 2 51329 23917
0 23919 5 1 1 23918
0 23920 7 3 2 62485 63831
0 23921 5 2 1 76028
0 23922 7 2 2 52969 63177
0 23923 5 2 1 76033
0 23924 7 1 2 72986 76034
0 23925 7 1 2 76029 23924
0 23926 5 1 1 23925
0 23927 7 1 2 23919 23926
0 23928 5 1 1 23927
0 23929 7 1 2 58030 23928
0 23930 5 1 1 23929
0 23931 7 1 2 23901 23930
0 23932 7 1 2 23854 23931
0 23933 7 1 2 23558 23932
0 23934 7 1 2 23403 23933
0 23935 5 1 1 23934
0 23936 7 1 2 51585 23935
0 23937 5 1 1 23936
0 23938 7 2 2 55022 57314
0 23939 7 1 2 72679 76037
0 23940 5 1 1 23939
0 23941 7 1 2 56107 61290
0 23942 5 1 1 23941
0 23943 7 1 2 58524 61257
0 23944 5 1 1 23943
0 23945 7 1 2 59182 23944
0 23946 5 1 1 23945
0 23947 7 1 2 23942 23946
0 23948 5 2 1 23947
0 23949 7 2 2 53175 76039
0 23950 5 1 1 76041
0 23951 7 1 2 51037 76042
0 23952 5 1 1 23951
0 23953 7 1 2 23940 23952
0 23954 5 2 1 23953
0 23955 7 1 2 75106 76043
0 23956 5 1 1 23955
0 23957 7 1 2 60049 65785
0 23958 5 1 1 23957
0 23959 7 1 2 48188 23958
0 23960 5 1 1 23959
0 23961 7 1 2 49332 61284
0 23962 5 1 1 23961
0 23963 7 1 2 23960 23962
0 23964 5 1 1 23963
0 23965 7 1 2 48384 23964
0 23966 5 1 1 23965
0 23967 7 1 2 58480 62266
0 23968 5 1 1 23967
0 23969 7 1 2 23966 23968
0 23970 5 1 1 23969
0 23971 7 1 2 56353 23970
0 23972 5 1 1 23971
0 23973 7 2 2 61608 61975
0 23974 5 1 1 76045
0 23975 7 4 2 61197 23974
0 23976 5 6 1 76047
0 23977 7 1 2 55908 76048
0 23978 5 2 1 23977
0 23979 7 1 2 56921 76057
0 23980 5 1 1 23979
0 23981 7 1 2 23972 23980
0 23982 5 1 1 23981
0 23983 7 1 2 51330 66900
0 23984 7 1 2 23982 23983
0 23985 5 1 1 23984
0 23986 7 1 2 23956 23985
0 23987 5 1 1 23986
0 23988 7 1 2 54661 23987
0 23989 5 1 1 23988
0 23990 7 3 2 48610 56205
0 23991 5 2 1 76059
0 23992 7 2 2 61969 62079
0 23993 5 3 1 76064
0 23994 7 1 2 73247 76065
0 23995 5 1 1 23994
0 23996 7 2 2 52508 23995
0 23997 5 1 1 76069
0 23998 7 1 2 55023 76070
0 23999 5 1 1 23998
0 24000 7 1 2 76062 23999
0 24001 5 1 1 24000
0 24002 7 1 2 50751 24001
0 24003 5 1 1 24002
0 24004 7 3 2 52394 51038
0 24005 7 1 2 48611 76071
0 24006 5 1 1 24005
0 24007 7 2 2 24003 24006
0 24008 5 1 1 76074
0 24009 7 1 2 75107 24008
0 24010 5 1 1 24009
0 24011 7 1 2 23989 24010
0 24012 5 1 1 24011
0 24013 7 1 2 53505 24012
0 24014 5 1 1 24013
0 24015 7 1 2 59788 75568
0 24016 5 1 1 24015
0 24017 7 1 2 48189 24016
0 24018 5 1 1 24017
0 24019 7 3 2 75320 24018
0 24020 5 1 1 76076
0 24021 7 1 2 52395 76077
0 24022 5 1 1 24021
0 24023 7 1 2 62486 63510
0 24024 7 1 2 24022 24023
0 24025 5 1 1 24024
0 24026 7 4 2 52509 52889
0 24027 5 1 1 76079
0 24028 7 1 2 75016 76080
0 24029 7 3 2 55024 72751
0 24030 7 1 2 76083 75841
0 24031 7 1 2 24028 24030
0 24032 5 1 1 24031
0 24033 7 1 2 24025 24032
0 24034 5 1 1 24033
0 24035 7 1 2 53176 24034
0 24036 5 1 1 24035
0 24037 7 2 2 49438 63511
0 24038 5 2 1 76086
0 24039 7 2 2 53095 68927
0 24040 7 1 2 60473 76090
0 24041 5 1 1 24040
0 24042 7 1 2 76088 24041
0 24043 5 1 1 24042
0 24044 7 1 2 62106 24043
0 24045 5 2 1 24044
0 24046 7 1 2 55909 76087
0 24047 5 1 1 24046
0 24048 7 1 2 76092 24047
0 24049 5 1 1 24048
0 24050 7 1 2 62487 24049
0 24051 5 1 1 24050
0 24052 7 1 2 24036 24051
0 24053 5 1 1 24052
0 24054 7 1 2 55354 24053
0 24055 5 1 1 24054
0 24056 7 1 2 62466 75541
0 24057 5 1 1 24056
0 24058 7 1 2 75268 24057
0 24059 5 1 1 24058
0 24060 7 1 2 69876 24059
0 24061 5 1 1 24060
0 24062 7 1 2 58941 75542
0 24063 5 1 1 24062
0 24064 7 1 2 75269 24063
0 24065 5 1 1 24064
0 24066 7 1 2 56737 24065
0 24067 5 1 1 24066
0 24068 7 1 2 24061 24067
0 24069 5 1 1 24068
0 24070 7 1 2 69506 24069
0 24071 5 1 1 24070
0 24072 7 1 2 24055 24071
0 24073 5 1 1 24072
0 24074 7 1 2 54037 24073
0 24075 5 1 1 24074
0 24076 7 1 2 66043 76049
0 24077 5 1 1 24076
0 24078 7 1 2 63512 24077
0 24079 5 1 1 24078
0 24080 7 7 2 52970 55025
0 24081 7 1 2 75809 76094
0 24082 5 1 1 24081
0 24083 7 1 2 55026 75960
0 24084 5 2 1 24083
0 24085 7 1 2 66904 76101
0 24086 7 1 2 24082 24085
0 24087 7 1 2 24079 24086
0 24088 5 1 1 24087
0 24089 7 1 2 51331 24088
0 24090 5 1 1 24089
0 24091 7 1 2 68391 75939
0 24092 7 1 2 71571 24091
0 24093 5 1 1 24092
0 24094 7 1 2 24090 24093
0 24095 5 1 1 24094
0 24096 7 1 2 75281 24095
0 24097 5 1 1 24096
0 24098 7 2 2 71186 68585
0 24099 7 1 2 63470 75339
0 24100 7 1 2 64522 24099
0 24101 7 1 2 76103 24100
0 24102 5 2 1 24101
0 24103 7 1 2 24097 76105
0 24104 7 1 2 24075 24103
0 24105 7 1 2 24014 24104
0 24106 5 1 1 24105
0 24107 7 1 2 53302 24106
0 24108 5 1 1 24107
0 24109 7 3 2 64276 71383
0 24110 5 1 1 76107
0 24111 7 1 2 52971 76108
0 24112 5 1 1 24111
0 24113 7 2 2 73135 72685
0 24114 7 1 2 63542 73433
0 24115 7 1 2 76110 24114
0 24116 5 1 1 24115
0 24117 7 1 2 24112 24116
0 24118 5 1 1 24117
0 24119 7 1 2 53506 24118
0 24120 5 1 1 24119
0 24121 7 4 2 51932 54038
0 24122 5 1 1 76112
0 24123 7 1 2 70272 76113
0 24124 7 1 2 76084 24123
0 24125 5 2 1 24124
0 24126 7 1 2 67342 76116
0 24127 5 1 1 24126
0 24128 7 1 2 73145 24127
0 24129 5 1 1 24128
0 24130 7 1 2 49557 72170
0 24131 5 1 1 24130
0 24132 7 1 2 24129 24131
0 24133 5 1 1 24132
0 24134 7 1 2 57315 24133
0 24135 5 1 1 24134
0 24136 7 1 2 24120 24135
0 24137 5 1 1 24136
0 24138 7 1 2 52640 24137
0 24139 5 1 1 24138
0 24140 7 1 2 63733 75974
0 24141 5 1 1 24140
0 24142 7 1 2 57316 66607
0 24143 7 1 2 67972 24142
0 24144 5 1 1 24143
0 24145 7 1 2 24141 24144
0 24146 7 2 2 24139 24145
0 24147 5 1 1 76118
0 24148 7 1 2 24108 76119
0 24149 5 1 1 24148
0 24150 7 1 2 51586 24149
0 24151 5 1 1 24150
0 24152 7 3 2 73674 69871
0 24153 5 1 1 76120
0 24154 7 1 2 75248 24153
0 24155 5 1 1 24154
0 24156 7 2 2 66509 24155
0 24157 7 1 2 75961 76123
0 24158 5 1 1 24157
0 24159 7 2 2 75940 75616
0 24160 5 1 1 76125
0 24161 7 1 2 23239 75958
0 24162 5 1 1 24161
0 24163 7 1 2 62082 73201
0 24164 7 1 2 24162 24163
0 24165 5 1 1 24164
0 24166 7 1 2 24160 24165
0 24167 7 1 2 24158 24166
0 24168 5 1 1 24167
0 24169 7 1 2 49755 24168
0 24170 5 1 1 24169
0 24171 7 1 2 52972 58031
0 24172 5 2 1 24171
0 24173 7 1 2 62368 76127
0 24174 5 2 1 24173
0 24175 7 1 2 66508 74972
0 24176 7 1 2 62167 24175
0 24177 7 1 2 76129 24176
0 24178 5 1 1 24177
0 24179 7 1 2 24170 24178
0 24180 5 1 1 24179
0 24181 7 1 2 51332 24180
0 24182 5 1 1 24181
0 24183 7 2 2 53909 58863
0 24184 5 1 1 76131
0 24185 7 3 2 7260 24184
0 24186 5 1 1 76133
0 24187 7 5 2 56738 24186
0 24188 5 1 1 76136
0 24189 7 3 2 52641 68928
0 24190 5 1 1 76141
0 24191 7 1 2 62770 75802
0 24192 7 1 2 76142 24191
0 24193 7 1 2 24188 24192
0 24194 5 1 1 24193
0 24195 7 1 2 24182 24194
0 24196 5 1 1 24195
0 24197 7 1 2 51587 24196
0 24198 5 1 1 24197
0 24199 7 3 2 53303 59023
0 24200 7 2 2 66216 76144
0 24201 7 4 2 53177 70589
0 24202 7 1 2 76147 76149
0 24203 5 1 1 24202
0 24204 7 1 2 24198 24203
0 24205 5 1 1 24204
0 24206 7 1 2 58525 24205
0 24207 5 1 1 24206
0 24208 7 2 2 49558 59221
0 24209 5 1 1 76153
0 24210 7 1 2 65128 24209
0 24211 5 1 1 24210
0 24212 7 1 2 59143 24211
0 24213 5 1 1 24212
0 24214 7 1 2 64517 63578
0 24215 5 1 1 24214
0 24216 7 1 2 24213 24215
0 24217 5 1 1 24216
0 24218 7 1 2 48612 24217
0 24219 5 1 1 24218
0 24220 7 1 2 65121 75617
0 24221 5 1 1 24220
0 24222 7 3 2 52642 63454
0 24223 7 1 2 56108 67253
0 24224 7 1 2 76155 24223
0 24225 5 1 1 24224
0 24226 7 1 2 24221 24225
0 24227 7 1 2 24219 24226
0 24228 5 1 1 24227
0 24229 7 1 2 56739 24228
0 24230 5 1 1 24229
0 24231 7 2 2 50752 67254
0 24232 5 1 1 76158
0 24233 7 1 2 66901 76159
0 24234 5 1 1 24233
0 24235 7 1 2 62655 67328
0 24236 5 1 1 24235
0 24237 7 1 2 24234 24236
0 24238 5 1 1 24237
0 24239 7 1 2 59108 24238
0 24240 5 1 1 24239
0 24241 7 6 2 48613 50753
0 24242 5 2 1 76160
0 24243 7 2 2 67329 76161
0 24244 5 3 1 76168
0 24245 7 2 2 52643 66828
0 24246 7 1 2 63953 76173
0 24247 5 1 1 24246
0 24248 7 1 2 76170 24247
0 24249 5 1 1 24248
0 24250 7 1 2 56354 24249
0 24251 5 1 1 24250
0 24252 7 3 2 62406 57101
0 24253 5 1 1 76175
0 24254 7 1 2 76156 76176
0 24255 5 1 1 24254
0 24256 7 1 2 24251 24255
0 24257 7 1 2 24240 24256
0 24258 5 1 1 24257
0 24259 7 1 2 69877 24258
0 24260 5 1 1 24259
0 24261 7 2 2 56355 70934
0 24262 5 1 1 76178
0 24263 7 1 2 76179 76169
0 24264 5 1 1 24263
0 24265 7 1 2 62010 76157
0 24266 5 1 1 24265
0 24267 7 1 2 76171 24266
0 24268 5 1 1 24267
0 24269 7 1 2 48503 24268
0 24270 5 1 1 24269
0 24271 7 4 2 51039 57939
0 24272 5 1 1 76180
0 24273 7 1 2 62648 76181
0 24274 5 1 1 24273
0 24275 7 1 2 56554 76174
0 24276 5 1 1 24275
0 24277 7 1 2 24274 24276
0 24278 7 1 2 24270 24277
0 24279 5 1 1 24278
0 24280 7 1 2 48385 24279
0 24281 5 1 1 24280
0 24282 7 1 2 24264 24281
0 24283 7 1 2 24260 24282
0 24284 7 1 2 24230 24283
0 24285 5 1 1 24284
0 24286 7 1 2 53507 24285
0 24287 5 1 1 24286
0 24288 7 1 2 69878 75610
0 24289 5 1 1 24288
0 24290 7 2 2 70391 75745
0 24291 5 2 1 76184
0 24292 7 1 2 67395 76185
0 24293 7 1 2 24289 24292
0 24294 5 1 1 24293
0 24295 7 1 2 50754 24294
0 24296 5 1 1 24295
0 24297 7 1 2 49559 60487
0 24298 5 1 1 24297
0 24299 7 1 2 24296 24298
0 24300 5 1 1 24299
0 24301 7 1 2 51040 24300
0 24302 5 1 1 24301
0 24303 7 2 2 57363 73770
0 24304 5 1 1 76188
0 24305 7 1 2 24302 24304
0 24306 5 1 1 24305
0 24307 7 1 2 75282 24306
0 24308 5 1 1 24307
0 24309 7 1 2 51333 24308
0 24310 7 1 2 24287 24309
0 24311 5 1 1 24310
0 24312 7 1 2 56206 75879
0 24313 5 2 1 24312
0 24314 7 1 2 53508 75227
0 24315 5 1 1 24314
0 24316 7 1 2 76190 24315
0 24317 5 1 1 24316
0 24318 7 1 2 52644 24317
0 24319 5 1 1 24318
0 24320 7 1 2 70105 76000
0 24321 5 2 1 24320
0 24322 7 1 2 24319 76192
0 24323 5 2 1 24322
0 24324 7 1 2 55910 76194
0 24325 5 1 1 24324
0 24326 7 4 2 53178 73820
0 24327 7 1 2 75543 76196
0 24328 5 1 1 24327
0 24329 7 1 2 24325 24328
0 24330 5 1 1 24329
0 24331 7 1 2 71494 24330
0 24332 5 1 1 24331
0 24333 7 2 2 74973 76095
0 24334 5 1 1 76200
0 24335 7 1 2 63579 76201
0 24336 7 1 2 70132 24335
0 24337 5 1 1 24336
0 24338 7 1 2 24332 24337
0 24339 5 1 1 24338
0 24340 7 1 2 62168 24339
0 24341 5 1 1 24340
0 24342 7 1 2 49756 75970
0 24343 5 1 1 24342
0 24344 7 6 2 48614 53509
0 24345 7 3 2 62150 70209
0 24346 5 1 1 76208
0 24347 7 1 2 76202 24346
0 24348 5 1 1 24347
0 24349 7 1 2 24343 24348
0 24350 5 1 1 24349
0 24351 7 1 2 53304 24350
0 24352 5 1 1 24351
0 24353 7 1 2 72314 75962
0 24354 5 1 1 24353
0 24355 7 1 2 58802 75941
0 24356 5 1 1 24355
0 24357 7 6 2 52973 49560
0 24358 7 1 2 53510 76211
0 24359 5 1 1 24358
0 24360 7 1 2 24356 24359
0 24361 5 1 1 24360
0 24362 7 1 2 75810 24361
0 24363 5 1 1 24362
0 24364 7 1 2 24354 24363
0 24365 7 1 2 24352 24364
0 24366 5 1 1 24365
0 24367 7 1 2 52645 24366
0 24368 5 1 1 24367
0 24369 7 3 2 73430 75942
0 24370 5 2 1 76217
0 24371 7 1 2 53305 71572
0 24372 7 1 2 75963 24371
0 24373 5 1 1 24372
0 24374 7 1 2 76220 24373
0 24375 5 1 1 24374
0 24376 7 1 2 48756 24375
0 24377 5 1 1 24376
0 24378 7 8 2 53179 49561
0 24379 5 1 1 76222
0 24380 7 1 2 76223 75465
0 24381 7 1 2 71573 24380
0 24382 5 1 1 24381
0 24383 7 1 2 24377 24382
0 24384 5 1 1 24383
0 24385 7 1 2 53511 24384
0 24386 5 1 1 24385
0 24387 7 1 2 24368 24386
0 24388 5 1 1 24387
0 24389 7 1 2 51041 24388
0 24390 5 1 1 24389
0 24391 7 1 2 63455 71187
0 24392 5 2 1 24391
0 24393 7 1 2 73434 71118
0 24394 7 1 2 57317 24393
0 24395 7 1 2 71241 24394
0 24396 5 1 1 24395
0 24397 7 1 2 76230 24396
0 24398 5 1 1 24397
0 24399 7 1 2 53512 24398
0 24400 5 1 1 24399
0 24401 7 1 2 73422 75858
0 24402 5 1 1 24401
0 24403 7 1 2 24400 24402
0 24404 5 1 1 24403
0 24405 7 1 2 52646 24404
0 24406 5 1 1 24405
0 24407 7 2 2 56207 56628
0 24408 7 1 2 75478 76145
0 24409 7 1 2 76232 24408
0 24410 5 1 1 24409
0 24411 7 1 2 24406 24410
0 24412 5 1 1 24411
0 24413 7 1 2 55911 24412
0 24414 5 1 1 24413
0 24415 7 1 2 59024 71255
0 24416 7 5 2 52974 53180
0 24417 5 1 1 76234
0 24418 7 1 2 76235 75544
0 24419 7 1 2 24415 24418
0 24420 5 1 1 24419
0 24421 7 1 2 55355 24420
0 24422 7 1 2 24414 24421
0 24423 7 1 2 24390 24422
0 24424 7 1 2 24341 24423
0 24425 5 1 1 24424
0 24426 7 1 2 51588 24425
0 24427 7 2 2 24311 24426
0 24428 5 1 1 76239
0 24429 7 1 2 24207 24428
0 24430 5 1 1 24429
0 24431 7 1 2 50206 24430
0 24432 5 1 1 24431
0 24433 7 2 2 73248 70590
0 24434 7 2 2 66217 76197
0 24435 7 1 2 76241 76243
0 24436 5 1 1 24435
0 24437 7 1 2 71111 73518
0 24438 5 1 1 24437
0 24439 7 1 2 73441 68929
0 24440 5 1 1 24439
0 24441 7 1 2 24438 24440
0 24442 5 1 1 24441
0 24443 7 1 2 48757 24442
0 24444 5 1 1 24443
0 24445 7 1 2 75155 76143
0 24446 5 1 1 24445
0 24447 7 1 2 24444 24446
0 24448 5 2 1 24447
0 24449 7 1 2 51334 76245
0 24450 5 1 1 24449
0 24451 7 2 2 62488 75826
0 24452 5 1 1 76247
0 24453 7 1 2 24450 24452
0 24454 5 1 1 24453
0 24455 7 1 2 57318 24454
0 24456 5 1 1 24455
0 24457 7 1 2 71224 68930
0 24458 5 1 1 24457
0 24459 7 1 2 76020 24458
0 24460 5 2 1 24459
0 24461 7 1 2 76104 76249
0 24462 5 1 1 24461
0 24463 7 1 2 53306 76012
0 24464 5 1 1 24463
0 24465 7 1 2 70812 72441
0 24466 5 1 1 24465
0 24467 7 1 2 24464 24466
0 24468 5 1 1 24467
0 24469 7 1 2 75283 24468
0 24470 5 1 1 24469
0 24471 7 1 2 24462 24470
0 24472 7 1 2 24456 24471
0 24473 5 1 1 24472
0 24474 7 1 2 51589 24473
0 24475 5 1 1 24474
0 24476 7 1 2 24436 24475
0 24477 5 1 1 24476
0 24478 7 1 2 75210 24477
0 24479 5 1 1 24478
0 24480 7 1 2 24432 24479
0 24481 7 1 2 24151 24480
0 24482 5 1 1 24481
0 24483 7 1 2 50445 24482
0 24484 5 1 1 24483
0 24485 7 4 2 48758 58032
0 24486 7 2 2 53513 68873
0 24487 5 2 1 76255
0 24488 7 1 2 54312 62090
0 24489 5 2 1 24488
0 24490 7 2 2 62767 76259
0 24491 7 1 2 53307 76261
0 24492 5 1 1 24491
0 24493 7 1 2 76257 24492
0 24494 5 1 1 24493
0 24495 7 1 2 76251 24494
0 24496 5 1 1 24495
0 24497 7 3 2 55027 63205
0 24498 5 1 1 76263
0 24499 7 1 2 62768 76212
0 24500 5 1 1 24499
0 24501 7 1 2 24498 24500
0 24502 5 1 1 24501
0 24503 7 1 2 52510 24502
0 24504 5 1 1 24503
0 24505 7 1 2 59362 75238
0 24506 7 1 2 73451 24505
0 24507 5 1 1 24506
0 24508 7 1 2 24504 24507
0 24509 5 1 1 24508
0 24510 7 1 2 75413 24509
0 24511 5 1 1 24510
0 24512 7 1 2 75228 76262
0 24513 5 1 1 24512
0 24514 7 3 2 50207 68931
0 24515 7 1 2 54313 62114
0 24516 5 2 1 24515
0 24517 7 1 2 76266 76269
0 24518 5 1 1 24517
0 24519 7 1 2 63562 24518
0 24520 5 1 1 24519
0 24521 7 1 2 75871 24520
0 24522 5 1 1 24521
0 24523 7 1 2 24513 24522
0 24524 7 1 2 24511 24523
0 24525 7 1 2 24496 24524
0 24526 5 1 1 24525
0 24527 7 1 2 52396 24526
0 24528 5 1 1 24527
0 24529 7 3 2 59881 70532
0 24530 7 2 2 62083 76271
0 24531 7 1 2 75229 76274
0 24532 5 1 1 24531
0 24533 7 1 2 53308 76275
0 24534 5 1 1 24533
0 24535 7 1 2 17756 24534
0 24536 5 1 1 24535
0 24537 7 1 2 76252 24536
0 24538 5 1 1 24537
0 24539 7 1 2 24532 24538
0 24540 5 1 1 24539
0 24541 7 1 2 50755 24540
0 24542 5 1 1 24541
0 24543 7 1 2 24528 24542
0 24544 5 1 1 24543
0 24545 7 1 2 53181 24544
0 24546 5 1 1 24545
0 24547 7 1 2 49562 73590
0 24548 5 1 1 24547
0 24549 7 1 2 75385 24548
0 24550 5 1 1 24549
0 24551 7 1 2 62169 24550
0 24552 5 1 1 24551
0 24553 7 2 2 70887 76270
0 24554 7 1 2 76096 76276
0 24555 5 1 1 24554
0 24556 7 1 2 63563 24555
0 24557 5 1 1 24556
0 24558 7 1 2 58033 24557
0 24559 5 1 1 24558
0 24560 7 1 2 59144 76213
0 24561 5 3 1 24560
0 24562 7 1 2 75386 76278
0 24563 5 1 1 24562
0 24564 7 1 2 62341 24563
0 24565 5 1 1 24564
0 24566 7 1 2 57781 75836
0 24567 5 1 1 24566
0 24568 7 2 2 49563 63640
0 24569 7 1 2 71201 76281
0 24570 5 1 1 24569
0 24571 7 1 2 24567 24570
0 24572 7 1 2 24565 24571
0 24573 7 1 2 24559 24572
0 24574 7 1 2 24552 24573
0 24575 5 1 1 24574
0 24576 7 1 2 53514 24575
0 24577 5 1 1 24576
0 24578 7 1 2 62170 73463
0 24579 5 2 1 24578
0 24580 7 1 2 62875 71608
0 24581 5 2 1 24580
0 24582 7 1 2 52975 76285
0 24583 5 1 1 24582
0 24584 7 1 2 76283 24583
0 24585 5 1 1 24584
0 24586 7 1 2 56455 62679
0 24587 7 1 2 24585 24586
0 24588 5 1 1 24587
0 24589 7 1 2 24577 24588
0 24590 5 1 1 24589
0 24591 7 1 2 48759 24590
0 24592 5 1 1 24591
0 24593 7 1 2 24546 24592
0 24594 5 1 1 24593
0 24595 7 1 2 51335 24594
0 24596 5 1 1 24595
0 24597 7 2 2 62084 76218
0 24598 5 1 1 76287
0 24599 7 1 2 48760 76288
0 24600 5 1 1 24599
0 24601 7 3 2 52511 75239
0 24602 5 4 1 76289
0 24603 7 1 2 48190 65560
0 24604 5 2 1 24603
0 24605 7 1 2 63943 59786
0 24606 5 1 1 24605
0 24607 7 2 2 76296 24606
0 24608 5 1 1 76298
0 24609 7 1 2 51933 76299
0 24610 5 1 1 24609
0 24611 7 1 2 50208 61470
0 24612 5 1 1 24611
0 24613 7 1 2 24610 24612
0 24614 5 3 1 24613
0 24615 7 1 2 52397 75258
0 24616 7 1 2 76300 24615
0 24617 5 1 1 24616
0 24618 7 1 2 76292 24617
0 24619 5 1 1 24618
0 24620 7 1 2 53182 24619
0 24621 5 1 1 24620
0 24622 7 2 2 73223 75211
0 24623 5 1 1 76303
0 24624 7 1 2 48761 76304
0 24625 5 1 1 24624
0 24626 7 1 2 24621 24625
0 24627 5 1 1 24626
0 24628 7 1 2 50756 24627
0 24629 5 1 1 24628
0 24630 7 1 2 49439 76066
0 24631 5 1 1 24630
0 24632 7 2 2 73420 24631
0 24633 5 1 1 76305
0 24634 7 1 2 48762 76306
0 24635 5 1 1 24634
0 24636 7 1 2 24629 24635
0 24637 5 1 1 24636
0 24638 7 1 2 50446 24637
0 24639 5 1 1 24638
0 24640 7 1 2 24600 24639
0 24641 5 1 1 24640
0 24642 7 1 2 72888 24641
0 24643 5 1 1 24642
0 24644 7 2 2 24596 24643
0 24645 5 1 1 76307
0 24646 7 1 2 75831 76301
0 24647 5 1 1 24646
0 24648 7 1 2 56555 24647
0 24649 5 1 1 24648
0 24650 7 1 2 53183 24649
0 24651 5 1 1 24650
0 24652 7 1 2 24623 24651
0 24653 5 1 1 24652
0 24654 7 1 2 50757 24653
0 24655 5 1 1 24654
0 24656 7 1 2 24633 24655
0 24657 5 1 1 24656
0 24658 7 1 2 50447 24657
0 24659 5 1 1 24658
0 24660 7 1 2 24598 24659
0 24661 5 1 1 24660
0 24662 7 2 2 51042 24661
0 24663 5 1 1 76309
0 24664 7 1 2 49757 76310
0 24665 5 1 1 24664
0 24666 7 1 2 48615 75139
0 24667 5 1 1 24666
0 24668 7 1 2 50448 75318
0 24669 5 1 1 24668
0 24670 7 1 2 48191 24669
0 24671 5 1 1 24670
0 24672 7 1 2 75190 24671
0 24673 5 1 1 24672
0 24674 7 1 2 65004 60641
0 24675 5 1 1 24674
0 24676 7 2 2 54662 24675
0 24677 5 1 1 76311
0 24678 7 1 2 24673 76312
0 24679 5 1 1 24678
0 24680 7 2 2 60580 24679
0 24681 7 1 2 52398 76313
0 24682 5 1 1 24681
0 24683 7 1 2 24667 24682
0 24684 5 1 1 24683
0 24685 7 1 2 53184 24684
0 24686 5 1 1 24685
0 24687 7 1 2 52976 58270
0 24688 7 1 2 60243 24687
0 24689 7 1 2 74857 24688
0 24690 5 1 1 24689
0 24691 7 1 2 75628 24690
0 24692 5 1 1 24691
0 24693 7 1 2 63513 24692
0 24694 5 1 1 24693
0 24695 7 4 2 50449 68932
0 24696 5 2 1 76315
0 24697 7 1 2 70888 76316
0 24698 5 1 1 24697
0 24699 7 1 2 24694 24698
0 24700 5 1 1 24699
0 24701 7 1 2 49440 24700
0 24702 5 1 1 24701
0 24703 7 4 2 51043 60203
0 24704 7 1 2 48616 76321
0 24705 5 1 1 24704
0 24706 7 1 2 52512 76314
0 24707 5 1 1 24706
0 24708 7 1 2 24705 24707
0 24709 7 1 2 24702 24708
0 24710 7 1 2 24686 24709
0 24711 5 1 1 24710
0 24712 7 1 2 53309 24711
0 24713 5 1 1 24712
0 24714 7 6 2 53185 55028
0 24715 5 1 1 76325
0 24716 7 2 2 76326 75721
0 24717 5 1 1 76331
0 24718 7 2 2 51044 76214
0 24719 7 1 2 52144 76333
0 24720 5 1 1 24719
0 24721 7 1 2 24717 24720
0 24722 5 1 1 24721
0 24723 7 1 2 52399 24722
0 24724 5 1 1 24723
0 24725 7 1 2 76279 24724
0 24726 5 2 1 24725
0 24727 7 1 2 62171 76335
0 24728 5 1 1 24727
0 24729 7 1 2 76280 76231
0 24730 5 1 1 24729
0 24731 7 1 2 52145 24730
0 24732 5 1 1 24731
0 24733 7 1 2 57319 67330
0 24734 5 1 1 24733
0 24735 7 1 2 71202 76332
0 24736 5 1 1 24735
0 24737 7 1 2 24734 24736
0 24738 7 1 2 24732 24737
0 24739 7 1 2 24728 24738
0 24740 5 1 1 24739
0 24741 7 1 2 50450 24740
0 24742 5 1 1 24741
0 24743 7 2 2 52400 60121
0 24744 7 5 2 52890 53186
0 24745 7 1 2 76339 75301
0 24746 7 1 2 75981 24745
0 24747 7 1 2 76337 24746
0 24748 5 1 1 24747
0 24749 7 1 2 24742 24748
0 24750 5 1 1 24749
0 24751 7 1 2 50209 24750
0 24752 5 1 1 24751
0 24753 7 1 2 76260 76334
0 24754 5 1 1 24753
0 24755 7 1 2 56208 60581
0 24756 7 1 2 24677 24755
0 24757 5 1 1 24756
0 24758 7 1 2 24754 24757
0 24759 5 1 1 24758
0 24760 7 1 2 52513 24759
0 24761 5 1 1 24760
0 24762 7 1 2 49441 61260
0 24763 5 1 1 24762
0 24764 7 1 2 50451 24763
0 24765 5 1 1 24764
0 24766 7 1 2 62172 73411
0 24767 5 1 1 24766
0 24768 7 1 2 24765 24767
0 24769 5 1 1 24768
0 24770 7 1 2 75618 24769
0 24771 5 1 1 24770
0 24772 7 1 2 24761 24771
0 24773 7 1 2 24752 24772
0 24774 7 1 2 24713 24773
0 24775 5 1 1 24774
0 24776 7 1 2 53515 24775
0 24777 5 1 1 24776
0 24778 7 1 2 55356 24777
0 24779 7 1 2 24665 24778
0 24780 5 1 1 24779
0 24781 7 1 2 50758 63027
0 24782 5 1 1 24781
0 24783 7 1 2 76284 24782
0 24784 5 1 1 24783
0 24785 7 1 2 49564 24784
0 24786 5 1 1 24785
0 24787 7 6 2 53187 54663
0 24788 5 1 1 76344
0 24789 7 4 2 54314 76345
0 24790 5 1 1 76350
0 24791 7 1 2 49565 65339
0 24792 5 1 1 24791
0 24793 7 1 2 24790 24792
0 24794 5 1 1 24793
0 24795 7 1 2 52401 24794
0 24796 5 1 1 24795
0 24797 7 1 2 58034 58687
0 24798 5 1 1 24797
0 24799 7 1 2 51045 24798
0 24800 7 1 2 24796 24799
0 24801 7 2 2 24786 24800
0 24802 5 1 1 76354
0 24803 7 1 2 54315 75412
0 24804 5 1 1 24803
0 24805 7 1 2 52402 24804
0 24806 5 1 1 24805
0 24807 7 1 2 54664 24806
0 24808 5 1 1 24807
0 24809 7 1 2 53188 58035
0 24810 7 1 2 24808 24809
0 24811 5 1 1 24810
0 24812 7 2 2 62326 75315
0 24813 5 1 1 76356
0 24814 7 1 2 54316 76357
0 24815 5 2 1 24814
0 24816 7 1 2 56456 76358
0 24817 5 1 1 24816
0 24818 7 1 2 76277 76130
0 24819 5 1 1 24818
0 24820 7 1 2 55029 24819
0 24821 7 1 2 24817 24820
0 24822 7 1 2 24811 24821
0 24823 5 2 1 24822
0 24824 7 1 2 49758 76360
0 24825 7 1 2 24802 24824
0 24826 5 1 1 24825
0 24827 7 3 2 49566 63456
0 24828 7 1 2 62771 76362
0 24829 7 1 2 76359 24828
0 24830 5 1 1 24829
0 24831 7 1 2 51336 24830
0 24832 7 1 2 24826 24831
0 24833 5 1 1 24832
0 24834 7 1 2 52647 24833
0 24835 7 1 2 24780 24834
0 24836 5 1 1 24835
0 24837 7 1 2 76308 24836
0 24838 5 1 1 24837
0 24839 7 1 2 51590 24838
0 24840 5 1 1 24839
0 24841 7 3 2 48504 60244
0 24842 5 4 1 76365
0 24843 7 1 2 52146 76368
0 24844 5 2 1 24843
0 24845 7 1 2 10199 76372
0 24846 5 2 1 24845
0 24847 7 1 2 62173 76374
0 24848 5 1 1 24847
0 24849 7 1 2 54317 63031
0 24850 5 1 1 24849
0 24851 7 1 2 52403 24850
0 24852 5 1 1 24851
0 24853 7 1 2 24848 24852
0 24854 5 1 1 24853
0 24855 7 2 2 66312 24854
0 24856 7 2 2 53189 75897
0 24857 7 1 2 76376 76378
0 24858 5 1 1 24857
0 24859 7 1 2 24840 24858
0 24860 5 1 1 24859
0 24861 7 1 2 57611 24860
0 24862 5 1 1 24861
0 24863 7 1 2 54665 24417
0 24864 5 4 1 24863
0 24865 7 1 2 50210 76124
0 24866 5 1 1 24865
0 24867 7 1 2 60642 75639
0 24868 5 1 1 24867
0 24869 7 1 2 24866 24868
0 24870 5 1 1 24869
0 24871 7 1 2 75822 24870
0 24872 5 1 1 24871
0 24873 7 2 2 50211 67331
0 24874 5 1 1 76384
0 24875 7 1 2 75850 76385
0 24876 5 1 1 24875
0 24877 7 1 2 48763 23660
0 24878 5 2 1 24877
0 24879 7 7 2 53310 73522
0 24880 5 1 1 76388
0 24881 7 1 2 62047 76389
0 24882 5 1 1 24881
0 24883 7 1 2 49567 71228
0 24884 5 1 1 24883
0 24885 7 1 2 24882 24884
0 24886 5 1 1 24885
0 24887 7 1 2 51934 24886
0 24888 5 1 1 24887
0 24889 7 2 2 52891 53311
0 24890 7 1 2 62097 73523
0 24891 7 1 2 76395 24890
0 24892 5 1 1 24891
0 24893 7 1 2 24888 24892
0 24894 5 1 1 24893
0 24895 7 1 2 76386 24894
0 24896 5 1 1 24895
0 24897 7 1 2 24876 24896
0 24898 7 1 2 24872 24897
0 24899 5 1 1 24898
0 24900 7 1 2 50452 24899
0 24901 5 1 1 24900
0 24902 7 2 2 58526 58072
0 24903 5 1 1 76397
0 24904 7 1 2 76121 76398
0 24905 5 1 1 24904
0 24906 7 1 2 24901 24905
0 24907 5 1 1 24906
0 24908 7 1 2 49759 24907
0 24909 5 1 1 24908
0 24910 7 6 2 63384 71208
0 24911 7 1 2 75343 76399
0 24912 5 1 1 24911
0 24913 7 1 2 58036 70739
0 24914 5 1 1 24913
0 24915 7 1 2 48505 24914
0 24916 5 1 1 24915
0 24917 7 1 2 75019 76122
0 24918 7 1 2 24916 24917
0 24919 5 1 1 24918
0 24920 7 1 2 24912 24919
0 24921 5 1 1 24920
0 24922 7 1 2 63206 24921
0 24923 5 1 1 24922
0 24924 7 1 2 24909 24923
0 24925 5 1 1 24924
0 24926 7 1 2 51337 24925
0 24927 5 1 1 24926
0 24928 7 1 2 62489 75755
0 24929 5 1 1 24928
0 24930 7 1 2 52404 70740
0 24931 5 1 1 24930
0 24932 7 1 2 70853 24931
0 24933 5 1 1 24932
0 24934 7 1 2 75406 24933
0 24935 5 1 1 24934
0 24936 7 1 2 24929 24935
0 24937 5 1 1 24936
0 24938 7 1 2 68392 24937
0 24939 5 1 1 24938
0 24940 7 2 2 24927 24939
0 24941 5 1 1 76405
0 24942 7 1 2 66889 75298
0 24943 5 1 1 24942
0 24944 7 2 2 55357 75284
0 24945 7 1 2 52514 76407
0 24946 5 1 1 24945
0 24947 7 2 2 48764 66890
0 24948 5 1 1 76409
0 24949 7 1 2 75122 76410
0 24950 5 1 1 24949
0 24951 7 1 2 53312 24950
0 24952 7 1 2 24946 24951
0 24953 5 1 1 24952
0 24954 7 3 2 49760 66891
0 24955 5 1 1 76411
0 24956 7 1 2 73859 76412
0 24957 5 1 1 24956
0 24958 7 6 2 52648 69801
0 24959 5 2 1 76414
0 24960 7 1 2 49568 76420
0 24961 7 1 2 24957 24960
0 24962 5 1 1 24961
0 24963 7 1 2 52405 24962
0 24964 7 1 2 24953 24963
0 24965 5 1 1 24964
0 24966 7 1 2 50212 73109
0 24967 7 1 2 75407 24966
0 24968 5 1 1 24967
0 24969 7 1 2 24965 24968
0 24970 5 1 1 24969
0 24971 7 1 2 59902 24970
0 24972 5 1 1 24971
0 24973 7 1 2 24943 24972
0 24974 5 2 1 24973
0 24975 7 1 2 52147 76422
0 24976 5 1 1 24975
0 24977 7 3 2 68393 75408
0 24978 7 1 2 70889 76424
0 24979 5 1 1 24978
0 24980 7 1 2 24976 24979
0 24981 5 1 1 24980
0 24982 7 1 2 58431 24981
0 24983 5 1 1 24982
0 24984 7 5 2 52406 52892
0 24985 7 4 2 52148 76427
0 24986 7 1 2 60680 76432
0 24987 7 1 2 75259 24986
0 24988 5 1 1 24987
0 24989 7 1 2 76293 24988
0 24990 5 1 1 24989
0 24991 7 1 2 62680 24990
0 24992 5 1 1 24991
0 24993 7 1 2 55030 22210
0 24994 5 1 1 24993
0 24995 7 1 2 71119 75285
0 24996 7 1 2 24994 24995
0 24997 5 1 1 24996
0 24998 7 1 2 24992 24997
0 24999 5 1 1 24998
0 25000 7 1 2 50453 24999
0 25001 5 1 1 25000
0 25002 7 2 2 55031 75286
0 25003 7 1 2 75832 76436
0 25004 5 1 1 25003
0 25005 7 1 2 25001 25004
0 25006 5 2 1 25005
0 25007 7 1 2 51338 76438
0 25008 5 1 1 25007
0 25009 7 1 2 51935 70890
0 25010 5 1 1 25009
0 25011 7 1 2 70751 76369
0 25012 5 1 1 25011
0 25013 7 1 2 25010 25012
0 25014 5 1 1 25013
0 25015 7 2 2 76425 25014
0 25016 5 1 1 76440
0 25017 7 1 2 25008 25016
0 25018 7 1 2 24983 25017
0 25019 5 1 1 25018
0 25020 7 1 2 57612 25019
0 25021 5 1 1 25020
0 25022 7 1 2 76406 25021
0 25023 5 1 1 25022
0 25024 7 1 2 51591 25023
0 25025 5 1 1 25024
0 25026 7 3 2 50213 58527
0 25027 5 1 1 76442
0 25028 7 3 2 73771 76443
0 25029 5 1 1 76445
0 25030 7 1 2 75887 76446
0 25031 5 1 1 25030
0 25032 7 3 2 52407 51339
0 25033 5 1 1 76448
0 25034 7 1 2 9587 25033
0 25035 5 1 1 25034
0 25036 7 1 2 55912 25035
0 25037 5 1 1 25036
0 25038 7 4 2 52408 52649
0 25039 5 2 1 76451
0 25040 7 1 2 55358 76455
0 25041 5 1 1 25040
0 25042 7 1 2 52515 25041
0 25043 5 1 1 25042
0 25044 7 1 2 25037 25043
0 25045 5 1 1 25044
0 25046 7 1 2 53313 73502
0 25047 7 1 2 25045 25046
0 25048 5 1 1 25047
0 25049 7 1 2 72442 76387
0 25050 5 1 1 25049
0 25051 7 1 2 49761 25050
0 25052 7 1 2 25048 25051
0 25053 5 1 1 25052
0 25054 7 3 2 51046 65005
0 25055 7 2 2 75508 76294
0 25056 5 2 1 76460
0 25057 7 2 2 55359 58528
0 25058 5 1 1 76464
0 25059 7 1 2 76462 76465
0 25060 5 1 1 25059
0 25061 7 3 2 48765 51340
0 25062 7 1 2 49569 76466
0 25063 5 1 1 25062
0 25064 7 1 2 53516 25063
0 25065 7 1 2 25060 25064
0 25066 5 1 1 25065
0 25067 7 1 2 76457 25066
0 25068 7 1 2 25053 25067
0 25069 5 1 1 25068
0 25070 7 1 2 25031 25069
0 25071 5 1 1 25070
0 25072 7 1 2 51592 25071
0 25073 5 1 1 25072
0 25074 7 3 2 73271 71303
0 25075 7 1 2 53314 63658
0 25076 7 1 2 66218 25075
0 25077 7 1 2 76469 25076
0 25078 5 1 1 25077
0 25079 7 1 2 25073 25078
0 25080 5 1 1 25079
0 25081 7 1 2 60983 25080
0 25082 5 1 1 25081
0 25083 7 3 2 53315 68394
0 25084 7 1 2 70152 76472
0 25085 5 1 1 25084
0 25086 7 1 2 58037 73120
0 25087 7 1 2 63806 25086
0 25088 5 1 1 25087
0 25089 7 1 2 25085 25088
0 25090 5 1 1 25089
0 25091 7 1 2 75287 25090
0 25092 5 1 1 25091
0 25093 7 1 2 52409 76248
0 25094 5 1 1 25093
0 25095 7 1 2 25092 25094
0 25096 5 1 1 25095
0 25097 7 1 2 57613 25096
0 25098 5 1 1 25097
0 25099 7 2 2 71214 76081
0 25100 5 1 1 76475
0 25101 7 1 2 73903 76476
0 25102 5 1 1 25101
0 25103 7 1 2 51341 73772
0 25104 5 1 1 25103
0 25105 7 1 2 25102 25104
0 25106 5 1 1 25105
0 25107 7 1 2 75288 25106
0 25108 5 1 1 25107
0 25109 7 2 2 64819 59353
0 25110 7 2 2 52650 52893
0 25111 5 1 1 76479
0 25112 7 2 2 50099 76480
0 25113 5 1 1 76481
0 25114 7 1 2 51936 76482
0 25115 7 1 2 76477 25114
0 25116 5 1 1 25115
0 25117 7 1 2 25108 25116
0 25118 5 1 1 25117
0 25119 7 1 2 58529 25118
0 25120 5 1 1 25119
0 25121 7 1 2 25098 25120
0 25122 5 2 1 25121
0 25123 7 1 2 51593 76483
0 25124 5 1 1 25123
0 25125 7 2 2 51937 71090
0 25126 7 1 2 76485 76082
0 25127 7 2 2 60098 75335
0 25128 7 2 2 66098 73821
0 25129 7 1 2 76487 76489
0 25130 7 2 2 25126 25129
0 25131 5 1 1 76491
0 25132 7 1 2 25124 25131
0 25133 5 1 1 25132
0 25134 7 1 2 60340 25133
0 25135 5 1 1 25134
0 25136 7 2 2 59354 75041
0 25137 7 2 2 73249 70601
0 25138 7 1 2 76493 76495
0 25139 5 1 1 25138
0 25140 7 1 2 58432 71505
0 25141 7 2 2 76338 25140
0 25142 7 1 2 76494 76497
0 25143 5 1 1 25142
0 25144 7 2 2 66118 73166
0 25145 7 1 2 70443 75988
0 25146 7 1 2 76499 25145
0 25147 5 1 1 25146
0 25148 7 1 2 25143 25147
0 25149 5 1 1 25148
0 25150 7 1 2 57614 25149
0 25151 5 1 1 25150
0 25152 7 1 2 25139 25151
0 25153 7 1 2 25135 25152
0 25154 7 1 2 25082 25153
0 25155 7 1 2 25025 25154
0 25156 5 1 1 25155
0 25157 7 1 2 76380 25156
0 25158 5 1 1 25157
0 25159 7 1 2 75260 76449
0 25160 5 1 1 25159
0 25161 7 4 2 70591 75803
0 25162 5 1 1 76501
0 25163 7 1 2 25160 25162
0 25164 5 1 1 25163
0 25165 7 1 2 49762 25164
0 25166 5 1 1 25165
0 25167 7 1 2 69802 76463
0 25168 5 1 1 25167
0 25169 7 1 2 25166 25168
0 25170 5 1 1 25169
0 25171 7 1 2 53190 25170
0 25172 5 1 1 25171
0 25173 7 1 2 48766 75880
0 25174 5 1 1 25173
0 25175 7 1 2 49763 75501
0 25176 5 1 1 25175
0 25177 7 1 2 25174 25176
0 25178 5 2 1 25177
0 25179 7 1 2 51342 76505
0 25180 5 1 1 25179
0 25181 7 1 2 25172 25180
0 25182 5 1 1 25181
0 25183 7 1 2 50759 25182
0 25184 5 1 1 25183
0 25185 7 2 2 64329 75435
0 25186 5 1 1 76507
0 25187 7 1 2 75235 25186
0 25188 5 1 1 25187
0 25189 7 2 2 69803 25188
0 25190 5 1 1 76509
0 25191 7 1 2 75636 76510
0 25192 5 1 1 25191
0 25193 7 1 2 25184 25192
0 25194 5 1 1 25193
0 25195 7 1 2 50214 25194
0 25196 5 1 1 25195
0 25197 7 1 2 53316 14010
0 25198 5 4 1 25197
0 25199 7 1 2 67977 76511
0 25200 5 1 1 25199
0 25201 7 1 2 76191 25200
0 25202 5 1 1 25201
0 25203 7 1 2 52651 25202
0 25204 5 1 1 25203
0 25205 7 1 2 76193 25204
0 25206 5 1 1 25205
0 25207 7 1 2 73110 25206
0 25208 5 1 1 25207
0 25209 7 1 2 25196 25208
0 25210 5 1 1 25209
0 25211 7 1 2 51047 25210
0 25212 5 1 1 25211
0 25213 7 1 2 61351 63207
0 25214 5 1 1 25213
0 25215 7 1 2 70341 25214
0 25216 5 1 1 25215
0 25217 7 1 2 65340 73129
0 25218 7 1 2 25216 25217
0 25219 5 1 1 25218
0 25220 7 1 2 25212 25219
0 25221 5 1 1 25220
0 25222 7 1 2 57615 25221
0 25223 5 1 1 25222
0 25224 7 1 2 68305 75798
0 25225 5 1 1 25224
0 25226 7 1 2 51343 75873
0 25227 5 1 1 25226
0 25228 7 1 2 25225 25227
0 25229 5 1 1 25228
0 25230 7 1 2 52652 25229
0 25231 5 1 1 25230
0 25232 7 1 2 67809 76290
0 25233 5 1 1 25232
0 25234 7 1 2 25231 25233
0 25235 5 1 1 25234
0 25236 7 1 2 70249 25235
0 25237 5 1 1 25236
0 25238 7 2 2 53191 63608
0 25239 5 2 1 76515
0 25240 7 1 2 52977 59761
0 25241 5 1 1 25240
0 25242 7 1 2 66355 25241
0 25243 5 1 1 25242
0 25244 7 1 2 52410 25243
0 25245 5 1 1 25244
0 25246 7 1 2 76517 25245
0 25247 5 1 1 25246
0 25248 7 1 2 75888 25247
0 25249 5 1 1 25248
0 25250 7 1 2 63178 63783
0 25251 7 1 2 75894 25250
0 25252 5 1 1 25251
0 25253 7 1 2 25249 25252
0 25254 5 1 1 25253
0 25255 7 1 2 58038 25254
0 25256 5 1 1 25255
0 25257 7 2 2 62490 64791
0 25258 5 1 1 76519
0 25259 7 4 2 52411 75853
0 25260 7 1 2 73364 76521
0 25261 5 2 1 25260
0 25262 7 1 2 25258 76525
0 25263 5 1 1 25262
0 25264 7 1 2 56457 25263
0 25265 5 1 1 25264
0 25266 7 3 2 52287 51344
0 25267 5 1 1 76527
0 25268 7 3 2 70772 76528
0 25269 5 1 1 76530
0 25270 7 1 2 75289 76531
0 25271 5 1 1 25270
0 25272 7 1 2 25265 25271
0 25273 5 1 1 25272
0 25274 7 1 2 63609 25273
0 25275 5 1 1 25274
0 25276 7 1 2 25256 25275
0 25277 7 1 2 25237 25276
0 25278 5 1 1 25277
0 25279 7 1 2 55032 25278
0 25280 5 1 1 25279
0 25281 7 4 2 48767 68586
0 25282 5 2 1 76533
0 25283 7 1 2 55913 76408
0 25284 5 1 1 25283
0 25285 7 1 2 76537 25284
0 25286 5 1 1 25285
0 25287 7 1 2 70113 25286
0 25288 5 1 1 25287
0 25289 7 1 2 72443 75931
0 25290 5 1 1 25289
0 25291 7 4 2 62972 9311
0 25292 7 1 2 73091 15707
0 25293 7 1 2 76539 25292
0 25294 5 1 1 25293
0 25295 7 1 2 25290 25294
0 25296 7 1 2 25288 25295
0 25297 5 1 1 25296
0 25298 7 1 2 65341 59145
0 25299 7 1 2 25297 25298
0 25300 5 1 1 25299
0 25301 7 1 2 25280 25300
0 25302 7 1 2 25223 25301
0 25303 5 2 1 25302
0 25304 7 1 2 51594 76543
0 25305 5 1 1 25304
0 25306 7 2 2 53192 76452
0 25307 5 1 1 76545
0 25308 7 2 2 73224 76546
0 25309 7 3 2 59355 66099
0 25310 5 1 1 76549
0 25311 7 1 2 60540 76550
0 25312 7 1 2 76547 25311
0 25313 5 1 1 25312
0 25314 7 4 2 52653 50215
0 25315 5 1 1 76552
0 25316 7 1 2 64463 76553
0 25317 7 1 2 70168 76551
0 25318 7 1 2 25316 25317
0 25319 5 1 1 25318
0 25320 7 1 2 25313 25319
0 25321 7 1 2 25305 25320
0 25322 5 1 1 25321
0 25323 7 1 2 62269 25322
0 25324 5 1 1 25323
0 25325 7 2 2 47931 62055
0 25326 5 1 1 76556
0 25327 7 8 2 61183 25326
0 25328 5 5 1 76558
0 25329 7 1 2 65295 75494
0 25330 5 1 1 25329
0 25331 7 2 2 48768 63659
0 25332 5 1 1 76571
0 25333 7 1 2 25330 25332
0 25334 5 1 1 25333
0 25335 7 1 2 52978 25334
0 25336 5 1 1 25335
0 25337 7 6 2 53317 60541
0 25338 7 1 2 75854 76573
0 25339 5 1 1 25338
0 25340 7 1 2 25336 25339
0 25341 5 1 1 25340
0 25342 7 1 2 52516 25341
0 25343 5 1 1 25342
0 25344 7 1 2 62369 10223
0 25345 5 3 1 25344
0 25346 7 1 2 76572 76579
0 25347 5 1 1 25346
0 25348 7 1 2 25343 25347
0 25349 5 1 1 25348
0 25350 7 1 2 63734 25349
0 25351 5 1 1 25350
0 25352 7 5 2 50216 55360
0 25353 7 1 2 51048 76582
0 25354 7 1 2 75868 25353
0 25355 5 1 1 25354
0 25356 7 1 2 25351 25355
0 25357 5 1 1 25356
0 25358 7 1 2 52412 25357
0 25359 5 1 1 25358
0 25360 7 4 2 55361 73822
0 25361 7 1 2 62633 76587
0 25362 5 1 1 25361
0 25363 7 1 2 58803 67528
0 25364 5 2 1 25363
0 25365 7 1 2 25362 76591
0 25366 5 1 1 25365
0 25367 7 1 2 52654 25366
0 25368 5 1 1 25367
0 25369 7 1 2 63208 73867
0 25370 5 1 1 25369
0 25371 7 1 2 25368 25370
0 25372 5 1 1 25371
0 25373 7 1 2 76097 25372
0 25374 5 1 1 25373
0 25375 7 1 2 76478 76554
0 25376 5 1 1 25375
0 25377 7 1 2 25374 25376
0 25378 5 1 1 25377
0 25379 7 1 2 57320 25378
0 25380 5 1 1 25379
0 25381 7 2 2 49442 63179
0 25382 5 1 1 76593
0 25383 7 2 2 63514 73823
0 25384 5 1 1 76595
0 25385 7 1 2 76594 76596
0 25386 5 1 1 25385
0 25387 7 1 2 59882 75484
0 25388 5 2 1 25387
0 25389 7 3 2 55033 68306
0 25390 7 1 2 65342 76599
0 25391 5 1 1 25390
0 25392 7 1 2 76597 25391
0 25393 5 1 1 25392
0 25394 7 1 2 71188 25393
0 25395 5 1 1 25394
0 25396 7 1 2 25386 25395
0 25397 5 1 1 25396
0 25398 7 1 2 55362 25397
0 25399 5 1 1 25398
0 25400 7 2 2 49764 63735
0 25401 7 2 2 53318 63610
0 25402 5 1 1 76604
0 25403 7 1 2 50454 75833
0 25404 5 1 1 25403
0 25405 7 1 2 25402 25404
0 25406 5 1 1 25405
0 25407 7 1 2 52979 25406
0 25408 5 1 1 25407
0 25409 7 1 2 71614 25408
0 25410 5 1 1 25409
0 25411 7 1 2 76602 25410
0 25412 5 1 1 25411
0 25413 7 1 2 25399 25412
0 25414 5 1 1 25413
0 25415 7 1 2 52655 25414
0 25416 5 1 1 25415
0 25417 7 1 2 73442 75240
0 25418 7 1 2 74979 25417
0 25419 5 1 1 25418
0 25420 7 1 2 25416 25419
0 25421 7 1 2 25380 25420
0 25422 7 1 2 25359 25421
0 25423 5 2 1 25422
0 25424 7 1 2 57616 76606
0 25425 5 1 1 25424
0 25426 7 1 2 63628 71609
0 25427 5 2 1 25426
0 25428 7 1 2 72444 76608
0 25429 5 1 1 25428
0 25430 7 1 2 63611 72623
0 25431 5 1 1 25430
0 25432 7 1 2 55363 10076
0 25433 7 1 2 25431 25432
0 25434 5 1 1 25433
0 25435 7 1 2 51345 22617
0 25436 5 1 1 25435
0 25437 7 1 2 55914 25436
0 25438 7 1 2 25434 25437
0 25439 5 1 1 25438
0 25440 7 1 2 25429 25439
0 25441 5 1 1 25440
0 25442 7 1 2 52980 25441
0 25443 5 1 1 25442
0 25444 7 1 2 53193 73749
0 25445 7 1 2 75790 25444
0 25446 5 1 1 25445
0 25447 7 1 2 25443 25446
0 25448 5 1 1 25447
0 25449 7 1 2 51049 25448
0 25450 5 1 1 25449
0 25451 7 2 2 67529 76189
0 25452 5 1 1 76610
0 25453 7 1 2 49765 25452
0 25454 7 1 2 25450 25453
0 25455 5 1 1 25454
0 25456 7 1 2 50217 75800
0 25457 5 1 1 25456
0 25458 7 10 2 49443 53319
0 25459 5 1 1 76612
0 25460 7 2 2 52981 76613
0 25461 7 1 2 62610 68395
0 25462 7 1 2 76622 25461
0 25463 5 1 1 25462
0 25464 7 1 2 25457 25463
0 25465 5 1 1 25464
0 25466 7 1 2 54666 25465
0 25467 5 1 1 25466
0 25468 7 1 2 52517 50455
0 25469 5 2 1 25468
0 25470 7 1 2 55915 76609
0 25471 5 1 1 25470
0 25472 7 1 2 76624 25471
0 25473 5 1 1 25472
0 25474 7 1 2 52982 25473
0 25475 5 1 1 25474
0 25476 7 1 2 72981 25475
0 25477 5 1 1 25476
0 25478 7 1 2 75827 25477
0 25479 5 1 1 25478
0 25480 7 1 2 53517 25479
0 25481 7 1 2 25467 25480
0 25482 5 1 1 25481
0 25483 7 1 2 52656 25482
0 25484 7 1 2 25455 25483
0 25485 5 1 1 25484
0 25486 7 1 2 75971 76588
0 25487 5 1 1 25486
0 25488 7 1 2 52983 75881
0 25489 5 1 1 25488
0 25490 7 1 2 75859 25489
0 25491 5 1 1 25490
0 25492 7 1 2 51346 58530
0 25493 7 1 2 25491 25492
0 25494 5 1 1 25493
0 25495 7 1 2 25487 25494
0 25496 5 1 1 25495
0 25497 7 1 2 50456 25496
0 25498 5 1 1 25497
0 25499 7 1 2 70114 75101
0 25500 5 1 1 25499
0 25501 7 1 2 49570 67810
0 25502 5 1 1 25501
0 25503 7 1 2 25500 25502
0 25504 5 1 1 25503
0 25505 7 1 2 74887 25504
0 25506 5 1 1 25505
0 25507 7 1 2 25498 25506
0 25508 5 1 1 25507
0 25509 7 1 2 51050 25508
0 25510 5 1 1 25509
0 25511 7 1 2 53518 76611
0 25512 5 1 1 25511
0 25513 7 1 2 25510 25512
0 25514 5 1 1 25513
0 25515 7 1 2 48769 25514
0 25516 5 1 1 25515
0 25517 7 3 2 52413 70250
0 25518 5 1 1 76626
0 25519 7 1 2 75102 76627
0 25520 5 1 1 25519
0 25521 7 1 2 55916 76413
0 25522 5 1 1 25521
0 25523 7 1 2 25520 25522
0 25524 5 1 1 25523
0 25525 7 1 2 76126 25524
0 25526 5 1 1 25525
0 25527 7 1 2 25516 25526
0 25528 7 2 2 25485 25527
0 25529 5 1 1 76629
0 25530 7 1 2 25425 76630
0 25531 5 1 1 25530
0 25532 7 1 2 51595 25531
0 25533 5 1 1 25532
0 25534 7 1 2 61137 25518
0 25535 5 1 1 25534
0 25536 7 2 2 66313 25535
0 25537 7 1 2 76379 76631
0 25538 5 1 1 25537
0 25539 7 1 2 25533 25538
0 25540 5 1 1 25539
0 25541 7 1 2 76559 25540
0 25542 5 1 1 25541
0 25543 7 3 2 71189 73481
0 25544 7 1 2 76148 76633
0 25545 5 1 1 25544
0 25546 7 3 2 67680 69410
0 25547 5 1 1 76636
0 25548 7 1 2 76219 76637
0 25549 5 1 1 25548
0 25550 7 2 2 49571 75964
0 25551 7 1 2 65987 76639
0 25552 5 1 1 25551
0 25553 7 5 2 53194 50100
0 25554 7 3 2 70540 76641
0 25555 7 3 2 51938 52518
0 25556 7 2 2 76646 76649
0 25557 7 1 2 75075 76652
0 25558 5 1 1 25557
0 25559 7 1 2 54667 66344
0 25560 5 1 1 25559
0 25561 7 1 2 25558 25560
0 25562 5 1 1 25561
0 25563 7 1 2 53320 24813
0 25564 7 1 2 25562 25563
0 25565 5 1 1 25564
0 25566 7 1 2 25552 25565
0 25567 5 1 1 25566
0 25568 7 1 2 51051 25567
0 25569 5 1 1 25568
0 25570 7 2 2 51596 76109
0 25571 5 1 1 76654
0 25572 7 1 2 25569 25571
0 25573 5 1 1 25572
0 25574 7 1 2 53519 25573
0 25575 5 1 1 25574
0 25576 7 1 2 25549 25575
0 25577 5 1 1 25576
0 25578 7 1 2 52657 25577
0 25579 5 1 1 25578
0 25580 7 1 2 60514 65988
0 25581 7 1 2 75479 25580
0 25582 7 1 2 59036 25581
0 25583 5 1 1 25582
0 25584 7 1 2 25579 25583
0 25585 5 1 1 25584
0 25586 7 1 2 58531 25585
0 25587 5 1 1 25586
0 25588 7 1 2 25545 25587
0 25589 7 1 2 25542 25588
0 25590 7 1 2 25324 25589
0 25591 7 1 2 25158 25590
0 25592 7 1 2 24862 25591
0 25593 7 1 2 24484 25592
0 25594 7 1 2 23937 25593
0 25595 7 1 2 22876 25594
0 25596 5 1 1 25595
0 25597 7 1 2 49936 25596
0 25598 5 1 1 25597
0 25599 7 6 2 49333 50457
0 25600 5 1 1 76656
0 25601 7 2 2 73921 25600
0 25602 5 3 1 76662
0 25603 7 4 2 52414 54668
0 25604 7 2 2 66040 76667
0 25605 7 1 2 76664 76671
0 25606 5 1 1 25605
0 25607 7 1 2 63186 62616
0 25608 5 3 1 25607
0 25609 7 3 2 75460 76673
0 25610 7 2 2 51939 76676
0 25611 5 1 1 76679
0 25612 7 1 2 53096 76680
0 25613 5 1 1 25612
0 25614 7 1 2 50458 55763
0 25615 5 2 1 25614
0 25616 7 2 2 50218 76681
0 25617 5 1 1 76683
0 25618 7 1 2 64875 59681
0 25619 7 1 2 76684 25618
0 25620 5 1 1 25619
0 25621 7 1 2 25613 25620
0 25622 5 1 1 25621
0 25623 7 1 2 49444 25622
0 25624 5 1 1 25623
0 25625 7 5 2 48506 53195
0 25626 5 3 1 76685
0 25627 7 1 2 63180 76686
0 25628 5 1 1 25627
0 25629 7 1 2 25624 25628
0 25630 5 1 1 25629
0 25631 7 1 2 52288 25630
0 25632 5 1 1 25631
0 25633 7 6 2 52415 49445
0 25634 5 2 1 76693
0 25635 7 2 2 76690 76699
0 25636 5 7 1 76701
0 25637 7 1 2 54318 59743
0 25638 5 1 1 25637
0 25639 7 1 2 25611 25638
0 25640 5 1 1 25639
0 25641 7 1 2 76703 25640
0 25642 5 1 1 25641
0 25643 7 2 2 59657 70541
0 25644 7 3 2 49446 50101
0 25645 7 1 2 48507 76712
0 25646 7 1 2 76710 25645
0 25647 5 1 1 25646
0 25648 7 1 2 25642 25647
0 25649 7 1 2 25632 25648
0 25650 5 1 1 25649
0 25651 7 1 2 50760 25650
0 25652 5 1 1 25651
0 25653 7 1 2 25606 25652
0 25654 5 2 1 25653
0 25655 7 1 2 53321 76715
0 25656 5 1 1 25655
0 25657 7 4 2 56209 75358
0 25658 5 1 1 76717
0 25659 7 1 2 63396 76718
0 25660 5 1 1 25659
0 25661 7 1 2 25656 25660
0 25662 5 1 1 25661
0 25663 7 1 2 57229 25662
0 25664 5 1 1 25663
0 25665 7 1 2 56109 62001
0 25666 5 1 1 25665
0 25667 7 2 2 74028 25666
0 25668 5 1 1 76721
0 25669 7 1 2 57617 76722
0 25670 5 2 1 25669
0 25671 7 1 2 72987 76723
0 25672 5 1 1 25671
0 25673 7 3 2 56356 70753
0 25674 5 1 1 76725
0 25675 7 3 2 54669 57011
0 25676 7 1 2 70626 76728
0 25677 7 1 2 25674 25676
0 25678 5 1 1 25677
0 25679 7 3 2 52149 62649
0 25680 5 1 1 76731
0 25681 7 1 2 53097 76732
0 25682 5 1 1 25681
0 25683 7 1 2 25678 25682
0 25684 5 1 1 25683
0 25685 7 1 2 51940 25684
0 25686 5 1 1 25685
0 25687 7 3 2 52150 54670
0 25688 7 1 2 56210 76734
0 25689 5 2 1 25688
0 25690 7 1 2 25686 76737
0 25691 5 1 1 25690
0 25692 7 1 2 52984 25691
0 25693 5 1 1 25692
0 25694 7 1 2 14203 25693
0 25695 5 1 1 25694
0 25696 7 1 2 70693 25695
0 25697 5 1 1 25696
0 25698 7 4 2 50761 57012
0 25699 5 4 1 76739
0 25700 7 2 2 76428 76642
0 25701 5 1 1 76747
0 25702 7 2 2 76743 25701
0 25703 5 1 1 76749
0 25704 7 1 2 56110 73458
0 25705 5 1 1 25704
0 25706 7 1 2 14280 25705
0 25707 7 1 2 25703 25706
0 25708 5 1 1 25707
0 25709 7 1 2 61054 62103
0 25710 5 1 1 25709
0 25711 7 3 2 50762 76704
0 25712 5 1 1 76751
0 25713 7 2 2 52894 76752
0 25714 7 1 2 25710 76754
0 25715 5 1 1 25714
0 25716 7 2 2 52895 72965
0 25717 5 1 1 76756
0 25718 7 1 2 76702 25717
0 25719 5 1 1 25718
0 25720 7 1 2 56740 60694
0 25721 5 4 1 25720
0 25722 7 1 2 59484 76758
0 25723 7 1 2 25719 25722
0 25724 5 1 1 25723
0 25725 7 4 2 50102 71418
0 25726 7 1 2 70632 76762
0 25727 5 1 1 25726
0 25728 7 1 2 25724 25727
0 25729 7 1 2 25715 25728
0 25730 5 1 1 25729
0 25731 7 1 2 57618 25730
0 25732 5 1 1 25731
0 25733 7 1 2 25708 25732
0 25734 7 1 2 25697 25733
0 25735 7 1 2 25672 25734
0 25736 5 1 1 25735
0 25737 7 1 2 54319 25736
0 25738 5 1 1 25737
0 25739 7 1 2 56741 62157
0 25740 5 2 1 25739
0 25741 7 1 2 62426 76766
0 25742 5 1 1 25741
0 25743 7 2 2 52416 49334
0 25744 7 1 2 53196 66251
0 25745 7 1 2 76768 25744
0 25746 7 1 2 25742 25745
0 25747 5 1 1 25746
0 25748 7 1 2 25738 25747
0 25749 5 2 1 25748
0 25750 7 1 2 53322 76770
0 25751 5 1 1 25750
0 25752 7 2 2 50219 60598
0 25753 7 4 2 50763 70767
0 25754 5 1 1 76774
0 25755 7 1 2 73265 76215
0 25756 7 1 2 76775 25755
0 25757 7 1 2 76772 25756
0 25758 5 1 1 25757
0 25759 7 1 2 25751 25758
0 25760 7 1 2 25664 25759
0 25761 5 1 1 25760
0 25762 7 1 2 51052 25761
0 25763 5 1 1 25762
0 25764 7 1 2 49213 74982
0 25765 5 4 1 25764
0 25766 7 1 2 54039 76755
0 25767 5 1 1 25766
0 25768 7 2 2 67396 70623
0 25769 7 1 2 54040 60775
0 25770 5 3 1 25769
0 25771 7 1 2 54671 76784
0 25772 7 1 2 76782 25771
0 25773 5 1 1 25772
0 25774 7 1 2 25767 25773
0 25775 5 2 1 25774
0 25776 7 1 2 53323 76787
0 25777 5 1 1 25776
0 25778 7 1 2 50220 63120
0 25779 5 1 1 25778
0 25780 7 1 2 13573 25779
0 25781 5 2 1 25780
0 25782 7 1 2 76719 76789
0 25783 5 1 1 25782
0 25784 7 1 2 25777 25783
0 25785 5 1 1 25784
0 25786 7 1 2 51053 25785
0 25787 5 1 1 25786
0 25788 7 2 2 60448 76267
0 25789 5 1 1 76791
0 25790 7 1 2 73298 76792
0 25791 5 1 1 25790
0 25792 7 1 2 25787 25791
0 25793 5 1 1 25792
0 25794 7 1 2 76778 25793
0 25795 5 1 1 25794
0 25796 7 2 2 49572 62357
0 25797 7 2 2 56629 71574
0 25798 7 2 2 76793 76795
0 25799 5 1 1 76797
0 25800 7 3 2 49335 60653
0 25801 5 2 1 76799
0 25802 7 2 2 52985 76802
0 25803 5 1 1 76804
0 25804 7 1 2 58892 76805
0 25805 5 1 1 25804
0 25806 7 1 2 66035 25805
0 25807 5 1 1 25806
0 25808 7 1 2 49447 25807
0 25809 5 1 1 25808
0 25810 7 4 2 48386 53197
0 25811 7 1 2 53098 76806
0 25812 7 1 2 76137 25811
0 25813 5 1 1 25812
0 25814 7 1 2 25809 25813
0 25815 5 1 1 25814
0 25816 7 1 2 50764 25815
0 25817 5 1 1 25816
0 25818 7 1 2 62216 72948
0 25819 7 1 2 76067 25818
0 25820 5 1 1 25819
0 25821 7 1 2 25817 25820
0 25822 5 1 1 25821
0 25823 7 1 2 54041 25822
0 25824 5 1 1 25823
0 25825 7 3 2 52986 49336
0 25826 5 1 1 76810
0 25827 7 1 2 76733 76811
0 25828 5 1 1 25827
0 25829 7 1 2 56357 60782
0 25830 5 1 1 25829
0 25831 7 1 2 9726 76729
0 25832 7 1 2 25830 25831
0 25833 5 1 1 25832
0 25834 7 1 2 25828 25833
0 25835 5 1 1 25834
0 25836 7 1 2 52289 25835
0 25837 5 1 1 25836
0 25838 7 1 2 59078 75316
0 25839 5 1 1 25838
0 25840 7 1 2 57502 62071
0 25841 5 1 1 25840
0 25842 7 1 2 1077 25841
0 25843 7 1 2 25839 25842
0 25844 5 1 1 25843
0 25845 7 1 2 50765 25844
0 25846 5 1 1 25845
0 25847 7 1 2 52417 70468
0 25848 7 1 2 61464 25847
0 25849 5 1 1 25848
0 25850 7 1 2 57743 66030
0 25851 5 1 1 25850
0 25852 7 1 2 75710 25851
0 25853 5 1 1 25852
0 25854 7 1 2 61976 25853
0 25855 5 1 1 25854
0 25856 7 1 2 49337 55764
0 25857 5 4 1 25856
0 25858 7 1 2 52418 64003
0 25859 7 1 2 76813 25858
0 25860 5 1 1 25859
0 25861 7 1 2 25855 25860
0 25862 7 1 2 25849 25861
0 25863 7 1 2 25846 25862
0 25864 5 1 1 25863
0 25865 7 1 2 53198 25864
0 25866 5 1 1 25865
0 25867 7 1 2 25837 25866
0 25868 5 1 1 25867
0 25869 7 1 2 50221 25868
0 25870 5 1 1 25869
0 25871 7 1 2 70469 70444
0 25872 5 1 1 25871
0 25873 7 1 2 4664 25872
0 25874 5 1 1 25873
0 25875 7 1 2 76705 25874
0 25876 5 1 1 25875
0 25877 7 3 2 49448 59744
0 25878 5 1 1 76817
0 25879 7 1 2 66689 76818
0 25880 5 1 1 25879
0 25881 7 1 2 56211 61025
0 25882 5 1 1 25881
0 25883 7 1 2 62193 60161
0 25884 7 1 2 60099 25883
0 25885 5 1 1 25884
0 25886 7 1 2 25882 25885
0 25887 5 1 1 25886
0 25888 7 1 2 51941 25887
0 25889 5 1 1 25888
0 25890 7 1 2 25880 25889
0 25891 7 1 2 25876 25890
0 25892 5 1 1 25891
0 25893 7 1 2 70367 25892
0 25894 5 1 1 25893
0 25895 7 1 2 52290 62085
0 25896 5 1 1 25895
0 25897 7 1 2 63612 25896
0 25898 5 1 1 25897
0 25899 7 1 2 72972 25898
0 25900 5 1 1 25899
0 25901 7 1 2 76706 25900
0 25902 5 1 1 25901
0 25903 7 2 2 53099 76346
0 25904 7 1 2 48387 71203
0 25905 7 1 2 76820 25904
0 25906 5 1 1 25905
0 25907 7 1 2 25902 25906
0 25908 7 1 2 25894 25907
0 25909 7 1 2 25870 25908
0 25910 7 1 2 25824 25909
0 25911 5 2 1 25910
0 25912 7 1 2 53324 76822
0 25913 5 1 1 25912
0 25914 7 1 2 25799 25913
0 25915 5 1 1 25914
0 25916 7 1 2 51054 25915
0 25917 5 1 1 25916
0 25918 7 1 2 25795 25917
0 25919 5 1 1 25918
0 25920 7 1 2 50459 25919
0 25921 5 1 1 25920
0 25922 7 1 2 63121 76753
0 25923 5 1 1 25922
0 25924 7 1 2 71091 76821
0 25925 5 1 1 25924
0 25926 7 1 2 25923 25925
0 25927 5 1 1 25926
0 25928 7 1 2 54320 25927
0 25929 5 1 1 25928
0 25930 7 1 2 57230 63988
0 25931 7 1 2 70624 25930
0 25932 7 1 2 73933 25931
0 25933 7 1 2 54672 67711
0 25934 5 2 1 25933
0 25935 7 1 2 49449 66036
0 25936 5 1 1 25935
0 25937 7 1 2 50766 25936
0 25938 5 1 1 25937
0 25939 7 1 2 76824 25938
0 25940 7 1 2 25932 25939
0 25941 5 1 1 25940
0 25942 7 1 2 25929 25941
0 25943 5 1 1 25942
0 25944 7 1 2 51942 25943
0 25945 5 1 1 25944
0 25946 7 2 2 59682 70251
0 25947 7 1 2 76672 76826
0 25948 5 1 1 25947
0 25949 7 1 2 62617 76035
0 25950 5 3 1 25949
0 25951 7 2 2 52151 76828
0 25952 5 1 1 76831
0 25953 7 1 2 56358 66645
0 25954 7 1 2 76832 25953
0 25955 5 1 1 25954
0 25956 7 1 2 50460 62194
0 25957 7 1 2 72680 25956
0 25958 5 1 1 25957
0 25959 7 1 2 25955 25958
0 25960 5 1 1 25959
0 25961 7 1 2 50767 25960
0 25962 5 1 1 25961
0 25963 7 1 2 25948 25962
0 25964 7 1 2 25945 25963
0 25965 5 2 1 25964
0 25966 7 1 2 53325 76833
0 25967 5 1 1 25966
0 25968 7 1 2 60453 71271
0 25969 5 1 1 25968
0 25970 7 1 2 61527 25969
0 25971 5 1 1 25970
0 25972 7 1 2 67463 25971
0 25973 5 1 1 25972
0 25974 7 1 2 76720 25973
0 25975 5 1 1 25974
0 25976 7 1 2 25967 25975
0 25977 5 1 1 25976
0 25978 7 1 2 51055 25977
0 25979 5 1 1 25978
0 25980 7 2 2 65296 76317
0 25981 7 1 2 60599 70879
0 25982 7 2 2 76835 25981
0 25983 5 1 1 76837
0 25984 7 1 2 53326 76838
0 25985 5 1 1 25984
0 25986 7 1 2 25979 25985
0 25987 5 1 1 25986
0 25988 7 1 2 58433 25987
0 25989 5 1 1 25988
0 25990 7 2 2 53327 57231
0 25991 7 1 2 63807 72648
0 25992 7 2 2 65938 25991
0 25993 5 1 1 76841
0 25994 7 2 2 56212 76842
0 25995 5 1 1 76843
0 25996 7 1 2 76839 76844
0 25997 5 1 1 25996
0 25998 7 1 2 54042 59821
0 25999 5 4 1 25998
0 26000 7 1 2 76738 25712
0 26001 5 1 1 26000
0 26002 7 1 2 54321 57619
0 26003 7 1 2 60943 26002
0 26004 7 1 2 26001 26003
0 26005 5 1 1 26004
0 26006 7 4 2 48192 58864
0 26007 5 8 1 76849
0 26008 7 1 2 62634 76853
0 26009 7 1 2 76783 26008
0 26010 5 1 1 26009
0 26011 7 1 2 26005 26010
0 26012 5 1 1 26011
0 26013 7 1 2 51056 26012
0 26014 5 1 1 26013
0 26015 7 4 2 51943 53199
0 26016 7 1 2 76433 76861
0 26017 7 1 2 74987 26016
0 26018 5 1 1 26017
0 26019 7 1 2 26014 26018
0 26020 5 2 1 26019
0 26021 7 1 2 53328 76865
0 26022 5 1 1 26021
0 26023 7 2 2 51944 60774
0 26024 5 1 1 76867
0 26025 7 1 2 56111 26024
0 26026 5 1 1 26025
0 26027 7 1 2 49573 59917
0 26028 7 1 2 71612 26027
0 26029 7 1 2 26026 26028
0 26030 5 1 1 26029
0 26031 7 1 2 26022 26030
0 26032 5 1 1 26031
0 26033 7 1 2 76845 26032
0 26034 5 1 1 26033
0 26035 7 1 2 25997 26034
0 26036 7 1 2 25989 26035
0 26037 7 1 2 25921 26036
0 26038 7 1 2 25763 26037
0 26039 5 1 1 26038
0 26040 7 1 2 48617 26039
0 26041 5 1 1 26040
0 26042 7 1 2 49338 72691
0 26043 5 2 1 26042
0 26044 7 1 2 56112 59798
0 26045 5 1 1 26044
0 26046 7 1 2 76869 26045
0 26047 5 1 1 26046
0 26048 7 1 2 54322 26047
0 26049 5 1 1 26048
0 26050 7 2 2 52291 55692
0 26051 5 2 1 76871
0 26052 7 1 2 76657 76873
0 26053 5 1 1 26052
0 26054 7 1 2 26049 26053
0 26055 5 1 1 26054
0 26056 7 1 2 52152 26055
0 26057 5 1 1 26056
0 26058 7 1 2 48193 58837
0 26059 7 1 2 76658 26058
0 26060 5 1 1 26059
0 26061 7 1 2 26057 26060
0 26062 5 1 1 26061
0 26063 7 1 2 52987 26062
0 26064 5 1 1 26063
0 26065 7 1 2 56630 61397
0 26066 5 1 1 26065
0 26067 7 2 2 65934 26066
0 26068 5 1 1 76875
0 26069 7 1 2 55765 62435
0 26070 5 1 1 26069
0 26071 7 1 2 26068 26070
0 26072 5 1 1 26071
0 26073 7 1 2 59658 26072
0 26074 5 1 1 26073
0 26075 7 1 2 52153 57782
0 26076 5 2 1 26075
0 26077 7 3 2 48194 53100
0 26078 5 1 1 76879
0 26079 7 1 2 71130 26078
0 26080 7 1 2 76877 26079
0 26081 5 1 1 26080
0 26082 7 1 2 26074 26081
0 26083 7 1 2 26064 26082
0 26084 5 1 1 26083
0 26085 7 1 2 50768 26084
0 26086 5 1 1 26085
0 26087 7 1 2 58818 62635
0 26088 7 1 2 58899 26087
0 26089 5 1 1 26088
0 26090 7 1 2 26086 26089
0 26091 5 1 1 26090
0 26092 7 1 2 49450 26091
0 26093 5 1 1 26092
0 26094 7 1 2 60167 63191
0 26095 5 1 1 26094
0 26096 7 1 2 58136 74873
0 26097 5 1 1 26096
0 26098 7 1 2 26095 26097
0 26099 5 1 1 26098
0 26100 7 1 2 60122 26099
0 26101 5 1 1 26100
0 26102 7 2 2 57620 59300
0 26103 7 2 2 62407 55766
0 26104 5 2 1 76884
0 26105 7 2 2 62151 76885
0 26106 5 1 1 76888
0 26107 7 1 2 76882 76889
0 26108 5 1 1 26107
0 26109 7 1 2 59079 59069
0 26110 5 1 1 26109
0 26111 7 1 2 26108 26110
0 26112 5 1 1 26111
0 26113 7 1 2 50461 26112
0 26114 5 1 1 26113
0 26115 7 1 2 26101 26114
0 26116 5 1 1 26115
0 26117 7 1 2 54673 26116
0 26118 5 1 1 26117
0 26119 7 1 2 67426 70419
0 26120 5 1 1 26119
0 26121 7 1 2 26118 26120
0 26122 5 1 1 26121
0 26123 7 1 2 53200 26122
0 26124 5 1 1 26123
0 26125 7 3 2 52896 49451
0 26126 7 2 2 59375 76890
0 26127 7 1 2 57621 58825
0 26128 7 1 2 76893 26127
0 26129 5 1 1 26128
0 26130 7 1 2 52988 66160
0 26131 7 1 2 76347 26130
0 26132 7 1 2 61123 26131
0 26133 7 1 2 71133 26132
0 26134 5 1 1 26133
0 26135 7 1 2 26129 26134
0 26136 5 1 1 26135
0 26137 7 1 2 52154 26136
0 26138 5 1 1 26137
0 26139 7 5 2 52292 49339
0 26140 5 1 1 76895
0 26141 7 1 2 63983 66350
0 26142 5 1 1 26141
0 26143 7 1 2 52989 76894
0 26144 5 1 1 26143
0 26145 7 1 2 26142 26144
0 26146 5 1 1 26145
0 26147 7 1 2 76896 26146
0 26148 5 1 1 26147
0 26149 7 1 2 62011 72608
0 26150 5 1 1 26149
0 26151 7 4 2 52293 49214
0 26152 5 1 1 76900
0 26153 7 2 2 52897 76901
0 26154 7 2 2 73919 76348
0 26155 7 1 2 76904 76906
0 26156 5 1 1 26155
0 26157 7 1 2 26150 26156
0 26158 5 1 1 26157
0 26159 7 1 2 48195 26158
0 26160 5 1 1 26159
0 26161 7 1 2 49215 70768
0 26162 7 1 2 63292 26161
0 26163 5 1 1 26162
0 26164 7 1 2 26160 26163
0 26165 7 1 2 26148 26164
0 26166 7 1 2 26138 26165
0 26167 5 1 1 26166
0 26168 7 1 2 51945 26167
0 26169 5 1 1 26168
0 26170 7 1 2 64330 72649
0 26171 5 1 1 26170
0 26172 7 1 2 63293 76340
0 26173 5 1 1 26172
0 26174 7 1 2 26171 26173
0 26175 5 1 1 26174
0 26176 7 1 2 60888 58826
0 26177 7 1 2 26175 26176
0 26178 5 1 1 26177
0 26179 7 1 2 52155 76902
0 26180 7 1 2 76907 26179
0 26181 5 1 1 26180
0 26182 7 2 2 60542 76812
0 26183 7 1 2 76908 76891
0 26184 5 1 1 26183
0 26185 7 1 2 26181 26184
0 26186 5 1 1 26185
0 26187 7 1 2 47932 26186
0 26188 5 1 1 26187
0 26189 7 7 2 49340 53201
0 26190 7 1 2 62636 76910
0 26191 7 1 2 76905 26190
0 26192 5 1 1 26191
0 26193 7 1 2 26188 26192
0 26194 7 1 2 26178 26193
0 26195 7 1 2 26169 26194
0 26196 5 1 1 26195
0 26197 7 1 2 50103 26196
0 26198 5 1 1 26197
0 26199 7 1 2 60944 65006
0 26200 7 1 2 76713 26199
0 26201 5 1 1 26200
0 26202 7 2 2 65153 74840
0 26203 5 1 1 76917
0 26204 7 1 2 48196 26203
0 26205 5 1 1 26204
0 26206 7 1 2 52156 60984
0 26207 5 2 1 26206
0 26208 7 1 2 75775 76919
0 26209 7 1 2 26205 26208
0 26210 5 1 1 26209
0 26211 7 1 2 26201 26210
0 26212 5 1 1 26211
0 26213 7 1 2 64301 72686
0 26214 7 1 2 26212 26213
0 26215 5 1 1 26214
0 26216 7 1 2 26198 26215
0 26217 7 1 2 26124 26216
0 26218 7 1 2 26093 26217
0 26219 5 1 1 26218
0 26220 7 1 2 50222 26219
0 26221 5 1 1 26220
0 26222 7 1 2 65786 76814
0 26223 5 1 1 26222
0 26224 7 1 2 48197 26223
0 26225 5 1 1 26224
0 26226 7 1 2 6184 26225
0 26227 5 1 1 26226
0 26228 7 1 2 76807 26227
0 26229 5 1 1 26228
0 26230 7 1 2 47933 62048
0 26231 5 1 1 26230
0 26232 7 2 2 51946 61184
0 26233 5 4 1 76921
0 26234 7 1 2 53101 68104
0 26235 7 1 2 76923 26234
0 26236 7 1 2 26231 26235
0 26237 5 1 1 26236
0 26238 7 1 2 76870 26237
0 26239 5 1 1 26238
0 26240 7 1 2 52990 26239
0 26241 5 1 1 26240
0 26242 7 1 2 62056 76800
0 26243 5 1 1 26242
0 26244 7 1 2 52294 61595
0 26245 7 1 2 61636 26244
0 26246 7 1 2 26243 26245
0 26247 5 1 1 26246
0 26248 7 1 2 26241 26247
0 26249 5 1 1 26248
0 26250 7 1 2 49452 26249
0 26251 5 1 1 26250
0 26252 7 1 2 26229 26251
0 26253 5 1 1 26252
0 26254 7 1 2 50769 26253
0 26255 5 1 1 26254
0 26256 7 1 2 58434 57172
0 26257 5 1 1 26256
0 26258 7 1 2 58400 60359
0 26259 5 1 1 26258
0 26260 7 1 2 57232 62072
0 26261 5 1 1 26260
0 26262 7 1 2 26259 26261
0 26263 5 1 1 26262
0 26264 7 1 2 56742 26263
0 26265 5 1 1 26264
0 26266 7 1 2 26257 26265
0 26267 5 1 1 26266
0 26268 7 5 2 52295 54674
0 26269 7 1 2 70769 76927
0 26270 7 1 2 26267 26269
0 26271 5 1 1 26270
0 26272 7 1 2 50462 26271
0 26273 7 1 2 26255 26272
0 26274 5 1 1 26273
0 26275 7 1 2 49341 76808
0 26276 7 1 2 70903 26275
0 26277 5 1 1 26276
0 26278 7 1 2 49216 62091
0 26279 5 1 1 26278
0 26280 7 1 2 58562 62041
0 26281 7 1 2 76854 26280
0 26282 7 1 2 26279 26281
0 26283 5 1 1 26282
0 26284 7 1 2 26277 26283
0 26285 5 1 1 26284
0 26286 7 1 2 50770 26285
0 26287 5 1 1 26286
0 26288 7 1 2 53910 58819
0 26289 7 1 2 76349 26288
0 26290 7 1 2 58900 26289
0 26291 5 1 1 26290
0 26292 7 1 2 54323 26291
0 26293 7 1 2 26287 26292
0 26294 5 1 1 26293
0 26295 7 1 2 54043 26294
0 26296 7 1 2 26274 26295
0 26297 5 1 1 26296
0 26298 7 2 2 56113 57622
0 26299 7 1 2 56743 61609
0 26300 5 2 1 26299
0 26301 7 3 2 49453 60543
0 26302 7 1 2 76934 76936
0 26303 5 1 1 26302
0 26304 7 1 2 59376 76138
0 26305 5 1 1 26304
0 26306 7 2 2 51947 59862
0 26307 5 1 1 76939
0 26308 7 1 2 667 26307
0 26309 5 1 1 26308
0 26310 7 1 2 52157 62637
0 26311 7 1 2 26309 26310
0 26312 5 1 1 26311
0 26313 7 1 2 26305 26312
0 26314 5 1 1 26313
0 26315 7 1 2 53202 26314
0 26316 5 1 1 26315
0 26317 7 1 2 26303 26316
0 26318 5 1 1 26317
0 26319 7 1 2 54044 26318
0 26320 5 1 1 26319
0 26321 7 2 2 53203 59377
0 26322 5 2 1 76941
0 26323 7 1 2 61479 76942
0 26324 5 1 1 26323
0 26325 7 1 2 26320 26324
0 26326 5 1 1 26325
0 26327 7 1 2 76932 26326
0 26328 5 1 1 26327
0 26329 7 1 2 70215 68867
0 26330 5 1 1 26329
0 26331 7 1 2 76665 26330
0 26332 5 1 1 26331
0 26333 7 2 2 49217 76659
0 26334 5 1 1 76945
0 26335 7 1 2 59548 76946
0 26336 5 1 1 26335
0 26337 7 1 2 26332 26336
0 26338 5 1 1 26337
0 26339 7 1 2 48388 62358
0 26340 7 1 2 26338 26339
0 26341 5 1 1 26340
0 26342 7 1 2 52419 26341
0 26343 7 1 2 26328 26342
0 26344 7 1 2 26297 26343
0 26345 7 1 2 26221 26344
0 26346 5 1 1 26345
0 26347 7 1 2 48389 50223
0 26348 5 2 1 26347
0 26349 7 1 2 61953 70726
0 26350 5 1 1 26349
0 26351 7 1 2 76947 26350
0 26352 5 1 1 26351
0 26353 7 1 2 55767 26352
0 26354 5 1 1 26353
0 26355 7 1 2 50224 76876
0 26356 5 1 1 26355
0 26357 7 1 2 47934 52158
0 26358 5 1 1 26357
0 26359 7 1 2 54045 60606
0 26360 7 1 2 26358 26359
0 26361 7 1 2 61679 26360
0 26362 5 1 1 26361
0 26363 7 1 2 26356 26362
0 26364 7 1 2 26354 26363
0 26365 5 1 1 26364
0 26366 7 1 2 53204 26365
0 26367 5 1 1 26366
0 26368 7 4 2 49454 50225
0 26369 7 1 2 59780 76949
0 26370 5 1 1 26369
0 26371 7 1 2 53205 65822
0 26372 5 1 1 26371
0 26373 7 1 2 26370 26372
0 26374 5 1 1 26373
0 26375 7 1 2 52296 26374
0 26376 5 1 1 26375
0 26377 7 3 2 52898 76714
0 26378 7 2 2 60474 76953
0 26379 5 1 1 76956
0 26380 7 4 2 53206 54046
0 26381 7 1 2 48390 76958
0 26382 5 1 1 26381
0 26383 7 1 2 26379 26382
0 26384 5 1 1 26383
0 26385 7 1 2 51948 26384
0 26386 5 1 1 26385
0 26387 7 1 2 70881 76950
0 26388 5 1 1 26387
0 26389 7 1 2 54047 76236
0 26390 7 1 2 65935 26389
0 26391 5 1 1 26390
0 26392 7 1 2 26388 26391
0 26393 7 1 2 26386 26392
0 26394 5 1 1 26393
0 26395 7 1 2 52159 26394
0 26396 5 1 1 26395
0 26397 7 1 2 26376 26396
0 26398 7 1 2 26367 26397
0 26399 5 1 1 26398
0 26400 7 1 2 53102 26399
0 26401 5 1 1 26400
0 26402 7 1 2 61820 76924
0 26403 5 1 1 26402
0 26404 7 1 2 52297 60301
0 26405 7 1 2 26403 26404
0 26406 5 1 1 26405
0 26407 7 1 2 52160 76874
0 26408 5 1 1 26407
0 26409 7 1 2 47935 55693
0 26410 5 1 1 26409
0 26411 7 1 2 26408 26410
0 26412 5 1 1 26411
0 26413 7 1 2 61528 26412
0 26414 5 1 1 26413
0 26415 7 3 2 49218 50226
0 26416 7 1 2 62098 76962
0 26417 5 1 1 26416
0 26418 7 1 2 54048 60475
0 26419 5 1 1 26418
0 26420 7 1 2 26417 26419
0 26421 5 1 1 26420
0 26422 7 1 2 60945 26421
0 26423 5 1 1 26422
0 26424 7 1 2 26414 26423
0 26425 7 1 2 26406 26424
0 26426 5 1 1 26425
0 26427 7 1 2 76911 26426
0 26428 5 1 1 26427
0 26429 7 1 2 26401 26428
0 26430 5 1 1 26429
0 26431 7 1 2 50463 26430
0 26432 5 1 1 26431
0 26433 7 5 2 53103 60681
0 26434 5 2 1 76965
0 26435 7 1 2 49219 76966
0 26436 5 1 1 26435
0 26437 7 1 2 49342 60695
0 26438 5 3 1 26437
0 26439 7 3 2 52899 76972
0 26440 7 1 2 59751 61045
0 26441 7 1 2 76975 26440
0 26442 5 1 1 26441
0 26443 7 1 2 26436 26442
0 26444 5 1 1 26443
0 26445 7 1 2 52298 26444
0 26446 5 1 1 26445
0 26447 7 1 2 48391 76940
0 26448 5 1 1 26447
0 26449 7 3 2 52299 54049
0 26450 5 1 1 76978
0 26451 7 1 2 26152 26450
0 26452 7 1 2 26448 26451
0 26453 5 1 1 26452
0 26454 7 1 2 54050 70883
0 26455 5 1 1 26454
0 26456 7 1 2 53104 26455
0 26457 7 1 2 26453 26456
0 26458 5 1 1 26457
0 26459 7 1 2 51949 76897
0 26460 7 1 2 70796 26459
0 26461 5 1 1 26460
0 26462 7 1 2 26458 26461
0 26463 5 1 1 26462
0 26464 7 1 2 52161 26463
0 26465 5 1 1 26464
0 26466 7 1 2 26446 26465
0 26467 5 1 1 26466
0 26468 7 1 2 75776 26467
0 26469 5 1 1 26468
0 26470 7 1 2 26432 26469
0 26471 5 1 1 26470
0 26472 7 1 2 50771 26471
0 26473 5 1 1 26472
0 26474 7 1 2 52991 72840
0 26475 5 1 1 26474
0 26476 7 1 2 17575 26475
0 26477 5 1 1 26476
0 26478 7 1 2 61628 26477
0 26479 5 1 1 26478
0 26480 7 1 2 71968 76829
0 26481 5 1 1 26480
0 26482 7 1 2 26479 26481
0 26483 5 1 1 26482
0 26484 7 1 2 73412 26483
0 26485 5 1 1 26484
0 26486 7 1 2 73754 76819
0 26487 5 1 1 26486
0 26488 7 1 2 26485 26487
0 26489 5 1 1 26488
0 26490 7 1 2 62427 26489
0 26491 5 1 1 26490
0 26492 7 1 2 48198 53207
0 26493 7 1 2 59937 26492
0 26494 7 1 2 76909 26493
0 26495 5 1 1 26494
0 26496 7 1 2 26491 26495
0 26497 5 1 1 26496
0 26498 7 1 2 58435 26497
0 26499 5 1 1 26498
0 26500 7 2 2 52900 76643
0 26501 7 1 2 70998 72841
0 26502 7 1 2 76981 26501
0 26503 5 1 1 26502
0 26504 7 1 2 48508 26503
0 26505 7 1 2 26499 26504
0 26506 7 1 2 26473 26505
0 26507 5 1 1 26506
0 26508 7 1 2 55034 26507
0 26509 7 1 2 26346 26508
0 26510 5 1 1 26509
0 26511 7 2 2 74003 76694
0 26512 5 1 1 76983
0 26513 7 1 2 49455 70639
0 26514 5 1 1 26513
0 26515 7 2 2 53208 61755
0 26516 5 1 1 76985
0 26517 7 1 2 49343 76986
0 26518 5 1 1 26517
0 26519 7 1 2 26514 26518
0 26520 5 1 1 26519
0 26521 7 1 2 48509 26520
0 26522 5 1 1 26521
0 26523 7 1 2 26512 26522
0 26524 5 1 1 26523
0 26525 7 1 2 51950 26524
0 26526 5 1 1 26525
0 26527 7 1 2 712 63126
0 26528 5 1 1 26527
0 26529 7 1 2 48510 76951
0 26530 7 1 2 26528 26529
0 26531 5 1 1 26530
0 26532 7 1 2 26526 26531
0 26533 5 1 1 26532
0 26534 7 1 2 54324 26533
0 26535 5 1 1 26534
0 26536 7 1 2 59993 70361
0 26537 5 1 1 26536
0 26538 7 1 2 56922 76660
0 26539 7 1 2 26537 26538
0 26540 5 1 1 26539
0 26541 7 1 2 26535 26540
0 26542 5 1 1 26541
0 26543 7 1 2 58436 26542
0 26544 5 1 1 26543
0 26545 7 1 2 66570 71028
0 26546 5 1 1 26545
0 26547 7 1 2 48392 65178
0 26548 5 1 1 26547
0 26549 7 1 2 26546 26548
0 26550 5 1 1 26549
0 26551 7 1 2 76912 26550
0 26552 5 1 1 26551
0 26553 7 1 2 56744 66588
0 26554 5 1 1 26553
0 26555 7 1 2 62436 76666
0 26556 5 1 1 26555
0 26557 7 1 2 52992 59618
0 26558 5 2 1 26557
0 26559 7 1 2 17952 76987
0 26560 7 1 2 26556 26559
0 26561 5 1 1 26560
0 26562 7 1 2 62728 26561
0 26563 5 1 1 26562
0 26564 7 1 2 26554 26563
0 26565 5 1 1 26564
0 26566 7 1 2 55768 26565
0 26567 5 2 1 26566
0 26568 7 1 2 63187 73961
0 26569 5 2 1 26568
0 26570 7 1 2 58401 76991
0 26571 5 1 1 26570
0 26572 7 1 2 26334 26571
0 26573 5 1 1 26572
0 26574 7 1 2 48199 26573
0 26575 5 1 1 26574
0 26576 7 1 2 76988 26575
0 26577 5 1 1 26576
0 26578 7 1 2 48393 26577
0 26579 5 1 1 26578
0 26580 7 1 2 56114 70234
0 26581 7 1 2 74004 26580
0 26582 5 1 1 26581
0 26583 7 1 2 63197 26582
0 26584 5 1 1 26583
0 26585 7 1 2 62057 26584
0 26586 5 1 1 26585
0 26587 7 1 2 52300 65405
0 26588 5 4 1 26587
0 26589 7 1 2 49344 63181
0 26590 5 1 1 26589
0 26591 7 1 2 49220 59641
0 26592 7 1 2 65751 26591
0 26593 5 1 1 26592
0 26594 7 1 2 26590 26593
0 26595 5 1 1 26594
0 26596 7 1 2 76993 26595
0 26597 5 1 1 26596
0 26598 7 2 2 26586 26597
0 26599 7 1 2 65757 76903
0 26600 5 1 1 26599
0 26601 7 1 2 76997 26600
0 26602 7 1 2 26579 26601
0 26603 7 1 2 76989 26602
0 26604 5 1 1 26603
0 26605 7 1 2 49456 26604
0 26606 5 1 1 26605
0 26607 7 1 2 26552 26606
0 26608 5 1 1 26607
0 26609 7 1 2 52420 26608
0 26610 5 1 1 26609
0 26611 7 1 2 62092 62611
0 26612 5 1 1 26611
0 26613 7 1 2 54325 62235
0 26614 5 1 1 26613
0 26615 7 1 2 26612 26614
0 26616 5 1 1 26615
0 26617 7 1 2 53105 26616
0 26618 5 1 1 26617
0 26619 7 1 2 49345 60204
0 26620 5 2 1 26619
0 26621 7 3 2 52162 72692
0 26622 7 1 2 50104 54326
0 26623 7 1 2 77001 26622
0 26624 5 1 1 26623
0 26625 7 1 2 76999 26624
0 26626 7 1 2 26618 26625
0 26627 5 1 1 26626
0 26628 7 1 2 52993 26627
0 26629 5 1 1 26628
0 26630 7 1 2 50227 76051
0 26631 5 1 1 26630
0 26632 7 1 2 49221 76979
0 26633 5 1 1 26632
0 26634 7 1 2 26631 26633
0 26635 5 1 1 26634
0 26636 7 1 2 59659 26635
0 26637 5 1 1 26636
0 26638 7 1 2 48394 70754
0 26639 5 1 1 26638
0 26640 7 1 2 51951 26639
0 26641 5 2 1 26640
0 26642 7 1 2 261 77004
0 26643 5 3 1 26642
0 26644 7 1 2 76827 77006
0 26645 5 1 1 26644
0 26646 7 1 2 52301 76663
0 26647 5 1 1 26646
0 26648 7 1 2 61773 59692
0 26649 7 1 2 26647 26648
0 26650 5 1 1 26649
0 26651 7 1 2 49457 26650
0 26652 7 1 2 26645 26651
0 26653 7 1 2 26637 26652
0 26654 7 1 2 26629 26653
0 26655 5 1 1 26654
0 26656 7 1 2 60396 76898
0 26657 5 1 1 26656
0 26658 7 1 2 53106 61730
0 26659 5 2 1 26658
0 26660 7 1 2 48395 62865
0 26661 7 1 2 77009 26660
0 26662 5 1 1 26661
0 26663 7 1 2 26657 26662
0 26664 5 1 1 26663
0 26665 7 1 2 49222 26664
0 26666 5 1 1 26665
0 26667 7 1 2 50228 65403
0 26668 5 1 1 26667
0 26669 7 1 2 25826 26668
0 26670 5 1 1 26669
0 26671 7 1 2 58171 26670
0 26672 5 1 1 26671
0 26673 7 1 2 53209 26672
0 26674 7 1 2 26666 26673
0 26675 7 1 2 76998 26674
0 26676 7 1 2 76990 26675
0 26677 5 1 1 26676
0 26678 7 1 2 48511 26677
0 26679 7 1 2 26655 26678
0 26680 5 1 1 26679
0 26681 7 1 2 54327 61452
0 26682 5 1 1 26681
0 26683 7 1 2 70727 76661
0 26684 5 1 1 26683
0 26685 7 1 2 49458 26684
0 26686 7 1 2 26682 26685
0 26687 5 1 1 26686
0 26688 7 1 2 53210 62792
0 26689 5 2 1 26688
0 26690 7 1 2 48512 66356
0 26691 7 1 2 77011 26690
0 26692 7 1 2 26687 26691
0 26693 5 1 1 26692
0 26694 7 1 2 54328 76984
0 26695 5 1 1 26694
0 26696 7 1 2 26693 26695
0 26697 5 1 1 26696
0 26698 7 1 2 61185 26697
0 26699 5 1 1 26698
0 26700 7 2 2 60205 61390
0 26701 5 1 1 77013
0 26702 7 1 2 67390 76880
0 26703 7 1 2 77014 26702
0 26704 5 1 1 26703
0 26705 7 1 2 54675 26704
0 26706 7 1 2 26699 26705
0 26707 7 1 2 26680 26706
0 26708 7 1 2 26610 26707
0 26709 7 1 2 26544 26708
0 26710 5 1 1 26709
0 26711 7 1 2 53911 62804
0 26712 5 1 1 26711
0 26713 7 1 2 62812 26712
0 26714 5 1 1 26713
0 26715 7 1 2 58865 26714
0 26716 5 1 1 26715
0 26717 7 2 2 54329 62805
0 26718 5 1 1 77015
0 26719 7 1 2 58271 58838
0 26720 5 1 1 26719
0 26721 7 1 2 73944 26720
0 26722 5 2 1 26721
0 26723 7 1 2 74157 74703
0 26724 5 1 1 26723
0 26725 7 1 2 77017 26724
0 26726 5 1 1 26725
0 26727 7 1 2 56115 26726
0 26728 5 1 1 26727
0 26729 7 1 2 26718 26728
0 26730 7 1 2 26716 26729
0 26731 5 1 1 26730
0 26732 7 1 2 49459 26731
0 26733 5 1 1 26732
0 26734 7 2 2 48396 76850
0 26735 7 1 2 74791 77019
0 26736 5 1 1 26735
0 26737 7 1 2 26733 26736
0 26738 5 1 1 26737
0 26739 7 1 2 48513 26738
0 26740 5 1 1 26739
0 26741 7 2 2 47936 61840
0 26742 5 1 1 77021
0 26743 7 1 2 49124 77022
0 26744 5 1 1 26743
0 26745 7 1 2 67304 26744
0 26746 5 3 1 26745
0 26747 7 1 2 53912 64894
0 26748 5 1 1 26747
0 26749 7 1 2 66646 26748
0 26750 5 1 1 26749
0 26751 7 1 2 77023 26750
0 26752 5 1 1 26751
0 26753 7 2 2 65912 76851
0 26754 5 1 1 77026
0 26755 7 1 2 64883 77027
0 26756 5 1 1 26755
0 26757 7 1 2 50772 26756
0 26758 7 1 2 26752 26757
0 26759 7 1 2 26740 26758
0 26760 5 1 1 26759
0 26761 7 1 2 51057 26760
0 26762 7 1 2 26710 26761
0 26763 5 1 1 26762
0 26764 7 1 2 53329 26763
0 26765 7 1 2 26510 26764
0 26766 5 1 1 26765
0 26767 7 1 2 51058 76771
0 26768 5 1 1 26767
0 26769 7 1 2 51059 76834
0 26770 5 1 1 26769
0 26771 7 1 2 25983 26770
0 26772 5 1 1 26771
0 26773 7 1 2 58437 26772
0 26774 5 1 1 26773
0 26775 7 1 2 76846 76866
0 26776 5 1 1 26775
0 26777 7 1 2 49574 26776
0 26778 7 1 2 26774 26777
0 26779 7 1 2 26768 26778
0 26780 7 1 2 51060 76788
0 26781 5 1 1 26780
0 26782 7 1 2 65222 73413
0 26783 7 1 2 73780 70891
0 26784 7 1 2 26782 26783
0 26785 5 1 1 26784
0 26786 7 1 2 26781 26785
0 26787 5 1 1 26786
0 26788 7 1 2 76779 26787
0 26789 5 1 1 26788
0 26790 7 1 2 51061 76823
0 26791 5 1 1 26790
0 26792 7 1 2 26789 26791
0 26793 5 1 1 26792
0 26794 7 1 2 50464 26793
0 26795 5 1 1 26794
0 26796 7 1 2 51062 76716
0 26797 5 1 1 26796
0 26798 7 1 2 25995 26797
0 26799 5 1 1 26798
0 26800 7 1 2 57233 26799
0 26801 5 1 1 26800
0 26802 7 1 2 26795 26801
0 26803 7 1 2 26779 26802
0 26804 5 1 1 26803
0 26805 7 1 2 52519 26804
0 26806 7 1 2 26766 26805
0 26807 5 1 1 26806
0 26808 7 1 2 63641 75756
0 26809 5 1 1 26808
0 26810 7 2 2 52901 65007
0 26811 5 1 1 77028
0 26812 7 2 2 56116 26811
0 26813 5 1 1 77030
0 26814 7 1 2 51952 26813
0 26815 5 1 1 26814
0 26816 7 1 2 54330 13571
0 26817 5 2 1 26816
0 26818 7 1 2 52302 77032
0 26819 5 1 1 26818
0 26820 7 1 2 26815 26819
0 26821 5 1 1 26820
0 26822 7 1 2 59683 26821
0 26823 5 1 1 26822
0 26824 7 1 2 74308 76881
0 26825 5 1 1 26824
0 26826 7 1 2 26823 26825
0 26827 5 1 1 26826
0 26828 7 1 2 26827 75381
0 26829 5 1 1 26828
0 26830 7 1 2 26809 26829
0 26831 5 1 1 26830
0 26832 7 1 2 76707 26831
0 26833 5 1 1 26832
0 26834 7 1 2 64530 72974
0 26835 7 1 2 60521 26834
0 26836 5 1 1 26835
0 26837 7 1 2 26833 26836
0 26838 5 1 1 26837
0 26839 7 1 2 50773 26838
0 26840 5 1 1 26839
0 26841 7 1 2 50465 76855
0 26842 7 1 2 76933 26841
0 26843 5 1 1 26842
0 26844 7 1 2 60946 58866
0 26845 7 1 2 75473 26844
0 26846 5 1 1 26845
0 26847 7 1 2 26843 26846
0 26848 5 1 1 26847
0 26849 7 1 2 63457 70169
0 26850 7 1 2 26848 26849
0 26851 5 1 1 26850
0 26852 7 1 2 26840 26851
0 26853 5 1 1 26852
0 26854 7 1 2 61561 76847
0 26855 7 1 2 26853 26854
0 26856 5 1 1 26855
0 26857 7 1 2 55364 26856
0 26858 7 1 2 26807 26857
0 26859 7 1 2 26041 26858
0 26860 5 1 1 26859
0 26861 7 2 2 61029 58502
0 26862 5 1 1 77034
0 26863 7 1 2 54051 60076
0 26864 5 1 1 26863
0 26865 7 1 2 61288 26864
0 26866 5 1 1 26865
0 26867 7 1 2 77035 26866
0 26868 5 1 1 26867
0 26869 7 1 2 60724 64055
0 26870 5 4 1 26869
0 26871 7 1 2 49346 77036
0 26872 5 1 1 26871
0 26873 7 1 2 47937 74768
0 26874 5 1 1 26873
0 26875 7 1 2 49347 60717
0 26876 5 2 1 26875
0 26877 7 1 2 26874 77040
0 26878 5 1 1 26877
0 26879 7 1 2 48397 26878
0 26880 5 1 1 26879
0 26881 7 1 2 26872 26880
0 26882 5 1 1 26881
0 26883 7 1 2 57173 26882
0 26884 5 1 1 26883
0 26885 7 1 2 48514 71021
0 26886 7 1 2 9707 26885
0 26887 5 1 1 26886
0 26888 7 1 2 50774 26887
0 26889 7 1 2 26884 26888
0 26890 7 1 2 26868 26889
0 26891 5 1 1 26890
0 26892 7 1 2 62408 8919
0 26893 5 1 1 26892
0 26894 7 1 2 59173 59729
0 26895 7 1 2 26893 26894
0 26896 5 1 1 26895
0 26897 7 1 2 50466 26896
0 26898 5 1 1 26897
0 26899 7 2 2 63253 55769
0 26900 5 2 1 77042
0 26901 7 1 2 64307 77043
0 26902 5 1 1 26901
0 26903 7 1 2 59619 26902
0 26904 5 1 1 26903
0 26905 7 1 2 58259 76963
0 26906 5 2 1 26905
0 26907 7 1 2 54676 77046
0 26908 7 1 2 26862 26907
0 26909 7 1 2 26904 26908
0 26910 7 1 2 26898 26909
0 26911 5 1 1 26910
0 26912 7 1 2 26891 26911
0 26913 5 1 1 26912
0 26914 7 1 2 48515 66252
0 26915 5 2 1 26914
0 26916 7 1 2 74965 77048
0 26917 5 2 1 26916
0 26918 7 1 2 47938 77050
0 26919 5 1 1 26918
0 26920 7 1 2 50467 64004
0 26921 5 1 1 26920
0 26922 7 1 2 63967 66253
0 26923 5 1 1 26922
0 26924 7 1 2 26921 26923
0 26925 7 1 2 26919 26924
0 26926 5 1 1 26925
0 26927 7 1 2 61977 26926
0 26928 5 1 1 26927
0 26929 7 2 2 47939 62638
0 26930 5 1 1 77052
0 26931 7 1 2 59174 65880
0 26932 5 1 1 26931
0 26933 7 1 2 50775 26932
0 26934 5 1 1 26933
0 26935 7 1 2 26930 26934
0 26936 5 1 1 26935
0 26937 7 1 2 54052 26936
0 26938 5 1 1 26937
0 26939 7 1 2 74966 26938
0 26940 5 1 1 26939
0 26941 7 1 2 55770 26940
0 26942 5 1 1 26941
0 26943 7 1 2 54053 62639
0 26944 5 2 1 26943
0 26945 7 1 2 61398 65803
0 26946 5 1 1 26945
0 26947 7 1 2 50776 63921
0 26948 7 1 2 26946 26947
0 26949 5 1 1 26948
0 26950 7 1 2 77054 26949
0 26951 5 1 1 26950
0 26952 7 1 2 58402 26951
0 26953 5 1 1 26952
0 26954 7 1 2 26942 26953
0 26955 5 1 1 26954
0 26956 7 1 2 56745 26955
0 26957 5 1 1 26956
0 26958 7 1 2 26928 26957
0 26959 7 1 2 26913 26958
0 26960 5 1 1 26959
0 26961 7 1 2 49460 26960
0 26962 5 1 1 26961
0 26963 7 3 2 48516 58719
0 26964 7 1 2 57756 74475
0 26965 5 2 1 26964
0 26966 7 1 2 77056 77059
0 26967 5 1 1 26966
0 26968 7 1 2 61859 76351
0 26969 5 1 1 26968
0 26970 7 1 2 26967 26969
0 26971 5 1 1 26970
0 26972 7 1 2 55771 26971
0 26973 5 1 1 26972
0 26974 7 1 2 60961 66254
0 26975 5 1 1 26974
0 26976 7 1 2 50468 65950
0 26977 5 2 1 26976
0 26978 7 1 2 26975 77061
0 26979 5 1 1 26978
0 26980 7 1 2 48517 26979
0 26981 5 1 1 26980
0 26982 7 1 2 26973 26981
0 26983 7 1 2 53211 61908
0 26984 5 2 1 26983
0 26985 7 1 2 4975 77063
0 26986 5 1 1 26985
0 26987 7 1 2 47940 26986
0 26988 5 1 1 26987
0 26989 7 1 2 77049 26988
0 26990 5 1 1 26989
0 26991 7 1 2 58260 26990
0 26992 5 1 1 26991
0 26993 7 1 2 50469 63347
0 26994 5 1 1 26993
0 26995 7 1 2 26992 26994
0 26996 5 1 1 26995
0 26997 7 1 2 58607 26996
0 26998 5 1 1 26997
0 26999 7 1 2 47941 60302
0 27000 7 1 2 62197 26999
0 27001 7 1 2 58287 27000
0 27002 5 2 1 27001
0 27003 7 1 2 76691 77065
0 27004 5 1 1 27003
0 27005 7 1 2 54677 27004
0 27006 5 1 1 27005
0 27007 7 3 2 48518 59994
0 27008 5 1 1 77067
0 27009 7 1 2 59436 59392
0 27010 7 1 2 77068 27009
0 27011 5 1 1 27010
0 27012 7 1 2 27006 27011
0 27013 5 1 1 27012
0 27014 7 1 2 54331 27013
0 27015 5 1 1 27014
0 27016 7 1 2 26998 27015
0 27017 7 1 2 26982 27016
0 27018 5 1 1 27017
0 27019 7 1 2 56117 27018
0 27020 5 1 1 27019
0 27021 7 1 2 47942 62612
0 27022 5 1 1 27021
0 27023 7 1 2 63188 27022
0 27024 5 2 1 27023
0 27025 7 1 2 56746 77070
0 27026 5 1 1 27025
0 27027 7 1 2 50470 61480
0 27028 5 1 1 27027
0 27029 7 1 2 27026 27028
0 27030 5 1 1 27029
0 27031 7 1 2 55772 27030
0 27032 5 1 1 27031
0 27033 7 1 2 50471 74785
0 27034 5 1 1 27033
0 27035 7 1 2 63182 76046
0 27036 5 1 1 27035
0 27037 7 1 2 27034 27036
0 27038 7 1 2 27032 27037
0 27039 5 1 1 27038
0 27040 7 1 2 63348 27039
0 27041 5 1 1 27040
0 27042 7 1 2 74309 74849
0 27043 5 1 1 27042
0 27044 7 1 2 57174 66690
0 27045 5 1 1 27044
0 27046 7 1 2 27043 27045
0 27047 5 1 1 27046
0 27048 7 1 2 55773 27047
0 27049 5 1 1 27048
0 27050 7 1 2 50777 58508
0 27051 5 1 1 27050
0 27052 7 1 2 77055 27051
0 27053 5 1 1 27052
0 27054 7 1 2 74583 27053
0 27055 5 1 1 27054
0 27056 7 1 2 76052 77051
0 27057 5 1 1 27056
0 27058 7 1 2 59720 62640
0 27059 5 1 1 27058
0 27060 7 1 2 65869 77057
0 27061 5 1 1 27060
0 27062 7 1 2 27059 27061
0 27063 7 1 2 27057 27062
0 27064 7 1 2 27055 27063
0 27065 7 1 2 27049 27064
0 27066 5 1 1 27065
0 27067 7 1 2 57503 27066
0 27068 5 1 1 27067
0 27069 7 1 2 27041 27068
0 27070 7 1 2 27020 27069
0 27071 7 1 2 26962 27070
0 27072 5 1 1 27071
0 27073 7 1 2 49575 27072
0 27074 5 1 1 27073
0 27075 7 1 2 50229 59449
0 27076 5 2 1 27075
0 27077 7 1 2 64989 74535
0 27078 7 2 2 77072 27077
0 27079 5 1 1 77074
0 27080 7 1 2 20983 27079
0 27081 5 1 1 27080
0 27082 7 2 2 56118 27081
0 27083 7 1 2 71848 77076
0 27084 5 1 1 27083
0 27085 7 3 2 50230 57504
0 27086 5 2 1 77078
0 27087 7 1 2 62238 77079
0 27088 5 2 1 27087
0 27089 7 1 2 27084 77083
0 27090 5 1 1 27089
0 27091 7 1 2 54332 27090
0 27092 5 1 1 27091
0 27093 7 1 2 50472 65392
0 27094 7 1 2 62158 27093
0 27095 5 2 1 27094
0 27096 7 1 2 27092 77085
0 27097 5 1 1 27096
0 27098 7 1 2 49223 27097
0 27099 5 1 1 27098
0 27100 7 1 2 53330 75592
0 27101 5 1 1 27100
0 27102 7 1 2 77081 27101
0 27103 5 1 1 27102
0 27104 7 1 2 57828 27103
0 27105 5 1 1 27104
0 27106 7 1 2 62866 72536
0 27107 5 2 1 27106
0 27108 7 1 2 27105 77087
0 27109 5 1 1 27108
0 27110 7 1 2 58608 27109
0 27111 5 1 1 27110
0 27112 7 2 2 47943 50231
0 27113 5 1 1 77089
0 27114 7 1 2 55694 27113
0 27115 5 1 1 27114
0 27116 7 1 2 71801 27115
0 27117 7 1 2 77071 27116
0 27118 5 2 1 27117
0 27119 7 1 2 27111 77091
0 27120 7 1 2 27099 27119
0 27121 5 1 1 27120
0 27122 7 1 2 65073 27121
0 27123 5 1 1 27122
0 27124 7 1 2 27074 27123
0 27125 5 1 1 27124
0 27126 7 1 2 48618 27125
0 27127 5 1 1 27126
0 27128 7 1 2 53212 61924
0 27129 5 2 1 27128
0 27130 7 2 2 59183 77093
0 27131 7 1 2 62143 77095
0 27132 5 1 1 27131
0 27133 7 1 2 50778 61949
0 27134 5 1 1 27133
0 27135 7 1 2 62195 70470
0 27136 5 1 1 27135
0 27137 7 1 2 27134 27136
0 27138 7 1 2 27132 27137
0 27139 5 1 1 27138
0 27140 7 1 2 54333 27139
0 27141 5 1 1 27140
0 27142 7 1 2 50779 66640
0 27143 5 1 1 27142
0 27144 7 1 2 27141 27143
0 27145 5 1 1 27144
0 27146 7 1 2 49576 27145
0 27147 5 1 1 27146
0 27148 7 1 2 65122 75705
0 27149 5 1 1 27148
0 27150 7 1 2 27147 27149
0 27151 5 1 1 27150
0 27152 7 1 2 48619 27151
0 27153 5 1 1 27152
0 27154 7 1 2 71956 75645
0 27155 5 1 1 27154
0 27156 7 1 2 27153 27155
0 27157 5 1 1 27156
0 27158 7 1 2 61261 27157
0 27159 5 1 1 27158
0 27160 7 2 2 56923 64237
0 27161 7 2 2 48620 54054
0 27162 5 1 1 77099
0 27163 7 1 2 77077 27162
0 27164 5 1 1 27163
0 27165 7 1 2 77084 27164
0 27166 5 1 1 27165
0 27167 7 1 2 54334 27166
0 27168 5 1 1 27167
0 27169 7 1 2 77086 27168
0 27170 5 1 1 27169
0 27171 7 1 2 49224 27170
0 27172 5 1 1 27171
0 27173 7 1 2 59080 75737
0 27174 5 1 1 27173
0 27175 7 1 2 77082 27174
0 27176 5 1 1 27175
0 27177 7 1 2 57829 27176
0 27178 5 1 1 27177
0 27179 7 1 2 77088 27178
0 27180 5 1 1 27179
0 27181 7 1 2 58609 27180
0 27182 5 1 1 27181
0 27183 7 1 2 77092 27182
0 27184 7 1 2 27172 27183
0 27185 5 1 1 27184
0 27186 7 1 2 77097 27185
0 27187 5 1 1 27186
0 27188 7 1 2 27159 27187
0 27189 7 1 2 27127 27188
0 27190 5 1 1 27189
0 27191 7 1 2 51063 27190
0 27192 5 1 1 27191
0 27193 7 1 2 59301 66937
0 27194 5 1 1 27193
0 27195 7 1 2 54055 27194
0 27196 5 1 1 27195
0 27197 7 1 2 57791 27196
0 27198 5 1 1 27197
0 27199 7 1 2 55774 27198
0 27200 5 1 1 27199
0 27201 7 1 2 61399 59789
0 27202 5 1 1 27201
0 27203 7 1 2 65208 27202
0 27204 5 1 1 27203
0 27205 7 1 2 59088 70758
0 27206 5 1 1 27205
0 27207 7 1 2 54335 27206
0 27208 5 1 1 27207
0 27209 7 1 2 64953 27208
0 27210 7 1 2 27204 27209
0 27211 7 1 2 27200 27210
0 27212 5 1 1 27211
0 27213 7 1 2 53213 27212
0 27214 5 1 1 27213
0 27215 7 1 2 59462 70368
0 27216 5 1 1 27215
0 27217 7 1 2 49348 27216
0 27218 5 1 1 27217
0 27219 7 1 2 55775 59109
0 27220 5 1 1 27219
0 27221 7 1 2 27218 27220
0 27222 5 1 1 27221
0 27223 7 1 2 60206 27222
0 27224 5 1 1 27223
0 27225 7 1 2 53214 65838
0 27226 5 1 1 27225
0 27227 7 1 2 26701 27226
0 27228 5 1 1 27227
0 27229 7 1 2 58307 27228
0 27230 5 1 1 27229
0 27231 7 3 2 56119 62729
0 27232 5 2 1 77101
0 27233 7 1 2 65412 77104
0 27234 5 1 1 27233
0 27235 7 1 2 53215 27234
0 27236 5 1 1 27235
0 27237 7 1 2 59081 72485
0 27238 5 1 1 27237
0 27239 7 1 2 27236 27238
0 27240 5 1 1 27239
0 27241 7 1 2 58610 27240
0 27242 5 1 1 27241
0 27243 7 2 2 60106 63586
0 27244 5 4 1 77106
0 27245 7 1 2 60207 77107
0 27246 5 1 1 27245
0 27247 7 2 2 48398 62730
0 27248 5 2 1 77112
0 27249 7 1 2 49461 61073
0 27250 7 1 2 77114 27249
0 27251 7 1 2 27246 27250
0 27252 5 1 1 27251
0 27253 7 1 2 27242 27252
0 27254 7 1 2 27230 27253
0 27255 7 1 2 27224 27254
0 27256 7 1 2 27214 27255
0 27257 5 1 1 27256
0 27258 7 1 2 48519 27257
0 27259 5 1 1 27258
0 27260 7 2 2 55776 60749
0 27261 5 1 1 77116
0 27262 7 1 2 59730 27261
0 27263 5 2 1 27262
0 27264 7 1 2 54056 77118
0 27265 5 1 1 27264
0 27266 7 1 2 59411 27265
0 27267 5 1 1 27266
0 27268 7 1 2 47944 27267
0 27269 5 1 1 27268
0 27270 7 1 2 61186 71405
0 27271 5 1 1 27270
0 27272 7 1 2 57772 27271
0 27273 5 1 1 27272
0 27274 7 2 2 27269 27273
0 27275 5 2 1 77120
0 27276 7 1 2 76809 77122
0 27277 5 1 1 27276
0 27278 7 1 2 58172 76959
0 27279 5 1 1 27278
0 27280 7 1 2 49462 60245
0 27281 5 10 1 27280
0 27282 7 1 2 47945 4429
0 27283 7 1 2 66357 27282
0 27284 7 1 2 77124 27283
0 27285 5 1 1 27284
0 27286 7 1 2 27279 27285
0 27287 5 1 1 27286
0 27288 7 1 2 48200 27287
0 27289 5 1 1 27288
0 27290 7 1 2 62731 76695
0 27291 5 1 1 27290
0 27292 7 1 2 27289 27291
0 27293 5 1 1 27292
0 27294 7 1 2 58611 27293
0 27295 5 1 1 27294
0 27296 7 1 2 60985 61187
0 27297 5 1 1 27296
0 27298 7 1 2 49225 27297
0 27299 5 1 1 27298
0 27300 7 1 2 63255 27299
0 27301 5 1 1 27300
0 27302 7 1 2 60208 27301
0 27303 5 1 1 27302
0 27304 7 2 2 48399 60209
0 27305 5 1 1 77134
0 27306 7 1 2 52421 65209
0 27307 5 1 1 27306
0 27308 7 1 2 27305 27307
0 27309 5 1 1 27308
0 27310 7 1 2 59829 27309
0 27311 5 1 1 27310
0 27312 7 1 2 58272 70919
0 27313 7 1 2 74021 27312
0 27314 5 1 1 27313
0 27315 7 1 2 52422 27314
0 27316 5 1 1 27315
0 27317 7 1 2 27311 27316
0 27318 7 1 2 27303 27317
0 27319 5 1 1 27318
0 27320 7 1 2 49463 27319
0 27321 5 1 1 27320
0 27322 7 1 2 27295 27321
0 27323 7 1 2 27277 27322
0 27324 5 1 1 27323
0 27325 7 1 2 49349 27324
0 27326 5 1 1 27325
0 27327 7 2 2 50232 59642
0 27328 5 1 1 77136
0 27329 7 2 2 58328 77137
0 27330 7 1 2 48201 77138
0 27331 5 1 1 27330
0 27332 7 2 2 48400 59660
0 27333 5 1 1 77140
0 27334 7 1 2 54057 77141
0 27335 5 1 1 27334
0 27336 7 1 2 27331 27335
0 27337 5 1 1 27336
0 27338 7 1 2 47946 27337
0 27339 5 1 1 27338
0 27340 7 2 2 54058 75624
0 27341 5 1 1 77142
0 27342 7 1 2 48202 77143
0 27343 5 1 1 27342
0 27344 7 1 2 27339 27343
0 27345 5 1 1 27344
0 27346 7 1 2 58612 27345
0 27347 5 1 1 27346
0 27348 7 1 2 60210 59454
0 27349 5 1 1 27348
0 27350 7 1 2 53107 76878
0 27351 7 1 2 76992 27350
0 27352 5 1 1 27351
0 27353 7 1 2 27349 27352
0 27354 5 1 1 27353
0 27355 7 1 2 48401 27354
0 27356 5 1 1 27355
0 27357 7 1 2 74515 71549
0 27358 5 1 1 27357
0 27359 7 1 2 27341 27358
0 27360 5 1 1 27359
0 27361 7 1 2 52303 58295
0 27362 5 2 1 27361
0 27363 7 1 2 27360 77144
0 27364 5 1 1 27363
0 27365 7 1 2 47947 75625
0 27366 5 1 1 27365
0 27367 7 1 2 27333 27366
0 27368 5 1 1 27367
0 27369 7 1 2 61821 27368
0 27370 5 1 1 27369
0 27371 7 1 2 57283 62437
0 27372 7 1 2 77139 27371
0 27373 5 1 1 27372
0 27374 7 1 2 27370 27373
0 27375 5 1 1 27374
0 27376 7 1 2 55777 27375
0 27377 5 1 1 27376
0 27378 7 1 2 27364 27377
0 27379 7 1 2 27356 27378
0 27380 7 1 2 27347 27379
0 27381 5 1 1 27380
0 27382 7 1 2 49464 27381
0 27383 5 1 1 27382
0 27384 7 1 2 27326 27383
0 27385 7 1 2 27259 27384
0 27386 5 1 1 27385
0 27387 7 1 2 54678 27386
0 27388 5 2 1 27387
0 27389 7 1 2 62350 69879
0 27390 5 1 1 27389
0 27391 7 1 2 57505 61841
0 27392 5 1 1 27391
0 27393 7 1 2 27390 27392
0 27394 5 1 1 27393
0 27395 7 1 2 64872 27394
0 27396 5 1 1 27395
0 27397 7 1 2 59184 70861
0 27398 5 1 1 27397
0 27399 7 2 2 52423 57792
0 27400 5 1 1 77148
0 27401 7 1 2 63224 27400
0 27402 5 1 1 27401
0 27403 7 1 2 27398 27402
0 27404 5 1 1 27403
0 27405 7 1 2 47948 27404
0 27406 5 1 1 27405
0 27407 7 2 2 58517 56747
0 27408 5 1 1 77150
0 27409 7 1 2 27406 27408
0 27410 5 1 1 27409
0 27411 7 1 2 55778 27410
0 27412 5 1 1 27411
0 27413 7 1 2 60341 60037
0 27414 5 3 1 27413
0 27415 7 1 2 48520 77152
0 27416 5 1 1 27415
0 27417 7 1 2 60303 61272
0 27418 5 1 1 27417
0 27419 7 1 2 27416 27418
0 27420 5 1 1 27419
0 27421 7 1 2 58613 27420
0 27422 5 1 1 27421
0 27423 7 1 2 63914 27008
0 27424 5 1 1 27423
0 27425 7 1 2 48203 27424
0 27426 5 1 1 27425
0 27427 7 1 2 64876 27426
0 27428 5 1 1 27427
0 27429 7 1 2 58308 27428
0 27430 5 1 1 27429
0 27431 7 1 2 48204 74814
0 27432 5 1 1 27431
0 27433 7 2 2 58181 27432
0 27434 5 2 1 77155
0 27435 7 1 2 61375 77157
0 27436 5 1 1 27435
0 27437 7 2 2 58518 62447
0 27438 5 1 1 77159
0 27439 7 1 2 27436 27438
0 27440 7 1 2 27430 27439
0 27441 7 1 2 27422 27440
0 27442 7 1 2 27412 27441
0 27443 5 1 1 27442
0 27444 7 1 2 49465 27443
0 27445 5 1 1 27444
0 27446 7 1 2 27396 27445
0 27447 5 1 1 27446
0 27448 7 1 2 50780 27447
0 27449 5 1 1 27448
0 27450 7 1 2 77146 27449
0 27451 5 1 1 27450
0 27452 7 1 2 49577 27451
0 27453 5 1 1 27452
0 27454 7 1 2 55779 69156
0 27455 5 1 1 27454
0 27456 7 1 2 23409 27455
0 27457 5 1 1 27456
0 27458 7 1 2 47949 27457
0 27459 5 1 1 27458
0 27460 7 2 2 71406 74826
0 27461 5 2 1 77161
0 27462 7 1 2 54336 77163
0 27463 5 1 1 27462
0 27464 7 1 2 27459 27463
0 27465 5 1 1 27464
0 27466 7 1 2 48205 27465
0 27467 5 1 1 27466
0 27468 7 1 2 63944 62073
0 27469 5 1 1 27468
0 27470 7 3 2 61943 27469
0 27471 5 5 1 77165
0 27472 7 1 2 57773 77168
0 27473 5 1 1 27472
0 27474 7 1 2 27467 27473
0 27475 5 2 1 27474
0 27476 7 1 2 65123 75436
0 27477 7 1 2 77173 27476
0 27478 5 1 1 27477
0 27479 7 1 2 27453 27478
0 27480 5 1 1 27479
0 27481 7 1 2 52520 27480
0 27482 5 1 1 27481
0 27483 7 2 2 56120 62758
0 27484 5 1 1 77175
0 27485 7 1 2 47950 70862
0 27486 5 1 1 27485
0 27487 7 1 2 27484 27486
0 27488 5 2 1 27487
0 27489 7 1 2 55780 77177
0 27490 5 1 1 27489
0 27491 7 1 2 65417 1064
0 27492 5 1 1 27491
0 27493 7 1 2 59582 27492
0 27494 5 1 1 27493
0 27495 7 1 2 58614 77153
0 27496 5 1 1 27495
0 27497 7 1 2 60421 58487
0 27498 5 1 1 27497
0 27499 7 1 2 48206 27498
0 27500 5 1 1 27499
0 27501 7 1 2 27496 27500
0 27502 7 2 2 27494 27501
0 27503 7 1 2 27490 77179
0 27504 5 1 1 27503
0 27505 7 1 2 56924 27504
0 27506 5 1 1 27505
0 27507 7 2 2 60962 63036
0 27508 5 1 1 77181
0 27509 7 1 2 49350 27508
0 27510 5 1 1 27509
0 27511 7 1 2 49226 67319
0 27512 5 1 1 27511
0 27513 7 1 2 59643 27512
0 27514 5 1 1 27513
0 27515 7 2 2 48207 27514
0 27516 5 1 1 77183
0 27517 7 1 2 49351 70235
0 27518 5 1 1 27517
0 27519 7 1 2 27516 27518
0 27520 5 2 1 27519
0 27521 7 1 2 69880 77185
0 27522 5 1 1 27521
0 27523 7 2 2 27510 27522
0 27524 5 1 1 77187
0 27525 7 1 2 48402 27524
0 27526 5 1 1 27525
0 27527 7 2 2 61756 62159
0 27528 5 1 1 77189
0 27529 7 1 2 61421 77190
0 27530 5 1 1 27529
0 27531 7 1 2 27526 27530
0 27532 5 1 1 27531
0 27533 7 1 2 56359 27532
0 27534 5 1 1 27533
0 27535 7 1 2 27506 27534
0 27536 5 1 1 27535
0 27537 7 1 2 50781 27536
0 27538 5 1 1 27537
0 27539 7 1 2 53331 27538
0 27540 7 1 2 77147 27539
0 27541 5 1 1 27540
0 27542 7 1 2 61703 62160
0 27543 5 1 1 27542
0 27544 7 1 2 55917 61996
0 27545 7 1 2 27543 27544
0 27546 5 3 1 27545
0 27547 7 1 2 53216 77191
0 27548 5 1 1 27547
0 27549 7 1 2 50782 27548
0 27550 5 1 1 27549
0 27551 7 2 2 56360 61704
0 27552 5 1 1 77194
0 27553 7 1 2 70937 27552
0 27554 5 1 1 27553
0 27555 7 1 2 54679 70839
0 27556 7 1 2 27554 27555
0 27557 5 1 1 27556
0 27558 7 1 2 48521 75131
0 27559 5 1 1 27558
0 27560 7 1 2 50783 27559
0 27561 5 1 1 27560
0 27562 7 1 2 49352 27561
0 27563 5 1 1 27562
0 27564 7 1 2 27557 27563
0 27565 7 1 2 27550 27564
0 27566 5 1 1 27565
0 27567 7 1 2 54337 27566
0 27568 5 1 1 27567
0 27569 7 1 2 50784 24020
0 27570 5 1 1 27569
0 27571 7 2 2 60476 62107
0 27572 5 2 1 77196
0 27573 7 2 2 50233 77198
0 27574 5 1 1 77200
0 27575 7 1 2 76668 77201
0 27576 5 1 1 27575
0 27577 7 1 2 27570 27576
0 27578 5 1 1 27577
0 27579 7 1 2 53217 27578
0 27580 5 1 1 27579
0 27581 7 1 2 52304 61692
0 27582 5 1 1 27581
0 27583 7 1 2 61508 27582
0 27584 5 1 1 27583
0 27585 7 1 2 55695 27584
0 27586 5 1 1 27585
0 27587 7 1 2 63629 27586
0 27588 5 1 1 27587
0 27589 7 1 2 49466 27588
0 27590 5 1 1 27589
0 27591 7 1 2 76669 76960
0 27592 5 2 1 27591
0 27593 7 1 2 27590 77202
0 27594 5 1 1 27593
0 27595 7 1 2 53108 27594
0 27596 5 1 1 27595
0 27597 7 1 2 60091 70369
0 27598 7 1 2 26106 27597
0 27599 5 1 1 27598
0 27600 7 1 2 62359 27599
0 27601 5 2 1 27600
0 27602 7 1 2 57013 70435
0 27603 5 1 1 27602
0 27604 7 1 2 56361 27603
0 27605 5 2 1 27604
0 27606 7 1 2 47951 70872
0 27607 5 1 1 27606
0 27608 7 1 2 54680 27607
0 27609 7 1 2 77206 27608
0 27610 5 1 1 27609
0 27611 7 1 2 77204 27610
0 27612 5 1 1 27611
0 27613 7 1 2 54059 27612
0 27614 5 1 1 27613
0 27615 7 1 2 59745 1834
0 27616 5 1 1 27615
0 27617 7 1 2 54681 27616
0 27618 5 1 1 27617
0 27619 7 1 2 76708 27618
0 27620 5 1 1 27619
0 27621 7 1 2 62650 72928
0 27622 5 1 1 27621
0 27623 7 1 2 50473 27622
0 27624 7 1 2 27620 27623
0 27625 7 1 2 27614 27624
0 27626 7 1 2 27596 27625
0 27627 7 1 2 27580 27626
0 27628 5 1 1 27627
0 27629 7 1 2 27568 27628
0 27630 5 1 1 27629
0 27631 7 3 2 53109 76687
0 27632 5 1 1 77208
0 27633 7 1 2 50785 77209
0 27634 5 1 1 27633
0 27635 7 1 2 49578 27634
0 27636 7 1 2 27630 27635
0 27637 5 1 1 27636
0 27638 7 1 2 48621 27637
0 27639 7 1 2 27541 27638
0 27640 5 1 1 27639
0 27641 7 1 2 52424 60852
0 27642 5 1 1 27641
0 27643 7 1 2 63769 59752
0 27644 5 1 1 27643
0 27645 7 1 2 52305 27644
0 27646 5 1 1 27645
0 27647 7 1 2 27642 27646
0 27648 7 1 2 63394 27647
0 27649 5 1 1 27648
0 27650 7 1 2 50786 27649
0 27651 5 1 1 27650
0 27652 7 1 2 52425 73934
0 27653 5 1 1 27652
0 27654 7 1 2 49467 27653
0 27655 7 1 2 27651 27654
0 27656 5 1 1 27655
0 27657 7 1 2 59620 70987
0 27658 5 1 1 27657
0 27659 7 2 2 53110 60211
0 27660 7 1 2 48522 77211
0 27661 5 1 1 27660
0 27662 7 1 2 53218 27661
0 27663 7 1 2 27658 27662
0 27664 5 1 1 27663
0 27665 7 1 2 27656 27664
0 27666 5 1 1 27665
0 27667 7 1 2 52426 75777
0 27668 5 2 1 27667
0 27669 7 1 2 50474 76913
0 27670 5 1 1 27669
0 27671 7 2 2 53111 70464
0 27672 5 1 1 77215
0 27673 7 1 2 57014 77216
0 27674 5 1 1 27673
0 27675 7 1 2 27670 27674
0 27676 5 1 1 27675
0 27677 7 1 2 50234 27676
0 27678 5 1 1 27677
0 27679 7 1 2 77213 27678
0 27680 5 1 1 27679
0 27681 7 1 2 52306 27680
0 27682 5 1 1 27681
0 27683 7 1 2 57623 74830
0 27684 5 1 1 27683
0 27685 7 2 2 56121 27684
0 27686 5 1 1 77217
0 27687 7 1 2 56362 77218
0 27688 5 1 1 27687
0 27689 7 1 2 54060 69662
0 27690 7 1 2 27688 27689
0 27691 5 1 1 27690
0 27692 7 1 2 27682 27691
0 27693 5 1 1 27692
0 27694 7 1 2 54682 27693
0 27695 5 1 1 27694
0 27696 7 1 2 27666 27695
0 27697 5 1 1 27696
0 27698 7 1 2 57940 27697
0 27699 5 1 1 27698
0 27700 7 2 2 49468 75757
0 27701 7 1 2 58182 61909
0 27702 7 1 2 73922 71610
0 27703 7 1 2 27701 27702
0 27704 7 1 2 77219 27703
0 27705 5 1 1 27704
0 27706 7 1 2 27699 27705
0 27707 5 1 1 27706
0 27708 7 1 2 57234 27707
0 27709 5 1 1 27708
0 27710 7 5 2 50235 57015
0 27711 5 2 1 77221
0 27712 7 1 2 61629 77222
0 27713 5 1 1 27712
0 27714 7 1 2 57351 27713
0 27715 5 1 1 27714
0 27716 7 1 2 53332 1445
0 27717 5 1 1 27716
0 27718 7 1 2 55696 27717
0 27719 7 1 2 27715 27718
0 27720 5 1 1 27719
0 27721 7 1 2 50236 57354
0 27722 7 1 2 67255 27721
0 27723 5 1 1 27722
0 27724 7 1 2 27720 27723
0 27725 5 1 1 27724
0 27726 7 1 2 48622 27725
0 27727 5 1 1 27726
0 27728 7 2 2 53112 54061
0 27729 5 2 1 77228
0 27730 7 2 2 70894 77230
0 27731 7 1 2 60853 77232
0 27732 7 1 2 75646 27731
0 27733 5 1 1 27732
0 27734 7 1 2 27727 27733
0 27735 5 1 1 27734
0 27736 7 1 2 54338 27735
0 27737 5 1 1 27736
0 27738 7 1 2 70931 76114
0 27739 5 1 1 27738
0 27740 7 1 2 49353 76647
0 27741 5 1 1 27740
0 27742 7 1 2 27739 27741
0 27743 5 1 1 27742
0 27744 7 3 2 48623 50475
0 27745 5 3 1 77234
0 27746 7 1 2 49579 77235
0 27747 7 1 2 27743 27746
0 27748 5 1 1 27747
0 27749 7 1 2 27737 27748
0 27750 5 1 1 27749
0 27751 7 1 2 54683 27750
0 27752 5 1 1 27751
0 27753 7 1 2 48523 70982
0 27754 5 1 1 27753
0 27755 7 1 2 50787 27754
0 27756 5 1 1 27755
0 27757 7 2 2 70445 71607
0 27758 5 1 1 77240
0 27759 7 1 2 49469 27758
0 27760 7 1 2 27756 27759
0 27761 5 1 1 27760
0 27762 7 1 2 57941 24788
0 27763 7 1 2 68008 27762
0 27764 7 1 2 27761 27763
0 27765 5 1 1 27764
0 27766 7 1 2 27752 27765
0 27767 5 1 1 27766
0 27768 7 1 2 70370 27767
0 27769 5 1 1 27768
0 27770 7 3 2 53333 56925
0 27771 7 1 2 70216 77242
0 27772 5 1 1 27771
0 27773 7 4 2 55697 60477
0 27774 5 1 1 77245
0 27775 7 1 2 56363 27774
0 27776 5 1 1 27775
0 27777 7 3 2 57016 27776
0 27778 7 1 2 56213 59863
0 27779 5 1 1 27778
0 27780 7 1 2 48208 27779
0 27781 5 1 1 27780
0 27782 7 1 2 49580 27781
0 27783 7 1 2 77249 27782
0 27784 5 1 1 27783
0 27785 7 1 2 27772 27784
0 27786 5 1 1 27785
0 27787 7 1 2 48624 27786
0 27788 5 1 1 27787
0 27789 7 1 2 48524 75647
0 27790 7 1 2 70217 27789
0 27791 5 1 1 27790
0 27792 7 1 2 27788 27791
0 27793 5 1 1 27792
0 27794 7 1 2 58688 27793
0 27795 5 1 1 27794
0 27796 7 1 2 52307 61471
0 27797 5 1 1 27796
0 27798 7 1 2 48525 27797
0 27799 5 1 1 27798
0 27800 7 1 2 64277 76162
0 27801 7 1 2 27799 27800
0 27802 5 1 1 27801
0 27803 7 1 2 27795 27802
0 27804 5 1 1 27803
0 27805 7 1 2 60013 27804
0 27806 5 1 1 27805
0 27807 7 2 2 50788 76688
0 27808 7 1 2 59266 75375
0 27809 7 1 2 77252 27808
0 27810 7 1 2 77169 27809
0 27811 5 1 1 27810
0 27812 7 1 2 27806 27811
0 27813 7 1 2 27769 27812
0 27814 7 1 2 27709 27813
0 27815 7 1 2 27640 27814
0 27816 7 1 2 27482 27815
0 27817 5 1 1 27816
0 27818 7 1 2 55035 27817
0 27819 5 1 1 27818
0 27820 7 1 2 58532 56631
0 27821 5 1 1 27820
0 27822 7 1 2 59185 27821
0 27823 5 2 1 27822
0 27824 7 1 2 49470 77254
0 27825 5 2 1 27824
0 27826 7 1 2 27632 77256
0 27827 5 1 1 27826
0 27828 7 1 2 73188 27827
0 27829 5 1 1 27828
0 27830 7 1 2 51953 76370
0 27831 5 1 1 27830
0 27832 7 1 2 10157 27831
0 27833 5 1 1 27832
0 27834 7 1 2 57235 27833
0 27835 5 1 1 27834
0 27836 7 3 2 57624 56632
0 27837 5 5 1 77258
0 27838 7 1 2 58519 77261
0 27839 5 2 1 27838
0 27840 7 1 2 50237 77266
0 27841 5 1 1 27840
0 27842 7 1 2 27835 27841
0 27843 5 1 1 27842
0 27844 7 1 2 49471 27843
0 27845 5 1 1 27844
0 27846 7 2 2 54339 76914
0 27847 7 1 2 61615 77268
0 27848 5 1 1 27847
0 27849 7 1 2 50789 27848
0 27850 7 1 2 27845 27849
0 27851 5 1 1 27850
0 27852 7 2 2 57017 70371
0 27853 5 1 1 77270
0 27854 7 1 2 77000 75629
0 27855 5 1 1 27854
0 27856 7 1 2 76862 27855
0 27857 5 1 1 27856
0 27858 7 1 2 75421 27857
0 27859 5 1 1 27858
0 27860 7 1 2 77271 27859
0 27861 5 1 1 27860
0 27862 7 2 2 73599 73920
0 27863 5 1 1 77272
0 27864 7 1 2 75148 27863
0 27865 5 1 1 27864
0 27866 7 1 2 70938 27865
0 27867 5 1 1 27866
0 27868 7 2 2 61006 76674
0 27869 5 1 1 77274
0 27870 7 1 2 27672 27869
0 27871 5 1 1 27870
0 27872 7 1 2 56214 27871
0 27873 5 1 1 27872
0 27874 7 1 2 54684 27873
0 27875 7 1 2 27867 27874
0 27876 7 1 2 27861 27875
0 27877 5 1 1 27876
0 27878 7 1 2 27851 27877
0 27879 5 1 1 27878
0 27880 7 1 2 27829 27879
0 27881 5 1 1 27880
0 27882 7 1 2 57942 27881
0 27883 5 1 1 27882
0 27884 7 3 2 48526 53113
0 27885 5 3 1 77276
0 27886 7 1 2 54062 76899
0 27887 5 1 1 27886
0 27888 7 1 2 77279 27887
0 27889 5 1 1 27888
0 27890 7 1 2 51954 27889
0 27891 5 1 1 27890
0 27892 7 1 2 73192 77233
0 27893 5 1 1 27892
0 27894 7 2 2 48527 50238
0 27895 7 1 2 52994 77282
0 27896 5 1 1 27895
0 27897 7 1 2 54340 27896
0 27898 7 1 2 27893 27897
0 27899 7 1 2 27891 27898
0 27900 5 1 1 27899
0 27901 7 1 2 50476 66238
0 27902 5 1 1 27901
0 27903 7 1 2 54685 27902
0 27904 7 1 2 77220 27903
0 27905 7 1 2 27900 27904
0 27906 5 1 1 27905
0 27907 7 1 2 27883 27906
0 27908 5 1 1 27907
0 27909 7 1 2 55036 27908
0 27910 5 1 1 27909
0 27911 7 2 2 54341 62012
0 27912 7 1 2 67346 72966
0 27913 7 1 2 77284 27912
0 27914 5 1 1 27913
0 27915 7 1 2 27910 27914
0 27916 5 1 1 27915
0 27917 7 1 2 58438 27916
0 27918 5 1 1 27917
0 27919 7 1 2 51347 27918
0 27920 7 1 2 27819 27919
0 27921 7 1 2 27192 27920
0 27922 5 1 1 27921
0 27923 7 1 2 26860 27922
0 27924 5 1 1 27923
0 27925 7 1 2 53520 27924
0 27926 5 1 1 27925
0 27927 7 2 2 57625 60397
0 27928 7 1 2 56633 77286
0 27929 5 2 1 27928
0 27930 7 1 2 54063 76058
0 27931 5 1 1 27930
0 27932 7 1 2 54342 77108
0 27933 5 1 1 27932
0 27934 7 1 2 52427 27933
0 27935 7 1 2 27931 27934
0 27936 5 1 1 27935
0 27937 7 1 2 53219 27936
0 27938 5 1 1 27937
0 27939 7 1 2 77288 27938
0 27940 5 1 1 27939
0 27941 7 1 2 75758 27940
0 27942 5 1 1 27941
0 27943 7 6 2 52521 49472
0 27944 5 1 1 77290
0 27945 7 1 2 76692 27944
0 27946 5 2 1 27945
0 27947 7 1 2 59314 77170
0 27948 5 2 1 27947
0 27949 7 1 2 56748 70946
0 27950 5 1 1 27949
0 27951 7 1 2 77298 27950
0 27952 5 1 1 27951
0 27953 7 1 2 77296 27952
0 27954 5 1 1 27953
0 27955 7 1 2 58554 75725
0 27956 5 2 1 27955
0 27957 7 1 2 27954 77300
0 27958 5 1 1 27957
0 27959 7 1 2 54343 27958
0 27960 5 1 1 27959
0 27961 7 1 2 57236 63712
0 27962 5 2 1 27961
0 27963 7 1 2 70947 77297
0 27964 7 1 2 77302 27963
0 27965 5 1 1 27964
0 27966 7 1 2 77301 27965
0 27967 5 1 1 27966
0 27968 7 1 2 54064 27967
0 27969 5 1 1 27968
0 27970 7 1 2 77037 23046
0 27971 7 1 2 62467 27970
0 27972 5 1 1 27971
0 27973 7 1 2 27969 27972
0 27974 7 1 2 27960 27973
0 27975 5 1 1 27974
0 27976 7 1 2 53334 27975
0 27977 5 1 1 27976
0 27978 7 1 2 27942 27977
0 27979 5 1 1 27978
0 27980 7 1 2 51064 27979
0 27981 5 1 1 27980
0 27982 7 2 2 73274 77269
0 27983 5 1 1 77304
0 27984 7 1 2 55037 77305
0 27985 5 1 1 27984
0 27986 7 1 2 52428 76224
0 27987 5 1 1 27986
0 27988 7 1 2 25459 27987
0 27989 5 3 1 27988
0 27990 7 2 2 48625 77306
0 27991 5 1 1 77309
0 27992 7 1 2 75649 27991
0 27993 5 2 1 27992
0 27994 7 1 2 63701 77311
0 27995 5 1 1 27994
0 27996 7 2 2 76327 75699
0 27997 5 1 1 77313
0 27998 7 2 2 54344 77314
0 27999 5 1 1 77315
0 28000 7 1 2 52522 77316
0 28001 5 1 1 28000
0 28002 7 1 2 27995 28001
0 28003 5 1 1 28002
0 28004 7 1 2 60986 28003
0 28005 5 1 1 28004
0 28006 7 1 2 27985 28005
0 28007 5 1 1 28006
0 28008 7 1 2 50239 28007
0 28009 5 1 1 28008
0 28010 7 1 2 50240 60987
0 28011 5 3 1 28010
0 28012 7 1 2 49354 77317
0 28013 5 1 1 28012
0 28014 7 6 2 55038 56634
0 28015 7 2 2 56215 77320
0 28016 5 1 1 77326
0 28017 7 1 2 4973 28016
0 28018 5 1 1 28017
0 28019 7 1 2 75759 28018
0 28020 5 1 1 28019
0 28021 7 3 2 49473 56458
0 28022 5 1 1 77328
0 28023 7 1 2 77321 77329
0 28024 5 1 1 28023
0 28025 7 1 2 56216 76182
0 28026 5 1 1 28025
0 28027 7 1 2 28024 28026
0 28028 7 1 2 28020 28027
0 28029 5 1 1 28028
0 28030 7 1 2 52308 28029
0 28031 5 1 1 28030
0 28032 7 1 2 76696 75837
0 28033 5 1 1 28032
0 28034 7 1 2 28031 28033
0 28035 5 1 1 28034
0 28036 7 1 2 28013 28035
0 28037 5 1 1 28036
0 28038 7 1 2 54345 70392
0 28039 7 1 2 77192 28038
0 28040 5 1 1 28039
0 28041 7 1 2 77280 28040
0 28042 5 1 1 28041
0 28043 7 1 2 56459 76328
0 28044 7 1 2 28042 28043
0 28045 5 1 1 28044
0 28046 7 1 2 66902 76614
0 28047 5 1 1 28046
0 28048 7 2 2 52163 76237
0 28049 5 1 1 77331
0 28050 7 3 2 71844 68295
0 28051 5 1 1 77333
0 28052 7 1 2 77332 77334
0 28053 5 1 1 28052
0 28054 7 1 2 76615 75424
0 28055 5 2 1 28054
0 28056 7 1 2 28053 77336
0 28057 5 1 1 28056
0 28058 7 1 2 52309 28057
0 28059 5 1 1 28058
0 28060 7 1 2 28047 28059
0 28061 7 1 2 70770 77335
0 28062 5 1 1 28061
0 28063 7 1 2 77337 28062
0 28064 5 1 1 28063
0 28065 7 1 2 56635 28064
0 28066 5 1 1 28065
0 28067 7 1 2 49581 66684
0 28068 5 1 1 28067
0 28069 7 1 2 27999 28068
0 28070 5 1 1 28069
0 28071 7 1 2 52523 28070
0 28072 5 1 1 28071
0 28073 7 1 2 28066 28072
0 28074 7 1 2 28060 28073
0 28075 5 1 1 28074
0 28076 7 1 2 52429 28075
0 28077 5 1 1 28076
0 28078 7 1 2 50790 28077
0 28079 7 1 2 28045 28078
0 28080 7 1 2 28037 28079
0 28081 7 1 2 28009 28080
0 28082 7 1 2 27981 28081
0 28083 5 1 1 28082
0 28084 7 1 2 54065 61262
0 28085 5 1 1 28084
0 28086 7 2 2 52310 28085
0 28087 5 1 1 77338
0 28088 7 1 2 56364 28087
0 28089 5 1 1 28088
0 28090 7 1 2 53114 28089
0 28091 5 1 1 28090
0 28092 7 4 2 76994 77005
0 28093 7 1 2 61562 62198
0 28094 7 1 2 77340 28093
0 28095 5 1 1 28094
0 28096 7 1 2 76948 26516
0 28097 5 1 1 28096
0 28098 7 1 2 76566 28097
0 28099 5 1 1 28098
0 28100 7 1 2 56217 66855
0 28101 5 1 1 28100
0 28102 7 2 2 57506 62161
0 28103 5 1 1 77344
0 28104 7 1 2 56926 77345
0 28105 5 1 1 28104
0 28106 7 1 2 28101 28105
0 28107 5 1 1 28106
0 28108 7 1 2 28099 28107
0 28109 7 1 2 28095 28108
0 28110 5 1 1 28109
0 28111 7 1 2 28091 28110
0 28112 5 1 1 28111
0 28113 7 1 2 61286 76961
0 28114 5 1 1 28113
0 28115 7 1 2 77066 28114
0 28116 5 1 1 28115
0 28117 7 1 2 48403 28116
0 28118 5 1 1 28117
0 28119 7 1 2 48209 59830
0 28120 5 1 1 28119
0 28121 7 1 2 61281 28120
0 28122 5 1 1 28121
0 28123 7 1 2 62861 28122
0 28124 5 1 1 28123
0 28125 7 1 2 28118 28124
0 28126 7 1 2 28112 28125
0 28127 5 1 1 28126
0 28128 7 1 2 54346 28127
0 28129 5 1 1 28128
0 28130 7 2 2 49474 77277
0 28131 5 1 1 77346
0 28132 7 1 2 28129 28131
0 28133 5 1 1 28132
0 28134 7 1 2 56460 28133
0 28135 5 1 1 28134
0 28136 7 1 2 76970 27853
0 28137 5 1 1 28136
0 28138 7 1 2 57018 76973
0 28139 5 1 1 28138
0 28140 7 1 2 72934 28139
0 28141 5 1 1 28140
0 28142 7 1 2 28137 28141
0 28143 5 1 1 28142
0 28144 7 1 2 56365 28143
0 28145 5 1 1 28144
0 28146 7 1 2 52902 28145
0 28147 5 1 1 28146
0 28148 7 1 2 50105 58923
0 28149 7 1 2 212 28148
0 28150 5 1 1 28149
0 28151 7 1 2 28147 28150
0 28152 5 1 1 28151
0 28153 7 1 2 51955 28152
0 28154 5 1 1 28153
0 28155 7 2 2 60854 70640
0 28156 5 1 1 77348
0 28157 7 1 2 57019 77349
0 28158 5 1 1 28157
0 28159 7 1 2 55781 64949
0 28160 5 1 1 28159
0 28161 7 1 2 56218 28160
0 28162 5 1 1 28161
0 28163 7 1 2 28158 28162
0 28164 7 1 2 28154 28163
0 28165 5 1 1 28164
0 28166 7 1 2 75760 28165
0 28167 5 1 1 28166
0 28168 7 5 2 70773 72929
0 28169 7 1 2 49582 50241
0 28170 7 1 2 60643 28169
0 28171 7 1 2 77350 28170
0 28172 5 1 1 28171
0 28173 7 1 2 28167 28172
0 28174 7 1 2 28135 28173
0 28175 5 1 1 28174
0 28176 7 1 2 51065 28175
0 28177 5 1 1 28176
0 28178 7 1 2 48404 76971
0 28179 5 1 1 28178
0 28180 7 1 2 76976 28179
0 28181 5 1 1 28180
0 28182 7 1 2 60107 28181
0 28183 5 1 1 28182
0 28184 7 1 2 51956 28183
0 28185 5 1 1 28184
0 28186 7 1 2 74896 28185
0 28187 5 1 1 28186
0 28188 7 1 2 56636 28187
0 28189 5 1 1 28188
0 28190 7 1 2 71014 74831
0 28191 5 1 1 28190
0 28192 7 1 2 28189 28191
0 28193 5 1 1 28192
0 28194 7 1 2 57020 28193
0 28195 5 1 1 28194
0 28196 7 1 2 60836 62152
0 28197 5 4 1 28196
0 28198 7 1 2 70393 77355
0 28199 5 1 1 28198
0 28200 7 3 2 59938 55698
0 28201 5 5 1 77359
0 28202 7 1 2 56122 77362
0 28203 7 1 2 28199 28202
0 28204 5 1 1 28203
0 28205 7 1 2 56219 28204
0 28206 5 1 1 28205
0 28207 7 1 2 28195 28206
0 28208 5 1 1 28207
0 28209 7 2 2 75680 28208
0 28210 7 1 2 75425 77367
0 28211 5 1 1 28210
0 28212 7 1 2 54686 28211
0 28213 7 1 2 28177 28212
0 28214 5 1 1 28213
0 28215 7 1 2 28083 28214
0 28216 5 1 1 28215
0 28217 7 1 2 76341 76085
0 28218 5 1 1 28217
0 28219 7 1 2 76089 28218
0 28220 5 1 1 28219
0 28221 7 1 2 49355 28220
0 28222 5 1 1 28221
0 28223 7 1 2 59939 67397
0 28224 5 1 1 28223
0 28225 7 1 2 59222 28224
0 28226 5 2 1 28225
0 28227 7 1 2 63458 77369
0 28228 5 1 1 28227
0 28229 7 1 2 28222 28228
0 28230 5 1 1 28229
0 28231 7 1 2 54347 28230
0 28232 5 1 1 28231
0 28233 7 1 2 58533 60855
0 28234 5 1 1 28233
0 28235 7 1 2 63131 60644
0 28236 5 2 1 28235
0 28237 7 1 2 28234 77371
0 28238 5 1 1 28237
0 28239 7 1 2 55039 62651
0 28240 7 1 2 28238 28239
0 28241 5 1 1 28240
0 28242 7 1 2 53335 28241
0 28243 7 1 2 28232 28242
0 28244 5 1 1 28243
0 28245 7 1 2 49475 59883
0 28246 5 1 1 28245
0 28247 7 1 2 55699 74908
0 28248 7 1 2 73234 28247
0 28249 5 1 1 28248
0 28250 7 1 2 28246 28249
0 28251 5 1 1 28250
0 28252 7 1 2 57626 28251
0 28253 5 1 1 28252
0 28254 7 1 2 73232 76954
0 28255 5 1 1 28254
0 28256 7 1 2 63415 66044
0 28257 5 1 1 28256
0 28258 7 1 2 28255 28257
0 28259 7 1 2 28253 28258
0 28260 5 1 1 28259
0 28261 7 1 2 50791 28260
0 28262 5 1 1 28261
0 28263 7 1 2 60014 70939
0 28264 5 1 1 28263
0 28265 7 1 2 56366 28264
0 28266 5 2 1 28265
0 28267 7 1 2 63515 77373
0 28268 5 1 1 28267
0 28269 7 1 2 49583 28268
0 28270 7 1 2 28262 28269
0 28271 5 1 1 28270
0 28272 7 1 2 52524 28271
0 28273 7 1 2 28244 28272
0 28274 5 1 1 28273
0 28275 7 1 2 53336 75562
0 28276 5 1 1 28275
0 28277 7 4 2 48626 53220
0 28278 5 1 1 77375
0 28279 7 1 2 76700 28278
0 28280 5 6 1 28279
0 28281 7 1 2 49584 77379
0 28282 7 1 2 58571 28281
0 28283 5 1 1 28282
0 28284 7 1 2 28276 28283
0 28285 5 1 1 28284
0 28286 7 1 2 59940 28285
0 28287 5 1 1 28286
0 28288 7 3 2 56556 57355
0 28289 7 1 2 77385 77287
0 28290 5 1 1 28289
0 28291 7 1 2 28287 28290
0 28292 5 1 1 28291
0 28293 7 1 2 55700 28292
0 28294 5 1 1 28293
0 28295 7 1 2 63132 77310
0 28296 5 1 1 28295
0 28297 7 1 2 28294 28296
0 28298 5 1 1 28297
0 28299 7 1 2 50792 28298
0 28300 5 1 1 28299
0 28301 7 5 2 48627 75437
0 28302 5 1 1 77388
0 28303 7 1 2 77389 77374
0 28304 5 1 1 28303
0 28305 7 1 2 28300 28304
0 28306 5 1 1 28305
0 28307 7 1 2 51066 28306
0 28308 5 1 1 28307
0 28309 7 1 2 55701 61453
0 28310 5 1 1 28309
0 28311 7 1 2 59768 28310
0 28312 5 1 1 28311
0 28313 7 2 2 56220 75551
0 28314 5 1 1 77393
0 28315 7 1 2 55040 77394
0 28316 7 1 2 28312 28315
0 28317 5 1 1 28316
0 28318 7 1 2 28308 28317
0 28319 7 2 2 28274 28318
0 28320 5 1 1 77395
0 28321 7 1 2 61499 76915
0 28322 5 1 1 28321
0 28323 7 1 2 71419 73250
0 28324 5 1 1 28323
0 28325 7 1 2 28322 28324
0 28326 5 1 1 28325
0 28327 7 1 2 54348 28326
0 28328 5 1 1 28327
0 28329 7 1 2 49476 61500
0 28330 5 1 1 28329
0 28331 7 1 2 50242 76352
0 28332 5 1 1 28331
0 28333 7 1 2 28330 28332
0 28334 5 1 1 28333
0 28335 7 1 2 58534 28334
0 28336 5 1 1 28335
0 28337 7 1 2 28328 28336
0 28338 5 1 1 28337
0 28339 7 1 2 53337 28338
0 28340 5 1 1 28339
0 28341 7 1 2 51957 73251
0 28342 7 1 2 76794 28341
0 28343 5 1 1 28342
0 28344 7 1 2 28340 28343
0 28345 5 1 1 28344
0 28346 7 1 2 55041 28345
0 28347 5 1 1 28346
0 28348 7 2 2 71420 70940
0 28349 5 1 1 77397
0 28350 7 2 2 59799 74268
0 28351 5 1 1 77399
0 28352 7 1 2 28349 28351
0 28353 5 1 1 28352
0 28354 7 1 2 67332 28353
0 28355 5 1 1 28354
0 28356 7 1 2 28347 28355
0 28357 5 1 1 28356
0 28358 7 1 2 52525 28357
0 28359 5 1 1 28358
0 28360 7 1 2 75515 77398
0 28361 5 1 1 28360
0 28362 7 1 2 77386 77400
0 28363 5 1 1 28362
0 28364 7 1 2 28361 28363
0 28365 5 1 1 28364
0 28366 7 1 2 51067 28365
0 28367 5 1 1 28366
0 28368 7 2 2 53338 66031
0 28369 7 1 2 60600 68933
0 28370 7 1 2 77376 28369
0 28371 7 1 2 77401 28370
0 28372 5 1 1 28371
0 28373 7 1 2 28367 28372
0 28374 7 1 2 28359 28373
0 28375 5 2 1 28374
0 28376 7 1 2 58439 77403
0 28377 5 1 1 28376
0 28378 7 1 2 77396 28377
0 28379 5 1 1 28378
0 28380 7 1 2 57237 28379
0 28381 5 1 1 28380
0 28382 7 3 2 52311 76935
0 28383 5 1 1 77405
0 28384 7 2 2 53115 60151
0 28385 5 1 1 77408
0 28386 7 1 2 56927 28385
0 28387 7 1 2 28383 28386
0 28388 5 1 1 28387
0 28389 7 2 2 50793 28388
0 28390 7 1 2 49227 76995
0 28391 5 1 1 28390
0 28392 7 1 2 56123 62058
0 28393 5 2 1 28392
0 28394 7 1 2 28391 77412
0 28395 5 1 1 28394
0 28396 7 1 2 59995 28395
0 28397 5 1 1 28396
0 28398 7 1 2 55782 62759
0 28399 7 1 2 72664 28398
0 28400 5 1 1 28399
0 28401 7 1 2 63256 74789
0 28402 5 1 1 28401
0 28403 7 1 2 49228 28402
0 28404 5 1 1 28403
0 28405 7 1 2 59194 28404
0 28406 7 1 2 28400 28405
0 28407 7 1 2 28397 28406
0 28408 5 1 1 28407
0 28409 7 1 2 77410 28408
0 28410 5 1 1 28409
0 28411 7 2 2 49477 77002
0 28412 7 1 2 76967 77414
0 28413 5 1 1 28412
0 28414 7 1 2 77203 28413
0 28415 5 1 1 28414
0 28416 7 1 2 52995 28415
0 28417 5 1 1 28416
0 28418 7 1 2 77231 24122
0 28419 7 1 2 27574 28418
0 28420 5 1 1 28419
0 28421 7 1 2 75781 28420
0 28422 5 1 1 28421
0 28423 7 1 2 25878 77064
0 28424 5 1 1 28423
0 28425 7 1 2 52430 28424
0 28426 5 1 1 28425
0 28427 7 1 2 50243 77210
0 28428 5 1 1 28427
0 28429 7 1 2 28426 28428
0 28430 5 1 1 28429
0 28431 7 1 2 63257 28430
0 28432 5 2 1 28431
0 28433 7 1 2 28422 77416
0 28434 7 1 2 28417 28433
0 28435 7 1 2 28410 28434
0 28436 5 1 1 28435
0 28437 7 1 2 52526 28436
0 28438 5 1 1 28437
0 28439 7 2 2 77250 75946
0 28440 5 1 1 77418
0 28441 7 1 2 77409 77419
0 28442 5 1 1 28441
0 28443 7 1 2 77406 76060
0 28444 5 1 1 28443
0 28445 7 1 2 28442 28444
0 28446 5 1 1 28445
0 28447 7 1 2 50794 28446
0 28448 5 1 1 28447
0 28449 7 2 2 52431 48628
0 28450 5 1 1 77420
0 28451 7 2 2 58820 77421
0 28452 7 1 2 58893 76648
0 28453 7 1 2 77422 28452
0 28454 5 1 1 28453
0 28455 7 2 2 28448 28454
0 28456 7 1 2 28438 77424
0 28457 5 1 1 28456
0 28458 7 1 2 53339 28457
0 28459 5 1 1 28458
0 28460 7 2 2 70153 76225
0 28461 5 1 1 77426
0 28462 7 1 2 22401 9427
0 28463 5 1 1 28462
0 28464 7 1 2 53116 28463
0 28465 5 1 1 28464
0 28466 7 1 2 50795 77407
0 28467 5 1 1 28466
0 28468 7 1 2 28465 28467
0 28469 5 1 1 28468
0 28470 7 1 2 77427 28469
0 28471 5 1 1 28470
0 28472 7 1 2 28459 28471
0 28473 5 1 1 28472
0 28474 7 1 2 55042 28473
0 28475 5 1 1 28474
0 28476 7 2 2 63516 75761
0 28477 7 1 2 60093 71050
0 28478 5 1 1 28477
0 28479 7 1 2 77428 28478
0 28480 5 1 1 28479
0 28481 7 1 2 61596 25803
0 28482 5 2 1 28481
0 28483 7 1 2 64711 75438
0 28484 7 1 2 77430 28483
0 28485 5 1 1 28484
0 28486 7 1 2 60152 63808
0 28487 7 1 2 75399 28486
0 28488 5 1 1 28487
0 28489 7 1 2 63543 28488
0 28490 5 1 1 28489
0 28491 7 1 2 49585 60069
0 28492 7 1 2 28490 28491
0 28493 5 1 1 28492
0 28494 7 1 2 52527 28493
0 28495 7 1 2 28485 28494
0 28496 5 1 1 28495
0 28497 7 2 2 53340 63517
0 28498 5 3 1 77432
0 28499 7 1 2 60070 77433
0 28500 5 1 1 28499
0 28501 7 1 2 48629 28500
0 28502 5 1 1 28501
0 28503 7 1 2 52312 28502
0 28504 7 1 2 28496 28503
0 28505 5 1 1 28504
0 28506 7 1 2 28480 28505
0 28507 5 1 1 28506
0 28508 7 1 2 57021 28507
0 28509 5 1 1 28508
0 28510 7 1 2 61291 75654
0 28511 5 1 1 28510
0 28512 7 2 2 56124 67212
0 28513 7 2 2 52903 62219
0 28514 5 2 1 77439
0 28515 7 1 2 61247 77440
0 28516 5 1 1 28515
0 28517 7 1 2 77437 28516
0 28518 5 1 1 28517
0 28519 7 2 2 28511 28518
0 28520 5 1 1 77443
0 28521 7 1 2 53341 77444
0 28522 5 1 1 28521
0 28523 7 1 2 52528 75770
0 28524 5 1 1 28523
0 28525 7 1 2 49586 28440
0 28526 7 1 2 28524 28525
0 28527 5 1 1 28526
0 28528 7 1 2 50244 28527
0 28529 7 1 2 28522 28528
0 28530 5 1 1 28529
0 28531 7 1 2 61610 70362
0 28532 5 2 1 28531
0 28533 7 1 2 77312 77445
0 28534 5 1 1 28533
0 28535 7 1 2 50796 28534
0 28536 7 1 2 28530 28535
0 28537 5 1 1 28536
0 28538 7 1 2 70501 76186
0 28539 5 1 1 28538
0 28540 7 1 2 58572 28539
0 28541 5 1 1 28540
0 28542 7 1 2 69881 28541
0 28543 5 1 1 28542
0 28544 7 1 2 56367 61600
0 28545 5 1 1 28544
0 28546 7 1 2 62347 28545
0 28547 5 1 1 28546
0 28548 7 1 2 48405 28547
0 28549 5 1 1 28548
0 28550 7 1 2 56368 62313
0 28551 5 1 1 28550
0 28552 7 1 2 57022 28551
0 28553 7 1 2 28549 28552
0 28554 7 2 2 28543 28553
0 28555 5 1 1 77447
0 28556 7 1 2 56461 28555
0 28557 5 1 1 28556
0 28558 7 2 2 61639 77246
0 28559 5 1 1 77449
0 28560 7 3 2 49587 57321
0 28561 5 2 1 77451
0 28562 7 1 2 75523 77454
0 28563 5 3 1 28562
0 28564 7 1 2 77450 77456
0 28565 5 1 1 28564
0 28566 7 1 2 54687 75767
0 28567 7 1 2 28565 28566
0 28568 7 1 2 28557 28567
0 28569 5 1 1 28568
0 28570 7 1 2 51068 28569
0 28571 7 1 2 28537 28570
0 28572 5 1 1 28571
0 28573 7 1 2 28509 28572
0 28574 7 1 2 28475 28573
0 28575 5 1 1 28574
0 28576 7 1 2 50477 28575
0 28577 5 1 1 28576
0 28578 7 1 2 28381 28577
0 28579 7 1 2 28216 28578
0 28580 5 1 1 28579
0 28581 7 1 2 51348 28580
0 28582 5 1 1 28581
0 28583 7 2 2 73217 73220
0 28584 5 1 1 77459
0 28585 7 2 2 53117 49588
0 28586 7 1 2 51069 77461
0 28587 5 1 1 28586
0 28588 7 1 2 27997 28587
0 28589 5 1 1 28588
0 28590 7 1 2 52529 28589
0 28591 5 1 1 28590
0 28592 7 1 2 70682 77387
0 28593 5 1 1 28592
0 28594 7 1 2 28591 28593
0 28595 5 1 1 28594
0 28596 7 1 2 59941 28595
0 28597 5 1 1 28596
0 28598 7 1 2 55043 77229
0 28599 5 1 1 28598
0 28600 7 1 2 75753 28599
0 28601 5 1 1 28600
0 28602 7 1 2 57023 4438
0 28603 7 1 2 28601 28602
0 28604 5 1 1 28603
0 28605 7 1 2 28597 28604
0 28606 5 1 1 28605
0 28607 7 1 2 54688 28606
0 28608 5 1 1 28607
0 28609 7 1 2 51958 70154
0 28610 7 1 2 73524 76616
0 28611 7 1 2 28609 28610
0 28612 5 1 1 28611
0 28613 7 1 2 28608 28612
0 28614 5 1 1 28613
0 28615 7 1 2 70372 28614
0 28616 5 1 1 28615
0 28617 7 3 2 50245 61630
0 28618 5 1 1 77463
0 28619 7 1 2 53342 76709
0 28620 5 1 1 28619
0 28621 7 1 2 72930 77307
0 28622 5 2 1 28621
0 28623 7 1 2 28620 77466
0 28624 5 1 1 28623
0 28625 7 1 2 52530 28624
0 28626 5 1 1 28625
0 28627 7 2 2 52164 71092
0 28628 7 1 2 76238 75516
0 28629 7 1 2 77468 28628
0 28630 5 2 1 28629
0 28631 7 1 2 28626 77470
0 28632 5 1 1 28631
0 28633 7 1 2 77464 28632
0 28634 5 1 1 28633
0 28635 7 1 2 61910 70170
0 28636 5 1 1 28635
0 28637 7 1 2 28634 28636
0 28638 5 1 1 28637
0 28639 7 1 2 55044 28638
0 28640 5 1 1 28639
0 28641 7 2 2 55045 71288
0 28642 5 2 1 77472
0 28643 7 1 2 67343 77474
0 28644 5 1 1 28643
0 28645 7 1 2 77380 77465
0 28646 7 1 2 28644 28645
0 28647 5 1 1 28646
0 28648 7 3 2 52313 75426
0 28649 5 1 1 77476
0 28650 7 1 2 66905 28649
0 28651 5 1 1 28650
0 28652 7 1 2 77308 28651
0 28653 5 1 1 28652
0 28654 7 1 2 67333 77291
0 28655 5 1 1 28654
0 28656 7 1 2 76061 77473
0 28657 5 1 1 28656
0 28658 7 1 2 28655 28657
0 28659 7 1 2 28653 28658
0 28660 7 1 2 28647 28659
0 28661 5 1 1 28660
0 28662 7 1 2 71495 28661
0 28663 5 1 1 28662
0 28664 7 1 2 28640 28663
0 28665 7 2 2 28616 28664
0 28666 5 1 1 77479
0 28667 7 1 2 71603 77381
0 28668 5 1 1 28667
0 28669 7 1 2 55046 70106
0 28670 5 1 1 28669
0 28671 7 1 2 28668 28670
0 28672 5 1 1 28671
0 28673 7 1 2 49589 28672
0 28674 5 1 1 28673
0 28675 7 1 2 53343 75947
0 28676 7 1 2 76038 28675
0 28677 5 1 1 28676
0 28678 7 1 2 28674 28677
0 28679 5 1 1 28678
0 28680 7 1 2 50797 28679
0 28681 5 1 1 28680
0 28682 7 1 2 63518 70436
0 28683 7 1 2 77457 28682
0 28684 5 1 1 28683
0 28685 7 1 2 28681 28684
0 28686 5 1 1 28685
0 28687 7 2 2 57238 28686
0 28688 7 1 2 60015 77481
0 28689 5 1 1 28688
0 28690 7 3 2 53344 56637
0 28691 5 1 1 77483
0 28692 7 1 2 61911 77484
0 28693 5 1 1 28692
0 28694 7 1 2 65223 75344
0 28695 7 1 2 70494 28694
0 28696 5 1 1 28695
0 28697 7 1 2 28693 28696
0 28698 5 1 1 28697
0 28699 7 2 2 77477 28698
0 28700 5 1 1 77486
0 28701 7 1 2 60016 77429
0 28702 5 1 1 28701
0 28703 7 1 2 28700 28702
0 28704 5 1 1 28703
0 28705 7 1 2 57024 28704
0 28706 5 1 1 28705
0 28707 7 1 2 28689 28706
0 28708 7 1 2 77480 28707
0 28709 5 1 1 28708
0 28710 7 1 2 51349 28709
0 28711 5 1 1 28710
0 28712 7 1 2 28584 28711
0 28713 5 1 1 28712
0 28714 7 1 2 58440 28713
0 28715 5 1 1 28714
0 28716 7 1 2 73525 71256
0 28717 5 1 1 28716
0 28718 7 2 2 49590 59903
0 28719 5 1 1 77488
0 28720 7 1 2 28717 28719
0 28721 5 1 1 28720
0 28722 7 1 2 77382 28721
0 28723 5 1 1 28722
0 28724 7 2 2 55047 57025
0 28725 7 1 2 60269 75230
0 28726 7 1 2 77490 28725
0 28727 5 1 1 28726
0 28728 7 1 2 28723 28727
0 28729 5 1 1 28728
0 28730 7 1 2 52314 28729
0 28731 5 1 1 28730
0 28732 7 1 2 28022 75768
0 28733 5 2 1 28732
0 28734 7 4 2 51959 55048
0 28735 7 1 2 77492 77494
0 28736 5 1 1 28735
0 28737 7 1 2 28731 28736
0 28738 5 1 1 28737
0 28739 7 1 2 50798 28738
0 28740 5 1 1 28739
0 28741 7 1 2 52531 76689
0 28742 7 1 2 76390 28741
0 28743 5 1 1 28742
0 28744 7 2 2 51070 76928
0 28745 5 1 1 77498
0 28746 7 1 2 60153 77499
0 28747 7 1 2 77458 28746
0 28748 5 1 1 28747
0 28749 7 1 2 28743 28748
0 28750 7 1 2 28740 28749
0 28751 5 1 1 28750
0 28752 7 1 2 53118 28751
0 28753 5 1 1 28752
0 28754 7 1 2 76916 76929
0 28755 5 1 1 28754
0 28756 7 1 2 25680 28755
0 28757 5 1 1 28756
0 28758 7 1 2 75838 28757
0 28759 5 1 1 28758
0 28760 7 1 2 73414 68934
0 28761 5 1 1 28760
0 28762 7 1 2 63544 28761
0 28763 5 1 1 28762
0 28764 7 3 2 53221 63519
0 28765 5 1 1 77500
0 28766 7 1 2 48528 28765
0 28767 5 1 1 28766
0 28768 7 1 2 75762 28767
0 28769 7 1 2 28763 28768
0 28770 5 1 1 28769
0 28771 7 1 2 28759 28770
0 28772 5 1 1 28771
0 28773 7 1 2 50246 28772
0 28774 5 1 1 28773
0 28775 7 1 2 28753 28774
0 28776 5 2 1 28775
0 28777 7 1 2 51350 77503
0 28778 5 1 1 28777
0 28779 7 2 2 73252 76650
0 28780 7 1 2 60515 72424
0 28781 7 1 2 77505 28780
0 28782 5 1 1 28781
0 28783 7 5 2 51960 53345
0 28784 5 1 1 77507
0 28785 7 2 2 67199 77508
0 28786 5 1 1 77512
0 28787 7 2 2 71821 77513
0 28788 5 2 1 77514
0 28789 7 2 2 71369 77383
0 28790 7 1 2 49591 77518
0 28791 5 1 1 28790
0 28792 7 1 2 77516 28791
0 28793 5 1 1 28792
0 28794 7 1 2 51351 28793
0 28795 5 1 1 28794
0 28796 7 3 2 59884 63784
0 28797 7 1 2 70171 77520
0 28798 5 1 1 28797
0 28799 7 1 2 28795 28798
0 28800 5 1 1 28799
0 28801 7 1 2 52165 28800
0 28802 5 1 1 28801
0 28803 7 1 2 63736 70892
0 28804 7 1 2 77330 28803
0 28805 5 1 1 28804
0 28806 7 1 2 28802 28805
0 28807 5 1 1 28806
0 28808 7 1 2 57627 28807
0 28809 5 1 1 28808
0 28810 7 1 2 28782 28809
0 28811 7 1 2 28778 28810
0 28812 5 1 1 28811
0 28813 7 1 2 59864 28812
0 28814 5 1 1 28813
0 28815 7 1 2 53222 61030
0 28816 5 1 1 28815
0 28817 7 1 2 53346 28816
0 28818 7 1 2 76825 28817
0 28819 5 1 1 28818
0 28820 7 1 2 25658 28819
0 28821 5 1 1 28820
0 28822 7 1 2 52532 28821
0 28823 5 1 1 28822
0 28824 7 1 2 28314 28823
0 28825 5 1 1 28824
0 28826 7 2 2 73526 28825
0 28827 5 1 1 77523
0 28828 7 1 2 75199 77384
0 28829 5 1 1 28828
0 28830 7 2 2 52166 57322
0 28831 5 1 1 77525
0 28832 7 1 2 71421 77526
0 28833 5 1 1 28832
0 28834 7 1 2 28829 28833
0 28835 5 1 1 28834
0 28836 7 1 2 49592 28835
0 28837 5 1 1 28836
0 28838 7 2 2 52167 48630
0 28839 7 1 2 75430 77527
0 28840 5 1 1 28839
0 28841 7 1 2 28837 28840
0 28842 5 1 1 28841
0 28843 7 1 2 51071 28842
0 28844 5 1 1 28843
0 28845 7 1 2 28844 77517
0 28846 5 1 1 28845
0 28847 7 1 2 53119 28846
0 28848 5 1 1 28847
0 28849 7 1 2 28827 28848
0 28850 5 1 1 28849
0 28851 7 1 2 51352 28850
0 28852 5 1 1 28851
0 28853 7 1 2 66032 68396
0 28854 7 1 2 60522 28853
0 28855 7 2 2 75200 28854
0 28856 5 1 1 77529
0 28857 7 1 2 28852 28856
0 28858 5 1 1 28857
0 28859 7 1 2 70907 28858
0 28860 5 1 1 28859
0 28861 7 3 2 52315 60168
0 28862 7 2 2 71190 77531
0 28863 7 5 2 50799 60682
0 28864 7 1 2 77536 76473
0 28865 7 1 2 77534 28864
0 28866 5 1 1 28865
0 28867 7 1 2 28860 28866
0 28868 7 1 2 28814 28867
0 28869 7 1 2 28715 28868
0 28870 5 1 1 28869
0 28871 7 1 2 50478 28870
0 28872 5 1 1 28871
0 28873 7 1 2 53120 69159
0 28874 5 1 1 28873
0 28875 7 1 2 70980 28874
0 28876 5 2 1 28875
0 28877 7 1 2 60478 75948
0 28878 7 1 2 67709 28877
0 28879 5 1 1 28878
0 28880 7 1 2 76063 28879
0 28881 5 1 1 28880
0 28882 7 1 2 50800 28881
0 28883 5 1 1 28882
0 28884 7 2 2 65079 57854
0 28885 7 1 2 52533 62370
0 28886 7 1 2 77543 28885
0 28887 5 1 1 28886
0 28888 7 1 2 28883 28887
0 28889 5 1 1 28888
0 28890 7 1 2 49593 28889
0 28891 5 1 1 28890
0 28892 7 1 2 62371 75517
0 28893 7 1 2 77544 28892
0 28894 5 1 1 28893
0 28895 7 1 2 28891 28894
0 28896 5 2 1 28895
0 28897 7 1 2 51072 77545
0 28898 5 1 1 28897
0 28899 7 1 2 70373 68935
0 28900 7 2 2 77493 28899
0 28901 5 1 1 77547
0 28902 7 1 2 28898 28901
0 28903 5 1 1 28902
0 28904 7 1 2 51353 28903
0 28905 5 1 1 28904
0 28906 7 1 2 70437 73218
0 28907 5 1 1 28906
0 28908 7 1 2 28905 28907
0 28909 5 1 1 28908
0 28910 7 1 2 77541 28909
0 28911 5 1 1 28910
0 28912 7 2 2 71215 77521
0 28913 7 1 2 71285 76342
0 28914 7 2 2 76486 28913
0 28915 7 1 2 57239 77551
0 28916 7 1 2 77549 28915
0 28917 5 1 1 28916
0 28918 7 1 2 49766 28917
0 28919 7 1 2 28911 28918
0 28920 7 1 2 28872 28919
0 28921 7 1 2 28582 28920
0 28922 5 1 1 28921
0 28923 7 1 2 52658 28922
0 28924 7 1 2 27926 28923
0 28925 5 1 1 28924
0 28926 7 1 2 57507 72780
0 28927 5 2 1 28926
0 28928 7 1 2 60696 74700
0 28929 5 1 1 28928
0 28930 7 1 2 21037 28929
0 28931 5 1 1 28930
0 28932 7 1 2 56125 28931
0 28933 5 1 1 28932
0 28934 7 2 2 77553 28933
0 28935 5 1 1 77555
0 28936 7 1 2 65469 77556
0 28937 5 1 1 28936
0 28938 7 1 2 61950 62162
0 28939 5 1 1 28938
0 28940 7 1 2 53121 77339
0 28941 5 1 1 28940
0 28942 7 1 2 28939 28941
0 28943 5 1 1 28942
0 28944 7 1 2 54689 28943
0 28945 5 1 1 28944
0 28946 7 2 2 59942 70438
0 28947 5 1 1 77557
0 28948 7 1 2 70299 77558
0 28949 5 1 1 28948
0 28950 7 1 2 54349 28949
0 28951 7 1 2 28945 28950
0 28952 7 1 2 28937 28951
0 28953 5 1 1 28952
0 28954 7 1 2 48529 70471
0 28955 5 1 1 28954
0 28956 7 2 2 59721 59588
0 28957 5 2 1 77559
0 28958 7 1 2 59186 76053
0 28959 5 1 1 28958
0 28960 7 2 2 77561 28959
0 28961 5 1 1 77563
0 28962 7 1 2 58535 77564
0 28963 5 1 1 28962
0 28964 7 1 2 66255 28963
0 28965 5 1 1 28964
0 28966 7 1 2 28955 28965
0 28967 7 1 2 28953 28966
0 28968 5 1 1 28967
0 28969 7 1 2 49478 28968
0 28970 5 1 1 28969
0 28971 7 1 2 76353 25027
0 28972 7 1 2 76040 28971
0 28973 5 1 1 28972
0 28974 7 1 2 28970 28973
0 28975 5 1 1 28974
0 28976 7 1 2 53521 28975
0 28977 5 1 1 28976
0 28978 7 2 2 53522 58689
0 28979 7 1 2 59223 76054
0 28980 5 1 1 28979
0 28981 7 1 2 77562 28980
0 28982 5 1 1 28981
0 28983 7 1 2 77565 28982
0 28984 5 1 1 28983
0 28985 7 1 2 58919 70374
0 28986 7 1 2 76522 28985
0 28987 7 2 2 50801 58441
0 28988 5 2 1 77567
0 28989 7 1 2 47952 77569
0 28990 5 1 1 28989
0 28991 7 1 2 72800 28990
0 28992 7 1 2 28986 28991
0 28993 5 1 1 28992
0 28994 7 1 2 28984 28993
0 28995 5 1 1 28994
0 28996 7 1 2 50247 28995
0 28997 5 1 1 28996
0 28998 7 1 2 64464 76523
0 28999 7 1 2 59309 28998
0 29000 5 1 1 28999
0 29001 7 1 2 28997 29000
0 29002 7 1 2 28977 29001
0 29003 5 1 1 29002
0 29004 7 1 2 52534 29003
0 29005 5 1 1 29004
0 29006 7 1 2 54066 76055
0 29007 5 1 1 29006
0 29008 7 1 2 54350 61263
0 29009 5 1 1 29008
0 29010 7 1 2 65470 70741
0 29011 7 1 2 29009 29010
0 29012 7 1 2 29007 29011
0 29013 5 1 1 29012
0 29014 7 1 2 77267 77356
0 29015 5 1 1 29014
0 29016 7 1 2 59187 77372
0 29017 7 1 2 29015 29016
0 29018 7 1 2 72786 29017
0 29019 5 1 1 29018
0 29020 7 1 2 53223 29019
0 29021 7 1 2 29013 29020
0 29022 5 1 1 29021
0 29023 7 1 2 50248 63713
0 29024 5 1 1 29023
0 29025 7 1 2 76068 29024
0 29026 5 1 1 29025
0 29027 7 1 2 76670 29026
0 29028 5 1 1 29027
0 29029 7 1 2 56638 74269
0 29030 5 1 1 29029
0 29031 7 1 2 29028 29030
0 29032 5 1 1 29031
0 29033 7 1 2 57628 29032
0 29034 5 1 1 29033
0 29035 7 1 2 58536 62372
0 29036 7 1 2 72788 29035
0 29037 5 1 1 29036
0 29038 7 3 2 50249 70375
0 29039 5 1 1 77571
0 29040 7 2 2 60988 77572
0 29041 5 1 1 77574
0 29042 7 1 2 62652 77575
0 29043 5 1 1 29042
0 29044 7 1 2 66033 76930
0 29045 7 1 2 77357 29044
0 29046 5 1 1 29045
0 29047 7 1 2 29043 29046
0 29048 7 1 2 29037 29047
0 29049 7 1 2 29034 29048
0 29050 7 1 2 29022 29049
0 29051 5 2 1 29050
0 29052 7 1 2 48631 77576
0 29053 5 1 1 29052
0 29054 7 1 2 70394 77299
0 29055 5 1 1 29054
0 29056 7 1 2 54351 29055
0 29057 5 1 1 29056
0 29058 7 1 2 72537 77303
0 29059 5 1 1 29058
0 29060 7 1 2 59110 77038
0 29061 5 1 1 29060
0 29062 7 1 2 29059 29061
0 29063 7 1 2 29057 29062
0 29064 5 1 1 29063
0 29065 7 1 2 77253 29064
0 29066 5 1 1 29065
0 29067 7 1 2 29053 29066
0 29068 5 1 1 29067
0 29069 7 1 2 53523 29068
0 29070 5 1 1 29069
0 29071 7 1 2 29005 29070
0 29072 5 1 1 29071
0 29073 7 1 2 53347 29072
0 29074 5 1 1 29073
0 29075 7 1 2 52535 77577
0 29076 5 1 1 29075
0 29077 7 1 2 56126 29041
0 29078 5 1 1 29077
0 29079 7 1 2 48632 29078
0 29080 5 1 1 29079
0 29081 7 1 2 50802 77289
0 29082 7 1 2 29080 29081
0 29083 5 1 1 29082
0 29084 7 1 2 50250 58905
0 29085 5 3 1 29084
0 29086 7 1 2 54690 77578
0 29087 5 1 1 29086
0 29088 7 1 2 56221 29087
0 29089 7 1 2 29083 29088
0 29090 5 1 1 29089
0 29091 7 1 2 29076 29090
0 29092 5 1 1 29091
0 29093 7 1 2 72315 29092
0 29094 5 1 1 29093
0 29095 7 1 2 29074 29094
0 29096 5 1 1 29095
0 29097 7 1 2 51073 29096
0 29098 5 1 1 29097
0 29099 7 1 2 56749 71950
0 29100 5 1 1 29099
0 29101 7 1 2 54352 29100
0 29102 7 1 2 77193 29101
0 29103 5 1 1 29102
0 29104 7 1 2 77281 29103
0 29105 5 1 1 29104
0 29106 7 1 2 53224 29105
0 29107 5 1 1 29106
0 29108 7 1 2 77257 29107
0 29109 5 1 1 29108
0 29110 7 1 2 53348 29109
0 29111 5 1 1 29110
0 29112 7 1 2 58821 76226
0 29113 7 1 2 77469 29112
0 29114 5 1 1 29113
0 29115 7 1 2 29111 29114
0 29116 5 1 1 29115
0 29117 7 1 2 52536 29116
0 29118 5 1 1 29117
0 29119 7 1 2 67250 68009
0 29120 5 1 1 29119
0 29121 7 1 2 77467 29120
0 29122 5 1 1 29121
0 29123 7 1 2 52537 29122
0 29124 5 1 1 29123
0 29125 7 1 2 77471 29124
0 29126 5 1 1 29125
0 29127 7 1 2 60989 29126
0 29128 5 1 1 29127
0 29129 7 1 2 27983 29128
0 29130 5 1 1 29129
0 29131 7 1 2 50251 29130
0 29132 5 1 1 29131
0 29133 7 1 2 73415 71289
0 29134 7 1 2 77423 29133
0 29135 5 1 1 29134
0 29136 7 1 2 29132 29135
0 29137 7 1 2 29118 29136
0 29138 5 1 1 29137
0 29139 7 1 2 50803 29138
0 29140 5 1 1 29139
0 29141 7 1 2 77368 75722
0 29142 5 1 1 29141
0 29143 7 1 2 29140 29142
0 29144 5 1 1 29143
0 29145 7 1 2 74287 29144
0 29146 5 1 1 29145
0 29147 7 1 2 29098 29146
0 29148 5 1 1 29147
0 29149 7 1 2 51354 29148
0 29150 5 1 1 29149
0 29151 7 1 2 70941 77431
0 29152 5 1 1 29151
0 29153 7 1 2 49356 60350
0 29154 5 1 1 29153
0 29155 7 1 2 56222 29154
0 29156 5 1 1 29155
0 29157 7 1 2 29152 29156
0 29158 5 1 1 29157
0 29159 7 1 2 54691 29158
0 29160 5 1 1 29159
0 29161 7 1 2 77205 29160
0 29162 5 1 1 29161
0 29163 7 1 2 54067 29162
0 29164 5 1 1 29163
0 29165 7 1 2 56223 76078
0 29166 5 3 1 29165
0 29167 7 1 2 77411 77581
0 29168 5 1 1 29167
0 29169 7 1 2 77199 75782
0 29170 5 1 1 29169
0 29171 7 1 2 58828 77415
0 29172 5 1 1 29171
0 29173 7 1 2 29170 29172
0 29174 5 1 1 29173
0 29175 7 1 2 50252 29174
0 29176 5 1 1 29175
0 29177 7 1 2 77417 29176
0 29178 7 1 2 29168 29177
0 29179 7 1 2 29164 29178
0 29180 5 1 1 29179
0 29181 7 1 2 52538 29180
0 29182 5 1 1 29181
0 29183 7 1 2 77425 29182
0 29184 5 1 1 29183
0 29185 7 1 2 74288 29184
0 29186 5 1 1 29185
0 29187 7 1 2 48633 62772
0 29188 5 1 1 29187
0 29189 7 1 2 75952 29188
0 29190 5 1 1 29189
0 29191 7 1 2 77446 29190
0 29192 5 1 1 29191
0 29193 7 1 2 53524 28520
0 29194 5 1 1 29193
0 29195 7 1 2 75953 29194
0 29196 5 1 1 29195
0 29197 7 1 2 50253 29196
0 29198 5 1 1 29197
0 29199 7 1 2 29192 29198
0 29200 5 1 1 29199
0 29201 7 1 2 50804 29200
0 29202 5 1 1 29201
0 29203 7 1 2 52539 77448
0 29204 5 1 1 29203
0 29205 7 1 2 57323 68307
0 29206 7 1 2 29204 29205
0 29207 5 1 1 29206
0 29208 7 2 2 54692 76203
0 29209 5 1 1 77584
0 29210 7 1 2 75954 29209
0 29211 5 1 1 29210
0 29212 7 1 2 77247 29211
0 29213 5 1 1 29212
0 29214 7 1 2 76730 76204
0 29215 5 1 1 29214
0 29216 7 1 2 29213 29215
0 29217 5 1 1 29216
0 29218 7 1 2 61640 29217
0 29219 5 1 1 29218
0 29220 7 1 2 62348 70759
0 29221 5 1 1 29220
0 29222 7 1 2 72922 29221
0 29223 5 1 1 29222
0 29224 7 1 2 77585 29223
0 29225 5 1 1 29224
0 29226 7 1 2 58804 73860
0 29227 7 1 2 77248 29226
0 29228 5 1 1 29227
0 29229 7 1 2 29225 29228
0 29230 5 1 1 29229
0 29231 7 1 2 57026 29230
0 29232 5 1 1 29231
0 29233 7 1 2 29219 29232
0 29234 7 1 2 29207 29233
0 29235 7 1 2 29202 29234
0 29236 5 1 1 29235
0 29237 7 1 2 51074 29236
0 29238 5 1 1 29237
0 29239 7 1 2 29186 29238
0 29240 5 1 1 29239
0 29241 7 1 2 53349 29240
0 29242 5 1 1 29241
0 29243 7 1 2 50254 75771
0 29244 5 2 1 29243
0 29245 7 1 2 53225 77586
0 29246 5 2 1 29245
0 29247 7 1 2 70363 77587
0 29248 5 1 1 29247
0 29249 7 1 2 77588 29248
0 29250 5 1 1 29249
0 29251 7 1 2 50805 29250
0 29252 5 1 1 29251
0 29253 7 1 2 56928 28559
0 29254 5 1 1 29253
0 29255 7 1 2 60304 63143
0 29256 7 1 2 70826 29255
0 29257 5 1 1 29256
0 29258 7 1 2 29254 29257
0 29259 5 1 1 29258
0 29260 7 1 2 59478 29259
0 29261 5 1 1 29260
0 29262 7 1 2 52540 29261
0 29263 7 1 2 29252 29262
0 29264 5 1 1 29263
0 29265 7 4 2 50106 54693
0 29266 7 1 2 72759 77590
0 29267 5 1 1 29266
0 29268 7 1 2 76166 29267
0 29269 5 1 1 29268
0 29270 7 1 2 51961 29269
0 29271 5 1 1 29270
0 29272 7 2 2 71422 76872
0 29273 5 1 1 77594
0 29274 7 1 2 76167 29273
0 29275 5 1 1 29274
0 29276 7 1 2 52168 29275
0 29277 5 1 1 29276
0 29278 7 1 2 29271 29277
0 29279 5 1 1 29278
0 29280 7 1 2 52996 29279
0 29281 5 1 1 29280
0 29282 7 1 2 60131 62129
0 29283 5 1 1 29282
0 29284 7 1 2 76163 29283
0 29285 5 1 1 29284
0 29286 7 1 2 29281 29285
0 29287 5 1 1 29286
0 29288 7 1 2 53226 29287
0 29289 5 1 1 29288
0 29290 7 1 2 63613 76957
0 29291 5 1 1 29290
0 29292 7 1 2 29289 29291
0 29293 5 1 1 29292
0 29294 7 1 2 52432 29293
0 29295 5 1 1 29294
0 29296 7 2 2 72693 77537
0 29297 7 1 2 52997 77377
0 29298 7 1 2 77596 29297
0 29299 5 1 1 29298
0 29300 7 1 2 29295 29299
0 29301 7 1 2 29264 29300
0 29302 5 1 1 29301
0 29303 7 1 2 51075 29302
0 29304 5 1 1 29303
0 29305 7 1 2 66199 76931
0 29306 5 1 1 29305
0 29307 7 1 2 61501 65481
0 29308 7 1 2 70877 29307
0 29309 5 1 1 29308
0 29310 7 1 2 29306 29309
0 29311 5 1 1 29310
0 29312 7 1 2 57240 29311
0 29313 5 1 1 29312
0 29314 7 1 2 75201 77251
0 29315 5 1 1 29314
0 29316 7 1 2 75170 70868
0 29317 5 1 1 29316
0 29318 7 1 2 29315 29317
0 29319 5 1 1 29318
0 29320 7 1 2 53122 29319
0 29321 5 1 1 29320
0 29322 7 1 2 62379 72931
0 29323 5 1 1 29322
0 29324 7 1 2 29321 29323
0 29325 5 1 1 29324
0 29326 7 1 2 55049 29325
0 29327 5 1 1 29326
0 29328 7 1 2 29313 29327
0 29329 5 1 1 29328
0 29330 7 1 2 52541 29329
0 29331 5 1 1 29330
0 29332 7 1 2 29304 29331
0 29333 5 1 1 29332
0 29334 7 1 2 72316 29333
0 29335 5 1 1 29334
0 29336 7 1 2 29242 29335
0 29337 5 1 1 29336
0 29338 7 1 2 51355 29337
0 29339 5 1 1 29338
0 29340 7 1 2 53525 77460
0 29341 5 1 1 29340
0 29342 7 1 2 53526 28666
0 29343 5 1 1 29342
0 29344 7 1 2 53527 77482
0 29345 5 1 1 29344
0 29346 7 2 2 72932 70155
0 29347 7 1 2 65476 75485
0 29348 7 1 2 77598 29347
0 29349 5 1 1 29348
0 29350 7 1 2 29345 29349
0 29351 5 1 1 29350
0 29352 7 1 2 60017 29351
0 29353 5 1 1 29352
0 29354 7 1 2 49594 68308
0 29355 5 2 1 29354
0 29356 7 1 2 62428 75495
0 29357 5 1 1 29356
0 29358 7 1 2 77600 29357
0 29359 5 1 1 29358
0 29360 7 1 2 52542 29359
0 29361 5 1 1 29360
0 29362 7 1 2 53528 77390
0 29363 5 1 1 29362
0 29364 7 1 2 29361 29363
0 29365 5 1 1 29364
0 29366 7 1 2 60018 29365
0 29367 5 1 1 29366
0 29368 7 2 2 51962 73431
0 29369 7 1 2 49767 71286
0 29370 7 1 2 70495 29369
0 29371 7 1 2 77602 29370
0 29372 5 1 1 29371
0 29373 7 1 2 29367 29372
0 29374 5 1 1 29373
0 29375 7 1 2 51076 29374
0 29376 5 1 1 29375
0 29377 7 1 2 53529 77487
0 29378 5 1 1 29377
0 29379 7 1 2 29376 29378
0 29380 5 1 1 29379
0 29381 7 1 2 57027 29380
0 29382 5 1 1 29381
0 29383 7 1 2 58805 66716
0 29384 5 2 1 29383
0 29385 7 1 2 61631 62681
0 29386 7 1 2 77573 29385
0 29387 5 1 1 29386
0 29388 7 1 2 77604 29387
0 29389 5 1 1 29388
0 29390 7 1 2 70172 29389
0 29391 5 1 1 29390
0 29392 7 1 2 29382 29391
0 29393 7 1 2 29353 29392
0 29394 7 1 2 29343 29393
0 29395 5 1 1 29394
0 29396 7 1 2 51356 29395
0 29397 5 1 1 29396
0 29398 7 1 2 29341 29397
0 29399 5 1 1 29398
0 29400 7 1 2 58442 29399
0 29401 5 1 1 29400
0 29402 7 1 2 53530 77504
0 29403 5 1 1 29402
0 29404 7 1 2 51963 58213
0 29405 7 1 2 65022 29404
0 29406 5 1 1 29405
0 29407 7 1 2 70840 29406
0 29408 5 1 1 29407
0 29409 7 1 2 62682 71292
0 29410 7 1 2 29408 29409
0 29411 5 1 1 29410
0 29412 7 1 2 29403 29411
0 29413 5 1 1 29412
0 29414 7 1 2 51357 29413
0 29415 5 1 1 29414
0 29416 7 2 2 53350 62360
0 29417 5 1 1 77606
0 29418 7 2 2 75194 77607
0 29419 7 1 2 77506 77608
0 29420 5 1 1 29419
0 29421 7 1 2 72993 71822
0 29422 5 1 1 29421
0 29423 7 1 2 15879 29422
0 29424 5 1 1 29423
0 29425 7 1 2 57076 29424
0 29426 5 1 1 29425
0 29427 7 1 2 72317 77519
0 29428 5 1 1 29427
0 29429 7 1 2 29426 29428
0 29430 5 1 1 29429
0 29431 7 1 2 51358 29430
0 29432 5 1 1 29431
0 29433 7 1 2 70107 72889
0 29434 7 1 2 76605 29433
0 29435 5 1 1 29434
0 29436 7 1 2 29432 29435
0 29437 5 1 1 29436
0 29438 7 1 2 52169 29437
0 29439 5 1 1 29438
0 29440 7 2 2 63737 70156
0 29441 7 1 2 63674 76617
0 29442 7 1 2 77610 29441
0 29443 5 1 1 29442
0 29444 7 1 2 29439 29443
0 29445 5 1 1 29444
0 29446 7 1 2 57629 29445
0 29447 5 1 1 29446
0 29448 7 1 2 29420 29447
0 29449 7 1 2 29415 29448
0 29450 5 1 1 29449
0 29451 7 1 2 59865 29450
0 29452 5 1 1 29451
0 29453 7 2 2 53531 77550
0 29454 7 1 2 77535 77612
0 29455 5 1 1 29454
0 29456 7 1 2 53532 77515
0 29457 5 1 1 29456
0 29458 7 1 2 75877 77601
0 29459 5 1 1 29458
0 29460 7 1 2 56224 29459
0 29461 5 1 1 29460
0 29462 7 1 2 68309 75763
0 29463 5 1 1 29462
0 29464 7 1 2 29461 29463
0 29465 5 1 1 29464
0 29466 7 1 2 60270 29465
0 29467 5 1 1 29466
0 29468 7 1 2 75943 22882
0 29469 5 1 1 29468
0 29470 7 1 2 57028 29469
0 29471 7 1 2 75202 29470
0 29472 7 1 2 75882 29471
0 29473 5 1 1 29472
0 29474 7 1 2 29467 29473
0 29475 5 1 1 29474
0 29476 7 1 2 51077 29475
0 29477 5 1 1 29476
0 29478 7 1 2 29457 29477
0 29479 5 1 1 29478
0 29480 7 1 2 53123 29479
0 29481 5 1 1 29480
0 29482 7 1 2 53533 77524
0 29483 5 1 1 29482
0 29484 7 1 2 29481 29483
0 29485 5 1 1 29484
0 29486 7 1 2 51359 29485
0 29487 5 1 1 29486
0 29488 7 1 2 53534 77530
0 29489 5 1 1 29488
0 29490 7 1 2 29487 29489
0 29491 5 1 1 29490
0 29492 7 1 2 70908 29491
0 29493 5 1 1 29492
0 29494 7 1 2 29455 29493
0 29495 7 1 2 29452 29494
0 29496 7 1 2 29401 29495
0 29497 7 1 2 29339 29496
0 29498 5 1 1 29497
0 29499 7 1 2 50479 29498
0 29500 5 1 1 29499
0 29501 7 1 2 53535 77546
0 29502 5 1 1 29501
0 29503 7 1 2 75466 75486
0 29504 7 1 2 77207 29503
0 29505 5 1 1 29504
0 29506 7 1 2 29502 29505
0 29507 5 1 1 29506
0 29508 7 1 2 51078 29507
0 29509 5 1 1 29508
0 29510 7 1 2 53536 77548
0 29511 5 1 1 29510
0 29512 7 1 2 29509 29511
0 29513 5 1 1 29512
0 29514 7 1 2 51360 29513
0 29515 5 1 1 29514
0 29516 7 1 2 77599 77609
0 29517 5 1 1 29516
0 29518 7 1 2 29515 29517
0 29519 5 1 1 29518
0 29520 7 1 2 77542 29519
0 29521 5 1 1 29520
0 29522 7 1 2 77552 77613
0 29523 5 1 1 29522
0 29524 7 1 2 53537 77404
0 29525 5 1 1 29524
0 29526 7 2 2 51079 64465
0 29527 7 2 2 56225 75487
0 29528 5 1 1 77616
0 29529 7 1 2 76651 77617
0 29530 7 1 2 77614 29529
0 29531 5 1 1 29530
0 29532 7 1 2 29525 29531
0 29533 5 1 1 29532
0 29534 7 1 2 58443 29533
0 29535 5 1 1 29534
0 29536 7 1 2 53538 28320
0 29537 5 1 1 29536
0 29538 7 1 2 55702 77370
0 29539 5 1 1 29538
0 29540 7 2 2 52433 63133
0 29541 7 1 2 53227 77618
0 29542 5 1 1 29541
0 29543 7 1 2 29539 29542
0 29544 5 1 1 29543
0 29545 7 1 2 75467 75991
0 29546 7 1 2 29544 29545
0 29547 5 1 1 29546
0 29548 7 1 2 29537 29547
0 29549 7 1 2 29535 29548
0 29550 5 1 1 29549
0 29551 7 1 2 51361 29550
0 29552 5 1 1 29551
0 29553 7 1 2 29523 29552
0 29554 5 1 1 29553
0 29555 7 1 2 57241 29554
0 29556 5 1 1 29555
0 29557 7 1 2 29521 29556
0 29558 7 1 2 29500 29557
0 29559 7 1 2 29150 29558
0 29560 5 1 1 29559
0 29561 7 1 2 48770 29560
0 29562 5 1 1 29561
0 29563 7 1 2 73962 76036
0 29564 5 1 1 29563
0 29565 7 1 2 48406 76567
0 29566 5 1 1 29565
0 29567 7 1 2 77278 29566
0 29568 5 1 1 29567
0 29569 7 1 2 65936 76769
0 29570 5 1 1 29569
0 29571 7 1 2 29568 29570
0 29572 5 1 1 29571
0 29573 7 1 2 74841 26140
0 29574 5 1 1 29573
0 29575 7 1 2 52170 29574
0 29576 5 1 1 29575
0 29577 7 1 2 29576 76415
0 29578 7 1 2 29572 29577
0 29579 5 1 1 29578
0 29580 7 1 2 74192 75290
0 29581 5 1 1 29580
0 29582 7 1 2 29579 29581
0 29583 5 1 1 29582
0 29584 7 1 2 53228 29583
0 29585 5 1 1 29584
0 29586 7 1 2 60132 62018
0 29587 5 1 1 29586
0 29588 7 1 2 52171 76918
0 29589 5 1 1 29588
0 29590 7 1 2 29587 29589
0 29591 5 1 1 29590
0 29592 7 1 2 62491 65660
0 29593 7 1 2 66034 29592
0 29594 7 1 2 29591 29593
0 29595 5 1 1 29594
0 29596 7 1 2 29585 29595
0 29597 5 1 1 29596
0 29598 7 1 2 68936 29597
0 29599 5 1 1 29598
0 29600 7 2 2 62270 73400
0 29601 7 2 2 53539 77620
0 29602 7 1 2 52659 77347
0 29603 7 1 2 77622 29602
0 29604 5 1 1 29603
0 29605 7 1 2 29599 29604
0 29606 5 1 1 29605
0 29607 7 1 2 53351 29606
0 29608 5 1 1 29607
0 29609 7 1 2 70621 75502
0 29610 7 1 2 77623 29609
0 29611 5 1 1 29610
0 29612 7 1 2 29608 29611
0 29613 5 1 1 29612
0 29614 7 1 2 52543 29613
0 29615 5 1 1 29614
0 29616 7 1 2 64313 73130
0 29617 5 1 1 29616
0 29618 7 1 2 77402 77621
0 29619 5 1 1 29618
0 29620 7 1 2 29617 29619
0 29621 5 1 1 29620
0 29622 7 4 2 52660 53229
0 29623 7 1 2 76205 77624
0 29624 7 1 2 29621 29623
0 29625 5 1 1 29624
0 29626 7 1 2 29615 29625
0 29627 5 1 1 29626
0 29628 7 1 2 29564 29627
0 29629 5 1 1 29628
0 29630 7 1 2 55545 29629
0 29631 7 1 2 29562 29630
0 29632 7 1 2 28925 29631
0 29633 5 1 1 29632
0 29634 7 1 2 53230 60832
0 29635 5 1 1 29634
0 29636 7 1 2 70307 29635
0 29637 5 1 1 29636
0 29638 7 1 2 52434 29637
0 29639 5 1 1 29638
0 29640 7 1 2 71449 76644
0 29641 7 1 2 77212 29640
0 29642 5 1 1 29641
0 29643 7 1 2 29639 29642
0 29644 5 1 1 29643
0 29645 7 1 2 58039 29644
0 29646 5 1 1 29645
0 29647 7 1 2 69666 77226
0 29648 7 1 2 60827 29647
0 29649 5 1 1 29648
0 29650 7 1 2 57630 29649
0 29651 5 1 1 29650
0 29652 7 1 2 54353 60654
0 29653 5 2 1 29652
0 29654 7 1 2 59762 77628
0 29655 5 1 1 29654
0 29656 7 1 2 56369 29655
0 29657 7 2 2 63770 61705
0 29658 5 1 1 77630
0 29659 7 1 2 66647 29658
0 29660 5 1 1 29659
0 29661 7 1 2 56929 60783
0 29662 5 2 1 29661
0 29663 7 1 2 70742 77632
0 29664 5 1 1 29663
0 29665 7 1 2 29660 29664
0 29666 7 1 2 29656 29665
0 29667 7 1 2 29651 29666
0 29668 5 1 1 29667
0 29669 7 1 2 56462 29668
0 29670 5 1 1 29669
0 29671 7 1 2 55365 29670
0 29672 7 1 2 29646 29671
0 29673 5 1 1 29672
0 29674 7 1 2 53352 75602
0 29675 5 1 1 29674
0 29676 7 1 2 60212 61481
0 29677 5 1 1 29676
0 29678 7 1 2 29675 29677
0 29679 5 1 1 29678
0 29680 7 1 2 59188 29679
0 29681 5 1 1 29680
0 29682 7 1 2 48530 72486
0 29683 5 1 1 29682
0 29684 7 1 2 23356 29683
0 29685 5 1 1 29684
0 29686 7 1 2 56127 29685
0 29687 5 1 1 29686
0 29688 7 1 2 29681 29687
0 29689 5 1 1 29688
0 29690 7 1 2 55783 29689
0 29691 5 1 1 29690
0 29692 7 2 2 53353 64873
0 29693 5 1 1 77634
0 29694 7 1 2 48531 60213
0 29695 5 1 1 29694
0 29696 7 1 2 65671 75669
0 29697 5 1 1 29696
0 29698 7 1 2 29695 29697
0 29699 5 1 1 29698
0 29700 7 1 2 58615 29699
0 29701 5 1 1 29700
0 29702 7 1 2 29693 29701
0 29703 5 1 1 29702
0 29704 7 1 2 56128 29703
0 29705 5 1 1 29704
0 29706 7 1 2 53354 75132
0 29707 5 1 1 29706
0 29708 7 1 2 19285 29707
0 29709 5 1 1 29708
0 29710 7 1 2 58348 61376
0 29711 7 1 2 29709 29710
0 29712 5 1 1 29711
0 29713 7 1 2 63192 77283
0 29714 5 1 1 29713
0 29715 7 1 2 75524 29714
0 29716 7 1 2 29712 29715
0 29717 7 1 2 29705 29716
0 29718 7 1 2 58616 67582
0 29719 5 1 1 29718
0 29720 7 1 2 63037 29719
0 29721 5 1 1 29720
0 29722 7 1 2 59189 29721
0 29723 5 1 1 29722
0 29724 7 1 2 53355 29723
0 29725 5 1 1 29724
0 29726 7 1 2 48532 57943
0 29727 7 1 2 77631 29726
0 29728 7 1 2 70287 29727
0 29729 5 1 1 29728
0 29730 7 1 2 29725 29729
0 29731 5 1 1 29730
0 29732 7 1 2 60326 61391
0 29733 5 1 1 29732
0 29734 7 1 2 66239 29733
0 29735 5 1 1 29734
0 29736 7 1 2 53356 29735
0 29737 5 1 1 29736
0 29738 7 1 2 48533 74591
0 29739 5 1 1 29738
0 29740 7 1 2 29737 29739
0 29741 5 1 1 29740
0 29742 7 1 2 58309 29741
0 29743 5 1 1 29742
0 29744 7 1 2 29731 29743
0 29745 7 1 2 29717 29744
0 29746 7 1 2 29691 29745
0 29747 5 1 1 29746
0 29748 7 1 2 49479 29747
0 29749 5 1 1 29748
0 29750 7 3 2 75525 24379
0 29751 5 1 1 77636
0 29752 7 1 2 53357 77160
0 29753 5 1 1 29752
0 29754 7 1 2 77637 29753
0 29755 5 1 1 29754
0 29756 7 1 2 63945 29755
0 29757 5 1 1 29756
0 29758 7 1 2 48534 53358
0 29759 7 2 2 58403 29758
0 29760 7 1 2 71453 77639
0 29761 5 1 1 29760
0 29762 7 1 2 29757 29761
0 29763 5 1 1 29762
0 29764 7 1 2 57830 29763
0 29765 5 1 1 29764
0 29766 7 1 2 48210 58288
0 29767 5 1 1 29766
0 29768 7 1 2 76883 77413
0 29769 7 1 2 29767 29768
0 29770 5 1 1 29769
0 29771 7 1 2 56557 29770
0 29772 5 1 1 29771
0 29773 7 1 2 60214 29772
0 29774 5 1 1 29773
0 29775 7 1 2 67373 75702
0 29776 5 1 1 29775
0 29777 7 1 2 62409 29751
0 29778 5 2 1 29777
0 29779 7 1 2 60246 77641
0 29780 7 1 2 29776 29779
0 29781 5 1 1 29780
0 29782 7 1 2 29774 29781
0 29783 5 1 1 29782
0 29784 7 2 2 52544 71954
0 29785 5 1 1 77643
0 29786 7 1 2 53359 77644
0 29787 5 1 1 29786
0 29788 7 2 2 64280 29787
0 29789 7 1 2 77645 75598
0 29790 5 1 1 29789
0 29791 7 1 2 54068 61405
0 29792 7 1 2 75681 29791
0 29793 5 1 1 29792
0 29794 7 1 2 56558 72487
0 29795 5 1 1 29794
0 29796 7 1 2 29793 29795
0 29797 5 1 1 29796
0 29798 7 1 2 62438 29797
0 29799 5 1 1 29798
0 29800 7 1 2 56463 4917
0 29801 5 1 1 29800
0 29802 7 1 2 64281 60398
0 29803 5 1 1 29802
0 29804 7 1 2 49357 72488
0 29805 5 1 1 29804
0 29806 7 1 2 29803 29805
0 29807 5 1 1 29806
0 29808 7 1 2 29801 29807
0 29809 5 1 1 29808
0 29810 7 1 2 29799 29809
0 29811 7 1 2 29790 29810
0 29812 5 1 1 29811
0 29813 7 1 2 55784 29812
0 29814 5 1 1 29813
0 29815 7 1 2 74550 77135
0 29816 5 1 1 29815
0 29817 7 1 2 77638 29816
0 29818 5 1 1 29817
0 29819 7 1 2 48535 29818
0 29820 5 1 1 29819
0 29821 7 1 2 69395 77646
0 29822 5 1 1 29821
0 29823 7 1 2 51362 29822
0 29824 7 1 2 29820 29823
0 29825 7 1 2 29814 29824
0 29826 7 1 2 29783 29825
0 29827 7 1 2 29765 29826
0 29828 7 1 2 29749 29827
0 29829 5 1 1 29828
0 29830 7 1 2 54694 29829
0 29831 7 1 2 29673 29830
0 29832 5 1 1 29831
0 29833 7 3 2 67256 67213
0 29834 5 3 1 77647
0 29835 7 1 2 60645 70395
0 29836 5 1 1 29835
0 29837 7 1 2 70654 29836
0 29838 5 1 1 29837
0 29839 7 1 2 77650 29838
0 29840 5 1 1 29839
0 29841 7 1 2 61352 58906
0 29842 5 1 1 29841
0 29843 7 1 2 29840 29842
0 29844 5 1 1 29843
0 29845 7 1 2 73111 29844
0 29846 5 1 1 29845
0 29847 7 1 2 47953 77119
0 29848 5 1 1 29847
0 29849 7 1 2 20003 29848
0 29850 5 1 1 29849
0 29851 7 1 2 29850 75659
0 29852 5 1 1 29851
0 29853 7 1 2 76050 75662
0 29854 5 1 1 29853
0 29855 7 1 2 57725 29854
0 29856 5 1 1 29855
0 29857 7 1 2 29852 29856
0 29858 5 1 1 29857
0 29859 7 1 2 51363 29858
0 29860 5 1 1 29859
0 29861 7 1 2 29846 29860
0 29862 5 1 1 29861
0 29863 7 1 2 54069 29862
0 29864 5 1 1 29863
0 29865 7 1 2 60637 75660
0 29866 5 1 1 29865
0 29867 7 1 2 57364 29866
0 29868 5 1 1 29867
0 29869 7 1 2 61292 29868
0 29870 5 1 1 29869
0 29871 7 1 2 56559 68013
0 29872 5 1 1 29871
0 29873 7 1 2 48536 77285
0 29874 5 1 1 29873
0 29875 7 1 2 29872 29874
0 29876 5 1 1 29875
0 29877 7 1 2 48407 61264
0 29878 7 1 2 29876 29877
0 29879 5 1 1 29878
0 29880 7 1 2 59684 61265
0 29881 5 2 1 29880
0 29882 7 1 2 59699 77653
0 29883 5 1 1 29882
0 29884 7 1 2 57374 29883
0 29885 5 1 1 29884
0 29886 7 1 2 59054 66169
0 29887 7 1 2 29885 29886
0 29888 7 1 2 29879 29887
0 29889 7 1 2 29870 29888
0 29890 5 1 1 29889
0 29891 7 1 2 76952 77255
0 29892 5 1 1 29891
0 29893 7 1 2 23997 29892
0 29894 5 1 1 29893
0 29895 7 1 2 50480 29894
0 29896 5 1 1 29895
0 29897 7 2 2 54354 57029
0 29898 7 1 2 59943 70641
0 29899 5 1 1 29898
0 29900 7 2 2 71006 29899
0 29901 5 1 1 77657
0 29902 7 1 2 48634 77658
0 29903 5 1 1 29902
0 29904 7 1 2 77655 29903
0 29905 5 1 1 29904
0 29906 7 1 2 29896 29905
0 29907 5 1 1 29906
0 29908 7 1 2 53360 29907
0 29909 5 1 1 29908
0 29910 7 1 2 52545 77656
0 29911 7 1 2 29901 29910
0 29912 5 1 1 29911
0 29913 7 1 2 55366 29912
0 29914 7 1 2 29909 29913
0 29915 5 1 1 29914
0 29916 7 1 2 29890 29915
0 29917 5 1 1 29916
0 29918 7 1 2 29864 29917
0 29919 5 1 1 29918
0 29920 7 1 2 50806 29919
0 29921 5 1 1 29920
0 29922 7 1 2 53231 72449
0 29923 5 1 1 29922
0 29924 7 1 2 29921 29923
0 29925 7 1 2 29832 29924
0 29926 5 1 1 29925
0 29927 7 1 2 49768 29926
0 29928 5 1 1 29927
0 29929 7 1 2 58555 65870
0 29930 7 1 2 74075 71239
0 29931 7 1 2 29929 29930
0 29932 5 1 1 29931
0 29933 7 1 2 60215 63984
0 29934 7 1 2 66013 29933
0 29935 5 1 1 29934
0 29936 7 1 2 29932 29935
0 29937 5 1 1 29936
0 29938 7 1 2 48537 29937
0 29939 5 1 1 29938
0 29940 7 1 2 66618 71423
0 29941 7 1 2 59267 29940
0 29942 5 1 1 29941
0 29943 7 1 2 29939 29942
0 29944 5 1 1 29943
0 29945 7 1 2 69882 29944
0 29946 5 1 1 29945
0 29947 7 1 2 57175 77039
0 29948 5 2 1 29947
0 29949 7 1 2 7150 77659
0 29950 5 1 1 29949
0 29951 7 1 2 50807 29950
0 29952 5 1 1 29951
0 29953 7 1 2 60216 58917
0 29954 5 1 1 29953
0 29955 7 1 2 29952 29954
0 29956 5 1 1 29955
0 29957 7 1 2 56129 29956
0 29958 5 1 1 29957
0 29959 7 1 2 48211 74828
0 29960 5 2 1 29959
0 29961 7 2 2 74023 77661
0 29962 5 1 1 77663
0 29963 7 1 2 54355 72781
0 29964 5 1 1 29963
0 29965 7 2 2 77664 29964
0 29966 7 1 2 50808 77665
0 29967 5 1 1 29966
0 29968 7 1 2 57508 74076
0 29969 7 1 2 29967 29968
0 29970 5 1 1 29969
0 29971 7 1 2 29958 29970
0 29972 5 1 1 29971
0 29973 7 1 2 56930 29972
0 29974 5 1 1 29973
0 29975 7 1 2 29946 29974
0 29976 5 1 1 29975
0 29977 7 1 2 66801 29976
0 29978 5 1 1 29977
0 29979 7 1 2 29928 29978
0 29980 5 1 1 29979
0 29981 7 1 2 48771 29980
0 29982 5 1 1 29981
0 29983 7 1 2 61563 62233
0 29984 5 1 1 29983
0 29985 7 1 2 62806 62059
0 29986 5 1 1 29985
0 29987 7 1 2 29984 29986
0 29988 5 1 1 29987
0 29989 7 1 2 56370 29988
0 29990 5 1 1 29989
0 29991 7 1 2 55918 61986
0 29992 5 1 1 29991
0 29993 7 1 2 56931 29992
0 29994 5 1 1 29993
0 29995 7 1 2 63929 77351
0 29996 5 1 1 29995
0 29997 7 1 2 48635 29996
0 29998 5 1 1 29997
0 29999 7 2 2 50481 29998
0 30000 5 1 1 77667
0 30001 7 1 2 29994 77668
0 30002 7 1 2 29990 30001
0 30003 5 1 1 30002
0 30004 7 1 2 48538 61796
0 30005 5 1 1 30004
0 30006 7 1 2 64732 30005
0 30007 5 2 1 30006
0 30008 7 1 2 76557 77669
0 30009 5 1 1 30008
0 30010 7 1 2 48539 62807
0 30011 5 1 1 30010
0 30012 7 1 2 58520 60133
0 30013 5 1 1 30012
0 30014 7 1 2 62276 30013
0 30015 5 1 1 30014
0 30016 7 1 2 61564 30015
0 30017 5 1 1 30016
0 30018 7 1 2 30011 30017
0 30019 7 1 2 30009 30018
0 30020 5 1 1 30019
0 30021 7 1 2 53232 30020
0 30022 5 1 1 30021
0 30023 7 1 2 54356 28450
0 30024 7 1 2 30022 30023
0 30025 5 1 1 30024
0 30026 7 1 2 30003 30025
0 30027 5 1 1 30026
0 30028 7 1 2 50809 30027
0 30029 5 1 1 30028
0 30030 7 1 2 49480 62760
0 30031 5 1 1 30030
0 30032 7 1 2 56130 70863
0 30033 5 2 1 30032
0 30034 7 1 2 59175 57793
0 30035 5 1 1 30034
0 30036 7 1 2 54070 30035
0 30037 5 1 1 30036
0 30038 7 1 2 77671 30037
0 30039 5 1 1 30038
0 30040 7 1 2 47954 30039
0 30041 5 1 1 30040
0 30042 7 1 2 30031 30041
0 30043 5 1 1 30042
0 30044 7 1 2 55785 30043
0 30045 5 1 1 30044
0 30046 7 2 2 59693 68011
0 30047 5 1 1 77673
0 30048 7 2 2 54071 30047
0 30049 5 1 1 77675
0 30050 7 1 2 61417 30049
0 30051 5 1 1 30050
0 30052 7 1 2 61978 30051
0 30053 5 1 1 30052
0 30054 7 1 2 56131 74665
0 30055 5 1 1 30054
0 30056 7 1 2 61138 66230
0 30057 5 1 1 30056
0 30058 7 1 2 52435 57242
0 30059 5 1 1 30058
0 30060 7 1 2 49481 30059
0 30061 5 1 1 30060
0 30062 7 1 2 58563 61124
0 30063 7 1 2 30061 30062
0 30064 7 1 2 30057 30063
0 30065 7 1 2 30055 30064
0 30066 7 1 2 30053 30065
0 30067 7 1 2 30045 30066
0 30068 5 1 1 30067
0 30069 7 1 2 52546 30068
0 30070 5 1 1 30069
0 30071 7 1 2 61139 28049
0 30072 5 1 1 30071
0 30073 7 1 2 48636 30072
0 30074 5 1 1 30073
0 30075 7 1 2 66351 28961
0 30076 5 1 1 30075
0 30077 7 1 2 30074 30076
0 30078 5 1 1 30077
0 30079 7 1 2 50255 30078
0 30080 5 1 1 30079
0 30081 7 1 2 64331 70446
0 30082 5 1 1 30081
0 30083 7 1 2 77237 30082
0 30084 5 1 1 30083
0 30085 7 1 2 61248 30084
0 30086 5 1 1 30085
0 30087 7 1 2 77238 25382
0 30088 5 1 1 30087
0 30089 7 1 2 52436 30088
0 30090 5 1 1 30089
0 30091 7 1 2 65193 60819
0 30092 5 1 1 30091
0 30093 7 1 2 48637 30092
0 30094 5 1 1 30093
0 30095 7 1 2 30090 30094
0 30096 7 1 2 30086 30095
0 30097 5 1 1 30096
0 30098 7 1 2 57631 30097
0 30099 5 1 1 30098
0 30100 7 4 2 70694 70300
0 30101 5 1 1 77677
0 30102 7 1 2 64332 77678
0 30103 5 1 1 30102
0 30104 7 1 2 48638 66352
0 30105 5 1 1 30104
0 30106 7 1 2 30103 30105
0 30107 5 1 1 30106
0 30108 7 1 2 51964 30107
0 30109 5 1 1 30108
0 30110 7 1 2 48540 60784
0 30111 5 3 1 30110
0 30112 7 1 2 50256 77236
0 30113 5 1 1 30112
0 30114 7 1 2 49482 74874
0 30115 5 1 1 30114
0 30116 7 1 2 30113 30115
0 30117 5 1 1 30116
0 30118 7 1 2 77681 30117
0 30119 5 1 1 30118
0 30120 7 1 2 49483 63771
0 30121 5 1 1 30120
0 30122 7 1 2 48639 30121
0 30123 5 1 1 30122
0 30124 7 2 2 63183 75914
0 30125 5 1 1 77684
0 30126 7 1 2 52172 77685
0 30127 5 1 1 30126
0 30128 7 1 2 30123 30127
0 30129 5 1 1 30128
0 30130 7 1 2 58537 30129
0 30131 5 1 1 30130
0 30132 7 1 2 54695 30131
0 30133 7 1 2 30119 30132
0 30134 7 1 2 30109 30133
0 30135 7 1 2 30099 30134
0 30136 7 1 2 30080 30135
0 30137 7 1 2 30070 30136
0 30138 5 1 1 30137
0 30139 7 1 2 30029 30138
0 30140 5 1 1 30139
0 30141 7 1 2 61172 62271
0 30142 5 1 1 30141
0 30143 7 1 2 61565 30142
0 30144 5 1 1 30143
0 30145 7 2 2 47955 61797
0 30146 5 1 1 77686
0 30147 7 1 2 62060 77687
0 30148 5 1 1 30147
0 30149 7 1 2 52437 62796
0 30150 7 1 2 30148 30149
0 30151 7 1 2 30144 30150
0 30152 5 1 1 30151
0 30153 7 1 2 54357 77292
0 30154 7 1 2 30152 30153
0 30155 5 1 1 30154
0 30156 7 1 2 30140 30155
0 30157 5 1 1 30156
0 30158 7 1 2 49595 30157
0 30159 5 1 1 30158
0 30160 7 1 2 53124 61808
0 30161 5 1 1 30160
0 30162 7 1 2 67214 30161
0 30163 5 1 1 30162
0 30164 7 2 2 65170 60058
0 30165 5 1 1 77688
0 30166 7 1 2 52547 30165
0 30167 5 3 1 30166
0 30168 7 1 2 57831 77690
0 30169 5 1 1 30168
0 30170 7 1 2 30163 30169
0 30171 5 1 1 30170
0 30172 7 1 2 48408 30171
0 30173 5 1 1 30172
0 30174 7 1 2 67215 74720
0 30175 5 1 1 30174
0 30176 7 1 2 57324 30175
0 30177 7 1 2 30173 30176
0 30178 5 1 1 30177
0 30179 7 1 2 54696 30178
0 30180 5 1 1 30179
0 30181 7 2 2 48409 64874
0 30182 5 1 1 77693
0 30183 7 1 2 77691 77694
0 30184 5 1 1 30183
0 30185 7 1 2 30180 30184
0 30186 5 1 1 30185
0 30187 7 1 2 48212 30186
0 30188 5 1 1 30187
0 30189 7 1 2 57509 67216
0 30190 5 1 1 30189
0 30191 7 2 2 57325 30190
0 30192 5 4 1 77695
0 30193 7 1 2 72075 77697
0 30194 5 1 1 30193
0 30195 7 1 2 53361 30194
0 30196 7 1 2 30188 30195
0 30197 5 1 1 30196
0 30198 7 1 2 48213 77670
0 30199 5 1 1 30198
0 30200 7 1 2 58521 61566
0 30201 5 1 1 30200
0 30202 7 1 2 30199 30201
0 30203 5 1 1 30202
0 30204 7 1 2 62361 30203
0 30205 5 1 1 30204
0 30206 7 2 2 61868 62669
0 30207 5 1 1 77701
0 30208 7 1 2 77293 30207
0 30209 5 1 1 30208
0 30210 7 1 2 30205 30209
0 30211 5 1 1 30210
0 30212 7 1 2 54358 30211
0 30213 5 1 1 30212
0 30214 7 1 2 56371 62621
0 30215 5 1 1 30214
0 30216 7 1 2 67200 30215
0 30217 5 1 1 30216
0 30218 7 1 2 47956 60544
0 30219 7 1 2 30217 30218
0 30220 5 1 1 30219
0 30221 7 1 2 49596 30220
0 30222 7 1 2 30213 30221
0 30223 5 1 1 30222
0 30224 7 1 2 30197 30223
0 30225 5 1 1 30224
0 30226 7 1 2 74310 76164
0 30227 7 1 2 77689 30226
0 30228 5 1 1 30227
0 30229 7 1 2 30225 30228
0 30230 5 1 1 30229
0 30231 7 1 2 55786 30230
0 30232 5 1 1 30231
0 30233 7 1 2 58581 60134
0 30234 5 1 1 30233
0 30235 7 1 2 59224 62267
0 30236 5 1 1 30235
0 30237 7 1 2 64005 62061
0 30238 5 2 1 30237
0 30239 7 1 2 30236 77703
0 30240 7 1 2 30234 30239
0 30241 5 1 1 30240
0 30242 7 1 2 54359 30241
0 30243 5 1 1 30242
0 30244 7 1 2 48214 62248
0 30245 5 1 1 30244
0 30246 7 1 2 30243 30245
0 30247 5 1 1 30246
0 30248 7 1 2 53362 30247
0 30249 5 1 1 30248
0 30250 7 1 2 57030 1464
0 30251 5 1 1 30250
0 30252 7 1 2 56372 60545
0 30253 7 1 2 30251 30252
0 30254 5 1 1 30253
0 30255 7 1 2 30249 30254
0 30256 5 1 1 30255
0 30257 7 1 2 48640 30256
0 30258 5 1 1 30257
0 30259 7 2 2 59549 60546
0 30260 5 1 1 77705
0 30261 7 1 2 23347 30260
0 30262 5 1 1 30261
0 30263 7 2 2 56132 57304
0 30264 5 1 1 77707
0 30265 7 1 2 30262 77708
0 30266 5 1 1 30265
0 30267 7 1 2 57744 75682
0 30268 7 1 2 77438 30267
0 30269 5 1 1 30268
0 30270 7 1 2 30266 30269
0 30271 5 1 1 30270
0 30272 7 1 2 55787 30271
0 30273 5 1 1 30272
0 30274 7 1 2 48215 74210
0 30275 5 1 1 30274
0 30276 7 1 2 77704 30275
0 30277 5 1 1 30276
0 30278 7 1 2 54360 30277
0 30279 5 1 1 30278
0 30280 7 1 2 67246 30279
0 30281 5 1 1 30280
0 30282 7 1 2 77243 30281
0 30283 5 1 1 30282
0 30284 7 1 2 30273 30283
0 30285 7 1 2 30258 30284
0 30286 5 1 1 30285
0 30287 7 1 2 61567 30286
0 30288 5 1 1 30287
0 30289 7 1 2 58690 76996
0 30290 5 1 1 30289
0 30291 7 1 2 56373 67431
0 30292 5 1 1 30291
0 30293 7 1 2 30290 30292
0 30294 5 1 1 30293
0 30295 7 1 2 53363 30294
0 30296 5 1 1 30295
0 30297 7 2 2 48216 75683
0 30298 7 1 2 67106 77709
0 30299 5 1 1 30298
0 30300 7 2 2 48410 60547
0 30301 5 1 1 77711
0 30302 7 1 2 61159 77712
0 30303 5 1 1 30302
0 30304 7 1 2 30299 30303
0 30305 5 1 1 30304
0 30306 7 1 2 55788 30305
0 30307 5 1 1 30306
0 30308 7 1 2 47957 75684
0 30309 5 1 1 30308
0 30310 7 1 2 30301 30309
0 30311 5 1 1 30310
0 30312 7 1 2 56374 62062
0 30313 7 1 2 30311 30312
0 30314 5 1 1 30313
0 30315 7 1 2 30307 30314
0 30316 7 1 2 30296 30315
0 30317 5 1 1 30316
0 30318 7 1 2 48641 30317
0 30319 5 1 1 30318
0 30320 7 1 2 52316 75396
0 30321 5 1 1 30320
0 30322 7 1 2 62137 77635
0 30323 7 1 2 30321 30322
0 30324 5 1 1 30323
0 30325 7 1 2 30319 30324
0 30326 5 1 1 30325
0 30327 7 1 2 62306 30326
0 30328 5 1 1 30327
0 30329 7 1 2 64267 76937
0 30330 5 1 1 30329
0 30331 7 1 2 58404 69006
0 30332 7 1 2 75666 30331
0 30333 5 1 1 30332
0 30334 7 1 2 30330 30333
0 30335 5 1 1 30334
0 30336 7 1 2 56133 30335
0 30337 5 1 1 30336
0 30338 7 1 2 59485 30182
0 30339 5 1 1 30338
0 30340 7 1 2 72370 30339
0 30341 5 1 1 30340
0 30342 7 2 2 54697 67217
0 30343 5 1 1 77713
0 30344 7 1 2 57774 66704
0 30345 5 1 1 30344
0 30346 7 1 2 30343 30345
0 30347 5 1 1 30346
0 30348 7 1 2 61717 30347
0 30349 5 1 1 30348
0 30350 7 1 2 30341 30349
0 30351 5 1 1 30350
0 30352 7 1 2 53364 30351
0 30353 5 1 1 30352
0 30354 7 1 2 48642 58491
0 30355 7 1 2 63590 30354
0 30356 5 1 1 30355
0 30357 7 1 2 30353 30356
0 30358 5 1 1 30357
0 30359 7 1 2 62063 30358
0 30360 5 1 1 30359
0 30361 7 1 2 30337 30360
0 30362 7 1 2 30328 30361
0 30363 7 1 2 53365 74425
0 30364 5 1 1 30363
0 30365 7 1 2 50482 76165
0 30366 5 1 1 30365
0 30367 7 1 2 30364 30366
0 30368 5 1 1 30367
0 30369 7 1 2 58509 30368
0 30370 5 1 1 30369
0 30371 7 1 2 63378 77710
0 30372 5 1 1 30371
0 30373 7 1 2 30370 30372
0 30374 5 1 1 30373
0 30375 7 1 2 55789 30374
0 30376 5 1 1 30375
0 30377 7 1 2 48541 60548
0 30378 5 1 1 30377
0 30379 7 1 2 53366 58188
0 30380 5 1 1 30379
0 30381 7 1 2 30378 30380
0 30382 5 1 1 30381
0 30383 7 1 2 62064 30382
0 30384 5 1 1 30383
0 30385 7 1 2 64877 58336
0 30386 5 1 1 30385
0 30387 7 1 2 53367 30386
0 30388 5 1 1 30387
0 30389 7 1 2 30384 30388
0 30390 5 1 1 30389
0 30391 7 1 2 48643 30390
0 30392 5 1 1 30391
0 30393 7 1 2 74426 77640
0 30394 5 1 1 30393
0 30395 7 1 2 30392 30394
0 30396 7 1 2 30376 30395
0 30397 5 1 1 30396
0 30398 7 1 2 77012 30397
0 30399 5 1 1 30398
0 30400 7 1 2 74792 75563
0 30401 5 1 1 30400
0 30402 7 1 2 60360 71407
0 30403 5 1 1 30402
0 30404 7 1 2 77698 30403
0 30405 5 1 1 30404
0 30406 7 1 2 48542 58329
0 30407 5 1 1 30406
0 30408 7 1 2 58405 74716
0 30409 5 1 1 30408
0 30410 7 1 2 30407 30409
0 30411 5 1 1 30410
0 30412 7 1 2 77692 30411
0 30413 5 1 1 30412
0 30414 7 1 2 64354 30413
0 30415 7 1 2 30405 30414
0 30416 5 1 1 30415
0 30417 7 1 2 54698 30416
0 30418 5 1 1 30417
0 30419 7 1 2 30401 30418
0 30420 5 1 1 30419
0 30421 7 1 2 53368 30420
0 30422 5 1 1 30421
0 30423 7 1 2 30399 30422
0 30424 7 1 2 30362 30423
0 30425 7 1 2 30288 30424
0 30426 7 1 2 30232 30425
0 30427 7 1 2 30159 30426
0 30428 5 1 1 30427
0 30429 7 1 2 55367 30428
0 30430 5 1 1 30429
0 30431 7 1 2 55919 61999
0 30432 5 1 1 30431
0 30433 7 1 2 56932 30432
0 30434 5 1 1 30433
0 30435 7 1 2 61568 62245
0 30436 5 1 1 30435
0 30437 7 1 2 62808 76568
0 30438 5 1 1 30437
0 30439 7 1 2 64733 30438
0 30440 7 1 2 30436 30439
0 30441 5 1 1 30440
0 30442 7 1 2 56375 30441
0 30443 5 1 1 30442
0 30444 7 1 2 30434 30443
0 30445 5 1 1 30444
0 30446 7 1 2 54361 30445
0 30447 5 1 1 30446
0 30448 7 1 2 58942 76139
0 30449 5 1 1 30448
0 30450 7 1 2 66648 30449
0 30451 5 2 1 30450
0 30452 7 1 2 54072 77715
0 30453 5 1 1 30452
0 30454 7 1 2 30447 30453
0 30455 5 1 1 30454
0 30456 7 1 2 57944 68701
0 30457 7 1 2 30455 30456
0 30458 5 1 1 30457
0 30459 7 1 2 30430 30458
0 30460 5 1 1 30459
0 30461 7 1 2 75291 30460
0 30462 5 1 1 30461
0 30463 7 2 2 54362 75204
0 30464 5 2 1 77717
0 30465 7 1 2 73840 77718
0 30466 5 1 1 30465
0 30467 7 1 2 67530 70533
0 30468 5 3 1 30467
0 30469 7 1 2 30466 77721
0 30470 5 1 1 30469
0 30471 7 1 2 56750 30470
0 30472 5 1 1 30471
0 30473 7 1 2 50483 77166
0 30474 5 1 1 30473
0 30475 7 1 2 57176 76416
0 30476 7 1 2 30474 30475
0 30477 5 1 1 30476
0 30478 7 1 2 30472 30477
0 30479 5 1 1 30478
0 30480 7 1 2 54699 30479
0 30481 5 1 1 30480
0 30482 7 1 2 73154 77174
0 30483 5 1 1 30482
0 30484 7 1 2 30481 30483
0 30485 5 1 1 30484
0 30486 7 1 2 56134 30485
0 30487 5 1 1 30486
0 30488 7 1 2 60697 68096
0 30489 5 1 1 30488
0 30490 7 1 2 57243 76856
0 30491 7 1 2 61676 30490
0 30492 7 4 2 30489 30491
0 30493 5 1 1 77724
0 30494 7 1 2 50484 77725
0 30495 5 1 1 30494
0 30496 7 1 2 73841 30495
0 30497 5 1 1 30496
0 30498 7 1 2 77722 30497
0 30499 5 1 1 30498
0 30500 7 1 2 54700 30499
0 30501 5 1 1 30500
0 30502 7 1 2 50485 76560
0 30503 5 1 1 30502
0 30504 7 1 2 61569 30503
0 30505 5 1 1 30504
0 30506 7 1 2 54363 70755
0 30507 5 1 1 30506
0 30508 7 1 2 74812 30507
0 30509 7 1 2 30505 30508
0 30510 5 1 1 30509
0 30511 7 1 2 73155 30510
0 30512 5 1 1 30511
0 30513 7 1 2 76569 76520
0 30514 5 1 1 30513
0 30515 7 1 2 62115 73156
0 30516 5 1 1 30515
0 30517 7 1 2 30514 30516
0 30518 5 1 1 30517
0 30519 7 1 2 61757 30518
0 30520 5 1 1 30519
0 30521 7 1 2 65029 61954
0 30522 7 1 2 76417 30521
0 30523 5 1 1 30522
0 30524 7 1 2 30520 30523
0 30525 7 1 2 30512 30524
0 30526 7 1 2 30501 30525
0 30527 5 1 1 30526
0 30528 7 1 2 57510 30527
0 30529 5 1 1 30528
0 30530 7 1 2 30487 30529
0 30531 5 1 1 30530
0 30532 7 1 2 56933 30531
0 30533 5 1 1 30532
0 30534 7 1 2 66649 68173
0 30535 5 2 1 30534
0 30536 7 1 2 60399 76418
0 30537 5 1 1 30536
0 30538 7 1 2 77723 30537
0 30539 5 1 1 30538
0 30540 7 1 2 62183 30539
0 30541 7 1 2 77728 30540
0 30542 5 1 1 30541
0 30543 7 1 2 30533 30542
0 30544 5 1 1 30543
0 30545 7 1 2 57945 30544
0 30546 5 1 1 30545
0 30547 7 5 2 49597 75292
0 30548 7 1 2 54364 76697
0 30549 5 1 1 30548
0 30550 7 8 2 50486 60666
0 30551 5 2 1 77735
0 30552 7 1 2 48644 77736
0 30553 5 1 1 30552
0 30554 7 1 2 30549 30553
0 30555 5 1 1 30554
0 30556 7 1 2 57632 30555
0 30557 5 1 1 30556
0 30558 7 1 2 23518 76625
0 30559 7 1 2 58538 30558
0 30560 7 1 2 65804 30559
0 30561 5 1 1 30560
0 30562 7 1 2 30557 30561
0 30563 5 1 1 30562
0 30564 7 1 2 77730 30563
0 30565 5 1 1 30564
0 30566 7 1 2 62918 70133
0 30567 7 1 2 60675 30566
0 30568 5 1 1 30567
0 30569 7 2 2 75488 75480
0 30570 5 1 1 77745
0 30571 7 2 2 49598 77378
0 30572 5 1 1 77747
0 30573 7 1 2 75293 77748
0 30574 5 1 1 30573
0 30575 7 1 2 30570 30574
0 30576 5 1 1 30575
0 30577 7 1 2 57031 63499
0 30578 7 1 2 30576 30577
0 30579 5 1 1 30578
0 30580 7 1 2 30568 30579
0 30581 7 1 2 30565 30580
0 30582 5 1 1 30581
0 30583 7 1 2 55368 30582
0 30584 5 1 1 30583
0 30585 7 1 2 64278 76534
0 30586 7 1 2 63500 30585
0 30587 5 1 1 30586
0 30588 7 1 2 30584 30587
0 30589 5 1 1 30588
0 30590 7 1 2 54701 30589
0 30591 5 1 1 30590
0 30592 7 2 2 63297 64099
0 30593 5 2 1 77749
0 30594 7 1 2 62919 77750
0 30595 5 1 1 30594
0 30596 7 1 2 48645 77731
0 30597 5 1 1 30596
0 30598 7 1 2 30595 30597
0 30599 5 2 1 30598
0 30600 7 1 2 60856 77753
0 30601 5 1 1 30600
0 30602 7 2 2 58040 70949
0 30603 7 1 2 62920 77360
0 30604 7 1 2 77755 30603
0 30605 5 1 1 30604
0 30606 7 1 2 30601 30605
0 30607 5 1 1 30606
0 30608 7 1 2 54365 30607
0 30609 5 1 1 30608
0 30610 7 1 2 70950 76115
0 30611 5 1 1 30610
0 30612 7 2 2 58539 76618
0 30613 7 1 2 70447 77757
0 30614 5 1 1 30613
0 30615 7 1 2 30611 30614
0 30616 5 1 1 30615
0 30617 7 1 2 70534 76253
0 30618 7 1 2 30616 30617
0 30619 5 1 1 30618
0 30620 7 1 2 30609 30619
0 30621 5 1 1 30620
0 30622 7 1 2 63785 30621
0 30623 5 1 1 30622
0 30624 7 1 2 30591 30623
0 30625 5 1 1 30624
0 30626 7 1 2 57244 30625
0 30627 5 1 1 30626
0 30628 7 1 2 62144 60573
0 30629 7 2 2 62290 30628
0 30630 7 1 2 48646 77759
0 30631 5 1 1 30630
0 30632 7 1 2 76892 75626
0 30633 7 1 2 77591 30632
0 30634 5 1 1 30633
0 30635 7 1 2 30631 30634
0 30636 5 1 1 30635
0 30637 7 1 2 77732 30636
0 30638 5 1 1 30637
0 30639 7 1 2 77592 76396
0 30640 5 1 1 30639
0 30641 7 1 2 76943 30640
0 30642 5 1 1 30641
0 30643 7 1 2 52438 30642
0 30644 5 1 1 30643
0 30645 7 1 2 53369 77760
0 30646 5 1 1 30645
0 30647 7 1 2 30644 30646
0 30648 5 1 1 30647
0 30649 7 1 2 52548 30648
0 30650 5 1 1 30649
0 30651 7 1 2 72988 75685
0 30652 5 1 1 30651
0 30653 7 1 2 30650 30652
0 30654 5 1 1 30653
0 30655 7 1 2 62921 30654
0 30656 5 1 1 30655
0 30657 7 1 2 30638 30656
0 30658 5 1 1 30657
0 30659 7 1 2 55369 30658
0 30660 5 1 1 30659
0 30661 7 1 2 67968 74251
0 30662 7 1 2 76955 30661
0 30663 5 1 1 30662
0 30664 7 1 2 30660 30663
0 30665 5 1 1 30664
0 30666 7 1 2 60893 30665
0 30667 5 1 1 30666
0 30668 7 1 2 30627 30667
0 30669 7 1 2 30546 30668
0 30670 7 1 2 30462 30669
0 30671 7 1 2 29982 30670
0 30672 5 1 1 30671
0 30673 7 1 2 55050 30672
0 30674 5 1 1 30673
0 30675 7 2 2 59294 65672
0 30676 5 1 1 77761
0 30677 7 1 2 23449 30676
0 30678 5 1 1 30677
0 30679 7 1 2 47958 30678
0 30680 5 1 1 30679
0 30681 7 1 2 56376 77176
0 30682 5 1 1 30681
0 30683 7 2 2 30680 30682
0 30684 5 1 1 77763
0 30685 7 1 2 55790 30684
0 30686 5 1 1 30685
0 30687 7 1 2 58582 59996
0 30688 5 2 1 30687
0 30689 7 1 2 60305 61203
0 30690 5 1 1 30689
0 30691 7 1 2 77765 30690
0 30692 5 1 1 30691
0 30693 7 1 2 58617 30692
0 30694 5 1 1 30693
0 30695 7 1 2 61380 77158
0 30696 5 1 1 30695
0 30697 7 1 2 56377 65419
0 30698 5 1 1 30697
0 30699 7 1 2 58173 62327
0 30700 5 2 1 30699
0 30701 7 1 2 30698 77767
0 30702 5 1 1 30701
0 30703 7 1 2 58310 30702
0 30704 5 1 1 30703
0 30705 7 1 2 50810 62462
0 30706 7 1 2 30704 30705
0 30707 7 1 2 30696 30706
0 30708 7 1 2 30694 30707
0 30709 7 1 2 30686 30708
0 30710 5 1 1 30709
0 30711 7 1 2 60837 59268
0 30712 5 1 1 30711
0 30713 7 1 2 52439 30712
0 30714 5 1 1 30713
0 30715 7 1 2 49484 30714
0 30716 7 1 2 75372 30715
0 30717 5 1 1 30716
0 30718 7 1 2 77589 30717
0 30719 5 1 1 30718
0 30720 7 1 2 62390 76767
0 30721 5 1 1 30720
0 30722 7 1 2 54073 30721
0 30723 5 1 1 30722
0 30724 7 1 2 52440 30723
0 30725 5 1 1 30724
0 30726 7 1 2 52549 30725
0 30727 5 1 1 30726
0 30728 7 1 2 54366 30727
0 30729 7 1 2 30719 30728
0 30730 5 1 1 30729
0 30731 7 1 2 57511 60655
0 30732 5 5 1 30731
0 30733 7 1 2 57245 77769
0 30734 5 1 1 30733
0 30735 7 1 2 58556 70827
0 30736 7 1 2 30734 30735
0 30737 5 1 1 30736
0 30738 7 1 2 54074 30737
0 30739 7 1 2 77582 30738
0 30740 5 1 1 30739
0 30741 7 1 2 50487 23950
0 30742 7 1 2 30740 30741
0 30743 5 1 1 30742
0 30744 7 1 2 30730 30743
0 30745 5 1 1 30744
0 30746 7 1 2 77109 77294
0 30747 5 1 1 30746
0 30748 7 1 2 54702 30747
0 30749 7 1 2 30745 30748
0 30750 5 1 1 30749
0 30751 7 1 2 30710 30750
0 30752 5 1 1 30751
0 30753 7 1 2 48543 77295
0 30754 5 1 1 30753
0 30755 7 1 2 53370 30754
0 30756 7 1 2 30752 30755
0 30757 5 1 1 30756
0 30758 7 1 2 55920 77125
0 30759 5 1 1 30758
0 30760 7 1 2 70960 30759
0 30761 5 1 1 30760
0 30762 7 1 2 64954 30761
0 30763 5 1 1 30762
0 30764 7 1 2 66358 30763
0 30765 5 1 1 30764
0 30766 7 1 2 30765 77770
0 30767 5 1 1 30766
0 30768 7 1 2 65301 2031
0 30769 5 1 1 30768
0 30770 7 1 2 52317 30769
0 30771 5 1 1 30770
0 30772 7 1 2 53125 65297
0 30773 5 2 1 30772
0 30774 7 1 2 60574 77774
0 30775 7 1 2 30771 30774
0 30776 5 1 1 30775
0 30777 7 1 2 51965 30776
0 30778 5 1 1 30777
0 30779 7 1 2 71624 30778
0 30780 7 1 2 30767 30779
0 30781 5 1 1 30780
0 30782 7 1 2 57246 30781
0 30783 5 1 1 30782
0 30784 7 1 2 53233 60725
0 30785 5 1 1 30784
0 30786 7 1 2 63630 30785
0 30787 5 1 1 30786
0 30788 7 1 2 51966 30787
0 30789 5 1 1 30788
0 30790 7 1 2 60575 30789
0 30791 5 2 1 30790
0 30792 7 1 2 70396 77776
0 30793 5 1 1 30792
0 30794 7 1 2 55921 60736
0 30795 5 1 1 30794
0 30796 7 1 2 60857 77126
0 30797 7 2 2 75733 30796
0 30798 5 1 1 77778
0 30799 7 1 2 54703 30798
0 30800 7 1 2 30795 30799
0 30801 5 1 1 30800
0 30802 7 1 2 77259 30801
0 30803 5 1 1 30802
0 30804 7 1 2 61509 65302
0 30805 5 4 1 30804
0 30806 7 1 2 55703 77780
0 30807 5 2 1 30806
0 30808 7 1 2 77784 77775
0 30809 5 1 1 30808
0 30810 7 1 2 50488 30809
0 30811 5 1 1 30810
0 30812 7 1 2 65224 71625
0 30813 5 1 1 30812
0 30814 7 1 2 52318 30813
0 30815 5 1 1 30814
0 30816 7 1 2 72801 77127
0 30817 5 1 1 30816
0 30818 7 1 2 55791 61860
0 30819 5 1 1 30818
0 30820 7 1 2 52550 30819
0 30821 5 1 1 30820
0 30822 7 1 2 30817 30821
0 30823 7 1 2 30815 30822
0 30824 7 1 2 30811 30823
0 30825 7 1 2 30803 30824
0 30826 7 1 2 30793 30825
0 30827 7 1 2 30783 30826
0 30828 5 1 1 30827
0 30829 7 1 2 52441 30828
0 30830 5 1 1 30829
0 30831 7 1 2 55922 77777
0 30832 5 1 1 30831
0 30833 7 1 2 63631 77785
0 30834 5 1 1 30833
0 30835 7 1 2 50489 30834
0 30836 5 1 1 30835
0 30837 7 1 2 52551 60858
0 30838 5 1 1 30837
0 30839 7 1 2 62373 30838
0 30840 7 1 2 30836 30839
0 30841 5 1 1 30840
0 30842 7 1 2 57633 30841
0 30843 5 1 1 30842
0 30844 7 1 2 30832 30843
0 30845 5 1 1 30844
0 30846 7 1 2 56639 30845
0 30847 5 1 1 30846
0 30848 7 1 2 52552 65805
0 30849 5 1 1 30848
0 30850 7 1 2 50811 77779
0 30851 5 1 1 30850
0 30852 7 1 2 30849 30851
0 30853 5 1 1 30852
0 30854 7 1 2 57634 30853
0 30855 5 1 1 30854
0 30856 7 3 2 48647 71626
0 30857 5 1 1 77786
0 30858 7 2 2 55923 30857
0 30859 5 1 1 77789
0 30860 7 2 2 66041 72755
0 30861 5 1 1 77791
0 30862 7 1 2 30861 24027
0 30863 5 1 1 30862
0 30864 7 1 2 60493 30863
0 30865 5 1 1 30864
0 30866 7 1 2 60726 67435
0 30867 5 1 1 30866
0 30868 7 1 2 30865 30867
0 30869 5 1 1 30868
0 30870 7 1 2 51967 30869
0 30871 5 1 1 30870
0 30872 7 1 2 30859 30871
0 30873 7 1 2 30855 30872
0 30874 5 1 1 30873
0 30875 7 1 2 57247 30874
0 30876 5 1 1 30875
0 30877 7 1 2 52553 60727
0 30878 5 1 1 30877
0 30879 7 1 2 76518 30878
0 30880 5 1 1 30879
0 30881 7 1 2 51968 30880
0 30882 5 1 1 30881
0 30883 7 1 2 72982 30882
0 30884 5 1 1 30883
0 30885 7 1 2 70397 30884
0 30886 5 1 1 30885
0 30887 7 1 2 60683 77792
0 30888 5 1 1 30887
0 30889 7 1 2 58564 71035
0 30890 5 1 1 30889
0 30891 7 1 2 30888 30890
0 30892 5 1 1 30891
0 30893 7 1 2 50490 30892
0 30894 5 1 1 30893
0 30895 7 1 2 71248 75949
0 30896 5 1 1 30895
0 30897 7 1 2 60422 30896
0 30898 5 1 1 30897
0 30899 7 2 2 52554 55704
0 30900 5 2 1 77793
0 30901 7 1 2 62374 77795
0 30902 5 1 1 30901
0 30903 7 1 2 55924 30902
0 30904 5 1 1 30903
0 30905 7 1 2 49599 30904
0 30906 7 1 2 30898 30905
0 30907 7 1 2 30894 30906
0 30908 7 1 2 30886 30907
0 30909 7 1 2 30876 30908
0 30910 7 1 2 30847 30909
0 30911 7 1 2 30830 30910
0 30912 5 1 1 30911
0 30913 7 1 2 51080 30912
0 30914 7 1 2 30757 30913
0 30915 5 1 1 30914
0 30916 7 2 2 54704 14978
0 30917 5 2 1 77797
0 30918 7 1 2 50257 63104
0 30919 5 1 1 30918
0 30920 7 1 2 48544 30919
0 30921 5 1 1 30920
0 30922 7 1 2 50491 30921
0 30923 5 1 1 30922
0 30924 7 1 2 77798 30923
0 30925 5 1 1 30924
0 30926 7 1 2 51081 30925
0 30927 5 1 1 30926
0 30928 7 1 2 59866 75081
0 30929 5 1 1 30928
0 30930 7 1 2 65446 70988
0 30931 5 1 1 30930
0 30932 7 1 2 739 30931
0 30933 7 1 2 30929 30932
0 30934 5 1 1 30933
0 30935 7 1 2 53234 30934
0 30936 5 1 1 30935
0 30937 7 1 2 30927 30936
0 30938 5 1 1 30937
0 30939 7 1 2 75764 30938
0 30940 5 1 1 30939
0 30941 7 1 2 48648 60516
0 30942 5 2 1 30941
0 30943 7 1 2 57032 75231
0 30944 5 1 1 30943
0 30945 7 1 2 77801 30944
0 30946 5 1 1 30945
0 30947 7 1 2 57635 75140
0 30948 7 1 2 30946 30947
0 30949 5 1 1 30948
0 30950 7 1 2 70157 71249
0 30951 5 1 1 30950
0 30952 7 2 2 63614 75376
0 30953 7 1 2 61472 77803
0 30954 7 1 2 30951 30953
0 30955 5 1 1 30954
0 30956 7 1 2 30949 30955
0 30957 7 1 2 30940 30956
0 30958 7 1 2 30915 30957
0 30959 5 1 1 30958
0 30960 7 1 2 55370 30959
0 30961 5 1 1 30960
0 30962 7 1 2 50492 77162
0 30963 5 1 1 30962
0 30964 7 1 2 49358 30963
0 30965 5 1 1 30964
0 30966 7 1 2 65915 30965
0 30967 5 1 1 30966
0 30968 7 1 2 48411 30967
0 30969 5 1 1 30968
0 30970 7 1 2 77188 30969
0 30971 5 1 1 30970
0 30972 7 1 2 54705 30971
0 30973 5 1 1 30972
0 30974 7 2 2 60059 58137
0 30975 5 2 1 77805
0 30976 7 1 2 58214 77807
0 30977 5 1 1 30976
0 30978 7 1 2 54367 30977
0 30979 5 1 1 30978
0 30980 7 1 2 54706 60698
0 30981 7 1 2 60077 30980
0 30982 5 1 1 30981
0 30983 7 1 2 30979 30982
0 30984 5 1 1 30983
0 30985 7 1 2 49125 30984
0 30986 5 1 1 30985
0 30987 7 2 2 54707 68165
0 30988 5 2 1 77809
0 30989 7 1 2 65255 59644
0 30990 5 1 1 30989
0 30991 7 1 2 61758 30990
0 30992 5 1 1 30991
0 30993 7 1 2 77811 30992
0 30994 5 2 1 30993
0 30995 7 1 2 48217 77813
0 30996 5 1 1 30995
0 30997 7 2 2 54708 61673
0 30998 5 1 1 77815
0 30999 7 1 2 49359 77816
0 31000 5 1 1 30999
0 31001 7 1 2 30996 31000
0 31002 7 1 2 30986 31001
0 31003 5 1 1 31002
0 31004 7 1 2 47959 31003
0 31005 5 1 1 31004
0 31006 7 1 2 49360 65030
0 31007 5 1 1 31006
0 31008 7 1 2 74086 31007
0 31009 5 1 1 31008
0 31010 7 1 2 61570 31009
0 31011 5 1 1 31010
0 31012 7 1 2 49126 77814
0 31013 5 1 1 31012
0 31014 7 1 2 59529 72077
0 31015 5 1 1 31014
0 31016 7 1 2 31013 31015
0 31017 7 1 2 31011 31016
0 31018 5 1 1 31017
0 31019 7 1 2 48218 31018
0 31020 5 1 1 31019
0 31021 7 1 2 61646 74855
0 31022 5 1 1 31021
0 31023 7 1 2 31020 31022
0 31024 7 1 2 31005 31023
0 31025 5 1 1 31024
0 31026 7 1 2 48412 31025
0 31027 5 1 1 31026
0 31028 7 1 2 30973 31027
0 31029 5 2 1 31028
0 31030 7 1 2 56378 77817
0 31031 5 1 1 31030
0 31032 7 1 2 54709 74732
0 31033 5 1 1 31032
0 31034 7 1 2 49485 77151
0 31035 5 1 1 31034
0 31036 7 1 2 31033 31035
0 31037 5 1 1 31036
0 31038 7 1 2 54075 31037
0 31039 5 1 1 31038
0 31040 7 1 2 56934 62459
0 31041 5 1 1 31040
0 31042 7 1 2 31039 31041
0 31043 5 1 1 31042
0 31044 7 1 2 47960 31043
0 31045 5 1 1 31044
0 31046 7 1 2 54368 62694
0 31047 5 1 1 31046
0 31048 7 2 2 23016 31047
0 31049 5 1 1 77819
0 31050 7 1 2 56935 31049
0 31051 5 1 1 31050
0 31052 7 1 2 31045 31051
0 31053 5 1 1 31052
0 31054 7 1 2 55792 31053
0 31055 5 1 1 31054
0 31056 7 1 2 56640 62859
0 31057 5 1 1 31056
0 31058 7 1 2 59997 31057
0 31059 5 1 1 31058
0 31060 7 1 2 57248 31059
0 31061 5 1 1 31060
0 31062 7 1 2 60903 31061
0 31063 5 1 1 31062
0 31064 7 1 2 57832 60078
0 31065 5 1 1 31064
0 31066 7 1 2 59333 31065
0 31067 5 1 1 31066
0 31068 7 1 2 63946 31067
0 31069 5 1 1 31068
0 31070 7 1 2 61102 75606
0 31071 5 1 1 31070
0 31072 7 1 2 74087 31071
0 31073 7 1 2 31069 31072
0 31074 7 1 2 31063 31073
0 31075 5 1 1 31074
0 31076 7 1 2 56936 31075
0 31077 5 1 1 31076
0 31078 7 1 2 61103 61989
0 31079 5 1 1 31078
0 31080 7 1 2 63038 74808
0 31081 7 1 2 74783 31080
0 31082 7 1 2 31079 31081
0 31083 5 1 1 31082
0 31084 7 1 2 56937 31083
0 31085 5 1 1 31084
0 31086 7 1 2 50812 31085
0 31087 5 1 1 31086
0 31088 7 1 2 48413 74799
0 31089 7 1 2 31087 31088
0 31090 5 1 1 31089
0 31091 7 1 2 31077 31090
0 31092 7 1 2 31055 31091
0 31093 7 1 2 31031 31092
0 31094 5 1 1 31093
0 31095 7 1 2 56560 31094
0 31096 5 1 1 31095
0 31097 7 2 2 61151 75595
0 31098 5 1 1 77821
0 31099 7 1 2 61927 62699
0 31100 5 1 1 31099
0 31101 7 1 2 47961 31100
0 31102 5 1 1 31101
0 31103 7 1 2 77820 31102
0 31104 5 1 1 31103
0 31105 7 1 2 55793 31104
0 31106 5 1 1 31105
0 31107 7 1 2 63930 60549
0 31108 7 1 2 72681 31107
0 31109 5 1 1 31108
0 31110 7 1 2 56379 31109
0 31111 5 1 1 31110
0 31112 7 1 2 61912 58618
0 31113 5 1 1 31112
0 31114 7 1 2 57033 31113
0 31115 7 1 2 61155 31114
0 31116 7 1 2 31111 31115
0 31117 7 1 2 31106 31116
0 31118 7 1 2 77822 31117
0 31119 5 1 1 31118
0 31120 7 1 2 57946 31119
0 31121 5 1 1 31120
0 31122 7 1 2 65816 74015
0 31123 5 1 1 31122
0 31124 7 1 2 61082 67446
0 31125 5 1 1 31124
0 31126 7 1 2 59195 31125
0 31127 7 1 2 31123 31126
0 31128 5 1 1 31127
0 31129 7 1 2 57947 31128
0 31130 5 1 1 31129
0 31131 7 2 2 58150 62214
0 31132 7 1 2 62781 69676
0 31133 7 1 2 77823 31132
0 31134 5 1 1 31133
0 31135 7 1 2 31130 31134
0 31136 5 1 1 31135
0 31137 7 1 2 48219 31136
0 31138 5 1 1 31137
0 31139 7 2 2 64333 61913
0 31140 7 1 2 62074 77825
0 31141 7 1 2 72642 31140
0 31142 5 1 1 31141
0 31143 7 1 2 31138 31142
0 31144 7 1 2 31121 31143
0 31145 7 1 2 31096 31144
0 31146 5 1 1 31145
0 31147 7 1 2 66608 31146
0 31148 5 1 1 31147
0 31149 7 1 2 30961 31148
0 31150 5 1 1 31149
0 31151 7 1 2 49769 31150
0 31152 5 1 1 31151
0 31153 7 1 2 61822 65817
0 31154 5 1 1 31153
0 31155 7 1 2 57177 61140
0 31156 5 1 1 31155
0 31157 7 1 2 77674 31156
0 31158 7 1 2 31154 31157
0 31159 5 1 1 31158
0 31160 7 1 2 54710 31159
0 31161 5 1 1 31160
0 31162 7 1 2 77764 31161
0 31163 5 1 1 31162
0 31164 7 1 2 57948 31163
0 31165 5 1 1 31164
0 31166 7 1 2 64853 66650
0 31167 5 1 1 31166
0 31168 7 1 2 64895 31167
0 31169 5 1 1 31168
0 31170 7 1 2 1619 31169
0 31171 5 1 1 31170
0 31172 7 1 2 54711 31171
0 31173 5 1 1 31172
0 31174 7 1 2 48414 77186
0 31175 5 1 1 31174
0 31176 7 1 2 64187 31175
0 31177 5 1 1 31176
0 31178 7 1 2 66975 31177
0 31179 5 1 1 31178
0 31180 7 1 2 31173 31179
0 31181 5 1 1 31180
0 31182 7 1 2 56561 31181
0 31183 5 1 1 31182
0 31184 7 1 2 31165 31183
0 31185 5 1 1 31184
0 31186 7 1 2 55794 31185
0 31187 5 1 1 31186
0 31188 7 1 2 49229 63147
0 31189 5 1 1 31188
0 31190 7 1 2 49230 74769
0 31191 5 1 1 31190
0 31192 7 1 2 65095 58619
0 31193 5 1 1 31192
0 31194 7 1 2 52319 31193
0 31195 7 1 2 31191 31194
0 31196 5 1 1 31195
0 31197 7 1 2 54369 61621
0 31198 7 1 2 31196 31197
0 31199 5 1 1 31198
0 31200 7 1 2 31189 31199
0 31201 5 1 1 31200
0 31202 7 1 2 54712 31201
0 31203 5 1 1 31202
0 31204 7 1 2 58620 67592
0 31205 5 1 1 31204
0 31206 7 1 2 49361 58333
0 31207 5 1 1 31206
0 31208 7 1 2 31205 31207
0 31209 5 1 1 31208
0 31210 7 1 2 60306 31209
0 31211 5 1 1 31210
0 31212 7 1 2 58183 57757
0 31213 5 2 1 31212
0 31214 7 1 2 62328 77827
0 31215 5 1 1 31214
0 31216 7 1 2 47962 58334
0 31217 5 1 1 31216
0 31218 7 1 2 31215 31217
0 31219 5 1 1 31218
0 31220 7 1 2 58311 31219
0 31221 5 1 1 31220
0 31222 7 1 2 31211 31221
0 31223 7 1 2 31203 31222
0 31224 5 1 1 31223
0 31225 7 1 2 56938 31224
0 31226 5 1 1 31225
0 31227 7 2 2 65096 59479
0 31228 5 1 1 77829
0 31229 7 1 2 57512 59417
0 31230 7 1 2 77830 31229
0 31231 5 1 1 31230
0 31232 7 1 2 31226 31231
0 31233 5 1 1 31232
0 31234 7 1 2 56562 31233
0 31235 5 1 1 31234
0 31236 7 1 2 65399 1813
0 31237 5 1 1 31236
0 31238 7 1 2 54370 31237
0 31239 5 1 1 31238
0 31240 7 1 2 59589 65951
0 31241 5 1 1 31240
0 31242 7 1 2 77766 31241
0 31243 7 1 2 31239 31242
0 31244 5 1 1 31243
0 31245 7 1 2 58621 31244
0 31246 5 1 1 31245
0 31247 7 1 2 58720 58647
0 31248 5 2 1 31247
0 31249 7 1 2 59998 77831
0 31250 5 1 1 31249
0 31251 7 1 2 57745 67467
0 31252 5 1 1 31251
0 31253 7 1 2 68018 77768
0 31254 7 1 2 31252 31253
0 31255 7 1 2 31250 31254
0 31256 5 1 1 31255
0 31257 7 1 2 58312 31256
0 31258 5 1 1 31257
0 31259 7 1 2 54713 70916
0 31260 5 1 1 31259
0 31261 7 1 2 56226 31260
0 31262 5 1 1 31261
0 31263 7 1 2 74145 31262
0 31264 5 1 1 31263
0 31265 7 2 2 54714 74748
0 31266 5 1 1 77833
0 31267 7 1 2 59225 77834
0 31268 5 1 1 31267
0 31269 7 1 2 58924 31268
0 31270 7 1 2 31264 31269
0 31271 7 1 2 31258 31270
0 31272 7 1 2 31246 31271
0 31273 5 1 1 31272
0 31274 7 1 2 57949 31273
0 31275 5 1 1 31274
0 31276 7 1 2 57950 65420
0 31277 5 1 1 31276
0 31278 7 1 2 48545 67307
0 31279 7 1 2 65839 31278
0 31280 5 1 1 31279
0 31281 7 1 2 31277 31280
0 31282 5 1 1 31281
0 31283 7 1 2 48415 31282
0 31284 5 1 1 31283
0 31285 7 1 2 57951 74375
0 31286 5 1 1 31285
0 31287 7 1 2 31284 31286
0 31288 5 1 1 31287
0 31289 7 1 2 58162 31288
0 31290 5 1 1 31289
0 31291 7 1 2 48649 58500
0 31292 5 1 1 31291
0 31293 7 1 2 63374 31292
0 31294 5 1 1 31293
0 31295 7 1 2 48546 74376
0 31296 5 1 1 31295
0 31297 7 1 2 59569 61930
0 31298 5 1 1 31297
0 31299 7 1 2 3150 4652
0 31300 7 1 2 31298 31299
0 31301 5 1 1 31300
0 31302 7 1 2 48416 31301
0 31303 5 1 1 31302
0 31304 7 1 2 31296 31303
0 31305 5 1 1 31304
0 31306 7 1 2 31294 31305
0 31307 5 1 1 31306
0 31308 7 1 2 31290 31307
0 31309 7 1 2 31275 31308
0 31310 7 1 2 31235 31309
0 31311 7 1 2 31187 31310
0 31312 5 1 1 31311
0 31313 7 1 2 69804 31312
0 31314 5 1 1 31313
0 31315 7 1 2 63381 68710
0 31316 7 1 2 63372 31315
0 31317 5 2 1 31316
0 31318 7 1 2 64268 64172
0 31319 7 1 2 68702 31318
0 31320 7 1 2 60838 31319
0 31321 7 1 2 72432 31320
0 31322 5 1 1 31321
0 31323 7 1 2 77835 31322
0 31324 7 1 2 31314 31323
0 31325 5 1 1 31324
0 31326 7 1 2 51082 31325
0 31327 5 1 1 31326
0 31328 7 1 2 31152 31327
0 31329 5 1 1 31328
0 31330 7 1 2 48772 31329
0 31331 5 1 1 31330
0 31332 7 2 2 48417 57775
0 31333 5 1 1 77837
0 31334 7 1 2 63276 77838
0 31335 5 1 1 31334
0 31336 7 1 2 11411 31335
0 31337 5 1 1 31336
0 31338 7 1 2 56563 31337
0 31339 5 1 1 31338
0 31340 7 1 2 54076 64741
0 31341 5 1 1 31340
0 31342 7 1 2 31339 31341
0 31343 5 1 1 31342
0 31344 7 1 2 54715 31343
0 31345 5 1 1 31344
0 31346 7 1 2 61162 31333
0 31347 5 1 1 31346
0 31348 7 1 2 48650 31347
0 31349 5 1 1 31348
0 31350 7 1 2 65547 62215
0 31351 5 1 1 31350
0 31352 7 1 2 31349 31351
0 31353 5 1 1 31352
0 31354 7 1 2 49600 31353
0 31355 5 1 1 31354
0 31356 7 1 2 31345 31355
0 31357 5 1 1 31356
0 31358 7 1 2 52661 31357
0 31359 5 1 1 31358
0 31360 7 1 2 59378 76619
0 31361 7 1 2 64309 31360
0 31362 5 1 1 31361
0 31363 7 1 2 31359 31362
0 31364 5 1 1 31363
0 31365 7 1 2 62065 31364
0 31366 5 1 1 31365
0 31367 7 1 2 49486 73432
0 31368 5 1 1 31367
0 31369 7 1 2 23088 31368
0 31370 5 1 1 31369
0 31371 7 1 2 48547 31370
0 31372 5 1 1 31371
0 31373 7 1 2 52662 76512
0 31374 5 1 1 31373
0 31375 7 1 2 31372 31374
0 31376 5 1 1 31375
0 31377 7 1 2 74752 31376
0 31378 5 1 1 31377
0 31379 7 1 2 53235 61928
0 31380 5 2 1 31379
0 31381 7 1 2 49601 77839
0 31382 5 1 1 31381
0 31383 7 1 2 62138 66236
0 31384 5 2 1 31383
0 31385 7 1 2 31382 77841
0 31386 5 2 1 31385
0 31387 7 1 2 52663 77843
0 31388 5 1 1 31387
0 31389 7 1 2 31378 31388
0 31390 5 1 1 31389
0 31391 7 1 2 48651 31390
0 31392 5 1 1 31391
0 31393 7 2 2 65024 77227
0 31394 5 1 1 77845
0 31395 7 1 2 74753 77846
0 31396 5 1 1 31395
0 31397 7 1 2 77842 31396
0 31398 5 1 1 31397
0 31399 7 1 2 75503 31398
0 31400 5 1 1 31399
0 31401 7 1 2 31392 31400
0 31402 5 1 1 31401
0 31403 7 1 2 71430 31402
0 31404 5 1 1 31403
0 31405 7 4 2 52664 58691
0 31406 5 2 1 77847
0 31407 7 2 2 56641 60601
0 31408 5 2 1 77853
0 31409 7 1 2 57952 77855
0 31410 5 1 1 31409
0 31411 7 1 2 61160 74754
0 31412 5 1 1 31411
0 31413 7 1 2 56939 77856
0 31414 5 1 1 31413
0 31415 7 1 2 31412 31414
0 31416 5 1 1 31415
0 31417 7 1 2 56564 31416
0 31418 5 1 1 31417
0 31419 7 1 2 31410 31418
0 31420 5 1 1 31419
0 31421 7 1 2 77848 31420
0 31422 5 1 1 31421
0 31423 7 1 2 31404 31422
0 31424 7 1 2 31366 31423
0 31425 5 1 1 31424
0 31426 7 1 2 49362 31425
0 31427 5 1 1 31426
0 31428 7 1 2 47963 77145
0 31429 5 2 1 31428
0 31430 7 1 2 48220 61784
0 31431 5 1 1 31430
0 31432 7 2 2 62659 31431
0 31433 5 2 1 77859
0 31434 7 1 2 77857 77860
0 31435 5 1 1 31434
0 31436 7 1 2 54716 31435
0 31437 5 1 1 31436
0 31438 7 1 2 53236 66228
0 31439 5 1 1 31438
0 31440 7 1 2 48418 31439
0 31441 5 1 1 31440
0 31442 7 2 2 50813 61959
0 31443 5 1 1 77863
0 31444 7 1 2 49487 31443
0 31445 5 1 1 31444
0 31446 7 1 2 62199 67080
0 31447 5 1 1 31446
0 31448 7 1 2 58622 31447
0 31449 5 1 1 31448
0 31450 7 1 2 31445 31449
0 31451 7 1 2 31441 31450
0 31452 7 1 2 31437 31451
0 31453 5 1 1 31452
0 31454 7 1 2 75547 31453
0 31455 5 1 1 31454
0 31456 7 1 2 61780 59389
0 31457 5 1 1 31456
0 31458 7 1 2 67308 31457
0 31459 5 1 1 31458
0 31460 7 1 2 63055 74694
0 31461 5 1 1 31460
0 31462 7 1 2 31459 31461
0 31463 5 1 1 31462
0 31464 7 1 2 52665 31463
0 31465 5 1 1 31464
0 31466 7 1 2 53371 63379
0 31467 7 1 2 59393 31466
0 31468 7 1 2 66224 31467
0 31469 5 1 1 31468
0 31470 7 1 2 31465 31469
0 31471 5 1 1 31470
0 31472 7 1 2 48221 31471
0 31473 5 1 1 31472
0 31474 7 1 2 62660 77858
0 31475 5 1 1 31474
0 31476 7 3 2 56565 63580
0 31477 7 1 2 31475 77865
0 31478 5 1 1 31477
0 31479 7 1 2 31473 31478
0 31480 5 1 1 31479
0 31481 7 1 2 49488 31480
0 31482 5 1 1 31481
0 31483 7 1 2 54077 58623
0 31484 5 2 1 31483
0 31485 7 1 2 52320 77864
0 31486 7 1 2 77868 31485
0 31487 5 1 1 31486
0 31488 7 1 2 75548 31487
0 31489 5 1 1 31488
0 31490 7 1 2 31482 31489
0 31491 5 1 1 31490
0 31492 7 1 2 48548 31491
0 31493 5 1 1 31492
0 31494 7 1 2 31455 31493
0 31495 7 1 2 31427 31494
0 31496 5 1 1 31495
0 31497 7 1 2 59685 31496
0 31498 5 1 1 31497
0 31499 7 1 2 77861 75590
0 31500 5 1 1 31499
0 31501 7 1 2 62130 63581
0 31502 7 1 2 56785 31501
0 31503 5 1 1 31502
0 31504 7 1 2 31500 31503
0 31505 5 1 1 31504
0 31506 7 1 2 47964 31505
0 31507 5 1 1 31506
0 31508 7 2 2 56380 63954
0 31509 5 1 1 77870
0 31510 7 2 2 57034 31509
0 31511 5 1 1 77872
0 31512 7 1 2 58041 77873
0 31513 5 1 1 31512
0 31514 7 1 2 77866 31513
0 31515 5 1 1 31514
0 31516 7 1 2 31507 31515
0 31517 5 1 1 31516
0 31518 7 1 2 54371 31517
0 31519 5 1 1 31518
0 31520 7 1 2 48652 77844
0 31521 5 1 1 31520
0 31522 7 1 2 64238 66705
0 31523 5 1 1 31522
0 31524 7 1 2 31521 31523
0 31525 5 3 1 31524
0 31526 7 1 2 77874 75537
0 31527 5 1 1 31526
0 31528 7 1 2 31519 31527
0 31529 5 1 1 31528
0 31530 7 1 2 49363 31529
0 31531 5 1 1 31530
0 31532 7 1 2 62439 77867
0 31533 5 1 1 31532
0 31534 7 1 2 66571 75577
0 31535 5 1 1 31534
0 31536 7 1 2 31533 31535
0 31537 5 1 1 31536
0 31538 7 1 2 49489 31537
0 31539 5 1 1 31538
0 31540 7 2 2 52666 72371
0 31541 7 1 2 71845 77877
0 31542 5 1 1 31541
0 31543 7 1 2 31539 31542
0 31544 5 1 1 31543
0 31545 7 1 2 48549 31544
0 31546 5 1 1 31545
0 31547 7 1 2 53237 63957
0 31548 5 1 1 31547
0 31549 7 1 2 62732 31548
0 31550 5 1 1 31549
0 31551 7 1 2 74696 31550
0 31552 5 1 1 31551
0 31553 7 1 2 75549 31552
0 31554 5 1 1 31553
0 31555 7 1 2 31546 31554
0 31556 5 1 1 31555
0 31557 7 1 2 59686 31556
0 31558 5 1 1 31557
0 31559 7 1 2 58349 56751
0 31560 7 1 2 77875 31559
0 31561 5 1 1 31560
0 31562 7 2 2 56381 62440
0 31563 7 1 2 62733 77879
0 31564 5 1 1 31563
0 31565 7 1 2 59486 5265
0 31566 7 1 2 31564 31565
0 31567 5 1 1 31566
0 31568 7 1 2 49602 31567
0 31569 5 1 1 31568
0 31570 7 1 2 65074 63955
0 31571 5 1 1 31570
0 31572 7 1 2 31569 31571
0 31573 5 1 1 31572
0 31574 7 1 2 48653 31573
0 31575 5 1 1 31574
0 31576 7 1 2 58231 62139
0 31577 7 1 2 64181 31576
0 31578 5 1 1 31577
0 31579 7 1 2 31575 31578
0 31580 7 1 2 31561 31579
0 31581 5 1 1 31580
0 31582 7 1 2 52667 31581
0 31583 5 1 1 31582
0 31584 7 1 2 31558 31583
0 31585 7 1 2 31531 31584
0 31586 5 1 1 31585
0 31587 7 1 2 55795 31586
0 31588 5 1 1 31587
0 31589 7 1 2 57326 65793
0 31590 5 1 1 31589
0 31591 7 1 2 67240 31590
0 31592 5 1 1 31591
0 31593 7 1 2 47965 75565
0 31594 5 1 1 31593
0 31595 7 1 2 31592 31594
0 31596 5 1 1 31595
0 31597 7 1 2 52668 31596
0 31598 5 1 1 31597
0 31599 7 1 2 71969 75518
0 31600 7 1 2 64339 31599
0 31601 5 1 1 31600
0 31602 7 1 2 31598 31601
0 31603 5 1 1 31602
0 31604 7 1 2 54078 31603
0 31605 5 1 1 31604
0 31606 7 1 2 57352 77878
0 31607 5 1 1 31606
0 31608 7 1 2 31605 31607
0 31609 5 1 1 31608
0 31610 7 1 2 48419 61979
0 31611 5 1 1 31610
0 31612 7 1 2 59731 31611
0 31613 5 1 1 31612
0 31614 7 1 2 31609 31613
0 31615 5 1 1 31614
0 31616 7 1 2 56382 28947
0 31617 5 1 1 31616
0 31618 7 1 2 65149 70364
0 31619 5 1 1 31618
0 31620 7 1 2 4909 31619
0 31621 7 1 2 31617 31620
0 31622 5 1 1 31621
0 31623 7 1 2 57953 31622
0 31624 5 1 1 31623
0 31625 7 1 2 59047 61392
0 31626 7 1 2 74584 31625
0 31627 5 1 1 31626
0 31628 7 1 2 31624 31627
0 31629 5 1 1 31628
0 31630 7 1 2 54717 31629
0 31631 5 1 1 31630
0 31632 7 1 2 59517 62217
0 31633 5 1 1 31632
0 31634 7 1 2 48222 31633
0 31635 5 1 1 31634
0 31636 7 1 2 59412 31635
0 31637 5 1 1 31636
0 31638 7 1 2 31637 77876
0 31639 5 1 1 31638
0 31640 7 1 2 64297 31639
0 31641 7 1 2 31631 31640
0 31642 5 1 1 31641
0 31643 7 1 2 52669 31642
0 31644 5 1 1 31643
0 31645 7 1 2 31615 31644
0 31646 7 1 2 31588 31645
0 31647 7 1 2 31498 31646
0 31648 5 1 1 31647
0 31649 7 1 2 55371 31648
0 31650 5 1 1 31649
0 31651 7 1 2 64269 64303
0 31652 7 1 2 64256 59837
0 31653 7 1 2 68711 31652
0 31654 7 1 2 31651 31653
0 31655 5 1 1 31654
0 31656 7 1 2 77836 31655
0 31657 7 1 2 31650 31656
0 31658 5 1 1 31657
0 31659 7 1 2 62683 31658
0 31660 5 1 1 31659
0 31661 7 2 2 60576 77799
0 31662 7 1 2 48654 77881
0 31663 5 1 1 31662
0 31664 7 4 2 49490 58692
0 31665 5 1 1 77883
0 31666 7 3 2 52173 58540
0 31667 7 1 2 77884 77887
0 31668 5 1 1 31667
0 31669 7 1 2 31663 31668
0 31670 5 1 1 31669
0 31671 7 1 2 77733 31670
0 31672 5 1 1 31671
0 31673 7 1 2 52442 77882
0 31674 5 1 1 31673
0 31675 7 1 2 76944 31674
0 31676 5 1 1 31675
0 31677 7 1 2 55925 31676
0 31678 5 1 1 31677
0 31679 7 1 2 54372 72989
0 31680 5 1 1 31679
0 31681 7 1 2 31678 31680
0 31682 5 1 1 31681
0 31683 7 1 2 58042 31682
0 31684 5 1 1 31683
0 31685 7 1 2 66651 76735
0 31686 5 1 1 31685
0 31687 7 1 2 59381 31686
0 31688 5 1 1 31687
0 31689 7 1 2 56464 31688
0 31690 5 1 1 31689
0 31691 7 1 2 31684 31690
0 31692 5 1 1 31691
0 31693 7 1 2 62922 31692
0 31694 5 1 1 31693
0 31695 7 1 2 31672 31694
0 31696 5 1 1 31695
0 31697 7 1 2 55051 31696
0 31698 5 1 1 31697
0 31699 7 1 2 76744 28831
0 31700 5 1 1 31699
0 31701 7 1 2 49603 31700
0 31702 5 1 1 31701
0 31703 7 1 2 71257 77885
0 31704 5 1 1 31703
0 31705 7 1 2 31702 31704
0 31706 5 1 1 31705
0 31707 7 1 2 62923 59918
0 31708 7 1 2 31706 31707
0 31709 5 1 1 31708
0 31710 7 1 2 31698 31709
0 31711 5 1 1 31710
0 31712 7 1 2 70728 31711
0 31713 5 1 1 31712
0 31714 7 2 2 61649 62877
0 31715 7 1 2 77754 77890
0 31716 5 1 1 31715
0 31717 7 2 2 62924 65772
0 31718 7 1 2 77758 77892
0 31719 5 1 1 31718
0 31720 7 1 2 31716 31719
0 31721 5 1 1 31720
0 31722 7 1 2 55052 31721
0 31723 5 1 1 31722
0 31724 7 1 2 67218 71250
0 31725 5 1 1 31724
0 31726 7 2 2 49604 31725
0 31727 5 1 1 77894
0 31728 7 1 2 77802 31727
0 31729 5 1 1 31728
0 31730 7 1 2 77893 31729
0 31731 5 1 1 31730
0 31732 7 1 2 31723 31731
0 31733 5 1 1 31732
0 31734 7 1 2 52174 31733
0 31735 5 1 1 31734
0 31736 7 1 2 52555 73067
0 31737 5 1 1 31736
0 31738 7 1 2 53238 73078
0 31739 5 1 1 31738
0 31740 7 1 2 31737 31739
0 31741 5 1 1 31740
0 31742 7 1 2 49605 31741
0 31743 5 1 1 31742
0 31744 7 1 2 73070 76620
0 31745 5 1 1 31744
0 31746 7 1 2 31743 31745
0 31747 5 1 1 31746
0 31748 7 1 2 58541 31747
0 31749 5 1 1 31748
0 31750 7 1 2 53239 73068
0 31751 5 1 1 31750
0 31752 7 1 2 73085 31751
0 31753 5 1 1 31752
0 31754 7 1 2 49606 75819
0 31755 5 1 1 31754
0 31756 7 1 2 56566 31755
0 31757 7 1 2 31753 31756
0 31758 5 1 1 31757
0 31759 7 1 2 31749 31758
0 31760 5 1 1 31759
0 31761 7 1 2 62925 31760
0 31762 5 1 1 31761
0 31763 7 1 2 31735 31762
0 31764 5 1 1 31763
0 31765 7 1 2 51969 31764
0 31766 5 1 1 31765
0 31767 7 1 2 58542 77746
0 31768 5 1 1 31767
0 31769 7 1 2 48773 72334
0 31770 7 1 2 75794 31769
0 31771 5 1 1 31770
0 31772 7 1 2 53240 62571
0 31773 7 1 2 58115 31772
0 31774 7 1 2 31771 31773
0 31775 5 1 1 31774
0 31776 7 1 2 31768 31775
0 31777 5 1 1 31776
0 31778 7 1 2 63459 31777
0 31779 5 1 1 31778
0 31780 7 2 2 59146 66652
0 31781 7 1 2 52175 49607
0 31782 7 1 2 62926 31781
0 31783 7 1 2 77896 31782
0 31784 5 1 1 31783
0 31785 7 1 2 31779 31784
0 31786 5 1 1 31785
0 31787 7 1 2 70252 31786
0 31788 5 1 1 31787
0 31789 7 1 2 52176 75823
0 31790 5 1 1 31789
0 31791 7 1 2 58522 62375
0 31792 5 1 1 31791
0 31793 7 1 2 77800 31792
0 31794 5 1 1 31793
0 31795 7 1 2 31790 31794
0 31796 5 1 1 31795
0 31797 7 1 2 62927 73392
0 31798 7 1 2 31796 31797
0 31799 5 1 1 31798
0 31800 7 1 2 77239 30125
0 31801 5 1 1 31800
0 31802 7 1 2 58543 63460
0 31803 7 1 2 75294 31802
0 31804 7 1 2 31801 31803
0 31805 5 1 1 31804
0 31806 7 1 2 31799 31805
0 31807 5 1 1 31806
0 31808 7 1 2 49608 31807
0 31809 5 1 1 31808
0 31810 7 1 2 62641 71176
0 31811 7 1 2 74635 75489
0 31812 7 1 2 75915 31811
0 31813 7 1 2 31810 31812
0 31814 5 1 1 31813
0 31815 7 1 2 31809 31814
0 31816 7 1 2 31788 31815
0 31817 7 1 2 31766 31816
0 31818 7 1 2 31713 31817
0 31819 5 1 1 31818
0 31820 7 1 2 55372 31819
0 31821 5 1 1 31820
0 31822 7 2 2 48774 64279
0 31823 7 1 2 63738 66379
0 31824 7 2 2 77898 31823
0 31825 7 1 2 73195 77900
0 31826 5 1 1 31825
0 31827 7 1 2 51970 77901
0 31828 5 1 1 31827
0 31829 7 1 2 57327 70253
0 31830 5 1 1 31829
0 31831 7 1 2 57035 73023
0 31832 5 1 1 31831
0 31833 7 1 2 71563 31832
0 31834 5 1 1 31833
0 31835 7 1 2 52177 31834
0 31836 5 1 1 31835
0 31837 7 1 2 73033 31836
0 31838 5 1 1 31837
0 31839 7 1 2 51971 31838
0 31840 5 1 1 31839
0 31841 7 1 2 31830 31840
0 31842 5 1 1 31841
0 31843 7 1 2 49609 31842
0 31844 5 1 1 31843
0 31845 7 2 2 54718 76621
0 31846 7 1 2 76830 77902
0 31847 5 1 1 31846
0 31848 7 1 2 31844 31847
0 31849 5 1 1 31848
0 31850 7 1 2 62928 31849
0 31851 5 1 1 31850
0 31852 7 1 2 51083 31851
0 31853 5 1 1 31852
0 31854 7 2 2 51972 77128
0 31855 5 1 1 77904
0 31856 7 1 2 65362 31855
0 31857 5 1 1 31856
0 31858 7 1 2 48655 31857
0 31859 5 1 1 31858
0 31860 7 1 2 64334 72975
0 31861 5 1 1 31860
0 31862 7 1 2 31859 31861
0 31863 5 1 1 31862
0 31864 7 1 2 77734 31863
0 31865 5 1 1 31864
0 31866 7 1 2 70134 73572
0 31867 5 1 1 31866
0 31868 7 1 2 28786 31867
0 31869 5 1 1 31868
0 31870 7 1 2 62929 31869
0 31871 5 1 1 31870
0 31872 7 1 2 31865 31871
0 31873 5 1 1 31872
0 31874 7 1 2 54719 31873
0 31875 5 1 1 31874
0 31876 7 1 2 74869 25952
0 31877 5 1 1 31876
0 31878 7 1 2 49770 76740
0 31879 7 1 2 76254 31878
0 31880 7 1 2 31877 31879
0 31881 5 1 1 31880
0 31882 7 1 2 55053 31881
0 31883 7 1 2 31875 31882
0 31884 5 1 1 31883
0 31885 7 1 2 55373 31884
0 31886 7 1 2 31853 31885
0 31887 5 1 1 31886
0 31888 7 1 2 31828 31887
0 31889 5 1 1 31888
0 31890 7 1 2 57636 31889
0 31891 5 1 1 31890
0 31892 7 1 2 31826 31891
0 31893 7 1 2 31821 31892
0 31894 5 1 1 31893
0 31895 7 1 2 58444 31894
0 31896 5 1 1 31895
0 31897 7 1 2 51597 31896
0 31898 7 1 2 31660 31897
0 31899 7 1 2 31331 31898
0 31900 7 1 2 30674 31899
0 31901 5 1 1 31900
0 31902 7 1 2 53695 31901
0 31903 7 1 2 29633 31902
0 31904 5 1 1 31903
0 31905 7 1 2 52811 31904
0 31906 7 1 2 25598 31905
0 31907 5 1 1 31906
0 31908 7 2 2 57365 75014
0 31909 7 2 2 60123 70448
0 31910 5 2 1 77908
0 31911 7 1 2 56135 77910
0 31912 5 1 1 31911
0 31913 7 1 2 75060 31912
0 31914 7 1 2 77906 31913
0 31915 5 1 1 31914
0 31916 7 2 2 58901 76968
0 31917 5 1 1 77912
0 31918 7 1 2 70135 77913
0 31919 5 1 1 31918
0 31920 7 1 2 70181 31919
0 31921 5 1 1 31920
0 31922 7 1 2 52998 58693
0 31923 7 1 2 31921 31922
0 31924 5 1 1 31923
0 31925 7 1 2 31915 31924
0 31926 5 1 1 31925
0 31927 7 1 2 68587 31926
0 31928 5 1 1 31927
0 31929 7 2 2 52999 54373
0 31930 7 3 2 68703 77914
0 31931 5 1 1 77916
0 31932 7 1 2 52443 75804
0 31933 7 1 2 75965 31932
0 31934 5 1 1 31933
0 31935 7 1 2 31931 31934
0 31936 5 1 1 31935
0 31937 7 1 2 55926 31936
0 31938 5 1 1 31937
0 31939 7 1 2 53372 2109
0 31940 5 1 1 31939
0 31941 7 1 2 50814 64727
0 31942 7 1 2 31940 31941
0 31943 5 1 1 31942
0 31944 7 1 2 31938 31943
0 31945 5 1 1 31944
0 31946 7 1 2 48775 31945
0 31947 5 1 1 31946
0 31948 7 1 2 63786 76227
0 31949 7 1 2 75851 31948
0 31950 5 1 1 31949
0 31951 7 1 2 31947 31950
0 31952 5 1 1 31951
0 31953 7 1 2 62108 31952
0 31954 5 1 1 31953
0 31955 7 2 2 58694 75519
0 31956 5 1 1 77919
0 31957 7 1 2 51364 77920
0 31958 7 1 2 58583 31957
0 31959 7 1 2 76140 31958
0 31960 5 1 1 31959
0 31961 7 1 2 31954 31960
0 31962 5 1 1 31961
0 31963 7 1 2 50258 31962
0 31964 5 1 1 31963
0 31965 7 1 2 59315 69883
0 31966 5 1 1 31965
0 31967 7 1 2 310 31966
0 31968 5 1 1 31967
0 31969 7 1 2 66706 31968
0 31970 5 1 1 31969
0 31971 7 1 2 57798 74030
0 31972 5 2 1 31971
0 31973 7 1 2 57036 77921
0 31974 5 1 1 31973
0 31975 7 1 2 54374 76724
0 31976 7 1 2 31974 31975
0 31977 5 1 1 31976
0 31978 7 1 2 31970 31977
0 31979 5 1 1 31978
0 31980 7 1 2 75520 31979
0 31981 5 1 1 31980
0 31982 7 1 2 53373 75612
0 31983 5 1 1 31982
0 31984 7 1 2 48776 10474
0 31985 7 1 2 31983 31984
0 31986 5 1 1 31985
0 31987 7 1 2 50815 31986
0 31988 7 1 2 31981 31987
0 31989 5 1 1 31988
0 31990 7 1 2 53000 57356
0 31991 5 1 1 31990
0 31992 7 1 2 64674 10246
0 31993 7 1 2 31991 31992
0 31994 5 1 1 31993
0 31995 7 1 2 64615 31994
0 31996 5 1 1 31995
0 31997 7 1 2 54720 31996
0 31998 5 1 1 31997
0 31999 7 1 2 51365 31998
0 32000 7 1 2 31989 31999
0 32001 5 1 1 32000
0 32002 7 1 2 31964 32001
0 32003 5 1 1 32002
0 32004 7 1 2 53540 32003
0 32005 5 1 1 32004
0 32006 7 1 2 31928 32005
0 32007 5 1 1 32006
0 32008 7 1 2 51084 32007
0 32009 5 1 1 32008
0 32010 7 2 2 64019 70136
0 32011 5 1 1 77923
0 32012 7 1 2 63209 63739
0 32013 7 1 2 77924 32012
0 32014 5 1 1 32013
0 32015 7 1 2 32009 32014
0 32016 5 1 1 32015
0 32017 7 1 2 53696 32016
0 32018 5 1 1 32017
0 32019 7 1 2 48656 29417
0 32020 5 1 1 32019
0 32021 7 2 2 76580 32020
0 32022 7 1 2 73253 77925
0 32023 5 1 1 32022
0 32024 7 1 2 76221 32023
0 32025 5 1 1 32024
0 32026 7 3 2 53697 60684
0 32027 7 2 2 55374 58839
0 32028 7 1 2 73313 77930
0 32029 7 1 2 77927 32028
0 32030 5 1 1 32029
0 32031 7 1 2 67894 32030
0 32032 5 1 1 32031
0 32033 7 1 2 32025 32032
0 32034 5 1 1 32033
0 32035 7 1 2 54079 64103
0 32036 5 1 1 32035
0 32037 7 1 2 49610 58589
0 32038 5 1 1 32037
0 32039 7 1 2 32036 32038
0 32040 5 1 1 32039
0 32041 7 1 2 69884 32040
0 32042 5 1 1 32041
0 32043 7 1 2 56752 63877
0 32044 5 1 1 32043
0 32045 7 1 2 2454 32044
0 32046 5 1 1 32045
0 32047 7 1 2 58584 32046
0 32048 5 1 1 32047
0 32049 7 1 2 53541 68026
0 32050 7 1 2 32048 32049
0 32051 7 1 2 32042 32050
0 32052 5 1 1 32051
0 32053 7 1 2 61211 76128
0 32054 5 1 1 32053
0 32055 7 1 2 54721 32054
0 32056 7 1 2 32052 32055
0 32057 5 1 1 32056
0 32058 7 1 2 77696 77922
0 32059 5 1 1 32058
0 32060 7 1 2 72318 32059
0 32061 5 1 1 32060
0 32062 7 1 2 59226 75496
0 32063 5 1 1 32062
0 32064 7 1 2 58808 67241
0 32065 5 1 1 32064
0 32066 7 3 2 64577 32065
0 32067 7 1 2 25668 77932
0 32068 5 1 1 32067
0 32069 7 1 2 32063 32068
0 32070 7 1 2 32061 32069
0 32071 7 1 2 32057 32070
0 32072 5 1 1 32071
0 32073 7 1 2 54375 32072
0 32074 5 1 1 32073
0 32075 7 2 2 72319 75676
0 32076 7 1 2 62761 77935
0 32077 5 1 1 32076
0 32078 7 1 2 56753 77933
0 32079 5 1 1 32078
0 32080 7 1 2 63985 72320
0 32081 7 1 2 58642 32080
0 32082 5 1 1 32081
0 32083 7 1 2 32079 32082
0 32084 5 1 1 32083
0 32085 7 1 2 77102 32084
0 32086 5 1 1 32085
0 32087 7 1 2 32077 32086
0 32088 5 1 1 32087
0 32089 7 1 2 55796 32088
0 32090 5 1 1 32089
0 32091 7 1 2 57328 75575
0 32092 5 1 1 32091
0 32093 7 1 2 49364 77871
0 32094 5 3 1 32093
0 32095 7 1 2 67201 77937
0 32096 5 1 1 32095
0 32097 7 1 2 63632 32096
0 32098 7 1 2 32092 32097
0 32099 5 1 1 32098
0 32100 7 1 2 53542 32099
0 32101 5 1 1 32100
0 32102 7 1 2 49771 65237
0 32103 5 1 1 32102
0 32104 7 1 2 49611 32103
0 32105 7 1 2 32101 32104
0 32106 5 1 1 32105
0 32107 7 1 2 59999 77936
0 32108 5 1 1 32107
0 32109 7 1 2 75593 77934
0 32110 5 1 1 32109
0 32111 7 1 2 32108 32110
0 32112 5 1 1 32111
0 32113 7 1 2 58624 32112
0 32114 5 1 1 32113
0 32115 7 1 2 54080 67219
0 32116 5 1 1 32115
0 32117 7 1 2 31228 32116
0 32118 5 1 1 32117
0 32119 7 1 2 72321 32118
0 32120 7 1 2 66187 32119
0 32121 5 1 1 32120
0 32122 7 1 2 66256 75490
0 32123 7 1 2 67415 32122
0 32124 5 1 1 32123
0 32125 7 1 2 32121 32124
0 32126 7 1 2 32114 32125
0 32127 7 1 2 32106 32126
0 32128 7 1 2 32090 32127
0 32129 7 1 2 32074 32128
0 32130 5 1 1 32129
0 32131 7 1 2 51366 32130
0 32132 5 1 1 32131
0 32133 7 1 2 75751 76589
0 32134 5 1 1 32133
0 32135 7 3 2 52444 53543
0 32136 7 1 2 64820 77940
0 32137 5 1 1 32136
0 32138 7 1 2 54722 72464
0 32139 5 1 1 32138
0 32140 7 1 2 32137 32139
0 32141 5 1 1 32140
0 32142 7 1 2 55927 32141
0 32143 5 1 1 32142
0 32144 7 1 2 25190 32143
0 32145 5 1 1 32144
0 32146 7 1 2 53001 32145
0 32147 5 1 1 32146
0 32148 7 1 2 3991 75359
0 32149 7 1 2 74415 32148
0 32150 5 1 1 32149
0 32151 7 1 2 32147 32150
0 32152 5 1 1 32151
0 32153 7 1 2 62109 32152
0 32154 5 1 1 32153
0 32155 7 1 2 69805 75779
0 32156 5 1 1 32155
0 32157 7 1 2 32154 32156
0 32158 5 1 1 32157
0 32159 7 1 2 50259 32158
0 32160 5 1 1 32159
0 32161 7 1 2 77528 76590
0 32162 5 1 1 32161
0 32163 7 1 2 75786 77917
0 32164 5 1 1 32163
0 32165 7 1 2 32162 32164
0 32166 5 1 1 32165
0 32167 7 1 2 53241 32166
0 32168 5 1 1 32167
0 32169 7 1 2 65495 66382
0 32170 7 1 2 74416 75765
0 32171 7 1 2 32169 32170
0 32172 5 1 1 32171
0 32173 7 1 2 32168 32172
0 32174 7 1 2 32160 32173
0 32175 7 1 2 32134 32174
0 32176 7 1 2 32132 32175
0 32177 5 1 1 32176
0 32178 7 1 2 53698 32177
0 32179 5 1 1 32178
0 32180 7 1 2 32034 32179
0 32181 5 1 1 32180
0 32182 7 1 2 51085 32181
0 32183 5 1 1 32182
0 32184 7 1 2 73139 68310
0 32185 5 1 1 32184
0 32186 7 1 2 53374 75651
0 32187 5 1 1 32186
0 32188 7 1 2 63947 76228
0 32189 5 1 1 32188
0 32190 7 1 2 32187 32189
0 32191 5 1 1 32190
0 32192 7 1 2 57833 32191
0 32193 5 1 1 32192
0 32194 7 2 2 64282 57805
0 32195 7 1 2 69396 77943
0 32196 5 1 1 32195
0 32197 7 1 2 2568 57375
0 32198 5 1 1 32197
0 32199 7 1 2 32196 32198
0 32200 7 1 2 32193 32199
0 32201 5 1 1 32200
0 32202 7 1 2 54723 32201
0 32203 5 1 1 32202
0 32204 7 2 2 54724 63887
0 32205 5 1 1 77945
0 32206 7 1 2 77944 77946
0 32207 5 1 1 32206
0 32208 7 1 2 57102 65889
0 32209 5 1 1 32208
0 32210 7 1 2 57366 32209
0 32211 5 1 1 32210
0 32212 7 1 2 66257 32211
0 32213 5 1 1 32212
0 32214 7 1 2 32207 32213
0 32215 5 1 1 32214
0 32216 7 1 2 56754 32215
0 32217 5 1 1 32216
0 32218 7 1 2 50816 57103
0 32219 7 1 2 74135 32218
0 32220 5 1 1 32219
0 32221 7 1 2 62782 76229
0 32222 5 1 1 32221
0 32223 7 1 2 32220 32222
0 32224 7 1 2 75707 32223
0 32225 7 1 2 32217 32224
0 32226 5 1 1 32225
0 32227 7 1 2 55797 32226
0 32228 5 1 1 32227
0 32229 7 1 2 62410 56940
0 32230 5 1 1 32229
0 32231 7 1 2 77938 32230
0 32232 5 1 1 32231
0 32233 7 1 2 53375 32232
0 32234 5 1 1 32233
0 32235 7 1 2 54725 77642
0 32236 7 1 2 32234 32235
0 32237 5 1 1 32236
0 32238 7 1 2 50817 64100
0 32239 5 1 1 32238
0 32240 7 1 2 60247 32239
0 32241 7 1 2 32237 32240
0 32242 5 1 1 32241
0 32243 7 1 2 53544 30572
0 32244 7 1 2 32242 32243
0 32245 7 1 2 75664 32244
0 32246 7 1 2 32228 32245
0 32247 7 1 2 32203 32246
0 32248 5 1 1 32247
0 32249 7 1 2 49772 32011
0 32250 5 1 1 32249
0 32251 7 1 2 51367 32250
0 32252 7 1 2 32248 32251
0 32253 5 1 1 32252
0 32254 7 1 2 32185 32253
0 32255 5 1 1 32254
0 32256 7 1 2 66764 32255
0 32257 5 1 1 32256
0 32258 7 1 2 32183 32257
0 32259 5 1 1 32258
0 32260 7 1 2 52670 32259
0 32261 5 1 1 32260
0 32262 7 1 2 74682 76216
0 32263 5 1 1 32262
0 32264 7 1 2 60577 76111
0 32265 5 1 1 32264
0 32266 7 1 2 32263 32265
0 32267 5 1 1 32266
0 32268 7 1 2 52671 32267
0 32269 5 1 1 32268
0 32270 7 1 2 75972 76467
0 32271 5 1 1 32270
0 32272 7 1 2 32269 32271
0 32273 5 1 1 32272
0 32274 7 1 2 73675 32273
0 32275 5 1 1 32274
0 32276 7 1 2 63597 75545
0 32277 5 1 1 32276
0 32278 7 1 2 48777 71980
0 32279 5 1 1 32278
0 32280 7 1 2 32277 32279
0 32281 5 1 1 32280
0 32282 7 1 2 51086 32281
0 32283 5 1 1 32282
0 32284 7 1 2 75936 76468
0 32285 5 1 1 32284
0 32286 7 1 2 57329 75108
0 32287 7 1 2 75890 32286
0 32288 5 1 1 32287
0 32289 7 1 2 32285 32288
0 32290 5 1 1 32289
0 32291 7 1 2 73676 32290
0 32292 5 1 1 32291
0 32293 7 1 2 32283 32292
0 32294 5 1 1 32293
0 32295 7 1 2 53376 32294
0 32296 5 1 1 32295
0 32297 7 1 2 32275 32296
0 32298 5 1 1 32297
0 32299 7 1 2 53545 32298
0 32300 5 1 1 32299
0 32301 7 1 2 52672 75847
0 32302 5 1 1 32301
0 32303 7 1 2 71097 76776
0 32304 5 1 1 32303
0 32305 7 1 2 32302 32304
0 32306 5 1 1 32305
0 32307 7 1 2 49773 75192
0 32308 7 1 2 32306 32307
0 32309 5 1 1 32308
0 32310 7 1 2 32300 32309
0 32311 5 1 1 32310
0 32312 7 1 2 53699 32311
0 32313 5 1 1 32312
0 32314 7 1 2 73352 76198
0 32315 7 1 2 76470 32314
0 32316 5 1 1 32315
0 32317 7 1 2 32313 32316
0 32318 5 1 1 32317
0 32319 7 1 2 62174 32318
0 32320 5 1 1 32319
0 32321 7 1 2 75295 76013
0 32322 5 1 1 32321
0 32323 7 1 2 62362 75156
0 32324 7 1 2 77611 32323
0 32325 5 1 1 32324
0 32326 7 1 2 32322 32325
0 32327 5 1 1 32326
0 32328 7 1 2 55928 32327
0 32329 5 1 1 32328
0 32330 7 1 2 76015 75926
0 32331 5 1 1 32330
0 32332 7 1 2 32329 32331
0 32333 5 1 1 32332
0 32334 7 1 2 53377 32333
0 32335 5 1 1 32334
0 32336 7 1 2 76025 32335
0 32337 5 1 1 32336
0 32338 7 1 2 53700 32337
0 32339 5 1 1 32338
0 32340 7 1 2 73499 71197
0 32341 7 1 2 75332 32340
0 32342 5 1 1 32341
0 32343 7 1 2 32339 32342
0 32344 7 1 2 32320 32343
0 32345 5 1 1 32344
0 32346 7 1 2 75414 32345
0 32347 5 1 1 32346
0 32348 7 1 2 32261 32347
0 32349 7 1 2 32018 32348
0 32350 5 1 1 32349
0 32351 7 1 2 51598 32350
0 32352 5 1 1 32351
0 32353 7 4 2 48778 53701
0 32354 7 1 2 76098 77947
0 32355 5 1 1 32354
0 32356 7 1 2 69310 76150
0 32357 5 1 1 32356
0 32358 7 1 2 32355 32357
0 32359 5 1 1 32358
0 32360 7 1 2 55929 32359
0 32361 5 1 1 32360
0 32362 7 1 2 71076 76151
0 32363 5 1 1 32362
0 32364 7 1 2 32361 32363
0 32365 5 1 1 32364
0 32366 7 1 2 52445 32365
0 32367 5 1 1 32366
0 32368 7 1 2 66045 77726
0 32369 5 1 1 32368
0 32370 7 1 2 54726 32369
0 32371 5 1 1 32370
0 32372 7 1 2 52556 32371
0 32373 5 2 1 32372
0 32374 7 1 2 51087 77951
0 32375 5 1 1 32374
0 32376 7 1 2 76102 32375
0 32377 5 1 1 32376
0 32378 7 1 2 48779 32377
0 32379 5 1 1 32378
0 32380 7 2 2 61602 70449
0 32381 5 1 1 77953
0 32382 7 1 2 70387 32381
0 32383 5 1 1 32382
0 32384 7 1 2 59111 77171
0 32385 5 1 1 32384
0 32386 7 1 2 32383 32385
0 32387 5 1 1 32386
0 32388 7 1 2 56383 32387
0 32389 5 1 1 32388
0 32390 7 1 2 55930 77727
0 32391 5 1 1 32390
0 32392 7 1 2 56941 32391
0 32393 5 1 1 32392
0 32394 7 1 2 32389 32393
0 32395 5 1 1 32394
0 32396 7 1 2 48657 63520
0 32397 7 1 2 32395 32396
0 32398 5 1 1 32397
0 32399 7 1 2 32379 32398
0 32400 5 1 1 32399
0 32401 7 1 2 53702 32400
0 32402 5 1 1 32401
0 32403 7 1 2 32367 32402
0 32404 5 1 1 32403
0 32405 7 1 2 51368 32404
0 32406 5 1 1 32405
0 32407 7 1 2 54727 76044
0 32408 5 1 1 32407
0 32409 7 1 2 58565 63521
0 32410 7 1 2 77583 32409
0 32411 5 1 1 32410
0 32412 7 1 2 76093 32411
0 32413 5 1 1 32412
0 32414 7 1 2 54081 32413
0 32415 5 1 1 32414
0 32416 7 1 2 76075 32415
0 32417 7 1 2 32408 32416
0 32418 5 1 1 32417
0 32419 7 1 2 52673 32418
0 32420 5 1 1 32419
0 32421 7 1 2 70078 76117
0 32422 5 1 1 32421
0 32423 7 1 2 55931 71191
0 32424 7 1 2 32422 32423
0 32425 5 1 1 32424
0 32426 7 1 2 32420 32425
0 32427 5 1 1 32426
0 32428 7 1 2 66476 32427
0 32429 5 1 1 32428
0 32430 7 1 2 32406 32429
0 32431 5 1 1 32430
0 32432 7 1 2 53546 32431
0 32433 5 1 1 32432
0 32434 7 1 2 68588 75824
0 32435 5 1 1 32434
0 32436 7 2 2 63598 71575
0 32437 7 1 2 60124 75738
0 32438 7 1 2 70989 32437
0 32439 7 1 2 77955 32438
0 32440 5 1 1 32439
0 32441 7 1 2 32435 32440
0 32442 5 1 1 32441
0 32443 7 1 2 53002 32442
0 32444 5 1 1 32443
0 32445 7 1 2 53242 73157
0 32446 5 1 1 32445
0 32447 7 1 2 32444 32446
0 32448 5 1 1 32447
0 32449 7 1 2 55054 32448
0 32450 5 1 1 32449
0 32451 7 1 2 51369 77952
0 32452 5 1 1 32451
0 32453 7 1 2 71192 73092
0 32454 5 1 1 32453
0 32455 7 1 2 32452 32454
0 32456 5 1 1 32455
0 32457 7 1 2 62684 32456
0 32458 5 1 1 32457
0 32459 7 1 2 32450 32458
0 32460 5 1 1 32459
0 32461 7 1 2 52674 32460
0 32462 5 1 1 32461
0 32463 7 1 2 76106 32462
0 32464 5 1 1 32463
0 32465 7 1 2 53703 32464
0 32466 5 1 1 32465
0 32467 7 1 2 32433 32466
0 32468 5 1 1 32467
0 32469 7 1 2 53378 32468
0 32470 5 1 1 32469
0 32471 7 1 2 53704 24147
0 32472 5 1 1 32471
0 32473 7 1 2 32470 32472
0 32474 5 1 1 32473
0 32475 7 1 2 51599 32474
0 32476 5 1 1 32475
0 32477 7 1 2 75932 76250
0 32478 5 1 1 32477
0 32479 7 1 2 57330 76246
0 32480 5 1 1 32479
0 32481 7 1 2 32478 32480
0 32482 5 1 1 32481
0 32483 7 1 2 53705 32482
0 32484 5 1 1 32483
0 32485 7 5 2 49937 62492
0 32486 5 1 1 77957
0 32487 7 1 2 53003 73215
0 32488 5 1 1 32487
0 32489 7 1 2 55932 71060
0 32490 5 1 1 32489
0 32491 7 1 2 32488 32490
0 32492 5 1 1 32491
0 32493 7 1 2 77958 32492
0 32494 5 1 1 32493
0 32495 7 1 2 32484 32494
0 32496 5 1 1 32495
0 32497 7 1 2 51370 32496
0 32498 5 1 1 32497
0 32499 7 3 2 55375 68980
0 32500 7 1 2 76195 77962
0 32501 5 1 1 32500
0 32502 7 1 2 32498 32501
0 32503 5 1 1 32502
0 32504 7 1 2 51600 32503
0 32505 5 1 1 32504
0 32506 7 4 2 53379 68751
0 32507 7 2 2 66219 77965
0 32508 7 1 2 76634 77969
0 32509 5 1 1 32508
0 32510 7 1 2 32505 32509
0 32511 5 1 1 32510
0 32512 7 1 2 75212 32511
0 32513 5 1 1 32512
0 32514 7 1 2 53706 76240
0 32515 5 1 1 32514
0 32516 7 1 2 68719 70592
0 32517 7 2 2 76244 32516
0 32518 5 1 1 77971
0 32519 7 2 2 73371 75157
0 32520 5 1 1 77973
0 32521 7 1 2 49491 63798
0 32522 5 1 1 32521
0 32523 7 1 2 32520 32522
0 32524 5 1 1 32523
0 32525 7 1 2 76840 32524
0 32526 5 1 1 32525
0 32527 7 1 2 51371 73314
0 32528 7 1 2 75966 32527
0 32529 5 1 1 32528
0 32530 7 1 2 32526 32529
0 32531 5 1 1 32530
0 32532 7 1 2 52675 32531
0 32533 5 1 1 32532
0 32534 7 1 2 63210 76581
0 32535 5 1 1 32534
0 32536 7 1 2 23230 75860
0 32537 5 1 1 32536
0 32538 7 1 2 52557 32537
0 32539 5 1 1 32538
0 32540 7 1 2 32535 32539
0 32541 5 1 1 32540
0 32542 7 1 2 73372 32541
0 32543 5 1 1 32542
0 32544 7 1 2 32533 32543
0 32545 5 1 1 32544
0 32546 7 1 2 66765 32545
0 32547 5 1 1 32546
0 32548 7 8 2 52676 68808
0 32549 5 3 1 77975
0 32550 7 3 2 66280 77976
0 32551 7 1 2 71258 75944
0 32552 7 1 2 77986 32551
0 32553 5 1 1 32552
0 32554 7 1 2 32547 32553
0 32555 5 1 1 32554
0 32556 7 1 2 62175 32555
0 32557 5 1 1 32556
0 32558 7 1 2 53380 69244
0 32559 7 2 2 68504 32558
0 32560 5 1 1 77989
0 32561 7 1 2 75967 77990
0 32562 5 1 1 32561
0 32563 7 2 2 49774 66552
0 32564 5 1 1 77991
0 32565 7 1 2 32486 32564
0 32566 5 1 1 32565
0 32567 7 1 2 75956 32566
0 32568 5 1 1 32567
0 32569 7 1 2 32562 32568
0 32570 5 1 1 32569
0 32571 7 1 2 66609 32570
0 32572 5 1 1 32571
0 32573 7 1 2 68937 75048
0 32574 7 1 2 73842 32573
0 32575 7 1 2 76623 32574
0 32576 5 1 1 32575
0 32577 7 1 2 32572 32576
0 32578 7 1 2 32557 32577
0 32579 5 1 1 32578
0 32580 7 1 2 51601 32579
0 32581 5 1 1 32580
0 32582 7 1 2 32518 32581
0 32583 5 1 1 32582
0 32584 7 1 2 58544 32583
0 32585 5 1 1 32584
0 32586 7 1 2 32515 32585
0 32587 5 1 1 32586
0 32588 7 1 2 50260 32587
0 32589 5 1 1 32588
0 32590 7 1 2 32513 32589
0 32591 7 1 2 32476 32590
0 32592 5 1 1 32591
0 32593 7 1 2 50493 32592
0 32594 5 1 1 32593
0 32595 7 1 2 53707 75475
0 32596 5 1 1 32595
0 32597 7 1 2 57954 75322
0 32598 5 1 1 32597
0 32599 7 1 2 58695 32598
0 32600 5 1 1 32599
0 32601 7 1 2 75364 32600
0 32602 5 1 1 32601
0 32603 7 1 2 75324 76291
0 32604 5 1 1 32603
0 32605 7 1 2 75270 32604
0 32606 5 1 1 32605
0 32607 7 1 2 32602 32606
0 32608 5 1 1 32607
0 32609 7 1 2 49612 31917
0 32610 5 1 1 32609
0 32611 7 1 2 52558 75061
0 32612 7 1 2 32610 32611
0 32613 5 1 1 32612
0 32614 7 1 2 60125 75241
0 32615 7 1 2 77679 32614
0 32616 5 1 1 32615
0 32617 7 1 2 32613 32616
0 32618 5 1 1 32617
0 32619 7 1 2 58806 32618
0 32620 5 1 1 32619
0 32621 7 1 2 32608 32620
0 32622 5 1 1 32621
0 32623 7 1 2 51088 32622
0 32624 5 1 1 32623
0 32625 7 1 2 75415 75463
0 32626 5 1 1 32625
0 32627 7 1 2 56567 32626
0 32628 5 1 1 32627
0 32629 7 1 2 76437 32628
0 32630 5 1 1 32629
0 32631 7 1 2 32624 32630
0 32632 5 1 1 32631
0 32633 7 1 2 53708 32632
0 32634 5 1 1 32633
0 32635 7 1 2 60307 60102
0 32636 5 1 1 32635
0 32637 7 1 2 60947 32636
0 32638 5 1 1 32637
0 32639 7 1 2 59753 76852
0 32640 5 1 1 32639
0 32641 7 1 2 76974 32640
0 32642 5 1 1 32641
0 32643 7 1 2 32638 32642
0 32644 5 2 1 32643
0 32645 7 2 2 52321 77993
0 32646 5 1 1 77995
0 32647 7 1 2 71557 77977
0 32648 7 1 2 77996 32647
0 32649 5 1 1 32648
0 32650 7 1 2 32634 32649
0 32651 5 1 1 32650
0 32652 7 1 2 51602 32651
0 32653 5 1 1 32652
0 32654 7 1 2 73443 69316
0 32655 5 1 1 32654
0 32656 7 1 2 70929 32655
0 32657 5 1 1 32656
0 32658 7 1 2 52677 32657
0 32659 5 1 1 32658
0 32660 7 2 2 48780 68752
0 32661 7 1 2 55055 77997
0 32662 5 1 1 32661
0 32663 7 1 2 32659 32662
0 32664 5 1 1 32663
0 32665 7 1 2 58043 32664
0 32666 5 1 1 32665
0 32667 7 1 2 53709 75266
0 32668 5 1 1 32667
0 32669 7 1 2 32666 32668
0 32670 5 1 1 32669
0 32671 7 1 2 51603 32670
0 32672 5 1 1 32671
0 32673 7 2 2 59037 65731
0 32674 7 1 2 75305 77999
0 32675 5 1 1 32674
0 32676 7 1 2 32672 32675
0 32677 5 1 1 32676
0 32678 7 1 2 52322 32677
0 32679 5 1 1 32678
0 32680 7 2 2 68809 69411
0 32681 5 1 1 78001
0 32682 7 1 2 71506 78002
0 32683 5 1 1 32682
0 32684 7 1 2 32679 32683
0 32685 5 1 1 32684
0 32686 7 1 2 75223 32685
0 32687 5 1 1 32686
0 32688 7 1 2 51089 75261
0 32689 5 1 1 32688
0 32690 7 4 2 55056 58765
0 32691 7 1 2 52323 78003
0 32692 5 1 1 32691
0 32693 7 1 2 32689 32692
0 32694 5 1 1 32693
0 32695 7 1 2 71153 32694
0 32696 5 1 1 32695
0 32697 7 1 2 15610 32696
0 32698 5 1 1 32697
0 32699 7 1 2 49775 32698
0 32700 5 1 1 32699
0 32701 7 2 2 50818 60479
0 32702 5 1 1 78007
0 32703 7 1 2 57955 32702
0 32704 5 1 1 32703
0 32705 7 1 2 76264 32704
0 32706 5 1 1 32705
0 32707 7 1 2 32700 32706
0 32708 5 1 1 32707
0 32709 7 1 2 53126 32708
0 32710 5 1 1 32709
0 32711 7 1 2 51090 76506
0 32712 5 1 1 32711
0 32713 7 1 2 32710 32712
0 32714 5 1 1 32713
0 32715 7 1 2 75213 32714
0 32716 5 1 1 32715
0 32717 7 1 2 75874 75328
0 32718 5 1 1 32717
0 32719 7 1 2 61571 75326
0 32720 5 1 1 32719
0 32721 7 1 2 67334 32720
0 32722 5 1 1 32721
0 32723 7 1 2 71015 73773
0 32724 5 1 1 32723
0 32725 7 1 2 32722 32724
0 32726 5 1 1 32725
0 32727 7 1 2 75296 32726
0 32728 5 1 1 32727
0 32729 7 1 2 32718 32728
0 32730 7 1 2 32716 32729
0 32731 5 1 1 32730
0 32732 7 1 2 53710 32731
0 32733 5 1 1 32732
0 32734 7 1 2 61661 74667
0 32735 5 1 1 32734
0 32736 7 3 2 71077 73824
0 32737 5 1 1 78009
0 32738 7 2 2 70593 78010
0 32739 7 1 2 70760 78012
0 32740 7 1 2 32735 32739
0 32741 5 1 1 32740
0 32742 7 1 2 67735 15859
0 32743 5 1 1 32742
0 32744 7 1 2 75400 77959
0 32745 7 1 2 32743 32744
0 32746 7 1 2 75214 32745
0 32747 5 1 1 32746
0 32748 7 1 2 32741 32747
0 32749 7 1 2 32733 32748
0 32750 5 1 1 32749
0 32751 7 1 2 51604 32750
0 32752 5 1 1 32751
0 32753 7 1 2 58822 70602
0 32754 7 1 2 78000 32753
0 32755 7 1 2 75215 32754
0 32756 5 1 1 32755
0 32757 7 1 2 32752 32756
0 32758 5 1 1 32757
0 32759 7 1 2 50494 32758
0 32760 5 1 1 32759
0 32761 7 1 2 32687 32760
0 32762 7 1 2 32653 32761
0 32763 5 1 1 32762
0 32764 7 1 2 51372 32763
0 32765 5 1 1 32764
0 32766 7 1 2 32596 32765
0 32767 5 1 1 32766
0 32768 7 1 2 57037 32767
0 32769 5 1 1 32768
0 32770 7 2 2 76152 77966
0 32771 7 1 2 76377 78014
0 32772 5 1 1 32771
0 32773 7 1 2 53711 24645
0 32774 5 1 1 32773
0 32775 7 4 2 51373 69311
0 32776 7 1 2 51091 58445
0 32777 5 1 1 32776
0 32778 7 1 2 50261 77794
0 32779 5 1 1 32778
0 32780 7 1 2 32777 32779
0 32781 5 1 1 32780
0 32782 7 1 2 51973 32781
0 32783 5 1 1 32782
0 32784 7 1 2 71232 32783
0 32785 5 1 1 32784
0 32786 7 1 2 78016 32785
0 32787 5 1 1 32786
0 32788 7 1 2 68788 77737
0 32789 5 1 1 32788
0 32790 7 3 2 66281 71078
0 32791 5 3 1 78020
0 32792 7 1 2 66766 76763
0 32793 7 1 2 77931 32792
0 32794 5 1 1 32793
0 32795 7 1 2 78023 32794
0 32796 5 1 1 32795
0 32797 7 1 2 53004 32796
0 32798 5 1 1 32797
0 32799 7 1 2 32789 32798
0 32800 7 1 2 32787 32799
0 32801 5 1 1 32800
0 32802 7 1 2 52178 32801
0 32803 5 1 1 32802
0 32804 7 2 2 64792 66767
0 32805 5 1 1 78026
0 32806 7 1 2 49938 66713
0 32807 5 1 1 32806
0 32808 7 1 2 32805 32807
0 32809 5 1 1 32808
0 32810 7 1 2 50819 32809
0 32811 5 1 1 32810
0 32812 7 1 2 53005 78021
0 32813 5 1 1 32812
0 32814 7 1 2 73305 72842
0 32815 5 1 1 32814
0 32816 7 1 2 32813 32815
0 32817 5 2 1 32816
0 32818 7 1 2 62176 78028
0 32819 5 1 1 32818
0 32820 7 1 2 66824 68874
0 32821 5 1 1 32820
0 32822 7 1 2 78024 32821
0 32823 5 1 1 32822
0 32824 7 1 2 61529 32823
0 32825 5 1 1 32824
0 32826 7 1 2 32819 32825
0 32827 7 1 2 32811 32826
0 32828 7 1 2 32803 32827
0 32829 5 1 1 32828
0 32830 7 1 2 52446 32829
0 32831 5 1 1 32830
0 32832 7 1 2 66483 70158
0 32833 5 1 1 32832
0 32834 7 1 2 52559 6976
0 32835 5 1 1 32834
0 32836 7 1 2 32833 32835
0 32837 7 1 2 75141 32836
0 32838 5 1 1 32837
0 32839 7 2 2 51374 71307
0 32840 7 1 2 72731 78030
0 32841 7 1 2 62177 32840
0 32842 5 1 1 32841
0 32843 7 1 2 32838 32842
0 32844 7 1 2 32831 32843
0 32845 5 1 1 32844
0 32846 7 1 2 53243 32845
0 32847 5 1 1 32846
0 32848 7 1 2 74870 75630
0 32849 5 1 1 32848
0 32850 7 1 2 66685 32849
0 32851 5 1 1 32850
0 32852 7 3 2 52179 70254
0 32853 5 1 1 78032
0 32854 7 1 2 74832 78033
0 32855 5 1 1 32854
0 32856 7 1 2 50495 70496
0 32857 5 1 1 32856
0 32858 7 1 2 32855 32857
0 32859 5 1 1 32858
0 32860 7 1 2 75427 32859
0 32861 5 1 1 32860
0 32862 7 1 2 32851 32861
0 32863 5 1 1 32862
0 32864 7 1 2 54728 32863
0 32865 5 1 1 32864
0 32866 7 1 2 52560 75984
0 32867 5 1 1 32866
0 32868 7 1 2 68938 76698
0 32869 5 1 1 32868
0 32870 7 1 2 66906 32869
0 32871 5 1 1 32870
0 32872 7 1 2 60217 32871
0 32873 5 1 1 32872
0 32874 7 1 2 32867 32873
0 32875 7 1 2 32865 32874
0 32876 5 1 1 32875
0 32877 7 1 2 66477 32876
0 32878 5 1 1 32877
0 32879 7 4 2 51375 71079
0 32880 5 1 1 78035
0 32881 7 2 2 75302 78036
0 32882 7 1 2 76286 78039
0 32883 5 1 1 32882
0 32884 7 1 2 54729 76373
0 32885 5 1 1 32884
0 32886 7 1 2 78040 32885
0 32887 5 1 1 32886
0 32888 7 1 2 64335 63702
0 32889 5 1 1 32888
0 32890 7 1 2 52561 68888
0 32891 5 1 1 32890
0 32892 7 1 2 32889 32891
0 32893 5 1 1 32892
0 32894 7 1 2 66825 32893
0 32895 5 1 1 32894
0 32896 7 1 2 32887 32895
0 32897 5 1 1 32896
0 32898 7 1 2 62178 32897
0 32899 5 1 1 32898
0 32900 7 1 2 32883 32899
0 32901 7 1 2 32878 32900
0 32902 7 1 2 32847 32901
0 32903 5 1 1 32902
0 32904 7 1 2 53381 32903
0 32905 5 1 1 32904
0 32906 7 1 2 60218 76336
0 32907 5 1 1 32906
0 32908 7 1 2 71177 76640
0 32909 5 1 1 32908
0 32910 7 1 2 32907 32909
0 32911 5 1 1 32910
0 32912 7 1 2 55376 32911
0 32913 5 1 1 32912
0 32914 7 1 2 24110 32913
0 32915 5 1 1 32914
0 32916 7 1 2 53712 32915
0 32917 5 1 1 32916
0 32918 7 1 2 75945 78022
0 32919 7 1 2 76375 32918
0 32920 5 1 1 32919
0 32921 7 1 2 32917 32920
0 32922 5 1 1 32921
0 32923 7 1 2 62179 32922
0 32924 5 1 1 32923
0 32925 7 1 2 62140 63740
0 32926 7 1 2 73948 32925
0 32927 5 1 1 32926
0 32928 7 1 2 56642 60667
0 32929 5 1 1 32928
0 32930 7 1 2 49492 32929
0 32931 5 1 1 32930
0 32932 7 1 2 50820 32931
0 32933 5 1 1 32932
0 32934 7 1 2 70841 32933
0 32935 5 1 1 32934
0 32936 7 1 2 50496 68397
0 32937 7 1 2 32935 32936
0 32938 5 1 1 32937
0 32939 7 1 2 32927 32938
0 32940 5 1 1 32939
0 32941 7 1 2 66553 32940
0 32942 5 1 1 32941
0 32943 7 1 2 62099 73306
0 32944 7 1 2 76757 32943
0 32945 5 1 1 32944
0 32946 7 1 2 78025 32945
0 32947 5 1 1 32946
0 32948 7 1 2 70255 32947
0 32949 5 1 1 32948
0 32950 7 1 2 71896 77891
0 32951 5 1 1 32950
0 32952 7 1 2 52180 78029
0 32953 5 1 1 32952
0 32954 7 1 2 32951 32953
0 32955 7 1 2 32949 32954
0 32956 5 1 1 32955
0 32957 7 1 2 56227 32956
0 32958 5 1 1 32957
0 32959 7 1 2 49613 64209
0 32960 7 1 2 77963 32959
0 32961 5 1 1 32960
0 32962 7 1 2 32958 32961
0 32963 5 1 1 32962
0 32964 7 1 2 52562 32963
0 32965 5 1 1 32964
0 32966 7 1 2 32942 32965
0 32967 7 1 2 32924 32966
0 32968 7 1 2 32905 32967
0 32969 5 1 1 32968
0 32970 7 1 2 53547 32969
0 32971 5 1 1 32970
0 32972 7 1 2 55377 24663
0 32973 5 1 1 32972
0 32974 7 1 2 51376 76355
0 32975 5 1 1 32974
0 32976 7 1 2 68831 76361
0 32977 7 1 2 32975 32976
0 32978 7 1 2 32973 32977
0 32979 5 1 1 32978
0 32980 7 1 2 32971 32979
0 32981 5 1 1 32980
0 32982 7 1 2 52678 32981
0 32983 5 1 1 32982
0 32984 7 1 2 32774 32983
0 32985 5 1 1 32984
0 32986 7 1 2 51605 32985
0 32987 5 1 1 32986
0 32988 7 1 2 32772 32987
0 32989 5 1 1 32988
0 32990 7 1 2 57637 32989
0 32991 5 1 1 32990
0 32992 7 1 2 53713 24941
0 32993 5 1 1 32992
0 32994 7 2 2 58957 67886
0 32995 7 2 2 56136 76366
0 32996 5 1 1 78043
0 32997 7 1 2 51092 32996
0 32998 5 1 1 32997
0 32999 7 1 2 73266 74657
0 33000 7 1 2 69847 32999
0 33001 5 1 1 33000
0 33002 7 1 2 32998 33001
0 33003 5 1 1 33002
0 33004 7 1 2 56465 33003
0 33005 5 1 1 33004
0 33006 7 1 2 73254 73079
0 33007 5 1 1 33006
0 33008 7 1 2 33005 33007
0 33009 5 1 1 33008
0 33010 7 1 2 78041 33009
0 33011 5 1 1 33010
0 33012 7 1 2 53714 76423
0 33013 5 1 1 33012
0 33014 7 1 2 58044 71276
0 33015 5 1 1 33014
0 33016 7 1 2 56568 33015
0 33017 5 2 1 33016
0 33018 7 1 2 51974 59356
0 33019 7 1 2 73471 33018
0 33020 7 1 2 78045 33019
0 33021 5 1 1 33020
0 33022 7 1 2 33013 33021
0 33023 5 1 1 33022
0 33024 7 1 2 52181 33023
0 33025 5 1 1 33024
0 33026 7 1 2 67811 71311
0 33027 5 2 1 33026
0 33028 7 1 2 52447 66478
0 33029 7 1 2 75409 33028
0 33030 5 1 1 33029
0 33031 7 1 2 78047 33030
0 33032 5 1 1 33031
0 33033 7 1 2 59885 33032
0 33034 5 1 1 33033
0 33035 7 1 2 33025 33034
0 33036 5 1 1 33035
0 33037 7 1 2 58446 33036
0 33038 5 1 1 33037
0 33039 7 1 2 53715 76441
0 33040 5 1 1 33039
0 33041 7 1 2 53716 76439
0 33042 5 1 1 33041
0 33043 7 1 2 62236 78046
0 33044 5 1 1 33043
0 33045 7 1 2 73861 77509
0 33046 5 1 1 33045
0 33047 7 1 2 33044 33046
0 33048 5 1 1 33047
0 33049 7 1 2 68810 75336
0 33050 7 1 2 33048 33049
0 33051 5 1 1 33050
0 33052 7 1 2 33042 33051
0 33053 5 1 1 33052
0 33054 7 1 2 51377 33053
0 33055 5 1 1 33054
0 33056 7 1 2 33040 33055
0 33057 7 1 2 33038 33056
0 33058 5 1 1 33057
0 33059 7 1 2 57638 33058
0 33060 5 1 1 33059
0 33061 7 1 2 33011 33060
0 33062 7 1 2 32993 33061
0 33063 5 1 1 33062
0 33064 7 1 2 51606 33063
0 33065 5 1 1 33064
0 33066 7 1 2 73255 75262
0 33067 5 1 1 33066
0 33068 7 1 2 76461 33067
0 33069 5 1 1 33068
0 33070 7 1 2 76458 33069
0 33071 5 1 1 33070
0 33072 7 1 2 52679 76447
0 33073 5 1 1 33072
0 33074 7 1 2 33071 33073
0 33075 5 1 1 33074
0 33076 7 1 2 49776 33075
0 33077 5 1 1 33076
0 33078 7 1 2 52182 76282
0 33079 5 1 1 33078
0 33080 7 1 2 25029 33079
0 33081 5 1 1 33080
0 33082 7 1 2 63211 33081
0 33083 5 1 1 33082
0 33084 7 1 2 33077 33083
0 33085 5 1 1 33084
0 33086 7 1 2 53717 33085
0 33087 5 1 1 33086
0 33088 7 3 2 52183 52680
0 33089 7 3 2 63642 68811
0 33090 7 1 2 78049 78052
0 33091 7 1 2 75791 33090
0 33092 5 1 1 33091
0 33093 7 1 2 33087 33092
0 33094 5 1 1 33093
0 33095 7 1 2 51378 33094
0 33096 5 1 1 33095
0 33097 7 1 2 68481 77888
0 33098 7 1 2 76426 33097
0 33099 5 1 1 33098
0 33100 7 1 2 33096 33099
0 33101 5 1 1 33100
0 33102 7 1 2 51607 33101
0 33103 5 1 1 33102
0 33104 7 1 2 50497 76471
0 33105 7 1 2 77970 33104
0 33106 5 1 1 33105
0 33107 7 1 2 33103 33106
0 33108 5 1 1 33107
0 33109 7 1 2 60990 33108
0 33110 5 1 1 33109
0 33111 7 1 2 53718 76484
0 33112 5 1 1 33111
0 33113 7 3 2 66610 77978
0 33114 7 1 2 74833 75792
0 33115 5 1 1 33114
0 33116 7 1 2 56466 57639
0 33117 5 1 1 33116
0 33118 7 1 2 33115 33117
0 33119 5 1 1 33118
0 33120 7 1 2 78055 33119
0 33121 5 1 1 33120
0 33122 7 1 2 33112 33121
0 33123 5 1 1 33122
0 33124 7 1 2 51608 33123
0 33125 5 1 1 33124
0 33126 7 1 2 53719 76492
0 33127 5 1 1 33126
0 33128 7 1 2 33125 33127
0 33129 5 1 1 33128
0 33130 7 1 2 60342 33129
0 33131 5 1 1 33130
0 33132 7 3 2 53548 65732
0 33133 7 2 2 73294 78058
0 33134 7 1 2 76496 78061
0 33135 5 1 1 33134
0 33136 7 1 2 76498 78062
0 33137 5 1 1 33136
0 33138 7 1 2 52904 75989
0 33139 7 1 2 77928 33138
0 33140 7 1 2 76500 33139
0 33141 5 1 1 33140
0 33142 7 1 2 33137 33141
0 33143 5 1 1 33142
0 33144 7 1 2 57640 33143
0 33145 5 1 1 33144
0 33146 7 1 2 33135 33145
0 33147 7 1 2 33131 33146
0 33148 7 1 2 33110 33147
0 33149 7 1 2 33065 33148
0 33150 5 1 1 33149
0 33151 7 1 2 76381 33150
0 33152 5 1 1 33151
0 33153 7 1 2 53720 76544
0 33154 5 1 1 33153
0 33155 7 1 2 59893 72983
0 33156 5 2 1 33155
0 33157 7 1 2 73225 78063
0 33158 5 1 1 33157
0 33159 7 2 2 65298 59147
0 33160 5 2 1 78065
0 33161 7 1 2 33158 78067
0 33162 5 1 1 33161
0 33163 7 1 2 59176 78042
0 33164 7 1 2 33162 33163
0 33165 5 1 1 33164
0 33166 7 1 2 70137 73393
0 33167 5 1 1 33166
0 33168 7 1 2 53382 71016
0 33169 7 1 2 70108 33168
0 33170 5 1 1 33169
0 33171 7 1 2 33167 33170
0 33172 5 1 1 33171
0 33173 7 1 2 77987 33172
0 33174 5 1 1 33173
0 33175 7 1 2 33165 33174
0 33176 7 1 2 33154 33175
0 33177 5 1 1 33176
0 33178 7 1 2 51609 33177
0 33179 5 1 1 33178
0 33180 7 1 2 77619 77972
0 33181 5 1 1 33180
0 33182 7 1 2 66314 68484
0 33183 7 1 2 76548 33182
0 33184 5 1 1 33183
0 33185 7 1 2 33181 33184
0 33186 7 1 2 33179 33185
0 33187 5 1 1 33186
0 33188 7 1 2 62272 33187
0 33189 5 1 1 33188
0 33190 7 1 2 76632 78015
0 33191 5 1 1 33190
0 33192 7 1 2 53721 76607
0 33193 5 1 1 33192
0 33194 7 1 2 70256 70173
0 33195 7 1 2 77988 33194
0 33196 5 1 1 33195
0 33197 7 1 2 33193 33196
0 33198 5 1 1 33197
0 33199 7 1 2 57641 33198
0 33200 5 1 1 33199
0 33201 7 1 2 50498 58545
0 33202 7 1 2 77926 33201
0 33203 5 1 1 33202
0 33204 7 1 2 61530 77907
0 33205 5 1 1 33204
0 33206 7 1 2 33203 33205
0 33207 5 1 1 33206
0 33208 7 1 2 33207 78056
0 33209 5 1 1 33208
0 33210 7 1 2 53722 25529
0 33211 5 1 1 33210
0 33212 7 1 2 33209 33211
0 33213 7 1 2 33200 33212
0 33214 5 1 1 33213
0 33215 7 1 2 51610 33214
0 33216 5 1 1 33215
0 33217 7 1 2 33191 33216
0 33218 5 1 1 33217
0 33219 7 1 2 76561 33218
0 33220 5 1 1 33219
0 33221 7 1 2 76653 78017
0 33222 5 1 1 33221
0 33223 7 2 2 66479 76508
0 33224 5 1 1 78069
0 33225 7 1 2 33222 33224
0 33226 5 1 1 33225
0 33227 7 1 2 52184 33226
0 33228 5 1 1 33227
0 33229 7 1 2 49614 66480
0 33230 5 1 1 33229
0 33231 7 1 2 67887 77510
0 33232 7 1 2 70543 33231
0 33233 5 1 1 33232
0 33234 7 1 2 33230 33233
0 33235 5 1 1 33234
0 33236 7 1 2 75968 33235
0 33237 5 1 1 33236
0 33238 7 1 2 27528 78070
0 33239 5 1 1 33238
0 33240 7 1 2 33237 33239
0 33241 7 1 2 33228 33240
0 33242 5 1 1 33241
0 33243 7 1 2 51611 33242
0 33244 5 1 1 33243
0 33245 7 1 2 73121 69712
0 33246 7 1 2 76343 33245
0 33247 7 1 2 73275 77929
0 33248 7 1 2 33246 33247
0 33249 5 1 1 33248
0 33250 7 1 2 33244 33249
0 33251 5 1 1 33250
0 33252 7 1 2 51093 33251
0 33253 5 1 1 33252
0 33254 7 1 2 53723 76655
0 33255 5 1 1 33254
0 33256 7 1 2 33253 33255
0 33257 5 1 1 33256
0 33258 7 1 2 53549 33257
0 33259 5 1 1 33258
0 33260 7 2 2 72527 77964
0 33261 7 1 2 53244 75875
0 33262 7 1 2 78071 33261
0 33263 5 1 1 33262
0 33264 7 1 2 33259 33263
0 33265 5 1 1 33264
0 33266 7 1 2 52681 33265
0 33267 5 1 1 33266
0 33268 7 1 2 75869 78072
0 33269 5 1 1 33268
0 33270 7 1 2 33267 33269
0 33271 5 1 1 33270
0 33272 7 1 2 58546 33271
0 33273 5 1 1 33272
0 33274 7 1 2 66315 77967
0 33275 7 1 2 76635 33274
0 33276 5 1 1 33275
0 33277 7 1 2 48953 33276
0 33278 7 1 2 33273 33277
0 33279 7 1 2 33220 33278
0 33280 7 1 2 33189 33279
0 33281 7 1 2 33152 33280
0 33282 7 1 2 32991 33281
0 33283 7 1 2 32769 33282
0 33284 7 1 2 32594 33283
0 33285 7 1 2 32352 33284
0 33286 5 1 1 33285
0 33287 7 1 2 55659 33286
0 33288 7 1 2 31907 33287
0 33289 5 1 1 33288
0 33290 7 1 2 49493 77818
0 33291 5 1 1 33290
0 33292 7 1 2 62163 62785
0 33293 5 1 1 33292
0 33294 7 1 2 33291 33293
0 33295 5 1 1 33294
0 33296 7 1 2 48550 33295
0 33297 5 1 1 33296
0 33298 7 1 2 66016 76209
0 33299 5 1 1 33298
0 33300 7 1 2 33297 33299
0 33301 5 1 1 33300
0 33302 7 1 2 56569 33301
0 33303 5 1 1 33302
0 33304 7 1 2 61572 77832
0 33305 5 1 1 33304
0 33306 7 2 2 56384 61759
0 33307 5 2 1 78073
0 33308 7 1 2 58206 64220
0 33309 5 1 1 33308
0 33310 7 1 2 78075 33309
0 33311 7 1 2 33305 33310
0 33312 5 1 1 33311
0 33313 7 1 2 56137 33312
0 33314 5 1 1 33313
0 33315 7 1 2 58925 4328
0 33316 7 1 2 33314 33315
0 33317 5 1 1 33316
0 33318 7 1 2 53913 33317
0 33319 5 1 1 33318
0 33320 7 1 2 61064 77195
0 33321 5 1 1 33320
0 33322 7 1 2 72080 30998
0 33323 5 1 1 33322
0 33324 7 1 2 59227 33323
0 33325 5 1 1 33324
0 33326 7 1 2 33321 33325
0 33327 7 1 2 33319 33326
0 33328 5 1 1 33327
0 33329 7 1 2 58867 33328
0 33330 5 1 1 33329
0 33331 7 1 2 59505 59240
0 33332 5 1 1 33331
0 33333 7 1 2 3830 23454
0 33334 5 1 1 33333
0 33335 7 1 2 56138 33334
0 33336 5 1 1 33335
0 33337 7 1 2 58926 33336
0 33338 7 1 2 33332 33337
0 33339 5 1 1 33338
0 33340 7 1 2 68143 33339
0 33341 5 1 1 33340
0 33342 7 1 2 56228 74175
0 33343 5 1 1 33342
0 33344 7 1 2 62411 33343
0 33345 5 1 1 33344
0 33346 7 1 2 68160 33345
0 33347 7 1 2 63042 33346
0 33348 5 1 1 33347
0 33349 7 1 2 54730 33348
0 33350 5 1 1 33349
0 33351 7 1 2 56229 68152
0 33352 5 1 1 33351
0 33353 7 1 2 55933 59507
0 33354 5 2 1 33353
0 33355 7 1 2 68084 78077
0 33356 7 1 2 33352 33355
0 33357 5 1 1 33356
0 33358 7 1 2 58927 33357
0 33359 5 1 1 33358
0 33360 7 1 2 56755 33359
0 33361 5 1 1 33360
0 33362 7 1 2 33350 33361
0 33363 7 1 2 56385 60750
0 33364 5 1 1 33363
0 33365 7 1 2 68107 33364
0 33366 5 1 1 33365
0 33367 7 1 2 56139 33366
0 33368 5 1 1 33367
0 33369 7 1 2 62249 68097
0 33370 5 1 1 33369
0 33371 7 1 2 33368 33370
0 33372 5 1 1 33371
0 33373 7 1 2 60699 33372
0 33374 5 1 1 33373
0 33375 7 1 2 50499 66653
0 33376 5 1 1 33375
0 33377 7 1 2 62468 33376
0 33378 5 1 1 33377
0 33379 7 1 2 33374 33378
0 33380 7 1 2 33362 33379
0 33381 7 1 2 33341 33380
0 33382 7 1 2 33330 33381
0 33383 5 1 1 33382
0 33384 7 1 2 57956 33383
0 33385 5 1 1 33384
0 33386 7 1 2 33303 33385
0 33387 5 1 1 33386
0 33388 7 1 2 55057 33387
0 33389 5 1 1 33388
0 33390 7 1 2 57957 62783
0 33391 7 1 2 77716 33390
0 33392 5 1 1 33391
0 33393 7 1 2 33389 33392
0 33394 5 1 1 33393
0 33395 7 1 2 48781 33394
0 33396 5 1 1 33395
0 33397 7 1 2 1909 64020
0 33398 5 1 1 33397
0 33399 7 1 2 74016 33398
0 33400 5 1 1 33399
0 33401 7 1 2 58215 63974
0 33402 5 1 1 33401
0 33403 7 1 2 61872 33402
0 33404 5 1 1 33403
0 33405 7 1 2 33400 33404
0 33406 5 1 1 33405
0 33407 7 1 2 54376 33406
0 33408 5 1 1 33407
0 33409 7 2 2 53127 65430
0 33410 5 1 1 78079
0 33411 7 1 2 48420 33410
0 33412 5 1 1 33411
0 33413 7 1 2 77808 33412
0 33414 5 1 1 33413
0 33415 7 1 2 48223 33414
0 33416 5 1 1 33415
0 33417 7 1 2 64028 33416
0 33418 5 1 1 33417
0 33419 7 1 2 58868 33418
0 33420 5 1 1 33419
0 33421 7 1 2 57513 61611
0 33422 7 1 2 61852 33421
0 33423 5 1 1 33422
0 33424 7 1 2 33420 33423
0 33425 5 1 1 33424
0 33426 7 1 2 54731 33425
0 33427 5 1 1 33426
0 33428 7 1 2 33408 33427
0 33429 5 1 1 33428
0 33430 7 1 2 49494 33429
0 33431 5 1 1 33430
0 33432 7 1 2 65927 33431
0 33433 5 1 1 33432
0 33434 7 1 2 48551 33433
0 33435 5 1 1 33434
0 33436 7 1 2 67317 33435
0 33437 5 1 1 33436
0 33438 7 1 2 55058 33437
0 33439 5 1 1 33438
0 33440 7 1 2 49495 66872
0 33441 5 1 1 33440
0 33442 7 1 2 63288 66324
0 33443 5 1 1 33442
0 33444 7 1 2 52682 33443
0 33445 5 1 1 33444
0 33446 7 1 2 62788 33445
0 33447 5 1 1 33446
0 33448 7 1 2 33441 33447
0 33449 5 1 1 33448
0 33450 7 1 2 48224 33449
0 33451 5 1 1 33450
0 33452 7 1 2 63289 64902
0 33453 5 1 1 33452
0 33454 7 1 2 61315 33453
0 33455 5 1 1 33454
0 33456 7 1 2 61706 33455
0 33457 5 1 1 33456
0 33458 7 1 2 65089 1981
0 33459 5 1 1 33458
0 33460 7 1 2 62314 33459
0 33461 5 1 1 33460
0 33462 7 1 2 33457 33461
0 33463 7 1 2 33451 33462
0 33464 5 1 1 33463
0 33465 7 1 2 54377 33464
0 33466 5 1 1 33465
0 33467 7 1 2 66510 33466
0 33468 5 1 1 33467
0 33469 7 1 2 47966 33468
0 33470 5 1 1 33469
0 33471 7 1 2 59316 66545
0 33472 5 1 1 33471
0 33473 7 1 2 65517 59269
0 33474 5 1 1 33473
0 33475 7 1 2 33472 33474
0 33476 5 1 1 33475
0 33477 7 1 2 54082 33476
0 33478 5 1 1 33477
0 33479 7 1 2 33470 33478
0 33480 5 1 1 33479
0 33481 7 1 2 55798 33480
0 33482 5 1 1 33481
0 33483 7 2 2 47967 65250
0 33484 5 1 1 78081
0 33485 7 1 2 48225 73997
0 33486 5 1 1 33485
0 33487 7 1 2 33484 33486
0 33488 5 1 1 33487
0 33489 7 1 2 49127 33488
0 33490 5 1 1 33489
0 33491 7 3 2 49128 56386
0 33492 5 1 1 78083
0 33493 7 1 2 61163 58648
0 33494 7 1 2 33492 33493
0 33495 7 1 2 32205 33494
0 33496 7 1 2 33490 33495
0 33497 5 1 1 33496
0 33498 7 1 2 49231 33497
0 33499 5 1 1 33498
0 33500 7 1 2 58696 60776
0 33501 5 1 1 33500
0 33502 7 1 2 50821 72896
0 33503 7 1 2 76857 33502
0 33504 5 1 1 33503
0 33505 7 1 2 56387 33504
0 33506 5 1 1 33505
0 33507 7 1 2 33501 33506
0 33508 7 1 2 33499 33507
0 33509 5 1 1 33508
0 33510 7 1 2 56140 33509
0 33511 5 1 1 33510
0 33512 7 1 2 58869 73991
0 33513 5 1 1 33512
0 33514 7 1 2 59196 33513
0 33515 5 1 1 33514
0 33516 7 1 2 56756 33515
0 33517 5 1 1 33516
0 33518 7 1 2 59197 4537
0 33519 5 1 1 33518
0 33520 7 1 2 54378 33519
0 33521 5 1 1 33520
0 33522 7 1 2 33517 33521
0 33523 5 1 1 33522
0 33524 7 1 2 54732 33523
0 33525 5 1 1 33524
0 33526 7 1 2 74864 75742
0 33527 5 1 1 33526
0 33528 7 1 2 59228 33527
0 33529 5 1 1 33528
0 33530 7 1 2 56230 65239
0 33531 5 1 1 33530
0 33532 7 1 2 55059 33531
0 33533 5 1 1 33532
0 33534 7 1 2 58928 33533
0 33535 7 1 2 33529 33534
0 33536 7 1 2 33525 33535
0 33537 7 1 2 33511 33536
0 33538 5 1 1 33537
0 33539 7 1 2 48782 33538
0 33540 5 1 1 33539
0 33541 7 1 2 33482 33540
0 33542 7 1 2 33439 33541
0 33543 5 1 1 33542
0 33544 7 1 2 56570 33543
0 33545 5 1 1 33544
0 33546 7 1 2 61074 62449
0 33547 5 1 1 33546
0 33548 7 1 2 50822 59274
0 33549 5 2 1 33548
0 33550 7 1 2 61309 78086
0 33551 7 1 2 33547 33550
0 33552 5 1 1 33551
0 33553 7 1 2 56231 33552
0 33554 5 1 1 33553
0 33555 7 1 2 48783 74131
0 33556 7 1 2 33554 33555
0 33557 5 1 1 33556
0 33558 7 2 2 66155 66999
0 33559 5 1 1 78088
0 33560 7 1 2 66839 33559
0 33561 5 1 1 33560
0 33562 7 1 2 54733 33561
0 33563 5 1 1 33562
0 33564 7 2 2 56141 61313
0 33565 5 1 1 78090
0 33566 7 1 2 33563 33565
0 33567 5 1 1 33566
0 33568 7 1 2 56757 33567
0 33569 5 1 1 33568
0 33570 7 1 2 66915 74608
0 33571 5 1 1 33570
0 33572 7 1 2 33569 33571
0 33573 7 1 2 33557 33572
0 33574 5 1 1 33573
0 33575 7 1 2 56571 33574
0 33576 5 1 1 33575
0 33577 7 1 2 54734 74526
0 33578 5 1 1 33577
0 33579 7 1 2 68019 33578
0 33580 5 1 1 33579
0 33581 7 1 2 48226 33580
0 33582 5 1 1 33581
0 33583 7 1 2 4615 33582
0 33584 5 1 1 33583
0 33585 7 1 2 55060 33584
0 33586 5 1 1 33585
0 33587 7 1 2 56942 57289
0 33588 5 1 1 33587
0 33589 7 1 2 33586 33588
0 33590 5 1 1 33589
0 33591 7 1 2 56142 33590
0 33592 5 1 1 33591
0 33593 7 1 2 60931 58174
0 33594 7 1 2 60886 33593
0 33595 5 1 1 33594
0 33596 7 2 2 55061 68098
0 33597 5 2 1 78092
0 33598 7 1 2 71993 78094
0 33599 7 1 2 33595 33598
0 33600 5 1 1 33599
0 33601 7 1 2 56388 33600
0 33602 5 1 1 33601
0 33603 7 1 2 57514 78093
0 33604 5 1 1 33603
0 33605 7 1 2 57642 7262
0 33606 5 1 1 33605
0 33607 7 1 2 56943 33606
0 33608 5 1 1 33607
0 33609 7 1 2 33604 33608
0 33610 7 1 2 33602 33609
0 33611 5 1 1 33610
0 33612 7 1 2 54735 33611
0 33613 5 1 1 33612
0 33614 7 1 2 3861 33613
0 33615 7 1 2 33592 33614
0 33616 5 1 1 33615
0 33617 7 1 2 58116 33616
0 33618 5 1 1 33617
0 33619 7 1 2 33576 33618
0 33620 5 1 1 33619
0 33621 7 1 2 60700 33620
0 33622 5 1 1 33621
0 33623 7 1 2 3379 77719
0 33624 5 1 1 33623
0 33625 7 1 2 55062 33624
0 33626 5 1 1 33625
0 33627 7 1 2 49129 74536
0 33628 5 1 1 33627
0 33629 7 3 2 50500 61669
0 33630 5 3 1 78096
0 33631 7 1 2 62743 78097
0 33632 7 1 2 33628 33631
0 33633 5 1 1 33632
0 33634 7 1 2 56944 33633
0 33635 5 1 1 33634
0 33636 7 1 2 33626 33635
0 33637 5 1 1 33636
0 33638 7 1 2 49232 33637
0 33639 5 1 1 33638
0 33640 7 1 2 59711 64511
0 33641 5 1 1 33640
0 33642 7 1 2 3544 33641
0 33643 5 1 1 33642
0 33644 7 1 2 64221 33643
0 33645 5 1 1 33644
0 33646 7 1 2 50501 60859
0 33647 5 1 1 33646
0 33648 7 1 2 65320 33647
0 33649 5 1 1 33648
0 33650 7 1 2 33645 33649
0 33651 7 1 2 33639 33650
0 33652 5 1 1 33651
0 33653 7 1 2 54736 33652
0 33654 5 1 1 33653
0 33655 7 2 2 50502 16209
0 33656 5 3 1 78102
0 33657 7 1 2 49130 78104
0 33658 5 1 1 33657
0 33659 7 1 2 64222 61055
0 33660 5 1 1 33659
0 33661 7 1 2 33658 33660
0 33662 5 1 1 33661
0 33663 7 1 2 48227 33662
0 33664 5 1 1 33663
0 33665 7 1 2 60423 26742
0 33666 5 2 1 33665
0 33667 7 1 2 55799 78107
0 33668 5 1 1 33667
0 33669 7 1 2 59437 78099
0 33670 5 1 1 33669
0 33671 7 1 2 76741 33670
0 33672 7 1 2 33668 33671
0 33673 7 1 2 33664 33672
0 33674 5 1 1 33673
0 33675 7 1 2 7178 77358
0 33676 5 1 1 33675
0 33677 7 1 2 58697 33676
0 33678 5 1 1 33677
0 33679 7 1 2 56232 33678
0 33680 5 1 1 33679
0 33681 7 1 2 55063 33680
0 33682 7 1 2 33674 33681
0 33683 5 1 1 33682
0 33684 7 1 2 66151 74816
0 33685 5 1 1 33684
0 33686 7 1 2 55800 65823
0 33687 7 1 2 66788 33686
0 33688 5 1 1 33687
0 33689 7 1 2 33685 33688
0 33690 7 1 2 33683 33689
0 33691 7 1 2 33654 33690
0 33692 5 1 1 33691
0 33693 7 1 2 56143 33692
0 33694 5 1 1 33693
0 33695 7 1 2 65129 64672
0 33696 5 1 1 33695
0 33697 7 1 2 47968 33696
0 33698 5 1 1 33697
0 33699 7 1 2 65111 61760
0 33700 5 1 1 33699
0 33701 7 1 2 33698 33700
0 33702 5 1 1 33701
0 33703 7 1 2 48228 33702
0 33704 5 1 1 33703
0 33705 7 1 2 56945 61573
0 33706 7 1 2 63968 33705
0 33707 5 1 1 33706
0 33708 7 1 2 33704 33707
0 33709 5 1 1 33708
0 33710 7 1 2 55801 33709
0 33711 5 1 1 33710
0 33712 7 1 2 62868 74859
0 33713 5 1 1 33712
0 33714 7 2 2 47969 59229
0 33715 5 1 1 78109
0 33716 7 1 2 58216 33715
0 33717 5 1 1 33716
0 33718 7 1 2 49131 64663
0 33719 7 1 2 33717 33718
0 33720 5 1 1 33719
0 33721 7 1 2 33713 33720
0 33722 5 1 1 33721
0 33723 7 1 2 61662 33722
0 33724 5 1 1 33723
0 33725 7 1 2 65060 78110
0 33726 5 1 1 33725
0 33727 7 1 2 65130 33726
0 33728 5 1 1 33727
0 33729 7 1 2 74017 33728
0 33730 5 1 1 33729
0 33731 7 1 2 62869 66177
0 33732 5 1 1 33731
0 33733 7 1 2 3708 3109
0 33734 7 1 2 33732 33733
0 33735 7 1 2 33730 33734
0 33736 7 1 2 33724 33735
0 33737 7 1 2 33711 33736
0 33738 5 1 1 33737
0 33739 7 1 2 54379 33738
0 33740 5 1 1 33739
0 33741 7 1 2 54083 65251
0 33742 5 1 1 33741
0 33743 7 1 2 63101 33742
0 33744 5 1 1 33743
0 33745 7 1 2 47970 33744
0 33746 5 1 1 33745
0 33747 7 1 2 74149 33746
0 33748 5 1 1 33747
0 33749 7 1 2 56389 33748
0 33750 5 1 1 33749
0 33751 7 1 2 61663 66863
0 33752 5 1 1 33751
0 33753 7 1 2 48552 75730
0 33754 5 1 1 33753
0 33755 7 1 2 33752 33754
0 33756 5 1 1 33755
0 33757 7 1 2 47971 33756
0 33758 5 1 1 33757
0 33759 7 1 2 54737 71807
0 33760 5 1 1 33759
0 33761 7 1 2 56946 70425
0 33762 5 1 1 33761
0 33763 7 1 2 33760 33762
0 33764 7 1 2 33758 33763
0 33765 7 1 2 33750 33764
0 33766 5 1 1 33765
0 33767 7 1 2 55064 33766
0 33768 5 1 1 33767
0 33769 7 1 2 65112 74860
0 33770 5 1 1 33769
0 33771 7 1 2 65131 33770
0 33772 5 1 1 33771
0 33773 7 1 2 54738 2095
0 33774 7 1 2 33772 33773
0 33775 5 1 1 33774
0 33776 7 1 2 62196 76132
0 33777 7 1 2 59277 33776
0 33778 5 1 1 33777
0 33779 7 1 2 33775 33778
0 33780 7 1 2 33768 33779
0 33781 7 1 2 33740 33780
0 33782 7 1 2 33694 33781
0 33783 5 1 1 33782
0 33784 7 1 2 58117 33783
0 33785 5 1 1 33784
0 33786 7 1 2 65524 5398
0 33787 5 1 1 33786
0 33788 7 1 2 64006 33787
0 33789 5 1 1 33788
0 33790 7 1 2 48784 61204
0 33791 5 1 1 33790
0 33792 7 1 2 33789 33791
0 33793 5 1 1 33792
0 33794 7 1 2 48229 33793
0 33795 5 1 1 33794
0 33796 7 1 2 66511 33795
0 33797 5 1 1 33796
0 33798 7 1 2 56572 33797
0 33799 5 1 1 33798
0 33800 7 1 2 58207 65514
0 33801 5 1 1 33800
0 33802 7 1 2 56390 74469
0 33803 5 1 1 33802
0 33804 7 1 2 33801 33803
0 33805 5 1 1 33804
0 33806 7 1 2 56144 33805
0 33807 5 1 1 33806
0 33808 7 1 2 65535 20211
0 33809 5 1 1 33808
0 33810 7 1 2 57515 33809
0 33811 5 1 1 33810
0 33812 7 1 2 64908 33811
0 33813 7 1 2 33807 33812
0 33814 5 1 1 33813
0 33815 7 1 2 58118 33814
0 33816 5 1 1 33815
0 33817 7 1 2 33799 33816
0 33818 5 1 1 33817
0 33819 7 1 2 65561 33818
0 33820 5 1 1 33819
0 33821 7 1 2 62412 67000
0 33822 5 1 1 33821
0 33823 7 1 2 66840 33822
0 33824 5 1 1 33823
0 33825 7 1 2 56573 33824
0 33826 5 1 1 33825
0 33827 7 1 2 56391 71797
0 33828 5 1 1 33827
0 33829 7 1 2 60079 66976
0 33830 5 1 1 33829
0 33831 7 1 2 2827 64926
0 33832 5 1 1 33831
0 33833 7 1 2 48421 33832
0 33834 5 1 1 33833
0 33835 7 1 2 33830 33834
0 33836 7 1 2 33828 33835
0 33837 5 1 1 33836
0 33838 7 1 2 58119 33837
0 33839 5 1 1 33838
0 33840 7 1 2 33826 33839
0 33841 5 1 1 33840
0 33842 7 1 2 54739 33841
0 33843 5 1 1 33842
0 33844 7 1 2 56574 78091
0 33845 5 1 1 33844
0 33846 7 1 2 33843 33845
0 33847 5 1 1 33846
0 33848 7 1 2 64052 33847
0 33849 5 1 1 33848
0 33850 7 1 2 62835 33849
0 33851 7 1 2 33820 33850
0 33852 7 1 2 33785 33851
0 33853 7 1 2 33622 33852
0 33854 7 1 2 33545 33853
0 33855 5 1 1 33854
0 33856 7 1 2 49777 33855
0 33857 5 1 1 33856
0 33858 7 1 2 51379 33857
0 33859 7 1 2 33396 33858
0 33860 5 1 1 33859
0 33861 7 1 2 67220 76574
0 33862 5 1 1 33861
0 33863 7 1 2 75509 33862
0 33864 5 1 1 33863
0 33865 7 1 2 56758 33864
0 33866 5 1 1 33865
0 33867 7 1 2 65608 63582
0 33868 5 1 1 33867
0 33869 7 1 2 33866 33868
0 33870 5 1 1 33869
0 33871 7 1 2 56145 33870
0 33872 5 1 1 33871
0 33873 7 1 2 65434 60550
0 33874 7 1 2 75670 33873
0 33875 5 1 1 33874
0 33876 7 1 2 77851 33875
0 33877 5 1 1 33876
0 33878 7 1 2 48553 33877
0 33879 5 1 1 33878
0 33880 7 1 2 52683 77886
0 33881 5 2 1 33880
0 33882 7 1 2 33879 78111
0 33883 7 1 2 33872 33882
0 33884 5 1 1 33883
0 33885 7 1 2 62413 33884
0 33886 5 1 1 33885
0 33887 7 1 2 59270 77849
0 33888 5 1 1 33887
0 33889 7 1 2 48658 76575
0 33890 5 1 1 33889
0 33891 7 1 2 75510 33890
0 33892 5 2 1 33891
0 33893 7 1 2 62414 78113
0 33894 5 1 1 33893
0 33895 7 1 2 76187 77850
0 33896 5 1 1 33895
0 33897 7 2 2 57516 58643
0 33898 7 1 2 49233 76576
0 33899 7 1 2 78115 33898
0 33900 5 1 1 33899
0 33901 7 1 2 33896 33900
0 33902 7 1 2 33894 33901
0 33903 5 1 1 33902
0 33904 7 1 2 60932 33903
0 33905 5 1 1 33904
0 33906 7 1 2 33888 33905
0 33907 7 1 2 33886 33906
0 33908 5 1 1 33907
0 33909 7 1 2 55065 33908
0 33910 5 1 1 33909
0 33911 7 1 2 71112 77699
0 33912 5 1 1 33911
0 33913 7 1 2 52684 76154
0 33914 5 1 1 33913
0 33915 7 1 2 33912 33914
0 33916 5 3 1 33915
0 33917 7 1 2 54740 78117
0 33918 5 1 1 33917
0 33919 7 1 2 66807 74117
0 33920 7 1 2 57376 33919
0 33921 5 1 1 33920
0 33922 7 1 2 33918 33921
0 33923 5 1 1 33922
0 33924 7 1 2 56759 33923
0 33925 5 1 1 33924
0 33926 7 1 2 58045 62464
0 33927 5 1 1 33926
0 33928 7 1 2 56575 59148
0 33929 7 1 2 33927 33928
0 33930 5 1 1 33929
0 33931 7 1 2 33925 33930
0 33932 5 1 1 33931
0 33933 7 1 2 54380 33932
0 33934 5 1 1 33933
0 33935 7 1 2 57178 59149
0 33936 7 1 2 65598 33935
0 33937 5 1 1 33936
0 33938 7 1 2 33934 33937
0 33939 7 1 2 33910 33938
0 33940 5 1 1 33939
0 33941 7 1 2 60701 33940
0 33942 5 1 1 33941
0 33943 7 1 2 65904 75671
0 33944 5 1 1 33943
0 33945 7 1 2 57517 75694
0 33946 5 1 1 33945
0 33947 7 1 2 33944 33946
0 33948 5 1 1 33947
0 33949 7 1 2 56760 33948
0 33950 5 1 1 33949
0 33951 7 1 2 31956 33950
0 33952 5 1 1 33951
0 33953 7 1 2 54084 33952
0 33954 5 1 1 33953
0 33955 7 1 2 61482 77391
0 33956 5 1 1 33955
0 33957 7 1 2 33954 33956
0 33958 5 1 1 33957
0 33959 7 1 2 56392 33958
0 33960 5 1 1 33959
0 33961 7 1 2 61273 75439
0 33962 5 1 1 33961
0 33963 7 1 2 57518 57746
0 33964 5 2 1 33963
0 33965 7 1 2 53383 78120
0 33966 5 1 1 33965
0 33967 7 1 2 2488 56761
0 33968 7 1 2 33966 33967
0 33969 5 1 1 33968
0 33970 7 1 2 33962 33969
0 33971 5 1 1 33970
0 33972 7 1 2 54085 33971
0 33973 5 1 1 33972
0 33974 7 1 2 71792 75440
0 33975 5 1 1 33974
0 33976 7 1 2 33973 33975
0 33977 5 1 1 33976
0 33978 7 1 2 67221 33977
0 33979 5 1 1 33978
0 33980 7 2 2 50823 56762
0 33981 7 1 2 56947 77100
0 33982 7 1 2 78122 33981
0 33983 5 1 1 33982
0 33984 7 1 2 33979 33983
0 33985 7 1 2 33960 33984
0 33986 5 1 1 33985
0 33987 7 1 2 51094 33986
0 33988 5 1 1 33987
0 33989 7 1 2 61164 73949
0 33990 5 1 1 33989
0 33991 7 2 2 54741 33990
0 33992 7 1 2 53384 78124
0 33993 5 1 1 33992
0 33994 7 1 2 24232 33993
0 33995 5 1 1 33994
0 33996 7 1 2 48659 33995
0 33997 5 1 1 33996
0 33998 7 1 2 75365 23358
0 33999 5 1 1 33998
0 34000 7 1 2 56948 33999
0 34001 5 1 1 34000
0 34002 7 1 2 33997 34001
0 34003 5 1 1 34002
0 34004 7 1 2 51095 34003
0 34005 5 1 1 34004
0 34006 7 1 2 75504 78125
0 34007 5 1 1 34006
0 34008 7 1 2 34005 34007
0 34009 5 1 1 34008
0 34010 7 1 2 56146 34009
0 34011 5 1 1 34010
0 34012 7 1 2 59230 75582
0 34013 7 1 2 78108 34012
0 34014 5 1 1 34013
0 34015 7 1 2 34011 34014
0 34016 7 1 2 33988 34015
0 34017 5 1 1 34016
0 34018 7 1 2 55802 34017
0 34019 5 1 1 34018
0 34020 7 2 2 48660 75360
0 34021 5 2 1 78126
0 34022 7 1 2 62283 75441
0 34023 7 1 2 71951 34022
0 34024 5 1 1 34023
0 34025 7 1 2 78128 34024
0 34026 5 1 1 34025
0 34027 7 1 2 57179 34026
0 34028 5 1 1 34027
0 34029 7 1 2 5075 34028
0 34030 5 1 1 34029
0 34031 7 1 2 49132 34030
0 34032 5 1 1 34031
0 34033 7 2 2 48422 63948
0 34034 5 1 1 78130
0 34035 7 1 2 61406 77903
0 34036 7 1 2 78131 34035
0 34037 5 1 1 34036
0 34038 7 1 2 78129 34037
0 34039 5 1 1 34038
0 34040 7 1 2 57249 71408
0 34041 5 1 1 34040
0 34042 7 1 2 78127 34041
0 34043 5 1 1 34042
0 34044 7 1 2 50503 34043
0 34045 5 1 1 34044
0 34046 7 1 2 47972 34045
0 34047 7 1 2 34039 34046
0 34048 5 1 1 34047
0 34049 7 1 2 65124 75695
0 34050 5 1 1 34049
0 34051 7 1 2 34048 34050
0 34052 7 1 2 34032 34051
0 34053 5 1 1 34052
0 34054 7 1 2 51096 34053
0 34055 5 1 1 34054
0 34056 7 1 2 58870 57284
0 34057 5 1 1 34056
0 34058 7 1 2 68071 34057
0 34059 5 1 1 34058
0 34060 7 1 2 75696 34059
0 34061 5 1 1 34060
0 34062 7 1 2 28302 34061
0 34063 5 1 1 34062
0 34064 7 1 2 51097 34063
0 34065 5 1 1 34064
0 34066 7 1 2 23096 34065
0 34067 5 1 1 34066
0 34068 7 1 2 58943 34067
0 34069 5 1 1 34068
0 34070 7 1 2 59732 69485
0 34071 5 1 1 34070
0 34072 7 1 2 51098 75521
0 34073 5 1 1 34072
0 34074 7 2 2 75511 34073
0 34075 5 3 1 78132
0 34076 7 1 2 54742 78134
0 34077 7 1 2 34071 34076
0 34078 5 1 1 34077
0 34079 7 1 2 76172 34078
0 34080 5 1 1 34079
0 34081 7 1 2 59231 34080
0 34082 5 1 1 34081
0 34083 7 1 2 48661 75583
0 34084 5 1 1 34083
0 34085 7 1 2 49778 34084
0 34086 7 1 2 34082 34085
0 34087 7 1 2 34069 34086
0 34088 7 1 2 34055 34087
0 34089 7 1 2 67969 73209
0 34090 7 1 2 57104 34089
0 34091 7 1 2 69491 34090
0 34092 5 1 1 34091
0 34093 7 1 2 64056 66161
0 34094 5 1 1 34093
0 34095 7 2 2 50824 56393
0 34096 7 1 2 59283 78137
0 34097 7 1 2 34094 34096
0 34098 5 1 1 34097
0 34099 7 1 2 34092 34098
0 34100 5 1 1 34099
0 34101 7 1 2 57180 34100
0 34102 5 1 1 34101
0 34103 7 2 2 56394 78135
0 34104 5 2 1 78139
0 34105 7 1 2 62857 78140
0 34106 5 1 1 34105
0 34107 7 1 2 63310 66808
0 34108 5 1 1 34107
0 34109 7 1 2 34106 34108
0 34110 7 1 2 34102 34109
0 34111 5 1 1 34110
0 34112 7 1 2 56147 34111
0 34113 5 1 1 34112
0 34114 7 3 2 48785 63522
0 34115 5 1 1 78143
0 34116 7 1 2 48786 60219
0 34117 5 1 1 34116
0 34118 7 5 2 49615 56643
0 34119 7 1 2 58698 60860
0 34120 7 1 2 78146 34119
0 34121 5 1 1 34120
0 34122 7 1 2 34117 34121
0 34123 5 1 1 34122
0 34124 7 1 2 55934 34123
0 34125 5 1 1 34124
0 34126 7 1 2 49616 60578
0 34127 5 2 1 34126
0 34128 7 1 2 48787 78151
0 34129 5 1 1 34128
0 34130 7 1 2 34125 34129
0 34131 5 1 1 34130
0 34132 7 1 2 55066 34131
0 34133 5 1 1 34132
0 34134 7 1 2 34115 34133
0 34135 5 1 1 34134
0 34136 7 1 2 57331 34135
0 34137 5 1 1 34136
0 34138 7 1 2 34113 34137
0 34139 7 1 2 34088 34138
0 34140 7 1 2 74072 75232
0 34141 5 2 1 34140
0 34142 7 1 2 48788 71242
0 34143 5 1 1 34142
0 34144 7 1 2 78153 34143
0 34145 5 1 1 34144
0 34146 7 1 2 71137 34145
0 34147 5 1 1 34146
0 34148 7 1 2 58046 74077
0 34149 5 1 1 34148
0 34150 7 1 2 61131 72667
0 34151 5 1 1 34150
0 34152 7 1 2 34149 34151
0 34153 5 1 1 34152
0 34154 7 1 2 48789 34153
0 34155 5 1 1 34154
0 34156 7 1 2 34147 34155
0 34157 5 1 1 34156
0 34158 7 1 2 55067 34157
0 34159 5 1 1 34158
0 34160 7 2 2 57519 71029
0 34161 5 1 1 78155
0 34162 7 1 2 78144 34161
0 34163 5 1 1 34162
0 34164 7 1 2 34159 34163
0 34165 5 1 1 34164
0 34166 7 1 2 57038 34165
0 34167 5 1 1 34166
0 34168 7 1 2 59063 59150
0 34169 5 1 1 34168
0 34170 7 1 2 59480 78136
0 34171 5 1 1 34170
0 34172 7 1 2 34169 34171
0 34173 5 1 1 34172
0 34174 7 1 2 56148 34173
0 34175 5 1 1 34174
0 34176 7 1 2 57181 78118
0 34177 5 1 1 34176
0 34178 7 1 2 52685 75655
0 34179 5 1 1 34178
0 34180 7 1 2 28461 34179
0 34181 5 1 1 34180
0 34182 7 1 2 55068 34181
0 34183 5 1 1 34182
0 34184 7 1 2 34177 34183
0 34185 5 1 1 34184
0 34186 7 1 2 54743 34185
0 34187 5 1 1 34186
0 34188 7 1 2 34175 34187
0 34189 5 1 1 34188
0 34190 7 1 2 60248 34189
0 34191 5 1 1 34190
0 34192 7 1 2 52324 77654
0 34193 5 1 1 34192
0 34194 7 1 2 60100 63587
0 34195 5 1 1 34194
0 34196 7 1 2 34193 34195
0 34197 5 1 1 34196
0 34198 7 1 2 54086 72625
0 34199 5 1 1 34198
0 34200 7 1 2 70174 34199
0 34201 7 1 2 74019 34200
0 34202 7 1 2 34197 34201
0 34203 7 1 2 77662 34202
0 34204 5 1 1 34203
0 34205 7 1 2 59151 34204
0 34206 5 1 1 34205
0 34207 7 1 2 55935 63523
0 34208 5 2 1 34207
0 34209 7 4 2 53128 55069
0 34210 7 1 2 71243 78159
0 34211 5 1 1 34210
0 34212 7 1 2 63545 34211
0 34213 5 1 1 34212
0 34214 7 1 2 63524 76815
0 34215 5 1 1 34214
0 34216 7 1 2 48423 34215
0 34217 5 2 1 34216
0 34218 7 1 2 50262 78163
0 34219 7 1 2 34213 34218
0 34220 5 1 1 34219
0 34221 7 1 2 78157 34220
0 34222 5 1 1 34221
0 34223 7 1 2 50504 34222
0 34224 5 1 1 34223
0 34225 7 1 2 63546 77475
0 34226 5 1 1 34225
0 34227 7 1 2 53129 34226
0 34228 5 1 1 34227
0 34229 7 1 2 28745 34228
0 34230 5 1 1 34229
0 34231 7 1 2 56644 34230
0 34232 5 1 1 34231
0 34233 7 1 2 78158 34232
0 34234 5 1 1 34233
0 34235 7 1 2 60861 34234
0 34236 5 1 1 34235
0 34237 7 1 2 34224 34236
0 34238 7 1 2 34206 34237
0 34239 5 1 1 34238
0 34240 7 1 2 48790 34239
0 34241 5 1 1 34240
0 34242 7 1 2 34191 34241
0 34243 7 1 2 34167 34242
0 34244 7 1 2 34139 34243
0 34245 7 1 2 34019 34244
0 34246 7 1 2 33942 34245
0 34247 7 1 2 73993 34034
0 34248 5 1 1 34247
0 34249 7 1 2 47973 34248
0 34250 5 1 1 34249
0 34251 7 1 2 75713 34250
0 34252 5 1 1 34251
0 34253 7 1 2 49365 34252
0 34254 5 1 1 34253
0 34255 7 2 2 58175 72894
0 34256 5 1 1 78165
0 34257 7 1 2 34254 34256
0 34258 5 1 1 34257
0 34259 7 1 2 56395 34258
0 34260 5 1 1 34259
0 34261 7 1 2 65189 61132
0 34262 5 2 1 34261
0 34263 7 1 2 56949 78167
0 34264 5 1 1 34263
0 34265 7 1 2 34260 34264
0 34266 5 1 1 34265
0 34267 7 1 2 56576 34266
0 34268 5 1 1 34267
0 34269 7 1 2 57958 78168
0 34270 5 1 1 34269
0 34271 7 1 2 34268 34270
0 34272 5 1 1 34271
0 34273 7 1 2 59152 34272
0 34274 5 1 1 34273
0 34275 7 1 2 77714 75672
0 34276 5 1 1 34275
0 34277 7 1 2 56396 75697
0 34278 5 1 1 34277
0 34279 7 1 2 34276 34278
0 34280 5 1 1 34279
0 34281 7 1 2 58176 34280
0 34282 5 1 1 34281
0 34283 7 1 2 56397 77392
0 34284 5 1 1 34283
0 34285 7 1 2 34282 34284
0 34286 5 1 1 34285
0 34287 7 1 2 51099 34286
0 34288 5 1 1 34287
0 34289 7 1 2 56233 58191
0 34290 5 1 1 34289
0 34291 7 1 2 75584 34290
0 34292 5 1 1 34291
0 34293 7 1 2 34288 34292
0 34294 5 1 1 34293
0 34295 7 1 2 74770 34294
0 34296 5 1 1 34295
0 34297 7 1 2 66156 78119
0 34298 5 1 1 34297
0 34299 7 1 2 51100 77244
0 34300 5 1 1 34299
0 34301 7 1 2 78133 34300
0 34302 5 1 1 34301
0 34303 7 1 2 61664 58151
0 34304 7 1 2 34302 34303
0 34305 5 1 1 34304
0 34306 7 1 2 78141 34305
0 34307 5 1 1 34306
0 34308 7 1 2 58350 34307
0 34309 5 1 1 34308
0 34310 7 1 2 34298 34309
0 34311 5 1 1 34310
0 34312 7 1 2 54744 34311
0 34313 5 1 1 34312
0 34314 7 1 2 34296 34313
0 34315 7 1 2 34274 34314
0 34316 5 1 1 34315
0 34317 7 1 2 56763 34316
0 34318 5 1 1 34317
0 34319 7 2 2 59621 58138
0 34320 5 1 1 78169
0 34321 7 1 2 77812 34320
0 34322 5 1 1 34321
0 34323 7 1 2 54087 34322
0 34324 5 1 1 34323
0 34325 7 1 2 49234 74084
0 34326 5 1 1 34325
0 34327 7 1 2 34324 34326
0 34328 5 1 1 34327
0 34329 7 1 2 48230 34328
0 34330 5 1 1 34329
0 34331 7 1 2 61925 74512
0 34332 5 1 1 34331
0 34333 7 1 2 49235 34332
0 34334 5 1 1 34333
0 34335 7 1 2 49366 73998
0 34336 5 1 1 34335
0 34337 7 1 2 34334 34336
0 34338 5 1 1 34337
0 34339 7 1 2 48424 34338
0 34340 5 1 1 34339
0 34341 7 1 2 74709 34340
0 34342 7 1 2 34330 34341
0 34343 5 1 1 34342
0 34344 7 1 2 58871 34343
0 34345 5 1 1 34344
0 34346 7 1 2 57643 78098
0 34347 5 1 1 34346
0 34348 7 1 2 64007 34347
0 34349 5 1 1 34348
0 34350 7 1 2 48425 65252
0 34351 5 2 1 34350
0 34352 7 1 2 74794 78171
0 34353 5 1 1 34352
0 34354 7 1 2 60933 34353
0 34355 5 1 1 34354
0 34356 7 1 2 59622 62657
0 34357 5 1 1 34356
0 34358 7 1 2 34355 34357
0 34359 7 1 2 34349 34358
0 34360 5 1 1 34359
0 34361 7 1 2 48231 34360
0 34362 5 1 1 34361
0 34363 7 2 2 54745 78100
0 34364 5 2 1 78173
0 34365 7 1 2 48426 65871
0 34366 5 1 1 34365
0 34367 7 1 2 78175 34366
0 34368 5 1 1 34367
0 34369 7 1 2 49367 34368
0 34370 5 1 1 34369
0 34371 7 1 2 48427 58699
0 34372 5 1 1 34371
0 34373 7 1 2 34370 34372
0 34374 5 1 1 34373
0 34375 7 1 2 49236 34374
0 34376 5 1 1 34375
0 34377 7 1 2 68105 78172
0 34378 5 1 1 34377
0 34379 7 1 2 58184 65256
0 34380 5 1 1 34379
0 34381 7 1 2 62307 34380
0 34382 7 1 2 34378 34381
0 34383 5 1 1 34382
0 34384 7 2 2 60934 61574
0 34385 5 1 1 78177
0 34386 7 1 2 56149 65253
0 34387 5 1 1 34386
0 34388 7 1 2 61125 34387
0 34389 5 1 1 34388
0 34390 7 1 2 78178 34389
0 34391 5 1 1 34390
0 34392 7 1 2 56467 34391
0 34393 7 1 2 34383 34392
0 34394 7 1 2 34376 34393
0 34395 7 1 2 34362 34394
0 34396 7 1 2 34345 34395
0 34397 5 1 1 34396
0 34398 7 1 2 52686 34397
0 34399 5 1 1 34398
0 34400 7 1 2 52687 74787
0 34401 5 1 1 34400
0 34402 7 1 2 49237 75700
0 34403 7 1 2 63591 34402
0 34404 5 1 1 34403
0 34405 7 1 2 34401 34404
0 34406 5 1 1 34405
0 34407 7 1 2 53914 34406
0 34408 5 1 1 34407
0 34409 7 1 2 52688 61647
0 34410 5 1 1 34409
0 34411 7 1 2 34408 34410
0 34412 5 1 1 34411
0 34413 7 1 2 77020 34412
0 34414 5 1 1 34413
0 34415 7 1 2 34399 34414
0 34416 5 1 1 34415
0 34417 7 1 2 56398 34416
0 34418 5 1 1 34417
0 34419 7 1 2 50825 77720
0 34420 5 1 1 34419
0 34421 7 1 2 49617 34420
0 34422 5 1 1 34421
0 34423 7 2 2 58406 58700
0 34424 5 1 1 78179
0 34425 7 1 2 72538 78180
0 34426 5 2 1 34425
0 34427 7 1 2 34422 78181
0 34428 5 1 1 34427
0 34429 7 1 2 56764 34428
0 34430 5 1 1 34429
0 34431 7 1 2 68126 70504
0 34432 5 1 1 34431
0 34433 7 1 2 54746 60108
0 34434 5 1 1 34433
0 34435 7 1 2 60135 59295
0 34436 5 1 1 34435
0 34437 7 1 2 52563 57644
0 34438 7 1 2 34436 34437
0 34439 7 1 2 34434 34438
0 34440 7 1 2 34432 34439
0 34441 5 1 1 34440
0 34442 7 1 2 49618 34441
0 34443 5 1 1 34442
0 34444 7 1 2 53915 67320
0 34445 5 1 1 34444
0 34446 7 1 2 50826 34445
0 34447 5 1 1 34446
0 34448 7 1 2 49619 34447
0 34449 5 1 1 34448
0 34450 7 1 2 57776 65686
0 34451 5 2 1 34450
0 34452 7 1 2 53916 71846
0 34453 5 1 1 34452
0 34454 7 1 2 78183 34453
0 34455 5 1 1 34454
0 34456 7 1 2 48428 34455
0 34457 5 1 1 34456
0 34458 7 1 2 34449 34457
0 34459 5 1 1 34458
0 34460 7 1 2 58872 34459
0 34461 5 1 1 34460
0 34462 7 1 2 50505 59440
0 34463 5 1 1 34462
0 34464 7 1 2 61718 72612
0 34465 5 1 1 34464
0 34466 7 1 2 64037 34465
0 34467 5 1 1 34466
0 34468 7 1 2 34463 34467
0 34469 5 1 1 34468
0 34470 7 1 2 54747 58481
0 34471 7 1 2 78166 34470
0 34472 5 1 1 34471
0 34473 7 1 2 34469 34472
0 34474 7 1 2 34461 34473
0 34475 7 1 2 34443 34474
0 34476 7 1 2 34430 34475
0 34477 5 1 1 34476
0 34478 7 1 2 52689 34477
0 34479 5 1 1 34478
0 34480 7 1 2 74011 76297
0 34481 5 1 1 34480
0 34482 7 1 2 54381 34481
0 34483 5 1 1 34482
0 34484 7 1 2 61083 72911
0 34485 5 1 1 34484
0 34486 7 1 2 47974 61707
0 34487 7 1 2 75458 34486
0 34488 5 1 1 34487
0 34489 7 1 2 62291 34488
0 34490 7 1 2 34485 34489
0 34491 7 1 2 34483 34490
0 34492 5 1 1 34491
0 34493 7 1 2 52690 34492
0 34494 5 1 1 34493
0 34495 7 1 2 61677 62450
0 34496 5 1 1 34495
0 34497 7 1 2 56150 76577
0 34498 7 1 2 34496 34497
0 34499 5 1 1 34498
0 34500 7 1 2 34494 34499
0 34501 5 1 1 34500
0 34502 7 1 2 67222 34501
0 34503 5 1 1 34502
0 34504 7 1 2 76938 75688
0 34505 5 1 1 34504
0 34506 7 1 2 77852 34505
0 34507 5 1 1 34506
0 34508 7 1 2 48554 34507
0 34509 5 1 1 34508
0 34510 7 1 2 48232 78114
0 34511 5 1 1 34510
0 34512 7 1 2 78112 34511
0 34513 7 1 2 34509 34512
0 34514 5 1 1 34513
0 34515 7 1 2 52325 78080
0 34516 5 1 1 34515
0 34517 7 1 2 58873 34516
0 34518 7 1 2 34514 34517
0 34519 5 1 1 34518
0 34520 7 1 2 34503 34519
0 34521 7 1 2 34479 34520
0 34522 7 1 2 34418 34521
0 34523 5 1 1 34522
0 34524 7 1 2 55070 34523
0 34525 5 1 1 34524
0 34526 7 1 2 34318 34525
0 34527 7 1 2 34246 34526
0 34528 5 1 1 34527
0 34529 7 2 2 49238 77363
0 34530 5 1 1 78185
0 34531 7 1 2 61944 34530
0 34532 7 1 2 74280 34531
0 34533 5 1 1 34532
0 34534 7 1 2 55071 34533
0 34535 5 1 1 34534
0 34536 7 1 2 76562 34535
0 34537 5 1 1 34536
0 34538 7 2 2 54748 65913
0 34539 5 1 1 78187
0 34540 7 1 2 51101 34539
0 34541 5 2 1 34540
0 34542 7 1 2 49368 78189
0 34543 7 1 2 34537 34542
0 34544 5 1 1 34543
0 34545 7 1 2 64223 69885
0 34546 5 1 1 34545
0 34547 7 1 2 59463 34546
0 34548 5 1 1 34547
0 34549 7 1 2 48233 34548
0 34550 5 1 1 34549
0 34551 7 1 2 65916 34550
0 34552 5 1 1 34551
0 34553 7 1 2 55072 34552
0 34554 5 1 1 34553
0 34555 7 1 2 59508 74005
0 34556 5 1 1 34555
0 34557 7 1 2 60935 62308
0 34558 7 1 2 34556 34557
0 34559 5 1 1 34558
0 34560 7 1 2 49369 66338
0 34561 5 1 1 34560
0 34562 7 1 2 51102 34561
0 34563 7 1 2 34559 34562
0 34564 5 1 1 34563
0 34565 7 1 2 55073 59687
0 34566 5 3 1 34565
0 34567 7 1 2 50827 78191
0 34568 5 1 1 34567
0 34569 7 1 2 48429 34568
0 34570 7 1 2 34564 34569
0 34571 5 1 1 34570
0 34572 7 1 2 65314 74128
0 34573 5 2 1 34572
0 34574 7 1 2 78192 78194
0 34575 5 1 1 34574
0 34576 7 1 2 48234 34575
0 34577 5 1 1 34576
0 34578 7 1 2 64151 69886
0 34579 5 1 1 34578
0 34580 7 1 2 34577 34579
0 34581 5 1 1 34580
0 34582 7 1 2 61575 34581
0 34583 5 1 1 34582
0 34584 7 1 2 34571 34583
0 34585 7 1 2 34554 34584
0 34586 7 1 2 34544 34585
0 34587 5 1 1 34586
0 34588 7 1 2 56950 34587
0 34589 5 1 1 34588
0 34590 7 1 2 56951 78101
0 34591 5 1 1 34590
0 34592 7 1 2 4713 34591
0 34593 5 1 1 34592
0 34594 7 1 2 61026 34593
0 34595 5 1 1 34594
0 34596 7 1 2 64909 34595
0 34597 5 1 1 34596
0 34598 7 1 2 56765 34597
0 34599 5 1 1 34598
0 34600 7 1 2 59712 58482
0 34601 5 1 1 34600
0 34602 7 1 2 60400 60080
0 34603 5 1 1 34602
0 34604 7 1 2 34601 34603
0 34605 5 1 1 34604
0 34606 7 1 2 54749 34605
0 34607 5 1 1 34606
0 34608 7 1 2 68061 34607
0 34609 5 1 1 34608
0 34610 7 1 2 56952 34609
0 34611 5 1 1 34610
0 34612 7 1 2 17051 34611
0 34613 7 1 2 34599 34612
0 34614 5 1 1 34613
0 34615 7 1 2 58874 34614
0 34616 5 1 1 34615
0 34617 7 1 2 56953 74259
0 34618 5 1 1 34617
0 34619 7 1 2 67568 74129
0 34620 5 1 1 34619
0 34621 7 1 2 34618 34620
0 34622 5 1 1 34621
0 34623 7 1 2 56766 34622
0 34624 5 1 1 34623
0 34625 7 1 2 8586 78184
0 34626 5 1 1 34625
0 34627 7 1 2 55074 34626
0 34628 5 1 1 34627
0 34629 7 1 2 34624 34628
0 34630 5 1 1 34629
0 34631 7 1 2 60702 34630
0 34632 5 1 1 34631
0 34633 7 1 2 49239 27328
0 34634 5 1 1 34633
0 34635 7 1 2 34385 34634
0 34636 5 1 1 34635
0 34637 7 1 2 77810 34636
0 34638 5 1 1 34637
0 34639 7 1 2 64668 34638
0 34640 5 1 1 34639
0 34641 7 1 2 56954 34640
0 34642 5 1 1 34641
0 34643 7 1 2 49240 64658
0 34644 7 1 2 74333 34643
0 34645 5 1 1 34644
0 34646 7 1 2 34642 34645
0 34647 5 1 1 34646
0 34648 7 1 2 48235 34647
0 34649 5 1 1 34648
0 34650 7 1 2 34632 34649
0 34651 7 1 2 34616 34650
0 34652 5 1 1 34651
0 34653 7 1 2 48430 34652
0 34654 5 1 1 34653
0 34655 7 1 2 34589 34654
0 34656 5 1 1 34655
0 34657 7 1 2 58120 34656
0 34658 5 1 1 34657
0 34659 7 1 2 59161 68195
0 34660 5 1 1 34659
0 34661 7 1 2 53550 34660
0 34662 7 1 2 34658 34661
0 34663 5 1 1 34662
0 34664 7 1 2 34528 34663
0 34665 5 1 1 34664
0 34666 7 1 2 55803 63902
0 34667 5 1 1 34666
0 34668 7 1 2 53245 75608
0 34669 7 1 2 64093 34668
0 34670 7 1 2 69486 34669
0 34671 7 1 2 34667 34670
0 34672 5 1 1 34671
0 34673 7 1 2 48791 34672
0 34674 5 1 1 34673
0 34675 7 1 2 65171 62261
0 34676 7 1 2 64531 34675
0 34677 5 1 1 34676
0 34678 7 1 2 34674 34677
0 34679 5 1 1 34678
0 34680 7 1 2 54750 34679
0 34681 5 1 1 34680
0 34682 7 1 2 66512 34681
0 34683 5 1 1 34682
0 34684 7 1 2 48555 34683
0 34685 5 1 1 34684
0 34686 7 1 2 55936 72897
0 34687 5 1 1 34686
0 34688 7 1 2 55075 34687
0 34689 5 1 1 34688
0 34690 7 1 2 47975 62042
0 34691 5 1 1 34690
0 34692 7 1 2 63236 34691
0 34693 5 1 1 34692
0 34694 7 1 2 55804 34693
0 34695 5 1 1 34694
0 34696 7 1 2 62043 69326
0 34697 5 1 1 34696
0 34698 7 2 2 59590 69157
0 34699 5 1 1 78196
0 34700 7 1 2 34697 34699
0 34701 7 1 2 34695 34700
0 34702 5 1 1 34701
0 34703 7 1 2 54751 34702
0 34704 5 1 1 34703
0 34705 7 1 2 34689 34704
0 34706 5 1 1 34705
0 34707 7 1 2 57182 34706
0 34708 5 1 1 34707
0 34709 7 1 2 3542 65760
0 34710 5 1 1 34709
0 34711 7 1 2 48431 34710
0 34712 5 1 1 34711
0 34713 7 1 2 60424 133
0 34714 5 2 1 34713
0 34715 7 1 2 49496 78198
0 34716 5 1 1 34715
0 34717 7 1 2 34712 34716
0 34718 5 1 1 34717
0 34719 7 1 2 54752 34718
0 34720 5 1 1 34719
0 34721 7 1 2 64712 66157
0 34722 5 1 1 34721
0 34723 7 1 2 34720 34722
0 34724 5 1 1 34723
0 34725 7 1 2 74983 34724
0 34726 5 1 1 34725
0 34727 7 1 2 59450 73080
0 34728 5 1 1 34727
0 34729 7 1 2 54753 65482
0 34730 7 1 2 34728 34729
0 34731 5 1 1 34730
0 34732 7 1 2 14024 34731
0 34733 5 1 1 34732
0 34734 7 1 2 56151 34733
0 34735 5 1 1 34734
0 34736 7 1 2 66158 77073
0 34737 5 1 1 34736
0 34738 7 1 2 62029 34737
0 34739 5 1 1 34738
0 34740 7 1 2 54754 62044
0 34741 7 1 2 34739 34740
0 34742 5 1 1 34741
0 34743 7 1 2 51103 34742
0 34744 5 1 1 34743
0 34745 7 1 2 47976 73999
0 34746 5 1 1 34745
0 34747 7 1 2 54755 63385
0 34748 5 1 1 34747
0 34749 7 1 2 62033 34748
0 34750 7 1 2 34746 34749
0 34751 5 1 1 34750
0 34752 7 1 2 34744 34751
0 34753 5 1 1 34752
0 34754 7 1 2 34735 34753
0 34755 7 1 2 34726 34754
0 34756 7 1 2 34708 34755
0 34757 5 1 1 34756
0 34758 7 1 2 48792 34757
0 34759 5 1 1 34758
0 34760 7 1 2 34685 34759
0 34761 5 1 1 34760
0 34762 7 1 2 53551 34761
0 34763 5 1 1 34762
0 34764 7 1 2 48793 59232
0 34765 5 1 1 34764
0 34766 7 1 2 65125 70035
0 34767 5 1 1 34766
0 34768 7 1 2 34765 34767
0 34769 5 1 1 34768
0 34770 7 1 2 58701 34769
0 34771 5 1 1 34770
0 34772 7 1 2 48794 64518
0 34773 5 1 1 34772
0 34774 7 1 2 34771 34773
0 34775 5 1 1 34774
0 34776 7 1 2 53552 34775
0 34777 5 1 1 34776
0 34778 7 2 2 56152 59169
0 34779 7 1 2 78200 78089
0 34780 5 1 1 34779
0 34781 7 1 2 34777 34780
0 34782 5 1 1 34781
0 34783 7 1 2 56767 34782
0 34784 5 1 1 34783
0 34785 7 1 2 49133 59591
0 34786 5 1 1 34785
0 34787 7 1 2 50828 34786
0 34788 5 1 1 34787
0 34789 7 1 2 48795 34788
0 34790 5 1 1 34789
0 34791 7 1 2 54382 64946
0 34792 5 1 1 34791
0 34793 7 1 2 19114 34792
0 34794 5 1 1 34793
0 34795 7 1 2 57183 34794
0 34796 5 1 1 34795
0 34797 7 1 2 34790 34796
0 34798 5 1 1 34797
0 34799 7 1 2 74289 34798
0 34800 5 1 1 34799
0 34801 7 1 2 34784 34800
0 34802 5 1 1 34801
0 34803 7 1 2 60703 34802
0 34804 5 1 1 34803
0 34805 7 1 2 55076 78078
0 34806 5 1 1 34805
0 34807 7 1 2 59233 78174
0 34808 5 1 1 34807
0 34809 7 1 2 34806 34808
0 34810 5 1 1 34809
0 34811 7 1 2 48796 34810
0 34812 5 1 1 34811
0 34813 7 1 2 65126 65165
0 34814 5 1 1 34813
0 34815 7 1 2 34812 34814
0 34816 5 1 1 34815
0 34817 7 1 2 53553 34816
0 34818 5 1 1 34817
0 34819 7 1 2 57039 16943
0 34820 5 1 1 34819
0 34821 7 1 2 59170 74636
0 34822 7 1 2 34820 34821
0 34823 5 1 1 34822
0 34824 7 1 2 34818 34823
0 34825 5 1 1 34824
0 34826 7 1 2 58875 34825
0 34827 5 1 1 34826
0 34828 7 1 2 56234 64082
0 34829 5 1 1 34828
0 34830 7 1 2 68311 34829
0 34831 5 1 1 34830
0 34832 7 1 2 4977 34831
0 34833 5 1 1 34832
0 34834 7 1 2 56153 34833
0 34835 5 1 1 34834
0 34836 7 1 2 59234 68085
0 34837 5 1 1 34836
0 34838 7 1 2 51104 34837
0 34839 5 1 1 34838
0 34840 7 1 2 68312 34839
0 34841 5 1 1 34840
0 34842 7 1 2 64896 59153
0 34843 5 1 1 34842
0 34844 7 1 2 58944 59395
0 34845 5 1 1 34844
0 34846 7 1 2 69684 34845
0 34847 5 1 1 34846
0 34848 7 1 2 68144 34847
0 34849 5 1 1 34848
0 34850 7 1 2 34843 34849
0 34851 7 1 2 34841 34850
0 34852 7 1 2 34835 34851
0 34853 5 1 1 34852
0 34854 7 1 2 48797 34853
0 34855 5 1 1 34854
0 34856 7 1 2 34827 34855
0 34857 5 1 1 34856
0 34858 7 1 2 56768 34857
0 34859 5 1 1 34858
0 34860 7 1 2 65075 71789
0 34861 5 1 1 34860
0 34862 7 1 2 52691 34861
0 34863 5 1 1 34862
0 34864 7 1 2 74290 34863
0 34865 5 1 1 34864
0 34866 7 1 2 67001 78201
0 34867 5 1 1 34866
0 34868 7 1 2 34865 34867
0 34869 5 1 1 34868
0 34870 7 1 2 57184 34869
0 34871 5 1 1 34870
0 34872 7 2 2 47977 58945
0 34873 5 1 1 78202
0 34874 7 1 2 59154 78203
0 34875 5 1 1 34874
0 34876 7 1 2 53554 64519
0 34877 5 1 1 34876
0 34878 7 1 2 34875 34877
0 34879 5 1 1 34878
0 34880 7 1 2 48798 34879
0 34881 5 1 1 34880
0 34882 7 1 2 34871 34881
0 34883 5 1 1 34882
0 34884 7 1 2 64053 34883
0 34885 5 1 1 34884
0 34886 7 1 2 49134 74136
0 34887 5 1 1 34886
0 34888 7 1 2 71794 34887
0 34889 5 1 1 34888
0 34890 7 1 2 56399 34889
0 34891 5 1 1 34890
0 34892 7 1 2 62415 58876
0 34893 5 1 1 34892
0 34894 7 1 2 59694 77033
0 34895 7 1 2 34893 34894
0 34896 5 1 1 34895
0 34897 7 1 2 56955 34896
0 34898 5 1 1 34897
0 34899 7 1 2 59688 31511
0 34900 5 1 1 34899
0 34901 7 1 2 70935 69667
0 34902 7 1 2 77880 34901
0 34903 5 1 1 34902
0 34904 7 1 2 34900 34903
0 34905 5 2 1 34904
0 34906 7 1 2 60704 78204
0 34907 5 1 1 34906
0 34908 7 1 2 34898 34907
0 34909 7 1 2 34891 34908
0 34910 5 1 1 34909
0 34911 7 1 2 51105 75313
0 34912 7 1 2 34910 34911
0 34913 5 1 1 34912
0 34914 7 1 2 34885 34913
0 34915 7 1 2 34859 34914
0 34916 7 1 2 34804 34915
0 34917 7 1 2 34763 34916
0 34918 5 1 1 34917
0 34919 7 1 2 56577 34918
0 34920 5 1 1 34919
0 34921 7 2 2 68181 75619
0 34922 5 2 1 78206
0 34923 7 1 2 61104 74705
0 34924 5 1 1 34923
0 34925 7 1 2 47978 77862
0 34926 5 1 1 34925
0 34927 7 1 2 50829 34926
0 34928 5 1 1 34927
0 34929 7 1 2 59623 34928
0 34930 5 1 1 34929
0 34931 7 1 2 34924 34930
0 34932 5 1 1 34931
0 34933 7 1 2 55805 34932
0 34934 5 1 1 34933
0 34935 7 1 2 48236 78186
0 34936 5 1 1 34935
0 34937 7 1 2 68868 34936
0 34938 5 1 1 34937
0 34939 7 1 2 54756 34938
0 34940 5 1 1 34939
0 34941 7 1 2 62131 76210
0 34942 5 1 1 34941
0 34943 7 1 2 34940 34942
0 34944 5 1 1 34943
0 34945 7 1 2 59689 34944
0 34946 5 1 1 34945
0 34947 7 1 2 64480 61035
0 34948 5 1 1 34947
0 34949 7 1 2 54383 62441
0 34950 5 1 1 34949
0 34951 7 1 2 57758 34950
0 34952 5 1 1 34951
0 34953 7 1 2 60060 34952
0 34954 5 1 1 34953
0 34955 7 1 2 34948 34954
0 34956 5 1 1 34955
0 34957 7 1 2 58407 34956
0 34958 5 1 1 34957
0 34959 7 1 2 61823 77828
0 34960 5 1 1 34959
0 34961 7 1 2 63156 58920
0 34962 7 1 2 63958 34961
0 34963 5 1 1 34962
0 34964 7 1 2 54384 34963
0 34965 5 1 1 34964
0 34966 7 1 2 34960 34965
0 34967 5 1 1 34966
0 34968 7 1 2 49370 34967
0 34969 5 1 1 34968
0 34970 7 1 2 34958 34969
0 34971 7 1 2 34946 34970
0 34972 7 1 2 34934 34971
0 34973 5 1 1 34972
0 34974 7 1 2 55077 59118
0 34975 7 1 2 34973 34974
0 34976 5 1 1 34975
0 34977 7 1 2 78208 34976
0 34978 5 1 1 34977
0 34979 7 1 2 56400 34978
0 34980 5 1 1 34979
0 34981 7 1 2 63765 70512
0 34982 5 2 1 34981
0 34983 7 1 2 49371 78210
0 34984 5 1 1 34983
0 34985 7 1 2 77666 34984
0 34986 5 1 1 34985
0 34987 7 1 2 63290 74291
0 34988 7 1 2 61367 34987
0 34989 5 1 1 34988
0 34990 7 1 2 78209 34989
0 34991 5 1 1 34990
0 34992 7 1 2 34986 34991
0 34993 5 1 1 34992
0 34994 7 1 2 48432 78207
0 34995 5 1 1 34994
0 34996 7 1 2 67485 76600
0 34997 5 1 1 34996
0 34998 7 1 2 34995 34997
0 34999 5 1 1 34998
0 35000 7 2 2 59661 61046
0 35001 5 1 1 78212
0 35002 7 1 2 70544 78213
0 35003 5 1 1 35002
0 35004 7 1 2 34999 35003
0 35005 5 1 1 35004
0 35006 7 1 2 55378 35005
0 35007 7 1 2 34993 35006
0 35008 7 1 2 34980 35007
0 35009 7 1 2 34920 35008
0 35010 7 1 2 34665 35009
0 35011 5 1 1 35010
0 35012 7 1 2 55546 35011
0 35013 7 1 2 33860 35012
0 35014 5 1 1 35013
0 35015 7 1 2 58877 16147
0 35016 5 1 1 35015
0 35017 7 2 2 65917 35016
0 35018 7 1 2 77018 78214
0 35019 5 1 1 35018
0 35020 7 1 2 49372 35019
0 35021 5 1 1 35020
0 35022 7 1 2 26754 35021
0 35023 5 1 1 35022
0 35024 7 1 2 48433 35023
0 35025 5 1 1 35024
0 35026 7 1 2 64183 58878
0 35027 5 1 1 35026
0 35028 7 1 2 35025 35027
0 35029 5 1 1 35028
0 35030 7 1 2 56401 35029
0 35031 5 1 1 35030
0 35032 7 1 2 32853 78105
0 35033 5 1 1 35032
0 35034 7 1 2 7056 35033
0 35035 5 1 1 35034
0 35036 7 1 2 58879 35035
0 35037 5 2 1 35036
0 35038 7 1 2 62391 61828
0 35039 5 2 1 35038
0 35040 7 1 2 54385 78218
0 35041 5 1 1 35040
0 35042 7 1 2 57645 35041
0 35043 7 1 2 78216 35042
0 35044 5 1 1 35043
0 35045 7 1 2 56956 35044
0 35046 5 1 1 35045
0 35047 7 1 2 53246 74513
0 35048 5 1 1 35047
0 35049 7 1 2 48556 35048
0 35050 5 1 1 35049
0 35051 7 1 2 6038 35050
0 35052 5 1 1 35051
0 35053 7 1 2 62661 68111
0 35054 5 1 1 35053
0 35055 7 1 2 61785 35054
0 35056 5 1 1 35055
0 35057 7 1 2 62262 74758
0 35058 5 1 1 35057
0 35059 7 2 2 35056 35058
0 35060 5 1 1 78220
0 35061 7 1 2 35052 35060
0 35062 5 1 1 35061
0 35063 7 1 2 64257 78084
0 35064 5 1 1 35063
0 35065 7 1 2 77651 35064
0 35066 5 1 1 35065
0 35067 7 1 2 61576 35066
0 35068 5 1 1 35067
0 35069 7 1 2 62132 65272
0 35070 5 1 1 35069
0 35071 7 1 2 77652 35070
0 35072 5 1 1 35071
0 35073 7 1 2 68121 35072
0 35074 5 1 1 35073
0 35075 7 1 2 35068 35074
0 35076 5 1 1 35075
0 35077 7 1 2 68166 35076
0 35078 5 1 1 35077
0 35079 7 1 2 35062 35078
0 35080 7 1 2 35046 35079
0 35081 7 1 2 35031 35080
0 35082 5 1 1 35081
0 35083 7 1 2 56578 35082
0 35084 5 1 1 35083
0 35085 7 1 2 50506 78221
0 35086 5 1 1 35085
0 35087 7 1 2 61781 61960
0 35088 5 1 1 35087
0 35089 7 1 2 35086 35088
0 35090 5 1 1 35089
0 35091 7 1 2 49373 58330
0 35092 5 1 1 35091
0 35093 7 1 2 56235 35092
0 35094 7 1 2 78217 35093
0 35095 7 1 2 35090 35094
0 35096 5 1 1 35095
0 35097 7 1 2 57959 35096
0 35098 5 1 1 35097
0 35099 7 1 2 35084 35098
0 35100 5 1 1 35099
0 35101 7 1 2 54757 35100
0 35102 5 1 1 35101
0 35103 7 1 2 63311 28935
0 35104 5 1 1 35103
0 35105 7 2 2 49620 77579
0 35106 5 1 1 78222
0 35107 7 1 2 57305 78223
0 35108 5 1 1 35107
0 35109 7 1 2 35104 35108
0 35110 5 1 1 35109
0 35111 7 1 2 54386 35110
0 35112 5 1 1 35111
0 35113 7 1 2 64298 35112
0 35114 7 1 2 35102 35113
0 35115 5 1 1 35114
0 35116 7 1 2 62930 66680
0 35117 7 1 2 35115 35116
0 35118 5 1 1 35117
0 35119 7 1 2 35014 35118
0 35120 5 1 1 35119
0 35121 7 1 2 73317 35120
0 35122 5 1 1 35121
0 35123 7 1 2 58721 75728
0 35124 5 2 1 35123
0 35125 7 2 2 62878 77570
0 35126 7 1 2 49241 78226
0 35127 5 1 1 35126
0 35128 7 2 2 54758 65020
0 35129 5 1 1 78228
0 35130 7 1 2 60425 78229
0 35131 5 1 1 35130
0 35132 7 1 2 35127 35131
0 35133 7 1 2 78224 35132
0 35134 5 1 1 35133
0 35135 7 1 2 57520 35134
0 35136 5 1 1 35135
0 35137 7 2 2 57834 65422
0 35138 5 1 1 78230
0 35139 7 1 2 50263 78231
0 35140 5 1 1 35139
0 35141 7 2 2 35136 35140
0 35142 5 1 1 78232
0 35143 7 2 2 49497 77058
0 35144 5 1 1 78234
0 35145 7 1 2 78233 35144
0 35146 5 1 1 35145
0 35147 7 1 2 51106 35146
0 35148 5 1 1 35147
0 35149 7 1 2 65263 66181
0 35150 5 1 1 35149
0 35151 7 1 2 52692 35150
0 35152 5 1 1 35151
0 35153 7 1 2 60763 70932
0 35154 5 2 1 35153
0 35155 7 1 2 57306 78236
0 35156 5 1 1 35155
0 35157 7 1 2 71131 35156
0 35158 5 1 1 35157
0 35159 7 3 2 49498 76367
0 35160 5 4 1 78238
0 35161 7 1 2 58829 77003
0 35162 5 1 1 35161
0 35163 7 1 2 48662 35162
0 35164 5 1 1 35163
0 35165 7 1 2 78241 35164
0 35166 5 2 1 35165
0 35167 7 1 2 56402 10279
0 35168 5 1 1 35167
0 35169 7 1 2 70974 35168
0 35170 5 1 1 35169
0 35171 7 1 2 54759 35170
0 35172 7 1 2 78245 35171
0 35173 7 1 2 35158 35172
0 35174 5 1 1 35173
0 35175 7 1 2 62613 70642
0 35176 5 1 1 35175
0 35177 7 1 2 56403 71007
0 35178 5 1 1 35177
0 35179 7 1 2 54387 35178
0 35180 5 1 1 35179
0 35181 7 1 2 50830 35180
0 35182 7 1 2 35176 35181
0 35183 5 1 1 35182
0 35184 7 1 2 55078 35183
0 35185 7 1 2 35174 35184
0 35186 5 1 1 35185
0 35187 7 1 2 35152 35186
0 35188 7 1 2 35148 35187
0 35189 5 1 1 35188
0 35190 7 1 2 68812 35189
0 35191 5 1 1 35190
0 35192 7 1 2 49242 59521
0 35193 5 1 1 35192
0 35194 7 1 2 23427 35129
0 35195 7 1 2 35193 35194
0 35196 5 1 1 35195
0 35197 7 1 2 57521 35196
0 35198 5 1 1 35197
0 35199 7 1 2 35138 35198
0 35200 5 1 1 35199
0 35201 7 1 2 65573 77948
0 35202 7 1 2 35200 35201
0 35203 5 1 1 35202
0 35204 7 1 2 35191 35203
0 35205 5 1 1 35204
0 35206 7 1 2 49621 35205
0 35207 5 1 1 35206
0 35208 7 3 2 52448 66353
0 35209 5 2 1 78247
0 35210 7 2 2 55079 78250
0 35211 5 1 1 78252
0 35212 7 1 2 60761 60889
0 35213 7 1 2 60897 35212
0 35214 5 1 1 35213
0 35215 7 1 2 67727 78237
0 35216 7 1 2 35214 35215
0 35217 5 1 1 35216
0 35218 7 1 2 52326 35217
0 35219 5 1 1 35218
0 35220 7 1 2 78253 35219
0 35221 5 1 1 35220
0 35222 7 1 2 64955 35221
0 35223 5 1 1 35222
0 35224 7 1 2 50831 69663
0 35225 5 2 1 35224
0 35226 7 2 2 66204 78254
0 35227 7 1 2 58047 78193
0 35228 5 1 1 35227
0 35229 7 1 2 51107 75461
0 35230 5 1 1 35229
0 35231 7 1 2 35228 35230
0 35232 7 1 2 78256 35231
0 35233 7 1 2 55080 10030
0 35234 5 1 1 35233
0 35235 7 1 2 50832 35234
0 35236 5 1 1 35235
0 35237 7 1 2 61353 64021
0 35238 5 1 1 35237
0 35239 7 1 2 35236 35238
0 35240 7 1 2 35232 35239
0 35241 7 1 2 48663 78239
0 35242 5 1 1 35241
0 35243 7 1 2 53385 35242
0 35244 5 1 1 35243
0 35245 7 1 2 78246 35244
0 35246 7 1 2 35240 35245
0 35247 7 1 2 35223 35246
0 35248 5 1 1 35247
0 35249 7 1 2 49779 35248
0 35250 5 1 1 35249
0 35251 7 1 2 62342 61126
0 35252 5 1 1 35251
0 35253 7 1 2 4288 35252
0 35254 5 1 1 35253
0 35255 7 1 2 67202 35254
0 35256 5 1 1 35255
0 35257 7 1 2 69782 35256
0 35258 5 1 1 35257
0 35259 7 1 2 35250 35258
0 35260 5 1 1 35259
0 35261 7 1 2 52693 35260
0 35262 5 1 1 35261
0 35263 7 1 2 67223 35142
0 35264 5 1 1 35263
0 35265 7 1 2 48664 78235
0 35266 5 1 1 35265
0 35267 7 1 2 35264 35266
0 35268 5 1 1 35267
0 35269 7 1 2 51108 35268
0 35270 5 1 1 35269
0 35271 7 1 2 61056 71802
0 35272 7 1 2 72843 35271
0 35273 5 1 1 35272
0 35274 7 1 2 74508 78170
0 35275 5 1 1 35274
0 35276 7 1 2 67203 35275
0 35277 5 1 1 35276
0 35278 7 1 2 50833 60800
0 35279 7 1 2 35277 35278
0 35280 5 1 1 35279
0 35281 7 1 2 35273 35280
0 35282 5 1 1 35281
0 35283 7 1 2 55081 35282
0 35284 5 1 1 35283
0 35285 7 1 2 64351 71134
0 35286 5 1 1 35285
0 35287 7 1 2 48799 35286
0 35288 5 1 1 35287
0 35289 7 2 2 51109 67224
0 35290 7 1 2 58408 78188
0 35291 7 1 2 78258 35290
0 35292 5 1 1 35291
0 35293 7 1 2 35288 35292
0 35294 7 1 2 35284 35293
0 35295 5 1 1 35294
0 35296 7 1 2 53386 35295
0 35297 5 1 1 35296
0 35298 7 1 2 51110 63102
0 35299 5 1 1 35298
0 35300 7 1 2 48665 35299
0 35301 5 1 1 35300
0 35302 7 1 2 63471 35301
0 35303 5 1 1 35302
0 35304 7 1 2 78257 35303
0 35305 5 1 1 35304
0 35306 7 1 2 48800 35305
0 35307 5 1 1 35306
0 35308 7 1 2 35297 35307
0 35309 7 1 2 35270 35308
0 35310 5 1 1 35309
0 35311 7 1 2 53555 35310
0 35312 5 1 1 35311
0 35313 7 1 2 70138 71234
0 35314 5 1 1 35313
0 35315 7 1 2 70182 35314
0 35316 5 1 1 35315
0 35317 7 1 2 50507 35316
0 35318 5 1 1 35317
0 35319 7 4 2 50107 76429
0 35320 5 1 1 78260
0 35321 7 2 2 54760 35320
0 35322 5 2 1 78264
0 35323 7 1 2 58048 77223
0 35324 5 1 1 35323
0 35325 7 1 2 78265 35324
0 35326 5 1 1 35325
0 35327 7 1 2 49622 77787
0 35328 5 1 1 35327
0 35329 7 1 2 56645 35328
0 35330 7 1 2 35326 35329
0 35331 5 1 1 35330
0 35332 7 1 2 58049 77682
0 35333 5 1 1 35332
0 35334 7 1 2 71154 73267
0 35335 5 1 1 35334
0 35336 7 1 2 35333 35335
0 35337 5 1 1 35336
0 35338 7 1 2 77129 35337
0 35339 5 1 1 35338
0 35340 7 1 2 49623 71627
0 35341 5 2 1 35340
0 35342 7 1 2 52564 78268
0 35343 5 1 1 35342
0 35344 7 1 2 65299 71064
0 35345 5 2 1 35344
0 35346 7 1 2 35343 78270
0 35347 7 1 2 35339 35346
0 35348 7 1 2 35331 35347
0 35349 5 1 1 35348
0 35350 7 1 2 51111 35349
0 35351 5 1 1 35350
0 35352 7 1 2 35318 35351
0 35353 5 1 1 35352
0 35354 7 1 2 57646 35353
0 35355 5 1 1 35354
0 35356 7 1 2 58050 71031
0 35357 5 1 1 35356
0 35358 7 1 2 60551 61829
0 35359 5 1 1 35358
0 35360 7 1 2 35357 35359
0 35361 5 1 1 35360
0 35362 7 1 2 51112 35361
0 35363 5 1 1 35362
0 35364 7 1 2 56468 60790
0 35365 5 1 1 35364
0 35366 7 1 2 35363 35365
0 35367 5 1 1 35366
0 35368 7 1 2 55937 35367
0 35369 5 1 1 35368
0 35370 7 1 2 52905 75354
0 35371 5 1 1 35370
0 35372 7 1 2 14627 35371
0 35373 5 1 1 35372
0 35374 7 1 2 67724 35373
0 35375 5 1 1 35374
0 35376 7 1 2 35369 35375
0 35377 5 1 1 35376
0 35378 7 1 2 57040 35377
0 35379 5 1 1 35378
0 35380 7 1 2 55938 68202
0 35381 5 2 1 35380
0 35382 7 1 2 74909 78272
0 35383 5 1 1 35382
0 35384 7 1 2 56236 35383
0 35385 5 1 1 35384
0 35386 7 1 2 60796 72682
0 35387 5 1 1 35386
0 35388 7 1 2 55082 35387
0 35389 5 1 1 35388
0 35390 7 1 2 76750 25100
0 35391 5 1 1 35390
0 35392 7 1 2 35389 35391
0 35393 5 1 1 35392
0 35394 7 1 2 35385 35393
0 35395 5 1 1 35394
0 35396 7 1 2 58051 35395
0 35397 5 1 1 35396
0 35398 7 1 2 50264 35211
0 35399 5 1 1 35398
0 35400 7 1 2 66205 67757
0 35401 7 1 2 76027 35400
0 35402 7 1 2 35399 35401
0 35403 7 1 2 78273 35402
0 35404 5 1 1 35403
0 35405 7 1 2 56469 35404
0 35406 5 1 1 35405
0 35407 7 1 2 55939 71043
0 35408 5 1 1 35407
0 35409 7 1 2 71564 35408
0 35410 5 1 1 35409
0 35411 7 1 2 51113 61354
0 35412 7 1 2 35410 35411
0 35413 5 1 1 35412
0 35414 7 1 2 35406 35413
0 35415 7 1 2 35397 35414
0 35416 7 1 2 35379 35415
0 35417 7 1 2 35355 35416
0 35418 5 1 1 35417
0 35419 7 1 2 49780 35418
0 35420 5 1 1 35419
0 35421 7 1 2 35312 35420
0 35422 7 1 2 35262 35421
0 35423 5 1 1 35422
0 35424 7 1 2 49939 35423
0 35425 5 1 1 35424
0 35426 7 1 2 35207 35425
0 35427 5 1 1 35426
0 35428 7 1 2 51380 35427
0 35429 5 1 1 35428
0 35430 7 1 2 62642 77680
0 35431 5 1 1 35430
0 35432 7 1 2 65872 77260
0 35433 7 1 2 71044 35432
0 35434 5 1 1 35433
0 35435 7 1 2 35431 35434
0 35436 5 1 1 35435
0 35437 7 1 2 57041 35436
0 35438 5 1 1 35437
0 35439 7 1 2 50508 70829
0 35440 5 1 1 35439
0 35441 7 1 2 28156 35440
0 35442 5 1 1 35441
0 35443 7 1 2 75783 35442
0 35444 5 1 1 35443
0 35445 7 1 2 35438 35444
0 35446 5 2 1 35445
0 35447 7 1 2 51114 78274
0 35448 5 1 1 35447
0 35449 7 1 2 76796 76836
0 35450 5 1 1 35449
0 35451 7 1 2 35448 35450
0 35452 5 1 1 35451
0 35453 7 1 2 58052 35452
0 35454 5 1 1 35453
0 35455 7 1 2 50265 63525
0 35456 5 1 1 35455
0 35457 7 1 2 60552 77491
0 35458 5 1 1 35457
0 35459 7 1 2 35456 35458
0 35460 5 1 1 35459
0 35461 7 1 2 57647 35460
0 35462 5 1 1 35461
0 35463 7 1 2 71093 78160
0 35464 7 1 2 65304 35463
0 35465 5 1 1 35464
0 35466 7 1 2 35462 35465
0 35467 5 1 1 35466
0 35468 7 1 2 56646 35467
0 35469 5 1 1 35468
0 35470 7 1 2 61593 76099
0 35471 7 1 2 78266 35470
0 35472 5 1 1 35471
0 35473 7 1 2 63547 35472
0 35474 5 1 1 35473
0 35475 7 1 2 77130 78164
0 35476 7 1 2 35474 35475
0 35477 5 1 1 35476
0 35478 7 1 2 66360 73781
0 35479 5 1 1 35478
0 35480 7 2 2 54761 59919
0 35481 5 1 1 78276
0 35482 7 1 2 35479 35481
0 35483 5 1 1 35482
0 35484 7 1 2 77683 35483
0 35485 5 1 1 35484
0 35486 7 1 2 64523 71032
0 35487 5 1 1 35486
0 35488 7 1 2 56404 35487
0 35489 5 1 1 35488
0 35490 7 1 2 55940 2819
0 35491 5 1 1 35490
0 35492 7 1 2 48557 65194
0 35493 7 1 2 35491 35492
0 35494 5 1 1 35493
0 35495 7 1 2 60584 59162
0 35496 7 1 2 35494 35495
0 35497 7 1 2 35489 35496
0 35498 5 1 1 35497
0 35499 7 1 2 35485 35498
0 35500 7 1 2 35477 35499
0 35501 7 1 2 35469 35500
0 35502 5 1 1 35501
0 35503 7 1 2 56470 35502
0 35504 5 1 1 35503
0 35505 7 1 2 35454 35504
0 35506 5 1 1 35505
0 35507 7 1 2 52694 35506
0 35508 5 1 1 35507
0 35509 7 1 2 58766 71235
0 35510 5 1 1 35509
0 35511 7 1 2 58121 35510
0 35512 5 1 1 35511
0 35513 7 1 2 69664 35512
0 35514 5 1 1 35513
0 35515 7 1 2 48801 78271
0 35516 5 1 1 35515
0 35517 7 1 2 3582 77796
0 35518 5 1 1 35517
0 35519 7 1 2 56647 35518
0 35520 5 1 1 35519
0 35521 7 1 2 70159 35520
0 35522 5 1 1 35521
0 35523 7 1 2 35516 35522
0 35524 5 1 1 35523
0 35525 7 1 2 14549 25113
0 35526 5 1 1 35525
0 35527 7 1 2 56648 35526
0 35528 5 1 1 35527
0 35529 7 1 2 76456 35528
0 35530 5 1 1 35529
0 35531 7 1 2 78269 35530
0 35532 5 1 1 35531
0 35533 7 1 2 58073 61693
0 35534 5 1 1 35533
0 35535 7 1 2 61531 70633
0 35536 5 1 1 35535
0 35537 7 1 2 78255 35536
0 35538 5 1 1 35537
0 35539 7 1 2 58767 35538
0 35540 5 1 1 35539
0 35541 7 1 2 35534 35540
0 35542 7 1 2 35532 35541
0 35543 7 1 2 35524 35542
0 35544 5 1 1 35543
0 35545 7 1 2 53130 35544
0 35546 5 1 1 35545
0 35547 7 1 2 35514 35546
0 35548 5 1 1 35547
0 35549 7 1 2 52327 35548
0 35550 5 1 1 35549
0 35551 7 1 2 58053 74088
0 35552 5 1 1 35551
0 35553 7 1 2 50834 71038
0 35554 5 1 1 35553
0 35555 7 1 2 35552 35554
0 35556 5 1 1 35555
0 35557 7 1 2 57042 35556
0 35558 5 1 1 35557
0 35559 7 1 2 58054 65305
0 35560 5 1 1 35559
0 35561 7 1 2 62383 35560
0 35562 5 1 1 35561
0 35563 7 1 2 50509 35562
0 35564 5 1 1 35563
0 35565 7 1 2 56579 35564
0 35566 7 1 2 35558 35565
0 35567 5 1 1 35566
0 35568 7 1 2 52695 35567
0 35569 5 1 1 35568
0 35570 7 1 2 55941 73888
0 35571 7 1 2 78267 35570
0 35572 5 1 1 35571
0 35573 7 1 2 24903 35572
0 35574 5 1 1 35573
0 35575 7 1 2 77131 35574
0 35576 5 1 1 35575
0 35577 7 1 2 71065 75468
0 35578 7 1 2 75746 35577
0 35579 7 1 2 24262 35578
0 35580 5 1 1 35579
0 35581 7 1 2 55083 35580
0 35582 7 1 2 35576 35581
0 35583 7 1 2 35569 35582
0 35584 7 1 2 35550 35583
0 35585 5 1 1 35584
0 35586 7 1 2 58055 78275
0 35587 5 1 1 35586
0 35588 7 1 2 56957 70831
0 35589 5 1 1 35588
0 35590 7 1 2 50510 35589
0 35591 5 1 1 35590
0 35592 7 1 2 66641 77262
0 35593 5 2 1 35592
0 35594 7 1 2 60862 78278
0 35595 5 1 1 35594
0 35596 7 1 2 54762 61321
0 35597 7 1 2 70948 35596
0 35598 7 1 2 35595 35597
0 35599 7 1 2 35591 35598
0 35600 5 1 1 35599
0 35601 7 1 2 48237 63888
0 35602 5 1 1 35601
0 35603 7 2 2 65459 35602
0 35604 7 1 2 57648 75469
0 35605 7 1 2 78280 35604
0 35606 5 1 1 35605
0 35607 7 1 2 52696 35606
0 35608 7 1 2 35600 35607
0 35609 5 1 1 35608
0 35610 7 1 2 67398 75361
0 35611 5 1 1 35610
0 35612 7 1 2 56405 60839
0 35613 5 1 1 35612
0 35614 7 1 2 66654 75442
0 35615 7 1 2 35613 35614
0 35616 5 1 1 35615
0 35617 7 1 2 35611 35616
0 35618 5 1 1 35617
0 35619 7 1 2 52565 35618
0 35620 5 1 1 35619
0 35621 7 1 2 51115 35620
0 35622 7 1 2 35609 35621
0 35623 7 1 2 77804 76233
0 35624 5 1 1 35623
0 35625 7 1 2 75443 77633
0 35626 5 1 1 35625
0 35627 7 1 2 56769 10074
0 35628 5 1 1 35627
0 35629 7 1 2 50266 73435
0 35630 7 1 2 78152 35629
0 35631 7 1 2 35628 35630
0 35632 5 1 1 35631
0 35633 7 1 2 35626 35632
0 35634 5 1 1 35633
0 35635 7 1 2 52566 35634
0 35636 5 1 1 35635
0 35637 7 1 2 35624 35636
0 35638 5 1 1 35637
0 35639 7 1 2 57649 35638
0 35640 5 1 1 35639
0 35641 7 1 2 61830 71247
0 35642 5 1 1 35641
0 35643 7 1 2 50267 67204
0 35644 5 1 1 35643
0 35645 7 1 2 35642 35644
0 35646 5 1 1 35645
0 35647 7 1 2 75362 35646
0 35648 5 1 1 35647
0 35649 7 1 2 60718 66642
0 35650 5 1 1 35649
0 35651 7 1 2 75450 35650
0 35652 5 1 1 35651
0 35653 7 1 2 35648 35652
0 35654 5 1 1 35653
0 35655 7 1 2 50511 35654
0 35656 5 1 1 35655
0 35657 7 1 2 35640 35656
0 35658 7 1 2 35622 35657
0 35659 7 1 2 35587 35658
0 35660 5 1 1 35659
0 35661 7 1 2 53556 35660
0 35662 7 1 2 35585 35661
0 35663 5 1 1 35662
0 35664 7 1 2 35508 35663
0 35665 5 1 1 35664
0 35666 7 1 2 55379 35665
0 35667 5 1 1 35666
0 35668 7 1 2 58056 61438
0 35669 5 1 1 35668
0 35670 7 1 2 76003 35669
0 35671 5 4 1 35670
0 35672 7 1 2 77224 78282
0 35673 5 1 1 35672
0 35674 7 1 2 70342 76004
0 35675 5 2 1 35674
0 35676 7 1 2 59769 77263
0 35677 5 2 1 35676
0 35678 7 1 2 63231 78288
0 35679 7 1 2 78286 35678
0 35680 5 1 1 35679
0 35681 7 1 2 35673 35680
0 35682 5 1 1 35681
0 35683 7 1 2 50512 35682
0 35684 5 1 1 35683
0 35685 7 1 2 67399 78283
0 35686 5 1 1 35685
0 35687 7 1 2 75404 35686
0 35688 7 1 2 35684 35687
0 35689 5 1 1 35688
0 35690 7 1 2 59155 35689
0 35691 5 1 1 35690
0 35692 7 1 2 35667 35691
0 35693 5 1 1 35692
0 35694 7 1 2 49940 35693
0 35695 5 1 1 35694
0 35696 7 1 2 35429 35695
0 35697 5 1 1 35696
0 35698 7 1 2 55547 35697
0 35699 5 1 1 35698
0 35700 7 3 2 60585 63867
0 35701 7 1 2 64724 78290
0 35702 5 1 1 35701
0 35703 7 1 2 66330 71384
0 35704 5 1 1 35703
0 35705 7 1 2 35702 35704
0 35706 5 1 1 35705
0 35707 7 1 2 66966 35706
0 35708 5 1 1 35707
0 35709 7 1 2 74044 72549
0 35710 5 1 1 35709
0 35711 7 1 2 35708 35710
0 35712 5 1 1 35711
0 35713 7 1 2 57185 35712
0 35714 5 1 1 35713
0 35715 7 2 2 66100 67438
0 35716 5 1 1 78293
0 35717 7 1 2 25547 35716
0 35718 5 1 1 35717
0 35719 7 1 2 47979 35718
0 35720 5 1 1 35719
0 35721 7 1 2 66101 66820
0 35722 5 2 1 35721
0 35723 7 1 2 35720 78295
0 35724 5 1 1 35723
0 35725 7 1 2 57960 35724
0 35726 5 1 1 35725
0 35727 7 2 2 62614 68939
0 35728 5 1 1 78297
0 35729 7 1 2 56580 72884
0 35730 7 1 2 78298 35729
0 35731 5 1 1 35730
0 35732 7 1 2 65749 68286
0 35733 5 1 1 35732
0 35734 7 1 2 57961 74450
0 35735 7 1 2 35733 35734
0 35736 5 1 1 35735
0 35737 7 1 2 35731 35736
0 35738 5 1 1 35737
0 35739 7 1 2 56770 35738
0 35740 5 1 1 35739
0 35741 7 1 2 35726 35740
0 35742 7 1 2 35714 35741
0 35743 5 1 1 35742
0 35744 7 1 2 56958 35743
0 35745 5 1 1 35744
0 35746 7 1 2 64771 71673
0 35747 7 1 2 78291 35746
0 35748 5 1 1 35747
0 35749 7 1 2 73621 78123
0 35750 7 1 2 66920 35749
0 35751 5 1 1 35750
0 35752 7 1 2 35748 35751
0 35753 7 1 2 35745 35752
0 35754 5 1 1 35753
0 35755 7 1 2 57522 35754
0 35756 5 1 1 35755
0 35757 7 1 2 62734 73899
0 35758 5 1 1 35757
0 35759 7 1 2 54088 76638
0 35760 5 1 1 35759
0 35761 7 1 2 78296 35760
0 35762 5 1 1 35761
0 35763 7 1 2 61002 35762
0 35764 5 1 1 35763
0 35765 7 1 2 35758 35764
0 35766 5 1 1 35765
0 35767 7 1 2 64291 35766
0 35768 5 1 1 35767
0 35769 7 1 2 51116 66380
0 35770 7 1 2 61813 35769
0 35771 7 1 2 66006 35770
0 35772 5 1 1 35771
0 35773 7 1 2 35768 35772
0 35774 7 1 2 35756 35773
0 35775 5 1 1 35774
0 35776 7 1 2 48802 35775
0 35777 5 1 1 35776
0 35778 7 1 2 67148 71981
0 35779 5 1 1 35778
0 35780 7 1 2 69769 35779
0 35781 5 1 1 35780
0 35782 7 1 2 52697 35781
0 35783 5 1 1 35782
0 35784 7 1 2 67225 75673
0 35785 7 1 2 76016 35784
0 35786 5 1 1 35785
0 35787 7 1 2 35783 35786
0 35788 5 1 1 35787
0 35789 7 1 2 55548 35788
0 35790 5 1 1 35789
0 35791 7 3 2 59064 65989
0 35792 5 1 1 78299
0 35793 7 1 2 67086 78300
0 35794 5 1 1 35793
0 35795 7 1 2 35790 35794
0 35796 5 1 1 35795
0 35797 7 1 2 53557 35796
0 35798 5 1 1 35797
0 35799 7 1 2 64922 71982
0 35800 5 1 1 35799
0 35801 7 1 2 73751 35800
0 35802 5 1 1 35801
0 35803 7 1 2 71910 35802
0 35804 5 1 1 35803
0 35805 7 1 2 57747 72130
0 35806 5 1 1 35805
0 35807 7 1 2 35804 35806
0 35808 5 1 1 35807
0 35809 7 1 2 57523 35808
0 35810 5 1 1 35809
0 35811 7 1 2 57748 70089
0 35812 7 1 2 69671 35811
0 35813 5 1 1 35812
0 35814 7 1 2 63787 66325
0 35815 7 1 2 66619 35814
0 35816 5 1 1 35815
0 35817 7 1 2 35813 35816
0 35818 5 1 1 35817
0 35819 7 1 2 57524 35818
0 35820 5 1 1 35819
0 35821 7 1 2 76538 35820
0 35822 5 1 1 35821
0 35823 7 1 2 56581 35822
0 35824 5 1 1 35823
0 35825 7 1 2 56959 72131
0 35826 5 1 1 35825
0 35827 7 1 2 53387 66844
0 35828 7 1 2 72954 35827
0 35829 5 1 1 35828
0 35830 7 1 2 35826 35829
0 35831 7 1 2 35824 35830
0 35832 7 1 2 35810 35831
0 35833 5 1 1 35832
0 35834 7 1 2 51612 35833
0 35835 5 1 1 35834
0 35836 7 1 2 35798 35835
0 35837 5 1 1 35836
0 35838 7 1 2 54089 35837
0 35839 5 1 1 35838
0 35840 7 1 2 75042 75703
0 35841 5 1 1 35840
0 35842 7 1 2 54388 78301
0 35843 5 1 1 35842
0 35844 7 1 2 35841 35843
0 35845 5 1 1 35844
0 35846 7 1 2 53558 35845
0 35847 5 1 1 35846
0 35848 7 1 2 72885 75686
0 35849 5 1 1 35848
0 35850 7 1 2 35847 35849
0 35851 5 1 1 35850
0 35852 7 1 2 55084 35851
0 35853 5 1 1 35852
0 35854 7 1 2 56582 63848
0 35855 7 1 2 64890 35854
0 35856 5 1 1 35855
0 35857 7 1 2 51381 67707
0 35858 5 1 1 35857
0 35859 7 1 2 7512 35858
0 35860 7 1 2 35856 35859
0 35861 5 1 1 35860
0 35862 7 1 2 62572 35861
0 35863 5 1 1 35862
0 35864 7 1 2 65574 75828
0 35865 5 1 1 35864
0 35866 7 2 2 51382 71716
0 35867 5 1 1 78302
0 35868 7 1 2 63407 78303
0 35869 5 1 1 35868
0 35870 7 1 2 35865 35869
0 35871 7 1 2 35863 35870
0 35872 5 1 1 35871
0 35873 7 1 2 51613 35872
0 35874 5 1 1 35873
0 35875 7 1 2 35853 35874
0 35876 5 1 1 35875
0 35877 7 1 2 54763 35876
0 35878 5 1 1 35877
0 35879 7 1 2 57713 75308
0 35880 5 1 1 35879
0 35881 7 1 2 62973 63319
0 35882 5 3 1 35881
0 35883 7 2 2 51614 78304
0 35884 7 1 2 55085 78307
0 35885 5 1 1 35884
0 35886 7 1 2 35880 35885
0 35887 5 1 1 35886
0 35888 7 1 2 74451 35887
0 35889 5 1 1 35888
0 35890 7 1 2 35878 35889
0 35891 7 1 2 35839 35890
0 35892 5 1 1 35891
0 35893 7 1 2 56771 35892
0 35894 5 1 1 35893
0 35895 7 1 2 68359 75534
0 35896 5 1 1 35895
0 35897 7 1 2 35792 35896
0 35898 5 1 1 35897
0 35899 7 1 2 57749 35898
0 35900 5 1 1 35899
0 35901 7 1 2 53388 62871
0 35902 7 1 2 72509 35901
0 35903 5 1 1 35902
0 35904 7 1 2 35900 35903
0 35905 5 1 1 35904
0 35906 7 1 2 55086 35905
0 35907 5 1 1 35906
0 35908 7 4 2 52698 50835
0 35909 7 1 2 68366 78309
0 35910 5 1 1 35909
0 35911 7 1 2 35907 35910
0 35912 5 1 1 35911
0 35913 7 1 2 53559 35912
0 35914 5 1 1 35913
0 35915 7 1 2 70090 74184
0 35916 5 1 1 35915
0 35917 7 2 2 57525 63526
0 35918 5 1 1 78313
0 35919 7 1 2 69511 78314
0 35920 5 1 1 35919
0 35921 7 1 2 35916 35920
0 35922 5 1 1 35921
0 35923 7 1 2 47980 35922
0 35924 5 1 1 35923
0 35925 7 1 2 63193 63853
0 35926 5 1 1 35925
0 35927 7 1 2 35924 35926
0 35928 5 1 1 35927
0 35929 7 1 2 63312 35928
0 35930 5 1 1 35929
0 35931 7 1 2 64760 78292
0 35932 5 1 1 35931
0 35933 7 1 2 72458 35932
0 35934 5 1 1 35933
0 35935 7 1 2 62573 35934
0 35936 5 1 1 35935
0 35937 7 2 2 55380 73202
0 35938 5 1 1 78315
0 35939 7 1 2 35938 35867
0 35940 5 1 1 35939
0 35941 7 1 2 69126 35940
0 35942 5 1 1 35941
0 35943 7 4 2 54389 63741
0 35944 7 1 2 65663 78317
0 35945 5 1 1 35944
0 35946 7 1 2 35942 35945
0 35947 5 1 1 35946
0 35948 7 1 2 54764 35947
0 35949 5 1 1 35948
0 35950 7 2 2 64270 64336
0 35951 7 1 2 75829 78321
0 35952 5 1 1 35951
0 35953 7 1 2 67002 76603
0 35954 5 1 1 35953
0 35955 7 1 2 35952 35954
0 35956 5 1 1 35955
0 35957 7 1 2 54090 35956
0 35958 5 1 1 35957
0 35959 7 1 2 35949 35958
0 35960 7 1 2 35936 35959
0 35961 7 1 2 35930 35960
0 35962 5 1 1 35961
0 35963 7 1 2 51615 35962
0 35964 5 1 1 35963
0 35965 7 1 2 35914 35964
0 35966 5 1 1 35965
0 35967 7 1 2 57186 35966
0 35968 5 1 1 35967
0 35969 7 2 2 59025 75093
0 35970 7 2 2 51117 78323
0 35971 5 1 1 78325
0 35972 7 1 2 54390 78326
0 35973 5 1 1 35972
0 35974 7 1 2 47981 67335
0 35975 5 1 1 35974
0 35976 7 1 2 69685 35975
0 35977 5 1 1 35976
0 35978 7 1 2 48666 35977
0 35979 5 1 1 35978
0 35980 7 1 2 64173 74292
0 35981 5 2 1 35980
0 35982 7 1 2 35979 78327
0 35983 5 1 1 35982
0 35984 7 1 2 56960 35983
0 35985 5 1 1 35984
0 35986 7 2 2 62574 64578
0 35987 5 1 1 78329
0 35988 7 2 2 72335 35987
0 35989 5 3 1 78331
0 35990 7 1 2 64152 78333
0 35991 5 1 1 35990
0 35992 7 1 2 35985 35991
0 35993 5 1 1 35992
0 35994 7 1 2 51616 64481
0 35995 7 1 2 35993 35994
0 35996 5 1 1 35995
0 35997 7 1 2 35973 35996
0 35998 5 1 1 35997
0 35999 7 1 2 55381 35998
0 36000 5 1 1 35999
0 36001 7 2 2 50836 71763
0 36002 7 2 2 73203 78336
0 36003 5 1 1 78338
0 36004 7 2 2 47982 78339
0 36005 5 1 1 78340
0 36006 7 1 2 64514 66866
0 36007 5 1 1 36006
0 36008 7 1 2 60401 36007
0 36009 5 1 1 36008
0 36010 7 1 2 63472 36009
0 36011 5 1 1 36010
0 36012 7 1 2 49624 71879
0 36013 7 1 2 36011 36012
0 36014 5 1 1 36013
0 36015 7 1 2 36005 36014
0 36016 5 1 1 36015
0 36017 7 1 2 67226 36016
0 36018 5 1 1 36017
0 36019 7 1 2 53389 64932
0 36020 5 1 1 36019
0 36021 7 2 2 47983 62493
0 36022 7 1 2 67617 78342
0 36023 5 2 1 36022
0 36024 7 1 2 71880 78322
0 36025 5 1 1 36024
0 36026 7 1 2 78344 36025
0 36027 5 1 1 36026
0 36028 7 1 2 36020 36027
0 36029 5 1 1 36028
0 36030 7 1 2 71717 74500
0 36031 5 1 1 36030
0 36032 7 1 2 62974 64355
0 36033 5 1 1 36032
0 36034 7 1 2 65507 65856
0 36035 7 1 2 36033 36034
0 36036 5 1 1 36035
0 36037 7 1 2 36031 36036
0 36038 5 1 1 36037
0 36039 7 1 2 51617 36038
0 36040 5 1 1 36039
0 36041 7 1 2 36029 36040
0 36042 7 1 2 36018 36041
0 36043 5 1 1 36042
0 36044 7 1 2 51383 36043
0 36045 5 1 1 36044
0 36046 7 1 2 61393 72385
0 36047 7 1 2 71962 36046
0 36048 5 1 1 36047
0 36049 7 1 2 5377 36048
0 36050 5 1 1 36049
0 36051 7 1 2 57285 36050
0 36052 5 1 1 36051
0 36053 7 4 2 55549 59357
0 36054 7 1 2 63195 77047
0 36055 5 1 1 36054
0 36056 7 1 2 78346 36055
0 36057 5 1 1 36056
0 36058 7 2 2 64812 71881
0 36059 5 2 1 78350
0 36060 7 1 2 61003 78351
0 36061 5 1 1 36060
0 36062 7 1 2 36057 36061
0 36063 5 1 1 36062
0 36064 7 1 2 54765 36063
0 36065 5 1 1 36064
0 36066 7 1 2 36052 36065
0 36067 5 1 1 36066
0 36068 7 1 2 51384 36067
0 36069 5 1 1 36068
0 36070 7 1 2 5237 73950
0 36071 5 1 1 36070
0 36072 7 5 2 55382 71882
0 36073 7 1 2 51118 78354
0 36074 7 1 2 36071 36073
0 36075 5 1 1 36074
0 36076 7 1 2 36069 36075
0 36077 5 1 1 36076
0 36078 7 1 2 57105 36077
0 36079 5 1 1 36078
0 36080 7 1 2 36045 36079
0 36081 7 1 2 36000 36080
0 36082 7 1 2 35968 36081
0 36083 7 1 2 35894 36082
0 36084 5 1 1 36083
0 36085 7 1 2 49941 36084
0 36086 5 1 1 36085
0 36087 7 1 2 35777 36086
0 36088 5 1 1 36087
0 36089 7 1 2 55806 36088
0 36090 5 1 1 36089
0 36091 7 1 2 62931 67583
0 36092 5 1 1 36091
0 36093 7 2 2 62575 67584
0 36094 5 1 1 78359
0 36095 7 1 2 65410 64198
0 36096 5 1 1 36095
0 36097 7 1 2 36094 36096
0 36098 5 1 1 36097
0 36099 7 1 2 65575 36098
0 36100 5 1 1 36099
0 36101 7 1 2 36092 36100
0 36102 5 1 1 36101
0 36103 7 1 2 51618 36102
0 36104 5 1 1 36103
0 36105 7 1 2 53390 72489
0 36106 5 1 1 36105
0 36107 7 1 2 22913 36106
0 36108 5 1 1 36107
0 36109 7 1 2 71722 36108
0 36110 5 1 1 36109
0 36111 7 1 2 36104 36110
0 36112 5 1 1 36111
0 36113 7 1 2 54766 36112
0 36114 5 1 1 36113
0 36115 7 1 2 65673 78341
0 36116 5 1 1 36115
0 36117 7 1 2 36114 36116
0 36118 5 1 1 36117
0 36119 7 1 2 57526 36118
0 36120 5 1 1 36119
0 36121 7 1 2 51619 64694
0 36122 7 1 2 78360 36121
0 36123 5 1 1 36122
0 36124 7 1 2 71113 71764
0 36125 7 1 2 65674 36124
0 36126 5 1 1 36125
0 36127 7 1 2 36123 36126
0 36128 5 1 1 36127
0 36129 7 1 2 54767 36128
0 36130 5 1 1 36129
0 36131 7 1 2 36003 36130
0 36132 5 1 1 36131
0 36133 7 1 2 67227 36132
0 36134 5 1 1 36133
0 36135 7 1 2 75094 72322
0 36136 7 1 2 65692 36135
0 36137 5 1 1 36136
0 36138 7 1 2 36134 36137
0 36139 7 1 2 36120 36138
0 36140 5 1 1 36139
0 36141 7 1 2 51385 36140
0 36142 5 1 1 36141
0 36143 7 2 2 68334 78343
0 36144 5 1 1 78361
0 36145 7 1 2 65497 70091
0 36146 5 1 1 36145
0 36147 7 1 2 61719 73750
0 36148 5 1 1 36147
0 36149 7 1 2 16780 36148
0 36150 5 1 1 36149
0 36151 7 1 2 63313 36150
0 36152 5 1 1 36151
0 36153 7 1 2 54391 76535
0 36154 5 1 1 36153
0 36155 7 1 2 60553 74742
0 36156 5 1 1 36155
0 36157 7 1 2 36154 36156
0 36158 7 1 2 36152 36157
0 36159 5 1 1 36158
0 36160 7 1 2 55087 36159
0 36161 5 1 1 36160
0 36162 7 1 2 36146 36161
0 36163 5 1 1 36162
0 36164 7 1 2 51620 36163
0 36165 5 1 1 36164
0 36166 7 1 2 36144 36165
0 36167 5 1 1 36166
0 36168 7 1 2 60308 36167
0 36169 5 1 1 36168
0 36170 7 1 2 72390 71965
0 36171 5 1 1 36170
0 36172 7 1 2 68646 36171
0 36173 5 1 1 36172
0 36174 7 1 2 60309 36173
0 36175 5 1 1 36174
0 36176 7 1 2 50268 78347
0 36177 5 1 1 36176
0 36178 7 1 2 78352 36177
0 36179 5 1 1 36178
0 36180 7 1 2 60000 58277
0 36181 7 1 2 36179 36180
0 36182 5 1 1 36181
0 36183 7 1 2 36175 36182
0 36184 5 1 1 36183
0 36185 7 1 2 51386 36184
0 36186 5 1 1 36185
0 36187 7 1 2 65708 71745
0 36188 7 1 2 58634 36187
0 36189 5 1 1 36188
0 36190 7 1 2 36186 36189
0 36191 5 1 1 36190
0 36192 7 1 2 57106 36191
0 36193 5 1 1 36192
0 36194 7 1 2 67347 66707
0 36195 5 1 1 36194
0 36196 7 5 2 64579 59289
0 36197 7 1 2 55088 67585
0 36198 7 1 2 78363 36197
0 36199 5 1 1 36198
0 36200 7 1 2 36195 36199
0 36201 5 1 1 36200
0 36202 7 1 2 54768 36201
0 36203 5 1 1 36202
0 36204 7 1 2 67602 72349
0 36205 5 1 1 36204
0 36206 7 1 2 36203 36205
0 36207 5 1 1 36206
0 36208 7 1 2 65990 36207
0 36209 5 1 1 36208
0 36210 7 1 2 36193 36209
0 36211 7 1 2 36169 36210
0 36212 7 1 2 36142 36211
0 36213 5 1 1 36212
0 36214 7 1 2 49942 36213
0 36215 5 1 1 36214
0 36216 7 1 2 67336 69512
0 36217 5 1 1 36216
0 36218 7 1 2 49625 71983
0 36219 5 1 1 36218
0 36220 7 1 2 73752 36219
0 36221 5 1 1 36220
0 36222 7 1 2 64813 36221
0 36223 5 1 1 36222
0 36224 7 1 2 36217 36223
0 36225 5 1 1 36224
0 36226 7 1 2 48238 36225
0 36227 5 1 1 36226
0 36228 7 2 2 63788 68875
0 36229 7 1 2 65896 78368
0 36230 5 1 1 36229
0 36231 7 1 2 36227 36230
0 36232 5 1 1 36231
0 36233 7 1 2 47984 36232
0 36234 5 1 1 36233
0 36235 7 1 2 51387 65511
0 36236 5 1 1 36235
0 36237 7 1 2 63849 71856
0 36238 7 1 2 36236 36237
0 36239 5 1 1 36238
0 36240 7 1 2 36234 36239
0 36241 5 1 1 36240
0 36242 7 1 2 64352 36241
0 36243 5 1 1 36242
0 36244 7 1 2 61720 67506
0 36245 7 1 2 67228 78369
0 36246 7 1 2 36244 36245
0 36247 5 1 1 36246
0 36248 7 1 2 36243 36247
0 36249 5 1 1 36248
0 36250 7 1 2 66967 36249
0 36251 5 1 1 36250
0 36252 7 1 2 65664 78294
0 36253 5 1 1 36252
0 36254 7 1 2 36251 36253
0 36255 5 1 1 36254
0 36256 7 1 2 48803 36255
0 36257 5 1 1 36256
0 36258 7 1 2 57107 69238
0 36259 5 1 1 36258
0 36260 7 1 2 56961 69247
0 36261 5 1 1 36260
0 36262 7 1 2 36259 36261
0 36263 5 1 1 36262
0 36264 7 1 2 71746 36263
0 36265 5 1 1 36264
0 36266 7 1 2 64616 66102
0 36267 7 1 2 67068 36266
0 36268 7 1 2 66193 36267
0 36269 5 1 1 36268
0 36270 7 1 2 36265 36269
0 36271 5 1 1 36270
0 36272 7 1 2 74615 36271
0 36273 5 1 1 36272
0 36274 7 1 2 36257 36273
0 36275 7 1 2 36215 36274
0 36276 5 1 1 36275
0 36277 7 1 2 58625 36276
0 36278 5 1 1 36277
0 36279 7 2 2 62494 64356
0 36280 5 3 1 78370
0 36281 7 1 2 53006 60871
0 36282 5 1 1 36281
0 36283 7 1 2 78240 36282
0 36284 5 1 1 36283
0 36285 7 1 2 55942 36284
0 36286 5 1 1 36285
0 36287 7 1 2 69668 36286
0 36288 5 1 1 36287
0 36289 7 1 2 65900 36288
0 36290 5 1 1 36289
0 36291 7 1 2 62932 76745
0 36292 7 1 2 36290 36291
0 36293 5 1 1 36292
0 36294 7 1 2 49626 36293
0 36295 5 1 1 36294
0 36296 7 2 2 54769 67367
0 36297 7 1 2 60310 78375
0 36298 5 1 1 36297
0 36299 7 1 2 54392 73459
0 36300 5 1 1 36299
0 36301 7 1 2 50837 36300
0 36302 5 2 1 36301
0 36303 7 1 2 57527 78377
0 36304 5 1 1 36303
0 36305 7 1 2 65690 36304
0 36306 7 1 2 36298 36305
0 36307 5 2 1 36306
0 36308 7 1 2 53391 78379
0 36309 5 1 1 36308
0 36310 7 1 2 77455 36309
0 36311 7 1 2 36295 36310
0 36312 5 1 1 36311
0 36313 7 1 2 78372 36312
0 36314 5 1 1 36313
0 36315 7 1 2 61869 66140
0 36316 5 1 1 36315
0 36317 7 2 2 60554 36316
0 36318 7 1 2 57528 78381
0 36319 5 1 1 36318
0 36320 7 1 2 53560 78380
0 36321 5 1 1 36320
0 36322 7 1 2 36319 36321
0 36323 5 1 1 36322
0 36324 7 1 2 67242 78371
0 36325 5 1 1 36324
0 36326 7 1 2 36323 36325
0 36327 5 1 1 36326
0 36328 7 1 2 67229 78330
0 36329 5 2 1 36328
0 36330 7 1 2 55383 78383
0 36331 7 1 2 36327 36330
0 36332 7 1 2 36314 36331
0 36333 5 1 1 36332
0 36334 7 1 2 73584 78305
0 36335 5 1 1 36334
0 36336 7 1 2 58289 65843
0 36337 7 1 2 61237 36336
0 36338 5 1 1 36337
0 36339 7 1 2 36335 36338
0 36340 5 1 1 36339
0 36341 7 1 2 54770 36340
0 36342 5 1 1 36341
0 36343 7 1 2 59403 78306
0 36344 5 1 1 36343
0 36345 7 1 2 73725 36344
0 36346 7 1 2 36342 36345
0 36347 5 1 1 36346
0 36348 7 1 2 55089 36347
0 36349 7 1 2 36333 36348
0 36350 5 1 1 36349
0 36351 7 1 2 57529 78376
0 36352 5 1 1 36351
0 36353 7 1 2 2369 36352
0 36354 5 1 1 36353
0 36355 7 1 2 60311 36354
0 36356 5 1 1 36355
0 36357 7 1 2 57650 74180
0 36358 7 1 2 74538 36357
0 36359 5 1 1 36358
0 36360 7 1 2 57108 36359
0 36361 5 1 1 36360
0 36362 7 1 2 64950 58278
0 36363 5 1 1 36362
0 36364 7 1 2 58057 36363
0 36365 7 1 2 36361 36364
0 36366 7 1 2 36356 36365
0 36367 5 1 1 36366
0 36368 7 1 2 62933 36367
0 36369 5 1 1 36368
0 36370 7 1 2 60426 64466
0 36371 7 1 2 78281 36370
0 36372 5 1 1 36371
0 36373 7 1 2 64292 36372
0 36374 5 1 1 36373
0 36375 7 1 2 65682 67365
0 36376 5 2 1 36375
0 36377 7 1 2 64409 67497
0 36378 7 1 2 78385 36377
0 36379 5 1 1 36378
0 36380 7 1 2 36374 36379
0 36381 5 1 1 36380
0 36382 7 1 2 62576 36381
0 36383 5 1 1 36382
0 36384 7 1 2 51388 36383
0 36385 7 1 2 36369 36384
0 36386 5 1 1 36385
0 36387 7 1 2 58217 66165
0 36388 5 1 1 36387
0 36389 7 1 2 47985 36388
0 36390 5 1 1 36389
0 36391 7 1 2 50513 61961
0 36392 5 1 1 36391
0 36393 7 1 2 54771 36392
0 36394 5 1 1 36393
0 36395 7 1 2 65395 36394
0 36396 7 1 2 36390 36395
0 36397 5 1 1 36396
0 36398 7 1 2 61238 36397
0 36399 5 1 1 36398
0 36400 7 1 2 58979 65923
0 36401 5 1 1 36400
0 36402 7 1 2 62495 65928
0 36403 5 1 1 36402
0 36404 7 1 2 59055 63006
0 36405 5 1 1 36404
0 36406 7 1 2 36403 36405
0 36407 5 2 1 36406
0 36408 7 1 2 36401 78387
0 36409 7 1 2 36399 36408
0 36410 5 1 1 36409
0 36411 7 1 2 51119 36410
0 36412 5 1 1 36411
0 36413 7 2 2 48804 75491
0 36414 5 3 1 78389
0 36415 7 1 2 55384 78391
0 36416 7 1 2 36412 36415
0 36417 5 1 1 36416
0 36418 7 1 2 36386 36417
0 36419 5 1 1 36418
0 36420 7 1 2 36350 36419
0 36421 5 1 1 36420
0 36422 7 1 2 49943 36421
0 36423 5 1 1 36422
0 36424 7 2 2 60402 63527
0 36425 7 1 2 59722 78394
0 36426 5 1 1 36425
0 36427 7 1 2 55090 78382
0 36428 5 1 1 36427
0 36429 7 1 2 36426 36428
0 36430 5 1 1 36429
0 36431 7 1 2 67244 36430
0 36432 5 1 1 36431
0 36433 7 1 2 64482 67337
0 36434 5 1 1 36433
0 36435 7 1 2 65897 76318
0 36436 5 1 1 36435
0 36437 7 1 2 51120 64239
0 36438 5 1 1 36437
0 36439 7 1 2 36436 36438
0 36440 5 1 1 36439
0 36441 7 1 2 61057 36440
0 36442 5 1 1 36441
0 36443 7 1 2 36434 36442
0 36444 5 1 1 36443
0 36445 7 1 2 48239 36444
0 36446 5 1 1 36445
0 36447 7 1 2 64814 60555
0 36448 5 2 1 36447
0 36449 7 1 2 28051 78396
0 36450 5 1 1 36449
0 36451 7 1 2 47986 36450
0 36452 5 1 1 36451
0 36453 7 1 2 64541 78395
0 36454 5 1 1 36453
0 36455 7 1 2 36452 36454
0 36456 5 1 1 36455
0 36457 7 1 2 61095 36456
0 36458 5 1 1 36457
0 36459 7 1 2 64960 67338
0 36460 5 1 1 36459
0 36461 7 1 2 36458 36460
0 36462 7 1 2 36446 36461
0 36463 5 1 1 36462
0 36464 7 1 2 55385 36463
0 36465 5 1 1 36464
0 36466 7 1 2 63368 71385
0 36467 7 1 2 77824 36466
0 36468 7 1 2 65840 36467
0 36469 5 1 1 36468
0 36470 7 1 2 36465 36469
0 36471 5 1 1 36470
0 36472 7 1 2 64353 36471
0 36473 5 1 1 36472
0 36474 7 1 2 36432 36473
0 36475 5 1 1 36474
0 36476 7 1 2 62934 36475
0 36477 5 1 1 36476
0 36478 7 1 2 36423 36477
0 36479 5 1 1 36478
0 36480 7 1 2 51621 36479
0 36481 5 1 1 36480
0 36482 7 1 2 57651 60963
0 36483 5 1 1 36482
0 36484 7 1 2 63660 68445
0 36485 5 3 1 36484
0 36486 7 1 2 64126 67698
0 36487 5 1 1 36486
0 36488 7 1 2 78398 36487
0 36489 5 2 1 36488
0 36490 7 1 2 57109 78401
0 36491 5 1 1 36490
0 36492 7 1 2 64293 72547
0 36493 5 1 1 36492
0 36494 7 1 2 36491 36493
0 36495 5 1 1 36494
0 36496 7 1 2 51121 36495
0 36497 5 1 1 36496
0 36498 7 1 2 63742 78308
0 36499 5 1 1 36498
0 36500 7 1 2 36497 36499
0 36501 5 1 1 36500
0 36502 7 1 2 49944 36501
0 36503 5 1 1 36502
0 36504 7 1 2 66586 74263
0 36505 5 1 1 36504
0 36506 7 1 2 21713 36505
0 36507 5 1 1 36506
0 36508 7 1 2 71668 36507
0 36509 5 1 1 36508
0 36510 7 1 2 36503 36509
0 36511 5 1 1 36510
0 36512 7 1 2 36483 36511
0 36513 5 1 1 36512
0 36514 7 1 2 74532 71963
0 36515 5 1 1 36514
0 36516 7 1 2 68647 36515
0 36517 5 1 1 36516
0 36518 7 1 2 57110 36517
0 36519 5 1 1 36518
0 36520 7 1 2 63314 73987
0 36521 5 1 1 36520
0 36522 7 1 2 65499 36521
0 36523 5 1 1 36522
0 36524 7 1 2 62577 36523
0 36525 5 1 1 36524
0 36526 7 1 2 62935 73988
0 36527 5 1 1 36526
0 36528 7 1 2 36525 36527
0 36529 5 1 1 36528
0 36530 7 1 2 51622 36529
0 36531 5 1 1 36530
0 36532 7 1 2 36519 36531
0 36533 5 1 1 36532
0 36534 7 1 2 49945 36533
0 36535 5 1 1 36534
0 36536 7 1 2 64271 67071
0 36537 7 1 2 72539 77899
0 36538 7 1 2 36536 36537
0 36539 5 1 1 36538
0 36540 7 1 2 36535 36539
0 36541 5 1 1 36540
0 36542 7 1 2 51389 36541
0 36543 5 1 1 36542
0 36544 7 1 2 49946 78362
0 36545 5 1 1 36544
0 36546 7 1 2 36543 36545
0 36547 5 1 1 36546
0 36548 7 1 2 59491 36547
0 36549 5 1 1 36548
0 36550 7 1 2 36513 36549
0 36551 7 1 2 36481 36550
0 36552 7 1 2 36278 36551
0 36553 7 1 2 36090 36552
0 36554 7 1 2 35699 36553
0 36555 7 1 2 66122 74277
0 36556 5 1 1 36555
0 36557 7 1 2 24272 36556
0 36558 5 1 1 36557
0 36559 7 1 2 49243 36558
0 36560 5 1 1 36559
0 36561 7 1 2 54091 67348
0 36562 5 1 1 36561
0 36563 7 1 2 36560 36562
0 36564 5 1 1 36563
0 36565 7 1 2 49135 36564
0 36566 5 1 1 36565
0 36567 7 1 2 67349 78106
0 36568 5 1 1 36567
0 36569 7 1 2 36566 36568
0 36570 5 1 1 36569
0 36571 7 1 2 47987 36570
0 36572 5 1 1 36571
0 36573 7 1 2 54393 70794
0 36574 5 1 1 36573
0 36575 7 1 2 74012 36574
0 36576 5 1 1 36575
0 36577 7 1 2 67350 36576
0 36578 5 1 1 36577
0 36579 7 1 2 36572 36578
0 36580 5 1 1 36579
0 36581 7 1 2 48240 36580
0 36582 5 1 1 36581
0 36583 7 1 2 59509 61774
0 36584 5 2 1 36583
0 36585 7 1 2 49136 78403
0 36586 5 1 1 36585
0 36587 7 1 2 73978 36586
0 36588 5 1 1 36587
0 36589 7 1 2 47988 36588
0 36590 5 1 1 36589
0 36591 7 1 2 60728 71409
0 36592 5 1 1 36591
0 36593 7 1 2 49244 36592
0 36594 5 1 1 36593
0 36595 7 1 2 50838 71033
0 36596 7 1 2 36594 36595
0 36597 7 1 2 36590 36596
0 36598 5 1 1 36597
0 36599 7 1 2 76183 36598
0 36600 5 1 1 36599
0 36601 7 1 2 36582 36600
0 36602 5 1 1 36601
0 36603 7 1 2 49499 36602
0 36604 5 1 1 36603
0 36605 7 1 2 62164 70864
0 36606 5 2 1 36605
0 36607 7 1 2 77182 78405
0 36608 5 2 1 36607
0 36609 7 1 2 63528 78407
0 36610 5 1 1 36609
0 36611 7 1 2 69425 72782
0 36612 5 2 1 36611
0 36613 7 1 2 36610 78409
0 36614 5 1 1 36613
0 36615 7 1 2 57962 36614
0 36616 5 1 1 36615
0 36617 7 1 2 36604 36616
0 36618 5 1 1 36617
0 36619 7 1 2 48558 36618
0 36620 5 1 1 36619
0 36621 7 1 2 55807 70865
0 36622 5 1 1 36621
0 36623 7 1 2 59733 36622
0 36624 5 1 1 36623
0 36625 7 1 2 47989 36624
0 36626 5 1 1 36625
0 36627 7 1 2 54394 65562
0 36628 5 1 1 36627
0 36629 7 1 2 61876 36628
0 36630 5 1 1 36629
0 36631 7 1 2 48241 36630
0 36632 5 1 1 36631
0 36633 7 1 2 75743 36632
0 36634 7 1 2 36626 36633
0 36635 5 1 1 36634
0 36636 7 1 2 63529 36635
0 36637 5 1 1 36636
0 36638 7 1 2 78410 36637
0 36639 5 1 1 36638
0 36640 7 1 2 49500 36639
0 36641 5 1 1 36640
0 36642 7 1 2 74776 69426
0 36643 5 1 1 36642
0 36644 7 1 2 36641 36643
0 36645 5 1 1 36644
0 36646 7 1 2 57963 36645
0 36647 5 1 1 36646
0 36648 7 1 2 36620 36647
0 36649 5 1 1 36648
0 36650 7 1 2 71674 36649
0 36651 5 1 1 36650
0 36652 7 1 2 64210 74009
0 36653 5 1 1 36652
0 36654 7 1 2 47990 36653
0 36655 5 1 1 36654
0 36656 7 1 2 57783 36655
0 36657 5 1 1 36656
0 36658 7 1 2 54772 36657
0 36659 5 1 1 36658
0 36660 7 1 2 57759 65918
0 36661 5 1 1 36660
0 36662 7 1 2 58409 36661
0 36663 5 1 1 36662
0 36664 7 1 2 54773 20610
0 36665 5 1 1 36664
0 36666 7 1 2 36663 36665
0 36667 5 1 1 36666
0 36668 7 1 2 48242 36667
0 36669 5 1 1 36668
0 36670 7 1 2 54395 64494
0 36671 5 1 1 36670
0 36672 7 1 2 74851 36671
0 36673 5 1 1 36672
0 36674 7 1 2 55808 36673
0 36675 5 1 1 36674
0 36676 7 1 2 36669 36675
0 36677 7 1 2 36659 36676
0 36678 5 1 1 36677
0 36679 7 1 2 65733 72455
0 36680 7 1 2 36678 36679
0 36681 5 1 1 36680
0 36682 7 1 2 36651 36681
0 36683 5 1 1 36682
0 36684 7 1 2 48805 36683
0 36685 5 1 1 36684
0 36686 7 1 2 57845 74396
0 36687 5 1 1 36686
0 36688 7 1 2 61577 36687
0 36689 5 2 1 36688
0 36690 7 1 2 68122 78404
0 36691 5 1 1 36690
0 36692 7 1 2 55809 62815
0 36693 5 1 1 36692
0 36694 7 1 2 36691 36693
0 36695 7 1 2 78215 36694
0 36696 7 2 2 78411 36695
0 36697 5 1 1 78413
0 36698 7 1 2 36697 78138
0 36699 5 1 1 36698
0 36700 7 1 2 59723 74312
0 36701 5 1 1 36700
0 36702 7 1 2 36699 36701
0 36703 5 1 1 36702
0 36704 7 1 2 55091 36703
0 36705 5 1 1 36704
0 36706 7 1 2 63473 67230
0 36707 7 1 2 64114 36706
0 36708 5 1 1 36707
0 36709 7 1 2 36705 36708
0 36710 5 1 1 36709
0 36711 7 1 2 53392 36710
0 36712 5 1 1 36711
0 36713 7 1 2 49627 64115
0 36714 5 1 1 36713
0 36715 7 1 2 63040 78406
0 36716 5 1 1 36715
0 36717 7 1 2 63461 36716
0 36718 5 1 1 36717
0 36719 7 1 2 36714 36718
0 36720 5 1 1 36719
0 36721 7 1 2 52699 36720
0 36722 5 1 1 36721
0 36723 7 1 2 36712 36722
0 36724 5 1 1 36723
0 36725 7 1 2 71765 36724
0 36726 5 1 1 36725
0 36727 7 1 2 65257 7137
0 36728 5 1 1 36727
0 36729 7 1 2 56406 36728
0 36730 5 1 1 36729
0 36731 7 1 2 48243 78190
0 36732 5 2 1 36731
0 36733 7 1 2 55092 61674
0 36734 5 1 1 36733
0 36735 7 1 2 78415 36734
0 36736 7 1 2 36730 36735
0 36737 5 1 1 36736
0 36738 7 1 2 58880 36737
0 36739 5 2 1 36738
0 36740 7 1 2 55093 73607
0 36741 5 2 1 36740
0 36742 7 1 2 65315 77024
0 36743 5 1 1 36742
0 36744 7 1 2 78419 36743
0 36745 7 1 2 60936 74847
0 36746 5 1 1 36745
0 36747 7 1 2 31266 36746
0 36748 5 1 1 36747
0 36749 7 1 2 56407 36748
0 36750 5 1 1 36749
0 36751 7 1 2 57835 78085
0 36752 5 1 1 36751
0 36753 7 1 2 51122 36752
0 36754 5 1 1 36753
0 36755 7 1 2 56772 36754
0 36756 5 1 1 36755
0 36757 7 1 2 48244 66212
0 36758 5 1 1 36757
0 36759 7 1 2 70037 36758
0 36760 7 1 2 36756 36759
0 36761 5 1 1 36760
0 36762 7 1 2 60705 36761
0 36763 5 1 1 36762
0 36764 7 1 2 36750 36763
0 36765 7 1 2 36744 36764
0 36766 7 1 2 78417 36765
0 36767 5 1 1 36766
0 36768 7 1 2 62936 36767
0 36769 5 1 1 36768
0 36770 7 1 2 68016 74701
0 36771 5 1 1 36770
0 36772 7 1 2 78095 36771
0 36773 5 1 1 36772
0 36774 7 1 2 60706 36773
0 36775 5 1 1 36774
0 36776 7 1 2 59550 59513
0 36777 5 2 1 36776
0 36778 7 1 2 56237 78421
0 36779 5 1 1 36778
0 36780 7 1 2 61578 36779
0 36781 5 1 1 36780
0 36782 7 1 2 68020 68112
0 36783 5 1 1 36782
0 36784 7 1 2 49245 66339
0 36785 5 1 1 36784
0 36786 7 1 2 56238 36785
0 36787 5 1 1 36786
0 36788 7 1 2 36783 36787
0 36789 5 1 1 36788
0 36790 7 1 2 36781 36789
0 36791 5 1 1 36790
0 36792 7 1 2 54774 36791
0 36793 5 1 1 36792
0 36794 7 1 2 60126 74928
0 36795 5 1 1 36794
0 36796 7 1 2 56962 36795
0 36797 5 1 1 36796
0 36798 7 1 2 48245 63269
0 36799 7 1 2 59455 36798
0 36800 5 1 1 36799
0 36801 7 1 2 78420 36800
0 36802 7 1 2 36797 36801
0 36803 7 1 2 36793 36802
0 36804 7 1 2 36775 36803
0 36805 7 1 2 78418 36804
0 36806 5 1 1 36805
0 36807 7 1 2 63000 36806
0 36808 5 1 1 36807
0 36809 7 1 2 36769 36808
0 36810 5 1 1 36809
0 36811 7 1 2 51623 36810
0 36812 5 1 1 36811
0 36813 7 1 2 64669 78416
0 36814 5 1 1 36813
0 36815 7 1 2 60656 36814
0 36816 5 1 1 36815
0 36817 7 1 2 64997 63032
0 36818 5 1 1 36817
0 36819 7 1 2 60556 77167
0 36820 5 1 1 36819
0 36821 7 1 2 55094 36820
0 36822 5 1 1 36821
0 36823 7 1 2 36818 36822
0 36824 7 1 2 36816 36823
0 36825 5 1 1 36824
0 36826 7 1 2 74774 36825
0 36827 5 1 1 36826
0 36828 7 2 2 55095 71883
0 36829 7 1 2 65258 65919
0 36830 5 1 1 36829
0 36831 7 1 2 60937 36830
0 36832 5 1 1 36831
0 36833 7 1 2 78176 36832
0 36834 5 1 1 36833
0 36835 7 1 2 48246 36834
0 36836 5 1 1 36835
0 36837 7 1 2 61683 68145
0 36838 7 1 2 73966 36837
0 36839 5 1 1 36838
0 36840 7 1 2 57784 36839
0 36841 5 1 1 36840
0 36842 7 1 2 54775 36841
0 36843 5 1 1 36842
0 36844 7 1 2 36836 36843
0 36845 7 1 2 74853 36844
0 36846 5 1 1 36845
0 36847 7 1 2 78423 36846
0 36848 5 1 1 36847
0 36849 7 1 2 68099 75309
0 36850 5 1 1 36849
0 36851 7 1 2 57290 78424
0 36852 5 1 1 36851
0 36853 7 1 2 36850 36852
0 36854 5 1 1 36853
0 36855 7 1 2 60707 36854
0 36856 5 1 1 36855
0 36857 7 1 2 58881 68040
0 36858 7 1 2 75310 36857
0 36859 5 1 1 36858
0 36860 7 1 2 67747 71766
0 36861 7 1 2 73608 36860
0 36862 5 1 1 36861
0 36863 7 1 2 36859 36862
0 36864 7 1 2 36856 36863
0 36865 7 1 2 36848 36864
0 36866 5 1 1 36865
0 36867 7 1 2 56408 36866
0 36868 5 1 1 36867
0 36869 7 1 2 36827 36868
0 36870 5 1 1 36869
0 36871 7 1 2 56583 36870
0 36872 5 1 1 36871
0 36873 7 1 2 36812 36872
0 36874 7 1 2 36726 36873
0 36875 5 1 1 36874
0 36876 7 1 2 51390 36875
0 36877 5 1 1 36876
0 36878 7 1 2 59570 78355
0 36879 5 1 1 36878
0 36880 7 2 2 63661 74264
0 36881 7 1 2 48247 78425
0 36882 5 1 1 36881
0 36883 7 1 2 36879 36882
0 36884 5 1 1 36883
0 36885 7 1 2 61579 36884
0 36886 5 1 1 36885
0 36887 7 4 2 55550 67812
0 36888 7 3 2 50839 59558
0 36889 5 1 1 78431
0 36890 7 1 2 61761 62879
0 36891 7 1 2 36889 36890
0 36892 5 1 1 36891
0 36893 7 1 2 74967 36892
0 36894 5 1 1 36893
0 36895 7 1 2 78427 36894
0 36896 5 1 1 36895
0 36897 7 1 2 71906 78356
0 36898 5 1 1 36897
0 36899 7 1 2 36896 36898
0 36900 7 1 2 36886 36899
0 36901 5 1 1 36900
0 36902 7 1 2 55810 36901
0 36903 5 1 1 36902
0 36904 7 1 2 74585 78426
0 36905 5 1 1 36904
0 36906 7 1 2 61980 78402
0 36907 5 1 1 36906
0 36908 7 1 2 36905 36907
0 36909 5 1 1 36908
0 36910 7 1 2 47991 36909
0 36911 5 1 1 36910
0 36912 7 1 2 61881 78357
0 36913 5 1 1 36912
0 36914 7 1 2 65385 77869
0 36915 5 1 1 36914
0 36916 7 1 2 78358 36915
0 36917 5 1 1 36916
0 36918 7 1 2 61762 78428
0 36919 7 1 2 78227 36918
0 36920 5 1 1 36919
0 36921 7 1 2 36917 36920
0 36922 5 1 1 36921
0 36923 7 1 2 48248 36922
0 36924 5 1 1 36923
0 36925 7 1 2 36913 36924
0 36926 7 1 2 36911 36925
0 36927 7 1 2 36903 36926
0 36928 5 1 1 36927
0 36929 7 1 2 51123 36928
0 36930 5 1 1 36929
0 36931 7 2 2 60403 68398
0 36932 5 1 1 78434
0 36933 7 1 2 68603 36932
0 36934 5 1 1 36933
0 36935 7 1 2 48806 36934
0 36936 5 1 1 36935
0 36937 7 2 2 54092 68296
0 36938 7 1 2 67681 78436
0 36939 5 1 1 36938
0 36940 7 1 2 36936 36939
0 36941 5 1 1 36940
0 36942 7 1 2 51624 36941
0 36943 5 1 1 36942
0 36944 7 2 2 74977 78348
0 36945 5 1 1 78438
0 36946 7 1 2 36943 36945
0 36947 5 1 1 36946
0 36948 7 1 2 797 36947
0 36949 5 1 1 36948
0 36950 7 1 2 51391 60820
0 36951 7 1 2 66987 36950
0 36952 5 1 1 36951
0 36953 7 1 2 36949 36952
0 36954 7 1 2 36930 36953
0 36955 5 1 1 36954
0 36956 7 1 2 57111 36955
0 36957 5 1 1 36956
0 36958 7 1 2 78211 78324
0 36959 5 1 1 36958
0 36960 7 1 2 50840 78414
0 36961 5 1 1 36960
0 36962 7 1 2 64294 36961
0 36963 5 1 1 36962
0 36964 7 1 2 56409 61228
0 36965 5 2 1 36964
0 36966 7 2 2 54776 58980
0 36967 7 3 2 56410 78442
0 36968 7 1 2 78408 78444
0 36969 5 1 1 36968
0 36970 7 1 2 78440 36969
0 36971 7 1 2 36963 36970
0 36972 5 1 1 36971
0 36973 7 1 2 51625 36972
0 36974 5 1 1 36973
0 36975 7 1 2 36959 36974
0 36976 5 1 1 36975
0 36977 7 1 2 51124 36976
0 36978 5 1 1 36977
0 36979 7 1 2 68171 75747
0 36980 5 1 1 36979
0 36981 7 1 2 58981 36980
0 36982 5 1 1 36981
0 36983 7 1 2 61096 66977
0 36984 7 1 2 75539 36983
0 36985 5 1 1 36984
0 36986 7 1 2 36982 36985
0 36987 5 1 1 36986
0 36988 7 1 2 60557 36987
0 36989 5 1 1 36988
0 36990 7 1 2 3522 78364
0 36991 5 1 1 36990
0 36992 7 1 2 59551 63335
0 36993 5 1 1 36992
0 36994 7 1 2 36991 36993
0 36995 5 1 1 36994
0 36996 7 1 2 58626 36995
0 36997 5 1 1 36996
0 36998 7 1 2 36989 36997
0 36999 7 1 2 77060 78365
0 37000 5 1 1 36999
0 37001 7 1 2 60558 61242
0 37002 5 2 1 37001
0 37003 7 1 2 57187 63336
0 37004 5 1 1 37003
0 37005 7 1 2 78447 37004
0 37006 7 1 2 37000 37005
0 37007 5 1 1 37006
0 37008 7 1 2 55811 37007
0 37009 5 1 1 37008
0 37010 7 1 2 59404 78366
0 37011 5 1 1 37010
0 37012 7 1 2 78448 37011
0 37013 5 1 1 37012
0 37014 7 1 2 60001 37013
0 37015 5 1 1 37014
0 37016 7 1 2 60327 66209
0 37017 5 1 1 37016
0 37018 7 1 2 57043 37017
0 37019 5 1 1 37018
0 37020 7 1 2 56584 68313
0 37021 7 1 2 37019 37020
0 37022 5 1 1 37021
0 37023 7 1 2 37022 78332
0 37024 5 1 1 37023
0 37025 7 1 2 50841 68021
0 37026 5 1 1 37025
0 37027 7 1 2 60801 37026
0 37028 7 1 2 37024 37027
0 37029 5 1 1 37028
0 37030 7 1 2 37015 37029
0 37031 7 1 2 37009 37030
0 37032 7 1 2 36998 37031
0 37033 5 1 1 37032
0 37034 7 1 2 67187 37033
0 37035 5 1 1 37034
0 37036 7 1 2 36978 37035
0 37037 5 1 1 37036
0 37038 7 1 2 55386 37037
0 37039 5 1 1 37038
0 37040 7 1 2 36957 37039
0 37041 7 1 2 36877 37040
0 37042 5 1 1 37041
0 37043 7 1 2 49947 37042
0 37044 5 1 1 37043
0 37045 7 1 2 36685 37044
0 37046 5 1 1 37045
0 37047 7 1 2 56154 37046
0 37048 5 1 1 37047
0 37049 7 1 2 70398 74479
0 37050 5 1 1 37049
0 37051 7 1 2 51125 58982
0 37052 7 1 2 37050 37051
0 37053 5 1 1 37052
0 37054 7 1 2 64678 74293
0 37055 7 1 2 74724 37054
0 37056 5 1 1 37055
0 37057 7 1 2 37053 37056
0 37058 5 1 1 37057
0 37059 7 1 2 65991 37058
0 37060 5 1 1 37059
0 37061 7 1 2 62735 67738
0 37062 5 1 1 37061
0 37063 7 1 2 66332 37062
0 37064 5 1 1 37063
0 37065 7 1 2 62578 37064
0 37066 5 1 1 37065
0 37067 7 1 2 62937 63889
0 37068 5 1 1 37067
0 37069 7 1 2 37066 37068
0 37070 5 1 1 37069
0 37071 7 1 2 51626 37070
0 37072 5 1 1 37071
0 37073 7 1 2 63969 78437
0 37074 5 1 1 37073
0 37075 7 1 2 7858 37074
0 37076 5 1 1 37075
0 37077 7 1 2 55551 73825
0 37078 7 1 2 37076 37077
0 37079 5 1 1 37078
0 37080 7 1 2 37072 37079
0 37081 5 1 1 37080
0 37082 7 1 2 49246 37081
0 37083 5 1 1 37082
0 37084 7 1 2 64418 66123
0 37085 5 1 1 37084
0 37086 7 1 2 67986 37085
0 37087 5 1 1 37086
0 37088 7 1 2 71884 37087
0 37089 5 1 1 37088
0 37090 7 2 2 57530 78349
0 37091 7 1 2 54093 23338
0 37092 5 1 1 37091
0 37093 7 1 2 61580 37092
0 37094 7 1 2 78449 37093
0 37095 5 1 1 37094
0 37096 7 1 2 37089 37095
0 37097 5 1 1 37096
0 37098 7 1 2 54396 37097
0 37099 5 1 1 37098
0 37100 7 1 2 68429 74759
0 37101 5 1 1 37100
0 37102 7 2 2 73527 71066
0 37103 5 1 1 78451
0 37104 7 1 2 71767 78452
0 37105 5 2 1 37104
0 37106 7 1 2 37101 78453
0 37107 7 1 2 37099 37106
0 37108 5 1 1 37107
0 37109 7 1 2 48249 37108
0 37110 5 1 1 37109
0 37111 7 1 2 63643 71768
0 37112 5 1 1 37111
0 37113 7 1 2 78353 37112
0 37114 5 1 1 37113
0 37115 7 1 2 56585 37114
0 37116 5 1 1 37115
0 37117 7 1 2 68741 78345
0 37118 5 1 1 37117
0 37119 7 1 2 54094 37118
0 37120 5 1 1 37119
0 37121 7 1 2 37116 37120
0 37122 7 1 2 37110 37121
0 37123 7 1 2 37083 37122
0 37124 5 1 1 37123
0 37125 7 1 2 51392 37124
0 37126 5 1 1 37125
0 37127 7 1 2 37060 37126
0 37128 5 1 1 37127
0 37129 7 1 2 54777 37128
0 37130 5 1 1 37129
0 37131 7 1 2 74448 76490
0 37132 5 1 1 37131
0 37133 7 1 2 50514 65992
0 37134 7 1 2 58983 37133
0 37135 7 1 2 61842 37134
0 37136 5 1 1 37135
0 37137 7 1 2 37132 37136
0 37138 5 1 1 37137
0 37139 7 1 2 50842 37138
0 37140 5 1 1 37139
0 37141 7 1 2 55387 78334
0 37142 5 1 1 37141
0 37143 7 1 2 56586 74760
0 37144 7 1 2 71902 37143
0 37145 5 1 1 37144
0 37146 7 1 2 37142 37145
0 37147 5 1 1 37146
0 37148 7 1 2 67699 37147
0 37149 5 1 1 37148
0 37150 7 1 2 37140 37149
0 37151 5 1 1 37150
0 37152 7 1 2 55096 37151
0 37153 5 1 1 37152
0 37154 7 1 2 66847 74124
0 37155 5 1 1 37154
0 37156 7 1 2 62579 65604
0 37157 5 1 1 37156
0 37158 7 1 2 37155 37157
0 37159 5 1 1 37158
0 37160 7 1 2 71747 37159
0 37161 5 1 1 37160
0 37162 7 1 2 53561 67664
0 37163 7 2 2 67098 37162
0 37164 5 1 1 78455
0 37165 7 1 2 47992 78456
0 37166 5 1 1 37165
0 37167 7 1 2 64542 68430
0 37168 5 1 1 37167
0 37169 7 1 2 37166 37168
0 37170 5 1 1 37169
0 37171 7 1 2 51393 61581
0 37172 7 1 2 37170 37171
0 37173 5 1 1 37172
0 37174 7 1 2 37161 37173
0 37175 7 1 2 37153 37174
0 37176 7 1 2 37130 37175
0 37177 5 1 1 37176
0 37178 7 1 2 49948 37177
0 37179 5 1 1 37178
0 37180 7 2 2 64474 70229
0 37181 5 1 1 78457
0 37182 7 1 2 61763 78458
0 37183 5 1 1 37182
0 37184 7 1 2 66867 37183
0 37185 5 1 1 37184
0 37186 7 1 2 48250 37185
0 37187 5 1 1 37186
0 37188 7 1 2 64421 37187
0 37189 5 1 1 37188
0 37190 7 1 2 51126 37189
0 37191 5 1 1 37190
0 37192 7 1 2 62852 68876
0 37193 7 1 2 63033 37192
0 37194 5 1 1 37193
0 37195 7 1 2 37191 37194
0 37196 5 1 1 37195
0 37197 7 1 2 71675 37196
0 37198 5 1 1 37197
0 37199 7 1 2 74092 72422
0 37200 5 1 1 37199
0 37201 7 1 2 37198 37200
0 37202 5 1 1 37201
0 37203 7 1 2 68196 37202
0 37204 5 1 1 37203
0 37205 7 1 2 37179 37204
0 37206 5 1 1 37205
0 37207 7 1 2 55812 37206
0 37208 5 1 1 37207
0 37209 7 2 2 60002 71849
0 37210 7 1 2 78450 78459
0 37211 5 1 1 37210
0 37212 7 1 2 63338 67188
0 37213 5 1 1 37212
0 37214 7 1 2 37211 37213
0 37215 5 1 1 37214
0 37216 7 1 2 54397 37215
0 37217 5 1 1 37216
0 37218 7 1 2 17912 37217
0 37219 5 1 1 37218
0 37220 7 1 2 49247 37219
0 37221 5 1 1 37220
0 37222 7 1 2 71723 75535
0 37223 5 1 1 37222
0 37224 7 1 2 68742 78454
0 37225 5 1 1 37224
0 37226 7 1 2 47993 37225
0 37227 5 1 1 37226
0 37228 7 1 2 37223 37227
0 37229 7 1 2 37221 37228
0 37230 5 1 1 37229
0 37231 7 1 2 54778 37230
0 37232 5 1 1 37231
0 37233 7 1 2 63970 68431
0 37234 5 1 1 37233
0 37235 7 1 2 37164 37234
0 37236 5 1 1 37235
0 37237 7 1 2 61582 37236
0 37238 5 1 1 37237
0 37239 7 1 2 64679 70236
0 37240 7 1 2 71885 37239
0 37241 5 1 1 37240
0 37242 7 1 2 73826 69713
0 37243 7 1 2 59074 37242
0 37244 7 1 2 67360 37243
0 37245 5 1 1 37244
0 37246 7 1 2 37241 37245
0 37247 5 1 1 37246
0 37248 7 1 2 55097 37247
0 37249 5 1 1 37248
0 37250 7 1 2 37238 37249
0 37251 7 1 2 37232 37250
0 37252 5 1 1 37251
0 37253 7 1 2 51394 37252
0 37254 5 1 1 37253
0 37255 7 1 2 57846 61775
0 37256 5 1 1 37255
0 37257 7 1 2 64410 74294
0 37258 7 1 2 37256 37257
0 37259 5 1 1 37258
0 37260 7 1 2 62601 37259
0 37261 5 1 1 37260
0 37262 7 1 2 56587 37261
0 37263 5 1 1 37262
0 37264 7 1 2 72078 72544
0 37265 5 1 1 37264
0 37266 7 1 2 60559 74519
0 37267 5 1 1 37266
0 37268 7 1 2 37265 37267
0 37269 5 2 1 37268
0 37270 7 1 2 47994 78461
0 37271 5 1 1 37270
0 37272 7 1 2 74224 37271
0 37273 5 1 1 37272
0 37274 7 1 2 58984 37273
0 37275 5 1 1 37274
0 37276 7 1 2 37263 37275
0 37277 5 1 1 37276
0 37278 7 1 2 65993 37277
0 37279 5 1 1 37278
0 37280 7 1 2 37254 37279
0 37281 5 1 1 37280
0 37282 7 1 2 49949 37281
0 37283 5 1 1 37282
0 37284 7 1 2 71676 78462
0 37285 5 1 1 37284
0 37286 7 1 2 58177 71830
0 37287 7 1 2 74750 37286
0 37288 5 1 1 37287
0 37289 7 1 2 37285 37288
0 37290 5 1 1 37289
0 37291 7 1 2 47995 37290
0 37292 5 1 1 37291
0 37293 7 1 2 71677 74222
0 37294 5 1 1 37293
0 37295 7 1 2 37292 37294
0 37296 5 1 1 37295
0 37297 7 1 2 68197 37296
0 37298 5 1 1 37297
0 37299 7 1 2 37283 37298
0 37300 5 1 1 37299
0 37301 7 1 2 62066 37300
0 37302 5 1 1 37301
0 37303 7 1 2 52700 67758
0 37304 5 1 1 37303
0 37305 7 1 2 49248 58722
0 37306 7 1 2 65873 37305
0 37307 5 1 1 37306
0 37308 7 1 2 75711 77062
0 37309 7 1 2 37307 37308
0 37310 7 1 2 78225 37309
0 37311 5 1 1 37310
0 37312 7 1 2 51127 37311
0 37313 5 1 1 37312
0 37314 7 1 2 37304 37313
0 37315 5 1 1 37314
0 37316 7 1 2 71769 37315
0 37317 5 1 1 37316
0 37318 7 2 2 64404 78412
0 37319 5 2 1 78463
0 37320 7 1 2 65905 78465
0 37321 5 1 1 37320
0 37322 7 1 2 52567 64670
0 37323 5 1 1 37322
0 37324 7 2 2 60427 62273
0 37325 5 1 1 78467
0 37326 7 1 2 50843 78468
0 37327 5 1 1 37326
0 37328 7 1 2 37323 37327
0 37329 5 1 1 37328
0 37330 7 1 2 63462 65092
0 37331 5 1 1 37330
0 37332 7 1 2 6006 37331
0 37333 7 1 2 37329 37332
0 37334 5 1 1 37333
0 37335 7 1 2 57531 37334
0 37336 5 1 1 37335
0 37337 7 1 2 52568 65408
0 37338 5 1 1 37337
0 37339 7 1 2 55098 37338
0 37340 5 1 1 37339
0 37341 7 1 2 62975 37340
0 37342 7 1 2 37336 37341
0 37343 7 1 2 37321 37342
0 37344 5 1 1 37343
0 37345 7 1 2 71886 37344
0 37346 5 1 1 37345
0 37347 7 1 2 37317 37346
0 37348 5 1 1 37347
0 37349 7 1 2 49628 37348
0 37350 5 1 1 37349
0 37351 7 1 2 48667 61583
0 37352 5 1 1 37351
0 37353 7 1 2 49249 59530
0 37354 7 1 2 62263 37353
0 37355 7 1 2 77113 37354
0 37356 5 2 1 37355
0 37357 7 1 2 37352 78469
0 37358 5 1 1 37357
0 37359 7 1 2 51128 37358
0 37360 5 1 1 37359
0 37361 7 1 2 73204 76964
0 37362 5 1 1 37361
0 37363 7 1 2 66907 37362
0 37364 5 1 1 37363
0 37365 7 1 2 60136 37364
0 37366 5 1 1 37365
0 37367 7 1 2 37360 37366
0 37368 5 1 1 37367
0 37369 7 1 2 50515 37368
0 37370 5 1 1 37369
0 37371 7 1 2 65097 71850
0 37372 7 1 2 59533 37371
0 37373 5 1 1 37372
0 37374 7 1 2 75526 37373
0 37375 5 1 1 37374
0 37376 7 1 2 68297 37375
0 37377 5 1 1 37376
0 37378 7 1 2 37370 37377
0 37379 5 1 1 37378
0 37380 7 1 2 71770 37379
0 37381 5 1 1 37380
0 37382 7 1 2 57652 78464
0 37383 5 1 1 37382
0 37384 7 1 2 62938 37383
0 37385 5 1 1 37384
0 37386 7 1 2 48251 23407
0 37387 5 2 1 37386
0 37388 7 1 2 57532 15232
0 37389 5 1 1 37388
0 37390 7 1 2 78471 37389
0 37391 5 1 1 37390
0 37392 7 1 2 48668 65508
0 37393 7 1 2 37391 37392
0 37394 5 1 1 37393
0 37395 7 1 2 37385 37394
0 37396 5 1 1 37395
0 37397 7 1 2 51627 37396
0 37398 5 1 1 37397
0 37399 7 1 2 37381 37398
0 37400 5 1 1 37399
0 37401 7 1 2 54779 37400
0 37402 5 1 1 37401
0 37403 7 1 2 57653 78422
0 37404 5 1 1 37403
0 37405 7 1 2 61584 37404
0 37406 5 1 1 37405
0 37407 7 1 2 52569 61127
0 37408 7 1 2 37406 37407
0 37409 5 1 1 37408
0 37410 7 1 2 73205 37409
0 37411 5 1 1 37410
0 37412 7 1 2 57533 66903
0 37413 5 1 1 37412
0 37414 7 1 2 37411 37413
0 37415 5 1 1 37414
0 37416 7 1 2 78337 37415
0 37417 5 1 1 37416
0 37418 7 1 2 65509 64260
0 37419 5 1 1 37418
0 37420 7 1 2 62976 37419
0 37421 5 1 1 37420
0 37422 7 1 2 67152 37421
0 37423 5 1 1 37422
0 37424 7 1 2 49250 76206
0 37425 7 1 2 68436 37424
0 37426 5 1 1 37425
0 37427 7 1 2 37423 37426
0 37428 5 1 1 37427
0 37429 7 1 2 37325 37428
0 37430 5 1 1 37429
0 37431 7 1 2 52570 71930
0 37432 5 1 1 37431
0 37433 7 1 2 71840 37432
0 37434 5 1 1 37433
0 37435 7 1 2 51395 37434
0 37436 7 1 2 37430 37435
0 37437 7 1 2 37417 37436
0 37438 7 1 2 37402 37437
0 37439 7 1 2 37350 37438
0 37440 5 1 1 37439
0 37441 7 1 2 63975 78472
0 37442 5 1 1 37441
0 37443 7 1 2 49251 58985
0 37444 7 1 2 37442 37443
0 37445 5 1 1 37444
0 37446 7 1 2 61219 37445
0 37447 5 1 1 37446
0 37448 7 1 2 54780 37447
0 37449 5 1 1 37448
0 37450 7 1 2 60973 71803
0 37451 7 1 2 74125 37450
0 37452 5 1 1 37451
0 37453 7 1 2 61220 37452
0 37454 5 1 1 37453
0 37455 7 1 2 61585 37454
0 37456 5 1 1 37455
0 37457 7 1 2 51129 2739
0 37458 7 1 2 37456 37457
0 37459 7 1 2 37449 37458
0 37460 5 1 1 37459
0 37461 7 1 2 64680 68314
0 37462 7 1 2 78466 37461
0 37463 5 1 1 37462
0 37464 7 1 2 65406 61776
0 37465 5 1 1 37464
0 37466 7 1 2 47996 37465
0 37467 5 1 1 37466
0 37468 7 1 2 57654 61870
0 37469 7 1 2 37467 37468
0 37470 5 1 1 37469
0 37471 7 1 2 60560 58986
0 37472 7 1 2 37470 37471
0 37473 5 1 1 37472
0 37474 7 1 2 78335 78378
0 37475 5 1 1 37474
0 37476 7 1 2 55099 37475
0 37477 7 1 2 37473 37476
0 37478 7 1 2 37463 37477
0 37479 5 1 1 37478
0 37480 7 1 2 51628 37479
0 37481 7 1 2 37460 37480
0 37482 5 1 1 37481
0 37483 7 1 2 55388 35971
0 37484 7 1 2 37482 37483
0 37485 5 1 1 37484
0 37486 7 1 2 49950 37485
0 37487 7 1 2 37440 37486
0 37488 5 1 1 37487
0 37489 7 1 2 66124 75394
0 37490 5 1 1 37489
0 37491 7 1 2 57964 62116
0 37492 5 1 1 37491
0 37493 7 1 2 37490 37492
0 37494 5 1 1 37493
0 37495 7 1 2 70092 37494
0 37496 5 1 1 37495
0 37497 7 1 2 58987 73401
0 37498 5 1 1 37497
0 37499 7 1 2 62117 76536
0 37500 5 1 1 37499
0 37501 7 1 2 37498 37500
0 37502 7 1 2 37496 37501
0 37503 5 1 1 37502
0 37504 7 1 2 49951 37503
0 37505 5 1 1 37504
0 37506 7 1 2 64621 66909
0 37507 5 1 1 37506
0 37508 7 1 2 37505 37507
0 37509 5 1 1 37508
0 37510 7 1 2 57534 37509
0 37511 5 1 1 37510
0 37512 7 1 2 68704 69103
0 37513 7 1 2 65150 37512
0 37514 7 1 2 63264 37513
0 37515 5 1 1 37514
0 37516 7 1 2 37511 37515
0 37517 5 1 1 37516
0 37518 7 1 2 51629 37517
0 37519 5 1 1 37518
0 37520 7 1 2 62496 69104
0 37521 5 1 1 37520
0 37522 7 1 2 59713 74237
0 37523 7 1 2 61721 37522
0 37524 7 1 2 68198 37523
0 37525 5 1 1 37524
0 37526 7 1 2 37521 37525
0 37527 5 1 1 37526
0 37528 7 1 2 54781 37527
0 37529 5 1 1 37528
0 37530 7 2 2 56588 59596
0 37531 7 1 2 69317 78473
0 37532 7 1 2 69887 37531
0 37533 5 1 1 37532
0 37534 7 1 2 37529 37533
0 37535 5 1 1 37534
0 37536 7 1 2 66103 37535
0 37537 5 1 1 37536
0 37538 7 1 2 37519 37537
0 37539 5 1 1 37538
0 37540 7 1 2 64224 37539
0 37541 5 1 1 37540
0 37542 7 1 2 61586 65031
0 37543 5 1 1 37542
0 37544 7 1 2 63989 37543
0 37545 5 1 1 37544
0 37546 7 1 2 57535 37545
0 37547 5 1 1 37546
0 37548 7 1 2 65264 37547
0 37549 5 1 1 37548
0 37550 7 1 2 51130 37549
0 37551 5 1 1 37550
0 37552 7 1 2 61966 69427
0 37553 5 1 1 37552
0 37554 7 1 2 37551 37553
0 37555 5 1 1 37554
0 37556 7 1 2 48252 37555
0 37557 5 1 1 37556
0 37558 7 1 2 35728 35918
0 37559 5 1 1 37558
0 37560 7 1 2 60351 37559
0 37561 5 1 1 37560
0 37562 7 1 2 78397 37561
0 37563 7 1 2 37557 37562
0 37564 5 1 1 37563
0 37565 7 1 2 64622 66367
0 37566 7 1 2 37564 37565
0 37567 5 1 1 37566
0 37568 7 1 2 37541 37567
0 37569 7 1 2 37488 37568
0 37570 7 1 2 37302 37569
0 37571 7 1 2 37208 37570
0 37572 5 1 1 37571
0 37573 7 1 2 56411 37572
0 37574 5 1 1 37573
0 37575 7 1 2 37048 37574
0 37576 7 1 2 36554 37575
0 37577 5 1 1 37576
0 37578 7 1 2 48954 37577
0 37579 5 1 1 37578
0 37580 7 1 2 70334 78328
0 37581 5 3 1 37580
0 37582 7 1 2 66655 78475
0 37583 5 1 1 37582
0 37584 7 1 2 58058 70787
0 37585 5 1 1 37584
0 37586 7 1 2 72914 37585
0 37587 5 1 1 37586
0 37588 7 1 2 49781 37587
0 37589 5 1 1 37588
0 37590 7 1 2 37583 37589
0 37591 5 1 1 37590
0 37592 7 1 2 51396 37591
0 37593 5 1 1 37592
0 37594 7 1 2 67400 72707
0 37595 5 1 1 37594
0 37596 7 1 2 58988 37595
0 37597 5 2 1 37596
0 37598 7 1 2 63832 78478
0 37599 5 1 1 37598
0 37600 7 1 2 37593 37599
0 37601 5 1 1 37600
0 37602 7 1 2 49952 37601
0 37603 5 1 1 37602
0 37604 7 2 2 55943 57044
0 37605 5 2 1 78480
0 37606 7 1 2 61322 78482
0 37607 5 2 1 37606
0 37608 7 2 2 63833 78484
0 37609 7 1 2 68842 78486
0 37610 5 1 1 37609
0 37611 7 1 2 37603 37610
0 37612 5 1 1 37611
0 37613 7 1 2 48955 37612
0 37614 5 1 1 37613
0 37615 7 7 2 68774 70615
0 37616 5 1 1 78488
0 37617 7 1 2 78489 78487
0 37618 5 1 1 37617
0 37619 7 1 2 37614 37618
0 37620 5 1 1 37619
0 37621 7 1 2 55552 37620
0 37622 5 1 1 37621
0 37623 7 1 2 64199 67682
0 37624 7 1 2 72353 37623
0 37625 5 1 1 37624
0 37626 7 1 2 37622 37625
0 37627 5 1 1 37626
0 37628 7 1 2 60863 37627
0 37629 5 1 1 37628
0 37630 7 1 2 72445 76677
0 37631 5 1 1 37630
0 37632 7 2 2 55389 57045
0 37633 7 3 2 60729 78495
0 37634 7 1 2 58768 78497
0 37635 5 1 1 37634
0 37636 7 1 2 37631 37635
0 37637 5 1 1 37636
0 37638 7 1 2 53562 37637
0 37639 5 1 1 37638
0 37640 7 1 2 70603 78498
0 37641 5 1 1 37640
0 37642 7 1 2 37639 37641
0 37643 5 1 1 37642
0 37644 7 1 2 55100 37643
0 37645 5 1 1 37644
0 37646 7 1 2 60730 68589
0 37647 7 1 2 72824 37646
0 37648 5 1 1 37647
0 37649 7 1 2 37645 37648
0 37650 5 1 1 37649
0 37651 7 1 2 49953 37650
0 37652 5 1 1 37651
0 37653 7 2 2 55101 78499
0 37654 7 1 2 68843 78500
0 37655 5 1 1 37654
0 37656 7 1 2 37652 37655
0 37657 5 1 1 37656
0 37658 7 1 2 48956 37657
0 37659 5 1 1 37658
0 37660 7 1 2 78490 78501
0 37661 5 1 1 37660
0 37662 7 1 2 37659 37661
0 37663 5 1 1 37662
0 37664 7 1 2 57655 37663
0 37665 5 1 1 37664
0 37666 7 4 2 60517 73256
0 37667 5 1 1 78502
0 37668 7 1 2 55390 37667
0 37669 5 1 1 37668
0 37670 7 1 2 52571 37669
0 37671 5 1 1 37670
0 37672 7 2 2 72553 25307
0 37673 5 1 1 78506
0 37674 7 1 2 55944 37673
0 37675 5 1 1 37674
0 37676 7 1 2 51397 57357
0 37677 5 1 1 37676
0 37678 7 1 2 37675 37677
0 37679 7 1 2 37671 37678
0 37680 5 1 1 37679
0 37681 7 1 2 49782 37680
0 37682 5 1 1 37681
0 37683 7 2 2 49629 69806
0 37684 5 2 1 78508
0 37685 7 1 2 66046 78509
0 37686 5 1 1 37685
0 37687 7 1 2 61444 78510
0 37688 5 4 1 37687
0 37689 7 1 2 52572 78512
0 37690 5 1 1 37689
0 37691 7 1 2 22708 37690
0 37692 5 2 1 37691
0 37693 7 1 2 66656 78516
0 37694 5 1 1 37693
0 37695 7 1 2 37686 37694
0 37696 7 1 2 37682 37695
0 37697 5 1 1 37696
0 37698 7 2 2 51131 69620
0 37699 7 1 2 60731 78518
0 37700 7 1 2 37697 37699
0 37701 5 1 1 37700
0 37702 7 1 2 37665 37701
0 37703 5 1 1 37702
0 37704 7 1 2 51975 37703
0 37705 5 1 1 37704
0 37706 7 2 2 62977 67853
0 37707 5 2 1 78520
0 37708 7 2 2 49954 72708
0 37709 5 2 1 78524
0 37710 7 1 2 67848 78526
0 37711 5 1 1 37710
0 37712 7 2 2 78522 37711
0 37713 7 1 2 66657 78528
0 37714 5 1 1 37713
0 37715 7 2 2 66047 67987
0 37716 5 1 1 78530
0 37717 7 1 2 69621 78531
0 37718 5 1 1 37717
0 37719 7 1 2 37714 37718
0 37720 5 1 1 37719
0 37721 7 1 2 55102 37720
0 37722 5 1 1 37721
0 37723 7 1 2 69622 72323
0 37724 7 1 2 57332 37723
0 37725 7 1 2 59920 37724
0 37726 5 1 1 37725
0 37727 7 1 2 37722 37726
0 37728 5 1 1 37727
0 37729 7 1 2 55391 37728
0 37730 5 1 1 37729
0 37731 7 1 2 58122 70183
0 37732 7 1 2 78507 37731
0 37733 5 1 1 37732
0 37734 7 1 2 49783 37733
0 37735 5 1 1 37734
0 37736 7 1 2 76005 37735
0 37737 5 1 1 37736
0 37738 7 1 2 59921 37737
0 37739 5 1 1 37738
0 37740 7 2 2 48807 77751
0 37741 7 1 2 49784 78532
0 37742 5 1 1 37741
0 37743 7 1 2 70093 37742
0 37744 5 1 1 37743
0 37745 7 1 2 37739 37744
0 37746 5 1 1 37745
0 37747 7 1 2 69623 37746
0 37748 5 1 1 37747
0 37749 7 1 2 37730 37748
0 37750 5 1 1 37749
0 37751 7 1 2 60220 37750
0 37752 5 1 1 37751
0 37753 7 2 2 62978 69624
0 37754 7 1 2 78435 78534
0 37755 7 1 2 77756 37754
0 37756 5 1 1 37755
0 37757 7 1 2 37752 37756
0 37758 5 1 1 37757
0 37759 7 1 2 55705 37758
0 37760 5 1 1 37759
0 37761 7 1 2 72939 71308
0 37762 7 1 2 70951 37761
0 37763 7 1 2 78517 37762
0 37764 5 1 1 37763
0 37765 7 1 2 37760 37764
0 37766 7 1 2 37705 37765
0 37767 5 1 1 37766
0 37768 7 1 2 55553 37767
0 37769 5 1 1 37768
0 37770 7 1 2 37629 37769
0 37771 5 1 1 37770
0 37772 7 1 2 50844 37771
0 37773 5 1 1 37772
0 37774 7 1 2 64174 75723
0 37775 5 2 1 37774
0 37776 7 1 2 75249 78536
0 37777 5 1 1 37776
0 37778 7 2 2 57046 37777
0 37779 5 1 1 78538
0 37780 7 1 2 60668 75242
0 37781 5 1 1 37780
0 37782 7 2 2 48808 50269
0 37783 5 1 1 78540
0 37784 7 1 2 74834 71857
0 37785 5 1 1 37784
0 37786 7 1 2 37783 37785
0 37787 5 1 1 37786
0 37788 7 1 2 57333 37787
0 37789 5 1 1 37788
0 37790 7 1 2 37781 37789
0 37791 5 1 1 37790
0 37792 7 1 2 50516 37791
0 37793 5 1 1 37792
0 37794 7 1 2 37779 37793
0 37795 5 1 1 37794
0 37796 7 1 2 55103 37795
0 37797 5 1 1 37796
0 37798 7 3 2 63530 65806
0 37799 5 1 1 78542
0 37800 7 1 2 48809 78543
0 37801 5 1 1 37800
0 37802 7 1 2 37797 37801
0 37803 5 1 1 37802
0 37804 7 1 2 67872 37803
0 37805 5 1 1 37804
0 37806 7 1 2 70139 78544
0 37807 5 1 1 37806
0 37808 7 2 2 52906 68877
0 37809 7 3 2 71216 78545
0 37810 5 1 1 78547
0 37811 7 1 2 51976 78548
0 37812 5 1 1 37811
0 37813 7 1 2 37103 37812
0 37814 5 1 1 37813
0 37815 7 1 2 71193 37814
0 37816 5 1 1 37815
0 37817 7 1 2 37807 37816
0 37818 5 1 1 37817
0 37819 7 1 2 62979 37818
0 37820 5 1 1 37819
0 37821 7 1 2 61355 77738
0 37822 5 1 1 37821
0 37823 7 1 2 77648 37822
0 37824 5 1 1 37823
0 37825 7 1 2 55104 37824
0 37826 5 1 1 37825
0 37827 7 1 2 37799 37826
0 37828 5 1 1 37827
0 37829 7 1 2 62497 37828
0 37830 5 1 1 37829
0 37831 7 1 2 37820 37830
0 37832 5 1 1 37831
0 37833 7 1 2 69625 37832
0 37834 5 1 1 37833
0 37835 7 1 2 37805 37834
0 37836 5 1 1 37835
0 37837 7 1 2 55392 37836
0 37838 5 1 1 37837
0 37839 7 2 2 51398 69626
0 37840 7 2 2 49785 67731
0 37841 7 1 2 65807 78552
0 37842 5 1 1 37841
0 37843 7 1 2 64240 74295
0 37844 5 3 1 37843
0 37845 7 1 2 70335 78554
0 37846 5 3 1 37845
0 37847 7 1 2 77739 78557
0 37848 5 1 1 37847
0 37849 7 1 2 37842 37848
0 37850 5 1 1 37849
0 37851 7 1 2 57047 37850
0 37852 5 1 1 37851
0 37853 7 1 2 61445 78555
0 37854 5 3 1 37853
0 37855 7 1 2 57334 78560
0 37856 5 1 1 37855
0 37857 7 1 2 23759 37856
0 37858 7 1 2 37852 37857
0 37859 5 1 1 37858
0 37860 7 1 2 78550 37859
0 37861 5 1 1 37860
0 37862 7 1 2 37838 37861
0 37863 5 1 1 37862
0 37864 7 1 2 57656 37863
0 37865 5 1 1 37864
0 37866 7 1 2 66643 77743
0 37867 5 2 1 37866
0 37868 7 1 2 70076 78563
0 37869 5 1 1 37868
0 37870 7 1 2 55105 60249
0 37871 7 1 2 65808 37870
0 37872 7 1 2 77895 37871
0 37873 5 1 1 37872
0 37874 7 1 2 37869 37873
0 37875 5 1 1 37874
0 37876 7 1 2 67873 37875
0 37877 5 1 1 37876
0 37878 7 1 2 67401 67988
0 37879 7 1 2 77740 37878
0 37880 5 1 1 37879
0 37881 7 1 2 72709 78564
0 37882 5 1 1 37881
0 37883 7 1 2 37716 37882
0 37884 7 1 2 37880 37883
0 37885 5 1 1 37884
0 37886 7 1 2 78519 37885
0 37887 5 1 1 37886
0 37888 7 1 2 37877 37887
0 37889 5 1 1 37888
0 37890 7 1 2 64598 37889
0 37891 5 1 1 37890
0 37892 7 1 2 55945 61356
0 37893 5 1 1 37892
0 37894 7 1 2 77649 37893
0 37895 5 1 1 37894
0 37896 7 1 2 77741 37895
0 37897 5 1 1 37896
0 37898 7 1 2 78533 37897
0 37899 5 1 1 37898
0 37900 7 1 2 49786 37899
0 37901 5 1 1 37900
0 37902 7 1 2 63217 37901
0 37903 5 1 1 37902
0 37904 7 1 2 63489 71080
0 37905 7 1 2 37903 37904
0 37906 5 1 1 37905
0 37907 7 1 2 37891 37906
0 37908 7 1 2 37865 37907
0 37909 5 1 1 37908
0 37910 7 1 2 55554 37909
0 37911 5 1 1 37910
0 37912 7 3 2 51630 64572
0 37913 5 1 1 78565
0 37914 7 3 2 69627 78566
0 37915 5 1 1 78568
0 37916 7 1 2 62580 67849
0 37917 5 1 1 37916
0 37918 7 5 2 21449 37917
0 37919 7 2 2 22299 78571
0 37920 7 1 2 53393 78576
0 37921 5 1 1 37920
0 37922 7 1 2 70594 72589
0 37923 5 1 1 37922
0 37924 7 1 2 37921 37923
0 37925 5 1 1 37924
0 37926 7 1 2 55555 37925
0 37927 5 1 1 37926
0 37928 7 1 2 37915 37927
0 37929 5 1 1 37928
0 37930 7 1 2 66658 37929
0 37931 5 1 1 37930
0 37932 7 1 2 66048 72136
0 37933 7 1 2 78525 37932
0 37934 5 1 1 37933
0 37935 7 1 2 37931 37934
0 37936 5 1 1 37935
0 37937 7 1 2 55393 37936
0 37938 5 1 1 37937
0 37939 7 1 2 57307 78483
0 37940 5 4 1 37939
0 37941 7 3 2 72324 78578
0 37942 7 2 2 69628 78582
0 37943 7 1 2 74265 78585
0 37944 5 1 1 37943
0 37945 7 1 2 37938 37944
0 37946 5 1 1 37945
0 37947 7 1 2 55106 37946
0 37948 5 1 1 37947
0 37949 7 1 2 58769 67402
0 37950 5 1 1 37949
0 37951 7 1 2 58123 37950
0 37952 5 1 1 37951
0 37953 7 1 2 49787 37952
0 37954 5 1 1 37953
0 37955 7 1 2 76006 37954
0 37956 5 1 1 37955
0 37957 7 1 2 75050 37956
0 37958 5 1 1 37957
0 37959 7 1 2 37948 37958
0 37960 5 1 1 37959
0 37961 7 1 2 65809 37960
0 37962 5 1 1 37961
0 37963 7 1 2 56963 77744
0 37964 5 1 1 37963
0 37965 7 2 2 63834 78567
0 37966 5 1 1 78587
0 37967 7 2 2 69629 78588
0 37968 7 1 2 57657 78589
0 37969 7 1 2 37964 37968
0 37970 5 1 1 37969
0 37971 7 1 2 37962 37970
0 37972 7 1 2 37911 37971
0 37973 7 1 2 37773 37972
0 37974 5 1 1 37973
0 37975 7 1 2 57250 37974
0 37976 5 1 1 37975
0 37977 7 1 2 68878 78529
0 37978 5 1 1 37977
0 37979 7 2 2 72960 68955
0 37980 7 1 2 54095 51132
0 37981 7 1 2 78591 37980
0 37982 7 1 2 67989 37981
0 37983 5 1 1 37982
0 37984 7 1 2 37978 37983
0 37985 5 1 1 37984
0 37986 7 1 2 55394 37985
0 37987 5 1 1 37986
0 37988 7 1 2 72961 68775
0 37989 7 1 2 73295 37988
0 37990 5 1 1 37989
0 37991 7 1 2 37987 37990
0 37992 5 1 1 37991
0 37993 7 1 2 50845 37992
0 37994 5 1 1 37993
0 37995 7 2 2 51399 67732
0 37996 7 1 2 50270 74546
0 37997 7 1 2 78593 37996
0 37998 5 1 1 37997
0 37999 7 1 2 37994 37998
0 38000 5 1 1 37999
0 38001 7 1 2 57048 38000
0 38002 5 1 1 38001
0 38003 7 1 2 73619 76578
0 38004 5 1 1 38003
0 38005 7 1 2 68796 38004
0 38006 5 1 1 38005
0 38007 7 1 2 48810 38006
0 38008 5 1 1 38007
0 38009 7 10 2 55395 62980
0 38010 7 1 2 75444 78595
0 38011 5 1 1 38010
0 38012 7 1 2 70292 78513
0 38013 5 1 1 38012
0 38014 7 1 2 38011 38013
0 38015 5 1 1 38014
0 38016 7 1 2 57335 38015
0 38017 5 1 1 38016
0 38018 7 1 2 63583 73136
0 38019 5 1 1 38018
0 38020 7 1 2 70293 75492
0 38021 5 1 1 38020
0 38022 7 1 2 74353 38021
0 38023 5 1 1 38022
0 38024 7 1 2 75922 38023
0 38025 5 1 1 38024
0 38026 7 1 2 38019 38025
0 38027 7 1 2 38017 38026
0 38028 5 1 1 38027
0 38029 7 1 2 49955 38028
0 38030 5 1 1 38029
0 38031 7 1 2 38008 38030
0 38032 5 1 1 38031
0 38033 7 1 2 50271 38032
0 38034 5 1 1 38033
0 38035 7 1 2 69312 73613
0 38036 7 1 2 73244 38035
0 38037 5 1 1 38036
0 38038 7 1 2 38034 38037
0 38039 5 1 1 38038
0 38040 7 1 2 51133 38039
0 38041 5 1 1 38040
0 38042 7 1 2 49630 64713
0 38043 5 1 1 38042
0 38044 7 1 2 53563 38043
0 38045 5 1 1 38044
0 38046 7 1 2 50517 78018
0 38047 7 1 2 38045 38046
0 38048 7 1 2 70958 38047
0 38049 5 1 1 38048
0 38050 7 1 2 38041 38049
0 38051 5 1 1 38050
0 38052 7 1 2 48957 38051
0 38053 5 1 1 38052
0 38054 7 1 2 71424 68399
0 38055 7 1 2 78491 38054
0 38056 5 1 1 38055
0 38057 7 1 2 38053 38056
0 38058 7 1 2 38002 38057
0 38059 5 1 1 38058
0 38060 7 1 2 57658 38059
0 38061 5 1 1 38060
0 38062 7 2 2 63835 67874
0 38063 7 1 2 64175 71425
0 38064 7 1 2 66049 38063
0 38065 5 1 1 38064
0 38066 7 1 2 48811 61502
0 38067 7 1 2 78485 38066
0 38068 5 1 1 38067
0 38069 7 1 2 38065 38068
0 38070 5 1 1 38069
0 38071 7 1 2 78605 38070
0 38072 5 1 1 38071
0 38073 7 1 2 63687 15456
0 38074 5 1 1 38073
0 38075 7 2 2 67403 38074
0 38076 5 1 1 78607
0 38077 7 1 2 63272 68022
0 38078 7 1 2 78481 38077
0 38079 5 1 1 38078
0 38080 7 1 2 70897 38079
0 38081 5 2 1 38080
0 38082 7 1 2 51977 78609
0 38083 5 1 1 38082
0 38084 7 1 2 2120 38083
0 38085 5 1 1 38084
0 38086 7 2 2 50846 38085
0 38087 5 1 1 78611
0 38088 7 1 2 25315 38087
0 38089 5 1 1 38088
0 38090 7 1 2 58059 38089
0 38091 5 1 1 38090
0 38092 7 1 2 38076 38091
0 38093 5 1 1 38092
0 38094 7 1 2 51400 38093
0 38095 5 1 1 38094
0 38096 7 3 2 51978 67531
0 38097 5 1 1 78613
0 38098 7 2 2 55946 70660
0 38099 5 1 1 78616
0 38100 7 1 2 38097 38099
0 38101 5 1 1 38100
0 38102 7 1 2 58770 60561
0 38103 7 1 2 38101 38102
0 38104 5 1 1 38103
0 38105 7 1 2 38095 38104
0 38106 5 1 1 38105
0 38107 7 1 2 49788 38106
0 38108 5 1 1 38107
0 38109 7 1 2 49631 73757
0 38110 5 2 1 38109
0 38111 7 1 2 52328 78161
0 38112 7 1 2 71194 38111
0 38113 7 1 2 78596 38112
0 38114 5 1 1 38113
0 38115 7 1 2 67817 38114
0 38116 5 1 1 38115
0 38117 7 1 2 78618 38116
0 38118 5 1 1 38117
0 38119 7 1 2 70554 77603
0 38120 5 1 1 38119
0 38121 7 1 2 62581 38120
0 38122 5 1 1 38121
0 38123 7 1 2 77956 38122
0 38124 5 1 1 38123
0 38125 7 1 2 68705 78583
0 38126 5 1 1 38125
0 38127 7 1 2 38124 38126
0 38128 5 1 1 38127
0 38129 7 1 2 55107 38128
0 38130 5 1 1 38129
0 38131 7 1 2 38118 38130
0 38132 5 1 1 38131
0 38133 7 1 2 50272 38132
0 38134 5 1 1 38133
0 38135 7 1 2 77495 78479
0 38136 5 1 1 38135
0 38137 7 2 2 61299 70661
0 38138 7 1 2 72325 78620
0 38139 5 1 1 38138
0 38140 7 1 2 38136 38139
0 38141 5 1 1 38140
0 38142 7 1 2 63789 38141
0 38143 5 1 1 38142
0 38144 7 1 2 38134 38143
0 38145 7 1 2 38108 38144
0 38146 5 1 1 38145
0 38147 7 1 2 69630 38146
0 38148 5 1 1 38147
0 38149 7 1 2 38072 38148
0 38150 7 1 2 38061 38149
0 38151 5 1 1 38150
0 38152 7 1 2 57251 38151
0 38153 5 1 1 38152
0 38154 7 1 2 75456 78004
0 38155 5 1 1 38154
0 38156 7 3 2 50518 59904
0 38157 5 1 1 78622
0 38158 7 2 2 58060 78623
0 38159 5 1 1 78625
0 38160 7 2 2 54782 78626
0 38161 5 1 1 78627
0 38162 7 1 2 70643 78628
0 38163 5 1 1 38162
0 38164 7 1 2 38155 38163
0 38165 5 1 1 38164
0 38166 7 1 2 50273 38165
0 38167 5 1 1 38166
0 38168 7 1 2 67725 70999
0 38169 5 2 1 38168
0 38170 7 1 2 73805 78629
0 38171 5 1 1 38170
0 38172 7 1 2 63531 38171
0 38173 5 1 1 38172
0 38174 7 1 2 58074 68879
0 38175 5 1 1 38174
0 38176 7 1 2 58075 77496
0 38177 5 1 1 38176
0 38178 7 1 2 50274 75614
0 38179 5 1 1 38178
0 38180 7 1 2 38177 38179
0 38181 5 1 1 38180
0 38182 7 1 2 70399 38181
0 38183 5 1 1 38182
0 38184 7 1 2 38175 38183
0 38185 7 1 2 38173 38184
0 38186 7 1 2 38167 38185
0 38187 5 1 1 38186
0 38188 7 1 2 53564 38187
0 38189 5 1 1 38188
0 38190 7 1 2 73765 78630
0 38191 5 1 1 38190
0 38192 7 1 2 63532 38191
0 38193 5 1 1 38192
0 38194 7 1 2 50847 75839
0 38195 5 1 1 38194
0 38196 7 1 2 38161 38195
0 38197 5 1 1 38196
0 38198 7 1 2 70644 38197
0 38199 5 1 1 38198
0 38200 7 1 2 60823 68880
0 38201 7 1 2 71293 38200
0 38202 5 1 1 38201
0 38203 7 1 2 38199 38202
0 38204 5 1 1 38203
0 38205 7 1 2 50275 38204
0 38206 5 1 1 38205
0 38207 7 1 2 38193 38206
0 38208 5 1 1 38207
0 38209 7 1 2 52701 38208
0 38210 5 1 1 38209
0 38211 7 1 2 38189 38210
0 38212 5 1 1 38211
0 38213 7 1 2 57049 38212
0 38214 5 1 1 38213
0 38215 7 1 2 55108 71480
0 38216 5 1 1 38215
0 38217 7 1 2 77434 38216
0 38218 5 1 1 38217
0 38219 7 1 2 63766 38218
0 38220 5 1 1 38219
0 38221 7 3 2 52702 50519
0 38222 5 1 1 78631
0 38223 7 1 2 77497 78632
0 38224 5 1 1 38223
0 38225 7 1 2 50848 76018
0 38226 5 1 1 38225
0 38227 7 1 2 38224 38226
0 38228 5 1 1 38227
0 38229 7 1 2 56649 38228
0 38230 5 1 1 38229
0 38231 7 1 2 24190 38230
0 38232 7 1 2 38220 38231
0 38233 5 1 1 38232
0 38234 7 1 2 50276 38233
0 38235 5 1 1 38234
0 38236 7 1 2 70683 75445
0 38237 7 1 2 72925 38236
0 38238 5 1 1 38237
0 38239 7 1 2 55109 73476
0 38240 5 1 1 38239
0 38241 7 1 2 77435 38240
0 38242 5 1 1 38241
0 38243 7 1 2 72920 38242
0 38244 5 1 1 38243
0 38245 7 1 2 55110 71300
0 38246 7 1 2 65356 38245
0 38247 5 1 1 38246
0 38248 7 1 2 38244 38247
0 38249 7 1 2 38238 38248
0 38250 7 1 2 38235 38249
0 38251 5 1 1 38250
0 38252 7 1 2 53565 38251
0 38253 5 1 1 38252
0 38254 7 1 2 54783 75059
0 38255 7 1 2 73012 38254
0 38256 5 1 1 38255
0 38257 7 1 2 38253 38256
0 38258 5 1 1 38257
0 38259 7 1 2 57336 38258
0 38260 5 1 1 38259
0 38261 7 1 2 51979 76391
0 38262 5 1 1 38261
0 38263 7 1 2 63548 38262
0 38264 5 1 1 38263
0 38265 7 1 2 70400 38264
0 38266 5 1 1 38265
0 38267 7 1 2 59944 63533
0 38268 5 2 1 38267
0 38269 7 1 2 38266 78634
0 38270 5 1 1 38269
0 38271 7 1 2 50520 38270
0 38272 5 1 1 38271
0 38273 7 1 2 72963 72967
0 38274 5 1 1 38273
0 38275 7 1 2 72912 73931
0 38276 5 1 1 38275
0 38277 7 1 2 73206 38276
0 38278 5 1 1 38277
0 38279 7 1 2 38274 38278
0 38280 7 1 2 38272 38279
0 38281 5 1 1 38280
0 38282 7 1 2 76540 38281
0 38283 5 1 1 38282
0 38284 7 1 2 55396 38283
0 38285 7 1 2 38260 38284
0 38286 7 1 2 38214 38285
0 38287 5 1 1 38286
0 38288 7 1 2 52703 78579
0 38289 5 1 1 38288
0 38290 7 1 2 73883 71630
0 38291 5 1 1 38290
0 38292 7 1 2 38289 38291
0 38293 5 1 1 38292
0 38294 7 1 2 49789 38293
0 38295 5 1 1 38294
0 38296 7 1 2 63463 78584
0 38297 5 1 1 38296
0 38298 7 1 2 38295 38297
0 38299 5 1 1 38298
0 38300 7 1 2 56650 38299
0 38301 5 1 1 38300
0 38302 7 1 2 75992 78580
0 38303 5 1 1 38302
0 38304 7 1 2 55111 28691
0 38305 5 2 1 38304
0 38306 7 1 2 49790 2519
0 38307 7 1 2 57050 38306
0 38308 7 1 2 77790 38307
0 38309 5 1 1 38308
0 38310 7 1 2 75929 38309
0 38311 5 1 1 38310
0 38312 7 1 2 78636 38311
0 38313 5 1 1 38312
0 38314 7 1 2 38303 38313
0 38315 7 1 2 38301 38314
0 38316 5 1 1 38315
0 38317 7 1 2 51980 38316
0 38318 5 1 1 38317
0 38319 7 1 2 2150 66059
0 38320 5 1 1 38319
0 38321 7 1 2 63615 38320
0 38322 5 1 1 38321
0 38323 7 1 2 38222 38322
0 38324 5 1 1 38323
0 38325 7 1 2 58061 38324
0 38326 5 1 1 38325
0 38327 7 1 2 50521 63703
0 38328 7 1 2 66050 38327
0 38329 5 1 1 38328
0 38330 7 1 2 38326 38329
0 38331 5 1 1 38330
0 38332 7 1 2 49791 38331
0 38333 5 1 1 38332
0 38334 7 1 2 252 63708
0 38335 5 1 1 38334
0 38336 7 1 2 49792 38335
0 38337 5 1 1 38336
0 38338 7 1 2 64241 76256
0 38339 5 1 1 38338
0 38340 7 1 2 38337 38339
0 38341 5 1 1 38340
0 38342 7 1 2 67404 38341
0 38343 5 1 1 38342
0 38344 7 1 2 64242 75428
0 38345 5 1 1 38344
0 38346 7 1 2 75250 38345
0 38347 5 1 1 38346
0 38348 7 1 2 63662 38347
0 38349 5 1 1 38348
0 38350 7 1 2 51401 38349
0 38351 7 1 2 38343 38350
0 38352 7 1 2 38333 38351
0 38353 7 1 2 38318 38352
0 38354 5 1 1 38353
0 38355 7 1 2 38287 38354
0 38356 5 1 1 38355
0 38357 7 1 2 73000 78553
0 38358 5 1 1 38357
0 38359 7 1 2 73573 78558
0 38360 5 1 1 38359
0 38361 7 1 2 38358 38360
0 38362 5 1 1 38361
0 38363 7 1 2 51402 38362
0 38364 5 1 1 38363
0 38365 7 2 2 59156 78284
0 38366 7 1 2 50277 78638
0 38367 5 1 1 38366
0 38368 7 1 2 38364 38367
0 38369 5 1 1 38368
0 38370 7 1 2 57051 38369
0 38371 5 1 1 38370
0 38372 7 1 2 48812 15509
0 38373 5 1 1 38372
0 38374 7 1 2 51981 38373
0 38375 5 1 1 38374
0 38376 7 1 2 63616 78637
0 38377 5 1 1 38376
0 38378 7 1 2 38375 38377
0 38379 5 1 1 38378
0 38380 7 1 2 57337 38379
0 38381 5 1 1 38380
0 38382 7 4 2 65343 60127
0 38383 5 2 1 78640
0 38384 7 1 2 54784 78644
0 38385 5 2 1 38384
0 38386 7 4 2 50278 78646
0 38387 5 1 1 78648
0 38388 7 1 2 71114 78649
0 38389 5 1 1 38388
0 38390 7 1 2 73174 28784
0 38391 5 1 1 38390
0 38392 7 1 2 75923 38391
0 38393 5 1 1 38392
0 38394 7 1 2 38389 38393
0 38395 7 1 2 38381 38394
0 38396 5 1 1 38395
0 38397 7 1 2 49793 38396
0 38398 5 1 1 38397
0 38399 7 2 2 69783 75345
0 38400 7 1 2 57338 78652
0 38401 5 1 1 38400
0 38402 7 1 2 73847 78147
0 38403 5 1 1 38402
0 38404 7 1 2 48813 77511
0 38405 5 1 1 38404
0 38406 7 1 2 38403 38405
0 38407 5 1 1 38406
0 38408 7 1 2 53566 38407
0 38409 5 1 1 38408
0 38410 7 1 2 38401 38409
0 38411 7 1 2 38398 38410
0 38412 5 1 1 38411
0 38413 7 1 2 51403 38412
0 38414 5 1 1 38413
0 38415 7 1 2 38371 38414
0 38416 5 1 1 38415
0 38417 7 1 2 57659 38416
0 38418 5 1 1 38417
0 38419 7 1 2 58771 78647
0 38420 5 1 1 38419
0 38421 7 1 2 38420 38159
0 38422 5 1 1 38421
0 38423 7 1 2 49794 38422
0 38424 5 1 1 38423
0 38425 7 1 2 50522 61254
0 38426 5 1 1 38425
0 38427 7 3 2 55112 72326
0 38428 7 1 2 62880 78654
0 38429 7 1 2 38426 38428
0 38430 5 1 1 38429
0 38431 7 1 2 38424 38430
0 38432 5 1 1 38431
0 38433 7 1 2 51404 38432
0 38434 5 1 1 38433
0 38435 7 1 2 56651 78639
0 38436 5 1 1 38435
0 38437 7 1 2 38434 38436
0 38438 5 1 1 38437
0 38439 7 1 2 50279 38438
0 38440 5 1 1 38439
0 38441 7 1 2 65344 73315
0 38442 7 1 2 78594 38441
0 38443 5 1 1 38442
0 38444 7 1 2 38440 38443
0 38445 5 1 1 38444
0 38446 7 1 2 66659 38445
0 38447 5 1 1 38446
0 38448 7 1 2 58772 73891
0 38449 7 1 2 77352 38448
0 38450 5 1 1 38449
0 38451 7 1 2 38447 38450
0 38452 7 1 2 38418 38451
0 38453 7 1 2 38356 38452
0 38454 5 1 1 38453
0 38455 7 1 2 69631 38454
0 38456 5 1 1 38455
0 38457 7 1 2 70645 71858
0 38458 5 1 1 38457
0 38459 7 1 2 70823 78541
0 38460 5 1 1 38459
0 38461 7 1 2 38458 38460
0 38462 5 1 1 38461
0 38463 7 1 2 50523 38462
0 38464 5 1 1 38463
0 38465 7 1 2 48814 63617
0 38466 5 1 1 38465
0 38467 7 1 2 64176 70472
0 38468 7 1 2 77854 38467
0 38469 5 1 1 38468
0 38470 7 1 2 38466 38469
0 38471 7 1 2 38464 38470
0 38472 5 1 1 38471
0 38473 7 1 2 57339 38472
0 38474 5 1 1 38473
0 38475 7 1 2 73936 75243
0 38476 5 1 1 38475
0 38477 7 1 2 63618 70646
0 38478 5 1 1 38477
0 38479 7 1 2 71017 78641
0 38480 5 1 1 38479
0 38481 7 1 2 38478 38480
0 38482 5 1 1 38481
0 38483 7 1 2 48815 38482
0 38484 5 1 1 38483
0 38485 7 1 2 75251 78154
0 38486 5 1 1 38485
0 38487 7 1 2 75454 38486
0 38488 5 1 1 38487
0 38489 7 1 2 38484 38488
0 38490 5 1 1 38489
0 38491 7 1 2 57052 38490
0 38492 5 1 1 38491
0 38493 7 1 2 38476 38492
0 38494 7 1 2 38474 38493
0 38495 5 1 1 38494
0 38496 7 1 2 55113 38495
0 38497 5 1 1 38496
0 38498 7 2 2 51982 66660
0 38499 5 1 1 78657
0 38500 7 1 2 73006 15216
0 38501 7 1 2 38499 38500
0 38502 5 1 1 38501
0 38503 7 1 2 78145 38502
0 38504 5 1 1 38503
0 38505 7 1 2 38497 38504
0 38506 5 1 1 38505
0 38507 7 1 2 55397 67875
0 38508 7 1 2 38506 38507
0 38509 5 1 1 38508
0 38510 7 1 2 38456 38509
0 38511 7 1 2 38153 38510
0 38512 5 1 1 38511
0 38513 7 1 2 55556 38512
0 38514 5 1 1 38513
0 38515 7 1 2 48816 78619
0 38516 5 2 1 38515
0 38517 7 1 2 78659 78537
0 38518 5 1 1 38517
0 38519 7 1 2 67876 38518
0 38520 5 1 1 38519
0 38521 7 1 2 70294 72710
0 38522 5 1 1 38521
0 38523 7 1 2 58989 38522
0 38524 5 1 1 38523
0 38525 7 1 2 69632 38524
0 38526 5 1 1 38525
0 38527 7 1 2 38520 38526
0 38528 5 1 1 38527
0 38529 7 1 2 76583 38528
0 38530 5 1 1 38529
0 38531 7 2 2 66282 72327
0 38532 7 1 2 78592 78661
0 38533 5 1 1 38532
0 38534 7 1 2 38530 38533
0 38535 5 1 1 38534
0 38536 7 1 2 55114 38535
0 38537 5 1 1 38536
0 38538 7 1 2 67733 78633
0 38539 5 1 1 38538
0 38540 7 2 2 51405 73803
0 38541 5 1 1 78663
0 38542 7 1 2 38539 38541
0 38543 5 1 1 38542
0 38544 7 1 2 49795 38543
0 38545 5 1 1 38544
0 38546 7 1 2 52573 64821
0 38547 5 1 1 38546
0 38548 7 1 2 75252 38547
0 38549 5 7 1 38548
0 38550 7 1 2 53567 63644
0 38551 7 1 2 78665 38550
0 38552 5 1 1 38551
0 38553 7 1 2 38545 38552
0 38554 5 1 1 38553
0 38555 7 1 2 48958 69313
0 38556 7 1 2 38554 38555
0 38557 5 1 1 38556
0 38558 7 1 2 38537 38557
0 38559 5 1 1 38558
0 38560 7 1 2 55557 38559
0 38561 5 1 1 38560
0 38562 7 1 2 65281 68676
0 38563 7 1 2 73536 38562
0 38564 5 1 1 38563
0 38565 7 1 2 38561 38564
0 38566 5 1 1 38565
0 38567 7 1 2 66661 38566
0 38568 5 1 1 38567
0 38569 7 2 2 67629 75346
0 38570 5 1 1 78672
0 38571 7 1 2 67901 73594
0 38572 7 1 2 78673 38571
0 38573 5 1 1 38572
0 38574 7 1 2 38568 38573
0 38575 5 1 1 38574
0 38576 7 1 2 57252 38575
0 38577 5 1 1 38576
0 38578 7 1 2 70401 78242
0 38579 5 1 1 38578
0 38580 7 1 2 71008 38579
0 38581 5 1 1 38580
0 38582 7 1 2 51983 38581
0 38583 5 1 1 38582
0 38584 7 1 2 50524 78279
0 38585 5 1 1 38584
0 38586 7 1 2 63633 38585
0 38587 7 1 2 38583 38586
0 38588 5 1 1 38587
0 38589 7 1 2 78590 38588
0 38590 5 1 1 38589
0 38591 7 1 2 38577 38590
0 38592 7 1 2 38514 38591
0 38593 5 1 1 38592
0 38594 7 1 2 58447 38593
0 38595 5 1 1 38594
0 38596 7 1 2 60497 73338
0 38597 5 1 1 38596
0 38598 7 1 2 50280 78011
0 38599 5 1 1 38598
0 38600 7 1 2 38597 38599
0 38601 5 1 1 38600
0 38602 7 1 2 48817 38601
0 38603 5 1 1 38602
0 38604 7 1 2 24874 37810
0 38605 5 1 1 38604
0 38606 7 1 2 69807 38605
0 38607 5 1 1 38606
0 38608 7 1 2 55398 78549
0 38609 5 1 1 38608
0 38610 7 1 2 51134 75123
0 38611 5 1 1 38610
0 38612 7 1 2 38609 38611
0 38613 5 1 1 38612
0 38614 7 1 2 52704 38613
0 38615 5 1 1 38614
0 38616 7 1 2 38607 38615
0 38617 5 2 1 38616
0 38618 7 1 2 52574 78674
0 38619 5 1 1 38618
0 38620 7 2 2 63809 73112
0 38621 7 1 2 53568 78676
0 38622 5 1 1 38621
0 38623 7 1 2 76598 38622
0 38624 5 2 1 38623
0 38625 7 1 2 52705 78678
0 38626 5 1 1 38625
0 38627 7 1 2 38619 38626
0 38628 5 1 1 38627
0 38629 7 1 2 49956 38628
0 38630 5 1 1 38629
0 38631 7 1 2 38603 38630
0 38632 5 1 1 38631
0 38633 7 1 2 48959 38632
0 38634 5 1 1 38633
0 38635 7 1 2 78492 78677
0 38636 5 1 1 38635
0 38637 7 1 2 38634 38636
0 38638 5 1 1 38637
0 38639 7 1 2 57053 38638
0 38640 5 1 1 38639
0 38641 7 1 2 66354 78261
0 38642 5 1 1 38641
0 38643 7 1 2 59894 38642
0 38644 5 1 1 38643
0 38645 7 1 2 58062 38644
0 38646 5 1 1 38645
0 38647 7 1 2 55706 58794
0 38648 5 1 1 38647
0 38649 7 1 2 65477 70893
0 38650 5 2 1 38649
0 38651 7 1 2 38648 78680
0 38652 7 1 2 38646 38651
0 38653 5 1 1 38652
0 38654 7 1 2 49796 38653
0 38655 5 1 1 38654
0 38656 7 1 2 54096 55707
0 38657 7 1 2 68881 72328
0 38658 7 1 2 38656 38657
0 38659 5 1 1 38658
0 38660 7 1 2 38655 38659
0 38661 5 1 1 38660
0 38662 7 1 2 78551 38661
0 38663 5 1 1 38662
0 38664 7 1 2 38640 38663
0 38665 5 1 1 38664
0 38666 7 1 2 70402 38665
0 38667 5 1 1 38666
0 38668 7 1 2 9960 70844
0 38669 5 1 1 38668
0 38670 7 2 2 63836 38669
0 38671 7 1 2 68844 78682
0 38672 5 1 1 38671
0 38673 7 1 2 71000 78675
0 38674 5 1 1 38673
0 38675 7 1 2 68590 76400
0 38676 5 3 1 38675
0 38677 7 1 2 74992 76584
0 38678 5 1 1 38677
0 38679 7 1 2 78684 38678
0 38680 7 1 2 38674 38679
0 38681 5 1 1 38680
0 38682 7 1 2 57340 38681
0 38683 5 1 1 38682
0 38684 7 1 2 70439 73356
0 38685 5 1 1 38684
0 38686 7 1 2 75340 38685
0 38687 5 1 1 38686
0 38688 7 1 2 58063 60498
0 38689 7 1 2 38687 38688
0 38690 5 1 1 38689
0 38691 7 2 2 53007 70684
0 38692 5 1 1 78687
0 38693 7 1 2 58894 78688
0 38694 5 1 1 38693
0 38695 7 1 2 58732 38694
0 38696 5 1 1 38695
0 38697 7 1 2 67532 38696
0 38698 5 1 1 38697
0 38699 7 1 2 49797 38698
0 38700 7 1 2 38690 38699
0 38701 5 1 1 38700
0 38702 7 1 2 76401 78666
0 38703 5 1 1 38702
0 38704 7 1 2 67533 72367
0 38705 5 2 1 38704
0 38706 7 1 2 53569 78689
0 38707 7 1 2 38703 38706
0 38708 5 1 1 38707
0 38709 7 1 2 57054 38708
0 38710 7 1 2 38701 38709
0 38711 5 1 1 38710
0 38712 7 4 2 50281 63837
0 38713 7 1 2 76541 78691
0 38714 5 1 1 38713
0 38715 7 1 2 78685 38714
0 38716 5 1 1 38715
0 38717 7 1 2 53394 38716
0 38718 5 1 1 38717
0 38719 7 1 2 75924 78679
0 38720 5 1 1 38719
0 38721 7 1 2 59886 76001
0 38722 5 1 1 38721
0 38723 7 1 2 50525 63838
0 38724 7 1 2 76982 38723
0 38725 7 1 2 76022 38724
0 38726 5 1 1 38725
0 38727 7 1 2 38722 38726
0 38728 7 1 2 38720 38727
0 38729 5 1 1 38728
0 38730 7 1 2 71001 38729
0 38731 5 1 1 38730
0 38732 7 1 2 38718 38731
0 38733 7 1 2 38711 38732
0 38734 7 1 2 38683 38733
0 38735 5 1 1 38734
0 38736 7 1 2 49957 38735
0 38737 5 1 1 38736
0 38738 7 1 2 38672 38737
0 38739 5 1 1 38738
0 38740 7 1 2 48960 38739
0 38741 5 1 1 38740
0 38742 7 1 2 78493 78683
0 38743 5 1 1 38742
0 38744 7 1 2 72711 78692
0 38745 5 1 1 38744
0 38746 7 1 2 38745 78686
0 38747 5 1 1 38746
0 38748 7 1 2 49958 38747
0 38749 5 1 1 38748
0 38750 7 1 2 68845 78693
0 38751 5 1 1 38750
0 38752 7 1 2 38749 38751
0 38753 5 1 1 38752
0 38754 7 1 2 48961 38753
0 38755 5 1 1 38754
0 38756 7 2 2 48818 59001
0 38757 5 1 1 78695
0 38758 7 1 2 69105 76585
0 38759 7 1 2 78696 38758
0 38760 5 1 1 38759
0 38761 7 1 2 38755 38760
0 38762 5 1 1 38761
0 38763 7 1 2 57055 38762
0 38764 5 1 1 38763
0 38765 7 1 2 76402 78514
0 38766 5 1 1 38765
0 38767 7 2 2 49798 67534
0 38768 5 2 1 78697
0 38769 7 1 2 53395 78698
0 38770 5 1 1 38769
0 38771 7 1 2 38766 38770
0 38772 5 1 1 38771
0 38773 7 1 2 57341 38772
0 38774 5 1 1 38773
0 38775 7 1 2 75244 76403
0 38776 5 1 1 38775
0 38777 7 1 2 78690 38776
0 38778 5 1 1 38777
0 38779 7 1 2 53570 38778
0 38780 5 1 1 38779
0 38781 7 1 2 53396 76404
0 38782 5 1 1 38781
0 38783 7 1 2 67537 38782
0 38784 5 1 1 38783
0 38785 7 1 2 75927 38784
0 38786 5 1 1 38785
0 38787 7 1 2 38780 38786
0 38788 7 1 2 38774 38787
0 38789 5 1 1 38788
0 38790 7 1 2 69633 38789
0 38791 5 1 1 38790
0 38792 7 1 2 38764 38791
0 38793 5 1 1 38792
0 38794 7 1 2 70647 38793
0 38795 5 1 1 38794
0 38796 7 1 2 38743 38795
0 38797 7 1 2 38741 38796
0 38798 7 1 2 38667 38797
0 38799 5 1 1 38798
0 38800 7 1 2 50849 38799
0 38801 5 1 1 38800
0 38802 7 1 2 57342 70648
0 38803 5 1 1 38802
0 38804 7 1 2 67231 38803
0 38805 5 1 1 38804
0 38806 7 1 2 64243 76678
0 38807 7 1 2 78606 38806
0 38808 7 1 2 38805 38807
0 38809 5 1 1 38808
0 38810 7 1 2 38801 38809
0 38811 5 1 1 38810
0 38812 7 1 2 55558 38811
0 38813 5 1 1 38812
0 38814 7 1 2 63790 73528
0 38815 7 1 2 78569 38814
0 38816 5 1 1 38815
0 38817 7 1 2 71259 76100
0 38818 5 1 1 38817
0 38819 7 1 2 63549 38818
0 38820 5 1 1 38819
0 38821 7 1 2 49959 76542
0 38822 5 1 1 38821
0 38823 7 1 2 68847 38822
0 38824 5 1 1 38823
0 38825 7 1 2 48962 38824
0 38826 5 1 1 38825
0 38827 7 1 2 37616 38826
0 38828 5 1 1 38827
0 38829 7 1 2 38820 38828
0 38830 5 1 1 38829
0 38831 7 1 2 77436 24334
0 38832 5 1 1 38831
0 38833 7 1 2 52706 38832
0 38834 5 1 1 38833
0 38835 7 1 2 25384 38834
0 38836 5 1 1 38835
0 38837 7 1 2 57343 69634
0 38838 7 1 2 38836 38837
0 38839 5 1 1 38838
0 38840 7 1 2 38830 38839
0 38841 5 1 1 38840
0 38842 7 1 2 55399 38841
0 38843 5 1 1 38842
0 38844 7 1 2 67736 15877
0 38845 5 1 1 38844
0 38846 7 1 2 49799 38845
0 38847 5 1 1 38846
0 38848 7 1 2 76601 78148
0 38849 5 1 1 38848
0 38850 7 1 2 38847 38849
0 38851 5 1 1 38850
0 38852 7 2 2 57056 69635
0 38853 7 1 2 51406 78701
0 38854 7 1 2 38851 38853
0 38855 5 1 1 38854
0 38856 7 1 2 38843 38855
0 38857 5 1 1 38856
0 38858 7 1 2 57660 38857
0 38859 5 1 1 38858
0 38860 7 1 2 63743 78586
0 38861 5 1 1 38860
0 38862 7 1 2 62582 77752
0 38863 5 1 1 38862
0 38864 7 1 2 78535 38863
0 38865 5 1 1 38864
0 38866 7 2 2 48819 67854
0 38867 5 1 1 78703
0 38868 7 1 2 49800 78704
0 38869 5 1 1 38868
0 38870 7 1 2 38865 38869
0 38871 5 1 1 38870
0 38872 7 1 2 56652 68400
0 38873 7 1 2 38871 38872
0 38874 5 1 1 38873
0 38875 7 1 2 38861 38874
0 38876 5 1 1 38875
0 38877 7 1 2 54785 38876
0 38878 5 1 1 38877
0 38879 7 1 2 53247 68591
0 38880 5 1 1 38879
0 38881 7 1 2 55400 24715
0 38882 5 1 1 38881
0 38883 7 1 2 52449 74417
0 38884 7 1 2 38882 38883
0 38885 5 1 1 38884
0 38886 7 1 2 38880 38885
0 38887 5 1 1 38886
0 38888 7 1 2 55947 38887
0 38889 5 1 1 38888
0 38890 7 2 2 56239 68592
0 38891 5 1 1 78705
0 38892 7 1 2 38889 38891
0 38893 5 1 1 38892
0 38894 7 1 2 58773 38893
0 38895 5 1 1 38894
0 38896 7 1 2 51407 78285
0 38897 5 1 1 38896
0 38898 7 3 2 63839 71507
0 38899 5 1 1 78707
0 38900 7 3 2 49801 66611
0 38901 5 1 1 78710
0 38902 7 1 2 56653 78711
0 38903 5 2 1 38902
0 38904 7 1 2 38899 78713
0 38905 5 1 1 38904
0 38906 7 1 2 66051 38905
0 38907 5 1 1 38906
0 38908 7 1 2 38897 38907
0 38909 7 1 2 38895 38908
0 38910 5 1 1 38909
0 38911 7 1 2 69636 38910
0 38912 5 1 1 38911
0 38913 7 1 2 38878 38912
0 38914 7 1 2 38859 38913
0 38915 5 1 1 38914
0 38916 7 1 2 55559 38915
0 38917 5 1 1 38916
0 38918 7 1 2 76031 78714
0 38919 5 1 1 38918
0 38920 7 1 2 73835 38919
0 38921 5 1 1 38920
0 38922 7 1 2 37966 38921
0 38923 5 1 1 38922
0 38924 7 1 2 49960 38923
0 38925 5 1 1 38924
0 38926 7 1 2 67621 78390
0 38927 5 1 1 38926
0 38928 7 1 2 38925 38927
0 38929 5 1 1 38928
0 38930 7 1 2 48963 38929
0 38931 5 1 1 38930
0 38932 7 1 2 63575 67902
0 38933 7 1 2 72407 75245
0 38934 7 1 2 38932 38933
0 38935 5 1 1 38934
0 38936 7 1 2 38931 38935
0 38937 5 1 1 38936
0 38938 7 1 2 66662 38937
0 38939 5 1 1 38938
0 38940 7 1 2 57661 66681
0 38941 7 1 2 74547 78149
0 38942 7 1 2 38940 38941
0 38943 5 1 1 38942
0 38944 7 1 2 38939 38943
0 38945 7 1 2 38917 38944
0 38946 5 1 1 38945
0 38947 7 1 2 60732 38946
0 38948 5 1 1 38947
0 38949 7 1 2 38816 38948
0 38950 7 1 2 38813 38949
0 38951 5 1 1 38950
0 38952 7 1 2 51984 38951
0 38953 5 1 1 38952
0 38954 7 1 2 68832 78694
0 38955 5 1 1 38954
0 38956 7 1 2 32737 38955
0 38957 5 1 1 38956
0 38958 7 1 2 48820 38957
0 38959 5 1 1 38958
0 38960 7 1 2 67344 24880
0 38961 5 1 1 38960
0 38962 7 1 2 69808 38961
0 38963 5 1 1 38962
0 38964 7 1 2 50282 78316
0 38965 5 1 1 38964
0 38966 7 1 2 62691 38965
0 38967 5 1 1 38966
0 38968 7 1 2 52707 38967
0 38969 5 1 1 38968
0 38970 7 1 2 38963 38969
0 38971 5 1 1 38970
0 38972 7 1 2 52575 38971
0 38973 5 1 1 38972
0 38974 7 2 2 69809 73529
0 38975 5 3 1 78715
0 38976 7 1 2 75994 78717
0 38977 5 1 1 38976
0 38978 7 1 2 52708 38977
0 38979 5 1 1 38978
0 38980 7 1 2 38973 38979
0 38981 5 1 1 38980
0 38982 7 1 2 49961 38981
0 38983 5 1 1 38982
0 38984 7 1 2 38959 38983
0 38985 5 1 1 38984
0 38986 7 1 2 50850 38985
0 38987 5 1 1 38986
0 38988 7 1 2 55708 78031
0 38989 7 1 2 78559 38988
0 38990 5 1 1 38989
0 38991 7 1 2 38987 38990
0 38992 5 1 1 38991
0 38993 7 1 2 50526 38992
0 38994 5 1 1 38993
0 38995 7 1 2 78019 78476
0 38996 5 1 1 38995
0 38997 7 1 2 38994 38996
0 38998 5 1 1 38997
0 38999 7 1 2 48964 38998
0 39000 5 1 1 38999
0 39001 7 1 2 63840 65773
0 39002 7 1 2 78494 39001
0 39003 5 1 1 39002
0 39004 7 1 2 39000 39003
0 39005 5 1 1 39004
0 39006 7 1 2 57057 39005
0 39007 5 1 1 39006
0 39008 7 2 2 63645 66283
0 39009 5 1 1 78720
0 39010 7 1 2 74548 78721
0 39011 5 1 1 39010
0 39012 7 2 2 63841 71045
0 39013 7 1 2 78722 78577
0 39014 5 1 1 39013
0 39015 7 1 2 39011 39014
0 39016 5 1 1 39015
0 39017 7 1 2 61357 39016
0 39018 5 1 1 39017
0 39019 7 1 2 65774 68593
0 39020 5 1 1 39019
0 39021 7 1 2 75382 78597
0 39022 7 1 2 71046 39021
0 39023 5 1 1 39022
0 39024 7 1 2 39020 39023
0 39025 5 1 1 39024
0 39026 7 1 2 53248 75834
0 39027 7 1 2 39025 39026
0 39028 5 1 1 39027
0 39029 7 1 2 51408 65775
0 39030 7 1 2 75621 39029
0 39031 5 1 1 39030
0 39032 7 1 2 39028 39031
0 39033 5 1 1 39032
0 39034 7 1 2 69637 39033
0 39035 5 1 1 39034
0 39036 7 1 2 39018 39035
0 39037 7 1 2 39007 39036
0 39038 5 1 1 39037
0 39039 7 1 2 55560 39038
0 39040 5 1 1 39039
0 39041 7 1 2 78723 78570
0 39042 5 1 1 39041
0 39043 7 1 2 64573 67048
0 39044 5 1 1 39043
0 39045 7 1 2 77983 39044
0 39046 5 1 1 39045
0 39047 7 1 2 52576 39046
0 39048 5 1 1 39047
0 39049 7 1 2 32560 39048
0 39050 5 1 1 39049
0 39051 7 1 2 78496 39050
0 39052 5 1 1 39051
0 39053 7 1 2 53571 74203
0 39054 7 1 2 77452 39053
0 39055 5 1 1 39054
0 39056 7 1 2 39052 39055
0 39057 5 1 1 39056
0 39058 7 1 2 48965 39057
0 39059 5 1 1 39058
0 39060 7 1 2 59002 67903
0 39061 7 1 2 78539 39060
0 39062 5 1 1 39061
0 39063 7 1 2 39059 39062
0 39064 5 1 1 39063
0 39065 7 1 2 55561 39064
0 39066 5 1 1 39065
0 39067 7 1 2 67742 78702
0 39068 5 1 1 39067
0 39069 7 1 2 39066 39068
0 39070 5 1 1 39069
0 39071 7 1 2 55115 39070
0 39072 5 1 1 39071
0 39073 7 1 2 75051 78287
0 39074 5 1 1 39073
0 39075 7 1 2 39072 39074
0 39076 5 1 1 39075
0 39077 7 1 2 60864 39076
0 39078 5 1 1 39077
0 39079 7 1 2 39042 39078
0 39080 7 1 2 39040 39079
0 39081 5 1 1 39080
0 39082 7 1 2 70403 39081
0 39083 5 1 1 39082
0 39084 7 1 2 63225 73788
0 39085 5 1 1 39084
0 39086 7 2 2 49962 69910
0 39087 7 2 2 65588 78724
0 39088 5 1 1 78726
0 39089 7 1 2 39085 39088
0 39090 5 1 1 39089
0 39091 7 1 2 54786 39090
0 39092 5 1 1 39091
0 39093 7 1 2 68348 71748
0 39094 5 1 1 39093
0 39095 7 1 2 39092 39094
0 39096 5 1 1 39095
0 39097 7 1 2 49802 39096
0 39098 5 1 1 39097
0 39099 7 2 2 53572 71309
0 39100 7 1 2 67268 78728
0 39101 5 1 1 39100
0 39102 7 1 2 39098 39101
0 39103 5 1 1 39102
0 39104 7 1 2 48253 39103
0 39105 5 1 1 39104
0 39106 7 1 2 56155 73641
0 39107 5 1 1 39106
0 39108 7 4 2 59326 65734
0 39109 5 1 1 78730
0 39110 7 1 2 57536 78731
0 39111 5 1 1 39110
0 39112 7 1 2 39107 39111
0 39113 5 1 1 39112
0 39114 7 1 2 67683 39113
0 39115 5 1 1 39114
0 39116 7 1 2 39105 39115
0 39117 5 1 1 39116
0 39118 7 1 2 54398 39117
0 39119 5 1 1 39118
0 39120 7 2 2 66522 71081
0 39121 5 1 1 78734
0 39122 7 1 2 67596 71867
0 39123 5 1 1 39122
0 39124 7 1 2 39121 39123
0 39125 5 1 1 39124
0 39126 7 1 2 67684 39125
0 39127 5 1 1 39126
0 39128 7 1 2 39119 39127
0 39129 5 1 1 39128
0 39130 7 1 2 47997 39129
0 39131 5 1 1 39130
0 39132 7 9 2 55562 69527
0 39133 7 2 2 49374 78736
0 39134 7 1 2 63254 78745
0 39135 5 1 1 39134
0 39136 7 1 2 15553 39135
0 39137 5 1 1 39136
0 39138 7 1 2 54787 39137
0 39139 5 1 1 39138
0 39140 7 7 2 67618 69528
0 39141 5 2 1 78747
0 39142 7 1 2 48254 73642
0 39143 5 1 1 39142
0 39144 7 1 2 78754 39143
0 39145 5 1 1 39144
0 39146 7 1 2 56156 39145
0 39147 5 1 1 39146
0 39148 7 1 2 39139 39147
0 39149 5 1 1 39148
0 39150 7 1 2 55401 39149
0 39151 5 1 1 39150
0 39152 7 1 2 58279 78727
0 39153 5 1 1 39152
0 39154 7 1 2 39151 39153
0 39155 5 1 1 39154
0 39156 7 1 2 54097 39155
0 39157 5 1 1 39156
0 39158 7 1 2 71655 71749
0 39159 5 1 1 39158
0 39160 7 1 2 39157 39159
0 39161 5 1 1 39160
0 39162 7 1 2 49803 39161
0 39163 5 1 1 39162
0 39164 7 1 2 39131 39163
0 39165 5 1 1 39164
0 39166 7 1 2 56964 39165
0 39167 5 1 1 39166
0 39168 7 1 2 72408 72525
0 39169 5 1 1 39168
0 39170 7 3 2 70477 72528
0 39171 5 3 1 78756
0 39172 7 1 2 71790 78757
0 39173 5 1 1 39172
0 39174 7 1 2 39169 39173
0 39175 5 1 1 39174
0 39176 7 1 2 73506 39175
0 39177 5 1 1 39176
0 39178 7 1 2 56157 77053
0 39179 5 1 1 39178
0 39180 7 1 2 62873 39179
0 39181 5 1 1 39180
0 39182 7 1 2 67455 71711
0 39183 7 1 2 39181 39182
0 39184 5 1 1 39183
0 39185 7 1 2 39177 39184
0 39186 5 1 1 39185
0 39187 7 1 2 60312 39186
0 39188 5 1 1 39187
0 39189 7 4 2 71664 69038
0 39190 7 1 2 60007 74427
0 39191 7 1 2 78762 39190
0 39192 5 1 1 39191
0 39193 7 1 2 39188 39192
0 39194 7 1 2 39167 39193
0 39195 5 1 1 39194
0 39196 7 1 2 58627 39195
0 39197 5 1 1 39196
0 39198 7 1 2 59552 63560
0 39199 5 1 1 39198
0 39200 7 1 2 76319 39199
0 39201 5 1 1 39200
0 39202 7 1 2 61798 39201
0 39203 5 1 1 39202
0 39204 7 1 2 62448 77103
0 39205 5 1 1 39204
0 39206 7 1 2 70404 39205
0 39207 5 1 1 39206
0 39208 7 1 2 54788 39207
0 39209 5 1 1 39208
0 39210 7 1 2 71990 39209
0 39211 5 1 1 39210
0 39212 7 1 2 51135 39211
0 39213 5 1 1 39212
0 39214 7 1 2 39203 39213
0 39215 5 1 1 39214
0 39216 7 1 2 67783 39215
0 39217 5 1 1 39216
0 39218 7 1 2 74711 78748
0 39219 5 1 1 39218
0 39220 7 1 2 67276 71868
0 39221 5 1 1 39220
0 39222 7 1 2 57836 73643
0 39223 5 1 1 39222
0 39224 7 1 2 39221 39223
0 39225 5 1 1 39224
0 39226 7 1 2 64008 39225
0 39227 5 1 1 39226
0 39228 7 1 2 58189 78746
0 39229 5 1 1 39228
0 39230 7 1 2 48255 70478
0 39231 7 2 2 72529 39230
0 39232 5 1 1 78766
0 39233 7 1 2 39229 39232
0 39234 5 1 1 39233
0 39235 7 1 2 55116 39234
0 39236 5 1 1 39235
0 39237 7 1 2 39227 39236
0 39238 5 1 1 39237
0 39239 7 1 2 61587 39238
0 39240 5 1 1 39239
0 39241 7 1 2 39219 39240
0 39242 7 1 2 39217 39241
0 39243 5 1 1 39242
0 39244 7 1 2 67685 39243
0 39245 5 1 1 39244
0 39246 7 2 2 66220 74962
0 39247 7 1 2 59271 68813
0 39248 7 1 2 78768 39247
0 39249 5 1 1 39248
0 39250 7 1 2 39245 39249
0 39251 5 1 1 39250
0 39252 7 1 2 55813 39251
0 39253 5 1 1 39252
0 39254 7 2 2 51409 78053
0 39255 7 1 2 68168 78770
0 39256 5 1 1 39255
0 39257 7 5 2 59003 73307
0 39258 5 1 1 78772
0 39259 7 1 2 65455 78773
0 39260 5 1 1 39259
0 39261 7 1 2 54399 66612
0 39262 7 2 2 78729 39261
0 39263 5 1 1 78777
0 39264 7 1 2 59456 78778
0 39265 5 1 1 39264
0 39266 7 1 2 39260 39265
0 39267 7 1 2 39256 39266
0 39268 5 1 1 39267
0 39269 7 1 2 49375 39268
0 39270 5 1 1 39269
0 39271 7 1 2 50527 66136
0 39272 5 1 1 39271
0 39273 7 1 2 47998 39272
0 39274 5 1 1 39273
0 39275 7 1 2 9806 39274
0 39276 5 1 1 39275
0 39277 7 1 2 78774 39276
0 39278 5 1 1 39277
0 39279 7 1 2 39270 39278
0 39280 5 1 1 39279
0 39281 7 1 2 48434 39280
0 39282 5 1 1 39281
0 39283 7 1 2 49252 74201
0 39284 5 1 1 39283
0 39285 7 1 2 64229 39284
0 39286 5 1 1 39285
0 39287 7 1 2 49376 39286
0 39288 5 1 1 39287
0 39289 7 1 2 65833 39288
0 39290 5 1 1 39289
0 39291 7 1 2 58313 78775
0 39292 7 1 2 39290 39291
0 39293 5 1 1 39292
0 39294 7 1 2 39282 39293
0 39295 5 1 1 39294
0 39296 7 1 2 55563 39295
0 39297 5 1 1 39296
0 39298 7 1 2 52329 61731
0 39299 5 2 1 39298
0 39300 7 1 2 58483 78779
0 39301 5 1 1 39300
0 39302 7 1 2 63915 39301
0 39303 5 1 1 39302
0 39304 7 1 2 48256 39303
0 39305 5 1 1 39304
0 39306 7 1 2 65781 77156
0 39307 5 1 1 39306
0 39308 7 1 2 58314 39307
0 39309 5 1 1 39308
0 39310 7 1 2 39305 39309
0 39311 5 1 1 39310
0 39312 7 1 2 68401 68629
0 39313 7 1 2 39311 39312
0 39314 5 1 1 39313
0 39315 7 1 2 39297 39314
0 39316 5 1 1 39315
0 39317 7 1 2 54789 39316
0 39318 5 1 1 39317
0 39319 7 1 2 48435 67322
0 39320 5 1 1 39319
0 39321 7 1 2 4734 39320
0 39322 5 1 1 39321
0 39323 7 1 2 48257 39322
0 39324 5 1 1 39323
0 39325 7 1 2 48436 65778
0 39326 5 1 1 39325
0 39327 7 1 2 39324 39326
0 39328 5 1 1 39327
0 39329 7 1 2 78749 39328
0 39330 5 1 1 39329
0 39331 7 1 2 59624 69688
0 39332 7 1 2 74527 39331
0 39333 5 1 1 39332
0 39334 7 1 2 76320 39333
0 39335 5 1 1 39334
0 39336 7 1 2 48437 39335
0 39337 5 1 1 39336
0 39338 7 1 2 49377 69428
0 39339 5 1 1 39338
0 39340 7 1 2 39337 39339
0 39341 5 1 1 39340
0 39342 7 1 2 60313 39341
0 39343 5 1 1 39342
0 39344 7 1 2 61058 63115
0 39345 5 1 1 39344
0 39346 7 1 2 57662 59464
0 39347 7 1 2 39345 39346
0 39348 5 1 1 39347
0 39349 7 1 2 69429 39348
0 39350 5 1 1 39349
0 39351 7 1 2 39343 39350
0 39352 5 1 1 39351
0 39353 7 1 2 67784 39352
0 39354 5 1 1 39353
0 39355 7 1 2 47999 78750
0 39356 5 1 1 39355
0 39357 7 2 2 69412 68956
0 39358 5 1 1 78781
0 39359 7 1 2 39356 39358
0 39360 5 2 1 39359
0 39361 7 1 2 64009 78783
0 39362 5 1 1 39361
0 39363 7 2 2 48000 78758
0 39364 5 1 1 78785
0 39365 7 1 2 67146 71692
0 39366 5 1 1 39365
0 39367 7 1 2 39364 39366
0 39368 5 1 1 39367
0 39369 7 1 2 55117 39368
0 39370 5 1 1 39369
0 39371 7 1 2 39362 39370
0 39372 5 1 1 39371
0 39373 7 1 2 60314 39372
0 39374 5 1 1 39373
0 39375 7 1 2 64162 78737
0 39376 5 1 1 39375
0 39377 7 1 2 57537 73644
0 39378 5 1 1 39377
0 39379 7 1 2 39376 39378
0 39380 5 1 1 39379
0 39381 7 1 2 63153 39380
0 39382 5 1 1 39381
0 39383 7 1 2 59553 64951
0 39384 7 1 2 78782 39383
0 39385 5 1 1 39384
0 39386 7 1 2 39382 39385
0 39387 7 1 2 39374 39386
0 39388 5 1 1 39387
0 39389 7 1 2 58628 39388
0 39390 5 1 1 39389
0 39391 7 1 2 39354 39390
0 39392 7 1 2 39330 39391
0 39393 5 1 1 39392
0 39394 7 1 2 67686 39393
0 39395 5 1 1 39394
0 39396 7 1 2 59597 71656
0 39397 7 1 2 59385 39396
0 39398 7 1 2 78769 39397
0 39399 5 1 1 39398
0 39400 7 1 2 39395 39399
0 39401 7 1 2 39318 39400
0 39402 7 1 2 39253 39401
0 39403 5 1 1 39402
0 39404 7 1 2 56412 39403
0 39405 5 1 1 39404
0 39406 7 2 2 68669 68833
0 39407 7 1 2 60271 57785
0 39408 5 1 1 39407
0 39409 7 1 2 71431 39408
0 39410 5 1 1 39409
0 39411 7 1 2 65827 39410
0 39412 5 1 1 39411
0 39413 7 1 2 55814 39412
0 39414 5 1 1 39413
0 39415 7 1 2 60315 78386
0 39416 5 1 1 39415
0 39417 7 1 2 39414 39416
0 39418 5 1 1 39417
0 39419 7 1 2 78787 39418
0 39420 5 1 1 39419
0 39421 7 1 2 39263 39420
0 39422 5 1 1 39421
0 39423 7 1 2 57538 39422
0 39424 5 1 1 39423
0 39425 7 1 2 73339 71696
0 39426 5 1 1 39425
0 39427 7 1 2 57539 78771
0 39428 5 1 1 39427
0 39429 7 1 2 39258 39428
0 39430 5 1 1 39429
0 39431 7 1 2 72783 39430
0 39432 5 1 1 39431
0 39433 7 1 2 39426 39432
0 39434 7 1 2 39424 39433
0 39435 5 1 1 39434
0 39436 7 1 2 54790 39435
0 39437 5 1 1 39436
0 39438 7 1 2 53573 66635
0 39439 7 2 2 71657 39438
0 39440 7 1 2 70866 78789
0 39441 5 1 1 39440
0 39442 7 1 2 59004 61708
0 39443 7 1 2 78027 39442
0 39444 5 1 1 39443
0 39445 7 1 2 39441 39444
0 39446 5 1 1 39445
0 39447 7 1 2 55815 39446
0 39448 5 1 1 39447
0 39449 7 2 2 66636 68814
0 39450 7 1 2 66021 78791
0 39451 5 1 1 39450
0 39452 7 1 2 39448 39451
0 39453 5 1 1 39452
0 39454 7 1 2 48001 39453
0 39455 5 1 1 39454
0 39456 7 1 2 74506 78776
0 39457 5 1 1 39456
0 39458 7 1 2 4496 78790
0 39459 5 1 1 39458
0 39460 7 1 2 39457 39459
0 39461 7 1 2 39455 39460
0 39462 7 1 2 39437 39461
0 39463 5 1 1 39462
0 39464 7 1 2 55564 39463
0 39465 5 1 1 39464
0 39466 7 1 2 48258 73984
0 39467 5 1 1 39466
0 39468 7 1 2 58702 77075
0 39469 5 1 1 39468
0 39470 7 1 2 39467 39469
0 39471 5 1 1 39470
0 39472 7 1 2 49253 39471
0 39473 5 1 1 39472
0 39474 7 1 2 63474 39473
0 39475 5 1 1 39474
0 39476 7 1 2 39475 78788
0 39477 5 1 1 39476
0 39478 7 1 2 60974 62643
0 39479 5 1 1 39478
0 39480 7 1 2 62080 76682
0 39481 7 1 2 77568 39480
0 39482 5 1 1 39481
0 39483 7 1 2 48259 62881
0 39484 7 1 2 25617 39483
0 39485 7 1 2 39482 39484
0 39486 5 1 1 39485
0 39487 7 1 2 39479 39486
0 39488 5 1 1 39487
0 39489 7 1 2 59399 78037
0 39490 7 1 2 39488 39489
0 39491 5 1 1 39490
0 39492 7 1 2 39477 39491
0 39493 5 1 1 39492
0 39494 7 1 2 55565 39493
0 39495 5 1 1 39494
0 39496 7 1 2 63890 71678
0 39497 5 1 1 39496
0 39498 7 1 2 78399 39497
0 39499 5 1 1 39498
0 39500 7 1 2 55816 39499
0 39501 5 1 1 39500
0 39502 7 1 2 63680 74388
0 39503 5 1 1 39502
0 39504 7 1 2 54400 74390
0 39505 7 1 2 39503 39504
0 39506 5 2 1 39505
0 39507 7 1 2 39501 78793
0 39508 5 1 1 39507
0 39509 7 1 2 71082 39508
0 39510 5 1 1 39509
0 39511 7 1 2 55817 78763
0 39512 5 1 1 39511
0 39513 7 1 2 39510 39512
0 39514 5 1 1 39513
0 39515 7 1 2 56773 39514
0 39516 5 1 1 39515
0 39517 7 1 2 50528 69872
0 39518 5 1 1 39517
0 39519 7 1 2 48260 39518
0 39520 5 1 1 39519
0 39521 7 1 2 71410 39520
0 39522 5 1 1 39521
0 39523 7 2 2 67785 68402
0 39524 7 1 2 73969 78795
0 39525 7 1 2 39522 39524
0 39526 5 1 1 39525
0 39527 7 1 2 39516 39526
0 39528 7 1 2 39495 39527
0 39529 5 1 1 39528
0 39530 7 1 2 56158 39529
0 39531 5 1 1 39530
0 39532 7 1 2 6783 78400
0 39533 5 1 1 39532
0 39534 7 1 2 48261 39533
0 39535 5 1 1 39534
0 39536 7 1 2 78794 39535
0 39537 5 1 1 39536
0 39538 7 1 2 71083 39537
0 39539 5 1 1 39538
0 39540 7 1 2 48262 78764
0 39541 5 1 1 39540
0 39542 7 1 2 39539 39541
0 39543 5 1 1 39542
0 39544 7 1 2 48002 39543
0 39545 5 1 1 39544
0 39546 7 1 2 65210 78765
0 39547 5 1 1 39546
0 39548 7 1 2 39545 39547
0 39549 5 1 1 39548
0 39550 7 1 2 59583 39549
0 39551 5 1 1 39550
0 39552 7 1 2 57540 67558
0 39553 7 1 2 64718 39552
0 39554 5 1 1 39553
0 39555 7 1 2 68410 39554
0 39556 5 1 1 39555
0 39557 7 1 2 56774 39556
0 39558 5 1 1 39557
0 39559 7 1 2 59272 78318
0 39560 5 1 1 39559
0 39561 7 1 2 62736 68403
0 39562 5 1 1 39561
0 39563 7 1 2 39560 39562
0 39564 7 1 2 39558 39563
0 39565 5 1 1 39564
0 39566 7 1 2 55818 39565
0 39567 5 1 1 39566
0 39568 7 1 2 63850 67538
0 39569 7 1 2 59571 39568
0 39570 7 1 2 67362 39569
0 39571 5 1 1 39570
0 39572 7 1 2 67451 78319
0 39573 5 1 1 39572
0 39574 7 1 2 62329 68404
0 39575 5 1 1 39574
0 39576 7 1 2 39573 39575
0 39577 7 1 2 39571 39576
0 39578 7 1 2 39567 39577
0 39579 5 1 1 39578
0 39580 7 1 2 54791 39579
0 39581 5 1 1 39580
0 39582 7 1 2 65008 69848
0 39583 5 1 1 39582
0 39584 7 1 2 57541 68405
0 39585 7 1 2 39583 39584
0 39586 5 1 1 39585
0 39587 7 1 2 39581 39586
0 39588 5 1 1 39587
0 39589 7 1 2 68630 39588
0 39590 5 1 1 39589
0 39591 7 1 2 49963 78439
0 39592 5 1 1 39591
0 39593 7 1 2 55402 67659
0 39594 7 1 2 78784 39593
0 39595 5 1 1 39594
0 39596 7 1 2 39592 39595
0 39597 5 1 1 39596
0 39598 7 1 2 55819 39597
0 39599 5 1 1 39598
0 39600 7 1 2 62685 74275
0 39601 5 1 1 39600
0 39602 7 1 2 39599 39601
0 39603 5 1 1 39602
0 39604 7 1 2 62416 39603
0 39605 5 1 1 39604
0 39606 7 1 2 39590 39605
0 39607 7 1 2 39551 39606
0 39608 7 1 2 39531 39607
0 39609 7 1 2 39465 39608
0 39610 5 1 1 39609
0 39611 7 1 2 56965 39610
0 39612 5 1 1 39611
0 39613 7 1 2 39405 39612
0 39614 7 1 2 39197 39613
0 39615 5 1 1 39614
0 39616 7 1 2 57965 39615
0 39617 5 1 1 39616
0 39618 7 2 2 67189 74278
0 39619 7 1 2 60954 71734
0 39620 7 1 2 78797 39619
0 39621 5 2 1 39620
0 39622 7 1 2 68080 74653
0 39623 7 1 2 78798 39622
0 39624 5 2 1 39623
0 39625 7 1 2 49254 73645
0 39626 5 1 1 39625
0 39627 7 1 2 78755 39626
0 39628 5 1 1 39627
0 39629 7 1 2 64985 39628
0 39630 5 1 1 39629
0 39631 7 1 2 67786 69430
0 39632 5 1 1 39631
0 39633 7 1 2 39630 39632
0 39634 5 1 1 39633
0 39635 7 1 2 54098 39634
0 39636 5 1 1 39635
0 39637 7 2 2 67049 72409
0 39638 5 1 1 78803
0 39639 7 1 2 78759 39638
0 39640 5 2 1 39639
0 39641 7 1 2 64664 78805
0 39642 5 1 1 39641
0 39643 7 1 2 39636 39642
0 39644 5 1 1 39643
0 39645 7 1 2 48263 39644
0 39646 5 1 1 39645
0 39647 7 1 2 57837 78732
0 39648 5 1 1 39647
0 39649 7 1 2 78760 39648
0 39650 5 1 1 39649
0 39651 7 1 2 66869 39650
0 39652 5 1 1 39651
0 39653 7 1 2 39646 39652
0 39654 5 1 1 39653
0 39655 7 1 2 55820 39654
0 39656 5 1 1 39655
0 39657 7 1 2 55566 74239
0 39658 7 1 2 78082 39657
0 39659 5 1 1 39658
0 39660 7 1 2 78761 39659
0 39661 5 1 1 39660
0 39662 7 1 2 48264 39661
0 39663 5 1 1 39662
0 39664 7 1 2 67018 66159
0 39665 7 1 2 69761 39664
0 39666 5 1 1 39665
0 39667 7 1 2 39663 39666
0 39668 5 1 1 39667
0 39669 7 1 2 54099 39668
0 39670 5 1 1 39669
0 39671 7 1 2 60975 78806
0 39672 5 1 1 39671
0 39673 7 1 2 39670 39672
0 39674 5 1 1 39673
0 39675 7 1 2 55118 39674
0 39676 5 1 1 39675
0 39677 7 1 2 65291 78735
0 39678 5 1 1 39677
0 39679 7 1 2 39676 39678
0 39680 5 1 1 39679
0 39681 7 1 2 49255 39680
0 39682 5 1 1 39681
0 39683 7 2 2 39656 39682
0 39684 7 1 2 60316 78786
0 39685 5 1 1 39684
0 39686 7 1 2 65098 78804
0 39687 5 1 1 39686
0 39688 7 1 2 39685 39687
0 39689 5 1 1 39688
0 39690 7 1 2 58629 39689
0 39691 5 1 1 39690
0 39692 7 1 2 62737 78767
0 39693 5 1 1 39692
0 39694 7 1 2 39691 39693
0 39695 5 1 1 39694
0 39696 7 2 2 55119 39695
0 39697 5 1 1 78809
0 39698 7 1 2 59048 78810
0 39699 5 1 1 39698
0 39700 7 1 2 67190 68349
0 39701 7 1 2 77706 39700
0 39702 5 1 1 39701
0 39703 7 1 2 39699 39702
0 39704 7 1 2 78807 39703
0 39705 5 1 1 39704
0 39706 7 1 2 49378 39705
0 39707 5 1 1 39706
0 39708 7 1 2 78801 39707
0 39709 5 1 1 39708
0 39710 7 1 2 48438 39709
0 39711 5 1 1 39710
0 39712 7 1 2 78799 39711
0 39713 5 1 1 39712
0 39714 7 1 2 58064 78800
0 39715 7 1 2 78802 39714
0 39716 7 1 2 39697 39715
0 39717 7 1 2 78808 39716
0 39718 5 1 1 39717
0 39719 7 1 2 63315 67687
0 39720 7 1 2 39718 39719
0 39721 7 1 2 39713 39720
0 39722 5 1 1 39721
0 39723 7 1 2 39617 39722
0 39724 5 1 1 39723
0 39725 7 1 2 48821 39724
0 39726 5 1 1 39725
0 39727 7 1 2 39083 39726
0 39728 7 1 2 38953 39727
0 39729 7 1 2 38595 39728
0 39730 7 1 2 37976 39729
0 39731 7 1 2 37579 39730
0 39732 7 1 2 35122 39731
0 39733 5 1 1 39732
0 39734 7 1 2 51771 39733
0 39735 5 1 1 39734
0 39736 7 1 2 53793 39735
0 39737 7 1 2 33289 39736
0 39738 5 1 1 39737
0 39739 7 1 2 74161 77025
0 39740 5 1 1 39739
0 39741 7 1 2 58882 73954
0 39742 5 1 1 39741
0 39743 7 1 2 57253 76759
0 39744 7 1 2 8695 39743
0 39745 5 1 1 39744
0 39746 7 1 2 61111 39745
0 39747 5 1 1 39746
0 39748 7 1 2 39742 39747
0 39749 7 1 2 39740 39748
0 39750 5 2 1 39749
0 39751 7 1 2 77098 78811
0 39752 5 1 1 39751
0 39753 7 1 2 61027 64076
0 39754 5 1 1 39753
0 39755 7 1 2 53397 39754
0 39756 5 1 1 39755
0 39757 7 1 2 61414 39756
0 39758 5 1 1 39757
0 39759 7 1 2 62141 64077
0 39760 5 1 1 39759
0 39761 7 1 2 2542 39760
0 39762 5 1 1 39761
0 39763 7 1 2 48003 39762
0 39764 5 1 1 39763
0 39765 7 3 2 62142 59625
0 39766 5 1 1 78813
0 39767 7 1 2 2811 2446
0 39768 5 1 1 39767
0 39769 7 1 2 58410 39768
0 39770 5 1 1 39769
0 39771 7 1 2 39766 39770
0 39772 7 1 2 39764 39771
0 39773 5 1 1 39772
0 39774 7 1 2 48439 39773
0 39775 5 1 1 39774
0 39776 7 1 2 39758 39775
0 39777 5 1 1 39776
0 39778 7 1 2 48559 39777
0 39779 5 1 1 39778
0 39780 7 1 2 1373 34424
0 39781 5 1 1 39780
0 39782 7 1 2 48004 39781
0 39783 5 1 1 39782
0 39784 7 1 2 61031 2546
0 39785 5 1 1 39784
0 39786 7 1 2 58411 39785
0 39787 5 1 1 39786
0 39788 7 1 2 65791 39787
0 39789 7 1 2 39783 39788
0 39790 5 1 1 39789
0 39791 7 1 2 48440 39790
0 39792 5 1 1 39791
0 39793 7 1 2 65378 59522
0 39794 7 1 2 9615 39793
0 39795 5 1 1 39794
0 39796 7 1 2 78195 39795
0 39797 7 1 2 39792 39796
0 39798 5 1 1 39797
0 39799 7 1 2 49632 39798
0 39800 5 1 1 39799
0 39801 7 1 2 39779 39800
0 39802 5 1 1 39801
0 39803 7 1 2 54100 39802
0 39804 5 1 1 39803
0 39805 7 1 2 67388 78814
0 39806 5 1 1 39805
0 39807 7 1 2 57058 78121
0 39808 5 1 1 39807
0 39809 7 1 2 54401 39808
0 39810 5 1 1 39809
0 39811 7 1 2 56159 65390
0 39812 5 1 1 39811
0 39813 7 1 2 37181 39812
0 39814 5 1 1 39813
0 39815 7 1 2 56413 39814
0 39816 5 1 1 39815
0 39817 7 1 2 39810 39816
0 39818 5 1 1 39817
0 39819 7 1 2 49633 39818
0 39820 5 1 1 39819
0 39821 7 1 2 39806 39820
0 39822 7 1 2 39804 39821
0 39823 5 1 1 39822
0 39824 7 1 2 56775 39823
0 39825 5 1 1 39824
0 39826 7 1 2 56414 65890
0 39827 5 1 1 39826
0 39828 7 2 2 57059 39827
0 39829 5 2 1 78816
0 39830 7 1 2 61824 78818
0 39831 5 1 1 39830
0 39832 7 1 2 56415 63903
0 39833 5 1 1 39832
0 39834 7 1 2 59235 75599
0 39835 5 1 1 39834
0 39836 7 1 2 71795 39835
0 39837 7 1 2 39833 39836
0 39838 5 1 1 39837
0 39839 7 1 2 54792 39838
0 39840 5 1 1 39839
0 39841 7 1 2 2548 39840
0 39842 7 1 2 39831 39841
0 39843 5 1 1 39842
0 39844 7 1 2 55821 39843
0 39845 5 1 1 39844
0 39846 7 1 2 63949 65818
0 39847 5 2 1 39846
0 39848 7 1 2 64094 78820
0 39849 5 1 1 39848
0 39850 7 1 2 49501 39849
0 39851 5 1 1 39850
0 39852 7 1 2 49256 63950
0 39853 7 1 2 66014 39852
0 39854 5 1 1 39853
0 39855 7 1 2 39851 39854
0 39856 5 1 1 39855
0 39857 7 1 2 54793 39856
0 39858 5 1 1 39857
0 39859 7 1 2 62417 62228
0 39860 5 1 1 39859
0 39861 7 1 2 53249 39860
0 39862 5 1 1 39861
0 39863 7 1 2 54794 39862
0 39864 5 1 1 39863
0 39865 7 1 2 49502 60618
0 39866 5 1 1 39865
0 39867 7 1 2 66748 39866
0 39868 5 1 1 39867
0 39869 7 1 2 54402 39868
0 39870 5 1 1 39869
0 39871 7 1 2 62695 78087
0 39872 5 1 1 39871
0 39873 7 1 2 39870 39872
0 39874 7 1 2 39864 39873
0 39875 5 1 1 39874
0 39876 7 1 2 48560 39875
0 39877 5 1 1 39876
0 39878 7 1 2 58723 62200
0 39879 5 2 1 39878
0 39880 7 1 2 62392 60991
0 39881 5 1 1 39880
0 39882 7 1 2 48561 39881
0 39883 5 1 1 39882
0 39884 7 1 2 59275 39883
0 39885 5 1 1 39884
0 39886 7 1 2 78822 39885
0 39887 5 1 1 39886
0 39888 7 1 2 39877 39887
0 39889 7 1 2 39858 39888
0 39890 7 1 2 39845 39889
0 39891 5 1 1 39890
0 39892 7 1 2 49634 39891
0 39893 5 1 1 39892
0 39894 7 1 2 71851 31665
0 39895 5 1 1 39894
0 39896 7 1 2 60976 39895
0 39897 5 1 1 39896
0 39898 7 1 2 60646 71852
0 39899 5 1 1 39898
0 39900 7 1 2 54403 76513
0 39901 7 1 2 39899 39900
0 39902 5 1 1 39901
0 39903 7 1 2 39897 39902
0 39904 5 1 1 39903
0 39905 7 1 2 48562 39904
0 39906 5 1 1 39905
0 39907 7 1 2 65151 78823
0 39908 5 1 1 39907
0 39909 7 1 2 62201 74835
0 39910 5 1 1 39909
0 39911 7 1 2 54404 77094
0 39912 7 1 2 39910 39911
0 39913 5 1 1 39912
0 39914 7 1 2 39908 39913
0 39915 5 1 1 39914
0 39916 7 1 2 49635 39915
0 39917 5 1 1 39916
0 39918 7 1 2 39906 39917
0 39919 5 1 1 39918
0 39920 7 1 2 59112 39919
0 39921 5 1 1 39920
0 39922 7 1 2 64851 61033
0 39923 5 1 1 39922
0 39924 7 1 2 55822 39923
0 39925 5 1 1 39924
0 39926 7 1 2 69391 39925
0 39927 5 1 1 39926
0 39928 7 1 2 64947 39927
0 39929 5 1 1 39928
0 39930 7 1 2 39921 39929
0 39931 7 1 2 39893 39930
0 39932 7 1 2 39825 39931
0 39933 5 1 1 39932
0 39934 7 1 2 48669 39933
0 39935 5 1 1 39934
0 39936 7 1 2 39752 39935
0 39937 5 1 1 39936
0 39938 7 1 2 77998 39937
0 39939 5 1 1 39938
0 39940 7 1 2 68838 77984
0 39941 5 6 1 39940
0 39942 7 2 2 56471 78824
0 39943 5 3 1 78830
0 39944 7 1 2 48966 78831
0 39945 5 1 1 39944
0 39946 7 1 2 56416 63872
0 39947 5 1 1 39946
0 39948 7 2 2 63898 39947
0 39949 7 1 2 67501 78835
0 39950 5 1 1 39949
0 39951 7 1 2 55823 39950
0 39952 5 1 1 39951
0 39953 7 1 2 61941 62250
0 39954 5 1 1 39953
0 39955 7 1 2 63274 66749
0 39956 5 1 1 39955
0 39957 7 1 2 74801 39956
0 39958 5 1 1 39957
0 39959 7 1 2 57542 77840
0 39960 5 1 1 39959
0 39961 7 1 2 56472 31394
0 39962 7 1 2 39960 39961
0 39963 7 1 2 39958 39962
0 39964 5 1 1 39963
0 39965 7 1 2 54405 39964
0 39966 5 1 1 39965
0 39967 7 1 2 39954 39966
0 39968 7 1 2 39952 39967
0 39969 5 1 1 39968
0 39970 7 1 2 56776 39969
0 39971 5 1 1 39970
0 39972 7 1 2 48005 62288
0 39973 5 1 1 39972
0 39974 7 1 2 77660 39973
0 39975 5 1 1 39974
0 39976 7 2 2 56160 39975
0 39977 5 1 1 78837
0 39978 7 1 2 57188 69888
0 39979 5 1 1 39978
0 39980 7 1 2 60404 74842
0 39981 5 1 1 39980
0 39982 7 1 2 39979 39981
0 39983 5 2 1 39982
0 39984 7 1 2 54795 78839
0 39985 5 1 1 39984
0 39986 7 1 2 53398 39985
0 39987 7 1 2 39977 39986
0 39988 5 1 1 39987
0 39989 7 1 2 56417 39988
0 39990 5 1 1 39989
0 39991 7 2 2 60657 77318
0 39992 7 1 2 61065 78841
0 39993 5 1 1 39992
0 39994 7 1 2 28103 39993
0 39995 5 1 1 39994
0 39996 7 1 2 57189 39995
0 39997 5 1 1 39996
0 39998 7 1 2 63912 76801
0 39999 5 1 1 39998
0 40000 7 1 2 39997 39999
0 40001 5 2 1 40000
0 40002 7 1 2 54796 78843
0 40003 5 1 1 40002
0 40004 7 1 2 48670 73300
0 40005 5 1 1 40004
0 40006 7 1 2 52709 40005
0 40007 7 1 2 40003 40006
0 40008 7 2 2 39990 40007
0 40009 5 1 1 78845
0 40010 7 1 2 56418 74314
0 40011 5 2 1 40010
0 40012 7 1 2 64976 67502
0 40013 5 1 1 40012
0 40014 7 1 2 48006 40013
0 40015 5 1 1 40014
0 40016 7 1 2 78847 40015
0 40017 5 1 1 40016
0 40018 7 1 2 61981 40017
0 40019 5 1 1 40018
0 40020 7 1 2 50283 77629
0 40021 5 1 1 40020
0 40022 7 1 2 57286 40021
0 40023 5 1 1 40022
0 40024 7 1 2 50851 40023
0 40025 5 2 1 40024
0 40026 7 1 2 57806 78849
0 40027 5 1 1 40026
0 40028 7 1 2 57077 59487
0 40029 5 1 1 40028
0 40030 7 1 2 56161 40029
0 40031 5 1 1 40030
0 40032 7 1 2 57190 62251
0 40033 5 1 1 40032
0 40034 7 1 2 40031 40033
0 40035 5 1 1 40034
0 40036 7 1 2 60250 40035
0 40037 5 1 1 40036
0 40038 7 1 2 53574 40037
0 40039 7 1 2 40027 40038
0 40040 7 1 2 40019 40039
0 40041 7 1 2 78846 40040
0 40042 7 1 2 39971 40041
0 40043 5 1 1 40042
0 40044 7 1 2 56473 67839
0 40045 5 1 1 40044
0 40046 7 1 2 78523 40045
0 40047 5 1 1 40046
0 40048 7 1 2 40043 40047
0 40049 5 1 1 40048
0 40050 7 1 2 39945 40049
0 40051 7 1 2 39939 40050
0 40052 5 1 1 40051
0 40053 7 1 2 51136 40052
0 40054 5 1 1 40053
0 40055 7 1 2 55824 70285
0 40056 5 1 1 40055
0 40057 7 1 2 70914 40056
0 40058 5 1 1 40057
0 40059 7 1 2 62583 40058
0 40060 5 1 1 40059
0 40061 7 1 2 49804 70210
0 40062 5 1 1 40061
0 40063 7 1 2 40060 40062
0 40064 5 1 1 40063
0 40065 7 1 2 52812 40064
0 40066 5 1 1 40065
0 40067 7 3 2 60221 63212
0 40068 5 1 1 78851
0 40069 7 1 2 70211 78852
0 40070 5 1 1 40069
0 40071 7 1 2 40066 40070
0 40072 5 1 1 40071
0 40073 7 1 2 56162 40072
0 40074 5 1 1 40073
0 40075 7 1 2 62584 65841
0 40076 5 1 1 40075
0 40077 7 1 2 48441 69127
0 40078 5 1 1 40077
0 40079 7 1 2 40076 40078
0 40080 5 1 1 40079
0 40081 7 1 2 52813 40080
0 40082 5 1 1 40081
0 40083 7 1 2 61394 78853
0 40084 5 1 1 40083
0 40085 7 1 2 40082 40084
0 40086 5 1 1 40085
0 40087 7 1 2 58315 40086
0 40088 5 1 1 40087
0 40089 7 1 2 54101 71697
0 40090 5 1 1 40089
0 40091 7 1 2 21077 40090
0 40092 5 1 1 40091
0 40093 7 1 2 48822 40092
0 40094 5 1 1 40093
0 40095 7 1 2 59005 78199
0 40096 5 1 1 40095
0 40097 7 1 2 40094 40096
0 40098 5 1 1 40097
0 40099 7 1 2 52330 18958
0 40100 5 1 1 40099
0 40101 7 1 2 40098 40100
0 40102 5 1 1 40101
0 40103 7 4 2 52814 62585
0 40104 7 1 2 74516 78854
0 40105 5 1 1 40104
0 40106 7 1 2 59013 40068
0 40107 5 3 1 40106
0 40108 7 1 2 50108 56654
0 40109 5 1 1 40108
0 40110 7 1 2 49379 40109
0 40111 7 1 2 78858 40110
0 40112 5 1 1 40111
0 40113 7 1 2 40105 40112
0 40114 5 1 1 40113
0 40115 7 1 2 48442 40114
0 40116 5 1 1 40115
0 40117 7 1 2 64419 61175
0 40118 5 1 1 40117
0 40119 7 1 2 68087 40118
0 40120 5 1 1 40119
0 40121 7 1 2 54406 78855
0 40122 7 1 2 40120 40121
0 40123 5 1 1 40122
0 40124 7 1 2 40116 40123
0 40125 7 1 2 40102 40124
0 40126 7 1 2 40088 40125
0 40127 7 1 2 40074 40126
0 40128 5 1 1 40127
0 40129 7 1 2 56419 40128
0 40130 5 1 1 40129
0 40131 7 1 2 48265 78859
0 40132 5 1 1 40131
0 40133 7 1 2 52815 65709
0 40134 5 1 1 40133
0 40135 7 1 2 40132 40134
0 40136 5 1 1 40135
0 40137 7 1 2 61166 40136
0 40138 5 1 1 40137
0 40139 7 1 2 65103 78856
0 40140 5 1 1 40139
0 40141 7 1 2 40138 40140
0 40142 5 1 1 40141
0 40143 7 1 2 58630 40142
0 40144 5 1 1 40143
0 40145 7 1 2 57543 78857
0 40146 7 1 2 77123 40145
0 40147 5 1 1 40146
0 40148 7 1 2 40144 40147
0 40149 7 1 2 40130 40148
0 40150 5 1 1 40149
0 40151 7 1 2 56589 40150
0 40152 5 1 1 40151
0 40153 7 1 2 65795 74576
0 40154 5 1 1 40153
0 40155 7 1 2 77121 40154
0 40156 5 1 1 40155
0 40157 7 1 2 61233 71693
0 40158 7 1 2 40156 40157
0 40159 5 1 1 40158
0 40160 7 1 2 40152 40159
0 40161 5 1 1 40160
0 40162 7 1 2 53724 40161
0 40163 5 1 1 40162
0 40164 7 1 2 63695 67840
0 40165 5 1 1 40164
0 40166 7 1 2 63316 78860
0 40167 5 1 1 40166
0 40168 7 1 2 48967 63696
0 40169 5 1 1 40168
0 40170 7 1 2 38757 40169
0 40171 7 1 2 40167 40170
0 40172 5 1 1 40171
0 40173 7 1 2 53725 40172
0 40174 5 1 1 40173
0 40175 7 1 2 40165 40174
0 40176 5 1 1 40175
0 40177 7 1 2 77110 40176
0 40178 5 1 1 40177
0 40179 7 1 2 52710 70578
0 40180 5 4 1 40179
0 40181 7 1 2 62981 65593
0 40182 5 1 1 40181
0 40183 7 1 2 62586 69529
0 40184 7 1 2 40182 40183
0 40185 5 1 1 40184
0 40186 7 1 2 78861 40185
0 40187 5 1 1 40186
0 40188 7 1 2 60251 40187
0 40189 5 1 1 40188
0 40190 7 1 2 67121 71459
0 40191 5 1 1 40190
0 40192 7 1 2 74932 40191
0 40193 5 8 1 40192
0 40194 7 1 2 60252 70195
0 40195 5 1 1 40194
0 40196 7 1 2 54102 71427
0 40197 5 1 1 40196
0 40198 7 1 2 57663 76675
0 40199 5 1 1 40198
0 40200 7 1 2 40197 40199
0 40201 7 1 2 40195 40200
0 40202 5 1 1 40201
0 40203 7 1 2 78865 40202
0 40204 5 1 1 40203
0 40205 7 1 2 40189 40204
0 40206 7 1 2 40178 40205
0 40207 7 1 2 40163 40206
0 40208 5 1 1 40207
0 40209 7 1 2 55120 40208
0 40210 5 1 1 40209
0 40211 7 1 2 48266 77016
0 40212 5 1 1 40211
0 40213 7 1 2 66834 40212
0 40214 5 1 1 40213
0 40215 7 1 2 59065 40214
0 40216 5 1 1 40215
0 40217 7 1 2 58273 30146
0 40218 5 1 1 40217
0 40219 7 1 2 61368 40218
0 40220 5 1 1 40219
0 40221 7 1 2 62816 68045
0 40222 5 1 1 40221
0 40223 7 1 2 40220 40222
0 40224 7 1 2 40216 40223
0 40225 5 1 1 40224
0 40226 7 1 2 55825 40225
0 40227 5 1 1 40226
0 40228 7 1 2 61410 61990
0 40229 5 1 1 40228
0 40230 7 1 2 59066 74218
0 40231 5 1 1 40230
0 40232 7 1 2 65379 61369
0 40233 5 1 1 40232
0 40234 7 1 2 40231 40233
0 40235 5 1 1 40234
0 40236 7 1 2 61843 40235
0 40237 5 1 1 40236
0 40238 7 1 2 54103 61483
0 40239 7 1 2 59067 40238
0 40240 5 1 1 40239
0 40241 7 1 2 61361 40240
0 40242 5 1 1 40241
0 40243 7 1 2 61066 40242
0 40244 5 1 1 40243
0 40245 7 1 2 59280 63878
0 40246 5 1 1 40245
0 40247 7 1 2 61861 68200
0 40248 5 1 1 40247
0 40249 7 1 2 68037 40248
0 40250 7 1 2 40246 40249
0 40251 7 1 2 40244 40250
0 40252 7 1 2 40237 40251
0 40253 7 1 2 40229 40252
0 40254 7 1 2 40227 40253
0 40255 5 1 1 40254
0 40256 7 1 2 74242 40255
0 40257 5 1 1 40256
0 40258 7 1 2 40210 40257
0 40259 5 1 1 40258
0 40260 7 1 2 54797 40259
0 40261 5 1 1 40260
0 40262 7 1 2 73326 74257
0 40263 5 7 1 40262
0 40264 7 2 2 56420 78873
0 40265 5 1 1 78880
0 40266 7 1 2 56590 67855
0 40267 5 2 1 40266
0 40268 7 1 2 40265 78882
0 40269 5 1 1 40268
0 40270 7 1 2 55121 40269
0 40271 5 1 1 40270
0 40272 7 1 2 69638 71508
0 40273 5 1 1 40272
0 40274 7 1 2 53575 38867
0 40275 7 1 2 40273 40274
0 40276 7 1 2 40271 40275
0 40277 5 1 1 40276
0 40278 7 3 2 58774 67856
0 40279 5 1 1 78884
0 40280 7 1 2 49805 40279
0 40281 5 1 1 40280
0 40282 7 1 2 60222 40281
0 40283 7 1 2 40277 40282
0 40284 5 1 1 40283
0 40285 7 1 2 57838 68028
0 40286 5 1 1 40285
0 40287 7 1 2 7135 40286
0 40288 5 1 1 40287
0 40289 7 1 2 55122 40288
0 40290 5 1 1 40289
0 40291 7 1 2 58775 78817
0 40292 5 1 1 40291
0 40293 7 1 2 54104 58124
0 40294 7 1 2 40292 40293
0 40295 5 1 1 40294
0 40296 7 1 2 40290 40295
0 40297 5 1 1 40296
0 40298 7 1 2 55826 40297
0 40299 5 1 1 40298
0 40300 7 1 2 58585 77010
0 40301 7 1 2 78780 40300
0 40302 5 1 1 40301
0 40303 7 1 2 57060 58776
0 40304 7 1 2 40302 40303
0 40305 5 1 1 40304
0 40306 7 1 2 58125 40305
0 40307 5 1 1 40306
0 40308 7 1 2 7931 40307
0 40309 5 1 1 40308
0 40310 7 1 2 52711 65594
0 40311 5 1 1 40310
0 40312 7 1 2 54407 40311
0 40313 7 1 2 40309 40312
0 40314 5 1 1 40313
0 40315 7 1 2 40299 40314
0 40316 5 1 1 40315
0 40317 7 1 2 56777 40316
0 40318 5 1 1 40317
0 40319 7 1 2 65099 58139
0 40320 5 1 1 40319
0 40321 7 1 2 77105 40320
0 40322 5 1 1 40321
0 40323 7 1 2 49137 40322
0 40324 5 1 1 40323
0 40325 7 1 2 56163 72895
0 40326 5 1 1 40325
0 40327 7 1 2 57664 40326
0 40328 7 2 2 40324 40327
0 40329 5 1 1 78887
0 40330 7 1 2 67970 78888
0 40331 5 1 1 40330
0 40332 7 1 2 67248 40331
0 40333 5 1 1 40332
0 40334 7 1 2 48671 67257
0 40335 7 1 2 40329 40334
0 40336 5 1 1 40335
0 40337 7 1 2 40333 40336
0 40338 5 1 1 40337
0 40339 7 1 2 55123 40338
0 40340 5 1 1 40339
0 40341 7 1 2 60253 67627
0 40342 5 1 1 40341
0 40343 7 1 2 48823 71120
0 40344 5 2 1 40343
0 40345 7 1 2 64200 70200
0 40346 5 1 1 40345
0 40347 7 1 2 59592 74637
0 40348 5 1 1 40347
0 40349 7 1 2 40346 40348
0 40350 5 1 1 40349
0 40351 7 1 2 59724 40350
0 40352 5 1 1 40351
0 40353 7 1 2 78889 40352
0 40354 5 1 1 40353
0 40355 7 1 2 56421 40354
0 40356 5 1 1 40355
0 40357 7 1 2 40342 40356
0 40358 7 1 2 40340 40357
0 40359 7 1 2 58946 74231
0 40360 5 1 1 40359
0 40361 7 1 2 66663 40360
0 40362 5 1 1 40361
0 40363 7 1 2 55124 40362
0 40364 5 1 1 40363
0 40365 7 1 2 19591 40364
0 40366 5 1 1 40365
0 40367 7 1 2 56591 40366
0 40368 5 1 1 40367
0 40369 7 1 2 55827 64512
0 40370 5 1 1 40369
0 40371 7 1 2 58929 40370
0 40372 5 1 1 40371
0 40373 7 1 2 54105 40372
0 40374 5 1 1 40373
0 40375 7 1 2 64524 40374
0 40376 5 1 1 40375
0 40377 7 1 2 58126 40376
0 40378 5 1 1 40377
0 40379 7 1 2 40368 40378
0 40380 5 1 1 40379
0 40381 7 1 2 57287 40380
0 40382 5 1 1 40381
0 40383 7 1 2 65155 69889
0 40384 5 1 1 40383
0 40385 7 1 2 58930 40384
0 40386 5 1 1 40385
0 40387 7 1 2 68911 40386
0 40388 5 1 1 40387
0 40389 7 1 2 48824 60658
0 40390 5 1 1 40389
0 40391 7 1 2 40388 40390
0 40392 5 1 1 40391
0 40393 7 1 2 56592 40392
0 40394 5 1 1 40393
0 40395 7 1 2 68155 77364
0 40396 5 1 1 40395
0 40397 7 1 2 77771 40396
0 40398 5 1 1 40397
0 40399 7 1 2 56422 40398
0 40400 5 1 1 40399
0 40401 7 1 2 56966 60659
0 40402 5 1 1 40401
0 40403 7 1 2 68913 40402
0 40404 7 1 2 40400 40403
0 40405 5 1 1 40404
0 40406 7 1 2 58127 40405
0 40407 5 1 1 40406
0 40408 7 1 2 40394 40407
0 40409 5 1 1 40408
0 40410 7 1 2 54408 40409
0 40411 5 1 1 40410
0 40412 7 1 2 40382 40411
0 40413 7 1 2 40358 40412
0 40414 7 1 2 49636 63226
0 40415 5 1 1 40414
0 40416 7 1 2 3806 40415
0 40417 5 1 1 40416
0 40418 7 1 2 48007 40417
0 40419 5 1 1 40418
0 40420 7 1 2 5958 40419
0 40421 5 1 1 40420
0 40422 7 1 2 59725 40421
0 40423 5 1 1 40422
0 40424 7 1 2 52712 64204
0 40425 7 1 2 40423 40424
0 40426 5 1 1 40425
0 40427 7 1 2 56423 40426
0 40428 5 1 1 40427
0 40429 7 1 2 78890 40428
0 40430 5 1 1 40429
0 40431 7 1 2 48672 40430
0 40432 5 1 1 40431
0 40433 7 2 2 58557 77069
0 40434 5 1 1 78891
0 40435 7 1 2 54106 64897
0 40436 5 1 1 40435
0 40437 7 1 2 40434 40436
0 40438 5 1 1 40437
0 40439 7 1 2 55125 40438
0 40440 5 1 1 40439
0 40441 7 1 2 48008 74638
0 40442 5 1 1 40441
0 40443 7 1 2 40440 40442
0 40444 5 1 1 40443
0 40445 7 1 2 56593 40444
0 40446 5 1 1 40445
0 40447 7 1 2 55126 61141
0 40448 5 1 1 40447
0 40449 7 1 2 34873 40448
0 40450 5 1 1 40449
0 40451 7 1 2 54107 40450
0 40452 5 1 1 40451
0 40453 7 1 2 48009 64520
0 40454 5 1 1 40453
0 40455 7 1 2 40452 40454
0 40456 5 1 1 40455
0 40457 7 1 2 58128 40456
0 40458 5 1 1 40457
0 40459 7 1 2 40446 40458
0 40460 5 1 1 40459
0 40461 7 1 2 61982 40460
0 40462 5 1 1 40461
0 40463 7 1 2 40432 40462
0 40464 7 1 2 40413 40463
0 40465 7 1 2 40318 40464
0 40466 5 1 1 40465
0 40467 7 1 2 69039 40466
0 40468 5 1 1 40467
0 40469 7 1 2 40284 40468
0 40470 7 2 2 40261 40469
0 40471 5 1 1 78893
0 40472 7 1 2 40054 78894
0 40473 5 1 1 40472
0 40474 7 1 2 51772 40473
0 40475 5 1 1 40474
0 40476 7 1 2 71509 69018
0 40477 5 1 1 40476
0 40478 7 1 2 7951 40477
0 40479 5 1 1 40478
0 40480 7 1 2 52816 40479
0 40481 5 1 1 40480
0 40482 7 8 2 61221 70481
0 40483 7 1 2 49964 78895
0 40484 5 2 1 40483
0 40485 7 1 2 49806 67122
0 40486 5 1 1 40485
0 40487 7 1 2 78903 40486
0 40488 5 3 1 40487
0 40489 7 1 2 51773 78905
0 40490 5 1 1 40489
0 40491 7 1 2 40481 40490
0 40492 5 5 1 40491
0 40493 7 1 2 56424 60811
0 40494 5 3 1 40493
0 40495 7 1 2 56240 63916
0 40496 5 1 1 40495
0 40497 7 1 2 49380 40496
0 40498 5 1 1 40497
0 40499 7 2 2 78913 40498
0 40500 7 1 2 51137 78916
0 40501 7 1 2 78908 40500
0 40502 5 1 1 40501
0 40503 7 1 2 40475 40502
0 40504 5 1 1 40503
0 40505 7 1 2 51631 40504
0 40506 5 1 1 40505
0 40507 7 2 2 60178 60767
0 40508 7 3 2 71432 78918
0 40509 5 1 1 78920
0 40510 7 2 2 60437 78921
0 40511 5 2 1 78923
0 40512 7 2 2 75898 78925
0 40513 5 1 1 78927
0 40514 7 1 2 48968 78928
0 40515 5 1 1 40514
0 40516 7 2 2 51138 78896
0 40517 7 1 2 51985 70261
0 40518 5 1 1 40517
0 40519 7 1 2 65449 40518
0 40520 5 1 1 40519
0 40521 7 1 2 55709 40520
0 40522 5 1 1 40521
0 40523 7 1 2 35001 40522
0 40524 5 1 1 40523
0 40525 7 1 2 52331 40524
0 40526 5 1 1 40525
0 40527 7 2 2 61532 59662
0 40528 5 1 1 78931
0 40529 7 1 2 55710 78932
0 40530 5 1 1 40529
0 40531 7 1 2 40526 40530
0 40532 5 1 1 40531
0 40533 7 1 2 52185 40532
0 40534 5 1 1 40533
0 40535 7 1 2 59663 59818
0 40536 7 1 2 72695 40535
0 40537 5 1 1 40536
0 40538 7 1 2 40534 40537
0 40539 5 2 1 40538
0 40540 7 1 2 78929 78933
0 40541 5 1 1 40540
0 40542 7 1 2 40515 40541
0 40543 5 1 1 40542
0 40544 7 1 2 56241 40543
0 40545 5 1 1 40544
0 40546 7 4 2 67961 73831
0 40547 5 2 1 78935
0 40548 7 1 2 70685 78936
0 40549 5 1 1 40548
0 40550 7 1 2 40545 40549
0 40551 5 1 1 40550
0 40552 7 1 2 53726 40551
0 40553 5 1 1 40552
0 40554 7 1 2 49637 29962
0 40555 5 1 1 40554
0 40556 7 1 2 61293 67232
0 40557 5 1 1 40556
0 40558 7 1 2 40555 40557
0 40559 5 1 1 40558
0 40560 7 1 2 56164 40559
0 40561 5 1 1 40560
0 40562 7 1 2 74779 77554
0 40563 5 1 1 40562
0 40564 7 1 2 57112 40563
0 40565 5 1 1 40564
0 40566 7 1 2 55711 71024
0 40567 5 1 1 40566
0 40568 7 1 2 48673 40567
0 40569 5 1 1 40568
0 40570 7 1 2 78470 35106
0 40571 7 1 2 40569 40570
0 40572 5 1 1 40571
0 40573 7 1 2 56425 40572
0 40574 5 1 1 40573
0 40575 7 1 2 40565 40574
0 40576 7 1 2 40561 40575
0 40577 5 1 1 40576
0 40578 7 1 2 51139 40577
0 40579 5 1 1 40578
0 40580 7 1 2 63227 78259
0 40581 5 1 1 40580
0 40582 7 1 2 59236 76392
0 40583 5 1 1 40582
0 40584 7 1 2 40581 40583
0 40585 5 1 1 40584
0 40586 7 1 2 76056 40585
0 40587 5 1 1 40586
0 40588 7 1 2 77453 78162
0 40589 5 1 1 40588
0 40590 7 1 2 76393 77560
0 40591 5 1 1 40590
0 40592 7 1 2 40589 40591
0 40593 7 1 2 40587 40592
0 40594 7 1 2 40579 40593
0 40595 5 1 1 40594
0 40596 7 1 2 50529 40595
0 40597 5 1 1 40596
0 40598 7 1 2 71115 75656
0 40599 5 1 1 40598
0 40600 7 1 2 75512 40599
0 40601 5 1 1 40600
0 40602 7 1 2 64848 40601
0 40603 5 1 1 40602
0 40604 7 1 2 24253 77939
0 40605 5 1 1 40604
0 40606 7 1 2 59887 40605
0 40607 5 1 1 40606
0 40608 7 1 2 40603 40607
0 40609 5 1 1 40608
0 40610 7 1 2 55828 40609
0 40611 5 1 1 40610
0 40612 7 1 2 52713 71847
0 40613 5 2 1 40612
0 40614 7 3 2 51140 57113
0 40615 7 1 2 73460 71853
0 40616 7 1 2 78943 40615
0 40617 5 1 1 40616
0 40618 7 1 2 78941 40617
0 40619 5 1 1 40618
0 40620 7 1 2 56165 40619
0 40621 5 1 1 40620
0 40622 7 1 2 51141 78460
0 40623 7 1 2 57807 40622
0 40624 5 1 1 40623
0 40625 7 1 2 78942 40624
0 40626 5 1 1 40625
0 40627 7 1 2 74586 40626
0 40628 5 1 1 40627
0 40629 7 1 2 77080 78944
0 40630 5 1 1 40629
0 40631 7 1 2 78142 40630
0 40632 7 1 2 40628 40631
0 40633 7 1 2 40621 40632
0 40634 7 1 2 40611 40633
0 40635 5 1 1 40634
0 40636 7 1 2 54409 40635
0 40637 5 1 1 40636
0 40638 7 1 2 50284 57344
0 40639 5 1 1 40638
0 40640 7 1 2 70873 40639
0 40641 5 1 1 40640
0 40642 7 1 2 77462 40641
0 40643 5 1 1 40642
0 40644 7 1 2 62034 77149
0 40645 5 1 1 40644
0 40646 7 1 2 54108 40645
0 40647 5 1 1 40646
0 40648 7 1 2 77672 40647
0 40649 5 1 1 40648
0 40650 7 1 2 69890 40649
0 40651 5 1 1 40650
0 40652 7 1 2 56778 77676
0 40653 5 1 1 40652
0 40654 7 1 2 56166 75749
0 40655 5 1 1 40654
0 40656 7 1 2 52577 40655
0 40657 7 1 2 63043 40656
0 40658 7 1 2 40653 40657
0 40659 7 1 2 40651 40658
0 40660 5 1 1 40659
0 40661 7 1 2 52714 40660
0 40662 5 1 1 40661
0 40663 7 1 2 40643 40662
0 40664 5 1 1 40663
0 40665 7 1 2 55127 40664
0 40666 5 1 1 40665
0 40667 7 1 2 40637 40666
0 40668 7 1 2 40597 40667
0 40669 5 1 1 40668
0 40670 7 1 2 54798 40669
0 40671 5 1 1 40670
0 40672 7 1 2 48674 63139
0 40673 7 1 2 603 40672
0 40674 5 1 1 40673
0 40675 7 1 2 64205 40674
0 40676 5 1 1 40675
0 40677 7 1 2 71225 70752
0 40678 5 1 1 40677
0 40679 7 1 2 40676 40678
0 40680 5 1 1 40679
0 40681 7 1 2 48825 40680
0 40682 5 1 1 40681
0 40683 7 1 2 69873 77353
0 40684 5 1 1 40683
0 40685 7 1 2 55128 40684
0 40686 5 1 1 40685
0 40687 7 1 2 52578 40686
0 40688 5 1 1 40687
0 40689 7 1 2 75505 40688
0 40690 5 1 1 40689
0 40691 7 1 2 50530 56594
0 40692 7 1 2 67562 40691
0 40693 5 1 1 40692
0 40694 7 1 2 40690 40693
0 40695 7 1 2 40682 40694
0 40696 7 1 2 40671 40695
0 40697 5 1 1 40696
0 40698 7 1 2 53576 40697
0 40699 5 1 1 40698
0 40700 7 1 2 29528 78556
0 40701 5 1 1 40700
0 40702 7 1 2 52579 40701
0 40703 5 1 1 40702
0 40704 7 1 2 56242 78561
0 40705 5 1 1 40704
0 40706 7 1 2 40703 40705
0 40707 5 1 1 40706
0 40708 7 1 2 78926 40707
0 40709 5 1 1 40708
0 40710 7 1 2 62686 77354
0 40711 5 1 1 40710
0 40712 7 1 2 76007 40711
0 40713 5 1 1 40712
0 40714 7 1 2 51986 40713
0 40715 5 1 1 40714
0 40716 7 1 2 71205 75855
0 40717 7 1 2 75355 40716
0 40718 5 1 1 40717
0 40719 7 1 2 76008 40718
0 40720 5 1 1 40719
0 40721 7 1 2 57665 40720
0 40722 5 1 1 40721
0 40723 7 1 2 40715 40722
0 40724 5 1 1 40723
0 40725 7 1 2 50531 40724
0 40726 5 1 1 40725
0 40727 7 4 2 76863 75811
0 40728 5 1 1 78946
0 40729 7 1 2 55712 62687
0 40730 7 1 2 78947 40729
0 40731 5 1 1 40730
0 40732 7 1 2 76009 40731
0 40733 5 1 1 40732
0 40734 7 1 2 73036 40733
0 40735 5 1 1 40734
0 40736 7 1 2 70690 71526
0 40737 5 1 1 40736
0 40738 7 1 2 70327 40737
0 40739 5 1 1 40738
0 40740 7 1 2 53727 40739
0 40741 7 1 2 40735 40740
0 40742 7 1 2 40726 40741
0 40743 7 1 2 40709 40742
0 40744 7 1 2 40699 40743
0 40745 5 1 1 40744
0 40746 7 5 2 51142 72712
0 40747 7 1 2 78950 78934
0 40748 5 1 1 40747
0 40749 7 1 2 40513 40748
0 40750 5 1 1 40749
0 40751 7 1 2 56243 40750
0 40752 5 1 1 40751
0 40753 7 1 2 59358 75064
0 40754 5 1 1 40753
0 40755 7 1 2 49965 40754
0 40756 7 1 2 40752 40755
0 40757 5 1 1 40756
0 40758 7 1 2 52817 40757
0 40759 7 1 2 40745 40758
0 40760 5 1 1 40759
0 40761 7 1 2 40553 40760
0 40762 5 1 1 40761
0 40763 7 2 2 67952 40762
0 40764 5 1 1 78955
0 40765 7 1 2 65735 78937
0 40766 5 1 1 40765
0 40767 7 1 2 53728 61439
0 40768 5 1 1 40767
0 40769 7 1 2 78832 40768
0 40770 5 1 1 40769
0 40771 7 2 2 52818 40770
0 40772 5 1 1 78957
0 40773 7 1 2 55567 78958
0 40774 5 1 1 40773
0 40775 7 1 2 40766 40774
0 40776 5 1 1 40775
0 40777 7 1 2 51774 40776
0 40778 5 1 1 40777
0 40779 7 1 2 50532 51632
0 40780 7 1 2 70456 40779
0 40781 7 1 2 78909 40780
0 40782 5 1 1 40781
0 40783 7 1 2 40778 40782
0 40784 5 1 1 40783
0 40785 7 1 2 63917 70778
0 40786 7 1 2 40784 40785
0 40787 5 1 1 40786
0 40788 7 1 2 40764 40787
0 40789 7 1 2 40506 40788
0 40790 5 1 1 40789
0 40791 7 1 2 51410 40790
0 40792 5 1 1 40791
0 40793 7 1 2 53008 62380
0 40794 5 1 1 40793
0 40795 7 1 2 66206 40794
0 40796 5 1 1 40795
0 40797 7 1 2 55948 40796
0 40798 5 1 1 40797
0 40799 7 1 2 9755 40798
0 40800 5 1 1 40799
0 40801 7 1 2 59945 40800
0 40802 5 1 1 40801
0 40803 7 1 2 53009 77897
0 40804 5 1 1 40803
0 40805 7 1 2 40802 40804
0 40806 5 1 1 40805
0 40807 7 1 2 50533 40806
0 40808 5 1 1 40807
0 40809 7 1 2 51987 78617
0 40810 5 2 1 40809
0 40811 7 1 2 40808 78959
0 40812 5 1 1 40811
0 40813 7 1 2 55403 40812
0 40814 5 1 1 40813
0 40815 7 2 2 63744 74073
0 40816 5 1 1 78961
0 40817 7 1 2 70257 78962
0 40818 5 1 1 40817
0 40819 7 1 2 66664 73181
0 40820 5 1 1 40819
0 40821 7 1 2 65345 67405
0 40822 5 1 1 40821
0 40823 7 1 2 40820 40822
0 40824 5 1 1 40823
0 40825 7 1 2 68406 40824
0 40826 5 1 1 40825
0 40827 7 1 2 63184 71386
0 40828 5 1 1 40827
0 40829 7 4 2 65939 70869
0 40830 5 1 1 78963
0 40831 7 1 2 63791 78964
0 40832 5 1 1 40831
0 40833 7 1 2 55129 77918
0 40834 5 1 1 40833
0 40835 7 1 2 40832 40834
0 40836 5 1 1 40835
0 40837 7 1 2 51988 40836
0 40838 5 1 1 40837
0 40839 7 1 2 40828 40838
0 40840 7 1 2 40826 40839
0 40841 5 1 1 40840
0 40842 7 1 2 52186 40841
0 40843 5 1 1 40842
0 40844 7 1 2 40818 40843
0 40845 7 1 2 40814 40844
0 40846 5 1 1 40845
0 40847 7 1 2 78866 40846
0 40848 5 1 1 40847
0 40849 7 1 2 67878 78904
0 40850 5 5 1 40849
0 40851 7 3 2 51411 78967
0 40852 7 1 2 57254 78612
0 40853 5 1 1 40852
0 40854 7 1 2 70870 72745
0 40855 5 1 1 40854
0 40856 7 1 2 59163 40855
0 40857 5 1 1 40856
0 40858 7 1 2 56655 40857
0 40859 5 1 1 40858
0 40860 7 1 2 57061 78624
0 40861 5 1 1 40860
0 40862 7 1 2 62384 38157
0 40863 5 2 1 40862
0 40864 7 1 2 55949 78975
0 40865 5 1 1 40864
0 40866 7 1 2 40861 40865
0 40867 7 1 2 40859 40866
0 40868 5 1 1 40867
0 40869 7 1 2 50285 40868
0 40870 5 1 1 40869
0 40871 7 1 2 65363 61687
0 40872 5 1 1 40871
0 40873 7 1 2 57062 40872
0 40874 5 1 1 40873
0 40875 7 3 2 51989 56244
0 40876 5 1 1 78977
0 40877 7 1 2 61300 56656
0 40878 5 1 1 40877
0 40879 7 1 2 40876 40878
0 40880 7 1 2 40874 40879
0 40881 5 1 1 40880
0 40882 7 1 2 51143 40881
0 40883 5 1 1 40882
0 40884 7 1 2 40870 40883
0 40885 7 1 2 40853 40884
0 40886 5 1 1 40885
0 40887 7 1 2 78972 40886
0 40888 5 1 1 40887
0 40889 7 2 2 64574 71869
0 40890 5 2 1 78980
0 40891 7 3 2 72702 78885
0 40892 5 1 1 78984
0 40893 7 1 2 78982 40892
0 40894 5 4 1 40893
0 40895 7 3 2 55404 78987
0 40896 5 1 1 78991
0 40897 7 3 2 50286 66665
0 40898 5 1 1 78994
0 40899 7 1 2 61510 40898
0 40900 5 1 1 40899
0 40901 7 1 2 57255 40900
0 40902 5 1 1 40901
0 40903 7 1 2 66666 73001
0 40904 5 1 1 40903
0 40905 7 1 2 38387 40904
0 40906 7 1 2 40902 40905
0 40907 5 1 1 40906
0 40908 7 1 2 78992 40907
0 40909 5 1 1 40908
0 40910 7 1 2 40888 40909
0 40911 7 1 2 40848 40910
0 40912 5 1 1 40911
0 40913 7 1 2 51633 40912
0 40914 5 1 1 40913
0 40915 7 1 2 68407 68315
0 40916 5 2 1 40915
0 40917 7 1 2 52187 75158
0 40918 7 1 2 73633 40917
0 40919 5 1 1 40918
0 40920 7 1 2 78997 40919
0 40921 5 1 1 40920
0 40922 7 1 2 58777 40921
0 40923 5 1 1 40922
0 40924 7 2 2 70595 76474
0 40925 5 1 1 78999
0 40926 7 2 2 51412 64201
0 40927 7 1 2 61694 63663
0 40928 7 1 2 79001 40927
0 40929 5 1 1 40928
0 40930 7 1 2 40925 40929
0 40931 5 1 1 40930
0 40932 7 1 2 54799 40931
0 40933 5 1 1 40932
0 40934 7 1 2 40923 40933
0 40935 5 1 1 40934
0 40936 7 1 2 51990 40935
0 40937 5 1 1 40936
0 40938 7 1 2 52580 67339
0 40939 5 3 1 40938
0 40940 7 1 2 73530 73804
0 40941 5 1 1 40940
0 40942 7 1 2 79003 40941
0 40943 5 1 1 40942
0 40944 7 1 2 55405 40943
0 40945 5 1 1 40944
0 40946 7 1 2 75641 40945
0 40947 5 1 1 40946
0 40948 7 1 2 50534 40947
0 40949 5 1 1 40948
0 40950 7 1 2 75347 78320
0 40951 5 1 1 40950
0 40952 7 1 2 40949 40951
0 40953 5 1 1 40952
0 40954 7 1 2 57256 40953
0 40955 5 1 1 40954
0 40956 7 2 2 63704 78667
0 40957 5 1 1 79006
0 40958 7 1 2 64177 63745
0 40959 5 2 1 40958
0 40960 7 1 2 40957 79008
0 40961 5 1 1 40960
0 40962 7 1 2 50287 40961
0 40963 5 1 1 40962
0 40964 7 1 2 40955 40963
0 40965 5 1 1 40964
0 40966 7 1 2 53577 40965
0 40967 5 1 1 40966
0 40968 7 2 2 51413 70328
0 40969 5 3 1 79010
0 40970 7 1 2 50288 79011
0 40971 5 1 1 40970
0 40972 7 2 2 73531 75109
0 40973 7 1 2 73871 79015
0 40974 5 1 1 40973
0 40975 7 1 2 79012 40974
0 40976 5 2 1 40975
0 40977 7 1 2 61603 79017
0 40978 5 1 1 40977
0 40979 7 1 2 40971 40978
0 40980 7 1 2 40967 40979
0 40981 5 1 1 40980
0 40982 7 1 2 50852 40981
0 40983 5 1 1 40982
0 40984 7 1 2 40937 40983
0 40985 5 1 1 40984
0 40986 7 1 2 53729 40985
0 40987 5 1 1 40986
0 40988 7 2 2 56474 77960
0 40989 7 1 2 73468 79019
0 40990 5 1 1 40989
0 40991 7 1 2 40987 40990
0 40992 5 1 1 40991
0 40993 7 1 2 66667 40992
0 40994 5 1 1 40993
0 40995 7 1 2 76363 78581
0 40996 5 2 1 40995
0 40997 7 1 2 78660 79021
0 40998 5 1 1 40997
0 40999 7 1 2 53578 40998
0 41000 5 1 1 40999
0 41001 7 1 2 6061 73758
0 41002 5 2 1 41001
0 41003 7 1 2 70329 79023
0 41004 5 1 1 41003
0 41005 7 1 2 41000 41004
0 41006 5 1 1 41005
0 41007 7 1 2 51414 41006
0 41008 5 1 1 41007
0 41009 7 3 2 63842 72713
0 41010 7 1 2 66052 79025
0 41011 5 1 1 41010
0 41012 7 1 2 41008 41011
0 41013 5 1 1 41012
0 41014 7 1 2 50289 41013
0 41015 5 1 1 41014
0 41016 7 5 2 72703 75002
0 41017 5 1 1 79028
0 41018 7 2 2 51991 79029
0 41019 5 1 1 79033
0 41020 7 1 2 55130 79034
0 41021 5 1 1 41020
0 41022 7 1 2 67704 41021
0 41023 5 1 1 41022
0 41024 7 1 2 67406 41023
0 41025 5 1 1 41024
0 41026 7 1 2 70336 78511
0 41027 5 1 1 41026
0 41028 7 1 2 78621 41027
0 41029 5 1 1 41028
0 41030 7 1 2 41025 41029
0 41031 5 1 1 41030
0 41032 7 1 2 50853 41031
0 41033 5 1 1 41032
0 41034 7 1 2 41015 41033
0 41035 5 1 1 41034
0 41036 7 1 2 57257 41035
0 41037 5 1 1 41036
0 41038 7 1 2 77322 78610
0 41039 5 1 1 41038
0 41040 7 2 2 59888 62644
0 41041 5 1 1 79035
0 41042 7 1 2 41039 41041
0 41043 5 1 1 41042
0 41044 7 1 2 51992 41043
0 41045 5 1 1 41044
0 41046 7 1 2 67407 76268
0 41047 5 1 1 41046
0 41048 7 2 2 56657 63534
0 41049 5 2 1 79037
0 41050 7 1 2 76329 75812
0 41051 5 1 1 41050
0 41052 7 1 2 79039 41051
0 41053 5 2 1 41052
0 41054 7 1 2 50535 79041
0 41055 5 1 1 41054
0 41056 7 1 2 41047 41055
0 41057 7 1 2 41045 41056
0 41058 5 1 1 41057
0 41059 7 1 2 58778 41058
0 41060 5 1 1 41059
0 41061 7 1 2 59889 76798
0 41062 5 1 1 41061
0 41063 7 1 2 55406 41062
0 41064 7 1 2 41060 41063
0 41065 5 1 1 41064
0 41066 7 1 2 75253 79022
0 41067 5 3 1 41066
0 41068 7 1 2 56658 79043
0 41069 5 1 1 41068
0 41070 7 1 2 70079 41069
0 41071 5 1 1 41070
0 41072 7 1 2 51993 41071
0 41073 5 1 1 41072
0 41074 7 1 2 50536 79044
0 41075 5 1 1 41074
0 41076 7 1 2 51415 41075
0 41077 7 1 2 41073 41076
0 41078 5 1 1 41077
0 41079 7 1 2 53579 41078
0 41080 7 1 2 41065 41079
0 41081 5 1 1 41080
0 41082 7 1 2 63843 77625
0 41083 5 1 1 41082
0 41084 7 1 2 68604 41083
0 41085 5 1 1 41084
0 41086 7 1 2 51994 41085
0 41087 5 1 1 41086
0 41088 7 1 2 49807 78066
0 41089 5 1 1 41088
0 41090 7 1 2 41087 41089
0 41091 5 1 1 41090
0 41092 7 1 2 56475 41091
0 41093 5 1 1 41092
0 41094 7 1 2 73125 78068
0 41095 5 1 1 41094
0 41096 7 1 2 52715 41095
0 41097 5 1 1 41096
0 41098 7 1 2 51416 71370
0 41099 5 1 1 41098
0 41100 7 1 2 41097 41099
0 41101 5 1 1 41100
0 41102 7 1 2 49808 41101
0 41103 5 1 1 41102
0 41104 7 1 2 41093 41103
0 41105 5 1 1 41104
0 41106 7 1 2 56659 41105
0 41107 5 1 1 41106
0 41108 7 1 2 73212 79016
0 41109 5 1 1 41108
0 41110 7 1 2 41107 41109
0 41111 5 1 1 41110
0 41112 7 1 2 75813 41111
0 41113 5 1 1 41112
0 41114 7 1 2 55131 73226
0 41115 7 1 2 75119 41114
0 41116 5 1 1 41115
0 41117 7 1 2 79013 41116
0 41118 5 1 1 41117
0 41119 7 1 2 67408 41118
0 41120 5 1 1 41119
0 41121 7 2 2 64599 70604
0 41122 5 3 1 79046
0 41123 7 1 2 76526 79048
0 41124 5 1 1 41123
0 41125 7 2 2 51144 72795
0 41126 7 1 2 41124 79051
0 41127 5 1 1 41126
0 41128 7 1 2 66053 78708
0 41129 5 1 1 41128
0 41130 7 1 2 41127 41129
0 41131 7 1 2 41120 41130
0 41132 5 1 1 41131
0 41133 7 1 2 50537 41132
0 41134 5 1 1 41133
0 41135 7 1 2 73806 71372
0 41136 5 1 1 41135
0 41137 7 1 2 77974 41136
0 41138 5 1 1 41137
0 41139 7 2 2 70596 76394
0 41140 5 1 1 79053
0 41141 7 1 2 63792 79054
0 41142 5 1 1 41141
0 41143 7 1 2 41138 41142
0 41144 5 1 1 41143
0 41145 7 1 2 53250 58547
0 41146 7 1 2 41144 41145
0 41147 5 1 1 41146
0 41148 7 1 2 62688 78664
0 41149 5 1 1 41148
0 41150 7 1 2 41147 41149
0 41151 7 1 2 41134 41150
0 41152 7 1 2 41113 41151
0 41153 7 1 2 41081 41152
0 41154 7 1 2 41037 41153
0 41155 5 1 1 41154
0 41156 7 1 2 53730 41155
0 41157 5 1 1 41156
0 41158 7 1 2 63619 78951
0 41159 5 1 1 41158
0 41160 7 1 2 73741 41159
0 41161 5 1 1 41160
0 41162 7 1 2 56660 41161
0 41163 5 1 1 41162
0 41164 7 2 2 63664 70605
0 41165 5 1 1 79055
0 41166 7 1 2 41163 41165
0 41167 5 1 1 41166
0 41168 7 1 2 67409 41167
0 41169 5 1 1 41168
0 41170 7 2 2 55950 72727
0 41171 5 1 1 79057
0 41172 7 1 2 73574 79058
0 41173 5 1 1 41172
0 41174 7 1 2 73742 41173
0 41175 5 1 1 41174
0 41176 7 1 2 51145 41175
0 41177 5 1 1 41176
0 41178 7 1 2 63682 71538
0 41179 5 1 1 41178
0 41180 7 1 2 63690 71510
0 41181 5 1 1 41180
0 41182 7 1 2 41179 41181
0 41183 5 1 1 41182
0 41184 7 2 2 67410 41183
0 41185 5 1 1 79059
0 41186 7 1 2 65776 73738
0 41187 5 1 1 41186
0 41188 7 1 2 41185 41187
0 41189 5 1 1 41188
0 41190 7 1 2 57258 41189
0 41191 5 1 1 41190
0 41192 7 1 2 41177 41191
0 41193 7 1 2 41169 41192
0 41194 5 1 1 41193
0 41195 7 1 2 51417 41194
0 41196 5 1 1 41195
0 41197 7 1 2 63683 76199
0 41198 7 2 2 76242 41197
0 41199 7 2 2 57259 79061
0 41200 5 1 1 79063
0 41201 7 2 2 75303 78050
0 41202 7 2 2 59157 63675
0 41203 7 1 2 79065 79067
0 41204 7 1 2 78503 41203
0 41205 5 1 1 41204
0 41206 7 1 2 41200 41205
0 41207 7 1 2 41196 41206
0 41208 5 1 1 41207
0 41209 7 1 2 49966 41208
0 41210 5 1 1 41209
0 41211 7 1 2 41157 41210
0 41212 7 1 2 40994 41211
0 41213 5 1 1 41212
0 41214 7 1 2 52819 41213
0 41215 5 1 1 41214
0 41216 7 1 2 53251 73575
0 41217 5 1 1 41216
0 41218 7 1 2 73175 41217
0 41219 5 1 1 41218
0 41220 7 1 2 52450 41219
0 41221 5 1 1 41220
0 41222 7 1 2 56661 76516
0 41223 5 1 1 41222
0 41224 7 1 2 41221 41223
0 41225 5 1 1 41224
0 41226 7 1 2 55951 41225
0 41227 5 1 1 41226
0 41228 7 1 2 74888 70634
0 41229 5 1 1 41228
0 41230 7 1 2 41227 41229
0 41231 5 1 1 41230
0 41232 7 1 2 78897 41231
0 41233 5 1 1 41232
0 41234 7 1 2 48969 73739
0 41235 5 2 1 41234
0 41236 7 1 2 41233 79069
0 41237 5 1 1 41236
0 41238 7 1 2 51146 41237
0 41239 5 1 1 41238
0 41240 7 2 2 58807 63646
0 41241 5 2 1 79071
0 41242 7 1 2 50290 63422
0 41243 5 1 1 41242
0 41244 7 1 2 79073 41243
0 41245 5 1 1 41244
0 41246 7 1 2 71511 41245
0 41247 5 1 1 41246
0 41248 7 2 2 58779 63423
0 41249 7 1 2 63684 79075
0 41250 5 1 1 41249
0 41251 7 1 2 41247 41250
0 41252 5 1 1 41251
0 41253 7 2 2 67411 41252
0 41254 5 1 1 79077
0 41255 7 3 2 52581 67962
0 41256 7 1 2 73189 76146
0 41257 7 1 2 79079 41256
0 41258 5 1 1 41257
0 41259 7 1 2 41254 41258
0 41260 5 1 1 41259
0 41261 7 1 2 57260 41260
0 41262 5 1 1 41261
0 41263 7 1 2 73002 78938
0 41264 7 1 2 67412 41263
0 41265 5 1 1 41264
0 41266 7 1 2 41262 41265
0 41267 7 1 2 41239 41266
0 41268 5 1 1 41267
0 41269 7 1 2 51418 41268
0 41270 5 1 1 41269
0 41271 7 1 2 48970 79064
0 41272 5 1 1 41271
0 41273 7 1 2 52188 73894
0 41274 7 1 2 70597 41273
0 41275 7 1 2 79068 41274
0 41276 7 1 2 78504 41275
0 41277 5 1 1 41276
0 41278 7 1 2 41272 41277
0 41279 7 1 2 41270 41278
0 41280 5 1 1 41279
0 41281 7 1 2 53731 41280
0 41282 5 1 1 41281
0 41283 7 5 2 70561 71512
0 41284 5 3 1 79082
0 41285 7 1 2 66668 79083
0 41286 7 1 2 73469 41285
0 41287 5 1 1 41286
0 41288 7 1 2 41282 41287
0 41289 7 1 2 41215 41288
0 41290 5 1 1 41289
0 41291 7 1 2 55568 41290
0 41292 5 1 1 41291
0 41293 7 1 2 40914 41292
0 41294 5 2 1 41293
0 41295 7 1 2 51775 79090
0 41296 5 1 1 41295
0 41297 7 9 2 68753 73657
0 41298 7 1 2 53252 73024
0 41299 5 1 1 41298
0 41300 7 1 2 71565 41299
0 41301 5 1 1 41300
0 41302 7 1 2 52451 41301
0 41303 5 1 1 41302
0 41304 7 1 2 50854 71621
0 41305 5 1 1 41304
0 41306 7 1 2 41303 41305
0 41307 5 1 1 41306
0 41308 7 1 2 51995 72677
0 41309 7 1 2 41307 41308
0 41310 5 1 1 41309
0 41311 7 2 2 65009 73384
0 41312 5 1 1 79101
0 41313 7 1 2 71616 41312
0 41314 7 1 2 41310 41313
0 41315 5 1 1 41314
0 41316 7 1 2 55952 41315
0 41317 5 1 1 41316
0 41318 7 1 2 55953 78243
0 41319 5 2 1 41318
0 41320 7 1 2 52452 77132
0 41321 5 3 1 41320
0 41322 7 1 2 71628 79105
0 41323 7 1 2 79103 41322
0 41324 5 1 1 41323
0 41325 7 1 2 51996 41324
0 41326 5 1 1 41325
0 41327 7 1 2 57063 65346
0 41328 5 1 1 41327
0 41329 7 1 2 73184 41328
0 41330 5 1 1 41329
0 41331 7 1 2 52189 41330
0 41332 5 1 1 41331
0 41333 7 1 2 72610 41332
0 41334 7 1 2 41326 41333
0 41335 5 1 1 41334
0 41336 7 1 2 51147 41335
0 41337 5 1 1 41336
0 41338 7 1 2 72976 71496
0 41339 7 1 2 71622 41338
0 41340 5 1 1 41339
0 41341 7 1 2 41337 41340
0 41342 7 1 2 41317 41341
0 41343 5 2 1 41342
0 41344 7 2 2 72293 79108
0 41345 7 1 2 79092 79110
0 41346 5 1 1 41345
0 41347 7 2 2 51419 58780
0 41348 5 2 1 79112
0 41349 7 3 2 56245 70606
0 41350 5 1 1 79116
0 41351 7 1 2 79114 41350
0 41352 5 1 1 41351
0 41353 7 1 2 49967 57064
0 41354 7 1 2 41352 41353
0 41355 5 1 1 41354
0 41356 7 2 2 55407 57345
0 41357 5 1 1 79119
0 41358 7 1 2 49638 41357
0 41359 5 1 1 41358
0 41360 7 1 2 53732 75062
0 41361 7 1 2 41359 41360
0 41362 5 1 1 41361
0 41363 7 1 2 41355 41362
0 41364 5 1 1 41363
0 41365 7 1 2 53580 41364
0 41366 5 1 1 41365
0 41367 7 1 2 68839 71315
0 41368 5 1 1 41367
0 41369 7 3 2 53733 56246
0 41370 7 1 2 70330 79121
0 41371 5 1 1 41370
0 41372 7 1 2 72554 41371
0 41373 5 1 1 41372
0 41374 7 1 2 41368 41373
0 41375 5 1 1 41374
0 41376 7 1 2 41366 41375
0 41377 5 1 1 41376
0 41378 7 1 2 60223 41377
0 41379 5 1 1 41378
0 41380 7 1 2 68840 78527
0 41381 5 1 1 41380
0 41382 7 1 2 51420 56247
0 41383 7 1 2 41381 41382
0 41384 5 2 1 41383
0 41385 7 1 2 41379 79124
0 41386 5 1 1 41385
0 41387 7 1 2 55569 41386
0 41388 5 1 1 41387
0 41389 7 1 2 70337 18401
0 41390 5 1 1 41389
0 41391 7 2 2 49968 41390
0 41392 7 1 2 60254 65706
0 41393 5 1 1 41392
0 41394 7 1 2 51634 41393
0 41395 7 1 2 79126 41394
0 41396 5 1 1 41395
0 41397 7 1 2 41388 41396
0 41398 5 1 1 41397
0 41399 7 1 2 52820 41398
0 41400 5 1 1 41399
0 41401 7 1 2 55570 76450
0 41402 7 1 2 78898 41401
0 41403 5 1 1 41402
0 41404 7 2 2 67141 71460
0 41405 5 1 1 79128
0 41406 7 1 2 41403 41405
0 41407 5 1 1 41406
0 41408 7 1 2 53734 41407
0 41409 5 1 1 41408
0 41410 7 1 2 74820 71312
0 41411 5 1 1 41410
0 41412 7 1 2 41409 41411
0 41413 5 1 1 41412
0 41414 7 1 2 77133 41413
0 41415 5 1 1 41414
0 41416 7 2 2 65736 71623
0 41417 5 1 1 79130
0 41418 7 1 2 48971 79131
0 41419 5 1 1 41418
0 41420 7 1 2 68566 41419
0 41421 5 1 1 41420
0 41422 7 1 2 75899 41421
0 41423 5 1 1 41422
0 41424 7 1 2 53735 79129
0 41425 5 2 1 41424
0 41426 7 1 2 41423 79132
0 41427 5 1 1 41426
0 41428 7 1 2 52453 41427
0 41429 5 1 1 41428
0 41430 7 1 2 67801 41417
0 41431 5 1 1 41430
0 41432 7 1 2 78899 41431
0 41433 5 1 1 41432
0 41434 7 1 2 66398 68834
0 41435 5 2 1 41434
0 41436 7 1 2 41433 79134
0 41437 5 1 1 41436
0 41438 7 1 2 51421 41437
0 41439 5 1 1 41438
0 41440 7 1 2 41429 41439
0 41441 7 1 2 41415 41440
0 41442 7 1 2 41400 41441
0 41443 5 1 1 41442
0 41444 7 1 2 61503 41443
0 41445 5 1 1 41444
0 41446 7 2 2 51635 78867
0 41447 7 1 2 56248 79136
0 41448 5 1 1 41447
0 41449 7 1 2 72714 78733
0 41450 5 1 1 41449
0 41451 7 1 2 41448 41450
0 41452 5 2 1 41451
0 41453 7 1 2 55408 79138
0 41454 5 1 1 41453
0 41455 7 3 2 51636 78968
0 41456 7 1 2 72551 79140
0 41457 5 1 1 41456
0 41458 7 1 2 41454 41457
0 41459 5 1 1 41458
0 41460 7 1 2 50291 41459
0 41461 5 1 1 41460
0 41462 7 1 2 41445 41461
0 41463 5 1 1 41462
0 41464 7 1 2 51148 41463
0 41465 5 1 1 41464
0 41466 7 1 2 56249 67787
0 41467 5 2 1 41466
0 41468 7 1 2 53736 75095
0 41469 5 1 1 41468
0 41470 7 1 2 79143 41469
0 41471 5 1 1 41470
0 41472 7 1 2 73833 75185
0 41473 7 1 2 41471 41472
0 41474 5 1 1 41473
0 41475 7 2 2 56476 72410
0 41476 5 1 1 79145
0 41477 7 1 2 56250 66399
0 41478 5 1 1 41477
0 41479 7 1 2 41476 41478
0 41480 5 1 1 41479
0 41481 7 1 2 78825 41480
0 41482 5 1 1 41481
0 41483 7 1 2 68631 79117
0 41484 5 1 1 41483
0 41485 7 1 2 54109 78655
0 41486 7 1 2 78738 41485
0 41487 5 1 1 41486
0 41488 7 1 2 41484 41487
0 41489 7 1 2 41482 41488
0 41490 7 1 2 41474 41489
0 41491 5 1 1 41490
0 41492 7 1 2 51422 41491
0 41493 5 1 1 41492
0 41494 7 1 2 57065 78751
0 41495 7 1 2 79030 41494
0 41496 5 1 1 41495
0 41497 7 1 2 41493 41496
0 41498 5 1 1 41497
0 41499 7 1 2 60562 41498
0 41500 5 1 1 41499
0 41501 7 1 2 41465 41500
0 41502 5 2 1 41501
0 41503 7 1 2 51776 79147
0 41504 5 1 1 41503
0 41505 7 1 2 52454 78064
0 41506 5 3 1 41505
0 41507 7 1 2 51149 77781
0 41508 5 1 1 41507
0 41509 7 1 2 79149 41508
0 41510 5 2 1 41509
0 41511 7 2 2 72294 79152
0 41512 7 1 2 79093 79154
0 41513 5 1 1 41512
0 41514 7 1 2 41504 41513
0 41515 5 1 1 41514
0 41516 7 1 2 57261 41515
0 41517 5 1 1 41516
0 41518 7 1 2 53737 78562
0 41519 5 1 1 41518
0 41520 7 1 2 78833 41519
0 41521 5 1 1 41520
0 41522 7 1 2 52821 41521
0 41523 5 1 1 41522
0 41524 7 1 2 79087 41523
0 41525 5 1 1 41524
0 41526 7 1 2 73686 41525
0 41527 5 1 1 41526
0 41528 7 1 2 51150 79141
0 41529 5 1 1 41528
0 41530 7 1 2 41527 41529
0 41531 5 1 1 41530
0 41532 7 1 2 51423 41531
0 41533 5 1 1 41532
0 41534 7 1 2 61695 73904
0 41535 7 1 2 79137 41534
0 41536 5 1 1 41535
0 41537 7 1 2 41533 41536
0 41538 5 1 1 41537
0 41539 7 1 2 50538 41538
0 41540 5 1 1 41539
0 41541 7 1 2 61047 73373
0 41542 7 1 2 79142 41541
0 41543 5 1 1 41542
0 41544 7 2 2 63620 65737
0 41545 7 1 2 73827 70616
0 41546 7 1 2 79156 41545
0 41547 5 1 1 41546
0 41548 7 1 2 41543 41547
0 41549 5 1 1 41548
0 41550 7 1 2 51151 41549
0 41551 5 1 1 41550
0 41552 7 1 2 73766 71373
0 41553 5 1 1 41552
0 41554 7 1 2 62982 41553
0 41555 5 1 1 41554
0 41556 7 1 2 51152 73863
0 41557 5 1 1 41556
0 41558 7 1 2 15574 41557
0 41559 7 1 2 41555 41558
0 41560 5 1 1 41559
0 41561 7 1 2 67857 41560
0 41562 5 1 1 41561
0 41563 7 1 2 59890 69314
0 41564 7 1 2 75900 41563
0 41565 5 1 1 41564
0 41566 7 1 2 41562 41565
0 41567 5 1 1 41566
0 41568 7 1 2 51637 41567
0 41569 5 1 1 41568
0 41570 7 2 2 58781 77323
0 41571 5 1 1 79158
0 41572 7 1 2 79004 41571
0 41573 5 2 1 41572
0 41574 7 1 2 53581 79160
0 41575 5 1 1 41574
0 41576 7 1 2 70607 79159
0 41577 5 1 1 41576
0 41578 7 1 2 41575 41577
0 41579 5 1 1 41578
0 41580 7 1 2 50292 69714
0 41581 7 1 2 41579 41580
0 41582 5 1 1 41581
0 41583 7 1 2 38570 41582
0 41584 5 1 1 41583
0 41585 7 1 2 69530 41584
0 41586 5 1 1 41585
0 41587 7 1 2 41569 41586
0 41588 5 1 1 41587
0 41589 7 1 2 55409 41588
0 41590 5 1 1 41589
0 41591 7 1 2 41551 41590
0 41592 7 1 2 41540 41591
0 41593 5 2 1 41592
0 41594 7 1 2 51777 79162
0 41595 5 1 1 41594
0 41596 7 2 2 73849 72876
0 41597 7 1 2 79094 79164
0 41598 5 1 1 41597
0 41599 7 1 2 41595 41598
0 41600 5 1 1 41599
0 41601 7 1 2 57066 41600
0 41602 5 1 1 41601
0 41603 7 3 2 51153 78868
0 41604 7 2 2 56251 79166
0 41605 7 1 2 73003 79169
0 41606 5 1 1 41605
0 41607 7 1 2 73576 78988
0 41608 5 1 1 41607
0 41609 7 1 2 41606 41608
0 41610 5 1 1 41609
0 41611 7 1 2 55410 41610
0 41612 5 1 1 41611
0 41613 7 1 2 56662 78976
0 41614 5 1 1 41613
0 41615 7 1 2 59164 41614
0 41616 5 1 1 41615
0 41617 7 3 2 50293 41616
0 41618 7 1 2 78969 79171
0 41619 5 1 1 41618
0 41620 7 2 2 69931 78869
0 41621 5 1 1 79174
0 41622 7 1 2 51997 79175
0 41623 5 1 1 41622
0 41624 7 1 2 41619 41623
0 41625 5 1 1 41624
0 41626 7 1 2 51424 41625
0 41627 5 1 1 41626
0 41628 7 1 2 41612 41627
0 41629 5 2 1 41628
0 41630 7 1 2 51778 79176
0 41631 5 1 1 41630
0 41632 7 2 2 68528 79172
0 41633 7 1 2 79095 79178
0 41634 5 1 1 41633
0 41635 7 1 2 41631 41634
0 41636 5 1 1 41635
0 41637 7 1 2 51638 41636
0 41638 5 1 1 41637
0 41639 7 1 2 78650 78952
0 41640 5 1 1 41639
0 41641 7 1 2 73743 41640
0 41642 5 1 1 41641
0 41643 7 1 2 56252 41642
0 41644 5 1 1 41643
0 41645 7 1 2 59026 73418
0 41646 7 1 2 79066 41645
0 41647 5 1 1 41646
0 41648 7 1 2 41644 41647
0 41649 5 1 1 41648
0 41650 7 1 2 67888 41649
0 41651 5 1 1 41650
0 41652 7 1 2 71277 76330
0 41653 5 1 1 41652
0 41654 7 1 2 79040 41653
0 41655 5 1 1 41654
0 41656 7 1 2 75003 41655
0 41657 5 1 1 41656
0 41658 7 1 2 57346 76364
0 41659 5 1 1 41658
0 41660 7 1 2 75254 41659
0 41661 5 1 1 41660
0 41662 7 1 2 51425 41661
0 41663 5 1 1 41662
0 41664 7 1 2 41657 41663
0 41665 5 1 1 41664
0 41666 7 1 2 53582 41665
0 41667 5 1 1 41666
0 41668 7 1 2 73634 76524
0 41669 5 1 1 41668
0 41670 7 1 2 79049 41669
0 41671 5 1 1 41670
0 41672 7 1 2 63705 41671
0 41673 5 1 1 41672
0 41674 7 1 2 56253 79018
0 41675 5 1 1 41674
0 41676 7 1 2 41673 41675
0 41677 7 1 2 41667 41676
0 41678 5 1 1 41677
0 41679 7 1 2 51998 41678
0 41680 5 1 1 41679
0 41681 7 3 2 69810 68882
0 41682 7 1 2 56254 79180
0 41683 5 1 1 41682
0 41684 7 1 2 76592 41683
0 41685 5 1 1 41684
0 41686 7 1 2 56663 41685
0 41687 5 1 1 41686
0 41688 7 2 2 62645 72890
0 41689 5 1 1 79183
0 41690 7 1 2 41687 41689
0 41691 5 1 1 41690
0 41692 7 1 2 58782 41691
0 41693 5 1 1 41692
0 41694 7 1 2 63185 78662
0 41695 5 1 1 41694
0 41696 7 2 2 63599 76023
0 41697 7 1 2 71067 79185
0 41698 5 1 1 41697
0 41699 7 1 2 41695 41698
0 41700 5 1 1 41699
0 41701 7 1 2 77324 41700
0 41702 5 1 1 41701
0 41703 7 1 2 63621 78706
0 41704 5 1 1 41703
0 41705 7 1 2 50539 79047
0 41706 5 1 1 41705
0 41707 7 1 2 41704 41706
0 41708 5 1 1 41707
0 41709 7 1 2 51154 41708
0 41710 5 1 1 41709
0 41711 7 1 2 41702 41710
0 41712 7 1 2 41693 41711
0 41713 7 1 2 41680 41712
0 41714 5 1 1 41713
0 41715 7 1 2 53738 41714
0 41716 5 1 1 41715
0 41717 7 1 2 41651 41716
0 41718 5 1 1 41717
0 41719 7 1 2 52822 41718
0 41720 5 1 1 41719
0 41721 7 1 2 78651 78930
0 41722 5 1 1 41721
0 41723 7 1 2 79070 41722
0 41724 5 1 1 41723
0 41725 7 1 2 56255 41724
0 41726 5 1 1 41725
0 41727 7 1 2 71595 77485
0 41728 7 1 2 79080 41727
0 41729 5 1 1 41728
0 41730 7 1 2 41726 41729
0 41731 5 1 1 41730
0 41732 7 1 2 69286 41731
0 41733 5 1 1 41732
0 41734 7 1 2 41720 41733
0 41735 5 1 1 41734
0 41736 7 2 2 67953 41735
0 41737 5 1 1 79187
0 41738 7 1 2 41638 41737
0 41739 7 1 2 41602 41738
0 41740 7 1 2 41517 41739
0 41741 5 1 1 41740
0 41742 7 1 2 57666 41741
0 41743 5 1 1 41742
0 41744 7 1 2 41346 41743
0 41745 7 1 2 41296 41744
0 41746 5 1 1 41745
0 41747 7 1 2 58448 41746
0 41748 5 1 1 41747
0 41749 7 2 2 51155 78310
0 41750 5 1 1 79189
0 41751 7 1 2 60343 59867
0 41752 5 1 1 41751
0 41753 7 1 2 74913 41752
0 41754 5 1 1 41753
0 41755 7 1 2 51999 41754
0 41756 5 1 1 41755
0 41757 7 1 2 65347 1486
0 41758 5 1 1 41757
0 41759 7 1 2 41756 41758
0 41760 5 1 1 41759
0 41761 7 1 2 57667 41760
0 41762 5 1 1 41761
0 41763 7 1 2 59868 70743
0 41764 5 1 1 41763
0 41765 7 1 2 59770 41764
0 41766 5 1 1 41765
0 41767 7 1 2 52190 41766
0 41768 5 1 1 41767
0 41769 7 2 2 65010 60685
0 41770 5 1 1 79191
0 41771 7 1 2 21274 41770
0 41772 5 1 1 41771
0 41773 7 1 2 52000 41772
0 41774 5 1 1 41773
0 41775 7 1 2 55954 58141
0 41776 5 1 1 41775
0 41777 7 1 2 70355 41776
0 41778 5 1 1 41777
0 41779 7 1 2 50294 41778
0 41780 5 1 1 41779
0 41781 7 1 2 61142 41780
0 41782 7 1 2 41774 41781
0 41783 7 1 2 41768 41782
0 41784 7 1 2 41762 41783
0 41785 5 1 1 41784
0 41786 7 1 2 50855 41785
0 41787 5 1 1 41786
0 41788 7 1 2 65450 60454
0 41789 5 1 1 41788
0 41790 7 1 2 52001 41789
0 41791 5 1 1 41790
0 41792 7 1 2 57668 78034
0 41793 5 1 1 41792
0 41794 7 1 2 41791 41793
0 41795 5 1 1 41794
0 41796 7 1 2 50856 41795
0 41797 5 1 1 41796
0 41798 7 1 2 59907 41797
0 41799 5 1 1 41798
0 41800 7 1 2 58449 41799
0 41801 5 1 1 41800
0 41802 7 1 2 55829 67354
0 41803 5 1 1 41802
0 41804 7 1 2 51156 41803
0 41805 5 1 1 41804
0 41806 7 1 2 41801 41805
0 41807 7 1 2 41787 41806
0 41808 5 1 1 41807
0 41809 7 1 2 51426 41808
0 41810 5 1 1 41809
0 41811 7 1 2 41750 41810
0 41812 5 1 1 41811
0 41813 7 1 2 49809 41812
0 41814 5 1 1 41813
0 41815 7 1 2 57669 76760
0 41816 5 1 1 41815
0 41817 7 1 2 53010 75167
0 41818 5 1 1 41817
0 41819 7 1 2 41816 41818
0 41820 5 1 1 41819
0 41821 7 1 2 52907 41820
0 41822 5 1 1 41821
0 41823 7 1 2 50295 59070
0 41824 5 1 1 41823
0 41825 7 1 2 41822 41824
0 41826 5 1 1 41825
0 41827 7 1 2 52002 41826
0 41828 5 1 1 41827
0 41829 7 2 2 50296 58142
0 41830 5 1 1 79193
0 41831 7 1 2 63122 79194
0 41832 5 1 1 41831
0 41833 7 1 2 74897 41832
0 41834 7 1 2 41828 41833
0 41835 5 1 1 41834
0 41836 7 1 2 63535 41835
0 41837 5 1 1 41836
0 41838 7 1 2 63536 9761
0 41839 5 1 1 41838
0 41840 7 1 2 63537 76785
0 41841 5 1 1 41840
0 41842 7 1 2 25789 41841
0 41843 5 1 1 41842
0 41844 7 1 2 76780 41843
0 41845 5 1 1 41844
0 41846 7 1 2 41839 41845
0 41847 5 1 1 41846
0 41848 7 1 2 50540 41847
0 41849 5 1 1 41848
0 41850 7 1 2 63538 70258
0 41851 5 1 1 41850
0 41852 7 1 2 52003 59165
0 41853 7 1 2 73074 41852
0 41854 5 1 1 41853
0 41855 7 1 2 41851 41854
0 41856 5 1 1 41855
0 41857 7 1 2 62229 41856
0 41858 5 1 1 41857
0 41859 7 1 2 61075 78277
0 41860 5 1 1 41859
0 41861 7 1 2 25993 41860
0 41862 5 1 1 41861
0 41863 7 1 2 57262 41862
0 41864 5 1 1 41863
0 41865 7 1 2 74994 41864
0 41866 7 1 2 41858 41865
0 41867 7 1 2 41849 41866
0 41868 7 1 2 41837 41867
0 41869 5 1 1 41868
0 41870 7 1 2 78598 41869
0 41871 5 1 1 41870
0 41872 7 1 2 41814 41871
0 41873 5 1 1 41872
0 41874 7 1 2 53253 41873
0 41875 5 1 1 41874
0 41876 7 1 2 58450 60154
0 41877 5 1 1 41876
0 41878 7 2 2 60874 41877
0 41879 7 1 2 63497 79195
0 41880 5 1 1 41879
0 41881 7 1 2 76030 41880
0 41882 5 1 1 41881
0 41883 7 1 2 50297 62241
0 41884 5 1 1 41883
0 41885 7 1 2 57670 62049
0 41886 5 1 1 41885
0 41887 7 1 2 74676 41886
0 41888 7 1 2 41884 41887
0 41889 5 1 1 41888
0 41890 7 1 2 52004 41889
0 41891 5 1 1 41890
0 41892 7 1 2 54110 62104
0 41893 5 1 1 41892
0 41894 7 1 2 54410 62225
0 41895 5 1 1 41894
0 41896 7 1 2 41893 41895
0 41897 5 1 1 41896
0 41898 7 1 2 57671 74669
0 41899 5 2 1 41898
0 41900 7 1 2 60638 77031
0 41901 7 1 2 79197 41900
0 41902 7 1 2 41897 41901
0 41903 7 1 2 41891 41902
0 41904 5 1 1 41903
0 41905 7 1 2 72171 41904
0 41906 5 1 1 41905
0 41907 7 1 2 41882 41906
0 41908 5 1 1 41907
0 41909 7 1 2 53011 41908
0 41910 5 1 1 41909
0 41911 7 1 2 41875 41910
0 41912 5 1 1 41911
0 41913 7 1 2 52455 41912
0 41914 5 1 1 41913
0 41915 7 1 2 55132 9292
0 41916 5 2 1 41915
0 41917 7 1 2 61188 70206
0 41918 5 3 1 41917
0 41919 7 1 2 59572 63140
0 41920 7 1 2 79201 41919
0 41921 5 1 1 41920
0 41922 7 1 2 73385 41921
0 41923 5 1 1 41922
0 41924 7 1 2 49503 41923
0 41925 5 1 1 41924
0 41926 7 1 2 79199 41925
0 41927 5 1 1 41926
0 41928 7 1 2 48826 41927
0 41929 5 1 1 41928
0 41930 7 1 2 50857 41929
0 41931 5 1 1 41930
0 41932 7 1 2 55133 22278
0 41933 7 1 2 64359 41932
0 41934 5 1 1 41933
0 41935 7 1 2 52716 41934
0 41936 5 1 1 41935
0 41937 7 1 2 65447 70813
0 41938 5 1 1 41937
0 41939 7 1 2 52717 59559
0 41940 5 1 1 41939
0 41941 7 1 2 72798 72772
0 41942 5 1 1 41941
0 41943 7 1 2 41940 41942
0 41944 5 1 1 41943
0 41945 7 1 2 70259 41944
0 41946 5 1 1 41945
0 41947 7 1 2 41938 41946
0 41948 7 1 2 41936 41947
0 41949 7 1 2 71438 25111
0 41950 5 1 1 41949
0 41951 7 1 2 52005 41950
0 41952 5 1 1 41951
0 41953 7 1 2 63647 72760
0 41954 5 1 1 41953
0 41955 7 1 2 41952 41954
0 41956 5 1 1 41955
0 41957 7 1 2 76761 41956
0 41958 5 1 1 41957
0 41959 7 1 2 48827 75137
0 41960 5 1 1 41959
0 41961 7 1 2 60840 57787
0 41962 5 1 1 41961
0 41963 7 1 2 57672 41962
0 41964 7 1 2 41960 41963
0 41965 5 1 1 41964
0 41966 7 1 2 41958 41965
0 41967 7 1 2 41948 41966
0 41968 7 1 2 41931 41967
0 41969 5 1 1 41968
0 41970 7 1 2 51427 41969
0 41971 5 1 1 41970
0 41972 7 1 2 57263 63397
0 41973 5 1 1 41972
0 41974 7 1 2 76781 76790
0 41975 5 1 1 41974
0 41976 7 1 2 71009 41975
0 41977 5 1 1 41976
0 41978 7 1 2 50541 41977
0 41979 5 1 1 41978
0 41980 7 1 2 71026 41979
0 41981 7 1 2 41973 41980
0 41982 5 1 1 41981
0 41983 7 1 2 79190 41982
0 41984 5 1 1 41983
0 41985 7 1 2 41971 41984
0 41986 5 1 1 41985
0 41987 7 1 2 49810 41986
0 41988 5 1 1 41987
0 41989 7 1 2 73099 73489
0 41990 5 1 1 41989
0 41991 7 1 2 73503 41990
0 41992 5 1 1 41991
0 41993 7 1 2 50298 41992
0 41994 5 1 1 41993
0 41995 7 1 2 39009 41994
0 41996 5 1 1 41995
0 41997 7 1 2 49811 41996
0 41998 5 1 1 41997
0 41999 7 1 2 73482 78716
0 42000 5 1 1 41999
0 42001 7 2 2 51428 57673
0 42002 7 1 2 62689 79204
0 42003 5 1 1 42002
0 42004 7 1 2 76032 42003
0 42005 5 1 1 42004
0 42006 7 1 2 70492 42005
0 42007 5 1 1 42006
0 42008 7 1 2 60224 61440
0 42009 7 1 2 77615 42008
0 42010 5 1 1 42009
0 42011 7 1 2 42007 42010
0 42012 5 1 1 42011
0 42013 7 1 2 52006 42012
0 42014 5 1 1 42013
0 42015 7 1 2 42000 42014
0 42016 7 1 2 41998 42015
0 42017 5 1 1 42016
0 42018 7 1 2 53012 42017
0 42019 5 1 1 42018
0 42020 7 1 2 73483 79181
0 42021 5 1 1 42020
0 42022 7 1 2 62363 70923
0 42023 5 1 1 42022
0 42024 7 1 2 48828 42023
0 42025 5 1 1 42024
0 42026 7 1 2 73122 42025
0 42027 5 1 1 42026
0 42028 7 1 2 73477 72732
0 42029 5 1 1 42028
0 42030 7 1 2 42027 42029
0 42031 5 1 1 42030
0 42032 7 1 2 52332 42031
0 42033 5 1 1 42032
0 42034 7 1 2 70993 73500
0 42035 5 1 1 42034
0 42036 7 1 2 42033 42035
0 42037 5 1 1 42036
0 42038 7 1 2 49812 42037
0 42039 5 1 1 42038
0 42040 7 1 2 42021 42039
0 42041 7 1 2 42019 42040
0 42042 5 1 1 42041
0 42043 7 1 2 58451 42042
0 42044 5 1 1 42043
0 42045 7 1 2 60739 63386
0 42046 5 1 1 42045
0 42047 7 1 2 63123 42046
0 42048 5 1 1 42047
0 42049 7 1 2 52007 76786
0 42050 5 2 1 42049
0 42051 7 1 2 60328 79206
0 42052 5 1 1 42051
0 42053 7 1 2 55955 42052
0 42054 5 1 1 42053
0 42055 7 1 2 60225 62242
0 42056 5 1 1 42055
0 42057 7 1 2 50858 75391
0 42058 5 1 1 42057
0 42059 7 1 2 42056 42058
0 42060 7 1 2 42054 42059
0 42061 7 1 2 42048 42060
0 42062 5 1 1 42061
0 42063 7 1 2 53013 42062
0 42064 5 1 1 42063
0 42065 7 1 2 9529 79207
0 42066 5 1 1 42065
0 42067 7 1 2 62220 42066
0 42068 5 1 1 42067
0 42069 7 1 2 55956 65828
0 42070 5 1 1 42069
0 42071 7 1 2 42068 42070
0 42072 5 1 1 42071
0 42073 7 1 2 50542 42072
0 42074 5 1 1 42073
0 42075 7 1 2 50109 71018
0 42076 7 1 2 76858 42075
0 42077 5 1 1 42076
0 42078 7 1 2 55134 42077
0 42079 7 1 2 42074 42078
0 42080 7 1 2 42064 42079
0 42081 5 1 1 42080
0 42082 7 1 2 59166 76419
0 42083 7 1 2 42081 42082
0 42084 5 1 1 42083
0 42085 7 1 2 42044 42084
0 42086 7 1 2 41988 42085
0 42087 7 1 2 41914 42086
0 42088 5 1 1 42087
0 42089 7 1 2 53739 42088
0 42090 5 1 1 42089
0 42091 7 1 2 52008 76977
0 42092 5 1 1 42091
0 42093 7 1 2 70266 42092
0 42094 5 1 1 42093
0 42095 7 1 2 52191 42094
0 42096 5 1 1 42095
0 42097 7 1 2 54411 41830
0 42098 5 1 1 42097
0 42099 7 1 2 53131 42098
0 42100 5 1 1 42099
0 42101 7 1 2 42096 42100
0 42102 5 1 1 42101
0 42103 7 1 2 52333 42102
0 42104 5 1 1 42103
0 42105 7 1 2 65353 77365
0 42106 5 1 1 42105
0 42107 7 1 2 61594 42106
0 42108 5 1 1 42107
0 42109 7 1 2 42104 42108
0 42110 5 1 1 42109
0 42111 7 1 2 52456 42110
0 42112 5 1 1 42111
0 42113 7 1 2 70657 76711
0 42114 5 1 1 42113
0 42115 7 1 2 42112 42114
0 42116 5 1 1 42115
0 42117 7 1 2 62364 42116
0 42118 5 1 1 42117
0 42119 7 1 2 73388 25754
0 42120 5 1 1 42119
0 42121 7 1 2 52334 42120
0 42122 5 1 1 42121
0 42123 7 1 2 38692 42122
0 42124 5 1 1 42123
0 42125 7 1 2 76371 42124
0 42126 5 1 1 42125
0 42127 7 1 2 71281 42126
0 42128 5 1 1 42127
0 42129 7 1 2 50110 42128
0 42130 5 1 1 42129
0 42131 7 1 2 62035 73182
0 42132 5 1 1 42131
0 42133 7 1 2 14921 42132
0 42134 5 1 1 42133
0 42135 7 1 2 52457 42134
0 42136 5 1 1 42135
0 42137 7 1 2 73386 73876
0 42138 5 1 1 42137
0 42139 7 1 2 42136 42138
0 42140 7 1 2 42130 42139
0 42141 5 1 1 42140
0 42142 7 1 2 52192 42141
0 42143 5 1 1 42142
0 42144 7 1 2 71209 70856
0 42145 5 1 1 42144
0 42146 7 2 2 50111 59158
0 42147 5 1 1 79208
0 42148 7 1 2 79150 42147
0 42149 5 1 1 42148
0 42150 7 1 2 57674 42149
0 42151 5 1 1 42150
0 42152 7 1 2 56256 60686
0 42153 5 1 1 42152
0 42154 7 1 2 55135 42153
0 42155 5 1 1 42154
0 42156 7 1 2 60563 42155
0 42157 5 1 1 42156
0 42158 7 1 2 42151 42157
0 42159 5 1 1 42158
0 42160 7 1 2 53014 42159
0 42161 5 1 1 42160
0 42162 7 1 2 42145 42161
0 42163 7 1 2 42143 42162
0 42164 5 1 1 42163
0 42165 7 1 2 60948 42164
0 42166 5 1 1 42165
0 42167 7 1 2 76645 76628
0 42168 5 1 1 42167
0 42169 7 1 2 73389 42168
0 42170 5 1 1 42169
0 42171 7 1 2 57675 42170
0 42172 5 1 1 42171
0 42173 7 1 2 56257 70744
0 42174 5 2 1 42173
0 42175 7 1 2 22578 79210
0 42176 5 1 1 42175
0 42177 7 1 2 53015 42176
0 42178 5 1 1 42177
0 42179 7 1 2 42172 42178
0 42180 5 1 1 42179
0 42181 7 1 2 50859 42180
0 42182 5 1 1 42181
0 42183 7 2 2 53016 60494
0 42184 5 1 1 79212
0 42185 7 1 2 49504 42184
0 42186 5 1 1 42185
0 42187 7 1 2 76072 42186
0 42188 5 1 1 42187
0 42189 7 1 2 42182 42188
0 42190 5 1 1 42189
0 42191 7 1 2 76859 42190
0 42192 5 1 1 42191
0 42193 7 3 2 52193 58840
0 42194 7 1 2 62298 78103
0 42195 5 1 1 42194
0 42196 7 1 2 13463 42195
0 42197 5 1 1 42196
0 42198 7 1 2 52335 42197
0 42199 5 1 1 42198
0 42200 7 1 2 42199 40528
0 42201 5 1 1 42200
0 42202 7 1 2 79214 42201
0 42203 5 1 1 42202
0 42204 7 1 2 53254 63910
0 42205 5 1 1 42204
0 42206 7 1 2 77911 79198
0 42207 7 1 2 61076 65901
0 42208 5 1 1 42207
0 42209 7 1 2 57676 79215
0 42210 5 1 1 42209
0 42211 7 1 2 42208 42210
0 42212 7 1 2 42206 42211
0 42213 5 1 1 42212
0 42214 7 1 2 53017 42213
0 42215 5 1 1 42214
0 42216 7 1 2 42205 42215
0 42217 5 1 1 42216
0 42218 7 1 2 52458 42217
0 42219 5 1 1 42218
0 42220 7 1 2 63134 61149
0 42221 5 1 1 42220
0 42222 7 1 2 50860 68031
0 42223 5 1 1 42222
0 42224 7 1 2 42221 42223
0 42225 5 1 1 42224
0 42226 7 1 2 53018 42225
0 42227 5 1 1 42226
0 42228 7 1 2 62376 42227
0 42229 7 1 2 42219 42228
0 42230 7 1 2 42203 42229
0 42231 5 1 1 42230
0 42232 7 1 2 51157 42231
0 42233 5 1 1 42232
0 42234 7 1 2 42192 42233
0 42235 7 1 2 42166 42234
0 42236 7 1 2 42118 42235
0 42237 5 2 1 42236
0 42238 7 2 2 62498 67889
0 42239 5 2 1 79219
0 42240 7 1 2 79217 79220
0 42241 5 1 1 42240
0 42242 7 1 2 42090 42241
0 42243 5 1 1 42242
0 42244 7 1 2 52823 42243
0 42245 5 1 1 42244
0 42246 7 1 2 75089 75164
0 42247 7 1 2 79218 42246
0 42248 5 1 1 42247
0 42249 7 1 2 17369 78862
0 42250 5 6 1 42249
0 42251 7 1 2 52194 62381
0 42252 5 1 1 42251
0 42253 7 1 2 9745 42252
0 42254 5 1 1 42253
0 42255 7 1 2 58841 42254
0 42256 5 1 1 42255
0 42257 7 1 2 58895 70686
0 42258 5 1 1 42257
0 42259 7 1 2 62385 42258
0 42260 5 1 1 42259
0 42261 7 1 2 57677 42260
0 42262 5 1 1 42261
0 42263 7 1 2 42256 42262
0 42264 5 1 1 42263
0 42265 7 1 2 50543 42264
0 42266 5 1 1 42265
0 42267 7 1 2 60949 71094
0 42268 7 1 2 76777 42267
0 42269 5 1 1 42268
0 42270 7 1 2 42266 42269
0 42271 5 1 1 42270
0 42272 7 1 2 79223 42271
0 42273 5 1 1 42272
0 42274 7 2 2 52718 68113
0 42275 7 1 2 74243 79229
0 42276 5 1 1 42275
0 42277 7 1 2 42273 42276
0 42278 5 1 1 42277
0 42279 7 1 2 51429 42278
0 42280 5 1 1 42279
0 42281 7 1 2 52908 78051
0 42282 7 1 2 59800 42281
0 42283 5 1 1 42282
0 42284 7 1 2 73486 42283
0 42285 5 1 1 42284
0 42286 7 1 2 42285 79072
0 42287 5 1 1 42286
0 42288 7 1 2 53583 78546
0 42289 5 1 1 42288
0 42290 7 1 2 73268 77501
0 42291 5 1 1 42290
0 42292 7 1 2 42289 42291
0 42293 5 1 1 42292
0 42294 7 1 2 52009 42293
0 42295 5 1 1 42294
0 42296 7 1 2 76430 77502
0 42297 5 1 1 42296
0 42298 7 1 2 76258 42297
0 42299 5 1 1 42298
0 42300 7 1 2 52195 42299
0 42301 5 1 1 42300
0 42302 7 1 2 42295 42301
0 42303 5 1 1 42302
0 42304 7 1 2 52719 42303
0 42305 5 1 1 42304
0 42306 7 1 2 68114 68316
0 42307 7 1 2 70662 42306
0 42308 5 1 1 42307
0 42309 7 1 2 42305 42308
0 42310 5 1 1 42309
0 42311 7 1 2 57678 42310
0 42312 5 1 1 42311
0 42313 7 1 2 55136 73290
0 42314 7 1 2 79230 42313
0 42315 5 1 1 42314
0 42316 7 1 2 63539 76860
0 42317 5 1 1 42316
0 42318 7 1 2 58902 76091
0 42319 5 1 1 42318
0 42320 7 1 2 42317 42319
0 42321 5 1 1 42320
0 42322 7 1 2 62983 78248
0 42323 7 1 2 42321 42322
0 42324 5 1 1 42323
0 42325 7 1 2 42315 42324
0 42326 7 1 2 42312 42325
0 42327 5 1 1 42326
0 42328 7 1 2 55411 42327
0 42329 5 1 1 42328
0 42330 7 1 2 42287 42329
0 42331 5 1 1 42330
0 42332 7 1 2 69531 42331
0 42333 5 1 1 42332
0 42334 7 1 2 42280 42333
0 42335 5 1 1 42334
0 42336 7 1 2 76848 42335
0 42337 5 1 1 42336
0 42338 7 1 2 55571 42337
0 42339 7 1 2 42248 42338
0 42340 7 1 2 42245 42339
0 42341 5 1 1 42340
0 42342 7 2 2 62984 68670
0 42343 5 2 1 79231
0 42344 7 1 2 73611 70482
0 42345 5 1 1 42344
0 42346 7 1 2 79233 42345
0 42347 5 2 1 42346
0 42348 7 1 2 58452 79235
0 42349 5 1 1 42348
0 42350 7 2 2 66613 70483
0 42351 7 2 2 60711 79237
0 42352 5 1 1 79239
0 42353 7 1 2 42349 42352
0 42354 5 1 1 42353
0 42355 7 1 2 49969 42354
0 42356 5 1 1 42355
0 42357 7 3 2 67858 78599
0 42358 7 2 2 52010 79241
0 42359 5 1 1 79244
0 42360 7 3 2 67123 78600
0 42361 5 2 1 79246
0 42362 7 1 2 58453 79247
0 42363 5 1 1 42362
0 42364 7 1 2 42359 42363
0 42365 7 1 2 42356 42364
0 42366 5 1 1 42365
0 42367 7 1 2 52196 42366
0 42368 5 1 1 42367
0 42369 7 3 2 62985 76586
0 42370 7 2 2 67859 79251
0 42371 5 1 1 79254
0 42372 7 1 2 42368 42371
0 42373 5 1 1 42372
0 42374 7 1 2 57679 42373
0 42375 5 1 1 42374
0 42376 7 2 2 62180 79252
0 42377 7 1 2 73162 79256
0 42378 5 1 1 42377
0 42379 7 1 2 54111 76920
0 42380 5 1 1 42379
0 42381 7 1 2 70687 76529
0 42382 7 1 2 70484 42381
0 42383 7 1 2 42380 42382
0 42384 5 1 1 42383
0 42385 7 1 2 42378 42384
0 42386 5 1 1 42385
0 42387 7 1 2 49970 42386
0 42388 5 1 1 42387
0 42389 7 1 2 52197 67124
0 42390 7 1 2 79257 42389
0 42391 5 1 1 42390
0 42392 7 1 2 42388 42391
0 42393 7 1 2 42375 42392
0 42394 5 1 1 42393
0 42395 7 1 2 50544 42394
0 42396 5 1 1 42395
0 42397 7 1 2 27686 79242
0 42398 5 1 1 42397
0 42399 7 2 2 52336 79238
0 42400 5 1 1 79258
0 42401 7 1 2 71072 74836
0 42402 7 1 2 79259 42401
0 42403 5 1 1 42402
0 42404 7 1 2 42398 42403
0 42405 5 1 1 42404
0 42406 7 1 2 60344 42405
0 42407 5 1 1 42406
0 42408 7 1 2 60155 61732
0 42409 5 2 1 42408
0 42410 7 1 2 70756 79260
0 42411 5 1 1 42410
0 42412 7 1 2 73093 78521
0 42413 7 1 2 42411 42412
0 42414 5 1 1 42413
0 42415 7 1 2 42407 42414
0 42416 7 1 2 42396 42415
0 42417 5 1 1 42416
0 42418 7 1 2 50861 42417
0 42419 5 1 1 42418
0 42420 7 1 2 74078 78572
0 42421 5 1 1 42420
0 42422 7 2 2 61461 70905
0 42423 5 1 1 79262
0 42424 7 1 2 49381 79263
0 42425 5 1 1 42424
0 42426 7 1 2 50299 42425
0 42427 5 1 1 42426
0 42428 7 2 2 58631 62067
0 42429 5 2 1 79264
0 42430 7 1 2 57680 79266
0 42431 5 1 1 42430
0 42432 7 1 2 50545 70218
0 42433 5 1 1 42432
0 42434 7 1 2 42431 42433
0 42435 7 1 2 42427 42434
0 42436 5 1 1 42435
0 42437 7 1 2 52011 42436
0 42438 5 1 1 42437
0 42439 7 1 2 57681 60865
0 42440 5 1 1 42439
0 42441 7 1 2 65380 42440
0 42442 5 1 1 42441
0 42443 7 1 2 57264 42442
0 42444 5 1 1 42443
0 42445 7 1 2 70405 69160
0 42446 5 1 1 42445
0 42447 7 1 2 70746 77264
0 42448 7 1 2 42446 42447
0 42449 7 1 2 42444 42448
0 42450 7 1 2 42438 42449
0 42451 5 2 1 42450
0 42452 7 1 2 50862 79268
0 42453 5 1 1 42452
0 42454 7 2 2 52337 75217
0 42455 5 1 1 79270
0 42456 7 1 2 42453 42455
0 42457 5 1 1 42456
0 42458 7 1 2 71084 70485
0 42459 7 1 2 42457 42458
0 42460 5 1 1 42459
0 42461 7 1 2 42421 42460
0 42462 5 1 1 42461
0 42463 7 1 2 51430 42462
0 42464 5 1 1 42463
0 42465 7 1 2 61189 71142
0 42466 5 1 1 42465
0 42467 7 1 2 61143 42466
0 42468 5 1 1 42467
0 42469 7 1 2 50300 42468
0 42470 5 1 1 42469
0 42471 7 1 2 50863 60895
0 42472 5 1 1 42471
0 42473 7 1 2 55137 42472
0 42474 7 1 2 42470 42473
0 42475 7 1 2 54800 9685
0 42476 5 1 1 42475
0 42477 7 1 2 50546 42476
0 42478 5 1 1 42477
0 42479 7 1 2 50547 61454
0 42480 5 1 1 42479
0 42481 7 1 2 50864 70729
0 42482 5 1 1 42481
0 42483 7 1 2 73335 42482
0 42484 7 1 2 42480 42483
0 42485 5 1 1 42484
0 42486 7 1 2 58454 42485
0 42487 5 1 1 42486
0 42488 7 1 2 42478 42487
0 42489 7 1 2 42474 42488
0 42490 5 1 1 42489
0 42491 7 1 2 79243 42490
0 42492 5 1 1 42491
0 42493 7 1 2 59457 71804
0 42494 5 1 1 42493
0 42495 7 1 2 71358 42494
0 42496 5 1 1 42495
0 42497 7 1 2 57682 76302
0 42498 5 1 1 42497
0 42499 7 1 2 52012 70219
0 42500 5 1 1 42499
0 42501 7 1 2 61825 79265
0 42502 7 1 2 42500 42501
0 42503 5 1 1 42502
0 42504 7 1 2 55957 42503
0 42505 5 1 1 42504
0 42506 7 1 2 42498 42505
0 42507 5 1 1 42506
0 42508 7 1 2 72425 42507
0 42509 5 1 1 42508
0 42510 7 1 2 42496 42509
0 42511 5 1 1 42510
0 42512 7 1 2 50548 42511
0 42513 5 1 1 42512
0 42514 7 1 2 73262 10358
0 42515 5 1 1 42514
0 42516 7 1 2 59869 42515
0 42517 5 1 1 42516
0 42518 7 1 2 73374 69932
0 42519 5 1 1 42518
0 42520 7 1 2 50112 69766
0 42521 7 1 2 74946 42520
0 42522 5 1 1 42521
0 42523 7 1 2 42519 42522
0 42524 7 1 2 42517 42523
0 42525 5 1 1 42524
0 42526 7 1 2 52013 42525
0 42527 5 1 1 42526
0 42528 7 1 2 70406 71355
0 42529 5 1 1 42528
0 42530 7 1 2 42527 42529
0 42531 5 1 1 42530
0 42532 7 1 2 50301 42531
0 42533 5 1 1 42532
0 42534 7 1 2 61618 77522
0 42535 5 1 1 42534
0 42536 7 1 2 70465 71387
0 42537 5 1 1 42536
0 42538 7 1 2 42535 42537
0 42539 5 1 1 42538
0 42540 7 1 2 74651 42539
0 42541 5 1 1 42540
0 42542 7 1 2 70502 71051
0 42543 5 1 1 42542
0 42544 7 1 2 58455 42543
0 42545 5 1 1 42544
0 42546 7 1 2 59082 75367
0 42547 5 1 1 42546
0 42548 7 1 2 75370 42547
0 42549 5 1 1 42548
0 42550 7 1 2 42545 42549
0 42551 5 1 1 42550
0 42552 7 1 2 71356 42551
0 42553 5 1 1 42552
0 42554 7 1 2 42541 42553
0 42555 7 1 2 42533 42554
0 42556 7 1 2 42513 42555
0 42557 5 1 1 42556
0 42558 7 1 2 73327 77985
0 42559 5 5 1 42558
0 42560 7 1 2 42557 79272
0 42561 5 1 1 42560
0 42562 7 1 2 42492 42561
0 42563 7 1 2 42464 42562
0 42564 5 1 1 42563
0 42565 7 1 2 52459 42564
0 42566 5 1 1 42565
0 42567 7 1 2 42419 42566
0 42568 5 1 1 42567
0 42569 7 1 2 53255 42568
0 42570 5 1 1 42569
0 42571 7 1 2 59810 62118
0 42572 7 1 2 63127 42571
0 42573 5 1 1 42572
0 42574 7 1 2 50302 42573
0 42575 5 1 1 42574
0 42576 7 1 2 70709 42575
0 42577 5 1 1 42576
0 42578 7 1 2 53019 42577
0 42579 5 1 1 42578
0 42580 7 1 2 61190 70231
0 42581 5 1 1 42580
0 42582 7 1 2 62119 75378
0 42583 5 1 1 42582
0 42584 7 1 2 50549 42583
0 42585 5 1 1 42584
0 42586 7 1 2 60439 42585
0 42587 7 1 2 42581 42586
0 42588 7 1 2 42579 42587
0 42589 5 1 1 42588
0 42590 7 1 2 51158 42589
0 42591 5 1 1 42590
0 42592 7 1 2 61637 70505
0 42593 5 1 1 42592
0 42594 7 1 2 52338 42593
0 42595 5 1 1 42594
0 42596 7 1 2 60255 61622
0 42597 5 1 1 42596
0 42598 7 1 2 52014 42597
0 42599 5 1 1 42598
0 42600 7 1 2 70270 42599
0 42601 7 1 2 42595 42600
0 42602 5 1 1 42601
0 42603 7 1 2 51159 42602
0 42604 5 1 1 42603
0 42605 7 1 2 54801 14738
0 42606 5 3 1 42605
0 42607 7 1 2 65940 79277
0 42608 5 1 1 42607
0 42609 7 1 2 10170 42608
0 42610 5 1 1 42609
0 42611 7 1 2 52015 60480
0 42612 7 1 2 42610 42611
0 42613 5 1 1 42612
0 42614 7 1 2 42604 42613
0 42615 5 1 1 42614
0 42616 7 1 2 58456 42615
0 42617 5 1 1 42616
0 42618 7 1 2 60156 72762
0 42619 5 1 1 42618
0 42620 7 1 2 60272 65231
0 42621 5 1 1 42620
0 42622 7 1 2 55138 42621
0 42623 5 1 1 42622
0 42624 7 1 2 77772 42623
0 42625 5 1 1 42624
0 42626 7 1 2 42619 42625
0 42627 5 1 1 42626
0 42628 7 1 2 50550 42627
0 42629 5 1 1 42628
0 42630 7 1 2 52460 79200
0 42631 5 1 1 42630
0 42632 7 1 2 42629 42631
0 42633 5 1 1 42632
0 42634 7 1 2 53020 42633
0 42635 5 1 1 42634
0 42636 7 1 2 42617 42635
0 42637 7 1 2 42591 42636
0 42638 5 1 1 42637
0 42639 7 1 2 55412 42638
0 42640 5 1 1 42639
0 42641 7 1 2 42640 40816
0 42642 5 1 1 42641
0 42643 7 1 2 62986 42642
0 42644 5 1 1 42643
0 42645 7 1 2 50551 72977
0 42646 5 1 1 42645
0 42647 7 1 2 65225 42646
0 42648 5 1 1 42647
0 42649 7 1 2 61533 42648
0 42650 5 1 1 42649
0 42651 7 1 2 50865 59664
0 42652 5 1 1 42651
0 42653 7 1 2 42650 42652
0 42654 7 1 2 73186 42653
0 42655 5 1 1 42654
0 42656 7 1 2 52198 42655
0 42657 5 1 1 42656
0 42658 7 1 2 59908 73179
0 42659 7 1 2 42657 42658
0 42660 5 1 1 42659
0 42661 7 1 2 58457 42660
0 42662 5 1 1 42661
0 42663 7 1 2 61191 61455
0 42664 5 1 1 42663
0 42665 7 1 2 59771 42664
0 42666 5 1 1 42665
0 42667 7 1 2 50866 42666
0 42668 5 1 1 42667
0 42669 7 1 2 54802 30101
0 42670 5 1 1 42669
0 42671 7 1 2 52199 64956
0 42672 7 1 2 42670 42671
0 42673 5 1 1 42672
0 42674 7 1 2 61511 70895
0 42675 5 1 1 42674
0 42676 7 1 2 62243 42675
0 42677 5 1 1 42676
0 42678 7 1 2 50867 60712
0 42679 5 1 1 42678
0 42680 7 1 2 42677 42679
0 42681 7 1 2 42673 42680
0 42682 5 1 1 42681
0 42683 7 1 2 50552 42682
0 42684 5 1 1 42683
0 42685 7 1 2 55139 42684
0 42686 7 1 2 42668 42685
0 42687 5 1 1 42686
0 42688 7 1 2 53021 42687
0 42689 5 1 1 42688
0 42690 7 1 2 52200 60733
0 42691 5 1 1 42690
0 42692 7 1 2 60501 42691
0 42693 5 1 1 42692
0 42694 7 2 2 52016 42693
0 42695 5 2 1 79280
0 42696 7 1 2 57683 79281
0 42697 5 1 1 42696
0 42698 7 1 2 55958 65810
0 42699 5 1 1 42698
0 42700 7 1 2 55140 42699
0 42701 7 1 2 42697 42700
0 42702 5 1 1 42701
0 42703 7 1 2 50868 42702
0 42704 5 1 1 42703
0 42705 7 1 2 65232 60872
0 42706 5 1 1 42705
0 42707 7 1 2 48267 78156
0 42708 5 1 1 42707
0 42709 7 1 2 51160 42708
0 42710 5 1 1 42709
0 42711 7 1 2 42706 42710
0 42712 7 1 2 42704 42711
0 42713 7 1 2 42689 42712
0 42714 7 1 2 42662 42713
0 42715 5 2 1 42714
0 42716 7 1 2 68594 79284
0 42717 5 1 1 42716
0 42718 7 1 2 76421 42717
0 42719 7 1 2 42644 42718
0 42720 5 1 1 42719
0 42721 7 1 2 73318 42720
0 42722 5 1 1 42721
0 42723 7 1 2 63490 77979
0 42724 7 1 2 79285 42723
0 42725 5 1 1 42724
0 42726 7 1 2 51639 42725
0 42727 7 1 2 42722 42726
0 42728 7 1 2 42570 42727
0 42729 5 1 1 42728
0 42730 7 2 2 42341 42729
0 42731 7 1 2 51779 79286
0 42732 5 1 1 42731
0 42733 7 1 2 75124 77044
0 42734 5 2 1 42733
0 42735 7 1 2 65158 77007
0 42736 5 1 1 42735
0 42737 7 1 2 79288 42736
0 42738 5 1 1 42737
0 42739 7 1 2 51640 42738
0 42740 5 1 1 42739
0 42741 7 2 2 66297 77115
0 42742 7 1 2 62499 79290
0 42743 5 1 1 42742
0 42744 7 1 2 42740 42743
0 42745 5 2 1 42744
0 42746 7 1 2 49971 79292
0 42747 5 1 1 42746
0 42748 7 1 2 68835 79291
0 42749 5 1 1 42748
0 42750 7 1 2 42747 42749
0 42751 5 1 1 42750
0 42752 7 1 2 51431 42751
0 42753 5 1 1 42752
0 42754 7 1 2 71474 77595
0 42755 5 1 1 42754
0 42756 7 1 2 74995 42755
0 42757 5 1 1 42756
0 42758 7 2 2 66487 42757
0 42759 5 1 1 79294
0 42760 7 1 2 42753 42759
0 42761 5 1 1 42760
0 42762 7 1 2 52824 42761
0 42763 5 1 1 42762
0 42764 7 1 2 53740 79293
0 42765 5 1 1 42764
0 42766 7 2 2 50303 77045
0 42767 7 3 2 62500 67788
0 42768 7 1 2 79296 79298
0 42769 5 1 1 42768
0 42770 7 1 2 42765 42769
0 42771 5 1 1 42770
0 42772 7 1 2 48972 42771
0 42773 5 1 1 42772
0 42774 7 1 2 71823 79299
0 42775 7 1 2 77008 42774
0 42776 5 1 1 42775
0 42777 7 1 2 42773 42776
0 42778 5 1 1 42777
0 42779 7 1 2 51432 42778
0 42780 5 1 1 42779
0 42781 7 1 2 42763 42780
0 42782 5 1 1 42781
0 42783 7 1 2 51780 42782
0 42784 5 1 1 42783
0 42785 7 1 2 52201 74186
0 42786 7 1 2 77980 42785
0 42787 5 1 1 42786
0 42788 7 1 2 60602 59006
0 42789 7 1 2 79157 42788
0 42790 5 1 1 42789
0 42791 7 1 2 42787 42790
0 42792 5 1 1 42791
0 42793 7 1 2 51433 42792
0 42794 5 1 1 42793
0 42795 7 3 2 61914 73677
0 42796 7 1 2 69911 79301
0 42797 5 1 1 42796
0 42798 7 2 2 50869 62987
0 42799 7 2 2 52339 75096
0 42800 7 1 2 53584 78614
0 42801 7 1 2 79306 42800
0 42802 5 1 1 42801
0 42803 7 1 2 66000 42802
0 42804 5 1 1 42803
0 42805 7 1 2 79304 42804
0 42806 5 1 1 42805
0 42807 7 1 2 42797 42806
0 42808 5 1 1 42807
0 42809 7 1 2 73319 42808
0 42810 5 1 1 42809
0 42811 7 1 2 42794 42810
0 42812 5 1 1 42811
0 42813 7 1 2 51781 42812
0 42814 5 1 1 42813
0 42815 7 3 2 50870 69912
0 42816 7 2 2 70486 79308
0 42817 7 1 2 49972 79311
0 42818 5 1 1 42817
0 42819 7 2 2 66427 76736
0 42820 7 1 2 70010 79313
0 42821 5 1 1 42820
0 42822 7 1 2 42818 42821
0 42823 5 1 1 42822
0 42824 7 1 2 51782 42823
0 42825 5 1 1 42824
0 42826 7 5 2 62501 69532
0 42827 7 1 2 72533 79315
0 42828 5 1 1 42827
0 42829 7 1 2 42825 42828
0 42830 5 2 1 42829
0 42831 7 1 2 51161 60030
0 42832 7 1 2 79320 42831
0 42833 5 1 1 42832
0 42834 7 1 2 42814 42833
0 42835 5 1 1 42834
0 42836 7 1 2 53022 42835
0 42837 5 1 1 42836
0 42838 7 2 2 54803 79253
0 42839 7 1 2 60603 79322
0 42840 5 1 1 42839
0 42841 7 1 2 68605 42840
0 42842 5 1 1 42841
0 42843 7 1 2 53741 42842
0 42844 5 1 1 42843
0 42845 7 1 2 79221 42844
0 42846 5 1 1 42845
0 42847 7 1 2 66298 42846
0 42848 5 1 1 42847
0 42849 7 2 2 52017 75125
0 42850 5 2 1 79324
0 42851 7 1 2 61915 73782
0 42852 5 1 1 42851
0 42853 7 1 2 79326 42852
0 42854 5 1 1 42853
0 42855 7 1 2 78725 42854
0 42856 5 1 1 42855
0 42857 7 1 2 42848 42856
0 42858 5 1 1 42857
0 42859 7 1 2 52825 42858
0 42860 5 1 1 42859
0 42861 7 1 2 59946 78826
0 42862 5 1 1 42861
0 42863 7 1 2 66624 76980
0 42864 5 1 1 42863
0 42865 7 1 2 42862 42864
0 42866 5 1 1 42865
0 42867 7 1 2 51641 42866
0 42868 5 1 1 42867
0 42869 7 1 2 74440 75097
0 42870 5 1 1 42869
0 42871 7 1 2 42868 42870
0 42872 5 1 1 42871
0 42873 7 1 2 48973 42872
0 42874 5 1 1 42873
0 42875 7 1 2 52340 74187
0 42876 7 1 2 77981 42875
0 42877 5 1 1 42876
0 42878 7 1 2 42874 42877
0 42879 5 1 1 42878
0 42880 7 1 2 51434 42879
0 42881 5 1 1 42880
0 42882 7 1 2 42860 42881
0 42883 5 1 1 42882
0 42884 7 1 2 51783 42883
0 42885 5 1 1 42884
0 42886 7 1 2 42837 42885
0 42887 5 1 1 42886
0 42888 7 1 2 58458 42887
0 42889 5 1 1 42888
0 42890 7 2 2 71475 74206
0 42891 7 1 2 62429 69533
0 42892 7 1 2 79328 42891
0 42893 5 1 1 42892
0 42894 7 1 2 65738 73492
0 42895 5 1 1 42894
0 42896 7 1 2 52720 73731
0 42897 5 1 1 42896
0 42898 7 1 2 42895 42897
0 42899 5 1 1 42898
0 42900 7 1 2 49813 42899
0 42901 5 1 1 42900
0 42902 7 1 2 67860 79307
0 42903 5 1 1 42902
0 42904 7 1 2 51162 72354
0 42905 5 1 1 42904
0 42906 7 1 2 42903 42905
0 42907 5 1 1 42906
0 42908 7 1 2 53585 42907
0 42909 5 1 1 42908
0 42910 7 1 2 42901 42909
0 42911 5 2 1 42910
0 42912 7 1 2 51435 71236
0 42913 7 1 2 79330 42912
0 42914 5 1 1 42913
0 42915 7 1 2 42893 42914
0 42916 5 1 1 42915
0 42917 7 1 2 51784 42916
0 42918 5 1 1 42917
0 42919 7 2 2 68987 79309
0 42920 7 2 2 53586 73648
0 42921 7 1 2 56664 79334
0 42922 7 1 2 79332 42921
0 42923 5 1 1 42922
0 42924 7 1 2 42918 42923
0 42925 5 1 1 42924
0 42926 7 1 2 60669 42925
0 42927 5 1 1 42926
0 42928 7 1 2 50871 79245
0 42929 5 1 1 42928
0 42930 7 2 2 48443 76925
0 42931 5 1 1 79336
0 42932 7 1 2 71359 79273
0 42933 7 1 2 42931 42932
0 42934 5 1 1 42933
0 42935 7 1 2 42929 42934
0 42936 5 1 1 42935
0 42937 7 1 2 51642 42936
0 42938 5 1 1 42937
0 42939 7 1 2 66104 77597
0 42940 7 1 2 79224 42939
0 42941 5 1 1 42940
0 42942 7 1 2 42938 42941
0 42943 5 1 1 42942
0 42944 7 1 2 51785 42943
0 42945 5 1 1 42944
0 42946 7 2 2 60607 60719
0 42947 5 1 1 79338
0 42948 7 1 2 51163 42947
0 42949 7 1 2 79321 42948
0 42950 5 1 1 42949
0 42951 7 1 2 42945 42950
0 42952 5 1 1 42951
0 42953 7 1 2 53023 42952
0 42954 5 1 1 42953
0 42955 7 1 2 42927 42954
0 42956 7 1 2 42889 42955
0 42957 7 1 2 42784 42956
0 42958 5 1 1 42957
0 42959 7 1 2 53132 42958
0 42960 5 1 1 42959
0 42961 7 1 2 61249 79323
0 42962 5 1 1 42961
0 42963 7 1 2 68606 42962
0 42964 5 1 1 42963
0 42965 7 1 2 53742 42964
0 42966 5 1 1 42965
0 42967 7 1 2 79222 42966
0 42968 5 1 1 42967
0 42969 7 1 2 52826 42968
0 42970 5 1 1 42969
0 42971 7 2 2 52721 63424
0 42972 5 1 1 79340
0 42973 7 1 2 69287 79341
0 42974 5 1 1 42973
0 42975 7 1 2 42970 42974
0 42976 5 1 1 42975
0 42977 7 2 2 66299 42976
0 42978 5 1 1 79342
0 42979 7 1 2 50872 79236
0 42980 5 1 1 42979
0 42981 7 1 2 73508 79302
0 42982 5 1 1 42981
0 42983 7 1 2 42980 42982
0 42984 5 1 1 42983
0 42985 7 1 2 49973 42984
0 42986 5 1 1 42985
0 42987 7 1 2 55413 79305
0 42988 5 1 1 42987
0 42989 7 1 2 65159 73375
0 42990 5 1 1 42989
0 42991 7 1 2 42988 42990
0 42992 5 1 1 42991
0 42993 7 1 2 67125 42992
0 42994 5 1 1 42993
0 42995 7 1 2 42986 42994
0 42996 5 1 1 42995
0 42997 7 1 2 53024 42996
0 42998 5 1 1 42997
0 42999 7 2 2 67535 78573
0 43000 5 1 1 79344
0 43001 7 1 2 52018 79345
0 43002 5 1 1 43001
0 43003 7 1 2 42998 43002
0 43004 5 2 1 43003
0 43005 7 1 2 51643 79346
0 43006 5 1 1 43005
0 43007 7 1 2 42978 43006
0 43008 5 1 1 43007
0 43009 7 1 2 52341 43008
0 43010 5 1 1 43009
0 43011 7 2 2 66221 74244
0 43012 5 1 1 79348
0 43013 7 2 2 71155 74821
0 43014 5 1 1 79350
0 43015 7 1 2 48829 43014
0 43016 5 1 1 43015
0 43017 7 1 2 65994 71156
0 43018 5 1 1 43017
0 43019 7 1 2 25310 43018
0 43020 5 2 1 43019
0 43021 7 1 2 67861 79352
0 43022 7 1 2 43016 43021
0 43023 5 1 1 43022
0 43024 7 1 2 43012 43023
0 43025 5 1 1 43024
0 43026 7 1 2 59947 43025
0 43027 5 1 1 43026
0 43028 7 3 2 53587 63844
0 43029 5 2 1 79354
0 43030 7 1 2 77605 79357
0 43031 5 1 1 43030
0 43032 7 1 2 69534 75098
0 43033 7 1 2 43031 43032
0 43034 5 1 1 43033
0 43035 7 2 2 43027 43034
0 43036 5 1 1 79359
0 43037 7 1 2 43010 79360
0 43038 5 1 1 43037
0 43039 7 1 2 51786 43038
0 43040 5 1 1 43039
0 43041 7 1 2 52019 71301
0 43042 7 2 2 69813 43041
0 43043 7 1 2 53025 69535
0 43044 7 1 2 71596 43043
0 43045 7 1 2 79361 43044
0 43046 5 1 1 43045
0 43047 7 1 2 43040 43046
0 43048 5 1 1 43047
0 43049 7 1 2 58459 43048
0 43050 5 1 1 43049
0 43051 7 1 2 69814 77532
0 43052 7 1 2 77538 79316
0 43053 7 2 2 43051 43052
0 43054 5 1 1 79363
0 43055 7 1 2 43050 43054
0 43056 7 1 2 42960 43055
0 43057 5 1 1 43056
0 43058 7 1 2 50553 43057
0 43059 5 1 1 43058
0 43060 7 2 2 61048 71824
0 43061 5 1 1 79365
0 43062 7 1 2 75126 43061
0 43063 5 2 1 43062
0 43064 7 1 2 61192 79367
0 43065 5 1 1 43064
0 43066 7 1 2 61916 75884
0 43067 7 1 2 76868 43066
0 43068 5 1 1 43067
0 43069 7 1 2 43065 43068
0 43070 5 1 1 43069
0 43071 7 1 2 51436 43070
0 43072 5 1 1 43071
0 43073 7 2 2 55414 78432
0 43074 7 1 2 73444 79369
0 43075 5 1 1 43074
0 43076 7 1 2 43072 43075
0 43077 5 1 1 43076
0 43078 7 1 2 53743 43077
0 43079 5 1 1 43078
0 43080 7 1 2 70789 78792
0 43081 5 1 1 43080
0 43082 7 1 2 43079 43081
0 43083 5 1 1 43082
0 43084 7 1 2 66400 43083
0 43085 5 1 1 43084
0 43086 7 1 2 48010 62330
0 43087 5 1 1 43086
0 43088 7 1 2 51437 43087
0 43089 7 1 2 70579 43088
0 43090 5 1 1 43089
0 43091 7 1 2 59030 69536
0 43092 7 1 2 7741 43091
0 43093 7 1 2 72668 43092
0 43094 5 1 1 43093
0 43095 7 1 2 43090 43094
0 43096 5 1 1 43095
0 43097 7 1 2 55572 43096
0 43098 5 1 1 43097
0 43099 7 2 2 55713 68776
0 43100 7 1 2 69913 74889
0 43101 7 1 2 79371 43100
0 43102 5 1 1 43101
0 43103 7 1 2 43098 43102
0 43104 5 1 1 43103
0 43105 7 1 2 51164 43104
0 43106 5 1 1 43105
0 43107 7 3 2 53744 75181
0 43108 7 1 2 71665 79373
0 43109 5 1 1 43108
0 43110 7 1 2 67862 79370
0 43111 5 1 1 43110
0 43112 7 1 2 74317 71388
0 43113 7 1 2 76922 43112
0 43114 5 1 1 43113
0 43115 7 1 2 43111 43114
0 43116 5 1 1 43115
0 43117 7 1 2 53026 43116
0 43118 5 1 1 43117
0 43119 7 1 2 61193 72957
0 43120 5 1 1 43119
0 43121 7 1 2 74837 79303
0 43122 5 1 1 43121
0 43123 7 1 2 43120 43122
0 43124 5 1 1 43123
0 43125 7 1 2 73349 43124
0 43126 5 1 1 43125
0 43127 7 1 2 43118 43126
0 43128 5 1 1 43127
0 43129 7 1 2 51644 43128
0 43130 5 1 1 43129
0 43131 7 1 2 43109 43130
0 43132 7 1 2 43106 43131
0 43133 5 1 1 43132
0 43134 7 1 2 52722 43133
0 43135 5 1 1 43134
0 43136 7 1 2 67789 68595
0 43137 5 2 1 43136
0 43138 7 1 2 51165 77593
0 43139 7 1 2 66433 43138
0 43140 7 1 2 75996 43139
0 43141 5 1 1 43140
0 43142 7 1 2 79376 43141
0 43143 5 1 1 43142
0 43144 7 1 2 52202 43143
0 43145 5 1 1 43144
0 43146 7 4 2 55573 68981
0 43147 5 1 1 79378
0 43148 7 1 2 55714 67790
0 43149 5 1 1 43148
0 43150 7 1 2 43147 43149
0 43151 5 1 1 43150
0 43152 7 1 2 68596 43151
0 43153 5 1 1 43152
0 43154 7 1 2 43145 43153
0 43155 5 1 1 43154
0 43156 7 1 2 50304 43155
0 43157 5 1 1 43156
0 43158 7 1 2 49974 79351
0 43159 5 1 1 43158
0 43160 7 1 2 65739 72172
0 43161 5 1 1 43160
0 43162 7 1 2 43159 43161
0 43163 5 1 1 43162
0 43164 7 1 2 59560 43163
0 43165 5 1 1 43164
0 43166 7 1 2 51645 63746
0 43167 7 1 2 72968 68350
0 43168 7 1 2 43166 43167
0 43169 7 1 2 61473 43168
0 43170 5 1 1 43169
0 43171 7 1 2 43165 43170
0 43172 7 1 2 43157 43171
0 43173 5 1 1 43172
0 43174 7 1 2 52827 43173
0 43175 5 1 1 43174
0 43176 7 1 2 43135 43175
0 43177 7 1 2 43085 43176
0 43178 5 1 1 43177
0 43179 7 1 2 52342 43178
0 43180 5 1 1 43179
0 43181 7 1 2 22495 79358
0 43182 5 1 1 43181
0 43183 7 1 2 59561 43182
0 43184 5 1 1 43183
0 43185 7 1 2 62690 70317
0 43186 5 1 1 43185
0 43187 7 1 2 78718 43186
0 43188 7 1 2 43184 43187
0 43189 5 1 1 43188
0 43190 7 1 2 78739 43189
0 43191 5 1 1 43190
0 43192 7 1 2 70450 79353
0 43193 5 1 1 43192
0 43194 7 1 2 11124 43193
0 43195 5 1 1 43194
0 43196 7 1 2 73320 43195
0 43197 5 1 1 43196
0 43198 7 1 2 72590 79310
0 43199 5 1 1 43198
0 43200 7 1 2 43197 43199
0 43201 7 1 2 43191 43200
0 43202 5 1 1 43201
0 43203 7 1 2 52723 43202
0 43204 5 1 1 43203
0 43205 7 1 2 60713 79349
0 43206 5 1 1 43205
0 43207 7 11 2 51646 67863
0 43208 7 1 2 55141 21142
0 43209 5 2 1 43208
0 43210 7 1 2 69811 79393
0 43211 5 1 1 43210
0 43212 7 1 2 14530 43211
0 43213 5 1 1 43212
0 43214 7 1 2 79382 43213
0 43215 5 1 1 43214
0 43216 7 1 2 43206 43215
0 43217 7 2 2 43204 43216
0 43218 5 1 1 79395
0 43219 7 1 2 43180 79396
0 43220 5 1 1 43219
0 43221 7 1 2 50554 43220
0 43222 5 1 1 43221
0 43223 7 1 2 77533 76488
0 43224 5 1 1 43223
0 43225 7 1 2 48974 43224
0 43226 5 1 1 43225
0 43227 7 1 2 49814 43226
0 43228 5 1 1 43227
0 43229 7 1 2 60488 71229
0 43230 5 1 1 43229
0 43231 7 1 2 48830 43230
0 43232 5 1 1 43231
0 43233 7 1 2 63425 43232
0 43234 5 1 1 43233
0 43235 7 1 2 43228 43234
0 43236 5 1 1 43235
0 43237 7 1 2 50873 43236
0 43238 5 1 1 43237
0 43239 7 3 2 64389 67569
0 43240 7 1 2 59790 63124
0 43241 7 1 2 79397 43240
0 43242 5 1 1 43241
0 43243 7 1 2 43238 43242
0 43244 5 1 1 43243
0 43245 7 1 2 52020 43244
0 43246 5 1 1 43245
0 43247 7 1 2 59014 42972
0 43248 5 4 1 43247
0 43249 7 1 2 50874 79400
0 43250 5 2 1 43249
0 43251 7 1 2 71002 79398
0 43252 5 1 1 43251
0 43253 7 1 2 79404 43252
0 43254 5 1 1 43253
0 43255 7 1 2 57265 43254
0 43256 5 1 1 43255
0 43257 7 1 2 43246 43256
0 43258 5 1 1 43257
0 43259 7 1 2 50305 43258
0 43260 5 1 1 43259
0 43261 7 1 2 13429 79401
0 43262 5 1 1 43261
0 43263 7 1 2 71440 79399
0 43264 5 1 1 43263
0 43265 7 1 2 79405 43264
0 43266 5 1 1 43265
0 43267 7 1 2 52343 43266
0 43268 5 1 1 43267
0 43269 7 1 2 43262 43268
0 43270 7 1 2 43260 43269
0 43271 5 1 1 43270
0 43272 7 1 2 49975 43271
0 43273 5 1 1 43272
0 43274 7 1 2 73678 75865
0 43275 5 1 1 43274
0 43276 7 1 2 58809 43275
0 43277 5 2 1 43276
0 43278 7 1 2 70497 79406
0 43279 5 1 1 43278
0 43280 7 1 2 67570 71441
0 43281 5 1 1 43280
0 43282 7 1 2 58810 43281
0 43283 5 2 1 43282
0 43284 7 1 2 60031 79408
0 43285 5 1 1 43284
0 43286 7 1 2 54412 73532
0 43287 7 1 2 72970 43286
0 43288 5 1 1 43287
0 43289 7 1 2 58811 43288
0 43290 5 1 1 43289
0 43291 7 1 2 60050 43290
0 43292 5 1 1 43291
0 43293 7 1 2 62692 43292
0 43294 7 1 2 43285 43293
0 43295 7 1 2 43279 43294
0 43296 5 1 1 43295
0 43297 7 1 2 67126 43296
0 43298 5 1 1 43297
0 43299 7 1 2 51647 43298
0 43300 7 1 2 43273 43299
0 43301 5 1 1 43300
0 43302 7 4 2 51166 79225
0 43303 7 1 2 59754 61176
0 43304 5 1 1 43303
0 43305 7 1 2 71298 43304
0 43306 5 1 1 43305
0 43307 7 1 2 59746 60647
0 43308 5 2 1 43307
0 43309 7 1 2 43306 79414
0 43310 5 1 1 43309
0 43311 7 1 2 79410 43310
0 43312 5 1 1 43311
0 43313 7 3 2 68836 73649
0 43314 5 1 1 79416
0 43315 7 1 2 55574 43314
0 43316 7 1 2 43312 43315
0 43317 5 1 1 43316
0 43318 7 1 2 51438 43317
0 43319 7 1 2 43301 43318
0 43320 5 1 1 43319
0 43321 7 2 2 62502 72411
0 43322 5 1 1 79419
0 43323 7 2 2 66768 79420
0 43324 5 2 1 79421
0 43325 7 3 2 51648 62988
0 43326 7 2 2 67864 79425
0 43327 7 1 2 78008 79428
0 43328 5 1 1 43327
0 43329 7 1 2 79423 43328
0 43330 5 1 1 43329
0 43331 7 1 2 60273 43330
0 43332 5 1 1 43331
0 43333 7 1 2 75333 79429
0 43334 5 1 1 43333
0 43335 7 1 2 73398 69780
0 43336 5 1 1 43335
0 43337 7 1 2 74996 43336
0 43338 5 1 1 43337
0 43339 7 2 2 57684 78740
0 43340 7 1 2 43338 79430
0 43341 5 1 1 43340
0 43342 7 1 2 43334 43341
0 43343 5 1 1 43342
0 43344 7 1 2 52021 43343
0 43345 5 1 1 43344
0 43346 7 1 2 43332 43345
0 43347 5 1 1 43346
0 43348 7 1 2 55415 43347
0 43349 5 1 1 43348
0 43350 7 1 2 61641 66300
0 43351 7 1 2 79226 43350
0 43352 5 1 1 43351
0 43353 7 1 2 68557 79274
0 43354 7 1 2 77273 43353
0 43355 5 1 1 43354
0 43356 7 1 2 43352 43355
0 43357 5 1 1 43356
0 43358 7 1 2 52344 43357
0 43359 5 1 1 43358
0 43360 7 1 2 61616 72530
0 43361 7 1 2 78574 43360
0 43362 5 1 1 43361
0 43363 7 1 2 43359 43362
0 43364 5 1 1 43363
0 43365 7 1 2 51439 43364
0 43366 5 1 1 43365
0 43367 7 2 2 55575 70376
0 43368 7 1 2 71371 79417
0 43369 7 1 2 79432 43368
0 43370 5 1 1 43369
0 43371 7 1 2 43366 43370
0 43372 7 1 2 43349 43371
0 43373 5 1 1 43372
0 43374 7 1 2 58460 43373
0 43375 5 1 1 43374
0 43376 7 1 2 69513 71483
0 43377 5 1 1 43376
0 43378 7 1 2 73614 76555
0 43379 5 1 1 43378
0 43380 7 1 2 43377 43379
0 43381 5 1 1 43380
0 43382 7 1 2 79379 43381
0 43383 5 1 1 43382
0 43384 7 1 2 79377 43383
0 43385 5 1 1 43384
0 43386 7 1 2 52828 43385
0 43387 5 1 1 43386
0 43388 7 1 2 48975 69914
0 43389 7 1 2 78827 43388
0 43390 5 1 1 43389
0 43391 7 1 2 43387 43390
0 43392 5 1 1 43391
0 43393 7 1 2 70420 43392
0 43394 5 1 1 43393
0 43395 7 1 2 73057 73555
0 43396 7 1 2 74963 43395
0 43397 7 1 2 79275 43396
0 43398 5 1 1 43397
0 43399 7 1 2 43394 43398
0 43400 5 1 1 43399
0 43401 7 1 2 59870 43400
0 43402 5 1 1 43401
0 43403 7 1 2 52909 73163
0 43404 7 1 2 76764 43403
0 43405 7 2 2 79380 43404
0 43406 5 1 1 79434
0 43407 7 1 2 61632 79435
0 43408 5 1 1 43407
0 43409 7 1 2 48268 21154
0 43410 5 1 1 43409
0 43411 7 1 2 50875 60019
0 43412 7 1 2 79383 43411
0 43413 7 1 2 43410 43412
0 43414 5 1 1 43413
0 43415 7 1 2 43408 43414
0 43416 5 1 1 43415
0 43417 7 1 2 60481 43416
0 43418 5 1 1 43417
0 43419 7 1 2 59922 72412
0 43420 7 1 2 67439 71171
0 43421 7 1 2 43419 43420
0 43422 5 1 1 43421
0 43423 7 1 2 51167 75392
0 43424 5 1 1 43423
0 43425 7 1 2 57544 43424
0 43426 5 1 1 43425
0 43427 7 1 2 65307 59781
0 43428 5 1 1 43427
0 43429 7 1 2 55142 43428
0 43430 5 2 1 43429
0 43431 7 1 2 79384 79436
0 43432 7 1 2 43426 43431
0 43433 5 1 1 43432
0 43434 7 1 2 43422 43433
0 43435 7 1 2 43418 43434
0 43436 5 1 1 43435
0 43437 7 1 2 62989 43436
0 43438 5 1 1 43437
0 43439 7 1 2 63754 79202
0 43440 5 1 1 43439
0 43441 7 1 2 79422 43440
0 43442 5 1 1 43441
0 43443 7 1 2 43438 43442
0 43444 5 1 1 43443
0 43445 7 1 2 55416 43444
0 43446 5 1 1 43445
0 43447 7 1 2 52022 70909
0 43448 5 1 1 43447
0 43449 7 1 2 59113 43448
0 43450 5 1 1 43449
0 43451 7 3 2 68437 79418
0 43452 5 1 1 79438
0 43453 7 1 2 63232 79439
0 43454 7 1 2 43450 43453
0 43455 5 1 1 43454
0 43456 7 1 2 43446 43455
0 43457 7 1 2 43402 43456
0 43458 7 1 2 43375 43457
0 43459 7 1 2 43320 43458
0 43460 7 1 2 43222 43459
0 43461 5 1 1 43460
0 43462 7 1 2 51787 43461
0 43463 5 1 1 43462
0 43464 7 2 2 51788 79440
0 43465 5 1 1 79441
0 43466 7 1 2 66105 79411
0 43467 5 1 1 43466
0 43468 7 1 2 79234 42400
0 43469 5 1 1 43468
0 43470 7 1 2 49976 43469
0 43471 5 1 1 43470
0 43472 7 1 2 79249 43471
0 43473 5 1 1 43472
0 43474 7 1 2 51649 71157
0 43475 7 1 2 43473 43474
0 43476 5 1 1 43475
0 43477 7 1 2 43467 43476
0 43478 5 2 1 43477
0 43479 7 1 2 51789 79443
0 43480 5 1 1 43479
0 43481 7 1 2 60482 79335
0 43482 7 1 2 79333 43481
0 43483 5 1 1 43482
0 43484 7 1 2 43480 43483
0 43485 5 1 1 43484
0 43486 7 1 2 52203 43485
0 43487 5 1 1 43486
0 43488 7 1 2 43465 43487
0 43489 5 1 1 43488
0 43490 7 1 2 50306 74571
0 43491 5 1 1 43490
0 43492 7 1 2 70983 43491
0 43493 5 3 1 43492
0 43494 7 1 2 43489 79445
0 43495 5 1 1 43494
0 43496 7 3 2 69815 79374
0 43497 7 1 2 53027 58842
0 43498 7 2 2 73484 43497
0 43499 7 1 2 77539 79451
0 43500 7 1 2 79448 43499
0 43501 5 1 1 43500
0 43502 7 1 2 43495 43501
0 43503 7 1 2 43463 43502
0 43504 7 1 2 43059 43503
0 43505 5 1 1 43504
0 43506 7 1 2 57067 43505
0 43507 5 1 1 43506
0 43508 7 1 2 52023 75219
0 43509 5 1 1 43508
0 43510 7 1 2 65370 77041
0 43511 5 1 1 43510
0 43512 7 1 2 43509 43511
0 43513 5 1 1 43512
0 43514 7 1 2 52204 43513
0 43515 5 1 1 43514
0 43516 7 1 2 53133 77742
0 43517 5 1 1 43516
0 43518 7 1 2 43515 43517
0 43519 5 1 1 43518
0 43520 7 1 2 52345 43519
0 43521 5 1 1 43520
0 43522 7 1 2 62086 65941
0 43523 5 1 1 43522
0 43524 7 2 2 43521 43523
0 43525 7 1 2 52461 79269
0 43526 5 1 1 43525
0 43527 7 1 2 79453 43526
0 43528 5 1 1 43527
0 43529 7 1 2 50876 43528
0 43530 5 1 1 43529
0 43531 7 1 2 52462 79271
0 43532 5 2 1 43531
0 43533 7 1 2 43530 79455
0 43534 5 1 1 43533
0 43535 7 1 2 77626 79449
0 43536 7 2 2 43534 43535
0 43537 5 1 1 79457
0 43538 7 1 2 78044 79282
0 43539 5 1 1 43538
0 43540 7 2 2 51168 43539
0 43541 5 1 1 79459
0 43542 7 1 2 60449 77241
0 43543 5 1 1 43542
0 43544 7 1 2 43541 43543
0 43545 5 1 1 43544
0 43546 7 1 2 78429 43545
0 43547 5 1 1 43546
0 43548 7 1 2 60814 77889
0 43549 5 1 1 43548
0 43550 7 1 2 55143 43549
0 43551 5 2 1 43550
0 43552 7 1 2 65995 79461
0 43553 5 1 1 43552
0 43554 7 1 2 43547 43553
0 43555 5 1 1 43554
0 43556 7 1 2 52724 43555
0 43557 5 1 1 43556
0 43558 7 1 2 53588 25058
0 43559 5 1 1 43558
0 43560 7 1 2 60804 67691
0 43561 7 1 2 43559 43560
0 43562 5 1 1 43561
0 43563 7 1 2 75196 43562
0 43564 5 1 1 43563
0 43565 7 1 2 51650 43564
0 43566 5 1 1 43565
0 43567 7 1 2 43557 43566
0 43568 5 1 1 43567
0 43569 7 1 2 67865 43568
0 43570 5 1 1 43569
0 43571 7 1 2 66401 77982
0 43572 5 1 1 43571
0 43573 7 2 2 59007 65740
0 43574 5 2 1 79463
0 43575 7 1 2 75814 79464
0 43576 5 1 1 43575
0 43577 7 2 2 43572 43576
0 43578 5 1 1 79467
0 43579 7 1 2 60805 43578
0 43580 5 1 1 43579
0 43581 7 1 2 60256 79283
0 43582 5 3 1 43581
0 43583 7 2 2 51651 70487
0 43584 7 2 2 75815 79472
0 43585 5 1 1 79474
0 43586 7 1 2 49977 79475
0 43587 7 1 2 79469 43586
0 43588 5 1 1 43587
0 43589 7 1 2 79465 43588
0 43590 5 1 1 43589
0 43591 7 1 2 79460 43590
0 43592 5 1 1 43591
0 43593 7 1 2 43580 43592
0 43594 5 1 1 43593
0 43595 7 1 2 51440 43594
0 43596 5 1 1 43595
0 43597 7 1 2 79205 79412
0 43598 5 1 1 43597
0 43599 7 4 2 53745 73650
0 43600 5 1 1 79476
0 43601 7 1 2 79355 79477
0 43602 5 2 1 43601
0 43603 7 1 2 43598 79480
0 43604 5 1 1 43603
0 43605 7 1 2 55576 43604
0 43606 5 1 1 43605
0 43607 7 2 2 78601 79385
0 43608 7 1 2 73257 79482
0 43609 5 1 1 43608
0 43610 7 1 2 43606 43609
0 43611 5 3 1 43610
0 43612 7 1 2 60875 65796
0 43613 5 2 1 43612
0 43614 7 1 2 79484 79487
0 43615 5 1 1 43614
0 43616 7 1 2 54112 76926
0 43617 5 2 1 43616
0 43618 7 1 2 49978 79232
0 43619 5 1 1 43618
0 43620 7 1 2 79250 43619
0 43621 5 1 1 43620
0 43622 7 1 2 79489 43621
0 43623 5 1 1 43622
0 43624 7 1 2 52205 49979
0 43625 7 1 2 79240 43624
0 43626 5 1 1 43625
0 43627 7 1 2 43623 43626
0 43628 5 2 1 43627
0 43629 7 1 2 50555 79491
0 43630 5 1 1 43629
0 43631 7 1 2 62110 79255
0 43632 5 1 1 43631
0 43633 7 1 2 43630 43632
0 43634 5 1 1 43633
0 43635 7 1 2 52463 43634
0 43636 5 1 1 43635
0 43637 7 1 2 73635 78575
0 43638 5 1 1 43637
0 43639 7 1 2 51652 43638
0 43640 7 1 2 43636 43639
0 43641 5 1 1 43640
0 43642 7 1 2 55577 79481
0 43643 5 1 1 43642
0 43644 7 1 2 57685 43643
0 43645 7 1 2 43641 43644
0 43646 5 1 1 43645
0 43647 7 1 2 43615 43646
0 43648 7 1 2 43596 43647
0 43649 7 1 2 43570 43648
0 43650 5 1 1 43649
0 43651 7 1 2 51790 43650
0 43652 5 1 1 43651
0 43653 7 1 2 60157 79485
0 43654 5 1 1 43653
0 43655 7 2 2 52829 75816
0 43656 5 1 1 79493
0 43657 7 1 2 55578 43656
0 43658 5 1 1 43657
0 43659 7 1 2 59948 72194
0 43660 7 1 2 43658 43659
0 43661 5 1 1 43660
0 43662 7 1 2 10982 43661
0 43663 5 1 1 43662
0 43664 7 1 2 78828 43663
0 43665 5 1 1 43664
0 43666 7 1 2 73732 75787
0 43667 7 1 2 61456 43666
0 43668 5 1 1 43667
0 43669 7 1 2 52464 60609
0 43670 5 1 1 43669
0 43671 7 1 2 55144 43670
0 43672 5 1 1 43671
0 43673 7 1 2 68754 72137
0 43674 7 1 2 43672 43673
0 43675 5 1 1 43674
0 43676 7 1 2 43668 43675
0 43677 5 1 1 43676
0 43678 7 1 2 52725 43677
0 43679 5 1 1 43678
0 43680 7 1 2 59949 59008
0 43681 5 1 1 43680
0 43682 7 1 2 72940 77941
0 43683 7 1 2 61457 43682
0 43684 5 1 1 43683
0 43685 7 1 2 43681 43684
0 43686 5 1 1 43685
0 43687 7 1 2 67791 43686
0 43688 5 1 1 43687
0 43689 7 1 2 43679 43688
0 43690 7 1 2 43665 43689
0 43691 5 1 1 43690
0 43692 7 1 2 51441 43691
0 43693 5 1 1 43692
0 43694 7 1 2 52024 76444
0 43695 5 1 1 43694
0 43696 7 1 2 59190 43695
0 43697 5 1 1 43696
0 43698 7 1 2 79483 43697
0 43699 5 1 1 43698
0 43700 7 1 2 43693 43699
0 43701 5 2 1 43700
0 43702 7 1 2 65011 79495
0 43703 5 1 1 43702
0 43704 7 1 2 43654 43703
0 43705 5 1 1 43704
0 43706 7 1 2 51791 43705
0 43707 5 1 1 43706
0 43708 7 2 2 77942 79478
0 43709 7 1 2 72466 76459
0 43710 7 1 2 79497 43709
0 43711 7 2 2 61458 43710
0 43712 5 1 1 79499
0 43713 7 1 2 43707 43712
0 43714 5 1 1 43713
0 43715 7 1 2 58461 43714
0 43716 5 1 1 43715
0 43717 7 1 2 53134 79470
0 43718 5 1 1 43717
0 43719 7 1 2 791 43718
0 43720 5 1 1 43719
0 43721 7 1 2 52346 43720
0 43722 5 1 1 43721
0 43723 7 1 2 76969 77029
0 43724 5 1 1 43723
0 43725 7 1 2 43722 43724
0 43726 5 1 1 43725
0 43727 7 1 2 76453 79450
0 43728 7 2 2 43726 43727
0 43729 5 1 1 79501
0 43730 7 1 2 43716 43729
0 43731 7 1 2 43652 43730
0 43732 5 1 1 43731
0 43733 7 1 2 76382 43732
0 43734 5 1 1 43733
0 43735 7 1 2 43537 43734
0 43736 7 1 2 43507 43735
0 43737 7 1 2 42732 43736
0 43738 5 1 1 43737
0 43739 7 1 2 58065 43738
0 43740 5 1 1 43739
0 43741 7 1 2 65357 76748
0 43742 5 1 1 43741
0 43743 7 1 2 71468 43742
0 43744 5 1 1 43743
0 43745 7 1 2 52025 43744
0 43746 5 1 1 43745
0 43747 7 1 2 60483 78249
0 43748 5 1 1 43747
0 43749 7 1 2 71469 43748
0 43750 5 1 1 43749
0 43751 7 1 2 52206 43750
0 43752 5 1 1 43751
0 43753 7 1 2 51169 70262
0 43754 5 1 1 43753
0 43755 7 1 2 71618 43754
0 43756 7 1 2 43752 43755
0 43757 7 1 2 43746 43756
0 43758 5 2 1 43757
0 43759 7 1 2 78910 79503
0 43760 5 1 1 43759
0 43761 7 1 2 60841 78205
0 43762 5 1 1 43761
0 43763 7 1 2 58947 77117
0 43764 5 1 1 43763
0 43765 7 1 2 43762 43764
0 43766 5 1 1 43765
0 43767 7 1 2 48011 43766
0 43768 5 1 1 43767
0 43769 7 2 2 57686 61474
0 43770 5 1 1 79505
0 43771 7 1 2 66644 43770
0 43772 5 1 1 43771
0 43773 7 1 2 48012 65321
0 43774 5 1 1 43773
0 43775 7 1 2 56967 65211
0 43776 5 1 1 43775
0 43777 7 1 2 48444 62331
0 43778 7 1 2 68017 43777
0 43779 5 1 1 43778
0 43780 7 1 2 43776 43779
0 43781 7 1 2 43774 43780
0 43782 5 1 1 43781
0 43783 7 1 2 58316 43782
0 43784 5 1 1 43783
0 43785 7 1 2 43772 43784
0 43786 7 1 2 43768 43785
0 43787 5 1 1 43786
0 43788 7 1 2 74296 43787
0 43789 5 1 1 43788
0 43790 7 1 2 59091 76886
0 43791 7 1 2 75570 43790
0 43792 5 1 1 43791
0 43793 7 1 2 76272 43792
0 43794 5 1 1 43793
0 43795 7 1 2 43789 43794
0 43796 5 1 1 43795
0 43797 7 1 2 56595 43796
0 43798 5 1 1 43797
0 43799 7 2 2 67980 76322
0 43800 5 1 1 79507
0 43801 7 1 2 77729 79508
0 43802 5 1 1 43801
0 43803 7 2 2 57966 74297
0 43804 7 1 2 77178 79509
0 43805 5 1 1 43804
0 43806 7 1 2 43802 43805
0 43807 5 1 1 43806
0 43808 7 1 2 55830 43807
0 43809 5 1 1 43808
0 43810 7 1 2 59302 63923
0 43811 7 1 2 65787 43810
0 43812 5 1 1 43811
0 43813 7 1 2 48269 43812
0 43814 5 1 1 43813
0 43815 7 1 2 65212 59584
0 43816 5 1 1 43815
0 43817 7 1 2 59198 43816
0 43818 7 1 2 43814 43817
0 43819 5 1 1 43818
0 43820 7 1 2 74298 43819
0 43821 5 1 1 43820
0 43822 7 2 2 65788 70649
0 43823 5 1 1 79511
0 43824 7 1 2 56968 76323
0 43825 7 1 2 43823 43824
0 43826 5 1 1 43825
0 43827 7 1 2 43821 43826
0 43828 5 1 1 43827
0 43829 7 1 2 67981 43828
0 43830 5 1 1 43829
0 43831 7 1 2 43809 43830
0 43832 7 1 2 43798 43831
0 43833 5 1 1 43832
0 43834 7 1 2 48831 43833
0 43835 5 1 1 43834
0 43836 7 1 2 76887 79512
0 43837 5 1 1 43836
0 43838 7 1 2 49505 43837
0 43839 5 1 1 43838
0 43840 7 1 2 63105 43839
0 43841 5 1 1 43840
0 43842 7 1 2 48563 43841
0 43843 5 1 1 43842
0 43844 7 1 2 59273 75731
0 43845 5 1 1 43844
0 43846 7 1 2 43843 43845
0 43847 5 1 1 43846
0 43848 7 1 2 57967 76273
0 43849 7 1 2 43847 43848
0 43850 5 1 1 43849
0 43851 7 1 2 55145 78474
0 43852 5 1 1 43851
0 43853 7 1 2 43800 43852
0 43854 5 1 1 43853
0 43855 7 1 2 48832 43854
0 43856 5 1 1 43855
0 43857 7 1 2 67290 73081
0 43858 5 1 1 43857
0 43859 7 1 2 43856 43858
0 43860 5 1 1 43859
0 43861 7 1 2 48013 43860
0 43862 5 1 1 43861
0 43863 7 1 2 63213 66126
0 43864 5 1 1 43863
0 43865 7 1 2 43862 43864
0 43866 5 1 1 43865
0 43867 7 1 2 48445 43866
0 43868 5 1 1 43867
0 43869 7 2 2 57297 76265
0 43870 7 1 2 62332 79513
0 43871 5 1 1 43870
0 43872 7 1 2 43868 43871
0 43873 5 1 1 43872
0 43874 7 1 2 67469 43873
0 43875 5 1 1 43874
0 43876 7 1 2 60317 79514
0 43877 5 1 1 43876
0 43878 7 2 2 63648 77090
0 43879 7 1 2 48270 79515
0 43880 7 1 2 67995 43879
0 43881 5 1 1 43880
0 43882 7 1 2 43877 43881
0 43883 5 1 1 43882
0 43884 7 1 2 58948 43883
0 43885 5 1 1 43884
0 43886 7 1 2 74299 78892
0 43887 5 1 1 43886
0 43888 7 1 2 67281 79516
0 43889 5 1 1 43888
0 43890 7 1 2 43887 43889
0 43891 5 1 1 43890
0 43892 7 1 2 56596 43891
0 43893 5 1 1 43892
0 43894 7 1 2 77154 79510
0 43895 5 1 1 43894
0 43896 7 1 2 43893 43895
0 43897 5 1 1 43896
0 43898 7 1 2 48833 43897
0 43899 5 1 1 43898
0 43900 7 1 2 43885 43899
0 43901 5 1 1 43900
0 43902 7 1 2 58632 43901
0 43903 5 1 1 43902
0 43904 7 1 2 43875 43903
0 43905 7 1 2 43850 43904
0 43906 7 1 2 43835 43905
0 43907 5 1 1 43906
0 43908 7 1 2 53746 43907
0 43909 5 1 1 43908
0 43910 7 1 2 69639 75901
0 43911 5 1 1 43910
0 43912 7 1 2 70175 77180
0 43913 5 1 1 43912
0 43914 7 1 2 55146 43913
0 43915 5 1 1 43914
0 43916 7 1 2 52726 43915
0 43917 5 1 1 43916
0 43918 7 1 2 53589 43917
0 43919 5 1 1 43918
0 43920 7 1 2 65819 74300
0 43921 5 1 1 43920
0 43922 7 1 2 57545 65273
0 43923 7 1 2 76324 43922
0 43924 5 1 1 43923
0 43925 7 1 2 43921 43924
0 43926 5 1 1 43925
0 43927 7 1 2 48271 43926
0 43928 5 1 1 43927
0 43929 7 1 2 62738 74301
0 43930 5 1 1 43929
0 43931 7 1 2 60226 78945
0 43932 5 1 1 43931
0 43933 7 1 2 43930 43932
0 43934 5 1 1 43933
0 43935 7 1 2 62418 43934
0 43936 5 1 1 43935
0 43937 7 1 2 48014 70237
0 43938 5 1 1 43937
0 43939 7 1 2 59303 43938
0 43940 5 1 1 43939
0 43941 7 1 2 74302 43940
0 43942 5 1 1 43941
0 43943 7 1 2 43936 43942
0 43944 7 1 2 43928 43943
0 43945 5 1 1 43944
0 43946 7 1 2 55831 43945
0 43947 5 1 1 43946
0 43948 7 1 2 58733 71632
0 43949 5 1 1 43948
0 43950 7 1 2 49815 43949
0 43951 5 1 1 43950
0 43952 7 1 2 60977 57808
0 43953 5 1 1 43952
0 43954 7 1 2 23285 43953
0 43955 5 1 1 43954
0 43956 7 1 2 56779 43955
0 43957 5 1 1 43956
0 43958 7 1 2 48015 76177
0 43959 5 1 1 43958
0 43960 7 1 2 60352 78116
0 43961 5 1 1 43960
0 43962 7 1 2 57715 43961
0 43963 7 1 2 43959 43962
0 43964 7 1 2 43957 43963
0 43965 5 1 1 43964
0 43966 7 1 2 73082 43965
0 43967 5 1 1 43966
0 43968 7 1 2 43951 43967
0 43969 7 1 2 43947 43968
0 43970 7 1 2 43919 43969
0 43971 5 1 1 43970
0 43972 7 1 2 73321 43971
0 43973 5 1 1 43972
0 43974 7 1 2 43911 43973
0 43975 7 1 2 43909 43974
0 43976 5 2 1 43975
0 43977 7 1 2 51792 79517
0 43978 5 1 1 43977
0 43979 7 1 2 43760 43978
0 43980 5 1 1 43979
0 43981 7 1 2 51442 43980
0 43982 5 1 1 43981
0 43983 7 1 2 48446 65364
0 43984 5 1 1 43983
0 43985 7 1 2 60428 5332
0 43986 7 2 2 43984 43985
0 43987 7 1 2 78911 79519
0 43988 5 1 1 43987
0 43989 7 1 2 73777 69030
0 43990 5 1 1 43989
0 43991 7 1 2 71513 69733
0 43992 5 1 1 43991
0 43993 7 1 2 43990 43992
0 43994 5 1 1 43993
0 43995 7 1 2 53590 43994
0 43996 5 1 1 43995
0 43997 7 1 2 71514 69034
0 43998 5 1 1 43997
0 43999 7 1 2 43996 43998
0 44000 5 1 1 43999
0 44001 7 1 2 60227 44000
0 44002 5 1 1 44001
0 44003 7 1 2 43988 44002
0 44004 5 1 1 44003
0 44005 7 1 2 51443 44004
0 44006 5 1 1 44005
0 44007 7 2 2 55417 78870
0 44008 7 1 2 50556 51793
0 44009 7 1 2 77197 44008
0 44010 7 1 2 79521 44009
0 44011 5 1 1 44010
0 44012 7 1 2 44006 44011
0 44013 5 1 1 44012
0 44014 7 1 2 70779 44013
0 44015 5 1 1 44014
0 44016 7 1 2 57546 61491
0 44017 5 1 1 44016
0 44018 7 1 2 64575 44017
0 44019 5 1 1 44018
0 44020 7 1 2 56258 62793
0 44021 5 4 1 44020
0 44022 7 1 2 77341 79523
0 44023 5 1 1 44022
0 44024 7 1 2 57803 44023
0 44025 5 1 1 44024
0 44026 7 1 2 48675 44025
0 44027 5 1 1 44026
0 44028 7 1 2 67233 74755
0 44029 5 1 1 44028
0 44030 7 1 2 57347 44029
0 44031 5 1 1 44030
0 44032 7 1 2 48016 44031
0 44033 5 1 1 44032
0 44034 7 1 2 48676 76726
0 44035 5 1 1 44034
0 44036 7 1 2 44033 44035
0 44037 5 1 1 44036
0 44038 7 1 2 62309 44037
0 44039 5 1 1 44038
0 44040 7 1 2 58492 66237
0 44041 7 1 2 77342 44040
0 44042 5 1 1 44041
0 44043 7 1 2 44039 44042
0 44044 7 1 2 44027 44043
0 44045 5 1 1 44044
0 44046 7 1 2 49639 44045
0 44047 5 1 1 44046
0 44048 7 1 2 76563 30264
0 44049 5 1 1 44048
0 44050 7 1 2 49640 77700
0 44051 7 1 2 44049 44050
0 44052 5 1 1 44051
0 44053 7 2 2 61316 58912
0 44054 7 1 2 57547 78373
0 44055 5 1 1 44054
0 44056 7 1 2 79527 44055
0 44057 5 1 1 44056
0 44058 7 1 2 76570 44057
0 44059 5 1 1 44058
0 44060 7 1 2 3819 44059
0 44061 7 1 2 44052 44060
0 44062 5 1 1 44061
0 44063 7 1 2 61588 44062
0 44064 5 1 1 44063
0 44065 7 1 2 74756 78374
0 44066 5 1 1 44065
0 44067 7 1 2 79528 44066
0 44068 5 1 1 44067
0 44069 7 1 2 48017 44068
0 44070 5 1 1 44069
0 44071 7 1 2 62587 76727
0 44072 5 1 1 44071
0 44073 7 1 2 44070 44072
0 44074 5 1 1 44073
0 44075 7 1 2 62310 44074
0 44076 5 1 1 44075
0 44077 7 1 2 62588 57799
0 44078 5 1 1 44077
0 44079 7 1 2 62589 79524
0 44080 5 1 1 44079
0 44081 7 1 2 48564 64261
0 44082 7 1 2 62204 44081
0 44083 5 1 1 44082
0 44084 7 1 2 44080 44083
0 44085 5 1 1 44084
0 44086 7 1 2 77343 44085
0 44087 5 1 1 44086
0 44088 7 1 2 44078 44087
0 44089 7 1 2 44076 44088
0 44090 7 1 2 44064 44089
0 44091 7 1 2 44047 44090
0 44092 5 1 1 44091
0 44093 7 1 2 50557 44092
0 44094 5 1 1 44093
0 44095 7 1 2 44019 44094
0 44096 5 1 1 44095
0 44097 7 1 2 71870 44096
0 44098 5 1 1 44097
0 44099 7 2 2 54413 61492
0 44100 5 1 1 79529
0 44101 7 1 2 57548 79530
0 44102 5 1 1 44101
0 44103 7 1 2 78985 44102
0 44104 5 1 1 44103
0 44105 7 2 2 44098 44104
0 44106 5 1 1 79531
0 44107 7 1 2 56665 62019
0 44108 5 1 1 44107
0 44109 7 1 2 70697 44108
0 44110 5 1 1 44109
0 44111 7 1 2 59665 44110
0 44112 5 1 1 44111
0 44113 7 1 2 56426 44112
0 44114 5 2 1 44113
0 44115 7 1 2 79167 79533
0 44116 5 1 1 44115
0 44117 7 1 2 79532 44116
0 44118 5 1 1 44117
0 44119 7 1 2 68964 44118
0 44120 5 1 1 44119
0 44121 7 1 2 44015 44120
0 44122 7 1 2 43982 44121
0 44123 5 1 1 44122
0 44124 7 1 2 51653 44123
0 44125 5 1 1 44124
0 44126 7 1 2 55418 79161
0 44127 5 1 1 44126
0 44128 7 1 2 75642 44127
0 44129 5 1 1 44128
0 44130 7 1 2 52347 44129
0 44131 5 1 1 44130
0 44132 7 1 2 79009 44131
0 44133 5 1 1 44132
0 44134 7 1 2 53591 44133
0 44135 5 1 1 44134
0 44136 7 1 2 52348 77325
0 44137 7 1 2 76502 44136
0 44138 5 1 1 44137
0 44139 7 1 2 79014 44138
0 44140 7 1 2 44135 44139
0 44141 5 1 1 44140
0 44142 7 1 2 53747 44141
0 44143 5 1 1 44142
0 44144 7 1 2 78048 44143
0 44145 5 1 1 44144
0 44146 7 1 2 55579 44145
0 44147 5 1 1 44146
0 44148 7 1 2 70377 71461
0 44149 7 1 2 78796 44148
0 44150 5 1 1 44149
0 44151 7 1 2 44147 44150
0 44152 5 1 1 44151
0 44153 7 1 2 60020 44152
0 44154 5 1 1 44153
0 44155 7 1 2 9423 28618
0 44156 5 3 1 44155
0 44157 7 1 2 51170 71462
0 44158 7 1 2 79535 44157
0 44159 5 1 1 44158
0 44160 7 1 2 72725 44159
0 44161 5 1 1 44160
0 44162 7 1 2 67904 44161
0 44163 5 1 1 44162
0 44164 7 1 2 12785 32880
0 44165 5 1 1 44164
0 44166 7 1 2 49816 44165
0 44167 5 1 1 44166
0 44168 7 1 2 51654 44167
0 44169 7 1 2 44163 44168
0 44170 5 1 1 44169
0 44171 7 1 2 70378 78005
0 44172 5 1 1 44171
0 44173 7 1 2 79005 44172
0 44174 5 1 1 44173
0 44175 7 1 2 55419 44174
0 44176 5 1 1 44175
0 44177 7 1 2 75643 44176
0 44178 5 1 1 44177
0 44179 7 1 2 53592 44178
0 44180 5 1 1 44179
0 44181 7 1 2 72933 78712
0 44182 5 1 1 44181
0 44183 7 1 2 70379 78709
0 44184 5 1 1 44183
0 44185 7 1 2 44182 44184
0 44186 7 1 2 44180 44185
0 44187 5 1 1 44186
0 44188 7 1 2 53135 44187
0 44189 5 1 1 44188
0 44190 7 1 2 53593 79007
0 44191 5 1 1 44190
0 44192 7 1 2 44189 44191
0 44193 5 1 1 44192
0 44194 7 1 2 59950 44193
0 44195 5 1 1 44194
0 44196 7 1 2 51444 70380
0 44197 7 1 2 78477 44196
0 44198 5 1 1 44197
0 44199 7 1 2 44195 44198
0 44200 5 1 1 44199
0 44201 7 1 2 53748 44200
0 44202 5 1 1 44201
0 44203 7 1 2 70381 75902
0 44204 5 1 1 44203
0 44205 7 1 2 56666 60610
0 44206 7 1 2 78953 44205
0 44207 5 1 1 44206
0 44208 7 1 2 44204 44207
0 44209 5 1 1 44208
0 44210 7 1 2 67890 44209
0 44211 5 1 1 44210
0 44212 7 1 2 55580 44211
0 44213 7 1 2 44202 44212
0 44214 5 1 1 44213
0 44215 7 1 2 44170 44214
0 44216 5 1 1 44215
0 44217 7 1 2 44154 44216
0 44218 5 1 1 44217
0 44219 7 1 2 52830 44218
0 44220 5 1 1 44219
0 44221 7 1 2 79431 79026
0 44222 5 1 1 44221
0 44223 7 1 2 64822 68755
0 44224 5 1 1 44223
0 44225 7 1 2 53399 55959
0 44226 7 1 2 73472 44225
0 44227 5 1 1 44226
0 44228 7 1 2 44224 44227
0 44229 5 1 1 44228
0 44230 7 1 2 52582 44229
0 44231 5 1 1 44230
0 44232 7 1 2 73828 77949
0 44233 5 1 1 44232
0 44234 7 1 2 44231 44233
0 44235 5 1 1 44234
0 44236 7 1 2 72413 44235
0 44237 5 1 1 44236
0 44238 7 1 2 71323 68731
0 44239 5 1 1 44238
0 44240 7 1 2 49980 74822
0 44241 5 1 1 44240
0 44242 7 1 2 44239 44241
0 44243 5 1 1 44242
0 44244 7 1 2 71535 44243
0 44245 5 1 1 44244
0 44246 7 2 2 66106 73291
0 44247 5 1 1 79538
0 44248 7 1 2 66001 44247
0 44249 5 1 1 44248
0 44250 7 1 2 78886 44249
0 44251 5 1 1 44250
0 44252 7 1 2 65996 70562
0 44253 5 1 1 44252
0 44254 7 1 2 44251 44253
0 44255 7 1 2 44245 44254
0 44256 7 1 2 44237 44255
0 44257 5 1 1 44256
0 44258 7 1 2 51171 44257
0 44259 5 1 1 44258
0 44260 7 1 2 44222 44259
0 44261 5 1 1 44260
0 44262 7 1 2 74838 44261
0 44263 5 1 1 44262
0 44264 7 1 2 57687 75182
0 44265 7 1 2 79381 44264
0 44266 7 1 2 78668 44265
0 44267 5 1 1 44266
0 44268 7 1 2 44263 44267
0 44269 5 1 1 44268
0 44270 7 1 2 50307 44269
0 44271 5 1 1 44270
0 44272 7 1 2 67645 75065
0 44273 5 1 1 44272
0 44274 7 1 2 32681 44273
0 44275 5 1 1 44274
0 44276 7 1 2 52349 44275
0 44277 5 1 1 44276
0 44278 7 1 2 71584 73646
0 44279 5 1 1 44278
0 44280 7 1 2 44277 44279
0 44281 5 1 1 44280
0 44282 7 1 2 55420 44281
0 44283 5 1 1 44282
0 44284 7 1 2 49641 67473
0 44285 5 1 1 44284
0 44286 7 1 2 71316 44285
0 44287 5 1 1 44286
0 44288 7 1 2 78430 44287
0 44289 5 1 1 44288
0 44290 7 1 2 44283 44289
0 44291 5 1 1 44290
0 44292 7 1 2 52831 44291
0 44293 5 1 1 44292
0 44294 7 1 2 59923 79386
0 44295 5 1 1 44294
0 44296 7 1 2 66769 71771
0 44297 7 1 2 73497 44296
0 44298 5 1 1 44297
0 44299 7 1 2 44295 44298
0 44300 5 1 1 44299
0 44301 7 1 2 55421 44300
0 44302 5 1 1 44301
0 44303 7 1 2 68597 78741
0 44304 5 2 1 44303
0 44305 7 1 2 44302 79540
0 44306 5 1 1 44305
0 44307 7 1 2 58783 44306
0 44308 5 1 1 44307
0 44309 7 1 2 69288 72138
0 44310 7 1 2 70608 44309
0 44311 5 1 1 44310
0 44312 7 1 2 59924 65997
0 44313 7 1 2 71318 44312
0 44314 5 1 1 44313
0 44315 7 1 2 44311 44314
0 44316 5 1 1 44315
0 44317 7 1 2 53594 44316
0 44318 5 1 1 44317
0 44319 7 1 2 44308 44318
0 44320 7 1 2 44293 44319
0 44321 7 1 2 44271 44320
0 44322 5 1 1 44321
0 44323 7 1 2 60880 44322
0 44324 5 1 1 44323
0 44325 7 1 2 66107 79084
0 44326 5 1 1 44325
0 44327 7 1 2 56477 69245
0 44328 5 1 1 44327
0 44329 7 1 2 68505 44328
0 44330 5 1 1 44329
0 44331 7 2 2 69579 44330
0 44332 7 3 2 65998 79542
0 44333 5 1 1 79544
0 44334 7 2 2 51172 70382
0 44335 7 1 2 79545 79547
0 44336 5 1 1 44335
0 44337 7 1 2 44326 44336
0 44338 5 1 1 44337
0 44339 7 1 2 60021 44338
0 44340 5 1 1 44339
0 44341 7 1 2 56667 65741
0 44342 7 1 2 60611 44341
0 44343 5 1 1 44342
0 44344 7 1 2 67802 44343
0 44345 5 1 1 44344
0 44346 7 1 2 78900 44345
0 44347 5 1 1 44346
0 44348 7 1 2 79135 44347
0 44349 5 1 1 44348
0 44350 7 1 2 51445 44349
0 44351 5 1 1 44350
0 44352 7 1 2 79546 79536
0 44353 5 1 1 44352
0 44354 7 1 2 44351 44353
0 44355 5 1 1 44354
0 44356 7 1 2 51173 44355
0 44357 5 1 1 44356
0 44358 7 5 2 52727 67813
0 44359 5 1 1 79549
0 44360 7 1 2 79433 79550
0 44361 5 1 1 44360
0 44362 7 1 2 51655 78602
0 44363 5 1 1 44362
0 44364 7 1 2 44361 44363
0 44365 5 1 1 44364
0 44366 7 1 2 56478 44365
0 44367 5 1 1 44366
0 44368 7 1 2 51656 73843
0 44369 5 1 1 44368
0 44370 7 1 2 44367 44369
0 44371 5 1 1 44370
0 44372 7 1 2 67127 44371
0 44373 5 1 1 44372
0 44374 7 1 2 44357 44373
0 44375 7 1 2 44340 44374
0 44376 7 1 2 44324 44375
0 44377 7 1 2 44220 44376
0 44378 5 2 1 44377
0 44379 7 1 2 51794 79554
0 44380 5 1 1 44379
0 44381 7 1 2 53400 67792
0 44382 5 1 1 44381
0 44383 7 1 2 53595 67092
0 44384 5 1 1 44383
0 44385 7 1 2 44382 44384
0 44386 5 1 1 44385
0 44387 7 1 2 52583 44386
0 44388 5 1 1 44387
0 44389 7 1 2 51657 73542
0 44390 5 1 1 44389
0 44391 7 1 2 44388 44390
0 44392 5 1 1 44391
0 44393 7 1 2 55422 44392
0 44394 5 1 1 44393
0 44395 7 1 2 65742 76002
0 44396 5 1 1 44395
0 44397 7 1 2 44394 44396
0 44398 5 1 1 44397
0 44399 7 1 2 52832 44398
0 44400 5 1 1 44399
0 44401 7 1 2 44333 44400
0 44402 5 1 1 44401
0 44403 7 1 2 56780 65898
0 44404 5 2 1 44403
0 44405 7 1 2 44402 79556
0 44406 5 1 1 44405
0 44407 7 1 2 55960 61831
0 44408 5 1 1 44407
0 44409 7 1 2 57688 70802
0 44410 5 1 1 44409
0 44411 7 1 2 44408 44410
0 44412 5 1 1 44411
0 44413 7 1 2 7787 73716
0 44414 5 1 1 44413
0 44415 7 1 2 70582 44414
0 44416 5 1 1 44415
0 44417 7 1 2 66108 44416
0 44418 7 1 2 44412 44417
0 44419 5 1 1 44418
0 44420 7 1 2 44406 44419
0 44421 5 1 1 44420
0 44422 7 1 2 51174 44421
0 44423 5 1 1 44422
0 44424 7 1 2 71772 43600
0 44425 7 1 2 73717 44424
0 44426 5 1 1 44425
0 44427 7 1 2 49817 73544
0 44428 7 1 2 73698 44427
0 44429 7 1 2 70803 44428
0 44430 5 1 1 44429
0 44431 7 1 2 44426 44430
0 44432 5 1 1 44431
0 44433 7 1 2 51446 44432
0 44434 5 1 1 44433
0 44435 7 2 2 63144 77265
0 44436 5 1 1 79558
0 44437 7 1 2 70798 79559
0 44438 5 2 1 44437
0 44439 7 1 2 76503 78752
0 44440 7 1 2 79560 44439
0 44441 5 1 1 44440
0 44442 7 1 2 44434 44441
0 44443 7 2 2 44423 44442
0 44444 5 1 1 79562
0 44445 7 3 2 67111 69537
0 44446 5 1 1 79564
0 44447 7 1 2 44436 79565
0 44448 5 1 1 44447
0 44449 7 1 2 70799 44448
0 44450 5 1 1 44449
0 44451 7 1 2 48976 73790
0 44452 5 1 1 44451
0 44453 7 1 2 44446 44452
0 44454 5 1 1 44453
0 44455 7 1 2 53596 44454
0 44456 7 1 2 44450 44455
0 44457 5 1 1 44456
0 44458 7 1 2 79541 44457
0 44459 5 1 1 44458
0 44460 7 1 2 58784 44459
0 44461 5 1 1 44460
0 44462 7 1 2 79563 44461
0 44463 5 1 1 44462
0 44464 7 1 2 51795 44463
0 44465 5 1 1 44464
0 44466 7 1 2 73545 68529
0 44467 7 1 2 79096 44466
0 44468 7 1 2 70804 44467
0 44469 5 1 1 44468
0 44470 7 1 2 44465 44469
0 44471 5 1 1 44470
0 44472 7 1 2 50558 44471
0 44473 5 1 1 44472
0 44474 7 3 2 75183 70609
0 44475 7 2 2 72297 79567
0 44476 5 1 1 79570
0 44477 7 1 2 44473 44476
0 44478 7 1 2 44380 44477
0 44479 5 1 1 44478
0 44480 7 1 2 57068 44479
0 44481 5 1 1 44480
0 44482 7 1 2 75910 41171
0 44483 5 1 1 44482
0 44484 7 1 2 67891 44483
0 44485 5 1 1 44484
0 44486 7 1 2 72698 79216
0 44487 5 1 1 44486
0 44488 7 1 2 75110 44487
0 44489 5 1 1 44488
0 44490 7 1 2 56597 77806
0 44491 5 1 1 44490
0 44492 7 1 2 58493 74645
0 44493 5 1 1 44492
0 44494 7 1 2 44491 44493
0 44495 5 1 1 44494
0 44496 7 1 2 48272 44495
0 44497 5 1 1 44496
0 44498 7 1 2 57377 68041
0 44499 5 1 1 44498
0 44500 7 1 2 44497 44499
0 44501 5 1 1 44500
0 44502 7 1 2 58883 44501
0 44503 5 1 1 44502
0 44504 7 1 2 57378 60081
0 44505 5 1 1 44504
0 44506 7 1 2 57114 59330
0 44507 5 1 1 44506
0 44508 7 1 2 57367 44507
0 44509 5 1 1 44508
0 44510 7 1 2 60938 44509
0 44511 5 1 1 44510
0 44512 7 1 2 56787 44511
0 44513 5 1 1 44512
0 44514 7 1 2 60708 44513
0 44515 5 1 1 44514
0 44516 7 1 2 44505 44515
0 44517 7 1 2 44503 44516
0 44518 5 1 1 44517
0 44519 7 1 2 51447 44518
0 44520 5 1 1 44519
0 44521 7 1 2 44489 44520
0 44522 5 1 1 44521
0 44523 7 1 2 48447 44522
0 44524 5 1 1 44523
0 44525 7 1 2 75111 77111
0 44526 5 1 1 44525
0 44527 7 1 2 57726 61709
0 44528 5 1 1 44527
0 44529 7 1 2 67499 68156
0 44530 5 1 1 44529
0 44531 7 1 2 44528 44530
0 44532 5 1 1 44531
0 44533 7 1 2 69891 44532
0 44534 5 1 1 44533
0 44535 7 1 2 61997 64101
0 44536 5 1 1 44535
0 44537 7 1 2 57727 44536
0 44538 5 1 1 44537
0 44539 7 1 2 44534 44538
0 44540 5 1 1 44539
0 44541 7 1 2 51448 44540
0 44542 5 1 1 44541
0 44543 7 1 2 44526 44542
0 44544 5 1 1 44543
0 44545 7 1 2 54414 44544
0 44546 5 1 1 44545
0 44547 7 1 2 75112 77366
0 44548 5 1 1 44547
0 44549 7 2 2 51449 57379
0 44550 7 1 2 77172 79572
0 44551 5 1 1 44550
0 44552 7 1 2 44548 44551
0 44553 5 1 1 44552
0 44554 7 1 2 49257 44553
0 44555 5 1 1 44554
0 44556 7 1 2 75113 78842
0 44557 5 1 1 44556
0 44558 7 1 2 44555 44557
0 44559 5 1 1 44558
0 44560 7 1 2 48273 44559
0 44561 5 1 1 44560
0 44562 7 1 2 53256 74024
0 44563 5 1 1 44562
0 44564 7 1 2 75114 44563
0 44565 5 1 1 44564
0 44566 7 1 2 75115 72784
0 44567 5 1 1 44566
0 44568 7 1 2 30493 79573
0 44569 5 1 1 44568
0 44570 7 1 2 44567 44569
0 44571 5 1 1 44570
0 44572 7 1 2 49382 44571
0 44573 5 1 1 44572
0 44574 7 1 2 19934 75116
0 44575 5 1 1 44574
0 44576 7 1 2 48677 44575
0 44577 5 1 1 44576
0 44578 7 1 2 53597 76295
0 44579 7 1 2 44577 44578
0 44580 7 1 2 75117 75796
0 44581 5 1 1 44580
0 44582 7 1 2 48565 44581
0 44583 5 1 1 44582
0 44584 7 1 2 56259 78669
0 44585 5 1 1 44584
0 44586 7 1 2 44583 44585
0 44587 7 1 2 44579 44586
0 44588 7 1 2 44573 44587
0 44589 7 1 2 44565 44588
0 44590 7 1 2 44561 44589
0 44591 7 1 2 44546 44590
0 44592 7 1 2 44524 44591
0 44593 5 1 1 44592
0 44594 7 1 2 72700 25269
0 44595 7 1 2 79115 44594
0 44596 5 1 1 44595
0 44597 7 1 2 53749 44596
0 44598 7 1 2 44593 44597
0 44599 5 1 1 44598
0 44600 7 1 2 44485 44599
0 44601 5 1 1 44600
0 44602 7 1 2 52833 44601
0 44603 5 1 1 44602
0 44604 7 1 2 53750 78515
0 44605 5 1 1 44604
0 44606 7 1 2 78834 44605
0 44607 5 1 1 44606
0 44608 7 1 2 56260 44607
0 44609 5 1 1 44608
0 44610 7 1 2 68756 78670
0 44611 5 1 1 44610
0 44612 7 1 2 44609 44611
0 44613 5 2 1 44612
0 44614 7 1 2 55961 79574
0 44615 5 1 1 44614
0 44616 7 1 2 79125 44615
0 44617 5 1 1 44616
0 44618 7 1 2 52834 44617
0 44619 5 1 1 44618
0 44620 7 1 2 15218 68607
0 44621 5 1 1 44620
0 44622 7 1 2 52728 44621
0 44623 5 1 1 44622
0 44624 7 1 2 75091 44623
0 44625 5 1 1 44624
0 44626 7 1 2 56479 44625
0 44627 5 1 1 44626
0 44628 7 1 2 48977 79551
0 44629 5 1 1 44628
0 44630 7 1 2 44627 44629
0 44631 5 2 1 44630
0 44632 7 1 2 79122 79576
0 44633 5 1 1 44632
0 44634 7 1 2 44619 44633
0 44635 5 1 1 44634
0 44636 7 1 2 70283 44635
0 44637 5 1 1 44636
0 44638 7 1 2 66054 78901
0 44639 5 1 1 44638
0 44640 7 1 2 78939 44639
0 44641 5 1 1 44640
0 44642 7 1 2 69289 44641
0 44643 5 1 1 44642
0 44644 7 1 2 44637 44643
0 44645 7 1 2 44603 44644
0 44646 5 1 1 44645
0 44647 7 1 2 51175 44646
0 44648 5 1 1 44647
0 44649 7 1 2 79088 40772
0 44650 5 1 1 44649
0 44651 7 1 2 56427 70506
0 44652 5 1 1 44651
0 44653 7 1 2 58573 44652
0 44654 5 1 1 44653
0 44655 7 1 2 70280 44654
0 44656 5 1 1 44655
0 44657 7 1 2 44650 44656
0 44658 5 1 1 44657
0 44659 7 1 2 58412 61207
0 44660 5 1 1 44659
0 44661 7 1 2 56428 61067
0 44662 5 1 1 44661
0 44663 7 1 2 44660 44662
0 44664 5 1 1 44663
0 44665 7 1 2 61844 44664
0 44666 5 1 1 44665
0 44667 7 1 2 67205 7113
0 44668 5 1 1 44667
0 44669 7 1 2 48018 44668
0 44670 5 1 1 44669
0 44671 7 1 2 56429 62818
0 44672 5 1 1 44671
0 44673 7 1 2 48448 79525
0 44674 5 1 1 44673
0 44675 7 1 2 70627 78076
0 44676 7 1 2 44674 44675
0 44677 5 1 1 44676
0 44678 7 1 2 58261 44677
0 44679 5 1 1 44678
0 44680 7 1 2 44672 44679
0 44681 7 1 2 44670 44680
0 44682 5 1 1 44681
0 44683 7 1 2 55832 44682
0 44684 5 1 1 44683
0 44685 7 1 2 61208 67301
0 44686 5 1 1 44685
0 44687 7 1 2 48566 66564
0 44688 5 1 1 44687
0 44689 7 1 2 53401 44688
0 44690 7 1 2 44686 44689
0 44691 7 1 2 61991 78819
0 44692 5 1 1 44691
0 44693 7 1 2 52584 62030
0 44694 5 1 1 44693
0 44695 7 1 2 30000 44694
0 44696 5 1 1 44695
0 44697 7 1 2 44692 44696
0 44698 7 1 2 44690 44697
0 44699 7 1 2 44684 44698
0 44700 7 1 2 44666 44699
0 44701 5 1 1 44700
0 44702 7 1 2 55962 77275
0 44703 5 1 1 44702
0 44704 7 1 2 49642 77214
0 44705 7 1 2 44703 44704
0 44706 7 1 2 74876 44705
0 44707 5 1 1 44706
0 44708 7 1 2 55147 44707
0 44709 7 1 2 44701 44708
0 44710 5 1 1 44709
0 44711 7 1 2 22878 44710
0 44712 5 1 1 44711
0 44713 7 1 2 79375 44712
0 44714 5 1 1 44713
0 44715 7 1 2 44658 44714
0 44716 5 1 1 44715
0 44717 7 1 2 51450 44716
0 44718 5 1 1 44717
0 44719 7 3 2 51451 44100
0 44720 7 1 2 79076 79578
0 44721 5 1 1 44720
0 44722 7 1 2 48978 60499
0 44723 7 1 2 73548 44722
0 44724 5 1 1 44723
0 44725 7 1 2 78699 44724
0 44726 5 1 1 44725
0 44727 7 1 2 52026 44726
0 44728 5 1 1 44727
0 44729 7 1 2 68598 70508
0 44730 5 1 1 44729
0 44731 7 1 2 44728 44730
0 44732 5 1 1 44731
0 44733 7 1 2 71515 44732
0 44734 5 1 1 44733
0 44735 7 1 2 44721 44734
0 44736 5 1 1 44735
0 44737 7 1 2 70818 44736
0 44738 5 1 1 44737
0 44739 7 2 2 51452 61832
0 44740 5 1 1 79581
0 44741 7 2 2 56480 67963
0 44742 5 1 1 79583
0 44743 7 1 2 63665 79584
0 44744 7 1 2 79582 44743
0 44745 5 1 1 44744
0 44746 7 1 2 44738 44745
0 44747 5 1 1 44746
0 44748 7 1 2 53751 44747
0 44749 5 1 1 44748
0 44750 7 5 2 58843 71210
0 44751 7 1 2 79120 79585
0 44752 5 1 1 44751
0 44753 7 1 2 7414 44752
0 44754 5 1 1 44753
0 44755 7 1 2 78150 44754
0 44756 5 1 1 44755
0 44757 7 1 2 61258 71116
0 44758 5 1 1 44757
0 44759 7 1 2 67539 44758
0 44760 5 1 1 44759
0 44761 7 1 2 48834 44760
0 44762 5 1 1 44761
0 44763 7 1 2 53752 44762
0 44764 7 1 2 44756 44763
0 44765 5 1 1 44764
0 44766 7 1 2 61250 76431
0 44767 7 1 2 71212 44766
0 44768 5 1 1 44767
0 44769 7 1 2 44740 44768
0 44770 5 2 1 44769
0 44771 7 1 2 71516 79590
0 44772 5 1 1 44771
0 44773 7 1 2 70663 79113
0 44774 5 1 1 44773
0 44775 7 1 2 49981 44774
0 44776 7 1 2 44772 44775
0 44777 5 1 1 44776
0 44778 7 1 2 50559 44777
0 44779 7 1 2 44765 44778
0 44780 5 1 1 44779
0 44781 7 1 2 61490 78038
0 44782 5 1 1 44781
0 44783 7 1 2 73311 44782
0 44784 5 1 1 44783
0 44785 7 1 2 56261 58785
0 44786 7 1 2 44784 44785
0 44787 5 1 1 44786
0 44788 7 1 2 44780 44787
0 44789 5 1 1 44788
0 44790 7 1 2 53598 44789
0 44791 5 1 1 44790
0 44792 7 1 2 58795 79591
0 44793 5 1 1 44792
0 44794 7 1 2 70664 79579
0 44795 5 1 1 44794
0 44796 7 1 2 44793 44795
0 44797 5 1 1 44796
0 44798 7 1 2 49818 44797
0 44799 5 1 1 44798
0 44800 7 1 2 73207 79186
0 44801 5 1 1 44800
0 44802 7 1 2 44799 44801
0 44803 5 1 1 44802
0 44804 7 1 2 53753 44803
0 44805 5 1 1 44804
0 44806 7 1 2 70819 71313
0 44807 7 1 2 79580 44806
0 44808 5 1 1 44807
0 44809 7 1 2 44805 44808
0 44810 7 1 2 44791 44809
0 44811 5 1 1 44810
0 44812 7 1 2 52835 44811
0 44813 5 1 1 44812
0 44814 7 1 2 44749 44813
0 44815 5 1 1 44814
0 44816 7 1 2 57689 44815
0 44817 5 1 1 44816
0 44818 7 1 2 56262 70509
0 44819 5 1 1 44818
0 44820 7 1 2 70846 44819
0 44821 5 1 1 44820
0 44822 7 1 2 69538 79027
0 44823 7 1 2 44821 44822
0 44824 5 1 1 44823
0 44825 7 1 2 44817 44824
0 44826 7 1 2 44718 44825
0 44827 7 1 2 44648 44826
0 44828 5 1 1 44827
0 44829 7 2 2 67954 44828
0 44830 5 1 1 79592
0 44831 7 1 2 66895 78960
0 44832 5 1 1 44831
0 44833 7 1 2 58786 44832
0 44834 5 1 1 44833
0 44835 7 1 2 66614 78978
0 44836 5 1 1 44835
0 44837 7 1 2 49819 44836
0 44838 7 1 2 44834 44837
0 44839 5 1 1 44838
0 44840 7 1 2 57348 77489
0 44841 5 1 1 44840
0 44842 7 1 2 50560 78006
0 44843 5 1 1 44842
0 44844 7 1 2 44841 44843
0 44845 5 1 1 44844
0 44846 7 1 2 55423 44845
0 44847 5 1 1 44846
0 44848 7 1 2 59905 75246
0 44849 5 1 1 44848
0 44850 7 1 2 44847 44849
0 44851 5 1 1 44850
0 44852 7 1 2 55963 44851
0 44853 5 1 1 44852
0 44854 7 1 2 53599 24948
0 44855 7 1 2 44853 44854
0 44856 5 1 1 44855
0 44857 7 1 2 44839 44856
0 44858 5 1 1 44857
0 44859 7 1 2 53402 73113
0 44860 7 1 2 73478 44859
0 44861 7 1 2 77478 44860
0 44862 5 1 1 44861
0 44863 7 1 2 53754 44862
0 44864 7 1 2 44858 44863
0 44865 5 1 1 44864
0 44866 7 6 2 51453 72715
0 44867 5 1 1 79594
0 44868 7 1 2 73292 71517
0 44869 5 1 1 44868
0 44870 7 1 2 44867 44869
0 44871 5 2 1 44870
0 44872 7 2 2 65478 72978
0 44873 7 1 2 79600 79602
0 44874 5 1 1 44873
0 44875 7 1 2 70610 71375
0 44876 5 1 1 44875
0 44877 7 1 2 49982 44876
0 44878 7 1 2 44874 44877
0 44879 5 1 1 44878
0 44880 7 1 2 55581 44879
0 44881 7 1 2 44865 44880
0 44882 5 1 1 44881
0 44883 7 1 2 59909 78251
0 44884 5 2 1 44883
0 44885 7 2 2 51658 79604
0 44886 7 1 2 64688 79606
0 44887 7 1 2 79127 44886
0 44888 5 1 1 44887
0 44889 7 1 2 44882 44888
0 44890 5 1 1 44889
0 44891 7 1 2 52836 44890
0 44892 5 1 1 44891
0 44893 7 1 2 75103 71319
0 44894 5 1 1 44893
0 44895 7 1 2 55964 66481
0 44896 5 1 1 44895
0 44897 7 1 2 67895 44896
0 44898 5 1 1 44897
0 44899 7 1 2 73778 44898
0 44900 5 1 1 44899
0 44901 7 1 2 44894 44900
0 44902 5 1 1 44901
0 44903 7 1 2 79607 44902
0 44904 5 1 1 44903
0 44905 7 1 2 79577 79603
0 44906 5 1 1 44905
0 44907 7 1 2 63491 79056
0 44908 5 1 1 44907
0 44909 7 1 2 44906 44908
0 44910 5 1 1 44909
0 44911 7 1 2 65743 44910
0 44912 5 1 1 44911
0 44913 7 1 2 44904 44912
0 44914 7 1 2 44892 44913
0 44915 5 1 1 44914
0 44916 7 1 2 50308 44915
0 44917 5 1 1 44916
0 44918 7 1 2 64178 79539
0 44919 5 1 1 44918
0 44920 7 1 2 55582 72728
0 44921 5 1 1 44920
0 44922 7 1 2 37913 44921
0 44923 5 1 1 44922
0 44924 7 1 2 55424 44923
0 44925 5 1 1 44924
0 44926 7 1 2 44919 44925
0 44927 5 1 1 44926
0 44928 7 1 2 55148 44927
0 44929 5 1 1 44928
0 44930 7 1 2 55583 73845
0 44931 5 1 1 44930
0 44932 7 1 2 53755 44931
0 44933 7 1 2 44929 44932
0 44934 5 1 1 44933
0 44935 7 1 2 65999 72716
0 44936 5 1 1 44935
0 44937 7 1 2 71518 71773
0 44938 5 1 1 44937
0 44939 7 1 2 51659 60590
0 44940 5 1 1 44939
0 44941 7 1 2 44938 44940
0 44942 5 1 1 44941
0 44943 7 1 2 73566 44942
0 44944 5 1 1 44943
0 44945 7 1 2 49983 44944
0 44946 7 1 2 44936 44945
0 44947 5 1 1 44946
0 44948 7 1 2 52837 44947
0 44949 7 1 2 44934 44948
0 44950 5 1 1 44949
0 44951 7 2 2 51454 78906
0 44952 7 1 2 66055 79608
0 44953 5 1 1 44952
0 44954 7 1 2 61222 79248
0 44955 5 2 1 44954
0 44956 7 1 2 44953 79610
0 44957 5 1 1 44956
0 44958 7 1 2 51660 44957
0 44959 5 1 1 44958
0 44960 7 1 2 52350 55584
0 44961 7 1 2 71262 44960
0 44962 7 1 2 69290 44961
0 44963 7 1 2 75903 44962
0 44964 5 1 1 44963
0 44965 7 1 2 44959 44964
0 44966 7 1 2 44950 44965
0 44967 7 1 2 44917 44966
0 44968 5 2 1 44967
0 44969 7 1 2 51796 79612
0 44970 5 1 1 44969
0 44971 7 1 2 14653 79211
0 44972 5 1 1 44971
0 44973 7 2 2 72467 79097
0 44974 7 2 2 44972 79614
0 44975 5 1 1 79616
0 44976 7 1 2 69539 79325
0 44977 5 1 1 44976
0 44978 7 1 2 70580 70820
0 44979 5 1 1 44978
0 44980 7 1 2 44977 44979
0 44981 5 1 1 44980
0 44982 7 1 2 58787 44981
0 44983 5 1 1 44982
0 44984 7 1 2 64202 71698
0 44985 5 1 1 44984
0 44986 7 1 2 44742 44985
0 44987 5 1 1 44986
0 44988 7 2 2 52027 63676
0 44989 5 1 1 79618
0 44990 7 1 2 44987 79619
0 44991 5 1 1 44990
0 44992 7 1 2 65479 75788
0 44993 7 1 2 71536 44992
0 44994 5 1 1 44993
0 44995 7 1 2 44991 44994
0 44996 5 1 1 44995
0 44997 7 1 2 53756 44996
0 44998 5 1 1 44997
0 44999 7 1 2 70672 44989
0 45000 5 1 1 44999
0 45001 7 1 2 67841 71519
0 45002 7 1 2 45000 45001
0 45003 5 1 1 45002
0 45004 7 1 2 44998 45003
0 45005 7 1 2 44983 45004
0 45006 5 1 1 45005
0 45007 7 2 2 67955 45006
0 45008 5 1 1 79620
0 45009 7 2 2 51661 73235
0 45010 7 1 2 78912 79622
0 45011 5 1 1 45010
0 45012 7 1 2 45008 45011
0 45013 5 1 1 45012
0 45014 7 1 2 51455 45013
0 45015 5 1 1 45014
0 45016 7 1 2 55585 79575
0 45017 5 1 1 45016
0 45018 7 1 2 71463 68563
0 45019 5 1 1 45018
0 45020 7 1 2 45017 45019
0 45021 5 1 1 45020
0 45022 7 1 2 52838 45021
0 45023 5 1 1 45022
0 45024 7 1 2 72139 79123
0 45025 5 1 1 45024
0 45026 7 1 2 68567 45025
0 45027 5 1 1 45026
0 45028 7 1 2 75904 45027
0 45029 5 1 1 45028
0 45030 7 1 2 79133 45029
0 45031 7 1 2 45023 45030
0 45032 5 2 1 45031
0 45033 7 2 2 51797 73083
0 45034 7 1 2 79624 79626
0 45035 5 1 1 45034
0 45036 7 1 2 45015 45035
0 45037 5 1 1 45036
0 45038 7 1 2 57690 45037
0 45039 5 1 1 45038
0 45040 7 1 2 44975 45039
0 45041 7 1 2 44970 45040
0 45042 5 1 1 45041
0 45043 7 1 2 61475 45042
0 45044 5 1 1 45043
0 45045 7 1 2 44830 45044
0 45046 7 1 2 44481 45045
0 45047 7 1 2 44125 45046
0 45048 5 1 1 45047
0 45049 7 1 2 50877 45048
0 45050 5 1 1 45049
0 45051 7 1 2 50878 69487
0 45052 5 1 1 45051
0 45053 7 1 2 57549 45052
0 45054 5 1 1 45053
0 45055 7 1 2 64111 45054
0 45056 5 1 1 45055
0 45057 7 1 2 49258 45056
0 45058 5 1 1 45057
0 45059 7 1 2 60061 74824
0 45060 5 1 1 45059
0 45061 7 1 2 45058 45060
0 45062 5 1 1 45061
0 45063 7 1 2 48274 45062
0 45064 5 1 1 45063
0 45065 7 1 2 59421 65866
0 45066 5 1 1 45065
0 45067 7 1 2 48275 45066
0 45068 5 1 1 45067
0 45069 7 1 2 59413 45068
0 45070 5 1 1 45069
0 45071 7 1 2 64010 45070
0 45072 5 1 1 45071
0 45073 7 1 2 50879 74026
0 45074 5 1 1 45073
0 45075 7 1 2 61274 45074
0 45076 5 1 1 45075
0 45077 7 1 2 45072 45076
0 45078 7 1 2 45064 45077
0 45079 5 1 1 45078
0 45080 7 1 2 58990 45079
0 45081 5 1 1 45080
0 45082 7 1 2 55965 71559
0 45083 5 1 1 45082
0 45084 7 1 2 61229 45083
0 45085 5 1 1 45084
0 45086 7 1 2 45081 45085
0 45087 5 1 1 45086
0 45088 7 1 2 56430 45087
0 45089 5 1 1 45088
0 45090 7 1 2 62590 62311
0 45091 5 1 1 45090
0 45092 7 1 2 74728 77826
0 45093 5 1 1 45092
0 45094 7 1 2 45091 45093
0 45095 5 1 1 45094
0 45096 7 1 2 56598 45095
0 45097 5 1 1 45096
0 45098 7 1 2 67712 76746
0 45099 7 1 2 78074 45098
0 45100 5 1 1 45099
0 45101 7 1 2 1375 45100
0 45102 5 1 1 45101
0 45103 7 1 2 58991 45102
0 45104 5 1 1 45103
0 45105 7 1 2 45097 45104
0 45106 5 1 1 45105
0 45107 7 1 2 48449 45106
0 45108 5 1 1 45107
0 45109 7 1 2 74717 78443
0 45110 5 1 1 45109
0 45111 7 1 2 61223 45110
0 45112 5 1 1 45111
0 45113 7 1 2 79526 45112
0 45114 5 1 1 45113
0 45115 7 1 2 65326 58992
0 45116 5 1 1 45115
0 45117 7 1 2 1928 45116
0 45118 5 1 1 45117
0 45119 7 1 2 62667 45118
0 45120 5 1 1 45119
0 45121 7 1 2 62789 61234
0 45122 5 1 1 45121
0 45123 7 1 2 77184 78445
0 45124 5 1 1 45123
0 45125 7 1 2 45122 45124
0 45126 7 1 2 45120 45125
0 45127 7 1 2 45114 45126
0 45128 7 1 2 45108 45127
0 45129 5 1 1 45128
0 45130 7 1 2 48019 45129
0 45131 5 1 1 45130
0 45132 7 1 2 61239 62671
0 45133 5 1 1 45132
0 45134 7 1 2 58949 58993
0 45135 5 1 1 45134
0 45136 7 1 2 61224 45135
0 45137 5 1 1 45136
0 45138 7 1 2 72082 45137
0 45139 5 1 1 45138
0 45140 7 1 2 45133 45139
0 45141 7 1 2 45131 45140
0 45142 5 1 1 45141
0 45143 7 1 2 55833 45142
0 45144 5 1 1 45143
0 45145 7 1 2 61078 78821
0 45146 5 1 1 45145
0 45147 7 1 2 56969 45146
0 45148 5 1 1 45147
0 45149 7 1 2 78182 45148
0 45150 5 1 1 45149
0 45151 7 1 2 49259 45150
0 45152 5 1 1 45151
0 45153 7 1 2 66708 74804
0 45154 5 1 1 45153
0 45155 7 1 2 45152 45154
0 45156 5 1 1 45155
0 45157 7 1 2 48276 45156
0 45158 5 1 1 45157
0 45159 7 1 2 56970 31098
0 45160 5 1 1 45159
0 45161 7 1 2 45158 45160
0 45162 5 1 1 45161
0 45163 7 1 2 58994 45162
0 45164 5 1 1 45163
0 45165 7 1 2 54113 71135
0 45166 5 1 1 45165
0 45167 7 1 2 61724 45166
0 45168 5 1 1 45167
0 45169 7 1 2 78446 45168
0 45170 5 1 1 45169
0 45171 7 1 2 63157 65882
0 45172 7 1 2 78441 45171
0 45173 5 1 1 45172
0 45174 7 1 2 61240 45173
0 45175 5 1 1 45174
0 45176 7 1 2 45170 45175
0 45177 5 1 1 45176
0 45178 7 1 2 61983 45177
0 45179 5 1 1 45178
0 45180 7 1 2 48020 75557
0 45181 5 1 1 45180
0 45182 7 1 2 1596 45181
0 45183 5 1 1 45182
0 45184 7 1 2 54114 45183
0 45185 5 1 1 45184
0 45186 7 1 2 50880 61278
0 45187 5 1 1 45186
0 45188 7 1 2 66774 45187
0 45189 5 1 1 45188
0 45190 7 1 2 74806 45189
0 45191 7 1 2 45185 45190
0 45192 5 1 1 45191
0 45193 7 1 2 61230 45192
0 45194 5 1 1 45193
0 45195 7 1 2 78388 45194
0 45196 7 1 2 45179 45195
0 45197 7 1 2 45164 45196
0 45198 7 1 2 45144 45197
0 45199 7 1 2 45089 45198
0 45200 5 1 1 45199
0 45201 7 2 2 69540 45200
0 45202 5 1 1 79628
0 45203 7 1 2 60440 72635
0 45204 5 1 1 45203
0 45205 7 1 2 70176 79276
0 45206 7 1 2 45204 45205
0 45207 5 1 1 45206
0 45208 7 1 2 78863 45207
0 45209 7 1 2 45202 45208
0 45210 5 1 1 45209
0 45211 7 1 2 51176 45210
0 45212 5 1 1 45211
0 45213 7 1 2 69874 77702
0 45214 5 1 1 45213
0 45215 7 1 2 78219 45214
0 45216 5 1 1 45215
0 45217 7 1 2 57691 45216
0 45218 5 1 1 45217
0 45219 7 1 2 54804 45218
0 45220 5 1 1 45219
0 45221 7 1 2 49138 60709
0 45222 5 1 1 45221
0 45223 7 1 2 1301 45222
0 45224 5 1 1 45223
0 45225 7 1 2 59317 45224
0 45226 5 1 1 45225
0 45227 7 1 2 54805 61992
0 45228 5 1 1 45227
0 45229 7 1 2 57692 45228
0 45230 7 1 2 45226 45229
0 45231 5 1 1 45230
0 45232 7 1 2 48021 45231
0 45233 5 1 1 45232
0 45234 7 1 2 56167 77164
0 45235 5 1 1 45234
0 45236 7 1 2 61650 45235
0 45237 5 1 1 45236
0 45238 7 1 2 48277 45237
0 45239 5 1 1 45238
0 45240 7 1 2 61878 76816
0 45241 5 1 1 45240
0 45242 7 1 2 48450 45241
0 45243 5 1 1 45242
0 45244 7 1 2 64475 61710
0 45245 7 1 2 77441 45244
0 45246 5 1 1 45245
0 45247 7 1 2 61764 74672
0 45248 5 1 1 45247
0 45249 7 1 2 74707 45248
0 45250 7 1 2 45246 45249
0 45251 7 1 2 45243 45250
0 45252 7 1 2 45239 45251
0 45253 7 1 2 45233 45252
0 45254 5 1 1 45253
0 45255 7 1 2 54415 45254
0 45256 5 1 1 45255
0 45257 7 1 2 45220 45256
0 45258 5 1 1 45257
0 45259 7 1 2 78367 45258
0 45260 5 1 1 45259
0 45261 7 2 2 59481 78812
0 45262 5 1 1 79630
0 45263 7 1 2 76207 79631
0 45264 5 1 1 45263
0 45265 7 1 2 54416 77580
0 45266 5 1 1 45265
0 45267 7 1 2 50881 45266
0 45268 5 1 1 45267
0 45269 7 1 2 64580 61243
0 45270 7 1 2 45268 45269
0 45271 5 1 1 45270
0 45272 7 1 2 78384 45271
0 45273 7 1 2 45264 45272
0 45274 7 2 2 45260 45273
0 45275 7 1 2 49820 7365
0 45276 5 1 1 45275
0 45277 7 1 2 52729 64357
0 45278 7 1 2 45262 45277
0 45279 5 1 1 45278
0 45280 7 1 2 53600 45279
0 45281 5 1 1 45280
0 45282 7 2 2 45276 45281
0 45283 5 1 1 79634
0 45284 7 1 2 49643 45283
0 45285 5 1 1 45284
0 45286 7 1 2 79632 45285
0 45287 5 1 1 45286
0 45288 7 1 2 55149 45287
0 45289 5 1 1 45288
0 45290 7 1 2 78392 45289
0 45291 5 1 1 45290
0 45292 7 1 2 69541 45291
0 45293 5 1 1 45292
0 45294 7 1 2 78864 78983
0 45295 5 1 1 45294
0 45296 7 1 2 78914 45295
0 45297 5 1 1 45296
0 45298 7 1 2 45293 45297
0 45299 7 1 2 45212 45298
0 45300 5 1 1 45299
0 45301 7 1 2 51662 45300
0 45302 5 1 1 45301
0 45303 7 1 2 52028 79042
0 45304 5 1 1 45303
0 45305 7 1 2 56168 60785
0 45306 5 1 1 45305
0 45307 7 1 2 56263 73533
0 45308 7 1 2 45306 45307
0 45309 5 1 1 45308
0 45310 7 1 2 45304 45309
0 45311 5 1 1 45310
0 45312 7 1 2 50561 45311
0 45313 5 1 1 45312
0 45314 7 1 2 73679 70428
0 45315 5 1 1 45314
0 45316 7 1 2 63550 45315
0 45317 5 1 1 45316
0 45318 7 1 2 56264 45317
0 45319 5 1 1 45318
0 45320 7 1 2 45313 45319
0 45321 5 2 1 45320
0 45322 7 1 2 78742 79636
0 45323 5 1 1 45322
0 45324 7 1 2 65533 60812
0 45325 5 2 1 45324
0 45326 7 1 2 79387 79638
0 45327 5 1 1 45326
0 45328 7 1 2 45323 45327
0 45329 5 1 1 45328
0 45330 7 1 2 56481 45329
0 45331 5 1 1 45330
0 45332 7 1 2 70673 73880
0 45333 5 1 1 45332
0 45334 7 1 2 52029 45333
0 45335 5 1 1 45334
0 45336 7 1 2 78681 45335
0 45337 5 1 1 45336
0 45338 7 1 2 50562 45337
0 45339 5 1 1 45338
0 45340 7 1 2 65480 59819
0 45341 7 1 2 76434 45340
0 45342 5 1 1 45341
0 45343 7 1 2 45339 45342
0 45344 5 1 1 45343
0 45345 7 1 2 57693 45344
0 45346 5 1 1 45345
0 45347 7 1 2 60441 78645
0 45348 5 1 1 45347
0 45349 7 2 2 56265 45348
0 45350 7 1 2 51177 79640
0 45351 5 1 1 45350
0 45352 7 1 2 45346 45351
0 45353 5 1 1 45352
0 45354 7 1 2 79388 45353
0 45355 5 1 1 45354
0 45356 7 1 2 56482 67021
0 45357 5 1 1 45356
0 45358 7 1 2 79144 45357
0 45359 5 1 1 45358
0 45360 7 1 2 79586 45359
0 45361 5 1 1 45360
0 45362 7 1 2 67646 73260
0 45363 5 1 1 45362
0 45364 7 1 2 45361 45363
0 45365 5 1 1 45364
0 45366 7 1 2 52839 45365
0 45367 5 1 1 45366
0 45368 7 2 2 76864 78262
0 45369 7 1 2 51663 71145
0 45370 7 1 2 79642 45369
0 45371 5 1 1 45370
0 45372 7 1 2 45367 45371
0 45373 5 2 1 45372
0 45374 7 1 2 73037 79644
0 45375 5 1 1 45374
0 45376 7 1 2 62744 63540
0 45377 5 1 1 45376
0 45378 7 1 2 52030 77327
0 45379 5 1 1 45378
0 45380 7 1 2 45377 45379
0 45381 5 1 1 45380
0 45382 7 1 2 50563 45381
0 45383 5 1 1 45382
0 45384 7 1 2 55715 79038
0 45385 5 1 1 45384
0 45386 7 1 2 45383 45385
0 45387 5 1 1 45386
0 45388 7 2 2 53757 79146
0 45389 7 1 2 45387 79646
0 45390 5 1 1 45389
0 45391 7 1 2 55716 73764
0 45392 5 1 1 45391
0 45393 7 1 2 70674 45392
0 45394 5 1 1 45393
0 45395 7 1 2 79389 45394
0 45396 5 1 1 45395
0 45397 7 1 2 63810 78979
0 45398 5 1 1 45397
0 45399 7 1 2 63551 45398
0 45400 5 2 1 45399
0 45401 7 1 2 79647 79648
0 45402 5 1 1 45401
0 45403 7 1 2 45396 45402
0 45404 5 2 1 45403
0 45405 7 1 2 73038 79650
0 45406 5 1 1 45405
0 45407 7 1 2 45390 45406
0 45408 5 1 1 45407
0 45409 7 1 2 57694 45408
0 45410 5 1 1 45409
0 45411 7 1 2 45375 45410
0 45412 7 1 2 45355 45411
0 45413 7 1 2 45331 45412
0 45414 5 1 1 45413
0 45415 7 1 2 62990 45414
0 45416 5 1 1 45415
0 45417 7 1 2 67793 70177
0 45418 5 1 1 45417
0 45419 7 1 2 39109 45418
0 45420 5 1 1 45419
0 45421 7 1 2 62503 45420
0 45422 5 1 1 45421
0 45423 7 1 2 70178 79390
0 45424 5 1 1 45423
0 45425 7 1 2 45422 45424
0 45426 5 3 1 45425
0 45427 7 2 2 51178 62745
0 45428 5 1 1 79655
0 45429 7 1 2 79652 79656
0 45430 5 1 1 45429
0 45431 7 1 2 56266 67647
0 45432 5 1 1 45431
0 45433 7 1 2 67803 45432
0 45434 5 2 1 45433
0 45435 7 1 2 62504 79657
0 45436 5 1 1 45435
0 45437 7 1 2 67191 77992
0 45438 5 1 1 45437
0 45439 7 1 2 45436 45438
0 45440 5 1 1 45439
0 45441 7 1 2 52840 45440
0 45442 5 1 1 45441
0 45443 7 1 2 70563 73813
0 45444 5 1 1 45443
0 45445 7 1 2 45442 45444
0 45446 5 1 1 45445
0 45447 7 1 2 61251 45446
0 45448 5 1 1 45447
0 45449 7 1 2 45430 45448
0 45450 5 1 1 45449
0 45451 7 1 2 50564 45450
0 45452 5 1 1 45451
0 45453 7 1 2 59782 71178
0 45454 7 1 2 79653 45453
0 45455 5 1 1 45454
0 45456 7 1 2 62505 60648
0 45457 5 1 1 45456
0 45458 7 1 2 71126 45457
0 45459 5 1 1 45458
0 45460 7 1 2 67866 45459
0 45461 5 1 1 45460
0 45462 7 1 2 56267 78013
0 45463 5 1 1 45462
0 45464 7 2 2 55717 69542
0 45465 7 1 2 63576 75348
0 45466 7 1 2 79659 45465
0 45467 5 1 1 45466
0 45468 7 1 2 45463 45467
0 45469 7 1 2 45461 45468
0 45470 5 1 1 45469
0 45471 7 1 2 51664 45470
0 45472 5 1 1 45471
0 45473 7 2 2 73651 78059
0 45474 7 1 2 79649 79661
0 45475 5 1 1 45474
0 45476 7 2 2 45472 45475
0 45477 5 1 1 79663
0 45478 7 1 2 73039 45477
0 45479 5 1 1 45478
0 45480 7 1 2 45455 45479
0 45481 7 1 2 45452 45480
0 45482 5 1 1 45481
0 45483 7 1 2 57695 45482
0 45484 5 1 1 45483
0 45485 7 1 2 61144 74901
0 45486 5 1 1 45485
0 45487 7 1 2 52207 45486
0 45488 5 1 1 45487
0 45489 7 1 2 55966 70185
0 45490 5 1 1 45489
0 45491 7 1 2 55150 45490
0 45492 7 1 2 45488 45491
0 45493 5 1 1 45492
0 45494 7 1 2 56268 59167
0 45495 7 1 2 45493 45494
0 45496 5 1 1 45495
0 45497 7 1 2 63541 72631
0 45498 5 1 1 45497
0 45499 7 1 2 75387 45498
0 45500 7 1 2 45496 45499
0 45501 5 1 1 45500
0 45502 7 1 2 79662 45501
0 45503 5 1 1 45502
0 45504 7 1 2 45484 45503
0 45505 7 1 2 45416 45504
0 45506 7 1 2 45302 45505
0 45507 5 1 1 45506
0 45508 7 1 2 68965 45507
0 45509 5 1 1 45508
0 45510 7 1 2 52031 76742
0 45511 5 1 1 45510
0 45512 7 1 2 70842 45511
0 45513 5 1 1 45512
0 45514 7 1 2 68883 45513
0 45515 5 1 1 45514
0 45516 7 1 2 78635 45515
0 45517 5 1 1 45516
0 45518 7 1 2 79031 45517
0 45519 5 1 1 45518
0 45520 7 1 2 50565 77782
0 45521 5 1 1 45520
0 45522 7 2 2 79106 45521
0 45523 5 2 1 79665
0 45524 7 1 2 70331 79667
0 45525 5 1 1 45524
0 45526 7 1 2 77788 79107
0 45527 5 1 1 45526
0 45528 7 1 2 54806 45527
0 45529 5 1 1 45528
0 45530 7 1 2 75471 45529
0 45531 5 1 1 45530
0 45532 7 1 2 64203 45531
0 45533 5 1 1 45532
0 45534 7 1 2 75255 45533
0 45535 5 1 1 45534
0 45536 7 1 2 53601 45535
0 45537 5 1 1 45536
0 45538 7 1 2 45525 45537
0 45539 5 1 1 45538
0 45540 7 1 2 51456 45539
0 45541 5 1 1 45540
0 45542 7 1 2 45519 45541
0 45543 5 1 1 45542
0 45544 7 1 2 53758 45543
0 45545 5 1 1 45544
0 45546 7 2 2 51457 79668
0 45547 7 1 2 79020 79669
0 45548 5 1 1 45547
0 45549 7 1 2 45545 45548
0 45550 5 1 1 45549
0 45551 7 1 2 52841 45550
0 45552 5 1 1 45551
0 45553 7 1 2 79085 79670
0 45554 5 1 1 45553
0 45555 7 1 2 45552 45554
0 45556 5 1 1 45555
0 45557 7 1 2 55586 57696
0 45558 7 1 2 45556 45557
0 45559 5 1 1 45558
0 45560 7 1 2 72717 78965
0 45561 5 1 1 45560
0 45562 7 1 2 75911 45561
0 45563 5 1 1 45562
0 45564 7 1 2 51179 45563
0 45565 5 1 1 45564
0 45566 7 1 2 52032 79060
0 45567 5 1 1 45566
0 45568 7 1 2 45565 45567
0 45569 5 1 1 45568
0 45570 7 1 2 51458 45569
0 45571 5 1 1 45570
0 45572 7 1 2 52033 79062
0 45573 5 1 1 45572
0 45574 7 1 2 55587 45573
0 45575 7 1 2 45571 45574
0 45576 5 1 1 45575
0 45577 7 1 2 58574 77225
0 45578 5 1 1 45577
0 45579 7 1 2 61504 66669
0 45580 5 1 1 45579
0 45581 7 1 2 45578 45580
0 45582 5 1 1 45581
0 45583 7 1 2 50566 45582
0 45584 5 1 1 45583
0 45585 7 1 2 66060 45584
0 45586 5 2 1 45585
0 45587 7 1 2 68408 79671
0 45588 5 1 1 45587
0 45589 7 1 2 67571 78615
0 45590 5 1 1 45589
0 45591 7 1 2 45588 45590
0 45592 5 2 1 45591
0 45593 7 1 2 71464 79673
0 45594 5 1 1 45593
0 45595 7 1 2 67705 41019
0 45596 5 1 1 45595
0 45597 7 1 2 78995 45596
0 45598 5 1 1 45597
0 45599 7 1 2 72173 79024
0 45600 5 1 1 45599
0 45601 7 1 2 51665 45600
0 45602 7 1 2 45598 45601
0 45603 7 1 2 45594 45602
0 45604 5 1 1 45603
0 45605 7 1 2 45576 45604
0 45606 5 1 1 45605
0 45607 7 1 2 49984 45606
0 45608 5 1 1 45607
0 45609 7 1 2 52034 78608
0 45610 5 1 1 45609
0 45611 7 1 2 58734 40830
0 45612 5 1 1 45611
0 45613 7 1 2 51180 45612
0 45614 5 1 1 45613
0 45615 7 1 2 49821 45614
0 45616 7 1 2 45610 45615
0 45617 5 1 1 45616
0 45618 7 1 2 59951 79045
0 45619 5 1 1 45618
0 45620 7 1 2 70081 45619
0 45621 5 1 1 45620
0 45622 7 1 2 51459 45621
0 45623 7 1 2 45617 45622
0 45624 5 1 1 45623
0 45625 7 1 2 78719 79074
0 45626 5 1 1 45625
0 45627 7 1 2 45626 78948
0 45628 5 1 1 45627
0 45629 7 1 2 50309 79184
0 45630 5 1 1 45629
0 45631 7 1 2 45628 45630
0 45632 5 1 1 45631
0 45633 7 1 2 58788 45632
0 45634 5 1 1 45633
0 45635 7 2 2 59159 63666
0 45636 7 1 2 49644 79675
0 45637 5 1 1 45636
0 45638 7 1 2 41140 45637
0 45639 5 1 1 45638
0 45640 7 1 2 78949 45639
0 45641 5 1 1 45640
0 45642 7 1 2 71520 79036
0 45643 5 1 1 45642
0 45644 7 1 2 45641 45643
0 45645 5 1 1 45644
0 45646 7 1 2 55425 45645
0 45647 5 1 1 45646
0 45648 7 1 2 45634 45647
0 45649 7 1 2 45624 45648
0 45650 5 1 1 45649
0 45651 7 1 2 55588 45650
0 45652 5 1 1 45651
0 45653 7 1 2 70295 78671
0 45654 5 1 1 45653
0 45655 7 1 2 54807 75004
0 45656 5 1 1 45655
0 45657 7 1 2 45654 45656
0 45658 5 1 1 45657
0 45659 7 1 2 53602 45658
0 45660 5 1 1 45659
0 45661 7 1 2 79050 45660
0 45662 5 1 1 45661
0 45663 7 1 2 66301 45662
0 45664 5 1 1 45663
0 45665 7 1 2 52035 73534
0 45666 7 1 2 67743 45665
0 45667 5 1 1 45666
0 45668 7 1 2 45664 45667
0 45669 5 1 1 45668
0 45670 7 1 2 66670 45669
0 45671 5 1 1 45670
0 45672 7 1 2 53759 45671
0 45673 7 1 2 45652 45672
0 45674 5 1 1 45673
0 45675 7 1 2 52842 45674
0 45676 7 1 2 45608 45675
0 45677 5 1 1 45676
0 45678 7 1 2 79543 79674
0 45679 5 1 1 45678
0 45680 7 1 2 71296 78658
0 45681 7 1 2 79032 45680
0 45682 5 1 1 45681
0 45683 7 1 2 79104 79666
0 45684 5 3 1 45683
0 45685 7 1 2 66615 79677
0 45686 7 1 2 78907 45685
0 45687 5 1 1 45686
0 45688 7 1 2 45682 45687
0 45689 7 1 2 45679 45688
0 45690 5 1 1 45689
0 45691 7 1 2 51666 45690
0 45692 5 1 1 45691
0 45693 7 1 2 78902 78966
0 45694 5 1 1 45693
0 45695 7 1 2 78940 45694
0 45696 5 1 1 45695
0 45697 7 1 2 51181 45696
0 45698 5 1 1 45697
0 45699 7 1 2 52036 79078
0 45700 5 1 1 45699
0 45701 7 1 2 45698 45700
0 45702 5 1 1 45701
0 45703 7 1 2 51460 45702
0 45704 5 1 1 45703
0 45705 7 1 2 52037 79081
0 45706 7 1 2 79676 45705
0 45707 7 1 2 78505 45706
0 45708 5 1 1 45707
0 45709 7 1 2 45704 45708
0 45710 5 1 1 45709
0 45711 7 1 2 65744 45710
0 45712 5 1 1 45711
0 45713 7 1 2 45692 45712
0 45714 7 1 2 45677 45713
0 45715 7 1 2 45559 45714
0 45716 5 2 1 45715
0 45717 7 1 2 51798 79680
0 45718 5 1 1 45717
0 45719 7 1 2 59952 79170
0 45720 5 1 1 45719
0 45721 7 1 2 78244 78989
0 45722 5 1 1 45721
0 45723 7 1 2 55426 45722
0 45724 7 1 2 45720 45723
0 45725 5 1 1 45724
0 45726 7 1 2 10630 79151
0 45727 5 2 1 45726
0 45728 7 2 2 52038 79682
0 45729 7 1 2 78970 79684
0 45730 5 1 1 45729
0 45731 7 1 2 51461 41621
0 45732 7 1 2 45730 45731
0 45733 5 1 1 45732
0 45734 7 1 2 51799 45733
0 45735 7 1 2 45725 45734
0 45736 5 1 1 45735
0 45737 7 1 2 52585 73652
0 45738 7 1 2 68530 45737
0 45739 7 1 2 77968 45738
0 45740 7 1 2 79685 45739
0 45741 5 1 1 45740
0 45742 7 1 2 45736 45741
0 45743 5 1 1 45742
0 45744 7 1 2 51667 57697
0 45745 7 1 2 45743 45744
0 45746 5 1 1 45745
0 45747 7 1 2 69816 79098
0 45748 7 1 2 79678 45747
0 45749 5 1 1 45748
0 45750 7 2 2 45746 45749
0 45751 5 1 1 79686
0 45752 7 1 2 45718 79687
0 45753 5 1 1 45752
0 45754 7 1 2 70220 45753
0 45755 5 1 1 45754
0 45756 7 1 2 60429 78973
0 45757 5 1 1 45756
0 45758 7 1 2 72632 79522
0 45759 5 1 1 45758
0 45760 7 1 2 45757 45759
0 45761 5 1 1 45760
0 45762 7 1 2 51182 45761
0 45763 5 1 1 45762
0 45764 7 1 2 40896 45763
0 45765 5 1 1 45764
0 45766 7 1 2 55967 45765
0 45767 5 1 1 45766
0 45768 7 1 2 60430 78990
0 45769 5 1 1 45768
0 45770 7 1 2 65358 70451
0 45771 7 1 2 79168 45770
0 45772 5 1 1 45771
0 45773 7 1 2 45769 45772
0 45774 5 1 1 45773
0 45775 7 1 2 55427 45774
0 45776 5 1 1 45775
0 45777 7 1 2 51183 40509
0 45778 7 1 2 78974 45777
0 45779 5 1 1 45778
0 45780 7 1 2 45776 45779
0 45781 5 1 1 45780
0 45782 7 1 2 57698 45781
0 45783 5 1 1 45782
0 45784 7 1 2 71360 78871
0 45785 5 1 1 45784
0 45786 7 1 2 51668 45785
0 45787 7 1 2 45783 45786
0 45788 7 1 2 45767 45787
0 45789 5 1 1 45788
0 45790 7 1 2 68599 72633
0 45791 5 1 1 45790
0 45792 7 1 2 78998 45791
0 45793 5 1 1 45792
0 45794 7 1 2 57699 45793
0 45795 5 1 1 45794
0 45796 7 1 2 50310 79182
0 45797 5 1 1 45796
0 45798 7 1 2 68608 45797
0 45799 5 1 1 45798
0 45800 7 1 2 55718 45799
0 45801 5 1 1 45800
0 45802 7 1 2 78700 45801
0 45803 5 1 1 45802
0 45804 7 1 2 56668 45803
0 45805 5 1 1 45804
0 45806 7 1 2 24955 45805
0 45807 5 1 1 45806
0 45808 7 1 2 72662 45807
0 45809 5 1 1 45808
0 45810 7 1 2 38901 45809
0 45811 7 1 2 45795 45810
0 45812 5 1 1 45811
0 45813 7 1 2 58789 45812
0 45814 5 1 1 45813
0 45815 7 1 2 61534 73680
0 45816 7 1 2 63390 45815
0 45817 5 1 1 45816
0 45818 7 1 2 63552 45817
0 45819 5 1 1 45818
0 45820 7 1 2 76504 45819
0 45821 5 1 1 45820
0 45822 7 1 2 59755 71052
0 45823 5 1 1 45822
0 45824 7 1 2 50567 45823
0 45825 5 1 1 45824
0 45826 7 1 2 73040 76803
0 45827 5 1 1 45826
0 45828 7 1 2 71444 45827
0 45829 7 1 2 45825 45828
0 45830 5 1 1 45829
0 45831 7 1 2 68706 78656
0 45832 7 1 2 45830 45831
0 45833 5 1 1 45832
0 45834 7 1 2 45821 45833
0 45835 5 1 1 45834
0 45836 7 1 2 52351 45835
0 45837 5 1 1 45836
0 45838 7 1 2 64600 75066
0 45839 5 1 1 45838
0 45840 7 1 2 67818 45839
0 45841 5 1 1 45840
0 45842 7 1 2 51184 45841
0 45843 5 1 1 45842
0 45844 7 1 2 73357 78653
0 45845 7 1 2 72629 45844
0 45846 5 1 1 45845
0 45847 7 1 2 45843 45846
0 45848 7 1 2 45837 45847
0 45849 7 1 2 45814 45848
0 45850 5 1 1 45849
0 45851 7 1 2 69543 45850
0 45852 5 1 1 45851
0 45853 7 1 2 61145 72627
0 45854 5 1 1 45853
0 45855 7 1 2 59801 45854
0 45856 5 1 1 45855
0 45857 7 1 2 65354 78919
0 45858 5 1 1 45857
0 45859 7 1 2 55968 45858
0 45860 5 1 1 45859
0 45861 7 1 2 55151 45860
0 45862 7 1 2 45856 45861
0 45863 5 1 1 45862
0 45864 7 1 2 49985 79568
0 45865 5 1 1 45864
0 45866 7 1 2 79089 45865
0 45867 5 1 1 45866
0 45868 7 1 2 51462 45867
0 45869 7 1 2 45863 45868
0 45870 5 1 1 45869
0 45871 7 1 2 55589 45870
0 45872 7 1 2 45852 45871
0 45873 5 1 1 45872
0 45874 7 2 2 45789 45873
0 45875 7 1 2 51800 79688
0 45876 5 1 1 45875
0 45877 7 1 2 60442 78922
0 45878 5 1 1 45877
0 45879 7 1 2 59925 79615
0 45880 7 2 2 45878 45879
0 45881 5 1 1 79690
0 45882 7 1 2 45876 45881
0 45883 5 1 1 45882
0 45884 7 1 2 57069 45883
0 45885 5 1 1 45884
0 45886 7 1 2 22257 79002
0 45887 5 1 1 45886
0 45888 7 1 2 74906 75005
0 45889 5 1 1 45888
0 45890 7 1 2 45887 45889
0 45891 5 1 1 45890
0 45892 7 1 2 53603 45891
0 45893 5 1 1 45892
0 45894 7 1 2 60431 79000
0 45895 5 1 1 45894
0 45896 7 1 2 45893 45895
0 45897 5 1 1 45896
0 45898 7 1 2 54808 45897
0 45899 5 1 1 45898
0 45900 7 1 2 49822 58796
0 45901 7 1 2 75171 45900
0 45902 5 1 1 45901
0 45903 7 1 2 76010 45902
0 45904 5 1 1 45903
0 45905 7 1 2 51463 45904
0 45906 5 1 1 45905
0 45907 7 1 2 45899 45906
0 45908 5 1 1 45907
0 45909 7 1 2 53760 45908
0 45910 5 1 1 45909
0 45911 7 1 2 49986 70598
0 45912 7 1 2 75168 45911
0 45913 7 1 2 71376 75978
0 45914 7 1 2 45912 45913
0 45915 5 1 1 45914
0 45916 7 1 2 45910 45915
0 45917 5 1 1 45916
0 45918 7 1 2 52843 45917
0 45919 5 1 1 45918
0 45920 7 1 2 66892 70513
0 45921 7 1 2 79086 45920
0 45922 5 1 1 45921
0 45923 7 1 2 45919 45922
0 45924 5 1 1 45923
0 45925 7 2 2 67956 45924
0 45926 5 1 1 79692
0 45927 7 1 2 73615 79102
0 45928 5 1 1 45927
0 45929 7 1 2 55152 77566
0 45930 5 1 1 45929
0 45931 7 1 2 45928 45930
0 45932 5 1 1 45931
0 45933 7 1 2 73699 45932
0 45934 5 1 1 45933
0 45935 7 1 2 60824 78054
0 45936 5 1 1 45935
0 45937 7 1 2 55153 67050
0 45938 5 1 1 45937
0 45939 7 1 2 45936 45938
0 45940 5 1 1 45939
0 45941 7 1 2 48979 45940
0 45942 5 1 1 45941
0 45943 7 1 2 67572 67842
0 45944 5 1 1 45943
0 45945 7 1 2 45942 45944
0 45946 5 1 1 45945
0 45947 7 1 2 58790 45946
0 45948 5 1 1 45947
0 45949 7 1 2 45934 45948
0 45950 5 1 1 45949
0 45951 7 1 2 51464 45950
0 45952 5 1 1 45951
0 45953 7 3 2 63891 60786
0 45954 5 2 1 79694
0 45955 7 1 2 78993 79697
0 45956 5 1 1 45955
0 45957 7 2 2 45952 45956
0 45958 5 1 1 79699
0 45959 7 1 2 79587 79609
0 45960 5 1 1 45959
0 45961 7 2 2 55719 75077
0 45962 7 1 2 49823 79701
0 45963 5 1 1 45962
0 45964 7 1 2 41017 45963
0 45965 5 1 1 45964
0 45966 7 1 2 49987 45965
0 45967 5 1 1 45966
0 45968 7 2 2 64576 73308
0 45969 5 1 1 79703
0 45970 7 1 2 45967 45969
0 45971 5 1 1 45970
0 45972 7 1 2 52844 45971
0 45973 5 1 1 45972
0 45974 7 1 2 79611 45973
0 45975 7 1 2 45960 45974
0 45976 5 1 1 45975
0 45977 7 1 2 73041 45976
0 45978 5 1 1 45977
0 45979 7 1 2 79700 45978
0 45980 5 1 1 45979
0 45981 7 1 2 51801 45980
0 45982 5 1 1 45981
0 45983 7 1 2 61049 63667
0 45984 7 1 2 73276 45983
0 45985 7 1 2 69367 79479
0 45986 7 1 2 45984 45985
0 45987 5 2 1 45986
0 45988 7 2 2 58844 73658
0 45989 7 2 2 73042 79707
0 45990 7 1 2 50113 68531
0 45991 7 1 2 74441 45990
0 45992 7 1 2 79709 45991
0 45993 5 1 1 45992
0 45994 7 1 2 79705 45993
0 45995 7 1 2 45982 45994
0 45996 5 1 1 45995
0 45997 7 1 2 51669 45996
0 45998 5 1 1 45997
0 45999 7 1 2 45926 45998
0 46000 5 1 1 45999
0 46001 7 1 2 66671 46000
0 46002 5 1 1 46001
0 46003 7 1 2 50073 46002
0 46004 7 1 2 45885 46003
0 46005 7 1 2 45755 46004
0 46006 7 1 2 45509 46005
0 46007 7 1 2 45050 46006
0 46008 7 1 2 43740 46007
0 46009 7 1 2 41748 46008
0 46010 7 1 2 40792 46009
0 46011 5 1 1 46010
0 46012 7 1 2 39738 46011
0 46013 5 1 1 46012
0 46014 7 1 2 52869 46013
0 46015 5 1 1 46014
0 46016 7 1 2 53794 79287
0 46017 5 1 1 46016
0 46018 7 1 2 59626 77319
0 46019 5 1 1 46018
0 46020 7 1 2 70383 46019
0 46021 5 1 1 46020
0 46022 7 1 2 58462 9238
0 46023 5 2 1 46022
0 46024 7 1 2 50311 77773
0 46025 5 1 1 46024
0 46026 7 1 2 63772 72935
0 46027 7 1 2 77442 46026
0 46028 7 1 2 46025 46027
0 46029 7 1 2 79711 46028
0 46030 5 1 1 46029
0 46031 7 1 2 57266 46030
0 46032 5 1 1 46031
0 46033 7 1 2 46021 46032
0 46034 5 1 1 46033
0 46035 7 1 2 52465 46034
0 46036 5 1 1 46035
0 46037 7 1 2 79454 46036
0 46038 5 1 1 46037
0 46039 7 1 2 50882 46038
0 46040 5 1 1 46039
0 46041 7 1 2 79456 46040
0 46042 5 1 1 46041
0 46043 7 1 2 71476 46042
0 46044 5 1 1 46043
0 46045 7 1 2 65797 71952
0 46046 7 1 2 79196 46045
0 46047 5 1 1 46046
0 46048 7 1 2 50883 46047
0 46049 5 1 1 46048
0 46050 7 1 2 50568 65829
0 46051 5 1 1 46050
0 46052 7 1 2 72582 79203
0 46053 7 1 2 46051 46052
0 46054 7 1 2 70288 79712
0 46055 7 1 2 46053 46054
0 46056 5 1 1 46055
0 46057 7 1 2 52466 46056
0 46058 5 1 1 46057
0 46059 7 1 2 46049 46058
0 46060 5 1 1 46059
0 46061 7 1 2 62506 46060
0 46062 5 1 1 46061
0 46063 7 1 2 46044 46062
0 46064 5 1 1 46063
0 46065 7 1 2 51465 46064
0 46066 5 1 1 46065
0 46067 7 1 2 70695 76134
0 46068 5 1 1 46067
0 46069 7 1 2 52352 70221
0 46070 5 1 1 46069
0 46071 7 1 2 24608 46070
0 46072 5 1 1 46071
0 46073 7 1 2 52039 46072
0 46074 5 1 1 46073
0 46075 7 1 2 48451 9425
0 46076 5 1 1 46075
0 46077 7 1 2 79267 46076
0 46078 5 1 1 46077
0 46079 7 1 2 29039 46078
0 46080 7 1 2 46074 46079
0 46081 5 1 1 46080
0 46082 7 1 2 53136 46081
0 46083 5 1 1 46082
0 46084 7 1 2 46068 46083
0 46085 5 1 1 46084
0 46086 7 1 2 50569 46085
0 46087 5 1 1 46086
0 46088 7 1 2 55969 77954
0 46089 5 1 1 46088
0 46090 7 1 2 46087 46089
0 46091 5 1 1 46090
0 46092 7 1 2 59038 76454
0 46093 7 1 2 46091 46092
0 46094 5 1 1 46093
0 46095 7 1 2 46066 46094
0 46096 5 1 1 46095
0 46097 7 1 2 53257 46096
0 46098 5 1 1 46097
0 46099 7 1 2 73177 79278
0 46100 5 1 1 46099
0 46101 7 1 2 70696 72747
0 46102 5 1 1 46101
0 46103 7 1 2 46100 46102
0 46104 5 1 1 46103
0 46105 7 1 2 58463 46104
0 46106 5 1 1 46105
0 46107 7 1 2 57700 60737
0 46108 5 1 1 46107
0 46109 7 1 2 74899 46108
0 46110 5 1 1 46109
0 46111 7 1 2 79279 46110
0 46112 5 1 1 46111
0 46113 7 1 2 58896 71047
0 46114 5 1 1 46113
0 46115 7 1 2 10275 46114
0 46116 5 1 1 46115
0 46117 7 1 2 53137 46116
0 46118 5 1 1 46117
0 46119 7 1 2 65012 72650
0 46120 5 1 1 46119
0 46121 7 1 2 59666 78263
0 46122 5 1 1 46121
0 46123 7 1 2 60274 72651
0 46124 5 1 1 46123
0 46125 7 1 2 46122 46124
0 46126 5 1 1 46125
0 46127 7 1 2 52040 46126
0 46128 5 1 1 46127
0 46129 7 1 2 46120 46128
0 46130 7 1 2 46118 46129
0 46131 7 1 2 46112 46130
0 46132 7 1 2 46106 46131
0 46133 5 1 1 46132
0 46134 7 1 2 53028 46133
0 46135 5 1 1 46134
0 46136 7 1 2 64970 61862
0 46137 7 1 2 62165 46136
0 46138 5 1 1 46137
0 46139 7 1 2 51185 46138
0 46140 5 1 1 46139
0 46141 7 1 2 46135 46140
0 46142 5 1 1 46141
0 46143 7 1 2 79552 46142
0 46144 5 1 1 46143
0 46145 7 1 2 66616 72990
0 46146 5 1 1 46145
0 46147 7 1 2 55428 71593
0 46148 5 1 1 46147
0 46149 7 1 2 70421 46148
0 46150 5 1 1 46149
0 46151 7 1 2 51466 71095
0 46152 5 1 1 46151
0 46153 7 1 2 46150 46152
0 46154 5 1 1 46153
0 46155 7 1 2 52730 73445
0 46156 7 1 2 46154 46155
0 46157 5 1 1 46156
0 46158 7 1 2 46146 46157
0 46159 5 1 1 46158
0 46160 7 1 2 62991 79446
0 46161 7 1 2 46159 46160
0 46162 5 1 1 46161
0 46163 7 1 2 46144 46162
0 46164 7 1 2 46098 46163
0 46165 5 1 1 46164
0 46166 7 7 2 71342 72192
0 46167 7 1 2 46165 79713
0 46168 5 1 1 46167
0 46169 7 1 2 46017 46168
0 46170 5 1 1 46169
0 46171 7 1 2 51802 46170
0 46172 5 1 1 46171
0 46173 7 1 2 58823 76765
0 46174 5 1 1 46173
0 46175 7 1 2 1905 46174
0 46176 5 1 1 46175
0 46177 7 1 2 52910 46176
0 46178 5 1 1 46177
0 46179 7 1 2 50114 74270
0 46180 5 1 1 46179
0 46181 7 1 2 46178 46180
0 46182 5 1 1 46181
0 46183 7 1 2 52353 46182
0 46184 5 1 1 46183
0 46185 7 1 2 63240 74572
0 46186 5 1 1 46185
0 46187 7 1 2 46184 46186
0 46188 5 1 1 46187
0 46189 7 1 2 52208 46188
0 46190 5 1 1 46189
0 46191 7 1 2 66258 77915
0 46192 7 1 2 62230 46191
0 46193 5 1 1 46192
0 46194 7 1 2 46190 46193
0 46195 5 1 1 46194
0 46196 7 1 2 52041 46195
0 46197 5 1 1 46196
0 46198 7 1 2 74271 79506
0 46199 5 1 1 46198
0 46200 7 1 2 46197 46199
0 46201 5 1 1 46200
0 46202 7 1 2 78603 46201
0 46203 5 1 1 46202
0 46204 7 1 2 53029 78311
0 46205 5 1 1 46204
0 46206 7 1 2 25267 46205
0 46207 5 2 1 46206
0 46208 7 1 2 52209 79720
0 46209 5 1 1 46208
0 46210 7 1 2 52731 72652
0 46211 5 1 1 46210
0 46212 7 1 2 46209 46211
0 46213 5 1 1 46212
0 46214 7 1 2 50312 46213
0 46215 5 1 1 46214
0 46216 7 1 2 21802 46215
0 46217 5 1 1 46216
0 46218 7 1 2 58464 46217
0 46219 5 1 1 46218
0 46220 7 1 2 52732 70422
0 46221 5 1 1 46220
0 46222 7 1 2 14892 46221
0 46223 5 1 1 46222
0 46224 7 1 2 62020 46223
0 46225 5 1 1 46224
0 46226 7 1 2 52354 60361
0 46227 5 1 1 46226
0 46228 7 1 2 60082 46227
0 46229 5 1 1 46228
0 46230 7 1 2 78312 46229
0 46231 5 1 1 46230
0 46232 7 1 2 46225 46231
0 46233 5 1 1 46232
0 46234 7 1 2 50313 46233
0 46235 5 1 1 46234
0 46236 7 1 2 52733 72768
0 46237 5 1 1 46236
0 46238 7 1 2 59953 79721
0 46239 5 1 1 46238
0 46240 7 1 2 73366 46239
0 46241 5 1 1 46240
0 46242 7 1 2 61194 46241
0 46243 5 1 1 46242
0 46244 7 1 2 46237 46243
0 46245 7 1 2 46235 46244
0 46246 7 1 2 46219 46245
0 46247 5 1 1 46246
0 46248 7 1 2 49824 46247
0 46249 5 1 1 46248
0 46250 7 1 2 46203 46249
0 46251 5 1 1 46250
0 46252 7 1 2 51186 46251
0 46253 5 1 1 46252
0 46254 7 1 2 57701 75397
0 46255 5 1 1 46254
0 46256 7 1 2 54115 46255
0 46257 5 1 1 46256
0 46258 7 1 2 74552 79337
0 46259 5 1 1 46258
0 46260 7 1 2 46257 46259
0 46261 5 1 1 46260
0 46262 7 1 2 64011 46261
0 46263 5 1 1 46262
0 46264 7 1 2 79356 46263
0 46265 5 1 1 46264
0 46266 7 1 2 68609 46265
0 46267 5 1 1 46266
0 46268 7 1 2 52734 46267
0 46269 5 1 1 46268
0 46270 7 1 2 46253 46269
0 46271 5 1 1 46270
0 46272 7 1 2 53761 46271
0 46273 5 1 1 46272
0 46274 7 1 2 32646 79415
0 46275 5 2 1 46274
0 46276 7 1 2 78057 79722
0 46277 5 1 1 46276
0 46278 7 1 2 46273 46277
0 46279 5 1 1 46278
0 46280 7 1 2 52845 46279
0 46281 5 1 1 46280
0 46282 7 1 2 62507 72941
0 46283 7 1 2 69291 46282
0 46284 7 1 2 79723 46283
0 46285 5 1 1 46284
0 46286 7 1 2 46281 46285
0 46287 5 1 1 46286
0 46288 7 1 2 69187 46287
0 46289 5 1 1 46288
0 46290 7 5 2 53795 67867
0 46291 7 3 2 55429 79724
0 46292 5 1 1 79729
0 46293 7 2 2 62992 79730
0 46294 7 1 2 71158 77994
0 46295 5 1 1 46294
0 46296 7 1 2 55154 46295
0 46297 5 1 1 46296
0 46298 7 1 2 52355 46297
0 46299 5 1 1 46298
0 46300 7 1 2 51187 75416
0 46301 5 1 1 46300
0 46302 7 1 2 49383 46301
0 46303 5 1 1 46302
0 46304 7 1 2 79437 46303
0 46305 5 1 1 46304
0 46306 7 1 2 46299 46305
0 46307 5 1 1 46306
0 46308 7 1 2 79732 46307
0 46309 5 1 1 46308
0 46310 7 3 2 67868 69933
0 46311 7 1 2 62274 79734
0 46312 5 1 1 46311
0 46313 7 1 2 61505 75337
0 46314 7 1 2 79372 46313
0 46315 5 1 1 46314
0 46316 7 1 2 46312 46315
0 46317 5 1 1 46316
0 46318 7 1 2 53030 46317
0 46319 5 1 1 46318
0 46320 7 1 2 76564 79735
0 46321 5 1 1 46320
0 46322 7 1 2 46319 46321
0 46323 5 1 1 46322
0 46324 7 1 2 53796 46323
0 46325 5 1 1 46324
0 46326 7 1 2 58845 75637
0 46327 7 1 2 75083 46326
0 46328 7 1 2 79209 46327
0 46329 5 1 1 46328
0 46330 7 1 2 46325 46329
0 46331 5 1 1 46330
0 46332 7 1 2 53138 46331
0 46333 5 1 1 46332
0 46334 7 2 2 53797 50115
0 46335 7 1 2 63588 79737
0 46336 7 1 2 79736 46335
0 46337 5 1 1 46336
0 46338 7 1 2 46333 46337
0 46339 5 1 1 46338
0 46340 7 1 2 52356 46339
0 46341 5 1 1 46340
0 46342 7 1 2 52042 79409
0 46343 5 1 1 46342
0 46344 7 1 2 49825 65309
0 46345 5 1 1 46344
0 46346 7 1 2 46343 46345
0 46347 5 1 1 46346
0 46348 7 1 2 79725 46347
0 46349 5 1 1 46348
0 46350 7 1 2 46341 46349
0 46351 5 1 1 46350
0 46352 7 1 2 50314 46351
0 46353 5 1 1 46352
0 46354 7 1 2 15669 72145
0 46355 5 4 1 46354
0 46356 7 1 2 52735 75417
0 46357 5 1 1 46356
0 46358 7 1 2 53139 71230
0 46359 7 1 2 76773 46358
0 46360 5 1 1 46359
0 46361 7 1 2 46357 46360
0 46362 5 1 1 46361
0 46363 7 1 2 71159 46362
0 46364 5 1 1 46363
0 46365 7 1 2 75341 46364
0 46366 5 1 1 46365
0 46367 7 1 2 79739 46366
0 46368 5 1 1 46367
0 46369 7 1 2 67573 72778
0 46370 5 1 1 46369
0 46371 7 1 2 73595 46370
0 46372 5 1 1 46371
0 46373 7 1 2 57702 46372
0 46374 5 1 1 46373
0 46375 7 1 2 60876 79261
0 46376 5 1 1 46375
0 46377 7 1 2 55155 75866
0 46378 5 1 1 46377
0 46379 7 1 2 73596 46378
0 46380 5 1 1 46379
0 46381 7 1 2 46376 46380
0 46382 5 1 1 46381
0 46383 7 1 2 71019 69934
0 46384 7 1 2 76565 46383
0 46385 5 1 1 46384
0 46386 7 1 2 46382 46385
0 46387 7 1 2 46374 46386
0 46388 5 1 1 46387
0 46389 7 1 2 69946 46388
0 46390 5 1 1 46389
0 46391 7 1 2 55970 75084
0 46392 7 1 2 77361 46391
0 46393 5 1 1 46392
0 46394 7 1 2 46390 46393
0 46395 5 1 1 46394
0 46396 7 1 2 52736 46395
0 46397 5 1 1 46396
0 46398 7 1 2 46368 46397
0 46399 5 1 1 46398
0 46400 7 1 2 53604 46399
0 46401 5 1 1 46400
0 46402 7 1 2 55156 70408
0 46403 5 1 1 46402
0 46404 7 1 2 49826 46403
0 46405 5 1 1 46404
0 46406 7 1 2 76135 79407
0 46407 5 1 1 46406
0 46408 7 1 2 46405 46407
0 46409 5 1 1 46408
0 46410 7 1 2 79726 46409
0 46411 5 1 1 46410
0 46412 7 1 2 46401 46411
0 46413 7 1 2 46353 46412
0 46414 5 1 1 46413
0 46415 7 1 2 51467 46414
0 46416 5 1 1 46415
0 46417 7 1 2 46309 46416
0 46418 5 1 1 46417
0 46419 7 1 2 51670 46418
0 46420 5 1 1 46419
0 46421 7 1 2 50315 79402
0 46422 5 1 1 46421
0 46423 7 1 2 64390 79366
0 46424 5 1 1 46423
0 46425 7 1 2 46422 46424
0 46426 5 1 1 46425
0 46427 7 1 2 49988 46426
0 46428 5 1 1 46427
0 46429 7 1 2 67128 79368
0 46430 5 1 1 46429
0 46431 7 1 2 46428 46430
0 46432 5 1 1 46431
0 46433 7 1 2 52210 46432
0 46434 5 1 1 46433
0 46435 7 2 2 61604 71825
0 46436 5 1 1 79743
0 46437 7 1 2 64391 79744
0 46438 5 1 1 46437
0 46439 7 1 2 52737 75186
0 46440 7 1 2 73452 46439
0 46441 5 1 1 46440
0 46442 7 1 2 59039 73895
0 46443 5 1 1 46442
0 46444 7 1 2 59015 46443
0 46445 7 1 2 46441 46444
0 46446 5 1 1 46445
0 46447 7 1 2 50316 46446
0 46448 5 1 1 46447
0 46449 7 1 2 46438 46448
0 46450 5 1 1 46449
0 46451 7 1 2 49989 46450
0 46452 5 1 1 46451
0 46453 7 1 2 75127 46436
0 46454 5 1 1 46453
0 46455 7 1 2 67129 46454
0 46456 5 1 1 46455
0 46457 7 1 2 46452 46456
0 46458 5 1 1 46457
0 46459 7 1 2 55720 46458
0 46460 5 1 1 46459
0 46461 7 1 2 46434 46460
0 46462 5 1 1 46461
0 46463 7 1 2 53798 46462
0 46464 5 1 1 46463
0 46465 7 1 2 62591 73449
0 46466 5 1 1 46465
0 46467 7 2 2 62993 46466
0 46468 7 2 2 50317 79745
0 46469 7 1 2 50074 79660
0 46470 7 1 2 79747 46469
0 46471 5 1 1 46470
0 46472 7 1 2 46464 46471
0 46473 5 1 1 46472
0 46474 7 1 2 51671 46473
0 46475 5 1 1 46474
0 46476 7 1 2 65830 69188
0 46477 7 1 2 79413 46476
0 46478 5 1 1 46477
0 46479 7 1 2 46475 46478
0 46480 5 1 1 46479
0 46481 7 1 2 51468 46480
0 46482 5 1 1 46481
0 46483 7 1 2 78433 79391
0 46484 5 1 1 46483
0 46485 7 1 2 43406 46484
0 46486 5 1 1 46485
0 46487 7 1 2 73395 46486
0 46488 5 1 1 46487
0 46489 7 1 2 79424 46488
0 46490 5 1 1 46489
0 46491 7 1 2 55430 46490
0 46492 5 1 1 46491
0 46493 7 1 2 43452 46492
0 46494 5 1 1 46493
0 46495 7 1 2 53799 46494
0 46496 5 1 1 46495
0 46497 7 1 2 46482 46496
0 46498 5 1 1 46497
0 46499 7 1 2 52357 46498
0 46500 5 1 1 46499
0 46501 7 1 2 53800 43218
0 46502 5 1 1 46501
0 46503 7 1 2 46500 46502
0 46504 5 1 1 46503
0 46505 7 1 2 50570 46504
0 46506 5 1 1 46505
0 46507 7 1 2 46420 46506
0 46508 7 1 2 46289 46507
0 46509 5 1 1 46508
0 46510 7 1 2 51803 46509
0 46511 5 1 1 46510
0 46512 7 1 2 53801 79347
0 46513 5 1 1 46512
0 46514 7 1 2 73123 72142
0 46515 7 1 2 79748 46514
0 46516 5 1 1 46515
0 46517 7 1 2 46513 46516
0 46518 5 1 1 46517
0 46519 7 1 2 51672 46518
0 46520 5 1 1 46519
0 46521 7 1 2 53802 79343
0 46522 5 1 1 46521
0 46523 7 1 2 46520 46522
0 46524 5 1 1 46523
0 46525 7 1 2 52358 46524
0 46526 5 1 1 46525
0 46527 7 1 2 53803 43036
0 46528 5 1 1 46527
0 46529 7 1 2 46526 46528
0 46530 5 1 1 46529
0 46531 7 1 2 51804 46530
0 46532 5 1 1 46531
0 46533 7 1 2 52846 63677
0 46534 7 3 2 53762 53804
0 46535 7 1 2 71160 79749
0 46536 7 1 2 46533 46535
0 46537 7 1 2 79362 46536
0 46538 5 1 1 46537
0 46539 7 1 2 46532 46538
0 46540 5 1 1 46539
0 46541 7 1 2 58465 46540
0 46542 5 1 1 46541
0 46543 7 1 2 71361 42423
0 46544 5 1 1 46543
0 46545 7 1 2 63793 73396
0 46546 5 1 1 46545
0 46547 7 1 2 46544 46546
0 46548 5 1 1 46547
0 46549 7 1 2 52043 46548
0 46550 5 1 1 46549
0 46551 7 1 2 65160 62430
0 46552 5 1 1 46551
0 46553 7 1 2 79289 46552
0 46554 5 1 1 46553
0 46555 7 1 2 51469 46554
0 46556 5 1 1 46555
0 46557 7 1 2 46550 46556
0 46558 5 1 1 46557
0 46559 7 1 2 51673 46558
0 46560 5 1 1 46559
0 46561 7 1 2 48452 45428
0 46562 5 1 1 46561
0 46563 7 1 2 55590 46562
0 46564 7 2 2 79394 46563
0 46565 7 1 2 79553 79752
0 46566 5 1 1 46565
0 46567 7 1 2 46560 46566
0 46568 5 1 1 46567
0 46569 7 1 2 67869 46568
0 46570 5 1 1 46569
0 46571 7 1 2 52847 79295
0 46572 5 1 1 46571
0 46573 7 1 2 57267 62021
0 46574 5 1 1 46573
0 46575 7 1 2 72923 46574
0 46576 5 1 1 46575
0 46577 7 1 2 65161 46576
0 46578 5 1 1 46577
0 46579 7 1 2 48980 79297
0 46580 5 1 1 46579
0 46581 7 1 2 46578 46580
0 46582 5 1 1 46581
0 46583 7 1 2 79300 46582
0 46584 5 1 1 46583
0 46585 7 1 2 69040 79753
0 46586 5 1 1 46585
0 46587 7 1 2 46584 46586
0 46588 5 1 1 46587
0 46589 7 1 2 51470 46588
0 46590 5 1 1 46589
0 46591 7 1 2 46572 46590
0 46592 7 1 2 46570 46591
0 46593 5 1 1 46592
0 46594 7 1 2 53805 46593
0 46595 5 1 1 46594
0 46596 7 2 2 69915 72143
0 46597 7 2 2 62508 79754
0 46598 7 1 2 58466 60032
0 46599 5 1 1 46598
0 46600 7 2 2 79339 46599
0 46601 5 1 1 79758
0 46602 7 1 2 70698 79759
0 46603 5 1 1 46602
0 46604 7 1 2 79756 46603
0 46605 5 1 1 46604
0 46606 7 1 2 46595 46605
0 46607 5 1 1 46606
0 46608 7 1 2 51805 46607
0 46609 5 1 1 46608
0 46610 7 1 2 53605 79750
0 46611 7 2 2 72295 46610
0 46612 7 1 2 50884 73653
0 46613 7 3 2 79760 46612
0 46614 5 1 1 79762
0 46615 7 1 2 63706 79763
0 46616 5 1 1 46615
0 46617 7 1 2 69434 79317
0 46618 5 2 1 46617
0 46619 7 1 2 53806 79331
0 46620 5 1 1 46619
0 46621 7 4 2 69544 69417
0 46622 7 1 2 62994 79767
0 46623 5 1 1 46622
0 46624 7 1 2 46620 46623
0 46625 5 1 1 46624
0 46626 7 1 2 71161 46625
0 46627 5 1 1 46626
0 46628 7 1 2 79765 46627
0 46629 5 1 1 46628
0 46630 7 1 2 73376 46629
0 46631 5 1 1 46630
0 46632 7 1 2 73493 79751
0 46633 7 1 2 79329 46632
0 46634 5 1 1 46633
0 46635 7 1 2 46631 46634
0 46636 5 1 1 46635
0 46637 7 1 2 51806 57268
0 46638 7 1 2 46636 46637
0 46639 5 1 1 46638
0 46640 7 1 2 46616 46639
0 46641 5 1 1 46640
0 46642 7 1 2 60670 46641
0 46643 5 1 1 46642
0 46644 7 1 2 65162 70384
0 46645 5 2 1 46644
0 46646 7 1 2 48981 59954
0 46647 5 1 1 46646
0 46648 7 1 2 79771 46647
0 46649 5 1 1 46648
0 46650 7 1 2 77961 46649
0 46651 5 1 1 46650
0 46652 7 1 2 79327 79772
0 46653 5 1 1 46652
0 46654 7 1 2 73322 46653
0 46655 5 1 1 46654
0 46656 7 1 2 46651 46655
0 46657 5 1 1 46656
0 46658 7 1 2 51674 46657
0 46659 5 1 1 46658
0 46660 7 1 2 60604 74890
0 46661 5 1 1 46660
0 46662 7 1 2 55157 46661
0 46663 5 1 1 46662
0 46664 7 1 2 55591 46663
0 46665 7 1 2 79227 46664
0 46666 5 1 1 46665
0 46667 7 1 2 46659 46666
0 46668 5 1 1 46667
0 46669 7 1 2 51471 46668
0 46670 5 1 1 46669
0 46671 7 1 2 67794 71162
0 46672 5 1 1 46671
0 46673 7 1 2 66302 71264
0 46674 7 1 2 72950 46673
0 46675 5 1 1 46674
0 46676 7 1 2 46672 46675
0 46677 5 1 1 46676
0 46678 7 1 2 52848 46677
0 46679 5 1 1 46678
0 46680 7 1 2 71163 75071
0 46681 5 1 1 46680
0 46682 7 1 2 46679 46681
0 46683 5 1 1 46682
0 46684 7 1 2 78604 46683
0 46685 5 1 1 46684
0 46686 7 1 2 46670 46685
0 46687 5 1 1 46686
0 46688 7 1 2 53807 51807
0 46689 7 1 2 58467 46688
0 46690 7 1 2 46687 46689
0 46691 5 1 1 46690
0 46692 7 1 2 53808 79314
0 46693 5 1 1 46692
0 46694 7 1 2 73912 72531
0 46695 5 1 1 46694
0 46696 7 1 2 46693 46695
0 46697 5 1 1 46696
0 46698 7 1 2 70011 46697
0 46699 5 1 1 46698
0 46700 7 1 2 69947 79312
0 46701 5 1 1 46700
0 46702 7 1 2 46699 46701
0 46703 5 1 1 46702
0 46704 7 1 2 51808 46703
0 46705 5 1 1 46704
0 46706 7 1 2 46614 46705
0 46707 5 1 1 46706
0 46708 7 1 2 73387 46601
0 46709 7 1 2 46707 46708
0 46710 5 1 1 46709
0 46711 7 1 2 46691 46710
0 46712 7 1 2 46643 46711
0 46713 7 1 2 46609 46712
0 46714 5 1 1 46713
0 46715 7 1 2 53140 46714
0 46716 5 1 1 46715
0 46717 7 1 2 53809 79364
0 46718 5 1 1 46717
0 46719 7 1 2 46716 46718
0 46720 7 1 2 46542 46719
0 46721 5 1 1 46720
0 46722 7 1 2 50571 46721
0 46723 5 1 1 46722
0 46724 7 1 2 53810 79444
0 46725 5 1 1 46724
0 46726 7 1 2 73494 72871
0 46727 7 1 2 79746 46726
0 46728 5 1 1 46727
0 46729 7 1 2 46725 46728
0 46730 5 1 1 46729
0 46731 7 1 2 51809 46730
0 46732 5 1 1 46731
0 46733 7 1 2 53031 71604
0 46734 7 1 2 79764 46733
0 46735 5 1 1 46734
0 46736 7 1 2 46732 46735
0 46737 5 1 1 46736
0 46738 7 1 2 52211 46737
0 46739 5 1 1 46738
0 46740 7 1 2 53811 79442
0 46741 5 1 1 46740
0 46742 7 1 2 46739 46741
0 46743 5 1 1 46742
0 46744 7 1 2 79447 46743
0 46745 5 1 1 46744
0 46746 7 1 2 53812 75184
0 46747 7 1 2 77540 46746
0 46748 7 1 2 72298 46747
0 46749 7 1 2 79452 46748
0 46750 5 1 1 46749
0 46751 7 1 2 46745 46750
0 46752 7 1 2 46723 46751
0 46753 7 1 2 46511 46752
0 46754 5 1 1 46753
0 46755 7 1 2 57070 46754
0 46756 5 1 1 46755
0 46757 7 1 2 53813 79458
0 46758 5 1 1 46757
0 46759 7 1 2 53814 79486
0 46760 5 1 1 46759
0 46761 7 1 2 58548 79757
0 46762 5 1 1 46761
0 46763 7 1 2 46760 46762
0 46764 5 2 1 46763
0 46765 7 1 2 60158 79773
0 46766 5 1 1 46765
0 46767 7 1 2 53815 79496
0 46768 5 1 1 46767
0 46769 7 1 2 62509 70207
0 46770 5 1 1 46769
0 46771 7 1 2 62995 76073
0 46772 7 1 2 61459 46771
0 46773 5 1 1 46772
0 46774 7 1 2 46770 46773
0 46775 5 1 1 46774
0 46776 7 1 2 79755 46775
0 46777 5 1 1 46776
0 46778 7 1 2 46768 46777
0 46779 5 1 1 46778
0 46780 7 1 2 65013 46779
0 46781 5 1 1 46780
0 46782 7 1 2 46766 46781
0 46783 5 1 1 46782
0 46784 7 1 2 51810 46783
0 46785 5 1 1 46784
0 46786 7 1 2 53816 79500
0 46787 5 1 1 46786
0 46788 7 1 2 46785 46787
0 46789 5 1 1 46788
0 46790 7 1 2 58468 46789
0 46791 5 1 1 46790
0 46792 7 1 2 53817 79502
0 46793 5 1 1 46792
0 46794 7 1 2 74411 79318
0 46795 5 1 1 46794
0 46796 7 1 2 52467 79492
0 46797 5 1 1 46796
0 46798 7 1 2 43000 46797
0 46799 5 1 1 46798
0 46800 7 1 2 53818 46799
0 46801 5 1 1 46800
0 46802 7 1 2 62510 79490
0 46803 5 1 1 46802
0 46804 7 1 2 76435 75356
0 46805 5 1 1 46804
0 46806 7 1 2 46803 46805
0 46807 5 1 1 46806
0 46808 7 1 2 72574 72144
0 46809 7 1 2 46807 46808
0 46810 5 1 1 46809
0 46811 7 1 2 46801 46810
0 46812 5 1 1 46811
0 46813 7 1 2 50572 46812
0 46814 5 1 1 46813
0 46815 7 1 2 73913 79319
0 46816 5 1 1 46815
0 46817 7 1 2 52468 79733
0 46818 5 1 1 46817
0 46819 7 1 2 46816 46818
0 46820 5 1 1 46819
0 46821 7 1 2 77909 46820
0 46822 5 1 1 46821
0 46823 7 1 2 73914 79498
0 46824 5 1 1 46823
0 46825 7 1 2 46822 46824
0 46826 7 1 2 46814 46825
0 46827 5 1 1 46826
0 46828 7 1 2 51675 46827
0 46829 5 1 1 46828
0 46830 7 1 2 46795 46829
0 46831 5 1 1 46830
0 46832 7 1 2 57703 46831
0 46833 5 1 1 46832
0 46834 7 1 2 43322 43585
0 46835 5 1 1 46834
0 46836 7 1 2 49990 46835
0 46837 5 1 1 46836
0 46838 7 1 2 65745 79403
0 46839 5 1 1 46838
0 46840 7 1 2 46837 46839
0 46841 5 1 1 46840
0 46842 7 1 2 53819 46841
0 46843 5 1 1 46842
0 46844 7 1 2 69435 68490
0 46845 7 1 2 79494 46844
0 46846 5 1 1 46845
0 46847 7 1 2 46843 46846
0 46848 5 1 1 46847
0 46849 7 1 2 79471 46848
0 46850 5 1 1 46849
0 46851 7 1 2 58549 69189
0 46852 7 1 2 79228 46851
0 46853 5 1 1 46852
0 46854 7 1 2 46850 46853
0 46855 5 1 1 46854
0 46856 7 1 2 51188 46855
0 46857 5 1 1 46856
0 46858 7 1 2 71774 71304
0 46859 5 1 1 46858
0 46860 7 1 2 66969 46859
0 46861 5 1 1 46860
0 46862 7 1 2 73323 46861
0 46863 5 1 1 46862
0 46864 7 1 2 79468 46863
0 46865 5 1 1 46864
0 46866 7 1 2 53820 46865
0 46867 5 1 1 46866
0 46868 7 1 2 79766 46867
0 46869 5 1 1 46868
0 46870 7 1 2 60806 46869
0 46871 5 1 1 46870
0 46872 7 1 2 46857 46871
0 46873 5 1 1 46872
0 46874 7 1 2 51472 46873
0 46875 5 1 1 46874
0 46876 7 1 2 79426 79731
0 46877 7 1 2 79462 46876
0 46878 5 1 1 46877
0 46879 7 1 2 79488 79774
0 46880 5 1 1 46879
0 46881 7 1 2 46878 46880
0 46882 7 1 2 46875 46881
0 46883 7 1 2 46833 46882
0 46884 5 1 1 46883
0 46885 7 1 2 51811 46884
0 46886 5 1 1 46885
0 46887 7 1 2 46793 46886
0 46888 7 1 2 46791 46887
0 46889 5 1 1 46888
0 46890 7 1 2 76383 46889
0 46891 5 1 1 46890
0 46892 7 1 2 46758 46891
0 46893 7 1 2 46756 46892
0 46894 7 1 2 46172 46893
0 46895 5 1 1 46894
0 46896 7 1 2 58066 46895
0 46897 5 1 1 46896
0 46898 7 1 2 53821 79518
0 46899 5 1 1 46898
0 46900 7 2 2 71343 79569
0 46901 5 2 1 79775
0 46902 7 1 2 46899 79777
0 46903 5 1 1 46902
0 46904 7 1 2 51473 46903
0 46905 5 1 1 46904
0 46906 7 1 2 69465 44106
0 46907 5 1 1 46906
0 46908 7 1 2 69466 78872
0 46909 5 1 1 46908
0 46910 7 1 2 79778 46909
0 46911 5 3 1 46910
0 46912 7 1 2 51189 79534
0 46913 7 1 2 79779 46912
0 46914 5 1 1 46913
0 46915 7 1 2 46907 46914
0 46916 7 1 2 46905 46915
0 46917 5 1 1 46916
0 46918 7 1 2 51812 46917
0 46919 5 1 1 46918
0 46920 7 1 2 71539 79740
0 46921 5 1 1 46920
0 46922 7 1 2 12193 72146
0 46923 5 1 1 46922
0 46924 7 1 2 70611 46923
0 46925 5 1 1 46924
0 46926 7 2 2 46921 46925
0 46927 5 1 1 79782
0 46928 7 1 2 49827 79727
0 46929 5 1 1 46928
0 46930 7 1 2 79783 46929
0 46931 5 1 1 46930
0 46932 7 1 2 51813 46931
0 46933 5 1 1 46932
0 46934 7 1 2 72473 79099
0 46935 5 2 1 46934
0 46936 7 1 2 46933 79784
0 46937 5 4 1 46936
0 46938 7 1 2 79520 79786
0 46939 5 1 1 46938
0 46940 7 1 2 51814 46927
0 46941 5 1 1 46940
0 46942 7 1 2 79785 46941
0 46943 5 1 1 46942
0 46944 7 1 2 60228 46943
0 46945 5 1 1 46944
0 46946 7 1 2 46939 46945
0 46947 5 1 1 46946
0 46948 7 1 2 70780 46947
0 46949 5 1 1 46948
0 46950 7 1 2 79504 79787
0 46951 5 1 1 46950
0 46952 7 1 2 46949 46951
0 46953 5 1 1 46952
0 46954 7 1 2 51474 46953
0 46955 5 1 1 46954
0 46956 7 1 2 51815 58903
0 46957 7 1 2 79213 46956
0 46958 7 1 2 70781 46957
0 46959 7 1 2 79780 46958
0 46960 5 1 1 46959
0 46961 7 1 2 46955 46960
0 46962 7 1 2 46919 46961
0 46963 5 1 1 46962
0 46964 7 1 2 51676 46963
0 46965 5 1 1 46964
0 46966 7 1 2 53822 79555
0 46967 5 1 1 46966
0 46968 7 1 2 53823 44444
0 46969 5 1 1 46968
0 46970 7 1 2 53824 79566
0 46971 5 1 1 46970
0 46972 7 1 2 73815 79741
0 46973 7 1 2 70805 46972
0 46974 5 1 1 46973
0 46975 7 1 2 46971 46974
0 46976 5 1 1 46975
0 46977 7 1 2 53606 79561
0 46978 7 1 2 46976 46977
0 46979 5 1 1 46978
0 46980 7 1 2 53825 66109
0 46981 7 1 2 74245 46980
0 46982 5 1 1 46981
0 46983 7 1 2 46979 46982
0 46984 5 1 1 46983
0 46985 7 1 2 58791 46984
0 46986 5 1 1 46985
0 46987 7 2 2 75068 70806
0 46988 7 1 2 72872 79790
0 46989 5 1 1 46988
0 46990 7 3 2 75905 79714
0 46991 5 1 1 79792
0 46992 7 1 2 51190 79557
0 46993 7 1 2 79793 46992
0 46994 5 1 1 46993
0 46995 7 1 2 46989 46994
0 46996 7 1 2 46986 46995
0 46997 7 1 2 46969 46996
0 46998 5 1 1 46997
0 46999 7 1 2 50573 46998
0 47000 5 1 1 46999
0 47001 7 1 2 62511 79537
0 47002 5 1 1 47001
0 47003 7 1 2 72580 47002
0 47004 5 1 1 47003
0 47005 7 1 2 56483 47004
0 47006 5 1 1 47005
0 47007 7 1 2 44359 47006
0 47008 5 1 1 47007
0 47009 7 1 2 79768 47008
0 47010 5 1 1 47009
0 47011 7 2 2 73659 69421
0 47012 7 1 2 57704 79795
0 47013 5 1 1 47012
0 47014 7 1 2 60687 69422
0 47015 7 1 2 79708 47014
0 47016 5 1 1 47015
0 47017 7 1 2 47013 47016
0 47018 5 1 1 47017
0 47019 7 1 2 60881 47018
0 47020 5 1 1 47019
0 47021 7 1 2 60022 79548
0 47022 7 1 2 79794 47021
0 47023 5 1 1 47022
0 47024 7 1 2 47020 47023
0 47025 7 1 2 47010 47024
0 47026 7 1 2 47000 47025
0 47027 7 1 2 46967 47026
0 47028 5 1 1 47027
0 47029 7 1 2 51816 47028
0 47030 5 1 1 47029
0 47031 7 1 2 53826 79571
0 47032 5 1 1 47031
0 47033 7 1 2 50574 79761
0 47034 7 1 2 79791 47033
0 47035 5 1 1 47034
0 47036 7 1 2 47032 47035
0 47037 7 1 2 47030 47036
0 47038 5 1 1 47037
0 47039 7 1 2 57071 47038
0 47040 5 1 1 47039
0 47041 7 1 2 53827 79593
0 47042 5 1 1 47041
0 47043 7 1 2 53828 79613
0 47044 5 1 1 47043
0 47045 7 1 2 72718 76532
0 47046 5 1 1 47045
0 47047 7 1 2 50318 79605
0 47048 7 1 2 79601 47047
0 47049 5 1 1 47048
0 47050 7 1 2 47046 47049
0 47051 5 1 1 47050
0 47052 7 1 2 79715 47051
0 47053 5 1 1 47052
0 47054 7 1 2 47044 47053
0 47055 5 1 1 47054
0 47056 7 1 2 51817 47055
0 47057 5 1 1 47056
0 47058 7 1 2 53829 79617
0 47059 5 1 1 47058
0 47060 7 1 2 79623 79788
0 47061 5 1 1 47060
0 47062 7 1 2 53830 79621
0 47063 5 1 1 47062
0 47064 7 1 2 47061 47063
0 47065 5 1 1 47064
0 47066 7 1 2 51475 47065
0 47067 5 1 1 47066
0 47068 7 1 2 53831 79625
0 47069 5 1 1 47068
0 47070 7 1 2 46991 47069
0 47071 5 1 1 47070
0 47072 7 1 2 79627 47071
0 47073 5 1 1 47072
0 47074 7 1 2 47067 47073
0 47075 5 1 1 47074
0 47076 7 1 2 57705 47075
0 47077 5 1 1 47076
0 47078 7 1 2 47059 47077
0 47079 7 1 2 47057 47078
0 47080 5 1 1 47079
0 47081 7 1 2 61476 47080
0 47082 5 1 1 47081
0 47083 7 1 2 47042 47082
0 47084 7 1 2 47040 47083
0 47085 7 1 2 46965 47084
0 47086 5 1 1 47085
0 47087 7 1 2 50885 47086
0 47088 5 1 1 47087
0 47089 7 1 2 79641 79781
0 47090 5 1 1 47089
0 47091 7 1 2 69467 79629
0 47092 5 1 1 47091
0 47093 7 1 2 47090 47092
0 47094 5 1 1 47093
0 47095 7 1 2 51191 47094
0 47096 5 1 1 47095
0 47097 7 1 2 78986 79639
0 47098 5 1 1 47097
0 47099 7 1 2 49828 78915
0 47100 5 1 1 47099
0 47101 7 1 2 79635 47100
0 47102 5 1 1 47101
0 47103 7 1 2 49645 47102
0 47104 5 1 1 47103
0 47105 7 1 2 79633 47104
0 47106 5 1 1 47105
0 47107 7 1 2 55158 47106
0 47108 5 1 1 47107
0 47109 7 1 2 78393 47108
0 47110 5 1 1 47109
0 47111 7 1 2 69545 47110
0 47112 5 1 1 47111
0 47113 7 1 2 47098 47112
0 47114 5 1 1 47113
0 47115 7 1 2 69468 47114
0 47116 5 1 1 47115
0 47117 7 1 2 47096 47116
0 47118 5 1 1 47117
0 47119 7 1 2 51677 47118
0 47120 5 1 1 47119
0 47121 7 1 2 14346 79695
0 47122 5 1 1 47121
0 47123 7 1 2 59199 47122
0 47124 5 1 1 47123
0 47125 7 1 2 73043 79643
0 47126 5 1 1 47125
0 47127 7 1 2 47124 47126
0 47128 5 1 1 47127
0 47129 7 1 2 79796 47128
0 47130 5 1 1 47129
0 47131 7 1 2 52849 79658
0 47132 5 1 1 47131
0 47133 7 1 2 21833 47132
0 47134 5 1 1 47133
0 47135 7 1 2 72719 47134
0 47136 5 1 1 47135
0 47137 7 1 2 51678 78981
0 47138 5 1 1 47137
0 47139 7 1 2 47136 47138
0 47140 5 1 1 47139
0 47141 7 1 2 78642 47140
0 47142 5 1 1 47141
0 47143 7 1 2 51192 79698
0 47144 7 1 2 79139 47143
0 47145 5 1 1 47144
0 47146 7 1 2 47142 47145
0 47147 5 1 1 47146
0 47148 7 1 2 57706 47147
0 47149 5 1 1 47148
0 47150 7 1 2 62996 79651
0 47151 5 1 1 47150
0 47152 7 1 2 79664 47151
0 47153 5 1 1 47152
0 47154 7 1 2 57707 47153
0 47155 5 1 1 47154
0 47156 7 1 2 62997 79645
0 47157 5 1 1 47156
0 47158 7 1 2 79588 79654
0 47159 5 1 1 47158
0 47160 7 1 2 53607 77627
0 47161 7 1 2 75817 47160
0 47162 7 1 2 78753 47161
0 47163 5 1 1 47162
0 47164 7 1 2 47159 47163
0 47165 7 1 2 47157 47164
0 47166 7 1 2 47155 47165
0 47167 5 1 1 47166
0 47168 7 1 2 73044 47167
0 47169 5 1 1 47168
0 47170 7 1 2 72720 79637
0 47171 5 1 1 47170
0 47172 7 1 2 55159 75906
0 47173 5 1 1 47172
0 47174 7 1 2 47171 47173
0 47175 5 1 1 47174
0 47176 7 1 2 78743 47175
0 47177 5 1 1 47176
0 47178 7 1 2 47169 47177
0 47179 7 1 2 47149 47178
0 47180 5 1 1 47179
0 47181 7 1 2 69469 47180
0 47182 5 1 1 47181
0 47183 7 1 2 47130 47182
0 47184 7 1 2 47120 47183
0 47185 5 1 1 47184
0 47186 7 1 2 51818 47185
0 47187 5 1 1 47186
0 47188 7 1 2 53832 79681
0 47189 5 1 1 47188
0 47190 7 1 2 79595 79683
0 47191 5 1 1 47190
0 47192 7 2 2 59359 79118
0 47193 7 1 2 50319 79797
0 47194 5 1 1 47193
0 47195 7 1 2 47191 47194
0 47196 5 1 1 47195
0 47197 7 1 2 52044 47196
0 47198 5 1 1 47197
0 47199 7 1 2 67814 71521
0 47200 5 1 1 47199
0 47201 7 1 2 47198 47200
0 47202 5 1 1 47201
0 47203 7 1 2 57708 47202
0 47204 5 1 1 47203
0 47205 7 1 2 67536 73740
0 47206 5 1 1 47205
0 47207 7 1 2 79596 79679
0 47208 5 1 1 47207
0 47209 7 1 2 75907 79672
0 47210 5 1 1 47209
0 47211 7 1 2 47208 47210
0 47212 5 1 1 47211
0 47213 7 1 2 51193 47212
0 47214 5 1 1 47213
0 47215 7 1 2 47206 47214
0 47216 7 1 2 47204 47215
0 47217 5 1 1 47216
0 47218 7 1 2 79716 47217
0 47219 5 1 1 47218
0 47220 7 1 2 47189 47219
0 47221 5 1 1 47220
0 47222 7 1 2 51819 47221
0 47223 5 1 1 47222
0 47224 7 1 2 53833 45751
0 47225 5 1 1 47224
0 47226 7 1 2 47223 47225
0 47227 5 1 1 47226
0 47228 7 1 2 70222 47227
0 47229 5 1 1 47228
0 47230 7 1 2 53834 79689
0 47231 5 1 1 47230
0 47232 7 1 2 62746 72575
0 47233 5 1 1 47232
0 47234 7 1 2 52738 73549
0 47235 7 1 2 70452 47234
0 47236 5 1 1 47235
0 47237 7 1 2 47233 47236
0 47238 5 1 1 47237
0 47239 7 1 2 57709 47238
0 47240 5 1 1 47239
0 47241 7 1 2 62512 60825
0 47242 5 1 1 47241
0 47243 7 1 2 55431 47242
0 47244 5 1 1 47243
0 47245 7 1 2 73281 47244
0 47246 5 1 1 47245
0 47247 7 1 2 47240 47246
0 47248 5 1 1 47247
0 47249 7 1 2 50575 47248
0 47250 5 1 1 47249
0 47251 7 1 2 55834 71022
0 47252 5 1 1 47251
0 47253 7 1 2 72576 78289
0 47254 7 1 2 47252 47253
0 47255 5 1 1 47254
0 47256 7 1 2 47250 47255
0 47257 5 1 1 47256
0 47258 7 1 2 56484 47257
0 47259 5 1 1 47258
0 47260 7 1 2 61689 75908
0 47261 5 1 1 47260
0 47262 7 1 2 57710 79597
0 47263 5 1 1 47262
0 47264 7 1 2 47261 47263
0 47265 5 1 1 47264
0 47266 7 1 2 73045 47265
0 47267 5 1 1 47266
0 47268 7 1 2 60443 79696
0 47269 5 1 1 47268
0 47270 7 1 2 67815 71481
0 47271 7 1 2 47269 47270
0 47272 5 1 1 47271
0 47273 7 1 2 47267 47272
0 47274 7 1 2 47259 47273
0 47275 5 1 1 47274
0 47276 7 1 2 79769 47275
0 47277 5 1 1 47276
0 47278 7 1 2 47231 47277
0 47279 5 1 1 47278
0 47280 7 1 2 51820 47279
0 47281 5 1 1 47280
0 47282 7 1 2 53835 79691
0 47283 5 1 1 47282
0 47284 7 1 2 47281 47283
0 47285 5 1 1 47284
0 47286 7 1 2 57072 47285
0 47287 5 1 1 47286
0 47288 7 1 2 53836 79693
0 47289 5 1 1 47288
0 47290 7 1 2 69019 75178
0 47291 7 1 2 79710 47290
0 47292 5 1 1 47291
0 47293 7 1 2 79706 47292
0 47294 5 1 1 47293
0 47295 7 1 2 53837 47294
0 47296 5 1 1 47295
0 47297 7 2 2 69546 73915
0 47298 7 1 2 79589 79799
0 47299 5 1 1 47298
0 47300 7 1 2 46292 47299
0 47301 5 1 1 47300
0 47302 7 1 2 72721 47301
0 47303 5 1 1 47302
0 47304 7 1 2 78971 79702
0 47305 5 1 1 47304
0 47306 7 1 2 52850 79704
0 47307 5 1 1 47306
0 47308 7 1 2 47305 47307
0 47309 5 1 1 47308
0 47310 7 1 2 53838 47309
0 47311 5 1 1 47310
0 47312 7 1 2 47303 47311
0 47313 5 1 1 47312
0 47314 7 1 2 73046 47313
0 47315 5 1 1 47314
0 47316 7 1 2 53839 45958
0 47317 5 1 1 47316
0 47318 7 1 2 78643 78954
0 47319 5 1 1 47318
0 47320 7 1 2 75912 47319
0 47321 5 1 1 47320
0 47322 7 1 2 79800 47321
0 47323 5 1 1 47322
0 47324 7 1 2 47317 47323
0 47325 7 1 2 47315 47324
0 47326 5 1 1 47325
0 47327 7 1 2 51821 47326
0 47328 5 1 1 47327
0 47329 7 1 2 47296 47328
0 47330 5 1 1 47329
0 47331 7 1 2 51679 47330
0 47332 5 1 1 47331
0 47333 7 1 2 47289 47332
0 47334 5 1 1 47333
0 47335 7 1 2 66672 47334
0 47336 5 1 1 47335
0 47337 7 1 2 49081 47336
0 47338 7 1 2 47287 47337
0 47339 7 1 2 47229 47338
0 47340 7 1 2 47187 47339
0 47341 7 1 2 47088 47340
0 47342 7 1 2 46897 47341
0 47343 7 1 2 53840 79091
0 47344 5 1 1 47343
0 47345 7 1 2 55971 73236
0 47346 5 1 1 47345
0 47347 7 1 2 66207 47346
0 47348 5 1 1 47347
0 47349 7 1 2 71497 47348
0 47350 5 1 1 47349
0 47351 7 1 2 67413 79052
0 47352 5 1 1 47351
0 47353 7 1 2 47350 47352
0 47354 5 1 1 47353
0 47355 7 1 2 50576 47354
0 47356 5 1 1 47355
0 47357 7 1 2 51476 73196
0 47358 5 1 1 47357
0 47359 7 1 2 71237 78996
0 47360 5 1 1 47359
0 47361 7 1 2 40728 47360
0 47362 5 1 1 47361
0 47363 7 1 2 51194 47362
0 47364 5 1 1 47363
0 47365 7 1 2 47358 47364
0 47366 7 1 2 47356 47365
0 47367 5 1 1 47366
0 47368 7 1 2 75909 47367
0 47369 5 1 1 47368
0 47370 7 1 2 79109 79598
0 47371 5 1 1 47370
0 47372 7 1 2 47369 47371
0 47373 5 1 1 47372
0 47374 7 1 2 79717 47373
0 47375 5 1 1 47374
0 47376 7 1 2 47344 47375
0 47377 5 1 1 47376
0 47378 7 1 2 51822 47377
0 47379 5 1 1 47378
0 47380 7 1 2 53841 79148
0 47381 5 1 1 47380
0 47382 7 1 2 79153 79599
0 47383 5 1 1 47382
0 47384 7 1 2 52469 77783
0 47385 5 1 1 47384
0 47386 7 1 2 50886 77905
0 47387 5 1 1 47386
0 47388 7 1 2 47385 47387
0 47389 5 1 1 47388
0 47390 7 1 2 59360 70612
0 47391 7 1 2 47389 47390
0 47392 5 1 1 47391
0 47393 7 1 2 47383 47392
0 47394 5 1 1 47393
0 47395 7 1 2 79718 47394
0 47396 5 1 1 47395
0 47397 7 1 2 47381 47396
0 47398 5 1 1 47397
0 47399 7 1 2 51823 47398
0 47400 5 1 1 47399
0 47401 7 4 2 53842 79100
0 47402 7 1 2 79155 79801
0 47403 5 1 1 47402
0 47404 7 1 2 47400 47403
0 47405 5 1 1 47404
0 47406 7 1 2 57269 47405
0 47407 5 1 1 47406
0 47408 7 1 2 53843 79163
0 47409 5 1 1 47408
0 47410 7 1 2 71540 73850
0 47411 5 1 1 47410
0 47412 7 1 2 61252 73331
0 47413 5 1 1 47412
0 47414 7 1 2 75073 47413
0 47415 5 1 1 47414
0 47416 7 1 2 71522 47415
0 47417 5 1 1 47416
0 47418 7 1 2 47411 47417
0 47419 5 1 1 47418
0 47420 7 1 2 79770 47419
0 47421 5 1 1 47420
0 47422 7 1 2 47409 47421
0 47423 5 1 1 47422
0 47424 7 1 2 51824 47423
0 47425 5 1 1 47424
0 47426 7 1 2 79165 79802
0 47427 5 1 1 47426
0 47428 7 1 2 47425 47427
0 47429 5 1 1 47428
0 47430 7 1 2 57073 47429
0 47431 5 1 1 47430
0 47432 7 1 2 53844 79188
0 47433 5 1 1 47432
0 47434 7 1 2 53845 79177
0 47435 5 1 1 47434
0 47436 7 1 2 72722 79173
0 47437 5 1 1 47436
0 47438 7 1 2 73744 47437
0 47439 5 1 1 47438
0 47440 7 1 2 51477 47439
0 47441 5 1 1 47440
0 47442 7 1 2 73004 79798
0 47443 5 1 1 47442
0 47444 7 1 2 47441 47443
0 47445 5 1 1 47444
0 47446 7 1 2 75085 47445
0 47447 5 1 1 47446
0 47448 7 1 2 47435 47447
0 47449 5 1 1 47448
0 47450 7 1 2 51825 47449
0 47451 5 1 1 47450
0 47452 7 1 2 79179 79803
0 47453 5 1 1 47452
0 47454 7 1 2 47451 47453
0 47455 5 1 1 47454
0 47456 7 1 2 51680 47455
0 47457 5 1 1 47456
0 47458 7 1 2 47433 47457
0 47459 7 1 2 47431 47458
0 47460 7 1 2 47407 47459
0 47461 5 1 1 47460
0 47462 7 1 2 57711 47461
0 47463 5 1 1 47462
0 47464 7 1 2 79111 79804
0 47465 5 1 1 47464
0 47466 7 1 2 47463 47465
0 47467 7 1 2 47379 47466
0 47468 5 1 1 47467
0 47469 7 1 2 58469 47468
0 47470 5 1 1 47469
0 47471 7 1 2 78917 79789
0 47472 5 1 1 47471
0 47473 7 1 2 52851 68351
0 47474 5 2 1 47473
0 47475 7 1 2 48982 54116
0 47476 5 2 1 47475
0 47477 7 1 2 63896 71873
0 47478 5 1 1 47477
0 47479 7 1 2 79807 47478
0 47480 5 1 1 47479
0 47481 7 1 2 53763 47480
0 47482 5 1 1 47481
0 47483 7 1 2 79805 47482
0 47484 5 1 1 47483
0 47485 7 1 2 56599 47484
0 47486 5 1 1 47485
0 47487 7 1 2 64967 78836
0 47488 5 1 1 47487
0 47489 7 1 2 78874 47488
0 47490 5 1 1 47489
0 47491 7 1 2 47486 47490
0 47492 5 1 1 47491
0 47493 7 1 2 55835 47492
0 47494 5 1 1 47493
0 47495 7 1 2 60003 78881
0 47496 5 1 1 47495
0 47497 7 1 2 63317 70617
0 47498 5 1 1 47497
0 47499 7 1 2 67850 47498
0 47500 5 1 1 47499
0 47501 7 1 2 66747 47500
0 47502 5 1 1 47501
0 47503 7 1 2 47496 47502
0 47504 5 1 1 47503
0 47505 7 1 2 74802 47504
0 47506 5 1 1 47505
0 47507 7 1 2 77096 78875
0 47508 5 1 1 47507
0 47509 7 1 2 61951 68182
0 47510 5 1 1 47509
0 47511 7 1 2 69547 47510
0 47512 5 1 1 47511
0 47513 7 1 2 76514 47512
0 47514 5 1 1 47513
0 47515 7 1 2 72807 71859
0 47516 5 1 1 47515
0 47517 7 1 2 69548 47516
0 47518 5 1 1 47517
0 47519 7 1 2 29785 47518
0 47520 5 1 1 47519
0 47521 7 1 2 47514 47520
0 47522 5 1 1 47521
0 47523 7 1 2 69656 47522
0 47524 5 1 1 47523
0 47525 7 1 2 47508 47524
0 47526 7 1 2 47506 47525
0 47527 5 1 1 47526
0 47528 7 1 2 54417 47527
0 47529 5 1 1 47528
0 47530 7 1 2 59237 78876
0 47531 5 1 1 47530
0 47532 7 2 2 48835 58232
0 47533 7 1 2 59045 67479
0 47534 7 1 2 79809 47533
0 47535 5 1 1 47534
0 47536 7 1 2 47531 47535
0 47537 5 1 1 47536
0 47538 7 1 2 58413 61917
0 47539 7 1 2 47537 47538
0 47540 5 1 1 47539
0 47541 7 1 2 47529 47540
0 47542 7 1 2 47494 47541
0 47543 5 1 1 47542
0 47544 7 1 2 56781 47543
0 47545 5 1 1 47544
0 47546 7 1 2 59049 78844
0 47547 5 1 1 47546
0 47548 7 1 2 59238 78840
0 47549 5 1 1 47548
0 47550 7 1 2 57191 78197
0 47551 5 1 1 47550
0 47552 7 1 2 55836 77762
0 47553 5 1 1 47552
0 47554 7 1 2 47551 47553
0 47555 7 1 2 47549 47554
0 47556 5 1 1 47555
0 47557 7 1 2 57968 47556
0 47558 5 1 1 47557
0 47559 7 1 2 47547 47558
0 47560 5 1 1 47559
0 47561 7 1 2 54809 47560
0 47562 5 1 1 47561
0 47563 7 1 2 61323 78838
0 47564 5 1 1 47563
0 47565 7 1 2 47562 47564
0 47566 5 1 1 47565
0 47567 7 1 2 77950 47566
0 47568 5 1 1 47567
0 47569 7 1 2 73324 40009
0 47570 5 1 1 47569
0 47571 7 1 2 54810 59241
0 47572 5 1 1 47571
0 47573 7 1 2 66673 47572
0 47574 5 1 1 47573
0 47575 7 1 2 78877 47574
0 47576 5 1 1 47575
0 47577 7 1 2 56169 67870
0 47578 5 1 1 47577
0 47579 7 1 2 58494 66821
0 47580 7 1 2 63362 47579
0 47581 5 1 1 47580
0 47582 7 1 2 47578 47581
0 47583 5 1 1 47582
0 47584 7 1 2 56600 47583
0 47585 5 1 1 47584
0 47586 7 1 2 47576 47585
0 47587 5 1 1 47586
0 47588 7 1 2 60257 47587
0 47589 5 1 1 47588
0 47590 7 1 2 48022 3123
0 47591 5 1 1 47590
0 47592 7 1 2 78848 47591
0 47593 5 1 1 47592
0 47594 7 1 2 78878 47593
0 47595 5 1 1 47594
0 47596 7 1 2 78815 79810
0 47597 5 1 1 47596
0 47598 7 1 2 79808 47597
0 47599 5 1 1 47598
0 47600 7 1 2 53764 47599
0 47601 5 1 1 47600
0 47602 7 1 2 79806 47601
0 47603 5 1 1 47602
0 47604 7 1 2 65605 47603
0 47605 5 1 1 47604
0 47606 7 1 2 47595 47605
0 47607 5 1 1 47606
0 47608 7 1 2 61984 47607
0 47609 5 1 1 47608
0 47610 7 1 2 58950 78879
0 47611 5 1 1 47610
0 47612 7 1 2 78883 47611
0 47613 5 1 1 47612
0 47614 7 1 2 78850 47613
0 47615 5 1 1 47614
0 47616 7 1 2 47609 47615
0 47617 7 1 2 47589 47616
0 47618 7 1 2 47570 47617
0 47619 7 1 2 47568 47618
0 47620 7 1 2 47545 47619
0 47621 5 1 1 47620
0 47622 7 1 2 53846 47621
0 47623 5 1 1 47622
0 47624 7 1 2 70613 79742
0 47625 5 1 1 47624
0 47626 7 1 2 47623 47625
0 47627 5 1 1 47626
0 47628 7 1 2 53608 47627
0 47629 5 1 1 47628
0 47630 7 1 2 70332 79728
0 47631 5 1 1 47630
0 47632 7 1 2 47629 47631
0 47633 5 1 1 47632
0 47634 7 1 2 51826 47633
0 47635 5 1 1 47634
0 47636 7 1 2 47472 47635
0 47637 5 1 1 47636
0 47638 7 1 2 51195 47637
0 47639 5 1 1 47638
0 47640 7 1 2 53847 40471
0 47641 5 1 1 47640
0 47642 7 1 2 71552 78924
0 47643 5 1 1 47642
0 47644 7 1 2 79776 47643
0 47645 5 1 1 47644
0 47646 7 1 2 47641 47645
0 47647 5 1 1 47646
0 47648 7 1 2 51827 47647
0 47649 5 1 1 47648
0 47650 7 1 2 47639 47649
0 47651 5 1 1 47650
0 47652 7 1 2 51681 47651
0 47653 5 1 1 47652
0 47654 7 1 2 53848 78956
0 47655 5 1 1 47654
0 47656 7 1 2 72355 75997
0 47657 7 1 2 79192 47656
0 47658 5 1 1 47657
0 47659 7 1 2 79466 47658
0 47660 5 1 1 47659
0 47661 7 1 2 52739 47660
0 47662 5 1 1 47661
0 47663 7 1 2 70535 75172
0 47664 7 1 2 79392 47663
0 47665 5 1 1 47664
0 47666 7 1 2 47662 47665
0 47667 5 1 1 47666
0 47668 7 1 2 52359 47667
0 47669 5 1 1 47668
0 47670 7 1 2 60432 61441
0 47671 7 1 2 78744 47670
0 47672 5 1 1 47671
0 47673 7 1 2 47669 47672
0 47674 5 1 1 47673
0 47675 7 1 2 53849 47674
0 47676 5 1 1 47675
0 47677 7 1 2 60778 71265
0 47678 7 1 2 74393 79427
0 47679 7 1 2 47677 47678
0 47680 5 1 1 47679
0 47681 7 2 2 53850 63918
0 47682 7 1 2 55592 78829
0 47683 7 1 2 79811 47682
0 47684 5 1 1 47683
0 47685 7 1 2 47680 47684
0 47686 5 1 1 47685
0 47687 7 1 2 52852 47686
0 47688 5 1 1 47687
0 47689 7 1 2 67964 78060
0 47690 5 1 1 47689
0 47691 7 1 2 70479 70546
0 47692 7 1 2 79473 47691
0 47693 5 1 1 47692
0 47694 7 1 2 47690 47693
0 47695 5 1 1 47694
0 47696 7 1 2 79812 47695
0 47697 5 1 1 47696
0 47698 7 1 2 47688 47697
0 47699 5 1 1 47698
0 47700 7 1 2 56485 47699
0 47701 5 1 1 47700
0 47702 7 1 2 52740 58897
0 47703 7 1 2 73667 47702
0 47704 7 1 2 70453 79719
0 47705 7 1 2 47703 47704
0 47706 5 1 1 47705
0 47707 7 1 2 47701 47706
0 47708 7 1 2 47676 47707
0 47709 5 1 1 47708
0 47710 7 1 2 51828 47709
0 47711 5 1 1 47710
0 47712 7 1 2 52911 73495
0 47713 7 1 2 79738 47712
0 47714 7 1 2 60797 72818
0 47715 7 1 2 75306 47714
0 47716 7 1 2 47713 47715
0 47717 5 1 1 47716
0 47718 7 1 2 47711 47717
0 47719 5 1 1 47718
0 47720 7 1 2 70782 47719
0 47721 5 1 1 47720
0 47722 7 1 2 47655 47721
0 47723 7 1 2 47653 47722
0 47724 5 1 1 47723
0 47725 7 1 2 51478 47724
0 47726 5 1 1 47725
0 47727 7 1 2 47470 47726
0 47728 7 1 2 47342 47727
0 47729 5 1 1 47728
0 47730 7 1 2 51 47729
0 47731 7 1 2 46015 47730
0 47732 5 1 1 47731
0 47733 7 1 2 22454 47732
3 129999 5 0 1 47733
