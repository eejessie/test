1 0 0 2 0
2 7 1 0
2 67 1 0
1 1 0 2 0
2 68 1 1
2 69 1 1
1 2 0 2 0
2 70 1 2
2 71 1 2
1 3 0 2 0
2 72 1 3
2 73 1 3
1 4 0 2 0
2 74 1 4
2 75 1 4
1 5 0 2 0
2 76 1 5
2 77 1 5
1 6 0 2 0
2 78 1 6
2 79 1 6
2 80 1 15
2 81 1 15
2 82 1 16
2 83 1 16
2 84 1 18
2 85 1 18
2 86 1 21
2 87 1 21
2 88 1 24
2 89 1 24
2 90 1 27
2 91 1 27
2 92 1 29
2 93 1 29
2 94 1 30
2 95 1 30
2 96 1 31
2 97 1 31
2 98 1 34
2 99 1 34
2 100 1 37
2 101 1 37
2 102 1 38
2 103 1 38
2 104 1 45
2 105 1 45
2 106 1 51
2 107 1 51
2 108 1 52
2 109 1 52
0 8 5 1 1 7
0 9 5 1 1 68
0 10 5 1 1 70
0 11 5 1 1 72
0 12 5 1 1 74
0 13 5 1 1 76
0 14 5 1 1 78
0 15 7 2 2 67 71
0 16 5 2 1 80
0 17 7 1 2 69 73
0 18 5 2 1 17
0 19 7 1 2 9 11
0 20 5 1 1 19
0 21 7 2 2 84 20
0 22 5 1 1 86
0 23 7 1 2 81 87
0 24 5 2 1 23
0 25 7 1 2 82 22
0 26 5 1 1 25
0 27 7 2 2 88 26
0 28 5 1 1 90
0 29 7 2 2 77 28
0 30 5 2 1 92
0 31 7 2 2 85 89
0 32 5 1 1 96
0 33 7 1 2 14 32
0 34 5 2 1 33
0 35 7 1 2 79 97
0 36 5 1 1 35
0 37 7 2 2 98 36
0 38 5 2 1 100
0 39 7 1 2 94 102
0 40 5 1 1 39
0 41 7 1 2 93 99
0 42 5 1 1 41
0 43 7 1 2 8 10
0 44 5 1 1 43
0 45 7 2 2 83 44
0 46 5 1 1 104
0 47 7 1 2 75 46
0 48 7 1 2 42 47
0 49 7 1 2 40 48
0 50 5 1 1 49
0 51 7 2 2 13 91
0 52 5 2 1 106
0 53 7 1 2 101 107
0 54 5 1 1 53
0 55 7 1 2 95 108
0 56 5 1 1 55
0 57 7 1 2 12 105
0 58 5 1 1 57
0 59 7 1 2 56 58
0 60 5 1 1 59
0 61 7 1 2 103 109
0 62 5 1 1 61
0 63 7 1 2 60 62
0 64 7 1 2 54 63
0 65 5 1 1 64
0 66 7 1 2 50 65
3 139 5 0 1 66
