1 0 0 2 0
2 49 1 0
2 739 1 0
1 1 0 2 0
2 740 1 1
2 741 1 1
1 2 0 2 0
2 742 1 2
2 743 1 2
1 3 0 2 0
2 744 1 3
2 745 1 3
1 4 0 2 0
2 746 1 4
2 747 1 4
1 5 0 2 0
2 748 1 5
2 749 1 5
1 6 0 2 0
2 750 1 6
2 751 1 6
1 7 0 2 0
2 752 1 7
2 753 1 7
1 8 0 2 0
2 754 1 8
2 755 1 8
1 9 0 2 0
2 756 1 9
2 757 1 9
1 10 0 2 0
2 758 1 10
2 759 1 10
1 11 0 2 0
2 760 1 11
2 761 1 11
1 12 0 2 0
2 762 1 12
2 763 1 12
1 13 0 2 0
2 764 1 13
2 765 1 13
1 14 0 2 0
2 766 1 14
2 767 1 14
1 15 0 2 0
2 768 1 15
2 769 1 15
1 16 0 2 0
2 770 1 16
2 771 1 16
1 17 0 2 0
2 772 1 17
2 773 1 17
1 18 0 2 0
2 774 1 18
2 775 1 18
1 19 0 2 0
2 776 1 19
2 777 1 19
1 20 0 2 0
2 778 1 20
2 779 1 20
1 21 0 2 0
2 780 1 21
2 781 1 21
1 22 0 2 0
2 782 1 22
2 783 1 22
1 23 0 2 0
2 784 1 23
2 785 1 23
1 24 0 2 0
2 786 1 24
2 787 1 24
1 25 0 2 0
2 788 1 25
2 789 1 25
1 26 0 2 0
2 790 1 26
2 791 1 26
1 27 0 2 0
2 792 1 27
2 793 1 27
1 28 0 2 0
2 794 1 28
2 795 1 28
1 29 0 2 0
2 796 1 29
2 797 1 29
1 30 0 2 0
2 798 1 30
2 799 1 30
1 31 0 2 0
2 800 1 31
2 801 1 31
1 32 0 2 0
2 802 1 32
2 803 1 32
1 33 0 3 0
2 804 1 33
2 805 1 33
2 806 1 33
1 34 0 2 0
2 807 1 34
2 808 1 34
1 35 0 2 0
2 809 1 35
2 810 1 35
1 36 0 2 0
2 811 1 36
2 812 1 36
1 37 0 2 0
2 813 1 37
2 814 1 37
1 38 0 2 0
2 815 1 38
2 816 1 38
1 39 0 2 0
2 817 1 39
2 818 1 39
1 40 0 2 0
2 819 1 40
2 820 1 40
1 41 0 2 0
2 821 1 41
2 822 1 41
1 42 0 2 0
2 823 1 42
2 824 1 42
1 43 0 2 0
2 825 1 43
2 826 1 43
1 44 0 2 0
2 827 1 44
2 828 1 44
1 45 0 2 0
2 829 1 45
2 830 1 45
1 46 0 2 0
2 831 1 46
2 832 1 46
1 47 0 2 0
2 833 1 47
2 834 1 47
1 48 0 2 0
2 835 1 48
2 836 1 48
2 837 1 69
2 838 1 69
2 839 1 70
2 840 1 70
2 841 1 71
2 842 1 71
2 843 1 72
2 844 1 72
2 845 1 73
2 846 1 73
2 847 1 74
2 848 1 74
2 849 1 75
2 850 1 75
2 851 1 76
2 852 1 76
2 853 1 77
2 854 1 77
2 855 1 78
2 856 1 78
2 857 1 79
2 858 1 79
2 859 1 80
2 860 1 80
2 861 1 100
2 862 1 100
2 863 1 102
2 864 1 102
2 865 1 104
2 866 1 104
2 867 1 106
2 868 1 106
2 869 1 108
2 870 1 108
2 871 1 110
2 872 1 110
2 873 1 111
2 874 1 111
2 875 1 112
2 876 1 112
2 877 1 112
2 878 1 115
2 879 1 115
2 880 1 116
2 881 1 116
2 882 1 119
2 883 1 119
2 884 1 122
2 885 1 122
2 886 1 124
2 887 1 124
2 888 1 127
2 889 1 127
2 890 1 130
2 891 1 130
2 892 1 132
2 893 1 132
2 894 1 135
2 895 1 135
2 896 1 138
2 897 1 138
2 898 1 140
2 899 1 140
2 900 1 143
2 901 1 143
2 902 1 146
2 903 1 146
2 904 1 148
2 905 1 148
2 906 1 151
2 907 1 151
2 908 1 154
2 909 1 154
2 910 1 156
2 911 1 156
2 912 1 159
2 913 1 159
2 914 1 162
2 915 1 162
2 916 1 164
2 917 1 164
2 918 1 167
2 919 1 167
2 920 1 170
2 921 1 170
2 922 1 172
2 923 1 172
2 924 1 175
2 925 1 175
2 926 1 178
2 927 1 178
2 928 1 180
2 929 1 180
2 930 1 183
2 931 1 183
2 932 1 186
2 933 1 186
2 934 1 188
2 935 1 188
2 936 1 191
2 937 1 191
2 938 1 194
2 939 1 194
2 940 1 196
2 941 1 196
2 942 1 199
2 943 1 199
2 944 1 202
2 945 1 202
2 946 1 204
2 947 1 204
2 948 1 207
2 949 1 207
2 950 1 210
2 951 1 210
2 952 1 212
2 953 1 212
2 954 1 215
2 955 1 215
2 956 1 216
2 957 1 216
2 958 1 219
2 959 1 219
2 960 1 221
2 961 1 221
2 962 1 222
2 963 1 222
2 964 1 222
2 965 1 223
2 966 1 223
2 967 1 224
2 968 1 224
2 969 1 225
2 970 1 225
2 971 1 231
2 972 1 231
2 973 1 234
2 974 1 234
2 975 1 234
2 976 1 234
2 977 1 236
2 978 1 236
2 979 1 236
2 980 1 237
2 981 1 237
2 982 1 243
2 983 1 243
2 984 1 246
2 985 1 246
2 986 1 246
2 987 1 246
2 988 1 248
2 989 1 248
2 990 1 248
2 991 1 249
2 992 1 249
2 993 1 255
2 994 1 255
2 995 1 258
2 996 1 258
2 997 1 258
2 998 1 258
2 999 1 260
2 1000 1 260
2 1001 1 260
2 1002 1 261
2 1003 1 261
2 1004 1 267
2 1005 1 267
2 1006 1 270
2 1007 1 270
2 1008 1 270
2 1009 1 270
2 1010 1 272
2 1011 1 272
2 1012 1 272
2 1013 1 273
2 1014 1 273
2 1015 1 279
2 1016 1 279
2 1017 1 282
2 1018 1 282
2 1019 1 282
2 1020 1 282
2 1021 1 284
2 1022 1 284
2 1023 1 284
2 1024 1 285
2 1025 1 285
2 1026 1 291
2 1027 1 291
2 1028 1 294
2 1029 1 294
2 1030 1 294
2 1031 1 296
2 1032 1 296
2 1033 1 296
2 1034 1 296
2 1035 1 297
2 1036 1 297
2 1037 1 303
2 1038 1 303
2 1039 1 306
2 1040 1 306
2 1041 1 306
2 1042 1 306
2 1043 1 307
2 1044 1 307
2 1045 1 313
2 1046 1 313
2 1047 1 316
2 1048 1 316
2 1049 1 316
2 1050 1 317
2 1051 1 317
2 1052 1 323
2 1053 1 323
2 1054 1 326
2 1055 1 326
2 1056 1 326
2 1057 1 326
2 1058 1 328
2 1059 1 328
2 1060 1 328
2 1061 1 329
2 1062 1 329
2 1063 1 335
2 1064 1 335
2 1065 1 337
2 1066 1 337
2 1067 1 338
2 1068 1 338
2 1069 1 338
2 1070 1 338
2 1071 1 339
2 1072 1 339
2 1073 1 345
2 1074 1 345
2 1075 1 348
2 1076 1 348
2 1077 1 348
2 1078 1 350
2 1079 1 350
2 1080 1 350
2 1081 1 351
2 1082 1 351
2 1083 1 357
2 1084 1 357
2 1085 1 360
2 1086 1 360
2 1087 1 360
2 1088 1 360
2 1089 1 362
2 1090 1 362
2 1091 1 362
2 1092 1 362
2 1093 1 363
2 1094 1 363
2 1095 1 369
2 1096 1 369
2 1097 1 372
2 1098 1 372
2 1099 1 372
2 1100 1 374
2 1101 1 374
2 1102 1 374
2 1103 1 375
2 1104 1 375
2 1105 1 381
2 1106 1 381
2 1107 1 384
2 1108 1 384
2 1109 1 384
2 1110 1 386
2 1111 1 386
2 1112 1 386
2 1113 1 387
2 1114 1 387
2 1115 1 388
2 1116 1 388
2 1117 1 393
2 1118 1 393
2 1119 1 398
2 1120 1 398
2 1121 1 401
2 1122 1 401
2 1123 1 406
2 1124 1 406
2 1125 1 406
2 1126 1 410
2 1127 1 410
2 1128 1 411
2 1129 1 411
2 1130 1 414
2 1131 1 414
2 1132 1 416
2 1133 1 416
2 1134 1 418
2 1135 1 418
2 1136 1 419
2 1137 1 419
2 1138 1 422
2 1139 1 422
2 1140 1 425
2 1141 1 425
2 1142 1 426
2 1143 1 426
2 1144 1 426
2 1145 1 428
2 1146 1 428
2 1147 1 430
2 1148 1 430
2 1149 1 431
2 1150 1 431
2 1151 1 433
2 1152 1 433
2 1153 1 433
2 1154 1 436
2 1155 1 436
2 1156 1 439
2 1157 1 439
2 1158 1 439
2 1159 1 441
2 1160 1 441
2 1161 1 447
2 1162 1 447
2 1163 1 454
2 1164 1 454
2 1165 1 456
2 1166 1 456
2 1167 1 460
2 1168 1 460
2 1169 1 464
2 1170 1 464
2 1171 1 468
2 1172 1 468
2 1173 1 472
2 1174 1 472
2 1175 1 473
2 1176 1 473
2 1177 1 478
2 1178 1 478
2 1179 1 479
2 1180 1 479
2 1181 1 482
2 1182 1 482
2 1183 1 483
2 1184 1 483
2 1185 1 488
2 1186 1 488
2 1187 1 488
2 1188 1 494
2 1189 1 494
2 1190 1 495
2 1191 1 495
2 1192 1 498
2 1193 1 498
2 1194 1 498
2 1195 1 504
2 1196 1 504
2 1197 1 505
2 1198 1 505
2 1199 1 508
2 1200 1 508
2 1201 1 508
2 1202 1 509
2 1203 1 509
2 1204 1 512
2 1205 1 512
2 1206 1 513
2 1207 1 513
2 1208 1 518
2 1209 1 518
2 1210 1 518
2 1211 1 519
2 1212 1 519
2 1213 1 525
2 1214 1 525
2 1215 1 528
2 1216 1 528
2 1217 1 528
2 1218 1 529
2 1219 1 529
2 1220 1 534
2 1221 1 534
2 1222 1 534
2 1223 1 535
2 1224 1 535
2 1225 1 583
2 1226 1 583
2 1227 1 584
2 1228 1 584
2 1229 1 587
2 1230 1 587
2 1231 1 587
2 1232 1 591
2 1233 1 591
2 1234 1 593
2 1235 1 593
2 1236 1 595
2 1237 1 595
2 1238 1 595
2 1239 1 599
2 1240 1 599
2 1241 1 600
2 1242 1 600
2 1243 1 603
2 1244 1 603
2 1245 1 607
2 1246 1 607
2 1247 1 608
2 1248 1 608
2 1249 1 611
2 1250 1 611
2 1251 1 612
2 1252 1 612
2 1253 1 615
2 1254 1 615
2 1255 1 616
2 1256 1 616
2 1257 1 619
2 1258 1 619
2 1259 1 620
2 1260 1 620
2 1261 1 623
2 1262 1 623
2 1263 1 624
2 1264 1 624
2 1265 1 627
2 1266 1 627
2 1267 1 628
2 1268 1 628
2 1269 1 631
2 1270 1 631
2 1271 1 632
2 1272 1 632
2 1273 1 636
2 1274 1 636
0 50 5 1 1 49
0 51 5 1 1 740
0 52 5 1 1 742
0 53 5 1 1 744
0 54 5 1 1 746
0 55 5 1 1 748
0 56 5 1 1 750
0 57 5 1 1 752
0 58 5 1 1 754
0 59 5 1 1 756
0 60 5 1 1 758
0 61 5 1 1 760
0 62 5 1 1 762
0 63 5 1 1 764
0 64 5 1 1 766
0 65 5 1 1 768
0 66 5 1 1 770
0 67 5 1 1 772
0 68 5 1 1 774
0 69 5 2 1 776
0 70 5 2 1 778
0 71 5 2 1 780
0 72 5 2 1 782
0 73 5 2 1 784
0 74 5 2 1 786
0 75 5 2 1 788
0 76 5 2 1 790
0 77 5 2 1 792
0 78 5 2 1 794
0 79 5 2 1 796
0 80 5 2 1 798
0 81 5 1 1 800
0 82 5 1 1 802
0 83 5 1 1 804
0 84 5 1 1 807
0 85 5 1 1 809
0 86 5 1 1 811
0 87 5 1 1 813
0 88 5 1 1 815
0 89 5 1 1 817
0 90 5 1 1 819
0 91 5 1 1 821
0 92 5 1 1 823
0 93 5 1 1 825
0 94 5 1 1 827
0 95 5 1 1 829
0 96 5 1 1 831
0 97 5 1 1 833
0 98 5 1 1 835
0 99 7 1 2 65 81
0 100 5 2 1 99
0 101 7 1 2 769 801
0 102 5 2 1 101
0 103 7 1 2 52 68
0 104 5 2 1 103
0 105 7 1 2 743 775
0 106 5 2 1 105
0 107 7 1 2 51 67
0 108 5 2 1 107
0 109 7 1 2 741 773
0 110 5 2 1 109
0 111 7 2 2 739 771
0 112 5 3 1 873
0 113 7 1 2 871 875
0 114 5 1 1 113
0 115 7 2 2 869 114
0 116 5 2 1 878
0 117 7 1 2 867 880
0 118 5 1 1 117
0 119 7 2 2 865 118
0 120 5 1 1 882
0 121 7 1 2 53 120
0 122 5 2 1 121
0 123 7 1 2 745 883
0 124 5 2 1 123
0 125 7 1 2 837 886
0 126 5 1 1 125
0 127 7 2 2 884 126
0 128 5 1 1 888
0 129 7 1 2 54 128
0 130 5 2 1 129
0 131 7 1 2 747 889
0 132 5 2 1 131
0 133 7 1 2 839 892
0 134 5 1 1 133
0 135 7 2 2 890 134
0 136 5 1 1 894
0 137 7 1 2 55 136
0 138 5 2 1 137
0 139 7 1 2 749 895
0 140 5 2 1 139
0 141 7 1 2 841 898
0 142 5 1 1 141
0 143 7 2 2 896 142
0 144 5 1 1 900
0 145 7 1 2 56 144
0 146 5 2 1 145
0 147 7 1 2 751 901
0 148 5 2 1 147
0 149 7 1 2 843 904
0 150 5 1 1 149
0 151 7 2 2 902 150
0 152 5 1 1 906
0 153 7 1 2 57 152
0 154 5 2 1 153
0 155 7 1 2 753 907
0 156 5 2 1 155
0 157 7 1 2 845 910
0 158 5 1 1 157
0 159 7 2 2 908 158
0 160 5 1 1 912
0 161 7 1 2 58 160
0 162 5 2 1 161
0 163 7 1 2 755 913
0 164 5 2 1 163
0 165 7 1 2 847 916
0 166 5 1 1 165
0 167 7 2 2 914 166
0 168 5 1 1 918
0 169 7 1 2 59 168
0 170 5 2 1 169
0 171 7 1 2 757 919
0 172 5 2 1 171
0 173 7 1 2 849 922
0 174 5 1 1 173
0 175 7 2 2 920 174
0 176 5 1 1 924
0 177 7 1 2 60 176
0 178 5 2 1 177
0 179 7 1 2 759 925
0 180 5 2 1 179
0 181 7 1 2 851 928
0 182 5 1 1 181
0 183 7 2 2 926 182
0 184 5 1 1 930
0 185 7 1 2 61 184
0 186 5 2 1 185
0 187 7 1 2 761 931
0 188 5 2 1 187
0 189 7 1 2 853 934
0 190 5 1 1 189
0 191 7 2 2 932 190
0 192 5 1 1 936
0 193 7 1 2 62 192
0 194 5 2 1 193
0 195 7 1 2 763 937
0 196 5 2 1 195
0 197 7 1 2 855 940
0 198 5 1 1 197
0 199 7 2 2 938 198
0 200 5 1 1 942
0 201 7 1 2 63 200
0 202 5 2 1 201
0 203 7 1 2 765 943
0 204 5 2 1 203
0 205 7 1 2 857 946
0 206 5 1 1 205
0 207 7 2 2 944 206
0 208 5 1 1 948
0 209 7 1 2 64 208
0 210 5 2 1 209
0 211 7 1 2 767 949
0 212 5 2 1 211
0 213 7 1 2 859 952
0 214 5 1 1 213
0 215 7 2 2 950 214
0 216 5 2 1 954
0 217 7 1 2 863 956
0 218 5 1 1 217
0 219 7 2 2 861 218
0 220 5 1 1 958
0 221 7 2 2 836 220
0 222 5 3 1 960
0 223 7 2 2 98 959
0 224 5 2 1 965
0 225 7 2 2 862 864
0 226 5 1 1 969
0 227 7 1 2 955 226
0 228 5 1 1 227
0 229 7 1 2 957 970
0 230 5 1 1 229
0 231 7 2 2 228 230
0 232 5 1 1 971
0 233 7 1 2 97 232
0 234 5 4 1 233
0 235 7 1 2 834 972
0 236 5 3 1 235
0 237 7 2 2 951 953
0 238 5 1 1 980
0 239 7 1 2 799 981
0 240 5 1 1 239
0 241 7 1 2 860 238
0 242 5 1 1 241
0 243 7 2 2 240 242
0 244 5 1 1 982
0 245 7 1 2 832 244
0 246 5 4 1 245
0 247 7 1 2 96 983
0 248 5 3 1 247
0 249 7 2 2 945 947
0 250 5 1 1 991
0 251 7 1 2 797 992
0 252 5 1 1 251
0 253 7 1 2 858 250
0 254 5 1 1 253
0 255 7 2 2 252 254
0 256 5 1 1 993
0 257 7 1 2 830 256
0 258 5 4 1 257
0 259 7 1 2 95 994
0 260 5 3 1 259
0 261 7 2 2 939 941
0 262 5 1 1 1002
0 263 7 1 2 795 1003
0 264 5 1 1 263
0 265 7 1 2 856 262
0 266 5 1 1 265
0 267 7 2 2 264 266
0 268 5 1 1 1004
0 269 7 1 2 828 268
0 270 5 4 1 269
0 271 7 1 2 94 1005
0 272 5 3 1 271
0 273 7 2 2 933 935
0 274 5 1 1 1013
0 275 7 1 2 793 1014
0 276 5 1 1 275
0 277 7 1 2 854 274
0 278 5 1 1 277
0 279 7 2 2 276 278
0 280 5 1 1 1015
0 281 7 1 2 826 280
0 282 5 4 1 281
0 283 7 1 2 93 1016
0 284 5 3 1 283
0 285 7 2 2 927 929
0 286 5 1 1 1024
0 287 7 1 2 791 1025
0 288 5 1 1 287
0 289 7 1 2 852 286
0 290 5 1 1 289
0 291 7 2 2 288 290
0 292 5 1 1 1026
0 293 7 1 2 92 1027
0 294 5 3 1 293
0 295 7 1 2 824 292
0 296 5 4 1 295
0 297 7 2 2 921 923
0 298 5 1 1 1035
0 299 7 1 2 789 1036
0 300 5 1 1 299
0 301 7 1 2 850 298
0 302 5 1 1 301
0 303 7 2 2 300 302
0 304 5 1 1 1037
0 305 7 1 2 822 304
0 306 5 4 1 305
0 307 7 2 2 915 917
0 308 5 1 1 1043
0 309 7 1 2 787 1044
0 310 5 1 1 309
0 311 7 1 2 848 308
0 312 5 1 1 311
0 313 7 2 2 310 312
0 314 5 1 1 1045
0 315 7 1 2 820 314
0 316 5 3 1 315
0 317 7 2 2 909 911
0 318 5 1 1 1050
0 319 7 1 2 785 1051
0 320 5 1 1 319
0 321 7 1 2 846 318
0 322 5 1 1 321
0 323 7 2 2 320 322
0 324 5 1 1 1052
0 325 7 1 2 818 324
0 326 5 4 1 325
0 327 7 1 2 89 1053
0 328 5 3 1 327
0 329 7 2 2 903 905
0 330 5 1 1 1061
0 331 7 1 2 783 1062
0 332 5 1 1 331
0 333 7 1 2 844 330
0 334 5 1 1 333
0 335 7 2 2 332 334
0 336 5 1 1 1063
0 337 7 2 2 816 336
0 338 5 4 1 1065
0 339 7 2 2 897 899
0 340 5 1 1 1071
0 341 7 1 2 781 1072
0 342 5 1 1 341
0 343 7 1 2 842 340
0 344 5 1 1 343
0 345 7 2 2 342 344
0 346 5 1 1 1073
0 347 7 1 2 814 346
0 348 5 3 1 347
0 349 7 1 2 87 1074
0 350 5 3 1 349
0 351 7 2 2 891 893
0 352 5 1 1 1081
0 353 7 1 2 779 1082
0 354 5 1 1 353
0 355 7 1 2 840 352
0 356 5 1 1 355
0 357 7 2 2 354 356
0 358 5 1 1 1083
0 359 7 1 2 812 358
0 360 5 4 1 359
0 361 7 1 2 86 1084
0 362 5 4 1 361
0 363 7 2 2 885 887
0 364 5 1 1 1093
0 365 7 1 2 777 1094
0 366 5 1 1 365
0 367 7 1 2 838 364
0 368 5 1 1 367
0 369 7 2 2 366 368
0 370 5 1 1 1095
0 371 7 1 2 85 1096
0 372 5 3 1 371
0 373 7 1 2 810 370
0 374 5 3 1 373
0 375 7 2 2 866 868
0 376 5 1 1 1103
0 377 7 1 2 879 376
0 378 5 1 1 377
0 379 7 1 2 881 1104
0 380 5 1 1 379
0 381 7 2 2 378 380
0 382 5 1 1 1105
0 383 7 1 2 84 382
0 384 5 3 1 383
0 385 7 1 2 808 1106
0 386 5 3 1 385
0 387 7 2 2 870 872
0 388 5 2 1 1113
0 389 7 1 2 874 1115
0 390 5 1 1 389
0 391 7 1 2 876 1114
0 392 5 1 1 391
0 393 7 2 2 390 392
0 394 5 1 1 1117
0 395 7 1 2 805 1118
0 396 5 1 1 395
0 397 7 1 2 83 394
0 398 5 2 1 397
0 399 7 1 2 50 66
0 400 5 1 1 399
0 401 7 2 2 877 400
0 402 5 1 1 1121
0 403 7 1 2 803 402
0 404 7 1 2 1119 403
0 405 5 1 1 404
0 406 7 3 2 396 405
0 407 5 1 1 1123
0 408 7 1 2 1110 1124
0 409 5 1 1 408
0 410 7 2 2 1107 409
0 411 5 2 1 1126
0 412 7 1 2 1100 1128
0 413 5 1 1 412
0 414 7 2 2 1097 413
0 415 5 1 1 1130
0 416 7 2 2 1089 1131
0 417 5 1 1 1132
0 418 7 2 2 1085 417
0 419 5 2 1 1134
0 420 7 1 2 1078 1136
0 421 5 1 1 420
0 422 7 2 2 1075 421
0 423 7 1 2 1067 1138
0 424 5 1 1 423
0 425 7 2 2 88 1064
0 426 5 3 1 1140
0 427 7 1 2 424 1142
0 428 7 2 2 1058 427
0 429 5 1 1 1145
0 430 7 2 2 1054 429
0 431 5 2 1 1147
0 432 7 1 2 90 1046
0 433 5 3 1 432
0 434 7 1 2 1149 1151
0 435 5 1 1 434
0 436 7 2 2 1047 435
0 437 5 1 1 1154
0 438 7 1 2 91 1038
0 439 5 3 1 438
0 440 7 1 2 437 1156
0 441 5 2 1 440
0 442 7 1 2 1039 1159
0 443 7 1 2 1031 442
0 444 5 1 1 443
0 445 7 1 2 1028 444
0 446 7 1 2 1021 445
0 447 5 2 1 446
0 448 7 1 2 1017 1161
0 449 5 1 1 448
0 450 7 1 2 1010 449
0 451 5 1 1 450
0 452 7 1 2 1006 451
0 453 5 1 1 452
0 454 7 2 2 999 453
0 455 5 1 1 1163
0 456 7 2 2 995 455
0 457 5 1 1 1165
0 458 7 1 2 988 457
0 459 5 1 1 458
0 460 7 2 2 984 459
0 461 5 1 1 1167
0 462 7 1 2 977 1168
0 463 5 1 1 462
0 464 7 2 2 973 463
0 465 5 1 1 1169
0 466 7 1 2 967 1170
0 467 5 1 1 466
0 468 7 2 2 962 467
0 469 5 1 1 1171
0 470 7 1 2 966 465
0 471 5 1 1 470
0 472 7 2 2 974 978
0 473 5 2 1 1173
0 474 7 1 2 985 1175
0 475 5 1 1 474
0 476 7 1 2 461 1174
0 477 5 1 1 476
0 478 7 2 2 986 989
0 479 5 2 1 1177
0 480 7 1 2 1166 1179
0 481 5 1 1 480
0 482 7 2 2 996 1000
0 483 5 2 1 1181
0 484 7 1 2 1007 1183
0 485 5 1 1 484
0 486 7 1 2 997 1164
0 487 5 1 1 486
0 488 7 3 2 1008 1011
0 489 5 1 1 1185
0 490 7 1 2 1162 1186
0 491 5 1 1 490
0 492 7 1 2 1018 491
0 493 5 1 1 492
0 494 7 2 2 1019 1022
0 495 5 2 1 1188
0 496 7 1 2 1032 1190
0 497 5 1 1 496
0 498 7 3 2 1029 1033
0 499 5 1 1 1192
0 500 7 1 2 1160 1193
0 501 5 1 1 500
0 502 7 1 2 1040 501
0 503 5 1 1 502
0 504 7 2 2 1041 1157
0 505 5 2 1 1195
0 506 7 1 2 1155 1197
0 507 5 1 1 506
0 508 7 3 2 1048 1152
0 509 5 2 1 1199
0 510 7 1 2 1148 1200
0 511 5 1 1 510
0 512 7 2 2 1055 1059
0 513 5 2 1 1204
0 514 7 1 2 1068 1206
0 515 5 1 1 514
0 516 7 1 2 1056 1146
0 517 5 1 1 516
0 518 7 3 2 1076 1079
0 519 5 2 1 1208
0 520 7 1 2 1135 1209
0 521 5 1 1 520
0 522 7 1 2 1086 1133
0 523 5 1 1 522
0 524 7 1 2 1087 1090
0 525 5 2 1 524
0 526 7 1 2 415 1213
0 527 5 1 1 526
0 528 7 3 2 1098 1101
0 529 5 2 1 1215
0 530 7 1 2 1129 1216
0 531 5 1 1 530
0 532 7 1 2 1127 1218
0 533 5 1 1 532
0 534 7 3 2 1108 1111
0 535 5 2 1 1220
0 536 7 1 2 1125 1221
0 537 5 1 1 536
0 538 7 1 2 407 1223
0 539 5 1 1 538
0 540 7 1 2 537 539
0 541 7 1 2 533 540
0 542 7 1 2 531 541
0 543 5 1 1 542
0 544 7 1 2 527 543
0 545 7 1 2 523 544
0 546 5 1 1 545
0 547 7 1 2 1137 1211
0 548 5 1 1 547
0 549 7 1 2 546 548
0 550 7 1 2 521 549
0 551 5 1 1 550
0 552 7 1 2 1069 1143
0 553 5 1 1 552
0 554 7 1 2 1139 553
0 555 5 1 1 554
0 556 7 1 2 551 555
0 557 7 1 2 517 556
0 558 7 1 2 515 557
0 559 5 1 1 558
0 560 7 1 2 1150 1202
0 561 5 1 1 560
0 562 7 1 2 559 561
0 563 7 1 2 511 562
0 564 5 1 1 563
0 565 7 1 2 507 564
0 566 7 1 2 503 565
0 567 7 1 2 497 566
0 568 7 1 2 493 567
0 569 7 1 2 487 568
0 570 7 1 2 485 569
0 571 7 1 2 963 570
0 572 7 1 2 481 571
0 573 7 1 2 477 572
0 574 7 1 2 475 573
0 575 7 1 2 471 574
0 576 7 1 2 1172 575
0 577 5 1 1 576
0 578 7 1 2 806 1116
0 579 5 1 1 578
0 580 7 1 2 82 1122
0 581 7 1 2 579 580
0 582 5 1 1 581
0 583 7 2 2 1120 582
0 584 5 2 1 1225
0 585 7 1 2 1112 1227
0 586 5 1 1 585
0 587 7 3 2 1109 586
0 588 5 1 1 1229
0 589 7 1 2 1099 1230
0 590 5 1 1 589
0 591 7 2 2 1102 590
0 592 5 1 1 1232
0 593 7 2 2 1088 1233
0 594 5 1 1 1234
0 595 7 3 2 1091 594
0 596 5 1 1 1236
0 597 7 1 2 1080 1237
0 598 5 1 1 597
0 599 7 2 2 1077 598
0 600 5 2 1 1239
0 601 7 1 2 1144 1241
0 602 5 1 1 601
0 603 7 2 2 1070 602
0 604 5 1 1 1243
0 605 7 1 2 1060 604
0 606 5 1 1 605
0 607 7 2 2 1057 606
0 608 5 2 1 1245
0 609 7 1 2 1153 1247
0 610 5 1 1 609
0 611 7 2 2 1049 610
0 612 5 2 1 1249
0 613 7 1 2 1158 1251
0 614 5 1 1 613
0 615 7 2 2 1042 614
0 616 5 2 1 1253
0 617 7 1 2 1030 1255
0 618 5 1 1 617
0 619 7 2 2 1034 618
0 620 5 2 1 1257
0 621 7 1 2 1023 1259
0 622 5 1 1 621
0 623 7 2 2 1020 622
0 624 5 2 1 1261
0 625 7 1 2 1012 1263
0 626 5 1 1 625
0 627 7 2 2 1009 626
0 628 5 2 1 1265
0 629 7 1 2 1001 1267
0 630 5 1 1 629
0 631 7 2 2 998 630
0 632 5 2 1 1269
0 633 7 1 2 990 1271
0 634 5 1 1 633
0 635 7 1 2 987 634
0 636 5 2 1 635
0 637 7 1 2 975 1273
0 638 5 1 1 637
0 639 7 1 2 979 964
0 640 7 1 2 638 639
0 641 5 1 1 640
0 642 7 1 2 1176 1274
0 643 5 1 1 642
0 644 7 1 2 976 961
0 645 5 1 1 644
0 646 7 1 2 1184 1266
0 647 5 1 1 646
0 648 7 1 2 1182 1268
0 649 5 1 1 648
0 650 7 1 2 647 649
0 651 5 1 1 650
0 652 7 1 2 1187 1262
0 653 5 1 1 652
0 654 7 1 2 489 1264
0 655 5 1 1 654
0 656 7 1 2 1191 1260
0 657 5 1 1 656
0 658 7 1 2 1189 1258
0 659 5 1 1 658
0 660 7 1 2 1194 1256
0 661 5 1 1 660
0 662 7 1 2 499 1254
0 663 5 1 1 662
0 664 7 1 2 661 663
0 665 5 1 1 664
0 666 7 1 2 1205 1244
0 667 5 1 1 666
0 668 7 1 2 1141 1240
0 669 5 1 1 668
0 670 7 1 2 1207 669
0 671 5 1 1 670
0 672 7 1 2 1066 1242
0 673 5 1 1 672
0 674 7 1 2 1210 1238
0 675 5 1 1 674
0 676 7 1 2 1092 1235
0 677 5 1 1 676
0 678 7 1 2 1214 592
0 679 5 1 1 678
0 680 7 1 2 1217 1231
0 681 5 1 1 680
0 682 7 1 2 1224 1226
0 683 5 1 1 682
0 684 7 1 2 1222 1228
0 685 5 1 1 684
0 686 7 1 2 683 685
0 687 5 1 1 686
0 688 7 1 2 1219 588
0 689 5 1 1 688
0 690 7 1 2 687 689
0 691 7 1 2 681 690
0 692 5 1 1 691
0 693 7 1 2 679 692
0 694 7 1 2 677 693
0 695 5 1 1 694
0 696 7 1 2 1212 596
0 697 5 1 1 696
0 698 7 1 2 695 697
0 699 7 1 2 675 698
0 700 5 1 1 699
0 701 7 1 2 673 700
0 702 7 1 2 671 701
0 703 7 1 2 667 702
0 704 5 1 1 703
0 705 7 1 2 1203 1248
0 706 5 1 1 705
0 707 7 1 2 1201 1246
0 708 5 1 1 707
0 709 7 1 2 706 708
0 710 5 1 1 709
0 711 7 1 2 704 710
0 712 5 1 1 711
0 713 7 1 2 1196 1252
0 714 5 1 1 713
0 715 7 1 2 1198 1250
0 716 5 1 1 715
0 717 7 1 2 714 716
0 718 5 1 1 717
0 719 7 1 2 712 718
0 720 7 1 2 665 719
0 721 7 1 2 659 720
0 722 7 1 2 657 721
0 723 7 1 2 655 722
0 724 7 1 2 653 723
0 725 7 1 2 651 724
0 726 7 1 2 968 725
0 727 7 1 2 645 726
0 728 7 1 2 1180 1272
0 729 5 1 1 728
0 730 7 1 2 1178 1270
0 731 5 1 1 730
0 732 7 1 2 729 731
0 733 7 1 2 727 732
0 734 7 1 2 643 733
0 735 7 1 2 641 734
0 736 7 1 2 469 735
0 737 5 1 1 736
0 738 7 1 2 577 737
3 1499 5 0 1 738
