1 0 0 2 0
2 13 1 0
2 172 1 0
1 1 0 2 0
2 173 1 1
2 174 1 1
1 2 0 2 0
2 175 1 2
2 176 1 2
1 3 0 2 0
2 177 1 3
2 178 1 3
1 4 0 2 0
2 179 1 4
2 180 1 4
1 5 0 2 0
2 181 1 5
2 182 1 5
1 6 0 2 0
2 183 1 6
2 184 1 6
1 7 0 2 0
2 185 1 7
2 186 1 7
1 8 0 2 0
2 187 1 8
2 188 1 8
1 9 0 2 0
2 189 1 9
2 190 1 9
1 10 0 2 0
2 191 1 10
2 192 1 10
1 11 0 2 0
2 193 1 11
2 194 1 11
1 12 0 2 0
2 195 1 12
2 196 1 12
2 197 1 28
2 198 1 28
2 199 1 30
2 200 1 30
2 201 1 32
2 202 1 32
2 203 1 34
2 204 1 34
2 205 1 36
2 206 1 36
2 207 1 38
2 208 1 38
2 209 1 39
2 210 1 39
2 211 1 40
2 212 1 40
2 213 1 40
2 214 1 43
2 215 1 43
2 216 1 44
2 217 1 44
2 218 1 47
2 219 1 47
2 220 1 48
2 221 1 48
2 222 1 51
2 223 1 51
2 224 1 53
2 225 1 53
2 226 1 54
2 227 1 54
2 228 1 55
2 229 1 55
2 230 1 61
2 231 1 61
2 232 1 64
2 233 1 64
2 234 1 64
2 235 1 66
2 236 1 66
2 237 1 66
2 238 1 67
2 239 1 67
2 240 1 73
2 241 1 73
2 242 1 76
2 243 1 76
2 244 1 76
2 245 1 78
2 246 1 78
2 247 1 78
2 248 1 79
2 249 1 79
2 250 1 85
2 251 1 85
2 252 1 88
2 253 1 88
2 254 1 90
2 255 1 90
2 256 1 93
2 257 1 93
2 258 1 98
2 259 1 98
2 260 1 99
2 261 1 99
2 262 1 102
2 263 1 102
2 264 1 103
2 265 1 103
2 266 1 106
2 267 1 106
2 268 1 114
2 269 1 114
2 270 1 115
2 271 1 115
2 272 1 120
2 273 1 120
2 274 1 121
2 275 1 121
2 276 1 124
2 277 1 124
2 278 1 125
2 279 1 125
2 280 1 128
2 281 1 128
2 282 1 132
2 283 1 132
2 284 1 134
2 285 1 134
2 286 1 134
2 287 1 135
2 288 1 135
2 289 1 142
2 290 1 142
2 291 1 143
2 292 1 143
2 293 1 145
2 294 1 145
0 14 5 1 1 13
0 15 5 1 1 173
0 16 5 1 1 175
0 17 5 1 1 177
0 18 5 1 1 179
0 19 5 1 1 181
0 20 5 1 1 183
0 21 5 1 1 185
0 22 5 1 1 187
0 23 5 1 1 189
0 24 5 1 1 191
0 25 5 1 1 193
0 26 5 1 1 195
0 27 7 1 2 17 21
0 28 5 2 1 27
0 29 7 1 2 178 186
0 30 5 2 1 29
0 31 7 1 2 16 20
0 32 5 2 1 31
0 33 7 1 2 176 184
0 34 5 2 1 33
0 35 7 1 2 15 19
0 36 5 2 1 35
0 37 7 1 2 174 182
0 38 5 2 1 37
0 39 7 2 2 172 180
0 40 5 3 1 209
0 41 7 1 2 207 211
0 42 5 1 1 41
0 43 7 2 2 205 42
0 44 5 2 1 214
0 45 7 1 2 203 216
0 46 5 1 1 45
0 47 7 2 2 201 46
0 48 5 2 1 218
0 49 7 1 2 199 220
0 50 5 1 1 49
0 51 7 2 2 197 50
0 52 5 1 1 222
0 53 7 2 2 196 52
0 54 5 2 1 224
0 55 7 2 2 198 200
0 56 5 1 1 228
0 57 7 1 2 219 56
0 58 5 1 1 57
0 59 7 1 2 221 229
0 60 5 1 1 59
0 61 7 2 2 58 60
0 62 5 1 1 230
0 63 7 1 2 25 62
0 64 5 3 1 63
0 65 7 1 2 194 231
0 66 5 3 1 65
0 67 7 2 2 202 204
0 68 5 1 1 238
0 69 7 1 2 215 68
0 70 5 1 1 69
0 71 7 1 2 217 239
0 72 5 1 1 71
0 73 7 2 2 70 72
0 74 5 1 1 240
0 75 7 1 2 24 74
0 76 5 3 1 75
0 77 7 1 2 192 241
0 78 5 3 1 77
0 79 7 2 2 206 208
0 80 5 1 1 248
0 81 7 1 2 210 80
0 82 5 1 1 81
0 83 7 1 2 212 249
0 84 5 1 1 83
0 85 7 2 2 82 84
0 86 5 1 1 250
0 87 7 1 2 190 251
0 88 5 2 1 87
0 89 7 1 2 23 86
0 90 5 2 1 89
0 91 7 1 2 14 18
0 92 5 1 1 91
0 93 7 2 2 213 92
0 94 5 1 1 256
0 95 7 1 2 22 257
0 96 5 1 1 95
0 97 7 1 2 254 96
0 98 5 2 1 97
0 99 7 2 2 252 258
0 100 7 1 2 245 260
0 101 5 1 1 100
0 102 7 2 2 242 101
0 103 5 2 1 262
0 104 7 1 2 235 264
0 105 5 1 1 104
0 106 7 2 2 232 105
0 107 5 1 1 266
0 108 7 1 2 226 267
0 109 5 1 1 108
0 110 7 1 2 225 107
0 111 5 1 1 110
0 112 7 1 2 109 111
0 113 5 1 1 112
0 114 7 2 2 26 223
0 115 5 2 1 268
0 116 7 1 2 188 94
0 117 5 1 1 116
0 118 7 1 2 253 117
0 119 5 1 1 118
0 120 7 2 2 255 119
0 121 5 2 1 272
0 122 7 1 2 246 274
0 123 5 1 1 122
0 124 7 2 2 243 123
0 125 5 2 1 276
0 126 7 1 2 236 278
0 127 5 1 1 126
0 128 7 2 2 233 127
0 129 5 1 1 280
0 130 7 1 2 270 281
0 131 5 1 1 130
0 132 7 2 2 227 131
0 133 5 1 1 282
0 134 7 3 2 234 237
0 135 5 2 1 284
0 136 7 1 2 265 287
0 137 5 1 1 136
0 138 7 1 2 263 285
0 139 5 1 1 138
0 140 7 1 2 137 139
0 141 5 1 1 140
0 142 7 2 2 244 247
0 143 5 2 1 289
0 144 7 1 2 273 291
0 145 5 2 1 144
0 146 7 1 2 261 290
0 147 5 1 1 146
0 148 7 1 2 271 147
0 149 7 1 2 293 148
0 150 7 1 2 141 149
0 151 7 1 2 133 150
0 152 7 1 2 113 151
0 153 5 1 1 152
0 154 7 1 2 269 129
0 155 5 1 1 154
0 156 7 1 2 277 286
0 157 5 1 1 156
0 158 7 1 2 259 292
0 159 5 1 1 158
0 160 7 1 2 275 159
0 161 5 1 1 160
0 162 7 1 2 294 161
0 163 5 1 1 162
0 164 7 1 2 279 288
0 165 5 1 1 164
0 166 7 1 2 163 165
0 167 7 1 2 157 166
0 168 7 1 2 155 167
0 169 7 1 2 283 168
0 170 5 1 1 169
0 171 7 1 2 153 170
3 399 5 0 1 171
