1 0 0 2 0
2 64 1 0
2 65 1 0
1 1 0 2 0
2 66 1 1
2 67 1 1
1 2 0 2 0
2 68 1 2
2 69 1 2
1 3 0 2 0
2 70 1 3
2 71 1 3
1 4 0 2 0
2 72 1 4
2 73 1 4
1 5 0 2 0
2 74 1 5
2 75 1 5
1 6 0 2 0
2 76 1 6
2 77 1 6
1 7 0 2 0
2 78 1 7
2 79 1 7
1 8 0 2 0
2 80 1 8
2 81 1 8
1 9 0 2 0
2 82 1 9
2 83 1 9
1 10 0 2 0
2 84 1 10
2 85 1 10
1 11 0 2 0
2 86 1 11
2 87 1 11
1 12 0 2 0
2 88 1 12
2 89 1 12
1 13 0 2 0
2 90 1 13
2 91 1 13
1 14 0 2 0
2 92 1 14
2 93 1 14
1 15 0 2 0
2 94 1 15
2 95 1 15
1 16 0 2 0
2 96 1 16
2 165 1 16
1 17 0 2 0
2 176 1 17
2 189 1 17
1 18 0 2 0
2 208 1 18
2 228 1 18
1 19 0 2 0
2 251 1 19
2 275 1 19
1 20 0 2 0
2 299 1 20
2 324 1 20
1 21 0 2 0
2 349 1 21
2 374 1 21
1 22 0 2 0
2 399 1 22
2 427 1 22
1 23 0 2 0
2 455 1 23
2 483 1 23
1 24 0 2 0
2 512 1 24
2 542 1 24
1 25 0 2 0
2 572 1 25
2 602 1 25
1 26 0 2 0
2 632 1 26
2 662 1 26
1 27 0 2 0
2 692 1 27
2 722 1 27
1 28 0 2 0
2 752 1 28
2 785 1 28
1 29 0 2 0
2 817 1 29
2 849 1 29
1 30 0 2 0
2 882 1 30
2 915 1 30
1 31 0 2 0
2 948 1 31
2 981 1 31
1 32 0 2 0
2 1012 1 32
2 1033 1 32
1 33 0 2 0
2 1034 1 33
2 1035 1 33
1 34 0 2 0
2 1036 1 34
2 1037 1 34
1 35 0 2 0
2 1038 1 35
2 1039 1 35
1 36 0 2 0
2 1040 1 36
2 1041 1 36
1 37 0 2 0
2 1042 1 37
2 1043 1 37
1 38 0 2 0
2 1044 1 38
2 1045 1 38
1 39 0 2 0
2 1046 1 39
2 1047 1 39
1 40 0 2 0
2 1048 1 40
2 1049 1 40
1 41 0 2 0
2 1050 1 41
2 1051 1 41
1 42 0 2 0
2 1052 1 42
2 1053 1 42
1 43 0 2 0
2 1054 1 43
2 1055 1 43
1 44 0 2 0
2 1056 1 44
2 1057 1 44
1 45 0 2 0
2 1058 1 45
2 1059 1 45
1 46 0 2 0
2 1060 1 46
2 1061 1 46
1 47 0 2 0
2 1062 1 47
2 1063 1 47
1 48 0 2 0
2 1064 1 48
2 1065 1 48
1 49 0 2 0
2 1066 1 49
2 1067 1 49
1 50 0 2 0
2 1068 1 50
2 1069 1 50
1 51 0 2 0
2 1070 1 51
2 1071 1 51
1 52 0 2 0
2 1072 1 52
2 1073 1 52
1 53 0 2 0
2 1074 1 53
2 1075 1 53
1 54 0 2 0
2 1076 1 54
2 1077 1 54
1 55 0 2 0
2 1078 1 55
2 1079 1 55
1 56 0 2 0
2 1080 1 56
2 1081 1 56
1 57 0 2 0
2 1082 1 57
2 1083 1 57
1 58 0 2 0
2 1084 1 58
2 1085 1 58
1 59 0 2 0
2 1086 1 59
2 1087 1 59
1 60 0 2 0
2 1088 1 60
2 1089 1 60
1 61 0 2 0
2 1090 1 61
2 1091 1 61
1 62 0 2 0
2 1092 1 62
2 1093 1 62
1 63 0 2 0
2 1094 1 63
2 1095 1 63
2 1096 1 161
2 1097 1 161
2 1098 1 162
2 1099 1 162
2 1100 1 167
2 1101 1 167
2 1102 1 167
2 1103 1 170
2 1104 1 170
2 1105 1 172
2 1106 1 172
2 1107 1 173
2 1108 1 173
2 1109 1 177
2 1110 1 177
2 1111 1 178
2 1112 1 178
2 1113 1 178
2 1114 1 180
2 1115 1 180
2 1116 1 180
2 1117 1 182
2 1118 1 182
2 1119 1 183
2 1120 1 183
2 1121 1 183
2 1122 1 183
2 1123 1 190
2 1124 1 190
2 1125 1 194
2 1126 1 194
2 1127 1 196
2 1128 1 196
2 1129 1 197
2 1130 1 197
2 1131 1 199
2 1132 1 199
2 1133 1 199
2 1134 1 201
2 1135 1 201
2 1136 1 202
2 1137 1 202
2 1138 1 202
2 1139 1 202
2 1140 1 209
2 1141 1 209
2 1142 1 214
2 1143 1 214
2 1144 1 216
2 1145 1 216
2 1146 1 217
2 1147 1 217
2 1148 1 219
2 1149 1 219
2 1150 1 219
2 1151 1 221
2 1152 1 221
2 1153 1 222
2 1154 1 222
2 1155 1 222
2 1156 1 222
2 1157 1 229
2 1158 1 229
2 1159 1 229
2 1160 1 236
2 1161 1 236
2 1162 1 239
2 1163 1 239
2 1164 1 240
2 1165 1 240
2 1166 1 242
2 1167 1 242
2 1168 1 242
2 1169 1 244
2 1170 1 244
2 1171 1 245
2 1172 1 245
2 1173 1 245
2 1174 1 245
2 1175 1 252
2 1176 1 252
2 1177 1 252
2 1178 1 260
2 1179 1 260
2 1180 1 263
2 1181 1 263
2 1182 1 264
2 1183 1 264
2 1184 1 266
2 1185 1 266
2 1186 1 266
2 1187 1 268
2 1188 1 268
2 1189 1 269
2 1190 1 269
2 1191 1 269
2 1192 1 269
2 1193 1 276
2 1194 1 276
2 1195 1 276
2 1196 1 284
2 1197 1 284
2 1198 1 287
2 1199 1 287
2 1200 1 288
2 1201 1 288
2 1202 1 288
2 1203 1 290
2 1204 1 290
2 1205 1 290
2 1206 1 292
2 1207 1 292
2 1208 1 293
2 1209 1 293
2 1210 1 293
2 1211 1 293
2 1212 1 300
2 1213 1 300
2 1214 1 300
2 1215 1 305
2 1216 1 305
2 1217 1 307
2 1218 1 307
2 1219 1 310
2 1220 1 310
2 1221 1 312
2 1222 1 312
2 1223 1 313
2 1224 1 313
2 1225 1 315
2 1226 1 315
2 1227 1 315
2 1228 1 317
2 1229 1 317
2 1230 1 318
2 1231 1 318
2 1232 1 318
2 1233 1 318
2 1234 1 326
2 1235 1 326
2 1236 1 326
2 1237 1 328
2 1238 1 328
2 1239 1 329
2 1240 1 329
2 1241 1 329
2 1242 1 329
2 1243 1 331
2 1244 1 331
2 1245 1 331
2 1246 1 336
2 1247 1 336
2 1248 1 338
2 1249 1 338
2 1250 1 341
2 1251 1 341
2 1252 1 343
2 1253 1 343
2 1254 1 344
2 1255 1 344
2 1256 1 351
2 1257 1 351
2 1258 1 351
2 1259 1 353
2 1260 1 353
2 1261 1 354
2 1262 1 354
2 1263 1 354
2 1264 1 354
2 1265 1 356
2 1266 1 356
2 1267 1 356
2 1268 1 361
2 1269 1 361
2 1270 1 363
2 1271 1 363
2 1272 1 366
2 1273 1 366
2 1274 1 368
2 1275 1 368
2 1276 1 369
2 1277 1 369
2 1278 1 376
2 1279 1 376
2 1280 1 376
2 1281 1 378
2 1282 1 378
2 1283 1 379
2 1284 1 379
2 1285 1 379
2 1286 1 379
2 1287 1 381
2 1288 1 381
2 1289 1 381
2 1290 1 386
2 1291 1 386
2 1292 1 388
2 1293 1 388
2 1294 1 390
2 1295 1 390
2 1296 1 393
2 1297 1 393
2 1298 1 394
2 1299 1 394
2 1300 1 394
2 1301 1 400
2 1302 1 400
2 1303 1 400
2 1304 1 401
2 1305 1 401
2 1306 1 401
2 1307 1 408
2 1308 1 408
2 1309 1 410
2 1310 1 410
2 1311 1 415
2 1312 1 415
2 1313 1 416
2 1314 1 416
2 1315 1 416
2 1316 1 418
2 1317 1 418
2 1318 1 418
2 1319 1 420
2 1320 1 420
2 1321 1 421
2 1322 1 421
2 1323 1 421
2 1324 1 421
2 1325 1 428
2 1326 1 428
2 1327 1 428
2 1328 1 429
2 1329 1 429
2 1330 1 429
2 1331 1 436
2 1332 1 436
2 1333 1 438
2 1334 1 438
2 1335 1 443
2 1336 1 443
2 1337 1 444
2 1338 1 444
2 1339 1 444
2 1340 1 446
2 1341 1 446
2 1342 1 446
2 1343 1 448
2 1344 1 448
2 1345 1 449
2 1346 1 449
2 1347 1 449
2 1348 1 449
2 1349 1 456
2 1350 1 456
2 1351 1 456
2 1352 1 457
2 1353 1 457
2 1354 1 457
2 1355 1 464
2 1356 1 464
2 1357 1 466
2 1358 1 466
2 1359 1 471
2 1360 1 471
2 1361 1 472
2 1362 1 472
2 1363 1 472
2 1364 1 474
2 1365 1 474
2 1366 1 474
2 1367 1 476
2 1368 1 476
2 1369 1 477
2 1370 1 477
2 1371 1 477
2 1372 1 477
2 1373 1 484
2 1374 1 484
2 1375 1 484
2 1376 1 485
2 1377 1 485
2 1378 1 485
2 1379 1 493
2 1380 1 493
2 1381 1 495
2 1382 1 495
2 1383 1 500
2 1384 1 500
2 1385 1 501
2 1386 1 501
2 1387 1 501
2 1388 1 503
2 1389 1 503
2 1390 1 503
2 1391 1 505
2 1392 1 505
2 1393 1 506
2 1394 1 506
2 1395 1 506
2 1396 1 506
2 1397 1 513
2 1398 1 513
2 1399 1 513
2 1400 1 518
2 1401 1 518
2 1402 1 520
2 1403 1 520
2 1404 1 522
2 1405 1 522
2 1406 1 522
2 1407 1 525
2 1408 1 525
2 1409 1 528
2 1410 1 528
2 1411 1 530
2 1412 1 530
2 1413 1 531
2 1414 1 531
2 1415 1 533
2 1416 1 533
2 1417 1 533
2 1418 1 535
2 1419 1 535
2 1420 1 536
2 1421 1 536
2 1422 1 536
2 1423 1 536
2 1424 1 543
2 1425 1 543
2 1426 1 543
2 1427 1 548
2 1428 1 548
2 1429 1 550
2 1430 1 550
2 1431 1 552
2 1432 1 552
2 1433 1 552
2 1434 1 555
2 1435 1 555
2 1436 1 558
2 1437 1 558
2 1438 1 560
2 1439 1 560
2 1440 1 563
2 1441 1 563
2 1442 1 563
2 1443 1 565
2 1444 1 565
2 1445 1 566
2 1446 1 566
2 1447 1 566
2 1448 1 566
2 1449 1 573
2 1450 1 573
2 1451 1 573
2 1452 1 578
2 1453 1 578
2 1454 1 580
2 1455 1 580
2 1456 1 582
2 1457 1 582
2 1458 1 582
2 1459 1 585
2 1460 1 585
2 1461 1 588
2 1462 1 588
2 1463 1 590
2 1464 1 590
2 1465 1 593
2 1466 1 593
2 1467 1 593
2 1468 1 595
2 1469 1 595
2 1470 1 596
2 1471 1 596
2 1472 1 596
2 1473 1 596
2 1474 1 603
2 1475 1 603
2 1476 1 603
2 1477 1 608
2 1478 1 608
2 1479 1 610
2 1480 1 610
2 1481 1 612
2 1482 1 612
2 1483 1 612
2 1484 1 615
2 1485 1 615
2 1486 1 617
2 1487 1 617
2 1488 1 620
2 1489 1 620
2 1490 1 623
2 1491 1 623
2 1492 1 623
2 1493 1 625
2 1494 1 625
2 1495 1 626
2 1496 1 626
2 1497 1 626
2 1498 1 626
2 1499 1 633
2 1500 1 633
2 1501 1 633
2 1502 1 638
2 1503 1 638
2 1504 1 640
2 1505 1 640
2 1506 1 642
2 1507 1 642
2 1508 1 642
2 1509 1 645
2 1510 1 645
2 1511 1 647
2 1512 1 647
2 1513 1 650
2 1514 1 650
2 1515 1 653
2 1516 1 653
2 1517 1 653
2 1518 1 655
2 1519 1 655
2 1520 1 656
2 1521 1 656
2 1522 1 656
2 1523 1 656
2 1524 1 663
2 1525 1 663
2 1526 1 663
2 1527 1 668
2 1528 1 668
2 1529 1 670
2 1530 1 670
2 1531 1 672
2 1532 1 672
2 1533 1 672
2 1534 1 675
2 1535 1 675
2 1536 1 677
2 1537 1 677
2 1538 1 680
2 1539 1 680
2 1540 1 683
2 1541 1 683
2 1542 1 683
2 1543 1 685
2 1544 1 685
2 1545 1 686
2 1546 1 686
2 1547 1 686
2 1548 1 686
2 1549 1 693
2 1550 1 693
2 1551 1 693
2 1552 1 698
2 1553 1 698
2 1554 1 700
2 1555 1 700
2 1556 1 702
2 1557 1 702
2 1558 1 702
2 1559 1 705
2 1560 1 705
2 1561 1 707
2 1562 1 707
2 1563 1 710
2 1564 1 710
2 1565 1 713
2 1566 1 713
2 1567 1 713
2 1568 1 715
2 1569 1 715
2 1570 1 716
2 1571 1 716
2 1572 1 716
2 1573 1 716
2 1574 1 723
2 1575 1 723
2 1576 1 723
2 1577 1 728
2 1578 1 728
2 1579 1 730
2 1580 1 730
2 1581 1 732
2 1582 1 732
2 1583 1 732
2 1584 1 735
2 1585 1 735
2 1586 1 737
2 1587 1 737
2 1588 1 740
2 1589 1 740
2 1590 1 743
2 1591 1 743
2 1592 1 743
2 1593 1 745
2 1594 1 745
2 1595 1 746
2 1596 1 746
2 1597 1 746
2 1598 1 746
2 1599 1 753
2 1600 1 753
2 1601 1 753
2 1602 1 753
2 1603 1 754
2 1604 1 754
2 1605 1 754
2 1606 1 755
2 1607 1 755
2 1608 1 755
2 1609 1 762
2 1610 1 762
2 1611 1 764
2 1612 1 764
2 1613 1 768
2 1614 1 768
2 1615 1 773
2 1616 1 773
2 1617 1 776
2 1618 1 776
2 1619 1 776
2 1620 1 778
2 1621 1 778
2 1622 1 779
2 1623 1 779
2 1624 1 779
2 1625 1 779
2 1626 1 787
2 1627 1 787
2 1628 1 787
2 1629 1 789
2 1630 1 789
2 1631 1 790
2 1632 1 790
2 1633 1 790
2 1634 1 790
2 1635 1 792
2 1636 1 792
2 1637 1 792
2 1638 1 793
2 1639 1 793
2 1640 1 793
2 1641 1 794
2 1642 1 794
2 1643 1 805
2 1644 1 805
2 1645 1 807
2 1646 1 807
2 1647 1 811
2 1648 1 811
2 1649 1 819
2 1650 1 819
2 1651 1 819
2 1652 1 821
2 1653 1 821
2 1654 1 822
2 1655 1 822
2 1656 1 822
2 1657 1 822
2 1658 1 824
2 1659 1 824
2 1660 1 824
2 1661 1 825
2 1662 1 825
2 1663 1 826
2 1664 1 826
2 1665 1 837
2 1666 1 837
2 1667 1 839
2 1668 1 839
2 1669 1 843
2 1670 1 843
2 1671 1 850
2 1672 1 850
2 1673 1 850
2 1674 1 850
2 1675 1 851
2 1676 1 851
2 1677 1 851
2 1678 1 852
2 1679 1 852
2 1680 1 865
2 1681 1 865
2 1682 1 866
2 1683 1 866
2 1684 1 870
2 1685 1 870
2 1686 1 873
2 1687 1 873
2 1688 1 873
2 1689 1 875
2 1690 1 875
2 1691 1 876
2 1692 1 876
2 1693 1 876
2 1694 1 876
2 1695 1 883
2 1696 1 883
2 1697 1 883
2 1698 1 884
2 1699 1 884
2 1700 1 884
2 1701 1 885
2 1702 1 885
2 1703 1 898
2 1704 1 898
2 1705 1 899
2 1706 1 899
2 1707 1 903
2 1708 1 903
2 1709 1 906
2 1710 1 906
2 1711 1 906
2 1712 1 908
2 1713 1 908
2 1714 1 909
2 1715 1 909
2 1716 1 909
2 1717 1 909
2 1718 1 916
2 1719 1 916
2 1720 1 916
2 1721 1 918
2 1722 1 918
2 1723 1 932
2 1724 1 932
2 1725 1 936
2 1726 1 936
2 1727 1 938
2 1728 1 938
2 1729 1 939
2 1730 1 939
2 1731 1 941
2 1732 1 941
2 1733 1 942
2 1734 1 942
2 1735 1 942
2 1736 1 942
2 1737 1 949
2 1738 1 949
2 1739 1 949
2 1740 1 950
2 1741 1 950
2 1742 1 951
2 1743 1 951
2 1744 1 966
2 1745 1 966
2 1746 1 969
2 1747 1 969
2 1748 1 972
2 1749 1 972
2 1750 1 972
2 1751 1 974
2 1752 1 974
2 1753 1 974
2 1754 1 975
2 1755 1 975
2 1756 1 975
2 1757 1 975
2 1758 1 982
2 1759 1 982
2 1760 1 983
2 1761 1 983
2 1762 1 984
2 1763 1 984
2 1764 1 1000
2 1765 1 1000
2 1766 1 1003
2 1767 1 1003
2 1768 1 1005
2 1769 1 1005
2 1770 1 1006
2 1771 1 1006
2 1772 1 1006
2 1773 1 1014
2 1774 1 1014
0 97 5 1 1 64
0 98 5 1 1 66
0 99 5 1 1 68
0 100 5 1 1 70
0 101 5 1 1 72
0 102 5 1 1 74
0 103 5 1 1 76
0 104 5 1 1 78
0 105 5 1 1 80
0 106 5 1 1 82
0 107 5 1 1 84
0 108 5 1 1 86
0 109 5 1 1 88
0 110 5 1 1 90
0 111 5 1 1 92
0 112 5 1 1 94
0 113 5 1 1 96
0 114 5 1 1 176
0 115 5 1 1 208
0 116 5 1 1 251
0 117 5 1 1 299
0 118 5 1 1 349
0 119 5 1 1 399
0 120 5 1 1 455
0 121 5 1 1 512
0 122 5 1 1 572
0 123 5 1 1 632
0 124 5 1 1 692
0 125 5 1 1 752
0 126 5 1 1 817
0 127 5 1 1 882
0 128 5 1 1 948
0 129 5 1 1 1012
0 130 5 1 1 1034
0 131 5 1 1 1036
0 132 5 1 1 1038
0 133 5 1 1 1040
0 134 5 1 1 1042
0 135 5 1 1 1044
0 136 5 1 1 1046
0 137 5 1 1 1048
0 138 5 1 1 1050
0 139 5 1 1 1052
0 140 5 1 1 1054
0 141 5 1 1 1056
0 142 5 1 1 1058
0 143 5 1 1 1060
0 144 5 1 1 1062
0 145 5 1 1 1064
0 146 5 1 1 1066
0 147 5 1 1 1068
0 148 5 1 1 1070
0 149 5 1 1 1072
0 150 5 1 1 1074
0 151 5 1 1 1076
0 152 5 1 1 1078
0 153 5 1 1 1080
0 154 5 1 1 1082
0 155 5 1 1 1084
0 156 5 1 1 1086
0 157 5 1 1 1088
0 158 5 1 1 1090
0 159 5 1 1 1092
0 160 5 1 1 1094
0 161 7 2 2 65 1033
0 162 5 2 1 1096
0 163 7 1 2 97 129
0 164 5 1 1 163
3 2067 7 0 2 1098 164
0 166 7 1 2 67 1035
0 167 5 3 1 166
0 168 7 1 2 98 130
0 169 5 1 1 168
0 170 7 2 2 1100 169
0 171 5 1 1 1103
0 172 7 2 2 1097 1104
0 173 5 2 1 1105
0 174 7 1 2 1099 171
0 175 5 1 1 174
3 2068 7 0 2 1107 175
0 177 7 2 2 1101 1108
0 178 5 3 1 1109
0 179 7 1 2 69 1037
0 180 5 3 1 179
0 181 7 1 2 99 131
0 182 5 2 1 181
0 183 7 4 2 1114 1117
0 184 5 1 1 1119
0 185 7 1 2 1110 184
0 186 5 1 1 185
0 187 7 1 2 1111 1120
0 188 5 1 1 187
3 2069 7 0 2 186 188
0 190 7 2 2 1106 1121
0 191 5 1 1 1123
0 192 7 1 2 1102 1115
0 193 5 1 1 192
0 194 7 2 2 1118 193
0 195 5 1 1 1125
0 196 7 2 2 191 195
0 197 5 2 1 1127
0 198 7 1 2 71 1039
0 199 5 3 1 198
0 200 7 1 2 100 132
0 201 5 2 1 200
0 202 7 4 2 1131 1134
0 203 5 1 1 1136
0 204 7 1 2 1129 1137
0 205 5 1 1 204
0 206 7 1 2 1128 203
0 207 5 1 1 206
3 2070 7 0 2 205 207
0 209 7 2 2 1122 1138
0 210 7 1 2 1112 1140
0 211 5 1 1 210
0 212 7 1 2 1116 1132
0 213 5 1 1 212
0 214 7 2 2 1135 213
0 215 5 1 1 1142
0 216 7 2 2 211 215
0 217 5 2 1 1144
0 218 7 1 2 73 1041
0 219 5 3 1 218
0 220 7 1 2 101 133
0 221 5 2 1 220
0 222 7 4 2 1148 1151
0 223 5 1 1 1153
0 224 7 1 2 1146 1154
0 225 5 1 1 224
0 226 7 1 2 1145 223
0 227 5 1 1 226
3 2071 7 0 2 225 227
0 229 7 3 2 1139 1155
0 230 7 1 2 1124 1157
0 231 5 1 1 230
0 232 7 1 2 1126 1158
0 233 5 1 1 232
0 234 7 1 2 1133 1149
0 235 5 1 1 234
0 236 7 2 2 1152 235
0 237 5 1 1 1160
0 238 7 1 2 233 237
0 239 7 2 2 231 238
0 240 5 2 1 1162
0 241 7 1 2 75 1043
0 242 5 3 1 241
0 243 7 1 2 102 134
0 244 5 2 1 243
0 245 7 4 2 1166 1169
0 246 5 1 1 1171
0 247 7 1 2 1164 1172
0 248 5 1 1 247
0 249 7 1 2 1163 246
0 250 5 1 1 249
3 2072 7 0 2 248 250
0 252 7 3 2 1156 1173
0 253 7 1 2 1141 1175
0 254 7 1 2 1113 253
0 255 5 1 1 254
0 256 7 1 2 1143 1176
0 257 5 1 1 256
0 258 7 1 2 1150 1167
0 259 5 1 1 258
0 260 7 2 2 1170 259
0 261 5 1 1 1178
0 262 7 1 2 257 261
0 263 7 2 2 255 262
0 264 5 2 1 1180
0 265 7 1 2 77 1045
0 266 5 3 1 265
0 267 7 1 2 103 135
0 268 5 2 1 267
0 269 7 4 2 1184 1187
0 270 5 1 1 1189
0 271 7 1 2 1182 1190
0 272 5 1 1 271
0 273 7 1 2 1181 270
0 274 5 1 1 273
3 2073 7 0 2 272 274
0 276 7 3 2 1174 1191
0 277 7 1 2 1159 1193
0 278 7 1 2 1130 277
0 279 5 1 1 278
0 280 7 1 2 1161 1194
0 281 5 1 1 280
0 282 7 1 2 1168 1185
0 283 5 1 1 282
0 284 7 2 2 1188 283
0 285 5 1 1 1196
0 286 7 1 2 281 285
0 287 7 2 2 279 286
0 288 5 3 1 1198
0 289 7 1 2 79 1047
0 290 5 3 1 289
0 291 7 1 2 104 136
0 292 5 2 1 291
0 293 7 4 2 1203 1206
0 294 5 1 1 1208
0 295 7 1 2 1200 1209
0 296 5 1 1 295
0 297 7 1 2 1199 294
0 298 5 1 1 297
3 2074 7 0 2 296 298
0 300 7 3 2 1192 1210
0 301 7 1 2 1179 1212
0 302 5 1 1 301
0 303 7 1 2 1186 1204
0 304 5 1 1 303
0 305 7 2 2 1207 304
0 306 5 1 1 1215
0 307 7 2 2 302 306
0 308 5 1 1 1217
0 309 7 1 2 1177 1213
0 310 7 2 2 1147 309
0 311 5 1 1 1219
0 312 7 2 2 1218 311
0 313 5 2 1 1221
0 314 7 1 2 81 1049
0 315 5 3 1 314
0 316 7 1 2 105 137
0 317 5 2 1 316
0 318 7 4 2 1225 1228
0 319 5 1 1 1230
0 320 7 1 2 1223 1231
0 321 5 1 1 320
0 322 7 1 2 1222 319
0 323 5 1 1 322
3 2075 7 0 2 321 323
0 325 7 1 2 83 1051
0 326 5 3 1 325
0 327 7 1 2 106 138
0 328 5 2 1 327
0 329 7 4 2 1234 1237
0 330 5 1 1 1239
0 331 7 3 2 1211 1232
0 332 7 1 2 1197 1243
0 333 5 1 1 332
0 334 7 1 2 1205 1226
0 335 5 1 1 334
0 336 7 2 2 1229 335
0 337 5 1 1 1246
0 338 7 2 2 333 337
0 339 5 1 1 1248
0 340 7 1 2 1195 1244
0 341 7 2 2 1165 340
0 342 5 1 1 1250
0 343 7 2 2 1249 342
0 344 5 2 1 1252
0 345 7 1 2 1240 1254
0 346 5 1 1 345
0 347 7 1 2 330 1253
0 348 5 1 1 347
3 2076 7 0 2 346 348
0 350 7 1 2 85 1053
0 351 5 3 1 350
0 352 7 1 2 107 139
0 353 5 2 1 352
0 354 7 4 2 1256 1259
0 355 5 1 1 1261
0 356 7 3 2 1233 1241
0 357 7 1 2 1216 1265
0 358 5 1 1 357
0 359 7 1 2 1227 1235
0 360 5 1 1 359
0 361 7 2 2 1238 360
0 362 5 1 1 1268
0 363 7 2 2 358 362
0 364 5 1 1 1270
0 365 7 1 2 1214 1266
0 366 7 2 2 1183 365
0 367 5 1 1 1272
0 368 7 2 2 1271 367
0 369 5 2 1 1274
0 370 7 1 2 1262 1276
0 371 5 1 1 370
0 372 7 1 2 355 1275
0 373 5 1 1 372
3 2077 7 0 2 371 373
0 375 7 1 2 87 1055
0 376 5 3 1 375
0 377 7 1 2 108 140
0 378 5 2 1 377
0 379 7 4 2 1278 1281
0 380 5 1 1 1283
0 381 7 3 2 1242 1263
0 382 7 1 2 1247 1287
0 383 5 1 1 382
0 384 7 1 2 1236 1257
0 385 5 1 1 384
0 386 7 2 2 1260 385
0 387 5 1 1 1290
0 388 7 2 2 383 387
0 389 5 1 1 1292
0 390 7 2 2 1245 1288
0 391 7 1 2 1201 1294
0 392 5 1 1 391
0 393 7 2 2 1293 392
0 394 5 3 1 1296
0 395 7 1 2 1284 1298
0 396 5 1 1 395
0 397 7 1 2 380 1297
0 398 5 1 1 397
3 2078 7 0 2 396 398
0 400 7 3 2 1264 1285
0 401 7 3 2 1267 1301
0 402 7 1 2 1220 1304
0 403 5 1 1 402
0 404 7 1 2 1269 1302
0 405 5 1 1 404
0 406 7 1 2 1258 1279
0 407 5 1 1 406
0 408 7 2 2 1282 407
0 409 5 1 1 1307
0 410 7 2 2 405 409
0 411 5 1 1 1309
0 412 7 1 2 308 1305
0 413 5 1 1 412
0 414 7 1 2 1310 413
0 415 7 2 2 403 414
0 416 5 3 1 1311
0 417 7 1 2 89 1057
0 418 5 3 1 417
0 419 7 1 2 109 141
0 420 5 2 1 419
0 421 7 4 2 1316 1319
0 422 5 1 1 1321
0 423 7 1 2 1313 1322
0 424 5 1 1 423
0 425 7 1 2 1312 422
0 426 5 1 1 425
3 2079 7 0 2 424 426
0 428 7 3 2 1286 1323
0 429 7 3 2 1289 1325
0 430 7 1 2 1251 1328
0 431 5 1 1 430
0 432 7 1 2 1291 1326
0 433 5 1 1 432
0 434 7 1 2 1280 1317
0 435 5 1 1 434
0 436 7 2 2 1320 435
0 437 5 1 1 1331
0 438 7 2 2 433 437
0 439 5 1 1 1333
0 440 7 1 2 339 1329
0 441 5 1 1 440
0 442 7 1 2 1334 441
0 443 7 2 2 431 442
0 444 5 3 1 1335
0 445 7 1 2 91 1059
0 446 5 3 1 445
0 447 7 1 2 110 142
0 448 5 2 1 447
0 449 7 4 2 1340 1343
0 450 5 1 1 1345
0 451 7 1 2 1337 1346
0 452 5 1 1 451
0 453 7 1 2 1336 450
0 454 5 1 1 453
3 2080 7 0 2 452 454
0 456 7 3 2 1324 1347
0 457 7 3 2 1303 1349
0 458 7 1 2 1273 1352
0 459 5 1 1 458
0 460 7 1 2 1308 1350
0 461 5 1 1 460
0 462 7 1 2 1318 1341
0 463 5 1 1 462
0 464 7 2 2 1344 463
0 465 5 1 1 1355
0 466 7 2 2 461 465
0 467 5 1 1 1357
0 468 7 1 2 364 1353
0 469 5 1 1 468
0 470 7 1 2 1358 469
0 471 7 2 2 459 470
0 472 5 3 1 1359
0 473 7 1 2 93 1061
0 474 5 3 1 473
0 475 7 1 2 111 143
0 476 5 2 1 475
0 477 7 4 2 1364 1367
0 478 5 1 1 1369
0 479 7 1 2 1361 1370
0 480 5 1 1 479
0 481 7 1 2 1360 478
0 482 5 1 1 481
3 2081 7 0 2 480 482
0 484 7 3 2 1348 1371
0 485 7 3 2 1327 1373
0 486 7 1 2 1295 1376
0 487 7 1 2 1202 486
0 488 5 1 1 487
0 489 7 1 2 1332 1374
0 490 5 1 1 489
0 491 7 1 2 1342 1365
0 492 5 1 1 491
0 493 7 2 2 1368 492
0 494 5 1 1 1379
0 495 7 2 2 490 494
0 496 5 1 1 1381
0 497 7 1 2 389 1377
0 498 5 1 1 497
0 499 7 1 2 1382 498
0 500 7 2 2 488 499
0 501 5 3 1 1383
0 502 7 1 2 95 1063
0 503 5 3 1 502
0 504 7 1 2 112 144
0 505 5 2 1 504
0 506 7 4 2 1388 1391
0 507 5 1 1 1393
0 508 7 1 2 1385 1394
0 509 5 1 1 508
0 510 7 1 2 1384 507
0 511 5 1 1 510
3 2082 7 0 2 509 511
0 513 7 3 2 1372 1395
0 514 7 1 2 1356 1397
0 515 5 1 1 514
0 516 7 1 2 1366 1389
0 517 5 1 1 516
0 518 7 2 2 1392 517
0 519 5 1 1 1400
0 520 7 2 2 515 519
0 521 5 1 1 1402
0 522 7 3 2 1351 1398
0 523 7 1 2 411 1404
0 524 5 1 1 523
0 525 7 2 2 1403 524
0 526 5 1 1 1407
0 527 7 1 2 1306 1405
0 528 7 2 2 1224 527
0 529 5 1 1 1409
0 530 7 2 2 1408 529
0 531 5 2 1 1411
0 532 7 1 2 165 1065
0 533 5 3 1 532
0 534 7 1 2 113 145
0 535 5 2 1 534
0 536 7 4 2 1415 1418
0 537 5 1 1 1420
0 538 7 1 2 1413 1421
0 539 5 1 1 538
0 540 7 1 2 1412 537
0 541 5 1 1 540
3 2083 7 0 2 539 541
0 543 7 3 2 1396 1422
0 544 7 1 2 1380 1424
0 545 5 1 1 544
0 546 7 1 2 1390 1416
0 547 5 1 1 546
0 548 7 2 2 1419 547
0 549 5 1 1 1427
0 550 7 2 2 545 549
0 551 5 1 1 1429
0 552 7 3 2 1375 1425
0 553 7 1 2 439 1431
0 554 5 1 1 553
0 555 7 2 2 1430 554
0 556 5 1 1 1434
0 557 7 1 2 1330 1432
0 558 7 2 2 1255 557
0 559 5 1 1 1436
0 560 7 2 2 1435 559
0 561 5 1 1 1438
0 562 7 1 2 189 1067
0 563 5 3 1 562
0 564 7 1 2 114 146
0 565 5 2 1 564
0 566 7 4 2 1440 1443
0 567 5 1 1 1445
0 568 7 1 2 561 1446
0 569 5 1 1 568
0 570 7 1 2 1439 567
0 571 5 1 1 570
3 2084 7 0 2 569 571
0 573 7 3 2 1423 1447
0 574 7 1 2 1401 1449
0 575 5 1 1 574
0 576 7 1 2 1417 1441
0 577 5 1 1 576
0 578 7 2 2 1444 577
0 579 5 1 1 1452
0 580 7 2 2 575 579
0 581 5 1 1 1454
0 582 7 3 2 1399 1450
0 583 7 1 2 467 1456
0 584 5 1 1 583
0 585 7 2 2 1455 584
0 586 5 1 1 1459
0 587 7 1 2 1354 1457
0 588 7 2 2 1277 587
0 589 5 1 1 1461
0 590 7 2 2 1460 589
0 591 5 1 1 1463
0 592 7 1 2 228 1069
0 593 5 3 1 592
0 594 7 1 2 115 147
0 595 5 2 1 594
0 596 7 4 2 1465 1468
0 597 5 1 1 1470
0 598 7 1 2 591 1471
0 599 5 1 1 598
0 600 7 1 2 1464 597
0 601 5 1 1 600
3 2085 7 0 2 599 601
0 603 7 3 2 1448 1472
0 604 7 1 2 1428 1474
0 605 5 1 1 604
0 606 7 1 2 1442 1466
0 607 5 1 1 606
0 608 7 2 2 1469 607
0 609 5 1 1 1477
0 610 7 2 2 605 609
0 611 5 1 1 1479
0 612 7 3 2 1426 1475
0 613 7 1 2 496 1481
0 614 5 1 1 613
0 615 7 2 2 1480 614
0 616 5 1 1 1484
0 617 7 2 2 1378 1482
0 618 7 1 2 1299 1486
0 619 5 1 1 618
0 620 7 2 2 1485 619
0 621 5 1 1 1488
0 622 7 1 2 275 1071
0 623 5 3 1 622
0 624 7 1 2 116 148
0 625 5 2 1 624
0 626 7 4 2 1490 1493
0 627 5 1 1 1495
0 628 7 1 2 621 1496
0 629 5 1 1 628
0 630 7 1 2 1489 627
0 631 5 1 1 630
3 2086 7 0 2 629 631
0 633 7 3 2 1473 1497
0 634 7 1 2 1453 1499
0 635 5 1 1 634
0 636 7 1 2 1467 1491
0 637 5 1 1 636
0 638 7 2 2 1494 637
0 639 5 1 1 1502
0 640 7 2 2 635 639
0 641 5 1 1 1504
0 642 7 3 2 1451 1500
0 643 7 1 2 521 1506
0 644 5 1 1 643
0 645 7 2 2 1505 644
0 646 5 1 1 1509
0 647 7 2 2 1406 1507
0 648 7 1 2 1314 1511
0 649 5 1 1 648
0 650 7 2 2 1510 649
0 651 5 1 1 1513
0 652 7 1 2 324 1073
0 653 5 3 1 652
0 654 7 1 2 117 149
0 655 5 2 1 654
0 656 7 4 2 1515 1518
0 657 5 1 1 1520
0 658 7 1 2 651 1521
0 659 5 1 1 658
0 660 7 1 2 1514 657
0 661 5 1 1 660
3 2087 7 0 2 659 661
0 663 7 3 2 1498 1522
0 664 7 1 2 1478 1524
0 665 5 1 1 664
0 666 7 1 2 1492 1516
0 667 5 1 1 666
0 668 7 2 2 1519 667
0 669 5 1 1 1527
0 670 7 2 2 665 669
0 671 5 1 1 1529
0 672 7 3 2 1476 1525
0 673 7 1 2 551 1531
0 674 5 1 1 673
0 675 7 2 2 1530 674
0 676 5 1 1 1534
0 677 7 2 2 1433 1532
0 678 7 1 2 1338 1536
0 679 5 1 1 678
0 680 7 2 2 1535 679
0 681 5 1 1 1538
0 682 7 1 2 374 1075
0 683 5 3 1 682
0 684 7 1 2 118 150
0 685 5 2 1 684
0 686 7 4 2 1540 1543
0 687 5 1 1 1545
0 688 7 1 2 681 1546
0 689 5 1 1 688
0 690 7 1 2 1539 687
0 691 5 1 1 690
3 2088 7 0 2 689 691
0 693 7 3 2 1523 1547
0 694 7 1 2 1503 1549
0 695 5 1 1 694
0 696 7 1 2 1517 1541
0 697 5 1 1 696
0 698 7 2 2 1544 697
0 699 5 1 1 1552
0 700 7 2 2 695 699
0 701 5 1 1 1554
0 702 7 3 2 1501 1550
0 703 7 1 2 581 1556
0 704 5 1 1 703
0 705 7 2 2 1555 704
0 706 5 1 1 1559
0 707 7 2 2 1458 1557
0 708 7 1 2 1362 1561
0 709 5 1 1 708
0 710 7 2 2 1560 709
0 711 5 1 1 1563
0 712 7 1 2 427 1077
0 713 5 3 1 712
0 714 7 1 2 119 151
0 715 5 2 1 714
0 716 7 4 2 1565 1568
0 717 5 1 1 1570
0 718 7 1 2 711 1571
0 719 5 1 1 718
0 720 7 1 2 1564 717
0 721 5 1 1 720
3 2089 7 0 2 719 721
0 723 7 3 2 1548 1572
0 724 7 1 2 1528 1574
0 725 5 1 1 724
0 726 7 1 2 1542 1566
0 727 5 1 1 726
0 728 7 2 2 1569 727
0 729 5 1 1 1577
0 730 7 2 2 725 729
0 731 5 1 1 1579
0 732 7 3 2 1526 1575
0 733 7 1 2 611 1581
0 734 5 1 1 733
0 735 7 2 2 1580 734
0 736 5 1 1 1584
0 737 7 2 2 1483 1582
0 738 7 1 2 1386 1586
0 739 5 1 1 738
0 740 7 2 2 1585 739
0 741 5 1 1 1588
0 742 7 1 2 483 1079
0 743 5 3 1 742
0 744 7 1 2 120 152
0 745 5 2 1 744
0 746 7 4 2 1590 1593
0 747 5 1 1 1595
0 748 7 1 2 741 1596
0 749 5 1 1 748
0 750 7 1 2 1589 747
0 751 5 1 1 750
3 2090 7 0 2 749 751
0 753 7 4 2 1573 1597
0 754 7 3 2 1551 1599
0 755 7 3 2 1508 1603
0 756 7 1 2 1410 1606
0 757 5 1 1 756
0 758 7 1 2 1553 1600
0 759 5 1 1 758
0 760 7 1 2 1567 1591
0 761 5 1 1 760
0 762 7 2 2 1594 761
0 763 5 1 1 1609
0 764 7 2 2 759 763
0 765 5 1 1 1611
0 766 7 1 2 641 1604
0 767 5 1 1 766
0 768 7 2 2 1612 767
0 769 5 1 1 1613
0 770 7 1 2 526 1607
0 771 5 1 1 770
0 772 7 1 2 1614 771
0 773 7 2 2 757 772
0 774 5 1 1 1615
0 775 7 1 2 542 1081
0 776 5 3 1 775
0 777 7 1 2 121 153
0 778 5 2 1 777
0 779 7 4 2 1617 1620
0 780 5 1 1 1622
0 781 7 1 2 774 1623
0 782 5 1 1 781
0 783 7 1 2 1616 780
0 784 5 1 1 783
3 2091 7 0 2 782 784
0 786 7 1 2 602 1083
0 787 5 3 1 786
0 788 7 1 2 122 154
0 789 5 2 1 788
0 790 7 4 2 1626 1629
0 791 5 1 1 1631
0 792 7 3 2 1598 1624
0 793 7 3 2 1576 1635
0 794 7 2 2 1533 1638
0 795 7 1 2 1437 1641
0 796 5 1 1 795
0 797 7 1 2 556 1642
0 798 5 1 1 797
0 799 7 1 2 671 1639
0 800 5 1 1 799
0 801 7 1 2 1578 1636
0 802 5 1 1 801
0 803 7 1 2 1592 1618
0 804 5 1 1 803
0 805 7 2 2 1621 804
0 806 5 1 1 1643
0 807 7 2 2 802 806
0 808 5 1 1 1645
0 809 7 1 2 800 1646
0 810 7 1 2 798 809
0 811 7 2 2 796 810
0 812 5 1 1 1647
0 813 7 1 2 1632 812
0 814 5 1 1 813
0 815 7 1 2 791 1648
0 816 5 1 1 815
3 2092 7 0 2 814 816
0 818 7 1 2 662 1085
0 819 5 3 1 818
0 820 7 1 2 123 155
0 821 5 2 1 820
0 822 7 4 2 1649 1652
0 823 5 1 1 1654
0 824 7 3 2 1625 1633
0 825 7 2 2 1601 1658
0 826 7 2 2 1558 1661
0 827 7 1 2 1462 1663
0 828 5 1 1 827
0 829 7 1 2 586 1664
0 830 5 1 1 829
0 831 7 1 2 701 1662
0 832 5 1 1 831
0 833 7 1 2 1610 1659
0 834 5 1 1 833
0 835 7 1 2 1619 1627
0 836 5 1 1 835
0 837 7 2 2 1630 836
0 838 5 1 1 1665
0 839 7 2 2 834 838
0 840 5 1 1 1667
0 841 7 1 2 832 1668
0 842 7 1 2 830 841
0 843 7 2 2 828 842
0 844 5 1 1 1669
0 845 7 1 2 1655 844
0 846 5 1 1 845
0 847 7 1 2 823 1670
0 848 5 1 1 847
3 2093 7 0 2 846 848
0 850 7 4 2 1634 1656
0 851 7 3 2 1637 1671
0 852 7 2 2 1583 1675
0 853 7 1 2 1487 1678
0 854 7 1 2 1300 853
0 855 5 1 1 854
0 856 7 1 2 616 1679
0 857 5 1 1 856
0 858 7 1 2 731 1676
0 859 5 1 1 858
0 860 7 1 2 1644 1672
0 861 5 1 1 860
0 862 7 1 2 1628 1650
0 863 5 1 1 862
0 864 7 1 2 1653 863
0 865 5 2 1 864
0 866 7 2 2 861 1680
0 867 5 1 1 1682
0 868 7 1 2 859 1683
0 869 7 1 2 857 868
0 870 7 2 2 855 869
0 871 5 1 1 1684
0 872 7 1 2 722 1087
0 873 5 3 1 872
0 874 7 1 2 124 156
0 875 5 2 1 874
0 876 7 4 2 1686 1689
0 877 5 1 1 1691
0 878 7 1 2 871 1692
0 879 5 1 1 878
0 880 7 1 2 1685 877
0 881 5 1 1 880
3 2094 7 0 2 879 881
0 883 7 3 2 1657 1693
0 884 7 3 2 1660 1695
0 885 7 2 2 1605 1698
0 886 7 1 2 1512 1701
0 887 7 1 2 1315 886
0 888 5 1 1 887
0 889 7 1 2 646 1702
0 890 5 1 1 889
0 891 7 1 2 765 1699
0 892 5 1 1 891
0 893 7 1 2 1666 1696
0 894 5 1 1 893
0 895 7 1 2 1651 1687
0 896 5 1 1 895
0 897 7 1 2 1690 896
0 898 5 2 1 897
0 899 7 2 2 894 1703
0 900 5 1 1 1705
0 901 7 1 2 892 1706
0 902 7 1 2 890 901
0 903 7 2 2 888 902
0 904 5 1 1 1707
0 905 7 1 2 785 1089
0 906 5 3 1 905
0 907 7 1 2 125 157
0 908 5 2 1 907
0 909 7 4 2 1709 1712
0 910 5 1 1 1714
0 911 7 1 2 904 1715
0 912 5 1 1 911
0 913 7 1 2 1708 910
0 914 5 1 1 913
3 2095 7 0 2 912 914
0 916 7 3 2 1694 1716
0 917 7 1 2 1673 1718
0 918 7 2 2 1640 917
0 919 7 1 2 1537 1721
0 920 7 1 2 1339 919
0 921 5 1 1 920
0 922 7 1 2 676 1722
0 923 5 1 1 922
0 924 7 1 2 808 1674
0 925 5 1 1 924
0 926 7 1 2 1681 925
0 927 5 1 1 926
0 928 7 1 2 1719 927
0 929 5 1 1 928
0 930 7 1 2 1688 1710
0 931 5 1 1 930
0 932 7 2 2 1713 931
0 933 5 1 1 1723
0 934 7 1 2 929 933
0 935 7 1 2 923 934
0 936 7 2 2 921 935
0 937 5 1 1 1725
0 938 7 2 2 849 1091
0 939 5 2 1 1727
0 940 7 1 2 126 158
0 941 5 2 1 940
0 942 7 4 2 1729 1731
0 943 5 1 1 1733
0 944 7 1 2 937 1734
0 945 5 1 1 944
0 946 7 1 2 1726 943
0 947 5 1 1 946
3 2096 7 0 2 945 947
0 949 7 3 2 1717 1735
0 950 7 2 2 1700 1737
0 951 7 2 2 1602 1740
0 952 7 1 2 1562 1742
0 953 7 1 2 1363 952
0 954 5 1 1 953
0 955 7 1 2 706 1743
0 956 5 1 1 955
0 957 7 1 2 840 1697
0 958 5 1 1 957
0 959 7 1 2 1704 958
0 960 5 1 1 959
0 961 7 1 2 1738 960
0 962 5 1 1 961
0 963 7 1 2 1711 1730
0 964 5 1 1 963
0 965 7 1 2 1732 964
0 966 5 2 1 965
0 967 7 1 2 962 1744
0 968 7 1 2 956 967
0 969 7 2 2 954 968
0 970 5 1 1 1746
0 971 7 1 2 915 1093
0 972 5 3 1 971
0 973 7 1 2 127 159
0 974 5 3 1 973
0 975 7 4 2 1748 1751
0 976 5 1 1 1754
0 977 7 1 2 970 1755
0 978 5 1 1 977
0 979 7 1 2 1747 976
0 980 5 1 1 979
3 2097 7 0 2 978 980
0 982 7 2 2 1736 1756
0 983 7 2 2 1720 1758
0 984 7 2 2 1677 1760
0 985 7 1 2 1587 1762
0 986 7 1 2 1387 985
0 987 5 1 1 986
0 988 7 1 2 736 1763
0 989 5 1 1 988
0 990 7 1 2 867 1761
0 991 5 1 1 990
0 992 7 1 2 1724 1759
0 993 5 1 1 992
0 994 7 1 2 1728 1752
0 995 5 1 1 994
0 996 7 1 2 1749 995
0 997 7 1 2 993 996
0 998 7 1 2 991 997
0 999 7 1 2 989 998
0 1000 7 2 2 987 999
0 1001 5 1 1 1764
0 1002 7 1 2 981 1095
0 1003 5 2 1 1002
0 1004 7 1 2 128 160
0 1005 5 2 1 1004
0 1006 7 3 2 1766 1768
0 1007 5 1 1 1770
0 1008 7 1 2 1001 1771
0 1009 5 1 1 1008
0 1010 7 1 2 1765 1007
0 1011 5 1 1 1010
3 2098 7 0 2 1009 1011
0 1013 7 1 2 1757 1772
0 1014 7 2 2 1741 1013
0 1015 7 1 2 1608 1773
0 1016 7 1 2 1414 1015
0 1017 5 1 1 1016
0 1018 7 1 2 769 1774
0 1019 5 1 1 1018
0 1020 7 1 2 900 1739
0 1021 5 1 1 1020
0 1022 7 1 2 1745 1021
0 1023 5 1 1 1022
0 1024 7 1 2 1753 1023
0 1025 5 1 1 1024
0 1026 7 1 2 1750 1767
0 1027 7 1 2 1025 1026
0 1028 5 1 1 1027
0 1029 7 1 2 1769 1028
0 1030 5 1 1 1029
0 1031 7 1 2 1019 1030
0 1032 7 1 2 1017 1031
3 2099 5 0 1 1032
