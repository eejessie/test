1 0 0 208 0
2 25 1 0
2 26 1 0
2 39926 1 0
2 39927 1 0
2 39928 1 0
2 39929 1 0
2 39930 1 0
2 39931 1 0
2 39932 1 0
2 39933 1 0
2 39934 1 0
2 39935 1 0
2 39936 1 0
2 39937 1 0
2 39938 1 0
2 39939 1 0
2 39940 1 0
2 39941 1 0
2 39942 1 0
2 39943 1 0
2 39944 1 0
2 39945 1 0
2 39946 1 0
2 39947 1 0
2 39948 1 0
2 39949 1 0
2 39950 1 0
2 39951 1 0
2 39952 1 0
2 39953 1 0
2 39954 1 0
2 39955 1 0
2 39956 1 0
2 39957 1 0
2 39958 1 0
2 39959 1 0
2 39960 1 0
2 39961 1 0
2 39962 1 0
2 39963 1 0
2 39964 1 0
2 39965 1 0
2 39966 1 0
2 39967 1 0
2 39968 1 0
2 39969 1 0
2 39970 1 0
2 39971 1 0
2 39972 1 0
2 39973 1 0
2 39974 1 0
2 39975 1 0
2 39976 1 0
2 39977 1 0
2 39978 1 0
2 39979 1 0
2 39980 1 0
2 39981 1 0
2 39982 1 0
2 39983 1 0
2 39984 1 0
2 39985 1 0
2 39986 1 0
2 39987 1 0
2 39988 1 0
2 39989 1 0
2 39990 1 0
2 39991 1 0
2 39992 1 0
2 39993 1 0
2 39994 1 0
2 39995 1 0
2 39996 1 0
2 39997 1 0
2 39998 1 0
2 39999 1 0
2 40000 1 0
2 40001 1 0
2 40002 1 0
2 40003 1 0
2 40004 1 0
2 40005 1 0
2 40006 1 0
2 40007 1 0
2 40008 1 0
2 40009 1 0
2 40010 1 0
2 40011 1 0
2 40012 1 0
2 40013 1 0
2 40014 1 0
2 40015 1 0
2 40016 1 0
2 40017 1 0
2 40018 1 0
2 40019 1 0
2 40020 1 0
2 40021 1 0
2 40022 1 0
2 40023 1 0
2 40024 1 0
2 40025 1 0
2 40026 1 0
2 40027 1 0
2 40028 1 0
2 40029 1 0
2 40030 1 0
2 40031 1 0
2 40032 1 0
2 40033 1 0
2 40034 1 0
2 40035 1 0
2 40036 1 0
2 40037 1 0
2 40038 1 0
2 40039 1 0
2 40040 1 0
2 40041 1 0
2 40042 1 0
2 40043 1 0
2 40044 1 0
2 40045 1 0
2 40046 1 0
2 40047 1 0
2 40048 1 0
2 40049 1 0
2 40050 1 0
2 40051 1 0
2 40052 1 0
2 40053 1 0
2 40054 1 0
2 40055 1 0
2 40056 1 0
2 40057 1 0
2 40058 1 0
2 40059 1 0
2 40060 1 0
2 40061 1 0
2 40062 1 0
2 40063 1 0
2 40064 1 0
2 40065 1 0
2 40066 1 0
2 40067 1 0
2 40068 1 0
2 40069 1 0
2 40070 1 0
2 40071 1 0
2 40072 1 0
2 40073 1 0
2 40074 1 0
2 40075 1 0
2 40076 1 0
2 40077 1 0
2 40078 1 0
2 40079 1 0
2 40080 1 0
2 40081 1 0
2 40082 1 0
2 40083 1 0
2 40084 1 0
2 40085 1 0
2 40086 1 0
2 40087 1 0
2 40088 1 0
2 40089 1 0
2 40090 1 0
2 40091 1 0
2 40092 1 0
2 40093 1 0
2 40094 1 0
2 40095 1 0
2 40096 1 0
2 40097 1 0
2 40098 1 0
2 40099 1 0
2 40100 1 0
2 40101 1 0
2 40102 1 0
2 40103 1 0
2 40104 1 0
2 40105 1 0
2 40106 1 0
2 40107 1 0
2 40108 1 0
2 40109 1 0
2 40110 1 0
2 40111 1 0
2 40112 1 0
2 40113 1 0
2 40114 1 0
2 40115 1 0
2 40116 1 0
2 40117 1 0
2 40118 1 0
2 40119 1 0
2 40120 1 0
2 40121 1 0
2 40122 1 0
2 40123 1 0
2 40124 1 0
2 40125 1 0
2 40126 1 0
2 40127 1 0
2 40128 1 0
2 40129 1 0
2 40130 1 0
2 40131 1 0
1 1 0 177 0
2 40132 1 1
2 40133 1 1
2 40134 1 1
2 40135 1 1
2 40136 1 1
2 40137 1 1
2 40138 1 1
2 40139 1 1
2 40140 1 1
2 40141 1 1
2 40142 1 1
2 40143 1 1
2 40144 1 1
2 40145 1 1
2 40146 1 1
2 40147 1 1
2 40148 1 1
2 40149 1 1
2 40150 1 1
2 40151 1 1
2 40152 1 1
2 40153 1 1
2 40154 1 1
2 40155 1 1
2 40156 1 1
2 40157 1 1
2 40158 1 1
2 40159 1 1
2 40160 1 1
2 40161 1 1
2 40162 1 1
2 40163 1 1
2 40164 1 1
2 40165 1 1
2 40166 1 1
2 40167 1 1
2 40168 1 1
2 40169 1 1
2 40170 1 1
2 40171 1 1
2 40172 1 1
2 40173 1 1
2 40174 1 1
2 40175 1 1
2 40176 1 1
2 40177 1 1
2 40178 1 1
2 40179 1 1
2 40180 1 1
2 40181 1 1
2 40182 1 1
2 40183 1 1
2 40184 1 1
2 40185 1 1
2 40186 1 1
2 40187 1 1
2 40188 1 1
2 40189 1 1
2 40190 1 1
2 40191 1 1
2 40192 1 1
2 40193 1 1
2 40194 1 1
2 40195 1 1
2 40196 1 1
2 40197 1 1
2 40198 1 1
2 40199 1 1
2 40200 1 1
2 40201 1 1
2 40202 1 1
2 40203 1 1
2 40204 1 1
2 40205 1 1
2 40206 1 1
2 40207 1 1
2 40208 1 1
2 40209 1 1
2 40210 1 1
2 40211 1 1
2 40212 1 1
2 40213 1 1
2 40214 1 1
2 40215 1 1
2 40216 1 1
2 40217 1 1
2 40218 1 1
2 40219 1 1
2 40220 1 1
2 40221 1 1
2 40222 1 1
2 40223 1 1
2 40224 1 1
2 40225 1 1
2 40226 1 1
2 40227 1 1
2 40228 1 1
2 40229 1 1
2 40230 1 1
2 40231 1 1
2 40232 1 1
2 40233 1 1
2 40234 1 1
2 40235 1 1
2 40236 1 1
2 40237 1 1
2 40238 1 1
2 40239 1 1
2 40240 1 1
2 40241 1 1
2 40242 1 1
2 40243 1 1
2 40244 1 1
2 40245 1 1
2 40246 1 1
2 40247 1 1
2 40248 1 1
2 40249 1 1
2 40250 1 1
2 40251 1 1
2 40252 1 1
2 40253 1 1
2 40254 1 1
2 40255 1 1
2 40256 1 1
2 40257 1 1
2 40258 1 1
2 40259 1 1
2 40260 1 1
2 40261 1 1
2 40262 1 1
2 40263 1 1
2 40264 1 1
2 40265 1 1
2 40266 1 1
2 40267 1 1
2 40268 1 1
2 40269 1 1
2 40270 1 1
2 40271 1 1
2 40272 1 1
2 40273 1 1
2 40274 1 1
2 40275 1 1
2 40276 1 1
2 40277 1 1
2 40278 1 1
2 40279 1 1
2 40280 1 1
2 40281 1 1
2 40282 1 1
2 40283 1 1
2 40284 1 1
2 40285 1 1
2 40286 1 1
2 40287 1 1
2 40288 1 1
2 40289 1 1
2 40290 1 1
2 40291 1 1
2 40292 1 1
2 40293 1 1
2 40294 1 1
2 40295 1 1
2 40296 1 1
2 40297 1 1
2 40298 1 1
2 40299 1 1
2 40300 1 1
2 40301 1 1
2 40302 1 1
2 40303 1 1
2 40304 1 1
2 40305 1 1
2 40306 1 1
2 40307 1 1
2 40308 1 1
1 2 0 233 0
2 40309 1 2
2 40310 1 2
2 40311 1 2
2 40312 1 2
2 40313 1 2
2 40314 1 2
2 40315 1 2
2 40316 1 2
2 40317 1 2
2 40318 1 2
2 40319 1 2
2 40320 1 2
2 40321 1 2
2 40322 1 2
2 40323 1 2
2 40324 1 2
2 40325 1 2
2 40326 1 2
2 40327 1 2
2 40328 1 2
2 40329 1 2
2 40330 1 2
2 40331 1 2
2 40332 1 2
2 40333 1 2
2 40334 1 2
2 40335 1 2
2 40336 1 2
2 40337 1 2
2 40338 1 2
2 40339 1 2
2 40340 1 2
2 40341 1 2
2 40342 1 2
2 40343 1 2
2 40344 1 2
2 40345 1 2
2 40346 1 2
2 40347 1 2
2 40348 1 2
2 40349 1 2
2 40350 1 2
2 40351 1 2
2 40352 1 2
2 40353 1 2
2 40354 1 2
2 40355 1 2
2 40356 1 2
2 40357 1 2
2 40358 1 2
2 40359 1 2
2 40360 1 2
2 40361 1 2
2 40362 1 2
2 40363 1 2
2 40364 1 2
2 40365 1 2
2 40366 1 2
2 40367 1 2
2 40368 1 2
2 40369 1 2
2 40370 1 2
2 40371 1 2
2 40372 1 2
2 40373 1 2
2 40374 1 2
2 40375 1 2
2 40376 1 2
2 40377 1 2
2 40378 1 2
2 40379 1 2
2 40380 1 2
2 40381 1 2
2 40382 1 2
2 40383 1 2
2 40384 1 2
2 40385 1 2
2 40386 1 2
2 40387 1 2
2 40388 1 2
2 40389 1 2
2 40390 1 2
2 40391 1 2
2 40392 1 2
2 40393 1 2
2 40394 1 2
2 40395 1 2
2 40396 1 2
2 40397 1 2
2 40398 1 2
2 40399 1 2
2 40400 1 2
2 40401 1 2
2 40402 1 2
2 40403 1 2
2 40404 1 2
2 40405 1 2
2 40406 1 2
2 40407 1 2
2 40408 1 2
2 40409 1 2
2 40410 1 2
2 40411 1 2
2 40412 1 2
2 40413 1 2
2 40414 1 2
2 40415 1 2
2 40416 1 2
2 40417 1 2
2 40418 1 2
2 40419 1 2
2 40420 1 2
2 40421 1 2
2 40422 1 2
2 40423 1 2
2 40424 1 2
2 40425 1 2
2 40426 1 2
2 40427 1 2
2 40428 1 2
2 40429 1 2
2 40430 1 2
2 40431 1 2
2 40432 1 2
2 40433 1 2
2 40434 1 2
2 40435 1 2
2 40436 1 2
2 40437 1 2
2 40438 1 2
2 40439 1 2
2 40440 1 2
2 40441 1 2
2 40442 1 2
2 40443 1 2
2 40444 1 2
2 40445 1 2
2 40446 1 2
2 40447 1 2
2 40448 1 2
2 40449 1 2
2 40450 1 2
2 40451 1 2
2 40452 1 2
2 40453 1 2
2 40454 1 2
2 40455 1 2
2 40456 1 2
2 40457 1 2
2 40458 1 2
2 40459 1 2
2 40460 1 2
2 40461 1 2
2 40462 1 2
2 40463 1 2
2 40464 1 2
2 40465 1 2
2 40466 1 2
2 40467 1 2
2 40468 1 2
2 40469 1 2
2 40470 1 2
2 40471 1 2
2 40472 1 2
2 40473 1 2
2 40474 1 2
2 40475 1 2
2 40476 1 2
2 40477 1 2
2 40478 1 2
2 40479 1 2
2 40480 1 2
2 40481 1 2
2 40482 1 2
2 40483 1 2
2 40484 1 2
2 40485 1 2
2 40486 1 2
2 40487 1 2
2 40488 1 2
2 40489 1 2
2 40490 1 2
2 40491 1 2
2 40492 1 2
2 40493 1 2
2 40494 1 2
2 40495 1 2
2 40496 1 2
2 40497 1 2
2 40498 1 2
2 40499 1 2
2 40500 1 2
2 40501 1 2
2 40502 1 2
2 40503 1 2
2 40504 1 2
2 40505 1 2
2 40506 1 2
2 40507 1 2
2 40508 1 2
2 40509 1 2
2 40510 1 2
2 40511 1 2
2 40512 1 2
2 40513 1 2
2 40514 1 2
2 40515 1 2
2 40516 1 2
2 40517 1 2
2 40518 1 2
2 40519 1 2
2 40520 1 2
2 40521 1 2
2 40522 1 2
2 40523 1 2
2 40524 1 2
2 40525 1 2
2 40526 1 2
2 40527 1 2
2 40528 1 2
2 40529 1 2
2 40530 1 2
2 40531 1 2
2 40532 1 2
2 40533 1 2
2 40534 1 2
2 40535 1 2
2 40536 1 2
2 40537 1 2
2 40538 1 2
2 40539 1 2
2 40540 1 2
2 40541 1 2
1 3 0 163 0
2 40542 1 3
2 40543 1 3
2 40544 1 3
2 40545 1 3
2 40546 1 3
2 40547 1 3
2 40548 1 3
2 40549 1 3
2 40550 1 3
2 40551 1 3
2 40552 1 3
2 40553 1 3
2 40554 1 3
2 40555 1 3
2 40556 1 3
2 40557 1 3
2 40558 1 3
2 40559 1 3
2 40560 1 3
2 40561 1 3
2 40562 1 3
2 40563 1 3
2 40564 1 3
2 40565 1 3
2 40566 1 3
2 40567 1 3
2 40568 1 3
2 40569 1 3
2 40570 1 3
2 40571 1 3
2 40572 1 3
2 40573 1 3
2 40574 1 3
2 40575 1 3
2 40576 1 3
2 40577 1 3
2 40578 1 3
2 40579 1 3
2 40580 1 3
2 40581 1 3
2 40582 1 3
2 40583 1 3
2 40584 1 3
2 40585 1 3
2 40586 1 3
2 40587 1 3
2 40588 1 3
2 40589 1 3
2 40590 1 3
2 40591 1 3
2 40592 1 3
2 40593 1 3
2 40594 1 3
2 40595 1 3
2 40596 1 3
2 40597 1 3
2 40598 1 3
2 40599 1 3
2 40600 1 3
2 40601 1 3
2 40602 1 3
2 40603 1 3
2 40604 1 3
2 40605 1 3
2 40606 1 3
2 40607 1 3
2 40608 1 3
2 40609 1 3
2 40610 1 3
2 40611 1 3
2 40612 1 3
2 40613 1 3
2 40614 1 3
2 40615 1 3
2 40616 1 3
2 40617 1 3
2 40618 1 3
2 40619 1 3
2 40620 1 3
2 40621 1 3
2 40622 1 3
2 40623 1 3
2 40624 1 3
2 40625 1 3
2 40626 1 3
2 40627 1 3
2 40628 1 3
2 40629 1 3
2 40630 1 3
2 40631 1 3
2 40632 1 3
2 40633 1 3
2 40634 1 3
2 40635 1 3
2 40636 1 3
2 40637 1 3
2 40638 1 3
2 40639 1 3
2 40640 1 3
2 40641 1 3
2 40642 1 3
2 40643 1 3
2 40644 1 3
2 40645 1 3
2 40646 1 3
2 40647 1 3
2 40648 1 3
2 40649 1 3
2 40650 1 3
2 40651 1 3
2 40652 1 3
2 40653 1 3
2 40654 1 3
2 40655 1 3
2 40656 1 3
2 40657 1 3
2 40658 1 3
2 40659 1 3
2 40660 1 3
2 40661 1 3
2 40662 1 3
2 40663 1 3
2 40664 1 3
2 40665 1 3
2 40666 1 3
2 40667 1 3
2 40668 1 3
2 40669 1 3
2 40670 1 3
2 40671 1 3
2 40672 1 3
2 40673 1 3
2 40674 1 3
2 40675 1 3
2 40676 1 3
2 40677 1 3
2 40678 1 3
2 40679 1 3
2 40680 1 3
2 40681 1 3
2 40682 1 3
2 40683 1 3
2 40684 1 3
2 40685 1 3
2 40686 1 3
2 40687 1 3
2 40688 1 3
2 40689 1 3
2 40690 1 3
2 40691 1 3
2 40692 1 3
2 40693 1 3
2 40694 1 3
2 40695 1 3
2 40696 1 3
2 40697 1 3
2 40698 1 3
2 40699 1 3
2 40700 1 3
2 40701 1 3
2 40702 1 3
2 40703 1 3
2 40704 1 3
1 4 0 195 0
2 40705 1 4
2 40706 1 4
2 40707 1 4
2 40708 1 4
2 40709 1 4
2 40710 1 4
2 40711 1 4
2 40712 1 4
2 40713 1 4
2 40714 1 4
2 40715 1 4
2 40716 1 4
2 40717 1 4
2 40718 1 4
2 40719 1 4
2 40720 1 4
2 40721 1 4
2 40722 1 4
2 40723 1 4
2 40724 1 4
2 40725 1 4
2 40726 1 4
2 40727 1 4
2 40728 1 4
2 40729 1 4
2 40730 1 4
2 40731 1 4
2 40732 1 4
2 40733 1 4
2 40734 1 4
2 40735 1 4
2 40736 1 4
2 40737 1 4
2 40738 1 4
2 40739 1 4
2 40740 1 4
2 40741 1 4
2 40742 1 4
2 40743 1 4
2 40744 1 4
2 40745 1 4
2 40746 1 4
2 40747 1 4
2 40748 1 4
2 40749 1 4
2 40750 1 4
2 40751 1 4
2 40752 1 4
2 40753 1 4
2 40754 1 4
2 40755 1 4
2 40756 1 4
2 40757 1 4
2 40758 1 4
2 40759 1 4
2 40760 1 4
2 40761 1 4
2 40762 1 4
2 40763 1 4
2 40764 1 4
2 40765 1 4
2 40766 1 4
2 40767 1 4
2 40768 1 4
2 40769 1 4
2 40770 1 4
2 40771 1 4
2 40772 1 4
2 40773 1 4
2 40774 1 4
2 40775 1 4
2 40776 1 4
2 40777 1 4
2 40778 1 4
2 40779 1 4
2 40780 1 4
2 40781 1 4
2 40782 1 4
2 40783 1 4
2 40784 1 4
2 40785 1 4
2 40786 1 4
2 40787 1 4
2 40788 1 4
2 40789 1 4
2 40790 1 4
2 40791 1 4
2 40792 1 4
2 40793 1 4
2 40794 1 4
2 40795 1 4
2 40796 1 4
2 40797 1 4
2 40798 1 4
2 40799 1 4
2 40800 1 4
2 40801 1 4
2 40802 1 4
2 40803 1 4
2 40804 1 4
2 40805 1 4
2 40806 1 4
2 40807 1 4
2 40808 1 4
2 40809 1 4
2 40810 1 4
2 40811 1 4
2 40812 1 4
2 40813 1 4
2 40814 1 4
2 40815 1 4
2 40816 1 4
2 40817 1 4
2 40818 1 4
2 40819 1 4
2 40820 1 4
2 40821 1 4
2 40822 1 4
2 40823 1 4
2 40824 1 4
2 40825 1 4
2 40826 1 4
2 40827 1 4
2 40828 1 4
2 40829 1 4
2 40830 1 4
2 40831 1 4
2 40832 1 4
2 40833 1 4
2 40834 1 4
2 40835 1 4
2 40836 1 4
2 40837 1 4
2 40838 1 4
2 40839 1 4
2 40840 1 4
2 40841 1 4
2 40842 1 4
2 40843 1 4
2 40844 1 4
2 40845 1 4
2 40846 1 4
2 40847 1 4
2 40848 1 4
2 40849 1 4
2 40850 1 4
2 40851 1 4
2 40852 1 4
2 40853 1 4
2 40854 1 4
2 40855 1 4
2 40856 1 4
2 40857 1 4
2 40858 1 4
2 40859 1 4
2 40860 1 4
2 40861 1 4
2 40862 1 4
2 40863 1 4
2 40864 1 4
2 40865 1 4
2 40866 1 4
2 40867 1 4
2 40868 1 4
2 40869 1 4
2 40870 1 4
2 40871 1 4
2 40872 1 4
2 40873 1 4
2 40874 1 4
2 40875 1 4
2 40876 1 4
2 40877 1 4
2 40878 1 4
2 40879 1 4
2 40880 1 4
2 40881 1 4
2 40882 1 4
2 40883 1 4
2 40884 1 4
2 40885 1 4
2 40886 1 4
2 40887 1 4
2 40888 1 4
2 40889 1 4
2 40890 1 4
2 40891 1 4
2 40892 1 4
2 40893 1 4
2 40894 1 4
2 40895 1 4
2 40896 1 4
2 40897 1 4
2 40898 1 4
2 40899 1 4
1 5 0 71 0
2 40900 1 5
2 40901 1 5
2 40902 1 5
2 40903 1 5
2 40904 1 5
2 40905 1 5
2 40906 1 5
2 40907 1 5
2 40908 1 5
2 40909 1 5
2 40910 1 5
2 40911 1 5
2 40912 1 5
2 40913 1 5
2 40914 1 5
2 40915 1 5
2 40916 1 5
2 40917 1 5
2 40918 1 5
2 40919 1 5
2 40920 1 5
2 40921 1 5
2 40922 1 5
2 40923 1 5
2 40924 1 5
2 40925 1 5
2 40926 1 5
2 40927 1 5
2 40928 1 5
2 40929 1 5
2 40930 1 5
2 40931 1 5
2 40932 1 5
2 40933 1 5
2 40934 1 5
2 40935 1 5
2 40936 1 5
2 40937 1 5
2 40938 1 5
2 40939 1 5
2 40940 1 5
2 40941 1 5
2 40942 1 5
2 40943 1 5
2 40944 1 5
2 40945 1 5
2 40946 1 5
2 40947 1 5
2 40948 1 5
2 40949 1 5
2 40950 1 5
2 40951 1 5
2 40952 1 5
2 40953 1 5
2 40954 1 5
2 40955 1 5
2 40956 1 5
2 40957 1 5
2 40958 1 5
2 40959 1 5
2 40960 1 5
2 40961 1 5
2 40962 1 5
2 40963 1 5
2 40964 1 5
2 40965 1 5
2 40966 1 5
2 40967 1 5
2 40968 1 5
2 40969 1 5
2 40970 1 5
1 6 0 67 0
2 40971 1 6
2 40972 1 6
2 40973 1 6
2 40974 1 6
2 40975 1 6
2 40976 1 6
2 40977 1 6
2 40978 1 6
2 40979 1 6
2 40980 1 6
2 40981 1 6
2 40982 1 6
2 40983 1 6
2 40984 1 6
2 40985 1 6
2 40986 1 6
2 40987 1 6
2 40988 1 6
2 40989 1 6
2 40990 1 6
2 40991 1 6
2 40992 1 6
2 40993 1 6
2 40994 1 6
2 40995 1 6
2 40996 1 6
2 40997 1 6
2 40998 1 6
2 40999 1 6
2 41000 1 6
2 41001 1 6
2 41002 1 6
2 41003 1 6
2 41004 1 6
2 41005 1 6
2 41006 1 6
2 41007 1 6
2 41008 1 6
2 41009 1 6
2 41010 1 6
2 41011 1 6
2 41012 1 6
2 41013 1 6
2 41014 1 6
2 41015 1 6
2 41016 1 6
2 41017 1 6
2 41018 1 6
2 41019 1 6
2 41020 1 6
2 41021 1 6
2 41022 1 6
2 41023 1 6
2 41024 1 6
2 41025 1 6
2 41026 1 6
2 41027 1 6
2 41028 1 6
2 41029 1 6
2 41030 1 6
2 41031 1 6
2 41032 1 6
2 41033 1 6
2 41034 1 6
2 41035 1 6
2 41036 1 6
2 41037 1 6
1 7 0 17 0
2 41038 1 7
2 41039 1 7
2 41040 1 7
2 41041 1 7
2 41042 1 7
2 41043 1 7
2 41044 1 7
2 41045 1 7
2 41046 1 7
2 41047 1 7
2 41048 1 7
2 41049 1 7
2 41050 1 7
2 41051 1 7
2 41052 1 7
2 41053 1 7
2 41054 1 7
1 8 0 102 0
2 41055 1 8
2 41056 1 8
2 41057 1 8
2 41058 1 8
2 41059 1 8
2 41060 1 8
2 41061 1 8
2 41062 1 8
2 41063 1 8
2 41064 1 8
2 41065 1 8
2 41066 1 8
2 41067 1 8
2 41068 1 8
2 41069 1 8
2 41070 1 8
2 41071 1 8
2 41072 1 8
2 41073 1 8
2 41074 1 8
2 41075 1 8
2 41076 1 8
2 41077 1 8
2 41078 1 8
2 41079 1 8
2 41080 1 8
2 41081 1 8
2 41082 1 8
2 41083 1 8
2 41084 1 8
2 41085 1 8
2 41086 1 8
2 41087 1 8
2 41088 1 8
2 41089 1 8
2 41090 1 8
2 41091 1 8
2 41092 1 8
2 41093 1 8
2 41094 1 8
2 41095 1 8
2 41096 1 8
2 41097 1 8
2 41098 1 8
2 41099 1 8
2 41100 1 8
2 41101 1 8
2 41102 1 8
2 41103 1 8
2 41104 1 8
2 41105 1 8
2 41106 1 8
2 41107 1 8
2 41108 1 8
2 41109 1 8
2 41110 1 8
2 41111 1 8
2 41112 1 8
2 41113 1 8
2 41114 1 8
2 41115 1 8
2 41116 1 8
2 41117 1 8
2 41118 1 8
2 41119 1 8
2 41120 1 8
2 41121 1 8
2 41122 1 8
2 41123 1 8
2 41124 1 8
2 41125 1 8
2 41126 1 8
2 41127 1 8
2 41128 1 8
2 41129 1 8
2 41130 1 8
2 41131 1 8
2 41132 1 8
2 41133 1 8
2 41134 1 8
2 41135 1 8
2 41136 1 8
2 41137 1 8
2 41138 1 8
2 41139 1 8
2 41140 1 8
2 41141 1 8
2 41142 1 8
2 41143 1 8
2 41144 1 8
2 41145 1 8
2 41146 1 8
2 41147 1 8
2 41148 1 8
2 41149 1 8
2 41150 1 8
2 41151 1 8
2 41152 1 8
2 41153 1 8
2 41154 1 8
2 41155 1 8
2 41156 1 8
1 9 0 128 0
2 41157 1 9
2 41158 1 9
2 41159 1 9
2 41160 1 9
2 41161 1 9
2 41162 1 9
2 41163 1 9
2 41164 1 9
2 41165 1 9
2 41166 1 9
2 41167 1 9
2 41168 1 9
2 41169 1 9
2 41170 1 9
2 41171 1 9
2 41172 1 9
2 41173 1 9
2 41174 1 9
2 41175 1 9
2 41176 1 9
2 41177 1 9
2 41178 1 9
2 41179 1 9
2 41180 1 9
2 41181 1 9
2 41182 1 9
2 41183 1 9
2 41184 1 9
2 41185 1 9
2 41186 1 9
2 41187 1 9
2 41188 1 9
2 41189 1 9
2 41190 1 9
2 41191 1 9
2 41192 1 9
2 41193 1 9
2 41194 1 9
2 41195 1 9
2 41196 1 9
2 41197 1 9
2 41198 1 9
2 41199 1 9
2 41200 1 9
2 41201 1 9
2 41202 1 9
2 41203 1 9
2 41204 1 9
2 41205 1 9
2 41206 1 9
2 41207 1 9
2 41208 1 9
2 41209 1 9
2 41210 1 9
2 41211 1 9
2 41212 1 9
2 41213 1 9
2 41214 1 9
2 41215 1 9
2 41216 1 9
2 41217 1 9
2 41218 1 9
2 41219 1 9
2 41220 1 9
2 41221 1 9
2 41222 1 9
2 41223 1 9
2 41224 1 9
2 41225 1 9
2 41226 1 9
2 41227 1 9
2 41228 1 9
2 41229 1 9
2 41230 1 9
2 41231 1 9
2 41232 1 9
2 41233 1 9
2 41234 1 9
2 41235 1 9
2 41236 1 9
2 41237 1 9
2 41238 1 9
2 41239 1 9
2 41240 1 9
2 41241 1 9
2 41242 1 9
2 41243 1 9
2 41244 1 9
2 41245 1 9
2 41246 1 9
2 41247 1 9
2 41248 1 9
2 41249 1 9
2 41250 1 9
2 41251 1 9
2 41252 1 9
2 41253 1 9
2 41254 1 9
2 41255 1 9
2 41256 1 9
2 41257 1 9
2 41258 1 9
2 41259 1 9
2 41260 1 9
2 41261 1 9
2 41262 1 9
2 41263 1 9
2 41264 1 9
2 41265 1 9
2 41266 1 9
2 41267 1 9
2 41268 1 9
2 41269 1 9
2 41270 1 9
2 41271 1 9
2 41272 1 9
2 41273 1 9
2 41274 1 9
2 41275 1 9
2 41276 1 9
2 41277 1 9
2 41278 1 9
2 41279 1 9
2 41280 1 9
2 41281 1 9
2 41282 1 9
2 41283 1 9
2 41284 1 9
1 10 0 124 0
2 41285 1 10
2 41286 1 10
2 41287 1 10
2 41288 1 10
2 41289 1 10
2 41290 1 10
2 41291 1 10
2 41292 1 10
2 41293 1 10
2 41294 1 10
2 41295 1 10
2 41296 1 10
2 41297 1 10
2 41298 1 10
2 41299 1 10
2 41300 1 10
2 41301 1 10
2 41302 1 10
2 41303 1 10
2 41304 1 10
2 41305 1 10
2 41306 1 10
2 41307 1 10
2 41308 1 10
2 41309 1 10
2 41310 1 10
2 41311 1 10
2 41312 1 10
2 41313 1 10
2 41314 1 10
2 41315 1 10
2 41316 1 10
2 41317 1 10
2 41318 1 10
2 41319 1 10
2 41320 1 10
2 41321 1 10
2 41322 1 10
2 41323 1 10
2 41324 1 10
2 41325 1 10
2 41326 1 10
2 41327 1 10
2 41328 1 10
2 41329 1 10
2 41330 1 10
2 41331 1 10
2 41332 1 10
2 41333 1 10
2 41334 1 10
2 41335 1 10
2 41336 1 10
2 41337 1 10
2 41338 1 10
2 41339 1 10
2 41340 1 10
2 41341 1 10
2 41342 1 10
2 41343 1 10
2 41344 1 10
2 41345 1 10
2 41346 1 10
2 41347 1 10
2 41348 1 10
2 41349 1 10
2 41350 1 10
2 41351 1 10
2 41352 1 10
2 41353 1 10
2 41354 1 10
2 41355 1 10
2 41356 1 10
2 41357 1 10
2 41358 1 10
2 41359 1 10
2 41360 1 10
2 41361 1 10
2 41362 1 10
2 41363 1 10
2 41364 1 10
2 41365 1 10
2 41366 1 10
2 41367 1 10
2 41368 1 10
2 41369 1 10
2 41370 1 10
2 41371 1 10
2 41372 1 10
2 41373 1 10
2 41374 1 10
2 41375 1 10
2 41376 1 10
2 41377 1 10
2 41378 1 10
2 41379 1 10
2 41380 1 10
2 41381 1 10
2 41382 1 10
2 41383 1 10
2 41384 1 10
2 41385 1 10
2 41386 1 10
2 41387 1 10
2 41388 1 10
2 41389 1 10
2 41390 1 10
2 41391 1 10
2 41392 1 10
2 41393 1 10
2 41394 1 10
2 41395 1 10
2 41396 1 10
2 41397 1 10
2 41398 1 10
2 41399 1 10
2 41400 1 10
2 41401 1 10
2 41402 1 10
2 41403 1 10
2 41404 1 10
2 41405 1 10
2 41406 1 10
2 41407 1 10
2 41408 1 10
1 11 0 135 0
2 41409 1 11
2 41410 1 11
2 41411 1 11
2 41412 1 11
2 41413 1 11
2 41414 1 11
2 41415 1 11
2 41416 1 11
2 41417 1 11
2 41418 1 11
2 41419 1 11
2 41420 1 11
2 41421 1 11
2 41422 1 11
2 41423 1 11
2 41424 1 11
2 41425 1 11
2 41426 1 11
2 41427 1 11
2 41428 1 11
2 41429 1 11
2 41430 1 11
2 41431 1 11
2 41432 1 11
2 41433 1 11
2 41434 1 11
2 41435 1 11
2 41436 1 11
2 41437 1 11
2 41438 1 11
2 41439 1 11
2 41440 1 11
2 41441 1 11
2 41442 1 11
2 41443 1 11
2 41444 1 11
2 41445 1 11
2 41446 1 11
2 41447 1 11
2 41448 1 11
2 41449 1 11
2 41450 1 11
2 41451 1 11
2 41452 1 11
2 41453 1 11
2 41454 1 11
2 41455 1 11
2 41456 1 11
2 41457 1 11
2 41458 1 11
2 41459 1 11
2 41460 1 11
2 41461 1 11
2 41462 1 11
2 41463 1 11
2 41464 1 11
2 41465 1 11
2 41466 1 11
2 41467 1 11
2 41468 1 11
2 41469 1 11
2 41470 1 11
2 41471 1 11
2 41472 1 11
2 41473 1 11
2 41474 1 11
2 41475 1 11
2 41476 1 11
2 41477 1 11
2 41478 1 11
2 41479 1 11
2 41480 1 11
2 41481 1 11
2 41482 1 11
2 41483 1 11
2 41484 1 11
2 41485 1 11
2 41486 1 11
2 41487 1 11
2 41488 1 11
2 41489 1 11
2 41490 1 11
2 41491 1 11
2 41492 1 11
2 41493 1 11
2 41494 1 11
2 41495 1 11
2 41496 1 11
2 41497 1 11
2 41498 1 11
2 41499 1 11
2 41500 1 11
2 41501 1 11
2 41502 1 11
2 41503 1 11
2 41504 1 11
2 41505 1 11
2 41506 1 11
2 41507 1 11
2 41508 1 11
2 41509 1 11
2 41510 1 11
2 41511 1 11
2 41512 1 11
2 41513 1 11
2 41514 1 11
2 41515 1 11
2 41516 1 11
2 41517 1 11
2 41518 1 11
2 41519 1 11
2 41520 1 11
2 41521 1 11
2 41522 1 11
2 41523 1 11
2 41524 1 11
2 41525 1 11
2 41526 1 11
2 41527 1 11
2 41528 1 11
2 41529 1 11
2 41530 1 11
2 41531 1 11
2 41532 1 11
2 41533 1 11
2 41534 1 11
2 41535 1 11
2 41536 1 11
2 41537 1 11
2 41538 1 11
2 41539 1 11
2 41540 1 11
2 41541 1 11
2 41542 1 11
2 41543 1 11
1 12 0 145 0
2 41544 1 12
2 41545 1 12
2 41546 1 12
2 41547 1 12
2 41548 1 12
2 41549 1 12
2 41550 1 12
2 41551 1 12
2 41552 1 12
2 41553 1 12
2 41554 1 12
2 41555 1 12
2 41556 1 12
2 41557 1 12
2 41558 1 12
2 41559 1 12
2 41560 1 12
2 41561 1 12
2 41562 1 12
2 41563 1 12
2 41564 1 12
2 41565 1 12
2 41566 1 12
2 41567 1 12
2 41568 1 12
2 41569 1 12
2 41570 1 12
2 41571 1 12
2 41572 1 12
2 41573 1 12
2 41574 1 12
2 41575 1 12
2 41576 1 12
2 41577 1 12
2 41578 1 12
2 41579 1 12
2 41580 1 12
2 41581 1 12
2 41582 1 12
2 41583 1 12
2 41584 1 12
2 41585 1 12
2 41586 1 12
2 41587 1 12
2 41588 1 12
2 41589 1 12
2 41590 1 12
2 41591 1 12
2 41592 1 12
2 41593 1 12
2 41594 1 12
2 41595 1 12
2 41596 1 12
2 41597 1 12
2 41598 1 12
2 41599 1 12
2 41600 1 12
2 41601 1 12
2 41602 1 12
2 41603 1 12
2 41604 1 12
2 41605 1 12
2 41606 1 12
2 41607 1 12
2 41608 1 12
2 41609 1 12
2 41610 1 12
2 41611 1 12
2 41612 1 12
2 41613 1 12
2 41614 1 12
2 41615 1 12
2 41616 1 12
2 41617 1 12
2 41618 1 12
2 41619 1 12
2 41620 1 12
2 41621 1 12
2 41622 1 12
2 41623 1 12
2 41624 1 12
2 41625 1 12
2 41626 1 12
2 41627 1 12
2 41628 1 12
2 41629 1 12
2 41630 1 12
2 41631 1 12
2 41632 1 12
2 41633 1 12
2 41634 1 12
2 41635 1 12
2 41636 1 12
2 41637 1 12
2 41638 1 12
2 41639 1 12
2 41640 1 12
2 41641 1 12
2 41642 1 12
2 41643 1 12
2 41644 1 12
2 41645 1 12
2 41646 1 12
2 41647 1 12
2 41648 1 12
2 41649 1 12
2 41650 1 12
2 41651 1 12
2 41652 1 12
2 41653 1 12
2 41654 1 12
2 41655 1 12
2 41656 1 12
2 41657 1 12
2 41658 1 12
2 41659 1 12
2 41660 1 12
2 41661 1 12
2 41662 1 12
2 41663 1 12
2 41664 1 12
2 41665 1 12
2 41666 1 12
2 41667 1 12
2 41668 1 12
2 41669 1 12
2 41670 1 12
2 41671 1 12
2 41672 1 12
2 41673 1 12
2 41674 1 12
2 41675 1 12
2 41676 1 12
2 41677 1 12
2 41678 1 12
2 41679 1 12
2 41680 1 12
2 41681 1 12
2 41682 1 12
2 41683 1 12
2 41684 1 12
2 41685 1 12
2 41686 1 12
2 41687 1 12
2 41688 1 12
1 13 0 81 0
2 41689 1 13
2 41690 1 13
2 41691 1 13
2 41692 1 13
2 41693 1 13
2 41694 1 13
2 41695 1 13
2 41696 1 13
2 41697 1 13
2 41698 1 13
2 41699 1 13
2 41700 1 13
2 41701 1 13
2 41702 1 13
2 41703 1 13
2 41704 1 13
2 41705 1 13
2 41706 1 13
2 41707 1 13
2 41708 1 13
2 41709 1 13
2 41710 1 13
2 41711 1 13
2 41712 1 13
2 41713 1 13
2 41714 1 13
2 41715 1 13
2 41716 1 13
2 41717 1 13
2 41718 1 13
2 41719 1 13
2 41720 1 13
2 41721 1 13
2 41722 1 13
2 41723 1 13
2 41724 1 13
2 41725 1 13
2 41726 1 13
2 41727 1 13
2 41728 1 13
2 41729 1 13
2 41730 1 13
2 41731 1 13
2 41732 1 13
2 41733 1 13
2 41734 1 13
2 41735 1 13
2 41736 1 13
2 41737 1 13
2 41738 1 13
2 41739 1 13
2 41740 1 13
2 41741 1 13
2 41742 1 13
2 41743 1 13
2 41744 1 13
2 41745 1 13
2 41746 1 13
2 41747 1 13
2 41748 1 13
2 41749 1 13
2 41750 1 13
2 41751 1 13
2 41752 1 13
2 41753 1 13
2 41754 1 13
2 41755 1 13
2 41756 1 13
2 41757 1 13
2 41758 1 13
2 41759 1 13
2 41760 1 13
2 41761 1 13
2 41762 1 13
2 41763 1 13
2 41764 1 13
2 41765 1 13
2 41766 1 13
2 41767 1 13
2 41768 1 13
2 41769 1 13
1 14 0 54 0
2 41770 1 14
2 41771 1 14
2 41772 1 14
2 41773 1 14
2 41774 1 14
2 41775 1 14
2 41776 1 14
2 41777 1 14
2 41778 1 14
2 41779 1 14
2 41780 1 14
2 41781 1 14
2 41782 1 14
2 41783 1 14
2 41784 1 14
2 41785 1 14
2 41786 1 14
2 41787 1 14
2 41788 1 14
2 41789 1 14
2 41790 1 14
2 41791 1 14
2 41792 1 14
2 41793 1 14
2 41794 1 14
2 41795 1 14
2 41796 1 14
2 41797 1 14
2 41798 1 14
2 41799 1 14
2 41800 1 14
2 41801 1 14
2 41802 1 14
2 41803 1 14
2 41804 1 14
2 41805 1 14
2 41806 1 14
2 41807 1 14
2 41808 1 14
2 41809 1 14
2 41810 1 14
2 41811 1 14
2 41812 1 14
2 41813 1 14
2 41814 1 14
2 41815 1 14
2 41816 1 14
2 41817 1 14
2 41818 1 14
2 41819 1 14
2 41820 1 14
2 41821 1 14
2 41822 1 14
2 41823 1 14
1 15 0 30 0
2 41824 1 15
2 41825 1 15
2 41826 1 15
2 41827 1 15
2 41828 1 15
2 41829 1 15
2 41830 1 15
2 41831 1 15
2 41832 1 15
2 41833 1 15
2 41834 1 15
2 41835 1 15
2 41836 1 15
2 41837 1 15
2 41838 1 15
2 41839 1 15
2 41840 1 15
2 41841 1 15
2 41842 1 15
2 41843 1 15
2 41844 1 15
2 41845 1 15
2 41846 1 15
2 41847 1 15
2 41848 1 15
2 41849 1 15
2 41850 1 15
2 41851 1 15
2 41852 1 15
2 41853 1 15
1 16 0 151 0
2 41854 1 16
2 41855 1 16
2 41856 1 16
2 41857 1 16
2 41858 1 16
2 41859 1 16
2 41860 1 16
2 41861 1 16
2 41862 1 16
2 41863 1 16
2 41864 1 16
2 41865 1 16
2 41866 1 16
2 41867 1 16
2 41868 1 16
2 41869 1 16
2 41870 1 16
2 41871 1 16
2 41872 1 16
2 41873 1 16
2 41874 1 16
2 41875 1 16
2 41876 1 16
2 41877 1 16
2 41878 1 16
2 41879 1 16
2 41880 1 16
2 41881 1 16
2 41882 1 16
2 41883 1 16
2 41884 1 16
2 41885 1 16
2 41886 1 16
2 41887 1 16
2 41888 1 16
2 41889 1 16
2 41890 1 16
2 41891 1 16
2 41892 1 16
2 41893 1 16
2 41894 1 16
2 41895 1 16
2 41896 1 16
2 41897 1 16
2 41898 1 16
2 41899 1 16
2 41900 1 16
2 41901 1 16
2 41902 1 16
2 41903 1 16
2 41904 1 16
2 41905 1 16
2 41906 1 16
2 41907 1 16
2 41908 1 16
2 41909 1 16
2 41910 1 16
2 41911 1 16
2 41912 1 16
2 41913 1 16
2 41914 1 16
2 41915 1 16
2 41916 1 16
2 41917 1 16
2 41918 1 16
2 41919 1 16
2 41920 1 16
2 41921 1 16
2 41922 1 16
2 41923 1 16
2 41924 1 16
2 41925 1 16
2 41926 1 16
2 41927 1 16
2 41928 1 16
2 41929 1 16
2 41930 1 16
2 41931 1 16
2 41932 1 16
2 41933 1 16
2 41934 1 16
2 41935 1 16
2 41936 1 16
2 41937 1 16
2 41938 1 16
2 41939 1 16
2 41940 1 16
2 41941 1 16
2 41942 1 16
2 41943 1 16
2 41944 1 16
2 41945 1 16
2 41946 1 16
2 41947 1 16
2 41948 1 16
2 41949 1 16
2 41950 1 16
2 41951 1 16
2 41952 1 16
2 41953 1 16
2 41954 1 16
2 41955 1 16
2 41956 1 16
2 41957 1 16
2 41958 1 16
2 41959 1 16
2 41960 1 16
2 41961 1 16
2 41962 1 16
2 41963 1 16
2 41964 1 16
2 41965 1 16
2 41966 1 16
2 41967 1 16
2 41968 1 16
2 41969 1 16
2 41970 1 16
2 41971 1 16
2 41972 1 16
2 41973 1 16
2 41974 1 16
2 41975 1 16
2 41976 1 16
2 41977 1 16
2 41978 1 16
2 41979 1 16
2 41980 1 16
2 41981 1 16
2 41982 1 16
2 41983 1 16
2 41984 1 16
2 41985 1 16
2 41986 1 16
2 41987 1 16
2 41988 1 16
2 41989 1 16
2 41990 1 16
2 41991 1 16
2 41992 1 16
2 41993 1 16
2 41994 1 16
2 41995 1 16
2 41996 1 16
2 41997 1 16
2 41998 1 16
2 41999 1 16
2 42000 1 16
2 42001 1 16
2 42002 1 16
2 42003 1 16
2 42004 1 16
1 17 0 208 0
2 42005 1 17
2 42006 1 17
2 42007 1 17
2 42008 1 17
2 42009 1 17
2 42010 1 17
2 42011 1 17
2 42012 1 17
2 42013 1 17
2 42014 1 17
2 42015 1 17
2 42016 1 17
2 42017 1 17
2 42018 1 17
2 42019 1 17
2 42020 1 17
2 42021 1 17
2 42022 1 17
2 42023 1 17
2 42024 1 17
2 42025 1 17
2 42026 1 17
2 42027 1 17
2 42028 1 17
2 42029 1 17
2 42030 1 17
2 42031 1 17
2 42032 1 17
2 42033 1 17
2 42034 1 17
2 42035 1 17
2 42036 1 17
2 42037 1 17
2 42038 1 17
2 42039 1 17
2 42040 1 17
2 42041 1 17
2 42042 1 17
2 42043 1 17
2 42044 1 17
2 42045 1 17
2 42046 1 17
2 42047 1 17
2 42048 1 17
2 42049 1 17
2 42050 1 17
2 42051 1 17
2 42052 1 17
2 42053 1 17
2 42054 1 17
2 42055 1 17
2 42056 1 17
2 42057 1 17
2 42058 1 17
2 42059 1 17
2 42060 1 17
2 42061 1 17
2 42062 1 17
2 42063 1 17
2 42064 1 17
2 42065 1 17
2 42066 1 17
2 42067 1 17
2 42068 1 17
2 42069 1 17
2 42070 1 17
2 42071 1 17
2 42072 1 17
2 42073 1 17
2 42074 1 17
2 42075 1 17
2 42076 1 17
2 42077 1 17
2 42078 1 17
2 42079 1 17
2 42080 1 17
2 42081 1 17
2 42082 1 17
2 42083 1 17
2 42084 1 17
2 42085 1 17
2 42086 1 17
2 42087 1 17
2 42088 1 17
2 42089 1 17
2 42090 1 17
2 42091 1 17
2 42092 1 17
2 42093 1 17
2 42094 1 17
2 42095 1 17
2 42096 1 17
2 42097 1 17
2 42098 1 17
2 42099 1 17
2 42100 1 17
2 42101 1 17
2 42102 1 17
2 42103 1 17
2 42104 1 17
2 42105 1 17
2 42106 1 17
2 42107 1 17
2 42108 1 17
2 42109 1 17
2 42110 1 17
2 42111 1 17
2 42112 1 17
2 42113 1 17
2 42114 1 17
2 42115 1 17
2 42116 1 17
2 42117 1 17
2 42118 1 17
2 42119 1 17
2 42120 1 17
2 42121 1 17
2 42122 1 17
2 42123 1 17
2 42124 1 17
2 42125 1 17
2 42126 1 17
2 42127 1 17
2 42128 1 17
2 42129 1 17
2 42130 1 17
2 42131 1 17
2 42132 1 17
2 42133 1 17
2 42134 1 17
2 42135 1 17
2 42136 1 17
2 42137 1 17
2 42138 1 17
2 42139 1 17
2 42140 1 17
2 42141 1 17
2 42142 1 17
2 42143 1 17
2 42144 1 17
2 42145 1 17
2 42146 1 17
2 42147 1 17
2 42148 1 17
2 42149 1 17
2 42150 1 17
2 42151 1 17
2 42152 1 17
2 42153 1 17
2 42154 1 17
2 42155 1 17
2 42156 1 17
2 42157 1 17
2 42158 1 17
2 42159 1 17
2 42160 1 17
2 42161 1 17
2 42162 1 17
2 42163 1 17
2 42164 1 17
2 42165 1 17
2 42166 1 17
2 42167 1 17
2 42168 1 17
2 42169 1 17
2 42170 1 17
2 42171 1 17
2 42172 1 17
2 42173 1 17
2 42174 1 17
2 42175 1 17
2 42176 1 17
2 42177 1 17
2 42178 1 17
2 42179 1 17
2 42180 1 17
2 42181 1 17
2 42182 1 17
2 42183 1 17
2 42184 1 17
2 42185 1 17
2 42186 1 17
2 42187 1 17
2 42188 1 17
2 42189 1 17
2 42190 1 17
2 42191 1 17
2 42192 1 17
2 42193 1 17
2 42194 1 17
2 42195 1 17
2 42196 1 17
2 42197 1 17
2 42198 1 17
2 42199 1 17
2 42200 1 17
2 42201 1 17
2 42202 1 17
2 42203 1 17
2 42204 1 17
2 42205 1 17
2 42206 1 17
2 42207 1 17
2 42208 1 17
2 42209 1 17
2 42210 1 17
2 42211 1 17
2 42212 1 17
1 18 0 237 0
2 42213 1 18
2 42214 1 18
2 42215 1 18
2 42216 1 18
2 42217 1 18
2 42218 1 18
2 42219 1 18
2 42220 1 18
2 42221 1 18
2 42222 1 18
2 42223 1 18
2 42224 1 18
2 42225 1 18
2 42226 1 18
2 42227 1 18
2 42228 1 18
2 42229 1 18
2 42230 1 18
2 42231 1 18
2 42232 1 18
2 42233 1 18
2 42234 1 18
2 42235 1 18
2 42236 1 18
2 42237 1 18
2 42238 1 18
2 42239 1 18
2 42240 1 18
2 42241 1 18
2 42242 1 18
2 42243 1 18
2 42244 1 18
2 42245 1 18
2 42246 1 18
2 42247 1 18
2 42248 1 18
2 42249 1 18
2 42250 1 18
2 42251 1 18
2 42252 1 18
2 42253 1 18
2 42254 1 18
2 42255 1 18
2 42256 1 18
2 42257 1 18
2 42258 1 18
2 42259 1 18
2 42260 1 18
2 42261 1 18
2 42262 1 18
2 42263 1 18
2 42264 1 18
2 42265 1 18
2 42266 1 18
2 42267 1 18
2 42268 1 18
2 42269 1 18
2 42270 1 18
2 42271 1 18
2 42272 1 18
2 42273 1 18
2 42274 1 18
2 42275 1 18
2 42276 1 18
2 42277 1 18
2 42278 1 18
2 42279 1 18
2 42280 1 18
2 42281 1 18
2 42282 1 18
2 42283 1 18
2 42284 1 18
2 42285 1 18
2 42286 1 18
2 42287 1 18
2 42288 1 18
2 42289 1 18
2 42290 1 18
2 42291 1 18
2 42292 1 18
2 42293 1 18
2 42294 1 18
2 42295 1 18
2 42296 1 18
2 42297 1 18
2 42298 1 18
2 42299 1 18
2 42300 1 18
2 42301 1 18
2 42302 1 18
2 42303 1 18
2 42304 1 18
2 42305 1 18
2 42306 1 18
2 42307 1 18
2 42308 1 18
2 42309 1 18
2 42310 1 18
2 42311 1 18
2 42312 1 18
2 42313 1 18
2 42314 1 18
2 42315 1 18
2 42316 1 18
2 42317 1 18
2 42318 1 18
2 42319 1 18
2 42320 1 18
2 42321 1 18
2 42322 1 18
2 42323 1 18
2 42324 1 18
2 42325 1 18
2 42326 1 18
2 42327 1 18
2 42328 1 18
2 42329 1 18
2 42330 1 18
2 42331 1 18
2 42332 1 18
2 42333 1 18
2 42334 1 18
2 42335 1 18
2 42336 1 18
2 42337 1 18
2 42338 1 18
2 42339 1 18
2 42340 1 18
2 42341 1 18
2 42342 1 18
2 42343 1 18
2 42344 1 18
2 42345 1 18
2 42346 1 18
2 42347 1 18
2 42348 1 18
2 42349 1 18
2 42350 1 18
2 42351 1 18
2 42352 1 18
2 42353 1 18
2 42354 1 18
2 42355 1 18
2 42356 1 18
2 42357 1 18
2 42358 1 18
2 42359 1 18
2 42360 1 18
2 42361 1 18
2 42362 1 18
2 42363 1 18
2 42364 1 18
2 42365 1 18
2 42366 1 18
2 42367 1 18
2 42368 1 18
2 42369 1 18
2 42370 1 18
2 42371 1 18
2 42372 1 18
2 42373 1 18
2 42374 1 18
2 42375 1 18
2 42376 1 18
2 42377 1 18
2 42378 1 18
2 42379 1 18
2 42380 1 18
2 42381 1 18
2 42382 1 18
2 42383 1 18
2 42384 1 18
2 42385 1 18
2 42386 1 18
2 42387 1 18
2 42388 1 18
2 42389 1 18
2 42390 1 18
2 42391 1 18
2 42392 1 18
2 42393 1 18
2 42394 1 18
2 42395 1 18
2 42396 1 18
2 42397 1 18
2 42398 1 18
2 42399 1 18
2 42400 1 18
2 42401 1 18
2 42402 1 18
2 42403 1 18
2 42404 1 18
2 42405 1 18
2 42406 1 18
2 42407 1 18
2 42408 1 18
2 42409 1 18
2 42410 1 18
2 42411 1 18
2 42412 1 18
2 42413 1 18
2 42414 1 18
2 42415 1 18
2 42416 1 18
2 42417 1 18
2 42418 1 18
2 42419 1 18
2 42420 1 18
2 42421 1 18
2 42422 1 18
2 42423 1 18
2 42424 1 18
2 42425 1 18
2 42426 1 18
2 42427 1 18
2 42428 1 18
2 42429 1 18
2 42430 1 18
2 42431 1 18
2 42432 1 18
2 42433 1 18
2 42434 1 18
2 42435 1 18
2 42436 1 18
2 42437 1 18
2 42438 1 18
2 42439 1 18
2 42440 1 18
2 42441 1 18
2 42442 1 18
2 42443 1 18
2 42444 1 18
2 42445 1 18
2 42446 1 18
2 42447 1 18
2 42448 1 18
2 42449 1 18
1 19 0 283 0
2 42450 1 19
2 42451 1 19
2 42452 1 19
2 42453 1 19
2 42454 1 19
2 42455 1 19
2 42456 1 19
2 42457 1 19
2 42458 1 19
2 42459 1 19
2 42460 1 19
2 42461 1 19
2 42462 1 19
2 42463 1 19
2 42464 1 19
2 42465 1 19
2 42466 1 19
2 42467 1 19
2 42468 1 19
2 42469 1 19
2 42470 1 19
2 42471 1 19
2 42472 1 19
2 42473 1 19
2 42474 1 19
2 42475 1 19
2 42476 1 19
2 42477 1 19
2 42478 1 19
2 42479 1 19
2 42480 1 19
2 42481 1 19
2 42482 1 19
2 42483 1 19
2 42484 1 19
2 42485 1 19
2 42486 1 19
2 42487 1 19
2 42488 1 19
2 42489 1 19
2 42490 1 19
2 42491 1 19
2 42492 1 19
2 42493 1 19
2 42494 1 19
2 42495 1 19
2 42496 1 19
2 42497 1 19
2 42498 1 19
2 42499 1 19
2 42500 1 19
2 42501 1 19
2 42502 1 19
2 42503 1 19
2 42504 1 19
2 42505 1 19
2 42506 1 19
2 42507 1 19
2 42508 1 19
2 42509 1 19
2 42510 1 19
2 42511 1 19
2 42512 1 19
2 42513 1 19
2 42514 1 19
2 42515 1 19
2 42516 1 19
2 42517 1 19
2 42518 1 19
2 42519 1 19
2 42520 1 19
2 42521 1 19
2 42522 1 19
2 42523 1 19
2 42524 1 19
2 42525 1 19
2 42526 1 19
2 42527 1 19
2 42528 1 19
2 42529 1 19
2 42530 1 19
2 42531 1 19
2 42532 1 19
2 42533 1 19
2 42534 1 19
2 42535 1 19
2 42536 1 19
2 42537 1 19
2 42538 1 19
2 42539 1 19
2 42540 1 19
2 42541 1 19
2 42542 1 19
2 42543 1 19
2 42544 1 19
2 42545 1 19
2 42546 1 19
2 42547 1 19
2 42548 1 19
2 42549 1 19
2 42550 1 19
2 42551 1 19
2 42552 1 19
2 42553 1 19
2 42554 1 19
2 42555 1 19
2 42556 1 19
2 42557 1 19
2 42558 1 19
2 42559 1 19
2 42560 1 19
2 42561 1 19
2 42562 1 19
2 42563 1 19
2 42564 1 19
2 42565 1 19
2 42566 1 19
2 42567 1 19
2 42568 1 19
2 42569 1 19
2 42570 1 19
2 42571 1 19
2 42572 1 19
2 42573 1 19
2 42574 1 19
2 42575 1 19
2 42576 1 19
2 42577 1 19
2 42578 1 19
2 42579 1 19
2 42580 1 19
2 42581 1 19
2 42582 1 19
2 42583 1 19
2 42584 1 19
2 42585 1 19
2 42586 1 19
2 42587 1 19
2 42588 1 19
2 42589 1 19
2 42590 1 19
2 42591 1 19
2 42592 1 19
2 42593 1 19
2 42594 1 19
2 42595 1 19
2 42596 1 19
2 42597 1 19
2 42598 1 19
2 42599 1 19
2 42600 1 19
2 42601 1 19
2 42602 1 19
2 42603 1 19
2 42604 1 19
2 42605 1 19
2 42606 1 19
2 42607 1 19
2 42608 1 19
2 42609 1 19
2 42610 1 19
2 42611 1 19
2 42612 1 19
2 42613 1 19
2 42614 1 19
2 42615 1 19
2 42616 1 19
2 42617 1 19
2 42618 1 19
2 42619 1 19
2 42620 1 19
2 42621 1 19
2 42622 1 19
2 42623 1 19
2 42624 1 19
2 42625 1 19
2 42626 1 19
2 42627 1 19
2 42628 1 19
2 42629 1 19
2 42630 1 19
2 42631 1 19
2 42632 1 19
2 42633 1 19
2 42634 1 19
2 42635 1 19
2 42636 1 19
2 42637 1 19
2 42638 1 19
2 42639 1 19
2 42640 1 19
2 42641 1 19
2 42642 1 19
2 42643 1 19
2 42644 1 19
2 42645 1 19
2 42646 1 19
2 42647 1 19
2 42648 1 19
2 42649 1 19
2 42650 1 19
2 42651 1 19
2 42652 1 19
2 42653 1 19
2 42654 1 19
2 42655 1 19
2 42656 1 19
2 42657 1 19
2 42658 1 19
2 42659 1 19
2 42660 1 19
2 42661 1 19
2 42662 1 19
2 42663 1 19
2 42664 1 19
2 42665 1 19
2 42666 1 19
2 42667 1 19
2 42668 1 19
2 42669 1 19
2 42670 1 19
2 42671 1 19
2 42672 1 19
2 42673 1 19
2 42674 1 19
2 42675 1 19
2 42676 1 19
2 42677 1 19
2 42678 1 19
2 42679 1 19
2 42680 1 19
2 42681 1 19
2 42682 1 19
2 42683 1 19
2 42684 1 19
2 42685 1 19
2 42686 1 19
2 42687 1 19
2 42688 1 19
2 42689 1 19
2 42690 1 19
2 42691 1 19
2 42692 1 19
2 42693 1 19
2 42694 1 19
2 42695 1 19
2 42696 1 19
2 42697 1 19
2 42698 1 19
2 42699 1 19
2 42700 1 19
2 42701 1 19
2 42702 1 19
2 42703 1 19
2 42704 1 19
2 42705 1 19
2 42706 1 19
2 42707 1 19
2 42708 1 19
2 42709 1 19
2 42710 1 19
2 42711 1 19
2 42712 1 19
2 42713 1 19
2 42714 1 19
2 42715 1 19
2 42716 1 19
2 42717 1 19
2 42718 1 19
2 42719 1 19
2 42720 1 19
2 42721 1 19
2 42722 1 19
2 42723 1 19
2 42724 1 19
2 42725 1 19
2 42726 1 19
2 42727 1 19
2 42728 1 19
2 42729 1 19
2 42730 1 19
2 42731 1 19
2 42732 1 19
1 20 0 166 0
2 42733 1 20
2 42734 1 20
2 42735 1 20
2 42736 1 20
2 42737 1 20
2 42738 1 20
2 42739 1 20
2 42740 1 20
2 42741 1 20
2 42742 1 20
2 42743 1 20
2 42744 1 20
2 42745 1 20
2 42746 1 20
2 42747 1 20
2 42748 1 20
2 42749 1 20
2 42750 1 20
2 42751 1 20
2 42752 1 20
2 42753 1 20
2 42754 1 20
2 42755 1 20
2 42756 1 20
2 42757 1 20
2 42758 1 20
2 42759 1 20
2 42760 1 20
2 42761 1 20
2 42762 1 20
2 42763 1 20
2 42764 1 20
2 42765 1 20
2 42766 1 20
2 42767 1 20
2 42768 1 20
2 42769 1 20
2 42770 1 20
2 42771 1 20
2 42772 1 20
2 42773 1 20
2 42774 1 20
2 42775 1 20
2 42776 1 20
2 42777 1 20
2 42778 1 20
2 42779 1 20
2 42780 1 20
2 42781 1 20
2 42782 1 20
2 42783 1 20
2 42784 1 20
2 42785 1 20
2 42786 1 20
2 42787 1 20
2 42788 1 20
2 42789 1 20
2 42790 1 20
2 42791 1 20
2 42792 1 20
2 42793 1 20
2 42794 1 20
2 42795 1 20
2 42796 1 20
2 42797 1 20
2 42798 1 20
2 42799 1 20
2 42800 1 20
2 42801 1 20
2 42802 1 20
2 42803 1 20
2 42804 1 20
2 42805 1 20
2 42806 1 20
2 42807 1 20
2 42808 1 20
2 42809 1 20
2 42810 1 20
2 42811 1 20
2 42812 1 20
2 42813 1 20
2 42814 1 20
2 42815 1 20
2 42816 1 20
2 42817 1 20
2 42818 1 20
2 42819 1 20
2 42820 1 20
2 42821 1 20
2 42822 1 20
2 42823 1 20
2 42824 1 20
2 42825 1 20
2 42826 1 20
2 42827 1 20
2 42828 1 20
2 42829 1 20
2 42830 1 20
2 42831 1 20
2 42832 1 20
2 42833 1 20
2 42834 1 20
2 42835 1 20
2 42836 1 20
2 42837 1 20
2 42838 1 20
2 42839 1 20
2 42840 1 20
2 42841 1 20
2 42842 1 20
2 42843 1 20
2 42844 1 20
2 42845 1 20
2 42846 1 20
2 42847 1 20
2 42848 1 20
2 42849 1 20
2 42850 1 20
2 42851 1 20
2 42852 1 20
2 42853 1 20
2 42854 1 20
2 42855 1 20
2 42856 1 20
2 42857 1 20
2 42858 1 20
2 42859 1 20
2 42860 1 20
2 42861 1 20
2 42862 1 20
2 42863 1 20
2 42864 1 20
2 42865 1 20
2 42866 1 20
2 42867 1 20
2 42868 1 20
2 42869 1 20
2 42870 1 20
2 42871 1 20
2 42872 1 20
2 42873 1 20
2 42874 1 20
2 42875 1 20
2 42876 1 20
2 42877 1 20
2 42878 1 20
2 42879 1 20
2 42880 1 20
2 42881 1 20
2 42882 1 20
2 42883 1 20
2 42884 1 20
2 42885 1 20
2 42886 1 20
2 42887 1 20
2 42888 1 20
2 42889 1 20
2 42890 1 20
2 42891 1 20
2 42892 1 20
2 42893 1 20
2 42894 1 20
2 42895 1 20
2 42896 1 20
2 42897 1 20
2 42898 1 20
1 21 0 150 0
2 42899 1 21
2 42900 1 21
2 42901 1 21
2 42902 1 21
2 42903 1 21
2 42904 1 21
2 42905 1 21
2 42906 1 21
2 42907 1 21
2 42908 1 21
2 42909 1 21
2 42910 1 21
2 42911 1 21
2 42912 1 21
2 42913 1 21
2 42914 1 21
2 42915 1 21
2 42916 1 21
2 42917 1 21
2 42918 1 21
2 42919 1 21
2 42920 1 21
2 42921 1 21
2 42922 1 21
2 42923 1 21
2 42924 1 21
2 42925 1 21
2 42926 1 21
2 42927 1 21
2 42928 1 21
2 42929 1 21
2 42930 1 21
2 42931 1 21
2 42932 1 21
2 42933 1 21
2 42934 1 21
2 42935 1 21
2 42936 1 21
2 42937 1 21
2 42938 1 21
2 42939 1 21
2 42940 1 21
2 42941 1 21
2 42942 1 21
2 42943 1 21
2 42944 1 21
2 42945 1 21
2 42946 1 21
2 42947 1 21
2 42948 1 21
2 42949 1 21
2 42950 1 21
2 42951 1 21
2 42952 1 21
2 42953 1 21
2 42954 1 21
2 42955 1 21
2 42956 1 21
2 42957 1 21
2 42958 1 21
2 42959 1 21
2 42960 1 21
2 42961 1 21
2 42962 1 21
2 42963 1 21
2 42964 1 21
2 42965 1 21
2 42966 1 21
2 42967 1 21
2 42968 1 21
2 42969 1 21
2 42970 1 21
2 42971 1 21
2 42972 1 21
2 42973 1 21
2 42974 1 21
2 42975 1 21
2 42976 1 21
2 42977 1 21
2 42978 1 21
2 42979 1 21
2 42980 1 21
2 42981 1 21
2 42982 1 21
2 42983 1 21
2 42984 1 21
2 42985 1 21
2 42986 1 21
2 42987 1 21
2 42988 1 21
2 42989 1 21
2 42990 1 21
2 42991 1 21
2 42992 1 21
2 42993 1 21
2 42994 1 21
2 42995 1 21
2 42996 1 21
2 42997 1 21
2 42998 1 21
2 42999 1 21
2 43000 1 21
2 43001 1 21
2 43002 1 21
2 43003 1 21
2 43004 1 21
2 43005 1 21
2 43006 1 21
2 43007 1 21
2 43008 1 21
2 43009 1 21
2 43010 1 21
2 43011 1 21
2 43012 1 21
2 43013 1 21
2 43014 1 21
2 43015 1 21
2 43016 1 21
2 43017 1 21
2 43018 1 21
2 43019 1 21
2 43020 1 21
2 43021 1 21
2 43022 1 21
2 43023 1 21
2 43024 1 21
2 43025 1 21
2 43026 1 21
2 43027 1 21
2 43028 1 21
2 43029 1 21
2 43030 1 21
2 43031 1 21
2 43032 1 21
2 43033 1 21
2 43034 1 21
2 43035 1 21
2 43036 1 21
2 43037 1 21
2 43038 1 21
2 43039 1 21
2 43040 1 21
2 43041 1 21
2 43042 1 21
2 43043 1 21
2 43044 1 21
2 43045 1 21
2 43046 1 21
2 43047 1 21
2 43048 1 21
1 22 0 117 0
2 43049 1 22
2 43050 1 22
2 43051 1 22
2 43052 1 22
2 43053 1 22
2 43054 1 22
2 43055 1 22
2 43056 1 22
2 43057 1 22
2 43058 1 22
2 43059 1 22
2 43060 1 22
2 43061 1 22
2 43062 1 22
2 43063 1 22
2 43064 1 22
2 43065 1 22
2 43066 1 22
2 43067 1 22
2 43068 1 22
2 43069 1 22
2 43070 1 22
2 43071 1 22
2 43072 1 22
2 43073 1 22
2 43074 1 22
2 43075 1 22
2 43076 1 22
2 43077 1 22
2 43078 1 22
2 43079 1 22
2 43080 1 22
2 43081 1 22
2 43082 1 22
2 43083 1 22
2 43084 1 22
2 43085 1 22
2 43086 1 22
2 43087 1 22
2 43088 1 22
2 43089 1 22
2 43090 1 22
2 43091 1 22
2 43092 1 22
2 43093 1 22
2 43094 1 22
2 43095 1 22
2 43096 1 22
2 43097 1 22
2 43098 1 22
2 43099 1 22
2 43100 1 22
2 43101 1 22
2 43102 1 22
2 43103 1 22
2 43104 1 22
2 43105 1 22
2 43106 1 22
2 43107 1 22
2 43108 1 22
2 43109 1 22
2 43110 1 22
2 43111 1 22
2 43112 1 22
2 43113 1 22
2 43114 1 22
2 43115 1 22
2 43116 1 22
2 43117 1 22
2 43118 1 22
2 43119 1 22
2 43120 1 22
2 43121 1 22
2 43122 1 22
2 43123 1 22
2 43124 1 22
2 43125 1 22
2 43126 1 22
2 43127 1 22
2 43128 1 22
2 43129 1 22
2 43130 1 22
2 43131 1 22
2 43132 1 22
2 43133 1 22
2 43134 1 22
2 43135 1 22
2 43136 1 22
2 43137 1 22
2 43138 1 22
2 43139 1 22
2 43140 1 22
2 43141 1 22
2 43142 1 22
2 43143 1 22
2 43144 1 22
2 43145 1 22
2 43146 1 22
2 43147 1 22
2 43148 1 22
2 43149 1 22
2 43150 1 22
2 43151 1 22
2 43152 1 22
2 43153 1 22
2 43154 1 22
2 43155 1 22
2 43156 1 22
2 43157 1 22
2 43158 1 22
2 43159 1 22
2 43160 1 22
2 43161 1 22
2 43162 1 22
2 43163 1 22
2 43164 1 22
2 43165 1 22
1 23 0 113 0
2 43166 1 23
2 43167 1 23
2 43168 1 23
2 43169 1 23
2 43170 1 23
2 43171 1 23
2 43172 1 23
2 43173 1 23
2 43174 1 23
2 43175 1 23
2 43176 1 23
2 43177 1 23
2 43178 1 23
2 43179 1 23
2 43180 1 23
2 43181 1 23
2 43182 1 23
2 43183 1 23
2 43184 1 23
2 43185 1 23
2 43186 1 23
2 43187 1 23
2 43188 1 23
2 43189 1 23
2 43190 1 23
2 43191 1 23
2 43192 1 23
2 43193 1 23
2 43194 1 23
2 43195 1 23
2 43196 1 23
2 43197 1 23
2 43198 1 23
2 43199 1 23
2 43200 1 23
2 43201 1 23
2 43202 1 23
2 43203 1 23
2 43204 1 23
2 43205 1 23
2 43206 1 23
2 43207 1 23
2 43208 1 23
2 43209 1 23
2 43210 1 23
2 43211 1 23
2 43212 1 23
2 43213 1 23
2 43214 1 23
2 43215 1 23
2 43216 1 23
2 43217 1 23
2 43218 1 23
2 43219 1 23
2 43220 1 23
2 43221 1 23
2 43222 1 23
2 43223 1 23
2 43224 1 23
2 43225 1 23
2 43226 1 23
2 43227 1 23
2 43228 1 23
2 43229 1 23
2 43230 1 23
2 43231 1 23
2 43232 1 23
2 43233 1 23
2 43234 1 23
2 43235 1 23
2 43236 1 23
2 43237 1 23
2 43238 1 23
2 43239 1 23
2 43240 1 23
2 43241 1 23
2 43242 1 23
2 43243 1 23
2 43244 1 23
2 43245 1 23
2 43246 1 23
2 43247 1 23
2 43248 1 23
2 43249 1 23
2 43250 1 23
2 43251 1 23
2 43252 1 23
2 43253 1 23
2 43254 1 23
2 43255 1 23
2 43256 1 23
2 43257 1 23
2 43258 1 23
2 43259 1 23
2 43260 1 23
2 43261 1 23
2 43262 1 23
2 43263 1 23
2 43264 1 23
2 43265 1 23
2 43266 1 23
2 43267 1 23
2 43268 1 23
2 43269 1 23
2 43270 1 23
2 43271 1 23
2 43272 1 23
2 43273 1 23
2 43274 1 23
2 43275 1 23
2 43276 1 23
2 43277 1 23
2 43278 1 23
1 24 0 6 0
2 43279 1 24
2 43280 1 24
2 43281 1 24
2 43282 1 24
2 43283 1 24
2 43284 1 24
2 43285 1 27
2 43286 1 27
2 43287 1 27
2 43288 1 27
2 43289 1 27
2 43290 1 27
2 43291 1 27
2 43292 1 27
2 43293 1 27
2 43294 1 27
2 43295 1 27
2 43296 1 27
2 43297 1 27
2 43298 1 27
2 43299 1 27
2 43300 1 27
2 43301 1 27
2 43302 1 27
2 43303 1 27
2 43304 1 27
2 43305 1 27
2 43306 1 27
2 43307 1 27
2 43308 1 27
2 43309 1 27
2 43310 1 27
2 43311 1 27
2 43312 1 27
2 43313 1 27
2 43314 1 27
2 43315 1 27
2 43316 1 27
2 43317 1 27
2 43318 1 27
2 43319 1 27
2 43320 1 27
2 43321 1 27
2 43322 1 27
2 43323 1 27
2 43324 1 27
2 43325 1 27
2 43326 1 27
2 43327 1 27
2 43328 1 27
2 43329 1 27
2 43330 1 27
2 43331 1 27
2 43332 1 27
2 43333 1 27
2 43334 1 27
2 43335 1 27
2 43336 1 27
2 43337 1 27
2 43338 1 27
2 43339 1 27
2 43340 1 27
2 43341 1 27
2 43342 1 27
2 43343 1 27
2 43344 1 27
2 43345 1 27
2 43346 1 27
2 43347 1 27
2 43348 1 27
2 43349 1 27
2 43350 1 27
2 43351 1 27
2 43352 1 27
2 43353 1 27
2 43354 1 27
2 43355 1 27
2 43356 1 27
2 43357 1 27
2 43358 1 27
2 43359 1 27
2 43360 1 27
2 43361 1 27
2 43362 1 27
2 43363 1 27
2 43364 1 27
2 43365 1 27
2 43366 1 27
2 43367 1 27
2 43368 1 27
2 43369 1 27
2 43370 1 27
2 43371 1 27
2 43372 1 27
2 43373 1 27
2 43374 1 27
2 43375 1 27
2 43376 1 27
2 43377 1 27
2 43378 1 27
2 43379 1 27
2 43380 1 27
2 43381 1 27
2 43382 1 27
2 43383 1 27
2 43384 1 27
2 43385 1 27
2 43386 1 27
2 43387 1 27
2 43388 1 27
2 43389 1 27
2 43390 1 27
2 43391 1 27
2 43392 1 27
2 43393 1 27
2 43394 1 27
2 43395 1 27
2 43396 1 27
2 43397 1 27
2 43398 1 27
2 43399 1 27
2 43400 1 27
2 43401 1 27
2 43402 1 27
2 43403 1 27
2 43404 1 27
2 43405 1 27
2 43406 1 27
2 43407 1 27
2 43408 1 27
2 43409 1 27
2 43410 1 27
2 43411 1 27
2 43412 1 27
2 43413 1 27
2 43414 1 27
2 43415 1 27
2 43416 1 27
2 43417 1 27
2 43418 1 27
2 43419 1 27
2 43420 1 27
2 43421 1 27
2 43422 1 27
2 43423 1 27
2 43424 1 27
2 43425 1 27
2 43426 1 27
2 43427 1 27
2 43428 1 27
2 43429 1 27
2 43430 1 27
2 43431 1 27
2 43432 1 27
2 43433 1 27
2 43434 1 27
2 43435 1 27
2 43436 1 27
2 43437 1 27
2 43438 1 27
2 43439 1 27
2 43440 1 27
2 43441 1 27
2 43442 1 27
2 43443 1 27
2 43444 1 27
2 43445 1 27
2 43446 1 27
2 43447 1 27
2 43448 1 27
2 43449 1 27
2 43450 1 27
2 43451 1 27
2 43452 1 27
2 43453 1 27
2 43454 1 27
2 43455 1 27
2 43456 1 27
2 43457 1 27
2 43458 1 27
2 43459 1 27
2 43460 1 27
2 43461 1 27
2 43462 1 27
2 43463 1 27
2 43464 1 27
2 43465 1 27
2 43466 1 27
2 43467 1 27
2 43468 1 28
2 43469 1 28
2 43470 1 28
2 43471 1 28
2 43472 1 28
2 43473 1 28
2 43474 1 28
2 43475 1 28
2 43476 1 28
2 43477 1 28
2 43478 1 28
2 43479 1 28
2 43480 1 28
2 43481 1 28
2 43482 1 28
2 43483 1 28
2 43484 1 28
2 43485 1 28
2 43486 1 28
2 43487 1 28
2 43488 1 28
2 43489 1 28
2 43490 1 28
2 43491 1 28
2 43492 1 28
2 43493 1 28
2 43494 1 28
2 43495 1 28
2 43496 1 28
2 43497 1 28
2 43498 1 28
2 43499 1 28
2 43500 1 28
2 43501 1 28
2 43502 1 28
2 43503 1 28
2 43504 1 28
2 43505 1 28
2 43506 1 28
2 43507 1 28
2 43508 1 28
2 43509 1 28
2 43510 1 28
2 43511 1 28
2 43512 1 28
2 43513 1 28
2 43514 1 28
2 43515 1 28
2 43516 1 28
2 43517 1 28
2 43518 1 28
2 43519 1 28
2 43520 1 28
2 43521 1 28
2 43522 1 28
2 43523 1 28
2 43524 1 28
2 43525 1 28
2 43526 1 28
2 43527 1 28
2 43528 1 28
2 43529 1 28
2 43530 1 28
2 43531 1 28
2 43532 1 28
2 43533 1 28
2 43534 1 28
2 43535 1 28
2 43536 1 28
2 43537 1 28
2 43538 1 28
2 43539 1 28
2 43540 1 28
2 43541 1 28
2 43542 1 28
2 43543 1 28
2 43544 1 28
2 43545 1 28
2 43546 1 28
2 43547 1 28
2 43548 1 28
2 43549 1 28
2 43550 1 28
2 43551 1 28
2 43552 1 28
2 43553 1 28
2 43554 1 28
2 43555 1 28
2 43556 1 28
2 43557 1 28
2 43558 1 28
2 43559 1 28
2 43560 1 28
2 43561 1 28
2 43562 1 28
2 43563 1 28
2 43564 1 28
2 43565 1 28
2 43566 1 28
2 43567 1 28
2 43568 1 28
2 43569 1 28
2 43570 1 28
2 43571 1 28
2 43572 1 28
2 43573 1 28
2 43574 1 28
2 43575 1 28
2 43576 1 28
2 43577 1 28
2 43578 1 28
2 43579 1 28
2 43580 1 28
2 43581 1 28
2 43582 1 28
2 43583 1 28
2 43584 1 28
2 43585 1 28
2 43586 1 28
2 43587 1 28
2 43588 1 28
2 43589 1 28
2 43590 1 28
2 43591 1 28
2 43592 1 28
2 43593 1 28
2 43594 1 28
2 43595 1 28
2 43596 1 28
2 43597 1 28
2 43598 1 28
2 43599 1 28
2 43600 1 28
2 43601 1 28
2 43602 1 28
2 43603 1 28
2 43604 1 28
2 43605 1 28
2 43606 1 28
2 43607 1 28
2 43608 1 28
2 43609 1 28
2 43610 1 28
2 43611 1 28
2 43612 1 28
2 43613 1 28
2 43614 1 28
2 43615 1 29
2 43616 1 29
2 43617 1 29
2 43618 1 29
2 43619 1 29
2 43620 1 29
2 43621 1 29
2 43622 1 29
2 43623 1 29
2 43624 1 29
2 43625 1 29
2 43626 1 29
2 43627 1 29
2 43628 1 29
2 43629 1 29
2 43630 1 29
2 43631 1 29
2 43632 1 29
2 43633 1 29
2 43634 1 29
2 43635 1 29
2 43636 1 29
2 43637 1 29
2 43638 1 29
2 43639 1 29
2 43640 1 29
2 43641 1 29
2 43642 1 29
2 43643 1 29
2 43644 1 29
2 43645 1 29
2 43646 1 29
2 43647 1 29
2 43648 1 29
2 43649 1 29
2 43650 1 29
2 43651 1 29
2 43652 1 29
2 43653 1 29
2 43654 1 29
2 43655 1 29
2 43656 1 29
2 43657 1 29
2 43658 1 29
2 43659 1 29
2 43660 1 29
2 43661 1 29
2 43662 1 29
2 43663 1 29
2 43664 1 29
2 43665 1 29
2 43666 1 29
2 43667 1 29
2 43668 1 29
2 43669 1 29
2 43670 1 29
2 43671 1 29
2 43672 1 29
2 43673 1 29
2 43674 1 29
2 43675 1 29
2 43676 1 29
2 43677 1 29
2 43678 1 29
2 43679 1 29
2 43680 1 29
2 43681 1 29
2 43682 1 29
2 43683 1 29
2 43684 1 29
2 43685 1 29
2 43686 1 29
2 43687 1 29
2 43688 1 29
2 43689 1 29
2 43690 1 29
2 43691 1 29
2 43692 1 29
2 43693 1 29
2 43694 1 29
2 43695 1 29
2 43696 1 29
2 43697 1 29
2 43698 1 29
2 43699 1 29
2 43700 1 29
2 43701 1 29
2 43702 1 29
2 43703 1 29
2 43704 1 29
2 43705 1 29
2 43706 1 29
2 43707 1 29
2 43708 1 29
2 43709 1 29
2 43710 1 29
2 43711 1 29
2 43712 1 29
2 43713 1 29
2 43714 1 29
2 43715 1 29
2 43716 1 29
2 43717 1 29
2 43718 1 29
2 43719 1 29
2 43720 1 29
2 43721 1 29
2 43722 1 29
2 43723 1 29
2 43724 1 29
2 43725 1 29
2 43726 1 29
2 43727 1 29
2 43728 1 29
2 43729 1 29
2 43730 1 29
2 43731 1 29
2 43732 1 29
2 43733 1 29
2 43734 1 29
2 43735 1 29
2 43736 1 29
2 43737 1 29
2 43738 1 29
2 43739 1 29
2 43740 1 29
2 43741 1 29
2 43742 1 29
2 43743 1 29
2 43744 1 29
2 43745 1 29
2 43746 1 29
2 43747 1 29
2 43748 1 29
2 43749 1 29
2 43750 1 29
2 43751 1 29
2 43752 1 29
2 43753 1 29
2 43754 1 29
2 43755 1 29
2 43756 1 29
2 43757 1 29
2 43758 1 29
2 43759 1 29
2 43760 1 29
2 43761 1 29
2 43762 1 29
2 43763 1 29
2 43764 1 29
2 43765 1 29
2 43766 1 29
2 43767 1 29
2 43768 1 29
2 43769 1 29
2 43770 1 29
2 43771 1 29
2 43772 1 29
2 43773 1 29
2 43774 1 29
2 43775 1 29
2 43776 1 29
2 43777 1 29
2 43778 1 29
2 43779 1 29
2 43780 1 29
2 43781 1 29
2 43782 1 29
2 43783 1 29
2 43784 1 29
2 43785 1 29
2 43786 1 29
2 43787 1 29
2 43788 1 29
2 43789 1 29
2 43790 1 29
2 43791 1 29
2 43792 1 29
2 43793 1 29
2 43794 1 29
2 43795 1 29
2 43796 1 29
2 43797 1 29
2 43798 1 29
2 43799 1 29
2 43800 1 29
2 43801 1 29
2 43802 1 29
2 43803 1 29
2 43804 1 29
2 43805 1 29
2 43806 1 29
2 43807 1 29
2 43808 1 29
2 43809 1 29
2 43810 1 29
2 43811 1 29
2 43812 1 29
2 43813 1 29
2 43814 1 29
2 43815 1 29
2 43816 1 29
2 43817 1 29
2 43818 1 29
2 43819 1 29
2 43820 1 29
2 43821 1 29
2 43822 1 29
2 43823 1 30
2 43824 1 30
2 43825 1 30
2 43826 1 30
2 43827 1 30
2 43828 1 30
2 43829 1 30
2 43830 1 30
2 43831 1 30
2 43832 1 30
2 43833 1 30
2 43834 1 30
2 43835 1 30
2 43836 1 30
2 43837 1 30
2 43838 1 30
2 43839 1 30
2 43840 1 30
2 43841 1 30
2 43842 1 30
2 43843 1 30
2 43844 1 30
2 43845 1 30
2 43846 1 30
2 43847 1 30
2 43848 1 30
2 43849 1 30
2 43850 1 30
2 43851 1 30
2 43852 1 30
2 43853 1 30
2 43854 1 30
2 43855 1 30
2 43856 1 30
2 43857 1 30
2 43858 1 30
2 43859 1 30
2 43860 1 30
2 43861 1 30
2 43862 1 30
2 43863 1 30
2 43864 1 30
2 43865 1 30
2 43866 1 30
2 43867 1 30
2 43868 1 30
2 43869 1 30
2 43870 1 30
2 43871 1 30
2 43872 1 30
2 43873 1 30
2 43874 1 30
2 43875 1 30
2 43876 1 30
2 43877 1 30
2 43878 1 30
2 43879 1 30
2 43880 1 30
2 43881 1 30
2 43882 1 30
2 43883 1 30
2 43884 1 30
2 43885 1 30
2 43886 1 30
2 43887 1 30
2 43888 1 30
2 43889 1 30
2 43890 1 30
2 43891 1 30
2 43892 1 30
2 43893 1 30
2 43894 1 30
2 43895 1 30
2 43896 1 30
2 43897 1 30
2 43898 1 30
2 43899 1 30
2 43900 1 30
2 43901 1 30
2 43902 1 30
2 43903 1 30
2 43904 1 30
2 43905 1 30
2 43906 1 30
2 43907 1 30
2 43908 1 30
2 43909 1 30
2 43910 1 30
2 43911 1 30
2 43912 1 30
2 43913 1 30
2 43914 1 30
2 43915 1 30
2 43916 1 30
2 43917 1 30
2 43918 1 30
2 43919 1 30
2 43920 1 30
2 43921 1 30
2 43922 1 30
2 43923 1 30
2 43924 1 30
2 43925 1 30
2 43926 1 30
2 43927 1 30
2 43928 1 30
2 43929 1 30
2 43930 1 30
2 43931 1 30
2 43932 1 30
2 43933 1 30
2 43934 1 30
2 43935 1 30
2 43936 1 30
2 43937 1 30
2 43938 1 30
2 43939 1 30
2 43940 1 30
2 43941 1 30
2 43942 1 30
2 43943 1 30
2 43944 1 30
2 43945 1 30
2 43946 1 30
2 43947 1 30
2 43948 1 30
2 43949 1 30
2 43950 1 30
2 43951 1 30
2 43952 1 30
2 43953 1 30
2 43954 1 30
2 43955 1 30
2 43956 1 30
2 43957 1 30
2 43958 1 30
2 43959 1 30
2 43960 1 30
2 43961 1 30
2 43962 1 30
2 43963 1 30
2 43964 1 30
2 43965 1 30
2 43966 1 30
2 43967 1 30
2 43968 1 30
2 43969 1 30
2 43970 1 30
2 43971 1 30
2 43972 1 30
2 43973 1 30
2 43974 1 30
2 43975 1 30
2 43976 1 30
2 43977 1 30
2 43978 1 30
2 43979 1 30
2 43980 1 30
2 43981 1 30
2 43982 1 31
2 43983 1 31
2 43984 1 31
2 43985 1 31
2 43986 1 31
2 43987 1 31
2 43988 1 31
2 43989 1 31
2 43990 1 31
2 43991 1 31
2 43992 1 31
2 43993 1 31
2 43994 1 31
2 43995 1 31
2 43996 1 31
2 43997 1 31
2 43998 1 31
2 43999 1 31
2 44000 1 31
2 44001 1 31
2 44002 1 31
2 44003 1 31
2 44004 1 31
2 44005 1 31
2 44006 1 31
2 44007 1 31
2 44008 1 31
2 44009 1 31
2 44010 1 31
2 44011 1 31
2 44012 1 31
2 44013 1 31
2 44014 1 31
2 44015 1 31
2 44016 1 31
2 44017 1 31
2 44018 1 31
2 44019 1 31
2 44020 1 31
2 44021 1 31
2 44022 1 31
2 44023 1 31
2 44024 1 31
2 44025 1 31
2 44026 1 31
2 44027 1 31
2 44028 1 31
2 44029 1 31
2 44030 1 31
2 44031 1 31
2 44032 1 31
2 44033 1 31
2 44034 1 31
2 44035 1 31
2 44036 1 31
2 44037 1 31
2 44038 1 31
2 44039 1 31
2 44040 1 31
2 44041 1 31
2 44042 1 31
2 44043 1 31
2 44044 1 31
2 44045 1 31
2 44046 1 31
2 44047 1 31
2 44048 1 31
2 44049 1 31
2 44050 1 31
2 44051 1 31
2 44052 1 31
2 44053 1 31
2 44054 1 31
2 44055 1 31
2 44056 1 31
2 44057 1 31
2 44058 1 31
2 44059 1 31
2 44060 1 31
2 44061 1 31
2 44062 1 31
2 44063 1 31
2 44064 1 31
2 44065 1 31
2 44066 1 31
2 44067 1 31
2 44068 1 31
2 44069 1 31
2 44070 1 31
2 44071 1 31
2 44072 1 31
2 44073 1 31
2 44074 1 31
2 44075 1 31
2 44076 1 31
2 44077 1 31
2 44078 1 31
2 44079 1 31
2 44080 1 31
2 44081 1 31
2 44082 1 31
2 44083 1 31
2 44084 1 31
2 44085 1 31
2 44086 1 31
2 44087 1 31
2 44088 1 31
2 44089 1 31
2 44090 1 31
2 44091 1 31
2 44092 1 31
2 44093 1 31
2 44094 1 31
2 44095 1 31
2 44096 1 31
2 44097 1 31
2 44098 1 31
2 44099 1 31
2 44100 1 31
2 44101 1 31
2 44102 1 31
2 44103 1 31
2 44104 1 31
2 44105 1 31
2 44106 1 31
2 44107 1 31
2 44108 1 31
2 44109 1 31
2 44110 1 31
2 44111 1 31
2 44112 1 31
2 44113 1 31
2 44114 1 31
2 44115 1 31
2 44116 1 31
2 44117 1 31
2 44118 1 31
2 44119 1 31
2 44120 1 31
2 44121 1 31
2 44122 1 31
2 44123 1 31
2 44124 1 31
2 44125 1 31
2 44126 1 31
2 44127 1 31
2 44128 1 31
2 44129 1 31
2 44130 1 31
2 44131 1 31
2 44132 1 31
2 44133 1 31
2 44134 1 31
2 44135 1 31
2 44136 1 31
2 44137 1 31
2 44138 1 31
2 44139 1 31
2 44140 1 31
2 44141 1 31
2 44142 1 31
2 44143 1 31
2 44144 1 31
2 44145 1 31
2 44146 1 31
2 44147 1 31
2 44148 1 31
2 44149 1 31
2 44150 1 31
2 44151 1 31
2 44152 1 31
2 44153 1 31
2 44154 1 31
2 44155 1 32
2 44156 1 32
2 44157 1 32
2 44158 1 32
2 44159 1 32
2 44160 1 32
2 44161 1 32
2 44162 1 32
2 44163 1 32
2 44164 1 32
2 44165 1 32
2 44166 1 32
2 44167 1 32
2 44168 1 32
2 44169 1 32
2 44170 1 32
2 44171 1 32
2 44172 1 32
2 44173 1 32
2 44174 1 32
2 44175 1 32
2 44176 1 32
2 44177 1 32
2 44178 1 32
2 44179 1 32
2 44180 1 32
2 44181 1 32
2 44182 1 32
2 44183 1 32
2 44184 1 32
2 44185 1 32
2 44186 1 32
2 44187 1 32
2 44188 1 32
2 44189 1 32
2 44190 1 32
2 44191 1 32
2 44192 1 32
2 44193 1 32
2 44194 1 32
2 44195 1 32
2 44196 1 32
2 44197 1 32
2 44198 1 32
2 44199 1 32
2 44200 1 32
2 44201 1 32
2 44202 1 32
2 44203 1 32
2 44204 1 32
2 44205 1 32
2 44206 1 32
2 44207 1 32
2 44208 1 32
2 44209 1 32
2 44210 1 32
2 44211 1 32
2 44212 1 32
2 44213 1 32
2 44214 1 32
2 44215 1 32
2 44216 1 32
2 44217 1 32
2 44218 1 32
2 44219 1 32
2 44220 1 32
2 44221 1 32
2 44222 1 32
2 44223 1 33
2 44224 1 33
2 44225 1 33
2 44226 1 33
2 44227 1 33
2 44228 1 33
2 44229 1 33
2 44230 1 33
2 44231 1 33
2 44232 1 33
2 44233 1 33
2 44234 1 33
2 44235 1 33
2 44236 1 33
2 44237 1 33
2 44238 1 33
2 44239 1 33
2 44240 1 33
2 44241 1 33
2 44242 1 33
2 44243 1 33
2 44244 1 33
2 44245 1 33
2 44246 1 33
2 44247 1 33
2 44248 1 33
2 44249 1 33
2 44250 1 33
2 44251 1 33
2 44252 1 33
2 44253 1 33
2 44254 1 33
2 44255 1 33
2 44256 1 33
2 44257 1 33
2 44258 1 33
2 44259 1 33
2 44260 1 33
2 44261 1 33
2 44262 1 33
2 44263 1 33
2 44264 1 33
2 44265 1 33
2 44266 1 33
2 44267 1 33
2 44268 1 33
2 44269 1 33
2 44270 1 33
2 44271 1 33
2 44272 1 33
2 44273 1 33
2 44274 1 33
2 44275 1 33
2 44276 1 33
2 44277 1 33
2 44278 1 33
2 44279 1 33
2 44280 1 33
2 44281 1 33
2 44282 1 33
2 44283 1 33
2 44284 1 33
2 44285 1 33
2 44286 1 33
2 44287 1 33
2 44288 1 33
2 44289 1 33
2 44290 1 33
2 44291 1 33
2 44292 1 33
2 44293 1 33
2 44294 1 33
2 44295 1 33
2 44296 1 33
2 44297 1 33
2 44298 1 33
2 44299 1 33
2 44300 1 33
2 44301 1 33
2 44302 1 33
2 44303 1 33
2 44304 1 33
2 44305 1 34
2 44306 1 34
2 44307 1 34
2 44308 1 34
2 44309 1 34
2 44310 1 34
2 44311 1 34
2 44312 1 34
2 44313 1 34
2 44314 1 34
2 44315 1 34
2 44316 1 34
2 44317 1 34
2 44318 1 34
2 44319 1 34
2 44320 1 34
2 44321 1 34
2 44322 1 34
2 44323 1 34
2 44324 1 34
2 44325 1 34
2 44326 1 34
2 44327 1 34
2 44328 1 34
2 44329 1 34
2 44330 1 34
2 44331 1 34
2 44332 1 34
2 44333 1 34
2 44334 1 34
2 44335 1 34
2 44336 1 34
2 44337 1 34
2 44338 1 34
2 44339 1 34
2 44340 1 34
2 44341 1 34
2 44342 1 34
2 44343 1 34
2 44344 1 34
2 44345 1 34
2 44346 1 34
2 44347 1 34
2 44348 1 34
2 44349 1 34
2 44350 1 34
2 44351 1 34
2 44352 1 34
2 44353 1 34
2 44354 1 34
2 44355 1 34
2 44356 1 34
2 44357 1 34
2 44358 1 34
2 44359 1 34
2 44360 1 34
2 44361 1 34
2 44362 1 34
2 44363 1 34
2 44364 1 34
2 44365 1 34
2 44366 1 34
2 44367 1 34
2 44368 1 34
2 44369 1 34
2 44370 1 34
2 44371 1 34
2 44372 1 34
2 44373 1 34
2 44374 1 34
2 44375 1 34
2 44376 1 35
2 44377 1 35
2 44378 1 35
2 44379 1 35
2 44380 1 35
2 44381 1 35
2 44382 1 35
2 44383 1 35
2 44384 1 35
2 44385 1 35
2 44386 1 35
2 44387 1 35
2 44388 1 35
2 44389 1 35
2 44390 1 35
2 44391 1 35
2 44392 1 35
2 44393 1 35
2 44394 1 35
2 44395 1 35
2 44396 1 35
2 44397 1 35
2 44398 1 35
2 44399 1 35
2 44400 1 35
2 44401 1 35
2 44402 1 35
2 44403 1 35
2 44404 1 35
2 44405 1 35
2 44406 1 35
2 44407 1 35
2 44408 1 35
2 44409 1 35
2 44410 1 35
2 44411 1 35
2 44412 1 35
2 44413 1 35
2 44414 1 35
2 44415 1 35
2 44416 1 35
2 44417 1 35
2 44418 1 35
2 44419 1 35
2 44420 1 35
2 44421 1 35
2 44422 1 35
2 44423 1 35
2 44424 1 35
2 44425 1 35
2 44426 1 35
2 44427 1 35
2 44428 1 35
2 44429 1 35
2 44430 1 35
2 44431 1 35
2 44432 1 35
2 44433 1 35
2 44434 1 35
2 44435 1 35
2 44436 1 35
2 44437 1 35
2 44438 1 35
2 44439 1 35
2 44440 1 35
2 44441 1 35
2 44442 1 35
2 44443 1 35
2 44444 1 35
2 44445 1 35
2 44446 1 35
2 44447 1 35
2 44448 1 35
2 44449 1 35
2 44450 1 35
2 44451 1 35
2 44452 1 35
2 44453 1 35
2 44454 1 35
2 44455 1 36
2 44456 1 36
2 44457 1 36
2 44458 1 36
2 44459 1 36
2 44460 1 36
2 44461 1 36
2 44462 1 36
2 44463 1 36
2 44464 1 36
2 44465 1 36
2 44466 1 36
2 44467 1 36
2 44468 1 36
2 44469 1 36
2 44470 1 36
2 44471 1 36
2 44472 1 36
2 44473 1 36
2 44474 1 36
2 44475 1 36
2 44476 1 36
2 44477 1 36
2 44478 1 36
2 44479 1 36
2 44480 1 36
2 44481 1 36
2 44482 1 36
2 44483 1 36
2 44484 1 36
2 44485 1 36
2 44486 1 36
2 44487 1 36
2 44488 1 36
2 44489 1 36
2 44490 1 36
2 44491 1 36
2 44492 1 36
2 44493 1 36
2 44494 1 36
2 44495 1 36
2 44496 1 36
2 44497 1 36
2 44498 1 36
2 44499 1 36
2 44500 1 36
2 44501 1 36
2 44502 1 36
2 44503 1 36
2 44504 1 36
2 44505 1 36
2 44506 1 36
2 44507 1 36
2 44508 1 36
2 44509 1 36
2 44510 1 36
2 44511 1 36
2 44512 1 36
2 44513 1 36
2 44514 1 36
2 44515 1 36
2 44516 1 36
2 44517 1 36
2 44518 1 36
2 44519 1 36
2 44520 1 36
2 44521 1 36
2 44522 1 36
2 44523 1 36
2 44524 1 36
2 44525 1 36
2 44526 1 36
2 44527 1 36
2 44528 1 36
2 44529 1 36
2 44530 1 36
2 44531 1 36
2 44532 1 36
2 44533 1 36
2 44534 1 36
2 44535 1 36
2 44536 1 36
2 44537 1 36
2 44538 1 36
2 44539 1 36
2 44540 1 36
2 44541 1 36
2 44542 1 36
2 44543 1 36
2 44544 1 36
2 44545 1 36
2 44546 1 36
2 44547 1 36
2 44548 1 36
2 44549 1 36
2 44550 1 36
2 44551 1 36
2 44552 1 36
2 44553 1 36
2 44554 1 36
2 44555 1 36
2 44556 1 36
2 44557 1 36
2 44558 1 36
2 44559 1 36
2 44560 1 36
2 44561 1 36
2 44562 1 36
2 44563 1 36
2 44564 1 36
2 44565 1 36
2 44566 1 36
2 44567 1 36
2 44568 1 36
2 44569 1 36
2 44570 1 36
2 44571 1 37
2 44572 1 37
2 44573 1 37
2 44574 1 37
2 44575 1 37
2 44576 1 37
2 44577 1 37
2 44578 1 37
2 44579 1 37
2 44580 1 37
2 44581 1 37
2 44582 1 37
2 44583 1 37
2 44584 1 37
2 44585 1 37
2 44586 1 37
2 44587 1 37
2 44588 1 37
2 44589 1 37
2 44590 1 37
2 44591 1 37
2 44592 1 37
2 44593 1 37
2 44594 1 37
2 44595 1 37
2 44596 1 37
2 44597 1 37
2 44598 1 37
2 44599 1 37
2 44600 1 37
2 44601 1 37
2 44602 1 37
2 44603 1 37
2 44604 1 37
2 44605 1 37
2 44606 1 37
2 44607 1 37
2 44608 1 37
2 44609 1 37
2 44610 1 37
2 44611 1 37
2 44612 1 37
2 44613 1 37
2 44614 1 37
2 44615 1 37
2 44616 1 37
2 44617 1 37
2 44618 1 37
2 44619 1 37
2 44620 1 37
2 44621 1 37
2 44622 1 37
2 44623 1 37
2 44624 1 37
2 44625 1 37
2 44626 1 37
2 44627 1 37
2 44628 1 37
2 44629 1 37
2 44630 1 37
2 44631 1 37
2 44632 1 37
2 44633 1 37
2 44634 1 37
2 44635 1 37
2 44636 1 37
2 44637 1 37
2 44638 1 37
2 44639 1 37
2 44640 1 37
2 44641 1 37
2 44642 1 37
2 44643 1 37
2 44644 1 37
2 44645 1 37
2 44646 1 37
2 44647 1 37
2 44648 1 37
2 44649 1 37
2 44650 1 37
2 44651 1 37
2 44652 1 37
2 44653 1 37
2 44654 1 37
2 44655 1 37
2 44656 1 37
2 44657 1 37
2 44658 1 37
2 44659 1 37
2 44660 1 37
2 44661 1 37
2 44662 1 37
2 44663 1 37
2 44664 1 37
2 44665 1 37
2 44666 1 37
2 44667 1 37
2 44668 1 37
2 44669 1 37
2 44670 1 37
2 44671 1 37
2 44672 1 37
2 44673 1 37
2 44674 1 37
2 44675 1 37
2 44676 1 37
2 44677 1 37
2 44678 1 37
2 44679 1 37
2 44680 1 37
2 44681 1 37
2 44682 1 37
2 44683 1 37
2 44684 1 37
2 44685 1 37
2 44686 1 37
2 44687 1 37
2 44688 1 37
2 44689 1 37
2 44690 1 37
2 44691 1 37
2 44692 1 37
2 44693 1 37
2 44694 1 37
2 44695 1 37
2 44696 1 37
2 44697 1 37
2 44698 1 37
2 44699 1 37
2 44700 1 37
2 44701 1 37
2 44702 1 37
2 44703 1 37
2 44704 1 37
2 44705 1 37
2 44706 1 37
2 44707 1 37
2 44708 1 38
2 44709 1 38
2 44710 1 38
2 44711 1 38
2 44712 1 38
2 44713 1 38
2 44714 1 38
2 44715 1 38
2 44716 1 38
2 44717 1 38
2 44718 1 38
2 44719 1 38
2 44720 1 38
2 44721 1 38
2 44722 1 38
2 44723 1 38
2 44724 1 38
2 44725 1 38
2 44726 1 38
2 44727 1 38
2 44728 1 38
2 44729 1 38
2 44730 1 38
2 44731 1 38
2 44732 1 38
2 44733 1 38
2 44734 1 38
2 44735 1 38
2 44736 1 38
2 44737 1 38
2 44738 1 38
2 44739 1 38
2 44740 1 38
2 44741 1 38
2 44742 1 38
2 44743 1 38
2 44744 1 38
2 44745 1 38
2 44746 1 38
2 44747 1 38
2 44748 1 38
2 44749 1 38
2 44750 1 38
2 44751 1 38
2 44752 1 38
2 44753 1 38
2 44754 1 38
2 44755 1 38
2 44756 1 38
2 44757 1 38
2 44758 1 38
2 44759 1 38
2 44760 1 38
2 44761 1 38
2 44762 1 38
2 44763 1 38
2 44764 1 38
2 44765 1 38
2 44766 1 38
2 44767 1 38
2 44768 1 38
2 44769 1 38
2 44770 1 38
2 44771 1 38
2 44772 1 38
2 44773 1 38
2 44774 1 38
2 44775 1 38
2 44776 1 38
2 44777 1 38
2 44778 1 38
2 44779 1 38
2 44780 1 38
2 44781 1 38
2 44782 1 38
2 44783 1 38
2 44784 1 38
2 44785 1 38
2 44786 1 38
2 44787 1 38
2 44788 1 38
2 44789 1 38
2 44790 1 38
2 44791 1 38
2 44792 1 38
2 44793 1 38
2 44794 1 38
2 44795 1 38
2 44796 1 38
2 44797 1 38
2 44798 1 38
2 44799 1 38
2 44800 1 38
2 44801 1 38
2 44802 1 38
2 44803 1 38
2 44804 1 38
2 44805 1 38
2 44806 1 38
2 44807 1 38
2 44808 1 38
2 44809 1 38
2 44810 1 38
2 44811 1 38
2 44812 1 38
2 44813 1 38
2 44814 1 38
2 44815 1 38
2 44816 1 38
2 44817 1 38
2 44818 1 38
2 44819 1 38
2 44820 1 38
2 44821 1 38
2 44822 1 38
2 44823 1 38
2 44824 1 38
2 44825 1 38
2 44826 1 38
2 44827 1 38
2 44828 1 38
2 44829 1 38
2 44830 1 38
2 44831 1 38
2 44832 1 38
2 44833 1 38
2 44834 1 38
2 44835 1 38
2 44836 1 38
2 44837 1 38
2 44838 1 38
2 44839 1 38
2 44840 1 38
2 44841 1 39
2 44842 1 39
2 44843 1 39
2 44844 1 39
2 44845 1 39
2 44846 1 39
2 44847 1 39
2 44848 1 39
2 44849 1 39
2 44850 1 39
2 44851 1 39
2 44852 1 39
2 44853 1 39
2 44854 1 39
2 44855 1 39
2 44856 1 39
2 44857 1 39
2 44858 1 39
2 44859 1 39
2 44860 1 39
2 44861 1 39
2 44862 1 39
2 44863 1 39
2 44864 1 39
2 44865 1 39
2 44866 1 39
2 44867 1 39
2 44868 1 39
2 44869 1 39
2 44870 1 39
2 44871 1 39
2 44872 1 39
2 44873 1 39
2 44874 1 39
2 44875 1 39
2 44876 1 39
2 44877 1 39
2 44878 1 39
2 44879 1 39
2 44880 1 39
2 44881 1 39
2 44882 1 39
2 44883 1 39
2 44884 1 39
2 44885 1 39
2 44886 1 39
2 44887 1 39
2 44888 1 39
2 44889 1 39
2 44890 1 39
2 44891 1 39
2 44892 1 39
2 44893 1 39
2 44894 1 39
2 44895 1 39
2 44896 1 39
2 44897 1 39
2 44898 1 39
2 44899 1 39
2 44900 1 39
2 44901 1 39
2 44902 1 39
2 44903 1 39
2 44904 1 39
2 44905 1 39
2 44906 1 39
2 44907 1 39
2 44908 1 39
2 44909 1 39
2 44910 1 39
2 44911 1 39
2 44912 1 39
2 44913 1 39
2 44914 1 39
2 44915 1 39
2 44916 1 39
2 44917 1 39
2 44918 1 39
2 44919 1 39
2 44920 1 39
2 44921 1 39
2 44922 1 39
2 44923 1 39
2 44924 1 39
2 44925 1 39
2 44926 1 39
2 44927 1 39
2 44928 1 39
2 44929 1 39
2 44930 1 39
2 44931 1 39
2 44932 1 39
2 44933 1 39
2 44934 1 39
2 44935 1 39
2 44936 1 39
2 44937 1 39
2 44938 1 39
2 44939 1 39
2 44940 1 39
2 44941 1 39
2 44942 1 39
2 44943 1 39
2 44944 1 39
2 44945 1 39
2 44946 1 39
2 44947 1 39
2 44948 1 39
2 44949 1 39
2 44950 1 39
2 44951 1 39
2 44952 1 39
2 44953 1 39
2 44954 1 39
2 44955 1 39
2 44956 1 39
2 44957 1 39
2 44958 1 39
2 44959 1 39
2 44960 1 39
2 44961 1 39
2 44962 1 39
2 44963 1 39
2 44964 1 39
2 44965 1 39
2 44966 1 39
2 44967 1 39
2 44968 1 39
2 44969 1 39
2 44970 1 39
2 44971 1 39
2 44972 1 39
2 44973 1 39
2 44974 1 39
2 44975 1 39
2 44976 1 39
2 44977 1 39
2 44978 1 39
2 44979 1 39
2 44980 1 39
2 44981 1 39
2 44982 1 39
2 44983 1 39
2 44984 1 40
2 44985 1 40
2 44986 1 40
2 44987 1 40
2 44988 1 40
2 44989 1 40
2 44990 1 40
2 44991 1 40
2 44992 1 40
2 44993 1 40
2 44994 1 40
2 44995 1 40
2 44996 1 40
2 44997 1 40
2 44998 1 40
2 44999 1 40
2 45000 1 40
2 45001 1 40
2 45002 1 40
2 45003 1 40
2 45004 1 40
2 45005 1 40
2 45006 1 40
2 45007 1 40
2 45008 1 40
2 45009 1 40
2 45010 1 40
2 45011 1 40
2 45012 1 40
2 45013 1 40
2 45014 1 40
2 45015 1 40
2 45016 1 40
2 45017 1 40
2 45018 1 40
2 45019 1 40
2 45020 1 40
2 45021 1 40
2 45022 1 40
2 45023 1 40
2 45024 1 40
2 45025 1 40
2 45026 1 40
2 45027 1 40
2 45028 1 40
2 45029 1 40
2 45030 1 40
2 45031 1 40
2 45032 1 40
2 45033 1 40
2 45034 1 40
2 45035 1 40
2 45036 1 40
2 45037 1 40
2 45038 1 40
2 45039 1 40
2 45040 1 40
2 45041 1 40
2 45042 1 40
2 45043 1 40
2 45044 1 40
2 45045 1 40
2 45046 1 40
2 45047 1 40
2 45048 1 40
2 45049 1 40
2 45050 1 40
2 45051 1 40
2 45052 1 40
2 45053 1 40
2 45054 1 40
2 45055 1 40
2 45056 1 40
2 45057 1 40
2 45058 1 40
2 45059 1 40
2 45060 1 40
2 45061 1 40
2 45062 1 40
2 45063 1 40
2 45064 1 40
2 45065 1 40
2 45066 1 41
2 45067 1 41
2 45068 1 41
2 45069 1 41
2 45070 1 41
2 45071 1 41
2 45072 1 41
2 45073 1 41
2 45074 1 41
2 45075 1 41
2 45076 1 41
2 45077 1 41
2 45078 1 41
2 45079 1 41
2 45080 1 41
2 45081 1 41
2 45082 1 41
2 45083 1 41
2 45084 1 41
2 45085 1 41
2 45086 1 41
2 45087 1 41
2 45088 1 41
2 45089 1 41
2 45090 1 41
2 45091 1 41
2 45092 1 41
2 45093 1 41
2 45094 1 41
2 45095 1 41
2 45096 1 41
2 45097 1 41
2 45098 1 41
2 45099 1 41
2 45100 1 41
2 45101 1 41
2 45102 1 41
2 45103 1 41
2 45104 1 41
2 45105 1 41
2 45106 1 41
2 45107 1 41
2 45108 1 41
2 45109 1 41
2 45110 1 41
2 45111 1 41
2 45112 1 41
2 45113 1 41
2 45114 1 41
2 45115 1 41
2 45116 1 41
2 45117 1 41
2 45118 1 41
2 45119 1 41
2 45120 1 41
2 45121 1 41
2 45122 1 41
2 45123 1 41
2 45124 1 41
2 45125 1 41
2 45126 1 41
2 45127 1 41
2 45128 1 41
2 45129 1 41
2 45130 1 41
2 45131 1 41
2 45132 1 41
2 45133 1 41
2 45134 1 41
2 45135 1 41
2 45136 1 41
2 45137 1 41
2 45138 1 41
2 45139 1 42
2 45140 1 42
2 45141 1 42
2 45142 1 42
2 45143 1 42
2 45144 1 42
2 45145 1 42
2 45146 1 42
2 45147 1 42
2 45148 1 42
2 45149 1 42
2 45150 1 42
2 45151 1 42
2 45152 1 42
2 45153 1 42
2 45154 1 42
2 45155 1 42
2 45156 1 42
2 45157 1 42
2 45158 1 42
2 45159 1 42
2 45160 1 42
2 45161 1 42
2 45162 1 42
2 45163 1 42
2 45164 1 42
2 45165 1 42
2 45166 1 42
2 45167 1 42
2 45168 1 42
2 45169 1 42
2 45170 1 42
2 45171 1 42
2 45172 1 42
2 45173 1 42
2 45174 1 42
2 45175 1 42
2 45176 1 42
2 45177 1 42
2 45178 1 42
2 45179 1 42
2 45180 1 42
2 45181 1 42
2 45182 1 42
2 45183 1 42
2 45184 1 42
2 45185 1 42
2 45186 1 42
2 45187 1 42
2 45188 1 42
2 45189 1 42
2 45190 1 42
2 45191 1 42
2 45192 1 42
2 45193 1 42
2 45194 1 42
2 45195 1 42
2 45196 1 42
2 45197 1 42
2 45198 1 42
2 45199 1 42
2 45200 1 42
2 45201 1 42
2 45202 1 42
2 45203 1 42
2 45204 1 42
2 45205 1 42
2 45206 1 42
2 45207 1 42
2 45208 1 43
2 45209 1 43
2 45210 1 43
2 45211 1 43
2 45212 1 43
2 45213 1 43
2 45214 1 43
2 45215 1 43
2 45216 1 43
2 45217 1 43
2 45218 1 43
2 45219 1 43
2 45220 1 43
2 45221 1 43
2 45222 1 43
2 45223 1 43
2 45224 1 43
2 45225 1 43
2 45226 1 43
2 45227 1 43
2 45228 1 43
2 45229 1 43
2 45230 1 43
2 45231 1 43
2 45232 1 43
2 45233 1 43
2 45234 1 43
2 45235 1 43
2 45236 1 43
2 45237 1 43
2 45238 1 43
2 45239 1 43
2 45240 1 43
2 45241 1 43
2 45242 1 43
2 45243 1 43
2 45244 1 43
2 45245 1 43
2 45246 1 43
2 45247 1 43
2 45248 1 43
2 45249 1 43
2 45250 1 43
2 45251 1 43
2 45252 1 43
2 45253 1 43
2 45254 1 43
2 45255 1 43
2 45256 1 43
2 45257 1 43
2 45258 1 43
2 45259 1 43
2 45260 1 43
2 45261 1 43
2 45262 1 43
2 45263 1 43
2 45264 1 43
2 45265 1 43
2 45266 1 43
2 45267 1 43
2 45268 1 43
2 45269 1 43
2 45270 1 43
2 45271 1 43
2 45272 1 43
2 45273 1 43
2 45274 1 43
2 45275 1 43
2 45276 1 43
2 45277 1 43
2 45278 1 43
2 45279 1 43
2 45280 1 43
2 45281 1 43
2 45282 1 43
2 45283 1 43
2 45284 1 43
2 45285 1 43
2 45286 1 43
2 45287 1 43
2 45288 1 43
2 45289 1 43
2 45290 1 43
2 45291 1 43
2 45292 1 43
2 45293 1 43
2 45294 1 43
2 45295 1 43
2 45296 1 43
2 45297 1 43
2 45298 1 43
2 45299 1 43
2 45300 1 43
2 45301 1 43
2 45302 1 43
2 45303 1 43
2 45304 1 43
2 45305 1 43
2 45306 1 43
2 45307 1 43
2 45308 1 43
2 45309 1 43
2 45310 1 43
2 45311 1 43
2 45312 1 43
2 45313 1 43
2 45314 1 43
2 45315 1 43
2 45316 1 43
2 45317 1 43
2 45318 1 43
2 45319 1 43
2 45320 1 43
2 45321 1 43
2 45322 1 43
2 45323 1 43
2 45324 1 43
2 45325 1 43
2 45326 1 43
2 45327 1 43
2 45328 1 43
2 45329 1 43
2 45330 1 43
2 45331 1 43
2 45332 1 43
2 45333 1 43
2 45334 1 43
2 45335 1 43
2 45336 1 43
2 45337 1 43
2 45338 1 43
2 45339 1 43
2 45340 1 43
2 45341 1 43
2 45342 1 43
2 45343 1 43
2 45344 1 43
2 45345 1 43
2 45346 1 43
2 45347 1 43
2 45348 1 43
2 45349 1 43
2 45350 1 43
2 45351 1 43
2 45352 1 43
2 45353 1 43
2 45354 1 43
2 45355 1 43
2 45356 1 43
2 45357 1 43
2 45358 1 43
2 45359 1 43
2 45360 1 43
2 45361 1 43
2 45362 1 43
2 45363 1 43
2 45364 1 44
2 45365 1 44
2 45366 1 44
2 45367 1 44
2 45368 1 44
2 45369 1 44
2 45370 1 44
2 45371 1 44
2 45372 1 44
2 45373 1 44
2 45374 1 44
2 45375 1 44
2 45376 1 44
2 45377 1 44
2 45378 1 44
2 45379 1 44
2 45380 1 44
2 45381 1 44
2 45382 1 44
2 45383 1 44
2 45384 1 44
2 45385 1 44
2 45386 1 44
2 45387 1 44
2 45388 1 44
2 45389 1 44
2 45390 1 44
2 45391 1 44
2 45392 1 44
2 45393 1 44
2 45394 1 44
2 45395 1 44
2 45396 1 44
2 45397 1 44
2 45398 1 44
2 45399 1 44
2 45400 1 44
2 45401 1 44
2 45402 1 44
2 45403 1 44
2 45404 1 44
2 45405 1 44
2 45406 1 44
2 45407 1 44
2 45408 1 44
2 45409 1 44
2 45410 1 44
2 45411 1 44
2 45412 1 44
2 45413 1 44
2 45414 1 44
2 45415 1 44
2 45416 1 44
2 45417 1 44
2 45418 1 44
2 45419 1 44
2 45420 1 44
2 45421 1 44
2 45422 1 44
2 45423 1 44
2 45424 1 44
2 45425 1 44
2 45426 1 44
2 45427 1 44
2 45428 1 44
2 45429 1 44
2 45430 1 44
2 45431 1 44
2 45432 1 44
2 45433 1 44
2 45434 1 44
2 45435 1 44
2 45436 1 44
2 45437 1 44
2 45438 1 44
2 45439 1 44
2 45440 1 44
2 45441 1 44
2 45442 1 44
2 45443 1 44
2 45444 1 44
2 45445 1 44
2 45446 1 44
2 45447 1 44
2 45448 1 44
2 45449 1 44
2 45450 1 44
2 45451 1 44
2 45452 1 44
2 45453 1 44
2 45454 1 44
2 45455 1 44
2 45456 1 44
2 45457 1 44
2 45458 1 44
2 45459 1 44
2 45460 1 44
2 45461 1 44
2 45462 1 44
2 45463 1 44
2 45464 1 44
2 45465 1 44
2 45466 1 44
2 45467 1 44
2 45468 1 44
2 45469 1 44
2 45470 1 44
2 45471 1 44
2 45472 1 44
2 45473 1 44
2 45474 1 44
2 45475 1 44
2 45476 1 44
2 45477 1 44
2 45478 1 44
2 45479 1 44
2 45480 1 44
2 45481 1 44
2 45482 1 44
2 45483 1 44
2 45484 1 44
2 45485 1 44
2 45486 1 44
2 45487 1 44
2 45488 1 44
2 45489 1 44
2 45490 1 44
2 45491 1 44
2 45492 1 44
2 45493 1 44
2 45494 1 44
2 45495 1 44
2 45496 1 44
2 45497 1 44
2 45498 1 44
2 45499 1 44
2 45500 1 44
2 45501 1 44
2 45502 1 44
2 45503 1 44
2 45504 1 44
2 45505 1 44
2 45506 1 44
2 45507 1 44
2 45508 1 44
2 45509 1 44
2 45510 1 44
2 45511 1 44
2 45512 1 44
2 45513 1 44
2 45514 1 44
2 45515 1 44
2 45516 1 44
2 45517 1 44
2 45518 1 44
2 45519 1 44
2 45520 1 44
2 45521 1 44
2 45522 1 44
2 45523 1 44
2 45524 1 44
2 45525 1 44
2 45526 1 44
2 45527 1 44
2 45528 1 44
2 45529 1 44
2 45530 1 44
2 45531 1 44
2 45532 1 44
2 45533 1 44
2 45534 1 44
2 45535 1 44
2 45536 1 44
2 45537 1 44
2 45538 1 44
2 45539 1 44
2 45540 1 44
2 45541 1 44
2 45542 1 44
2 45543 1 44
2 45544 1 45
2 45545 1 45
2 45546 1 45
2 45547 1 45
2 45548 1 45
2 45549 1 45
2 45550 1 45
2 45551 1 45
2 45552 1 45
2 45553 1 45
2 45554 1 45
2 45555 1 45
2 45556 1 45
2 45557 1 45
2 45558 1 45
2 45559 1 45
2 45560 1 45
2 45561 1 45
2 45562 1 45
2 45563 1 45
2 45564 1 45
2 45565 1 45
2 45566 1 45
2 45567 1 45
2 45568 1 45
2 45569 1 45
2 45570 1 45
2 45571 1 45
2 45572 1 45
2 45573 1 45
2 45574 1 45
2 45575 1 45
2 45576 1 45
2 45577 1 45
2 45578 1 45
2 45579 1 45
2 45580 1 45
2 45581 1 45
2 45582 1 45
2 45583 1 45
2 45584 1 45
2 45585 1 45
2 45586 1 45
2 45587 1 45
2 45588 1 45
2 45589 1 45
2 45590 1 45
2 45591 1 45
2 45592 1 45
2 45593 1 45
2 45594 1 45
2 45595 1 45
2 45596 1 45
2 45597 1 45
2 45598 1 45
2 45599 1 45
2 45600 1 45
2 45601 1 45
2 45602 1 45
2 45603 1 45
2 45604 1 45
2 45605 1 45
2 45606 1 45
2 45607 1 45
2 45608 1 45
2 45609 1 45
2 45610 1 45
2 45611 1 45
2 45612 1 45
2 45613 1 45
2 45614 1 45
2 45615 1 45
2 45616 1 45
2 45617 1 45
2 45618 1 45
2 45619 1 45
2 45620 1 45
2 45621 1 45
2 45622 1 45
2 45623 1 45
2 45624 1 45
2 45625 1 45
2 45626 1 45
2 45627 1 45
2 45628 1 45
2 45629 1 45
2 45630 1 45
2 45631 1 45
2 45632 1 45
2 45633 1 45
2 45634 1 45
2 45635 1 45
2 45636 1 45
2 45637 1 45
2 45638 1 45
2 45639 1 45
2 45640 1 45
2 45641 1 45
2 45642 1 45
2 45643 1 45
2 45644 1 45
2 45645 1 45
2 45646 1 45
2 45647 1 45
2 45648 1 45
2 45649 1 45
2 45650 1 45
2 45651 1 45
2 45652 1 45
2 45653 1 45
2 45654 1 45
2 45655 1 45
2 45656 1 45
2 45657 1 45
2 45658 1 45
2 45659 1 45
2 45660 1 45
2 45661 1 45
2 45662 1 45
2 45663 1 45
2 45664 1 45
2 45665 1 45
2 45666 1 45
2 45667 1 45
2 45668 1 45
2 45669 1 45
2 45670 1 45
2 45671 1 45
2 45672 1 45
2 45673 1 45
2 45674 1 45
2 45675 1 45
2 45676 1 45
2 45677 1 45
2 45678 1 45
2 45679 1 45
2 45680 1 45
2 45681 1 45
2 45682 1 45
2 45683 1 45
2 45684 1 45
2 45685 1 45
2 45686 1 45
2 45687 1 45
2 45688 1 45
2 45689 1 45
2 45690 1 45
2 45691 1 45
2 45692 1 45
2 45693 1 45
2 45694 1 45
2 45695 1 45
2 45696 1 45
2 45697 1 45
2 45698 1 45
2 45699 1 45
2 45700 1 45
2 45701 1 45
2 45702 1 45
2 45703 1 45
2 45704 1 45
2 45705 1 45
2 45706 1 45
2 45707 1 45
2 45708 1 45
2 45709 1 45
2 45710 1 45
2 45711 1 45
2 45712 1 45
2 45713 1 45
2 45714 1 45
2 45715 1 45
2 45716 1 45
2 45717 1 45
2 45718 1 45
2 45719 1 45
2 45720 1 45
2 45721 1 45
2 45722 1 45
2 45723 1 45
2 45724 1 45
2 45725 1 45
2 45726 1 45
2 45727 1 45
2 45728 1 45
2 45729 1 45
2 45730 1 45
2 45731 1 45
2 45732 1 45
2 45733 1 45
2 45734 1 45
2 45735 1 45
2 45736 1 45
2 45737 1 45
2 45738 1 45
2 45739 1 45
2 45740 1 45
2 45741 1 45
2 45742 1 45
2 45743 1 45
2 45744 1 45
2 45745 1 45
2 45746 1 45
2 45747 1 45
2 45748 1 45
2 45749 1 45
2 45750 1 45
2 45751 1 45
2 45752 1 45
2 45753 1 45
2 45754 1 45
2 45755 1 45
2 45756 1 45
2 45757 1 45
2 45758 1 45
2 45759 1 45
2 45760 1 45
2 45761 1 45
2 45762 1 45
2 45763 1 45
2 45764 1 45
2 45765 1 45
2 45766 1 45
2 45767 1 45
2 45768 1 45
2 45769 1 45
2 45770 1 45
2 45771 1 45
2 45772 1 45
2 45773 1 45
2 45774 1 45
2 45775 1 45
2 45776 1 45
2 45777 1 45
2 45778 1 45
2 45779 1 45
2 45780 1 45
2 45781 1 45
2 45782 1 45
2 45783 1 45
2 45784 1 45
2 45785 1 45
2 45786 1 45
2 45787 1 45
2 45788 1 45
2 45789 1 45
2 45790 1 45
2 45791 1 46
2 45792 1 46
2 45793 1 46
2 45794 1 46
2 45795 1 46
2 45796 1 46
2 45797 1 46
2 45798 1 46
2 45799 1 46
2 45800 1 46
2 45801 1 46
2 45802 1 46
2 45803 1 46
2 45804 1 46
2 45805 1 46
2 45806 1 46
2 45807 1 46
2 45808 1 46
2 45809 1 46
2 45810 1 46
2 45811 1 46
2 45812 1 46
2 45813 1 46
2 45814 1 46
2 45815 1 46
2 45816 1 46
2 45817 1 46
2 45818 1 46
2 45819 1 46
2 45820 1 46
2 45821 1 46
2 45822 1 46
2 45823 1 46
2 45824 1 46
2 45825 1 46
2 45826 1 46
2 45827 1 46
2 45828 1 46
2 45829 1 46
2 45830 1 46
2 45831 1 46
2 45832 1 46
2 45833 1 46
2 45834 1 46
2 45835 1 46
2 45836 1 46
2 45837 1 46
2 45838 1 46
2 45839 1 46
2 45840 1 46
2 45841 1 46
2 45842 1 46
2 45843 1 46
2 45844 1 46
2 45845 1 46
2 45846 1 46
2 45847 1 46
2 45848 1 46
2 45849 1 46
2 45850 1 46
2 45851 1 46
2 45852 1 46
2 45853 1 46
2 45854 1 46
2 45855 1 46
2 45856 1 46
2 45857 1 46
2 45858 1 46
2 45859 1 46
2 45860 1 46
2 45861 1 46
2 45862 1 46
2 45863 1 46
2 45864 1 46
2 45865 1 46
2 45866 1 46
2 45867 1 46
2 45868 1 46
2 45869 1 46
2 45870 1 46
2 45871 1 46
2 45872 1 46
2 45873 1 46
2 45874 1 46
2 45875 1 46
2 45876 1 46
2 45877 1 46
2 45878 1 46
2 45879 1 46
2 45880 1 46
2 45881 1 46
2 45882 1 46
2 45883 1 46
2 45884 1 46
2 45885 1 46
2 45886 1 46
2 45887 1 46
2 45888 1 46
2 45889 1 46
2 45890 1 46
2 45891 1 46
2 45892 1 46
2 45893 1 46
2 45894 1 46
2 45895 1 46
2 45896 1 46
2 45897 1 46
2 45898 1 46
2 45899 1 46
2 45900 1 46
2 45901 1 46
2 45902 1 46
2 45903 1 46
2 45904 1 46
2 45905 1 46
2 45906 1 46
2 45907 1 46
2 45908 1 46
2 45909 1 46
2 45910 1 46
2 45911 1 46
2 45912 1 46
2 45913 1 46
2 45914 1 46
2 45915 1 46
2 45916 1 46
2 45917 1 46
2 45918 1 46
2 45919 1 46
2 45920 1 46
2 45921 1 46
2 45922 1 46
2 45923 1 46
2 45924 1 46
2 45925 1 46
2 45926 1 46
2 45927 1 46
2 45928 1 46
2 45929 1 46
2 45930 1 46
2 45931 1 46
2 45932 1 46
2 45933 1 46
2 45934 1 46
2 45935 1 46
2 45936 1 46
2 45937 1 46
2 45938 1 46
2 45939 1 46
2 45940 1 46
2 45941 1 46
2 45942 1 46
2 45943 1 46
2 45944 1 46
2 45945 1 46
2 45946 1 46
2 45947 1 46
2 45948 1 46
2 45949 1 46
2 45950 1 46
2 45951 1 46
2 45952 1 46
2 45953 1 46
2 45954 1 46
2 45955 1 46
2 45956 1 46
2 45957 1 46
2 45958 1 46
2 45959 1 46
2 45960 1 46
2 45961 1 46
2 45962 1 46
2 45963 1 46
2 45964 1 46
2 45965 1 46
2 45966 1 46
2 45967 1 46
2 45968 1 46
2 45969 1 46
2 45970 1 46
2 45971 1 46
2 45972 1 46
2 45973 1 46
2 45974 1 46
2 45975 1 46
2 45976 1 46
2 45977 1 46
2 45978 1 46
2 45979 1 46
2 45980 1 46
2 45981 1 46
2 45982 1 46
2 45983 1 46
2 45984 1 46
2 45985 1 46
2 45986 1 46
2 45987 1 46
2 45988 1 46
2 45989 1 46
2 45990 1 46
2 45991 1 46
2 45992 1 46
2 45993 1 46
2 45994 1 46
2 45995 1 46
2 45996 1 46
2 45997 1 46
2 45998 1 46
2 45999 1 46
2 46000 1 46
2 46001 1 46
2 46002 1 46
2 46003 1 46
2 46004 1 46
2 46005 1 46
2 46006 1 46
2 46007 1 47
2 46008 1 47
2 46009 1 47
2 46010 1 47
2 46011 1 47
2 46012 1 47
2 46013 1 47
2 46014 1 47
2 46015 1 47
2 46016 1 47
2 46017 1 47
2 46018 1 47
2 46019 1 47
2 46020 1 47
2 46021 1 47
2 46022 1 47
2 46023 1 47
2 46024 1 47
2 46025 1 47
2 46026 1 47
2 46027 1 47
2 46028 1 47
2 46029 1 47
2 46030 1 47
2 46031 1 47
2 46032 1 47
2 46033 1 47
2 46034 1 47
2 46035 1 47
2 46036 1 47
2 46037 1 47
2 46038 1 47
2 46039 1 47
2 46040 1 47
2 46041 1 47
2 46042 1 47
2 46043 1 47
2 46044 1 47
2 46045 1 47
2 46046 1 47
2 46047 1 47
2 46048 1 47
2 46049 1 47
2 46050 1 47
2 46051 1 47
2 46052 1 47
2 46053 1 47
2 46054 1 47
2 46055 1 47
2 46056 1 47
2 46057 1 47
2 46058 1 47
2 46059 1 47
2 46060 1 47
2 46061 1 47
2 46062 1 47
2 46063 1 47
2 46064 1 47
2 46065 1 47
2 46066 1 47
2 46067 1 47
2 46068 1 47
2 46069 1 47
2 46070 1 47
2 46071 1 47
2 46072 1 47
2 46073 1 47
2 46074 1 47
2 46075 1 47
2 46076 1 47
2 46077 1 47
2 46078 1 47
2 46079 1 47
2 46080 1 47
2 46081 1 47
2 46082 1 47
2 46083 1 47
2 46084 1 47
2 46085 1 47
2 46086 1 47
2 46087 1 47
2 46088 1 47
2 46089 1 47
2 46090 1 47
2 46091 1 47
2 46092 1 47
2 46093 1 47
2 46094 1 47
2 46095 1 47
2 46096 1 47
2 46097 1 47
2 46098 1 47
2 46099 1 47
2 46100 1 47
2 46101 1 47
2 46102 1 47
2 46103 1 47
2 46104 1 47
2 46105 1 47
2 46106 1 47
2 46107 1 47
2 46108 1 47
2 46109 1 47
2 46110 1 47
2 46111 1 47
2 46112 1 47
2 46113 1 47
2 46114 1 47
2 46115 1 47
2 46116 1 47
2 46117 1 47
2 46118 1 47
2 46119 1 47
2 46120 1 47
2 46121 1 47
2 46122 1 47
2 46123 1 47
2 46124 1 47
2 46125 1 47
2 46126 1 47
2 46127 1 47
2 46128 1 47
2 46129 1 47
2 46130 1 47
2 46131 1 47
2 46132 1 47
2 46133 1 47
2 46134 1 47
2 46135 1 47
2 46136 1 47
2 46137 1 47
2 46138 1 47
2 46139 1 47
2 46140 1 47
2 46141 1 47
2 46142 1 47
2 46143 1 47
2 46144 1 47
2 46145 1 47
2 46146 1 47
2 46147 1 47
2 46148 1 47
2 46149 1 47
2 46150 1 47
2 46151 1 47
2 46152 1 47
2 46153 1 47
2 46154 1 47
2 46155 1 47
2 46156 1 47
2 46157 1 47
2 46158 1 47
2 46159 1 47
2 46160 1 47
2 46161 1 47
2 46162 1 47
2 46163 1 47
2 46164 1 47
2 46165 1 47
2 46166 1 47
2 46167 1 47
2 46168 1 47
2 46169 1 47
2 46170 1 47
2 46171 1 47
2 46172 1 47
2 46173 1 47
2 46174 1 47
2 46175 1 47
2 46176 1 47
2 46177 1 47
2 46178 1 47
2 46179 1 47
2 46180 1 48
2 46181 1 48
2 46182 1 48
2 46183 1 48
2 46184 1 48
2 46185 1 48
2 46186 1 48
2 46187 1 48
2 46188 1 48
2 46189 1 48
2 46190 1 48
2 46191 1 48
2 46192 1 48
2 46193 1 48
2 46194 1 48
2 46195 1 48
2 46196 1 48
2 46197 1 48
2 46198 1 48
2 46199 1 48
2 46200 1 48
2 46201 1 48
2 46202 1 48
2 46203 1 48
2 46204 1 48
2 46205 1 48
2 46206 1 48
2 46207 1 48
2 46208 1 48
2 46209 1 48
2 46210 1 48
2 46211 1 48
2 46212 1 48
2 46213 1 48
2 46214 1 48
2 46215 1 48
2 46216 1 48
2 46217 1 48
2 46218 1 48
2 46219 1 48
2 46220 1 48
2 46221 1 48
2 46222 1 48
2 46223 1 48
2 46224 1 48
2 46225 1 48
2 46226 1 48
2 46227 1 48
2 46228 1 48
2 46229 1 48
2 46230 1 48
2 46231 1 48
2 46232 1 48
2 46233 1 48
2 46234 1 48
2 46235 1 48
2 46236 1 48
2 46237 1 48
2 46238 1 48
2 46239 1 48
2 46240 1 48
2 46241 1 48
2 46242 1 48
2 46243 1 48
2 46244 1 48
2 46245 1 48
2 46246 1 48
2 46247 1 48
2 46248 1 48
2 46249 1 48
2 46250 1 48
2 46251 1 48
2 46252 1 48
2 46253 1 48
2 46254 1 48
2 46255 1 48
2 46256 1 48
2 46257 1 48
2 46258 1 48
2 46259 1 48
2 46260 1 48
2 46261 1 48
2 46262 1 48
2 46263 1 48
2 46264 1 48
2 46265 1 48
2 46266 1 48
2 46267 1 48
2 46268 1 48
2 46269 1 48
2 46270 1 48
2 46271 1 48
2 46272 1 48
2 46273 1 48
2 46274 1 48
2 46275 1 48
2 46276 1 48
2 46277 1 48
2 46278 1 48
2 46279 1 48
2 46280 1 48
2 46281 1 48
2 46282 1 48
2 46283 1 48
2 46284 1 48
2 46285 1 48
2 46286 1 48
2 46287 1 48
2 46288 1 48
2 46289 1 48
2 46290 1 48
2 46291 1 48
2 46292 1 48
2 46293 1 48
2 46294 1 48
2 46295 1 48
2 46296 1 48
2 46297 1 48
2 46298 1 48
2 46299 1 48
2 46300 1 48
2 46301 1 48
2 46302 1 48
2 46303 1 48
2 46304 1 48
2 46305 1 48
2 46306 1 48
2 46307 1 48
2 46308 1 48
2 46309 1 48
2 46310 1 48
2 46311 1 48
2 46312 1 48
2 46313 1 48
2 46314 1 48
2 46315 1 48
2 46316 1 48
2 46317 1 48
2 46318 1 48
2 46319 1 48
2 46320 1 48
2 46321 1 48
2 46322 1 49
2 46323 1 49
2 46324 1 49
2 46325 1 49
2 46326 1 49
2 46327 1 49
2 46328 1 49
2 46329 1 49
2 46330 1 49
2 46331 1 49
2 46332 1 49
2 46333 1 49
2 46334 1 49
2 46335 1 49
2 46336 1 49
2 46337 1 49
2 46338 1 49
2 46339 1 49
2 46340 1 49
2 46341 1 49
2 46342 1 49
2 46343 1 49
2 46344 1 49
2 46345 1 49
2 46346 1 49
2 46347 1 49
2 46348 1 49
2 46349 1 49
2 46350 1 49
2 46351 1 49
2 46352 1 49
2 46353 1 49
2 46354 1 49
2 46355 1 49
2 46356 1 49
2 46357 1 49
2 46358 1 49
2 46359 1 49
2 46360 1 49
2 46361 1 49
2 46362 1 49
2 46363 1 49
2 46364 1 49
2 46365 1 49
2 46366 1 49
2 46367 1 49
2 46368 1 49
2 46369 1 49
2 46370 1 49
2 46371 1 49
2 46372 1 49
2 46373 1 49
2 46374 1 49
2 46375 1 49
2 46376 1 49
2 46377 1 49
2 46378 1 49
2 46379 1 49
2 46380 1 49
2 46381 1 49
2 46382 1 49
2 46383 1 49
2 46384 1 49
2 46385 1 49
2 46386 1 49
2 46387 1 49
2 46388 1 49
2 46389 1 49
2 46390 1 49
2 46391 1 49
2 46392 1 49
2 46393 1 49
2 46394 1 49
2 46395 1 49
2 46396 1 49
2 46397 1 49
2 46398 1 49
2 46399 1 49
2 46400 1 49
2 46401 1 49
2 46402 1 49
2 46403 1 49
2 46404 1 49
2 46405 1 49
2 46406 1 49
2 46407 1 49
2 46408 1 49
2 46409 1 49
2 46410 1 49
2 46411 1 49
2 46412 1 49
2 46413 1 49
2 46414 1 49
2 46415 1 49
2 46416 1 49
2 46417 1 49
2 46418 1 49
2 46419 1 49
2 46420 1 49
2 46421 1 49
2 46422 1 49
2 46423 1 49
2 46424 1 49
2 46425 1 49
2 46426 1 49
2 46427 1 49
2 46428 1 49
2 46429 1 49
2 46430 1 49
2 46431 1 49
2 46432 1 49
2 46433 1 49
2 46434 1 49
2 46435 1 49
2 46436 1 49
2 46437 1 49
2 46438 1 49
2 46439 1 49
2 46440 1 49
2 46441 1 49
2 46442 1 49
2 46443 1 49
2 46444 1 49
2 46445 1 50
2 46446 1 50
2 46447 1 50
2 46448 1 50
2 46449 1 50
2 46450 1 50
2 46451 1 50
2 46452 1 50
2 46453 1 50
2 46454 1 50
2 46455 1 50
2 46456 1 50
2 46457 1 50
2 46458 1 50
2 46459 1 50
2 46460 1 50
2 46461 1 50
2 46462 1 50
2 46463 1 50
2 46464 1 50
2 46465 1 50
2 46466 1 50
2 46467 1 50
2 46468 1 50
2 46469 1 50
2 46470 1 50
2 46471 1 50
2 46472 1 50
2 46473 1 50
2 46474 1 50
2 46475 1 50
2 46476 1 50
2 46477 1 50
2 46478 1 50
2 46479 1 50
2 46480 1 50
2 46481 1 50
2 46482 1 50
2 46483 1 50
2 46484 1 50
2 46485 1 50
2 46486 1 50
2 46487 1 50
2 46488 1 50
2 46489 1 50
2 46490 1 50
2 46491 1 50
2 46492 1 50
2 46493 1 50
2 46494 1 50
2 46495 1 50
2 46496 1 50
2 46497 1 50
2 46498 1 50
2 46499 1 50
2 46500 1 50
2 46501 1 50
2 46502 1 50
2 46503 1 50
2 46504 1 50
2 46505 1 50
2 46506 1 50
2 46507 1 50
2 46508 1 50
2 46509 1 50
2 46510 1 50
2 46511 1 50
2 46512 1 50
2 46513 1 50
2 46514 1 50
2 46515 1 50
2 46516 1 50
2 46517 1 50
2 46518 1 50
2 46519 1 50
2 46520 1 50
2 46521 1 50
2 46522 1 50
2 46523 1 50
2 46524 1 50
2 46525 1 50
2 46526 1 50
2 46527 1 50
2 46528 1 51
2 46529 1 51
2 46530 1 51
2 46531 1 51
2 46532 1 51
2 46533 1 51
2 46534 1 51
2 46535 1 51
2 46536 1 51
2 46537 1 51
2 46538 1 52
2 46539 1 52
2 46540 1 52
2 46541 1 52
2 46542 1 52
2 46543 1 52
2 46544 1 52
2 46545 1 52
2 46546 1 52
2 46547 1 52
2 46548 1 52
2 46549 1 52
2 46550 1 52
2 46551 1 52
2 46552 1 52
2 46553 1 54
2 46554 1 54
2 46555 1 54
2 46556 1 56
2 46557 1 56
2 46558 1 57
2 46559 1 57
2 46560 1 57
2 46561 1 57
2 46562 1 57
2 46563 1 57
2 46564 1 57
2 46565 1 57
2 46566 1 57
2 46567 1 57
2 46568 1 57
2 46569 1 57
2 46570 1 57
2 46571 1 57
2 46572 1 57
2 46573 1 57
2 46574 1 57
2 46575 1 57
2 46576 1 57
2 46577 1 57
2 46578 1 57
2 46579 1 57
2 46580 1 57
2 46581 1 57
2 46582 1 57
2 46583 1 57
2 46584 1 57
2 46585 1 57
2 46586 1 57
2 46587 1 57
2 46588 1 57
2 46589 1 57
2 46590 1 57
2 46591 1 57
2 46592 1 57
2 46593 1 57
2 46594 1 57
2 46595 1 57
2 46596 1 57
2 46597 1 57
2 46598 1 57
2 46599 1 57
2 46600 1 57
2 46601 1 57
2 46602 1 58
2 46603 1 58
2 46604 1 58
2 46605 1 58
2 46606 1 58
2 46607 1 58
2 46608 1 58
2 46609 1 58
2 46610 1 58
2 46611 1 58
2 46612 1 58
2 46613 1 58
2 46614 1 58
2 46615 1 58
2 46616 1 58
2 46617 1 58
2 46618 1 58
2 46619 1 58
2 46620 1 58
2 46621 1 58
2 46622 1 58
2 46623 1 58
2 46624 1 58
2 46625 1 58
2 46626 1 58
2 46627 1 58
2 46628 1 58
2 46629 1 58
2 46630 1 58
2 46631 1 58
2 46632 1 58
2 46633 1 58
2 46634 1 58
2 46635 1 58
2 46636 1 58
2 46637 1 58
2 46638 1 58
2 46639 1 58
2 46640 1 58
2 46641 1 58
2 46642 1 58
2 46643 1 58
2 46644 1 58
2 46645 1 59
2 46646 1 59
2 46647 1 59
2 46648 1 59
2 46649 1 59
2 46650 1 60
2 46651 1 60
2 46652 1 60
2 46653 1 60
2 46654 1 60
2 46655 1 60
2 46656 1 60
2 46657 1 60
2 46658 1 60
2 46659 1 60
2 46660 1 60
2 46661 1 60
2 46662 1 60
2 46663 1 60
2 46664 1 60
2 46665 1 60
2 46666 1 60
2 46667 1 60
2 46668 1 60
2 46669 1 60
2 46670 1 60
2 46671 1 60
2 46672 1 60
2 46673 1 60
2 46674 1 60
2 46675 1 60
2 46676 1 60
2 46677 1 60
2 46678 1 60
2 46679 1 60
2 46680 1 60
2 46681 1 60
2 46682 1 60
2 46683 1 60
2 46684 1 60
2 46685 1 60
2 46686 1 60
2 46687 1 60
2 46688 1 60
2 46689 1 60
2 46690 1 60
2 46691 1 60
2 46692 1 60
2 46693 1 60
2 46694 1 60
2 46695 1 60
2 46696 1 60
2 46697 1 60
2 46698 1 60
2 46699 1 60
2 46700 1 62
2 46701 1 62
2 46702 1 62
2 46703 1 62
2 46704 1 62
2 46705 1 62
2 46706 1 62
2 46707 1 62
2 46708 1 62
2 46709 1 62
2 46710 1 62
2 46711 1 62
2 46712 1 62
2 46713 1 62
2 46714 1 62
2 46715 1 62
2 46716 1 62
2 46717 1 62
2 46718 1 62
2 46719 1 62
2 46720 1 62
2 46721 1 62
2 46722 1 62
2 46723 1 62
2 46724 1 62
2 46725 1 63
2 46726 1 63
2 46727 1 63
2 46728 1 63
2 46729 1 63
2 46730 1 63
2 46731 1 63
2 46732 1 63
2 46733 1 63
2 46734 1 63
2 46735 1 63
2 46736 1 63
2 46737 1 63
2 46738 1 63
2 46739 1 63
2 46740 1 63
2 46741 1 63
2 46742 1 63
2 46743 1 63
2 46744 1 63
2 46745 1 63
2 46746 1 63
2 46747 1 63
2 46748 1 63
2 46749 1 63
2 46750 1 63
2 46751 1 63
2 46752 1 63
2 46753 1 63
2 46754 1 63
2 46755 1 63
2 46756 1 63
2 46757 1 63
2 46758 1 63
2 46759 1 63
2 46760 1 63
2 46761 1 63
2 46762 1 63
2 46763 1 63
2 46764 1 63
2 46765 1 63
2 46766 1 63
2 46767 1 63
2 46768 1 63
2 46769 1 63
2 46770 1 63
2 46771 1 63
2 46772 1 64
2 46773 1 64
2 46774 1 64
2 46775 1 65
2 46776 1 65
2 46777 1 65
2 46778 1 65
2 46779 1 65
2 46780 1 65
2 46781 1 66
2 46782 1 66
2 46783 1 66
2 46784 1 66
2 46785 1 66
2 46786 1 66
2 46787 1 66
2 46788 1 66
2 46789 1 66
2 46790 1 66
2 46791 1 66
2 46792 1 66
2 46793 1 66
2 46794 1 66
2 46795 1 66
2 46796 1 66
2 46797 1 66
2 46798 1 66
2 46799 1 66
2 46800 1 66
2 46801 1 66
2 46802 1 66
2 46803 1 66
2 46804 1 66
2 46805 1 66
2 46806 1 66
2 46807 1 66
2 46808 1 66
2 46809 1 66
2 46810 1 66
2 46811 1 66
2 46812 1 66
2 46813 1 66
2 46814 1 66
2 46815 1 66
2 46816 1 66
2 46817 1 66
2 46818 1 66
2 46819 1 66
2 46820 1 67
2 46821 1 67
2 46822 1 67
2 46823 1 67
2 46824 1 67
2 46825 1 67
2 46826 1 67
2 46827 1 67
2 46828 1 67
2 46829 1 67
2 46830 1 67
2 46831 1 67
2 46832 1 67
2 46833 1 67
2 46834 1 67
2 46835 1 67
2 46836 1 67
2 46837 1 67
2 46838 1 67
2 46839 1 67
2 46840 1 67
2 46841 1 67
2 46842 1 67
2 46843 1 67
2 46844 1 67
2 46845 1 67
2 46846 1 67
2 46847 1 67
2 46848 1 67
2 46849 1 67
2 46850 1 67
2 46851 1 67
2 46852 1 67
2 46853 1 67
2 46854 1 67
2 46855 1 68
2 46856 1 68
2 46857 1 68
2 46858 1 69
2 46859 1 69
2 46860 1 69
2 46861 1 69
2 46862 1 69
2 46863 1 69
2 46864 1 69
2 46865 1 70
2 46866 1 70
2 46867 1 72
2 46868 1 72
2 46869 1 72
2 46870 1 72
2 46871 1 72
2 46872 1 72
2 46873 1 72
2 46874 1 73
2 46875 1 73
2 46876 1 73
2 46877 1 73
2 46878 1 73
2 46879 1 73
2 46880 1 74
2 46881 1 74
2 46882 1 75
2 46883 1 75
2 46884 1 77
2 46885 1 77
2 46886 1 78
2 46887 1 78
2 46888 1 78
2 46889 1 78
2 46890 1 78
2 46891 1 78
2 46892 1 78
2 46893 1 78
2 46894 1 78
2 46895 1 78
2 46896 1 78
2 46897 1 79
2 46898 1 79
2 46899 1 79
2 46900 1 79
2 46901 1 80
2 46902 1 80
2 46903 1 80
2 46904 1 81
2 46905 1 81
2 46906 1 81
2 46907 1 82
2 46908 1 82
2 46909 1 83
2 46910 1 83
2 46911 1 83
2 46912 1 83
2 46913 1 85
2 46914 1 85
2 46915 1 86
2 46916 1 86
2 46917 1 86
2 46918 1 86
2 46919 1 86
2 46920 1 86
2 46921 1 86
2 46922 1 87
2 46923 1 87
2 46924 1 88
2 46925 1 88
2 46926 1 89
2 46927 1 89
2 46928 1 89
2 46929 1 89
2 46930 1 89
2 46931 1 92
2 46932 1 92
2 46933 1 92
2 46934 1 92
2 46935 1 95
2 46936 1 95
2 46937 1 97
2 46938 1 97
2 46939 1 98
2 46940 1 98
2 46941 1 98
2 46942 1 98
2 46943 1 98
2 46944 1 98
2 46945 1 99
2 46946 1 99
2 46947 1 100
2 46948 1 100
2 46949 1 100
2 46950 1 100
2 46951 1 100
2 46952 1 100
2 46953 1 100
2 46954 1 100
2 46955 1 101
2 46956 1 101
2 46957 1 101
2 46958 1 103
2 46959 1 103
2 46960 1 103
2 46961 1 103
2 46962 1 103
2 46963 1 103
2 46964 1 105
2 46965 1 105
2 46966 1 105
2 46967 1 105
2 46968 1 105
2 46969 1 106
2 46970 1 106
2 46971 1 106
2 46972 1 106
2 46973 1 106
2 46974 1 106
2 46975 1 106
2 46976 1 106
2 46977 1 106
2 46978 1 106
2 46979 1 106
2 46980 1 106
2 46981 1 106
2 46982 1 106
2 46983 1 106
2 46984 1 106
2 46985 1 106
2 46986 1 106
2 46987 1 107
2 46988 1 107
2 46989 1 107
2 46990 1 107
2 46991 1 107
2 46992 1 107
2 46993 1 118
2 46994 1 118
2 46995 1 118
2 46996 1 118
2 46997 1 118
2 46998 1 118
2 46999 1 118
2 47000 1 118
2 47001 1 118
2 47002 1 118
2 47003 1 118
2 47004 1 118
2 47005 1 118
2 47006 1 118
2 47007 1 118
2 47008 1 118
2 47009 1 118
2 47010 1 118
2 47011 1 118
2 47012 1 118
2 47013 1 118
2 47014 1 118
2 47015 1 118
2 47016 1 118
2 47017 1 118
2 47018 1 118
2 47019 1 118
2 47020 1 118
2 47021 1 118
2 47022 1 118
2 47023 1 118
2 47024 1 118
2 47025 1 118
2 47026 1 118
2 47027 1 119
2 47028 1 119
2 47029 1 119
2 47030 1 119
2 47031 1 119
2 47032 1 119
2 47033 1 119
2 47034 1 119
2 47035 1 119
2 47036 1 119
2 47037 1 119
2 47038 1 119
2 47039 1 119
2 47040 1 119
2 47041 1 119
2 47042 1 119
2 47043 1 119
2 47044 1 119
2 47045 1 119
2 47046 1 119
2 47047 1 119
2 47048 1 119
2 47049 1 119
2 47050 1 119
2 47051 1 119
2 47052 1 119
2 47053 1 119
2 47054 1 119
2 47055 1 119
2 47056 1 119
2 47057 1 119
2 47058 1 119
2 47059 1 119
2 47060 1 119
2 47061 1 119
2 47062 1 120
2 47063 1 120
2 47064 1 120
2 47065 1 121
2 47066 1 121
2 47067 1 121
2 47068 1 121
2 47069 1 121
2 47070 1 121
2 47071 1 121
2 47072 1 121
2 47073 1 121
2 47074 1 122
2 47075 1 122
2 47076 1 122
2 47077 1 122
2 47078 1 122
2 47079 1 122
2 47080 1 122
2 47081 1 122
2 47082 1 122
2 47083 1 122
2 47084 1 122
2 47085 1 122
2 47086 1 122
2 47087 1 122
2 47088 1 122
2 47089 1 122
2 47090 1 122
2 47091 1 122
2 47092 1 122
2 47093 1 122
2 47094 1 122
2 47095 1 122
2 47096 1 122
2 47097 1 122
2 47098 1 122
2 47099 1 122
2 47100 1 122
2 47101 1 122
2 47102 1 122
2 47103 1 122
2 47104 1 122
2 47105 1 122
2 47106 1 122
2 47107 1 123
2 47108 1 123
2 47109 1 123
2 47110 1 123
2 47111 1 123
2 47112 1 123
2 47113 1 123
2 47114 1 123
2 47115 1 123
2 47116 1 123
2 47117 1 123
2 47118 1 123
2 47119 1 123
2 47120 1 123
2 47121 1 123
2 47122 1 123
2 47123 1 123
2 47124 1 123
2 47125 1 123
2 47126 1 123
2 47127 1 123
2 47128 1 123
2 47129 1 123
2 47130 1 123
2 47131 1 123
2 47132 1 123
2 47133 1 123
2 47134 1 123
2 47135 1 123
2 47136 1 123
2 47137 1 123
2 47138 1 124
2 47139 1 124
2 47140 1 124
2 47141 1 125
2 47142 1 125
2 47143 1 125
2 47144 1 125
2 47145 1 125
2 47146 1 125
2 47147 1 125
2 47148 1 125
2 47149 1 125
2 47150 1 125
2 47151 1 125
2 47152 1 125
2 47153 1 125
2 47154 1 125
2 47155 1 125
2 47156 1 125
2 47157 1 125
2 47158 1 125
2 47159 1 127
2 47160 1 127
2 47161 1 132
2 47162 1 132
2 47163 1 132
2 47164 1 132
2 47165 1 133
2 47166 1 133
2 47167 1 133
2 47168 1 133
2 47169 1 133
2 47170 1 134
2 47171 1 134
2 47172 1 136
2 47173 1 136
2 47174 1 147
2 47175 1 147
2 47176 1 147
2 47177 1 149
2 47178 1 149
2 47179 1 149
2 47180 1 149
2 47181 1 149
2 47182 1 149
2 47183 1 149
2 47184 1 149
2 47185 1 149
2 47186 1 150
2 47187 1 150
2 47188 1 150
2 47189 1 150
2 47190 1 150
2 47191 1 151
2 47192 1 151
2 47193 1 151
2 47194 1 151
2 47195 1 151
2 47196 1 153
2 47197 1 153
2 47198 1 154
2 47199 1 154
2 47200 1 154
2 47201 1 155
2 47202 1 155
2 47203 1 155
2 47204 1 156
2 47205 1 156
2 47206 1 156
2 47207 1 156
2 47208 1 167
2 47209 1 167
2 47210 1 167
2 47211 1 167
2 47212 1 167
2 47213 1 167
2 47214 1 167
2 47215 1 167
2 47216 1 167
2 47217 1 167
2 47218 1 167
2 47219 1 167
2 47220 1 167
2 47221 1 167
2 47222 1 167
2 47223 1 167
2 47224 1 167
2 47225 1 167
2 47226 1 167
2 47227 1 167
2 47228 1 167
2 47229 1 167
2 47230 1 167
2 47231 1 167
2 47232 1 167
2 47233 1 167
2 47234 1 167
2 47235 1 167
2 47236 1 167
2 47237 1 167
2 47238 1 167
2 47239 1 168
2 47240 1 168
2 47241 1 168
2 47242 1 168
2 47243 1 168
2 47244 1 168
2 47245 1 168
2 47246 1 168
2 47247 1 168
2 47248 1 169
2 47249 1 169
2 47250 1 171
2 47251 1 171
2 47252 1 172
2 47253 1 172
2 47254 1 172
2 47255 1 172
2 47256 1 173
2 47257 1 173
2 47258 1 175
2 47259 1 175
2 47260 1 175
2 47261 1 175
2 47262 1 175
2 47263 1 175
2 47264 1 175
2 47265 1 175
2 47266 1 175
2 47267 1 175
2 47268 1 175
2 47269 1 175
2 47270 1 175
2 47271 1 175
2 47272 1 175
2 47273 1 175
2 47274 1 175
2 47275 1 175
2 47276 1 175
2 47277 1 175
2 47278 1 175
2 47279 1 175
2 47280 1 175
2 47281 1 175
2 47282 1 175
2 47283 1 175
2 47284 1 175
2 47285 1 175
2 47286 1 175
2 47287 1 175
2 47288 1 175
2 47289 1 175
2 47290 1 175
2 47291 1 175
2 47292 1 175
2 47293 1 175
2 47294 1 175
2 47295 1 175
2 47296 1 175
2 47297 1 175
2 47298 1 175
2 47299 1 175
2 47300 1 175
2 47301 1 175
2 47302 1 175
2 47303 1 175
2 47304 1 175
2 47305 1 176
2 47306 1 176
2 47307 1 176
2 47308 1 176
2 47309 1 176
2 47310 1 176
2 47311 1 176
2 47312 1 176
2 47313 1 176
2 47314 1 176
2 47315 1 176
2 47316 1 176
2 47317 1 176
2 47318 1 176
2 47319 1 176
2 47320 1 176
2 47321 1 176
2 47322 1 176
2 47323 1 176
2 47324 1 176
2 47325 1 176
2 47326 1 176
2 47327 1 176
2 47328 1 176
2 47329 1 176
2 47330 1 176
2 47331 1 176
2 47332 1 176
2 47333 1 176
2 47334 1 176
2 47335 1 176
2 47336 1 176
2 47337 1 176
2 47338 1 176
2 47339 1 176
2 47340 1 176
2 47341 1 176
2 47342 1 176
2 47343 1 176
2 47344 1 176
2 47345 1 176
2 47346 1 176
2 47347 1 176
2 47348 1 176
2 47349 1 176
2 47350 1 176
2 47351 1 176
2 47352 1 176
2 47353 1 176
2 47354 1 176
2 47355 1 176
2 47356 1 176
2 47357 1 176
2 47358 1 176
2 47359 1 176
2 47360 1 176
2 47361 1 176
2 47362 1 176
2 47363 1 176
2 47364 1 176
2 47365 1 176
2 47366 1 176
2 47367 1 176
2 47368 1 176
2 47369 1 176
2 47370 1 176
2 47371 1 177
2 47372 1 177
2 47373 1 177
2 47374 1 177
2 47375 1 177
2 47376 1 177
2 47377 1 177
2 47378 1 177
2 47379 1 177
2 47380 1 177
2 47381 1 177
2 47382 1 177
2 47383 1 177
2 47384 1 177
2 47385 1 177
2 47386 1 177
2 47387 1 177
2 47388 1 177
2 47389 1 177
2 47390 1 177
2 47391 1 177
2 47392 1 177
2 47393 1 177
2 47394 1 177
2 47395 1 177
2 47396 1 177
2 47397 1 177
2 47398 1 177
2 47399 1 177
2 47400 1 177
2 47401 1 177
2 47402 1 177
2 47403 1 177
2 47404 1 177
2 47405 1 177
2 47406 1 177
2 47407 1 177
2 47408 1 177
2 47409 1 177
2 47410 1 177
2 47411 1 177
2 47412 1 177
2 47413 1 177
2 47414 1 177
2 47415 1 177
2 47416 1 177
2 47417 1 177
2 47418 1 177
2 47419 1 177
2 47420 1 177
2 47421 1 177
2 47422 1 177
2 47423 1 177
2 47424 1 177
2 47425 1 177
2 47426 1 177
2 47427 1 177
2 47428 1 177
2 47429 1 177
2 47430 1 177
2 47431 1 177
2 47432 1 177
2 47433 1 177
2 47434 1 177
2 47435 1 177
2 47436 1 177
2 47437 1 177
2 47438 1 177
2 47439 1 177
2 47440 1 177
2 47441 1 177
2 47442 1 178
2 47443 1 178
2 47444 1 178
2 47445 1 178
2 47446 1 178
2 47447 1 178
2 47448 1 178
2 47449 1 178
2 47450 1 178
2 47451 1 178
2 47452 1 178
2 47453 1 178
2 47454 1 178
2 47455 1 178
2 47456 1 178
2 47457 1 178
2 47458 1 178
2 47459 1 178
2 47460 1 178
2 47461 1 178
2 47462 1 178
2 47463 1 178
2 47464 1 178
2 47465 1 178
2 47466 1 178
2 47467 1 178
2 47468 1 178
2 47469 1 178
2 47470 1 178
2 47471 1 178
2 47472 1 178
2 47473 1 178
2 47474 1 178
2 47475 1 178
2 47476 1 178
2 47477 1 178
2 47478 1 178
2 47479 1 178
2 47480 1 178
2 47481 1 178
2 47482 1 178
2 47483 1 178
2 47484 1 178
2 47485 1 178
2 47486 1 178
2 47487 1 178
2 47488 1 178
2 47489 1 178
2 47490 1 178
2 47491 1 178
2 47492 1 178
2 47493 1 178
2 47494 1 178
2 47495 1 178
2 47496 1 178
2 47497 1 178
2 47498 1 178
2 47499 1 178
2 47500 1 178
2 47501 1 178
2 47502 1 178
2 47503 1 178
2 47504 1 178
2 47505 1 178
2 47506 1 178
2 47507 1 178
2 47508 1 178
2 47509 1 178
2 47510 1 178
2 47511 1 179
2 47512 1 179
2 47513 1 179
2 47514 1 179
2 47515 1 179
2 47516 1 179
2 47517 1 179
2 47518 1 179
2 47519 1 179
2 47520 1 179
2 47521 1 179
2 47522 1 179
2 47523 1 179
2 47524 1 179
2 47525 1 179
2 47526 1 180
2 47527 1 180
2 47528 1 180
2 47529 1 180
2 47530 1 180
2 47531 1 180
2 47532 1 180
2 47533 1 180
2 47534 1 180
2 47535 1 180
2 47536 1 180
2 47537 1 180
2 47538 1 181
2 47539 1 181
2 47540 1 181
2 47541 1 181
2 47542 1 181
2 47543 1 182
2 47544 1 182
2 47545 1 182
2 47546 1 182
2 47547 1 182
2 47548 1 182
2 47549 1 182
2 47550 1 182
2 47551 1 182
2 47552 1 182
2 47553 1 182
2 47554 1 182
2 47555 1 182
2 47556 1 182
2 47557 1 182
2 47558 1 182
2 47559 1 182
2 47560 1 182
2 47561 1 182
2 47562 1 183
2 47563 1 183
2 47564 1 184
2 47565 1 184
2 47566 1 184
2 47567 1 184
2 47568 1 184
2 47569 1 184
2 47570 1 186
2 47571 1 186
2 47572 1 186
2 47573 1 186
2 47574 1 191
2 47575 1 191
2 47576 1 191
2 47577 1 191
2 47578 1 191
2 47579 1 191
2 47580 1 191
2 47581 1 191
2 47582 1 191
2 47583 1 191
2 47584 1 191
2 47585 1 191
2 47586 1 191
2 47587 1 191
2 47588 1 191
2 47589 1 191
2 47590 1 191
2 47591 1 191
2 47592 1 191
2 47593 1 191
2 47594 1 191
2 47595 1 191
2 47596 1 191
2 47597 1 191
2 47598 1 191
2 47599 1 191
2 47600 1 191
2 47601 1 191
2 47602 1 191
2 47603 1 191
2 47604 1 192
2 47605 1 192
2 47606 1 192
2 47607 1 192
2 47608 1 192
2 47609 1 192
2 47610 1 192
2 47611 1 192
2 47612 1 192
2 47613 1 192
2 47614 1 192
2 47615 1 192
2 47616 1 192
2 47617 1 192
2 47618 1 192
2 47619 1 192
2 47620 1 192
2 47621 1 192
2 47622 1 192
2 47623 1 192
2 47624 1 192
2 47625 1 192
2 47626 1 192
2 47627 1 192
2 47628 1 192
2 47629 1 192
2 47630 1 192
2 47631 1 192
2 47632 1 192
2 47633 1 192
2 47634 1 192
2 47635 1 192
2 47636 1 192
2 47637 1 192
2 47638 1 192
2 47639 1 192
2 47640 1 192
2 47641 1 192
2 47642 1 192
2 47643 1 192
2 47644 1 192
2 47645 1 192
2 47646 1 192
2 47647 1 192
2 47648 1 192
2 47649 1 192
2 47650 1 192
2 47651 1 192
2 47652 1 192
2 47653 1 192
2 47654 1 192
2 47655 1 192
2 47656 1 192
2 47657 1 192
2 47658 1 192
2 47659 1 192
2 47660 1 192
2 47661 1 192
2 47662 1 192
2 47663 1 192
2 47664 1 192
2 47665 1 192
2 47666 1 192
2 47667 1 192
2 47668 1 192
2 47669 1 192
2 47670 1 192
2 47671 1 192
2 47672 1 192
2 47673 1 192
2 47674 1 192
2 47675 1 192
2 47676 1 192
2 47677 1 192
2 47678 1 192
2 47679 1 192
2 47680 1 192
2 47681 1 192
2 47682 1 192
2 47683 1 192
2 47684 1 192
2 47685 1 192
2 47686 1 192
2 47687 1 192
2 47688 1 192
2 47689 1 192
2 47690 1 192
2 47691 1 193
2 47692 1 193
2 47693 1 193
2 47694 1 193
2 47695 1 193
2 47696 1 193
2 47697 1 193
2 47698 1 193
2 47699 1 193
2 47700 1 193
2 47701 1 193
2 47702 1 193
2 47703 1 193
2 47704 1 193
2 47705 1 193
2 47706 1 193
2 47707 1 193
2 47708 1 193
2 47709 1 193
2 47710 1 193
2 47711 1 193
2 47712 1 193
2 47713 1 193
2 47714 1 193
2 47715 1 193
2 47716 1 193
2 47717 1 193
2 47718 1 193
2 47719 1 193
2 47720 1 193
2 47721 1 193
2 47722 1 193
2 47723 1 193
2 47724 1 193
2 47725 1 193
2 47726 1 193
2 47727 1 193
2 47728 1 193
2 47729 1 193
2 47730 1 193
2 47731 1 193
2 47732 1 193
2 47733 1 193
2 47734 1 193
2 47735 1 193
2 47736 1 193
2 47737 1 193
2 47738 1 193
2 47739 1 193
2 47740 1 193
2 47741 1 193
2 47742 1 193
2 47743 1 193
2 47744 1 193
2 47745 1 193
2 47746 1 193
2 47747 1 193
2 47748 1 193
2 47749 1 193
2 47750 1 194
2 47751 1 194
2 47752 1 194
2 47753 1 194
2 47754 1 194
2 47755 1 194
2 47756 1 194
2 47757 1 194
2 47758 1 194
2 47759 1 194
2 47760 1 194
2 47761 1 194
2 47762 1 194
2 47763 1 194
2 47764 1 194
2 47765 1 194
2 47766 1 194
2 47767 1 194
2 47768 1 194
2 47769 1 194
2 47770 1 194
2 47771 1 194
2 47772 1 194
2 47773 1 194
2 47774 1 194
2 47775 1 194
2 47776 1 194
2 47777 1 194
2 47778 1 194
2 47779 1 194
2 47780 1 194
2 47781 1 194
2 47782 1 194
2 47783 1 194
2 47784 1 194
2 47785 1 194
2 47786 1 194
2 47787 1 194
2 47788 1 194
2 47789 1 194
2 47790 1 194
2 47791 1 194
2 47792 1 194
2 47793 1 194
2 47794 1 194
2 47795 1 194
2 47796 1 194
2 47797 1 194
2 47798 1 194
2 47799 1 194
2 47800 1 194
2 47801 1 194
2 47802 1 194
2 47803 1 194
2 47804 1 194
2 47805 1 194
2 47806 1 194
2 47807 1 194
2 47808 1 194
2 47809 1 194
2 47810 1 194
2 47811 1 194
2 47812 1 194
2 47813 1 194
2 47814 1 194
2 47815 1 194
2 47816 1 194
2 47817 1 194
2 47818 1 194
2 47819 1 194
2 47820 1 194
2 47821 1 194
2 47822 1 194
2 47823 1 194
2 47824 1 194
2 47825 1 194
2 47826 1 194
2 47827 1 194
2 47828 1 194
2 47829 1 194
2 47830 1 194
2 47831 1 194
2 47832 1 196
2 47833 1 196
2 47834 1 196
2 47835 1 197
2 47836 1 197
2 47837 1 197
2 47838 1 197
2 47839 1 200
2 47840 1 200
2 47841 1 201
2 47842 1 201
2 47843 1 215
2 47844 1 215
2 47845 1 215
2 47846 1 215
2 47847 1 215
2 47848 1 215
2 47849 1 215
2 47850 1 215
2 47851 1 215
2 47852 1 215
2 47853 1 215
2 47854 1 217
2 47855 1 217
2 47856 1 217
2 47857 1 217
2 47858 1 217
2 47859 1 217
2 47860 1 217
2 47861 1 217
2 47862 1 219
2 47863 1 219
2 47864 1 220
2 47865 1 220
2 47866 1 220
2 47867 1 227
2 47868 1 227
2 47869 1 227
2 47870 1 233
2 47871 1 233
2 47872 1 233
2 47873 1 233
2 47874 1 233
2 47875 1 233
2 47876 1 233
2 47877 1 233
2 47878 1 233
2 47879 1 233
2 47880 1 233
2 47881 1 235
2 47882 1 235
2 47883 1 235
2 47884 1 235
2 47885 1 236
2 47886 1 236
2 47887 1 236
2 47888 1 246
2 47889 1 246
2 47890 1 246
2 47891 1 246
2 47892 1 246
2 47893 1 246
2 47894 1 246
2 47895 1 247
2 47896 1 247
2 47897 1 247
2 47898 1 247
2 47899 1 247
2 47900 1 247
2 47901 1 248
2 47902 1 248
2 47903 1 248
2 47904 1 248
2 47905 1 248
2 47906 1 248
2 47907 1 248
2 47908 1 248
2 47909 1 248
2 47910 1 248
2 47911 1 248
2 47912 1 248
2 47913 1 248
2 47914 1 248
2 47915 1 248
2 47916 1 248
2 47917 1 248
2 47918 1 248
2 47919 1 248
2 47920 1 248
2 47921 1 248
2 47922 1 248
2 47923 1 248
2 47924 1 248
2 47925 1 249
2 47926 1 249
2 47927 1 251
2 47928 1 251
2 47929 1 251
2 47930 1 251
2 47931 1 251
2 47932 1 251
2 47933 1 251
2 47934 1 251
2 47935 1 251
2 47936 1 251
2 47937 1 251
2 47938 1 252
2 47939 1 252
2 47940 1 252
2 47941 1 253
2 47942 1 253
2 47943 1 253
2 47944 1 253
2 47945 1 255
2 47946 1 255
2 47947 1 255
2 47948 1 255
2 47949 1 255
2 47950 1 255
2 47951 1 255
2 47952 1 256
2 47953 1 256
2 47954 1 256
2 47955 1 256
2 47956 1 256
2 47957 1 256
2 47958 1 256
2 47959 1 256
2 47960 1 256
2 47961 1 256
2 47962 1 266
2 47963 1 266
2 47964 1 266
2 47965 1 266
2 47966 1 266
2 47967 1 266
2 47968 1 266
2 47969 1 266
2 47970 1 266
2 47971 1 266
2 47972 1 266
2 47973 1 266
2 47974 1 266
2 47975 1 266
2 47976 1 266
2 47977 1 266
2 47978 1 266
2 47979 1 267
2 47980 1 267
2 47981 1 268
2 47982 1 268
2 47983 1 270
2 47984 1 270
2 47985 1 270
2 47986 1 271
2 47987 1 271
2 47988 1 271
2 47989 1 271
2 47990 1 271
2 47991 1 271
2 47992 1 271
2 47993 1 271
2 47994 1 271
2 47995 1 271
2 47996 1 271
2 47997 1 271
2 47998 1 271
2 47999 1 272
2 48000 1 272
2 48001 1 272
2 48002 1 273
2 48003 1 273
2 48004 1 273
2 48005 1 273
2 48006 1 273
2 48007 1 273
2 48008 1 273
2 48009 1 273
2 48010 1 273
2 48011 1 273
2 48012 1 275
2 48013 1 275
2 48014 1 276
2 48015 1 276
2 48016 1 277
2 48017 1 277
2 48018 1 280
2 48019 1 280
2 48020 1 280
2 48021 1 287
2 48022 1 287
2 48023 1 287
2 48024 1 287
2 48025 1 287
2 48026 1 288
2 48027 1 288
2 48028 1 288
2 48029 1 288
2 48030 1 288
2 48031 1 288
2 48032 1 289
2 48033 1 289
2 48034 1 290
2 48035 1 290
2 48036 1 290
2 48037 1 291
2 48038 1 291
2 48039 1 292
2 48040 1 292
2 48041 1 294
2 48042 1 294
2 48043 1 296
2 48044 1 296
2 48045 1 297
2 48046 1 297
2 48047 1 297
2 48048 1 297
2 48049 1 297
2 48050 1 297
2 48051 1 297
2 48052 1 297
2 48053 1 297
2 48054 1 297
2 48055 1 297
2 48056 1 297
2 48057 1 297
2 48058 1 297
2 48059 1 297
2 48060 1 297
2 48061 1 297
2 48062 1 297
2 48063 1 297
2 48064 1 297
2 48065 1 297
2 48066 1 297
2 48067 1 297
2 48068 1 297
2 48069 1 297
2 48070 1 297
2 48071 1 297
2 48072 1 297
2 48073 1 297
2 48074 1 297
2 48075 1 297
2 48076 1 297
2 48077 1 297
2 48078 1 297
2 48079 1 297
2 48080 1 297
2 48081 1 297
2 48082 1 297
2 48083 1 297
2 48084 1 297
2 48085 1 297
2 48086 1 297
2 48087 1 298
2 48088 1 298
2 48089 1 299
2 48090 1 299
2 48091 1 299
2 48092 1 299
2 48093 1 299
2 48094 1 299
2 48095 1 299
2 48096 1 299
2 48097 1 299
2 48098 1 299
2 48099 1 299
2 48100 1 299
2 48101 1 299
2 48102 1 299
2 48103 1 299
2 48104 1 299
2 48105 1 299
2 48106 1 299
2 48107 1 299
2 48108 1 299
2 48109 1 299
2 48110 1 299
2 48111 1 299
2 48112 1 299
2 48113 1 299
2 48114 1 299
2 48115 1 299
2 48116 1 299
2 48117 1 299
2 48118 1 299
2 48119 1 299
2 48120 1 299
2 48121 1 299
2 48122 1 299
2 48123 1 299
2 48124 1 299
2 48125 1 299
2 48126 1 299
2 48127 1 299
2 48128 1 299
2 48129 1 299
2 48130 1 299
2 48131 1 299
2 48132 1 299
2 48133 1 299
2 48134 1 299
2 48135 1 299
2 48136 1 300
2 48137 1 300
2 48138 1 300
2 48139 1 300
2 48140 1 307
2 48141 1 307
2 48142 1 307
2 48143 1 307
2 48144 1 307
2 48145 1 307
2 48146 1 308
2 48147 1 308
2 48148 1 309
2 48149 1 309
2 48150 1 312
2 48151 1 312
2 48152 1 312
2 48153 1 312
2 48154 1 312
2 48155 1 312
2 48156 1 312
2 48157 1 312
2 48158 1 312
2 48159 1 312
2 48160 1 312
2 48161 1 312
2 48162 1 312
2 48163 1 312
2 48164 1 312
2 48165 1 312
2 48166 1 312
2 48167 1 312
2 48168 1 312
2 48169 1 312
2 48170 1 312
2 48171 1 312
2 48172 1 313
2 48173 1 313
2 48174 1 313
2 48175 1 313
2 48176 1 313
2 48177 1 313
2 48178 1 314
2 48179 1 314
2 48180 1 314
2 48181 1 314
2 48182 1 315
2 48183 1 315
2 48184 1 315
2 48185 1 315
2 48186 1 316
2 48187 1 316
2 48188 1 316
2 48189 1 316
2 48190 1 316
2 48191 1 316
2 48192 1 316
2 48193 1 317
2 48194 1 317
2 48195 1 317
2 48196 1 317
2 48197 1 318
2 48198 1 318
2 48199 1 318
2 48200 1 318
2 48201 1 318
2 48202 1 318
2 48203 1 318
2 48204 1 318
2 48205 1 318
2 48206 1 318
2 48207 1 318
2 48208 1 318
2 48209 1 318
2 48210 1 318
2 48211 1 318
2 48212 1 318
2 48213 1 318
2 48214 1 318
2 48215 1 318
2 48216 1 318
2 48217 1 318
2 48218 1 318
2 48219 1 318
2 48220 1 318
2 48221 1 318
2 48222 1 318
2 48223 1 318
2 48224 1 318
2 48225 1 318
2 48226 1 318
2 48227 1 318
2 48228 1 318
2 48229 1 318
2 48230 1 318
2 48231 1 318
2 48232 1 318
2 48233 1 318
2 48234 1 318
2 48235 1 318
2 48236 1 318
2 48237 1 318
2 48238 1 318
2 48239 1 318
2 48240 1 318
2 48241 1 318
2 48242 1 318
2 48243 1 318
2 48244 1 318
2 48245 1 318
2 48246 1 318
2 48247 1 319
2 48248 1 319
2 48249 1 319
2 48250 1 319
2 48251 1 319
2 48252 1 319
2 48253 1 319
2 48254 1 319
2 48255 1 319
2 48256 1 319
2 48257 1 322
2 48258 1 322
2 48259 1 322
2 48260 1 322
2 48261 1 322
2 48262 1 322
2 48263 1 322
2 48264 1 322
2 48265 1 322
2 48266 1 322
2 48267 1 322
2 48268 1 322
2 48269 1 322
2 48270 1 322
2 48271 1 322
2 48272 1 322
2 48273 1 322
2 48274 1 322
2 48275 1 322
2 48276 1 322
2 48277 1 322
2 48278 1 322
2 48279 1 322
2 48280 1 322
2 48281 1 322
2 48282 1 322
2 48283 1 322
2 48284 1 322
2 48285 1 322
2 48286 1 322
2 48287 1 322
2 48288 1 322
2 48289 1 322
2 48290 1 322
2 48291 1 324
2 48292 1 324
2 48293 1 325
2 48294 1 325
2 48295 1 325
2 48296 1 325
2 48297 1 325
2 48298 1 325
2 48299 1 325
2 48300 1 330
2 48301 1 330
2 48302 1 330
2 48303 1 330
2 48304 1 330
2 48305 1 330
2 48306 1 330
2 48307 1 330
2 48308 1 330
2 48309 1 333
2 48310 1 333
2 48311 1 333
2 48312 1 333
2 48313 1 333
2 48314 1 333
2 48315 1 333
2 48316 1 335
2 48317 1 335
2 48318 1 335
2 48319 1 335
2 48320 1 336
2 48321 1 336
2 48322 1 336
2 48323 1 336
2 48324 1 336
2 48325 1 336
2 48326 1 336
2 48327 1 336
2 48328 1 336
2 48329 1 336
2 48330 1 348
2 48331 1 348
2 48332 1 348
2 48333 1 348
2 48334 1 348
2 48335 1 348
2 48336 1 348
2 48337 1 348
2 48338 1 348
2 48339 1 348
2 48340 1 348
2 48341 1 348
2 48342 1 348
2 48343 1 348
2 48344 1 348
2 48345 1 348
2 48346 1 348
2 48347 1 349
2 48348 1 349
2 48349 1 349
2 48350 1 350
2 48351 1 350
2 48352 1 350
2 48353 1 350
2 48354 1 351
2 48355 1 351
2 48356 1 351
2 48357 1 351
2 48358 1 351
2 48359 1 351
2 48360 1 351
2 48361 1 351
2 48362 1 351
2 48363 1 351
2 48364 1 360
2 48365 1 360
2 48366 1 360
2 48367 1 360
2 48368 1 360
2 48369 1 360
2 48370 1 360
2 48371 1 360
2 48372 1 360
2 48373 1 360
2 48374 1 360
2 48375 1 360
2 48376 1 360
2 48377 1 360
2 48378 1 360
2 48379 1 360
2 48380 1 361
2 48381 1 361
2 48382 1 361
2 48383 1 361
2 48384 1 361
2 48385 1 362
2 48386 1 362
2 48387 1 362
2 48388 1 362
2 48389 1 362
2 48390 1 362
2 48391 1 362
2 48392 1 362
2 48393 1 362
2 48394 1 363
2 48395 1 363
2 48396 1 371
2 48397 1 371
2 48398 1 371
2 48399 1 371
2 48400 1 371
2 48401 1 371
2 48402 1 371
2 48403 1 371
2 48404 1 371
2 48405 1 371
2 48406 1 371
2 48407 1 372
2 48408 1 372
2 48409 1 373
2 48410 1 373
2 48411 1 374
2 48412 1 374
2 48413 1 374
2 48414 1 375
2 48415 1 375
2 48416 1 375
2 48417 1 376
2 48418 1 376
2 48419 1 383
2 48420 1 383
2 48421 1 383
2 48422 1 383
2 48423 1 384
2 48424 1 384
2 48425 1 397
2 48426 1 397
2 48427 1 397
2 48428 1 397
2 48429 1 397
2 48430 1 397
2 48431 1 397
2 48432 1 397
2 48433 1 397
2 48434 1 397
2 48435 1 397
2 48436 1 397
2 48437 1 397
2 48438 1 397
2 48439 1 397
2 48440 1 397
2 48441 1 397
2 48442 1 397
2 48443 1 397
2 48444 1 397
2 48445 1 397
2 48446 1 397
2 48447 1 398
2 48448 1 398
2 48449 1 399
2 48450 1 399
2 48451 1 400
2 48452 1 400
2 48453 1 400
2 48454 1 400
2 48455 1 400
2 48456 1 400
2 48457 1 400
2 48458 1 400
2 48459 1 400
2 48460 1 400
2 48461 1 400
2 48462 1 400
2 48463 1 400
2 48464 1 400
2 48465 1 400
2 48466 1 400
2 48467 1 400
2 48468 1 400
2 48469 1 400
2 48470 1 400
2 48471 1 400
2 48472 1 400
2 48473 1 400
2 48474 1 400
2 48475 1 400
2 48476 1 400
2 48477 1 400
2 48478 1 400
2 48479 1 400
2 48480 1 400
2 48481 1 400
2 48482 1 400
2 48483 1 400
2 48484 1 400
2 48485 1 400
2 48486 1 400
2 48487 1 400
2 48488 1 400
2 48489 1 400
2 48490 1 400
2 48491 1 400
2 48492 1 400
2 48493 1 400
2 48494 1 400
2 48495 1 400
2 48496 1 400
2 48497 1 400
2 48498 1 400
2 48499 1 400
2 48500 1 400
2 48501 1 400
2 48502 1 400
2 48503 1 400
2 48504 1 400
2 48505 1 400
2 48506 1 400
2 48507 1 400
2 48508 1 400
2 48509 1 400
2 48510 1 400
2 48511 1 400
2 48512 1 400
2 48513 1 400
2 48514 1 400
2 48515 1 400
2 48516 1 400
2 48517 1 400
2 48518 1 400
2 48519 1 400
2 48520 1 400
2 48521 1 400
2 48522 1 400
2 48523 1 400
2 48524 1 400
2 48525 1 400
2 48526 1 400
2 48527 1 400
2 48528 1 400
2 48529 1 401
2 48530 1 401
2 48531 1 401
2 48532 1 401
2 48533 1 401
2 48534 1 401
2 48535 1 401
2 48536 1 401
2 48537 1 401
2 48538 1 401
2 48539 1 401
2 48540 1 401
2 48541 1 401
2 48542 1 401
2 48543 1 401
2 48544 1 401
2 48545 1 401
2 48546 1 401
2 48547 1 401
2 48548 1 401
2 48549 1 401
2 48550 1 401
2 48551 1 401
2 48552 1 401
2 48553 1 401
2 48554 1 401
2 48555 1 401
2 48556 1 401
2 48557 1 401
2 48558 1 401
2 48559 1 401
2 48560 1 401
2 48561 1 401
2 48562 1 401
2 48563 1 401
2 48564 1 401
2 48565 1 401
2 48566 1 402
2 48567 1 402
2 48568 1 402
2 48569 1 402
2 48570 1 402
2 48571 1 402
2 48572 1 402
2 48573 1 402
2 48574 1 402
2 48575 1 402
2 48576 1 402
2 48577 1 402
2 48578 1 402
2 48579 1 402
2 48580 1 402
2 48581 1 402
2 48582 1 402
2 48583 1 402
2 48584 1 402
2 48585 1 402
2 48586 1 402
2 48587 1 402
2 48588 1 402
2 48589 1 402
2 48590 1 402
2 48591 1 402
2 48592 1 402
2 48593 1 402
2 48594 1 402
2 48595 1 402
2 48596 1 404
2 48597 1 404
2 48598 1 411
2 48599 1 411
2 48600 1 411
2 48601 1 411
2 48602 1 411
2 48603 1 411
2 48604 1 411
2 48605 1 411
2 48606 1 411
2 48607 1 413
2 48608 1 413
2 48609 1 413
2 48610 1 413
2 48611 1 413
2 48612 1 413
2 48613 1 413
2 48614 1 413
2 48615 1 413
2 48616 1 413
2 48617 1 413
2 48618 1 413
2 48619 1 413
2 48620 1 414
2 48621 1 414
2 48622 1 414
2 48623 1 414
2 48624 1 414
2 48625 1 414
2 48626 1 414
2 48627 1 414
2 48628 1 414
2 48629 1 414
2 48630 1 414
2 48631 1 414
2 48632 1 414
2 48633 1 414
2 48634 1 414
2 48635 1 414
2 48636 1 414
2 48637 1 414
2 48638 1 414
2 48639 1 414
2 48640 1 414
2 48641 1 414
2 48642 1 415
2 48643 1 415
2 48644 1 415
2 48645 1 415
2 48646 1 415
2 48647 1 415
2 48648 1 415
2 48649 1 415
2 48650 1 415
2 48651 1 415
2 48652 1 415
2 48653 1 415
2 48654 1 415
2 48655 1 415
2 48656 1 415
2 48657 1 415
2 48658 1 415
2 48659 1 415
2 48660 1 415
2 48661 1 415
2 48662 1 415
2 48663 1 415
2 48664 1 415
2 48665 1 415
2 48666 1 415
2 48667 1 415
2 48668 1 415
2 48669 1 415
2 48670 1 415
2 48671 1 415
2 48672 1 415
2 48673 1 415
2 48674 1 415
2 48675 1 415
2 48676 1 415
2 48677 1 415
2 48678 1 415
2 48679 1 415
2 48680 1 415
2 48681 1 415
2 48682 1 415
2 48683 1 415
2 48684 1 415
2 48685 1 415
2 48686 1 415
2 48687 1 415
2 48688 1 415
2 48689 1 415
2 48690 1 415
2 48691 1 415
2 48692 1 415
2 48693 1 415
2 48694 1 415
2 48695 1 415
2 48696 1 415
2 48697 1 415
2 48698 1 415
2 48699 1 415
2 48700 1 415
2 48701 1 415
2 48702 1 415
2 48703 1 415
2 48704 1 415
2 48705 1 415
2 48706 1 415
2 48707 1 415
2 48708 1 415
2 48709 1 415
2 48710 1 415
2 48711 1 415
2 48712 1 416
2 48713 1 416
2 48714 1 416
2 48715 1 416
2 48716 1 416
2 48717 1 416
2 48718 1 416
2 48719 1 416
2 48720 1 416
2 48721 1 416
2 48722 1 416
2 48723 1 416
2 48724 1 416
2 48725 1 416
2 48726 1 416
2 48727 1 416
2 48728 1 416
2 48729 1 416
2 48730 1 416
2 48731 1 416
2 48732 1 416
2 48733 1 416
2 48734 1 416
2 48735 1 416
2 48736 1 416
2 48737 1 416
2 48738 1 416
2 48739 1 416
2 48740 1 416
2 48741 1 416
2 48742 1 416
2 48743 1 416
2 48744 1 416
2 48745 1 416
2 48746 1 416
2 48747 1 416
2 48748 1 416
2 48749 1 416
2 48750 1 416
2 48751 1 416
2 48752 1 416
2 48753 1 416
2 48754 1 416
2 48755 1 416
2 48756 1 416
2 48757 1 416
2 48758 1 416
2 48759 1 416
2 48760 1 416
2 48761 1 416
2 48762 1 416
2 48763 1 416
2 48764 1 416
2 48765 1 416
2 48766 1 416
2 48767 1 416
2 48768 1 416
2 48769 1 416
2 48770 1 416
2 48771 1 416
2 48772 1 416
2 48773 1 416
2 48774 1 416
2 48775 1 417
2 48776 1 417
2 48777 1 417
2 48778 1 417
2 48779 1 417
2 48780 1 417
2 48781 1 417
2 48782 1 417
2 48783 1 417
2 48784 1 417
2 48785 1 418
2 48786 1 418
2 48787 1 418
2 48788 1 418
2 48789 1 419
2 48790 1 419
2 48791 1 420
2 48792 1 420
2 48793 1 423
2 48794 1 423
2 48795 1 423
2 48796 1 424
2 48797 1 424
2 48798 1 428
2 48799 1 428
2 48800 1 428
2 48801 1 428
2 48802 1 428
2 48803 1 429
2 48804 1 429
2 48805 1 429
2 48806 1 429
2 48807 1 429
2 48808 1 429
2 48809 1 429
2 48810 1 429
2 48811 1 429
2 48812 1 429
2 48813 1 429
2 48814 1 429
2 48815 1 429
2 48816 1 429
2 48817 1 429
2 48818 1 429
2 48819 1 429
2 48820 1 429
2 48821 1 429
2 48822 1 429
2 48823 1 429
2 48824 1 429
2 48825 1 429
2 48826 1 429
2 48827 1 429
2 48828 1 429
2 48829 1 429
2 48830 1 429
2 48831 1 429
2 48832 1 429
2 48833 1 429
2 48834 1 429
2 48835 1 429
2 48836 1 429
2 48837 1 429
2 48838 1 429
2 48839 1 429
2 48840 1 429
2 48841 1 429
2 48842 1 429
2 48843 1 430
2 48844 1 430
2 48845 1 430
2 48846 1 430
2 48847 1 430
2 48848 1 430
2 48849 1 430
2 48850 1 430
2 48851 1 430
2 48852 1 430
2 48853 1 430
2 48854 1 430
2 48855 1 430
2 48856 1 430
2 48857 1 430
2 48858 1 430
2 48859 1 430
2 48860 1 430
2 48861 1 430
2 48862 1 430
2 48863 1 430
2 48864 1 430
2 48865 1 431
2 48866 1 431
2 48867 1 431
2 48868 1 431
2 48869 1 431
2 48870 1 431
2 48871 1 432
2 48872 1 432
2 48873 1 432
2 48874 1 432
2 48875 1 432
2 48876 1 432
2 48877 1 432
2 48878 1 432
2 48879 1 432
2 48880 1 433
2 48881 1 433
2 48882 1 433
2 48883 1 433
2 48884 1 433
2 48885 1 440
2 48886 1 440
2 48887 1 440
2 48888 1 440
2 48889 1 440
2 48890 1 440
2 48891 1 440
2 48892 1 440
2 48893 1 440
2 48894 1 440
2 48895 1 440
2 48896 1 440
2 48897 1 440
2 48898 1 440
2 48899 1 440
2 48900 1 440
2 48901 1 440
2 48902 1 440
2 48903 1 440
2 48904 1 440
2 48905 1 440
2 48906 1 440
2 48907 1 440
2 48908 1 440
2 48909 1 440
2 48910 1 440
2 48911 1 440
2 48912 1 440
2 48913 1 440
2 48914 1 440
2 48915 1 440
2 48916 1 440
2 48917 1 440
2 48918 1 440
2 48919 1 440
2 48920 1 440
2 48921 1 440
2 48922 1 440
2 48923 1 440
2 48924 1 440
2 48925 1 440
2 48926 1 440
2 48927 1 440
2 48928 1 440
2 48929 1 440
2 48930 1 440
2 48931 1 440
2 48932 1 440
2 48933 1 440
2 48934 1 440
2 48935 1 440
2 48936 1 440
2 48937 1 440
2 48938 1 440
2 48939 1 440
2 48940 1 440
2 48941 1 440
2 48942 1 440
2 48943 1 440
2 48944 1 440
2 48945 1 440
2 48946 1 440
2 48947 1 440
2 48948 1 440
2 48949 1 441
2 48950 1 441
2 48951 1 442
2 48952 1 442
2 48953 1 442
2 48954 1 442
2 48955 1 442
2 48956 1 442
2 48957 1 442
2 48958 1 442
2 48959 1 442
2 48960 1 442
2 48961 1 442
2 48962 1 442
2 48963 1 442
2 48964 1 442
2 48965 1 442
2 48966 1 442
2 48967 1 442
2 48968 1 442
2 48969 1 442
2 48970 1 442
2 48971 1 442
2 48972 1 443
2 48973 1 443
2 48974 1 446
2 48975 1 446
2 48976 1 446
2 48977 1 446
2 48978 1 446
2 48979 1 446
2 48980 1 448
2 48981 1 448
2 48982 1 448
2 48983 1 448
2 48984 1 448
2 48985 1 448
2 48986 1 448
2 48987 1 448
2 48988 1 448
2 48989 1 450
2 48990 1 450
2 48991 1 451
2 48992 1 451
2 48993 1 451
2 48994 1 451
2 48995 1 451
2 48996 1 451
2 48997 1 451
2 48998 1 451
2 48999 1 451
2 49000 1 451
2 49001 1 451
2 49002 1 451
2 49003 1 451
2 49004 1 451
2 49005 1 451
2 49006 1 451
2 49007 1 451
2 49008 1 451
2 49009 1 451
2 49010 1 451
2 49011 1 451
2 49012 1 451
2 49013 1 451
2 49014 1 451
2 49015 1 451
2 49016 1 451
2 49017 1 451
2 49018 1 451
2 49019 1 451
2 49020 1 451
2 49021 1 451
2 49022 1 451
2 49023 1 451
2 49024 1 451
2 49025 1 451
2 49026 1 451
2 49027 1 451
2 49028 1 451
2 49029 1 451
2 49030 1 451
2 49031 1 451
2 49032 1 451
2 49033 1 451
2 49034 1 451
2 49035 1 451
2 49036 1 451
2 49037 1 451
2 49038 1 451
2 49039 1 451
2 49040 1 451
2 49041 1 451
2 49042 1 451
2 49043 1 451
2 49044 1 451
2 49045 1 451
2 49046 1 451
2 49047 1 451
2 49048 1 451
2 49049 1 451
2 49050 1 451
2 49051 1 451
2 49052 1 451
2 49053 1 451
2 49054 1 451
2 49055 1 451
2 49056 1 451
2 49057 1 451
2 49058 1 451
2 49059 1 451
2 49060 1 451
2 49061 1 451
2 49062 1 451
2 49063 1 451
2 49064 1 451
2 49065 1 451
2 49066 1 451
2 49067 1 451
2 49068 1 452
2 49069 1 452
2 49070 1 452
2 49071 1 452
2 49072 1 452
2 49073 1 452
2 49074 1 452
2 49075 1 452
2 49076 1 452
2 49077 1 452
2 49078 1 452
2 49079 1 452
2 49080 1 452
2 49081 1 452
2 49082 1 452
2 49083 1 452
2 49084 1 452
2 49085 1 452
2 49086 1 452
2 49087 1 452
2 49088 1 452
2 49089 1 452
2 49090 1 452
2 49091 1 452
2 49092 1 452
2 49093 1 452
2 49094 1 452
2 49095 1 452
2 49096 1 452
2 49097 1 453
2 49098 1 453
2 49099 1 459
2 49100 1 459
2 49101 1 460
2 49102 1 460
2 49103 1 460
2 49104 1 460
2 49105 1 460
2 49106 1 460
2 49107 1 460
2 49108 1 460
2 49109 1 460
2 49110 1 460
2 49111 1 460
2 49112 1 460
2 49113 1 460
2 49114 1 460
2 49115 1 460
2 49116 1 460
2 49117 1 460
2 49118 1 460
2 49119 1 460
2 49120 1 460
2 49121 1 460
2 49122 1 460
2 49123 1 460
2 49124 1 461
2 49125 1 461
2 49126 1 461
2 49127 1 461
2 49128 1 461
2 49129 1 461
2 49130 1 461
2 49131 1 461
2 49132 1 470
2 49133 1 470
2 49134 1 470
2 49135 1 470
2 49136 1 470
2 49137 1 470
2 49138 1 471
2 49139 1 471
2 49140 1 471
2 49141 1 472
2 49142 1 472
2 49143 1 472
2 49144 1 472
2 49145 1 472
2 49146 1 472
2 49147 1 474
2 49148 1 474
2 49149 1 474
2 49150 1 474
2 49151 1 474
2 49152 1 476
2 49153 1 476
2 49154 1 476
2 49155 1 477
2 49156 1 477
2 49157 1 477
2 49158 1 478
2 49159 1 478
2 49160 1 478
2 49161 1 478
2 49162 1 478
2 49163 1 478
2 49164 1 478
2 49165 1 478
2 49166 1 478
2 49167 1 478
2 49168 1 478
2 49169 1 480
2 49170 1 480
2 49171 1 480
2 49172 1 480
2 49173 1 480
2 49174 1 481
2 49175 1 481
2 49176 1 481
2 49177 1 481
2 49178 1 481
2 49179 1 481
2 49180 1 481
2 49181 1 481
2 49182 1 481
2 49183 1 481
2 49184 1 481
2 49185 1 481
2 49186 1 481
2 49187 1 481
2 49188 1 481
2 49189 1 481
2 49190 1 481
2 49191 1 481
2 49192 1 481
2 49193 1 481
2 49194 1 481
2 49195 1 481
2 49196 1 481
2 49197 1 481
2 49198 1 481
2 49199 1 481
2 49200 1 481
2 49201 1 481
2 49202 1 481
2 49203 1 481
2 49204 1 481
2 49205 1 481
2 49206 1 481
2 49207 1 481
2 49208 1 481
2 49209 1 481
2 49210 1 481
2 49211 1 481
2 49212 1 481
2 49213 1 481
2 49214 1 481
2 49215 1 481
2 49216 1 481
2 49217 1 481
2 49218 1 481
2 49219 1 481
2 49220 1 481
2 49221 1 481
2 49222 1 481
2 49223 1 481
2 49224 1 481
2 49225 1 481
2 49226 1 481
2 49227 1 481
2 49228 1 481
2 49229 1 481
2 49230 1 481
2 49231 1 481
2 49232 1 481
2 49233 1 481
2 49234 1 481
2 49235 1 481
2 49236 1 481
2 49237 1 481
2 49238 1 481
2 49239 1 482
2 49240 1 482
2 49241 1 482
2 49242 1 482
2 49243 1 482
2 49244 1 482
2 49245 1 482
2 49246 1 482
2 49247 1 482
2 49248 1 482
2 49249 1 482
2 49250 1 482
2 49251 1 482
2 49252 1 482
2 49253 1 482
2 49254 1 482
2 49255 1 486
2 49256 1 486
2 49257 1 486
2 49258 1 487
2 49259 1 487
2 49260 1 487
2 49261 1 499
2 49262 1 499
2 49263 1 499
2 49264 1 499
2 49265 1 499
2 49266 1 499
2 49267 1 499
2 49268 1 499
2 49269 1 499
2 49270 1 499
2 49271 1 499
2 49272 1 501
2 49273 1 501
2 49274 1 501
2 49275 1 501
2 49276 1 501
2 49277 1 501
2 49278 1 501
2 49279 1 501
2 49280 1 501
2 49281 1 501
2 49282 1 501
2 49283 1 501
2 49284 1 501
2 49285 1 501
2 49286 1 503
2 49287 1 503
2 49288 1 504
2 49289 1 504
2 49290 1 504
2 49291 1 516
2 49292 1 516
2 49293 1 516
2 49294 1 516
2 49295 1 516
2 49296 1 517
2 49297 1 517
2 49298 1 517
2 49299 1 517
2 49300 1 518
2 49301 1 518
2 49302 1 519
2 49303 1 519
2 49304 1 520
2 49305 1 520
2 49306 1 520
2 49307 1 520
2 49308 1 520
2 49309 1 520
2 49310 1 521
2 49311 1 521
2 49312 1 528
2 49313 1 528
2 49314 1 528
2 49315 1 528
2 49316 1 528
2 49317 1 528
2 49318 1 529
2 49319 1 529
2 49320 1 529
2 49321 1 529
2 49322 1 529
2 49323 1 529
2 49324 1 529
2 49325 1 529
2 49326 1 530
2 49327 1 530
2 49328 1 530
2 49329 1 532
2 49330 1 532
2 49331 1 532
2 49332 1 532
2 49333 1 532
2 49334 1 532
2 49335 1 532
2 49336 1 534
2 49337 1 534
2 49338 1 537
2 49339 1 537
2 49340 1 537
2 49341 1 540
2 49342 1 540
2 49343 1 540
2 49344 1 541
2 49345 1 541
2 49346 1 541
2 49347 1 541
2 49348 1 546
2 49349 1 546
2 49350 1 557
2 49351 1 557
2 49352 1 557
2 49353 1 557
2 49354 1 557
2 49355 1 557
2 49356 1 557
2 49357 1 557
2 49358 1 557
2 49359 1 557
2 49360 1 565
2 49361 1 565
2 49362 1 565
2 49363 1 565
2 49364 1 565
2 49365 1 565
2 49366 1 565
2 49367 1 566
2 49368 1 566
2 49369 1 566
2 49370 1 566
2 49371 1 566
2 49372 1 566
2 49373 1 566
2 49374 1 566
2 49375 1 566
2 49376 1 566
2 49377 1 566
2 49378 1 575
2 49379 1 575
2 49380 1 575
2 49381 1 575
2 49382 1 576
2 49383 1 576
2 49384 1 576
2 49385 1 576
2 49386 1 576
2 49387 1 576
2 49388 1 578
2 49389 1 578
2 49390 1 578
2 49391 1 578
2 49392 1 578
2 49393 1 578
2 49394 1 578
2 49395 1 578
2 49396 1 578
2 49397 1 578
2 49398 1 578
2 49399 1 578
2 49400 1 578
2 49401 1 578
2 49402 1 578
2 49403 1 578
2 49404 1 578
2 49405 1 578
2 49406 1 578
2 49407 1 578
2 49408 1 578
2 49409 1 578
2 49410 1 578
2 49411 1 578
2 49412 1 578
2 49413 1 578
2 49414 1 578
2 49415 1 578
2 49416 1 578
2 49417 1 578
2 49418 1 578
2 49419 1 578
2 49420 1 578
2 49421 1 578
2 49422 1 578
2 49423 1 578
2 49424 1 578
2 49425 1 578
2 49426 1 578
2 49427 1 578
2 49428 1 578
2 49429 1 578
2 49430 1 578
2 49431 1 578
2 49432 1 578
2 49433 1 578
2 49434 1 578
2 49435 1 578
2 49436 1 578
2 49437 1 578
2 49438 1 578
2 49439 1 578
2 49440 1 578
2 49441 1 578
2 49442 1 578
2 49443 1 578
2 49444 1 578
2 49445 1 578
2 49446 1 578
2 49447 1 578
2 49448 1 578
2 49449 1 578
2 49450 1 578
2 49451 1 578
2 49452 1 578
2 49453 1 578
2 49454 1 578
2 49455 1 578
2 49456 1 579
2 49457 1 579
2 49458 1 579
2 49459 1 579
2 49460 1 579
2 49461 1 579
2 49462 1 579
2 49463 1 579
2 49464 1 579
2 49465 1 579
2 49466 1 579
2 49467 1 579
2 49468 1 579
2 49469 1 579
2 49470 1 579
2 49471 1 579
2 49472 1 579
2 49473 1 579
2 49474 1 579
2 49475 1 579
2 49476 1 579
2 49477 1 579
2 49478 1 579
2 49479 1 579
2 49480 1 579
2 49481 1 579
2 49482 1 579
2 49483 1 579
2 49484 1 579
2 49485 1 579
2 49486 1 579
2 49487 1 579
2 49488 1 579
2 49489 1 579
2 49490 1 579
2 49491 1 579
2 49492 1 579
2 49493 1 579
2 49494 1 579
2 49495 1 579
2 49496 1 579
2 49497 1 579
2 49498 1 579
2 49499 1 579
2 49500 1 579
2 49501 1 579
2 49502 1 579
2 49503 1 579
2 49504 1 579
2 49505 1 579
2 49506 1 579
2 49507 1 579
2 49508 1 579
2 49509 1 579
2 49510 1 579
2 49511 1 579
2 49512 1 579
2 49513 1 579
2 49514 1 579
2 49515 1 579
2 49516 1 579
2 49517 1 579
2 49518 1 579
2 49519 1 579
2 49520 1 579
2 49521 1 579
2 49522 1 579
2 49523 1 579
2 49524 1 579
2 49525 1 579
2 49526 1 579
2 49527 1 579
2 49528 1 579
2 49529 1 579
2 49530 1 579
2 49531 1 579
2 49532 1 579
2 49533 1 579
2 49534 1 579
2 49535 1 579
2 49536 1 579
2 49537 1 579
2 49538 1 579
2 49539 1 579
2 49540 1 579
2 49541 1 579
2 49542 1 579
2 49543 1 579
2 49544 1 579
2 49545 1 580
2 49546 1 580
2 49547 1 580
2 49548 1 580
2 49549 1 582
2 49550 1 582
2 49551 1 582
2 49552 1 585
2 49553 1 585
2 49554 1 585
2 49555 1 585
2 49556 1 585
2 49557 1 585
2 49558 1 585
2 49559 1 585
2 49560 1 585
2 49561 1 585
2 49562 1 585
2 49563 1 585
2 49564 1 585
2 49565 1 585
2 49566 1 585
2 49567 1 585
2 49568 1 585
2 49569 1 585
2 49570 1 585
2 49571 1 585
2 49572 1 585
2 49573 1 585
2 49574 1 585
2 49575 1 585
2 49576 1 585
2 49577 1 585
2 49578 1 585
2 49579 1 585
2 49580 1 585
2 49581 1 585
2 49582 1 585
2 49583 1 585
2 49584 1 585
2 49585 1 585
2 49586 1 585
2 49587 1 585
2 49588 1 585
2 49589 1 585
2 49590 1 585
2 49591 1 585
2 49592 1 585
2 49593 1 585
2 49594 1 585
2 49595 1 585
2 49596 1 585
2 49597 1 585
2 49598 1 585
2 49599 1 585
2 49600 1 585
2 49601 1 585
2 49602 1 585
2 49603 1 585
2 49604 1 585
2 49605 1 585
2 49606 1 585
2 49607 1 585
2 49608 1 585
2 49609 1 585
2 49610 1 585
2 49611 1 585
2 49612 1 585
2 49613 1 585
2 49614 1 585
2 49615 1 585
2 49616 1 585
2 49617 1 585
2 49618 1 585
2 49619 1 585
2 49620 1 585
2 49621 1 585
2 49622 1 585
2 49623 1 586
2 49624 1 586
2 49625 1 586
2 49626 1 586
2 49627 1 586
2 49628 1 586
2 49629 1 586
2 49630 1 586
2 49631 1 586
2 49632 1 586
2 49633 1 586
2 49634 1 586
2 49635 1 586
2 49636 1 586
2 49637 1 586
2 49638 1 586
2 49639 1 586
2 49640 1 586
2 49641 1 586
2 49642 1 586
2 49643 1 586
2 49644 1 586
2 49645 1 586
2 49646 1 586
2 49647 1 586
2 49648 1 586
2 49649 1 586
2 49650 1 586
2 49651 1 586
2 49652 1 586
2 49653 1 586
2 49654 1 586
2 49655 1 586
2 49656 1 586
2 49657 1 586
2 49658 1 586
2 49659 1 586
2 49660 1 586
2 49661 1 586
2 49662 1 586
2 49663 1 586
2 49664 1 586
2 49665 1 586
2 49666 1 586
2 49667 1 586
2 49668 1 586
2 49669 1 586
2 49670 1 586
2 49671 1 586
2 49672 1 586
2 49673 1 586
2 49674 1 586
2 49675 1 586
2 49676 1 586
2 49677 1 586
2 49678 1 587
2 49679 1 587
2 49680 1 587
2 49681 1 587
2 49682 1 587
2 49683 1 587
2 49684 1 587
2 49685 1 587
2 49686 1 587
2 49687 1 587
2 49688 1 587
2 49689 1 588
2 49690 1 588
2 49691 1 588
2 49692 1 588
2 49693 1 588
2 49694 1 588
2 49695 1 588
2 49696 1 588
2 49697 1 589
2 49698 1 589
2 49699 1 590
2 49700 1 590
2 49701 1 591
2 49702 1 591
2 49703 1 593
2 49704 1 593
2 49705 1 594
2 49706 1 594
2 49707 1 595
2 49708 1 595
2 49709 1 595
2 49710 1 595
2 49711 1 595
2 49712 1 595
2 49713 1 595
2 49714 1 595
2 49715 1 595
2 49716 1 596
2 49717 1 596
2 49718 1 596
2 49719 1 596
2 49720 1 596
2 49721 1 596
2 49722 1 596
2 49723 1 596
2 49724 1 596
2 49725 1 598
2 49726 1 598
2 49727 1 608
2 49728 1 608
2 49729 1 608
2 49730 1 608
2 49731 1 608
2 49732 1 608
2 49733 1 608
2 49734 1 609
2 49735 1 609
2 49736 1 609
2 49737 1 610
2 49738 1 610
2 49739 1 610
2 49740 1 611
2 49741 1 611
2 49742 1 613
2 49743 1 613
2 49744 1 613
2 49745 1 613
2 49746 1 620
2 49747 1 620
2 49748 1 620
2 49749 1 620
2 49750 1 620
2 49751 1 620
2 49752 1 620
2 49753 1 620
2 49754 1 620
2 49755 1 620
2 49756 1 621
2 49757 1 621
2 49758 1 622
2 49759 1 622
2 49760 1 622
2 49761 1 622
2 49762 1 622
2 49763 1 622
2 49764 1 622
2 49765 1 622
2 49766 1 622
2 49767 1 623
2 49768 1 623
2 49769 1 623
2 49770 1 623
2 49771 1 623
2 49772 1 623
2 49773 1 623
2 49774 1 623
2 49775 1 623
2 49776 1 623
2 49777 1 623
2 49778 1 623
2 49779 1 623
2 49780 1 623
2 49781 1 623
2 49782 1 624
2 49783 1 624
2 49784 1 624
2 49785 1 624
2 49786 1 625
2 49787 1 625
2 49788 1 625
2 49789 1 625
2 49790 1 625
2 49791 1 625
2 49792 1 625
2 49793 1 626
2 49794 1 626
2 49795 1 635
2 49796 1 635
2 49797 1 635
2 49798 1 635
2 49799 1 635
2 49800 1 635
2 49801 1 635
2 49802 1 635
2 49803 1 635
2 49804 1 635
2 49805 1 635
2 49806 1 635
2 49807 1 635
2 49808 1 635
2 49809 1 635
2 49810 1 635
2 49811 1 635
2 49812 1 635
2 49813 1 635
2 49814 1 635
2 49815 1 635
2 49816 1 635
2 49817 1 636
2 49818 1 636
2 49819 1 636
2 49820 1 636
2 49821 1 637
2 49822 1 637
2 49823 1 637
2 49824 1 637
2 49825 1 637
2 49826 1 637
2 49827 1 637
2 49828 1 637
2 49829 1 638
2 49830 1 638
2 49831 1 638
2 49832 1 639
2 49833 1 639
2 49834 1 639
2 49835 1 639
2 49836 1 639
2 49837 1 639
2 49838 1 639
2 49839 1 639
2 49840 1 639
2 49841 1 639
2 49842 1 639
2 49843 1 640
2 49844 1 640
2 49845 1 640
2 49846 1 641
2 49847 1 641
2 49848 1 641
2 49849 1 641
2 49850 1 641
2 49851 1 641
2 49852 1 641
2 49853 1 641
2 49854 1 641
2 49855 1 641
2 49856 1 641
2 49857 1 642
2 49858 1 642
2 49859 1 651
2 49860 1 651
2 49861 1 651
2 49862 1 651
2 49863 1 651
2 49864 1 651
2 49865 1 651
2 49866 1 651
2 49867 1 651
2 49868 1 651
2 49869 1 652
2 49870 1 652
2 49871 1 652
2 49872 1 652
2 49873 1 652
2 49874 1 652
2 49875 1 652
2 49876 1 652
2 49877 1 652
2 49878 1 652
2 49879 1 652
2 49880 1 652
2 49881 1 652
2 49882 1 652
2 49883 1 652
2 49884 1 652
2 49885 1 652
2 49886 1 652
2 49887 1 652
2 49888 1 652
2 49889 1 652
2 49890 1 652
2 49891 1 652
2 49892 1 652
2 49893 1 652
2 49894 1 652
2 49895 1 652
2 49896 1 652
2 49897 1 652
2 49898 1 652
2 49899 1 652
2 49900 1 652
2 49901 1 652
2 49902 1 652
2 49903 1 652
2 49904 1 652
2 49905 1 652
2 49906 1 652
2 49907 1 652
2 49908 1 652
2 49909 1 652
2 49910 1 653
2 49911 1 653
2 49912 1 654
2 49913 1 654
2 49914 1 654
2 49915 1 654
2 49916 1 654
2 49917 1 654
2 49918 1 655
2 49919 1 655
2 49920 1 655
2 49921 1 655
2 49922 1 655
2 49923 1 656
2 49924 1 656
2 49925 1 656
2 49926 1 656
2 49927 1 657
2 49928 1 657
2 49929 1 657
2 49930 1 657
2 49931 1 657
2 49932 1 657
2 49933 1 657
2 49934 1 657
2 49935 1 657
2 49936 1 657
2 49937 1 657
2 49938 1 657
2 49939 1 657
2 49940 1 657
2 49941 1 657
2 49942 1 659
2 49943 1 659
2 49944 1 659
2 49945 1 659
2 49946 1 659
2 49947 1 660
2 49948 1 660
2 49949 1 660
2 49950 1 660
2 49951 1 660
2 49952 1 660
2 49953 1 660
2 49954 1 660
2 49955 1 661
2 49956 1 661
2 49957 1 661
2 49958 1 661
2 49959 1 661
2 49960 1 661
2 49961 1 663
2 49962 1 663
2 49963 1 663
2 49964 1 663
2 49965 1 663
2 49966 1 663
2 49967 1 663
2 49968 1 664
2 49969 1 664
2 49970 1 664
2 49971 1 664
2 49972 1 664
2 49973 1 664
2 49974 1 664
2 49975 1 664
2 49976 1 664
2 49977 1 664
2 49978 1 664
2 49979 1 664
2 49980 1 664
2 49981 1 664
2 49982 1 664
2 49983 1 664
2 49984 1 664
2 49985 1 664
2 49986 1 664
2 49987 1 664
2 49988 1 664
2 49989 1 664
2 49990 1 666
2 49991 1 666
2 49992 1 666
2 49993 1 666
2 49994 1 666
2 49995 1 666
2 49996 1 666
2 49997 1 666
2 49998 1 666
2 49999 1 666
2 50000 1 666
2 50001 1 666
2 50002 1 666
2 50003 1 666
2 50004 1 666
2 50005 1 666
2 50006 1 666
2 50007 1 666
2 50008 1 666
2 50009 1 666
2 50010 1 666
2 50011 1 666
2 50012 1 666
2 50013 1 667
2 50014 1 667
2 50015 1 667
2 50016 1 667
2 50017 1 669
2 50018 1 669
2 50019 1 669
2 50020 1 669
2 50021 1 669
2 50022 1 669
2 50023 1 669
2 50024 1 669
2 50025 1 669
2 50026 1 674
2 50027 1 674
2 50028 1 674
2 50029 1 674
2 50030 1 674
2 50031 1 674
2 50032 1 674
2 50033 1 674
2 50034 1 674
2 50035 1 674
2 50036 1 675
2 50037 1 675
2 50038 1 677
2 50039 1 677
2 50040 1 677
2 50041 1 678
2 50042 1 678
2 50043 1 678
2 50044 1 678
2 50045 1 678
2 50046 1 679
2 50047 1 679
2 50048 1 679
2 50049 1 680
2 50050 1 680
2 50051 1 681
2 50052 1 681
2 50053 1 686
2 50054 1 686
2 50055 1 686
2 50056 1 686
2 50057 1 686
2 50058 1 686
2 50059 1 686
2 50060 1 686
2 50061 1 686
2 50062 1 686
2 50063 1 687
2 50064 1 687
2 50065 1 687
2 50066 1 687
2 50067 1 687
2 50068 1 687
2 50069 1 687
2 50070 1 687
2 50071 1 687
2 50072 1 687
2 50073 1 687
2 50074 1 687
2 50075 1 687
2 50076 1 695
2 50077 1 695
2 50078 1 697
2 50079 1 697
2 50080 1 697
2 50081 1 706
2 50082 1 706
2 50083 1 708
2 50084 1 708
2 50085 1 708
2 50086 1 708
2 50087 1 708
2 50088 1 708
2 50089 1 708
2 50090 1 708
2 50091 1 709
2 50092 1 709
2 50093 1 709
2 50094 1 710
2 50095 1 710
2 50096 1 710
2 50097 1 710
2 50098 1 710
2 50099 1 710
2 50100 1 711
2 50101 1 711
2 50102 1 713
2 50103 1 713
2 50104 1 713
2 50105 1 713
2 50106 1 713
2 50107 1 713
2 50108 1 713
2 50109 1 713
2 50110 1 713
2 50111 1 714
2 50112 1 714
2 50113 1 714
2 50114 1 725
2 50115 1 725
2 50116 1 726
2 50117 1 726
2 50118 1 726
2 50119 1 726
2 50120 1 726
2 50121 1 726
2 50122 1 727
2 50123 1 727
2 50124 1 727
2 50125 1 728
2 50126 1 728
2 50127 1 728
2 50128 1 728
2 50129 1 728
2 50130 1 728
2 50131 1 728
2 50132 1 728
2 50133 1 728
2 50134 1 728
2 50135 1 728
2 50136 1 728
2 50137 1 728
2 50138 1 729
2 50139 1 729
2 50140 1 729
2 50141 1 739
2 50142 1 739
2 50143 1 739
2 50144 1 739
2 50145 1 739
2 50146 1 739
2 50147 1 739
2 50148 1 739
2 50149 1 739
2 50150 1 740
2 50151 1 740
2 50152 1 740
2 50153 1 740
2 50154 1 740
2 50155 1 740
2 50156 1 742
2 50157 1 742
2 50158 1 742
2 50159 1 742
2 50160 1 742
2 50161 1 742
2 50162 1 742
2 50163 1 743
2 50164 1 743
2 50165 1 743
2 50166 1 743
2 50167 1 743
2 50168 1 743
2 50169 1 745
2 50170 1 745
2 50171 1 747
2 50172 1 747
2 50173 1 748
2 50174 1 748
2 50175 1 748
2 50176 1 748
2 50177 1 748
2 50178 1 748
2 50179 1 748
2 50180 1 748
2 50181 1 748
2 50182 1 748
2 50183 1 748
2 50184 1 748
2 50185 1 748
2 50186 1 748
2 50187 1 748
2 50188 1 749
2 50189 1 749
2 50190 1 750
2 50191 1 750
2 50192 1 750
2 50193 1 750
2 50194 1 750
2 50195 1 750
2 50196 1 750
2 50197 1 751
2 50198 1 751
2 50199 1 751
2 50200 1 751
2 50201 1 751
2 50202 1 751
2 50203 1 751
2 50204 1 751
2 50205 1 751
2 50206 1 751
2 50207 1 751
2 50208 1 751
2 50209 1 751
2 50210 1 751
2 50211 1 751
2 50212 1 751
2 50213 1 751
2 50214 1 751
2 50215 1 751
2 50216 1 751
2 50217 1 751
2 50218 1 751
2 50219 1 753
2 50220 1 753
2 50221 1 754
2 50222 1 754
2 50223 1 754
2 50224 1 754
2 50225 1 754
2 50226 1 754
2 50227 1 754
2 50228 1 754
2 50229 1 754
2 50230 1 754
2 50231 1 754
2 50232 1 754
2 50233 1 754
2 50234 1 754
2 50235 1 755
2 50236 1 755
2 50237 1 755
2 50238 1 755
2 50239 1 755
2 50240 1 755
2 50241 1 755
2 50242 1 756
2 50243 1 756
2 50244 1 756
2 50245 1 756
2 50246 1 756
2 50247 1 757
2 50248 1 757
2 50249 1 757
2 50250 1 763
2 50251 1 763
2 50252 1 763
2 50253 1 770
2 50254 1 770
2 50255 1 770
2 50256 1 770
2 50257 1 770
2 50258 1 771
2 50259 1 771
2 50260 1 771
2 50261 1 771
2 50262 1 771
2 50263 1 771
2 50264 1 771
2 50265 1 771
2 50266 1 772
2 50267 1 772
2 50268 1 773
2 50269 1 773
2 50270 1 776
2 50271 1 776
2 50272 1 776
2 50273 1 776
2 50274 1 776
2 50275 1 776
2 50276 1 776
2 50277 1 776
2 50278 1 776
2 50279 1 776
2 50280 1 776
2 50281 1 776
2 50282 1 776
2 50283 1 776
2 50284 1 776
2 50285 1 776
2 50286 1 776
2 50287 1 776
2 50288 1 776
2 50289 1 776
2 50290 1 776
2 50291 1 776
2 50292 1 776
2 50293 1 776
2 50294 1 777
2 50295 1 777
2 50296 1 778
2 50297 1 778
2 50298 1 778
2 50299 1 778
2 50300 1 778
2 50301 1 778
2 50302 1 785
2 50303 1 785
2 50304 1 785
2 50305 1 785
2 50306 1 785
2 50307 1 785
2 50308 1 785
2 50309 1 786
2 50310 1 786
2 50311 1 786
2 50312 1 786
2 50313 1 786
2 50314 1 786
2 50315 1 787
2 50316 1 787
2 50317 1 787
2 50318 1 787
2 50319 1 787
2 50320 1 787
2 50321 1 787
2 50322 1 787
2 50323 1 787
2 50324 1 787
2 50325 1 787
2 50326 1 787
2 50327 1 787
2 50328 1 787
2 50329 1 787
2 50330 1 787
2 50331 1 787
2 50332 1 787
2 50333 1 787
2 50334 1 787
2 50335 1 787
2 50336 1 788
2 50337 1 788
2 50338 1 788
2 50339 1 788
2 50340 1 788
2 50341 1 797
2 50342 1 797
2 50343 1 797
2 50344 1 797
2 50345 1 797
2 50346 1 797
2 50347 1 797
2 50348 1 798
2 50349 1 798
2 50350 1 798
2 50351 1 798
2 50352 1 798
2 50353 1 798
2 50354 1 798
2 50355 1 798
2 50356 1 798
2 50357 1 798
2 50358 1 798
2 50359 1 799
2 50360 1 799
2 50361 1 799
2 50362 1 799
2 50363 1 799
2 50364 1 801
2 50365 1 801
2 50366 1 803
2 50367 1 803
2 50368 1 803
2 50369 1 803
2 50370 1 803
2 50371 1 803
2 50372 1 803
2 50373 1 803
2 50374 1 803
2 50375 1 803
2 50376 1 803
2 50377 1 804
2 50378 1 804
2 50379 1 804
2 50380 1 804
2 50381 1 804
2 50382 1 804
2 50383 1 804
2 50384 1 804
2 50385 1 804
2 50386 1 804
2 50387 1 804
2 50388 1 804
2 50389 1 804
2 50390 1 804
2 50391 1 805
2 50392 1 805
2 50393 1 805
2 50394 1 805
2 50395 1 805
2 50396 1 805
2 50397 1 805
2 50398 1 805
2 50399 1 805
2 50400 1 805
2 50401 1 805
2 50402 1 805
2 50403 1 805
2 50404 1 806
2 50405 1 806
2 50406 1 813
2 50407 1 813
2 50408 1 813
2 50409 1 813
2 50410 1 813
2 50411 1 814
2 50412 1 814
2 50413 1 815
2 50414 1 815
2 50415 1 815
2 50416 1 815
2 50417 1 815
2 50418 1 815
2 50419 1 815
2 50420 1 815
2 50421 1 815
2 50422 1 815
2 50423 1 816
2 50424 1 816
2 50425 1 816
2 50426 1 816
2 50427 1 817
2 50428 1 817
2 50429 1 817
2 50430 1 817
2 50431 1 817
2 50432 1 817
2 50433 1 817
2 50434 1 817
2 50435 1 817
2 50436 1 817
2 50437 1 817
2 50438 1 817
2 50439 1 817
2 50440 1 817
2 50441 1 817
2 50442 1 817
2 50443 1 817
2 50444 1 817
2 50445 1 817
2 50446 1 817
2 50447 1 817
2 50448 1 818
2 50449 1 818
2 50450 1 818
2 50451 1 818
2 50452 1 818
2 50453 1 818
2 50454 1 818
2 50455 1 818
2 50456 1 818
2 50457 1 818
2 50458 1 818
2 50459 1 818
2 50460 1 818
2 50461 1 819
2 50462 1 819
2 50463 1 820
2 50464 1 820
2 50465 1 822
2 50466 1 822
2 50467 1 822
2 50468 1 825
2 50469 1 825
2 50470 1 825
2 50471 1 825
2 50472 1 825
2 50473 1 825
2 50474 1 825
2 50475 1 825
2 50476 1 825
2 50477 1 825
2 50478 1 825
2 50479 1 825
2 50480 1 825
2 50481 1 825
2 50482 1 825
2 50483 1 825
2 50484 1 825
2 50485 1 825
2 50486 1 825
2 50487 1 825
2 50488 1 825
2 50489 1 826
2 50490 1 826
2 50491 1 826
2 50492 1 827
2 50493 1 827
2 50494 1 827
2 50495 1 827
2 50496 1 828
2 50497 1 828
2 50498 1 828
2 50499 1 828
2 50500 1 828
2 50501 1 829
2 50502 1 829
2 50503 1 830
2 50504 1 830
2 50505 1 830
2 50506 1 830
2 50507 1 830
2 50508 1 830
2 50509 1 830
2 50510 1 830
2 50511 1 830
2 50512 1 830
2 50513 1 830
2 50514 1 830
2 50515 1 830
2 50516 1 830
2 50517 1 830
2 50518 1 830
2 50519 1 830
2 50520 1 830
2 50521 1 831
2 50522 1 831
2 50523 1 831
2 50524 1 831
2 50525 1 831
2 50526 1 832
2 50527 1 832
2 50528 1 832
2 50529 1 832
2 50530 1 841
2 50531 1 841
2 50532 1 841
2 50533 1 841
2 50534 1 842
2 50535 1 842
2 50536 1 847
2 50537 1 847
2 50538 1 847
2 50539 1 847
2 50540 1 847
2 50541 1 847
2 50542 1 855
2 50543 1 855
2 50544 1 857
2 50545 1 857
2 50546 1 857
2 50547 1 857
2 50548 1 858
2 50549 1 858
2 50550 1 858
2 50551 1 858
2 50552 1 858
2 50553 1 858
2 50554 1 858
2 50555 1 859
2 50556 1 859
2 50557 1 859
2 50558 1 859
2 50559 1 859
2 50560 1 859
2 50561 1 859
2 50562 1 859
2 50563 1 859
2 50564 1 859
2 50565 1 860
2 50566 1 860
2 50567 1 860
2 50568 1 860
2 50569 1 861
2 50570 1 861
2 50571 1 862
2 50572 1 862
2 50573 1 862
2 50574 1 866
2 50575 1 866
2 50576 1 866
2 50577 1 866
2 50578 1 866
2 50579 1 866
2 50580 1 866
2 50581 1 866
2 50582 1 866
2 50583 1 866
2 50584 1 866
2 50585 1 866
2 50586 1 866
2 50587 1 866
2 50588 1 866
2 50589 1 866
2 50590 1 866
2 50591 1 866
2 50592 1 866
2 50593 1 866
2 50594 1 866
2 50595 1 866
2 50596 1 866
2 50597 1 866
2 50598 1 866
2 50599 1 866
2 50600 1 867
2 50601 1 867
2 50602 1 867
2 50603 1 867
2 50604 1 867
2 50605 1 867
2 50606 1 867
2 50607 1 867
2 50608 1 868
2 50609 1 868
2 50610 1 869
2 50611 1 869
2 50612 1 882
2 50613 1 882
2 50614 1 882
2 50615 1 882
2 50616 1 883
2 50617 1 883
2 50618 1 883
2 50619 1 883
2 50620 1 883
2 50621 1 883
2 50622 1 883
2 50623 1 883
2 50624 1 883
2 50625 1 883
2 50626 1 884
2 50627 1 884
2 50628 1 893
2 50629 1 893
2 50630 1 893
2 50631 1 893
2 50632 1 893
2 50633 1 893
2 50634 1 895
2 50635 1 895
2 50636 1 895
2 50637 1 895
2 50638 1 895
2 50639 1 895
2 50640 1 895
2 50641 1 895
2 50642 1 895
2 50643 1 895
2 50644 1 895
2 50645 1 896
2 50646 1 896
2 50647 1 898
2 50648 1 898
2 50649 1 898
2 50650 1 898
2 50651 1 898
2 50652 1 898
2 50653 1 898
2 50654 1 898
2 50655 1 898
2 50656 1 898
2 50657 1 906
2 50658 1 906
2 50659 1 906
2 50660 1 906
2 50661 1 906
2 50662 1 906
2 50663 1 906
2 50664 1 906
2 50665 1 906
2 50666 1 907
2 50667 1 907
2 50668 1 907
2 50669 1 908
2 50670 1 908
2 50671 1 908
2 50672 1 908
2 50673 1 908
2 50674 1 908
2 50675 1 908
2 50676 1 908
2 50677 1 909
2 50678 1 909
2 50679 1 909
2 50680 1 909
2 50681 1 909
2 50682 1 909
2 50683 1 909
2 50684 1 909
2 50685 1 910
2 50686 1 910
2 50687 1 910
2 50688 1 910
2 50689 1 910
2 50690 1 910
2 50691 1 910
2 50692 1 910
2 50693 1 910
2 50694 1 910
2 50695 1 910
2 50696 1 910
2 50697 1 910
2 50698 1 910
2 50699 1 910
2 50700 1 910
2 50701 1 910
2 50702 1 910
2 50703 1 910
2 50704 1 910
2 50705 1 910
2 50706 1 910
2 50707 1 911
2 50708 1 911
2 50709 1 911
2 50710 1 911
2 50711 1 911
2 50712 1 911
2 50713 1 911
2 50714 1 911
2 50715 1 911
2 50716 1 911
2 50717 1 911
2 50718 1 911
2 50719 1 911
2 50720 1 911
2 50721 1 911
2 50722 1 911
2 50723 1 912
2 50724 1 912
2 50725 1 914
2 50726 1 914
2 50727 1 916
2 50728 1 916
2 50729 1 916
2 50730 1 916
2 50731 1 916
2 50732 1 916
2 50733 1 916
2 50734 1 916
2 50735 1 916
2 50736 1 916
2 50737 1 916
2 50738 1 916
2 50739 1 916
2 50740 1 916
2 50741 1 925
2 50742 1 925
2 50743 1 926
2 50744 1 926
2 50745 1 926
2 50746 1 926
2 50747 1 926
2 50748 1 926
2 50749 1 926
2 50750 1 926
2 50751 1 926
2 50752 1 926
2 50753 1 926
2 50754 1 926
2 50755 1 929
2 50756 1 929
2 50757 1 929
2 50758 1 929
2 50759 1 929
2 50760 1 929
2 50761 1 929
2 50762 1 929
2 50763 1 929
2 50764 1 929
2 50765 1 929
2 50766 1 929
2 50767 1 929
2 50768 1 930
2 50769 1 930
2 50770 1 930
2 50771 1 930
2 50772 1 930
2 50773 1 939
2 50774 1 939
2 50775 1 939
2 50776 1 939
2 50777 1 939
2 50778 1 939
2 50779 1 939
2 50780 1 939
2 50781 1 940
2 50782 1 940
2 50783 1 940
2 50784 1 940
2 50785 1 940
2 50786 1 940
2 50787 1 940
2 50788 1 942
2 50789 1 942
2 50790 1 944
2 50791 1 944
2 50792 1 944
2 50793 1 944
2 50794 1 944
2 50795 1 944
2 50796 1 944
2 50797 1 944
2 50798 1 944
2 50799 1 944
2 50800 1 945
2 50801 1 945
2 50802 1 952
2 50803 1 952
2 50804 1 952
2 50805 1 952
2 50806 1 952
2 50807 1 952
2 50808 1 952
2 50809 1 952
2 50810 1 952
2 50811 1 952
2 50812 1 952
2 50813 1 952
2 50814 1 952
2 50815 1 952
2 50816 1 952
2 50817 1 952
2 50818 1 952
2 50819 1 953
2 50820 1 953
2 50821 1 954
2 50822 1 954
2 50823 1 954
2 50824 1 954
2 50825 1 954
2 50826 1 955
2 50827 1 955
2 50828 1 955
2 50829 1 956
2 50830 1 956
2 50831 1 956
2 50832 1 956
2 50833 1 956
2 50834 1 956
2 50835 1 956
2 50836 1 956
2 50837 1 956
2 50838 1 956
2 50839 1 956
2 50840 1 957
2 50841 1 957
2 50842 1 957
2 50843 1 957
2 50844 1 957
2 50845 1 957
2 50846 1 957
2 50847 1 957
2 50848 1 957
2 50849 1 957
2 50850 1 957
2 50851 1 957
2 50852 1 957
2 50853 1 957
2 50854 1 957
2 50855 1 959
2 50856 1 959
2 50857 1 959
2 50858 1 963
2 50859 1 963
2 50860 1 963
2 50861 1 963
2 50862 1 963
2 50863 1 970
2 50864 1 970
2 50865 1 970
2 50866 1 970
2 50867 1 970
2 50868 1 970
2 50869 1 970
2 50870 1 971
2 50871 1 971
2 50872 1 971
2 50873 1 971
2 50874 1 971
2 50875 1 971
2 50876 1 971
2 50877 1 971
2 50878 1 971
2 50879 1 971
2 50880 1 971
2 50881 1 971
2 50882 1 971
2 50883 1 971
2 50884 1 972
2 50885 1 972
2 50886 1 972
2 50887 1 973
2 50888 1 973
2 50889 1 973
2 50890 1 973
2 50891 1 973
2 50892 1 973
2 50893 1 973
2 50894 1 973
2 50895 1 974
2 50896 1 974
2 50897 1 974
2 50898 1 974
2 50899 1 976
2 50900 1 976
2 50901 1 976
2 50902 1 976
2 50903 1 976
2 50904 1 976
2 50905 1 977
2 50906 1 977
2 50907 1 977
2 50908 1 980
2 50909 1 980
2 50910 1 980
2 50911 1 980
2 50912 1 980
2 50913 1 981
2 50914 1 981
2 50915 1 992
2 50916 1 992
2 50917 1 992
2 50918 1 992
2 50919 1 992
2 50920 1 992
2 50921 1 992
2 50922 1 992
2 50923 1 992
2 50924 1 992
2 50925 1 993
2 50926 1 993
2 50927 1 993
2 50928 1 993
2 50929 1 993
2 50930 1 993
2 50931 1 993
2 50932 1 993
2 50933 1 994
2 50934 1 994
2 50935 1 994
2 50936 1 994
2 50937 1 995
2 50938 1 995
2 50939 1 998
2 50940 1 998
2 50941 1 998
2 50942 1 998
2 50943 1 998
2 50944 1 998
2 50945 1 998
2 50946 1 999
2 50947 1 999
2 50948 1 999
2 50949 1 999
2 50950 1 1000
2 50951 1 1000
2 50952 1 1000
2 50953 1 1003
2 50954 1 1003
2 50955 1 1003
2 50956 1 1003
2 50957 1 1003
2 50958 1 1003
2 50959 1 1003
2 50960 1 1003
2 50961 1 1004
2 50962 1 1004
2 50963 1 1004
2 50964 1 1004
2 50965 1 1017
2 50966 1 1017
2 50967 1 1017
2 50968 1 1017
2 50969 1 1018
2 50970 1 1018
2 50971 1 1018
2 50972 1 1018
2 50973 1 1018
2 50974 1 1018
2 50975 1 1018
2 50976 1 1027
2 50977 1 1027
2 50978 1 1027
2 50979 1 1027
2 50980 1 1027
2 50981 1 1028
2 50982 1 1028
2 50983 1 1028
2 50984 1 1028
2 50985 1 1028
2 50986 1 1028
2 50987 1 1028
2 50988 1 1029
2 50989 1 1029
2 50990 1 1030
2 50991 1 1030
2 50992 1 1032
2 50993 1 1032
2 50994 1 1032
2 50995 1 1032
2 50996 1 1033
2 50997 1 1033
2 50998 1 1033
2 50999 1 1033
2 51000 1 1033
2 51001 1 1033
2 51002 1 1034
2 51003 1 1034
2 51004 1 1044
2 51005 1 1044
2 51006 1 1044
2 51007 1 1045
2 51008 1 1045
2 51009 1 1056
2 51010 1 1056
2 51011 1 1056
2 51012 1 1056
2 51013 1 1056
2 51014 1 1056
2 51015 1 1057
2 51016 1 1057
2 51017 1 1058
2 51018 1 1058
2 51019 1 1058
2 51020 1 1058
2 51021 1 1058
2 51022 1 1058
2 51023 1 1058
2 51024 1 1058
2 51025 1 1058
2 51026 1 1058
2 51027 1 1058
2 51028 1 1058
2 51029 1 1058
2 51030 1 1058
2 51031 1 1058
2 51032 1 1058
2 51033 1 1058
2 51034 1 1058
2 51035 1 1058
2 51036 1 1058
2 51037 1 1058
2 51038 1 1058
2 51039 1 1058
2 51040 1 1058
2 51041 1 1058
2 51042 1 1058
2 51043 1 1058
2 51044 1 1058
2 51045 1 1058
2 51046 1 1058
2 51047 1 1058
2 51048 1 1058
2 51049 1 1058
2 51050 1 1058
2 51051 1 1058
2 51052 1 1058
2 51053 1 1058
2 51054 1 1058
2 51055 1 1058
2 51056 1 1059
2 51057 1 1059
2 51058 1 1059
2 51059 1 1059
2 51060 1 1059
2 51061 1 1059
2 51062 1 1059
2 51063 1 1059
2 51064 1 1059
2 51065 1 1059
2 51066 1 1060
2 51067 1 1060
2 51068 1 1060
2 51069 1 1060
2 51070 1 1062
2 51071 1 1062
2 51072 1 1072
2 51073 1 1072
2 51074 1 1072
2 51075 1 1072
2 51076 1 1072
2 51077 1 1072
2 51078 1 1073
2 51079 1 1073
2 51080 1 1073
2 51081 1 1073
2 51082 1 1073
2 51083 1 1073
2 51084 1 1073
2 51085 1 1076
2 51086 1 1076
2 51087 1 1076
2 51088 1 1076
2 51089 1 1076
2 51090 1 1077
2 51091 1 1077
2 51092 1 1077
2 51093 1 1077
2 51094 1 1077
2 51095 1 1078
2 51096 1 1078
2 51097 1 1078
2 51098 1 1078
2 51099 1 1079
2 51100 1 1079
2 51101 1 1079
2 51102 1 1084
2 51103 1 1084
2 51104 1 1084
2 51105 1 1087
2 51106 1 1087
2 51107 1 1089
2 51108 1 1089
2 51109 1 1092
2 51110 1 1092
2 51111 1 1101
2 51112 1 1101
2 51113 1 1102
2 51114 1 1102
2 51115 1 1105
2 51116 1 1105
2 51117 1 1105
2 51118 1 1105
2 51119 1 1106
2 51120 1 1106
2 51121 1 1107
2 51122 1 1107
2 51123 1 1107
2 51124 1 1107
2 51125 1 1107
2 51126 1 1107
2 51127 1 1107
2 51128 1 1108
2 51129 1 1108
2 51130 1 1116
2 51131 1 1116
2 51132 1 1116
2 51133 1 1118
2 51134 1 1118
2 51135 1 1119
2 51136 1 1119
2 51137 1 1121
2 51138 1 1121
2 51139 1 1128
2 51140 1 1128
2 51141 1 1151
2 51142 1 1151
2 51143 1 1151
2 51144 1 1151
2 51145 1 1152
2 51146 1 1152
2 51147 1 1152
2 51148 1 1152
2 51149 1 1152
2 51150 1 1153
2 51151 1 1153
2 51152 1 1153
2 51153 1 1153
2 51154 1 1154
2 51155 1 1154
2 51156 1 1155
2 51157 1 1155
2 51158 1 1155
2 51159 1 1155
2 51160 1 1155
2 51161 1 1155
2 51162 1 1156
2 51163 1 1156
2 51164 1 1156
2 51165 1 1156
2 51166 1 1156
2 51167 1 1157
2 51168 1 1157
2 51169 1 1157
2 51170 1 1157
2 51171 1 1157
2 51172 1 1157
2 51173 1 1157
2 51174 1 1157
2 51175 1 1157
2 51176 1 1157
2 51177 1 1161
2 51178 1 1161
2 51179 1 1161
2 51180 1 1168
2 51181 1 1168
2 51182 1 1181
2 51183 1 1181
2 51184 1 1181
2 51185 1 1181
2 51186 1 1181
2 51187 1 1182
2 51188 1 1182
2 51189 1 1183
2 51190 1 1183
2 51191 1 1184
2 51192 1 1184
2 51193 1 1185
2 51194 1 1185
2 51195 1 1185
2 51196 1 1186
2 51197 1 1186
2 51198 1 1186
2 51199 1 1186
2 51200 1 1186
2 51201 1 1186
2 51202 1 1186
2 51203 1 1186
2 51204 1 1188
2 51205 1 1188
2 51206 1 1189
2 51207 1 1189
2 51208 1 1190
2 51209 1 1190
2 51210 1 1192
2 51211 1 1192
2 51212 1 1202
2 51213 1 1202
2 51214 1 1202
2 51215 1 1202
2 51216 1 1202
2 51217 1 1202
2 51218 1 1202
2 51219 1 1202
2 51220 1 1202
2 51221 1 1202
2 51222 1 1202
2 51223 1 1202
2 51224 1 1202
2 51225 1 1202
2 51226 1 1202
2 51227 1 1202
2 51228 1 1203
2 51229 1 1203
2 51230 1 1203
2 51231 1 1206
2 51232 1 1206
2 51233 1 1206
2 51234 1 1206
2 51235 1 1206
2 51236 1 1207
2 51237 1 1207
2 51238 1 1207
2 51239 1 1207
2 51240 1 1209
2 51241 1 1209
2 51242 1 1209
2 51243 1 1209
2 51244 1 1211
2 51245 1 1211
2 51246 1 1212
2 51247 1 1212
2 51248 1 1212
2 51249 1 1213
2 51250 1 1213
2 51251 1 1213
2 51252 1 1213
2 51253 1 1213
2 51254 1 1213
2 51255 1 1213
2 51256 1 1214
2 51257 1 1214
2 51258 1 1221
2 51259 1 1221
2 51260 1 1221
2 51261 1 1221
2 51262 1 1222
2 51263 1 1222
2 51264 1 1222
2 51265 1 1223
2 51266 1 1223
2 51267 1 1223
2 51268 1 1225
2 51269 1 1225
2 51270 1 1225
2 51271 1 1225
2 51272 1 1225
2 51273 1 1225
2 51274 1 1225
2 51275 1 1225
2 51276 1 1225
2 51277 1 1225
2 51278 1 1225
2 51279 1 1225
2 51280 1 1225
2 51281 1 1225
2 51282 1 1226
2 51283 1 1226
2 51284 1 1226
2 51285 1 1229
2 51286 1 1229
2 51287 1 1229
2 51288 1 1229
2 51289 1 1229
2 51290 1 1229
2 51291 1 1229
2 51292 1 1229
2 51293 1 1229
2 51294 1 1229
2 51295 1 1229
2 51296 1 1245
2 51297 1 1245
2 51298 1 1245
2 51299 1 1245
2 51300 1 1245
2 51301 1 1245
2 51302 1 1245
2 51303 1 1245
2 51304 1 1256
2 51305 1 1256
2 51306 1 1259
2 51307 1 1259
2 51308 1 1259
2 51309 1 1259
2 51310 1 1259
2 51311 1 1259
2 51312 1 1260
2 51313 1 1260
2 51314 1 1267
2 51315 1 1267
2 51316 1 1267
2 51317 1 1267
2 51318 1 1267
2 51319 1 1267
2 51320 1 1268
2 51321 1 1268
2 51322 1 1268
2 51323 1 1268
2 51324 1 1268
2 51325 1 1268
2 51326 1 1268
2 51327 1 1268
2 51328 1 1268
2 51329 1 1268
2 51330 1 1268
2 51331 1 1276
2 51332 1 1276
2 51333 1 1276
2 51334 1 1276
2 51335 1 1276
2 51336 1 1276
2 51337 1 1276
2 51338 1 1276
2 51339 1 1276
2 51340 1 1276
2 51341 1 1276
2 51342 1 1277
2 51343 1 1277
2 51344 1 1277
2 51345 1 1277
2 51346 1 1277
2 51347 1 1285
2 51348 1 1285
2 51349 1 1286
2 51350 1 1286
2 51351 1 1286
2 51352 1 1287
2 51353 1 1287
2 51354 1 1287
2 51355 1 1288
2 51356 1 1288
2 51357 1 1289
2 51358 1 1289
2 51359 1 1290
2 51360 1 1290
2 51361 1 1291
2 51362 1 1291
2 51363 1 1291
2 51364 1 1291
2 51365 1 1291
2 51366 1 1291
2 51367 1 1291
2 51368 1 1291
2 51369 1 1291
2 51370 1 1291
2 51371 1 1291
2 51372 1 1291
2 51373 1 1292
2 51374 1 1292
2 51375 1 1292
2 51376 1 1293
2 51377 1 1293
2 51378 1 1293
2 51379 1 1294
2 51380 1 1294
2 51381 1 1294
2 51382 1 1294
2 51383 1 1294
2 51384 1 1294
2 51385 1 1294
2 51386 1 1294
2 51387 1 1294
2 51388 1 1304
2 51389 1 1304
2 51390 1 1304
2 51391 1 1304
2 51392 1 1304
2 51393 1 1304
2 51394 1 1304
2 51395 1 1304
2 51396 1 1304
2 51397 1 1304
2 51398 1 1304
2 51399 1 1304
2 51400 1 1304
2 51401 1 1304
2 51402 1 1304
2 51403 1 1304
2 51404 1 1306
2 51405 1 1306
2 51406 1 1306
2 51407 1 1306
2 51408 1 1306
2 51409 1 1306
2 51410 1 1307
2 51411 1 1307
2 51412 1 1307
2 51413 1 1310
2 51414 1 1310
2 51415 1 1310
2 51416 1 1310
2 51417 1 1310
2 51418 1 1310
2 51419 1 1310
2 51420 1 1315
2 51421 1 1315
2 51422 1 1315
2 51423 1 1315
2 51424 1 1315
2 51425 1 1315
2 51426 1 1315
2 51427 1 1315
2 51428 1 1323
2 51429 1 1323
2 51430 1 1323
2 51431 1 1323
2 51432 1 1323
2 51433 1 1323
2 51434 1 1324
2 51435 1 1324
2 51436 1 1324
2 51437 1 1324
2 51438 1 1324
2 51439 1 1324
2 51440 1 1325
2 51441 1 1325
2 51442 1 1325
2 51443 1 1333
2 51444 1 1333
2 51445 1 1333
2 51446 1 1333
2 51447 1 1334
2 51448 1 1334
2 51449 1 1336
2 51450 1 1336
2 51451 1 1336
2 51452 1 1336
2 51453 1 1336
2 51454 1 1336
2 51455 1 1336
2 51456 1 1336
2 51457 1 1336
2 51458 1 1336
2 51459 1 1336
2 51460 1 1336
2 51461 1 1336
2 51462 1 1336
2 51463 1 1336
2 51464 1 1338
2 51465 1 1338
2 51466 1 1338
2 51467 1 1338
2 51468 1 1338
2 51469 1 1338
2 51470 1 1338
2 51471 1 1338
2 51472 1 1338
2 51473 1 1338
2 51474 1 1338
2 51475 1 1338
2 51476 1 1339
2 51477 1 1339
2 51478 1 1342
2 51479 1 1342
2 51480 1 1342
2 51481 1 1351
2 51482 1 1351
2 51483 1 1351
2 51484 1 1351
2 51485 1 1351
2 51486 1 1351
2 51487 1 1351
2 51488 1 1351
2 51489 1 1351
2 51490 1 1351
2 51491 1 1351
2 51492 1 1351
2 51493 1 1352
2 51494 1 1352
2 51495 1 1352
2 51496 1 1355
2 51497 1 1355
2 51498 1 1355
2 51499 1 1363
2 51500 1 1363
2 51501 1 1363
2 51502 1 1363
2 51503 1 1364
2 51504 1 1364
2 51505 1 1370
2 51506 1 1370
2 51507 1 1370
2 51508 1 1370
2 51509 1 1370
2 51510 1 1371
2 51511 1 1371
2 51512 1 1373
2 51513 1 1373
2 51514 1 1373
2 51515 1 1373
2 51516 1 1373
2 51517 1 1373
2 51518 1 1373
2 51519 1 1373
2 51520 1 1373
2 51521 1 1373
2 51522 1 1373
2 51523 1 1373
2 51524 1 1373
2 51525 1 1373
2 51526 1 1373
2 51527 1 1373
2 51528 1 1373
2 51529 1 1373
2 51530 1 1373
2 51531 1 1373
2 51532 1 1373
2 51533 1 1373
2 51534 1 1373
2 51535 1 1373
2 51536 1 1373
2 51537 1 1373
2 51538 1 1373
2 51539 1 1373
2 51540 1 1373
2 51541 1 1373
2 51542 1 1373
2 51543 1 1373
2 51544 1 1373
2 51545 1 1373
2 51546 1 1373
2 51547 1 1373
2 51548 1 1373
2 51549 1 1373
2 51550 1 1373
2 51551 1 1373
2 51552 1 1373
2 51553 1 1373
2 51554 1 1373
2 51555 1 1373
2 51556 1 1373
2 51557 1 1373
2 51558 1 1373
2 51559 1 1373
2 51560 1 1373
2 51561 1 1373
2 51562 1 1373
2 51563 1 1373
2 51564 1 1373
2 51565 1 1373
2 51566 1 1373
2 51567 1 1373
2 51568 1 1373
2 51569 1 1373
2 51570 1 1373
2 51571 1 1373
2 51572 1 1374
2 51573 1 1374
2 51574 1 1374
2 51575 1 1382
2 51576 1 1382
2 51577 1 1382
2 51578 1 1382
2 51579 1 1383
2 51580 1 1383
2 51581 1 1383
2 51582 1 1383
2 51583 1 1384
2 51584 1 1384
2 51585 1 1384
2 51586 1 1385
2 51587 1 1385
2 51588 1 1386
2 51589 1 1386
2 51590 1 1386
2 51591 1 1386
2 51592 1 1386
2 51593 1 1386
2 51594 1 1386
2 51595 1 1386
2 51596 1 1387
2 51597 1 1387
2 51598 1 1388
2 51599 1 1388
2 51600 1 1391
2 51601 1 1391
2 51602 1 1391
2 51603 1 1391
2 51604 1 1391
2 51605 1 1391
2 51606 1 1391
2 51607 1 1391
2 51608 1 1391
2 51609 1 1391
2 51610 1 1391
2 51611 1 1391
2 51612 1 1391
2 51613 1 1391
2 51614 1 1391
2 51615 1 1391
2 51616 1 1391
2 51617 1 1393
2 51618 1 1393
2 51619 1 1393
2 51620 1 1394
2 51621 1 1394
2 51622 1 1394
2 51623 1 1394
2 51624 1 1394
2 51625 1 1394
2 51626 1 1394
2 51627 1 1394
2 51628 1 1394
2 51629 1 1394
2 51630 1 1394
2 51631 1 1394
2 51632 1 1395
2 51633 1 1395
2 51634 1 1395
2 51635 1 1396
2 51636 1 1396
2 51637 1 1397
2 51638 1 1397
2 51639 1 1407
2 51640 1 1407
2 51641 1 1407
2 51642 1 1407
2 51643 1 1407
2 51644 1 1407
2 51645 1 1407
2 51646 1 1407
2 51647 1 1408
2 51648 1 1408
2 51649 1 1415
2 51650 1 1415
2 51651 1 1416
2 51652 1 1416
2 51653 1 1416
2 51654 1 1416
2 51655 1 1416
2 51656 1 1416
2 51657 1 1416
2 51658 1 1432
2 51659 1 1432
2 51660 1 1432
2 51661 1 1433
2 51662 1 1433
2 51663 1 1446
2 51664 1 1446
2 51665 1 1446
2 51666 1 1446
2 51667 1 1447
2 51668 1 1447
2 51669 1 1447
2 51670 1 1447
2 51671 1 1447
2 51672 1 1447
2 51673 1 1447
2 51674 1 1447
2 51675 1 1448
2 51676 1 1448
2 51677 1 1449
2 51678 1 1449
2 51679 1 1450
2 51680 1 1450
2 51681 1 1464
2 51682 1 1464
2 51683 1 1464
2 51684 1 1464
2 51685 1 1464
2 51686 1 1464
2 51687 1 1464
2 51688 1 1464
2 51689 1 1464
2 51690 1 1467
2 51691 1 1467
2 51692 1 1478
2 51693 1 1478
2 51694 1 1478
2 51695 1 1479
2 51696 1 1479
2 51697 1 1479
2 51698 1 1479
2 51699 1 1479
2 51700 1 1479
2 51701 1 1479
2 51702 1 1480
2 51703 1 1480
2 51704 1 1480
2 51705 1 1480
2 51706 1 1480
2 51707 1 1480
2 51708 1 1480
2 51709 1 1481
2 51710 1 1481
2 51711 1 1481
2 51712 1 1481
2 51713 1 1482
2 51714 1 1482
2 51715 1 1482
2 51716 1 1484
2 51717 1 1484
2 51718 1 1511
2 51719 1 1511
2 51720 1 1512
2 51721 1 1512
2 51722 1 1512
2 51723 1 1512
2 51724 1 1512
2 51725 1 1512
2 51726 1 1512
2 51727 1 1512
2 51728 1 1512
2 51729 1 1512
2 51730 1 1512
2 51731 1 1512
2 51732 1 1516
2 51733 1 1516
2 51734 1 1518
2 51735 1 1518
2 51736 1 1519
2 51737 1 1519
2 51738 1 1519
2 51739 1 1519
2 51740 1 1519
2 51741 1 1519
2 51742 1 1519
2 51743 1 1519
2 51744 1 1519
2 51745 1 1519
2 51746 1 1519
2 51747 1 1520
2 51748 1 1520
2 51749 1 1521
2 51750 1 1521
2 51751 1 1525
2 51752 1 1525
2 51753 1 1525
2 51754 1 1525
2 51755 1 1525
2 51756 1 1525
2 51757 1 1526
2 51758 1 1526
2 51759 1 1526
2 51760 1 1526
2 51761 1 1526
2 51762 1 1526
2 51763 1 1526
2 51764 1 1526
2 51765 1 1526
2 51766 1 1534
2 51767 1 1534
2 51768 1 1534
2 51769 1 1536
2 51770 1 1536
2 51771 1 1537
2 51772 1 1537
2 51773 1 1540
2 51774 1 1540
2 51775 1 1540
2 51776 1 1540
2 51777 1 1541
2 51778 1 1541
2 51779 1 1541
2 51780 1 1541
2 51781 1 1541
2 51782 1 1541
2 51783 1 1542
2 51784 1 1542
2 51785 1 1542
2 51786 1 1547
2 51787 1 1547
2 51788 1 1550
2 51789 1 1550
2 51790 1 1550
2 51791 1 1550
2 51792 1 1550
2 51793 1 1550
2 51794 1 1550
2 51795 1 1551
2 51796 1 1551
2 51797 1 1551
2 51798 1 1552
2 51799 1 1552
2 51800 1 1552
2 51801 1 1553
2 51802 1 1553
2 51803 1 1553
2 51804 1 1553
2 51805 1 1555
2 51806 1 1555
2 51807 1 1559
2 51808 1 1559
2 51809 1 1560
2 51810 1 1560
2 51811 1 1560
2 51812 1 1561
2 51813 1 1561
2 51814 1 1561
2 51815 1 1561
2 51816 1 1561
2 51817 1 1561
2 51818 1 1561
2 51819 1 1561
2 51820 1 1561
2 51821 1 1561
2 51822 1 1561
2 51823 1 1561
2 51824 1 1561
2 51825 1 1561
2 51826 1 1562
2 51827 1 1562
2 51828 1 1562
2 51829 1 1562
2 51830 1 1565
2 51831 1 1565
2 51832 1 1565
2 51833 1 1565
2 51834 1 1565
2 51835 1 1567
2 51836 1 1567
2 51837 1 1577
2 51838 1 1577
2 51839 1 1578
2 51840 1 1578
2 51841 1 1578
2 51842 1 1579
2 51843 1 1579
2 51844 1 1579
2 51845 1 1579
2 51846 1 1579
2 51847 1 1579
2 51848 1 1579
2 51849 1 1580
2 51850 1 1580
2 51851 1 1580
2 51852 1 1580
2 51853 1 1580
2 51854 1 1580
2 51855 1 1580
2 51856 1 1580
2 51857 1 1580
2 51858 1 1580
2 51859 1 1580
2 51860 1 1580
2 51861 1 1580
2 51862 1 1580
2 51863 1 1581
2 51864 1 1581
2 51865 1 1581
2 51866 1 1581
2 51867 1 1581
2 51868 1 1581
2 51869 1 1582
2 51870 1 1582
2 51871 1 1582
2 51872 1 1582
2 51873 1 1582
2 51874 1 1582
2 51875 1 1582
2 51876 1 1582
2 51877 1 1583
2 51878 1 1583
2 51879 1 1583
2 51880 1 1583
2 51881 1 1583
2 51882 1 1583
2 51883 1 1583
2 51884 1 1583
2 51885 1 1583
2 51886 1 1583
2 51887 1 1583
2 51888 1 1583
2 51889 1 1583
2 51890 1 1583
2 51891 1 1583
2 51892 1 1583
2 51893 1 1583
2 51894 1 1586
2 51895 1 1586
2 51896 1 1586
2 51897 1 1586
2 51898 1 1587
2 51899 1 1587
2 51900 1 1587
2 51901 1 1587
2 51902 1 1589
2 51903 1 1589
2 51904 1 1602
2 51905 1 1602
2 51906 1 1603
2 51907 1 1603
2 51908 1 1603
2 51909 1 1603
2 51910 1 1603
2 51911 1 1603
2 51912 1 1603
2 51913 1 1603
2 51914 1 1603
2 51915 1 1603
2 51916 1 1603
2 51917 1 1603
2 51918 1 1603
2 51919 1 1603
2 51920 1 1603
2 51921 1 1603
2 51922 1 1603
2 51923 1 1603
2 51924 1 1603
2 51925 1 1603
2 51926 1 1603
2 51927 1 1603
2 51928 1 1603
2 51929 1 1603
2 51930 1 1603
2 51931 1 1603
2 51932 1 1603
2 51933 1 1603
2 51934 1 1603
2 51935 1 1603
2 51936 1 1603
2 51937 1 1603
2 51938 1 1603
2 51939 1 1604
2 51940 1 1604
2 51941 1 1604
2 51942 1 1608
2 51943 1 1608
2 51944 1 1609
2 51945 1 1609
2 51946 1 1609
2 51947 1 1609
2 51948 1 1610
2 51949 1 1610
2 51950 1 1610
2 51951 1 1610
2 51952 1 1611
2 51953 1 1611
2 51954 1 1611
2 51955 1 1611
2 51956 1 1612
2 51957 1 1612
2 51958 1 1612
2 51959 1 1612
2 51960 1 1612
2 51961 1 1612
2 51962 1 1613
2 51963 1 1613
2 51964 1 1613
2 51965 1 1614
2 51966 1 1614
2 51967 1 1614
2 51968 1 1614
2 51969 1 1627
2 51970 1 1627
2 51971 1 1627
2 51972 1 1627
2 51973 1 1627
2 51974 1 1627
2 51975 1 1627
2 51976 1 1627
2 51977 1 1627
2 51978 1 1627
2 51979 1 1627
2 51980 1 1629
2 51981 1 1629
2 51982 1 1629
2 51983 1 1629
2 51984 1 1629
2 51985 1 1629
2 51986 1 1629
2 51987 1 1629
2 51988 1 1629
2 51989 1 1629
2 51990 1 1629
2 51991 1 1629
2 51992 1 1629
2 51993 1 1629
2 51994 1 1629
2 51995 1 1629
2 51996 1 1629
2 51997 1 1629
2 51998 1 1629
2 51999 1 1629
2 52000 1 1629
2 52001 1 1629
2 52002 1 1629
2 52003 1 1629
2 52004 1 1629
2 52005 1 1629
2 52006 1 1629
2 52007 1 1629
2 52008 1 1629
2 52009 1 1629
2 52010 1 1629
2 52011 1 1629
2 52012 1 1629
2 52013 1 1629
2 52014 1 1629
2 52015 1 1629
2 52016 1 1630
2 52017 1 1630
2 52018 1 1630
2 52019 1 1630
2 52020 1 1630
2 52021 1 1630
2 52022 1 1630
2 52023 1 1630
2 52024 1 1630
2 52025 1 1630
2 52026 1 1630
2 52027 1 1630
2 52028 1 1630
2 52029 1 1630
2 52030 1 1630
2 52031 1 1630
2 52032 1 1630
2 52033 1 1630
2 52034 1 1630
2 52035 1 1630
2 52036 1 1631
2 52037 1 1631
2 52038 1 1631
2 52039 1 1631
2 52040 1 1632
2 52041 1 1632
2 52042 1 1632
2 52043 1 1632
2 52044 1 1632
2 52045 1 1633
2 52046 1 1633
2 52047 1 1634
2 52048 1 1634
2 52049 1 1634
2 52050 1 1634
2 52051 1 1634
2 52052 1 1634
2 52053 1 1634
2 52054 1 1634
2 52055 1 1634
2 52056 1 1634
2 52057 1 1634
2 52058 1 1634
2 52059 1 1634
2 52060 1 1636
2 52061 1 1636
2 52062 1 1637
2 52063 1 1637
2 52064 1 1637
2 52065 1 1637
2 52066 1 1637
2 52067 1 1637
2 52068 1 1637
2 52069 1 1637
2 52070 1 1637
2 52071 1 1638
2 52072 1 1638
2 52073 1 1638
2 52074 1 1638
2 52075 1 1638
2 52076 1 1639
2 52077 1 1639
2 52078 1 1640
2 52079 1 1640
2 52080 1 1640
2 52081 1 1640
2 52082 1 1642
2 52083 1 1642
2 52084 1 1642
2 52085 1 1644
2 52086 1 1644
2 52087 1 1647
2 52088 1 1647
2 52089 1 1647
2 52090 1 1648
2 52091 1 1648
2 52092 1 1648
2 52093 1 1648
2 52094 1 1648
2 52095 1 1648
2 52096 1 1648
2 52097 1 1648
2 52098 1 1648
2 52099 1 1648
2 52100 1 1648
2 52101 1 1648
2 52102 1 1648
2 52103 1 1648
2 52104 1 1648
2 52105 1 1648
2 52106 1 1648
2 52107 1 1648
2 52108 1 1648
2 52109 1 1648
2 52110 1 1648
2 52111 1 1648
2 52112 1 1648
2 52113 1 1648
2 52114 1 1650
2 52115 1 1650
2 52116 1 1651
2 52117 1 1651
2 52118 1 1651
2 52119 1 1652
2 52120 1 1652
2 52121 1 1657
2 52122 1 1657
2 52123 1 1657
2 52124 1 1657
2 52125 1 1657
2 52126 1 1657
2 52127 1 1657
2 52128 1 1657
2 52129 1 1668
2 52130 1 1668
2 52131 1 1668
2 52132 1 1668
2 52133 1 1668
2 52134 1 1668
2 52135 1 1668
2 52136 1 1668
2 52137 1 1668
2 52138 1 1671
2 52139 1 1671
2 52140 1 1671
2 52141 1 1671
2 52142 1 1671
2 52143 1 1671
2 52144 1 1671
2 52145 1 1671
2 52146 1 1671
2 52147 1 1671
2 52148 1 1672
2 52149 1 1672
2 52150 1 1672
2 52151 1 1674
2 52152 1 1674
2 52153 1 1674
2 52154 1 1674
2 52155 1 1674
2 52156 1 1674
2 52157 1 1674
2 52158 1 1674
2 52159 1 1674
2 52160 1 1674
2 52161 1 1675
2 52162 1 1675
2 52163 1 1675
2 52164 1 1675
2 52165 1 1675
2 52166 1 1675
2 52167 1 1675
2 52168 1 1675
2 52169 1 1683
2 52170 1 1683
2 52171 1 1683
2 52172 1 1683
2 52173 1 1683
2 52174 1 1683
2 52175 1 1683
2 52176 1 1683
2 52177 1 1683
2 52178 1 1683
2 52179 1 1683
2 52180 1 1683
2 52181 1 1683
2 52182 1 1683
2 52183 1 1683
2 52184 1 1683
2 52185 1 1683
2 52186 1 1683
2 52187 1 1683
2 52188 1 1683
2 52189 1 1683
2 52190 1 1683
2 52191 1 1683
2 52192 1 1685
2 52193 1 1685
2 52194 1 1685
2 52195 1 1685
2 52196 1 1685
2 52197 1 1686
2 52198 1 1686
2 52199 1 1686
2 52200 1 1686
2 52201 1 1686
2 52202 1 1697
2 52203 1 1697
2 52204 1 1697
2 52205 1 1697
2 52206 1 1697
2 52207 1 1697
2 52208 1 1697
2 52209 1 1697
2 52210 1 1702
2 52211 1 1702
2 52212 1 1702
2 52213 1 1702
2 52214 1 1702
2 52215 1 1702
2 52216 1 1703
2 52217 1 1703
2 52218 1 1703
2 52219 1 1703
2 52220 1 1703
2 52221 1 1703
2 52222 1 1704
2 52223 1 1704
2 52224 1 1708
2 52225 1 1708
2 52226 1 1708
2 52227 1 1708
2 52228 1 1708
2 52229 1 1708
2 52230 1 1708
2 52231 1 1708
2 52232 1 1708
2 52233 1 1708
2 52234 1 1708
2 52235 1 1708
2 52236 1 1709
2 52237 1 1709
2 52238 1 1709
2 52239 1 1709
2 52240 1 1709
2 52241 1 1709
2 52242 1 1709
2 52243 1 1709
2 52244 1 1709
2 52245 1 1709
2 52246 1 1710
2 52247 1 1710
2 52248 1 1710
2 52249 1 1711
2 52250 1 1711
2 52251 1 1711
2 52252 1 1712
2 52253 1 1712
2 52254 1 1712
2 52255 1 1712
2 52256 1 1712
2 52257 1 1713
2 52258 1 1713
2 52259 1 1713
2 52260 1 1713
2 52261 1 1713
2 52262 1 1713
2 52263 1 1713
2 52264 1 1714
2 52265 1 1714
2 52266 1 1714
2 52267 1 1714
2 52268 1 1714
2 52269 1 1714
2 52270 1 1714
2 52271 1 1716
2 52272 1 1716
2 52273 1 1716
2 52274 1 1716
2 52275 1 1716
2 52276 1 1718
2 52277 1 1718
2 52278 1 1720
2 52279 1 1720
2 52280 1 1725
2 52281 1 1725
2 52282 1 1725
2 52283 1 1725
2 52284 1 1725
2 52285 1 1725
2 52286 1 1725
2 52287 1 1725
2 52288 1 1725
2 52289 1 1725
2 52290 1 1726
2 52291 1 1726
2 52292 1 1726
2 52293 1 1726
2 52294 1 1726
2 52295 1 1729
2 52296 1 1729
2 52297 1 1732
2 52298 1 1732
2 52299 1 1732
2 52300 1 1732
2 52301 1 1732
2 52302 1 1732
2 52303 1 1734
2 52304 1 1734
2 52305 1 1734
2 52306 1 1734
2 52307 1 1735
2 52308 1 1735
2 52309 1 1736
2 52310 1 1736
2 52311 1 1736
2 52312 1 1737
2 52313 1 1737
2 52314 1 1737
2 52315 1 1742
2 52316 1 1742
2 52317 1 1742
2 52318 1 1742
2 52319 1 1742
2 52320 1 1742
2 52321 1 1742
2 52322 1 1742
2 52323 1 1742
2 52324 1 1742
2 52325 1 1742
2 52326 1 1742
2 52327 1 1742
2 52328 1 1742
2 52329 1 1742
2 52330 1 1742
2 52331 1 1742
2 52332 1 1742
2 52333 1 1742
2 52334 1 1742
2 52335 1 1743
2 52336 1 1743
2 52337 1 1743
2 52338 1 1743
2 52339 1 1743
2 52340 1 1743
2 52341 1 1744
2 52342 1 1744
2 52343 1 1744
2 52344 1 1744
2 52345 1 1744
2 52346 1 1745
2 52347 1 1745
2 52348 1 1745
2 52349 1 1745
2 52350 1 1745
2 52351 1 1745
2 52352 1 1745
2 52353 1 1745
2 52354 1 1752
2 52355 1 1752
2 52356 1 1752
2 52357 1 1752
2 52358 1 1752
2 52359 1 1752
2 52360 1 1752
2 52361 1 1752
2 52362 1 1752
2 52363 1 1752
2 52364 1 1753
2 52365 1 1753
2 52366 1 1754
2 52367 1 1754
2 52368 1 1759
2 52369 1 1759
2 52370 1 1760
2 52371 1 1760
2 52372 1 1760
2 52373 1 1760
2 52374 1 1760
2 52375 1 1760
2 52376 1 1761
2 52377 1 1761
2 52378 1 1770
2 52379 1 1770
2 52380 1 1770
2 52381 1 1770
2 52382 1 1770
2 52383 1 1770
2 52384 1 1770
2 52385 1 1770
2 52386 1 1770
2 52387 1 1783
2 52388 1 1783
2 52389 1 1783
2 52390 1 1783
2 52391 1 1783
2 52392 1 1783
2 52393 1 1783
2 52394 1 1783
2 52395 1 1783
2 52396 1 1783
2 52397 1 1783
2 52398 1 1783
2 52399 1 1783
2 52400 1 1783
2 52401 1 1783
2 52402 1 1784
2 52403 1 1784
2 52404 1 1784
2 52405 1 1784
2 52406 1 1784
2 52407 1 1784
2 52408 1 1784
2 52409 1 1784
2 52410 1 1784
2 52411 1 1785
2 52412 1 1785
2 52413 1 1785
2 52414 1 1785
2 52415 1 1785
2 52416 1 1785
2 52417 1 1786
2 52418 1 1786
2 52419 1 1786
2 52420 1 1786
2 52421 1 1786
2 52422 1 1786
2 52423 1 1786
2 52424 1 1786
2 52425 1 1786
2 52426 1 1786
2 52427 1 1786
2 52428 1 1786
2 52429 1 1799
2 52430 1 1799
2 52431 1 1799
2 52432 1 1799
2 52433 1 1799
2 52434 1 1799
2 52435 1 1799
2 52436 1 1799
2 52437 1 1799
2 52438 1 1799
2 52439 1 1799
2 52440 1 1799
2 52441 1 1799
2 52442 1 1799
2 52443 1 1799
2 52444 1 1799
2 52445 1 1799
2 52446 1 1799
2 52447 1 1799
2 52448 1 1799
2 52449 1 1799
2 52450 1 1799
2 52451 1 1799
2 52452 1 1799
2 52453 1 1799
2 52454 1 1799
2 52455 1 1799
2 52456 1 1799
2 52457 1 1799
2 52458 1 1799
2 52459 1 1799
2 52460 1 1799
2 52461 1 1799
2 52462 1 1799
2 52463 1 1799
2 52464 1 1799
2 52465 1 1800
2 52466 1 1800
2 52467 1 1800
2 52468 1 1801
2 52469 1 1801
2 52470 1 1801
2 52471 1 1801
2 52472 1 1801
2 52473 1 1802
2 52474 1 1802
2 52475 1 1802
2 52476 1 1802
2 52477 1 1803
2 52478 1 1803
2 52479 1 1803
2 52480 1 1803
2 52481 1 1803
2 52482 1 1804
2 52483 1 1804
2 52484 1 1804
2 52485 1 1804
2 52486 1 1804
2 52487 1 1804
2 52488 1 1804
2 52489 1 1804
2 52490 1 1805
2 52491 1 1805
2 52492 1 1805
2 52493 1 1805
2 52494 1 1805
2 52495 1 1805
2 52496 1 1805
2 52497 1 1805
2 52498 1 1805
2 52499 1 1805
2 52500 1 1805
2 52501 1 1805
2 52502 1 1805
2 52503 1 1805
2 52504 1 1807
2 52505 1 1807
2 52506 1 1814
2 52507 1 1814
2 52508 1 1814
2 52509 1 1814
2 52510 1 1814
2 52511 1 1814
2 52512 1 1814
2 52513 1 1814
2 52514 1 1814
2 52515 1 1814
2 52516 1 1814
2 52517 1 1814
2 52518 1 1817
2 52519 1 1817
2 52520 1 1817
2 52521 1 1822
2 52522 1 1822
2 52523 1 1828
2 52524 1 1828
2 52525 1 1828
2 52526 1 1828
2 52527 1 1828
2 52528 1 1828
2 52529 1 1828
2 52530 1 1828
2 52531 1 1840
2 52532 1 1840
2 52533 1 1840
2 52534 1 1840
2 52535 1 1840
2 52536 1 1840
2 52537 1 1840
2 52538 1 1840
2 52539 1 1841
2 52540 1 1841
2 52541 1 1841
2 52542 1 1842
2 52543 1 1842
2 52544 1 1843
2 52545 1 1843
2 52546 1 1850
2 52547 1 1850
2 52548 1 1850
2 52549 1 1850
2 52550 1 1850
2 52551 1 1850
2 52552 1 1850
2 52553 1 1850
2 52554 1 1851
2 52555 1 1851
2 52556 1 1851
2 52557 1 1851
2 52558 1 1852
2 52559 1 1852
2 52560 1 1856
2 52561 1 1856
2 52562 1 1856
2 52563 1 1856
2 52564 1 1870
2 52565 1 1870
2 52566 1 1870
2 52567 1 1870
2 52568 1 1870
2 52569 1 1881
2 52570 1 1881
2 52571 1 1881
2 52572 1 1881
2 52573 1 1881
2 52574 1 1881
2 52575 1 1882
2 52576 1 1882
2 52577 1 1882
2 52578 1 1883
2 52579 1 1883
2 52580 1 1886
2 52581 1 1886
2 52582 1 1886
2 52583 1 1886
2 52584 1 1886
2 52585 1 1886
2 52586 1 1886
2 52587 1 1886
2 52588 1 1886
2 52589 1 1886
2 52590 1 1887
2 52591 1 1887
2 52592 1 1887
2 52593 1 1889
2 52594 1 1889
2 52595 1 1891
2 52596 1 1891
2 52597 1 1898
2 52598 1 1898
2 52599 1 1898
2 52600 1 1898
2 52601 1 1900
2 52602 1 1900
2 52603 1 1900
2 52604 1 1900
2 52605 1 1900
2 52606 1 1900
2 52607 1 1900
2 52608 1 1900
2 52609 1 1900
2 52610 1 1900
2 52611 1 1900
2 52612 1 1900
2 52613 1 1900
2 52614 1 1900
2 52615 1 1900
2 52616 1 1900
2 52617 1 1900
2 52618 1 1901
2 52619 1 1901
2 52620 1 1901
2 52621 1 1901
2 52622 1 1902
2 52623 1 1902
2 52624 1 1902
2 52625 1 1902
2 52626 1 1902
2 52627 1 1902
2 52628 1 1902
2 52629 1 1911
2 52630 1 1911
2 52631 1 1911
2 52632 1 1911
2 52633 1 1911
2 52634 1 1911
2 52635 1 1911
2 52636 1 1911
2 52637 1 1911
2 52638 1 1911
2 52639 1 1911
2 52640 1 1911
2 52641 1 1911
2 52642 1 1911
2 52643 1 1911
2 52644 1 1911
2 52645 1 1911
2 52646 1 1911
2 52647 1 1912
2 52648 1 1912
2 52649 1 1912
2 52650 1 1912
2 52651 1 1913
2 52652 1 1913
2 52653 1 1914
2 52654 1 1914
2 52655 1 1914
2 52656 1 1914
2 52657 1 1917
2 52658 1 1917
2 52659 1 1928
2 52660 1 1928
2 52661 1 1928
2 52662 1 1928
2 52663 1 1928
2 52664 1 1932
2 52665 1 1932
2 52666 1 1935
2 52667 1 1935
2 52668 1 1935
2 52669 1 1935
2 52670 1 1935
2 52671 1 1936
2 52672 1 1936
2 52673 1 1937
2 52674 1 1937
2 52675 1 1937
2 52676 1 1937
2 52677 1 1937
2 52678 1 1937
2 52679 1 1938
2 52680 1 1938
2 52681 1 1938
2 52682 1 1938
2 52683 1 1938
2 52684 1 1939
2 52685 1 1939
2 52686 1 1939
2 52687 1 1939
2 52688 1 1939
2 52689 1 1939
2 52690 1 1939
2 52691 1 1939
2 52692 1 1939
2 52693 1 1939
2 52694 1 1939
2 52695 1 1939
2 52696 1 1939
2 52697 1 1939
2 52698 1 1939
2 52699 1 1940
2 52700 1 1940
2 52701 1 1940
2 52702 1 1940
2 52703 1 1940
2 52704 1 1940
2 52705 1 1948
2 52706 1 1948
2 52707 1 1948
2 52708 1 1948
2 52709 1 1948
2 52710 1 1948
2 52711 1 1948
2 52712 1 1950
2 52713 1 1950
2 52714 1 1953
2 52715 1 1953
2 52716 1 1953
2 52717 1 1953
2 52718 1 1960
2 52719 1 1960
2 52720 1 1960
2 52721 1 1972
2 52722 1 1972
2 52723 1 1972
2 52724 1 1973
2 52725 1 1973
2 52726 1 1973
2 52727 1 1973
2 52728 1 1975
2 52729 1 1975
2 52730 1 1975
2 52731 1 1975
2 52732 1 1975
2 52733 1 1978
2 52734 1 1978
2 52735 1 1993
2 52736 1 1993
2 52737 1 1996
2 52738 1 1996
2 52739 1 1996
2 52740 1 1996
2 52741 1 1996
2 52742 1 1996
2 52743 1 1996
2 52744 1 2006
2 52745 1 2006
2 52746 1 2006
2 52747 1 2007
2 52748 1 2007
2 52749 1 2007
2 52750 1 2010
2 52751 1 2010
2 52752 1 2011
2 52753 1 2011
2 52754 1 2031
2 52755 1 2031
2 52756 1 2031
2 52757 1 2033
2 52758 1 2033
2 52759 1 2033
2 52760 1 2033
2 52761 1 2033
2 52762 1 2034
2 52763 1 2034
2 52764 1 2034
2 52765 1 2037
2 52766 1 2037
2 52767 1 2038
2 52768 1 2038
2 52769 1 2038
2 52770 1 2038
2 52771 1 2038
2 52772 1 2038
2 52773 1 2041
2 52774 1 2041
2 52775 1 2041
2 52776 1 2041
2 52777 1 2041
2 52778 1 2042
2 52779 1 2042
2 52780 1 2042
2 52781 1 2043
2 52782 1 2043
2 52783 1 2049
2 52784 1 2049
2 52785 1 2049
2 52786 1 2049
2 52787 1 2049
2 52788 1 2050
2 52789 1 2050
2 52790 1 2050
2 52791 1 2050
2 52792 1 2050
2 52793 1 2058
2 52794 1 2058
2 52795 1 2058
2 52796 1 2058
2 52797 1 2058
2 52798 1 2066
2 52799 1 2066
2 52800 1 2066
2 52801 1 2066
2 52802 1 2066
2 52803 1 2066
2 52804 1 2066
2 52805 1 2066
2 52806 1 2067
2 52807 1 2067
2 52808 1 2067
2 52809 1 2067
2 52810 1 2067
2 52811 1 2067
2 52812 1 2067
2 52813 1 2067
2 52814 1 2067
2 52815 1 2067
2 52816 1 2067
2 52817 1 2068
2 52818 1 2068
2 52819 1 2069
2 52820 1 2069
2 52821 1 2082
2 52822 1 2082
2 52823 1 2082
2 52824 1 2083
2 52825 1 2083
2 52826 1 2097
2 52827 1 2097
2 52828 1 2106
2 52829 1 2106
2 52830 1 2107
2 52831 1 2107
2 52832 1 2118
2 52833 1 2118
2 52834 1 2118
2 52835 1 2118
2 52836 1 2119
2 52837 1 2119
2 52838 1 2120
2 52839 1 2120
2 52840 1 2128
2 52841 1 2128
2 52842 1 2132
2 52843 1 2132
2 52844 1 2132
2 52845 1 2133
2 52846 1 2133
2 52847 1 2133
2 52848 1 2133
2 52849 1 2133
2 52850 1 2133
2 52851 1 2135
2 52852 1 2135
2 52853 1 2143
2 52854 1 2143
2 52855 1 2143
2 52856 1 2143
2 52857 1 2143
2 52858 1 2143
2 52859 1 2143
2 52860 1 2143
2 52861 1 2145
2 52862 1 2145
2 52863 1 2145
2 52864 1 2145
2 52865 1 2145
2 52866 1 2145
2 52867 1 2145
2 52868 1 2145
2 52869 1 2145
2 52870 1 2145
2 52871 1 2145
2 52872 1 2145
2 52873 1 2147
2 52874 1 2147
2 52875 1 2147
2 52876 1 2147
2 52877 1 2147
2 52878 1 2147
2 52879 1 2147
2 52880 1 2151
2 52881 1 2151
2 52882 1 2159
2 52883 1 2159
2 52884 1 2159
2 52885 1 2159
2 52886 1 2159
2 52887 1 2159
2 52888 1 2160
2 52889 1 2160
2 52890 1 2161
2 52891 1 2161
2 52892 1 2166
2 52893 1 2166
2 52894 1 2166
2 52895 1 2166
2 52896 1 2166
2 52897 1 2166
2 52898 1 2170
2 52899 1 2170
2 52900 1 2170
2 52901 1 2170
2 52902 1 2170
2 52903 1 2170
2 52904 1 2170
2 52905 1 2170
2 52906 1 2170
2 52907 1 2170
2 52908 1 2170
2 52909 1 2170
2 52910 1 2170
2 52911 1 2170
2 52912 1 2170
2 52913 1 2170
2 52914 1 2170
2 52915 1 2170
2 52916 1 2170
2 52917 1 2170
2 52918 1 2170
2 52919 1 2170
2 52920 1 2170
2 52921 1 2170
2 52922 1 2170
2 52923 1 2170
2 52924 1 2170
2 52925 1 2170
2 52926 1 2170
2 52927 1 2170
2 52928 1 2170
2 52929 1 2170
2 52930 1 2170
2 52931 1 2170
2 52932 1 2170
2 52933 1 2170
2 52934 1 2170
2 52935 1 2170
2 52936 1 2170
2 52937 1 2170
2 52938 1 2170
2 52939 1 2170
2 52940 1 2170
2 52941 1 2170
2 52942 1 2170
2 52943 1 2170
2 52944 1 2170
2 52945 1 2170
2 52946 1 2170
2 52947 1 2170
2 52948 1 2170
2 52949 1 2170
2 52950 1 2170
2 52951 1 2171
2 52952 1 2171
2 52953 1 2171
2 52954 1 2171
2 52955 1 2172
2 52956 1 2172
2 52957 1 2172
2 52958 1 2172
2 52959 1 2172
2 52960 1 2172
2 52961 1 2172
2 52962 1 2172
2 52963 1 2172
2 52964 1 2172
2 52965 1 2172
2 52966 1 2173
2 52967 1 2173
2 52968 1 2173
2 52969 1 2175
2 52970 1 2175
2 52971 1 2175
2 52972 1 2176
2 52973 1 2176
2 52974 1 2186
2 52975 1 2186
2 52976 1 2186
2 52977 1 2186
2 52978 1 2186
2 52979 1 2186
2 52980 1 2188
2 52981 1 2188
2 52982 1 2191
2 52983 1 2191
2 52984 1 2191
2 52985 1 2192
2 52986 1 2192
2 52987 1 2192
2 52988 1 2192
2 52989 1 2193
2 52990 1 2193
2 52991 1 2193
2 52992 1 2194
2 52993 1 2194
2 52994 1 2195
2 52995 1 2195
2 52996 1 2198
2 52997 1 2198
2 52998 1 2198
2 52999 1 2200
2 53000 1 2200
2 53001 1 2205
2 53002 1 2205
2 53003 1 2205
2 53004 1 2205
2 53005 1 2205
2 53006 1 2205
2 53007 1 2212
2 53008 1 2212
2 53009 1 2212
2 53010 1 2212
2 53011 1 2212
2 53012 1 2212
2 53013 1 2212
2 53014 1 2213
2 53015 1 2213
2 53016 1 2218
2 53017 1 2218
2 53018 1 2225
2 53019 1 2225
2 53020 1 2231
2 53021 1 2231
2 53022 1 2233
2 53023 1 2233
2 53024 1 2233
2 53025 1 2237
2 53026 1 2237
2 53027 1 2241
2 53028 1 2241
2 53029 1 2252
2 53030 1 2252
2 53031 1 2252
2 53032 1 2252
2 53033 1 2252
2 53034 1 2252
2 53035 1 2252
2 53036 1 2252
2 53037 1 2252
2 53038 1 2254
2 53039 1 2254
2 53040 1 2255
2 53041 1 2255
2 53042 1 2257
2 53043 1 2257
2 53044 1 2259
2 53045 1 2259
2 53046 1 2268
2 53047 1 2268
2 53048 1 2268
2 53049 1 2268
2 53050 1 2269
2 53051 1 2269
2 53052 1 2270
2 53053 1 2270
2 53054 1 2289
2 53055 1 2289
2 53056 1 2289
2 53057 1 2289
2 53058 1 2290
2 53059 1 2290
2 53060 1 2290
2 53061 1 2290
2 53062 1 2290
2 53063 1 2290
2 53064 1 2290
2 53065 1 2290
2 53066 1 2290
2 53067 1 2290
2 53068 1 2291
2 53069 1 2291
2 53070 1 2298
2 53071 1 2298
2 53072 1 2298
2 53073 1 2298
2 53074 1 2298
2 53075 1 2298
2 53076 1 2298
2 53077 1 2298
2 53078 1 2298
2 53079 1 2299
2 53080 1 2299
2 53081 1 2299
2 53082 1 2299
2 53083 1 2299
2 53084 1 2299
2 53085 1 2300
2 53086 1 2300
2 53087 1 2300
2 53088 1 2300
2 53089 1 2300
2 53090 1 2300
2 53091 1 2300
2 53092 1 2301
2 53093 1 2301
2 53094 1 2301
2 53095 1 2301
2 53096 1 2301
2 53097 1 2301
2 53098 1 2301
2 53099 1 2301
2 53100 1 2309
2 53101 1 2309
2 53102 1 2310
2 53103 1 2310
2 53104 1 2311
2 53105 1 2311
2 53106 1 2333
2 53107 1 2333
2 53108 1 2336
2 53109 1 2336
2 53110 1 2344
2 53111 1 2344
2 53112 1 2344
2 53113 1 2363
2 53114 1 2363
2 53115 1 2363
2 53116 1 2364
2 53117 1 2364
2 53118 1 2367
2 53119 1 2367
2 53120 1 2368
2 53121 1 2368
2 53122 1 2378
2 53123 1 2378
2 53124 1 2378
2 53125 1 2378
2 53126 1 2378
2 53127 1 2378
2 53128 1 2381
2 53129 1 2381
2 53130 1 2381
2 53131 1 2381
2 53132 1 2381
2 53133 1 2384
2 53134 1 2384
2 53135 1 2384
2 53136 1 2384
2 53137 1 2384
2 53138 1 2384
2 53139 1 2384
2 53140 1 2384
2 53141 1 2384
2 53142 1 2384
2 53143 1 2384
2 53144 1 2385
2 53145 1 2385
2 53146 1 2385
2 53147 1 2385
2 53148 1 2385
2 53149 1 2394
2 53150 1 2394
2 53151 1 2395
2 53152 1 2395
2 53153 1 2395
2 53154 1 2395
2 53155 1 2397
2 53156 1 2397
2 53157 1 2398
2 53158 1 2398
2 53159 1 2401
2 53160 1 2401
2 53161 1 2404
2 53162 1 2404
2 53163 1 2404
2 53164 1 2404
2 53165 1 2405
2 53166 1 2405
2 53167 1 2408
2 53168 1 2408
2 53169 1 2408
2 53170 1 2409
2 53171 1 2409
2 53172 1 2410
2 53173 1 2410
2 53174 1 2410
2 53175 1 2410
2 53176 1 2410
2 53177 1 2410
2 53178 1 2410
2 53179 1 2410
2 53180 1 2410
2 53181 1 2410
2 53182 1 2410
2 53183 1 2410
2 53184 1 2424
2 53185 1 2424
2 53186 1 2424
2 53187 1 2424
2 53188 1 2424
2 53189 1 2424
2 53190 1 2424
2 53191 1 2424
2 53192 1 2425
2 53193 1 2425
2 53194 1 2440
2 53195 1 2440
2 53196 1 2440
2 53197 1 2440
2 53198 1 2441
2 53199 1 2441
2 53200 1 2441
2 53201 1 2446
2 53202 1 2446
2 53203 1 2446
2 53204 1 2446
2 53205 1 2446
2 53206 1 2446
2 53207 1 2446
2 53208 1 2446
2 53209 1 2446
2 53210 1 2446
2 53211 1 2446
2 53212 1 2446
2 53213 1 2446
2 53214 1 2446
2 53215 1 2446
2 53216 1 2446
2 53217 1 2446
2 53218 1 2446
2 53219 1 2447
2 53220 1 2447
2 53221 1 2447
2 53222 1 2449
2 53223 1 2449
2 53224 1 2454
2 53225 1 2454
2 53226 1 2454
2 53227 1 2454
2 53228 1 2454
2 53229 1 2454
2 53230 1 2454
2 53231 1 2454
2 53232 1 2454
2 53233 1 2454
2 53234 1 2454
2 53235 1 2454
2 53236 1 2454
2 53237 1 2454
2 53238 1 2454
2 53239 1 2454
2 53240 1 2454
2 53241 1 2456
2 53242 1 2456
2 53243 1 2456
2 53244 1 2456
2 53245 1 2456
2 53246 1 2457
2 53247 1 2457
2 53248 1 2459
2 53249 1 2459
2 53250 1 2459
2 53251 1 2459
2 53252 1 2459
2 53253 1 2459
2 53254 1 2459
2 53255 1 2460
2 53256 1 2460
2 53257 1 2460
2 53258 1 2460
2 53259 1 2460
2 53260 1 2460
2 53261 1 2460
2 53262 1 2460
2 53263 1 2460
2 53264 1 2460
2 53265 1 2460
2 53266 1 2460
2 53267 1 2460
2 53268 1 2460
2 53269 1 2460
2 53270 1 2460
2 53271 1 2460
2 53272 1 2468
2 53273 1 2468
2 53274 1 2468
2 53275 1 2468
2 53276 1 2468
2 53277 1 2468
2 53278 1 2468
2 53279 1 2468
2 53280 1 2468
2 53281 1 2468
2 53282 1 2468
2 53283 1 2468
2 53284 1 2468
2 53285 1 2468
2 53286 1 2468
2 53287 1 2468
2 53288 1 2468
2 53289 1 2468
2 53290 1 2468
2 53291 1 2468
2 53292 1 2468
2 53293 1 2468
2 53294 1 2468
2 53295 1 2468
2 53296 1 2468
2 53297 1 2468
2 53298 1 2468
2 53299 1 2469
2 53300 1 2469
2 53301 1 2470
2 53302 1 2470
2 53303 1 2470
2 53304 1 2470
2 53305 1 2470
2 53306 1 2470
2 53307 1 2470
2 53308 1 2471
2 53309 1 2471
2 53310 1 2472
2 53311 1 2472
2 53312 1 2472
2 53313 1 2472
2 53314 1 2472
2 53315 1 2472
2 53316 1 2473
2 53317 1 2473
2 53318 1 2473
2 53319 1 2473
2 53320 1 2473
2 53321 1 2473
2 53322 1 2473
2 53323 1 2473
2 53324 1 2473
2 53325 1 2473
2 53326 1 2482
2 53327 1 2482
2 53328 1 2482
2 53329 1 2482
2 53330 1 2482
2 53331 1 2482
2 53332 1 2482
2 53333 1 2482
2 53334 1 2482
2 53335 1 2482
2 53336 1 2482
2 53337 1 2490
2 53338 1 2490
2 53339 1 2490
2 53340 1 2490
2 53341 1 2490
2 53342 1 2490
2 53343 1 2490
2 53344 1 2490
2 53345 1 2490
2 53346 1 2500
2 53347 1 2500
2 53348 1 2506
2 53349 1 2506
2 53350 1 2507
2 53351 1 2507
2 53352 1 2513
2 53353 1 2513
2 53354 1 2519
2 53355 1 2519
2 53356 1 2519
2 53357 1 2519
2 53358 1 2519
2 53359 1 2519
2 53360 1 2519
2 53361 1 2519
2 53362 1 2520
2 53363 1 2520
2 53364 1 2521
2 53365 1 2521
2 53366 1 2521
2 53367 1 2521
2 53368 1 2521
2 53369 1 2523
2 53370 1 2523
2 53371 1 2524
2 53372 1 2524
2 53373 1 2540
2 53374 1 2540
2 53375 1 2540
2 53376 1 2544
2 53377 1 2544
2 53378 1 2551
2 53379 1 2551
2 53380 1 2551
2 53381 1 2551
2 53382 1 2551
2 53383 1 2553
2 53384 1 2553
2 53385 1 2575
2 53386 1 2575
2 53387 1 2575
2 53388 1 2575
2 53389 1 2576
2 53390 1 2576
2 53391 1 2576
2 53392 1 2576
2 53393 1 2576
2 53394 1 2576
2 53395 1 2577
2 53396 1 2577
2 53397 1 2578
2 53398 1 2578
2 53399 1 2579
2 53400 1 2579
2 53401 1 2580
2 53402 1 2580
2 53403 1 2580
2 53404 1 2584
2 53405 1 2584
2 53406 1 2585
2 53407 1 2585
2 53408 1 2585
2 53409 1 2585
2 53410 1 2586
2 53411 1 2586
2 53412 1 2586
2 53413 1 2586
2 53414 1 2592
2 53415 1 2592
2 53416 1 2592
2 53417 1 2594
2 53418 1 2594
2 53419 1 2601
2 53420 1 2601
2 53421 1 2601
2 53422 1 2601
2 53423 1 2601
2 53424 1 2601
2 53425 1 2602
2 53426 1 2602
2 53427 1 2602
2 53428 1 2610
2 53429 1 2610
2 53430 1 2610
2 53431 1 2610
2 53432 1 2610
2 53433 1 2610
2 53434 1 2610
2 53435 1 2610
2 53436 1 2610
2 53437 1 2610
2 53438 1 2611
2 53439 1 2611
2 53440 1 2611
2 53441 1 2611
2 53442 1 2612
2 53443 1 2612
2 53444 1 2620
2 53445 1 2620
2 53446 1 2620
2 53447 1 2620
2 53448 1 2620
2 53449 1 2620
2 53450 1 2620
2 53451 1 2620
2 53452 1 2620
2 53453 1 2620
2 53454 1 2620
2 53455 1 2620
2 53456 1 2620
2 53457 1 2620
2 53458 1 2620
2 53459 1 2620
2 53460 1 2620
2 53461 1 2620
2 53462 1 2620
2 53463 1 2620
2 53464 1 2620
2 53465 1 2620
2 53466 1 2620
2 53467 1 2620
2 53468 1 2620
2 53469 1 2620
2 53470 1 2622
2 53471 1 2622
2 53472 1 2622
2 53473 1 2622
2 53474 1 2622
2 53475 1 2622
2 53476 1 2622
2 53477 1 2622
2 53478 1 2622
2 53479 1 2635
2 53480 1 2635
2 53481 1 2635
2 53482 1 2635
2 53483 1 2637
2 53484 1 2637
2 53485 1 2637
2 53486 1 2639
2 53487 1 2639
2 53488 1 2639
2 53489 1 2640
2 53490 1 2640
2 53491 1 2641
2 53492 1 2641
2 53493 1 2641
2 53494 1 2641
2 53495 1 2641
2 53496 1 2641
2 53497 1 2641
2 53498 1 2641
2 53499 1 2642
2 53500 1 2642
2 53501 1 2642
2 53502 1 2652
2 53503 1 2652
2 53504 1 2653
2 53505 1 2653
2 53506 1 2653
2 53507 1 2654
2 53508 1 2654
2 53509 1 2655
2 53510 1 2655
2 53511 1 2655
2 53512 1 2655
2 53513 1 2655
2 53514 1 2655
2 53515 1 2655
2 53516 1 2655
2 53517 1 2657
2 53518 1 2657
2 53519 1 2657
2 53520 1 2657
2 53521 1 2658
2 53522 1 2658
2 53523 1 2658
2 53524 1 2660
2 53525 1 2660
2 53526 1 2660
2 53527 1 2660
2 53528 1 2660
2 53529 1 2660
2 53530 1 2660
2 53531 1 2660
2 53532 1 2660
2 53533 1 2660
2 53534 1 2660
2 53535 1 2660
2 53536 1 2660
2 53537 1 2661
2 53538 1 2661
2 53539 1 2661
2 53540 1 2661
2 53541 1 2661
2 53542 1 2661
2 53543 1 2661
2 53544 1 2661
2 53545 1 2661
2 53546 1 2661
2 53547 1 2661
2 53548 1 2661
2 53549 1 2661
2 53550 1 2668
2 53551 1 2668
2 53552 1 2672
2 53553 1 2672
2 53554 1 2673
2 53555 1 2673
2 53556 1 2673
2 53557 1 2673
2 53558 1 2673
2 53559 1 2673
2 53560 1 2673
2 53561 1 2673
2 53562 1 2673
2 53563 1 2674
2 53564 1 2674
2 53565 1 2674
2 53566 1 2674
2 53567 1 2675
2 53568 1 2675
2 53569 1 2675
2 53570 1 2676
2 53571 1 2676
2 53572 1 2678
2 53573 1 2678
2 53574 1 2678
2 53575 1 2679
2 53576 1 2679
2 53577 1 2696
2 53578 1 2696
2 53579 1 2696
2 53580 1 2696
2 53581 1 2696
2 53582 1 2696
2 53583 1 2696
2 53584 1 2696
2 53585 1 2708
2 53586 1 2708
2 53587 1 2708
2 53588 1 2709
2 53589 1 2709
2 53590 1 2713
2 53591 1 2713
2 53592 1 2713
2 53593 1 2714
2 53594 1 2714
2 53595 1 2714
2 53596 1 2714
2 53597 1 2714
2 53598 1 2714
2 53599 1 2714
2 53600 1 2714
2 53601 1 2714
2 53602 1 2714
2 53603 1 2714
2 53604 1 2715
2 53605 1 2715
2 53606 1 2715
2 53607 1 2715
2 53608 1 2715
2 53609 1 2715
2 53610 1 2715
2 53611 1 2715
2 53612 1 2715
2 53613 1 2715
2 53614 1 2715
2 53615 1 2715
2 53616 1 2715
2 53617 1 2715
2 53618 1 2716
2 53619 1 2716
2 53620 1 2724
2 53621 1 2724
2 53622 1 2724
2 53623 1 2724
2 53624 1 2724
2 53625 1 2724
2 53626 1 2724
2 53627 1 2724
2 53628 1 2724
2 53629 1 2724
2 53630 1 2724
2 53631 1 2724
2 53632 1 2724
2 53633 1 2724
2 53634 1 2724
2 53635 1 2724
2 53636 1 2724
2 53637 1 2724
2 53638 1 2724
2 53639 1 2724
2 53640 1 2724
2 53641 1 2724
2 53642 1 2724
2 53643 1 2724
2 53644 1 2724
2 53645 1 2724
2 53646 1 2724
2 53647 1 2724
2 53648 1 2724
2 53649 1 2724
2 53650 1 2724
2 53651 1 2724
2 53652 1 2724
2 53653 1 2724
2 53654 1 2724
2 53655 1 2724
2 53656 1 2724
2 53657 1 2724
2 53658 1 2724
2 53659 1 2724
2 53660 1 2724
2 53661 1 2724
2 53662 1 2724
2 53663 1 2724
2 53664 1 2724
2 53665 1 2725
2 53666 1 2725
2 53667 1 2725
2 53668 1 2725
2 53669 1 2725
2 53670 1 2725
2 53671 1 2734
2 53672 1 2734
2 53673 1 2734
2 53674 1 2734
2 53675 1 2735
2 53676 1 2735
2 53677 1 2735
2 53678 1 2736
2 53679 1 2736
2 53680 1 2736
2 53681 1 2736
2 53682 1 2736
2 53683 1 2736
2 53684 1 2736
2 53685 1 2736
2 53686 1 2736
2 53687 1 2736
2 53688 1 2736
2 53689 1 2736
2 53690 1 2737
2 53691 1 2737
2 53692 1 2737
2 53693 1 2737
2 53694 1 2737
2 53695 1 2738
2 53696 1 2738
2 53697 1 2739
2 53698 1 2739
2 53699 1 2739
2 53700 1 2739
2 53701 1 2739
2 53702 1 2739
2 53703 1 2739
2 53704 1 2739
2 53705 1 2739
2 53706 1 2739
2 53707 1 2739
2 53708 1 2739
2 53709 1 2739
2 53710 1 2739
2 53711 1 2739
2 53712 1 2740
2 53713 1 2740
2 53714 1 2744
2 53715 1 2744
2 53716 1 2747
2 53717 1 2747
2 53718 1 2747
2 53719 1 2747
2 53720 1 2747
2 53721 1 2747
2 53722 1 2747
2 53723 1 2747
2 53724 1 2747
2 53725 1 2747
2 53726 1 2747
2 53727 1 2748
2 53728 1 2748
2 53729 1 2748
2 53730 1 2749
2 53731 1 2749
2 53732 1 2750
2 53733 1 2750
2 53734 1 2754
2 53735 1 2754
2 53736 1 2764
2 53737 1 2764
2 53738 1 2764
2 53739 1 2764
2 53740 1 2765
2 53741 1 2765
2 53742 1 2765
2 53743 1 2767
2 53744 1 2767
2 53745 1 2772
2 53746 1 2772
2 53747 1 2772
2 53748 1 2772
2 53749 1 2772
2 53750 1 2773
2 53751 1 2773
2 53752 1 2773
2 53753 1 2773
2 53754 1 2773
2 53755 1 2773
2 53756 1 2773
2 53757 1 2775
2 53758 1 2775
2 53759 1 2775
2 53760 1 2775
2 53761 1 2775
2 53762 1 2775
2 53763 1 2775
2 53764 1 2775
2 53765 1 2775
2 53766 1 2775
2 53767 1 2775
2 53768 1 2775
2 53769 1 2775
2 53770 1 2775
2 53771 1 2775
2 53772 1 2775
2 53773 1 2775
2 53774 1 2775
2 53775 1 2775
2 53776 1 2775
2 53777 1 2775
2 53778 1 2775
2 53779 1 2775
2 53780 1 2775
2 53781 1 2775
2 53782 1 2775
2 53783 1 2776
2 53784 1 2776
2 53785 1 2776
2 53786 1 2777
2 53787 1 2777
2 53788 1 2777
2 53789 1 2777
2 53790 1 2777
2 53791 1 2777
2 53792 1 2779
2 53793 1 2779
2 53794 1 2779
2 53795 1 2779
2 53796 1 2780
2 53797 1 2780
2 53798 1 2781
2 53799 1 2781
2 53800 1 2788
2 53801 1 2788
2 53802 1 2791
2 53803 1 2791
2 53804 1 2791
2 53805 1 2791
2 53806 1 2791
2 53807 1 2791
2 53808 1 2791
2 53809 1 2791
2 53810 1 2791
2 53811 1 2791
2 53812 1 2791
2 53813 1 2791
2 53814 1 2791
2 53815 1 2791
2 53816 1 2791
2 53817 1 2791
2 53818 1 2791
2 53819 1 2791
2 53820 1 2791
2 53821 1 2791
2 53822 1 2791
2 53823 1 2791
2 53824 1 2791
2 53825 1 2791
2 53826 1 2791
2 53827 1 2791
2 53828 1 2791
2 53829 1 2791
2 53830 1 2791
2 53831 1 2791
2 53832 1 2791
2 53833 1 2791
2 53834 1 2791
2 53835 1 2791
2 53836 1 2791
2 53837 1 2791
2 53838 1 2791
2 53839 1 2791
2 53840 1 2791
2 53841 1 2791
2 53842 1 2791
2 53843 1 2791
2 53844 1 2791
2 53845 1 2792
2 53846 1 2792
2 53847 1 2792
2 53848 1 2793
2 53849 1 2793
2 53850 1 2793
2 53851 1 2793
2 53852 1 2793
2 53853 1 2794
2 53854 1 2794
2 53855 1 2795
2 53856 1 2795
2 53857 1 2795
2 53858 1 2795
2 53859 1 2795
2 53860 1 2807
2 53861 1 2807
2 53862 1 2807
2 53863 1 2807
2 53864 1 2807
2 53865 1 2807
2 53866 1 2807
2 53867 1 2807
2 53868 1 2807
2 53869 1 2807
2 53870 1 2807
2 53871 1 2807
2 53872 1 2807
2 53873 1 2807
2 53874 1 2807
2 53875 1 2807
2 53876 1 2807
2 53877 1 2807
2 53878 1 2807
2 53879 1 2807
2 53880 1 2807
2 53881 1 2807
2 53882 1 2807
2 53883 1 2807
2 53884 1 2807
2 53885 1 2807
2 53886 1 2807
2 53887 1 2807
2 53888 1 2807
2 53889 1 2807
2 53890 1 2807
2 53891 1 2807
2 53892 1 2807
2 53893 1 2807
2 53894 1 2807
2 53895 1 2807
2 53896 1 2807
2 53897 1 2807
2 53898 1 2807
2 53899 1 2807
2 53900 1 2807
2 53901 1 2807
2 53902 1 2807
2 53903 1 2807
2 53904 1 2807
2 53905 1 2807
2 53906 1 2807
2 53907 1 2807
2 53908 1 2807
2 53909 1 2807
2 53910 1 2807
2 53911 1 2807
2 53912 1 2807
2 53913 1 2807
2 53914 1 2807
2 53915 1 2807
2 53916 1 2807
2 53917 1 2807
2 53918 1 2807
2 53919 1 2807
2 53920 1 2807
2 53921 1 2807
2 53922 1 2807
2 53923 1 2807
2 53924 1 2807
2 53925 1 2807
2 53926 1 2807
2 53927 1 2807
2 53928 1 2807
2 53929 1 2807
2 53930 1 2807
2 53931 1 2807
2 53932 1 2807
2 53933 1 2807
2 53934 1 2809
2 53935 1 2809
2 53936 1 2809
2 53937 1 2809
2 53938 1 2809
2 53939 1 2809
2 53940 1 2809
2 53941 1 2809
2 53942 1 2809
2 53943 1 2809
2 53944 1 2809
2 53945 1 2809
2 53946 1 2809
2 53947 1 2809
2 53948 1 2809
2 53949 1 2809
2 53950 1 2809
2 53951 1 2809
2 53952 1 2809
2 53953 1 2809
2 53954 1 2809
2 53955 1 2809
2 53956 1 2809
2 53957 1 2809
2 53958 1 2809
2 53959 1 2809
2 53960 1 2809
2 53961 1 2809
2 53962 1 2809
2 53963 1 2809
2 53964 1 2809
2 53965 1 2809
2 53966 1 2809
2 53967 1 2809
2 53968 1 2809
2 53969 1 2809
2 53970 1 2809
2 53971 1 2809
2 53972 1 2809
2 53973 1 2809
2 53974 1 2809
2 53975 1 2809
2 53976 1 2809
2 53977 1 2809
2 53978 1 2809
2 53979 1 2809
2 53980 1 2809
2 53981 1 2809
2 53982 1 2809
2 53983 1 2809
2 53984 1 2809
2 53985 1 2809
2 53986 1 2809
2 53987 1 2809
2 53988 1 2809
2 53989 1 2809
2 53990 1 2809
2 53991 1 2809
2 53992 1 2809
2 53993 1 2809
2 53994 1 2809
2 53995 1 2809
2 53996 1 2809
2 53997 1 2809
2 53998 1 2809
2 53999 1 2809
2 54000 1 2809
2 54001 1 2809
2 54002 1 2809
2 54003 1 2809
2 54004 1 2809
2 54005 1 2809
2 54006 1 2809
2 54007 1 2809
2 54008 1 2809
2 54009 1 2809
2 54010 1 2809
2 54011 1 2809
2 54012 1 2809
2 54013 1 2809
2 54014 1 2809
2 54015 1 2809
2 54016 1 2809
2 54017 1 2809
2 54018 1 2809
2 54019 1 2809
2 54020 1 2809
2 54021 1 2809
2 54022 1 2809
2 54023 1 2810
2 54024 1 2810
2 54025 1 2810
2 54026 1 2810
2 54027 1 2810
2 54028 1 2810
2 54029 1 2810
2 54030 1 2810
2 54031 1 2815
2 54032 1 2815
2 54033 1 2823
2 54034 1 2823
2 54035 1 2823
2 54036 1 2823
2 54037 1 2823
2 54038 1 2823
2 54039 1 2823
2 54040 1 2823
2 54041 1 2823
2 54042 1 2823
2 54043 1 2823
2 54044 1 2823
2 54045 1 2823
2 54046 1 2823
2 54047 1 2824
2 54048 1 2824
2 54049 1 2824
2 54050 1 2824
2 54051 1 2837
2 54052 1 2837
2 54053 1 2837
2 54054 1 2838
2 54055 1 2838
2 54056 1 2838
2 54057 1 2838
2 54058 1 2838
2 54059 1 2838
2 54060 1 2838
2 54061 1 2843
2 54062 1 2843
2 54063 1 2843
2 54064 1 2843
2 54065 1 2849
2 54066 1 2849
2 54067 1 2849
2 54068 1 2849
2 54069 1 2849
2 54070 1 2849
2 54071 1 2849
2 54072 1 2849
2 54073 1 2849
2 54074 1 2849
2 54075 1 2849
2 54076 1 2849
2 54077 1 2849
2 54078 1 2849
2 54079 1 2849
2 54080 1 2849
2 54081 1 2849
2 54082 1 2850
2 54083 1 2850
2 54084 1 2850
2 54085 1 2850
2 54086 1 2850
2 54087 1 2850
2 54088 1 2850
2 54089 1 2850
2 54090 1 2850
2 54091 1 2850
2 54092 1 2850
2 54093 1 2850
2 54094 1 2850
2 54095 1 2850
2 54096 1 2850
2 54097 1 2850
2 54098 1 2850
2 54099 1 2850
2 54100 1 2850
2 54101 1 2850
2 54102 1 2850
2 54103 1 2850
2 54104 1 2850
2 54105 1 2850
2 54106 1 2850
2 54107 1 2850
2 54108 1 2850
2 54109 1 2853
2 54110 1 2853
2 54111 1 2853
2 54112 1 2853
2 54113 1 2853
2 54114 1 2854
2 54115 1 2854
2 54116 1 2854
2 54117 1 2854
2 54118 1 2854
2 54119 1 2854
2 54120 1 2854
2 54121 1 2854
2 54122 1 2854
2 54123 1 2854
2 54124 1 2854
2 54125 1 2854
2 54126 1 2854
2 54127 1 2854
2 54128 1 2855
2 54129 1 2855
2 54130 1 2865
2 54131 1 2865
2 54132 1 2865
2 54133 1 2865
2 54134 1 2865
2 54135 1 2865
2 54136 1 2865
2 54137 1 2865
2 54138 1 2865
2 54139 1 2865
2 54140 1 2865
2 54141 1 2865
2 54142 1 2865
2 54143 1 2865
2 54144 1 2865
2 54145 1 2865
2 54146 1 2865
2 54147 1 2865
2 54148 1 2865
2 54149 1 2865
2 54150 1 2865
2 54151 1 2865
2 54152 1 2865
2 54153 1 2865
2 54154 1 2865
2 54155 1 2865
2 54156 1 2865
2 54157 1 2865
2 54158 1 2865
2 54159 1 2865
2 54160 1 2865
2 54161 1 2865
2 54162 1 2865
2 54163 1 2865
2 54164 1 2865
2 54165 1 2865
2 54166 1 2865
2 54167 1 2865
2 54168 1 2865
2 54169 1 2865
2 54170 1 2865
2 54171 1 2865
2 54172 1 2865
2 54173 1 2865
2 54174 1 2865
2 54175 1 2865
2 54176 1 2865
2 54177 1 2865
2 54178 1 2865
2 54179 1 2865
2 54180 1 2865
2 54181 1 2865
2 54182 1 2865
2 54183 1 2865
2 54184 1 2865
2 54185 1 2865
2 54186 1 2865
2 54187 1 2865
2 54188 1 2865
2 54189 1 2865
2 54190 1 2865
2 54191 1 2865
2 54192 1 2865
2 54193 1 2865
2 54194 1 2865
2 54195 1 2865
2 54196 1 2865
2 54197 1 2865
2 54198 1 2865
2 54199 1 2865
2 54200 1 2865
2 54201 1 2865
2 54202 1 2865
2 54203 1 2865
2 54204 1 2865
2 54205 1 2865
2 54206 1 2865
2 54207 1 2867
2 54208 1 2867
2 54209 1 2870
2 54210 1 2870
2 54211 1 2870
2 54212 1 2870
2 54213 1 2870
2 54214 1 2877
2 54215 1 2877
2 54216 1 2877
2 54217 1 2877
2 54218 1 2877
2 54219 1 2878
2 54220 1 2878
2 54221 1 2878
2 54222 1 2878
2 54223 1 2878
2 54224 1 2879
2 54225 1 2879
2 54226 1 2885
2 54227 1 2885
2 54228 1 2886
2 54229 1 2886
2 54230 1 2886
2 54231 1 2886
2 54232 1 2886
2 54233 1 2893
2 54234 1 2893
2 54235 1 2896
2 54236 1 2896
2 54237 1 2896
2 54238 1 2900
2 54239 1 2900
2 54240 1 2900
2 54241 1 2900
2 54242 1 2900
2 54243 1 2901
2 54244 1 2901
2 54245 1 2901
2 54246 1 2906
2 54247 1 2906
2 54248 1 2906
2 54249 1 2911
2 54250 1 2911
2 54251 1 2912
2 54252 1 2912
2 54253 1 2912
2 54254 1 2912
2 54255 1 2912
2 54256 1 2912
2 54257 1 2912
2 54258 1 2913
2 54259 1 2913
2 54260 1 2913
2 54261 1 2913
2 54262 1 2928
2 54263 1 2928
2 54264 1 2928
2 54265 1 2928
2 54266 1 2928
2 54267 1 2928
2 54268 1 2928
2 54269 1 2928
2 54270 1 2928
2 54271 1 2928
2 54272 1 2928
2 54273 1 2928
2 54274 1 2928
2 54275 1 2928
2 54276 1 2928
2 54277 1 2928
2 54278 1 2928
2 54279 1 2928
2 54280 1 2928
2 54281 1 2928
2 54282 1 2928
2 54283 1 2928
2 54284 1 2928
2 54285 1 2928
2 54286 1 2928
2 54287 1 2929
2 54288 1 2929
2 54289 1 2930
2 54290 1 2930
2 54291 1 2930
2 54292 1 2930
2 54293 1 2930
2 54294 1 2930
2 54295 1 2930
2 54296 1 2931
2 54297 1 2931
2 54298 1 2931
2 54299 1 2934
2 54300 1 2934
2 54301 1 2934
2 54302 1 2934
2 54303 1 2935
2 54304 1 2935
2 54305 1 2935
2 54306 1 2942
2 54307 1 2942
2 54308 1 2942
2 54309 1 2942
2 54310 1 2942
2 54311 1 2942
2 54312 1 2942
2 54313 1 2942
2 54314 1 2942
2 54315 1 2942
2 54316 1 2942
2 54317 1 2942
2 54318 1 2942
2 54319 1 2942
2 54320 1 2942
2 54321 1 2942
2 54322 1 2942
2 54323 1 2942
2 54324 1 2942
2 54325 1 2942
2 54326 1 2942
2 54327 1 2942
2 54328 1 2943
2 54329 1 2943
2 54330 1 2943
2 54331 1 2943
2 54332 1 2943
2 54333 1 2943
2 54334 1 2943
2 54335 1 2943
2 54336 1 2944
2 54337 1 2944
2 54338 1 2945
2 54339 1 2945
2 54340 1 2945
2 54341 1 2945
2 54342 1 2945
2 54343 1 2945
2 54344 1 2945
2 54345 1 2945
2 54346 1 2945
2 54347 1 2945
2 54348 1 2945
2 54349 1 2945
2 54350 1 2945
2 54351 1 2945
2 54352 1 2945
2 54353 1 2945
2 54354 1 2945
2 54355 1 2945
2 54356 1 2945
2 54357 1 2945
2 54358 1 2945
2 54359 1 2945
2 54360 1 2945
2 54361 1 2945
2 54362 1 2945
2 54363 1 2945
2 54364 1 2945
2 54365 1 2945
2 54366 1 2945
2 54367 1 2945
2 54368 1 2945
2 54369 1 2945
2 54370 1 2945
2 54371 1 2945
2 54372 1 2945
2 54373 1 2945
2 54374 1 2945
2 54375 1 2945
2 54376 1 2946
2 54377 1 2946
2 54378 1 2954
2 54379 1 2954
2 54380 1 2954
2 54381 1 2954
2 54382 1 2954
2 54383 1 2954
2 54384 1 2954
2 54385 1 2954
2 54386 1 2954
2 54387 1 2954
2 54388 1 2954
2 54389 1 2954
2 54390 1 2954
2 54391 1 2954
2 54392 1 2954
2 54393 1 2954
2 54394 1 2954
2 54395 1 2954
2 54396 1 2957
2 54397 1 2957
2 54398 1 2957
2 54399 1 2957
2 54400 1 2957
2 54401 1 2957
2 54402 1 2957
2 54403 1 2957
2 54404 1 2957
2 54405 1 2957
2 54406 1 2957
2 54407 1 2957
2 54408 1 2957
2 54409 1 2957
2 54410 1 2957
2 54411 1 2957
2 54412 1 2957
2 54413 1 2957
2 54414 1 2957
2 54415 1 2957
2 54416 1 2957
2 54417 1 2957
2 54418 1 2957
2 54419 1 2958
2 54420 1 2958
2 54421 1 2962
2 54422 1 2962
2 54423 1 2962
2 54424 1 2962
2 54425 1 2962
2 54426 1 2962
2 54427 1 2962
2 54428 1 2962
2 54429 1 2962
2 54430 1 2962
2 54431 1 2962
2 54432 1 2962
2 54433 1 2962
2 54434 1 2962
2 54435 1 2962
2 54436 1 2962
2 54437 1 2963
2 54438 1 2963
2 54439 1 2963
2 54440 1 2963
2 54441 1 2963
2 54442 1 2963
2 54443 1 2963
2 54444 1 2963
2 54445 1 2963
2 54446 1 2963
2 54447 1 2963
2 54448 1 2963
2 54449 1 2963
2 54450 1 2963
2 54451 1 2963
2 54452 1 2963
2 54453 1 2964
2 54454 1 2964
2 54455 1 2964
2 54456 1 2964
2 54457 1 2964
2 54458 1 2964
2 54459 1 2964
2 54460 1 2964
2 54461 1 2972
2 54462 1 2972
2 54463 1 2972
2 54464 1 2973
2 54465 1 2973
2 54466 1 2973
2 54467 1 2984
2 54468 1 2984
2 54469 1 2984
2 54470 1 2984
2 54471 1 2984
2 54472 1 2984
2 54473 1 2984
2 54474 1 2984
2 54475 1 2984
2 54476 1 2984
2 54477 1 2984
2 54478 1 2991
2 54479 1 2991
2 54480 1 2991
2 54481 1 2991
2 54482 1 2991
2 54483 1 2997
2 54484 1 2997
2 54485 1 3010
2 54486 1 3010
2 54487 1 3010
2 54488 1 3010
2 54489 1 3010
2 54490 1 3010
2 54491 1 3010
2 54492 1 3010
2 54493 1 3010
2 54494 1 3010
2 54495 1 3010
2 54496 1 3010
2 54497 1 3010
2 54498 1 3010
2 54499 1 3010
2 54500 1 3010
2 54501 1 3010
2 54502 1 3010
2 54503 1 3010
2 54504 1 3010
2 54505 1 3010
2 54506 1 3010
2 54507 1 3010
2 54508 1 3011
2 54509 1 3011
2 54510 1 3011
2 54511 1 3011
2 54512 1 3011
2 54513 1 3012
2 54514 1 3012
2 54515 1 3012
2 54516 1 3013
2 54517 1 3013
2 54518 1 3013
2 54519 1 3021
2 54520 1 3021
2 54521 1 3021
2 54522 1 3021
2 54523 1 3038
2 54524 1 3038
2 54525 1 3049
2 54526 1 3049
2 54527 1 3049
2 54528 1 3049
2 54529 1 3049
2 54530 1 3049
2 54531 1 3049
2 54532 1 3049
2 54533 1 3049
2 54534 1 3049
2 54535 1 3049
2 54536 1 3049
2 54537 1 3050
2 54538 1 3050
2 54539 1 3050
2 54540 1 3050
2 54541 1 3050
2 54542 1 3050
2 54543 1 3050
2 54544 1 3058
2 54545 1 3058
2 54546 1 3058
2 54547 1 3058
2 54548 1 3058
2 54549 1 3058
2 54550 1 3058
2 54551 1 3058
2 54552 1 3058
2 54553 1 3058
2 54554 1 3058
2 54555 1 3059
2 54556 1 3059
2 54557 1 3060
2 54558 1 3060
2 54559 1 3061
2 54560 1 3061
2 54561 1 3061
2 54562 1 3061
2 54563 1 3061
2 54564 1 3062
2 54565 1 3062
2 54566 1 3062
2 54567 1 3062
2 54568 1 3062
2 54569 1 3062
2 54570 1 3062
2 54571 1 3062
2 54572 1 3063
2 54573 1 3063
2 54574 1 3063
2 54575 1 3063
2 54576 1 3063
2 54577 1 3071
2 54578 1 3071
2 54579 1 3071
2 54580 1 3071
2 54581 1 3071
2 54582 1 3071
2 54583 1 3071
2 54584 1 3071
2 54585 1 3071
2 54586 1 3071
2 54587 1 3071
2 54588 1 3075
2 54589 1 3075
2 54590 1 3075
2 54591 1 3075
2 54592 1 3075
2 54593 1 3075
2 54594 1 3075
2 54595 1 3075
2 54596 1 3075
2 54597 1 3075
2 54598 1 3075
2 54599 1 3075
2 54600 1 3075
2 54601 1 3075
2 54602 1 3075
2 54603 1 3075
2 54604 1 3075
2 54605 1 3075
2 54606 1 3075
2 54607 1 3075
2 54608 1 3075
2 54609 1 3075
2 54610 1 3075
2 54611 1 3075
2 54612 1 3075
2 54613 1 3075
2 54614 1 3075
2 54615 1 3075
2 54616 1 3075
2 54617 1 3075
2 54618 1 3075
2 54619 1 3075
2 54620 1 3075
2 54621 1 3075
2 54622 1 3075
2 54623 1 3075
2 54624 1 3075
2 54625 1 3075
2 54626 1 3075
2 54627 1 3075
2 54628 1 3075
2 54629 1 3077
2 54630 1 3077
2 54631 1 3077
2 54632 1 3077
2 54633 1 3077
2 54634 1 3085
2 54635 1 3085
2 54636 1 3085
2 54637 1 3085
2 54638 1 3085
2 54639 1 3086
2 54640 1 3086
2 54641 1 3089
2 54642 1 3089
2 54643 1 3089
2 54644 1 3089
2 54645 1 3096
2 54646 1 3096
2 54647 1 3096
2 54648 1 3096
2 54649 1 3096
2 54650 1 3096
2 54651 1 3096
2 54652 1 3096
2 54653 1 3096
2 54654 1 3096
2 54655 1 3096
2 54656 1 3096
2 54657 1 3096
2 54658 1 3096
2 54659 1 3096
2 54660 1 3098
2 54661 1 3098
2 54662 1 3098
2 54663 1 3111
2 54664 1 3111
2 54665 1 3111
2 54666 1 3111
2 54667 1 3111
2 54668 1 3111
2 54669 1 3111
2 54670 1 3111
2 54671 1 3111
2 54672 1 3112
2 54673 1 3112
2 54674 1 3112
2 54675 1 3112
2 54676 1 3121
2 54677 1 3121
2 54678 1 3121
2 54679 1 3121
2 54680 1 3121
2 54681 1 3121
2 54682 1 3121
2 54683 1 3121
2 54684 1 3121
2 54685 1 3121
2 54686 1 3121
2 54687 1 3121
2 54688 1 3121
2 54689 1 3121
2 54690 1 3122
2 54691 1 3122
2 54692 1 3123
2 54693 1 3123
2 54694 1 3124
2 54695 1 3124
2 54696 1 3124
2 54697 1 3133
2 54698 1 3133
2 54699 1 3133
2 54700 1 3133
2 54701 1 3133
2 54702 1 3133
2 54703 1 3133
2 54704 1 3133
2 54705 1 3133
2 54706 1 3133
2 54707 1 3133
2 54708 1 3141
2 54709 1 3141
2 54710 1 3142
2 54711 1 3142
2 54712 1 3142
2 54713 1 3142
2 54714 1 3144
2 54715 1 3144
2 54716 1 3151
2 54717 1 3151
2 54718 1 3151
2 54719 1 3151
2 54720 1 3151
2 54721 1 3152
2 54722 1 3152
2 54723 1 3161
2 54724 1 3161
2 54725 1 3161
2 54726 1 3161
2 54727 1 3161
2 54728 1 3161
2 54729 1 3161
2 54730 1 3163
2 54731 1 3163
2 54732 1 3163
2 54733 1 3163
2 54734 1 3164
2 54735 1 3164
2 54736 1 3172
2 54737 1 3172
2 54738 1 3173
2 54739 1 3173
2 54740 1 3178
2 54741 1 3178
2 54742 1 3178
2 54743 1 3197
2 54744 1 3197
2 54745 1 3198
2 54746 1 3198
2 54747 1 3199
2 54748 1 3199
2 54749 1 3199
2 54750 1 3199
2 54751 1 3199
2 54752 1 3199
2 54753 1 3199
2 54754 1 3199
2 54755 1 3199
2 54756 1 3199
2 54757 1 3199
2 54758 1 3199
2 54759 1 3200
2 54760 1 3200
2 54761 1 3200
2 54762 1 3200
2 54763 1 3200
2 54764 1 3201
2 54765 1 3201
2 54766 1 3202
2 54767 1 3202
2 54768 1 3203
2 54769 1 3203
2 54770 1 3210
2 54771 1 3210
2 54772 1 3210
2 54773 1 3218
2 54774 1 3218
2 54775 1 3218
2 54776 1 3218
2 54777 1 3218
2 54778 1 3218
2 54779 1 3218
2 54780 1 3218
2 54781 1 3218
2 54782 1 3218
2 54783 1 3218
2 54784 1 3218
2 54785 1 3219
2 54786 1 3219
2 54787 1 3219
2 54788 1 3219
2 54789 1 3219
2 54790 1 3219
2 54791 1 3220
2 54792 1 3220
2 54793 1 3220
2 54794 1 3220
2 54795 1 3220
2 54796 1 3220
2 54797 1 3221
2 54798 1 3221
2 54799 1 3222
2 54800 1 3222
2 54801 1 3222
2 54802 1 3222
2 54803 1 3222
2 54804 1 3222
2 54805 1 3222
2 54806 1 3222
2 54807 1 3222
2 54808 1 3223
2 54809 1 3223
2 54810 1 3223
2 54811 1 3224
2 54812 1 3224
2 54813 1 3224
2 54814 1 3224
2 54815 1 3224
2 54816 1 3226
2 54817 1 3226
2 54818 1 3231
2 54819 1 3231
2 54820 1 3231
2 54821 1 3231
2 54822 1 3231
2 54823 1 3231
2 54824 1 3231
2 54825 1 3231
2 54826 1 3231
2 54827 1 3231
2 54828 1 3231
2 54829 1 3231
2 54830 1 3231
2 54831 1 3231
2 54832 1 3232
2 54833 1 3232
2 54834 1 3232
2 54835 1 3233
2 54836 1 3233
2 54837 1 3234
2 54838 1 3234
2 54839 1 3234
2 54840 1 3234
2 54841 1 3238
2 54842 1 3238
2 54843 1 3238
2 54844 1 3238
2 54845 1 3238
2 54846 1 3238
2 54847 1 3238
2 54848 1 3238
2 54849 1 3238
2 54850 1 3239
2 54851 1 3239
2 54852 1 3239
2 54853 1 3239
2 54854 1 3240
2 54855 1 3240
2 54856 1 3241
2 54857 1 3241
2 54858 1 3241
2 54859 1 3241
2 54860 1 3241
2 54861 1 3241
2 54862 1 3241
2 54863 1 3241
2 54864 1 3241
2 54865 1 3241
2 54866 1 3242
2 54867 1 3242
2 54868 1 3250
2 54869 1 3250
2 54870 1 3250
2 54871 1 3250
2 54872 1 3250
2 54873 1 3250
2 54874 1 3250
2 54875 1 3250
2 54876 1 3250
2 54877 1 3250
2 54878 1 3251
2 54879 1 3251
2 54880 1 3251
2 54881 1 3251
2 54882 1 3251
2 54883 1 3251
2 54884 1 3252
2 54885 1 3252
2 54886 1 3253
2 54887 1 3253
2 54888 1 3253
2 54889 1 3256
2 54890 1 3256
2 54891 1 3258
2 54892 1 3258
2 54893 1 3258
2 54894 1 3260
2 54895 1 3260
2 54896 1 3261
2 54897 1 3261
2 54898 1 3269
2 54899 1 3269
2 54900 1 3270
2 54901 1 3270
2 54902 1 3270
2 54903 1 3270
2 54904 1 3272
2 54905 1 3272
2 54906 1 3281
2 54907 1 3281
2 54908 1 3281
2 54909 1 3282
2 54910 1 3282
2 54911 1 3282
2 54912 1 3284
2 54913 1 3284
2 54914 1 3284
2 54915 1 3289
2 54916 1 3289
2 54917 1 3289
2 54918 1 3289
2 54919 1 3289
2 54920 1 3289
2 54921 1 3289
2 54922 1 3290
2 54923 1 3290
2 54924 1 3290
2 54925 1 3290
2 54926 1 3292
2 54927 1 3292
2 54928 1 3300
2 54929 1 3300
2 54930 1 3300
2 54931 1 3300
2 54932 1 3300
2 54933 1 3300
2 54934 1 3300
2 54935 1 3300
2 54936 1 3301
2 54937 1 3301
2 54938 1 3302
2 54939 1 3302
2 54940 1 3320
2 54941 1 3320
2 54942 1 3322
2 54943 1 3322
2 54944 1 3322
2 54945 1 3322
2 54946 1 3322
2 54947 1 3322
2 54948 1 3324
2 54949 1 3324
2 54950 1 3324
2 54951 1 3324
2 54952 1 3335
2 54953 1 3335
2 54954 1 3335
2 54955 1 3343
2 54956 1 3343
2 54957 1 3343
2 54958 1 3343
2 54959 1 3344
2 54960 1 3344
2 54961 1 3348
2 54962 1 3348
2 54963 1 3348
2 54964 1 3349
2 54965 1 3349
2 54966 1 3349
2 54967 1 3349
2 54968 1 3350
2 54969 1 3350
2 54970 1 3351
2 54971 1 3351
2 54972 1 3351
2 54973 1 3351
2 54974 1 3351
2 54975 1 3359
2 54976 1 3359
2 54977 1 3359
2 54978 1 3359
2 54979 1 3359
2 54980 1 3359
2 54981 1 3359
2 54982 1 3359
2 54983 1 3359
2 54984 1 3359
2 54985 1 3359
2 54986 1 3359
2 54987 1 3359
2 54988 1 3359
2 54989 1 3359
2 54990 1 3360
2 54991 1 3360
2 54992 1 3360
2 54993 1 3360
2 54994 1 3363
2 54995 1 3363
2 54996 1 3363
2 54997 1 3363
2 54998 1 3363
2 54999 1 3363
2 55000 1 3363
2 55001 1 3363
2 55002 1 3363
2 55003 1 3363
2 55004 1 3364
2 55005 1 3364
2 55006 1 3364
2 55007 1 3365
2 55008 1 3365
2 55009 1 3366
2 55010 1 3366
2 55011 1 3369
2 55012 1 3369
2 55013 1 3391
2 55014 1 3391
2 55015 1 3391
2 55016 1 3393
2 55017 1 3393
2 55018 1 3393
2 55019 1 3393
2 55020 1 3393
2 55021 1 3393
2 55022 1 3393
2 55023 1 3395
2 55024 1 3395
2 55025 1 3395
2 55026 1 3395
2 55027 1 3395
2 55028 1 3396
2 55029 1 3396
2 55030 1 3396
2 55031 1 3396
2 55032 1 3396
2 55033 1 3396
2 55034 1 3396
2 55035 1 3396
2 55036 1 3396
2 55037 1 3396
2 55038 1 3396
2 55039 1 3396
2 55040 1 3396
2 55041 1 3396
2 55042 1 3396
2 55043 1 3396
2 55044 1 3396
2 55045 1 3396
2 55046 1 3396
2 55047 1 3396
2 55048 1 3396
2 55049 1 3396
2 55050 1 3396
2 55051 1 3396
2 55052 1 3396
2 55053 1 3396
2 55054 1 3396
2 55055 1 3396
2 55056 1 3396
2 55057 1 3396
2 55058 1 3396
2 55059 1 3396
2 55060 1 3396
2 55061 1 3396
2 55062 1 3396
2 55063 1 3396
2 55064 1 3396
2 55065 1 3396
2 55066 1 3396
2 55067 1 3396
2 55068 1 3396
2 55069 1 3396
2 55070 1 3396
2 55071 1 3396
2 55072 1 3396
2 55073 1 3396
2 55074 1 3396
2 55075 1 3396
2 55076 1 3396
2 55077 1 3396
2 55078 1 3396
2 55079 1 3396
2 55080 1 3396
2 55081 1 3396
2 55082 1 3396
2 55083 1 3396
2 55084 1 3396
2 55085 1 3396
2 55086 1 3396
2 55087 1 3396
2 55088 1 3396
2 55089 1 3396
2 55090 1 3396
2 55091 1 3396
2 55092 1 3396
2 55093 1 3396
2 55094 1 3396
2 55095 1 3396
2 55096 1 3396
2 55097 1 3396
2 55098 1 3396
2 55099 1 3396
2 55100 1 3396
2 55101 1 3396
2 55102 1 3396
2 55103 1 3396
2 55104 1 3396
2 55105 1 3396
2 55106 1 3396
2 55107 1 3396
2 55108 1 3396
2 55109 1 3396
2 55110 1 3396
2 55111 1 3396
2 55112 1 3396
2 55113 1 3396
2 55114 1 3396
2 55115 1 3396
2 55116 1 3396
2 55117 1 3396
2 55118 1 3396
2 55119 1 3396
2 55120 1 3396
2 55121 1 3396
2 55122 1 3396
2 55123 1 3396
2 55124 1 3396
2 55125 1 3396
2 55126 1 3396
2 55127 1 3396
2 55128 1 3396
2 55129 1 3396
2 55130 1 3396
2 55131 1 3396
2 55132 1 3396
2 55133 1 3396
2 55134 1 3396
2 55135 1 3397
2 55136 1 3397
2 55137 1 3397
2 55138 1 3397
2 55139 1 3397
2 55140 1 3397
2 55141 1 3397
2 55142 1 3397
2 55143 1 3398
2 55144 1 3398
2 55145 1 3399
2 55146 1 3399
2 55147 1 3399
2 55148 1 3399
2 55149 1 3399
2 55150 1 3399
2 55151 1 3399
2 55152 1 3399
2 55153 1 3399
2 55154 1 3400
2 55155 1 3400
2 55156 1 3400
2 55157 1 3400
2 55158 1 3400
2 55159 1 3400
2 55160 1 3400
2 55161 1 3400
2 55162 1 3401
2 55163 1 3401
2 55164 1 3401
2 55165 1 3401
2 55166 1 3403
2 55167 1 3403
2 55168 1 3403
2 55169 1 3403
2 55170 1 3403
2 55171 1 3403
2 55172 1 3403
2 55173 1 3403
2 55174 1 3403
2 55175 1 3403
2 55176 1 3403
2 55177 1 3403
2 55178 1 3404
2 55179 1 3404
2 55180 1 3404
2 55181 1 3404
2 55182 1 3404
2 55183 1 3404
2 55184 1 3404
2 55185 1 3404
2 55186 1 3404
2 55187 1 3407
2 55188 1 3407
2 55189 1 3407
2 55190 1 3407
2 55191 1 3407
2 55192 1 3407
2 55193 1 3407
2 55194 1 3409
2 55195 1 3409
2 55196 1 3409
2 55197 1 3410
2 55198 1 3410
2 55199 1 3410
2 55200 1 3410
2 55201 1 3410
2 55202 1 3410
2 55203 1 3410
2 55204 1 3410
2 55205 1 3411
2 55206 1 3411
2 55207 1 3413
2 55208 1 3413
2 55209 1 3416
2 55210 1 3416
2 55211 1 3416
2 55212 1 3416
2 55213 1 3416
2 55214 1 3416
2 55215 1 3416
2 55216 1 3416
2 55217 1 3424
2 55218 1 3424
2 55219 1 3426
2 55220 1 3426
2 55221 1 3426
2 55222 1 3426
2 55223 1 3426
2 55224 1 3426
2 55225 1 3426
2 55226 1 3426
2 55227 1 3426
2 55228 1 3426
2 55229 1 3426
2 55230 1 3426
2 55231 1 3426
2 55232 1 3426
2 55233 1 3426
2 55234 1 3426
2 55235 1 3426
2 55236 1 3426
2 55237 1 3426
2 55238 1 3426
2 55239 1 3426
2 55240 1 3426
2 55241 1 3426
2 55242 1 3426
2 55243 1 3426
2 55244 1 3426
2 55245 1 3426
2 55246 1 3426
2 55247 1 3426
2 55248 1 3426
2 55249 1 3426
2 55250 1 3426
2 55251 1 3426
2 55252 1 3426
2 55253 1 3426
2 55254 1 3426
2 55255 1 3426
2 55256 1 3426
2 55257 1 3426
2 55258 1 3426
2 55259 1 3426
2 55260 1 3426
2 55261 1 3426
2 55262 1 3426
2 55263 1 3426
2 55264 1 3429
2 55265 1 3429
2 55266 1 3429
2 55267 1 3429
2 55268 1 3431
2 55269 1 3431
2 55270 1 3431
2 55271 1 3438
2 55272 1 3438
2 55273 1 3438
2 55274 1 3438
2 55275 1 3438
2 55276 1 3438
2 55277 1 3438
2 55278 1 3439
2 55279 1 3439
2 55280 1 3439
2 55281 1 3451
2 55282 1 3451
2 55283 1 3451
2 55284 1 3452
2 55285 1 3452
2 55286 1 3453
2 55287 1 3453
2 55288 1 3453
2 55289 1 3453
2 55290 1 3453
2 55291 1 3453
2 55292 1 3453
2 55293 1 3453
2 55294 1 3457
2 55295 1 3457
2 55296 1 3457
2 55297 1 3457
2 55298 1 3457
2 55299 1 3457
2 55300 1 3457
2 55301 1 3457
2 55302 1 3457
2 55303 1 3457
2 55304 1 3457
2 55305 1 3457
2 55306 1 3458
2 55307 1 3458
2 55308 1 3458
2 55309 1 3458
2 55310 1 3460
2 55311 1 3460
2 55312 1 3460
2 55313 1 3460
2 55314 1 3460
2 55315 1 3460
2 55316 1 3460
2 55317 1 3460
2 55318 1 3460
2 55319 1 3460
2 55320 1 3460
2 55321 1 3460
2 55322 1 3461
2 55323 1 3461
2 55324 1 3463
2 55325 1 3463
2 55326 1 3463
2 55327 1 3463
2 55328 1 3463
2 55329 1 3463
2 55330 1 3463
2 55331 1 3463
2 55332 1 3463
2 55333 1 3463
2 55334 1 3463
2 55335 1 3463
2 55336 1 3472
2 55337 1 3472
2 55338 1 3472
2 55339 1 3472
2 55340 1 3472
2 55341 1 3472
2 55342 1 3472
2 55343 1 3472
2 55344 1 3472
2 55345 1 3472
2 55346 1 3472
2 55347 1 3472
2 55348 1 3474
2 55349 1 3474
2 55350 1 3478
2 55351 1 3478
2 55352 1 3478
2 55353 1 3478
2 55354 1 3478
2 55355 1 3478
2 55356 1 3480
2 55357 1 3480
2 55358 1 3480
2 55359 1 3483
2 55360 1 3483
2 55361 1 3484
2 55362 1 3484
2 55363 1 3492
2 55364 1 3492
2 55365 1 3492
2 55366 1 3492
2 55367 1 3492
2 55368 1 3492
2 55369 1 3492
2 55370 1 3492
2 55371 1 3492
2 55372 1 3492
2 55373 1 3492
2 55374 1 3492
2 55375 1 3492
2 55376 1 3492
2 55377 1 3492
2 55378 1 3492
2 55379 1 3492
2 55380 1 3492
2 55381 1 3492
2 55382 1 3492
2 55383 1 3492
2 55384 1 3493
2 55385 1 3493
2 55386 1 3494
2 55387 1 3494
2 55388 1 3494
2 55389 1 3494
2 55390 1 3494
2 55391 1 3494
2 55392 1 3494
2 55393 1 3494
2 55394 1 3495
2 55395 1 3495
2 55396 1 3495
2 55397 1 3496
2 55398 1 3496
2 55399 1 3496
2 55400 1 3496
2 55401 1 3496
2 55402 1 3496
2 55403 1 3516
2 55404 1 3516
2 55405 1 3516
2 55406 1 3516
2 55407 1 3516
2 55408 1 3516
2 55409 1 3516
2 55410 1 3516
2 55411 1 3516
2 55412 1 3516
2 55413 1 3516
2 55414 1 3516
2 55415 1 3517
2 55416 1 3517
2 55417 1 3517
2 55418 1 3517
2 55419 1 3517
2 55420 1 3517
2 55421 1 3517
2 55422 1 3517
2 55423 1 3517
2 55424 1 3517
2 55425 1 3518
2 55426 1 3518
2 55427 1 3518
2 55428 1 3518
2 55429 1 3518
2 55430 1 3518
2 55431 1 3518
2 55432 1 3518
2 55433 1 3518
2 55434 1 3519
2 55435 1 3519
2 55436 1 3519
2 55437 1 3520
2 55438 1 3520
2 55439 1 3520
2 55440 1 3520
2 55441 1 3523
2 55442 1 3523
2 55443 1 3530
2 55444 1 3530
2 55445 1 3531
2 55446 1 3531
2 55447 1 3532
2 55448 1 3532
2 55449 1 3532
2 55450 1 3544
2 55451 1 3544
2 55452 1 3544
2 55453 1 3544
2 55454 1 3544
2 55455 1 3544
2 55456 1 3544
2 55457 1 3544
2 55458 1 3544
2 55459 1 3544
2 55460 1 3544
2 55461 1 3544
2 55462 1 3544
2 55463 1 3544
2 55464 1 3544
2 55465 1 3544
2 55466 1 3550
2 55467 1 3550
2 55468 1 3550
2 55469 1 3550
2 55470 1 3550
2 55471 1 3550
2 55472 1 3550
2 55473 1 3551
2 55474 1 3551
2 55475 1 3552
2 55476 1 3552
2 55477 1 3559
2 55478 1 3559
2 55479 1 3559
2 55480 1 3559
2 55481 1 3559
2 55482 1 3559
2 55483 1 3569
2 55484 1 3569
2 55485 1 3569
2 55486 1 3570
2 55487 1 3570
2 55488 1 3570
2 55489 1 3570
2 55490 1 3570
2 55491 1 3570
2 55492 1 3570
2 55493 1 3570
2 55494 1 3571
2 55495 1 3571
2 55496 1 3571
2 55497 1 3571
2 55498 1 3571
2 55499 1 3571
2 55500 1 3571
2 55501 1 3571
2 55502 1 3571
2 55503 1 3571
2 55504 1 3572
2 55505 1 3572
2 55506 1 3572
2 55507 1 3573
2 55508 1 3573
2 55509 1 3581
2 55510 1 3581
2 55511 1 3581
2 55512 1 3581
2 55513 1 3584
2 55514 1 3584
2 55515 1 3586
2 55516 1 3586
2 55517 1 3586
2 55518 1 3586
2 55519 1 3586
2 55520 1 3586
2 55521 1 3586
2 55522 1 3586
2 55523 1 3586
2 55524 1 3586
2 55525 1 3586
2 55526 1 3586
2 55527 1 3587
2 55528 1 3587
2 55529 1 3590
2 55530 1 3590
2 55531 1 3590
2 55532 1 3591
2 55533 1 3591
2 55534 1 3601
2 55535 1 3601
2 55536 1 3601
2 55537 1 3601
2 55538 1 3601
2 55539 1 3601
2 55540 1 3601
2 55541 1 3601
2 55542 1 3601
2 55543 1 3601
2 55544 1 3601
2 55545 1 3612
2 55546 1 3612
2 55547 1 3613
2 55548 1 3613
2 55549 1 3619
2 55550 1 3619
2 55551 1 3619
2 55552 1 3619
2 55553 1 3619
2 55554 1 3619
2 55555 1 3619
2 55556 1 3629
2 55557 1 3629
2 55558 1 3629
2 55559 1 3631
2 55560 1 3631
2 55561 1 3642
2 55562 1 3642
2 55563 1 3642
2 55564 1 3650
2 55565 1 3650
2 55566 1 3650
2 55567 1 3654
2 55568 1 3654
2 55569 1 3654
2 55570 1 3654
2 55571 1 3654
2 55572 1 3654
2 55573 1 3654
2 55574 1 3663
2 55575 1 3663
2 55576 1 3663
2 55577 1 3663
2 55578 1 3663
2 55579 1 3663
2 55580 1 3663
2 55581 1 3665
2 55582 1 3665
2 55583 1 3672
2 55584 1 3672
2 55585 1 3679
2 55586 1 3679
2 55587 1 3679
2 55588 1 3679
2 55589 1 3679
2 55590 1 3679
2 55591 1 3679
2 55592 1 3695
2 55593 1 3695
2 55594 1 3695
2 55595 1 3695
2 55596 1 3695
2 55597 1 3695
2 55598 1 3695
2 55599 1 3695
2 55600 1 3696
2 55601 1 3696
2 55602 1 3696
2 55603 1 3696
2 55604 1 3696
2 55605 1 3696
2 55606 1 3696
2 55607 1 3696
2 55608 1 3696
2 55609 1 3703
2 55610 1 3703
2 55611 1 3704
2 55612 1 3704
2 55613 1 3704
2 55614 1 3704
2 55615 1 3704
2 55616 1 3704
2 55617 1 3704
2 55618 1 3704
2 55619 1 3707
2 55620 1 3707
2 55621 1 3707
2 55622 1 3707
2 55623 1 3708
2 55624 1 3708
2 55625 1 3719
2 55626 1 3719
2 55627 1 3720
2 55628 1 3720
2 55629 1 3721
2 55630 1 3721
2 55631 1 3722
2 55632 1 3722
2 55633 1 3723
2 55634 1 3723
2 55635 1 3723
2 55636 1 3723
2 55637 1 3724
2 55638 1 3724
2 55639 1 3727
2 55640 1 3727
2 55641 1 3727
2 55642 1 3727
2 55643 1 3727
2 55644 1 3727
2 55645 1 3727
2 55646 1 3736
2 55647 1 3736
2 55648 1 3736
2 55649 1 3739
2 55650 1 3739
2 55651 1 3739
2 55652 1 3739
2 55653 1 3739
2 55654 1 3747
2 55655 1 3747
2 55656 1 3747
2 55657 1 3747
2 55658 1 3749
2 55659 1 3749
2 55660 1 3751
2 55661 1 3751
2 55662 1 3755
2 55663 1 3755
2 55664 1 3765
2 55665 1 3765
2 55666 1 3765
2 55667 1 3765
2 55668 1 3765
2 55669 1 3765
2 55670 1 3765
2 55671 1 3765
2 55672 1 3765
2 55673 1 3765
2 55674 1 3765
2 55675 1 3765
2 55676 1 3765
2 55677 1 3765
2 55678 1 3765
2 55679 1 3765
2 55680 1 3765
2 55681 1 3765
2 55682 1 3766
2 55683 1 3766
2 55684 1 3766
2 55685 1 3766
2 55686 1 3766
2 55687 1 3766
2 55688 1 3766
2 55689 1 3766
2 55690 1 3767
2 55691 1 3767
2 55692 1 3767
2 55693 1 3770
2 55694 1 3770
2 55695 1 3775
2 55696 1 3775
2 55697 1 3775
2 55698 1 3775
2 55699 1 3775
2 55700 1 3777
2 55701 1 3777
2 55702 1 3778
2 55703 1 3778
2 55704 1 3778
2 55705 1 3778
2 55706 1 3780
2 55707 1 3780
2 55708 1 3781
2 55709 1 3781
2 55710 1 3781
2 55711 1 3781
2 55712 1 3781
2 55713 1 3781
2 55714 1 3785
2 55715 1 3785
2 55716 1 3785
2 55717 1 3796
2 55718 1 3796
2 55719 1 3796
2 55720 1 3796
2 55721 1 3796
2 55722 1 3798
2 55723 1 3798
2 55724 1 3798
2 55725 1 3798
2 55726 1 3798
2 55727 1 3799
2 55728 1 3799
2 55729 1 3799
2 55730 1 3799
2 55731 1 3799
2 55732 1 3806
2 55733 1 3806
2 55734 1 3813
2 55735 1 3813
2 55736 1 3813
2 55737 1 3813
2 55738 1 3813
2 55739 1 3813
2 55740 1 3813
2 55741 1 3813
2 55742 1 3813
2 55743 1 3813
2 55744 1 3813
2 55745 1 3814
2 55746 1 3814
2 55747 1 3816
2 55748 1 3816
2 55749 1 3816
2 55750 1 3816
2 55751 1 3816
2 55752 1 3816
2 55753 1 3816
2 55754 1 3816
2 55755 1 3816
2 55756 1 3816
2 55757 1 3816
2 55758 1 3820
2 55759 1 3820
2 55760 1 3828
2 55761 1 3828
2 55762 1 3828
2 55763 1 3828
2 55764 1 3828
2 55765 1 3828
2 55766 1 3828
2 55767 1 3828
2 55768 1 3828
2 55769 1 3829
2 55770 1 3829
2 55771 1 3835
2 55772 1 3835
2 55773 1 3835
2 55774 1 3835
2 55775 1 3835
2 55776 1 3835
2 55777 1 3835
2 55778 1 3835
2 55779 1 3835
2 55780 1 3835
2 55781 1 3836
2 55782 1 3836
2 55783 1 3838
2 55784 1 3838
2 55785 1 3844
2 55786 1 3844
2 55787 1 3844
2 55788 1 3844
2 55789 1 3844
2 55790 1 3845
2 55791 1 3845
2 55792 1 3845
2 55793 1 3845
2 55794 1 3845
2 55795 1 3846
2 55796 1 3846
2 55797 1 3846
2 55798 1 3847
2 55799 1 3847
2 55800 1 3848
2 55801 1 3848
2 55802 1 3850
2 55803 1 3850
2 55804 1 3850
2 55805 1 3850
2 55806 1 3850
2 55807 1 3854
2 55808 1 3854
2 55809 1 3858
2 55810 1 3858
2 55811 1 3858
2 55812 1 3858
2 55813 1 3865
2 55814 1 3865
2 55815 1 3865
2 55816 1 3865
2 55817 1 3865
2 55818 1 3865
2 55819 1 3865
2 55820 1 3865
2 55821 1 3865
2 55822 1 3865
2 55823 1 3865
2 55824 1 3865
2 55825 1 3865
2 55826 1 3877
2 55827 1 3877
2 55828 1 3877
2 55829 1 3877
2 55830 1 3878
2 55831 1 3878
2 55832 1 3878
2 55833 1 3878
2 55834 1 3878
2 55835 1 3879
2 55836 1 3879
2 55837 1 3879
2 55838 1 3880
2 55839 1 3880
2 55840 1 3880
2 55841 1 3880
2 55842 1 3880
2 55843 1 3880
2 55844 1 3881
2 55845 1 3881
2 55846 1 3892
2 55847 1 3892
2 55848 1 3892
2 55849 1 3894
2 55850 1 3894
2 55851 1 3894
2 55852 1 3904
2 55853 1 3904
2 55854 1 3904
2 55855 1 3904
2 55856 1 3904
2 55857 1 3904
2 55858 1 3904
2 55859 1 3904
2 55860 1 3905
2 55861 1 3905
2 55862 1 3908
2 55863 1 3908
2 55864 1 3908
2 55865 1 3908
2 55866 1 3908
2 55867 1 3908
2 55868 1 3909
2 55869 1 3909
2 55870 1 3909
2 55871 1 3911
2 55872 1 3911
2 55873 1 3911
2 55874 1 3911
2 55875 1 3920
2 55876 1 3920
2 55877 1 3921
2 55878 1 3921
2 55879 1 3921
2 55880 1 3922
2 55881 1 3922
2 55882 1 3922
2 55883 1 3950
2 55884 1 3950
2 55885 1 3950
2 55886 1 3950
2 55887 1 3950
2 55888 1 3950
2 55889 1 3950
2 55890 1 3950
2 55891 1 3950
2 55892 1 3950
2 55893 1 3951
2 55894 1 3951
2 55895 1 3951
2 55896 1 3952
2 55897 1 3952
2 55898 1 3953
2 55899 1 3953
2 55900 1 3959
2 55901 1 3959
2 55902 1 3960
2 55903 1 3960
2 55904 1 3960
2 55905 1 3960
2 55906 1 3962
2 55907 1 3962
2 55908 1 3966
2 55909 1 3966
2 55910 1 3969
2 55911 1 3969
2 55912 1 3973
2 55913 1 3973
2 55914 1 3978
2 55915 1 3978
2 55916 1 3990
2 55917 1 3990
2 55918 1 3990
2 55919 1 3990
2 55920 1 3991
2 55921 1 3991
2 55922 1 3992
2 55923 1 3992
2 55924 1 3993
2 55925 1 3993
2 55926 1 3995
2 55927 1 3995
2 55928 1 3995
2 55929 1 3997
2 55930 1 3997
2 55931 1 3997
2 55932 1 4001
2 55933 1 4001
2 55934 1 4006
2 55935 1 4006
2 55936 1 4008
2 55937 1 4008
2 55938 1 4023
2 55939 1 4023
2 55940 1 4023
2 55941 1 4023
2 55942 1 4024
2 55943 1 4024
2 55944 1 4024
2 55945 1 4025
2 55946 1 4025
2 55947 1 4026
2 55948 1 4026
2 55949 1 4026
2 55950 1 4028
2 55951 1 4028
2 55952 1 4054
2 55953 1 4054
2 55954 1 4069
2 55955 1 4069
2 55956 1 4069
2 55957 1 4070
2 55958 1 4070
2 55959 1 4071
2 55960 1 4071
2 55961 1 4078
2 55962 1 4078
2 55963 1 4078
2 55964 1 4078
2 55965 1 4079
2 55966 1 4079
2 55967 1 4100
2 55968 1 4100
2 55969 1 4106
2 55970 1 4106
2 55971 1 4120
2 55972 1 4120
2 55973 1 4120
2 55974 1 4121
2 55975 1 4121
2 55976 1 4125
2 55977 1 4125
2 55978 1 4125
2 55979 1 4137
2 55980 1 4137
2 55981 1 4137
2 55982 1 4138
2 55983 1 4138
2 55984 1 4138
2 55985 1 4138
2 55986 1 4138
2 55987 1 4147
2 55988 1 4147
2 55989 1 4147
2 55990 1 4147
2 55991 1 4147
2 55992 1 4147
2 55993 1 4148
2 55994 1 4148
2 55995 1 4149
2 55996 1 4149
2 55997 1 4152
2 55998 1 4152
2 55999 1 4152
2 56000 1 4152
2 56001 1 4152
2 56002 1 4152
2 56003 1 4152
2 56004 1 4152
2 56005 1 4152
2 56006 1 4161
2 56007 1 4161
2 56008 1 4161
2 56009 1 4161
2 56010 1 4161
2 56011 1 4161
2 56012 1 4161
2 56013 1 4161
2 56014 1 4161
2 56015 1 4161
2 56016 1 4161
2 56017 1 4163
2 56018 1 4163
2 56019 1 4187
2 56020 1 4187
2 56021 1 4187
2 56022 1 4188
2 56023 1 4188
2 56024 1 4201
2 56025 1 4201
2 56026 1 4201
2 56027 1 4201
2 56028 1 4201
2 56029 1 4201
2 56030 1 4201
2 56031 1 4201
2 56032 1 4201
2 56033 1 4201
2 56034 1 4201
2 56035 1 4213
2 56036 1 4213
2 56037 1 4213
2 56038 1 4213
2 56039 1 4213
2 56040 1 4213
2 56041 1 4214
2 56042 1 4214
2 56043 1 4214
2 56044 1 4214
2 56045 1 4214
2 56046 1 4215
2 56047 1 4215
2 56048 1 4215
2 56049 1 4215
2 56050 1 4215
2 56051 1 4215
2 56052 1 4222
2 56053 1 4222
2 56054 1 4222
2 56055 1 4222
2 56056 1 4223
2 56057 1 4223
2 56058 1 4231
2 56059 1 4231
2 56060 1 4231
2 56061 1 4231
2 56062 1 4231
2 56063 1 4231
2 56064 1 4232
2 56065 1 4232
2 56066 1 4232
2 56067 1 4232
2 56068 1 4232
2 56069 1 4232
2 56070 1 4232
2 56071 1 4232
2 56072 1 4232
2 56073 1 4232
2 56074 1 4232
2 56075 1 4232
2 56076 1 4232
2 56077 1 4232
2 56078 1 4232
2 56079 1 4232
2 56080 1 4232
2 56081 1 4233
2 56082 1 4233
2 56083 1 4233
2 56084 1 4233
2 56085 1 4235
2 56086 1 4235
2 56087 1 4242
2 56088 1 4242
2 56089 1 4242
2 56090 1 4242
2 56091 1 4242
2 56092 1 4242
2 56093 1 4242
2 56094 1 4242
2 56095 1 4242
2 56096 1 4242
2 56097 1 4242
2 56098 1 4243
2 56099 1 4243
2 56100 1 4243
2 56101 1 4243
2 56102 1 4248
2 56103 1 4248
2 56104 1 4252
2 56105 1 4252
2 56106 1 4253
2 56107 1 4253
2 56108 1 4254
2 56109 1 4254
2 56110 1 4255
2 56111 1 4255
2 56112 1 4262
2 56113 1 4262
2 56114 1 4264
2 56115 1 4264
2 56116 1 4264
2 56117 1 4264
2 56118 1 4264
2 56119 1 4264
2 56120 1 4264
2 56121 1 4264
2 56122 1 4305
2 56123 1 4305
2 56124 1 4305
2 56125 1 4312
2 56126 1 4312
2 56127 1 4312
2 56128 1 4312
2 56129 1 4312
2 56130 1 4313
2 56131 1 4313
2 56132 1 4322
2 56133 1 4322
2 56134 1 4322
2 56135 1 4322
2 56136 1 4323
2 56137 1 4323
2 56138 1 4323
2 56139 1 4323
2 56140 1 4323
2 56141 1 4323
2 56142 1 4324
2 56143 1 4324
2 56144 1 4325
2 56145 1 4325
2 56146 1 4328
2 56147 1 4328
2 56148 1 4328
2 56149 1 4328
2 56150 1 4328
2 56151 1 4328
2 56152 1 4328
2 56153 1 4328
2 56154 1 4329
2 56155 1 4329
2 56156 1 4331
2 56157 1 4331
2 56158 1 4334
2 56159 1 4334
2 56160 1 4334
2 56161 1 4334
2 56162 1 4335
2 56163 1 4335
2 56164 1 4342
2 56165 1 4342
2 56166 1 4342
2 56167 1 4342
2 56168 1 4342
2 56169 1 4342
2 56170 1 4342
2 56171 1 4354
2 56172 1 4354
2 56173 1 4368
2 56174 1 4368
2 56175 1 4368
2 56176 1 4368
2 56177 1 4368
2 56178 1 4368
2 56179 1 4368
2 56180 1 4368
2 56181 1 4368
2 56182 1 4368
2 56183 1 4368
2 56184 1 4368
2 56185 1 4368
2 56186 1 4369
2 56187 1 4369
2 56188 1 4369
2 56189 1 4369
2 56190 1 4370
2 56191 1 4370
2 56192 1 4370
2 56193 1 4408
2 56194 1 4408
2 56195 1 4408
2 56196 1 4408
2 56197 1 4408
2 56198 1 4408
2 56199 1 4409
2 56200 1 4409
2 56201 1 4409
2 56202 1 4409
2 56203 1 4409
2 56204 1 4409
2 56205 1 4409
2 56206 1 4409
2 56207 1 4409
2 56208 1 4409
2 56209 1 4409
2 56210 1 4409
2 56211 1 4416
2 56212 1 4416
2 56213 1 4416
2 56214 1 4416
2 56215 1 4448
2 56216 1 4448
2 56217 1 4459
2 56218 1 4459
2 56219 1 4459
2 56220 1 4459
2 56221 1 4459
2 56222 1 4459
2 56223 1 4459
2 56224 1 4492
2 56225 1 4492
2 56226 1 4492
2 56227 1 4492
2 56228 1 4492
2 56229 1 4495
2 56230 1 4495
2 56231 1 4495
2 56232 1 4495
2 56233 1 4511
2 56234 1 4511
2 56235 1 4511
2 56236 1 4511
2 56237 1 4511
2 56238 1 4511
2 56239 1 4512
2 56240 1 4512
2 56241 1 4512
2 56242 1 4514
2 56243 1 4514
2 56244 1 4514
2 56245 1 4518
2 56246 1 4518
2 56247 1 4527
2 56248 1 4527
2 56249 1 4527
2 56250 1 4528
2 56251 1 4528
2 56252 1 4532
2 56253 1 4532
2 56254 1 4532
2 56255 1 4532
2 56256 1 4532
2 56257 1 4532
2 56258 1 4532
2 56259 1 4532
2 56260 1 4532
2 56261 1 4532
2 56262 1 4532
2 56263 1 4532
2 56264 1 4532
2 56265 1 4533
2 56266 1 4533
2 56267 1 4534
2 56268 1 4534
2 56269 1 4534
2 56270 1 4534
2 56271 1 4534
2 56272 1 4547
2 56273 1 4547
2 56274 1 4548
2 56275 1 4548
2 56276 1 4548
2 56277 1 4549
2 56278 1 4549
2 56279 1 4549
2 56280 1 4549
2 56281 1 4549
2 56282 1 4549
2 56283 1 4549
2 56284 1 4549
2 56285 1 4549
2 56286 1 4549
2 56287 1 4549
2 56288 1 4549
2 56289 1 4549
2 56290 1 4549
2 56291 1 4549
2 56292 1 4549
2 56293 1 4549
2 56294 1 4549
2 56295 1 4549
2 56296 1 4549
2 56297 1 4553
2 56298 1 4553
2 56299 1 4554
2 56300 1 4554
2 56301 1 4555
2 56302 1 4555
2 56303 1 4561
2 56304 1 4561
2 56305 1 4561
2 56306 1 4561
2 56307 1 4562
2 56308 1 4562
2 56309 1 4585
2 56310 1 4585
2 56311 1 4585
2 56312 1 4585
2 56313 1 4590
2 56314 1 4590
2 56315 1 4600
2 56316 1 4600
2 56317 1 4603
2 56318 1 4603
2 56319 1 4604
2 56320 1 4604
2 56321 1 4605
2 56322 1 4605
2 56323 1 4605
2 56324 1 4609
2 56325 1 4609
2 56326 1 4609
2 56327 1 4613
2 56328 1 4613
2 56329 1 4613
2 56330 1 4613
2 56331 1 4613
2 56332 1 4613
2 56333 1 4613
2 56334 1 4622
2 56335 1 4622
2 56336 1 4622
2 56337 1 4622
2 56338 1 4622
2 56339 1 4622
2 56340 1 4623
2 56341 1 4623
2 56342 1 4623
2 56343 1 4626
2 56344 1 4626
2 56345 1 4626
2 56346 1 4626
2 56347 1 4626
2 56348 1 4626
2 56349 1 4626
2 56350 1 4626
2 56351 1 4626
2 56352 1 4626
2 56353 1 4626
2 56354 1 4626
2 56355 1 4626
2 56356 1 4626
2 56357 1 4626
2 56358 1 4626
2 56359 1 4631
2 56360 1 4631
2 56361 1 4631
2 56362 1 4631
2 56363 1 4636
2 56364 1 4636
2 56365 1 4644
2 56366 1 4644
2 56367 1 4646
2 56368 1 4646
2 56369 1 4646
2 56370 1 4646
2 56371 1 4646
2 56372 1 4658
2 56373 1 4658
2 56374 1 4658
2 56375 1 4668
2 56376 1 4668
2 56377 1 4676
2 56378 1 4676
2 56379 1 4676
2 56380 1 4676
2 56381 1 4676
2 56382 1 4676
2 56383 1 4676
2 56384 1 4676
2 56385 1 4676
2 56386 1 4677
2 56387 1 4677
2 56388 1 4686
2 56389 1 4686
2 56390 1 4686
2 56391 1 4686
2 56392 1 4686
2 56393 1 4687
2 56394 1 4687
2 56395 1 4687
2 56396 1 4688
2 56397 1 4688
2 56398 1 4699
2 56399 1 4699
2 56400 1 4700
2 56401 1 4700
2 56402 1 4700
2 56403 1 4700
2 56404 1 4700
2 56405 1 4700
2 56406 1 4701
2 56407 1 4701
2 56408 1 4701
2 56409 1 4710
2 56410 1 4710
2 56411 1 4717
2 56412 1 4717
2 56413 1 4717
2 56414 1 4717
2 56415 1 4718
2 56416 1 4718
2 56417 1 4722
2 56418 1 4722
2 56419 1 4729
2 56420 1 4729
2 56421 1 4736
2 56422 1 4736
2 56423 1 4765
2 56424 1 4765
2 56425 1 4765
2 56426 1 4765
2 56427 1 4772
2 56428 1 4772
2 56429 1 4780
2 56430 1 4780
2 56431 1 4780
2 56432 1 4780
2 56433 1 4780
2 56434 1 4780
2 56435 1 4800
2 56436 1 4800
2 56437 1 4800
2 56438 1 4800
2 56439 1 4813
2 56440 1 4813
2 56441 1 4813
2 56442 1 4813
2 56443 1 4813
2 56444 1 4813
2 56445 1 4813
2 56446 1 4813
2 56447 1 4814
2 56448 1 4814
2 56449 1 4814
2 56450 1 4814
2 56451 1 4814
2 56452 1 4815
2 56453 1 4815
2 56454 1 4820
2 56455 1 4820
2 56456 1 4820
2 56457 1 4820
2 56458 1 4820
2 56459 1 4822
2 56460 1 4822
2 56461 1 4822
2 56462 1 4826
2 56463 1 4826
2 56464 1 4837
2 56465 1 4837
2 56466 1 4837
2 56467 1 4837
2 56468 1 4838
2 56469 1 4838
2 56470 1 4839
2 56471 1 4839
2 56472 1 4849
2 56473 1 4849
2 56474 1 4849
2 56475 1 4858
2 56476 1 4858
2 56477 1 4858
2 56478 1 4858
2 56479 1 4858
2 56480 1 4880
2 56481 1 4880
2 56482 1 4880
2 56483 1 4880
2 56484 1 4880
2 56485 1 4881
2 56486 1 4881
2 56487 1 4881
2 56488 1 4881
2 56489 1 4881
2 56490 1 4886
2 56491 1 4886
2 56492 1 4886
2 56493 1 4886
2 56494 1 4887
2 56495 1 4887
2 56496 1 4895
2 56497 1 4895
2 56498 1 4895
2 56499 1 4895
2 56500 1 4895
2 56501 1 4903
2 56502 1 4903
2 56503 1 4903
2 56504 1 4943
2 56505 1 4943
2 56506 1 4943
2 56507 1 4943
2 56508 1 4943
2 56509 1 4943
2 56510 1 4943
2 56511 1 4944
2 56512 1 4944
2 56513 1 4945
2 56514 1 4945
2 56515 1 4947
2 56516 1 4947
2 56517 1 4950
2 56518 1 4950
2 56519 1 4950
2 56520 1 4950
2 56521 1 4963
2 56522 1 4963
2 56523 1 4963
2 56524 1 4963
2 56525 1 4963
2 56526 1 4963
2 56527 1 4965
2 56528 1 4965
2 56529 1 4965
2 56530 1 4965
2 56531 1 4972
2 56532 1 4972
2 56533 1 4972
2 56534 1 4973
2 56535 1 4973
2 56536 1 4980
2 56537 1 4980
2 56538 1 4988
2 56539 1 4988
2 56540 1 4988
2 56541 1 4988
2 56542 1 4988
2 56543 1 4988
2 56544 1 4988
2 56545 1 4988
2 56546 1 4988
2 56547 1 4988
2 56548 1 4988
2 56549 1 4989
2 56550 1 4989
2 56551 1 4989
2 56552 1 4989
2 56553 1 4990
2 56554 1 4990
2 56555 1 4991
2 56556 1 4991
2 56557 1 4991
2 56558 1 4991
2 56559 1 4991
2 56560 1 4991
2 56561 1 4992
2 56562 1 4992
2 56563 1 4992
2 56564 1 4992
2 56565 1 4992
2 56566 1 4992
2 56567 1 4992
2 56568 1 4992
2 56569 1 4992
2 56570 1 5001
2 56571 1 5001
2 56572 1 5001
2 56573 1 5001
2 56574 1 5001
2 56575 1 5002
2 56576 1 5002
2 56577 1 5002
2 56578 1 5003
2 56579 1 5003
2 56580 1 5003
2 56581 1 5003
2 56582 1 5003
2 56583 1 5003
2 56584 1 5003
2 56585 1 5003
2 56586 1 5003
2 56587 1 5003
2 56588 1 5003
2 56589 1 5005
2 56590 1 5005
2 56591 1 5006
2 56592 1 5006
2 56593 1 5006
2 56594 1 5006
2 56595 1 5006
2 56596 1 5006
2 56597 1 5006
2 56598 1 5007
2 56599 1 5007
2 56600 1 5008
2 56601 1 5008
2 56602 1 5016
2 56603 1 5016
2 56604 1 5016
2 56605 1 5016
2 56606 1 5016
2 56607 1 5017
2 56608 1 5017
2 56609 1 5017
2 56610 1 5017
2 56611 1 5017
2 56612 1 5017
2 56613 1 5017
2 56614 1 5017
2 56615 1 5024
2 56616 1 5024
2 56617 1 5024
2 56618 1 5024
2 56619 1 5024
2 56620 1 5024
2 56621 1 5036
2 56622 1 5036
2 56623 1 5036
2 56624 1 5036
2 56625 1 5036
2 56626 1 5036
2 56627 1 5036
2 56628 1 5036
2 56629 1 5036
2 56630 1 5036
2 56631 1 5036
2 56632 1 5047
2 56633 1 5047
2 56634 1 5047
2 56635 1 5047
2 56636 1 5047
2 56637 1 5047
2 56638 1 5047
2 56639 1 5050
2 56640 1 5050
2 56641 1 5057
2 56642 1 5057
2 56643 1 5057
2 56644 1 5057
2 56645 1 5057
2 56646 1 5057
2 56647 1 5066
2 56648 1 5066
2 56649 1 5067
2 56650 1 5067
2 56651 1 5068
2 56652 1 5068
2 56653 1 5068
2 56654 1 5080
2 56655 1 5080
2 56656 1 5080
2 56657 1 5080
2 56658 1 5080
2 56659 1 5080
2 56660 1 5080
2 56661 1 5080
2 56662 1 5080
2 56663 1 5080
2 56664 1 5080
2 56665 1 5081
2 56666 1 5081
2 56667 1 5081
2 56668 1 5092
2 56669 1 5092
2 56670 1 5092
2 56671 1 5092
2 56672 1 5092
2 56673 1 5092
2 56674 1 5092
2 56675 1 5092
2 56676 1 5092
2 56677 1 5092
2 56678 1 5092
2 56679 1 5092
2 56680 1 5092
2 56681 1 5092
2 56682 1 5092
2 56683 1 5092
2 56684 1 5092
2 56685 1 5093
2 56686 1 5093
2 56687 1 5093
2 56688 1 5093
2 56689 1 5093
2 56690 1 5093
2 56691 1 5093
2 56692 1 5094
2 56693 1 5094
2 56694 1 5094
2 56695 1 5094
2 56696 1 5094
2 56697 1 5094
2 56698 1 5094
2 56699 1 5096
2 56700 1 5096
2 56701 1 5107
2 56702 1 5107
2 56703 1 5107
2 56704 1 5107
2 56705 1 5107
2 56706 1 5107
2 56707 1 5107
2 56708 1 5107
2 56709 1 5107
2 56710 1 5107
2 56711 1 5108
2 56712 1 5108
2 56713 1 5108
2 56714 1 5108
2 56715 1 5108
2 56716 1 5108
2 56717 1 5108
2 56718 1 5108
2 56719 1 5108
2 56720 1 5108
2 56721 1 5108
2 56722 1 5108
2 56723 1 5109
2 56724 1 5109
2 56725 1 5110
2 56726 1 5110
2 56727 1 5111
2 56728 1 5111
2 56729 1 5115
2 56730 1 5115
2 56731 1 5116
2 56732 1 5116
2 56733 1 5116
2 56734 1 5116
2 56735 1 5116
2 56736 1 5116
2 56737 1 5117
2 56738 1 5117
2 56739 1 5117
2 56740 1 5120
2 56741 1 5120
2 56742 1 5120
2 56743 1 5127
2 56744 1 5127
2 56745 1 5127
2 56746 1 5127
2 56747 1 5127
2 56748 1 5127
2 56749 1 5130
2 56750 1 5130
2 56751 1 5130
2 56752 1 5130
2 56753 1 5130
2 56754 1 5130
2 56755 1 5130
2 56756 1 5130
2 56757 1 5130
2 56758 1 5130
2 56759 1 5130
2 56760 1 5130
2 56761 1 5130
2 56762 1 5131
2 56763 1 5131
2 56764 1 5140
2 56765 1 5140
2 56766 1 5140
2 56767 1 5140
2 56768 1 5140
2 56769 1 5140
2 56770 1 5141
2 56771 1 5141
2 56772 1 5141
2 56773 1 5141
2 56774 1 5141
2 56775 1 5141
2 56776 1 5141
2 56777 1 5141
2 56778 1 5142
2 56779 1 5142
2 56780 1 5142
2 56781 1 5150
2 56782 1 5150
2 56783 1 5150
2 56784 1 5150
2 56785 1 5150
2 56786 1 5150
2 56787 1 5154
2 56788 1 5154
2 56789 1 5154
2 56790 1 5154
2 56791 1 5155
2 56792 1 5155
2 56793 1 5155
2 56794 1 5155
2 56795 1 5155
2 56796 1 5155
2 56797 1 5155
2 56798 1 5155
2 56799 1 5155
2 56800 1 5155
2 56801 1 5155
2 56802 1 5155
2 56803 1 5155
2 56804 1 5155
2 56805 1 5156
2 56806 1 5156
2 56807 1 5158
2 56808 1 5158
2 56809 1 5159
2 56810 1 5159
2 56811 1 5159
2 56812 1 5171
2 56813 1 5171
2 56814 1 5171
2 56815 1 5171
2 56816 1 5171
2 56817 1 5171
2 56818 1 5171
2 56819 1 5171
2 56820 1 5171
2 56821 1 5172
2 56822 1 5172
2 56823 1 5172
2 56824 1 5176
2 56825 1 5176
2 56826 1 5176
2 56827 1 5180
2 56828 1 5180
2 56829 1 5180
2 56830 1 5180
2 56831 1 5180
2 56832 1 5180
2 56833 1 5180
2 56834 1 5180
2 56835 1 5188
2 56836 1 5188
2 56837 1 5190
2 56838 1 5190
2 56839 1 5190
2 56840 1 5190
2 56841 1 5190
2 56842 1 5190
2 56843 1 5190
2 56844 1 5190
2 56845 1 5190
2 56846 1 5190
2 56847 1 5190
2 56848 1 5190
2 56849 1 5198
2 56850 1 5198
2 56851 1 5200
2 56852 1 5200
2 56853 1 5206
2 56854 1 5206
2 56855 1 5206
2 56856 1 5206
2 56857 1 5206
2 56858 1 5206
2 56859 1 5206
2 56860 1 5206
2 56861 1 5206
2 56862 1 5206
2 56863 1 5206
2 56864 1 5206
2 56865 1 5206
2 56866 1 5206
2 56867 1 5206
2 56868 1 5206
2 56869 1 5206
2 56870 1 5206
2 56871 1 5207
2 56872 1 5207
2 56873 1 5207
2 56874 1 5214
2 56875 1 5214
2 56876 1 5215
2 56877 1 5215
2 56878 1 5226
2 56879 1 5226
2 56880 1 5227
2 56881 1 5227
2 56882 1 5227
2 56883 1 5227
2 56884 1 5227
2 56885 1 5227
2 56886 1 5227
2 56887 1 5227
2 56888 1 5227
2 56889 1 5227
2 56890 1 5227
2 56891 1 5227
2 56892 1 5227
2 56893 1 5227
2 56894 1 5233
2 56895 1 5233
2 56896 1 5248
2 56897 1 5248
2 56898 1 5248
2 56899 1 5248
2 56900 1 5248
2 56901 1 5248
2 56902 1 5249
2 56903 1 5249
2 56904 1 5249
2 56905 1 5249
2 56906 1 5249
2 56907 1 5249
2 56908 1 5250
2 56909 1 5250
2 56910 1 5250
2 56911 1 5250
2 56912 1 5250
2 56913 1 5265
2 56914 1 5265
2 56915 1 5265
2 56916 1 5265
2 56917 1 5265
2 56918 1 5265
2 56919 1 5265
2 56920 1 5266
2 56921 1 5266
2 56922 1 5269
2 56923 1 5269
2 56924 1 5271
2 56925 1 5271
2 56926 1 5272
2 56927 1 5272
2 56928 1 5273
2 56929 1 5273
2 56930 1 5281
2 56931 1 5281
2 56932 1 5281
2 56933 1 5282
2 56934 1 5282
2 56935 1 5289
2 56936 1 5289
2 56937 1 5289
2 56938 1 5289
2 56939 1 5289
2 56940 1 5289
2 56941 1 5289
2 56942 1 5293
2 56943 1 5293
2 56944 1 5303
2 56945 1 5303
2 56946 1 5303
2 56947 1 5303
2 56948 1 5304
2 56949 1 5304
2 56950 1 5304
2 56951 1 5304
2 56952 1 5304
2 56953 1 5304
2 56954 1 5304
2 56955 1 5304
2 56956 1 5312
2 56957 1 5312
2 56958 1 5312
2 56959 1 5312
2 56960 1 5312
2 56961 1 5312
2 56962 1 5312
2 56963 1 5312
2 56964 1 5312
2 56965 1 5312
2 56966 1 5312
2 56967 1 5313
2 56968 1 5313
2 56969 1 5313
2 56970 1 5313
2 56971 1 5313
2 56972 1 5313
2 56973 1 5313
2 56974 1 5314
2 56975 1 5314
2 56976 1 5314
2 56977 1 5314
2 56978 1 5315
2 56979 1 5315
2 56980 1 5319
2 56981 1 5319
2 56982 1 5319
2 56983 1 5319
2 56984 1 5319
2 56985 1 5319
2 56986 1 5319
2 56987 1 5319
2 56988 1 5319
2 56989 1 5319
2 56990 1 5319
2 56991 1 5319
2 56992 1 5319
2 56993 1 5319
2 56994 1 5319
2 56995 1 5319
2 56996 1 5331
2 56997 1 5331
2 56998 1 5331
2 56999 1 5332
2 57000 1 5332
2 57001 1 5335
2 57002 1 5335
2 57003 1 5335
2 57004 1 5335
2 57005 1 5336
2 57006 1 5336
2 57007 1 5336
2 57008 1 5336
2 57009 1 5336
2 57010 1 5336
2 57011 1 5336
2 57012 1 5336
2 57013 1 5336
2 57014 1 5336
2 57015 1 5336
2 57016 1 5336
2 57017 1 5336
2 57018 1 5336
2 57019 1 5336
2 57020 1 5336
2 57021 1 5338
2 57022 1 5338
2 57023 1 5338
2 57024 1 5341
2 57025 1 5341
2 57026 1 5341
2 57027 1 5341
2 57028 1 5341
2 57029 1 5341
2 57030 1 5341
2 57031 1 5341
2 57032 1 5341
2 57033 1 5341
2 57034 1 5341
2 57035 1 5341
2 57036 1 5348
2 57037 1 5348
2 57038 1 5348
2 57039 1 5348
2 57040 1 5348
2 57041 1 5348
2 57042 1 5348
2 57043 1 5348
2 57044 1 5348
2 57045 1 5348
2 57046 1 5348
2 57047 1 5348
2 57048 1 5348
2 57049 1 5348
2 57050 1 5348
2 57051 1 5348
2 57052 1 5348
2 57053 1 5348
2 57054 1 5348
2 57055 1 5348
2 57056 1 5348
2 57057 1 5348
2 57058 1 5348
2 57059 1 5348
2 57060 1 5348
2 57061 1 5348
2 57062 1 5348
2 57063 1 5348
2 57064 1 5348
2 57065 1 5348
2 57066 1 5348
2 57067 1 5348
2 57068 1 5348
2 57069 1 5348
2 57070 1 5348
2 57071 1 5348
2 57072 1 5348
2 57073 1 5348
2 57074 1 5349
2 57075 1 5349
2 57076 1 5349
2 57077 1 5349
2 57078 1 5349
2 57079 1 5349
2 57080 1 5349
2 57081 1 5349
2 57082 1 5349
2 57083 1 5349
2 57084 1 5349
2 57085 1 5350
2 57086 1 5350
2 57087 1 5350
2 57088 1 5353
2 57089 1 5353
2 57090 1 5353
2 57091 1 5353
2 57092 1 5353
2 57093 1 5353
2 57094 1 5353
2 57095 1 5353
2 57096 1 5353
2 57097 1 5353
2 57098 1 5353
2 57099 1 5354
2 57100 1 5354
2 57101 1 5354
2 57102 1 5354
2 57103 1 5354
2 57104 1 5354
2 57105 1 5354
2 57106 1 5358
2 57107 1 5358
2 57108 1 5358
2 57109 1 5361
2 57110 1 5361
2 57111 1 5362
2 57112 1 5362
2 57113 1 5362
2 57114 1 5366
2 57115 1 5366
2 57116 1 5366
2 57117 1 5366
2 57118 1 5379
2 57119 1 5379
2 57120 1 5380
2 57121 1 5380
2 57122 1 5380
2 57123 1 5384
2 57124 1 5384
2 57125 1 5384
2 57126 1 5384
2 57127 1 5384
2 57128 1 5398
2 57129 1 5398
2 57130 1 5398
2 57131 1 5402
2 57132 1 5402
2 57133 1 5402
2 57134 1 5402
2 57135 1 5402
2 57136 1 5402
2 57137 1 5402
2 57138 1 5403
2 57139 1 5403
2 57140 1 5403
2 57141 1 5404
2 57142 1 5404
2 57143 1 5411
2 57144 1 5411
2 57145 1 5411
2 57146 1 5411
2 57147 1 5411
2 57148 1 5411
2 57149 1 5412
2 57150 1 5412
2 57151 1 5412
2 57152 1 5412
2 57153 1 5412
2 57154 1 5412
2 57155 1 5412
2 57156 1 5415
2 57157 1 5415
2 57158 1 5415
2 57159 1 5415
2 57160 1 5415
2 57161 1 5416
2 57162 1 5416
2 57163 1 5416
2 57164 1 5416
2 57165 1 5416
2 57166 1 5417
2 57167 1 5417
2 57168 1 5417
2 57169 1 5417
2 57170 1 5417
2 57171 1 5417
2 57172 1 5417
2 57173 1 5417
2 57174 1 5417
2 57175 1 5418
2 57176 1 5418
2 57177 1 5418
2 57178 1 5418
2 57179 1 5418
2 57180 1 5418
2 57181 1 5418
2 57182 1 5426
2 57183 1 5426
2 57184 1 5427
2 57185 1 5427
2 57186 1 5427
2 57187 1 5427
2 57188 1 5427
2 57189 1 5443
2 57190 1 5443
2 57191 1 5443
2 57192 1 5443
2 57193 1 5443
2 57194 1 5443
2 57195 1 5443
2 57196 1 5443
2 57197 1 5443
2 57198 1 5443
2 57199 1 5443
2 57200 1 5443
2 57201 1 5443
2 57202 1 5443
2 57203 1 5443
2 57204 1 5443
2 57205 1 5443
2 57206 1 5443
2 57207 1 5443
2 57208 1 5443
2 57209 1 5443
2 57210 1 5443
2 57211 1 5443
2 57212 1 5443
2 57213 1 5443
2 57214 1 5443
2 57215 1 5443
2 57216 1 5443
2 57217 1 5443
2 57218 1 5443
2 57219 1 5443
2 57220 1 5443
2 57221 1 5444
2 57222 1 5444
2 57223 1 5444
2 57224 1 5444
2 57225 1 5445
2 57226 1 5445
2 57227 1 5445
2 57228 1 5445
2 57229 1 5448
2 57230 1 5448
2 57231 1 5448
2 57232 1 5448
2 57233 1 5448
2 57234 1 5448
2 57235 1 5448
2 57236 1 5448
2 57237 1 5448
2 57238 1 5448
2 57239 1 5448
2 57240 1 5449
2 57241 1 5449
2 57242 1 5449
2 57243 1 5449
2 57244 1 5449
2 57245 1 5449
2 57246 1 5449
2 57247 1 5449
2 57248 1 5449
2 57249 1 5449
2 57250 1 5449
2 57251 1 5449
2 57252 1 5449
2 57253 1 5449
2 57254 1 5449
2 57255 1 5449
2 57256 1 5449
2 57257 1 5449
2 57258 1 5449
2 57259 1 5449
2 57260 1 5449
2 57261 1 5449
2 57262 1 5449
2 57263 1 5449
2 57264 1 5449
2 57265 1 5449
2 57266 1 5449
2 57267 1 5449
2 57268 1 5449
2 57269 1 5449
2 57270 1 5449
2 57271 1 5449
2 57272 1 5449
2 57273 1 5449
2 57274 1 5449
2 57275 1 5449
2 57276 1 5449
2 57277 1 5449
2 57278 1 5449
2 57279 1 5449
2 57280 1 5449
2 57281 1 5450
2 57282 1 5450
2 57283 1 5450
2 57284 1 5450
2 57285 1 5454
2 57286 1 5454
2 57287 1 5457
2 57288 1 5457
2 57289 1 5457
2 57290 1 5457
2 57291 1 5457
2 57292 1 5457
2 57293 1 5457
2 57294 1 5457
2 57295 1 5457
2 57296 1 5457
2 57297 1 5465
2 57298 1 5465
2 57299 1 5465
2 57300 1 5465
2 57301 1 5465
2 57302 1 5465
2 57303 1 5465
2 57304 1 5465
2 57305 1 5465
2 57306 1 5465
2 57307 1 5465
2 57308 1 5474
2 57309 1 5474
2 57310 1 5475
2 57311 1 5475
2 57312 1 5475
2 57313 1 5475
2 57314 1 5475
2 57315 1 5475
2 57316 1 5476
2 57317 1 5476
2 57318 1 5482
2 57319 1 5482
2 57320 1 5484
2 57321 1 5484
2 57322 1 5485
2 57323 1 5485
2 57324 1 5485
2 57325 1 5485
2 57326 1 5485
2 57327 1 5486
2 57328 1 5486
2 57329 1 5486
2 57330 1 5486
2 57331 1 5486
2 57332 1 5486
2 57333 1 5494
2 57334 1 5494
2 57335 1 5494
2 57336 1 5495
2 57337 1 5495
2 57338 1 5495
2 57339 1 5495
2 57340 1 5498
2 57341 1 5498
2 57342 1 5498
2 57343 1 5498
2 57344 1 5499
2 57345 1 5499
2 57346 1 5507
2 57347 1 5507
2 57348 1 5507
2 57349 1 5508
2 57350 1 5508
2 57351 1 5510
2 57352 1 5510
2 57353 1 5516
2 57354 1 5516
2 57355 1 5517
2 57356 1 5517
2 57357 1 5525
2 57358 1 5525
2 57359 1 5525
2 57360 1 5525
2 57361 1 5525
2 57362 1 5525
2 57363 1 5526
2 57364 1 5526
2 57365 1 5526
2 57366 1 5526
2 57367 1 5526
2 57368 1 5527
2 57369 1 5527
2 57370 1 5532
2 57371 1 5532
2 57372 1 5539
2 57373 1 5539
2 57374 1 5542
2 57375 1 5542
2 57376 1 5542
2 57377 1 5542
2 57378 1 5542
2 57379 1 5543
2 57380 1 5543
2 57381 1 5546
2 57382 1 5546
2 57383 1 5546
2 57384 1 5546
2 57385 1 5547
2 57386 1 5547
2 57387 1 5558
2 57388 1 5558
2 57389 1 5558
2 57390 1 5558
2 57391 1 5558
2 57392 1 5558
2 57393 1 5558
2 57394 1 5558
2 57395 1 5558
2 57396 1 5559
2 57397 1 5559
2 57398 1 5560
2 57399 1 5560
2 57400 1 5560
2 57401 1 5571
2 57402 1 5571
2 57403 1 5571
2 57404 1 5571
2 57405 1 5571
2 57406 1 5571
2 57407 1 5578
2 57408 1 5578
2 57409 1 5579
2 57410 1 5579
2 57411 1 5579
2 57412 1 5579
2 57413 1 5579
2 57414 1 5580
2 57415 1 5580
2 57416 1 5581
2 57417 1 5581
2 57418 1 5582
2 57419 1 5582
2 57420 1 5588
2 57421 1 5588
2 57422 1 5598
2 57423 1 5598
2 57424 1 5606
2 57425 1 5606
2 57426 1 5606
2 57427 1 5606
2 57428 1 5606
2 57429 1 5606
2 57430 1 5606
2 57431 1 5606
2 57432 1 5613
2 57433 1 5613
2 57434 1 5613
2 57435 1 5613
2 57436 1 5613
2 57437 1 5613
2 57438 1 5613
2 57439 1 5614
2 57440 1 5614
2 57441 1 5614
2 57442 1 5621
2 57443 1 5621
2 57444 1 5621
2 57445 1 5621
2 57446 1 5621
2 57447 1 5621
2 57448 1 5636
2 57449 1 5636
2 57450 1 5636
2 57451 1 5636
2 57452 1 5636
2 57453 1 5636
2 57454 1 5636
2 57455 1 5636
2 57456 1 5637
2 57457 1 5637
2 57458 1 5640
2 57459 1 5640
2 57460 1 5641
2 57461 1 5641
2 57462 1 5643
2 57463 1 5643
2 57464 1 5646
2 57465 1 5646
2 57466 1 5646
2 57467 1 5647
2 57468 1 5647
2 57469 1 5647
2 57470 1 5647
2 57471 1 5647
2 57472 1 5647
2 57473 1 5649
2 57474 1 5649
2 57475 1 5649
2 57476 1 5649
2 57477 1 5649
2 57478 1 5649
2 57479 1 5649
2 57480 1 5649
2 57481 1 5649
2 57482 1 5649
2 57483 1 5649
2 57484 1 5649
2 57485 1 5649
2 57486 1 5649
2 57487 1 5649
2 57488 1 5649
2 57489 1 5649
2 57490 1 5650
2 57491 1 5650
2 57492 1 5651
2 57493 1 5651
2 57494 1 5655
2 57495 1 5655
2 57496 1 5662
2 57497 1 5662
2 57498 1 5662
2 57499 1 5663
2 57500 1 5663
2 57501 1 5663
2 57502 1 5663
2 57503 1 5663
2 57504 1 5663
2 57505 1 5663
2 57506 1 5663
2 57507 1 5663
2 57508 1 5667
2 57509 1 5667
2 57510 1 5671
2 57511 1 5671
2 57512 1 5671
2 57513 1 5673
2 57514 1 5673
2 57515 1 5677
2 57516 1 5677
2 57517 1 5677
2 57518 1 5677
2 57519 1 5702
2 57520 1 5702
2 57521 1 5702
2 57522 1 5715
2 57523 1 5715
2 57524 1 5715
2 57525 1 5715
2 57526 1 5715
2 57527 1 5729
2 57528 1 5729
2 57529 1 5735
2 57530 1 5735
2 57531 1 5735
2 57532 1 5736
2 57533 1 5736
2 57534 1 5757
2 57535 1 5757
2 57536 1 5757
2 57537 1 5759
2 57538 1 5759
2 57539 1 5762
2 57540 1 5762
2 57541 1 5762
2 57542 1 5762
2 57543 1 5762
2 57544 1 5762
2 57545 1 5765
2 57546 1 5765
2 57547 1 5765
2 57548 1 5765
2 57549 1 5765
2 57550 1 5765
2 57551 1 5766
2 57552 1 5766
2 57553 1 5770
2 57554 1 5770
2 57555 1 5771
2 57556 1 5771
2 57557 1 5790
2 57558 1 5790
2 57559 1 5797
2 57560 1 5797
2 57561 1 5814
2 57562 1 5814
2 57563 1 5815
2 57564 1 5815
2 57565 1 5818
2 57566 1 5818
2 57567 1 5818
2 57568 1 5818
2 57569 1 5818
2 57570 1 5818
2 57571 1 5818
2 57572 1 5818
2 57573 1 5818
2 57574 1 5818
2 57575 1 5818
2 57576 1 5818
2 57577 1 5818
2 57578 1 5818
2 57579 1 5819
2 57580 1 5819
2 57581 1 5819
2 57582 1 5819
2 57583 1 5820
2 57584 1 5820
2 57585 1 5837
2 57586 1 5837
2 57587 1 5837
2 57588 1 5837
2 57589 1 5837
2 57590 1 5844
2 57591 1 5844
2 57592 1 5844
2 57593 1 5844
2 57594 1 5844
2 57595 1 5844
2 57596 1 5844
2 57597 1 5844
2 57598 1 5844
2 57599 1 5844
2 57600 1 5844
2 57601 1 5844
2 57602 1 5844
2 57603 1 5844
2 57604 1 5844
2 57605 1 5849
2 57606 1 5849
2 57607 1 5863
2 57608 1 5863
2 57609 1 5863
2 57610 1 5863
2 57611 1 5866
2 57612 1 5866
2 57613 1 5866
2 57614 1 5867
2 57615 1 5867
2 57616 1 5867
2 57617 1 5867
2 57618 1 5867
2 57619 1 5878
2 57620 1 5878
2 57621 1 5878
2 57622 1 5878
2 57623 1 5878
2 57624 1 5878
2 57625 1 5878
2 57626 1 5878
2 57627 1 5878
2 57628 1 5878
2 57629 1 5878
2 57630 1 5878
2 57631 1 5878
2 57632 1 5878
2 57633 1 5878
2 57634 1 5878
2 57635 1 5878
2 57636 1 5878
2 57637 1 5878
2 57638 1 5878
2 57639 1 5878
2 57640 1 5878
2 57641 1 5878
2 57642 1 5878
2 57643 1 5878
2 57644 1 5878
2 57645 1 5878
2 57646 1 5878
2 57647 1 5878
2 57648 1 5878
2 57649 1 5878
2 57650 1 5878
2 57651 1 5878
2 57652 1 5878
2 57653 1 5878
2 57654 1 5878
2 57655 1 5878
2 57656 1 5878
2 57657 1 5878
2 57658 1 5878
2 57659 1 5878
2 57660 1 5878
2 57661 1 5878
2 57662 1 5878
2 57663 1 5878
2 57664 1 5878
2 57665 1 5878
2 57666 1 5878
2 57667 1 5878
2 57668 1 5879
2 57669 1 5879
2 57670 1 5879
2 57671 1 5879
2 57672 1 5879
2 57673 1 5896
2 57674 1 5896
2 57675 1 5906
2 57676 1 5906
2 57677 1 5911
2 57678 1 5911
2 57679 1 5911
2 57680 1 5911
2 57681 1 5911
2 57682 1 5911
2 57683 1 5911
2 57684 1 5911
2 57685 1 5911
2 57686 1 5911
2 57687 1 5911
2 57688 1 5911
2 57689 1 5911
2 57690 1 5923
2 57691 1 5923
2 57692 1 5923
2 57693 1 5949
2 57694 1 5949
2 57695 1 5949
2 57696 1 5949
2 57697 1 5949
2 57698 1 5950
2 57699 1 5950
2 57700 1 5950
2 57701 1 5952
2 57702 1 5952
2 57703 1 5954
2 57704 1 5954
2 57705 1 5954
2 57706 1 5954
2 57707 1 5959
2 57708 1 5959
2 57709 1 5960
2 57710 1 5960
2 57711 1 5960
2 57712 1 5960
2 57713 1 5960
2 57714 1 5960
2 57715 1 5960
2 57716 1 5963
2 57717 1 5963
2 57718 1 5963
2 57719 1 5963
2 57720 1 5963
2 57721 1 5966
2 57722 1 5966
2 57723 1 5966
2 57724 1 5966
2 57725 1 5966
2 57726 1 5966
2 57727 1 5966
2 57728 1 5966
2 57729 1 5966
2 57730 1 5966
2 57731 1 5967
2 57732 1 5967
2 57733 1 5967
2 57734 1 5971
2 57735 1 5971
2 57736 1 5977
2 57737 1 5977
2 57738 1 5985
2 57739 1 5985
2 57740 1 5985
2 57741 1 5985
2 57742 1 5986
2 57743 1 5986
2 57744 1 5988
2 57745 1 5988
2 57746 1 5988
2 57747 1 5989
2 57748 1 5989
2 57749 1 5992
2 57750 1 5992
2 57751 1 5993
2 57752 1 5993
2 57753 1 5993
2 57754 1 5993
2 57755 1 5993
2 57756 1 5995
2 57757 1 5995
2 57758 1 6000
2 57759 1 6000
2 57760 1 6000
2 57761 1 6002
2 57762 1 6002
2 57763 1 6002
2 57764 1 6002
2 57765 1 6002
2 57766 1 6003
2 57767 1 6003
2 57768 1 6003
2 57769 1 6003
2 57770 1 6003
2 57771 1 6011
2 57772 1 6011
2 57773 1 6012
2 57774 1 6012
2 57775 1 6012
2 57776 1 6021
2 57777 1 6021
2 57778 1 6021
2 57779 1 6023
2 57780 1 6023
2 57781 1 6023
2 57782 1 6023
2 57783 1 6024
2 57784 1 6024
2 57785 1 6034
2 57786 1 6034
2 57787 1 6034
2 57788 1 6034
2 57789 1 6034
2 57790 1 6034
2 57791 1 6035
2 57792 1 6035
2 57793 1 6036
2 57794 1 6036
2 57795 1 6042
2 57796 1 6042
2 57797 1 6042
2 57798 1 6042
2 57799 1 6042
2 57800 1 6043
2 57801 1 6043
2 57802 1 6043
2 57803 1 6047
2 57804 1 6047
2 57805 1 6048
2 57806 1 6048
2 57807 1 6048
2 57808 1 6048
2 57809 1 6048
2 57810 1 6048
2 57811 1 6048
2 57812 1 6048
2 57813 1 6048
2 57814 1 6048
2 57815 1 6048
2 57816 1 6048
2 57817 1 6050
2 57818 1 6050
2 57819 1 6052
2 57820 1 6052
2 57821 1 6052
2 57822 1 6052
2 57823 1 6052
2 57824 1 6052
2 57825 1 6052
2 57826 1 6052
2 57827 1 6053
2 57828 1 6053
2 57829 1 6053
2 57830 1 6053
2 57831 1 6069
2 57832 1 6069
2 57833 1 6069
2 57834 1 6069
2 57835 1 6069
2 57836 1 6069
2 57837 1 6070
2 57838 1 6070
2 57839 1 6070
2 57840 1 6070
2 57841 1 6071
2 57842 1 6071
2 57843 1 6071
2 57844 1 6073
2 57845 1 6073
2 57846 1 6075
2 57847 1 6075
2 57848 1 6075
2 57849 1 6075
2 57850 1 6076
2 57851 1 6076
2 57852 1 6076
2 57853 1 6076
2 57854 1 6080
2 57855 1 6080
2 57856 1 6080
2 57857 1 6080
2 57858 1 6080
2 57859 1 6080
2 57860 1 6080
2 57861 1 6080
2 57862 1 6080
2 57863 1 6080
2 57864 1 6081
2 57865 1 6081
2 57866 1 6084
2 57867 1 6084
2 57868 1 6113
2 57869 1 6113
2 57870 1 6113
2 57871 1 6115
2 57872 1 6115
2 57873 1 6127
2 57874 1 6127
2 57875 1 6129
2 57876 1 6129
2 57877 1 6130
2 57878 1 6130
2 57879 1 6132
2 57880 1 6132
2 57881 1 6149
2 57882 1 6149
2 57883 1 6156
2 57884 1 6156
2 57885 1 6162
2 57886 1 6162
2 57887 1 6162
2 57888 1 6162
2 57889 1 6162
2 57890 1 6162
2 57891 1 6162
2 57892 1 6166
2 57893 1 6166
2 57894 1 6166
2 57895 1 6167
2 57896 1 6167
2 57897 1 6172
2 57898 1 6172
2 57899 1 6173
2 57900 1 6173
2 57901 1 6173
2 57902 1 6174
2 57903 1 6174
2 57904 1 6181
2 57905 1 6181
2 57906 1 6181
2 57907 1 6181
2 57908 1 6181
2 57909 1 6181
2 57910 1 6182
2 57911 1 6182
2 57912 1 6183
2 57913 1 6183
2 57914 1 6183
2 57915 1 6183
2 57916 1 6183
2 57917 1 6183
2 57918 1 6183
2 57919 1 6183
2 57920 1 6183
2 57921 1 6184
2 57922 1 6184
2 57923 1 6185
2 57924 1 6185
2 57925 1 6193
2 57926 1 6193
2 57927 1 6202
2 57928 1 6202
2 57929 1 6202
2 57930 1 6202
2 57931 1 6203
2 57932 1 6203
2 57933 1 6203
2 57934 1 6205
2 57935 1 6205
2 57936 1 6205
2 57937 1 6205
2 57938 1 6205
2 57939 1 6205
2 57940 1 6205
2 57941 1 6217
2 57942 1 6217
2 57943 1 6217
2 57944 1 6218
2 57945 1 6218
2 57946 1 6218
2 57947 1 6218
2 57948 1 6218
2 57949 1 6219
2 57950 1 6219
2 57951 1 6219
2 57952 1 6220
2 57953 1 6220
2 57954 1 6220
2 57955 1 6235
2 57956 1 6235
2 57957 1 6235
2 57958 1 6235
2 57959 1 6235
2 57960 1 6235
2 57961 1 6235
2 57962 1 6235
2 57963 1 6235
2 57964 1 6235
2 57965 1 6236
2 57966 1 6236
2 57967 1 6236
2 57968 1 6236
2 57969 1 6236
2 57970 1 6236
2 57971 1 6237
2 57972 1 6237
2 57973 1 6237
2 57974 1 6237
2 57975 1 6237
2 57976 1 6237
2 57977 1 6237
2 57978 1 6237
2 57979 1 6237
2 57980 1 6237
2 57981 1 6238
2 57982 1 6238
2 57983 1 6238
2 57984 1 6240
2 57985 1 6240
2 57986 1 6241
2 57987 1 6241
2 57988 1 6241
2 57989 1 6241
2 57990 1 6241
2 57991 1 6242
2 57992 1 6242
2 57993 1 6242
2 57994 1 6254
2 57995 1 6254
2 57996 1 6254
2 57997 1 6254
2 57998 1 6254
2 57999 1 6254
2 58000 1 6254
2 58001 1 6254
2 58002 1 6254
2 58003 1 6254
2 58004 1 6254
2 58005 1 6256
2 58006 1 6256
2 58007 1 6256
2 58008 1 6256
2 58009 1 6256
2 58010 1 6256
2 58011 1 6256
2 58012 1 6256
2 58013 1 6256
2 58014 1 6256
2 58015 1 6258
2 58016 1 6258
2 58017 1 6259
2 58018 1 6259
2 58019 1 6259
2 58020 1 6259
2 58021 1 6259
2 58022 1 6259
2 58023 1 6259
2 58024 1 6259
2 58025 1 6259
2 58026 1 6259
2 58027 1 6259
2 58028 1 6259
2 58029 1 6259
2 58030 1 6259
2 58031 1 6259
2 58032 1 6259
2 58033 1 6259
2 58034 1 6259
2 58035 1 6259
2 58036 1 6259
2 58037 1 6259
2 58038 1 6259
2 58039 1 6259
2 58040 1 6259
2 58041 1 6259
2 58042 1 6259
2 58043 1 6259
2 58044 1 6259
2 58045 1 6259
2 58046 1 6259
2 58047 1 6259
2 58048 1 6259
2 58049 1 6259
2 58050 1 6259
2 58051 1 6259
2 58052 1 6259
2 58053 1 6259
2 58054 1 6259
2 58055 1 6259
2 58056 1 6259
2 58057 1 6259
2 58058 1 6259
2 58059 1 6259
2 58060 1 6259
2 58061 1 6259
2 58062 1 6259
2 58063 1 6259
2 58064 1 6259
2 58065 1 6266
2 58066 1 6266
2 58067 1 6267
2 58068 1 6267
2 58069 1 6267
2 58070 1 6267
2 58071 1 6275
2 58072 1 6275
2 58073 1 6282
2 58074 1 6282
2 58075 1 6282
2 58076 1 6293
2 58077 1 6293
2 58078 1 6293
2 58079 1 6302
2 58080 1 6302
2 58081 1 6302
2 58082 1 6302
2 58083 1 6302
2 58084 1 6302
2 58085 1 6304
2 58086 1 6304
2 58087 1 6304
2 58088 1 6304
2 58089 1 6304
2 58090 1 6305
2 58091 1 6305
2 58092 1 6306
2 58093 1 6306
2 58094 1 6309
2 58095 1 6309
2 58096 1 6309
2 58097 1 6310
2 58098 1 6310
2 58099 1 6310
2 58100 1 6310
2 58101 1 6320
2 58102 1 6320
2 58103 1 6320
2 58104 1 6321
2 58105 1 6321
2 58106 1 6321
2 58107 1 6322
2 58108 1 6322
2 58109 1 6322
2 58110 1 6322
2 58111 1 6322
2 58112 1 6339
2 58113 1 6339
2 58114 1 6360
2 58115 1 6360
2 58116 1 6360
2 58117 1 6360
2 58118 1 6364
2 58119 1 6364
2 58120 1 6371
2 58121 1 6371
2 58122 1 6372
2 58123 1 6372
2 58124 1 6372
2 58125 1 6379
2 58126 1 6379
2 58127 1 6379
2 58128 1 6380
2 58129 1 6380
2 58130 1 6392
2 58131 1 6392
2 58132 1 6392
2 58133 1 6392
2 58134 1 6392
2 58135 1 6409
2 58136 1 6409
2 58137 1 6409
2 58138 1 6410
2 58139 1 6410
2 58140 1 6410
2 58141 1 6410
2 58142 1 6410
2 58143 1 6410
2 58144 1 6414
2 58145 1 6414
2 58146 1 6415
2 58147 1 6415
2 58148 1 6416
2 58149 1 6416
2 58150 1 6424
2 58151 1 6424
2 58152 1 6424
2 58153 1 6425
2 58154 1 6425
2 58155 1 6443
2 58156 1 6443
2 58157 1 6443
2 58158 1 6443
2 58159 1 6444
2 58160 1 6444
2 58161 1 6446
2 58162 1 6446
2 58163 1 6446
2 58164 1 6446
2 58165 1 6448
2 58166 1 6448
2 58167 1 6463
2 58168 1 6463
2 58169 1 6464
2 58170 1 6464
2 58171 1 6466
2 58172 1 6466
2 58173 1 6466
2 58174 1 6467
2 58175 1 6467
2 58176 1 6482
2 58177 1 6482
2 58178 1 6482
2 58179 1 6482
2 58180 1 6490
2 58181 1 6490
2 58182 1 6490
2 58183 1 6490
2 58184 1 6491
2 58185 1 6491
2 58186 1 6491
2 58187 1 6500
2 58188 1 6500
2 58189 1 6500
2 58190 1 6502
2 58191 1 6502
2 58192 1 6502
2 58193 1 6502
2 58194 1 6505
2 58195 1 6505
2 58196 1 6508
2 58197 1 6508
2 58198 1 6510
2 58199 1 6510
2 58200 1 6511
2 58201 1 6511
2 58202 1 6517
2 58203 1 6517
2 58204 1 6518
2 58205 1 6518
2 58206 1 6525
2 58207 1 6525
2 58208 1 6538
2 58209 1 6538
2 58210 1 6538
2 58211 1 6538
2 58212 1 6538
2 58213 1 6539
2 58214 1 6539
2 58215 1 6539
2 58216 1 6539
2 58217 1 6539
2 58218 1 6541
2 58219 1 6541
2 58220 1 6545
2 58221 1 6545
2 58222 1 6546
2 58223 1 6546
2 58224 1 6546
2 58225 1 6546
2 58226 1 6549
2 58227 1 6549
2 58228 1 6561
2 58229 1 6561
2 58230 1 6562
2 58231 1 6562
2 58232 1 6566
2 58233 1 6566
2 58234 1 6599
2 58235 1 6599
2 58236 1 6600
2 58237 1 6600
2 58238 1 6608
2 58239 1 6608
2 58240 1 6608
2 58241 1 6608
2 58242 1 6608
2 58243 1 6608
2 58244 1 6608
2 58245 1 6611
2 58246 1 6611
2 58247 1 6611
2 58248 1 6611
2 58249 1 6611
2 58250 1 6611
2 58251 1 6611
2 58252 1 6611
2 58253 1 6611
2 58254 1 6611
2 58255 1 6612
2 58256 1 6612
2 58257 1 6612
2 58258 1 6612
2 58259 1 6625
2 58260 1 6625
2 58261 1 6625
2 58262 1 6625
2 58263 1 6626
2 58264 1 6626
2 58265 1 6626
2 58266 1 6627
2 58267 1 6627
2 58268 1 6627
2 58269 1 6627
2 58270 1 6627
2 58271 1 6627
2 58272 1 6627
2 58273 1 6627
2 58274 1 6628
2 58275 1 6628
2 58276 1 6628
2 58277 1 6628
2 58278 1 6628
2 58279 1 6628
2 58280 1 6628
2 58281 1 6632
2 58282 1 6632
2 58283 1 6632
2 58284 1 6632
2 58285 1 6632
2 58286 1 6632
2 58287 1 6632
2 58288 1 6633
2 58289 1 6633
2 58290 1 6634
2 58291 1 6634
2 58292 1 6635
2 58293 1 6635
2 58294 1 6635
2 58295 1 6635
2 58296 1 6635
2 58297 1 6636
2 58298 1 6636
2 58299 1 6636
2 58300 1 6636
2 58301 1 6636
2 58302 1 6636
2 58303 1 6636
2 58304 1 6636
2 58305 1 6636
2 58306 1 6636
2 58307 1 6636
2 58308 1 6636
2 58309 1 6636
2 58310 1 6636
2 58311 1 6661
2 58312 1 6661
2 58313 1 6664
2 58314 1 6664
2 58315 1 6665
2 58316 1 6665
2 58317 1 6673
2 58318 1 6673
2 58319 1 6673
2 58320 1 6674
2 58321 1 6674
2 58322 1 6689
2 58323 1 6689
2 58324 1 6691
2 58325 1 6691
2 58326 1 6691
2 58327 1 6705
2 58328 1 6705
2 58329 1 6732
2 58330 1 6732
2 58331 1 6732
2 58332 1 6732
2 58333 1 6733
2 58334 1 6733
2 58335 1 6733
2 58336 1 6733
2 58337 1 6733
2 58338 1 6733
2 58339 1 6734
2 58340 1 6734
2 58341 1 6743
2 58342 1 6743
2 58343 1 6743
2 58344 1 6745
2 58345 1 6745
2 58346 1 6753
2 58347 1 6753
2 58348 1 6754
2 58349 1 6754
2 58350 1 6767
2 58351 1 6767
2 58352 1 6775
2 58353 1 6775
2 58354 1 6775
2 58355 1 6775
2 58356 1 6777
2 58357 1 6777
2 58358 1 6777
2 58359 1 6796
2 58360 1 6796
2 58361 1 6797
2 58362 1 6797
2 58363 1 6803
2 58364 1 6803
2 58365 1 6814
2 58366 1 6814
2 58367 1 6818
2 58368 1 6818
2 58369 1 6819
2 58370 1 6819
2 58371 1 6819
2 58372 1 6820
2 58373 1 6820
2 58374 1 6820
2 58375 1 6827
2 58376 1 6827
2 58377 1 6833
2 58378 1 6833
2 58379 1 6837
2 58380 1 6837
2 58381 1 6840
2 58382 1 6840
2 58383 1 6840
2 58384 1 6840
2 58385 1 6843
2 58386 1 6843
2 58387 1 6848
2 58388 1 6848
2 58389 1 6848
2 58390 1 6849
2 58391 1 6849
2 58392 1 6849
2 58393 1 6849
2 58394 1 6849
2 58395 1 6850
2 58396 1 6850
2 58397 1 6850
2 58398 1 6850
2 58399 1 6854
2 58400 1 6854
2 58401 1 6855
2 58402 1 6855
2 58403 1 6859
2 58404 1 6859
2 58405 1 6859
2 58406 1 6860
2 58407 1 6860
2 58408 1 6860
2 58409 1 6892
2 58410 1 6892
2 58411 1 6892
2 58412 1 6892
2 58413 1 6892
2 58414 1 6892
2 58415 1 6892
2 58416 1 6892
2 58417 1 6892
2 58418 1 6892
2 58419 1 6892
2 58420 1 6894
2 58421 1 6894
2 58422 1 6897
2 58423 1 6897
2 58424 1 6897
2 58425 1 6897
2 58426 1 6897
2 58427 1 6897
2 58428 1 6897
2 58429 1 6897
2 58430 1 6897
2 58431 1 6899
2 58432 1 6899
2 58433 1 6900
2 58434 1 6900
2 58435 1 6900
2 58436 1 6900
2 58437 1 6900
2 58438 1 6901
2 58439 1 6901
2 58440 1 6901
2 58441 1 6901
2 58442 1 6901
2 58443 1 6903
2 58444 1 6903
2 58445 1 6905
2 58446 1 6905
2 58447 1 6905
2 58448 1 6905
2 58449 1 6905
2 58450 1 6905
2 58451 1 6906
2 58452 1 6906
2 58453 1 6908
2 58454 1 6908
2 58455 1 6909
2 58456 1 6909
2 58457 1 6909
2 58458 1 6911
2 58459 1 6911
2 58460 1 6911
2 58461 1 6915
2 58462 1 6915
2 58463 1 6918
2 58464 1 6918
2 58465 1 6918
2 58466 1 6919
2 58467 1 6919
2 58468 1 6937
2 58469 1 6937
2 58470 1 6948
2 58471 1 6948
2 58472 1 6948
2 58473 1 6948
2 58474 1 6949
2 58475 1 6949
2 58476 1 6951
2 58477 1 6951
2 58478 1 6953
2 58479 1 6953
2 58480 1 6955
2 58481 1 6955
2 58482 1 6956
2 58483 1 6956
2 58484 1 6960
2 58485 1 6960
2 58486 1 6963
2 58487 1 6963
2 58488 1 6963
2 58489 1 6964
2 58490 1 6964
2 58491 1 6969
2 58492 1 6969
2 58493 1 6979
2 58494 1 6979
2 58495 1 6979
2 58496 1 6979
2 58497 1 6987
2 58498 1 6987
2 58499 1 6988
2 58500 1 6988
2 58501 1 6997
2 58502 1 6997
2 58503 1 6997
2 58504 1 6999
2 58505 1 6999
2 58506 1 6999
2 58507 1 6999
2 58508 1 7013
2 58509 1 7013
2 58510 1 7013
2 58511 1 7024
2 58512 1 7024
2 58513 1 7031
2 58514 1 7031
2 58515 1 7031
2 58516 1 7032
2 58517 1 7032
2 58518 1 7032
2 58519 1 7041
2 58520 1 7041
2 58521 1 7056
2 58522 1 7056
2 58523 1 7056
2 58524 1 7062
2 58525 1 7062
2 58526 1 7062
2 58527 1 7063
2 58528 1 7063
2 58529 1 7063
2 58530 1 7066
2 58531 1 7066
2 58532 1 7066
2 58533 1 7070
2 58534 1 7070
2 58535 1 7071
2 58536 1 7071
2 58537 1 7084
2 58538 1 7084
2 58539 1 7084
2 58540 1 7084
2 58541 1 7084
2 58542 1 7084
2 58543 1 7084
2 58544 1 7084
2 58545 1 7084
2 58546 1 7084
2 58547 1 7084
2 58548 1 7084
2 58549 1 7084
2 58550 1 7084
2 58551 1 7084
2 58552 1 7084
2 58553 1 7084
2 58554 1 7084
2 58555 1 7084
2 58556 1 7084
2 58557 1 7084
2 58558 1 7085
2 58559 1 7085
2 58560 1 7088
2 58561 1 7088
2 58562 1 7088
2 58563 1 7088
2 58564 1 7088
2 58565 1 7088
2 58566 1 7088
2 58567 1 7088
2 58568 1 7088
2 58569 1 7088
2 58570 1 7088
2 58571 1 7088
2 58572 1 7088
2 58573 1 7088
2 58574 1 7088
2 58575 1 7088
2 58576 1 7088
2 58577 1 7088
2 58578 1 7089
2 58579 1 7089
2 58580 1 7089
2 58581 1 7089
2 58582 1 7089
2 58583 1 7089
2 58584 1 7089
2 58585 1 7090
2 58586 1 7090
2 58587 1 7097
2 58588 1 7097
2 58589 1 7097
2 58590 1 7097
2 58591 1 7097
2 58592 1 7104
2 58593 1 7104
2 58594 1 7104
2 58595 1 7104
2 58596 1 7106
2 58597 1 7106
2 58598 1 7106
2 58599 1 7107
2 58600 1 7107
2 58601 1 7108
2 58602 1 7108
2 58603 1 7108
2 58604 1 7111
2 58605 1 7111
2 58606 1 7118
2 58607 1 7118
2 58608 1 7118
2 58609 1 7118
2 58610 1 7118
2 58611 1 7118
2 58612 1 7118
2 58613 1 7119
2 58614 1 7119
2 58615 1 7120
2 58616 1 7120
2 58617 1 7127
2 58618 1 7127
2 58619 1 7127
2 58620 1 7127
2 58621 1 7127
2 58622 1 7139
2 58623 1 7139
2 58624 1 7139
2 58625 1 7139
2 58626 1 7139
2 58627 1 7140
2 58628 1 7140
2 58629 1 7145
2 58630 1 7145
2 58631 1 7145
2 58632 1 7145
2 58633 1 7148
2 58634 1 7148
2 58635 1 7148
2 58636 1 7148
2 58637 1 7156
2 58638 1 7156
2 58639 1 7156
2 58640 1 7157
2 58641 1 7157
2 58642 1 7157
2 58643 1 7174
2 58644 1 7174
2 58645 1 7188
2 58646 1 7188
2 58647 1 7188
2 58648 1 7189
2 58649 1 7189
2 58650 1 7190
2 58651 1 7190
2 58652 1 7190
2 58653 1 7190
2 58654 1 7199
2 58655 1 7199
2 58656 1 7199
2 58657 1 7199
2 58658 1 7199
2 58659 1 7199
2 58660 1 7199
2 58661 1 7199
2 58662 1 7199
2 58663 1 7199
2 58664 1 7199
2 58665 1 7200
2 58666 1 7200
2 58667 1 7200
2 58668 1 7200
2 58669 1 7200
2 58670 1 7200
2 58671 1 7200
2 58672 1 7200
2 58673 1 7200
2 58674 1 7200
2 58675 1 7200
2 58676 1 7200
2 58677 1 7201
2 58678 1 7201
2 58679 1 7209
2 58680 1 7209
2 58681 1 7209
2 58682 1 7209
2 58683 1 7209
2 58684 1 7209
2 58685 1 7209
2 58686 1 7209
2 58687 1 7209
2 58688 1 7210
2 58689 1 7210
2 58690 1 7210
2 58691 1 7211
2 58692 1 7211
2 58693 1 7211
2 58694 1 7211
2 58695 1 7231
2 58696 1 7231
2 58697 1 7243
2 58698 1 7243
2 58699 1 7243
2 58700 1 7250
2 58701 1 7250
2 58702 1 7250
2 58703 1 7259
2 58704 1 7259
2 58705 1 7259
2 58706 1 7259
2 58707 1 7282
2 58708 1 7282
2 58709 1 7282
2 58710 1 7282
2 58711 1 7282
2 58712 1 7283
2 58713 1 7283
2 58714 1 7283
2 58715 1 7283
2 58716 1 7284
2 58717 1 7284
2 58718 1 7298
2 58719 1 7298
2 58720 1 7298
2 58721 1 7298
2 58722 1 7298
2 58723 1 7298
2 58724 1 7298
2 58725 1 7298
2 58726 1 7298
2 58727 1 7298
2 58728 1 7298
2 58729 1 7299
2 58730 1 7299
2 58731 1 7303
2 58732 1 7303
2 58733 1 7303
2 58734 1 7309
2 58735 1 7309
2 58736 1 7330
2 58737 1 7330
2 58738 1 7331
2 58739 1 7331
2 58740 1 7338
2 58741 1 7338
2 58742 1 7341
2 58743 1 7341
2 58744 1 7341
2 58745 1 7341
2 58746 1 7341
2 58747 1 7341
2 58748 1 7341
2 58749 1 7341
2 58750 1 7342
2 58751 1 7342
2 58752 1 7343
2 58753 1 7343
2 58754 1 7343
2 58755 1 7350
2 58756 1 7350
2 58757 1 7350
2 58758 1 7350
2 58759 1 7351
2 58760 1 7351
2 58761 1 7351
2 58762 1 7352
2 58763 1 7352
2 58764 1 7352
2 58765 1 7352
2 58766 1 7353
2 58767 1 7353
2 58768 1 7360
2 58769 1 7360
2 58770 1 7360
2 58771 1 7360
2 58772 1 7360
2 58773 1 7360
2 58774 1 7360
2 58775 1 7361
2 58776 1 7361
2 58777 1 7361
2 58778 1 7388
2 58779 1 7388
2 58780 1 7389
2 58781 1 7389
2 58782 1 7389
2 58783 1 7389
2 58784 1 7389
2 58785 1 7389
2 58786 1 7389
2 58787 1 7396
2 58788 1 7396
2 58789 1 7396
2 58790 1 7396
2 58791 1 7396
2 58792 1 7396
2 58793 1 7396
2 58794 1 7396
2 58795 1 7397
2 58796 1 7397
2 58797 1 7397
2 58798 1 7397
2 58799 1 7397
2 58800 1 7397
2 58801 1 7406
2 58802 1 7406
2 58803 1 7409
2 58804 1 7409
2 58805 1 7409
2 58806 1 7422
2 58807 1 7422
2 58808 1 7422
2 58809 1 7425
2 58810 1 7425
2 58811 1 7425
2 58812 1 7425
2 58813 1 7447
2 58814 1 7447
2 58815 1 7447
2 58816 1 7447
2 58817 1 7448
2 58818 1 7448
2 58819 1 7448
2 58820 1 7449
2 58821 1 7449
2 58822 1 7450
2 58823 1 7450
2 58824 1 7450
2 58825 1 7459
2 58826 1 7459
2 58827 1 7459
2 58828 1 7459
2 58829 1 7460
2 58830 1 7460
2 58831 1 7460
2 58832 1 7460
2 58833 1 7463
2 58834 1 7463
2 58835 1 7475
2 58836 1 7475
2 58837 1 7475
2 58838 1 7484
2 58839 1 7484
2 58840 1 7485
2 58841 1 7485
2 58842 1 7486
2 58843 1 7486
2 58844 1 7497
2 58845 1 7497
2 58846 1 7498
2 58847 1 7498
2 58848 1 7501
2 58849 1 7501
2 58850 1 7502
2 58851 1 7502
2 58852 1 7502
2 58853 1 7502
2 58854 1 7503
2 58855 1 7503
2 58856 1 7514
2 58857 1 7514
2 58858 1 7514
2 58859 1 7514
2 58860 1 7514
2 58861 1 7514
2 58862 1 7514
2 58863 1 7514
2 58864 1 7531
2 58865 1 7531
2 58866 1 7531
2 58867 1 7531
2 58868 1 7531
2 58869 1 7532
2 58870 1 7532
2 58871 1 7532
2 58872 1 7532
2 58873 1 7536
2 58874 1 7536
2 58875 1 7563
2 58876 1 7563
2 58877 1 7571
2 58878 1 7571
2 58879 1 7571
2 58880 1 7571
2 58881 1 7571
2 58882 1 7573
2 58883 1 7573
2 58884 1 7574
2 58885 1 7574
2 58886 1 7574
2 58887 1 7574
2 58888 1 7574
2 58889 1 7574
2 58890 1 7574
2 58891 1 7574
2 58892 1 7574
2 58893 1 7574
2 58894 1 7574
2 58895 1 7574
2 58896 1 7574
2 58897 1 7574
2 58898 1 7574
2 58899 1 7574
2 58900 1 7574
2 58901 1 7574
2 58902 1 7574
2 58903 1 7574
2 58904 1 7575
2 58905 1 7575
2 58906 1 7575
2 58907 1 7575
2 58908 1 7577
2 58909 1 7577
2 58910 1 7577
2 58911 1 7580
2 58912 1 7580
2 58913 1 7580
2 58914 1 7580
2 58915 1 7580
2 58916 1 7580
2 58917 1 7580
2 58918 1 7580
2 58919 1 7580
2 58920 1 7590
2 58921 1 7590
2 58922 1 7590
2 58923 1 7597
2 58924 1 7597
2 58925 1 7597
2 58926 1 7597
2 58927 1 7597
2 58928 1 7597
2 58929 1 7598
2 58930 1 7598
2 58931 1 7598
2 58932 1 7598
2 58933 1 7598
2 58934 1 7605
2 58935 1 7605
2 58936 1 7605
2 58937 1 7605
2 58938 1 7605
2 58939 1 7606
2 58940 1 7606
2 58941 1 7606
2 58942 1 7606
2 58943 1 7606
2 58944 1 7606
2 58945 1 7613
2 58946 1 7613
2 58947 1 7614
2 58948 1 7614
2 58949 1 7614
2 58950 1 7626
2 58951 1 7626
2 58952 1 7633
2 58953 1 7633
2 58954 1 7639
2 58955 1 7639
2 58956 1 7639
2 58957 1 7646
2 58958 1 7646
2 58959 1 7646
2 58960 1 7646
2 58961 1 7646
2 58962 1 7646
2 58963 1 7657
2 58964 1 7657
2 58965 1 7657
2 58966 1 7657
2 58967 1 7658
2 58968 1 7658
2 58969 1 7658
2 58970 1 7659
2 58971 1 7659
2 58972 1 7661
2 58973 1 7661
2 58974 1 7661
2 58975 1 7684
2 58976 1 7684
2 58977 1 7685
2 58978 1 7685
2 58979 1 7685
2 58980 1 7685
2 58981 1 7686
2 58982 1 7686
2 58983 1 7686
2 58984 1 7686
2 58985 1 7686
2 58986 1 7686
2 58987 1 7686
2 58988 1 7686
2 58989 1 7686
2 58990 1 7686
2 58991 1 7686
2 58992 1 7690
2 58993 1 7690
2 58994 1 7697
2 58995 1 7697
2 58996 1 7698
2 58997 1 7698
2 58998 1 7698
2 58999 1 7698
2 59000 1 7698
2 59001 1 7698
2 59002 1 7698
2 59003 1 7698
2 59004 1 7698
2 59005 1 7698
2 59006 1 7698
2 59007 1 7698
2 59008 1 7698
2 59009 1 7717
2 59010 1 7717
2 59011 1 7720
2 59012 1 7720
2 59013 1 7720
2 59014 1 7720
2 59015 1 7720
2 59016 1 7720
2 59017 1 7720
2 59018 1 7724
2 59019 1 7724
2 59020 1 7724
2 59021 1 7724
2 59022 1 7728
2 59023 1 7728
2 59024 1 7728
2 59025 1 7728
2 59026 1 7729
2 59027 1 7729
2 59028 1 7730
2 59029 1 7730
2 59030 1 7730
2 59031 1 7730
2 59032 1 7732
2 59033 1 7732
2 59034 1 7732
2 59035 1 7732
2 59036 1 7732
2 59037 1 7740
2 59038 1 7740
2 59039 1 7741
2 59040 1 7741
2 59041 1 7741
2 59042 1 7741
2 59043 1 7741
2 59044 1 7741
2 59045 1 7741
2 59046 1 7741
2 59047 1 7741
2 59048 1 7741
2 59049 1 7741
2 59050 1 7741
2 59051 1 7741
2 59052 1 7741
2 59053 1 7741
2 59054 1 7741
2 59055 1 7741
2 59056 1 7741
2 59057 1 7741
2 59058 1 7741
2 59059 1 7741
2 59060 1 7742
2 59061 1 7742
2 59062 1 7743
2 59063 1 7743
2 59064 1 7743
2 59065 1 7743
2 59066 1 7743
2 59067 1 7743
2 59068 1 7743
2 59069 1 7744
2 59070 1 7744
2 59071 1 7744
2 59072 1 7753
2 59073 1 7753
2 59074 1 7753
2 59075 1 7755
2 59076 1 7755
2 59077 1 7755
2 59078 1 7756
2 59079 1 7756
2 59080 1 7756
2 59081 1 7756
2 59082 1 7756
2 59083 1 7770
2 59084 1 7770
2 59085 1 7770
2 59086 1 7770
2 59087 1 7771
2 59088 1 7771
2 59089 1 7771
2 59090 1 7771
2 59091 1 7771
2 59092 1 7771
2 59093 1 7771
2 59094 1 7771
2 59095 1 7772
2 59096 1 7772
2 59097 1 7772
2 59098 1 7775
2 59099 1 7775
2 59100 1 7775
2 59101 1 7775
2 59102 1 7775
2 59103 1 7778
2 59104 1 7778
2 59105 1 7779
2 59106 1 7779
2 59107 1 7783
2 59108 1 7783
2 59109 1 7789
2 59110 1 7789
2 59111 1 7814
2 59112 1 7814
2 59113 1 7844
2 59114 1 7844
2 59115 1 7844
2 59116 1 7844
2 59117 1 7844
2 59118 1 7844
2 59119 1 7844
2 59120 1 7844
2 59121 1 7844
2 59122 1 7844
2 59123 1 7844
2 59124 1 7845
2 59125 1 7845
2 59126 1 7845
2 59127 1 7846
2 59128 1 7846
2 59129 1 7847
2 59130 1 7847
2 59131 1 7848
2 59132 1 7848
2 59133 1 7851
2 59134 1 7851
2 59135 1 7851
2 59136 1 7851
2 59137 1 7851
2 59138 1 7851
2 59139 1 7851
2 59140 1 7851
2 59141 1 7851
2 59142 1 7851
2 59143 1 7851
2 59144 1 7851
2 59145 1 7851
2 59146 1 7851
2 59147 1 7851
2 59148 1 7851
2 59149 1 7852
2 59150 1 7852
2 59151 1 7852
2 59152 1 7852
2 59153 1 7852
2 59154 1 7852
2 59155 1 7852
2 59156 1 7853
2 59157 1 7853
2 59158 1 7854
2 59159 1 7854
2 59160 1 7854
2 59161 1 7859
2 59162 1 7859
2 59163 1 7859
2 59164 1 7884
2 59165 1 7884
2 59166 1 7891
2 59167 1 7891
2 59168 1 7901
2 59169 1 7901
2 59170 1 7901
2 59171 1 7907
2 59172 1 7907
2 59173 1 7926
2 59174 1 7926
2 59175 1 7934
2 59176 1 7934
2 59177 1 7934
2 59178 1 7934
2 59179 1 7934
2 59180 1 7934
2 59181 1 7934
2 59182 1 7935
2 59183 1 7935
2 59184 1 7935
2 59185 1 7935
2 59186 1 7935
2 59187 1 7935
2 59188 1 7935
2 59189 1 7946
2 59190 1 7946
2 59191 1 7947
2 59192 1 7947
2 59193 1 7947
2 59194 1 7950
2 59195 1 7950
2 59196 1 7950
2 59197 1 7950
2 59198 1 7953
2 59199 1 7953
2 59200 1 7953
2 59201 1 7970
2 59202 1 7970
2 59203 1 7970
2 59204 1 7970
2 59205 1 7970
2 59206 1 7970
2 59207 1 7970
2 59208 1 7970
2 59209 1 7971
2 59210 1 7971
2 59211 1 7971
2 59212 1 7974
2 59213 1 7974
2 59214 1 7982
2 59215 1 7982
2 59216 1 7982
2 59217 1 7982
2 59218 1 7982
2 59219 1 7982
2 59220 1 7982
2 59221 1 7982
2 59222 1 7983
2 59223 1 7983
2 59224 1 7983
2 59225 1 7983
2 59226 1 7985
2 59227 1 7985
2 59228 1 7988
2 59229 1 7988
2 59230 1 7991
2 59231 1 7991
2 59232 1 7992
2 59233 1 7992
2 59234 1 7993
2 59235 1 7993
2 59236 1 8014
2 59237 1 8014
2 59238 1 8015
2 59239 1 8015
2 59240 1 8015
2 59241 1 8015
2 59242 1 8016
2 59243 1 8016
2 59244 1 8016
2 59245 1 8016
2 59246 1 8020
2 59247 1 8020
2 59248 1 8031
2 59249 1 8031
2 59250 1 8031
2 59251 1 8031
2 59252 1 8049
2 59253 1 8049
2 59254 1 8049
2 59255 1 8049
2 59256 1 8049
2 59257 1 8049
2 59258 1 8049
2 59259 1 8056
2 59260 1 8056
2 59261 1 8056
2 59262 1 8056
2 59263 1 8057
2 59264 1 8057
2 59265 1 8057
2 59266 1 8058
2 59267 1 8058
2 59268 1 8097
2 59269 1 8097
2 59270 1 8097
2 59271 1 8097
2 59272 1 8097
2 59273 1 8097
2 59274 1 8097
2 59275 1 8097
2 59276 1 8098
2 59277 1 8098
2 59278 1 8101
2 59279 1 8101
2 59280 1 8101
2 59281 1 8108
2 59282 1 8108
2 59283 1 8109
2 59284 1 8109
2 59285 1 8109
2 59286 1 8109
2 59287 1 8109
2 59288 1 8109
2 59289 1 8117
2 59290 1 8117
2 59291 1 8117
2 59292 1 8117
2 59293 1 8117
2 59294 1 8117
2 59295 1 8117
2 59296 1 8117
2 59297 1 8125
2 59298 1 8125
2 59299 1 8125
2 59300 1 8125
2 59301 1 8125
2 59302 1 8125
2 59303 1 8125
2 59304 1 8125
2 59305 1 8127
2 59306 1 8127
2 59307 1 8127
2 59308 1 8127
2 59309 1 8127
2 59310 1 8127
2 59311 1 8129
2 59312 1 8129
2 59313 1 8129
2 59314 1 8129
2 59315 1 8129
2 59316 1 8130
2 59317 1 8130
2 59318 1 8131
2 59319 1 8131
2 59320 1 8138
2 59321 1 8138
2 59322 1 8138
2 59323 1 8138
2 59324 1 8138
2 59325 1 8139
2 59326 1 8139
2 59327 1 8139
2 59328 1 8139
2 59329 1 8139
2 59330 1 8139
2 59331 1 8142
2 59332 1 8142
2 59333 1 8142
2 59334 1 8142
2 59335 1 8142
2 59336 1 8142
2 59337 1 8142
2 59338 1 8144
2 59339 1 8144
2 59340 1 8152
2 59341 1 8152
2 59342 1 8152
2 59343 1 8152
2 59344 1 8152
2 59345 1 8152
2 59346 1 8152
2 59347 1 8153
2 59348 1 8153
2 59349 1 8153
2 59350 1 8153
2 59351 1 8153
2 59352 1 8154
2 59353 1 8154
2 59354 1 8164
2 59355 1 8164
2 59356 1 8164
2 59357 1 8164
2 59358 1 8165
2 59359 1 8165
2 59360 1 8165
2 59361 1 8165
2 59362 1 8165
2 59363 1 8165
2 59364 1 8165
2 59365 1 8165
2 59366 1 8165
2 59367 1 8165
2 59368 1 8169
2 59369 1 8169
2 59370 1 8169
2 59371 1 8169
2 59372 1 8194
2 59373 1 8194
2 59374 1 8194
2 59375 1 8194
2 59376 1 8195
2 59377 1 8195
2 59378 1 8195
2 59379 1 8195
2 59380 1 8196
2 59381 1 8196
2 59382 1 8197
2 59383 1 8197
2 59384 1 8206
2 59385 1 8206
2 59386 1 8206
2 59387 1 8206
2 59388 1 8206
2 59389 1 8206
2 59390 1 8206
2 59391 1 8207
2 59392 1 8207
2 59393 1 8207
2 59394 1 8207
2 59395 1 8207
2 59396 1 8207
2 59397 1 8207
2 59398 1 8207
2 59399 1 8207
2 59400 1 8207
2 59401 1 8209
2 59402 1 8209
2 59403 1 8226
2 59404 1 8226
2 59405 1 8226
2 59406 1 8227
2 59407 1 8227
2 59408 1 8227
2 59409 1 8242
2 59410 1 8242
2 59411 1 8242
2 59412 1 8242
2 59413 1 8245
2 59414 1 8245
2 59415 1 8259
2 59416 1 8259
2 59417 1 8259
2 59418 1 8260
2 59419 1 8260
2 59420 1 8260
2 59421 1 8260
2 59422 1 8260
2 59423 1 8260
2 59424 1 8260
2 59425 1 8260
2 59426 1 8260
2 59427 1 8260
2 59428 1 8260
2 59429 1 8260
2 59430 1 8260
2 59431 1 8260
2 59432 1 8261
2 59433 1 8261
2 59434 1 8270
2 59435 1 8270
2 59436 1 8270
2 59437 1 8271
2 59438 1 8271
2 59439 1 8277
2 59440 1 8277
2 59441 1 8277
2 59442 1 8277
2 59443 1 8277
2 59444 1 8277
2 59445 1 8277
2 59446 1 8277
2 59447 1 8277
2 59448 1 8277
2 59449 1 8277
2 59450 1 8277
2 59451 1 8277
2 59452 1 8277
2 59453 1 8277
2 59454 1 8277
2 59455 1 8277
2 59456 1 8277
2 59457 1 8277
2 59458 1 8277
2 59459 1 8277
2 59460 1 8277
2 59461 1 8277
2 59462 1 8277
2 59463 1 8277
2 59464 1 8277
2 59465 1 8277
2 59466 1 8277
2 59467 1 8277
2 59468 1 8277
2 59469 1 8277
2 59470 1 8277
2 59471 1 8277
2 59472 1 8277
2 59473 1 8277
2 59474 1 8277
2 59475 1 8277
2 59476 1 8277
2 59477 1 8277
2 59478 1 8277
2 59479 1 8277
2 59480 1 8277
2 59481 1 8277
2 59482 1 8277
2 59483 1 8277
2 59484 1 8277
2 59485 1 8277
2 59486 1 8277
2 59487 1 8277
2 59488 1 8277
2 59489 1 8277
2 59490 1 8277
2 59491 1 8277
2 59492 1 8277
2 59493 1 8277
2 59494 1 8278
2 59495 1 8278
2 59496 1 8278
2 59497 1 8278
2 59498 1 8279
2 59499 1 8279
2 59500 1 8289
2 59501 1 8289
2 59502 1 8290
2 59503 1 8290
2 59504 1 8290
2 59505 1 8290
2 59506 1 8290
2 59507 1 8290
2 59508 1 8290
2 59509 1 8290
2 59510 1 8290
2 59511 1 8290
2 59512 1 8290
2 59513 1 8290
2 59514 1 8295
2 59515 1 8295
2 59516 1 8295
2 59517 1 8295
2 59518 1 8295
2 59519 1 8295
2 59520 1 8295
2 59521 1 8296
2 59522 1 8296
2 59523 1 8296
2 59524 1 8296
2 59525 1 8296
2 59526 1 8313
2 59527 1 8313
2 59528 1 8313
2 59529 1 8313
2 59530 1 8313
2 59531 1 8313
2 59532 1 8313
2 59533 1 8313
2 59534 1 8313
2 59535 1 8313
2 59536 1 8313
2 59537 1 8313
2 59538 1 8313
2 59539 1 8313
2 59540 1 8313
2 59541 1 8313
2 59542 1 8313
2 59543 1 8313
2 59544 1 8313
2 59545 1 8313
2 59546 1 8313
2 59547 1 8313
2 59548 1 8313
2 59549 1 8317
2 59550 1 8317
2 59551 1 8318
2 59552 1 8318
2 59553 1 8319
2 59554 1 8319
2 59555 1 8319
2 59556 1 8319
2 59557 1 8321
2 59558 1 8321
2 59559 1 8321
2 59560 1 8322
2 59561 1 8322
2 59562 1 8329
2 59563 1 8329
2 59564 1 8329
2 59565 1 8336
2 59566 1 8336
2 59567 1 8336
2 59568 1 8345
2 59569 1 8345
2 59570 1 8345
2 59571 1 8345
2 59572 1 8345
2 59573 1 8345
2 59574 1 8346
2 59575 1 8346
2 59576 1 8348
2 59577 1 8348
2 59578 1 8349
2 59579 1 8349
2 59580 1 8352
2 59581 1 8352
2 59582 1 8354
2 59583 1 8354
2 59584 1 8354
2 59585 1 8362
2 59586 1 8362
2 59587 1 8390
2 59588 1 8390
2 59589 1 8394
2 59590 1 8394
2 59591 1 8397
2 59592 1 8397
2 59593 1 8400
2 59594 1 8400
2 59595 1 8400
2 59596 1 8400
2 59597 1 8400
2 59598 1 8401
2 59599 1 8401
2 59600 1 8402
2 59601 1 8402
2 59602 1 8403
2 59603 1 8403
2 59604 1 8412
2 59605 1 8412
2 59606 1 8412
2 59607 1 8412
2 59608 1 8412
2 59609 1 8412
2 59610 1 8412
2 59611 1 8412
2 59612 1 8415
2 59613 1 8415
2 59614 1 8415
2 59615 1 8416
2 59616 1 8416
2 59617 1 8429
2 59618 1 8429
2 59619 1 8429
2 59620 1 8429
2 59621 1 8429
2 59622 1 8429
2 59623 1 8429
2 59624 1 8429
2 59625 1 8429
2 59626 1 8451
2 59627 1 8451
2 59628 1 8457
2 59629 1 8457
2 59630 1 8457
2 59631 1 8457
2 59632 1 8457
2 59633 1 8457
2 59634 1 8457
2 59635 1 8457
2 59636 1 8458
2 59637 1 8458
2 59638 1 8458
2 59639 1 8467
2 59640 1 8467
2 59641 1 8467
2 59642 1 8467
2 59643 1 8469
2 59644 1 8469
2 59645 1 8469
2 59646 1 8480
2 59647 1 8480
2 59648 1 8480
2 59649 1 8480
2 59650 1 8480
2 59651 1 8480
2 59652 1 8482
2 59653 1 8482
2 59654 1 8492
2 59655 1 8492
2 59656 1 8492
2 59657 1 8492
2 59658 1 8492
2 59659 1 8492
2 59660 1 8492
2 59661 1 8492
2 59662 1 8492
2 59663 1 8492
2 59664 1 8492
2 59665 1 8493
2 59666 1 8493
2 59667 1 8493
2 59668 1 8493
2 59669 1 8494
2 59670 1 8494
2 59671 1 8494
2 59672 1 8494
2 59673 1 8495
2 59674 1 8495
2 59675 1 8506
2 59676 1 8506
2 59677 1 8511
2 59678 1 8511
2 59679 1 8511
2 59680 1 8511
2 59681 1 8511
2 59682 1 8511
2 59683 1 8511
2 59684 1 8511
2 59685 1 8511
2 59686 1 8511
2 59687 1 8511
2 59688 1 8511
2 59689 1 8511
2 59690 1 8511
2 59691 1 8511
2 59692 1 8511
2 59693 1 8511
2 59694 1 8511
2 59695 1 8511
2 59696 1 8511
2 59697 1 8511
2 59698 1 8511
2 59699 1 8511
2 59700 1 8511
2 59701 1 8511
2 59702 1 8511
2 59703 1 8511
2 59704 1 8511
2 59705 1 8511
2 59706 1 8511
2 59707 1 8511
2 59708 1 8511
2 59709 1 8511
2 59710 1 8511
2 59711 1 8511
2 59712 1 8511
2 59713 1 8511
2 59714 1 8511
2 59715 1 8511
2 59716 1 8511
2 59717 1 8511
2 59718 1 8511
2 59719 1 8511
2 59720 1 8511
2 59721 1 8512
2 59722 1 8512
2 59723 1 8512
2 59724 1 8525
2 59725 1 8525
2 59726 1 8525
2 59727 1 8525
2 59728 1 8525
2 59729 1 8525
2 59730 1 8525
2 59731 1 8535
2 59732 1 8535
2 59733 1 8535
2 59734 1 8535
2 59735 1 8536
2 59736 1 8536
2 59737 1 8543
2 59738 1 8543
2 59739 1 8543
2 59740 1 8543
2 59741 1 8543
2 59742 1 8543
2 59743 1 8543
2 59744 1 8543
2 59745 1 8558
2 59746 1 8558
2 59747 1 8558
2 59748 1 8558
2 59749 1 8558
2 59750 1 8558
2 59751 1 8558
2 59752 1 8558
2 59753 1 8559
2 59754 1 8559
2 59755 1 8559
2 59756 1 8570
2 59757 1 8570
2 59758 1 8578
2 59759 1 8578
2 59760 1 8579
2 59761 1 8579
2 59762 1 8599
2 59763 1 8599
2 59764 1 8599
2 59765 1 8599
2 59766 1 8615
2 59767 1 8615
2 59768 1 8620
2 59769 1 8620
2 59770 1 8623
2 59771 1 8623
2 59772 1 8628
2 59773 1 8628
2 59774 1 8630
2 59775 1 8630
2 59776 1 8630
2 59777 1 8630
2 59778 1 8630
2 59779 1 8630
2 59780 1 8647
2 59781 1 8647
2 59782 1 8647
2 59783 1 8647
2 59784 1 8647
2 59785 1 8647
2 59786 1 8650
2 59787 1 8650
2 59788 1 8651
2 59789 1 8651
2 59790 1 8651
2 59791 1 8654
2 59792 1 8654
2 59793 1 8665
2 59794 1 8665
2 59795 1 8668
2 59796 1 8668
2 59797 1 8676
2 59798 1 8676
2 59799 1 8676
2 59800 1 8677
2 59801 1 8677
2 59802 1 8677
2 59803 1 8678
2 59804 1 8678
2 59805 1 8682
2 59806 1 8682
2 59807 1 8692
2 59808 1 8692
2 59809 1 8720
2 59810 1 8720
2 59811 1 8720
2 59812 1 8723
2 59813 1 8723
2 59814 1 8729
2 59815 1 8729
2 59816 1 8734
2 59817 1 8734
2 59818 1 8734
2 59819 1 8734
2 59820 1 8734
2 59821 1 8734
2 59822 1 8741
2 59823 1 8741
2 59824 1 8741
2 59825 1 8741
2 59826 1 8742
2 59827 1 8742
2 59828 1 8744
2 59829 1 8744
2 59830 1 8751
2 59831 1 8751
2 59832 1 8752
2 59833 1 8752
2 59834 1 8760
2 59835 1 8760
2 59836 1 8787
2 59837 1 8787
2 59838 1 8802
2 59839 1 8802
2 59840 1 8806
2 59841 1 8806
2 59842 1 8807
2 59843 1 8807
2 59844 1 8821
2 59845 1 8821
2 59846 1 8822
2 59847 1 8822
2 59848 1 8822
2 59849 1 8822
2 59850 1 8822
2 59851 1 8843
2 59852 1 8843
2 59853 1 8843
2 59854 1 8843
2 59855 1 8847
2 59856 1 8847
2 59857 1 8847
2 59858 1 8847
2 59859 1 8848
2 59860 1 8848
2 59861 1 8862
2 59862 1 8862
2 59863 1 8865
2 59864 1 8865
2 59865 1 8865
2 59866 1 8866
2 59867 1 8866
2 59868 1 8866
2 59869 1 8866
2 59870 1 8866
2 59871 1 8867
2 59872 1 8867
2 59873 1 8867
2 59874 1 8867
2 59875 1 8882
2 59876 1 8882
2 59877 1 8883
2 59878 1 8883
2 59879 1 8901
2 59880 1 8901
2 59881 1 8901
2 59882 1 8913
2 59883 1 8913
2 59884 1 8913
2 59885 1 8913
2 59886 1 8915
2 59887 1 8915
2 59888 1 8919
2 59889 1 8919
2 59890 1 8919
2 59891 1 8919
2 59892 1 8935
2 59893 1 8935
2 59894 1 8936
2 59895 1 8936
2 59896 1 8936
2 59897 1 8957
2 59898 1 8957
2 59899 1 8973
2 59900 1 8973
2 59901 1 8981
2 59902 1 8981
2 59903 1 8992
2 59904 1 8992
2 59905 1 8992
2 59906 1 8993
2 59907 1 8993
2 59908 1 9019
2 59909 1 9019
2 59910 1 9019
2 59911 1 9019
2 59912 1 9019
2 59913 1 9019
2 59914 1 9019
2 59915 1 9020
2 59916 1 9020
2 59917 1 9028
2 59918 1 9028
2 59919 1 9028
2 59920 1 9028
2 59921 1 9031
2 59922 1 9031
2 59923 1 9032
2 59924 1 9032
2 59925 1 9032
2 59926 1 9061
2 59927 1 9061
2 59928 1 9061
2 59929 1 9061
2 59930 1 9061
2 59931 1 9061
2 59932 1 9061
2 59933 1 9061
2 59934 1 9062
2 59935 1 9062
2 59936 1 9062
2 59937 1 9062
2 59938 1 9062
2 59939 1 9062
2 59940 1 9063
2 59941 1 9063
2 59942 1 9077
2 59943 1 9077
2 59944 1 9077
2 59945 1 9080
2 59946 1 9080
2 59947 1 9090
2 59948 1 9090
2 59949 1 9090
2 59950 1 9090
2 59951 1 9090
2 59952 1 9090
2 59953 1 9090
2 59954 1 9090
2 59955 1 9090
2 59956 1 9090
2 59957 1 9090
2 59958 1 9090
2 59959 1 9090
2 59960 1 9090
2 59961 1 9090
2 59962 1 9090
2 59963 1 9090
2 59964 1 9090
2 59965 1 9090
2 59966 1 9090
2 59967 1 9091
2 59968 1 9091
2 59969 1 9091
2 59970 1 9091
2 59971 1 9091
2 59972 1 9091
2 59973 1 9092
2 59974 1 9092
2 59975 1 9092
2 59976 1 9092
2 59977 1 9092
2 59978 1 9092
2 59979 1 9093
2 59980 1 9093
2 59981 1 9093
2 59982 1 9093
2 59983 1 9093
2 59984 1 9099
2 59985 1 9099
2 59986 1 9112
2 59987 1 9112
2 59988 1 9112
2 59989 1 9112
2 59990 1 9112
2 59991 1 9112
2 59992 1 9112
2 59993 1 9112
2 59994 1 9112
2 59995 1 9112
2 59996 1 9113
2 59997 1 9113
2 59998 1 9113
2 59999 1 9113
2 60000 1 9114
2 60001 1 9114
2 60002 1 9118
2 60003 1 9118
2 60004 1 9118
2 60005 1 9118
2 60006 1 9118
2 60007 1 9124
2 60008 1 9124
2 60009 1 9124
2 60010 1 9137
2 60011 1 9137
2 60012 1 9137
2 60013 1 9137
2 60014 1 9137
2 60015 1 9138
2 60016 1 9138
2 60017 1 9138
2 60018 1 9146
2 60019 1 9146
2 60020 1 9147
2 60021 1 9147
2 60022 1 9147
2 60023 1 9147
2 60024 1 9147
2 60025 1 9147
2 60026 1 9148
2 60027 1 9148
2 60028 1 9148
2 60029 1 9148
2 60030 1 9175
2 60031 1 9175
2 60032 1 9175
2 60033 1 9175
2 60034 1 9176
2 60035 1 9176
2 60036 1 9177
2 60037 1 9177
2 60038 1 9178
2 60039 1 9178
2 60040 1 9178
2 60041 1 9178
2 60042 1 9189
2 60043 1 9189
2 60044 1 9189
2 60045 1 9189
2 60046 1 9192
2 60047 1 9192
2 60048 1 9192
2 60049 1 9192
2 60050 1 9192
2 60051 1 9192
2 60052 1 9192
2 60053 1 9205
2 60054 1 9205
2 60055 1 9205
2 60056 1 9210
2 60057 1 9210
2 60058 1 9210
2 60059 1 9210
2 60060 1 9210
2 60061 1 9226
2 60062 1 9226
2 60063 1 9227
2 60064 1 9227
2 60065 1 9228
2 60066 1 9228
2 60067 1 9236
2 60068 1 9236
2 60069 1 9236
2 60070 1 9236
2 60071 1 9236
2 60072 1 9236
2 60073 1 9236
2 60074 1 9236
2 60075 1 9236
2 60076 1 9247
2 60077 1 9247
2 60078 1 9247
2 60079 1 9248
2 60080 1 9248
2 60081 1 9248
2 60082 1 9251
2 60083 1 9251
2 60084 1 9251
2 60085 1 9251
2 60086 1 9251
2 60087 1 9251
2 60088 1 9251
2 60089 1 9251
2 60090 1 9251
2 60091 1 9251
2 60092 1 9253
2 60093 1 9253
2 60094 1 9255
2 60095 1 9255
2 60096 1 9255
2 60097 1 9256
2 60098 1 9256
2 60099 1 9256
2 60100 1 9256
2 60101 1 9265
2 60102 1 9265
2 60103 1 9265
2 60104 1 9265
2 60105 1 9265
2 60106 1 9265
2 60107 1 9266
2 60108 1 9266
2 60109 1 9266
2 60110 1 9266
2 60111 1 9266
2 60112 1 9266
2 60113 1 9266
2 60114 1 9266
2 60115 1 9266
2 60116 1 9266
2 60117 1 9266
2 60118 1 9266
2 60119 1 9266
2 60120 1 9266
2 60121 1 9267
2 60122 1 9267
2 60123 1 9274
2 60124 1 9274
2 60125 1 9275
2 60126 1 9275
2 60127 1 9275
2 60128 1 9275
2 60129 1 9275
2 60130 1 9276
2 60131 1 9276
2 60132 1 9284
2 60133 1 9284
2 60134 1 9284
2 60135 1 9284
2 60136 1 9284
2 60137 1 9284
2 60138 1 9285
2 60139 1 9285
2 60140 1 9285
2 60141 1 9285
2 60142 1 9285
2 60143 1 9285
2 60144 1 9298
2 60145 1 9298
2 60146 1 9298
2 60147 1 9298
2 60148 1 9298
2 60149 1 9298
2 60150 1 9298
2 60151 1 9299
2 60152 1 9299
2 60153 1 9299
2 60154 1 9300
2 60155 1 9300
2 60156 1 9300
2 60157 1 9300
2 60158 1 9301
2 60159 1 9301
2 60160 1 9308
2 60161 1 9308
2 60162 1 9315
2 60163 1 9315
2 60164 1 9315
2 60165 1 9315
2 60166 1 9315
2 60167 1 9315
2 60168 1 9315
2 60169 1 9315
2 60170 1 9315
2 60171 1 9315
2 60172 1 9316
2 60173 1 9316
2 60174 1 9316
2 60175 1 9316
2 60176 1 9316
2 60177 1 9316
2 60178 1 9316
2 60179 1 9318
2 60180 1 9318
2 60181 1 9318
2 60182 1 9323
2 60183 1 9323
2 60184 1 9323
2 60185 1 9323
2 60186 1 9323
2 60187 1 9323
2 60188 1 9323
2 60189 1 9324
2 60190 1 9324
2 60191 1 9355
2 60192 1 9355
2 60193 1 9355
2 60194 1 9355
2 60195 1 9355
2 60196 1 9355
2 60197 1 9355
2 60198 1 9355
2 60199 1 9357
2 60200 1 9357
2 60201 1 9357
2 60202 1 9359
2 60203 1 9359
2 60204 1 9360
2 60205 1 9360
2 60206 1 9361
2 60207 1 9361
2 60208 1 9361
2 60209 1 9361
2 60210 1 9361
2 60211 1 9361
2 60212 1 9361
2 60213 1 9361
2 60214 1 9369
2 60215 1 9369
2 60216 1 9378
2 60217 1 9378
2 60218 1 9381
2 60219 1 9381
2 60220 1 9381
2 60221 1 9381
2 60222 1 9381
2 60223 1 9381
2 60224 1 9381
2 60225 1 9381
2 60226 1 9381
2 60227 1 9381
2 60228 1 9383
2 60229 1 9383
2 60230 1 9383
2 60231 1 9383
2 60232 1 9386
2 60233 1 9386
2 60234 1 9386
2 60235 1 9386
2 60236 1 9387
2 60237 1 9387
2 60238 1 9387
2 60239 1 9387
2 60240 1 9387
2 60241 1 9387
2 60242 1 9387
2 60243 1 9387
2 60244 1 9387
2 60245 1 9406
2 60246 1 9406
2 60247 1 9406
2 60248 1 9406
2 60249 1 9420
2 60250 1 9420
2 60251 1 9438
2 60252 1 9438
2 60253 1 9438
2 60254 1 9438
2 60255 1 9438
2 60256 1 9438
2 60257 1 9438
2 60258 1 9438
2 60259 1 9438
2 60260 1 9438
2 60261 1 9438
2 60262 1 9438
2 60263 1 9438
2 60264 1 9438
2 60265 1 9438
2 60266 1 9438
2 60267 1 9438
2 60268 1 9438
2 60269 1 9438
2 60270 1 9438
2 60271 1 9438
2 60272 1 9438
2 60273 1 9438
2 60274 1 9438
2 60275 1 9438
2 60276 1 9438
2 60277 1 9438
2 60278 1 9438
2 60279 1 9438
2 60280 1 9438
2 60281 1 9438
2 60282 1 9438
2 60283 1 9438
2 60284 1 9438
2 60285 1 9438
2 60286 1 9438
2 60287 1 9438
2 60288 1 9438
2 60289 1 9438
2 60290 1 9438
2 60291 1 9438
2 60292 1 9438
2 60293 1 9438
2 60294 1 9438
2 60295 1 9438
2 60296 1 9438
2 60297 1 9438
2 60298 1 9438
2 60299 1 9438
2 60300 1 9438
2 60301 1 9438
2 60302 1 9438
2 60303 1 9438
2 60304 1 9438
2 60305 1 9438
2 60306 1 9438
2 60307 1 9438
2 60308 1 9438
2 60309 1 9438
2 60310 1 9438
2 60311 1 9438
2 60312 1 9438
2 60313 1 9438
2 60314 1 9438
2 60315 1 9440
2 60316 1 9440
2 60317 1 9442
2 60318 1 9442
2 60319 1 9458
2 60320 1 9458
2 60321 1 9458
2 60322 1 9458
2 60323 1 9458
2 60324 1 9458
2 60325 1 9458
2 60326 1 9458
2 60327 1 9458
2 60328 1 9458
2 60329 1 9458
2 60330 1 9458
2 60331 1 9458
2 60332 1 9458
2 60333 1 9459
2 60334 1 9459
2 60335 1 9459
2 60336 1 9460
2 60337 1 9460
2 60338 1 9460
2 60339 1 9460
2 60340 1 9460
2 60341 1 9460
2 60342 1 9460
2 60343 1 9460
2 60344 1 9460
2 60345 1 9460
2 60346 1 9460
2 60347 1 9460
2 60348 1 9463
2 60349 1 9463
2 60350 1 9468
2 60351 1 9468
2 60352 1 9468
2 60353 1 9468
2 60354 1 9468
2 60355 1 9468
2 60356 1 9468
2 60357 1 9469
2 60358 1 9469
2 60359 1 9469
2 60360 1 9470
2 60361 1 9470
2 60362 1 9470
2 60363 1 9479
2 60364 1 9479
2 60365 1 9479
2 60366 1 9479
2 60367 1 9479
2 60368 1 9479
2 60369 1 9479
2 60370 1 9479
2 60371 1 9479
2 60372 1 9479
2 60373 1 9479
2 60374 1 9480
2 60375 1 9480
2 60376 1 9482
2 60377 1 9482
2 60378 1 9483
2 60379 1 9483
2 60380 1 9483
2 60381 1 9483
2 60382 1 9483
2 60383 1 9483
2 60384 1 9484
2 60385 1 9484
2 60386 1 9484
2 60387 1 9492
2 60388 1 9492
2 60389 1 9492
2 60390 1 9493
2 60391 1 9493
2 60392 1 9505
2 60393 1 9505
2 60394 1 9505
2 60395 1 9505
2 60396 1 9505
2 60397 1 9505
2 60398 1 9505
2 60399 1 9505
2 60400 1 9505
2 60401 1 9505
2 60402 1 9505
2 60403 1 9505
2 60404 1 9505
2 60405 1 9505
2 60406 1 9505
2 60407 1 9506
2 60408 1 9506
2 60409 1 9506
2 60410 1 9506
2 60411 1 9506
2 60412 1 9566
2 60413 1 9566
2 60414 1 9566
2 60415 1 9567
2 60416 1 9567
2 60417 1 9569
2 60418 1 9569
2 60419 1 9596
2 60420 1 9596
2 60421 1 9597
2 60422 1 9597
2 60423 1 9597
2 60424 1 9597
2 60425 1 9597
2 60426 1 9600
2 60427 1 9600
2 60428 1 9600
2 60429 1 9600
2 60430 1 9601
2 60431 1 9601
2 60432 1 9603
2 60433 1 9603
2 60434 1 9603
2 60435 1 9603
2 60436 1 9603
2 60437 1 9603
2 60438 1 9603
2 60439 1 9605
2 60440 1 9605
2 60441 1 9607
2 60442 1 9607
2 60443 1 9607
2 60444 1 9610
2 60445 1 9610
2 60446 1 9611
2 60447 1 9611
2 60448 1 9611
2 60449 1 9611
2 60450 1 9611
2 60451 1 9611
2 60452 1 9611
2 60453 1 9611
2 60454 1 9611
2 60455 1 9611
2 60456 1 9611
2 60457 1 9611
2 60458 1 9611
2 60459 1 9611
2 60460 1 9611
2 60461 1 9611
2 60462 1 9611
2 60463 1 9611
2 60464 1 9611
2 60465 1 9611
2 60466 1 9611
2 60467 1 9611
2 60468 1 9611
2 60469 1 9611
2 60470 1 9611
2 60471 1 9611
2 60472 1 9611
2 60473 1 9611
2 60474 1 9612
2 60475 1 9612
2 60476 1 9612
2 60477 1 9612
2 60478 1 9612
2 60479 1 9612
2 60480 1 9620
2 60481 1 9620
2 60482 1 9622
2 60483 1 9622
2 60484 1 9629
2 60485 1 9629
2 60486 1 9629
2 60487 1 9637
2 60488 1 9637
2 60489 1 9653
2 60490 1 9653
2 60491 1 9657
2 60492 1 9657
2 60493 1 9661
2 60494 1 9661
2 60495 1 9662
2 60496 1 9662
2 60497 1 9663
2 60498 1 9663
2 60499 1 9672
2 60500 1 9672
2 60501 1 9672
2 60502 1 9675
2 60503 1 9675
2 60504 1 9692
2 60505 1 9692
2 60506 1 9692
2 60507 1 9692
2 60508 1 9692
2 60509 1 9692
2 60510 1 9692
2 60511 1 9692
2 60512 1 9692
2 60513 1 9692
2 60514 1 9692
2 60515 1 9692
2 60516 1 9692
2 60517 1 9692
2 60518 1 9692
2 60519 1 9692
2 60520 1 9692
2 60521 1 9737
2 60522 1 9737
2 60523 1 9738
2 60524 1 9738
2 60525 1 9749
2 60526 1 9749
2 60527 1 9761
2 60528 1 9761
2 60529 1 9761
2 60530 1 9761
2 60531 1 9761
2 60532 1 9761
2 60533 1 9761
2 60534 1 9761
2 60535 1 9770
2 60536 1 9770
2 60537 1 9770
2 60538 1 9788
2 60539 1 9788
2 60540 1 9791
2 60541 1 9791
2 60542 1 9801
2 60543 1 9801
2 60544 1 9801
2 60545 1 9801
2 60546 1 9803
2 60547 1 9803
2 60548 1 9803
2 60549 1 9818
2 60550 1 9818
2 60551 1 9821
2 60552 1 9821
2 60553 1 9827
2 60554 1 9827
2 60555 1 9837
2 60556 1 9837
2 60557 1 9837
2 60558 1 9837
2 60559 1 9838
2 60560 1 9838
2 60561 1 9838
2 60562 1 9865
2 60563 1 9865
2 60564 1 9865
2 60565 1 9865
2 60566 1 9865
2 60567 1 9865
2 60568 1 9865
2 60569 1 9865
2 60570 1 9865
2 60571 1 9865
2 60572 1 9877
2 60573 1 9877
2 60574 1 9877
2 60575 1 9877
2 60576 1 9877
2 60577 1 9877
2 60578 1 9877
2 60579 1 9877
2 60580 1 9877
2 60581 1 9877
2 60582 1 9877
2 60583 1 9877
2 60584 1 9878
2 60585 1 9878
2 60586 1 9878
2 60587 1 9886
2 60588 1 9886
2 60589 1 9886
2 60590 1 9886
2 60591 1 9886
2 60592 1 9886
2 60593 1 9886
2 60594 1 9886
2 60595 1 9887
2 60596 1 9887
2 60597 1 9890
2 60598 1 9890
2 60599 1 9890
2 60600 1 9890
2 60601 1 9890
2 60602 1 9890
2 60603 1 9891
2 60604 1 9891
2 60605 1 9898
2 60606 1 9898
2 60607 1 9900
2 60608 1 9900
2 60609 1 9910
2 60610 1 9910
2 60611 1 9910
2 60612 1 9950
2 60613 1 9950
2 60614 1 9950
2 60615 1 9950
2 60616 1 9950
2 60617 1 9951
2 60618 1 9951
2 60619 1 9951
2 60620 1 9951
2 60621 1 9951
2 60622 1 9952
2 60623 1 9952
2 60624 1 9955
2 60625 1 9955
2 60626 1 9960
2 60627 1 9960
2 60628 1 9977
2 60629 1 9977
2 60630 1 9977
2 60631 1 9979
2 60632 1 9979
2 60633 1 9980
2 60634 1 9980
2 60635 1 9980
2 60636 1 9980
2 60637 1 9980
2 60638 1 9980
2 60639 1 9983
2 60640 1 9983
2 60641 1 9985
2 60642 1 9985
2 60643 1 9987
2 60644 1 9987
2 60645 1 9989
2 60646 1 9989
2 60647 1 9992
2 60648 1 9992
2 60649 1 9992
2 60650 1 9992
2 60651 1 9993
2 60652 1 9993
2 60653 1 10000
2 60654 1 10000
2 60655 1 10000
2 60656 1 10000
2 60657 1 10000
2 60658 1 10039
2 60659 1 10039
2 60660 1 10040
2 60661 1 10040
2 60662 1 10062
2 60663 1 10062
2 60664 1 10062
2 60665 1 10070
2 60666 1 10070
2 60667 1 10070
2 60668 1 10070
2 60669 1 10070
2 60670 1 10070
2 60671 1 10071
2 60672 1 10071
2 60673 1 10071
2 60674 1 10072
2 60675 1 10072
2 60676 1 10090
2 60677 1 10090
2 60678 1 10090
2 60679 1 10090
2 60680 1 10090
2 60681 1 10090
2 60682 1 10117
2 60683 1 10117
2 60684 1 10117
2 60685 1 10117
2 60686 1 10117
2 60687 1 10117
2 60688 1 10138
2 60689 1 10138
2 60690 1 10138
2 60691 1 10138
2 60692 1 10138
2 60693 1 10139
2 60694 1 10139
2 60695 1 10140
2 60696 1 10140
2 60697 1 10147
2 60698 1 10147
2 60699 1 10147
2 60700 1 10148
2 60701 1 10148
2 60702 1 10148
2 60703 1 10150
2 60704 1 10150
2 60705 1 10150
2 60706 1 10150
2 60707 1 10150
2 60708 1 10150
2 60709 1 10150
2 60710 1 10151
2 60711 1 10151
2 60712 1 10151
2 60713 1 10151
2 60714 1 10151
2 60715 1 10151
2 60716 1 10151
2 60717 1 10161
2 60718 1 10161
2 60719 1 10163
2 60720 1 10163
2 60721 1 10165
2 60722 1 10165
2 60723 1 10166
2 60724 1 10166
2 60725 1 10167
2 60726 1 10167
2 60727 1 10172
2 60728 1 10172
2 60729 1 10172
2 60730 1 10173
2 60731 1 10173
2 60732 1 10177
2 60733 1 10177
2 60734 1 10182
2 60735 1 10182
2 60736 1 10182
2 60737 1 10182
2 60738 1 10193
2 60739 1 10193
2 60740 1 10193
2 60741 1 10193
2 60742 1 10193
2 60743 1 10193
2 60744 1 10194
2 60745 1 10194
2 60746 1 10194
2 60747 1 10196
2 60748 1 10196
2 60749 1 10196
2 60750 1 10196
2 60751 1 10196
2 60752 1 10204
2 60753 1 10204
2 60754 1 10218
2 60755 1 10218
2 60756 1 10238
2 60757 1 10238
2 60758 1 10238
2 60759 1 10248
2 60760 1 10248
2 60761 1 10248
2 60762 1 10249
2 60763 1 10249
2 60764 1 10250
2 60765 1 10250
2 60766 1 10250
2 60767 1 10250
2 60768 1 10251
2 60769 1 10251
2 60770 1 10251
2 60771 1 10251
2 60772 1 10251
2 60773 1 10251
2 60774 1 10251
2 60775 1 10251
2 60776 1 10261
2 60777 1 10261
2 60778 1 10261
2 60779 1 10261
2 60780 1 10261
2 60781 1 10262
2 60782 1 10262
2 60783 1 10262
2 60784 1 10263
2 60785 1 10263
2 60786 1 10264
2 60787 1 10264
2 60788 1 10275
2 60789 1 10275
2 60790 1 10275
2 60791 1 10275
2 60792 1 10275
2 60793 1 10278
2 60794 1 10278
2 60795 1 10281
2 60796 1 10281
2 60797 1 10288
2 60798 1 10288
2 60799 1 10289
2 60800 1 10289
2 60801 1 10290
2 60802 1 10290
2 60803 1 10290
2 60804 1 10290
2 60805 1 10298
2 60806 1 10298
2 60807 1 10310
2 60808 1 10310
2 60809 1 10310
2 60810 1 10310
2 60811 1 10310
2 60812 1 10313
2 60813 1 10313
2 60814 1 10316
2 60815 1 10316
2 60816 1 10318
2 60817 1 10318
2 60818 1 10318
2 60819 1 10318
2 60820 1 10318
2 60821 1 10318
2 60822 1 10318
2 60823 1 10321
2 60824 1 10321
2 60825 1 10321
2 60826 1 10324
2 60827 1 10324
2 60828 1 10325
2 60829 1 10325
2 60830 1 10325
2 60831 1 10329
2 60832 1 10329
2 60833 1 10329
2 60834 1 10330
2 60835 1 10330
2 60836 1 10331
2 60837 1 10331
2 60838 1 10331
2 60839 1 10332
2 60840 1 10332
2 60841 1 10342
2 60842 1 10342
2 60843 1 10342
2 60844 1 10355
2 60845 1 10355
2 60846 1 10356
2 60847 1 10356
2 60848 1 10371
2 60849 1 10371
2 60850 1 10371
2 60851 1 10371
2 60852 1 10371
2 60853 1 10422
2 60854 1 10422
2 60855 1 10423
2 60856 1 10423
2 60857 1 10434
2 60858 1 10434
2 60859 1 10434
2 60860 1 10434
2 60861 1 10451
2 60862 1 10451
2 60863 1 10451
2 60864 1 10504
2 60865 1 10504
2 60866 1 10504
2 60867 1 10505
2 60868 1 10505
2 60869 1 10505
2 60870 1 10509
2 60871 1 10509
2 60872 1 10512
2 60873 1 10512
2 60874 1 10513
2 60875 1 10513
2 60876 1 10518
2 60877 1 10518
2 60878 1 10518
2 60879 1 10526
2 60880 1 10526
2 60881 1 10526
2 60882 1 10526
2 60883 1 10526
2 60884 1 10526
2 60885 1 10527
2 60886 1 10527
2 60887 1 10527
2 60888 1 10542
2 60889 1 10542
2 60890 1 10542
2 60891 1 10542
2 60892 1 10546
2 60893 1 10546
2 60894 1 10557
2 60895 1 10557
2 60896 1 10579
2 60897 1 10579
2 60898 1 10587
2 60899 1 10587
2 60900 1 10587
2 60901 1 10587
2 60902 1 10587
2 60903 1 10588
2 60904 1 10588
2 60905 1 10590
2 60906 1 10590
2 60907 1 10607
2 60908 1 10607
2 60909 1 10607
2 60910 1 10607
2 60911 1 10607
2 60912 1 10607
2 60913 1 10607
2 60914 1 10613
2 60915 1 10613
2 60916 1 10626
2 60917 1 10626
2 60918 1 10656
2 60919 1 10656
2 60920 1 10656
2 60921 1 10657
2 60922 1 10657
2 60923 1 10657
2 60924 1 10657
2 60925 1 10672
2 60926 1 10672
2 60927 1 10674
2 60928 1 10674
2 60929 1 10674
2 60930 1 10674
2 60931 1 10677
2 60932 1 10677
2 60933 1 10690
2 60934 1 10690
2 60935 1 10690
2 60936 1 10692
2 60937 1 10692
2 60938 1 10695
2 60939 1 10695
2 60940 1 10698
2 60941 1 10698
2 60942 1 10698
2 60943 1 10698
2 60944 1 10699
2 60945 1 10699
2 60946 1 10707
2 60947 1 10707
2 60948 1 10712
2 60949 1 10712
2 60950 1 10712
2 60951 1 10712
2 60952 1 10712
2 60953 1 10713
2 60954 1 10713
2 60955 1 10713
2 60956 1 10719
2 60957 1 10719
2 60958 1 10719
2 60959 1 10719
2 60960 1 10719
2 60961 1 10719
2 60962 1 10719
2 60963 1 10730
2 60964 1 10730
2 60965 1 10734
2 60966 1 10734
2 60967 1 10737
2 60968 1 10737
2 60969 1 10737
2 60970 1 10737
2 60971 1 10737
2 60972 1 10737
2 60973 1 10737
2 60974 1 10737
2 60975 1 10737
2 60976 1 10737
2 60977 1 10737
2 60978 1 10737
2 60979 1 10737
2 60980 1 10737
2 60981 1 10737
2 60982 1 10737
2 60983 1 10737
2 60984 1 10738
2 60985 1 10738
2 60986 1 10738
2 60987 1 10738
2 60988 1 10741
2 60989 1 10741
2 60990 1 10744
2 60991 1 10744
2 60992 1 10747
2 60993 1 10747
2 60994 1 10749
2 60995 1 10749
2 60996 1 10765
2 60997 1 10765
2 60998 1 10779
2 60999 1 10779
2 61000 1 10792
2 61001 1 10792
2 61002 1 10792
2 61003 1 10795
2 61004 1 10795
2 61005 1 10798
2 61006 1 10798
2 61007 1 10802
2 61008 1 10802
2 61009 1 10807
2 61010 1 10807
2 61011 1 10814
2 61012 1 10814
2 61013 1 10822
2 61014 1 10822
2 61015 1 10822
2 61016 1 10823
2 61017 1 10823
2 61018 1 10823
2 61019 1 10823
2 61020 1 10823
2 61021 1 10856
2 61022 1 10856
2 61023 1 10856
2 61024 1 10856
2 61025 1 10864
2 61026 1 10864
2 61027 1 10868
2 61028 1 10868
2 61029 1 10868
2 61030 1 10892
2 61031 1 10892
2 61032 1 10893
2 61033 1 10893
2 61034 1 10902
2 61035 1 10902
2 61036 1 10910
2 61037 1 10910
2 61038 1 10912
2 61039 1 10912
2 61040 1 10914
2 61041 1 10914
2 61042 1 10916
2 61043 1 10916
2 61044 1 10916
2 61045 1 10916
2 61046 1 10917
2 61047 1 10917
2 61048 1 10923
2 61049 1 10923
2 61050 1 10928
2 61051 1 10928
2 61052 1 10930
2 61053 1 10930
2 61054 1 10933
2 61055 1 10933
2 61056 1 10956
2 61057 1 10956
2 61058 1 10958
2 61059 1 10958
2 61060 1 10966
2 61061 1 10966
2 61062 1 10966
2 61063 1 10966
2 61064 1 10966
2 61065 1 10971
2 61066 1 10971
2 61067 1 10976
2 61068 1 10976
2 61069 1 10977
2 61070 1 10977
2 61071 1 10978
2 61072 1 10978
2 61073 1 10985
2 61074 1 10985
2 61075 1 10985
2 61076 1 10985
2 61077 1 10986
2 61078 1 10986
2 61079 1 10993
2 61080 1 10993
2 61081 1 10993
2 61082 1 10993
2 61083 1 10994
2 61084 1 10994
2 61085 1 10995
2 61086 1 10995
2 61087 1 11038
2 61088 1 11038
2 61089 1 11039
2 61090 1 11039
2 61091 1 11051
2 61092 1 11051
2 61093 1 11051
2 61094 1 11051
2 61095 1 11051
2 61096 1 11051
2 61097 1 11051
2 61098 1 11051
2 61099 1 11054
2 61100 1 11054
2 61101 1 11054
2 61102 1 11059
2 61103 1 11059
2 61104 1 11061
2 61105 1 11061
2 61106 1 11064
2 61107 1 11064
2 61108 1 11072
2 61109 1 11072
2 61110 1 11074
2 61111 1 11074
2 61112 1 11074
2 61113 1 11074
2 61114 1 11083
2 61115 1 11083
2 61116 1 11085
2 61117 1 11085
2 61118 1 11086
2 61119 1 11086
2 61120 1 11119
2 61121 1 11119
2 61122 1 11132
2 61123 1 11132
2 61124 1 11132
2 61125 1 11132
2 61126 1 11132
2 61127 1 11133
2 61128 1 11133
2 61129 1 11133
2 61130 1 11146
2 61131 1 11146
2 61132 1 11146
2 61133 1 11147
2 61134 1 11147
2 61135 1 11147
2 61136 1 11155
2 61137 1 11155
2 61138 1 11158
2 61139 1 11158
2 61140 1 11158
2 61141 1 11158
2 61142 1 11158
2 61143 1 11168
2 61144 1 11168
2 61145 1 11169
2 61146 1 11169
2 61147 1 11169
2 61148 1 11171
2 61149 1 11171
2 61150 1 11177
2 61151 1 11177
2 61152 1 11177
2 61153 1 11194
2 61154 1 11194
2 61155 1 11194
2 61156 1 11194
2 61157 1 11195
2 61158 1 11195
2 61159 1 11195
2 61160 1 11195
2 61161 1 11196
2 61162 1 11196
2 61163 1 11196
2 61164 1 11196
2 61165 1 11196
2 61166 1 11197
2 61167 1 11197
2 61168 1 11197
2 61169 1 11201
2 61170 1 11201
2 61171 1 11211
2 61172 1 11211
2 61173 1 11220
2 61174 1 11220
2 61175 1 11220
2 61176 1 11235
2 61177 1 11235
2 61178 1 11235
2 61179 1 11235
2 61180 1 11235
2 61181 1 11240
2 61182 1 11240
2 61183 1 11253
2 61184 1 11253
2 61185 1 11264
2 61186 1 11264
2 61187 1 11264
2 61188 1 11264
2 61189 1 11265
2 61190 1 11265
2 61191 1 11265
2 61192 1 11265
2 61193 1 11265
2 61194 1 11265
2 61195 1 11265
2 61196 1 11266
2 61197 1 11266
2 61198 1 11266
2 61199 1 11290
2 61200 1 11290
2 61201 1 11298
2 61202 1 11298
2 61203 1 11312
2 61204 1 11312
2 61205 1 11322
2 61206 1 11322
2 61207 1 11322
2 61208 1 11325
2 61209 1 11325
2 61210 1 11333
2 61211 1 11333
2 61212 1 11333
2 61213 1 11333
2 61214 1 11333
2 61215 1 11334
2 61216 1 11334
2 61217 1 11345
2 61218 1 11345
2 61219 1 11345
2 61220 1 11345
2 61221 1 11345
2 61222 1 11346
2 61223 1 11346
2 61224 1 11379
2 61225 1 11379
2 61226 1 11379
2 61227 1 11390
2 61228 1 11390
2 61229 1 11393
2 61230 1 11393
2 61231 1 11394
2 61232 1 11394
2 61233 1 11397
2 61234 1 11397
2 61235 1 11409
2 61236 1 11409
2 61237 1 11414
2 61238 1 11414
2 61239 1 11414
2 61240 1 11414
2 61241 1 11445
2 61242 1 11445
2 61243 1 11455
2 61244 1 11455
2 61245 1 11464
2 61246 1 11464
2 61247 1 11474
2 61248 1 11474
2 61249 1 11474
2 61250 1 11474
2 61251 1 11475
2 61252 1 11475
2 61253 1 11476
2 61254 1 11476
2 61255 1 11476
2 61256 1 11477
2 61257 1 11477
2 61258 1 11477
2 61259 1 11478
2 61260 1 11478
2 61261 1 11478
2 61262 1 11479
2 61263 1 11479
2 61264 1 11479
2 61265 1 11490
2 61266 1 11490
2 61267 1 11490
2 61268 1 11498
2 61269 1 11498
2 61270 1 11498
2 61271 1 11498
2 61272 1 11508
2 61273 1 11508
2 61274 1 11510
2 61275 1 11510
2 61276 1 11516
2 61277 1 11516
2 61278 1 11516
2 61279 1 11520
2 61280 1 11520
2 61281 1 11520
2 61282 1 11520
2 61283 1 11520
2 61284 1 11520
2 61285 1 11520
2 61286 1 11520
2 61287 1 11520
2 61288 1 11520
2 61289 1 11520
2 61290 1 11520
2 61291 1 11520
2 61292 1 11520
2 61293 1 11520
2 61294 1 11520
2 61295 1 11520
2 61296 1 11528
2 61297 1 11528
2 61298 1 11531
2 61299 1 11531
2 61300 1 11531
2 61301 1 11532
2 61302 1 11532
2 61303 1 11558
2 61304 1 11558
2 61305 1 11569
2 61306 1 11569
2 61307 1 11570
2 61308 1 11570
2 61309 1 11580
2 61310 1 11580
2 61311 1 11587
2 61312 1 11587
2 61313 1 11587
2 61314 1 11587
2 61315 1 11587
2 61316 1 11587
2 61317 1 11587
2 61318 1 11588
2 61319 1 11588
2 61320 1 11588
2 61321 1 11588
2 61322 1 11589
2 61323 1 11589
2 61324 1 11589
2 61325 1 11590
2 61326 1 11590
2 61327 1 11590
2 61328 1 11590
2 61329 1 11591
2 61330 1 11591
2 61331 1 11591
2 61332 1 11591
2 61333 1 11591
2 61334 1 11592
2 61335 1 11592
2 61336 1 11592
2 61337 1 11600
2 61338 1 11600
2 61339 1 11600
2 61340 1 11601
2 61341 1 11601
2 61342 1 11602
2 61343 1 11602
2 61344 1 11602
2 61345 1 11618
2 61346 1 11618
2 61347 1 11638
2 61348 1 11638
2 61349 1 11638
2 61350 1 11643
2 61351 1 11643
2 61352 1 11645
2 61353 1 11645
2 61354 1 11648
2 61355 1 11648
2 61356 1 11648
2 61357 1 11648
2 61358 1 11648
2 61359 1 11657
2 61360 1 11657
2 61361 1 11660
2 61362 1 11660
2 61363 1 11697
2 61364 1 11697
2 61365 1 11697
2 61366 1 11697
2 61367 1 11697
2 61368 1 11698
2 61369 1 11698
2 61370 1 11698
2 61371 1 11698
2 61372 1 11725
2 61373 1 11725
2 61374 1 11729
2 61375 1 11729
2 61376 1 11729
2 61377 1 11730
2 61378 1 11730
2 61379 1 11730
2 61380 1 11739
2 61381 1 11739
2 61382 1 11763
2 61383 1 11763
2 61384 1 11773
2 61385 1 11773
2 61386 1 11782
2 61387 1 11782
2 61388 1 11782
2 61389 1 11783
2 61390 1 11783
2 61391 1 11783
2 61392 1 11791
2 61393 1 11791
2 61394 1 11791
2 61395 1 11795
2 61396 1 11795
2 61397 1 11796
2 61398 1 11796
2 61399 1 11796
2 61400 1 11801
2 61401 1 11801
2 61402 1 11802
2 61403 1 11802
2 61404 1 11802
2 61405 1 11805
2 61406 1 11805
2 61407 1 11806
2 61408 1 11806
2 61409 1 11806
2 61410 1 11806
2 61411 1 11807
2 61412 1 11807
2 61413 1 11808
2 61414 1 11808
2 61415 1 11808
2 61416 1 11808
2 61417 1 11824
2 61418 1 11824
2 61419 1 11824
2 61420 1 11824
2 61421 1 11824
2 61422 1 11824
2 61423 1 11824
2 61424 1 11824
2 61425 1 11824
2 61426 1 11824
2 61427 1 11824
2 61428 1 11824
2 61429 1 11857
2 61430 1 11857
2 61431 1 11857
2 61432 1 11857
2 61433 1 11857
2 61434 1 11857
2 61435 1 11857
2 61436 1 11858
2 61437 1 11858
2 61438 1 11866
2 61439 1 11866
2 61440 1 11868
2 61441 1 11868
2 61442 1 11868
2 61443 1 11869
2 61444 1 11869
2 61445 1 11869
2 61446 1 11870
2 61447 1 11870
2 61448 1 11870
2 61449 1 11871
2 61450 1 11871
2 61451 1 11874
2 61452 1 11874
2 61453 1 11882
2 61454 1 11882
2 61455 1 11882
2 61456 1 11888
2 61457 1 11888
2 61458 1 11902
2 61459 1 11902
2 61460 1 11904
2 61461 1 11904
2 61462 1 11908
2 61463 1 11908
2 61464 1 11909
2 61465 1 11909
2 61466 1 11911
2 61467 1 11911
2 61468 1 11916
2 61469 1 11916
2 61470 1 11917
2 61471 1 11917
2 61472 1 11927
2 61473 1 11927
2 61474 1 11929
2 61475 1 11929
2 61476 1 11939
2 61477 1 11939
2 61478 1 11939
2 61479 1 11941
2 61480 1 11941
2 61481 1 11942
2 61482 1 11942
2 61483 1 11942
2 61484 1 11943
2 61485 1 11943
2 61486 1 11947
2 61487 1 11947
2 61488 1 11948
2 61489 1 11948
2 61490 1 11957
2 61491 1 11957
2 61492 1 11957
2 61493 1 11957
2 61494 1 11958
2 61495 1 11958
2 61496 1 11958
2 61497 1 11960
2 61498 1 11960
2 61499 1 11960
2 61500 1 11960
2 61501 1 11962
2 61502 1 11962
2 61503 1 11975
2 61504 1 11975
2 61505 1 11980
2 61506 1 11980
2 61507 1 11985
2 61508 1 11985
2 61509 1 11987
2 61510 1 11987
2 61511 1 11989
2 61512 1 11989
2 61513 1 12005
2 61514 1 12005
2 61515 1 12016
2 61516 1 12016
2 61517 1 12033
2 61518 1 12033
2 61519 1 12033
2 61520 1 12033
2 61521 1 12033
2 61522 1 12033
2 61523 1 12034
2 61524 1 12034
2 61525 1 12034
2 61526 1 12034
2 61527 1 12035
2 61528 1 12035
2 61529 1 12036
2 61530 1 12036
2 61531 1 12036
2 61532 1 12040
2 61533 1 12040
2 61534 1 12040
2 61535 1 12043
2 61536 1 12043
2 61537 1 12047
2 61538 1 12047
2 61539 1 12065
2 61540 1 12065
2 61541 1 12065
2 61542 1 12065
2 61543 1 12065
2 61544 1 12065
2 61545 1 12066
2 61546 1 12066
2 61547 1 12066
2 61548 1 12066
2 61549 1 12067
2 61550 1 12067
2 61551 1 12067
2 61552 1 12067
2 61553 1 12067
2 61554 1 12067
2 61555 1 12067
2 61556 1 12067
2 61557 1 12071
2 61558 1 12071
2 61559 1 12071
2 61560 1 12071
2 61561 1 12073
2 61562 1 12073
2 61563 1 12073
2 61564 1 12073
2 61565 1 12073
2 61566 1 12073
2 61567 1 12073
2 61568 1 12074
2 61569 1 12074
2 61570 1 12074
2 61571 1 12074
2 61572 1 12076
2 61573 1 12076
2 61574 1 12076
2 61575 1 12076
2 61576 1 12076
2 61577 1 12076
2 61578 1 12076
2 61579 1 12076
2 61580 1 12076
2 61581 1 12076
2 61582 1 12076
2 61583 1 12076
2 61584 1 12076
2 61585 1 12076
2 61586 1 12076
2 61587 1 12077
2 61588 1 12077
2 61589 1 12077
2 61590 1 12077
2 61591 1 12077
2 61592 1 12077
2 61593 1 12077
2 61594 1 12077
2 61595 1 12077
2 61596 1 12077
2 61597 1 12079
2 61598 1 12079
2 61599 1 12082
2 61600 1 12082
2 61601 1 12082
2 61602 1 12082
2 61603 1 12082
2 61604 1 12082
2 61605 1 12087
2 61606 1 12087
2 61607 1 12095
2 61608 1 12095
2 61609 1 12096
2 61610 1 12096
2 61611 1 12109
2 61612 1 12109
2 61613 1 12109
2 61614 1 12110
2 61615 1 12110
2 61616 1 12110
2 61617 1 12110
2 61618 1 12110
2 61619 1 12110
2 61620 1 12111
2 61621 1 12111
2 61622 1 12111
2 61623 1 12132
2 61624 1 12132
2 61625 1 12132
2 61626 1 12135
2 61627 1 12135
2 61628 1 12153
2 61629 1 12153
2 61630 1 12153
2 61631 1 12153
2 61632 1 12156
2 61633 1 12156
2 61634 1 12156
2 61635 1 12157
2 61636 1 12157
2 61637 1 12158
2 61638 1 12158
2 61639 1 12161
2 61640 1 12161
2 61641 1 12161
2 61642 1 12184
2 61643 1 12184
2 61644 1 12185
2 61645 1 12185
2 61646 1 12188
2 61647 1 12188
2 61648 1 12188
2 61649 1 12188
2 61650 1 12189
2 61651 1 12189
2 61652 1 12191
2 61653 1 12191
2 61654 1 12204
2 61655 1 12204
2 61656 1 12204
2 61657 1 12204
2 61658 1 12207
2 61659 1 12207
2 61660 1 12207
2 61661 1 12219
2 61662 1 12219
2 61663 1 12219
2 61664 1 12219
2 61665 1 12219
2 61666 1 12219
2 61667 1 12219
2 61668 1 12219
2 61669 1 12219
2 61670 1 12219
2 61671 1 12219
2 61672 1 12219
2 61673 1 12219
2 61674 1 12219
2 61675 1 12219
2 61676 1 12219
2 61677 1 12219
2 61678 1 12219
2 61679 1 12219
2 61680 1 12219
2 61681 1 12219
2 61682 1 12219
2 61683 1 12220
2 61684 1 12220
2 61685 1 12220
2 61686 1 12220
2 61687 1 12220
2 61688 1 12220
2 61689 1 12220
2 61690 1 12220
2 61691 1 12220
2 61692 1 12228
2 61693 1 12228
2 61694 1 12230
2 61695 1 12230
2 61696 1 12232
2 61697 1 12232
2 61698 1 12233
2 61699 1 12233
2 61700 1 12233
2 61701 1 12235
2 61702 1 12235
2 61703 1 12237
2 61704 1 12237
2 61705 1 12238
2 61706 1 12238
2 61707 1 12239
2 61708 1 12239
2 61709 1 12245
2 61710 1 12245
2 61711 1 12272
2 61712 1 12272
2 61713 1 12272
2 61714 1 12272
2 61715 1 12272
2 61716 1 12272
2 61717 1 12273
2 61718 1 12273
2 61719 1 12286
2 61720 1 12286
2 61721 1 12286
2 61722 1 12286
2 61723 1 12286
2 61724 1 12287
2 61725 1 12287
2 61726 1 12292
2 61727 1 12292
2 61728 1 12295
2 61729 1 12295
2 61730 1 12299
2 61731 1 12299
2 61732 1 12312
2 61733 1 12312
2 61734 1 12316
2 61735 1 12316
2 61736 1 12323
2 61737 1 12323
2 61738 1 12323
2 61739 1 12323
2 61740 1 12323
2 61741 1 12323
2 61742 1 12323
2 61743 1 12323
2 61744 1 12323
2 61745 1 12323
2 61746 1 12323
2 61747 1 12323
2 61748 1 12323
2 61749 1 12323
2 61750 1 12323
2 61751 1 12323
2 61752 1 12323
2 61753 1 12323
2 61754 1 12323
2 61755 1 12323
2 61756 1 12323
2 61757 1 12323
2 61758 1 12323
2 61759 1 12324
2 61760 1 12324
2 61761 1 12324
2 61762 1 12324
2 61763 1 12324
2 61764 1 12325
2 61765 1 12325
2 61766 1 12325
2 61767 1 12325
2 61768 1 12325
2 61769 1 12326
2 61770 1 12326
2 61771 1 12347
2 61772 1 12347
2 61773 1 12347
2 61774 1 12347
2 61775 1 12363
2 61776 1 12363
2 61777 1 12363
2 61778 1 12363
2 61779 1 12363
2 61780 1 12363
2 61781 1 12405
2 61782 1 12405
2 61783 1 12422
2 61784 1 12422
2 61785 1 12422
2 61786 1 12422
2 61787 1 12423
2 61788 1 12423
2 61789 1 12436
2 61790 1 12436
2 61791 1 12457
2 61792 1 12457
2 61793 1 12457
2 61794 1 12457
2 61795 1 12460
2 61796 1 12460
2 61797 1 12460
2 61798 1 12460
2 61799 1 12460
2 61800 1 12468
2 61801 1 12468
2 61802 1 12468
2 61803 1 12468
2 61804 1 12468
2 61805 1 12469
2 61806 1 12469
2 61807 1 12496
2 61808 1 12496
2 61809 1 12496
2 61810 1 12496
2 61811 1 12496
2 61812 1 12496
2 61813 1 12497
2 61814 1 12497
2 61815 1 12497
2 61816 1 12497
2 61817 1 12498
2 61818 1 12498
2 61819 1 12499
2 61820 1 12499
2 61821 1 12499
2 61822 1 12499
2 61823 1 12501
2 61824 1 12501
2 61825 1 12517
2 61826 1 12517
2 61827 1 12518
2 61828 1 12518
2 61829 1 12518
2 61830 1 12518
2 61831 1 12518
2 61832 1 12518
2 61833 1 12519
2 61834 1 12519
2 61835 1 12531
2 61836 1 12531
2 61837 1 12532
2 61838 1 12532
2 61839 1 12532
2 61840 1 12532
2 61841 1 12532
2 61842 1 12532
2 61843 1 12548
2 61844 1 12548
2 61845 1 12548
2 61846 1 12548
2 61847 1 12550
2 61848 1 12550
2 61849 1 12550
2 61850 1 12551
2 61851 1 12551
2 61852 1 12553
2 61853 1 12553
2 61854 1 12554
2 61855 1 12554
2 61856 1 12554
2 61857 1 12554
2 61858 1 12555
2 61859 1 12555
2 61860 1 12556
2 61861 1 12556
2 61862 1 12565
2 61863 1 12565
2 61864 1 12565
2 61865 1 12565
2 61866 1 12565
2 61867 1 12565
2 61868 1 12565
2 61869 1 12565
2 61870 1 12565
2 61871 1 12565
2 61872 1 12566
2 61873 1 12566
2 61874 1 12566
2 61875 1 12567
2 61876 1 12567
2 61877 1 12567
2 61878 1 12567
2 61879 1 12567
2 61880 1 12567
2 61881 1 12567
2 61882 1 12576
2 61883 1 12576
2 61884 1 12576
2 61885 1 12577
2 61886 1 12577
2 61887 1 12577
2 61888 1 12577
2 61889 1 12577
2 61890 1 12577
2 61891 1 12577
2 61892 1 12578
2 61893 1 12578
2 61894 1 12578
2 61895 1 12578
2 61896 1 12578
2 61897 1 12578
2 61898 1 12579
2 61899 1 12579
2 61900 1 12579
2 61901 1 12579
2 61902 1 12579
2 61903 1 12581
2 61904 1 12581
2 61905 1 12583
2 61906 1 12583
2 61907 1 12585
2 61908 1 12585
2 61909 1 12601
2 61910 1 12601
2 61911 1 12601
2 61912 1 12606
2 61913 1 12606
2 61914 1 12606
2 61915 1 12607
2 61916 1 12607
2 61917 1 12608
2 61918 1 12608
2 61919 1 12608
2 61920 1 12608
2 61921 1 12608
2 61922 1 12608
2 61923 1 12608
2 61924 1 12608
2 61925 1 12608
2 61926 1 12608
2 61927 1 12619
2 61928 1 12619
2 61929 1 12619
2 61930 1 12619
2 61931 1 12619
2 61932 1 12619
2 61933 1 12619
2 61934 1 12619
2 61935 1 12619
2 61936 1 12619
2 61937 1 12619
2 61938 1 12620
2 61939 1 12620
2 61940 1 12620
2 61941 1 12621
2 61942 1 12621
2 61943 1 12621
2 61944 1 12621
2 61945 1 12630
2 61946 1 12630
2 61947 1 12633
2 61948 1 12633
2 61949 1 12638
2 61950 1 12638
2 61951 1 12638
2 61952 1 12638
2 61953 1 12638
2 61954 1 12638
2 61955 1 12638
2 61956 1 12638
2 61957 1 12638
2 61958 1 12648
2 61959 1 12648
2 61960 1 12648
2 61961 1 12648
2 61962 1 12648
2 61963 1 12648
2 61964 1 12648
2 61965 1 12648
2 61966 1 12648
2 61967 1 12648
2 61968 1 12648
2 61969 1 12649
2 61970 1 12649
2 61971 1 12650
2 61972 1 12650
2 61973 1 12650
2 61974 1 12651
2 61975 1 12651
2 61976 1 12651
2 61977 1 12651
2 61978 1 12651
2 61979 1 12651
2 61980 1 12651
2 61981 1 12653
2 61982 1 12653
2 61983 1 12655
2 61984 1 12655
2 61985 1 12655
2 61986 1 12655
2 61987 1 12655
2 61988 1 12655
2 61989 1 12662
2 61990 1 12662
2 61991 1 12662
2 61992 1 12662
2 61993 1 12663
2 61994 1 12663
2 61995 1 12665
2 61996 1 12665
2 61997 1 12665
2 61998 1 12672
2 61999 1 12672
2 62000 1 12672
2 62001 1 12672
2 62002 1 12672
2 62003 1 12673
2 62004 1 12673
2 62005 1 12673
2 62006 1 12673
2 62007 1 12673
2 62008 1 12682
2 62009 1 12682
2 62010 1 12682
2 62011 1 12683
2 62012 1 12683
2 62013 1 12686
2 62014 1 12686
2 62015 1 12686
2 62016 1 12688
2 62017 1 12688
2 62018 1 12688
2 62019 1 12688
2 62020 1 12688
2 62021 1 12688
2 62022 1 12688
2 62023 1 12688
2 62024 1 12689
2 62025 1 12689
2 62026 1 12689
2 62027 1 12689
2 62028 1 12690
2 62029 1 12690
2 62030 1 12691
2 62031 1 12691
2 62032 1 12692
2 62033 1 12692
2 62034 1 12705
2 62035 1 12705
2 62036 1 12705
2 62037 1 12705
2 62038 1 12705
2 62039 1 12705
2 62040 1 12705
2 62041 1 12705
2 62042 1 12705
2 62043 1 12706
2 62044 1 12706
2 62045 1 12706
2 62046 1 12706
2 62047 1 12706
2 62048 1 12709
2 62049 1 12709
2 62050 1 12711
2 62051 1 12711
2 62052 1 12711
2 62053 1 12711
2 62054 1 12711
2 62055 1 12711
2 62056 1 12711
2 62057 1 12712
2 62058 1 12712
2 62059 1 12712
2 62060 1 12721
2 62061 1 12721
2 62062 1 12721
2 62063 1 12721
2 62064 1 12722
2 62065 1 12722
2 62066 1 12722
2 62067 1 12722
2 62068 1 12722
2 62069 1 12752
2 62070 1 12752
2 62071 1 12752
2 62072 1 12755
2 62073 1 12755
2 62074 1 12759
2 62075 1 12759
2 62076 1 12762
2 62077 1 12762
2 62078 1 12762
2 62079 1 12762
2 62080 1 12762
2 62081 1 12762
2 62082 1 12764
2 62083 1 12764
2 62084 1 12764
2 62085 1 12765
2 62086 1 12765
2 62087 1 12767
2 62088 1 12767
2 62089 1 12767
2 62090 1 12791
2 62091 1 12791
2 62092 1 12791
2 62093 1 12791
2 62094 1 12791
2 62095 1 12791
2 62096 1 12793
2 62097 1 12793
2 62098 1 12793
2 62099 1 12794
2 62100 1 12794
2 62101 1 12808
2 62102 1 12808
2 62103 1 12811
2 62104 1 12811
2 62105 1 12811
2 62106 1 12811
2 62107 1 12811
2 62108 1 12818
2 62109 1 12818
2 62110 1 12819
2 62111 1 12819
2 62112 1 12822
2 62113 1 12822
2 62114 1 12823
2 62115 1 12823
2 62116 1 12824
2 62117 1 12824
2 62118 1 12824
2 62119 1 12824
2 62120 1 12824
2 62121 1 12824
2 62122 1 12824
2 62123 1 12824
2 62124 1 12824
2 62125 1 12824
2 62126 1 12824
2 62127 1 12824
2 62128 1 12824
2 62129 1 12825
2 62130 1 12825
2 62131 1 12850
2 62132 1 12850
2 62133 1 12850
2 62134 1 12850
2 62135 1 12851
2 62136 1 12851
2 62137 1 12851
2 62138 1 12852
2 62139 1 12852
2 62140 1 12855
2 62141 1 12855
2 62142 1 12855
2 62143 1 12859
2 62144 1 12859
2 62145 1 12863
2 62146 1 12863
2 62147 1 12863
2 62148 1 12863
2 62149 1 12864
2 62150 1 12864
2 62151 1 12884
2 62152 1 12884
2 62153 1 12884
2 62154 1 12884
2 62155 1 12885
2 62156 1 12885
2 62157 1 12895
2 62158 1 12895
2 62159 1 12895
2 62160 1 12896
2 62161 1 12896
2 62162 1 12896
2 62163 1 12896
2 62164 1 12897
2 62165 1 12897
2 62166 1 12931
2 62167 1 12931
2 62168 1 12934
2 62169 1 12934
2 62170 1 12949
2 62171 1 12949
2 62172 1 12950
2 62173 1 12950
2 62174 1 12950
2 62175 1 12950
2 62176 1 12950
2 62177 1 12976
2 62178 1 12976
2 62179 1 12999
2 62180 1 12999
2 62181 1 12999
2 62182 1 13038
2 62183 1 13038
2 62184 1 13045
2 62185 1 13045
2 62186 1 13053
2 62187 1 13053
2 62188 1 13056
2 62189 1 13056
2 62190 1 13056
2 62191 1 13067
2 62192 1 13067
2 62193 1 13067
2 62194 1 13067
2 62195 1 13076
2 62196 1 13076
2 62197 1 13085
2 62198 1 13085
2 62199 1 13085
2 62200 1 13094
2 62201 1 13094
2 62202 1 13098
2 62203 1 13098
2 62204 1 13098
2 62205 1 13108
2 62206 1 13108
2 62207 1 13108
2 62208 1 13108
2 62209 1 13109
2 62210 1 13109
2 62211 1 13109
2 62212 1 13130
2 62213 1 13130
2 62214 1 13130
2 62215 1 13152
2 62216 1 13152
2 62217 1 13162
2 62218 1 13162
2 62219 1 13162
2 62220 1 13162
2 62221 1 13162
2 62222 1 13165
2 62223 1 13165
2 62224 1 13172
2 62225 1 13172
2 62226 1 13172
2 62227 1 13172
2 62228 1 13172
2 62229 1 13178
2 62230 1 13178
2 62231 1 13178
2 62232 1 13179
2 62233 1 13179
2 62234 1 13179
2 62235 1 13179
2 62236 1 13193
2 62237 1 13193
2 62238 1 13194
2 62239 1 13194
2 62240 1 13194
2 62241 1 13194
2 62242 1 13194
2 62243 1 13194
2 62244 1 13215
2 62245 1 13215
2 62246 1 13215
2 62247 1 13215
2 62248 1 13215
2 62249 1 13216
2 62250 1 13216
2 62251 1 13216
2 62252 1 13216
2 62253 1 13217
2 62254 1 13217
2 62255 1 13218
2 62256 1 13218
2 62257 1 13218
2 62258 1 13218
2 62259 1 13218
2 62260 1 13219
2 62261 1 13219
2 62262 1 13227
2 62263 1 13227
2 62264 1 13236
2 62265 1 13236
2 62266 1 13238
2 62267 1 13238
2 62268 1 13250
2 62269 1 13250
2 62270 1 13250
2 62271 1 13250
2 62272 1 13250
2 62273 1 13250
2 62274 1 13253
2 62275 1 13253
2 62276 1 13253
2 62277 1 13254
2 62278 1 13254
2 62279 1 13254
2 62280 1 13254
2 62281 1 13254
2 62282 1 13279
2 62283 1 13279
2 62284 1 13293
2 62285 1 13293
2 62286 1 13293
2 62287 1 13293
2 62288 1 13298
2 62289 1 13298
2 62290 1 13298
2 62291 1 13298
2 62292 1 13299
2 62293 1 13299
2 62294 1 13299
2 62295 1 13299
2 62296 1 13300
2 62297 1 13300
2 62298 1 13302
2 62299 1 13302
2 62300 1 13302
2 62301 1 13306
2 62302 1 13306
2 62303 1 13306
2 62304 1 13306
2 62305 1 13306
2 62306 1 13307
2 62307 1 13307
2 62308 1 13307
2 62309 1 13320
2 62310 1 13320
2 62311 1 13320
2 62312 1 13321
2 62313 1 13321
2 62314 1 13321
2 62315 1 13322
2 62316 1 13322
2 62317 1 13325
2 62318 1 13325
2 62319 1 13333
2 62320 1 13333
2 62321 1 13334
2 62322 1 13334
2 62323 1 13334
2 62324 1 13343
2 62325 1 13343
2 62326 1 13344
2 62327 1 13344
2 62328 1 13345
2 62329 1 13345
2 62330 1 13347
2 62331 1 13347
2 62332 1 13353
2 62333 1 13353
2 62334 1 13353
2 62335 1 13353
2 62336 1 13354
2 62337 1 13354
2 62338 1 13354
2 62339 1 13355
2 62340 1 13355
2 62341 1 13356
2 62342 1 13356
2 62343 1 13356
2 62344 1 13357
2 62345 1 13357
2 62346 1 13366
2 62347 1 13366
2 62348 1 13366
2 62349 1 13366
2 62350 1 13382
2 62351 1 13382
2 62352 1 13382
2 62353 1 13382
2 62354 1 13387
2 62355 1 13387
2 62356 1 13389
2 62357 1 13389
2 62358 1 13399
2 62359 1 13399
2 62360 1 13399
2 62361 1 13409
2 62362 1 13409
2 62363 1 13412
2 62364 1 13412
2 62365 1 13412
2 62366 1 13412
2 62367 1 13412
2 62368 1 13412
2 62369 1 13417
2 62370 1 13417
2 62371 1 13417
2 62372 1 13417
2 62373 1 13417
2 62374 1 13418
2 62375 1 13418
2 62376 1 13418
2 62377 1 13418
2 62378 1 13426
2 62379 1 13426
2 62380 1 13426
2 62381 1 13426
2 62382 1 13426
2 62383 1 13426
2 62384 1 13426
2 62385 1 13430
2 62386 1 13430
2 62387 1 13430
2 62388 1 13430
2 62389 1 13431
2 62390 1 13431
2 62391 1 13432
2 62392 1 13432
2 62393 1 13440
2 62394 1 13440
2 62395 1 13440
2 62396 1 13440
2 62397 1 13440
2 62398 1 13440
2 62399 1 13440
2 62400 1 13440
2 62401 1 13440
2 62402 1 13440
2 62403 1 13453
2 62404 1 13453
2 62405 1 13453
2 62406 1 13453
2 62407 1 13455
2 62408 1 13455
2 62409 1 13470
2 62410 1 13470
2 62411 1 13470
2 62412 1 13470
2 62413 1 13471
2 62414 1 13471
2 62415 1 13472
2 62416 1 13472
2 62417 1 13476
2 62418 1 13476
2 62419 1 13476
2 62420 1 13476
2 62421 1 13477
2 62422 1 13477
2 62423 1 13487
2 62424 1 13487
2 62425 1 13487
2 62426 1 13490
2 62427 1 13490
2 62428 1 13503
2 62429 1 13503
2 62430 1 13503
2 62431 1 13503
2 62432 1 13519
2 62433 1 13519
2 62434 1 13519
2 62435 1 13519
2 62436 1 13528
2 62437 1 13528
2 62438 1 13528
2 62439 1 13528
2 62440 1 13528
2 62441 1 13528
2 62442 1 13528
2 62443 1 13548
2 62444 1 13548
2 62445 1 13556
2 62446 1 13556
2 62447 1 13556
2 62448 1 13556
2 62449 1 13564
2 62450 1 13564
2 62451 1 13572
2 62452 1 13572
2 62453 1 13602
2 62454 1 13602
2 62455 1 13602
2 62456 1 13602
2 62457 1 13602
2 62458 1 13602
2 62459 1 13603
2 62460 1 13603
2 62461 1 13603
2 62462 1 13616
2 62463 1 13616
2 62464 1 13617
2 62465 1 13617
2 62466 1 13646
2 62467 1 13646
2 62468 1 13646
2 62469 1 13649
2 62470 1 13649
2 62471 1 13650
2 62472 1 13650
2 62473 1 13664
2 62474 1 13664
2 62475 1 13664
2 62476 1 13665
2 62477 1 13665
2 62478 1 13685
2 62479 1 13685
2 62480 1 13686
2 62481 1 13686
2 62482 1 13686
2 62483 1 13686
2 62484 1 13686
2 62485 1 13686
2 62486 1 13689
2 62487 1 13689
2 62488 1 13689
2 62489 1 13690
2 62490 1 13690
2 62491 1 13691
2 62492 1 13691
2 62493 1 13704
2 62494 1 13704
2 62495 1 13704
2 62496 1 13704
2 62497 1 13705
2 62498 1 13705
2 62499 1 13708
2 62500 1 13708
2 62501 1 13708
2 62502 1 13708
2 62503 1 13711
2 62504 1 13711
2 62505 1 13711
2 62506 1 13712
2 62507 1 13712
2 62508 1 13712
2 62509 1 13757
2 62510 1 13757
2 62511 1 13782
2 62512 1 13782
2 62513 1 13796
2 62514 1 13796
2 62515 1 13796
2 62516 1 13796
2 62517 1 13796
2 62518 1 13796
2 62519 1 13796
2 62520 1 13796
2 62521 1 13796
2 62522 1 13796
2 62523 1 13796
2 62524 1 13796
2 62525 1 13796
2 62526 1 13797
2 62527 1 13797
2 62528 1 13800
2 62529 1 13800
2 62530 1 13800
2 62531 1 13801
2 62532 1 13801
2 62533 1 13802
2 62534 1 13802
2 62535 1 13802
2 62536 1 13802
2 62537 1 13802
2 62538 1 13802
2 62539 1 13803
2 62540 1 13803
2 62541 1 13804
2 62542 1 13804
2 62543 1 13808
2 62544 1 13808
2 62545 1 13809
2 62546 1 13809
2 62547 1 13812
2 62548 1 13812
2 62549 1 13813
2 62550 1 13813
2 62551 1 13820
2 62552 1 13820
2 62553 1 13820
2 62554 1 13820
2 62555 1 13820
2 62556 1 13820
2 62557 1 13821
2 62558 1 13821
2 62559 1 13821
2 62560 1 13822
2 62561 1 13822
2 62562 1 13843
2 62563 1 13843
2 62564 1 13843
2 62565 1 13843
2 62566 1 13849
2 62567 1 13849
2 62568 1 13869
2 62569 1 13869
2 62570 1 13891
2 62571 1 13891
2 62572 1 13892
2 62573 1 13892
2 62574 1 13892
2 62575 1 13896
2 62576 1 13896
2 62577 1 13896
2 62578 1 13896
2 62579 1 13896
2 62580 1 13896
2 62581 1 13903
2 62582 1 13903
2 62583 1 13903
2 62584 1 13911
2 62585 1 13911
2 62586 1 13914
2 62587 1 13914
2 62588 1 13919
2 62589 1 13919
2 62590 1 13919
2 62591 1 13922
2 62592 1 13922
2 62593 1 13933
2 62594 1 13933
2 62595 1 13944
2 62596 1 13944
2 62597 1 13955
2 62598 1 13955
2 62599 1 13963
2 62600 1 13963
2 62601 1 14020
2 62602 1 14020
2 62603 1 14020
2 62604 1 14033
2 62605 1 14033
2 62606 1 14033
2 62607 1 14033
2 62608 1 14033
2 62609 1 14043
2 62610 1 14043
2 62611 1 14043
2 62612 1 14043
2 62613 1 14043
2 62614 1 14063
2 62615 1 14063
2 62616 1 14063
2 62617 1 14063
2 62618 1 14063
2 62619 1 14064
2 62620 1 14064
2 62621 1 14065
2 62622 1 14065
2 62623 1 14065
2 62624 1 14087
2 62625 1 14087
2 62626 1 14106
2 62627 1 14106
2 62628 1 14106
2 62629 1 14108
2 62630 1 14108
2 62631 1 14108
2 62632 1 14108
2 62633 1 14130
2 62634 1 14130
2 62635 1 14130
2 62636 1 14130
2 62637 1 14143
2 62638 1 14143
2 62639 1 14143
2 62640 1 14174
2 62641 1 14174
2 62642 1 14174
2 62643 1 14175
2 62644 1 14175
2 62645 1 14175
2 62646 1 14190
2 62647 1 14190
2 62648 1 14190
2 62649 1 14190
2 62650 1 14190
2 62651 1 14205
2 62652 1 14205
2 62653 1 14206
2 62654 1 14206
2 62655 1 14214
2 62656 1 14214
2 62657 1 14214
2 62658 1 14219
2 62659 1 14219
2 62660 1 14219
2 62661 1 14222
2 62662 1 14222
2 62663 1 14223
2 62664 1 14223
2 62665 1 14224
2 62666 1 14224
2 62667 1 14235
2 62668 1 14235
2 62669 1 14235
2 62670 1 14237
2 62671 1 14237
2 62672 1 14248
2 62673 1 14248
2 62674 1 14248
2 62675 1 14255
2 62676 1 14255
2 62677 1 14255
2 62678 1 14255
2 62679 1 14255
2 62680 1 14256
2 62681 1 14256
2 62682 1 14256
2 62683 1 14298
2 62684 1 14298
2 62685 1 14310
2 62686 1 14310
2 62687 1 14313
2 62688 1 14313
2 62689 1 14313
2 62690 1 14321
2 62691 1 14321
2 62692 1 14321
2 62693 1 14338
2 62694 1 14338
2 62695 1 14346
2 62696 1 14346
2 62697 1 14346
2 62698 1 14346
2 62699 1 14362
2 62700 1 14362
2 62701 1 14373
2 62702 1 14373
2 62703 1 14373
2 62704 1 14373
2 62705 1 14374
2 62706 1 14374
2 62707 1 14374
2 62708 1 14374
2 62709 1 14374
2 62710 1 14374
2 62711 1 14374
2 62712 1 14410
2 62713 1 14410
2 62714 1 14430
2 62715 1 14430
2 62716 1 14439
2 62717 1 14439
2 62718 1 14462
2 62719 1 14462
2 62720 1 14462
2 62721 1 14468
2 62722 1 14468
2 62723 1 14471
2 62724 1 14471
2 62725 1 14471
2 62726 1 14475
2 62727 1 14475
2 62728 1 14478
2 62729 1 14478
2 62730 1 14478
2 62731 1 14478
2 62732 1 14478
2 62733 1 14481
2 62734 1 14481
2 62735 1 14481
2 62736 1 14481
2 62737 1 14481
2 62738 1 14482
2 62739 1 14482
2 62740 1 14488
2 62741 1 14488
2 62742 1 14488
2 62743 1 14492
2 62744 1 14492
2 62745 1 14493
2 62746 1 14493
2 62747 1 14493
2 62748 1 14493
2 62749 1 14505
2 62750 1 14505
2 62751 1 14505
2 62752 1 14510
2 62753 1 14510
2 62754 1 14510
2 62755 1 14510
2 62756 1 14510
2 62757 1 14510
2 62758 1 14510
2 62759 1 14529
2 62760 1 14529
2 62761 1 14529
2 62762 1 14529
2 62763 1 14529
2 62764 1 14529
2 62765 1 14529
2 62766 1 14529
2 62767 1 14529
2 62768 1 14529
2 62769 1 14529
2 62770 1 14529
2 62771 1 14529
2 62772 1 14530
2 62773 1 14530
2 62774 1 14530
2 62775 1 14539
2 62776 1 14539
2 62777 1 14540
2 62778 1 14540
2 62779 1 14540
2 62780 1 14540
2 62781 1 14540
2 62782 1 14562
2 62783 1 14562
2 62784 1 14564
2 62785 1 14564
2 62786 1 14564
2 62787 1 14564
2 62788 1 14565
2 62789 1 14565
2 62790 1 14577
2 62791 1 14577
2 62792 1 14580
2 62793 1 14580
2 62794 1 14580
2 62795 1 14580
2 62796 1 14580
2 62797 1 14580
2 62798 1 14580
2 62799 1 14580
2 62800 1 14580
2 62801 1 14580
2 62802 1 14580
2 62803 1 14580
2 62804 1 14580
2 62805 1 14580
2 62806 1 14580
2 62807 1 14580
2 62808 1 14580
2 62809 1 14581
2 62810 1 14581
2 62811 1 14581
2 62812 1 14581
2 62813 1 14581
2 62814 1 14581
2 62815 1 14581
2 62816 1 14581
2 62817 1 14581
2 62818 1 14581
2 62819 1 14581
2 62820 1 14581
2 62821 1 14581
2 62822 1 14581
2 62823 1 14581
2 62824 1 14581
2 62825 1 14581
2 62826 1 14581
2 62827 1 14581
2 62828 1 14581
2 62829 1 14581
2 62830 1 14581
2 62831 1 14581
2 62832 1 14582
2 62833 1 14582
2 62834 1 14584
2 62835 1 14584
2 62836 1 14596
2 62837 1 14596
2 62838 1 14596
2 62839 1 14597
2 62840 1 14597
2 62841 1 14599
2 62842 1 14599
2 62843 1 14599
2 62844 1 14599
2 62845 1 14606
2 62846 1 14606
2 62847 1 14606
2 62848 1 14606
2 62849 1 14606
2 62850 1 14606
2 62851 1 14623
2 62852 1 14623
2 62853 1 14623
2 62854 1 14649
2 62855 1 14649
2 62856 1 14650
2 62857 1 14650
2 62858 1 14650
2 62859 1 14650
2 62860 1 14650
2 62861 1 14650
2 62862 1 14650
2 62863 1 14679
2 62864 1 14679
2 62865 1 14686
2 62866 1 14686
2 62867 1 14687
2 62868 1 14687
2 62869 1 14722
2 62870 1 14722
2 62871 1 14727
2 62872 1 14727
2 62873 1 14734
2 62874 1 14734
2 62875 1 14737
2 62876 1 14737
2 62877 1 14753
2 62878 1 14753
2 62879 1 14753
2 62880 1 14753
2 62881 1 14753
2 62882 1 14753
2 62883 1 14755
2 62884 1 14755
2 62885 1 14755
2 62886 1 14764
2 62887 1 14764
2 62888 1 14764
2 62889 1 14764
2 62890 1 14765
2 62891 1 14765
2 62892 1 14765
2 62893 1 14765
2 62894 1 14769
2 62895 1 14769
2 62896 1 14772
2 62897 1 14772
2 62898 1 14785
2 62899 1 14785
2 62900 1 14785
2 62901 1 14787
2 62902 1 14787
2 62903 1 14787
2 62904 1 14805
2 62905 1 14805
2 62906 1 14805
2 62907 1 14805
2 62908 1 14806
2 62909 1 14806
2 62910 1 14806
2 62911 1 14832
2 62912 1 14832
2 62913 1 14853
2 62914 1 14853
2 62915 1 14853
2 62916 1 14869
2 62917 1 14869
2 62918 1 14902
2 62919 1 14902
2 62920 1 14906
2 62921 1 14906
2 62922 1 14925
2 62923 1 14925
2 62924 1 14925
2 62925 1 14925
2 62926 1 14925
2 62927 1 14925
2 62928 1 14925
2 62929 1 14925
2 62930 1 14926
2 62931 1 14926
2 62932 1 14926
2 62933 1 14928
2 62934 1 14928
2 62935 1 14932
2 62936 1 14932
2 62937 1 14933
2 62938 1 14933
2 62939 1 14957
2 62940 1 14957
2 62941 1 14958
2 62942 1 14958
2 62943 1 14977
2 62944 1 14977
2 62945 1 14977
2 62946 1 14977
2 62947 1 14977
2 62948 1 14997
2 62949 1 14997
2 62950 1 14997
2 62951 1 14998
2 62952 1 14998
2 62953 1 15015
2 62954 1 15015
2 62955 1 15020
2 62956 1 15020
2 62957 1 15021
2 62958 1 15021
2 62959 1 15050
2 62960 1 15050
2 62961 1 15064
2 62962 1 15064
2 62963 1 15064
2 62964 1 15064
2 62965 1 15064
2 62966 1 15064
2 62967 1 15064
2 62968 1 15064
2 62969 1 15066
2 62970 1 15066
2 62971 1 15074
2 62972 1 15074
2 62973 1 15074
2 62974 1 15074
2 62975 1 15074
2 62976 1 15074
2 62977 1 15074
2 62978 1 15074
2 62979 1 15075
2 62980 1 15075
2 62981 1 15075
2 62982 1 15075
2 62983 1 15075
2 62984 1 15083
2 62985 1 15083
2 62986 1 15091
2 62987 1 15091
2 62988 1 15091
2 62989 1 15096
2 62990 1 15096
2 62991 1 15096
2 62992 1 15096
2 62993 1 15096
2 62994 1 15104
2 62995 1 15104
2 62996 1 15110
2 62997 1 15110
2 62998 1 15148
2 62999 1 15148
2 63000 1 15148
2 63001 1 15148
2 63002 1 15148
2 63003 1 15148
2 63004 1 15152
2 63005 1 15152
2 63006 1 15176
2 63007 1 15176
2 63008 1 15176
2 63009 1 15176
2 63010 1 15176
2 63011 1 15176
2 63012 1 15176
2 63013 1 15178
2 63014 1 15178
2 63015 1 15200
2 63016 1 15200
2 63017 1 15201
2 63018 1 15201
2 63019 1 15212
2 63020 1 15212
2 63021 1 15220
2 63022 1 15220
2 63023 1 15232
2 63024 1 15232
2 63025 1 15255
2 63026 1 15255
2 63027 1 15255
2 63028 1 15301
2 63029 1 15301
2 63030 1 15301
2 63031 1 15301
2 63032 1 15301
2 63033 1 15301
2 63034 1 15302
2 63035 1 15302
2 63036 1 15302
2 63037 1 15312
2 63038 1 15312
2 63039 1 15315
2 63040 1 15315
2 63041 1 15323
2 63042 1 15323
2 63043 1 15323
2 63044 1 15323
2 63045 1 15324
2 63046 1 15324
2 63047 1 15332
2 63048 1 15332
2 63049 1 15337
2 63050 1 15337
2 63051 1 15337
2 63052 1 15337
2 63053 1 15353
2 63054 1 15353
2 63055 1 15361
2 63056 1 15361
2 63057 1 15361
2 63058 1 15361
2 63059 1 15361
2 63060 1 15361
2 63061 1 15362
2 63062 1 15362
2 63063 1 15369
2 63064 1 15369
2 63065 1 15369
2 63066 1 15369
2 63067 1 15369
2 63068 1 15395
2 63069 1 15395
2 63070 1 15395
2 63071 1 15395
2 63072 1 15396
2 63073 1 15396
2 63074 1 15396
2 63075 1 15396
2 63076 1 15396
2 63077 1 15396
2 63078 1 15396
2 63079 1 15396
2 63080 1 15396
2 63081 1 15396
2 63082 1 15397
2 63083 1 15397
2 63084 1 15397
2 63085 1 15397
2 63086 1 15397
2 63087 1 15397
2 63088 1 15398
2 63089 1 15398
2 63090 1 15411
2 63091 1 15411
2 63092 1 15416
2 63093 1 15416
2 63094 1 15416
2 63095 1 15417
2 63096 1 15417
2 63097 1 15417
2 63098 1 15417
2 63099 1 15444
2 63100 1 15444
2 63101 1 15456
2 63102 1 15456
2 63103 1 15456
2 63104 1 15501
2 63105 1 15501
2 63106 1 15501
2 63107 1 15501
2 63108 1 15501
2 63109 1 15501
2 63110 1 15502
2 63111 1 15502
2 63112 1 15503
2 63113 1 15503
2 63114 1 15503
2 63115 1 15536
2 63116 1 15536
2 63117 1 15574
2 63118 1 15574
2 63119 1 15574
2 63120 1 15575
2 63121 1 15575
2 63122 1 15617
2 63123 1 15617
2 63124 1 15630
2 63125 1 15630
2 63126 1 15653
2 63127 1 15653
2 63128 1 15653
2 63129 1 15653
2 63130 1 15653
2 63131 1 15656
2 63132 1 15656
2 63133 1 15657
2 63134 1 15657
2 63135 1 15657
2 63136 1 15721
2 63137 1 15721
2 63138 1 15721
2 63139 1 15723
2 63140 1 15723
2 63141 1 15726
2 63142 1 15726
2 63143 1 15726
2 63144 1 15726
2 63145 1 15781
2 63146 1 15781
2 63147 1 15782
2 63148 1 15782
2 63149 1 15782
2 63150 1 15782
2 63151 1 15783
2 63152 1 15783
2 63153 1 15795
2 63154 1 15795
2 63155 1 15795
2 63156 1 15795
2 63157 1 15808
2 63158 1 15808
2 63159 1 15808
2 63160 1 15811
2 63161 1 15811
2 63162 1 15811
2 63163 1 15811
2 63164 1 15812
2 63165 1 15812
2 63166 1 15812
2 63167 1 15827
2 63168 1 15827
2 63169 1 15829
2 63170 1 15829
2 63171 1 15849
2 63172 1 15849
2 63173 1 15884
2 63174 1 15884
2 63175 1 15924
2 63176 1 15924
2 63177 1 15947
2 63178 1 15947
2 63179 1 15958
2 63180 1 15958
2 63181 1 15973
2 63182 1 15973
2 63183 1 15973
2 63184 1 16018
2 63185 1 16018
2 63186 1 16018
2 63187 1 16018
2 63188 1 16020
2 63189 1 16020
2 63190 1 16020
2 63191 1 16020
2 63192 1 16031
2 63193 1 16031
2 63194 1 16065
2 63195 1 16065
2 63196 1 16065
2 63197 1 16065
2 63198 1 16065
2 63199 1 16065
2 63200 1 16065
2 63201 1 16065
2 63202 1 16065
2 63203 1 16078
2 63204 1 16078
2 63205 1 16079
2 63206 1 16079
2 63207 1 16091
2 63208 1 16091
2 63209 1 16126
2 63210 1 16126
2 63211 1 16126
2 63212 1 16134
2 63213 1 16134
2 63214 1 16134
2 63215 1 16134
2 63216 1 16141
2 63217 1 16141
2 63218 1 16141
2 63219 1 16144
2 63220 1 16144
2 63221 1 16145
2 63222 1 16145
2 63223 1 16154
2 63224 1 16154
2 63225 1 16154
2 63226 1 16154
2 63227 1 16193
2 63228 1 16193
2 63229 1 16193
2 63230 1 16197
2 63231 1 16197
2 63232 1 16197
2 63233 1 16217
2 63234 1 16217
2 63235 1 16217
2 63236 1 16217
2 63237 1 16217
2 63238 1 16217
2 63239 1 16219
2 63240 1 16219
2 63241 1 16222
2 63242 1 16222
2 63243 1 16222
2 63244 1 16222
2 63245 1 16229
2 63246 1 16229
2 63247 1 16229
2 63248 1 16251
2 63249 1 16251
2 63250 1 16259
2 63251 1 16259
2 63252 1 16260
2 63253 1 16260
2 63254 1 16260
2 63255 1 16261
2 63256 1 16261
2 63257 1 16262
2 63258 1 16262
2 63259 1 16282
2 63260 1 16282
2 63261 1 16282
2 63262 1 16290
2 63263 1 16290
2 63264 1 16291
2 63265 1 16291
2 63266 1 16299
2 63267 1 16299
2 63268 1 16299
2 63269 1 16299
2 63270 1 16308
2 63271 1 16308
2 63272 1 16308
2 63273 1 16308
2 63274 1 16322
2 63275 1 16322
2 63276 1 16325
2 63277 1 16325
2 63278 1 16325
2 63279 1 16335
2 63280 1 16335
2 63281 1 16335
2 63282 1 16335
2 63283 1 16335
2 63284 1 16335
2 63285 1 16335
2 63286 1 16335
2 63287 1 16335
2 63288 1 16336
2 63289 1 16336
2 63290 1 16336
2 63291 1 16336
2 63292 1 16336
2 63293 1 16341
2 63294 1 16341
2 63295 1 16341
2 63296 1 16341
2 63297 1 16349
2 63298 1 16349
2 63299 1 16349
2 63300 1 16349
2 63301 1 16349
2 63302 1 16349
2 63303 1 16351
2 63304 1 16351
2 63305 1 16351
2 63306 1 16354
2 63307 1 16354
2 63308 1 16355
2 63309 1 16355
2 63310 1 16359
2 63311 1 16359
2 63312 1 16373
2 63313 1 16373
2 63314 1 16373
2 63315 1 16373
2 63316 1 16373
2 63317 1 16373
2 63318 1 16374
2 63319 1 16374
2 63320 1 16374
2 63321 1 16375
2 63322 1 16375
2 63323 1 16376
2 63324 1 16376
2 63325 1 16405
2 63326 1 16405
2 63327 1 16406
2 63328 1 16406
2 63329 1 16406
2 63330 1 16409
2 63331 1 16409
2 63332 1 16410
2 63333 1 16410
2 63334 1 16411
2 63335 1 16411
2 63336 1 16411
2 63337 1 16428
2 63338 1 16428
2 63339 1 16429
2 63340 1 16429
2 63341 1 16429
2 63342 1 16429
2 63343 1 16429
2 63344 1 16440
2 63345 1 16440
2 63346 1 16440
2 63347 1 16440
2 63348 1 16440
2 63349 1 16531
2 63350 1 16531
2 63351 1 16541
2 63352 1 16541
2 63353 1 16541
2 63354 1 16561
2 63355 1 16561
2 63356 1 16574
2 63357 1 16574
2 63358 1 16574
2 63359 1 16575
2 63360 1 16575
2 63361 1 16609
2 63362 1 16609
2 63363 1 16613
2 63364 1 16613
2 63365 1 16618
2 63366 1 16618
2 63367 1 16650
2 63368 1 16650
2 63369 1 16650
2 63370 1 16650
2 63371 1 16651
2 63372 1 16651
2 63373 1 16652
2 63374 1 16652
2 63375 1 16668
2 63376 1 16668
2 63377 1 16693
2 63378 1 16693
2 63379 1 16726
2 63380 1 16726
2 63381 1 16726
2 63382 1 16785
2 63383 1 16785
2 63384 1 16806
2 63385 1 16806
2 63386 1 16814
2 63387 1 16814
2 63388 1 16814
2 63389 1 16814
2 63390 1 16839
2 63391 1 16839
2 63392 1 16859
2 63393 1 16859
2 63394 1 16903
2 63395 1 16903
2 63396 1 16905
2 63397 1 16905
2 63398 1 16906
2 63399 1 16906
2 63400 1 16914
2 63401 1 16914
2 63402 1 16914
2 63403 1 16916
2 63404 1 16916
2 63405 1 16916
2 63406 1 16926
2 63407 1 16926
2 63408 1 16949
2 63409 1 16949
2 63410 1 16962
2 63411 1 16962
2 63412 1 16977
2 63413 1 16977
2 63414 1 16977
2 63415 1 16977
2 63416 1 16977
2 63417 1 16977
2 63418 1 16998
2 63419 1 16998
2 63420 1 16998
2 63421 1 16998
2 63422 1 16999
2 63423 1 16999
2 63424 1 16999
2 63425 1 16999
2 63426 1 17000
2 63427 1 17000
2 63428 1 17000
2 63429 1 17000
2 63430 1 17000
2 63431 1 17009
2 63432 1 17009
2 63433 1 17009
2 63434 1 17009
2 63435 1 17009
2 63436 1 17009
2 63437 1 17009
2 63438 1 17010
2 63439 1 17010
2 63440 1 17010
2 63441 1 17010
2 63442 1 17011
2 63443 1 17011
2 63444 1 17011
2 63445 1 17022
2 63446 1 17022
2 63447 1 17023
2 63448 1 17023
2 63449 1 17035
2 63450 1 17035
2 63451 1 17060
2 63452 1 17060
2 63453 1 17064
2 63454 1 17064
2 63455 1 17076
2 63456 1 17076
2 63457 1 17081
2 63458 1 17081
2 63459 1 17095
2 63460 1 17095
2 63461 1 17095
2 63462 1 17096
2 63463 1 17096
2 63464 1 17103
2 63465 1 17103
2 63466 1 17118
2 63467 1 17118
2 63468 1 17125
2 63469 1 17125
2 63470 1 17125
2 63471 1 17133
2 63472 1 17133
2 63473 1 17133
2 63474 1 17140
2 63475 1 17140
2 63476 1 17169
2 63477 1 17169
2 63478 1 17169
2 63479 1 17169
2 63480 1 17169
2 63481 1 17169
2 63482 1 17173
2 63483 1 17173
2 63484 1 17182
2 63485 1 17182
2 63486 1 17182
2 63487 1 17182
2 63488 1 17182
2 63489 1 17182
2 63490 1 17206
2 63491 1 17206
2 63492 1 17206
2 63493 1 17206
2 63494 1 17207
2 63495 1 17207
2 63496 1 17207
2 63497 1 17238
2 63498 1 17238
2 63499 1 17241
2 63500 1 17241
2 63501 1 17241
2 63502 1 17242
2 63503 1 17242
2 63504 1 17243
2 63505 1 17243
2 63506 1 17244
2 63507 1 17244
2 63508 1 17244
2 63509 1 17270
2 63510 1 17270
2 63511 1 17291
2 63512 1 17291
2 63513 1 17292
2 63514 1 17292
2 63515 1 17294
2 63516 1 17294
2 63517 1 17305
2 63518 1 17305
2 63519 1 17316
2 63520 1 17316
2 63521 1 17316
2 63522 1 17316
2 63523 1 17324
2 63524 1 17324
2 63525 1 17324
2 63526 1 17324
2 63527 1 17325
2 63528 1 17325
2 63529 1 17326
2 63530 1 17326
2 63531 1 17347
2 63532 1 17347
2 63533 1 17348
2 63534 1 17348
2 63535 1 17352
2 63536 1 17352
2 63537 1 17352
2 63538 1 17352
2 63539 1 17352
2 63540 1 17352
2 63541 1 17352
2 63542 1 17352
2 63543 1 17363
2 63544 1 17363
2 63545 1 17366
2 63546 1 17366
2 63547 1 17445
2 63548 1 17445
2 63549 1 17448
2 63550 1 17448
2 63551 1 17448
2 63552 1 17448
2 63553 1 17449
2 63554 1 17449
2 63555 1 17463
2 63556 1 17463
2 63557 1 17470
2 63558 1 17470
2 63559 1 17471
2 63560 1 17471
2 63561 1 17471
2 63562 1 17475
2 63563 1 17475
2 63564 1 17477
2 63565 1 17477
2 63566 1 17495
2 63567 1 17495
2 63568 1 17496
2 63569 1 17496
2 63570 1 17498
2 63571 1 17498
2 63572 1 17499
2 63573 1 17499
2 63574 1 17499
2 63575 1 17499
2 63576 1 17499
2 63577 1 17499
2 63578 1 17499
2 63579 1 17499
2 63580 1 17499
2 63581 1 17499
2 63582 1 17499
2 63583 1 17499
2 63584 1 17503
2 63585 1 17503
2 63586 1 17525
2 63587 1 17525
2 63588 1 17526
2 63589 1 17526
2 63590 1 17526
2 63591 1 17527
2 63592 1 17527
2 63593 1 17527
2 63594 1 17527
2 63595 1 17528
2 63596 1 17528
2 63597 1 17531
2 63598 1 17531
2 63599 1 17532
2 63600 1 17532
2 63601 1 17533
2 63602 1 17533
2 63603 1 17533
2 63604 1 17533
2 63605 1 17533
2 63606 1 17534
2 63607 1 17534
2 63608 1 17534
2 63609 1 17537
2 63610 1 17537
2 63611 1 17541
2 63612 1 17541
2 63613 1 17542
2 63614 1 17542
2 63615 1 17542
2 63616 1 17542
2 63617 1 17545
2 63618 1 17545
2 63619 1 17545
2 63620 1 17545
2 63621 1 17545
2 63622 1 17546
2 63623 1 17546
2 63624 1 17561
2 63625 1 17561
2 63626 1 17566
2 63627 1 17566
2 63628 1 17567
2 63629 1 17567
2 63630 1 17567
2 63631 1 17567
2 63632 1 17568
2 63633 1 17568
2 63634 1 17579
2 63635 1 17579
2 63636 1 17579
2 63637 1 17580
2 63638 1 17580
2 63639 1 17580
2 63640 1 17580
2 63641 1 17590
2 63642 1 17590
2 63643 1 17590
2 63644 1 17590
2 63645 1 17590
2 63646 1 17590
2 63647 1 17605
2 63648 1 17605
2 63649 1 17605
2 63650 1 17609
2 63651 1 17609
2 63652 1 17623
2 63653 1 17623
2 63654 1 17623
2 63655 1 17623
2 63656 1 17624
2 63657 1 17624
2 63658 1 17625
2 63659 1 17625
2 63660 1 17627
2 63661 1 17627
2 63662 1 17628
2 63663 1 17628
2 63664 1 17628
2 63665 1 17628
2 63666 1 17628
2 63667 1 17628
2 63668 1 17628
2 63669 1 17628
2 63670 1 17636
2 63671 1 17636
2 63672 1 17637
2 63673 1 17637
2 63674 1 17650
2 63675 1 17650
2 63676 1 17650
2 63677 1 17679
2 63678 1 17679
2 63679 1 17679
2 63680 1 17679
2 63681 1 17679
2 63682 1 17679
2 63683 1 17702
2 63684 1 17702
2 63685 1 17706
2 63686 1 17706
2 63687 1 17718
2 63688 1 17718
2 63689 1 17718
2 63690 1 17731
2 63691 1 17731
2 63692 1 17734
2 63693 1 17734
2 63694 1 17742
2 63695 1 17742
2 63696 1 17743
2 63697 1 17743
2 63698 1 17743
2 63699 1 17744
2 63700 1 17744
2 63701 1 17747
2 63702 1 17747
2 63703 1 17749
2 63704 1 17749
2 63705 1 17765
2 63706 1 17765
2 63707 1 17765
2 63708 1 17765
2 63709 1 17765
2 63710 1 17765
2 63711 1 17775
2 63712 1 17775
2 63713 1 17776
2 63714 1 17776
2 63715 1 17780
2 63716 1 17780
2 63717 1 17781
2 63718 1 17781
2 63719 1 17784
2 63720 1 17784
2 63721 1 17784
2 63722 1 17804
2 63723 1 17804
2 63724 1 17804
2 63725 1 17804
2 63726 1 17807
2 63727 1 17807
2 63728 1 17824
2 63729 1 17824
2 63730 1 17825
2 63731 1 17825
2 63732 1 17829
2 63733 1 17829
2 63734 1 17829
2 63735 1 17829
2 63736 1 17829
2 63737 1 17831
2 63738 1 17831
2 63739 1 17847
2 63740 1 17847
2 63741 1 17847
2 63742 1 17847
2 63743 1 17850
2 63744 1 17850
2 63745 1 17852
2 63746 1 17852
2 63747 1 17859
2 63748 1 17859
2 63749 1 17866
2 63750 1 17866
2 63751 1 17871
2 63752 1 17871
2 63753 1 17919
2 63754 1 17919
2 63755 1 17919
2 63756 1 17919
2 63757 1 17919
2 63758 1 17929
2 63759 1 17929
2 63760 1 17930
2 63761 1 17930
2 63762 1 17930
2 63763 1 17947
2 63764 1 17947
2 63765 1 17947
2 63766 1 17947
2 63767 1 17947
2 63768 1 17947
2 63769 1 17947
2 63770 1 17947
2 63771 1 17947
2 63772 1 17948
2 63773 1 17948
2 63774 1 17948
2 63775 1 17948
2 63776 1 17948
2 63777 1 17948
2 63778 1 17948
2 63779 1 17975
2 63780 1 17975
2 63781 1 17976
2 63782 1 17976
2 63783 1 17997
2 63784 1 17997
2 63785 1 17997
2 63786 1 17997
2 63787 1 17997
2 63788 1 17997
2 63789 1 17997
2 63790 1 17997
2 63791 1 17997
2 63792 1 17997
2 63793 1 17998
2 63794 1 17998
2 63795 1 17998
2 63796 1 17998
2 63797 1 17998
2 63798 1 17998
2 63799 1 17998
2 63800 1 18001
2 63801 1 18001
2 63802 1 18024
2 63803 1 18024
2 63804 1 18028
2 63805 1 18028
2 63806 1 18028
2 63807 1 18028
2 63808 1 18031
2 63809 1 18031
2 63810 1 18042
2 63811 1 18042
2 63812 1 18077
2 63813 1 18077
2 63814 1 18077
2 63815 1 18077
2 63816 1 18077
2 63817 1 18078
2 63818 1 18078
2 63819 1 18088
2 63820 1 18088
2 63821 1 18091
2 63822 1 18091
2 63823 1 18105
2 63824 1 18105
2 63825 1 18105
2 63826 1 18106
2 63827 1 18106
2 63828 1 18113
2 63829 1 18113
2 63830 1 18123
2 63831 1 18123
2 63832 1 18123
2 63833 1 18123
2 63834 1 18123
2 63835 1 18123
2 63836 1 18123
2 63837 1 18132
2 63838 1 18132
2 63839 1 18137
2 63840 1 18137
2 63841 1 18137
2 63842 1 18137
2 63843 1 18137
2 63844 1 18137
2 63845 1 18137
2 63846 1 18149
2 63847 1 18149
2 63848 1 18157
2 63849 1 18157
2 63850 1 18207
2 63851 1 18207
2 63852 1 18224
2 63853 1 18224
2 63854 1 18224
2 63855 1 18224
2 63856 1 18224
2 63857 1 18224
2 63858 1 18224
2 63859 1 18249
2 63860 1 18249
2 63861 1 18302
2 63862 1 18302
2 63863 1 18307
2 63864 1 18307
2 63865 1 18309
2 63866 1 18309
2 63867 1 18332
2 63868 1 18332
2 63869 1 18341
2 63870 1 18341
2 63871 1 18344
2 63872 1 18344
2 63873 1 18359
2 63874 1 18359
2 63875 1 18360
2 63876 1 18360
2 63877 1 18377
2 63878 1 18377
2 63879 1 18378
2 63880 1 18378
2 63881 1 18383
2 63882 1 18383
2 63883 1 18390
2 63884 1 18390
2 63885 1 18390
2 63886 1 18393
2 63887 1 18393
2 63888 1 18393
2 63889 1 18393
2 63890 1 18393
2 63891 1 18393
2 63892 1 18393
2 63893 1 18393
2 63894 1 18393
2 63895 1 18409
2 63896 1 18409
2 63897 1 18409
2 63898 1 18417
2 63899 1 18417
2 63900 1 18439
2 63901 1 18439
2 63902 1 18445
2 63903 1 18445
2 63904 1 18445
2 63905 1 18458
2 63906 1 18458
2 63907 1 18458
2 63908 1 18458
2 63909 1 18458
2 63910 1 18458
2 63911 1 18458
2 63912 1 18458
2 63913 1 18459
2 63914 1 18459
2 63915 1 18460
2 63916 1 18460
2 63917 1 18469
2 63918 1 18469
2 63919 1 18469
2 63920 1 18469
2 63921 1 18469
2 63922 1 18469
2 63923 1 18478
2 63924 1 18478
2 63925 1 18487
2 63926 1 18487
2 63927 1 18487
2 63928 1 18487
2 63929 1 18487
2 63930 1 18490
2 63931 1 18490
2 63932 1 18505
2 63933 1 18505
2 63934 1 18512
2 63935 1 18512
2 63936 1 18532
2 63937 1 18532
2 63938 1 18533
2 63939 1 18533
2 63940 1 18537
2 63941 1 18537
2 63942 1 18546
2 63943 1 18546
2 63944 1 18548
2 63945 1 18548
2 63946 1 18554
2 63947 1 18554
2 63948 1 18565
2 63949 1 18565
2 63950 1 18565
2 63951 1 18565
2 63952 1 18567
2 63953 1 18567
2 63954 1 18571
2 63955 1 18571
2 63956 1 18571
2 63957 1 18594
2 63958 1 18594
2 63959 1 18594
2 63960 1 18598
2 63961 1 18598
2 63962 1 18611
2 63963 1 18611
2 63964 1 18634
2 63965 1 18634
2 63966 1 18635
2 63967 1 18635
2 63968 1 18635
2 63969 1 18642
2 63970 1 18642
2 63971 1 18642
2 63972 1 18642
2 63973 1 18642
2 63974 1 18642
2 63975 1 18642
2 63976 1 18685
2 63977 1 18685
2 63978 1 18690
2 63979 1 18690
2 63980 1 18697
2 63981 1 18697
2 63982 1 18700
2 63983 1 18700
2 63984 1 18717
2 63985 1 18717
2 63986 1 18746
2 63987 1 18746
2 63988 1 18778
2 63989 1 18778
2 63990 1 18791
2 63991 1 18791
2 63992 1 18802
2 63993 1 18802
2 63994 1 18818
2 63995 1 18818
2 63996 1 18818
2 63997 1 18819
2 63998 1 18819
2 63999 1 18836
2 64000 1 18836
2 64001 1 18837
2 64002 1 18837
2 64003 1 18844
2 64004 1 18844
2 64005 1 18844
2 64006 1 18867
2 64007 1 18867
2 64008 1 18871
2 64009 1 18871
2 64010 1 18879
2 64011 1 18879
2 64012 1 18892
2 64013 1 18892
2 64014 1 18892
2 64015 1 18892
2 64016 1 18892
2 64017 1 18892
2 64018 1 18892
2 64019 1 18892
2 64020 1 18892
2 64021 1 18892
2 64022 1 18892
2 64023 1 18938
2 64024 1 18938
2 64025 1 18938
2 64026 1 18939
2 64027 1 18939
2 64028 1 18947
2 64029 1 18947
2 64030 1 18973
2 64031 1 18973
2 64032 1 18974
2 64033 1 18974
2 64034 1 18974
2 64035 1 18983
2 64036 1 18983
2 64037 1 19001
2 64038 1 19001
2 64039 1 19001
2 64040 1 19001
2 64041 1 19001
2 64042 1 19004
2 64043 1 19004
2 64044 1 19005
2 64045 1 19005
2 64046 1 19005
2 64047 1 19005
2 64048 1 19005
2 64049 1 19005
2 64050 1 19006
2 64051 1 19006
2 64052 1 19006
2 64053 1 19006
2 64054 1 19016
2 64055 1 19016
2 64056 1 19018
2 64057 1 19018
2 64058 1 19018
2 64059 1 19018
2 64060 1 19023
2 64061 1 19023
2 64062 1 19023
2 64063 1 19024
2 64064 1 19024
2 64065 1 19024
2 64066 1 19033
2 64067 1 19033
2 64068 1 19043
2 64069 1 19043
2 64070 1 19045
2 64071 1 19045
2 64072 1 19045
2 64073 1 19045
2 64074 1 19045
2 64075 1 19062
2 64076 1 19062
2 64077 1 19062
2 64078 1 19062
2 64079 1 19065
2 64080 1 19065
2 64081 1 19092
2 64082 1 19092
2 64083 1 19093
2 64084 1 19093
2 64085 1 19110
2 64086 1 19110
2 64087 1 19118
2 64088 1 19118
2 64089 1 19118
2 64090 1 19119
2 64091 1 19119
2 64092 1 19121
2 64093 1 19121
2 64094 1 19122
2 64095 1 19122
2 64096 1 19169
2 64097 1 19169
2 64098 1 19169
2 64099 1 19202
2 64100 1 19202
2 64101 1 19202
2 64102 1 19202
2 64103 1 19202
2 64104 1 19203
2 64105 1 19203
2 64106 1 19203
2 64107 1 19203
2 64108 1 19203
2 64109 1 19210
2 64110 1 19210
2 64111 1 19220
2 64112 1 19220
2 64113 1 19227
2 64114 1 19227
2 64115 1 19227
2 64116 1 19228
2 64117 1 19228
2 64118 1 19229
2 64119 1 19229
2 64120 1 19229
2 64121 1 19229
2 64122 1 19229
2 64123 1 19240
2 64124 1 19240
2 64125 1 19240
2 64126 1 19240
2 64127 1 19240
2 64128 1 19244
2 64129 1 19244
2 64130 1 19245
2 64131 1 19245
2 64132 1 19246
2 64133 1 19246
2 64134 1 19252
2 64135 1 19252
2 64136 1 19252
2 64137 1 19252
2 64138 1 19252
2 64139 1 19252
2 64140 1 19252
2 64141 1 19262
2 64142 1 19262
2 64143 1 19263
2 64144 1 19263
2 64145 1 19265
2 64146 1 19265
2 64147 1 19273
2 64148 1 19273
2 64149 1 19274
2 64150 1 19274
2 64151 1 19274
2 64152 1 19274
2 64153 1 19274
2 64154 1 19274
2 64155 1 19288
2 64156 1 19288
2 64157 1 19288
2 64158 1 19289
2 64159 1 19289
2 64160 1 19297
2 64161 1 19297
2 64162 1 19313
2 64163 1 19313
2 64164 1 19313
2 64165 1 19313
2 64166 1 19313
2 64167 1 19314
2 64168 1 19314
2 64169 1 19314
2 64170 1 19319
2 64171 1 19319
2 64172 1 19324
2 64173 1 19324
2 64174 1 19336
2 64175 1 19336
2 64176 1 19336
2 64177 1 19336
2 64178 1 19336
2 64179 1 19358
2 64180 1 19358
2 64181 1 19358
2 64182 1 19359
2 64183 1 19359
2 64184 1 19382
2 64185 1 19382
2 64186 1 19391
2 64187 1 19391
2 64188 1 19399
2 64189 1 19399
2 64190 1 19399
2 64191 1 19408
2 64192 1 19408
2 64193 1 19417
2 64194 1 19417
2 64195 1 19440
2 64196 1 19440
2 64197 1 19440
2 64198 1 19446
2 64199 1 19446
2 64200 1 19447
2 64201 1 19447
2 64202 1 19455
2 64203 1 19455
2 64204 1 19464
2 64205 1 19464
2 64206 1 19472
2 64207 1 19472
2 64208 1 19472
2 64209 1 19475
2 64210 1 19475
2 64211 1 19475
2 64212 1 19475
2 64213 1 19475
2 64214 1 19475
2 64215 1 19478
2 64216 1 19478
2 64217 1 19486
2 64218 1 19486
2 64219 1 19488
2 64220 1 19488
2 64221 1 19501
2 64222 1 19501
2 64223 1 19502
2 64224 1 19502
2 64225 1 19502
2 64226 1 19502
2 64227 1 19502
2 64228 1 19510
2 64229 1 19510
2 64230 1 19527
2 64231 1 19527
2 64232 1 19544
2 64233 1 19544
2 64234 1 19554
2 64235 1 19554
2 64236 1 19577
2 64237 1 19577
2 64238 1 19577
2 64239 1 19585
2 64240 1 19585
2 64241 1 19625
2 64242 1 19625
2 64243 1 19625
2 64244 1 19638
2 64245 1 19638
2 64246 1 19638
2 64247 1 19653
2 64248 1 19653
2 64249 1 19665
2 64250 1 19665
2 64251 1 19672
2 64252 1 19672
2 64253 1 19686
2 64254 1 19686
2 64255 1 19686
2 64256 1 19689
2 64257 1 19689
2 64258 1 19689
2 64259 1 19691
2 64260 1 19691
2 64261 1 19691
2 64262 1 19691
2 64263 1 19691
2 64264 1 19691
2 64265 1 19691
2 64266 1 19691
2 64267 1 19691
2 64268 1 19692
2 64269 1 19692
2 64270 1 19703
2 64271 1 19703
2 64272 1 19704
2 64273 1 19704
2 64274 1 19705
2 64275 1 19705
2 64276 1 19705
2 64277 1 19712
2 64278 1 19712
2 64279 1 19712
2 64280 1 19736
2 64281 1 19736
2 64282 1 19744
2 64283 1 19744
2 64284 1 19744
2 64285 1 19758
2 64286 1 19758
2 64287 1 19760
2 64288 1 19760
2 64289 1 19760
2 64290 1 19760
2 64291 1 19760
2 64292 1 19779
2 64293 1 19779
2 64294 1 19779
2 64295 1 19786
2 64296 1 19786
2 64297 1 19786
2 64298 1 19797
2 64299 1 19797
2 64300 1 19822
2 64301 1 19822
2 64302 1 19822
2 64303 1 19828
2 64304 1 19828
2 64305 1 19830
2 64306 1 19830
2 64307 1 19831
2 64308 1 19831
2 64309 1 19831
2 64310 1 19831
2 64311 1 19831
2 64312 1 19831
2 64313 1 19831
2 64314 1 19832
2 64315 1 19832
2 64316 1 19839
2 64317 1 19839
2 64318 1 19847
2 64319 1 19847
2 64320 1 19847
2 64321 1 19856
2 64322 1 19856
2 64323 1 19858
2 64324 1 19858
2 64325 1 19858
2 64326 1 19859
2 64327 1 19859
2 64328 1 19862
2 64329 1 19862
2 64330 1 19863
2 64331 1 19863
2 64332 1 19881
2 64333 1 19881
2 64334 1 19882
2 64335 1 19882
2 64336 1 19882
2 64337 1 19882
2 64338 1 19896
2 64339 1 19896
2 64340 1 19899
2 64341 1 19899
2 64342 1 19899
2 64343 1 19919
2 64344 1 19919
2 64345 1 19919
2 64346 1 19926
2 64347 1 19926
2 64348 1 19934
2 64349 1 19934
2 64350 1 19934
2 64351 1 19934
2 64352 1 19934
2 64353 1 19934
2 64354 1 19935
2 64355 1 19935
2 64356 1 19943
2 64357 1 19943
2 64358 1 19943
2 64359 1 19943
2 64360 1 19981
2 64361 1 19981
2 64362 1 19981
2 64363 1 19981
2 64364 1 20001
2 64365 1 20001
2 64366 1 20001
2 64367 1 20001
2 64368 1 20001
2 64369 1 20003
2 64370 1 20003
2 64371 1 20009
2 64372 1 20009
2 64373 1 20034
2 64374 1 20034
2 64375 1 20034
2 64376 1 20066
2 64377 1 20066
2 64378 1 20087
2 64379 1 20087
2 64380 1 20106
2 64381 1 20106
2 64382 1 20121
2 64383 1 20121
2 64384 1 20121
2 64385 1 20121
2 64386 1 20121
2 64387 1 20121
2 64388 1 20126
2 64389 1 20126
2 64390 1 20139
2 64391 1 20139
2 64392 1 20147
2 64393 1 20147
2 64394 1 20172
2 64395 1 20172
2 64396 1 20189
2 64397 1 20189
2 64398 1 20189
2 64399 1 20189
2 64400 1 20189
2 64401 1 20191
2 64402 1 20191
2 64403 1 20229
2 64404 1 20229
2 64405 1 20229
2 64406 1 20229
2 64407 1 20229
2 64408 1 20232
2 64409 1 20232
2 64410 1 20250
2 64411 1 20250
2 64412 1 20286
2 64413 1 20286
2 64414 1 20297
2 64415 1 20297
2 64416 1 20297
2 64417 1 20297
2 64418 1 20297
2 64419 1 20297
2 64420 1 20297
2 64421 1 20297
2 64422 1 20298
2 64423 1 20298
2 64424 1 20331
2 64425 1 20331
2 64426 1 20372
2 64427 1 20372
2 64428 1 20373
2 64429 1 20373
2 64430 1 20374
2 64431 1 20374
2 64432 1 20375
2 64433 1 20375
2 64434 1 20405
2 64435 1 20405
2 64436 1 20425
2 64437 1 20425
2 64438 1 20434
2 64439 1 20434
2 64440 1 20435
2 64441 1 20435
2 64442 1 20435
2 64443 1 20462
2 64444 1 20462
2 64445 1 20469
2 64446 1 20469
2 64447 1 20470
2 64448 1 20470
2 64449 1 20614
2 64450 1 20614
2 64451 1 20631
2 64452 1 20631
2 64453 1 20632
2 64454 1 20632
2 64455 1 20632
2 64456 1 20632
2 64457 1 20636
2 64458 1 20636
2 64459 1 20638
2 64460 1 20638
2 64461 1 20647
2 64462 1 20647
2 64463 1 20647
2 64464 1 20654
2 64465 1 20654
2 64466 1 20698
2 64467 1 20698
2 64468 1 20751
2 64469 1 20751
2 64470 1 20754
2 64471 1 20754
2 64472 1 20764
2 64473 1 20764
2 64474 1 20764
2 64475 1 20764
2 64476 1 20764
2 64477 1 20764
2 64478 1 20764
2 64479 1 20767
2 64480 1 20767
2 64481 1 20782
2 64482 1 20782
2 64483 1 20803
2 64484 1 20803
2 64485 1 20846
2 64486 1 20846
2 64487 1 20860
2 64488 1 20860
2 64489 1 20860
2 64490 1 20866
2 64491 1 20866
2 64492 1 20876
2 64493 1 20876
2 64494 1 20880
2 64495 1 20880
2 64496 1 20883
2 64497 1 20883
2 64498 1 20884
2 64499 1 20884
2 64500 1 20892
2 64501 1 20892
2 64502 1 20893
2 64503 1 20893
2 64504 1 20893
2 64505 1 20893
2 64506 1 20893
2 64507 1 20893
2 64508 1 20893
2 64509 1 20944
2 64510 1 20944
2 64511 1 20944
2 64512 1 20944
2 64513 1 20944
2 64514 1 20946
2 64515 1 20946
2 64516 1 20964
2 64517 1 20964
2 64518 1 20965
2 64519 1 20965
2 64520 1 21006
2 64521 1 21006
2 64522 1 21006
2 64523 1 21007
2 64524 1 21007
2 64525 1 21008
2 64526 1 21008
2 64527 1 21009
2 64528 1 21009
2 64529 1 21030
2 64530 1 21030
2 64531 1 21040
2 64532 1 21040
2 64533 1 21061
2 64534 1 21061
2 64535 1 21100
2 64536 1 21100
2 64537 1 21100
2 64538 1 21100
2 64539 1 21100
2 64540 1 21109
2 64541 1 21109
2 64542 1 21110
2 64543 1 21110
2 64544 1 21118
2 64545 1 21118
2 64546 1 21127
2 64547 1 21127
2 64548 1 21140
2 64549 1 21140
2 64550 1 21171
2 64551 1 21171
2 64552 1 21171
2 64553 1 21174
2 64554 1 21174
2 64555 1 21175
2 64556 1 21175
2 64557 1 21183
2 64558 1 21183
2 64559 1 21184
2 64560 1 21184
2 64561 1 21205
2 64562 1 21205
2 64563 1 21220
2 64564 1 21220
2 64565 1 21260
2 64566 1 21260
2 64567 1 21268
2 64568 1 21268
2 64569 1 21268
2 64570 1 21350
2 64571 1 21350
2 64572 1 21369
2 64573 1 21369
2 64574 1 21386
2 64575 1 21386
2 64576 1 21409
2 64577 1 21409
2 64578 1 21409
2 64579 1 21409
2 64580 1 21440
2 64581 1 21440
2 64582 1 21487
2 64583 1 21487
2 64584 1 21497
2 64585 1 21497
2 64586 1 21497
2 64587 1 21527
2 64588 1 21527
2 64589 1 21530
2 64590 1 21530
2 64591 1 21639
2 64592 1 21639
2 64593 1 21639
2 64594 1 21640
2 64595 1 21640
2 64596 1 21660
2 64597 1 21660
2 64598 1 21660
2 64599 1 21661
2 64600 1 21661
2 64601 1 21661
2 64602 1 21664
2 64603 1 21664
2 64604 1 21665
2 64605 1 21665
2 64606 1 21666
2 64607 1 21666
2 64608 1 21666
2 64609 1 21666
2 64610 1 21681
2 64611 1 21681
2 64612 1 21684
2 64613 1 21684
2 64614 1 21707
2 64615 1 21707
2 64616 1 21721
2 64617 1 21721
2 64618 1 21721
2 64619 1 21721
2 64620 1 21738
2 64621 1 21738
2 64622 1 21747
2 64623 1 21747
2 64624 1 21747
2 64625 1 21747
2 64626 1 21770
2 64627 1 21770
2 64628 1 21772
2 64629 1 21772
2 64630 1 21810
2 64631 1 21810
2 64632 1 21827
2 64633 1 21827
2 64634 1 21846
2 64635 1 21846
2 64636 1 21848
2 64637 1 21848
2 64638 1 21853
2 64639 1 21853
2 64640 1 21896
2 64641 1 21896
2 64642 1 21917
2 64643 1 21917
2 64644 1 21917
2 64645 1 21917
2 64646 1 21917
2 64647 1 21917
2 64648 1 21954
2 64649 1 21954
2 64650 1 21954
2 64651 1 21955
2 64652 1 21955
2 64653 1 21958
2 64654 1 21958
2 64655 1 21958
2 64656 1 21958
2 64657 1 21958
2 64658 1 21959
2 64659 1 21959
2 64660 1 21972
2 64661 1 21972
2 64662 1 21972
2 64663 1 21972
2 64664 1 21972
2 64665 1 21972
2 64666 1 21972
2 64667 1 21972
2 64668 1 21972
2 64669 1 21972
2 64670 1 21972
2 64671 1 21972
2 64672 1 21972
2 64673 1 21972
2 64674 1 21972
2 64675 1 21972
2 64676 1 21972
2 64677 1 21972
2 64678 1 21972
2 64679 1 21972
2 64680 1 21972
2 64681 1 21972
2 64682 1 21972
2 64683 1 21972
2 64684 1 21972
2 64685 1 21972
2 64686 1 21972
2 64687 1 21972
2 64688 1 21972
2 64689 1 21972
2 64690 1 21972
2 64691 1 21972
2 64692 1 21972
2 64693 1 21972
2 64694 1 21972
2 64695 1 21972
2 64696 1 21974
2 64697 1 21974
2 64698 1 21974
2 64699 1 21974
2 64700 1 21981
2 64701 1 21981
2 64702 1 21981
2 64703 1 21981
2 64704 1 21995
2 64705 1 21995
2 64706 1 22043
2 64707 1 22043
2 64708 1 22055
2 64709 1 22055
2 64710 1 22056
2 64711 1 22056
2 64712 1 22060
2 64713 1 22060
2 64714 1 22062
2 64715 1 22062
2 64716 1 22076
2 64717 1 22076
2 64718 1 22099
2 64719 1 22099
2 64720 1 22102
2 64721 1 22102
2 64722 1 22102
2 64723 1 22140
2 64724 1 22140
2 64725 1 22168
2 64726 1 22168
2 64727 1 22169
2 64728 1 22169
2 64729 1 22179
2 64730 1 22179
2 64731 1 22183
2 64732 1 22183
2 64733 1 22184
2 64734 1 22184
2 64735 1 22184
2 64736 1 22193
2 64737 1 22193
2 64738 1 22193
2 64739 1 22193
2 64740 1 22193
2 64741 1 22258
2 64742 1 22258
2 64743 1 22278
2 64744 1 22278
2 64745 1 22304
2 64746 1 22304
2 64747 1 22304
2 64748 1 22330
2 64749 1 22330
2 64750 1 22339
2 64751 1 22339
2 64752 1 22373
2 64753 1 22373
2 64754 1 22373
2 64755 1 22374
2 64756 1 22374
2 64757 1 22376
2 64758 1 22376
2 64759 1 22402
2 64760 1 22402
2 64761 1 22403
2 64762 1 22403
2 64763 1 22440
2 64764 1 22440
2 64765 1 22482
2 64766 1 22482
2 64767 1 22484
2 64768 1 22484
2 64769 1 22484
2 64770 1 22494
2 64771 1 22494
2 64772 1 22513
2 64773 1 22513
2 64774 1 22532
2 64775 1 22532
2 64776 1 22538
2 64777 1 22538
2 64778 1 22543
2 64779 1 22543
2 64780 1 22547
2 64781 1 22547
2 64782 1 22578
2 64783 1 22578
2 64784 1 22596
2 64785 1 22596
2 64786 1 22597
2 64787 1 22597
2 64788 1 22597
2 64789 1 22597
2 64790 1 22597
2 64791 1 22597
2 64792 1 22651
2 64793 1 22651
2 64794 1 22696
2 64795 1 22696
2 64796 1 22696
2 64797 1 22747
2 64798 1 22747
2 64799 1 22749
2 64800 1 22749
2 64801 1 22749
2 64802 1 22750
2 64803 1 22750
2 64804 1 22769
2 64805 1 22769
2 64806 1 22807
2 64807 1 22807
2 64808 1 22810
2 64809 1 22810
2 64810 1 22819
2 64811 1 22819
2 64812 1 22819
2 64813 1 22830
2 64814 1 22830
2 64815 1 22830
2 64816 1 22833
2 64817 1 22833
2 64818 1 22841
2 64819 1 22841
2 64820 1 22846
2 64821 1 22846
2 64822 1 22852
2 64823 1 22852
2 64824 1 22855
2 64825 1 22855
2 64826 1 22858
2 64827 1 22858
2 64828 1 22862
2 64829 1 22862
2 64830 1 22863
2 64831 1 22863
2 64832 1 22863
2 64833 1 22866
2 64834 1 22866
2 64835 1 22866
2 64836 1 22866
2 64837 1 22866
2 64838 1 22869
2 64839 1 22869
2 64840 1 22869
2 64841 1 22869
2 64842 1 22873
2 64843 1 22873
2 64844 1 22873
2 64845 1 22873
2 64846 1 22873
2 64847 1 22873
2 64848 1 22874
2 64849 1 22874
2 64850 1 22874
2 64851 1 22877
2 64852 1 22877
2 64853 1 22881
2 64854 1 22881
2 64855 1 22881
2 64856 1 22884
2 64857 1 22884
2 64858 1 22885
2 64859 1 22885
2 64860 1 22890
2 64861 1 22890
2 64862 1 22891
2 64863 1 22891
2 64864 1 22891
2 64865 1 22891
2 64866 1 22908
2 64867 1 22908
2 64868 1 22936
2 64869 1 22936
2 64870 1 22943
2 64871 1 22943
2 64872 1 22968
2 64873 1 22968
2 64874 1 22969
2 64875 1 22969
2 64876 1 22972
2 64877 1 22972
2 64878 1 22972
2 64879 1 22972
2 64880 1 22972
2 64881 1 22973
2 64882 1 22973
2 64883 1 22977
2 64884 1 22977
2 64885 1 22977
2 64886 1 22983
2 64887 1 22983
2 64888 1 22983
2 64889 1 22983
2 64890 1 22984
2 64891 1 22984
2 64892 1 22984
2 64893 1 22985
2 64894 1 22985
2 64895 1 22985
2 64896 1 22985
2 64897 1 22986
2 64898 1 22986
2 64899 1 22986
2 64900 1 22986
2 64901 1 22989
2 64902 1 22989
2 64903 1 22991
2 64904 1 22991
2 64905 1 22993
2 64906 1 22993
2 64907 1 22994
2 64908 1 22994
2 64909 1 22994
2 64910 1 22999
2 64911 1 22999
2 64912 1 23007
2 64913 1 23007
2 64914 1 23010
2 64915 1 23010
2 64916 1 23011
2 64917 1 23011
2 64918 1 23011
2 64919 1 23023
2 64920 1 23023
2 64921 1 23031
2 64922 1 23031
2 64923 1 23038
2 64924 1 23038
2 64925 1 23039
2 64926 1 23039
2 64927 1 23040
2 64928 1 23040
2 64929 1 23040
2 64930 1 23041
2 64931 1 23041
2 64932 1 23041
2 64933 1 23041
2 64934 1 23041
2 64935 1 23047
2 64936 1 23047
2 64937 1 23066
2 64938 1 23066
2 64939 1 23066
2 64940 1 23067
2 64941 1 23067
2 64942 1 23067
2 64943 1 23082
2 64944 1 23082
2 64945 1 23089
2 64946 1 23089
2 64947 1 23090
2 64948 1 23090
2 64949 1 23090
2 64950 1 23092
2 64951 1 23092
2 64952 1 23103
2 64953 1 23103
2 64954 1 23106
2 64955 1 23106
2 64956 1 23108
2 64957 1 23108
2 64958 1 23108
2 64959 1 23116
2 64960 1 23116
2 64961 1 23120
2 64962 1 23120
2 64963 1 23120
2 64964 1 23120
2 64965 1 23120
2 64966 1 23120
2 64967 1 23129
2 64968 1 23129
2 64969 1 23129
2 64970 1 23129
2 64971 1 23130
2 64972 1 23130
2 64973 1 23148
2 64974 1 23148
2 64975 1 23157
2 64976 1 23157
2 64977 1 23158
2 64978 1 23158
2 64979 1 23159
2 64980 1 23159
2 64981 1 23169
2 64982 1 23169
2 64983 1 23170
2 64984 1 23170
2 64985 1 23228
2 64986 1 23228
2 64987 1 23229
2 64988 1 23229
2 64989 1 23231
2 64990 1 23231
2 64991 1 23231
2 64992 1 23232
2 64993 1 23232
2 64994 1 23233
2 64995 1 23233
2 64996 1 23247
2 64997 1 23247
2 64998 1 23248
2 64999 1 23248
2 65000 1 23249
2 65001 1 23249
2 65002 1 23250
2 65003 1 23250
2 65004 1 23251
2 65005 1 23251
2 65006 1 23253
2 65007 1 23253
2 65008 1 23253
2 65009 1 23261
2 65010 1 23261
2 65011 1 23261
2 65012 1 23269
2 65013 1 23269
2 65014 1 23271
2 65015 1 23271
2 65016 1 23271
2 65017 1 23274
2 65018 1 23274
2 65019 1 23275
2 65020 1 23275
2 65021 1 23275
2 65022 1 23279
2 65023 1 23279
2 65024 1 23305
2 65025 1 23305
2 65026 1 23307
2 65027 1 23307
2 65028 1 23307
2 65029 1 23307
2 65030 1 23307
2 65031 1 23307
2 65032 1 23333
2 65033 1 23333
2 65034 1 23341
2 65035 1 23341
2 65036 1 23391
2 65037 1 23391
2 65038 1 23391
2 65039 1 23392
2 65040 1 23392
2 65041 1 23393
2 65042 1 23393
2 65043 1 23394
2 65044 1 23394
2 65045 1 23395
2 65046 1 23395
2 65047 1 23395
2 65048 1 23395
2 65049 1 23395
2 65050 1 23395
2 65051 1 23395
2 65052 1 23395
2 65053 1 23395
2 65054 1 23395
2 65055 1 23404
2 65056 1 23404
2 65057 1 23409
2 65058 1 23409
2 65059 1 23409
2 65060 1 23410
2 65061 1 23410
2 65062 1 23410
2 65063 1 23415
2 65064 1 23415
2 65065 1 23429
2 65066 1 23429
2 65067 1 23432
2 65068 1 23432
2 65069 1 23438
2 65070 1 23438
2 65071 1 23438
2 65072 1 23447
2 65073 1 23447
2 65074 1 23447
2 65075 1 23447
2 65076 1 23447
2 65077 1 23447
2 65078 1 23447
2 65079 1 23447
2 65080 1 23448
2 65081 1 23448
2 65082 1 23448
2 65083 1 23456
2 65084 1 23456
2 65085 1 23457
2 65086 1 23457
2 65087 1 23457
2 65088 1 23457
2 65089 1 23457
2 65090 1 23457
2 65091 1 23457
2 65092 1 23457
2 65093 1 23457
2 65094 1 23457
2 65095 1 23457
2 65096 1 23457
2 65097 1 23457
2 65098 1 23458
2 65099 1 23458
2 65100 1 23458
2 65101 1 23470
2 65102 1 23470
2 65103 1 23470
2 65104 1 23470
2 65105 1 23470
2 65106 1 23470
2 65107 1 23470
2 65108 1 23470
2 65109 1 23478
2 65110 1 23478
2 65111 1 23478
2 65112 1 23478
2 65113 1 23478
2 65114 1 23478
2 65115 1 23494
2 65116 1 23494
2 65117 1 23494
2 65118 1 23494
2 65119 1 23494
2 65120 1 23496
2 65121 1 23496
2 65122 1 23499
2 65123 1 23499
2 65124 1 23509
2 65125 1 23509
2 65126 1 23510
2 65127 1 23510
2 65128 1 23518
2 65129 1 23518
2 65130 1 23546
2 65131 1 23546
2 65132 1 23573
2 65133 1 23573
2 65134 1 23573
2 65135 1 23573
2 65136 1 23573
2 65137 1 23573
2 65138 1 23574
2 65139 1 23574
2 65140 1 23582
2 65141 1 23582
2 65142 1 23598
2 65143 1 23598
2 65144 1 23598
2 65145 1 23598
2 65146 1 23598
2 65147 1 23598
2 65148 1 23599
2 65149 1 23599
2 65150 1 23602
2 65151 1 23602
2 65152 1 23616
2 65153 1 23616
2 65154 1 23619
2 65155 1 23619
2 65156 1 23619
2 65157 1 23619
2 65158 1 23619
2 65159 1 23619
2 65160 1 23619
2 65161 1 23619
2 65162 1 23635
2 65163 1 23635
2 65164 1 23636
2 65165 1 23636
2 65166 1 23665
2 65167 1 23665
2 65168 1 23665
2 65169 1 23668
2 65170 1 23668
2 65171 1 23668
2 65172 1 23669
2 65173 1 23669
2 65174 1 23669
2 65175 1 23669
2 65176 1 23677
2 65177 1 23677
2 65178 1 23677
2 65179 1 23677
2 65180 1 23678
2 65181 1 23678
2 65182 1 23678
2 65183 1 23692
2 65184 1 23692
2 65185 1 23693
2 65186 1 23693
2 65187 1 23699
2 65188 1 23699
2 65189 1 23702
2 65190 1 23702
2 65191 1 23706
2 65192 1 23706
2 65193 1 23730
2 65194 1 23730
2 65195 1 23730
2 65196 1 23733
2 65197 1 23733
2 65198 1 23746
2 65199 1 23746
2 65200 1 23746
2 65201 1 23754
2 65202 1 23754
2 65203 1 23763
2 65204 1 23763
2 65205 1 23763
2 65206 1 23763
2 65207 1 23763
2 65208 1 23765
2 65209 1 23765
2 65210 1 23767
2 65211 1 23767
2 65212 1 23769
2 65213 1 23769
2 65214 1 23770
2 65215 1 23770
2 65216 1 23770
2 65217 1 23770
2 65218 1 23771
2 65219 1 23771
2 65220 1 23771
2 65221 1 23772
2 65222 1 23772
2 65223 1 23772
2 65224 1 23772
2 65225 1 23772
2 65226 1 23772
2 65227 1 23772
2 65228 1 23772
2 65229 1 23772
2 65230 1 23772
2 65231 1 23774
2 65232 1 23774
2 65233 1 23780
2 65234 1 23780
2 65235 1 23780
2 65236 1 23780
2 65237 1 23781
2 65238 1 23781
2 65239 1 23781
2 65240 1 23789
2 65241 1 23789
2 65242 1 23791
2 65243 1 23791
2 65244 1 23813
2 65245 1 23813
2 65246 1 23815
2 65247 1 23815
2 65248 1 23816
2 65249 1 23816
2 65250 1 23816
2 65251 1 23843
2 65252 1 23843
2 65253 1 23843
2 65254 1 23845
2 65255 1 23845
2 65256 1 23845
2 65257 1 23845
2 65258 1 23846
2 65259 1 23846
2 65260 1 23879
2 65261 1 23879
2 65262 1 23879
2 65263 1 23889
2 65264 1 23889
2 65265 1 23889
2 65266 1 23897
2 65267 1 23897
2 65268 1 23899
2 65269 1 23899
2 65270 1 23899
2 65271 1 23899
2 65272 1 23899
2 65273 1 23899
2 65274 1 23899
2 65275 1 23899
2 65276 1 23899
2 65277 1 23899
2 65278 1 23900
2 65279 1 23900
2 65280 1 23924
2 65281 1 23924
2 65282 1 23924
2 65283 1 23924
2 65284 1 23924
2 65285 1 23924
2 65286 1 23924
2 65287 1 23924
2 65288 1 23924
2 65289 1 23925
2 65290 1 23925
2 65291 1 23925
2 65292 1 23929
2 65293 1 23929
2 65294 1 23938
2 65295 1 23938
2 65296 1 23940
2 65297 1 23940
2 65298 1 23943
2 65299 1 23943
2 65300 1 23943
2 65301 1 23943
2 65302 1 23944
2 65303 1 23944
2 65304 1 23944
2 65305 1 23953
2 65306 1 23953
2 65307 1 23955
2 65308 1 23955
2 65309 1 23955
2 65310 1 23955
2 65311 1 23955
2 65312 1 23955
2 65313 1 23955
2 65314 1 23955
2 65315 1 23958
2 65316 1 23958
2 65317 1 23958
2 65318 1 23958
2 65319 1 23958
2 65320 1 23958
2 65321 1 23958
2 65322 1 23958
2 65323 1 23958
2 65324 1 23958
2 65325 1 23958
2 65326 1 23959
2 65327 1 23959
2 65328 1 23961
2 65329 1 23961
2 65330 1 23987
2 65331 1 23987
2 65332 1 24024
2 65333 1 24024
2 65334 1 24024
2 65335 1 24024
2 65336 1 24033
2 65337 1 24033
2 65338 1 24034
2 65339 1 24034
2 65340 1 24034
2 65341 1 24034
2 65342 1 24037
2 65343 1 24037
2 65344 1 24043
2 65345 1 24043
2 65346 1 24043
2 65347 1 24043
2 65348 1 24044
2 65349 1 24044
2 65350 1 24045
2 65351 1 24045
2 65352 1 24045
2 65353 1 24045
2 65354 1 24048
2 65355 1 24048
2 65356 1 24048
2 65357 1 24049
2 65358 1 24049
2 65359 1 24049
2 65360 1 24049
2 65361 1 24049
2 65362 1 24049
2 65363 1 24052
2 65364 1 24052
2 65365 1 24052
2 65366 1 24060
2 65367 1 24060
2 65368 1 24060
2 65369 1 24088
2 65370 1 24088
2 65371 1 24088
2 65372 1 24088
2 65373 1 24088
2 65374 1 24089
2 65375 1 24089
2 65376 1 24089
2 65377 1 24090
2 65378 1 24090
2 65379 1 24091
2 65380 1 24091
2 65381 1 24091
2 65382 1 24091
2 65383 1 24091
2 65384 1 24099
2 65385 1 24099
2 65386 1 24099
2 65387 1 24099
2 65388 1 24099
2 65389 1 24106
2 65390 1 24106
2 65391 1 24106
2 65392 1 24107
2 65393 1 24107
2 65394 1 24107
2 65395 1 24120
2 65396 1 24120
2 65397 1 24136
2 65398 1 24136
2 65399 1 24136
2 65400 1 24136
2 65401 1 24136
2 65402 1 24136
2 65403 1 24142
2 65404 1 24142
2 65405 1 24142
2 65406 1 24142
2 65407 1 24142
2 65408 1 24142
2 65409 1 24142
2 65410 1 24150
2 65411 1 24150
2 65412 1 24150
2 65413 1 24159
2 65414 1 24159
2 65415 1 24159
2 65416 1 24188
2 65417 1 24188
2 65418 1 24215
2 65419 1 24215
2 65420 1 24220
2 65421 1 24220
2 65422 1 24220
2 65423 1 24247
2 65424 1 24247
2 65425 1 24247
2 65426 1 24250
2 65427 1 24250
2 65428 1 24256
2 65429 1 24256
2 65430 1 24256
2 65431 1 24256
2 65432 1 24256
2 65433 1 24257
2 65434 1 24257
2 65435 1 24258
2 65436 1 24258
2 65437 1 24264
2 65438 1 24264
2 65439 1 24274
2 65440 1 24274
2 65441 1 24280
2 65442 1 24280
2 65443 1 24283
2 65444 1 24283
2 65445 1 24283
2 65446 1 24283
2 65447 1 24283
2 65448 1 24283
2 65449 1 24283
2 65450 1 24284
2 65451 1 24284
2 65452 1 24284
2 65453 1 24288
2 65454 1 24288
2 65455 1 24295
2 65456 1 24295
2 65457 1 24295
2 65458 1 24296
2 65459 1 24296
2 65460 1 24297
2 65461 1 24297
2 65462 1 24299
2 65463 1 24299
2 65464 1 24299
2 65465 1 24299
2 65466 1 24302
2 65467 1 24302
2 65468 1 24303
2 65469 1 24303
2 65470 1 24305
2 65471 1 24305
2 65472 1 24307
2 65473 1 24307
2 65474 1 24310
2 65475 1 24310
2 65476 1 24313
2 65477 1 24313
2 65478 1 24313
2 65479 1 24313
2 65480 1 24314
2 65481 1 24314
2 65482 1 24315
2 65483 1 24315
2 65484 1 24317
2 65485 1 24317
2 65486 1 24318
2 65487 1 24318
2 65488 1 24318
2 65489 1 24318
2 65490 1 24318
2 65491 1 24318
2 65492 1 24318
2 65493 1 24318
2 65494 1 24318
2 65495 1 24351
2 65496 1 24351
2 65497 1 24351
2 65498 1 24355
2 65499 1 24355
2 65500 1 24358
2 65501 1 24358
2 65502 1 24362
2 65503 1 24362
2 65504 1 24362
2 65505 1 24362
2 65506 1 24376
2 65507 1 24376
2 65508 1 24376
2 65509 1 24376
2 65510 1 24392
2 65511 1 24392
2 65512 1 24392
2 65513 1 24392
2 65514 1 24396
2 65515 1 24396
2 65516 1 24401
2 65517 1 24401
2 65518 1 24401
2 65519 1 24401
2 65520 1 24401
2 65521 1 24411
2 65522 1 24411
2 65523 1 24416
2 65524 1 24416
2 65525 1 24418
2 65526 1 24418
2 65527 1 24432
2 65528 1 24432
2 65529 1 24441
2 65530 1 24441
2 65531 1 24452
2 65532 1 24452
2 65533 1 24452
2 65534 1 24452
2 65535 1 24453
2 65536 1 24453
2 65537 1 24453
2 65538 1 24453
2 65539 1 24454
2 65540 1 24454
2 65541 1 24464
2 65542 1 24464
2 65543 1 24464
2 65544 1 24464
2 65545 1 24481
2 65546 1 24481
2 65547 1 24488
2 65548 1 24488
2 65549 1 24497
2 65550 1 24497
2 65551 1 24497
2 65552 1 24497
2 65553 1 24497
2 65554 1 24497
2 65555 1 24497
2 65556 1 24497
2 65557 1 24497
2 65558 1 24497
2 65559 1 24497
2 65560 1 24497
2 65561 1 24497
2 65562 1 24499
2 65563 1 24499
2 65564 1 24500
2 65565 1 24500
2 65566 1 24501
2 65567 1 24501
2 65568 1 24501
2 65569 1 24516
2 65570 1 24516
2 65571 1 24516
2 65572 1 24516
2 65573 1 24516
2 65574 1 24518
2 65575 1 24518
2 65576 1 24521
2 65577 1 24521
2 65578 1 24521
2 65579 1 24521
2 65580 1 24521
2 65581 1 24521
2 65582 1 24521
2 65583 1 24521
2 65584 1 24521
2 65585 1 24521
2 65586 1 24521
2 65587 1 24525
2 65588 1 24525
2 65589 1 24525
2 65590 1 24525
2 65591 1 24525
2 65592 1 24534
2 65593 1 24534
2 65594 1 24543
2 65595 1 24543
2 65596 1 24565
2 65597 1 24565
2 65598 1 24565
2 65599 1 24569
2 65600 1 24569
2 65601 1 24572
2 65602 1 24572
2 65603 1 24572
2 65604 1 24585
2 65605 1 24585
2 65606 1 24586
2 65607 1 24586
2 65608 1 24599
2 65609 1 24599
2 65610 1 24599
2 65611 1 24621
2 65612 1 24621
2 65613 1 24649
2 65614 1 24649
2 65615 1 24649
2 65616 1 24649
2 65617 1 24653
2 65618 1 24653
2 65619 1 24653
2 65620 1 24654
2 65621 1 24654
2 65622 1 24663
2 65623 1 24663
2 65624 1 24667
2 65625 1 24667
2 65626 1 24668
2 65627 1 24668
2 65628 1 24669
2 65629 1 24669
2 65630 1 24669
2 65631 1 24686
2 65632 1 24686
2 65633 1 24698
2 65634 1 24698
2 65635 1 24698
2 65636 1 24698
2 65637 1 24716
2 65638 1 24716
2 65639 1 24719
2 65640 1 24719
2 65641 1 24722
2 65642 1 24722
2 65643 1 24731
2 65644 1 24731
2 65645 1 24731
2 65646 1 24732
2 65647 1 24732
2 65648 1 24748
2 65649 1 24748
2 65650 1 24750
2 65651 1 24750
2 65652 1 24750
2 65653 1 24751
2 65654 1 24751
2 65655 1 24765
2 65656 1 24765
2 65657 1 24766
2 65658 1 24766
2 65659 1 24766
2 65660 1 24776
2 65661 1 24776
2 65662 1 24780
2 65663 1 24780
2 65664 1 24792
2 65665 1 24792
2 65666 1 24810
2 65667 1 24810
2 65668 1 24816
2 65669 1 24816
2 65670 1 24835
2 65671 1 24835
2 65672 1 24872
2 65673 1 24872
2 65674 1 24877
2 65675 1 24877
2 65676 1 24880
2 65677 1 24880
2 65678 1 24903
2 65679 1 24903
2 65680 1 24904
2 65681 1 24904
2 65682 1 24911
2 65683 1 24911
2 65684 1 24930
2 65685 1 24930
2 65686 1 24930
2 65687 1 24940
2 65688 1 24940
2 65689 1 24960
2 65690 1 24960
2 65691 1 24962
2 65692 1 24962
2 65693 1 24977
2 65694 1 24977
2 65695 1 24977
2 65696 1 24990
2 65697 1 24990
2 65698 1 25000
2 65699 1 25000
2 65700 1 25010
2 65701 1 25010
2 65702 1 25010
2 65703 1 25010
2 65704 1 25010
2 65705 1 25014
2 65706 1 25014
2 65707 1 25018
2 65708 1 25018
2 65709 1 25018
2 65710 1 25033
2 65711 1 25033
2 65712 1 25033
2 65713 1 25034
2 65714 1 25034
2 65715 1 25034
2 65716 1 25056
2 65717 1 25056
2 65718 1 25068
2 65719 1 25068
2 65720 1 25068
2 65721 1 25113
2 65722 1 25113
2 65723 1 25118
2 65724 1 25118
2 65725 1 25120
2 65726 1 25120
2 65727 1 25169
2 65728 1 25169
2 65729 1 25174
2 65730 1 25174
2 65731 1 25206
2 65732 1 25206
2 65733 1 25206
2 65734 1 25207
2 65735 1 25207
2 65736 1 25225
2 65737 1 25225
2 65738 1 25245
2 65739 1 25245
2 65740 1 25300
2 65741 1 25300
2 65742 1 25303
2 65743 1 25303
2 65744 1 25305
2 65745 1 25305
2 65746 1 25306
2 65747 1 25306
2 65748 1 25314
2 65749 1 25314
2 65750 1 25353
2 65751 1 25353
2 65752 1 25363
2 65753 1 25363
2 65754 1 25370
2 65755 1 25370
2 65756 1 25387
2 65757 1 25387
2 65758 1 25401
2 65759 1 25401
2 65760 1 25411
2 65761 1 25411
2 65762 1 25411
2 65763 1 25413
2 65764 1 25413
2 65765 1 25418
2 65766 1 25418
2 65767 1 25436
2 65768 1 25436
2 65769 1 25436
2 65770 1 25445
2 65771 1 25445
2 65772 1 25445
2 65773 1 25445
2 65774 1 25445
2 65775 1 25446
2 65776 1 25446
2 65777 1 25455
2 65778 1 25455
2 65779 1 25469
2 65780 1 25469
2 65781 1 25470
2 65782 1 25470
2 65783 1 25470
2 65784 1 25495
2 65785 1 25495
2 65786 1 25496
2 65787 1 25496
2 65788 1 25496
2 65789 1 25496
2 65790 1 25496
2 65791 1 25496
2 65792 1 25496
2 65793 1 25496
2 65794 1 25496
2 65795 1 25496
2 65796 1 25496
2 65797 1 25496
2 65798 1 25507
2 65799 1 25507
2 65800 1 25510
2 65801 1 25510
2 65802 1 25510
2 65803 1 25517
2 65804 1 25517
2 65805 1 25517
2 65806 1 25517
2 65807 1 25525
2 65808 1 25525
2 65809 1 25526
2 65810 1 25526
2 65811 1 25526
2 65812 1 25537
2 65813 1 25537
2 65814 1 25540
2 65815 1 25540
2 65816 1 25554
2 65817 1 25554
2 65818 1 25558
2 65819 1 25558
2 65820 1 25566
2 65821 1 25566
2 65822 1 25581
2 65823 1 25581
2 65824 1 25590
2 65825 1 25590
2 65826 1 25594
2 65827 1 25594
2 65828 1 25596
2 65829 1 25596
2 65830 1 25602
2 65831 1 25602
2 65832 1 25602
2 65833 1 25613
2 65834 1 25613
2 65835 1 25614
2 65836 1 25614
2 65837 1 25623
2 65838 1 25623
2 65839 1 25636
2 65840 1 25636
2 65841 1 25636
2 65842 1 25638
2 65843 1 25638
2 65844 1 25638
2 65845 1 25638
2 65846 1 25641
2 65847 1 25641
2 65848 1 25642
2 65849 1 25642
2 65850 1 25646
2 65851 1 25646
2 65852 1 25649
2 65853 1 25649
2 65854 1 25650
2 65855 1 25650
2 65856 1 25650
2 65857 1 25678
2 65858 1 25678
2 65859 1 25679
2 65860 1 25679
2 65861 1 25679
2 65862 1 25679
2 65863 1 25679
2 65864 1 25695
2 65865 1 25695
2 65866 1 25696
2 65867 1 25696
2 65868 1 25697
2 65869 1 25697
2 65870 1 25698
2 65871 1 25698
2 65872 1 25717
2 65873 1 25717
2 65874 1 25718
2 65875 1 25718
2 65876 1 25733
2 65877 1 25733
2 65878 1 25757
2 65879 1 25757
2 65880 1 25770
2 65881 1 25770
2 65882 1 25770
2 65883 1 25770
2 65884 1 25788
2 65885 1 25788
2 65886 1 25788
2 65887 1 25789
2 65888 1 25789
2 65889 1 25805
2 65890 1 25805
2 65891 1 25806
2 65892 1 25806
2 65893 1 25807
2 65894 1 25807
2 65895 1 25832
2 65896 1 25832
2 65897 1 25832
2 65898 1 25842
2 65899 1 25842
2 65900 1 25864
2 65901 1 25864
2 65902 1 25866
2 65903 1 25866
2 65904 1 25869
2 65905 1 25869
2 65906 1 25896
2 65907 1 25896
2 65908 1 25896
2 65909 1 25897
2 65910 1 25897
2 65911 1 25917
2 65912 1 25917
2 65913 1 25926
2 65914 1 25926
2 65915 1 25951
2 65916 1 25951
2 65917 1 25952
2 65918 1 25952
2 65919 1 25974
2 65920 1 25974
2 65921 1 25974
2 65922 1 25979
2 65923 1 25979
2 65924 1 25991
2 65925 1 25991
2 65926 1 26029
2 65927 1 26029
2 65928 1 26029
2 65929 1 26029
2 65930 1 26029
2 65931 1 26029
2 65932 1 26029
2 65933 1 26030
2 65934 1 26030
2 65935 1 26039
2 65936 1 26039
2 65937 1 26039
2 65938 1 26050
2 65939 1 26050
2 65940 1 26051
2 65941 1 26051
2 65942 1 26053
2 65943 1 26053
2 65944 1 26093
2 65945 1 26093
2 65946 1 26111
2 65947 1 26111
2 65948 1 26145
2 65949 1 26145
2 65950 1 26183
2 65951 1 26183
2 65952 1 26183
2 65953 1 26183
2 65954 1 26184
2 65955 1 26184
2 65956 1 26191
2 65957 1 26191
2 65958 1 26226
2 65959 1 26226
2 65960 1 26249
2 65961 1 26249
2 65962 1 26252
2 65963 1 26252
2 65964 1 26252
2 65965 1 26253
2 65966 1 26253
2 65967 1 26253
2 65968 1 26253
2 65969 1 26253
2 65970 1 26256
2 65971 1 26256
2 65972 1 26256
2 65973 1 26256
2 65974 1 26256
2 65975 1 26256
2 65976 1 26261
2 65977 1 26261
2 65978 1 26280
2 65979 1 26280
2 65980 1 26293
2 65981 1 26293
2 65982 1 26327
2 65983 1 26327
2 65984 1 26332
2 65985 1 26332
2 65986 1 26349
2 65987 1 26349
2 65988 1 26375
2 65989 1 26375
2 65990 1 26375
2 65991 1 26375
2 65992 1 26406
2 65993 1 26406
2 65994 1 26406
2 65995 1 26406
2 65996 1 26508
2 65997 1 26508
2 65998 1 26514
2 65999 1 26514
2 66000 1 26514
2 66001 1 26515
2 66002 1 26515
2 66003 1 26519
2 66004 1 26519
2 66005 1 26533
2 66006 1 26533
2 66007 1 26533
2 66008 1 26534
2 66009 1 26534
2 66010 1 26535
2 66011 1 26535
2 66012 1 26544
2 66013 1 26544
2 66014 1 26544
2 66015 1 26544
2 66016 1 26563
2 66017 1 26563
2 66018 1 26564
2 66019 1 26564
2 66020 1 26572
2 66021 1 26572
2 66022 1 26586
2 66023 1 26586
2 66024 1 26586
2 66025 1 26586
2 66026 1 26586
2 66027 1 26624
2 66028 1 26624
2 66029 1 26624
2 66030 1 26626
2 66031 1 26626
2 66032 1 26640
2 66033 1 26640
2 66034 1 26648
2 66035 1 26648
2 66036 1 26657
2 66037 1 26657
2 66038 1 26791
2 66039 1 26791
2 66040 1 26791
2 66041 1 26796
2 66042 1 26796
2 66043 1 26813
2 66044 1 26813
2 66045 1 26826
2 66046 1 26826
2 66047 1 26826
2 66048 1 26826
2 66049 1 26829
2 66050 1 26829
2 66051 1 26829
2 66052 1 26850
2 66053 1 26850
2 66054 1 26850
2 66055 1 26850
2 66056 1 26850
2 66057 1 26851
2 66058 1 26851
2 66059 1 26862
2 66060 1 26862
2 66061 1 26863
2 66062 1 26863
2 66063 1 26865
2 66064 1 26865
2 66065 1 26865
2 66066 1 26865
2 66067 1 26865
2 66068 1 26870
2 66069 1 26870
2 66070 1 26898
2 66071 1 26898
2 66072 1 26901
2 66073 1 26901
2 66074 1 26904
2 66075 1 26904
2 66076 1 26953
2 66077 1 26953
2 66078 1 26961
2 66079 1 26961
2 66080 1 26963
2 66081 1 26963
2 66082 1 26963
2 66083 1 26982
2 66084 1 26982
2 66085 1 27009
2 66086 1 27009
2 66087 1 27032
2 66088 1 27032
2 66089 1 27040
2 66090 1 27040
2 66091 1 27053
2 66092 1 27053
2 66093 1 27069
2 66094 1 27069
2 66095 1 27069
2 66096 1 27098
2 66097 1 27098
2 66098 1 27098
2 66099 1 27100
2 66100 1 27100
2 66101 1 27111
2 66102 1 27111
2 66103 1 27111
2 66104 1 27161
2 66105 1 27161
2 66106 1 27179
2 66107 1 27179
2 66108 1 27208
2 66109 1 27208
2 66110 1 27244
2 66111 1 27244
2 66112 1 27274
2 66113 1 27274
2 66114 1 27301
2 66115 1 27301
2 66116 1 27319
2 66117 1 27319
2 66118 1 27339
2 66119 1 27339
2 66120 1 27343
2 66121 1 27343
2 66122 1 27375
2 66123 1 27375
2 66124 1 27376
2 66125 1 27376
2 66126 1 27390
2 66127 1 27390
2 66128 1 27402
2 66129 1 27402
2 66130 1 27421
2 66131 1 27421
2 66132 1 27421
2 66133 1 27421
2 66134 1 27421
2 66135 1 27421
2 66136 1 27478
2 66137 1 27478
2 66138 1 27478
2 66139 1 27479
2 66140 1 27479
2 66141 1 27486
2 66142 1 27486
2 66143 1 27486
2 66144 1 27497
2 66145 1 27497
2 66146 1 27497
2 66147 1 27497
2 66148 1 27500
2 66149 1 27500
2 66150 1 27502
2 66151 1 27502
2 66152 1 27523
2 66153 1 27523
2 66154 1 27552
2 66155 1 27552
2 66156 1 27556
2 66157 1 27556
2 66158 1 27578
2 66159 1 27578
2 66160 1 27580
2 66161 1 27580
2 66162 1 27607
2 66163 1 27607
2 66164 1 27614
2 66165 1 27614
2 66166 1 27619
2 66167 1 27619
2 66168 1 27626
2 66169 1 27626
2 66170 1 27633
2 66171 1 27633
2 66172 1 27701
2 66173 1 27701
2 66174 1 27702
2 66175 1 27702
2 66176 1 27735
2 66177 1 27735
2 66178 1 27746
2 66179 1 27746
2 66180 1 27747
2 66181 1 27747
2 66182 1 27747
2 66183 1 27762
2 66184 1 27762
2 66185 1 27803
2 66186 1 27803
2 66187 1 27803
2 66188 1 27807
2 66189 1 27807
2 66190 1 27822
2 66191 1 27822
2 66192 1 27854
2 66193 1 27854
2 66194 1 27861
2 66195 1 27861
2 66196 1 27907
2 66197 1 27907
2 66198 1 27931
2 66199 1 27931
2 66200 1 27931
2 66201 1 27931
2 66202 1 27945
2 66203 1 27945
2 66204 1 27945
2 66205 1 27945
2 66206 1 27968
2 66207 1 27968
2 66208 1 28011
2 66209 1 28011
2 66210 1 28011
2 66211 1 28038
2 66212 1 28038
2 66213 1 28038
2 66214 1 28039
2 66215 1 28039
2 66216 1 28069
2 66217 1 28069
2 66218 1 28069
2 66219 1 28069
2 66220 1 28139
2 66221 1 28139
2 66222 1 28163
2 66223 1 28163
2 66224 1 28170
2 66225 1 28170
2 66226 1 28177
2 66227 1 28177
2 66228 1 28233
2 66229 1 28233
2 66230 1 28269
2 66231 1 28269
2 66232 1 28277
2 66233 1 28277
2 66234 1 28277
2 66235 1 28286
2 66236 1 28286
2 66237 1 28287
2 66238 1 28287
2 66239 1 28303
2 66240 1 28303
2 66241 1 28309
2 66242 1 28309
2 66243 1 28309
2 66244 1 28321
2 66245 1 28321
2 66246 1 28321
2 66247 1 28331
2 66248 1 28331
2 66249 1 28331
2 66250 1 28331
2 66251 1 28338
2 66252 1 28338
2 66253 1 28354
2 66254 1 28354
2 66255 1 28355
2 66256 1 28355
2 66257 1 28375
2 66258 1 28375
2 66259 1 28381
2 66260 1 28381
2 66261 1 28392
2 66262 1 28392
2 66263 1 28392
2 66264 1 28392
2 66265 1 28392
2 66266 1 28392
2 66267 1 28403
2 66268 1 28403
2 66269 1 28403
2 66270 1 28405
2 66271 1 28405
2 66272 1 28406
2 66273 1 28406
2 66274 1 28406
2 66275 1 28406
2 66276 1 28406
2 66277 1 28426
2 66278 1 28426
2 66279 1 28459
2 66280 1 28459
2 66281 1 28479
2 66282 1 28479
2 66283 1 28487
2 66284 1 28487
2 66285 1 28487
2 66286 1 28487
2 66287 1 28487
2 66288 1 28487
2 66289 1 28487
2 66290 1 28487
2 66291 1 28487
2 66292 1 28488
2 66293 1 28488
2 66294 1 28492
2 66295 1 28492
2 66296 1 28492
2 66297 1 28493
2 66298 1 28493
2 66299 1 28495
2 66300 1 28495
2 66301 1 28503
2 66302 1 28503
2 66303 1 28541
2 66304 1 28541
2 66305 1 28550
2 66306 1 28550
2 66307 1 28559
2 66308 1 28559
2 66309 1 28559
2 66310 1 28559
2 66311 1 28570
2 66312 1 28570
2 66313 1 28577
2 66314 1 28577
2 66315 1 28587
2 66316 1 28587
2 66317 1 28599
2 66318 1 28599
2 66319 1 28615
2 66320 1 28615
2 66321 1 28616
2 66322 1 28616
2 66323 1 28616
2 66324 1 28617
2 66325 1 28617
2 66326 1 28625
2 66327 1 28625
2 66328 1 28635
2 66329 1 28635
2 66330 1 28643
2 66331 1 28643
2 66332 1 28643
2 66333 1 28643
2 66334 1 28643
2 66335 1 28643
2 66336 1 28643
2 66337 1 28643
2 66338 1 28643
2 66339 1 28643
2 66340 1 28643
2 66341 1 28643
2 66342 1 28643
2 66343 1 28643
2 66344 1 28643
2 66345 1 28644
2 66346 1 28644
2 66347 1 28646
2 66348 1 28646
2 66349 1 28648
2 66350 1 28648
2 66351 1 28649
2 66352 1 28649
2 66353 1 28653
2 66354 1 28653
2 66355 1 28662
2 66356 1 28662
2 66357 1 28670
2 66358 1 28670
2 66359 1 28675
2 66360 1 28675
2 66361 1 28678
2 66362 1 28678
2 66363 1 28678
2 66364 1 28699
2 66365 1 28699
2 66366 1 28709
2 66367 1 28709
2 66368 1 28710
2 66369 1 28710
2 66370 1 28711
2 66371 1 28711
2 66372 1 28720
2 66373 1 28720
2 66374 1 28733
2 66375 1 28733
2 66376 1 28734
2 66377 1 28734
2 66378 1 28734
2 66379 1 28742
2 66380 1 28742
2 66381 1 28761
2 66382 1 28761
2 66383 1 28778
2 66384 1 28778
2 66385 1 28814
2 66386 1 28814
2 66387 1 28828
2 66388 1 28828
2 66389 1 28828
2 66390 1 28843
2 66391 1 28843
2 66392 1 28851
2 66393 1 28851
2 66394 1 28857
2 66395 1 28857
2 66396 1 28860
2 66397 1 28860
2 66398 1 28861
2 66399 1 28861
2 66400 1 28863
2 66401 1 28863
2 66402 1 28863
2 66403 1 28863
2 66404 1 28863
2 66405 1 28863
2 66406 1 28879
2 66407 1 28879
2 66408 1 28897
2 66409 1 28897
2 66410 1 28897
2 66411 1 28897
2 66412 1 28897
2 66413 1 28898
2 66414 1 28898
2 66415 1 28902
2 66416 1 28902
2 66417 1 28918
2 66418 1 28918
2 66419 1 28925
2 66420 1 28925
2 66421 1 28939
2 66422 1 28939
2 66423 1 28939
2 66424 1 28956
2 66425 1 28956
2 66426 1 28956
2 66427 1 28956
2 66428 1 28986
2 66429 1 28986
2 66430 1 28986
2 66431 1 28986
2 66432 1 28986
2 66433 1 28987
2 66434 1 28987
2 66435 1 28987
2 66436 1 28988
2 66437 1 28988
2 66438 1 29002
2 66439 1 29002
2 66440 1 29002
2 66441 1 29003
2 66442 1 29003
2 66443 1 29012
2 66444 1 29012
2 66445 1 29019
2 66446 1 29019
2 66447 1 29019
2 66448 1 29019
2 66449 1 29029
2 66450 1 29029
2 66451 1 29034
2 66452 1 29034
2 66453 1 29034
2 66454 1 29034
2 66455 1 29035
2 66456 1 29035
2 66457 1 29040
2 66458 1 29040
2 66459 1 29052
2 66460 1 29052
2 66461 1 29060
2 66462 1 29060
2 66463 1 29060
2 66464 1 29062
2 66465 1 29062
2 66466 1 29091
2 66467 1 29091
2 66468 1 29092
2 66469 1 29092
2 66470 1 29137
2 66471 1 29137
2 66472 1 29161
2 66473 1 29161
2 66474 1 29162
2 66475 1 29162
2 66476 1 29162
2 66477 1 29162
2 66478 1 29163
2 66479 1 29163
2 66480 1 29178
2 66481 1 29178
2 66482 1 29180
2 66483 1 29180
2 66484 1 29189
2 66485 1 29189
2 66486 1 29210
2 66487 1 29210
2 66488 1 29211
2 66489 1 29211
2 66490 1 29219
2 66491 1 29219
2 66492 1 29229
2 66493 1 29229
2 66494 1 29232
2 66495 1 29232
2 66496 1 29249
2 66497 1 29249
2 66498 1 29249
2 66499 1 29286
2 66500 1 29286
2 66501 1 29287
2 66502 1 29287
2 66503 1 29295
2 66504 1 29295
2 66505 1 29295
2 66506 1 29304
2 66507 1 29304
2 66508 1 29307
2 66509 1 29307
2 66510 1 29317
2 66511 1 29317
2 66512 1 29326
2 66513 1 29326
2 66514 1 29333
2 66515 1 29333
2 66516 1 29340
2 66517 1 29340
2 66518 1 29340
2 66519 1 29363
2 66520 1 29363
2 66521 1 29367
2 66522 1 29367
2 66523 1 29400
2 66524 1 29400
2 66525 1 29410
2 66526 1 29410
2 66527 1 29410
2 66528 1 29411
2 66529 1 29411
2 66530 1 29411
2 66531 1 29412
2 66532 1 29412
2 66533 1 29412
2 66534 1 29435
2 66535 1 29435
2 66536 1 29447
2 66537 1 29447
2 66538 1 29447
2 66539 1 29454
2 66540 1 29454
2 66541 1 29455
2 66542 1 29455
2 66543 1 29461
2 66544 1 29461
2 66545 1 29481
2 66546 1 29481
2 66547 1 29500
2 66548 1 29500
2 66549 1 29501
2 66550 1 29501
2 66551 1 29533
2 66552 1 29533
2 66553 1 29534
2 66554 1 29534
2 66555 1 29602
2 66556 1 29602
2 66557 1 29602
2 66558 1 29602
2 66559 1 29603
2 66560 1 29603
2 66561 1 29605
2 66562 1 29605
2 66563 1 29618
2 66564 1 29618
2 66565 1 29640
2 66566 1 29640
2 66567 1 29640
2 66568 1 29679
2 66569 1 29679
2 66570 1 29691
2 66571 1 29691
2 66572 1 29711
2 66573 1 29711
2 66574 1 29711
2 66575 1 29728
2 66576 1 29728
2 66577 1 29737
2 66578 1 29737
2 66579 1 29773
2 66580 1 29773
2 66581 1 29781
2 66582 1 29781
2 66583 1 29781
2 66584 1 29798
2 66585 1 29798
2 66586 1 29801
2 66587 1 29801
2 66588 1 29801
2 66589 1 29801
2 66590 1 29801
2 66591 1 29801
2 66592 1 29801
2 66593 1 29822
2 66594 1 29822
2 66595 1 29823
2 66596 1 29823
2 66597 1 29830
2 66598 1 29830
2 66599 1 29854
2 66600 1 29854
2 66601 1 29854
2 66602 1 29854
2 66603 1 29854
2 66604 1 29854
2 66605 1 29854
2 66606 1 29854
2 66607 1 29854
2 66608 1 29854
2 66609 1 29854
2 66610 1 29854
2 66611 1 29855
2 66612 1 29855
2 66613 1 29879
2 66614 1 29879
2 66615 1 29879
2 66616 1 29898
2 66617 1 29898
2 66618 1 29898
2 66619 1 29898
2 66620 1 29916
2 66621 1 29916
2 66622 1 29916
2 66623 1 29917
2 66624 1 29917
2 66625 1 29938
2 66626 1 29938
2 66627 1 29938
2 66628 1 29941
2 66629 1 29941
2 66630 1 29941
2 66631 1 29941
2 66632 1 29989
2 66633 1 29989
2 66634 1 30038
2 66635 1 30038
2 66636 1 30044
2 66637 1 30044
2 66638 1 30059
2 66639 1 30059
2 66640 1 30094
2 66641 1 30094
2 66642 1 30116
2 66643 1 30116
2 66644 1 30122
2 66645 1 30122
2 66646 1 30122
2 66647 1 30139
2 66648 1 30139
2 66649 1 30169
2 66650 1 30169
2 66651 1 30189
2 66652 1 30189
2 66653 1 30226
2 66654 1 30226
2 66655 1 30234
2 66656 1 30234
2 66657 1 30243
2 66658 1 30243
2 66659 1 30257
2 66660 1 30257
2 66661 1 30262
2 66662 1 30262
2 66663 1 30268
2 66664 1 30268
2 66665 1 30275
2 66666 1 30275
2 66667 1 30289
2 66668 1 30289
2 66669 1 30289
2 66670 1 30289
2 66671 1 30309
2 66672 1 30309
2 66673 1 30319
2 66674 1 30319
2 66675 1 30319
2 66676 1 30377
2 66677 1 30377
2 66678 1 30384
2 66679 1 30384
2 66680 1 30392
2 66681 1 30392
2 66682 1 30402
2 66683 1 30402
2 66684 1 30416
2 66685 1 30416
2 66686 1 30424
2 66687 1 30424
2 66688 1 30433
2 66689 1 30433
2 66690 1 30433
2 66691 1 30436
2 66692 1 30436
2 66693 1 30436
2 66694 1 30436
2 66695 1 30455
2 66696 1 30455
2 66697 1 30455
2 66698 1 30459
2 66699 1 30459
2 66700 1 30475
2 66701 1 30475
2 66702 1 30476
2 66703 1 30476
2 66704 1 30476
2 66705 1 30507
2 66706 1 30507
2 66707 1 30516
2 66708 1 30516
2 66709 1 30592
2 66710 1 30592
2 66711 1 30656
2 66712 1 30656
2 66713 1 30656
2 66714 1 30704
2 66715 1 30704
2 66716 1 30706
2 66717 1 30706
2 66718 1 30735
2 66719 1 30735
2 66720 1 30735
2 66721 1 30749
2 66722 1 30749
2 66723 1 30788
2 66724 1 30788
2 66725 1 30823
2 66726 1 30823
2 66727 1 30831
2 66728 1 30831
2 66729 1 30919
2 66730 1 30919
2 66731 1 30929
2 66732 1 30929
2 66733 1 31029
2 66734 1 31029
2 66735 1 31029
2 66736 1 31042
2 66737 1 31042
2 66738 1 31042
2 66739 1 31051
2 66740 1 31051
2 66741 1 31076
2 66742 1 31076
2 66743 1 31080
2 66744 1 31080
2 66745 1 31081
2 66746 1 31081
2 66747 1 31081
2 66748 1 31081
2 66749 1 31102
2 66750 1 31102
2 66751 1 31171
2 66752 1 31171
2 66753 1 31216
2 66754 1 31216
2 66755 1 31216
2 66756 1 31217
2 66757 1 31217
2 66758 1 31231
2 66759 1 31231
2 66760 1 31231
2 66761 1 31232
2 66762 1 31232
2 66763 1 31244
2 66764 1 31244
2 66765 1 31264
2 66766 1 31264
2 66767 1 31269
2 66768 1 31269
2 66769 1 31273
2 66770 1 31273
2 66771 1 31274
2 66772 1 31274
2 66773 1 31285
2 66774 1 31285
2 66775 1 31285
2 66776 1 31289
2 66777 1 31289
2 66778 1 31307
2 66779 1 31307
2 66780 1 31308
2 66781 1 31308
2 66782 1 31311
2 66783 1 31311
2 66784 1 31312
2 66785 1 31312
2 66786 1 31313
2 66787 1 31313
2 66788 1 31333
2 66789 1 31333
2 66790 1 31333
2 66791 1 31334
2 66792 1 31334
2 66793 1 31334
2 66794 1 31336
2 66795 1 31336
2 66796 1 31336
2 66797 1 31343
2 66798 1 31343
2 66799 1 31343
2 66800 1 31360
2 66801 1 31360
2 66802 1 31401
2 66803 1 31401
2 66804 1 31401
2 66805 1 31403
2 66806 1 31403
2 66807 1 31403
2 66808 1 31403
2 66809 1 31403
2 66810 1 31415
2 66811 1 31415
2 66812 1 31428
2 66813 1 31428
2 66814 1 31431
2 66815 1 31431
2 66816 1 31461
2 66817 1 31461
2 66818 1 31471
2 66819 1 31471
2 66820 1 31498
2 66821 1 31498
2 66822 1 31534
2 66823 1 31534
2 66824 1 31535
2 66825 1 31535
2 66826 1 31573
2 66827 1 31573
2 66828 1 31581
2 66829 1 31581
2 66830 1 31587
2 66831 1 31587
2 66832 1 31588
2 66833 1 31588
2 66834 1 31593
2 66835 1 31593
2 66836 1 31596
2 66837 1 31596
2 66838 1 31597
2 66839 1 31597
2 66840 1 31602
2 66841 1 31602
2 66842 1 31603
2 66843 1 31603
2 66844 1 31603
2 66845 1 31604
2 66846 1 31604
2 66847 1 31621
2 66848 1 31621
2 66849 1 31621
2 66850 1 31638
2 66851 1 31638
2 66852 1 31645
2 66853 1 31645
2 66854 1 31645
2 66855 1 31663
2 66856 1 31663
2 66857 1 31668
2 66858 1 31668
2 66859 1 31669
2 66860 1 31669
2 66861 1 31672
2 66862 1 31672
2 66863 1 31681
2 66864 1 31681
2 66865 1 31733
2 66866 1 31733
2 66867 1 31775
2 66868 1 31775
2 66869 1 31775
2 66870 1 31797
2 66871 1 31797
2 66872 1 31797
2 66873 1 31798
2 66874 1 31798
2 66875 1 31803
2 66876 1 31803
2 66877 1 31814
2 66878 1 31814
2 66879 1 31814
2 66880 1 31851
2 66881 1 31851
2 66882 1 31852
2 66883 1 31852
2 66884 1 31852
2 66885 1 31852
2 66886 1 31852
2 66887 1 31852
2 66888 1 31853
2 66889 1 31853
2 66890 1 31853
2 66891 1 31853
2 66892 1 31853
2 66893 1 31869
2 66894 1 31869
2 66895 1 31870
2 66896 1 31870
2 66897 1 31871
2 66898 1 31871
2 66899 1 31871
2 66900 1 31872
2 66901 1 31872
2 66902 1 31878
2 66903 1 31878
2 66904 1 31884
2 66905 1 31884
2 66906 1 31949
2 66907 1 31949
2 66908 1 31949
2 66909 1 31997
2 66910 1 31997
2 66911 1 31997
2 66912 1 32009
2 66913 1 32009
2 66914 1 32027
2 66915 1 32027
2 66916 1 32065
2 66917 1 32065
2 66918 1 32074
2 66919 1 32074
2 66920 1 32112
2 66921 1 32112
2 66922 1 32116
2 66923 1 32116
2 66924 1 32120
2 66925 1 32120
2 66926 1 32125
2 66927 1 32125
2 66928 1 32138
2 66929 1 32138
2 66930 1 32149
2 66931 1 32149
2 66932 1 32160
2 66933 1 32160
2 66934 1 32207
2 66935 1 32207
2 66936 1 32210
2 66937 1 32210
2 66938 1 32212
2 66939 1 32212
2 66940 1 32228
2 66941 1 32228
2 66942 1 32245
2 66943 1 32245
2 66944 1 32267
2 66945 1 32267
2 66946 1 32268
2 66947 1 32268
2 66948 1 32268
2 66949 1 32322
2 66950 1 32322
2 66951 1 32322
2 66952 1 32331
2 66953 1 32331
2 66954 1 32339
2 66955 1 32339
2 66956 1 32344
2 66957 1 32344
2 66958 1 32386
2 66959 1 32386
2 66960 1 32386
2 66961 1 32416
2 66962 1 32416
2 66963 1 32425
2 66964 1 32425
2 66965 1 32426
2 66966 1 32426
2 66967 1 32430
2 66968 1 32430
2 66969 1 32430
2 66970 1 32430
2 66971 1 32439
2 66972 1 32439
2 66973 1 32440
2 66974 1 32440
2 66975 1 32441
2 66976 1 32441
2 66977 1 32441
2 66978 1 32461
2 66979 1 32461
2 66980 1 32461
2 66981 1 32461
2 66982 1 32461
2 66983 1 32462
2 66984 1 32462
2 66985 1 32482
2 66986 1 32482
2 66987 1 32517
2 66988 1 32517
2 66989 1 32517
2 66990 1 32518
2 66991 1 32518
2 66992 1 32547
2 66993 1 32547
2 66994 1 32547
2 66995 1 32547
2 66996 1 32548
2 66997 1 32548
2 66998 1 32549
2 66999 1 32549
2 67000 1 32583
2 67001 1 32583
2 67002 1 32594
2 67003 1 32594
2 67004 1 32636
2 67005 1 32636
2 67006 1 32647
2 67007 1 32647
2 67008 1 32704
2 67009 1 32704
2 67010 1 32704
2 67011 1 32784
2 67012 1 32784
2 67013 1 32802
2 67014 1 32802
2 67015 1 32814
2 67016 1 32814
2 67017 1 32817
2 67018 1 32817
2 67019 1 32836
2 67020 1 32836
2 67021 1 32837
2 67022 1 32837
2 67023 1 32865
2 67024 1 32865
2 67025 1 32872
2 67026 1 32872
2 67027 1 32884
2 67028 1 32884
2 67029 1 32923
2 67030 1 32923
2 67031 1 33012
2 67032 1 33012
2 67033 1 33012
2 67034 1 33015
2 67035 1 33015
2 67036 1 33015
2 67037 1 33027
2 67038 1 33027
2 67039 1 33048
2 67040 1 33048
2 67041 1 33105
2 67042 1 33105
2 67043 1 33105
2 67044 1 33105
2 67045 1 33129
2 67046 1 33129
2 67047 1 33145
2 67048 1 33145
2 67049 1 33193
2 67050 1 33193
2 67051 1 33195
2 67052 1 33195
2 67053 1 33202
2 67054 1 33202
2 67055 1 33209
2 67056 1 33209
2 67057 1 33221
2 67058 1 33221
2 67059 1 33221
2 67060 1 33239
2 67061 1 33239
2 67062 1 33239
2 67063 1 33262
2 67064 1 33262
2 67065 1 33294
2 67066 1 33294
2 67067 1 33305
2 67068 1 33305
2 67069 1 33308
2 67070 1 33308
2 67071 1 33315
2 67072 1 33315
2 67073 1 33324
2 67074 1 33324
2 67075 1 33379
2 67076 1 33379
2 67077 1 33379
2 67078 1 33380
2 67079 1 33380
2 67080 1 33380
2 67081 1 33381
2 67082 1 33381
2 67083 1 33384
2 67084 1 33384
2 67085 1 33385
2 67086 1 33385
2 67087 1 33393
2 67088 1 33393
2 67089 1 33394
2 67090 1 33394
2 67091 1 33405
2 67092 1 33405
2 67093 1 33405
2 67094 1 33417
2 67095 1 33417
2 67096 1 33456
2 67097 1 33456
2 67098 1 33498
2 67099 1 33498
2 67100 1 33498
2 67101 1 33522
2 67102 1 33522
2 67103 1 33525
2 67104 1 33525
2 67105 1 33553
2 67106 1 33553
2 67107 1 33576
2 67108 1 33576
2 67109 1 33598
2 67110 1 33598
2 67111 1 33607
2 67112 1 33607
2 67113 1 33626
2 67114 1 33626
2 67115 1 33627
2 67116 1 33627
2 67117 1 33657
2 67118 1 33657
2 67119 1 33758
2 67120 1 33758
2 67121 1 33778
2 67122 1 33778
2 67123 1 33831
2 67124 1 33831
2 67125 1 33832
2 67126 1 33832
2 67127 1 33835
2 67128 1 33835
2 67129 1 33835
2 67130 1 33835
2 67131 1 33848
2 67132 1 33848
2 67133 1 33868
2 67134 1 33868
2 67135 1 33873
2 67136 1 33873
2 67137 1 33873
2 67138 1 33873
2 67139 1 33873
2 67140 1 33884
2 67141 1 33884
2 67142 1 33891
2 67143 1 33891
2 67144 1 33899
2 67145 1 33899
2 67146 1 33959
2 67147 1 33959
2 67148 1 33959
2 67149 1 34013
2 67150 1 34013
2 67151 1 34013
2 67152 1 34013
2 67153 1 34013
2 67154 1 34013
2 67155 1 34013
2 67156 1 34013
2 67157 1 34013
2 67158 1 34018
2 67159 1 34018
2 67160 1 34081
2 67161 1 34081
2 67162 1 34090
2 67163 1 34090
2 67164 1 34090
2 67165 1 34096
2 67166 1 34096
2 67167 1 34112
2 67168 1 34112
2 67169 1 34189
2 67170 1 34189
2 67171 1 34192
2 67172 1 34192
2 67173 1 34193
2 67174 1 34193
2 67175 1 34204
2 67176 1 34204
2 67177 1 34204
2 67178 1 34233
2 67179 1 34233
2 67180 1 34250
2 67181 1 34250
2 67182 1 34251
2 67183 1 34251
2 67184 1 34282
2 67185 1 34282
2 67186 1 34285
2 67187 1 34285
2 67188 1 34286
2 67189 1 34286
2 67190 1 34308
2 67191 1 34308
2 67192 1 34351
2 67193 1 34351
2 67194 1 34396
2 67195 1 34396
2 67196 1 34413
2 67197 1 34413
2 67198 1 34431
2 67199 1 34431
2 67200 1 34438
2 67201 1 34438
2 67202 1 34438
2 67203 1 34440
2 67204 1 34440
2 67205 1 34479
2 67206 1 34479
2 67207 1 34568
2 67208 1 34568
2 67209 1 34587
2 67210 1 34587
2 67211 1 34602
2 67212 1 34602
2 67213 1 34642
2 67214 1 34642
2 67215 1 34660
2 67216 1 34660
2 67217 1 34673
2 67218 1 34673
2 67219 1 34698
2 67220 1 34698
2 67221 1 34717
2 67222 1 34717
2 67223 1 34740
2 67224 1 34740
2 67225 1 34741
2 67226 1 34741
2 67227 1 34765
2 67228 1 34765
2 67229 1 34805
2 67230 1 34805
2 67231 1 34812
2 67232 1 34812
2 67233 1 34845
2 67234 1 34845
2 67235 1 34870
2 67236 1 34870
2 67237 1 34915
2 67238 1 34915
2 67239 1 34927
2 67240 1 34927
2 67241 1 34935
2 67242 1 34935
2 67243 1 34936
2 67244 1 34936
2 67245 1 34941
2 67246 1 34941
2 67247 1 34974
2 67248 1 34974
2 67249 1 34979
2 67250 1 34979
2 67251 1 35034
2 67252 1 35034
2 67253 1 35039
2 67254 1 35039
2 67255 1 35054
2 67256 1 35054
2 67257 1 35220
2 67258 1 35220
2 67259 1 35250
2 67260 1 35250
2 67261 1 35263
2 67262 1 35263
2 67263 1 35338
2 67264 1 35338
2 67265 1 35349
2 67266 1 35349
2 67267 1 35349
2 67268 1 35401
2 67269 1 35401
2 67270 1 35412
2 67271 1 35412
2 67272 1 35412
2 67273 1 35430
2 67274 1 35430
2 67275 1 35431
2 67276 1 35431
2 67277 1 35459
2 67278 1 35459
2 67279 1 35524
2 67280 1 35524
2 67281 1 35524
2 67282 1 35524
2 67283 1 35524
2 67284 1 35524
2 67285 1 35524
2 67286 1 35524
2 67287 1 35529
2 67288 1 35529
2 67289 1 35537
2 67290 1 35537
2 67291 1 35541
2 67292 1 35541
2 67293 1 35542
2 67294 1 35542
2 67295 1 35542
2 67296 1 35542
2 67297 1 35542
2 67298 1 35544
2 67299 1 35544
2 67300 1 35544
2 67301 1 35545
2 67302 1 35545
2 67303 1 35578
2 67304 1 35578
2 67305 1 35620
2 67306 1 35620
2 67307 1 35653
2 67308 1 35653
2 67309 1 35659
2 67310 1 35659
2 67311 1 35659
2 67312 1 35659
2 67313 1 35669
2 67314 1 35669
2 67315 1 35706
2 67316 1 35706
2 67317 1 35706
2 67318 1 35717
2 67319 1 35717
2 67320 1 35814
2 67321 1 35814
2 67322 1 35864
2 67323 1 35864
2 67324 1 35866
2 67325 1 35866
2 67326 1 35884
2 67327 1 35884
2 67328 1 35884
2 67329 1 35884
2 67330 1 35884
2 67331 1 35884
2 67332 1 35884
2 67333 1 35884
2 67334 1 35884
2 67335 1 35886
2 67336 1 35886
2 67337 1 35886
2 67338 1 35886
2 67339 1 35886
2 67340 1 35886
2 67341 1 35886
2 67342 1 35887
2 67343 1 35887
2 67344 1 35892
2 67345 1 35892
2 67346 1 35892
2 67347 1 35892
2 67348 1 35894
2 67349 1 35894
2 67350 1 35904
2 67351 1 35904
2 67352 1 35952
2 67353 1 35952
2 67354 1 35958
2 67355 1 35958
2 67356 1 35958
2 67357 1 35985
2 67358 1 35985
2 67359 1 35985
2 67360 1 35985
2 67361 1 35985
2 67362 1 35985
2 67363 1 35985
2 67364 1 35985
2 67365 1 35985
2 67366 1 35994
2 67367 1 35994
2 67368 1 35994
2 67369 1 35994
2 67370 1 35994
2 67371 1 35994
2 67372 1 35994
2 67373 1 35994
2 67374 1 35994
2 67375 1 35994
2 67376 1 35994
2 67377 1 35994
2 67378 1 35994
2 67379 1 35994
2 67380 1 35994
2 67381 1 35994
2 67382 1 35994
2 67383 1 35996
2 67384 1 35996
2 67385 1 35996
2 67386 1 36002
2 67387 1 36002
2 67388 1 36016
2 67389 1 36016
2 67390 1 36034
2 67391 1 36034
2 67392 1 36042
2 67393 1 36042
2 67394 1 36052
2 67395 1 36052
2 67396 1 36063
2 67397 1 36063
2 67398 1 36063
2 67399 1 36063
2 67400 1 36063
2 67401 1 36065
2 67402 1 36065
2 67403 1 36071
2 67404 1 36071
2 67405 1 36072
2 67406 1 36072
2 67407 1 36094
2 67408 1 36094
2 67409 1 36095
2 67410 1 36095
2 67411 1 36095
2 67412 1 36095
2 67413 1 36119
2 67414 1 36119
2 67415 1 36133
2 67416 1 36133
2 67417 1 36133
2 67418 1 36133
2 67419 1 36134
2 67420 1 36134
2 67421 1 36145
2 67422 1 36145
2 67423 1 36150
2 67424 1 36150
2 67425 1 36173
2 67426 1 36173
2 67427 1 36173
2 67428 1 36200
2 67429 1 36200
2 67430 1 36211
2 67431 1 36211
2 67432 1 36211
2 67433 1 36223
2 67434 1 36223
2 67435 1 36223
2 67436 1 36233
2 67437 1 36233
2 67438 1 36304
2 67439 1 36304
2 67440 1 36315
2 67441 1 36315
2 67442 1 36317
2 67443 1 36317
2 67444 1 36324
2 67445 1 36324
2 67446 1 36327
2 67447 1 36327
2 67448 1 36327
2 67449 1 36350
2 67450 1 36350
2 67451 1 36350
2 67452 1 36388
2 67453 1 36388
2 67454 1 36389
2 67455 1 36389
2 67456 1 36391
2 67457 1 36391
2 67458 1 36392
2 67459 1 36392
2 67460 1 36392
2 67461 1 36392
2 67462 1 36392
2 67463 1 36392
2 67464 1 36392
2 67465 1 36395
2 67466 1 36395
2 67467 1 36398
2 67468 1 36398
2 67469 1 36416
2 67470 1 36416
2 67471 1 36418
2 67472 1 36418
2 67473 1 36418
2 67474 1 36467
2 67475 1 36467
2 67476 1 36475
2 67477 1 36475
2 67478 1 36485
2 67479 1 36485
2 67480 1 36506
2 67481 1 36506
2 67482 1 36536
2 67483 1 36536
2 67484 1 36547
2 67485 1 36547
2 67486 1 36558
2 67487 1 36558
2 67488 1 36570
2 67489 1 36570
2 67490 1 36571
2 67491 1 36571
2 67492 1 36586
2 67493 1 36586
2 67494 1 36614
2 67495 1 36614
2 67496 1 36654
2 67497 1 36654
2 67498 1 36665
2 67499 1 36665
2 67500 1 36666
2 67501 1 36666
2 67502 1 36666
2 67503 1 36681
2 67504 1 36681
2 67505 1 36744
2 67506 1 36744
2 67507 1 36867
2 67508 1 36867
2 67509 1 36876
2 67510 1 36876
2 67511 1 36884
2 67512 1 36884
2 67513 1 36901
2 67514 1 36901
2 67515 1 36911
2 67516 1 36911
2 67517 1 36924
2 67518 1 36924
2 67519 1 36944
2 67520 1 36944
2 67521 1 36981
2 67522 1 36981
2 67523 1 36995
2 67524 1 36995
2 67525 1 36997
2 67526 1 36997
2 67527 1 36998
2 67528 1 36998
2 67529 1 36999
2 67530 1 36999
2 67531 1 37002
2 67532 1 37002
2 67533 1 37017
2 67534 1 37017
2 67535 1 37030
2 67536 1 37030
2 67537 1 37031
2 67538 1 37031
2 67539 1 37045
2 67540 1 37045
2 67541 1 37045
2 67542 1 37052
2 67543 1 37052
2 67544 1 37074
2 67545 1 37074
2 67546 1 37085
2 67547 1 37085
2 67548 1 37105
2 67549 1 37105
2 67550 1 37106
2 67551 1 37106
2 67552 1 37110
2 67553 1 37110
2 67554 1 37112
2 67555 1 37112
2 67556 1 37116
2 67557 1 37116
2 67558 1 37120
2 67559 1 37120
2 67560 1 37122
2 67561 1 37122
2 67562 1 37134
2 67563 1 37134
2 67564 1 37151
2 67565 1 37151
2 67566 1 37152
2 67567 1 37152
2 67568 1 37152
2 67569 1 37207
2 67570 1 37207
2 67571 1 37255
2 67572 1 37255
2 67573 1 37265
2 67574 1 37265
2 67575 1 37328
2 67576 1 37328
2 67577 1 37435
2 67578 1 37435
2 67579 1 37436
2 67580 1 37436
2 67581 1 37438
2 67582 1 37438
2 67583 1 37438
2 67584 1 37441
2 67585 1 37441
2 67586 1 37446
2 67587 1 37446
2 67588 1 37498
2 67589 1 37498
2 67590 1 37502
2 67591 1 37502
2 67592 1 37515
2 67593 1 37515
2 67594 1 37529
2 67595 1 37529
2 67596 1 37533
2 67597 1 37533
2 67598 1 37594
2 67599 1 37594
2 67600 1 37641
2 67601 1 37641
2 67602 1 37696
2 67603 1 37696
2 67604 1 37696
2 67605 1 37734
2 67606 1 37734
2 67607 1 37851
2 67608 1 37851
2 67609 1 37852
2 67610 1 37852
2 67611 1 37881
2 67612 1 37881
2 67613 1 37895
2 67614 1 37895
2 67615 1 37896
2 67616 1 37896
2 67617 1 37900
2 67618 1 37900
2 67619 1 37920
2 67620 1 37920
2 67621 1 37928
2 67622 1 37928
2 67623 1 37952
2 67624 1 37952
2 67625 1 38020
2 67626 1 38020
2 67627 1 38080
2 67628 1 38080
2 67629 1 38082
2 67630 1 38082
2 67631 1 38090
2 67632 1 38090
2 67633 1 38090
2 67634 1 38090
2 67635 1 38091
2 67636 1 38091
2 67637 1 38091
2 67638 1 38091
2 67639 1 38091
2 67640 1 38091
2 67641 1 38091
2 67642 1 38091
2 67643 1 38091
2 67644 1 38092
2 67645 1 38092
2 67646 1 38105
2 67647 1 38105
2 67648 1 38105
2 67649 1 38105
2 67650 1 38105
2 67651 1 38122
2 67652 1 38122
2 67653 1 38142
2 67654 1 38142
2 67655 1 38142
2 67656 1 38142
2 67657 1 38150
2 67658 1 38150
2 67659 1 38159
2 67660 1 38159
2 67661 1 38159
2 67662 1 38159
2 67663 1 38163
2 67664 1 38163
2 67665 1 38182
2 67666 1 38182
2 67667 1 38186
2 67668 1 38186
2 67669 1 38196
2 67670 1 38196
2 67671 1 38206
2 67672 1 38206
2 67673 1 38221
2 67674 1 38221
2 67675 1 38230
2 67676 1 38230
2 67677 1 38246
2 67678 1 38246
2 67679 1 38248
2 67680 1 38248
2 67681 1 38280
2 67682 1 38280
2 67683 1 38280
2 67684 1 38284
2 67685 1 38284
2 67686 1 38342
2 67687 1 38342
2 67688 1 38342
2 67689 1 38352
2 67690 1 38352
2 67691 1 38405
2 67692 1 38405
2 67693 1 38520
2 67694 1 38520
2 67695 1 38520
2 67696 1 38520
2 67697 1 38520
2 67698 1 38546
2 67699 1 38546
2 67700 1 38556
2 67701 1 38556
2 67702 1 38557
2 67703 1 38557
2 67704 1 38673
2 67705 1 38673
2 67706 1 38675
2 67707 1 38675
2 67708 1 38852
2 67709 1 38852
2 67710 1 38852
2 67711 1 38861
2 67712 1 38861
2 67713 1 38869
2 67714 1 38869
2 67715 1 38929
2 67716 1 38929
2 67717 1 38950
2 67718 1 38950
2 67719 1 38958
2 67720 1 38958
2 67721 1 38964
2 67722 1 38964
2 67723 1 38964
2 67724 1 38964
2 67725 1 38974
2 67726 1 38974
2 67727 1 39063
2 67728 1 39063
2 67729 1 39063
2 67730 1 39066
2 67731 1 39066
2 67732 1 39126
2 67733 1 39126
2 67734 1 39142
2 67735 1 39142
2 67736 1 39198
2 67737 1 39198
2 67738 1 39220
2 67739 1 39220
2 67740 1 39220
2 67741 1 39276
2 67742 1 39276
2 67743 1 39277
2 67744 1 39277
2 67745 1 39279
2 67746 1 39279
2 67747 1 39280
2 67748 1 39280
2 67749 1 39280
2 67750 1 39280
2 67751 1 39297
2 67752 1 39297
2 67753 1 39310
2 67754 1 39310
2 67755 1 39327
2 67756 1 39327
2 67757 1 39401
2 67758 1 39401
2 67759 1 39401
2 67760 1 39472
2 67761 1 39472
2 67762 1 39479
2 67763 1 39479
2 67764 1 39503
2 67765 1 39503
2 67766 1 39544
2 67767 1 39544
2 67768 1 39545
2 67769 1 39545
2 67770 1 39549
2 67771 1 39549
2 67772 1 39579
2 67773 1 39579
2 67774 1 39580
2 67775 1 39580
2 67776 1 39580
2 67777 1 39854
2 67778 1 39854
0 27 5 183 1 25
0 28 5 147 1 40132
0 29 5 208 1 40309
0 30 5 159 1 40542
0 31 5 173 1 40705
0 32 5 68 1 40900
0 33 5 82 1 40971
0 34 5 71 1 41038
0 35 5 79 1 41055
0 36 5 116 1 41157
0 37 5 137 1 41285
0 38 5 133 1 41409
0 39 5 143 1 41544
0 40 5 82 1 41689
0 41 5 73 1 41770
0 42 5 69 1 41824
0 43 5 156 1 41854
0 44 5 180 1 42005
0 45 5 247 1 42213
0 46 5 216 1 42450
0 47 5 173 1 42733
0 48 5 142 1 42899
0 49 5 123 1 43049
0 50 5 83 1 43166
0 51 5 10 1 43279
0 52 7 15 2 41039 45139
0 53 5 1 1 46538
0 54 7 3 2 44305 41825
0 55 5 1 1 46553
0 56 7 2 2 53 55
0 57 5 44 1 46556
0 58 7 43 2 40972 41771
0 59 5 5 1 46602
0 60 7 50 2 44841 46007
0 61 5 1 1 46650
0 62 7 25 2 44376 41855
0 63 5 47 1 46700
0 64 7 3 2 41158 46725
0 65 5 6 1 46772
0 66 7 39 2 41056 45208
0 67 5 35 1 46781
0 68 7 3 2 44455 46820
0 69 5 7 1 46855
0 70 7 2 2 26 46858
0 71 5 1 1 46865
0 72 7 7 2 46775 71
0 73 5 6 1 46867
0 74 7 2 2 40310 46874
0 75 5 2 1 46880
0 76 7 1 2 43468 46882
0 77 5 2 1 76
0 78 7 11 2 41159 45209
0 79 5 4 1 46886
0 80 7 3 2 41057 46887
0 81 5 3 1 46901
0 82 7 2 2 43615 46904
0 83 5 4 1 46907
0 84 7 1 2 39926 46909
0 85 5 2 1 84
0 86 7 7 2 44456 41856
0 87 5 2 1 46915
0 88 7 2 2 44377 46916
0 89 5 5 1 46924
0 90 7 1 2 40311 46926
0 91 5 1 1 90
0 92 7 4 2 46913 91
0 93 5 1 1 46931
0 94 7 1 2 46884 93
0 95 5 2 1 94
0 96 7 1 2 45544 46935
0 97 5 2 1 96
0 98 7 6 2 41058 41857
0 99 5 2 1 46939
0 100 7 8 2 45210 42006
0 101 5 3 1 46947
0 102 7 1 2 46945 46955
0 103 5 6 1 102
0 104 7 1 2 39927 46958
0 105 5 5 1 104
0 106 7 18 2 43616 44457
0 107 5 6 1 46969
0 108 7 1 2 42007 46987
0 109 5 1 1 108
0 110 7 1 2 46964 109
0 111 5 1 1 110
0 112 7 1 2 42214 111
0 113 5 1 1 112
0 114 7 1 2 46937 113
0 115 5 1 1 114
0 116 7 1 2 44571 115
0 117 5 1 1 116
0 118 7 34 2 41160 45364
0 119 5 35 1 46993
0 120 7 3 2 43617 47027
0 121 5 9 1 47062
0 122 7 33 2 44458 42008
0 123 5 31 1 47074
0 124 7 3 2 40312 47107
0 125 5 18 1 47138
0 126 7 1 2 46701 47141
0 127 5 2 1 126
0 128 7 1 2 47065 47159
0 129 5 1 1 128
0 130 7 1 2 43285 129
0 131 5 1 1 130
0 132 7 4 2 42009 46821
0 133 5 5 1 47161
0 134 7 2 2 47165 46859
0 135 7 1 2 47108 47170
0 136 5 2 1 135
0 137 7 1 2 43618 47172
0 138 5 1 1 137
0 139 7 1 2 131 138
0 140 5 1 1 139
0 141 7 1 2 43469 140
0 142 5 1 1 141
0 143 7 1 2 42010 46856
0 144 5 1 1 143
0 145 7 1 2 39928 144
0 146 5 1 1 145
0 147 7 3 2 42011 46776
0 148 5 1 1 47174
0 149 7 9 2 44378 44459
0 150 5 5 1 47177
0 151 7 5 2 41858 47178
0 152 5 1 1 47191
0 153 7 2 2 148 152
0 154 5 3 1 47196
0 155 7 3 2 146 47198
0 156 5 4 1 47201
0 157 7 1 2 43619 47202
0 158 5 1 1 157
0 159 7 1 2 142 158
0 160 5 1 1 159
0 161 7 1 2 45545 160
0 162 5 1 1 161
0 163 7 1 2 117 162
0 164 5 1 1 163
0 165 7 1 2 46651 164
0 166 5 1 1 165
0 167 7 31 2 41545 42734
0 168 5 9 1 47208
0 169 7 2 2 43470 47142
0 170 5 1 1 47248
0 171 7 2 2 47066 170
0 172 5 4 1 47250
0 173 7 2 2 45546 47252
0 174 5 1 1 47256
0 175 7 47 2 39929 41059
0 176 5 66 1 47258
0 177 7 71 2 43286 44379
0 178 5 69 1 47371
0 179 7 15 2 45211 47442
0 180 5 12 1 47511
0 181 7 5 2 47305 47526
0 182 5 19 1 47538
0 183 7 2 2 40133 47109
0 184 5 6 1 47562
0 185 7 1 2 47063 47564
0 186 5 4 1 185
0 187 7 1 2 47543 47570
0 188 5 1 1 187
0 189 7 1 2 47257 188
0 190 5 1 1 189
0 191 7 30 2 40134 41161
0 192 5 87 1 47574
0 193 7 59 2 43471 44460
0 194 5 82 1 47691
0 195 7 1 2 47750 47544
0 196 5 3 1 195
0 197 7 4 2 47604 47832
0 198 5 1 1 47835
0 199 7 1 2 45547 47836
0 200 5 2 1 199
0 201 7 2 2 42215 46988
0 202 5 1 1 47841
0 203 7 1 2 47839 202
0 204 5 1 1 203
0 205 7 1 2 44572 204
0 206 5 1 1 205
0 207 7 1 2 190 206
0 208 5 1 1 207
0 209 7 1 2 47209 208
0 210 5 1 1 209
0 211 7 1 2 166 210
0 212 5 1 1 211
0 213 7 1 2 44708 212
0 214 5 1 1 213
0 215 7 11 2 41859 42735
0 216 5 1 1 47843
0 217 7 8 2 44380 41546
0 218 7 1 2 47844 47854
0 219 5 2 1 218
0 220 7 3 2 44381 47210
0 221 5 1 1 47864
0 222 7 1 2 45212 221
0 223 5 1 1 222
0 224 7 1 2 44382 46652
0 225 5 1 1 224
0 226 7 1 2 47239 225
0 227 5 3 1 226
0 228 7 1 2 43287 47867
0 229 7 1 2 223 228
0 230 5 1 1 229
0 231 7 1 2 47862 230
0 232 5 1 1 231
0 233 7 11 2 43620 45548
0 234 5 1 1 47870
0 235 7 4 2 43472 44573
0 236 7 3 2 47075 47881
0 237 5 1 1 47885
0 238 7 1 2 47871 47886
0 239 7 1 2 232 238
0 240 5 1 1 239
0 241 7 1 2 214 240
0 242 5 1 1 241
0 243 7 1 2 43982 242
0 244 5 1 1 243
0 245 7 1 2 43288 46822
0 246 5 7 1 245
0 247 7 6 2 46726 47888
0 248 5 24 1 47895
0 249 7 2 2 43621 47901
0 250 5 1 1 47925
0 251 7 11 2 44461 44574
0 252 5 3 1 47927
0 253 7 4 2 45549 47928
0 254 5 1 1 47941
0 255 7 7 2 43473 40706
0 256 7 10 2 42012 42736
0 257 7 1 2 44842 47952
0 258 7 1 2 47945 257
0 259 7 1 2 47942 258
0 260 7 1 2 47926 259
0 261 5 1 1 260
0 262 7 1 2 244 261
0 263 5 1 1 262
0 264 7 1 2 46180 263
0 265 5 1 1 264
0 266 7 17 2 45213 42216
0 267 5 2 1 47962
0 268 7 2 2 47372 47963
0 269 5 1 1 47981
0 270 7 3 2 44575 47028
0 271 5 13 1 47983
0 272 7 3 2 41286 47110
0 273 5 10 1 47999
0 274 7 1 2 43474 48002
0 275 5 2 1 274
0 276 7 2 2 47986 48012
0 277 5 2 1 48014
0 278 7 1 2 47982 48016
0 279 5 1 1 278
0 280 7 3 2 45550 47539
0 281 7 1 2 47887 48018
0 282 5 1 1 281
0 283 7 1 2 279 282
0 284 5 1 1 283
0 285 7 1 2 43622 284
0 286 5 1 1 285
0 287 7 5 2 42217 46948
0 288 7 6 2 44383 44576
0 289 5 2 1 48026
0 290 7 3 2 43289 48027
0 291 5 2 1 48034
0 292 7 2 2 47692 48035
0 293 7 1 2 48021 48039
0 294 5 2 1 293
0 295 7 1 2 286 48041
0 296 5 2 1 295
0 297 7 42 2 40707 41547
0 298 5 2 1 48045
0 299 7 47 2 46008 42900
0 300 7 4 2 48046 48089
0 301 7 1 2 48043 48136
0 302 5 1 1 301
0 303 7 1 2 265 302
0 304 5 1 1 303
0 305 7 1 2 43823 304
0 306 5 1 1 305
0 307 7 6 2 40708 48090
0 308 5 2 1 48140
0 309 7 2 2 47964 47855
0 310 7 1 2 48141 48148
0 311 5 1 1 310
0 312 7 22 2 42013 45551
0 313 5 6 1 48150
0 314 7 4 2 44462 48151
0 315 5 4 1 48178
0 316 7 7 2 41548 48091
0 317 5 4 1 48186
0 318 7 50 2 42737 46181
0 319 7 10 2 44843 48197
0 320 5 1 1 48247
0 321 7 1 2 48193 320
0 322 5 34 1 321
0 323 7 1 2 40709 48257
0 324 5 2 1 323
0 325 7 7 2 43983 48198
0 326 5 1 1 48293
0 327 7 1 2 41549 48294
0 328 5 1 1 327
0 329 7 1 2 48291 328
0 330 5 9 1 329
0 331 7 1 2 46823 48300
0 332 5 1 1 331
0 333 7 7 2 43984 44384
0 334 5 1 1 48309
0 335 7 4 2 44844 48310
0 336 7 10 2 41860 46182
0 337 7 1 2 46009 48320
0 338 7 1 2 48316 337
0 339 5 1 1 338
0 340 7 1 2 332 339
0 341 5 1 1 340
0 342 7 1 2 48179 341
0 343 5 1 1 342
0 344 7 1 2 311 343
0 345 5 1 1 344
0 346 7 1 2 43475 345
0 347 5 1 1 346
0 348 7 17 2 42218 46010
0 349 7 3 2 42901 48330
0 350 7 4 2 40710 44385
0 351 7 10 2 41550 45214
0 352 7 1 2 47029 48354
0 353 7 1 2 48350 352
0 354 7 1 2 48347 353
0 355 5 1 1 354
0 356 7 1 2 347 355
0 357 5 1 1 356
0 358 7 1 2 43290 357
0 359 5 1 1 358
0 360 7 16 2 43476 44386
0 361 5 5 1 48364
0 362 7 9 2 41861 48365
0 363 5 2 1 48385
0 364 7 1 2 48386 48180
0 365 7 1 2 48301 364
0 366 5 1 1 365
0 367 7 1 2 359 366
0 368 5 1 1 367
0 369 7 1 2 44577 368
0 370 5 1 1 369
0 371 7 11 2 41551 42902
0 372 7 2 2 48331 48396
0 373 7 2 2 46949 48407
0 374 7 3 2 43291 47693
0 375 5 3 1 48411
0 376 7 2 2 48351 48412
0 377 7 1 2 48409 48417
0 378 5 1 1 377
0 379 7 1 2 370 378
0 380 5 1 1 379
0 381 7 1 2 43623 380
0 382 5 1 1 381
0 383 7 4 2 44387 47929
0 384 5 2 1 48419
0 385 7 1 2 43292 47946
0 386 7 1 2 48420 385
0 387 7 1 2 48410 386
0 388 5 1 1 387
0 389 7 1 2 382 388
0 390 5 1 1 389
0 391 7 1 2 44709 390
0 392 5 1 1 391
0 393 7 1 2 306 392
0 394 5 1 1 393
0 395 7 1 2 44984 394
0 396 5 1 1 395
0 397 7 22 2 40711 44845
0 398 5 2 1 48425
0 399 7 2 2 41690 48426
0 400 7 78 2 40543 41410
0 401 5 37 1 48451
0 402 7 30 2 42738 42903
0 403 7 1 2 48529 48566
0 404 7 2 2 48044 403
0 405 7 1 2 48449 48596
0 406 5 1 1 405
0 407 7 1 2 396 406
0 408 5 1 1 407
0 409 7 1 2 44155 408
0 410 5 1 1 409
0 411 7 9 2 43985 44710
0 412 5 1 1 48598
0 413 7 13 2 43293 43477
0 414 5 22 1 48607
0 415 7 70 2 40313 41287
0 416 5 63 1 48642
0 417 7 10 2 41162 45552
0 418 5 4 1 48775
0 419 7 2 2 48643 48776
0 420 7 2 2 48620 48789
0 421 7 1 2 48599 48791
0 422 5 1 1 421
0 423 7 3 2 41862 47605
0 424 5 2 1 48793
0 425 7 1 2 47306 48794
0 426 5 1 1 425
0 427 7 1 2 47751 426
0 428 5 5 1 427
0 429 7 40 2 44578 42219
0 430 5 22 1 48803
0 431 7 6 2 43624 48804
0 432 5 9 1 48865
0 433 7 5 2 40712 48530
0 434 5 1 1 48880
0 435 7 1 2 48866 48881
0 436 7 1 2 48798 435
0 437 5 1 1 436
0 438 7 1 2 422 437
0 439 5 1 1 438
0 440 7 64 2 44156 44985
0 441 5 2 1 48885
0 442 7 21 2 44846 42739
0 443 5 2 1 48951
0 444 7 1 2 48949 48972
0 445 5 1 1 444
0 446 7 6 2 44157 41691
0 447 5 1 1 48974
0 448 7 9 2 40901 44986
0 449 5 1 1 48980
0 450 7 2 2 447 449
0 451 5 77 1 48989
0 452 7 29 2 41552 46011
0 453 5 2 1 49068
0 454 7 1 2 48990 49097
0 455 5 1 1 454
0 456 7 1 2 445 455
0 457 7 1 2 439 456
0 458 5 1 1 457
0 459 7 2 2 44987 48792
0 460 7 23 2 40713 44158
0 461 7 8 2 48452 49101
0 462 5 1 1 49124
0 463 7 1 2 48952 49125
0 464 7 1 2 49099 463
0 465 5 1 1 464
0 466 7 1 2 458 465
0 467 5 1 1 466
0 468 7 1 2 42904 467
0 469 5 1 1 468
0 470 7 6 2 43824 44847
0 471 7 3 2 46012 49132
0 472 7 6 2 48600 49138
0 473 5 1 1 49141
0 474 7 5 2 44579 48531
0 475 5 1 1 49147
0 476 7 3 2 43294 47606
0 477 5 3 1 49152
0 478 7 11 2 43986 41553
0 479 5 1 1 49158
0 480 7 5 2 48447 479
0 481 5 65 1 49169
0 482 7 16 2 42740 49174
0 483 5 1 1 49239
0 484 7 1 2 49153 49240
0 485 5 1 1 484
0 486 7 3 2 43478 43987
0 487 7 3 2 44463 46653
0 488 5 1 1 49258
0 489 7 1 2 49255 49259
0 490 5 1 1 489
0 491 7 1 2 485 490
0 492 5 1 1 491
0 493 7 1 2 49148 492
0 494 5 1 1 493
0 495 7 1 2 473 494
0 496 5 1 1 495
0 497 7 1 2 43625 496
0 498 5 1 1 497
0 499 7 11 2 43825 43988
0 500 5 1 1 49261
0 501 7 14 2 44711 49262
0 502 7 1 2 47694 46654
0 503 5 2 1 502
0 504 7 3 2 43295 47211
0 505 5 1 1 49288
0 506 7 1 2 47607 49289
0 507 5 1 1 506
0 508 7 1 2 49286 507
0 509 5 1 1 508
0 510 7 1 2 49272 509
0 511 5 1 1 510
0 512 7 1 2 498 511
0 513 5 1 1 512
0 514 7 1 2 46824 513
0 515 5 1 1 514
0 516 7 5 2 39930 47575
0 517 5 4 1 49291
0 518 7 2 2 49296 48712
0 519 5 2 1 49300
0 520 7 6 2 40314 41060
0 521 5 2 1 49304
0 522 7 1 2 44580 49310
0 523 5 1 1 522
0 524 7 1 2 49302 523
0 525 5 1 1 524
0 526 7 1 2 49142 525
0 527 5 1 1 526
0 528 7 6 2 40135 46727
0 529 5 8 1 49312
0 530 7 3 2 49318 46777
0 531 5 1 1 49326
0 532 7 7 2 47608 49327
0 533 5 1 1 49329
0 534 7 2 2 43296 46655
0 535 5 1 1 49336
0 536 7 1 2 47240 535
0 537 5 3 1 536
0 538 7 1 2 49273 49338
0 539 5 1 1 538
0 540 7 3 2 40714 48953
0 541 5 4 1 49341
0 542 7 1 2 43989 49339
0 543 5 1 1 542
0 544 7 1 2 49344 543
0 545 5 1 1 544
0 546 7 2 2 43626 545
0 547 5 1 1 49348
0 548 7 1 2 49349 49149
0 549 5 1 1 548
0 550 7 1 2 539 549
0 551 5 1 1 550
0 552 7 1 2 49330 551
0 553 5 1 1 552
0 554 7 1 2 527 553
0 555 7 1 2 515 554
0 556 5 1 1 555
0 557 7 10 2 46183 48886
0 558 7 1 2 42220 49350
0 559 7 1 2 556 558
0 560 5 1 1 559
0 561 7 1 2 469 560
0 562 5 1 1 561
0 563 7 1 2 45365 562
0 564 5 1 1 563
0 565 7 7 2 44848 44988
0 566 7 11 2 40715 40902
0 567 5 1 1 49367
0 568 7 1 2 49360 49368
0 569 7 1 2 48597 568
0 570 5 1 1 569
0 571 7 1 2 45791 570
0 572 7 1 2 564 571
0 573 7 1 2 410 572
0 574 5 1 1 573
0 575 7 4 2 41411 41863
0 576 7 6 2 43297 44464
0 577 5 1 1 49382
0 578 7 68 2 43627 44581
0 579 5 89 1 49388
0 580 7 4 2 49383 49389
0 581 5 1 1 49545
0 582 7 3 2 48366 49546
0 583 7 1 2 49378 49549
0 584 5 1 1 583
0 585 7 71 2 43826 44712
0 586 5 55 1 49552
0 587 7 11 2 40136 47443
0 588 5 8 1 49678
0 589 7 2 2 49679 46888
0 590 5 2 1 49697
0 591 7 2 2 48713 49699
0 592 5 1 1 49701
0 593 7 2 2 41163 49456
0 594 5 2 1 49703
0 595 7 9 2 39931 45215
0 596 5 9 1 49707
0 597 7 1 2 49708 49457
0 598 5 2 1 597
0 599 7 1 2 49705 49725
0 600 7 1 2 49702 599
0 601 5 1 1 600
0 602 7 1 2 49553 601
0 603 5 1 1 602
0 604 7 1 2 584 603
0 605 5 1 1 604
0 606 7 1 2 46656 605
0 607 5 1 1 606
0 608 7 7 2 44582 41412
0 609 7 3 2 46970 49727
0 610 7 3 2 43479 49734
0 611 7 2 2 41554 49737
0 612 5 1 1 49740
0 613 7 4 2 42741 47902
0 614 7 1 2 49741 49742
0 615 5 1 1 614
0 616 7 1 2 607 615
0 617 5 1 1 616
0 618 7 1 2 45553 617
0 619 5 1 1 618
0 620 7 10 2 43628 43827
0 621 5 2 1 49746
0 622 7 9 2 43480 47373
0 623 5 15 1 49758
0 624 7 4 2 49747 49759
0 625 7 7 2 44583 44713
0 626 7 2 2 44465 49786
0 627 7 1 2 41864 49069
0 628 7 1 2 49793 627
0 629 7 1 2 49782 628
0 630 5 1 1 629
0 631 7 1 2 619 630
0 632 5 1 1 631
0 633 7 1 2 44989 632
0 634 5 1 1 633
0 635 7 22 2 43481 43629
0 636 5 4 1 49795
0 637 7 8 2 44466 49796
0 638 5 3 1 49821
0 639 7 11 2 43828 44584
0 640 7 3 2 49822 49832
0 641 7 11 2 44849 41692
0 642 7 2 2 44714 49846
0 643 5 1 1 49857
0 644 7 1 2 49843 49858
0 645 7 1 2 49743 644
0 646 5 1 1 645
0 647 7 1 2 634 646
0 648 5 1 1 647
0 649 7 1 2 46184 648
0 650 5 1 1 649
0 651 7 10 2 40315 47752
0 652 5 41 1 49859
0 653 7 2 2 41288 47753
0 654 5 6 1 49910
0 655 7 5 2 49869 49912
0 656 5 4 1 49918
0 657 7 15 2 48714 49919
0 658 5 1 1 49927
0 659 7 5 2 39932 46728
0 660 5 8 1 49942
0 661 7 6 2 46825 49947
0 662 5 1 1 49955
0 663 7 7 2 43829 46013
0 664 7 22 2 44990 46185
0 665 5 1 1 49968
0 666 7 23 2 41693 42905
0 667 5 4 1 49990
0 668 7 1 2 665 50013
0 669 5 9 1 668
0 670 7 1 2 49961 50017
0 671 7 1 2 49956 670
0 672 7 1 2 49928 671
0 673 5 1 1 672
0 674 7 10 2 41061 41289
0 675 7 2 2 40316 50026
0 676 5 1 1 50036
0 677 7 3 2 47374 48715
0 678 5 5 1 50038
0 679 7 3 2 43482 48716
0 680 5 2 1 50046
0 681 7 2 2 50041 50049
0 682 7 1 2 49704 50051
0 683 5 1 1 682
0 684 7 1 2 676 683
0 685 5 1 1 684
0 686 7 10 2 41865 42906
0 687 7 13 2 41694 42742
0 688 7 1 2 50053 50063
0 689 7 1 2 685 688
0 690 5 1 1 689
0 691 7 1 2 673 690
0 692 5 1 1 691
0 693 7 1 2 41555 692
0 694 5 1 1 693
0 695 7 2 2 47540 49929
0 696 5 1 1 50076
0 697 7 3 2 48199 49847
0 698 5 1 1 50078
0 699 7 1 2 43830 50079
0 700 7 1 2 50077 699
0 701 5 1 1 700
0 702 7 1 2 694 701
0 703 5 1 1 702
0 704 7 1 2 44715 703
0 705 5 1 1 704
0 706 7 2 2 49920 50039
0 707 5 1 1 50081
0 708 7 8 2 41413 44991
0 709 7 3 2 46186 50083
0 710 7 6 2 40544 44850
0 711 7 2 2 46014 50094
0 712 5 1 1 50100
0 713 7 9 2 45216 42743
0 714 7 3 2 41556 50102
0 715 5 1 1 50111
0 716 7 1 2 712 715
0 717 5 1 1 716
0 718 7 1 2 50091 717
0 719 7 1 2 50082 718
0 720 5 1 1 719
0 721 7 1 2 705 720
0 722 5 1 1 721
0 723 7 1 2 42221 722
0 724 5 1 1 723
0 725 7 2 2 48092 47903
0 726 7 6 2 43483 43831
0 727 7 3 2 50116 46971
0 728 7 13 2 44585 41557
0 729 7 3 2 44716 41695
0 730 7 1 2 50125 50138
0 731 7 1 2 50122 730
0 732 7 1 2 50114 731
0 733 5 1 1 732
0 734 7 1 2 724 733
0 735 7 1 2 650 734
0 736 5 1 1 735
0 737 7 1 2 42014 736
0 738 5 1 1 737
0 739 7 9 2 41290 44851
0 740 7 6 2 39933 46940
0 741 5 1 1 50150
0 742 7 7 2 43630 45366
0 743 5 6 1 50156
0 744 7 1 2 741 50163
0 745 5 2 1 744
0 746 7 1 2 45554 50169
0 747 5 2 1 746
0 748 7 15 2 40317 41164
0 749 5 2 1 50173
0 750 7 7 2 43631 47609
0 751 5 22 1 50190
0 752 7 1 2 39934 50197
0 753 5 2 1 752
0 754 7 14 2 41062 41165
0 755 5 7 1 50221
0 756 7 5 2 40137 50222
0 757 5 3 1 50242
0 758 7 1 2 50219 50247
0 759 5 1 1 758
0 760 7 1 2 45217 759
0 761 5 1 1 760
0 762 7 1 2 50188 761
0 763 5 3 1 762
0 764 7 1 2 42222 50250
0 765 5 1 1 764
0 766 7 1 2 50171 765
0 767 5 1 1 766
0 768 7 1 2 50141 767
0 769 5 1 1 768
0 770 7 5 2 44586 49797
0 771 7 8 2 41558 42223
0 772 5 2 1 50258
0 773 7 2 2 44467 50259
0 774 7 1 2 50253 50268
0 775 5 1 1 774
0 776 7 24 2 41291 45367
0 777 5 2 1 50270
0 778 7 6 2 45555 50271
0 779 7 1 2 44852 50296
0 780 5 1 1 779
0 781 7 1 2 775 780
0 782 5 1 1 781
0 783 7 1 2 47307 782
0 784 5 1 1 783
0 785 7 7 2 43484 46972
0 786 5 6 1 50302
0 787 7 21 2 41866 42224
0 788 5 5 1 50315
0 789 7 1 2 50316 50126
0 790 7 1 2 50303 789
0 791 5 1 1 790
0 792 7 1 2 784 791
0 793 7 1 2 769 792
0 794 5 1 1 793
0 795 7 1 2 49554 794
0 796 5 1 1 795
0 797 7 7 2 43632 42225
0 798 5 11 1 50341
0 799 7 5 2 43485 47930
0 800 5 1 1 50359
0 801 7 2 2 50342 50360
0 802 5 1 1 50364
0 803 7 11 2 39935 46782
0 804 5 14 1 50366
0 805 7 13 2 41414 44853
0 806 7 2 2 50377 50391
0 807 7 1 2 45368 50404
0 808 7 1 2 50365 807
0 809 5 1 1 808
0 810 7 1 2 46015 809
0 811 7 1 2 796 810
0 812 5 1 1 811
0 813 7 5 2 41559 49555
0 814 5 2 1 50406
0 815 7 10 2 40318 45556
0 816 5 4 1 50413
0 817 7 21 2 45218 45369
0 818 5 13 1 50427
0 819 7 2 2 41166 50428
0 820 5 2 1 50461
0 821 7 1 2 50423 50463
0 822 5 3 1 821
0 823 7 1 2 50407 50465
0 824 5 1 1 823
0 825 7 21 2 45370 45557
0 826 5 3 1 50468
0 827 7 4 2 41167 50469
0 828 5 5 1 50492
0 829 7 2 2 42226 47030
0 830 5 18 1 50501
0 831 7 5 2 40138 50503
0 832 5 4 1 50521
0 833 7 1 2 48785 50526
0 834 5 1 1 833
0 835 7 1 2 49709 834
0 836 5 1 1 835
0 837 7 1 2 50496 836
0 838 5 1 1 837
0 839 7 1 2 41063 838
0 840 5 1 1 839
0 841 7 4 2 40139 46889
0 842 5 2 1 50530
0 843 7 1 2 45558 50531
0 844 5 1 1 843
0 845 7 1 2 840 844
0 846 5 1 1 845
0 847 7 6 2 40319 44854
0 848 7 1 2 49623 50536
0 849 7 1 2 846 848
0 850 5 1 1 849
0 851 7 1 2 824 850
0 852 5 1 1 851
0 853 7 1 2 41292 852
0 854 5 1 1 853
0 855 7 2 2 43832 41168
0 856 5 1 1 50542
0 857 7 4 2 44717 50543
0 858 7 7 2 43486 47308
0 859 5 10 1 50548
0 860 7 4 2 45219 50555
0 861 5 2 1 50565
0 862 7 3 2 45559 50566
0 863 5 1 1 50571
0 864 7 1 2 50544 50572
0 865 5 1 1 864
0 866 7 26 2 45371 42227
0 867 5 8 1 50574
0 868 7 2 2 43487 50575
0 869 5 2 1 50608
0 870 7 1 2 50609 49735
0 871 5 1 1 870
0 872 7 1 2 865 871
0 873 5 1 1 872
0 874 7 1 2 41560 873
0 875 5 1 1 874
0 876 7 1 2 42744 875
0 877 7 1 2 854 876
0 878 5 1 1 877
0 879 7 1 2 44992 878
0 880 7 1 2 812 879
0 881 5 1 1 880
0 882 7 4 2 41696 42228
0 883 7 10 2 44718 42745
0 884 7 2 2 50612 50616
0 885 5 1 1 50626
0 886 7 1 2 44855 50627
0 887 7 1 2 49844 886
0 888 5 1 1 887
0 889 7 1 2 881 888
0 890 5 1 1 889
0 891 7 1 2 46187 890
0 892 5 1 1 891
0 893 7 6 2 46188 49556
0 894 5 1 1 50628
0 895 7 11 2 41561 44993
0 896 7 2 2 50629 50634
0 897 5 1 1 50645
0 898 7 10 2 45560 49624
0 899 7 1 2 50018 50142
0 900 7 1 2 50647 899
0 901 5 1 1 900
0 902 7 1 2 897 901
0 903 5 1 1 902
0 904 7 1 2 46994 903
0 905 5 1 1 904
0 906 7 9 2 43833 45561
0 907 5 3 1 50657
0 908 7 8 2 41293 42229
0 909 5 8 1 50669
0 910 7 22 2 41867 42015
0 911 5 16 1 50685
0 912 7 2 2 50670 50686
0 913 5 1 1 50723
0 914 7 2 2 50666 913
0 915 5 1 1 50725
0 916 7 14 2 44719 41562
0 917 5 1 1 50727
0 918 7 1 2 49991 50728
0 919 7 1 2 915 918
0 920 5 1 1 919
0 921 7 1 2 905 920
0 922 5 1 1 921
0 923 7 1 2 42746 922
0 924 5 1 1 923
0 925 7 2 2 42907 49625
0 926 7 12 2 41294 44994
0 927 5 1 1 50743
0 928 7 1 2 45372 50744
0 929 7 13 2 45562 46016
0 930 7 5 2 41169 41563
0 931 7 1 2 50755 50768
0 932 7 1 2 928 931
0 933 7 1 2 50741 932
0 934 5 1 1 933
0 935 7 1 2 924 934
0 936 5 1 1 935
0 937 7 1 2 40320 936
0 938 5 1 1 937
0 939 7 8 2 43834 41295
0 940 7 7 2 46189 50617
0 941 5 1 1 50781
0 942 7 2 2 50773 50782
0 943 5 1 1 50788
0 944 7 10 2 41564 45563
0 945 7 2 2 44995 50790
0 946 7 1 2 50789 50800
0 947 5 1 1 946
0 948 7 1 2 938 947
0 949 5 1 1 948
0 950 7 1 2 48621 949
0 951 5 1 1 950
0 952 7 17 2 46017 49557
0 953 5 2 1 50802
0 954 7 5 2 43298 41868
0 955 5 3 1 50821
0 956 7 11 2 44388 50822
0 957 5 15 1 50829
0 958 7 1 2 45373 50840
0 959 5 3 1 958
0 960 7 1 2 50855 49969
0 961 5 1 1 960
0 962 7 1 2 45374 47896
0 963 5 5 1 962
0 964 7 1 2 49992 50858
0 965 5 1 1 964
0 966 7 1 2 961 965
0 967 5 1 1 966
0 968 7 1 2 50803 967
0 969 5 1 1 968
0 970 7 7 2 41415 42747
0 971 7 14 2 41869 45375
0 972 5 3 1 50870
0 973 7 8 2 44389 45220
0 974 5 4 1 50887
0 975 7 1 2 50884 50895
0 976 5 6 1 975
0 977 7 3 2 49948 50899
0 978 7 1 2 50905 49970
0 979 5 1 1 978
0 980 7 5 2 42016 42908
0 981 7 2 2 41697 50908
0 982 5 1 1 50913
0 983 7 1 2 45221 50914
0 984 5 1 1 983
0 985 7 1 2 979 984
0 986 5 1 1 985
0 987 7 1 2 50863 986
0 988 5 1 1 987
0 989 7 1 2 41565 988
0 990 7 1 2 969 989
0 991 5 1 1 990
0 992 7 10 2 42230 49390
0 993 5 8 1 50915
0 994 7 4 2 43835 50139
0 995 7 2 2 48200 50859
0 996 7 1 2 50933 50937
0 997 5 1 1 996
0 998 7 7 2 41416 46018
0 999 7 4 2 43299 45376
0 1000 7 3 2 46702 50946
0 1001 7 1 2 49971 50950
0 1002 5 1 1 1001
0 1003 7 8 2 40545 42017
0 1004 5 4 1 50953
0 1005 7 1 2 50954 49993
0 1006 5 1 1 1005
0 1007 7 1 2 1002 1006
0 1008 5 1 1 1007
0 1009 7 1 2 50939 1008
0 1010 5 1 1 1009
0 1011 7 1 2 44856 1010
0 1012 7 1 2 997 1011
0 1013 5 1 1 1012
0 1014 7 1 2 50916 1013
0 1015 7 1 2 991 1014
0 1016 5 1 1 1015
0 1017 7 4 2 44996 50470
0 1018 7 7 2 41296 44720
0 1019 7 1 2 46190 50969
0 1020 7 1 2 50965 1019
0 1021 7 1 2 49139 1020
0 1022 5 1 1 1021
0 1023 7 1 2 1016 1022
0 1024 5 1 1 1023
0 1025 7 1 2 47610 1024
0 1026 5 1 1 1025
0 1027 7 5 2 47695 49391
0 1028 5 7 1 50976
0 1029 7 2 2 46019 50977
0 1030 7 2 2 42231 50988
0 1031 5 1 1 50990
0 1032 7 4 2 45377 49458
0 1033 5 6 1 50992
0 1034 7 2 2 50993 50052
0 1035 5 1 1 51002
0 1036 7 1 2 41064 50414
0 1037 5 1 1 1036
0 1038 7 1 2 1035 1037
0 1039 5 1 1 1038
0 1040 7 1 2 42748 1039
0 1041 5 1 1 1040
0 1042 7 1 2 1031 1041
0 1043 5 1 1 1042
0 1044 7 3 2 43836 41566
0 1045 7 2 2 44721 49994
0 1046 7 1 2 51004 51007
0 1047 7 1 2 1043 1046
0 1048 5 1 1 1047
0 1049 7 1 2 43990 1048
0 1050 7 1 2 1026 1049
0 1051 7 1 2 951 1050
0 1052 7 1 2 892 1051
0 1053 7 1 2 738 1052
0 1054 5 1 1 1053
0 1055 7 1 2 43837 41870
0 1056 5 6 1 1055
0 1057 7 2 2 49957 51009
0 1058 7 39 2 42018 42232
0 1059 5 10 1 51017
0 1060 7 4 2 47696 51018
0 1061 5 1 1 51066
0 1062 7 2 2 51015 51067
0 1063 5 1 1 51070
0 1064 7 1 2 47162 51010
0 1065 5 1 1 1064
0 1066 7 1 2 47611 50900
0 1067 5 1 1 1066
0 1068 7 1 2 1065 1067
0 1069 5 1 1 1068
0 1070 7 1 2 43300 1069
0 1071 5 1 1 1070
0 1072 7 6 2 42019 47612
0 1073 5 7 1 51072
0 1074 7 1 2 51078 531
0 1075 5 1 1 1074
0 1076 7 5 2 43838 42020
0 1077 5 5 1 51085
0 1078 7 4 2 40140 46995
0 1079 5 3 1 51095
0 1080 7 1 2 51090 51099
0 1081 7 1 2 1075 1080
0 1082 5 1 1 1081
0 1083 7 1 2 1071 1082
0 1084 5 3 1 1083
0 1085 7 1 2 42233 51102
0 1086 5 1 1 1085
0 1087 7 2 2 42021 48019
0 1088 5 1 1 51105
0 1089 7 2 2 44468 51106
0 1090 5 1 1 51107
0 1091 7 1 2 43488 51108
0 1092 5 2 1 1091
0 1093 7 1 2 1086 51109
0 1094 5 1 1 1093
0 1095 7 1 2 49392 1094
0 1096 5 1 1 1095
0 1097 7 1 2 1063 1096
0 1098 5 1 1 1097
0 1099 7 1 2 50092 1098
0 1100 5 1 1 1099
0 1101 7 2 2 43489 46917
0 1102 5 2 1 51111
0 1103 7 1 2 40546 51112
0 1104 5 1 1 1103
0 1105 7 4 2 47375 47613
0 1106 5 2 1 51115
0 1107 7 7 2 45222 47754
0 1108 5 2 1 51121
0 1109 7 1 2 51128 51011
0 1110 7 1 2 51116 1109
0 1111 5 1 1 1110
0 1112 7 1 2 1104 1111
0 1113 5 1 1 1112
0 1114 7 1 2 51019 1113
0 1115 5 1 1 1114
0 1116 7 3 2 42234 50707
0 1117 5 1 1 51130
0 1118 7 2 2 46729 46996
0 1119 5 2 1 51133
0 1120 7 1 2 47889 51134
0 1121 5 2 1 1120
0 1122 7 1 2 51131 51137
0 1123 5 1 1 1122
0 1124 7 1 2 1090 1123
0 1125 5 1 1 1124
0 1126 7 1 2 43490 1125
0 1127 5 1 1 1126
0 1128 7 2 2 47527 51012
0 1129 7 1 2 42022 51139
0 1130 5 1 1 1129
0 1131 7 1 2 44469 50708
0 1132 7 1 2 50860 1131
0 1133 5 1 1 1132
0 1134 7 1 2 1130 1133
0 1135 5 1 1 1134
0 1136 7 1 2 42235 1135
0 1137 5 1 1 1136
0 1138 7 1 2 1127 1137
0 1139 5 1 1 1138
0 1140 7 1 2 49393 1139
0 1141 5 1 1 1140
0 1142 7 1 2 1115 1141
0 1143 5 1 1 1142
0 1144 7 1 2 41417 49995
0 1145 7 1 2 1143 1144
0 1146 5 1 1 1145
0 1147 7 1 2 1100 1146
0 1148 5 1 1 1147
0 1149 7 1 2 48717 1148
0 1150 5 1 1 1149
0 1151 7 4 2 44390 48608
0 1152 5 5 1 51141
0 1153 7 4 2 40321 51145
0 1154 5 2 1 51150
0 1155 7 6 2 43839 45378
0 1156 5 5 1 51156
0 1157 7 10 2 42236 50687
0 1158 7 1 2 41170 51167
0 1159 5 1 1 1158
0 1160 7 1 2 51162 1159
0 1161 5 3 1 1160
0 1162 7 1 2 49680 51177
0 1163 5 1 1 1162
0 1164 7 1 2 50726 1163
0 1165 5 1 1 1164
0 1166 7 1 2 51151 1165
0 1167 5 1 1 1166
0 1168 7 2 2 43633 49689
0 1169 5 1 1 51180
0 1170 7 1 2 41297 1169
0 1171 7 1 2 51178 1170
0 1172 5 1 1 1171
0 1173 7 1 2 1167 1172
0 1174 5 1 1 1173
0 1175 7 1 2 51008 1174
0 1176 5 1 1 1175
0 1177 7 1 2 1150 1176
0 1178 5 1 1 1177
0 1179 7 1 2 44857 1178
0 1180 5 1 1 1179
0 1181 7 5 2 44470 42237
0 1182 5 2 1 51182
0 1183 7 2 2 43491 51183
0 1184 5 2 1 51189
0 1185 7 3 2 45564 47111
0 1186 5 8 1 51193
0 1187 7 1 2 43492 51196
0 1188 5 2 1 1187
0 1189 7 2 2 51187 51204
0 1190 5 2 1 51206
0 1191 7 1 2 47904 51208
0 1192 5 2 1 1191
0 1193 7 1 2 51191 51210
0 1194 5 1 1 1193
0 1195 7 1 2 49394 50646
0 1196 7 1 2 1194 1195
0 1197 5 1 1 1196
0 1198 7 1 2 1180 1197
0 1199 5 1 1 1198
0 1200 7 1 2 42749 1199
0 1201 5 1 1 1200
0 1202 7 16 2 41418 41567
0 1203 7 3 2 42909 51212
0 1204 7 1 2 51228 51103
0 1205 5 1 1 1204
0 1206 7 5 2 44722 44858
0 1207 7 4 2 43840 51231
0 1208 7 1 2 46703 49384
0 1209 5 4 1 1208
0 1210 7 1 2 43493 46868
0 1211 5 2 1 1210
0 1212 7 3 2 51240 51244
0 1213 5 7 1 51246
0 1214 7 2 2 46191 51249
0 1215 7 1 2 51236 51256
0 1216 5 1 1 1215
0 1217 7 1 2 1205 1216
0 1218 5 1 1 1217
0 1219 7 1 2 42238 1218
0 1220 5 1 1 1219
0 1221 7 4 2 42023 47309
0 1222 5 3 1 51258
0 1223 7 3 2 47697 51259
0 1224 5 1 1 51265
0 1225 7 14 2 44859 46192
0 1226 7 3 2 49558 50830
0 1227 7 1 2 51268 51282
0 1228 5 1 1 1227
0 1229 7 11 2 45565 42910
0 1230 7 1 2 51285 51213
0 1231 7 1 2 47528 1230
0 1232 5 1 1 1231
0 1233 7 1 2 1228 1232
0 1234 5 1 1 1233
0 1235 7 1 2 51266 1234
0 1236 5 1 1 1235
0 1237 7 1 2 1220 1236
0 1238 5 1 1 1237
0 1239 7 1 2 49395 1238
0 1240 5 1 1 1239
0 1241 7 1 2 51229 51071
0 1242 5 1 1 1241
0 1243 7 1 2 1240 1242
0 1244 5 1 1 1243
0 1245 7 8 2 44997 46020
0 1246 7 1 2 48718 51296
0 1247 7 1 2 1244 1246
0 1248 5 1 1 1247
0 1249 7 1 2 40716 1248
0 1250 7 1 2 1201 1249
0 1251 5 1 1 1250
0 1252 7 1 2 1054 1251
0 1253 5 1 1 1252
0 1254 7 1 2 44159 1253
0 1255 5 1 1 1254
0 1256 7 2 2 43991 44587
0 1257 7 1 2 46021 51304
0 1258 5 1 1 1257
0 1259 7 6 2 43301 40717
0 1260 7 2 2 44391 51306
0 1261 7 1 2 47845 51312
0 1262 5 1 1 1261
0 1263 7 1 2 1258 1262
0 1264 5 1 1 1263
0 1265 7 1 2 40547 1264
0 1266 5 1 1 1265
0 1267 7 6 2 44588 45223
0 1268 7 11 2 40718 42750
0 1269 5 1 1 51320
0 1270 7 1 2 51314 51321
0 1271 5 1 1 1270
0 1272 7 1 2 1266 1271
0 1273 5 1 1 1272
0 1274 7 1 2 42024 1273
0 1275 5 1 1 1274
0 1276 7 11 2 45379 42751
0 1277 7 5 2 40719 44589
0 1278 7 1 2 51331 51342
0 1279 7 1 2 47905 1278
0 1280 5 1 1 1279
0 1281 7 1 2 1275 1280
0 1282 5 1 1 1281
0 1283 7 1 2 50084 1282
0 1284 5 1 1 1283
0 1285 7 2 2 45380 46730
0 1286 5 3 1 51347
0 1287 7 3 2 47890 51348
0 1288 5 2 1 51352
0 1289 7 2 2 44590 51355
0 1290 5 2 1 51357
0 1291 7 12 2 43302 42025
0 1292 5 3 1 51361
0 1293 7 3 2 46704 51362
0 1294 5 9 1 51376
0 1295 7 1 2 51359 51379
0 1296 5 1 1 1295
0 1297 7 1 2 50064 49274
0 1298 7 1 2 1296 1297
0 1299 5 1 1 1298
0 1300 7 1 2 1284 1299
0 1301 5 1 1 1300
0 1302 7 1 2 44860 1301
0 1303 5 1 1 1302
0 1304 7 16 2 44723 46022
0 1305 5 1 1 51388
0 1306 7 6 2 43841 51389
0 1307 5 3 1 51404
0 1308 7 1 2 51405 50861
0 1309 5 1 1 1308
0 1310 7 7 2 41419 45224
0 1311 7 1 2 47953 51413
0 1312 5 1 1 1311
0 1313 7 1 2 1309 1312
0 1314 5 1 1 1313
0 1315 7 8 2 44591 44998
0 1316 7 1 2 51420 49159
0 1317 7 1 2 1314 1316
0 1318 5 1 1 1317
0 1319 7 1 2 1303 1318
0 1320 5 1 1 1319
0 1321 7 1 2 42911 1320
0 1322 5 1 1 1321
0 1323 7 6 2 44592 44861
0 1324 7 6 2 44724 44999
0 1325 7 3 2 51428 51434
0 1326 7 1 2 49263 51440
0 1327 7 1 2 50938 1326
0 1328 5 1 1 1327
0 1329 7 1 2 1322 1328
0 1330 5 1 1 1329
0 1331 7 1 2 43634 1330
0 1332 5 1 1 1331
0 1333 7 4 2 43992 41698
0 1334 7 2 2 49559 51443
0 1335 5 1 1 51447
0 1336 7 15 2 40548 40720
0 1337 5 1 1 51449
0 1338 7 12 2 41420 51450
0 1339 7 2 2 45000 51464
0 1340 5 1 1 51476
0 1341 7 1 2 1335 1340
0 1342 5 3 1 1341
0 1343 7 1 2 48567 51429
0 1344 7 1 2 51377 1343
0 1345 7 1 2 51478 1344
0 1346 5 1 1 1345
0 1347 7 1 2 1332 1346
0 1348 5 1 1 1347
0 1349 7 1 2 47614 1348
0 1350 5 1 1 1349
0 1351 7 12 2 40721 41421
0 1352 7 3 2 42912 51481
0 1353 7 1 2 51493 51140
0 1354 5 1 1 1353
0 1355 7 3 2 46193 47906
0 1356 5 1 1 51496
0 1357 7 1 2 49275 51497
0 1358 5 1 1 1357
0 1359 7 1 2 1354 1358
0 1360 5 1 1 1359
0 1361 7 1 2 48954 1360
0 1362 5 1 1 1361
0 1363 7 4 2 49264 50729
0 1364 7 2 2 51499 50115
0 1365 5 1 1 51503
0 1366 7 1 2 1362 1365
0 1367 5 1 1 1366
0 1368 7 1 2 45001 1367
0 1369 5 1 1 1368
0 1370 7 5 2 41699 48568
0 1371 7 2 2 49560 51505
0 1372 5 1 1 51510
0 1373 7 60 2 43993 44862
0 1374 5 3 1 51512
0 1375 7 1 2 47529 51513
0 1376 7 1 2 51511 1375
0 1377 5 1 1 1376
0 1378 7 1 2 1369 1377
0 1379 5 1 1 1378
0 1380 7 1 2 49930 1379
0 1381 5 1 1 1380
0 1382 7 4 2 44593 47615
0 1383 5 4 1 51575
0 1384 7 3 2 50198 51579
0 1385 5 2 1 51583
0 1386 7 8 2 49459 51584
0 1387 5 2 1 51588
0 1388 7 2 2 47444 51589
0 1389 5 1 1 51598
0 1390 7 1 2 47755 48644
0 1391 5 17 1 1390
0 1392 7 1 2 1389 51600
0 1393 5 3 1 1392
0 1394 7 12 2 45002 41871
0 1395 5 3 1 51620
0 1396 7 2 2 44725 51621
0 1397 7 2 2 48569 49175
0 1398 7 1 2 51635 51637
0 1399 7 1 2 51617 1398
0 1400 5 1 1 1399
0 1401 7 1 2 1381 1400
0 1402 5 1 1 1401
0 1403 7 1 2 42026 1402
0 1404 5 1 1 1403
0 1405 7 1 2 50019 48955
0 1406 5 1 1 1405
0 1407 7 8 2 42913 49070
0 1408 5 2 1 51639
0 1409 7 1 2 45003 51640
0 1410 5 1 1 1409
0 1411 7 1 2 1406 1410
0 1412 5 1 1 1411
0 1413 7 1 2 49276 1412
0 1414 5 1 1 1413
0 1415 7 2 2 40722 48570
0 1416 7 7 2 44863 45381
0 1417 5 1 1 51651
0 1418 7 1 2 50085 51652
0 1419 7 1 2 51649 1418
0 1420 5 1 1 1419
0 1421 7 1 2 1414 1420
0 1422 5 1 1 1421
0 1423 7 1 2 50978 1422
0 1424 5 1 1 1423
0 1425 7 1 2 1404 1424
0 1426 7 1 2 1350 1425
0 1427 5 1 1 1426
0 1428 7 1 2 42239 1427
0 1429 5 1 1 1428
0 1430 7 1 2 49561 51003
0 1431 5 1 1 1430
0 1432 7 3 2 42027 49958
0 1433 5 2 1 51658
0 1434 7 1 2 49738 51659
0 1435 5 1 1 1434
0 1436 7 1 2 49562 51152
0 1437 5 1 1 1436
0 1438 7 1 2 1435 1437
0 1439 5 1 1 1438
0 1440 7 1 2 45566 1439
0 1441 5 1 1 1440
0 1442 7 1 2 1431 1441
0 1443 5 1 1 1442
0 1444 7 1 2 40723 1443
0 1445 5 1 1 1444
0 1446 7 4 2 43994 41298
0 1447 7 8 2 40322 46997
0 1448 5 2 1 51667
0 1449 7 2 2 51663 51668
0 1450 7 2 2 48622 50648
0 1451 5 1 1 51679
0 1452 7 1 2 51677 51680
0 1453 5 1 1 1452
0 1454 7 1 2 1445 1453
0 1455 5 1 1 1454
0 1456 7 1 2 44864 1455
0 1457 5 1 1 1456
0 1458 7 1 2 40141 50994
0 1459 5 1 1 1458
0 1460 7 1 2 50424 1459
0 1461 5 1 1 1460
0 1462 7 1 2 47445 1461
0 1463 5 1 1 1462
0 1464 7 9 2 40142 45567
0 1465 5 1 1 51681
0 1466 7 1 2 50294 1465
0 1467 5 2 1 1466
0 1468 7 1 2 40323 51690
0 1469 5 1 1 1468
0 1470 7 1 2 1463 1469
0 1471 5 1 1 1470
0 1472 7 1 2 51500 1471
0 1473 5 1 1 1472
0 1474 7 1 2 1457 1473
0 1475 5 1 1 1474
0 1476 7 1 2 42914 1475
0 1477 5 1 1 1476
0 1478 7 3 2 44865 49265
0 1479 7 7 2 44726 51692
0 1480 7 7 2 43494 47076
0 1481 5 4 1 51702
0 1482 7 3 2 49396 51703
0 1483 5 1 1 51713
0 1484 7 2 2 51695 51714
0 1485 7 1 2 51498 51716
0 1486 5 1 1 1485
0 1487 7 1 2 1477 1486
0 1488 5 1 1 1487
0 1489 7 1 2 42752 1488
0 1490 5 1 1 1489
0 1491 7 1 2 51504 51715
0 1492 5 1 1 1491
0 1493 7 1 2 1490 1492
0 1494 5 1 1 1493
0 1495 7 1 2 45004 1494
0 1496 5 1 1 1495
0 1497 7 1 2 47907 51506
0 1498 7 1 2 51717 1497
0 1499 5 1 1 1498
0 1500 7 1 2 40903 1499
0 1501 7 1 2 1496 1500
0 1502 7 1 2 1429 1501
0 1503 5 1 1 1502
0 1504 7 1 2 1255 1503
0 1505 5 1 1 1504
0 1506 7 1 2 42451 1505
0 1507 5 1 1 1506
0 1508 7 1 2 46322 1507
0 1509 7 1 2 574 1508
0 1510 5 1 1 1509
0 1511 7 2 2 41700 48532
0 1512 7 12 2 44866 45792
0 1513 7 1 2 39936 50896
0 1514 5 1 1 1513
0 1515 7 1 2 50709 51349
0 1516 7 2 2 1514 1515
0 1517 7 1 2 49931 51732
0 1518 5 2 1 1517
0 1519 7 11 2 41065 45382
0 1520 5 2 1 51736
0 1521 7 2 2 47756 49710
0 1522 5 1 1 51749
0 1523 7 1 2 51737 51750
0 1524 5 1 1 1523
0 1525 7 6 2 47616 49397
0 1526 5 9 1 51751
0 1527 7 1 2 50710 51752
0 1528 7 1 2 1524 1527
0 1529 5 1 1 1528
0 1530 7 1 2 51734 1529
0 1531 5 1 1 1530
0 1532 7 1 2 42240 1531
0 1533 5 1 1 1532
0 1534 7 3 2 47077 46705
0 1535 5 1 1 51766
0 1536 7 2 2 43303 51767
0 1537 5 2 1 51769
0 1538 7 1 2 43495 47203
0 1539 5 1 1 1538
0 1540 7 4 2 51771 1539
0 1541 5 6 1 51773
0 1542 7 3 2 45568 49398
0 1543 5 1 1 51783
0 1544 7 1 2 51777 51784
0 1545 5 1 1 1544
0 1546 7 1 2 1533 1545
0 1547 5 2 1 1546
0 1548 7 1 2 51720 51786
0 1549 5 1 1 1548
0 1550 7 7 2 42028 49870
0 1551 5 3 1 51788
0 1552 7 3 2 45383 47757
0 1553 5 4 1 51798
0 1554 7 1 2 51801 51117
0 1555 5 2 1 1554
0 1556 7 1 2 51795 51805
0 1557 5 1 1 1556
0 1558 7 1 2 45569 1557
0 1559 5 2 1 1558
0 1560 7 3 2 47446 47576
0 1561 5 14 1 51809
0 1562 7 4 2 45570 48719
0 1563 5 1 1 51826
0 1564 7 1 2 50600 1563
0 1565 5 5 1 1564
0 1566 7 1 2 51812 51830
0 1567 5 2 1 1566
0 1568 7 1 2 44392 46973
0 1569 5 1 1 1568
0 1570 7 1 2 51020 1569
0 1571 5 1 1 1570
0 1572 7 1 2 51835 1571
0 1573 7 1 2 51807 1572
0 1574 5 1 1 1573
0 1575 7 1 2 41872 1574
0 1576 5 1 1 1575
0 1577 7 2 2 43496 47031
0 1578 5 3 1 51837
0 1579 7 7 2 47112 51839
0 1580 7 14 2 40143 45384
0 1581 5 6 1 51849
0 1582 7 8 2 41171 51850
0 1583 5 17 1 51869
0 1584 7 1 2 47310 51877
0 1585 5 1 1 1584
0 1586 7 4 2 51842 1585
0 1587 5 4 1 51894
0 1588 7 1 2 45571 51898
0 1589 5 2 1 1588
0 1590 7 1 2 50601 51902
0 1591 5 1 1 1590
0 1592 7 1 2 48720 1591
0 1593 5 1 1 1592
0 1594 7 1 2 49460 1224
0 1595 5 1 1 1594
0 1596 7 1 2 45572 1595
0 1597 5 1 1 1596
0 1598 7 1 2 1593 1597
0 1599 7 1 2 1576 1598
0 1600 5 1 1 1599
0 1601 7 1 2 45793 1600
0 1602 5 2 1 1601
0 1603 7 33 2 42241 45794
0 1604 5 3 1 51906
0 1605 7 1 2 48645 51895
0 1606 5 1 1 1605
0 1607 7 1 2 51907 1606
0 1608 5 2 1 1607
0 1609 7 4 2 40144 42452
0 1610 7 4 2 41299 47447
0 1611 5 4 1 51948
0 1612 7 6 2 41066 45573
0 1613 7 3 2 39937 51956
0 1614 5 4 1 51962
0 1615 7 1 2 51952 51965
0 1616 5 1 1 1615
0 1617 7 1 2 51944 1616
0 1618 5 1 1 1617
0 1619 7 1 2 51942 1618
0 1620 5 1 1 1619
0 1621 7 1 2 45225 1620
0 1622 5 1 1 1621
0 1623 7 1 2 51904 1622
0 1624 5 1 1 1623
0 1625 7 1 2 44867 1624
0 1626 5 1 1 1625
0 1627 7 11 2 41568 42453
0 1628 5 1 1 51969
0 1629 7 36 2 41300 45574
0 1630 5 20 1 51980
0 1631 7 4 2 43635 52016
0 1632 5 5 1 52036
0 1633 7 2 2 52040 48843
0 1634 5 13 1 52045
0 1635 7 1 2 52047 51778
0 1636 5 2 1 1635
0 1637 7 9 2 40145 46783
0 1638 5 5 1 52062
0 1639 7 2 2 52071 47032
0 1640 5 4 1 52076
0 1641 7 1 2 39938 52078
0 1642 5 3 1 1641
0 1643 7 1 2 46731 51096
0 1644 5 2 1 1643
0 1645 7 1 2 52082 52085
0 1646 5 1 1 1645
0 1647 7 3 2 43497 46826
0 1648 5 24 1 52087
0 1649 7 1 2 47113 52090
0 1650 7 2 2 1646 1649
0 1651 5 3 1 52114
0 1652 7 2 2 49399 52116
0 1653 5 1 1 52119
0 1654 7 1 2 42242 52120
0 1655 5 1 1 1654
0 1656 7 1 2 52060 1655
0 1657 5 8 1 1656
0 1658 7 1 2 51970 52121
0 1659 5 1 1 1658
0 1660 7 1 2 1626 1659
0 1661 5 1 1 1660
0 1662 7 1 2 49563 1661
0 1663 5 1 1 1662
0 1664 7 1 2 1549 1663
0 1665 5 1 1 1664
0 1666 7 1 2 51718 1665
0 1667 5 1 1 1666
0 1668 7 9 2 44868 42454
0 1669 7 1 2 52129 50934
0 1670 5 1 1 1669
0 1671 7 10 2 40549 50392
0 1672 5 3 1 52138
0 1673 7 1 2 52148 917
0 1674 5 10 1 1673
0 1675 7 8 2 45005 45795
0 1676 7 1 2 52161 51669
0 1677 7 1 2 52151 1676
0 1678 5 1 1 1677
0 1679 7 1 2 1670 1678
0 1680 5 1 1 1679
0 1681 7 1 2 51981 1680
0 1682 5 1 1 1681
0 1683 7 23 2 42029 45796
0 1684 5 1 1 52169
0 1685 7 5 2 41873 52170
0 1686 7 5 2 44869 42243
0 1687 7 1 2 52192 52197
0 1688 7 1 2 50935 1687
0 1689 5 1 1 1688
0 1690 7 1 2 1682 1689
0 1691 5 1 1 1690
0 1692 7 1 2 48623 1691
0 1693 5 1 1 1692
0 1694 7 1 2 46023 1693
0 1695 7 1 2 1667 1694
0 1696 5 1 1 1695
0 1697 7 8 2 40550 50086
0 1698 7 1 2 41569 52202
0 1699 5 1 1 1698
0 1700 7 1 2 643 1699
0 1701 5 1 1 1700
0 1702 7 6 2 40324 51982
0 1703 5 6 1 52210
0 1704 7 2 2 46998 52211
0 1705 5 1 1 52222
0 1706 7 1 2 1701 52223
0 1707 5 1 1 1706
0 1708 7 12 2 41570 41701
0 1709 7 10 2 43636 47078
0 1710 5 3 1 52236
0 1711 7 3 2 43637 52072
0 1712 5 5 1 52249
0 1713 7 7 2 43498 46706
0 1714 5 7 1 52257
0 1715 7 1 2 40325 52264
0 1716 5 5 1 1715
0 1717 7 1 2 43304 52271
0 1718 5 2 1 1717
0 1719 7 1 2 52252 52276
0 1720 5 2 1 1719
0 1721 7 1 2 47033 52278
0 1722 5 1 1 1721
0 1723 7 1 2 40146 50841
0 1724 5 1 1 1723
0 1725 7 10 2 50378 1724
0 1726 5 5 1 52280
0 1727 7 1 2 47143 52281
0 1728 5 1 1 1727
0 1729 7 2 2 1722 1728
0 1730 5 1 1 52295
0 1731 7 1 2 52246 52296
0 1732 5 6 1 1731
0 1733 7 1 2 41422 48844
0 1734 5 4 1 1733
0 1735 7 2 2 40551 48845
0 1736 5 3 1 52307
0 1737 7 3 2 52303 52309
0 1738 5 1 1 52312
0 1739 7 1 2 48533 52313
0 1740 7 1 2 52297 1739
0 1741 5 1 1 1740
0 1742 7 20 2 40147 45226
0 1743 5 6 1 52315
0 1744 7 5 2 47259 52316
0 1745 5 8 1 52341
0 1746 7 1 2 47034 52346
0 1747 5 1 1 1746
0 1748 7 1 2 47139 1747
0 1749 5 1 1 1748
0 1750 7 1 2 49564 1749
0 1751 5 1 1 1750
0 1752 7 10 2 42030 46974
0 1753 7 2 2 48534 52354
0 1754 5 2 1 52364
0 1755 7 1 2 49626 52366
0 1756 5 1 1 1755
0 1757 7 1 2 52282 1756
0 1758 5 1 1 1757
0 1759 7 2 2 48535 49798
0 1760 7 6 2 41874 47035
0 1761 5 2 1 52370
0 1762 7 1 2 47376 52371
0 1763 7 1 2 52368 1762
0 1764 5 1 1 1763
0 1765 7 1 2 1758 1764
0 1766 7 1 2 1751 1765
0 1767 5 1 1 1766
0 1768 7 1 2 52017 1767
0 1769 5 1 1 1768
0 1770 7 9 2 44727 42244
0 1771 5 1 1 52378
0 1772 7 1 2 52379 49833
0 1773 5 1 1 1772
0 1774 7 1 2 1769 1773
0 1775 7 1 2 1741 1774
0 1776 5 1 1 1775
0 1777 7 1 2 52224 1776
0 1778 5 1 1 1777
0 1779 7 1 2 1707 1778
0 1780 5 1 1 1779
0 1781 7 1 2 45797 1780
0 1782 5 1 1 1781
0 1783 7 15 2 40148 41067
0 1784 5 9 1 52387
0 1785 7 6 2 39939 52388
0 1786 5 12 1 52411
0 1787 7 1 2 44594 52417
0 1788 5 1 1 1787
0 1789 7 1 2 42455 50791
0 1790 7 1 2 50936 1789
0 1791 7 1 2 1788 1790
0 1792 5 1 1 1791
0 1793 7 1 2 42753 1792
0 1794 7 1 2 1782 1793
0 1795 5 1 1 1794
0 1796 7 1 2 46194 1795
0 1797 7 1 2 1696 1796
0 1798 5 1 1 1797
0 1799 7 36 2 45575 42456
0 1800 5 3 1 52429
0 1801 7 5 2 52430 50272
0 1802 5 4 1 52468
0 1803 7 5 2 50317 52171
0 1804 5 8 1 52477
0 1805 7 14 2 45385 42457
0 1806 5 1 1 52490
0 1807 7 2 2 45227 52491
0 1808 7 1 2 51957 52504
0 1809 5 1 1 1808
0 1810 7 1 2 52482 1809
0 1811 5 1 1 1810
0 1812 7 1 2 39940 1811
0 1813 5 1 1 1812
0 1814 7 12 2 41301 45228
0 1815 5 1 1 52506
0 1816 7 1 2 52507 52492
0 1817 5 3 1 1816
0 1818 7 1 2 52518 52483
0 1819 5 1 1 1818
0 1820 7 1 2 41068 1819
0 1821 5 1 1 1820
0 1822 7 2 2 1813 1821
0 1823 5 1 1 52521
0 1824 7 1 2 52473 52522
0 1825 5 1 1 1824
0 1826 7 1 2 40149 1825
0 1827 5 1 1 1826
0 1828 7 8 2 45386 52431
0 1829 5 1 1 52523
0 1830 7 1 2 39941 52524
0 1831 5 1 1 1830
0 1832 7 1 2 52484 1831
0 1833 5 1 1 1832
0 1834 7 1 2 41302 1833
0 1835 5 1 1 1834
0 1836 7 1 2 1827 1835
0 1837 5 1 1 1836
0 1838 7 1 2 41172 1837
0 1839 5 1 1 1838
0 1840 7 8 2 41303 45798
0 1841 7 3 2 41875 51021
0 1842 5 2 1 52539
0 1843 7 2 2 52531 52540
0 1844 7 1 2 49767 52544
0 1845 5 1 1 1844
0 1846 7 1 2 1839 1845
0 1847 5 1 1 1846
0 1848 7 1 2 49972 1847
0 1849 5 1 1 1848
0 1850 7 8 2 39942 47758
0 1851 5 4 1 52546
0 1852 7 2 2 52547 52478
0 1853 5 1 1 52558
0 1854 7 1 2 41069 52559
0 1855 5 1 1 1854
0 1856 7 4 2 42458 46999
0 1857 5 1 1 52560
0 1858 7 1 2 51983 52561
0 1859 5 1 1 1858
0 1860 7 1 2 1855 1859
0 1861 5 1 1 1860
0 1862 7 1 2 49996 1861
0 1863 5 1 1 1862
0 1864 7 1 2 1849 1863
0 1865 5 1 1 1864
0 1866 7 1 2 40326 1865
0 1867 5 1 1 1866
0 1868 7 1 2 51810 49973
0 1869 5 1 1 1868
0 1870 7 5 2 47759 47260
0 1871 7 1 2 52564 49997
0 1872 5 1 1 1871
0 1873 7 1 2 1869 1872
0 1874 5 1 1 1873
0 1875 7 1 2 52545 1874
0 1876 5 1 1 1875
0 1877 7 1 2 1867 1876
0 1878 5 1 1 1877
0 1879 7 1 2 49071 1878
0 1880 5 1 1 1879
0 1881 7 6 2 42031 51908
0 1882 5 3 1 52569
0 1883 7 2 2 49923 52570
0 1884 7 1 2 50151 52578
0 1885 5 1 1 1884
0 1886 7 10 2 41304 50174
0 1887 7 3 2 42459 52580
0 1888 7 1 2 50471 52590
0 1889 5 2 1 1888
0 1890 7 1 2 1885 52593
0 1891 5 2 1 1890
0 1892 7 1 2 50080 52595
0 1893 5 1 1 1892
0 1894 7 1 2 1880 1893
0 1895 5 1 1 1894
0 1896 7 1 2 49627 1895
0 1897 5 1 1 1896
0 1898 7 4 2 46024 52225
0 1899 5 1 1 52597
0 1900 7 17 2 45799 42915
0 1901 7 4 2 52601 51984
0 1902 7 7 2 40327 44728
0 1903 7 1 2 47000 52622
0 1904 7 1 2 52618 1903
0 1905 7 1 2 52598 1904
0 1906 5 1 1 1905
0 1907 7 1 2 43995 1906
0 1908 7 1 2 1897 1907
0 1909 7 1 2 1798 1908
0 1910 5 1 1 1909
0 1911 7 18 2 46025 46195
0 1912 7 4 2 44870 52629
0 1913 7 2 2 41305 50711
0 1914 5 4 1 52651
0 1915 7 1 2 43638 52653
0 1916 5 1 1 1915
0 1917 7 2 2 51774 1916
0 1918 5 1 1 52657
0 1919 7 1 2 52647 1918
0 1920 5 1 1 1919
0 1921 7 1 2 41306 51670
0 1922 7 1 2 48258 1921
0 1923 5 1 1 1922
0 1924 7 1 2 1920 1923
0 1925 5 1 1 1924
0 1926 7 1 2 45576 1925
0 1927 5 1 1 1926
0 1928 7 5 2 45387 46026
0 1929 7 1 2 44871 52659
0 1930 5 1 1 1929
0 1931 7 1 2 47241 1930
0 1932 5 2 1 1931
0 1933 7 1 2 51813 52664
0 1934 5 1 1 1933
0 1935 7 5 2 43639 44393
0 1936 7 2 2 44471 48609
0 1937 7 6 2 52666 52671
0 1938 5 5 1 52673
0 1939 7 15 2 42032 46027
0 1940 7 6 2 44872 52684
0 1941 5 1 1 52699
0 1942 7 1 2 52679 52700
0 1943 5 1 1 1942
0 1944 7 1 2 1934 1943
0 1945 5 1 1 1944
0 1946 7 1 2 41876 1945
0 1947 5 1 1 1946
0 1948 7 7 2 45229 46028
0 1949 5 1 1 52705
0 1950 7 2 2 44873 52706
0 1951 5 1 1 52712
0 1952 7 1 2 47242 1951
0 1953 5 4 1 1952
0 1954 7 1 2 52714 51899
0 1955 5 1 1 1954
0 1956 7 1 2 1947 1955
0 1957 5 1 1 1956
0 1958 7 1 2 42245 1957
0 1959 5 1 1 1958
0 1960 7 3 2 49461 51775
0 1961 5 1 1 52718
0 1962 7 1 2 47212 1961
0 1963 5 1 1 1962
0 1964 7 1 2 1959 1963
0 1965 5 1 1 1964
0 1966 7 1 2 46196 1965
0 1967 5 1 1 1966
0 1968 7 1 2 1927 1967
0 1969 5 1 1 1968
0 1970 7 1 2 45006 1969
0 1971 5 1 1 1970
0 1972 7 3 2 43499 42033
0 1973 5 4 1 52721
0 1974 7 1 2 45577 52724
0 1975 5 5 1 1974
0 1976 7 1 2 46778 52728
0 1977 5 1 1 1976
0 1978 7 2 2 45578 46927
0 1979 5 1 1 52733
0 1980 7 1 2 43305 52701
0 1981 5 1 1 1980
0 1982 7 1 2 40150 1981
0 1983 5 1 1 1982
0 1984 7 1 2 1979 1983
0 1985 5 1 1 1984
0 1986 7 1 2 1977 1985
0 1987 5 1 1 1986
0 1988 7 1 2 49340 1987
0 1989 5 1 1 1988
0 1990 7 1 2 43500 46657
0 1991 5 1 1 1990
0 1992 7 1 2 505 1991
0 1993 5 2 1 1992
0 1994 7 1 2 51197 52735
0 1995 5 1 1 1994
0 1996 7 7 2 44874 48332
0 1997 7 1 2 44472 52737
0 1998 5 1 1 1997
0 1999 7 1 2 51838 49290
0 2000 5 1 1 1999
0 2001 7 1 2 1998 2000
0 2002 7 1 2 1995 2001
0 2003 5 1 1 2002
0 2004 7 1 2 46827 2003
0 2005 5 1 1 2004
0 2006 7 3 2 41571 47954
0 2007 5 3 1 52744
0 2008 7 1 2 46925 52745
0 2009 5 1 1 2008
0 2010 7 2 2 42754 50472
0 2011 5 2 1 52750
0 2012 7 1 2 52581 52751
0 2013 5 1 1 2012
0 2014 7 1 2 50248 48333
0 2015 7 1 2 51802 2014
0 2016 5 1 1 2015
0 2017 7 1 2 2013 2016
0 2018 5 1 1 2017
0 2019 7 1 2 44875 2018
0 2020 5 1 1 2019
0 2021 7 1 2 2009 2020
0 2022 7 1 2 2005 2021
0 2023 7 1 2 1989 2022
0 2024 5 1 1 2023
0 2025 7 1 2 49998 2024
0 2026 5 1 1 2025
0 2027 7 1 2 1971 2026
0 2028 5 1 1 2027
0 2029 7 1 2 41423 2028
0 2030 5 1 1 2029
0 2031 7 3 2 48093 49848
0 2032 5 1 1 52754
0 2033 7 5 2 45007 42755
0 2034 7 3 2 46197 52757
0 2035 7 1 2 41572 52762
0 2036 5 1 1 2035
0 2037 7 2 2 2032 2036
0 2038 5 6 1 52765
0 2039 7 1 2 52548 52767
0 2040 5 1 1 2039
0 2041 7 5 2 41173 45008
0 2042 7 3 2 40151 52773
0 2043 7 2 2 52648 52778
0 2044 5 1 1 52781
0 2045 7 1 2 2040 2044
0 2046 5 1 1 2045
0 2047 7 1 2 41877 2046
0 2048 5 1 1 2047
0 2049 7 5 2 45230 42916
0 2050 7 5 2 40152 41573
0 2051 7 1 2 50065 52788
0 2052 7 1 2 52783 2051
0 2053 5 1 1 2052
0 2054 7 1 2 2048 2053
0 2055 5 1 1 2054
0 2056 7 1 2 41070 2055
0 2057 5 1 1 2056
0 2058 7 5 2 39943 41878
0 2059 5 1 1 52793
0 2060 7 1 2 52794 52782
0 2061 5 1 1 2060
0 2062 7 1 2 2057 2061
0 2063 5 1 1 2062
0 2064 7 1 2 49462 2063
0 2065 5 1 1 2064
0 2066 7 8 2 47377 47698
0 2067 5 11 1 52798
0 2068 7 2 2 52630 52806
0 2069 7 2 2 44876 48646
0 2070 7 1 2 51622 52819
0 2071 7 1 2 52817 2070
0 2072 5 1 1 2071
0 2073 7 1 2 2065 2072
0 2074 5 1 1 2073
0 2075 7 1 2 51022 2074
0 2076 5 1 1 2075
0 2077 7 1 2 2030 2076
0 2078 5 1 1 2077
0 2079 7 1 2 40552 2078
0 2080 5 1 1 2079
0 2081 7 1 2 49565 48201
0 2082 5 3 1 2081
0 2083 7 2 2 42917 49463
0 2084 7 1 2 52565 50940
0 2085 7 1 2 52824 2084
0 2086 5 1 1 2085
0 2087 7 1 2 52821 2086
0 2088 5 1 1 2087
0 2089 7 1 2 44877 2088
0 2090 5 1 1 2089
0 2091 7 1 2 50804 48397
0 2092 5 1 1 2091
0 2093 7 1 2 2090 2092
0 2094 5 1 1 2093
0 2095 7 1 2 41702 2094
0 2096 5 1 1 2095
0 2097 7 2 2 47261 49464
0 2098 7 1 2 47213 52826
0 2099 5 1 1 2098
0 2100 7 1 2 48647 46658
0 2101 5 1 1 2100
0 2102 7 1 2 2099 2101
0 2103 5 1 1 2102
0 2104 7 1 2 47760 2103
0 2105 5 1 1 2104
0 2106 7 2 2 47448 46659
0 2107 5 2 1 52828
0 2108 7 1 2 51590 52829
0 2109 5 1 1 2108
0 2110 7 1 2 2105 2109
0 2111 5 1 1 2110
0 2112 7 1 2 50093 2111
0 2113 5 1 1 2112
0 2114 7 1 2 2096 2113
0 2115 5 1 1 2114
0 2116 7 1 2 41879 2115
0 2117 5 1 1 2116
0 2118 7 4 2 41703 45231
0 2119 7 2 2 42756 51214
0 2120 7 2 2 52832 52836
0 2121 7 1 2 52389 52825
0 2122 7 1 2 52838 2121
0 2123 5 1 1 2122
0 2124 7 1 2 2117 2123
0 2125 5 1 1 2124
0 2126 7 1 2 51023 2125
0 2127 5 1 1 2126
0 2128 7 2 2 41574 49974
0 2129 7 1 2 51814 52660
0 2130 7 1 2 52840 2129
0 2131 5 1 1 2130
0 2132 7 3 2 41174 47449
0 2133 5 6 1 52842
0 2134 7 1 2 51851 52843
0 2135 5 2 1 2134
0 2136 7 1 2 41704 48259
0 2137 7 1 2 52851 2136
0 2138 5 1 1 2137
0 2139 7 1 2 2131 2138
0 2140 5 1 1 2139
0 2141 7 1 2 41880 2140
0 2142 5 1 1 2141
0 2143 7 8 2 41705 46198
0 2144 5 1 1 52853
0 2145 7 12 2 45009 42918
0 2146 5 1 1 52861
0 2147 7 7 2 2144 2146
0 2148 7 1 2 49072 52873
0 2149 5 1 1 2148
0 2150 7 1 2 698 2149
0 2151 5 2 1 2150
0 2152 7 1 2 51632 51900
0 2153 7 1 2 52880 2152
0 2154 5 1 1 2153
0 2155 7 1 2 2142 2154
0 2156 5 1 1 2155
0 2157 7 1 2 42246 2156
0 2158 5 1 1 2157
0 2159 7 6 2 45010 42247
0 2160 5 2 1 52882
0 2161 7 2 2 51779 52881
0 2162 7 1 2 52888 52890
0 2163 5 1 1 2162
0 2164 7 1 2 2158 2163
0 2165 5 1 1 2164
0 2166 7 6 2 48536 49400
0 2167 7 1 2 2165 52892
0 2168 5 1 1 2167
0 2169 7 1 2 47243 61
0 2170 5 53 1 2169
0 2171 7 4 2 46199 52898
0 2172 7 11 2 41175 44729
0 2173 7 3 2 48648 52955
0 2174 5 1 1 52966
0 2175 7 3 2 46029 48610
0 2176 5 2 1 52969
0 2177 7 1 2 52972 50966
0 2178 7 1 2 52967 2177
0 2179 7 1 2 52951 2178
0 2180 5 1 1 2179
0 2181 7 1 2 45800 2180
0 2182 7 1 2 2168 2181
0 2183 7 1 2 2127 2182
0 2184 7 1 2 2080 2183
0 2185 5 1 1 2184
0 2186 7 6 2 45388 50175
0 2187 5 1 1 52974
0 2188 7 2 2 49628 52975
0 2189 5 1 1 52980
0 2190 7 1 2 48537 2189
0 2191 5 3 1 2190
0 2192 7 4 2 40153 41307
0 2193 7 3 2 46784 52985
0 2194 5 2 1 52989
0 2195 7 2 2 41308 48624
0 2196 5 1 1 52994
0 2197 7 1 2 52347 2196
0 2198 5 3 1 2197
0 2199 7 1 2 45579 52996
0 2200 5 2 1 2199
0 2201 7 1 2 52992 52999
0 2202 5 1 1 2201
0 2203 7 1 2 46660 2202
0 2204 5 1 1 2203
0 2205 7 6 2 41309 42757
0 2206 7 1 2 53001 50792
0 2207 5 1 1 2206
0 2208 7 1 2 2204 2207
0 2209 5 1 1 2208
0 2210 7 1 2 52982 2209
0 2211 5 1 1 2210
0 2212 7 7 2 39944 44730
0 2213 7 2 2 47761 51168
0 2214 5 1 1 53014
0 2215 7 1 2 51163 2214
0 2216 5 1 1 2215
0 2217 7 1 2 49465 2216
0 2218 5 2 1 2217
0 2219 7 1 2 43842 51870
0 2220 5 1 1 2219
0 2221 7 1 2 53016 2220
0 2222 5 1 1 2221
0 2223 7 1 2 41071 2222
0 2224 5 1 1 2223
0 2225 7 2 2 40154 50774
0 2226 7 1 2 45232 53018
0 2227 5 1 1 2226
0 2228 7 1 2 2224 2227
0 2229 5 1 1 2228
0 2230 7 1 2 53007 2229
0 2231 5 2 1 2230
0 2232 7 1 2 47114 52290
0 2233 5 3 1 2232
0 2234 7 1 2 42248 53022
0 2235 5 1 1 2234
0 2236 7 1 2 47079 52283
0 2237 5 2 1 2236
0 2238 7 1 2 42249 52073
0 2239 5 1 1 2238
0 2240 7 1 2 39945 2239
0 2241 5 2 1 2240
0 2242 7 1 2 45580 52265
0 2243 5 1 1 2242
0 2244 7 1 2 47036 2243
0 2245 7 1 2 53027 2244
0 2246 5 1 1 2245
0 2247 7 1 2 53025 2246
0 2248 7 1 2 2235 2247
0 2249 5 1 1 2248
0 2250 7 1 2 49401 2249
0 2251 5 1 1 2250
0 2252 7 9 2 43843 42250
0 2253 5 1 1 53029
0 2254 7 2 2 53030 50688
0 2255 5 2 1 53038
0 2256 7 1 2 2251 53040
0 2257 5 2 1 2256
0 2258 7 1 2 41424 53042
0 2259 5 2 1 2258
0 2260 7 1 2 53020 53044
0 2261 5 1 1 2260
0 2262 7 1 2 49073 2261
0 2263 5 1 1 2262
0 2264 7 1 2 2211 2263
0 2265 5 1 1 2264
0 2266 7 1 2 45011 2265
0 2267 5 1 1 2266
0 2268 7 4 2 44878 50066
0 2269 5 2 1 53046
0 2270 7 2 2 43844 50504
0 2271 5 1 1 53052
0 2272 7 1 2 40155 53053
0 2273 5 1 1 2272
0 2274 7 1 2 53017 2273
0 2275 5 1 1 2274
0 2276 7 1 2 44731 47262
0 2277 7 1 2 2275 2276
0 2278 5 1 1 2277
0 2279 7 1 2 53045 2278
0 2280 5 1 1 2279
0 2281 7 1 2 53047 2280
0 2282 5 1 1 2281
0 2283 7 1 2 2267 2282
0 2284 5 1 1 2283
0 2285 7 1 2 46200 2284
0 2286 5 1 1 2285
0 2287 7 1 2 46030 53043
0 2288 5 1 1 2287
0 2289 7 4 2 42758 49466
0 2290 7 10 2 39946 40553
0 2291 7 2 2 47762 53058
0 2292 7 1 2 53054 53068
0 2293 5 1 1 2292
0 2294 7 1 2 2288 2293
0 2295 5 1 1 2294
0 2296 7 1 2 41425 2295
0 2297 5 1 1 2296
0 2298 7 9 2 40554 50864
0 2299 5 6 1 53070
0 2300 7 7 2 44732 41881
0 2301 7 8 2 39947 46031
0 2302 7 1 2 51024 53092
0 2303 7 1 2 53085 2302
0 2304 5 1 1 2303
0 2305 7 1 2 53079 2304
0 2306 5 1 1 2305
0 2307 7 1 2 49924 2306
0 2308 5 1 1 2307
0 2309 7 2 2 50996 50527
0 2310 5 2 1 53100
0 2311 7 2 2 49566 53093
0 2312 5 1 1 53104
0 2313 7 1 2 45233 53071
0 2314 5 1 1 2313
0 2315 7 1 2 2312 2314
0 2316 5 1 1 2315
0 2317 7 1 2 53102 2316
0 2318 5 1 1 2317
0 2319 7 1 2 2308 2318
0 2320 5 1 1 2319
0 2321 7 1 2 41072 2320
0 2322 5 1 1 2321
0 2323 7 1 2 2297 2322
0 2324 5 1 1 2323
0 2325 7 1 2 41575 49999
0 2326 7 1 2 2324 2325
0 2327 5 1 1 2326
0 2328 7 1 2 42460 2327
0 2329 7 1 2 2286 2328
0 2330 5 1 1 2329
0 2331 7 1 2 2185 2330
0 2332 5 1 1 2331
0 2333 7 2 2 48538 51780
0 2334 7 1 2 50067 53106
0 2335 5 1 1 2334
0 2336 7 2 2 46032 50712
0 2337 5 1 1 53108
0 2338 7 1 2 52203 53109
0 2339 5 1 1 2338
0 2340 7 1 2 2335 2339
0 2341 5 1 1 2340
0 2342 7 1 2 44879 2341
0 2343 5 1 1 2342
0 2344 7 3 2 46033 47699
0 2345 7 1 2 48539 53110
0 2346 7 1 2 51733 2345
0 2347 5 1 1 2346
0 2348 7 1 2 53080 2347
0 2349 5 1 1 2348
0 2350 7 1 2 50635 2349
0 2351 5 1 1 2350
0 2352 7 1 2 2343 2351
0 2353 5 1 1 2352
0 2354 7 1 2 46201 2353
0 2355 5 1 1 2354
0 2356 7 1 2 50000 49074
0 2357 7 1 2 53107 2356
0 2358 5 1 1 2357
0 2359 7 1 2 2355 2358
0 2360 5 1 1 2359
0 2361 7 1 2 42251 2360
0 2362 5 1 1 2361
0 2363 7 3 2 41576 47846
0 2364 5 2 1 53113
0 2365 7 1 2 50001 53114
0 2366 5 1 1 2365
0 2367 7 2 2 45581 52631
0 2368 7 2 2 49361 53118
0 2369 5 1 1 53120
0 2370 7 1 2 52766 2369
0 2371 5 1 1 2370
0 2372 7 1 2 51878 2371
0 2373 5 1 1 2372
0 2374 7 1 2 2366 2373
0 2375 5 1 1 2374
0 2376 7 1 2 47311 2375
0 2377 5 1 1 2376
0 2378 7 6 2 45012 48321
0 2379 5 1 1 53122
0 2380 7 1 2 50014 2379
0 2381 5 5 1 2380
0 2382 7 1 2 47214 53128
0 2383 5 1 1 2382
0 2384 7 11 2 41882 46034
0 2385 7 5 2 44880 53133
0 2386 5 1 1 53144
0 2387 7 1 2 52889 53145
0 2388 7 1 2 52874 2387
0 2389 5 1 1 2388
0 2390 7 1 2 2383 2389
0 2391 5 1 1 2390
0 2392 7 1 2 51815 2391
0 2393 5 1 1 2392
0 2394 7 2 2 40156 50713
0 2395 5 4 1 53149
0 2396 7 1 2 41176 50714
0 2397 5 2 1 2396
0 2398 7 2 2 53151 53155
0 2399 5 1 1 53157
0 2400 7 1 2 51079 2399
0 2401 5 2 1 2400
0 2402 7 1 2 52768 53159
0 2403 5 1 1 2402
0 2404 7 4 2 41706 42034
0 2405 7 2 2 41577 53161
0 2406 7 1 2 48571 53165
0 2407 5 1 1 2406
0 2408 7 3 2 41177 52725
0 2409 5 2 1 53167
0 2410 7 12 2 51863 53170
0 2411 7 1 2 53172 53121
0 2412 5 1 1 2411
0 2413 7 1 2 2407 2412
0 2414 7 1 2 2403 2413
0 2415 7 1 2 2393 2414
0 2416 7 1 2 2377 2415
0 2417 5 1 1 2416
0 2418 7 1 2 48453 2417
0 2419 5 1 1 2418
0 2420 7 1 2 2362 2419
0 2421 5 1 1 2420
0 2422 7 1 2 45801 2421
0 2423 5 1 1 2422
0 2424 7 8 2 41426 42252
0 2425 7 2 2 42461 53184
0 2426 5 1 1 53192
0 2427 7 1 2 53193 52891
0 2428 5 1 1 2427
0 2429 7 1 2 2423 2428
0 2430 5 1 1 2429
0 2431 7 1 2 48721 2430
0 2432 5 1 1 2431
0 2433 7 1 2 40724 2432
0 2434 7 1 2 2332 2433
0 2435 5 1 1 2434
0 2436 7 1 2 1910 2435
0 2437 5 1 1 2436
0 2438 7 1 2 40904 2437
0 2439 5 1 1 2438
0 2440 7 4 2 52493 48777
0 2441 5 3 1 53194
0 2442 7 1 2 52485 53198
0 2443 5 1 1 2442
0 2444 7 1 2 49629 2443
0 2445 5 1 1 2444
0 2446 7 18 2 44733 45802
0 2447 5 3 1 53201
0 2448 7 1 2 53202 50493
0 2449 5 2 1 2448
0 2450 7 1 2 2445 53222
0 2451 5 1 1 2450
0 2452 7 1 2 49176 2451
0 2453 5 1 1 2452
0 2454 7 17 2 45389 45803
0 2455 5 1 1 53224
0 2456 7 5 2 44881 45582
0 2457 7 2 2 53225 53241
0 2458 5 1 1 53246
0 2459 7 7 2 41178 41427
0 2460 7 17 2 40555 43996
0 2461 7 1 2 53248 53255
0 2462 7 1 2 53247 2461
0 2463 5 1 1 2462
0 2464 7 1 2 2453 2463
0 2465 5 1 1 2464
0 2466 7 1 2 41707 2465
0 2467 5 1 1 2466
0 2468 7 27 2 41428 45804
0 2469 5 2 1 53272
0 2470 7 7 2 45013 45390
0 2471 7 2 2 53273 53301
0 2472 7 6 2 40725 45583
0 2473 7 10 2 40556 41179
0 2474 7 1 2 41578 53316
0 2475 7 1 2 53310 2474
0 2476 7 1 2 53308 2475
0 2477 5 1 1 2476
0 2478 7 1 2 2467 2477
0 2479 5 1 1 2478
0 2480 7 1 2 40328 2479
0 2481 5 1 1 2480
0 2482 7 11 2 40557 51482
0 2483 7 1 2 52432 49849
0 2484 7 1 2 53326 2483
0 2485 5 1 1 2484
0 2486 7 1 2 2481 2485
0 2487 5 1 1 2486
0 2488 7 1 2 41310 2487
0 2489 5 1 1 2488
0 2490 7 9 2 41708 41883
0 2491 7 1 2 48454 53337
0 2492 7 1 2 48427 2491
0 2493 7 1 2 52571 2492
0 2494 5 1 1 2493
0 2495 7 1 2 2489 2494
0 2496 5 1 1 2495
0 2497 7 1 2 48625 2496
0 2498 5 1 1 2497
0 2499 7 1 2 43845 50689
0 2500 5 2 1 2499
0 2501 7 1 2 1653 53346
0 2502 5 1 1 2501
0 2503 7 1 2 42253 2502
0 2504 5 1 1 2503
0 2505 7 1 2 52061 2504
0 2506 5 2 1 2505
0 2507 7 2 2 41429 53348
0 2508 5 1 1 53350
0 2509 7 1 2 42462 53021
0 2510 7 1 2 2508 2509
0 2511 5 1 1 2510
0 2512 7 1 2 48540 51787
0 2513 5 2 1 2512
0 2514 7 1 2 45805 53352
0 2515 5 1 1 2514
0 2516 7 1 2 41579 2515
0 2517 7 1 2 2511 2516
0 2518 5 1 1 2517
0 2519 7 8 2 44882 48455
0 2520 5 2 1 53354
0 2521 7 5 2 39948 45584
0 2522 5 1 1 53364
0 2523 7 2 2 44595 2522
0 2524 5 2 1 53369
0 2525 7 1 2 41073 51945
0 2526 7 1 2 53371 2525
0 2527 5 1 1 2526
0 2528 7 1 2 51943 2527
0 2529 5 1 1 2528
0 2530 7 1 2 45234 2529
0 2531 5 1 1 2530
0 2532 7 1 2 51905 2531
0 2533 5 1 1 2532
0 2534 7 1 2 53355 2533
0 2535 5 1 1 2534
0 2536 7 1 2 2518 2535
0 2537 5 1 1 2536
0 2538 7 1 2 40726 2537
0 2539 5 1 1 2538
0 2540 7 3 2 49630 49177
0 2541 5 1 1 53373
0 2542 7 1 2 40329 1823
0 2543 5 1 1 2542
0 2544 7 2 2 45806 47450
0 2545 7 1 2 50724 53376
0 2546 5 1 1 2545
0 2547 7 1 2 2543 2546
0 2548 5 1 1 2547
0 2549 7 1 2 40157 2548
0 2550 5 1 1 2549
0 2551 7 5 2 41311 41884
0 2552 5 1 1 53378
0 2553 7 2 2 40330 53379
0 2554 5 1 1 53383
0 2555 7 1 2 52572 53384
0 2556 5 1 1 2555
0 2557 7 1 2 2550 2556
0 2558 5 1 1 2557
0 2559 7 1 2 41180 2558
0 2560 5 1 1 2559
0 2561 7 1 2 50037 52479
0 2562 5 1 1 2561
0 2563 7 1 2 2560 2562
0 2564 5 1 1 2563
0 2565 7 1 2 53374 2564
0 2566 5 1 1 2565
0 2567 7 1 2 2539 2566
0 2568 5 1 1 2567
0 2569 7 1 2 41709 2568
0 2570 5 1 1 2569
0 2571 7 1 2 2498 2570
0 2572 5 1 1 2571
0 2573 7 1 2 46035 2572
0 2574 5 1 1 2573
0 2575 7 4 2 41312 52433
0 2576 5 6 1 53385
0 2577 7 2 2 41885 51816
0 2578 5 2 1 53395
0 2579 7 2 2 51896 53397
0 2580 5 3 1 53399
0 2581 7 1 2 42254 53401
0 2582 5 1 1 2581
0 2583 7 1 2 48649 2582
0 2584 5 2 1 2583
0 2585 7 4 2 45585 50715
0 2586 5 4 1 53406
0 2587 7 1 2 53407 53400
0 2588 5 1 1 2587
0 2589 7 1 2 53404 2588
0 2590 5 1 1 2589
0 2591 7 1 2 52719 2590
0 2592 5 3 1 2591
0 2593 7 1 2 45807 53414
0 2594 5 2 1 2593
0 2595 7 1 2 53389 53417
0 2596 5 1 1 2595
0 2597 7 1 2 48456 2596
0 2598 5 1 1 2597
0 2599 7 1 2 49631 52596
0 2600 5 1 1 2599
0 2601 7 6 2 40331 50970
0 2602 7 3 2 53226 48778
0 2603 7 1 2 53419 53425
0 2604 5 1 1 2603
0 2605 7 1 2 2600 2604
0 2606 7 1 2 2598 2605
0 2607 5 1 1 2606
0 2608 7 1 2 41580 2607
0 2609 5 1 1 2608
0 2610 7 10 2 40558 41313
0 2611 7 4 2 50176 53428
0 2612 7 2 2 44883 53438
0 2613 7 1 2 53274 50473
0 2614 7 1 2 53442 2613
0 2615 5 1 1 2614
0 2616 7 1 2 2609 2615
0 2617 5 1 1 2616
0 2618 7 1 2 40727 2617
0 2619 5 1 1 2618
0 2620 7 26 2 45586 45808
0 2621 5 1 1 53444
0 2622 7 9 2 45391 53445
0 2623 7 1 2 43997 51215
0 2624 7 1 2 53470 2623
0 2625 7 1 2 53439 2624
0 2626 5 1 1 2625
0 2627 7 1 2 2619 2626
0 2628 5 1 1 2627
0 2629 7 1 2 50068 2628
0 2630 5 1 1 2629
0 2631 7 1 2 2574 2630
0 2632 5 1 1 2631
0 2633 7 1 2 46202 2632
0 2634 5 1 1 2633
0 2635 7 4 2 48094 53446
0 2636 5 1 1 53479
0 2637 7 3 2 40332 51451
0 2638 7 1 2 53480 53483
0 2639 7 3 2 41710 45392
0 2640 7 2 2 41581 53486
0 2641 7 8 2 41314 41430
0 2642 7 3 2 41181 53491
0 2643 7 1 2 53489 53499
0 2644 7 1 2 2638 2643
0 2645 5 1 1 2644
0 2646 7 1 2 44160 2645
0 2647 7 1 2 2634 2646
0 2648 5 1 1 2647
0 2649 7 1 2 43050 2648
0 2650 7 1 2 2439 2649
0 2651 5 1 1 2650
0 2652 7 2 2 43998 41431
0 2653 7 3 2 40559 53502
0 2654 5 2 1 53504
0 2655 7 8 2 40728 44734
0 2656 5 1 1 53509
0 2657 7 4 2 43846 53510
0 2658 5 3 1 53517
0 2659 7 1 2 53507 53521
0 2660 5 13 1 2659
0 2661 7 13 2 43051 52632
0 2662 7 1 2 48722 53402
0 2663 5 1 1 2662
0 2664 7 1 2 53447 2663
0 2665 7 1 2 52658 2664
0 2666 5 1 1 2665
0 2667 7 1 2 45235 51901
0 2668 5 2 1 2667
0 2669 7 1 2 48650 53550
0 2670 5 1 1 2669
0 2671 7 1 2 50716 2670
0 2672 5 2 1 2671
0 2673 7 9 2 41182 42035
0 2674 5 4 1 53554
0 2675 7 3 2 42036 47451
0 2676 5 2 1 53567
0 2677 7 1 2 45393 51817
0 2678 5 3 1 2677
0 2679 7 2 2 53570 53572
0 2680 7 1 2 53563 53575
0 2681 5 1 1 2680
0 2682 7 1 2 41886 2681
0 2683 5 1 1 2682
0 2684 7 1 2 42255 2683
0 2685 7 1 2 53552 2684
0 2686 5 1 1 2685
0 2687 7 1 2 42463 53000
0 2688 5 1 1 2687
0 2689 7 1 2 2686 2688
0 2690 7 1 2 2666 2689
0 2691 5 1 1 2690
0 2692 7 1 2 1857 52486
0 2693 5 1 1 2692
0 2694 7 1 2 40333 2693
0 2695 5 1 1 2694
0 2696 7 8 2 45236 42464
0 2697 7 1 2 50027 53577
0 2698 5 1 1 2697
0 2699 7 1 2 52487 2698
0 2700 5 1 1 2699
0 2701 7 1 2 40158 2700
0 2702 5 1 1 2701
0 2703 7 1 2 2695 2702
0 2704 7 1 2 2691 2703
0 2705 5 1 1 2704
0 2706 7 1 2 53537 2705
0 2707 5 1 1 2706
0 2708 7 3 2 47763 51119
0 2709 5 2 1 53585
0 2710 7 1 2 48723 53588
0 2711 5 1 1 2710
0 2712 7 1 2 49467 2711
0 2713 5 3 1 2712
0 2714 7 11 2 41887 42465
0 2715 7 14 2 46323 48572
0 2716 7 2 2 51025 53604
0 2717 7 1 2 53593 53618
0 2718 7 1 2 53590 2717
0 2719 5 1 1 2718
0 2720 7 1 2 2707 2719
0 2721 5 1 1 2720
0 2722 7 1 2 41582 2721
0 2723 5 1 1 2722
0 2724 7 45 2 42919 46324
0 2725 7 6 2 44884 53620
0 2726 7 1 2 48037 250
0 2727 5 1 1 2726
0 2728 7 1 2 45587 2727
0 2729 5 1 1 2728
0 2730 7 1 2 2729 269
0 2731 5 1 1 2730
0 2732 7 1 2 51879 2731
0 2733 5 1 1 2732
0 2734 7 4 2 43640 48152
0 2735 5 3 1 53671
0 2736 7 12 2 44596 45588
0 2737 5 5 1 53678
0 2738 7 2 2 50602 53690
0 2739 5 15 1 53695
0 2740 7 2 2 47312 53697
0 2741 7 1 2 41888 53712
0 2742 5 1 1 2741
0 2743 7 1 2 53675 2742
0 2744 5 2 1 2743
0 2745 7 1 2 44473 53714
0 2746 5 1 1 2745
0 2747 7 11 2 41889 47313
0 2748 5 3 1 53716
0 2749 7 2 2 41183 53727
0 2750 5 2 1 53730
0 2751 7 1 2 53698 53732
0 2752 5 1 1 2751
0 2753 7 1 2 40334 47545
0 2754 5 2 1 2753
0 2755 7 1 2 45589 47037
0 2756 7 1 2 47144 2755
0 2757 7 1 2 53734 2756
0 2758 5 1 1 2757
0 2759 7 1 2 2752 2758
0 2760 5 1 1 2759
0 2761 7 1 2 43501 2760
0 2762 5 1 1 2761
0 2763 7 1 2 2746 2762
0 2764 7 4 2 2733 2763
0 2765 5 3 1 53736
0 2766 7 1 2 48805 47186
0 2767 5 2 1 2766
0 2768 7 1 2 53737 53743
0 2769 5 1 1 2768
0 2770 7 1 2 45809 2769
0 2771 5 1 1 2770
0 2772 7 5 2 44597 51909
0 2773 5 7 1 53745
0 2774 7 1 2 53390 53750
0 2775 5 26 1 2774
0 2776 7 3 2 40335 53757
0 2777 5 6 1 53783
0 2778 7 1 2 52018 51675
0 2779 5 4 1 2778
0 2780 7 2 2 42466 53792
0 2781 5 2 1 53796
0 2782 7 1 2 53751 53798
0 2783 5 1 1 2782
0 2784 7 1 2 48626 2783
0 2785 5 1 1 2784
0 2786 7 1 2 53786 2785
0 2787 7 1 2 2771 2786
0 2788 5 2 1 2787
0 2789 7 1 2 42759 53800
0 2790 5 1 1 2789
0 2791 7 43 2 42467 46036
0 2792 5 3 1 53802
0 2793 7 5 2 42037 53803
0 2794 7 2 2 50318 53848
0 2795 7 5 2 47314 49932
0 2796 5 1 1 53855
0 2797 7 1 2 53853 53856
0 2798 5 1 1 2797
0 2799 7 1 2 2790 2798
0 2800 5 1 1 2799
0 2801 7 1 2 53665 2800
0 2802 5 1 1 2801
0 2803 7 1 2 2723 2802
0 2804 5 1 1 2803
0 2805 7 1 2 48991 2804
0 2806 5 1 1 2805
0 2807 7 74 2 40905 41711
0 2808 5 1 1 53860
0 2809 7 89 2 43052 53861
0 2810 5 8 1 53934
0 2811 7 1 2 53799 53418
0 2812 5 1 1 2811
0 2813 7 1 2 53935 2812
0 2814 5 1 1 2813
0 2815 7 2 2 49871 47541
0 2816 5 1 1 54031
0 2817 7 1 2 42038 54032
0 2818 5 1 1 2817
0 2819 7 1 2 50309 2818
0 2820 5 1 1 2819
0 2821 7 1 2 45590 2820
0 2822 5 1 1 2821
0 2823 7 14 2 43641 42039
0 2824 5 4 1 54033
0 2825 7 1 2 50042 54047
0 2826 5 1 1 2825
0 2827 7 1 2 45591 2826
0 2828 5 1 1 2827
0 2829 7 1 2 53717 51831
0 2830 5 1 1 2829
0 2831 7 1 2 2828 2830
0 2832 5 1 1 2831
0 2833 7 1 2 47617 2832
0 2834 5 1 1 2833
0 2835 7 1 2 42256 46975
0 2836 5 1 1 2835
0 2837 7 3 2 45592 47764
0 2838 5 7 1 54051
0 2839 7 1 2 44598 54054
0 2840 7 1 2 2836 2839
0 2841 5 1 1 2840
0 2842 7 1 2 47700 50576
0 2843 5 4 1 2842
0 2844 7 1 2 45810 54061
0 2845 7 1 2 2841 2844
0 2846 7 1 2 2834 2845
0 2847 7 1 2 2822 2846
0 2848 5 1 1 2847
0 2849 7 17 2 45014 46325
0 2850 7 27 2 44161 54065
0 2851 7 1 2 48627 53793
0 2852 5 1 1 2851
0 2853 7 5 2 45593 48651
0 2854 5 14 1 54109
0 2855 7 2 2 42468 54114
0 2856 7 1 2 2852 54128
0 2857 5 1 1 2856
0 2858 7 1 2 54082 2857
0 2859 7 1 2 2848 2858
0 2860 5 1 1 2859
0 2861 7 1 2 2814 2860
0 2862 5 1 1 2861
0 2863 7 1 2 48260 2862
0 2864 5 1 1 2863
0 2865 7 77 2 46326 48887
0 2866 5 1 1 54130
0 2867 7 2 2 45237 51880
0 2868 7 1 2 48187 54207
0 2869 5 1 1 2868
0 2870 7 5 2 45394 47618
0 2871 7 1 2 48248 54209
0 2872 5 1 1 2871
0 2873 7 1 2 2869 2872
0 2874 5 1 1 2873
0 2875 7 1 2 42257 2874
0 2876 5 1 1 2875
0 2877 7 5 2 42920 50756
0 2878 7 5 2 41583 42040
0 2879 7 2 2 44599 54219
0 2880 7 1 2 54214 54224
0 2881 5 1 1 2880
0 2882 7 1 2 2876 2881
0 2883 5 1 1 2882
0 2884 7 1 2 47378 2883
0 2885 5 2 1 2884
0 2886 7 5 2 39949 44600
0 2887 7 1 2 54228 48408
0 2888 5 1 1 2887
0 2889 7 1 2 54226 2888
0 2890 5 1 1 2889
0 2891 7 1 2 45811 2890
0 2892 5 1 1 2891
0 2893 7 2 2 45812 50260
0 2894 7 1 2 44601 48095
0 2895 7 1 2 54233 2894
0 2896 5 3 1 2895
0 2897 7 1 2 43306 54235
0 2898 5 1 1 2897
0 2899 7 1 2 41184 52434
0 2900 7 5 2 44885 45238
0 2901 7 3 2 48202 54238
0 2902 5 1 1 54243
0 2903 7 1 2 2899 54244
0 2904 5 1 1 2903
0 2905 7 1 2 54236 2904
0 2906 5 3 1 2905
0 2907 7 1 2 41074 54246
0 2908 7 1 2 2898 2907
0 2909 5 1 1 2908
0 2910 7 1 2 40159 54247
0 2911 5 2 1 2910
0 2912 7 7 2 41185 42469
0 2913 7 4 2 50273 54251
0 2914 5 1 1 54258
0 2915 7 1 2 54259 54245
0 2916 5 1 1 2915
0 2917 7 1 2 54249 2916
0 2918 7 1 2 2909 2917
0 2919 7 1 2 2892 2918
0 2920 5 1 1 2919
0 2921 7 1 2 54131 2920
0 2922 5 1 1 2921
0 2923 7 1 2 2864 2922
0 2924 7 1 2 2806 2923
0 2925 5 1 1 2924
0 2926 7 1 2 53524 2925
0 2927 5 1 1 2926
0 2928 7 25 2 44735 42470
0 2929 5 2 1 54262
0 2930 7 7 2 40729 54263
0 2931 5 3 1 54289
0 2932 7 1 2 54290 51209
0 2933 5 1 1 2932
0 2934 7 4 2 45813 47701
0 2935 7 3 2 43999 48153
0 2936 7 1 2 54299 54303
0 2937 5 1 1 2936
0 2938 7 1 2 2933 2937
0 2939 5 1 1 2938
0 2940 7 1 2 43847 2939
0 2941 5 1 1 2940
0 2942 7 22 2 41432 42471
0 2943 5 8 1 54306
0 2944 7 2 2 53219 54328
0 2945 5 38 1 54336
0 2946 7 2 2 45594 54338
0 2947 7 1 2 44000 51704
0 2948 7 1 2 54376 2947
0 2949 5 1 1 2948
0 2950 7 1 2 2941 2949
0 2951 5 1 1 2950
0 2952 7 1 2 47908 2951
0 2953 5 1 1 2952
0 2954 7 18 2 45814 48541
0 2955 5 1 1 54378
0 2956 7 1 2 54329 2955
0 2957 5 23 1 2956
0 2958 7 2 2 44001 54396
0 2959 5 1 1 54419
0 2960 7 1 2 54208 54420
0 2961 5 1 1 2960
0 2962 7 16 2 42041 42472
0 2963 7 16 2 43848 40730
0 2964 7 8 2 44736 54437
0 2965 5 1 1 54453
0 2966 7 1 2 54421 54454
0 2967 5 1 1 2966
0 2968 7 1 2 2961 2967
0 2969 5 1 1 2968
0 2970 7 1 2 47379 2969
0 2971 5 1 1 2970
0 2972 7 3 2 54264 54438
0 2973 5 3 1 54461
0 2974 7 1 2 53173 54462
0 2975 5 1 1 2974
0 2976 7 1 2 2971 2975
0 2977 5 1 1 2976
0 2978 7 1 2 42258 2977
0 2979 5 1 1 2978
0 2980 7 1 2 2953 2979
0 2981 5 1 1 2980
0 2982 7 1 2 44602 2981
0 2983 5 1 1 2982
0 2984 7 11 2 44002 45815
0 2985 7 1 2 45239 54467
0 2986 5 1 1 2985
0 2987 7 1 2 54296 2986
0 2988 5 1 1 2987
0 2989 7 1 2 43849 2988
0 2990 5 1 1 2989
0 2991 7 5 2 44003 45240
0 2992 5 1 1 54478
0 2993 7 1 2 54339 54479
0 2994 5 1 1 2993
0 2995 7 1 2 2990 2994
0 2996 5 1 1 2995
0 2997 7 2 2 51026 2996
0 2998 7 1 2 52799 54483
0 2999 5 1 1 2998
0 3000 7 1 2 2983 2999
0 3001 5 1 1 3000
0 3002 7 1 2 43642 3001
0 3003 5 1 1 3002
0 3004 7 1 2 48040 54484
0 3005 5 1 1 3004
0 3006 7 1 2 3003 3005
0 3007 5 1 1 3006
0 3008 7 1 2 41712 3007
0 3009 5 1 1 3008
0 3010 7 23 2 40731 42473
0 3011 5 5 1 54485
0 3012 7 3 2 44004 53275
0 3013 5 3 1 54513
0 3014 7 1 2 54508 54516
0 3015 5 1 1 3014
0 3016 7 1 2 40560 3015
0 3017 5 1 1 3016
0 3018 7 1 2 40732 54340
0 3019 5 1 1 3018
0 3020 7 1 2 3017 3019
0 3021 5 4 1 3020
0 3022 7 1 2 49100 54519
0 3023 5 1 1 3022
0 3024 7 1 2 48867 51444
0 3025 7 1 2 54397 3024
0 3026 7 1 2 48799 3025
0 3027 5 1 1 3026
0 3028 7 1 2 3023 3027
0 3029 5 1 1 3028
0 3030 7 1 2 45395 3029
0 3031 5 1 1 3030
0 3032 7 1 2 3009 3031
0 3033 5 1 1 3032
0 3034 7 1 2 42921 3033
0 3035 5 1 1 3034
0 3036 7 1 2 47380 53518
0 3037 5 1 1 3036
0 3038 7 2 2 47315 53525
0 3039 7 1 2 41890 54523
0 3040 5 1 1 3039
0 3041 7 1 2 3037 3040
0 3042 5 1 1 3041
0 3043 7 1 2 49933 3042
0 3044 5 1 1 3043
0 3045 7 1 2 51753 53526
0 3046 5 1 1 3045
0 3047 7 1 2 3044 3046
0 3048 5 1 1 3047
0 3049 7 12 2 42259 42474
0 3050 7 7 2 42042 54525
0 3051 7 1 2 54537 49975
0 3052 7 1 2 3048 3051
0 3053 5 1 1 3052
0 3054 7 1 2 3035 3053
0 3055 5 1 1 3054
0 3056 7 1 2 46327 3055
0 3057 5 1 1 3056
0 3058 7 11 2 43053 52854
0 3059 5 2 1 54544
0 3060 7 2 2 54486 54545
0 3061 7 5 2 41433 53317
0 3062 7 8 2 40336 45396
0 3063 5 5 1 54564
0 3064 7 1 2 54559 54565
0 3065 7 1 2 54557 3064
0 3066 5 1 1 3065
0 3067 7 1 2 3057 3066
0 3068 5 1 1 3067
0 3069 7 1 2 44162 3068
0 3070 5 1 1 3069
0 3071 7 11 2 44163 46328
0 3072 7 1 2 42922 54577
0 3073 7 1 2 53801 3072
0 3074 5 1 1 3073
0 3075 7 41 2 46203 43054
0 3076 7 1 2 42475 54588
0 3077 7 5 2 40906 41186
0 3078 7 1 2 54566 54629
0 3079 7 1 2 3076 3078
0 3080 5 1 1 3079
0 3081 7 1 2 3074 3080
0 3082 5 1 1 3081
0 3083 7 1 2 51479 3082
0 3084 5 1 1 3083
0 3085 7 5 2 41713 54589
0 3086 5 2 1 54634
0 3087 7 1 2 52390 54635
0 3088 5 1 1 3087
0 3089 7 4 2 40337 46329
0 3090 7 1 2 54641 52862
0 3091 5 1 1 3090
0 3092 7 1 2 3088 3091
0 3093 5 1 1 3092
0 3094 7 1 2 39950 3093
0 3095 5 1 1 3094
0 3096 7 15 2 40160 40338
0 3097 5 1 1 54645
0 3098 7 3 2 42923 54646
0 3099 7 1 2 54066 54660
0 3100 5 1 1 3099
0 3101 7 1 2 3095 3100
0 3102 5 1 1 3101
0 3103 7 1 2 41187 3102
0 3104 5 1 1 3103
0 3105 7 1 2 54636 52827
0 3106 5 1 1 3105
0 3107 7 1 2 3104 3106
0 3108 5 1 1 3107
0 3109 7 1 2 45397 3108
0 3110 5 1 1 3109
0 3111 7 9 2 46330 52863
0 3112 7 4 2 43643 48611
0 3113 5 1 1 54672
0 3114 7 1 2 51985 3113
0 3115 7 1 2 54663 3114
0 3116 5 1 1 3115
0 3117 7 1 2 3110 3116
0 3118 5 1 1 3117
0 3119 7 1 2 43850 3118
0 3120 5 1 1 3119
0 3121 7 14 2 41714 43055
0 3122 7 2 2 54676 48322
0 3123 5 2 1 54690
0 3124 7 3 2 51027 49468
0 3125 5 1 1 54694
0 3126 7 1 2 52566 54695
0 3127 7 1 2 54691 3126
0 3128 5 1 1 3127
0 3129 7 1 2 3120 3128
0 3130 5 1 1 3129
0 3131 7 1 2 42476 3130
0 3132 5 1 1 3131
0 3133 7 11 2 45241 47381
0 3134 5 1 1 54697
0 3135 7 1 2 51028 54698
0 3136 5 1 1 3135
0 3137 7 1 2 50667 3136
0 3138 5 1 1 3137
0 3139 7 1 2 48724 3138
0 3140 5 1 1 3139
0 3141 7 2 2 40561 49469
0 3142 5 4 1 54708
0 3143 7 1 2 50603 1088
0 3144 5 2 1 3143
0 3145 7 1 2 54710 54714
0 3146 5 1 1 3145
0 3147 7 1 2 3140 3146
0 3148 5 1 1 3147
0 3149 7 1 2 47702 3148
0 3150 5 1 1 3149
0 3151 7 5 2 43307 50888
0 3152 5 2 1 54716
0 3153 7 1 2 48806 54717
0 3154 5 1 1 3153
0 3155 7 1 2 43851 48020
0 3156 5 1 1 3155
0 3157 7 1 2 3154 3156
0 3158 5 1 1 3157
0 3159 7 1 2 43644 3158
0 3160 5 1 1 3159
0 3161 7 7 2 43308 43852
0 3162 7 1 2 47979 53691
0 3163 5 4 1 3162
0 3164 7 2 2 44394 54730
0 3165 5 1 1 54734
0 3166 7 1 2 54723 54735
0 3167 5 1 1 3166
0 3168 7 1 2 3160 3167
0 3169 5 1 1 3168
0 3170 7 1 2 51881 3169
0 3171 5 1 1 3170
0 3172 7 2 2 44603 52680
0 3173 5 2 1 54736
0 3174 7 1 2 53031 54737
0 3175 5 1 1 3174
0 3176 7 1 2 43853 53715
0 3177 5 1 1 3176
0 3178 7 3 2 50577 49402
0 3179 5 1 1 54740
0 3180 7 1 2 54741 53718
0 3181 5 1 1 3180
0 3182 7 1 2 3177 3181
0 3183 5 1 1 3182
0 3184 7 1 2 47619 3183
0 3185 5 1 1 3184
0 3186 7 1 2 3175 3185
0 3187 7 1 2 3171 3186
0 3188 7 1 2 3150 3187
0 3189 5 1 1 3188
0 3190 7 1 2 53621 52162
0 3191 7 1 2 3189 3190
0 3192 5 1 1 3191
0 3193 7 1 2 3132 3192
0 3194 5 1 1 3193
0 3195 7 1 2 44737 3194
0 3196 5 1 1 3195
0 3197 7 2 2 43309 48725
0 3198 5 2 1 54743
0 3199 7 12 2 42043 47703
0 3200 5 5 1 54747
0 3201 7 2 2 50889 54748
0 3202 5 2 1 54764
0 3203 7 2 2 51882 50901
0 3204 7 1 2 49403 54768
0 3205 5 1 1 3204
0 3206 7 1 2 54766 3205
0 3207 5 1 1 3206
0 3208 7 1 2 54744 3207
0 3209 5 1 1 3208
0 3210 7 3 2 45398 49331
0 3211 5 1 1 54770
0 3212 7 1 2 49404 54771
0 3213 5 1 1 3212
0 3214 7 1 2 3209 3213
0 3215 5 1 1 3214
0 3216 7 1 2 42260 3215
0 3217 5 1 1 3216
0 3218 7 12 2 41891 45595
0 3219 5 6 1 54773
0 3220 7 6 2 44474 48367
0 3221 5 2 1 54791
0 3222 7 9 2 44604 42044
0 3223 5 3 1 54799
0 3224 7 5 2 43645 54800
0 3225 5 1 1 54811
0 3226 7 2 2 54792 54812
0 3227 7 1 2 54774 54816
0 3228 5 1 1 3227
0 3229 7 1 2 3217 3228
0 3230 5 1 1 3229
0 3231 7 14 2 43854 45816
0 3232 5 3 1 54818
0 3233 7 2 2 54330 54832
0 3234 5 4 1 54835
0 3235 7 1 2 54067 54837
0 3236 7 1 2 3230 3235
0 3237 5 1 1 3236
0 3238 7 9 2 41188 41315
0 3239 7 4 2 40339 48457
0 3240 7 2 2 54841 54850
0 3241 7 10 2 41715 45817
0 3242 7 2 2 43056 54856
0 3243 7 1 2 50474 54866
0 3244 7 1 2 54854 3243
0 3245 5 1 1 3244
0 3246 7 1 2 3237 3245
0 3247 5 1 1 3246
0 3248 7 1 2 42924 3247
0 3249 5 1 1 3248
0 3250 7 10 2 42477 46204
0 3251 7 6 2 41434 41716
0 3252 7 2 2 43057 54878
0 3253 7 3 2 54868 54884
0 3254 5 1 1 54886
0 3255 7 1 2 43502 47199
0 3256 5 2 1 3255
0 3257 7 1 2 1535 54889
0 3258 5 3 1 3257
0 3259 7 1 2 52048 54891
0 3260 5 2 1 3259
0 3261 7 2 2 49405 52086
0 3262 5 1 1 54896
0 3263 7 1 2 42261 54897
0 3264 5 1 1 3263
0 3265 7 1 2 54894 3264
0 3266 5 1 1 3265
0 3267 7 1 2 43310 3266
0 3268 5 1 1 3267
0 3269 7 2 2 44605 47064
0 3270 5 4 1 54898
0 3271 7 1 2 47565 54899
0 3272 5 2 1 3271
0 3273 7 1 2 53347 54904
0 3274 5 1 1 3273
0 3275 7 1 2 42262 3274
0 3276 5 1 1 3275
0 3277 7 1 2 3268 3276
0 3278 5 1 1 3277
0 3279 7 1 2 54887 3278
0 3280 5 1 1 3279
0 3281 7 3 2 46828 48726
0 3282 5 3 1 54906
0 3283 7 1 2 47038 50917
0 3284 5 3 1 3283
0 3285 7 1 2 1061 54912
0 3286 5 1 1 3285
0 3287 7 1 2 3286 54888
0 3288 5 1 1 3287
0 3289 7 7 2 45015 45596
0 3290 7 4 2 53622 54915
0 3291 5 1 1 54922
0 3292 7 2 2 43311 54923
0 3293 5 1 1 54926
0 3294 7 1 2 54838 54927
0 3295 5 1 1 3294
0 3296 7 1 2 3254 3295
0 3297 5 1 1 3296
0 3298 7 1 2 47080 3297
0 3299 5 1 1 3298
0 3300 7 8 2 42263 46205
0 3301 7 2 2 54677 54928
0 3302 5 2 1 54936
0 3303 7 1 2 54307 54937
0 3304 5 1 1 3303
0 3305 7 1 2 3299 3304
0 3306 5 1 1 3305
0 3307 7 1 2 50254 3306
0 3308 5 1 1 3307
0 3309 7 1 2 3288 3308
0 3310 5 1 1 3309
0 3311 7 1 2 54907 3310
0 3312 5 1 1 3311
0 3313 7 1 2 44005 3312
0 3314 7 1 2 3280 3313
0 3315 7 1 2 3249 3314
0 3316 7 1 2 3196 3315
0 3317 5 1 1 3316
0 3318 7 1 2 50630 52122
0 3319 5 1 1 3318
0 3320 7 2 2 48458 51986
0 3321 5 1 1 54940
0 3322 7 6 2 42264 48542
0 3323 5 1 1 54942
0 3324 7 4 2 3323 475
0 3325 7 1 2 52981 54948
0 3326 5 1 1 3325
0 3327 7 1 2 3321 3326
0 3328 5 1 1 3327
0 3329 7 1 2 42925 3328
0 3330 5 1 1 3329
0 3331 7 1 2 3319 3330
0 3332 5 1 1 3331
0 3333 7 1 2 54678 3332
0 3334 5 1 1 3333
0 3335 7 3 2 42265 51818
0 3336 5 1 1 54952
0 3337 7 1 2 51803 54953
0 3338 5 1 1 3337
0 3339 7 1 2 51211 3338
0 3340 5 1 1 3339
0 3341 7 1 2 49406 3340
0 3342 5 1 1 3341
0 3343 7 4 2 44475 51029
0 3344 7 2 2 49760 54955
0 3345 5 1 1 54959
0 3346 7 1 2 3342 3345
0 3347 5 1 1 3346
0 3348 7 3 2 43855 48727
0 3349 5 4 1 54961
0 3350 7 2 2 44738 54962
0 3351 5 5 1 54968
0 3352 7 1 2 54664 54969
0 3353 7 1 2 3347 3352
0 3354 5 1 1 3353
0 3355 7 1 2 3334 3354
0 3356 5 1 1 3355
0 3357 7 1 2 42478 3356
0 3358 5 1 1 3357
0 3359 7 15 2 42926 43058
0 3360 7 4 2 54857 54975
0 3361 7 1 2 48459 52049
0 3362 5 1 1 3361
0 3363 7 10 2 44739 45597
0 3364 7 3 2 41316 54994
0 3365 5 2 1 55004
0 3366 7 2 2 50177 55005
0 3367 5 1 1 55009
0 3368 7 1 2 45399 55010
0 3369 5 2 1 3368
0 3370 7 1 2 3362 55011
0 3371 5 1 1 3370
0 3372 7 1 2 54990 3371
0 3373 5 1 1 3372
0 3374 7 1 2 40733 3373
0 3375 7 1 2 3358 3374
0 3376 5 1 1 3375
0 3377 7 1 2 40907 3376
0 3378 7 1 2 3317 3377
0 3379 5 1 1 3378
0 3380 7 1 2 3084 3379
0 3381 7 1 2 3070 3380
0 3382 5 1 1 3381
0 3383 7 1 2 52899 3382
0 3384 5 1 1 3383
0 3385 7 1 2 2927 3384
0 3386 7 1 2 2651 3385
0 3387 7 1 2 1510 3386
0 3388 5 1 1 3387
0 3389 7 1 2 46603 3388
0 3390 5 1 1 3389
0 3391 7 3 2 44223 41772
0 3392 5 1 1 55013
0 3393 7 7 2 40973 45066
0 3394 5 1 1 55016
0 3395 7 5 2 3392 3394
0 3396 5 107 1 55023
0 3397 7 8 2 43503 41892
0 3398 5 2 1 55135
0 3399 7 9 2 55136 47382
0 3400 5 8 1 55145
0 3401 7 4 2 48047 48992
0 3402 5 1 1 55162
0 3403 7 12 2 44006 40908
0 3404 7 9 2 55166 49850
0 3405 5 1 1 55178
0 3406 7 1 2 3402 3405
0 3407 5 7 1 3406
0 3408 7 1 2 46037 52619
0 3409 5 3 1 3408
0 3410 7 8 2 42479 48203
0 3411 5 2 1 55197
0 3412 7 1 2 55194 55205
0 3413 5 2 1 3412
0 3414 7 1 2 52976 55207
0 3415 5 1 1 3414
0 3416 7 8 2 42480 51987
0 3417 5 1 1 55209
0 3418 7 1 2 48204 55210
0 3419 5 1 1 3418
0 3420 7 1 2 3415 3419
0 3421 5 1 1 3420
0 3422 7 1 2 55187 3421
0 3423 5 1 1 3422
0 3424 7 2 2 53804 51988
0 3425 5 1 1 55217
0 3426 7 45 2 45818 42760
0 3427 5 1 1 55219
0 3428 7 1 2 55220 51989
0 3429 5 4 1 3428
0 3430 7 1 2 53845 55264
0 3431 5 3 1 3430
0 3432 7 1 2 51671 55268
0 3433 5 1 1 3432
0 3434 7 1 2 3425 3433
0 3435 5 1 1 3434
0 3436 7 1 2 49178 3435
0 3437 5 1 1 3436
0 3438 7 7 2 40734 47215
0 3439 5 3 1 55271
0 3440 7 1 2 55272 53797
0 3441 5 1 1 3440
0 3442 7 1 2 3437 3441
0 3443 5 1 1 3442
0 3444 7 1 2 40909 50002
0 3445 7 1 2 3443 3444
0 3446 5 1 1 3445
0 3447 7 1 2 3423 3446
0 3448 5 1 1 3447
0 3449 7 1 2 41435 3448
0 3450 5 1 1 3449
0 3451 7 3 2 40735 46661
0 3452 5 2 1 55281
0 3453 7 8 2 44007 49075
0 3454 5 1 1 55286
0 3455 7 1 2 3454 55278
0 3456 7 1 2 55284 3455
0 3457 5 12 1 3456
0 3458 7 4 2 42927 55294
0 3459 5 1 1 55306
0 3460 7 12 2 40340 42481
0 3461 7 2 2 55310 50274
0 3462 5 1 1 55322
0 3463 7 12 2 41717 45598
0 3464 7 1 2 55324 54630
0 3465 7 1 2 55323 3464
0 3466 7 1 2 55307 3465
0 3467 5 1 1 3466
0 3468 7 1 2 3450 3467
0 3469 5 1 1 3468
0 3470 7 1 2 40562 3469
0 3471 5 1 1 3470
0 3472 7 12 2 42482 49567
0 3473 5 1 1 55336
0 3474 7 2 2 55337 48302
0 3475 5 1 1 55348
0 3476 7 1 2 51990 55349
0 3477 5 1 1 3476
0 3478 7 6 2 43856 42483
0 3479 5 1 1 55350
0 3480 7 3 2 48205 55351
0 3481 5 1 1 55356
0 3482 7 1 2 44740 55357
0 3483 5 2 1 3482
0 3484 7 2 2 54341 51991
0 3485 5 1 1 55361
0 3486 7 1 2 48096 55362
0 3487 5 1 1 3486
0 3488 7 1 2 55359 3487
0 3489 5 1 1 3488
0 3490 7 1 2 49179 3489
0 3491 5 1 1 3490
0 3492 7 21 2 42928 48048
0 3493 5 2 1 55363
0 3494 7 8 2 54265 49962
0 3495 5 3 1 55386
0 3496 7 6 2 42761 54342
0 3497 5 1 1 55397
0 3498 7 1 2 51992 55398
0 3499 5 1 1 3498
0 3500 7 1 2 55394 3499
0 3501 5 1 1 3500
0 3502 7 1 2 55364 3501
0 3503 5 1 1 3502
0 3504 7 1 2 3491 3503
0 3505 5 1 1 3504
0 3506 7 1 2 52977 3505
0 3507 5 1 1 3506
0 3508 7 1 2 3477 3507
0 3509 5 1 1 3508
0 3510 7 1 2 53862 3509
0 3511 5 1 1 3510
0 3512 7 1 2 3471 3511
0 3513 5 1 1 3512
0 3514 7 1 2 46331 3513
0 3515 5 1 1 3514
0 3516 7 12 2 45819 46038
0 3517 7 10 2 55403 54590
0 3518 7 9 2 40563 40910
0 3519 7 3 2 55425 51483
0 3520 7 4 2 41584 45400
0 3521 7 1 2 55325 55437
0 3522 7 1 2 52582 3521
0 3523 7 2 2 55434 3522
0 3524 7 1 2 55415 55441
0 3525 5 1 1 3524
0 3526 7 1 2 3515 3525
0 3527 5 1 1 3526
0 3528 7 1 2 55154 3527
0 3529 5 1 1 3528
0 3530 7 2 2 40341 47987
0 3531 5 2 1 55443
0 3532 7 3 2 40161 54842
0 3533 5 1 1 55447
0 3534 7 1 2 55445 3533
0 3535 5 1 1 3534
0 3536 7 1 2 47512 3535
0 3537 5 1 1 3536
0 3538 7 1 2 50556 51672
0 3539 5 1 1 3538
0 3540 7 1 2 3537 3539
0 3541 5 1 1 3540
0 3542 7 1 2 42484 3541
0 3543 5 1 1 3542
0 3544 7 16 2 44606 45820
0 3545 7 1 2 55450 50170
0 3546 5 1 1 3545
0 3547 7 1 2 42266 3546
0 3548 7 1 2 3543 3547
0 3549 5 1 1 3548
0 3550 7 7 2 41893 45821
0 3551 7 2 2 44607 55466
0 3552 5 2 1 55473
0 3553 7 1 2 41317 52494
0 3554 5 1 1 3553
0 3555 7 1 2 55475 3554
0 3556 5 1 1 3555
0 3557 7 1 2 43646 3556
0 3558 5 1 1 3557
0 3559 7 6 2 39951 50028
0 3560 5 1 1 55477
0 3561 7 1 2 53594 55478
0 3562 5 1 1 3561
0 3563 7 1 2 45599 3562
0 3564 7 1 2 3558 3563
0 3565 5 1 1 3564
0 3566 7 1 2 46039 3565
0 3567 7 1 2 3549 3566
0 3568 5 1 1 3567
0 3569 7 3 2 52088 49949
0 3570 5 8 1 55483
0 3571 7 10 2 45600 47001
0 3572 7 3 2 55221 55494
0 3573 5 2 1 55504
0 3574 7 1 2 48652 55505
0 3575 7 1 2 55486 3574
0 3576 5 1 1 3575
0 3577 7 1 2 3568 3576
0 3578 5 1 1 3577
0 3579 7 1 2 44886 3578
0 3580 5 1 1 3579
0 3581 7 4 2 45601 55222
0 3582 5 1 1 55509
0 3583 7 1 2 53805 48807
0 3584 5 2 1 3583
0 3585 7 1 2 3582 55513
0 3586 5 12 1 3585
0 3587 7 2 2 43312 47856
0 3588 7 1 2 55515 55527
0 3589 5 1 1 3588
0 3590 7 3 2 44887 53448
0 3591 5 2 1 55529
0 3592 7 1 2 53111 55530
0 3593 5 1 1 3592
0 3594 7 1 2 3589 3593
0 3595 5 1 1 3594
0 3596 7 1 2 43647 3595
0 3597 5 1 1 3596
0 3598 7 1 2 51939 51754
0 3599 5 1 1 3598
0 3600 7 1 2 52465 53752
0 3601 5 11 1 3600
0 3602 7 1 2 47513 55534
0 3603 7 1 2 3599 3602
0 3604 5 1 1 3603
0 3605 7 1 2 53787 3604
0 3606 5 1 1 3605
0 3607 7 1 2 46662 3606
0 3608 5 1 1 3607
0 3609 7 1 2 3597 3608
0 3610 5 1 1 3609
0 3611 7 1 2 42045 3610
0 3612 5 2 1 3611
0 3613 7 2 2 52435 50223
0 3614 5 1 1 55547
0 3615 7 1 2 53753 3614
0 3616 5 1 1 3615
0 3617 7 1 2 39952 3616
0 3618 5 1 1 3617
0 3619 7 7 2 45822 48808
0 3620 7 1 2 41075 55549
0 3621 5 1 1 3620
0 3622 7 1 2 54252 51691
0 3623 5 1 1 3622
0 3624 7 1 2 3621 3623
0 3625 7 1 2 3618 3624
0 3626 5 1 1 3625
0 3627 7 1 2 45242 3626
0 3628 5 1 1 3627
0 3629 7 3 2 45823 47263
0 3630 7 1 2 48809 55556
0 3631 5 2 1 3630
0 3632 7 1 2 55559 53788
0 3633 7 1 2 3628 3632
0 3634 5 1 1 3633
0 3635 7 1 2 47216 3634
0 3636 5 1 1 3635
0 3637 7 1 2 55545 3636
0 3638 7 1 2 3580 3637
0 3639 5 1 1 3638
0 3640 7 1 2 41436 3639
0 3641 5 1 1 3640
0 3642 7 3 2 42762 55438
0 3643 5 1 1 55561
0 3644 7 1 2 52317 52702
0 3645 5 1 1 3644
0 3646 7 1 2 3643 3645
0 3647 5 1 1 3646
0 3648 7 1 2 47452 3647
0 3649 5 1 1 3648
0 3650 7 3 2 40162 47217
0 3651 5 1 1 55564
0 3652 7 1 2 50717 55565
0 3653 5 1 1 3652
0 3654 7 7 2 44888 41894
0 3655 7 1 2 51738 53094
0 3656 7 1 2 55567 3655
0 3657 5 1 1 3656
0 3658 7 1 2 3653 3657
0 3659 7 1 2 3649 3658
0 3660 5 1 1 3659
0 3661 7 1 2 45602 3660
0 3662 5 1 1 3661
0 3663 7 7 2 45401 47264
0 3664 5 1 1 55574
0 3665 7 2 2 50103 52789
0 3666 5 1 1 55581
0 3667 7 1 2 55575 55582
0 3668 5 1 1 3667
0 3669 7 1 2 3662 3668
0 3670 5 1 1 3669
0 3671 7 1 2 3670 52591
0 3672 5 2 1 3671
0 3673 7 1 2 3641 55583
0 3674 5 1 1 3673
0 3675 7 1 2 40564 3674
0 3676 5 1 1 3675
0 3677 7 1 2 48460 52738
0 3678 5 1 1 3677
0 3679 7 7 2 42763 49632
0 3680 7 1 2 50367 50793
0 3681 7 1 2 55585 3680
0 3682 5 1 1 3681
0 3683 7 1 2 3678 3682
0 3684 5 1 1 3683
0 3685 7 1 2 42485 3684
0 3686 5 1 1 3685
0 3687 7 1 2 46040 53471
0 3688 7 1 2 47514 51237
0 3689 7 1 2 3687 3688
0 3690 5 1 1 3689
0 3691 7 1 2 3686 3690
0 3692 5 1 1 3691
0 3693 7 1 2 41318 3692
0 3694 5 1 1 3693
0 3695 7 8 2 46041 48461
0 3696 7 9 2 44889 42046
0 3697 7 1 2 52436 55600
0 3698 7 1 2 55592 3697
0 3699 5 1 1 3698
0 3700 7 1 2 3694 3699
0 3701 5 1 1 3700
0 3702 7 1 2 40342 3701
0 3703 5 2 1 3702
0 3704 7 8 2 42764 51910
0 3705 7 1 2 55611 50127
0 3706 5 1 1 3705
0 3707 7 4 2 46042 53758
0 3708 7 2 2 55619 55601
0 3709 5 1 1 55623
0 3710 7 1 2 3706 3709
0 3711 5 1 1 3710
0 3712 7 1 2 48462 3711
0 3713 5 1 1 3712
0 3714 7 1 2 55609 3713
0 3715 5 1 1 3714
0 3716 7 1 2 47765 3715
0 3717 5 1 1 3716
0 3718 7 1 2 51747 52335
0 3719 5 2 1 3718
0 3720 7 2 2 55625 50448
0 3721 7 2 2 39953 55627
0 3722 5 2 1 55629
0 3723 7 4 2 40163 42047
0 3724 7 2 2 46785 55633
0 3725 5 1 1 55637
0 3726 7 1 2 55631 3725
0 3727 5 7 1 3726
0 3728 7 1 2 55639 46663
0 3729 5 1 1 3728
0 3730 7 1 2 45402 55566
0 3731 5 1 1 3730
0 3732 7 1 2 3729 3731
0 3733 5 1 1 3732
0 3734 7 1 2 54343 3733
0 3735 5 1 1 3734
0 3736 7 3 2 45403 55404
0 3737 7 1 2 51238 55646
0 3738 5 1 1 3737
0 3739 7 5 2 50865 51971
0 3740 5 1 1 55649
0 3741 7 1 2 45243 55650
0 3742 5 1 1 3741
0 3743 7 1 2 3738 3742
0 3744 5 1 1 3743
0 3745 7 1 2 40164 3744
0 3746 5 1 1 3745
0 3747 7 4 2 45244 45824
0 3748 7 1 2 44741 55654
0 3749 5 2 1 3748
0 3750 7 1 2 54331 55658
0 3751 5 2 1 3750
0 3752 7 1 2 47453 55660
0 3753 5 1 1 3752
0 3754 7 1 2 53203 47265
0 3755 5 2 1 3754
0 3756 7 1 2 3753 55662
0 3757 5 1 1 3756
0 3758 7 1 2 55562 3757
0 3759 5 1 1 3758
0 3760 7 1 2 3746 3759
0 3761 7 1 2 3735 3760
0 3762 5 1 1 3761
0 3763 7 1 2 45603 3762
0 3764 5 1 1 3763
0 3765 7 18 2 39954 40165
0 3766 5 8 1 55664
0 3767 7 3 2 45404 55665
0 3768 7 1 2 46786 55690
0 3769 7 1 2 55651 3768
0 3770 5 2 1 3769
0 3771 7 1 2 3764 55693
0 3772 5 1 1 3771
0 3773 7 1 2 52583 3772
0 3774 5 1 1 3773
0 3775 7 5 2 44395 42048
0 3776 5 1 1 55695
0 3777 7 2 2 43313 55696
0 3778 5 4 1 55700
0 3779 7 1 2 45604 55702
0 3780 5 2 1 3779
0 3781 7 6 2 51056 55706
0 3782 5 1 1 55708
0 3783 7 1 2 49872 53356
0 3784 5 1 1 3783
0 3785 7 3 2 44476 50128
0 3786 7 1 2 55714 52369
0 3787 5 1 1 3786
0 3788 7 1 2 45825 3787
0 3789 7 1 2 3784 3788
0 3790 5 1 1 3789
0 3791 7 1 2 42486 612
0 3792 5 1 1 3791
0 3793 7 1 2 53134 3792
0 3794 7 1 2 3790 3793
0 3795 5 1 1 3794
0 3796 7 5 2 40565 55223
0 3797 5 1 1 55717
0 3798 7 5 2 43504 41437
0 3799 7 5 2 44477 41585
0 3800 7 1 2 55722 55727
0 3801 7 1 2 55718 3800
0 3802 5 1 1 3801
0 3803 7 1 2 3795 3802
0 3804 5 1 1 3803
0 3805 7 1 2 55709 3804
0 3806 5 2 1 3805
0 3807 7 1 2 3774 55732
0 3808 7 1 2 3717 3807
0 3809 7 1 2 3676 3808
0 3810 5 1 1 3809
0 3811 7 1 2 40736 3810
0 3812 5 1 1 3811
0 3813 7 11 2 42487 49633
0 3814 5 2 1 55734
0 3815 7 1 2 53220 55745
0 3816 5 11 1 3815
0 3817 7 1 2 55640 55747
0 3818 5 1 1 3817
0 3819 7 1 2 43505 47530
0 3820 5 2 1 3819
0 3821 7 1 2 49568 53227
0 3822 7 1 2 55758 3821
0 3823 5 1 1 3822
0 3824 7 1 2 3818 3823
0 3825 5 1 1 3824
0 3826 7 1 2 41189 3825
0 3827 5 1 1 3826
0 3828 7 9 2 40166 43857
0 3829 7 2 2 44742 55760
0 3830 7 1 2 53228 47515
0 3831 7 1 2 55769 3830
0 3832 5 1 1 3831
0 3833 7 1 2 3827 3832
0 3834 5 1 1 3833
0 3835 7 10 2 40343 44008
0 3836 7 2 2 51993 55771
0 3837 7 1 2 49076 55781
0 3838 7 2 2 3834 3837
0 3839 5 1 1 55783
0 3840 7 1 2 3812 3839
0 3841 5 1 1 3840
0 3842 7 1 2 49976 3841
0 3843 5 1 1 3842
0 3844 7 5 2 43648 40737
0 3845 7 5 2 44608 55785
0 3846 7 3 2 43314 45245
0 3847 5 2 1 55795
0 3848 7 2 2 55796 55697
0 3849 5 1 1 55800
0 3850 7 5 2 42765 54526
0 3851 7 1 2 55802 50393
0 3852 7 1 2 55801 3851
0 3853 5 1 1 3852
0 3854 7 2 2 42766 54398
0 3855 5 1 1 55807
0 3856 7 1 2 51057 55808
0 3857 5 1 1 3856
0 3858 7 4 2 46043 53595
0 3859 7 1 2 49569 55809
0 3860 5 1 1 3859
0 3861 7 1 2 3857 3860
0 3862 5 1 1 3861
0 3863 7 1 2 44890 3862
0 3864 5 1 1 3863
0 3865 7 13 2 42488 42767
0 3866 7 1 2 55813 50408
0 3867 5 1 1 3866
0 3868 7 1 2 3864 3867
0 3869 5 1 1 3868
0 3870 7 1 2 47704 55707
0 3871 7 1 2 3869 3870
0 3872 5 1 1 3871
0 3873 7 1 2 3853 3872
0 3874 5 1 1 3873
0 3875 7 1 2 55790 3874
0 3876 5 1 1 3875
0 3877 7 4 2 44609 42489
0 3878 7 5 2 43649 55826
0 3879 7 3 2 55830 50805
0 3880 7 6 2 42049 47383
0 3881 5 2 1 55838
0 3882 7 1 2 45605 51113
0 3883 5 1 1 3882
0 3884 7 1 2 55839 3883
0 3885 5 1 1 3884
0 3886 7 1 2 41895 51190
0 3887 5 1 1 3886
0 3888 7 1 2 3885 3887
0 3889 5 1 1 3888
0 3890 7 1 2 55835 3889
0 3891 5 1 1 3890
0 3892 7 3 2 41438 53578
0 3893 5 1 1 55846
0 3894 7 3 2 47384 51030
0 3895 7 1 2 55847 55849
0 3896 5 1 1 3895
0 3897 7 1 2 54344 47705
0 3898 7 1 2 55710 3897
0 3899 5 1 1 3898
0 3900 7 1 2 3896 3899
0 3901 5 1 1 3900
0 3902 7 1 2 49407 3901
0 3903 5 1 1 3902
0 3904 7 8 2 45826 49408
0 3905 7 2 2 47706 55852
0 3906 7 1 2 55860 55711
0 3907 5 1 1 3906
0 3908 7 6 2 44478 45405
0 3909 5 3 1 55862
0 3910 7 1 2 43506 55863
0 3911 5 4 1 3910
0 3912 7 1 2 50304 49959
0 3913 5 1 1 3912
0 3914 7 1 2 44610 3913
0 3915 5 1 1 3914
0 3916 7 1 2 55871 3915
0 3917 5 1 1 3916
0 3918 7 1 2 42267 3917
0 3919 5 1 1 3918
0 3920 7 2 2 45606 47385
0 3921 7 3 2 49873 55875
0 3922 5 3 1 55877
0 3923 7 1 2 42050 55878
0 3924 5 1 1 3923
0 3925 7 1 2 45827 3924
0 3926 7 1 2 3919 3925
0 3927 5 1 1 3926
0 3928 7 1 2 41190 50573
0 3929 5 1 1 3928
0 3930 7 1 2 41319 50466
0 3931 5 1 1 3930
0 3932 7 1 2 42490 3931
0 3933 7 1 2 3929 3932
0 3934 5 1 1 3933
0 3935 7 1 2 44743 3934
0 3936 7 1 2 3927 3935
0 3937 5 1 1 3936
0 3938 7 1 2 3907 3937
0 3939 5 1 1 3938
0 3940 7 1 2 43858 3939
0 3941 5 1 1 3940
0 3942 7 1 2 3903 3941
0 3943 5 1 1 3942
0 3944 7 1 2 42768 3943
0 3945 5 1 1 3944
0 3946 7 1 2 3891 3945
0 3947 5 1 1 3946
0 3948 7 1 2 41586 3947
0 3949 5 1 1 3948
0 3950 7 10 2 44611 41896
0 3951 5 3 1 55883
0 3952 7 2 2 43650 55884
0 3953 7 2 2 47707 55896
0 3954 7 1 2 55712 55898
0 3955 5 1 1 3954
0 3956 7 1 2 46829 50305
0 3957 5 1 1 3956
0 3958 7 1 2 42051 3957
0 3959 5 2 1 3958
0 3960 7 4 2 46965 55900
0 3961 5 1 1 55902
0 3962 7 2 2 50164 55903
0 3963 5 1 1 55906
0 3964 7 1 2 44612 3963
0 3965 5 1 1 3964
0 3966 7 2 2 45406 49874
0 3967 7 1 2 41897 55908
0 3968 5 1 1 3967
0 3969 7 2 2 3965 3968
0 3970 7 1 2 42268 55910
0 3971 5 1 1 3970
0 3972 7 1 2 49875 55840
0 3973 5 2 1 3972
0 3974 7 1 2 49470 55912
0 3975 5 1 1 3974
0 3976 7 1 2 41898 3975
0 3977 5 1 1 3976
0 3978 7 2 2 47708 54034
0 3979 5 1 1 55914
0 3980 7 1 2 45607 3979
0 3981 7 1 2 3977 3980
0 3982 5 1 1 3981
0 3983 7 1 2 49570 3982
0 3984 7 1 2 3971 3983
0 3985 5 1 1 3984
0 3986 7 1 2 3955 3985
0 3987 5 1 1 3986
0 3988 7 1 2 54379 3987
0 3989 5 1 1 3988
0 3990 7 4 2 41899 49876
0 3991 5 2 1 55916
0 3992 7 2 2 40344 47454
0 3993 5 2 1 55922
0 3994 7 1 2 49877 55924
0 3995 7 3 2 51819 3994
0 3996 5 1 1 55926
0 3997 7 3 2 55920 3996
0 3998 7 1 2 42269 55929
0 3999 5 1 1 3998
0 4000 7 1 2 51958 52795
0 4001 5 2 1 4000
0 4002 7 1 2 3999 55932
0 4003 5 1 1 4002
0 4004 7 1 2 41320 4003
0 4005 5 1 1 4004
0 4006 7 2 2 41321 47872
0 4007 5 1 1 55934
0 4008 7 2 2 42270 50178
0 4009 5 1 1 55936
0 4010 7 1 2 55487 55937
0 4011 5 1 1 4010
0 4012 7 1 2 4007 4011
0 4013 5 1 1 4012
0 4014 7 1 2 45407 4013
0 4015 5 1 1 4014
0 4016 7 1 2 4005 4015
0 4017 5 1 1 4016
0 4018 7 1 2 49571 4017
0 4019 5 1 1 4018
0 4020 7 1 2 45408 50319
0 4021 7 1 2 49739 4020
0 4022 5 1 1 4021
0 4023 7 4 2 41439 47386
0 4024 7 3 2 49409 55938
0 4025 7 2 2 40566 42271
0 4026 5 3 1 55945
0 4027 7 1 2 47709 54775
0 4028 5 2 1 4027
0 4029 7 1 2 55947 55950
0 4030 5 1 1 4029
0 4031 7 1 2 55942 4030
0 4032 5 1 1 4031
0 4033 7 1 2 47516 51757
0 4034 5 1 1 4033
0 4035 7 1 2 49934 4034
0 4036 5 1 1 4035
0 4037 7 1 2 43859 54995
0 4038 7 1 2 4036 4037
0 4039 5 1 1 4038
0 4040 7 1 2 4032 4039
0 4041 5 1 1 4040
0 4042 7 1 2 42052 4041
0 4043 5 1 1 4042
0 4044 7 1 2 4022 4043
0 4045 7 1 2 4019 4044
0 4046 5 1 1 4045
0 4047 7 1 2 42491 4046
0 4048 5 1 1 4047
0 4049 7 1 2 46044 4048
0 4050 7 1 2 3989 4049
0 4051 5 1 1 4050
0 4052 7 1 2 55735 50567
0 4053 5 1 1 4052
0 4054 7 2 2 40167 55748
0 4055 5 1 1 55952
0 4056 7 1 2 55746 55659
0 4057 5 1 1 4056
0 4058 7 1 2 47455 4057
0 4059 5 1 1 4058
0 4060 7 1 2 55663 4059
0 4061 7 1 2 4055 4060
0 4062 5 1 1 4061
0 4063 7 1 2 45409 4062
0 4064 5 1 1 4063
0 4065 7 1 2 4053 4064
0 4066 5 1 1 4065
0 4067 7 1 2 45608 4066
0 4068 5 1 1 4067
0 4069 7 3 2 39955 52318
0 4070 5 2 1 55954
0 4071 7 2 2 51739 55955
0 4072 7 1 2 55736 55959
0 4073 5 1 1 4072
0 4074 7 1 2 4068 4073
0 4075 5 1 1 4074
0 4076 7 1 2 41191 4075
0 4077 5 1 1 4076
0 4078 7 4 2 49634 46787
0 4079 7 2 2 45609 55961
0 4080 7 1 2 39956 51946
0 4081 7 1 2 55965 4080
0 4082 5 1 1 4081
0 4083 7 1 2 4077 4082
0 4084 5 1 1 4083
0 4085 7 1 2 48653 4084
0 4086 5 1 1 4085
0 4087 7 1 2 42769 4086
0 4088 5 1 1 4087
0 4089 7 1 2 44891 4088
0 4090 7 1 2 4051 4089
0 4091 5 1 1 4090
0 4092 7 1 2 3949 4091
0 4093 5 1 1 4092
0 4094 7 1 2 44009 4093
0 4095 5 1 1 4094
0 4096 7 1 2 3876 4095
0 4097 5 1 1 4096
0 4098 7 1 2 46206 4097
0 4099 5 1 1 4098
0 4100 7 2 2 43315 50336
0 4101 7 1 2 55698 55967
0 4102 7 1 2 54055 4101
0 4103 5 1 1 4102
0 4104 7 1 2 54062 4103
0 4105 5 1 1 4104
0 4106 7 2 2 55786 50129
0 4107 7 1 2 48097 55969
0 4108 7 1 2 54399 4107
0 4109 7 1 2 4105 4108
0 4110 5 1 1 4109
0 4111 7 1 2 4099 4110
0 4112 5 1 1 4111
0 4113 7 1 2 41718 4112
0 4114 5 1 1 4113
0 4115 7 1 2 3843 4114
0 4116 5 1 1 4115
0 4117 7 1 2 40911 4116
0 4118 5 1 1 4117
0 4119 7 1 2 44479 50578
0 4120 5 3 1 4119
0 4121 7 2 2 55971 53676
0 4122 5 1 1 55974
0 4123 7 1 2 43507 4122
0 4124 5 1 1 4123
0 4125 7 3 2 43651 48003
0 4126 5 1 1 55976
0 4127 7 1 2 45610 55977
0 4128 5 1 1 4127
0 4129 7 1 2 4124 4128
0 4130 5 1 1 4129
0 4131 7 1 2 45828 4130
0 4132 5 1 1 4131
0 4133 7 1 2 52474 4132
0 4134 5 1 1 4133
0 4135 7 1 2 44892 4134
0 4136 5 1 1 4135
0 4137 7 3 2 50320 54422
0 4138 7 5 2 41587 49410
0 4139 5 1 1 55982
0 4140 7 1 2 55979 55983
0 4141 5 1 1 4140
0 4142 7 1 2 4136 4141
0 4143 5 1 1 4142
0 4144 7 1 2 46045 4143
0 4145 5 1 1 4144
0 4146 7 1 2 50604 48182
0 4147 5 6 1 4146
0 4148 7 2 2 43508 55987
0 4149 5 2 1 55993
0 4150 7 1 2 55995 55975
0 4151 5 1 1 4150
0 4152 7 9 2 41588 45829
0 4153 5 1 1 55997
0 4154 7 1 2 47847 55998
0 4155 7 1 2 4151 4154
0 4156 5 1 1 4155
0 4157 7 1 2 4145 4156
0 4158 5 1 1 4157
0 4159 7 1 2 40567 4158
0 4160 5 1 1 4159
0 4161 7 11 2 42272 53806
0 4162 5 1 1 56006
0 4163 7 2 2 50979 55439
0 4164 7 1 2 56007 56017
0 4165 5 1 1 4164
0 4166 7 1 2 4160 4165
0 4167 5 1 1 4166
0 4168 7 1 2 41440 4167
0 4169 5 1 1 4168
0 4170 7 1 2 55405 54943
0 4171 7 1 2 56018 4170
0 4172 5 1 1 4171
0 4173 7 1 2 4169 4172
0 4174 5 1 1 4173
0 4175 7 1 2 48993 4174
0 4176 5 1 1 4175
0 4177 7 1 2 44893 55988
0 4178 7 1 2 54400 4177
0 4179 5 1 1 4178
0 4180 7 1 2 54266 51005
0 4181 7 1 2 51198 4180
0 4182 5 1 1 4181
0 4183 7 1 2 4179 4182
0 4184 5 1 1 4183
0 4185 7 1 2 43509 4184
0 4186 5 1 1 4185
0 4187 7 3 2 44744 51972
0 4188 5 2 1 56019
0 4189 7 1 2 45410 51721
0 4190 5 1 1 4189
0 4191 7 1 2 56022 4190
0 4192 5 1 1 4191
0 4193 7 1 2 43860 4192
0 4194 5 1 1 4193
0 4195 7 1 2 54345 51653
0 4196 5 1 1 4195
0 4197 7 1 2 4194 4196
0 4198 5 1 1 4197
0 4199 7 1 2 44480 4198
0 4200 5 1 1 4199
0 4201 7 11 2 40568 54308
0 4202 5 1 1 56024
0 4203 7 1 2 55602 56025
0 4204 5 1 1 4203
0 4205 7 1 2 4200 4204
0 4206 5 1 1 4205
0 4207 7 1 2 42273 4206
0 4208 5 1 1 4207
0 4209 7 1 2 4186 4208
0 4210 5 1 1 4209
0 4211 7 1 2 47848 4210
0 4212 5 1 1 4211
0 4213 7 6 2 43510 42492
0 4214 7 5 2 43861 44481
0 4215 7 6 2 44745 56041
0 4216 5 1 1 56046
0 4217 7 1 2 56035 56047
0 4218 7 1 2 52739 4217
0 4219 5 1 1 4218
0 4220 7 1 2 4212 4219
0 4221 5 1 1 4220
0 4222 7 4 2 43652 40912
0 4223 7 2 2 44613 41719
0 4224 7 1 2 56052 56056
0 4225 7 1 2 4221 4224
0 4226 5 1 1 4225
0 4227 7 1 2 4176 4226
0 4228 5 1 1 4227
0 4229 7 1 2 40738 4228
0 4230 5 1 1 4229
0 4231 7 6 2 41720 55167
0 4232 7 17 2 45611 42770
0 4233 7 4 2 41589 50690
0 4234 7 1 2 56064 56081
0 4235 5 2 1 4234
0 4236 7 1 2 45411 52740
0 4237 5 1 1 4236
0 4238 7 1 2 56085 4237
0 4239 5 1 1 4238
0 4240 7 1 2 47710 4239
0 4241 5 1 1 4240
0 4242 7 11 2 42274 42771
0 4243 7 4 2 41590 50871
0 4244 7 1 2 56087 56098
0 4245 5 1 1 4244
0 4246 7 1 2 4241 4245
0 4247 5 1 1 4246
0 4248 7 2 2 47620 4247
0 4249 7 1 2 54309 49411
0 4250 5 1 1 4249
0 4251 7 1 2 41441 49471
0 4252 5 2 1 4251
0 4253 7 2 2 54711 56104
0 4254 5 2 1 56106
0 4255 7 2 2 48543 56107
0 4256 7 1 2 45830 56110
0 4257 5 1 1 4256
0 4258 7 1 2 4250 4257
0 4259 5 1 1 4258
0 4260 7 1 2 56102 4259
0 4261 5 1 1 4260
0 4262 7 2 2 54527 55715
0 4263 5 1 1 56112
0 4264 7 8 2 45831 48154
0 4265 7 1 2 44894 56114
0 4266 5 1 1 4265
0 4267 7 1 2 4263 4266
0 4268 5 1 1 4267
0 4269 7 1 2 43511 4268
0 4270 5 1 1 4269
0 4271 7 1 2 41591 55980
0 4272 5 1 1 4271
0 4273 7 1 2 55532 4272
0 4274 5 1 1 4273
0 4275 7 1 2 44614 4274
0 4276 5 1 1 4275
0 4277 7 1 2 48181 51722
0 4278 5 1 1 4277
0 4279 7 1 2 4276 4278
0 4280 7 1 2 4270 4279
0 4281 5 1 1 4280
0 4282 7 1 2 46046 4281
0 4283 5 1 1 4282
0 4284 7 1 2 55510 56082
0 4285 5 1 1 4284
0 4286 7 1 2 4283 4285
0 4287 5 1 1 4286
0 4288 7 1 2 43653 4287
0 4289 5 1 1 4288
0 4290 7 1 2 52469 46664
0 4291 5 1 1 4290
0 4292 7 1 2 4289 4291
0 4293 5 1 1 4292
0 4294 7 1 2 49572 4293
0 4295 5 1 1 4294
0 4296 7 1 2 4261 4295
0 4297 5 1 1 4296
0 4298 7 1 2 56058 4297
0 4299 5 1 1 4298
0 4300 7 1 2 4230 4299
0 4301 5 1 1 4300
0 4302 7 1 2 46207 4301
0 4303 5 1 1 4302
0 4304 7 1 2 55972 55996
0 4305 5 3 1 4304
0 4306 7 1 2 56122 54401
0 4307 5 1 1 4306
0 4308 7 1 2 51031 56026
0 4309 5 1 1 4308
0 4310 7 1 2 4307 4309
0 4311 5 1 1 4310
0 4312 7 5 2 40913 52226
0 4313 7 2 2 56125 55791
0 4314 7 1 2 42929 53135
0 4315 7 1 2 56130 4314
0 4316 7 1 2 4311 4315
0 4317 5 1 1 4316
0 4318 7 1 2 4303 4317
0 4319 5 1 1 4318
0 4320 7 1 2 47316 4319
0 4321 5 1 1 4320
0 4322 7 4 2 44164 46208
0 4323 7 6 2 40569 44615
0 4324 7 2 2 56136 51216
0 4325 7 2 2 51911 50069
0 4326 7 1 2 56142 56144
0 4327 5 1 1 4326
0 4328 7 8 2 45832 51994
0 4329 7 2 2 50070 50730
0 4330 5 1 1 56154
0 4331 7 2 2 41592 51297
0 4332 5 1 1 56156
0 4333 7 1 2 53050 4332
0 4334 5 4 1 4333
0 4335 7 2 2 41442 56158
0 4336 7 1 2 40570 56162
0 4337 5 1 1 4336
0 4338 7 1 2 4330 4337
0 4339 5 1 1 4338
0 4340 7 1 2 56146 4339
0 4341 5 1 1 4340
0 4342 7 7 2 41721 42493
0 4343 7 1 2 48334 56164
0 4344 7 1 2 52139 4343
0 4345 5 1 1 4344
0 4346 7 1 2 4341 4345
0 4347 5 1 1 4346
0 4348 7 1 2 52978 4347
0 4349 5 1 1 4348
0 4350 7 1 2 4327 4349
0 4351 5 1 1 4350
0 4352 7 1 2 55488 4351
0 4353 5 1 1 4352
0 4354 7 2 2 47456 47965
0 4355 5 1 1 56171
0 4356 7 1 2 50199 56172
0 4357 5 1 1 4356
0 4358 7 1 2 50172 4357
0 4359 5 1 1 4358
0 4360 7 1 2 46665 4359
0 4361 5 1 1 4360
0 4362 7 1 2 47218 50467
0 4363 5 1 1 4362
0 4364 7 1 2 4361 4363
0 4365 5 1 1 4364
0 4366 7 1 2 41322 4365
0 4367 5 1 1 4366
0 4368 7 13 2 45246 45612
0 4369 5 4 1 56173
0 4370 7 3 2 42772 56174
0 4371 7 1 2 50557 50769
0 4372 7 1 2 56190 4371
0 4373 5 1 1 4372
0 4374 7 1 2 4367 4373
0 4375 5 1 1 4374
0 4376 7 1 2 42494 4375
0 4377 5 1 1 4376
0 4378 7 1 2 50321 47266
0 4379 5 1 1 4378
0 4380 7 1 2 43654 51058
0 4381 7 1 2 56186 4380
0 4382 5 1 1 4381
0 4383 7 1 2 4379 4382
0 4384 5 1 1 4383
0 4385 7 1 2 46666 4384
0 4386 5 1 1 4385
0 4387 7 1 2 47219 47842
0 4388 5 1 1 4387
0 4389 7 1 2 4386 4388
0 4390 5 1 1 4389
0 4391 7 1 2 55451 4390
0 4392 5 1 1 4391
0 4393 7 1 2 55546 4392
0 4394 7 1 2 4377 4393
0 4395 5 1 1 4394
0 4396 7 1 2 41443 4395
0 4397 5 1 1 4396
0 4398 7 1 2 55584 4397
0 4399 5 1 1 4398
0 4400 7 1 2 40571 4399
0 4401 5 1 1 4400
0 4402 7 1 2 48463 55624
0 4403 5 1 1 4402
0 4404 7 1 2 55610 4403
0 4405 5 1 1 4404
0 4406 7 1 2 47766 4405
0 4407 5 1 1 4406
0 4408 7 6 2 45412 47457
0 4409 5 12 1 56193
0 4410 7 1 2 56199 53152
0 4411 5 1 1 4410
0 4412 7 1 2 55652 4411
0 4413 5 1 1 4412
0 4414 7 1 2 54346 55641
0 4415 5 1 1 4414
0 4416 7 4 2 44746 53229
0 4417 5 1 1 56211
0 4418 7 1 2 55761 56212
0 4419 5 1 1 4418
0 4420 7 1 2 4415 4419
0 4421 5 1 1 4420
0 4422 7 1 2 46667 4421
0 4423 5 1 1 4422
0 4424 7 1 2 4413 4423
0 4425 5 1 1 4424
0 4426 7 1 2 45613 4425
0 4427 5 1 1 4426
0 4428 7 1 2 55694 4427
0 4429 5 1 1 4428
0 4430 7 1 2 52584 4429
0 4431 5 1 1 4430
0 4432 7 1 2 55733 4431
0 4433 7 1 2 4407 4432
0 4434 7 1 2 4401 4433
0 4435 5 1 1 4434
0 4436 7 1 2 41722 4435
0 4437 5 1 1 4436
0 4438 7 1 2 4353 4437
0 4439 5 1 1 4438
0 4440 7 1 2 40739 4439
0 4441 5 1 1 4440
0 4442 7 1 2 41723 55784
0 4443 5 1 1 4442
0 4444 7 1 2 4441 4443
0 4445 5 1 1 4444
0 4446 7 1 2 56132 4445
0 4447 5 1 1 4446
0 4448 7 2 2 42275 52807
0 4449 7 1 2 44616 56215
0 4450 5 1 1 4449
0 4451 7 1 2 53738 4450
0 4452 5 1 1 4451
0 4453 7 1 2 45833 4452
0 4454 5 1 1 4453
0 4455 7 1 2 53789 4454
0 4456 5 1 1 4455
0 4457 7 1 2 51641 4456
0 4458 5 1 1 4457
0 4459 7 7 2 46209 48956
0 4460 5 1 1 56217
0 4461 7 1 2 47840 4355
0 4462 5 1 1 4461
0 4463 7 1 2 44617 4462
0 4464 5 1 1 4463
0 4465 7 1 2 42276 54210
0 4466 5 1 1 4465
0 4467 7 1 2 174 4466
0 4468 5 1 1 4467
0 4469 7 1 2 47909 4468
0 4470 5 1 1 4469
0 4471 7 1 2 47873 53174
0 4472 5 1 1 4471
0 4473 7 1 2 54063 4472
0 4474 7 1 2 4470 4473
0 4475 7 1 2 4464 4474
0 4476 5 1 1 4475
0 4477 7 1 2 45834 4476
0 4478 5 1 1 4477
0 4479 7 1 2 53754 52519
0 4480 5 1 1 4479
0 4481 7 1 2 41192 4480
0 4482 5 1 1 4481
0 4483 7 1 2 53790 4482
0 4484 7 1 2 4478 4483
0 4485 5 1 1 4484
0 4486 7 1 2 56218 4485
0 4487 5 1 1 4486
0 4488 7 1 2 4458 4487
0 4489 5 1 1 4488
0 4490 7 1 2 53863 4489
0 4491 5 1 1 4490
0 4492 7 5 2 40914 49851
0 4493 7 1 2 56224 56191
0 4494 5 1 1 4493
0 4495 7 4 2 40345 41593
0 4496 7 1 2 46047 50579
0 4497 7 1 2 56229 4496
0 4498 7 1 2 48994 4497
0 4499 5 1 1 4498
0 4500 7 1 2 4494 4499
0 4501 5 1 1 4500
0 4502 7 1 2 54253 4501
0 4503 5 1 1 4502
0 4504 7 1 2 40915 51430
0 4505 7 1 2 56145 4504
0 4506 5 1 1 4505
0 4507 7 1 2 4503 4506
0 4508 5 1 1 4507
0 4509 7 1 2 50558 4508
0 4510 5 1 1 4509
0 4511 7 6 2 49305 49292
0 4512 5 3 1 56233
0 4513 7 1 2 45413 56239
0 4514 5 3 1 4513
0 4515 7 1 2 56242 55904
0 4516 5 1 1 4515
0 4517 7 1 2 42277 4516
0 4518 5 2 1 4517
0 4519 7 1 2 56245 46938
0 4520 5 1 1 4519
0 4521 7 1 2 44618 4520
0 4522 5 1 1 4521
0 4523 7 1 2 51059 52729
0 4524 7 1 2 46932 4523
0 4525 5 1 1 4524
0 4526 7 1 2 50605 234
0 4527 5 3 1 4526
0 4528 7 2 2 56247 51864
0 4529 5 1 1 56250
0 4530 7 1 2 46869 56251
0 4531 5 1 1 4530
0 4532 7 13 2 43316 46707
0 4533 5 2 1 56252
0 4534 7 5 2 44482 45614
0 4535 5 1 1 56267
0 4536 7 1 2 56253 56268
0 4537 5 1 1 4536
0 4538 7 1 2 50610 4537
0 4539 5 1 1 4538
0 4540 7 1 2 43655 4539
0 4541 5 1 1 4540
0 4542 7 1 2 45835 4541
0 4543 7 1 2 4531 4542
0 4544 7 1 2 4525 4543
0 4545 7 1 2 4522 4544
0 4546 5 1 1 4545
0 4547 7 2 2 48995 49077
0 4548 7 3 2 50677 48172
0 4549 5 20 1 56274
0 4550 7 1 2 56277 55930
0 4551 5 1 1 4550
0 4552 7 1 2 42053 50310
0 4553 5 2 1 4552
0 4554 7 2 2 41900 47267
0 4555 5 2 1 56299
0 4556 7 1 2 56297 56301
0 4557 7 1 2 56243 4556
0 4558 5 1 1 4557
0 4559 7 1 2 51995 4558
0 4560 5 1 1 4559
0 4561 7 4 2 41323 48155
0 4562 5 2 1 56303
0 4563 7 1 2 42278 51673
0 4564 5 1 1 4563
0 4565 7 1 2 56307 4564
0 4566 5 1 1 4565
0 4567 7 1 2 47517 4566
0 4568 5 1 1 4567
0 4569 7 1 2 42495 4568
0 4570 7 1 2 4560 4569
0 4571 7 1 2 4551 4570
0 4572 5 1 1 4571
0 4573 7 1 2 56272 4572
0 4574 7 1 2 4546 4573
0 4575 5 1 1 4574
0 4576 7 1 2 4510 4575
0 4577 5 1 1 4576
0 4578 7 1 2 46210 4577
0 4579 5 1 1 4578
0 4580 7 1 2 4491 4579
0 4581 5 1 1 4580
0 4582 7 1 2 53527 4581
0 4583 5 1 1 4582
0 4584 7 1 2 47767 55703
0 4585 5 4 1 4584
0 4586 7 1 2 44619 56309
0 4587 5 1 1 4586
0 4588 7 1 2 47571 4587
0 4589 7 1 2 51586 47910
0 4590 5 2 1 4589
0 4591 7 1 2 47911 51789
0 4592 5 1 1 4591
0 4593 7 1 2 56313 4592
0 4594 7 1 2 4588 4593
0 4595 5 1 1 4594
0 4596 7 1 2 45615 4595
0 4597 5 1 1 4596
0 4598 7 1 2 43317 54769
0 4599 5 1 1 4598
0 4600 7 2 2 4599 3211
0 4601 5 1 1 56315
0 4602 7 1 2 42279 4601
0 4603 5 2 1 4602
0 4604 7 2 2 48810 52681
0 4605 5 3 1 56319
0 4606 7 1 2 56317 56321
0 4607 7 1 2 4597 4606
0 4608 5 1 1 4607
0 4609 7 3 2 40740 53864
0 4610 7 1 2 42930 56324
0 4611 7 1 2 4608 4610
0 4612 5 1 1 4611
0 4613 7 7 2 45616 46211
0 4614 7 1 2 56327 48996
0 4615 7 1 2 55489 4614
0 4616 7 1 2 51678 4615
0 4617 5 1 1 4616
0 4618 7 1 2 4612 4617
0 4619 5 1 1 4618
0 4620 7 1 2 45836 4619
0 4621 5 1 1 4620
0 4622 7 6 2 40346 40741
0 4623 7 3 2 41324 56334
0 4624 7 1 2 51286 56340
0 4625 5 1 1 4624
0 4626 7 16 2 44010 46212
0 4627 7 1 2 41901 53857
0 4628 5 1 1 4627
0 4629 7 1 2 51758 4628
0 4630 5 1 1 4629
0 4631 7 4 2 51032 4630
0 4632 7 1 2 56343 56359
0 4633 5 1 1 4632
0 4634 7 1 2 4625 4633
0 4635 5 1 1 4634
0 4636 7 2 2 40916 42496
0 4637 7 1 2 41724 56363
0 4638 7 1 2 4635 4637
0 4639 5 1 1 4638
0 4640 7 1 2 4621 4639
0 4641 5 1 1 4640
0 4642 7 1 2 48464 4641
0 4643 5 1 1 4642
0 4644 7 2 2 51759 696
0 4645 5 1 1 56365
0 4646 7 5 2 43862 40917
0 4647 7 1 2 56367 52855
0 4648 7 1 2 53511 4647
0 4649 7 1 2 54538 4648
0 4650 7 1 2 4645 4649
0 4651 5 1 1 4650
0 4652 7 1 2 4643 4651
0 4653 5 1 1 4652
0 4654 7 1 2 52900 4653
0 4655 5 1 1 4654
0 4656 7 1 2 4583 4655
0 4657 7 1 2 4447 4656
0 4658 7 3 2 46213 53357
0 4659 7 1 2 54916 56372
0 4660 5 1 1 4659
0 4661 7 1 2 50909 48149
0 4662 7 1 2 51719 4661
0 4663 5 1 1 4662
0 4664 7 1 2 4660 4663
0 4665 5 1 1 4664
0 4666 7 1 2 43318 4665
0 4667 5 1 1 4666
0 4668 7 2 2 49977 53242
0 4669 7 1 2 48465 46830
0 4670 7 1 2 56375 4669
0 4671 5 1 1 4670
0 4672 7 1 2 4667 4671
0 4673 5 1 1 4672
0 4674 7 1 2 40918 4673
0 4675 5 1 1 4674
0 4676 7 9 2 40572 45617
0 4677 7 2 2 44165 52856
0 4678 5 1 1 56386
0 4679 7 1 2 56377 56387
0 4680 7 1 2 50405 4679
0 4681 5 1 1 4680
0 4682 7 1 2 4675 4681
0 4683 5 1 1 4682
0 4684 7 1 2 44483 4683
0 4685 5 1 1 4684
0 4686 7 5 2 45618 50842
0 4687 5 3 1 56388
0 4688 7 2 2 51060 56393
0 4689 7 1 2 48997 56373
0 4690 7 1 2 56396 4689
0 4691 5 1 1 4690
0 4692 7 1 2 4685 4691
0 4693 5 1 1 4692
0 4694 7 1 2 46048 4693
0 4695 5 1 1 4694
0 4696 7 1 2 47891 46773
0 4697 5 1 1 4696
0 4698 7 1 2 46214 48466
0 4699 7 2 2 48998 4698
0 4700 7 6 2 41594 56065
0 4701 5 3 1 56400
0 4702 7 1 2 56398 56401
0 4703 7 1 2 4697 4702
0 4704 5 1 1 4703
0 4705 7 1 2 4695 4704
0 4706 5 1 1 4705
0 4707 7 1 2 43512 4706
0 4708 5 1 1 4707
0 4709 7 1 2 46668 56397
0 4710 5 2 1 4709
0 4711 7 1 2 47912 56402
0 4712 5 1 1 4711
0 4713 7 1 2 56409 4712
0 4714 5 1 1 4713
0 4715 7 1 2 44484 4714
0 4716 5 1 1 4715
0 4717 7 4 2 46049 47317
0 4718 7 2 2 42280 51654
0 4719 7 1 2 56411 56415
0 4720 5 1 1 4719
0 4721 7 1 2 4716 4720
0 4722 5 2 1 4721
0 4723 7 1 2 56399 56417
0 4724 5 1 1 4723
0 4725 7 1 2 4708 4724
0 4726 5 1 1 4725
0 4727 7 1 2 40742 4726
0 4728 5 1 1 4727
0 4729 7 2 2 50631 56059
0 4730 7 1 2 47833 56403
0 4731 5 1 1 4730
0 4732 7 1 2 56410 4731
0 4733 5 1 1 4732
0 4734 7 1 2 47621 4733
0 4735 5 1 1 4734
0 4736 7 2 2 51061 54056
0 4737 7 1 2 47318 56421
0 4738 5 1 1 4737
0 4739 7 1 2 55951 4738
0 4740 5 1 1 4739
0 4741 7 1 2 46669 4740
0 4742 5 1 1 4741
0 4743 7 1 2 4735 4742
0 4744 5 1 1 4743
0 4745 7 1 2 56419 4744
0 4746 5 1 1 4745
0 4747 7 1 2 4728 4746
0 4748 5 1 1 4747
0 4749 7 1 2 45837 4748
0 4750 5 1 1 4749
0 4751 7 1 2 46050 46831
0 4752 7 1 2 51480 4751
0 4753 5 1 1 4752
0 4754 7 1 2 51414 48311
0 4755 7 1 2 50071 4754
0 4756 5 1 1 4755
0 4757 7 1 2 4753 4756
0 4758 5 1 1 4757
0 4759 7 1 2 41595 4758
0 4760 5 1 1 4759
0 4761 7 1 2 50104 48352
0 4762 5 1 1 4761
0 4763 7 1 2 216 334
0 4764 5 1 1 4763
0 4765 7 4 2 44011 42773
0 4766 5 1 1 56423
0 4767 7 1 2 40573 4766
0 4768 7 1 2 4764 4767
0 4769 5 1 1 4768
0 4770 7 1 2 4762 4769
0 4771 5 1 1 4770
0 4772 7 2 2 44895 4771
0 4773 5 1 1 56427
0 4774 7 1 2 54879 56428
0 4775 5 1 1 4774
0 4776 7 1 2 4760 4775
0 4777 5 1 1 4776
0 4778 7 1 2 43319 4777
0 4779 5 1 1 4778
0 4780 7 6 2 41725 46051
0 4781 7 1 2 56429 51501
0 4782 5 1 1 4781
0 4783 7 1 2 51452 56163
0 4784 5 1 1 4783
0 4785 7 1 2 4782 4784
0 4786 5 1 1 4785
0 4787 7 1 2 46708 4786
0 4788 5 1 1 4787
0 4789 7 1 2 4779 4788
0 4790 5 1 1 4789
0 4791 7 1 2 40919 4790
0 4792 5 1 1 4791
0 4793 7 1 2 49126 52599
0 4794 7 1 2 47913 4793
0 4795 5 1 1 4794
0 4796 7 1 2 4792 4795
0 4797 5 1 1 4796
0 4798 7 1 2 46215 4797
0 4799 5 1 1 4798
0 4800 7 4 2 48398 50941
0 4801 7 1 2 56435 56325
0 4802 7 1 2 51016 4801
0 4803 5 1 1 4802
0 4804 7 1 2 4799 4803
0 4805 5 1 1 4804
0 4806 7 1 2 47711 54539
0 4807 7 1 2 4805 4806
0 4808 5 1 1 4807
0 4809 7 1 2 4750 4808
0 4810 5 1 1 4809
0 4811 7 1 2 48728 4810
0 4812 5 1 1 4811
0 4813 7 8 2 40920 44747
0 4814 7 5 2 43863 56439
0 4815 7 2 2 49078 51445
0 4816 7 1 2 56447 56452
0 4817 5 1 1 4816
0 4818 7 1 2 40921 56159
0 4819 5 1 1 4818
0 4820 7 5 2 44166 41596
0 4821 5 1 1 56454
0 4822 7 3 2 41726 56455
0 4823 7 1 2 46052 56459
0 4824 5 1 1 4823
0 4825 7 1 2 4819 4824
0 4826 5 2 1 4825
0 4827 7 1 2 51465 56462
0 4828 5 1 1 4827
0 4829 7 1 2 4817 4828
0 4830 5 1 1 4829
0 4831 7 1 2 54423 4830
0 4832 5 1 1 4831
0 4833 7 1 2 4417 3893
0 4834 5 1 1 4833
0 4835 7 1 2 42774 4834
0 4836 5 1 1 4835
0 4837 7 4 2 45414 55224
0 4838 5 2 1 56464
0 4839 7 2 2 53807 53086
0 4840 5 1 1 56470
0 4841 7 1 2 56468 4840
0 4842 5 1 1 4841
0 4843 7 1 2 43864 4842
0 4844 5 1 1 4843
0 4845 7 1 2 4836 4844
0 4846 5 1 1 4845
0 4847 7 1 2 49180 4846
0 4848 5 1 1 4847
0 4849 7 3 2 44012 55568
0 4850 7 1 2 56472 55647
0 4851 5 1 1 4850
0 4852 7 1 2 47220 54291
0 4853 5 1 1 4852
0 4854 7 1 2 4851 4853
0 4855 5 1 1 4854
0 4856 7 1 2 43865 4855
0 4857 5 1 1 4856
0 4858 7 5 2 46053 54347
0 4859 5 1 1 56475
0 4860 7 1 2 50872 51514
0 4861 7 1 2 56476 4860
0 4862 5 1 1 4861
0 4863 7 1 2 4857 4862
0 4864 7 1 2 4848 4863
0 4865 5 1 1 4864
0 4866 7 1 2 53865 4865
0 4867 5 1 1 4866
0 4868 7 1 2 45415 53136
0 4869 7 1 2 54402 4868
0 4870 7 1 2 55163 4869
0 4871 5 1 1 4870
0 4872 7 1 2 4867 4871
0 4873 5 1 1 4872
0 4874 7 1 2 47387 4873
0 4875 5 1 1 4874
0 4876 7 1 2 4832 4875
0 4877 5 1 1 4876
0 4878 7 1 2 42281 4877
0 4879 5 1 1 4878
0 4880 7 5 2 43866 48601
0 4881 7 5 2 53866 56480
0 4882 5 1 1 56485
0 4883 7 1 2 48999 51466
0 4884 5 1 1 4883
0 4885 7 1 2 4882 4884
0 4886 5 4 1 4885
0 4887 7 2 2 50757 51723
0 4888 7 1 2 56490 56494
0 4889 5 1 1 4888
0 4890 7 1 2 4879 4889
0 4891 5 1 1 4890
0 4892 7 1 2 44620 4891
0 4893 5 1 1 4892
0 4894 7 1 2 47244 2386
0 4895 5 5 1 4894
0 4896 7 1 2 56115 56496
0 4897 7 1 2 56491 4896
0 4898 5 1 1 4897
0 4899 7 1 2 4893 4898
0 4900 5 1 1 4899
0 4901 7 1 2 43656 4900
0 4902 5 1 1 4901
0 4903 7 3 2 46054 51996
0 4904 7 1 2 52130 56501
0 4905 5 1 1 4904
0 4906 7 1 2 51912 47388
0 4907 7 1 2 56497 4906
0 4908 5 1 1 4907
0 4909 7 1 2 4905 4908
0 4910 5 1 1 4909
0 4911 7 1 2 45416 56492
0 4912 7 1 2 4910 4911
0 4913 5 1 1 4912
0 4914 7 1 2 4902 4913
0 4915 5 1 1 4914
0 4916 7 1 2 46216 4915
0 4917 5 1 1 4916
0 4918 7 1 2 54380 54699
0 4919 5 1 1 4918
0 4920 7 1 2 54332 4919
0 4921 5 1 1 4920
0 4922 7 1 2 50961 54721
0 4923 5 1 1 4922
0 4924 7 1 2 56131 48348
0 4925 7 1 2 4923 4924
0 4926 7 1 2 4921 4925
0 4927 5 1 1 4926
0 4928 7 1 2 4917 4927
0 4929 5 1 1 4928
0 4930 7 1 2 47622 4929
0 4931 5 1 1 4930
0 4932 7 1 2 4812 4931
0 4933 7 1 2 4657 4932
0 4934 7 1 2 4321 4933
0 4935 7 1 2 4118 4934
0 4936 5 1 1 4935
0 4937 7 1 2 46332 4936
0 4938 5 1 1 4937
0 4939 7 1 2 3529 4938
0 4940 5 1 1 4939
0 4941 7 1 2 55028 4940
0 4942 5 1 1 4941
0 4943 7 7 2 43867 53808
0 4944 5 2 1 56504
0 4945 7 2 2 56505 56278
0 4946 5 1 1 56513
0 4947 7 2 2 53809 53032
0 4948 5 1 1 56515
0 4949 7 1 2 55265 4948
0 4950 5 4 1 4949
0 4951 7 1 2 47002 56517
0 4952 5 1 1 4951
0 4953 7 1 2 4946 4952
0 4954 5 1 1 4953
0 4955 7 1 2 40347 4954
0 4956 5 1 1 4955
0 4957 7 1 2 55620 51086
0 4958 5 1 1 4957
0 4959 7 1 2 4956 4958
0 4960 5 1 1 4959
0 4961 7 1 2 44896 4960
0 4962 5 1 1 4961
0 4963 7 6 2 42282 49834
0 4964 5 1 1 56521
0 4965 7 4 2 42775 55999
0 4966 7 1 2 56522 56527
0 4967 5 1 1 4966
0 4968 7 1 2 4962 4967
0 4969 5 1 1 4968
0 4970 7 1 2 44748 4969
0 4971 5 1 1 4970
0 4972 7 3 2 40574 49728
0 4973 7 2 2 55225 52198
0 4974 7 1 2 56531 56534
0 4975 5 1 1 4974
0 4976 7 1 2 4971 4975
0 4977 5 1 1 4976
0 4978 7 1 2 44013 4977
0 4979 5 1 1 4978
0 4980 7 2 2 49573 51343
0 4981 7 1 2 56536 56535
0 4982 5 1 1 4981
0 4983 7 1 2 4979 4982
0 4984 5 1 1 4983
0 4985 7 1 2 54068 56133
0 4986 7 1 2 4984 4985
0 4987 5 1 1 4986
0 4988 7 11 2 41193 42283
0 4989 7 4 2 52172 56538
0 4990 5 2 1 56549
0 4991 7 6 2 43059 48573
0 4992 7 9 2 49369 52227
0 4993 7 1 2 56555 56561
0 4994 7 1 2 56550 4993
0 4995 7 1 2 56108 4994
0 4996 5 1 1 4995
0 4997 7 1 2 4987 4996
0 4998 5 1 1 4997
0 4999 7 1 2 46604 4998
0 5000 5 1 1 4999
0 5001 7 5 2 46333 52633
0 5002 7 3 2 53449 56570
0 5003 7 11 2 41597 45067
0 5004 7 1 2 56578 53487
0 5005 7 2 2 56575 5004
0 5006 7 7 2 44224 41194
0 5007 7 2 2 56591 53492
0 5008 7 2 2 55426 56335
0 5009 7 1 2 56598 56600
0 5010 7 1 2 56589 5009
0 5011 5 1 1 5010
0 5012 7 1 2 5000 5011
0 5013 5 1 1 5012
0 5014 7 1 2 52091 5013
0 5015 5 1 1 5014
0 5016 7 5 2 42284 48206
0 5017 7 8 2 39957 43868
0 5018 7 1 2 53204 56607
0 5019 7 1 2 51421 5018
0 5020 7 1 2 56602 5019
0 5021 5 1 1 5020
0 5022 7 1 2 48098 52204
0 5023 5 1 1 5022
0 5024 7 6 2 42776 49574
0 5025 7 1 2 56615 52875
0 5026 5 1 1 5025
0 5027 7 1 2 5023 5026
0 5028 5 1 1 5027
0 5029 7 1 2 54254 54567
0 5030 7 1 2 5028 5029
0 5031 5 1 1 5030
0 5032 7 1 2 5021 5031
0 5033 5 1 1 5032
0 5034 7 1 2 46334 5033
0 5035 5 1 1 5034
0 5036 7 11 2 42497 46335
0 5037 7 1 2 48099 52983
0 5038 5 1 1 5037
0 5039 7 1 2 52822 5038
0 5040 5 1 1 5039
0 5041 7 1 2 45016 5040
0 5042 5 1 1 5041
0 5043 7 1 2 1372 5042
0 5044 5 1 1 5043
0 5045 7 1 2 56621 5044
0 5046 5 1 1 5045
0 5047 7 7 2 45017 53623
0 5048 5 1 1 56632
0 5049 7 1 2 54639 5048
0 5050 5 2 1 5049
0 5051 7 1 2 51390 56639
0 5052 5 1 1 5051
0 5053 7 1 2 53605 52205
0 5054 5 1 1 5053
0 5055 7 1 2 5052 5054
0 5056 5 1 1 5055
0 5057 7 6 2 41195 45838
0 5058 5 1 1 56641
0 5059 7 1 2 56642 54568
0 5060 7 1 2 5056 5059
0 5061 5 1 1 5060
0 5062 7 1 2 5046 5061
0 5063 5 1 1 5062
0 5064 7 1 2 45619 5063
0 5065 5 1 1 5064
0 5066 7 2 2 53538 52984
0 5067 7 2 2 42285 55682
0 5068 5 3 1 56649
0 5069 7 1 2 56165 56651
0 5070 7 1 2 56647 5069
0 5071 5 1 1 5070
0 5072 7 1 2 5065 5071
0 5073 5 1 1 5072
0 5074 7 1 2 41325 5073
0 5075 5 1 1 5074
0 5076 7 1 2 5035 5075
0 5077 5 1 1 5076
0 5078 7 1 2 44167 5077
0 5079 5 1 1 5078
0 5080 7 11 2 42777 53624
0 5081 7 3 2 49575 56654
0 5082 5 1 1 56665
0 5083 7 1 2 56666 53794
0 5084 5 1 1 5083
0 5085 7 1 2 41326 56652
0 5086 7 1 2 56648 5085
0 5087 5 1 1 5086
0 5088 7 1 2 5084 5087
0 5089 5 1 1 5088
0 5090 7 1 2 42498 5089
0 5091 5 1 1 5090
0 5092 7 17 2 46055 43060
0 5093 7 7 2 45839 56668
0 5094 7 7 2 56685 56328
0 5095 5 1 1 56692
0 5096 7 2 2 47003 53420
0 5097 7 1 2 56693 56699
0 5098 5 1 1 5097
0 5099 7 1 2 5091 5098
0 5100 5 1 1 5099
0 5101 7 1 2 48981 5100
0 5102 5 1 1 5101
0 5103 7 1 2 5079 5102
0 5104 5 1 1 5103
0 5105 7 1 2 49181 5104
0 5106 5 1 1 5105
0 5107 7 10 2 41327 42499
0 5108 7 12 2 41444 45620
0 5109 5 2 1 56711
0 5110 7 2 2 40575 56712
0 5111 5 2 1 56725
0 5112 7 1 2 56701 56726
0 5113 5 1 1 5112
0 5114 7 1 2 53205 51997
0 5115 5 2 1 5114
0 5116 7 6 2 49635 54949
0 5117 7 3 2 42500 56731
0 5118 5 1 1 56737
0 5119 7 1 2 56729 5118
0 5120 5 3 1 5119
0 5121 7 1 2 51674 56740
0 5122 5 1 1 5121
0 5123 7 1 2 5113 5122
0 5124 5 1 1 5123
0 5125 7 1 2 49000 51515
0 5126 5 1 1 5125
0 5127 7 6 2 49102 50636
0 5128 5 1 1 56743
0 5129 7 1 2 5126 5128
0 5130 5 13 1 5129
0 5131 7 2 2 46336 56749
0 5132 7 1 2 5124 56762
0 5133 5 1 1 5132
0 5134 7 1 2 49636 52579
0 5135 5 1 1 5134
0 5136 7 1 2 56027 53103
0 5137 5 1 1 5136
0 5138 7 1 2 5135 5137
0 5139 5 1 1 5138
0 5140 7 6 2 39958 40743
0 5141 7 8 2 40922 41598
0 5142 7 3 2 54679 56770
0 5143 7 1 2 56764 56778
0 5144 7 1 2 5139 5143
0 5145 5 1 1 5144
0 5146 7 1 2 5133 5145
0 5147 5 1 1 5146
0 5148 7 1 2 42778 5147
0 5149 5 1 1 5148
0 5150 7 6 2 46056 46337
0 5151 7 1 2 55338 53795
0 5152 7 1 2 56750 5151
0 5153 5 1 1 5152
0 5154 7 4 2 44014 50394
0 5155 7 14 2 40348 40576
0 5156 5 2 1 56791
0 5157 7 1 2 45018 56792
0 5158 7 2 2 56787 5157
0 5159 7 3 2 44168 54843
0 5160 7 1 2 56809 53472
0 5161 7 1 2 56807 5160
0 5162 5 1 1 5161
0 5163 7 1 2 5153 5162
0 5164 5 1 1 5163
0 5165 7 1 2 56781 5164
0 5166 5 1 1 5165
0 5167 7 1 2 5149 5166
0 5168 5 1 1 5167
0 5169 7 1 2 42931 5168
0 5170 5 1 1 5169
0 5171 7 9 2 45621 43061
0 5172 7 3 2 56812 53488
0 5173 7 1 2 46057 56821
0 5174 7 1 2 54855 5173
0 5175 5 1 1 5174
0 5176 7 3 2 56137 53185
0 5177 5 1 1 56824
0 5178 7 1 2 5177 55012
0 5179 5 1 1 5178
0 5180 7 8 2 39959 46338
0 5181 7 1 2 56827 52758
0 5182 7 1 2 5179 5181
0 5183 5 1 1 5182
0 5184 7 1 2 5175 5183
0 5185 5 1 1 5184
0 5186 7 1 2 44169 5185
0 5187 5 1 1 5186
0 5188 7 2 2 45622 48982
0 5189 5 1 1 56835
0 5190 7 12 2 45417 43062
0 5191 7 1 2 56837 50942
0 5192 7 1 2 53440 5191
0 5193 7 1 2 56836 5192
0 5194 5 1 1 5193
0 5195 7 1 2 45840 5194
0 5196 7 1 2 5187 5195
0 5197 5 1 1 5196
0 5198 7 2 2 46058 52380
0 5199 5 1 1 56849
0 5200 7 2 2 56608 56850
0 5201 5 1 1 56851
0 5202 7 1 2 5201 53081
0 5203 5 1 1 5202
0 5204 7 1 2 52979 5203
0 5205 5 1 1 5204
0 5206 7 18 2 42779 48467
0 5207 5 3 1 56853
0 5208 7 1 2 51998 56854
0 5209 5 1 1 5208
0 5210 7 1 2 5205 5209
0 5211 5 1 1 5210
0 5212 7 1 2 54132 5211
0 5213 5 1 1 5212
0 5214 7 2 2 56669 55326
0 5215 7 2 2 56448 56874
0 5216 5 1 1 56876
0 5217 7 1 2 41328 56877
0 5218 5 1 1 5217
0 5219 7 1 2 42501 5218
0 5220 7 1 2 5213 5219
0 5221 5 1 1 5220
0 5222 7 1 2 51516 5221
0 5223 7 1 2 5197 5222
0 5224 5 1 1 5223
0 5225 7 1 2 49001 55339
0 5226 5 2 1 5225
0 5227 7 14 2 40349 44170
0 5228 7 1 2 53318 56880
0 5229 7 1 2 53309 5228
0 5230 5 1 1 5229
0 5231 7 1 2 56878 5230
0 5232 5 1 1 5231
0 5233 7 2 2 40744 41329
0 5234 5 1 1 56894
0 5235 7 1 2 56813 56895
0 5236 7 1 2 49079 5235
0 5237 7 1 2 5232 5236
0 5238 5 1 1 5237
0 5239 7 1 2 5224 5238
0 5240 5 1 1 5239
0 5241 7 1 2 46217 5240
0 5242 5 1 1 5241
0 5243 7 1 2 5170 5242
0 5244 7 1 2 5106 5243
0 5245 5 1 1 5244
0 5246 7 1 2 46605 5245
0 5247 5 1 1 5246
0 5248 7 6 2 39960 56793
0 5249 7 6 2 40923 44225
0 5250 7 5 2 40745 56902
0 5251 7 1 2 56896 56908
0 5252 7 1 2 53500 5251
0 5253 7 1 2 56590 5252
0 5254 5 1 1 5253
0 5255 7 1 2 5247 5254
0 5256 5 1 1 5255
0 5257 7 1 2 46732 5256
0 5258 5 1 1 5257
0 5259 7 1 2 5015 5258
0 5260 7 1 2 4942 5259
0 5261 7 1 2 3390 5260
0 5262 5 1 1 5261
0 5263 7 1 2 46445 5262
0 5264 5 1 1 5263
0 5265 7 7 2 42502 46446
0 5266 7 2 2 42932 56855
0 5267 7 1 2 56920 56230
0 5268 5 1 1 5267
0 5269 7 2 2 44749 48261
0 5270 5 1 1 56922
0 5271 7 2 2 43869 56923
0 5272 5 2 1 56924
0 5273 7 2 2 49711 56925
0 5274 5 1 1 56928
0 5275 7 1 2 40168 56929
0 5276 5 1 1 5275
0 5277 7 1 2 5268 5276
0 5278 5 1 1 5277
0 5279 7 1 2 40746 5278
0 5280 5 1 1 5279
0 5281 7 3 2 48207 51502
0 5282 5 2 1 56930
0 5283 7 1 2 55956 56931
0 5284 5 1 1 5283
0 5285 7 1 2 5280 5284
0 5286 5 1 1 5285
0 5287 7 1 2 53936 5286
0 5288 5 1 1 5287
0 5289 7 7 2 42933 49002
0 5290 5 1 1 56935
0 5291 7 1 2 43657 52418
0 5292 5 1 1 5291
0 5293 7 2 2 45247 5292
0 5294 5 1 1 56942
0 5295 7 1 2 56936 56943
0 5296 5 1 1 5295
0 5297 7 1 2 54647 49351
0 5298 5 1 1 5297
0 5299 7 1 2 5296 5298
0 5300 5 1 1 5299
0 5301 7 1 2 56616 5300
0 5302 5 1 1 5301
0 5303 7 4 2 42934 50943
0 5304 7 8 2 40169 56794
0 5305 7 1 2 48888 56948
0 5306 7 1 2 56944 5305
0 5307 5 1 1 5306
0 5308 7 1 2 5302 5307
0 5309 5 1 1 5308
0 5310 7 1 2 49182 5309
0 5311 5 1 1 5310
0 5312 7 11 2 44015 48468
0 5313 7 7 2 44171 44897
0 5314 7 4 2 45019 56967
0 5315 7 2 2 56956 56974
0 5316 7 1 2 48208 56978
0 5317 5 1 1 5316
0 5318 7 1 2 56871 50819
0 5319 5 16 1 5318
0 5320 7 1 2 42935 56980
0 5321 7 1 2 56751 5320
0 5322 5 1 1 5321
0 5323 7 1 2 5317 5322
0 5324 5 1 1 5323
0 5325 7 1 2 54648 5324
0 5326 5 1 1 5325
0 5327 7 1 2 5311 5326
0 5328 5 1 1 5327
0 5329 7 1 2 46339 5328
0 5330 5 1 1 5329
0 5331 7 3 2 39961 48574
0 5332 7 2 2 48469 56763
0 5333 7 1 2 56996 56999
0 5334 5 1 1 5333
0 5335 7 4 2 46340 49576
0 5336 7 16 2 44016 44172
0 5337 5 1 1 57005
0 5338 7 3 2 39962 57006
0 5339 7 1 2 57001 57021
0 5340 5 1 1 5339
0 5341 7 12 2 40924 43063
0 5342 7 1 2 57024 53327
0 5343 5 1 1 5342
0 5344 7 1 2 5340 5343
0 5345 5 1 1 5344
0 5346 7 1 2 52769 5345
0 5347 5 1 1 5346
0 5348 7 38 2 40925 54680
0 5349 5 11 1 57036
0 5350 7 3 2 48889 56828
0 5351 5 1 1 57085
0 5352 7 1 2 57074 5351
0 5353 5 11 1 5352
0 5354 7 7 2 48262 53528
0 5355 5 1 1 57099
0 5356 7 1 2 57088 57100
0 5357 5 1 1 5356
0 5358 7 3 2 49266 56440
0 5359 5 1 1 57106
0 5360 7 1 2 462 5359
0 5361 5 2 1 5360
0 5362 7 3 2 39963 46670
0 5363 5 1 1 57111
0 5364 7 1 2 57112 54665
0 5365 5 1 1 5364
0 5366 7 4 2 54591 52228
0 5367 7 1 2 42780 57114
0 5368 5 1 1 5367
0 5369 7 1 2 5365 5368
0 5370 5 1 1 5369
0 5371 7 1 2 57109 5370
0 5372 5 1 1 5371
0 5373 7 1 2 5357 5372
0 5374 7 1 2 5347 5373
0 5375 7 1 2 5334 5374
0 5376 5 1 1 5375
0 5377 7 1 2 52253 5376
0 5378 5 1 1 5377
0 5379 7 2 2 42936 54642
0 5380 7 3 2 52901 51467
0 5381 5 1 1 57120
0 5382 7 1 2 44173 57121
0 5383 5 1 1 5382
0 5384 7 5 2 44898 55168
0 5385 7 1 2 56981 57123
0 5386 5 1 1 5385
0 5387 7 1 2 5383 5386
0 5388 5 1 1 5387
0 5389 7 1 2 45020 5388
0 5390 5 1 1 5389
0 5391 7 1 2 48975 48957
0 5392 7 1 2 53505 5391
0 5393 5 1 1 5392
0 5394 7 1 2 5390 5393
0 5395 5 1 1 5394
0 5396 7 1 2 57118 5395
0 5397 5 1 1 5396
0 5398 7 3 2 46341 53529
0 5399 7 1 2 40350 48890
0 5400 7 1 2 57128 5399
0 5401 5 1 1 5400
0 5402 7 7 2 40170 44017
0 5403 7 3 2 53059 57131
0 5404 7 2 2 57025 54880
0 5405 7 1 2 57138 57141
0 5406 5 1 1 5405
0 5407 7 1 2 5401 5406
0 5408 5 1 1 5407
0 5409 7 1 2 48263 5408
0 5410 5 1 1 5409
0 5411 7 6 2 43870 44174
0 5412 7 7 2 48602 57143
0 5413 7 1 2 54643 57149
0 5414 5 1 1 5413
0 5415 7 5 2 40926 41445
0 5416 7 5 2 40747 57156
0 5417 7 9 2 40171 40577
0 5418 7 7 2 39964 43064
0 5419 7 1 2 57166 57175
0 5420 7 1 2 57161 5419
0 5421 5 1 1 5420
0 5422 7 1 2 5414 5421
0 5423 5 1 1 5422
0 5424 7 1 2 52770 5423
0 5425 5 1 1 5424
0 5426 7 2 2 52229 49127
0 5427 7 5 2 42781 54592
0 5428 7 1 2 55666 57184
0 5429 7 1 2 57182 5428
0 5430 5 1 1 5429
0 5431 7 1 2 5425 5430
0 5432 7 1 2 5410 5431
0 5433 7 1 2 5397 5432
0 5434 5 1 1 5433
0 5435 7 1 2 46733 5434
0 5436 5 1 1 5435
0 5437 7 1 2 5378 5436
0 5438 7 1 2 5330 5437
0 5439 7 1 2 5288 5438
0 5440 5 1 1 5439
0 5441 7 1 2 56913 5440
0 5442 5 1 1 5441
0 5443 7 32 2 43065 46447
0 5444 7 4 2 44899 42937
0 5445 7 4 2 57189 57221
0 5446 7 1 2 50105 57225
0 5447 5 1 1 5446
0 5448 7 11 2 41599 46218
0 5449 7 41 2 46342 43167
0 5450 7 4 2 46059 57240
0 5451 7 1 2 57229 57281
0 5452 5 1 1 5451
0 5453 7 1 2 5447 5452
0 5454 5 2 1 5453
0 5455 7 1 2 53276 57285
0 5456 5 1 1 5455
0 5457 7 10 2 46448 54976
0 5458 7 1 2 57287 53579
0 5459 7 1 2 52902 5458
0 5460 5 1 1 5459
0 5461 7 1 2 5456 5460
0 5462 5 1 1 5461
0 5463 7 1 2 41076 5462
0 5464 5 1 1 5463
0 5465 7 11 2 52634 57241
0 5466 7 1 2 53277 48355
0 5467 7 1 2 57297 5466
0 5468 5 1 1 5467
0 5469 7 1 2 5464 5468
0 5470 5 1 1 5469
0 5471 7 1 2 40748 5470
0 5472 5 1 1 5471
0 5473 7 1 2 53278 52903
0 5474 5 2 1 5473
0 5475 7 6 2 41600 53810
0 5476 5 2 1 57310
0 5477 7 1 2 57308 57316
0 5478 5 1 1 5477
0 5479 7 1 2 42938 5478
0 5480 5 1 1 5479
0 5481 7 1 2 48209 52131
0 5482 5 2 1 5481
0 5483 7 1 2 5480 57318
0 5484 5 2 1 5483
0 5485 7 5 2 44018 41077
0 5486 7 6 2 45248 57190
0 5487 7 1 2 57322 57327
0 5488 7 1 2 57320 5487
0 5489 5 1 1 5488
0 5490 7 1 2 5472 5489
0 5491 5 1 1 5490
0 5492 7 1 2 40578 5491
0 5493 5 1 1 5492
0 5494 7 3 2 41078 57328
0 5495 7 4 2 48210 51517
0 5496 5 1 1 57336
0 5497 7 1 2 3459 5496
0 5498 5 4 1 5497
0 5499 7 2 2 54348 57340
0 5500 5 1 1 57344
0 5501 7 1 2 57333 57345
0 5502 5 1 1 5501
0 5503 7 1 2 5493 5502
0 5504 5 1 1 5503
0 5505 7 1 2 53867 5504
0 5506 5 1 1 5505
0 5507 7 3 2 48100 53279
0 5508 5 2 1 57346
0 5509 7 1 2 57349 55206
0 5510 5 2 1 5509
0 5511 7 1 2 40579 57351
0 5512 5 1 1 5511
0 5513 7 1 2 54349 48211
0 5514 5 1 1 5513
0 5515 7 1 2 5512 5514
0 5516 5 2 1 5515
0 5517 7 2 2 41601 57353
0 5518 5 1 1 57355
0 5519 7 1 2 55226 56374
0 5520 5 1 1 5519
0 5521 7 1 2 5518 5520
0 5522 5 1 1 5521
0 5523 7 1 2 40749 5522
0 5524 5 1 1 5523
0 5525 7 6 2 40580 41602
0 5526 7 5 2 45841 53503
0 5527 7 2 2 57357 57363
0 5528 5 1 1 57368
0 5529 7 1 2 48212 57369
0 5530 5 1 1 5529
0 5531 7 1 2 5524 5530
0 5532 5 2 1 5531
0 5533 7 1 2 49003 57334
0 5534 7 1 2 57370 5533
0 5535 5 1 1 5534
0 5536 7 1 2 5506 5535
0 5537 5 1 1 5536
0 5538 7 1 2 40172 5537
0 5539 5 2 1 5538
0 5540 7 1 2 40173 57286
0 5541 5 1 1 5540
0 5542 7 5 2 40174 46449
0 5543 7 2 2 54977 48958
0 5544 7 1 2 57374 57379
0 5545 5 1 1 5544
0 5546 7 4 2 41603 57242
0 5547 7 2 2 46219 57381
0 5548 7 1 2 52707 57385
0 5549 5 1 1 5548
0 5550 7 1 2 5545 5549
0 5551 5 1 1 5550
0 5552 7 1 2 41079 5551
0 5553 5 1 1 5552
0 5554 7 1 2 5541 5553
0 5555 5 1 1 5554
0 5556 7 1 2 53280 5555
0 5557 5 1 1 5556
0 5558 7 9 2 42939 57191
0 5559 7 2 2 49313 57387
0 5560 7 3 2 42503 52904
0 5561 7 1 2 57396 57398
0 5562 5 1 1 5561
0 5563 7 1 2 5557 5562
0 5564 5 1 1 5563
0 5565 7 1 2 51453 5564
0 5566 5 1 1 5565
0 5567 7 1 2 53256 57321
0 5568 5 1 1 5567
0 5569 7 1 2 5500 5568
0 5570 5 1 1 5569
0 5571 7 6 2 43066 46734
0 5572 7 1 2 57401 57375
0 5573 7 1 2 5570 5572
0 5574 5 1 1 5573
0 5575 7 1 2 5566 5574
0 5576 5 1 1 5575
0 5577 7 1 2 41727 5576
0 5578 5 2 1 5577
0 5579 7 5 2 40175 45021
0 5580 7 2 2 46450 57409
0 5581 7 2 2 46220 57402
0 5582 7 2 2 41446 51724
0 5583 5 1 1 57418
0 5584 7 1 2 1628 5583
0 5585 5 1 1 5584
0 5586 7 1 2 40581 5585
0 5587 5 1 1 5586
0 5588 7 2 2 41604 54350
0 5589 5 1 1 57420
0 5590 7 1 2 5587 5589
0 5591 5 1 1 5590
0 5592 7 1 2 40750 5591
0 5593 5 1 1 5592
0 5594 7 1 2 5528 5593
0 5595 5 1 1 5594
0 5596 7 1 2 57416 5595
0 5597 5 1 1 5596
0 5598 7 2 2 53625 57323
0 5599 7 1 2 57422 54239
0 5600 7 1 2 55749 5599
0 5601 5 1 1 5600
0 5602 7 1 2 5597 5601
0 5603 5 1 1 5602
0 5604 7 1 2 42782 5603
0 5605 5 1 1 5604
0 5606 7 8 2 44900 56344
0 5607 7 1 2 45249 57424
0 5608 5 1 1 5607
0 5609 7 1 2 55384 5608
0 5610 5 1 1 5609
0 5611 7 1 2 48470 5610
0 5612 5 1 1 5611
0 5613 7 7 2 44750 45250
0 5614 7 3 2 46221 49183
0 5615 7 1 2 57432 57439
0 5616 5 1 1 5615
0 5617 7 1 2 5612 5616
0 5618 5 1 1 5617
0 5619 7 1 2 41080 5618
0 5620 5 1 1 5619
0 5621 7 6 2 42940 51468
0 5622 7 1 2 48356 57442
0 5623 5 1 1 5622
0 5624 7 1 2 5620 5623
0 5625 5 1 1 5624
0 5626 7 1 2 56686 5625
0 5627 5 1 1 5626
0 5628 7 1 2 5605 5627
0 5629 5 1 1 5628
0 5630 7 1 2 57414 5629
0 5631 5 1 1 5630
0 5632 7 1 2 57407 5631
0 5633 5 1 1 5632
0 5634 7 1 2 40927 5633
0 5635 5 1 1 5634
0 5636 7 8 2 40176 44175
0 5637 7 2 2 46451 57448
0 5638 7 1 2 41728 57403
0 5639 7 1 2 57371 5638
0 5640 5 2 1 5639
0 5641 7 2 2 44019 49852
0 5642 5 1 1 57460
0 5643 7 2 2 40751 50637
0 5644 5 1 1 57462
0 5645 7 1 2 5642 5644
0 5646 5 3 1 5645
0 5647 7 6 2 48575 56622
0 5648 5 1 1 57467
0 5649 7 17 2 46060 54593
0 5650 7 2 2 53281 57473
0 5651 5 2 1 57490
0 5652 7 1 2 5648 57492
0 5653 5 1 1 5652
0 5654 7 1 2 40582 5653
0 5655 5 2 1 5654
0 5656 7 1 2 53626 55399
0 5657 5 1 1 5656
0 5658 7 1 2 57494 5657
0 5659 5 1 1 5658
0 5660 7 1 2 57464 5659
0 5661 5 1 1 5660
0 5662 7 3 2 46343 52163
0 5663 7 9 2 42941 51518
0 5664 7 1 2 55593 57499
0 5665 7 1 2 57496 5664
0 5666 5 1 1 5665
0 5667 7 2 2 5661 5666
0 5668 7 1 2 55416 50140
0 5669 5 1 1 5668
0 5670 7 1 2 41447 55227
0 5671 5 3 1 5670
0 5672 7 1 2 57510 53846
0 5673 5 2 1 5672
0 5674 7 1 2 40583 57513
0 5675 5 1 1 5674
0 5676 7 1 2 4859 5675
0 5677 5 4 1 5676
0 5678 7 1 2 54666 57515
0 5679 5 1 1 5678
0 5680 7 1 2 5669 5679
0 5681 5 1 1 5680
0 5682 7 1 2 49184 5681
0 5683 5 1 1 5682
0 5684 7 1 2 57508 5683
0 5685 5 1 1 5684
0 5686 7 1 2 46788 5685
0 5687 5 1 1 5686
0 5688 7 1 2 57458 5687
0 5689 5 1 1 5688
0 5690 7 1 2 57456 5689
0 5691 5 1 1 5690
0 5692 7 1 2 5635 5691
0 5693 5 1 1 5692
0 5694 7 1 2 39965 5693
0 5695 5 1 1 5694
0 5696 7 1 2 57372 5695
0 5697 5 1 1 5696
0 5698 7 1 2 40351 5697
0 5699 5 1 1 5698
0 5700 7 1 2 57037 53328
0 5701 5 1 1 5700
0 5702 7 3 2 45022 49128
0 5703 5 1 1 57519
0 5704 7 1 2 49004 49277
0 5705 5 1 1 5704
0 5706 7 1 2 5703 5705
0 5707 5 1 1 5706
0 5708 7 1 2 46344 55155
0 5709 7 1 2 5707 5708
0 5710 5 1 1 5709
0 5711 7 1 2 5701 5710
0 5712 5 1 1 5711
0 5713 7 1 2 52905 5712
0 5714 5 1 1 5713
0 5715 7 5 2 45023 56456
0 5716 7 1 2 52708 57522
0 5717 5 1 1 5716
0 5718 7 1 2 55156 48959
0 5719 7 1 2 49005 5718
0 5720 5 1 1 5719
0 5721 7 1 2 5717 5720
0 5722 5 1 1 5721
0 5723 7 1 2 57129 5722
0 5724 5 1 1 5723
0 5725 7 1 2 5714 5724
0 5726 5 1 1 5725
0 5727 7 1 2 42942 5726
0 5728 5 1 1 5727
0 5729 7 2 2 54133 51146
0 5730 5 1 1 57527
0 5731 7 1 2 54023 5730
0 5732 5 1 1 5731
0 5733 7 1 2 57101 5732
0 5734 5 1 1 5733
0 5735 7 3 2 41605 48213
0 5736 7 2 2 43067 56493
0 5737 5 1 1 57532
0 5738 7 1 2 56481 57528
0 5739 5 1 1 5738
0 5740 7 1 2 5737 5739
0 5741 5 1 1 5740
0 5742 7 1 2 57529 5741
0 5743 5 1 1 5742
0 5744 7 1 2 5734 5743
0 5745 7 1 2 5728 5744
0 5746 5 1 1 5745
0 5747 7 1 2 56914 5746
0 5748 5 1 1 5747
0 5749 7 1 2 5699 5748
0 5750 5 1 1 5749
0 5751 7 1 2 47004 5750
0 5752 5 1 1 5751
0 5753 7 1 2 5442 5752
0 5754 5 1 1 5753
0 5755 7 1 2 46606 5754
0 5756 5 1 1 5755
0 5757 7 3 2 46452 46645
0 5758 7 1 2 49768 47067
0 5759 5 2 1 5758
0 5760 7 1 2 5294 57537
0 5761 5 1 1 5760
0 5762 7 6 2 46222 55814
0 5763 7 1 2 49170 53362
0 5764 5 1 1 5763
0 5765 7 6 2 2541 5764
0 5766 7 2 2 57539 57545
0 5767 7 1 2 5761 57551
0 5768 5 1 1 5767
0 5769 7 1 2 53811 50409
0 5770 5 2 1 5769
0 5771 7 2 2 41081 53249
0 5772 7 1 2 57167 54240
0 5773 7 1 2 56465 5772
0 5774 7 1 2 57555 5773
0 5775 5 1 1 5774
0 5776 7 1 2 57553 5775
0 5777 5 1 1 5776
0 5778 7 1 2 40752 5777
0 5779 5 1 1 5778
0 5780 7 1 2 51871 55962
0 5781 5 1 1 5780
0 5782 7 1 2 48544 5781
0 5783 5 1 1 5782
0 5784 7 1 2 42504 5783
0 5785 5 1 1 5784
0 5786 7 1 2 45251 50243
0 5787 7 1 2 56213 5786
0 5788 5 1 1 5787
0 5789 7 1 2 5785 5788
0 5790 5 2 1 5789
0 5791 7 1 2 55287 57557
0 5792 5 1 1 5791
0 5793 7 1 2 5779 5792
0 5794 5 1 1 5793
0 5795 7 1 2 39966 5794
0 5796 5 1 1 5795
0 5797 7 2 2 53530 57311
0 5798 7 1 2 52266 57559
0 5799 5 1 1 5798
0 5800 7 1 2 5796 5799
0 5801 5 1 1 5800
0 5802 7 1 2 40352 5801
0 5803 5 1 1 5802
0 5804 7 1 2 52267 47005
0 5805 5 1 1 5804
0 5806 7 1 2 52083 5805
0 5807 5 1 1 5806
0 5808 7 1 2 57560 5807
0 5809 5 1 1 5808
0 5810 7 1 2 55157 47068
0 5811 5 1 1 5810
0 5812 7 1 2 52348 5811
0 5813 5 1 1 5812
0 5814 7 2 2 48471 54487
0 5815 5 2 1 57561
0 5816 7 1 2 5813 57562
0 5817 5 1 1 5816
0 5818 7 14 2 39967 40353
0 5819 7 4 2 52063 47006
0 5820 5 2 1 57579
0 5821 7 1 2 57565 57580
0 5822 7 1 2 54520 5821
0 5823 5 1 1 5822
0 5824 7 1 2 5817 5823
0 5825 5 1 1 5824
0 5826 7 1 2 52906 5825
0 5827 5 1 1 5826
0 5828 7 1 2 5809 5827
0 5829 7 1 2 5803 5828
0 5830 5 1 1 5829
0 5831 7 1 2 42943 5830
0 5832 5 1 1 5831
0 5833 7 1 2 5768 5832
0 5834 5 1 1 5833
0 5835 7 1 2 41729 5834
0 5836 5 1 1 5835
0 5837 7 5 2 40354 45252
0 5838 5 1 1 57585
0 5839 7 1 2 52349 5838
0 5840 7 1 2 57538 5839
0 5841 5 1 1 5840
0 5842 7 1 2 57540 5841
0 5843 5 1 1 5842
0 5844 7 15 2 45842 48101
0 5845 7 1 2 50179 57590
0 5846 7 1 2 55960 5845
0 5847 5 1 1 5846
0 5848 7 1 2 5843 5847
0 5849 5 2 1 5848
0 5850 7 1 2 41606 51477
0 5851 7 1 2 57605 5850
0 5852 5 1 1 5851
0 5853 7 1 2 5836 5852
0 5854 5 1 1 5853
0 5855 7 1 2 40928 5854
0 5856 5 1 1 5855
0 5857 7 1 2 57183 57606
0 5858 5 1 1 5857
0 5859 7 1 2 5856 5858
0 5860 5 1 1 5859
0 5861 7 1 2 46345 5860
0 5862 5 1 1 5861
0 5863 7 4 2 57566 57168
0 5864 7 1 2 51740 56643
0 5865 7 1 2 57607 5864
0 5866 7 3 2 40753 51217
0 5867 7 5 2 40929 52833
0 5868 7 1 2 53539 57614
0 5869 7 1 2 57611 5868
0 5870 7 1 2 5865 5869
0 5871 5 1 1 5870
0 5872 7 1 2 5862 5871
0 5873 5 1 1 5872
0 5874 7 1 2 57534 5873
0 5875 5 1 1 5874
0 5876 7 1 2 5756 5875
0 5877 5 1 1 5876
0 5878 7 49 2 44226 45068
0 5879 5 5 1 57619
0 5880 7 1 2 57668 48846
0 5881 7 1 2 5877 5880
0 5882 5 1 1 5881
0 5883 7 1 2 46061 49171
0 5884 5 1 1 5883
0 5885 7 1 2 48087 1949
0 5886 5 1 1 5885
0 5887 7 1 2 41082 5886
0 5888 7 1 2 5884 5887
0 5889 5 1 1 5888
0 5890 7 1 2 51322 48357
0 5891 5 1 1 5890
0 5892 7 1 2 5889 5891
0 5893 5 1 1 5892
0 5894 7 1 2 54594 5893
0 5895 5 1 1 5894
0 5896 7 2 2 44901 57324
0 5897 7 1 2 53627 50106
0 5898 7 1 2 57673 5897
0 5899 5 1 1 5898
0 5900 7 1 2 5895 5899
0 5901 5 1 1 5900
0 5902 7 1 2 55750 5901
0 5903 5 1 1 5902
0 5904 7 1 2 46735 48303
0 5905 5 1 1 5904
0 5906 7 2 2 41083 52713
0 5907 7 1 2 56345 57675
0 5908 5 1 1 5907
0 5909 7 1 2 5905 5908
0 5910 5 1 1 5909
0 5911 7 13 2 45843 43068
0 5912 7 1 2 48472 57677
0 5913 7 1 2 5910 5912
0 5914 5 1 1 5913
0 5915 7 1 2 5903 5914
0 5916 5 1 1 5915
0 5917 7 1 2 57415 5916
0 5918 5 1 1 5917
0 5919 7 1 2 57408 5918
0 5920 5 1 1 5919
0 5921 7 1 2 40930 5920
0 5922 5 1 1 5921
0 5923 7 3 2 55228 53628
0 5924 7 1 2 57690 52206
0 5925 5 1 1 5924
0 5926 7 1 2 46062 55751
0 5927 7 1 2 56640 5926
0 5928 5 1 1 5927
0 5929 7 1 2 5925 5928
0 5930 5 1 1 5929
0 5931 7 1 2 49185 5930
0 5932 5 1 1 5931
0 5933 7 1 2 5932 57509
0 5934 5 1 1 5933
0 5935 7 1 2 46789 5934
0 5936 5 1 1 5935
0 5937 7 1 2 5936 57459
0 5938 5 1 1 5937
0 5939 7 1 2 57457 5938
0 5940 5 1 1 5939
0 5941 7 1 2 5922 5940
0 5942 5 1 1 5941
0 5943 7 1 2 39968 5942
0 5944 5 1 1 5943
0 5945 7 1 2 5944 57373
0 5946 5 1 1 5945
0 5947 7 1 2 41330 5946
0 5948 5 1 1 5947
0 5949 7 5 2 44751 56609
0 5950 7 3 2 41084 46346
0 5951 5 1 1 57698
0 5952 7 2 2 48891 57699
0 5953 5 1 1 57701
0 5954 7 4 2 41902 51519
0 5955 7 1 2 57702 57703
0 5956 7 1 2 57693 5955
0 5957 5 1 1 5956
0 5958 7 1 2 48473 49186
0 5959 5 2 1 5958
0 5960 7 7 2 54439 50731
0 5961 5 1 1 57709
0 5962 7 1 2 57707 5961
0 5963 5 5 1 5962
0 5964 7 1 2 49006 57716
0 5965 5 1 1 5964
0 5966 7 10 2 40931 44902
0 5967 7 3 2 57721 49278
0 5968 7 1 2 41730 57731
0 5969 5 1 1 5968
0 5970 7 1 2 5965 5969
0 5971 5 2 1 5970
0 5972 7 1 2 43069 55158
0 5973 7 1 2 57734 5972
0 5974 5 1 1 5973
0 5975 7 1 2 5957 5974
0 5976 5 1 1 5975
0 5977 7 2 2 46063 46453
0 5978 7 1 2 54869 57736
0 5979 7 1 2 5976 5978
0 5980 5 1 1 5979
0 5981 7 1 2 5948 5980
0 5982 5 1 1 5981
0 5983 7 1 2 45623 5982
0 5984 5 1 1 5983
0 5985 7 4 2 41085 53937
0 5986 5 2 1 57738
0 5987 7 1 2 57075 5953
0 5988 5 3 1 5987
0 5989 7 2 2 39969 57744
0 5990 5 1 1 57747
0 5991 7 1 2 57742 5990
0 5992 5 2 1 5991
0 5993 7 5 2 44903 48102
0 5994 7 1 2 48474 57751
0 5995 5 2 1 5994
0 5996 7 1 2 56926 57756
0 5997 5 1 1 5996
0 5998 7 1 2 57749 5997
0 5999 5 1 1 5998
0 6000 7 3 2 56655 50638
0 6001 5 1 1 57758
0 6002 7 5 2 44176 41086
0 6003 7 5 2 39970 57761
0 6004 7 1 2 48475 57766
0 6005 7 1 2 57759 6004
0 6006 5 1 1 6005
0 6007 7 1 2 5999 6006
0 6008 5 1 1 6007
0 6009 7 1 2 45253 6008
0 6010 5 1 1 6009
0 6011 7 2 2 46064 54978
0 6012 7 3 2 41087 41448
0 6013 7 1 2 53060 57773
0 6014 7 1 2 56225 6013
0 6015 7 1 2 57771 6014
0 6016 5 1 1 6015
0 6017 7 1 2 6010 6016
0 6018 5 1 1 6017
0 6019 7 1 2 40754 6018
0 6020 5 1 1 6019
0 6021 7 3 2 53629 50618
0 6022 5 1 1 57776
0 6023 7 4 2 43871 41088
0 6024 7 2 2 45254 57779
0 6025 5 1 1 57783
0 6026 7 1 2 57777 57784
0 6027 5 1 1 6026
0 6028 7 1 2 55594 57417
0 6029 5 1 1 6028
0 6030 7 1 2 6027 6029
0 6031 5 1 1 6030
0 6032 7 1 2 39971 6031
0 6033 5 1 1 6032
0 6034 7 6 2 48476 57474
0 6035 5 2 1 57785
0 6036 7 2 2 46790 57786
0 6037 5 1 1 57793
0 6038 7 1 2 6033 6037
0 6039 5 1 1 6038
0 6040 7 1 2 49187 6039
0 6041 5 1 1 6040
0 6042 7 5 2 48049 48477
0 6043 7 3 2 57185 57795
0 6044 5 1 1 57800
0 6045 7 1 2 47268 57801
0 6046 5 1 1 6045
0 6047 7 2 2 45255 56982
0 6048 7 12 2 53630 51520
0 6049 5 1 1 57805
0 6050 7 2 2 47269 57806
0 6051 5 1 1 57817
0 6052 7 8 2 48050 54595
0 6053 5 4 1 57819
0 6054 7 1 2 47458 57820
0 6055 5 1 1 6054
0 6056 7 1 2 6051 6055
0 6057 5 1 1 6056
0 6058 7 1 2 57803 6057
0 6059 5 1 1 6058
0 6060 7 1 2 6046 6059
0 6061 7 1 2 6041 6060
0 6062 5 1 1 6061
0 6063 7 1 2 49007 6062
0 6064 5 1 1 6063
0 6065 7 1 2 6020 6064
0 6066 5 1 1 6065
0 6067 7 1 2 40177 6066
0 6068 5 1 1 6067
0 6069 7 6 2 45256 48892
0 6070 7 4 2 57831 57700
0 6071 5 3 1 57837
0 6072 7 1 2 53868 57404
0 6073 5 2 1 6072
0 6074 7 1 2 57841 57844
0 6075 5 4 1 6074
0 6076 7 4 2 57169 50866
0 6077 5 1 1 57850
0 6078 7 1 2 57846 57851
0 6079 5 1 1 6078
0 6080 7 10 2 42286 46347
0 6081 7 2 2 48893 57854
0 6082 7 1 2 50029 57864
0 6083 5 1 1 6082
0 6084 7 2 2 52319 57038
0 6085 5 1 1 57866
0 6086 7 1 2 6083 6085
0 6087 5 1 1 6086
0 6088 7 1 2 50806 6087
0 6089 5 1 1 6088
0 6090 7 1 2 6079 6089
0 6091 5 1 1 6090
0 6092 7 1 2 39972 6091
0 6093 5 1 1 6092
0 6094 7 1 2 50775 51391
0 6095 5 1 1 6094
0 6096 7 1 2 52391 57804
0 6097 5 1 1 6096
0 6098 7 1 2 6095 6097
0 6099 5 1 1 6098
0 6100 7 1 2 53938 6099
0 6101 5 1 1 6100
0 6102 7 1 2 6093 6101
0 6103 5 1 1 6102
0 6104 7 1 2 44904 6103
0 6105 5 1 1 6104
0 6106 7 1 2 55770 50112
0 6107 7 1 2 57750 6106
0 6108 5 1 1 6107
0 6109 7 1 2 6105 6108
0 6110 5 1 1 6109
0 6111 7 1 2 46223 6110
0 6112 5 1 1 6111
0 6113 7 3 2 40932 46791
0 6114 7 1 2 54681 57868
0 6115 5 2 1 6114
0 6116 7 1 2 39973 57847
0 6117 5 1 1 6116
0 6118 7 1 2 57871 6117
0 6119 5 1 1 6118
0 6120 7 1 2 57170 56436
0 6121 7 1 2 6119 6120
0 6122 5 1 1 6121
0 6123 7 1 2 6112 6122
0 6124 5 1 1 6123
0 6125 7 1 2 44020 6124
0 6126 5 1 1 6125
0 6127 7 2 2 49188 57787
0 6128 5 1 1 57873
0 6129 7 2 2 49080 53519
0 6130 5 2 1 57875
0 6131 7 1 2 54596 57876
0 6132 5 2 1 6131
0 6133 7 1 2 6128 57879
0 6134 5 1 1 6133
0 6135 7 1 2 41331 49008
0 6136 7 1 2 6134 6135
0 6137 5 1 1 6136
0 6138 7 1 2 6126 6137
0 6139 7 1 2 6068 6138
0 6140 5 1 1 6139
0 6141 7 1 2 56915 6140
0 6142 5 1 1 6141
0 6143 7 1 2 5984 6142
0 6144 5 1 1 6143
0 6145 7 1 2 40974 6144
0 6146 5 1 1 6145
0 6147 7 1 2 55024 6146
0 6148 5 1 1 6147
0 6149 7 2 2 55295 50649
0 6150 7 1 2 41332 57881
0 6151 5 1 1 6150
0 6152 7 1 2 6151 5381
0 6153 5 1 1 6152
0 6154 7 1 2 42944 6153
0 6155 5 1 1 6154
0 6156 7 2 2 5355 56933
0 6157 7 1 2 6155 57883
0 6158 5 1 1 6157
0 6159 7 1 2 42505 6158
0 6160 5 1 1 6159
0 6161 7 1 2 53508 2656
0 6162 5 7 1 6161
0 6163 7 1 2 52907 57885
0 6164 5 1 1 6163
0 6165 7 1 2 56856 48428
0 6166 5 3 1 6165
0 6167 7 2 2 6164 57892
0 6168 5 1 1 57895
0 6169 7 1 2 44752 55288
0 6170 5 1 1 6169
0 6171 7 1 2 57896 6170
0 6172 5 2 1 6171
0 6173 7 3 2 42945 57897
0 6174 5 2 1 57899
0 6175 7 1 2 56147 57900
0 6176 5 1 1 6175
0 6177 7 1 2 6160 6176
0 6178 5 1 1 6177
0 6179 7 1 2 52320 6178
0 6180 5 1 1 6179
0 6181 7 6 2 44905 54870
0 6182 7 2 2 50678 54785
0 6183 5 9 1 57910
0 6184 7 2 2 46065 57912
0 6185 7 2 2 57904 57921
0 6186 5 1 1 57923
0 6187 7 1 2 49279 57924
0 6188 5 1 1 6187
0 6189 7 1 2 6180 6188
0 6190 5 1 1 6189
0 6191 7 1 2 53869 6190
0 6192 5 1 1 6191
0 6193 7 2 2 45257 55208
0 6194 7 1 2 52790 57925
0 6195 5 1 1 6194
0 6196 7 1 2 6186 6195
0 6197 5 1 1 6196
0 6198 7 1 2 51469 6197
0 6199 5 1 1 6198
0 6200 7 1 2 53812 57230
0 6201 7 1 2 57913 6200
0 6202 7 4 2 40755 49637
0 6203 5 3 1 57927
0 6204 7 1 2 44021 48545
0 6205 5 7 1 6204
0 6206 7 1 2 57931 57934
0 6207 7 1 2 6201 6206
0 6208 5 1 1 6207
0 6209 7 1 2 6199 6208
0 6210 5 1 1 6209
0 6211 7 1 2 49009 6210
0 6212 5 1 1 6211
0 6213 7 1 2 6192 6212
0 6214 5 1 1 6213
0 6215 7 1 2 46348 6214
0 6216 5 1 1 6215
0 6217 7 3 2 45844 52635
0 6218 7 5 2 40178 43070
0 6219 7 3 2 57941 57944
0 6220 7 3 2 52508 56713
0 6221 7 1 2 57952 51454
0 6222 7 1 2 56126 6221
0 6223 7 1 2 57949 6222
0 6224 5 1 1 6223
0 6225 7 1 2 6216 6224
0 6226 5 1 1 6225
0 6227 7 1 2 46454 47270
0 6228 7 1 2 6226 6227
0 6229 5 1 1 6228
0 6230 7 1 2 46646 6229
0 6231 5 1 1 6230
0 6232 7 1 2 47069 6231
0 6233 7 1 2 6148 6232
0 6234 5 1 1 6233
0 6235 7 10 2 46224 46349
0 6236 7 6 2 43168 57955
0 6237 7 10 2 45624 55406
0 6238 7 3 2 57965 57971
0 6239 5 1 1 57981
0 6240 7 2 2 40975 41731
0 6241 7 5 2 41196 41773
0 6242 7 3 2 57984 57986
0 6243 7 1 2 50275 51218
0 6244 7 1 2 57991 6243
0 6245 7 1 2 56601 6244
0 6246 7 1 2 57982 6245
0 6247 5 1 1 6246
0 6248 7 1 2 6234 6247
0 6249 7 1 2 5882 6248
0 6250 7 1 2 5264 6249
0 6251 5 1 1 6250
0 6252 7 1 2 46558 6251
0 6253 5 1 1 6252
0 6254 7 11 2 43872 41449
0 6255 5 1 1 57994
0 6256 7 10 2 40584 44753
0 6257 5 1 1 58005
0 6258 7 2 2 6255 6257
0 6259 5 48 1 58015
0 6260 7 1 2 54424 50261
0 6261 5 1 1 6260
0 6262 7 1 2 2458 6261
0 6263 5 1 1 6262
0 6264 7 1 2 41333 6263
0 6265 5 1 1 6264
0 6266 7 2 2 43658 53679
0 6267 5 4 1 58065
0 6268 7 1 2 42287 50951
0 6269 5 1 1 6268
0 6270 7 1 2 48654 6269
0 6271 5 1 1 6270
0 6272 7 1 2 54776 56200
0 6273 5 1 1 6272
0 6274 7 1 2 50606 6273
0 6275 5 2 1 6274
0 6276 7 1 2 6271 58071
0 6277 5 1 1 6276
0 6278 7 1 2 58067 6277
0 6279 5 1 1 6278
0 6280 7 1 2 42506 6279
0 6281 5 1 1 6280
0 6282 7 3 2 41903 54035
0 6283 7 1 2 55550 58073
0 6284 5 1 1 6283
0 6285 7 1 2 6281 6284
0 6286 5 1 1 6285
0 6287 7 1 2 41607 6286
0 6288 5 1 1 6287
0 6289 7 1 2 6265 6288
0 6290 5 1 1 6289
0 6291 7 1 2 40756 6290
0 6292 5 1 1 6291
0 6293 7 3 2 41334 41608
0 6294 7 1 2 50475 54468
0 6295 7 1 2 58076 6294
0 6296 5 1 1 6295
0 6297 7 1 2 6292 6296
0 6298 5 1 1 6297
0 6299 7 1 2 47623 6298
0 6300 5 1 1 6299
0 6301 7 1 2 47459 51122
0 6302 5 6 1 6301
0 6303 7 1 2 47624 58079
0 6304 5 5 1 6303
0 6305 7 2 2 40355 58085
0 6306 5 2 1 58090
0 6307 7 1 2 52470 58091
0 6308 5 1 1 6307
0 6309 7 3 2 47039 47566
0 6310 5 4 1 58094
0 6311 7 1 2 3560 53735
0 6312 5 1 1 6311
0 6313 7 1 2 42288 6312
0 6314 5 1 1 6313
0 6315 7 1 2 55933 6314
0 6316 5 1 1 6315
0 6317 7 1 2 58097 6316
0 6318 5 1 1 6317
0 6319 7 1 2 47577 54569
0 6320 5 3 1 6319
0 6321 7 3 2 47712 46832
0 6322 5 5 1 58104
0 6323 7 1 2 49950 58105
0 6324 5 1 1 6323
0 6325 7 1 2 40356 6324
0 6326 5 1 1 6325
0 6327 7 1 2 49700 6326
0 6328 5 1 1 6327
0 6329 7 1 2 41335 6328
0 6330 5 1 1 6329
0 6331 7 1 2 58101 6330
0 6332 5 1 1 6331
0 6333 7 1 2 42289 6332
0 6334 5 1 1 6333
0 6335 7 1 2 42054 592
0 6336 5 1 1 6335
0 6337 7 1 2 42055 58107
0 6338 5 1 1 6337
0 6339 7 2 2 6338 46966
0 6340 7 1 2 50165 58112
0 6341 5 1 1 6340
0 6342 7 1 2 49472 6341
0 6343 5 1 1 6342
0 6344 7 1 2 6336 6343
0 6345 5 1 1 6344
0 6346 7 1 2 45625 6345
0 6347 5 1 1 6346
0 6348 7 1 2 6334 6347
0 6349 7 1 2 6318 6348
0 6350 5 1 1 6349
0 6351 7 1 2 45845 6350
0 6352 5 1 1 6351
0 6353 7 1 2 6308 6352
0 6354 5 1 1 6353
0 6355 7 1 2 49189 6354
0 6356 5 1 1 6355
0 6357 7 1 2 42290 55907
0 6358 5 1 1 6357
0 6359 7 1 2 40357 55704
0 6360 5 4 1 6359
0 6361 7 1 2 41904 58114
0 6362 5 1 1 6361
0 6363 7 1 2 47713 50449
0 6364 5 2 1 6363
0 6365 7 1 2 45626 58118
0 6366 7 1 2 6362 6365
0 6367 5 1 1 6366
0 6368 7 1 2 44621 6367
0 6369 7 1 2 6358 6368
0 6370 5 1 1 6369
0 6371 7 2 2 47714 47874
0 6372 5 3 1 58120
0 6373 7 1 2 49878 55713
0 6374 5 1 1 6373
0 6375 7 1 2 58122 6374
0 6376 5 1 1 6375
0 6377 7 1 2 41905 6376
0 6378 5 1 1 6377
0 6379 7 3 2 43320 50671
0 6380 5 2 1 58125
0 6381 7 1 2 44396 58126
0 6382 5 1 1 6381
0 6383 7 1 2 58123 6382
0 6384 5 1 1 6383
0 6385 7 1 2 42056 6384
0 6386 5 1 1 6385
0 6387 7 1 2 6378 6386
0 6388 7 1 2 6370 6387
0 6389 5 1 1 6388
0 6390 7 1 2 42507 6389
0 6391 5 1 1 6390
0 6392 7 5 2 45846 51033
0 6393 7 1 2 50831 49935
0 6394 5 1 1 6393
0 6395 7 1 2 50981 6394
0 6396 5 1 1 6395
0 6397 7 1 2 58130 6396
0 6398 5 1 1 6397
0 6399 7 1 2 6391 6398
0 6400 5 1 1 6399
0 6401 7 1 2 48051 6400
0 6402 5 1 1 6401
0 6403 7 1 2 6356 6402
0 6404 7 1 2 6300 6403
0 6405 5 1 1 6404
0 6406 7 1 2 46066 6405
0 6407 5 1 1 6406
0 6408 7 1 2 40358 48847
0 6409 5 3 1 6408
0 6410 7 6 2 52019 58135
0 6411 7 1 2 58098 48871
0 6412 5 1 1 6411
0 6413 7 1 2 58138 6412
0 6414 5 2 1 6413
0 6415 7 2 2 47546 58144
0 6416 7 2 2 55229 58146
0 6417 5 1 1 58148
0 6418 7 1 2 48052 58149
0 6419 5 1 1 6418
0 6420 7 1 2 6407 6419
0 6421 5 1 1 6420
0 6422 7 1 2 49010 6421
0 6423 5 1 1 6422
0 6424 7 3 2 42057 51820
0 6425 5 2 1 58150
0 6426 7 1 2 55853 58151
0 6427 5 1 1 6426
0 6428 7 1 2 55868 54722
0 6429 5 1 1 6428
0 6430 7 1 2 43513 6429
0 6431 5 1 1 6430
0 6432 7 1 2 47040 54700
0 6433 5 1 1 6432
0 6434 7 1 2 54738 6433
0 6435 7 1 2 6431 6434
0 6436 5 1 1 6435
0 6437 7 1 2 42508 6436
0 6438 5 1 1 6437
0 6439 7 1 2 6427 6438
0 6440 5 1 1 6439
0 6441 7 1 2 42291 6440
0 6442 5 1 1 6441
0 6443 7 4 2 44485 47389
0 6444 5 2 1 58155
0 6445 7 1 2 40359 58159
0 6446 5 4 1 6445
0 6447 7 1 2 40179 46989
0 6448 5 2 1 6447
0 6449 7 1 2 42058 52437
0 6450 7 1 2 58165 6449
0 6451 7 1 2 58161 6450
0 6452 5 1 1 6451
0 6453 7 1 2 6442 6452
0 6454 5 1 1 6453
0 6455 7 1 2 41609 6454
0 6456 5 1 1 6455
0 6457 7 1 2 51725 58147
0 6458 5 1 1 6457
0 6459 7 1 2 6456 6458
0 6460 5 1 1 6459
0 6461 7 1 2 44022 6460
0 6462 5 1 1 6461
0 6463 7 2 2 52173 51184
0 6464 5 2 1 58167
0 6465 7 1 2 52466 58169
0 6466 5 3 1 6465
0 6467 7 2 2 43514 58171
0 6468 5 1 1 58174
0 6469 7 1 2 52438 47041
0 6470 5 1 1 6469
0 6471 7 1 2 6468 6470
0 6472 5 1 1 6471
0 6473 7 1 2 49160 6472
0 6474 5 1 1 6473
0 6475 7 1 2 51913 48429
0 6476 7 1 2 51705 6475
0 6477 5 1 1 6476
0 6478 7 1 2 6474 6477
0 6479 5 1 1 6478
0 6480 7 1 2 47390 6479
0 6481 5 1 1 6480
0 6482 7 4 2 44023 44486
0 6483 7 1 2 56036 58176
0 6484 7 1 2 50794 6483
0 6485 5 1 1 6484
0 6486 7 1 2 6481 6485
0 6487 5 1 1 6486
0 6488 7 1 2 48729 6487
0 6489 5 1 1 6488
0 6490 7 4 2 51914 51363
0 6491 7 3 2 44397 44906
0 6492 7 1 2 58184 55792
0 6493 7 1 2 58180 6492
0 6494 5 1 1 6493
0 6495 7 1 2 6489 6494
0 6496 7 1 2 6462 6495
0 6497 5 1 1 6496
0 6498 7 1 2 40933 6497
0 6499 5 1 1 6498
0 6500 7 3 2 41610 49103
0 6501 7 1 2 48848 47988
0 6502 7 4 2 50505 6501
0 6503 5 1 1 58190
0 6504 7 1 2 58136 2187
0 6505 7 2 2 6503 6504
0 6506 5 1 1 58194
0 6507 7 1 2 40180 6506
0 6508 5 2 1 6507
0 6509 7 1 2 47115 48849
0 6510 5 2 1 6509
0 6511 7 2 2 52020 58198
0 6512 5 1 1 58200
0 6513 7 1 2 52247 52041
0 6514 7 1 2 6512 6513
0 6515 5 1 1 6514
0 6516 7 1 2 58196 6515
0 6517 5 2 1 6516
0 6518 7 2 2 45847 58202
0 6519 7 1 2 58187 58204
0 6520 5 1 1 6519
0 6521 7 1 2 6499 6520
0 6522 5 1 1 6521
0 6523 7 1 2 42783 6522
0 6524 5 1 1 6523
0 6525 7 2 2 55169 46671
0 6526 7 1 2 41906 55927
0 6527 5 1 1 6526
0 6528 7 1 2 49829 6527
0 6529 5 1 1 6528
0 6530 7 1 2 45627 6529
0 6531 5 1 1 6530
0 6532 7 1 2 41336 54954
0 6533 5 1 1 6532
0 6534 7 1 2 6531 6533
0 6535 5 1 1 6534
0 6536 7 1 2 42059 6535
0 6537 5 1 1 6536
0 6538 7 5 2 40181 50180
0 6539 5 5 1 58208
0 6540 7 1 2 45418 58213
0 6541 5 2 1 6540
0 6542 7 1 2 42292 58218
0 6543 7 1 2 55905 6542
0 6544 5 1 1 6543
0 6545 7 2 2 51840 47140
0 6546 5 4 1 58220
0 6547 7 1 2 47391 51883
0 6548 5 1 1 6547
0 6549 7 2 2 58221 6548
0 6550 5 1 1 58226
0 6551 7 1 2 41907 6550
0 6552 5 1 1 6551
0 6553 7 1 2 47145 58166
0 6554 5 1 1 6553
0 6555 7 1 2 45628 6554
0 6556 7 1 2 6552 6555
0 6557 5 1 1 6556
0 6558 7 1 2 44622 6557
0 6559 7 1 2 6544 6558
0 6560 5 1 1 6559
0 6561 7 2 2 42293 47625
0 6562 5 2 1 58228
0 6563 7 1 2 50157 58229
0 6564 5 1 1 6563
0 6565 7 1 2 43659 50580
0 6566 5 2 1 6565
0 6567 7 1 2 58232 53586
0 6568 5 1 1 6567
0 6569 7 1 2 41908 56248
0 6570 7 1 2 6568 6569
0 6571 5 1 1 6570
0 6572 7 1 2 6564 6571
0 6573 7 1 2 6560 6572
0 6574 7 1 2 6537 6573
0 6575 5 1 1 6574
0 6576 7 1 2 42509 6575
0 6577 5 1 1 6576
0 6578 7 1 2 51760 707
0 6579 5 1 1 6578
0 6580 7 1 2 41909 6579
0 6581 5 1 1 6580
0 6582 7 1 2 50982 6581
0 6583 5 1 1 6582
0 6584 7 1 2 58131 6583
0 6585 5 1 1 6584
0 6586 7 1 2 6577 6585
0 6587 5 1 1 6586
0 6588 7 1 2 58206 6587
0 6589 5 1 1 6588
0 6590 7 1 2 6524 6589
0 6591 5 1 1 6590
0 6592 7 1 2 41732 6591
0 6593 5 1 1 6592
0 6594 7 1 2 6423 6593
0 6595 5 1 1 6594
0 6596 7 1 2 46225 6595
0 6597 5 1 1 6596
0 6598 7 1 2 50843 58145
0 6599 5 2 1 6598
0 6600 7 2 2 50368 50925
0 6601 5 1 1 58236
0 6602 7 1 2 54759 58237
0 6603 5 1 1 6602
0 6604 7 1 2 58234 6603
0 6605 5 1 1 6604
0 6606 7 1 2 55296 6605
0 6607 5 1 1 6606
0 6608 7 7 2 45419 47578
0 6609 7 1 2 48872 46672
0 6610 5 1 1 6609
0 6611 7 10 2 45258 47271
0 6612 5 4 1 58245
0 6613 7 1 2 58246 52908
0 6614 5 1 1 6613
0 6615 7 1 2 6610 6614
0 6616 5 1 1 6615
0 6617 7 1 2 58238 6616
0 6618 5 1 1 6617
0 6619 7 1 2 46673 54110
0 6620 5 1 1 6619
0 6621 7 1 2 6618 6620
0 6622 5 1 1 6621
0 6623 7 1 2 40757 6622
0 6624 5 1 1 6623
0 6625 7 4 2 45629 49473
0 6626 5 3 1 58259
0 6627 7 8 2 48730 58263
0 6628 5 7 1 58266
0 6629 7 1 2 54760 55282
0 6630 7 1 2 58274 6629
0 6631 5 1 1 6630
0 6632 7 7 2 39974 45420
0 6633 5 2 1 58281
0 6634 7 2 2 58282 46902
0 6635 5 5 1 58290
0 6636 7 14 2 44024 46067
0 6637 5 1 1 58297
0 6638 7 1 2 58298 52791
0 6639 7 1 2 58291 6638
0 6640 5 1 1 6639
0 6641 7 1 2 6631 6640
0 6642 7 1 2 6624 6641
0 6643 7 1 2 6607 6642
0 6644 5 1 1 6643
0 6645 7 1 2 53870 52602
0 6646 7 1 2 6644 6645
0 6647 5 1 1 6646
0 6648 7 1 2 6597 6647
0 6649 5 1 1 6648
0 6650 7 1 2 55029 6649
0 6651 5 1 1 6650
0 6652 7 1 2 56254 54211
0 6653 5 1 1 6652
0 6654 7 1 2 41337 58152
0 6655 5 1 1 6654
0 6656 7 1 2 6653 6655
0 6657 7 1 2 55911 6656
0 6658 5 1 1 6657
0 6659 7 1 2 42510 6658
0 6660 5 1 1 6659
0 6661 7 2 2 41910 49690
0 6662 5 1 1 58311
0 6663 7 1 2 41197 6662
0 6664 5 2 1 6663
0 6665 7 2 2 52336 58313
0 6666 7 1 2 45848 54813
0 6667 7 1 2 58315 6666
0 6668 5 1 1 6667
0 6669 7 1 2 6660 6668
0 6670 5 1 1 6669
0 6671 7 1 2 42294 6670
0 6672 5 1 1 6671
0 6673 7 3 2 56255 54749
0 6674 5 2 1 58317
0 6675 7 1 2 49412 50534
0 6676 5 1 1 6675
0 6677 7 1 2 58320 6676
0 6678 5 1 1 6677
0 6679 7 1 2 52439 6678
0 6680 5 1 1 6679
0 6681 7 1 2 6672 6680
0 6682 5 1 1 6681
0 6683 7 1 2 46068 6682
0 6684 5 1 1 6683
0 6685 7 1 2 6417 6684
0 6686 5 1 1 6685
0 6687 7 1 2 44907 6686
0 6688 5 1 1 6687
0 6689 7 2 2 42511 52682
0 6690 5 1 1 58322
0 6691 7 3 2 43321 52667
0 6692 7 1 2 52174 58324
0 6693 5 1 1 6692
0 6694 7 1 2 6690 6693
0 6695 5 1 1 6694
0 6696 7 1 2 56088 50130
0 6697 7 1 2 6695 6696
0 6698 5 1 1 6697
0 6699 7 1 2 6688 6698
0 6700 5 1 1 6699
0 6701 7 1 2 44025 6700
0 6702 5 1 1 6701
0 6703 7 1 2 47626 58072
0 6704 5 1 1 6703
0 6705 7 2 2 51380 58119
0 6706 5 1 1 58327
0 6707 7 1 2 45630 6706
0 6708 5 1 1 6707
0 6709 7 1 2 6704 6708
0 6710 5 1 1 6709
0 6711 7 1 2 42512 6710
0 6712 5 1 1 6711
0 6713 7 1 2 52800 52480
0 6714 5 1 1 6713
0 6715 7 1 2 6712 6714
0 6716 5 1 1 6715
0 6717 7 1 2 46674 6716
0 6718 5 1 1 6717
0 6719 7 1 2 56528 54960
0 6720 5 1 1 6719
0 6721 7 1 2 6718 6720
0 6722 5 1 1 6721
0 6723 7 1 2 44026 6722
0 6724 5 1 1 6723
0 6725 7 1 2 55612 55603
0 6726 7 1 2 48418 6725
0 6727 5 1 1 6726
0 6728 7 1 2 6724 6727
0 6729 5 1 1 6728
0 6730 7 1 2 48731 6729
0 6731 5 1 1 6730
0 6732 7 4 2 47392 49413
0 6733 7 6 2 40758 45849
0 6734 7 2 2 56089 55604
0 6735 7 1 2 58333 58339
0 6736 7 1 2 58329 6735
0 6737 5 1 1 6736
0 6738 7 1 2 6731 6737
0 6739 7 1 2 6702 6738
0 6740 5 1 1 6739
0 6741 7 1 2 49352 6740
0 6742 5 1 1 6741
0 6743 7 3 2 52175 48335
0 6744 7 1 2 49414 51521
0 6745 7 2 2 58341 6744
0 6746 5 1 1 58344
0 6747 7 1 2 47627 58345
0 6748 5 1 1 6747
0 6749 7 1 2 40360 51080
0 6750 5 1 1 6749
0 6751 7 1 2 54731 6750
0 6752 5 1 1 6751
0 6753 7 2 2 42060 49547
0 6754 5 2 1 58346
0 6755 7 1 2 48387 58347
0 6756 5 1 1 6755
0 6757 7 1 2 52654 6756
0 6758 5 1 1 6757
0 6759 7 1 2 50166 6758
0 6760 5 1 1 6759
0 6761 7 1 2 42295 6760
0 6762 5 1 1 6761
0 6763 7 1 2 6752 6762
0 6764 5 1 1 6763
0 6765 7 1 2 49241 6764
0 6766 5 1 1 6765
0 6767 7 2 2 51884 52216
0 6768 5 1 1 58350
0 6769 7 1 2 54701 58351
0 6770 5 1 1 6769
0 6771 7 1 2 42296 55872
0 6772 7 1 2 54739 6771
0 6773 7 1 2 6770 6772
0 6774 5 1 1 6773
0 6775 7 4 2 46069 51522
0 6776 7 1 2 51709 6768
0 6777 5 3 1 6776
0 6778 7 1 2 47393 58356
0 6779 5 1 1 6778
0 6780 7 1 2 45631 800
0 6781 7 1 2 47572 6780
0 6782 7 1 2 6779 6781
0 6783 5 1 1 6782
0 6784 7 1 2 58352 6783
0 6785 7 1 2 6774 6784
0 6786 5 1 1 6785
0 6787 7 1 2 6766 6786
0 6788 5 1 1 6787
0 6789 7 1 2 42513 6788
0 6790 5 1 1 6789
0 6791 7 1 2 6748 6790
0 6792 5 1 1 6791
0 6793 7 1 2 49011 6792
0 6794 5 1 1 6793
0 6795 7 1 2 42514 55876
0 6796 5 2 1 6795
0 6797 7 2 2 51915 54036
0 6798 5 1 1 58361
0 6799 7 1 2 58359 6798
0 6800 5 1 1 6799
0 6801 7 1 2 44623 6800
0 6802 5 1 1 6801
0 6803 7 2 2 47394 50425
0 6804 5 1 1 58363
0 6805 7 1 2 50337 58364
0 6806 5 1 1 6805
0 6807 7 1 2 53677 6806
0 6808 5 1 1 6807
0 6809 7 1 2 42515 6808
0 6810 5 1 1 6809
0 6811 7 1 2 6802 6810
0 6812 5 1 1 6811
0 6813 7 1 2 47628 6812
0 6814 5 2 1 6813
0 6815 7 1 2 3849 55873
0 6816 5 1 1 6815
0 6817 7 1 2 42297 6816
0 6818 5 2 1 6817
0 6819 7 3 2 47081 49761
0 6820 5 3 1 58369
0 6821 7 1 2 48732 56310
0 6822 5 1 1 6821
0 6823 7 1 2 58372 6822
0 6824 5 1 1 6823
0 6825 7 1 2 45632 6824
0 6826 5 1 1 6825
0 6827 7 2 2 58367 6826
0 6828 5 1 1 58375
0 6829 7 1 2 42516 6828
0 6830 5 1 1 6829
0 6831 7 1 2 58365 6830
0 6832 5 1 1 6831
0 6833 7 2 2 56771 56424
0 6834 7 1 2 6832 58377
0 6835 5 1 1 6834
0 6836 7 1 2 43322 51135
0 6837 5 2 1 6836
0 6838 7 1 2 51136 47173
0 6839 5 1 1 6838
0 6840 7 4 2 58379 6839
0 6841 5 1 1 58381
0 6842 7 1 2 40182 47204
0 6843 5 2 1 6842
0 6844 7 1 2 6841 58385
0 6845 5 1 1 6844
0 6846 7 1 2 48873 6845
0 6847 5 1 1 6846
0 6848 7 3 2 42298 48733
0 6849 5 5 1 58387
0 6850 7 4 2 49474 58390
0 6851 5 1 1 58395
0 6852 7 1 2 58321 58396
0 6853 5 1 1 6852
0 6854 7 2 2 52412 50462
0 6855 5 2 1 58399
0 6856 7 1 2 52217 58401
0 6857 7 1 2 6853 6856
0 6858 7 1 2 6847 6857
0 6859 5 3 1 6858
0 6860 7 3 2 45850 49104
0 6861 7 1 2 52909 58406
0 6862 7 1 2 58403 6861
0 6863 5 1 1 6862
0 6864 7 1 2 6835 6863
0 6865 5 1 1 6864
0 6866 7 1 2 45024 6865
0 6867 5 1 1 6866
0 6868 7 1 2 50918 51100
0 6869 5 1 1 6868
0 6870 7 1 2 50369 54761
0 6871 7 1 2 6869 6870
0 6872 5 1 1 6871
0 6873 7 1 2 58235 6872
0 6874 5 1 1 6873
0 6875 7 1 2 54858 57007
0 6876 7 1 2 48960 6875
0 6877 7 1 2 6874 6876
0 6878 5 1 1 6877
0 6879 7 1 2 6867 6878
0 6880 7 1 2 6794 6879
0 6881 5 1 1 6880
0 6882 7 1 2 42946 6881
0 6883 5 1 1 6882
0 6884 7 1 2 6742 6883
0 6885 5 1 1 6884
0 6886 7 1 2 46607 6885
0 6887 5 1 1 6886
0 6888 7 1 2 6651 6887
0 6889 5 1 1 6888
0 6890 7 1 2 46350 6889
0 6891 5 1 1 6890
0 6892 7 11 2 43071 46608
0 6893 5 1 1 58409
0 6894 7 2 2 50322 52685
0 6895 7 1 2 55970 58420
0 6896 5 1 1 6895
0 6897 7 9 2 46070 49190
0 6898 7 1 2 41911 56201
0 6899 5 2 1 6898
0 6900 7 5 2 51262 58431
0 6901 5 5 1 58433
0 6902 7 1 2 47768 58434
0 6903 5 2 1 6902
0 6904 7 1 2 46792 58283
0 6905 5 6 1 6904
0 6906 7 2 2 42299 58445
0 6907 5 1 1 58451
0 6908 7 2 2 51381 6907
0 6909 5 3 1 58453
0 6910 7 1 2 41198 53150
0 6911 5 3 1 6910
0 6912 7 1 2 58458 54057
0 6913 7 1 2 58455 6912
0 6914 7 1 2 58443 6913
0 6915 5 2 1 6914
0 6916 7 1 2 58422 58461
0 6917 5 1 1 6916
0 6918 7 3 2 42784 58086
0 6919 7 2 2 48053 58463
0 6920 5 1 1 58466
0 6921 7 1 2 6917 6920
0 6922 5 1 1 6921
0 6923 7 1 2 49475 6922
0 6924 5 1 1 6923
0 6925 7 1 2 45633 47205
0 6926 5 1 1 6925
0 6927 7 1 2 58292 6926
0 6928 5 1 1 6927
0 6929 7 1 2 40183 6928
0 6930 5 1 1 6929
0 6931 7 1 2 48655 52542
0 6932 5 1 1 6931
0 6933 7 1 2 45634 58382
0 6934 5 1 1 6933
0 6935 7 1 2 6932 6934
0 6936 7 1 2 6930 6935
0 6937 5 2 1 6936
0 6938 7 1 2 58423 58468
0 6939 5 1 1 6938
0 6940 7 1 2 6924 6939
0 6941 5 1 1 6940
0 6942 7 1 2 45851 6941
0 6943 5 1 1 6942
0 6944 7 1 2 6896 6943
0 6945 5 1 1 6944
0 6946 7 1 2 49012 6945
0 6947 5 1 1 6946
0 6948 7 4 2 51199 50528
0 6949 5 2 1 58470
0 6950 7 1 2 50997 58471
0 6951 5 2 1 6950
0 6952 7 1 2 47547 58476
0 6953 5 2 1 6952
0 6954 7 1 2 49476 51799
0 6955 5 2 1 6954
0 6956 7 2 2 48734 58480
0 6957 5 1 1 58482
0 6958 7 1 2 45635 54905
0 6959 5 1 1 6958
0 6960 7 2 2 58483 6959
0 6961 5 1 1 58484
0 6962 7 1 2 58478 58485
0 6963 5 3 1 6962
0 6964 7 2 2 58407 58486
0 6965 5 1 1 58489
0 6966 7 1 2 47221 58490
0 6967 5 1 1 6966
0 6968 7 1 2 42300 52845
0 6969 5 2 1 6968
0 6970 7 1 2 51205 58491
0 6971 5 1 1 6970
0 6972 7 1 2 41912 6971
0 6973 5 1 1 6972
0 6974 7 1 2 53175 56394
0 6975 5 1 1 6974
0 6976 7 1 2 49477 6975
0 6977 7 1 2 6973 6976
0 6978 5 1 1 6977
0 6979 7 4 2 42785 51973
0 6980 5 1 1 58493
0 6981 7 1 2 45852 52543
0 6982 5 1 1 6981
0 6983 7 1 2 46675 6982
0 6984 5 1 1 6983
0 6985 7 1 2 6980 6984
0 6986 5 1 1 6985
0 6987 7 2 2 45853 49478
0 6988 5 2 1 58497
0 6989 7 1 2 58499 55170
0 6990 7 1 2 6986 6989
0 6991 7 1 2 6978 6990
0 6992 5 1 1 6991
0 6993 7 1 2 6967 6992
0 6994 5 1 1 6993
0 6995 7 1 2 41733 6994
0 6996 5 1 1 6995
0 6997 7 3 2 44027 57722
0 6998 5 1 1 58501
0 6999 7 4 2 58502 56166
0 7000 5 1 1 58504
0 7001 7 1 2 55188 55850
0 7002 5 1 1 7001
0 7003 7 1 2 7000 7002
0 7004 5 1 1 7003
0 7005 7 1 2 46071 7004
0 7006 5 1 1 7005
0 7007 7 1 2 56167 58378
0 7008 5 1 1 7007
0 7009 7 1 2 7006 7008
0 7010 5 1 1 7009
0 7011 7 1 2 41913 7010
0 7012 5 1 1 7011
0 7013 7 3 2 42061 56060
0 7014 7 1 2 58508 57399
0 7015 5 1 1 7014
0 7016 7 1 2 7012 7015
0 7017 5 1 1 7016
0 7018 7 1 2 47629 7017
0 7019 5 1 1 7018
0 7020 7 1 2 58432 54052
0 7021 5 1 1 7020
0 7022 7 1 2 57400 7021
0 7023 5 1 1 7022
0 7024 7 2 2 53137 51068
0 7025 7 1 2 44908 58511
0 7026 5 1 1 7025
0 7027 7 1 2 7023 7026
0 7028 5 1 1 7027
0 7029 7 1 2 51446 7028
0 7030 5 1 1 7029
0 7031 7 3 2 42062 48336
0 7032 7 3 2 40759 55728
0 7033 7 1 2 43515 51623
0 7034 7 1 2 58516 7033
0 7035 7 1 2 58513 7034
0 7036 5 1 1 7035
0 7037 7 1 2 7030 7036
0 7038 5 1 1 7037
0 7039 7 1 2 40934 7038
0 7040 5 1 1 7039
0 7041 7 2 2 53338 47947
0 7042 7 1 2 44177 55729
0 7043 7 1 2 58519 7042
0 7044 7 1 2 58514 7043
0 7045 5 1 1 7044
0 7046 7 1 2 7040 7045
0 7047 7 1 2 7019 7046
0 7048 5 1 1 7047
0 7049 7 1 2 48735 7048
0 7050 5 1 1 7049
0 7051 7 1 2 6996 7050
0 7052 7 1 2 6947 7051
0 7053 5 1 1 7052
0 7054 7 1 2 46226 7053
0 7055 5 1 1 7054
0 7056 7 3 2 42301 58095
0 7057 5 1 1 58521
0 7058 7 1 2 58080 58522
0 7059 5 1 1 7058
0 7060 7 1 2 49479 7059
0 7061 5 1 1 7060
0 7062 7 3 2 45636 51081
0 7063 5 3 1 58524
0 7064 7 1 2 47769 58525
0 7065 5 1 1 7064
0 7066 7 3 2 48736 7065
0 7067 5 1 1 58530
0 7068 7 1 2 58479 58531
0 7069 7 1 2 7061 7068
0 7070 5 2 1 7069
0 7071 7 2 2 40935 42947
0 7072 7 1 2 55407 58535
0 7073 7 1 2 48450 7072
0 7074 7 1 2 58533 7073
0 7075 5 1 1 7074
0 7076 7 1 2 7055 7075
0 7077 5 1 1 7076
0 7078 7 1 2 58410 7077
0 7079 5 1 1 7078
0 7080 7 1 2 6891 7079
0 7081 5 1 1 7080
0 7082 7 1 2 46559 7081
0 7083 5 1 1 7082
0 7084 7 21 2 41040 41826
0 7085 5 2 1 58537
0 7086 7 1 2 55417 58462
0 7087 5 1 1 7086
0 7088 7 18 2 42786 46351
0 7089 7 7 2 42517 58560
0 7090 7 2 2 50323 50910
0 7091 7 1 2 58578 58585
0 7092 5 1 1 7091
0 7093 7 1 2 7087 7092
0 7094 5 1 1 7093
0 7095 7 1 2 49191 7094
0 7096 5 1 1 7095
0 7097 7 5 2 45854 54597
0 7098 7 1 2 58587 58467
0 7099 5 1 1 7098
0 7100 7 1 2 7096 7099
0 7101 5 1 1 7100
0 7102 7 1 2 49013 7101
0 7103 5 1 1 7102
0 7104 7 4 2 44178 42787
0 7105 5 1 1 58592
0 7106 7 3 2 46227 58593
0 7107 7 2 2 45025 51523
0 7108 7 3 2 46352 7057
0 7109 7 1 2 58599 58601
0 7110 5 1 1 7109
0 7111 7 2 2 41734 56838
0 7112 7 1 2 48054 58604
0 7113 5 1 1 7112
0 7114 7 1 2 7110 7113
0 7115 5 1 1 7114
0 7116 7 1 2 58596 7115
0 7117 5 1 1 7116
0 7118 7 7 2 45421 42948
0 7119 7 2 2 56670 49370
0 7120 7 2 2 49853 58613
0 7121 7 1 2 58606 58615
0 7122 5 1 1 7121
0 7123 7 1 2 7117 7122
0 7124 5 1 1 7123
0 7125 7 1 2 39975 7124
0 7126 5 1 1 7125
0 7127 7 5 2 44028 56968
0 7128 7 1 2 58617 51507
0 7129 7 1 2 58602 7128
0 7130 5 1 1 7129
0 7131 7 1 2 7126 7130
0 7132 5 1 1 7131
0 7133 7 1 2 46736 7132
0 7134 5 1 1 7133
0 7135 7 1 2 45422 58108
0 7136 5 1 1 7135
0 7137 7 1 2 42302 7136
0 7138 5 1 1 7137
0 7139 7 5 2 40760 43072
0 7140 7 2 2 48103 57723
0 7141 5 1 1 58627
0 7142 7 1 2 44179 57530
0 7143 5 1 1 7142
0 7144 7 1 2 7141 7143
0 7145 5 4 1 7144
0 7146 7 1 2 58622 58629
0 7147 5 1 1 7146
0 7148 7 4 2 53631 48961
0 7149 5 1 1 58633
0 7150 7 1 2 58634 57022
0 7151 5 1 1 7150
0 7152 7 1 2 7147 7151
0 7153 5 1 1 7152
0 7154 7 1 2 7138 7153
0 7155 5 1 1 7154
0 7156 7 3 2 52092 46860
0 7157 7 3 2 47770 58637
0 7158 5 1 1 58640
0 7159 7 1 2 7158 1522
0 7160 5 1 1 7159
0 7161 7 1 2 58614 7160
0 7162 5 1 1 7161
0 7163 7 1 2 58561 57023
0 7164 7 1 2 58641 7163
0 7165 5 1 1 7164
0 7166 7 1 2 7162 7165
0 7167 5 1 1 7166
0 7168 7 1 2 57222 7167
0 7169 5 1 1 7168
0 7170 7 1 2 7155 7169
0 7171 5 1 1 7170
0 7172 7 1 2 41735 7171
0 7173 5 1 1 7172
0 7174 7 2 2 57325 56969
0 7175 7 1 2 45259 52763
0 7176 7 1 2 58643 7175
0 7177 7 1 2 58603 7176
0 7178 5 1 1 7177
0 7179 7 1 2 7173 7178
0 7180 7 1 2 7134 7179
0 7181 5 1 1 7180
0 7182 7 1 2 45855 7181
0 7183 5 1 1 7182
0 7184 7 1 2 7103 7183
0 7185 5 1 1 7184
0 7186 7 1 2 45069 7185
0 7187 5 1 1 7186
0 7188 7 3 2 52603 56671
0 7189 7 2 2 58087 58645
0 7190 7 4 2 41774 49362
0 7191 5 1 1 58650
0 7192 7 1 2 49105 58651
0 7193 7 1 2 58648 7192
0 7194 5 1 1 7193
0 7195 7 1 2 7187 7194
0 7196 5 1 1 7195
0 7197 7 1 2 44227 7196
0 7198 5 1 1 7197
0 7199 7 11 2 45026 45070
0 7200 7 12 2 44180 40976
0 7201 7 2 2 58654 58665
0 7202 7 1 2 48430 58677
0 7203 7 1 2 58649 7202
0 7204 5 1 1 7203
0 7205 7 1 2 7198 7204
0 7206 5 1 1 7205
0 7207 7 1 2 49480 7206
0 7208 5 1 1 7207
0 7209 7 9 2 44029 46353
0 7210 7 3 2 41914 47395
0 7211 5 4 1 58688
0 7212 7 1 2 41736 58689
0 7213 5 1 1 7212
0 7214 7 1 2 52876 7213
0 7215 7 1 2 1356 7214
0 7216 7 1 2 7067 7215
0 7217 5 1 1 7216
0 7218 7 1 2 58247 50003
0 7219 7 1 2 58474 7218
0 7220 5 1 1 7219
0 7221 7 1 2 7217 7220
0 7222 5 1 1 7221
0 7223 7 1 2 55230 7222
0 7224 5 1 1 7223
0 7225 7 1 2 41089 53123
0 7226 5 1 1 7225
0 7227 7 1 2 50015 7226
0 7228 5 1 1 7227
0 7229 7 1 2 39976 7228
0 7230 5 1 1 7229
0 7231 7 2 2 48368 46976
0 7232 5 1 1 58695
0 7233 7 1 2 7232 50004
0 7234 5 1 1 7233
0 7235 7 1 2 50158 49978
0 7236 5 1 1 7235
0 7237 7 1 2 7234 7236
0 7238 7 1 2 7230 7237
0 7239 5 1 1 7238
0 7240 7 1 2 44624 7239
0 7241 5 1 1 7240
0 7242 7 1 2 41737 52784
0 7243 5 3 1 7242
0 7244 7 1 2 41338 49979
0 7245 5 1 1 7244
0 7246 7 1 2 58697 7245
0 7247 5 1 1 7246
0 7248 7 1 2 47396 7247
0 7249 5 1 1 7248
0 7250 7 3 2 44625 49980
0 7251 5 1 1 58700
0 7252 7 1 2 47531 50306
0 7253 5 1 1 7252
0 7254 7 1 2 58701 7253
0 7255 5 1 1 7254
0 7256 7 1 2 42063 7255
0 7257 7 1 2 7249 7256
0 7258 5 1 1 7257
0 7259 7 4 2 46228 49879
0 7260 7 1 2 51624 58703
0 7261 5 1 1 7260
0 7262 7 1 2 47715 50005
0 7263 5 1 1 7262
0 7264 7 1 2 45423 7263
0 7265 7 1 2 7261 7264
0 7266 5 1 1 7265
0 7267 7 1 2 7258 7266
0 7268 5 1 1 7267
0 7269 7 1 2 42303 7268
0 7270 7 1 2 7241 7269
0 7271 5 1 1 7270
0 7272 7 1 2 58370 53129
0 7273 5 1 1 7272
0 7274 7 1 2 49415 53124
0 7275 5 1 1 7274
0 7276 7 1 2 45637 7275
0 7277 7 1 2 7273 7276
0 7278 5 1 1 7277
0 7279 7 1 2 42518 7278
0 7280 7 1 2 7271 7279
0 7281 5 1 1 7280
0 7282 7 5 2 47771 50844
0 7283 5 4 1 58707
0 7284 7 2 2 42064 58712
0 7285 5 1 1 58716
0 7286 7 1 2 46229 52883
0 7287 7 1 2 55854 7286
0 7288 7 1 2 58717 7287
0 7289 5 1 1 7288
0 7290 7 1 2 7281 7289
0 7291 5 1 1 7290
0 7292 7 1 2 46072 7291
0 7293 5 1 1 7292
0 7294 7 1 2 7224 7293
0 7295 5 1 1 7294
0 7296 7 1 2 44909 7295
0 7297 5 1 1 7296
0 7298 7 11 2 42519 42949
0 7299 7 2 2 55327 58718
0 7300 5 1 1 58729
0 7301 7 1 2 49416 58730
0 7302 5 1 1 7301
0 7303 7 3 2 52176 49981
0 7304 7 1 2 58330 58731
0 7305 5 1 1 7304
0 7306 7 1 2 40361 58702
0 7307 5 1 1 7306
0 7308 7 1 2 927 52808
0 7309 7 2 2 42950 50718
0 7310 5 1 1 58734
0 7311 7 1 2 50020 7310
0 7312 7 1 2 7308 7311
0 7313 5 1 1 7312
0 7314 7 1 2 7307 7313
0 7315 5 1 1 7314
0 7316 7 1 2 42520 7315
0 7317 5 1 1 7316
0 7318 7 1 2 7305 7317
0 7319 5 1 1 7318
0 7320 7 1 2 42304 7319
0 7321 5 1 1 7320
0 7322 7 1 2 7302 7321
0 7323 5 1 1 7322
0 7324 7 1 2 47222 7323
0 7325 5 1 1 7324
0 7326 7 1 2 7297 7325
0 7327 5 1 1 7326
0 7328 7 1 2 58679 7327
0 7329 5 1 1 7328
0 7330 7 2 2 55418 58469
0 7331 5 2 1 58736
0 7332 7 1 2 41738 49192
0 7333 7 1 2 58737 7332
0 7334 5 1 1 7333
0 7335 7 1 2 47548 58475
0 7336 5 1 1 7335
0 7337 7 1 2 58532 7336
0 7338 5 2 1 7337
0 7339 7 1 2 55231 58740
0 7340 5 1 1 7339
0 7341 7 8 2 43660 41915
0 7342 5 2 1 58742
0 7343 7 3 2 48811 52686
0 7344 7 1 2 58743 58752
0 7345 5 1 1 7344
0 7346 7 1 2 7340 7345
0 7347 5 1 1 7346
0 7348 7 1 2 57115 7347
0 7349 5 1 1 7348
0 7350 7 4 2 44398 42305
0 7351 5 3 1 58755
0 7352 7 4 2 43323 58756
0 7353 5 2 1 58762
0 7354 7 1 2 58732 58763
0 7355 5 1 1 7354
0 7356 7 1 2 7355 7300
0 7357 5 1 1 7356
0 7358 7 1 2 49417 7357
0 7359 5 1 1 7358
0 7360 7 7 2 42306 42951
0 7361 7 3 2 54425 58768
0 7362 7 1 2 53339 52809
0 7363 7 1 2 58775 7362
0 7364 5 1 1 7363
0 7365 7 1 2 7359 7364
0 7366 5 1 1 7365
0 7367 7 1 2 44910 58562
0 7368 7 1 2 7366 7367
0 7369 5 1 1 7368
0 7370 7 1 2 7349 7369
0 7371 5 1 1 7370
0 7372 7 1 2 40761 7371
0 7373 5 1 1 7372
0 7374 7 1 2 44181 7373
0 7375 7 1 2 7334 7374
0 7376 7 1 2 7329 7375
0 7377 5 1 1 7376
0 7378 7 1 2 50691 56216
0 7379 5 1 1 7378
0 7380 7 1 2 58068 7379
0 7381 5 1 1 7380
0 7382 7 1 2 57468 7381
0 7383 5 1 1 7382
0 7384 7 1 2 58738 7383
0 7385 5 1 1 7384
0 7386 7 1 2 41611 7385
0 7387 5 1 1 7386
0 7388 7 2 2 46354 52683
0 7389 7 7 2 44626 54528
0 7390 7 1 2 57752 58780
0 7391 7 1 2 58778 7390
0 7392 5 1 1 7391
0 7393 7 1 2 44030 7392
0 7394 7 1 2 7387 7393
0 7395 5 1 1 7394
0 7396 7 8 2 42521 48576
0 7397 7 6 2 42065 46355
0 7398 7 1 2 50324 58795
0 7399 7 1 2 52810 7398
0 7400 7 1 2 58787 7399
0 7401 5 1 1 7400
0 7402 7 1 2 58739 7401
0 7403 5 1 1 7402
0 7404 7 1 2 44911 7403
0 7405 5 1 1 7404
0 7406 7 2 2 54598 48337
0 7407 7 1 2 56083 58801
0 7408 5 1 1 7407
0 7409 7 3 2 45638 55815
0 7410 7 1 2 53666 58803
0 7411 5 1 1 7410
0 7412 7 1 2 7408 7411
0 7413 5 1 1 7412
0 7414 7 1 2 49418 7413
0 7415 5 1 1 7414
0 7416 7 1 2 40762 7415
0 7417 7 1 2 7405 7416
0 7418 5 1 1 7417
0 7419 7 1 2 45027 7418
0 7420 7 1 2 7395 7419
0 7421 5 1 1 7420
0 7422 7 3 2 40763 52604
0 7423 7 1 2 58806 58741
0 7424 5 1 1 7423
0 7425 7 4 2 43661 51034
0 7426 7 1 2 55885 56346
0 7427 7 1 2 58809 7426
0 7428 5 1 1 7427
0 7429 7 1 2 7424 7428
0 7430 5 1 1 7429
0 7431 7 1 2 56672 49854
0 7432 7 1 2 7430 7431
0 7433 5 1 1 7432
0 7434 7 1 2 40936 7433
0 7435 7 1 2 7421 7434
0 7436 5 1 1 7435
0 7437 7 1 2 7377 7436
0 7438 5 1 1 7437
0 7439 7 1 2 52801 58733
0 7440 5 1 1 7439
0 7441 7 1 2 56168 58735
0 7442 5 1 1 7441
0 7443 7 1 2 7440 7442
0 7444 5 1 1 7443
0 7445 7 1 2 49242 7444
0 7446 5 1 1 7445
0 7447 7 4 2 49762 46918
0 7448 5 3 1 58813
0 7449 7 2 2 46230 55605
0 7450 7 3 2 46073 52164
0 7451 7 1 2 44031 58822
0 7452 7 1 2 58820 7451
0 7453 7 1 2 58814 7452
0 7454 5 1 1 7453
0 7455 7 1 2 7446 7454
0 7456 5 1 1 7455
0 7457 7 1 2 42307 7456
0 7458 5 1 1 7457
0 7459 7 4 2 45639 53813
0 7460 7 4 2 51524 58825
0 7461 7 1 2 56311 53130
0 7462 5 1 1 7461
0 7463 7 2 2 47716 49982
0 7464 5 1 1 58833
0 7465 7 1 2 42066 58834
0 7466 5 1 1 7465
0 7467 7 1 2 7462 7466
0 7468 5 1 1 7467
0 7469 7 1 2 58829 7468
0 7470 5 1 1 7469
0 7471 7 1 2 7458 7470
0 7472 5 1 1 7471
0 7473 7 1 2 44182 7472
0 7474 5 1 1 7473
0 7475 7 3 2 42308 58719
0 7476 7 1 2 50719 48983
0 7477 7 1 2 58835 7476
0 7478 7 1 2 49243 7477
0 7479 5 1 1 7478
0 7480 7 1 2 7474 7479
0 7481 5 1 1 7480
0 7482 7 1 2 46356 7481
0 7483 5 1 1 7482
0 7484 7 2 2 43073 55189
0 7485 5 2 1 58838
0 7486 7 2 2 46231 58839
0 7487 7 1 2 58842 58512
0 7488 5 1 1 7487
0 7489 7 1 2 7483 7488
0 7490 5 1 1 7489
0 7491 7 1 2 48737 7490
0 7492 5 1 1 7491
0 7493 7 1 2 45071 7492
0 7494 7 1 2 7438 7493
0 7495 5 1 1 7494
0 7496 7 1 2 54048 6804
0 7497 5 2 1 7496
0 7498 7 2 2 58788 58844
0 7499 7 1 2 56460 58846
0 7500 5 1 1 7499
0 7501 7 2 2 51035 55569
0 7502 7 4 2 44183 44627
0 7503 7 2 2 52636 58850
0 7504 7 1 2 58848 58854
0 7505 5 1 1 7504
0 7506 7 1 2 54129 58630
0 7507 5 1 1 7506
0 7508 7 1 2 7505 7507
0 7509 5 1 1 7508
0 7510 7 1 2 47717 7509
0 7511 5 1 1 7510
0 7512 7 1 2 56498 58536
0 7513 5 1 1 7512
0 7514 7 8 2 41612 41916
0 7515 7 1 2 58856 58597
0 7516 5 1 1 7515
0 7517 7 1 2 7513 7516
0 7518 5 1 1 7517
0 7519 7 1 2 42522 58845
0 7520 7 1 2 7518 7519
0 7521 5 1 1 7520
0 7522 7 1 2 7511 7521
0 7523 5 1 1 7522
0 7524 7 1 2 45028 7523
0 7525 5 1 1 7524
0 7526 7 1 2 7500 7525
0 7527 5 1 1 7526
0 7528 7 1 2 44032 7527
0 7529 5 1 1 7528
0 7530 7 1 2 45029 51169
0 7531 7 5 2 43662 51525
0 7532 7 4 2 44184 52637
0 7533 7 1 2 58864 58869
0 7534 7 1 2 7530 7533
0 7535 5 1 1 7534
0 7536 7 2 2 49193 49014
0 7537 7 1 2 42952 58873
0 7538 5 1 1 7537
0 7539 7 1 2 44033 56457
0 7540 7 1 2 53125 7539
0 7541 5 1 1 7540
0 7542 7 1 2 7538 7541
0 7543 5 1 1 7542
0 7544 7 1 2 42788 7543
0 7545 5 1 1 7544
0 7546 7 1 2 48104 51625
0 7547 7 1 2 58503 7546
0 7548 5 1 1 7547
0 7549 7 1 2 7545 7548
0 7550 5 1 1 7549
0 7551 7 1 2 42523 56202
0 7552 7 1 2 7550 7551
0 7553 5 1 1 7552
0 7554 7 1 2 7535 7553
0 7555 5 1 1 7554
0 7556 7 1 2 49913 7555
0 7557 5 1 1 7556
0 7558 7 1 2 48431 49015
0 7559 7 1 2 58847 7558
0 7560 5 1 1 7559
0 7561 7 1 2 7557 7560
0 7562 7 1 2 7529 7561
0 7563 5 2 1 7562
0 7564 7 1 2 43074 58875
0 7565 5 1 1 7564
0 7566 7 1 2 41775 7565
0 7567 5 1 1 7566
0 7568 7 1 2 44228 7567
0 7569 7 1 2 7495 7568
0 7570 5 1 1 7569
0 7571 7 5 2 42789 48432
0 7572 5 1 1 58877
0 7573 7 2 2 56937 58878
0 7574 7 20 2 43075 55030
0 7575 5 4 1 58884
0 7576 7 1 2 52212 55705
0 7577 5 3 1 7576
0 7578 7 1 2 58885 58908
0 7579 5 1 1 7578
0 7580 7 9 2 46357 57620
0 7581 7 1 2 42067 58911
0 7582 7 1 2 54732 7581
0 7583 5 1 1 7582
0 7584 7 1 2 7579 7583
0 7585 5 1 1 7584
0 7586 7 1 2 58882 7585
0 7587 5 1 1 7586
0 7588 7 1 2 55570 58870
0 7589 5 1 1 7588
0 7590 7 3 2 40937 48577
0 7591 7 1 2 41613 58920
0 7592 5 1 1 7591
0 7593 7 1 2 7589 7592
0 7594 5 1 1 7593
0 7595 7 1 2 56203 7594
0 7596 5 1 1 7595
0 7597 7 6 2 40938 44399
0 7598 7 5 2 43324 58923
0 7599 7 1 2 58929 57753
0 7600 5 1 1 7599
0 7601 7 1 2 7596 7600
0 7602 5 1 1 7601
0 7603 7 1 2 45030 7602
0 7604 5 1 1 7603
0 7605 7 5 2 44185 44400
0 7606 7 6 2 43325 58934
0 7607 7 1 2 52755 58939
0 7608 5 1 1 7607
0 7609 7 1 2 7604 7608
0 7610 5 1 1 7609
0 7611 7 1 2 48738 7610
0 7612 5 1 1 7611
0 7613 7 2 2 43663 44912
0 7614 7 3 2 46074 58945
0 7615 5 1 1 58947
0 7616 7 1 2 982 7251
0 7617 5 1 1 7616
0 7618 7 1 2 58948 7617
0 7619 5 1 1 7618
0 7620 7 1 2 51508 54225
0 7621 5 1 1 7620
0 7622 7 1 2 7619 7621
0 7623 5 1 1 7622
0 7624 7 1 2 44186 7623
0 7625 5 1 1 7624
0 7626 7 2 2 45031 58628
0 7627 7 1 2 54037 58950
0 7628 5 1 1 7627
0 7629 7 1 2 45640 7628
0 7630 7 1 2 7625 7629
0 7631 7 1 2 7612 7630
0 7632 5 1 1 7631
0 7633 7 2 2 47397 46676
0 7634 5 1 1 58952
0 7635 7 1 2 7634 52747
0 7636 5 1 1 7635
0 7637 7 1 2 49016 7636
0 7638 5 1 1 7637
0 7639 7 3 2 41614 52759
0 7640 7 1 2 58930 58954
0 7641 5 1 1 7640
0 7642 7 1 2 7638 7641
0 7643 5 1 1 7642
0 7644 7 1 2 52785 7643
0 7645 5 1 1 7644
0 7646 7 6 2 45032 42068
0 7647 7 1 2 50143 58957
0 7648 7 1 2 58871 7647
0 7649 5 1 1 7648
0 7650 7 1 2 42309 7649
0 7651 7 1 2 7645 7650
0 7652 5 1 1 7651
0 7653 7 1 2 46358 7652
0 7654 7 1 2 7632 7653
0 7655 5 1 1 7654
0 7656 7 1 2 42310 50450
0 7657 5 4 1 7656
0 7658 7 3 2 41917 48739
0 7659 5 2 1 58967
0 7660 7 1 2 58963 58970
0 7661 5 3 1 7660
0 7662 7 1 2 57039 52952
0 7663 7 1 2 58972 7662
0 7664 5 1 1 7663
0 7665 7 1 2 7655 7664
0 7666 5 1 1 7665
0 7667 7 1 2 57621 7666
0 7668 5 1 1 7667
0 7669 7 1 2 56938 58909
0 7670 5 1 1 7669
0 7671 7 1 2 49353 58973
0 7672 5 1 1 7671
0 7673 7 1 2 7670 7672
0 7674 5 1 1 7673
0 7675 7 1 2 47223 7674
0 7676 5 1 1 7675
0 7677 7 1 2 58974 58951
0 7678 5 1 1 7677
0 7679 7 1 2 7676 7678
0 7680 5 1 1 7679
0 7681 7 1 2 58886 7680
0 7682 5 1 1 7681
0 7683 7 1 2 50845 48656
0 7684 5 2 1 7683
0 7685 7 4 2 42069 43076
0 7686 7 11 2 53871 57622
0 7687 5 1 1 58981
0 7688 7 1 2 58982 52953
0 7689 5 1 1 7688
0 7690 7 2 2 45033 55031
0 7691 7 1 2 58631 58992
0 7692 5 1 1 7691
0 7693 7 1 2 7689 7692
0 7694 5 1 1 7693
0 7695 7 1 2 58977 7694
0 7696 5 1 1 7695
0 7697 7 2 2 58655 51269
0 7698 7 13 2 44187 44229
0 7699 7 1 2 58996 57855
0 7700 7 1 2 52661 7699
0 7701 7 1 2 58994 7700
0 7702 5 1 1 7701
0 7703 7 1 2 7696 7702
0 7704 5 1 1 7703
0 7705 7 1 2 58975 7704
0 7706 5 1 1 7705
0 7707 7 1 2 7682 7706
0 7708 7 1 2 7668 7707
0 7709 5 1 1 7708
0 7710 7 1 2 44034 7709
0 7711 5 1 1 7710
0 7712 7 1 2 7587 7711
0 7713 5 1 1 7712
0 7714 7 1 2 42524 7713
0 7715 5 1 1 7714
0 7716 7 1 2 45072 55190
0 7717 5 2 1 7716
0 7718 7 1 2 55025 59009
0 7719 5 1 1 7718
0 7720 7 7 2 57008 49363
0 7721 5 1 1 59011
0 7722 7 1 2 55032 7721
0 7723 5 1 1 7722
0 7724 7 4 2 7719 7723
0 7725 7 1 2 43077 50040
0 7726 7 1 2 59018 7725
0 7727 5 1 1 7726
0 7728 7 4 2 43664 44230
0 7729 7 2 2 51526 59022
0 7730 7 4 2 54069 58851
0 7731 5 1 1 59028
0 7732 7 5 2 45073 45856
0 7733 7 1 2 59029 59032
0 7734 7 1 2 59026 7733
0 7735 5 1 1 7734
0 7736 7 1 2 7727 7735
0 7737 5 1 1 7736
0 7738 7 1 2 48323 7737
0 7739 5 1 1 7738
0 7740 7 2 2 43665 56939
0 7741 7 21 2 45074 46359
0 7742 5 2 1 59039
0 7743 7 7 2 44035 44231
0 7744 7 3 2 59040 59062
0 7745 7 1 2 44628 51726
0 7746 7 1 2 59069 7745
0 7747 7 1 2 59037 7746
0 7748 5 1 1 7747
0 7749 7 1 2 7739 7748
0 7750 5 1 1 7749
0 7751 7 1 2 46075 7750
0 7752 5 1 1 7751
0 7753 7 3 2 49161 56656
0 7754 5 1 1 59072
0 7755 7 3 2 45857 57623
0 7756 7 5 2 40939 44629
0 7757 7 1 2 43666 45034
0 7758 7 1 2 59078 7757
0 7759 7 1 2 59075 7758
0 7760 7 1 2 59073 7759
0 7761 5 1 1 7760
0 7762 7 1 2 7752 7761
0 7763 5 1 1 7762
0 7764 7 1 2 51036 7763
0 7765 5 1 1 7764
0 7766 7 1 2 7715 7765
0 7767 5 1 1 7766
0 7768 7 1 2 47630 7767
0 7769 5 1 1 7768
0 7770 7 4 2 45075 43078
0 7771 7 8 2 40977 59083
0 7772 5 3 1 59087
0 7773 7 1 2 59088 58876
0 7774 5 1 1 7773
0 7775 7 5 2 42525 55171
0 7776 5 1 1 59098
0 7777 7 1 2 3291 54555
0 7778 5 2 1 7777
0 7779 7 2 2 48740 59103
0 7780 5 1 1 59105
0 7781 7 1 2 50581 56633
0 7782 5 1 1 7781
0 7783 7 2 2 7780 7782
0 7784 5 1 1 59107
0 7785 7 1 2 47718 7784
0 7786 5 1 1 7785
0 7787 7 1 2 53410 54546
0 7788 5 1 1 7787
0 7789 7 2 2 46360 51287
0 7790 7 1 2 59109 58958
0 7791 5 1 1 7790
0 7792 7 1 2 54692 7791
0 7793 5 1 1 7792
0 7794 7 1 2 47398 7793
0 7795 5 1 1 7794
0 7796 7 1 2 7788 7795
0 7797 7 1 2 7786 7796
0 7798 5 1 1 7797
0 7799 7 1 2 51601 7798
0 7800 5 1 1 7799
0 7801 7 1 2 49419 54547
0 7802 5 1 1 7801
0 7803 7 1 2 46950 56634
0 7804 5 1 1 7803
0 7805 7 1 2 54693 7804
0 7806 5 1 1 7805
0 7807 7 1 2 58764 7806
0 7808 5 1 1 7807
0 7809 7 1 2 7802 7808
0 7810 7 1 2 7800 7809
0 7811 5 1 1 7810
0 7812 7 1 2 59099 7811
0 7813 5 1 1 7812
0 7814 7 2 2 53632 49106
0 7815 7 1 2 52165 59111
0 7816 7 1 2 58404 7815
0 7817 5 1 1 7816
0 7818 7 1 2 7813 7817
0 7819 5 1 1 7818
0 7820 7 1 2 57624 7819
0 7821 5 1 1 7820
0 7822 7 1 2 59100 52050
0 7823 5 1 1 7822
0 7824 7 1 2 6965 7823
0 7825 5 1 1 7824
0 7826 7 1 2 54979 58993
0 7827 7 1 2 7825 7826
0 7828 5 1 1 7827
0 7829 7 1 2 7821 7828
0 7830 5 1 1 7829
0 7831 7 1 2 52910 7830
0 7832 5 1 1 7831
0 7833 7 1 2 7774 7832
0 7834 7 1 2 7769 7833
0 7835 7 1 2 7570 7834
0 7836 7 1 2 7208 7835
0 7837 5 1 1 7836
0 7838 7 1 2 58538 7837
0 7839 5 1 1 7838
0 7840 7 1 2 7083 7839
0 7841 5 1 1 7840
0 7842 7 1 2 46455 7841
0 7843 5 1 1 7842
0 7844 7 11 2 44036 40978
0 7845 7 3 2 41776 59113
0 7846 7 2 2 54599 52911
0 7847 7 2 2 42526 59127
0 7848 7 2 2 59129 58357
0 7849 7 1 2 59124 59131
0 7850 5 1 1 7849
0 7851 7 16 2 46361 55033
0 7852 7 7 2 46076 48055
0 7853 7 2 2 41918 51832
0 7854 7 3 2 58720 59156
0 7855 7 1 2 59149 59158
0 7856 5 1 1 7855
0 7857 7 1 2 49244 59157
0 7858 5 1 1 7857
0 7859 7 3 2 58299 55606
0 7860 7 1 2 59161 51827
0 7861 5 1 1 7860
0 7862 7 1 2 7858 7861
0 7863 5 1 1 7862
0 7864 7 1 2 42527 7863
0 7865 5 1 1 7864
0 7866 7 1 2 6746 7865
0 7867 5 1 1 7866
0 7868 7 1 2 46232 7867
0 7869 5 1 1 7868
0 7870 7 1 2 7856 7869
0 7871 5 1 1 7870
0 7872 7 1 2 47631 7871
0 7873 5 1 1 7872
0 7874 7 1 2 53699 46677
0 7875 5 1 1 7874
0 7876 7 1 2 56086 7875
0 7877 5 1 1 7876
0 7878 7 1 2 49880 7877
0 7879 5 1 1 7878
0 7880 7 1 2 42311 54808
0 7881 7 1 2 52655 7880
0 7882 5 1 1 7881
0 7883 7 1 2 58124 7882
0 7884 5 2 1 7883
0 7885 7 1 2 46678 59164
0 7886 5 1 1 7885
0 7887 7 1 2 7879 7886
0 7888 5 1 1 7887
0 7889 7 1 2 42528 7888
0 7890 5 1 1 7889
0 7891 7 2 2 49936 52573
0 7892 5 1 1 59166
0 7893 7 1 2 53115 59167
0 7894 5 1 1 7893
0 7895 7 1 2 7890 7894
0 7896 5 1 1 7895
0 7897 7 1 2 44037 7896
0 7898 5 1 1 7897
0 7899 7 1 2 49881 55535
0 7900 5 1 1 7899
0 7901 7 3 2 45858 49823
0 7902 5 1 1 59168
0 7903 7 1 2 42312 59169
0 7904 5 1 1 7903
0 7905 7 1 2 7900 7904
0 7906 5 1 1 7905
0 7907 7 2 2 50692 7906
0 7908 7 1 2 58879 59171
0 7909 5 1 1 7908
0 7910 7 1 2 7898 7909
0 7911 5 1 1 7910
0 7912 7 1 2 46233 7911
0 7913 5 1 1 7912
0 7914 7 1 2 48137 59172
0 7915 5 1 1 7914
0 7916 7 1 2 7913 7915
0 7917 7 1 2 7873 7916
0 7918 5 1 1 7917
0 7919 7 1 2 59133 7918
0 7920 5 1 1 7919
0 7921 7 1 2 7850 7920
0 7922 5 1 1 7921
0 7923 7 1 2 41739 7922
0 7924 5 1 1 7923
0 7925 7 1 2 47632 54115
0 7926 5 2 1 7925
0 7927 7 1 2 51796 59173
0 7928 5 1 1 7927
0 7929 7 1 2 42529 51062
0 7930 7 1 2 7928 7929
0 7931 5 1 1 7930
0 7932 7 1 2 7892 7931
0 7933 5 1 1 7932
0 7934 7 7 2 41777 48578
0 7935 7 7 2 40979 45035
0 7936 7 1 2 59182 58680
0 7937 7 1 2 58857 7936
0 7938 7 1 2 59175 7937
0 7939 7 1 2 7933 7938
0 7940 5 1 1 7939
0 7941 7 1 2 7924 7940
0 7942 5 1 1 7941
0 7943 7 1 2 40940 7942
0 7944 5 1 1 7943
0 7945 7 1 2 44630 52440
0 7946 5 2 1 7945
0 7947 7 3 2 43667 55536
0 7948 5 1 1 59191
0 7949 7 1 2 59189 7948
0 7950 5 4 1 7949
0 7951 7 1 2 47633 59194
0 7952 5 1 1 7951
0 7953 7 3 2 41339 50325
0 7954 5 1 1 59198
0 7955 7 1 2 42530 59199
0 7956 5 1 1 7955
0 7957 7 1 2 7952 7956
0 7958 5 1 1 7957
0 7959 7 1 2 42070 7958
0 7960 5 1 1 7959
0 7961 7 1 2 51602 54058
0 7962 7 1 2 51833 7961
0 7963 5 1 1 7962
0 7964 7 1 2 1543 7963
0 7965 5 1 1 7964
0 7966 7 1 2 42531 7965
0 7967 5 1 1 7966
0 7968 7 1 2 7960 7967
0 7969 5 1 1 7968
0 7970 7 8 2 45036 41778
0 7971 7 3 2 44188 59201
0 7972 5 1 1 59209
0 7973 7 1 2 44913 59114
0 7974 7 2 2 59210 7973
0 7975 7 1 2 56571 59212
0 7976 7 1 2 7969 7975
0 7977 5 1 1 7976
0 7978 7 1 2 7944 7977
0 7979 5 1 1 7978
0 7980 7 1 2 46560 7979
0 7981 5 1 1 7980
0 7982 7 8 2 41740 45076
0 7983 7 4 2 40941 59214
0 7984 5 1 1 59222
0 7985 7 2 2 59223 59063
0 7986 7 1 2 59226 59132
0 7987 5 1 1 7986
0 7988 7 2 2 53814 56329
0 7989 7 1 2 56970 59228
0 7990 5 1 1 7989
0 7991 7 2 2 42953 56090
0 7992 7 2 2 40942 44487
0 7993 7 2 2 59230 59232
0 7994 7 1 2 41919 56000
0 7995 7 1 2 59234 7994
0 7996 5 1 1 7995
0 7997 7 1 2 7990 7996
0 7998 5 1 1 7997
0 7999 7 1 2 52722 7998
0 8000 5 1 1 7999
0 8001 7 1 2 56416 58872
0 8002 5 1 1 8001
0 8003 7 1 2 54777 55730
0 8004 7 1 2 58921 8003
0 8005 5 1 1 8004
0 8006 7 1 2 8002 8005
0 8007 5 1 1 8006
0 8008 7 1 2 42532 8007
0 8009 5 1 1 8008
0 8010 7 1 2 8000 8009
0 8011 5 1 1 8010
0 8012 7 1 2 48741 8011
0 8013 5 1 1 8012
0 8014 7 2 2 54929 51727
0 8015 7 4 2 44631 46077
0 8016 7 4 2 43668 44189
0 8017 7 1 2 59238 59242
0 8018 7 1 2 59236 8017
0 8019 5 1 1 8018
0 8020 7 2 2 42954 55816
0 8021 7 1 2 41920 50795
0 8022 7 1 2 59233 8021
0 8023 7 1 2 59246 8022
0 8024 5 1 1 8023
0 8025 7 1 2 8019 8024
0 8026 5 1 1 8025
0 8027 7 1 2 43516 8026
0 8028 5 1 1 8027
0 8029 7 1 2 254 7954
0 8030 5 1 1 8029
0 8031 7 4 2 44914 53815
0 8032 5 1 1 59248
0 8033 7 1 2 59249 56134
0 8034 7 1 2 8030 8033
0 8035 5 1 1 8034
0 8036 7 1 2 8028 8035
0 8037 5 1 1 8036
0 8038 7 1 2 42071 8037
0 8039 5 1 1 8038
0 8040 7 1 2 56099 59235
0 8041 5 1 1 8040
0 8042 7 1 2 43669 53243
0 8043 7 1 2 58855 8042
0 8044 5 1 1 8043
0 8045 7 1 2 8041 8044
0 8046 5 1 1 8045
0 8047 7 1 2 42533 8046
0 8048 5 1 1 8047
0 8049 7 7 2 44190 44488
0 8050 7 1 2 52649 59252
0 8051 5 1 1 8050
0 8052 7 1 2 58858 58922
0 8053 5 1 1 8052
0 8054 7 1 2 8051 8053
0 8055 5 1 1 8054
0 8056 7 4 2 43517 45641
0 8057 7 3 2 44632 59259
0 8058 5 2 1 59263
0 8059 7 1 2 59266 4529
0 8060 5 1 1 8059
0 8061 7 1 2 42534 8060
0 8062 5 1 1 8061
0 8063 7 1 2 44633 58362
0 8064 5 1 1 8063
0 8065 7 1 2 8062 8064
0 8066 5 1 1 8065
0 8067 7 1 2 8055 8066
0 8068 5 1 1 8067
0 8069 7 1 2 8048 8068
0 8070 7 1 2 8039 8069
0 8071 7 1 2 8013 8070
0 8072 5 1 1 8071
0 8073 7 1 2 59070 8072
0 8074 5 1 1 8073
0 8075 7 1 2 44038 58632
0 8076 5 1 1 8075
0 8077 7 1 2 49107 48264
0 8078 5 1 1 8077
0 8079 7 1 2 8076 8078
0 8080 5 1 1 8079
0 8081 7 1 2 42535 58887
0 8082 7 1 2 58358 8081
0 8083 7 1 2 8080 8082
0 8084 5 1 1 8083
0 8085 7 1 2 8074 8084
0 8086 5 1 1 8085
0 8087 7 1 2 45037 8086
0 8088 5 1 1 8087
0 8089 7 1 2 7987 8088
0 8090 5 1 1 8089
0 8091 7 1 2 58539 8090
0 8092 5 1 1 8091
0 8093 7 1 2 7981 8092
0 8094 5 1 1 8093
0 8095 7 1 2 46456 8094
0 8096 5 1 1 8095
0 8097 7 8 2 44915 41779
0 8098 7 2 2 49937 58586
0 8099 7 1 2 59268 59276
0 8100 5 1 1 8099
0 8101 7 3 2 45077 57231
0 8102 7 1 2 50297 59278
0 8103 5 1 1 8102
0 8104 7 1 2 8100 8103
0 8105 5 1 1 8104
0 8106 7 1 2 40980 8105
0 8107 5 1 1 8106
0 8108 7 2 2 44232 56330
0 8109 7 6 2 41780 45424
0 8110 7 1 2 59283 58077
0 8111 7 1 2 59281 8110
0 8112 5 1 1 8111
0 8113 7 1 2 8107 8112
0 8114 5 1 1 8113
0 8115 7 1 2 44039 8114
0 8116 5 1 1 8115
0 8117 7 8 2 46234 55034
0 8118 7 1 2 48433 50298
0 8119 7 1 2 59289 8118
0 8120 5 1 1 8119
0 8121 7 1 2 8116 8120
0 8122 5 1 1 8121
0 8123 7 1 2 46561 8122
0 8124 5 1 1 8123
0 8125 7 8 2 45078 41827
0 8126 5 1 1 59297
0 8127 7 6 2 44233 59298
0 8128 5 1 1 59305
0 8129 7 5 2 41041 44916
0 8130 7 2 2 44040 59311
0 8131 7 2 2 59306 59316
0 8132 7 1 2 59318 59277
0 8133 5 1 1 8132
0 8134 7 1 2 8124 8133
0 8135 5 1 1 8134
0 8136 7 1 2 57737 8135
0 8137 5 1 1 8136
0 8138 7 5 2 44489 44917
0 8139 7 6 2 43670 45260
0 8140 7 1 2 51332 59325
0 8141 7 1 2 59320 8140
0 8142 7 7 2 43169 58540
0 8143 5 1 1 59331
0 8144 7 2 2 42955 46609
0 8145 7 1 2 59264 59338
0 8146 7 1 2 59332 8145
0 8147 7 1 2 8141 8146
0 8148 5 1 1 8147
0 8149 7 1 2 45859 8148
0 8150 7 1 2 8137 8149
0 8151 5 1 1 8150
0 8152 7 7 2 46457 46562
0 8153 7 5 2 45079 48056
0 8154 7 2 2 46078 59347
0 8155 7 1 2 58704 59352
0 8156 5 1 1 8155
0 8157 7 1 2 50693 49194
0 8158 7 1 2 59176 8157
0 8159 5 1 1 8158
0 8160 7 1 2 8156 8159
0 8161 5 1 1 8160
0 8162 7 1 2 44634 8161
0 8163 5 1 1 8162
0 8164 7 4 2 43671 48057
0 8165 7 10 2 45080 46235
0 8166 7 1 2 47719 59358
0 8167 7 1 2 59354 8166
0 8168 5 1 1 8167
0 8169 7 4 2 41781 51527
0 8170 7 1 2 50054 59368
0 8171 7 1 2 51790 8170
0 8172 5 1 1 8171
0 8173 7 1 2 8168 8172
0 8174 5 1 1 8173
0 8175 7 1 2 46079 8174
0 8176 5 1 1 8175
0 8177 7 1 2 8163 8176
0 8178 5 1 1 8177
0 8179 7 1 2 45642 8178
0 8180 5 1 1 8179
0 8181 7 1 2 45425 51603
0 8182 5 1 1 8181
0 8183 7 1 2 42072 53380
0 8184 5 1 1 8183
0 8185 7 1 2 8182 8184
0 8186 5 1 1 8185
0 8187 7 1 2 54930 59353
0 8188 7 1 2 8186 8187
0 8189 5 1 1 8188
0 8190 7 1 2 8180 8189
0 8191 5 1 1 8190
0 8192 7 1 2 59340 8191
0 8193 5 1 1 8192
0 8194 7 4 2 42956 52912
0 8195 7 4 2 44041 41828
0 8196 7 2 2 41782 42313
0 8197 7 2 2 41042 43170
0 8198 7 1 2 59380 59382
0 8199 7 1 2 59376 8198
0 8200 7 1 2 59372 8199
0 8201 5 1 1 8200
0 8202 7 1 2 8193 8201
0 8203 5 1 1 8202
0 8204 7 1 2 40981 8203
0 8205 5 1 1 8204
0 8206 7 7 2 44234 46458
0 8207 7 10 2 46236 48058
0 8208 7 1 2 41783 46563
0 8209 7 2 2 59391 8208
0 8210 7 1 2 53700 59401
0 8211 5 1 1 8210
0 8212 7 1 2 59299 50055
0 8213 7 1 2 59312 8212
0 8214 7 1 2 54304 8213
0 8215 5 1 1 8214
0 8216 7 1 2 8211 8215
0 8217 5 1 1 8216
0 8218 7 1 2 49882 8217
0 8219 5 1 1 8218
0 8220 7 1 2 59165 59402
0 8221 5 1 1 8220
0 8222 7 1 2 8219 8221
0 8223 5 1 1 8222
0 8224 7 1 2 46080 8223
0 8225 5 1 1 8224
0 8226 7 3 2 45643 55886
0 8227 7 3 2 45081 42073
0 8228 7 1 2 59406 58541
0 8229 7 1 2 59403 8228
0 8230 7 1 2 51638 8229
0 8231 5 1 1 8230
0 8232 7 1 2 8225 8231
0 8233 5 1 1 8232
0 8234 7 1 2 59384 8233
0 8235 5 1 1 8234
0 8236 7 1 2 42536 8235
0 8237 7 1 2 8205 8236
0 8238 5 1 1 8237
0 8239 7 1 2 46362 8238
0 8240 7 1 2 8151 8239
0 8241 5 1 1 8240
0 8242 7 4 2 59269 59115
0 8243 7 1 2 59409 59159
0 8244 5 1 1 8243
0 8245 7 2 2 40764 54220
0 8246 7 1 2 59290 59413
0 8247 7 1 2 59195 8246
0 8248 5 1 1 8247
0 8249 7 1 2 8244 8248
0 8250 5 1 1 8249
0 8251 7 1 2 46564 8250
0 8252 5 1 1 8251
0 8253 7 1 2 59160 59319
0 8254 5 1 1 8253
0 8255 7 1 2 8252 8254
0 8256 5 1 1 8255
0 8257 7 1 2 56782 8256
0 8258 5 1 1 8257
0 8259 7 3 2 55035 49195
0 8260 7 14 2 42537 43079
0 8261 7 2 2 59418 58542
0 8262 7 1 2 50056 47955
0 8263 7 1 2 59432 8262
0 8264 7 1 2 59415 8263
0 8265 5 1 1 8264
0 8266 7 1 2 8258 8265
0 8267 5 1 1 8266
0 8268 7 1 2 46459 8267
0 8269 5 1 1 8268
0 8270 7 3 2 40765 54600
0 8271 7 2 2 49081 59434
0 8272 5 1 1 59437
0 8273 7 1 2 58681 59373
0 8274 5 1 1 8273
0 8275 7 1 2 8272 8274
0 8276 5 1 1 8275
0 8277 7 55 2 43171 46610
0 8278 5 4 1 59439
0 8279 7 2 2 59440 58543
0 8280 5 1 1 59498
0 8281 7 1 2 54426 59499
0 8282 7 1 2 8276 8281
0 8283 5 1 1 8282
0 8284 7 1 2 8269 8283
0 8285 5 1 1 8284
0 8286 7 1 2 47634 8285
0 8287 5 1 1 8286
0 8288 7 1 2 49911 50415
0 8289 5 2 1 8288
0 8290 7 12 2 42790 46460
0 8291 7 1 2 59502 50057
0 8292 7 1 2 59416 8291
0 8293 7 1 2 59500 8292
0 8294 5 1 1 8293
0 8295 7 7 2 43172 59392
0 8296 7 5 2 40982 59381
0 8297 7 1 2 46081 59521
0 8298 7 1 2 59514 8297
0 8299 5 1 1 8298
0 8300 7 1 2 8294 8299
0 8301 5 1 1 8300
0 8302 7 1 2 59433 8301
0 8303 5 1 1 8302
0 8304 7 1 2 8287 8303
0 8305 7 1 2 8241 8304
0 8306 5 1 1 8305
0 8307 7 1 2 49017 8306
0 8308 5 1 1 8307
0 8309 7 1 2 8096 8308
0 8310 5 1 1 8309
0 8311 7 1 2 47319 8310
0 8312 5 1 1 8311
0 8313 7 23 2 45140 46461
0 8314 5 1 1 59526
0 8315 7 1 2 59527 53740
0 8316 5 1 1 8315
0 8317 7 2 2 42074 48742
0 8318 5 2 1 59549
0 8319 7 4 2 58391 59551
0 8320 7 1 2 51207 59553
0 8321 5 3 1 8320
0 8322 7 2 2 43173 59557
0 8323 7 1 2 41829 59560
0 8324 5 1 1 8323
0 8325 7 1 2 8316 8324
0 8326 5 1 1 8325
0 8327 7 1 2 41043 8326
0 8328 5 1 1 8327
0 8329 7 3 2 46462 46554
0 8330 7 1 2 53741 59562
0 8331 5 1 1 8330
0 8332 7 1 2 8328 8331
0 8333 5 1 1 8332
0 8334 7 1 2 49245 8333
0 8335 5 1 1 8334
0 8336 7 3 2 41830 51528
0 8337 7 1 2 41044 46082
0 8338 7 1 2 59565 8337
0 8339 7 1 2 59561 8338
0 8340 5 1 1 8339
0 8341 7 1 2 8335 8340
0 8342 5 1 1 8341
0 8343 7 1 2 42538 8342
0 8344 5 1 1 8343
0 8345 7 6 2 41831 45644
0 8346 7 2 2 41045 59568
0 8347 7 1 2 49420 56204
0 8348 5 2 1 8347
0 8349 7 2 2 43174 59576
0 8350 7 1 2 59574 59578
0 8351 5 1 1 8350
0 8352 7 2 2 48743 49706
0 8353 5 1 1 59580
0 8354 7 3 2 50998 59581
0 8355 7 1 2 40184 54900
0 8356 5 1 1 8355
0 8357 7 1 2 59582 8356
0 8358 5 1 1 8357
0 8359 7 1 2 45645 8358
0 8360 5 1 1 8359
0 8361 7 1 2 47007 52986
0 8362 5 2 1 8361
0 8363 7 1 2 40362 48015
0 8364 5 1 1 8363
0 8365 7 1 2 59585 8364
0 8366 7 1 2 8360 8365
0 8367 5 1 1 8366
0 8368 7 1 2 59341 8367
0 8369 5 1 1 8368
0 8370 7 1 2 8351 8369
0 8371 5 1 1 8370
0 8372 7 1 2 51529 8371
0 8373 5 1 1 8372
0 8374 7 1 2 51572 59342
0 8375 7 1 2 56360 8374
0 8376 5 1 1 8375
0 8377 7 1 2 8373 8376
0 8378 5 1 1 8377
0 8379 7 1 2 48088 55232
0 8380 7 1 2 8378 8379
0 8381 5 1 1 8380
0 8382 7 1 2 8344 8381
0 8383 5 1 1 8382
0 8384 7 1 2 46611 8383
0 8385 5 1 1 8384
0 8386 7 1 2 42539 53742
0 8387 5 1 1 8386
0 8388 7 1 2 45860 56361
0 8389 5 1 1 8388
0 8390 7 2 2 8387 8389
0 8391 5 1 1 59587
0 8392 7 1 2 51573 59588
0 8393 5 1 1 8392
0 8394 7 2 2 44042 58203
0 8395 5 1 1 59589
0 8396 7 1 2 45861 59590
0 8397 5 2 1 8396
0 8398 7 1 2 49172 59591
0 8399 5 1 1 8398
0 8400 7 5 2 44235 41046
0 8401 7 2 2 41832 42791
0 8402 7 2 2 46463 59598
0 8403 7 2 2 59593 59600
0 8404 7 1 2 45082 59602
0 8405 7 1 2 8399 8404
0 8406 7 1 2 8393 8405
0 8407 5 1 1 8406
0 8408 7 1 2 8385 8407
0 8409 5 1 1 8408
0 8410 7 1 2 54578 8409
0 8411 5 1 1 8410
0 8412 7 8 2 40766 56772
0 8413 7 1 2 46555 59604
0 8414 5 1 1 8413
0 8415 7 3 2 45141 48059
0 8416 7 2 2 40943 41047
0 8417 7 1 2 59612 59615
0 8418 5 1 1 8417
0 8419 7 1 2 8414 8418
0 8420 5 1 1 8419
0 8421 7 1 2 58563 8420
0 8422 7 1 2 58205 8421
0 8423 5 1 1 8422
0 8424 7 1 2 58353 52298
0 8425 5 1 1 8424
0 8426 7 1 2 44043 52913
0 8427 5 1 1 8426
0 8428 7 1 2 49345 8427
0 8429 5 9 1 8428
0 8430 7 1 2 43672 59617
0 8431 5 1 1 8430
0 8432 7 1 2 58354 53403
0 8433 5 1 1 8432
0 8434 7 1 2 8431 8433
0 8435 5 1 1 8434
0 8436 7 1 2 52021 8435
0 8437 5 1 1 8436
0 8438 7 1 2 42314 59618
0 8439 5 1 1 8438
0 8440 7 1 2 41921 59162
0 8441 5 1 1 8440
0 8442 7 1 2 8439 8441
0 8443 5 1 1 8442
0 8444 7 1 2 44635 8443
0 8445 5 1 1 8444
0 8446 7 1 2 8437 8445
0 8447 7 1 2 8425 8446
0 8448 5 1 1 8447
0 8449 7 1 2 42540 8448
0 8450 5 1 1 8449
0 8451 7 2 2 54469 58487
0 8452 5 1 1 59626
0 8453 7 1 2 48962 59627
0 8454 5 1 1 8453
0 8455 7 1 2 8450 8454
0 8456 5 1 1 8455
0 8457 7 8 2 41833 43080
0 8458 7 3 2 44191 41048
0 8459 7 1 2 59628 59636
0 8460 7 1 2 8456 8459
0 8461 5 1 1 8460
0 8462 7 1 2 8423 8461
0 8463 5 1 1 8462
0 8464 7 1 2 46464 8463
0 8465 5 1 1 8464
0 8466 7 1 2 47772 58454
0 8467 5 4 1 8466
0 8468 7 1 2 56205 58255
0 8469 5 3 1 8468
0 8470 7 1 2 45646 59643
0 8471 5 1 1 8470
0 8472 7 1 2 51755 8471
0 8473 5 1 1 8472
0 8474 7 1 2 58964 8473
0 8475 5 1 1 8474
0 8476 7 1 2 59639 8475
0 8477 5 1 1 8476
0 8478 7 1 2 49196 8477
0 8479 5 1 1 8478
0 8480 7 6 2 45261 50476
0 8481 5 1 1 59646
0 8482 7 2 2 49550 59647
0 8483 5 1 1 59652
0 8484 7 1 2 41615 59653
0 8485 5 1 1 8484
0 8486 7 1 2 8479 8485
0 8487 5 1 1 8486
0 8488 7 1 2 45862 8487
0 8489 5 1 1 8488
0 8490 7 1 2 40767 59558
0 8491 5 1 1 8490
0 8492 7 11 2 41090 55667
0 8493 5 4 1 59654
0 8494 7 4 2 59655 52585
0 8495 5 2 1 59669
0 8496 7 1 2 48022 59670
0 8497 5 1 1 8496
0 8498 7 1 2 8491 8497
0 8499 5 1 1 8498
0 8500 7 1 2 51974 8499
0 8501 5 1 1 8500
0 8502 7 1 2 8489 8501
0 8503 5 1 1 8502
0 8504 7 1 2 46083 8503
0 8505 5 1 1 8504
0 8506 7 2 2 53450 59577
0 8507 7 1 2 55273 59675
0 8508 5 1 1 8507
0 8509 7 1 2 8505 8508
0 8510 5 1 1 8509
0 8511 7 44 2 41834 43175
0 8512 5 3 1 59677
0 8513 7 1 2 46363 59678
0 8514 7 1 2 59616 8513
0 8515 7 1 2 8510 8514
0 8516 5 1 1 8515
0 8517 7 1 2 8465 8516
0 8518 5 1 1 8517
0 8519 7 1 2 55036 8518
0 8520 5 1 1 8519
0 8521 7 1 2 59679 50983
0 8522 7 1 2 58424 8521
0 8523 5 1 1 8522
0 8524 7 1 2 40185 48060
0 8525 7 7 2 41199 45142
0 8526 7 1 2 59724 59503
0 8527 7 1 2 8524 8526
0 8528 5 1 1 8527
0 8529 7 1 2 8523 8528
0 8530 5 1 1 8529
0 8531 7 1 2 45647 8530
0 8532 5 1 1 8531
0 8533 7 1 2 59528 6957
0 8534 5 1 1 8533
0 8535 7 4 2 45426 46465
0 8536 7 2 2 45143 59731
0 8537 5 1 1 59735
0 8538 7 1 2 59721 8537
0 8539 5 1 1 8538
0 8540 7 1 2 47773 8539
0 8541 5 1 1 8540
0 8542 7 1 2 59722 8314
0 8543 5 8 1 8542
0 8544 7 1 2 49481 59737
0 8545 5 1 1 8544
0 8546 7 1 2 8541 8545
0 8547 5 1 1 8546
0 8548 7 1 2 45648 8547
0 8549 5 1 1 8548
0 8550 7 1 2 8534 8549
0 8551 5 1 1 8550
0 8552 7 1 2 55274 8551
0 8553 5 1 1 8552
0 8554 7 1 2 8532 8553
0 8555 5 1 1 8554
0 8556 7 1 2 41049 8555
0 8557 5 1 1 8556
0 8558 7 8 2 46084 43176
0 8559 7 3 2 45649 59745
0 8560 7 1 2 41835 59313
0 8561 7 1 2 59753 8560
0 8562 5 1 1 8561
0 8563 7 1 2 47224 59343
0 8564 7 1 2 58477 8563
0 8565 5 1 1 8564
0 8566 7 1 2 8562 8565
0 8567 5 1 1 8566
0 8568 7 1 2 40768 8567
0 8569 5 1 1 8568
0 8570 7 2 2 45650 49082
0 8571 7 1 2 44044 59333
0 8572 7 1 2 59756 8571
0 8573 5 1 1 8572
0 8574 7 1 2 8569 8573
0 8575 5 1 1 8574
0 8576 7 1 2 47549 8575
0 8577 5 1 1 8576
0 8578 7 2 2 40769 44306
0 8579 7 2 2 41616 59758
0 8580 7 1 2 59760 59601
0 8581 7 1 2 6961 8580
0 8582 5 1 1 8581
0 8583 7 1 2 8577 8582
0 8584 7 1 2 8557 8583
0 8585 5 1 1 8584
0 8586 7 1 2 46612 8585
0 8587 5 1 1 8586
0 8588 7 1 2 59348 59603
0 8589 7 1 2 58488 8588
0 8590 5 1 1 8589
0 8591 7 1 2 8587 8590
0 8592 5 1 1 8591
0 8593 7 1 2 45863 8592
0 8594 5 1 1 8593
0 8595 7 1 2 46647 58558
0 8596 5 1 1 8595
0 8597 7 1 2 57669 46557
0 8598 5 1 1 8597
0 8599 7 4 2 8596 8598
0 8600 7 1 2 56916 59150
0 8601 7 1 2 59762 8600
0 8602 7 1 2 53415 8601
0 8603 5 1 1 8602
0 8604 7 1 2 8594 8603
0 8605 5 1 1 8604
0 8606 7 1 2 57026 8605
0 8607 5 1 1 8606
0 8608 7 1 2 8520 8607
0 8609 7 1 2 8411 8608
0 8610 5 1 1 8609
0 8611 7 1 2 52877 8610
0 8612 5 1 1 8611
0 8613 7 1 2 44045 51821
0 8614 5 1 1 8613
0 8615 7 2 2 47720 50919
0 8616 5 1 1 59766
0 8617 7 1 2 47399 59767
0 8618 5 1 1 8617
0 8619 7 1 2 8614 8618
0 8620 5 2 1 8619
0 8621 7 1 2 42075 59768
0 8622 5 1 1 8621
0 8623 7 2 2 44046 48744
0 8624 5 1 1 59770
0 8625 7 1 2 41617 8624
0 8626 7 1 2 8622 8625
0 8627 5 1 1 8626
0 8628 7 2 2 47550 58099
0 8629 5 1 1 59772
0 8630 7 6 2 42315 48657
0 8631 7 1 2 59773 59774
0 8632 5 1 1 8631
0 8633 7 1 2 40770 55701
0 8634 5 1 1 8633
0 8635 7 1 2 44918 8634
0 8636 7 1 2 8632 8635
0 8637 5 1 1 8636
0 8638 7 1 2 56169 8637
0 8639 7 1 2 8627 8638
0 8640 5 1 1 8639
0 8641 7 1 2 53451 57463
0 8642 7 1 2 47551 8641
0 8643 5 1 1 8642
0 8644 7 1 2 42792 8643
0 8645 7 1 2 8640 8644
0 8646 5 1 1 8645
0 8647 7 6 2 50451 47552
0 8648 7 1 2 59780 47563
0 8649 5 1 1 8648
0 8650 7 2 2 41200 41922
0 8651 7 3 2 59786 55576
0 8652 5 1 1 59788
0 8653 7 1 2 8649 8652
0 8654 5 2 1 8653
0 8655 7 1 2 59791 59775
0 8656 5 1 1 8655
0 8657 7 1 2 47635 53411
0 8658 5 1 1 8657
0 8659 7 1 2 59554 8658
0 8660 7 1 2 7285 8659
0 8661 5 1 1 8660
0 8662 7 1 2 40771 8661
0 8663 5 1 1 8662
0 8664 7 1 2 8656 8663
0 8665 5 2 1 8664
0 8666 7 1 2 50639 59793
0 8667 5 1 1 8666
0 8668 7 2 2 41923 59769
0 8669 5 1 1 59795
0 8670 7 1 2 44047 51604
0 8671 5 1 1 8670
0 8672 7 1 2 8669 8671
0 8673 5 1 1 8672
0 8674 7 1 2 42076 8673
0 8675 5 1 1 8674
0 8676 7 3 2 47579 48658
0 8677 5 3 1 59797
0 8678 7 2 2 44048 42316
0 8679 7 1 2 59800 59803
0 8680 5 1 1 8679
0 8681 7 1 2 8675 8680
0 8682 5 2 1 8681
0 8683 7 1 2 49855 59805
0 8684 5 1 1 8683
0 8685 7 1 2 8667 8684
0 8686 5 1 1 8685
0 8687 7 1 2 42541 8686
0 8688 5 1 1 8687
0 8689 7 1 2 58081 51756
0 8690 5 1 1 8689
0 8691 7 1 2 53230 49197
0 8692 7 2 2 8690 8691
0 8693 5 1 1 59807
0 8694 7 1 2 45038 59808
0 8695 5 1 1 8694
0 8696 7 1 2 46085 8695
0 8697 7 1 2 8688 8696
0 8698 5 1 1 8697
0 8699 7 1 2 8646 8698
0 8700 5 1 1 8699
0 8701 7 1 2 40944 8700
0 8702 5 1 1 8701
0 8703 7 1 2 51975 59794
0 8704 5 1 1 8703
0 8705 7 1 2 8693 8704
0 8706 5 1 1 8705
0 8707 7 1 2 56430 8706
0 8708 5 1 1 8707
0 8709 7 1 2 44192 8708
0 8710 5 1 1 8709
0 8711 7 1 2 43081 8710
0 8712 7 1 2 8702 8711
0 8713 5 1 1 8712
0 8714 7 1 2 48659 55844
0 8715 5 1 1 8714
0 8716 7 1 2 47636 8715
0 8717 5 1 1 8716
0 8718 7 1 2 49482 58766
0 8719 7 1 2 8717 8718
0 8720 5 3 1 8719
0 8721 7 1 2 54488 59809
0 8722 5 1 1 8721
0 8723 7 2 2 45864 59552
0 8724 5 1 1 59812
0 8725 7 1 2 50043 51761
0 8726 5 1 1 8725
0 8727 7 1 2 49921 8726
0 8728 5 1 1 8727
0 8729 7 2 2 59813 8728
0 8730 7 1 2 44049 59814
0 8731 5 1 1 8730
0 8732 7 1 2 8722 8731
0 8733 5 1 1 8732
0 8734 7 6 2 45039 58564
0 8735 7 1 2 56971 59816
0 8736 7 1 2 8733 8735
0 8737 5 1 1 8736
0 8738 7 1 2 46237 8737
0 8739 7 1 2 8713 8738
0 8740 5 1 1 8739
0 8741 7 4 2 47460 52321
0 8742 5 2 1 59822
0 8743 7 1 2 44050 53231
0 8744 5 2 1 8743
0 8745 7 1 2 51037 52592
0 8746 5 1 1 8745
0 8747 7 1 2 59828 8746
0 8748 5 1 1 8747
0 8749 7 1 2 59823 8748
0 8750 5 1 1 8749
0 8751 7 2 2 44051 53452
0 8752 5 2 1 59830
0 8753 7 1 2 53596 59776
0 8754 7 1 2 58100 8753
0 8755 5 1 1 8754
0 8756 7 1 2 59832 8755
0 8757 5 1 1 8756
0 8758 7 1 2 47272 8757
0 8759 5 1 1 8758
0 8760 7 2 2 48786 50999
0 8761 5 1 1 59834
0 8762 7 1 2 55759 50506
0 8763 5 1 1 8762
0 8764 7 1 2 59835 8763
0 8765 5 1 1 8764
0 8766 7 1 2 54470 8765
0 8767 5 1 1 8766
0 8768 7 1 2 8759 8767
0 8769 7 1 2 8750 8768
0 8770 5 1 1 8769
0 8771 7 1 2 42793 8770
0 8772 5 1 1 8771
0 8773 7 1 2 55810 59771
0 8774 5 1 1 8773
0 8775 7 1 2 8772 8774
0 8776 5 1 1 8775
0 8777 7 1 2 49018 8776
0 8778 5 1 1 8777
0 8779 7 1 2 47580 58965
0 8780 5 1 1 8779
0 8781 7 1 2 51966 51000
0 8782 5 1 1 8781
0 8783 7 1 2 45262 8782
0 8784 5 1 1 8783
0 8785 7 1 2 8780 8784
0 8786 7 1 2 59640 8785
0 8787 5 2 1 8786
0 8788 7 1 2 58823 59836
0 8789 5 1 1 8788
0 8790 7 1 2 42542 50694
0 8791 7 1 2 50072 8790
0 8792 7 1 2 51822 8791
0 8793 5 1 1 8792
0 8794 7 1 2 8789 8793
0 8795 5 1 1 8794
0 8796 7 1 2 49108 8795
0 8797 5 1 1 8796
0 8798 7 1 2 8778 8797
0 8799 5 1 1 8798
0 8800 7 1 2 44919 8799
0 8801 5 1 1 8800
0 8802 7 2 2 40772 55233
0 8803 5 1 1 59838
0 8804 7 1 2 51123 59839
0 8805 5 1 1 8804
0 8806 7 2 2 40186 48660
0 8807 5 2 1 59840
0 8808 7 1 2 55811 56539
0 8809 7 1 2 59841 8808
0 8810 5 1 1 8809
0 8811 7 1 2 8805 8810
0 8812 5 1 1 8811
0 8813 7 1 2 45427 8812
0 8814 5 1 1 8813
0 8815 7 1 2 58334 56192
0 8816 5 1 1 8815
0 8817 7 1 2 8814 8816
0 8818 5 1 1 8817
0 8819 7 1 2 47461 8818
0 8820 5 1 1 8819
0 8821 7 2 2 44490 47320
0 8822 5 5 1 59844
0 8823 7 1 2 45651 59846
0 8824 5 1 1 8823
0 8825 7 1 2 53101 8824
0 8826 5 1 1 8825
0 8827 7 1 2 55234 8826
0 8828 5 1 1 8827
0 8829 7 1 2 53816 58968
0 8830 5 1 1 8829
0 8831 7 1 2 8828 8830
0 8832 5 1 1 8831
0 8833 7 1 2 40773 8832
0 8834 5 1 1 8833
0 8835 7 1 2 8820 8834
0 8836 5 1 1 8835
0 8837 7 1 2 57523 8836
0 8838 5 1 1 8837
0 8839 7 1 2 8801 8838
0 8840 5 1 1 8839
0 8841 7 1 2 46364 8840
0 8842 5 1 1 8841
0 8843 7 4 2 53817 50672
0 8844 7 1 2 59851 51710
0 8845 5 1 1 8844
0 8846 7 1 2 4162 55266
0 8847 5 4 1 8846
0 8848 7 2 2 47008 59855
0 8849 7 1 2 40187 59859
0 8850 5 1 1 8849
0 8851 7 1 2 8845 8850
0 8852 5 1 1 8851
0 8853 7 1 2 58248 8852
0 8854 5 1 1 8853
0 8855 7 1 2 59852 51082
0 8856 7 1 2 58708 8855
0 8857 5 1 1 8856
0 8858 7 1 2 8854 8857
0 8859 5 1 1 8858
0 8860 7 1 2 40363 8859
0 8861 5 1 1 8860
0 8862 7 2 2 40774 56066
0 8863 7 1 2 53377 59861
0 8864 5 1 1 8863
0 8865 7 3 2 45263 50276
0 8866 7 5 2 47581 47273
0 8867 5 4 1 59866
0 8868 7 1 2 56008 59867
0 8869 7 1 2 59863 8868
0 8870 5 1 1 8869
0 8871 7 1 2 8864 8870
0 8872 7 1 2 8861 8871
0 8873 5 1 1 8872
0 8874 7 1 2 56779 8873
0 8875 5 1 1 8874
0 8876 7 1 2 42957 8875
0 8877 7 1 2 8842 8876
0 8878 5 1 1 8877
0 8879 7 1 2 41784 8878
0 8880 7 1 2 8740 8879
0 8881 5 1 1 8880
0 8882 7 2 2 41741 59798
0 8883 7 2 2 53597 58769
0 8884 7 1 2 59875 59877
0 8885 5 1 1 8884
0 8886 7 1 2 52166 56347
0 8887 7 1 2 51762 8886
0 8888 5 1 1 8887
0 8889 7 1 2 8885 8888
0 8890 5 1 1 8889
0 8891 7 1 2 46086 8890
0 8892 5 1 1 8891
0 8893 7 1 2 42958 54859
0 8894 7 1 2 51323 8893
0 8895 7 1 2 51124 8894
0 8896 5 1 1 8895
0 8897 7 1 2 8892 8896
0 8898 5 1 1 8897
0 8899 7 1 2 45428 8898
0 8900 5 1 1 8899
0 8901 7 3 2 46238 47774
0 8902 7 1 2 45040 59879
0 8903 5 1 1 8902
0 8904 7 1 2 58698 8903
0 8905 5 1 1 8904
0 8906 7 1 2 56067 58335
0 8907 7 1 2 8905 8906
0 8908 5 1 1 8907
0 8909 7 1 2 8900 8908
0 8910 5 1 1 8909
0 8911 7 1 2 47462 8910
0 8912 5 1 1 8911
0 8913 7 4 2 44052 45429
0 8914 5 1 1 59882
0 8915 7 2 2 46087 49483
0 8916 7 1 2 59883 59886
0 8917 5 1 1 8916
0 8918 7 1 2 42317 50379
0 8919 5 4 1 8918
0 8920 7 1 2 42077 56187
0 8921 5 1 1 8920
0 8922 7 1 2 51324 8921
0 8923 7 1 2 59888 8922
0 8924 5 1 1 8923
0 8925 7 1 2 8917 8924
0 8926 5 1 1 8925
0 8927 7 1 2 49983 8926
0 8928 5 1 1 8927
0 8929 7 1 2 53311 51509
0 8930 5 1 1 8929
0 8931 7 1 2 8928 8930
0 8932 5 1 1 8931
0 8933 7 1 2 47775 8932
0 8934 5 1 1 8933
0 8935 7 2 2 46239 51298
0 8936 7 3 2 41340 55772
0 8937 7 1 2 59892 59894
0 8938 5 1 1 8937
0 8939 7 1 2 56331 52779
0 8940 5 1 1 8939
0 8941 7 1 2 45430 51763
0 8942 5 1 1 8941
0 8943 7 1 2 51967 8942
0 8944 5 1 1 8943
0 8945 7 1 2 51633 52878
0 8946 7 1 2 8944 8945
0 8947 5 1 1 8946
0 8948 7 1 2 8940 8947
0 8949 5 1 1 8948
0 8950 7 1 2 51325 8949
0 8951 5 1 1 8950
0 8952 7 1 2 8938 8951
0 8953 7 1 2 8934 8952
0 8954 5 1 1 8953
0 8955 7 1 2 45865 8954
0 8956 5 1 1 8955
0 8957 7 2 2 41742 50058
0 8958 5 1 1 59897
0 8959 7 1 2 48661 58153
0 8960 5 1 1 8959
0 8961 7 1 2 59898 8960
0 8962 5 1 1 8961
0 8963 7 1 2 49984 59810
0 8964 5 1 1 8963
0 8965 7 1 2 8962 8964
0 8966 5 1 1 8965
0 8967 7 1 2 46088 54489
0 8968 7 1 2 8966 8967
0 8969 5 1 1 8968
0 8970 7 1 2 8956 8969
0 8971 7 1 2 8912 8970
0 8972 5 1 1 8971
0 8973 7 2 2 46365 8972
0 8974 7 1 2 40945 56579
0 8975 7 1 2 59899 8974
0 8976 5 1 1 8975
0 8977 7 1 2 8881 8976
0 8978 5 1 1 8977
0 8979 7 1 2 40983 8978
0 8980 5 1 1 8979
0 8981 7 2 2 51852 48779
0 8982 5 1 1 59901
0 8983 7 1 2 48745 8982
0 8984 5 1 1 8983
0 8985 7 1 2 49484 3336
0 8986 7 1 2 8984 8985
0 8987 5 1 1 8986
0 8988 7 1 2 59101 8987
0 8989 5 1 1 8988
0 8990 7 1 2 56194 58230
0 8991 5 1 1 8990
0 8992 7 3 2 40188 48780
0 8993 5 2 1 59903
0 8994 7 1 2 59906 58267
0 8995 7 1 2 8991 8994
0 8996 7 1 2 51885 51968
0 8997 5 1 1 8996
0 8998 7 1 2 45264 8997
0 8999 5 1 1 8998
0 9000 7 1 2 50995 58817
0 9001 5 1 1 9000
0 9002 7 1 2 8999 9001
0 9003 7 1 2 8995 9002
0 9004 7 1 2 59641 9003
0 9005 5 1 1 9004
0 9006 7 1 2 58408 9005
0 9007 5 1 1 9006
0 9008 7 1 2 8989 9007
0 9009 5 1 1 9008
0 9010 7 1 2 41743 9009
0 9011 5 1 1 9010
0 9012 7 1 2 40775 48984
0 9013 7 1 2 59815 9012
0 9014 5 1 1 9013
0 9015 7 1 2 9011 9014
0 9016 5 1 1 9015
0 9017 7 1 2 55037 9016
0 9018 5 1 1 9017
0 9019 7 7 2 41785 42543
0 9020 7 2 2 57009 59908
0 9021 7 1 2 59183 59915
0 9022 7 1 2 59811 9021
0 9023 5 1 1 9022
0 9024 7 1 2 9018 9023
0 9025 5 1 1 9024
0 9026 7 1 2 46366 9025
0 9027 5 1 1 9026
0 9028 7 4 2 43673 47931
0 9029 5 1 1 59917
0 9030 7 1 2 55484 59918
0 9031 5 2 1 9030
0 9032 7 3 2 45866 55328
0 9033 7 1 2 58411 49109
0 9034 7 1 2 59923 9033
0 9035 7 1 2 59921 9034
0 9036 5 1 1 9035
0 9037 7 1 2 9027 9036
0 9038 5 1 1 9037
0 9039 7 1 2 46240 9038
0 9040 5 1 1 9039
0 9041 7 1 2 49110 59676
0 9042 5 1 1 9041
0 9043 7 1 2 56364 59806
0 9044 5 1 1 9043
0 9045 7 1 2 9042 9044
0 9046 5 1 1 9045
0 9047 7 1 2 45041 9046
0 9048 5 1 1 9047
0 9049 7 1 2 54427 48976
0 9050 7 1 2 59796 9049
0 9051 5 1 1 9050
0 9052 7 1 2 9048 9051
0 9053 5 1 1 9052
0 9054 7 1 2 53633 46613
0 9055 7 1 2 9053 9054
0 9056 5 1 1 9055
0 9057 7 1 2 9040 9056
0 9058 5 1 1 9057
0 9059 7 1 2 52914 9058
0 9060 5 1 1 9059
0 9061 7 8 2 41924 43082
0 9062 7 6 2 41786 42959
0 9063 7 2 2 59926 59934
0 9064 7 1 2 59940 53162
0 9065 5 1 1 9064
0 9066 7 1 2 51605 53126
0 9067 5 1 1 9066
0 9068 7 1 2 58526 9067
0 9069 5 1 1 9068
0 9070 7 1 2 59041 53131
0 9071 7 1 2 9069 9070
0 9072 5 1 1 9071
0 9073 7 1 2 9065 9072
0 9074 5 1 1 9073
0 9075 7 1 2 54490 9074
0 9076 5 1 1 9075
0 9077 7 3 2 43083 59284
0 9078 5 1 1 59942
0 9079 7 1 2 45867 59943
0 9080 7 2 2 58066 9079
0 9081 7 1 2 7464 8958
0 9082 5 1 1 9081
0 9083 7 1 2 47637 9082
0 9084 7 1 2 59945 9083
0 9085 5 1 1 9084
0 9086 7 1 2 9076 9085
0 9087 5 1 1 9086
0 9088 7 1 2 41618 9087
0 9089 5 1 1 9088
0 9090 7 20 2 41787 43084
0 9091 5 6 1 59947
0 9092 7 6 2 41925 46367
0 9093 7 5 2 45083 59973
0 9094 5 1 1 59979
0 9095 7 1 2 59967 9094
0 9096 5 1 1 9095
0 9097 7 1 2 58527 9096
0 9098 5 1 1 9097
0 9099 7 2 2 59042 51606
0 9100 5 1 1 59984
0 9101 7 1 2 41926 59985
0 9102 5 1 1 9101
0 9103 7 1 2 9098 9102
0 9104 5 1 1 9103
0 9105 7 1 2 57425 56170
0 9106 7 1 2 9104 9105
0 9107 5 1 1 9106
0 9108 7 1 2 9089 9107
0 9109 5 1 1 9108
0 9110 7 1 2 40984 9109
0 9111 5 1 1 9110
0 9112 7 10 2 40776 48399
0 9113 5 4 1 59986
0 9114 7 2 2 41744 58528
0 9115 7 1 2 59987 60000
0 9116 5 1 1 9115
0 9117 7 1 2 51843 52213
0 9118 5 5 1 9117
0 9119 7 1 2 48324 57465
0 9120 7 1 2 60002 9119
0 9121 5 1 1 9120
0 9122 7 1 2 9116 9121
0 9123 5 1 1 9122
0 9124 7 3 2 46368 59909
0 9125 7 1 2 44236 60007
0 9126 7 1 2 9123 9125
0 9127 5 1 1 9126
0 9128 7 1 2 9111 9127
0 9129 5 1 1 9128
0 9130 7 1 2 46089 9129
0 9131 5 1 1 9130
0 9132 7 1 2 44053 59134
0 9133 7 1 2 60003 9132
0 9134 5 1 1 9133
0 9135 7 1 2 40777 802
0 9136 5 1 1 9135
0 9137 7 5 2 41788 42078
0 9138 7 3 2 40985 60010
0 9139 7 1 2 43085 60015
0 9140 7 1 2 9136 9139
0 9141 5 1 1 9140
0 9142 7 1 2 9134 9141
0 9143 5 1 1 9142
0 9144 7 1 2 41619 9143
0 9145 5 1 1 9144
0 9146 7 2 2 41789 58978
0 9147 7 6 2 40986 44920
0 9148 7 4 2 40778 60020
0 9149 7 1 2 60018 60026
0 9150 5 1 1 9149
0 9151 7 1 2 9145 9150
0 9152 5 1 1 9151
0 9153 7 1 2 53340 57541
0 9154 7 1 2 9152 9153
0 9155 5 1 1 9154
0 9156 7 1 2 9131 9155
0 9157 5 1 1 9156
0 9158 7 1 2 40946 9157
0 9159 5 1 1 9158
0 9160 7 1 2 59619 53127
0 9161 7 1 2 60004 9160
0 9162 5 1 1 9161
0 9163 7 1 2 48579 48434
0 9164 7 1 2 60001 9163
0 9165 5 1 1 9164
0 9166 7 1 2 9162 9165
0 9167 5 1 1 9166
0 9168 7 1 2 58666 60008
0 9169 7 1 2 9167 9168
0 9170 5 1 1 9169
0 9171 7 1 2 9159 9170
0 9172 5 1 1 9171
0 9173 7 1 2 47321 9172
0 9174 5 1 1 9173
0 9175 7 4 2 41091 47776
0 9176 5 2 1 60030
0 9177 7 2 2 52554 60034
0 9178 7 4 2 47638 60036
0 9179 7 1 2 53132 59946
0 9180 5 1 1 9179
0 9181 7 1 2 40779 53598
0 9182 7 1 2 53634 59215
0 9183 7 1 2 9181 9182
0 9184 5 1 1 9183
0 9185 7 1 2 9180 9184
0 9186 5 1 1 9185
0 9187 7 1 2 41620 9186
0 9188 5 1 1 9187
0 9189 7 4 2 58682 52132
0 9190 7 1 2 50059 59202
0 9191 5 1 1 9190
0 9192 7 7 2 42079 46241
0 9193 7 1 2 60046 59216
0 9194 5 1 1 9193
0 9195 7 1 2 9191 9194
0 9196 5 1 1 9195
0 9197 7 1 2 60042 9196
0 9198 5 1 1 9197
0 9199 7 1 2 9188 9198
0 9200 5 1 1 9199
0 9201 7 1 2 40987 9200
0 9202 5 1 1 9201
0 9203 7 1 2 51530 60047
0 9204 5 1 1 9203
0 9205 7 3 2 40780 58859
0 9206 7 1 2 42960 60053
0 9207 5 1 1 9206
0 9208 7 1 2 9204 9207
0 9209 5 1 1 9208
0 9210 7 5 2 44237 41745
0 9211 7 1 2 60056 60009
0 9212 7 1 2 9209 9211
0 9213 5 1 1 9212
0 9214 7 1 2 9202 9213
0 9215 5 1 1 9214
0 9216 7 1 2 46090 9215
0 9217 5 1 1 9216
0 9218 7 1 2 49162 53163
0 9219 7 1 2 55198 9218
0 9220 7 1 2 59135 9219
0 9221 5 1 1 9220
0 9222 7 1 2 9217 9221
0 9223 5 1 1 9222
0 9224 7 1 2 40947 9223
0 9225 5 1 1 9224
0 9226 7 2 2 53818 53635
0 9227 7 2 2 41790 41927
0 9228 7 2 2 58667 60063
0 9229 7 1 2 60061 60065
0 9230 7 1 2 57466 9229
0 9231 5 1 1 9230
0 9232 7 1 2 9225 9231
0 9233 5 1 1 9232
0 9234 7 1 2 60038 9233
0 9235 5 1 1 9234
0 9236 7 9 2 41621 41791
0 9237 7 1 2 56903 60067
0 9238 7 1 2 59900 9237
0 9239 5 1 1 9238
0 9240 7 1 2 9235 9239
0 9241 7 1 2 9174 9240
0 9242 7 1 2 9060 9241
0 9243 7 1 2 8980 9242
0 9244 5 1 1 9243
0 9245 7 1 2 59334 9244
0 9246 5 1 1 9245
0 9247 7 3 2 41792 45144
0 9248 7 3 2 40988 60076
0 9249 5 1 1 60079
0 9250 7 1 2 8128 9249
0 9251 5 10 1 9250
0 9252 7 1 2 55172 54867
0 9253 7 2 2 58534 9252
0 9254 5 1 1 60092
0 9255 7 3 2 42318 49111
0 9256 7 4 2 45042 42544
0 9257 7 1 2 44636 60097
0 9258 7 1 2 60094 9257
0 9259 7 1 2 58779 9258
0 9260 5 1 1 9259
0 9261 7 1 2 9254 9260
0 9262 5 1 1 9261
0 9263 7 1 2 60082 9262
0 9264 5 1 1 9263
0 9265 7 6 2 45145 53872
0 9266 7 14 2 46369 60101
0 9267 7 2 2 51073 50920
0 9268 7 1 2 40781 60121
0 9269 5 1 1 9268
0 9270 7 1 2 8395 9269
0 9271 5 1 1 9270
0 9272 7 1 2 60107 9271
0 9273 5 1 1 9272
0 9274 7 2 2 43086 49485
0 9275 7 5 2 45043 41836
0 9276 7 2 2 60125 57010
0 9277 7 1 2 60123 60130
0 9278 7 1 2 58088 9277
0 9279 5 1 1 9278
0 9280 7 1 2 9273 9279
0 9281 5 1 1 9280
0 9282 7 1 2 45868 9281
0 9283 5 1 1 9282
0 9284 7 6 2 44193 60126
0 9285 7 6 2 60132 59927
0 9286 5 1 1 60138
0 9287 7 1 2 51200 60139
0 9288 5 1 1 9287
0 9289 7 1 2 53692 3782
0 9290 5 1 1 9289
0 9291 7 1 2 44491 60108
0 9292 7 1 2 9290 9291
0 9293 5 1 1 9292
0 9294 7 1 2 9288 9293
0 9295 5 1 1 9294
0 9296 7 1 2 43518 9295
0 9297 5 1 1 9296
0 9298 7 7 2 45146 45652
0 9299 7 3 2 41746 46370
0 9300 7 4 2 40948 60151
0 9301 7 2 2 47400 60154
0 9302 7 1 2 60144 60158
0 9303 5 1 1 9302
0 9304 7 1 2 9286 9303
0 9305 5 1 1 9304
0 9306 7 1 2 48746 9305
0 9307 5 1 1 9306
0 9308 7 2 2 45147 47966
0 9309 7 1 2 60160 60159
0 9310 5 1 1 9309
0 9311 7 1 2 9307 9310
0 9312 5 1 1 9311
0 9313 7 1 2 51886 9312
0 9314 5 1 1 9313
0 9315 7 10 2 48894 59629
0 9316 5 7 1 60162
0 9317 7 1 2 41341 56389
0 9318 5 3 1 9317
0 9319 7 1 2 60163 60179
0 9320 5 1 1 9319
0 9321 7 1 2 40364 9320
0 9322 5 1 1 9321
0 9323 7 7 2 46371 53873
0 9324 7 2 2 60182 60145
0 9325 5 1 1 60189
0 9326 7 1 2 60172 9325
0 9327 5 1 1 9326
0 9328 7 1 2 53176 9327
0 9329 7 1 2 9322 9328
0 9330 5 1 1 9329
0 9331 7 1 2 60109 56320
0 9332 5 1 1 9331
0 9333 7 1 2 50044 58492
0 9334 5 1 1 9333
0 9335 7 1 2 60140 9334
0 9336 5 1 1 9335
0 9337 7 1 2 9332 9336
0 9338 7 1 2 9330 9337
0 9339 7 1 2 9314 9338
0 9340 7 1 2 9297 9339
0 9341 5 1 1 9340
0 9342 7 1 2 54491 9341
0 9343 5 1 1 9342
0 9344 7 1 2 9283 9343
0 9345 5 1 1 9344
0 9346 7 1 2 55038 9345
0 9347 5 1 1 9346
0 9348 7 1 2 9264 9347
0 9349 5 1 1 9348
0 9350 7 1 2 46466 9349
0 9351 5 1 1 9350
0 9352 7 1 2 57011 57497
0 9353 7 1 2 59837 9352
0 9354 5 1 1 9353
0 9355 7 8 2 41201 54649
0 9356 5 1 1 60191
0 9357 7 3 2 50673 60192
0 9358 5 1 1 60199
0 9359 7 2 2 53874 56839
0 9360 5 2 1 60202
0 9361 7 8 2 45265 46372
0 9362 7 1 2 60206 58959
0 9363 7 1 2 57767 9362
0 9364 5 1 1 9363
0 9365 7 1 2 60204 9364
0 9366 5 1 1 9365
0 9367 7 1 2 60200 9366
0 9368 5 1 1 9367
0 9369 7 2 2 54682 49371
0 9370 7 1 2 47116 48662
0 9371 5 1 1 9370
0 9372 7 1 2 60214 9371
0 9373 5 1 1 9372
0 9374 7 1 2 9368 9373
0 9375 5 1 1 9374
0 9376 7 1 2 42545 9375
0 9377 5 1 1 9376
0 9378 7 2 2 42080 59419
0 9379 7 1 2 60216 56326
0 9380 5 1 1 9379
0 9381 7 10 2 43326 43674
0 9382 5 1 1 60218
0 9383 7 4 2 44492 60219
0 9384 5 1 1 60228
0 9385 7 1 2 60229 48028
0 9386 7 4 2 54579 52167
0 9387 7 9 2 45653 50429
0 9388 5 1 1 60236
0 9389 7 1 2 60232 60237
0 9390 7 1 2 9385 9389
0 9391 5 1 1 9390
0 9392 7 1 2 9380 9391
0 9393 5 1 1 9392
0 9394 7 1 2 43519 9393
0 9395 5 1 1 9394
0 9396 7 1 2 9377 9395
0 9397 7 1 2 9354 9396
0 9398 5 1 1 9397
0 9399 7 1 2 59680 46614
0 9400 7 1 2 9398 9399
0 9401 5 1 1 9400
0 9402 7 1 2 9351 9401
0 9403 5 1 1 9402
0 9404 7 1 2 41050 9403
0 9405 5 1 1 9404
0 9406 7 4 2 55039 53875
0 9407 5 1 1 60245
0 9408 7 1 2 56322 58376
0 9409 5 1 1 9408
0 9410 7 1 2 42546 9409
0 9411 5 1 1 9410
0 9412 7 1 2 58366 9411
0 9413 5 1 1 9412
0 9414 7 1 2 40782 9413
0 9415 5 1 1 9414
0 9416 7 1 2 9415 59592
0 9417 5 1 1 9416
0 9418 7 1 2 60246 9417
0 9419 5 1 1 9418
0 9420 7 2 2 51422 46615
0 9421 7 1 2 60095 60249
0 9422 7 1 2 58323 9421
0 9423 5 1 1 9422
0 9424 7 1 2 9419 9423
0 9425 5 1 1 9424
0 9426 7 1 2 46373 9425
0 9427 5 1 1 9426
0 9428 7 1 2 46616 60093
0 9429 5 1 1 9428
0 9430 7 1 2 9427 9429
0 9431 5 1 1 9430
0 9432 7 1 2 59563 9431
0 9433 5 1 1 9432
0 9434 7 1 2 9405 9433
0 9435 5 1 1 9434
0 9436 7 1 2 48265 9435
0 9437 5 1 1 9436
0 9438 7 64 2 46467 57625
0 9439 5 1 1 60251
0 9440 7 2 2 44054 58405
0 9441 5 1 1 60315
0 9442 7 2 2 55137 47322
0 9443 5 1 1 60317
0 9444 7 1 2 54956 51344
0 9445 7 1 2 60318 9444
0 9446 5 1 1 9445
0 9447 7 1 2 9441 9446
0 9448 5 1 1 9447
0 9449 7 1 2 60252 9448
0 9450 5 1 1 9449
0 9451 7 1 2 45654 59125
0 9452 7 1 2 59579 9451
0 9453 5 1 1 9452
0 9454 7 1 2 9450 9453
0 9455 5 1 1 9454
0 9456 7 1 2 54667 9455
0 9457 5 1 1 9456
0 9458 7 14 2 45084 46468
0 9459 7 3 2 54070 60319
0 9460 7 12 2 40783 44238
0 9461 7 1 2 42961 51038
0 9462 7 1 2 60336 9461
0 9463 7 2 2 60333 9462
0 9464 5 1 1 60348
0 9465 7 1 2 41928 49914
0 9466 7 1 2 60349 9465
0 9467 5 1 1 9466
0 9468 7 7 2 45655 43177
0 9469 7 3 2 46617 60350
0 9470 5 3 1 60357
0 9471 7 1 2 56840 52857
0 9472 7 1 2 50361 9471
0 9473 7 1 2 60358 9472
0 9474 5 1 1 9473
0 9475 7 1 2 9467 9474
0 9476 5 1 1 9475
0 9477 7 1 2 47323 9476
0 9478 5 1 1 9477
0 9479 7 11 2 43087 43178
0 9480 7 2 2 45431 60363
0 9481 7 1 2 45656 48325
0 9482 7 2 2 60374 9481
0 9483 7 6 2 41747 41793
0 9484 7 3 2 40989 47401
0 9485 7 1 2 60378 60384
0 9486 7 1 2 60376 9485
0 9487 5 1 1 9486
0 9488 7 1 2 9464 9487
0 9489 5 1 1 9488
0 9490 7 1 2 47639 9489
0 9491 5 1 1 9490
0 9492 7 3 2 40990 44493
0 9493 7 2 2 60379 60387
0 9494 7 1 2 43520 60390
0 9495 7 1 2 60377 9494
0 9496 5 1 1 9495
0 9497 7 1 2 9491 9496
0 9498 5 1 1 9497
0 9499 7 1 2 44637 9498
0 9500 5 1 1 9499
0 9501 7 1 2 9478 9500
0 9502 5 1 1 9501
0 9503 7 1 2 43675 9502
0 9504 5 1 1 9503
0 9505 7 15 2 41794 43179
0 9506 7 5 2 60392 59116
0 9507 7 1 2 54601 55329
0 9508 7 1 2 60407 9507
0 9509 7 1 2 59922 9508
0 9510 5 1 1 9509
0 9511 7 1 2 9504 9510
0 9512 7 1 2 9457 9511
0 9513 5 1 1 9512
0 9514 7 1 2 45869 9513
0 9515 5 1 1 9514
0 9516 7 1 2 53713 54668
0 9517 5 1 1 9516
0 9518 7 1 2 54938 9517
0 9519 5 1 1 9518
0 9520 7 1 2 41929 9519
0 9521 5 1 1 9520
0 9522 7 1 2 54548 60180
0 9523 5 1 1 9522
0 9524 7 1 2 40365 9523
0 9525 5 1 1 9524
0 9526 7 1 2 42081 59104
0 9527 7 1 2 9525 9526
0 9528 5 1 1 9527
0 9529 7 1 2 9521 9528
0 9530 5 1 1 9529
0 9531 7 1 2 47640 9530
0 9532 5 1 1 9531
0 9533 7 1 2 50832 54116
0 9534 5 1 1 9533
0 9535 7 1 2 58397 9534
0 9536 5 1 1 9535
0 9537 7 1 2 54549 9536
0 9538 5 1 1 9537
0 9539 7 1 2 9532 9538
0 9540 7 1 2 54640 3293
0 9541 5 1 1 9540
0 9542 7 1 2 46833 9541
0 9543 5 1 1 9542
0 9544 7 1 2 43327 54637
0 9545 5 1 1 9544
0 9546 7 1 2 46709 54924
0 9547 5 1 1 9546
0 9548 7 1 2 9545 9547
0 9549 7 1 2 9543 9548
0 9550 5 1 1 9549
0 9551 7 1 2 42082 9550
0 9552 5 1 1 9551
0 9553 7 1 2 45657 56265
0 9554 5 1 1 9553
0 9555 7 1 2 54550 9554
0 9556 5 1 1 9555
0 9557 7 1 2 59108 9556
0 9558 7 1 2 9552 9557
0 9559 5 1 1 9558
0 9560 7 1 2 47721 9559
0 9561 5 1 1 9560
0 9562 7 1 2 41092 54556
0 9563 5 1 1 9562
0 9564 7 1 2 59106 9563
0 9565 5 1 1 9564
0 9566 7 3 2 43676 54778
0 9567 5 2 1 60412
0 9568 7 1 2 44401 47967
0 9569 5 2 1 9568
0 9570 7 1 2 60415 60417
0 9571 5 1 1 9570
0 9572 7 1 2 54669 9571
0 9573 5 1 1 9572
0 9574 7 1 2 54939 9573
0 9575 7 1 2 9565 9574
0 9576 5 1 1 9575
0 9577 7 1 2 43328 9576
0 9578 5 1 1 9577
0 9579 7 1 2 58759 54909
0 9580 5 1 1 9579
0 9581 7 1 2 54551 9580
0 9582 5 1 1 9581
0 9583 7 1 2 44402 60413
0 9584 7 1 2 54670 9583
0 9585 5 1 1 9584
0 9586 7 1 2 9582 9585
0 9587 7 1 2 9578 9586
0 9588 5 1 1 9587
0 9589 7 1 2 51887 9588
0 9590 5 1 1 9589
0 9591 7 1 2 9561 9590
0 9592 7 1 2 9539 9591
0 9593 5 1 1 9592
0 9594 7 1 2 60253 9593
0 9595 5 1 1 9594
0 9596 7 2 2 47582 46737
0 9597 5 5 1 60419
0 9598 7 1 2 39977 58638
0 9599 5 1 1 9598
0 9600 7 4 2 60421 9599
0 9601 5 2 1 60426
0 9602 7 1 2 47777 60430
0 9603 5 7 1 9602
0 9604 7 1 2 42083 60432
0 9605 5 2 1 9604
0 9606 7 1 2 42319 59871
0 9607 5 3 1 9606
0 9608 7 1 2 59555 60441
0 9609 7 1 2 60439 9608
0 9610 5 2 1 9609
0 9611 7 28 2 40991 60393
0 9612 5 6 1 60446
0 9613 7 1 2 60447 56635
0 9614 7 1 2 60444 9613
0 9615 5 1 1 9614
0 9616 7 1 2 9595 9615
0 9617 5 1 1 9616
0 9618 7 1 2 54492 9617
0 9619 5 1 1 9618
0 9620 7 2 2 57192 52864
0 9621 7 1 2 54493 52051
0 9622 5 2 1 9621
0 9623 7 1 2 8452 60482
0 9624 5 1 1 9623
0 9625 7 1 2 60480 9624
0 9626 5 1 1 9625
0 9627 7 1 2 52268 8761
0 9628 5 1 1 9627
0 9629 7 3 2 43521 47179
0 9630 7 1 2 48747 60484
0 9631 5 1 1 9630
0 9632 7 1 2 59556 9631
0 9633 5 1 1 9632
0 9634 7 1 2 49314 50507
0 9635 5 1 1 9634
0 9636 7 1 2 49486 50508
0 9637 5 2 1 9636
0 9638 7 1 2 9635 60487
0 9639 7 1 2 9633 9638
0 9640 7 1 2 9628 9639
0 9641 5 1 1 9640
0 9642 7 1 2 44055 9641
0 9643 5 1 1 9642
0 9644 7 1 2 9643 8483
0 9645 5 1 1 9644
0 9646 7 1 2 45870 9645
0 9647 5 1 1 9646
0 9648 7 1 2 53719 60005
0 9649 5 1 1 9648
0 9650 7 1 2 47641 58910
0 9651 5 1 1 9650
0 9652 7 1 2 42084 51607
0 9653 5 2 1 9652
0 9654 7 1 2 58275 58767
0 9655 7 1 2 60489 9654
0 9656 7 1 2 9651 9655
0 9657 7 2 2 9649 9656
0 9658 5 1 1 60491
0 9659 7 1 2 54494 9658
0 9660 5 1 1 9659
0 9661 7 2 2 41342 54529
0 9662 5 2 1 60493
0 9663 7 2 2 42085 52322
0 9664 7 1 2 50224 60497
0 9665 7 1 2 60494 9664
0 9666 5 1 1 9665
0 9667 7 1 2 59829 9666
0 9668 5 1 1 9667
0 9669 7 1 2 40366 9668
0 9670 5 1 1 9669
0 9671 7 1 2 44638 46905
0 9672 5 3 1 9671
0 9673 7 1 2 45432 60499
0 9674 5 1 1 9673
0 9675 7 2 2 42320 51865
0 9676 5 1 1 60502
0 9677 7 1 2 46857 52730
0 9678 5 1 1 9677
0 9679 7 1 2 9676 9678
0 9680 5 1 1 9679
0 9681 7 1 2 9674 9680
0 9682 5 1 1 9681
0 9683 7 1 2 54471 9682
0 9684 5 1 1 9683
0 9685 7 1 2 9670 9684
0 9686 5 1 1 9685
0 9687 7 1 2 39978 9686
0 9688 5 1 1 9687
0 9689 7 1 2 9660 9688
0 9690 7 1 2 9647 9689
0 9691 5 1 1 9690
0 9692 7 17 2 46242 57243
0 9693 7 1 2 41748 60504
0 9694 7 1 2 9691 9693
0 9695 5 1 1 9694
0 9696 7 1 2 9626 9695
0 9697 5 1 1 9696
0 9698 7 1 2 55040 9697
0 9699 5 1 1 9698
0 9700 7 1 2 9619 9699
0 9701 7 1 2 9515 9700
0 9702 5 1 1 9701
0 9703 7 1 2 58544 9702
0 9704 5 1 1 9703
0 9705 7 1 2 53416 54558
0 9706 5 1 1 9705
0 9707 7 1 2 40784 8391
0 9708 5 1 1 9707
0 9709 7 1 2 45871 60316
0 9710 5 1 1 9709
0 9711 7 1 2 9708 9710
0 9712 5 1 1 9711
0 9713 7 1 2 54671 9712
0 9714 5 1 1 9713
0 9715 7 1 2 9706 9714
0 9716 5 1 1 9715
0 9717 7 1 2 46618 59344
0 9718 7 1 2 9716 9717
0 9719 5 1 1 9718
0 9720 7 1 2 9704 9719
0 9721 5 1 1 9720
0 9722 7 1 2 4821 48973
0 9723 5 1 1 9722
0 9724 7 1 2 7105 9723
0 9725 7 1 2 9721 9724
0 9726 5 1 1 9725
0 9727 7 1 2 9437 9726
0 9728 7 1 2 9246 9727
0 9729 7 1 2 8612 9728
0 9730 7 1 2 8312 9729
0 9731 7 1 2 7843 9730
0 9732 5 1 1 9731
0 9733 7 1 2 58017 9732
0 9734 5 1 1 9733
0 9735 7 1 2 45658 51776
0 9736 5 1 1 9735
0 9737 7 2 2 41093 42086
0 9738 5 2 1 60521
0 9739 7 1 2 60523 53573
0 9740 5 1 1 9739
0 9741 7 1 2 41930 9740
0 9742 5 1 1 9741
0 9743 7 1 2 42321 53551
0 9744 7 1 2 9742 9743
0 9745 5 1 1 9744
0 9746 7 1 2 45872 9745
0 9747 7 1 2 9736 9746
0 9748 5 1 1 9747
0 9749 7 2 2 52441 54901
0 9750 5 1 1 60525
0 9751 7 1 2 40189 60526
0 9752 5 1 1 9751
0 9753 7 1 2 50311 52481
0 9754 5 1 1 9753
0 9755 7 1 2 9752 9754
0 9756 7 1 2 9748 9755
0 9757 5 1 1 9756
0 9758 7 1 2 46679 9757
0 9759 5 1 1 9758
0 9760 7 1 2 47245 5363
0 9761 5 8 1 9760
0 9762 7 1 2 52250 47984
0 9763 5 1 1 9762
0 9764 7 1 2 52442 9763
0 9765 5 1 1 9764
0 9766 7 1 2 52488 9765
0 9767 5 1 1 9766
0 9768 7 1 2 60527 9767
0 9769 5 1 1 9768
0 9770 7 3 2 47324 50856
0 9771 7 1 2 60535 54059
0 9772 5 1 1 9771
0 9773 7 1 2 53408 51382
0 9774 5 1 1 9773
0 9775 7 1 2 47642 9774
0 9776 7 1 2 59642 9775
0 9777 5 1 1 9776
0 9778 7 1 2 9772 9777
0 9779 5 1 1 9778
0 9780 7 1 2 56529 9779
0 9781 5 1 1 9780
0 9782 7 1 2 9769 9781
0 9783 7 1 2 9759 9782
0 9784 5 1 1 9783
0 9785 7 1 2 53939 9784
0 9786 5 1 1 9785
0 9787 7 1 2 42322 55957
0 9788 5 2 1 9787
0 9789 7 1 2 41094 60538
0 9790 5 1 1 9789
0 9791 7 2 2 48628 48874
0 9792 5 1 1 60540
0 9793 7 1 2 9790 9792
0 9794 5 1 1 9793
0 9795 7 1 2 45433 9794
0 9796 5 1 1 9795
0 9797 7 1 2 863 9796
0 9798 5 1 1 9797
0 9799 7 1 2 47225 9798
0 9800 5 1 1 9799
0 9801 7 4 2 39979 51741
0 9802 5 1 1 60542
0 9803 7 3 2 57914 60543
0 9804 5 1 1 60546
0 9805 7 1 2 43677 56308
0 9806 7 1 2 59826 9805
0 9807 5 1 1 9806
0 9808 7 1 2 56279 9807
0 9809 5 1 1 9808
0 9810 7 1 2 9804 9809
0 9811 5 1 1 9810
0 9812 7 1 2 46680 9811
0 9813 5 1 1 9812
0 9814 7 1 2 9800 9813
0 9815 5 1 1 9814
0 9816 7 1 2 41202 9815
0 9817 5 1 1 9816
0 9818 7 2 2 50299 46681
0 9819 7 1 2 59872 60549
0 9820 5 1 1 9819
0 9821 7 2 2 39980 49487
0 9822 7 1 2 60551 58392
0 9823 5 1 1 9822
0 9824 7 1 2 43522 9823
0 9825 5 1 1 9824
0 9826 7 1 2 58139 6601
0 9827 5 2 1 9826
0 9828 7 1 2 47226 60553
0 9829 7 1 2 9825 9828
0 9830 5 1 1 9829
0 9831 7 1 2 9820 9830
0 9832 7 1 2 9817 9831
0 9833 5 1 1 9832
0 9834 7 1 2 42547 9833
0 9835 5 1 1 9834
0 9836 7 1 2 47246 1941
0 9837 5 4 1 9836
0 9838 7 3 2 55452 56540
0 9839 5 1 1 60559
0 9840 7 1 2 9839 53791
0 9841 5 1 1 9840
0 9842 7 1 2 60555 9841
0 9843 5 1 1 9842
0 9844 7 1 2 47402 56123
0 9845 5 1 1 9844
0 9846 7 1 2 54064 9845
0 9847 5 1 1 9846
0 9848 7 1 2 56499 9847
0 9849 5 1 1 9848
0 9850 7 1 2 47325 56103
0 9851 5 1 1 9850
0 9852 7 1 2 9849 9851
0 9853 5 1 1 9852
0 9854 7 1 2 45873 9853
0 9855 5 1 1 9854
0 9856 7 1 2 9843 9855
0 9857 7 1 2 9835 9856
0 9858 5 1 1 9857
0 9859 7 1 2 54134 9858
0 9860 5 1 1 9859
0 9861 7 1 2 9786 9860
0 9862 5 1 1 9861
0 9863 7 1 2 43873 9862
0 9864 5 1 1 9863
0 9865 7 10 2 45266 52392
0 9866 5 1 1 60562
0 9867 7 1 2 40367 58191
0 9868 5 1 1 9867
0 9869 7 1 2 41343 55495
0 9870 5 1 1 9869
0 9871 7 1 2 9868 9870
0 9872 5 1 1 9871
0 9873 7 1 2 60563 9872
0 9874 5 1 1 9873
0 9875 7 1 2 1705 9874
0 9876 5 1 1 9875
0 9877 7 12 2 42794 43088
0 9878 7 3 2 60572 54860
0 9879 7 1 2 57724 60584
0 9880 7 1 2 9876 9879
0 9881 5 1 1 9880
0 9882 7 1 2 9864 9881
0 9883 5 1 1 9882
0 9884 7 1 2 44754 9883
0 9885 5 1 1 9884
0 9886 7 8 2 40949 53341
0 9887 7 2 2 51916 58979
0 9888 7 1 2 60587 60595
0 9889 5 1 1 9888
0 9890 7 6 2 44194 50745
0 9891 7 2 2 56175 60597
0 9892 7 1 2 56623 60603
0 9893 5 1 1 9892
0 9894 7 1 2 9889 9893
0 9895 5 1 1 9894
0 9896 7 1 2 47778 9895
0 9897 5 1 1 9896
0 9898 7 2 2 53302 56624
0 9899 7 1 2 57449 54844
0 9900 7 2 2 60605 9899
0 9901 5 1 1 60607
0 9902 7 1 2 45267 60608
0 9903 5 1 1 9902
0 9904 7 1 2 9897 9903
0 9905 5 1 1 9904
0 9906 7 1 2 39981 9905
0 9907 5 1 1 9906
0 9908 7 1 2 57867 58192
0 9909 5 1 1 9908
0 9910 7 3 2 56810 50967
0 9911 7 1 2 46374 60609
0 9912 5 1 1 9911
0 9913 7 1 2 9909 9912
0 9914 5 1 1 9913
0 9915 7 1 2 42548 9914
0 9916 5 1 1 9915
0 9917 7 1 2 9907 9916
0 9918 5 1 1 9917
0 9919 7 1 2 40368 9918
0 9920 5 1 1 9919
0 9921 7 1 2 52323 53195
0 9922 5 1 1 9921
0 9923 7 1 2 1853 9922
0 9924 5 1 1 9923
0 9925 7 1 2 41344 53940
0 9926 7 1 2 9924 9925
0 9927 5 1 1 9926
0 9928 7 1 2 9920 9927
0 9929 5 1 1 9928
0 9930 7 1 2 41095 9929
0 9931 5 1 1 9930
0 9932 7 1 2 58288 53153
0 9933 5 1 1 9932
0 9934 7 1 2 54135 9933
0 9935 5 1 1 9934
0 9936 7 1 2 60205 9935
0 9937 5 1 1 9936
0 9938 7 1 2 50181 55211
0 9939 7 1 2 9937 9938
0 9940 5 1 1 9939
0 9941 7 1 2 9931 9940
0 9942 5 1 1 9941
0 9943 7 1 2 44921 55586
0 9944 7 1 2 9942 9943
0 9945 5 1 1 9944
0 9946 7 1 2 9885 9945
0 9947 5 1 1 9946
0 9948 7 1 2 44056 9947
0 9949 5 1 1 9948
0 9950 7 5 2 53876 58980
0 9951 5 5 1 60612
0 9952 7 2 2 42795 54381
0 9953 5 1 1 60622
0 9954 7 1 2 55395 9953
0 9955 5 2 1 9954
0 9956 7 1 2 60613 60624
0 9957 5 1 1 9956
0 9958 7 1 2 47403 54382
0 9959 5 1 1 9958
0 9960 7 2 2 47326 54403
0 9961 7 1 2 41931 60626
0 9962 5 1 1 9961
0 9963 7 1 2 9959 9962
0 9964 5 1 1 9963
0 9965 7 1 2 51333 9964
0 9966 5 1 1 9965
0 9967 7 1 2 55387 50857
0 9968 5 1 1 9967
0 9969 7 1 2 9966 9968
0 9970 5 1 1 9969
0 9971 7 1 2 54136 9970
0 9972 5 1 1 9971
0 9973 7 1 2 9957 9972
0 9974 5 1 1 9973
0 9975 7 1 2 47643 9974
0 9976 5 1 1 9975
0 9977 7 3 2 41749 59928
0 9978 7 1 2 58931 60628
0 9979 5 2 1 9978
0 9980 7 6 2 45434 46375
0 9981 5 1 1 60633
0 9982 7 1 2 48895 60634
0 9983 5 2 1 9982
0 9984 7 1 2 57076 60639
0 9985 5 2 1 9984
0 9986 7 1 2 47722 60641
0 9987 5 2 1 9986
0 9988 7 1 2 60631 60643
0 9989 5 2 1 9988
0 9990 7 1 2 55235 60645
0 9991 5 1 1 9990
0 9992 7 4 2 44755 53819
0 9993 5 2 1 60647
0 9994 7 1 2 53941 58713
0 9995 5 1 1 9994
0 9996 7 1 2 46834 52555
0 9997 7 1 2 51804 9996
0 9998 5 1 1 9997
0 9999 7 1 2 44403 50695
0 10000 5 5 1 9999
0 10001 7 1 2 60653 48414
0 10002 7 1 2 9998 10001
0 10003 5 1 1 10002
0 10004 7 1 2 54137 10003
0 10005 5 1 1 10004
0 10006 7 1 2 9995 10005
0 10007 5 1 1 10006
0 10008 7 1 2 60648 10007
0 10009 5 1 1 10008
0 10010 7 1 2 9991 10009
0 10011 5 1 1 10010
0 10012 7 1 2 43874 10011
0 10013 5 1 1 10012
0 10014 7 1 2 53206 60646
0 10015 5 1 1 10014
0 10016 7 1 2 59253 55723
0 10017 7 1 2 60606 10016
0 10018 5 1 1 10017
0 10019 7 1 2 10015 10018
0 10020 5 1 1 10019
0 10021 7 1 2 42796 10020
0 10022 5 1 1 10021
0 10023 7 1 2 57040 58256
0 10024 7 1 2 60625 10023
0 10025 5 1 1 10024
0 10026 7 1 2 58579 57832
0 10027 7 1 2 55939 10026
0 10028 5 1 1 10027
0 10029 7 1 2 10025 10028
0 10030 5 1 1 10029
0 10031 7 1 2 51888 10030
0 10032 5 1 1 10031
0 10033 7 1 2 10022 10032
0 10034 7 1 2 10013 10033
0 10035 7 1 2 9976 10034
0 10036 5 1 1 10035
0 10037 7 1 2 44057 10036
0 10038 5 1 1 10037
0 10039 7 2 2 44195 52760
0 10040 7 2 2 56625 60658
0 10041 7 1 2 54455 60660
0 10042 7 1 2 47837 10041
0 10043 5 1 1 10042
0 10044 7 1 2 41622 10043
0 10045 7 1 2 10038 10044
0 10046 5 1 1 10045
0 10047 7 1 2 54310 51104
0 10048 5 1 1 10047
0 10049 7 1 2 54383 54212
0 10050 7 1 2 47834 10049
0 10051 5 1 1 10050
0 10052 7 1 2 10048 10051
0 10053 5 1 1 10052
0 10054 7 1 2 42797 10053
0 10055 5 1 1 10054
0 10056 7 1 2 55388 51250
0 10057 5 1 1 10056
0 10058 7 1 2 10055 10057
0 10059 5 1 1 10058
0 10060 7 1 2 40785 10059
0 10061 5 1 1 10060
0 10062 7 3 2 45874 49577
0 10063 5 1 1 60662
0 10064 7 1 2 54404 51251
0 10065 5 1 1 10064
0 10066 7 1 2 10063 10065
0 10067 5 1 1 10066
0 10068 7 1 2 45435 10067
0 10069 5 1 1 10068
0 10070 7 6 2 43329 40585
0 10071 7 3 2 44404 60665
0 10072 7 2 2 41450 54428
0 10073 7 1 2 60671 60674
0 10074 5 1 1 10073
0 10075 7 1 2 10069 10074
0 10076 5 1 1 10075
0 10077 7 1 2 58300 10076
0 10078 5 1 1 10077
0 10079 7 1 2 10061 10078
0 10080 5 1 1 10079
0 10081 7 1 2 54138 10080
0 10082 5 1 1 10081
0 10083 7 1 2 41932 52852
0 10084 5 1 1 10083
0 10085 7 1 2 51897 10084
0 10086 5 1 1 10085
0 10087 7 1 2 53138 53574
0 10088 5 1 1 10087
0 10089 7 1 2 1269 6637
0 10090 5 6 1 10089
0 10091 7 1 2 54384 60676
0 10092 7 1 2 10088 10091
0 10093 7 1 2 10086 10092
0 10094 5 1 1 10093
0 10095 7 1 2 50867 54495
0 10096 7 1 2 52117 10095
0 10097 5 1 1 10096
0 10098 7 1 2 10094 10097
0 10099 5 1 1 10098
0 10100 7 1 2 53942 10099
0 10101 5 1 1 10100
0 10102 7 1 2 44922 10101
0 10103 7 1 2 10082 10102
0 10104 5 1 1 10103
0 10105 7 1 2 42323 10104
0 10106 7 1 2 10046 10105
0 10107 5 1 1 10106
0 10108 7 1 2 53943 51326
0 10109 5 1 1 10108
0 10110 7 1 2 46091 54139
0 10111 7 1 2 54305 10110
0 10112 5 1 1 10111
0 10113 7 1 2 10109 10112
0 10114 5 1 1 10113
0 10115 7 1 2 43330 10114
0 10116 5 1 1 10115
0 10117 7 6 2 48896 58796
0 10118 5 1 1 60682
0 10119 7 1 2 60683 59862
0 10120 5 1 1 10119
0 10121 7 1 2 10116 10120
0 10122 5 1 1 10121
0 10123 7 1 2 44923 10122
0 10124 5 1 1 10123
0 10125 7 1 2 44058 60684
0 10126 7 1 2 56404 10125
0 10127 5 1 1 10126
0 10128 7 1 2 10124 10127
0 10129 5 1 1 10128
0 10130 7 1 2 54405 10129
0 10131 5 1 1 10130
0 10132 7 1 2 43331 58425
0 10133 5 1 1 10132
0 10134 7 1 2 55279 10133
0 10135 5 1 1 10134
0 10136 7 1 2 60685 10135
0 10137 5 1 1 10136
0 10138 7 5 2 43332 44059
0 10139 7 2 2 41750 56773
0 10140 7 2 2 56673 60693
0 10141 7 1 2 60688 60695
0 10142 5 1 1 10141
0 10143 7 1 2 10137 10142
0 10144 5 1 1 10143
0 10145 7 1 2 55340 10144
0 10146 5 1 1 10145
0 10147 7 3 2 44924 50758
0 10148 5 3 1 60697
0 10149 7 1 2 47247 60700
0 10150 5 7 1 10149
0 10151 7 7 2 57027 54861
0 10152 7 1 2 48546 60689
0 10153 7 1 2 60710 10152
0 10154 7 1 2 60703 10153
0 10155 5 1 1 10154
0 10156 7 1 2 10146 10155
0 10157 7 1 2 10131 10156
0 10158 5 1 1 10157
0 10159 7 1 2 47192 10158
0 10160 5 1 1 10159
0 10161 7 2 2 50759 52168
0 10162 7 1 2 57144 58683
0 10163 7 2 2 51232 10162
0 10164 7 1 2 60717 60719
0 10165 5 2 1 10164
0 10166 7 2 2 50410 58301
0 10167 5 2 1 60723
0 10168 7 1 2 41451 58880
0 10169 5 1 1 10168
0 10170 7 1 2 60725 10169
0 10171 5 1 1 10170
0 10172 7 3 2 42549 10171
0 10173 5 2 1 60727
0 10174 7 1 2 44060 60704
0 10175 5 1 1 10174
0 10176 7 1 2 49346 10175
0 10177 5 2 1 10176
0 10178 7 1 2 54385 60732
0 10179 5 1 1 10178
0 10180 7 1 2 60730 10179
0 10181 5 1 1 10180
0 10182 7 4 2 43333 53944
0 10183 7 1 2 47175 60734
0 10184 7 1 2 10181 10183
0 10185 5 1 1 10184
0 10186 7 1 2 60721 10185
0 10187 7 1 2 10160 10186
0 10188 5 1 1 10187
0 10189 7 1 2 43523 10188
0 10190 5 1 1 10189
0 10191 7 1 2 57041 54386
0 10192 5 1 1 10191
0 10193 7 6 2 45659 46376
0 10194 7 3 2 43334 45044
0 10195 5 1 1 60744
0 10196 7 5 2 44196 60745
0 10197 7 1 2 60738 60747
0 10198 7 1 2 54406 10197
0 10199 5 1 1 10198
0 10200 7 1 2 10192 10199
0 10201 5 1 1 10200
0 10202 7 1 2 49198 10201
0 10203 5 1 1 10202
0 10204 7 2 2 60748 57002
0 10205 5 1 1 60752
0 10206 7 1 2 41623 60753
0 10207 5 1 1 10206
0 10208 7 1 2 53945 50395
0 10209 5 1 1 10208
0 10210 7 1 2 10207 10209
0 10211 5 1 1 10210
0 10212 7 1 2 54496 10211
0 10213 5 1 1 10212
0 10214 7 1 2 10203 10213
0 10215 5 1 1 10214
0 10216 7 1 2 42798 10215
0 10217 5 1 1 10216
0 10218 7 2 2 53946 58302
0 10219 5 1 1 60754
0 10220 7 1 2 56023 55533
0 10221 5 1 1 10220
0 10222 7 1 2 43875 10221
0 10223 5 1 1 10222
0 10224 7 1 2 54996 51728
0 10225 5 1 1 10224
0 10226 7 1 2 10223 10225
0 10227 5 1 1 10226
0 10228 7 1 2 60755 10227
0 10229 5 1 1 10228
0 10230 7 1 2 10217 10229
0 10231 5 1 1 10230
0 10232 7 1 2 54750 10231
0 10233 5 1 1 10232
0 10234 7 1 2 60722 10233
0 10235 5 1 1 10234
0 10236 7 1 2 46835 10235
0 10237 5 1 1 10236
0 10238 7 3 2 48547 51770
0 10239 5 1 1 60756
0 10240 7 1 2 60733 60757
0 10241 5 1 1 10240
0 10242 7 1 2 49280 60705
0 10243 5 1 1 10242
0 10244 7 1 2 10241 10243
0 10245 5 1 1 10244
0 10246 7 1 2 53947 10245
0 10247 5 1 1 10246
0 10248 7 3 2 50658 51392
0 10249 5 2 1 60759
0 10250 7 4 2 46377 49364
0 10251 7 8 2 39982 41203
0 10252 5 1 1 60768
0 10253 7 1 2 10252 57012
0 10254 7 1 2 60764 10253
0 10255 7 1 2 60760 10254
0 10256 5 1 1 10255
0 10257 7 1 2 10247 10256
0 10258 5 1 1 10257
0 10259 7 1 2 45875 10258
0 10260 5 1 1 10259
0 10261 7 5 2 41933 47082
0 10262 7 3 2 43089 47404
0 10263 7 2 2 53877 60781
0 10264 5 2 1 60784
0 10265 7 1 2 60776 60785
0 10266 7 1 2 60728 10265
0 10267 5 1 1 10266
0 10268 7 1 2 10260 10267
0 10269 7 1 2 10237 10268
0 10270 7 1 2 10190 10269
0 10271 7 1 2 10107 10270
0 10272 5 1 1 10271
0 10273 7 1 2 44639 10272
0 10274 5 1 1 10273
0 10275 7 5 2 41934 51917
0 10276 5 1 1 60788
0 10277 7 1 2 10276 53391
0 10278 5 2 1 10277
0 10279 7 1 2 45436 60793
0 10280 5 1 1 10279
0 10281 7 2 2 45876 60433
0 10282 7 1 2 48156 60795
0 10283 5 1 1 10282
0 10284 7 1 2 10280 10283
0 10285 5 1 1 10284
0 10286 7 1 2 46682 10285
0 10287 5 1 1 10286
0 10288 7 2 2 47892 60420
0 10289 5 2 1 60797
0 10290 7 4 2 42799 48157
0 10291 7 1 2 60801 56001
0 10292 7 1 2 60799 10291
0 10293 5 1 1 10292
0 10294 7 1 2 10287 10293
0 10295 5 1 1 10294
0 10296 7 1 2 54140 10295
0 10297 5 1 1 10296
0 10298 7 2 2 53342 57725
0 10299 7 1 2 56674 56116
0 10300 7 1 2 60805 10299
0 10301 5 1 1 10300
0 10302 7 1 2 10297 10301
0 10303 5 1 1 10302
0 10304 7 1 2 49281 10303
0 10305 5 1 1 10304
0 10306 7 1 2 10274 10305
0 10307 5 1 1 10306
0 10308 7 1 2 43678 10307
0 10309 5 1 1 10308
0 10310 7 5 2 40586 51219
0 10311 7 1 2 56881 52532
0 10312 7 1 2 51299 10311
0 10313 7 2 2 60807 10312
0 10314 5 1 1 60812
0 10315 7 1 2 46793 50522
0 10316 5 2 1 10315
0 10317 7 1 2 50497 60814
0 10318 5 7 1 10317
0 10319 7 1 2 60813 60816
0 10320 5 1 1 10319
0 10321 7 3 2 40587 45268
0 10322 7 1 2 41624 60823
0 10323 7 1 2 57556 10322
0 10324 7 2 2 45045 57450
0 10325 7 3 2 53232 50760
0 10326 7 1 2 60826 60828
0 10327 7 1 2 10323 10326
0 10328 5 1 1 10327
0 10329 7 3 2 43876 45269
0 10330 5 2 1 60831
0 10331 7 3 2 41096 50326
0 10332 5 2 1 60836
0 10333 7 1 2 42087 60837
0 10334 5 1 1 10333
0 10335 7 1 2 60834 10334
0 10336 5 1 1 10335
0 10337 7 1 2 40190 10336
0 10338 5 1 1 10337
0 10339 7 1 2 41097 51179
0 10340 5 1 1 10339
0 10341 7 1 2 10338 10340
0 10342 5 3 1 10341
0 10343 7 1 2 53878 54267
0 10344 7 1 2 48963 10343
0 10345 7 1 2 60841 10344
0 10346 5 1 1 10345
0 10347 7 1 2 10328 10346
0 10348 5 1 1 10347
0 10349 7 1 2 49488 10348
0 10350 5 1 1 10349
0 10351 7 1 2 10320 10350
0 10352 5 1 1 10351
0 10353 7 1 2 39983 10352
0 10354 5 1 1 10353
0 10355 7 2 2 56811 56949
0 10356 7 2 2 41452 50640
0 10357 7 1 2 60846 60829
0 10358 7 1 2 60844 10357
0 10359 5 1 1 10358
0 10360 7 1 2 56368 49856
0 10361 7 1 2 51170 10360
0 10362 7 1 2 55400 10361
0 10363 5 1 1 10362
0 10364 7 1 2 10359 10363
0 10365 7 1 2 10354 10364
0 10366 5 1 1 10365
0 10367 7 1 2 58623 10366
0 10368 5 1 1 10367
0 10369 7 1 2 50380 49246
0 10370 5 1 1 10369
0 10371 7 5 2 45270 51531
0 10372 7 1 2 56412 60848
0 10373 5 1 1 10372
0 10374 7 1 2 10370 10373
0 10375 5 1 1 10374
0 10376 7 1 2 42088 10375
0 10377 5 1 1 10376
0 10378 7 1 2 44061 52665
0 10379 5 1 1 10378
0 10380 7 1 2 7572 10379
0 10381 5 1 1 10380
0 10382 7 1 2 50833 10381
0 10383 5 1 1 10382
0 10384 7 1 2 10377 10383
0 10385 5 1 1 10384
0 10386 7 1 2 54387 10385
0 10387 5 1 1 10386
0 10388 7 1 2 58438 60729
0 10389 5 1 1 10388
0 10390 7 1 2 10387 10389
0 10391 5 1 1 10390
0 10392 7 1 2 53948 10391
0 10393 5 1 1 10392
0 10394 7 1 2 48312 50113
0 10395 5 1 1 10394
0 10396 7 1 2 4773 10395
0 10397 5 1 1 10396
0 10398 7 1 2 41453 10397
0 10399 5 1 1 10398
0 10400 7 1 2 46836 60724
0 10401 5 1 1 10400
0 10402 7 1 2 10399 10401
0 10403 5 1 1 10402
0 10404 7 1 2 43335 10403
0 10405 5 1 1 10404
0 10406 7 1 2 57893 60726
0 10407 5 1 1 10406
0 10408 7 1 2 46710 10407
0 10409 5 1 1 10408
0 10410 7 1 2 10405 10409
0 10411 5 1 1 10410
0 10412 7 1 2 54429 54141
0 10413 7 1 2 10411 10412
0 10414 5 1 1 10413
0 10415 7 1 2 10393 10414
0 10416 5 1 1 10415
0 10417 7 1 2 44494 10416
0 10418 5 1 1 10417
0 10419 7 1 2 54388 49247
0 10420 5 1 1 10419
0 10421 7 1 2 60731 10420
0 10422 5 2 1 10421
0 10423 7 2 2 50834 60614
0 10424 7 1 2 60853 60855
0 10425 5 1 1 10424
0 10426 7 1 2 53233 51300
0 10427 7 1 2 60720 10426
0 10428 5 1 1 10427
0 10429 7 1 2 10425 10428
0 10430 7 1 2 10418 10429
0 10431 5 1 1 10430
0 10432 7 1 2 42324 10431
0 10433 5 1 1 10432
0 10434 7 4 2 48897 60739
0 10435 5 1 1 60857
0 10436 7 1 2 52846 56500
0 10437 5 1 1 10436
0 10438 7 1 2 488 53116
0 10439 5 1 1 10438
0 10440 7 1 2 47327 10439
0 10441 5 1 1 10440
0 10442 7 1 2 10437 10441
0 10443 5 1 1 10442
0 10444 7 1 2 60858 10443
0 10445 5 1 1 10444
0 10446 7 1 2 53949 58293
0 10447 7 1 2 60706 10446
0 10448 5 1 1 10447
0 10449 7 1 2 10445 10448
0 10450 5 1 1 10449
0 10451 7 3 2 49578 54472
0 10452 7 1 2 10450 60861
0 10453 5 1 1 10452
0 10454 7 1 2 10433 10453
0 10455 5 1 1 10454
0 10456 7 1 2 43524 10455
0 10457 5 1 1 10456
0 10458 7 1 2 60536 60707
0 10459 5 1 1 10458
0 10460 7 1 2 44925 2337
0 10461 5 1 1 10460
0 10462 7 1 2 53412 49098
0 10463 7 1 2 10461 10462
0 10464 5 1 1 10463
0 10465 7 1 2 10459 10464
0 10466 5 1 1 10465
0 10467 7 1 2 60862 10466
0 10468 5 1 1 10467
0 10469 7 1 2 47405 51171
0 10470 7 1 2 60854 10469
0 10471 5 1 1 10470
0 10472 7 1 2 58446 60863
0 10473 7 1 2 60708 10472
0 10474 5 1 1 10473
0 10475 7 1 2 10471 10474
0 10476 5 1 1 10475
0 10477 7 1 2 44495 10476
0 10478 5 1 1 10477
0 10479 7 1 2 10468 10478
0 10480 5 1 1 10479
0 10481 7 1 2 53950 10480
0 10482 5 1 1 10481
0 10483 7 1 2 57150 57498
0 10484 7 1 2 56418 10483
0 10485 5 1 1 10484
0 10486 7 1 2 10482 10485
0 10487 7 1 2 10457 10486
0 10488 5 1 1 10487
0 10489 7 1 2 48748 10488
0 10490 5 1 1 10489
0 10491 7 1 2 10368 10490
0 10492 7 1 2 10309 10491
0 10493 7 1 2 9949 10492
0 10494 5 1 1 10493
0 10495 7 1 2 46469 10494
0 10496 5 1 1 10495
0 10497 7 1 2 55408 57244
0 10498 7 1 2 55442 10497
0 10499 5 1 1 10498
0 10500 7 1 2 10496 10499
0 10501 5 1 1 10500
0 10502 7 1 2 57626 10501
0 10503 5 1 1 10502
0 10504 7 3 2 40786 42325
0 10505 5 3 1 60864
0 10506 7 1 2 56138 59648
0 10507 5 1 1 10506
0 10508 7 1 2 60867 10507
0 10509 5 2 1 10508
0 10510 7 1 2 43679 60870
0 10511 5 1 1 10510
0 10512 7 2 2 40787 48812
0 10513 5 2 1 60872
0 10514 7 1 2 10511 60874
0 10515 5 1 1 10514
0 10516 7 1 2 41454 10515
0 10517 5 1 1 10516
0 10518 7 3 2 45271 51157
0 10519 5 1 1 60876
0 10520 7 1 2 53312 60877
0 10521 5 1 1 10520
0 10522 7 1 2 10517 10521
0 10523 5 1 1 10522
0 10524 7 1 2 44496 10523
0 10525 5 1 1 10524
0 10526 7 6 2 41455 42089
0 10527 5 3 1 60879
0 10528 7 1 2 40788 60880
0 10529 7 1 2 52052 10528
0 10530 5 1 1 10529
0 10531 7 1 2 10525 10530
0 10532 5 1 1 10531
0 10533 7 1 2 44405 10532
0 10534 5 1 1 10533
0 10535 7 1 2 52372 51484
0 10536 7 1 2 58268 10535
0 10537 5 1 1 10536
0 10538 7 1 2 10534 10537
0 10539 5 1 1 10538
0 10540 7 1 2 42550 10539
0 10541 5 1 1 10540
0 10542 7 4 2 45877 54440
0 10543 7 1 2 50502 54908
0 10544 5 1 1 10543
0 10545 7 1 2 52376 3776
0 10546 5 2 1 10545
0 10547 7 1 2 49421 60892
0 10548 5 1 1 10547
0 10549 7 1 2 10544 10548
0 10550 5 1 1 10549
0 10551 7 1 2 60888 10550
0 10552 5 1 1 10551
0 10553 7 1 2 10541 10552
0 10554 5 1 1 10553
0 10555 7 1 2 43336 10554
0 10556 5 1 1 10555
0 10557 7 2 2 40789 54839
0 10558 7 1 2 58140 47200
0 10559 5 1 1 10558
0 10560 7 1 2 50926 10559
0 10561 5 1 1 10560
0 10562 7 1 2 60894 10561
0 10563 5 1 1 10562
0 10564 7 1 2 10556 10563
0 10565 5 1 1 10564
0 10566 7 1 2 43525 10565
0 10567 5 1 1 10566
0 10568 7 1 2 658 56314
0 10569 5 1 1 10568
0 10570 7 1 2 42090 10569
0 10571 5 1 1 10570
0 10572 7 1 2 56366 10571
0 10573 5 1 1 10572
0 10574 7 1 2 45878 10573
0 10575 5 1 1 10574
0 10576 7 1 2 49489 48629
0 10577 5 1 1 10576
0 10578 7 1 2 52350 10577
0 10579 5 2 1 10578
0 10580 7 1 2 41204 54430
0 10581 7 1 2 60896 10580
0 10582 5 1 1 10581
0 10583 7 1 2 10575 10582
0 10584 5 1 1 10583
0 10585 7 1 2 42326 10584
0 10586 5 1 1 10585
0 10587 7 5 2 42551 50477
0 10588 7 2 2 50890 60898
0 10589 5 1 1 60903
0 10590 7 2 2 47644 47163
0 10591 5 1 1 60905
0 10592 7 1 2 10591 51114
0 10593 5 1 1 10592
0 10594 7 1 2 55453 10593
0 10595 5 1 1 10594
0 10596 7 1 2 10589 10595
0 10597 5 1 1 10596
0 10598 7 1 2 49915 60904
0 10599 5 1 1 10598
0 10600 7 1 2 40369 10599
0 10601 5 1 1 10600
0 10602 7 1 2 43337 10601
0 10603 7 1 2 10597 10602
0 10604 5 1 1 10603
0 10605 7 1 2 55855 54892
0 10606 5 1 1 10605
0 10607 7 7 2 47406 51608
0 10608 5 1 1 60907
0 10609 7 1 2 51063 10608
0 10610 5 1 1 10609
0 10611 7 1 2 45879 10610
0 10612 5 1 1 10611
0 10613 7 2 2 42552 51853
0 10614 7 1 2 49490 60914
0 10615 5 1 1 10614
0 10616 7 1 2 10612 10615
0 10617 5 1 1 10616
0 10618 7 1 2 43877 10617
0 10619 5 1 1 10618
0 10620 7 1 2 10606 10619
0 10621 7 1 2 10604 10620
0 10622 7 1 2 10586 10621
0 10623 5 1 1 10622
0 10624 7 1 2 40790 10623
0 10625 5 1 1 10624
0 10626 7 2 2 45437 54497
0 10627 5 1 1 60916
0 10628 7 1 2 52586 58132
0 10629 5 1 1 10628
0 10630 7 1 2 10627 10629
0 10631 5 1 1 10630
0 10632 7 1 2 60564 10631
0 10633 5 1 1 10632
0 10634 7 1 2 49491 60917
0 10635 5 1 1 10634
0 10636 7 1 2 10633 10635
0 10637 5 1 1 10636
0 10638 7 1 2 56610 10637
0 10639 5 1 1 10638
0 10640 7 1 2 10625 10639
0 10641 5 1 1 10640
0 10642 7 1 2 44756 10641
0 10643 5 1 1 10642
0 10644 7 1 2 47083 6851
0 10645 5 1 1 10644
0 10646 7 1 2 48875 10645
0 10647 5 1 1 10646
0 10648 7 1 2 47914 10647
0 10649 5 1 1 10648
0 10650 7 1 2 54913 10649
0 10651 5 1 1 10650
0 10652 7 1 2 54840 10651
0 10653 5 1 1 10652
0 10654 7 1 2 57995 54540
0 10655 5 1 1 10654
0 10656 7 3 2 43338 52443
0 10657 7 4 2 44406 50430
0 10658 5 1 1 60921
0 10659 7 1 2 54963 60922
0 10660 7 1 2 60918 10659
0 10661 5 1 1 10660
0 10662 7 1 2 10655 10661
0 10663 7 1 2 10653 10662
0 10664 5 1 1 10663
0 10665 7 1 2 40791 10664
0 10666 5 1 1 10665
0 10667 7 1 2 10643 10666
0 10668 7 1 2 10567 10667
0 10669 5 1 1 10668
0 10670 7 1 2 54142 10669
0 10671 5 1 1 10670
0 10672 7 2 2 48663 55752
0 10673 7 1 2 52351 48787
0 10674 5 4 1 10673
0 10675 7 1 2 60925 60927
0 10676 5 1 1 10675
0 10677 7 2 2 60908 51415
0 10678 5 1 1 60931
0 10679 7 1 2 53453 60932
0 10680 5 1 1 10679
0 10681 7 1 2 10676 10680
0 10682 5 1 1 10681
0 10683 7 1 2 54143 10682
0 10684 5 1 1 10683
0 10685 7 1 2 41345 46881
0 10686 5 1 1 10685
0 10687 7 1 2 43526 10686
0 10688 5 1 1 10687
0 10689 7 1 2 48664 46928
0 10690 5 3 1 10689
0 10691 7 1 2 43339 60933
0 10692 5 2 1 10691
0 10693 7 1 2 49492 46910
0 10694 7 1 2 60500 10693
0 10695 7 2 2 60936 10694
0 10696 5 1 1 60938
0 10697 7 1 2 10688 60939
0 10698 5 4 1 10697
0 10699 7 2 2 57678 55330
0 10700 7 1 2 57157 60944
0 10701 7 1 2 60940 10700
0 10702 5 1 1 10701
0 10703 7 1 2 10684 10702
0 10704 5 1 1 10703
0 10705 7 1 2 45438 10704
0 10706 5 1 1 10705
0 10707 7 2 2 56702 53951
0 10708 7 1 2 54851 60946
0 10709 5 1 1 10708
0 10710 7 1 2 48665 57042
0 10711 5 1 1 10710
0 10712 7 5 2 44197 41205
0 10713 7 3 2 46378 58960
0 10714 7 1 2 60948 60953
0 10715 7 1 2 60897 10714
0 10716 5 1 1 10715
0 10717 7 1 2 10711 10716
0 10718 5 1 1 10717
0 10719 7 7 2 45880 49638
0 10720 5 1 1 60956
0 10721 7 1 2 42327 60957
0 10722 7 1 2 10718 10721
0 10723 5 1 1 10722
0 10724 7 1 2 10709 10723
0 10725 7 1 2 10706 10724
0 10726 5 1 1 10725
0 10727 7 1 2 44062 10726
0 10728 5 1 1 10727
0 10729 7 1 2 58170 1829
0 10730 5 2 1 10729
0 10731 7 1 2 43527 60963
0 10732 5 1 1 10731
0 10733 7 1 2 52444 55864
0 10734 5 2 1 10733
0 10735 7 1 2 10732 60965
0 10736 5 1 1 10735
0 10737 7 17 2 43680 40588
0 10738 7 4 2 60967 49729
0 10739 5 1 1 60984
0 10740 7 1 2 10739 434
0 10741 5 2 1 10740
0 10742 7 1 2 10736 60988
0 10743 5 1 1 10742
0 10744 7 2 2 48749 54407
0 10745 7 1 2 58472 60990
0 10746 5 1 1 10745
0 10747 7 2 2 48548 55856
0 10748 5 1 1 60992
0 10749 7 2 2 49493 51192
0 10750 5 1 1 60994
0 10751 7 1 2 54311 10750
0 10752 5 1 1 10751
0 10753 7 1 2 10748 10752
0 10754 5 1 1 10753
0 10755 7 1 2 42091 10754
0 10756 5 1 1 10755
0 10757 7 1 2 10746 10756
0 10758 5 1 1 10757
0 10759 7 1 2 40792 10758
0 10760 5 1 1 10759
0 10761 7 1 2 10743 10760
0 10762 5 1 1 10761
0 10763 7 1 2 43340 10762
0 10764 5 1 1 10763
0 10765 7 2 2 44757 51609
0 10766 5 1 1 60996
0 10767 7 1 2 60889 60997
0 10768 5 1 1 10767
0 10769 7 1 2 10764 10768
0 10770 5 1 1 10769
0 10771 7 1 2 46837 10770
0 10772 5 1 1 10771
0 10773 7 1 2 60503 60991
0 10774 5 1 1 10773
0 10775 7 1 2 54312 54814
0 10776 5 1 1 10775
0 10777 7 1 2 54038 49150
0 10778 5 1 1 10777
0 10779 7 2 2 43341 50117
0 10780 7 1 2 44758 60998
0 10781 5 1 1 10780
0 10782 7 1 2 10778 10781
0 10783 5 1 1 10782
0 10784 7 1 2 45881 10783
0 10785 5 1 1 10784
0 10786 7 1 2 10776 10785
0 10787 7 1 2 10774 10786
0 10788 5 1 1 10787
0 10789 7 1 2 46779 10788
0 10790 5 1 1 10789
0 10791 7 1 2 41346 46929
0 10792 5 3 1 10791
0 10793 7 1 2 43681 61000
0 10794 5 1 1 10793
0 10795 7 2 2 55887 47180
0 10796 5 1 1 61003
0 10797 7 1 2 10794 10796
0 10798 5 2 1 10797
0 10799 7 1 2 54408 52731
0 10800 7 1 2 61005 10799
0 10801 5 1 1 10800
0 10802 7 2 2 43528 51039
0 10803 5 1 1 61007
0 10804 7 1 2 49639 10803
0 10805 5 1 1 10804
0 10806 7 1 2 41347 50200
0 10807 5 2 1 10806
0 10808 7 1 2 9356 54389
0 10809 7 1 2 61009 10808
0 10810 7 1 2 10805 10809
0 10811 5 1 1 10810
0 10812 7 1 2 54541 55724
0 10813 5 1 1 10812
0 10814 7 2 2 43342 53207
0 10815 5 1 1 61011
0 10816 7 1 2 43878 61012
0 10817 5 1 1 10816
0 10818 7 1 2 10813 10817
0 10819 5 1 1 10818
0 10820 7 1 2 60934 10819
0 10821 5 1 1 10820
0 10822 7 3 2 44759 48750
0 10823 5 5 1 61013
0 10824 7 1 2 42553 54944
0 10825 7 1 2 61016 10824
0 10826 5 1 1 10825
0 10827 7 1 2 10821 10826
0 10828 7 1 2 10811 10827
0 10829 7 1 2 10801 10828
0 10830 7 1 2 10790 10829
0 10831 5 1 1 10830
0 10832 7 1 2 40793 10831
0 10833 5 1 1 10832
0 10834 7 1 2 46711 60964
0 10835 5 1 1 10834
0 10836 7 1 2 60966 10835
0 10837 5 1 1 10836
0 10838 7 1 2 43529 10837
0 10839 5 1 1 10838
0 10840 7 1 2 60899 47193
0 10841 5 1 1 10840
0 10842 7 1 2 10839 10841
0 10843 5 1 1 10842
0 10844 7 1 2 60989 10843
0 10845 5 1 1 10844
0 10846 7 1 2 10833 10845
0 10847 7 1 2 10772 10846
0 10848 5 1 1 10847
0 10849 7 1 2 53952 10848
0 10850 5 1 1 10849
0 10851 7 1 2 10728 10850
0 10852 7 1 2 10671 10851
0 10853 5 1 1 10852
0 10854 7 1 2 42800 10853
0 10855 5 1 1 10854
0 10856 7 4 2 53879 56675
0 10857 7 1 2 43530 51001
0 10858 7 1 2 10696 10857
0 10859 5 1 1 10858
0 10860 7 1 2 3225 10859
0 10861 5 1 1 10860
0 10862 7 1 2 42328 10861
0 10863 5 1 1 10862
0 10864 7 2 2 50823 48421
0 10865 5 1 1 61025
0 10866 7 1 2 39984 60501
0 10867 5 1 1 10866
0 10868 7 3 2 61001 10867
0 10869 5 1 1 61027
0 10870 7 1 2 43682 61028
0 10871 5 1 1 10870
0 10872 7 1 2 10865 10871
0 10873 7 1 2 10863 10872
0 10874 5 1 1 10873
0 10875 7 1 2 40794 52732
0 10876 7 1 2 10874 10875
0 10877 5 1 1 10876
0 10878 7 1 2 47875 50947
0 10879 7 1 2 61004 10878
0 10880 5 1 1 10879
0 10881 7 1 2 44063 50489
0 10882 5 1 1 10881
0 10883 7 1 2 51866 10882
0 10884 7 1 2 58141 10883
0 10885 7 1 2 46870 10884
0 10886 5 1 1 10885
0 10887 7 1 2 10880 10886
0 10888 7 1 2 10877 10887
0 10889 5 1 1 10888
0 10890 7 1 2 42554 10889
0 10891 5 1 1 10890
0 10892 7 2 2 44640 50696
0 10893 7 2 2 51918 61030
0 10894 5 1 1 61032
0 10895 7 1 2 52674 61033
0 10896 5 1 1 10895
0 10897 7 1 2 10891 10896
0 10898 5 1 1 10897
0 10899 7 1 2 49579 10898
0 10900 5 1 1 10899
0 10901 7 1 2 44641 46871
0 10902 5 2 1 10901
0 10903 7 1 2 43531 61029
0 10904 5 1 1 10903
0 10905 7 1 2 61034 10904
0 10906 5 1 1 10905
0 10907 7 1 2 43683 10906
0 10908 5 1 1 10907
0 10909 7 1 2 43532 61026
0 10910 5 2 1 10909
0 10911 7 1 2 10908 61036
0 10912 5 2 1 10911
0 10913 7 1 2 60881 61038
0 10914 5 2 1 10913
0 10915 7 1 2 52402 52556
0 10916 5 4 1 10915
0 10917 7 2 2 45272 61042
0 10918 5 1 1 61046
0 10919 7 1 2 10918 49422
0 10920 5 1 1 10919
0 10921 7 1 2 44760 10920
0 10922 5 1 1 10921
0 10923 7 2 2 45660 60941
0 10924 5 1 1 61048
0 10925 7 1 2 10922 10924
0 10926 5 1 1 10925
0 10927 7 1 2 43879 10926
0 10928 5 2 1 10927
0 10929 7 1 2 51252 56105
0 10930 5 2 1 10929
0 10931 7 1 2 49494 54910
0 10932 7 1 2 49303 10931
0 10933 5 2 1 10932
0 10934 7 1 2 44761 61054
0 10935 5 1 1 10934
0 10936 7 1 2 61052 10935
0 10937 5 1 1 10936
0 10938 7 1 2 45661 10937
0 10939 5 1 1 10938
0 10940 7 1 2 61050 10939
0 10941 5 1 1 10940
0 10942 7 1 2 45439 10941
0 10943 5 1 1 10942
0 10944 7 1 2 61040 10943
0 10945 5 1 1 10944
0 10946 7 1 2 42555 10945
0 10947 5 1 1 10946
0 10948 7 1 2 48549 61039
0 10949 5 1 1 10948
0 10950 7 1 2 49580 60434
0 10951 5 1 1 10950
0 10952 7 1 2 10949 10951
0 10953 5 1 1 10952
0 10954 7 1 2 52177 10953
0 10955 5 1 1 10954
0 10956 7 2 2 48751 58386
0 10957 7 1 2 58380 47171
0 10958 7 2 2 47206 10957
0 10959 5 1 1 61058
0 10960 7 1 2 47117 61059
0 10961 5 1 1 10960
0 10962 7 1 2 61056 10961
0 10963 5 1 1 10962
0 10964 7 1 2 49423 57583
0 10965 5 1 1 10964
0 10966 7 5 2 46712 54751
0 10967 5 1 1 61060
0 10968 7 1 2 49495 10967
0 10969 5 1 1 10968
0 10970 7 1 2 43343 10969
0 10971 5 2 1 10970
0 10972 7 1 2 10965 61065
0 10973 7 1 2 10963 10972
0 10974 5 1 1 10973
0 10975 7 1 2 54409 10974
0 10976 5 2 1 10975
0 10977 7 2 2 52074 49424
0 10978 5 2 1 61069
0 10979 7 1 2 42092 61071
0 10980 5 1 1 10979
0 10981 7 1 2 55632 10980
0 10982 5 1 1 10981
0 10983 7 1 2 41206 10982
0 10984 5 1 1 10983
0 10985 7 4 2 40370 42093
0 10986 5 2 1 61073
0 10987 7 1 2 41348 61074
0 10988 5 1 1 10987
0 10989 7 1 2 10984 10988
0 10990 5 1 1 10989
0 10991 7 1 2 42556 10990
0 10992 5 1 1 10991
0 10993 7 4 2 39985 54650
0 10994 7 2 2 50277 46890
0 10995 7 2 2 61079 61083
0 10996 7 1 2 41098 61085
0 10997 5 1 1 10996
0 10998 7 1 2 54819 10997
0 10999 5 1 1 10998
0 11000 7 1 2 10992 10999
0 11001 5 1 1 11000
0 11002 7 1 2 44762 11001
0 11003 5 1 1 11002
0 11004 7 1 2 55857 58318
0 11005 5 1 1 11004
0 11006 7 1 2 42557 57996
0 11007 7 1 2 50452 11006
0 11008 5 1 1 11007
0 11009 7 1 2 11005 11008
0 11010 7 1 2 11003 11009
0 11011 7 1 2 61067 11010
0 11012 5 1 1 11011
0 11013 7 1 2 42329 11012
0 11014 5 1 1 11013
0 11015 7 1 2 10955 11014
0 11016 7 1 2 10947 11015
0 11017 5 1 1 11016
0 11018 7 1 2 44064 11017
0 11019 5 1 1 11018
0 11020 7 1 2 10900 11019
0 11021 5 1 1 11020
0 11022 7 1 2 61021 11021
0 11023 5 1 1 11022
0 11024 7 1 2 10855 11023
0 11025 5 1 1 11024
0 11026 7 1 2 44926 11025
0 11027 5 1 1 11026
0 11028 7 1 2 50862 57865
0 11029 5 1 1 11028
0 11030 7 1 2 53953 58456
0 11031 5 1 1 11030
0 11032 7 1 2 11029 11031
0 11033 5 1 1 11032
0 11034 7 1 2 48752 11033
0 11035 5 1 1 11034
0 11036 7 1 2 42330 60856
0 11037 5 1 1 11036
0 11038 7 2 2 45440 53728
0 11039 5 2 1 61087
0 11040 7 1 2 54144 61089
0 11041 5 1 1 11040
0 11042 7 1 2 60617 11041
0 11043 5 1 1 11042
0 11044 7 1 2 49425 11043
0 11045 5 1 1 11044
0 11046 7 1 2 11037 11045
0 11047 7 1 2 11035 11046
0 11048 5 1 1 11047
0 11049 7 1 2 41625 11048
0 11050 5 1 1 11049
0 11051 7 8 2 46379 57833
0 11052 5 1 1 61091
0 11053 7 1 2 57077 11052
0 11054 5 3 1 11053
0 11055 7 1 2 41099 54024
0 11056 5 1 1 11055
0 11057 7 1 2 43344 11056
0 11058 7 1 2 61099 11057
0 11059 5 2 1 11058
0 11060 7 1 2 46838 57043
0 11061 5 2 1 11060
0 11062 7 1 2 61102 61104
0 11063 5 1 1 11062
0 11064 7 2 2 50159 53680
0 11065 5 1 1 61106
0 11066 7 1 2 11063 61107
0 11067 5 1 1 11066
0 11068 7 1 2 11050 11067
0 11069 5 1 1 11068
0 11070 7 1 2 44763 11069
0 11071 5 1 1 11070
0 11072 7 2 2 40950 48029
0 11073 7 1 2 58744 51040
0 11074 7 4 2 43345 41626
0 11075 7 1 2 54683 61110
0 11076 7 1 2 11073 11075
0 11077 7 1 2 61108 11076
0 11078 5 1 1 11077
0 11079 7 1 2 11071 11078
0 11080 5 1 1 11079
0 11081 7 1 2 46092 11080
0 11082 5 1 1 11081
0 11083 7 2 2 60573 60694
0 11084 5 1 1 61114
0 11085 7 2 2 45662 61115
0 11086 5 2 1 61116
0 11087 7 1 2 45441 61117
0 11088 5 1 1 11087
0 11089 7 1 2 11082 11088
0 11090 5 1 1 11089
0 11091 7 1 2 43880 11090
0 11092 5 1 1 11091
0 11093 7 1 2 58331 58421
0 11094 5 1 1 11093
0 11095 7 1 2 52752 11094
0 11096 5 1 1 11095
0 11097 7 1 2 44764 11096
0 11098 5 1 1 11097
0 11099 7 1 2 51661 58393
0 11100 5 1 1 11099
0 11101 7 1 2 41456 54117
0 11102 7 1 2 11100 11101
0 11103 5 1 1 11102
0 11104 7 1 2 11065 11103
0 11105 5 1 1 11104
0 11106 7 1 2 42801 11105
0 11107 5 1 1 11106
0 11108 7 1 2 11098 11107
0 11109 5 1 1 11108
0 11110 7 1 2 56780 11109
0 11111 5 1 1 11110
0 11112 7 1 2 11092 11111
0 11113 5 1 1 11112
0 11114 7 1 2 42558 11113
0 11115 5 1 1 11114
0 11116 7 1 2 49426 48338
0 11117 7 1 2 51283 11116
0 11118 5 1 1 11117
0 11119 7 2 2 41457 52308
0 11120 5 1 1 61120
0 11121 7 1 2 43684 11120
0 11122 5 1 1 11121
0 11123 7 1 2 54950 11122
0 11124 5 1 1 11123
0 11125 7 1 2 47532 47227
0 11126 7 1 2 11124 11125
0 11127 5 1 1 11126
0 11128 7 1 2 11118 11127
0 11129 5 1 1 11128
0 11130 7 1 2 51260 11129
0 11131 5 1 1 11130
0 11132 7 5 2 54964 61017
0 11133 5 3 1 61122
0 11134 7 1 2 42802 50262
0 11135 7 1 2 61127 11134
0 11136 5 1 1 11135
0 11137 7 1 2 11131 11136
0 11138 5 1 1 11137
0 11139 7 1 2 60711 11138
0 11140 5 1 1 11139
0 11141 7 1 2 11115 11140
0 11142 5 1 1 11141
0 11143 7 1 2 47723 11142
0 11144 5 1 1 11143
0 11145 7 1 2 41349 60654
0 11146 5 3 1 11145
0 11147 7 3 2 43346 44765
0 11148 7 1 2 53820 61133
0 11149 5 1 1 11148
0 11150 7 1 2 3427 11149
0 11151 5 1 1 11150
0 11152 7 1 2 43881 11151
0 11153 5 1 1 11152
0 11154 7 1 2 3497 11153
0 11155 5 2 1 11154
0 11156 7 1 2 61130 61136
0 11157 5 1 1 11156
0 11158 7 5 2 43882 49787
0 11159 7 1 2 53849 61138
0 11160 5 1 1 11159
0 11161 7 1 2 11157 11160
0 11162 5 1 1 11161
0 11163 7 1 2 43685 11162
0 11164 5 1 1 11163
0 11165 7 1 2 46713 54801
0 11166 7 1 2 54410 11165
0 11167 5 1 1 11166
0 11168 7 2 2 43883 54351
0 11169 5 3 1 61143
0 11170 7 1 2 55311 50971
0 11171 5 2 1 11170
0 11172 7 1 2 61145 61148
0 11173 7 1 2 11167 11172
0 11174 5 1 1 11173
0 11175 7 1 2 42803 11174
0 11176 5 1 1 11175
0 11177 7 3 2 43884 53087
0 11178 5 1 1 61150
0 11179 7 1 2 53850 61151
0 11180 7 1 2 48036 11179
0 11181 5 1 1 11180
0 11182 7 1 2 11176 11181
0 11183 7 1 2 11164 11182
0 11184 5 1 1 11183
0 11185 7 1 2 53954 11184
0 11186 5 1 1 11185
0 11187 7 1 2 54083 51350
0 11188 7 1 2 55836 11187
0 11189 5 1 1 11188
0 11190 7 1 2 11186 11189
0 11191 5 1 1 11190
0 11192 7 1 2 42331 11191
0 11193 5 1 1 11192
0 11194 7 4 2 43885 45046
0 11195 7 4 2 44198 44766
0 11196 7 5 2 61153 61157
0 11197 7 3 2 42559 56783
0 11198 7 1 2 48813 61166
0 11199 7 1 2 61161 11198
0 11200 5 1 1 11199
0 11201 7 2 2 52022 53955
0 11202 5 1 1 61169
0 11203 7 1 2 54411 47956
0 11204 7 1 2 61170 11203
0 11205 5 1 1 11204
0 11206 7 1 2 11200 11205
0 11207 5 1 1 11206
0 11208 7 1 2 43347 11207
0 11209 5 1 1 11208
0 11210 7 1 2 59079 50613
0 11211 7 2 2 55341 11210
0 11212 7 1 2 56676 61171
0 11213 5 1 1 11212
0 11214 7 1 2 11209 11213
0 11215 5 1 1 11214
0 11216 7 1 2 43686 11215
0 11217 5 1 1 11216
0 11218 7 1 2 54390 52314
0 11219 5 1 1 11218
0 11220 7 3 2 44642 53186
0 11221 5 1 1 61173
0 11222 7 1 2 42560 61174
0 11223 5 1 1 11222
0 11224 7 1 2 11219 11223
0 11225 5 1 1 11224
0 11226 7 1 2 47957 60735
0 11227 7 1 2 11225 11226
0 11228 5 1 1 11227
0 11229 7 1 2 11217 11228
0 11230 5 1 1 11229
0 11231 7 1 2 46839 11230
0 11232 5 1 1 11231
0 11233 7 1 2 49427 61137
0 11234 5 1 1 11233
0 11235 7 5 2 44767 55236
0 11236 7 1 2 43886 61176
0 11237 5 1 1 11236
0 11238 7 1 2 11234 11237
0 11239 5 1 1 11238
0 11240 7 2 2 59929 53164
0 11241 7 1 2 58924 61181
0 11242 7 1 2 11239 11241
0 11243 5 1 1 11242
0 11244 7 1 2 11232 11243
0 11245 7 1 2 11193 11244
0 11246 5 1 1 11245
0 11247 7 1 2 41627 11246
0 11248 5 1 1 11247
0 11249 7 1 2 11144 11248
0 11250 5 1 1 11249
0 11251 7 1 2 44065 11250
0 11252 5 1 1 11251
0 11253 7 2 2 48313 54724
0 11254 7 1 2 61183 56471
0 11255 5 1 1 11254
0 11256 7 1 2 2959 54464
0 11257 5 1 1 11256
0 11258 7 1 2 49744 11257
0 11259 5 1 1 11258
0 11260 7 1 2 11255 11259
0 11261 5 1 1 11260
0 11262 7 1 2 48753 11261
0 11263 5 1 1 11262
0 11264 7 4 2 44643 53821
0 11265 7 7 2 43687 44066
0 11266 7 3 2 49581 61189
0 11267 7 1 2 61185 61196
0 11268 5 1 1 11267
0 11269 7 1 2 11263 11268
0 11270 5 1 1 11269
0 11271 7 1 2 42332 11270
0 11272 5 1 1 11271
0 11273 7 1 2 49428 57932
0 11274 5 1 1 11273
0 11275 7 1 2 57935 11274
0 11276 5 1 1 11275
0 11277 7 1 2 52525 49745
0 11278 7 1 2 11276 11277
0 11279 5 1 1 11278
0 11280 7 1 2 11272 11279
0 11281 5 1 1 11280
0 11282 7 1 2 53956 11281
0 11283 5 1 1 11282
0 11284 7 1 2 55389 50381
0 11285 5 1 1 11284
0 11286 7 1 2 3855 11285
0 11287 5 1 1 11286
0 11288 7 1 2 53957 11287
0 11289 5 1 1 11288
0 11290 7 2 2 46380 47915
0 11291 7 1 2 48898 55390
0 11292 7 1 2 61199 11291
0 11293 5 1 1 11292
0 11294 7 1 2 11289 11293
0 11295 5 1 1 11294
0 11296 7 1 2 44067 11295
0 11297 5 1 1 11296
0 11298 7 2 2 41751 55817
0 11299 7 1 2 57028 54456
0 11300 7 1 2 61201 11299
0 11301 5 1 1 11300
0 11302 7 1 2 11297 11301
0 11303 5 1 1 11302
0 11304 7 1 2 52053 11303
0 11305 5 1 1 11304
0 11306 7 1 2 57107 60585
0 11307 5 1 1 11306
0 11308 7 1 2 11305 11307
0 11309 5 1 1 11308
0 11310 7 1 2 42094 11309
0 11311 5 1 1 11310
0 11312 7 2 2 58852 52884
0 11313 7 1 2 61167 61197
0 11314 7 1 2 61203 11313
0 11315 5 1 1 11314
0 11316 7 1 2 11311 11315
0 11317 7 1 2 11283 11316
0 11318 5 1 1 11317
0 11319 7 1 2 41628 11318
0 11320 5 1 1 11319
0 11321 7 1 2 52445 50873
0 11322 7 3 2 44407 44768
0 11323 7 1 2 61205 58303
0 11324 7 1 2 11321 11323
0 11325 7 2 2 49429 54725
0 11326 7 1 2 57044 61208
0 11327 7 1 2 11324 11326
0 11328 5 1 1 11327
0 11329 7 1 2 11320 11328
0 11330 5 1 1 11329
0 11331 7 1 2 47645 11330
0 11332 5 1 1 11331
0 11333 7 5 2 43688 45882
0 11334 7 2 2 48814 61210
0 11335 5 1 1 61215
0 11336 7 1 2 54509 11335
0 11337 5 1 1 11336
0 11338 7 1 2 47724 54118
0 11339 7 1 2 11337 11338
0 11340 5 1 1 11339
0 11341 7 1 2 60483 11340
0 11342 5 1 1 11341
0 11343 7 1 2 51660 11342
0 11344 5 1 1 11343
0 11345 7 5 2 44644 45442
0 11346 7 2 2 45663 61217
0 11347 5 1 1 61222
0 11348 7 1 2 11347 60868
0 11349 5 1 1 11348
0 11350 7 1 2 43689 11349
0 11351 5 1 1 11350
0 11352 7 1 2 60875 11351
0 11353 5 1 1 11352
0 11354 7 1 2 47725 11353
0 11355 5 1 1 11354
0 11356 7 1 2 40795 48868
0 11357 5 1 1 11356
0 11358 7 1 2 11355 11357
0 11359 5 1 1 11358
0 11360 7 1 2 42561 11359
0 11361 5 1 1 11360
0 11362 7 1 2 11344 11361
0 11363 5 1 1 11362
0 11364 7 1 2 43090 56369
0 11365 7 1 2 56155 11364
0 11366 7 1 2 11363 11365
0 11367 5 1 1 11366
0 11368 7 1 2 11332 11367
0 11369 7 1 2 11252 11368
0 11370 7 1 2 11027 11369
0 11371 5 1 1 11370
0 11372 7 1 2 59441 11371
0 11373 5 1 1 11372
0 11374 7 1 2 10503 11373
0 11375 5 1 1 11374
0 11376 7 1 2 46243 11375
0 11377 5 1 1 11376
0 11378 7 1 2 47646 58439
0 11379 5 3 1 11378
0 11380 7 1 2 48754 59907
0 11381 5 1 1 11380
0 11382 7 1 2 49496 51383
0 11383 7 1 2 60442 11382
0 11384 7 1 2 11381 11383
0 11385 7 1 2 61224 11384
0 11386 5 1 1 11385
0 11387 7 1 2 44769 11386
0 11388 5 1 1 11387
0 11389 7 1 2 51764 2796
0 11390 5 2 1 11389
0 11391 7 1 2 42333 61227
0 11392 5 1 1 11391
0 11393 7 2 2 47407 48795
0 11394 5 2 1 61229
0 11395 7 1 2 52054 61230
0 11396 5 1 1 11395
0 11397 7 2 2 42095 54119
0 11398 7 1 2 58818 58398
0 11399 5 1 1 11398
0 11400 7 1 2 61233 11399
0 11401 7 1 2 60427 11400
0 11402 5 1 1 11401
0 11403 7 1 2 11396 11402
0 11404 7 1 2 11392 11403
0 11405 7 1 2 11388 11404
0 11406 5 1 1 11405
0 11407 7 1 2 45883 11406
0 11408 5 1 1 11407
0 11409 7 2 2 42562 58260
0 11410 5 1 1 61235
0 11411 7 1 2 44770 61236
0 11412 5 1 1 11411
0 11413 7 1 2 44771 52023
0 11414 5 4 1 11413
0 11415 7 1 2 49860 61237
0 11416 5 1 1 11415
0 11417 7 1 2 52304 11416
0 11418 5 1 1 11417
0 11419 7 1 2 49824 52024
0 11420 5 1 1 11419
0 11421 7 1 2 11418 11420
0 11422 5 1 1 11421
0 11423 7 1 2 45884 11422
0 11424 5 1 1 11423
0 11425 7 1 2 2426 11424
0 11426 5 1 1 11425
0 11427 7 1 2 50453 11426
0 11428 5 1 1 11427
0 11429 7 1 2 11412 11428
0 11430 7 1 2 11408 11429
0 11431 5 1 1 11430
0 11432 7 1 2 59442 11431
0 11433 5 1 1 11432
0 11434 7 1 2 56318 51110
0 11435 5 1 1 11434
0 11436 7 1 2 44645 11435
0 11437 5 1 1 11436
0 11438 7 1 2 48023 52802
0 11439 5 1 1 11438
0 11440 7 1 2 11437 11439
0 11441 5 1 1 11440
0 11442 7 1 2 43690 11441
0 11443 5 1 1 11442
0 11444 7 1 2 48042 11443
0 11445 5 2 1 11444
0 11446 7 1 2 45885 61241
0 11447 5 1 1 11446
0 11448 7 1 2 45886 56323
0 11449 7 1 2 53739 11448
0 11450 5 1 1 11449
0 11451 7 1 2 44772 11450
0 11452 5 1 1 11451
0 11453 7 1 2 11447 11452
0 11454 5 1 1 11453
0 11455 7 2 2 60565 54914
0 11456 5 1 1 61243
0 11457 7 1 2 39986 61244
0 11458 5 1 1 11457
0 11459 7 1 2 47042 58264
0 11460 5 1 1 11459
0 11461 7 1 2 60541 11460
0 11462 5 1 1 11461
0 11463 7 1 2 54120 11462
0 11464 7 2 2 11458 11463
0 11465 7 1 2 42563 61245
0 11466 5 1 1 11465
0 11467 7 1 2 60254 11466
0 11468 7 1 2 11454 11467
0 11469 5 1 1 11468
0 11470 7 1 2 11433 11469
0 11471 5 1 1 11470
0 11472 7 1 2 43887 11471
0 11473 5 1 1 11472
0 11474 7 4 2 43691 40992
0 11475 7 2 2 60394 61247
0 11476 5 3 1 61251
0 11477 7 3 2 41935 46619
0 11478 7 3 2 43180 61256
0 11479 5 3 1 61259
0 11480 7 1 2 60255 59326
0 11481 5 1 1 11480
0 11482 7 1 2 61262 11481
0 11483 5 1 1 11482
0 11484 7 1 2 48369 11483
0 11485 5 1 1 11484
0 11486 7 1 2 61253 11485
0 11487 5 1 1 11486
0 11488 7 1 2 43348 11487
0 11489 5 1 1 11488
0 11490 7 3 2 43533 60448
0 11491 5 1 1 61265
0 11492 7 1 2 43692 61266
0 11493 5 1 1 11492
0 11494 7 1 2 11489 11493
0 11495 5 1 1 11494
0 11496 7 1 2 48004 11495
0 11497 5 1 1 11496
0 11498 7 4 2 60320 59023
0 11499 5 1 1 61268
0 11500 7 1 2 61269 54772
0 11501 5 1 1 11500
0 11502 7 1 2 47084 61267
0 11503 5 1 1 11502
0 11504 7 1 2 11501 11503
0 11505 5 1 1 11504
0 11506 7 1 2 44646 11505
0 11507 5 1 1 11506
0 11508 7 2 2 44497 54802
0 11509 5 1 1 61272
0 11510 7 2 2 43693 52258
0 11511 5 1 1 61274
0 11512 7 1 2 11509 11511
0 11513 5 1 1 11512
0 11514 7 1 2 59443 11513
0 11515 5 1 1 11514
0 11516 7 3 2 43694 50874
0 11517 5 1 1 61276
0 11518 7 1 2 54767 11517
0 11519 5 1 1 11518
0 11520 7 17 2 44239 60321
0 11521 7 1 2 51576 61279
0 11522 7 1 2 11519 11521
0 11523 5 1 1 11522
0 11524 7 1 2 11515 11523
0 11525 5 1 1 11524
0 11526 7 1 2 43349 11525
0 11527 5 1 1 11526
0 11528 7 2 2 48755 59444
0 11529 7 1 2 49319 61296
0 11530 5 1 1 11529
0 11531 7 3 2 44240 44408
0 11532 7 2 2 43695 61298
0 11533 7 1 2 51315 60322
0 11534 7 1 2 61301 11533
0 11535 5 1 1 11534
0 11536 7 1 2 11530 11535
0 11537 5 1 1 11536
0 11538 7 1 2 43350 11537
0 11539 5 1 1 11538
0 11540 7 1 2 49430 60449
0 11541 5 1 1 11540
0 11542 7 1 2 11539 11541
0 11543 5 1 1 11542
0 11544 7 1 2 47043 11543
0 11545 5 1 1 11544
0 11546 7 1 2 11527 11545
0 11547 7 1 2 11507 11546
0 11548 7 1 2 11497 11547
0 11549 5 1 1 11548
0 11550 7 1 2 42334 11549
0 11551 5 1 1 11550
0 11552 7 1 2 46714 50362
0 11553 5 1 1 11552
0 11554 7 1 2 44647 46780
0 11555 5 1 1 11554
0 11556 7 1 2 40191 11555
0 11557 5 1 1 11556
0 11558 7 2 2 61002 11557
0 11559 7 1 2 43696 61303
0 11560 5 1 1 11559
0 11561 7 1 2 11553 11560
0 11562 5 1 1 11561
0 11563 7 1 2 43351 11562
0 11564 5 1 1 11563
0 11565 7 1 2 50984 11564
0 11566 5 1 1 11565
0 11567 7 1 2 59445 11566
0 11568 5 1 1 11567
0 11569 7 2 2 41936 49799
0 11570 7 2 2 44241 47181
0 11571 7 1 2 60323 53681
0 11572 7 1 2 61307 11571
0 11573 7 1 2 61305 11572
0 11574 5 1 1 11573
0 11575 7 1 2 11568 11574
0 11576 5 1 1 11575
0 11577 7 1 2 42096 11576
0 11578 5 1 1 11577
0 11579 7 1 2 52037 58199
0 11580 5 2 1 11579
0 11581 7 1 2 48815 53177
0 11582 5 1 1 11581
0 11583 7 1 2 61309 11582
0 11584 5 1 1 11583
0 11585 7 1 2 59446 11584
0 11586 5 1 1 11585
0 11587 7 7 2 42335 43181
0 11588 7 4 2 46620 61311
0 11589 5 3 1 61318
0 11590 7 4 2 45664 46470
0 11591 7 5 2 57627 61325
0 11592 5 3 1 61329
0 11593 7 1 2 43352 54803
0 11594 7 1 2 61330 11593
0 11595 5 1 1 11594
0 11596 7 1 2 61322 11595
0 11597 5 1 1 11596
0 11598 7 1 2 44498 11597
0 11599 5 1 1 11598
0 11600 7 3 2 42097 43182
0 11601 7 2 2 46621 61337
0 11602 5 3 1 61340
0 11603 7 1 2 52025 61341
0 11604 5 1 1 11603
0 11605 7 1 2 11599 11604
0 11606 5 1 1 11605
0 11607 7 1 2 49800 11606
0 11608 5 1 1 11607
0 11609 7 1 2 11586 11608
0 11610 5 1 1 11609
0 11611 7 1 2 46840 11610
0 11612 5 1 1 11611
0 11613 7 1 2 11578 11612
0 11614 7 1 2 11551 11613
0 11615 5 1 1 11614
0 11616 7 1 2 54352 11615
0 11617 5 1 1 11616
0 11618 7 2 2 50835 55861
0 11619 5 1 1 61345
0 11620 7 1 2 11619 61149
0 11621 5 1 1 11620
0 11622 7 1 2 51041 11621
0 11623 5 1 1 11622
0 11624 7 1 2 55858 53088
0 11625 7 1 2 60039 11624
0 11626 5 1 1 11625
0 11627 7 1 2 11623 11626
0 11628 5 1 1 11627
0 11629 7 1 2 59447 11628
0 11630 5 1 1 11629
0 11631 7 1 2 11617 11630
0 11632 7 1 2 11473 11631
0 11633 5 1 1 11632
0 11634 7 1 2 46381 11633
0 11635 5 1 1 11634
0 11636 7 1 2 61072 50509
0 11637 5 1 1 11636
0 11638 7 3 2 48756 50498
0 11639 5 1 1 61347
0 11640 7 1 2 11637 61348
0 11641 5 1 1 11640
0 11642 7 1 2 42564 11641
0 11643 5 2 1 11642
0 11644 7 1 2 45887 52055
0 11645 5 2 1 11644
0 11646 7 1 2 61350 61352
0 11647 5 1 1 11646
0 11648 7 5 2 55041 57193
0 11649 7 1 2 49582 61354
0 11650 7 1 2 11647 11649
0 11651 5 1 1 11650
0 11652 7 1 2 11635 11651
0 11653 5 1 1 11652
0 11654 7 1 2 44068 11653
0 11655 5 1 1 11654
0 11656 7 1 2 61263 11499
0 11657 5 2 1 11656
0 11658 7 1 2 52026 61359
0 11659 5 1 1 11658
0 11660 7 2 2 48816 61280
0 11661 5 1 1 61361
0 11662 7 1 2 11659 11661
0 11663 5 1 1 11662
0 11664 7 1 2 47408 11663
0 11665 5 1 1 11664
0 11666 7 1 2 48817 59448
0 11667 5 1 1 11666
0 11668 7 1 2 61252 60181
0 11669 5 1 1 11668
0 11670 7 1 2 11667 11669
0 11671 7 1 2 11665 11670
0 11672 5 1 1 11671
0 11673 7 1 2 47726 11672
0 11674 5 1 1 11673
0 11675 7 1 2 51823 61360
0 11676 5 1 1 11675
0 11677 7 1 2 61254 11676
0 11678 5 1 1 11677
0 11679 7 1 2 48818 11678
0 11680 5 1 1 11679
0 11681 7 1 2 52038 60450
0 11682 7 1 2 53396 11681
0 11683 5 1 1 11682
0 11684 7 1 2 11680 11683
0 11685 7 1 2 11674 11684
0 11686 5 1 1 11685
0 11687 7 1 2 42098 11686
0 11688 5 1 1 11687
0 11689 7 1 2 55138 60256
0 11690 5 1 1 11689
0 11691 7 1 2 59494 11690
0 11692 5 1 1 11691
0 11693 7 1 2 51201 11692
0 11694 5 1 1 11693
0 11695 7 1 2 60451 52723
0 11696 5 1 1 11695
0 11697 7 5 2 45085 41937
0 11698 7 4 2 44242 61363
0 11699 7 1 2 46471 51185
0 11700 7 1 2 61368 11699
0 11701 5 1 1 11700
0 11702 7 1 2 11696 11701
0 11703 7 1 2 11694 11702
0 11704 5 1 1 11703
0 11705 7 1 2 49431 11704
0 11706 5 1 1 11705
0 11707 7 1 2 58523 61297
0 11708 5 1 1 11707
0 11709 7 1 2 11706 11708
0 11710 5 1 1 11709
0 11711 7 1 2 47328 11710
0 11712 5 1 1 11711
0 11713 7 1 2 44648 61281
0 11714 5 1 1 11713
0 11715 7 1 2 61264 11714
0 11716 5 1 1 11715
0 11717 7 1 2 53589 11716
0 11718 5 1 1 11717
0 11719 7 1 2 51577 60452
0 11720 5 1 1 11719
0 11721 7 1 2 11718 11720
0 11722 5 1 1 11721
0 11723 7 1 2 43697 11722
0 11724 5 1 1 11723
0 11725 7 2 2 55888 59449
0 11726 5 1 1 61372
0 11727 7 1 2 11724 11726
0 11728 5 1 1 11727
0 11729 7 3 2 40371 53587
0 11730 5 3 1 61374
0 11731 7 1 2 42336 61377
0 11732 7 1 2 11728 11731
0 11733 5 1 1 11732
0 11734 7 1 2 11712 11733
0 11735 7 1 2 11688 11734
0 11736 5 1 1 11735
0 11737 7 1 2 54498 11736
0 11738 5 1 1 11737
0 11739 7 2 2 42337 52675
0 11740 5 1 1 61380
0 11741 7 1 2 52178 61373
0 11742 7 1 2 61381 11741
0 11743 5 1 1 11742
0 11744 7 1 2 11738 11743
0 11745 5 1 1 11744
0 11746 7 1 2 57003 11745
0 11747 5 1 1 11746
0 11748 7 1 2 42962 11747
0 11749 7 1 2 11655 11748
0 11750 5 1 1 11749
0 11751 7 1 2 47009 61238
0 11752 5 1 1 11751
0 11753 7 1 2 52305 11752
0 11754 5 1 1 11753
0 11755 7 1 2 40372 11754
0 11756 5 1 1 11755
0 11757 7 1 2 41458 58193
0 11758 5 1 1 11757
0 11759 7 1 2 11756 11758
0 11760 5 1 1 11759
0 11761 7 1 2 40589 11760
0 11762 5 1 1 11761
0 11763 7 2 2 50278 50416
0 11764 7 1 2 53250 61382
0 11765 5 1 1 11764
0 11766 7 1 2 11762 11765
0 11767 5 1 1 11766
0 11768 7 1 2 54499 11767
0 11769 5 1 1 11768
0 11770 7 1 2 45443 57886
0 11771 7 1 2 60928 11770
0 11772 5 1 1 11771
0 11773 7 2 2 48024 59656
0 11774 5 1 1 61384
0 11775 7 1 2 41207 57936
0 11776 7 1 2 61385 11775
0 11777 5 1 1 11776
0 11778 7 1 2 11772 11777
0 11779 5 1 1 11778
0 11780 7 1 2 41350 11779
0 11781 5 1 1 11780
0 11782 7 3 2 49640 48630
0 11783 7 3 2 40796 42099
0 11784 7 1 2 56541 61389
0 11785 7 1 2 61386 11784
0 11786 5 1 1 11785
0 11787 7 1 2 11781 11786
0 11788 5 1 1 11787
0 11789 7 1 2 40373 11788
0 11790 5 1 1 11789
0 11791 7 3 2 50478 60909
0 11792 5 1 1 61392
0 11793 7 1 2 45273 61393
0 11794 5 1 1 11793
0 11795 7 2 2 40374 198
0 11796 5 3 1 61395
0 11797 7 1 2 41351 61396
0 11798 5 1 1 11797
0 11799 7 1 2 42100 11798
0 11800 5 1 1 11799
0 11801 7 2 2 47329 51610
0 11802 5 3 1 61400
0 11803 7 1 2 41938 61401
0 11804 5 1 1 11803
0 11805 7 2 2 51591 11804
0 11806 7 4 2 47893 49315
0 11807 5 2 1 61407
0 11808 7 4 2 40375 54845
0 11809 7 1 2 61408 61413
0 11810 5 1 1 11809
0 11811 7 1 2 42338 11810
0 11812 5 1 1 11811
0 11813 7 1 2 61405 11812
0 11814 7 1 2 11800 11813
0 11815 5 1 1 11814
0 11816 7 1 2 40590 11815
0 11817 5 1 1 11816
0 11818 7 1 2 11794 11817
0 11819 5 1 1 11818
0 11820 7 1 2 41459 11819
0 11821 5 1 1 11820
0 11822 7 1 2 58006 59649
0 11823 5 1 1 11822
0 11824 7 12 2 42339 49641
0 11825 5 1 1 61417
0 11826 7 1 2 53555 61418
0 11827 7 1 2 52997 11826
0 11828 5 1 1 11827
0 11829 7 1 2 11823 11828
0 11830 7 1 2 11821 11829
0 11831 5 1 1 11830
0 11832 7 1 2 40797 11831
0 11833 5 1 1 11832
0 11834 7 1 2 11790 11833
0 11835 5 1 1 11834
0 11836 7 1 2 45888 11835
0 11837 5 1 1 11836
0 11838 7 1 2 11769 11837
0 11839 5 1 1 11838
0 11840 7 1 2 59136 11839
0 11841 5 1 1 11840
0 11842 7 1 2 53473 60942
0 11843 5 1 1 11842
0 11844 7 1 2 42565 58269
0 11845 5 1 1 11844
0 11846 7 1 2 40591 8724
0 11847 7 1 2 11845 11846
0 11848 5 1 1 11847
0 11849 7 1 2 11843 11848
0 11850 5 1 1 11849
0 11851 7 1 2 41460 11850
0 11852 5 1 1 11851
0 11853 7 1 2 58007 53474
0 11854 5 1 1 11853
0 11855 7 1 2 11852 11854
0 11856 5 1 1 11855
0 11857 7 7 2 40993 59948
0 11858 5 2 1 61429
0 11859 7 1 2 40798 61430
0 11860 7 1 2 11856 11859
0 11861 5 1 1 11860
0 11862 7 1 2 11841 11861
0 11863 5 1 1 11862
0 11864 7 1 2 43183 11863
0 11865 5 1 1 11864
0 11866 7 2 2 48666 57581
0 11867 5 1 1 61438
0 11868 7 3 2 41208 50279
0 11869 5 3 1 61440
0 11870 7 3 2 55446 61443
0 11871 5 2 1 61446
0 11872 7 1 2 52064 54902
0 11873 5 1 1 11872
0 11874 7 2 2 61447 11873
0 11875 5 1 1 61451
0 11876 7 1 2 41461 11875
0 11877 5 1 1 11876
0 11878 7 1 2 11867 11877
0 11879 5 1 1 11878
0 11880 7 1 2 40592 11879
0 11881 5 1 1 11880
0 11882 7 3 2 52393 50182
0 11883 7 1 2 41462 61453
0 11884 7 1 2 59864 11883
0 11885 5 1 1 11884
0 11886 7 1 2 11881 11885
0 11887 5 1 1 11886
0 11888 7 2 2 59420 60324
0 11889 7 1 2 60337 61456
0 11890 7 1 2 11887 11889
0 11891 5 1 1 11890
0 11892 7 1 2 46244 11891
0 11893 7 1 2 11865 11892
0 11894 5 1 1 11893
0 11895 7 1 2 49019 11894
0 11896 7 1 2 11750 11895
0 11897 5 1 1 11896
0 11898 7 1 2 51091 3262
0 11899 5 1 1 11898
0 11900 7 1 2 42340 11899
0 11901 5 1 1 11900
0 11902 7 2 2 54895 11901
0 11903 7 1 2 49497 51844
0 11904 5 2 1 11903
0 11905 7 1 2 58388 61460
0 11906 5 1 1 11905
0 11907 7 1 2 49432 51074
0 11908 5 2 1 11907
0 11909 7 2 2 11906 61462
0 11910 5 1 1 61464
0 11911 7 2 2 44409 11910
0 11912 5 1 1 61466
0 11913 7 1 2 51845 50927
0 11914 5 1 1 11913
0 11915 7 1 2 41939 58270
0 11916 7 2 2 11914 11915
0 11917 5 2 1 61468
0 11918 7 1 2 11912 61470
0 11919 5 1 1 11918
0 11920 7 1 2 43353 11919
0 11921 5 1 1 11920
0 11922 7 1 2 61458 11921
0 11923 5 1 1 11922
0 11924 7 1 2 41463 11923
0 11925 5 1 1 11924
0 11926 7 1 2 43888 51611
0 11927 5 2 1 11926
0 11928 7 1 2 50985 61472
0 11929 5 2 1 11928
0 11930 7 1 2 50479 54718
0 11931 7 1 2 61474 11930
0 11932 5 1 1 11931
0 11933 7 1 2 11925 11932
0 11934 5 1 1 11933
0 11935 7 1 2 42566 11934
0 11936 5 1 1 11935
0 11937 7 1 2 47897 54762
0 11938 5 1 1 11937
0 11939 7 3 2 53178 11938
0 11940 7 1 2 52056 61476
0 11941 5 2 1 11940
0 11942 7 3 2 47898 58239
0 11943 5 2 1 61481
0 11944 7 1 2 61484 50921
0 11945 5 1 1 11944
0 11946 7 1 2 61479 11945
0 11947 5 2 1 11946
0 11948 7 2 2 45889 61486
0 11949 7 1 2 43889 61488
0 11950 5 1 1 11949
0 11951 7 1 2 45444 60910
0 11952 5 1 1 11951
0 11953 7 1 2 856 11952
0 11954 5 1 1 11953
0 11955 7 1 2 45665 11954
0 11956 5 1 1 11955
0 11957 7 4 2 41209 51042
0 11958 5 3 1 61490
0 11959 7 1 2 51164 61494
0 11960 5 4 1 11959
0 11961 7 1 2 59657 61497
0 11962 5 2 1 11961
0 11963 7 1 2 11956 61501
0 11964 5 1 1 11963
0 11965 7 1 2 45274 11964
0 11966 5 1 1 11965
0 11967 7 1 2 43890 11639
0 11968 5 1 1 11967
0 11969 7 1 2 42567 11968
0 11970 7 1 2 11966 11969
0 11971 5 1 1 11970
0 11972 7 1 2 47253 52310
0 11973 5 1 1 11972
0 11974 7 1 2 40593 52046
0 11975 5 2 1 11974
0 11976 7 1 2 53179 61503
0 11977 5 1 1 11976
0 11978 7 1 2 43891 54121
0 11979 5 1 1 11978
0 11980 7 2 2 50928 11979
0 11981 7 1 2 11977 61505
0 11982 5 1 1 11981
0 11983 7 1 2 47916 11982
0 11984 5 1 1 11983
0 11985 7 2 2 11973 11984
0 11986 7 1 2 40594 52248
0 11987 5 2 1 11986
0 11988 7 1 2 43534 61509
0 11989 5 2 1 11988
0 11990 7 1 2 43892 51676
0 11991 5 1 1 11990
0 11992 7 1 2 61511 11991
0 11993 5 1 1 11992
0 11994 7 1 2 52027 11993
0 11995 5 1 1 11994
0 11996 7 1 2 45890 4964
0 11997 7 1 2 11995 11996
0 11998 7 1 2 61507 11997
0 11999 5 1 1 11998
0 12000 7 1 2 44773 11999
0 12001 7 1 2 11971 12000
0 12002 5 1 1 12001
0 12003 7 1 2 11950 12002
0 12004 7 1 2 11936 12003
0 12005 5 2 1 12004
0 12006 7 1 2 54145 61513
0 12007 5 1 1 12006
0 12008 7 1 2 49498 58400
0 12009 5 1 1 12008
0 12010 7 1 2 61014 12009
0 12011 5 1 1 12010
0 12012 7 1 2 61053 12011
0 12013 5 1 1 12012
0 12014 7 1 2 43893 12013
0 12015 5 1 1 12014
0 12016 7 2 2 43698 51253
0 12017 7 1 2 49788 61515
0 12018 5 1 1 12017
0 12019 7 1 2 12015 12018
0 12020 5 1 1 12019
0 12021 7 1 2 45891 12020
0 12022 5 1 1 12021
0 12023 7 1 2 52446 50545
0 12024 5 1 1 12023
0 12025 7 1 2 12022 12024
0 12026 5 1 1 12025
0 12027 7 1 2 53958 12026
0 12028 5 1 1 12027
0 12029 7 1 2 12007 12028
0 12030 5 1 1 12029
0 12031 7 1 2 59450 12030
0 12032 5 1 1 12031
0 12033 7 6 2 40595 46382
0 12034 7 4 2 44199 41464
0 12035 7 2 2 45047 61523
0 12036 7 3 2 61517 61527
0 12037 5 1 1 61529
0 12038 7 1 2 56362 61530
0 12039 5 1 1 12038
0 12040 7 3 2 50697 53187
0 12041 5 1 1 61532
0 12042 7 1 2 48757 57584
0 12043 5 2 1 12042
0 12044 7 1 2 44774 61535
0 12045 5 1 1 12044
0 12046 7 1 2 12041 12045
0 12047 5 2 1 12046
0 12048 7 1 2 43894 61537
0 12049 5 1 1 12048
0 12050 7 1 2 41465 52123
0 12051 5 1 1 12050
0 12052 7 1 2 12049 12051
0 12053 5 1 1 12052
0 12054 7 1 2 53959 12053
0 12055 5 1 1 12054
0 12056 7 1 2 12039 12055
0 12057 5 1 1 12056
0 12058 7 1 2 42568 60257
0 12059 7 1 2 12057 12058
0 12060 5 1 1 12059
0 12061 7 1 2 12032 12060
0 12062 5 1 1 12061
0 12063 7 1 2 44069 12062
0 12064 5 1 1 12063
0 12065 7 6 2 41752 56904
0 12066 7 4 2 45086 57194
0 12067 7 8 2 61539 61545
0 12068 5 1 1 61549
0 12069 7 1 2 61550 54752
0 12070 5 1 1 12069
0 12071 7 4 2 40994 48899
0 12072 5 1 1 61557
0 12073 7 7 2 41795 46383
0 12074 7 4 2 43184 61561
0 12075 5 1 1 61568
0 12076 7 15 2 61558 61569
0 12077 5 10 1 61572
0 12078 7 1 2 44410 61573
0 12079 5 2 1 12078
0 12080 7 1 2 39987 61597
0 12081 5 1 1 12080
0 12082 7 6 2 44411 53960
0 12083 5 1 1 61599
0 12084 7 1 2 60258 61600
0 12085 5 1 1 12084
0 12086 7 1 2 61587 12085
0 12087 5 2 1 12086
0 12088 7 1 2 53180 61605
0 12089 7 1 2 12081 12088
0 12090 5 1 1 12089
0 12091 7 1 2 12070 12090
0 12092 5 1 1 12091
0 12093 7 1 2 41940 12092
0 12094 5 1 1 12093
0 12095 7 2 2 44499 53961
0 12096 5 2 1 61607
0 12097 7 1 2 60259 61608
0 12098 5 1 1 12097
0 12099 7 1 2 61598 12098
0 12100 5 1 1 12099
0 12101 7 1 2 43354 12100
0 12102 5 1 1 12101
0 12103 7 1 2 44500 61606
0 12104 5 1 1 12103
0 12105 7 1 2 12102 12104
0 12106 5 1 1 12105
0 12107 7 1 2 43535 12106
0 12108 5 1 1 12107
0 12109 7 3 2 47182 58668
0 12110 7 6 2 43355 43185
0 12111 7 3 2 61562 61614
0 12112 5 1 1 61620
0 12113 7 1 2 45048 61621
0 12114 7 1 2 61611 12113
0 12115 5 1 1 12114
0 12116 7 1 2 12108 12115
0 12117 5 1 1 12116
0 12118 7 1 2 42101 12117
0 12119 5 1 1 12118
0 12120 7 1 2 12094 12119
0 12121 5 1 1 12120
0 12122 7 1 2 52057 12121
0 12123 5 1 1 12122
0 12124 7 1 2 54084 60777
0 12125 5 1 1 12124
0 12126 7 1 2 44649 57045
0 12127 5 1 1 12126
0 12128 7 1 2 12125 12127
0 12129 5 1 1 12128
0 12130 7 1 2 43536 12129
0 12131 5 1 1 12130
0 12132 7 3 2 54580 51626
0 12133 5 1 1 61623
0 12134 7 1 2 54025 12133
0 12135 5 2 1 12134
0 12136 7 1 2 42102 61626
0 12137 5 1 1 12136
0 12138 7 1 2 61609 12137
0 12139 5 1 1 12138
0 12140 7 1 2 44650 12139
0 12141 5 1 1 12140
0 12142 7 1 2 12131 12141
0 12143 5 1 1 12142
0 12144 7 1 2 60260 12143
0 12145 5 1 1 12144
0 12146 7 1 2 51423 57245
0 12147 7 1 2 60066 12146
0 12148 5 1 1 12147
0 12149 7 1 2 12145 12148
0 12150 5 1 1 12149
0 12151 7 1 2 47330 12150
0 12152 5 1 1 12151
0 12153 7 4 2 42103 60261
0 12154 5 1 1 61628
0 12155 7 1 2 60474 12154
0 12156 5 3 1 12155
0 12157 7 2 2 54071 61632
0 12158 7 2 2 58935 48413
0 12159 7 1 2 61635 61637
0 12160 5 1 1 12159
0 12161 7 3 2 41941 61551
0 12162 5 1 1 61639
0 12163 7 1 2 54085 61633
0 12164 5 1 1 12163
0 12165 7 1 2 12162 12164
0 12166 5 1 1 12165
0 12167 7 1 2 51824 12166
0 12168 5 1 1 12167
0 12169 7 1 2 42104 61574
0 12170 5 1 1 12169
0 12171 7 1 2 57046 60262
0 12172 7 1 2 53160 12171
0 12173 5 1 1 12172
0 12174 7 1 2 12170 12173
0 12175 7 1 2 12168 12174
0 12176 5 1 1 12175
0 12177 7 1 2 44651 12176
0 12178 5 1 1 12177
0 12179 7 1 2 12160 12178
0 12180 7 1 2 12152 12179
0 12181 5 1 1 12180
0 12182 7 1 2 43699 12181
0 12183 5 1 1 12182
0 12184 7 2 2 48030 59254
0 12185 7 2 2 48612 61642
0 12186 7 1 2 61636 61644
0 12187 5 1 1 12186
0 12188 7 4 2 45049 59974
0 12189 7 2 2 61646 59255
0 12190 5 1 1 61650
0 12191 7 2 2 44652 50549
0 12192 7 1 2 61652 61629
0 12193 7 1 2 61651 12192
0 12194 5 1 1 12193
0 12195 7 1 2 12187 12194
0 12196 7 1 2 12183 12195
0 12197 5 1 1 12196
0 12198 7 1 2 42341 12197
0 12199 5 1 1 12198
0 12200 7 1 2 12123 12199
0 12201 5 1 1 12200
0 12202 7 1 2 40799 12201
0 12203 5 1 1 12202
0 12204 7 4 2 41796 45275
0 12205 7 1 2 51424 61654
0 12206 7 1 2 54673 12205
0 12207 7 3 2 50480 57246
0 12208 7 1 2 61612 61658
0 12209 7 1 2 12206 12208
0 12210 5 1 1 12209
0 12211 7 1 2 12203 12210
0 12212 5 1 1 12211
0 12213 7 1 2 55342 12212
0 12214 5 1 1 12213
0 12215 7 1 2 12064 12214
0 12216 5 1 1 12215
0 12217 7 1 2 46245 12216
0 12218 5 1 1 12217
0 12219 7 22 2 53880 57247
0 12220 5 9 1 61661
0 12221 7 1 2 44070 61514
0 12222 5 1 1 12221
0 12223 7 1 2 47917 58201
0 12224 5 1 1 12223
0 12225 7 1 2 42342 47985
0 12226 5 1 1 12225
0 12227 7 1 2 12224 12226
0 12228 5 2 1 12227
0 12229 7 1 2 40800 61692
0 12230 5 2 1 12229
0 12231 7 1 2 48850 47197
0 12232 5 2 1 12231
0 12233 7 3 2 40801 52028
0 12234 7 1 2 61696 61698
0 12235 5 2 1 12234
0 12236 7 1 2 52373 61699
0 12237 5 2 1 12236
0 12238 7 2 2 56176 61218
0 12239 5 2 1 61705
0 12240 7 1 2 61707 60869
0 12241 5 1 1 12240
0 12242 7 1 2 44501 12241
0 12243 5 1 1 12242
0 12244 7 1 2 42105 61700
0 12245 5 2 1 12244
0 12246 7 1 2 12243 61709
0 12247 5 1 1 12246
0 12248 7 1 2 44412 12247
0 12249 5 1 1 12248
0 12250 7 1 2 61703 12249
0 12251 5 1 1 12250
0 12252 7 1 2 43356 12251
0 12253 5 1 1 12252
0 12254 7 1 2 61701 12253
0 12255 5 1 1 12254
0 12256 7 1 2 43537 12255
0 12257 5 1 1 12256
0 12258 7 1 2 61694 12257
0 12259 5 1 1 12258
0 12260 7 1 2 43700 12259
0 12261 5 1 1 12260
0 12262 7 1 2 60873 61477
0 12263 5 1 1 12262
0 12264 7 1 2 12261 12263
0 12265 5 1 1 12264
0 12266 7 1 2 55343 12265
0 12267 5 1 1 12266
0 12268 7 1 2 12222 12267
0 12269 5 1 1 12268
0 12270 7 1 2 61662 12269
0 12271 5 1 1 12270
0 12272 7 6 2 46472 59421
0 12273 7 2 2 48900 61711
0 12274 7 1 2 49267 61538
0 12275 5 1 1 12274
0 12276 7 1 2 412 57933
0 12277 7 1 2 52124 12276
0 12278 5 1 1 12277
0 12279 7 1 2 12275 12278
0 12280 5 1 1 12279
0 12281 7 1 2 61717 12280
0 12282 5 1 1 12281
0 12283 7 1 2 46246 12282
0 12284 7 1 2 12271 12283
0 12285 5 1 1 12284
0 12286 7 5 2 43186 60152
0 12287 7 2 2 49372 61719
0 12288 7 1 2 54333 52575
0 12289 5 1 1 12288
0 12290 7 1 2 48667 12289
0 12291 5 1 1 12290
0 12292 7 2 2 50431 54997
0 12293 5 1 1 61726
0 12294 7 1 2 58328 60443
0 12295 7 2 2 61225 12294
0 12296 7 1 2 48758 8481
0 12297 5 1 1 12296
0 12298 7 1 2 61728 12297
0 12299 5 2 1 12298
0 12300 7 1 2 41466 61730
0 12301 5 1 1 12300
0 12302 7 1 2 12293 12301
0 12303 5 1 1 12302
0 12304 7 1 2 45892 12303
0 12305 5 1 1 12304
0 12306 7 1 2 12291 12305
0 12307 5 1 1 12306
0 12308 7 1 2 40596 12307
0 12309 5 1 1 12308
0 12310 7 1 2 50674 61075
0 12311 5 1 1 12310
0 12312 7 2 2 45666 51596
0 12313 7 1 2 50432 61732
0 12314 5 1 1 12313
0 12315 7 1 2 12311 12314
0 12316 5 2 1 12315
0 12317 7 1 2 53282 61734
0 12318 5 1 1 12317
0 12319 7 1 2 12309 12318
0 12320 5 1 1 12319
0 12321 7 1 2 61724 12320
0 12322 5 1 1 12321
0 12323 7 23 2 48901 57195
0 12324 7 5 2 40376 56703
0 12325 5 5 1 61759
0 12326 7 2 2 61760 60817
0 12327 5 1 1 61769
0 12328 7 1 2 60815 61349
0 12329 5 1 1 12328
0 12330 7 1 2 42569 12329
0 12331 5 1 1 12330
0 12332 7 1 2 61353 12331
0 12333 5 1 1 12332
0 12334 7 1 2 41467 12333
0 12335 5 1 1 12334
0 12336 7 1 2 12327 12335
0 12337 5 1 1 12336
0 12338 7 1 2 40597 12337
0 12339 5 1 1 12338
0 12340 7 1 2 54353 48668
0 12341 7 1 2 60818 12340
0 12342 5 1 1 12341
0 12343 7 1 2 12339 12342
0 12344 5 1 1 12343
0 12345 7 1 2 40802 12344
0 12346 5 1 1 12345
0 12347 7 4 2 40377 53429
0 12348 7 1 2 61771 54514
0 12349 7 1 2 60819 12348
0 12350 5 1 1 12349
0 12351 7 1 2 12346 12350
0 12352 5 1 1 12351
0 12353 7 1 2 61736 12352
0 12354 5 1 1 12353
0 12355 7 1 2 42963 12354
0 12356 7 1 2 12322 12355
0 12357 5 1 1 12356
0 12358 7 1 2 55042 12357
0 12359 7 1 2 12285 12358
0 12360 5 1 1 12359
0 12361 7 1 2 48819 61531
0 12362 5 1 1 12361
0 12363 7 6 2 40951 41352
0 12364 7 1 2 52956 61775
0 12365 7 1 2 56822 12364
0 12366 5 1 1 12365
0 12367 7 1 2 12362 12366
0 12368 5 1 1 12367
0 12369 7 1 2 40378 12368
0 12370 5 1 1 12369
0 12371 7 1 2 41942 53701
0 12372 5 1 1 12371
0 12373 7 1 2 3165 12372
0 12374 5 1 1 12373
0 12375 7 1 2 47647 12374
0 12376 5 1 1 12375
0 12377 7 1 2 58109 48032
0 12378 5 1 1 12377
0 12379 7 1 2 45667 12378
0 12380 5 1 1 12379
0 12381 7 1 2 60418 12380
0 12382 5 1 1 12381
0 12383 7 1 2 42106 12382
0 12384 5 1 1 12383
0 12385 7 1 2 12376 12384
0 12386 5 1 1 12385
0 12387 7 1 2 43357 12386
0 12388 5 1 1 12387
0 12389 7 1 2 53702 49332
0 12390 5 1 1 12389
0 12391 7 1 2 42107 54779
0 12392 7 1 2 54793 12391
0 12393 5 1 1 12392
0 12394 7 1 2 53744 12393
0 12395 7 1 2 12390 12394
0 12396 7 1 2 12388 12395
0 12397 5 1 1 12396
0 12398 7 1 2 54086 12397
0 12399 5 1 1 12398
0 12400 7 1 2 48820 57047
0 12401 5 1 1 12400
0 12402 7 1 2 51889 47918
0 12403 5 1 1 12402
0 12404 7 1 2 51846 12403
0 12405 5 2 1 12404
0 12406 7 1 2 60859 61781
0 12407 5 1 1 12406
0 12408 7 1 2 11202 12407
0 12409 5 1 1 12408
0 12410 7 1 2 43701 12409
0 12411 5 1 1 12410
0 12412 7 1 2 12401 12411
0 12413 7 1 2 12399 12412
0 12414 5 1 1 12413
0 12415 7 1 2 48478 12414
0 12416 5 1 1 12415
0 12417 7 1 2 12370 12416
0 12418 5 1 1 12417
0 12419 7 1 2 60263 12418
0 12420 5 1 1 12419
0 12421 7 1 2 40192 53731
0 12422 5 4 1 12421
0 12423 7 2 2 42108 61783
0 12424 5 1 1 61787
0 12425 7 1 2 53962 61788
0 12426 5 1 1 12425
0 12427 7 1 2 58971 58394
0 12428 7 1 2 61729 12427
0 12429 5 1 1 12428
0 12430 7 1 2 54087 12429
0 12431 5 1 1 12430
0 12432 7 1 2 12426 12431
0 12433 5 1 1 12432
0 12434 7 1 2 41468 12433
0 12435 5 1 1 12434
0 12436 7 2 2 45445 54998
0 12437 5 1 1 61789
0 12438 7 1 2 47968 59658
0 12439 5 1 1 12438
0 12440 7 1 2 12437 12439
0 12441 5 1 1 12440
0 12442 7 1 2 53963 12441
0 12443 5 1 1 12442
0 12444 7 1 2 54088 61727
0 12445 5 1 1 12444
0 12446 7 1 2 57078 10118
0 12447 5 1 1 12446
0 12448 7 1 2 54122 61018
0 12449 7 1 2 12447 12448
0 12450 5 1 1 12449
0 12451 7 1 2 12445 12450
0 12452 7 1 2 12443 12451
0 12453 7 1 2 12435 12452
0 12454 5 1 1 12453
0 12455 7 1 2 40598 12454
0 12456 5 1 1 12455
0 12457 7 4 2 54072 61524
0 12458 7 1 2 61791 61735
0 12459 5 1 1 12458
0 12460 7 5 2 40379 53493
0 12461 5 1 1 61795
0 12462 7 1 2 52342 61019
0 12463 5 1 1 12462
0 12464 7 1 2 12461 12463
0 12465 5 1 1 12464
0 12466 7 1 2 42343 12465
0 12467 5 1 1 12466
0 12468 7 5 2 41469 45446
0 12469 7 2 2 45668 48800
0 12470 7 1 2 61800 61805
0 12471 5 1 1 12470
0 12472 7 1 2 12467 12471
0 12473 5 1 1 12472
0 12474 7 1 2 53964 12473
0 12475 5 1 1 12474
0 12476 7 1 2 12459 12475
0 12477 7 1 2 12456 12476
0 12478 5 1 1 12477
0 12479 7 1 2 59451 12478
0 12480 5 1 1 12479
0 12481 7 1 2 45893 12480
0 12482 7 1 2 12420 12481
0 12483 5 1 1 12482
0 12484 7 1 2 59495 9439
0 12485 5 1 1 12484
0 12486 7 1 2 57048 12485
0 12487 5 1 1 12486
0 12488 7 1 2 60475 61334
0 12489 5 1 1 12488
0 12490 7 1 2 54146 12489
0 12491 5 1 1 12490
0 12492 7 1 2 12487 12491
0 12493 5 1 1 12492
0 12494 7 1 2 41470 12493
0 12495 5 1 1 12494
0 12496 7 6 2 39988 40995
0 12497 7 4 2 61807 60395
0 12498 5 2 1 61813
0 12499 7 4 2 52065 61814
0 12500 5 1 1 61819
0 12501 7 2 2 47010 60264
0 12502 5 1 1 61823
0 12503 7 1 2 45669 61824
0 12504 5 1 1 12503
0 12505 7 1 2 12500 12504
0 12506 5 1 1 12505
0 12507 7 1 2 53965 12506
0 12508 5 1 1 12507
0 12509 7 1 2 12495 12508
0 12510 5 1 1 12509
0 12511 7 1 2 40599 12510
0 12512 5 1 1 12511
0 12513 7 1 2 44775 50499
0 12514 5 1 1 12513
0 12515 7 1 2 61820 12514
0 12516 5 1 1 12515
0 12517 7 2 2 44243 53251
0 12518 7 6 2 45087 45670
0 12519 7 2 2 61827 59732
0 12520 7 1 2 61825 61833
0 12521 5 1 1 12520
0 12522 7 1 2 12516 12521
0 12523 5 1 1 12522
0 12524 7 1 2 53966 12523
0 12525 5 1 1 12524
0 12526 7 1 2 12512 12525
0 12527 5 1 1 12526
0 12528 7 1 2 48669 12527
0 12529 5 1 1 12528
0 12530 7 1 2 48550 50500
0 12531 5 2 1 12530
0 12532 7 6 2 49642 61835
0 12533 7 1 2 61837 61821
0 12534 5 1 1 12533
0 12535 7 1 2 44244 54560
0 12536 7 1 2 61834 12535
0 12537 5 1 1 12536
0 12538 7 1 2 12534 12537
0 12539 5 1 1 12538
0 12540 7 1 2 53967 12539
0 12541 5 1 1 12540
0 12542 7 1 2 42570 12541
0 12543 7 1 2 12529 12542
0 12544 5 1 1 12543
0 12545 7 1 2 40803 12544
0 12546 7 1 2 12483 12545
0 12547 5 1 1 12546
0 12548 7 4 2 52533 54852
0 12549 5 1 1 61843
0 12550 7 3 2 53881 58412
0 12551 5 2 1 61847
0 12552 7 1 2 61312 61848
0 12553 5 2 1 12552
0 12554 7 4 2 44245 45050
0 12555 7 2 2 61854 57013
0 12556 7 2 2 59043 61326
0 12557 7 1 2 61858 61860
0 12558 5 1 1 12557
0 12559 7 1 2 61852 12558
0 12560 5 1 1 12559
0 12561 7 1 2 61844 12560
0 12562 5 1 1 12561
0 12563 7 1 2 60712 61319
0 12564 5 1 1 12563
0 12565 7 10 2 46384 46473
0 12566 7 3 2 42571 61862
0 12567 7 7 2 40600 44200
0 12568 7 1 2 61828 61875
0 12569 7 1 2 61855 12568
0 12570 7 1 2 61872 12569
0 12571 5 1 1 12570
0 12572 7 1 2 12564 12571
0 12573 5 1 1 12572
0 12574 7 1 2 61020 12573
0 12575 5 1 1 12574
0 12576 7 3 2 40601 46622
0 12577 7 7 2 45894 43187
0 12578 7 6 2 42344 43091
0 12579 7 5 2 53882 61892
0 12580 7 1 2 61885 61898
0 12581 7 2 2 61882 12580
0 12582 5 1 1 61903
0 12583 7 2 2 57628 50746
0 12584 7 1 2 56882 61863
0 12585 7 2 2 61905 12584
0 12586 5 1 1 61907
0 12587 7 1 2 54377 61908
0 12588 5 1 1 12587
0 12589 7 1 2 12582 12588
0 12590 7 1 2 12575 12589
0 12591 5 1 1 12590
0 12592 7 1 2 40804 12591
0 12593 5 1 1 12592
0 12594 7 1 2 12562 12593
0 12595 5 1 1 12594
0 12596 7 1 2 47011 12595
0 12597 5 1 1 12596
0 12598 7 1 2 48670 54521
0 12599 5 1 1 12598
0 12600 7 1 2 57563 12599
0 12601 5 3 1 12600
0 12602 7 1 2 52066 61282
0 12603 7 1 2 57089 12602
0 12604 7 1 2 61909 12603
0 12605 5 1 1 12604
0 12606 7 3 2 40805 59452
0 12607 7 2 2 53883 61912
0 12608 7 10 2 49643 61123
0 12609 7 1 2 59422 61917
0 12610 7 1 2 61915 12609
0 12611 5 1 1 12610
0 12612 7 1 2 12605 12611
0 12613 7 1 2 12597 12612
0 12614 5 1 1 12613
0 12615 7 1 2 50510 12614
0 12616 5 1 1 12615
0 12617 7 1 2 61764 53755
0 12618 5 1 1 12617
0 12619 7 11 2 44246 41471
0 12620 7 3 2 61927 51455
0 12621 7 4 2 44201 60334
0 12622 7 1 2 61938 61941
0 12623 7 1 2 12618 12622
0 12624 5 1 1 12623
0 12625 7 1 2 12616 12624
0 12626 5 1 1 12625
0 12627 7 1 2 48631 12626
0 12628 5 1 1 12627
0 12629 7 1 2 51940 53199
0 12630 5 2 1 12629
0 12631 7 1 2 61945 61822
0 12632 5 1 1 12631
0 12633 7 2 2 44071 60265
0 12634 7 1 2 61947 53426
0 12635 5 1 1 12634
0 12636 7 1 2 12632 12635
0 12637 5 1 1 12636
0 12638 7 9 2 48479 48671
0 12639 5 1 1 61949
0 12640 7 1 2 53968 61950
0 12641 7 1 2 12637 12640
0 12642 5 1 1 12641
0 12643 7 1 2 12628 12642
0 12644 7 1 2 12547 12643
0 12645 5 1 1 12644
0 12646 7 1 2 42964 12645
0 12647 5 1 1 12646
0 12648 7 11 2 40806 42965
0 12649 7 2 2 45276 60364
0 12650 7 3 2 40952 40996
0 12651 7 7 2 60380 61971
0 12652 7 1 2 52394 61974
0 12653 7 2 2 61969 12652
0 12654 5 1 1 61981
0 12655 7 6 2 61928 60325
0 12656 7 1 2 54089 61983
0 12657 5 1 1 12656
0 12658 7 1 2 12654 12657
0 12659 5 1 1 12658
0 12660 7 1 2 39989 12659
0 12661 5 1 1 12660
0 12662 7 4 2 54581 57410
0 12663 5 2 1 61989
0 12664 7 1 2 57079 61993
0 12665 5 3 1 12664
0 12666 7 1 2 61984 61995
0 12667 5 1 1 12666
0 12668 7 1 2 12661 12667
0 12669 5 1 1 12668
0 12670 7 1 2 40602 12669
0 12671 5 1 1 12670
0 12672 7 5 2 57029 52834
0 12673 5 5 1 61998
0 12674 7 1 2 55668 57774
0 12675 7 1 2 61999 12674
0 12676 7 1 2 60453 12675
0 12677 5 1 1 12676
0 12678 7 1 2 12671 12677
0 12679 5 1 1 12678
0 12680 7 1 2 50511 12679
0 12681 5 1 1 12680
0 12682 7 3 2 40603 40997
0 12683 7 2 2 60396 62008
0 12684 7 1 2 61792 62011
0 12685 5 1 1 12684
0 12686 7 3 2 48480 59453
0 12687 5 1 1 62013
0 12688 7 8 2 40193 44247
0 12689 7 4 2 45088 45277
0 12690 5 2 1 62024
0 12691 7 2 2 62016 62025
0 12692 7 2 2 41210 49644
0 12693 7 1 2 41100 59733
0 12694 7 1 2 62032 12693
0 12695 7 1 2 62030 12694
0 12696 5 1 1 12695
0 12697 7 1 2 12687 12696
0 12698 5 1 1 12697
0 12699 7 1 2 53969 12698
0 12700 5 1 1 12699
0 12701 7 1 2 12685 12700
0 12702 5 1 1 12701
0 12703 7 1 2 45671 12702
0 12704 5 1 1 12703
0 12705 7 9 2 53970 60454
0 12706 5 5 1 62034
0 12707 7 1 2 48632 62035
0 12708 5 1 1 12707
0 12709 7 2 2 45278 61990
0 12710 5 1 1 62048
0 12711 7 7 2 44248 41101
0 12712 7 3 2 62050 60326
0 12713 5 1 1 62057
0 12714 7 1 2 39990 62058
0 12715 7 1 2 62049 12714
0 12716 5 1 1 12715
0 12717 7 1 2 12708 12716
0 12718 5 1 1 12717
0 12719 7 1 2 61838 12718
0 12720 5 1 1 12719
0 12721 7 4 2 49645 47012
0 12722 7 5 2 46794 51682
0 12723 5 1 1 62064
0 12724 7 1 2 48551 12723
0 12725 5 1 1 12724
0 12726 7 1 2 62060 12725
0 12727 5 1 1 12726
0 12728 7 1 2 56727 12727
0 12729 5 1 1 12728
0 12730 7 1 2 61737 12729
0 12731 5 1 1 12730
0 12732 7 1 2 56378 57158
0 12733 7 1 2 61720 12732
0 12734 5 1 1 12733
0 12735 7 1 2 12731 12734
0 12736 5 1 1 12735
0 12737 7 1 2 55043 12736
0 12738 5 1 1 12737
0 12739 7 1 2 12720 12738
0 12740 7 1 2 12704 12739
0 12741 7 1 2 12681 12740
0 12742 5 1 1 12741
0 12743 7 1 2 61958 12742
0 12744 5 1 1 12743
0 12745 7 1 2 45447 48415
0 12746 5 1 1 12745
0 12747 7 1 2 42345 12746
0 12748 5 1 1 12747
0 12749 7 1 2 61570 12748
0 12750 5 1 1 12749
0 12751 7 1 2 39991 55626
0 12752 5 3 1 12751
0 12753 7 1 2 62069 52077
0 12754 5 1 1 12753
0 12755 7 2 2 57196 12754
0 12756 7 1 2 45089 62072
0 12757 5 1 1 12756
0 12758 7 1 2 12750 12757
0 12759 5 2 1 12758
0 12760 7 1 2 44249 62074
0 12761 5 1 1 12760
0 12762 7 6 2 40998 43188
0 12763 7 1 2 59968 59060
0 12764 5 3 1 12763
0 12765 7 2 2 45672 62082
0 12766 5 1 1 62085
0 12767 7 3 2 45090 60635
0 12768 5 1 1 62087
0 12769 7 1 2 62088 48416
0 12770 5 1 1 12769
0 12771 7 1 2 12766 12770
0 12772 5 1 1 12771
0 12773 7 1 2 62076 12772
0 12774 5 1 1 12773
0 12775 7 1 2 12761 12774
0 12776 5 1 1 12775
0 12777 7 1 2 53884 12776
0 12778 5 1 1 12777
0 12779 7 1 2 40999 62075
0 12780 5 1 1 12779
0 12781 7 1 2 55014 62073
0 12782 5 1 1 12781
0 12783 7 1 2 12780 12782
0 12784 5 1 1 12783
0 12785 7 1 2 48902 12784
0 12786 5 1 1 12785
0 12787 7 1 2 12778 12786
0 12788 5 1 1 12787
0 12789 7 1 2 43895 12788
0 12790 5 1 1 12789
0 12791 7 6 2 41102 45051
0 12792 5 1 1 62090
0 12793 7 3 2 44202 62091
0 12794 7 2 2 62096 59930
0 12795 7 1 2 46474 62099
0 12796 5 1 1 12795
0 12797 7 1 2 61683 12796
0 12798 5 1 1 12797
0 12799 7 1 2 55044 12798
0 12800 5 1 1 12799
0 12801 7 1 2 41103 61640
0 12802 5 1 1 12801
0 12803 7 1 2 61588 12802
0 12804 7 1 2 12800 12803
0 12805 5 1 1 12804
0 12806 7 1 2 60769 12805
0 12807 5 1 1 12806
0 12808 7 2 2 57197 51627
0 12809 7 1 2 57768 62101
0 12810 5 1 1 12809
0 12811 7 5 2 41753 57248
0 12812 7 1 2 54631 62103
0 12813 5 1 1 12812
0 12814 7 1 2 12810 12813
0 12815 5 1 1 12814
0 12816 7 1 2 55045 12815
0 12817 5 1 1 12816
0 12818 7 2 2 41000 41211
0 12819 7 2 2 60397 62108
0 12820 5 1 1 62110
0 12821 7 1 2 54147 62111
0 12822 5 2 1 12821
0 12823 7 2 2 57198 61364
0 12824 7 13 2 39992 40953
0 12825 7 2 2 62116 62051
0 12826 7 1 2 41754 62129
0 12827 7 1 2 62114 12826
0 12828 5 1 1 12827
0 12829 7 1 2 62112 12828
0 12830 7 1 2 12817 12829
0 12831 5 1 1 12830
0 12832 7 1 2 40194 12831
0 12833 5 1 1 12832
0 12834 7 1 2 12807 12833
0 12835 5 1 1 12834
0 12836 7 1 2 51043 12835
0 12837 5 1 1 12836
0 12838 7 1 2 12790 12837
0 12839 5 1 1 12838
0 12840 7 1 2 44776 56348
0 12841 7 1 2 12839 12840
0 12842 5 1 1 12841
0 12843 7 1 2 12744 12842
0 12844 5 1 1 12843
0 12845 7 1 2 42572 12844
0 12846 5 1 1 12845
0 12847 7 1 2 61899 61387
0 12848 7 1 2 61913 12847
0 12849 5 1 1 12848
0 12850 7 4 2 57629 53971
0 12851 5 3 1 62131
0 12852 7 2 2 39993 59044
0 12853 5 1 1 62138
0 12854 7 1 2 59969 12853
0 12855 5 3 1 12854
0 12856 7 1 2 44250 62140
0 12857 5 1 1 12856
0 12858 7 1 2 59095 12857
0 12859 5 2 1 12858
0 12860 7 1 2 48903 62143
0 12861 5 1 1 12860
0 12862 7 1 2 62135 12861
0 12863 5 4 1 12862
0 12864 7 2 2 56177 59734
0 12865 7 1 2 50244 62149
0 12866 7 1 2 57887 12865
0 12867 7 1 2 62145 12866
0 12868 5 1 1 12867
0 12869 7 1 2 12849 12868
0 12870 5 1 1 12869
0 12871 7 1 2 52605 12870
0 12872 5 1 1 12871
0 12873 7 1 2 12846 12872
0 12874 5 1 1 12873
0 12875 7 1 2 49499 12874
0 12876 5 1 1 12875
0 12877 7 1 2 12647 12876
0 12878 7 1 2 12360 12877
0 12879 7 1 2 12218 12878
0 12880 7 1 2 11897 12879
0 12881 5 1 1 12880
0 12882 7 1 2 52915 12881
0 12883 5 1 1 12882
0 12884 7 4 2 41755 56370
0 12885 7 2 2 43092 54354
0 12886 7 1 2 62151 62155
0 12887 5 1 1 12886
0 12888 7 1 2 54148 56028
0 12889 7 1 2 53858 12888
0 12890 5 1 1 12889
0 12891 7 1 2 12887 12890
0 12892 5 1 1 12891
0 12893 7 1 2 41943 12892
0 12894 5 1 1 12893
0 12895 7 3 2 47648 60968
0 12896 7 4 2 45052 58853
0 12897 7 2 2 46385 54313
0 12898 7 1 2 62160 62164
0 12899 7 1 2 62157 12898
0 12900 5 1 1 12899
0 12901 7 1 2 12894 12900
0 12902 5 1 1 12901
0 12903 7 1 2 51044 12902
0 12904 5 1 1 12903
0 12905 7 1 2 59030 50902
0 12906 5 1 1 12905
0 12907 7 1 2 53972 61131
0 12908 5 1 1 12907
0 12909 7 1 2 12906 12908
0 12910 5 1 1 12909
0 12911 7 1 2 43702 12910
0 12912 5 1 1 12911
0 12913 7 1 2 61109 61182
0 12914 5 1 1 12913
0 12915 7 1 2 12912 12914
0 12916 5 1 1 12915
0 12917 7 1 2 47649 12916
0 12918 5 1 1 12917
0 12919 7 1 2 60686 50891
0 12920 5 1 1 12919
0 12921 7 1 2 53973 51351
0 12922 5 1 1 12921
0 12923 7 1 2 12920 12922
0 12924 5 1 1 12923
0 12925 7 1 2 49938 12924
0 12926 5 1 1 12925
0 12927 7 1 2 12918 12926
0 12928 5 1 1 12927
0 12929 7 1 2 43358 12928
0 12930 5 1 1 12929
0 12931 7 2 2 54073 58936
0 12932 5 1 1 62166
0 12933 7 1 2 50875 62167
0 12934 5 2 1 12933
0 12935 7 1 2 60618 62168
0 12936 5 1 1 12935
0 12937 7 1 2 47650 12936
0 12938 5 1 1 12937
0 12939 7 1 2 60644 12938
0 12940 5 1 1 12939
0 12941 7 1 2 49433 12940
0 12942 5 1 1 12941
0 12943 7 1 2 12930 12942
0 12944 5 1 1 12943
0 12945 7 1 2 42346 12944
0 12946 5 1 1 12945
0 12947 7 1 2 60736 54893
0 12948 5 1 1 12947
0 12949 7 2 2 44203 51628
0 12950 7 5 2 42109 60740
0 12951 7 1 2 54794 62172
0 12952 7 1 2 62170 12951
0 12953 5 1 1 12952
0 12954 7 1 2 12948 12953
0 12955 5 1 1 12954
0 12956 7 1 2 49434 12955
0 12957 5 1 1 12956
0 12958 7 1 2 12946 12957
0 12959 5 1 1 12958
0 12960 7 1 2 54412 12959
0 12961 5 1 1 12960
0 12962 7 1 2 12904 12961
0 12963 5 1 1 12962
0 12964 7 1 2 41629 12963
0 12965 5 1 1 12964
0 12966 7 1 2 55683 52218
0 12967 5 1 1 12966
0 12968 7 1 2 55159 12967
0 12969 5 1 1 12968
0 12970 7 1 2 47044 12969
0 12971 5 1 1 12970
0 12972 7 1 2 41212 58760
0 12973 5 1 1 12972
0 12974 7 1 2 12973 61234
0 12975 5 1 1 12974
0 12976 7 2 2 43359 49320
0 12977 5 1 1 62177
0 12978 7 1 2 47118 52214
0 12979 5 1 1 12978
0 12980 7 1 2 62178 12979
0 12981 5 1 1 12980
0 12982 7 1 2 12975 12981
0 12983 7 1 2 12971 12982
0 12984 5 1 1 12983
0 12985 7 1 2 60713 52140
0 12986 7 1 2 12984 12985
0 12987 5 1 1 12986
0 12988 7 1 2 12965 12987
0 12989 5 1 1 12988
0 12990 7 1 2 46093 12989
0 12991 5 1 1 12990
0 12992 7 1 2 42110 60935
0 12993 5 1 1 12992
0 12994 7 1 2 60422 54123
0 12995 5 1 1 12994
0 12996 7 1 2 12993 12995
0 12997 7 1 2 54890 12996
0 12998 5 1 1 12997
0 12999 7 3 2 48481 56774
0 13000 7 1 2 62179 60586
0 13001 7 1 2 12998 13000
0 13002 5 1 1 13001
0 13003 7 1 2 12991 13002
0 13004 5 1 1 13003
0 13005 7 1 2 40807 13004
0 13006 5 1 1 13005
0 13007 7 1 2 48759 52141
0 13008 5 1 1 13007
0 13009 7 1 2 50263 52893
0 13010 5 1 1 13009
0 13011 7 1 2 13008 13010
0 13012 5 1 1 13011
0 13013 7 1 2 46094 13012
0 13014 5 1 1 13013
0 13015 7 1 2 43538 60666
0 13016 7 1 2 52837 13015
0 13017 5 1 1 13016
0 13018 7 1 2 13014 13017
0 13019 5 1 1 13018
0 13020 7 1 2 45895 13019
0 13021 5 1 1 13020
0 13022 7 1 2 49083 53188
0 13023 7 1 2 55831 13022
0 13024 5 1 1 13023
0 13025 7 1 2 13021 13024
0 13026 5 1 1 13025
0 13027 7 1 2 47045 13026
0 13028 5 1 1 13027
0 13029 7 1 2 48482 52736
0 13030 5 1 1 13029
0 13031 7 1 2 54753 49084
0 13032 7 1 2 54945 13031
0 13033 5 1 1 13032
0 13034 7 1 2 13030 13033
0 13035 5 1 1 13034
0 13036 7 1 2 45896 13035
0 13037 5 1 1 13036
0 13038 7 2 2 54314 49085
0 13039 7 1 2 51069 62182
0 13040 5 1 1 13039
0 13041 7 1 2 13037 13040
0 13042 5 1 1 13041
0 13043 7 1 2 48760 13042
0 13044 5 1 1 13043
0 13045 7 2 2 55409 51186
0 13046 7 1 2 53358 62184
0 13047 5 1 1 13046
0 13048 7 1 2 13044 13047
0 13049 7 1 2 13028 13048
0 13050 5 1 1 13049
0 13051 7 1 2 58624 13050
0 13052 5 1 1 13051
0 13053 7 2 2 43360 42804
0 13054 7 1 2 57679 57796
0 13055 5 1 1 13054
0 13056 7 3 2 43539 44777
0 13057 7 1 2 46386 62188
0 13058 7 1 2 55832 13057
0 13059 7 1 2 51693 13058
0 13060 5 1 1 13059
0 13061 7 1 2 13055 13060
0 13062 5 1 1 13061
0 13063 7 1 2 62186 13062
0 13064 5 1 1 13063
0 13065 7 1 2 54391 55984
0 13066 5 1 1 13065
0 13067 7 4 2 40604 45897
0 13068 5 1 1 62191
0 13069 7 1 2 4139 13068
0 13070 5 1 1 13069
0 13071 7 1 2 41472 4153
0 13072 7 1 2 13070 13071
0 13073 5 1 1 13072
0 13074 7 1 2 13066 13073
0 13075 5 1 1 13074
0 13076 7 2 2 46095 58625
0 13077 7 1 2 43540 62195
0 13078 7 1 2 13075 13077
0 13079 5 1 1 13078
0 13080 7 1 2 13064 13079
0 13081 5 1 1 13080
0 13082 7 1 2 51202 13081
0 13083 5 1 1 13082
0 13084 7 1 2 58580 52381
0 13085 7 3 2 44072 59321
0 13086 7 1 2 62197 61209
0 13087 7 1 2 13084 13086
0 13088 5 1 1 13087
0 13089 7 1 2 13083 13088
0 13090 7 1 2 13052 13089
0 13091 5 1 1 13090
0 13092 7 1 2 53885 13091
0 13093 5 1 1 13092
0 13094 7 2 2 40808 59256
0 13095 7 1 2 45673 50131
0 13096 7 1 2 62200 13095
0 13097 7 1 2 60954 13096
0 13098 7 3 2 43703 52970
0 13099 7 1 2 54413 62202
0 13100 7 1 2 13097 13099
0 13101 5 1 1 13100
0 13102 7 1 2 13093 13101
0 13103 5 1 1 13102
0 13104 7 1 2 46841 13103
0 13105 5 1 1 13104
0 13106 7 1 2 57090 60820
0 13107 5 1 1 13106
0 13108 7 4 2 40195 60949
0 13109 7 3 2 54074 62205
0 13110 5 1 1 62209
0 13111 7 1 2 50481 62210
0 13112 5 1 1 13111
0 13113 7 1 2 13107 13112
0 13114 5 1 1 13113
0 13115 7 1 2 53283 49342
0 13116 5 1 1 13115
0 13117 7 1 2 44073 57312
0 13118 5 1 1 13117
0 13119 7 1 2 13116 13118
0 13120 5 1 1 13119
0 13121 7 1 2 40605 13120
0 13122 5 1 1 13121
0 13123 7 1 2 58304 57421
0 13124 5 1 1 13123
0 13125 7 1 2 13122 13124
0 13126 5 1 1 13125
0 13127 7 1 2 48672 13126
0 13128 7 1 2 13114 13127
0 13129 5 1 1 13128
0 13130 7 3 2 49769 49500
0 13131 5 1 1 62212
0 13132 7 1 2 46897 13131
0 13133 5 1 1 13132
0 13134 7 1 2 49501 46922
0 13135 5 1 1 13134
0 13136 7 1 2 49691 13135
0 13137 5 1 1 13136
0 13138 7 1 2 13133 13137
0 13139 5 1 1 13138
0 13140 7 1 2 59550 13139
0 13141 5 1 1 13140
0 13142 7 1 2 49435 49333
0 13143 5 1 1 13142
0 13144 7 1 2 13141 13143
0 13145 5 1 1 13144
0 13146 7 1 2 42347 13145
0 13147 5 1 1 13146
0 13148 7 1 2 49436 61061
0 13149 5 1 1 13148
0 13150 7 1 2 13147 13149
0 13151 5 1 1 13150
0 13152 7 2 2 58565 52133
0 13153 7 1 2 56486 62215
0 13154 7 1 2 13151 13153
0 13155 5 1 1 13154
0 13156 7 1 2 13129 13155
0 13157 7 1 2 13105 13156
0 13158 7 1 2 13006 13157
0 13159 5 1 1 13158
0 13160 7 1 2 60266 13159
0 13161 5 1 1 13160
0 13162 7 5 2 45279 61552
0 13163 5 1 1 62217
0 13164 7 1 2 52395 62218
0 13165 5 2 1 13164
0 13166 7 1 2 47013 61575
0 13167 5 1 1 13166
0 13168 7 1 2 62222 13167
0 13169 5 1 1 13168
0 13170 7 1 2 53822 13169
0 13171 5 1 1 13170
0 13172 7 5 2 42805 53454
0 13173 5 1 1 62224
0 13174 7 1 2 61817 12502
0 13175 5 1 1 13174
0 13176 7 1 2 53974 13175
0 13177 5 1 1 13176
0 13178 7 3 2 41213 46475
0 13179 7 4 2 57630 62229
0 13180 5 1 1 62232
0 13181 7 1 2 59496 13180
0 13182 5 1 1 13181
0 13183 7 1 2 58284 13182
0 13184 5 1 1 13183
0 13185 7 1 2 13184 12820
0 13186 5 1 1 13185
0 13187 7 1 2 54149 13186
0 13188 5 1 1 13187
0 13189 7 1 2 13177 13188
0 13190 5 1 1 13189
0 13191 7 1 2 46795 13190
0 13192 5 1 1 13191
0 13193 7 2 2 53886 59949
0 13194 7 6 2 45448 43189
0 13195 7 1 2 62238 62109
0 13196 7 1 2 62236 13195
0 13197 5 1 1 13196
0 13198 7 1 2 13192 13197
0 13199 5 1 1 13198
0 13200 7 1 2 40196 13199
0 13201 5 1 1 13200
0 13202 7 1 2 62117 57992
0 13203 7 1 2 60375 13202
0 13204 5 1 1 13203
0 13205 7 1 2 13201 13204
0 13206 5 1 1 13205
0 13207 7 1 2 62225 13206
0 13208 5 1 1 13207
0 13209 7 1 2 13171 13208
0 13210 5 1 1 13209
0 13211 7 1 2 48483 13210
0 13212 5 1 1 13211
0 13213 7 1 2 40197 61576
0 13214 5 1 1 13213
0 13215 7 5 2 57631 57199
0 13216 7 4 2 42111 47779
0 13217 5 2 1 62249
0 13218 7 5 2 41104 41756
0 13219 7 2 2 40954 62255
0 13220 7 1 2 62250 62260
0 13221 7 1 2 62244 13220
0 13222 5 1 1 13221
0 13223 7 1 2 13214 13222
0 13224 5 1 1 13223
0 13225 7 1 2 41944 13224
0 13226 5 1 1 13225
0 13227 7 2 2 42112 46796
0 13228 5 1 1 62262
0 13229 7 1 2 61577 62263
0 13230 5 1 1 13229
0 13231 7 1 2 13226 13230
0 13232 5 1 1 13231
0 13233 7 1 2 39994 13232
0 13234 5 1 1 13233
0 13235 7 1 2 52774 58669
0 13236 7 2 2 61571 13235
0 13237 7 1 2 46956 50885
0 13238 5 2 1 13237
0 13239 7 1 2 62264 62266
0 13240 5 1 1 13239
0 13241 7 1 2 13234 13240
0 13242 5 1 1 13241
0 13243 7 1 2 48339 60958
0 13244 7 1 2 13242 13243
0 13245 5 1 1 13244
0 13246 7 1 2 13212 13245
0 13247 5 1 1 13246
0 13248 7 1 2 44927 13247
0 13249 5 1 1 13248
0 13250 7 6 2 41001 41473
0 13251 7 1 2 47014 62268
0 13252 7 1 2 55613 13251
0 13253 7 3 2 60381 60365
0 13254 7 5 2 39995 57171
0 13255 7 1 2 57869 62277
0 13256 7 1 2 62274 13255
0 13257 7 1 2 13252 13256
0 13258 5 1 1 13257
0 13259 7 1 2 13249 13258
0 13260 5 1 1 13259
0 13261 7 1 2 40809 13260
0 13262 5 1 1 13261
0 13263 7 1 2 60267 60842
0 13264 5 1 1 13263
0 13265 7 1 2 61323 13264
0 13266 5 1 1 13265
0 13267 7 1 2 53512 13266
0 13268 5 1 1 13267
0 13269 7 1 2 52079 50650
0 13270 5 1 1 13269
0 13271 7 1 2 48552 13270
0 13272 5 1 1 13271
0 13273 7 1 2 60408 13272
0 13274 5 1 1 13273
0 13275 7 1 2 13268 13274
0 13276 5 1 1 13275
0 13277 7 1 2 42573 13276
0 13278 5 1 1 13277
0 13279 7 2 2 42113 61365
0 13280 5 1 1 62282
0 13281 7 1 2 60031 59385
0 13282 7 1 2 62283 13281
0 13283 5 1 1 13282
0 13284 7 1 2 60476 13283
0 13285 5 1 1 13284
0 13286 7 1 2 54473 61419
0 13287 7 1 2 13285 13286
0 13288 5 1 1 13287
0 13289 7 1 2 13278 13288
0 13290 5 1 1 13289
0 13291 7 1 2 53975 13290
0 13292 5 1 1 13291
0 13293 7 4 2 44074 49646
0 13294 5 1 1 62284
0 13295 7 1 2 45898 62285
0 13296 5 1 1 13295
0 13297 7 1 2 54297 13296
0 13298 5 4 1 13297
0 13299 7 4 2 40198 41945
0 13300 5 2 1 62292
0 13301 7 1 2 62296 13228
0 13302 5 3 1 13301
0 13303 7 1 2 61320 62298
0 13304 7 1 2 62288 13303
0 13305 5 1 1 13304
0 13306 7 5 2 41214 45091
0 13307 7 3 2 62052 62301
0 13308 7 1 2 62306 57132
0 13309 7 1 2 62150 13308
0 13310 7 1 2 55753 13309
0 13311 5 1 1 13310
0 13312 7 1 2 13305 13311
0 13313 5 1 1 13312
0 13314 7 1 2 54150 13313
0 13315 5 1 1 13314
0 13316 7 1 2 13292 13315
0 13317 5 1 1 13316
0 13318 7 1 2 39996 13317
0 13319 5 1 1 13318
0 13320 7 3 2 40199 40955
0 13321 7 3 2 54684 62309
0 13322 5 2 1 62312
0 13323 7 1 2 62313 61946
0 13324 5 1 1 13323
0 13325 7 2 2 56542 62267
0 13326 5 1 1 62317
0 13327 7 1 2 60233 62318
0 13328 5 1 1 13327
0 13329 7 1 2 13324 13328
0 13330 5 1 1 13329
0 13331 7 1 2 59454 13330
0 13332 5 1 1 13331
0 13333 7 2 2 58983 57335
0 13334 5 3 1 62319
0 13335 7 1 2 47583 52526
0 13336 7 1 2 62320 13335
0 13337 5 1 1 13336
0 13338 7 1 2 13332 13337
0 13339 5 1 1 13338
0 13340 7 1 2 49647 13339
0 13341 5 1 1 13340
0 13342 7 1 2 60455 56029
0 13343 5 2 1 13342
0 13344 7 2 2 56644 60327
0 13345 7 2 2 45280 62053
0 13346 7 1 2 62326 62328
0 13347 7 2 2 61790 13346
0 13348 5 1 1 62330
0 13349 7 1 2 62324 13348
0 13350 5 1 1 13349
0 13351 7 1 2 62314 13350
0 13352 5 1 1 13351
0 13353 7 4 2 41474 41797
0 13354 7 3 2 40606 62332
0 13355 7 2 2 47015 62336
0 13356 7 3 2 44204 59184
0 13357 7 2 2 43190 56626
0 13358 7 1 2 62341 62344
0 13359 7 1 2 62339 13358
0 13360 5 1 1 13359
0 13361 7 1 2 13352 13360
0 13362 7 1 2 13341 13361
0 13363 5 1 1 13362
0 13364 7 1 2 44075 13363
0 13365 5 1 1 13364
0 13366 7 4 2 40200 42348
0 13367 7 1 2 53976 62346
0 13368 5 1 1 13367
0 13369 7 1 2 10519 13326
0 13370 5 1 1 13369
0 13371 7 1 2 54151 13370
0 13372 5 1 1 13371
0 13373 7 1 2 13368 13372
0 13374 5 1 1 13373
0 13375 7 1 2 60456 54292
0 13376 7 1 2 13374 13375
0 13377 5 1 1 13376
0 13378 7 1 2 46096 13377
0 13379 7 1 2 13365 13378
0 13380 7 1 2 13319 13379
0 13381 5 1 1 13380
0 13382 7 4 2 42114 49648
0 13383 7 1 2 62223 62113
0 13384 5 1 1 13383
0 13385 7 1 2 62350 13384
0 13386 5 1 1 13385
0 13387 7 2 2 41798 60366
0 13388 7 1 2 57615 62354
0 13389 7 2 2 41002 50225
0 13390 7 1 2 55691 62356
0 13391 7 1 2 13388 13390
0 13392 5 1 1 13391
0 13393 7 1 2 13386 13392
0 13394 5 1 1 13393
0 13395 7 1 2 42349 13394
0 13396 5 1 1 13395
0 13397 7 1 2 39997 60642
0 13398 5 1 1 13397
0 13399 7 3 2 45053 60950
0 13400 7 1 2 46387 62358
0 13401 5 1 1 13400
0 13402 7 1 2 13398 13401
0 13403 5 1 1 13402
0 13404 7 1 2 46797 13403
0 13405 5 1 1 13404
0 13406 7 1 2 47016 53977
0 13407 5 1 1 13406
0 13408 7 1 2 13405 13407
0 13409 5 2 1 13408
0 13410 7 1 2 40201 62361
0 13411 5 1 1 13410
0 13412 7 6 2 41215 58285
0 13413 7 1 2 62363 57049
0 13414 5 1 1 13413
0 13415 7 1 2 13411 13414
0 13416 5 1 1 13415
0 13417 7 5 2 41003 44778
0 13418 7 4 2 60398 62369
0 13419 7 1 2 45674 62374
0 13420 7 1 2 13416 13419
0 13421 5 1 1 13420
0 13422 7 1 2 13396 13421
0 13423 5 1 1 13422
0 13424 7 1 2 40810 13423
0 13425 5 1 1 13424
0 13426 7 7 2 44076 45675
0 13427 5 1 1 62378
0 13428 7 1 2 62379 62362
0 13429 5 1 1 13428
0 13430 7 4 2 49712 50226
0 13431 5 2 1 62385
0 13432 7 2 2 61900 62386
0 13433 5 1 1 62391
0 13434 7 1 2 45449 62392
0 13435 5 1 1 13434
0 13436 7 1 2 13429 13435
0 13437 5 1 1 13436
0 13438 7 1 2 40202 13437
0 13439 5 1 1 13438
0 13440 7 10 2 39998 44077
0 13441 7 1 2 54632 62393
0 13442 7 1 2 56823 13441
0 13443 5 1 1 13442
0 13444 7 1 2 13439 13443
0 13445 5 1 1 13444
0 13446 7 1 2 62014 13445
0 13447 5 1 1 13446
0 13448 7 1 2 13425 13447
0 13449 5 1 1 13448
0 13450 7 1 2 45899 13449
0 13451 5 1 1 13450
0 13452 7 1 2 41105 50433
0 13453 5 4 1 13452
0 13454 7 1 2 62403 60037
0 13455 5 2 1 13454
0 13456 7 1 2 61540 51470
0 13457 7 1 2 61457 13456
0 13458 7 1 2 62407 13457
0 13459 5 1 1 13458
0 13460 7 1 2 42806 13459
0 13461 7 1 2 13451 13460
0 13462 5 1 1 13461
0 13463 7 1 2 41630 13462
0 13464 7 1 2 13381 13463
0 13465 5 1 1 13464
0 13466 7 1 2 13262 13465
0 13467 5 1 1 13466
0 13468 7 1 2 49502 13467
0 13469 5 1 1 13468
0 13470 7 4 2 43896 46476
0 13471 7 2 2 44078 62409
0 13472 7 2 2 48964 62413
0 13473 7 1 2 52885 61158
0 13474 7 1 2 62415 13473
0 13475 5 1 1 13474
0 13476 7 4 2 44413 41475
0 13477 7 2 2 40956 62417
0 13478 7 1 2 50761 52835
0 13479 7 1 2 61615 57358
0 13480 7 1 2 13478 13479
0 13481 7 1 2 62421 13480
0 13482 5 1 1 13481
0 13483 7 1 2 13475 13482
0 13484 5 1 1 13483
0 13485 7 1 2 43541 13484
0 13486 5 1 1 13485
0 13487 7 3 2 56562 59746
0 13488 7 1 2 41476 62423
0 13489 5 1 1 13488
0 13490 7 2 2 58937 51636
0 13491 7 1 2 62426 62416
0 13492 5 1 1 13491
0 13493 7 1 2 13489 13492
0 13494 5 1 1 13493
0 13495 7 1 2 42350 13494
0 13496 5 1 1 13495
0 13497 7 1 2 13486 13496
0 13498 5 1 1 13497
0 13499 7 1 2 43093 13498
0 13500 5 1 1 13499
0 13501 7 1 2 48965 56487
0 13502 5 1 1 13501
0 13503 7 4 2 40811 61525
0 13504 7 1 2 56157 62428
0 13505 5 1 1 13504
0 13506 7 1 2 13502 13505
0 13507 5 1 1 13506
0 13508 7 1 2 57249 56650
0 13509 7 1 2 13507 13508
0 13510 5 1 1 13509
0 13511 7 1 2 13500 13510
0 13512 5 1 1 13511
0 13513 7 1 2 42574 13512
0 13514 5 1 1 13513
0 13515 7 1 2 54152 55684
0 13516 5 1 1 13515
0 13517 7 1 2 54026 13516
0 13518 5 1 1 13517
0 13519 7 4 2 42351 61886
0 13520 7 1 2 62432 49086
0 13521 7 1 2 48882 13520
0 13522 7 1 2 13518 13521
0 13523 5 1 1 13522
0 13524 7 1 2 13514 13523
0 13525 5 1 1 13524
0 13526 7 1 2 47146 13525
0 13527 5 1 1 13526
0 13528 7 7 2 40607 44502
0 13529 7 1 2 49763 62436
0 13530 7 1 2 61533 13529
0 13531 5 1 1 13530
0 13532 7 1 2 53522 13531
0 13533 5 1 1 13532
0 13534 7 1 2 43704 13533
0 13535 5 1 1 13534
0 13536 7 1 2 49583 51825
0 13537 5 1 1 13536
0 13538 7 1 2 55146 54946
0 13539 5 1 1 13538
0 13540 7 1 2 13537 13539
0 13541 5 1 1 13540
0 13542 7 1 2 40812 13541
0 13543 5 1 1 13542
0 13544 7 1 2 13535 13543
0 13545 5 1 1 13544
0 13546 7 1 2 45900 13545
0 13547 5 1 1 13546
0 13548 7 2 2 41946 55725
0 13549 7 1 2 54500 62443
0 13550 7 1 2 58765 13549
0 13551 5 1 1 13550
0 13552 7 1 2 13547 13551
0 13553 5 1 1 13552
0 13554 7 1 2 46097 13553
0 13555 5 1 1 13554
0 13556 7 4 2 49801 62437
0 13557 5 1 1 62445
0 13558 7 1 2 53823 62446
0 13559 5 1 1 13558
0 13560 7 1 2 8803 13559
0 13561 5 1 1 13560
0 13562 7 1 2 41477 13561
0 13563 5 1 1 13562
0 13564 7 2 2 48553 53824
0 13565 5 1 1 62449
0 13566 7 1 2 40813 62450
0 13567 5 1 1 13566
0 13568 7 1 2 13563 13567
0 13569 5 1 1 13568
0 13570 7 1 2 47331 13569
0 13571 5 1 1 13570
0 13572 7 2 2 47409 57364
0 13573 5 1 1 62451
0 13574 7 1 2 48554 54501
0 13575 5 1 1 13574
0 13576 7 1 2 54517 13575
0 13577 5 1 1 13576
0 13578 7 1 2 58214 13577
0 13579 5 1 1 13578
0 13580 7 1 2 13573 13579
0 13581 5 1 1 13580
0 13582 7 1 2 46098 13581
0 13583 5 1 1 13582
0 13584 7 1 2 13571 13583
0 13585 5 1 1 13584
0 13586 7 1 2 60238 13585
0 13587 5 1 1 13586
0 13588 7 1 2 13555 13587
0 13589 5 1 1 13588
0 13590 7 1 2 41631 13589
0 13591 5 1 1 13590
0 13592 7 1 2 51307 50396
0 13593 7 1 2 60923 13592
0 13594 7 1 2 57972 13593
0 13595 5 1 1 13594
0 13596 7 1 2 13591 13595
0 13597 5 1 1 13596
0 13598 7 1 2 48904 13597
0 13599 5 1 1 13598
0 13600 7 1 2 3473 52367
0 13601 5 1 1 13600
0 13602 7 6 2 41947 48613
0 13603 7 3 2 58757 62453
0 13604 7 1 2 57124 50073
0 13605 7 1 2 10720 13604
0 13606 7 1 2 62459 13605
0 13607 7 1 2 13601 13606
0 13608 5 1 1 13607
0 13609 7 1 2 13599 13608
0 13610 5 1 1 13609
0 13611 7 1 2 46388 13610
0 13612 5 1 1 13611
0 13613 7 1 2 48370 60865
0 13614 7 1 2 54414 13613
0 13615 5 1 1 13614
0 13616 7 2 2 41478 60969
0 13617 7 2 2 50559 59847
0 13618 5 1 1 62464
0 13619 7 1 2 13618 60900
0 13620 5 1 1 13619
0 13621 7 1 2 54795 58133
0 13622 5 1 1 13621
0 13623 7 1 2 13620 13622
0 13624 5 1 1 13623
0 13625 7 1 2 62462 13624
0 13626 5 1 1 13625
0 13627 7 1 2 13615 13626
0 13628 5 1 1 13627
0 13629 7 1 2 41948 13628
0 13630 5 1 1 13629
0 13631 7 1 2 52447 61801
0 13632 7 1 2 62447 13631
0 13633 5 1 1 13632
0 13634 7 1 2 13630 13633
0 13635 5 1 1 13634
0 13636 7 1 2 60696 13635
0 13637 5 1 1 13636
0 13638 7 1 2 13612 13637
0 13639 5 1 1 13638
0 13640 7 1 2 43191 13639
0 13641 5 1 1 13640
0 13642 7 1 2 13527 13641
0 13643 5 1 1 13642
0 13644 7 1 2 44653 13643
0 13645 5 1 1 13644
0 13646 7 3 2 54582 60746
0 13647 5 1 1 62466
0 13648 7 1 2 57080 13647
0 13649 5 2 1 13648
0 13650 7 2 2 41949 48555
0 13651 7 1 2 54039 62471
0 13652 7 1 2 62469 13651
0 13653 5 1 1 13652
0 13654 7 1 2 10205 13653
0 13655 5 1 1 13654
0 13656 7 1 2 44503 13655
0 13657 5 1 1 13656
0 13658 7 1 2 56449 60629
0 13659 5 1 1 13658
0 13660 7 1 2 13657 13659
0 13661 5 1 1 13660
0 13662 7 1 2 44414 13661
0 13663 5 1 1 13662
0 13664 7 3 2 54075 59243
0 13665 5 2 1 62473
0 13666 7 1 2 62476 61610
0 13667 5 1 1 13666
0 13668 7 1 2 49584 13667
0 13669 5 1 1 13668
0 13670 7 1 2 13663 13669
0 13671 5 1 1 13670
0 13672 7 1 2 43542 13671
0 13673 5 1 1 13672
0 13674 7 1 2 52847 62474
0 13675 5 1 1 13674
0 13676 7 1 2 46919 61601
0 13677 5 1 1 13676
0 13678 7 1 2 13675 13677
0 13679 5 1 1 13678
0 13680 7 1 2 49585 13679
0 13681 5 1 1 13680
0 13682 7 1 2 45901 13681
0 13683 7 1 2 13673 13682
0 13684 5 1 1 13683
0 13685 7 2 2 45450 48556
0 13686 7 6 2 47780 62465
0 13687 7 1 2 49586 62480
0 13688 5 1 1 13687
0 13689 7 3 2 50201 47274
0 13690 5 2 1 62486
0 13691 7 2 2 49883 62489
0 13692 7 1 2 45676 62491
0 13693 5 1 1 13692
0 13694 7 1 2 13688 13693
0 13695 5 1 1 13694
0 13696 7 1 2 61092 13695
0 13697 5 1 1 13696
0 13698 7 1 2 53978 61806
0 13699 5 1 1 13698
0 13700 7 1 2 13697 13699
0 13701 5 1 1 13700
0 13702 7 1 2 62478 13701
0 13703 5 1 1 13702
0 13704 7 4 2 43705 41479
0 13705 7 2 2 60778 62493
0 13706 5 1 1 62497
0 13707 7 1 2 54027 12932
0 13708 5 4 1 13707
0 13709 7 1 2 62498 62499
0 13710 5 1 1 13709
0 13711 7 3 2 41757 58925
0 13712 7 3 2 45281 48557
0 13713 7 1 2 56814 62506
0 13714 7 1 2 62503 13713
0 13715 5 1 1 13714
0 13716 7 1 2 13710 13715
0 13717 5 1 1 13716
0 13718 7 1 2 43361 13717
0 13719 5 1 1 13718
0 13720 7 1 2 60615 62494
0 13721 7 1 2 47194 13720
0 13722 5 1 1 13721
0 13723 7 1 2 13719 13722
0 13724 5 1 1 13723
0 13725 7 1 2 43543 13724
0 13726 5 1 1 13725
0 13727 7 1 2 42575 13726
0 13728 7 1 2 13703 13727
0 13729 5 1 1 13728
0 13730 7 1 2 13684 13729
0 13731 5 1 1 13730
0 13732 7 1 2 40814 13731
0 13733 5 1 1 13732
0 13734 7 1 2 53455 49334
0 13735 5 1 1 13734
0 13736 7 1 2 40608 48633
0 13737 5 1 1 13736
0 13738 7 1 2 39999 62065
0 13739 5 1 1 13738
0 13740 7 1 2 13737 13739
0 13741 5 1 1 13740
0 13742 7 1 2 54255 13741
0 13743 5 1 1 13742
0 13744 7 1 2 13735 13743
0 13745 5 1 1 13744
0 13746 7 1 2 41480 13745
0 13747 5 1 1 13746
0 13748 7 1 2 54256 53061
0 13749 7 1 2 62066 13748
0 13750 5 1 1 13749
0 13751 7 1 2 13747 13750
0 13752 5 1 1 13751
0 13753 7 1 2 53979 13752
0 13754 5 1 1 13753
0 13755 7 1 2 62481 60926
0 13756 5 1 1 13755
0 13757 7 2 2 41481 53456
0 13758 7 1 2 55928 62509
0 13759 5 1 1 13758
0 13760 7 1 2 13756 13759
0 13761 5 1 1 13760
0 13762 7 1 2 45282 13761
0 13763 5 1 1 13762
0 13764 7 1 2 55754 48790
0 13765 5 1 1 13764
0 13766 7 1 2 13763 13765
0 13767 5 1 1 13766
0 13768 7 1 2 54153 13767
0 13769 5 1 1 13768
0 13770 7 1 2 13754 13769
0 13771 5 1 1 13770
0 13772 7 1 2 45451 13771
0 13773 5 1 1 13772
0 13774 7 1 2 48558 1451
0 13775 5 1 1 13774
0 13776 7 1 2 53980 13775
0 13777 5 1 1 13776
0 13778 7 1 2 12037 13777
0 13779 5 1 1 13778
0 13780 7 1 2 48673 13779
0 13781 5 1 1 13780
0 13782 7 2 2 40000 62000
0 13783 5 1 1 62511
0 13784 7 1 2 48484 52396
0 13785 7 1 2 62512 13784
0 13786 5 1 1 13785
0 13787 7 1 2 13781 13786
0 13788 5 1 1 13787
0 13789 7 1 2 42576 13788
0 13790 5 1 1 13789
0 13791 7 1 2 44079 13790
0 13792 7 1 2 13773 13791
0 13793 5 1 1 13792
0 13794 7 1 2 13733 13793
0 13795 5 1 1 13794
0 13796 7 13 2 40380 43897
0 13797 7 2 2 50972 62513
0 13798 5 1 1 62526
0 13799 7 1 2 13798 13294
0 13800 5 3 1 13799
0 13801 7 2 2 47584 47166
0 13802 7 6 2 40001 42115
0 13803 5 2 1 62533
0 13804 7 2 2 41950 47463
0 13805 5 1 1 62541
0 13806 7 1 2 62539 13805
0 13807 5 1 1 13806
0 13808 7 2 2 62531 13807
0 13809 5 2 1 62543
0 13810 7 1 2 62528 62544
0 13811 5 1 1 13810
0 13812 7 2 2 50454 48674
0 13813 5 2 1 62547
0 13814 7 1 2 62286 62548
0 13815 5 1 1 13814
0 13816 7 1 2 13811 13815
0 13817 5 1 1 13816
0 13818 7 1 2 54154 13817
0 13819 5 1 1 13818
0 13820 7 6 2 49649 48675
0 13821 7 3 2 44080 62551
0 13822 5 2 1 62557
0 13823 7 1 2 52377 62529
0 13824 7 1 2 43544 52848
0 13825 5 1 1 13824
0 13826 7 1 2 47332 53171
0 13827 5 1 1 13826
0 13828 7 1 2 13825 13827
0 13829 7 1 2 13823 13828
0 13830 5 1 1 13829
0 13831 7 1 2 62560 13830
0 13832 5 1 1 13831
0 13833 7 1 2 53981 13832
0 13834 5 1 1 13833
0 13835 7 1 2 13819 13834
0 13836 5 1 1 13835
0 13837 7 1 2 45902 13836
0 13838 5 1 1 13837
0 13839 7 1 2 62545 62549
0 13840 5 1 1 13839
0 13841 7 1 2 54268 13840
0 13842 5 1 1 13841
0 13843 7 4 2 46977 50550
0 13844 5 1 1 62562
0 13845 7 1 2 13844 51013
0 13846 5 1 1 13845
0 13847 7 1 2 54355 13846
0 13848 5 1 1 13847
0 13849 7 2 2 43545 49748
0 13850 7 1 2 45903 59845
0 13851 7 1 2 62566 13850
0 13852 5 1 1 13851
0 13853 7 1 2 13848 13852
0 13854 7 1 2 13842 13853
0 13855 5 1 1 13854
0 13856 7 1 2 54155 13855
0 13857 5 1 1 13856
0 13858 7 1 2 43362 51791
0 13859 5 1 1 13858
0 13860 7 1 2 41951 50191
0 13861 5 1 1 13860
0 13862 7 1 2 13859 13861
0 13863 5 1 1 13862
0 13864 7 1 2 44415 13863
0 13865 5 1 1 13864
0 13866 7 1 2 48485 50312
0 13867 7 1 2 13865 13866
0 13868 5 1 1 13867
0 13869 7 2 2 51890 52084
0 13870 5 1 1 62568
0 13871 7 1 2 61015 62569
0 13872 5 1 1 13871
0 13873 7 1 2 42577 13872
0 13874 7 1 2 13868 13873
0 13875 5 1 1 13874
0 13876 7 1 2 50192 54392
0 13877 7 1 2 49328 13876
0 13878 5 1 1 13877
0 13879 7 1 2 13875 13878
0 13880 5 1 1 13879
0 13881 7 1 2 53982 13880
0 13882 5 1 1 13881
0 13883 7 1 2 13857 13882
0 13884 5 1 1 13883
0 13885 7 1 2 40815 13884
0 13886 5 1 1 13885
0 13887 7 1 2 13838 13886
0 13888 5 1 1 13887
0 13889 7 1 2 42352 13888
0 13890 5 1 1 13889
0 13891 7 2 2 57567 55762
0 13892 7 3 2 41106 44779
0 13893 7 1 2 61441 62572
0 13894 7 1 2 62570 13893
0 13895 5 1 1 13894
0 13896 7 6 2 47085 60970
0 13897 5 1 1 62575
0 13898 7 1 2 48614 62418
0 13899 7 1 2 62576 13898
0 13900 5 1 1 13899
0 13901 7 1 2 13895 13900
0 13902 5 1 1 13901
0 13903 7 3 2 45677 59423
0 13904 7 1 2 62581 57616
0 13905 7 1 2 13902 13904
0 13906 5 1 1 13905
0 13907 7 1 2 41632 13906
0 13908 7 1 2 13890 13907
0 13909 7 1 2 13795 13908
0 13910 5 1 1 13909
0 13911 7 2 2 42116 49716
0 13912 5 1 1 62584
0 13913 7 1 2 41107 13912
0 13914 5 2 1 13913
0 13915 7 1 2 52337 62586
0 13916 5 1 1 13915
0 13917 7 1 2 61901 13916
0 13918 5 1 1 13917
0 13919 7 3 2 44081 46798
0 13920 5 1 1 62588
0 13921 7 1 2 40203 50327
0 13922 5 2 1 13921
0 13923 7 1 2 13920 62591
0 13924 5 1 1 13923
0 13925 7 1 2 40002 13924
0 13926 5 1 1 13925
0 13927 7 1 2 2992 60839
0 13928 5 1 1 13927
0 13929 7 1 2 40204 13928
0 13930 5 1 1 13929
0 13931 7 1 2 13427 13930
0 13932 7 1 2 13926 13931
0 13933 5 2 1 13932
0 13934 7 1 2 45452 62593
0 13935 5 1 1 13934
0 13936 7 1 2 13935 11774
0 13937 5 1 1 13936
0 13938 7 1 2 54156 13937
0 13939 5 1 1 13938
0 13940 7 1 2 13918 13939
0 13941 5 1 1 13940
0 13942 7 1 2 41216 13941
0 13943 5 1 1 13942
0 13944 7 2 2 45453 57133
0 13945 7 1 2 54157 58249
0 13946 7 1 2 62595 13945
0 13947 5 1 1 13946
0 13948 7 1 2 13943 13947
0 13949 5 1 1 13948
0 13950 7 1 2 61951 13949
0 13951 5 1 1 13950
0 13952 7 1 2 61093 59659
0 13953 5 1 1 13952
0 13954 7 1 2 42353 50569
0 13955 5 2 1 13954
0 13956 7 1 2 41217 54158
0 13957 7 1 2 62597 13956
0 13958 5 1 1 13957
0 13959 7 1 2 13953 13958
0 13960 5 1 1 13959
0 13961 7 1 2 53421 13960
0 13962 5 1 1 13961
0 13963 7 2 2 45678 51120
0 13964 5 1 1 62599
0 13965 7 1 2 42354 50235
0 13966 5 1 1 13965
0 13967 7 1 2 57050 13966
0 13968 7 1 2 13964 13967
0 13969 5 1 1 13968
0 13970 7 1 2 45283 55880
0 13971 5 1 1 13970
0 13972 7 1 2 54786 54090
0 13973 7 1 2 53398 13972
0 13974 7 1 2 13971 13973
0 13975 5 1 1 13974
0 13976 7 1 2 13969 13975
0 13977 5 1 1 13976
0 13978 7 1 2 41482 13977
0 13979 5 1 1 13978
0 13980 7 1 2 49681 61624
0 13981 5 1 1 13980
0 13982 7 1 2 57743 13981
0 13983 5 1 1 13982
0 13984 7 1 2 54965 56543
0 13985 7 1 2 13983 13984
0 13986 5 1 1 13985
0 13987 7 1 2 13979 13986
0 13988 7 1 2 13962 13987
0 13989 5 1 1 13988
0 13990 7 1 2 45454 13989
0 13991 5 1 1 13990
0 13992 7 1 2 61625 62552
0 13993 5 1 1 13992
0 13994 7 1 2 57051 50560
0 13995 5 1 1 13994
0 13996 7 1 2 47275 57451
0 13997 7 1 2 60955 13996
0 13998 5 1 1 13997
0 13999 7 1 2 13995 13998
0 14000 5 1 1 13999
0 14001 7 1 2 46891 54970
0 14002 7 1 2 14000 14001
0 14003 5 1 1 14002
0 14004 7 1 2 13993 14003
0 14005 5 1 1 14004
0 14006 7 1 2 42355 14005
0 14007 5 1 1 14006
0 14008 7 1 2 48486 51364
0 14009 7 1 2 61602 14008
0 14010 5 1 1 14009
0 14011 7 1 2 14007 14010
0 14012 7 1 2 13991 14011
0 14013 5 1 1 14012
0 14014 7 1 2 40816 14013
0 14015 5 1 1 14014
0 14016 7 1 2 13951 14015
0 14017 5 1 1 14016
0 14018 7 1 2 45904 14017
0 14019 5 1 1 14018
0 14020 7 3 2 54076 49112
0 14021 7 1 2 62601 53196
0 14022 7 1 2 61918 14021
0 14023 5 1 1 14022
0 14024 7 1 2 44928 14023
0 14025 7 1 2 14019 14024
0 14026 5 1 1 14025
0 14027 7 1 2 13910 14026
0 14028 5 1 1 14027
0 14029 7 1 2 46099 14028
0 14030 5 1 1 14029
0 14031 7 1 2 40609 50732
0 14032 5 1 1 14031
0 14033 7 5 2 52397 57568
0 14034 5 1 1 62604
0 14035 7 1 2 62605 50144
0 14036 7 1 2 62061 14035
0 14037 5 1 1 14036
0 14038 7 1 2 14032 14037
0 14039 5 1 1 14038
0 14040 7 1 2 40817 45284
0 14041 7 1 2 14039 14040
0 14042 5 1 1 14041
0 14043 7 5 2 40818 50733
0 14044 5 1 1 62609
0 14045 7 1 2 14044 57708
0 14046 5 1 1 14045
0 14047 7 1 2 43363 59842
0 14048 5 1 1 14047
0 14049 7 1 2 61536 14048
0 14050 7 1 2 14046 14049
0 14051 5 1 1 14050
0 14052 7 1 2 14042 14051
0 14053 5 1 1 14052
0 14054 7 1 2 45679 14053
0 14055 5 1 1 14054
0 14056 7 1 2 59777 53329
0 14057 7 1 2 13870 14056
0 14058 5 1 1 14057
0 14059 7 1 2 14055 14058
0 14060 5 1 1 14059
0 14061 7 1 2 45905 14060
0 14062 5 1 1 14061
0 14063 7 5 2 53430 51485
0 14064 7 2 2 41218 62614
0 14065 7 3 2 52448 50434
0 14066 7 1 2 62606 62621
0 14067 7 1 2 62619 14066
0 14068 5 1 1 14067
0 14069 7 1 2 14062 14068
0 14070 5 1 1 14069
0 14071 7 1 2 43094 14070
0 14072 5 1 1 14071
0 14073 7 1 2 57680 56178
0 14074 7 1 2 57612 14073
0 14075 5 1 1 14074
0 14076 7 1 2 56048 60043
0 14077 7 1 2 58074 14076
0 14078 5 1 1 14077
0 14079 7 1 2 14075 14078
0 14080 5 1 1 14079
0 14081 7 1 2 51142 14080
0 14082 5 1 1 14081
0 14083 7 1 2 14072 14082
0 14084 5 1 1 14083
0 14085 7 1 2 53887 14084
0 14086 5 1 1 14085
0 14087 7 2 2 47333 56714
0 14088 7 1 2 49884 62624
0 14089 5 1 1 14088
0 14090 7 1 2 61043 53422
0 14091 5 1 1 14090
0 14092 7 1 2 14089 14091
0 14093 5 1 1 14092
0 14094 7 1 2 45455 14093
0 14095 5 1 1 14094
0 14096 7 1 2 51045 51811
0 14097 7 1 2 54971 14096
0 14098 5 1 1 14097
0 14099 7 1 2 14095 14098
0 14100 5 1 1 14099
0 14101 7 1 2 45285 14100
0 14102 5 1 1 14101
0 14103 7 1 2 59789 61420
0 14104 5 1 1 14103
0 14105 7 1 2 62364 60838
0 14106 5 3 1 14105
0 14107 7 1 2 44504 58289
0 14108 5 4 1 14107
0 14109 7 1 2 54999 62629
0 14110 5 1 1 14109
0 14111 7 1 2 62626 14110
0 14112 5 1 1 14111
0 14113 7 1 2 48676 14112
0 14114 5 1 1 14113
0 14115 7 1 2 14104 14114
0 14116 7 1 2 14102 14115
0 14117 5 1 1 14116
0 14118 7 1 2 41633 14117
0 14119 5 1 1 14118
0 14120 7 1 2 1417 61495
0 14121 5 1 1 14120
0 14122 7 1 2 49682 14121
0 14123 5 1 1 14122
0 14124 7 1 2 44929 62365
0 14125 5 1 1 14124
0 14126 7 1 2 14123 14125
0 14127 5 1 1 14126
0 14128 7 1 2 45286 14127
0 14129 5 1 1 14128
0 14130 7 4 2 45680 62630
0 14131 5 1 1 62633
0 14132 7 1 2 44930 62634
0 14133 5 1 1 14132
0 14134 7 1 2 62627 14133
0 14135 7 1 2 14129 14134
0 14136 5 1 1 14135
0 14137 7 1 2 61952 14136
0 14138 5 1 1 14137
0 14139 7 1 2 14119 14138
0 14140 5 1 1 14139
0 14141 7 1 2 40819 14140
0 14142 5 1 1 14141
0 14143 7 3 2 48677 60808
0 14144 7 1 2 8914 61496
0 14145 5 1 1 14144
0 14146 7 1 2 49683 14145
0 14147 5 1 1 14146
0 14148 7 1 2 44082 62366
0 14149 5 1 1 14148
0 14150 7 1 2 14147 14149
0 14151 5 1 1 14150
0 14152 7 1 2 45287 14151
0 14153 5 1 1 14152
0 14154 7 1 2 44083 62635
0 14155 5 1 1 14154
0 14156 7 1 2 62628 14155
0 14157 7 1 2 14153 14156
0 14158 5 1 1 14157
0 14159 7 1 2 62637 14158
0 14160 5 1 1 14159
0 14161 7 1 2 14142 14160
0 14162 5 1 1 14161
0 14163 7 1 2 60234 14162
0 14164 5 1 1 14163
0 14165 7 1 2 42807 14164
0 14166 7 1 2 14086 14165
0 14167 5 1 1 14166
0 14168 7 1 2 43192 14167
0 14169 7 1 2 14030 14168
0 14170 5 1 1 14169
0 14171 7 1 2 54862 59747
0 14172 7 1 2 59605 14171
0 14173 5 1 1 14172
0 14174 7 3 2 42578 59504
0 14175 7 3 2 44505 44780
0 14176 7 1 2 59012 62643
0 14177 7 1 2 62640 14176
0 14178 5 1 1 14177
0 14179 7 1 2 14173 14178
0 14180 5 1 1 14179
0 14181 7 1 2 43898 14180
0 14182 5 1 1 14181
0 14183 7 1 2 54356 62424
0 14184 5 1 1 14183
0 14185 7 1 2 14182 14184
0 14186 5 1 1 14185
0 14187 7 1 2 49321 14186
0 14188 5 1 1 14187
0 14189 7 1 2 41219 50826
0 14190 5 5 1 14189
0 14191 7 1 2 54315 62646
0 14192 5 1 1 14191
0 14193 7 1 2 44506 54393
0 14194 5 1 1 14193
0 14195 7 1 2 14192 14194
0 14196 5 1 1 14195
0 14197 7 1 2 62425 14196
0 14198 5 1 1 14197
0 14199 7 1 2 14188 14198
0 14200 5 1 1 14199
0 14201 7 1 2 43095 14200
0 14202 5 1 1 14201
0 14203 7 1 2 53221 54836
0 14204 5 1 1 14203
0 14205 7 2 2 57250 14204
0 14206 7 2 2 59151 62651
0 14207 7 1 2 48905 62653
0 14208 5 1 1 14207
0 14209 7 1 2 43364 61738
0 14210 5 1 1 14209
0 14211 7 1 2 61684 14210
0 14212 5 1 1 14211
0 14213 7 1 2 44084 50619
0 14214 7 3 2 52134 14213
0 14215 7 1 2 43899 62655
0 14216 7 1 2 14212 14215
0 14217 5 1 1 14216
0 14218 7 1 2 14208 14217
0 14219 5 3 1 14218
0 14220 7 1 2 44507 62658
0 14221 5 1 1 14220
0 14222 7 2 2 57681 59748
0 14223 7 2 2 48559 62661
0 14224 7 2 2 43365 56563
0 14225 7 1 2 62663 62665
0 14226 5 1 1 14225
0 14227 7 1 2 14221 14226
0 14228 5 1 1 14227
0 14229 7 1 2 46842 14228
0 14230 5 1 1 14229
0 14231 7 1 2 14202 14230
0 14232 5 1 1 14231
0 14233 7 1 2 42117 14232
0 14234 5 1 1 14233
0 14235 7 3 2 40820 56458
0 14236 5 1 1 62667
0 14237 7 2 2 62668 58824
0 14238 5 1 1 62670
0 14239 7 1 2 50620 58505
0 14240 5 1 1 14239
0 14241 7 1 2 14238 14240
0 14242 5 1 1 14241
0 14243 7 1 2 43900 14242
0 14244 5 1 1 14243
0 14245 7 1 2 56744 56477
0 14246 5 1 1 14245
0 14247 7 1 2 14244 14246
0 14248 5 3 1 14247
0 14249 7 1 2 49692 57251
0 14250 7 1 2 62672 14249
0 14251 5 1 1 14250
0 14252 7 1 2 46477 56037
0 14253 7 1 2 48966 51435
0 14254 7 1 2 14252 14253
0 14255 7 5 2 43096 47334
0 14256 7 3 2 44205 49268
0 14257 7 1 2 62675 62680
0 14258 7 1 2 14254 14257
0 14259 5 1 1 14258
0 14260 7 1 2 14251 14259
0 14261 5 1 1 14260
0 14262 7 1 2 41952 14261
0 14263 5 1 1 14262
0 14264 7 1 2 47410 61739
0 14265 5 1 1 14264
0 14266 7 1 2 61685 14265
0 14267 5 1 1 14266
0 14268 7 1 2 50118 47335
0 14269 7 1 2 62656 14268
0 14270 7 1 2 14267 14269
0 14271 5 1 1 14270
0 14272 7 1 2 14263 14271
0 14273 5 1 1 14272
0 14274 7 1 2 47046 14273
0 14275 5 1 1 14274
0 14276 7 1 2 55147 62673
0 14277 5 1 1 14276
0 14278 7 1 2 44508 55685
0 14279 7 1 2 62674 14278
0 14280 5 1 1 14279
0 14281 7 1 2 46100 47948
0 14282 7 1 2 57524 14281
0 14283 7 1 2 60627 14282
0 14284 5 1 1 14283
0 14285 7 1 2 14280 14284
0 14286 5 1 1 14285
0 14287 7 1 2 42118 14286
0 14288 5 1 1 14287
0 14289 7 1 2 14277 14288
0 14290 5 1 1 14289
0 14291 7 1 2 57252 14290
0 14292 5 1 1 14291
0 14293 7 1 2 14275 14292
0 14294 7 1 2 14234 14293
0 14295 5 1 1 14294
0 14296 7 1 2 43706 14295
0 14297 5 1 1 14296
0 14298 7 2 2 58926 60630
0 14299 5 1 1 62683
0 14300 7 1 2 46715 54091
0 14301 5 1 1 14300
0 14302 7 1 2 61105 14301
0 14303 5 1 1 14302
0 14304 7 1 2 43366 14303
0 14305 5 1 1 14304
0 14306 7 1 2 14299 14305
0 14307 5 1 1 14306
0 14308 7 1 2 54394 14307
0 14309 5 1 1 14308
0 14310 7 2 2 42579 49379
0 14311 7 1 2 40003 12083
0 14312 5 1 1 14311
0 14313 7 3 2 62500 14312
0 14314 7 1 2 62685 62687
0 14315 5 1 1 14314
0 14316 7 1 2 14309 14315
0 14317 5 1 1 14316
0 14318 7 1 2 59152 14317
0 14319 5 1 1 14318
0 14320 7 1 2 58581 61206
0 14321 7 3 2 43367 49269
0 14322 7 1 2 62690 60806
0 14323 7 1 2 14320 14322
0 14324 5 1 1 14323
0 14325 7 1 2 14319 14324
0 14326 5 1 1 14325
0 14327 7 1 2 43193 54754
0 14328 7 1 2 14326 14327
0 14329 5 1 1 14328
0 14330 7 1 2 14297 14329
0 14331 5 1 1 14330
0 14332 7 1 2 52029 14331
0 14333 5 1 1 14332
0 14334 7 1 2 40381 12977
0 14335 5 1 1 14334
0 14336 7 1 2 62654 14335
0 14337 5 1 1 14336
0 14338 7 2 2 43901 57200
0 14339 7 1 2 52272 62693
0 14340 7 1 2 62657 14339
0 14341 5 1 1 14340
0 14342 7 1 2 14337 14341
0 14343 5 1 1 14342
0 14344 7 1 2 48906 14343
0 14345 5 1 1 14344
0 14346 7 4 2 43194 53888
0 14347 7 1 2 48061 56687
0 14348 5 1 1 14347
0 14349 7 1 2 43368 48603
0 14350 7 1 2 62216 14349
0 14351 5 1 1 14350
0 14352 7 1 2 14348 14351
0 14353 5 1 1 14352
0 14354 7 1 2 43902 14353
0 14355 5 1 1 14354
0 14356 7 1 2 59153 62156
0 14357 5 1 1 14356
0 14358 7 1 2 14355 14357
0 14359 5 1 1 14358
0 14360 7 1 2 49322 14359
0 14361 5 1 1 14360
0 14362 7 2 2 44931 61198
0 14363 7 1 2 58582 62699
0 14364 5 1 1 14363
0 14365 7 1 2 14361 14364
0 14366 5 1 1 14365
0 14367 7 1 2 62695 14366
0 14368 5 1 1 14367
0 14369 7 1 2 14345 14368
0 14370 5 1 1 14369
0 14371 7 1 2 42356 14370
0 14372 5 1 1 14371
0 14373 7 4 2 43369 60971
0 14374 7 7 2 45288 43097
0 14375 7 1 2 62705 60351
0 14376 7 1 2 62701 14375
0 14377 7 1 2 62504 62183
0 14378 7 1 2 14376 14377
0 14379 5 1 1 14378
0 14380 7 1 2 14372 14379
0 14381 5 1 1 14380
0 14382 7 1 2 44654 14381
0 14383 5 1 1 14382
0 14384 7 1 2 57511 13565
0 14385 5 1 1 14384
0 14386 7 1 2 55331 62706
0 14387 7 1 2 61616 56775
0 14388 7 1 2 48353 14387
0 14389 7 1 2 14386 14388
0 14390 7 1 2 14385 14389
0 14391 5 1 1 14390
0 14392 7 1 2 14383 14391
0 14393 5 1 1 14392
0 14394 7 1 2 47047 14393
0 14395 5 1 1 14394
0 14396 7 1 2 54804 62659
0 14397 5 1 1 14396
0 14398 7 1 2 43195 56677
0 14399 7 1 2 54415 14398
0 14400 7 1 2 62666 14399
0 14401 5 1 1 14400
0 14402 7 1 2 14397 14401
0 14403 5 1 1 14402
0 14404 7 1 2 58389 14403
0 14405 5 1 1 14404
0 14406 7 1 2 62380 61802
0 14407 5 1 1 14406
0 14408 7 1 2 2965 14407
0 14409 5 1 1 14408
0 14410 7 2 2 43370 56127
0 14411 7 1 2 62662 62712
0 14412 7 1 2 14409 14411
0 14413 5 1 1 14412
0 14414 7 1 2 14405 14413
0 14415 5 1 1 14414
0 14416 7 1 2 47651 14415
0 14417 5 1 1 14416
0 14418 7 1 2 49885 62660
0 14419 5 1 1 14418
0 14420 7 1 2 54300 60972
0 14421 5 1 1 14420
0 14422 7 1 2 54510 14421
0 14423 5 1 1 14422
0 14424 7 1 2 41483 14423
0 14425 5 1 1 14424
0 14426 7 1 2 40821 54395
0 14427 5 1 1 14426
0 14428 7 1 2 14425 14427
0 14429 5 1 1 14428
0 14430 7 2 2 43196 52687
0 14431 7 1 2 43098 62714
0 14432 7 1 2 62713 14431
0 14433 7 1 2 14429 14432
0 14434 5 1 1 14433
0 14435 7 1 2 14419 14434
0 14436 5 1 1 14435
0 14437 7 1 2 48821 14436
0 14438 5 1 1 14437
0 14439 7 2 2 40957 55787
0 14440 7 1 2 52672 62716
0 14441 7 1 2 53166 14440
0 14442 7 1 2 62664 14441
0 14443 5 1 1 14442
0 14444 7 1 2 14438 14443
0 14445 7 1 2 14417 14444
0 14446 5 1 1 14445
0 14447 7 1 2 46843 14446
0 14448 5 1 1 14447
0 14449 7 1 2 14395 14448
0 14450 7 1 2 14333 14449
0 14451 7 1 2 14170 14450
0 14452 7 1 2 13645 14451
0 14453 5 1 1 14452
0 14454 7 1 2 46623 14453
0 14455 5 1 1 14454
0 14456 7 1 2 13469 14455
0 14457 7 1 2 13161 14456
0 14458 5 1 1 14457
0 14459 7 1 2 42966 14458
0 14460 5 1 1 14459
0 14461 7 1 2 7972 7984
0 14462 5 3 1 14461
0 14463 7 1 2 48062 62718
0 14464 5 1 1 14463
0 14465 7 1 2 49020 59369
0 14466 5 1 1 14465
0 14467 7 1 2 14464 14466
0 14468 5 2 1 14467
0 14469 7 1 2 41004 62721
0 14470 5 1 1 14469
0 14471 7 3 2 41634 60382
0 14472 7 1 2 56909 62723
0 14473 5 1 1 14472
0 14474 7 1 2 14470 14473
0 14475 5 2 1 14474
0 14476 7 1 2 54269 62726
0 14477 5 1 1 14476
0 14478 7 5 2 59203 58670
0 14479 5 1 1 62728
0 14480 7 1 2 9407 14479
0 14481 5 5 1 14480
0 14482 7 2 2 49199 60959
0 14483 5 1 1 62738
0 14484 7 1 2 62733 62739
0 14485 5 1 1 14484
0 14486 7 1 2 14477 14485
0 14487 5 1 1 14486
0 14488 7 3 2 40205 43197
0 14489 7 1 2 58770 62740
0 14490 7 1 2 14487 14489
0 14491 5 1 1 14490
0 14492 7 2 2 46247 55344
0 14493 7 4 2 44932 58656
0 14494 7 1 2 58997 62394
0 14495 7 1 2 61327 14494
0 14496 7 1 2 62745 14495
0 14497 7 1 2 62743 14496
0 14498 5 1 1 14497
0 14499 7 1 2 14491 14498
0 14500 5 1 1 14499
0 14501 7 1 2 46101 14500
0 14502 5 1 1 14501
0 14503 7 1 2 60960 62727
0 14504 5 1 1 14503
0 14505 7 3 2 59910 62370
0 14506 7 1 2 62749 58874
0 14507 5 1 1 14506
0 14508 7 1 2 14504 14507
0 14509 5 1 1 14508
0 14510 7 7 2 42808 43198
0 14511 7 1 2 40004 58771
0 14512 7 1 2 62752 14511
0 14513 7 1 2 14509 14512
0 14514 5 1 1 14513
0 14515 7 1 2 14502 14514
0 14516 5 1 1 14515
0 14517 7 1 2 46389 14516
0 14518 5 1 1 14517
0 14519 7 1 2 44781 58506
0 14520 5 1 1 14519
0 14521 7 1 2 40822 56020
0 14522 5 1 1 14521
0 14523 7 1 2 14483 14522
0 14524 5 1 1 14523
0 14525 7 1 2 49021 14524
0 14526 5 1 1 14525
0 14527 7 1 2 14520 14526
0 14528 5 1 1 14527
0 14529 7 13 2 46248 43199
0 14530 7 3 2 56678 62759
0 14531 7 1 2 40005 62772
0 14532 7 1 2 59522 14531
0 14533 7 1 2 14528 14532
0 14534 5 1 1 14533
0 14535 7 1 2 14518 14534
0 14536 5 1 1 14535
0 14537 7 1 2 49503 14536
0 14538 5 1 1 14537
0 14539 7 2 2 58657 57014
0 14540 7 5 2 44251 44655
0 14541 7 1 2 62777 61864
0 14542 7 1 2 62775 14541
0 14543 7 1 2 53105 59237
0 14544 7 1 2 14542 14543
0 14545 5 1 1 14544
0 14546 7 1 2 14538 14545
0 14547 5 1 1 14546
0 14548 7 1 2 46959 14547
0 14549 5 1 1 14548
0 14550 7 1 2 62132 50382
0 14551 5 1 1 14550
0 14552 7 1 2 45681 59980
0 14553 5 1 1 14552
0 14554 7 1 2 59970 14553
0 14555 5 1 1 14554
0 14556 7 1 2 44252 14555
0 14557 5 1 1 14556
0 14558 7 1 2 59096 14557
0 14559 5 1 1 14558
0 14560 7 1 2 47336 14559
0 14561 5 1 1 14560
0 14562 7 2 2 55046 59931
0 14563 5 1 1 62782
0 14564 7 4 2 43371 61299
0 14565 7 2 2 45092 60741
0 14566 7 1 2 62784 62788
0 14567 5 1 1 14566
0 14568 7 1 2 14563 14567
0 14569 7 1 2 14561 14568
0 14570 5 1 1 14569
0 14571 7 1 2 48907 14570
0 14572 5 1 1 14571
0 14573 7 1 2 14551 14572
0 14574 5 1 1 14573
0 14575 7 1 2 49886 14574
0 14576 5 1 1 14575
0 14577 7 2 2 55047 48908
0 14578 5 1 1 62790
0 14579 7 1 2 14578 7687
0 14580 5 17 1 14579
0 14581 7 23 2 43099 62792
0 14582 7 2 2 62809 55889
0 14583 5 1 1 62832
0 14584 7 2 2 62793 62676
0 14585 5 1 1 62834
0 14586 7 1 2 52030 62835
0 14587 5 1 1 14586
0 14588 7 1 2 14583 14587
0 14589 7 1 2 14576 14588
0 14590 5 1 1 14589
0 14591 7 1 2 42119 14590
0 14592 5 1 1 14591
0 14593 7 1 2 44253 53889
0 14594 5 1 1 14593
0 14595 7 1 2 14594 12072
0 14596 5 3 1 14595
0 14597 7 2 2 59084 62836
0 14598 5 1 1 62839
0 14599 7 4 2 44206 61856
0 14600 7 1 2 59950 62841
0 14601 5 1 1 14600
0 14602 7 1 2 14598 14601
0 14603 5 1 1 14602
0 14604 7 1 2 52219 14603
0 14605 5 1 1 14604
0 14606 7 6 2 44254 48909
0 14607 7 1 2 62845 59981
0 14608 7 1 2 51834 14607
0 14609 5 1 1 14608
0 14610 7 1 2 14605 14609
0 14611 5 1 1 14610
0 14612 7 1 2 47337 14611
0 14613 5 1 1 14612
0 14614 7 1 2 50455 52220
0 14615 5 1 1 14614
0 14616 7 1 2 51384 14615
0 14617 5 1 1 14616
0 14618 7 1 2 62810 14617
0 14619 5 1 1 14618
0 14620 7 1 2 59045 62842
0 14621 7 1 2 53672 14620
0 14622 5 1 1 14621
0 14623 7 3 2 59046 54917
0 14624 7 1 2 44255 48761
0 14625 7 1 2 58940 14624
0 14626 7 1 2 62851 14625
0 14627 5 1 1 14626
0 14628 7 1 2 14622 14627
0 14629 7 1 2 14619 14628
0 14630 7 1 2 14613 14629
0 14631 5 1 1 14630
0 14632 7 1 2 47652 14631
0 14633 5 1 1 14632
0 14634 7 1 2 47781 56390
0 14635 5 1 1 14634
0 14636 7 1 2 48762 14635
0 14637 5 1 1 14636
0 14638 7 1 2 50836 54060
0 14639 5 1 1 14638
0 14640 7 1 2 60995 14639
0 14641 7 1 2 14637 14640
0 14642 5 1 1 14641
0 14643 7 1 2 62811 14642
0 14644 5 1 1 14643
0 14645 7 1 2 44656 46990
0 14646 5 1 1 14645
0 14647 7 1 2 55874 14646
0 14648 5 1 1 14647
0 14649 7 2 2 48910 57632
0 14650 7 7 2 46390 62854
0 14651 7 1 2 42357 62856
0 14652 7 1 2 14648 14651
0 14653 5 1 1 14652
0 14654 7 1 2 47727 48763
0 14655 7 1 2 58998 14654
0 14656 7 1 2 62852 14655
0 14657 5 1 1 14656
0 14658 7 1 2 45906 14657
0 14659 7 1 2 14653 14658
0 14660 7 1 2 14644 14659
0 14661 7 1 2 14633 14660
0 14662 7 1 2 14592 14661
0 14663 5 1 1 14662
0 14664 7 1 2 58195 11456
0 14665 5 1 1 14664
0 14666 7 1 2 62146 14665
0 14667 5 1 1 14666
0 14668 7 1 2 54124 58197
0 14669 5 1 1 14668
0 14670 7 1 2 62857 14669
0 14671 5 1 1 14670
0 14672 7 1 2 42580 14671
0 14673 7 1 2 14667 14672
0 14674 5 1 1 14673
0 14675 7 1 2 14663 14674
0 14676 5 1 1 14675
0 14677 7 1 2 46478 14676
0 14678 5 1 1 14677
0 14679 7 2 2 40958 57985
0 14680 7 1 2 59951 60800
0 14681 5 1 1 14680
0 14682 7 1 2 9100 14681
0 14683 5 1 1 14682
0 14684 7 1 2 42120 14683
0 14685 5 1 1 14684
0 14686 7 2 2 45093 42358
0 14687 7 2 2 46391 62865
0 14688 7 1 2 59801 62867
0 14689 5 1 1 14688
0 14690 7 1 2 14685 14689
0 14691 5 1 1 14690
0 14692 7 1 2 45907 14691
0 14693 5 1 1 14692
0 14694 7 1 2 41220 13280
0 14695 5 1 1 14694
0 14696 7 1 2 49437 14695
0 14697 5 1 1 14696
0 14698 7 1 2 42581 62086
0 14699 7 1 2 14697 14698
0 14700 5 1 1 14699
0 14701 7 1 2 14693 14700
0 14702 5 1 1 14701
0 14703 7 1 2 62863 14702
0 14704 5 1 1 14703
0 14705 7 1 2 45908 59559
0 14706 5 1 1 14705
0 14707 7 1 2 49438 53156
0 14708 5 1 1 14707
0 14709 7 1 2 52449 14708
0 14710 5 1 1 14709
0 14711 7 1 2 14706 14710
0 14712 5 1 1 14711
0 14713 7 1 2 62837 61563
0 14714 7 1 2 14712 14713
0 14715 5 1 1 14714
0 14716 7 1 2 43200 14715
0 14717 7 1 2 14704 14716
0 14718 5 1 1 14717
0 14719 7 1 2 48266 14718
0 14720 7 1 2 14678 14719
0 14721 5 1 1 14720
0 14722 7 2 2 59177 60021
0 14723 5 1 1 62869
0 14724 7 1 2 45909 61731
0 14725 5 1 1 14724
0 14726 7 1 2 52450 9029
0 14727 5 2 1 14726
0 14728 7 1 2 14725 62871
0 14729 5 1 1 14728
0 14730 7 1 2 62870 14729
0 14731 5 1 1 14730
0 14732 7 1 2 45910 60492
0 14733 5 1 1 14732
0 14734 7 2 2 59291 49087
0 14735 7 1 2 41221 53409
0 14736 5 1 1 14735
0 14737 7 2 2 42582 48764
0 14738 5 1 1 62875
0 14739 7 1 2 62876 60488
0 14740 7 1 2 14736 14739
0 14741 5 1 1 14740
0 14742 7 1 2 62873 14741
0 14743 7 1 2 14733 14742
0 14744 5 1 1 14743
0 14745 7 1 2 14731 14744
0 14746 5 1 1 14745
0 14747 7 1 2 46392 14746
0 14748 5 1 1 14747
0 14749 7 1 2 45911 60445
0 14750 5 1 1 14749
0 14751 7 1 2 62872 14750
0 14752 5 1 1 14751
0 14753 7 6 2 41005 43100
0 14754 5 1 1 62877
0 14755 7 3 2 41799 46249
0 14756 7 1 2 49088 62883
0 14757 7 1 2 62878 14756
0 14758 7 1 2 14752 14757
0 14759 5 1 1 14758
0 14760 7 1 2 14748 14759
0 14761 5 1 1 14760
0 14762 7 1 2 43201 14761
0 14763 5 1 1 14762
0 14764 7 4 2 54602 49089
0 14765 5 4 1 62886
0 14766 7 1 2 56657 55571
0 14767 5 1 1 14766
0 14768 7 1 2 62890 14767
0 14769 5 2 1 14768
0 14770 7 1 2 51828 62894
0 14771 5 1 1 14770
0 14772 7 2 2 53636 51655
0 14773 7 1 2 47849 62896
0 14774 5 1 1 14773
0 14775 7 1 2 57475 48358
0 14776 5 1 1 14775
0 14777 7 1 2 14774 14776
0 14778 5 1 1 14777
0 14779 7 1 2 42359 14778
0 14780 5 1 1 14779
0 14781 7 1 2 14771 14780
0 14782 5 1 1 14781
0 14783 7 1 2 47338 14782
0 14784 5 1 1 14783
0 14785 7 3 2 57476 58860
0 14786 5 1 1 62898
0 14787 7 3 2 48580 58797
0 14788 7 1 2 44933 62901
0 14789 5 1 1 14788
0 14790 7 1 2 14786 14789
0 14791 5 1 1 14790
0 14792 7 1 2 43707 14791
0 14793 5 1 1 14792
0 14794 7 1 2 50456 50132
0 14795 7 1 2 53540 14794
0 14796 5 1 1 14795
0 14797 7 1 2 14793 14796
0 14798 5 1 1 14797
0 14799 7 1 2 45682 14798
0 14800 5 1 1 14799
0 14801 7 1 2 56100 58802
0 14802 5 1 1 14801
0 14803 7 1 2 57477 54221
0 14804 5 1 1 14803
0 14805 7 4 2 43372 44934
0 14806 7 3 2 44416 62904
0 14807 7 1 2 53606 62908
0 14808 5 1 1 14807
0 14809 7 1 2 14804 14808
0 14810 5 1 1 14809
0 14811 7 1 2 50338 50426
0 14812 7 1 2 14810 14811
0 14813 5 1 1 14812
0 14814 7 1 2 14802 14813
0 14815 7 1 2 14800 14814
0 14816 7 1 2 14784 14815
0 14817 5 1 1 14816
0 14818 7 1 2 47653 14817
0 14819 5 1 1 14818
0 14820 7 1 2 48038 2816
0 14821 5 1 1 14820
0 14822 7 1 2 42121 14821
0 14823 5 1 1 14822
0 14824 7 1 2 50313 14823
0 14825 5 1 1 14824
0 14826 7 1 2 45683 14825
0 14827 5 1 1 14826
0 14828 7 1 2 58368 14827
0 14829 5 1 1 14828
0 14830 7 1 2 58635 14829
0 14831 5 1 1 14830
0 14832 7 2 2 50339 47339
0 14833 7 1 2 59501 62911
0 14834 5 1 1 14833
0 14835 7 1 2 60416 14834
0 14836 5 1 1 14835
0 14837 7 1 2 42122 14836
0 14838 5 1 1 14837
0 14839 7 1 2 50340 48765
0 14840 7 1 2 56395 14839
0 14841 5 1 1 14840
0 14842 7 1 2 56422 58976
0 14843 5 1 1 14842
0 14844 7 1 2 47728 47969
0 14845 5 1 1 14844
0 14846 7 1 2 58069 14845
0 14847 7 1 2 14843 14846
0 14848 7 1 2 14841 14847
0 14849 7 1 2 14838 14848
0 14850 5 1 1 14849
0 14851 7 1 2 62887 14850
0 14852 5 1 1 14851
0 14853 7 3 2 42123 62899
0 14854 5 1 1 62913
0 14855 7 1 2 56658 51431
0 14856 5 1 1 14855
0 14857 7 1 2 14854 14856
0 14858 5 1 1 14857
0 14859 7 1 2 47782 62600
0 14860 5 1 1 14859
0 14861 7 1 2 11740 14860
0 14862 7 1 2 14858 14861
0 14863 5 1 1 14862
0 14864 7 1 2 45912 14863
0 14865 7 1 2 14852 14864
0 14866 7 1 2 14831 14865
0 14867 7 1 2 14819 14866
0 14868 5 1 1 14867
0 14869 7 2 2 51172 53591
0 14870 5 1 1 62916
0 14871 7 1 2 41635 14870
0 14872 5 1 1 14871
0 14873 7 1 2 44935 61246
0 14874 5 1 1 14873
0 14875 7 1 2 42809 14874
0 14876 7 1 2 14872 14875
0 14877 5 1 1 14876
0 14878 7 1 2 46102 58849
0 14879 7 1 2 53859 14878
0 14880 5 1 1 14879
0 14881 7 1 2 14877 14880
0 14882 5 1 1 14881
0 14883 7 1 2 53637 14882
0 14884 5 1 1 14883
0 14885 7 1 2 48634 54903
0 14886 5 1 1 14885
0 14887 7 1 2 52352 14886
0 14888 5 1 1 14887
0 14889 7 1 2 45684 14888
0 14890 5 1 1 14889
0 14891 7 1 2 61452 14890
0 14892 5 1 1 14891
0 14893 7 1 2 62888 14892
0 14894 5 1 1 14893
0 14895 7 1 2 42583 14894
0 14896 7 1 2 14884 14895
0 14897 5 1 1 14896
0 14898 7 1 2 14868 14897
0 14899 5 1 1 14898
0 14900 7 1 2 57633 14899
0 14901 5 1 1 14900
0 14902 7 2 2 59174 60490
0 14903 5 1 1 62918
0 14904 7 1 2 47919 60006
0 14905 5 1 1 14904
0 14906 7 2 2 62919 14905
0 14907 5 1 1 62920
0 14908 7 1 2 58276 62921
0 14909 5 1 1 14908
0 14910 7 1 2 45913 14909
0 14911 5 1 1 14910
0 14912 7 1 2 61351 14911
0 14913 5 1 1 14912
0 14914 7 1 2 57380 14913
0 14915 5 1 1 14914
0 14916 7 1 2 57670 14915
0 14917 5 1 1 14916
0 14918 7 1 2 57535 14917
0 14919 7 1 2 14901 14918
0 14920 5 1 1 14919
0 14921 7 1 2 14763 14920
0 14922 5 1 1 14921
0 14923 7 1 2 49022 14922
0 14924 5 1 1 14923
0 14925 7 8 2 43202 55048
0 14926 7 3 2 53890 62922
0 14927 5 1 1 62930
0 14928 7 2 2 61559 60399
0 14929 5 1 1 62933
0 14930 7 1 2 14927 14929
0 14931 5 1 1 14930
0 14932 7 2 2 48105 56002
0 14933 7 2 2 47340 58529
0 14934 5 1 1 62937
0 14935 7 1 2 41353 58227
0 14936 5 1 1 14935
0 14937 7 1 2 41953 14936
0 14938 5 1 1 14937
0 14939 7 1 2 14934 14938
0 14940 5 1 1 14939
0 14941 7 1 2 62935 14940
0 14942 5 1 1 14941
0 14943 7 1 2 47533 62938
0 14944 5 1 1 14943
0 14945 7 1 2 45914 61406
0 14946 7 1 2 14944 14945
0 14947 5 1 1 14946
0 14948 7 1 2 42584 61448
0 14949 5 1 1 14948
0 14950 7 1 2 56219 14949
0 14951 7 1 2 14947 14950
0 14952 5 1 1 14951
0 14953 7 1 2 14942 14952
0 14954 5 1 1 14953
0 14955 7 1 2 14931 14954
0 14956 5 1 1 14955
0 14957 7 2 2 41108 44657
0 14958 7 2 2 42360 62939
0 14959 7 1 2 62941 48188
0 14960 5 1 1 14959
0 14961 7 1 2 54227 14960
0 14962 5 1 1 14961
0 14963 7 1 2 45915 14962
0 14964 5 1 1 14963
0 14965 7 1 2 44417 54237
0 14966 5 1 1 14965
0 14967 7 1 2 40006 54248
0 14968 7 1 2 14966 14967
0 14969 5 1 1 14968
0 14970 7 1 2 45456 48249
0 14971 7 1 2 55548 14970
0 14972 5 1 1 14971
0 14973 7 1 2 54250 14972
0 14974 7 1 2 14969 14973
0 14975 7 1 2 14964 14974
0 14976 5 1 1 14975
0 14977 7 5 2 46479 48911
0 14978 7 1 2 57634 62943
0 14979 7 1 2 14976 14978
0 14980 5 1 1 14979
0 14981 7 1 2 14956 14980
0 14982 5 1 1 14981
0 14983 7 1 2 46393 14982
0 14984 5 1 1 14983
0 14985 7 1 2 42124 48250
0 14986 5 1 1 14985
0 14987 7 1 2 48194 14986
0 14988 5 1 1 14987
0 14989 7 1 2 48766 14988
0 14990 5 1 1 14989
0 14991 7 1 2 42361 48251
0 14992 5 1 1 14991
0 14993 7 1 2 14990 14992
0 14994 5 1 1 14993
0 14995 7 1 2 45916 14994
0 14996 5 1 1 14995
0 14997 7 3 2 42585 48106
0 14998 7 2 2 45685 62948
0 14999 7 1 2 41636 49770
0 15000 7 1 2 62951 14999
0 15001 5 1 1 15000
0 15002 7 1 2 14996 15001
0 15003 5 1 1 15002
0 15004 7 1 2 62036 15003
0 15005 5 1 1 15004
0 15006 7 1 2 14984 15005
0 15007 7 1 2 14924 15006
0 15008 7 1 2 14721 15007
0 15009 5 1 1 15008
0 15010 7 1 2 53531 15009
0 15011 5 1 1 15010
0 15012 7 1 2 14549 15011
0 15013 7 1 2 14460 15012
0 15014 7 1 2 12883 15013
0 15015 7 2 2 45917 60911
0 15016 5 1 1 62953
0 15017 7 1 2 50482 62954
0 15018 5 1 1 15017
0 15019 7 1 2 3462 56553
0 15020 5 2 1 15019
0 15021 7 2 2 41109 62955
0 15022 7 1 2 55669 62957
0 15023 5 1 1 15022
0 15024 7 1 2 15018 15023
0 15025 5 1 1 15024
0 15026 7 1 2 45289 15025
0 15027 5 1 1 15026
0 15028 7 1 2 52594 15027
0 15029 5 1 1 15028
0 15030 7 1 2 44085 15029
0 15031 5 1 1 15030
0 15032 7 1 2 44509 60871
0 15033 5 1 1 15032
0 15034 7 1 2 61710 15033
0 15035 5 1 1 15034
0 15036 7 1 2 44418 15035
0 15037 5 1 1 15036
0 15038 7 1 2 61704 15037
0 15039 5 1 1 15038
0 15040 7 1 2 43373 15039
0 15041 5 1 1 15040
0 15042 7 1 2 61702 15041
0 15043 5 1 1 15042
0 15044 7 1 2 43546 15043
0 15045 5 1 1 15044
0 15046 7 1 2 61695 15045
0 15047 5 1 1 15046
0 15048 7 1 2 43708 15047
0 15049 5 1 1 15048
0 15050 7 2 2 44658 61478
0 15051 5 1 1 62959
0 15052 7 1 2 51092 15051
0 15053 5 1 1 15052
0 15054 7 1 2 60866 15053
0 15055 5 1 1 15054
0 15056 7 1 2 15049 15055
0 15057 5 1 1 15056
0 15058 7 1 2 42586 15057
0 15059 5 1 1 15058
0 15060 7 1 2 15031 15059
0 15061 5 1 1 15060
0 15062 7 1 2 46250 15061
0 15063 5 1 1 15062
0 15064 7 8 2 45457 54846
0 15065 5 1 1 62961
0 15066 7 2 2 56795 62962
0 15067 7 1 2 51288 58336
0 15068 7 1 2 62969 15067
0 15069 5 1 1 15068
0 15070 7 1 2 15063 15069
0 15071 5 1 1 15070
0 15072 7 1 2 57382 15071
0 15073 5 1 1 15072
0 15074 7 8 2 42967 46480
0 15075 7 5 2 51532 62971
0 15076 7 1 2 59424 62979
0 15077 7 1 2 53349 15076
0 15078 5 1 1 15077
0 15079 7 1 2 46103 15078
0 15080 7 1 2 15073 15079
0 15081 5 1 1 15080
0 15082 7 1 2 52820 60821
0 15083 5 2 1 15082
0 15084 7 1 2 49439 61485
0 15085 5 1 1 15084
0 15086 7 1 2 51093 15085
0 15087 5 1 1 15086
0 15088 7 1 2 42362 15087
0 15089 5 1 1 15088
0 15090 7 1 2 61480 15089
0 15091 5 3 1 15090
0 15092 7 1 2 41637 62986
0 15093 5 1 1 15092
0 15094 7 1 2 62984 15093
0 15095 5 1 1 15094
0 15096 7 5 2 44086 42587
0 15097 5 1 1 62989
0 15098 7 1 2 57288 62990
0 15099 7 1 2 15095 15098
0 15100 5 1 1 15099
0 15101 7 1 2 57388 52135
0 15102 7 1 2 62987 15101
0 15103 5 1 1 15102
0 15104 7 2 2 52343 61491
0 15105 5 1 1 62994
0 15106 7 1 2 51656 60929
0 15107 5 1 1 15106
0 15108 7 1 2 15105 15107
0 15109 5 1 1 15108
0 15110 7 2 2 56796 52534
0 15111 7 1 2 60505 62996
0 15112 7 1 2 15109 15111
0 15113 5 1 1 15112
0 15114 7 1 2 15103 15113
0 15115 5 1 1 15114
0 15116 7 1 2 40823 15115
0 15117 5 1 1 15116
0 15118 7 1 2 42810 15117
0 15119 7 1 2 15100 15118
0 15120 5 1 1 15119
0 15121 7 1 2 41484 15120
0 15122 7 1 2 15081 15121
0 15123 5 1 1 15122
0 15124 7 1 2 43903 62995
0 15125 5 1 1 15124
0 15126 7 1 2 59884 60930
0 15127 5 1 1 15126
0 15128 7 1 2 15125 15127
0 15129 5 1 1 15128
0 15130 7 1 2 48678 15129
0 15131 5 1 1 15130
0 15132 7 1 2 61465 61473
0 15133 5 1 1 15132
0 15134 7 1 2 44419 15133
0 15135 5 1 1 15134
0 15136 7 1 2 61471 15135
0 15137 5 1 1 15136
0 15138 7 1 2 43374 15137
0 15139 5 1 1 15138
0 15140 7 1 2 61459 15139
0 15141 5 1 1 15140
0 15142 7 1 2 40824 15141
0 15143 5 1 1 15142
0 15144 7 1 2 15131 15143
0 15145 5 1 1 15144
0 15146 7 1 2 57386 15145
0 15147 5 1 1 15146
0 15148 7 6 2 51533 57389
0 15149 5 1 1 62998
0 15150 7 1 2 52279 52311
0 15151 5 1 1 15150
0 15152 7 2 2 60220 48388
0 15153 5 1 1 63004
0 15154 7 1 2 40610 15153
0 15155 5 1 1 15154
0 15156 7 1 2 52031 52353
0 15157 7 1 2 15155 15156
0 15158 5 1 1 15157
0 15159 7 1 2 15151 15158
0 15160 5 1 1 15159
0 15161 7 1 2 47048 15160
0 15162 5 1 1 15161
0 15163 7 1 2 53026 61506
0 15164 5 1 1 15163
0 15165 7 1 2 53023 61504
0 15166 7 1 2 15164 15165
0 15167 5 1 1 15166
0 15168 7 1 2 15162 15167
0 15169 5 1 1 15168
0 15170 7 1 2 62999 15169
0 15171 5 1 1 15170
0 15172 7 1 2 15147 15171
0 15173 5 1 1 15172
0 15174 7 1 2 46104 15173
0 15175 5 1 1 15174
0 15176 7 7 2 60574 62972
0 15177 7 1 2 43904 47049
0 15178 5 2 1 15177
0 15179 7 1 2 63013 61512
0 15180 5 1 1 15179
0 15181 7 1 2 52032 15180
0 15182 5 1 1 15181
0 15183 7 1 2 61508 15182
0 15184 5 1 1 15183
0 15185 7 1 2 41638 15184
0 15186 5 1 1 15185
0 15187 7 1 2 62985 15186
0 15188 5 1 1 15187
0 15189 7 1 2 44087 15188
0 15190 5 1 1 15189
0 15191 7 1 2 48435 62988
0 15192 5 1 1 15191
0 15193 7 1 2 15190 15192
0 15194 5 1 1 15193
0 15195 7 1 2 63006 15194
0 15196 5 1 1 15195
0 15197 7 1 2 45918 15196
0 15198 7 1 2 15175 15197
0 15199 5 1 1 15198
0 15200 7 2 2 63007 61487
0 15201 7 2 2 43905 63015
0 15202 5 1 1 63017
0 15203 7 1 2 11792 61502
0 15204 5 1 1 15203
0 15205 7 1 2 60506 52709
0 15206 7 1 2 15204 15205
0 15207 5 1 1 15206
0 15208 7 1 2 15202 15207
0 15209 5 1 1 15208
0 15210 7 1 2 41639 15209
0 15211 5 1 1 15210
0 15212 7 2 2 48107 57201
0 15213 7 1 2 49133 63019
0 15214 7 1 2 52125 15213
0 15215 5 1 1 15214
0 15216 7 1 2 15211 15215
0 15217 5 1 1 15216
0 15218 7 1 2 40825 15217
0 15219 5 1 1 15218
0 15220 7 2 2 44088 48267
0 15221 5 1 1 63021
0 15222 7 1 2 63022 62694
0 15223 7 1 2 52126 15222
0 15224 5 1 1 15223
0 15225 7 1 2 42588 15224
0 15226 7 1 2 15219 15225
0 15227 5 1 1 15226
0 15228 7 1 2 44782 15227
0 15229 7 1 2 15199 15228
0 15230 5 1 1 15229
0 15231 7 1 2 46920 50551
0 15232 5 2 1 15231
0 15233 7 1 2 42125 47838
0 15234 5 1 1 15233
0 15235 7 1 2 63023 15234
0 15236 5 1 1 15235
0 15237 7 1 2 49440 15236
0 15238 5 1 1 15237
0 15239 7 1 2 61411 59583
0 15240 5 1 1 15239
0 15241 7 1 2 47920 50047
0 15242 5 1 1 15241
0 15243 7 1 2 49504 15242
0 15244 5 1 1 15243
0 15245 7 1 2 47050 15244
0 15246 5 1 1 15245
0 15247 7 1 2 15240 15246
0 15248 5 1 1 15247
0 15249 7 1 2 42363 15248
0 15250 5 1 1 15249
0 15251 7 1 2 15238 15250
0 15252 5 1 1 15251
0 15253 7 1 2 60890 15252
0 15254 5 1 1 15253
0 15255 7 3 2 50183 53257
0 15256 7 1 2 52471 63025
0 15257 5 1 1 15256
0 15258 7 1 2 57139 62958
0 15259 5 1 1 15258
0 15260 7 1 2 52527 54441
0 15261 7 1 2 60912 15260
0 15262 5 1 1 15261
0 15263 7 1 2 15259 15262
0 15264 5 1 1 15263
0 15265 7 1 2 45290 15264
0 15266 5 1 1 15265
0 15267 7 1 2 15257 15266
0 15268 7 1 2 15254 15267
0 15269 5 1 1 15268
0 15270 7 1 2 57298 15269
0 15271 5 1 1 15270
0 15272 7 1 2 54474 63018
0 15273 5 1 1 15272
0 15274 7 1 2 15271 15273
0 15275 5 1 1 15274
0 15276 7 1 2 41640 15275
0 15277 5 1 1 15276
0 15278 7 1 2 53258 61770
0 15279 5 1 1 15278
0 15280 7 1 2 54442 61489
0 15281 5 1 1 15280
0 15282 7 1 2 15279 15281
0 15283 5 1 1 15282
0 15284 7 1 2 42811 15283
0 15285 5 1 1 15284
0 15286 7 1 2 54820 58305
0 15287 7 1 2 52127 15286
0 15288 5 1 1 15287
0 15289 7 1 2 15285 15288
0 15290 5 1 1 15289
0 15291 7 1 2 57226 15290
0 15292 5 1 1 15291
0 15293 7 1 2 15277 15292
0 15294 7 1 2 15230 15293
0 15295 7 1 2 15123 15294
0 15296 5 1 1 15295
0 15297 7 1 2 55049 15296
0 15298 5 1 1 15297
0 15299 7 1 2 47464 60457
0 15300 5 1 1 15299
0 15301 7 6 2 40007 50227
0 15302 5 3 1 63028
0 15303 7 1 2 63029 61283
0 15304 5 1 1 15303
0 15305 7 1 2 15300 15304
0 15306 5 1 1 15305
0 15307 7 1 2 45291 15306
0 15308 5 1 1 15307
0 15309 7 1 2 60268 48781
0 15310 5 1 1 15309
0 15311 7 1 2 15308 15310
0 15312 5 2 1 15311
0 15313 7 1 2 46683 63037
0 15314 5 1 1 15313
0 15315 7 2 2 62026 59505
0 15316 7 1 2 62054 50770
0 15317 7 1 2 63039 15316
0 15318 5 1 1 15317
0 15319 7 1 2 15314 15318
0 15320 5 1 1 15319
0 15321 7 1 2 40206 15320
0 15322 5 1 1 15321
0 15323 7 4 2 41222 44936
0 15324 7 2 2 63041 61655
0 15325 7 1 2 61808 59749
0 15326 7 1 2 63045 15325
0 15327 5 1 1 15326
0 15328 7 1 2 15322 15327
0 15329 5 1 1 15328
0 15330 7 1 2 57888 15329
0 15331 5 1 1 15330
0 15332 7 2 2 43203 60064
0 15333 7 1 2 61809 48340
0 15334 7 1 2 57937 15333
0 15335 7 1 2 63047 15334
0 15336 5 1 1 15335
0 15337 7 4 2 62017 60328
0 15338 5 1 1 63049
0 15339 7 1 2 50107 51471
0 15340 7 1 2 63050 15339
0 15341 5 1 1 15340
0 15342 7 1 2 15336 15341
0 15343 5 1 1 15342
0 15344 7 1 2 44937 50228
0 15345 7 1 2 15343 15344
0 15346 5 1 1 15345
0 15347 7 1 2 15331 15346
0 15348 5 1 1 15347
0 15349 7 1 2 45458 15348
0 15350 5 1 1 15349
0 15351 7 1 2 48436 60458
0 15352 5 1 1 15351
0 15353 7 2 2 46481 49200
0 15354 7 1 2 52811 61369
0 15355 7 1 2 63053 15354
0 15356 5 1 1 15355
0 15357 7 1 2 15352 15356
0 15358 5 1 1 15357
0 15359 7 1 2 52688 15358
0 15360 5 1 1 15359
0 15361 7 6 2 41006 60068
0 15362 7 2 2 62753 63055
0 15363 7 1 2 40826 63061
0 15364 5 1 1 15363
0 15365 7 1 2 15360 15364
0 15366 5 1 1 15365
0 15367 7 1 2 49650 15366
0 15368 5 1 1 15367
0 15369 7 5 2 40207 41007
0 15370 7 1 2 63063 59750
0 15371 7 1 2 53568 15370
0 15372 7 1 2 57938 63046
0 15373 7 1 2 15371 15372
0 15374 5 1 1 15373
0 15375 7 1 2 15368 15374
0 15376 5 1 1 15375
0 15377 7 1 2 42364 15376
0 15378 5 1 1 15377
0 15379 7 1 2 15350 15378
0 15380 5 1 1 15379
0 15381 7 1 2 46251 15380
0 15382 5 1 1 15381
0 15383 7 1 2 60528 57889
0 15384 5 1 1 15383
0 15385 7 1 2 57894 15384
0 15386 5 1 1 15385
0 15387 7 1 2 46252 15386
0 15388 5 1 1 15387
0 15389 7 1 2 55595 59988
0 15390 5 1 1 15389
0 15391 7 1 2 15388 15390
0 15392 5 1 1 15391
0 15393 7 1 2 61331 15392
0 15394 5 1 1 15393
0 15395 7 4 2 40827 53062
0 15396 7 10 2 42968 43204
0 15397 7 6 2 46105 63072
0 15398 7 2 2 41008 41641
0 15399 7 1 2 62333 63088
0 15400 7 1 2 63082 15399
0 15401 7 1 2 63068 15400
0 15402 5 1 1 15401
0 15403 7 1 2 15394 15402
0 15404 5 1 1 15403
0 15405 7 1 2 52080 15404
0 15406 5 1 1 15405
0 15407 7 1 2 53154 62587
0 15408 5 1 1 15407
0 15409 7 1 2 59455 15408
0 15410 5 1 1 15409
0 15411 7 2 2 51742 52324
0 15412 7 1 2 63090 60269
0 15413 5 1 1 15412
0 15414 7 1 2 15410 15413
0 15415 5 1 1 15414
0 15416 7 3 2 40828 50771
0 15417 7 4 2 48487 48108
0 15418 5 1 1 63095
0 15419 7 1 2 63092 63096
0 15420 7 1 2 15415 15419
0 15421 5 1 1 15420
0 15422 7 1 2 15406 15421
0 15423 7 1 2 15382 15422
0 15424 5 1 1 15423
0 15425 7 1 2 41354 15424
0 15426 5 1 1 15425
0 15427 7 1 2 46253 48437
0 15428 7 1 2 61284 15427
0 15429 7 1 2 51173 55596
0 15430 7 1 2 15428 15429
0 15431 5 1 1 15430
0 15432 7 1 2 15426 15431
0 15433 5 1 1 15432
0 15434 7 1 2 40382 15433
0 15435 5 1 1 15434
0 15436 7 1 2 62253 53576
0 15437 5 1 1 15436
0 15438 7 1 2 41954 15437
0 15439 5 1 1 15438
0 15440 7 1 2 53553 15439
0 15441 5 1 1 15440
0 15442 7 1 2 61985 15441
0 15443 5 1 1 15442
0 15444 7 2 2 41223 55642
0 15445 5 1 1 63099
0 15446 7 1 2 41485 59673
0 15447 5 1 1 15446
0 15448 7 1 2 15445 15447
0 15449 5 1 1 15448
0 15450 7 1 2 59456 15449
0 15451 5 1 1 15450
0 15452 7 1 2 15443 15451
0 15453 5 1 1 15452
0 15454 7 1 2 40611 15453
0 15455 5 1 1 15454
0 15456 7 3 2 43205 55643
0 15457 7 1 2 57987 62269
0 15458 7 1 2 63101 15457
0 15459 5 1 1 15458
0 15460 7 1 2 15455 15459
0 15461 5 1 1 15460
0 15462 7 1 2 42365 15461
0 15463 5 1 1 15462
0 15464 7 1 2 60270 51829
0 15465 5 1 1 15464
0 15466 7 1 2 61342 15465
0 15467 5 1 1 15466
0 15468 7 1 2 60435 15467
0 15469 5 1 1 15468
0 15470 7 1 2 41955 58162
0 15471 5 1 1 15470
0 15472 7 1 2 48767 59873
0 15473 5 1 1 15472
0 15474 7 1 2 15471 15473
0 15475 7 1 2 51245 15474
0 15476 5 1 1 15475
0 15477 7 1 2 42126 15476
0 15478 5 1 1 15477
0 15479 7 1 2 49505 58819
0 15480 7 1 2 15478 15479
0 15481 5 1 1 15480
0 15482 7 1 2 61332 15481
0 15483 5 1 1 15482
0 15484 7 1 2 15469 15483
0 15485 5 1 1 15484
0 15486 7 1 2 48488 15485
0 15487 5 1 1 15486
0 15488 7 1 2 44938 15487
0 15489 7 1 2 15463 15488
0 15490 5 1 1 15489
0 15491 7 1 2 47411 51064
0 15492 7 1 2 58142 15491
0 15493 5 1 1 15492
0 15494 7 1 2 42127 51785
0 15495 5 1 1 15494
0 15496 7 1 2 15493 15495
0 15497 5 1 1 15496
0 15498 7 1 2 47729 61285
0 15499 7 1 2 15497 15498
0 15500 5 1 1 15499
0 15501 7 6 2 43375 45094
0 15502 7 2 2 63104 59386
0 15503 7 3 2 44659 50582
0 15504 7 1 2 52668 63112
0 15505 7 1 2 63110 15504
0 15506 5 1 1 15505
0 15507 7 1 2 60459 49789
0 15508 5 1 1 15507
0 15509 7 1 2 49887 62375
0 15510 5 1 1 15509
0 15511 7 1 2 15508 15510
0 15512 7 1 2 15506 15511
0 15513 7 1 2 15500 15512
0 15514 5 1 1 15513
0 15515 7 1 2 41956 15514
0 15516 5 1 1 15515
0 15517 7 1 2 47730 58137
0 15518 7 1 2 54733 15517
0 15519 5 1 1 15518
0 15520 7 1 2 45292 50922
0 15521 5 1 1 15520
0 15522 7 1 2 15519 15521
0 15523 5 1 1 15522
0 15524 7 1 2 51261 15523
0 15525 5 1 1 15524
0 15526 7 1 2 47970 50980
0 15527 5 1 1 15526
0 15528 7 1 2 15525 15527
0 15529 5 1 1 15528
0 15530 7 1 2 60271 15529
0 15531 5 1 1 15530
0 15532 7 1 2 15516 15531
0 15533 5 1 1 15532
0 15534 7 1 2 43906 15533
0 15535 5 1 1 15534
0 15536 7 2 2 49825 51316
0 15537 5 1 1 63115
0 15538 7 1 2 15537 51735
0 15539 5 1 1 15538
0 15540 7 1 2 42366 15539
0 15541 5 1 1 15540
0 15542 7 1 2 49826 53682
0 15543 7 1 2 58440 15542
0 15544 5 1 1 15543
0 15545 7 1 2 15541 15544
0 15546 5 1 1 15545
0 15547 7 1 2 44783 60272
0 15548 7 1 2 15546 15547
0 15549 5 1 1 15548
0 15550 7 1 2 60460 51284
0 15551 5 1 1 15550
0 15552 7 1 2 62404 51132
0 15553 5 1 1 15552
0 15554 7 1 2 45686 60655
0 15555 5 1 1 15554
0 15556 7 1 2 55968 15555
0 15557 5 1 1 15556
0 15558 7 1 2 15553 15557
0 15559 5 1 1 15558
0 15560 7 1 2 60273 52894
0 15561 7 1 2 15559 15560
0 15562 5 1 1 15561
0 15563 7 1 2 15551 15562
0 15564 5 1 1 15563
0 15565 7 1 2 47654 15564
0 15566 5 1 1 15565
0 15567 7 1 2 41642 15566
0 15568 7 1 2 15549 15567
0 15569 7 1 2 15535 15568
0 15570 5 1 1 15569
0 15571 7 1 2 46106 15570
0 15572 7 1 2 15490 15571
0 15573 5 1 1 15572
0 15574 7 3 2 48489 47228
0 15575 5 2 1 63117
0 15576 7 1 2 59457 51365
0 15577 5 1 1 15576
0 15578 7 1 2 60274 14903
0 15579 5 1 1 15578
0 15580 7 1 2 15577 15579
0 15581 5 1 1 15580
0 15582 7 1 2 46844 15581
0 15583 5 1 1 15582
0 15584 7 1 2 54053 54745
0 15585 5 1 1 15584
0 15586 7 1 2 40008 58761
0 15587 5 1 1 15586
0 15588 7 1 2 42128 15587
0 15589 7 1 2 15585 15588
0 15590 5 1 1 15589
0 15591 7 1 2 48679 56391
0 15592 5 1 1 15591
0 15593 7 1 2 51847 58277
0 15594 5 1 1 15593
0 15595 7 1 2 15592 15594
0 15596 5 1 1 15595
0 15597 7 1 2 15590 15596
0 15598 5 1 1 15597
0 15599 7 1 2 60275 15598
0 15600 5 1 1 15599
0 15601 7 1 2 52221 63111
0 15602 5 1 1 15601
0 15603 7 1 2 61343 15602
0 15604 5 1 1 15603
0 15605 7 1 2 60423 15604
0 15606 5 1 1 15605
0 15607 7 1 2 61324 15606
0 15608 7 1 2 15600 15607
0 15609 7 1 2 15583 15608
0 15610 5 1 1 15609
0 15611 7 1 2 63118 15610
0 15612 5 1 1 15611
0 15613 7 1 2 15573 15612
0 15614 5 1 1 15613
0 15615 7 1 2 40829 15614
0 15616 5 1 1 15615
0 15617 7 2 2 59285 59117
0 15618 7 1 2 51220 59754
0 15619 7 1 2 63122 15618
0 15620 7 1 2 60943 15619
0 15621 5 1 1 15620
0 15622 7 1 2 15616 15621
0 15623 5 1 1 15622
0 15624 7 1 2 46254 15623
0 15625 5 1 1 15624
0 15626 7 1 2 15435 15625
0 15627 5 1 1 15626
0 15628 7 1 2 45919 15627
0 15629 5 1 1 15628
0 15630 7 2 2 50651 61124
0 15631 7 1 2 60529 52081
0 15632 5 1 1 15631
0 15633 7 1 2 46684 51097
0 15634 5 1 1 15633
0 15635 7 1 2 15632 15634
0 15636 5 1 1 15635
0 15637 7 1 2 63124 15636
0 15638 5 1 1 15637
0 15639 7 1 2 49090 53351
0 15640 5 1 1 15639
0 15641 7 1 2 15638 15640
0 15642 5 1 1 15641
0 15643 7 1 2 40830 15642
0 15644 5 1 1 15643
0 15645 7 1 2 49651 55289
0 15646 7 1 2 61439 15645
0 15647 5 1 1 15646
0 15648 7 1 2 15644 15647
0 15649 5 1 1 15648
0 15650 7 1 2 54871 60276
0 15651 7 1 2 15649 15650
0 15652 5 1 1 15651
0 15653 7 5 2 40831 41009
0 15654 7 1 2 63126 61656
0 15655 7 1 2 57608 15654
0 15656 7 2 2 50796 61803
0 15657 7 3 2 41110 54847
0 15658 7 1 2 63133 63083
0 15659 7 1 2 63131 15658
0 15660 7 1 2 15655 15659
0 15661 5 1 1 15660
0 15662 7 1 2 15652 15661
0 15663 7 1 2 15629 15662
0 15664 5 1 1 15663
0 15665 7 1 2 43101 15664
0 15666 5 1 1 15665
0 15667 7 1 2 47731 58271
0 15668 5 1 1 15667
0 15669 7 1 2 50929 15668
0 15670 5 1 1 15669
0 15671 7 1 2 51662 8616
0 15672 5 1 1 15671
0 15673 7 1 2 41643 15672
0 15674 7 1 2 15670 15673
0 15675 5 1 1 15674
0 15676 7 1 2 50537 52995
0 15677 5 1 1 15676
0 15678 7 1 2 15675 15677
0 15679 5 1 1 15678
0 15680 7 1 2 60277 15679
0 15681 5 1 1 15680
0 15682 7 1 2 44939 62482
0 15683 5 1 1 15682
0 15684 7 1 2 53683 62563
0 15685 5 1 1 15684
0 15686 7 1 2 15683 15685
0 15687 5 1 1 15686
0 15688 7 1 2 50435 15687
0 15689 5 1 1 15688
0 15690 7 1 2 51612 55851
0 15691 5 1 1 15690
0 15692 7 1 2 50986 15691
0 15693 5 1 1 15692
0 15694 7 1 2 41957 15693
0 15695 5 1 1 15694
0 15696 7 1 2 49939 58457
0 15697 5 1 1 15696
0 15698 7 1 2 1483 15697
0 15699 7 1 2 15695 15698
0 15700 5 1 1 15699
0 15701 7 1 2 41644 15700
0 15702 5 1 1 15701
0 15703 7 1 2 15689 15702
0 15704 5 1 1 15703
0 15705 7 1 2 59458 15704
0 15706 5 1 1 15705
0 15707 7 1 2 15681 15706
0 15708 5 1 1 15707
0 15709 7 1 2 46107 15708
0 15710 5 1 1 15709
0 15711 7 1 2 61044 50436
0 15712 5 1 1 15711
0 15713 7 1 2 48788 15712
0 15714 5 1 1 15713
0 15715 7 1 2 63062 15714
0 15716 5 1 1 15715
0 15717 7 1 2 15710 15716
0 15718 5 1 1 15717
0 15719 7 1 2 44089 15718
0 15720 5 1 1 15719
0 15721 7 3 2 41355 57635
0 15722 7 1 2 40383 49201
0 15723 7 2 2 63136 15722
0 15724 7 1 2 59506 63139
0 15725 5 1 1 15724
0 15726 7 4 2 44090 63042
0 15727 7 1 2 59459 50762
0 15728 7 1 2 63141 15727
0 15729 5 1 1 15728
0 15730 7 1 2 15725 15729
0 15731 5 1 1 15730
0 15732 7 1 2 50720 15731
0 15733 5 1 1 15732
0 15734 7 1 2 47341 52715
0 15735 5 1 1 15734
0 15736 7 1 2 53117 15735
0 15737 5 1 1 15736
0 15738 7 1 2 50483 15737
0 15739 5 1 1 15738
0 15740 7 1 2 48438 53139
0 15741 5 1 1 15740
0 15742 7 1 2 15739 15741
0 15743 5 1 1 15742
0 15744 7 1 2 60400 60388
0 15745 7 1 2 50255 15744
0 15746 7 1 2 15743 15745
0 15747 5 1 1 15746
0 15748 7 1 2 15733 15747
0 15749 7 1 2 15720 15748
0 15750 5 1 1 15749
0 15751 7 1 2 43907 15750
0 15752 5 1 1 15751
0 15753 7 1 2 46108 53033
0 15754 7 1 2 58441 15753
0 15755 5 1 1 15754
0 15756 7 1 2 52753 15755
0 15757 5 1 1 15756
0 15758 7 1 2 41645 15757
0 15759 5 1 1 15758
0 15760 7 1 2 46685 59650
0 15761 5 1 1 15760
0 15762 7 1 2 15759 15761
0 15763 5 1 1 15762
0 15764 7 1 2 48768 15763
0 15765 5 1 1 15764
0 15766 7 1 2 56068 50952
0 15767 5 1 1 15766
0 15768 7 1 2 45687 58435
0 15769 5 1 1 15768
0 15770 7 1 2 49441 49963
0 15771 7 1 2 15769 15770
0 15772 5 1 1 15771
0 15773 7 1 2 15767 15772
0 15774 5 1 1 15773
0 15775 7 1 2 41646 15774
0 15776 5 1 1 15775
0 15777 7 1 2 15765 15776
0 15778 5 1 1 15777
0 15779 7 1 2 59460 15778
0 15780 5 1 1 15779
0 15781 7 2 2 49964 50343
0 15782 7 4 2 44256 41647
0 15783 7 2 2 60329 63147
0 15784 7 1 2 63145 63151
0 15785 7 1 2 51358 15784
0 15786 5 1 1 15785
0 15787 7 1 2 15780 15786
0 15788 5 1 1 15787
0 15789 7 1 2 44091 15788
0 15790 5 1 1 15789
0 15791 7 1 2 45459 56405
0 15792 5 1 1 15791
0 15793 7 1 2 55285 15792
0 15794 5 1 1 15793
0 15795 7 4 2 43908 41010
0 15796 7 1 2 63153 58332
0 15797 7 1 2 63048 15796
0 15798 7 1 2 15794 15797
0 15799 5 1 1 15798
0 15800 7 1 2 15790 15799
0 15801 5 1 1 15800
0 15802 7 1 2 47655 15801
0 15803 5 1 1 15802
0 15804 7 1 2 60401 62395
0 15805 7 1 2 56101 15804
0 15806 7 1 2 62357 15805
0 15807 5 1 1 15806
0 15808 7 3 2 41958 46482
0 15809 7 1 2 63157 63140
0 15810 5 1 1 15809
0 15811 7 4 2 43206 60069
0 15812 7 3 2 44092 41224
0 15813 7 1 2 41011 63164
0 15814 7 1 2 59824 15813
0 15815 7 1 2 63160 15814
0 15816 5 1 1 15815
0 15817 7 1 2 15810 15816
0 15818 5 1 1 15817
0 15819 7 1 2 42129 52812
0 15820 7 1 2 15818 15819
0 15821 5 1 1 15820
0 15822 7 1 2 15807 15821
0 15823 5 1 1 15822
0 15824 7 1 2 42367 15823
0 15825 5 1 1 15824
0 15826 7 1 2 50484 59118
0 15827 7 2 2 63161 15826
0 15828 7 1 2 49506 50370
0 15829 5 2 1 15828
0 15830 7 1 2 51613 63169
0 15831 7 1 2 63167 15830
0 15832 5 1 1 15831
0 15833 7 1 2 15825 15832
0 15834 5 1 1 15833
0 15835 7 1 2 42812 15834
0 15836 5 1 1 15835
0 15837 7 1 2 2554 62546
0 15838 5 1 1 15837
0 15839 7 1 2 42368 15838
0 15840 5 1 1 15839
0 15841 7 1 2 49507 61402
0 15842 5 1 1 15841
0 15843 7 1 2 60239 15842
0 15844 5 1 1 15843
0 15845 7 1 2 15840 15844
0 15846 5 1 1 15845
0 15847 7 1 2 44940 15846
0 15848 5 1 1 15847
0 15849 7 2 2 52676 51174
0 15850 7 1 2 63171 50133
0 15851 5 1 1 15850
0 15852 7 1 2 15848 15851
0 15853 5 1 1 15852
0 15854 7 1 2 46109 60409
0 15855 7 1 2 15853 15854
0 15856 5 1 1 15855
0 15857 7 1 2 15836 15856
0 15858 7 1 2 15803 15857
0 15859 7 1 2 15752 15858
0 15860 5 1 1 15859
0 15861 7 1 2 44784 15860
0 15862 5 1 1 15861
0 15863 7 1 2 40832 62917
0 15864 5 1 1 15863
0 15865 7 1 2 48635 59895
0 15866 5 1 1 15865
0 15867 7 1 2 15864 15866
0 15868 5 1 1 15867
0 15869 7 1 2 40612 15868
0 15870 5 1 1 15869
0 15871 7 1 2 47732 54715
0 15872 5 1 1 15871
0 15873 7 1 2 50583 53720
0 15874 5 1 1 15873
0 15875 7 1 2 15872 15874
0 15876 5 1 1 15875
0 15877 7 1 2 50193 51345
0 15878 7 1 2 15876 15877
0 15879 5 1 1 15878
0 15880 7 1 2 15870 15879
0 15881 5 1 1 15880
0 15882 7 1 2 41486 15881
0 15883 5 1 1 15882
0 15884 7 2 2 47585 60544
0 15885 7 1 2 63173 62558
0 15886 5 1 1 15885
0 15887 7 1 2 43709 48017
0 15888 5 1 1 15887
0 15889 7 1 2 237 15888
0 15890 5 1 1 15889
0 15891 7 1 2 47412 15890
0 15892 5 1 1 15891
0 15893 7 1 2 61463 15892
0 15894 5 1 1 15893
0 15895 7 1 2 40833 53189
0 15896 7 1 2 15894 15895
0 15897 5 1 1 15896
0 15898 7 1 2 15886 15897
0 15899 5 1 1 15898
0 15900 7 1 2 45293 15899
0 15901 5 1 1 15900
0 15902 7 1 2 15883 15901
0 15903 5 1 1 15902
0 15904 7 1 2 44941 15903
0 15905 5 1 1 15904
0 15906 7 1 2 49163 51416
0 15907 7 1 2 60122 15906
0 15908 5 1 1 15907
0 15909 7 1 2 15905 15908
0 15910 5 1 1 15909
0 15911 7 1 2 60278 15910
0 15912 5 1 1 15911
0 15913 7 1 2 43909 61055
0 15914 5 1 1 15913
0 15915 7 1 2 51247 15914
0 15916 5 1 1 15915
0 15917 7 1 2 54712 63168
0 15918 7 1 2 15916 15917
0 15919 5 1 1 15918
0 15920 7 1 2 15912 15919
0 15921 5 1 1 15920
0 15922 7 1 2 42813 15921
0 15923 5 1 1 15922
0 15924 7 2 2 43710 49835
0 15925 5 1 1 63175
0 15926 7 1 2 47342 61475
0 15927 5 1 1 15926
0 15928 7 1 2 15925 15927
0 15929 5 1 1 15928
0 15930 7 1 2 60240 15929
0 15931 5 1 1 15930
0 15932 7 1 2 41487 55899
0 15933 5 1 1 15932
0 15934 7 1 2 41959 55943
0 15935 5 1 1 15934
0 15936 7 1 2 45688 60878
0 15937 5 1 1 15936
0 15938 7 1 2 15935 15937
0 15939 5 1 1 15938
0 15940 7 1 2 51587 15939
0 15941 5 1 1 15940
0 15942 7 1 2 15933 15941
0 15943 7 1 2 15931 15942
0 15944 5 1 1 15943
0 15945 7 1 2 59461 15944
0 15946 5 1 1 15945
0 15947 7 2 2 42130 48490
0 15948 5 1 1 63177
0 15949 7 1 2 50194 63178
0 15950 7 1 2 61362 15949
0 15951 5 1 1 15950
0 15952 7 1 2 15946 15951
0 15953 5 1 1 15952
0 15954 7 1 2 44942 15953
0 15955 5 1 1 15954
0 15956 7 1 2 44660 47183
0 15957 7 1 2 54674 15956
0 15958 7 2 2 62077 60070
0 15959 7 1 2 63179 53039
0 15960 7 1 2 15957 15959
0 15961 5 1 1 15960
0 15962 7 1 2 15955 15961
0 15963 5 1 1 15962
0 15964 7 1 2 58306 15963
0 15965 5 1 1 15964
0 15966 7 1 2 42589 15965
0 15967 7 1 2 15923 15966
0 15968 7 1 2 15862 15967
0 15969 5 1 1 15968
0 15970 7 1 2 53423 62631
0 15971 5 1 1 15970
0 15972 7 1 2 51592 61403
0 15973 5 3 1 15972
0 15974 7 1 2 45460 51417
0 15975 7 1 2 63181 15974
0 15976 5 1 1 15975
0 15977 7 1 2 15971 15976
0 15978 5 1 1 15977
0 15979 7 1 2 62381 15978
0 15980 5 1 1 15979
0 15981 7 1 2 55793 62472
0 15982 7 1 2 60040 15981
0 15983 5 1 1 15982
0 15984 7 1 2 15980 15983
0 15985 5 1 1 15984
0 15986 7 1 2 59462 15985
0 15987 5 1 1 15986
0 15988 7 1 2 61286 48883
0 15989 7 1 2 61242 15988
0 15990 5 1 1 15989
0 15991 7 1 2 15987 15990
0 15992 5 1 1 15991
0 15993 7 1 2 44943 15992
0 15994 5 1 1 15993
0 15995 7 1 2 47733 56111
0 15996 5 1 1 15995
0 15997 7 1 2 54972 15996
0 15998 5 1 1 15997
0 15999 7 1 2 47343 59119
0 16000 7 1 2 63162 15999
0 16001 7 1 2 15998 16000
0 16002 5 1 1 16001
0 16003 7 1 2 15994 16002
0 16004 5 1 1 16003
0 16005 7 1 2 42814 16004
0 16006 5 1 1 16005
0 16007 7 1 2 50987 10766
0 16008 5 1 1 16007
0 16009 7 1 2 49134 16008
0 16010 5 1 1 16009
0 16011 7 1 2 41648 53041
0 16012 5 1 1 16011
0 16013 7 1 2 62644 50256
0 16014 7 1 2 16012 16013
0 16015 5 1 1 16014
0 16016 7 1 2 16010 16015
0 16017 5 1 1 16016
0 16018 7 4 2 41800 46110
0 16019 5 1 1 63184
0 16020 7 4 2 43207 63185
0 16021 7 1 2 44093 60385
0 16022 7 1 2 63188 16021
0 16023 7 1 2 16017 16022
0 16024 5 1 1 16023
0 16025 7 1 2 45920 16024
0 16026 7 1 2 16006 16025
0 16027 5 1 1 16026
0 16028 7 1 2 42969 16027
0 16029 7 1 2 15969 16028
0 16030 5 1 1 16029
0 16031 7 2 2 47051 59463
0 16032 5 1 1 63192
0 16033 7 1 2 44510 61630
0 16034 5 1 1 16033
0 16035 7 1 2 16032 16034
0 16036 5 1 1 16035
0 16037 7 1 2 55485 16036
0 16038 5 1 1 16037
0 16039 7 1 2 47086 60461
0 16040 7 1 2 61412 16039
0 16041 5 1 1 16040
0 16042 7 1 2 16038 16041
0 16043 5 1 1 16042
0 16044 7 1 2 52058 16043
0 16045 5 1 1 16044
0 16046 7 1 2 60279 61782
0 16047 5 1 1 16046
0 16048 7 1 2 59464 51138
0 16049 5 1 1 16048
0 16050 7 1 2 11491 16049
0 16051 7 1 2 16047 16050
0 16052 5 1 1 16051
0 16053 7 1 2 48869 16052
0 16054 5 1 1 16053
0 16055 7 1 2 16045 16054
0 16056 5 1 1 16055
0 16057 7 1 2 51696 55199
0 16058 7 1 2 16056 16057
0 16059 5 1 1 16058
0 16060 7 1 2 16030 16059
0 16061 5 1 1 16060
0 16062 7 1 2 46394 16061
0 16063 5 1 1 16062
0 16064 7 1 2 7149 62891
0 16065 5 9 1 16064
0 16066 7 1 2 40208 63038
0 16067 5 1 1 16066
0 16068 7 1 2 45294 59465
0 16069 5 1 1 16068
0 16070 7 1 2 61335 16069
0 16071 5 1 1 16070
0 16072 7 1 2 60770 16071
0 16073 5 1 1 16072
0 16074 7 1 2 16067 16073
0 16075 5 1 1 16074
0 16076 7 1 2 45461 16075
0 16077 5 1 1 16076
0 16078 7 2 2 62055 55670
0 16079 7 2 2 45295 46483
0 16080 7 1 2 61829 63205
0 16081 7 1 2 63203 16080
0 16082 5 1 1 16081
0 16083 7 1 2 16077 16082
0 16084 5 1 1 16083
0 16085 7 1 2 53208 16084
0 16086 5 1 1 16085
0 16087 7 1 2 62325 16086
0 16088 5 1 1 16087
0 16089 7 1 2 41356 16088
0 16090 5 1 1 16089
0 16091 7 2 2 42590 50437
0 16092 7 1 2 61045 63207
0 16093 5 1 1 16092
0 16094 7 1 2 52576 16093
0 16095 5 1 1 16094
0 16096 7 1 2 41357 16095
0 16097 5 1 1 16096
0 16098 7 1 2 56554 16097
0 16099 5 1 1 16098
0 16100 7 1 2 59466 16099
0 16101 5 1 1 16100
0 16102 7 1 2 47989 60566
0 16103 5 1 1 16102
0 16104 7 1 2 61444 16103
0 16105 5 1 1 16104
0 16106 7 1 2 40009 16105
0 16107 5 1 1 16106
0 16108 7 1 2 59586 16107
0 16109 5 1 1 16108
0 16110 7 1 2 52451 60280
0 16111 7 1 2 16109 16110
0 16112 5 1 1 16111
0 16113 7 1 2 16101 16112
0 16114 5 1 1 16113
0 16115 7 1 2 49652 16114
0 16116 5 1 1 16115
0 16117 7 1 2 55671 62331
0 16118 5 1 1 16117
0 16119 7 1 2 16116 16118
0 16120 7 1 2 16090 16119
0 16121 5 1 1 16120
0 16122 7 1 2 40384 16121
0 16123 5 1 1 16122
0 16124 7 1 2 62433 60016
0 16125 5 1 1 16124
0 16126 7 3 2 45689 56917
0 16127 7 1 2 55577 63209
0 16128 7 1 2 62031 16127
0 16129 5 1 1 16128
0 16130 7 1 2 16125 16129
0 16131 5 1 1 16130
0 16132 7 1 2 41358 16131
0 16133 5 1 1 16132
0 16134 7 4 2 45921 59523
0 16135 7 1 2 63212 63102
0 16136 5 1 1 16135
0 16137 7 1 2 16133 16136
0 16138 5 1 1 16137
0 16139 7 1 2 62033 16138
0 16140 5 1 1 16139
0 16141 7 3 2 44785 45095
0 16142 7 1 2 46484 63216
0 16143 7 1 2 53475 16142
0 16144 7 2 2 50030 46892
0 16145 7 2 2 40010 62018
0 16146 7 1 2 63219 63221
0 16147 7 1 2 16143 16146
0 16148 5 1 1 16147
0 16149 7 1 2 16140 16148
0 16150 7 1 2 16123 16149
0 16151 5 1 1 16150
0 16152 7 1 2 44094 16151
0 16153 5 1 1 16152
0 16154 7 4 2 42131 54270
0 16155 7 1 2 63223 8353
0 16156 5 1 1 16155
0 16157 7 1 2 61068 16156
0 16158 5 1 1 16157
0 16159 7 1 2 42369 16158
0 16160 5 1 1 16159
0 16161 7 1 2 49653 60440
0 16162 5 1 1 16161
0 16163 7 1 2 52895 16162
0 16164 5 1 1 16163
0 16165 7 1 2 51585 61404
0 16166 5 1 1 16165
0 16167 7 1 2 49587 16166
0 16168 5 1 1 16167
0 16169 7 1 2 50048 60758
0 16170 5 1 1 16169
0 16171 7 1 2 45922 16170
0 16172 7 1 2 16168 16171
0 16173 7 1 2 16164 16172
0 16174 5 1 1 16173
0 16175 7 1 2 44786 61049
0 16176 5 1 1 16175
0 16177 7 1 2 61051 16176
0 16178 5 1 1 16177
0 16179 7 1 2 45462 16178
0 16180 5 1 1 16179
0 16181 7 1 2 42591 61041
0 16182 7 1 2 16180 16181
0 16183 5 1 1 16182
0 16184 7 1 2 16174 16183
0 16185 5 1 1 16184
0 16186 7 1 2 16160 16185
0 16187 5 1 1 16186
0 16188 7 1 2 40834 16187
0 16189 5 1 1 16188
0 16190 7 1 2 52535 62514
0 16191 5 1 1 16190
0 16192 7 1 2 54511 16191
0 16193 5 3 1 16192
0 16194 7 1 2 52957 63227
0 16195 7 1 2 55644 16194
0 16196 5 1 1 16195
0 16197 7 3 2 48371 60667
0 16198 7 1 2 63230 52193
0 16199 7 1 2 49736 16198
0 16200 5 1 1 16199
0 16201 7 1 2 16196 16200
0 16202 5 1 1 16201
0 16203 7 1 2 42370 16202
0 16204 5 1 1 16203
0 16205 7 1 2 60901 60985
0 16206 7 1 2 51254 16205
0 16207 5 1 1 16206
0 16208 7 1 2 16204 16207
0 16209 7 1 2 16189 16208
0 16210 5 1 1 16209
0 16211 7 1 2 59467 16210
0 16212 5 1 1 16211
0 16213 7 1 2 16153 16212
0 16214 5 1 1 16213
0 16215 7 1 2 63194 16214
0 16216 5 1 1 16215
0 16217 7 6 2 45923 46255
0 16218 5 1 1 63233
0 16219 7 2 2 63234 61388
0 16220 7 1 2 56580 63239
0 16221 5 1 1 16220
0 16222 7 4 2 58721 59270
0 16223 7 1 2 57433 63241
0 16224 5 1 1 16223
0 16225 7 1 2 16221 16224
0 16226 5 1 1 16225
0 16227 7 1 2 42132 16226
0 16228 5 1 1 16227
0 16229 7 3 2 44787 50876
0 16230 7 1 2 63245 63242
0 16231 5 1 1 16230
0 16232 7 1 2 16228 16231
0 16233 5 1 1 16232
0 16234 7 1 2 41225 16233
0 16235 5 1 1 16234
0 16236 7 1 2 53008 63243
0 16237 7 1 2 62299 16236
0 16238 5 1 1 16237
0 16239 7 1 2 16235 16238
0 16240 5 1 1 16239
0 16241 7 1 2 41012 16240
0 16242 5 1 1 16241
0 16243 7 1 2 44257 53556
0 16244 7 1 2 60071 16243
0 16245 7 1 2 63240 16244
0 16246 5 1 1 16245
0 16247 7 1 2 16242 16246
0 16248 5 1 1 16247
0 16249 7 1 2 44095 16248
0 16250 5 1 1 16249
0 16251 7 2 2 48636 59292
0 16252 7 1 2 63093 63224
0 16253 7 1 2 63248 16252
0 16254 5 1 1 16253
0 16255 7 1 2 16250 16254
0 16256 5 1 1 16255
0 16257 7 1 2 42371 16256
0 16258 5 1 1 16257
0 16259 7 2 2 49588 52495
0 16260 7 3 2 51534 59935
0 16261 5 2 1 63252
0 16262 7 2 2 41013 63253
0 16263 7 1 2 45296 63257
0 16264 5 1 1 16263
0 16265 7 1 2 48063 63249
0 16266 5 1 1 16265
0 16267 7 1 2 16264 16266
0 16268 5 1 1 16267
0 16269 7 1 2 63250 16268
0 16270 5 1 1 16269
0 16271 7 1 2 16258 16270
0 16272 5 1 1 16271
0 16273 7 1 2 46111 16272
0 16274 5 1 1 16273
0 16275 7 1 2 51976 61498
0 16276 5 1 1 16275
0 16277 7 1 2 60567 55531
0 16278 7 1 2 62632 16277
0 16279 5 1 1 16278
0 16280 7 1 2 16276 16279
0 16281 5 1 1 16280
0 16282 7 3 2 44096 62371
0 16283 7 1 2 59178 63259
0 16284 7 1 2 16281 16283
0 16285 5 1 1 16284
0 16286 7 1 2 16274 16285
0 16287 5 1 1 16286
0 16288 7 1 2 46395 16287
0 16289 5 1 1 16288
0 16290 7 2 2 49654 53541
0 16291 7 2 2 63127 60011
0 16292 7 1 2 51919 63043
0 16293 7 1 2 63264 16292
0 16294 7 1 2 63262 16293
0 16295 5 1 1 16294
0 16296 7 1 2 43208 16295
0 16297 7 1 2 16289 16296
0 16298 5 1 1 16297
0 16299 7 4 2 42970 55050
0 16300 7 1 2 54316 62408
0 16301 5 1 1 16300
0 16302 7 1 2 52067 52574
0 16303 5 1 1 16302
0 16304 7 1 2 16301 16303
0 16305 5 1 1 16304
0 16306 7 1 2 40613 16305
0 16307 5 1 1 16306
0 16308 7 4 2 42372 53284
0 16309 5 1 1 63270
0 16310 7 1 2 55638 63271
0 16311 5 1 1 16310
0 16312 7 1 2 16307 16311
0 16313 5 1 1 16312
0 16314 7 1 2 42815 16313
0 16315 5 1 1 16314
0 16316 7 1 2 55391 60568
0 16317 5 1 1 16316
0 16318 7 1 2 16315 16317
0 16319 5 1 1 16318
0 16320 7 1 2 63266 16319
0 16321 5 1 1 16320
0 16322 7 2 2 50438 62056
0 16323 7 1 2 41488 62302
0 16324 7 1 2 63274 16323
0 16325 7 3 2 63235 50763
0 16326 7 1 2 62278 63276
0 16327 7 1 2 16324 16326
0 16328 5 1 1 16327
0 16329 7 1 2 16321 16328
0 16330 5 1 1 16329
0 16331 7 1 2 44097 16330
0 16332 5 1 1 16331
0 16333 7 1 2 40011 57558
0 16334 5 1 1 16333
0 16335 7 9 2 42592 48491
0 16336 5 5 1 63279
0 16337 7 1 2 40209 63280
0 16338 5 1 1 16337
0 16339 7 1 2 16334 16338
0 16340 5 1 1 16339
0 16341 7 4 2 59359 60338
0 16342 7 1 2 50764 63293
0 16343 7 1 2 16340 16342
0 16344 5 1 1 16343
0 16345 7 1 2 16332 16344
0 16346 5 1 1 16345
0 16347 7 1 2 44944 16346
0 16348 5 1 1 16347
0 16349 7 6 2 55051 57500
0 16350 5 1 1 63297
0 16351 7 3 2 60339 59279
0 16352 5 1 1 63303
0 16353 7 1 2 16350 16352
0 16354 5 2 1 16353
0 16355 7 2 2 46112 53009
0 16356 5 1 1 63308
0 16357 7 1 2 63309 60843
0 16358 5 1 1 16357
0 16359 7 2 2 56069 58240
0 16360 7 1 2 63310 55963
0 16361 5 1 1 16360
0 16362 7 1 2 16358 16361
0 16363 5 1 1 16362
0 16364 7 1 2 42593 16363
0 16365 5 1 1 16364
0 16366 7 1 2 53209 56070
0 16367 7 1 2 57582 16366
0 16368 5 1 1 16367
0 16369 7 1 2 16365 16368
0 16370 5 1 1 16369
0 16371 7 1 2 63306 16370
0 16372 5 1 1 16371
0 16373 7 6 2 56581 60340
0 16374 7 3 2 41111 45924
0 16375 7 2 2 42816 59880
0 16376 7 2 2 40012 42373
0 16377 7 1 2 63323 50698
0 16378 7 1 2 63321 16377
0 16379 5 1 1 16378
0 16380 7 1 2 45297 56945
0 16381 7 1 2 59902 16380
0 16382 5 1 1 16381
0 16383 7 1 2 16379 16382
0 16384 5 1 1 16383
0 16385 7 1 2 63318 16384
0 16386 5 1 1 16385
0 16387 7 1 2 56715 55200
0 16388 5 1 1 16387
0 16389 7 1 2 16386 16388
0 16390 5 1 1 16389
0 16391 7 1 2 40614 16390
0 16392 5 1 1 16391
0 16393 7 1 2 55557 61534
0 16394 7 1 2 63322 16393
0 16395 5 1 1 16394
0 16396 7 1 2 16392 16395
0 16397 5 1 1 16396
0 16398 7 1 2 63312 16397
0 16399 5 1 1 16398
0 16400 7 1 2 16372 16399
0 16401 7 1 2 16348 16400
0 16402 5 1 1 16401
0 16403 7 1 2 43102 16402
0 16404 5 1 1 16403
0 16405 7 2 2 55052 47783
0 16406 7 3 2 54271 48581
0 16407 7 1 2 63325 63327
0 16408 5 1 1 16407
0 16409 7 2 2 49655 52638
0 16410 7 2 2 56592 61366
0 16411 7 3 2 40210 45925
0 16412 7 1 2 63332 63334
0 16413 7 1 2 63330 16412
0 16414 5 1 1 16413
0 16415 7 1 2 16408 16414
0 16416 5 1 1 16415
0 16417 7 1 2 43103 16416
0 16418 5 1 1 16417
0 16419 7 1 2 41226 53599
0 16420 7 1 2 62019 63217
0 16421 7 1 2 16419 16420
0 16422 7 1 2 53607 16421
0 16423 5 1 1 16422
0 16424 7 1 2 16418 16423
0 16425 5 1 1 16424
0 16426 7 1 2 51046 16425
0 16427 5 1 1 16426
0 16428 7 2 2 43910 53608
0 16429 7 5 2 44788 57636
0 16430 7 1 2 63339 60915
0 16431 7 1 2 63337 16430
0 16432 5 1 1 16431
0 16433 7 1 2 16427 16432
0 16434 5 1 1 16433
0 16435 7 1 2 47465 16434
0 16436 5 1 1 16435
0 16437 7 1 2 44789 60012
0 16438 7 1 2 58836 16437
0 16439 5 1 1 16438
0 16440 7 5 2 40615 41112
0 16441 7 1 2 53285 63344
0 16442 7 1 2 59360 16441
0 16443 7 1 2 59651 16442
0 16444 5 1 1 16443
0 16445 7 1 2 16439 16444
0 16446 5 1 1 16445
0 16447 7 1 2 44258 16446
0 16448 5 1 1 16447
0 16449 7 1 2 41014 63218
0 16450 7 1 2 58776 16449
0 16451 5 1 1 16450
0 16452 7 1 2 16448 16451
0 16453 5 1 1 16452
0 16454 7 1 2 47586 60575
0 16455 7 1 2 16453 16454
0 16456 5 1 1 16455
0 16457 7 1 2 16436 16456
0 16458 5 1 1 16457
0 16459 7 1 2 49202 16458
0 16460 5 1 1 16459
0 16461 7 1 2 46485 16460
0 16462 7 1 2 16404 16461
0 16463 5 1 1 16462
0 16464 7 1 2 49508 16463
0 16465 7 1 2 16298 16464
0 16466 5 1 1 16465
0 16467 7 1 2 16216 16466
0 16468 7 1 2 16063 16467
0 16469 7 1 2 15666 16468
0 16470 7 1 2 15298 16469
0 16471 5 1 1 16470
0 16472 7 1 2 49023 16471
0 16473 5 1 1 16472
0 16474 7 1 2 51697 63016
0 16475 5 1 1 16474
0 16476 7 1 2 43376 61304
0 16477 5 1 1 16476
0 16478 7 1 2 46845 51578
0 16479 5 1 1 16478
0 16480 7 1 2 16477 16479
0 16481 5 1 1 16480
0 16482 7 1 2 43711 16481
0 16483 5 1 1 16482
0 16484 7 1 2 61037 16483
0 16485 5 1 1 16484
0 16486 7 1 2 42133 16485
0 16487 5 1 1 16486
0 16488 7 1 2 55897 60041
0 16489 5 1 1 16488
0 16490 7 1 2 16487 16489
0 16491 5 1 1 16490
0 16492 7 1 2 41489 16491
0 16493 5 1 1 16492
0 16494 7 1 2 56179 63182
0 16495 5 1 1 16494
0 16496 7 1 2 60835 60840
0 16497 5 1 1 16496
0 16498 7 1 2 40211 16497
0 16499 5 1 1 16498
0 16500 7 1 2 6025 62592
0 16501 5 1 1 16500
0 16502 7 1 2 40013 16501
0 16503 5 1 1 16502
0 16504 7 1 2 16499 16503
0 16505 5 1 1 16504
0 16506 7 1 2 52958 16505
0 16507 5 1 1 16506
0 16508 7 1 2 16495 16507
0 16509 5 1 1 16508
0 16510 7 1 2 62479 16509
0 16511 5 1 1 16510
0 16512 7 1 2 61057 10959
0 16513 5 1 1 16512
0 16514 7 1 2 46846 49442
0 16515 5 1 1 16514
0 16516 7 1 2 41490 51014
0 16517 7 1 2 16515 16516
0 16518 7 1 2 61066 16517
0 16519 7 1 2 16513 16518
0 16520 5 1 1 16519
0 16521 7 1 2 44790 62550
0 16522 5 1 1 16521
0 16523 7 1 2 42374 16522
0 16524 7 1 2 16520 16523
0 16525 5 1 1 16524
0 16526 7 1 2 16511 16525
0 16527 7 1 2 16493 16526
0 16528 5 1 1 16527
0 16529 7 1 2 41649 16528
0 16530 5 1 1 16529
0 16531 7 2 2 54561 51657
0 16532 5 1 1 63349
0 16533 7 1 2 45690 63350
0 16534 5 1 1 16533
0 16535 7 1 2 16530 16534
0 16536 5 1 1 16535
0 16537 7 1 2 48109 16536
0 16538 5 1 1 16537
0 16539 7 1 2 43377 61467
0 16540 5 1 1 16539
0 16541 7 3 2 43911 51047
0 16542 5 1 1 63351
0 16543 7 1 2 47344 61469
0 16544 5 1 1 16543
0 16545 7 1 2 16542 16544
0 16546 7 1 2 16540 16545
0 16547 5 1 1 16546
0 16548 7 1 2 41491 16547
0 16549 5 1 1 16548
0 16550 7 1 2 62507 61394
0 16551 5 1 1 16550
0 16552 7 1 2 16549 16551
0 16553 5 1 1 16552
0 16554 7 1 2 56220 16553
0 16555 5 1 1 16554
0 16556 7 1 2 16538 16555
0 16557 5 1 1 16556
0 16558 7 1 2 40835 16557
0 16559 5 1 1 16558
0 16560 7 1 2 48492 48189
0 16561 5 2 1 16560
0 16562 7 1 2 48190 50568
0 16563 5 1 1 16562
0 16564 7 1 2 45691 48252
0 16565 5 1 1 16564
0 16566 7 1 2 16563 16565
0 16567 5 1 1 16566
0 16568 7 1 2 62062 16567
0 16569 5 1 1 16568
0 16570 7 1 2 63354 16569
0 16571 5 1 1 16570
0 16572 7 1 2 48680 16571
0 16573 5 1 1 16572
0 16574 7 3 2 49589 52639
0 16575 7 2 2 41650 52033
0 16576 7 1 2 61697 63359
0 16577 5 1 1 16576
0 16578 7 1 2 61708 50266
0 16579 5 1 1 16578
0 16580 7 1 2 47184 16579
0 16581 5 1 1 16580
0 16582 7 1 2 60893 63360
0 16583 5 1 1 16582
0 16584 7 1 2 16581 16583
0 16585 5 1 1 16584
0 16586 7 1 2 43378 16585
0 16587 5 1 1 16586
0 16588 7 1 2 16577 16587
0 16589 5 1 1 16588
0 16590 7 1 2 43547 16589
0 16591 5 1 1 16590
0 16592 7 1 2 41651 61693
0 16593 5 1 1 16592
0 16594 7 1 2 16591 16593
0 16595 5 1 1 16594
0 16596 7 1 2 43712 16595
0 16597 5 1 1 16596
0 16598 7 1 2 50264 62960
0 16599 5 1 1 16598
0 16600 7 1 2 16597 16599
0 16601 5 1 1 16600
0 16602 7 1 2 63356 16601
0 16603 5 1 1 16602
0 16604 7 1 2 16573 16603
0 16605 5 1 1 16604
0 16606 7 1 2 44098 16605
0 16607 5 1 1 16606
0 16608 7 1 2 48110 47857
0 16609 5 2 1 16608
0 16610 7 1 2 44420 48253
0 16611 5 1 1 16610
0 16612 7 1 2 51647 16611
0 16613 5 2 1 16612
0 16614 7 1 2 43379 63363
0 16615 5 1 1 16614
0 16616 7 1 2 63361 16615
0 16617 5 1 1 16616
0 16618 7 2 2 62438 49730
0 16619 7 1 2 49802 63365
0 16620 7 1 2 60241 16619
0 16621 7 1 2 16617 16620
0 16622 5 1 1 16621
0 16623 7 1 2 16607 16622
0 16624 7 1 2 16559 16623
0 16625 5 1 1 16624
0 16626 7 1 2 57253 16625
0 16627 5 1 1 16626
0 16628 7 1 2 16475 16627
0 16629 5 1 1 16628
0 16630 7 1 2 53891 16629
0 16631 5 1 1 16630
0 16632 7 1 2 57478 61111
0 16633 5 1 1 16632
0 16634 7 1 2 49943 62892
0 16635 5 1 1 16634
0 16636 7 1 2 46847 63195
0 16637 7 1 2 16635 16636
0 16638 5 1 1 16637
0 16639 7 1 2 16633 16638
0 16640 5 1 1 16639
0 16641 7 1 2 42134 16640
0 16642 5 1 1 16641
0 16643 7 1 2 54603 53140
0 16644 7 1 2 55528 16643
0 16645 5 1 1 16644
0 16646 7 1 2 16642 16645
0 16647 5 1 1 16646
0 16648 7 1 2 44511 16647
0 16649 5 1 1 16648
0 16650 7 4 2 42135 54604
0 16651 7 2 2 46716 61112
0 16652 7 2 2 46113 63371
0 16653 7 1 2 63367 63373
0 16654 5 1 1 16653
0 16655 7 1 2 16649 16654
0 16656 5 1 1 16655
0 16657 7 1 2 43548 16656
0 16658 5 1 1 16657
0 16659 7 1 2 58156 62914
0 16660 5 1 1 16659
0 16661 7 1 2 16658 16660
0 16662 5 1 1 16661
0 16663 7 1 2 49443 16662
0 16664 5 1 1 16663
0 16665 7 1 2 56659 58185
0 16666 5 1 1 16665
0 16667 7 1 2 62893 16666
0 16668 5 2 1 16667
0 16669 7 1 2 47734 63375
0 16670 5 1 1 16669
0 16671 7 1 2 47656 46717
0 16672 7 1 2 63196 16671
0 16673 5 1 1 16672
0 16674 7 1 2 16670 16673
0 16675 5 1 1 16674
0 16676 7 1 2 43380 16675
0 16677 5 1 1 16676
0 16678 7 1 2 58106 62895
0 16679 5 1 1 16678
0 16680 7 1 2 16677 16679
0 16681 5 1 1 16680
0 16682 7 1 2 42136 16681
0 16683 5 1 1 16682
0 16684 7 1 2 52803 62900
0 16685 5 1 1 16684
0 16686 7 1 2 16683 16685
0 16687 5 1 1 16686
0 16688 7 1 2 48769 16687
0 16689 5 1 1 16688
0 16690 7 1 2 51748 62889
0 16691 5 1 1 16690
0 16692 7 1 2 45463 50827
0 16693 5 2 1 16692
0 16694 7 1 2 58636 63377
0 16695 5 1 1 16694
0 16696 7 1 2 16691 16695
0 16697 5 1 1 16696
0 16698 7 1 2 47657 16697
0 16699 5 1 1 16698
0 16700 7 1 2 47587 51373
0 16701 5 1 1 16700
0 16702 7 1 2 49717 16701
0 16703 7 1 2 63376 16702
0 16704 5 1 1 16703
0 16705 7 1 2 63197 53158
0 16706 5 1 1 16705
0 16707 7 1 2 57479 47858
0 16708 7 1 2 63378 16707
0 16709 5 1 1 16708
0 16710 7 1 2 16706 16709
0 16711 7 1 2 16704 16710
0 16712 7 1 2 16699 16711
0 16713 5 1 1 16712
0 16714 7 1 2 49444 16713
0 16715 5 1 1 16714
0 16716 7 1 2 16689 16715
0 16717 5 1 1 16716
0 16718 7 1 2 42375 16717
0 16719 5 1 1 16718
0 16720 7 1 2 54605 58241
0 16721 7 1 2 60698 16720
0 16722 5 1 1 16721
0 16723 7 1 2 16719 16722
0 16724 7 1 2 16664 16723
0 16725 5 1 1 16724
0 16726 7 3 2 45054 46486
0 16727 7 1 2 63379 57151
0 16728 7 1 2 16725 16727
0 16729 5 1 1 16728
0 16730 7 1 2 16631 16729
0 16731 5 1 1 16730
0 16732 7 1 2 42594 16731
0 16733 5 1 1 16732
0 16734 7 1 2 53443 62594
0 16735 5 1 1 16734
0 16736 7 1 2 45298 49164
0 16737 7 1 2 61733 16736
0 16738 5 1 1 16737
0 16739 7 1 2 16735 16738
0 16740 5 1 1 16739
0 16741 7 1 2 41492 16740
0 16742 5 1 1 16741
0 16743 7 1 2 48448 50411
0 16744 5 1 1 16743
0 16745 7 1 2 47588 59778
0 16746 7 1 2 62542 16745
0 16747 7 1 2 16744 16746
0 16748 5 1 1 16747
0 16749 7 1 2 16742 16748
0 16750 5 1 1 16749
0 16751 7 1 2 45464 16750
0 16752 5 1 1 16751
0 16753 7 1 2 51255 61128
0 16754 5 1 1 16753
0 16755 7 1 2 11178 16754
0 16756 5 1 1 16755
0 16757 7 1 2 42376 16756
0 16758 5 1 1 16757
0 16759 7 1 2 49656 10239
0 16760 5 1 1 16759
0 16761 7 1 2 43549 16760
0 16762 5 1 1 16761
0 16763 7 1 2 4216 16762
0 16764 5 1 1 16763
0 16765 7 1 2 48770 16764
0 16766 5 1 1 16765
0 16767 7 1 2 41960 56312
0 16768 5 1 1 16767
0 16769 7 1 2 49657 59889
0 16770 7 1 2 16768 16769
0 16771 7 1 2 61226 16770
0 16772 5 1 1 16771
0 16773 7 1 2 52896 16772
0 16774 5 1 1 16773
0 16775 7 1 2 16766 16774
0 16776 7 1 2 16758 16775
0 16777 5 1 1 16776
0 16778 7 1 2 40836 16777
0 16779 5 1 1 16778
0 16780 7 1 2 54911 60937
0 16781 5 1 1 16780
0 16782 7 1 2 43550 16781
0 16783 5 1 1 16782
0 16784 7 1 2 43713 46872
0 16785 5 2 1 16784
0 16786 7 1 2 63382 61035
0 16787 7 1 2 16783 16786
0 16788 5 1 1 16787
0 16789 7 1 2 48884 16788
0 16790 5 1 1 16789
0 16791 7 1 2 60986 58815
0 16792 5 1 1 16791
0 16793 7 1 2 62561 16792
0 16794 7 1 2 16790 16793
0 16795 5 1 1 16794
0 16796 7 1 2 51048 16795
0 16797 5 1 1 16796
0 16798 7 1 2 16779 16797
0 16799 5 1 1 16798
0 16800 7 1 2 41652 16799
0 16801 5 1 1 16800
0 16802 7 1 2 16752 16801
0 16803 5 1 1 16802
0 16804 7 1 2 61663 16803
0 16805 5 1 1 16804
0 16806 7 2 2 40837 61740
0 16807 7 1 2 52403 53359
0 16808 5 1 1 16807
0 16809 7 1 2 48560 61275
0 16810 5 1 1 16809
0 16811 7 1 2 41653 16810
0 16812 5 1 1 16811
0 16813 7 1 2 44945 48561
0 16814 5 4 1 16813
0 16815 7 1 2 43381 63386
0 16816 7 1 2 16812 16815
0 16817 5 1 1 16816
0 16818 7 1 2 16808 16817
0 16819 5 1 1 16818
0 16820 7 1 2 47052 16819
0 16821 5 1 1 16820
0 16822 7 1 2 41654 52365
0 16823 5 1 1 16822
0 16824 7 1 2 52149 16823
0 16825 5 1 1 16824
0 16826 7 1 2 52284 16825
0 16827 5 1 1 16826
0 16828 7 1 2 50457 62439
0 16829 7 1 2 50397 16828
0 16830 5 1 1 16829
0 16831 7 1 2 16827 16830
0 16832 7 1 2 16821 16831
0 16833 5 1 1 16832
0 16834 7 1 2 52034 16833
0 16835 5 1 1 16834
0 16836 7 1 2 50134 54947
0 16837 5 1 1 16836
0 16838 7 1 2 52150 16837
0 16839 5 2 1 16838
0 16840 7 1 2 46978 63390
0 16841 5 1 1 16840
0 16842 7 1 2 55890 53360
0 16843 5 1 1 16842
0 16844 7 1 2 16841 16843
0 16845 5 1 1 16844
0 16846 7 1 2 42137 16845
0 16847 5 1 1 16846
0 16848 7 1 2 1730 63391
0 16849 5 1 1 16848
0 16850 7 1 2 16847 16849
0 16851 7 1 2 16835 16850
0 16852 5 1 1 16851
0 16853 7 1 2 63384 16852
0 16854 5 1 1 16853
0 16855 7 1 2 16805 16854
0 16856 5 1 1 16855
0 16857 7 1 2 42971 16856
0 16858 5 1 1 16857
0 16859 7 2 2 57202 51535
0 16860 7 1 2 49590 51175
0 16861 7 1 2 63392 16860
0 16862 5 1 1 16861
0 16863 7 1 2 41655 61659
0 16864 7 1 2 62620 16863
0 16865 5 1 1 16864
0 16866 7 1 2 16862 16865
0 16867 5 1 1 16866
0 16868 7 1 2 40385 16867
0 16869 5 1 1 16868
0 16870 7 1 2 51049 54797
0 16871 5 1 1 16870
0 16872 7 1 2 51836 16871
0 16873 7 1 2 51808 16872
0 16874 5 1 1 16873
0 16875 7 1 2 41961 16874
0 16876 5 1 1 16875
0 16877 7 1 2 1117 51903
0 16878 5 1 1 16877
0 16879 7 1 2 48771 16878
0 16880 5 1 1 16879
0 16881 7 1 2 58473 62912
0 16882 5 1 1 16881
0 16883 7 1 2 47971 53181
0 16884 5 1 1 16883
0 16885 7 1 2 58070 16884
0 16886 7 1 2 16882 16885
0 16887 7 1 2 16880 16886
0 16888 7 1 2 16876 16887
0 16889 5 1 1 16888
0 16890 7 1 2 49591 16889
0 16891 5 1 1 16890
0 16892 7 1 2 53353 16891
0 16893 5 1 1 16892
0 16894 7 1 2 63393 16893
0 16895 5 1 1 16894
0 16896 7 1 2 16869 16895
0 16897 5 1 1 16896
0 16898 7 1 2 49354 16897
0 16899 5 1 1 16898
0 16900 7 1 2 46114 16899
0 16901 7 1 2 16858 16900
0 16902 5 1 1 16901
0 16903 7 2 2 42972 61953
0 16904 7 1 2 61741 60822
0 16905 5 2 1 16904
0 16906 7 2 2 62256 62310
0 16907 7 1 2 50439 57254
0 16908 7 1 2 63398 16907
0 16909 5 1 1 16908
0 16910 7 1 2 63396 16909
0 16911 5 1 1 16910
0 16912 7 1 2 63394 16911
0 16913 5 1 1 16912
0 16914 7 3 2 44791 42138
0 16915 5 1 1 63400
0 16916 7 3 2 43912 63401
0 16917 5 1 1 63403
0 16918 7 1 2 47921 61129
0 16919 7 1 2 61461 16918
0 16920 5 1 1 16919
0 16921 7 1 2 16917 16920
0 16922 5 1 1 16921
0 16923 7 1 2 42377 16922
0 16924 5 1 1 16923
0 16925 7 1 2 49951 60906
0 16926 5 2 1 16925
0 16927 7 1 2 63406 63024
0 16928 5 1 1 16927
0 16929 7 1 2 52897 16928
0 16930 5 1 1 16929
0 16931 7 1 2 16924 16930
0 16932 5 1 1 16931
0 16933 7 1 2 53892 57966
0 16934 7 1 2 16932 16933
0 16935 5 1 1 16934
0 16936 7 1 2 16913 16935
0 16937 5 1 1 16936
0 16938 7 1 2 44946 16937
0 16939 5 1 1 16938
0 16940 7 1 2 50328 50229
0 16941 7 1 2 54973 16940
0 16942 5 1 1 16941
0 16943 7 1 2 45692 53424
0 16944 5 1 1 16943
0 16945 7 1 2 16942 16944
0 16946 5 1 1 16945
0 16947 7 1 2 40014 16946
0 16948 5 1 1 16947
0 16949 7 2 2 41359 53010
0 16950 7 1 2 49861 63408
0 16951 5 1 1 16950
0 16952 7 1 2 51614 62625
0 16953 5 1 1 16952
0 16954 7 1 2 16951 16953
0 16955 5 1 1 16954
0 16956 7 1 2 45299 16955
0 16957 5 1 1 16956
0 16958 7 1 2 16948 16957
0 16959 5 1 1 16958
0 16960 7 1 2 45465 16959
0 16961 5 1 1 16960
0 16962 7 2 2 52325 62534
0 16963 7 1 2 63410 61421
0 16964 5 1 1 16963
0 16965 7 1 2 50607 48681
0 16966 7 1 2 56723 16965
0 16967 7 1 2 60539 16966
0 16968 5 1 1 16967
0 16969 7 1 2 16964 16968
0 16970 5 1 1 16969
0 16971 7 1 2 41227 16970
0 16972 5 1 1 16971
0 16973 7 1 2 16961 16972
0 16974 5 1 1 16973
0 16975 7 1 2 61664 16974
0 16976 5 1 1 16975
0 16977 7 6 2 50087 61876
0 16978 7 1 2 57203 63412
0 16979 7 1 2 14907 16978
0 16980 5 1 1 16979
0 16981 7 1 2 16976 16980
0 16982 5 1 1 16981
0 16983 7 1 2 41656 16982
0 16984 5 1 1 16983
0 16985 7 1 2 53893 61518
0 16986 7 1 2 53190 16985
0 16987 7 1 2 61414 16986
0 16988 7 1 2 63103 16987
0 16989 5 1 1 16988
0 16990 7 1 2 16984 16989
0 16991 5 1 1 16990
0 16992 7 1 2 42973 16991
0 16993 5 1 1 16992
0 16994 7 1 2 16939 16993
0 16995 5 1 1 16994
0 16996 7 1 2 40838 16995
0 16997 5 1 1 16996
0 16998 7 4 2 46487 54606
0 16999 7 4 2 44099 61162
0 17000 7 5 2 63418 63422
0 17001 7 1 2 45693 52115
0 17002 5 1 1 17001
0 17003 7 1 2 53405 17002
0 17004 5 1 1 17003
0 17005 7 1 2 52720 17004
0 17006 5 1 1 17005
0 17007 7 1 2 63426 17006
0 17008 5 1 1 17007
0 17009 7 7 2 43209 53638
0 17010 7 4 2 53894 63431
0 17011 7 3 2 42378 48493
0 17012 7 1 2 63442 61415
0 17013 7 1 2 63438 17012
0 17014 7 1 2 55630 17013
0 17015 5 1 1 17014
0 17016 7 1 2 17008 17015
0 17017 5 1 1 17016
0 17018 7 1 2 41657 17017
0 17019 5 1 1 17018
0 17020 7 1 2 2174 10678
0 17021 5 1 1 17020
0 17022 7 2 2 55179 60507
0 17023 5 2 1 63445
0 17024 7 1 2 50485 63446
0 17025 7 1 2 17021 17024
0 17026 5 1 1 17025
0 17027 7 1 2 42817 17026
0 17028 7 1 2 17019 17027
0 17029 7 1 2 16997 17028
0 17030 5 1 1 17029
0 17031 7 1 2 45926 17030
0 17032 7 1 2 16902 17031
0 17033 5 1 1 17032
0 17034 7 1 2 48111 48359
0 17035 5 2 1 17034
0 17036 7 1 2 48637 56221
0 17037 5 1 1 17036
0 17038 7 1 2 63449 17037
0 17039 5 1 1 17038
0 17040 7 1 2 61492 62289
0 17041 5 1 1 17040
0 17042 7 1 2 45466 54463
0 17043 5 1 1 17042
0 17044 7 1 2 17041 17043
0 17045 5 1 1 17044
0 17046 7 1 2 17039 17045
0 17047 5 1 1 17046
0 17048 7 1 2 45467 53146
0 17049 5 1 1 17048
0 17050 7 1 2 52748 17049
0 17051 5 1 1 17050
0 17052 7 1 2 41228 17051
0 17053 5 1 1 17052
0 17054 7 1 2 55672 53147
0 17055 5 1 1 17054
0 17056 7 1 2 17053 17055
0 17057 5 1 1 17056
0 17058 7 1 2 61422 17057
0 17059 5 1 1 17058
0 17060 7 2 2 49658 48341
0 17061 7 1 2 59848 55607
0 17062 7 1 2 63451 17061
0 17063 5 1 1 17062
0 17064 7 2 2 42818 62636
0 17065 7 1 2 52398 52152
0 17066 7 1 2 63453 17065
0 17067 5 1 1 17066
0 17068 7 1 2 17063 17067
0 17069 5 1 1 17068
0 17070 7 1 2 45300 17069
0 17071 5 1 1 17070
0 17072 7 1 2 17059 17071
0 17073 5 1 1 17072
0 17074 7 1 2 45927 17073
0 17075 5 1 1 17074
0 17076 7 2 2 41962 47017
0 17077 5 1 1 63455
0 17078 7 1 2 40015 62300
0 17079 5 1 1 17078
0 17080 7 1 2 17077 17079
0 17081 5 2 1 17080
0 17082 7 1 2 42379 50734
0 17083 7 1 2 63457 17082
0 17084 5 1 1 17083
0 17085 7 1 2 16532 17084
0 17086 5 1 1 17085
0 17087 7 1 2 53825 17086
0 17088 5 1 1 17087
0 17089 7 1 2 17075 17088
0 17090 5 1 1 17089
0 17091 7 1 2 40839 17090
0 17092 5 1 1 17091
0 17093 7 1 2 63452 63458
0 17094 5 1 1 17093
0 17095 7 3 2 41493 63345
0 17096 7 2 2 52326 63459
0 17097 7 1 2 63462 63454
0 17098 5 1 1 17097
0 17099 7 1 2 17094 17098
0 17100 5 1 1 17099
0 17101 7 1 2 45928 17100
0 17102 5 1 1 17101
0 17103 7 2 2 45468 53826
0 17104 7 1 2 63464 54562
0 17105 5 1 1 17104
0 17106 7 1 2 17102 17105
0 17107 5 1 1 17106
0 17108 7 1 2 49165 17107
0 17109 5 1 1 17108
0 17110 7 1 2 17092 17109
0 17111 5 1 1 17110
0 17112 7 1 2 42974 17111
0 17113 5 1 1 17112
0 17114 7 1 2 17047 17113
0 17115 5 1 1 17114
0 17116 7 1 2 61665 17115
0 17117 5 1 1 17116
0 17118 7 2 2 40016 55572
0 17119 7 1 2 63466 58342
0 17120 5 1 1 17119
0 17121 7 1 2 3740 17120
0 17122 5 1 1 17121
0 17123 7 1 2 47784 17122
0 17124 5 1 1 17123
0 17125 7 3 2 41658 51050
0 17126 5 1 1 63468
0 17127 7 1 2 55496 50398
0 17128 5 1 1 17127
0 17129 7 1 2 17126 17128
0 17130 5 1 1 17129
0 17131 7 1 2 63335 17130
0 17132 5 1 1 17131
0 17133 7 3 2 42595 61804
0 17134 7 1 2 41659 63471
0 17135 5 1 1 17134
0 17136 7 1 2 17132 17135
0 17137 5 1 1 17136
0 17138 7 1 2 42819 17137
0 17139 5 1 1 17138
0 17140 7 2 2 53827 50399
0 17141 5 1 1 63474
0 17142 7 1 2 40212 63475
0 17143 5 1 1 17142
0 17144 7 1 2 17139 17143
0 17145 5 1 1 17144
0 17146 7 1 2 45301 17145
0 17147 5 1 1 17146
0 17148 7 1 2 17124 17147
0 17149 5 1 1 17148
0 17150 7 1 2 40616 17149
0 17151 5 1 1 17150
0 17152 7 1 2 52549 53148
0 17153 5 1 1 17152
0 17154 7 1 2 3666 17153
0 17155 5 1 1 17154
0 17156 7 1 2 52179 53191
0 17157 7 1 2 17155 17156
0 17158 5 1 1 17157
0 17159 7 1 2 17151 17158
0 17160 5 1 1 17159
0 17161 7 1 2 41113 17160
0 17162 5 1 1 17161
0 17163 7 1 2 55653 53069
0 17164 5 1 1 17163
0 17165 7 1 2 17162 17164
0 17166 5 1 1 17165
0 17167 7 1 2 61959 17166
0 17168 5 1 1 17167
0 17169 7 6 2 46256 53828
0 17170 7 1 2 49135 55000
0 17171 7 1 2 57134 17170
0 17172 7 1 2 63476 17171
0 17173 5 2 1 17172
0 17174 7 1 2 53015 62290
0 17175 5 1 1 17174
0 17176 7 1 2 52496 54457
0 17177 5 1 1 17176
0 17178 7 1 2 17175 17177
0 17179 5 1 1 17178
0 17180 7 1 2 41114 17179
0 17181 5 1 1 17180
0 17182 7 6 2 40213 44792
0 17183 7 1 2 53580 63484
0 17184 7 1 2 54443 17183
0 17185 5 1 1 17184
0 17186 7 1 2 17181 17185
0 17187 5 1 1 17186
0 17188 7 1 2 40017 17187
0 17189 5 1 1 17188
0 17190 7 1 2 55497 62589
0 17191 7 1 2 55953 17190
0 17192 5 1 1 17191
0 17193 7 1 2 17189 17192
0 17194 5 1 1 17193
0 17195 7 1 2 48268 17194
0 17196 5 1 1 17195
0 17197 7 1 2 63482 17196
0 17198 7 1 2 17168 17197
0 17199 5 1 1 17198
0 17200 7 1 2 61742 17199
0 17201 5 1 1 17200
0 17202 7 1 2 17117 17201
0 17203 5 1 1 17202
0 17204 7 1 2 49509 17203
0 17205 5 1 1 17204
0 17206 7 4 2 47589 50371
0 17207 5 3 1 63490
0 17208 7 1 2 63491 63228
0 17209 5 1 1 17208
0 17210 7 1 2 58337 49940
0 17211 5 1 1 17210
0 17212 7 1 2 17209 17211
0 17213 5 1 1 17212
0 17214 7 1 2 44793 17213
0 17215 5 1 1 17214
0 17216 7 1 2 49941 60895
0 17217 5 1 1 17216
0 17218 7 1 2 17215 17217
0 17219 5 1 1 17218
0 17220 7 1 2 61666 17219
0 17221 5 1 1 17220
0 17222 7 1 2 54317 53592
0 17223 5 1 1 17222
0 17224 7 1 2 61146 17223
0 17225 5 1 1 17224
0 17226 7 1 2 41963 17225
0 17227 5 1 1 17226
0 17228 7 1 2 54318 61228
0 17229 5 1 1 17228
0 17230 7 1 2 17227 17229
0 17231 5 1 1 17230
0 17232 7 1 2 17231 63385
0 17233 5 1 1 17232
0 17234 7 1 2 17221 17233
0 17235 5 1 1 17234
0 17236 7 1 2 42139 17235
0 17237 5 1 1 17236
0 17238 7 2 2 54319 62102
0 17239 7 1 2 61638 63497
0 17240 5 1 1 17239
0 17241 7 3 2 44207 50088
0 17242 7 2 2 63499 61712
0 17243 7 2 2 47658 50383
0 17244 5 3 1 63504
0 17245 7 1 2 63506 58709
0 17246 5 1 1 17245
0 17247 7 1 2 63502 17246
0 17248 5 1 1 17247
0 17249 7 1 2 53895 47659
0 17250 7 1 2 62652 17249
0 17251 5 1 1 17250
0 17252 7 1 2 17248 17251
0 17253 5 1 1 17252
0 17254 7 1 2 44661 17253
0 17255 5 1 1 17254
0 17256 7 1 2 17240 17255
0 17257 5 1 1 17256
0 17258 7 1 2 43714 17257
0 17259 5 1 1 17258
0 17260 7 1 2 61645 63498
0 17261 5 1 1 17260
0 17262 7 1 2 17259 17261
0 17263 5 1 1 17262
0 17264 7 1 2 40840 17263
0 17265 5 1 1 17264
0 17266 7 1 2 17237 17265
0 17267 5 1 1 17266
0 17268 7 1 2 42380 17267
0 17269 5 1 1 17268
0 17270 7 2 2 47413 49592
0 17271 5 1 1 63509
0 17272 7 1 2 51706 49151
0 17273 5 1 1 17272
0 17274 7 1 2 17271 17273
0 17275 5 1 1 17274
0 17276 7 1 2 45929 17275
0 17277 5 1 1 17276
0 17278 7 1 2 50363 60675
0 17279 5 1 1 17278
0 17280 7 1 2 17277 17279
0 17281 5 1 1 17280
0 17282 7 1 2 61667 17281
0 17283 5 1 1 17282
0 17284 7 1 2 49731 61718
0 17285 7 1 2 51781 17284
0 17286 5 1 1 17285
0 17287 7 1 2 17283 17286
0 17288 5 1 1 17287
0 17289 7 1 2 43715 17288
0 17290 5 1 1 17289
0 17291 7 2 2 61721 56450
0 17292 7 2 2 59660 63208
0 17293 5 1 1 63513
0 17294 7 2 2 45930 49916
0 17295 7 1 2 47414 63515
0 17296 5 1 1 17295
0 17297 7 1 2 17293 17296
0 17298 5 1 1 17297
0 17299 7 1 2 63511 17298
0 17300 5 1 1 17299
0 17301 7 1 2 17290 17300
0 17302 5 1 1 17301
0 17303 7 1 2 40841 17302
0 17304 5 1 1 17303
0 17305 7 2 2 57204 50512
0 17306 7 1 2 55312 60598
0 17307 7 1 2 63517 17306
0 17308 5 1 1 17307
0 17309 7 1 2 56829 62696
0 17310 7 1 2 62956 17309
0 17311 5 1 1 17310
0 17312 7 1 2 17308 17311
0 17313 5 1 1 17312
0 17314 7 1 2 60569 17313
0 17315 5 1 1 17314
0 17316 7 4 2 56883 57205
0 17317 7 1 2 54260 54918
0 17318 7 1 2 63519 17317
0 17319 5 1 1 17318
0 17320 7 1 2 17315 17319
0 17321 5 1 1 17320
0 17322 7 1 2 49659 17321
0 17323 5 1 1 17322
0 17324 7 4 2 52536 52623
0 17325 5 2 1 63523
0 17326 7 2 2 52399 62118
0 17327 7 1 2 50440 63529
0 17328 7 1 2 61722 17327
0 17329 5 1 1 17328
0 17330 7 1 2 63397 17329
0 17331 5 1 1 17330
0 17332 7 1 2 63524 17331
0 17333 5 1 1 17332
0 17334 7 1 2 17323 17333
0 17335 5 1 1 17334
0 17336 7 1 2 44100 17335
0 17337 5 1 1 17336
0 17338 7 1 2 17304 17337
0 17339 7 1 2 17269 17338
0 17340 5 1 1 17339
0 17341 7 1 2 48269 17340
0 17342 5 1 1 17341
0 17343 7 1 2 52489 9750
0 17344 5 1 1 17343
0 17345 7 1 2 63427 17344
0 17346 5 1 1 17345
0 17347 7 2 2 55427 61796
0 17348 7 2 2 57255 50006
0 17349 7 1 2 53234 63533
0 17350 7 1 2 63531 17349
0 17351 5 1 1 17350
0 17352 7 8 2 46257 57206
0 17353 7 1 2 52452 63535
0 17354 7 1 2 61163 17353
0 17355 5 1 1 17354
0 17356 7 1 2 17351 17355
0 17357 5 1 1 17356
0 17358 7 1 2 44101 17357
0 17359 5 1 1 17358
0 17360 7 1 2 40842 54974
0 17361 5 1 1 17360
0 17362 7 1 2 12639 17361
0 17363 5 2 1 17362
0 17364 7 1 2 63543 61493
0 17365 5 1 1 17364
0 17366 7 2 2 45469 50973
0 17367 7 1 2 63545 56336
0 17368 5 1 1 17367
0 17369 7 1 2 17365 17368
0 17370 5 1 1 17369
0 17371 7 1 2 52606 61668
0 17372 7 1 2 17370 17371
0 17373 5 1 1 17372
0 17374 7 1 2 17359 17373
0 17375 5 1 1 17374
0 17376 7 1 2 60570 17375
0 17377 5 1 1 17376
0 17378 7 1 2 17346 17377
0 17379 5 1 1 17378
0 17380 7 1 2 60530 17379
0 17381 5 1 1 17380
0 17382 7 1 2 60789 49684
0 17383 5 1 1 17382
0 17384 7 1 2 45694 61761
0 17385 5 1 1 17384
0 17386 7 1 2 17383 17385
0 17387 5 1 1 17386
0 17388 7 1 2 47018 17387
0 17389 5 1 1 17388
0 17390 7 1 2 60790 48682
0 17391 5 1 1 17390
0 17392 7 1 2 17389 17391
0 17393 5 1 1 17392
0 17394 7 1 2 49660 17393
0 17395 5 1 1 17394
0 17396 7 1 2 50561 52968
0 17397 5 1 1 17396
0 17398 7 1 2 56716 60913
0 17399 5 1 1 17398
0 17400 7 1 2 17397 17399
0 17401 5 1 1 17400
0 17402 7 1 2 45302 17401
0 17403 5 1 1 17402
0 17404 7 1 2 3367 17403
0 17405 5 1 1 17404
0 17406 7 1 2 53235 17405
0 17407 5 1 1 17406
0 17408 7 1 2 17395 17407
0 17409 5 1 1 17408
0 17410 7 1 2 46115 17409
0 17411 5 1 1 17410
0 17412 7 1 2 52550 50441
0 17413 5 1 1 17412
0 17414 7 1 2 14131 17413
0 17415 5 1 1 17414
0 17416 7 1 2 55237 61954
0 17417 7 1 2 17415 17416
0 17418 5 1 1 17417
0 17419 7 1 2 17411 17418
0 17420 5 1 1 17419
0 17421 7 1 2 63439 17420
0 17422 5 1 1 17421
0 17423 7 1 2 54607 62944
0 17424 7 1 2 60623 17423
0 17425 7 1 2 52128 17424
0 17426 5 1 1 17425
0 17427 7 1 2 17422 17426
0 17428 5 1 1 17427
0 17429 7 1 2 49203 17428
0 17430 5 1 1 17429
0 17431 7 1 2 17381 17430
0 17432 7 1 2 17342 17431
0 17433 7 1 2 17205 17432
0 17434 7 1 2 17033 17433
0 17435 7 1 2 16733 17434
0 17436 5 1 1 17435
0 17437 7 1 2 55053 17436
0 17438 5 1 1 17437
0 17439 7 1 2 16473 17438
0 17440 7 1 2 15014 17439
0 17441 7 1 2 11377 17440
0 17442 5 1 1 17441
0 17443 7 1 2 58545 17442
0 17444 5 1 1 17443
0 17445 7 2 2 40018 59137
0 17446 5 1 1 63547
0 17447 7 1 2 61436 17446
0 17448 5 4 1 17447
0 17449 7 2 2 43210 63549
0 17450 5 1 1 63553
0 17451 7 1 2 61546 63222
0 17452 5 1 1 17451
0 17453 7 1 2 17450 17452
0 17454 5 1 1 17453
0 17455 7 1 2 55737 17454
0 17456 5 1 1 17455
0 17457 7 1 2 60367 63213
0 17458 5 1 1 17457
0 17459 7 1 2 17456 17458
0 17460 5 1 1 17459
0 17461 7 1 2 41660 17460
0 17462 5 1 1 17461
0 17463 7 2 2 45931 61893
0 17464 7 1 2 63555 62015
0 17465 5 1 1 17464
0 17466 7 1 2 17462 17465
0 17467 5 1 1 17466
0 17468 7 1 2 53896 17467
0 17469 5 1 1 17468
0 17470 7 2 2 46624 57256
0 17471 5 3 1 63557
0 17472 7 1 2 58888 57376
0 17473 5 1 1 17472
0 17474 7 1 2 63559 17473
0 17475 5 2 1 17474
0 17476 7 1 2 40019 63562
0 17477 5 2 1 17476
0 17478 7 1 2 60281 60742
0 17479 5 1 1 17478
0 17480 7 1 2 63564 17479
0 17481 5 1 1 17480
0 17482 7 1 2 55738 57525
0 17483 7 1 2 17481 17482
0 17484 5 1 1 17483
0 17485 7 1 2 17469 17484
0 17486 5 1 1 17485
0 17487 7 1 2 40843 17486
0 17488 5 1 1 17487
0 17489 7 1 2 51221 61904
0 17490 5 1 1 17489
0 17491 7 1 2 17488 17490
0 17492 5 1 1 17491
0 17493 7 1 2 40386 17492
0 17494 5 1 1 17493
0 17495 7 2 2 42596 48064
0 17496 7 2 2 54159 60282
0 17497 7 1 2 48494 63568
0 17498 5 2 1 17497
0 17499 7 12 2 43104 48912
0 17500 7 1 2 63572 57377
0 17501 5 1 1 17500
0 17502 7 1 2 61686 17501
0 17503 5 2 1 17502
0 17504 7 1 2 55054 63584
0 17505 5 1 1 17504
0 17506 7 1 2 40214 61553
0 17507 5 1 1 17506
0 17508 7 1 2 61589 17507
0 17509 7 1 2 17505 17508
0 17510 5 1 1 17509
0 17511 7 1 2 40020 17510
0 17512 5 1 1 17511
0 17513 7 1 2 62043 17512
0 17514 5 1 1 17513
0 17515 7 1 2 50652 17514
0 17516 5 1 1 17515
0 17517 7 1 2 63570 17516
0 17518 5 1 1 17517
0 17519 7 1 2 63566 17518
0 17520 5 1 1 17519
0 17521 7 1 2 17494 17520
0 17522 5 1 1 17521
0 17523 7 1 2 42975 17522
0 17524 5 1 1 17523
0 17525 7 2 2 54872 51536
0 17526 7 3 2 40021 41758
0 17527 7 4 2 57030 63588
0 17528 5 2 1 63591
0 17529 7 1 2 60283 63592
0 17530 5 1 1 17529
0 17531 7 2 2 61590 17530
0 17532 5 2 1 63597
0 17533 7 5 2 46488 57176
0 17534 7 3 2 48913 63601
0 17535 5 1 1 63606
0 17536 7 1 2 61687 17535
0 17537 5 2 1 17536
0 17538 7 1 2 55055 63609
0 17539 5 1 1 17538
0 17540 7 1 2 63598 17539
0 17541 5 2 1 17540
0 17542 7 4 2 40215 50348
0 17543 7 1 2 63611 63613
0 17544 5 1 1 17543
0 17545 7 5 2 41759 62119
0 17546 7 2 2 58413 63617
0 17547 7 1 2 60352 63622
0 17548 5 1 1 17547
0 17549 7 1 2 17544 17548
0 17550 5 1 1 17549
0 17551 7 1 2 49661 17550
0 17552 5 1 1 17551
0 17553 7 1 2 63571 17552
0 17554 5 1 1 17553
0 17555 7 1 2 63586 17554
0 17556 5 1 1 17555
0 17557 7 1 2 17524 17556
0 17558 5 1 1 17557
0 17559 7 1 2 42820 17558
0 17560 5 1 1 17559
0 17561 7 2 2 60576 62760
0 17562 7 1 2 57569 56226
0 17563 7 1 2 63624 17562
0 17564 7 1 2 63214 17563
0 17565 5 1 1 17564
0 17566 7 2 2 61857 62669
0 17567 7 4 2 46489 53639
0 17568 7 2 2 45096 53829
0 17569 7 1 2 63628 63632
0 17570 7 1 2 63626 17569
0 17571 5 1 1 17570
0 17572 7 1 2 17565 17571
0 17573 5 1 1 17572
0 17574 7 1 2 43913 17573
0 17575 5 1 1 17574
0 17576 7 1 2 40022 57426
0 17577 5 1 1 17576
0 17578 7 1 2 59996 17577
0 17579 5 3 1 17578
0 17580 7 4 2 40387 44259
0 17581 7 1 2 63637 61942
0 17582 5 1 1 17581
0 17583 7 1 2 62044 17582
0 17584 5 1 1 17583
0 17585 7 1 2 63634 17584
0 17586 5 1 1 17585
0 17587 7 1 2 44102 51270
0 17588 5 1 1 17587
0 17589 7 1 2 59997 17588
0 17590 5 6 1 17589
0 17591 7 1 2 40216 63641
0 17592 7 1 2 63612 17591
0 17593 5 1 1 17592
0 17594 7 1 2 17586 17593
0 17595 5 1 1 17594
0 17596 7 1 2 45695 17595
0 17597 5 1 1 17596
0 17598 7 1 2 63607 63642
0 17599 5 1 1 17598
0 17600 7 1 2 17599 63447
0 17601 5 1 1 17600
0 17602 7 1 2 55056 17601
0 17603 5 1 1 17602
0 17604 7 1 2 44260 61547
0 17605 7 3 2 63618 17604
0 17606 7 1 2 63643 63647
0 17607 5 1 1 17606
0 17608 7 1 2 60508 59213
0 17609 5 2 1 17608
0 17610 7 1 2 17607 63650
0 17611 7 1 2 17603 17610
0 17612 5 1 1 17611
0 17613 7 1 2 54651 17612
0 17614 5 1 1 17613
0 17615 7 1 2 17597 17614
0 17616 5 1 1 17615
0 17617 7 1 2 55238 17616
0 17618 5 1 1 17617
0 17619 7 1 2 17575 17618
0 17620 5 1 1 17619
0 17621 7 1 2 44794 17620
0 17622 5 1 1 17621
0 17623 7 4 2 42597 53640
0 17624 7 2 2 40217 50538
0 17625 7 2 2 63652 63656
0 17626 5 1 1 63658
0 17627 7 2 2 53286 54608
0 17628 7 8 2 40023 41661
0 17629 7 1 2 50349 63662
0 17630 7 1 2 63660 17629
0 17631 5 1 1 17630
0 17632 7 1 2 17626 17631
0 17633 5 1 1 17632
0 17634 7 1 2 40844 17633
0 17635 5 1 1 17634
0 17636 7 2 2 56717 51729
0 17637 7 2 2 53641 57135
0 17638 7 1 2 63670 63672
0 17639 5 1 1 17638
0 17640 7 1 2 17635 17639
0 17641 5 1 1 17640
0 17642 7 1 2 48914 17641
0 17643 5 1 1 17642
0 17644 7 1 2 62396 62510
0 17645 5 1 1 17644
0 17646 7 1 2 40845 55313
0 17647 5 1 1 17646
0 17648 7 1 2 17645 17647
0 17649 5 1 1 17648
0 17650 7 3 2 43105 50007
0 17651 7 1 2 57726 63674
0 17652 7 1 2 17649 17651
0 17653 5 1 1 17652
0 17654 7 1 2 17643 17653
0 17655 5 1 1 17654
0 17656 7 1 2 46625 17655
0 17657 5 1 1 17656
0 17658 7 1 2 60155 52136
0 17659 7 1 2 54661 17658
0 17660 5 1 1 17659
0 17661 7 1 2 61994 63595
0 17662 5 1 1 17661
0 17663 7 1 2 53287 50350
0 17664 7 1 2 57232 17663
0 17665 7 1 2 17662 17664
0 17666 5 1 1 17665
0 17667 7 1 2 17660 17666
0 17668 5 1 1 17667
0 17669 7 1 2 40846 17668
0 17670 5 1 1 17669
0 17671 7 1 2 41494 57727
0 17672 7 1 2 59924 17671
0 17673 7 1 2 63673 17672
0 17674 5 1 1 17673
0 17675 7 1 2 17670 17674
0 17676 5 1 1 17675
0 17677 7 1 2 55057 17676
0 17678 5 1 1 17677
0 17679 7 6 2 61541 59349
0 17680 5 1 1 63677
0 17681 7 1 2 53288 57956
0 17682 7 1 2 63614 17681
0 17683 7 1 2 63678 17682
0 17684 5 1 1 17683
0 17685 7 1 2 17678 17684
0 17686 7 1 2 17657 17685
0 17687 5 1 1 17686
0 17688 7 1 2 40617 17687
0 17689 5 1 1 17688
0 17690 7 1 2 60247 51486
0 17691 7 1 2 63659 17690
0 17692 5 1 1 17691
0 17693 7 1 2 62270 56337
0 17694 7 1 2 63244 17693
0 17695 7 1 2 61996 17694
0 17696 5 1 1 17695
0 17697 7 1 2 17692 17696
0 17698 7 1 2 17689 17697
0 17699 5 1 1 17698
0 17700 7 1 2 43211 17699
0 17701 5 1 1 17700
0 17702 7 2 2 40024 62812
0 17703 5 1 1 63683
0 17704 7 1 2 63684 63615
0 17705 5 1 1 17704
0 17706 7 2 2 40388 58999
0 17707 7 1 2 63685 62853
0 17708 5 1 1 17707
0 17709 7 1 2 17705 17708
0 17710 5 1 1 17709
0 17711 7 1 2 57501 17710
0 17712 5 1 1 17711
0 17713 7 1 2 63573 50417
0 17714 7 1 2 63304 17713
0 17715 5 1 1 17714
0 17716 7 1 2 17712 17715
0 17717 5 1 1 17716
0 17718 7 3 2 45932 46490
0 17719 7 1 2 48495 63687
0 17720 7 1 2 17717 17719
0 17721 5 1 1 17720
0 17722 7 1 2 17701 17721
0 17723 5 1 1 17722
0 17724 7 1 2 46116 17723
0 17725 5 1 1 17724
0 17726 7 1 2 17622 17725
0 17727 7 1 2 17560 17726
0 17728 5 1 1 17727
0 17729 7 1 2 41229 17728
0 17730 5 1 1 17729
0 17731 7 2 2 48400 51327
0 17732 7 1 2 53063 63503
0 17733 5 1 1 17732
0 17734 7 2 2 40389 56441
0 17735 7 1 2 53457 62104
0 17736 7 1 2 63692 17735
0 17737 5 1 1 17736
0 17738 7 1 2 17733 17737
0 17739 5 1 1 17738
0 17740 7 1 2 55058 17739
0 17741 5 1 1 17740
0 17742 7 2 2 61713 59217
0 17743 7 3 2 40618 61929
0 17744 7 2 2 62120 63696
0 17745 7 1 2 63694 63699
0 17746 5 1 1 17745
0 17747 7 2 2 60402 60743
0 17748 5 1 1 63701
0 17749 7 2 2 41015 51436
0 17750 7 1 2 45933 56884
0 17751 7 1 2 63703 17750
0 17752 7 1 2 63702 17751
0 17753 5 1 1 17752
0 17754 7 1 2 17746 17753
0 17755 7 1 2 17741 17754
0 17756 5 1 1 17755
0 17757 7 1 2 63690 17756
0 17758 5 1 1 17757
0 17759 7 1 2 55059 62105
0 17760 7 1 2 63477 17759
0 17761 7 1 2 57732 17760
0 17762 5 1 1 17761
0 17763 7 1 2 59271 60098
0 17764 7 1 2 62372 17763
0 17765 7 6 2 43914 57015
0 17766 7 1 2 57299 63705
0 17767 7 1 2 17764 17766
0 17768 5 1 1 17767
0 17769 7 1 2 17762 17768
0 17770 7 1 2 17758 17769
0 17771 7 1 2 17730 17770
0 17772 5 1 1 17771
0 17773 7 1 2 45470 17772
0 17774 5 1 1 17773
0 17775 7 2 2 47785 60509
0 17776 7 2 2 49662 63711
0 17777 7 1 2 51051 55180
0 17778 7 1 2 63713 17777
0 17779 5 1 1 17778
0 17780 7 2 2 50202 57257
0 17781 7 2 2 55332 56442
0 17782 7 1 2 63715 63717
0 17783 5 1 1 17782
0 17784 7 3 2 62251 61423
0 17785 7 1 2 61743 63719
0 17786 5 1 1 17785
0 17787 7 1 2 17783 17786
0 17788 5 1 1 17787
0 17789 7 1 2 63663 61960
0 17790 7 1 2 17788 17789
0 17791 5 1 1 17790
0 17792 7 1 2 17779 17791
0 17793 5 1 1 17792
0 17794 7 1 2 55239 17793
0 17795 5 1 1 17794
0 17796 7 1 2 52382 59250
0 17797 7 1 2 58509 17796
0 17798 7 1 2 63712 17797
0 17799 5 1 1 17798
0 17800 7 1 2 17795 17799
0 17801 5 1 1 17800
0 17802 7 1 2 55060 17801
0 17803 5 1 1 17802
0 17804 7 4 2 47786 51052
0 17805 5 1 1 63722
0 17806 7 1 2 57967 51393
0 17807 7 2 2 58671 62991
0 17808 5 1 1 63726
0 17809 7 1 2 58652 63727
0 17810 7 1 2 17806 17809
0 17811 5 1 1 17810
0 17812 7 1 2 59989 63648
0 17813 5 1 1 17812
0 17814 7 1 2 63651 17813
0 17815 5 1 1 17814
0 17816 7 1 2 42821 60961
0 17817 7 1 2 17815 17816
0 17818 5 1 1 17817
0 17819 7 1 2 17811 17818
0 17820 5 1 1 17819
0 17821 7 1 2 63723 17820
0 17822 5 1 1 17821
0 17823 7 1 2 50203 62373
0 17824 7 2 2 43212 52607
0 17825 7 2 2 60072 56765
0 17826 7 1 2 63728 63730
0 17827 7 1 2 17823 17826
0 17828 5 1 1 17827
0 17829 7 5 2 44947 45097
0 17830 7 1 2 46258 56918
0 17831 7 2 2 63732 17830
0 17832 7 1 2 61930 53259
0 17833 7 1 2 63737 17832
0 17834 5 1 1 17833
0 17835 7 1 2 17828 17834
0 17836 5 1 1 17835
0 17837 7 1 2 56071 54160
0 17838 7 1 2 17836 17837
0 17839 5 1 1 17838
0 17840 7 1 2 17822 17839
0 17841 7 1 2 17803 17840
0 17842 7 1 2 17774 17841
0 17843 5 1 1 17842
0 17844 7 1 2 41360 17843
0 17845 5 1 1 17844
0 17846 7 1 2 60477 15338
0 17847 5 4 1 17846
0 17848 7 1 2 48562 61445
0 17849 5 1 1 17848
0 17850 7 2 2 55587 17849
0 17851 5 1 1 63743
0 17852 7 2 2 50351 63744
0 17853 5 1 1 63745
0 17854 7 1 2 63739 63746
0 17855 5 1 1 17854
0 17856 7 1 2 60284 58242
0 17857 5 1 1 17856
0 17858 7 1 2 60360 17857
0 17859 5 2 1 17858
0 17860 7 1 2 50807 63747
0 17861 5 1 1 17860
0 17862 7 1 2 17855 17861
0 17863 5 1 1 17862
0 17864 7 1 2 42598 17863
0 17865 5 1 1 17864
0 17866 7 2 2 50280 52959
0 17867 5 1 1 63749
0 17868 7 1 2 61287 63616
0 17869 5 1 1 17868
0 17870 7 1 2 60361 17869
0 17871 5 2 1 17870
0 17872 7 1 2 63750 63751
0 17873 5 1 1 17872
0 17874 7 1 2 49593 15065
0 17875 5 1 1 17874
0 17876 7 1 2 40390 61321
0 17877 7 1 2 17875 17876
0 17878 5 1 1 17877
0 17879 7 1 2 17873 17878
0 17880 5 1 1 17879
0 17881 7 1 2 55240 17880
0 17882 5 1 1 17881
0 17883 7 1 2 17865 17882
0 17884 5 1 1 17883
0 17885 7 1 2 46259 17884
0 17886 5 1 1 17885
0 17887 7 1 2 45471 53431
0 17888 7 1 2 53252 17887
0 17889 7 1 2 57591 17888
0 17890 7 1 2 63752 17889
0 17891 5 1 1 17890
0 17892 7 1 2 17886 17891
0 17893 5 1 1 17892
0 17894 7 1 2 41662 17893
0 17895 5 1 1 17894
0 17896 7 1 2 42822 63272
0 17897 5 1 1 17896
0 17898 7 1 2 8032 17897
0 17899 5 1 1 17898
0 17900 7 1 2 40619 17899
0 17901 5 1 1 17900
0 17902 7 1 2 17901 17141
0 17903 5 1 1 17902
0 17904 7 1 2 40391 46626
0 17905 7 1 2 62761 17904
0 17906 7 1 2 61442 17905
0 17907 7 1 2 17903 17906
0 17908 5 1 1 17907
0 17909 7 1 2 17895 17908
0 17910 5 1 1 17909
0 17911 7 1 2 40847 17910
0 17912 5 1 1 17911
0 17913 7 1 2 46686 62382
0 17914 5 1 1 17913
0 17915 7 1 2 56091 56231
0 17916 5 1 1 17915
0 17917 7 1 2 17914 17916
0 17918 5 1 1 17917
0 17919 7 5 2 48496 46627
0 17920 7 1 2 50281 56645
0 17921 7 1 2 62762 17920
0 17922 7 1 2 63753 17921
0 17923 7 1 2 17918 17922
0 17924 5 1 1 17923
0 17925 7 1 2 17912 17924
0 17926 5 1 1 17925
0 17927 7 1 2 43106 17926
0 17928 5 1 1 17927
0 17929 7 2 2 63288 63527
0 17930 5 3 1 63758
0 17931 7 1 2 58498 63485
0 17932 5 1 1 17931
0 17933 7 1 2 50282 55739
0 17934 5 1 1 17933
0 17935 7 1 2 17932 17934
0 17936 5 1 1 17935
0 17937 7 1 2 41230 17936
0 17938 5 1 1 17937
0 17939 7 1 2 63759 17938
0 17940 5 1 1 17939
0 17941 7 1 2 45696 17940
0 17942 5 1 1 17941
0 17943 7 1 2 42599 54853
0 17944 5 1 1 17943
0 17945 7 1 2 17942 17944
0 17946 5 1 1 17945
0 17947 7 9 2 41016 59272
0 17948 7 7 2 42976 57258
0 17949 7 1 2 63772 56425
0 17950 7 1 2 63763 17949
0 17951 7 1 2 17946 17950
0 17952 5 1 1 17951
0 17953 7 1 2 17928 17952
0 17954 5 1 1 17953
0 17955 7 1 2 40025 17954
0 17956 5 1 1 17955
0 17957 7 1 2 51410 17851
0 17958 5 1 1 17957
0 17959 7 1 2 57807 17958
0 17960 5 1 1 17959
0 17961 7 1 2 57880 17960
0 17962 5 1 1 17961
0 17963 7 1 2 42600 17962
0 17964 5 1 1 17963
0 17965 7 1 2 57791 6022
0 17966 5 1 1 17965
0 17967 7 1 2 45934 51537
0 17968 7 1 2 62963 17967
0 17969 7 1 2 17966 17968
0 17970 5 1 1 17969
0 17971 7 1 2 17964 17970
0 17972 5 1 1 17971
0 17973 7 1 2 60285 17972
0 17974 5 1 1 17973
0 17975 7 2 2 58566 63729
0 17976 7 2 2 51233 63779
0 17977 7 1 2 51580 63123
0 17978 7 1 2 63781 17977
0 17979 5 1 1 17978
0 17980 7 1 2 17974 17979
0 17981 5 1 1 17980
0 17982 7 1 2 40392 17981
0 17983 5 1 1 17982
0 17984 7 1 2 54848 56466
0 17985 5 1 1 17984
0 17986 7 1 2 56511 17985
0 17987 5 1 1 17986
0 17988 7 1 2 41017 63486
0 17989 7 1 2 63432 17988
0 17990 7 1 2 59370 17989
0 17991 7 1 2 17987 17990
0 17992 5 1 1 17991
0 17993 7 1 2 17983 17992
0 17994 5 1 1 17993
0 17995 7 1 2 45697 17994
0 17996 5 1 1 17995
0 17997 7 10 2 46396 59515
0 17998 5 7 1 63783
0 17999 7 1 2 55588 56551
0 18000 5 1 1 17999
0 18001 7 2 2 51394 61499
0 18002 7 1 2 42601 63800
0 18003 5 1 1 18002
0 18004 7 1 2 18000 18003
0 18005 5 1 1 18004
0 18006 7 1 2 63784 18005
0 18007 5 1 1 18006
0 18008 7 1 2 49663 56552
0 18009 5 1 1 18008
0 18010 7 1 2 40620 63472
0 18011 5 1 1 18010
0 18012 7 1 2 18009 18011
0 18013 5 1 1 18012
0 18014 7 1 2 48967 62397
0 18015 7 1 2 57289 18014
0 18016 7 1 2 18013 18015
0 18017 5 1 1 18016
0 18018 7 1 2 18007 18017
0 18019 5 1 1 18018
0 18020 7 1 2 49510 18019
0 18021 5 1 1 18020
0 18022 7 1 2 48065 50783
0 18023 5 1 1 18022
0 18024 7 2 2 46117 63644
0 18025 7 1 2 48497 63802
0 18026 5 1 1 18025
0 18027 7 1 2 18023 18026
0 18028 5 4 1 18027
0 18029 7 1 2 57259 63804
0 18030 5 1 1 18029
0 18031 7 2 2 51538 53011
0 18032 7 1 2 63008 63808
0 18033 5 1 1 18032
0 18034 7 1 2 18030 18033
0 18035 5 1 1 18034
0 18036 7 1 2 62964 50352
0 18037 7 1 2 18035 18036
0 18038 5 1 1 18037
0 18039 7 1 2 63602 57502
0 18040 5 1 1 18039
0 18041 7 1 2 63793 18040
0 18042 5 2 1 18041
0 18043 7 1 2 55589 54696
0 18044 7 1 2 63810 18043
0 18045 5 1 1 18044
0 18046 7 1 2 45935 18045
0 18047 7 1 2 18038 18046
0 18048 5 1 1 18047
0 18049 7 1 2 2271 3125
0 18050 5 1 1 18049
0 18051 7 1 2 51395 18050
0 18052 5 1 1 18051
0 18053 7 1 2 17853 18052
0 18054 5 1 1 18053
0 18055 7 1 2 63785 18054
0 18056 5 1 1 18055
0 18057 7 1 2 56983 50513
0 18058 5 1 1 18057
0 18059 7 1 2 53002 50353
0 18060 7 1 2 62063 18059
0 18061 5 1 1 18060
0 18062 7 1 2 18058 18061
0 18063 5 1 1 18062
0 18064 7 1 2 57227 62398
0 18065 7 1 2 18063 18064
0 18066 5 1 1 18065
0 18067 7 1 2 42602 18066
0 18068 7 1 2 18056 18067
0 18069 5 1 1 18068
0 18070 7 1 2 40218 18069
0 18071 7 1 2 18048 18070
0 18072 5 1 1 18071
0 18073 7 1 2 18021 18072
0 18074 5 1 1 18073
0 18075 7 1 2 55061 18074
0 18076 5 1 1 18075
0 18077 7 5 2 44261 59047
0 18078 7 2 2 63812 62980
0 18079 7 1 2 54261 56984
0 18080 7 1 2 63817 18079
0 18081 5 1 1 18080
0 18082 7 1 2 18076 18081
0 18083 7 1 2 17996 18082
0 18084 7 1 2 17956 18083
0 18085 5 1 1 18084
0 18086 7 1 2 49024 18085
0 18087 5 1 1 18086
0 18088 7 2 2 46118 61839
0 18089 7 1 2 44208 63819
0 18090 5 1 1 18089
0 18091 7 2 2 42823 56443
0 18092 7 1 2 51053 63821
0 18093 5 1 1 18092
0 18094 7 1 2 18090 18093
0 18095 5 1 1 18094
0 18096 7 1 2 40219 18095
0 18097 5 1 1 18096
0 18098 7 1 2 61500 63822
0 18099 5 1 1 18098
0 18100 7 1 2 18097 18099
0 18101 5 1 1 18100
0 18102 7 1 2 42603 18101
0 18103 5 1 1 18102
0 18104 7 1 2 1305 53082
0 18105 5 3 1 18104
0 18106 7 2 2 53427 63823
0 18107 7 1 2 57452 63826
0 18108 5 1 1 18107
0 18109 7 1 2 18103 18108
0 18110 5 1 1 18109
0 18111 7 1 2 46260 18110
0 18112 5 1 1 18111
0 18113 7 2 2 53289 55428
0 18114 7 1 2 59904 63828
0 18115 7 1 2 56997 18114
0 18116 5 1 1 18115
0 18117 7 1 2 18112 18116
0 18118 5 1 1 18117
0 18119 7 1 2 61723 18118
0 18120 5 1 1 18119
0 18121 7 1 2 63714 58343
0 18122 5 1 1 18121
0 18123 7 7 2 57207 59247
0 18124 7 1 2 51158 53012
0 18125 7 1 2 63830 18124
0 18126 5 1 1 18125
0 18127 7 1 2 18122 18126
0 18128 5 1 1 18127
0 18129 7 1 2 49025 18128
0 18130 5 1 1 18129
0 18131 7 1 2 48498 53830
0 18132 5 2 1 18131
0 18133 7 1 2 55498 57516
0 18134 5 1 1 18133
0 18135 7 1 2 63837 18134
0 18136 5 1 1 18135
0 18137 7 7 2 40026 44209
0 18138 7 1 2 63839 57411
0 18139 7 1 2 57290 18138
0 18140 7 1 2 18136 18139
0 18141 5 1 1 18140
0 18142 7 1 2 18130 18141
0 18143 7 1 2 18120 18142
0 18144 5 1 1 18143
0 18145 7 1 2 55062 18144
0 18146 5 1 1 18145
0 18147 7 1 2 54077 56617
0 18148 5 1 1 18147
0 18149 7 2 2 40027 50653
0 18150 7 1 2 57945 56431
0 18151 7 1 2 63846 18150
0 18152 5 1 1 18151
0 18153 7 1 2 18148 18152
0 18154 5 1 1 18153
0 18155 7 1 2 47019 18154
0 18156 5 1 1 18155
0 18157 7 2 2 58567 51437
0 18158 7 1 2 50659 63848
0 18159 5 1 1 18158
0 18160 7 1 2 18156 18159
0 18161 5 1 1 18160
0 18162 7 1 2 40959 18161
0 18163 5 1 1 18162
0 18164 7 1 2 56784 63413
0 18165 7 1 2 50514 18164
0 18166 5 1 1 18165
0 18167 7 1 2 18163 18166
0 18168 5 1 1 18167
0 18169 7 1 2 42977 18168
0 18170 5 1 1 18169
0 18171 7 1 2 48977 56653
0 18172 5 1 1 18171
0 18173 7 1 2 5189 18172
0 18174 5 1 1 18173
0 18175 7 1 2 57788 18174
0 18176 5 1 1 18175
0 18177 7 1 2 18170 18176
0 18178 5 1 1 18177
0 18179 7 1 2 42604 18178
0 18180 5 1 1 18179
0 18181 7 1 2 48112 56444
0 18182 5 1 1 18181
0 18183 7 1 2 48499 58598
0 18184 5 1 1 18183
0 18185 7 1 2 18182 18184
0 18186 5 1 1 18185
0 18187 7 1 2 56841 54863
0 18188 7 1 2 55673 48782
0 18189 7 1 2 18187 18188
0 18190 7 1 2 18186 18189
0 18191 5 1 1 18190
0 18192 7 1 2 18180 18191
0 18193 5 1 1 18192
0 18194 7 1 2 60286 18193
0 18195 5 1 1 18194
0 18196 7 1 2 51165 17805
0 18197 5 1 1 18196
0 18198 7 1 2 18197 63849
0 18199 5 1 1 18198
0 18200 7 1 2 53095 54685
0 18201 7 1 2 61840 18200
0 18202 5 1 1 18201
0 18203 7 1 2 18199 18202
0 18204 5 1 1 18203
0 18205 7 1 2 44210 18204
0 18206 5 1 1 18205
0 18207 7 2 2 43107 62121
0 18208 7 1 2 45055 63820
0 18209 5 1 1 18208
0 18210 7 1 2 885 18209
0 18211 5 1 1 18210
0 18212 7 1 2 63850 18211
0 18213 5 1 1 18212
0 18214 7 1 2 18206 18213
0 18215 5 1 1 18214
0 18216 7 1 2 46261 18215
0 18217 5 1 1 18216
0 18218 7 1 2 48113 61997
0 18219 7 1 2 61841 18218
0 18220 5 1 1 18219
0 18221 7 1 2 42605 18220
0 18222 7 1 2 18217 18221
0 18223 5 1 1 18222
0 18224 7 7 2 40220 46397
0 18225 7 1 2 52865 63852
0 18226 5 1 1 18225
0 18227 7 1 2 40028 54552
0 18228 5 1 1 18227
0 18229 7 1 2 18226 18228
0 18230 5 1 1 18229
0 18231 7 1 2 44211 63824
0 18232 7 1 2 18230 18231
0 18233 5 1 1 18232
0 18234 7 1 2 57031 10195
0 18235 7 1 2 50021 18234
0 18236 7 1 2 53072 18235
0 18237 5 1 1 18236
0 18238 7 1 2 18233 18237
0 18239 5 1 1 18238
0 18240 7 1 2 45472 18239
0 18241 5 1 1 18240
0 18242 7 1 2 63414 63853
0 18243 7 1 2 56998 18242
0 18244 5 1 1 18243
0 18245 7 1 2 18241 18244
0 18246 5 1 1 18245
0 18247 7 1 2 48783 18246
0 18248 5 1 1 18247
0 18249 7 2 2 49664 48349
0 18250 7 1 2 53983 63859
0 18251 5 1 1 18250
0 18252 7 1 2 45936 18251
0 18253 7 1 2 18248 18252
0 18254 5 1 1 18253
0 18255 7 1 2 59468 18254
0 18256 7 1 2 18223 18255
0 18257 5 1 1 18256
0 18258 7 1 2 52960 60462
0 18259 7 1 2 60830 18258
0 18260 5 1 1 18259
0 18261 7 1 2 53847 55507
0 18262 5 1 1 18261
0 18263 7 1 2 57172 61986
0 18264 7 1 2 18262 18263
0 18265 5 1 1 18264
0 18266 7 1 2 18260 18265
0 18267 5 1 1 18266
0 18268 7 1 2 63851 18267
0 18269 5 1 1 18268
0 18270 7 1 2 45098 49594
0 18271 7 1 2 59387 58594
0 18272 7 1 2 18270 18271
0 18273 7 1 2 50515 18272
0 18274 5 1 1 18273
0 18275 7 1 2 40960 46119
0 18276 7 1 2 49665 18275
0 18277 7 1 2 62741 18276
0 18278 7 1 2 55063 18277
0 18279 7 1 2 61836 18278
0 18280 5 1 1 18279
0 18281 7 1 2 18274 18280
0 18282 5 1 1 18281
0 18283 7 1 2 42606 18282
0 18284 5 1 1 18283
0 18285 7 1 2 62311 62923
0 18286 7 1 2 63827 18285
0 18287 5 1 1 18286
0 18288 7 1 2 18284 18287
0 18289 5 1 1 18288
0 18290 7 1 2 46398 18289
0 18291 5 1 1 18290
0 18292 7 1 2 18269 18291
0 18293 5 1 1 18292
0 18294 7 1 2 52879 18293
0 18295 5 1 1 18294
0 18296 7 1 2 18257 18295
0 18297 7 1 2 18195 18296
0 18298 7 1 2 18146 18297
0 18299 5 1 1 18298
0 18300 7 1 2 49511 18299
0 18301 5 1 1 18300
0 18302 7 2 2 63340 60599
0 18303 7 1 2 62515 62641
0 18304 7 1 2 63861 18303
0 18305 5 1 1 18304
0 18306 7 1 2 61154 58595
0 18307 7 2 2 62750 18306
0 18308 5 1 1 63863
0 18309 7 2 2 56451 61202
0 18310 5 1 1 63865
0 18311 7 1 2 48683 57517
0 18312 5 1 1 18311
0 18313 7 1 2 63838 18312
0 18314 5 1 1 18313
0 18315 7 1 2 49026 18314
0 18316 5 1 1 18315
0 18317 7 1 2 18310 18316
0 18318 5 1 1 18317
0 18319 7 1 2 55064 18318
0 18320 5 1 1 18319
0 18321 7 1 2 18308 18320
0 18322 5 1 1 18321
0 18323 7 1 2 43213 50523
0 18324 7 1 2 18322 18323
0 18325 5 1 1 18324
0 18326 7 1 2 18305 18325
0 18327 5 1 1 18326
0 18328 7 1 2 46399 18327
0 18329 5 1 1 18328
0 18330 7 1 2 52562 62037
0 18331 5 1 1 18330
0 18332 7 2 2 58658 62778
0 18333 7 1 2 45937 61865
0 18334 7 1 2 57145 18333
0 18335 7 1 2 63867 18334
0 18336 5 1 1 18335
0 18337 7 1 2 18331 18336
0 18338 5 1 1 18337
0 18339 7 1 2 42381 18338
0 18340 5 1 1 18339
0 18341 7 2 2 43915 59425
0 18342 7 1 2 61975 60353
0 18343 5 1 1 18342
0 18344 7 2 2 46491 50524
0 18345 7 1 2 62794 63871
0 18346 5 1 1 18345
0 18347 7 1 2 18343 18346
0 18348 5 1 1 18347
0 18349 7 1 2 63869 18348
0 18350 5 1 1 18349
0 18351 7 1 2 18340 18350
0 18352 5 1 1 18351
0 18353 7 1 2 44795 18352
0 18354 5 1 1 18353
0 18355 7 1 2 60287 50525
0 18356 5 1 1 18355
0 18357 7 1 2 60362 18356
0 18358 5 1 1 18357
0 18359 7 2 2 45938 49027
0 18360 7 2 2 61955 63873
0 18361 5 1 1 63875
0 18362 7 1 2 43108 63876
0 18363 7 1 2 18358 18362
0 18364 5 1 1 18363
0 18365 7 1 2 18354 18364
0 18366 5 1 1 18365
0 18367 7 1 2 42824 18366
0 18368 5 1 1 18367
0 18369 7 1 2 61919 63748
0 18370 5 1 1 18369
0 18371 7 1 2 62078 62340
0 18372 5 1 1 18371
0 18373 7 1 2 18370 18372
0 18374 5 1 1 18373
0 18375 7 1 2 42607 18374
0 18376 5 1 1 18375
0 18377 7 2 2 45698 63525
0 18378 5 2 1 63877
0 18379 7 1 2 59469 63878
0 18380 5 1 1 18379
0 18381 7 1 2 18376 18380
0 18382 5 1 1 18381
0 18383 7 2 2 56679 49028
0 18384 7 1 2 18382 63881
0 18385 5 1 1 18384
0 18386 7 1 2 18368 18385
0 18387 5 1 1 18386
0 18388 7 1 2 40029 18387
0 18389 5 1 1 18388
0 18390 7 3 2 55740 61125
0 18391 5 1 1 63883
0 18392 7 1 2 63528 18391
0 18393 5 9 1 18392
0 18394 7 1 2 60288 50494
0 18395 7 1 2 63882 18394
0 18396 7 1 2 63886 18395
0 18397 5 1 1 18396
0 18398 7 1 2 18389 18397
0 18399 7 1 2 18329 18398
0 18400 5 1 1 18399
0 18401 7 1 2 46262 18400
0 18402 5 1 1 18401
0 18403 7 1 2 59085 63872
0 18404 5 1 1 18403
0 18405 7 1 2 17748 18404
0 18406 5 1 1 18405
0 18407 7 1 2 44262 18406
0 18408 5 1 1 18407
0 18409 7 3 2 45699 57260
0 18410 7 1 2 55017 63895
0 18411 5 1 1 18410
0 18412 7 1 2 18408 18411
0 18413 5 1 1 18412
0 18414 7 1 2 40030 18413
0 18415 5 1 1 18414
0 18416 7 1 2 46400 55026
0 18417 5 2 1 18416
0 18418 7 1 2 9981 46648
0 18419 5 1 1 18418
0 18420 7 1 2 60354 18419
0 18421 7 1 2 63898 18420
0 18422 5 1 1 18421
0 18423 7 1 2 18415 18422
0 18424 5 1 1 18423
0 18425 7 1 2 53897 18424
0 18426 5 1 1 18425
0 18427 7 1 2 62729 61660
0 18428 5 1 1 18427
0 18429 7 1 2 18426 18428
0 18430 5 1 1 18429
0 18431 7 1 2 61845 18430
0 18432 5 1 1 18431
0 18433 7 1 2 60636 62233
0 18434 5 1 1 18433
0 18435 7 1 2 63565 18434
0 18436 5 1 1 18435
0 18437 7 1 2 45700 18436
0 18438 5 1 1 18437
0 18439 7 2 2 40031 61355
0 18440 5 1 1 63900
0 18441 7 1 2 51872 63901
0 18442 5 1 1 18441
0 18443 7 1 2 18438 18442
0 18444 5 1 1 18443
0 18445 7 3 2 40393 61877
0 18446 7 1 2 53290 50747
0 18447 7 1 2 63902 18446
0 18448 5 1 1 18447
0 18449 7 1 2 56879 18448
0 18450 5 1 1 18449
0 18451 7 1 2 18444 18450
0 18452 5 1 1 18451
0 18453 7 1 2 42825 18452
0 18454 7 1 2 18432 18453
0 18455 5 1 1 18454
0 18456 7 1 2 63608 63887
0 18457 5 1 1 18456
0 18458 7 8 2 40621 42608
0 18459 5 2 1 63905
0 18460 7 2 2 57159 62106
0 18461 7 1 2 63906 63915
0 18462 5 1 1 18461
0 18463 7 1 2 18457 18462
0 18464 5 1 1 18463
0 18465 7 1 2 55065 18464
0 18466 5 1 1 18465
0 18467 7 1 2 63888 63649
0 18468 5 1 1 18467
0 18469 7 6 2 63907 60463
0 18470 5 1 1 63917
0 18471 7 1 2 61793 63918
0 18472 5 1 1 18471
0 18473 7 1 2 18468 18472
0 18474 7 1 2 18466 18473
0 18475 5 1 1 18474
0 18476 7 1 2 50516 18475
0 18477 5 1 1 18476
0 18478 7 2 2 57261 62734
0 18479 5 1 1 63923
0 18480 7 1 2 54111 55755
0 18481 7 1 2 63924 18480
0 18482 5 1 1 18481
0 18483 7 1 2 18477 18482
0 18484 5 1 1 18483
0 18485 7 1 2 40221 18484
0 18486 5 1 1 18485
0 18487 7 5 2 59000 61866
0 18488 7 1 2 53303 62303
0 18489 7 1 2 63925 18488
0 18490 5 2 1 18489
0 18491 7 1 2 62045 63930
0 18492 5 1 1 18491
0 18493 7 1 2 55741 18492
0 18494 5 1 1 18493
0 18495 7 1 2 53984 61815
0 18496 5 1 1 18495
0 18497 7 1 2 63931 18496
0 18498 5 1 1 18497
0 18499 7 1 2 53210 18498
0 18500 5 1 1 18499
0 18501 7 1 2 18494 18500
0 18502 5 1 1 18501
0 18503 7 1 2 45701 18502
0 18504 5 1 1 18503
0 18505 7 2 2 48500 62855
0 18506 7 1 2 61873 63932
0 18507 5 1 1 18506
0 18508 7 1 2 18504 18507
0 18509 5 1 1 18508
0 18510 7 1 2 48684 18509
0 18511 5 1 1 18510
0 18512 7 2 2 62858 61328
0 18513 5 1 1 63934
0 18514 7 1 2 62046 18513
0 18515 5 1 1 18514
0 18516 7 1 2 53319 63473
0 18517 7 1 2 18515 18516
0 18518 5 1 1 18517
0 18519 7 1 2 46120 18518
0 18520 7 1 2 18511 18519
0 18521 7 1 2 18486 18520
0 18522 5 1 1 18521
0 18523 7 1 2 42978 18522
0 18524 7 1 2 18455 18523
0 18525 5 1 1 18524
0 18526 7 1 2 18402 18525
0 18527 7 1 2 18301 18526
0 18528 5 1 1 18527
0 18529 7 1 2 49204 18528
0 18530 5 1 1 18529
0 18531 7 1 2 941 15418
0 18532 5 2 1 18531
0 18533 7 2 2 51539 63936
0 18534 5 1 1 63938
0 18535 7 1 2 63854 63939
0 18536 5 1 1 18535
0 18537 7 2 2 40032 48501
0 18538 5 1 1 63940
0 18539 7 1 2 63941 59438
0 18540 5 1 1 18539
0 18541 7 1 2 18536 18540
0 18542 5 1 1 18541
0 18543 7 1 2 62719 18542
0 18544 5 1 1 18543
0 18545 7 1 2 48582 62610
0 18546 5 2 1 18545
0 18547 7 1 2 18534 63942
0 18548 5 2 1 18547
0 18549 7 1 2 43382 63943
0 18550 5 1 1 18549
0 18551 7 1 2 62237 18550
0 18552 7 1 2 63944 18551
0 18553 5 1 1 18552
0 18554 7 2 2 45099 52640
0 18555 7 1 2 50089 49113
0 18556 7 1 2 57359 63855
0 18557 7 1 2 18555 18556
0 18558 7 1 2 63946 18557
0 18559 5 1 1 18558
0 18560 7 1 2 18553 18559
0 18561 7 1 2 18544 18560
0 18562 5 1 1 18561
0 18563 7 1 2 50418 18562
0 18564 5 1 1 18563
0 18565 7 4 2 41801 42826
0 18566 7 1 2 53985 61424
0 18567 7 2 2 63635 18566
0 18568 5 1 1 63952
0 18569 7 1 2 63948 63953
0 18570 5 1 1 18569
0 18571 7 3 2 40222 59048
0 18572 5 1 1 63954
0 18573 7 1 2 40033 59952
0 18574 5 1 1 18573
0 18575 7 1 2 18572 18574
0 18576 5 1 1 18575
0 18577 7 1 2 50419 18576
0 18578 7 1 2 63805 18577
0 18579 5 1 1 18578
0 18580 7 1 2 57186 61425
0 18581 7 1 2 63731 18580
0 18582 5 1 1 18581
0 18583 7 1 2 18579 18582
0 18584 5 1 1 18583
0 18585 7 1 2 49029 18584
0 18586 5 1 1 18585
0 18587 7 1 2 18570 18586
0 18588 7 1 2 18564 18587
0 18589 5 1 1 18588
0 18590 7 1 2 41018 18589
0 18591 5 1 1 18590
0 18592 7 1 2 49030 63806
0 18593 5 1 1 18592
0 18594 7 3 2 52858 57125
0 18595 5 1 1 63957
0 18596 7 1 2 63958 50621
0 18597 5 1 1 18596
0 18598 7 2 2 50008 57126
0 18599 5 1 1 63960
0 18600 7 1 2 49114 52841
0 18601 5 1 1 18600
0 18602 7 1 2 18599 18601
0 18603 5 1 1 18602
0 18604 7 1 2 55597 18603
0 18605 5 1 1 18604
0 18606 7 1 2 18597 18605
0 18607 7 1 2 18593 18606
0 18608 5 1 1 18607
0 18609 7 1 2 41802 18608
0 18610 5 1 1 18609
0 18611 7 2 2 55429 54881
0 18612 7 1 2 59361 63962
0 18613 7 1 2 59154 18612
0 18614 5 1 1 18613
0 18615 7 1 2 18610 18614
0 18616 5 1 1 18615
0 18617 7 1 2 63856 18616
0 18618 5 1 1 18617
0 18619 7 1 2 53064 57480
0 18620 7 1 2 57162 62724
0 18621 7 1 2 18619 18620
0 18622 5 1 1 18621
0 18623 7 1 2 18618 18622
0 18624 5 1 1 18623
0 18625 7 1 2 45702 63638
0 18626 7 1 2 18624 18625
0 18627 5 1 1 18626
0 18628 7 1 2 18591 18627
0 18629 5 1 1 18628
0 18630 7 1 2 43214 18629
0 18631 5 1 1 18630
0 18632 7 1 2 59350 63937
0 18633 5 1 1 18632
0 18634 7 2 2 42827 63254
0 18635 5 3 1 63964
0 18636 7 1 2 44796 63965
0 18637 5 1 1 18636
0 18638 7 1 2 18633 18637
0 18639 5 1 1 18638
0 18640 7 1 2 44263 18639
0 18641 5 1 1 18640
0 18642 7 7 2 45100 42979
0 18643 7 1 2 63969 48968
0 18644 7 1 2 63260 18643
0 18645 5 1 1 18644
0 18646 7 1 2 18641 18645
0 18647 5 1 1 18646
0 18648 7 1 2 49031 18647
0 18649 5 1 1 18648
0 18650 7 1 2 62795 63945
0 18651 5 1 1 18650
0 18652 7 1 2 18649 18651
0 18653 5 1 1 18652
0 18654 7 1 2 50420 57177
0 18655 7 1 2 57378 18654
0 18656 7 1 2 18653 18655
0 18657 5 1 1 18656
0 18658 7 1 2 45939 18657
0 18659 7 1 2 18631 18658
0 18660 5 1 1 18659
0 18661 7 1 2 56752 63563
0 18662 5 1 1 18661
0 18663 7 1 2 57946 60330
0 18664 5 1 1 18663
0 18665 7 1 2 12075 18664
0 18666 5 1 1 18665
0 18667 7 1 2 44264 18666
0 18668 5 1 1 18667
0 18669 7 1 2 55018 57262
0 18670 5 1 1 18669
0 18671 7 1 2 18668 18670
0 18672 5 1 1 18671
0 18673 7 1 2 56564 18672
0 18674 5 1 1 18673
0 18675 7 1 2 18662 18674
0 18676 5 1 1 18675
0 18677 7 1 2 18676 63847
0 18678 5 1 1 18677
0 18679 7 1 2 61288 57000
0 18680 5 1 1 18679
0 18681 7 1 2 18678 18680
0 18682 5 1 1 18681
0 18683 7 1 2 40394 18682
0 18684 5 1 1 18683
0 18685 7 2 2 46401 48502
0 18686 7 1 2 61818 61336
0 18687 5 1 1 18686
0 18688 7 1 2 56753 18687
0 18689 5 1 1 18688
0 18690 7 2 2 48066 62924
0 18691 7 1 2 63978 63619
0 18692 5 1 1 18691
0 18693 7 1 2 18689 18692
0 18694 5 1 1 18693
0 18695 7 1 2 63976 18694
0 18696 5 1 1 18695
0 18697 7 2 2 40395 50654
0 18698 5 1 1 63980
0 18699 7 1 2 48563 18698
0 18700 5 2 1 18699
0 18701 7 1 2 41019 59606
0 18702 7 1 2 62275 18701
0 18703 7 1 2 63982 18702
0 18704 5 1 1 18703
0 18705 7 1 2 42980 18704
0 18706 7 1 2 18696 18705
0 18707 7 1 2 18684 18706
0 18708 5 1 1 18707
0 18709 7 1 2 57178 63740
0 18710 5 1 1 18709
0 18711 7 1 2 62925 63857
0 18712 5 1 1 18711
0 18713 7 1 2 18710 18712
0 18714 5 1 1 18713
0 18715 7 1 2 55191 18714
0 18716 5 1 1 18715
0 18717 7 2 2 57412 58618
0 18718 7 1 2 63560 18440
0 18719 5 1 1 18718
0 18720 7 1 2 63984 18719
0 18721 5 1 1 18720
0 18722 7 1 2 18716 18721
0 18723 5 1 1 18722
0 18724 7 1 2 63983 18723
0 18725 5 1 1 18724
0 18726 7 1 2 45101 63926
0 18727 7 1 2 56808 18726
0 18728 5 1 1 18727
0 18729 7 1 2 46263 18728
0 18730 7 1 2 18725 18729
0 18731 5 1 1 18730
0 18732 7 1 2 42828 18731
0 18733 7 1 2 18708 18732
0 18734 5 1 1 18733
0 18735 7 1 2 61313 59936
0 18736 7 1 2 56565 18735
0 18737 5 1 1 18736
0 18738 7 1 2 46264 61830
0 18739 7 1 2 56975 18738
0 18740 7 1 2 62414 18739
0 18741 5 1 1 18740
0 18742 7 1 2 18737 18741
0 18743 5 1 1 18742
0 18744 7 1 2 41020 18743
0 18745 5 1 1 18744
0 18746 7 2 2 41803 59013
0 18747 5 1 1 63986
0 18748 7 1 2 59010 18747
0 18749 5 1 1 18748
0 18750 7 1 2 62410 59282
0 18751 7 1 2 18749 18750
0 18752 5 1 1 18751
0 18753 7 1 2 18745 18752
0 18754 5 1 1 18753
0 18755 7 1 2 43109 18754
0 18756 5 1 1 18755
0 18757 7 1 2 42981 50354
0 18758 7 1 2 56754 18757
0 18759 5 1 1 18758
0 18760 7 1 2 57570 54931
0 18761 7 1 2 59014 18760
0 18762 5 1 1 18761
0 18763 7 1 2 18759 18762
0 18764 5 1 1 18763
0 18765 7 1 2 63813 62411
0 18766 7 1 2 18764 18765
0 18767 5 1 1 18766
0 18768 7 1 2 18756 18767
0 18769 5 1 1 18768
0 18770 7 1 2 51396 18769
0 18771 5 1 1 18770
0 18772 7 1 2 42609 18771
0 18773 7 1 2 18734 18772
0 18774 5 1 1 18773
0 18775 7 1 2 47990 18774
0 18776 7 1 2 18660 18775
0 18777 5 1 1 18776
0 18778 7 2 2 56857 50355
0 18779 5 1 1 63988
0 18780 7 1 2 60762 18779
0 18781 5 1 1 18780
0 18782 7 1 2 63593 18781
0 18783 5 1 1 18782
0 18784 7 1 2 44797 58515
0 18785 5 1 1 18784
0 18786 7 1 2 53083 18785
0 18787 5 1 1 18786
0 18788 7 1 2 40396 18787
0 18789 5 1 1 18788
0 18790 7 1 2 48503 56072
0 18791 5 2 1 18790
0 18792 7 1 2 51406 50517
0 18793 5 1 1 18792
0 18794 7 1 2 63990 18793
0 18795 7 1 2 18789 18794
0 18796 5 1 1 18795
0 18797 7 1 2 40223 18796
0 18798 5 1 1 18797
0 18799 7 1 2 40397 63801
0 18800 5 1 1 18799
0 18801 7 1 2 18798 18800
0 18802 5 2 1 18801
0 18803 7 1 2 54161 63992
0 18804 5 1 1 18803
0 18805 7 1 2 18783 18804
0 18806 5 1 1 18805
0 18807 7 1 2 56349 18806
0 18808 5 1 1 18807
0 18809 7 1 2 51289 51472
0 18810 7 1 2 61022 18809
0 18811 5 1 1 18810
0 18812 7 1 2 18808 18811
0 18813 5 1 1 18812
0 18814 7 1 2 44948 18813
0 18815 5 1 1 18814
0 18816 7 1 2 57091 63989
0 18817 5 1 1 18816
0 18818 7 3 2 40398 53898
0 18819 7 2 2 61894 63994
0 18820 5 1 1 63997
0 18821 7 1 2 61155 54583
0 18822 7 1 2 51683 18821
0 18823 5 1 1 18822
0 18824 7 1 2 18820 18823
0 18825 5 1 1 18824
0 18826 7 1 2 51397 18825
0 18827 5 1 1 18826
0 18828 7 1 2 18817 18827
0 18829 5 1 1 18828
0 18830 7 1 2 55365 18829
0 18831 5 1 1 18830
0 18832 7 1 2 18815 18831
0 18833 5 1 1 18832
0 18834 7 1 2 59470 18833
0 18835 5 1 1 18834
0 18836 7 2 2 51271 55773
0 18837 5 2 1 63999
0 18838 7 1 2 55674 59990
0 18839 5 1 1 18838
0 18840 7 1 2 64001 18839
0 18841 5 1 1 18840
0 18842 7 1 2 60761 18841
0 18843 5 1 1 18842
0 18844 7 3 2 41663 58607
0 18845 7 1 2 40848 41231
0 18846 7 1 2 64003 18845
0 18847 5 1 1 18846
0 18848 7 1 2 64002 18847
0 18849 5 1 1 18848
0 18850 7 1 2 40224 18849
0 18851 5 1 1 18850
0 18852 7 1 2 56338 64004
0 18853 5 1 1 18852
0 18854 7 1 2 18851 18853
0 18855 5 1 1 18854
0 18856 7 1 2 40034 53073
0 18857 7 1 2 18855 18856
0 18858 5 1 1 18857
0 18859 7 1 2 18843 18858
0 18860 5 1 1 18859
0 18861 7 1 2 53986 18860
0 18862 5 1 1 18861
0 18863 7 1 2 50546 52662
0 18864 5 1 1 18863
0 18865 7 1 2 63991 18864
0 18866 5 1 1 18865
0 18867 7 2 2 55675 18866
0 18868 5 1 1 64006
0 18869 7 1 2 53987 64007
0 18870 5 1 1 18869
0 18871 7 2 2 58568 54919
0 18872 7 1 2 41495 64008
0 18873 7 1 2 63903 18872
0 18874 5 1 1 18873
0 18875 7 1 2 18870 18874
0 18876 5 1 1 18875
0 18877 7 1 2 63645 18876
0 18878 5 1 1 18877
0 18879 7 2 2 56885 54458
0 18880 7 1 2 56636 59757
0 18881 7 1 2 64010 18880
0 18882 5 1 1 18881
0 18883 7 1 2 18878 18882
0 18884 7 1 2 18862 18883
0 18885 5 1 1 18884
0 18886 7 1 2 60289 18885
0 18887 5 1 1 18886
0 18888 7 1 2 18835 18887
0 18889 5 1 1 18888
0 18890 7 1 2 42610 18889
0 18891 5 1 1 18890
0 18892 7 11 2 46265 51540
0 18893 7 1 2 61669 63993
0 18894 5 1 1 18893
0 18895 7 1 2 55676 53074
0 18896 5 1 1 18895
0 18897 7 1 2 60763 18896
0 18898 5 1 1 18897
0 18899 7 1 2 40399 18898
0 18900 5 1 1 18899
0 18901 7 1 2 18868 18900
0 18902 5 1 1 18901
0 18903 7 1 2 61744 18902
0 18904 5 1 1 18903
0 18905 7 1 2 18894 18904
0 18906 5 1 1 18905
0 18907 7 1 2 64012 18906
0 18908 5 1 1 18907
0 18909 7 1 2 54572 50529
0 18910 5 1 1 18909
0 18911 7 1 2 61745 18910
0 18912 5 1 1 18911
0 18913 7 1 2 50356 61670
0 18914 5 1 1 18913
0 18915 7 1 2 18912 18914
0 18916 5 1 1 18915
0 18917 7 1 2 56858 18916
0 18918 5 1 1 18917
0 18919 7 1 2 55763 51301
0 18920 7 1 2 61159 18919
0 18921 7 1 2 63518 18920
0 18922 5 1 1 18921
0 18923 7 1 2 18918 18922
0 18924 5 1 1 18923
0 18925 7 1 2 40035 18924
0 18926 5 1 1 18925
0 18927 7 1 2 55764 57282
0 18928 7 1 2 63718 18927
0 18929 5 1 1 18928
0 18930 7 1 2 18926 18929
0 18931 5 1 1 18930
0 18932 7 1 2 55366 18931
0 18933 5 1 1 18932
0 18934 7 1 2 18908 18933
0 18935 5 1 1 18934
0 18936 7 1 2 42611 18935
0 18937 5 1 1 18936
0 18938 7 3 2 40400 55241
0 18939 7 2 2 63664 49115
0 18940 7 1 2 64026 60481
0 18941 5 1 1 18940
0 18942 7 1 2 63448 18941
0 18943 5 1 1 18942
0 18944 7 1 2 63720 18943
0 18945 5 1 1 18944
0 18946 7 1 2 63773 51684
0 18947 7 2 2 52961 51374
0 18948 7 1 2 56566 64028
0 18949 7 1 2 18946 18948
0 18950 5 1 1 18949
0 18951 7 1 2 18945 18950
0 18952 5 1 1 18951
0 18953 7 1 2 64023 18952
0 18954 5 1 1 18953
0 18955 7 1 2 18937 18954
0 18956 5 1 1 18955
0 18957 7 1 2 55066 18956
0 18958 5 1 1 18957
0 18959 7 1 2 64013 63721
0 18960 5 1 1 18959
0 18961 7 1 2 59991 51685
0 18962 7 1 2 64029 18961
0 18963 5 1 1 18962
0 18964 7 1 2 18960 18963
0 18965 5 1 1 18964
0 18966 7 1 2 54162 18965
0 18967 5 1 1 18966
0 18968 7 1 2 18568 18967
0 18969 5 1 1 18968
0 18970 7 1 2 59471 18969
0 18971 5 1 1 18970
0 18972 7 1 2 63724 57179
0 18973 7 2 2 56905 52230
0 18974 7 3 2 46492 63970
0 18975 7 1 2 64032 57928
0 18976 7 1 2 64030 18975
0 18977 7 1 2 18972 18976
0 18978 5 1 1 18977
0 18979 7 1 2 18971 18978
0 18980 5 1 1 18979
0 18981 7 1 2 40401 18980
0 18982 5 1 1 18981
0 18983 7 2 2 40036 53260
0 18984 7 1 2 61175 64035
0 18985 7 1 2 58995 63927
0 18986 7 1 2 18984 18985
0 18987 5 1 1 18986
0 18988 7 1 2 18982 18987
0 18989 5 1 1 18988
0 18990 7 1 2 55242 18989
0 18991 5 1 1 18990
0 18992 7 1 2 18958 18991
0 18993 7 1 2 18891 18992
0 18994 7 1 2 18777 18993
0 18995 7 1 2 18530 18994
0 18996 7 1 2 18087 18995
0 18997 7 1 2 17845 18996
0 18998 5 1 1 18997
0 18999 7 1 2 58546 18998
0 19000 5 1 1 18999
0 19001 7 5 2 40622 49373
0 19002 7 1 2 64037 53501
0 19003 7 1 2 62725 19002
0 19004 7 2 2 61867 63277
0 19005 7 6 2 40402 44307
0 19006 7 4 2 45148 45473
0 19007 7 1 2 61810 64050
0 19008 7 1 2 64044 19007
0 19009 7 1 2 64042 19008
0 19010 7 1 2 19003 19009
0 19011 5 1 1 19010
0 19012 7 1 2 19000 19011
0 19013 5 1 1 19012
0 19014 7 1 2 46738 19013
0 19015 5 1 1 19014
0 19016 7 2 2 63069 61797
0 19017 5 1 1 64054
0 19018 7 4 2 53494 53484
0 19019 7 1 2 46739 64056
0 19020 5 1 1 19019
0 19021 7 1 2 19017 19020
0 19022 5 1 1 19021
0 19023 7 3 2 56680 53458
0 19024 7 3 2 64060 57233
0 19025 7 1 2 19022 64063
0 19026 5 1 1 19025
0 19027 7 1 2 59374 56732
0 19028 5 1 1 19027
0 19029 7 1 2 56927 19028
0 19030 5 1 1 19029
0 19031 7 1 2 42612 19030
0 19032 5 1 1 19031
0 19033 7 2 2 44798 52916
0 19034 5 1 1 64066
0 19035 7 1 2 44949 53075
0 19036 5 1 1 19035
0 19037 7 1 2 19034 19036
0 19038 5 1 1 19037
0 19039 7 1 2 52620 19038
0 19040 5 1 1 19039
0 19041 7 1 2 19032 19040
0 19042 5 1 1 19041
0 19043 7 2 2 40849 19042
0 19044 5 1 1 64068
0 19045 7 5 2 41361 53459
0 19046 7 1 2 64070 52917
0 19047 5 1 1 19046
0 19048 7 1 2 57317 19047
0 19049 5 1 1 19048
0 19050 7 1 2 42982 19049
0 19051 5 1 1 19050
0 19052 7 1 2 57319 19051
0 19053 5 1 1 19052
0 19054 7 1 2 41496 19053
0 19055 5 1 1 19054
0 19056 7 1 2 55212 51642
0 19057 5 1 1 19056
0 19058 7 1 2 19055 19057
0 19059 5 1 1 19058
0 19060 7 1 2 40623 19059
0 19061 5 1 1 19060
0 19062 7 4 2 40037 44950
0 19063 7 1 2 64075 56518
0 19064 5 1 1 19063
0 19065 7 2 2 41664 55818
0 19066 7 1 2 43916 64079
0 19067 5 1 1 19066
0 19068 7 1 2 19064 19067
0 19069 5 1 1 19068
0 19070 7 1 2 46266 19069
0 19071 5 1 1 19070
0 19072 7 1 2 56148 51643
0 19073 5 1 1 19072
0 19074 7 1 2 19071 19073
0 19075 5 1 1 19074
0 19076 7 1 2 44799 19075
0 19077 5 1 1 19076
0 19078 7 1 2 56718 58078
0 19079 7 1 2 62949 19078
0 19080 5 1 1 19079
0 19081 7 1 2 19077 19080
0 19082 7 1 2 19061 19081
0 19083 5 1 1 19082
0 19084 7 1 2 44103 19083
0 19085 5 1 1 19084
0 19086 7 1 2 19044 19085
0 19087 5 1 1 19086
0 19088 7 1 2 46740 19087
0 19089 5 1 1 19088
0 19090 7 1 2 40038 64069
0 19091 5 1 1 19090
0 19092 7 2 2 42829 63665
0 19093 5 2 1 64081
0 19094 7 1 2 46799 52741
0 19095 5 1 1 19094
0 19096 7 1 2 64083 19095
0 19097 5 1 1 19096
0 19098 7 1 2 49595 19097
0 19099 5 1 1 19098
0 19100 7 1 2 51949 50655
0 19101 5 1 1 19100
0 19102 7 1 2 18538 19101
0 19103 5 1 1 19102
0 19104 7 1 2 48969 19103
0 19105 5 1 1 19104
0 19106 7 1 2 19099 19105
0 19107 5 1 1 19106
0 19108 7 1 2 46267 19107
0 19109 5 1 1 19108
0 19110 7 2 2 48114 63666
0 19111 5 1 1 64085
0 19112 7 1 2 56733 64086
0 19113 5 1 1 19112
0 19114 7 1 2 19109 19113
0 19115 5 1 1 19114
0 19116 7 1 2 42613 19115
0 19117 5 1 1 19116
0 19118 7 3 2 44800 46800
0 19119 7 2 2 48254 64087
0 19120 5 1 1 64090
0 19121 7 2 2 48504 52918
0 19122 5 2 1 64092
0 19123 7 1 2 46121 50735
0 19124 5 1 1 19123
0 19125 7 1 2 64094 19124
0 19126 5 1 1 19125
0 19127 7 1 2 40039 42983
0 19128 7 1 2 19126 19127
0 19129 5 1 1 19128
0 19130 7 1 2 19120 19129
0 19131 5 1 1 19130
0 19132 7 1 2 56149 19131
0 19133 5 1 1 19132
0 19134 7 1 2 19117 19133
0 19135 5 1 1 19134
0 19136 7 1 2 44104 19135
0 19137 5 1 1 19136
0 19138 7 1 2 19091 19137
0 19139 7 1 2 19089 19138
0 19140 5 1 1 19139
0 19141 7 1 2 40403 19140
0 19142 5 1 1 19141
0 19143 7 1 2 57341 61121
0 19144 5 1 1 19143
0 19145 7 1 2 48851 49248
0 19146 5 1 1 19145
0 19147 7 1 2 57922 57674
0 19148 5 1 1 19147
0 19149 7 1 2 19146 19148
0 19150 5 1 1 19149
0 19151 7 1 2 46268 19150
0 19152 5 1 1 19151
0 19153 7 1 2 48852 48138
0 19154 5 1 1 19153
0 19155 7 1 2 19152 19154
0 19156 5 1 1 19155
0 19157 7 1 2 49596 19156
0 19158 5 1 1 19157
0 19159 7 1 2 19144 19158
0 19160 5 1 1 19159
0 19161 7 1 2 40040 19160
0 19162 5 1 1 19161
0 19163 7 1 2 48853 63097
0 19164 5 1 1 19163
0 19165 7 1 2 943 19164
0 19166 5 1 1 19165
0 19167 7 1 2 49205 19166
0 19168 5 1 1 19167
0 19169 7 3 2 48854 56985
0 19170 7 1 2 55367 64096
0 19171 5 1 1 19170
0 19172 7 1 2 48214 51664
0 19173 7 1 2 52142 19172
0 19174 5 1 1 19173
0 19175 7 1 2 19171 19174
0 19176 7 1 2 19168 19175
0 19177 5 1 1 19176
0 19178 7 1 2 46741 19177
0 19179 5 1 1 19178
0 19180 7 1 2 48215 51959
0 19181 7 1 2 57546 19180
0 19182 5 1 1 19181
0 19183 7 1 2 19179 19182
0 19184 7 1 2 19162 19183
0 19185 5 1 1 19184
0 19186 7 1 2 42614 19185
0 19187 5 1 1 19186
0 19188 7 1 2 19142 19187
0 19189 5 1 1 19188
0 19190 7 1 2 46402 19189
0 19191 5 1 1 19190
0 19192 7 1 2 19026 19191
0 19193 5 1 1 19192
0 19194 7 1 2 40225 19193
0 19195 5 1 1 19194
0 19196 7 1 2 48505 55297
0 19197 5 1 1 19196
0 19198 7 1 2 57877 19197
0 19199 5 1 1 19198
0 19200 7 1 2 60554 19199
0 19201 5 1 1 19200
0 19202 7 5 2 41115 57571
0 19203 7 5 2 64099 52509
0 19204 7 1 2 64104 57882
0 19205 5 1 1 19204
0 19206 7 1 2 19201 19205
0 19207 5 1 1 19206
0 19208 7 1 2 42615 19207
0 19209 5 1 1 19208
0 19210 7 2 2 45940 57572
0 19211 7 1 2 46801 51999
0 19212 7 1 2 64109 19211
0 19213 7 1 2 57898 19212
0 19214 5 1 1 19213
0 19215 7 1 2 19209 19214
0 19216 5 1 1 19215
0 19217 7 1 2 42984 19216
0 19218 5 1 1 19217
0 19219 7 1 2 58272 63170
0 19220 5 2 1 19219
0 19221 7 1 2 57552 64111
0 19222 5 1 1 19221
0 19223 7 1 2 19218 19222
0 19224 5 1 1 19223
0 19225 7 1 2 46403 19224
0 19226 5 1 1 19225
0 19227 7 3 2 45303 57821
0 19228 5 2 1 64113
0 19229 7 5 2 41497 52000
0 19230 7 1 2 46122 63319
0 19231 7 1 2 56897 19230
0 19232 7 1 2 64118 19231
0 19233 7 1 2 64114 19232
0 19234 5 1 1 19233
0 19235 7 1 2 19226 19234
0 19236 7 1 2 19195 19235
0 19237 5 1 1 19236
0 19238 7 1 2 53899 19237
0 19239 5 1 1 19238
0 19240 7 5 2 44212 51456
0 19241 7 1 2 49306 57953
0 19242 7 1 2 64123 19241
0 19243 5 1 1 19242
0 19244 7 2 2 40850 53495
0 19245 7 2 2 56886 53065
0 19246 7 2 2 45703 46742
0 19247 7 1 2 64130 64132
0 19248 7 1 2 64128 19247
0 19249 5 1 1 19248
0 19250 7 1 2 19243 19249
0 19251 5 1 1 19250
0 19252 7 7 2 56785 63236
0 19253 7 1 2 40226 50641
0 19254 7 1 2 64134 19253
0 19255 7 1 2 19251 19254
0 19256 5 1 1 19255
0 19257 7 1 2 19239 19256
0 19258 5 1 1 19257
0 19259 7 1 2 46565 19258
0 19260 5 1 1 19259
0 19261 7 1 2 52919 61910
0 19262 5 2 1 19261
0 19263 7 2 2 55243 50400
0 19264 5 1 1 64143
0 19265 7 2 2 61772 64144
0 19266 5 1 1 64145
0 19267 7 1 2 40851 64146
0 19268 5 1 1 19267
0 19269 7 1 2 64141 19268
0 19270 5 1 1 19269
0 19271 7 1 2 45704 19270
0 19272 5 1 1 19271
0 19273 7 2 2 44951 51457
0 19274 7 6 2 42616 49512
0 19275 7 1 2 64149 50944
0 19276 7 1 2 64147 19275
0 19277 5 1 1 19276
0 19278 7 1 2 19272 19277
0 19279 5 1 1 19278
0 19280 7 1 2 42985 19279
0 19281 5 1 1 19280
0 19282 7 1 2 44105 63889
0 19283 5 1 1 19282
0 19284 7 1 2 54465 19283
0 19285 5 1 1 19284
0 19286 7 1 2 45705 19285
0 19287 5 1 1 19286
0 19288 7 3 2 49513 56030
0 19289 5 2 1 64155
0 19290 7 1 2 44106 64156
0 19291 5 1 1 19290
0 19292 7 1 2 19287 19291
0 19293 5 1 1 19292
0 19294 7 1 2 48270 19293
0 19295 5 1 1 19294
0 19296 7 1 2 52453 56932
0 19297 5 2 1 19296
0 19298 7 1 2 19295 64160
0 19299 7 1 2 19281 19298
0 19300 5 1 1 19299
0 19301 7 1 2 40041 19300
0 19302 5 1 1 19301
0 19303 7 1 2 63483 19302
0 19304 5 1 1 19303
0 19305 7 1 2 46743 19304
0 19306 5 1 1 19305
0 19307 7 1 2 48401 57852
0 19308 5 1 1 19307
0 19309 7 1 2 5274 19308
0 19310 5 1 1 19309
0 19311 7 1 2 40852 19310
0 19312 5 1 1 19311
0 19313 7 5 2 49597 56350
0 19314 7 3 2 45304 52920
0 19315 5 1 1 64167
0 19316 7 1 2 40042 64168
0 19317 5 1 1 19316
0 19318 7 1 2 60701 19317
0 19319 5 2 1 19318
0 19320 7 1 2 64162 64170
0 19321 5 1 1 19320
0 19322 7 1 2 19312 19321
0 19323 5 1 1 19322
0 19324 7 2 2 49514 19323
0 19325 5 1 1 64172
0 19326 7 1 2 42617 64173
0 19327 5 1 1 19326
0 19328 7 1 2 49515 64163
0 19329 5 1 1 19328
0 19330 7 1 2 61961 63125
0 19331 5 1 1 19330
0 19332 7 1 2 19329 19331
0 19333 5 1 1 19332
0 19334 7 1 2 42618 19333
0 19335 5 1 1 19334
0 19336 7 5 2 45706 52608
0 19337 7 1 2 64174 48685
0 19338 7 1 2 57890 19337
0 19339 5 1 1 19338
0 19340 7 1 2 19335 19339
0 19341 5 1 1 19340
0 19342 7 1 2 52921 19341
0 19343 5 1 1 19342
0 19344 7 1 2 48876 53532
0 19345 5 1 1 19344
0 19346 7 1 2 45707 62559
0 19347 5 1 1 19346
0 19348 7 1 2 19345 19347
0 19349 5 1 1 19348
0 19350 7 1 2 42619 19349
0 19351 5 1 1 19350
0 19352 7 1 2 53211 55782
0 19353 5 1 1 19352
0 19354 7 1 2 19351 19353
0 19355 5 1 1 19354
0 19356 7 1 2 48271 19355
0 19357 5 1 1 19356
0 19358 7 3 2 41362 53831
0 19359 5 2 1 64179
0 19360 7 1 2 40404 55269
0 19361 5 1 1 19360
0 19362 7 1 2 64182 19361
0 19363 5 1 1 19362
0 19364 7 1 2 57443 19363
0 19365 5 1 1 19364
0 19366 7 1 2 49598 62399
0 19367 7 1 2 59229 19366
0 19368 5 1 1 19367
0 19369 7 1 2 19365 19368
0 19370 5 1 1 19369
0 19371 7 1 2 44952 19370
0 19372 5 1 1 19371
0 19373 7 1 2 64161 19372
0 19374 7 1 2 19357 19373
0 19375 7 1 2 19343 19374
0 19376 5 1 1 19375
0 19377 7 1 2 52093 19376
0 19378 5 1 1 19377
0 19379 7 1 2 19327 19378
0 19380 7 1 2 19306 19379
0 19381 5 1 1 19380
0 19382 7 2 2 45056 59630
0 19383 7 1 2 64184 59637
0 19384 7 1 2 19381 19383
0 19385 5 1 1 19384
0 19386 7 1 2 19260 19385
0 19387 5 1 1 19386
0 19388 7 1 2 46493 19387
0 19389 5 1 1 19388
0 19390 7 1 2 44662 50384
0 19391 5 2 1 19390
0 19392 7 1 2 55774 55756
0 19393 7 1 2 64186 19392
0 19394 5 1 1 19393
0 19395 7 1 2 54466 19394
0 19396 5 1 1 19395
0 19397 7 1 2 40227 19396
0 19398 5 1 1 19397
0 19399 7 3 2 42620 47466
0 19400 7 1 2 64188 54459
0 19401 5 1 1 19400
0 19402 7 1 2 19398 19401
0 19403 5 1 1 19402
0 19404 7 1 2 45708 19403
0 19405 5 1 1 19404
0 19406 7 1 2 1815 3097
0 19407 5 1 1 19406
0 19408 7 2 2 54320 53261
0 19409 7 1 2 19407 64191
0 19410 5 1 1 19409
0 19411 7 1 2 19405 19410
0 19412 5 1 1 19411
0 19413 7 1 2 48272 19412
0 19414 5 1 1 19413
0 19415 7 1 2 56734 63657
0 19416 5 1 1 19415
0 19417 7 2 2 50329 50736
0 19418 7 1 2 64193 62213
0 19419 5 1 1 19418
0 19420 7 1 2 19416 19419
0 19421 5 1 1 19420
0 19422 7 1 2 54502 19421
0 19423 5 1 1 19422
0 19424 7 1 2 50330 53375
0 19425 7 1 2 62214 19424
0 19426 5 1 1 19425
0 19427 7 1 2 54652 53244
0 19428 7 1 2 57891 19427
0 19429 7 1 2 64187 19428
0 19430 5 1 1 19429
0 19431 7 1 2 19426 19430
0 19432 5 1 1 19431
0 19433 7 1 2 45941 19432
0 19434 5 1 1 19433
0 19435 7 1 2 19423 19434
0 19436 5 1 1 19435
0 19437 7 1 2 46123 19436
0 19438 5 1 1 19437
0 19439 7 1 2 51574 57939
0 19440 7 3 2 63387 19439
0 19441 7 1 2 48686 64195
0 19442 5 1 1 19441
0 19443 7 1 2 48067 49666
0 19444 5 1 1 19443
0 19445 7 1 2 19442 19444
0 19446 5 2 1 19445
0 19447 7 2 2 47276 62293
0 19448 7 1 2 55614 64200
0 19449 7 1 2 64198 19448
0 19450 5 1 1 19449
0 19451 7 1 2 19438 19450
0 19452 5 1 1 19451
0 19453 7 1 2 42986 19452
0 19454 5 1 1 19453
0 19455 7 2 2 49771 52922
0 19456 7 1 2 52454 64164
0 19457 7 1 2 64202 19456
0 19458 5 1 1 19457
0 19459 7 1 2 19454 19458
0 19460 7 1 2 19414 19459
0 19461 5 1 1 19460
0 19462 7 1 2 53900 19461
0 19463 5 1 1 19462
0 19464 7 2 2 60600 57613
0 19465 7 1 2 56950 63278
0 19466 7 1 2 64204 19465
0 19467 5 1 1 19466
0 19468 7 1 2 19463 19467
0 19469 5 1 1 19468
0 19470 7 1 2 46404 19469
0 19471 5 1 1 19470
0 19472 7 3 2 48115 48439
0 19473 5 1 1 64206
0 19474 7 1 2 15221 19473
0 19475 5 6 1 19474
0 19476 7 1 2 64209 56741
0 19477 5 1 1 19476
0 19478 7 2 2 48116 51730
0 19479 7 1 2 64119 53262
0 19480 7 1 2 64215 19479
0 19481 5 1 1 19480
0 19482 7 1 2 19477 19481
0 19483 5 1 1 19482
0 19484 7 1 2 40043 19483
0 19485 5 1 1 19484
0 19486 7 2 2 54503 47229
0 19487 5 1 1 64217
0 19488 7 2 2 50742 54951
0 19489 7 1 2 64218 64219
0 19490 5 1 1 19489
0 19491 7 1 2 19485 19490
0 19492 5 1 1 19491
0 19493 7 1 2 46405 19492
0 19494 5 1 1 19493
0 19495 7 1 2 62615 64064
0 19496 5 1 1 19495
0 19497 7 1 2 19494 19496
0 19498 5 1 1 19497
0 19499 7 1 2 53901 19498
0 19500 5 1 1 19499
0 19501 7 2 2 64135 50801
0 19502 7 5 2 40044 41363
0 19503 7 1 2 64223 49129
0 19504 7 1 2 64221 19503
0 19505 5 1 1 19504
0 19506 7 1 2 19500 19505
0 19507 5 1 1 19506
0 19508 7 1 2 52254 19507
0 19509 5 1 1 19508
0 19510 7 2 2 48506 59251
0 19511 5 1 1 64228
0 19512 7 1 2 53642 64229
0 19513 5 1 1 19512
0 19514 7 1 2 54321 56660
0 19515 5 1 1 19514
0 19516 7 1 2 57495 19515
0 19517 5 1 1 19516
0 19518 7 1 2 41665 61080
0 19519 7 1 2 19517 19518
0 19520 5 1 1 19519
0 19521 7 1 2 19513 19520
0 19522 5 1 1 19521
0 19523 7 1 2 46744 19522
0 19524 5 1 1 19523
0 19525 7 1 2 52973 64093
0 19526 5 1 1 19525
0 19527 7 2 2 46802 60531
0 19528 5 1 1 64230
0 19529 7 1 2 49667 54653
0 19530 7 1 2 64231 19529
0 19531 5 1 1 19530
0 19532 7 1 2 19526 19531
0 19533 5 1 1 19532
0 19534 7 1 2 63653 19533
0 19535 5 1 1 19534
0 19536 7 1 2 56232 63336
0 19537 7 1 2 57794 19536
0 19538 5 1 1 19537
0 19539 7 1 2 19535 19538
0 19540 7 1 2 19524 19539
0 19541 5 1 1 19540
0 19542 7 1 2 40853 19541
0 19543 5 1 1 19542
0 19544 7 2 2 48507 48273
0 19545 5 1 1 64232
0 19546 7 1 2 42621 58684
0 19547 7 1 2 49772 19546
0 19548 7 1 2 64233 19547
0 19549 5 1 1 19548
0 19550 7 1 2 19543 19549
0 19551 5 1 1 19550
0 19552 7 1 2 53902 19551
0 19553 5 1 1 19552
0 19554 7 2 2 45305 62097
0 19555 7 1 2 64136 61081
0 19556 7 1 2 57797 19555
0 19557 7 1 2 64234 19556
0 19558 5 1 1 19557
0 19559 7 1 2 19553 19558
0 19560 5 1 1 19559
0 19561 7 1 2 48855 19560
0 19562 5 1 1 19561
0 19563 7 1 2 55677 55275
0 19564 5 1 1 19563
0 19565 7 1 2 40405 58426
0 19566 5 1 1 19565
0 19567 7 1 2 19564 19566
0 19568 5 1 1 19567
0 19569 7 1 2 42987 19568
0 19570 5 1 1 19569
0 19571 7 1 2 42830 64000
0 19572 5 1 1 19571
0 19573 7 1 2 19570 19572
0 19574 5 1 1 19573
0 19575 7 1 2 56738 19574
0 19576 5 1 1 19575
0 19577 7 3 2 48687 53460
0 19578 7 1 2 5270 57757
0 19579 5 1 1 19578
0 19580 7 1 2 44107 19579
0 19581 5 1 1 19580
0 19582 7 1 2 53513 57754
0 19583 5 1 1 19582
0 19584 7 1 2 19581 19583
0 19585 5 2 1 19584
0 19586 7 1 2 64236 64239
0 19587 5 1 1 19586
0 19588 7 1 2 19576 19587
0 19589 5 1 1 19588
0 19590 7 1 2 46406 19589
0 19591 5 1 1 19590
0 19592 7 1 2 62279 64129
0 19593 7 1 2 64065 19592
0 19594 5 1 1 19593
0 19595 7 1 2 19591 19594
0 19596 5 1 1 19595
0 19597 7 1 2 53903 19596
0 19598 5 1 1 19597
0 19599 7 1 2 64124 61798
0 19600 7 1 2 64222 19599
0 19601 5 1 1 19600
0 19602 7 1 2 19598 19601
0 19603 5 1 1 19602
0 19604 7 1 2 46745 19603
0 19605 5 1 1 19604
0 19606 7 1 2 19562 19605
0 19607 7 1 2 19509 19606
0 19608 7 1 2 19471 19607
0 19609 5 1 1 19608
0 19610 7 1 2 59335 19609
0 19611 5 1 1 19610
0 19612 7 1 2 19389 19611
0 19613 5 1 1 19612
0 19614 7 1 2 55067 19613
0 19615 5 1 1 19614
0 19616 7 1 2 49599 63198
0 19617 5 1 1 19616
0 19618 7 1 2 54609 46687
0 19619 7 1 2 57940 19618
0 19620 5 1 1 19619
0 19621 7 1 2 19617 19620
0 19622 5 1 1 19621
0 19623 7 1 2 41964 19622
0 19624 5 1 1 19623
0 19625 7 3 2 43110 48216
0 19626 7 1 2 64241 64196
0 19627 5 1 1 19626
0 19628 7 1 2 19624 19627
0 19629 5 1 1 19628
0 19630 7 1 2 51920 19629
0 19631 5 1 1 19630
0 19632 7 1 2 57929 59130
0 19633 5 1 1 19632
0 19634 7 1 2 19631 19633
0 19635 5 1 1 19634
0 19636 7 1 2 41116 19635
0 19637 5 1 1 19636
0 19638 7 3 2 45306 46269
0 19639 7 1 2 55615 63388
0 19640 5 1 1 19639
0 19641 7 1 2 55742 52923
0 19642 5 1 1 19641
0 19643 7 1 2 19640 19642
0 19644 5 1 1 19643
0 19645 7 1 2 64244 19644
0 19646 5 1 1 19645
0 19647 7 1 2 57592 60809
0 19648 5 1 1 19647
0 19649 7 1 2 19646 19648
0 19650 5 1 1 19649
0 19651 7 1 2 40854 19650
0 19652 5 1 1 19651
0 19653 7 2 2 50108 57234
0 19654 7 1 2 40624 64247
0 19655 7 1 2 63273 19654
0 19656 5 1 1 19655
0 19657 7 1 2 19652 19656
0 19658 5 1 1 19657
0 19659 7 1 2 43111 19658
0 19660 5 1 1 19659
0 19661 7 1 2 19637 19660
0 19662 5 1 1 19661
0 19663 7 1 2 41364 19662
0 19664 5 1 1 19663
0 19665 7 2 2 57942 56788
0 19666 5 1 1 64249
0 19667 7 1 2 40625 64250
0 19668 5 1 1 19667
0 19669 7 1 2 40855 57356
0 19670 5 1 1 19669
0 19671 7 1 2 19668 19670
0 19672 5 2 1 19671
0 19673 7 1 2 43112 64251
0 19674 5 1 1 19673
0 19675 7 1 2 49668 51541
0 19676 7 1 2 57469 19675
0 19677 5 1 1 19676
0 19678 7 1 2 19674 19677
0 19679 5 1 1 19678
0 19680 7 1 2 64133 19679
0 19681 5 1 1 19680
0 19682 7 1 2 19664 19681
0 19683 5 1 1 19682
0 19684 7 1 2 40406 19683
0 19685 5 1 1 19684
0 19686 7 3 2 40626 57593
0 19687 5 1 1 64253
0 19688 7 1 2 64254 64120
0 19689 5 3 1 19688
0 19690 7 1 2 51941 53392
0 19691 5 9 1 19690
0 19692 7 2 2 49669 64259
0 19693 5 1 1 64268
0 19694 7 1 2 63289 56730
0 19695 7 1 2 19693 19694
0 19696 5 1 1 19695
0 19697 7 1 2 48217 19696
0 19698 5 1 1 19697
0 19699 7 1 2 64256 19698
0 19700 5 1 1 19699
0 19701 7 1 2 48068 19700
0 19702 5 1 1 19701
0 19703 7 2 2 56719 50145
0 19704 5 2 1 64270
0 19705 7 3 2 57943 64271
0 19706 7 1 2 53263 64274
0 19707 5 1 1 19706
0 19708 7 1 2 19702 19707
0 19709 5 1 1 19708
0 19710 7 1 2 46746 19709
0 19711 5 1 1 19710
0 19712 7 3 2 40856 41117
0 19713 7 1 2 64277 63478
0 19714 7 1 2 64194 19713
0 19715 5 1 1 19714
0 19716 7 1 2 19711 19715
0 19717 5 1 1 19716
0 19718 7 1 2 43113 19717
0 19719 5 1 1 19718
0 19720 7 1 2 49670 60794
0 19721 5 1 1 19720
0 19722 7 1 2 63290 19721
0 19723 5 1 1 19722
0 19724 7 1 2 46747 58569
0 19725 7 1 2 57503 19724
0 19726 7 1 2 19723 19725
0 19727 5 1 1 19726
0 19728 7 1 2 19719 19727
0 19729 7 1 2 19685 19728
0 19730 5 1 1 19729
0 19731 7 1 2 40045 19730
0 19732 5 1 1 19731
0 19733 7 1 2 53600 48342
0 19734 7 1 2 57808 19733
0 19735 5 1 1 19734
0 19736 7 2 2 64278 48360
0 19737 7 1 2 56073 58588
0 19738 7 1 2 64280 19737
0 19739 5 1 1 19738
0 19740 7 1 2 19735 19739
0 19741 5 1 1 19740
0 19742 7 1 2 44801 19741
0 19743 5 1 1 19742
0 19744 7 3 2 45709 46803
0 19745 5 1 1 64282
0 19746 7 1 2 48069 57352
0 19747 5 1 1 19746
0 19748 7 1 2 19666 19747
0 19749 5 1 1 19748
0 19750 7 1 2 43114 19749
0 19751 5 1 1 19750
0 19752 7 1 2 48583 60044
0 19753 5 1 1 19752
0 19754 7 1 2 19751 19753
0 19755 5 1 1 19754
0 19756 7 1 2 40627 19755
0 19757 5 1 1 19756
0 19758 7 2 2 41498 55819
0 19759 7 1 2 57827 6049
0 19760 5 5 1 19759
0 19761 7 1 2 64285 64287
0 19762 5 1 1 19761
0 19763 7 1 2 19757 19762
0 19764 5 1 1 19763
0 19765 7 1 2 64283 19764
0 19766 5 1 1 19765
0 19767 7 1 2 19743 19766
0 19768 5 1 1 19767
0 19769 7 1 2 49516 19768
0 19770 5 1 1 19769
0 19771 7 1 2 56341 63263
0 19772 5 1 1 19771
0 19773 7 1 2 53609 56957
0 19774 5 1 1 19773
0 19775 7 1 2 19772 19774
0 19776 5 1 1 19775
0 19777 7 1 2 46804 19776
0 19778 5 1 1 19777
0 19779 7 3 2 53643 50765
0 19780 7 1 2 56482 64292
0 19781 5 1 1 19780
0 19782 7 1 2 19778 19781
0 19783 5 1 1 19782
0 19784 7 1 2 44953 19783
0 19785 5 1 1 19784
0 19786 7 3 2 55590 61126
0 19787 5 1 1 64295
0 19788 7 1 2 54610 64281
0 19789 7 1 2 64296 19788
0 19790 5 1 1 19789
0 19791 7 1 2 19785 19790
0 19792 5 1 1 19791
0 19793 7 1 2 42622 19792
0 19794 5 1 1 19793
0 19795 7 1 2 64248 61426
0 19796 5 1 1 19795
0 19797 7 2 2 48218 47972
0 19798 5 1 1 64298
0 19799 7 1 2 19798 63355
0 19800 5 1 1 19799
0 19801 7 1 2 48688 63389
0 19802 7 1 2 19800 19801
0 19803 5 1 1 19802
0 19804 7 1 2 19796 19803
0 19805 5 1 1 19804
0 19806 7 1 2 40857 19805
0 19807 5 1 1 19806
0 19808 7 1 2 64299 62638
0 19809 5 1 1 19808
0 19810 7 1 2 19807 19809
0 19811 5 1 1 19810
0 19812 7 1 2 41118 57682
0 19813 7 1 2 19811 19812
0 19814 5 1 1 19813
0 19815 7 1 2 19794 19814
0 19816 7 1 2 19770 19815
0 19817 7 1 2 19732 19816
0 19818 5 1 1 19817
0 19819 7 1 2 41804 19818
0 19820 5 1 1 19819
0 19821 7 1 2 50820 19787
0 19822 5 3 1 19821
0 19823 7 1 2 42623 64300
0 19824 5 1 1 19823
0 19825 7 1 2 48689 61177
0 19826 5 1 1 19825
0 19827 7 1 2 19824 19826
0 19828 5 2 1 19827
0 19829 7 1 2 45710 64303
0 19830 5 2 1 19829
0 19831 7 7 2 40046 42831
0 19832 7 2 2 46805 64307
0 19833 7 1 2 63884 64314
0 19834 5 1 1 19833
0 19835 7 1 2 64305 19834
0 19836 5 1 1 19835
0 19837 7 1 2 46270 19836
0 19838 5 1 1 19837
0 19839 7 2 2 57594 61956
0 19840 5 1 1 64316
0 19841 7 1 2 59890 64317
0 19842 5 1 1 19841
0 19843 7 1 2 19838 19842
0 19844 5 1 1 19843
0 19845 7 1 2 41666 19844
0 19846 5 1 1 19845
0 19847 7 3 2 42624 57573
0 19848 7 1 2 50031 54241
0 19849 7 1 2 64318 19848
0 19850 7 1 2 63331 19849
0 19851 5 1 1 19850
0 19852 7 1 2 19846 19851
0 19853 5 1 1 19852
0 19854 7 1 2 40858 19853
0 19855 5 1 1 19854
0 19856 7 2 2 55775 64275
0 19857 7 1 2 40628 64321
0 19858 5 3 1 19857
0 19859 7 2 2 53330 58494
0 19860 5 1 1 64326
0 19861 7 1 2 46271 64327
0 19862 5 2 1 19861
0 19863 7 2 2 45711 64252
0 19864 7 1 2 58250 64330
0 19865 5 1 1 19864
0 19866 7 1 2 64328 19865
0 19867 5 1 1 19866
0 19868 7 1 2 49517 19867
0 19869 5 1 1 19868
0 19870 7 1 2 64323 19869
0 19871 7 1 2 19855 19870
0 19872 5 1 1 19871
0 19873 7 1 2 59049 19872
0 19874 5 1 1 19873
0 19875 7 1 2 19820 19874
0 19876 5 1 1 19875
0 19877 7 1 2 40228 19876
0 19878 5 1 1 19877
0 19879 7 1 2 57595 50797
0 19880 7 1 2 64057 19879
0 19881 5 2 1 19880
0 19882 7 4 2 44108 50146
0 19883 7 1 2 57973 64334
0 19884 5 1 1 19883
0 19885 7 1 2 19487 19884
0 19886 5 1 1 19885
0 19887 7 1 2 40407 19886
0 19888 5 1 1 19887
0 19889 7 1 2 48856 54504
0 19890 7 1 2 60709 19889
0 19891 5 1 1 19890
0 19892 7 1 2 19888 19891
0 19893 5 1 1 19892
0 19894 7 1 2 48508 19893
0 19895 5 1 1 19894
0 19896 7 2 2 42832 48070
0 19897 5 1 1 64338
0 19898 7 1 2 41365 51921
0 19899 5 3 1 19898
0 19900 7 1 2 43716 64340
0 19901 5 1 1 19900
0 19902 7 1 2 64269 19901
0 19903 5 1 1 19902
0 19904 7 1 2 63879 19903
0 19905 5 1 1 19904
0 19906 7 1 2 64339 19905
0 19907 5 1 1 19906
0 19908 7 1 2 19895 19907
0 19909 5 1 1 19908
0 19910 7 1 2 46272 19909
0 19911 5 1 1 19910
0 19912 7 1 2 64332 19911
0 19913 5 1 1 19912
0 19914 7 1 2 59953 19913
0 19915 5 1 1 19914
0 19916 7 1 2 56180 59362
0 19917 7 1 2 55283 19916
0 19918 5 1 1 19917
0 19919 7 3 2 62027 59393
0 19920 5 1 1 64343
0 19921 7 1 2 45712 64344
0 19922 5 1 1 19921
0 19923 7 1 2 49445 19922
0 19924 5 1 1 19923
0 19925 7 1 2 63255 19920
0 19926 5 2 1 19925
0 19927 7 1 2 42833 64346
0 19928 7 1 2 19924 19927
0 19929 5 1 1 19928
0 19930 7 1 2 19918 19929
0 19931 5 1 1 19930
0 19932 7 1 2 42625 19931
0 19933 5 1 1 19932
0 19934 7 6 2 40408 45102
0 19935 7 2 2 64348 56150
0 19936 7 1 2 45307 64354
0 19937 7 1 2 63803 19936
0 19938 5 1 1 19937
0 19939 7 1 2 19933 19938
0 19940 5 1 1 19939
0 19941 7 1 2 41499 19940
0 19942 5 1 1 19941
0 19943 7 4 2 42834 52001
0 19944 7 1 2 55314 64356
0 19945 7 1 2 64347 19944
0 19946 5 1 1 19945
0 19947 7 1 2 19942 19946
0 19948 5 1 1 19947
0 19949 7 1 2 40629 19948
0 19950 5 1 1 19949
0 19951 7 1 2 49143 59937
0 19952 5 1 1 19951
0 19953 7 1 2 45103 59394
0 19954 7 1 2 64301 19953
0 19955 5 1 1 19954
0 19956 7 1 2 19952 19955
0 19957 5 1 1 19956
0 19958 7 1 2 45713 19957
0 19959 5 1 1 19958
0 19960 7 1 2 40859 56859
0 19961 7 1 2 59280 19960
0 19962 5 1 1 19961
0 19963 7 1 2 44802 58772
0 19964 7 1 2 63186 19963
0 19965 7 1 2 57704 19964
0 19966 5 1 1 19965
0 19967 7 1 2 19962 19966
0 19968 5 1 1 19967
0 19969 7 1 2 49518 19968
0 19970 5 1 1 19969
0 19971 7 1 2 19959 19970
0 19972 5 1 1 19971
0 19973 7 1 2 42626 19972
0 19974 5 1 1 19973
0 19975 7 1 2 64355 63807
0 19976 5 1 1 19975
0 19977 7 1 2 19974 19976
0 19978 5 1 1 19977
0 19979 7 1 2 47467 19978
0 19980 5 1 1 19979
0 19981 7 4 2 56074 48690
0 19982 7 1 2 54357 64345
0 19983 5 1 1 19982
0 19984 7 1 2 41805 58722
0 19985 7 1 2 56789 19984
0 19986 5 1 1 19985
0 19987 7 1 2 19983 19986
0 19988 5 1 1 19987
0 19989 7 1 2 64360 19988
0 19990 5 1 1 19989
0 19991 7 1 2 19980 19990
0 19992 7 1 2 19950 19991
0 19993 5 1 1 19992
0 19994 7 1 2 46407 19993
0 19995 5 1 1 19994
0 19996 7 1 2 19915 19995
0 19997 7 1 2 19878 19996
0 19998 5 1 1 19997
0 19999 7 1 2 41021 19998
0 20000 5 1 1 19999
0 20001 7 5 2 44265 61564
0 20002 5 1 1 64364
0 20003 7 2 2 53055 56031
0 20004 5 1 1 64369
0 20005 7 1 2 20004 64306
0 20006 5 1 1 20005
0 20007 7 1 2 46273 20006
0 20008 5 1 1 20007
0 20009 7 2 2 45714 57347
0 20010 7 1 2 61773 64371
0 20011 5 1 1 20010
0 20012 7 1 2 20008 20011
0 20013 5 1 1 20012
0 20014 7 1 2 48071 20013
0 20015 5 1 1 20014
0 20016 7 1 2 20015 64324
0 20017 5 1 1 20016
0 20018 7 1 2 49773 20017
0 20019 5 1 1 20018
0 20020 7 1 2 59661 64331
0 20021 5 1 1 20020
0 20022 7 1 2 64329 20021
0 20023 5 1 1 20022
0 20024 7 1 2 49519 20023
0 20025 5 1 1 20024
0 20026 7 1 2 55201 61920
0 20027 5 1 1 20026
0 20028 7 1 2 19840 20027
0 20029 5 1 1 20028
0 20030 7 1 2 42382 52419
0 20031 5 1 1 20030
0 20032 7 1 2 20029 20031
0 20033 5 1 1 20032
0 20034 7 3 2 53212 64361
0 20035 5 1 1 64373
0 20036 7 1 2 46274 64374
0 20037 5 1 1 20036
0 20038 7 1 2 20033 20037
0 20039 5 1 1 20038
0 20040 7 1 2 41667 20039
0 20041 5 1 1 20040
0 20042 7 1 2 52413 62553
0 20043 5 1 1 20042
0 20044 7 1 2 56728 20043
0 20045 5 1 1 20044
0 20046 7 1 2 54873 46688
0 20047 7 1 2 20045 20046
0 20048 5 1 1 20047
0 20049 7 1 2 20041 20048
0 20050 5 1 1 20049
0 20051 7 1 2 40860 20050
0 20052 5 1 1 20051
0 20053 7 1 2 64325 20052
0 20054 7 1 2 20025 20053
0 20055 5 1 1 20054
0 20056 7 1 2 45308 20055
0 20057 5 1 1 20056
0 20058 7 1 2 20019 20057
0 20059 5 1 1 20058
0 20060 7 1 2 64365 20059
0 20061 5 1 1 20060
0 20062 7 1 2 43215 20061
0 20063 7 1 2 20000 20062
0 20064 5 1 1 20063
0 20065 7 1 2 42835 56735
0 20066 5 2 1 20065
0 20067 7 1 2 51411 64376
0 20068 5 1 1 20067
0 20069 7 1 2 42627 20068
0 20070 5 1 1 20069
0 20071 7 1 2 53213 64357
0 20072 5 1 1 20071
0 20073 7 1 2 20070 20072
0 20074 5 1 1 20073
0 20075 7 1 2 43383 57828
0 20076 5 1 1 20075
0 20077 7 1 2 64288 20076
0 20078 7 1 2 20074 20077
0 20079 5 1 1 20078
0 20080 7 1 2 56688 54941
0 20081 7 1 2 63636 20080
0 20082 5 1 1 20081
0 20083 7 1 2 20079 20082
0 20084 5 1 1 20083
0 20085 7 1 2 40409 20084
0 20086 5 1 1 20085
0 20087 7 2 2 56986 57809
0 20088 7 1 2 40047 64378
0 20089 5 1 1 20088
0 20090 7 1 2 6044 20089
0 20091 5 1 1 20090
0 20092 7 1 2 48857 20091
0 20093 5 1 1 20092
0 20094 7 1 2 53542 57710
0 20095 7 1 2 53372 20094
0 20096 5 1 1 20095
0 20097 7 1 2 20093 20096
0 20098 5 1 1 20097
0 20099 7 1 2 42628 20098
0 20100 5 1 1 20099
0 20101 7 1 2 20086 20100
0 20102 5 1 1 20101
0 20103 7 1 2 57637 20102
0 20104 5 1 1 20103
0 20105 7 1 2 45715 64297
0 20106 5 2 1 20105
0 20107 7 1 2 51412 64380
0 20108 5 1 1 20107
0 20109 7 1 2 42629 48877
0 20110 7 1 2 20108 20109
0 20111 5 1 1 20110
0 20112 7 1 2 20035 20111
0 20113 5 1 1 20112
0 20114 7 1 2 43115 63298
0 20115 7 1 2 20113 20114
0 20116 5 1 1 20115
0 20117 7 1 2 20104 20116
0 20118 5 1 1 20117
0 20119 7 1 2 52094 20118
0 20120 5 1 1 20119
0 20121 7 6 2 41500 45104
0 20122 7 1 2 62020 64382
0 20123 7 1 2 57481 20122
0 20124 7 1 2 62997 20123
0 20125 5 1 1 20124
0 20126 7 2 2 62021 59050
0 20127 5 1 1 64388
0 20128 7 1 2 40048 58889
0 20129 5 1 1 20128
0 20130 7 1 2 20127 20129
0 20131 5 1 1 20130
0 20132 7 1 2 42988 20131
0 20133 7 1 2 64304 20132
0 20134 5 1 1 20133
0 20135 7 1 2 20125 20134
0 20136 5 1 1 20135
0 20137 7 1 2 51542 20136
0 20138 5 1 1 20137
0 20139 7 2 2 64308 63890
0 20140 5 1 1 64390
0 20141 7 1 2 51407 51947
0 20142 5 1 1 20141
0 20143 7 1 2 20140 20142
0 20144 5 1 1 20143
0 20145 7 1 2 46275 20144
0 20146 5 1 1 20145
0 20147 7 2 2 48691 53066
0 20148 7 1 2 57348 64392
0 20149 5 1 1 20148
0 20150 7 1 2 20146 20149
0 20151 5 1 1 20150
0 20152 7 1 2 43116 63313
0 20153 7 1 2 20151 20152
0 20154 5 1 1 20153
0 20155 7 1 2 20138 20154
0 20156 5 1 1 20155
0 20157 7 1 2 45716 20156
0 20158 5 1 1 20157
0 20159 7 1 2 40229 64379
0 20160 5 1 1 20159
0 20161 7 1 2 40049 57802
0 20162 5 1 1 20161
0 20163 7 1 2 20160 20162
0 20164 5 1 1 20163
0 20165 7 1 2 57638 64150
0 20166 7 1 2 20164 20165
0 20167 5 1 1 20166
0 20168 7 1 2 20158 20167
0 20169 5 1 1 20168
0 20170 7 1 2 46748 20169
0 20171 5 1 1 20170
0 20172 7 2 2 52042 64097
0 20173 5 1 1 64394
0 20174 7 1 2 58912 64395
0 20175 5 1 1 20174
0 20176 7 1 2 52710 57694
0 20177 5 1 1 20176
0 20178 7 1 2 6077 20177
0 20179 5 1 1 20178
0 20180 7 1 2 49520 58890
0 20181 7 1 2 20179 20180
0 20182 5 1 1 20181
0 20183 7 1 2 20175 20182
0 20184 5 1 1 20183
0 20185 7 1 2 57504 20184
0 20186 5 1 1 20185
0 20187 7 1 2 58265 49726
0 20188 5 1 1 20187
0 20189 7 5 2 41668 54444
0 20190 7 1 2 44803 64396
0 20191 7 2 2 20188 20190
0 20192 7 1 2 57639 57482
0 20193 7 1 2 64401 20192
0 20194 5 1 1 20193
0 20195 7 1 2 20186 20194
0 20196 5 1 1 20195
0 20197 7 1 2 42630 20196
0 20198 5 1 1 20197
0 20199 7 1 2 46494 20198
0 20200 7 1 2 20171 20199
0 20201 7 1 2 20120 20200
0 20202 5 1 1 20201
0 20203 7 1 2 58547 20202
0 20204 7 1 2 20064 20203
0 20205 5 1 1 20204
0 20206 7 1 2 44663 50570
0 20207 7 1 2 51181 20206
0 20208 5 1 1 20207
0 20209 7 1 2 46408 48878
0 20210 7 1 2 62598 20209
0 20211 7 1 2 59763 20210
0 20212 7 1 2 20208 20211
0 20213 5 1 1 20212
0 20214 7 1 2 58891 59575
0 20215 7 1 2 55490 20214
0 20216 5 1 1 20215
0 20217 7 1 2 20213 20216
0 20218 5 1 1 20217
0 20219 7 1 2 62412 20218
0 20220 5 1 1 20219
0 20221 7 1 2 57263 58548
0 20222 7 1 2 59524 20221
0 20223 7 1 2 64201 20222
0 20224 5 1 1 20223
0 20225 7 1 2 20220 20224
0 20226 5 1 1 20225
0 20227 7 1 2 63328 20226
0 20228 5 1 1 20227
0 20229 7 5 2 44804 53461
0 20230 7 1 2 53381 64403
0 20231 5 1 1 20230
0 20232 7 2 2 42383 56032
0 20233 5 1 1 64408
0 20234 7 1 2 20231 20233
0 20235 5 1 1 20234
0 20236 7 1 2 40410 20235
0 20237 5 1 1 20236
0 20238 7 1 2 63281 57915
0 20239 5 1 1 20238
0 20240 7 1 2 20237 20239
0 20241 5 1 1 20240
0 20242 7 1 2 41119 20241
0 20243 5 1 1 20242
0 20244 7 1 2 57586 64409
0 20245 5 1 1 20244
0 20246 7 1 2 20243 20245
0 20247 5 1 1 20246
0 20248 7 1 2 40050 20247
0 20249 5 1 1 20248
0 20250 7 2 2 54530 51418
0 20251 5 1 1 64410
0 20252 7 1 2 40630 49307
0 20253 7 1 2 64411 20252
0 20254 5 1 1 20253
0 20255 7 1 2 20249 20254
0 20256 5 1 1 20255
0 20257 7 1 2 59138 20256
0 20258 5 1 1 20257
0 20259 7 1 2 56392 63760
0 20260 5 1 1 20259
0 20261 7 1 2 20260 64158
0 20262 5 1 1 20261
0 20263 7 1 2 58414 20262
0 20264 5 1 1 20263
0 20265 7 1 2 20258 20264
0 20266 5 1 1 20265
0 20267 7 1 2 40230 20266
0 20268 5 1 1 20267
0 20269 7 1 2 57434 64237
0 20270 5 1 1 20269
0 20271 7 1 2 49446 56188
0 20272 5 1 1 20271
0 20273 7 1 2 63282 20272
0 20274 5 1 1 20273
0 20275 7 1 2 20270 20274
0 20276 5 1 1 20275
0 20277 7 1 2 41120 20276
0 20278 5 1 1 20277
0 20279 7 1 2 54709 55848
0 20280 5 1 1 20279
0 20281 7 1 2 20278 20280
0 20282 5 1 1 20281
0 20283 7 1 2 40051 20282
0 20284 5 1 1 20283
0 20285 7 1 2 42384 46848
0 20286 5 2 1 20285
0 20287 7 1 2 64412 64157
0 20288 5 1 1 20287
0 20289 7 1 2 20284 20288
0 20290 5 1 1 20289
0 20291 7 1 2 58415 20290
0 20292 5 1 1 20291
0 20293 7 1 2 20268 20292
0 20294 5 1 1 20293
0 20295 7 1 2 46566 20294
0 20296 5 1 1 20295
0 20297 7 8 2 57640 58549
0 20298 7 2 2 43117 64414
0 20299 7 1 2 53365 63761
0 20300 5 1 1 20299
0 20301 7 1 2 64159 20300
0 20302 5 1 1 20301
0 20303 7 1 2 52095 20302
0 20304 5 1 1 20303
0 20305 7 1 2 63283 58261
0 20306 5 1 1 20305
0 20307 7 1 2 51686 63762
0 20308 5 1 1 20307
0 20309 7 1 2 63284 60552
0 20310 5 1 1 20309
0 20311 7 1 2 20308 20310
0 20312 5 1 1 20311
0 20313 7 1 2 46749 20312
0 20314 5 1 1 20313
0 20315 7 1 2 20306 20314
0 20316 7 1 2 20304 20315
0 20317 5 1 1 20316
0 20318 7 1 2 64422 20317
0 20319 5 1 1 20318
0 20320 7 1 2 20296 20319
0 20321 5 1 1 20320
0 20322 7 1 2 46495 20321
0 20323 5 1 1 20322
0 20324 7 1 2 57435 51687
0 20325 7 1 2 63320 20324
0 20326 5 1 1 20325
0 20327 7 1 2 4202 20326
0 20328 5 1 1 20327
0 20329 7 1 2 63550 20328
0 20330 5 1 1 20329
0 20331 7 2 2 46628 57180
0 20332 7 1 2 49316 64404
0 20333 7 1 2 64424 20332
0 20334 5 1 1 20333
0 20335 7 1 2 48394 56033
0 20336 7 1 2 59139 20335
0 20337 5 1 1 20336
0 20338 7 1 2 20334 20337
0 20339 7 1 2 20330 20338
0 20340 5 1 1 20339
0 20341 7 1 2 49521 20340
0 20342 5 1 1 20341
0 20343 7 1 2 42631 63463
0 20344 5 1 1 20343
0 20345 7 1 2 20344 63880
0 20346 5 1 1 20345
0 20347 7 1 2 63551 20346
0 20348 5 1 1 20347
0 20349 7 1 2 52269 63526
0 20350 5 1 1 20349
0 20351 7 1 2 49774 56034
0 20352 5 1 1 20351
0 20353 7 1 2 20350 20352
0 20354 5 1 1 20353
0 20355 7 1 2 45717 59140
0 20356 7 1 2 20354 20355
0 20357 5 1 1 20356
0 20358 7 1 2 40231 59426
0 20359 7 1 2 49944 20358
0 20360 7 1 2 63754 20359
0 20361 5 1 1 20360
0 20362 7 1 2 20357 20361
0 20363 7 1 2 20348 20362
0 20364 7 1 2 20342 20363
0 20365 5 1 1 20364
0 20366 7 1 2 59336 20365
0 20367 5 1 1 20366
0 20368 7 1 2 49323 58257
0 20369 5 1 1 20368
0 20370 7 1 2 61431 20369
0 20371 5 1 1 20370
0 20372 7 2 2 44421 45105
0 20373 5 2 1 64426
0 20374 7 2 2 64428 62028
0 20375 7 2 2 41022 62083
0 20376 5 1 1 64432
0 20377 7 1 2 64430 64433
0 20378 5 1 1 20377
0 20379 7 1 2 46941 64366
0 20380 5 1 1 20379
0 20381 7 1 2 20378 20380
0 20382 5 1 1 20381
0 20383 7 1 2 55678 20382
0 20384 5 1 1 20383
0 20385 7 1 2 20371 20384
0 20386 5 1 1 20385
0 20387 7 1 2 46567 20386
0 20388 5 1 1 20387
0 20389 7 1 2 52291 64423
0 20390 5 1 1 20389
0 20391 7 1 2 20388 20390
0 20392 5 1 1 20391
0 20393 7 1 2 46496 20392
0 20394 5 1 1 20393
0 20395 7 1 2 55160 59141
0 20396 5 1 1 20395
0 20397 7 1 2 61437 20396
0 20398 5 1 1 20397
0 20399 7 1 2 59337 20398
0 20400 5 1 1 20399
0 20401 7 1 2 20394 20400
0 20402 5 1 1 20401
0 20403 7 1 2 48692 20402
0 20404 5 1 1 20403
0 20405 7 2 2 41806 57405
0 20406 5 1 1 64434
0 20407 7 1 2 46806 59051
0 20408 5 1 1 20407
0 20409 7 1 2 20406 20408
0 20410 5 1 1 20409
0 20411 7 1 2 41023 20410
0 20412 5 1 1 20411
0 20413 7 1 2 46807 64367
0 20414 5 1 1 20413
0 20415 7 1 2 20412 20414
0 20416 5 1 1 20415
0 20417 7 1 2 40052 20416
0 20418 5 1 1 20417
0 20419 7 1 2 46808 61432
0 20420 5 1 1 20419
0 20421 7 1 2 20418 20420
0 20422 5 1 1 20421
0 20423 7 1 2 40232 41051
0 20424 7 1 2 49522 20423
0 20425 7 2 2 59681 20424
0 20426 7 1 2 20422 64436
0 20427 5 1 1 20426
0 20428 7 1 2 20404 20427
0 20429 5 1 1 20428
0 20430 7 1 2 52455 20429
0 20431 5 1 1 20430
0 20432 7 1 2 50331 63064
0 20433 7 1 2 58550 20432
0 20434 7 2 2 41807 47277
0 20435 7 3 2 43216 57683
0 20436 7 1 2 64438 64440
0 20437 7 1 2 20433 20436
0 20438 5 1 1 20437
0 20439 7 1 2 20431 20438
0 20440 5 1 1 20439
0 20441 7 1 2 49671 20440
0 20442 5 1 1 20441
0 20443 7 1 2 20367 20442
0 20444 7 1 2 20323 20443
0 20445 5 1 1 20444
0 20446 7 1 2 46124 20445
0 20447 5 1 1 20446
0 20448 7 1 2 59682 52998
0 20449 5 1 1 20448
0 20450 7 1 2 52990 59529
0 20451 5 1 1 20450
0 20452 7 1 2 20449 20451
0 20453 5 1 1 20452
0 20454 7 1 2 41052 20453
0 20455 5 1 1 20454
0 20456 7 1 2 52991 59564
0 20457 5 1 1 20456
0 20458 7 1 2 20455 20457
0 20459 5 1 1 20458
0 20460 7 1 2 59142 20459
0 20461 5 1 1 20460
0 20462 7 2 2 46497 52096
0 20463 7 1 2 59764 64443
0 20464 5 1 1 20463
0 20465 7 1 2 20464 8280
0 20466 5 1 1 20465
0 20467 7 1 2 41366 20466
0 20468 5 1 1 20467
0 20469 7 2 2 45309 58551
0 20470 7 2 2 40233 64445
0 20471 7 1 2 41121 60464
0 20472 7 1 2 64447 20471
0 20473 5 1 1 20472
0 20474 7 1 2 20468 20473
0 20475 5 1 1 20474
0 20476 7 1 2 43118 20475
0 20477 5 1 1 20476
0 20478 7 1 2 20461 20477
0 20479 5 1 1 20478
0 20480 7 1 2 40411 20479
0 20481 5 1 1 20480
0 20482 7 1 2 55679 59345
0 20483 5 1 1 20482
0 20484 7 1 2 8143 20483
0 20485 5 1 1 20484
0 20486 7 1 2 59143 20485
0 20487 5 1 1 20486
0 20488 7 1 2 63603 59765
0 20489 5 1 1 20488
0 20490 7 1 2 20487 20489
0 20491 5 1 1 20490
0 20492 7 1 2 48693 20491
0 20493 5 1 1 20492
0 20494 7 1 2 64425 64437
0 20495 5 1 1 20494
0 20496 7 1 2 20493 20495
0 20497 5 1 1 20496
0 20498 7 1 2 46750 20497
0 20499 5 1 1 20498
0 20500 7 1 2 50032 64448
0 20501 7 1 2 63554 20500
0 20502 5 1 1 20501
0 20503 7 1 2 20499 20502
0 20504 7 1 2 20481 20503
0 20505 5 1 1 20504
0 20506 7 1 2 48509 55511
0 20507 7 1 2 20505 20506
0 20508 5 1 1 20507
0 20509 7 1 2 20447 20508
0 20510 5 1 1 20509
0 20511 7 1 2 46276 20510
0 20512 5 1 1 20511
0 20513 7 1 2 20228 20512
0 20514 5 1 1 20513
0 20515 7 1 2 49206 20514
0 20516 5 1 1 20515
0 20517 7 1 2 53003 63981
0 20518 5 1 1 20517
0 20519 7 1 2 56987 50930
0 20520 5 1 1 20519
0 20521 7 1 2 20518 20520
0 20522 5 1 1 20521
0 20523 7 1 2 52292 20522
0 20524 5 1 1 20523
0 20525 7 1 2 20524 20173
0 20526 5 1 1 20525
0 20527 7 1 2 42632 20526
0 20528 5 1 1 20527
0 20529 7 1 2 52293 64375
0 20530 5 1 1 20529
0 20531 7 1 2 20528 20530
0 20532 5 1 1 20531
0 20533 7 1 2 20532 63258
0 20534 5 1 1 20533
0 20535 7 1 2 48858 57542
0 20536 5 1 1 20535
0 20537 7 1 2 47278 57926
0 20538 5 1 1 20537
0 20539 7 1 2 20536 20538
0 20540 5 1 1 20539
0 20541 7 1 2 40412 20540
0 20542 5 1 1 20541
0 20543 7 1 2 56704 48219
0 20544 7 1 2 59891 20543
0 20545 5 1 1 20544
0 20546 7 1 2 20542 20545
0 20547 5 1 1 20546
0 20548 7 1 2 57798 20547
0 20549 5 1 1 20548
0 20550 7 1 2 57436 56519
0 20551 5 1 1 20550
0 20552 7 1 2 55213 55591
0 20553 5 1 1 20552
0 20554 7 1 2 20551 20553
0 20555 5 1 1 20554
0 20556 7 1 2 41122 20555
0 20557 5 1 1 20556
0 20558 7 1 2 64309 56739
0 20559 5 1 1 20558
0 20560 7 1 2 20557 20559
0 20561 5 1 1 20560
0 20562 7 1 2 40413 20561
0 20563 5 1 1 20562
0 20564 7 1 2 57780 51398
0 20565 7 1 2 57916 20564
0 20566 5 1 1 20565
0 20567 7 1 2 48859 53076
0 20568 5 1 1 20567
0 20569 7 1 2 20566 20568
0 20570 5 1 1 20569
0 20571 7 1 2 40053 20570
0 20572 5 1 1 20571
0 20573 7 1 2 56075 63460
0 20574 5 1 1 20573
0 20575 7 1 2 20572 20574
0 20576 5 1 1 20575
0 20577 7 1 2 42633 20576
0 20578 5 1 1 20577
0 20579 7 1 2 20563 20578
0 20580 5 1 1 20579
0 20581 7 1 2 46277 20580
0 20582 5 1 1 20581
0 20583 7 1 2 64393 64372
0 20584 5 1 1 20583
0 20585 7 1 2 20582 20584
0 20586 5 1 1 20585
0 20587 7 1 2 48072 20586
0 20588 5 1 1 20587
0 20589 7 1 2 53013 56520
0 20590 5 1 1 20589
0 20591 7 1 2 42634 53077
0 20592 5 1 1 20591
0 20593 7 1 2 20590 20592
0 20594 5 1 1 20593
0 20595 7 1 2 46278 20594
0 20596 5 1 1 20595
0 20597 7 1 2 64257 20596
0 20598 5 1 1 20597
0 20599 7 1 2 48073 20598
0 20600 5 1 1 20599
0 20601 7 1 2 64276 64036
0 20602 5 1 1 20601
0 20603 7 1 2 20600 20602
0 20604 5 1 1 20603
0 20605 7 1 2 40414 20604
0 20606 5 1 1 20605
0 20607 7 1 2 54874 47230
0 20608 7 1 2 62616 20607
0 20609 5 1 1 20608
0 20610 7 1 2 20606 20609
0 20611 5 1 1 20610
0 20612 7 1 2 46751 20611
0 20613 5 1 1 20612
0 20614 7 2 2 41123 60824
0 20615 7 1 2 64449 64322
0 20616 5 1 1 20615
0 20617 7 1 2 20613 20616
0 20618 7 1 2 20588 20617
0 20619 5 1 1 20618
0 20620 7 1 2 40234 20619
0 20621 5 1 1 20620
0 20622 7 1 2 20549 20621
0 20623 5 1 1 20622
0 20624 7 1 2 55068 20623
0 20625 5 1 1 20624
0 20626 7 1 2 20534 20625
0 20627 5 1 1 20626
0 20628 7 1 2 46409 20627
0 20629 5 1 1 20628
0 20630 7 1 2 54445 56021
0 20631 5 2 1 20630
0 20632 7 4 2 44109 56797
0 20633 7 1 2 53291 50147
0 20634 7 1 2 64453 20633
0 20635 5 1 1 20634
0 20636 7 2 2 64451 20635
0 20637 5 1 1 64457
0 20638 7 2 2 46125 20637
0 20639 7 1 2 40235 64459
0 20640 5 1 1 20639
0 20641 7 1 2 48074 64391
0 20642 5 1 1 20641
0 20643 7 1 2 20640 20642
0 20644 5 1 1 20643
0 20645 7 1 2 45718 20644
0 20646 5 1 1 20645
0 20647 7 3 2 41669 56766
0 20648 7 1 2 64461 64370
0 20649 5 1 1 20648
0 20650 7 1 2 20646 20649
0 20651 5 1 1 20650
0 20652 7 1 2 46279 20651
0 20653 5 1 1 20652
0 20654 7 2 2 56720 57360
0 20655 7 1 2 64224 56339
0 20656 7 1 2 57596 20655
0 20657 7 1 2 64464 20656
0 20658 5 1 1 20657
0 20659 7 1 2 20653 20658
0 20660 5 1 1 20659
0 20661 7 1 2 46752 20660
0 20662 5 1 1 20661
0 20663 7 1 2 55276 63891
0 20664 5 1 1 20663
0 20665 7 1 2 40054 64460
0 20666 5 1 1 20665
0 20667 7 1 2 20664 20666
0 20668 5 1 1 20667
0 20669 7 1 2 45719 20668
0 20670 5 1 1 20669
0 20671 7 1 2 48075 64151
0 20672 7 1 2 56988 20671
0 20673 5 1 1 20672
0 20674 7 1 2 20670 20673
0 20675 5 1 1 20674
0 20676 7 1 2 46280 20675
0 20677 5 1 1 20676
0 20678 7 1 2 20677 64333
0 20679 5 1 1 20678
0 20680 7 1 2 52097 20679
0 20681 5 1 1 20680
0 20682 7 1 2 63479 64402
0 20683 5 1 1 20682
0 20684 7 1 2 20681 20683
0 20685 7 1 2 20662 20684
0 20686 5 1 1 20685
0 20687 7 1 2 58416 20686
0 20688 5 1 1 20687
0 20689 7 1 2 20629 20688
0 20690 5 1 1 20689
0 20691 7 1 2 59346 20690
0 20692 5 1 1 20691
0 20693 7 1 2 20516 20692
0 20694 7 1 2 20205 20693
0 20695 5 1 1 20694
0 20696 7 1 2 49032 20695
0 20697 5 1 1 20696
0 20698 7 2 2 48440 63098
0 20699 5 1 1 64466
0 20700 7 1 2 57884 20699
0 20701 5 1 1 20700
0 20702 7 1 2 48879 20701
0 20703 5 1 1 20702
0 20704 7 1 2 48694 50656
0 20705 7 1 2 48274 20704
0 20706 5 1 1 20705
0 20707 7 1 2 43717 53370
0 20708 5 1 1 20707
0 20709 7 1 2 50808 51272
0 20710 7 1 2 20708 20709
0 20711 5 1 1 20710
0 20712 7 1 2 20706 20711
0 20713 5 1 1 20712
0 20714 7 1 2 44110 20713
0 20715 5 1 1 20714
0 20716 7 1 2 52924 62554
0 20717 5 1 1 20716
0 20718 7 1 2 63120 20717
0 20719 5 1 1 20718
0 20720 7 1 2 42989 53313
0 20721 7 1 2 20719 20720
0 20722 5 1 1 20721
0 20723 7 1 2 20715 20722
0 20724 7 1 2 20703 20723
0 20725 5 1 1 20724
0 20726 7 1 2 52098 20725
0 20727 5 1 1 20726
0 20728 7 1 2 19325 20727
0 20729 5 1 1 20728
0 20730 7 1 2 53988 20729
0 20731 5 1 1 20730
0 20732 7 1 2 48117 61921
0 20733 5 1 1 20732
0 20734 7 1 2 52823 20733
0 20735 5 1 1 20734
0 20736 7 1 2 40055 20735
0 20737 5 1 1 20736
0 20738 7 1 2 57781 50784
0 20739 5 1 1 20738
0 20740 7 1 2 20737 20739
0 20741 5 1 1 20740
0 20742 7 1 2 44954 20741
0 20743 5 1 1 20742
0 20744 7 1 2 42990 63667
0 20745 7 1 2 64302 20744
0 20746 5 1 1 20745
0 20747 7 1 2 20743 20746
0 20748 5 1 1 20747
0 20749 7 1 2 40236 20748
0 20750 5 1 1 20749
0 20751 7 2 2 52925 61922
0 20752 5 1 1 64468
0 20753 7 1 2 49600 49091
0 20754 5 2 1 20753
0 20755 7 1 2 20752 64470
0 20756 5 1 1 20755
0 20757 7 1 2 47279 52786
0 20758 7 1 2 20756 20757
0 20759 5 1 1 20758
0 20760 7 1 2 20750 20759
0 20761 5 1 1 20760
0 20762 7 1 2 45720 20761
0 20763 5 1 1 20762
0 20764 7 7 2 40056 52099
0 20765 7 1 2 49523 64472
0 20766 5 1 1 20765
0 20767 7 2 2 58273 20766
0 20768 5 1 1 64479
0 20769 7 1 2 64095 64471
0 20770 5 1 1 20769
0 20771 7 1 2 42991 20770
0 20772 5 1 1 20771
0 20773 7 1 2 49601 56222
0 20774 5 1 1 20773
0 20775 7 1 2 20772 20774
0 20776 5 1 1 20775
0 20777 7 1 2 20768 20776
0 20778 5 1 1 20777
0 20779 7 1 2 40861 20778
0 20780 7 1 2 20763 20779
0 20781 5 1 1 20780
0 20782 7 2 2 40057 57917
0 20783 5 1 1 64481
0 20784 7 1 2 40415 47973
0 20785 5 1 1 20784
0 20786 7 1 2 20783 20785
0 20787 5 1 1 20786
0 20788 7 1 2 50809 20787
0 20789 5 1 1 20788
0 20790 7 1 2 64381 20789
0 20791 5 1 1 20790
0 20792 7 1 2 41124 20791
0 20793 5 1 1 20792
0 20794 7 1 2 41501 50931
0 20795 5 1 1 20794
0 20796 7 1 2 54125 20795
0 20797 5 1 1 20796
0 20798 7 1 2 40631 20797
0 20799 5 1 1 20798
0 20800 7 1 2 45721 61799
0 20801 5 1 1 20800
0 20802 7 1 2 20799 20801
0 20803 5 2 1 20802
0 20804 7 1 2 64310 64483
0 20805 5 1 1 20804
0 20806 7 1 2 20793 20805
0 20807 5 1 1 20806
0 20808 7 1 2 40237 20807
0 20809 5 1 1 20808
0 20810 7 1 2 56860 64112
0 20811 5 1 1 20810
0 20812 7 1 2 44955 20811
0 20813 7 1 2 20809 20812
0 20814 5 1 1 20813
0 20815 7 1 2 45722 49685
0 20816 5 1 1 20815
0 20817 7 1 2 64480 20816
0 20818 5 1 1 20817
0 20819 7 1 2 56618 20818
0 20820 5 1 1 20819
0 20821 7 1 2 41670 20820
0 20822 5 1 1 20821
0 20823 7 1 2 46281 20822
0 20824 7 1 2 20814 20823
0 20825 5 1 1 20824
0 20826 7 1 2 64473 64484
0 20827 5 1 1 20826
0 20828 7 1 2 48510 58278
0 20829 5 1 1 20828
0 20830 7 1 2 20827 20829
0 20831 5 1 1 20830
0 20832 7 1 2 51644 20831
0 20833 5 1 1 20832
0 20834 7 1 2 44111 20833
0 20835 7 1 2 20825 20834
0 20836 5 1 1 20835
0 20837 7 1 2 54163 20836
0 20838 7 1 2 20781 20837
0 20839 5 1 1 20838
0 20840 7 1 2 20731 20839
0 20841 5 1 1 20840
0 20842 7 1 2 42635 20841
0 20843 5 1 1 20842
0 20844 7 1 2 57092 57901
0 20845 5 1 1 20844
0 20846 7 2 2 63415 56767
0 20847 7 1 2 49092 64485
0 20848 5 1 1 20847
0 20849 7 1 2 44805 55173
0 20850 7 1 2 53048 20849
0 20851 5 1 1 20850
0 20852 7 1 2 20848 20851
0 20853 5 1 1 20852
0 20854 7 1 2 54611 20853
0 20855 5 1 1 20854
0 20856 7 1 2 20845 20855
0 20857 5 1 1 20856
0 20858 7 1 2 52100 20857
0 20859 5 1 1 20858
0 20860 7 3 2 42836 57957
0 20861 7 1 2 64487 64088
0 20862 7 1 2 63985 20861
0 20863 5 1 1 20862
0 20864 7 1 2 20859 20863
0 20865 5 1 1 20864
0 20866 7 2 2 40416 20865
0 20867 7 1 2 64071 64490
0 20868 5 1 1 20867
0 20869 7 1 2 20843 20868
0 20870 5 1 1 20869
0 20871 7 1 2 46498 20870
0 20872 5 1 1 20871
0 20873 7 1 2 52068 58279
0 20874 5 1 1 20873
0 20875 7 1 2 54126 20874
0 20876 5 2 1 20875
0 20877 7 1 2 40058 64492
0 20878 5 1 1 20877
0 20879 7 1 2 52987 50421
0 20880 5 2 1 20879
0 20881 7 1 2 20878 64494
0 20882 5 1 1 20881
0 20883 7 2 2 48511 20882
0 20884 7 2 2 55410 60510
0 20885 7 1 2 56567 64498
0 20886 7 1 2 64496 20885
0 20887 5 1 1 20886
0 20888 7 1 2 20872 20887
0 20889 5 1 1 20888
0 20890 7 1 2 46629 20889
0 20891 5 1 1 20890
0 20892 7 2 2 40238 46689
0 20893 7 7 2 40417 42385
0 20894 5 1 1 64502
0 20895 7 1 2 54164 64503
0 20896 7 1 2 64500 20895
0 20897 5 1 1 20896
0 20898 7 1 2 61118 20897
0 20899 5 1 1 20898
0 20900 7 1 2 64165 20899
0 20901 5 1 1 20900
0 20902 7 1 2 45723 64469
0 20903 5 1 1 20902
0 20904 7 1 2 52143 59887
0 20905 5 1 1 20904
0 20906 7 1 2 20903 20905
0 20907 5 1 1 20906
0 20908 7 1 2 57052 61962
0 20909 7 1 2 20907 20908
0 20910 5 1 1 20909
0 20911 7 1 2 20901 20910
0 20912 5 1 1 20911
0 20913 7 1 2 40059 20912
0 20914 5 1 1 20913
0 20915 7 1 2 42992 57122
0 20916 5 1 1 20915
0 20917 7 1 2 56934 20916
0 20918 5 1 1 20917
0 20919 7 1 2 49524 20918
0 20920 5 1 1 20919
0 20921 7 1 2 55298 61923
0 20922 5 1 1 20921
0 20923 7 1 2 57878 20922
0 20924 5 1 1 20923
0 20925 7 1 2 51290 20924
0 20926 5 1 1 20925
0 20927 7 1 2 20920 20926
0 20928 5 1 1 20927
0 20929 7 1 2 54165 20928
0 20930 5 1 1 20929
0 20931 7 1 2 55333 53543
0 20932 7 1 2 57733 20931
0 20933 5 1 1 20932
0 20934 7 1 2 20930 20933
0 20935 5 1 1 20934
0 20936 7 1 2 40239 20935
0 20937 5 1 1 20936
0 20938 7 1 2 20914 20937
0 20939 5 1 1 20938
0 20940 7 1 2 42636 20939
0 20941 5 1 1 20940
0 20942 7 1 2 61991 53533
0 20943 5 1 1 20942
0 20944 7 5 2 54686 55430
0 20945 5 1 1 64509
0 20946 7 2 2 41502 64510
0 20947 7 1 2 64514 62400
0 20948 5 1 1 20947
0 20949 7 1 2 20943 20948
0 20950 5 1 1 20949
0 20951 7 1 2 49525 20950
0 20952 5 1 1 20951
0 20953 7 1 2 44112 61924
0 20954 5 1 1 20953
0 20955 7 1 2 53523 20954
0 20956 5 1 1 20955
0 20957 7 1 2 56815 63620
0 20958 7 1 2 20956 20957
0 20959 5 1 1 20958
0 20960 7 1 2 20952 20959
0 20961 5 1 1 20960
0 20962 7 1 2 42637 20961
0 20963 5 1 1 20962
0 20964 7 2 2 44113 61776
0 20965 7 2 2 45724 52624
0 20966 7 1 2 54864 57181
0 20967 7 1 2 64518 20966
0 20968 7 1 2 64516 20967
0 20969 5 1 1 20968
0 20970 7 1 2 20963 20969
0 20971 5 1 1 20970
0 20972 7 1 2 48275 20971
0 20973 5 1 1 20972
0 20974 7 1 2 48220 63809
0 20975 5 1 1 20974
0 20976 7 1 2 57902 20975
0 20977 5 1 1 20976
0 20978 7 1 2 46410 20977
0 20979 5 1 1 20978
0 20980 7 1 2 48076 57789
0 20981 5 1 1 20980
0 20982 7 1 2 20979 20981
0 20983 5 1 1 20982
0 20984 7 1 2 60827 20983
0 20985 5 1 1 20984
0 20986 7 1 2 62122 63675
0 20987 7 1 2 6168 20986
0 20988 5 1 1 20987
0 20989 7 1 2 20985 20988
0 20990 5 1 1 20989
0 20991 7 1 2 64238 20990
0 20992 5 1 1 20991
0 20993 7 1 2 20973 20992
0 20994 7 1 2 20941 20993
0 20995 5 1 1 20994
0 20996 7 1 2 46499 20995
0 20997 5 1 1 20996
0 20998 7 1 2 57300 56776
0 20999 7 1 2 59925 20998
0 21000 7 1 2 64058 20999
0 21001 5 1 1 21000
0 21002 7 1 2 20997 21001
0 21003 5 1 1 21002
0 21004 7 1 2 46630 21003
0 21005 5 1 1 21004
0 21006 7 3 2 56572 63688
0 21007 7 2 2 64225 64520
0 21008 7 2 2 54654 52231
0 21009 7 2 2 41503 60341
0 21010 7 1 2 61831 55431
0 21011 7 1 2 64527 21010
0 21012 7 1 2 64525 21011
0 21013 7 1 2 64523 21012
0 21014 5 1 1 21013
0 21015 7 1 2 21005 21014
0 21016 5 1 1 21015
0 21017 7 1 2 46753 21016
0 21018 5 1 1 21017
0 21019 7 1 2 64349 62617
0 21020 7 1 2 62067 64031
0 21021 7 1 2 21019 21020
0 21022 7 1 2 64521 21021
0 21023 5 1 1 21022
0 21024 7 1 2 21018 21023
0 21025 7 1 2 20891 21024
0 21026 5 1 1 21025
0 21027 7 1 2 46568 21026
0 21028 5 1 1 21027
0 21029 7 1 2 326 48146
0 21030 5 2 1 21029
0 21031 7 1 2 49602 64529
0 21032 5 1 1 21031
0 21033 7 1 2 60677 64220
0 21034 5 1 1 21033
0 21035 7 1 2 21032 21034
0 21036 5 1 1 21035
0 21037 7 1 2 42638 21036
0 21038 5 1 1 21037
0 21039 7 1 2 40862 50622
0 21040 5 2 1 21039
0 21041 7 1 2 44114 63825
0 21042 5 1 1 21041
0 21043 7 1 2 64531 21042
0 21044 5 1 1 21043
0 21045 7 1 2 52621 21044
0 21046 5 1 1 21045
0 21047 7 1 2 21038 21046
0 21048 5 1 1 21047
0 21049 7 1 2 60290 21048
0 21050 5 1 1 21049
0 21051 7 1 2 60465 56768
0 21052 7 1 2 58789 21051
0 21053 7 1 2 1738 21052
0 21054 5 1 1 21053
0 21055 7 1 2 21050 21054
0 21056 5 1 1 21055
0 21057 7 1 2 46411 21056
0 21058 5 1 1 21057
0 21059 7 1 2 48860 61816
0 21060 5 1 1 21059
0 21061 7 2 2 52002 61289
0 21062 5 1 1 64533
0 21063 7 1 2 21060 21062
0 21064 5 1 1 21063
0 21065 7 1 2 51487 62192
0 21066 7 1 2 53544 21065
0 21067 7 1 2 21064 21066
0 21068 5 1 1 21067
0 21069 7 1 2 21058 21068
0 21070 5 1 1 21069
0 21071 7 1 2 48915 21070
0 21072 5 1 1 21071
0 21073 7 1 2 53084 16356
0 21074 5 1 1 21073
0 21075 7 1 2 44115 21074
0 21076 5 1 1 21075
0 21077 7 1 2 64532 21076
0 21078 5 1 1 21077
0 21079 7 1 2 45942 21078
0 21080 5 1 1 21079
0 21081 7 1 2 55743 60678
0 21082 5 1 1 21081
0 21083 7 1 2 21080 21082
0 21084 5 1 1 21083
0 21085 7 1 2 45725 21084
0 21086 5 1 1 21085
0 21087 7 1 2 54512 16309
0 21088 5 1 1 21087
0 21089 7 1 2 40632 21088
0 21090 5 1 1 21089
0 21091 7 1 2 40863 54287
0 21092 7 1 2 2621 21091
0 21093 5 1 1 21092
0 21094 7 1 2 21090 21093
0 21095 5 1 1 21094
0 21096 7 1 2 53004 21095
0 21097 5 1 1 21096
0 21098 7 1 2 21086 21097
0 21099 5 1 1 21098
0 21100 7 5 2 43217 54980
0 21101 7 1 2 61976 64535
0 21102 7 1 2 21099 21101
0 21103 5 1 1 21102
0 21104 7 1 2 41671 21103
0 21105 7 1 2 21072 21104
0 21106 5 1 1 21105
0 21107 7 1 2 62038 57354
0 21108 5 1 1 21107
0 21109 7 2 2 52537 63341
0 21110 7 2 2 46282 61868
0 21111 7 1 2 60659 64542
0 21112 7 1 2 64540 21111
0 21113 5 1 1 21112
0 21114 7 1 2 21108 21113
0 21115 5 1 1 21114
0 21116 7 1 2 45726 21115
0 21117 5 1 1 21116
0 21118 7 2 2 44266 46283
0 21119 7 1 2 52383 64544
0 21120 7 1 2 56506 21119
0 21121 7 1 2 61943 21120
0 21122 5 1 1 21121
0 21123 7 1 2 21117 21122
0 21124 5 1 1 21123
0 21125 7 1 2 44116 21124
0 21126 5 1 1 21125
0 21127 7 2 2 48118 53314
0 21128 5 1 1 64546
0 21129 7 1 2 50776 56603
0 21130 5 1 1 21129
0 21131 7 1 2 21128 21130
0 21132 5 1 1 21131
0 21133 7 1 2 60714 62376
0 21134 7 1 2 21132 21133
0 21135 5 1 1 21134
0 21136 7 1 2 21126 21135
0 21137 5 1 1 21136
0 21138 7 1 2 40060 21137
0 21139 5 1 1 21138
0 21140 7 2 2 48221 62992
0 21141 5 1 1 64548
0 21142 7 1 2 40864 55270
0 21143 5 1 1 21142
0 21144 7 1 2 51665 57974
0 21145 5 1 1 21144
0 21146 7 1 2 21143 21145
0 21147 5 1 1 21146
0 21148 7 1 2 42993 21147
0 21149 5 1 1 21148
0 21150 7 1 2 21141 21149
0 21151 5 1 1 21150
0 21152 7 1 2 41504 21151
0 21153 5 1 1 21152
0 21154 7 1 2 53386 48142
0 21155 5 1 1 21154
0 21156 7 1 2 21153 21155
0 21157 5 1 1 21156
0 21158 7 1 2 21157 63569
0 21159 5 1 1 21158
0 21160 7 1 2 45727 57514
0 21161 5 1 1 21160
0 21162 7 1 2 64183 21161
0 21163 5 1 1 21162
0 21164 7 1 2 54981 61916
0 21165 7 1 2 21163 21164
0 21166 5 1 1 21165
0 21167 7 1 2 21159 21166
0 21168 5 1 1 21167
0 21169 7 1 2 40633 21168
0 21170 5 1 1 21169
0 21171 7 3 2 50748 59001
0 21172 7 1 2 64550 61861
0 21173 5 1 1 21172
0 21174 7 2 2 43119 48861
0 21175 7 2 2 53904 64553
0 21176 5 1 1 64555
0 21177 7 1 2 64556 60466
0 21178 5 1 1 21177
0 21179 7 1 2 21173 21178
0 21180 5 1 1 21179
0 21181 7 1 2 56946 21180
0 21182 5 1 1 21181
0 21183 7 2 2 45106 42837
0 21184 7 2 2 44267 64557
0 21185 7 1 2 61164 64559
0 21186 7 1 2 64543 21185
0 21187 5 1 1 21186
0 21188 7 1 2 21182 21187
0 21189 5 1 1 21188
0 21190 7 1 2 42639 21189
0 21191 5 1 1 21190
0 21192 7 1 2 57975 63629
0 21193 7 1 2 63862 21192
0 21194 5 1 1 21193
0 21195 7 1 2 21191 21194
0 21196 5 1 1 21195
0 21197 7 1 2 40865 21196
0 21198 5 1 1 21197
0 21199 7 1 2 44956 21198
0 21200 7 1 2 21170 21199
0 21201 7 1 2 21139 21200
0 21202 5 1 1 21201
0 21203 7 1 2 21106 21202
0 21204 5 1 1 21203
0 21205 7 2 2 60577 63073
0 21206 7 1 2 53905 64561
0 21207 7 1 2 62618 21206
0 21208 7 1 2 63215 21207
0 21209 5 1 1 21208
0 21210 7 1 2 21204 21209
0 21211 5 1 1 21210
0 21212 7 1 2 40418 21211
0 21213 5 1 1 21212
0 21214 7 1 2 5199 64377
0 21215 5 1 1 21214
0 21216 7 1 2 62039 21215
0 21217 5 1 1 21216
0 21218 7 1 2 60291 64098
0 21219 5 1 1 21218
0 21220 7 2 2 43218 56736
0 21221 7 1 2 61811 63949
0 21222 7 1 2 64563 21221
0 21223 5 1 1 21222
0 21224 7 1 2 21219 21223
0 21225 5 1 1 21224
0 21226 7 1 2 54166 21225
0 21227 5 1 1 21226
0 21228 7 1 2 21217 21227
0 21229 5 1 1 21228
0 21230 7 1 2 55368 21229
0 21231 5 1 1 21230
0 21232 7 1 2 62040 61239
0 21233 5 1 1 21232
0 21234 7 1 2 48862 61931
0 21235 7 1 2 61944 21234
0 21236 5 1 1 21235
0 21237 7 1 2 21233 21236
0 21238 5 1 1 21237
0 21239 7 1 2 40634 21238
0 21240 5 1 1 21239
0 21241 7 1 2 64121 62041
0 21242 5 1 1 21241
0 21243 7 1 2 21240 21242
0 21244 5 1 1 21243
0 21245 7 1 2 48119 21244
0 21246 5 1 1 21245
0 21247 7 1 2 61314 63623
0 21248 5 1 1 21247
0 21249 7 1 2 59002 50777
0 21250 7 1 2 60335 21249
0 21251 5 1 1 21250
0 21252 7 1 2 21248 21251
0 21253 5 1 1 21252
0 21254 7 1 2 50785 21253
0 21255 5 1 1 21254
0 21256 7 1 2 21246 21255
0 21257 5 1 1 21256
0 21258 7 1 2 49207 21257
0 21259 5 1 1 21258
0 21260 7 2 2 44213 41367
0 21261 7 1 2 58570 64565
0 21262 7 1 2 52207 21261
0 21263 5 1 1 21262
0 21264 7 1 2 5216 21263
0 21265 5 1 1 21264
0 21266 7 1 2 60292 21265
0 21267 5 1 1 21266
0 21268 7 3 2 43120 61972
0 21269 7 1 2 60383 64311
0 21270 7 1 2 64567 21269
0 21271 7 1 2 64564 21270
0 21272 5 1 1 21271
0 21273 7 1 2 21267 21272
0 21274 5 1 1 21273
0 21275 7 1 2 64014 21274
0 21276 5 1 1 21275
0 21277 7 1 2 21259 21276
0 21278 7 1 2 21231 21277
0 21279 5 1 1 21278
0 21280 7 1 2 42640 21279
0 21281 5 1 1 21280
0 21282 7 1 2 50267 64272
0 21283 5 1 1 21282
0 21284 7 1 2 40635 21283
0 21285 5 1 1 21284
0 21286 7 1 2 41672 56724
0 21287 7 1 2 61240 21286
0 21288 5 1 1 21287
0 21289 7 1 2 21285 21288
0 21290 5 1 1 21289
0 21291 7 1 2 42838 21290
0 21292 5 1 1 21291
0 21293 7 1 2 60699 63409
0 21294 5 1 1 21293
0 21295 7 1 2 21292 21294
0 21296 5 1 1 21295
0 21297 7 1 2 40866 21296
0 21298 5 1 1 21297
0 21299 7 1 2 53096 52153
0 21300 5 1 1 21299
0 21301 7 1 2 21300 63121
0 21302 5 1 1 21301
0 21303 7 1 2 41368 62383
0 21304 7 1 2 21302 21303
0 21305 5 1 1 21304
0 21306 7 1 2 21298 21305
0 21307 5 1 1 21306
0 21308 7 1 2 42994 21307
0 21309 5 1 1 21308
0 21310 7 1 2 55007 11825
0 21311 5 1 1 21310
0 21312 7 1 2 48255 62401
0 21313 7 1 2 21311 21312
0 21314 5 1 1 21313
0 21315 7 1 2 21309 21314
0 21316 5 1 1 21315
0 21317 7 1 2 53906 21316
0 21318 5 1 1 21317
0 21319 7 1 2 53067 53119
0 21320 7 1 2 64205 21319
0 21321 5 1 1 21320
0 21322 7 1 2 21318 21321
0 21323 5 1 1 21322
0 21324 7 1 2 57684 59472
0 21325 7 1 2 21323 21324
0 21326 5 1 1 21325
0 21327 7 1 2 21281 21326
0 21328 7 1 2 21213 21327
0 21329 5 1 1 21328
0 21330 7 1 2 40240 21329
0 21331 5 1 1 21330
0 21332 7 1 2 64059 64499
0 21333 5 1 1 21332
0 21334 7 1 2 61963 63892
0 21335 5 1 1 21334
0 21336 7 1 2 12549 894
0 21337 5 1 1 21336
0 21338 7 1 2 44117 16218
0 21339 7 1 2 21337 21338
0 21340 5 1 1 21339
0 21341 7 1 2 21335 21340
0 21342 5 1 1 21341
0 21343 7 1 2 42839 63604
0 21344 7 1 2 21342 21343
0 21345 5 1 1 21344
0 21346 7 1 2 21333 21345
0 21347 5 1 1 21346
0 21348 7 1 2 41673 21347
0 21349 5 1 1 21348
0 21350 7 2 2 55411 56958
0 21351 5 1 1 64570
0 21352 7 1 2 40867 57518
0 21353 5 1 1 21352
0 21354 7 1 2 21351 21353
0 21355 5 1 1 21354
0 21356 7 1 2 48695 21355
0 21357 5 1 1 21356
0 21358 7 1 2 53832 51473
0 21359 5 1 1 21358
0 21360 7 1 2 21357 21359
0 21361 5 1 1 21360
0 21362 7 1 2 57291 64076
0 21363 7 1 2 21361 21362
0 21364 5 1 1 21363
0 21365 7 1 2 21349 21364
0 21366 5 1 1 21365
0 21367 7 1 2 58984 21366
0 21368 5 1 1 21367
0 21369 7 2 2 62730 46690
0 21370 5 1 1 64572
0 21371 7 1 2 63774 64573
0 21372 7 1 2 61911 21371
0 21373 5 1 1 21372
0 21374 7 1 2 21368 21373
0 21375 5 1 1 21374
0 21376 7 1 2 45728 21375
0 21377 5 1 1 21376
0 21378 7 1 2 40419 56742
0 21379 5 1 1 21378
0 21380 7 1 2 63908 53496
0 21381 5 1 1 21380
0 21382 7 1 2 21379 21381
0 21383 5 1 1 21382
0 21384 7 1 2 63599 21383
0 21385 5 1 1 21384
0 21386 7 2 2 45729 63695
0 21387 7 1 2 64574 63700
0 21388 5 1 1 21387
0 21389 7 1 2 21385 21388
0 21390 5 1 1 21389
0 21391 7 1 2 44118 21390
0 21392 5 1 1 21391
0 21393 7 1 2 56910 57695
0 21394 7 1 2 64575 21393
0 21395 5 1 1 21394
0 21396 7 1 2 21392 21395
0 21397 5 1 1 21396
0 21398 7 1 2 48276 21397
0 21399 5 1 1 21398
0 21400 7 1 2 64152 64467
0 21401 7 1 2 63600 21400
0 21402 5 1 1 21401
0 21403 7 1 2 21399 21402
0 21404 7 1 2 21377 21403
0 21405 7 1 2 21331 21404
0 21406 5 1 1 21405
0 21407 7 1 2 58552 21406
0 21408 5 1 1 21407
0 21409 7 4 2 44308 41760
0 21410 7 1 2 63065 64576
0 21411 7 1 2 60073 21410
0 21412 7 1 2 56798 60146
0 21413 7 1 2 57163 21412
0 21414 7 1 2 21411 21413
0 21415 7 1 2 64524 21414
0 21416 5 1 1 21415
0 21417 7 1 2 21408 21416
0 21418 5 1 1 21417
0 21419 7 1 2 46754 21418
0 21420 5 1 1 21419
0 21421 7 1 2 64474 51328
0 21422 5 1 1 21421
0 21423 7 1 2 52069 58307
0 21424 5 1 1 21423
0 21425 7 1 2 21422 21424
0 21426 5 1 1 21425
0 21427 7 1 2 52154 21426
0 21428 5 1 1 21427
0 21429 7 1 2 46691 53514
0 21430 7 1 2 52070 21429
0 21431 5 1 1 21430
0 21432 7 1 2 52101 56959
0 21433 7 1 2 64082 21432
0 21434 5 1 1 21433
0 21435 7 1 2 21431 21434
0 21436 7 1 2 21428 21435
0 21437 5 1 1 21436
0 21438 7 1 2 42995 21437
0 21439 5 1 1 21438
0 21440 7 2 2 48256 57136
0 21441 5 1 1 64580
0 21442 7 1 2 64089 64581
0 21443 5 1 1 21442
0 21444 7 1 2 21439 21443
0 21445 5 1 1 21444
0 21446 7 1 2 49526 21445
0 21447 5 1 1 21446
0 21448 7 1 2 51543 50786
0 21449 5 1 1 21448
0 21450 7 1 2 57903 21449
0 21451 5 1 1 21450
0 21452 7 1 2 48696 21451
0 21453 5 1 1 21452
0 21454 7 1 2 45730 21453
0 21455 7 1 2 21447 21454
0 21456 5 1 1 21455
0 21457 7 1 2 48195 2902
0 21458 5 1 1 21457
0 21459 7 1 2 41125 21458
0 21460 5 1 1 21459
0 21461 7 1 2 19111 21460
0 21462 5 1 1 21461
0 21463 7 1 2 62530 21462
0 21464 5 1 1 21463
0 21465 7 1 2 52830 64084
0 21466 5 1 1 21465
0 21467 7 1 2 63544 21466
0 21468 5 1 1 21467
0 21469 7 1 2 42840 64055
0 21470 5 1 1 21469
0 21471 7 1 2 21468 21470
0 21472 5 1 1 21471
0 21473 7 1 2 42996 21472
0 21474 5 1 1 21473
0 21475 7 1 2 21464 21474
0 21476 5 1 1 21475
0 21477 7 1 2 40241 21476
0 21478 5 1 1 21477
0 21479 7 1 2 49527 57342
0 21480 5 1 1 21479
0 21481 7 1 2 55369 64315
0 21482 5 1 1 21481
0 21483 7 1 2 21480 21482
0 21484 5 1 1 21483
0 21485 7 1 2 49672 21484
0 21486 5 1 1 21485
0 21487 7 2 2 48584 64197
0 21488 7 1 2 64105 64582
0 21489 5 1 1 21488
0 21490 7 1 2 42386 21489
0 21491 7 1 2 21486 21490
0 21492 7 1 2 21478 21491
0 21493 5 1 1 21492
0 21494 7 1 2 53907 21493
0 21495 7 1 2 21456 21494
0 21496 5 1 1 21495
0 21497 7 3 2 52208 58188
0 21498 5 1 1 64584
0 21499 7 1 2 52641 64585
0 21500 7 1 2 64493 21499
0 21501 5 1 1 21500
0 21502 7 1 2 21496 21501
0 21503 5 1 1 21502
0 21504 7 1 2 43121 21503
0 21505 5 1 1 21504
0 21506 7 1 2 52155 62068
0 21507 5 1 1 21506
0 21508 7 1 2 58861 61427
0 21509 5 1 1 21508
0 21510 7 1 2 21507 21509
0 21511 5 1 1 21510
0 21512 7 1 2 48120 21511
0 21513 5 1 1 21512
0 21514 7 1 2 51688 64091
0 21515 5 1 1 21514
0 21516 7 1 2 21513 21515
0 21517 5 1 1 21516
0 21518 7 1 2 40061 21517
0 21519 5 1 1 21518
0 21520 7 1 2 48380 58862
0 21521 7 1 2 63860 21520
0 21522 5 1 1 21521
0 21523 7 1 2 21519 21522
0 21524 5 1 1 21523
0 21525 7 1 2 44119 21524
0 21526 5 1 1 21525
0 21527 7 2 2 50332 49775
0 21528 7 1 2 49673 64587
0 21529 5 1 1 21528
0 21530 7 2 2 44806 56181
0 21531 5 1 1 64589
0 21532 7 1 2 52414 64590
0 21533 5 1 1 21532
0 21534 7 1 2 21529 21533
0 21535 5 1 1 21534
0 21536 7 1 2 64207 21535
0 21537 5 1 1 21536
0 21538 7 1 2 21526 21537
0 21539 5 1 1 21538
0 21540 7 1 2 49528 21539
0 21541 5 1 1 21540
0 21542 7 1 2 45731 48638
0 21543 7 1 2 64240 21542
0 21544 5 1 1 21543
0 21545 7 1 2 56300 62347
0 21546 7 1 2 64583 21545
0 21547 5 1 1 21546
0 21548 7 1 2 21544 21547
0 21549 5 1 1 21548
0 21550 7 1 2 48697 21549
0 21551 5 1 1 21550
0 21552 7 1 2 47850 59662
0 21553 7 1 2 55370 61428
0 21554 7 1 2 21552 21553
0 21555 5 1 1 21554
0 21556 7 1 2 21551 21555
0 21557 7 1 2 21541 21556
0 21558 5 1 1 21557
0 21559 7 1 2 54167 21558
0 21560 5 1 1 21559
0 21561 7 1 2 21505 21560
0 21562 5 1 1 21561
0 21563 7 1 2 46631 21562
0 21564 5 1 1 21563
0 21565 7 1 2 56573 63679
0 21566 7 1 2 64497 21565
0 21567 5 1 1 21566
0 21568 7 1 2 21564 21567
0 21569 5 1 1 21568
0 21570 7 1 2 43219 21569
0 21571 5 1 1 21570
0 21572 7 1 2 64534 64491
0 21573 5 1 1 21572
0 21574 7 1 2 45943 21573
0 21575 7 1 2 21571 21574
0 21576 5 1 1 21575
0 21577 7 1 2 64203 60359
0 21578 5 1 1 21577
0 21579 7 1 2 50033 52742
0 21580 5 1 1 21579
0 21581 7 1 2 56406 21580
0 21582 5 1 1 21581
0 21583 7 1 2 40062 21582
0 21584 5 1 1 21583
0 21585 7 1 2 57587 52743
0 21586 5 1 1 21585
0 21587 7 1 2 56407 21586
0 21588 5 1 1 21587
0 21589 7 1 2 41126 21588
0 21590 5 1 1 21589
0 21591 7 1 2 21584 21590
0 21592 5 1 1 21591
0 21593 7 1 2 40242 21592
0 21594 5 1 1 21593
0 21595 7 1 2 48698 47231
0 21596 5 1 1 21595
0 21597 7 1 2 21594 21596
0 21598 5 1 1 21597
0 21599 7 1 2 60293 21598
0 21600 5 1 1 21599
0 21601 7 1 2 21578 21600
0 21602 5 1 1 21601
0 21603 7 1 2 44120 21602
0 21604 5 1 1 21603
0 21605 7 1 2 47468 63741
0 21606 5 1 1 21605
0 21607 7 1 2 40243 59473
0 21608 5 1 1 21607
0 21609 7 1 2 21606 21608
0 21610 5 1 1 21609
0 21611 7 1 2 45732 21610
0 21612 5 1 1 21611
0 21613 7 1 2 48699 61290
0 21614 5 1 1 21613
0 21615 7 1 2 21612 21614
0 21616 5 1 1 21615
0 21617 7 1 2 58881 21616
0 21618 5 1 1 21617
0 21619 7 1 2 21604 21618
0 21620 5 1 1 21619
0 21621 7 1 2 54168 21620
0 21622 5 1 1 21621
0 21623 7 1 2 44121 60532
0 21624 5 1 1 21623
0 21625 7 1 2 49347 21624
0 21626 5 1 1 21625
0 21627 7 1 2 58985 56816
0 21628 7 1 2 64444 21627
0 21629 7 1 2 21626 21628
0 21630 5 1 1 21629
0 21631 7 1 2 21622 21630
0 21632 5 1 1 21631
0 21633 7 1 2 46284 21632
0 21634 5 1 1 21633
0 21635 7 1 2 12068 61591
0 21636 5 1 1 21635
0 21637 7 1 2 40244 21636
0 21638 5 1 1 21637
0 21639 7 3 2 57264 59204
0 21640 7 2 2 47469 64591
0 21641 7 1 2 58672 64594
0 21642 5 1 1 21641
0 21643 7 1 2 62321 21642
0 21644 7 1 2 21638 21643
0 21645 5 1 1 21644
0 21646 7 1 2 45733 21645
0 21647 5 1 1 21646
0 21648 7 1 2 12586 21647
0 21649 5 1 1 21648
0 21650 7 1 2 48139 21649
0 21651 5 1 1 21650
0 21652 7 1 2 21634 21651
0 21653 5 1 1 21652
0 21654 7 1 2 43917 21653
0 21655 5 1 1 21654
0 21656 7 1 2 52102 57093
0 21657 5 1 1 21656
0 21658 7 1 2 21657 13783
0 21659 5 1 1 21658
0 21660 7 3 2 43918 45107
0 21661 7 3 2 64596 59388
0 21662 7 1 2 51645 64599
0 21663 5 1 1 21662
0 21664 7 2 2 46285 46500
0 21665 7 2 2 42841 64602
0 21666 7 4 2 43919 44268
0 21667 7 1 2 63733 64606
0 21668 7 1 2 64604 21667
0 21669 5 1 1 21668
0 21670 7 1 2 21663 21669
0 21671 5 1 1 21670
0 21672 7 1 2 21659 21671
0 21673 5 1 1 21672
0 21674 7 1 2 48191 61578
0 21675 7 1 2 64588 21674
0 21676 5 1 1 21675
0 21677 7 1 2 21673 21676
0 21678 5 1 1 21677
0 21679 7 1 2 40868 21678
0 21680 5 1 1 21679
0 21681 7 2 2 40063 58571
0 21682 7 1 2 64610 57526
0 21683 5 1 1 21682
0 21684 7 2 2 57053 52926
0 21685 5 1 1 64612
0 21686 7 1 2 21683 21685
0 21687 5 1 1 21686
0 21688 7 1 2 52103 21687
0 21689 5 1 1 21688
0 21690 7 1 2 53989 64171
0 21691 5 1 1 21690
0 21692 7 1 2 21689 21691
0 21693 5 1 1 21692
0 21694 7 1 2 56351 64600
0 21695 7 1 2 21693 21694
0 21696 5 1 1 21695
0 21697 7 1 2 21680 21696
0 21698 5 1 1 21697
0 21699 7 1 2 49529 21698
0 21700 5 1 1 21699
0 21701 7 1 2 43920 63935
0 21702 5 1 1 21701
0 21703 7 1 2 21702 61853
0 21704 5 1 1 21703
0 21705 7 1 2 52104 55371
0 21706 5 1 1 21705
0 21707 7 2 2 44957 48326
0 21708 7 1 2 41127 57137
0 21709 7 1 2 64614 21708
0 21710 5 1 1 21709
0 21711 7 1 2 21706 21710
0 21712 5 1 1 21711
0 21713 7 1 2 40064 21712
0 21714 5 1 1 21713
0 21715 7 1 2 49530 55372
0 21716 5 1 1 21715
0 21717 7 1 2 21714 21716
0 21718 5 1 1 21717
0 21719 7 1 2 46126 21718
0 21720 5 1 1 21719
0 21721 7 4 2 48222 49208
0 21722 7 1 2 49531 64616
0 21723 5 1 1 21722
0 21724 7 1 2 21720 21723
0 21725 5 1 1 21724
0 21726 7 1 2 21704 21725
0 21727 5 1 1 21726
0 21728 7 1 2 42387 64617
0 21729 7 1 2 61982 21728
0 21730 5 1 1 21729
0 21731 7 1 2 21727 21730
0 21732 7 1 2 21700 21731
0 21733 7 1 2 21655 21732
0 21734 5 1 1 21733
0 21735 7 1 2 44807 21734
0 21736 5 1 1 21735
0 21737 7 1 2 45734 48381
0 21738 5 2 1 21737
0 21739 7 1 2 64620 53028
0 21740 5 1 1 21739
0 21741 7 1 2 41505 21740
0 21742 5 1 1 21741
0 21743 7 1 2 64495 21742
0 21744 5 1 1 21743
0 21745 7 1 2 59474 21744
0 21746 5 1 1 21745
0 21747 7 4 2 40420 41506
0 21748 5 1 1 64622
0 21749 7 1 2 46501 64623
0 21750 7 1 2 63137 21749
0 21751 5 1 1 21750
0 21752 7 1 2 21746 21751
0 21753 5 1 1 21752
0 21754 7 1 2 54169 21753
0 21755 5 1 1 21754
0 21756 7 1 2 60467 57142
0 21757 7 1 2 64475 21756
0 21758 5 1 1 21757
0 21759 7 1 2 21755 21758
0 21760 5 1 1 21759
0 21761 7 1 2 40636 21760
0 21762 5 1 1 21761
0 21763 7 1 2 54655 64122
0 21764 7 1 2 61579 21763
0 21765 5 1 1 21764
0 21766 7 1 2 21762 21765
0 21767 5 1 1 21766
0 21768 7 1 2 55290 21767
0 21769 5 1 1 21768
0 21770 7 2 2 61869 64383
0 21771 7 1 2 56799 64626
0 21772 7 2 2 64551 21771
0 21773 5 1 1 64628
0 21774 7 1 2 52927 64629
0 21775 5 1 1 21774
0 21776 7 1 2 60702 19528
0 21777 5 1 1 21776
0 21778 7 1 2 40245 21777
0 21779 5 1 1 21778
0 21780 7 1 2 56408 21779
0 21781 5 1 1 21780
0 21782 7 1 2 54170 21781
0 21783 5 1 1 21782
0 21784 7 1 2 64476 64613
0 21785 5 1 1 21784
0 21786 7 1 2 61119 21785
0 21787 7 1 2 21783 21786
0 21788 5 1 1 21787
0 21789 7 1 2 60468 61925
0 21790 7 1 2 21788 21789
0 21791 5 1 1 21790
0 21792 7 1 2 21775 21791
0 21793 5 1 1 21792
0 21794 7 1 2 40869 21793
0 21795 5 1 1 21794
0 21796 7 1 2 21769 21795
0 21797 5 1 1 21796
0 21798 7 1 2 42997 21797
0 21799 5 1 1 21798
0 21800 7 1 2 57094 64210
0 21801 5 1 1 21800
0 21802 7 1 2 53644 52761
0 21803 7 1 2 64027 21802
0 21804 5 1 1 21803
0 21805 7 1 2 21801 21804
0 21806 5 1 1 21805
0 21807 7 1 2 21806 61987
0 21808 5 1 1 21807
0 21809 7 1 2 51291 62276
0 21810 7 2 2 55299 21809
0 21811 7 1 2 40065 61973
0 21812 7 1 2 64630 21811
0 21813 5 1 1 21812
0 21814 7 1 2 21808 21813
0 21815 5 1 1 21814
0 21816 7 1 2 40637 21815
0 21817 5 1 1 21816
0 21818 7 1 2 62123 62271
0 21819 7 1 2 64631 21818
0 21820 5 1 1 21819
0 21821 7 1 2 21817 21820
0 21822 5 1 1 21821
0 21823 7 1 2 52105 21822
0 21824 5 1 1 21823
0 21825 7 1 2 56379 61988
0 21826 5 1 1 21825
0 21827 7 2 2 48512 48639
0 21828 5 1 1 64632
0 21829 7 1 2 55680 55966
0 21830 5 1 1 21829
0 21831 7 1 2 21828 21830
0 21832 5 1 1 21831
0 21833 7 1 2 59475 21832
0 21834 5 1 1 21833
0 21835 7 1 2 21826 21834
0 21836 5 1 1 21835
0 21837 7 1 2 54171 21836
0 21838 5 1 1 21837
0 21839 7 1 2 55432 59476
0 21840 7 1 2 54885 21839
0 21841 5 1 1 21840
0 21842 7 1 2 21838 21841
0 21843 5 1 1 21842
0 21844 7 1 2 64211 21843
0 21845 5 1 1 21844
0 21846 7 2 2 57127 54553
0 21847 5 1 1 64634
0 21848 7 2 2 52866 58189
0 21849 5 1 1 64636
0 21850 7 1 2 46412 64637
0 21851 5 1 1 21850
0 21852 7 1 2 21847 21851
0 21853 5 2 1 21852
0 21854 7 1 2 51689 55964
0 21855 7 1 2 64638 21854
0 21856 5 1 1 21855
0 21857 7 1 2 54028 2866
0 21858 5 1 1 21857
0 21859 7 1 2 41674 57444
0 21860 7 1 2 21858 21859
0 21861 5 1 1 21860
0 21862 7 1 2 21856 21861
0 21863 5 1 1 21862
0 21864 7 1 2 59477 21863
0 21865 5 1 1 21864
0 21866 7 1 2 10435 62315
0 21867 5 1 1 21866
0 21868 7 1 2 62973 56582
0 21869 7 1 2 61939 21868
0 21870 7 1 2 21867 21869
0 21871 5 1 1 21870
0 21872 7 1 2 21865 21871
0 21873 5 1 1 21872
0 21874 7 1 2 42842 21873
0 21875 5 1 1 21874
0 21876 7 1 2 21845 21875
0 21877 7 1 2 21824 21876
0 21878 5 1 1 21877
0 21879 7 1 2 49532 21878
0 21880 5 1 1 21879
0 21881 7 1 2 52106 55308
0 21882 5 1 1 21881
0 21883 7 1 2 21882 21441
0 21884 5 1 1 21883
0 21885 7 1 2 60294 21884
0 21886 5 1 1 21885
0 21887 7 1 2 42998 60027
0 21888 7 1 2 63189 21887
0 21889 5 1 1 21888
0 21890 7 1 2 21886 21889
0 21891 5 1 1 21890
0 21892 7 1 2 48513 21891
0 21893 5 1 1 21892
0 21894 7 1 2 64212 63742
0 21895 5 1 1 21894
0 21896 7 2 2 46809 55291
0 21897 5 1 1 64640
0 21898 7 1 2 41128 64169
0 21899 5 1 1 21898
0 21900 7 1 2 3651 21899
0 21901 5 1 1 21900
0 21902 7 1 2 40870 21901
0 21903 5 1 1 21902
0 21904 7 1 2 21897 21903
0 21905 5 1 1 21904
0 21906 7 1 2 42999 61291
0 21907 7 1 2 21905 21906
0 21908 5 1 1 21907
0 21909 7 1 2 21895 21908
0 21910 5 1 1 21909
0 21911 7 1 2 62555 21910
0 21912 5 1 1 21911
0 21913 7 1 2 21893 21912
0 21914 5 1 1 21913
0 21915 7 1 2 45735 21914
0 21916 5 1 1 21915
0 21917 7 6 2 41808 62763
0 21918 7 1 2 60022 64642
0 21919 7 1 2 57853 62590
0 21920 7 1 2 21918 21919
0 21921 5 1 1 21920
0 21922 7 1 2 21916 21921
0 21923 5 1 1 21922
0 21924 7 1 2 57095 21923
0 21925 5 1 1 21924
0 21926 7 1 2 60478 12713
0 21927 5 1 1 21926
0 21928 7 1 2 61992 21927
0 21929 5 1 1 21928
0 21930 7 1 2 62322 21929
0 21931 5 1 1 21930
0 21932 7 1 2 61926 21931
0 21933 5 1 1 21932
0 21934 7 1 2 61878 62272
0 21935 7 1 2 64595 21934
0 21936 5 1 1 21935
0 21937 7 1 2 21933 21936
0 21938 5 1 1 21937
0 21939 7 1 2 45736 21938
0 21940 5 1 1 21939
0 21941 7 1 2 21773 21940
0 21942 5 1 1 21941
0 21943 7 1 2 57337 21942
0 21944 5 1 1 21943
0 21945 7 1 2 42641 21944
0 21946 7 1 2 21925 21945
0 21947 7 1 2 21880 21946
0 21948 7 1 2 21799 21947
0 21949 7 1 2 21736 21948
0 21950 5 1 1 21949
0 21951 7 1 2 58553 21950
0 21952 7 1 2 21576 21951
0 21953 5 1 1 21952
0 21954 7 3 2 45149 45310
0 21955 7 2 2 41809 64648
0 21956 7 1 2 53331 64651
0 21957 7 1 2 64526 21956
0 21958 7 5 2 41024 44309
0 21959 7 2 2 40961 64653
0 21960 7 1 2 50034 64658
0 21961 7 1 2 64043 21960
0 21962 7 1 2 21957 21961
0 21963 5 1 1 21962
0 21964 7 1 2 21953 21963
0 21965 7 1 2 21420 21964
0 21966 7 1 2 21028 21965
0 21967 7 1 2 20697 21966
0 21968 7 1 2 19615 21967
0 21969 5 1 1 21968
0 21970 7 1 2 47119 21969
0 21971 5 1 1 21970
0 21972 7 36 2 44310 45150
0 21973 5 1 1 64660
0 21974 7 4 2 53908 64661
0 21975 7 1 2 60074 63128
0 21976 7 1 2 64696 21975
0 21977 7 1 2 55499 61957
0 21978 7 1 2 21976 21977
0 21979 7 1 2 64522 21978
0 21980 5 1 1 21979
0 21981 7 4 2 46413 62735
0 21982 7 1 2 40066 64700
0 21983 5 1 1 21982
0 21984 7 1 2 61850 21983
0 21985 5 1 1 21984
0 21986 7 1 2 56989 21985
0 21987 5 1 1 21986
0 21988 7 1 2 64312 62556
0 21989 7 1 2 64701 21988
0 21990 5 1 1 21989
0 21991 7 1 2 21987 21990
0 21992 5 1 1 21991
0 21993 7 1 2 42642 21992
0 21994 5 1 1 21993
0 21995 7 2 2 42843 64702
0 21996 7 1 2 50974 64110
0 21997 7 1 2 64704 21996
0 21998 5 1 1 21997
0 21999 7 1 2 21994 21998
0 22000 5 1 1 21999
0 22001 7 1 2 44958 22000
0 22002 5 1 1 22001
0 22003 7 1 2 51977 57696
0 22004 7 1 2 64705 22003
0 22005 5 1 1 22004
0 22006 7 1 2 22002 22005
0 22007 5 1 1 22006
0 22008 7 1 2 44122 22007
0 22009 5 1 1 22008
0 22010 7 1 2 57554 19266
0 22011 5 1 1 22010
0 22012 7 1 2 40871 22011
0 22013 5 1 1 22012
0 22014 7 1 2 55292 63893
0 22015 5 1 1 22014
0 22016 7 1 2 22013 22015
0 22017 7 1 2 64142 22016
0 22018 5 1 1 22017
0 22019 7 1 2 63548 22018
0 22020 5 1 1 22019
0 22021 7 1 2 49209 63894
0 22022 5 1 1 22021
0 22023 7 1 2 64458 22022
0 22024 5 1 1 22023
0 22025 7 1 2 46127 22024
0 22026 5 1 1 22025
0 22027 7 1 2 55277 63885
0 22028 5 1 1 22027
0 22029 7 1 2 22026 22028
0 22030 5 1 1 22029
0 22031 7 1 2 58417 22030
0 22032 5 1 1 22031
0 22033 7 1 2 22020 22032
0 22034 5 1 1 22033
0 22035 7 1 2 49033 22034
0 22036 5 1 1 22035
0 22037 7 1 2 44959 63866
0 22038 5 1 1 22037
0 22039 7 1 2 22038 10314
0 22040 5 1 1 22039
0 22041 7 1 2 55069 22040
0 22042 5 1 1 22041
0 22043 7 2 2 44960 63864
0 22044 5 1 1 64706
0 22045 7 1 2 46128 59033
0 22046 7 1 2 61542 22045
0 22047 7 1 2 62639 22046
0 22048 5 1 1 22047
0 22049 7 1 2 22044 22048
0 22050 7 1 2 22042 22049
0 22051 5 1 1 22050
0 22052 7 1 2 56830 22051
0 22053 5 1 1 22052
0 22054 7 1 2 41025 53497
0 22055 7 2 2 56689 22054
0 22056 7 2 2 41675 59205
0 22057 7 1 2 64710 63904
0 22058 7 1 2 64708 22057
0 22059 5 1 1 22058
0 22060 7 2 2 56681 52232
0 22061 5 1 1 64712
0 22062 7 2 2 45944 55070
0 22063 7 1 2 64713 64714
0 22064 7 1 2 63532 22063
0 22065 5 1 1 22064
0 22066 7 1 2 22059 22065
0 22067 7 1 2 22053 22066
0 22068 5 1 1 22067
0 22069 7 1 2 40872 22068
0 22070 5 1 1 22069
0 22071 7 1 2 22036 22070
0 22072 7 1 2 22009 22071
0 22073 5 1 1 22072
0 22074 7 1 2 50518 22073
0 22075 5 1 1 22074
0 22076 7 2 2 53909 55345
0 22077 5 1 1 64716
0 22078 7 1 2 22077 18361
0 22079 5 1 1 22078
0 22080 7 1 2 49210 22079
0 22081 5 1 1 22080
0 22082 7 1 2 55181 55757
0 22083 5 1 1 22082
0 22084 7 1 2 53214 55164
0 22085 5 1 1 22084
0 22086 7 1 2 22083 22085
0 22087 5 1 1 22086
0 22088 7 1 2 48700 22087
0 22089 5 1 1 22088
0 22090 7 1 2 22081 22089
0 22091 5 1 1 22090
0 22092 7 1 2 56076 58418
0 22093 7 1 2 22091 22092
0 22094 5 1 1 22093
0 22095 7 1 2 22075 22094
0 22096 5 1 1 22095
0 22097 7 1 2 43220 22096
0 22098 5 1 1 22097
0 22099 7 2 2 58659 59507
0 22100 7 1 2 61139 64718
0 22101 5 1 1 22100
0 22102 7 3 2 49533 62351
0 22103 7 1 2 63589 63190
0 22104 7 1 2 64720 22103
0 22105 5 1 1 22104
0 22106 7 1 2 22101 22105
0 22107 5 1 1 22106
0 22108 7 1 2 40873 22107
0 22109 5 1 1 22108
0 22110 7 1 2 49732 53264
0 22111 7 1 2 64719 22110
0 22112 5 1 1 22111
0 22113 7 1 2 22109 22112
0 22114 5 1 1 22113
0 22115 7 1 2 44961 22114
0 22116 5 1 1 22115
0 22117 7 1 2 63590 60075
0 22118 7 1 2 61338 22117
0 22119 7 1 2 60679 22118
0 22120 7 1 2 56109 22119
0 22121 5 1 1 22120
0 22122 7 1 2 22116 22121
0 22123 5 1 1 22122
0 22124 7 1 2 44269 22123
0 22125 5 1 1 22124
0 22126 7 1 2 59218 55300
0 22127 5 1 1 22126
0 22128 7 1 2 63950 58600
0 22129 5 1 1 22128
0 22130 7 1 2 22127 22129
0 22131 5 1 1 22130
0 22132 7 1 2 40067 62079
0 22133 7 1 2 64721 22132
0 22134 7 1 2 22131 22133
0 22135 5 1 1 22134
0 22136 7 1 2 22125 22135
0 22137 5 1 1 22136
0 22138 7 1 2 44214 22137
0 22139 5 1 1 22138
0 22140 7 2 2 45057 55301
0 22141 5 1 1 64723
0 22142 7 1 2 42844 57461
0 22143 5 1 1 22142
0 22144 7 1 2 22141 22143
0 22145 5 1 1 22144
0 22146 7 1 2 62124 62926
0 22147 7 1 2 64722 22146
0 22148 7 1 2 22145 22147
0 22149 5 1 1 22148
0 22150 7 1 2 22139 22149
0 22151 5 1 1 22150
0 22152 7 1 2 45945 22151
0 22153 5 1 1 22152
0 22154 7 1 2 47991 64601
0 22155 5 1 1 22154
0 22156 7 1 2 62535 60469
0 22157 5 1 1 22156
0 22158 7 1 2 22155 22157
0 22159 5 1 1 22158
0 22160 7 1 2 48916 22159
0 22161 5 1 1 22160
0 22162 7 1 2 62536 62931
0 22163 5 1 1 22162
0 22164 7 1 2 22161 22163
0 22165 5 1 1 22164
0 22166 7 1 2 51544 22165
0 22167 5 1 1 22166
0 22168 7 2 2 55071 56769
0 22169 7 2 2 43221 49034
0 22170 7 1 2 64727 54222
0 22171 7 1 2 64725 22170
0 22172 5 1 1 22171
0 22173 7 1 2 22167 22172
0 22174 5 1 1 22173
0 22175 7 1 2 40421 22174
0 22176 5 1 1 22175
0 22177 7 1 2 55072 55192
0 22178 5 1 1 22177
0 22179 7 2 2 48917 59410
0 22180 5 1 1 64729
0 22181 7 1 2 22178 22180
0 22182 5 1 1 22181
0 22183 7 2 2 43222 22182
0 22184 7 3 2 41369 42140
0 22185 5 1 1 64733
0 22186 7 1 2 40068 64734
0 22187 7 1 2 64731 22186
0 22188 5 1 1 22187
0 22189 7 1 2 22176 22188
0 22190 5 1 1 22189
0 22191 7 1 2 46129 22190
0 22192 5 1 1 22191
0 22193 7 5 2 43223 62736
0 22194 7 1 2 62537 49211
0 22195 7 1 2 53056 22194
0 22196 7 1 2 64736 22195
0 22197 5 1 1 22196
0 22198 7 1 2 22192 22197
0 22199 5 1 1 22198
0 22200 7 1 2 54272 22199
0 22201 5 1 1 22200
0 22202 7 1 2 22153 22201
0 22203 5 1 1 22202
0 22204 7 1 2 46414 22203
0 22205 5 1 1 22204
0 22206 7 1 2 52689 50642
0 22207 5 1 1 22206
0 22208 7 1 2 53051 22207
0 22209 5 1 1 22208
0 22210 7 1 2 40962 22209
0 22211 5 1 1 22210
0 22212 7 1 2 52690 56461
0 22213 5 1 1 22212
0 22214 7 1 2 22211 22213
0 22215 5 1 1 22214
0 22216 7 1 2 22215 62291
0 22217 5 1 1 22216
0 22218 7 1 2 57930 63874
0 22219 5 1 1 22218
0 22220 7 1 2 54273 56061
0 22221 5 1 1 22220
0 22222 7 1 2 22219 22221
0 22223 5 1 1 22222
0 22224 7 1 2 60556 22223
0 22225 5 1 1 22224
0 22226 7 1 2 22217 22225
0 22227 5 1 1 22226
0 22228 7 1 2 49534 22227
0 22229 5 1 1 22228
0 22230 7 1 2 44962 63229
0 22231 5 1 1 22230
0 22232 7 1 2 42643 49166
0 22233 5 1 1 22232
0 22234 7 1 2 22231 22233
0 22235 5 1 1 22234
0 22236 7 1 2 44808 22235
0 22237 5 1 1 22236
0 22238 7 1 2 51545 60962
0 22239 5 1 1 22238
0 22240 7 1 2 22237 22239
0 22241 5 1 1 22240
0 22242 7 1 2 53910 22241
0 22243 5 1 1 22242
0 22244 7 1 2 45946 2808
0 22245 7 1 2 64199 22244
0 22246 5 1 1 22245
0 22247 7 1 2 22243 22246
0 22248 5 1 1 22247
0 22249 7 1 2 41232 48950
0 22250 7 1 2 51334 22249
0 22251 7 1 2 22248 22250
0 22252 5 1 1 22251
0 22253 7 1 2 22229 22252
0 22254 5 1 1 22253
0 22255 7 1 2 60403 62879
0 22256 7 1 2 22254 22255
0 22257 5 1 1 22256
0 22258 7 2 2 58660 56483
0 22259 7 1 2 55454 63928
0 22260 7 1 2 64741 22259
0 22261 7 1 2 60557 22260
0 22262 5 1 1 22261
0 22263 7 1 2 22257 22262
0 22264 7 1 2 22205 22263
0 22265 5 1 1 22264
0 22266 7 1 2 42388 22265
0 22267 5 1 1 22266
0 22268 7 1 2 44270 56831
0 22269 5 1 1 22268
0 22270 7 1 2 14754 22269
0 22271 5 1 1 22270
0 22272 7 1 2 55500 54522
0 22273 5 1 1 22272
0 22274 7 1 2 57564 22273
0 22275 5 1 1 22274
0 22276 7 1 2 49035 52928
0 22277 7 1 2 22275 22276
0 22278 5 2 1 22277
0 22279 7 1 2 42644 61842
0 22280 5 1 1 22279
0 22281 7 1 2 53223 22280
0 22282 5 1 1 22281
0 22283 7 1 2 57016 52600
0 22284 7 1 2 22282 22283
0 22285 5 1 1 22284
0 22286 7 1 2 64743 22285
0 22287 5 1 1 22286
0 22288 7 1 2 22271 22287
0 22289 5 1 1 22288
0 22290 7 1 2 64061 64038
0 22291 7 1 2 53490 61826
0 22292 7 1 2 22290 22291
0 22293 5 1 1 22292
0 22294 7 1 2 22289 22293
0 22295 5 1 1 22294
0 22296 7 1 2 41810 22295
0 22297 5 1 1 22296
0 22298 7 1 2 53292 56911
0 22299 5 1 1 22298
0 22300 7 1 2 17808 22299
0 22301 5 1 1 22300
0 22302 7 1 2 56832 22301
0 22303 5 1 1 22302
0 22304 7 3 2 45947 51488
0 22305 7 1 2 64568 64745
0 22306 5 1 1 22305
0 22307 7 1 2 22303 22306
0 22308 5 1 1 22307
0 22309 7 1 2 40638 22308
0 22310 5 1 1 22309
0 22311 7 1 2 46415 63840
0 22312 7 1 2 59120 22311
0 22313 7 1 2 54358 22312
0 22314 5 1 1 22313
0 22315 7 1 2 22310 22314
0 22316 5 1 1 22315
0 22317 7 1 2 55501 22316
0 22318 5 1 1 22317
0 22319 7 1 2 56833 58673
0 22320 7 1 2 64192 22319
0 22321 5 1 1 22320
0 22322 7 1 2 22318 22321
0 22323 5 1 1 22322
0 22324 7 1 2 7191 1899
0 22325 5 1 1 22324
0 22326 7 1 2 16019 22325
0 22327 7 1 2 22323 22326
0 22328 5 1 1 22327
0 22329 7 1 2 40963 53253
0 22330 7 2 2 64148 22329
0 22331 7 1 2 53304 55512
0 22332 7 1 2 64748 22331
0 22333 5 1 1 22332
0 22334 7 1 2 64744 22333
0 22335 5 1 1 22334
0 22336 7 1 2 41026 62139
0 22337 7 1 2 22335 22336
0 22338 5 1 1 22337
0 22339 7 2 2 53293 49116
0 22340 5 1 1 64750
0 22341 7 1 2 7776 22340
0 22342 5 1 1 22341
0 22343 7 1 2 40639 22342
0 22344 5 1 1 22343
0 22345 7 1 2 54359 55174
0 22346 5 1 1 22345
0 22347 7 1 2 22344 22346
0 22348 5 1 1 22347
0 22349 7 1 2 55502 22348
0 22350 5 1 1 22349
0 22351 7 1 2 63285 55175
0 22352 5 1 1 22351
0 22353 7 1 2 22350 22352
0 22354 5 1 1 22353
0 22355 7 1 2 56160 63552
0 22356 7 1 2 22354 22355
0 22357 5 1 1 22356
0 22358 7 1 2 22338 22357
0 22359 7 1 2 22328 22358
0 22360 7 1 2 22297 22359
0 22361 5 1 1 22360
0 22362 7 1 2 43224 22361
0 22363 5 1 1 22362
0 22364 7 1 2 53833 63402
0 22365 7 1 2 63706 22364
0 22366 7 1 2 60765 61333
0 22367 7 1 2 22365 22366
0 22368 5 1 1 22367
0 22369 7 1 2 22363 22368
0 22370 5 1 1 22369
0 22371 7 1 2 49535 22370
0 22372 5 1 1 22371
0 22373 7 3 2 53305 61832
0 22374 7 2 2 55776 50148
0 22375 7 1 2 64752 64755
0 22376 7 2 2 55244 52962
0 22377 7 1 2 64757 63929
0 22378 7 1 2 22375 22377
0 22379 5 1 1 22378
0 22380 7 1 2 46286 22379
0 22381 7 1 2 22372 22380
0 22382 7 1 2 22267 22381
0 22383 7 1 2 22098 22382
0 22384 5 1 1 22383
0 22385 7 1 2 57283 63070
0 22386 7 1 2 63132 22385
0 22387 5 1 1 22386
0 22388 7 1 2 57208 62287
0 22389 7 1 2 58340 22388
0 22390 5 1 1 22389
0 22391 7 1 2 22387 22390
0 22392 5 1 1 22391
0 22393 7 1 2 56646 22392
0 22394 5 1 1 22393
0 22395 7 1 2 60578 63251
0 22396 7 1 2 63054 22395
0 22397 5 1 1 22396
0 22398 7 1 2 22394 22397
0 22399 5 1 1 22398
0 22400 7 1 2 55073 22399
0 22401 5 1 1 22400
0 22402 7 2 2 44809 57856
0 22403 7 2 2 55820 55608
0 22404 7 1 2 64759 64761
0 22405 5 1 1 22404
0 22406 7 1 2 56690 60810
0 22407 7 1 2 50495 22406
0 22408 5 1 1 22407
0 22409 7 1 2 22405 22408
0 22410 5 1 1 22409
0 22411 7 1 2 40874 22410
0 22412 5 1 1 22411
0 22413 7 1 2 50265 63225
0 22414 5 1 1 22413
0 22415 7 1 2 52577 53200
0 22416 5 1 1 22415
0 22417 7 1 2 49674 22416
0 22418 5 1 1 22417
0 22419 7 1 2 53236 52963
0 22420 7 1 2 53366 22419
0 22421 5 1 1 22420
0 22422 7 1 2 63291 22421
0 22423 7 1 2 22418 22422
0 22424 5 1 1 22423
0 22425 7 1 2 44963 22424
0 22426 5 1 1 22425
0 22427 7 1 2 22414 22426
0 22428 5 1 1 22427
0 22429 7 1 2 42845 58685
0 22430 7 1 2 22428 22429
0 22431 5 1 1 22430
0 22432 7 1 2 22412 22431
0 22433 5 1 1 22432
0 22434 7 1 2 59478 22433
0 22435 5 1 1 22434
0 22436 7 1 2 22401 22435
0 22437 5 1 1 22436
0 22438 7 1 2 49536 22437
0 22439 5 1 1 22438
0 22440 7 2 2 55821 46632
0 22441 7 1 2 51546 64763
0 22442 5 1 1 22441
0 22443 7 1 2 53294 49093
0 22444 7 1 2 64726 22443
0 22445 5 1 1 22444
0 22446 7 1 2 22442 22445
0 22447 5 1 1 22446
0 22448 7 1 2 40640 22447
0 22449 5 1 1 22448
0 22450 7 1 2 59411 55401
0 22451 5 1 1 22450
0 22452 7 1 2 22449 22451
0 22453 5 1 1 22452
0 22454 7 1 2 48701 22453
0 22455 5 1 1 22454
0 22456 7 1 2 57547 64764
0 22457 5 1 1 22456
0 22458 7 1 2 22455 22457
0 22459 5 1 1 22458
0 22460 7 1 2 50519 22459
0 22461 5 1 1 22460
0 22462 7 1 2 56611 59273
0 22463 7 1 2 58826 22462
0 22464 7 1 2 63261 22463
0 22465 5 1 1 22464
0 22466 7 1 2 22461 22465
0 22467 5 1 1 22466
0 22468 7 1 2 46416 22467
0 22469 5 1 1 22468
0 22470 7 1 2 41811 50798
0 22471 7 1 2 53485 22470
0 22472 7 1 2 64709 22471
0 22473 5 1 1 22472
0 22474 7 1 2 22469 22473
0 22475 5 1 1 22474
0 22476 7 1 2 43225 22475
0 22477 5 1 1 22476
0 22478 7 1 2 22439 22477
0 22479 5 1 1 22478
0 22480 7 1 2 49036 22479
0 22481 5 1 1 22480
0 22482 7 2 2 56502 62402
0 22483 5 1 1 64765
0 22484 7 3 2 54746 58280
0 22485 7 1 2 51329 64767
0 22486 5 1 1 22485
0 22487 7 1 2 22483 22486
0 22488 5 1 1 22487
0 22489 7 1 2 52156 22488
0 22490 5 1 1 22489
0 22491 7 1 2 53515 64077
0 22492 7 1 2 56503 22491
0 22493 5 1 1 22492
0 22494 7 2 2 44123 63119
0 22495 5 1 1 64770
0 22496 7 1 2 64771 64768
0 22497 5 1 1 22496
0 22498 7 1 2 22493 22497
0 22499 7 1 2 22490 22498
0 22500 5 1 1 22499
0 22501 7 1 2 54172 22500
0 22502 5 1 1 22501
0 22503 7 1 2 55006 58616
0 22504 5 1 1 22503
0 22505 7 1 2 56875 64517
0 22506 7 1 2 52157 22505
0 22507 5 1 1 22506
0 22508 7 1 2 22504 22507
0 22509 7 1 2 22502 22508
0 22510 5 1 1 22509
0 22511 7 1 2 47020 22510
0 22512 5 1 1 22511
0 22513 7 2 2 54173 47232
0 22514 7 1 2 56960 54112
0 22515 7 1 2 64772 22514
0 22516 5 1 1 22515
0 22517 7 1 2 48702 49117
0 22518 7 1 2 64009 22517
0 22519 7 1 2 52158 22518
0 22520 5 1 1 22519
0 22521 7 1 2 22516 22520
0 22522 7 1 2 22512 22521
0 22523 5 1 1 22522
0 22524 7 1 2 45948 22523
0 22525 5 1 1 22524
0 22526 7 1 2 53097 55001
0 22527 7 1 2 64397 22526
0 22528 5 1 1 22527
0 22529 7 1 2 40069 58427
0 22530 5 1 1 22529
0 22531 7 1 2 55280 22530
0 22532 5 2 1 22531
0 22533 7 1 2 48514 50357
0 22534 7 1 2 64774 22533
0 22535 5 1 1 22534
0 22536 7 1 2 22528 22535
0 22537 5 1 1 22536
0 22538 7 2 2 42645 22537
0 22539 5 1 1 64776
0 22540 7 1 2 54174 64777
0 22541 5 1 1 22540
0 22542 7 1 2 58583 64586
0 22543 5 2 1 22542
0 22544 7 1 2 40422 64405
0 22545 5 1 1 22544
0 22546 7 1 2 63292 22545
0 22547 5 2 1 22546
0 22548 7 1 2 57086 64780
0 22549 5 1 1 22548
0 22550 7 1 2 63693 60945
0 22551 5 1 1 22550
0 22552 7 1 2 22549 22551
0 22553 5 1 1 22552
0 22554 7 1 2 49212 22553
0 22555 5 1 1 22554
0 22556 7 1 2 56380 50539
0 22557 7 1 2 57365 22556
0 22558 7 1 2 57096 22557
0 22559 5 1 1 22558
0 22560 7 1 2 22555 22559
0 22561 5 1 1 22560
0 22562 7 1 2 46130 22561
0 22563 5 1 1 22562
0 22564 7 1 2 64778 22563
0 22565 5 1 1 22564
0 22566 7 1 2 47992 22565
0 22567 5 1 1 22566
0 22568 7 1 2 22541 22567
0 22569 7 1 2 22525 22568
0 22570 5 1 1 22569
0 22571 7 1 2 59479 22570
0 22572 5 1 1 22571
0 22573 7 1 2 53197 64775
0 22574 5 1 1 22573
0 22575 7 1 2 55616 59414
0 22576 5 1 1 22575
0 22577 7 1 2 22574 22576
0 22578 5 2 1 22577
0 22579 7 1 2 61671 64782
0 22580 5 1 1 22579
0 22581 7 1 2 60579 62230
0 22582 7 1 2 56745 22581
0 22583 7 1 2 58134 22582
0 22584 5 1 1 22583
0 22585 7 1 2 22580 22584
0 22586 5 1 1 22585
0 22587 7 1 2 49537 22586
0 22588 5 1 1 22587
0 22589 7 1 2 53367 55293
0 22590 5 1 1 22589
0 22591 7 1 2 40875 50520
0 22592 7 1 2 60533 22591
0 22593 5 1 1 22592
0 22594 7 1 2 22590 22593
0 22595 5 1 1 22594
0 22596 7 2 2 62345 22595
0 22597 7 6 2 41761 61777
0 22598 7 1 2 40423 64786
0 22599 7 1 2 64784 22598
0 22600 5 1 1 22599
0 22601 7 1 2 22588 22600
0 22602 5 1 1 22601
0 22603 7 1 2 49675 22602
0 22604 5 1 1 22603
0 22605 7 1 2 51330 52159
0 22606 5 1 1 22605
0 22607 7 1 2 22606 22495
0 22608 5 1 1 22607
0 22609 7 1 2 47021 64769
0 22610 5 1 1 22609
0 22611 7 1 2 54127 22610
0 22612 5 1 1 22611
0 22613 7 1 2 22608 22612
0 22614 5 1 1 22613
0 22615 7 1 2 47022 52160
0 22616 7 1 2 64766 22615
0 22617 5 1 1 22616
0 22618 7 1 2 60771 53516
0 22619 7 1 2 60550 22618
0 22620 5 1 1 22619
0 22621 7 1 2 22617 22620
0 22622 7 1 2 22614 22621
0 22623 5 1 1 22622
0 22624 7 1 2 45949 22623
0 22625 5 1 1 22624
0 22626 7 1 2 49213 64781
0 22627 5 1 1 22626
0 22628 7 1 2 64454 63671
0 22629 5 1 1 22628
0 22630 7 1 2 22627 22629
0 22631 5 1 1 22630
0 22632 7 1 2 53098 22631
0 22633 5 1 1 22632
0 22634 7 1 2 19860 22633
0 22635 5 1 1 22634
0 22636 7 1 2 47993 22635
0 22637 5 1 1 22636
0 22638 7 1 2 22539 22637
0 22639 7 1 2 22625 22638
0 22640 5 1 1 22639
0 22641 7 1 2 61672 22640
0 22642 5 1 1 22641
0 22643 7 1 2 22604 22642
0 22644 5 1 1 22643
0 22645 7 1 2 55074 22644
0 22646 5 1 1 22645
0 22647 7 1 2 61580 64783
0 22648 5 1 1 22647
0 22649 7 1 2 53557 59508
0 22650 7 1 2 59219 22649
0 22651 7 2 2 57032 60342
0 22652 7 1 2 64792 54234
0 22653 7 1 2 22650 22652
0 22654 5 1 1 22653
0 22655 7 1 2 22648 22654
0 22656 5 1 1 22655
0 22657 7 1 2 49538 22656
0 22658 5 1 1 22657
0 22659 7 1 2 48703 62731
0 22660 7 1 2 64785 22659
0 22661 5 1 1 22660
0 22662 7 1 2 22658 22661
0 22663 5 1 1 22662
0 22664 7 1 2 49676 22663
0 22665 5 1 1 22664
0 22666 7 1 2 43000 22665
0 22667 7 1 2 22646 22666
0 22668 7 1 2 22572 22667
0 22669 7 1 2 22481 22668
0 22670 5 1 1 22669
0 22671 7 1 2 58554 22670
0 22672 7 1 2 22384 22671
0 22673 5 1 1 22672
0 22674 7 1 2 21980 22673
0 22675 5 1 1 22674
0 22676 7 1 2 52107 22675
0 22677 5 1 1 22676
0 22678 7 1 2 21971 22677
0 22679 7 1 2 19015 22678
0 22680 7 1 2 17444 22679
0 22681 7 1 2 9734 22680
0 22682 7 1 2 6253 22681
0 22683 5 1 1 22682
0 22684 7 1 2 43280 22683
0 22685 5 1 1 22684
0 22686 7 1 2 53581 62352
0 22687 5 1 1 22686
0 22688 7 1 2 45950 63246
0 22689 5 1 1 22688
0 22690 7 1 2 22687 22689
0 22691 5 1 1 22690
0 22692 7 1 2 47470 22691
0 22693 5 1 1 22692
0 22694 7 1 2 52180 57437
0 22695 5 1 1 22694
0 22696 7 3 2 41965 55744
0 22697 5 1 1 64794
0 22698 7 1 2 22695 22697
0 22699 5 1 1 22698
0 22700 7 1 2 47280 22699
0 22701 5 1 1 22700
0 22702 7 1 2 22693 22701
0 22703 5 1 1 22702
0 22704 7 1 2 41233 22703
0 22705 5 1 1 22704
0 22706 7 1 2 55578 64795
0 22707 5 1 1 22706
0 22708 7 1 2 22705 22707
0 22709 5 1 1 22708
0 22710 7 1 2 40246 22709
0 22711 5 1 1 22710
0 22712 7 1 2 49677 59790
0 22713 5 1 1 22712
0 22714 7 1 2 15948 22713
0 22715 5 1 1 22714
0 22716 7 1 2 42646 22715
0 22717 5 1 1 22716
0 22718 7 1 2 22711 22717
0 22719 5 1 1 22718
0 22720 7 1 2 40424 22719
0 22721 5 1 1 22720
0 22722 7 1 2 56244 58113
0 22723 5 1 1 22722
0 22724 7 1 2 63286 22723
0 22725 5 1 1 22724
0 22726 7 1 2 22721 22725
0 22727 5 1 1 22726
0 22728 7 1 2 41370 22727
0 22729 5 1 1 22728
0 22730 7 1 2 47938 47160
0 22731 5 1 1 22730
0 22732 7 1 2 43384 22731
0 22733 5 1 1 22732
0 22734 7 1 2 48423 4126
0 22735 7 1 2 22733 22734
0 22736 5 1 1 22735
0 22737 7 1 2 44664 50236
0 22738 5 1 1 22737
0 22739 7 1 2 40070 22738
0 22740 5 1 1 22739
0 22741 7 1 2 55978 22740
0 22742 5 1 1 22741
0 22743 7 1 2 40247 22742
0 22744 5 1 1 22743
0 22745 7 1 2 45951 22744
0 22746 7 1 2 22736 22745
0 22747 5 2 1 22746
0 22748 7 1 2 50204 59781
0 22749 5 3 1 22748
0 22750 7 2 2 46942 58286
0 22751 5 1 1 64802
0 22752 7 1 2 22751 61077
0 22753 5 1 1 22752
0 22754 7 1 2 47787 22753
0 22755 5 1 1 22754
0 22756 7 1 2 64799 22755
0 22757 5 1 1 22756
0 22758 7 1 2 42647 22757
0 22759 5 1 1 22758
0 22760 7 1 2 64797 22759
0 22761 5 1 1 22760
0 22762 7 1 2 48515 22761
0 22763 5 1 1 22762
0 22764 7 1 2 22729 22763
0 22765 5 1 1 22764
0 22766 7 1 2 45737 22765
0 22767 5 1 1 22766
0 22768 7 1 2 44665 52181
0 22769 5 2 1 22768
0 22770 7 1 2 61010 58222
0 22771 5 1 1 22770
0 22772 7 1 2 42648 22771
0 22773 5 1 1 22772
0 22774 7 1 2 64804 22773
0 22775 5 1 1 22774
0 22776 7 1 2 47471 22775
0 22777 5 1 1 22776
0 22778 7 1 2 53237 63183
0 22779 5 1 1 22778
0 22780 7 1 2 22777 22779
0 22781 5 1 1 22780
0 22782 7 1 2 45311 22781
0 22783 5 1 1 22782
0 22784 7 1 2 56206 62564
0 22785 5 1 1 22784
0 22786 7 1 2 41966 22785
0 22787 5 1 1 22786
0 22788 7 1 2 22787 56298
0 22789 5 1 1 22788
0 22790 7 1 2 55455 22789
0 22791 5 1 1 22790
0 22792 7 1 2 51597 58481
0 22793 5 1 1 22792
0 22794 7 1 2 47281 22793
0 22795 5 1 1 22794
0 22796 7 1 2 58102 51615
0 22797 7 1 2 22795 22796
0 22798 5 1 1 22797
0 22799 7 1 2 42649 22798
0 22800 5 1 1 22799
0 22801 7 1 2 22791 22800
0 22802 7 1 2 22783 22801
0 22803 5 1 1 22802
0 22804 7 1 2 63443 22803
0 22805 5 1 1 22804
0 22806 7 1 2 22767 22805
0 22807 5 2 1 22806
0 22808 7 1 2 46131 64806
0 22809 5 1 1 22808
0 22810 7 2 2 56077 61846
0 22811 7 1 2 51891 8629
0 22812 5 1 1 22811
0 22813 7 1 2 64808 22812
0 22814 5 1 1 22813
0 22815 7 1 2 22809 22814
0 22816 5 1 1 22815
0 22817 7 1 2 43001 22816
0 22818 5 1 1 22817
0 22819 7 3 2 44512 45312
0 22820 7 1 2 61219 64810
0 22821 7 1 2 54416 22820
0 22822 5 1 1 22821
0 22823 7 1 2 40641 48005
0 22824 7 1 2 62686 22823
0 22825 5 1 1 22824
0 22826 7 1 2 22822 22825
0 22827 5 1 1 22826
0 22828 7 1 2 58325 22827
0 22829 5 1 1 22828
0 22830 7 3 2 43718 63034
0 22831 5 1 1 64813
0 22832 7 1 2 22831 51241
0 22833 5 2 1 22832
0 22834 7 1 2 54431 56532
0 22835 7 1 2 64816 22834
0 22836 5 1 1 22835
0 22837 7 1 2 22829 22836
0 22838 5 1 1 22837
0 22839 7 1 2 43551 22838
0 22840 5 1 1 22839
0 22841 7 2 2 60221 54432
0 22842 7 1 2 64818 63366
0 22843 5 1 1 22842
0 22844 7 1 2 22840 22843
0 22845 5 1 1 22844
0 22846 7 2 2 56604 22845
0 22847 5 1 1 64820
0 22848 7 1 2 22818 22847
0 22849 5 1 1 22848
0 22850 7 1 2 62813 22849
0 22851 5 1 1 22850
0 22852 7 2 2 51083 55491
0 22853 5 1 1 64822
0 22854 7 1 2 58082 22853
0 22855 5 2 1 22854
0 22856 7 1 2 43719 64824
0 22857 5 1 1 22856
0 22858 7 2 2 46943 62538
0 22859 5 1 1 64826
0 22860 7 1 2 47788 64827
0 22861 5 1 1 22860
0 22862 7 2 2 40425 46921
0 22863 5 3 1 64828
0 22864 7 1 2 22861 64830
0 22865 7 1 2 22857 22864
0 22866 5 5 1 22865
0 22867 7 1 2 53759 64833
0 22868 5 1 1 22867
0 22869 7 4 2 42389 47553
0 22870 5 1 1 64838
0 22871 7 1 2 51873 64839
0 22872 5 1 1 22871
0 22873 7 6 2 48863 53413
0 22874 7 3 2 64842 52567
0 22875 5 1 1 64848
0 22876 7 1 2 22872 22875
0 22877 5 2 1 22876
0 22878 7 1 2 55315 64851
0 22879 5 1 1 22878
0 22880 7 1 2 22868 22879
0 22881 5 3 1 22880
0 22882 7 1 2 46132 64853
0 22883 5 1 1 22882
0 22884 7 2 2 55245 50486
0 22885 7 2 2 59799 64856
0 22886 5 1 1 64858
0 22887 7 1 2 47554 64859
0 22888 5 1 1 22887
0 22889 7 1 2 22883 22888
0 22890 5 2 1 22889
0 22891 7 4 2 57641 53645
0 22892 7 1 2 64862 63416
0 22893 7 1 2 64860 22892
0 22894 5 1 1 22893
0 22895 7 1 2 22851 22894
0 22896 5 1 1 22895
0 22897 7 1 2 46569 22896
0 22898 5 1 1 22897
0 22899 7 1 2 59954 64807
0 22900 5 1 1 22899
0 22901 7 1 2 48516 59052
0 22902 7 1 2 64854 22901
0 22903 5 1 1 22902
0 22904 7 1 2 22900 22903
0 22905 5 1 1 22904
0 22906 7 1 2 41027 22905
0 22907 5 1 1 22906
0 22908 7 2 2 64855 61565
0 22909 7 1 2 63697 64866
0 22910 5 1 1 22909
0 22911 7 1 2 22907 22910
0 22912 5 1 1 22911
0 22913 7 1 2 53911 22912
0 22914 5 1 1 22913
0 22915 7 1 2 48517 61560
0 22916 7 1 2 64867 22915
0 22917 5 1 1 22916
0 22918 7 1 2 22914 22917
0 22919 5 1 1 22918
0 22920 7 1 2 46133 22919
0 22921 5 1 1 22920
0 22922 7 1 2 12768 59971
0 22923 5 1 1 22922
0 22924 7 1 2 41234 22923
0 22925 5 1 1 22924
0 22926 7 1 2 9078 22925
0 22927 5 1 1 22926
0 22928 7 1 2 41028 22927
0 22929 5 1 1 22928
0 22930 7 1 2 47023 64368
0 22931 5 1 1 22930
0 22932 7 1 2 22929 22931
0 22933 5 1 1 22932
0 22934 7 1 2 53912 22933
0 22935 5 1 1 22934
0 22936 7 2 2 60637 46633
0 22937 7 1 2 64868 62359
0 22938 5 1 1 22937
0 22939 7 1 2 22935 22938
0 22940 5 1 1 22939
0 22941 7 1 2 61409 22940
0 22942 5 1 1 22941
0 22943 7 2 2 40964 56842
0 22944 7 1 2 64870 57993
0 22945 7 1 2 55492 22944
0 22946 5 1 1 22945
0 22947 7 1 2 22942 22946
0 22948 5 1 1 22947
0 22949 7 1 2 64809 22948
0 22950 5 1 1 22949
0 22951 7 1 2 22921 22950
0 22952 5 1 1 22951
0 22953 7 1 2 43002 22952
0 22954 5 1 1 22953
0 22955 7 1 2 64821 61849
0 22956 5 1 1 22955
0 22957 7 1 2 22954 22956
0 22958 5 1 1 22957
0 22959 7 1 2 64662 22958
0 22960 5 1 1 22959
0 22961 7 1 2 22898 22960
0 22962 5 1 1 22961
0 22963 7 1 2 43226 22962
0 22964 5 1 1 22963
0 22965 7 1 2 40248 58383
0 22966 5 1 1 22965
0 22967 7 1 2 22966 58294
0 22968 5 2 1 22967
0 22969 7 2 2 64024 52003
0 22970 7 1 2 64872 64874
0 22971 5 1 1 22970
0 22972 7 5 2 40426 41967
0 22973 5 2 1 64876
0 22974 7 1 2 64881 10658
0 22975 5 1 1 22974
0 22976 7 1 2 43385 22975
0 22977 5 3 1 22976
0 22978 7 1 2 40071 58110
0 22979 5 1 1 22978
0 22980 7 1 2 49335 22979
0 22981 5 1 1 22980
0 22982 7 1 2 42141 22981
0 22983 5 4 1 22982
0 22984 7 3 2 40427 44513
0 22985 5 4 1 64890
0 22986 7 4 2 43720 52813
0 22987 5 1 1 64897
0 22988 7 1 2 45474 64898
0 22989 5 2 1 22988
0 22990 7 1 2 64893 64901
0 22991 7 2 2 64886 22990
0 22992 5 1 1 64903
0 22993 7 2 2 64883 64904
0 22994 5 3 1 64905
0 22995 7 1 2 45738 64906
0 22996 5 1 1 22995
0 22997 7 1 2 46883 46933
0 22998 5 1 1 22997
0 22999 7 2 2 46885 22998
0 23000 5 1 1 64910
0 23001 7 1 2 42390 23000
0 23002 5 1 1 23001
0 23003 7 1 2 41371 23002
0 23004 7 1 2 22996 23003
0 23005 5 1 1 23004
0 23006 7 1 2 50490 51188
0 23007 7 2 2 64413 23006
0 23008 7 1 2 40249 64912
0 23009 5 1 1 23008
0 23010 7 2 2 46810 50584
0 23011 5 3 1 64914
0 23012 7 1 2 41235 64915
0 23013 5 1 1 23012
0 23014 7 1 2 23009 23013
0 23015 5 1 1 23014
0 23016 7 1 2 40072 23015
0 23017 5 1 1 23016
0 23018 7 1 2 55634 52734
0 23019 5 1 1 23018
0 23020 7 1 2 40250 50585
0 23021 5 1 1 23020
0 23022 7 1 2 48173 23021
0 23023 5 2 1 23022
0 23024 7 1 2 46875 64919
0 23025 5 1 1 23024
0 23026 7 1 2 23019 23025
0 23027 7 1 2 23017 23026
0 23028 5 1 1 23027
0 23029 7 1 2 40428 23028
0 23030 5 1 1 23029
0 23031 7 2 2 46893 59663
0 23032 7 1 2 48158 64921
0 23033 5 1 1 23032
0 23034 7 1 2 42650 23033
0 23035 7 1 2 23030 23034
0 23036 7 1 2 23005 23035
0 23037 5 1 1 23036
0 23038 7 2 2 50586 51317
0 23039 5 2 1 64923
0 23040 7 3 2 52035 58966
0 23041 7 5 2 49888 64927
0 23042 5 1 1 64930
0 23043 7 1 2 64925 23042
0 23044 5 1 1 23043
0 23045 7 1 2 44422 23044
0 23046 5 1 1 23045
0 23047 7 2 2 40429 50333
0 23048 7 1 2 44666 64935
0 23049 5 1 1 23048
0 23050 7 1 2 23046 23049
0 23051 5 1 1 23050
0 23052 7 1 2 43386 23051
0 23053 5 1 1 23052
0 23054 7 1 2 48822 22992
0 23055 5 1 1 23054
0 23056 7 1 2 45952 23055
0 23057 7 1 2 23053 23056
0 23058 5 1 1 23057
0 23059 7 1 2 46134 23058
0 23060 7 1 2 23037 23059
0 23061 5 1 1 23060
0 23062 7 1 2 22971 23061
0 23063 5 1 1 23062
0 23064 7 1 2 54612 23063
0 23065 5 1 1 23064
0 23066 7 3 2 43387 49447
0 23067 7 3 2 48372 64937
0 23068 7 1 2 62902 54531
0 23069 7 1 2 64940 23068
0 23070 5 1 1 23069
0 23071 7 1 2 23065 23070
0 23072 5 1 1 23071
0 23073 7 1 2 40642 23072
0 23074 5 1 1 23073
0 23075 7 1 2 63113 56661
0 23076 7 1 2 52677 23075
0 23077 5 1 1 23076
0 23078 7 1 2 57483 56304
0 23079 7 1 2 56234 23078
0 23080 5 1 1 23079
0 23081 7 1 2 23077 23080
0 23082 5 2 1 23081
0 23083 7 1 2 53582 64943
0 23084 5 1 1 23083
0 23085 7 1 2 23074 23084
0 23086 5 1 1 23085
0 23087 7 1 2 45108 23086
0 23088 5 1 1 23087
0 23089 7 2 2 49448 62440
0 23090 7 3 2 51054 64945
0 23091 5 1 1 64947
0 23092 7 2 2 2253 58143
0 23093 7 1 2 47087 64950
0 23094 5 1 1 23093
0 23095 7 1 2 23094 3179
0 23096 5 1 1 23095
0 23097 7 1 2 48389 23096
0 23098 5 1 1 23097
0 23099 7 1 2 23091 23098
0 23100 5 1 1 23099
0 23101 7 1 2 43388 23100
0 23102 5 1 1 23101
0 23103 7 2 2 43552 48823
0 23104 7 1 2 64952 62577
0 23105 5 1 1 23104
0 23106 7 2 2 23102 23105
0 23107 5 1 1 64954
0 23108 7 3 2 23107 59427
0 23109 5 1 1 64956
0 23110 7 1 2 64957 59179
0 23111 5 1 1 23110
0 23112 7 1 2 23088 23111
0 23113 5 1 1 23112
0 23114 7 1 2 41507 23113
0 23115 5 1 1 23114
0 23116 7 2 2 48564 59180
0 23117 7 1 2 64959 61346
0 23118 5 1 1 23117
0 23119 7 1 2 53299 64245
0 23120 7 6 2 45109 46135
0 23121 7 1 2 3479 64961
0 23122 7 1 2 23119 23121
0 23123 7 1 2 59671 23122
0 23124 5 1 1 23123
0 23125 7 1 2 23118 23124
0 23126 5 1 1 23125
0 23127 7 1 2 45739 23126
0 23128 5 1 1 23127
0 23129 7 4 2 44810 41812
0 23130 7 2 2 44667 64967
0 23131 7 1 2 47185 55352
0 23132 7 1 2 50060 23131
0 23133 7 1 2 64971 23132
0 23134 7 1 2 62203 23133
0 23135 5 1 1 23134
0 23136 7 1 2 23128 23135
0 23137 5 1 1 23136
0 23138 7 1 2 42142 23137
0 23139 5 1 1 23138
0 23140 7 1 2 60651 56469
0 23141 5 1 1 23140
0 23142 7 1 2 43921 23141
0 23143 5 1 1 23142
0 23144 7 1 2 42846 56214
0 23145 5 1 1 23144
0 23146 7 1 2 23143 23145
0 23147 5 1 1 23146
0 23148 7 2 2 48390 64938
0 23149 7 1 2 41813 58773
0 23150 7 1 2 64973 23149
0 23151 7 1 2 23147 23150
0 23152 5 1 1 23151
0 23153 7 1 2 23139 23152
0 23154 5 1 1 23153
0 23155 7 1 2 43122 23154
0 23156 5 1 1 23155
0 23157 7 2 2 47415 53610
0 23158 7 2 2 49803 64975
0 23159 7 2 2 47932 50587
0 23160 7 1 2 62508 59034
0 23161 7 1 2 64979 23160
0 23162 7 1 2 64977 23161
0 23163 5 1 1 23162
0 23164 7 1 2 23156 23163
0 23165 7 1 2 23115 23164
0 23166 5 1 1 23165
0 23167 7 1 2 44271 23166
0 23168 5 1 1 23167
0 23169 7 2 2 55019 54982
0 23170 7 2 2 50868 54542
0 23171 7 1 2 64946 64983
0 23172 5 1 1 23171
0 23173 7 1 2 54322 64951
0 23174 5 1 1 23173
0 23175 7 1 2 45740 60993
0 23176 5 1 1 23175
0 23177 7 1 2 23174 23176
0 23178 5 1 1 23177
0 23179 7 1 2 47088 23178
0 23180 5 1 1 23179
0 23181 7 1 2 54742 54417
0 23182 5 1 1 23181
0 23183 7 1 2 23180 23182
0 23184 5 1 1 23183
0 23185 7 1 2 42847 23184
0 23186 5 1 1 23185
0 23187 7 1 2 51203 55837
0 23188 5 1 1 23187
0 23189 7 1 2 23186 23188
0 23190 5 1 1 23189
0 23191 7 1 2 48391 23190
0 23192 5 1 1 23191
0 23193 7 1 2 23172 23192
0 23194 5 1 1 23193
0 23195 7 1 2 43389 23194
0 23196 5 1 1 23195
0 23197 7 1 2 44668 62448
0 23198 7 1 2 64984 23197
0 23199 5 1 1 23198
0 23200 7 1 2 23196 23199
0 23201 5 1 1 23200
0 23202 7 1 2 64981 23201
0 23203 5 1 1 23202
0 23204 7 1 2 23168 23203
0 23205 5 1 1 23204
0 23206 7 1 2 46570 23205
0 23207 5 1 1 23206
0 23208 7 1 2 58810 57470
0 23209 5 1 1 23208
0 23210 7 1 2 44514 56694
0 23211 5 1 1 23210
0 23212 7 1 2 23209 23211
0 23213 5 1 1 23212
0 23214 7 1 2 43553 23213
0 23215 5 1 1 23214
0 23216 7 1 2 43721 56695
0 23217 5 1 1 23216
0 23218 7 1 2 23215 23217
0 23219 5 1 1 23218
0 23220 7 1 2 44423 23219
0 23221 5 1 1 23220
0 23222 7 1 2 55419 64936
0 23223 5 1 1 23222
0 23224 7 1 2 23221 23223
0 23225 5 1 1 23224
0 23226 7 1 2 43390 23225
0 23227 5 1 1 23226
0 23228 7 2 2 51922 53545
0 23229 7 2 2 41236 55635
0 23230 5 1 1 64987
0 23231 7 3 2 64894 23230
0 23232 5 2 1 64989
0 23233 7 2 2 47735 56207
0 23234 5 1 1 64994
0 23235 7 1 2 54573 55845
0 23236 7 1 2 23234 23235
0 23237 5 1 1 23236
0 23238 7 1 2 64990 23237
0 23239 5 1 1 23238
0 23240 7 1 2 64985 23239
0 23241 5 1 1 23240
0 23242 7 1 2 23227 23241
0 23243 5 1 1 23242
0 23244 7 1 2 44669 23243
0 23245 5 1 1 23244
0 23246 7 1 2 64857 55448
0 23247 5 2 1 23246
0 23248 7 2 2 47789 56280
0 23249 5 2 1 64998
0 23250 7 2 2 56544 51854
0 23251 5 2 1 65002
0 23252 7 1 2 65000 65004
0 23253 5 3 1 23252
0 23254 7 1 2 53834 65006
0 23255 5 1 1 23254
0 23256 7 1 2 64996 23255
0 23257 5 1 1 23256
0 23258 7 1 2 40430 23257
0 23259 5 1 1 23258
0 23260 7 1 2 50167 62254
0 23261 5 3 1 23260
0 23262 7 1 2 65009 55218
0 23263 5 1 1 23262
0 23264 7 1 2 23259 23263
0 23265 5 1 1 23264
0 23266 7 1 2 47472 23265
0 23267 5 1 1 23266
0 23268 7 1 2 48159 60193
0 23269 5 2 1 23268
0 23270 7 1 2 53564 50168
0 23271 5 3 1 23270
0 23272 7 1 2 51841 65014
0 23273 5 1 1 23272
0 23274 7 2 2 40431 62647
0 23275 5 3 1 65017
0 23276 7 1 2 45741 65019
0 23277 7 1 2 23273 23276
0 23278 5 1 1 23277
0 23279 7 2 2 42391 58215
0 23280 5 1 1 65022
0 23281 7 1 2 41372 23280
0 23282 7 1 2 23278 23281
0 23283 5 1 1 23282
0 23284 7 1 2 65012 23283
0 23285 5 1 1 23284
0 23286 7 1 2 53835 23285
0 23287 5 1 1 23286
0 23288 7 1 2 23267 23287
0 23289 5 1 1 23288
0 23290 7 1 2 54613 23289
0 23291 5 1 1 23290
0 23292 7 1 2 23245 23291
0 23293 5 1 1 23292
0 23294 7 1 2 48518 23293
0 23295 5 1 1 23294
0 23296 7 1 2 55316 62483
0 23297 5 1 1 23296
0 23298 7 1 2 23297 15016
0 23299 5 1 1 23298
0 23300 7 1 2 45475 23299
0 23301 5 1 1 23300
0 23302 7 1 2 64153 59868
0 23303 5 1 1 23302
0 23304 7 1 2 61765 64805
0 23305 5 2 1 23304
0 23306 7 1 2 44515 50552
0 23307 5 6 1 23306
0 23308 7 1 2 65024 65026
0 23309 5 1 1 23308
0 23310 7 1 2 23303 23309
0 23311 7 1 2 23301 23310
0 23312 5 1 1 23311
0 23313 7 1 2 57790 23312
0 23314 5 1 1 23313
0 23315 7 1 2 47933 53238
0 23316 7 1 2 56662 23315
0 23317 7 1 2 49783 23316
0 23318 5 1 1 23317
0 23319 7 1 2 23314 23318
0 23320 5 1 1 23319
0 23321 7 1 2 42392 23320
0 23322 5 1 1 23321
0 23323 7 1 2 54360 64944
0 23324 5 1 1 23323
0 23325 7 1 2 62490 49922
0 23326 5 1 1 23325
0 23327 7 1 2 41508 23326
0 23328 5 1 1 23327
0 23329 7 1 2 59674 23328
0 23330 5 1 1 23329
0 23331 7 1 2 53851 23330
0 23332 5 1 1 23331
0 23333 7 2 2 51743 64226
0 23334 5 1 1 65032
0 23335 7 1 2 55246 49862
0 23336 7 1 2 65033 23335
0 23337 5 1 1 23336
0 23338 7 1 2 53836 56208
0 23339 5 1 1 23338
0 23340 7 1 2 55247 60194
0 23341 5 2 1 23340
0 23342 7 1 2 23339 65034
0 23343 5 1 1 23342
0 23344 7 1 2 41373 51263
0 23345 7 1 2 23343 23344
0 23346 5 1 1 23345
0 23347 7 1 2 23337 23346
0 23348 5 1 1 23347
0 23349 7 1 2 41509 23348
0 23350 5 1 1 23349
0 23351 7 1 2 23332 23350
0 23352 5 1 1 23351
0 23353 7 1 2 54614 56381
0 23354 7 1 2 23352 23353
0 23355 5 1 1 23354
0 23356 7 1 2 23324 23355
0 23357 7 1 2 23322 23356
0 23358 5 1 1 23357
0 23359 7 1 2 45313 23358
0 23360 5 1 1 23359
0 23361 7 1 2 23295 23360
0 23362 5 1 1 23361
0 23363 7 1 2 46634 23362
0 23364 5 1 1 23363
0 23365 7 1 2 63977 59293
0 23366 7 1 2 64861 23365
0 23367 5 1 1 23366
0 23368 7 1 2 23364 23367
0 23369 5 1 1 23368
0 23370 7 1 2 64663 23369
0 23371 5 1 1 23370
0 23372 7 1 2 23207 23371
0 23373 5 1 1 23372
0 23374 7 1 2 43227 23373
0 23375 5 1 1 23374
0 23376 7 1 2 60242 58589
0 23377 7 1 2 59672 23376
0 23378 5 1 1 23377
0 23379 7 1 2 53646 55981
0 23380 7 1 2 49551 23379
0 23381 5 1 1 23380
0 23382 7 1 2 23378 23381
0 23383 5 1 1 23382
0 23384 7 1 2 42848 23383
0 23385 5 1 1 23384
0 23386 7 1 2 43391 52108
0 23387 5 1 1 23386
0 23388 7 1 2 52075 62294
0 23389 5 1 1 23388
0 23390 7 1 2 9866 49945
0 23391 5 3 1 23390
0 23392 7 2 2 23389 65036
0 23393 5 2 1 65039
0 23394 7 2 2 23387 65040
0 23395 5 10 1 65043
0 23396 7 1 2 45476 65045
0 23397 5 1 1 23396
0 23398 7 1 2 55636 47899
0 23399 5 1 1 23398
0 23400 7 1 2 23397 23399
0 23401 5 1 1 23400
0 23402 7 1 2 41237 23401
0 23403 5 1 1 23402
0 23404 7 2 2 46898 61410
0 23405 5 1 1 65055
0 23406 7 1 2 45477 65056
0 23407 5 1 1 23406
0 23408 7 1 2 23403 23407
0 23409 5 3 1 23408
0 23410 7 3 2 49539 48772
0 23411 7 1 2 65057 65060
0 23412 5 1 1 23411
0 23413 7 1 2 47089 55493
0 23414 5 1 1 23413
0 23415 7 2 2 43554 45478
0 23416 7 1 2 56256 65063
0 23417 5 1 1 23416
0 23418 7 1 2 23414 23417
0 23419 5 1 1 23418
0 23420 7 1 2 48704 23419
0 23421 5 1 1 23420
0 23422 7 1 2 23412 23421
0 23423 5 1 1 23422
0 23424 7 1 2 45742 23423
0 23425 5 1 1 23424
0 23426 7 1 2 47790 59644
0 23427 5 1 1 23426
0 23428 7 1 2 47590 51385
0 23429 5 2 1 23428
0 23430 7 1 2 23427 65065
0 23431 5 1 1 23430
0 23432 7 2 2 23431 64504
0 23433 7 1 2 41374 65067
0 23434 5 1 1 23433
0 23435 7 1 2 42651 23434
0 23436 7 1 2 23425 23435
0 23437 5 1 1 23436
0 23438 7 3 2 47120 55681
0 23439 7 1 2 62942 65069
0 23440 5 1 1 23439
0 23441 7 1 2 56305 52804
0 23442 5 1 1 23441
0 23443 7 1 2 23440 23442
0 23444 5 1 1 23443
0 23445 7 1 2 43722 23444
0 23446 5 1 1 23445
0 23447 7 8 2 43555 40432
0 23448 7 3 2 43392 65072
0 23449 7 1 2 61220 58758
0 23450 7 1 2 65080 23449
0 23451 5 1 1 23450
0 23452 7 1 2 23446 23451
0 23453 5 1 1 23452
0 23454 7 1 2 41968 23453
0 23455 5 1 1 23454
0 23456 7 2 2 53565 55869
0 23457 5 13 1 65083
0 23458 7 3 2 47473 65085
0 23459 7 1 2 52327 48870
0 23460 7 1 2 65098 23459
0 23461 5 1 1 23460
0 23462 7 1 2 45953 23461
0 23463 7 1 2 23455 23462
0 23464 5 1 1 23463
0 23465 7 1 2 53546 23464
0 23466 7 1 2 23437 23465
0 23467 5 1 1 23466
0 23468 7 1 2 23385 23467
0 23469 5 1 1 23468
0 23470 7 8 2 64664 60295
0 23471 7 1 2 48519 65101
0 23472 7 1 2 23469 23471
0 23473 5 1 1 23472
0 23474 7 1 2 23375 23473
0 23475 5 1 1 23474
0 23476 7 1 2 49037 23475
0 23477 5 1 1 23476
0 23478 7 6 2 40251 43723
0 23479 7 1 2 65109 64072
0 23480 5 1 1 23479
0 23481 7 1 2 64260 60195
0 23482 7 1 2 47555 23481
0 23483 5 1 1 23482
0 23484 7 1 2 23480 23483
0 23485 5 1 1 23484
0 23486 7 1 2 45479 23485
0 23487 5 1 1 23486
0 23488 7 1 2 51356 58083
0 23489 5 1 1 23488
0 23490 7 1 2 55935 23489
0 23491 5 1 1 23490
0 23492 7 1 2 52043 64849
0 23493 5 1 1 23492
0 23494 7 5 2 43724 41238
0 23495 5 1 1 65115
0 23496 7 2 2 40252 65116
0 23497 5 1 1 65120
0 23498 7 1 2 64831 23497
0 23499 5 2 1 23498
0 23500 7 1 2 52004 65122
0 23501 5 1 1 23500
0 23502 7 1 2 23493 23501
0 23503 7 1 2 23491 23502
0 23504 5 1 1 23503
0 23505 7 1 2 45954 23504
0 23506 5 1 1 23505
0 23507 7 1 2 23487 23506
0 23508 5 1 1 23507
0 23509 7 2 2 45151 57265
0 23510 7 2 2 52642 65124
0 23511 7 1 2 23508 65126
0 23512 5 1 1 23511
0 23513 7 1 2 47121 50562
0 23514 5 1 1 23513
0 23515 7 1 2 52420 23514
0 23516 5 1 1 23515
0 23517 7 1 2 45314 23516
0 23518 5 2 1 23517
0 23519 7 1 2 51892 65128
0 23520 5 1 1 23519
0 23521 7 1 2 43725 23520
0 23522 5 1 1 23521
0 23523 7 1 2 52374 58373
0 23524 5 1 1 23523
0 23525 7 1 2 50721 52285
0 23526 5 1 1 23525
0 23527 7 1 2 23524 23526
0 23528 5 1 1 23527
0 23529 7 1 2 40433 23528
0 23530 5 1 1 23529
0 23531 7 1 2 47791 50160
0 23532 5 1 1 23531
0 23533 7 1 2 41969 64988
0 23534 5 1 1 23533
0 23535 7 1 2 23532 23534
0 23536 5 1 1 23535
0 23537 7 1 2 47474 23536
0 23538 5 1 1 23537
0 23539 7 1 2 23530 23538
0 23540 7 1 2 23522 23539
0 23541 5 1 1 23540
0 23542 7 1 2 59530 23541
0 23543 5 1 1 23542
0 23544 7 1 2 45480 49311
0 23545 5 1 1 23544
0 23546 7 2 2 46967 23545
0 23547 7 1 2 65130 55901
0 23548 5 1 1 23547
0 23549 7 1 2 59683 23548
0 23550 5 1 1 23549
0 23551 7 1 2 23543 23550
0 23552 5 1 1 23551
0 23553 7 1 2 44670 23552
0 23554 5 1 1 23553
0 23555 7 1 2 58163 50877
0 23556 5 1 1 23555
0 23557 7 1 2 47282 46991
0 23558 5 1 1 23557
0 23559 7 1 2 45315 47147
0 23560 7 1 2 23558 23559
0 23561 5 1 1 23560
0 23562 7 1 2 23556 23561
0 23563 5 1 1 23562
0 23564 7 1 2 43556 23563
0 23565 5 1 1 23564
0 23566 7 1 2 52849 61277
0 23567 5 1 1 23566
0 23568 7 1 2 23565 23567
0 23569 5 1 1 23568
0 23570 7 1 2 41375 59531
0 23571 7 1 2 23569 23570
0 23572 5 1 1 23571
0 23573 7 6 2 41837 62239
0 23574 5 2 1 65132
0 23575 7 1 2 55148 65133
0 23576 5 1 1 23575
0 23577 7 1 2 23572 23576
0 23578 7 1 2 23554 23577
0 23579 5 1 1 23578
0 23580 7 1 2 42652 23579
0 23581 5 1 1 23580
0 23582 7 2 2 41838 61617
0 23583 5 1 1 65140
0 23584 7 1 2 46502 46755
0 23585 5 1 1 23584
0 23586 7 1 2 43557 59738
0 23587 7 1 2 23585 23586
0 23588 5 1 1 23587
0 23589 7 1 2 23583 23588
0 23590 5 1 1 23589
0 23591 7 1 2 55456 52355
0 23592 7 1 2 23590 23591
0 23593 5 1 1 23592
0 23594 7 1 2 23581 23593
0 23595 5 1 1 23594
0 23596 7 1 2 42393 23595
0 23597 5 1 1 23596
0 23598 7 6 2 43393 45152
0 23599 7 2 2 63210 65142
0 23600 7 1 2 65148 54765
0 23601 5 1 1 23600
0 23602 7 2 2 45481 54532
0 23603 5 1 1 65150
0 23604 7 1 2 56257 58175
0 23605 5 1 1 23604
0 23606 7 1 2 23603 23605
0 23607 5 1 1 23606
0 23608 7 1 2 49297 59684
0 23609 7 1 2 23607 23608
0 23610 5 1 1 23609
0 23611 7 1 2 23601 23610
0 23612 5 1 1 23611
0 23613 7 1 2 48773 23612
0 23614 5 1 1 23613
0 23615 7 1 2 50886 55798
0 23616 5 2 1 23615
0 23617 7 1 2 48031 65152
0 23618 5 1 1 23617
0 23619 7 8 2 44516 41376
0 23620 7 1 2 50699 65154
0 23621 5 1 1 23620
0 23622 7 1 2 23618 23621
0 23623 5 1 1 23622
0 23624 7 1 2 59532 23623
0 23625 5 1 1 23624
0 23626 7 1 2 47090 59685
0 23627 5 1 1 23626
0 23628 7 1 2 23625 23627
0 23629 5 1 1 23628
0 23630 7 1 2 43558 23629
0 23631 5 1 1 23630
0 23632 7 1 2 48006 65141
0 23633 5 1 1 23632
0 23634 7 1 2 44671 59686
0 23635 5 2 1 23634
0 23636 7 2 2 54809 50295
0 23637 7 1 2 65143 60524
0 23638 7 1 2 63158 23637
0 23639 7 1 2 65164 23638
0 23640 5 1 1 23639
0 23641 7 1 2 65162 23640
0 23642 5 1 1 23641
0 23643 7 1 2 47660 23642
0 23644 5 1 1 23643
0 23645 7 1 2 23633 23644
0 23646 7 1 2 23631 23645
0 23647 5 1 1 23646
0 23648 7 1 2 43726 23647
0 23649 5 1 1 23648
0 23650 7 1 2 59687 58319
0 23651 5 1 1 23650
0 23652 7 1 2 23649 23651
0 23653 5 1 1 23652
0 23654 7 1 2 52456 23653
0 23655 5 1 1 23654
0 23656 7 1 2 23614 23655
0 23657 7 1 2 23597 23656
0 23658 5 1 1 23657
0 23659 7 1 2 56556 23658
0 23660 5 1 1 23659
0 23661 7 1 2 23512 23660
0 23662 5 1 1 23661
0 23663 7 1 2 55075 23662
0 23664 5 1 1 23663
0 23665 7 3 2 44672 41839
0 23666 7 1 2 62434 65166
0 23667 5 1 1 23666
0 23668 7 3 2 44517 46503
0 23669 7 4 2 45153 41970
0 23670 7 1 2 65169 65172
0 23671 7 1 2 53760 23670
0 23672 5 1 1 23671
0 23673 7 1 2 23667 23672
0 23674 5 1 1 23673
0 23675 7 1 2 64978 23674
0 23676 5 1 1 23675
0 23677 7 4 2 43228 54615
0 23678 7 3 2 41840 45955
0 23679 7 1 2 50766 65180
0 23680 7 1 2 65176 23679
0 23681 7 1 2 64911 23680
0 23682 5 1 1 23681
0 23683 7 1 2 23676 23682
0 23684 5 1 1 23683
0 23685 7 1 2 42143 23684
0 23686 5 1 1 23685
0 23687 7 1 2 64931 64976
0 23688 5 1 1 23687
0 23689 7 1 2 40253 46876
0 23690 5 1 1 23689
0 23691 7 1 2 23690 62389
0 23692 5 2 1 23691
0 23693 7 2 2 65183 61383
0 23694 7 1 2 53547 65185
0 23695 5 1 1 23694
0 23696 7 1 2 23688 23695
0 23697 5 1 1 23696
0 23698 7 1 2 42653 23697
0 23699 5 2 1 23698
0 23700 7 1 2 40254 10869
0 23701 5 1 1 23700
0 23702 7 2 2 58295 23701
0 23703 5 1 1 65189
0 23704 7 1 2 44673 51867
0 23705 5 1 1 23704
0 23706 7 2 2 46877 23705
0 23707 5 1 1 65191
0 23708 7 1 2 65190 23707
0 23709 5 1 1 23708
0 23710 7 1 2 40434 23709
0 23711 5 1 1 23710
0 23712 7 1 2 52510 59869
0 23713 5 1 1 23712
0 23714 7 1 2 23711 23713
0 23715 5 1 1 23714
0 23716 7 1 2 64986 23715
0 23717 5 1 1 23716
0 23718 7 1 2 65187 23717
0 23719 5 1 1 23718
0 23720 7 1 2 59688 23719
0 23721 5 1 1 23720
0 23722 7 1 2 23686 23721
0 23723 5 1 1 23722
0 23724 7 1 2 57642 23723
0 23725 5 1 1 23724
0 23726 7 1 2 64941 53619
0 23727 5 1 1 23726
0 23728 7 1 2 42394 23703
0 23729 5 1 1 23728
0 23730 7 3 2 40255 51242
0 23731 5 1 1 65193
0 23732 7 1 2 46873 23731
0 23733 5 2 1 23732
0 23734 7 1 2 48160 65196
0 23735 5 1 1 23734
0 23736 7 1 2 42395 65192
0 23737 5 1 1 23736
0 23738 7 1 2 23735 23737
0 23739 7 1 2 23729 23738
0 23740 5 1 1 23739
0 23741 7 1 2 40435 23740
0 23742 5 1 1 23741
0 23743 7 1 2 56281 64922
0 23744 5 1 1 23743
0 23745 7 1 2 23742 23744
0 23746 5 3 1 23745
0 23747 7 1 2 53548 65198
0 23748 5 1 1 23747
0 23749 7 1 2 23727 23748
0 23750 5 1 1 23749
0 23751 7 1 2 45956 23750
0 23752 5 1 1 23751
0 23753 7 1 2 65188 23752
0 23754 5 2 1 23753
0 23755 7 1 2 45154 59480
0 23756 7 1 2 65201 23755
0 23757 5 1 1 23756
0 23758 7 1 2 23725 23757
0 23759 7 1 2 23664 23758
0 23760 5 1 1 23759
0 23761 7 1 2 44311 23760
0 23762 5 1 1 23761
0 23763 7 5 2 42654 48824
0 23764 7 1 2 53611 65203
0 23765 5 2 1 23764
0 23766 7 1 2 53549 56151
0 23767 5 2 1 23766
0 23768 7 1 2 65208 65210
0 23769 5 2 1 23768
0 23770 7 4 2 64665 60470
0 23771 5 3 1 65214
0 23772 7 10 2 43229 46539
0 23773 5 1 1 65221
0 23774 7 2 2 65222 57643
0 23775 5 1 1 65231
0 23776 7 1 2 65218 23775
0 23777 5 1 1 23776
0 23778 7 1 2 64907 23777
0 23779 5 1 1 23778
0 23780 7 4 2 44312 57644
0 23781 7 3 2 45155 63159
0 23782 7 1 2 65073 65237
0 23783 5 1 1 23782
0 23784 7 1 2 45316 59689
0 23785 5 1 1 23784
0 23786 7 1 2 23783 23785
0 23787 5 1 1 23786
0 23788 7 1 2 47416 23787
0 23789 5 2 1 23788
0 23790 7 1 2 41239 59690
0 23791 5 2 1 23790
0 23792 7 1 2 47475 64811
0 23793 5 1 1 23792
0 23794 7 1 2 56302 23793
0 23795 5 1 1 23794
0 23796 7 1 2 40256 23795
0 23797 5 1 1 23796
0 23798 7 1 2 41841 51147
0 23799 5 1 1 23798
0 23800 7 1 2 23797 23799
0 23801 5 1 1 23800
0 23802 7 1 2 59739 23801
0 23803 5 1 1 23802
0 23804 7 1 2 65242 23803
0 23805 5 1 1 23804
0 23806 7 1 2 43727 23805
0 23807 5 1 1 23806
0 23808 7 1 2 65240 23807
0 23809 5 1 1 23808
0 23810 7 1 2 45482 23809
0 23811 5 1 1 23810
0 23812 7 1 2 64887 65020
0 23813 5 2 1 23812
0 23814 7 1 2 59691 65244
0 23815 5 2 1 23814
0 23816 7 3 2 46504 59782
0 23817 7 1 2 59725 65110
0 23818 7 1 2 65248 23817
0 23819 5 1 1 23818
0 23820 7 1 2 65246 23819
0 23821 7 1 2 23811 23820
0 23822 5 1 1 23821
0 23823 7 1 2 65233 23822
0 23824 5 1 1 23823
0 23825 7 1 2 23779 23824
0 23826 5 1 1 23825
0 23827 7 1 2 65212 23826
0 23828 5 1 1 23827
0 23829 7 1 2 44272 65202
0 23830 5 1 1 23829
0 23831 7 1 2 55027 23830
0 23832 5 1 1 23831
0 23833 7 1 2 52273 55989
0 23834 5 1 1 23833
0 23835 7 1 2 47876 48392
0 23836 5 1 1 23835
0 23837 7 1 2 23834 23836
0 23838 5 1 1 23837
0 23839 7 1 2 43394 23838
0 23840 5 1 1 23839
0 23841 7 1 2 43728 56124
0 23842 5 1 1 23841
0 23843 7 3 2 23840 23842
0 23844 5 1 1 65251
0 23845 7 4 2 50220 52274
0 23846 7 2 2 45743 65254
0 23847 5 1 1 65258
0 23848 7 1 2 23847 56246
0 23849 5 1 1 23848
0 23850 7 1 2 44674 23849
0 23851 5 1 1 23850
0 23852 7 1 2 65252 23851
0 23853 5 1 1 23852
0 23854 7 1 2 42655 23853
0 23855 5 1 1 23854
0 23856 7 1 2 55161 49540
0 23857 5 1 1 23856
0 23858 7 1 2 48774 55686
0 23859 7 1 2 58168 23858
0 23860 7 1 2 23857 23859
0 23861 5 1 1 23860
0 23862 7 1 2 23855 23861
0 23863 5 1 1 23862
0 23864 7 1 2 56557 23863
0 23865 5 1 1 23864
0 23866 7 1 2 57671 23865
0 23867 5 1 1 23866
0 23868 7 1 2 65223 23867
0 23869 7 1 2 23832 23868
0 23870 5 1 1 23869
0 23871 7 1 2 23828 23870
0 23872 7 1 2 23762 23871
0 23873 5 1 1 23872
0 23874 7 1 2 49038 23873
0 23875 5 1 1 23874
0 23876 7 1 2 45744 46951
0 23877 5 1 1 23876
0 23878 7 1 2 50679 23877
0 23879 5 3 1 23878
0 23880 7 1 2 47283 65260
0 23881 5 1 1 23880
0 23882 7 1 2 47476 50722
0 23883 7 1 2 57918 23882
0 23884 5 1 1 23883
0 23885 7 1 2 23881 23884
0 23886 5 1 1 23885
0 23887 7 1 2 47591 23886
0 23888 5 1 1 23887
0 23889 7 3 2 50283 56182
0 23890 7 1 2 47345 65263
0 23891 5 1 1 23890
0 23892 7 1 2 23888 23891
0 23893 5 1 1 23892
0 23894 7 1 2 62796 46571
0 23895 5 1 1 23894
0 23896 7 1 2 64666 61977
0 23897 5 2 1 23896
0 23898 7 1 2 23895 65266
0 23899 5 10 1 23898
0 23900 7 2 2 64441 65268
0 23901 7 1 2 23893 65278
0 23902 5 1 1 23901
0 23903 7 1 2 45745 50458
0 23904 7 1 2 60656 23903
0 23905 5 1 1 23904
0 23906 7 1 2 50680 23905
0 23907 5 1 1 23906
0 23908 7 1 2 57947 23907
0 23909 5 1 1 23908
0 23910 7 1 2 42396 46923
0 23911 5 1 1 23910
0 23912 7 1 2 47176 23911
0 23913 5 1 1 23912
0 23914 7 1 2 47187 64554
0 23915 7 1 2 9388 23914
0 23916 7 1 2 23913 23915
0 23917 5 1 1 23916
0 23918 7 1 2 23909 23917
0 23919 5 1 1 23918
0 23920 7 1 2 65269 23919
0 23921 5 1 1 23920
0 23922 7 1 2 64843 60110
0 23923 5 1 1 23922
0 23924 7 9 2 41842 48918
0 23925 7 3 2 62707 65280
0 23926 7 1 2 50588 65289
0 23927 5 1 1 23926
0 23928 7 1 2 23923 23927
0 23929 5 2 1 23928
0 23930 7 1 2 41240 65292
0 23931 5 1 1 23930
0 23932 7 1 2 60164 65261
0 23933 5 1 1 23932
0 23934 7 1 2 23931 23933
0 23935 5 1 1 23934
0 23936 7 1 2 44313 23935
0 23937 5 1 1 23936
0 23938 7 2 2 41241 50589
0 23939 5 1 1 65294
0 23940 7 2 2 48174 23939
0 23941 5 1 1 65296
0 23942 7 1 2 50681 65297
0 23943 5 4 1 23942
0 23944 7 3 2 46540 63574
0 23945 7 1 2 55893 54787
0 23946 7 1 2 65302 23945
0 23947 7 1 2 65298 23946
0 23948 5 1 1 23947
0 23949 7 1 2 23937 23948
0 23950 5 1 1 23949
0 23951 7 1 2 55076 23950
0 23952 5 1 1 23951
0 23953 7 2 2 57645 46572
0 23954 5 1 1 65305
0 23955 7 8 2 60077 64654
0 23956 5 1 1 65307
0 23957 7 1 2 23954 23956
0 23958 5 11 1 23957
0 23959 7 2 2 64844 54092
0 23960 5 1 1 65326
0 23961 7 2 2 45483 61895
0 23962 7 1 2 57617 65328
0 23963 5 1 1 23962
0 23964 7 1 2 23960 23963
0 23965 5 1 1 23964
0 23966 7 1 2 41242 23965
0 23967 5 1 1 23966
0 23968 7 1 2 53990 65262
0 23969 5 1 1 23968
0 23970 7 1 2 23967 23969
0 23971 5 1 1 23970
0 23972 7 1 2 65315 23971
0 23973 5 1 1 23972
0 23974 7 1 2 23952 23973
0 23975 5 1 1 23974
0 23976 7 1 2 41129 23975
0 23977 5 1 1 23976
0 23978 7 1 2 41130 65293
0 23979 5 1 1 23978
0 23980 7 1 2 45746 60141
0 23981 5 1 1 23980
0 23982 7 1 2 23979 23981
0 23983 5 1 1 23982
0 23984 7 1 2 44314 23983
0 23985 5 1 1 23984
0 23986 7 1 2 54788 64916
0 23987 5 2 1 23986
0 23988 7 1 2 65303 65330
0 23989 5 1 1 23988
0 23990 7 1 2 23985 23989
0 23991 5 1 1 23990
0 23992 7 1 2 55077 23991
0 23993 5 1 1 23992
0 23994 7 1 2 41131 65327
0 23995 5 1 1 23994
0 23996 7 1 2 57054 65331
0 23997 5 1 1 23996
0 23998 7 1 2 23995 23997
0 23999 5 1 1 23998
0 24000 7 1 2 65316 23999
0 24001 5 1 1 24000
0 24002 7 1 2 23993 24001
0 24003 5 1 1 24002
0 24004 7 1 2 40257 24003
0 24005 5 1 1 24004
0 24006 7 1 2 42397 52652
0 24007 5 1 1 24006
0 24008 7 1 2 41971 51194
0 24009 5 1 1 24008
0 24010 7 1 2 24007 24009
0 24011 5 1 1 24010
0 24012 7 1 2 43123 24011
0 24013 7 1 2 65270 24012
0 24014 5 1 1 24013
0 24015 7 1 2 24005 24014
0 24016 7 1 2 23977 24015
0 24017 5 1 1 24016
0 24018 7 1 2 40073 24017
0 24019 5 1 1 24018
0 24020 7 1 2 23921 24019
0 24021 5 1 1 24020
0 24022 7 1 2 45957 24021
0 24023 5 1 1 24022
0 24024 7 4 2 43124 47792
0 24025 7 1 2 65332 65264
0 24026 7 1 2 64189 24025
0 24027 7 1 2 65271 24026
0 24028 5 1 1 24027
0 24029 7 1 2 24023 24028
0 24030 5 1 1 24029
0 24031 7 1 2 43230 24030
0 24032 5 1 1 24031
0 24033 7 2 2 46417 46756
0 24034 7 4 2 47894 65336
0 24035 7 1 2 45156 62737
0 24036 5 1 1 24035
0 24037 7 2 2 57646 60133
0 24038 5 1 1 65342
0 24039 7 1 2 24036 24038
0 24040 5 1 1 24039
0 24041 7 1 2 44315 24040
0 24042 5 1 1 24041
0 24043 7 4 2 45157 58661
0 24044 7 2 2 44215 59594
0 24045 7 4 2 65344 65348
0 24046 5 1 1 65350
0 24047 7 1 2 24042 24046
0 24048 5 3 1 24047
0 24049 7 6 2 43231 65354
0 24050 7 1 2 65338 65357
0 24051 5 1 1 24050
0 24052 7 3 2 44316 59533
0 24053 7 1 2 50372 65363
0 24054 7 1 2 62814 24053
0 24055 5 1 1 24054
0 24056 7 1 2 24051 24055
0 24057 5 1 1 24056
0 24058 7 1 2 64261 24057
0 24059 5 1 1 24058
0 24060 7 3 2 51923 50846
0 24061 5 1 1 65366
0 24062 7 1 2 24061 53393
0 24063 5 1 1 24062
0 24064 7 1 2 60368 24063
0 24065 7 1 2 65272 24064
0 24066 5 1 1 24065
0 24067 7 1 2 24059 24066
0 24068 5 1 1 24067
0 24069 7 1 2 45484 24068
0 24070 5 1 1 24069
0 24071 7 1 2 54789 22870
0 24072 5 1 1 24071
0 24073 7 1 2 65279 24072
0 24074 5 1 1 24073
0 24075 7 1 2 24070 24074
0 24076 5 1 1 24075
0 24077 7 1 2 47592 24076
0 24078 5 1 1 24077
0 24079 7 1 2 24032 24078
0 24080 5 1 1 24079
0 24081 7 1 2 40436 24080
0 24082 5 1 1 24081
0 24083 7 1 2 23902 24082
0 24084 5 1 1 24083
0 24085 7 1 2 48121 24084
0 24086 5 1 1 24085
0 24087 7 1 2 50897 2552
0 24088 5 5 1 24087
0 24089 7 3 2 46505 65369
0 24090 7 2 2 49952 65374
0 24091 7 5 2 45158 42144
0 24092 7 1 2 43559 65379
0 24093 7 1 2 65377 24092
0 24094 5 1 1 24093
0 24095 7 1 2 65163 24094
0 24096 5 1 1 24095
0 24097 7 1 2 45747 24096
0 24098 5 1 1 24097
0 24099 7 5 2 45317 50590
0 24100 7 1 2 59692 65384
0 24101 5 1 1 24100
0 24102 7 1 2 24098 24101
0 24103 5 1 1 24102
0 24104 7 1 2 44518 24103
0 24105 5 1 1 24104
0 24106 7 3 2 41843 42398
0 24107 7 3 2 43232 65389
0 24108 7 1 2 55894 46957
0 24109 7 1 2 65392 24108
0 24110 7 1 2 59827 24109
0 24111 5 1 1 24110
0 24112 7 1 2 24105 24111
0 24113 5 1 1 24112
0 24114 7 1 2 58892 24113
0 24115 5 1 1 24114
0 24116 7 1 2 56195 47943
0 24117 5 1 1 24116
0 24118 7 1 2 41377 55990
0 24119 5 1 1 24118
0 24120 7 2 2 41243 53684
0 24121 5 1 1 65395
0 24122 7 1 2 24119 24121
0 24123 5 1 1 24122
0 24124 7 1 2 47417 24123
0 24125 5 1 1 24124
0 24126 7 1 2 24117 24125
0 24127 5 1 1 24126
0 24128 7 1 2 41972 24127
0 24129 5 1 1 24128
0 24130 7 1 2 58157 61706
0 24131 5 1 1 24130
0 24132 7 1 2 24129 24131
0 24133 5 1 1 24132
0 24134 7 1 2 43560 24133
0 24135 5 1 1 24134
0 24136 7 6 2 40258 44519
0 24137 7 1 2 53685 65397
0 24138 7 1 2 56258 24137
0 24139 5 1 1 24138
0 24140 7 1 2 24135 24139
0 24141 5 1 1 24140
0 24142 7 7 2 45159 46418
0 24143 7 1 2 65403 60296
0 24144 7 1 2 24141 24143
0 24145 5 1 1 24144
0 24146 7 1 2 24115 24145
0 24147 5 1 1 24146
0 24148 7 1 2 43729 24147
0 24149 5 1 1 24148
0 24150 7 3 2 59631 62927
0 24151 7 1 2 48615 65385
0 24152 5 1 1 24151
0 24153 7 1 2 42145 59404
0 24154 5 1 1 24153
0 24155 7 1 2 24152 24154
0 24156 5 1 1 24155
0 24157 7 1 2 44520 24156
0 24158 5 1 1 24157
0 24159 7 3 2 44675 50442
0 24160 5 1 1 65413
0 24161 7 1 2 43561 53382
0 24162 5 1 1 24161
0 24163 7 1 2 24160 24162
0 24164 5 1 1 24163
0 24165 7 1 2 43395 24164
0 24166 5 1 1 24165
0 24167 7 1 2 43562 64735
0 24168 5 1 1 24167
0 24169 7 1 2 24166 24168
0 24170 5 1 1 24169
0 24171 7 1 2 42399 24170
0 24172 5 1 1 24171
0 24173 7 1 2 24158 24172
0 24174 5 1 1 24173
0 24175 7 1 2 44424 24174
0 24176 5 1 1 24175
0 24177 7 1 2 51075 58127
0 24178 5 1 1 24177
0 24179 7 1 2 24176 24178
0 24180 5 1 1 24179
0 24181 7 1 2 65410 24180
0 24182 5 1 1 24181
0 24183 7 1 2 24149 24182
0 24184 5 1 1 24183
0 24185 7 1 2 48919 24184
0 24186 5 1 1 24185
0 24187 7 1 2 43730 50443
0 24188 5 2 1 24187
0 24189 7 1 2 43563 60924
0 24190 5 1 1 24189
0 24191 7 1 2 22185 24190
0 24192 5 1 1 24191
0 24193 7 1 2 43396 24192
0 24194 5 1 1 24193
0 24195 7 1 2 65416 24194
0 24196 5 1 1 24195
0 24197 7 1 2 44521 24196
0 24198 5 1 1 24197
0 24199 7 1 2 43564 60537
0 24200 5 1 1 24199
0 24201 7 1 2 58750 24200
0 24202 5 1 1 24201
0 24203 7 1 2 41378 24202
0 24204 5 1 1 24203
0 24205 7 1 2 49817 50045
0 24206 5 1 1 24205
0 24207 7 1 2 50444 24206
0 24208 5 1 1 24207
0 24209 7 1 2 24204 24208
0 24210 7 1 2 24198 24209
0 24211 5 1 1 24210
0 24212 7 1 2 42400 24211
0 24213 5 1 1 24212
0 24214 7 1 2 40437 60657
0 24215 5 2 1 24214
0 24216 7 1 2 47944 65418
0 24217 5 1 1 24216
0 24218 7 1 2 24213 24217
0 24219 5 1 1 24218
0 24220 7 3 2 43233 24219
0 24221 7 1 2 41844 65420
0 24222 5 1 1 24221
0 24223 7 1 2 60147 55915
0 24224 7 1 2 65378 24223
0 24225 5 1 1 24224
0 24226 7 1 2 24222 24225
0 24227 5 1 1 24226
0 24228 7 1 2 57647 24227
0 24229 5 1 1 24228
0 24230 7 1 2 60080 65421
0 24231 5 1 1 24230
0 24232 7 1 2 24229 24231
0 24233 5 1 1 24232
0 24234 7 1 2 53991 24233
0 24235 5 1 1 24234
0 24236 7 1 2 24186 24235
0 24237 5 1 1 24236
0 24238 7 1 2 44317 24237
0 24239 5 1 1 24238
0 24240 7 1 2 46541 62815
0 24241 7 1 2 65422 24240
0 24242 5 1 1 24241
0 24243 7 1 2 24239 24242
0 24244 5 1 1 24243
0 24245 7 1 2 42656 24244
0 24246 5 1 1 24245
0 24247 7 3 2 44318 44522
0 24248 7 1 2 65238 65423
0 24249 5 1 1 24248
0 24250 7 2 2 46573 61618
0 24251 5 1 1 65426
0 24252 7 1 2 24249 24251
0 24253 5 1 1 24252
0 24254 7 1 2 62797 24253
0 24255 5 1 1 24254
0 24256 7 5 2 41762 45160
0 24257 7 2 2 41814 65428
0 24258 7 2 2 43234 65433
0 24259 7 1 2 43397 64659
0 24260 7 1 2 65435 24259
0 24261 5 1 1 24260
0 24262 7 1 2 24255 24261
0 24263 5 1 1 24262
0 24264 7 2 2 48373 49449
0 24265 7 1 2 60596 65437
0 24266 7 1 2 24263 24265
0 24267 5 1 1 24266
0 24268 7 1 2 24246 24267
0 24269 5 1 1 24268
0 24270 7 1 2 48223 24269
0 24271 5 1 1 24270
0 24272 7 1 2 64834 65358
0 24273 5 1 1 24272
0 24274 7 2 2 41132 47122
0 24275 7 1 2 65439 52796
0 24276 5 1 1 24275
0 24277 7 1 2 45318 65099
0 24278 5 1 1 24277
0 24279 7 1 2 24276 24278
0 24280 5 2 1 24279
0 24281 7 1 2 65111 65441
0 24282 5 1 1 24281
0 24283 7 7 2 43398 40438
0 24284 7 3 2 48374 65443
0 24285 7 1 2 50878 65450
0 24286 5 1 1 24285
0 24287 7 1 2 24282 24286
0 24288 5 2 1 24287
0 24289 7 1 2 48920 65102
0 24290 7 1 2 65453 24289
0 24291 5 1 1 24290
0 24292 7 1 2 46419 24291
0 24293 7 1 2 24273 24292
0 24294 5 1 1 24293
0 24295 7 3 2 42849 48825
0 24296 7 2 2 54875 65455
0 24297 5 2 1 65458
0 24298 7 1 2 65460 55195
0 24299 5 4 1 24298
0 24300 7 1 2 50824 65086
0 24301 5 1 1 24300
0 24302 7 2 2 43565 50906
0 24303 5 2 1 65466
0 24304 7 1 2 24301 65468
0 24305 5 2 1 24304
0 24306 7 1 2 40439 65470
0 24307 5 2 1 24306
0 24308 7 1 2 47053 52421
0 24309 5 1 1 24308
0 24310 7 2 2 45319 24309
0 24311 5 1 1 65474
0 24312 7 1 2 53024 24311
0 24313 5 4 1 24312
0 24314 7 2 2 43731 65476
0 24315 5 2 1 65480
0 24316 7 1 2 65472 65482
0 24317 5 2 1 24316
0 24318 7 9 2 46506 64667
0 24319 7 1 2 62798 65486
0 24320 7 1 2 65484 24319
0 24321 5 1 1 24320
0 24322 7 1 2 42146 65027
0 24323 5 1 1 24322
0 24324 7 1 2 45320 58219
0 24325 7 1 2 24323 24324
0 24326 5 1 1 24325
0 24327 7 1 2 47477 51711
0 24328 5 1 1 24327
0 24329 7 1 2 58745 58096
0 24330 7 1 2 24328 24329
0 24331 5 1 1 24330
0 24332 7 1 2 24326 24331
0 24333 5 1 1 24332
0 24334 7 1 2 61078 24333
0 24335 5 1 1 24334
0 24336 7 1 2 43235 65273
0 24337 7 1 2 24335 24336
0 24338 5 1 1 24337
0 24339 7 1 2 43125 24338
0 24340 7 1 2 24321 24339
0 24341 5 1 1 24340
0 24342 7 1 2 65462 24341
0 24343 7 1 2 24294 24342
0 24344 5 1 1 24343
0 24345 7 1 2 24271 24344
0 24346 7 1 2 24086 24345
0 24347 7 1 2 23875 24346
0 24348 5 1 1 24347
0 24349 7 1 2 58018 24348
0 24350 5 1 1 24349
0 24351 7 3 2 43732 41133
0 24352 5 1 1 65495
0 24353 7 1 2 65070 65496
0 24354 5 1 1 24353
0 24355 7 2 2 54570 51143
0 24356 5 1 1 65498
0 24357 7 1 2 24354 24356
0 24358 5 2 1 24357
0 24359 7 1 2 65500 62859
0 24360 5 1 1 24359
0 24361 7 1 2 48382 49155
0 24362 5 4 1 24361
0 24363 7 1 2 45485 65502
0 24364 5 1 1 24363
0 24365 7 1 2 41244 51366
0 24366 5 1 1 24365
0 24367 7 1 2 24364 24366
0 24368 5 1 1 24367
0 24369 7 1 2 40440 62816
0 24370 7 1 2 24368 24369
0 24371 5 1 1 24370
0 24372 7 1 2 24360 24371
0 24373 5 1 1 24372
0 24374 7 1 2 53761 24373
0 24375 5 1 1 24374
0 24376 7 4 2 43399 59053
0 24377 5 1 1 65506
0 24378 7 1 2 44425 65507
0 24379 7 1 2 62843 24378
0 24380 5 1 1 24379
0 24381 7 1 2 14585 24380
0 24382 5 1 1 24381
0 24383 7 1 2 49804 65155
0 24384 7 1 2 56117 24383
0 24385 7 1 2 24382 24384
0 24386 5 1 1 24385
0 24387 7 1 2 24375 24386
0 24388 5 1 1 24387
0 24389 7 1 2 48122 24388
0 24390 5 1 1 24389
0 24391 7 1 2 59972 24377
0 24392 5 4 1 24391
0 24393 7 1 2 44273 65510
0 24394 5 1 1 24393
0 24395 7 1 2 59097 24394
0 24396 5 2 1 24395
0 24397 7 1 2 48921 65514
0 24398 5 1 1 24397
0 24399 7 1 2 62136 24398
0 24400 5 1 1 24399
0 24401 7 5 2 56092 54876
0 24402 5 1 1 65516
0 24403 7 1 2 65517 54817
0 24404 7 1 2 24400 24403
0 24405 5 1 1 24404
0 24406 7 1 2 24390 24405
0 24407 5 1 1 24406
0 24408 7 1 2 41973 24407
0 24409 5 1 1 24408
0 24410 7 1 2 50892 65081
0 24411 5 2 1 24410
0 24412 7 1 2 65483 65521
0 24413 5 1 1 24412
0 24414 7 1 2 53762 24413
0 24415 5 1 1 24414
0 24416 7 2 2 43400 52237
0 24417 5 1 1 65523
0 24418 7 2 2 48375 65524
0 24419 7 1 2 53462 65525
0 24420 5 1 1 24419
0 24421 7 1 2 64505 52415
0 24422 7 1 2 52563 24421
0 24423 5 1 1 24422
0 24424 7 1 2 24420 24423
0 24425 5 1 1 24424
0 24426 7 1 2 45321 24425
0 24427 5 1 1 24426
0 24428 7 1 2 24415 24427
0 24429 5 1 1 24428
0 24430 7 1 2 46136 24429
0 24431 5 1 1 24430
0 24432 7 2 2 55248 59865
0 24433 5 1 1 65527
0 24434 7 1 2 60196 51963
0 24435 7 1 2 65528 24434
0 24436 5 1 1 24435
0 24437 7 1 2 24431 24436
0 24438 5 1 1 24437
0 24439 7 1 2 62817 24438
0 24440 5 1 1 24439
0 24441 7 2 2 43733 57834
0 24442 7 1 2 65100 64389
0 24443 7 1 2 65529 24442
0 24444 7 1 2 55621 24443
0 24445 5 1 1 24444
0 24446 7 1 2 24440 24445
0 24447 5 1 1 24446
0 24448 7 1 2 43003 24447
0 24449 5 1 1 24448
0 24450 7 1 2 24409 24449
0 24451 5 1 1 24450
0 24452 7 4 2 41510 45161
0 24453 7 4 2 40643 44319
0 24454 7 2 2 46507 65535
0 24455 7 1 2 65531 65539
0 24456 7 1 2 24451 24455
0 24457 5 1 1 24456
0 24458 7 1 2 24350 24457
0 24459 7 1 2 23477 24458
0 24460 7 1 2 22964 24459
0 24461 5 1 1 24460
0 24462 7 1 2 49214 24461
0 24463 5 1 1 24462
0 24464 7 4 2 45958 58019
0 24465 7 1 2 57648 60207
0 24466 5 1 1 24465
0 24467 7 1 2 58904 24466
0 24468 5 1 1 24467
0 24469 7 1 2 48922 24468
0 24470 5 1 1 24469
0 24471 7 1 2 24470 62137
0 24472 5 1 1 24471
0 24473 7 1 2 65541 24472
0 24474 5 1 1 24473
0 24475 7 1 2 62818 63287
0 24476 5 1 1 24475
0 24477 7 1 2 24474 24476
0 24478 5 1 1 24477
0 24479 7 1 2 42850 24478
0 24480 5 1 1 24479
0 24481 7 2 2 62819 55392
0 24482 5 1 1 65545
0 24483 7 1 2 24480 24482
0 24484 5 1 1 24483
0 24485 7 1 2 49541 24484
0 24486 5 1 1 24485
0 24487 7 1 2 56800 58584
0 24488 7 2 2 45110 61932
0 24489 7 1 2 65547 57835
0 24490 7 1 2 24487 24489
0 24491 5 1 1 24490
0 24492 7 1 2 24486 24491
0 24493 5 1 1 24492
0 24494 7 1 2 42401 24493
0 24495 5 1 1 24494
0 24496 7 1 2 57512 60652
0 24497 5 13 1 24496
0 24498 7 1 2 43922 65549
0 24499 5 2 1 24498
0 24500 7 2 2 42851 54966
0 24501 7 3 2 55317 53432
0 24502 5 1 1 65566
0 24503 7 1 2 54337 24502
0 24504 5 1 1 24503
0 24505 7 1 2 65564 24504
0 24506 5 1 1 24505
0 24507 7 1 2 65562 24506
0 24508 5 1 1 24507
0 24509 7 1 2 62820 54780
0 24510 7 1 2 24508 24509
0 24511 5 1 1 24510
0 24512 7 1 2 24495 24511
0 24513 5 1 1 24512
0 24514 7 1 2 47284 24513
0 24515 5 1 1 24514
0 24516 7 5 2 43923 53295
0 24517 5 1 1 65569
0 24518 7 2 2 40644 54361
0 24519 5 1 1 65574
0 24520 7 1 2 24517 24519
0 24521 5 11 1 24520
0 24522 7 1 2 42852 65576
0 24523 5 1 1 24522
0 24524 7 1 2 55396 24523
0 24525 5 5 1 24524
0 24526 7 1 2 47974 55923
0 24527 7 1 2 62821 24526
0 24528 7 1 2 65587 24527
0 24529 5 1 1 24528
0 24530 7 1 2 24515 24529
0 24531 5 1 1 24530
0 24532 7 1 2 40259 24531
0 24533 5 1 1 24532
0 24534 7 2 2 58572 56887
0 24535 7 1 2 58020 61906
0 24536 7 1 2 65592 24535
0 24537 7 1 2 65367 24536
0 24538 5 1 1 24537
0 24539 7 1 2 24533 24538
0 24540 5 1 1 24539
0 24541 7 1 2 43004 24540
0 24542 5 1 1 24541
0 24543 7 2 2 59003 50090
0 24544 7 1 2 41134 45111
0 24545 7 1 2 52511 24544
0 24546 7 1 2 65594 24545
0 24547 7 1 2 57609 24546
0 24548 7 1 2 56696 24547
0 24549 5 1 1 24548
0 24550 7 1 2 24542 24549
0 24551 5 1 1 24550
0 24552 7 1 2 47123 24551
0 24553 5 1 1 24552
0 24554 7 1 2 40645 46960
0 24555 5 1 1 24554
0 24556 7 1 2 51848 60832
0 24557 5 1 1 24556
0 24558 7 1 2 41135 63456
0 24559 5 1 1 24558
0 24560 7 1 2 24557 24559
0 24561 5 1 1 24560
0 24562 7 1 2 41379 24561
0 24563 5 1 1 24562
0 24564 7 1 2 24555 24563
0 24565 5 3 1 24564
0 24566 7 1 2 40074 65596
0 24567 5 1 1 24566
0 24568 7 1 2 53566 51166
0 24569 5 2 1 24568
0 24570 7 1 2 43924 52993
0 24571 5 1 1 24570
0 24572 7 3 2 65599 24571
0 24573 5 1 1 65601
0 24574 7 1 2 24567 24573
0 24575 5 1 1 24574
0 24576 7 1 2 40441 24575
0 24577 5 1 1 24576
0 24578 7 1 2 40646 63100
0 24579 5 1 1 24578
0 24580 7 1 2 24577 24579
0 24581 5 1 1 24580
0 24582 7 1 2 45748 24581
0 24583 5 1 1 24582
0 24584 7 1 2 62070 52251
0 24585 5 2 1 24584
0 24586 7 2 2 65604 50675
0 24587 5 1 1 65606
0 24588 7 1 2 65607 53320
0 24589 5 1 1 24588
0 24590 7 1 2 42853 24589
0 24591 7 1 2 24583 24590
0 24592 5 1 1 24591
0 24593 7 1 2 46137 64955
0 24594 5 1 1 24593
0 24595 7 1 2 42657 24594
0 24596 7 1 2 24592 24595
0 24597 5 1 1 24596
0 24598 7 1 2 56512 3797
0 24599 5 3 1 24598
0 24600 7 1 2 56249 52259
0 24601 5 1 1 24600
0 24602 7 1 2 58233 24601
0 24603 5 1 1 24602
0 24604 7 1 2 43401 24603
0 24605 5 1 1 24604
0 24606 7 1 2 41245 50611
0 24607 5 1 1 24606
0 24608 7 1 2 52039 51065
0 24609 7 1 2 24607 24608
0 24610 5 1 1 24609
0 24611 7 1 2 24605 24610
0 24612 5 1 1 24611
0 24613 7 1 2 65608 24612
0 24614 5 1 1 24613
0 24615 7 1 2 50251 56078
0 24616 5 1 1 24615
0 24617 7 1 2 43566 64817
0 24618 5 1 1 24617
0 24619 7 1 2 9384 24618
0 24620 5 1 1 24619
0 24621 7 2 2 24620 59239
0 24622 7 1 2 42402 65611
0 24623 5 1 1 24622
0 24624 7 1 2 24616 24623
0 24625 5 1 1 24624
0 24626 7 1 2 42147 24625
0 24627 5 1 1 24626
0 24628 7 1 2 45749 64803
0 24629 5 1 1 24628
0 24630 7 1 2 24587 24629
0 24631 5 1 1 24630
0 24632 7 1 2 41246 24631
0 24633 5 1 1 24632
0 24634 7 1 2 64100 54781
0 24635 5 1 1 24634
0 24636 7 1 2 24633 24635
0 24637 5 1 1 24636
0 24638 7 1 2 42854 24637
0 24639 5 1 1 24638
0 24640 7 1 2 24627 24639
0 24641 5 1 1 24640
0 24642 7 1 2 54821 24641
0 24643 5 1 1 24642
0 24644 7 1 2 24614 24643
0 24645 7 1 2 24597 24644
0 24646 5 1 1 24645
0 24647 7 1 2 41511 24646
0 24648 5 1 1 24647
0 24649 7 4 2 41974 55412
0 24650 7 1 2 61273 65613
0 24651 7 1 2 49784 24650
0 24652 5 1 1 24651
0 24653 7 3 2 41247 56801
0 24654 7 2 2 53005 65617
0 24655 5 1 1 65620
0 24656 7 1 2 42658 65621
0 24657 7 1 2 55645 24656
0 24658 5 1 1 24657
0 24659 7 1 2 24652 24658
0 24660 5 1 1 24659
0 24661 7 1 2 45750 24660
0 24662 5 1 1 24661
0 24663 7 2 2 45959 56413
0 24664 7 1 2 50123 64924
0 24665 7 1 2 65622 24664
0 24666 5 1 1 24665
0 24667 7 2 2 24662 24666
0 24668 5 2 1 65624
0 24669 7 3 2 41248 65605
0 24670 7 1 2 65628 53006
0 24671 5 1 1 24670
0 24672 7 1 2 42148 65612
0 24673 5 1 1 24672
0 24674 7 1 2 24671 24673
0 24675 5 1 1 24674
0 24676 7 1 2 45960 24675
0 24677 5 1 1 24676
0 24678 7 1 2 63465 65255
0 24679 5 1 1 24678
0 24680 7 1 2 24677 24679
0 24681 5 1 1 24680
0 24682 7 1 2 40647 24681
0 24683 5 1 1 24682
0 24684 7 1 2 45486 65623
0 24685 7 1 2 63116 24684
0 24686 5 2 1 24685
0 24687 7 1 2 42403 65631
0 24688 7 1 2 24683 24687
0 24689 5 1 1 24688
0 24690 7 1 2 1684 2914
0 24691 5 1 1 24690
0 24692 7 1 2 56898 24691
0 24693 5 1 1 24692
0 24694 7 1 2 48705 2455
0 24695 5 1 1 24694
0 24696 7 1 2 50962 24695
0 24697 5 1 1 24696
0 24698 7 4 2 40648 45487
0 24699 5 1 1 65633
0 24700 7 1 2 5058 24699
0 24701 5 1 1 24700
0 24702 7 1 2 49686 24701
0 24703 7 1 2 24697 24702
0 24704 5 1 1 24703
0 24705 7 1 2 24693 24704
0 24706 5 1 1 24705
0 24707 7 1 2 45322 24706
0 24708 5 1 1 24707
0 24709 7 1 2 65618 52182
0 24710 5 1 1 24709
0 24711 7 1 2 24708 24710
0 24712 5 1 1 24711
0 24713 7 1 2 42855 24712
0 24714 5 1 1 24713
0 24715 7 1 2 47934 52183
0 24716 5 2 1 24715
0 24717 7 1 2 63913 65637
0 24718 5 1 1 24717
0 24719 7 2 2 52669 52971
0 24720 7 1 2 24718 65639
0 24721 5 1 1 24720
0 24722 7 2 2 47285 65565
0 24723 7 1 2 45961 63014
0 24724 7 1 2 47070 24723
0 24725 7 1 2 65641 24724
0 24726 5 1 1 24725
0 24727 7 1 2 24721 24726
0 24728 5 1 1 24727
0 24729 7 1 2 41975 24728
0 24730 5 1 1 24729
0 24731 7 3 2 46138 55833
0 24732 7 2 2 44523 65643
0 24733 5 1 1 65646
0 24734 7 1 2 40649 65647
0 24735 5 1 1 24734
0 24736 7 1 2 45751 24735
0 24737 7 1 2 24730 24736
0 24738 7 1 2 24714 24737
0 24739 5 1 1 24738
0 24740 7 1 2 44811 24739
0 24741 7 1 2 24689 24740
0 24742 5 1 1 24741
0 24743 7 1 2 65625 24742
0 24744 7 1 2 24648 24743
0 24745 5 1 1 24744
0 24746 7 1 2 43005 24745
0 24747 5 1 1 24746
0 24748 7 2 2 48520 64175
0 24749 5 1 1 65648
0 24750 7 3 2 44426 46287
0 24751 7 2 2 54274 65650
0 24752 7 1 2 50334 50119
0 24753 7 1 2 65653 24752
0 24754 5 1 1 24753
0 24755 7 1 2 24749 24754
0 24756 5 1 1 24755
0 24757 7 1 2 42856 24756
0 24758 5 1 1 24757
0 24759 7 1 2 48376 60791
0 24760 5 1 1 24759
0 24761 7 1 2 52467 24760
0 24762 5 1 1 24761
0 24763 7 1 2 58021 24762
0 24764 5 1 1 24763
0 24765 7 2 2 53215 50660
0 24766 5 3 1 65655
0 24767 7 1 2 24764 65657
0 24768 5 1 1 24767
0 24769 7 1 2 48123 24768
0 24770 5 1 1 24769
0 24771 7 1 2 24758 24770
0 24772 5 1 1 24771
0 24773 7 1 2 43402 24772
0 24774 5 1 1 24773
0 24775 7 1 2 40650 65550
0 24776 5 2 1 24775
0 24777 7 1 2 46139 61144
0 24778 5 1 1 24777
0 24779 7 1 2 65660 24778
0 24780 5 2 1 24779
0 24781 7 1 2 43006 59260
0 24782 7 1 2 65662 24781
0 24783 5 1 1 24782
0 24784 7 1 2 24774 24783
0 24785 5 1 1 24784
0 24786 7 1 2 43734 24785
0 24787 5 1 1 24786
0 24788 7 1 2 41512 56507
0 24789 5 1 1 24788
0 24790 7 1 2 65661 24789
0 24791 5 1 1 24790
0 24792 7 2 2 45752 55149
0 24793 5 1 1 65664
0 24794 7 1 2 43007 65665
0 24795 7 1 2 24791 24794
0 24796 5 1 1 24795
0 24797 7 1 2 24787 24796
0 24798 5 1 1 24797
0 24799 7 1 2 48007 24798
0 24800 5 1 1 24799
0 24801 7 1 2 45323 62492
0 24802 5 1 1 24801
0 24803 7 1 2 49713 61454
0 24804 5 1 1 24803
0 24805 7 1 2 44676 50847
0 24806 7 1 2 24804 24805
0 24807 5 1 1 24806
0 24808 7 1 2 24802 24807
0 24809 5 1 1 24808
0 24810 7 2 2 45488 24809
0 24811 5 1 1 65666
0 24812 7 1 2 55891 49830
0 24813 5 1 1 24812
0 24814 7 1 2 24811 24813
0 24815 5 1 1 24814
0 24816 7 2 2 45962 24815
0 24817 5 1 1 65668
0 24818 7 1 2 56705 65629
0 24819 5 1 1 24818
0 24820 7 1 2 24817 24819
0 24821 5 1 1 24820
0 24822 7 1 2 48124 24821
0 24823 5 1 1 24822
0 24824 7 1 2 45489 58160
0 24825 5 1 1 24824
0 24826 7 1 2 64814 24825
0 24827 5 1 1 24826
0 24828 7 1 2 24827 51772
0 24829 5 1 1 24828
0 24830 7 1 2 43567 24829
0 24831 5 1 1 24830
0 24832 7 1 2 24831 24417
0 24833 5 1 1 24832
0 24834 7 1 2 44677 48224
0 24835 7 2 2 24833 24834
0 24836 5 1 1 65670
0 24837 7 1 2 42659 65671
0 24838 5 1 1 24837
0 24839 7 1 2 24823 24838
0 24840 5 1 1 24839
0 24841 7 1 2 42404 24840
0 24842 5 1 1 24841
0 24843 7 1 2 53837 56240
0 24844 5 1 1 24843
0 24845 7 1 2 64025 61047
0 24846 5 1 1 24845
0 24847 7 1 2 24844 24846
0 24848 5 1 1 24847
0 24849 7 1 2 41380 24848
0 24850 5 1 1 24849
0 24851 7 1 2 63030 55812
0 24852 5 1 1 24851
0 24853 7 1 2 24850 24852
0 24854 5 1 1 24853
0 24855 7 1 2 45490 24854
0 24856 5 1 1 24855
0 24857 7 1 2 42660 50252
0 24858 5 1 1 24857
0 24859 7 1 2 50837 54301
0 24860 5 1 1 24859
0 24861 7 1 2 24858 24860
0 24862 5 1 1 24861
0 24863 7 1 2 42149 24862
0 24864 5 1 1 24863
0 24865 7 1 2 50152 55318
0 24866 5 1 1 24865
0 24867 7 1 2 44427 58746
0 24868 5 1 1 24867
0 24869 7 1 2 47939 24868
0 24870 5 1 1 24869
0 24871 7 1 2 43403 24870
0 24872 5 2 1 24871
0 24873 7 1 2 48424 65672
0 24874 5 1 1 24873
0 24875 7 1 2 43568 24874
0 24876 5 1 1 24875
0 24877 7 2 2 43735 50237
0 24878 5 1 1 65674
0 24879 7 1 2 44678 65675
0 24880 5 2 1 24879
0 24881 7 1 2 24876 65676
0 24882 5 1 1 24881
0 24883 7 1 2 45963 24882
0 24884 5 1 1 24883
0 24885 7 1 2 24866 24884
0 24886 7 1 2 24864 24885
0 24887 5 1 1 24886
0 24888 7 1 2 46140 24887
0 24889 5 1 1 24888
0 24890 7 1 2 24856 24889
0 24891 5 1 1 24890
0 24892 7 1 2 51292 24891
0 24893 5 1 1 24892
0 24894 7 1 2 24842 24893
0 24895 5 1 1 24894
0 24896 7 1 2 49603 24895
0 24897 5 1 1 24896
0 24898 7 1 2 24800 24897
0 24899 7 1 2 24747 24898
0 24900 5 1 1 24899
0 24901 7 1 2 62822 24900
0 24902 5 1 1 24901
0 24903 7 2 2 46420 58662
0 24904 7 2 2 40260 59004
0 24905 7 1 2 65678 65680
0 24906 5 1 1 24905
0 24907 7 1 2 17703 24906
0 24908 5 1 1 24907
0 24909 7 1 2 55444 24908
0 24910 5 1 1 24909
0 24911 7 2 2 50749 56593
0 24912 7 1 2 57453 62089
0 24913 7 1 2 65682 24912
0 24914 5 1 1 24913
0 24915 7 1 2 24910 24914
0 24916 5 1 1 24915
0 24917 7 1 2 55249 24916
0 24918 5 1 1 24917
0 24919 7 1 2 61168 63841
0 24920 7 1 2 63868 24919
0 24921 7 1 2 65010 24920
0 24922 5 1 1 24921
0 24923 7 1 2 24918 24922
0 24924 5 1 1 24923
0 24925 7 1 2 42405 24924
0 24926 5 1 1 24925
0 24927 7 1 2 40075 55457
0 24928 5 1 1 24927
0 24929 7 1 2 61766 24928
0 24930 5 3 1 24929
0 24931 7 1 2 58573 62022
0 24932 7 1 2 60951 24931
0 24933 7 1 2 64753 24932
0 24934 7 1 2 65684 24933
0 24935 5 1 1 24934
0 24936 7 1 2 24926 24935
0 24937 5 1 1 24936
0 24938 7 1 2 58022 24937
0 24939 5 1 1 24938
0 24940 7 2 2 47994 59955
0 24941 5 1 1 65687
0 24942 7 1 2 47024 63955
0 24943 5 1 1 24942
0 24944 7 1 2 24941 24943
0 24945 5 1 1 24944
0 24946 7 1 2 56852 24945
0 24947 5 1 1 24946
0 24948 7 1 2 59054 65007
0 24949 5 1 1 24948
0 24950 7 1 2 65688 63324
0 24951 5 1 1 24950
0 24952 7 1 2 24949 24951
0 24953 5 1 1 24952
0 24954 7 1 2 24953 56861
0 24955 5 1 1 24954
0 24956 7 1 2 24947 24955
0 24957 5 1 1 24956
0 24958 7 1 2 44274 24957
0 24959 5 1 1 24958
0 24960 7 2 2 43126 47995
0 24961 7 1 2 62866 65689
0 24962 7 2 2 56990 24961
0 24963 7 1 2 61812 65691
0 24964 5 1 1 24963
0 24965 7 1 2 24959 24964
0 24966 5 1 1 24965
0 24967 7 1 2 48923 24966
0 24968 5 1 1 24967
0 24969 7 1 2 40076 61543
0 24970 7 1 2 65692 24969
0 24971 5 1 1 24970
0 24972 7 1 2 24968 24971
0 24973 5 1 1 24972
0 24974 7 1 2 42661 24973
0 24975 5 1 1 24974
0 24976 7 1 2 45491 50661
0 24977 7 3 2 57454 52775
0 24978 7 1 2 24976 65693
0 24979 7 1 2 64611 24978
0 24980 7 1 2 64541 24979
0 24981 5 1 1 24980
0 24982 7 1 2 24975 24981
0 24983 5 1 1 24982
0 24984 7 1 2 40442 24983
0 24985 5 1 1 24984
0 24986 7 1 2 24939 24985
0 24987 5 1 1 24986
0 24988 7 1 2 43008 24987
0 24989 5 1 1 24988
0 24990 7 2 2 64754 55420
0 24991 7 1 2 61933 60845
0 24992 7 1 2 65696 24991
0 24993 5 1 1 24992
0 24994 7 1 2 24989 24993
0 24995 5 1 1 24994
0 24996 7 1 2 46757 24995
0 24997 5 1 1 24996
0 24998 7 1 2 65546 65299
0 24999 5 1 1 24998
0 25000 7 2 2 44812 62823
0 25001 7 1 2 65698 56118
0 25002 5 1 1 25001
0 25003 7 1 2 54323 65300
0 25004 7 1 2 62147 25003
0 25005 5 1 1 25004
0 25006 7 1 2 25002 25005
0 25007 5 1 1 25006
0 25008 7 1 2 40651 25007
0 25009 5 1 1 25008
0 25010 7 5 2 45492 64262
0 25011 7 1 2 41249 65700
0 25012 5 1 1 25011
0 25013 7 1 2 64341 25012
0 25014 5 2 1 25013
0 25015 7 1 2 58023 65705
0 25016 7 1 2 62148 25015
0 25017 5 1 1 25016
0 25018 7 3 2 50662 57685
0 25019 7 1 2 60885 17867
0 25020 5 1 1 25019
0 25021 7 1 2 65707 25020
0 25022 7 1 2 62799 25021
0 25023 5 1 1 25022
0 25024 7 1 2 25017 25023
0 25025 7 1 2 25009 25024
0 25026 5 1 1 25025
0 25027 7 1 2 42857 25026
0 25028 5 1 1 25027
0 25029 7 1 2 24999 25028
0 25030 5 1 1 25029
0 25031 7 1 2 40443 25030
0 25032 5 1 1 25031
0 25033 7 3 2 46421 58024
0 25034 7 3 2 45112 45493
0 25035 7 1 2 63842 65713
0 25036 7 1 2 65683 25035
0 25037 7 1 2 55617 25036
0 25038 7 1 2 65710 25037
0 25039 5 1 1 25038
0 25040 7 1 2 25032 25039
0 25041 5 1 1 25040
0 25042 7 1 2 43009 25041
0 25043 5 1 1 25042
0 25044 7 1 2 56599 64131
0 25045 7 1 2 65697 25044
0 25046 5 1 1 25045
0 25047 7 1 2 25043 25046
0 25048 5 1 1 25047
0 25049 7 1 2 52109 25048
0 25050 5 1 1 25049
0 25051 7 1 2 51953 58164
0 25052 5 1 1 25051
0 25053 7 1 2 42150 25052
0 25054 5 1 1 25053
0 25055 7 1 2 50230 65414
0 25056 5 2 1 25055
0 25057 7 1 2 25054 65716
0 25058 5 1 1 25057
0 25059 7 1 2 41513 25058
0 25060 5 1 1 25059
0 25061 7 1 2 46811 56700
0 25062 5 1 1 25061
0 25063 7 1 2 25060 25062
0 25064 5 1 1 25063
0 25065 7 1 2 40261 25064
0 25066 5 1 1 25065
0 25067 7 1 2 55925 51954
0 25068 5 3 1 25067
0 25069 7 1 2 41250 60882
0 25070 7 1 2 65718 25069
0 25071 5 1 1 25070
0 25072 7 1 2 25066 25071
0 25073 5 1 1 25072
0 25074 7 1 2 45753 25073
0 25075 5 1 1 25074
0 25076 7 1 2 41514 60201
0 25077 5 1 1 25076
0 25078 7 1 2 43925 25077
0 25079 7 1 2 25075 25078
0 25080 5 1 1 25079
0 25081 7 1 2 47793 65719
0 25082 5 1 1 25081
0 25083 7 1 2 58216 25082
0 25084 5 1 1 25083
0 25085 7 1 2 42151 25084
0 25086 5 1 1 25085
0 25087 7 1 2 50245 65415
0 25088 5 1 1 25087
0 25089 7 1 2 25086 25088
0 25090 5 1 1 25089
0 25091 7 1 2 45754 25090
0 25092 5 1 1 25091
0 25093 7 1 2 25092 9358
0 25094 5 1 1 25093
0 25095 7 1 2 44813 25094
0 25096 5 1 1 25095
0 25097 7 1 2 55940 64932
0 25098 5 1 1 25097
0 25099 7 1 2 40652 25098
0 25100 7 1 2 25096 25099
0 25101 5 1 1 25100
0 25102 7 1 2 42858 25101
0 25103 7 1 2 25080 25102
0 25104 5 1 1 25103
0 25105 7 1 2 48183 64917
0 25106 5 1 1 25105
0 25107 7 1 2 43736 25106
0 25108 5 1 1 25107
0 25109 7 1 2 60032 48025
0 25110 5 1 1 25109
0 25111 7 1 2 25108 25110
0 25112 5 1 1 25111
0 25113 7 2 2 44679 25112
0 25114 7 1 2 58025 65721
0 25115 5 1 1 25114
0 25116 7 1 2 47975 51874
0 25117 5 1 1 25116
0 25118 7 2 2 47794 64845
0 25119 5 1 1 65723
0 25120 7 2 2 40077 65724
0 25121 5 1 1 65725
0 25122 7 1 2 25117 25121
0 25123 5 1 1 25122
0 25124 7 1 2 57782 52625
0 25125 7 1 2 25123 25124
0 25126 5 1 1 25125
0 25127 7 1 2 46141 25126
0 25128 7 1 2 25115 25127
0 25129 5 1 1 25128
0 25130 7 1 2 42662 25129
0 25131 5 1 1 25130
0 25132 7 1 2 25104 25131
0 25133 5 1 1 25132
0 25134 7 1 2 55946 53254
0 25135 5 1 1 25134
0 25136 7 1 2 58016 60886
0 25137 5 1 1 25136
0 25138 7 1 2 40444 51195
0 25139 7 1 2 25137 25138
0 25140 5 1 1 25139
0 25141 7 1 2 25135 25140
0 25142 5 1 1 25141
0 25143 7 1 2 41381 25142
0 25144 5 1 1 25143
0 25145 7 1 2 48161 54563
0 25146 5 1 1 25145
0 25147 7 1 2 25144 25146
0 25148 5 1 1 25147
0 25149 7 1 2 25148 52344
0 25150 5 1 1 25149
0 25151 7 1 2 50184 56282
0 25152 7 1 2 64633 25151
0 25153 5 1 1 25152
0 25154 7 1 2 25153 55822
0 25155 7 1 2 25150 25154
0 25156 5 1 1 25155
0 25157 7 1 2 48924 64863
0 25158 7 1 2 25156 25157
0 25159 7 1 2 25133 25158
0 25160 5 1 1 25159
0 25161 7 1 2 25050 25160
0 25162 7 1 2 24997 25161
0 25163 7 1 2 24902 25162
0 25164 7 1 2 24553 25163
0 25165 5 1 1 25164
0 25166 7 1 2 65224 25165
0 25167 5 1 1 25166
0 25168 7 1 2 45494 64840
0 25169 5 2 1 25168
0 25170 7 1 2 56275 65727
0 25171 5 1 1 25170
0 25172 7 1 2 25171 62840
0 25173 5 1 1 25172
0 25174 7 2 2 62141 64429
0 25175 7 1 2 41382 65729
0 25176 5 1 1 25175
0 25177 7 1 2 59956 51353
0 25178 5 1 1 25177
0 25179 7 1 2 25176 25178
0 25180 5 1 1 25179
0 25181 7 1 2 42406 25180
0 25182 5 1 1 25181
0 25183 7 1 2 48162 62029
0 25184 7 1 2 65730 25183
0 25185 5 1 1 25184
0 25186 7 1 2 25182 25185
0 25187 5 1 1 25186
0 25188 7 1 2 62846 25187
0 25189 5 1 1 25188
0 25190 7 1 2 25173 25189
0 25191 5 1 1 25190
0 25192 7 1 2 40445 25191
0 25193 5 1 1 25192
0 25194 7 1 2 62824 60547
0 25195 5 1 1 25194
0 25196 7 1 2 25193 25195
0 25197 5 1 1 25196
0 25198 7 1 2 42663 25197
0 25199 5 1 1 25198
0 25200 7 1 2 51924 62833
0 25201 5 1 1 25200
0 25202 7 1 2 25199 25201
0 25203 5 1 1 25202
0 25204 7 1 2 46142 25203
0 25205 5 1 1 25204
0 25206 7 3 2 53239 56183
0 25207 7 2 2 40446 60580
0 25208 7 1 2 51950 65734
0 25209 7 1 2 65731 25208
0 25210 7 1 2 62800 25209
0 25211 5 1 1 25210
0 25212 7 1 2 25205 25211
0 25213 5 1 1 25212
0 25214 7 1 2 47795 25213
0 25215 5 1 1 25214
0 25216 7 1 2 62801 60124
0 25217 5 1 1 25216
0 25218 7 1 2 53306 59055
0 25219 7 1 2 63686 25218
0 25220 5 1 1 25219
0 25221 7 1 2 25217 25220
0 25222 5 1 1 25221
0 25223 7 1 2 56009 25222
0 25224 5 1 1 25223
0 25225 7 2 2 50284 54920
0 25226 7 1 2 65593 65736
0 25227 7 1 2 59076 25226
0 25228 5 1 1 25227
0 25229 7 1 2 25224 25228
0 25230 5 1 1 25229
0 25231 7 1 2 60798 25230
0 25232 5 1 1 25231
0 25233 7 1 2 45964 65667
0 25234 5 1 1 25233
0 25235 7 1 2 42664 51875
0 25236 5 1 1 25235
0 25237 7 1 2 55476 25236
0 25238 5 1 1 25237
0 25239 7 1 2 40447 25238
0 25240 5 1 1 25239
0 25241 7 1 2 42407 25240
0 25242 7 1 2 25234 25241
0 25243 5 1 1 25242
0 25244 7 1 2 56241 50285
0 25245 5 2 1 25244
0 25246 7 1 2 64800 65738
0 25247 5 1 1 25246
0 25248 7 1 2 42665 25247
0 25249 5 1 1 25248
0 25250 7 1 2 45755 25249
0 25251 7 1 2 64798 25250
0 25252 5 1 1 25251
0 25253 7 1 2 46143 25252
0 25254 7 1 2 25243 25253
0 25255 5 1 1 25254
0 25256 7 1 2 40448 64180
0 25257 7 1 2 64841 25256
0 25258 5 1 1 25257
0 25259 7 1 2 22886 25258
0 25260 7 1 2 25255 25259
0 25261 5 1 1 25260
0 25262 7 1 2 62825 25261
0 25263 5 1 1 25262
0 25264 7 1 2 25232 25263
0 25265 7 1 2 25215 25264
0 25266 5 1 1 25265
0 25267 7 1 2 43010 25266
0 25268 5 1 1 25267
0 25269 7 1 2 58158 61031
0 25270 5 1 1 25269
0 25271 7 1 2 41251 55895
0 25272 5 1 1 25271
0 25273 7 1 2 47418 52656
0 25274 7 1 2 25272 25273
0 25275 5 1 1 25274
0 25276 7 1 2 54810 25275
0 25277 5 1 1 25276
0 25278 7 1 2 64815 25277
0 25279 5 1 1 25278
0 25280 7 1 2 25270 25279
0 25281 5 1 1 25280
0 25282 7 1 2 43569 25281
0 25283 5 1 1 25282
0 25284 7 1 2 58348 25283
0 25285 5 1 1 25284
0 25286 7 1 2 62826 65518
0 25287 7 1 2 25285 25286
0 25288 5 1 1 25287
0 25289 7 1 2 25268 25288
0 25290 5 1 1 25289
0 25291 7 1 2 59693 25290
0 25292 5 1 1 25291
0 25293 7 1 2 40449 51360
0 25294 5 1 1 25293
0 25295 7 1 2 25294 23334
0 25296 5 1 1 25295
0 25297 7 1 2 47796 25296
0 25298 5 1 1 25297
0 25299 7 1 2 53729 51599
0 25300 5 2 1 25299
0 25301 7 1 2 58103 65740
0 25302 7 1 2 25298 25301
0 25303 5 2 1 25302
0 25304 7 1 2 48125 65742
0 25305 5 2 1 25304
0 25306 7 2 2 48225 46899
0 25307 7 1 2 65746 64942
0 25308 5 1 1 25307
0 25309 7 1 2 65744 25308
0 25310 5 1 1 25309
0 25311 7 1 2 42666 25310
0 25312 5 1 1 25311
0 25313 7 1 2 48126 65669
0 25314 5 2 1 25313
0 25315 7 1 2 25312 65748
0 25316 5 1 1 25315
0 25317 7 1 2 42408 25316
0 25318 5 1 1 25317
0 25319 7 1 2 40450 47188
0 25320 5 1 1 25319
0 25321 7 1 2 44680 25320
0 25322 5 1 1 25321
0 25323 7 1 2 65673 25322
0 25324 5 1 1 25323
0 25325 7 1 2 43570 25324
0 25326 5 1 1 25325
0 25327 7 1 2 63035 49450
0 25328 5 1 1 25327
0 25329 7 1 2 45965 25328
0 25330 7 1 2 25326 25329
0 25331 5 1 1 25330
0 25332 7 1 2 50153 47573
0 25333 5 1 1 25332
0 25334 7 1 2 42667 65739
0 25335 7 1 2 25333 25334
0 25336 5 1 1 25335
0 25337 7 1 2 46144 25336
0 25338 7 1 2 25331 25337
0 25339 5 1 1 25338
0 25340 7 1 2 48706 53240
0 25341 7 1 2 58464 25340
0 25342 5 1 1 25341
0 25343 7 1 2 25339 25342
0 25344 5 1 1 25343
0 25345 7 1 2 51293 25344
0 25346 5 1 1 25345
0 25347 7 1 2 25318 25346
0 25348 5 1 1 25347
0 25349 7 1 2 59957 25348
0 25350 5 1 1 25349
0 25351 7 1 2 55479 56010
0 25352 5 1 1 25351
0 25353 7 2 2 47556 59860
0 25354 5 1 1 65750
0 25355 7 1 2 25352 25354
0 25356 5 1 1 25355
0 25357 7 1 2 40262 25356
0 25358 5 1 1 25357
0 25359 7 1 2 63031 59853
0 25360 5 1 1 25359
0 25361 7 1 2 25358 25360
0 25362 5 1 1 25361
0 25363 7 2 2 53647 25362
0 25364 7 1 2 64350 65752
0 25365 5 1 1 25364
0 25366 7 1 2 25350 25365
0 25367 5 1 1 25366
0 25368 7 1 2 41029 25367
0 25369 5 1 1 25368
0 25370 7 2 2 41815 65753
0 25371 7 1 2 63639 65754
0 25372 5 1 1 25371
0 25373 7 1 2 25369 25372
0 25374 5 1 1 25373
0 25375 7 1 2 53913 25374
0 25376 5 1 1 25375
0 25377 7 1 2 56888 59185
0 25378 7 1 2 65755 25377
0 25379 5 1 1 25378
0 25380 7 1 2 25376 25379
0 25381 5 1 1 25380
0 25382 7 1 2 43236 25381
0 25383 5 1 1 25382
0 25384 7 1 2 43404 61006
0 25385 5 1 1 25384
0 25386 7 1 2 65677 25385
0 25387 5 2 1 25386
0 25388 7 1 2 43571 65756
0 25389 5 1 1 25388
0 25390 7 1 2 581 25389
0 25391 5 1 1 25390
0 25392 7 1 2 56605 25391
0 25393 5 1 1 25392
0 25394 7 1 2 55931 54215
0 25395 5 1 1 25394
0 25396 7 1 2 25393 25395
0 25397 5 1 1 25396
0 25398 7 1 2 42668 25397
0 25399 5 1 1 25398
0 25400 7 1 2 49818 52277
0 25401 5 2 1 25400
0 25402 7 1 2 56269 57597
0 25403 7 1 2 65758 25402
0 25404 5 1 1 25403
0 25405 7 1 2 25399 25404
0 25406 5 1 1 25405
0 25407 7 1 2 59481 25406
0 25408 5 1 1 25407
0 25409 7 1 2 46718 65459
0 25410 5 1 1 25409
0 25411 7 3 2 45756 48127
0 25412 7 1 2 45966 65370
0 25413 7 2 2 49953 25412
0 25414 7 1 2 65760 65763
0 25415 5 1 1 25414
0 25416 7 1 2 25410 25415
0 25417 5 1 1 25416
0 25418 7 2 2 49827 25417
0 25419 7 1 2 61292 65765
0 25420 5 1 1 25419
0 25421 7 1 2 25408 25420
0 25422 5 1 1 25421
0 25423 7 1 2 53914 25422
0 25424 5 1 1 25423
0 25425 7 1 2 46508 62791
0 25426 7 1 2 65766 25425
0 25427 5 1 1 25426
0 25428 7 1 2 25424 25427
0 25429 5 1 1 25428
0 25430 7 1 2 43127 25429
0 25431 5 1 1 25430
0 25432 7 1 2 42669 62080
0 25433 7 1 2 49863 25432
0 25434 7 1 2 64439 25433
0 25435 5 1 1 25434
0 25436 7 3 2 45113 48616
0 25437 7 1 2 63689 65156
0 25438 7 1 2 65767 25437
0 25439 7 1 2 61302 25438
0 25440 5 1 1 25439
0 25441 7 1 2 25435 25440
0 25442 5 1 1 25441
0 25443 7 1 2 54216 25442
0 25444 5 1 1 25443
0 25445 7 5 2 54877 59509
0 25446 7 2 2 44681 65770
0 25447 7 1 2 50344 65768
0 25448 7 1 2 61308 25447
0 25449 7 1 2 65775 25448
0 25450 5 1 1 25449
0 25451 7 1 2 25444 25450
0 25452 5 1 1 25451
0 25453 7 1 2 48925 25452
0 25454 5 1 1 25453
0 25455 7 2 2 49308 62125
0 25456 7 1 2 53838 55334
0 25457 7 1 2 63074 25456
0 25458 7 1 2 65777 25457
0 25459 7 1 2 63326 25458
0 25460 5 1 1 25459
0 25461 7 1 2 25454 25460
0 25462 5 1 1 25461
0 25463 7 1 2 59975 25462
0 25464 5 1 1 25463
0 25465 7 1 2 25431 25464
0 25466 5 1 1 25465
0 25467 7 1 2 42152 25466
0 25468 5 1 1 25467
0 25469 7 2 2 40451 63492
0 25470 7 3 2 57209 58608
0 25471 7 1 2 59856 65781
0 25472 7 1 2 62802 25471
0 25473 7 1 2 65779 25472
0 25474 5 1 1 25473
0 25475 7 1 2 25468 25474
0 25476 7 1 2 25383 25475
0 25477 5 1 1 25476
0 25478 7 1 2 45162 25477
0 25479 5 1 1 25478
0 25480 7 1 2 25292 25479
0 25481 5 1 1 25480
0 25482 7 1 2 43926 25481
0 25483 5 1 1 25482
0 25484 7 1 2 59792 64362
0 25485 5 1 1 25484
0 25486 7 1 2 47346 65386
0 25487 5 1 1 25486
0 25488 7 1 2 45757 51378
0 25489 5 1 1 25488
0 25490 7 1 2 25487 25489
0 25491 5 1 1 25490
0 25492 7 1 2 25491 50989
0 25493 5 1 1 25492
0 25494 7 1 2 25485 25493
0 25495 5 2 1 25494
0 25496 7 12 2 43237 60083
0 25497 7 1 2 65786 60715
0 25498 5 1 1 25497
0 25499 7 1 2 45967 48926
0 25500 7 1 2 65411 25499
0 25501 5 1 1 25500
0 25502 7 1 2 25498 25501
0 25503 5 1 1 25502
0 25504 7 1 2 65784 25503
0 25505 5 1 1 25504
0 25506 7 1 2 48175 64918
0 25507 5 2 1 25506
0 25508 7 1 2 60111 65798
0 25509 5 1 1 25508
0 25510 7 3 2 51744 60165
0 25511 7 1 2 42409 65800
0 25512 5 1 1 25511
0 25513 7 1 2 25509 25512
0 25514 5 1 1 25513
0 25515 7 1 2 41383 25514
0 25516 5 1 1 25515
0 25517 7 4 2 41136 50879
0 25518 7 1 2 60134 56817
0 25519 7 1 2 65803 25518
0 25520 5 1 1 25519
0 25521 7 1 2 25516 25520
0 25522 5 1 1 25521
0 25523 7 1 2 47797 25522
0 25524 5 1 1 25523
0 25525 7 2 2 44682 60183
0 25526 7 3 2 45163 65807
0 25527 5 1 1 65809
0 25528 7 1 2 50487 65810
0 25529 5 1 1 25528
0 25530 7 1 2 41845 61896
0 25531 7 1 2 60601 25530
0 25532 5 1 1 25531
0 25533 7 1 2 25529 25532
0 25534 5 1 1 25533
0 25535 7 1 2 46758 25534
0 25536 5 1 1 25535
0 25537 7 2 2 46961 56818
0 25538 7 1 2 65281 65812
0 25539 5 1 1 25538
0 25540 7 2 2 47167 57857
0 25541 7 1 2 61778 65429
0 25542 7 1 2 65814 25541
0 25543 5 1 1 25542
0 25544 7 1 2 25539 25543
0 25545 7 1 2 25536 25544
0 25546 5 1 1 25545
0 25547 7 1 2 47593 25546
0 25548 5 1 1 25547
0 25549 7 1 2 25524 25548
0 25550 5 1 1 25549
0 25551 7 1 2 40078 25550
0 25552 5 1 1 25551
0 25553 7 1 2 56283 65290
0 25554 5 2 1 25553
0 25555 7 1 2 44683 56184
0 25556 5 1 1 25555
0 25557 7 1 2 50682 25556
0 25558 5 2 1 25557
0 25559 7 1 2 60184 64051
0 25560 7 1 2 65818 25559
0 25561 5 1 1 25560
0 25562 7 1 2 65816 25561
0 25563 5 1 1 25562
0 25564 7 1 2 41252 25563
0 25565 5 1 1 25564
0 25566 7 2 2 48163 65404
0 25567 7 1 2 64787 65820
0 25568 5 1 1 25567
0 25569 7 1 2 25565 25568
0 25570 5 1 1 25569
0 25571 7 1 2 41137 25570
0 25572 5 1 1 25571
0 25573 7 1 2 47025 57858
0 25574 7 1 2 64649 25573
0 25575 7 1 2 64788 25574
0 25576 5 1 1 25575
0 25577 7 1 2 25572 25576
0 25578 5 1 1 25577
0 25579 7 1 2 40263 25578
0 25580 5 1 1 25579
0 25581 7 2 2 62257 61779
0 25582 7 1 2 41253 65822
0 25583 7 1 2 65821 25582
0 25584 5 1 1 25583
0 25585 7 1 2 25580 25584
0 25586 7 1 2 25552 25585
0 25587 5 1 1 25586
0 25588 7 1 2 61887 25587
0 25589 5 1 1 25588
0 25590 7 2 2 59569 62100
0 25591 5 1 1 65824
0 25592 7 1 2 40079 65825
0 25593 5 1 1 25592
0 25594 7 2 2 47286 51581
0 25595 5 1 1 65826
0 25596 7 2 2 60208 60102
0 25597 5 1 1 65828
0 25598 7 1 2 60173 25597
0 25599 5 1 1 25598
0 25600 7 1 2 65827 25599
0 25601 5 1 1 25600
0 25602 7 3 2 65405 64789
0 25603 5 1 1 65830
0 25604 7 1 2 65831 51125
0 25605 5 1 1 25604
0 25606 7 1 2 25601 25605
0 25607 5 1 1 25606
0 25608 7 1 2 42410 25607
0 25609 5 1 1 25608
0 25610 7 1 2 25593 25609
0 25611 7 1 2 65282 65333
0 25612 5 1 1 25611
0 25613 7 2 2 40264 60112
0 25614 5 2 1 65833
0 25615 7 1 2 41254 65834
0 25616 5 1 1 25615
0 25617 7 1 2 25612 25616
0 25618 5 1 1 25617
0 25619 7 1 2 56284 25618
0 25620 5 1 1 25619
0 25621 7 1 2 64999 60113
0 25622 5 1 1 25621
0 25623 7 2 2 47976 59632
0 25624 7 1 2 65694 65837
0 25625 5 1 1 25624
0 25626 7 1 2 65817 25625
0 25627 7 1 2 25622 25626
0 25628 5 1 1 25627
0 25629 7 1 2 47478 25628
0 25630 5 1 1 25629
0 25631 7 1 2 25620 25630
0 25632 7 1 2 25610 25631
0 25633 5 1 1 25632
0 25634 7 1 2 61888 25633
0 25635 5 1 1 25634
0 25636 7 3 2 64185 57762
0 25637 5 1 1 65839
0 25638 7 4 2 45164 62261
0 25639 7 1 2 46422 65842
0 25640 5 1 1 25639
0 25641 7 2 2 60174 25640
0 25642 5 2 1 65846
0 25643 7 1 2 40080 65848
0 25644 5 1 1 25643
0 25645 7 1 2 25637 25644
0 25646 5 2 1 25645
0 25647 7 1 2 47798 65850
0 25648 5 1 1 25647
0 25649 7 2 2 41763 65406
0 25650 7 3 2 40265 54633
0 25651 7 1 2 65852 65854
0 25652 5 1 1 25651
0 25653 7 1 2 25648 25652
0 25654 5 1 1 25653
0 25655 7 1 2 45324 25654
0 25656 5 1 1 25655
0 25657 7 1 2 47479 60114
0 25658 5 1 1 25657
0 25659 7 1 2 60175 25658
0 25660 5 1 1 25659
0 25661 7 1 2 47594 25660
0 25662 5 1 1 25661
0 25663 7 1 2 65832 58691
0 25664 5 1 1 25663
0 25665 7 1 2 43128 60127
0 25666 7 1 2 57763 25665
0 25667 7 1 2 52551 25666
0 25668 5 1 1 25667
0 25669 7 1 2 25664 25668
0 25670 5 1 1 25669
0 25671 7 1 2 51925 25670
0 25672 5 1 1 25671
0 25673 7 1 2 25662 25672
0 25674 7 1 2 25656 25673
0 25675 5 1 1 25674
0 25676 7 1 2 43238 25675
0 25677 5 1 1 25676
0 25678 7 2 2 49293 57764
0 25679 7 5 2 62708 63380
0 25680 7 1 2 45165 65859
0 25681 7 1 2 65857 25680
0 25682 5 1 1 25681
0 25683 7 1 2 25677 25682
0 25684 5 1 1 25683
0 25685 7 1 2 65701 25684
0 25686 5 1 1 25685
0 25687 7 1 2 25635 25686
0 25688 5 1 1 25687
0 25689 7 1 2 40452 25688
0 25690 5 1 1 25689
0 25691 7 1 2 25589 25690
0 25692 5 1 1 25691
0 25693 7 1 2 55078 25692
0 25694 5 1 1 25693
0 25695 7 2 2 41384 61094
0 25696 5 2 1 65864
0 25697 7 2 2 41138 61100
0 25698 7 2 2 40081 65868
0 25699 5 1 1 65870
0 25700 7 1 2 40266 65871
0 25701 5 1 1 25700
0 25702 7 1 2 65866 25701
0 25703 5 1 1 25702
0 25704 7 1 2 47124 25703
0 25705 5 1 1 25704
0 25706 7 1 2 65855 58605
0 25707 5 1 1 25706
0 25708 7 1 2 12710 25699
0 25709 5 1 1 25708
0 25710 7 1 2 47996 25709
0 25711 5 1 1 25710
0 25712 7 1 2 25707 25711
0 25713 7 1 2 25705 25712
0 25714 5 1 1 25713
0 25715 7 1 2 42411 25714
0 25716 5 1 1 25715
0 25717 7 2 2 53343 57033
0 25718 5 2 1 65872
0 25719 7 1 2 51964 65873
0 25720 5 1 1 25719
0 25721 7 1 2 47799 53992
0 25722 5 1 1 25721
0 25723 7 1 2 13110 25722
0 25724 5 1 1 25723
0 25725 7 1 2 56285 25724
0 25726 5 1 1 25725
0 25727 7 1 2 25720 25726
0 25728 7 1 2 25716 25727
0 25729 5 1 1 25728
0 25730 7 1 2 40453 25729
0 25731 5 1 1 25730
0 25732 7 1 2 54175 61223
0 25733 5 2 1 25732
0 25734 7 1 2 41385 61902
0 25735 5 1 1 25734
0 25736 7 1 2 65876 25735
0 25737 5 1 1 25736
0 25738 7 1 2 46759 25737
0 25739 5 1 1 25738
0 25740 7 1 2 53915 65813
0 25741 5 1 1 25740
0 25742 7 1 2 60602 65815
0 25743 5 1 1 25742
0 25744 7 1 2 25741 25743
0 25745 7 1 2 25739 25744
0 25746 5 1 1 25745
0 25747 7 1 2 60772 25746
0 25748 5 1 1 25747
0 25749 7 1 2 65295 65865
0 25750 5 1 1 25749
0 25751 7 1 2 56286 57055
0 25752 5 1 1 25751
0 25753 7 1 2 65877 25752
0 25754 5 1 1 25753
0 25755 7 1 2 45325 25754
0 25756 5 1 1 25755
0 25757 7 2 2 50750 54584
0 25758 5 1 1 65878
0 25759 7 1 2 50591 65879
0 25760 5 1 1 25759
0 25761 7 1 2 25756 25760
0 25762 5 1 1 25761
0 25763 7 1 2 50231 25762
0 25764 5 1 1 25763
0 25765 7 1 2 25750 25764
0 25766 7 1 2 25748 25765
0 25767 5 1 1 25766
0 25768 7 1 2 40267 25767
0 25769 5 1 1 25768
0 25770 7 4 2 47480 54093
0 25771 5 1 1 65880
0 25772 7 1 2 56306 65881
0 25773 5 1 1 25772
0 25774 7 1 2 65867 21176
0 25775 5 1 1 25774
0 25776 7 1 2 60545 56189
0 25777 7 1 2 25775 25776
0 25778 5 1 1 25777
0 25779 7 1 2 25773 25778
0 25780 7 1 2 25769 25779
0 25781 5 1 1 25780
0 25782 7 1 2 47800 25781
0 25783 5 1 1 25782
0 25784 7 1 2 25731 25783
0 25785 5 1 1 25784
0 25786 7 1 2 45968 25785
0 25787 5 1 1 25786
0 25788 7 3 2 50445 53993
0 25789 5 2 1 65884
0 25790 7 1 2 64263 65885
0 25791 5 1 1 25790
0 25792 7 1 2 56287 60235
0 25793 5 1 1 25792
0 25794 7 1 2 25791 25793
0 25795 5 1 1 25794
0 25796 7 1 2 47801 25795
0 25797 5 1 1 25796
0 25798 7 1 2 52184 62001
0 25799 5 1 1 25798
0 25800 7 1 2 25799 9901
0 25801 5 1 1 25800
0 25802 7 1 2 45758 25801
0 25803 5 1 1 25802
0 25804 7 1 2 62003 60640
0 25805 5 2 1 25804
0 25806 7 2 2 42412 51582
0 25807 5 2 1 65891
0 25808 7 1 2 45969 65892
0 25809 7 1 2 65889 25808
0 25810 5 1 1 25809
0 25811 7 1 2 25803 25810
0 25812 7 1 2 25797 25811
0 25813 5 1 1 25812
0 25814 7 1 2 47481 25813
0 25815 5 1 1 25814
0 25816 7 1 2 61095 62484
0 25817 5 1 1 25816
0 25818 7 1 2 54687 65856
0 25819 5 1 1 25818
0 25820 7 1 2 25817 25819
0 25821 5 1 1 25820
0 25822 7 1 2 52472 25821
0 25823 5 1 1 25822
0 25824 7 1 2 25815 25823
0 25825 5 1 1 25824
0 25826 7 1 2 40454 25825
0 25827 5 1 1 25826
0 25828 7 1 2 25787 25827
0 25829 5 1 1 25828
0 25830 7 1 2 65787 25829
0 25831 5 1 1 25830
0 25832 7 3 2 40455 64650
0 25833 7 1 2 64264 65895
0 25834 7 1 2 61554 63174
0 25835 7 1 2 25833 25834
0 25836 5 1 1 25835
0 25837 7 1 2 42859 25836
0 25838 7 1 2 25831 25837
0 25839 7 1 2 25694 25838
0 25840 5 1 1 25839
0 25841 7 1 2 48184 65728
0 25842 5 2 1 25841
0 25843 7 1 2 60115 65898
0 25844 5 1 1 25843
0 25845 7 1 2 49298 59570
0 25846 7 1 2 63575 25845
0 25847 5 1 1 25846
0 25848 7 1 2 25844 25847
0 25849 5 1 1 25848
0 25850 7 1 2 44684 25849
0 25851 5 1 1 25850
0 25852 7 1 2 55991 55687
0 25853 5 1 1 25852
0 25854 7 1 2 24793 55973
0 25855 7 1 2 25853 25854
0 25856 5 1 1 25855
0 25857 7 1 2 60166 25856
0 25858 5 1 1 25857
0 25859 7 1 2 25851 25858
0 25860 5 1 1 25859
0 25861 7 1 2 43737 25860
0 25862 5 1 1 25861
0 25863 7 1 2 48185 53696
0 25864 5 2 1 25863
0 25865 7 1 2 43129 55150
0 25866 7 2 2 65900 25865
0 25867 7 1 2 60135 65902
0 25868 5 1 1 25867
0 25869 7 2 2 63725 65339
0 25870 7 1 2 65430 59080
0 25871 7 1 2 65904 25870
0 25872 5 1 1 25871
0 25873 7 1 2 25868 25872
0 25874 7 1 2 25862 25873
0 25875 5 1 1 25874
0 25876 7 1 2 43239 25875
0 25877 5 1 1 25876
0 25878 7 1 2 56270 65380
0 25879 7 1 2 63576 25878
0 25880 7 1 2 54675 25879
0 25881 7 1 2 65375 25880
0 25882 5 1 1 25881
0 25883 7 1 2 25877 25882
0 25884 5 1 1 25883
0 25885 7 1 2 42670 25884
0 25886 5 1 1 25885
0 25887 7 1 2 42153 65757
0 25888 5 1 1 25887
0 25889 7 1 2 49451 56259
0 25890 5 1 1 25889
0 25891 7 1 2 25888 25890
0 25892 5 1 1 25891
0 25893 7 1 2 43572 25892
0 25894 5 1 1 25893
0 25895 7 1 2 25894 58349
0 25896 5 3 1 25895
0 25897 7 2 2 48927 65390
0 25898 7 1 2 65909 64442
0 25899 7 1 2 65906 25898
0 25900 5 1 1 25899
0 25901 7 1 2 25886 25900
0 25902 5 1 1 25901
0 25903 7 1 2 55079 25902
0 25904 5 1 1 25903
0 25905 7 1 2 53916 65903
0 25906 5 1 1 25905
0 25907 7 1 2 65905 62161
0 25908 5 1 1 25907
0 25909 7 1 2 25906 25908
0 25910 5 1 1 25909
0 25911 7 1 2 65788 25910
0 25912 5 1 1 25911
0 25913 7 1 2 48000 52270
0 25914 5 1 1 25913
0 25915 7 1 2 65789 25914
0 25916 5 1 1 25915
0 25917 7 2 2 57649 47736
0 25918 7 1 2 65381 65911
0 25919 7 1 2 65376 25918
0 25920 5 1 1 25919
0 25921 7 1 2 25916 25920
0 25922 5 1 1 25921
0 25923 7 1 2 43405 25922
0 25924 5 1 1 25923
0 25925 7 1 2 47940 48013
0 25926 5 2 1 25925
0 25927 7 1 2 65913 65790
0 25928 5 1 1 25927
0 25929 7 1 2 25924 25928
0 25930 5 1 1 25929
0 25931 7 1 2 45759 25930
0 25932 5 1 1 25931
0 25933 7 1 2 49299 50592
0 25934 7 1 2 65791 25933
0 25935 5 1 1 25934
0 25936 7 1 2 25932 25935
0 25937 5 1 1 25936
0 25938 7 1 2 53994 25937
0 25939 5 1 1 25938
0 25940 7 1 2 59031 65792
0 25941 7 1 2 65899 25940
0 25942 5 1 1 25941
0 25943 7 1 2 25939 25942
0 25944 5 1 1 25943
0 25945 7 1 2 43738 25944
0 25946 5 1 1 25945
0 25947 7 1 2 25912 25946
0 25948 5 1 1 25947
0 25949 7 1 2 42671 25948
0 25950 5 1 1 25949
0 25951 7 2 2 45970 57034
0 25952 7 2 2 61315 65915
0 25953 7 1 2 41764 60084
0 25954 7 1 2 65917 25953
0 25955 7 1 2 65907 25954
0 25956 5 1 1 25955
0 25957 7 1 2 46145 25956
0 25958 7 1 2 25950 25957
0 25959 7 1 2 25904 25958
0 25960 5 1 1 25959
0 25961 7 1 2 40653 25960
0 25962 7 1 2 25840 25961
0 25963 5 1 1 25962
0 25964 7 1 2 25505 25963
0 25965 5 1 1 25964
0 25966 7 1 2 43011 25965
0 25967 5 1 1 25966
0 25968 7 1 2 25483 25967
0 25969 5 1 1 25968
0 25970 7 1 2 44814 25969
0 25971 5 1 1 25970
0 25972 7 1 2 56697 62970
0 25973 5 1 1 25972
0 25974 7 3 2 48343 54433
0 25975 5 1 1 65919
0 25976 7 1 2 55508 25975
0 25977 5 1 1 25976
0 25978 7 1 2 54229 25977
0 25979 5 2 1 25978
0 25980 7 1 2 51926 62965
0 25981 5 1 1 25980
0 25982 7 1 2 43739 25981
0 25983 5 1 1 25982
0 25984 7 1 2 42860 25983
0 25985 7 1 2 65706 25984
0 25986 5 1 1 25985
0 25987 7 1 2 65922 25986
0 25988 5 1 1 25987
0 25989 7 1 2 43927 25988
0 25990 5 1 1 25989
0 25991 7 2 2 40456 63909
0 25992 7 1 2 42861 65924
0 25993 7 1 2 65301 25992
0 25994 5 1 1 25993
0 25995 7 1 2 25990 25994
0 25996 5 1 1 25995
0 25997 7 1 2 53648 25996
0 25998 5 1 1 25997
0 25999 7 1 2 25973 25998
0 26000 5 1 1 25999
0 26001 7 1 2 53917 26000
0 26002 5 1 1 26001
0 26003 7 1 2 56899 64137
0 26004 7 1 2 60610 26003
0 26005 5 1 1 26004
0 26006 7 1 2 26002 26005
0 26007 5 1 1 26006
0 26008 7 1 2 40268 26007
0 26009 5 1 1 26008
0 26010 7 1 2 53099 49836
0 26011 7 1 2 65015 26010
0 26012 5 1 1 26011
0 26013 7 1 2 24655 26012
0 26014 5 1 1 26013
0 26015 7 1 2 42413 26014
0 26016 5 1 1 26015
0 26017 7 1 2 65619 60802
0 26018 5 1 1 26017
0 26019 7 1 2 26016 26018
0 26020 5 1 1 26019
0 26021 7 1 2 53918 63654
0 26022 7 1 2 26020 26021
0 26023 5 1 1 26022
0 26024 7 1 2 26009 26023
0 26025 5 1 1 26024
0 26026 7 1 2 45166 26025
0 26027 5 1 1 26026
0 26028 7 1 2 54833 63914
0 26029 5 7 1 26028
0 26030 7 2 2 65690 65926
0 26031 7 1 2 57574 48585
0 26032 7 1 2 65910 26031
0 26033 7 1 2 65933 26032
0 26034 5 1 1 26033
0 26035 7 1 2 26027 26034
0 26036 5 1 1 26035
0 26037 7 1 2 55080 26036
0 26038 5 1 1 26037
0 26039 7 3 2 42862 56288
0 26040 7 1 2 56802 65935
0 26041 5 1 1 26040
0 26042 7 1 2 56612 58753
0 26043 5 1 1 26042
0 26044 7 1 2 26041 26043
0 26045 5 1 1 26044
0 26046 7 1 2 47802 26045
0 26047 5 1 1 26046
0 26048 7 1 2 54230 63146
0 26049 5 1 1 26048
0 26050 7 2 2 43928 52005
0 26051 5 2 1 65938
0 26052 7 1 2 55948 65940
0 26053 5 2 1 26052
0 26054 7 1 2 42863 58209
0 26055 7 1 2 65942 26054
0 26056 5 1 1 26055
0 26057 7 1 2 26049 26056
0 26058 5 1 1 26057
0 26059 7 1 2 45495 26058
0 26060 5 1 1 26059
0 26061 7 1 2 26047 26060
0 26062 5 1 1 26061
0 26063 7 1 2 42672 26062
0 26064 5 1 1 26063
0 26065 7 1 2 42414 61449
0 26066 5 1 1 26065
0 26067 7 1 2 54231 55503
0 26068 5 1 1 26067
0 26069 7 1 2 26066 26068
0 26070 5 1 1 26069
0 26071 7 1 2 55250 55765
0 26072 7 1 2 26070 26071
0 26073 5 1 1 26072
0 26074 7 1 2 26064 26073
0 26075 5 1 1 26074
0 26076 7 1 2 54176 26075
0 26077 5 1 1 26076
0 26078 7 1 2 53919 57575
0 26079 7 1 2 56093 26078
0 26080 7 1 2 65934 26079
0 26081 5 1 1 26080
0 26082 7 1 2 26077 26081
0 26083 5 1 1 26082
0 26084 7 1 2 43012 26083
0 26085 5 1 1 26084
0 26086 7 1 2 56951 55421
0 26087 7 1 2 60611 26086
0 26088 5 1 1 26087
0 26089 7 1 2 26085 26088
0 26090 5 1 1 26089
0 26091 7 1 2 60085 26090
0 26092 5 1 1 26091
0 26093 7 2 2 50286 59726
0 26094 7 1 2 58986 57610
0 26095 7 1 2 65944 26094
0 26096 7 1 2 56576 26095
0 26097 5 1 1 26096
0 26098 7 1 2 26092 26097
0 26099 7 1 2 26038 26098
0 26100 5 1 1 26099
0 26101 7 1 2 46760 26100
0 26102 5 1 1 26101
0 26103 7 1 2 60498 65849
0 26104 5 1 1 26103
0 26105 7 1 2 41976 65801
0 26106 5 1 1 26105
0 26107 7 1 2 26104 26106
0 26108 5 1 1 26107
0 26109 7 1 2 40082 26108
0 26110 5 1 1 26109
0 26111 7 2 2 57455 62092
0 26112 7 1 2 46952 59633
0 26113 7 1 2 65946 26112
0 26114 5 1 1 26113
0 26115 7 1 2 26110 26114
0 26116 5 1 1 26115
0 26117 7 1 2 53321 26116
0 26118 5 1 1 26117
0 26119 7 1 2 65602 60116
0 26120 5 1 1 26119
0 26121 7 1 2 65597 60167
0 26122 5 1 1 26121
0 26123 7 1 2 26120 26122
0 26124 5 1 1 26123
0 26125 7 1 2 40083 26124
0 26126 5 1 1 26125
0 26127 7 1 2 40269 52512
0 26128 7 1 2 65600 26127
0 26129 7 1 2 65840 26128
0 26130 5 1 1 26129
0 26131 7 1 2 60176 65835
0 26132 5 1 1 26131
0 26133 7 1 2 40654 53558
0 26134 7 1 2 26132 26133
0 26135 5 1 1 26134
0 26136 7 1 2 26130 26135
0 26137 7 1 2 26126 26136
0 26138 5 1 1 26137
0 26139 7 1 2 40457 26138
0 26140 5 1 1 26139
0 26141 7 1 2 26118 26140
0 26142 5 1 1 26141
0 26143 7 1 2 45760 26142
0 26144 5 1 1 26143
0 26145 7 2 2 53433 56545
0 26146 7 1 2 52328 65851
0 26147 5 1 1 26146
0 26148 7 1 2 40084 65802
0 26149 5 1 1 26148
0 26150 7 1 2 48640 60117
0 26151 5 1 1 26150
0 26152 7 1 2 60177 26151
0 26153 5 1 1 26152
0 26154 7 1 2 40458 26153
0 26155 5 1 1 26154
0 26156 7 1 2 26149 26155
0 26157 7 1 2 26147 26156
0 26158 5 1 1 26157
0 26159 7 1 2 65948 26158
0 26160 5 1 1 26159
0 26161 7 1 2 26144 26160
0 26162 5 1 1 26161
0 26163 7 1 2 42673 26162
0 26164 5 1 1 26163
0 26165 7 1 2 43573 60142
0 26166 5 1 1 26165
0 26167 7 1 2 26166 25527
0 26168 5 1 1 26167
0 26169 7 1 2 43740 26168
0 26170 5 1 1 26169
0 26171 7 1 2 44524 65811
0 26172 5 1 1 26171
0 26173 7 1 2 48008 60143
0 26174 5 1 1 26173
0 26175 7 1 2 26172 26174
0 26176 5 1 1 26175
0 26177 7 1 2 43574 26176
0 26178 5 1 1 26177
0 26179 7 1 2 26170 26178
0 26180 5 1 1 26179
0 26181 7 1 2 44428 26180
0 26182 5 1 1 26181
0 26183 7 4 2 43130 48009
0 26184 7 2 2 60128 59244
0 26185 7 1 2 65950 65954
0 26186 5 1 1 26185
0 26187 7 1 2 26182 26186
0 26188 5 1 1 26187
0 26189 7 1 2 43406 26188
0 26190 5 1 1 26189
0 26191 7 2 2 43131 65914
0 26192 7 1 2 65956 65955
0 26193 5 1 1 26192
0 26194 7 1 2 40655 26193
0 26195 7 1 2 26190 26194
0 26196 5 1 1 26195
0 26197 7 1 2 40270 65291
0 26198 5 1 1 26197
0 26199 7 1 2 26198 25603
0 26200 5 1 1 26199
0 26201 7 1 2 41139 26200
0 26202 5 1 1 26201
0 26203 7 1 2 65847 65836
0 26204 5 1 1 26203
0 26205 7 1 2 40459 26204
0 26206 5 1 1 26205
0 26207 7 1 2 26202 26206
0 26208 5 1 1 26207
0 26209 7 1 2 41255 26208
0 26210 5 1 1 26209
0 26211 7 1 2 49542 65407
0 26212 7 1 2 63399 26211
0 26213 5 1 1 26212
0 26214 7 1 2 26210 26213
0 26215 5 1 1 26214
0 26216 7 1 2 42154 26215
0 26217 5 1 1 26216
0 26218 7 1 2 58798 60103
0 26219 7 1 2 49925 26218
0 26220 5 1 1 26219
0 26221 7 1 2 40460 46962
0 26222 5 1 1 26221
0 26223 7 1 2 41256 55628
0 26224 5 1 1 26223
0 26225 7 1 2 26222 26224
0 26226 5 2 1 26225
0 26227 7 1 2 60168 65958
0 26228 5 1 1 26227
0 26229 7 1 2 26220 26228
0 26230 5 1 1 26229
0 26231 7 1 2 40085 26230
0 26232 5 1 1 26231
0 26233 7 1 2 59727 63091
0 26234 7 1 2 65808 26233
0 26235 5 1 1 26234
0 26236 7 1 2 43929 26235
0 26237 7 1 2 26232 26236
0 26238 7 1 2 26217 26237
0 26239 5 1 1 26238
0 26240 7 1 2 26196 26239
0 26241 5 1 1 26240
0 26242 7 1 2 45761 26241
0 26243 5 1 1 26242
0 26244 7 1 2 65634 65256
0 26245 5 1 1 26244
0 26246 7 1 2 65630 50778
0 26247 5 1 1 26246
0 26248 7 1 2 26245 26247
0 26249 5 2 1 26248
0 26250 7 1 2 60169 65960
0 26251 5 1 1 26250
0 26252 7 3 2 47595 62516
0 26253 5 5 1 65962
0 26254 7 1 2 41386 65963
0 26255 5 1 1 26254
0 26256 7 6 2 40656 44429
0 26257 7 1 2 55797 65970
0 26258 7 1 2 55909 26257
0 26259 5 1 1 26258
0 26260 7 1 2 26255 26259
0 26261 5 2 1 26260
0 26262 7 1 2 65976 60118
0 26263 5 1 1 26262
0 26264 7 1 2 42415 26263
0 26265 7 1 2 26251 26264
0 26266 5 1 1 26265
0 26267 7 1 2 45971 26266
0 26268 7 1 2 26243 26267
0 26269 5 1 1 26268
0 26270 7 1 2 42864 26269
0 26271 7 1 2 26164 26270
0 26272 5 1 1 26271
0 26273 7 1 2 44685 65259
0 26274 5 1 1 26273
0 26275 7 1 2 65253 26274
0 26276 5 1 1 26275
0 26277 7 1 2 60170 26276
0 26278 5 1 1 26277
0 26279 7 1 2 42416 60209
0 26280 7 2 2 65011 26279
0 26281 7 1 2 65978 65843
0 26282 5 1 1 26281
0 26283 7 1 2 52356 60190
0 26284 5 1 1 26283
0 26285 7 1 2 26282 26284
0 26286 5 1 1 26285
0 26287 7 1 2 44686 26286
0 26288 5 1 1 26287
0 26289 7 1 2 26278 26288
0 26290 5 1 1 26289
0 26291 7 1 2 42674 26290
0 26292 5 1 1 26291
0 26293 7 2 2 63556 65908
0 26294 5 1 1 65980
0 26295 7 1 2 65981 65283
0 26296 5 1 1 26295
0 26297 7 1 2 26292 26296
0 26298 5 1 1 26297
0 26299 7 1 2 43930 26298
0 26300 5 1 1 26299
0 26301 7 1 2 64958 65284
0 26302 5 1 1 26301
0 26303 7 1 2 46146 26302
0 26304 7 1 2 26300 26303
0 26305 5 1 1 26304
0 26306 7 1 2 43013 26305
0 26307 7 1 2 26272 26306
0 26308 5 1 1 26307
0 26309 7 1 2 45167 57588
0 26310 7 1 2 63346 26309
0 26311 7 1 2 64138 62206
0 26312 7 1 2 65737 26311
0 26313 7 1 2 26310 26312
0 26314 5 1 1 26313
0 26315 7 1 2 26308 26314
0 26316 5 1 1 26315
0 26317 7 1 2 55081 26316
0 26318 5 1 1 26317
0 26319 7 1 2 65598 57056
0 26320 5 1 1 26319
0 26321 7 1 2 65603 54094
0 26322 5 1 1 26321
0 26323 7 1 2 26320 26322
0 26324 5 1 1 26323
0 26325 7 1 2 40086 26324
0 26326 5 1 1 26325
0 26327 7 2 2 62709 65823
0 26328 5 1 1 65982
0 26329 7 1 2 45496 55766
0 26330 7 1 2 65983 26329
0 26331 5 1 1 26330
0 26332 7 2 2 48928 61519
0 26333 5 1 1 65984
0 26334 7 1 2 26328 26333
0 26335 5 1 1 26334
0 26336 7 1 2 40271 26335
0 26337 5 1 1 26336
0 26338 7 1 2 26337 20945
0 26339 5 1 1 26338
0 26340 7 1 2 53559 26339
0 26341 5 1 1 26340
0 26342 7 1 2 26331 26341
0 26343 7 1 2 26326 26342
0 26344 5 1 1 26343
0 26345 7 1 2 40461 26344
0 26346 5 1 1 26345
0 26347 7 1 2 53995 65804
0 26348 5 1 1 26347
0 26349 7 2 2 52329 57745
0 26350 5 1 1 65986
0 26351 7 1 2 42155 65987
0 26352 5 1 1 26351
0 26353 7 1 2 26348 26352
0 26354 5 1 1 26353
0 26355 7 1 2 40087 26354
0 26356 5 1 1 26355
0 26357 7 1 2 60571 60616
0 26358 5 1 1 26357
0 26359 7 1 2 26356 26358
0 26360 5 1 1 26359
0 26361 7 1 2 53322 26360
0 26362 5 1 1 26361
0 26363 7 1 2 26346 26362
0 26364 5 1 1 26363
0 26365 7 1 2 45762 26364
0 26366 5 1 1 26365
0 26367 7 1 2 62258 64871
0 26368 5 1 1 26367
0 26369 7 1 2 26350 26368
0 26370 5 1 1 26369
0 26371 7 1 2 40088 26370
0 26372 5 1 1 26371
0 26373 7 1 2 52255 57057
0 26374 5 1 1 26373
0 26375 7 4 2 56889 54078
0 26376 5 1 1 65988
0 26377 7 1 2 48641 65989
0 26378 5 1 1 26377
0 26379 7 1 2 26374 26378
0 26380 7 1 2 26372 26379
0 26381 5 1 1 26380
0 26382 7 1 2 65949 26381
0 26383 5 1 1 26382
0 26384 7 1 2 26366 26383
0 26385 5 1 1 26384
0 26386 7 1 2 42675 26385
0 26387 5 1 1 26386
0 26388 7 1 2 60588 65951
0 26389 5 1 1 26388
0 26390 7 1 2 47935 54177
0 26391 5 1 1 26390
0 26392 7 1 2 26389 26391
0 26393 5 1 1 26392
0 26394 7 1 2 43575 26393
0 26395 5 1 1 26394
0 26396 7 1 2 55139 57058
0 26397 5 1 1 26396
0 26398 7 1 2 7731 26397
0 26399 5 1 1 26398
0 26400 7 1 2 43741 26399
0 26401 5 1 1 26400
0 26402 7 1 2 26395 26401
0 26403 5 1 1 26402
0 26404 7 1 2 44430 26403
0 26405 5 1 1 26404
0 26406 7 4 2 41765 56053
0 26407 7 1 2 65992 65952
0 26408 5 1 1 26407
0 26409 7 1 2 26405 26408
0 26410 5 1 1 26409
0 26411 7 1 2 43407 26410
0 26412 5 1 1 26411
0 26413 7 1 2 65993 65957
0 26414 5 1 1 26413
0 26415 7 1 2 40657 26414
0 26416 7 1 2 26412 26415
0 26417 5 1 1 26416
0 26418 7 1 2 26376 57872
0 26419 5 1 1 26418
0 26420 7 1 2 40272 26419
0 26421 5 1 1 26420
0 26422 7 1 2 54095 50035
0 26423 5 1 1 26422
0 26424 7 1 2 40462 57746
0 26425 5 1 1 26424
0 26426 7 1 2 26423 26425
0 26427 7 1 2 26421 26426
0 26428 5 1 1 26427
0 26429 7 1 2 41257 26428
0 26430 5 1 1 26429
0 26431 7 1 2 46423 49543
0 26432 7 1 2 65947 26431
0 26433 5 1 1 26432
0 26434 7 1 2 26430 26433
0 26435 5 1 1 26434
0 26436 7 1 2 42156 26435
0 26437 5 1 1 26436
0 26438 7 1 2 49926 60687
0 26439 5 1 1 26438
0 26440 7 1 2 57059 65959
0 26441 5 1 1 26440
0 26442 7 1 2 26439 26441
0 26443 5 1 1 26442
0 26444 7 1 2 40089 26443
0 26445 5 1 1 26444
0 26446 7 1 2 51745 60210
0 26447 7 1 2 51425 26446
0 26448 7 1 2 62207 26447
0 26449 5 1 1 26448
0 26450 7 1 2 43931 26449
0 26451 7 1 2 26445 26450
0 26452 7 1 2 26437 26451
0 26453 5 1 1 26452
0 26454 7 1 2 26417 26453
0 26455 5 1 1 26454
0 26456 7 1 2 45763 26455
0 26457 5 1 1 26456
0 26458 7 1 2 57060 65961
0 26459 5 1 1 26458
0 26460 7 1 2 54096 65977
0 26461 5 1 1 26460
0 26462 7 1 2 42417 26461
0 26463 7 1 2 26459 26462
0 26464 5 1 1 26463
0 26465 7 1 2 45972 26464
0 26466 7 1 2 26457 26465
0 26467 5 1 1 26466
0 26468 7 1 2 26387 26467
0 26469 5 1 1 26468
0 26470 7 1 2 42865 26469
0 26471 5 1 1 26470
0 26472 7 1 2 59428 23844
0 26473 5 1 1 26472
0 26474 7 1 2 26294 26473
0 26475 5 1 1 26474
0 26476 7 1 2 43932 26475
0 26477 5 1 1 26476
0 26478 7 1 2 23109 26477
0 26479 5 1 1 26478
0 26480 7 1 2 53920 26479
0 26481 5 1 1 26480
0 26482 7 1 2 65257 57061
0 26483 5 1 1 26482
0 26484 7 1 2 52238 54097
0 26485 5 1 1 26484
0 26486 7 1 2 26483 26485
0 26487 5 1 1 26486
0 26488 7 1 2 45764 26487
0 26489 5 1 1 26488
0 26490 7 1 2 62098 65979
0 26491 5 1 1 26490
0 26492 7 1 2 26489 26491
0 26493 5 1 1 26492
0 26494 7 1 2 43933 55827
0 26495 7 1 2 26493 26494
0 26496 5 1 1 26495
0 26497 7 1 2 26481 26496
0 26498 5 1 1 26497
0 26499 7 1 2 46147 26498
0 26500 5 1 1 26499
0 26501 7 1 2 26471 26500
0 26502 5 1 1 26501
0 26503 7 1 2 43014 60086
0 26504 7 1 2 26502 26503
0 26505 5 1 1 26504
0 26506 7 1 2 47026 65943
0 26507 5 1 1 26506
0 26508 7 2 2 40658 56289
0 26509 5 1 1 65996
0 26510 7 1 2 26507 26509
0 26511 5 1 1 26510
0 26512 7 1 2 42676 26511
0 26513 5 1 1 26512
0 26514 7 3 2 43934 51927
0 26515 5 2 1 65998
0 26516 7 1 2 47997 65999
0 26517 5 1 1 26516
0 26518 7 1 2 26513 26517
0 26519 5 2 1 26518
0 26520 7 1 2 62126 65853
0 26521 5 1 1 26520
0 26522 7 1 2 26521 60178
0 26523 5 1 1 26522
0 26524 7 1 2 66003 26523
0 26525 5 1 1 26524
0 26526 7 1 2 42157 65708
0 26527 7 1 2 60136 26526
0 26528 5 1 1 26527
0 26529 7 1 2 26525 26528
0 26530 5 1 1 26529
0 26531 7 1 2 48586 26530
0 26532 5 1 1 26531
0 26533 7 3 2 45168 46288
0 26534 7 2 2 56691 66005
0 26535 7 2 2 50287 55335
0 26536 7 1 2 53323 62127
0 26537 7 1 2 66010 26536
0 26538 7 1 2 66008 26537
0 26539 5 1 1 26538
0 26540 7 1 2 26532 26539
0 26541 5 1 1 26540
0 26542 7 1 2 40463 26541
0 26543 5 1 1 26542
0 26544 7 4 2 41387 45169
0 26545 7 1 2 42418 66012
0 26546 7 1 2 57691 26545
0 26547 7 1 2 62367 62152
0 26548 7 1 2 26546 26547
0 26549 5 1 1 26548
0 26550 7 1 2 26543 26549
0 26551 5 1 1 26550
0 26552 7 1 2 55082 26551
0 26553 5 1 1 26552
0 26554 7 1 2 66004 57097
0 26555 5 1 1 26554
0 26556 7 1 2 48164 57686
0 26557 7 1 2 62153 26556
0 26558 5 1 1 26557
0 26559 7 1 2 26555 26558
0 26560 5 1 1 26559
0 26561 7 1 2 48587 26560
0 26562 5 1 1 26561
0 26563 7 2 2 57484 53476
0 26564 7 2 2 50751 61879
0 26565 7 1 2 60773 66018
0 26566 7 1 2 66016 26565
0 26567 5 1 1 26566
0 26568 7 1 2 26562 26567
0 26569 5 1 1 26568
0 26570 7 1 2 40464 26569
0 26571 5 1 1 26570
0 26572 7 2 2 55618 62966
0 26573 5 1 1 66020
0 26574 7 1 2 63843 53649
0 26575 7 1 2 61156 26574
0 26576 7 1 2 66021 26575
0 26577 5 1 1 26576
0 26578 7 1 2 26571 26577
0 26579 5 1 1 26578
0 26580 7 1 2 60087 26579
0 26581 5 1 1 26580
0 26582 7 1 2 26553 26581
0 26583 5 1 1 26582
0 26584 7 1 2 52110 26583
0 26585 5 1 1 26584
0 26586 7 5 2 45114 45170
0 26587 7 1 2 55433 66022
0 26588 7 1 2 63275 26587
0 26589 7 1 2 56577 26588
0 26590 7 1 2 59876 26589
0 26591 5 1 1 26590
0 26592 7 1 2 26585 26591
0 26593 7 1 2 26505 26592
0 26594 7 1 2 26318 26593
0 26595 7 1 2 26102 26594
0 26596 5 1 1 26595
0 26597 7 1 2 41515 26596
0 26598 5 1 1 26597
0 26599 7 1 2 46812 60119
0 26600 5 1 1 26599
0 26601 7 1 2 65285 57406
0 26602 5 1 1 26601
0 26603 7 1 2 26600 26602
0 26604 5 1 1 26603
0 26605 7 1 2 40465 26604
0 26606 5 1 1 26605
0 26607 7 1 2 41388 65841
0 26608 5 1 1 26607
0 26609 7 1 2 26606 26608
0 26610 5 1 1 26609
0 26611 7 1 2 42419 26610
0 26612 5 1 1 26611
0 26613 7 1 2 25591 26612
0 26614 5 1 1 26613
0 26615 7 1 2 40090 26614
0 26616 5 1 1 26615
0 26617 7 1 2 56890 62093
0 26618 7 1 2 65838 26617
0 26619 5 1 1 26618
0 26620 7 1 2 26616 26619
0 26621 5 1 1 26620
0 26622 7 1 2 65927 26621
0 26623 5 1 1 26622
0 26624 7 3 2 54782 59429
0 26625 5 1 1 66027
0 26626 7 2 2 60137 66028
0 26627 7 1 2 40466 66030
0 26628 5 1 1 26627
0 26629 7 1 2 45973 53034
0 26630 7 1 2 65829 26629
0 26631 5 1 1 26630
0 26632 7 1 2 26628 26631
0 26633 5 1 1 26632
0 26634 7 1 2 55480 26633
0 26635 5 1 1 26634
0 26636 7 1 2 26623 26635
0 26637 5 1 1 26636
0 26638 7 1 2 41516 26637
0 26639 5 1 1 26638
0 26640 7 2 2 40091 63347
0 26641 7 1 2 48707 66032
0 26642 7 1 2 66031 26641
0 26643 5 1 1 26642
0 26644 7 1 2 26639 26643
0 26645 5 1 1 26644
0 26646 7 1 2 40273 26645
0 26647 5 1 1 26646
0 26648 7 2 2 65368 62517
0 26649 7 1 2 53498 60120
0 26650 7 1 2 66034 26649
0 26651 5 1 1 26650
0 26652 7 1 2 26647 26651
0 26653 5 1 1 26652
0 26654 7 1 2 48588 26653
0 26655 5 1 1 26654
0 26656 7 1 2 56900 57954
0 26657 7 2 2 57950 26656
0 26658 7 1 2 65844 66036
0 26659 5 1 1 26658
0 26660 7 1 2 26655 26659
0 26661 5 1 1 26660
0 26662 7 1 2 55083 26661
0 26663 5 1 1 26662
0 26664 7 1 2 40467 57848
0 26665 5 1 1 26664
0 26666 7 1 2 41389 57739
0 26667 5 1 1 26666
0 26668 7 1 2 26665 26667
0 26669 5 1 1 26668
0 26670 7 1 2 42420 26669
0 26671 5 1 1 26670
0 26672 7 1 2 54783 57740
0 26673 5 1 1 26672
0 26674 7 1 2 26671 26673
0 26675 5 1 1 26674
0 26676 7 1 2 40092 26675
0 26677 5 1 1 26676
0 26678 7 1 2 46813 63998
0 26679 5 1 1 26678
0 26680 7 1 2 26677 26679
0 26681 5 1 1 26680
0 26682 7 1 2 65928 26681
0 26683 5 1 1 26682
0 26684 7 1 2 66000 61096
0 26685 5 1 1 26684
0 26686 7 1 2 66029 63995
0 26687 5 1 1 26686
0 26688 7 1 2 26685 26687
0 26689 5 1 1 26688
0 26690 7 1 2 55481 26689
0 26691 5 1 1 26690
0 26692 7 1 2 26683 26691
0 26693 5 1 1 26692
0 26694 7 1 2 41517 26693
0 26695 5 1 1 26694
0 26696 7 1 2 53434 53344
0 26697 7 1 2 62582 26696
0 26698 7 1 2 65778 26697
0 26699 5 1 1 26698
0 26700 7 1 2 26695 26699
0 26701 5 1 1 26700
0 26702 7 1 2 40274 26701
0 26703 5 1 1 26702
0 26704 7 1 2 41390 61794
0 26705 7 1 2 66035 26704
0 26706 5 1 1 26705
0 26707 7 1 2 26703 26706
0 26708 5 1 1 26707
0 26709 7 1 2 48589 26708
0 26710 5 1 1 26709
0 26711 7 1 2 63500 56382
0 26712 7 1 2 57951 26711
0 26713 7 1 2 64106 26712
0 26714 5 1 1 26713
0 26715 7 1 2 26710 26714
0 26716 5 1 1 26715
0 26717 7 1 2 60088 26716
0 26718 5 1 1 26717
0 26719 7 1 2 26663 26718
0 26720 5 1 1 26719
0 26721 7 1 2 47125 26720
0 26722 5 1 1 26721
0 26723 7 1 2 65626 60171
0 26724 5 1 1 26723
0 26725 7 1 2 52457 58574
0 26726 7 1 2 63411 26725
0 26727 7 1 2 53441 26726
0 26728 7 1 2 65845 26727
0 26729 5 1 1 26728
0 26730 7 1 2 26724 26729
0 26731 5 1 1 26730
0 26732 7 1 2 55084 26731
0 26733 5 1 1 26732
0 26734 7 1 2 65627 57062
0 26735 5 1 1 26734
0 26736 7 1 2 60803 56627
0 26737 7 1 2 66019 26736
0 26738 7 1 2 65780 26737
0 26739 5 1 1 26738
0 26740 7 1 2 26735 26739
0 26741 5 1 1 26740
0 26742 7 1 2 60089 26741
0 26743 5 1 1 26742
0 26744 7 1 2 26733 26743
0 26745 5 1 1 26744
0 26746 7 1 2 43015 26745
0 26747 5 1 1 26746
0 26748 7 1 2 26722 26747
0 26749 7 1 2 26598 26748
0 26750 5 1 1 26749
0 26751 7 1 2 43240 26750
0 26752 5 1 1 26751
0 26753 7 1 2 65567 50109
0 26754 5 1 1 26753
0 26755 7 1 2 60230 65371
0 26756 7 1 2 65609 26755
0 26757 5 1 1 26756
0 26758 7 1 2 26754 26757
0 26759 5 1 1 26758
0 26760 7 1 2 43576 26759
0 26761 5 1 1 26760
0 26762 7 1 2 63910 47851
0 26763 7 1 2 51618 26762
0 26764 5 1 1 26763
0 26765 7 1 2 26761 26764
0 26766 5 1 1 26765
0 26767 7 1 2 42158 26766
0 26768 5 1 1 26767
0 26769 7 1 2 60833 62607
0 26770 5 1 1 26769
0 26771 7 1 2 49776 60973
0 26772 5 1 1 26771
0 26773 7 1 2 26770 26772
0 26774 5 1 1 26773
0 26775 7 1 2 55823 62967
0 26776 7 1 2 26774 26775
0 26777 5 1 1 26776
0 26778 7 1 2 26768 26777
0 26779 5 1 1 26778
0 26780 7 1 2 45765 26779
0 26781 5 1 1 26780
0 26782 7 1 2 64101 52505
0 26783 5 1 1 26782
0 26784 7 1 2 47482 14738
0 26785 7 1 2 58500 26784
0 26786 5 1 1 26785
0 26787 7 1 2 26783 26786
0 26788 5 1 1 26787
0 26789 7 1 2 40275 26788
0 26790 5 1 1 26789
0 26791 7 3 2 41977 65444
0 26792 5 1 1 66038
0 26793 7 1 2 42159 66039
0 26794 5 1 1 26793
0 26795 7 1 2 65417 26794
0 26796 5 2 1 26795
0 26797 7 1 2 55458 66041
0 26798 5 1 1 26797
0 26799 7 1 2 26790 26798
0 26800 5 1 1 26799
0 26801 7 1 2 40659 26800
0 26802 5 1 1 26801
0 26803 7 1 2 51746 55655
0 26804 7 1 2 62571 26803
0 26805 5 1 1 26804
0 26806 7 1 2 26802 26805
0 26807 5 1 1 26806
0 26808 7 1 2 42866 56546
0 26809 7 1 2 26807 26808
0 26810 5 1 1 26809
0 26811 7 1 2 26781 26810
0 26812 5 1 1 26811
0 26813 7 2 2 65532 57292
0 26814 7 1 2 62803 66043
0 26815 7 1 2 26812 26814
0 26816 5 1 1 26815
0 26817 7 1 2 26752 26816
0 26818 7 1 2 25971 26817
0 26819 5 1 1 26818
0 26820 7 1 2 44320 26819
0 26821 5 1 1 26820
0 26822 7 1 2 25167 26821
0 26823 5 1 1 26822
0 26824 7 1 2 48077 26823
0 26825 5 1 1 26824
0 26826 7 4 2 43241 65181
0 26827 7 1 2 65785 66045
0 26828 5 1 1 26827
0 26829 7 3 2 43242 55537
0 26830 5 1 1 66049
0 26831 7 1 2 56260 62435
0 26832 5 1 1 26831
0 26833 7 1 2 26830 26832
0 26834 5 1 1 26833
0 26835 7 1 2 41846 26834
0 26836 5 1 1 26835
0 26837 7 1 2 65372 65149
0 26838 5 1 1 26837
0 26839 7 1 2 26836 26838
0 26840 5 1 1 26839
0 26841 7 1 2 44525 26840
0 26842 5 1 1 26841
0 26843 7 1 2 47347 48826
0 26844 7 1 2 66046 26843
0 26845 5 1 1 26844
0 26846 7 1 2 26842 26845
0 26847 5 1 1 26846
0 26848 7 1 2 42160 26847
0 26849 5 1 1 26848
0 26850 7 5 2 42677 53703
0 26851 5 2 1 66052
0 26852 7 1 2 58690 55538
0 26853 5 1 1 26852
0 26854 7 1 2 66057 26853
0 26855 5 1 1 26854
0 26856 7 1 2 59694 26855
0 26857 5 1 1 26856
0 26858 7 1 2 26849 26857
0 26859 5 1 1 26858
0 26860 7 1 2 43577 26859
0 26861 5 1 1 26860
0 26862 7 2 2 47091 55539
0 26863 5 2 1 66059
0 26864 7 1 2 66058 66061
0 26865 5 5 1 26864
0 26866 7 1 2 44526 66053
0 26867 5 1 1 26866
0 26868 7 1 2 40093 26867
0 26869 5 1 1 26868
0 26870 7 2 2 66063 26869
0 26871 7 1 2 59695 66068
0 26872 5 1 1 26871
0 26873 7 1 2 26861 26872
0 26874 5 1 1 26873
0 26875 7 1 2 43742 26874
0 26876 5 1 1 26875
0 26877 7 1 2 55151 59696
0 26878 7 1 2 66064 26877
0 26879 5 1 1 26878
0 26880 7 1 2 46148 26879
0 26881 7 1 2 26876 26880
0 26882 5 1 1 26881
0 26883 7 1 2 45171 50238
0 26884 5 1 1 26883
0 26885 7 1 2 40276 59740
0 26886 7 1 2 26884 26885
0 26887 5 1 1 26886
0 26888 7 1 2 65243 26887
0 26889 5 1 1 26888
0 26890 7 1 2 40094 26889
0 26891 5 1 1 26890
0 26892 7 1 2 60033 59697
0 26893 5 1 1 26892
0 26894 7 1 2 26891 26893
0 26895 5 1 1 26894
0 26896 7 1 2 45326 26895
0 26897 5 1 1 26896
0 26898 7 2 2 47596 59698
0 26899 5 1 1 66070
0 26900 7 1 2 26897 26899
0 26901 5 2 1 26900
0 26902 7 1 2 64265 66072
0 26903 5 1 1 26902
0 26904 7 2 2 47803 65393
0 26905 7 1 2 55558 66074
0 26906 5 1 1 26905
0 26907 7 1 2 26903 26906
0 26908 5 1 1 26907
0 26909 7 1 2 45497 26908
0 26910 5 1 1 26909
0 26911 7 1 2 48176 65893
0 26912 5 1 1 26911
0 26913 7 1 2 47518 26912
0 26914 5 1 1 26913
0 26915 7 1 2 54790 65894
0 26916 5 1 1 26915
0 26917 7 1 2 47287 26916
0 26918 5 1 1 26917
0 26919 7 1 2 65001 26918
0 26920 7 1 2 26914 26919
0 26921 5 1 1 26920
0 26922 7 1 2 66047 26921
0 26923 5 1 1 26922
0 26924 7 1 2 26910 26923
0 26925 5 1 1 26924
0 26926 7 1 2 40468 26925
0 26927 5 1 1 26926
0 26928 7 1 2 41258 60548
0 26929 5 1 1 26928
0 26930 7 1 2 65440 64482
0 26931 5 1 1 26930
0 26932 7 1 2 41259 56290
0 26933 7 1 2 47519 26932
0 26934 5 1 1 26933
0 26935 7 1 2 26931 26934
0 26936 5 1 1 26935
0 26937 7 1 2 40277 26936
0 26938 5 1 1 26937
0 26939 7 1 2 26929 26938
0 26940 5 1 1 26939
0 26941 7 1 2 66048 26940
0 26942 5 1 1 26941
0 26943 7 1 2 42867 26942
0 26944 7 1 2 26927 26943
0 26945 5 1 1 26944
0 26946 7 1 2 40660 26945
0 26947 7 1 2 26882 26946
0 26948 5 1 1 26947
0 26949 7 1 2 26828 26948
0 26950 5 1 1 26949
0 26951 7 1 2 58893 26950
0 26952 5 1 1 26951
0 26953 7 2 2 55251 48708
0 26954 5 1 1 66076
0 26955 7 1 2 54232 53852
0 26956 5 1 1 26955
0 26957 7 1 2 26954 26956
0 26958 5 1 1 26957
0 26959 7 1 2 47804 26958
0 26960 5 1 1 26959
0 26961 7 2 2 55252 51593
0 26962 5 1 1 66078
0 26963 7 3 2 40095 43743
0 26964 7 1 2 61186 66080
0 26965 5 1 1 26964
0 26966 7 1 2 26962 26965
0 26967 5 1 1 26966
0 26968 7 1 2 45498 26967
0 26969 5 1 1 26968
0 26970 7 1 2 26960 26969
0 26971 5 1 1 26970
0 26972 7 1 2 42421 26971
0 26973 5 1 1 26972
0 26974 7 1 2 65685 63311
0 26975 5 1 1 26974
0 26976 7 1 2 26973 26975
0 26977 5 1 1 26976
0 26978 7 1 2 46761 26977
0 26979 5 1 1 26978
0 26980 7 1 2 46149 65722
0 26981 5 1 1 26980
0 26982 7 2 2 57576 51335
0 26983 7 1 2 52006 66083
0 26984 7 1 2 58642 26983
0 26985 5 1 1 26984
0 26986 7 1 2 26981 26985
0 26987 5 1 1 26986
0 26988 7 1 2 42678 26987
0 26989 5 1 1 26988
0 26990 7 1 2 47805 65799
0 26991 5 1 1 26990
0 26992 7 1 2 42422 62532
0 26993 5 1 1 26992
0 26994 7 1 2 26991 26993
0 26995 5 1 1 26994
0 26996 7 1 2 49544 26995
0 26997 5 1 1 26996
0 26998 7 1 2 46849 54755
0 26999 5 1 1 26998
0 27000 7 1 2 59779 26999
0 27001 5 1 1 27000
0 27002 7 1 2 26997 27001
0 27003 5 1 1 27002
0 27004 7 1 2 40096 27003
0 27005 5 1 1 27004
0 27006 7 1 2 41140 53560
0 27007 7 1 2 58262 27006
0 27008 5 1 1 27007
0 27009 7 2 2 42161 51960
0 27010 5 1 1 66085
0 27011 7 1 2 4009 27010
0 27012 5 1 1 27011
0 27013 7 1 2 41391 27012
0 27014 5 1 1 27013
0 27015 7 1 2 47189 61076
0 27016 5 1 1 27015
0 27017 7 1 2 65717 27016
0 27018 5 1 1 27017
0 27019 7 1 2 45766 27018
0 27020 5 1 1 27019
0 27021 7 1 2 27014 27020
0 27022 5 1 1 27021
0 27023 7 1 2 40278 27022
0 27024 5 1 1 27023
0 27025 7 1 2 27008 27024
0 27026 7 1 2 27005 27025
0 27027 5 1 1 27026
0 27028 7 1 2 55253 27027
0 27029 5 1 1 27028
0 27030 7 1 2 26989 27029
0 27031 7 1 2 26979 27030
0 27032 5 2 1 27031
0 27033 7 1 2 61520 65793
0 27034 7 1 2 66087 27033
0 27035 5 1 1 27034
0 27036 7 1 2 26952 27035
0 27037 5 1 1 27036
0 27038 7 1 2 43016 27037
0 27039 5 1 1 27038
0 27040 7 2 2 65394 57543
0 27041 7 1 2 44687 66089
0 27042 5 1 1 27041
0 27043 7 1 2 60148 65157
0 27044 7 1 2 62974 27043
0 27045 7 1 2 65614 27044
0 27046 5 1 1 27045
0 27047 7 1 2 27042 27046
0 27048 5 1 1 27047
0 27049 7 1 2 47348 27048
0 27050 5 1 1 27049
0 27051 7 1 2 41978 66090
0 27052 5 1 1 27051
0 27053 7 2 2 45172 56185
0 27054 7 1 2 55413 62975
0 27055 7 1 2 66091 27054
0 27056 5 1 1 27055
0 27057 7 1 2 27052 27056
0 27058 5 1 1 27057
0 27059 7 1 2 43408 27058
0 27060 5 1 1 27059
0 27061 7 1 2 48827 65173
0 27062 7 1 2 65771 27061
0 27063 5 1 1 27062
0 27064 7 1 2 27060 27063
0 27065 5 1 1 27064
0 27066 7 1 2 44431 27065
0 27067 5 1 1 27066
0 27068 7 1 2 65461 2636
0 27069 5 3 1 27068
0 27070 7 1 2 59699 66093
0 27071 5 1 1 27070
0 27072 7 1 2 27067 27071
0 27073 5 1 1 27072
0 27074 7 1 2 44527 27073
0 27075 5 1 1 27074
0 27076 7 1 2 27050 27075
0 27077 5 1 1 27076
0 27078 7 1 2 42162 27077
0 27079 5 1 1 27078
0 27080 7 1 2 65747 65204
0 27081 5 1 1 27080
0 27082 7 1 2 55467 54217
0 27083 5 1 1 27082
0 27084 7 1 2 27081 27083
0 27085 5 1 1 27084
0 27086 7 1 2 47419 27085
0 27087 5 1 1 27086
0 27088 7 1 2 64928 57598
0 27089 5 1 1 27088
0 27090 7 1 2 27087 27089
0 27091 5 1 1 27090
0 27092 7 1 2 59700 27091
0 27093 5 1 1 27092
0 27094 7 1 2 27079 27093
0 27095 5 1 1 27094
0 27096 7 1 2 58894 27095
0 27097 5 1 1 27096
0 27098 7 3 2 43409 65408
0 27099 5 1 1 66096
0 27100 7 2 2 60331 66097
0 27101 7 1 2 61300 60779
0 27102 7 1 2 66099 27101
0 27103 7 1 2 65463 27102
0 27104 5 1 1 27103
0 27105 7 1 2 27097 27104
0 27106 5 1 1 27105
0 27107 7 1 2 43578 27106
0 27108 5 1 1 27107
0 27109 7 1 2 63036 64929
0 27110 5 1 1 27109
0 27111 7 3 2 56271 51367
0 27112 5 1 1 66101
0 27113 7 1 2 64926 27112
0 27114 7 1 2 27110 27113
0 27115 5 1 1 27114
0 27116 7 1 2 45974 27115
0 27117 5 1 1 27116
0 27118 7 1 2 52475 27117
0 27119 5 1 1 27118
0 27120 7 1 2 48128 27119
0 27121 5 1 1 27120
0 27122 7 1 2 47936 51368
0 27123 7 1 2 65519 27122
0 27124 5 1 1 27123
0 27125 7 1 2 27121 27124
0 27126 5 1 1 27125
0 27127 7 1 2 65412 27126
0 27128 5 1 1 27127
0 27129 7 1 2 27108 27128
0 27130 5 1 1 27129
0 27131 7 1 2 43744 27130
0 27132 5 1 1 27131
0 27133 7 1 2 59857 66073
0 27134 5 1 1 27133
0 27135 7 1 2 53839 47288
0 27136 7 1 2 66075 27135
0 27137 5 1 1 27136
0 27138 7 1 2 27134 27137
0 27139 5 1 1 27138
0 27140 7 1 2 40469 27139
0 27141 5 1 1 27140
0 27142 7 1 2 52007 59874
0 27143 5 1 1 27142
0 27144 7 1 2 57919 52568
0 27145 5 1 1 27144
0 27146 7 1 2 27143 27145
0 27147 5 1 1 27146
0 27148 7 1 2 42679 27147
0 27149 5 1 1 27148
0 27150 7 1 2 47483 55892
0 27151 5 1 1 27150
0 27152 7 1 2 45327 49917
0 27153 7 1 2 25595 27152
0 27154 5 1 1 27153
0 27155 7 1 2 27151 27154
0 27156 5 1 1 27155
0 27157 7 1 2 51928 27156
0 27158 5 1 1 27157
0 27159 7 1 2 27149 27158
0 27160 5 1 1 27159
0 27161 7 2 2 46150 59701
0 27162 7 1 2 27160 66104
0 27163 5 1 1 27162
0 27164 7 1 2 27141 27163
0 27165 5 1 1 27164
0 27166 7 1 2 45499 27165
0 27167 5 1 1 27166
0 27168 7 1 2 65741 51616
0 27169 5 1 1 27168
0 27170 7 1 2 42680 27169
0 27171 5 1 1 27170
0 27172 7 1 2 49831 55474
0 27173 5 1 1 27172
0 27174 7 1 2 42423 27173
0 27175 7 1 2 27171 27174
0 27176 5 1 1 27175
0 27177 7 1 2 42163 49864
0 27178 5 1 1 27177
0 27179 7 2 2 64801 27178
0 27180 5 1 1 66106
0 27181 7 1 2 42681 27180
0 27182 5 1 1 27181
0 27183 7 1 2 40097 48033
0 27184 5 1 1 27183
0 27185 7 1 2 54302 27184
0 27186 7 1 2 61132 27185
0 27187 5 1 1 27186
0 27188 7 1 2 45767 27187
0 27189 7 1 2 27182 27188
0 27190 5 1 1 27189
0 27191 7 1 2 66105 27190
0 27192 7 1 2 27176 27191
0 27193 5 1 1 27192
0 27194 7 1 2 27167 27193
0 27195 5 1 1 27194
0 27196 7 1 2 43017 27195
0 27197 5 1 1 27196
0 27198 7 1 2 55824 65167
0 27199 7 1 2 62764 27198
0 27200 7 1 2 52805 51176
0 27201 7 1 2 27199 27200
0 27202 5 1 1 27201
0 27203 7 1 2 27197 27202
0 27204 5 1 1 27203
0 27205 7 1 2 58895 27204
0 27206 5 1 1 27205
0 27207 7 1 2 65005 25119
0 27208 5 2 1 27207
0 27209 7 1 2 53840 66108
0 27210 5 1 1 27209
0 27211 7 1 2 64997 27210
0 27212 5 1 1 27211
0 27213 7 1 2 47289 27212
0 27214 5 1 1 27213
0 27215 7 1 2 56196 50532
0 27216 7 1 2 59858 27215
0 27217 5 1 1 27216
0 27218 7 1 2 27214 27217
0 27219 5 1 1 27218
0 27220 7 1 2 65794 57119
0 27221 7 1 2 27219 27220
0 27222 5 1 1 27221
0 27223 7 1 2 27206 27222
0 27224 7 1 2 27132 27223
0 27225 5 1 1 27224
0 27226 7 1 2 43935 27225
0 27227 5 1 1 27226
0 27228 7 1 2 27039 27227
0 27229 5 1 1 27228
0 27230 7 1 2 44321 27229
0 27231 5 1 1 27230
0 27232 7 1 2 24836 65745
0 27233 5 1 1 27232
0 27234 7 1 2 42682 27233
0 27235 5 1 1 27234
0 27236 7 1 2 65749 27235
0 27237 5 1 1 27236
0 27238 7 1 2 43936 27237
0 27239 5 1 1 27238
0 27240 7 1 2 65638 1806
0 27241 5 1 1 27240
0 27242 7 1 2 65759 27241
0 27243 5 1 1 27242
0 27244 7 2 2 42683 55865
0 27245 5 1 1 66110
0 27246 7 1 2 52185 61653
0 27247 5 1 1 27246
0 27248 7 1 2 27245 27247
0 27249 5 1 1 27248
0 27250 7 1 2 43745 27249
0 27251 5 1 1 27250
0 27252 7 1 2 27243 27251
0 27253 5 1 1 27252
0 27254 7 1 2 46151 27253
0 27255 5 1 1 27254
0 27256 7 1 2 55254 65743
0 27257 5 1 1 27256
0 27258 7 1 2 27255 27257
0 27259 5 1 1 27258
0 27260 7 1 2 40661 27259
0 27261 5 1 1 27260
0 27262 7 1 2 65632 27261
0 27263 5 1 1 27262
0 27264 7 1 2 43018 27263
0 27265 5 1 1 27264
0 27266 7 1 2 27239 27265
0 27267 5 1 1 27266
0 27268 7 1 2 42424 27267
0 27269 5 1 1 27268
0 27270 7 1 2 53601 65761
0 27271 7 1 2 63231 27270
0 27272 5 1 1 27271
0 27273 7 1 2 19687 3481
0 27274 5 2 1 27273
0 27275 7 1 2 66112 62460
0 27276 5 1 1 27275
0 27277 7 1 2 65929 54218
0 27278 5 1 1 27277
0 27279 7 1 2 27276 27278
0 27280 5 1 1 27279
0 27281 7 1 2 43746 55688
0 27282 7 1 2 27280 27281
0 27283 5 1 1 27282
0 27284 7 1 2 27272 27283
0 27285 5 1 1 27284
0 27286 7 1 2 48010 27285
0 27287 5 1 1 27286
0 27288 7 1 2 41392 50249
0 27289 5 1 1 27288
0 27290 7 1 2 47806 50154
0 27291 5 1 1 27290
0 27292 7 1 2 27289 27291
0 27293 5 1 1 27292
0 27294 7 1 2 45500 27293
0 27295 5 1 1 27294
0 27296 7 1 2 66107 27295
0 27297 5 1 1 27296
0 27298 7 1 2 43937 27297
0 27299 5 1 1 27298
0 27300 7 1 2 43938 50288
0 27301 5 2 1 27300
0 27302 7 1 2 65971 61306
0 27303 5 1 1 27302
0 27304 7 1 2 66114 27303
0 27305 5 1 1 27304
0 27306 7 1 2 43410 27305
0 27307 5 1 1 27306
0 27308 7 1 2 44528 56139
0 27309 5 1 1 27308
0 27310 7 1 2 66115 27309
0 27311 5 1 1 27310
0 27312 7 1 2 43747 27311
0 27313 5 1 1 27312
0 27314 7 1 2 27307 27313
0 27315 7 1 2 27299 27314
0 27316 5 1 1 27315
0 27317 7 1 2 46152 27316
0 27318 5 1 1 27317
0 27319 7 2 2 50289 58465
0 27320 7 1 2 56803 66116
0 27321 5 1 1 27320
0 27322 7 1 2 42684 27321
0 27323 7 1 2 27318 27322
0 27324 5 1 1 27323
0 27325 7 1 2 40470 66117
0 27326 5 1 1 27325
0 27327 7 1 2 24878 65028
0 27328 5 1 1 27327
0 27329 7 1 2 59240 27328
0 27330 5 1 1 27329
0 27331 7 1 2 27326 27330
0 27332 5 1 1 27331
0 27333 7 1 2 43939 27332
0 27334 5 1 1 27333
0 27335 7 1 2 56805 53182
0 27336 5 1 1 27335
0 27337 7 1 2 65642 27336
0 27338 5 1 1 27337
0 27339 7 2 2 44688 52357
0 27340 5 1 1 66118
0 27341 7 1 2 40662 27340
0 27342 5 1 1 27341
0 27343 7 2 2 44432 46153
0 27344 7 1 2 48617 66120
0 27345 7 1 2 47148 27344
0 27346 7 1 2 27342 27345
0 27347 5 1 1 27346
0 27348 7 1 2 27338 27347
0 27349 5 1 1 27348
0 27350 7 1 2 41979 27349
0 27351 5 1 1 27350
0 27352 7 1 2 40663 49865
0 27353 5 1 1 27352
0 27354 7 1 2 47661 56806
0 27355 5 1 1 27354
0 27356 7 1 2 54967 47520
0 27357 7 1 2 27355 27356
0 27358 5 1 1 27357
0 27359 7 1 2 27353 27358
0 27360 5 1 1 27359
0 27361 7 1 2 47958 27360
0 27362 5 1 1 27361
0 27363 7 1 2 45975 27362
0 27364 7 1 2 27351 27363
0 27365 7 1 2 27334 27364
0 27366 5 1 1 27365
0 27367 7 1 2 51294 27366
0 27368 7 1 2 27324 27367
0 27369 5 1 1 27368
0 27370 7 1 2 27287 27369
0 27371 7 1 2 27269 27370
0 27372 5 1 1 27371
0 27373 7 1 2 58896 27372
0 27374 5 1 1 27373
0 27375 7 2 2 53841 54805
0 27376 5 2 1 66122
0 27377 7 1 2 24433 66124
0 27378 5 1 1 27377
0 27379 7 1 2 47290 27378
0 27380 5 1 1 27379
0 27381 7 1 2 47521 66123
0 27382 5 1 1 27381
0 27383 7 1 2 46762 66077
0 27384 5 1 1 27383
0 27385 7 1 2 27382 27384
0 27386 7 1 2 27380 27385
0 27387 5 1 1 27386
0 27388 7 1 2 42425 27387
0 27389 5 1 1 27388
0 27390 7 2 2 52186 64358
0 27391 5 1 1 66126
0 27392 7 1 2 40098 66127
0 27393 5 1 1 27392
0 27394 7 1 2 52187 51961
0 27395 7 1 2 53057 27394
0 27396 5 1 1 27395
0 27397 7 1 2 27393 27396
0 27398 7 1 2 27389 27397
0 27399 5 1 1 27398
0 27400 7 1 2 40664 27399
0 27401 5 1 1 27400
0 27402 7 2 2 64266 51336
0 27403 7 1 2 60825 66128
0 27404 5 1 1 27403
0 27405 7 1 2 56508 64846
0 27406 5 1 1 27405
0 27407 7 1 2 27404 27406
0 27408 5 1 1 27407
0 27409 7 1 2 41141 27408
0 27410 5 1 1 27409
0 27411 7 1 2 55719 56291
0 27412 5 1 1 27411
0 27413 7 1 2 27410 27412
0 27414 5 1 1 27413
0 27415 7 1 2 57577 27414
0 27416 5 1 1 27415
0 27417 7 1 2 27401 27416
0 27418 5 1 1 27417
0 27419 7 1 2 47807 27418
0 27420 5 1 1 27419
0 27421 7 6 2 43940 54656
0 27422 7 1 2 65751 66130
0 27423 5 1 1 27422
0 27424 7 1 2 65644 47557
0 27425 5 1 1 27424
0 27426 7 1 2 58692 66079
0 27427 5 1 1 27426
0 27428 7 1 2 27425 27427
0 27429 5 1 1 27428
0 27430 7 1 2 45501 27429
0 27431 5 1 1 27430
0 27432 7 1 2 51594 58251
0 27433 5 1 1 27432
0 27434 7 1 2 59802 27433
0 27435 5 1 1 27434
0 27436 7 1 2 55255 27435
0 27437 5 1 1 27436
0 27438 7 1 2 42426 27437
0 27439 7 1 2 27431 27438
0 27440 5 1 1 27439
0 27441 7 1 2 46763 65686
0 27442 5 1 1 27441
0 27443 7 1 2 40099 61762
0 27444 5 1 1 27443
0 27445 7 1 2 46814 55459
0 27446 5 1 1 27445
0 27447 7 1 2 27444 27446
0 27448 7 1 2 27442 27447
0 27449 5 1 1 27448
0 27450 7 1 2 47597 51337
0 27451 7 1 2 27449 27450
0 27452 5 1 1 27451
0 27453 7 1 2 24733 65035
0 27454 5 1 1 27453
0 27455 7 1 2 42164 27454
0 27456 5 1 1 27455
0 27457 7 1 2 45768 27456
0 27458 7 1 2 27452 27457
0 27459 5 1 1 27458
0 27460 7 1 2 40665 27459
0 27461 7 1 2 27440 27460
0 27462 5 1 1 27461
0 27463 7 1 2 27423 27462
0 27464 7 1 2 27420 27463
0 27465 5 1 1 27464
0 27466 7 1 2 64864 27465
0 27467 5 1 1 27466
0 27468 7 1 2 27374 27467
0 27469 5 1 1 27468
0 27470 7 1 2 65225 27469
0 27471 5 1 1 27470
0 27472 7 1 2 27231 27471
0 27473 5 1 1 27472
0 27474 7 1 2 44815 27473
0 27475 5 1 1 27474
0 27476 7 1 2 43941 66088
0 27477 5 1 1 27476
0 27478 7 3 2 48165 55825
0 27479 7 2 2 52513 66136
0 27480 7 1 2 56235 66139
0 27481 5 1 1 27480
0 27482 7 1 2 27477 27481
0 27483 5 1 1 27482
0 27484 7 1 2 41518 27483
0 27485 5 1 1 27484
0 27486 7 3 2 40471 50232
0 27487 5 1 1 66141
0 27488 7 1 2 66142 62280
0 27489 7 1 2 66140 27488
0 27490 5 1 1 27489
0 27491 7 1 2 27485 27490
0 27492 5 1 1 27491
0 27493 7 1 2 58913 27492
0 27494 5 1 1 27493
0 27495 7 1 2 41519 66069
0 27496 5 1 1 27495
0 27497 7 4 2 41520 52458
0 27498 5 1 1 66144
0 27499 7 1 2 44529 50446
0 27500 5 2 1 27499
0 27501 7 1 2 60887 66148
0 27502 5 2 1 27501
0 27503 7 1 2 47349 66150
0 27504 5 1 1 27503
0 27505 7 1 2 47126 58693
0 27506 5 1 1 27505
0 27507 7 1 2 41521 27506
0 27508 5 1 1 27507
0 27509 7 1 2 27504 27508
0 27510 5 1 1 27509
0 27511 7 1 2 42427 27510
0 27512 5 1 1 27511
0 27513 7 1 2 46719 66102
0 27514 5 1 1 27513
0 27515 7 1 2 27512 27514
0 27516 5 1 1 27515
0 27517 7 1 2 45976 27516
0 27518 5 1 1 27517
0 27519 7 1 2 27498 27518
0 27520 5 1 1 27519
0 27521 7 1 2 44689 27520
0 27522 5 1 1 27521
0 27523 7 2 2 42685 55992
0 27524 5 1 1 66152
0 27525 7 1 2 56261 58172
0 27526 5 1 1 27525
0 27527 7 1 2 27524 27526
0 27528 5 1 1 27527
0 27529 7 1 2 41522 27528
0 27530 5 1 1 27529
0 27531 7 1 2 27522 27530
0 27532 5 1 1 27531
0 27533 7 1 2 43579 27532
0 27534 5 1 1 27533
0 27535 7 1 2 27496 27534
0 27536 5 1 1 27535
0 27537 7 1 2 43748 27536
0 27538 5 1 1 27537
0 27539 7 1 2 62454 62419
0 27540 7 1 2 66065 27539
0 27541 5 1 1 27540
0 27542 7 1 2 27538 27541
0 27543 5 1 1 27542
0 27544 7 1 2 43942 27543
0 27545 5 1 1 27544
0 27546 7 1 2 55140 55944
0 27547 7 1 2 66153 27546
0 27548 5 1 1 27547
0 27549 7 1 2 46154 27548
0 27550 7 1 2 27545 27549
0 27551 5 1 1 27550
0 27552 7 2 2 54822 56292
0 27553 5 1 1 66154
0 27554 7 1 2 66155 64624
0 27555 5 1 1 27554
0 27556 7 2 2 41980 55214
0 27557 5 1 1 66156
0 27558 7 1 2 66001 27557
0 27559 5 1 1 27558
0 27560 7 1 2 40472 27559
0 27561 5 1 1 27560
0 27562 7 1 2 54823 57920
0 27563 5 1 1 27562
0 27564 7 1 2 27561 27563
0 27565 5 1 1 27564
0 27566 7 1 2 41523 27565
0 27567 5 1 1 27566
0 27568 7 1 2 54784 65568
0 27569 5 1 1 27568
0 27570 7 1 2 27567 27569
0 27571 5 1 1 27570
0 27572 7 1 2 55579 27571
0 27573 5 1 1 27572
0 27574 7 1 2 27555 27573
0 27575 5 1 1 27574
0 27576 7 1 2 47808 27575
0 27577 5 1 1 27576
0 27578 7 2 2 56706 48166
0 27579 5 1 1 66158
0 27580 7 2 2 50185 57173
0 27581 7 1 2 66159 66160
0 27582 5 1 1 27581
0 27583 7 1 2 45977 56293
0 27584 5 1 1 27583
0 27585 7 1 2 47809 65702
0 27586 5 1 1 27585
0 27587 7 1 2 27584 27586
0 27588 5 1 1 27587
0 27589 7 1 2 62518 27588
0 27590 5 1 1 27589
0 27591 7 1 2 66002 27579
0 27592 5 1 1 27591
0 27593 7 1 2 40473 27592
0 27594 5 1 1 27593
0 27595 7 1 2 27594 27553
0 27596 5 1 1 27595
0 27597 7 1 2 47598 27596
0 27598 5 1 1 27597
0 27599 7 1 2 27590 27598
0 27600 5 1 1 27599
0 27601 7 1 2 41524 27600
0 27602 5 1 1 27601
0 27603 7 1 2 27582 27602
0 27604 5 1 1 27603
0 27605 7 1 2 47522 27604
0 27606 5 1 1 27605
0 27607 7 2 2 50186 62348
0 27608 5 1 1 66162
0 27609 7 1 2 57911 27608
0 27610 5 1 1 27609
0 27611 7 1 2 62487 27610
0 27612 5 1 1 27611
0 27613 7 1 2 51876 64506
0 27614 5 2 1 27613
0 27615 7 1 2 27612 66164
0 27616 5 1 1 27615
0 27617 7 1 2 45978 27616
0 27618 5 1 1 27617
0 27619 7 2 2 54657 62968
0 27620 7 1 2 52459 66166
0 27621 5 1 1 27620
0 27622 7 1 2 27618 27621
0 27623 5 1 1 27622
0 27624 7 1 2 43943 27623
0 27625 5 1 1 27624
0 27626 7 2 2 59787 55215
0 27627 7 1 2 62608 66168
0 27628 5 1 1 27627
0 27629 7 1 2 27625 27628
0 27630 5 1 1 27629
0 27631 7 1 2 41525 27630
0 27632 5 1 1 27631
0 27633 7 2 2 52400 56901
0 27634 7 1 2 66169 66170
0 27635 5 1 1 27634
0 27636 7 1 2 42868 27635
0 27637 7 1 2 27632 27636
0 27638 7 1 2 27606 27637
0 27639 7 1 2 27577 27638
0 27640 5 1 1 27639
0 27641 7 1 2 58897 27640
0 27642 7 1 2 27551 27641
0 27643 5 1 1 27642
0 27644 7 1 2 27494 27643
0 27645 5 1 1 27644
0 27646 7 1 2 43019 27645
0 27647 5 1 1 27646
0 27648 7 1 2 66037 62307
0 27649 5 1 1 27648
0 27650 7 1 2 27647 27649
0 27651 5 1 1 27650
0 27652 7 1 2 46574 27651
0 27653 5 1 1 27652
0 27654 7 1 2 51159 53650
0 27655 7 1 2 56266 27654
0 27656 7 1 2 64286 27655
0 27657 5 1 1 27656
0 27658 7 1 2 62353 57471
0 27659 5 1 1 27658
0 27660 7 1 2 58590 55598
0 27661 5 1 1 27660
0 27662 7 1 2 27659 27661
0 27663 5 1 1 27662
0 27664 7 1 2 50373 27663
0 27665 5 1 1 27664
0 27666 7 1 2 27657 27665
0 27667 5 1 1 27666
0 27668 7 1 2 52008 27667
0 27669 5 1 1 27668
0 27670 7 1 2 42428 58436
0 27671 5 1 1 27670
0 27672 7 1 2 56276 27671
0 27673 5 1 1 27672
0 27674 7 1 2 57997 57692
0 27675 7 1 2 27673 27674
0 27676 5 1 1 27675
0 27677 7 1 2 27669 27676
0 27678 5 1 1 27677
0 27679 7 1 2 41260 27678
0 27680 5 1 1 27679
0 27681 7 1 2 55482 62622
0 27682 5 1 1 27681
0 27683 7 1 2 41393 58694
0 27684 5 1 1 27683
0 27685 7 1 2 58452 27684
0 27686 5 1 1 27685
0 27687 7 1 2 45769 53571
0 27688 5 1 1 27687
0 27689 7 1 2 45979 27688
0 27690 7 1 2 27686 27689
0 27691 5 1 1 27690
0 27692 7 1 2 27682 27691
0 27693 5 1 1 27692
0 27694 7 1 2 57998 53612
0 27695 7 1 2 27693 27694
0 27696 5 1 1 27695
0 27697 7 1 2 27680 27696
0 27698 5 1 1 27697
0 27699 7 1 2 40474 27698
0 27700 5 1 1 27699
0 27701 7 2 2 57999 53651
0 27702 7 2 2 48001 55256
0 27703 7 1 2 40100 66174
0 27704 5 1 1 27703
0 27705 7 1 2 66125 27704
0 27706 5 1 1 27705
0 27707 7 1 2 42429 27706
0 27708 5 1 1 27707
0 27709 7 1 2 44690 55506
0 27710 5 1 1 27709
0 27711 7 1 2 27708 27710
0 27712 5 1 1 27711
0 27713 7 1 2 45328 27712
0 27714 5 1 1 27713
0 27715 7 1 2 27391 27714
0 27716 5 1 1 27715
0 27717 7 1 2 41142 27716
0 27718 5 1 1 27717
0 27719 7 1 2 65923 26573
0 27720 5 1 1 27719
0 27721 7 1 2 46764 27720
0 27722 5 1 1 27721
0 27723 7 1 2 52538 64313
0 27724 7 1 2 23941 27723
0 27725 5 1 1 27724
0 27726 7 1 2 27722 27725
0 27727 7 1 2 27718 27726
0 27728 5 1 1 27727
0 27729 7 1 2 66172 27728
0 27730 5 1 1 27729
0 27731 7 1 2 27700 27730
0 27732 5 1 1 27731
0 27733 7 1 2 40279 27732
0 27734 5 1 1 27733
0 27735 7 2 2 65016 61187
0 27736 5 1 1 66176
0 27737 7 1 2 40101 55257
0 27738 7 1 2 61450 27737
0 27739 5 1 1 27738
0 27740 7 1 2 27736 27739
0 27741 5 1 1 27740
0 27742 7 1 2 46815 27741
0 27743 5 1 1 27742
0 27744 7 1 2 49946 66177
0 27745 5 1 1 27744
0 27746 7 2 2 40475 50848
0 27747 5 3 1 66178
0 27748 7 1 2 66175 66179
0 27749 5 1 1 27748
0 27750 7 1 2 42430 27749
0 27751 7 1 2 27745 27750
0 27752 7 1 2 27743 27751
0 27753 5 1 1 27752
0 27754 7 1 2 66084 63220
0 27755 5 1 1 27754
0 27756 7 1 2 46155 66119
0 27757 5 1 1 27756
0 27758 7 1 2 27755 27757
0 27759 5 1 1 27758
0 27760 7 1 2 42686 27759
0 27761 5 1 1 27760
0 27762 7 2 2 42165 55258
0 27763 7 1 2 41261 66183
0 27764 7 1 2 65720 27763
0 27765 5 1 1 27764
0 27766 7 1 2 45770 27765
0 27767 7 1 2 27761 27766
0 27768 5 1 1 27767
0 27769 7 1 2 66173 27768
0 27770 7 1 2 27753 27769
0 27771 5 1 1 27770
0 27772 7 1 2 27734 27771
0 27773 5 1 1 27772
0 27774 7 1 2 65308 27773
0 27775 5 1 1 27774
0 27776 7 1 2 27653 27775
0 27777 5 1 1 27776
0 27778 7 1 2 43243 27777
0 27779 5 1 1 27778
0 27780 7 1 2 56236 66129
0 27781 5 1 1 27780
0 27782 7 1 2 65526 58827
0 27783 5 1 1 27782
0 27784 7 1 2 27781 27783
0 27785 5 1 1 27784
0 27786 7 1 2 45329 27785
0 27787 5 1 1 27786
0 27788 7 1 2 47092 62204
0 27789 7 1 2 66157 27788
0 27790 5 1 1 27789
0 27791 7 1 2 27787 27790
0 27792 5 1 1 27791
0 27793 7 1 2 43944 44322
0 27794 7 1 2 55085 27793
0 27795 7 1 2 66044 27794
0 27796 7 1 2 27792 27795
0 27797 5 1 1 27796
0 27798 7 1 2 27779 27797
0 27799 7 1 2 27475 27798
0 27800 5 1 1 27799
0 27801 7 1 2 51547 27800
0 27802 5 1 1 27801
0 27803 7 3 2 47093 48828
0 27804 5 1 1 66185
0 27805 7 1 2 27804 61310
0 27806 5 1 1 27805
0 27807 7 2 2 52239 48829
0 27808 5 1 1 66188
0 27809 7 1 2 48395 27808
0 27810 5 1 1 27809
0 27811 7 1 2 43411 27810
0 27812 7 1 2 27806 27811
0 27813 5 1 1 27812
0 27814 7 1 2 49805 66186
0 27815 5 1 1 27814
0 27816 7 1 2 27813 27815
0 27817 5 1 1 27816
0 27818 7 1 2 42687 54983
0 27819 7 1 2 46575 27818
0 27820 7 1 2 27817 27819
0 27821 5 1 1 27820
0 27822 7 2 2 40280 46289
0 27823 7 1 2 53463 64045
0 27824 7 1 2 66190 27823
0 27825 7 1 2 65945 27824
0 27826 7 1 2 65340 27825
0 27827 5 1 1 27826
0 27828 7 1 2 27821 27827
0 27829 5 1 1 27828
0 27830 7 1 2 44816 27829
0 27831 5 1 1 27830
0 27832 7 1 2 65703 49698
0 27833 5 1 1 27832
0 27834 7 1 2 45980 66109
0 27835 5 1 1 27834
0 27836 7 1 2 55449 60902
0 27837 5 1 1 27836
0 27838 7 1 2 27835 27837
0 27839 5 1 1 27838
0 27840 7 1 2 47291 27839
0 27841 5 1 1 27840
0 27842 7 1 2 27833 27841
0 27843 5 1 1 27842
0 27844 7 1 2 65533 64046
0 27845 7 1 2 57958 27844
0 27846 7 1 2 27843 27845
0 27847 5 1 1 27846
0 27848 7 1 2 27831 27847
0 27849 5 1 1 27848
0 27850 7 1 2 43945 27849
0 27851 5 1 1 27850
0 27852 7 1 2 54362 64852
0 27853 5 1 1 27852
0 27854 7 2 2 52460 47558
0 27855 5 1 1 66192
0 27856 7 1 2 50975 58243
0 27857 7 1 2 66193 27856
0 27858 5 1 1 27857
0 27859 7 1 2 27853 27858
0 27860 5 1 1 27859
0 27861 7 2 2 46424 64668
0 27862 7 1 2 46290 56804
0 27863 7 1 2 66194 27862
0 27864 7 1 2 27860 27863
0 27865 5 1 1 27864
0 27866 7 1 2 27851 27865
0 27867 5 1 1 27866
0 27868 7 1 2 42869 27867
0 27869 5 1 1 27868
0 27870 7 1 2 41394 65649
0 27871 5 1 1 27870
0 27872 7 1 2 54533 50632
0 27873 5 1 1 27872
0 27874 7 1 2 27871 27873
0 27875 5 1 1 27874
0 27876 7 1 2 27875 61482
0 27877 5 1 1 27876
0 27878 7 1 2 41143 62744
0 27879 7 1 2 65726 27878
0 27880 5 1 1 27879
0 27881 7 1 2 27877 27880
0 27882 5 1 1 27881
0 27883 7 1 2 46156 65409
0 27884 7 1 2 64047 27883
0 27885 7 1 2 27882 27884
0 27886 5 1 1 27885
0 27887 7 1 2 27869 27886
0 27888 5 1 1 27887
0 27889 7 1 2 55086 27888
0 27890 5 1 1 27889
0 27891 7 1 2 58000 51929
0 27892 5 1 1 27891
0 27893 7 1 2 63911 46894
0 27894 7 1 2 66086 27893
0 27895 5 1 1 27894
0 27896 7 1 2 27892 27895
0 27897 5 1 1 27896
0 27898 7 1 2 40281 27897
0 27899 5 1 1 27898
0 27900 7 1 2 53324 62573
0 27901 7 1 2 62623 27900
0 27902 5 1 1 27901
0 27903 7 1 2 27899 27902
0 27904 5 1 1 27903
0 27905 7 1 2 40102 27904
0 27906 5 1 1 27905
0 27907 7 2 2 51930 46930
0 27908 7 1 2 41526 55767
0 27909 7 1 2 66196 27908
0 27910 5 1 1 27909
0 27911 7 1 2 27906 27910
0 27912 5 1 1 27911
0 27913 7 1 2 41395 27912
0 27914 5 1 1 27913
0 27915 7 1 2 51243 65997
0 27916 5 1 1 27915
0 27917 7 1 2 52514 48167
0 27918 7 1 2 63032 27917
0 27919 5 1 1 27918
0 27920 7 1 2 27916 27919
0 27921 5 1 1 27920
0 27922 7 1 2 40282 27921
0 27923 5 1 1 27922
0 27924 7 1 2 50233 56613
0 27925 7 1 2 65265 27924
0 27926 5 1 1 27925
0 27927 7 1 2 27923 27926
0 27928 5 1 1 27927
0 27929 7 1 2 54363 27928
0 27930 5 1 1 27929
0 27931 7 4 2 42166 54824
0 27932 7 1 2 56721 66198
0 27933 7 1 2 65194 27932
0 27934 5 1 1 27933
0 27935 7 1 2 27930 27934
0 27936 7 1 2 27914 27935
0 27937 5 1 1 27936
0 27938 7 1 2 42870 27937
0 27939 5 1 1 27938
0 27940 7 1 2 65588 56294
0 27941 5 1 1 27940
0 27942 7 1 2 40666 54275
0 27943 5 1 1 27942
0 27944 7 1 2 61147 27943
0 27945 5 4 1 27944
0 27946 7 1 2 51855 64359
0 27947 7 1 2 66202 27946
0 27948 5 1 1 27947
0 27949 7 1 2 27941 27948
0 27950 5 1 1 27949
0 27951 7 1 2 46878 27950
0 27952 5 1 1 27951
0 27953 7 1 2 44817 65195
0 27954 7 1 2 56514 27953
0 27955 5 1 1 27954
0 27956 7 1 2 27952 27955
0 27957 7 1 2 27939 27956
0 27958 5 1 1 27957
0 27959 7 1 2 40476 27958
0 27960 5 1 1 27959
0 27961 7 1 2 49294 63348
0 27962 7 1 2 65936 27961
0 27963 5 1 1 27962
0 27964 7 1 2 47737 54713
0 27965 5 1 1 27964
0 27966 7 1 2 49756 27965
0 27967 5 1 1 27966
0 27968 7 2 2 46157 47420
0 27969 7 1 2 50593 66206
0 27970 7 1 2 27967 27969
0 27971 5 1 1 27970
0 27972 7 1 2 27963 27971
0 27973 5 1 1 27972
0 27974 7 1 2 45330 27973
0 27975 5 1 1 27974
0 27976 7 1 2 45771 56042
0 27977 5 1 1 27976
0 27978 7 1 2 40667 58811
0 27979 5 1 1 27978
0 27980 7 1 2 27977 27979
0 27981 5 1 1 27980
0 27982 7 1 2 43580 27981
0 27983 5 1 1 27982
0 27984 7 1 2 43946 47877
0 27985 5 1 1 27984
0 27986 7 1 2 27983 27985
0 27987 5 1 1 27986
0 27988 7 1 2 47421 59241
0 27989 7 1 2 27987 27988
0 27990 5 1 1 27989
0 27991 7 1 2 27975 27990
0 27992 5 1 1 27991
0 27993 7 1 2 54364 27992
0 27994 5 1 1 27993
0 27995 7 1 2 43947 56295
0 27996 7 1 2 59870 27995
0 27997 5 1 1 27996
0 27998 7 1 2 49889 50594
0 27999 7 1 2 60672 27998
0 28000 5 1 1 27999
0 28001 7 1 2 27997 28000
0 28002 5 1 1 28001
0 28003 7 1 2 45331 28002
0 28004 5 1 1 28003
0 28005 7 1 2 56140 55879
0 28006 5 1 1 28005
0 28007 7 1 2 28004 28006
0 28008 5 1 1 28007
0 28009 7 1 2 65551 28008
0 28010 5 1 1 28009
0 28011 7 3 2 46158 49749
0 28012 7 1 2 49764 66208
0 28013 7 1 2 55551 28012
0 28014 7 1 2 66151 28013
0 28015 5 1 1 28014
0 28016 7 1 2 28010 28015
0 28017 7 1 2 27994 28016
0 28018 7 1 2 27960 28017
0 28019 5 1 1 28018
0 28020 7 1 2 46291 28019
0 28021 5 1 1 28020
0 28022 7 1 2 65589 54932
0 28023 5 1 1 28022
0 28024 7 1 2 64258 28023
0 28025 5 1 1 28024
0 28026 7 1 2 40477 64873
0 28027 7 1 2 28025 28026
0 28028 5 1 1 28027
0 28029 7 1 2 28021 28028
0 28030 5 1 1 28029
0 28031 7 1 2 43132 65317
0 28032 7 1 2 28030 28031
0 28033 5 1 1 28032
0 28034 7 1 2 27890 28033
0 28035 5 1 1 28034
0 28036 7 1 2 43244 28035
0 28037 5 1 1 28036
0 28038 7 3 2 50120 60222
0 28039 7 2 2 48422 66211
0 28040 7 1 2 54434 47852
0 28041 7 1 2 64760 28040
0 28042 7 1 2 66214 28041
0 28043 5 1 1 28042
0 28044 7 1 2 63461 64062
0 28045 7 1 2 61086 28044
0 28046 5 1 1 28045
0 28047 7 1 2 28043 28046
0 28048 5 1 1 28047
0 28049 7 1 2 43020 28048
0 28050 5 1 1 28049
0 28051 7 1 2 47484 65819
0 28052 5 1 1 28051
0 28053 7 1 2 62940 53368
0 28054 5 1 1 28053
0 28055 7 1 2 28052 28054
0 28056 5 1 1 28055
0 28057 7 1 2 42688 28056
0 28058 5 1 1 28057
0 28059 7 1 2 43412 55552
0 28060 5 1 1 28059
0 28061 7 1 2 3417 28060
0 28062 5 1 1 28061
0 28063 7 1 2 52260 28062
0 28064 5 1 1 28063
0 28065 7 1 2 28058 28064
0 28066 5 1 1 28065
0 28067 7 1 2 43749 28066
0 28068 5 1 1 28067
0 28069 7 4 2 40478 44691
0 28070 5 1 1 66216
0 28071 7 1 2 47980 28070
0 28072 5 1 1 28071
0 28073 7 1 2 47422 48864
0 28074 7 1 2 56038 28073
0 28075 7 1 2 28072 28074
0 28076 5 1 1 28075
0 28077 7 1 2 28068 28076
0 28078 5 1 1 28077
0 28079 7 1 2 44530 28078
0 28080 5 1 1 28079
0 28081 7 1 2 42689 58326
0 28082 7 1 2 65396 28081
0 28083 5 1 1 28082
0 28084 7 1 2 28080 28083
0 28085 5 1 1 28084
0 28086 7 1 2 42167 28085
0 28087 5 1 1 28086
0 28088 7 1 2 64974 52528
0 28089 5 1 1 28088
0 28090 7 1 2 28087 28089
0 28091 5 1 1 28090
0 28092 7 1 2 58008 28091
0 28093 5 1 1 28092
0 28094 7 1 2 55152 52529
0 28095 5 1 1 28094
0 28096 7 1 2 45981 62461
0 28097 5 1 1 28096
0 28098 7 1 2 44531 27855
0 28099 7 1 2 28097 28098
0 28100 5 1 1 28099
0 28101 7 1 2 41262 58360
0 28102 5 1 1 28101
0 28103 7 1 2 42168 28102
0 28104 7 1 2 28100 28103
0 28105 5 1 1 28104
0 28106 7 1 2 28095 28105
0 28107 5 1 1 28106
0 28108 7 1 2 41527 28107
0 28109 5 1 1 28108
0 28110 7 1 2 51931 63487
0 28111 7 1 2 65442 28110
0 28112 5 1 1 28111
0 28113 7 1 2 28109 28112
0 28114 5 1 1 28113
0 28115 7 1 2 43750 28114
0 28116 5 1 1 28115
0 28117 7 1 2 54324 50422
0 28118 7 1 2 58371 28117
0 28119 5 1 1 28118
0 28120 7 1 2 44692 28119
0 28121 7 1 2 28116 28120
0 28122 5 1 1 28121
0 28123 7 1 2 58747 64406
0 28124 5 1 1 28123
0 28125 7 1 2 28124 20251
0 28126 5 1 1 28125
0 28127 7 1 2 43413 28126
0 28128 5 1 1 28127
0 28129 7 1 2 58748 66145
0 28130 5 1 1 28129
0 28131 7 1 2 28128 28130
0 28132 5 1 1 28131
0 28133 7 1 2 48377 28132
0 28134 5 1 1 28133
0 28135 7 1 2 50563 64519
0 28136 5 1 1 28135
0 28137 7 1 2 50358 21531
0 28138 5 1 1 28137
0 28139 7 2 2 43751 44818
0 28140 5 1 1 66220
0 28141 7 1 2 47485 28140
0 28142 7 1 2 28138 28141
0 28143 5 1 1 28142
0 28144 7 1 2 28136 28143
0 28145 5 1 1 28144
0 28146 7 1 2 42690 28145
0 28147 5 1 1 28146
0 28148 7 1 2 28134 28147
0 28149 5 1 1 28148
0 28150 7 1 2 47094 28149
0 28151 5 1 1 28150
0 28152 7 1 2 54276 65068
0 28153 5 1 1 28152
0 28154 7 1 2 41396 28153
0 28155 7 1 2 28151 28154
0 28156 5 1 1 28155
0 28157 7 1 2 43948 28156
0 28158 7 1 2 28122 28157
0 28159 5 1 1 28158
0 28160 7 1 2 28093 28159
0 28161 5 1 1 28160
0 28162 7 1 2 46159 28161
0 28163 5 2 1 28162
0 28164 7 1 2 52626 50903
0 28165 5 1 1 28164
0 28166 7 1 2 28165 13706
0 28167 5 1 1 28166
0 28168 7 1 2 41397 28167
0 28169 5 1 1 28168
0 28170 7 2 2 41528 50893
0 28171 7 1 2 52358 66224
0 28172 5 1 1 28171
0 28173 7 1 2 28169 28172
0 28174 5 1 1 28173
0 28175 7 1 2 43581 28174
0 28176 5 1 1 28175
0 28177 7 2 2 40479 65158
0 28178 5 1 1 66226
0 28179 7 1 2 63247 66227
0 28180 5 1 1 28179
0 28181 7 1 2 28176 28180
0 28182 5 1 1 28181
0 28183 7 1 2 43414 28182
0 28184 5 1 1 28183
0 28185 7 1 2 65029 59327
0 28186 5 1 1 28185
0 28187 7 1 2 40480 52261
0 28188 5 1 1 28187
0 28189 7 1 2 28186 28188
0 28190 5 1 1 28189
0 28191 7 1 2 63546 28190
0 28192 5 1 1 28191
0 28193 7 1 2 28184 28192
0 28194 5 1 1 28193
0 28195 7 1 2 40668 28194
0 28196 5 1 1 28195
0 28197 7 1 2 47423 65074
0 28198 7 1 2 51419 28197
0 28199 5 1 1 28198
0 28200 7 1 2 47810 62495
0 28201 5 1 1 28200
0 28202 7 1 2 44819 58217
0 28203 5 1 1 28202
0 28204 7 1 2 47292 21748
0 28205 7 1 2 28203 28204
0 28206 5 1 1 28205
0 28207 7 1 2 28201 28206
0 28208 5 1 1 28207
0 28209 7 1 2 45332 28208
0 28210 5 1 1 28209
0 28211 7 1 2 40481 49380
0 28212 7 1 2 65503 28211
0 28213 5 1 1 28212
0 28214 7 1 2 28210 28213
0 28215 5 1 1 28214
0 28216 7 1 2 45502 28215
0 28217 5 1 1 28216
0 28218 7 1 2 28199 28217
0 28219 5 1 1 28218
0 28220 7 1 2 50779 28219
0 28221 5 1 1 28220
0 28222 7 1 2 28196 28221
0 28223 5 1 1 28222
0 28224 7 1 2 45982 28223
0 28225 5 1 1 28224
0 28226 7 1 2 58026 61416
0 28227 7 1 2 63514 28226
0 28228 5 1 1 28227
0 28229 7 1 2 28225 28228
0 28230 5 1 1 28229
0 28231 7 1 2 45772 28230
0 28232 5 1 1 28231
0 28233 7 2 2 56237 65387
0 28234 7 1 2 65577 66228
0 28235 5 1 1 28234
0 28236 7 1 2 28232 28235
0 28237 5 1 1 28236
0 28238 7 1 2 42871 28237
0 28239 5 1 1 28238
0 28240 7 1 2 66222 28239
0 28241 5 1 1 28240
0 28242 7 1 2 54616 28241
0 28243 5 1 1 28242
0 28244 7 1 2 28050 28243
0 28245 5 1 1 28244
0 28246 7 1 2 65103 28245
0 28247 5 1 1 28246
0 28248 7 1 2 28037 28247
0 28249 5 1 1 28248
0 28250 7 1 2 48078 28249
0 28251 5 1 1 28250
0 28252 7 1 2 65485 63000
0 28253 5 1 1 28252
0 28254 7 1 2 64835 63786
0 28255 5 1 1 28254
0 28256 7 1 2 28253 28255
0 28257 5 1 1 28256
0 28258 7 1 2 44820 28257
0 28259 5 1 1 28258
0 28260 7 1 2 44124 46720
0 28261 7 1 2 60883 28260
0 28262 7 1 2 50307 57228
0 28263 7 1 2 28261 28262
0 28264 5 1 1 28263
0 28265 7 1 2 28259 28264
0 28266 5 1 1 28265
0 28267 7 1 2 43949 28266
0 28268 5 1 1 28267
0 28269 7 2 2 44821 60974
0 28270 7 1 2 63001 66230
0 28271 7 1 2 61062 28270
0 28272 5 1 1 28271
0 28273 7 1 2 28268 28272
0 28274 5 1 1 28273
0 28275 7 1 2 46160 28274
0 28276 5 1 1 28275
0 28277 7 3 2 46425 64836
0 28278 7 1 2 62754 57235
0 28279 7 1 2 53332 28278
0 28280 7 1 2 66232 28279
0 28281 5 1 1 28280
0 28282 7 1 2 28276 28281
0 28283 5 1 1 28282
0 28284 7 1 2 45173 28283
0 28285 5 1 1 28284
0 28286 7 2 2 48129 60369
0 28287 7 2 2 3961 66235
0 28288 7 1 2 49604 59566
0 28289 7 1 2 66237 28288
0 28290 5 1 1 28289
0 28291 7 1 2 28285 28290
0 28292 5 1 1 28291
0 28293 7 1 2 44323 28292
0 28294 5 1 1 28293
0 28295 7 1 2 46542 51698
0 28296 7 1 2 66238 28295
0 28297 5 1 1 28296
0 28298 7 1 2 28294 28297
0 28299 5 1 1 28298
0 28300 7 1 2 55087 28299
0 28301 5 1 1 28300
0 28302 7 1 2 53652 59741
0 28303 7 2 2 60849 28302
0 28304 5 1 1 66239
0 28305 7 1 2 65398 66240
0 28306 5 1 1 28305
0 28307 7 1 2 45174 28306
0 28308 5 1 1 28307
0 28309 7 3 2 60370 59395
0 28310 5 1 1 66241
0 28311 7 1 2 28304 28310
0 28312 5 1 1 28311
0 28313 7 1 2 47486 28312
0 28314 7 1 2 28308 28313
0 28315 5 1 1 28314
0 28316 7 1 2 46509 62297
0 28317 5 1 1 28316
0 28318 7 1 2 59742 28317
0 28319 7 1 2 57818 28318
0 28320 5 1 1 28319
0 28321 7 3 2 54617 59702
0 28322 7 1 2 63094 66244
0 28323 5 1 1 28322
0 28324 7 1 2 28320 28323
0 28325 7 1 2 28315 28324
0 28326 5 1 1 28325
0 28327 7 1 2 43752 28326
0 28328 5 1 1 28327
0 28329 7 1 2 65239 65451
0 28330 5 1 1 28329
0 28331 7 4 2 43753 41847
0 28332 7 1 2 66247 62742
0 28333 5 1 1 28332
0 28334 7 1 2 28330 28333
0 28335 5 1 1 28334
0 28336 7 1 2 64289 28335
0 28337 5 1 1 28336
0 28338 7 2 2 47859 51308
0 28339 7 1 2 45333 66245
0 28340 7 1 2 66251 28339
0 28341 5 1 1 28340
0 28342 7 1 2 28337 28341
0 28343 7 1 2 28328 28342
0 28344 5 1 1 28343
0 28345 7 1 2 45503 28344
0 28346 5 1 1 28345
0 28347 7 1 2 63467 57423
0 28348 5 1 1 28347
0 28349 7 1 2 28348 64116
0 28350 5 1 1 28349
0 28351 7 1 2 42169 28350
0 28352 5 1 1 28351
0 28353 7 1 2 48079 63368
0 28354 5 2 1 28353
0 28355 7 2 2 53653 58946
0 28356 7 1 2 54480 66255
0 28357 5 1 1 28356
0 28358 7 1 2 66253 28357
0 28359 5 1 1 28358
0 28360 7 1 2 47487 28359
0 28361 5 1 1 28360
0 28362 7 1 2 28352 28361
0 28363 5 1 1 28362
0 28364 7 1 2 47811 28363
0 28365 5 1 1 28364
0 28366 7 1 2 62648 57822
0 28367 5 1 1 28366
0 28368 7 1 2 43021 59976
0 28369 7 1 2 62198 28368
0 28370 5 1 1 28369
0 28371 7 1 2 28367 28370
0 28372 5 1 1 28371
0 28373 7 1 2 40482 28372
0 28374 5 1 1 28373
0 28375 7 2 2 53667 61190
0 28376 5 1 1 66257
0 28377 7 1 2 66254 28376
0 28378 5 1 1 28377
0 28379 7 1 2 47599 28378
0 28380 5 1 1 28379
0 28381 7 2 2 64279 63668
0 28382 7 1 2 46953 54618
0 28383 7 1 2 66259 28382
0 28384 5 1 1 28383
0 28385 7 1 2 28380 28384
0 28386 7 1 2 28374 28385
0 28387 7 1 2 28365 28386
0 28388 5 1 1 28387
0 28389 7 1 2 59703 28388
0 28390 5 1 1 28389
0 28391 7 1 2 44125 43022
0 28392 7 6 2 46426 28391
0 28393 7 1 2 44964 45175
0 28394 7 1 2 65121 28393
0 28395 7 1 2 66261 28394
0 28396 7 1 2 65249 28395
0 28397 5 1 1 28396
0 28398 7 1 2 28390 28397
0 28399 7 1 2 28346 28398
0 28400 5 1 1 28399
0 28401 7 1 2 44822 28400
0 28402 5 1 1 28401
0 28403 7 3 2 43415 49806
0 28404 7 1 2 58799 62976
0 28405 7 2 2 66267 28404
0 28406 7 5 2 44532 41529
0 28407 7 1 2 65174 66272
0 28408 7 1 2 48317 28407
0 28409 7 1 2 66270 28408
0 28410 5 1 1 28409
0 28411 7 1 2 28402 28410
0 28412 5 1 1 28411
0 28413 7 1 2 43950 28412
0 28414 5 1 1 28413
0 28415 7 1 2 45176 58009
0 28416 7 1 2 51548 28415
0 28417 7 1 2 47195 28416
0 28418 7 1 2 66271 28417
0 28419 5 1 1 28418
0 28420 7 1 2 28414 28419
0 28421 5 1 1 28420
0 28422 7 1 2 46161 28421
0 28423 5 1 1 28422
0 28424 7 1 2 45504 54719
0 28425 5 1 1 28424
0 28426 7 2 2 64888 28425
0 28427 5 1 1 66277
0 28428 7 1 2 64902 66278
0 28429 5 1 1 28428
0 28430 7 1 2 59704 28429
0 28431 5 1 1 28430
0 28432 7 1 2 59534 65481
0 28433 5 1 1 28432
0 28434 7 1 2 59535 65471
0 28435 5 1 1 28434
0 28436 7 1 2 59705 62649
0 28437 5 1 1 28436
0 28438 7 1 2 28435 28437
0 28439 5 1 1 28438
0 28440 7 1 2 40483 28439
0 28441 5 1 1 28440
0 28442 7 1 2 28433 28441
0 28443 7 1 2 28431 28442
0 28444 5 1 1 28443
0 28445 7 1 2 56862 57823
0 28446 7 1 2 28444 28445
0 28447 5 1 1 28446
0 28448 7 1 2 28423 28447
0 28449 5 1 1 28448
0 28450 7 1 2 44324 28449
0 28451 5 1 1 28450
0 28452 7 1 2 43023 49144
0 28453 7 1 2 66233 28452
0 28454 5 1 1 28453
0 28455 7 1 2 56991 57824
0 28456 7 1 2 64908 28455
0 28457 5 1 1 28456
0 28458 7 1 2 28454 28457
0 28459 5 2 1 28458
0 28460 7 1 2 65226 66279
0 28461 5 1 1 28460
0 28462 7 1 2 28451 28461
0 28463 5 1 1 28462
0 28464 7 1 2 57650 28463
0 28465 5 1 1 28464
0 28466 7 1 2 65215 66280
0 28467 5 1 1 28466
0 28468 7 1 2 28465 28467
0 28469 7 1 2 28301 28468
0 28470 5 1 1 28469
0 28471 7 1 2 53763 28470
0 28472 5 1 1 28471
0 28473 7 1 2 28251 28472
0 28474 7 1 2 27802 28473
0 28475 5 1 1 28474
0 28476 7 1 2 49039 28475
0 28477 5 1 1 28476
0 28478 7 1 2 54334 10815
0 28479 5 2 1 28478
0 28480 7 1 2 62827 64015
0 28481 5 1 1 28480
0 28482 7 1 2 57651 54619
0 28483 7 1 2 55165 28482
0 28484 5 1 1 28483
0 28485 7 1 2 28481 28484
0 28486 5 1 1 28485
0 28487 7 9 2 46510 65087
0 28488 7 2 2 64669 66283
0 28489 7 1 2 62519 66292
0 28490 7 1 2 28486 28489
0 28491 5 1 1 28490
0 28492 7 3 2 57266 55373
0 28493 7 2 2 65355 66294
0 28494 5 1 1 66297
0 28495 7 2 2 43245 65306
0 28496 5 1 1 66299
0 28497 7 1 2 57810 66300
0 28498 5 1 1 28497
0 28499 7 1 2 65309 51549
0 28500 7 1 2 63433 28499
0 28501 5 1 1 28500
0 28502 7 1 2 28498 28501
0 28503 5 2 1 28502
0 28504 7 1 2 49040 66301
0 28505 5 1 1 28504
0 28506 7 1 2 28494 28505
0 28507 5 1 1 28506
0 28508 7 1 2 49757 61510
0 28509 7 1 2 28507 28508
0 28510 5 1 1 28509
0 28511 7 1 2 28491 28510
0 28512 5 1 1 28511
0 28513 7 1 2 66281 28512
0 28514 5 1 1 28513
0 28515 7 1 2 59056 66199
0 28516 5 1 1 28515
0 28517 7 1 2 42691 59944
0 28518 5 1 1 28517
0 28519 7 1 2 28516 28518
0 28520 5 1 1 28519
0 28521 7 1 2 44533 28520
0 28522 5 1 1 28521
0 28523 7 1 2 40669 41816
0 28524 7 1 2 60217 28523
0 28525 5 1 1 28524
0 28526 7 1 2 28522 28525
0 28527 5 1 1 28526
0 28528 7 1 2 56755 28527
0 28529 5 1 1 28528
0 28530 7 1 2 47054 54505
0 28531 7 1 2 56583 51094
0 28532 7 1 2 28530 28531
0 28533 7 1 2 53996 28532
0 28534 5 1 1 28533
0 28535 7 1 2 28529 28534
0 28536 5 1 1 28535
0 28537 7 1 2 43024 28536
0 28538 5 1 1 28537
0 28539 7 1 2 45983 58800
0 28540 7 1 2 51550 56043
0 28541 7 2 2 28539 28540
0 28542 7 1 2 45115 49355
0 28543 7 1 2 66303 28542
0 28544 5 1 1 28543
0 28545 7 1 2 28538 28544
0 28546 5 1 1 28545
0 28547 7 1 2 44275 28546
0 28548 5 1 1 28547
0 28549 7 1 2 50963 55870
0 28550 5 2 1 28549
0 28551 7 1 2 59089 58723
0 28552 7 1 2 66305 28551
0 28553 7 1 2 56756 28552
0 28554 5 1 1 28553
0 28555 7 1 2 28548 28554
0 28556 5 1 1 28555
0 28557 7 1 2 43416 28556
0 28558 5 1 1 28557
0 28559 7 4 2 43951 47095
0 28560 7 1 2 58591 66307
0 28561 7 1 2 59019 28560
0 28562 5 1 1 28561
0 28563 7 1 2 28558 28562
0 28564 5 1 1 28563
0 28565 7 1 2 46576 28564
0 28566 5 1 1 28565
0 28567 7 1 2 40965 50022
0 28568 5 1 1 28567
0 28569 7 1 2 4678 28568
0 28570 5 2 1 28569
0 28571 7 1 2 45116 66311
0 28572 5 1 1 28571
0 28573 7 1 2 48929 59938
0 28574 5 1 1 28573
0 28575 7 1 2 28572 28574
0 28576 5 1 1 28575
0 28577 7 2 2 46427 66200
0 28578 7 1 2 28576 66313
0 28579 5 1 1 28578
0 28580 7 1 2 59286 58724
0 28581 7 1 2 57063 28580
0 28582 5 1 1 28581
0 28583 7 1 2 28579 28582
0 28584 5 1 1 28583
0 28585 7 1 2 44534 28584
0 28586 5 1 1 28585
0 28587 7 2 2 50911 59911
0 28588 7 1 2 64511 66315
0 28589 5 1 1 28588
0 28590 7 1 2 28586 28589
0 28591 5 1 1 28590
0 28592 7 1 2 48080 28591
0 28593 5 1 1 28592
0 28594 7 1 2 40966 52867
0 28595 5 1 1 28594
0 28596 7 1 2 44216 50023
0 28597 5 1 1 28596
0 28598 7 1 2 28595 28597
0 28599 5 2 1 28598
0 28600 7 1 2 41817 66317
0 28601 5 1 1 28600
0 28602 7 1 2 53921 59363
0 28603 5 1 1 28602
0 28604 7 1 2 28601 28603
0 28605 5 1 1 28604
0 28606 7 1 2 66304 28605
0 28607 5 1 1 28606
0 28608 7 1 2 28593 28607
0 28609 5 1 1 28608
0 28610 7 1 2 41030 28609
0 28611 5 1 1 28610
0 28612 7 1 2 48081 66312
0 28613 5 1 1 28612
0 28614 7 1 2 28613 18595
0 28615 5 2 1 28614
0 28616 7 3 2 44535 41818
0 28617 7 2 2 44276 66321
0 28618 7 1 2 66314 66324
0 28619 7 1 2 66319 28618
0 28620 5 1 1 28619
0 28621 7 1 2 28611 28620
0 28622 5 1 1 28621
0 28623 7 1 2 43417 28622
0 28624 5 1 1 28623
0 28625 7 2 2 52188 66322
0 28626 7 1 2 63154 66326
0 28627 7 1 2 58843 28626
0 28628 5 1 1 28627
0 28629 7 1 2 28624 28628
0 28630 5 1 1 28629
0 28631 7 1 2 64670 28630
0 28632 5 1 1 28631
0 28633 7 1 2 28566 28632
0 28634 5 1 1 28633
0 28635 7 2 2 43754 43246
0 28636 7 1 2 41530 66328
0 28637 7 1 2 28634 28636
0 28638 5 1 1 28637
0 28639 7 1 2 28514 28638
0 28640 5 1 1 28639
0 28641 7 1 2 42431 28640
0 28642 5 1 1 28641
0 28643 7 15 2 43247 65318
0 28644 7 2 2 57811 66330
0 28645 5 1 1 66345
0 28646 7 2 2 47096 66346
0 28647 5 1 1 66347
0 28648 7 2 2 55866 63314
0 28649 7 2 2 54620 65487
0 28650 7 1 2 66349 66351
0 28651 5 1 1 28650
0 28652 7 1 2 28645 28651
0 28653 5 2 1 28652
0 28654 7 1 2 43755 66353
0 28655 5 1 1 28654
0 28656 7 1 2 28647 28655
0 28657 5 1 1 28656
0 28658 7 1 2 49041 28657
0 28659 5 1 1 28658
0 28660 7 1 2 47149 66298
0 28661 5 1 1 28660
0 28662 7 2 2 62804 63419
0 28663 7 1 2 64671 55867
0 28664 7 1 2 58865 28663
0 28665 7 1 2 66355 28664
0 28666 5 1 1 28665
0 28667 7 1 2 28661 28666
0 28668 7 1 2 28659 28667
0 28669 5 1 1 28668
0 28670 7 2 2 58027 28669
0 28671 5 1 1 66357
0 28672 7 1 2 55088 56757
0 28673 5 1 1 28672
0 28674 7 1 2 28673 17680
0 28675 5 2 1 28674
0 28676 7 1 2 46577 66359
0 28677 5 1 1 28676
0 28678 7 3 2 48082 64672
0 28679 7 1 2 61978 66361
0 28680 5 1 1 28679
0 28681 7 1 2 28677 28680
0 28682 5 1 1 28681
0 28683 7 1 2 43952 66273
0 28684 7 1 2 64536 28683
0 28685 7 1 2 28682 28684
0 28686 5 1 1 28685
0 28687 7 1 2 28671 28686
0 28688 5 1 1 28687
0 28689 7 1 2 60919 28688
0 28690 5 1 1 28689
0 28691 7 1 2 28642 28690
0 28692 5 1 1 28691
0 28693 7 1 2 44693 28692
0 28694 5 1 1 28693
0 28695 7 1 2 42432 66358
0 28696 5 1 1 28695
0 28697 7 1 2 59607 63534
0 28698 5 1 1 28697
0 28699 7 2 2 58177 56972
0 28700 7 1 2 53307 66364
0 28701 7 1 2 63536 28700
0 28702 5 1 1 28701
0 28703 7 1 2 28698 28702
0 28704 5 1 1 28703
0 28705 7 1 2 55089 28704
0 28706 5 1 1 28705
0 28707 7 1 2 62732 66295
0 28708 5 1 1 28707
0 28709 7 2 2 55176 54638
0 28710 7 2 2 44277 59322
0 28711 7 2 2 65714 66368
0 28712 7 1 2 46511 66370
0 28713 7 1 2 66366 28712
0 28714 5 1 1 28713
0 28715 7 1 2 28708 28714
0 28716 7 1 2 28706 28715
0 28717 5 1 1 28716
0 28718 7 1 2 45177 28717
0 28719 5 1 1 28718
0 28720 7 2 2 59300 63627
0 28721 7 1 2 63775 66372
0 28722 5 1 1 28721
0 28723 7 1 2 28719 28722
0 28724 5 1 1 28723
0 28725 7 1 2 44325 28724
0 28726 5 1 1 28725
0 28727 7 1 2 65351 66296
0 28728 5 1 1 28727
0 28729 7 1 2 49042 66354
0 28730 5 1 1 28729
0 28731 7 1 2 28728 28730
0 28732 7 1 2 28726 28731
0 28733 5 2 1 28732
0 28734 7 3 2 43953 65445
0 28735 7 1 2 55002 66376
0 28736 7 1 2 66374 28735
0 28737 5 1 1 28736
0 28738 7 1 2 28696 28737
0 28739 5 1 1 28738
0 28740 7 1 2 41398 28739
0 28741 5 1 1 28740
0 28742 7 2 2 58010 53673
0 28743 7 1 2 63814 66379
0 28744 5 1 1 28743
0 28745 7 1 2 58001 50595
0 28746 7 1 2 58898 28745
0 28747 5 1 1 28746
0 28748 7 1 2 28744 28747
0 28749 5 1 1 28748
0 28750 7 1 2 46578 28749
0 28751 5 1 1 28750
0 28752 7 1 2 65310 66231
0 28753 7 1 2 62173 28752
0 28754 5 1 1 28753
0 28755 7 1 2 28751 28754
0 28756 5 1 1 28755
0 28757 7 1 2 56758 28756
0 28758 5 1 1 28757
0 28759 7 1 2 66380 59144
0 28760 5 1 1 28759
0 28761 7 2 2 61897 59287
0 28762 5 1 1 66381
0 28763 7 1 2 43954 62273
0 28764 7 1 2 66382 28763
0 28765 5 1 1 28764
0 28766 7 1 2 28760 28765
0 28767 5 1 1 28766
0 28768 7 1 2 45178 28767
0 28769 5 1 1 28768
0 28770 7 1 2 53035 61934
0 28771 7 1 2 59301 56843
0 28772 7 1 2 28770 28771
0 28773 5 1 1 28772
0 28774 7 1 2 28769 28773
0 28775 5 1 1 28774
0 28776 7 1 2 44326 28775
0 28777 5 1 1 28776
0 28778 7 2 2 46543 61935
0 28779 7 1 2 65329 64597
0 28780 7 1 2 66383 28779
0 28781 5 1 1 28780
0 28782 7 1 2 28777 28781
0 28783 5 1 1 28782
0 28784 7 1 2 56568 28783
0 28785 5 1 1 28784
0 28786 7 1 2 28758 28785
0 28787 5 1 1 28786
0 28788 7 1 2 49385 63075
0 28789 7 1 2 28787 28788
0 28790 5 1 1 28789
0 28791 7 1 2 28741 28790
0 28792 5 1 1 28791
0 28793 7 1 2 42692 28792
0 28794 5 1 1 28793
0 28795 7 1 2 28694 28794
0 28796 5 1 1 28795
0 28797 7 1 2 46162 28796
0 28798 5 1 1 28797
0 28799 7 1 2 59958 50948
0 28800 5 1 1 28799
0 28801 7 1 2 61521 59407
0 28802 5 1 1 28801
0 28803 7 1 2 28800 28802
0 28804 5 1 1 28803
0 28805 7 1 2 48830 28804
0 28806 5 1 1 28805
0 28807 7 1 2 62174 64598
0 28808 5 1 1 28807
0 28809 7 1 2 28806 28808
0 28810 5 1 1 28809
0 28811 7 1 2 56940 28810
0 28812 5 1 1 28811
0 28813 7 1 2 45117 60668
0 28814 7 2 2 62162 28813
0 28815 7 1 2 57859 66385
0 28816 5 1 1 28815
0 28817 7 1 2 43133 50663
0 28818 7 1 2 62720 28817
0 28819 5 1 1 28818
0 28820 7 1 2 28816 28819
0 28821 5 1 1 28820
0 28822 7 1 2 60048 28821
0 28823 5 1 1 28822
0 28824 7 1 2 28812 28823
0 28825 5 1 1 28824
0 28826 7 1 2 44278 28825
0 28827 5 1 1 28826
0 28828 7 3 2 42170 56332
0 28829 7 1 2 45058 57146
0 28830 7 1 2 66387 28829
0 28831 5 1 1 28830
0 28832 7 1 2 43418 63114
0 28833 7 1 2 56941 28832
0 28834 5 1 1 28833
0 28835 7 1 2 28831 28834
0 28836 5 1 1 28835
0 28837 7 1 2 59090 28836
0 28838 5 1 1 28837
0 28839 7 1 2 28827 28838
0 28840 5 1 1 28839
0 28841 7 1 2 49249 28840
0 28842 5 1 1 28841
0 28843 7 2 2 54079 62905
0 28844 7 1 2 57017 66390
0 28845 5 1 1 28844
0 28846 7 1 2 58840 28845
0 28847 5 1 1 28846
0 28848 7 1 2 45118 28847
0 28849 5 1 1 28848
0 28850 7 1 2 43134 63987
0 28851 5 2 1 28850
0 28852 7 1 2 28849 66392
0 28853 5 1 1 28852
0 28854 7 1 2 44279 28853
0 28855 5 1 1 28854
0 28856 7 1 2 59091 59015
0 28857 5 2 1 28856
0 28858 7 1 2 28855 66394
0 28859 5 1 1 28858
0 28860 7 2 2 40670 48831
0 28861 5 2 1 66396
0 28862 7 1 2 50668 66398
0 28863 5 6 1 28862
0 28864 7 1 2 46292 66400
0 28865 7 1 2 28859 28864
0 28866 5 1 1 28865
0 28867 7 1 2 56906 62691
0 28868 7 1 2 59110 62746
0 28869 7 1 2 28867 28868
0 28870 5 1 1 28869
0 28871 7 1 2 28866 28870
0 28872 5 1 1 28871
0 28873 7 1 2 52691 28872
0 28874 5 1 1 28873
0 28875 7 1 2 28842 28874
0 28876 5 1 1 28875
0 28877 7 1 2 43756 28876
0 28878 5 1 1 28877
0 28879 7 2 2 49043 59417
0 28880 7 1 2 53704 54726
0 28881 7 1 2 56558 28880
0 28882 7 1 2 66406 28881
0 28883 5 1 1 28882
0 28884 7 1 2 28878 28883
0 28885 5 1 1 28884
0 28886 7 1 2 44536 28885
0 28887 5 1 1 28886
0 28888 7 1 2 54806 60581
0 28889 7 1 2 58774 28888
0 28890 7 1 2 62702 28889
0 28891 7 1 2 66407 28890
0 28892 5 1 1 28891
0 28893 7 1 2 28887 28892
0 28894 5 1 1 28893
0 28895 7 1 2 46579 28894
0 28896 5 1 1 28895
0 28897 7 5 2 43419 46428
0 28898 7 2 2 55090 66408
0 28899 5 1 1 66413
0 28900 7 1 2 6893 28899
0 28901 5 1 1 28900
0 28902 7 2 2 46293 28901
0 28903 7 1 2 49094 66415
0 28904 5 1 1 28903
0 28905 7 1 2 56663 63764
0 28906 5 1 1 28905
0 28907 7 1 2 28904 28906
0 28908 5 1 1 28907
0 28909 7 1 2 40876 28908
0 28910 5 1 1 28909
0 28911 7 1 2 48590 58686
0 28912 7 1 2 63056 28911
0 28913 5 1 1 28912
0 28914 7 1 2 28910 28913
0 28915 5 1 1 28914
0 28916 7 1 2 49044 28915
0 28917 5 1 1 28916
0 28918 7 2 2 55091 52929
0 28919 7 1 2 53922 66417
0 28920 5 1 1 28919
0 28921 7 1 2 21370 28920
0 28922 5 1 1 28921
0 28923 7 1 2 66409 28922
0 28924 5 1 1 28923
0 28925 7 2 2 56682 59274
0 28926 5 1 1 66419
0 28927 7 1 2 66420 62864
0 28928 5 1 1 28927
0 28929 7 1 2 28924 28928
0 28930 5 1 1 28929
0 28931 7 1 2 56352 28930
0 28932 5 1 1 28931
0 28933 7 1 2 28917 28932
0 28934 5 1 1 28933
0 28935 7 1 2 66401 28934
0 28936 5 1 1 28935
0 28937 7 1 2 50664 57064
0 28938 5 1 1 28937
0 28939 7 3 2 43420 61880
0 28940 7 1 2 51426 57860
0 28941 7 1 2 66421 28940
0 28942 5 1 1 28941
0 28943 7 1 2 28938 28942
0 28944 5 1 1 28943
0 28945 7 1 2 64618 28944
0 28946 5 1 1 28945
0 28947 7 1 2 54727 54925
0 28948 7 1 2 58207 28947
0 28949 5 1 1 28948
0 28950 7 1 2 28946 28949
0 28951 5 1 1 28950
0 28952 7 1 2 41819 28951
0 28953 5 1 1 28952
0 28954 7 1 2 48226 57861
0 28955 7 1 2 51432 28954
0 28956 7 4 2 43421 51458
0 28957 7 1 2 59224 66424
0 28958 7 1 2 28955 28957
0 28959 5 1 1 28958
0 28960 7 1 2 28953 28959
0 28961 5 1 1 28960
0 28962 7 1 2 41031 28961
0 28963 5 1 1 28962
0 28964 7 1 2 62884 57728
0 28965 7 1 2 60153 28964
0 28966 7 1 2 62779 56094
0 28967 7 1 2 66425 28966
0 28968 7 1 2 28965 28967
0 28969 5 1 1 28968
0 28970 7 1 2 28963 28969
0 28971 7 1 2 28936 28970
0 28972 5 1 1 28971
0 28973 7 1 2 52240 64673
0 28974 7 1 2 28972 28973
0 28975 5 1 1 28974
0 28976 7 1 2 28896 28975
0 28977 5 1 1 28976
0 28978 7 1 2 43248 28977
0 28979 5 1 1 28978
0 28980 7 1 2 43422 62874
0 28981 5 1 1 28980
0 28982 7 1 2 28981 14723
0 28983 5 1 1 28982
0 28984 7 1 2 43249 28983
0 28985 5 1 1 28984
0 28986 7 5 2 43025 66284
0 28987 7 3 2 43423 44280
0 28988 7 2 2 42872 63734
0 28989 7 1 2 66433 66436
0 28990 7 1 2 66428 28989
0 28991 5 1 1 28990
0 28992 7 1 2 28985 28991
0 28993 5 1 1 28992
0 28994 7 1 2 46429 28993
0 28995 5 1 1 28994
0 28996 7 1 2 63057 62773
0 28997 5 1 1 28996
0 28998 7 1 2 28995 28997
0 28999 5 1 1 28998
0 29000 7 1 2 49045 28999
0 29001 5 1 1 29000
0 29002 7 3 2 53654 66285
0 29003 7 2 2 46163 63105
0 29004 7 1 2 59005 50643
0 29005 7 1 2 66441 29004
0 29006 7 1 2 66438 29005
0 29007 5 1 1 29006
0 29008 7 1 2 29001 29007
0 29009 5 1 1 29008
0 29010 7 1 2 45179 29009
0 29011 5 1 1 29010
0 29012 7 2 2 63199 64728
0 29013 7 1 2 59307 66443
0 29014 5 1 1 29013
0 29015 7 1 2 29011 29014
0 29016 5 1 1 29015
0 29017 7 1 2 44327 29016
0 29018 5 1 1 29017
0 29019 7 4 2 66023 59595
0 29020 7 1 2 66444 66445
0 29021 5 1 1 29020
0 29022 7 1 2 29018 29021
0 29023 5 1 1 29022
0 29024 7 1 2 55949 53693
0 29025 7 1 2 500 5234
0 29026 7 1 2 29024 29025
0 29027 7 1 2 29023 29026
0 29028 5 1 1 29027
0 29029 7 2 2 56079 53435
0 29030 5 1 1 66449
0 29031 7 1 2 48344 49837
0 29032 5 1 1 29031
0 29033 7 1 2 29030 29032
0 29034 5 4 1 29033
0 29035 7 2 2 43135 66451
0 29036 7 1 2 66455 60131
0 29037 5 1 1 29036
0 29038 7 1 2 56523 50074
0 29039 5 1 1 29038
0 29040 7 2 2 46164 53436
0 29041 7 1 2 54921 66457
0 29042 5 1 1 29041
0 29043 7 1 2 29039 29042
0 29044 5 1 1 29043
0 29045 7 1 2 66098 49374
0 29046 7 1 2 29044 29045
0 29047 5 1 1 29046
0 29048 7 1 2 29037 29047
0 29049 5 1 1 29048
0 29050 7 1 2 44328 29049
0 29051 5 1 1 29050
0 29052 7 2 2 45059 46544
0 29053 7 1 2 57018 66459
0 29054 7 1 2 66456 29053
0 29055 5 1 1 29054
0 29056 7 1 2 29051 29055
0 29057 5 1 1 29056
0 29058 7 1 2 51273 29057
0 29059 5 1 1 29058
0 29060 7 3 2 40967 51459
0 29061 7 1 2 52009 64674
0 29062 7 2 2 66461 29061
0 29063 7 1 2 53613 52233
0 29064 7 1 2 66464 29063
0 29065 5 1 1 29064
0 29066 7 1 2 29059 29065
0 29067 5 1 1 29066
0 29068 7 1 2 55092 29067
0 29069 5 1 1 29068
0 29070 7 1 2 51295 66458
0 29071 5 1 1 29070
0 29072 7 1 2 49838 56606
0 29073 5 1 1 29072
0 29074 7 1 2 29071 29073
0 29075 5 1 1 29074
0 29076 7 1 2 66391 29075
0 29077 5 1 1 29076
0 29078 7 1 2 66450 57116
0 29079 5 1 1 29078
0 29080 7 1 2 29077 29079
0 29081 5 1 1 29080
0 29082 7 1 2 40877 29081
0 29083 5 1 1 29082
0 29084 7 1 2 49839 50614
0 29085 7 1 2 59074 29084
0 29086 5 1 1 29085
0 29087 7 1 2 29083 29086
0 29088 5 1 1 29087
0 29089 7 1 2 44217 29088
0 29090 5 1 1 29089
0 29091 7 2 2 56227 57187
0 29092 5 2 1 66466
0 29093 7 1 2 56383 51666
0 29094 7 1 2 66467 29093
0 29095 5 1 1 29094
0 29096 7 1 2 29090 29095
0 29097 5 1 1 29096
0 29098 7 1 2 65319 29097
0 29099 5 1 1 29098
0 29100 7 1 2 29069 29099
0 29101 5 1 1 29100
0 29102 7 1 2 43250 29101
0 29103 5 1 1 29102
0 29104 7 1 2 55177 56524
0 29105 5 1 1 29104
0 29106 7 1 2 52010 64125
0 29107 5 1 1 29106
0 29108 7 1 2 29105 29107
0 29109 5 1 1 29108
0 29110 7 1 2 54688 52650
0 29111 5 1 1 29110
0 29112 7 1 2 6001 29111
0 29113 5 1 1 29112
0 29114 7 1 2 65320 29113
0 29115 5 1 1 29114
0 29116 7 1 2 65144 57959
0 29117 7 1 2 64577 29116
0 29118 7 1 2 66418 29117
0 29119 5 1 1 29118
0 29120 7 1 2 29115 29119
0 29121 5 1 1 29120
0 29122 7 1 2 43251 29121
0 29123 5 1 1 29122
0 29124 7 1 2 65508 52930
0 29125 5 1 1 29124
0 29126 7 1 2 29125 28926
0 29127 5 1 1 29126
0 29128 7 1 2 52868 29127
0 29129 5 1 1 29128
0 29130 7 1 2 57117 64558
0 29131 5 1 1 29130
0 29132 7 1 2 29129 29131
0 29133 5 1 1 29132
0 29134 7 1 2 44281 29133
0 29135 5 1 1 29134
0 29136 7 1 2 59186 46692
0 29137 7 2 2 63971 29136
0 29138 5 1 1 66470
0 29139 7 1 2 43136 66471
0 29140 5 1 1 29139
0 29141 7 1 2 29135 29140
0 29142 5 1 1 29141
0 29143 7 1 2 66293 29142
0 29144 5 1 1 29143
0 29145 7 1 2 29123 29144
0 29146 5 1 1 29145
0 29147 7 1 2 29109 29146
0 29148 5 1 1 29147
0 29149 7 1 2 43137 52011
0 29150 7 1 2 64039 29149
0 29151 5 1 1 29150
0 29152 7 1 2 48832 54585
0 29153 7 1 2 62692 29152
0 29154 5 1 1 29153
0 29155 7 1 2 29151 29154
0 29156 5 1 1 29155
0 29157 7 1 2 49985 29156
0 29158 7 1 2 66331 29157
0 29159 5 1 1 29158
0 29160 7 1 2 42433 66024
0 29161 7 2 2 66439 29160
0 29162 7 4 2 44282 44329
0 29163 7 2 2 57019 66474
0 29164 7 1 2 56057 54728
0 29165 7 1 2 66478 29164
0 29166 7 1 2 66472 29165
0 29167 5 1 1 29166
0 29168 7 1 2 29159 29167
0 29169 5 1 1 29168
0 29170 7 1 2 52931 29169
0 29171 5 1 1 29170
0 29172 7 1 2 66442 57440
0 29173 5 1 1 29172
0 29174 7 1 2 29173 63966
0 29175 5 1 1 29174
0 29176 7 1 2 44283 29175
0 29177 5 1 1 29176
0 29178 7 2 2 63735 59121
0 29179 7 1 2 48591 66480
0 29180 5 2 1 29179
0 29181 7 1 2 29177 66482
0 29182 5 1 1 29181
0 29183 7 1 2 49046 29182
0 29184 5 1 1 29183
0 29185 7 1 2 62805 63691
0 29186 5 1 1 29185
0 29187 7 1 2 29184 29186
0 29188 5 1 1 29187
0 29189 7 2 2 65159 64052
0 29190 7 1 2 56819 65540
0 29191 7 1 2 66484 29190
0 29192 7 1 2 29188 29191
0 29193 5 1 1 29192
0 29194 7 1 2 29171 29193
0 29195 7 1 2 29148 29194
0 29196 7 1 2 29103 29195
0 29197 7 1 2 29028 29196
0 29198 5 1 1 29197
0 29199 7 1 2 40484 29198
0 29200 5 1 1 29199
0 29201 7 1 2 66308 55788
0 29202 5 1 1 29201
0 29203 7 1 2 44126 61774
0 29204 5 1 1 29203
0 29205 7 1 2 29202 29204
0 29206 5 1 1 29205
0 29207 7 1 2 66410 29206
0 29208 7 1 2 65359 29207
0 29209 5 1 1 29208
0 29210 7 2 2 62828 66286
0 29211 7 2 2 66013 64048
0 29212 7 1 2 66488 53265
0 29213 7 1 2 66486 29212
0 29214 5 1 1 29213
0 29215 7 1 2 29209 29214
0 29216 5 1 1 29215
0 29217 7 1 2 45773 29216
0 29218 5 1 1 29217
0 29219 7 2 2 48833 62520
0 29220 5 1 1 66490
0 29221 7 1 2 45180 59759
0 29222 7 1 2 66491 29221
0 29223 7 1 2 66487 29222
0 29224 5 1 1 29223
0 29225 7 1 2 29218 29224
0 29226 5 1 1 29225
0 29227 7 1 2 48277 29226
0 29228 5 1 1 29227
0 29229 7 2 2 60223 62175
0 29230 7 1 2 65795 66492
0 29231 5 1 1 29230
0 29232 7 2 2 42434 61356
0 29233 7 1 2 64053 66217
0 29234 7 1 2 66494 29233
0 29235 5 1 1 29234
0 29236 7 1 2 29231 29235
0 29237 5 1 1 29236
0 29238 7 1 2 44537 29237
0 29239 5 1 1 29238
0 29240 7 1 2 42171 59728
0 29241 7 1 2 66218 29240
0 29242 7 1 2 66495 29241
0 29243 5 1 1 29242
0 29244 7 1 2 29239 29243
0 29245 5 1 1 29244
0 29246 7 1 2 44330 29245
0 29247 5 1 1 29246
0 29248 7 1 2 60231 59596
0 29249 7 3 2 45119 65382
0 29250 7 1 2 63896 66496
0 29251 7 1 2 29248 29250
0 29252 5 1 1 29251
0 29253 7 1 2 29247 29252
0 29254 5 1 1 29253
0 29255 7 1 2 62681 29254
0 29256 5 1 1 29255
0 29257 7 1 2 65088 62245
0 29258 5 1 1 29257
0 29259 7 1 2 43252 66414
0 29260 5 1 1 29259
0 29261 7 1 2 29258 29260
0 29262 5 1 1 29261
0 29263 7 1 2 40485 66465
0 29264 7 1 2 29262 29263
0 29265 5 1 1 29264
0 29266 7 1 2 29256 29265
0 29267 5 1 1 29266
0 29268 7 1 2 52771 29267
0 29269 5 1 1 29268
0 29270 7 1 2 29228 29269
0 29271 7 1 2 29200 29270
0 29272 7 1 2 28979 29271
0 29273 5 1 1 29272
0 29274 7 1 2 54365 29273
0 29275 5 1 1 29274
0 29276 7 1 2 60224 54446
0 29277 7 1 2 56113 29276
0 29278 5 1 1 29277
0 29279 7 1 2 44965 56152
0 29280 7 1 2 63026 29279
0 29281 5 1 1 29280
0 29282 7 1 2 29278 29281
0 29283 5 1 1 29282
0 29284 7 1 2 61357 29283
0 29285 5 1 1 29284
0 29286 7 2 2 57267 65205
0 29287 7 2 2 66323 66499
0 29288 7 1 2 64398 61248
0 29289 7 1 2 66501 29288
0 29290 5 1 1 29289
0 29291 7 1 2 29285 29290
0 29292 5 1 1 29291
0 29293 7 1 2 43026 29292
0 29294 5 1 1 29293
0 29295 7 3 2 43424 49750
0 29296 7 1 2 51274 59122
0 29297 7 1 2 66503 29296
0 29298 7 1 2 66502 29297
0 29299 5 1 1 29298
0 29300 7 1 2 29294 29299
0 29301 5 1 1 29300
0 29302 7 1 2 45181 29301
0 29303 5 1 1 29302
0 29304 7 2 2 62906 56353
0 29305 5 1 1 66506
0 29306 7 1 2 55385 29305
0 29307 5 2 1 29306
0 29308 7 1 2 59302 56044
0 29309 7 1 2 59024 29308
0 29310 7 1 2 66500 29309
0 29311 7 1 2 66508 29310
0 29312 5 1 1 29311
0 29313 7 1 2 29303 29312
0 29314 5 1 1 29313
0 29315 7 1 2 44823 29314
0 29316 5 1 1 29315
0 29317 7 2 2 65796 53668
0 29318 7 1 2 46979 53464
0 29319 7 1 2 56961 29318
0 29320 7 1 2 66510 29319
0 29321 5 1 1 29320
0 29322 7 1 2 29316 29321
0 29323 5 1 1 29322
0 29324 7 1 2 42172 29323
0 29325 5 1 1 29324
0 29326 7 2 2 66006 57210
0 29327 7 1 2 66350 66512
0 29328 5 1 1 29327
0 29329 7 1 2 44127 66511
0 29330 5 1 1 29329
0 29331 7 1 2 29328 29330
0 29332 5 1 1 29331
0 29333 7 2 2 65570 54113
0 29334 7 1 2 29332 66514
0 29335 5 1 1 29334
0 29336 7 1 2 29325 29335
0 29337 5 1 1 29336
0 29338 7 1 2 44331 29337
0 29339 5 1 1 29338
0 29340 7 3 2 53266 50401
0 29341 7 1 2 64176 66516
0 29342 5 1 1 29341
0 29343 7 1 2 54277 56525
0 29344 7 1 2 66509 29343
0 29345 5 1 1 29344
0 29346 7 1 2 29342 29345
0 29347 5 1 1 29346
0 29348 7 1 2 52359 29347
0 29349 5 1 1 29348
0 29350 7 1 2 64177 58002
0 29351 7 1 2 64756 29350
0 29352 5 1 1 29351
0 29353 7 1 2 29349 29352
0 29354 5 1 1 29353
0 29355 7 1 2 65227 58914
0 29356 7 1 2 29354 29355
0 29357 5 1 1 29356
0 29358 7 1 2 29339 29357
0 29359 5 1 1 29358
0 29360 7 1 2 49047 29359
0 29361 5 1 1 29360
0 29362 7 1 2 56722 56003
0 29363 7 2 2 63776 29362
0 29364 7 1 2 56342 66519
0 29365 5 1 1 29364
0 29366 7 1 2 15149 63794
0 29367 5 2 1 29366
0 29368 7 1 2 54278 64939
0 29369 7 1 2 54957 29368
0 29370 7 1 2 66521 29369
0 29371 5 1 1 29370
0 29372 7 1 2 29365 29371
0 29373 5 1 1 29372
0 29374 7 1 2 53923 29373
0 29375 5 1 1 29374
0 29376 7 1 2 63237 65160
0 29377 7 1 2 50968 29376
0 29378 7 1 2 63520 56790
0 29379 7 1 2 29377 29378
0 29380 5 1 1 29379
0 29381 7 1 2 29375 29380
0 29382 5 1 1 29381
0 29383 7 1 2 43955 29382
0 29384 5 1 1 29383
0 29385 7 1 2 46980 63916
0 29386 5 1 1 29385
0 29387 7 1 2 50752 52964
0 29388 7 1 2 63521 29387
0 29389 5 1 1 29388
0 29390 7 1 2 29386 29389
0 29391 5 1 1 29390
0 29392 7 1 2 48083 50955
0 29393 7 1 2 64178 29392
0 29394 7 1 2 29391 29393
0 29395 5 1 1 29394
0 29396 7 1 2 29384 29395
0 29397 5 1 1 29396
0 29398 7 1 2 45182 29397
0 29399 5 1 1 29398
0 29400 7 2 2 59919 63707
0 29401 7 1 2 60129 57268
0 29402 7 1 2 51234 29401
0 29403 7 1 2 58777 29402
0 29404 7 1 2 66523 29403
0 29405 5 1 1 29404
0 29406 7 1 2 29399 29405
0 29407 5 1 1 29406
0 29408 7 1 2 44332 29407
0 29409 5 1 1 29408
0 29410 7 3 2 43757 45183
0 29411 7 3 2 41053 66525
0 29412 7 3 2 44538 66528
0 29413 7 1 2 54543 63434
0 29414 7 1 2 63708 51441
0 29415 7 1 2 29413 29414
0 29416 7 1 2 66531 29415
0 29417 5 1 1 29416
0 29418 7 1 2 29409 29417
0 29419 5 1 1 29418
0 29420 7 1 2 55093 29419
0 29421 5 1 1 29420
0 29422 7 1 2 57652 66532
0 29423 5 1 1 29422
0 29424 7 1 2 44333 46981
0 29425 7 1 2 60081 29424
0 29426 5 1 1 29425
0 29427 7 1 2 29423 29426
0 29428 5 1 1 29427
0 29429 7 1 2 60749 66522
0 29430 5 1 1 29429
0 29431 7 1 2 57269 63961
0 29432 5 1 1 29431
0 29433 7 1 2 29430 29432
0 29434 5 1 1 29433
0 29435 7 2 2 54534 29434
0 29436 7 1 2 61140 66534
0 29437 5 1 1 29436
0 29438 7 1 2 45060 64126
0 29439 7 1 2 66520 29438
0 29440 5 1 1 29439
0 29441 7 1 2 29437 29440
0 29442 5 1 1 29441
0 29443 7 1 2 29428 29442
0 29444 5 1 1 29443
0 29445 7 1 2 44539 65182
0 29446 7 1 2 63435 29445
0 29447 7 3 2 43758 49118
0 29448 7 1 2 60847 66536
0 29449 7 1 2 29446 29448
0 29450 5 1 1 29449
0 29451 7 1 2 48084 56445
0 29452 7 1 2 54991 29451
0 29453 5 1 1 29452
0 29454 7 2 2 42693 57960
0 29455 7 2 2 60690 66539
0 29456 7 1 2 44966 61528
0 29457 7 1 2 66541 29456
0 29458 5 1 1 29457
0 29459 7 1 2 29453 29458
0 29460 5 1 1 29459
0 29461 7 2 2 46512 59729
0 29462 7 1 2 48709 66543
0 29463 7 1 2 29460 29462
0 29464 5 1 1 29463
0 29465 7 1 2 29450 29464
0 29466 5 1 1 29465
0 29467 7 1 2 56384 29466
0 29468 5 1 1 29467
0 29469 7 1 2 43759 65168
0 29470 7 1 2 56049 29469
0 29471 7 1 2 66535 29470
0 29472 5 1 1 29471
0 29473 7 1 2 29468 29472
0 29474 5 1 1 29473
0 29475 7 1 2 65234 29474
0 29476 5 1 1 29475
0 29477 7 1 2 29444 29476
0 29478 5 1 1 29477
0 29479 7 1 2 42173 29478
0 29480 5 1 1 29479
0 29481 7 2 2 53655 66332
0 29482 7 1 2 56746 66545
0 29483 5 1 1 29482
0 29484 7 1 2 45505 65431
0 29485 7 1 2 58178 57729
0 29486 7 1 2 29484 29485
0 29487 7 1 2 65235 63537
0 29488 7 1 2 29486 29487
0 29489 5 1 1 29488
0 29490 7 1 2 29483 29489
0 29491 5 1 1 29490
0 29492 7 1 2 66515 29491
0 29493 5 1 1 29492
0 29494 7 1 2 29480 29493
0 29495 7 1 2 29421 29494
0 29496 7 1 2 29361 29495
0 29497 5 1 1 29496
0 29498 7 1 2 42873 29497
0 29499 5 1 1 29498
0 29500 7 2 2 55094 53705
0 29501 7 2 2 57223 66547
0 29502 7 1 2 60691 66549
0 29503 5 1 1 29502
0 29504 7 1 2 57653 48168
0 29505 7 1 2 57236 55789
0 29506 7 1 2 29504 29505
0 29507 5 1 1 29506
0 29508 7 1 2 29503 29507
0 29509 5 1 1 29508
0 29510 7 1 2 49048 29509
0 29511 5 1 1 29510
0 29512 7 1 2 58866 66388
0 29513 5 1 1 29512
0 29514 7 1 2 51309 48402
0 29515 7 1 2 53706 29514
0 29516 5 1 1 29515
0 29517 7 1 2 29513 29516
0 29518 5 1 1 29517
0 29519 7 1 2 62806 29518
0 29520 5 1 1 29519
0 29521 7 1 2 29511 29520
0 29522 5 1 1 29521
0 29523 7 1 2 40671 29522
0 29524 5 1 1 29523
0 29525 7 1 2 51087 50923
0 29526 7 1 2 57441 29525
0 29527 7 1 2 62807 29526
0 29528 5 1 1 29527
0 29529 7 1 2 29524 29528
0 29530 5 1 1 29529
0 29531 7 1 2 43138 29530
0 29532 5 1 1 29531
0 29533 7 2 2 43956 49215
0 29534 7 2 2 48834 66551
0 29535 5 1 1 66553
0 29536 7 1 2 46294 60750
0 29537 5 1 1 29536
0 29538 7 1 2 5290 29537
0 29539 5 1 1 29538
0 29540 7 1 2 66554 29539
0 29541 5 1 1 29540
0 29542 7 1 2 44128 66422
0 29543 7 1 2 56376 29542
0 29544 5 1 1 29543
0 29545 7 1 2 29541 29544
0 29546 5 1 1 29545
0 29547 7 1 2 54040 58915
0 29548 7 1 2 29546 29547
0 29549 5 1 1 29548
0 29550 7 1 2 29532 29549
0 29551 5 1 1 29550
0 29552 7 1 2 46580 29551
0 29553 5 1 1 29552
0 29554 7 1 2 41676 56385
0 29555 7 1 2 66416 29554
0 29556 5 1 1 29555
0 29557 7 1 2 49840 53669
0 29558 7 1 2 59525 29557
0 29559 5 1 1 29558
0 29560 7 1 2 29556 29559
0 29561 5 1 1 29560
0 29562 7 1 2 40878 29561
0 29563 5 1 1 29562
0 29564 7 1 2 53036 46635
0 29565 7 1 2 50135 29564
0 29566 7 1 2 66262 29565
0 29567 5 1 1 29566
0 29568 7 1 2 29563 29567
0 29569 5 1 1 29568
0 29570 7 1 2 49049 29569
0 29571 5 1 1 29570
0 29572 7 1 2 43425 64703
0 29573 5 1 1 29572
0 29574 7 1 2 61851 29573
0 29575 5 1 1 29574
0 29576 7 1 2 50095 62384
0 29577 5 1 1 29576
0 29578 7 1 2 29535 29577
0 29579 5 1 1 29578
0 29580 7 1 2 46295 29579
0 29581 7 1 2 29575 29580
0 29582 5 1 1 29581
0 29583 7 1 2 29571 29582
0 29584 5 1 1 29583
0 29585 7 1 2 54041 29584
0 29586 5 1 1 29585
0 29587 7 1 2 60669 50009
0 29588 7 1 2 53707 29587
0 29589 7 1 2 58419 59608
0 29590 7 1 2 29588 29589
0 29591 5 1 1 29590
0 29592 7 1 2 29586 29591
0 29593 5 1 1 29592
0 29594 7 1 2 64675 29593
0 29595 5 1 1 29594
0 29596 7 1 2 29553 29595
0 29597 5 1 1 29596
0 29598 7 1 2 44540 43253
0 29599 7 1 2 29597 29598
0 29600 5 1 1 29599
0 29601 7 1 2 65941 66399
0 29602 5 4 1 29601
0 29603 7 2 2 40486 66555
0 29604 7 1 2 59706 57427
0 29605 5 2 1 29604
0 29606 7 1 2 60049 63142
0 29607 5 1 1 29606
0 29608 7 1 2 65089 55374
0 29609 5 1 1 29608
0 29610 7 1 2 29607 29609
0 29611 5 1 1 29610
0 29612 7 1 2 59536 29611
0 29613 5 1 1 29612
0 29614 7 1 2 66561 29613
0 29615 5 1 1 29614
0 29616 7 1 2 59086 29615
0 29617 5 1 1 29616
0 29618 7 2 2 43254 60078
0 29619 7 1 2 46430 66563
0 29620 7 1 2 66507 29619
0 29621 5 1 1 29620
0 29622 7 1 2 29617 29621
0 29623 5 1 1 29622
0 29624 7 1 2 44334 29623
0 29625 5 1 1 29624
0 29626 7 1 2 46545 60371
0 29627 7 1 2 51551 59364
0 29628 7 1 2 29626 29627
0 29629 5 1 1 29628
0 29630 7 1 2 29625 29629
0 29631 5 1 1 29630
0 29632 7 1 2 62838 29631
0 29633 5 1 1 29632
0 29634 7 1 2 66429 59613
0 29635 5 1 1 29634
0 29636 7 1 2 29635 66562
0 29637 5 1 1 29636
0 29638 7 1 2 44335 29637
0 29639 5 1 1 29638
0 29640 7 3 2 45184 62765
0 29641 7 1 2 59317 66565
0 29642 5 1 1 29641
0 29643 7 1 2 29639 29642
0 29644 5 1 1 29643
0 29645 7 1 2 62847 29644
0 29646 5 1 1 29645
0 29647 7 1 2 64655 55182
0 29648 7 1 2 66566 29647
0 29649 5 1 1 29648
0 29650 7 1 2 29646 29649
0 29651 5 1 1 29650
0 29652 7 1 2 65511 29651
0 29653 5 1 1 29652
0 29654 7 1 2 44336 62844
0 29655 7 1 2 64016 66544
0 29656 7 1 2 60019 29655
0 29657 7 1 2 29654 29656
0 29658 5 1 1 29657
0 29659 7 1 2 29653 29658
0 29660 7 1 2 29633 29659
0 29661 7 1 2 66246 63315
0 29662 5 1 1 29661
0 29663 7 1 2 41032 59516
0 29664 5 1 1 29663
0 29665 7 1 2 57224 59064
0 29666 7 1 2 66287 29665
0 29667 5 1 1 29666
0 29668 7 1 2 29664 29667
0 29669 5 1 1 29668
0 29670 7 1 2 65512 29669
0 29671 5 1 1 29670
0 29672 7 1 2 53561 61548
0 29673 5 1 1 29672
0 29674 7 1 2 29673 12112
0 29675 5 1 1 29674
0 29676 7 1 2 57237 60343
0 29677 7 1 2 29675 29676
0 29678 5 1 1 29677
0 29679 7 2 2 57293 65090
0 29680 7 1 2 66481 66568
0 29681 5 1 1 29680
0 29682 7 1 2 29678 29681
0 29683 7 1 2 29671 29682
0 29684 5 1 1 29683
0 29685 7 1 2 45185 29684
0 29686 5 1 1 29685
0 29687 7 1 2 29662 29686
0 29688 5 1 1 29687
0 29689 7 1 2 44337 29688
0 29690 5 1 1 29689
0 29691 7 2 2 66025 60344
0 29692 7 1 2 41677 54621
0 29693 7 1 2 59383 29692
0 29694 7 1 2 66570 29693
0 29695 5 1 1 29694
0 29696 7 1 2 29690 29695
0 29697 5 1 1 29696
0 29698 7 1 2 49050 29697
0 29699 5 1 1 29698
0 29700 7 1 2 66375 66397
0 29701 5 1 1 29700
0 29702 7 1 2 29699 29701
0 29703 7 1 2 29660 29702
0 29704 5 1 1 29703
0 29705 7 1 2 66559 29704
0 29706 5 1 1 29705
0 29707 7 1 2 29600 29706
0 29708 5 1 1 29707
0 29709 7 1 2 65552 29708
0 29710 5 1 1 29709
0 29711 7 3 2 59959 59707
0 29712 7 1 2 53216 66572
0 29713 5 1 1 29712
0 29714 7 1 2 54325 65091
0 29715 7 1 2 66100 29714
0 29716 5 1 1 29715
0 29717 7 1 2 29713 29716
0 29718 5 1 1 29717
0 29719 7 1 2 64507 29718
0 29720 5 1 1 29719
0 29721 7 1 2 43760 66146
0 29722 7 1 2 66573 29721
0 29723 5 1 1 29722
0 29724 7 1 2 29720 29723
0 29725 5 1 1 29724
0 29726 7 1 2 43957 29725
0 29727 5 1 1 29726
0 29728 7 2 2 43139 64968
0 29729 7 1 2 60975 59708
0 29730 7 1 2 66575 29729
0 29731 7 1 2 58173 29730
0 29732 5 1 1 29731
0 29733 7 1 2 29727 29732
0 29734 5 1 1 29733
0 29735 7 1 2 44694 29734
0 29736 5 1 1 29735
0 29737 7 2 2 46513 58028
0 29738 7 1 2 50290 65145
0 29739 7 1 2 62868 29738
0 29740 7 1 2 66577 29739
0 29741 5 1 1 29740
0 29742 7 1 2 58011 48169
0 29743 7 1 2 66574 29742
0 29744 5 1 1 29743
0 29745 7 1 2 29741 29744
0 29746 5 1 1 29745
0 29747 7 1 2 46982 29746
0 29748 5 1 1 29747
0 29749 7 1 2 59571 62355
0 29750 7 1 2 62527 29749
0 29751 5 1 1 29750
0 29752 7 1 2 29748 29751
0 29753 5 1 1 29752
0 29754 7 1 2 42694 29753
0 29755 5 1 1 29754
0 29756 7 1 2 29736 29755
0 29757 5 1 1 29756
0 29758 7 1 2 48227 29757
0 29759 5 1 1 29758
0 29760 7 1 2 53481 66377
0 29761 7 1 2 66485 64627
0 29762 7 1 2 29760 29761
0 29763 5 1 1 29762
0 29764 7 1 2 29759 29763
0 29765 5 1 1 29764
0 29766 7 1 2 44338 29765
0 29767 5 1 1 29766
0 29768 7 1 2 66062 59190
0 29769 5 1 1 29768
0 29770 7 1 2 60976 29769
0 29771 5 1 1 29770
0 29772 7 1 2 62521 53764
0 29773 5 2 1 29772
0 29774 7 1 2 29771 66579
0 29775 5 1 1 29774
0 29776 7 1 2 44824 29775
0 29777 5 1 1 29776
0 29778 7 1 2 66147 63176
0 29779 5 1 1 29778
0 29780 7 1 2 29777 29779
0 29781 5 3 1 29780
0 29782 7 1 2 46546 63951
0 29783 7 1 2 65177 29782
0 29784 7 1 2 66581 29783
0 29785 5 1 1 29784
0 29786 7 1 2 29767 29785
0 29787 5 1 1 29786
0 29788 7 1 2 44284 29787
0 29789 5 1 1 29788
0 29790 7 1 2 55020 46581
0 29791 7 1 2 63625 29790
0 29792 7 1 2 66582 29791
0 29793 5 1 1 29792
0 29794 7 1 2 29789 29793
0 29795 5 1 1 29794
0 29796 7 1 2 48930 29795
0 29797 5 1 1 29796
0 29798 7 2 2 54279 48228
0 29799 5 1 1 66584
0 29800 7 1 2 57350 29799
0 29801 5 7 1 29800
0 29802 7 1 2 61619 60156
0 29803 5 1 1 29802
0 29804 7 1 2 63577 66288
0 29805 5 1 1 29804
0 29806 7 1 2 29803 29805
0 29807 5 1 1 29806
0 29808 7 1 2 55095 29807
0 29809 5 1 1 29808
0 29810 7 1 2 44541 59497
0 29811 5 1 1 29810
0 29812 7 1 2 62467 29811
0 29813 7 1 2 61634 29812
0 29814 5 1 1 29813
0 29815 7 1 2 62133 66289
0 29816 5 1 1 29815
0 29817 7 1 2 29814 29816
0 29818 7 1 2 29809 29817
0 29819 5 1 1 29818
0 29820 7 1 2 45186 29819
0 29821 5 1 1 29820
0 29822 7 2 2 59709 62860
0 29823 5 2 1 66593
0 29824 7 1 2 43426 66594
0 29825 5 1 1 29824
0 29826 7 1 2 29821 29825
0 29827 5 1 1 29826
0 29828 7 1 2 44339 29827
0 29829 5 1 1 29828
0 29830 7 2 2 48931 63106
0 29831 7 1 2 65125 59597
0 29832 7 1 2 66597 29831
0 29833 5 1 1 29832
0 29834 7 1 2 29829 29833
0 29835 5 1 1 29834
0 29836 7 1 2 66556 29835
0 29837 5 1 1 29836
0 29838 7 1 2 61870 66475
0 29839 7 1 2 64980 29838
0 29840 7 1 2 65345 66423
0 29841 7 1 2 29839 29840
0 29842 5 1 1 29841
0 29843 7 1 2 29837 29842
0 29844 5 1 1 29843
0 29845 7 1 2 40487 29844
0 29846 5 1 1 29845
0 29847 7 1 2 62441 66493
0 29848 7 1 2 65360 29847
0 29849 5 1 1 29848
0 29850 7 1 2 29846 29849
0 29851 5 1 1 29850
0 29852 7 1 2 66586 29851
0 29853 5 1 1 29852
0 29854 7 12 2 43255 46582
0 29855 7 2 2 40672 62645
0 29856 7 1 2 52461 66611
0 29857 5 1 1 29856
0 29858 7 1 2 54825 47055
0 29859 7 1 2 50345 16915
0 29860 7 1 2 29858 29859
0 29861 5 1 1 29860
0 29862 7 1 2 29857 29861
0 29863 5 1 1 29862
0 29864 7 1 2 44695 29863
0 29865 5 1 1 29864
0 29866 7 1 2 65151 66612
0 29867 5 1 1 29866
0 29868 7 1 2 29865 29867
0 29869 5 1 1 29868
0 29870 7 1 2 66599 29869
0 29871 5 1 1 29870
0 29872 7 1 2 54326 65488
0 29873 7 1 2 64948 29872
0 29874 5 1 1 29873
0 29875 7 1 2 29871 29874
0 29876 5 1 1 29875
0 29877 7 1 2 43427 29876
0 29878 5 1 1 29877
0 29879 7 3 2 44340 44696
0 29880 7 1 2 45774 66613
0 29881 7 1 2 66526 29880
0 29882 7 1 2 66111 29881
0 29883 7 1 2 66578 29882
0 29884 5 1 1 29883
0 29885 7 1 2 29878 29884
0 29886 5 1 1 29885
0 29887 7 1 2 56559 29886
0 29888 5 1 1 29887
0 29889 7 1 2 65534 65424
0 29890 7 1 2 56119 29889
0 29891 7 1 2 57301 62703
0 29892 7 1 2 29890 29891
0 29893 5 1 1 29892
0 29894 7 1 2 29888 29893
0 29895 5 1 1 29894
0 29896 7 1 2 55096 29895
0 29897 5 1 1 29896
0 29898 7 4 2 43428 41531
0 29899 7 1 2 57302 66616
0 29900 7 1 2 66557 29899
0 29901 5 1 1 29900
0 29902 7 1 2 56526 50623
0 29903 7 1 2 66569 29902
0 29904 5 1 1 29903
0 29905 7 1 2 29901 29904
0 29906 5 1 1 29905
0 29907 7 1 2 45984 29906
0 29908 5 1 1 29907
0 29909 7 1 2 50300 56050
0 29910 7 1 2 63831 29909
0 29911 5 1 1 29910
0 29912 7 1 2 29908 29911
0 29913 5 1 1 29912
0 29914 7 1 2 55097 29913
0 29915 5 1 1 29914
0 29916 7 3 2 54622 60297
0 29917 7 2 2 53437 48784
0 29918 7 1 2 52692 66623
0 29919 7 1 2 66282 29918
0 29920 7 1 2 66620 29919
0 29921 5 1 1 29920
0 29922 7 1 2 29915 29921
0 29923 5 1 1 29922
0 29924 7 1 2 64676 29923
0 29925 5 1 1 29924
0 29926 7 1 2 65146 66290
0 29927 5 1 1 29926
0 29928 7 1 2 59723 29927
0 29929 5 1 1 29928
0 29930 7 1 2 44341 29929
0 29931 5 1 1 29930
0 29932 7 1 2 23773 29931
0 29933 5 1 1 29932
0 29934 7 1 2 57654 29933
0 29935 5 1 1 29934
0 29936 7 1 2 65219 29935
0 29937 5 1 1 29936
0 29938 7 3 2 54280 53614
0 29939 5 1 1 66625
0 29940 7 1 2 57493 29939
0 29941 5 4 1 29940
0 29942 7 1 2 66558 66628
0 29943 7 1 2 29937 29942
0 29944 5 1 1 29943
0 29945 7 1 2 29925 29944
0 29946 5 1 1 29945
0 29947 7 1 2 40488 29946
0 29948 5 1 1 29947
0 29949 7 1 2 62578 60355
0 29950 7 1 2 65321 29949
0 29951 7 1 2 66629 29950
0 29952 5 1 1 29951
0 29953 7 1 2 29948 29952
0 29954 7 1 2 29897 29953
0 29955 5 1 1 29954
0 29956 7 1 2 49051 29955
0 29957 5 1 1 29956
0 29958 7 1 2 48229 53997
0 29959 7 1 2 66333 29958
0 29960 7 1 2 66583 29959
0 29961 5 1 1 29960
0 29962 7 1 2 29957 29961
0 29963 7 1 2 29853 29962
0 29964 7 1 2 29797 29963
0 29965 5 1 1 29964
0 29966 7 1 2 49216 29965
0 29967 5 1 1 29966
0 29968 7 1 2 29710 29967
0 29969 7 1 2 29499 29968
0 29970 7 1 2 29275 29969
0 29971 7 1 2 28798 29970
0 29972 5 1 1 29971
0 29973 7 1 2 49324 29972
0 29974 5 1 1 29973
0 29975 7 1 2 47738 65882
0 29976 5 1 1 29975
0 29977 7 1 2 53998 65504
0 29978 5 1 1 29977
0 29979 7 1 2 29976 29978
0 29980 5 1 1 29979
0 29981 7 1 2 45775 29980
0 29982 5 1 1 29981
0 29983 7 1 2 65695 57862
0 29984 5 1 1 29983
0 29985 7 1 2 29982 29984
0 29986 5 1 1 29985
0 29987 7 1 2 41981 29986
0 29988 5 1 1 29987
0 29989 7 2 2 43429 40283
0 29990 7 1 2 56547 66632
0 29991 5 1 1 29990
0 29992 7 1 2 52404 60774
0 29993 5 1 1 29992
0 29994 7 1 2 44542 49687
0 29995 5 1 1 29994
0 29996 7 1 2 29993 29995
0 29997 5 1 1 29996
0 29998 7 1 2 42435 29997
0 29999 5 1 1 29998
0 30000 7 1 2 50239 4535
0 30001 5 1 1 30000
0 30002 7 1 2 43430 30001
0 30003 7 1 2 64621 30002
0 30004 5 1 1 30003
0 30005 7 1 2 29999 30004
0 30006 5 1 1 30005
0 30007 7 1 2 45334 30006
0 30008 5 1 1 30007
0 30009 7 1 2 29991 30008
0 30010 5 1 1 30009
0 30011 7 1 2 54178 30010
0 30012 5 1 1 30011
0 30013 7 1 2 29988 30012
0 30014 5 1 1 30013
0 30015 7 1 2 41399 30014
0 30016 5 1 1 30015
0 30017 7 1 2 47534 46774
0 30018 5 1 1 30017
0 30019 7 1 2 46900 46866
0 30020 5 1 1 30019
0 30021 7 1 2 30018 30020
0 30022 5 1 1 30021
0 30023 7 1 2 44697 60860
0 30024 7 1 2 30022 30023
0 30025 5 1 1 30024
0 30026 7 1 2 13433 30025
0 30027 5 1 1 30026
0 30028 7 1 2 40284 30027
0 30029 5 1 1 30028
0 30030 7 1 2 54098 62387
0 30031 7 1 2 59265 30030
0 30032 5 1 1 30031
0 30033 7 1 2 30029 30032
0 30034 7 1 2 30016 30033
0 30035 5 1 1 30034
0 30036 7 1 2 59537 30035
0 30037 5 1 1 30036
0 30038 7 2 2 57842 63596
0 30039 5 1 1 66634
0 30040 7 1 2 46765 57098
0 30041 5 1 1 30040
0 30042 7 1 2 66635 30041
0 30043 5 1 1 30042
0 30044 7 2 2 61316 30043
0 30045 7 1 2 41848 47600
0 30046 7 1 2 66636 30045
0 30047 5 1 1 30046
0 30048 7 1 2 30037 30047
0 30049 5 1 1 30048
0 30050 7 1 2 44342 30049
0 30051 5 1 1 30050
0 30052 7 1 2 46547 47601
0 30053 7 1 2 66637 30052
0 30054 5 1 1 30053
0 30055 7 1 2 30051 30054
0 30056 5 1 1 30055
0 30057 7 1 2 42695 30056
0 30058 5 1 1 30057
0 30059 7 2 2 44543 65883
0 30060 5 1 1 66638
0 30061 7 1 2 54029 30060
0 30062 5 1 1 30061
0 30063 7 1 2 50553 30062
0 30064 5 1 1 30063
0 30065 7 1 2 44544 60737
0 30066 5 1 1 30065
0 30067 7 1 2 30064 30066
0 30068 5 1 1 30067
0 30069 7 1 2 41982 30068
0 30070 5 1 1 30069
0 30071 7 1 2 57836 66411
0 30072 7 1 2 54796 30071
0 30073 5 1 1 30072
0 30074 7 1 2 30070 30073
0 30075 5 1 1 30074
0 30076 7 1 2 53746 65364
0 30077 7 1 2 30075 30076
0 30078 5 1 1 30077
0 30079 7 1 2 30058 30078
0 30080 5 1 1 30079
0 30081 7 1 2 48230 30080
0 30082 5 1 1 30081
0 30083 7 1 2 57081 25771
0 30084 5 1 1 30083
0 30085 7 1 2 66600 30084
0 30086 5 1 1 30085
0 30087 7 1 2 41144 65489
0 30088 7 1 2 63594 30087
0 30089 5 1 1 30088
0 30090 7 1 2 30086 30089
0 30091 5 1 1 30090
0 30092 7 1 2 45335 30091
0 30093 5 1 1 30092
0 30094 7 2 2 46431 66601
0 30095 7 1 2 63844 62094
0 30096 7 1 2 66640 30095
0 30097 5 1 1 30096
0 30098 7 1 2 30093 30097
0 30099 5 1 1 30098
0 30100 7 1 2 41400 57599
0 30101 7 1 2 59905 30100
0 30102 7 1 2 30099 30101
0 30103 5 1 1 30102
0 30104 7 1 2 30082 30103
0 30105 5 1 1 30104
0 30106 7 1 2 57655 30105
0 30107 5 1 1 30106
0 30108 7 1 2 24402 55196
0 30109 5 1 1 30108
0 30110 7 1 2 54179 47559
0 30111 5 1 1 30110
0 30112 7 1 2 62004 30111
0 30113 5 1 1 30112
0 30114 7 1 2 30109 30113
0 30115 5 1 1 30114
0 30116 7 2 2 47488 54623
0 30117 7 1 2 53924 66642
0 30118 7 1 2 55803 30117
0 30119 5 1 1 30118
0 30120 7 1 2 30115 30119
0 30121 5 1 1 30120
0 30122 7 3 2 44343 41263
0 30123 7 1 2 63066 66644
0 30124 7 1 2 66564 30123
0 30125 7 1 2 30121 30124
0 30126 5 1 1 30125
0 30127 7 1 2 30107 30126
0 30128 5 1 1 30127
0 30129 7 1 2 40489 30128
0 30130 5 1 1 30129
0 30131 7 1 2 57838 65399
0 30132 5 1 1 30131
0 30133 7 1 2 52111 57065
0 30134 5 1 1 30133
0 30135 7 1 2 30132 30134
0 30136 5 1 1 30135
0 30137 7 1 2 59538 30136
0 30138 5 1 1 30137
0 30139 7 2 2 48932 65337
0 30140 5 1 1 66647
0 30141 7 1 2 57082 30140
0 30142 5 1 1 30141
0 30143 7 1 2 59710 30142
0 30144 5 1 1 30143
0 30145 7 1 2 30138 30144
0 30146 5 1 1 30145
0 30147 7 1 2 40103 30146
0 30148 5 1 1 30147
0 30149 7 1 2 59711 65869
0 30150 5 1 1 30149
0 30151 7 1 2 57741 59539
0 30152 5 1 1 30151
0 30153 7 1 2 65286 57270
0 30154 5 1 1 30153
0 30155 7 1 2 30152 30154
0 30156 5 1 1 30155
0 30157 7 1 2 40285 30156
0 30158 5 1 1 30157
0 30159 7 1 2 30150 30158
0 30160 7 1 2 30148 30159
0 30161 5 1 1 30160
0 30162 7 1 2 44344 30161
0 30163 5 1 1 30162
0 30164 7 1 2 47489 61101
0 30165 5 1 1 30164
0 30166 7 1 2 54180 50564
0 30167 5 1 1 30166
0 30168 7 1 2 30165 30167
0 30169 5 2 1 30168
0 30170 7 1 2 65228 66649
0 30171 5 1 1 30170
0 30172 7 1 2 30163 30171
0 30173 5 1 1 30172
0 30174 7 1 2 53765 30173
0 30175 5 1 1 30174
0 30176 7 1 2 52338 64477
0 30177 5 1 1 30176
0 30178 7 1 2 47535 49317
0 30179 5 1 1 30178
0 30180 7 1 2 30177 30179
0 30181 5 1 1 30180
0 30182 7 1 2 44345 50753
0 30183 7 1 2 60952 60149
0 30184 7 1 2 30182 30183
0 30185 7 1 2 61874 30184
0 30186 7 1 2 30181 30185
0 30187 5 1 1 30186
0 30188 7 1 2 41766 58932
0 30189 7 2 2 61970 30188
0 30190 7 1 2 51932 46583
0 30191 7 1 2 66651 30190
0 30192 5 1 1 30191
0 30193 7 1 2 30187 30192
0 30194 7 1 2 30175 30193
0 30195 5 1 1 30194
0 30196 7 1 2 57656 30195
0 30197 5 1 1 30196
0 30198 7 1 2 64652 64578
0 30199 7 1 2 60386 30198
0 30200 7 1 2 65918 30199
0 30201 5 1 1 30200
0 30202 7 1 2 53766 65216
0 30203 7 1 2 66650 30202
0 30204 5 1 1 30203
0 30205 7 1 2 30201 30204
0 30206 7 1 2 30197 30205
0 30207 5 1 1 30206
0 30208 7 1 2 43761 30207
0 30209 5 1 1 30208
0 30210 7 1 2 42436 63516
0 30211 5 1 1 30210
0 30212 7 1 2 53394 30211
0 30213 5 1 1 30212
0 30214 7 1 2 65322 66652
0 30215 7 1 2 30213 30214
0 30216 5 1 1 30215
0 30217 7 1 2 30209 30216
0 30218 5 1 1 30217
0 30219 7 1 2 48231 30218
0 30220 5 1 1 30219
0 30221 7 1 2 30130 30220
0 30222 5 1 1 30221
0 30223 7 1 2 45506 30222
0 30224 5 1 1 30223
0 30225 7 1 2 47567 62405
0 30226 5 2 1 30225
0 30227 7 1 2 40104 66653
0 30228 5 1 1 30227
0 30229 7 1 2 50464 30228
0 30230 5 1 1 30229
0 30231 7 1 2 43762 30230
0 30232 5 1 1 30231
0 30233 7 1 2 65473 30232
0 30234 5 2 1 30233
0 30235 7 1 2 42696 66655
0 30236 5 1 1 30235
0 30237 7 1 2 62565 52194
0 30238 5 1 1 30237
0 30239 7 1 2 30236 30238
0 30240 5 1 1 30239
0 30241 7 1 2 41401 30240
0 30242 5 1 1 30241
0 30243 7 2 2 47424 49807
0 30244 7 1 2 52189 64812
0 30245 7 1 2 66657 30244
0 30246 5 1 1 30245
0 30247 7 1 2 30242 30246
0 30248 5 1 1 30247
0 30249 7 1 2 59540 30248
0 30250 5 1 1 30249
0 30251 7 1 2 50161 51951
0 30252 5 1 1 30251
0 30253 7 1 2 49452 63494
0 30254 5 1 1 30253
0 30255 7 1 2 42174 63507
0 30256 7 1 2 30254 30255
0 30257 5 2 1 30256
0 30258 7 1 2 30252 66659
0 30259 5 1 1 30258
0 30260 7 1 2 42697 30259
0 30261 5 1 1 30260
0 30262 7 2 2 55460 51144
0 30263 5 1 1 66661
0 30264 7 1 2 61767 30263
0 30265 5 1 1 30264
0 30266 7 1 2 44545 30265
0 30267 5 1 1 30266
0 30268 7 2 2 43763 55461
0 30269 5 1 1 66663
0 30270 7 1 2 30269 52520
0 30271 5 1 1 30270
0 30272 7 1 2 44433 30271
0 30273 5 1 1 30272
0 30274 7 1 2 56707 64877
0 30275 5 2 1 30274
0 30276 7 1 2 30273 66665
0 30277 5 1 1 30276
0 30278 7 1 2 43431 30277
0 30279 5 1 1 30278
0 30280 7 1 2 30267 30279
0 30281 7 1 2 30261 30280
0 30282 5 1 1 30281
0 30283 7 1 2 59712 30282
0 30284 5 1 1 30283
0 30285 7 1 2 30250 30284
0 30286 5 1 1 30285
0 30287 7 1 2 48232 30286
0 30288 5 1 1 30287
0 30289 7 4 2 54658 57600
0 30290 7 1 2 45187 47350
0 30291 5 1 1 30290
0 30292 7 1 2 59743 61084
0 30293 7 1 2 30291 30292
0 30294 7 1 2 66667 30293
0 30295 5 1 1 30294
0 30296 7 1 2 30288 30295
0 30297 5 1 1 30296
0 30298 7 1 2 45776 30297
0 30299 5 1 1 30298
0 30300 7 1 2 59541 66656
0 30301 5 1 1 30300
0 30302 7 1 2 45507 24352
0 30303 7 1 2 3134 30302
0 30304 5 1 1 30303
0 30305 7 1 2 51084 30304
0 30306 5 1 1 30305
0 30307 7 1 2 40105 54574
0 30308 7 1 2 47168 30307
0 30309 5 2 1 30308
0 30310 7 1 2 65021 66671
0 30311 7 1 2 30306 30310
0 30312 5 1 1 30311
0 30313 7 1 2 59713 30312
0 30314 5 1 1 30313
0 30315 7 1 2 30301 30314
0 30316 5 1 1 30315
0 30317 7 1 2 44698 30316
0 30318 5 1 1 30317
0 30319 7 3 2 49890 54702
0 30320 5 1 1 66673
0 30321 7 1 2 65134 66674
0 30322 5 1 1 30321
0 30323 7 1 2 45985 30322
0 30324 7 1 2 30318 30323
0 30325 5 1 1 30324
0 30326 7 1 2 58210 59736
0 30327 5 1 1 30326
0 30328 7 1 2 59714 51595
0 30329 5 1 1 30328
0 30330 7 1 2 30327 30329
0 30331 5 1 1 30330
0 30332 7 1 2 46816 30331
0 30333 5 1 1 30332
0 30334 7 1 2 58211 65135
0 30335 5 1 1 30334
0 30336 7 1 2 30333 30335
0 30337 5 1 1 30336
0 30338 7 1 2 40106 30337
0 30339 5 1 1 30338
0 30340 7 1 2 48710 66071
0 30341 5 1 1 30340
0 30342 7 1 2 42698 30341
0 30343 7 1 2 30339 30342
0 30344 5 1 1 30343
0 30345 7 1 2 42874 30344
0 30346 7 1 2 30325 30345
0 30347 5 1 1 30346
0 30348 7 1 2 65645 59542
0 30349 7 1 2 61063 30348
0 30350 5 1 1 30349
0 30351 7 1 2 30347 30350
0 30352 5 1 1 30351
0 30353 7 1 2 54933 30352
0 30354 5 1 1 30353
0 30355 7 1 2 30299 30354
0 30356 5 1 1 30355
0 30357 7 1 2 63578 30356
0 30358 5 1 1 30357
0 30359 7 1 2 43764 66654
0 30360 5 1 1 30359
0 30361 7 1 2 64832 30360
0 30362 5 1 1 30361
0 30363 7 1 2 53767 30362
0 30364 5 1 1 30363
0 30365 7 1 2 47977 52497
0 30366 7 1 2 61455 30365
0 30367 5 1 1 30366
0 30368 7 1 2 30364 30367
0 30369 5 1 1 30368
0 30370 7 1 2 48233 30369
0 30371 5 1 1 30370
0 30372 7 1 2 60243 63134
0 30373 7 1 2 66668 30372
0 30374 5 1 1 30373
0 30375 7 1 2 30371 30374
0 30376 5 1 1 30375
0 30377 7 2 2 60104 57271
0 30378 7 1 2 30376 66676
0 30379 5 1 1 30378
0 30380 7 1 2 30358 30379
0 30381 5 1 1 30380
0 30382 7 1 2 44346 30381
0 30383 5 1 1 30382
0 30384 7 2 2 50488 57601
0 30385 7 1 2 52330 52587
0 30386 7 1 2 66678 30385
0 30387 5 1 1 30386
0 30388 7 1 2 45508 65497
0 30389 5 1 1 30388
0 30390 7 1 2 64991 30389
0 30391 7 1 2 66672 30390
0 30392 7 2 2 64884 30391
0 30393 5 1 1 66680
0 30394 7 1 2 42437 30393
0 30395 5 1 1 30394
0 30396 7 1 2 55881 30395
0 30397 5 1 1 30396
0 30398 7 1 2 44699 30397
0 30399 5 1 1 30398
0 30400 7 1 2 50596 66675
0 30401 5 1 1 30400
0 30402 7 2 2 45986 30401
0 30403 7 1 2 30399 66682
0 30404 5 1 1 30403
0 30405 7 1 2 45777 66681
0 30406 5 1 1 30405
0 30407 7 1 2 45336 62488
0 30408 5 1 1 30407
0 30409 7 1 2 65023 30408
0 30410 5 1 1 30409
0 30411 7 1 2 41402 30410
0 30412 7 1 2 30406 30411
0 30413 5 1 1 30412
0 30414 7 1 2 50205 46817
0 30415 7 1 2 48177 20894
0 30416 5 2 1 30415
0 30417 7 1 2 58231 66684
0 30418 7 1 2 30414 30417
0 30419 5 1 1 30418
0 30420 7 1 2 66165 30419
0 30421 5 1 1 30420
0 30422 7 1 2 40107 30421
0 30423 5 1 1 30422
0 30424 7 2 2 42699 65013
0 30425 7 1 2 30423 66686
0 30426 7 1 2 30413 30425
0 30427 5 1 1 30426
0 30428 7 1 2 48234 30427
0 30429 7 1 2 30404 30428
0 30430 5 1 1 30429
0 30431 7 1 2 30387 30430
0 30432 5 1 1 30431
0 30433 7 3 2 43256 65304
0 30434 7 1 2 30432 66688
0 30435 5 1 1 30434
0 30436 7 4 2 63579 46584
0 30437 7 1 2 54575 51375
0 30438 7 1 2 53768 30437
0 30439 5 1 1 30438
0 30440 7 1 2 48835 62406
0 30441 5 1 1 30440
0 30442 7 1 2 50491 64319
0 30443 7 1 2 30441 30442
0 30444 5 1 1 30443
0 30445 7 1 2 30439 30444
0 30446 5 1 1 30445
0 30447 7 1 2 48235 30446
0 30448 5 1 1 30447
0 30449 7 1 2 64107 66679
0 30450 5 1 1 30449
0 30451 7 1 2 30448 30450
0 30452 5 1 1 30451
0 30453 7 1 2 66691 30452
0 30454 5 1 1 30453
0 30455 7 3 2 47490 59328
0 30456 5 1 1 66695
0 30457 7 1 2 53769 66696
0 30458 5 1 1 30457
0 30459 7 2 2 42700 52044
0 30460 7 1 2 64847 66698
0 30461 5 1 1 30460
0 30462 7 1 2 10894 30461
0 30463 5 1 1 30462
0 30464 7 1 2 47293 30463
0 30465 5 1 1 30464
0 30466 7 1 2 30458 30465
0 30467 5 1 1 30466
0 30468 7 1 2 64488 64697
0 30469 7 1 2 30467 30468
0 30470 5 1 1 30469
0 30471 7 1 2 30454 30470
0 30472 5 1 1 30471
0 30473 7 1 2 43257 30472
0 30474 5 1 1 30473
0 30475 7 2 2 53770 63420
0 30476 7 3 2 64677 66081
0 30477 7 1 2 42875 66702
0 30478 7 1 2 64235 30477
0 30479 7 1 2 66700 30478
0 30480 5 1 1 30479
0 30481 7 1 2 30474 30480
0 30482 5 1 1 30481
0 30483 7 1 2 47812 30482
0 30484 5 1 1 30483
0 30485 7 1 2 62252 66692
0 30486 5 1 1 30485
0 30487 7 1 2 45509 60185
0 30488 7 1 2 66703 30487
0 30489 5 1 1 30488
0 30490 7 1 2 30486 30489
0 30491 5 1 1 30490
0 30492 7 1 2 53771 30491
0 30493 5 1 1 30492
0 30494 7 1 2 65008 66693
0 30495 5 1 1 30494
0 30496 7 1 2 65003 56834
0 30497 7 1 2 64698 30496
0 30498 5 1 1 30497
0 30499 7 1 2 30495 30498
0 30500 5 1 1 30499
0 30501 7 1 2 55319 30500
0 30502 5 1 1 30501
0 30503 7 1 2 30493 30502
0 30504 5 1 1 30503
0 30505 7 1 2 48236 30504
0 30506 5 1 1 30505
0 30507 7 2 2 60186 64678
0 30508 7 1 2 60775 50301
0 30509 7 1 2 66669 30508
0 30510 7 1 2 66705 30509
0 30511 5 1 1 30510
0 30512 7 1 2 30506 30511
0 30513 5 1 1 30512
0 30514 7 1 2 43258 30513
0 30515 5 1 1 30514
0 30516 7 2 2 48933 65112
0 30517 7 1 2 47127 48237
0 30518 7 1 2 57211 64679
0 30519 7 1 2 30517 30518
0 30520 7 1 2 66707 30519
0 30521 7 1 2 53772 30520
0 30522 5 1 1 30521
0 30523 7 1 2 30515 30522
0 30524 5 1 1 30523
0 30525 7 1 2 46766 30524
0 30526 5 1 1 30525
0 30527 7 1 2 30484 30526
0 30528 7 1 2 30435 30527
0 30529 7 1 2 30383 30528
0 30530 5 1 1 30529
0 30531 7 1 2 55098 30530
0 30532 5 1 1 30531
0 30533 7 1 2 42175 49819
0 30534 5 1 1 30533
0 30535 7 1 2 42438 30534
0 30536 7 1 2 65131 30535
0 30537 5 1 1 30536
0 30538 7 1 2 45778 46992
0 30539 5 1 1 30538
0 30540 7 1 2 44700 30539
0 30541 7 1 2 30537 30540
0 30542 5 1 1 30541
0 30543 7 1 2 50838 55994
0 30544 5 1 1 30543
0 30545 7 1 2 30542 30544
0 30546 5 1 1 30545
0 30547 7 1 2 45987 30546
0 30548 5 1 1 30547
0 30549 7 1 2 40108 51800
0 30550 5 1 1 30549
0 30551 7 1 2 50535 30550
0 30552 5 1 1 30551
0 30553 7 1 2 41403 30552
0 30554 5 1 1 30553
0 30555 7 1 2 57589 53168
0 30556 5 1 1 30555
0 30557 7 1 2 30554 30556
0 30558 5 1 1 30557
0 30559 7 1 2 41145 30558
0 30560 5 1 1 30559
0 30561 7 1 2 42439 59843
0 30562 7 1 2 30560 30561
0 30563 5 1 1 30562
0 30564 7 1 2 44701 46908
0 30565 5 1 1 30564
0 30566 7 1 2 42176 50050
0 30567 7 1 2 30565 30566
0 30568 5 1 1 30567
0 30569 7 1 2 46963 51765
0 30570 5 1 1 30569
0 30571 7 1 2 47813 65805
0 30572 5 1 1 30571
0 30573 7 1 2 30570 30572
0 30574 5 1 1 30573
0 30575 7 1 2 40109 30574
0 30576 5 1 1 30575
0 30577 7 1 2 50291 27487
0 30578 5 1 1 30577
0 30579 7 1 2 45779 30578
0 30580 7 1 2 30576 30579
0 30581 7 1 2 30568 30580
0 30582 5 1 1 30581
0 30583 7 1 2 42701 30582
0 30584 7 1 2 30563 30583
0 30585 5 1 1 30584
0 30586 7 1 2 30548 30585
0 30587 5 1 1 30586
0 30588 7 1 2 42876 30587
0 30589 5 1 1 30588
0 30590 7 1 2 55259 53686
0 30591 5 1 1 30590
0 30592 7 2 2 42177 55516
0 30593 7 1 2 44546 66709
0 30594 5 1 1 30593
0 30595 7 1 2 30591 30594
0 30596 5 1 1 30595
0 30597 7 1 2 43765 30596
0 30598 5 1 1 30597
0 30599 7 1 2 50292 58804
0 30600 5 1 1 30599
0 30601 7 1 2 30598 30600
0 30602 5 1 1 30601
0 30603 7 1 2 55689 30602
0 30604 5 1 1 30603
0 30605 7 1 2 47097 56011
0 30606 5 1 1 30605
0 30607 7 1 2 13173 30606
0 30608 5 1 1 30607
0 30609 7 1 2 55153 30608
0 30610 5 1 1 30609
0 30611 7 1 2 42440 56467
0 30612 5 1 1 30611
0 30613 7 1 2 30610 30612
0 30614 5 1 1 30613
0 30615 7 1 2 49301 30614
0 30616 5 1 1 30615
0 30617 7 1 2 30604 30616
0 30618 7 1 2 30589 30617
0 30619 5 1 1 30618
0 30620 7 1 2 66602 30619
0 30621 5 1 1 30620
0 30622 7 1 2 53602 51619
0 30623 5 1 1 30622
0 30624 7 1 2 46983 65764
0 30625 5 1 1 30624
0 30626 7 1 2 45337 61763
0 30627 5 1 1 30626
0 30628 7 1 2 30625 30627
0 30629 5 1 1 30628
0 30630 7 1 2 43582 30629
0 30631 5 1 1 30630
0 30632 7 1 2 30623 30631
0 30633 5 1 1 30632
0 30634 7 1 2 42178 30633
0 30635 5 1 1 30634
0 30636 7 1 2 47056 55958
0 30637 5 1 1 30636
0 30638 7 1 2 41146 30637
0 30639 5 1 1 30638
0 30640 7 1 2 30639 58459
0 30641 5 1 1 30640
0 30642 7 1 2 43766 56708
0 30643 7 1 2 30641 30642
0 30644 5 1 1 30643
0 30645 7 1 2 30635 30644
0 30646 5 1 1 30645
0 30647 7 1 2 45780 30646
0 30648 5 1 1 30647
0 30649 7 1 2 51868 46906
0 30650 5 1 1 30649
0 30651 7 1 2 66082 30650
0 30652 5 1 1 30651
0 30653 7 1 2 49386 50880
0 30654 5 1 1 30653
0 30655 7 1 2 65469 30654
0 30656 5 3 1 30655
0 30657 7 1 2 40490 66711
0 30658 5 1 1 30657
0 30659 7 1 2 30652 30658
0 30660 5 1 1 30659
0 30661 7 1 2 53773 30660
0 30662 5 1 1 30661
0 30663 7 1 2 41264 66042
0 30664 5 1 1 30663
0 30665 7 1 2 55580 59329
0 30666 5 1 1 30665
0 30667 7 1 2 30664 30666
0 30668 5 1 1 30667
0 30669 7 1 2 55462 30668
0 30670 5 1 1 30669
0 30671 7 1 2 51955 58447
0 30672 5 1 1 30671
0 30673 7 1 2 42702 60197
0 30674 7 1 2 30672 30673
0 30675 5 1 1 30674
0 30676 7 1 2 30670 30675
0 30677 5 1 1 30676
0 30678 7 1 2 42441 30677
0 30679 5 1 1 30678
0 30680 7 1 2 30662 30679
0 30681 7 1 2 30648 30680
0 30682 5 1 1 30681
0 30683 7 1 2 42877 30682
0 30684 5 1 1 30683
0 30685 7 1 2 44547 65438
0 30686 7 1 2 53854 30685
0 30687 5 1 1 30686
0 30688 7 1 2 30684 30687
0 30689 5 1 1 30688
0 30690 7 1 2 65490 30689
0 30691 5 1 1 30690
0 30692 7 1 2 30621 30691
0 30693 5 1 1 30692
0 30694 7 1 2 54984 30693
0 30695 5 1 1 30694
0 30696 7 1 2 50246 65732
0 30697 7 1 2 57303 66489
0 30698 7 1 2 30696 30697
0 30699 5 1 1 30698
0 30700 7 1 2 30695 30699
0 30701 5 1 1 30700
0 30702 7 1 2 55099 30701
0 30703 5 1 1 30702
0 30704 7 2 2 66603 64320
0 30705 5 1 1 66714
0 30706 7 2 2 46514 66527
0 30707 7 1 2 45988 66614
0 30708 7 1 2 66716 30707
0 30709 5 1 1 30708
0 30710 7 1 2 30705 30709
0 30711 5 1 1 30710
0 30712 7 1 2 47128 30711
0 30713 5 1 1 30712
0 30714 7 1 2 54257 64227
0 30715 7 1 2 66604 30714
0 30716 5 1 1 30715
0 30717 7 1 2 30713 30716
0 30718 5 1 1 30717
0 30719 7 1 2 40286 30718
0 30720 5 1 1 30719
0 30721 7 1 2 47998 66715
0 30722 5 1 1 30721
0 30723 7 1 2 30720 30722
0 30724 5 1 1 30723
0 30725 7 1 2 42442 30724
0 30726 5 1 1 30725
0 30727 7 1 2 50293 64680
0 30728 7 1 2 65113 30727
0 30729 7 1 2 63211 30728
0 30730 5 1 1 30729
0 30731 7 1 2 30726 30730
0 30732 5 1 1 30731
0 30733 7 1 2 56560 30732
0 30734 5 1 1 30733
0 30735 7 3 2 53477 61082
0 30736 7 1 2 66014 66645
0 30737 7 1 2 57304 30736
0 30738 7 1 2 66718 30737
0 30739 5 1 1 30738
0 30740 7 1 2 30734 30739
0 30741 5 1 1 30740
0 30742 7 1 2 55100 30741
0 30743 5 1 1 30742
0 30744 7 1 2 56698 66167
0 30745 5 1 1 30744
0 30746 7 1 2 56296 66699
0 30747 5 1 1 30746
0 30748 7 1 2 51933 54807
0 30749 5 2 1 30748
0 30750 7 1 2 30747 66721
0 30751 5 1 1 30750
0 30752 7 1 2 47814 30751
0 30753 5 1 1 30752
0 30754 7 1 2 52498 66163
0 30755 5 1 1 30754
0 30756 7 1 2 30753 30755
0 30757 5 1 1 30756
0 30758 7 1 2 53615 30757
0 30759 5 1 1 30758
0 30760 7 1 2 30745 30759
0 30761 5 1 1 30760
0 30762 7 1 2 66334 30761
0 30763 5 1 1 30762
0 30764 7 1 2 30743 30763
0 30765 5 1 1 30764
0 30766 7 1 2 46767 30765
0 30767 5 1 1 30766
0 30768 7 1 2 57485 63138
0 30769 7 1 2 66719 30768
0 30770 5 1 1 30769
0 30771 7 1 2 41404 66685
0 30772 5 1 1 30771
0 30773 7 1 2 40491 64920
0 30774 5 1 1 30773
0 30775 7 1 2 30772 30774
0 30776 5 1 1 30775
0 30777 7 1 2 42703 30776
0 30778 5 1 1 30777
0 30779 7 1 2 66722 30778
0 30780 5 1 1 30779
0 30781 7 1 2 62144 48592
0 30782 7 1 2 30780 30781
0 30783 5 1 1 30782
0 30784 7 1 2 30770 30783
0 30785 5 1 1 30784
0 30786 7 1 2 46585 30785
0 30787 5 1 1 30786
0 30788 7 2 2 42443 57472
0 30789 5 1 1 66723
0 30790 7 1 2 65211 30789
0 30791 5 1 1 30790
0 30792 7 1 2 51856 30791
0 30793 5 1 1 30792
0 30794 7 1 2 63655 65937
0 30795 5 1 1 30794
0 30796 7 1 2 30793 30795
0 30797 5 1 1 30796
0 30798 7 1 2 40492 30797
0 30799 5 1 1 30798
0 30800 7 1 2 53774 62903
0 30801 5 1 1 30800
0 30802 7 1 2 30799 30801
0 30803 5 1 1 30802
0 30804 7 1 2 40110 65311
0 30805 7 1 2 30803 30804
0 30806 5 1 1 30805
0 30807 7 1 2 30787 30806
0 30808 5 1 1 30807
0 30809 7 1 2 43259 30808
0 30810 5 1 1 30809
0 30811 7 1 2 40287 55553
0 30812 5 1 1 30811
0 30813 7 1 2 52476 30812
0 30814 5 1 1 30813
0 30815 7 1 2 55101 66704
0 30816 7 1 2 63009 30815
0 30817 7 1 2 30814 30816
0 30818 5 1 1 30817
0 30819 7 1 2 30810 30818
0 30820 5 1 1 30819
0 30821 7 1 2 46861 30820
0 30822 5 1 1 30821
0 30823 7 2 2 64885 64895
0 30824 7 1 2 577 54576
0 30825 7 1 2 52726 30824
0 30826 5 1 1 30825
0 30827 7 1 2 48383 50162
0 30828 5 1 1 30827
0 30829 7 1 2 30826 30828
0 30830 7 1 2 66725 30829
0 30831 5 2 1 30830
0 30832 7 1 2 42444 66727
0 30833 5 1 1 30832
0 30834 7 1 2 55882 30833
0 30835 5 1 1 30834
0 30836 7 1 2 44702 30835
0 30837 5 1 1 30836
0 30838 7 1 2 66683 30837
0 30839 5 1 1 30838
0 30840 7 1 2 45781 66728
0 30841 5 1 1 30840
0 30842 7 1 2 50189 46914
0 30843 5 1 1 30842
0 30844 7 1 2 62349 30843
0 30845 5 1 1 30844
0 30846 7 1 2 30841 30845
0 30847 5 1 1 30846
0 30848 7 1 2 41405 30847
0 30849 5 1 1 30848
0 30850 7 1 2 40493 64913
0 30851 5 1 1 30850
0 30852 7 1 2 53562 64284
0 30853 5 1 1 30852
0 30854 7 1 2 30851 30853
0 30855 5 1 1 30854
0 30856 7 1 2 40288 30855
0 30857 5 1 1 30856
0 30858 7 1 2 65388 66143
0 30859 5 1 1 30858
0 30860 7 1 2 30857 30859
0 30861 5 1 1 30860
0 30862 7 1 2 40111 30861
0 30863 5 1 1 30862
0 30864 7 1 2 66687 30863
0 30865 7 1 2 30849 30864
0 30866 5 1 1 30865
0 30867 7 1 2 53616 30866
0 30868 7 1 2 30839 30867
0 30869 5 1 1 30868
0 30870 7 1 2 41265 66017
0 30871 7 1 2 64108 30870
0 30872 5 1 1 30871
0 30873 7 1 2 30869 30872
0 30874 5 1 1 30873
0 30875 7 1 2 66335 30874
0 30876 5 1 1 30875
0 30877 7 1 2 53775 65454
0 30878 5 1 1 30877
0 30879 7 1 2 50700 64073
0 30880 7 1 2 52678 30879
0 30881 5 1 1 30880
0 30882 7 1 2 30878 30881
0 30883 5 1 1 30882
0 30884 7 1 2 42878 30883
0 30885 5 1 1 30884
0 30886 7 1 2 61188 63172
0 30887 5 1 1 30886
0 30888 7 1 2 30885 30887
0 30889 5 1 1 30888
0 30890 7 1 2 64865 65491
0 30891 7 1 2 30889 30890
0 30892 5 1 1 30891
0 30893 7 1 2 30876 30892
0 30894 7 1 2 30822 30893
0 30895 7 1 2 30767 30894
0 30896 7 1 2 30703 30895
0 30897 5 1 1 30896
0 30898 7 1 2 49052 30897
0 30899 5 1 1 30898
0 30900 7 1 2 25758 65887
0 30901 5 1 1 30900
0 30902 7 1 2 47294 30901
0 30903 5 1 1 30902
0 30904 7 1 2 52515 57066
0 30905 5 1 1 30904
0 30906 7 1 2 30903 30905
0 30907 5 1 1 30906
0 30908 7 1 2 55320 30907
0 30909 5 1 1 30908
0 30910 7 1 2 55859 60203
0 30911 5 1 1 30910
0 30912 7 1 2 30909 30911
0 30913 5 1 1 30912
0 30914 7 1 2 42445 30913
0 30915 5 1 1 30914
0 30916 7 1 2 45338 57083
0 30917 5 1 1 30916
0 30918 7 1 2 57748 30917
0 30919 5 2 1 30918
0 30920 7 1 2 57845 66729
0 30921 5 1 1 30920
0 30922 7 1 2 53756 11410
0 30923 5 1 1 30922
0 30924 7 1 2 42179 30923
0 30925 7 1 2 30921 30924
0 30926 5 1 1 30925
0 30927 7 1 2 64508 60947
0 30928 5 1 1 30927
0 30929 7 2 2 46432 53776
0 30930 7 1 2 65530 66731
0 30931 5 1 1 30930
0 30932 7 1 2 30928 30931
0 30933 5 1 1 30932
0 30934 7 1 2 47491 30933
0 30935 5 1 1 30934
0 30936 7 1 2 56054 59430
0 30937 7 1 2 66011 30936
0 30938 5 1 1 30937
0 30939 7 1 2 30935 30938
0 30940 7 1 2 30926 30939
0 30941 7 1 2 30915 30940
0 30942 5 1 1 30941
0 30943 7 1 2 48238 30942
0 30944 5 1 1 30943
0 30945 7 1 2 64102 64790
0 30946 7 1 2 60244 58646
0 30947 7 1 2 30945 30946
0 30948 5 1 1 30947
0 30949 7 1 2 30944 30948
0 30950 5 1 1 30949
0 30951 7 1 2 66336 30950
0 30952 5 1 1 30951
0 30953 7 1 2 57578 56628
0 30954 7 1 2 64566 52886
0 30955 7 1 2 30953 30954
0 30956 7 1 2 65806 30955
0 30957 5 1 1 30956
0 30958 7 1 2 62710 65994
0 30959 7 1 2 51264 30958
0 30960 7 1 2 53777 30959
0 30961 5 1 1 30960
0 30962 7 1 2 30957 30961
0 30963 5 1 1 30962
0 30964 7 1 2 48239 65104
0 30965 7 1 2 30963 30964
0 30966 5 1 1 30965
0 30967 7 1 2 30952 30966
0 30968 5 1 1 30967
0 30969 7 1 2 47815 30968
0 30970 5 1 1 30969
0 30971 7 1 2 28178 66660
0 30972 5 1 1 30971
0 30973 7 1 2 42704 30972
0 30974 5 1 1 30973
0 30975 7 1 2 44434 55463
0 30976 7 1 2 49891 30975
0 30977 5 1 1 30976
0 30978 7 1 2 66666 30977
0 30979 5 1 1 30978
0 30980 7 1 2 43432 30979
0 30981 5 1 1 30980
0 30982 7 1 2 45782 30981
0 30983 7 1 2 30974 30982
0 30984 5 1 1 30983
0 30985 7 1 2 65025 63508
0 30986 5 1 1 30985
0 30987 7 1 2 42446 30986
0 30988 7 1 2 63493 64154
0 30989 5 1 1 30988
0 30990 7 1 2 55464 65018
0 30991 5 1 1 30990
0 30992 7 1 2 30989 30991
0 30993 7 1 2 30987 30992
0 30994 5 1 1 30993
0 30995 7 1 2 57067 30994
0 30996 7 1 2 30984 30995
0 30997 5 1 1 30996
0 30998 7 1 2 48934 65123
0 30999 7 1 2 66732 30998
0 31000 5 1 1 30999
0 31001 7 1 2 30997 31000
0 31002 5 1 1 31001
0 31003 7 1 2 66337 31002
0 31004 5 1 1 31003
0 31005 7 1 2 65373 59170
0 31006 5 1 1 31005
0 31007 7 1 2 53603 52588
0 31008 5 1 1 31007
0 31009 7 1 2 31006 31008
0 31010 5 1 1 31009
0 31011 7 1 2 45783 31010
0 31012 5 1 1 31011
0 31013 7 1 2 64878 60560
0 31014 5 1 1 31013
0 31015 7 1 2 31012 31014
0 31016 5 1 1 31015
0 31017 7 1 2 43433 31016
0 31018 5 1 1 31017
0 31019 7 1 2 52012 55468
0 31020 7 1 2 58696 31019
0 31021 5 1 1 31020
0 31022 7 1 2 31018 31021
0 31023 5 1 1 31022
0 31024 7 1 2 53999 31023
0 31025 5 1 1 31024
0 31026 7 1 2 41147 48618
0 31027 7 1 2 60561 31026
0 31028 5 1 1 31027
0 31029 7 3 2 52462 65161
0 31030 5 1 1 66733
0 31031 7 1 2 48378 53747
0 31032 5 1 1 31031
0 31033 7 1 2 31030 31032
0 31034 5 1 1 31033
0 31035 7 1 2 40112 47190
0 31036 7 1 2 31034 31035
0 31037 5 1 1 31036
0 31038 7 1 2 31028 31037
0 31039 5 1 1 31038
0 31040 7 1 2 41983 31039
0 31041 5 1 1 31040
0 31042 7 3 2 47492 52422
0 31043 7 1 2 66736 66734
0 31044 5 1 1 31043
0 31045 7 1 2 56548 66662
0 31046 5 1 1 31045
0 31047 7 1 2 31044 31046
0 31048 5 1 1 31047
0 31049 7 1 2 45339 31048
0 31050 5 1 1 31049
0 31051 7 2 2 40289 49718
0 31052 5 1 1 66739
0 31053 7 1 2 66735 66740
0 31054 5 1 1 31053
0 31055 7 1 2 31050 31054
0 31056 7 1 2 31041 31055
0 31057 5 1 1 31056
0 31058 7 1 2 40494 31057
0 31059 5 1 1 31058
0 31060 7 1 2 47493 53387
0 31061 5 1 1 31060
0 31062 7 1 2 55560 31061
0 31063 5 1 1 31062
0 31064 7 1 2 52331 65117
0 31065 7 1 2 31063 31064
0 31066 5 1 1 31065
0 31067 7 1 2 31059 31066
0 31068 5 1 1 31067
0 31069 7 1 2 54181 31068
0 31070 5 1 1 31069
0 31071 7 1 2 31025 31070
0 31072 5 1 1 31071
0 31073 7 1 2 42180 31072
0 31074 5 1 1 31073
0 31075 7 1 2 50206 53778
0 31076 7 2 2 50849 54000
0 31077 7 1 2 66741 51154
0 31078 7 1 2 31075 31077
0 31079 5 1 1 31078
0 31080 7 2 2 44435 65446
0 31081 7 4 2 47816 47662
0 31082 7 1 2 66743 66745
0 31083 5 1 1 31082
0 31084 7 1 2 63033 65114
0 31085 5 1 1 31084
0 31086 7 1 2 31083 31085
0 31087 5 1 1 31086
0 31088 7 1 2 44218 55216
0 31089 7 1 2 61647 31088
0 31090 7 1 2 31087 31089
0 31091 5 1 1 31090
0 31092 7 1 2 31079 31091
0 31093 7 1 2 31074 31092
0 31094 5 1 1 31093
0 31095 7 1 2 65105 31094
0 31096 5 1 1 31095
0 31097 7 1 2 31004 31096
0 31098 5 1 1 31097
0 31099 7 1 2 42879 31098
0 31100 5 1 1 31099
0 31101 7 1 2 61544 50701
0 31102 7 2 2 64427 64681
0 31103 7 1 2 61714 66749
0 31104 7 1 2 31101 31103
0 31105 7 1 2 50991 31104
0 31106 5 1 1 31105
0 31107 7 1 2 31100 31106
0 31108 5 1 1 31107
0 31109 7 1 2 46296 31108
0 31110 5 1 1 31109
0 31111 7 1 2 30970 31110
0 31112 7 1 2 30899 31111
0 31113 7 1 2 30532 31112
0 31114 7 1 2 30224 31113
0 31115 5 1 1 31114
0 31116 7 1 2 31115 57548
0 31117 5 1 1 31116
0 31118 7 1 2 58186 59817
0 31119 5 1 1 31118
0 31120 7 1 2 31119 22061
0 31121 5 1 1 31120
0 31122 7 1 2 40968 31121
0 31123 5 1 1 31122
0 31124 7 1 2 44436 54586
0 31125 7 1 2 56161 31124
0 31126 5 1 1 31125
0 31127 7 1 2 31123 31126
0 31128 5 1 1 31127
0 31129 7 1 2 44129 31128
0 31130 5 1 1 31129
0 31131 7 1 2 48441 61023
0 31132 5 1 1 31131
0 31133 7 1 2 31130 31132
0 31134 5 1 1 31133
0 31135 7 1 2 43434 31134
0 31136 5 1 1 31135
0 31137 7 1 2 44437 58428
0 31138 5 1 1 31137
0 31139 7 1 2 19897 31138
0 31140 5 1 1 31139
0 31141 7 1 2 57068 31140
0 31142 5 1 1 31141
0 31143 7 1 2 31136 31142
0 31144 5 1 1 31143
0 31145 7 1 2 49605 31144
0 31146 5 1 1 31145
0 31147 7 1 2 56414 51552
0 31148 5 1 1 31147
0 31149 7 1 2 483 31148
0 31150 5 1 1 31149
0 31151 7 1 2 64515 31150
0 31152 5 1 1 31151
0 31153 7 1 2 31146 31152
0 31154 5 1 1 31153
0 31155 7 1 2 65206 31154
0 31156 5 1 1 31155
0 31157 7 1 2 40879 58781
0 31158 5 1 1 31157
0 31159 7 1 2 59833 31158
0 31160 5 1 1 31159
0 31161 7 1 2 48521 31160
0 31162 5 1 1 31161
0 31163 7 1 2 40880 65656
0 31164 5 1 1 31163
0 31165 7 1 2 31162 31164
0 31166 5 1 1 31165
0 31167 7 1 2 62677 56273
0 31168 5 1 1 31167
0 31169 7 1 2 44967 58941
0 31170 7 1 2 59818 31169
0 31171 5 2 1 31170
0 31172 7 1 2 31168 66751
0 31173 5 1 1 31172
0 31174 7 1 2 31166 31173
0 31175 5 1 1 31174
0 31176 7 1 2 56080 51731
0 31177 7 1 2 54001 31176
0 31178 7 1 2 54524 31177
0 31179 5 1 1 31178
0 31180 7 1 2 31175 31179
0 31181 7 1 2 31156 31180
0 31182 5 1 1 31181
0 31183 7 1 2 41984 31182
0 31184 5 1 1 31183
0 31185 7 1 2 47922 57533
0 31186 5 1 1 31185
0 31187 7 1 2 47425 61648
0 31188 7 1 2 57152 31187
0 31189 5 1 1 31188
0 31190 7 1 2 31186 31189
0 31191 5 1 1 31190
0 31192 7 1 2 53465 31191
0 31193 5 1 1 31192
0 31194 7 1 2 46721 60751
0 31195 7 1 2 58782 31194
0 31196 7 1 2 57130 31195
0 31197 5 1 1 31196
0 31198 7 1 2 31193 31197
0 31199 5 1 1 31198
0 31200 7 1 2 52932 31199
0 31201 5 1 1 31200
0 31202 7 1 2 58429 61172
0 31203 5 1 1 31202
0 31204 7 1 2 53466 53534
0 31205 7 1 2 56463 31204
0 31206 5 1 1 31205
0 31207 7 1 2 31203 31206
0 31208 5 1 1 31207
0 31209 7 1 2 60782 31208
0 31210 5 1 1 31209
0 31211 7 1 2 31201 31210
0 31212 7 1 2 31184 31211
0 31213 5 1 1 31212
0 31214 7 1 2 43583 31213
0 31215 5 1 1 31214
0 31216 7 3 2 55828 56095
0 31217 7 2 2 57717 66753
0 31218 5 1 1 66756
0 31219 7 1 2 60589 60783
0 31220 7 1 2 66757 31219
0 31221 5 1 1 31220
0 31222 7 1 2 31215 31221
0 31223 5 1 1 31222
0 31224 7 1 2 65323 31223
0 31225 5 1 1 31224
0 31226 7 1 2 46297 31225
0 31227 5 1 1 31226
0 31228 7 1 2 52209 57976
0 31229 7 1 2 58942 31228
0 31230 5 1 1 31229
0 31231 7 3 2 49606 55517
0 31232 5 2 1 66758
0 31233 7 1 2 56533 55804
0 31234 5 1 1 31233
0 31235 7 1 2 66761 31234
0 31236 5 1 1 31235
0 31237 7 1 2 47351 49053
0 31238 7 1 2 31236 31237
0 31239 5 1 1 31238
0 31240 7 1 2 31230 31239
0 31241 5 1 1 31240
0 31242 7 1 2 41985 31241
0 31243 5 1 1 31242
0 31244 7 2 2 49054 63510
0 31245 7 1 2 55518 66763
0 31246 5 1 1 31245
0 31247 7 1 2 31243 31246
0 31248 5 1 1 31247
0 31249 7 1 2 49217 31248
0 31250 5 1 1 31249
0 31251 7 1 2 66764 56473
0 31252 5 1 1 31251
0 31253 7 1 2 48935 56262
0 31254 7 1 2 57711 31253
0 31255 5 1 1 31254
0 31256 7 1 2 31252 31255
0 31257 5 1 1 31256
0 31258 7 1 2 57977 31257
0 31259 5 1 1 31258
0 31260 7 1 2 55519 66517
0 31261 5 1 1 31260
0 31262 7 1 2 56096 51978
0 31263 7 1 2 56537 31262
0 31264 5 2 1 31263
0 31265 7 1 2 31261 66765
0 31266 5 1 1 31265
0 31267 7 1 2 49055 31266
0 31268 5 1 1 31267
0 31269 7 2 2 48522 55520
0 31270 5 1 1 66767
0 31271 7 1 2 56747 66768
0 31272 5 1 1 31271
0 31273 7 2 2 54535 53049
0 31274 7 2 2 59081 49282
0 31275 7 1 2 66769 66771
0 31276 5 1 1 31275
0 31277 7 1 2 31272 31276
0 31278 7 1 2 31268 31277
0 31279 5 1 1 31278
0 31280 7 1 2 47923 31279
0 31281 5 1 1 31280
0 31282 7 1 2 31259 31281
0 31283 7 1 2 31250 31282
0 31284 5 1 1 31283
0 31285 7 3 2 43584 46433
0 31286 7 1 2 65324 66773
0 31287 7 1 2 31284 31286
0 31288 5 1 1 31287
0 31289 7 2 2 53467 55302
0 31290 7 1 2 64699 63755
0 31291 5 1 1 31290
0 31292 7 1 2 46586 63698
0 31293 7 1 2 59225 31292
0 31294 5 1 1 31293
0 31295 7 1 2 31291 31294
0 31296 5 1 1 31295
0 31297 7 1 2 66776 31296
0 31298 5 1 1 31297
0 31299 7 1 2 64730 66754
0 31300 5 1 1 31299
0 31301 7 1 2 63680 57978
0 31302 5 1 1 31301
0 31303 7 1 2 31300 31302
0 31304 5 1 1 31303
0 31305 7 1 2 46587 31304
0 31306 5 1 1 31305
0 31307 7 2 2 65434 57979
0 31308 7 2 2 64656 66778
0 31309 7 1 2 59609 66780
0 31310 5 1 1 31309
0 31311 7 2 2 44130 59006
0 31312 7 2 2 59314 66782
0 31313 7 2 2 41849 58663
0 31314 7 1 2 66786 66755
0 31315 7 1 2 66784 31314
0 31316 5 1 1 31315
0 31317 7 1 2 31310 31316
0 31318 7 1 2 31306 31317
0 31319 5 1 1 31318
0 31320 7 1 2 49607 31319
0 31321 5 1 1 31320
0 31322 7 1 2 31298 31321
0 31323 5 1 1 31322
0 31324 7 1 2 43140 52286
0 31325 7 1 2 31323 31324
0 31326 5 1 1 31325
0 31327 7 1 2 43027 31326
0 31328 7 1 2 31288 31327
0 31329 5 1 1 31328
0 31330 7 1 2 43260 31329
0 31331 7 1 2 31227 31330
0 31332 5 1 1 31331
0 31333 7 3 2 59510 58837
0 31334 7 3 2 43141 66788
0 31335 7 1 2 62455 63709
0 31336 7 3 2 45188 64657
0 31337 7 1 2 66794 58653
0 31338 7 1 2 31335 31337
0 31339 7 1 2 66791 31338
0 31340 5 1 1 31339
0 31341 7 1 2 51629 52199
0 31342 7 1 2 65769 31341
0 31343 7 3 2 57147 59065
0 31344 7 1 2 46588 66797
0 31345 7 1 2 31342 31344
0 31346 7 1 2 63832 31345
0 31347 5 1 1 31346
0 31348 7 1 2 31340 31347
0 31349 5 1 1 31348
0 31350 7 1 2 44438 49790
0 31351 7 1 2 31349 31350
0 31352 5 1 1 31351
0 31353 7 1 2 31332 31352
0 31354 5 1 1 31353
0 31355 7 1 2 43767 31354
0 31356 5 1 1 31355
0 31357 7 1 2 59261 59715
0 31358 7 1 2 63200 31357
0 31359 5 1 1 31358
0 31360 7 2 2 48345 63538
0 31361 7 1 2 66015 48361
0 31362 7 1 2 66800 31361
0 31363 5 1 1 31362
0 31364 7 1 2 31359 31363
0 31365 5 1 1 31364
0 31366 7 1 2 43768 31365
0 31367 5 1 1 31366
0 31368 7 1 2 65896 50136
0 31369 7 1 2 66801 31368
0 31370 5 1 1 31369
0 31371 7 1 2 31367 31370
0 31372 5 1 1 31371
0 31373 7 1 2 42705 31372
0 31374 5 1 1 31373
0 31375 7 1 2 66513 48362
0 31376 7 1 2 64875 31375
0 31377 5 1 1 31376
0 31378 7 1 2 31374 31377
0 31379 5 1 1 31378
0 31380 7 1 2 40881 31379
0 31381 5 1 1 31380
0 31382 7 1 2 41986 59196
0 31383 5 1 1 31382
0 31384 7 1 2 60495 31383
0 31385 5 1 1 31384
0 31386 7 1 2 46693 31385
0 31387 5 1 1 31386
0 31388 7 1 2 47878 64080
0 31389 5 1 1 31388
0 31390 7 1 2 31387 31389
0 31391 5 1 1 31390
0 31392 7 1 2 63076 66774
0 31393 7 1 2 59377 31392
0 31394 7 1 2 31391 31393
0 31395 5 1 1 31394
0 31396 7 1 2 31381 31395
0 31397 5 1 1 31396
0 31398 7 1 2 44439 31397
0 31399 5 1 1 31398
0 31400 7 1 2 40882 63201
0 31401 5 3 1 31400
0 31402 7 1 2 7754 66802
0 31403 5 5 1 31402
0 31404 7 1 2 59192 66805
0 31405 5 1 1 31404
0 31406 7 1 2 42447 64335
0 31407 7 1 2 60062 31406
0 31408 5 1 1 31407
0 31409 7 1 2 31405 31408
0 31410 5 1 1 31409
0 31411 7 1 2 55141 31410
0 31412 5 1 1 31411
0 31413 7 1 2 55834 50767
0 31414 7 1 2 57812 31413
0 31415 5 2 1 31414
0 31416 7 1 2 31412 66810
0 31417 5 1 1 31416
0 31418 7 1 2 59716 31417
0 31419 5 1 1 31418
0 31420 7 1 2 31399 31419
0 31421 5 1 1 31420
0 31422 7 1 2 44347 31421
0 31423 5 1 1 31422
0 31424 7 1 2 47879 66806
0 31425 5 1 1 31424
0 31426 7 1 2 53656 48346
0 31427 7 1 2 64336 31426
0 31428 5 2 1 31427
0 31429 7 1 2 31425 66812
0 31430 5 1 1 31429
0 31431 7 2 2 46850 31430
0 31432 5 1 1 66814
0 31433 7 1 2 48318 58969
0 31434 7 1 2 64293 31433
0 31435 5 1 1 31434
0 31436 7 1 2 31432 31435
0 31437 5 1 1 31436
0 31438 7 1 2 42706 31437
0 31439 5 1 1 31438
0 31440 7 1 2 66263 47868
0 31441 5 1 1 31440
0 31442 7 1 2 66803 31441
0 31443 5 1 1 31442
0 31444 7 1 2 50335 66664
0 31445 7 1 2 31443 31444
0 31446 5 1 1 31445
0 31447 7 1 2 31439 31446
0 31448 5 1 1 31447
0 31449 7 1 2 43585 31448
0 31450 5 1 1 31449
0 31451 7 1 2 66811 31450
0 31452 5 1 1 31451
0 31453 7 1 2 65229 31452
0 31454 5 1 1 31453
0 31455 7 1 2 31423 31454
0 31456 5 1 1 31455
0 31457 7 1 2 43435 31456
0 31458 5 1 1 31457
0 31459 7 1 2 44703 58830
0 31460 5 1 1 31459
0 31461 7 2 2 44440 47853
0 31462 7 1 2 49218 66816
0 31463 7 1 2 55540 31462
0 31464 5 1 1 31463
0 31465 7 1 2 31460 31464
0 31466 5 1 1 31465
0 31467 7 1 2 43586 31466
0 31468 5 1 1 31467
0 31469 7 1 2 42707 19745
0 31470 7 1 2 50683 53694
0 31471 5 2 1 31470
0 31472 7 1 2 58355 66818
0 31473 7 1 2 31469 31472
0 31474 5 1 1 31473
0 31475 7 1 2 31468 31474
0 31476 5 1 1 31475
0 31477 7 1 2 43769 31476
0 31478 5 1 1 31477
0 31479 7 1 2 52262 56012
0 31480 7 1 2 64337 31479
0 31481 5 1 1 31480
0 31482 7 1 2 31478 31481
0 31483 5 1 1 31482
0 31484 7 1 2 53657 31483
0 31485 5 1 1 31484
0 31486 7 1 2 48379 57486
0 31487 7 1 2 60054 31486
0 31488 7 1 2 59193 31487
0 31489 5 1 1 31488
0 31490 7 1 2 31485 31489
0 31491 5 1 1 31490
0 31492 7 1 2 66605 31491
0 31493 5 1 1 31492
0 31494 7 1 2 31458 31493
0 31495 5 1 1 31494
0 31496 7 1 2 57657 31495
0 31497 5 1 1 31496
0 31498 7 2 2 55142 61216
0 31499 7 1 2 47352 66807
0 31500 5 1 1 31499
0 31501 7 1 2 66264 58953
0 31502 5 1 1 31501
0 31503 7 1 2 31500 31502
0 31504 5 1 1 31503
0 31505 7 1 2 66820 31504
0 31506 5 1 1 31505
0 31507 7 1 2 49337 51305
0 31508 5 1 1 31507
0 31509 7 1 2 547 31508
0 31510 5 1 1 31509
0 31511 7 1 2 53658 31510
0 31512 5 1 1 31511
0 31513 7 1 2 57487 59355
0 31514 5 1 1 31513
0 31515 7 1 2 31512 31514
0 31516 5 1 1 31515
0 31517 7 1 2 45784 31516
0 31518 5 1 1 31517
0 31519 7 1 2 66813 31518
0 31520 5 1 1 31519
0 31521 7 1 2 46722 31520
0 31522 5 1 1 31521
0 31523 7 1 2 43436 66815
0 31524 5 1 1 31523
0 31525 7 1 2 31522 31524
0 31526 5 1 1 31525
0 31527 7 1 2 43587 31526
0 31528 5 1 1 31527
0 31529 7 1 2 64294 61070
0 31530 5 1 1 31529
0 31531 7 1 2 43437 53687
0 31532 5 1 1 31531
0 31533 7 1 2 50684 31532
0 31534 5 2 1 31533
0 31535 7 2 2 46165 53659
0 31536 7 1 2 43770 66824
0 31537 7 1 2 66822 31536
0 31538 5 1 1 31537
0 31539 7 1 2 31530 31538
0 31540 5 1 1 31539
0 31541 7 1 2 51553 31540
0 31542 5 1 1 31541
0 31543 7 1 2 31528 31542
0 31544 5 1 1 31543
0 31545 7 1 2 42708 31544
0 31546 5 1 1 31545
0 31547 7 1 2 31506 31546
0 31548 5 1 1 31547
0 31549 7 1 2 65217 31548
0 31550 5 1 1 31549
0 31551 7 1 2 31497 31550
0 31552 5 1 1 31551
0 31553 7 1 2 49056 31552
0 31554 5 1 1 31553
0 31555 7 1 2 56333 59717
0 31556 7 1 2 56039 61191
0 31557 7 1 2 31555 31556
0 31558 5 1 1 31557
0 31559 7 1 2 56153 61964
0 31560 5 1 1 31559
0 31561 7 1 2 44131 55829
0 31562 7 1 2 54934 31561
0 31563 5 1 1 31562
0 31564 7 1 2 31560 31563
0 31565 5 1 1 31564
0 31566 7 1 2 46515 65897
0 31567 7 1 2 31565 31566
0 31568 5 1 1 31567
0 31569 7 1 2 31558 31568
0 31570 5 1 1 31569
0 31571 7 1 2 44441 31570
0 31572 5 1 1 31571
0 31573 7 2 2 49808 48327
0 31574 7 1 2 59378 66826
0 31575 7 1 2 66050 31574
0 31576 5 1 1 31575
0 31577 7 1 2 31572 31576
0 31578 5 1 1 31577
0 31579 7 1 2 44348 31578
0 31580 5 1 1 31579
0 31581 7 2 2 41987 55541
0 31582 5 1 1 66828
0 31583 7 1 2 44442 52463
0 31584 5 1 1 31583
0 31585 7 1 2 31582 31584
0 31586 5 1 1 31585
0 31587 7 2 2 44132 49809
0 31588 7 2 2 46298 66830
0 31589 7 1 2 65230 66832
0 31590 7 1 2 31586 31589
0 31591 5 1 1 31590
0 31592 7 1 2 31580 31591
0 31593 5 2 1 31592
0 31594 7 1 2 54002 66834
0 31595 5 1 1 31594
0 31596 7 2 2 44443 49810
0 31597 7 2 2 66836 66829
0 31598 5 1 1 66838
0 31599 7 1 2 40495 58783
0 31600 5 1 1 31599
0 31601 7 1 2 31598 31600
0 31602 5 2 1 31601
0 31603 7 3 2 44133 62766
0 31604 7 2 2 46589 66842
0 31605 7 1 2 54099 66845
0 31606 7 1 2 66840 31605
0 31607 5 1 1 31606
0 31608 7 1 2 31595 31607
0 31609 5 1 1 31608
0 31610 7 1 2 43438 31609
0 31611 5 1 1 31610
0 31612 7 1 2 43142 52405
0 31613 7 1 2 48836 55469
0 31614 7 1 2 31612 31613
0 31615 5 1 1 31614
0 31616 7 1 2 26625 31615
0 31617 5 1 1 31616
0 31618 7 1 2 49811 62505
0 31619 7 1 2 31617 31618
0 31620 5 1 1 31619
0 31621 7 3 2 40496 52406
0 31622 5 1 1 66847
0 31623 7 1 2 56629 66848
0 31624 7 1 2 61204 31623
0 31625 5 1 1 31624
0 31626 7 1 2 31620 31625
0 31627 5 1 1 31626
0 31628 7 1 2 66846 31627
0 31629 5 1 1 31628
0 31630 7 1 2 31611 31629
0 31631 5 1 1 31630
0 31632 7 1 2 57658 31631
0 31633 5 1 1 31632
0 31634 7 1 2 66821 62688
0 31635 5 1 1 31634
0 31636 7 1 2 49765 60414
0 31637 5 1 1 31636
0 31638 7 2 2 40497 52423
0 31639 7 1 2 48837 66850
0 31640 5 1 1 31639
0 31641 7 1 2 31637 31640
0 31642 5 1 1 31641
0 31643 7 1 2 54100 31642
0 31644 5 1 1 31643
0 31645 7 3 2 53925 49812
0 31646 7 1 2 56820 66852
0 31647 7 1 2 49960 31646
0 31648 5 1 1 31647
0 31649 7 1 2 31644 31648
0 31650 5 1 1 31649
0 31651 7 1 2 42709 31650
0 31652 5 1 1 31651
0 31653 7 1 2 31635 31652
0 31654 5 1 1 31653
0 31655 7 1 2 60404 56354
0 31656 7 1 2 66795 31655
0 31657 7 1 2 31654 31656
0 31658 5 1 1 31657
0 31659 7 1 2 31633 31658
0 31660 5 1 1 31659
0 31661 7 1 2 52933 31660
0 31662 5 1 1 31661
0 31663 7 2 2 52215 54475
0 31664 5 1 1 66855
0 31665 7 1 2 48936 66856
0 31666 7 1 2 66641 31665
0 31667 5 1 1 31666
0 31668 7 2 2 59977 66051
0 31669 7 2 2 49813 66857
0 31670 7 1 2 65287 66859
0 31671 5 1 1 31670
0 31672 7 2 2 47978 61715
0 31673 7 1 2 60105 66219
0 31674 7 1 2 66861 31673
0 31675 5 1 1 31674
0 31676 7 1 2 31671 31675
0 31677 5 1 1 31676
0 31678 7 1 2 40883 31677
0 31679 5 1 1 31678
0 31680 7 1 2 46516 57687
0 31681 7 2 2 55777 31680
0 31682 7 1 2 64791 66092
0 31683 7 1 2 66863 31682
0 31684 5 1 1 31683
0 31685 7 1 2 31679 31684
0 31686 5 1 1 31685
0 31687 7 1 2 44349 31686
0 31688 5 1 1 31687
0 31689 7 1 2 49119 66460
0 31690 7 1 2 66860 31689
0 31691 5 1 1 31690
0 31692 7 1 2 31688 31691
0 31693 5 1 1 31692
0 31694 7 1 2 47426 31693
0 31695 5 1 1 31694
0 31696 7 1 2 31667 31695
0 31697 5 1 1 31696
0 31698 7 1 2 57659 52424
0 31699 7 1 2 31697 31698
0 31700 5 1 1 31699
0 31701 7 1 2 51310 66839
0 31702 5 1 1 31701
0 31703 7 1 2 31664 31702
0 31704 5 1 1 31703
0 31705 7 1 2 64682 59665
0 31706 7 1 2 61581 31705
0 31707 7 1 2 31704 31706
0 31708 5 1 1 31707
0 31709 7 1 2 31700 31708
0 31710 5 1 1 31709
0 31711 7 1 2 48278 31710
0 31712 5 1 1 31711
0 31713 7 1 2 65464 50540
0 31714 5 1 1 31713
0 31715 7 1 2 55985 62952
0 31716 5 1 1 31715
0 31717 7 1 2 31714 31716
0 31718 5 1 1 31717
0 31719 7 1 2 52425 31718
0 31720 5 1 1 31719
0 31721 7 1 2 51153 9443
0 31722 5 1 1 31721
0 31723 7 1 2 50676 31722
0 31724 5 1 1 31723
0 31725 7 1 2 59405 51155
0 31726 5 1 1 31725
0 31727 7 1 2 31724 31726
0 31728 5 1 1 31727
0 31729 7 1 2 42710 48192
0 31730 7 1 2 31728 31729
0 31731 5 1 1 31730
0 31732 7 1 2 31720 31731
0 31733 5 2 1 31732
0 31734 7 1 2 66865 62602
0 31735 5 1 1 31734
0 31736 7 1 2 47880 48442
0 31737 7 1 2 47924 31736
0 31738 5 1 1 31737
0 31739 7 1 2 53688 49219
0 31740 7 1 2 47542 31739
0 31741 5 1 1 31740
0 31742 7 1 2 31738 31741
0 31743 5 1 1 31742
0 31744 7 1 2 43588 31743
0 31745 5 1 1 31744
0 31746 7 1 2 49693 49220
0 31747 7 1 2 59200 31746
0 31748 5 1 1 31747
0 31749 7 1 2 31745 31748
0 31750 5 1 1 31749
0 31751 7 1 2 48240 31750
0 31752 5 1 1 31751
0 31753 7 1 2 43771 41678
0 31754 7 1 2 64547 31753
0 31755 7 1 2 52287 31754
0 31756 5 1 1 31755
0 31757 7 1 2 31752 31756
0 31758 5 1 1 31757
0 31759 7 1 2 42711 31758
0 31760 5 1 1 31759
0 31761 7 1 2 43589 56223
0 31762 5 1 1 31761
0 31763 7 1 2 63362 31762
0 31764 5 1 1 31763
0 31765 7 1 2 43439 31764
0 31766 5 1 1 31765
0 31767 7 1 2 43590 63364
0 31768 5 1 1 31767
0 31769 7 1 2 31766 31768
0 31770 5 1 1 31769
0 31771 7 1 2 60792 55794
0 31772 7 1 2 31770 31771
0 31773 5 1 1 31772
0 31774 7 1 2 31760 31773
0 31775 5 3 1 31774
0 31776 7 1 2 54003 66867
0 31777 5 1 1 31776
0 31778 7 1 2 31735 31777
0 31779 5 1 1 31778
0 31780 7 1 2 66338 31779
0 31781 5 1 1 31780
0 31782 7 1 2 60225 66121
0 31783 7 1 2 64579 50149
0 31784 7 1 2 31782 31783
0 31785 7 1 2 59102 60161
0 31786 7 1 2 31784 31785
0 31787 7 1 2 66621 31786
0 31788 5 1 1 31787
0 31789 7 1 2 31781 31788
0 31790 7 1 2 31712 31789
0 31791 7 1 2 31662 31790
0 31792 7 1 2 31554 31791
0 31793 5 1 1 31792
0 31794 7 1 2 58029 31793
0 31795 5 1 1 31794
0 31796 7 1 2 46434 52426
0 31797 7 3 2 66339 31796
0 31798 7 2 2 48130 66870
0 31799 7 1 2 51699 66873
0 31800 5 1 1 31799
0 31801 7 1 2 45189 47860
0 31802 7 1 2 64384 31801
0 31803 7 2 2 48241 66476
0 31804 7 1 2 66426 66875
0 31805 7 1 2 57329 31804
0 31806 7 1 2 31802 31805
0 31807 5 1 1 31806
0 31808 7 1 2 31800 31807
0 31809 5 1 1 31808
0 31810 7 1 2 49057 31809
0 31811 5 1 1 31810
0 31812 7 1 2 56907 54882
0 31813 7 1 2 66750 31812
0 31814 7 3 2 57212 52787
0 31815 7 1 2 66427 66877
0 31816 7 1 2 31813 31815
0 31817 5 1 1 31816
0 31818 7 1 2 49986 57153
0 31819 7 1 2 66871 31818
0 31820 5 1 1 31819
0 31821 7 1 2 31817 31820
0 31822 5 1 1 31821
0 31823 7 1 2 52934 31822
0 31824 5 1 1 31823
0 31825 7 1 2 48937 66872
0 31826 5 1 1 31825
0 31827 7 1 2 65432 65236
0 31828 7 1 2 58933 57330
0 31829 7 1 2 31827 31828
0 31830 5 1 1 31829
0 31831 7 1 2 31826 31830
0 31832 5 1 1 31831
0 31833 7 1 2 57102 31832
0 31834 5 1 1 31833
0 31835 7 1 2 44134 49608
0 31836 7 1 2 54703 31835
0 31837 7 1 2 64560 56128
0 31838 7 1 2 31836 31837
0 31839 7 1 2 66352 31838
0 31840 5 1 1 31839
0 31841 7 1 2 49365 49130
0 31842 7 1 2 66874 31841
0 31843 5 1 1 31842
0 31844 7 1 2 31840 31843
0 31845 7 1 2 31834 31844
0 31846 7 1 2 31824 31845
0 31847 7 1 2 31811 31846
0 31848 5 1 1 31847
0 31849 7 1 2 53784 31848
0 31850 5 1 1 31849
0 31851 7 2 2 57272 56420
0 31852 5 6 1 66880
0 31853 7 5 2 52869 57331
0 31854 7 1 2 62420 64127
0 31855 7 1 2 66888 31854
0 31856 5 1 1 31855
0 31857 7 1 2 66882 31856
0 31858 5 1 1 31857
0 31859 7 1 2 43440 31858
0 31860 5 1 1 31859
0 31861 7 1 2 46435 52407
0 31862 7 1 2 62767 31861
0 31863 7 1 2 56488 31862
0 31864 5 1 1 31863
0 31865 7 1 2 31860 31864
0 31866 5 1 1 31865
0 31867 7 1 2 52935 31866
0 31868 5 1 1 31867
0 31869 7 2 2 66462 50402
0 31870 7 2 2 63777 56432
0 31871 7 3 2 66893 66895
0 31872 5 2 1 66897
0 31873 7 1 2 48242 50737
0 31874 7 1 2 65860 31873
0 31875 7 1 2 62682 31874
0 31876 5 1 1 31875
0 31877 7 1 2 66900 31876
0 31878 5 2 1 31877
0 31879 7 1 2 41148 66901
0 31880 5 1 1 31879
0 31881 7 1 2 43441 31880
0 31882 7 1 2 66902 31881
0 31883 5 1 1 31882
0 31884 7 2 2 65861 58943
0 31885 5 1 1 66904
0 31886 7 1 2 52427 61673
0 31887 5 1 1 31886
0 31888 7 1 2 31885 31887
0 31889 5 1 1 31888
0 31890 7 1 2 57103 31889
0 31891 5 1 1 31890
0 31892 7 1 2 52408 57273
0 31893 7 1 2 52756 31892
0 31894 7 1 2 55435 31893
0 31895 5 1 1 31894
0 31896 7 1 2 31891 31895
0 31897 7 1 2 31883 31896
0 31898 7 1 2 31868 31897
0 31899 5 1 1 31898
0 31900 7 1 2 53785 31899
0 31901 5 1 1 31900
0 31902 7 1 2 51433 49283
0 31903 7 1 2 66792 31902
0 31904 5 1 1 31903
0 31905 7 1 2 50810 53468
0 31906 5 1 1 31905
0 31907 7 1 2 31270 31906
0 31908 5 1 1 31907
0 31909 7 1 2 51554 31908
0 31910 5 1 1 31909
0 31911 7 1 2 66766 31910
0 31912 5 1 1 31911
0 31913 7 1 2 46299 31912
0 31914 5 1 1 31913
0 31915 7 1 2 48523 66094
0 31916 5 1 1 31915
0 31917 7 1 2 46300 66759
0 31918 5 1 1 31917
0 31919 7 1 2 31916 31918
0 31920 5 1 1 31919
0 31921 7 1 2 49221 31920
0 31922 5 1 1 31921
0 31923 7 1 2 53482 57712
0 31924 5 1 1 31923
0 31925 7 1 2 31922 31924
0 31926 7 1 2 31914 31925
0 31927 5 1 1 31926
0 31928 7 1 2 57274 31927
0 31929 5 1 1 31928
0 31930 7 1 2 31904 31929
0 31931 5 1 1 31930
0 31932 7 1 2 56263 31931
0 31933 5 1 1 31932
0 31934 7 1 2 47536 63436
0 31935 7 1 2 57799 31934
0 31936 7 1 2 55521 31935
0 31937 5 1 1 31936
0 31938 7 1 2 31933 31937
0 31939 5 1 1 31938
0 31940 7 1 2 47353 66853
0 31941 7 1 2 31939 31940
0 31942 5 1 1 31941
0 31943 7 1 2 31901 31942
0 31944 5 1 1 31943
0 31945 7 1 2 45190 31944
0 31946 5 1 1 31945
0 31947 7 1 2 55522 57549
0 31948 5 1 1 31947
0 31949 7 3 2 49136 51399
0 31950 7 1 2 66906 59831
0 31951 5 1 1 31950
0 31952 7 1 2 31948 31951
0 31953 5 1 1 31952
0 31954 7 1 2 47354 31953
0 31955 5 1 1 31954
0 31956 7 1 2 31218 31955
0 31957 5 1 1 31956
0 31958 7 1 2 41988 31957
0 31959 5 1 1 31958
0 31960 7 1 2 49222 55523
0 31961 5 1 1 31960
0 31962 7 1 2 44135 56495
0 31963 5 1 1 31962
0 31964 7 1 2 31961 31963
0 31965 5 1 1 31964
0 31966 7 1 2 49609 31965
0 31967 5 1 1 31966
0 31968 7 1 2 62226 66518
0 31969 5 1 1 31968
0 31970 7 1 2 31967 31969
0 31971 5 1 1 31970
0 31972 7 1 2 47427 31971
0 31973 5 1 1 31972
0 31974 7 1 2 31959 31973
0 31975 5 1 1 31974
0 31976 7 1 2 49356 31975
0 31977 5 1 1 31976
0 31978 7 1 2 65456 58507
0 31979 5 1 1 31978
0 31980 7 1 2 45785 62671
0 31981 5 1 1 31980
0 31982 7 1 2 31979 31981
0 31983 5 1 1 31982
0 31984 7 1 2 49610 31983
0 31985 5 1 1 31984
0 31986 7 1 2 63417 66777
0 31987 5 1 1 31986
0 31988 7 1 2 31985 31987
0 31989 5 1 1 31988
0 31990 7 1 2 43028 50385
0 31991 7 1 2 31989 31990
0 31992 5 1 1 31991
0 31993 7 1 2 31977 31992
0 31994 5 1 1 31993
0 31995 7 1 2 43143 31994
0 31996 5 1 1 31995
0 31997 7 3 2 61160 60099
0 31998 7 1 2 49841 51555
0 31999 7 1 2 59231 31998
0 32000 7 1 2 66909 31999
0 32001 7 1 2 61200 32000
0 32002 5 1 1 32001
0 32003 7 1 2 31996 32002
0 32004 5 1 1 32003
0 32005 7 1 2 43591 32004
0 32006 5 1 1 32005
0 32007 7 1 2 66095 57718
0 32008 5 1 1 32007
0 32009 7 2 2 51650 60811
0 32010 7 1 2 53469 66912
0 32011 5 1 1 32010
0 32012 7 1 2 32008 32011
0 32013 5 1 1 32012
0 32014 7 1 2 48938 32013
0 32015 5 1 1 32014
0 32016 7 1 2 44968 50615
0 32017 7 1 2 58790 32016
0 32018 7 1 2 66772 32017
0 32019 5 1 1 32018
0 32020 7 1 2 32015 32019
0 32021 5 1 1 32020
0 32022 7 1 2 47428 59932
0 32023 7 1 2 32021 32022
0 32024 5 1 1 32023
0 32025 7 1 2 32006 32024
0 32026 5 1 1 32025
0 32027 7 2 2 43261 32026
0 32028 7 1 2 66248 66914
0 32029 5 1 1 32028
0 32030 7 1 2 31946 32029
0 32031 5 1 1 32030
0 32032 7 1 2 44350 32031
0 32033 5 1 1 32032
0 32034 7 1 2 66529 66915
0 32035 5 1 1 32034
0 32036 7 1 2 66854 66858
0 32037 5 1 1 32036
0 32038 7 1 2 56891 51427
0 32039 7 1 2 66862 32038
0 32040 5 1 1 32039
0 32041 7 1 2 32037 32040
0 32042 5 1 1 32041
0 32043 7 1 2 40884 32042
0 32044 5 1 1 32043
0 32045 7 1 2 60604 66864
0 32046 5 1 1 32045
0 32047 7 1 2 32044 32046
0 32048 5 1 1 32047
0 32049 7 1 2 47429 32048
0 32050 5 1 1 32049
0 32051 7 1 2 61780 54865
0 32052 7 1 2 55778 32051
0 32053 7 1 2 63897 32052
0 32054 5 1 1 32053
0 32055 7 1 2 32050 32054
0 32056 5 1 1 32055
0 32057 7 1 2 59666 48279
0 32058 7 1 2 32056 32057
0 32059 5 1 1 32058
0 32060 7 1 2 61725 66866
0 32061 5 1 1 32060
0 32062 7 1 2 50754 53583
0 32063 7 1 2 61192 52200
0 32064 7 1 2 32062 32063
0 32065 7 2 2 52643 57213
0 32066 7 1 2 58944 66916
0 32067 7 1 2 32064 32066
0 32068 5 1 1 32067
0 32069 7 1 2 32061 32068
0 32070 7 1 2 32059 32069
0 32071 5 1 1 32070
0 32072 7 1 2 45191 32071
0 32073 5 1 1 32072
0 32074 7 2 2 59718 63580
0 32075 7 1 2 66918 66868
0 32076 5 1 1 32075
0 32077 7 1 2 32073 32076
0 32078 5 1 1 32077
0 32079 7 1 2 44351 32078
0 32080 5 1 1 32079
0 32081 7 1 2 66689 66869
0 32082 5 1 1 32081
0 32083 7 1 2 43442 66835
0 32084 5 1 1 32083
0 32085 7 1 2 48314 66827
0 32086 7 1 2 55542 32085
0 32087 7 1 2 66606 32086
0 32088 5 1 1 32087
0 32089 7 1 2 32084 32088
0 32090 5 1 1 32089
0 32091 7 1 2 63581 32090
0 32092 5 1 1 32091
0 32093 7 1 2 43443 66841
0 32094 5 1 1 32093
0 32095 7 1 2 65207 66849
0 32096 5 1 1 32095
0 32097 7 1 2 32094 32096
0 32098 5 1 1 32097
0 32099 7 1 2 64683 60511
0 32100 7 1 2 56062 32099
0 32101 7 1 2 32098 32100
0 32102 5 1 1 32101
0 32103 7 1 2 32092 32102
0 32104 5 1 1 32103
0 32105 7 1 2 52936 32104
0 32106 5 1 1 32105
0 32107 7 1 2 32082 32106
0 32108 7 1 2 32080 32107
0 32109 5 1 1 32108
0 32110 7 1 2 58030 32109
0 32111 5 1 1 32110
0 32112 7 2 2 58031 58805
0 32113 5 1 1 66920
0 32114 7 1 2 66762 32113
0 32115 5 1 1 32114
0 32116 7 2 2 52288 64537
0 32117 7 1 2 66760 66921
0 32118 5 1 1 32117
0 32119 7 1 2 66922 32118
0 32120 7 2 2 32115 32119
0 32121 7 1 2 66530 66924
0 32122 5 1 1 32121
0 32123 7 1 2 66249 66925
0 32124 5 1 1 32123
0 32125 7 2 2 63010 58784
0 32126 5 1 1 66926
0 32127 7 1 2 6239 32126
0 32128 5 1 1 32127
0 32129 7 1 2 62444 32128
0 32130 5 1 1 32129
0 32131 7 1 2 51318 55003
0 32132 7 1 2 63833 32131
0 32133 5 1 1 32132
0 32134 7 1 2 32130 32133
0 32135 5 1 1 32134
0 32136 7 1 2 44444 32135
0 32137 5 1 1 32136
0 32138 7 2 2 52384 63834
0 32139 7 1 2 52516 66928
0 32140 5 1 1 32139
0 32141 7 1 2 43772 32140
0 32142 7 1 2 32137 32141
0 32143 5 1 1 32142
0 32144 7 1 2 40113 31622
0 32145 5 1 1 32144
0 32146 7 1 2 41532 53748
0 32147 5 1 1 32146
0 32148 7 1 2 3485 32147
0 32149 5 2 1 32148
0 32150 7 1 2 57305 66930
0 32151 5 1 1 32150
0 32152 7 1 2 51319 66929
0 32153 5 1 1 32152
0 32154 7 1 2 9382 32153
0 32155 7 1 2 32151 32154
0 32156 5 1 1 32155
0 32157 7 1 2 32145 32156
0 32158 7 1 2 32143 32157
0 32159 5 1 1 32158
0 32160 7 2 2 41406 57438
0 32161 7 1 2 52670 66932
0 32162 7 1 2 66793 32161
0 32163 5 1 1 32162
0 32164 7 1 2 40673 32163
0 32165 7 1 2 32159 32164
0 32166 5 1 1 32165
0 32167 7 1 2 45340 66927
0 32168 5 1 1 32167
0 32169 7 1 2 64074 57306
0 32170 5 1 1 32169
0 32171 7 1 2 32168 32170
0 32172 5 1 1 32171
0 32173 7 1 2 32172 66851
0 32174 5 1 1 32173
0 32175 7 1 2 59330 63835
0 32176 7 1 2 41149 58128
0 32177 5 1 1 32176
0 32178 7 1 2 66823 32177
0 32179 7 1 2 32175 32178
0 32180 5 1 1 32179
0 32181 7 1 2 32174 32180
0 32182 5 1 1 32181
0 32183 7 1 2 41533 32182
0 32184 5 1 1 32183
0 32185 7 1 2 52627 50894
0 32186 7 1 2 62187 32185
0 32187 7 1 2 57294 32186
0 32188 7 1 2 53779 32187
0 32189 5 1 1 32188
0 32190 7 1 2 43958 32189
0 32191 7 1 2 32184 32190
0 32192 5 1 1 32191
0 32193 7 1 2 45192 32192
0 32194 7 1 2 32166 32193
0 32195 5 1 1 32194
0 32196 7 1 2 32124 32195
0 32197 5 1 1 32196
0 32198 7 1 2 44352 32197
0 32199 5 1 1 32198
0 32200 7 1 2 32122 32199
0 32201 5 1 1 32200
0 32202 7 1 2 49223 32201
0 32203 5 1 1 32202
0 32204 7 1 2 51556 66587
0 32205 5 1 1 32204
0 32206 7 1 2 62611 58791
0 32207 5 2 1 32206
0 32208 7 1 2 32205 66934
0 32209 5 1 1 32208
0 32210 7 2 2 43959 32209
0 32211 5 1 1 66936
0 32212 7 2 2 40674 48604
0 32213 7 1 2 66938 64216
0 32214 5 1 1 32213
0 32215 7 1 2 32211 32214
0 32216 5 1 1 32215
0 32217 7 1 2 58312 32216
0 32218 5 1 1 32217
0 32219 7 1 2 50554 57713
0 32220 7 1 2 58792 32219
0 32221 5 1 1 32220
0 32222 7 1 2 32218 32221
0 32223 5 1 1 32222
0 32224 7 1 2 66607 32223
0 32225 5 1 1 32224
0 32226 7 1 2 65175 61207
0 32227 7 1 2 59761 32226
0 32228 7 2 2 59511 58725
0 32229 7 1 2 60999 66940
0 32230 7 1 2 32227 32229
0 32231 5 1 1 32230
0 32232 7 1 2 32225 32231
0 32233 5 1 1 32232
0 32234 7 1 2 43144 32233
0 32235 5 1 1 32234
0 32236 7 1 2 54826 66617
0 32237 7 1 2 48393 32236
0 32238 7 1 2 57307 66362
0 32239 7 1 2 32237 32238
0 32240 5 1 1 32239
0 32241 7 1 2 32235 32240
0 32242 5 1 1 32241
0 32243 7 1 2 50924 32242
0 32244 5 1 1 32243
0 32245 7 2 2 60850 57390
0 32246 5 1 1 66942
0 32247 7 1 2 66744 66452
0 32248 7 1 2 66943 32247
0 32249 5 1 1 32248
0 32250 7 1 2 66402 63005
0 32251 5 1 1 32250
0 32252 7 1 2 29220 32251
0 32253 5 1 1 32252
0 32254 7 1 2 46166 32253
0 32255 5 1 1 32254
0 32256 7 1 2 40675 64363
0 32257 5 1 1 32256
0 32258 7 1 2 32255 32257
0 32259 5 1 1 32258
0 32260 7 1 2 59667 63787
0 32261 7 1 2 32259 32260
0 32262 5 1 1 32261
0 32263 7 1 2 32249 32262
0 32264 5 1 1 32263
0 32265 7 1 2 64684 32264
0 32266 5 1 1 32265
0 32267 7 2 2 45786 66923
0 32268 7 3 2 46590 51557
0 32269 7 1 2 66209 66946
0 32270 7 1 2 66944 32269
0 32271 5 1 1 32270
0 32272 7 1 2 32266 32271
0 32273 5 1 1 32272
0 32274 7 1 2 54366 32273
0 32275 5 1 1 32274
0 32276 7 1 2 48319 66878
0 32277 5 1 1 32276
0 32278 7 1 2 63795 32277
0 32279 5 1 1 32278
0 32280 7 1 2 43444 32279
0 32281 5 1 1 32280
0 32282 7 1 2 52409 63788
0 32283 5 1 1 32282
0 32284 7 1 2 32281 32283
0 32285 5 1 1 32284
0 32286 7 1 2 66560 32285
0 32287 5 1 1 32286
0 32288 7 1 2 65972 53315
0 32289 7 1 2 58863 32288
0 32290 7 1 2 66268 60512
0 32291 7 1 2 32289 32290
0 32292 5 1 1 32291
0 32293 7 1 2 32287 32292
0 32294 5 1 1 32293
0 32295 7 1 2 64685 32294
0 32296 5 1 1 32295
0 32297 7 1 2 60977 66947
0 32298 7 1 2 66945 32297
0 32299 5 1 1 32298
0 32300 7 1 2 32296 32299
0 32301 5 1 1 32300
0 32302 7 1 2 65553 32301
0 32303 5 1 1 32302
0 32304 7 1 2 32275 32303
0 32305 7 1 2 32244 32304
0 32306 7 1 2 32203 32305
0 32307 5 1 1 32306
0 32308 7 1 2 49058 32307
0 32309 5 1 1 32308
0 32310 7 1 2 32111 32309
0 32311 7 1 2 32035 32310
0 32312 7 1 2 32033 32311
0 32313 5 1 1 32312
0 32314 7 1 2 55102 32313
0 32315 5 1 1 32314
0 32316 7 1 2 31850 32315
0 32317 7 1 2 31795 32316
0 32318 7 1 2 31356 32317
0 32319 5 1 1 32318
0 32320 7 1 2 47057 32319
0 32321 5 1 1 32320
0 32322 7 3 2 65046 64033
0 32323 7 1 2 66949 49284
0 32324 5 1 1 32323
0 32325 7 1 2 53333 64643
0 32326 5 1 1 32325
0 32327 7 1 2 32324 32326
0 32328 5 1 1 32327
0 32329 7 1 2 44285 32328
0 32330 5 1 1 32329
0 32331 7 2 2 40676 63129
0 32332 7 1 2 62768 64385
0 32333 7 1 2 66952 32332
0 32334 5 1 1 32333
0 32335 7 1 2 32330 32334
0 32336 5 1 1 32335
0 32337 7 1 2 49059 32336
0 32338 5 1 1 32337
0 32339 7 2 2 46301 62928
0 32340 7 1 2 56489 66954
0 32341 5 1 1 32340
0 32342 7 1 2 66950 61940
0 32343 5 1 1 32342
0 32344 7 2 2 63155 66843
0 32345 7 1 2 64969 66956
0 32346 5 1 1 32345
0 32347 7 1 2 32343 32346
0 32348 5 1 1 32347
0 32349 7 1 2 48939 32348
0 32350 5 1 1 32349
0 32351 7 1 2 32341 32350
0 32352 7 1 2 32338 32351
0 32353 5 1 1 32352
0 32354 7 1 2 45193 32353
0 32355 5 1 1 32354
0 32356 7 1 2 49611 59007
0 32357 7 1 2 66844 32356
0 32358 7 1 2 66787 32357
0 32359 5 1 1 32358
0 32360 7 1 2 32355 32359
0 32361 5 1 1 32360
0 32362 7 1 2 44353 32361
0 32363 5 1 1 32362
0 32364 7 1 2 65349 66567
0 32365 7 1 2 64742 32364
0 32366 5 1 1 32365
0 32367 7 1 2 32363 32366
0 32368 5 1 1 32367
0 32369 7 1 2 52937 32368
0 32370 5 1 1 32369
0 32371 7 1 2 48970 66951
0 32372 5 1 1 32371
0 32373 7 1 2 52644 63163
0 32374 5 1 1 32373
0 32375 7 1 2 32372 32374
0 32376 5 1 1 32375
0 32377 7 1 2 44286 32376
0 32378 5 1 1 32377
0 32379 7 1 2 62081 59365
0 32380 7 1 2 49095 32379
0 32381 5 1 1 32380
0 32382 7 1 2 32378 32381
0 32383 5 1 1 32382
0 32384 7 1 2 53535 32383
0 32385 5 1 1 32384
0 32386 7 3 2 49285 63084
0 32387 7 1 2 63765 66958
0 32388 5 1 1 32387
0 32389 7 1 2 32385 32388
0 32390 5 1 1 32389
0 32391 7 1 2 45194 32390
0 32392 5 1 1 32391
0 32393 7 1 2 44969 59308
0 32394 7 1 2 66959 32393
0 32395 5 1 1 32394
0 32396 7 1 2 32392 32395
0 32397 5 1 1 32396
0 32398 7 1 2 44354 32397
0 32399 5 1 1 32398
0 32400 7 1 2 44970 66446
0 32401 7 1 2 66960 32400
0 32402 5 1 1 32401
0 32403 7 1 2 32399 32402
0 32404 5 1 1 32403
0 32405 7 1 2 49060 32404
0 32406 5 1 1 32405
0 32407 7 1 2 52144 61914
0 32408 5 1 1 32407
0 32409 7 1 2 53536 63152
0 32410 7 1 2 65047 32409
0 32411 5 1 1 32410
0 32412 7 1 2 32408 32411
0 32413 5 1 1 32412
0 32414 7 1 2 48940 32413
0 32415 5 1 1 32414
0 32416 7 2 2 41767 62929
0 32417 7 1 2 66961 66894
0 32418 5 1 1 32417
0 32419 7 1 2 32415 32418
0 32420 5 1 1 32419
0 32421 7 1 2 43029 32420
0 32422 5 1 1 32421
0 32423 7 1 2 49325 64478
0 32424 5 1 1 32423
0 32425 7 2 2 46946 50898
0 32426 5 2 1 66963
0 32427 7 1 2 66633 66965
0 32428 5 1 1 32427
0 32429 7 1 2 32424 32428
0 32430 5 4 1 32429
0 32431 7 1 2 60298 49357
0 32432 7 1 2 51700 32431
0 32433 7 1 2 66967 32432
0 32434 5 1 1 32433
0 32435 7 1 2 32422 32434
0 32436 5 1 1 32435
0 32437 7 1 2 45195 32436
0 32438 5 1 1 32437
0 32439 7 2 2 40677 49120
0 32440 7 2 2 63077 66971
0 32441 7 3 2 59303 49366
0 32442 7 1 2 61936 66975
0 32443 7 1 2 66973 32442
0 32444 5 1 1 32443
0 32445 7 1 2 32438 32444
0 32446 5 1 1 32445
0 32447 7 1 2 44355 32446
0 32448 5 1 1 32447
0 32449 7 1 2 66384 62747
0 32450 7 1 2 66974 32449
0 32451 5 1 1 32450
0 32452 7 1 2 32448 32451
0 32453 5 1 1 32452
0 32454 7 1 2 46167 32453
0 32455 5 1 1 32454
0 32456 7 1 2 32406 32455
0 32457 7 1 2 32370 32456
0 32458 5 1 1 32457
0 32459 7 1 2 46436 32458
0 32460 5 1 1 32459
0 32461 7 5 2 43145 49777
0 32462 7 2 2 58987 66978
0 32463 5 1 1 66983
0 32464 7 1 2 46517 66984
0 32465 5 1 1 32464
0 32466 7 1 2 49778 61746
0 32467 5 1 1 32466
0 32468 7 1 2 61688 32467
0 32469 5 1 1 32468
0 32470 7 1 2 55103 32469
0 32471 5 1 1 32470
0 32472 7 1 2 32471 61592
0 32473 7 1 2 32465 32472
0 32474 5 1 1 32473
0 32475 7 1 2 45196 32474
0 32476 5 1 1 32475
0 32477 7 1 2 66595 32476
0 32478 5 1 1 32477
0 32479 7 1 2 44356 32478
0 32480 5 1 1 32479
0 32481 7 1 2 54182 65232
0 32482 5 2 1 32481
0 32483 7 1 2 32480 66985
0 32484 5 1 1 32483
0 32485 7 1 2 57104 32484
0 32486 5 1 1 32485
0 32487 7 1 2 59220 57531
0 32488 5 1 1 32487
0 32489 7 1 2 59206 57755
0 32490 5 1 1 32489
0 32491 7 1 2 32488 32490
0 32492 5 1 1 32491
0 32493 7 1 2 44287 32492
0 32494 5 1 1 32493
0 32495 7 1 2 29138 32494
0 32496 5 1 1 32495
0 32497 7 1 2 57110 32496
0 32498 5 1 1 32497
0 32499 7 1 2 55104 57154
0 32500 5 1 1 32499
0 32501 7 1 2 65548 64040
0 32502 5 1 1 32501
0 32503 7 1 2 32500 32502
0 32504 5 1 1 32503
0 32505 7 1 2 52772 32504
0 32506 5 1 1 32505
0 32507 7 1 2 32498 32506
0 32508 5 1 1 32507
0 32509 7 1 2 65365 66979
0 32510 7 1 2 32508 32509
0 32511 5 1 1 32510
0 32512 7 1 2 32486 32511
0 32513 7 1 2 32460 32512
0 32514 5 1 1 32513
0 32515 7 1 2 53780 32514
0 32516 5 1 1 32515
0 32517 7 3 2 49779 48593
0 32518 7 2 2 52234 66987
0 32519 5 1 1 66990
0 32520 7 1 2 44971 59893
0 32521 7 1 2 65048 32520
0 32522 5 1 1 32521
0 32523 7 1 2 32519 32522
0 32524 5 1 1 32523
0 32525 7 1 2 44219 32524
0 32526 5 1 1 32525
0 32527 7 1 2 45061 56777
0 32528 7 1 2 66988 32527
0 32529 5 1 1 32528
0 32530 7 1 2 32526 32529
0 32531 5 1 1 32530
0 32532 7 1 2 44136 32531
0 32533 5 1 1 32532
0 32534 7 1 2 49780 58883
0 32535 5 1 1 32534
0 32536 7 1 2 32533 32535
0 32537 5 1 1 32536
0 32538 7 1 2 49612 32537
0 32539 5 1 1 32538
0 32540 7 1 2 48524 66989
0 32541 7 1 2 56759 32540
0 32542 5 1 1 32541
0 32543 7 1 2 32539 32542
0 32544 5 1 1 32543
0 32545 7 1 2 45989 32544
0 32546 5 1 1 32545
0 32547 7 4 2 58032 49224
0 32548 7 2 2 49061 66992
0 32549 7 2 2 48594 53584
0 32550 7 1 2 66996 66998
0 32551 5 1 1 32550
0 32552 7 1 2 32546 32551
0 32553 5 1 1 32552
0 32554 7 1 2 48838 32553
0 32555 5 1 1 32554
0 32556 7 1 2 49062 57550
0 32557 5 1 1 32556
0 32558 7 1 2 32557 21498
0 32559 5 1 1 32558
0 32560 7 1 2 52013 66999
0 32561 7 1 2 32559 32560
0 32562 5 1 1 32561
0 32563 7 1 2 32555 32562
0 32564 5 1 1 32563
0 32565 7 1 2 57214 32564
0 32566 5 1 1 32565
0 32567 7 1 2 41407 57983
0 32568 7 1 2 66997 32567
0 32569 5 1 1 32568
0 32570 7 1 2 32566 32569
0 32571 5 1 1 32570
0 32572 7 1 2 55105 32571
0 32573 5 1 1 32572
0 32574 7 1 2 66991 55436
0 32575 5 1 1 32574
0 32576 7 1 2 55193 63357
0 32577 7 1 2 65049 32576
0 32578 5 1 1 32577
0 32579 7 1 2 32575 32578
0 32580 5 1 1 32579
0 32581 7 1 2 43146 32580
0 32582 5 1 1 32581
0 32583 7 2 2 64489 66968
0 32584 7 1 2 67000 56979
0 32585 5 1 1 32584
0 32586 7 1 2 32582 32585
0 32587 5 1 1 32586
0 32588 7 1 2 55554 32587
0 32589 5 1 1 32588
0 32590 7 1 2 55555 61165
0 32591 7 1 2 67001 32590
0 32592 5 1 1 32591
0 32593 7 1 2 58033 65213
0 32594 5 2 1 32593
0 32595 7 1 2 55422 56825
0 32596 5 1 1 32595
0 32597 7 1 2 67002 32596
0 32598 5 1 1 32597
0 32599 7 1 2 49063 65050
0 32600 7 1 2 32598 32599
0 32601 5 1 1 32600
0 32602 7 1 2 32592 32601
0 32603 5 1 1 32602
0 32604 7 1 2 49225 32603
0 32605 5 1 1 32604
0 32606 7 1 2 52517 50075
0 32607 7 1 2 62583 32606
0 32608 7 1 2 64041 51230
0 32609 7 1 2 32607 32608
0 32610 5 1 1 32609
0 32611 7 1 2 32605 32610
0 32612 7 1 2 32589 32611
0 32613 5 1 1 32612
0 32614 7 1 2 60299 32613
0 32615 5 1 1 32614
0 32616 7 1 2 32573 32615
0 32617 5 1 1 32616
0 32618 7 1 2 64686 32617
0 32619 5 1 1 32618
0 32620 7 1 2 66191 51630
0 32621 5 1 1 32620
0 32622 7 1 2 58699 32621
0 32623 5 1 1 32622
0 32624 7 1 2 41150 32623
0 32625 5 1 1 32624
0 32626 7 1 2 40290 12792
0 32627 7 1 2 51634 32626
0 32628 7 1 2 50024 32627
0 32629 5 1 1 32628
0 32630 7 1 2 32625 32629
0 32631 5 1 1 32630
0 32632 7 1 2 43445 32631
0 32633 5 1 1 32632
0 32634 7 1 2 62295 50010
0 32635 5 1 1 32634
0 32636 7 2 2 41151 50011
0 32637 5 1 1 67004
0 32638 7 1 2 65651 57413
0 32639 5 1 1 32638
0 32640 7 1 2 32637 32639
0 32641 5 1 1 32640
0 32642 7 1 2 41989 32641
0 32643 5 1 1 32642
0 32644 7 1 2 41152 49987
0 32645 5 1 1 32644
0 32646 7 1 2 50016 32645
0 32647 5 2 1 32646
0 32648 7 1 2 45341 52410
0 32649 7 1 2 67006 32648
0 32650 5 1 1 32649
0 32651 7 1 2 32643 32650
0 32652 5 1 1 32651
0 32653 7 1 2 40114 32652
0 32654 5 1 1 32653
0 32655 7 1 2 32635 32654
0 32656 7 1 2 32633 32655
0 32657 5 1 1 32656
0 32658 7 1 2 58619 32657
0 32659 5 1 1 32658
0 32660 7 1 2 5337 52870
0 32661 7 1 2 567 32660
0 32662 7 1 2 49173 32661
0 32663 7 1 2 65051 32662
0 32664 5 1 1 32663
0 32665 7 1 2 32659 32664
0 32666 5 1 1 32665
0 32667 7 1 2 46437 32666
0 32668 5 1 1 32667
0 32669 7 1 2 66320 66980
0 32670 5 1 1 32669
0 32671 7 1 2 57660 32670
0 32672 7 1 2 32668 32671
0 32673 5 1 1 32672
0 32674 7 1 2 51558 66318
0 32675 5 1 1 32674
0 32676 7 1 2 32675 21849
0 32677 5 1 1 32676
0 32678 7 1 2 66981 32677
0 32679 5 1 1 32678
0 32680 7 1 2 57672 32679
0 32681 5 1 1 32680
0 32682 7 1 2 32681 57536
0 32683 7 1 2 32673 32682
0 32684 5 1 1 32683
0 32685 7 1 2 57961 64732
0 32686 5 1 1 32685
0 32687 7 1 2 32684 32686
0 32688 5 1 1 32687
0 32689 7 1 2 45197 32688
0 32690 5 1 1 32689
0 32691 7 1 2 59309 59016
0 32692 7 1 2 60513 32691
0 32693 5 1 1 32692
0 32694 7 1 2 32690 32693
0 32695 5 1 1 32694
0 32696 7 1 2 44357 32695
0 32697 5 1 1 32696
0 32698 7 1 2 65346 60514
0 32699 7 1 2 66785 32698
0 32700 5 1 1 32699
0 32701 7 1 2 32697 32700
0 32702 5 1 1 32701
0 32703 7 1 2 55267 55514
0 32704 5 3 1 32703
0 32705 7 1 2 58034 67008
0 32706 7 1 2 32702 32705
0 32707 5 1 1 32706
0 32708 7 1 2 65052 63815
0 32709 5 1 1 32708
0 32710 7 1 2 55106 66982
0 32711 5 1 1 32710
0 32712 7 1 2 32709 32711
0 32713 5 1 1 32712
0 32714 7 1 2 48941 32713
0 32715 5 1 1 32714
0 32716 7 1 2 32463 32715
0 32717 5 1 1 32716
0 32718 7 1 2 46518 32717
0 32719 5 1 1 32718
0 32720 7 1 2 32719 18479
0 32721 5 1 1 32720
0 32722 7 1 2 45198 32721
0 32723 5 1 1 32722
0 32724 7 1 2 66596 32723
0 32725 5 1 1 32724
0 32726 7 1 2 44358 32725
0 32727 5 1 1 32726
0 32728 7 1 2 66986 32727
0 32729 5 1 1 32728
0 32730 7 1 2 65465 66993
0 32731 7 1 2 32729 32730
0 32732 5 1 1 32731
0 32733 7 1 2 32707 32732
0 32734 7 1 2 32619 32733
0 32735 7 1 2 32516 32734
0 32736 5 1 1 32735
0 32737 7 1 2 47071 47150
0 32738 7 1 2 32736 32737
0 32739 5 1 1 32738
0 32740 7 1 2 65071 62574
0 32741 5 1 1 32740
0 32742 7 1 2 55941 51707
0 32743 5 1 1 32742
0 32744 7 1 2 32741 32743
0 32745 5 1 1 32744
0 32746 7 1 2 59057 32745
0 32747 5 1 1 32746
0 32748 7 1 2 59960 60884
0 32749 7 1 2 60485 32748
0 32750 5 1 1 32749
0 32751 7 1 2 32747 32750
0 32752 5 1 1 32751
0 32753 7 1 2 41990 32752
0 32754 5 1 1 32753
0 32755 7 1 2 65477 66576
0 32756 5 1 1 32755
0 32757 7 1 2 32754 32756
0 32758 5 1 1 32757
0 32759 7 1 2 40678 32758
0 32760 5 1 1 32759
0 32761 7 1 2 59961 52294
0 32762 5 1 1 32761
0 32763 7 1 2 52416 59982
0 32764 5 1 1 32763
0 32765 7 1 2 32762 32764
0 32766 5 1 1 32765
0 32767 7 1 2 47129 32766
0 32768 5 1 1 32767
0 32769 7 1 2 59962 65475
0 32770 5 1 1 32769
0 32771 7 1 2 32768 32770
0 32772 5 1 1 32771
0 32773 7 1 2 58003 32772
0 32774 5 1 1 32773
0 32775 7 1 2 32760 32774
0 32776 5 1 1 32775
0 32777 7 1 2 44288 32776
0 32778 5 1 1 32777
0 32779 7 1 2 58035 65478
0 32780 5 1 1 32779
0 32781 7 1 2 43592 50702
0 32782 7 1 2 65973 66274
0 32783 7 1 2 32781 32782
0 32784 5 2 1 32783
0 32785 7 1 2 32780 67011
0 32786 5 1 1 32785
0 32787 7 1 2 59092 32786
0 32788 5 1 1 32787
0 32789 7 1 2 32778 32788
0 32790 5 1 1 32789
0 32791 7 1 2 52871 32790
0 32792 5 1 1 32791
0 32793 7 1 2 41991 52850
0 32794 5 1 1 32793
0 32795 7 1 2 59849 32794
0 32796 5 1 1 32795
0 32797 7 1 2 56209 32796
0 32798 5 1 1 32797
0 32799 7 1 2 40291 32798
0 32800 5 1 1 32799
0 32801 7 1 2 62390 32800
0 32802 5 2 1 32801
0 32803 7 1 2 58036 67013
0 32804 5 1 1 32803
0 32805 7 1 2 67012 32804
0 32806 5 1 1 32805
0 32807 7 1 2 57661 54554
0 32808 7 1 2 32806 32807
0 32809 5 1 1 32808
0 32810 7 1 2 32792 32809
0 32811 5 1 1 32810
0 32812 7 1 2 46519 32811
0 32813 5 1 1 32812
0 32814 7 2 2 43262 58037
0 32815 7 1 2 64825 59145
0 32816 5 1 1 32815
0 32817 7 2 2 56844 46636
0 32818 5 1 1 67017
0 32819 7 1 2 52814 67018
0 32820 5 1 1 32819
0 32821 7 1 2 32816 32820
0 32822 5 1 1 32821
0 32823 7 1 2 52859 32822
0 32824 5 1 1 32823
0 32825 7 1 2 47817 52872
0 32826 7 1 2 64869 32825
0 32827 5 1 1 32826
0 32828 7 1 2 32824 32827
0 32829 5 1 1 32828
0 32830 7 1 2 67015 32829
0 32831 5 1 1 32830
0 32832 7 1 2 44220 32831
0 32833 7 1 2 32813 32832
0 32834 5 1 1 32833
0 32835 7 1 2 59187 64644
0 32836 5 2 1 32835
0 32837 7 2 2 57662 63206
0 32838 5 1 1 67021
0 32839 7 1 2 67005 67022
0 32840 5 1 1 32839
0 32841 7 1 2 67019 32840
0 32842 5 1 1 32841
0 32843 7 1 2 40115 32842
0 32844 5 1 1 32843
0 32845 7 1 2 59482 67007
0 32846 5 1 1 32845
0 32847 7 1 2 45342 60057
0 32848 7 1 2 64034 32847
0 32849 5 1 1 32848
0 32850 7 1 2 67020 32849
0 32851 5 1 1 32850
0 32852 7 1 2 47818 32851
0 32853 5 1 1 32852
0 32854 7 1 2 32846 32853
0 32855 7 1 2 32844 32854
0 32856 5 1 1 32855
0 32857 7 1 2 43147 32856
0 32858 5 1 1 32857
0 32859 7 1 2 47560 49988
0 32860 5 1 1 32859
0 32861 7 1 2 41266 50012
0 32862 5 1 1 32861
0 32863 7 1 2 32860 32862
0 32864 5 1 1 32863
0 32865 7 2 2 55107 57275
0 32866 7 1 2 32864 67023
0 32867 5 1 1 32866
0 32868 7 1 2 32858 32867
0 32869 5 1 1 32868
0 32870 7 1 2 45510 32869
0 32871 5 1 1 32870
0 32872 7 2 2 54080 58089
0 32873 7 1 2 66955 67025
0 32874 5 1 1 32873
0 32875 7 1 2 32871 32874
0 32876 5 1 1 32875
0 32877 7 1 2 58038 32876
0 32878 5 1 1 32877
0 32879 7 1 2 40969 32878
0 32880 5 1 1 32879
0 32881 7 1 2 48085 32880
0 32882 7 1 2 32834 32881
0 32883 5 1 1 32882
0 32884 7 2 2 58039 51559
0 32885 7 1 2 58988 66643
0 32886 5 1 1 32885
0 32887 7 1 2 44221 62259
0 32888 7 1 2 59983 32887
0 32889 5 1 1 32888
0 32890 7 1 2 48985 64431
0 32891 7 1 2 62084 32890
0 32892 5 1 1 32891
0 32893 7 1 2 32889 32892
0 32894 5 1 1 32893
0 32895 7 1 2 40116 32894
0 32896 5 1 1 32895
0 32897 7 1 2 48986 64435
0 32898 5 1 1 32897
0 32899 7 1 2 32896 32898
0 32900 5 1 1 32899
0 32901 7 1 2 44289 32900
0 32902 5 1 1 32901
0 32903 7 1 2 50850 58664
0 32904 7 1 2 64569 32903
0 32905 5 1 1 32904
0 32906 7 1 2 32902 32905
0 32907 5 1 1 32906
0 32908 7 1 2 43030 32907
0 32909 5 1 1 32908
0 32910 7 1 2 32886 32909
0 32911 5 1 1 32910
0 32912 7 1 2 46520 32911
0 32913 5 1 1 32912
0 32914 7 1 2 60248 60515
0 32915 5 1 1 32914
0 32916 7 1 2 32913 32915
0 32917 5 1 1 32916
0 32918 7 1 2 40292 32917
0 32919 5 1 1 32918
0 32920 7 1 2 47494 57962
0 32921 7 1 2 64737 32920
0 32922 5 1 1 32921
0 32923 7 2 2 55108 57391
0 32924 7 1 2 62128 62095
0 32925 7 1 2 67029 32924
0 32926 5 1 1 32925
0 32927 7 1 2 32922 32926
0 32928 5 1 1 32927
0 32929 7 1 2 45343 32928
0 32930 5 1 1 32929
0 32931 7 1 2 32919 32930
0 32932 5 1 1 32931
0 32933 7 1 2 47130 32932
0 32934 5 1 1 32933
0 32935 7 1 2 59850 62246
0 32936 5 1 1 32935
0 32937 7 1 2 47495 67024
0 32938 5 1 1 32937
0 32939 7 1 2 32936 32938
0 32940 5 1 1 32939
0 32941 7 1 2 40293 32940
0 32942 5 1 1 32941
0 32943 7 1 2 62308 63605
0 32944 5 1 1 32943
0 32945 7 1 2 32942 32944
0 32946 5 1 1 32945
0 32947 7 1 2 45344 32946
0 32948 5 1 1 32947
0 32949 7 1 2 54798 61433
0 32950 5 1 1 32949
0 32951 7 1 2 5951 46649
0 32952 5 1 1 32951
0 32953 7 1 2 40117 32952
0 32954 7 1 2 63899 32953
0 32955 5 1 1 32954
0 32956 7 1 2 32950 32955
0 32957 5 1 1 32956
0 32958 7 1 2 62240 32957
0 32959 5 1 1 32958
0 32960 7 1 2 32948 32959
0 32961 5 1 1 32960
0 32962 7 1 2 53926 32961
0 32963 5 1 1 32962
0 32964 7 1 2 40294 46862
0 32965 5 1 1 32964
0 32966 7 1 2 62071 32965
0 32967 5 1 1 32966
0 32968 7 1 2 61582 32967
0 32969 5 1 1 32968
0 32970 7 1 2 32963 32969
0 32971 5 1 1 32970
0 32972 7 1 2 46302 32971
0 32973 5 1 1 32972
0 32974 7 1 2 47819 48987
0 32975 5 1 1 32974
0 32976 7 1 2 41267 48978
0 32977 5 1 1 32976
0 32978 7 1 2 32975 32977
0 32979 5 1 1 32978
0 32980 7 1 2 63558 32979
0 32981 5 1 1 32980
0 32982 7 1 2 48979 65030
0 32983 5 1 1 32982
0 32984 7 1 2 41268 48988
0 32985 5 1 1 32984
0 32986 7 1 2 32983 32985
0 32987 5 1 1 32986
0 32988 7 1 2 45345 61358
0 32989 7 1 2 32987 32988
0 32990 5 1 1 32989
0 32991 7 1 2 32981 32990
0 32992 5 1 1 32991
0 32993 7 1 2 45511 32992
0 32994 5 1 1 32993
0 32995 7 1 2 55109 65862
0 32996 7 1 2 63530 32995
0 32997 5 1 1 32996
0 32998 7 1 2 32994 32997
0 32999 5 1 1 32998
0 33000 7 1 2 43031 32999
0 33001 5 1 1 33000
0 33002 7 1 2 32973 33001
0 33003 7 1 2 32934 33002
0 33004 5 1 1 33003
0 33005 7 1 2 67027 33004
0 33006 5 1 1 33005
0 33007 7 1 2 32883 33006
0 33008 5 1 1 33007
0 33009 7 1 2 64687 33008
0 33010 5 1 1 33009
0 33011 7 1 2 57276 56973
0 33012 7 3 2 62596 33011
0 33013 7 1 2 59310 67031
0 33014 5 1 1 33013
0 33015 7 3 2 45120 63148
0 33016 7 1 2 49375 67034
0 33017 5 1 1 33016
0 33018 7 1 2 55110 58620
0 33019 5 1 1 33018
0 33020 7 1 2 33017 33019
0 33021 5 1 1 33020
0 33022 7 1 2 57215 33021
0 33023 7 1 2 67014 33022
0 33024 5 1 1 33023
0 33025 7 1 2 46637 67032
0 33026 5 1 1 33025
0 33027 7 2 2 55111 49376
0 33028 7 1 2 51857 57383
0 33029 7 1 2 67037 33028
0 33030 5 1 1 33029
0 33031 7 1 2 33026 33030
0 33032 7 1 2 33024 33031
0 33033 5 1 1 33032
0 33034 7 1 2 45199 33033
0 33035 5 1 1 33034
0 33036 7 1 2 33014 33035
0 33037 5 1 1 33036
0 33038 7 1 2 44359 33037
0 33039 5 1 1 33038
0 33040 7 1 2 66447 67033
0 33041 5 1 1 33040
0 33042 7 1 2 33039 33041
0 33043 5 1 1 33042
0 33044 7 1 2 58040 33043
0 33045 5 1 1 33044
0 33046 7 1 2 57216 47949
0 33047 7 1 2 51768 33046
0 33048 7 2 2 66026 66477
0 33049 7 1 2 62180 67039
0 33050 7 1 2 33047 33049
0 33051 5 1 1 33050
0 33052 7 1 2 33045 33051
0 33053 5 1 1 33052
0 33054 7 1 2 50025 33053
0 33055 5 1 1 33054
0 33056 7 1 2 41269 63816
0 33057 5 1 1 33056
0 33058 7 1 2 58905 33057
0 33059 5 1 1 33058
0 33060 7 1 2 58621 33059
0 33061 5 1 1 33060
0 33062 7 1 2 56584 64793
0 33063 5 1 1 33062
0 33064 7 1 2 33061 33063
0 33065 5 1 1 33064
0 33066 7 1 2 41768 33065
0 33067 5 1 1 33066
0 33068 7 1 2 47820 58916
0 33069 5 1 1 33068
0 33070 7 1 2 58906 33069
0 33071 5 1 1 33070
0 33072 7 1 2 14236 6998
0 33073 5 1 1 33072
0 33074 7 1 2 45062 33073
0 33075 7 1 2 33071 33074
0 33076 5 1 1 33075
0 33077 7 1 2 33067 33076
0 33078 5 1 1 33077
0 33079 7 1 2 58609 33078
0 33080 5 1 1 33079
0 33081 7 1 2 60211 59017
0 33082 5 1 1 33081
0 33083 7 1 2 58841 33082
0 33084 5 1 1 33083
0 33085 7 1 2 45121 33084
0 33086 5 1 1 33085
0 33087 7 1 2 66393 33086
0 33088 5 1 1 33087
0 33089 7 1 2 44290 33088
0 33090 5 1 1 33089
0 33091 7 1 2 66395 33090
0 33092 5 1 1 33091
0 33093 7 1 2 47496 33092
0 33094 5 1 1 33093
0 33095 7 1 2 47295 51560
0 33096 7 1 2 62861 33095
0 33097 5 1 1 33096
0 33098 7 1 2 65334 59020
0 33099 5 1 1 33098
0 33100 7 1 2 33097 33099
0 33101 7 1 2 33094 33100
0 33102 5 1 1 33101
0 33103 7 1 2 45512 33102
0 33104 5 1 1 33103
0 33105 7 4 2 63736 59066
0 33106 7 1 2 44222 67041
0 33107 7 1 2 67026 33106
0 33108 5 1 1 33107
0 33109 7 1 2 33104 33108
0 33110 5 1 1 33109
0 33111 7 1 2 46303 33110
0 33112 5 1 1 33111
0 33113 7 1 2 33080 33112
0 33114 5 1 1 33113
0 33115 7 1 2 58041 66608
0 33116 7 1 2 33114 33115
0 33117 5 1 1 33116
0 33118 7 1 2 33055 33117
0 33119 7 1 2 33010 33118
0 33120 5 1 1 33119
0 33121 7 1 2 43773 33120
0 33122 5 1 1 33121
0 33123 7 1 2 65082 66966
0 33124 5 1 1 33123
0 33125 7 1 2 40118 52256
0 33126 7 1 2 52275 33125
0 33127 5 1 1 33126
0 33128 7 1 2 33124 33127
0 33129 5 2 1 33128
0 33130 7 1 2 49358 67045
0 33131 5 1 1 33130
0 33132 7 1 2 59825 59038
0 33133 5 1 1 33132
0 33134 7 1 2 33131 33133
0 33135 5 1 1 33134
0 33136 7 1 2 51561 33135
0 33137 5 1 1 33136
0 33138 7 1 2 47523 66708
0 33139 7 1 2 55375 33138
0 33140 5 1 1 33139
0 33141 7 1 2 33137 33140
0 33142 5 1 1 33141
0 33143 7 1 2 46438 33142
0 33144 5 1 1 33143
0 33145 7 2 2 54004 59992
0 33146 7 1 2 66040 67047
0 33147 5 1 1 33146
0 33148 7 1 2 33144 33147
0 33149 5 1 1 33148
0 33150 7 1 2 45122 33149
0 33151 5 1 1 33150
0 33152 7 1 2 65447 59941
0 33153 7 1 2 56760 33152
0 33154 5 1 1 33153
0 33155 7 1 2 33151 33154
0 33156 5 1 1 33155
0 33157 7 1 2 59543 33156
0 33158 5 1 1 33157
0 33159 7 1 2 41850 64538
0 33160 7 1 2 62722 33159
0 33161 5 1 1 33160
0 33162 7 1 2 44291 33161
0 33163 7 1 2 33158 33162
0 33164 5 1 1 33163
0 33165 7 1 2 65436 59610
0 33166 5 1 1 33165
0 33167 7 1 2 46521 26792
0 33168 5 1 1 33167
0 33169 7 1 2 45123 59744
0 33170 7 1 2 33168 33169
0 33171 7 1 2 56761 33170
0 33172 5 1 1 33171
0 33173 7 1 2 33166 33172
0 33174 5 1 1 33173
0 33175 7 1 2 54985 33174
0 33176 5 1 1 33175
0 33177 7 1 2 41033 33176
0 33178 5 1 1 33177
0 33179 7 1 2 44360 33178
0 33180 7 1 2 33164 33179
0 33181 5 1 1 33180
0 33182 7 1 2 46548 64539
0 33183 7 1 2 66360 33182
0 33184 5 1 1 33183
0 33185 7 1 2 33181 33184
0 33186 5 1 1 33185
0 33187 7 1 2 65092 33186
0 33188 5 1 1 33187
0 33189 7 1 2 43774 52089
0 33190 5 1 1 33189
0 33191 7 1 2 42181 33190
0 33192 5 1 1 33191
0 33193 7 2 2 46968 33192
0 33194 5 1 1 67049
0 33195 7 2 2 45513 52428
0 33196 5 1 1 67051
0 33197 7 1 2 67050 33196
0 33198 5 1 1 33197
0 33199 7 1 2 33198 63299
0 33200 5 1 1 33199
0 33201 7 1 2 64889 66726
0 33202 5 2 1 33201
0 33203 7 1 2 67053 63305
0 33204 5 1 1 33203
0 33205 7 1 2 33200 33204
0 33206 5 1 1 33205
0 33207 7 1 2 43148 33206
0 33208 5 1 1 33207
0 33209 7 2 2 53660 64992
0 33210 7 1 2 67042 67055
0 33211 5 1 1 33210
0 33212 7 1 2 33208 33211
0 33213 5 1 1 33212
0 33214 7 1 2 46591 33213
0 33215 5 1 1 33214
0 33216 7 1 2 61434 67054
0 33217 5 1 1 33216
0 33218 7 1 2 52552 60522
0 33219 5 1 1 33218
0 33220 7 1 2 64896 33219
0 33221 5 3 1 33220
0 33222 7 1 2 41992 59146
0 33223 7 1 2 67057 33222
0 33224 5 1 1 33223
0 33225 7 1 2 33217 33224
0 33226 5 1 1 33225
0 33227 7 1 2 59396 33226
0 33228 5 1 1 33227
0 33229 7 1 2 59412 67056
0 33230 5 1 1 33229
0 33231 7 1 2 33228 33230
0 33232 5 1 1 33231
0 33233 7 1 2 64688 33232
0 33234 5 1 1 33233
0 33235 7 1 2 33215 33234
0 33236 5 1 1 33235
0 33237 7 1 2 43263 33236
0 33238 5 1 1 33237
0 33239 7 3 2 59544 64049
0 33240 7 1 2 51369 57825
0 33241 7 1 2 63333 33240
0 33242 5 1 1 33241
0 33243 7 1 2 58899 50907
0 33244 5 1 1 33243
0 33245 7 1 2 59058 50881
0 33246 7 1 2 62785 33245
0 33247 5 1 1 33246
0 33248 7 1 2 33244 33247
0 33249 5 1 1 33248
0 33250 7 1 2 43593 57505
0 33251 7 1 2 33249 33250
0 33252 5 1 1 33251
0 33253 7 1 2 33242 33252
0 33254 5 1 1 33253
0 33255 7 1 2 67060 33254
0 33256 5 1 1 33255
0 33257 7 1 2 33238 33256
0 33258 5 1 1 33257
0 33259 7 1 2 49064 33258
0 33260 5 1 1 33259
0 33261 7 1 2 51129 63505
0 33262 5 2 1 33261
0 33263 7 1 2 64017 67063
0 33264 5 1 1 33263
0 33265 7 1 2 40295 55376
0 33266 5 1 1 33265
0 33267 7 1 2 61965 48363
0 33268 5 1 1 33267
0 33269 7 1 2 51562 59881
0 33270 5 1 1 33269
0 33271 7 1 2 33268 33270
0 33272 5 1 1 33271
0 33273 7 1 2 47497 33272
0 33274 5 1 1 33273
0 33275 7 1 2 33266 33274
0 33276 7 1 2 33264 33275
0 33277 5 1 1 33276
0 33278 7 1 2 42182 33277
0 33279 5 1 1 33278
0 33280 7 1 2 47296 59993
0 33281 5 1 1 33280
0 33282 7 1 2 65448 57428
0 33283 5 1 1 33282
0 33284 7 1 2 33281 33283
0 33285 5 1 1 33284
0 33286 7 1 2 41993 33285
0 33287 5 1 1 33286
0 33288 7 1 2 54720 57429
0 33289 5 1 1 33288
0 33290 7 1 2 59998 33289
0 33291 5 1 1 33290
0 33292 7 1 2 67052 33291
0 33293 5 1 1 33292
0 33294 7 2 2 48403 61390
0 33295 5 1 1 67065
0 33296 7 1 2 46304 62199
0 33297 5 1 1 33296
0 33298 7 1 2 33295 33297
0 33299 5 1 1 33298
0 33300 7 1 2 40498 33299
0 33301 5 1 1 33300
0 33302 7 1 2 33293 33301
0 33303 7 1 2 33287 33302
0 33304 7 1 2 33279 33303
0 33305 5 2 1 33304
0 33306 7 1 2 66694 67067
0 33307 5 1 1 33306
0 33308 7 2 2 51563 48328
0 33309 5 1 1 67069
0 33310 7 1 2 67058 67070
0 33311 5 1 1 33310
0 33312 7 1 2 64993 55377
0 33313 5 1 1 33312
0 33314 7 1 2 33311 33313
0 33315 5 2 1 33314
0 33316 7 1 2 66706 67071
0 33317 5 1 1 33316
0 33318 7 1 2 33307 33317
0 33319 5 1 1 33318
0 33320 7 1 2 43264 33319
0 33321 5 1 1 33320
0 33322 7 1 2 65467 55378
0 33323 5 1 1 33322
0 33324 7 2 2 43446 63165
0 33325 7 1 2 55573 60050
0 33326 7 1 2 67073 33325
0 33327 5 1 1 33326
0 33328 7 1 2 33323 33327
0 33329 5 1 1 33328
0 33330 7 1 2 63582 67061
0 33331 7 1 2 33329 33330
0 33332 5 1 1 33331
0 33333 7 1 2 33321 33332
0 33334 5 1 1 33333
0 33335 7 1 2 55112 33334
0 33336 5 1 1 33335
0 33337 7 1 2 54005 67068
0 33338 5 1 1 33337
0 33339 7 1 2 54183 67072
0 33340 5 1 1 33339
0 33341 7 1 2 33338 33340
0 33342 5 1 1 33341
0 33343 7 1 2 66340 33342
0 33344 5 1 1 33343
0 33345 7 1 2 60590 63369
0 33346 7 1 2 63143 33345
0 33347 5 1 1 33346
0 33348 7 1 2 54006 50904
0 33349 5 1 1 33348
0 33350 7 1 2 62169 33349
0 33351 5 1 1 33350
0 33352 7 1 2 48404 47950
0 33353 7 1 2 33351 33352
0 33354 5 1 1 33353
0 33355 7 1 2 33347 33354
0 33356 5 1 1 33355
0 33357 7 1 2 43447 33356
0 33358 5 1 1 33357
0 33359 7 1 2 56845 58927
0 33360 7 1 2 48405 33359
0 33361 7 1 2 58520 33360
0 33362 5 1 1 33361
0 33363 7 1 2 33358 33362
0 33364 5 1 1 33363
0 33365 7 1 2 40499 65106
0 33366 7 1 2 33364 33365
0 33367 5 1 1 33366
0 33368 7 1 2 33344 33367
0 33369 7 1 2 33336 33368
0 33370 7 1 2 33260 33369
0 33371 7 1 2 33188 33370
0 33372 5 1 1 33371
0 33373 7 1 2 58042 33372
0 33374 5 1 1 33373
0 33375 7 1 2 33122 33374
0 33376 5 1 1 33375
0 33377 7 1 2 67009 33376
0 33378 5 1 1 33377
0 33379 7 3 2 47561 63780
0 33380 7 3 2 45514 67075
0 33381 7 2 2 52235 67078
0 33382 7 1 2 57164 67081
0 33383 5 1 1 33382
0 33384 7 2 2 53842 63539
0 33385 7 2 2 65058 67083
0 33386 7 1 2 48605 56976
0 33387 7 1 2 67085 33386
0 33388 5 1 1 33387
0 33389 7 1 2 33383 33388
0 33390 5 1 1 33389
0 33391 7 1 2 55113 33390
0 33392 5 1 1 33391
0 33393 7 2 2 67079 64711
0 33394 7 2 2 61526 63130
0 33395 7 1 2 67087 67089
0 33396 5 1 1 33395
0 33397 7 1 2 63342 55183
0 33398 7 1 2 67086 33397
0 33399 5 1 1 33398
0 33400 7 1 2 33396 33399
0 33401 7 1 2 33392 33400
0 33402 5 1 1 33401
0 33403 7 1 2 43960 33402
0 33404 5 1 1 33403
0 33405 7 3 2 44825 51460
0 33406 7 1 2 58674 67091
0 33407 7 1 2 67088 33406
0 33408 5 1 1 33407
0 33409 7 1 2 58012 67038
0 33410 7 1 2 67082 33409
0 33411 5 1 1 33410
0 33412 7 1 2 33408 33411
0 33413 7 1 2 33404 33412
0 33414 5 1 1 33413
0 33415 7 1 2 45200 33414
0 33416 5 1 1 33415
0 33417 7 2 2 58043 67080
0 33418 7 1 2 66373 67094
0 33419 5 1 1 33418
0 33420 7 1 2 33416 33419
0 33421 5 1 1 33420
0 33422 7 1 2 44361 33421
0 33423 5 1 1 33422
0 33424 7 1 2 41534 66948
0 33425 7 1 2 67076 33424
0 33426 5 1 1 33425
0 33427 7 1 2 41270 65053
0 33428 5 1 1 33427
0 33429 7 1 2 23405 33428
0 33430 5 1 1 33429
0 33431 7 1 2 64689 62612
0 33432 7 1 2 67084 33431
0 33433 7 1 2 33430 33432
0 33434 5 1 1 33433
0 33435 7 1 2 33426 33434
0 33436 5 1 1 33435
0 33437 7 1 2 43961 33436
0 33438 5 1 1 33437
0 33439 7 1 2 46592 53267
0 33440 7 1 2 662 33439
0 33441 7 1 2 63782 33440
0 33442 5 1 1 33441
0 33443 7 1 2 33438 33442
0 33444 5 1 1 33443
0 33445 7 1 2 57663 33444
0 33446 5 1 1 33445
0 33447 7 1 2 65312 67028
0 33448 7 1 2 67077 33447
0 33449 5 1 1 33448
0 33450 7 1 2 33446 33449
0 33451 5 1 1 33450
0 33452 7 1 2 45515 33451
0 33453 5 1 1 33452
0 33454 7 1 2 54624 55768
0 33455 7 1 2 66646 33454
0 33456 7 2 2 53843 50738
0 33457 5 1 1 67096
0 33458 7 1 2 66571 67097
0 33459 7 1 2 33455 33458
0 33460 7 1 2 65250 33459
0 33461 5 1 1 33460
0 33462 7 1 2 33453 33461
0 33463 5 1 1 33462
0 33464 7 1 2 49065 33463
0 33465 5 1 1 33464
0 33466 7 1 2 56748 66448
0 33467 7 1 2 67095 33466
0 33468 5 1 1 33467
0 33469 7 1 2 33465 33468
0 33470 7 1 2 33423 33469
0 33471 5 1 1 33470
0 33472 7 1 2 45787 33471
0 33473 5 1 1 33472
0 33474 7 1 2 58044 64690
0 33475 7 1 2 56013 63540
0 33476 7 1 2 33474 33475
0 33477 7 1 2 66712 33476
0 33478 7 1 2 59021 33477
0 33479 5 1 1 33478
0 33480 7 1 2 33473 33479
0 33481 5 1 1 33480
0 33482 7 1 2 65061 33481
0 33483 5 1 1 33482
0 33484 7 1 2 59719 64899
0 33485 5 1 1 33484
0 33486 7 1 2 65241 33485
0 33487 5 1 1 33486
0 33488 7 1 2 45516 33487
0 33489 5 1 1 33488
0 33490 7 1 2 65247 33489
0 33491 5 1 1 33490
0 33492 7 1 2 63583 33491
0 33493 5 1 1 33492
0 33494 7 1 2 64837 66677
0 33495 5 1 1 33494
0 33496 7 1 2 33493 33495
0 33497 5 1 1 33496
0 33498 7 3 2 50811 57430
0 33499 7 1 2 33497 67098
0 33500 5 1 1 33499
0 33501 7 1 2 58045 61064
0 33502 5 1 1 33501
0 33503 7 1 2 49613 65479
0 33504 5 1 1 33503
0 33505 7 1 2 33502 33504
0 33506 5 1 1 33505
0 33507 7 1 2 61747 33506
0 33508 5 1 1 33507
0 33509 7 1 2 47537 47568
0 33510 7 1 2 3664 33509
0 33511 5 1 1 33510
0 33512 7 1 2 54763 63512
0 33513 7 1 2 33511 33512
0 33514 5 1 1 33513
0 33515 7 1 2 33508 33514
0 33516 5 1 1 33515
0 33517 7 1 2 46168 33516
0 33518 5 1 1 33517
0 33519 7 1 2 40296 56197
0 33520 5 1 1 33519
0 33521 7 1 2 65129 33520
0 33522 5 2 1 33521
0 33523 7 1 2 61748 67101
0 33524 5 1 1 33523
0 33525 7 2 2 60638 62697
0 33526 5 1 1 67103
0 33527 7 1 2 52815 67104
0 33528 5 1 1 33527
0 33529 7 1 2 33524 33528
0 33530 5 1 1 33529
0 33531 7 1 2 56863 33530
0 33532 5 1 1 33531
0 33533 7 1 2 33518 33532
0 33534 5 1 1 33533
0 33535 7 1 2 43775 33534
0 33536 5 1 1 33535
0 33537 7 1 2 66713 61749
0 33538 5 1 1 33537
0 33539 7 1 2 62650 61674
0 33540 5 1 1 33539
0 33541 7 1 2 33538 33540
0 33542 5 1 1 33541
0 33543 7 1 2 40500 33542
0 33544 5 1 1 33543
0 33545 7 1 2 28427 61675
0 33546 5 1 1 33545
0 33547 7 1 2 33544 33546
0 33548 5 1 1 33547
0 33549 7 1 2 56864 33548
0 33550 5 1 1 33549
0 33551 7 1 2 61676 67059
0 33552 5 1 1 33551
0 33553 7 2 2 65064 62678
0 33554 7 1 2 56892 63381
0 33555 7 1 2 67105 33554
0 33556 5 1 1 33555
0 33557 7 1 2 33552 33556
0 33558 5 1 1 33557
0 33559 7 1 2 41994 33558
0 33560 5 1 1 33559
0 33561 7 1 2 65075 66905
0 33562 5 1 1 33561
0 33563 7 1 2 33560 33562
0 33564 5 1 1 33563
0 33565 7 1 2 50812 33564
0 33566 5 1 1 33565
0 33567 7 1 2 33550 33566
0 33568 7 1 2 33536 33567
0 33569 5 1 1 33568
0 33570 7 1 2 45201 33569
0 33571 5 1 1 33570
0 33572 7 1 2 52693 50547
0 33573 5 1 1 33572
0 33574 7 1 2 56992 33194
0 33575 5 1 1 33574
0 33576 7 2 2 33573 33575
0 33577 5 1 1 67107
0 33578 7 1 2 48525 51338
0 33579 7 1 2 14034 33578
0 33580 5 1 1 33579
0 33581 7 1 2 67108 33580
0 33582 5 1 1 33581
0 33583 7 1 2 66919 33582
0 33584 5 1 1 33583
0 33585 7 1 2 33571 33584
0 33586 5 1 1 33585
0 33587 7 1 2 55379 33586
0 33588 5 1 1 33587
0 33589 7 1 2 33500 33588
0 33590 5 1 1 33589
0 33591 7 1 2 44362 33590
0 33592 5 1 1 33591
0 33593 7 1 2 55380 33577
0 33594 5 1 1 33593
0 33595 7 1 2 65245 67099
0 33596 5 1 1 33595
0 33597 7 1 2 56865 55381
0 33598 5 2 1 33597
0 33599 7 1 2 65652 54481
0 33600 7 1 2 66907 33599
0 33601 5 1 1 33600
0 33602 7 1 2 67109 33601
0 33603 5 1 1 33602
0 33604 7 1 2 43448 33603
0 33605 5 1 1 33604
0 33606 7 1 2 40297 49309
0 33607 5 2 1 33606
0 33608 7 1 2 66913 67111
0 33609 5 1 1 33608
0 33610 7 1 2 52818 62700
0 33611 5 1 1 33610
0 33612 7 1 2 33609 33611
0 33613 7 1 2 33605 33612
0 33614 5 1 1 33613
0 33615 7 1 2 45517 33614
0 33616 5 1 1 33615
0 33617 7 1 2 33596 33616
0 33618 7 1 2 33594 33617
0 33619 5 1 1 33618
0 33620 7 1 2 66690 33619
0 33621 5 1 1 33620
0 33622 7 1 2 33592 33621
0 33623 5 1 1 33622
0 33624 7 1 2 55114 33623
0 33625 5 1 1 33624
0 33626 7 2 2 62522 61134
0 33627 7 2 2 59545 53141
0 33628 7 1 2 67113 67115
0 33629 5 1 1 33628
0 33630 7 1 2 56866 59720
0 33631 5 1 1 33630
0 33632 7 1 2 33629 33631
0 33633 5 1 1 33632
0 33634 7 1 2 59093 33633
0 33635 5 1 1 33634
0 33636 7 1 2 59963 53142
0 33637 7 1 2 67114 33636
0 33638 5 1 1 33637
0 33639 7 1 2 63956 66697
0 33640 7 1 2 56993 33639
0 33641 5 1 1 33640
0 33642 7 1 2 33638 33641
0 33643 5 1 1 33642
0 33644 7 1 2 59546 33643
0 33645 5 1 1 33644
0 33646 7 1 2 59634 62755
0 33647 7 1 2 62337 33646
0 33648 5 1 1 33647
0 33649 7 1 2 33645 33648
0 33650 5 1 1 33649
0 33651 7 1 2 44292 33650
0 33652 5 1 1 33651
0 33653 7 1 2 33635 33652
0 33654 5 1 1 33653
0 33655 7 1 2 55382 33654
0 33656 5 1 1 33655
0 33657 7 2 2 46522 66007
0 33658 7 1 2 66908 59071
0 33659 7 1 2 67117 33658
0 33660 7 1 2 67046 33659
0 33661 5 1 1 33660
0 33662 7 1 2 33656 33661
0 33663 5 1 1 33662
0 33664 7 1 2 48942 33663
0 33665 5 1 1 33664
0 33666 7 1 2 56867 65797
0 33667 5 1 1 33666
0 33668 7 1 2 63343 66378
0 33669 7 1 2 67116 33668
0 33670 5 1 1 33669
0 33671 7 1 2 33667 33670
0 33672 5 1 1 33671
0 33673 7 1 2 67048 33672
0 33674 5 1 1 33673
0 33675 7 1 2 33665 33674
0 33676 5 1 1 33675
0 33677 7 1 2 44363 33676
0 33678 5 1 1 33677
0 33679 7 1 2 41679 46549
0 33680 7 1 2 51474 33679
0 33681 7 1 2 64562 33680
0 33682 7 1 2 62808 33681
0 33683 5 1 1 33682
0 33684 7 1 2 33678 33683
0 33685 5 1 1 33684
0 33686 7 1 2 65093 33685
0 33687 5 1 1 33686
0 33688 7 1 2 65220 28496
0 33689 5 1 1 33688
0 33690 7 1 2 54007 64909
0 33691 5 1 1 33690
0 33692 7 1 2 48943 66234
0 33693 5 1 1 33692
0 33694 7 1 2 33691 33693
0 33695 5 1 1 33694
0 33696 7 1 2 33689 33695
0 33697 5 1 1 33696
0 33698 7 1 2 57069 65492
0 33699 7 1 2 61370 33698
0 33700 7 1 2 65499 33699
0 33701 5 1 1 33700
0 33702 7 1 2 33697 33701
0 33703 5 1 1 33702
0 33704 7 1 2 67100 33703
0 33705 5 1 1 33704
0 33706 7 1 2 63996 67106
0 33707 5 1 1 33706
0 33708 7 1 2 54101 65501
0 33709 5 1 1 33708
0 33710 7 1 2 33707 33709
0 33711 5 1 1 33710
0 33712 7 1 2 56994 33711
0 33713 5 1 1 33712
0 33714 7 1 2 65735 50949
0 33715 7 1 2 63963 33714
0 33716 5 1 1 33715
0 33717 7 1 2 58046 52694
0 33718 7 1 2 66837 33717
0 33719 7 1 2 62470 33718
0 33720 5 1 1 33719
0 33721 7 1 2 33716 33720
0 33722 5 1 1 33721
0 33723 7 1 2 44548 33722
0 33724 5 1 1 33723
0 33725 7 1 2 33713 33724
0 33726 5 1 1 33725
0 33727 7 1 2 41995 33726
0 33728 5 1 1 33727
0 33729 7 1 2 43776 67102
0 33730 5 1 1 33729
0 33731 7 1 2 65522 33730
0 33732 5 1 1 33731
0 33733 7 1 2 56995 33732
0 33734 5 1 1 33733
0 33735 7 1 2 50459 49694
0 33736 5 1 1 33735
0 33737 7 1 2 52965 66210
0 33738 7 1 2 33736 33737
0 33739 5 1 1 33738
0 33740 7 1 2 33734 33739
0 33741 5 1 1 33740
0 33742 7 1 2 54008 33741
0 33743 5 1 1 33742
0 33744 7 1 2 33728 33743
0 33745 5 1 1 33744
0 33746 7 1 2 65107 33745
0 33747 5 1 1 33746
0 33748 7 1 2 54102 64900
0 33749 5 1 1 33748
0 33750 7 1 2 54009 67112
0 33751 5 1 1 33750
0 33752 7 1 2 45518 33751
0 33753 7 1 2 33749 33752
0 33754 7 1 2 61103 33753
0 33755 5 1 1 33754
0 33756 7 1 2 54184 67064
0 33757 5 1 1 33756
0 33758 7 2 2 47821 54103
0 33759 5 1 1 67119
0 33760 7 1 2 62005 33759
0 33761 5 1 1 33760
0 33762 7 1 2 47498 33761
0 33763 5 1 1 33762
0 33764 7 1 2 42183 62316
0 33765 7 1 2 33763 33764
0 33766 7 1 2 33757 33765
0 33767 5 1 1 33766
0 33768 7 1 2 33755 33767
0 33769 5 1 1 33768
0 33770 7 1 2 47297 57070
0 33771 5 1 1 33770
0 33772 7 1 2 54104 65449
0 33773 5 1 1 33772
0 33774 7 1 2 33771 33773
0 33775 5 1 1 33774
0 33776 7 1 2 41996 33775
0 33777 5 1 1 33776
0 33778 7 2 2 54081 59257
0 33779 5 1 1 67121
0 33780 7 1 2 60619 33779
0 33781 5 1 1 33780
0 33782 7 1 2 40501 33781
0 33783 5 1 1 33782
0 33784 7 1 2 33777 33783
0 33785 7 1 2 33769 33784
0 33786 5 1 1 33785
0 33787 7 1 2 56868 33786
0 33788 5 1 1 33787
0 33789 7 1 2 22859 30456
0 33790 5 1 1 33789
0 33791 7 1 2 54185 33790
0 33792 5 1 1 33791
0 33793 7 1 2 60620 33792
0 33794 5 1 1 33793
0 33795 7 1 2 47822 33794
0 33796 5 1 1 33795
0 33797 7 1 2 64823 62475
0 33798 5 1 1 33797
0 33799 7 1 2 54010 59783
0 33800 5 1 1 33799
0 33801 7 1 2 60621 12190
0 33802 5 1 1 33801
0 33803 7 1 2 40502 33802
0 33804 5 1 1 33803
0 33805 7 1 2 33800 33804
0 33806 7 1 2 33798 33805
0 33807 7 1 2 33796 33806
0 33808 5 1 1 33807
0 33809 7 1 2 50813 33808
0 33810 5 1 1 33809
0 33811 7 1 2 33788 33810
0 33812 5 1 1 33811
0 33813 7 1 2 66341 33812
0 33814 5 1 1 33813
0 33815 7 1 2 33747 33814
0 33816 5 1 1 33815
0 33817 7 1 2 55383 33816
0 33818 5 1 1 33817
0 33819 7 1 2 33705 33818
0 33820 7 1 2 33687 33819
0 33821 7 1 2 33625 33820
0 33822 5 1 1 33821
0 33823 7 1 2 53781 33822
0 33824 5 1 1 33823
0 33825 7 1 2 33483 33824
0 33826 7 1 2 33378 33825
0 33827 7 1 2 32739 33826
0 33828 7 1 2 32321 33827
0 33829 7 1 2 31117 33828
0 33830 7 1 2 29974 33829
0 33831 7 2 2 43032 66609
0 33832 7 2 2 55260 67123
0 33833 7 1 2 67125 64465
0 33834 5 1 1 33833
0 33835 7 4 2 51370 59547
0 33836 7 1 2 49614 52954
0 33837 5 1 1 33836
0 33838 7 1 2 19545 33837
0 33839 5 1 1 33838
0 33840 7 1 2 67127 33839
0 33841 5 1 1 33840
0 33842 7 1 2 65136 56437
0 33843 5 1 1 33842
0 33844 7 1 2 33841 33843
0 33845 5 1 1 33844
0 33846 7 1 2 44364 33845
0 33847 5 1 1 33846
0 33848 7 2 2 46550 62241
0 33849 5 1 1 67131
0 33850 7 1 2 56438 67132
0 33851 5 1 1 33850
0 33852 7 1 2 33847 33851
0 33853 5 1 1 33852
0 33854 7 1 2 42712 50346
0 33855 7 1 2 33853 33854
0 33856 5 1 1 33855
0 33857 7 1 2 33834 33856
0 33858 5 1 1 33857
0 33859 7 1 2 44704 33858
0 33860 5 1 1 33859
0 33861 7 1 2 63444 55440
0 33862 7 1 2 67126 33861
0 33863 5 1 1 33862
0 33864 7 1 2 33860 33863
0 33865 5 1 1 33864
0 33866 7 1 2 40885 33865
0 33867 5 1 1 33866
0 33868 7 2 2 63085 63567
0 33869 7 1 2 59572 67133
0 33870 5 1 1 33869
0 33871 7 1 2 58181 48304
0 33872 5 1 1 33871
0 33873 7 5 2 45519 46305
0 33874 7 1 2 58831 67135
0 33875 5 1 1 33874
0 33876 7 1 2 33872 33875
0 33877 5 1 1 33876
0 33878 7 1 2 66717 33877
0 33879 5 1 1 33878
0 33880 7 1 2 33870 33879
0 33881 5 1 1 33880
0 33882 7 1 2 44705 33881
0 33883 5 1 1 33882
0 33884 7 2 2 45520 65391
0 33885 7 1 2 67140 67134
0 33886 5 1 1 33885
0 33887 7 1 2 33883 33886
0 33888 5 1 1 33887
0 33889 7 1 2 44365 33888
0 33890 5 1 1 33889
0 33891 7 2 2 46551 63078
0 33892 7 1 2 67142 59155
0 33893 7 1 2 66054 33892
0 33894 5 1 1 33893
0 33895 7 1 2 33890 33894
0 33896 5 1 1 33895
0 33897 7 1 2 58047 33896
0 33898 5 1 1 33897
0 33899 7 2 2 44366 65147
0 33900 7 1 2 59804 54223
0 33901 7 1 2 62463 33900
0 33902 7 1 2 67144 33901
0 33903 7 1 2 65776 33902
0 33904 5 1 1 33903
0 33905 7 1 2 33898 33904
0 33906 7 1 2 33867 33905
0 33907 5 1 1 33906
0 33908 7 1 2 44549 33907
0 33909 5 1 1 33908
0 33910 7 1 2 65920 53334
0 33911 7 1 2 55986 33910
0 33912 7 1 2 67124 33911
0 33913 5 1 1 33912
0 33914 7 1 2 33909 33913
0 33915 5 1 1 33914
0 33916 7 1 2 48944 33915
0 33917 5 1 1 33916
0 33918 7 1 2 49615 49453
0 33919 7 1 2 65383 65425
0 33920 7 1 2 33918 33919
0 33921 7 1 2 55184 33920
0 33922 7 1 2 66789 33921
0 33923 5 1 1 33922
0 33924 7 1 2 33917 33923
0 33925 5 1 1 33924
0 33926 7 1 2 55115 33925
0 33927 5 1 1 33926
0 33928 7 1 2 66055 66342
0 33929 5 1 1 33928
0 33930 7 1 2 46523 49454
0 33931 7 1 2 67040 33930
0 33932 7 1 2 58182 33931
0 33933 5 1 1 33932
0 33934 7 1 2 33929 33933
0 33935 5 1 1 33934
0 33936 7 1 2 58048 33935
0 33937 5 1 1 33936
0 33938 7 1 2 40679 67128
0 33939 5 1 1 33938
0 33940 7 1 2 65138 33939
0 33941 5 1 1 33940
0 33942 7 1 2 44367 33941
0 33943 5 1 1 33942
0 33944 7 1 2 33849 33943
0 33945 5 1 1 33944
0 33946 7 1 2 57664 33945
0 33947 5 1 1 33946
0 33948 7 1 2 62242 65313
0 33949 5 1 1 33948
0 33950 7 1 2 33947 33949
0 33951 5 1 1 33950
0 33952 7 1 2 62496 58785
0 33953 7 1 2 33951 33952
0 33954 5 1 1 33953
0 33955 7 1 2 33937 33954
0 33956 5 1 1 33955
0 33957 7 1 2 46169 33956
0 33958 5 1 1 33957
0 33959 7 3 2 48526 55261
0 33960 7 1 2 53708 67146
0 33961 7 1 2 66343 33960
0 33962 5 1 1 33961
0 33963 7 1 2 33958 33962
0 33964 5 1 1 33963
0 33965 7 1 2 44550 33964
0 33966 5 1 1 33965
0 33967 7 1 2 65921 60987
0 33968 7 1 2 66344 33967
0 33969 5 1 1 33968
0 33970 7 1 2 33966 33969
0 33971 5 1 1 33970
0 33972 7 1 2 56569 33971
0 33973 5 1 1 33972
0 33974 7 1 2 44972 59512
0 33975 7 1 2 52887 33974
0 33976 7 1 2 63226 33975
0 33977 7 1 2 66524 33976
0 33978 7 1 2 65325 33977
0 33979 5 1 1 33978
0 33980 7 1 2 33973 33979
0 33981 5 1 1 33980
0 33982 7 1 2 43033 33981
0 33983 5 1 1 33982
0 33984 7 1 2 49250 58183
0 33985 5 1 1 33984
0 33986 7 1 2 45521 58832
0 33987 5 1 1 33986
0 33988 7 1 2 33985 33987
0 33989 5 1 1 33988
0 33990 7 1 2 58049 33989
0 33991 5 1 1 33990
0 33992 7 1 2 42880 57719
0 33993 5 1 1 33992
0 33994 7 1 2 50814 48443
0 33995 5 1 1 33994
0 33996 7 1 2 33993 33995
0 33997 5 1 1 33996
0 33998 7 1 2 51371 54536
0 33999 7 1 2 33997 33998
0 34000 5 1 1 33999
0 34001 7 1 2 33991 34000
0 34002 5 1 1 34001
0 34003 7 1 2 46984 66615
0 34004 7 1 2 58989 34003
0 34005 7 1 2 67118 34004
0 34006 7 1 2 34002 34005
0 34007 5 1 1 34006
0 34008 7 1 2 43149 34007
0 34009 7 1 2 33983 34008
0 34010 7 1 2 33927 34009
0 34011 5 1 1 34010
0 34012 7 1 2 54298 54518
0 34013 5 9 1 34012
0 34014 7 1 2 48711 67149
0 34015 5 1 1 34014
0 34016 7 1 2 53217 52241
0 34017 5 1 1 34016
0 34018 7 2 2 42713 59584
0 34019 7 1 2 41535 67158
0 34020 5 1 1 34019
0 34021 7 1 2 34017 34020
0 34022 5 1 1 34021
0 34023 7 1 2 40886 34022
0 34024 5 1 1 34023
0 34025 7 1 2 34015 34024
0 34026 5 1 1 34025
0 34027 7 1 2 43962 34026
0 34028 5 1 1 34027
0 34029 7 1 2 67092 67159
0 34030 5 1 1 34029
0 34031 7 1 2 34028 34030
0 34032 5 1 1 34031
0 34033 7 1 2 48131 34032
0 34034 5 1 1 34033
0 34035 7 1 2 52242 48295
0 34036 7 1 2 66203 34035
0 34037 5 1 1 34036
0 34038 7 1 2 34034 34037
0 34039 5 1 1 34038
0 34040 7 1 2 45788 34039
0 34041 5 1 1 34040
0 34042 7 1 2 65542 64530
0 34043 5 1 1 34042
0 34044 7 1 2 53506 55202
0 34045 5 1 1 34044
0 34046 7 1 2 34043 34045
0 34047 5 1 1 34046
0 34048 7 1 2 66189 34047
0 34049 5 1 1 34048
0 34050 7 1 2 34041 34049
0 34051 5 1 1 34050
0 34052 7 1 2 41680 34051
0 34053 5 1 1 34052
0 34054 7 1 2 62227 56962
0 34055 5 1 1 34054
0 34056 7 1 2 52385 51346
0 34057 7 1 2 56509 34056
0 34058 5 1 1 34057
0 34059 7 1 2 34055 34058
0 34060 5 1 1 34059
0 34061 7 1 2 52360 51275
0 34062 7 1 2 34060 34061
0 34063 5 1 1 34062
0 34064 7 1 2 34053 34063
0 34065 5 1 1 34064
0 34066 7 1 2 65361 34065
0 34067 5 1 1 34066
0 34068 7 1 2 46306 49791
0 34069 7 1 2 52201 34068
0 34070 7 1 2 64738 34069
0 34071 5 1 1 34070
0 34072 7 1 2 64386 50799
0 34073 7 1 2 64552 34072
0 34074 7 1 2 66430 34073
0 34075 5 1 1 34074
0 34076 7 1 2 34071 34075
0 34077 5 1 1 34076
0 34078 7 1 2 40503 34077
0 34079 5 1 1 34078
0 34080 7 1 2 1771 52361
0 34081 7 2 2 52306 34080
0 34082 5 1 1 67160
0 34083 7 1 2 51276 67161
0 34084 7 1 2 64739 34083
0 34085 5 1 1 34084
0 34086 7 1 2 34079 34085
0 34087 5 1 1 34086
0 34088 7 1 2 45202 34087
0 34089 5 1 1 34088
0 34090 7 3 2 40504 48839
0 34091 5 1 1 67162
0 34092 7 1 2 44826 67163
0 34093 5 1 1 34092
0 34094 7 1 2 34082 34093
0 34095 5 1 1 34094
0 34096 7 2 2 62769 34095
0 34097 7 1 2 59008 66976
0 34098 7 1 2 67165 34097
0 34099 5 1 1 34098
0 34100 7 1 2 34089 34099
0 34101 5 1 1 34100
0 34102 7 1 2 44368 34101
0 34103 5 1 1 34102
0 34104 7 1 2 44973 65352
0 34105 7 1 2 67166 34104
0 34106 5 1 1 34105
0 34107 7 1 2 34103 34106
0 34108 5 1 1 34107
0 34109 7 1 2 65930 34108
0 34110 5 1 1 34109
0 34111 7 1 2 52386 50137
0 34112 5 2 1 34111
0 34113 7 1 2 41536 53245
0 34114 5 1 1 34113
0 34115 7 1 2 67167 34114
0 34116 5 1 1 34115
0 34117 7 1 2 55353 34116
0 34118 5 1 1 34117
0 34119 7 1 2 44827 50096
0 34120 7 1 2 53749 34119
0 34121 5 1 1 34120
0 34122 7 1 2 34118 34121
0 34123 5 1 1 34122
0 34124 7 1 2 52362 62770
0 34125 7 1 2 34123 34124
0 34126 7 1 2 65356 34125
0 34127 5 1 1 34126
0 34128 7 1 2 34110 34127
0 34129 5 1 1 34128
0 34130 7 1 2 60680 34129
0 34131 5 1 1 34130
0 34132 7 1 2 56120 61249
0 34133 7 1 2 63086 62338
0 34134 7 1 2 34132 34133
0 34135 5 1 1 34134
0 34136 7 1 2 57665 50597
0 34137 7 1 2 58050 34136
0 34138 7 1 2 65772 65062
0 34139 7 1 2 34137 34138
0 34140 5 1 1 34139
0 34141 7 1 2 34135 34140
0 34142 5 1 1 34141
0 34143 7 1 2 48945 34142
0 34144 5 1 1 34143
0 34145 7 1 2 65762 54042
0 34146 7 1 2 63829 34145
0 34147 7 1 2 66962 34146
0 34148 5 1 1 34147
0 34149 7 1 2 34144 34148
0 34150 5 1 1 34149
0 34151 7 1 2 44551 34150
0 34152 5 1 1 34151
0 34153 7 1 2 58828 63395
0 34154 7 1 2 64740 34153
0 34155 5 1 1 34154
0 34156 7 1 2 34152 34155
0 34157 5 1 1 34156
0 34158 7 1 2 64691 34157
0 34159 5 1 1 34158
0 34160 7 1 2 45990 52243
0 34161 5 1 1 34160
0 34162 7 1 2 61768 34161
0 34163 5 1 1 34162
0 34164 7 1 2 48132 21973
0 34165 7 1 2 60356 34164
0 34166 7 1 2 63933 34165
0 34167 7 1 2 34163 34166
0 34168 5 1 1 34167
0 34169 7 1 2 34159 34168
0 34170 5 1 1 34169
0 34171 7 1 2 49226 58559
0 34172 7 1 2 34170 34171
0 34173 5 1 1 34172
0 34174 7 1 2 65925 62231
0 34175 7 1 2 66497 51442
0 34176 7 1 2 66876 60096
0 34177 7 1 2 34175 34176
0 34178 7 1 2 34174 34177
0 34179 5 1 1 34178
0 34180 7 1 2 46439 34179
0 34181 7 1 2 34173 34180
0 34182 7 1 2 34131 34181
0 34183 7 1 2 34067 34182
0 34184 5 1 1 34183
0 34185 7 1 2 34011 34184
0 34186 5 1 1 34185
0 34187 7 1 2 64273 67168
0 34188 5 1 1 34187
0 34189 7 2 2 64962 66431
0 34190 7 1 2 60345 67169
0 34191 5 1 1 34190
0 34192 7 2 2 48243 60410
0 34193 5 2 1 67171
0 34194 7 1 2 34191 67173
0 34195 5 1 1 34194
0 34196 7 1 2 48946 34195
0 34197 5 1 1 34196
0 34198 7 1 2 48296 62932
0 34199 5 1 1 34198
0 34200 7 1 2 34197 34199
0 34201 5 1 1 34200
0 34202 7 1 2 45203 34201
0 34203 5 1 1 34202
0 34204 7 3 2 42881 62771
0 34205 7 1 2 59304 61859
0 34206 7 1 2 67175 34205
0 34207 5 1 1 34206
0 34208 7 1 2 34203 34207
0 34209 5 1 1 34208
0 34210 7 1 2 44369 34209
0 34211 5 1 1 34210
0 34212 7 1 2 59067 59638
0 34213 7 1 2 65347 34212
0 34214 7 1 2 67176 34213
0 34215 5 1 1 34214
0 34216 7 1 2 34211 34215
0 34217 5 1 1 34216
0 34218 7 1 2 65931 34217
0 34219 5 1 1 34218
0 34220 7 1 2 54827 48143
0 34221 7 1 2 65362 34220
0 34222 5 1 1 34221
0 34223 7 1 2 40680 52776
0 34224 7 1 2 65773 34223
0 34225 7 1 2 66479 66498
0 34226 7 1 2 34224 34225
0 34227 5 1 1 34226
0 34228 7 1 2 34222 34227
0 34229 7 1 2 34219 34228
0 34230 5 1 1 34229
0 34231 7 1 2 54644 34230
0 34232 5 1 1 34231
0 34233 7 2 2 54043 67145
0 34234 7 1 2 56510 58179
0 34235 7 1 2 67178 34234
0 34236 7 1 2 66356 34235
0 34237 5 1 1 34236
0 34238 7 1 2 34232 34237
0 34239 5 1 1 34238
0 34240 7 1 2 34188 34239
0 34241 5 1 1 34240
0 34242 7 1 2 55008 11221
0 34243 5 1 1 34242
0 34244 7 1 2 49227 66113
0 34245 5 1 1 34244
0 34246 7 1 2 65610 64018
0 34247 5 1 1 34246
0 34248 7 1 2 34245 34247
0 34249 5 1 1 34248
0 34250 7 2 2 57277 34249
0 34251 7 2 2 40505 67180
0 34252 7 1 2 53927 67182
0 34253 5 1 1 34252
0 34254 7 1 2 45063 54435
0 34255 7 1 2 66365 34254
0 34256 7 1 2 62704 66917
0 34257 7 1 2 34255 34256
0 34258 5 1 1 34257
0 34259 7 1 2 34253 34258
0 34260 5 1 1 34259
0 34261 7 1 2 55116 34260
0 34262 5 1 1 34261
0 34263 7 1 2 63149 67170
0 34264 5 1 1 34263
0 34265 7 1 2 63766 67177
0 34266 5 1 1 34265
0 34267 7 1 2 34264 34266
0 34268 5 1 1 34267
0 34269 7 1 2 54834 1337
0 34270 7 1 2 15097 34269
0 34271 7 1 2 34268 34270
0 34272 5 1 1 34271
0 34273 7 1 2 59912 66957
0 34274 5 1 1 34273
0 34275 7 1 2 59077 51461
0 34276 7 1 2 66432 34275
0 34277 5 1 1 34276
0 34278 7 1 2 34274 34277
0 34279 5 1 1 34278
0 34280 7 1 2 52938 34279
0 34281 5 1 1 34280
0 34282 7 2 2 52609 59751
0 34283 7 1 2 61883 67184
0 34284 5 1 1 34283
0 34285 7 2 2 54436 64605
0 34286 7 2 2 62304 64607
0 34287 7 1 2 67186 67188
0 34288 5 1 1 34287
0 34289 7 1 2 34284 34288
0 34290 5 1 1 34289
0 34291 7 1 2 49228 34290
0 34292 5 1 1 34291
0 34293 7 1 2 34281 34292
0 34294 7 1 2 34272 34293
0 34295 5 1 1 34294
0 34296 7 1 2 65990 34295
0 34297 5 1 1 34296
0 34298 7 1 2 65170 56355
0 34299 7 1 2 64819 34298
0 34300 7 1 2 50101 34299
0 34301 7 1 2 62134 34300
0 34302 5 1 1 34301
0 34303 7 1 2 34297 34302
0 34304 7 1 2 34262 34303
0 34305 5 1 1 34304
0 34306 7 1 2 45204 34305
0 34307 5 1 1 34306
0 34308 7 2 2 62848 64351
0 34309 7 1 2 41851 67190
0 34310 7 1 2 67181 34309
0 34311 5 1 1 34310
0 34312 7 1 2 34307 34311
0 34313 5 1 1 34312
0 34314 7 1 2 44370 34313
0 34315 5 1 1 34314
0 34316 7 1 2 65353 67183
0 34317 5 1 1 34316
0 34318 7 1 2 34315 34317
0 34319 5 1 1 34318
0 34320 7 1 2 34243 34319
0 34321 5 1 1 34320
0 34322 7 1 2 34241 34321
0 34323 7 1 2 34186 34322
0 34324 5 1 1 34323
0 34325 7 1 2 43594 34324
0 34326 5 1 1 34325
0 34327 7 1 2 58051 67129
0 34328 5 1 1 34327
0 34329 7 1 2 48565 65137
0 34330 5 1 1 34329
0 34331 7 1 2 34328 34330
0 34332 5 1 1 34331
0 34333 7 1 2 45991 34332
0 34334 5 1 1 34333
0 34335 7 1 2 50956 59548
0 34336 5 1 1 34335
0 34337 7 1 2 65139 34336
0 34338 5 1 1 34337
0 34339 7 1 2 54327 34338
0 34340 5 1 1 34339
0 34341 7 1 2 34334 34340
0 34342 5 1 1 34341
0 34343 7 1 2 42882 34342
0 34344 5 1 1 34343
0 34345 7 1 2 55393 67130
0 34346 5 1 1 34345
0 34347 7 1 2 34344 34346
0 34348 5 1 1 34347
0 34349 7 1 2 50347 34348
0 34350 5 1 1 34349
0 34351 7 2 2 66204 62756
0 34352 7 1 2 59573 67192
0 34353 5 1 1 34352
0 34354 7 1 2 34350 34353
0 34355 5 1 1 34354
0 34356 7 1 2 44706 34355
0 34357 5 1 1 34356
0 34358 7 1 2 67193 67141
0 34359 5 1 1 34358
0 34360 7 1 2 34357 34359
0 34361 5 1 1 34360
0 34362 7 1 2 44552 34361
0 34363 5 1 1 34362
0 34364 7 1 2 61317 59599
0 34365 7 1 2 54815 34364
0 34366 7 1 2 65578 34365
0 34367 5 1 1 34366
0 34368 7 1 2 34363 34367
0 34369 5 1 1 34368
0 34370 7 1 2 54986 34369
0 34371 5 1 1 34370
0 34372 7 1 2 40681 66931
0 34373 5 1 1 34372
0 34374 7 1 2 53296 65939
0 34375 5 1 1 34374
0 34376 7 1 2 34373 34375
0 34377 5 1 1 34376
0 34378 7 1 2 40506 34377
0 34379 5 1 1 34378
0 34380 7 1 2 66275 62193
0 34381 7 1 2 53674 34380
0 34382 5 1 1 34381
0 34383 7 1 2 34379 34382
0 34384 5 1 1 34383
0 34385 7 1 2 65127 34384
0 34386 5 1 1 34385
0 34387 7 1 2 34371 34386
0 34388 5 1 1 34387
0 34389 7 1 2 55117 34388
0 34390 5 1 1 34389
0 34391 7 1 2 53782 56667
0 34392 5 1 1 34391
0 34393 7 1 2 67003 34392
0 34394 5 1 1 34393
0 34395 7 1 2 64352 59389
0 34396 7 2 2 65094 34395
0 34397 7 1 2 45205 67194
0 34398 7 1 2 34394 34397
0 34399 5 1 1 34398
0 34400 7 1 2 34390 34399
0 34401 5 1 1 34400
0 34402 7 1 2 43595 34401
0 34403 5 1 1 34402
0 34404 7 1 2 58052 55543
0 34405 5 1 1 34404
0 34406 7 1 2 65658 34405
0 34407 5 1 1 34406
0 34408 7 1 2 42883 34407
0 34409 5 1 1 34408
0 34410 7 1 2 56014 61141
0 34411 5 1 1 34410
0 34412 7 1 2 34409 34411
0 34413 5 2 1 34412
0 34414 7 1 2 60090 66412
0 34415 5 1 1 34414
0 34416 7 1 2 41852 58900
0 34417 5 1 1 34416
0 34418 7 1 2 34415 34417
0 34419 5 1 1 34418
0 34420 7 1 2 67196 34419
0 34421 5 1 1 34420
0 34422 7 1 2 55015 59635
0 34423 5 1 1 34422
0 34424 7 1 2 8126 27099
0 34425 5 1 1 34424
0 34426 7 1 2 41034 59061
0 34427 7 1 2 34425 34426
0 34428 5 1 1 34427
0 34429 7 1 2 34423 34428
0 34430 5 1 1 34429
0 34431 7 2 2 56869 58786
0 34432 7 1 2 34430 67198
0 34433 5 1 1 34432
0 34434 7 1 2 34421 34433
0 34435 5 1 1 34434
0 34436 7 1 2 47098 34435
0 34437 5 1 1 34436
0 34438 7 3 2 55118 60582
0 34439 7 1 2 53709 67200
0 34440 7 2 2 66205 34439
0 34441 7 1 2 41853 67203
0 34442 5 1 1 34441
0 34443 7 1 2 34437 34442
0 34444 5 1 1 34443
0 34445 7 1 2 43034 34444
0 34446 5 1 1 34445
0 34447 7 1 2 66103 63756
0 34448 7 1 2 66009 34447
0 34449 5 1 1 34448
0 34450 7 1 2 34446 34449
0 34451 5 1 1 34450
0 34452 7 1 2 66329 34451
0 34453 5 1 1 34452
0 34454 7 1 2 34403 34453
0 34455 5 1 1 34454
0 34456 7 1 2 44371 34455
0 34457 5 1 1 34456
0 34458 7 1 2 65515 67197
0 34459 5 1 1 34458
0 34460 7 1 2 58901 67199
0 34461 5 1 1 34460
0 34462 7 1 2 34459 34461
0 34463 5 1 1 34462
0 34464 7 1 2 42184 34463
0 34465 5 1 1 34464
0 34466 7 1 2 50598 47882
0 34467 7 1 2 54418 34466
0 34468 7 1 2 67201 34467
0 34469 5 1 1 34468
0 34470 7 1 2 34465 34469
0 34471 5 1 1 34470
0 34472 7 1 2 44553 34471
0 34473 5 1 1 34472
0 34474 7 1 2 43963 53710
0 34475 5 1 1 34474
0 34476 7 1 2 56141 61008
0 34477 5 1 1 34476
0 34478 7 1 2 34475 34477
0 34479 5 2 1 34478
0 34480 7 1 2 54367 67205
0 34481 5 1 1 34480
0 34482 7 1 2 58013 66056
0 34483 5 1 1 34482
0 34484 7 1 2 55465 55726
0 34485 7 1 2 63352 34484
0 34486 5 1 1 34485
0 34487 7 1 2 34483 34486
0 34488 7 1 2 34481 34487
0 34489 5 1 1 34488
0 34490 7 1 2 67202 34489
0 34491 5 1 1 34490
0 34492 7 1 2 34473 34491
0 34493 5 1 1 34492
0 34494 7 1 2 43777 34493
0 34495 5 1 1 34494
0 34496 7 1 2 47739 67204
0 34497 5 1 1 34496
0 34498 7 1 2 34495 34497
0 34499 5 1 1 34498
0 34500 7 1 2 34499 67143
0 34501 5 1 1 34500
0 34502 7 1 2 34457 34501
0 34503 5 1 1 34502
0 34504 7 1 2 49229 34503
0 34505 5 1 1 34504
0 34506 7 1 2 61522 63107
0 34507 7 1 2 55524 34506
0 34508 5 1 1 34507
0 34509 7 1 2 41820 51934
0 34510 7 1 2 56683 49842
0 34511 7 1 2 34509 34510
0 34512 5 1 1 34511
0 34513 7 1 2 34508 34512
0 34514 5 1 1 34513
0 34515 7 1 2 42185 34514
0 34516 5 1 1 34515
0 34517 7 1 2 45522 59964
0 34518 7 1 2 47883 34517
0 34519 7 1 2 56015 34518
0 34520 5 1 1 34519
0 34521 7 1 2 34516 34520
0 34522 5 1 1 34521
0 34523 7 1 2 44554 34522
0 34524 5 1 1 34523
0 34525 7 1 2 59431 63187
0 34526 7 1 2 67206 34525
0 34527 5 1 1 34526
0 34528 7 1 2 34524 34527
0 34529 5 1 1 34528
0 34530 7 1 2 44293 34529
0 34531 5 1 1 34530
0 34532 7 1 2 56040 66306
0 34533 5 1 1 34532
0 34534 7 1 2 45992 66309
0 34535 5 1 1 34534
0 34536 7 1 2 34533 34535
0 34537 5 1 1 34536
0 34538 7 1 2 42448 34537
0 34539 5 1 1 34538
0 34540 7 1 2 42714 50665
0 34541 5 1 1 34540
0 34542 7 1 2 34539 34541
0 34543 5 1 1 34542
0 34544 7 1 2 44707 34543
0 34545 5 1 1 34544
0 34546 7 1 2 53037 52499
0 34547 5 1 1 34546
0 34548 7 1 2 34545 34547
0 34549 5 1 1 34548
0 34550 7 1 2 64963 62880
0 34551 7 1 2 34549 34550
0 34552 5 1 1 34551
0 34553 7 1 2 34531 34552
0 34554 5 1 1 34553
0 34555 7 1 2 43778 34554
0 34556 5 1 1 34555
0 34557 7 1 2 63870 53112
0 34558 7 1 2 66548 34557
0 34559 5 1 1 34558
0 34560 7 1 2 34556 34559
0 34561 5 1 1 34560
0 34562 7 1 2 41537 34561
0 34563 5 1 1 34562
0 34564 7 1 2 52464 62579
0 34565 5 1 1 34564
0 34566 7 1 2 66580 34565
0 34567 5 1 1 34566
0 34568 7 2 2 43596 58917
0 34569 5 1 1 67207
0 34570 7 1 2 51400 67208
0 34571 7 1 2 34567 34570
0 34572 5 1 1 34571
0 34573 7 1 2 34563 34572
0 34574 5 1 1 34573
0 34575 7 1 2 43035 34574
0 34576 5 1 1 34575
0 34577 7 1 2 58907 34569
0 34578 5 1 1 34577
0 34579 7 1 2 65520 59920
0 34580 7 1 2 63404 34579
0 34581 7 1 2 34578 34580
0 34582 5 1 1 34581
0 34583 7 1 2 34576 34582
0 34584 5 1 1 34583
0 34585 7 1 2 51564 34584
0 34586 5 1 1 34585
0 34587 7 2 2 56097 58726
0 34588 7 1 2 64972 67209
0 34589 5 1 1 34588
0 34590 7 1 2 66618 63947
0 34591 7 1 2 55544 34590
0 34592 5 1 1 34591
0 34593 7 1 2 34589 34592
0 34594 5 1 1 34593
0 34595 7 1 2 44294 34594
0 34596 5 1 1 34595
0 34597 7 1 2 55021 49792
0 34598 7 1 2 67210 34597
0 34599 5 1 1 34598
0 34600 7 1 2 34596 34599
0 34601 5 1 1 34600
0 34602 7 2 2 43150 47099
0 34603 7 1 2 43779 64399
0 34604 7 1 2 67211 34603
0 34605 7 1 2 34601 34604
0 34606 5 1 1 34605
0 34607 7 1 2 34586 34606
0 34608 5 1 1 34607
0 34609 7 1 2 46593 34608
0 34610 5 1 1 34609
0 34611 7 1 2 55525 66619
0 34612 5 1 1 34611
0 34613 7 1 2 59262 60649
0 34614 5 1 1 34613
0 34615 7 1 2 34612 34614
0 34616 5 1 1 34615
0 34617 7 1 2 62580 34616
0 34618 5 1 1 34617
0 34619 7 1 2 62523 62189
0 34620 7 1 2 55622 34619
0 34621 5 1 1 34620
0 34622 7 1 2 34618 34621
0 34623 5 1 1 34622
0 34624 7 1 2 43036 34623
0 34625 5 1 1 34624
0 34626 7 1 2 51055 66585
0 34627 7 1 2 49845 34626
0 34628 5 1 1 34627
0 34629 7 1 2 34625 34628
0 34630 5 1 1 34629
0 34631 7 1 2 51565 34630
0 34632 5 1 1 34631
0 34633 7 1 2 55805 66504
0 34634 7 1 2 67066 49794
0 34635 7 1 2 34633 34634
0 34636 5 1 1 34635
0 34637 7 1 2 34632 34636
0 34638 5 1 1 34637
0 34639 7 1 2 46440 34638
0 34640 5 1 1 34639
0 34641 7 1 2 55423 66505
0 34642 7 2 2 47937 51489
0 34643 7 1 2 63469 67213
0 34644 7 1 2 34641 34643
0 34645 5 1 1 34644
0 34646 7 1 2 34640 34645
0 34647 5 1 1 34646
0 34648 7 1 2 41821 34647
0 34649 5 1 1 34648
0 34650 7 1 2 49814 56585
0 34651 7 1 2 64139 34650
0 34652 7 1 2 63353 67214
0 34653 7 1 2 34651 34652
0 34654 5 1 1 34653
0 34655 7 1 2 34649 34654
0 34656 5 1 1 34655
0 34657 7 1 2 41035 34656
0 34658 5 1 1 34657
0 34659 7 1 2 64140 49733
0 34660 7 2 2 49815 54447
0 34661 7 1 2 66325 63470
0 34662 7 1 2 67215 34661
0 34663 7 1 2 34659 34662
0 34664 5 1 1 34663
0 34665 7 1 2 34658 34664
0 34666 5 1 1 34665
0 34667 7 1 2 64692 34666
0 34668 5 1 1 34667
0 34669 7 1 2 34610 34668
0 34670 5 1 1 34669
0 34671 7 1 2 43265 34670
0 34672 5 1 1 34671
0 34673 7 2 2 59567 63267
0 34674 7 1 2 48011 67217
0 34675 5 1 1 34674
0 34676 7 1 2 49387 57238
0 34677 7 1 2 61391 34676
0 34678 7 1 2 60091 34677
0 34679 5 1 1 34678
0 34680 7 1 2 34675 34679
0 34681 5 1 1 34680
0 34682 7 1 2 45789 34681
0 34683 5 1 1 34682
0 34684 7 1 2 50599 67218
0 34685 5 1 1 34684
0 34686 7 1 2 34683 34685
0 34687 5 1 1 34686
0 34688 7 1 2 43780 34687
0 34689 5 1 1 34688
0 34690 7 1 2 47740 59379
0 34691 7 1 2 66550 34690
0 34692 5 1 1 34691
0 34693 7 1 2 34689 34692
0 34694 5 1 1 34693
0 34695 7 1 2 43151 34694
0 34696 5 1 1 34695
0 34697 7 1 2 46985 48170
0 34698 5 2 1 34697
0 34699 7 1 2 34091 67219
0 34700 5 1 1 34699
0 34701 7 1 2 59614 66775
0 34702 7 1 2 59294 34701
0 34703 7 1 2 34700 34702
0 34704 5 1 1 34703
0 34705 7 1 2 34696 34704
0 34706 5 1 1 34705
0 34707 7 1 2 43266 34706
0 34708 5 1 1 34707
0 34709 7 1 2 62780 65076
0 34710 7 1 2 51566 34709
0 34711 7 1 2 66473 34710
0 34712 5 1 1 34711
0 34713 7 1 2 34708 34712
0 34714 5 1 1 34713
0 34715 7 1 2 40682 34714
0 34716 5 1 1 34715
0 34717 7 2 2 63972 59068
0 34718 7 1 2 44974 67221
0 34719 7 1 2 66291 34718
0 34720 5 1 1 34719
0 34721 7 1 2 55119 59517
0 34722 5 1 1 34721
0 34723 7 1 2 34720 34722
0 34724 5 1 1 34723
0 34725 7 1 2 46441 50780
0 34726 7 1 2 60150 65077
0 34727 7 1 2 34725 34726
0 34728 7 1 2 34724 34727
0 34729 5 1 1 34728
0 34730 7 1 2 34716 34729
0 34731 5 1 1 34730
0 34732 7 1 2 44372 34731
0 34733 5 1 1 34732
0 34734 7 1 2 49892 53711
0 34735 5 1 1 34734
0 34736 7 1 2 67220 34735
0 34737 5 1 1 34736
0 34738 7 1 2 63300 34737
0 34739 5 1 1 34738
0 34740 7 2 2 44295 44555
0 34741 7 2 2 40887 67223
0 34742 7 1 2 60226 56586
0 34743 7 1 2 66389 34742
0 34744 7 1 2 67225 34743
0 34745 5 1 1 34744
0 34746 7 1 2 34739 34745
0 34747 5 1 1 34746
0 34748 7 1 2 40683 46552
0 34749 7 1 2 60372 34748
0 34750 7 1 2 34747 34749
0 34751 5 1 1 34750
0 34752 7 1 2 34733 34751
0 34753 5 1 1 34752
0 34754 7 1 2 65554 34753
0 34755 5 1 1 34754
0 34756 7 1 2 40507 66453
0 34757 5 1 1 34756
0 34758 7 1 2 46986 52695
0 34759 7 1 2 66403 34758
0 34760 5 1 1 34759
0 34761 7 1 2 34757 34760
0 34762 5 1 1 34761
0 34763 7 1 2 63789 34762
0 34764 5 1 1 34763
0 34765 7 2 2 44975 60692
0 34766 7 1 2 63020 67227
0 34767 7 1 2 64949 34766
0 34768 5 1 1 34767
0 34769 7 1 2 34764 34768
0 34770 5 1 1 34769
0 34771 7 1 2 55120 34770
0 34772 5 1 1 34771
0 34773 7 1 2 66454 67195
0 34774 5 1 1 34773
0 34775 7 1 2 56045 61250
0 34776 7 1 2 60013 34775
0 34777 7 1 2 59755 34776
0 34778 5 1 1 34777
0 34779 7 1 2 34774 34778
0 34780 5 1 1 34779
0 34781 7 1 2 57813 34780
0 34782 5 1 1 34781
0 34783 7 1 2 34772 34782
0 34784 5 1 1 34783
0 34785 7 1 2 43597 34784
0 34786 5 1 1 34785
0 34787 7 1 2 60227 55731
0 34788 7 1 2 62774 34787
0 34789 7 1 2 63265 34788
0 34790 7 1 2 66404 34789
0 34791 5 1 1 34790
0 34792 7 1 2 34786 34791
0 34793 5 1 1 34792
0 34794 7 1 2 45206 34793
0 34795 5 1 1 34794
0 34796 7 1 2 58902 66405
0 34797 5 1 1 34796
0 34798 7 1 2 44296 50121
0 34799 7 1 2 62789 34798
0 34800 5 1 1 34799
0 34801 7 1 2 34797 34800
0 34802 5 1 1 34801
0 34803 7 1 2 57506 34802
0 34804 5 1 1 34803
0 34805 7 2 2 60670 56587
0 34806 7 1 2 62781 54935
0 34807 7 1 2 58626 34806
0 34808 7 1 2 67229 34807
0 34809 5 1 1 34808
0 34810 7 1 2 34804 34809
0 34811 5 1 1 34810
0 34812 7 2 2 62715 34811
0 34813 7 1 2 44556 66250
0 34814 7 1 2 67231 34813
0 34815 5 1 1 34814
0 34816 7 1 2 34795 34815
0 34817 5 1 1 34816
0 34818 7 1 2 44373 34817
0 34819 5 1 1 34818
0 34820 7 1 2 66533 67232
0 34821 5 1 1 34820
0 34822 7 1 2 34819 34821
0 34823 5 1 1 34822
0 34824 7 1 2 54368 34823
0 34825 5 1 1 34824
0 34826 7 1 2 58129 59267
0 34827 5 1 1 34826
0 34828 7 1 2 47151 34827
0 34829 5 1 1 34828
0 34830 7 1 2 43449 67164
0 34831 5 1 1 34830
0 34832 7 1 2 34829 34831
0 34833 5 1 1 34832
0 34834 7 1 2 66302 34833
0 34835 5 1 1 34834
0 34836 7 1 2 62540 65165
0 34837 7 1 2 66363 58121
0 34838 7 1 2 34836 34837
0 34839 7 1 2 66622 34838
0 34840 5 1 1 34839
0 34841 7 1 2 34835 34840
0 34842 5 1 1 34841
0 34843 7 1 2 42715 34842
0 34844 5 1 1 34843
0 34845 7 2 2 51935 50257
0 34846 7 1 2 66348 67233
0 34847 5 1 1 34846
0 34848 7 1 2 34844 34847
0 34849 5 1 1 34848
0 34850 7 1 2 46170 34849
0 34851 5 1 1 34850
0 34852 7 1 2 62228 62907
0 34853 7 1 2 59896 34852
0 34854 7 1 2 66546 34853
0 34855 5 1 1 34854
0 34856 7 1 2 34851 34855
0 34857 5 1 1 34856
0 34858 7 1 2 58053 34857
0 34859 5 1 1 34858
0 34860 7 1 2 67230 64528
0 34861 7 1 2 63480 34860
0 34862 5 1 1 34861
0 34863 7 1 2 40119 66935
0 34864 5 1 1 34863
0 34865 7 1 2 55121 34864
0 34866 7 1 2 66937 34865
0 34867 5 1 1 34866
0 34868 7 1 2 34862 34867
0 34869 5 1 1 34868
0 34870 7 2 2 49816 48840
0 34871 5 1 1 67235
0 34872 7 1 2 65493 67212
0 34873 7 1 2 67236 34872
0 34874 7 1 2 34869 34873
0 34875 5 1 1 34874
0 34876 7 1 2 34859 34875
0 34877 7 1 2 34825 34876
0 34878 7 1 2 34755 34877
0 34879 7 1 2 34672 34878
0 34880 7 1 2 34505 34879
0 34881 5 1 1 34880
0 34882 7 1 2 49066 34881
0 34883 5 1 1 34882
0 34884 7 1 2 45124 57735
0 34885 5 1 1 34884
0 34886 7 1 2 59275 63423
0 34887 5 1 1 34886
0 34888 7 1 2 34885 34887
0 34889 5 1 1 34888
0 34890 7 1 2 44297 34889
0 34891 5 1 1 34890
0 34892 7 1 2 51701 58678
0 34893 5 1 1 34892
0 34894 7 1 2 34891 34893
0 34895 5 1 1 34894
0 34896 7 1 2 5095 65209
0 34897 5 1 1 34896
0 34898 7 1 2 54044 65427
0 34899 7 1 2 34897 34898
0 34900 5 1 1 34899
0 34901 7 1 2 64693 65078
0 34902 7 1 2 52663 34901
0 34903 7 1 2 66701 34902
0 34904 5 1 1 34903
0 34905 7 1 2 34900 34904
0 34906 5 1 1 34905
0 34907 7 1 2 44557 34906
0 34908 5 1 1 34907
0 34909 7 1 2 51936 47884
0 34910 5 1 1 34909
0 34911 7 1 2 43450 53388
0 34912 5 1 1 34911
0 34913 7 1 2 34910 34912
0 34914 5 1 1 34913
0 34915 7 2 2 54625 52696
0 34916 7 1 2 41271 67062
0 34917 7 1 2 67237 34916
0 34918 7 1 2 34914 34917
0 34919 5 1 1 34918
0 34920 7 1 2 34908 34919
0 34921 5 1 1 34920
0 34922 7 1 2 34895 34921
0 34923 5 1 1 34922
0 34924 7 1 2 62829 66066
0 34925 5 1 1 34924
0 34926 7 1 2 56709 57863
0 34927 7 2 2 63108 34926
0 34928 5 1 1 67239
0 34929 7 1 2 62849 67240
0 34930 5 1 1 34929
0 34931 7 1 2 34925 34930
0 34932 5 1 1 34931
0 34933 7 1 2 58054 34932
0 34934 5 1 1 34933
0 34935 7 2 2 42716 56826
0 34936 5 2 1 67241
0 34937 7 1 2 65659 67243
0 34938 5 1 1 34937
0 34939 7 1 2 62830 34938
0 34940 5 1 1 34939
0 34941 7 2 2 44298 62165
0 34942 7 1 2 42449 66386
0 34943 7 1 2 67245 34942
0 34944 5 1 1 34943
0 34945 7 1 2 34940 34944
0 34946 5 1 1 34945
0 34947 7 1 2 47100 34946
0 34948 5 1 1 34947
0 34949 7 1 2 34934 34948
0 34950 5 1 1 34949
0 34951 7 1 2 46171 34950
0 34952 5 1 1 34951
0 34953 7 1 2 62831 65901
0 34954 5 1 1 34953
0 34955 7 1 2 62176 67224
0 34956 7 1 2 66598 34955
0 34957 5 1 1 34956
0 34958 7 1 2 34954 34957
0 34959 5 1 1 34958
0 34960 7 1 2 67147 34959
0 34961 5 1 1 34960
0 34962 7 1 2 34952 34961
0 34963 5 1 1 34962
0 34964 7 1 2 43037 34963
0 34965 5 1 1 34964
0 34966 7 1 2 55358 66187
0 34967 7 1 2 65699 34966
0 34968 5 1 1 34967
0 34969 7 1 2 34965 34968
0 34970 5 1 1 34969
0 34971 7 1 2 43781 34970
0 34972 5 1 1 34971
0 34973 7 1 2 40508 67010
0 34974 5 2 1 34973
0 34975 7 1 2 64181 54958
0 34976 5 1 1 34975
0 34977 7 1 2 67247 34976
0 34978 5 1 1 34977
0 34979 7 2 2 65711 34978
0 34980 7 1 2 43451 63973
0 34981 7 1 2 62850 34980
0 34982 7 1 2 67249 34981
0 34983 5 1 1 34982
0 34984 7 1 2 34972 34983
0 34985 5 1 1 34984
0 34986 7 1 2 46594 34985
0 34987 5 1 1 34986
0 34988 7 1 2 59965 66067
0 34989 5 1 1 34988
0 34990 7 1 2 34928 34989
0 34991 5 1 1 34990
0 34992 7 1 2 58055 34991
0 34993 5 1 1 34992
0 34994 7 1 2 65513 67242
0 34995 5 1 1 34994
0 34996 7 1 2 65709 64970
0 34997 5 1 1 34996
0 34998 7 1 2 34995 34997
0 34999 5 1 1 34998
0 35000 7 1 2 47101 34999
0 35001 5 1 1 35000
0 35002 7 1 2 34993 35001
0 35003 5 1 1 35002
0 35004 7 1 2 46172 35003
0 35005 5 1 1 35004
0 35006 7 1 2 47102 65509
0 35007 5 1 1 35006
0 35008 7 1 2 41822 65953
0 35009 5 1 1 35008
0 35010 7 1 2 35007 35009
0 35011 5 1 1 35010
0 35012 7 1 2 45790 35011
0 35013 5 1 1 35012
0 35014 7 1 2 28762 35013
0 35015 5 1 1 35014
0 35016 7 1 2 67148 35015
0 35017 5 1 1 35016
0 35018 7 1 2 35005 35017
0 35019 5 1 1 35018
0 35020 7 1 2 43782 35019
0 35021 5 1 1 35020
0 35022 7 1 2 63109 67250
0 35023 5 1 1 35022
0 35024 7 1 2 35021 35023
0 35025 5 1 1 35024
0 35026 7 1 2 41036 35025
0 35027 5 1 1 35026
0 35028 7 1 2 47152 59854
0 35029 5 1 1 35028
0 35030 7 1 2 67248 35029
0 35031 5 1 1 35030
0 35032 7 1 2 58056 35031
0 35033 5 1 1 35032
0 35034 7 2 2 60978 66276
0 35035 7 1 2 66710 67251
0 35036 5 1 1 35035
0 35037 7 1 2 35033 35036
0 35038 5 1 1 35037
0 35039 7 2 2 61566 35038
0 35040 7 1 2 66434 67253
0 35041 5 1 1 35040
0 35042 7 1 2 35027 35041
0 35043 5 1 1 35042
0 35044 7 1 2 53928 35043
0 35045 5 1 1 35044
0 35046 7 1 2 43452 62342
0 35047 7 1 2 67254 35046
0 35048 5 1 1 35047
0 35049 7 1 2 35045 35048
0 35050 5 1 1 35049
0 35051 7 1 2 43038 35050
0 35052 5 1 1 35051
0 35053 7 1 2 42717 58812
0 35054 7 2 2 49616 59082
0 35055 7 1 2 64242 67255
0 35056 7 1 2 60391 35055
0 35057 7 1 2 35053 35056
0 35058 5 1 1 35057
0 35059 7 1 2 35052 35058
0 35060 5 1 1 35059
0 35061 7 1 2 64694 35060
0 35062 5 1 1 35061
0 35063 7 1 2 34987 35062
0 35064 5 1 1 35063
0 35065 7 1 2 41681 35064
0 35066 5 1 1 35065
0 35067 7 1 2 43453 59197
0 35068 5 1 1 35067
0 35069 7 1 2 60496 35068
0 35070 5 1 1 35069
0 35071 7 1 2 47103 35070
0 35072 5 1 1 35071
0 35073 7 1 2 49455 60920
0 35074 5 1 1 35073
0 35075 7 1 2 35072 35074
0 35076 5 1 1 35075
0 35077 7 1 2 58057 35076
0 35078 5 1 1 35077
0 35079 7 1 2 64407 54729
0 35080 5 1 1 35079
0 35081 7 1 2 67244 35080
0 35082 5 1 1 35081
0 35083 7 1 2 52363 35082
0 35084 5 1 1 35083
0 35085 7 1 2 35078 35084
0 35086 5 1 1 35085
0 35087 7 1 2 42884 35086
0 35088 5 1 1 35087
0 35089 7 1 2 49548 56016
0 35090 7 1 2 63405 35089
0 35091 5 1 1 35090
0 35092 7 1 2 35088 35091
0 35093 5 1 1 35092
0 35094 7 1 2 46307 35093
0 35095 5 1 1 35094
0 35096 7 1 2 48171 57602
0 35097 7 1 2 67252 35096
0 35098 5 1 1 35097
0 35099 7 1 2 35095 35098
0 35100 5 1 1 35099
0 35101 7 1 2 44976 43152
0 35102 7 1 2 65274 35101
0 35103 7 1 2 35100 35102
0 35104 5 1 1 35103
0 35105 7 1 2 40888 35104
0 35106 7 1 2 35066 35105
0 35107 5 1 1 35106
0 35108 7 1 2 53363 50412
0 35109 5 1 1 35108
0 35110 7 1 2 55526 35109
0 35111 7 1 2 65275 35110
0 35112 5 1 1 35111
0 35113 7 1 2 49617 57730
0 35114 7 1 2 66781 35113
0 35115 5 1 1 35114
0 35116 7 1 2 35112 35115
0 35117 5 1 1 35116
0 35118 7 1 2 43454 35117
0 35119 5 1 1 35118
0 35120 7 1 2 55806 56143
0 35121 7 1 2 65276 35120
0 35122 5 1 1 35121
0 35123 7 1 2 46308 35122
0 35124 7 1 2 35119 35123
0 35125 5 1 1 35124
0 35126 7 1 2 66770 67256
0 35127 5 1 1 35126
0 35128 7 1 2 61881 51222
0 35129 7 1 2 60718 35128
0 35130 5 1 1 35129
0 35131 7 1 2 35127 35130
0 35132 5 1 1 35131
0 35133 7 1 2 55122 35132
0 35134 5 1 1 35133
0 35135 7 1 2 48841 64707
0 35136 5 1 1 35135
0 35137 7 1 2 45125 60058
0 35138 7 1 2 57980 35137
0 35139 7 1 2 62181 35138
0 35140 5 1 1 35139
0 35141 7 1 2 35136 35140
0 35142 7 1 2 35134 35141
0 35143 5 1 1 35142
0 35144 7 1 2 46595 35143
0 35145 5 1 1 35144
0 35146 7 1 2 65457 59315
0 35147 7 1 2 55346 35146
0 35148 7 1 2 65343 35147
0 35149 5 1 1 35148
0 35150 7 1 2 65536 57160
0 35151 7 1 2 63089 35150
0 35152 7 1 2 66779 35151
0 35153 5 1 1 35152
0 35154 7 1 2 43039 35153
0 35155 7 1 2 35149 35154
0 35156 7 1 2 35145 35155
0 35157 5 1 1 35156
0 35158 7 1 2 52244 35157
0 35159 7 1 2 35125 35158
0 35160 5 1 1 35159
0 35161 7 1 2 66060 52939
0 35162 5 1 1 35161
0 35163 7 1 2 53689 58495
0 35164 5 1 1 35163
0 35165 7 1 2 35162 35164
0 35166 5 1 1 35165
0 35167 7 1 2 43783 35166
0 35168 5 1 1 35167
0 35169 7 1 2 66137 55716
0 35170 5 1 1 35169
0 35171 7 1 2 35168 35170
0 35172 5 1 1 35171
0 35173 7 1 2 43455 35172
0 35174 5 1 1 35173
0 35175 7 1 2 56710 47959
0 35176 7 1 2 50269 35175
0 35177 5 1 1 35176
0 35178 7 1 2 35174 35177
0 35179 5 1 1 35178
0 35180 7 1 2 46309 58058
0 35181 7 1 2 65277 35180
0 35182 7 1 2 35179 35181
0 35183 5 1 1 35182
0 35184 7 1 2 35160 35183
0 35185 5 1 1 35184
0 35186 7 1 2 43153 35185
0 35187 5 1 1 35186
0 35188 7 1 2 61979 59323
0 35189 7 1 2 61142 35188
0 35190 7 1 2 66724 67179
0 35191 7 1 2 35189 35190
0 35192 5 1 1 35191
0 35193 7 1 2 44137 35192
0 35194 7 1 2 35187 35193
0 35195 5 1 1 35194
0 35196 7 1 2 43267 35195
0 35197 7 1 2 35107 35196
0 35198 5 1 1 35197
0 35199 7 1 2 34923 35198
0 35200 7 1 2 34883 35199
0 35201 7 1 2 34326 35200
0 35202 5 1 1 35201
0 35203 7 1 2 46851 35202
0 35204 5 1 1 35203
0 35205 7 1 2 54849 66138
0 35206 7 1 2 66171 35205
0 35207 5 1 1 35206
0 35208 7 1 2 61221 62185
0 35209 7 1 2 49785 35208
0 35210 5 1 1 35209
0 35211 7 1 2 35207 35210
0 35212 5 1 1 35211
0 35213 7 1 2 64246 35212
0 35214 5 1 1 35213
0 35215 7 1 2 55354 65199
0 35216 5 1 1 35215
0 35217 7 1 2 64933 65932
0 35218 5 1 1 35217
0 35219 7 1 2 50964 66149
0 35220 5 2 1 35219
0 35221 7 1 2 67234 67257
0 35222 5 1 1 35221
0 35223 7 1 2 35218 35222
0 35224 5 1 1 35223
0 35225 7 1 2 47430 35224
0 35226 5 1 1 35225
0 35227 7 1 2 46173 35226
0 35228 7 1 2 35216 35227
0 35229 5 1 1 35228
0 35230 7 1 2 40298 65704
0 35231 5 1 1 35230
0 35232 7 1 2 64342 35231
0 35233 5 1 1 35232
0 35234 7 1 2 40684 35233
0 35235 5 1 1 35234
0 35236 7 1 2 53478 53019
0 35237 5 1 1 35236
0 35238 7 1 2 35235 35237
0 35239 5 1 1 35238
0 35240 7 1 2 46879 35239
0 35241 5 1 1 35240
0 35242 7 1 2 40299 51937
0 35243 5 1 1 35242
0 35244 7 1 2 46903 52530
0 35245 5 1 1 35244
0 35246 7 1 2 35243 35245
0 35247 5 1 1 35246
0 35248 7 1 2 40685 35247
0 35249 5 1 1 35248
0 35250 7 2 2 43964 50234
0 35251 7 1 2 65733 67259
0 35252 5 1 1 35251
0 35253 7 1 2 35249 35252
0 35254 5 1 1 35253
0 35255 7 1 2 40120 35254
0 35256 5 1 1 35255
0 35257 7 1 2 57174 66197
0 35258 5 1 1 35257
0 35259 7 1 2 35256 35258
0 35260 5 1 1 35259
0 35261 7 1 2 41408 35260
0 35262 5 1 1 35261
0 35263 7 2 2 45346 51938
0 35264 7 1 2 66033 53169
0 35265 7 1 2 67261 35264
0 35266 5 1 1 35265
0 35267 7 1 2 35262 35266
0 35268 7 1 2 35241 35267
0 35269 5 1 1 35268
0 35270 7 1 2 40509 35269
0 35271 5 1 1 35270
0 35272 7 1 2 40686 65197
0 35273 5 1 1 35272
0 35274 7 1 2 52988 62388
0 35275 5 1 1 35274
0 35276 7 1 2 35273 35275
0 35277 5 1 1 35276
0 35278 7 1 2 40510 35277
0 35279 5 1 1 35278
0 35280 7 1 2 49295 64450
0 35281 5 1 1 35280
0 35282 7 1 2 35279 35281
0 35283 5 1 1 35282
0 35284 7 1 2 56121 35283
0 35285 5 1 1 35284
0 35286 7 1 2 62281 63135
0 35287 7 1 2 67262 35286
0 35288 5 1 1 35287
0 35289 7 1 2 42885 35288
0 35290 7 1 2 35285 35289
0 35291 7 1 2 35271 35290
0 35292 5 1 1 35291
0 35293 7 1 2 46310 35292
0 35294 7 1 2 35229 35293
0 35295 5 1 1 35294
0 35296 7 1 2 44828 35295
0 35297 5 1 1 35296
0 35298 7 1 2 42886 65200
0 35299 5 1 1 35298
0 35300 7 1 2 58754 66658
0 35301 5 1 1 35300
0 35302 7 1 2 45993 35301
0 35303 7 1 2 35299 35302
0 35304 5 1 1 35303
0 35305 7 1 2 42887 65186
0 35306 5 1 1 35305
0 35307 7 1 2 64934 66207
0 35308 5 1 1 35307
0 35309 7 1 2 42718 35308
0 35310 7 1 2 35306 35309
0 35311 5 1 1 35310
0 35312 7 1 2 43965 35311
0 35313 7 1 2 35304 35312
0 35314 5 1 1 35313
0 35315 7 1 2 52345 60804
0 35316 7 1 2 52589 35315
0 35317 5 1 1 35316
0 35318 7 1 2 48842 65640
0 35319 7 1 2 67258 35318
0 35320 5 1 1 35319
0 35321 7 1 2 35317 35320
0 35322 5 1 1 35321
0 35323 7 1 2 42719 35322
0 35324 5 1 1 35323
0 35325 7 1 2 41538 35324
0 35326 7 1 2 35314 35325
0 35327 5 1 1 35326
0 35328 7 1 2 46311 35327
0 35329 5 1 1 35328
0 35330 7 1 2 59645 66624
0 35331 7 1 2 66670 35330
0 35332 5 1 1 35331
0 35333 7 1 2 35329 35332
0 35334 5 1 1 35333
0 35335 7 1 2 35297 35334
0 35336 5 1 1 35335
0 35337 7 1 2 35214 35336
0 35338 5 2 1 35337
0 35339 7 1 2 48947 67263
0 35340 5 1 1 35339
0 35341 7 1 2 52263 52059
0 35342 5 1 1 35341
0 35343 7 1 2 50932 35342
0 35344 5 1 1 35343
0 35345 7 1 2 43456 35344
0 35346 5 1 1 35345
0 35347 7 1 2 34871 35346
0 35348 5 1 1 35347
0 35349 7 3 2 58727 35348
0 35350 7 1 2 53929 66310
0 35351 7 1 2 67265 35350
0 35352 5 1 1 35351
0 35353 7 1 2 47431 49751
0 35354 7 1 2 58728 35353
0 35355 7 1 2 64953 60591
0 35356 7 1 2 35354 35355
0 35357 5 1 1 35356
0 35358 7 1 2 35352 35357
0 35359 5 1 1 35358
0 35360 7 1 2 50624 35359
0 35361 5 1 1 35360
0 35362 7 1 2 35340 35361
0 35363 5 1 1 35362
0 35364 7 1 2 66610 35363
0 35365 5 1 1 35364
0 35366 7 1 2 65031 61211
0 35367 5 1 1 35366
0 35368 7 1 2 42720 56238
0 35369 5 1 1 35368
0 35370 7 1 2 35367 35369
0 35371 5 1 1 35370
0 35372 7 1 2 45347 35371
0 35373 5 1 1 35372
0 35374 7 1 2 40511 55470
0 35375 7 1 2 65505 35374
0 35376 5 1 1 35375
0 35377 7 1 2 35373 35376
0 35378 5 1 1 35377
0 35379 7 1 2 45523 35378
0 35380 5 1 1 35379
0 35381 7 1 2 55656 65452
0 35382 5 1 1 35381
0 35383 7 1 2 35380 35382
0 35384 5 1 1 35383
0 35385 7 1 2 52014 35384
0 35386 5 1 1 35385
0 35387 7 1 2 45994 66229
0 35388 5 1 1 35387
0 35389 7 1 2 35386 35388
0 35390 5 1 1 35389
0 35391 7 1 2 58059 35390
0 35392 5 1 1 35391
0 35393 7 1 2 66933 67260
0 35394 7 1 2 66720 35393
0 35395 5 1 1 35394
0 35396 7 1 2 35392 35395
0 35397 5 1 1 35396
0 35398 7 1 2 42888 35397
0 35399 5 1 1 35398
0 35400 7 1 2 66223 35399
0 35401 5 2 1 35400
0 35402 7 1 2 65494 49359
0 35403 7 1 2 67268 35402
0 35404 5 1 1 35403
0 35405 7 1 2 35365 35404
0 35406 5 1 1 35405
0 35407 7 1 2 43154 35406
0 35408 5 1 1 35407
0 35409 7 1 2 40687 61178
0 35410 5 1 1 35409
0 35411 7 1 2 65563 35410
0 35412 5 3 1 35411
0 35413 7 1 2 64850 67270
0 35414 5 1 1 35413
0 35415 7 1 2 58060 64267
0 35416 5 1 1 35415
0 35417 7 1 2 52015 60663
0 35418 5 1 1 35417
0 35419 7 1 2 35416 35418
0 35420 5 1 1 35419
0 35421 7 1 2 42889 35420
0 35422 5 1 1 35421
0 35423 7 1 2 44829 56516
0 35424 5 1 1 35423
0 35425 7 1 2 35422 35424
0 35426 5 1 1 35425
0 35427 7 1 2 61483 35426
0 35428 5 1 1 35427
0 35429 7 1 2 35414 35428
0 35430 5 2 1 35429
0 35431 7 2 2 40512 40970
0 35432 7 1 2 43268 52860
0 35433 7 1 2 67275 35432
0 35434 7 1 2 67273 35433
0 35435 5 1 1 35434
0 35436 7 1 2 53089 58961
0 35437 7 1 2 66212 35436
0 35438 7 1 2 61643 35437
0 35439 7 1 2 66790 35438
0 35440 5 1 1 35439
0 35441 7 1 2 35435 35440
0 35442 5 1 1 35441
0 35443 7 1 2 66195 35442
0 35444 5 1 1 35443
0 35445 7 1 2 35408 35444
0 35446 5 1 1 35445
0 35447 7 1 2 55123 35446
0 35448 5 1 1 35447
0 35449 7 1 2 58990 46596
0 35450 5 1 1 35449
0 35451 7 1 2 65267 35450
0 35452 5 1 1 35451
0 35453 7 1 2 67264 35452
0 35454 5 1 1 35453
0 35455 7 1 2 43966 59258
0 35456 7 1 2 58962 35455
0 35457 7 1 2 67266 35456
0 35458 5 1 1 35457
0 35459 7 2 2 44445 59878
0 35460 7 1 2 62163 66213
0 35461 7 1 2 67277 35460
0 35462 5 1 1 35461
0 35463 7 1 2 35458 35462
0 35464 5 1 1 35463
0 35465 7 1 2 64415 35464
0 35466 5 1 1 35465
0 35467 7 1 2 66269 60250
0 35468 7 1 2 67278 35467
0 35469 5 1 1 35468
0 35470 7 1 2 45064 60014
0 35471 7 1 2 60389 35470
0 35472 7 1 2 67267 35471
0 35473 5 1 1 35472
0 35474 7 1 2 35469 35473
0 35475 5 1 1 35474
0 35476 7 1 2 46597 57148
0 35477 7 1 2 35475 35476
0 35478 5 1 1 35477
0 35479 7 1 2 35466 35478
0 35480 5 1 1 35479
0 35481 7 1 2 50625 35480
0 35482 5 1 1 35481
0 35483 7 1 2 35454 35482
0 35484 5 1 1 35483
0 35485 7 1 2 43155 35484
0 35486 5 1 1 35485
0 35487 7 1 2 46598 67191
0 35488 5 1 1 35487
0 35489 7 1 2 56893 59207
0 35490 7 1 2 66796 35489
0 35491 5 1 1 35490
0 35492 7 1 2 35488 35491
0 35493 5 1 1 35492
0 35494 7 1 2 57963 35493
0 35495 7 1 2 67274 35494
0 35496 5 1 1 35495
0 35497 7 1 2 35486 35496
0 35498 5 1 1 35497
0 35499 7 1 2 43269 35498
0 35500 5 1 1 35499
0 35501 7 1 2 54626 67269
0 35502 5 1 1 35501
0 35503 7 1 2 66215 52541
0 35504 7 1 2 66626 35503
0 35505 5 1 1 35504
0 35506 7 1 2 35502 35505
0 35507 5 1 1 35506
0 35508 7 1 2 53930 65108
0 35509 7 1 2 35507 35508
0 35510 5 1 1 35509
0 35511 7 1 2 35500 35510
0 35512 7 1 2 35448 35511
0 35513 5 1 1 35512
0 35514 7 1 2 51567 35513
0 35515 5 1 1 35514
0 35516 7 1 2 35204 35515
0 35517 7 1 2 33830 35516
0 35518 7 1 2 28477 35517
0 35519 7 1 2 26825 35518
0 35520 7 1 2 24463 35519
0 35521 5 1 1 35520
0 35522 7 1 2 46528 35521
0 35523 5 1 1 35522
0 35524 7 8 2 43270 46529
0 35525 7 1 2 45995 52299
0 35526 5 1 1 35525
0 35527 7 1 2 50240 52557
0 35528 5 1 1 35527
0 35529 7 2 2 45348 35528
0 35530 5 1 1 67287
0 35531 7 1 2 55321 67288
0 35532 5 1 1 35531
0 35533 7 1 2 35526 35532
0 35534 5 1 1 35533
0 35535 7 1 2 49140 35534
0 35536 5 1 1 35535
0 35537 7 2 2 47663 58115
0 35538 5 1 1 67289
0 35539 7 1 2 53721 58223
0 35540 5 1 1 35539
0 35541 7 2 2 35538 35540
0 35542 5 5 1 67291
0 35543 7 1 2 51797 67292
0 35544 5 3 1 35543
0 35545 7 2 2 42890 67298
0 35546 7 1 2 40688 51979
0 35547 7 1 2 67301 35546
0 35548 5 1 1 35547
0 35549 7 1 2 35536 35548
0 35550 5 1 1 35549
0 35551 7 1 2 44830 35550
0 35552 5 1 1 35551
0 35553 7 1 2 53297 50097
0 35554 7 1 2 67302 35553
0 35555 5 1 1 35554
0 35556 7 1 2 35552 35555
0 35557 5 1 1 35556
0 35558 7 1 2 53661 35557
0 35559 5 1 1 35558
0 35560 7 1 2 57491 57361
0 35561 7 1 2 67299 35560
0 35562 5 1 1 35561
0 35563 7 1 2 35559 35562
0 35564 5 1 1 35563
0 35565 7 1 2 44138 35564
0 35566 5 1 1 35565
0 35567 7 1 2 64746 59128
0 35568 5 1 1 35567
0 35569 7 1 2 63202 67150
0 35570 5 1 1 35569
0 35571 7 1 2 49167 66627
0 35572 5 1 1 35571
0 35573 7 1 2 35570 35572
0 35574 7 1 2 35568 35573
0 35575 5 1 1 35574
0 35576 7 1 2 49866 35575
0 35577 5 1 1 35576
0 35578 7 2 2 50207 46768
0 35579 7 1 2 66265 60534
0 35580 5 1 1 35579
0 35581 7 1 2 66804 35580
0 35582 5 1 1 35581
0 35583 7 1 2 54281 35582
0 35584 5 1 1 35583
0 35585 7 1 2 55303 63661
0 35586 5 1 1 35585
0 35587 7 1 2 35584 35586
0 35588 5 1 1 35587
0 35589 7 1 2 67303 35588
0 35590 5 1 1 35589
0 35591 7 1 2 35577 35590
0 35592 5 1 1 35591
0 35593 7 1 2 43967 35592
0 35594 5 1 1 35593
0 35595 7 1 2 67304 60045
0 35596 7 1 2 56921 35595
0 35597 5 1 1 35596
0 35598 7 1 2 35594 35597
0 35599 5 1 1 35598
0 35600 7 1 2 45524 35599
0 35601 5 1 1 35600
0 35602 7 1 2 33457 57309
0 35603 5 1 1 35602
0 35604 7 1 2 54627 35603
0 35605 5 1 1 35604
0 35606 7 1 2 52137 57778
0 35607 5 1 1 35606
0 35608 7 1 2 35605 35607
0 35609 5 1 1 35608
0 35610 7 1 2 51462 67300
0 35611 7 1 2 35609 35610
0 35612 5 1 1 35611
0 35613 7 1 2 35601 35612
0 35614 7 1 2 35566 35613
0 35615 5 1 1 35614
0 35616 7 1 2 45126 35615
0 35617 5 1 1 35616
0 35618 7 1 2 59966 63329
0 35619 5 1 1 35618
0 35620 7 2 2 40121 45127
0 35621 7 1 2 66630 67305
0 35622 5 1 1 35621
0 35623 7 1 2 35619 35622
0 35624 5 1 1 35623
0 35625 7 1 2 49230 35624
0 35626 5 1 1 35625
0 35627 7 1 2 59366 64462
0 35628 5 1 1 35627
0 35629 7 1 2 63256 35628
0 35630 5 1 1 35629
0 35631 7 1 2 43156 65555
0 35632 7 1 2 35630 35631
0 35633 5 1 1 35632
0 35634 7 1 2 63488 57814
0 35635 7 1 2 63633 35634
0 35636 5 1 1 35635
0 35637 7 1 2 35633 35636
0 35638 7 1 2 35626 35637
0 35639 5 1 1 35638
0 35640 7 1 2 43968 35639
0 35641 5 1 1 35640
0 35642 7 1 2 62993 67306
0 35643 7 1 2 53617 35642
0 35644 7 1 2 52145 35643
0 35645 5 1 1 35644
0 35646 7 1 2 35641 35645
0 35647 5 1 1 35646
0 35648 7 1 2 46911 35647
0 35649 5 1 1 35648
0 35650 7 1 2 42721 64067
0 35651 5 1 1 35650
0 35652 7 1 2 19264 35651
0 35653 5 2 1 35652
0 35654 7 1 2 44139 67307
0 35655 5 1 1 35654
0 35656 7 1 2 54282 49343
0 35657 5 1 1 35656
0 35658 7 1 2 35655 35657
0 35659 5 4 1 35658
0 35660 7 1 2 43969 54987
0 35661 7 1 2 61657 35660
0 35662 7 1 2 52553 35661
0 35663 7 1 2 67309 35662
0 35664 5 1 1 35663
0 35665 7 1 2 35649 35664
0 35666 5 1 1 35665
0 35667 7 1 2 45525 35666
0 35668 5 1 1 35667
0 35669 7 2 2 50957 67310
0 35670 7 1 2 50386 67313
0 35671 5 1 1 35670
0 35672 7 1 2 65615 51235
0 35673 7 1 2 61184 35672
0 35674 5 1 1 35673
0 35675 7 1 2 35671 35674
0 35676 5 1 1 35675
0 35677 7 1 2 47664 35676
0 35678 5 1 1 35677
0 35679 7 1 2 56264 67314
0 35680 5 1 1 35679
0 35681 7 1 2 50958 67308
0 35682 5 1 1 35681
0 35683 7 1 2 65616 51239
0 35684 5 1 1 35683
0 35685 7 1 2 35682 35684
0 35686 5 1 1 35685
0 35687 7 1 2 44140 35686
0 35688 5 1 1 35687
0 35689 7 1 2 67093 64762
0 35690 5 1 1 35689
0 35691 7 1 2 35688 35690
0 35692 5 1 1 35691
0 35693 7 1 2 49893 35692
0 35694 5 1 1 35693
0 35695 7 1 2 35680 35694
0 35696 7 1 2 35678 35695
0 35697 5 1 1 35696
0 35698 7 1 2 43157 59939
0 35699 7 1 2 35697 35698
0 35700 5 1 1 35699
0 35701 7 1 2 35668 35700
0 35702 7 1 2 35617 35701
0 35703 5 1 1 35702
0 35704 7 1 2 44299 35703
0 35705 5 1 1 35704
0 35706 7 3 2 59367 55304
0 35707 7 1 2 41153 67315
0 35708 5 1 1 35707
0 35709 7 1 2 63967 35708
0 35710 5 1 1 35709
0 35711 7 1 2 44300 35710
0 35712 5 1 1 35711
0 35713 7 1 2 66483 35712
0 35714 5 1 1 35713
0 35715 7 1 2 40122 35714
0 35716 5 1 1 35715
0 35717 7 2 2 48971 63268
0 35718 5 1 1 67318
0 35719 7 1 2 57326 67319
0 35720 5 1 1 35719
0 35721 7 1 2 35716 35720
0 35722 5 1 1 35721
0 35723 7 1 2 45349 35722
0 35724 5 1 1 35723
0 35725 7 1 2 63640 67316
0 35726 5 1 1 35725
0 35727 7 1 2 35724 35726
0 35728 5 1 1 35727
0 35729 7 1 2 43158 35728
0 35730 5 1 1 35729
0 35731 7 1 2 58575 50541
0 35732 7 1 2 67222 35731
0 35733 5 1 1 35732
0 35734 7 1 2 35730 35733
0 35735 5 1 1 35734
0 35736 7 1 2 47823 35735
0 35737 5 1 1 35736
0 35738 7 1 2 50851 52645
0 35739 7 1 2 67035 35738
0 35740 5 1 1 35739
0 35741 7 1 2 35718 35740
0 35742 5 1 1 35741
0 35743 7 1 2 44141 35742
0 35744 5 1 1 35743
0 35745 7 1 2 50852 52940
0 35746 7 1 2 63294 35745
0 35747 5 1 1 35746
0 35748 7 1 2 35744 35747
0 35749 5 1 1 35748
0 35750 7 1 2 43159 50208
0 35751 7 1 2 35749 35750
0 35752 5 1 1 35751
0 35753 7 1 2 35737 35752
0 35754 5 1 1 35753
0 35755 7 1 2 65635 35754
0 35756 5 1 1 35755
0 35757 7 1 2 49894 58918
0 35758 7 1 2 49251 35757
0 35759 5 1 1 35758
0 35760 7 1 2 40513 58710
0 35761 5 1 1 35760
0 35762 7 1 2 58903 59620
0 35763 7 1 2 35761 35762
0 35764 5 1 1 35763
0 35765 7 1 2 35759 35764
0 35766 5 1 1 35765
0 35767 7 1 2 43040 35766
0 35768 5 1 1 35767
0 35769 7 1 2 67036 62196
0 35770 7 1 2 58705 35769
0 35771 5 1 1 35770
0 35772 7 1 2 35768 35771
0 35773 5 1 1 35772
0 35774 7 1 2 42186 35773
0 35775 5 1 1 35774
0 35776 7 1 2 58224 61371
0 35777 7 1 2 66808 35776
0 35778 5 1 1 35777
0 35779 7 1 2 43160 51076
0 35780 7 1 2 63269 35779
0 35781 7 1 2 59621 35780
0 35782 5 1 1 35781
0 35783 7 1 2 35778 35782
0 35784 5 1 1 35783
0 35785 7 1 2 47355 35784
0 35786 5 1 1 35785
0 35787 7 1 2 50912 62783
0 35788 7 1 2 59622 35787
0 35789 5 1 1 35788
0 35790 7 1 2 57666 58116
0 35791 7 1 2 66809 35790
0 35792 5 1 1 35791
0 35793 7 1 2 35789 35792
0 35794 5 1 1 35793
0 35795 7 1 2 47665 35794
0 35796 5 1 1 35795
0 35797 7 1 2 35786 35796
0 35798 7 1 2 35775 35797
0 35799 5 1 1 35798
0 35800 7 1 2 43970 35799
0 35801 5 1 1 35800
0 35802 7 1 2 35756 35801
0 35803 5 1 1 35802
0 35804 7 1 2 54369 35803
0 35805 5 1 1 35804
0 35806 7 1 2 62142 49252
0 35807 5 1 1 35806
0 35808 7 1 2 56684 59371
0 35809 5 1 1 35808
0 35810 7 1 2 35807 35809
0 35811 5 1 1 35810
0 35812 7 1 2 51858 35811
0 35813 5 1 1 35812
0 35814 7 2 2 40514 51568
0 35815 7 1 2 45128 56786
0 35816 7 1 2 52727 35815
0 35817 7 1 2 67320 35816
0 35818 5 1 1 35817
0 35819 7 1 2 35813 35818
0 35820 5 1 1 35819
0 35821 7 1 2 43041 35820
0 35822 5 1 1 35821
0 35823 7 1 2 57488 59351
0 35824 7 1 2 55692 35823
0 35825 5 1 1 35824
0 35826 7 1 2 35822 35825
0 35827 5 1 1 35826
0 35828 7 1 2 54283 35827
0 35829 5 1 1 35828
0 35830 7 1 2 40123 67317
0 35831 5 1 1 35830
0 35832 7 1 2 63968 35831
0 35833 5 1 1 35832
0 35834 7 1 2 41539 51859
0 35835 7 1 2 57688 35834
0 35836 7 1 2 35833 35835
0 35837 5 1 1 35836
0 35838 7 1 2 35829 35837
0 35839 5 1 1 35838
0 35840 7 1 2 44301 35839
0 35841 5 1 1 35840
0 35842 7 1 2 43042 51860
0 35843 7 1 2 59094 35842
0 35844 7 1 2 67311 35843
0 35845 5 1 1 35844
0 35846 7 1 2 35841 35845
0 35847 5 1 1 35846
0 35848 7 1 2 43971 35847
0 35849 5 1 1 35848
0 35850 7 1 2 44977 65715
0 35851 7 1 2 48595 35850
0 35852 7 1 2 57140 35851
0 35853 7 1 2 67246 35852
0 35854 5 1 1 35853
0 35855 7 1 2 35849 35854
0 35856 5 1 1 35855
0 35857 7 1 2 46863 35856
0 35858 5 1 1 35857
0 35859 7 1 2 43784 35530
0 35860 5 1 1 35859
0 35861 7 1 2 51160 35860
0 35862 5 1 1 35861
0 35863 7 1 2 49867 60431
0 35864 5 2 1 35863
0 35865 7 1 2 50959 67322
0 35866 5 2 1 35865
0 35867 7 1 2 35862 67324
0 35868 5 1 1 35867
0 35869 7 1 2 67312 35868
0 35870 5 1 1 35869
0 35871 7 1 2 55471 49145
0 35872 7 1 2 61378 35871
0 35873 5 1 1 35872
0 35874 7 1 2 35870 35873
0 35875 5 1 1 35874
0 35876 7 1 2 64982 35875
0 35877 5 1 1 35876
0 35878 7 1 2 35858 35877
0 35879 7 1 2 35805 35878
0 35880 7 1 2 35705 35879
0 35881 5 1 1 35880
0 35882 7 1 2 67279 35881
0 35883 5 1 1 35882
0 35884 7 9 2 46524 43281
0 35885 7 1 2 40515 12424
0 35886 5 7 1 35885
0 35887 7 2 2 59181 67335
0 35888 7 1 2 44831 63156
0 35889 7 1 2 67342 35888
0 35890 5 1 1 35889
0 35891 7 1 2 50195 58084
0 35892 5 4 1 35891
0 35893 7 1 2 51161 67344
0 35894 5 2 1 35893
0 35895 7 1 2 67325 67348
0 35896 5 1 1 35895
0 35897 7 1 2 59295 50945
0 35898 7 1 2 35896 35897
0 35899 5 1 1 35898
0 35900 7 1 2 35890 35899
0 35901 5 1 1 35900
0 35902 7 1 2 49231 35901
0 35903 5 1 1 35902
0 35904 7 2 2 55124 59397
0 35905 7 1 2 43457 51408
0 35906 5 1 1 35905
0 35907 7 1 2 56872 35906
0 35908 5 1 1 35907
0 35909 7 1 2 60424 35908
0 35910 5 1 1 35909
0 35911 7 1 2 47741 50815
0 35912 5 1 1 35911
0 35913 7 1 2 47666 51409
0 35914 5 1 1 35913
0 35915 7 1 2 43458 56870
0 35916 5 1 1 35915
0 35917 7 1 2 35914 35916
0 35918 5 1 1 35917
0 35919 7 1 2 46852 35918
0 35920 5 1 1 35919
0 35921 7 1 2 35912 35920
0 35922 7 1 2 35910 35921
0 35923 5 1 1 35922
0 35924 7 1 2 42187 35923
0 35925 5 1 1 35924
0 35926 7 1 2 60979 50869
0 35927 5 1 1 35926
0 35928 7 1 2 35925 35927
0 35929 5 1 1 35928
0 35930 7 1 2 67350 35929
0 35931 5 1 1 35930
0 35932 7 1 2 60023 56963
0 35933 7 1 2 67343 35932
0 35934 5 1 1 35933
0 35935 7 1 2 35931 35934
0 35936 7 1 2 35903 35935
0 35937 5 1 1 35936
0 35938 7 1 2 46442 35937
0 35939 5 1 1 35938
0 35940 7 1 2 50703 57874
0 35941 5 1 1 35940
0 35942 7 1 2 53520 62915
0 35943 5 1 1 35942
0 35944 7 1 2 35941 35943
0 35945 5 1 1 35944
0 35946 7 1 2 46638 35945
0 35947 5 1 1 35946
0 35948 7 1 2 35939 35947
0 35949 5 1 1 35948
0 35950 7 1 2 45996 35949
0 35951 5 1 1 35950
0 35952 7 2 2 40689 54045
0 35953 5 1 1 67352
0 35954 7 1 2 67349 35953
0 35955 5 1 1 35954
0 35956 7 1 2 67351 35955
0 35957 5 1 1 35956
0 35958 7 3 2 43043 67336
0 35959 7 1 2 63767 53268
0 35960 7 1 2 67354 35959
0 35961 5 1 1 35960
0 35962 7 1 2 35957 35961
0 35963 5 1 1 35962
0 35964 7 1 2 56630 51401
0 35965 7 1 2 35963 35964
0 35966 5 1 1 35965
0 35967 7 1 2 35951 35966
0 35968 5 1 1 35967
0 35969 7 1 2 67326 35968
0 35970 5 1 1 35969
0 35971 7 1 2 51088 59356
0 35972 5 1 1 35971
0 35973 7 1 2 65636 49232
0 35974 7 1 2 67345 35973
0 35975 5 1 1 35974
0 35976 7 1 2 35972 35975
0 35977 5 1 1 35976
0 35978 7 1 2 59296 35977
0 35979 5 1 1 35978
0 35980 7 1 2 49270 63768
0 35981 7 1 2 67355 35980
0 35982 5 1 1 35981
0 35983 7 1 2 35979 35982
0 35984 5 1 1 35983
0 35985 7 9 2 46443 67327
0 35986 7 1 2 67357 56478
0 35987 7 1 2 35984 35986
0 35988 5 1 1 35987
0 35989 7 1 2 35970 35988
0 35990 7 1 2 35883 35989
0 35991 5 1 1 35990
0 35992 7 1 2 46599 35991
0 35993 5 1 1 35992
0 35994 7 17 2 46530 64695
0 35995 7 1 2 57792 5082
0 35996 5 3 1 35995
0 35997 7 1 2 45997 67383
0 35998 5 1 1 35997
0 35999 7 1 2 65712 58793
0 36000 5 1 1 35999
0 36001 7 1 2 35998 36000
0 36002 5 2 1 36001
0 36003 7 1 2 47742 50882
0 36004 5 1 1 36003
0 36005 7 1 2 44558 65044
0 36006 5 1 1 36005
0 36007 7 1 2 42188 58314
0 36008 7 1 2 36006 36007
0 36009 5 1 1 36008
0 36010 7 1 2 36004 36009
0 36011 5 1 1 36010
0 36012 7 1 2 43785 36011
0 36013 5 1 1 36012
0 36014 7 1 2 43598 64829
0 36015 7 1 2 55841 36014
0 36016 5 2 1 36015
0 36017 7 1 2 36013 67388
0 36018 5 1 1 36017
0 36019 7 1 2 67386 36018
0 36020 5 1 1 36019
0 36021 7 1 2 65543 57489
0 36022 5 1 1 36021
0 36023 7 1 2 58794 57004
0 36024 5 1 1 36023
0 36025 7 1 2 36022 36024
0 36026 5 1 1 36025
0 36027 7 1 2 40516 36026
0 36028 7 1 2 65059 36027
0 36029 5 1 1 36028
0 36030 7 1 2 36020 36029
0 36031 5 1 1 36030
0 36032 7 1 2 67366 36031
0 36033 5 1 1 36032
0 36034 7 2 2 44832 49752
0 36035 7 1 2 56664 67390
0 36036 5 1 1 36035
0 36037 7 1 2 40690 49381
0 36038 7 1 2 67238 36037
0 36039 5 1 1 36038
0 36040 7 1 2 36036 36039
0 36041 5 1 1 36040
0 36042 7 2 2 43282 58555
0 36043 7 1 2 45998 67392
0 36044 7 1 2 36041 36043
0 36045 5 1 1 36044
0 36046 7 1 2 36033 36045
0 36047 5 1 1 36046
0 36048 7 1 2 45129 36047
0 36049 5 1 1 36048
0 36050 7 1 2 47298 47251
0 36051 5 1 1 36050
0 36052 7 2 2 58225 36051
0 36053 5 1 1 67394
0 36054 7 1 2 42722 67395
0 36055 5 1 1 36054
0 36056 7 1 2 45999 55913
0 36057 5 1 1 36056
0 36058 7 1 2 45350 36057
0 36059 7 1 2 36055 36058
0 36060 5 1 1 36059
0 36061 7 1 2 52500 61375
0 36062 5 1 1 36061
0 36063 7 5 2 58374 53183
0 36064 7 1 2 61212 67396
0 36065 5 2 1 36064
0 36066 7 1 2 36062 67401
0 36067 7 1 2 36060 36066
0 36068 5 1 1 36067
0 36069 7 1 2 49618 36068
0 36070 5 1 1 36069
0 36071 7 2 2 43599 64891
0 36072 5 2 1 67403
0 36073 7 1 2 22987 67405
0 36074 5 1 1 36073
0 36075 7 1 2 42189 64796
0 36076 7 1 2 36074 36075
0 36077 5 1 1 36076
0 36078 7 1 2 36070 36077
0 36079 5 1 1 36078
0 36080 7 1 2 43161 67367
0 36081 7 1 2 64960 36080
0 36082 7 1 2 36079 36081
0 36083 5 1 1 36082
0 36084 7 1 2 36049 36083
0 36085 5 1 1 36084
0 36086 7 1 2 46525 36085
0 36087 5 1 1 36086
0 36088 7 1 2 50209 47900
0 36089 5 1 1 36088
0 36090 7 1 2 49895 36089
0 36091 5 1 1 36090
0 36092 7 1 2 45526 36091
0 36093 5 1 1 36092
0 36094 7 2 2 58092 36093
0 36095 5 4 1 67407
0 36096 7 1 2 65571 67409
0 36097 5 1 1 36096
0 36098 7 1 2 53300 67408
0 36099 5 1 1 36098
0 36100 7 1 2 55917 56210
0 36101 5 1 1 36100
0 36102 7 1 2 53298 50314
0 36103 7 1 2 36101 36102
0 36104 5 1 1 36103
0 36105 7 1 2 40691 54288
0 36106 7 1 2 36104 36105
0 36107 7 1 2 36099 36106
0 36108 5 1 1 36107
0 36109 7 1 2 36097 36108
0 36110 5 1 1 36109
0 36111 7 1 2 56574 60405
0 36112 7 1 2 67368 36111
0 36113 7 1 2 36110 36112
0 36114 5 1 1 36113
0 36115 7 1 2 36087 36114
0 36116 5 1 1 36115
0 36117 7 1 2 44302 36116
0 36118 5 1 1 36117
0 36119 7 2 2 57392 56619
0 36120 7 1 2 58448 58460
0 36121 7 1 2 58444 36120
0 36122 5 1 1 36121
0 36123 7 1 2 40517 36122
0 36124 5 1 1 36123
0 36125 7 1 2 58402 36124
0 36126 5 1 1 36125
0 36127 7 1 2 42723 36126
0 36128 5 1 1 36127
0 36129 7 1 2 67402 36128
0 36130 5 1 1 36129
0 36131 7 1 2 67413 36130
0 36132 5 1 1 36131
0 36133 7 4 2 55599 60516
0 36134 5 2 1 67415
0 36135 7 1 2 42724 67410
0 36136 5 1 1 36135
0 36137 7 1 2 7902 36136
0 36138 5 1 1 36137
0 36139 7 1 2 67416 36138
0 36140 5 1 1 36139
0 36141 7 1 2 36132 36140
0 36142 5 1 1 36141
0 36143 7 1 2 45130 36142
0 36144 5 1 1 36143
0 36145 7 2 2 41997 67417
0 36146 5 1 1 67421
0 36147 7 1 2 54704 67414
0 36148 5 1 1 36147
0 36149 7 1 2 36146 36148
0 36150 5 2 1 36149
0 36151 7 1 2 42190 67423
0 36152 5 1 1 36151
0 36153 7 1 2 47432 67422
0 36154 5 1 1 36153
0 36155 7 1 2 36152 36154
0 36156 5 1 1 36155
0 36157 7 1 2 45131 36156
0 36158 5 1 1 36157
0 36159 7 1 2 41823 61339
0 36160 7 1 2 67384 36159
0 36161 5 1 1 36160
0 36162 7 1 2 36158 36161
0 36163 5 1 1 36162
0 36164 7 1 2 46000 36163
0 36165 5 1 1 36164
0 36166 7 1 2 58576 66316
0 36167 7 1 2 67016 36166
0 36168 5 1 1 36167
0 36169 7 1 2 36165 36168
0 36170 5 1 1 36169
0 36171 7 1 2 49896 36170
0 36172 5 1 1 36171
0 36173 7 3 2 64645 55648
0 36174 7 1 2 65184 67425
0 36175 5 1 1 36174
0 36176 7 1 2 40518 67426
0 36177 5 1 1 36176
0 36178 7 1 2 45132 66941
0 36179 7 1 2 58075 36178
0 36180 5 1 1 36179
0 36181 7 1 2 36177 36180
0 36182 5 1 1 36181
0 36183 7 1 2 52816 36182
0 36184 5 1 1 36183
0 36185 7 1 2 45351 67427
0 36186 5 1 1 36185
0 36187 7 1 2 43600 63974
0 36188 7 1 2 60780 36187
0 36189 7 1 2 62642 36188
0 36190 5 1 1 36189
0 36191 7 1 2 36186 36190
0 36192 5 1 1 36191
0 36193 7 1 2 40519 36192
0 36194 5 1 1 36193
0 36195 7 1 2 36184 36194
0 36196 7 1 2 36175 36195
0 36197 5 1 1 36196
0 36198 7 1 2 43162 36197
0 36199 5 1 1 36198
0 36200 7 2 2 57278 67411
0 36201 7 1 2 63238 64964
0 36202 7 1 2 67428 36201
0 36203 5 1 1 36202
0 36204 7 1 2 36199 36203
0 36205 5 1 1 36204
0 36206 7 1 2 58061 36205
0 36207 5 1 1 36206
0 36208 7 1 2 40300 63383
0 36209 5 1 1 36208
0 36210 7 1 2 46934 36209
0 36211 5 3 1 36210
0 36212 7 1 2 52501 60406
0 36213 7 1 2 67385 36212
0 36214 7 1 2 67430 36213
0 36215 5 1 1 36214
0 36216 7 1 2 36207 36215
0 36217 7 1 2 36172 36216
0 36218 7 1 2 36144 36217
0 36219 5 1 1 36218
0 36220 7 1 2 41037 67369
0 36221 7 1 2 36219 36220
0 36222 5 1 1 36221
0 36223 7 3 2 43786 65095
0 36224 5 1 1 67433
0 36225 7 1 2 61293 67434
0 36226 5 1 1 36225
0 36227 7 1 2 52375 60471
0 36228 5 1 1 36227
0 36229 7 1 2 36226 36228
0 36230 5 1 1 36229
0 36231 7 1 2 43601 36230
0 36232 5 1 1 36231
0 36233 7 2 2 43271 47153
0 36234 7 1 2 61257 67436
0 36235 5 1 1 36234
0 36236 7 1 2 36232 36235
0 36237 5 1 1 36236
0 36238 7 1 2 67387 36237
0 36239 5 1 1 36238
0 36240 7 1 2 62524 53090
0 36241 7 1 2 63011 36240
0 36242 5 1 1 36241
0 36243 7 1 2 67419 36242
0 36244 5 1 1 36243
0 36245 7 1 2 54756 36244
0 36246 5 1 1 36245
0 36247 7 1 2 47131 63012
0 36248 7 1 2 61152 36247
0 36249 5 1 1 36248
0 36250 7 1 2 67420 36249
0 36251 5 1 1 36250
0 36252 7 1 2 43787 51893
0 36253 7 1 2 36251 36252
0 36254 5 1 1 36253
0 36255 7 1 2 36246 36254
0 36256 5 1 1 36255
0 36257 7 1 2 64715 36256
0 36258 5 1 1 36257
0 36259 7 1 2 36239 36258
0 36260 5 1 1 36259
0 36261 7 1 2 47356 36260
0 36262 5 1 1 36261
0 36263 7 1 2 61213 67424
0 36264 5 1 1 36263
0 36265 7 1 2 46001 67418
0 36266 5 1 1 36265
0 36267 7 1 2 58062 58751
0 36268 7 1 2 63836 36267
0 36269 5 1 1 36268
0 36270 7 1 2 36266 36269
0 36271 5 1 1 36270
0 36272 7 1 2 42191 66180
0 36273 7 1 2 36271 36272
0 36274 5 1 1 36273
0 36275 7 1 2 36264 36274
0 36276 5 1 1 36275
0 36277 7 1 2 55125 36276
0 36278 5 1 1 36277
0 36279 7 1 2 61294 61278
0 36280 5 1 1 36279
0 36281 7 1 2 61344 36280
0 36282 5 1 1 36281
0 36283 7 1 2 47433 36282
0 36284 5 1 1 36283
0 36285 7 1 2 36284 61255
0 36286 5 1 1 36285
0 36287 7 1 2 40692 66631
0 36288 5 1 1 36287
0 36289 7 1 2 54370 63338
0 36290 5 1 1 36289
0 36291 7 1 2 36288 36290
0 36292 5 1 1 36291
0 36293 7 1 2 36286 36292
0 36294 5 1 1 36293
0 36295 7 1 2 36278 36294
0 36296 5 1 1 36295
0 36297 7 1 2 47667 36296
0 36298 5 1 1 36297
0 36299 7 1 2 36262 36298
0 36300 5 1 1 36299
0 36301 7 1 2 67370 36300
0 36302 5 1 1 36301
0 36303 7 1 2 49619 66184
0 36304 7 2 2 53662 67328
0 36305 7 1 2 64416 67438
0 36306 7 1 2 36303 36305
0 36307 7 1 2 61784 36306
0 36308 5 1 1 36307
0 36309 7 1 2 36302 36308
0 36310 7 1 2 36222 36309
0 36311 7 1 2 36118 36310
0 36312 5 1 1 36311
0 36313 7 1 2 49233 36312
0 36314 5 1 1 36313
0 36315 7 2 2 67356 67358
0 36316 7 1 2 51569 64417
0 36317 7 2 2 67440 36316
0 36318 5 1 1 67442
0 36319 7 1 2 40693 67443
0 36320 5 1 1 36319
0 36321 7 1 2 20002 20376
0 36322 5 1 1 36321
0 36323 7 1 2 59518 36322
0 36324 5 2 1 36323
0 36325 7 1 2 65041 58919
0 36326 5 1 1 36325
0 36327 7 3 2 43163 55143
0 36328 7 1 2 55126 67446
0 36329 5 1 1 36328
0 36330 7 1 2 36326 36329
0 36331 5 1 1 36330
0 36332 7 1 2 46526 36331
0 36333 5 1 1 36332
0 36334 7 1 2 63561 36333
0 36335 5 1 1 36334
0 36336 7 1 2 57507 36335
0 36337 5 1 1 36336
0 36338 7 1 2 67444 36337
0 36339 5 1 1 36338
0 36340 7 1 2 41272 36339
0 36341 5 1 1 36340
0 36342 7 1 2 47299 59147
0 36343 5 1 1 36342
0 36344 7 1 2 46639 67447
0 36345 5 1 1 36344
0 36346 7 1 2 36343 36345
0 36347 5 1 1 36346
0 36348 7 1 2 59398 36347
0 36349 5 1 1 36348
0 36350 7 3 2 53670 59126
0 36351 7 1 2 40301 67449
0 36352 5 1 1 36351
0 36353 7 1 2 36349 36352
0 36354 5 1 1 36353
0 36355 7 1 2 43272 36354
0 36356 5 1 1 36355
0 36357 7 1 2 36341 36356
0 36358 5 1 1 36357
0 36359 7 1 2 45527 36358
0 36360 5 1 1 36359
0 36361 7 1 2 49714 63790
0 36362 5 1 1 36361
0 36363 7 1 2 51570 57397
0 36364 5 1 1 36363
0 36365 7 1 2 36362 36364
0 36366 5 1 1 36365
0 36367 7 1 2 55127 36366
0 36368 5 1 1 36367
0 36369 7 1 2 45133 63630
0 36370 7 1 2 57705 63204
0 36371 7 1 2 36369 36370
0 36372 5 1 1 36371
0 36373 7 1 2 36368 36372
0 36374 5 1 1 36373
0 36375 7 1 2 47132 36374
0 36376 5 1 1 36375
0 36377 7 1 2 44142 54242
0 36378 7 1 2 59664 36377
0 36379 7 1 2 67030 36378
0 36380 5 1 1 36379
0 36381 7 1 2 36376 36380
0 36382 7 1 2 36360 36381
0 36383 5 1 1 36382
0 36384 7 1 2 40520 36383
0 36385 5 1 1 36384
0 36386 7 1 2 46895 46640
0 36387 7 1 2 66242 36386
0 36388 5 2 1 36387
0 36389 7 2 2 59519 62881
0 36390 7 1 2 57988 67454
0 36391 5 2 1 36390
0 36392 7 7 2 59520 61435
0 36393 5 1 1 67458
0 36394 7 1 2 45352 67459
0 36395 5 2 1 36394
0 36396 7 1 2 63796 32246
0 36397 5 1 1 36396
0 36398 7 2 2 55128 36397
0 36399 5 1 1 67467
0 36400 7 1 2 41273 67468
0 36401 5 1 1 36400
0 36402 7 1 2 67465 36401
0 36403 5 1 1 36402
0 36404 7 1 2 40124 36403
0 36405 5 1 1 36404
0 36406 7 1 2 67456 36405
0 36407 5 1 1 36406
0 36408 7 1 2 41154 36407
0 36409 5 1 1 36408
0 36410 7 1 2 67452 36409
0 36411 5 1 1 36410
0 36412 7 1 2 51861 36411
0 36413 5 1 1 36412
0 36414 7 1 2 62368 59435
0 36415 7 1 2 63180 36414
0 36416 5 2 1 36415
0 36417 7 1 2 45134 58610
0 36418 7 3 2 61871 36417
0 36419 7 1 2 56594 67228
0 36420 7 1 2 67471 36419
0 36421 5 1 1 36420
0 36422 7 1 2 55129 47133
0 36423 7 1 2 63811 36422
0 36424 5 1 1 36423
0 36425 7 1 2 36421 36424
0 36426 5 1 1 36425
0 36427 7 1 2 40521 36426
0 36428 5 1 1 36427
0 36429 7 1 2 67469 36428
0 36430 5 1 1 36429
0 36431 7 1 2 52112 36430
0 36432 5 1 1 36431
0 36433 7 1 2 52332 47072
0 36434 7 1 2 63791 36433
0 36435 5 1 1 36434
0 36436 7 1 2 63044 55779
0 36437 7 1 2 65782 36436
0 36438 5 1 1 36437
0 36439 7 1 2 36435 36438
0 36440 5 1 1 36439
0 36441 7 1 2 55130 36440
0 36442 5 1 1 36441
0 36443 7 1 2 59288 67455
0 36444 5 1 1 36443
0 36445 7 1 2 45135 62023
0 36446 7 1 2 60851 36445
0 36447 7 1 2 66440 36446
0 36448 5 1 1 36447
0 36449 7 1 2 36444 36448
0 36450 5 1 1 36449
0 36451 7 1 2 40522 36450
0 36452 5 1 1 36451
0 36453 7 1 2 36442 36452
0 36454 5 1 1 36453
0 36455 7 1 2 47499 36454
0 36456 5 1 1 36455
0 36457 7 1 2 43972 36456
0 36458 7 1 2 36432 36457
0 36459 7 1 2 36413 36458
0 36460 7 1 2 36385 36459
0 36461 5 1 1 36460
0 36462 7 1 2 67460 61397
0 36463 5 1 1 36462
0 36464 7 1 2 44559 65037
0 36465 5 1 1 36464
0 36466 7 1 2 47668 50241
0 36467 7 2 2 36465 36466
0 36468 5 1 1 67474
0 36469 7 1 2 40125 48796
0 36470 5 1 1 36469
0 36471 7 1 2 60425 58111
0 36472 7 1 2 36470 36471
0 36473 5 1 1 36472
0 36474 7 1 2 36468 36473
0 36475 5 2 1 36474
0 36476 7 1 2 57815 67476
0 36477 5 1 1 36476
0 36478 7 1 2 65335 59399
0 36479 7 1 2 61785 36478
0 36480 5 1 1 36479
0 36481 7 1 2 36477 36480
0 36482 5 1 1 36481
0 36483 7 1 2 43788 36482
0 36484 5 1 1 36483
0 36485 7 2 2 66266 62909
0 36486 5 1 1 67478
0 36487 7 1 2 57829 36486
0 36488 5 1 1 36487
0 36489 7 1 2 53722 67404
0 36490 7 1 2 36488 36489
0 36491 5 1 1 36490
0 36492 7 1 2 36484 36491
0 36493 5 1 1 36492
0 36494 7 1 2 60300 36493
0 36495 5 1 1 36494
0 36496 7 1 2 36463 36495
0 36497 5 1 1 36496
0 36498 7 1 2 42192 36497
0 36499 5 1 1 36498
0 36500 7 1 2 65783 57706
0 36501 5 1 1 36500
0 36502 7 1 2 63797 36501
0 36503 5 1 1 36502
0 36504 7 1 2 47669 36503
0 36505 5 1 1 36504
0 36506 7 2 2 59933 62977
0 36507 7 1 2 63144 67480
0 36508 5 1 1 36507
0 36509 7 1 2 63798 36508
0 36510 5 1 1 36509
0 36511 7 1 2 42193 36510
0 36512 5 1 1 36511
0 36513 7 1 2 36505 36512
0 36514 5 1 1 36513
0 36515 7 1 2 43789 36514
0 36516 5 1 1 36515
0 36517 7 1 2 67481 67321
0 36518 5 1 1 36517
0 36519 7 1 2 63799 36518
0 36520 5 1 1 36519
0 36521 7 1 2 54757 36520
0 36522 5 1 1 36521
0 36523 7 1 2 36516 36522
0 36524 5 1 1 36523
0 36525 7 1 2 47357 36524
0 36526 5 1 1 36525
0 36527 7 1 2 63002 67397
0 36528 5 1 1 36527
0 36529 7 1 2 57279 60051
0 36530 7 1 2 58517 36529
0 36531 5 1 1 36530
0 36532 7 1 2 36528 36531
0 36533 5 1 1 36532
0 36534 7 1 2 43790 36533
0 36535 5 1 1 36534
0 36536 7 2 2 43602 62711
0 36537 7 1 2 67482 62981
0 36538 5 1 1 36537
0 36539 7 1 2 60517 60055
0 36540 5 1 1 36539
0 36541 7 1 2 36538 36540
0 36542 5 1 1 36541
0 36543 7 1 2 47434 36542
0 36544 5 1 1 36543
0 36545 7 1 2 47951 48329
0 36546 7 1 2 57384 36545
0 36547 5 2 1 36546
0 36548 7 1 2 36544 67484
0 36549 5 1 1 36548
0 36550 7 1 2 47154 36549
0 36551 5 1 1 36550
0 36552 7 1 2 58867 66879
0 36553 5 1 1 36552
0 36554 7 1 2 67485 36553
0 36555 5 1 1 36554
0 36556 7 1 2 47435 36555
0 36557 5 1 1 36556
0 36558 7 2 2 52339 57968
0 36559 7 1 2 59357 67486
0 36560 5 1 1 36559
0 36561 7 1 2 36557 36560
0 36562 5 1 1 36561
0 36563 7 1 2 47058 36562
0 36564 5 1 1 36563
0 36565 7 1 2 36551 36564
0 36566 7 1 2 36535 36565
0 36567 7 1 2 36526 36566
0 36568 5 1 1 36567
0 36569 7 1 2 55131 36568
0 36570 5 2 1 36569
0 36571 7 2 2 41998 67472
0 36572 7 1 2 51571 62786
0 36573 7 1 2 67490 36572
0 36574 5 1 1 36573
0 36575 7 1 2 36393 36574
0 36576 5 1 1 36575
0 36577 7 1 2 47670 36576
0 36578 5 1 1 36577
0 36579 7 1 2 66369 49256
0 36580 7 1 2 67491 36579
0 36581 5 1 1 36580
0 36582 7 1 2 36578 36581
0 36583 5 1 1 36582
0 36584 7 1 2 43791 36583
0 36585 5 1 1 36584
0 36586 7 2 2 65178 61258
0 36587 7 1 2 48086 67492
0 36588 5 1 1 36587
0 36589 7 1 2 67473 59027
0 36590 5 1 1 36589
0 36591 7 1 2 36588 36590
0 36592 5 1 1 36591
0 36593 7 1 2 47743 36592
0 36594 5 1 1 36593
0 36595 7 1 2 58749 67461
0 36596 5 1 1 36595
0 36597 7 1 2 36594 36596
0 36598 5 1 1 36597
0 36599 7 1 2 47358 36598
0 36600 5 1 1 36599
0 36601 7 1 2 40694 36600
0 36602 7 1 2 36585 36601
0 36603 7 1 2 67488 36602
0 36604 7 1 2 36499 36603
0 36605 5 1 1 36604
0 36606 7 1 2 67371 36605
0 36607 7 1 2 36461 36606
0 36608 5 1 1 36607
0 36609 7 1 2 36320 36608
0 36610 5 1 1 36609
0 36611 7 1 2 65556 36610
0 36612 5 1 1 36611
0 36613 7 1 2 44446 67462
0 36614 5 2 1 36613
0 36615 7 1 2 66258 62234
0 36616 5 1 1 36615
0 36617 7 1 2 67494 36616
0 36618 5 1 1 36617
0 36619 7 1 2 43603 36618
0 36620 5 1 1 36619
0 36621 7 1 2 44143 66256
0 36622 7 1 2 63051 36621
0 36623 5 1 1 36622
0 36624 7 1 2 67495 36623
0 36625 5 1 1 36624
0 36626 7 1 2 44560 36625
0 36627 5 1 1 36626
0 36628 7 1 2 36620 36627
0 36629 5 1 1 36628
0 36630 7 1 2 42194 36629
0 36631 5 1 1 36630
0 36632 7 1 2 66831 63631
0 36633 7 1 2 66371 36632
0 36634 5 1 1 36633
0 36635 7 1 2 36631 36634
0 36636 5 1 1 36635
0 36637 7 1 2 49719 36636
0 36638 5 1 1 36637
0 36639 7 1 2 66243 60017
0 36640 5 1 1 36639
0 36641 7 1 2 47359 67463
0 36642 5 1 1 36641
0 36643 7 1 2 40523 61631
0 36644 7 1 2 67479 36643
0 36645 5 1 1 36644
0 36646 7 1 2 36642 36645
0 36647 5 1 1 36646
0 36648 7 1 2 41999 36647
0 36649 5 1 1 36648
0 36650 7 1 2 36640 36649
0 36651 5 1 1 36650
0 36652 7 1 2 44561 36651
0 36653 5 1 1 36652
0 36654 7 2 2 50704 51311
0 36655 7 1 2 65179 63058
0 36656 7 1 2 67496 36655
0 36657 5 1 1 36656
0 36658 7 1 2 36653 36657
0 36659 5 1 1 36658
0 36660 7 1 2 43604 36659
0 36661 5 1 1 36660
0 36662 7 1 2 51372 58518
0 36663 7 1 2 67493 36662
0 36664 5 1 1 36663
0 36665 7 2 2 40302 50828
0 36666 5 3 1 67498
0 36667 7 1 2 65096 67500
0 36668 5 1 1 36667
0 36669 7 1 2 45528 62456
0 36670 5 1 1 36669
0 36671 7 1 2 36668 36670
0 36672 5 1 1 36671
0 36673 7 1 2 44447 36672
0 36674 5 1 1 36673
0 36675 7 1 2 43459 46818
0 36676 5 1 1 36675
0 36677 7 1 2 65038 36676
0 36678 5 1 1 36677
0 36679 7 1 2 47104 36678
0 36680 5 1 1 36679
0 36681 7 2 2 36674 36680
0 36682 5 1 1 67503
0 36683 7 1 2 36682 63818
0 36684 5 1 1 36683
0 36685 7 1 2 47602 61088
0 36686 5 1 1 36685
0 36687 7 1 2 67464 36686
0 36688 5 1 1 36687
0 36689 7 1 2 36684 36688
0 36690 5 1 1 36689
0 36691 7 1 2 43792 36690
0 36692 5 1 1 36691
0 36693 7 1 2 36664 36692
0 36694 7 1 2 36661 36693
0 36695 7 1 2 36638 36694
0 36696 7 1 2 67489 36695
0 36697 5 1 1 36696
0 36698 7 1 2 67372 36697
0 36699 5 1 1 36698
0 36700 7 1 2 36699 36318
0 36701 5 1 1 36700
0 36702 7 1 2 49965 36701
0 36703 5 1 1 36702
0 36704 7 1 2 60301 64115
0 36705 5 1 1 36704
0 36706 7 1 2 36399 36705
0 36707 5 1 1 36706
0 36708 7 1 2 41274 36707
0 36709 5 1 1 36708
0 36710 7 1 2 67466 36709
0 36711 5 1 1 36710
0 36712 7 1 2 40126 36711
0 36713 5 1 1 36712
0 36714 7 1 2 36713 67457
0 36715 5 1 1 36714
0 36716 7 1 2 41155 36715
0 36717 5 1 1 36716
0 36718 7 1 2 36717 67453
0 36719 5 1 1 36718
0 36720 7 1 2 51862 36719
0 36721 5 1 1 36720
0 36722 7 1 2 63307 67448
0 36723 5 1 1 36722
0 36724 7 1 2 53663 67043
0 36725 7 1 2 65042 36724
0 36726 5 1 1 36725
0 36727 7 1 2 36723 36726
0 36728 5 1 1 36727
0 36729 7 1 2 46527 36728
0 36730 5 1 1 36729
0 36731 7 1 2 43273 67450
0 36732 5 1 1 36731
0 36733 7 1 2 67445 36732
0 36734 7 1 2 36730 36733
0 36735 5 1 1 36734
0 36736 7 1 2 41275 36735
0 36737 5 1 1 36736
0 36738 7 1 2 57948 62982
0 36739 5 1 1 36738
0 36740 7 1 2 60518 64463
0 36741 5 1 1 36740
0 36742 7 1 2 36739 36741
0 36743 5 1 1 36742
0 36744 7 2 2 55132 36743
0 36745 5 1 1 67505
0 36746 7 1 2 41156 67506
0 36747 5 1 1 36746
0 36748 7 1 2 40303 64290
0 36749 5 1 1 36748
0 36750 7 1 2 64117 36749
0 36751 5 1 1 36750
0 36752 7 1 2 59483 36751
0 36753 5 1 1 36752
0 36754 7 1 2 36747 36753
0 36755 7 1 2 36737 36754
0 36756 5 1 1 36755
0 36757 7 1 2 45529 36756
0 36758 5 1 1 36757
0 36759 7 1 2 57826 63052
0 36760 5 1 1 36759
0 36761 7 1 2 36745 36760
0 36762 5 1 1 36761
0 36763 7 1 2 45353 36762
0 36764 5 1 1 36763
0 36765 7 1 2 2059 57830
0 36766 5 1 1 36765
0 36767 7 1 2 52401 60302
0 36768 7 1 2 64291 36767
0 36769 7 1 2 36766 36768
0 36770 5 1 1 36769
0 36771 7 1 2 36764 36770
0 36772 5 1 1 36771
0 36773 7 1 2 47134 36772
0 36774 5 1 1 36773
0 36775 7 1 2 52792 63295
0 36776 5 1 1 36775
0 36777 7 1 2 47824 63301
0 36778 5 1 1 36777
0 36779 7 1 2 36776 36778
0 36780 5 1 1 36779
0 36781 7 1 2 57217 58252
0 36782 7 1 2 36780 36781
0 36783 5 1 1 36782
0 36784 7 1 2 36774 36783
0 36785 7 1 2 36758 36784
0 36786 5 1 1 36785
0 36787 7 1 2 40524 36786
0 36788 5 1 1 36787
0 36789 7 1 2 47135 63792
0 36790 5 1 1 36789
0 36791 7 1 2 58287 63003
0 36792 5 1 1 36791
0 36793 7 1 2 36790 36792
0 36794 5 1 1 36793
0 36795 7 1 2 55133 36794
0 36796 5 1 1 36795
0 36797 7 1 2 67074 62897
0 36798 5 1 1 36797
0 36799 7 1 2 47136 63669
0 36800 7 1 2 59436 36799
0 36801 5 1 1 36800
0 36802 7 1 2 36798 36801
0 36803 5 1 1 36802
0 36804 7 1 2 60303 36803
0 36805 5 1 1 36804
0 36806 7 1 2 36796 36805
0 36807 5 1 1 36806
0 36808 7 1 2 40525 36807
0 36809 5 1 1 36808
0 36810 7 1 2 36809 67470
0 36811 5 1 1 36810
0 36812 7 1 2 52113 36811
0 36813 5 1 1 36812
0 36814 7 1 2 52333 59148
0 36815 5 1 1 36814
0 36816 7 1 2 32818 36815
0 36817 5 1 1 36816
0 36818 7 1 2 43274 36817
0 36819 5 1 1 36818
0 36820 7 1 2 56846 62235
0 36821 5 1 1 36820
0 36822 7 1 2 36819 36821
0 36823 5 1 1 36822
0 36824 7 1 2 59400 36823
0 36825 5 1 1 36824
0 36826 7 1 2 56847 57989
0 36827 5 1 1 36826
0 36828 7 1 2 52334 59059
0 36829 7 1 2 65097 36828
0 36830 5 1 1 36829
0 36831 7 1 2 36827 36830
0 36832 5 1 1 36831
0 36833 7 1 2 44303 36832
0 36834 5 1 1 36833
0 36835 7 1 2 41276 55022
0 36836 7 1 2 56848 36835
0 36837 5 1 1 36836
0 36838 7 1 2 36834 36837
0 36839 5 1 1 36838
0 36840 7 1 2 62983 36839
0 36841 5 1 1 36840
0 36842 7 1 2 36825 36841
0 36843 5 1 1 36842
0 36844 7 1 2 40526 36843
0 36845 5 1 1 36844
0 36846 7 1 2 46896 67136
0 36847 7 1 2 63858 36846
0 36848 7 1 2 63979 36847
0 36849 5 1 1 36848
0 36850 7 1 2 36845 36849
0 36851 5 1 1 36850
0 36852 7 1 2 47500 36851
0 36853 5 1 1 36852
0 36854 7 1 2 36813 36853
0 36855 7 1 2 36788 36854
0 36856 7 1 2 36721 36855
0 36857 5 1 1 36856
0 36858 7 1 2 45207 42891
0 36859 7 1 2 46531 36858
0 36860 7 1 2 65537 36859
0 36861 7 1 2 36857 36860
0 36862 5 1 1 36861
0 36863 7 1 2 36703 36862
0 36864 5 1 1 36863
0 36865 7 1 2 54371 36864
0 36866 5 1 1 36865
0 36867 7 2 2 51223 63296
0 36868 7 1 2 43973 67507
0 36869 5 1 1 36868
0 36870 7 1 2 58014 63302
0 36871 5 1 1 36870
0 36872 7 1 2 36869 36871
0 36873 5 1 1 36872
0 36874 7 1 2 41277 36873
0 36875 5 1 1 36874
0 36876 7 2 2 54448 67137
0 36877 7 1 2 61937 56588
0 36878 7 1 2 67509 36877
0 36879 5 1 1 36878
0 36880 7 1 2 36875 36879
0 36881 5 1 1 36880
0 36882 7 1 2 40304 36881
0 36883 5 1 1 36882
0 36884 7 2 2 45136 51224
0 36885 7 1 2 56595 67510
0 36886 7 1 2 67511 36885
0 36887 5 1 1 36886
0 36888 7 1 2 36883 36887
0 36889 5 1 1 36888
0 36890 7 1 2 40527 36889
0 36891 5 1 1 36890
0 36892 7 1 2 46312 67226
0 36893 7 1 2 67353 67512
0 36894 7 1 2 36892 36893
0 36895 5 1 1 36894
0 36896 7 1 2 36891 36895
0 36897 5 1 1 36896
0 36898 7 1 2 47501 36897
0 36899 5 1 1 36898
0 36900 7 1 2 60673 47254
0 36901 5 2 1 36900
0 36902 7 1 2 43974 36053
0 36903 5 1 1 36902
0 36904 7 1 2 67513 36903
0 36905 5 1 1 36904
0 36906 7 1 2 45354 36905
0 36907 5 1 1 36906
0 36908 7 1 2 60980 48801
0 36909 5 1 1 36908
0 36910 7 1 2 65965 36909
0 36911 5 2 1 36910
0 36912 7 1 2 45530 67515
0 36913 5 1 1 36912
0 36914 7 1 2 36907 36913
0 36915 5 1 1 36914
0 36916 7 1 2 67508 36915
0 36917 5 1 1 36916
0 36918 7 1 2 36899 36917
0 36919 5 1 1 36918
0 36920 7 1 2 42892 36919
0 36921 5 1 1 36920
0 36922 7 1 2 43605 65084
0 36923 5 1 1 36922
0 36924 7 2 2 47569 36923
0 36925 7 1 2 49720 67517
0 36926 5 1 1 36925
0 36927 7 1 2 67504 36926
0 36928 5 1 1 36927
0 36929 7 1 2 43793 36928
0 36930 5 1 1 36929
0 36931 7 1 2 67389 36930
0 36932 5 1 1 36931
0 36933 7 1 2 63316 63358
0 36934 7 1 2 36932 36933
0 36935 5 1 1 36934
0 36936 7 1 2 36921 36935
0 36937 5 1 1 36936
0 36938 7 1 2 57218 36937
0 36939 5 1 1 36938
0 36940 7 1 2 47155 67501
0 36941 5 1 1 36940
0 36942 7 1 2 47059 62457
0 36943 5 1 1 36942
0 36944 7 2 2 47073 36943
0 36945 5 1 1 67519
0 36946 7 1 2 36941 67520
0 36947 5 1 1 36946
0 36948 7 1 2 44448 50816
0 36949 5 1 1 36948
0 36950 7 1 2 56873 36949
0 36951 5 1 1 36950
0 36952 7 1 2 36947 36951
0 36953 5 1 1 36952
0 36954 7 1 2 45531 49715
0 36955 5 1 1 36954
0 36956 7 1 2 49753 51402
0 36957 7 1 2 36955 36956
0 36958 5 1 1 36957
0 36959 7 1 2 41540 49721
0 36960 7 1 2 65974 47960
0 36961 7 1 2 36959 36960
0 36962 5 1 1 36961
0 36963 7 1 2 36958 36962
0 36964 5 1 1 36963
0 36965 7 1 2 47671 36964
0 36966 5 1 1 36965
0 36967 7 1 2 49828 50817
0 36968 5 1 1 36967
0 36969 7 1 2 46723 53078
0 36970 5 1 1 36969
0 36971 7 1 2 50818 62585
0 36972 5 1 1 36971
0 36973 7 1 2 36970 36972
0 36974 5 1 1 36973
0 36975 7 1 2 49897 36974
0 36976 5 1 1 36975
0 36977 7 1 2 36968 36976
0 36978 7 1 2 36966 36977
0 36979 7 1 2 36953 36978
0 36980 5 1 1 36979
0 36981 7 2 2 43275 36980
0 36982 7 1 2 67451 67521
0 36983 5 1 1 36982
0 36984 7 1 2 46002 36983
0 36985 7 1 2 36939 36984
0 36986 5 1 1 36985
0 36987 7 1 2 50210 51354
0 36988 5 1 1 36987
0 36989 7 1 2 58093 36988
0 36990 5 1 1 36989
0 36991 7 1 2 57816 62377
0 36992 7 1 2 36990 36991
0 36993 5 1 1 36992
0 36994 7 1 2 23495 67406
0 36995 5 2 1 36994
0 36996 7 1 2 53723 67523
0 36997 5 2 1 36996
0 36998 7 2 2 43794 66746
0 36999 5 2 1 67527
0 37000 7 1 2 67525 67529
0 37001 5 1 1 37000
0 37002 7 2 2 51490 63150
0 37003 7 1 2 60332 63370
0 37004 7 1 2 67531 37003
0 37005 7 1 2 37001 37004
0 37006 5 1 1 37005
0 37007 7 1 2 36993 37006
0 37008 5 1 1 37007
0 37009 7 1 2 49966 37008
0 37010 5 1 1 37009
0 37011 7 1 2 50211 50853
0 37012 5 1 1 37011
0 37013 7 1 2 47825 50374
0 37014 5 1 1 37013
0 37015 7 1 2 37012 37014
0 37016 5 1 1 37015
0 37017 7 2 2 43276 58577
0 37018 7 1 2 58611 60024
0 37019 7 1 2 53269 62334
0 37020 7 1 2 37018 37019
0 37021 7 1 2 67533 37020
0 37022 7 1 2 37016 37021
0 37023 5 1 1 37022
0 37024 7 1 2 42725 37023
0 37025 7 1 2 37010 37024
0 37026 5 1 1 37025
0 37027 7 1 2 67373 37026
0 37028 7 1 2 36986 37027
0 37029 5 1 1 37028
0 37030 7 2 2 50705 67329
0 37031 7 2 2 55424 67535
0 37032 7 1 2 57714 64418
0 37033 7 1 2 67537 37032
0 37034 5 1 1 37033
0 37035 7 1 2 37029 37034
0 37036 7 1 2 36866 37035
0 37037 7 1 2 36612 37036
0 37038 7 1 2 36314 37037
0 37039 7 1 2 35993 37038
0 37040 5 1 1 37039
0 37041 7 1 2 49067 37040
0 37042 5 1 1 37041
0 37043 7 1 2 43460 66964
0 37044 5 1 1 37043
0 37045 7 3 2 49954 37044
0 37046 7 1 2 66747 67539
0 37047 5 1 1 37046
0 37048 7 1 2 47744 50375
0 37049 5 1 1 37048
0 37050 7 1 2 37047 37049
0 37051 5 1 1 37050
0 37052 7 2 2 60304 37051
0 37053 7 1 2 43795 58308
0 37054 7 1 2 67542 37053
0 37055 5 1 1 37054
0 37056 7 1 2 43796 63495
0 37057 5 1 1 37056
0 37058 7 1 2 51248 37057
0 37059 5 1 1 37058
0 37060 7 1 2 59484 60681
0 37061 7 1 2 37059 37060
0 37062 5 1 1 37061
0 37063 7 1 2 37055 37062
0 37064 5 1 1 37063
0 37065 7 1 2 54186 37064
0 37066 5 1 1 37065
0 37067 7 1 2 61024 60411
0 37068 7 1 2 61398 37067
0 37069 5 1 1 37068
0 37070 7 1 2 37066 37069
0 37071 5 1 1 37070
0 37072 7 1 2 51277 37071
0 37073 5 1 1 37072
0 37074 7 2 2 59668 66639
0 37075 5 1 1 67544
0 37076 7 1 2 48144 67545
0 37077 5 1 1 37076
0 37078 7 1 2 43461 48297
0 37079 7 1 2 61603 37078
0 37080 5 1 1 37079
0 37081 7 1 2 37077 37080
0 37082 5 1 1 37081
0 37083 7 1 2 45355 37082
0 37084 5 1 1 37083
0 37085 7 2 2 57188 56063
0 37086 5 1 1 67546
0 37087 7 1 2 51148 67547
0 37088 5 1 1 37087
0 37089 7 1 2 50155 51302
0 37090 7 1 2 59112 37089
0 37091 5 1 1 37090
0 37092 7 1 2 37088 37091
0 37093 5 1 1 37092
0 37094 7 1 2 44562 37093
0 37095 5 1 1 37094
0 37096 7 1 2 44449 63166
0 37097 7 1 2 60592 37096
0 37098 7 1 2 64243 37097
0 37099 5 1 1 37098
0 37100 7 1 2 37095 37099
0 37101 7 1 2 37084 37100
0 37102 5 1 1 37101
0 37103 7 1 2 43797 37102
0 37104 5 1 1 37103
0 37105 7 2 2 40889 58938
0 37106 7 2 2 53664 51303
0 37107 7 1 2 67548 67550
0 37108 5 1 1 37107
0 37109 7 1 2 37108 37086
0 37110 5 2 1 37109
0 37111 7 1 2 43606 65118
0 37112 5 2 1 37111
0 37113 7 1 2 50825 67524
0 37114 5 1 1 37113
0 37115 7 1 2 67554 37114
0 37116 5 2 1 37115
0 37117 7 1 2 67552 67556
0 37118 5 1 1 37117
0 37119 7 1 2 55799 64882
0 37120 5 2 1 37119
0 37121 7 1 2 54011 60486
0 37122 7 2 2 67558 37121
0 37123 5 1 1 67560
0 37124 7 1 2 48298 67561
0 37125 5 1 1 37124
0 37126 7 1 2 37118 37125
0 37127 7 1 2 37104 37126
0 37128 5 1 1 37127
0 37129 7 1 2 60305 37128
0 37130 5 1 1 37129
0 37131 7 1 2 44563 67172
0 37132 5 1 1 37131
0 37133 7 1 2 64965 62978
0 37134 7 2 2 60346 37133
0 37135 7 1 2 65119 67562
0 37136 5 1 1 37135
0 37137 7 1 2 37132 37136
0 37138 5 1 1 37137
0 37139 7 1 2 43607 37138
0 37140 5 1 1 37139
0 37141 7 1 2 65400 67563
0 37142 5 1 1 37141
0 37143 7 1 2 67174 37142
0 37144 5 1 1 37143
0 37145 7 1 2 43798 37144
0 37146 5 1 1 37145
0 37147 7 1 2 37140 37146
0 37148 5 1 1 37147
0 37149 7 1 2 54187 37148
0 37150 5 1 1 37149
0 37151 7 2 2 54988 56433
0 37152 7 3 2 43277 47672
0 37153 7 1 2 46641 49377
0 37154 7 1 2 67566 37153
0 37155 7 1 2 67564 37154
0 37156 5 1 1 37155
0 37157 7 1 2 37150 37156
0 37158 5 1 1 37157
0 37159 7 1 2 49722 37158
0 37160 5 1 1 37159
0 37161 7 1 2 40890 58928
0 37162 7 1 2 67565 37161
0 37163 5 1 1 37162
0 37164 7 1 2 54105 48299
0 37165 7 1 2 66181 37164
0 37166 5 1 1 37165
0 37167 7 1 2 37163 37166
0 37168 5 1 1 37167
0 37169 7 1 2 47673 37168
0 37170 5 1 1 37169
0 37171 7 1 2 62501 56426
0 37172 7 1 2 58706 37171
0 37173 5 1 1 37172
0 37174 7 1 2 60593 57772
0 37175 7 1 2 51313 37174
0 37176 5 1 1 37175
0 37177 7 1 2 37173 37176
0 37178 7 1 2 37170 37177
0 37179 5 1 1 37178
0 37180 7 1 2 59485 37179
0 37181 5 1 1 37180
0 37182 7 1 2 37160 37181
0 37183 7 1 2 37130 37182
0 37184 5 1 1 37183
0 37185 7 1 2 41682 37184
0 37186 5 1 1 37185
0 37187 7 1 2 37073 37186
0 37188 5 1 1 37187
0 37189 7 1 2 42195 37188
0 37190 5 1 1 37189
0 37191 7 1 2 63769 59752
0 37192 5 1 1 37191
0 37193 7 1 2 47861 66435
0 37194 7 1 2 63040 37193
0 37195 5 1 1 37194
0 37196 7 1 2 37192 37195
0 37197 5 1 1 37196
0 37198 7 1 2 54012 37197
0 37199 5 1 1 37198
0 37200 7 1 2 50387 52941
0 37201 7 1 2 61583 37200
0 37202 5 1 1 37201
0 37203 7 1 2 37199 37202
0 37204 5 1 1 37203
0 37205 7 1 2 44144 37204
0 37206 5 1 1 37205
0 37207 7 2 2 59211 60028
0 37208 7 1 2 50388 67534
0 37209 7 1 2 67569 37208
0 37210 5 1 1 37209
0 37211 7 1 2 37206 37210
0 37212 5 1 1 37211
0 37213 7 1 2 47674 37212
0 37214 5 1 1 37213
0 37215 7 1 2 54188 58714
0 37216 7 1 2 59623 37215
0 37217 5 1 1 37216
0 37218 7 1 2 62679 53143
0 37219 7 1 2 55185 37218
0 37220 5 1 1 37219
0 37221 7 1 2 37217 37220
0 37222 5 1 1 37221
0 37223 7 1 2 59486 37222
0 37224 5 1 1 37223
0 37225 7 1 2 37214 37224
0 37226 5 1 1 37225
0 37227 7 1 2 43799 37226
0 37228 5 1 1 37227
0 37229 7 1 2 46694 62689
0 37230 5 1 1 37229
0 37231 7 1 2 47436 64773
0 37232 5 1 1 37231
0 37233 7 1 2 44145 37232
0 37234 7 1 2 37230 37233
0 37235 5 1 1 37234
0 37236 7 1 2 40891 66752
0 37237 5 1 1 37236
0 37238 7 1 2 47745 61260
0 37239 7 1 2 37237 37238
0 37240 7 1 2 37235 37239
0 37241 5 1 1 37240
0 37242 7 1 2 37228 37241
0 37243 5 1 1 37242
0 37244 7 1 2 46313 37243
0 37245 5 1 1 37244
0 37246 7 1 2 37190 37245
0 37247 5 1 1 37246
0 37248 7 1 2 67374 37247
0 37249 5 1 1 37248
0 37250 7 1 2 47233 67337
0 37251 5 1 1 37250
0 37252 7 1 2 43800 52703
0 37253 5 1 1 37252
0 37254 7 1 2 37251 37253
0 37255 5 2 1 37254
0 37256 7 1 2 58556 64545
0 37257 7 1 2 67359 37256
0 37258 7 1 2 62776 37257
0 37259 7 1 2 67571 37258
0 37260 5 1 1 37259
0 37261 7 1 2 37249 37260
0 37262 5 1 1 37261
0 37263 7 1 2 43975 37262
0 37264 5 1 1 37263
0 37265 7 2 2 30320 67526
0 37266 7 1 2 67555 67573
0 37267 5 1 1 37266
0 37268 7 1 2 42196 37267
0 37269 5 1 1 37268
0 37270 7 1 2 52245 51149
0 37271 5 1 1 37270
0 37272 7 1 2 50196 54705
0 37273 5 1 1 37272
0 37274 7 1 2 37271 37273
0 37275 7 1 2 37269 37274
0 37276 5 1 1 37275
0 37277 7 1 2 54449 37276
0 37278 5 1 1 37277
0 37279 7 1 2 50533 64455
0 37280 5 1 1 37279
0 37281 7 1 2 49688 63027
0 37282 5 1 1 37281
0 37283 7 1 2 37280 37282
0 37284 7 1 2 37278 37283
0 37285 5 1 1 37284
0 37286 7 1 2 44374 43164
0 37287 7 1 2 46532 37286
0 37288 7 1 2 60106 37287
0 37289 7 1 2 37285 37288
0 37290 5 1 1 37289
0 37291 7 1 2 54106 54450
0 37292 7 1 2 67393 37291
0 37293 7 1 2 67338 37292
0 37294 5 1 1 37293
0 37295 7 1 2 37290 37294
0 37296 5 1 1 37295
0 37297 7 1 2 60306 37296
0 37298 5 1 1 37297
0 37299 7 1 2 62211 64456
0 37300 5 1 1 37299
0 37301 7 1 2 57071 54451
0 37302 7 1 2 51792 37301
0 37303 5 1 1 37302
0 37304 7 1 2 37300 37303
0 37305 5 1 1 37304
0 37306 7 1 2 65314 67280
0 37307 7 1 2 37305 37306
0 37308 5 1 1 37307
0 37309 7 1 2 37298 37308
0 37310 5 1 1 37309
0 37311 7 1 2 48280 37310
0 37312 5 1 1 37311
0 37313 7 1 2 67570 57284
0 37314 5 1 1 37313
0 37315 7 1 2 52831 19315
0 37316 5 1 1 37315
0 37317 7 1 2 37316 60215
0 37318 5 1 1 37317
0 37319 7 1 2 59784 54587
0 37320 7 1 2 64724 37319
0 37321 5 1 1 37320
0 37322 7 1 2 37318 37321
0 37323 5 1 1 37322
0 37324 7 1 2 60307 37323
0 37325 5 1 1 37324
0 37326 7 1 2 37314 37325
0 37327 5 1 1 37326
0 37328 7 2 2 46533 59730
0 37329 7 1 2 65538 67575
0 37330 7 1 2 54662 37329
0 37331 7 1 2 37327 37330
0 37332 5 1 1 37331
0 37333 7 1 2 37312 37332
0 37334 7 1 2 37264 37333
0 37335 5 1 1 37334
0 37336 7 1 2 54372 37335
0 37337 5 1 1 37336
0 37338 7 1 2 45532 61555
0 37339 5 1 1 37338
0 37340 7 1 2 60212 62934
0 37341 5 1 1 37340
0 37342 7 1 2 37339 37341
0 37343 5 1 1 37342
0 37344 7 1 2 65579 64213
0 37345 5 1 1 37344
0 37346 7 1 2 3475 37345
0 37347 5 1 1 37346
0 37348 7 1 2 37343 37347
0 37349 5 1 1 37348
0 37350 7 1 2 56631 60025
0 37351 7 1 2 52711 37350
0 37352 7 1 2 64646 37351
0 37353 7 1 2 63424 37352
0 37354 5 1 1 37353
0 37355 7 1 2 51339 57393
0 37356 7 1 2 63681 37355
0 37357 7 1 2 65580 37356
0 37358 5 1 1 37357
0 37359 7 1 2 37354 37358
0 37360 7 1 2 37349 37359
0 37361 5 1 1 37360
0 37362 7 1 2 40528 37361
0 37363 5 1 1 37362
0 37364 7 1 2 41683 65590
0 37365 5 1 1 37364
0 37366 7 1 2 37365 19511
0 37367 5 1 1 37366
0 37368 7 1 2 40892 37367
0 37369 5 1 1 37368
0 37370 7 1 2 56964 57313
0 37371 5 1 1 37370
0 37372 7 1 2 37369 37371
0 37373 5 1 1 37372
0 37374 7 1 2 46642 63079
0 37375 7 1 2 65886 37374
0 37376 7 1 2 37373 37375
0 37377 5 1 1 37376
0 37378 7 1 2 37363 37377
0 37379 5 1 1 37378
0 37380 7 1 2 67375 37379
0 37381 5 1 1 37380
0 37382 7 1 2 60650 67138
0 37383 7 1 2 62748 66798
0 37384 7 1 2 67360 64446
0 37385 7 1 2 37383 37384
0 37386 7 1 2 37382 37385
0 37387 5 1 1 37386
0 37388 7 1 2 37381 37387
0 37389 5 1 1 37388
0 37390 7 1 2 47502 37389
0 37391 5 1 1 37390
0 37392 7 1 2 45533 61584
0 37393 5 1 1 37392
0 37394 7 1 2 45356 62006
0 37395 5 1 1 37394
0 37396 7 1 2 47300 65890
0 37397 7 1 2 37395 37396
0 37398 5 1 1 37397
0 37399 7 1 2 65888 37398
0 37400 5 1 1 37399
0 37401 7 1 2 60308 37400
0 37402 5 1 1 37401
0 37403 7 1 2 37393 37402
0 37404 5 1 1 37403
0 37405 7 1 2 55309 37404
0 37406 5 1 1 37405
0 37407 7 1 2 60479 32838
0 37408 5 1 1 37407
0 37409 7 1 2 54013 37408
0 37410 5 1 1 37409
0 37411 7 1 2 61593 37410
0 37412 5 1 1 37411
0 37413 7 1 2 45534 37412
0 37414 5 1 1 37413
0 37415 7 1 2 59221 57332
0 37416 7 1 2 62130 37415
0 37417 5 1 1 37416
0 37418 7 1 2 37414 37417
0 37419 5 1 1 37418
0 37420 7 1 2 57338 37419
0 37421 5 1 1 37420
0 37422 7 1 2 37406 37421
0 37423 5 1 1 37422
0 37424 7 1 2 40529 37423
0 37425 5 1 1 37424
0 37426 7 1 2 51340 62882
0 37427 7 1 2 58253 37426
0 37428 7 1 2 55186 64647
0 37429 7 1 2 37427 37428
0 37430 5 1 1 37429
0 37431 7 1 2 37425 37430
0 37432 5 1 1 37431
0 37433 7 1 2 65581 37432
0 37434 5 1 1 37433
0 37435 7 2 2 54628 59624
0 37436 7 2 2 53931 67577
0 37437 5 1 1 67579
0 37438 7 3 2 52942 56356
0 37439 5 1 1 67581
0 37440 7 1 2 48292 37439
0 37441 5 2 1 37440
0 37442 7 1 2 54189 67584
0 37443 5 1 1 37442
0 37444 7 1 2 37437 37443
0 37445 5 1 1 37444
0 37446 7 2 2 55347 37445
0 37447 5 1 1 67586
0 37448 7 1 2 40530 67587
0 37449 5 1 1 37448
0 37450 7 1 2 65916 56434
0 37451 7 1 2 66994 37450
0 37452 5 1 1 37451
0 37453 7 1 2 64779 37452
0 37454 5 1 1 37453
0 37455 7 1 2 43044 37454
0 37456 5 1 1 37455
0 37457 7 1 2 67578 64717
0 37458 5 1 1 37457
0 37459 7 1 2 37456 37458
0 37460 5 1 1 37459
0 37461 7 1 2 58254 37460
0 37462 5 1 1 37461
0 37463 7 1 2 37449 37462
0 37464 5 1 1 37463
0 37465 7 1 2 59487 37464
0 37466 5 1 1 37465
0 37467 7 1 2 62002 48305
0 37468 5 1 1 37467
0 37469 7 1 2 66260 66825
0 37470 7 1 2 62171 37469
0 37471 5 1 1 37470
0 37472 7 1 2 37468 37471
0 37473 5 1 1 37472
0 37474 7 1 2 52628 55355
0 37475 7 1 2 60309 37474
0 37476 7 1 2 37473 37475
0 37477 5 1 1 37476
0 37478 7 1 2 37466 37477
0 37479 5 1 1 37478
0 37480 7 1 2 45535 37479
0 37481 5 1 1 37480
0 37482 7 1 2 64353 56446
0 37483 7 1 2 60059 37482
0 37484 7 1 2 46819 56614
0 37485 7 1 2 61716 37484
0 37486 7 1 2 37483 37485
0 37487 7 1 2 48306 37486
0 37488 5 1 1 37487
0 37489 7 1 2 37481 37488
0 37490 7 1 2 37434 37489
0 37491 5 1 1 37490
0 37492 7 1 2 67376 37491
0 37493 5 1 1 37492
0 37494 7 1 2 37391 37493
0 37495 5 1 1 37494
0 37496 7 1 2 47826 37495
0 37497 5 1 1 37496
0 37498 7 2 2 49898 54014
0 37499 5 1 1 67588
0 37500 7 1 2 67151 67589
0 37501 5 1 1 37500
0 37502 7 2 2 49899 58258
0 37503 5 1 1 67590
0 37504 7 1 2 49820 61231
0 37505 7 1 2 37503 37504
0 37506 5 1 1 37505
0 37507 7 1 2 54190 54515
0 37508 7 1 2 37506 37507
0 37509 5 1 1 37508
0 37510 7 1 2 37501 37509
0 37511 5 1 1 37510
0 37512 7 1 2 62012 37511
0 37513 5 1 1 37512
0 37514 7 1 2 67530 67574
0 37515 5 2 1 37514
0 37516 7 1 2 64512 67592
0 37517 5 1 1 37516
0 37518 7 1 2 60981 52289
0 37519 5 1 1 37518
0 37520 7 1 2 47524 66131
0 37521 5 1 1 37520
0 37522 7 1 2 37519 37521
0 37523 5 1 1 37522
0 37524 7 1 2 41278 37523
0 37525 5 1 1 37524
0 37526 7 1 2 55144 66737
0 37527 5 1 1 37526
0 37528 7 1 2 31052 37527
0 37529 5 2 1 37528
0 37530 7 1 2 43801 67594
0 37531 5 1 1 37530
0 37532 7 1 2 49766 64879
0 37533 5 2 1 37532
0 37534 7 1 2 37531 67596
0 37535 5 1 1 37534
0 37536 7 1 2 62442 37535
0 37537 5 1 1 37536
0 37538 7 1 2 37525 37537
0 37539 5 1 1 37538
0 37540 7 1 2 54191 37539
0 37541 5 1 1 37540
0 37542 7 1 2 37517 37541
0 37543 5 1 1 37542
0 37544 7 1 2 54293 37543
0 37545 5 1 1 37544
0 37546 7 1 2 60716 56965
0 37547 7 1 2 67593 37546
0 37548 5 1 1 37547
0 37549 7 1 2 37545 37548
0 37550 5 1 1 37549
0 37551 7 1 2 60310 37550
0 37552 5 1 1 37551
0 37553 7 1 2 37513 37552
0 37554 5 1 1 37553
0 37555 7 1 2 42197 37554
0 37556 5 1 1 37555
0 37557 7 1 2 49156 58639
0 37558 7 1 2 58711 37557
0 37559 5 1 1 37558
0 37560 7 1 2 61585 37559
0 37561 5 1 1 37560
0 37562 7 1 2 44450 49154
0 37563 7 1 2 62219 37562
0 37564 5 1 1 37563
0 37565 7 1 2 37561 37564
0 37566 5 1 1 37565
0 37567 7 1 2 43802 37566
0 37568 5 1 1 37567
0 37569 7 1 2 61586 58816
0 37570 5 1 1 37569
0 37571 7 1 2 37568 37570
0 37572 5 1 1 37571
0 37573 7 1 2 40695 37572
0 37574 5 1 1 37573
0 37575 7 1 2 65964 62220
0 37576 5 1 1 37575
0 37577 7 1 2 37574 37576
0 37578 5 1 1 37577
0 37579 7 1 2 57366 37578
0 37580 5 1 1 37579
0 37581 7 1 2 47437 62158
0 37582 5 1 1 37581
0 37583 7 1 2 65966 37582
0 37584 5 1 1 37583
0 37585 7 1 2 62221 37584
0 37586 5 1 1 37585
0 37587 7 1 2 66132 62265
0 37588 5 1 1 37587
0 37589 7 1 2 37586 37588
0 37590 5 1 1 37589
0 37591 7 1 2 54294 37590
0 37592 5 1 1 37591
0 37593 7 1 2 13897 65967
0 37594 5 2 1 37593
0 37595 7 1 2 60472 57367
0 37596 5 1 1 37595
0 37597 7 1 2 52797 54295
0 37598 7 1 2 62059 37597
0 37599 5 1 1 37598
0 37600 7 1 2 37596 37599
0 37601 5 1 1 37600
0 37602 7 1 2 54192 37601
0 37603 5 1 1 37602
0 37604 7 1 2 47503 54015
0 37605 7 1 2 61295 37604
0 37606 7 1 2 67152 37605
0 37607 5 1 1 37606
0 37608 7 1 2 37603 37607
0 37609 5 1 1 37608
0 37610 7 1 2 67598 37609
0 37611 5 1 1 37610
0 37612 7 1 2 37592 37611
0 37613 7 1 2 37580 37612
0 37614 7 1 2 37556 37613
0 37615 5 1 1 37614
0 37616 7 1 2 67377 37615
0 37617 5 1 1 37616
0 37618 7 1 2 65985 67330
0 37619 7 1 2 64419 37618
0 37620 7 1 2 67153 37619
0 37621 7 1 2 67339 37620
0 37622 5 1 1 37621
0 37623 7 1 2 37617 37622
0 37624 5 1 1 37623
0 37625 7 1 2 48281 37624
0 37626 5 1 1 37625
0 37627 7 1 2 37497 37626
0 37628 7 1 2 61594 13163
0 37629 5 1 1 37628
0 37630 7 1 2 64214 37629
0 37631 5 1 1 37630
0 37632 7 1 2 42893 57618
0 37633 7 1 2 62247 59994
0 37634 7 1 2 37632 37633
0 37635 5 1 1 37634
0 37636 7 1 2 37631 37635
0 37637 5 1 1 37636
0 37638 7 1 2 47301 37637
0 37639 5 1 1 37638
0 37640 7 1 2 54193 57676
0 37641 5 2 1 37640
0 37642 7 1 2 11084 67600
0 37643 5 1 1 37642
0 37644 7 1 2 40893 37643
0 37645 5 1 1 37644
0 37646 7 1 2 54194 64641
0 37647 5 1 1 37646
0 37648 7 1 2 37645 37647
0 37649 5 1 1 37648
0 37650 7 1 2 43045 37649
0 37651 5 1 1 37650
0 37652 7 1 2 57849 57339
0 37653 5 1 1 37652
0 37654 7 1 2 61097 48282
0 37655 5 1 1 37654
0 37656 7 1 2 66468 37655
0 37657 5 1 1 37656
0 37658 7 1 2 44146 37657
0 37659 5 1 1 37658
0 37660 7 1 2 61098 64208
0 37661 5 1 1 37660
0 37662 7 1 2 37659 37661
0 37663 5 1 1 37662
0 37664 7 1 2 40127 37663
0 37665 5 1 1 37664
0 37666 7 1 2 37653 37665
0 37667 7 1 2 37651 37666
0 37668 5 1 1 37667
0 37669 7 1 2 59488 37668
0 37670 5 1 1 37669
0 37671 7 1 2 37639 37670
0 37672 5 1 1 37671
0 37673 7 1 2 65582 37672
0 37674 5 1 1 37673
0 37675 7 1 2 60473 66648
0 37676 5 1 1 37675
0 37677 7 1 2 62323 37676
0 37678 5 1 1 37677
0 37679 7 1 2 40128 37678
0 37680 5 1 1 37679
0 37681 7 1 2 57839 59489
0 37682 5 1 1 37681
0 37683 7 1 2 37680 37682
0 37684 5 1 1 37683
0 37685 7 1 2 48307 37684
0 37686 5 1 1 37685
0 37687 7 1 2 66742 59625
0 37688 5 1 1 37687
0 37689 7 1 2 56977 58309
0 37690 7 1 2 65341 37689
0 37691 5 1 1 37690
0 37692 7 1 2 37688 37691
0 37693 5 1 1 37692
0 37694 7 1 2 46314 37693
0 37695 5 1 1 37694
0 37696 7 3 2 59611 63676
0 37697 5 1 1 67602
0 37698 7 1 2 46174 67603
0 37699 5 1 1 37698
0 37700 7 1 2 37695 37699
0 37701 5 1 1 37700
0 37702 7 1 2 59490 37701
0 37703 5 1 1 37702
0 37704 7 1 2 37686 37703
0 37705 5 1 1 37704
0 37706 7 1 2 49620 37705
0 37707 5 1 1 37706
0 37708 7 1 2 54016 58430
0 37709 5 1 1 37708
0 37710 7 1 2 46444 49121
0 37711 7 1 2 50854 37710
0 37712 7 1 2 58955 37711
0 37713 5 1 1 37712
0 37714 7 1 2 37709 37713
0 37715 5 1 1 37714
0 37716 7 1 2 63080 63757
0 37717 7 1 2 37715 37716
0 37718 5 1 1 37717
0 37719 7 1 2 37707 37718
0 37720 5 1 1 37719
0 37721 7 1 2 42726 37720
0 37722 5 1 1 37721
0 37723 7 1 2 55657 61980
0 37724 7 1 2 66236 37723
0 37725 7 1 2 66995 37724
0 37726 5 1 1 37725
0 37727 7 1 2 37722 37726
0 37728 7 1 2 37674 37727
0 37729 5 1 1 37728
0 37730 7 1 2 50212 37729
0 37731 5 1 1 37730
0 37732 7 1 2 66161 52943
0 37733 5 1 1 37732
0 37734 7 2 2 49754 48802
0 37735 7 1 2 49096 67605
0 37736 5 1 1 37735
0 37737 7 1 2 37733 37736
0 37738 5 1 1 37737
0 37739 7 1 2 61966 37738
0 37740 5 1 1 37739
0 37741 7 1 2 64619 67606
0 37742 5 1 1 37741
0 37743 7 1 2 4460 51648
0 37744 5 1 1 37743
0 37745 7 1 2 58212 53270
0 37746 7 1 2 37744 37745
0 37747 5 1 1 37746
0 37748 7 1 2 37742 37747
0 37749 7 1 2 37740 37748
0 37750 5 1 1 37749
0 37751 7 1 2 54373 37750
0 37752 5 1 1 37751
0 37753 7 1 2 64747 59375
0 37754 5 1 1 37753
0 37755 7 1 2 50739 64549
0 37756 5 1 1 37755
0 37757 7 1 2 48283 67154
0 37758 5 1 1 37757
0 37759 7 1 2 37756 37758
0 37760 7 1 2 37754 37759
0 37761 5 1 1 37760
0 37762 7 1 2 67516 37761
0 37763 5 1 1 37762
0 37764 7 1 2 49146 61214
0 37765 7 1 2 51257 37764
0 37766 5 1 1 37765
0 37767 7 1 2 37763 37766
0 37768 7 1 2 37752 37767
0 37769 5 1 1 37768
0 37770 7 1 2 54017 37769
0 37771 5 1 1 37770
0 37772 7 1 2 41684 65663
0 37773 5 1 1 37772
0 37774 7 1 2 55414 53361
0 37775 5 1 1 37774
0 37776 7 1 2 37773 37775
0 37777 5 1 1 37776
0 37778 7 1 2 40894 37777
0 37779 5 1 1 37778
0 37780 7 1 2 41685 64571
0 37781 5 1 1 37780
0 37782 7 1 2 37779 37781
0 37783 5 1 1 37782
0 37784 7 1 2 61516 37783
0 37785 5 1 1 37784
0 37786 7 1 2 41279 67595
0 37787 5 1 1 37786
0 37788 7 1 2 47525 65401
0 37789 5 1 1 37788
0 37790 7 1 2 37787 37789
0 37791 5 1 1 37790
0 37792 7 1 2 65583 55305
0 37793 5 1 1 37792
0 37794 7 1 2 57314 54460
0 37795 5 1 1 37794
0 37796 7 1 2 37793 37795
0 37797 5 1 1 37796
0 37798 7 1 2 40531 37797
0 37799 7 1 2 37791 37798
0 37800 5 1 1 37799
0 37801 7 1 2 43046 37800
0 37802 7 1 2 37785 37801
0 37803 5 1 1 37802
0 37804 7 1 2 44978 56479
0 37805 5 1 1 37804
0 37806 7 1 2 41686 61179
0 37807 5 1 1 37806
0 37808 7 1 2 37805 37807
0 37809 5 1 1 37808
0 37810 7 1 2 50124 37809
0 37811 5 1 1 37810
0 37812 7 1 2 65968 13557
0 37813 5 1 1 37812
0 37814 7 1 2 65557 37813
0 37815 5 1 1 37814
0 37816 7 1 2 56952 64758
0 37817 5 1 1 37816
0 37818 7 1 2 37815 37817
0 37819 5 1 1 37818
0 37820 7 1 2 44979 37819
0 37821 5 1 1 37820
0 37822 7 1 2 37811 37821
0 37823 5 1 1 37822
0 37824 7 1 2 44147 37823
0 37825 5 1 1 37824
0 37826 7 1 2 59324 67216
0 37827 7 1 2 61180 37826
0 37828 5 1 1 37827
0 37829 7 1 2 37825 37828
0 37830 5 1 1 37829
0 37831 7 1 2 67540 37830
0 37832 5 1 1 37831
0 37833 7 1 2 64103 60852
0 37834 7 1 2 66748 37833
0 37835 7 1 2 67271 37834
0 37836 5 1 1 37835
0 37837 7 1 2 46315 37836
0 37838 7 1 2 37832 37837
0 37839 5 1 1 37838
0 37840 7 1 2 54195 37839
0 37841 7 1 2 37803 37840
0 37842 5 1 1 37841
0 37843 7 1 2 37771 37842
0 37844 5 1 1 37843
0 37845 7 1 2 60311 37844
0 37846 5 1 1 37845
0 37847 7 1 2 37731 37846
0 37848 5 1 1 37847
0 37849 7 1 2 67378 37848
0 37850 5 1 1 37849
0 37851 7 2 2 63481 67361
0 37852 7 2 2 41054 44833
0 37853 7 1 2 50213 67609
0 37854 7 1 2 66977 66799
0 37855 7 1 2 37853 37854
0 37856 7 1 2 67607 37855
0 37857 5 1 1 37856
0 37858 7 1 2 37850 37857
0 37859 5 1 1 37858
0 37860 7 1 2 45536 37859
0 37861 5 1 1 37860
0 37862 7 1 2 56953 52844
0 37863 7 1 2 58807 37862
0 37864 5 1 1 37863
0 37865 7 1 2 47504 67599
0 37866 5 1 1 37865
0 37867 7 1 2 65969 67514
0 37868 5 1 1 37867
0 37869 7 1 2 45357 37868
0 37870 5 1 1 37869
0 37871 7 1 2 37866 37870
0 37872 5 1 1 37871
0 37873 7 1 2 42727 56357
0 37874 7 1 2 37872 37873
0 37875 5 1 1 37874
0 37876 7 1 2 37864 37875
0 37877 5 1 1 37876
0 37878 7 1 2 60312 37877
0 37879 5 1 1 37878
0 37880 7 1 2 61889 62885
0 37881 7 2 2 67293 37880
0 37882 7 1 2 43976 59123
0 37883 7 1 2 67611 37882
0 37884 5 1 1 37883
0 37885 7 1 2 37879 37884
0 37886 5 1 1 37885
0 37887 7 1 2 41687 37886
0 37888 5 1 1 37887
0 37889 7 1 2 43977 60029
0 37890 7 1 2 67612 37889
0 37891 5 1 1 37890
0 37892 7 1 2 42894 37891
0 37893 7 1 2 37888 37892
0 37894 5 1 1 37893
0 37895 7 2 2 43803 64608
0 37896 7 2 2 67613 62327
0 37897 5 1 1 67615
0 37898 7 1 2 44451 67616
0 37899 5 1 1 37898
0 37900 7 2 2 59035 65171
0 37901 7 1 2 44452 65079
0 37902 7 1 2 64609 37901
0 37903 7 1 2 67617 37902
0 37904 5 1 1 37903
0 37905 7 1 2 18470 37904
0 37906 5 1 1 37905
0 37907 7 1 2 47675 37906
0 37908 5 1 1 37907
0 37909 7 1 2 37899 37908
0 37910 5 1 1 37909
0 37911 7 1 2 42000 37910
0 37912 5 1 1 37911
0 37913 7 1 2 49755 67618
0 37914 7 1 2 62329 37913
0 37915 5 1 1 37914
0 37916 7 1 2 37912 37915
0 37917 5 1 1 37916
0 37918 7 1 2 43462 37917
0 37919 5 1 1 37918
0 37920 7 2 2 54828 61270
0 37921 7 1 2 67475 67619
0 37922 5 1 1 37921
0 37923 7 1 2 37919 37922
0 37924 5 1 1 37923
0 37925 7 1 2 64019 37924
0 37926 5 1 1 37925
0 37927 7 1 2 44453 63919
0 37928 5 2 1 37927
0 37929 7 1 2 37897 67621
0 37930 5 1 1 37929
0 37931 7 1 2 43608 37930
0 37932 5 1 1 37931
0 37933 7 1 2 40305 67620
0 37934 5 1 1 37933
0 37935 7 1 2 67622 37934
0 37936 5 1 1 37935
0 37937 7 1 2 44564 37936
0 37938 5 1 1 37937
0 37939 7 1 2 37932 37938
0 37940 5 1 1 37939
0 37941 7 1 2 64020 37940
0 37942 5 1 1 37941
0 37943 7 1 2 59913 48406
0 37944 7 1 2 66953 37943
0 37945 7 1 2 67567 37944
0 37946 5 1 1 37945
0 37947 7 1 2 37942 37946
0 37948 5 1 1 37947
0 37949 7 1 2 49723 37948
0 37950 5 1 1 37949
0 37951 7 1 2 41280 67499
0 37952 5 2 1 37951
0 37953 7 1 2 65975 63081
0 37954 7 1 2 54506 37953
0 37955 7 1 2 63059 37954
0 37956 7 1 2 67623 37955
0 37957 5 1 1 37956
0 37958 7 1 2 37950 37957
0 37959 7 1 2 37926 37958
0 37960 5 1 1 37959
0 37961 7 1 2 42198 37960
0 37962 5 1 1 37961
0 37963 7 1 2 54829 59995
0 37964 5 1 1 37963
0 37965 7 1 2 47360 53271
0 37966 7 1 2 57905 37965
0 37967 5 1 1 37966
0 37968 7 1 2 37964 37967
0 37969 5 1 1 37968
0 37970 7 1 2 49900 37969
0 37971 5 1 1 37970
0 37972 7 1 2 52610 64400
0 37973 7 1 2 51118 37972
0 37974 5 1 1 37973
0 37975 7 1 2 37971 37974
0 37976 5 1 1 37975
0 37977 7 1 2 42001 37976
0 37978 5 1 1 37977
0 37979 7 1 2 62159 63587
0 37980 5 1 1 37979
0 37981 7 1 2 37978 37980
0 37982 5 1 1 37981
0 37983 7 1 2 59491 37982
0 37984 5 1 1 37983
0 37985 7 1 2 46175 37984
0 37986 7 1 2 37962 37985
0 37987 5 1 1 37986
0 37988 7 1 2 37894 37987
0 37989 5 1 1 37988
0 37990 7 1 2 44834 37989
0 37991 5 1 1 37990
0 37992 7 1 2 55720 63193
0 37993 5 1 1 37992
0 37994 7 1 2 53844 64892
0 37995 7 1 2 51089 37994
0 37996 7 1 2 60313 37995
0 37997 5 1 1 37996
0 37998 7 1 2 37993 37997
0 37999 5 1 1 37998
0 38000 7 1 2 43609 37999
0 38001 5 1 1 38000
0 38002 7 1 2 52697 56919
0 38003 7 1 2 67189 38002
0 38004 5 1 1 38003
0 38005 7 1 2 46003 62757
0 38006 7 1 2 61884 38005
0 38007 5 1 1 38006
0 38008 7 1 2 38004 38007
0 38009 5 1 1 38008
0 38010 7 1 2 43804 38009
0 38011 5 1 1 38010
0 38012 7 1 2 62758 62009
0 38013 7 1 2 66327 38012
0 38014 5 1 1 38013
0 38015 7 1 2 38011 38014
0 38016 7 1 2 38001 38015
0 38017 5 1 1 38016
0 38018 7 1 2 64615 38017
0 38019 5 1 1 38018
0 38020 7 2 2 46643 57362
0 38021 7 1 2 48133 52190
0 38022 7 1 2 67568 38021
0 38023 7 1 2 67625 38022
0 38024 5 1 1 38023
0 38025 7 1 2 38019 38024
0 38026 5 1 1 38025
0 38027 7 1 2 47361 38026
0 38028 5 1 1 38027
0 38029 7 1 2 56596 62567
0 38030 5 1 1 38029
0 38031 7 1 2 65402 67614
0 38032 5 1 1 38031
0 38033 7 1 2 38030 38032
0 38034 5 1 1 38033
0 38035 7 1 2 42199 63738
0 38036 7 1 2 38034 38035
0 38037 5 1 1 38036
0 38038 7 1 2 61376 58154
0 38039 5 1 1 38038
0 38040 7 1 2 61890 50061
0 38041 7 1 2 67626 38040
0 38042 7 1 2 38039 38041
0 38043 5 1 1 38042
0 38044 7 1 2 38037 38043
0 38045 5 1 1 38044
0 38046 7 1 2 46176 38045
0 38047 5 1 1 38046
0 38048 7 1 2 55721 51278
0 38049 7 1 2 59492 38048
0 38050 7 1 2 67290 38049
0 38051 5 1 1 38050
0 38052 7 1 2 38047 38051
0 38053 7 1 2 38028 38052
0 38054 5 1 1 38053
0 38055 7 1 2 44148 38054
0 38056 5 1 1 38055
0 38057 7 1 2 48444 64255
0 38058 7 1 2 61261 38057
0 38059 7 1 2 61379 38058
0 38060 5 1 1 38059
0 38061 7 1 2 41541 38060
0 38062 7 1 2 38056 38061
0 38063 5 1 1 38062
0 38064 7 1 2 67379 38063
0 38065 7 1 2 37991 38064
0 38066 5 1 1 38065
0 38067 7 1 2 52646 58557
0 38068 7 1 2 67044 38067
0 38069 7 1 2 60664 67536
0 38070 7 1 2 38068 38069
0 38071 5 1 1 38070
0 38072 7 1 2 38066 38071
0 38073 5 1 1 38072
0 38074 7 1 2 54018 38073
0 38075 5 1 1 38074
0 38076 7 1 2 37861 38075
0 38077 7 1 2 37627 38076
0 38078 7 1 2 37337 38077
0 38079 7 1 2 43283 59513
0 38080 7 2 2 63060 38079
0 38081 5 1 1 67627
0 38082 7 2 2 52944 61367
0 38083 7 1 2 62787 67281
0 38084 7 1 2 67629 38083
0 38085 5 1 1 38084
0 38086 7 1 2 38081 38085
0 38087 5 1 1 38086
0 38088 7 1 2 47676 38087
0 38089 5 1 1 38088
0 38090 7 4 2 44304 67282
0 38091 7 9 2 45137 67631
0 38092 7 2 2 52945 67635
0 38093 7 1 2 47746 67644
0 38094 5 1 1 38093
0 38095 7 1 2 42002 67628
0 38096 5 1 1 38095
0 38097 7 1 2 38094 38096
0 38098 5 1 1 38097
0 38099 7 1 2 47362 38098
0 38100 5 1 1 38099
0 38101 7 1 2 38089 38100
0 38102 5 1 1 38101
0 38103 7 1 2 42200 38102
0 38104 5 1 1 38103
0 38105 7 5 2 46644 67331
0 38106 7 1 2 60558 67646
0 38107 5 1 1 38106
0 38108 7 1 2 67645 52118
0 38109 5 1 1 38108
0 38110 7 1 2 38107 38109
0 38111 5 1 1 38110
0 38112 7 1 2 43805 38111
0 38113 5 1 1 38112
0 38114 7 1 2 64995 67632
0 38115 7 1 2 67630 38114
0 38116 5 1 1 38115
0 38117 7 1 2 38113 38116
0 38118 7 1 2 38104 38117
0 38119 5 1 1 38118
0 38120 7 1 2 44149 38119
0 38121 5 1 1 38120
0 38122 7 2 2 67283 52300
0 38123 7 1 2 60347 66437
0 38124 7 1 2 67651 38123
0 38125 5 1 1 38124
0 38126 7 1 2 38121 38125
0 38127 5 1 1 38126
0 38128 7 1 2 54196 38127
0 38129 5 1 1 38128
0 38130 7 1 2 46695 61090
0 38131 5 1 1 38130
0 38132 7 1 2 52749 38131
0 38133 5 1 1 38132
0 38134 7 1 2 49901 38133
0 38135 5 1 1 38134
0 38136 7 1 2 50214 63407
0 38137 5 1 1 38136
0 38138 7 1 2 46696 38137
0 38139 5 1 1 38138
0 38140 7 1 2 38135 38139
0 38141 5 1 1 38140
0 38142 7 4 2 46534 60373
0 38143 7 1 2 67653 59227
0 38144 7 1 2 38141 38143
0 38145 5 1 1 38144
0 38146 7 1 2 38129 38145
0 38147 5 1 1 38146
0 38148 7 1 2 46316 38147
0 38149 5 1 1 38148
0 38150 7 2 2 54989 67284
0 38151 7 1 2 52698 67657
0 38152 7 1 2 63682 38151
0 38153 7 1 2 60428 38152
0 38154 5 1 1 38153
0 38155 7 1 2 38149 38154
0 38156 5 1 1 38155
0 38157 7 1 2 43978 38156
0 38158 5 1 1 38157
0 38159 7 4 2 58991 67654
0 38160 7 1 2 44565 67659
0 38161 5 1 1 38160
0 38162 7 1 2 61567 67332
0 38163 7 2 2 62343 38162
0 38164 5 1 1 67663
0 38165 7 1 2 38161 38164
0 38166 5 1 1 38165
0 38167 7 1 2 43610 38166
0 38168 5 1 1 38167
0 38169 7 1 2 43806 67660
0 38170 5 1 1 38169
0 38171 7 1 2 54197 67647
0 38172 7 1 2 53733 38171
0 38173 5 1 1 38172
0 38174 7 1 2 38170 38173
0 38175 7 1 2 38168 38174
0 38176 5 1 1 38175
0 38177 7 1 2 42201 38176
0 38178 5 1 1 38177
0 38179 7 1 2 43807 67664
0 38180 5 1 1 38179
0 38181 7 1 2 38178 38180
0 38182 5 2 1 38181
0 38183 7 1 2 54452 67665
0 38184 5 1 1 38183
0 38185 7 1 2 65679 56954
0 38186 7 2 2 41281 67285
0 38187 7 1 2 66783 67667
0 38188 7 1 2 38185 38187
0 38189 5 1 1 38188
0 38190 7 1 2 38184 38189
0 38191 5 1 1 38190
0 38192 7 1 2 48284 38191
0 38193 5 1 1 38192
0 38194 7 1 2 44980 64966
0 38195 7 1 2 67286 38194
0 38196 7 2 2 56637 38195
0 38197 7 1 2 56597 49122
0 38198 7 1 2 56955 38197
0 38199 7 1 2 67669 38198
0 38200 5 1 1 38199
0 38201 7 1 2 38193 38200
0 38202 7 1 2 38158 38201
0 38203 5 1 1 38202
0 38204 7 1 2 54374 38203
0 38205 5 1 1 38204
0 38206 7 2 2 65558 51279
0 38207 7 1 2 43463 67671
0 38208 5 1 1 38207
0 38209 7 1 2 57603 51225
0 38210 5 1 1 38209
0 38211 7 1 2 38208 38210
0 38212 5 1 1 38211
0 38213 7 1 2 44150 38212
0 38214 5 1 1 38213
0 38215 7 1 2 62613 62950
0 38216 5 1 1 38215
0 38217 7 1 2 38214 38216
0 38218 5 1 1 38217
0 38219 7 1 2 46853 38218
0 38220 5 1 1 38219
0 38221 7 2 2 43047 67155
0 38222 7 1 2 61113 67673
0 38223 5 1 1 38222
0 38224 7 1 2 65654 56474
0 38225 5 1 1 38224
0 38226 7 1 2 38223 38225
0 38227 5 1 1 38226
0 38228 7 1 2 46177 38227
0 38229 5 1 1 38228
0 38230 7 2 2 48244 48315
0 38231 5 1 1 67675
0 38232 7 1 2 55472 50403
0 38233 7 1 2 67676 38232
0 38234 5 1 1 38233
0 38235 7 1 2 38229 38234
0 38236 7 1 2 38220 38235
0 38237 5 1 1 38236
0 38238 7 1 2 47677 38237
0 38239 5 1 1 38238
0 38240 7 1 2 67674 63374
0 38241 5 1 1 38240
0 38242 7 1 2 38239 38241
0 38243 5 1 1 38242
0 38244 7 1 2 67661 38243
0 38245 5 1 1 38244
0 38246 7 2 2 49168 67648
0 38247 5 1 1 67677
0 38248 7 2 2 48445 67636
0 38249 7 1 2 66182 67679
0 38250 5 1 1 38249
0 38251 7 1 2 38247 38250
0 38252 5 1 1 38251
0 38253 7 1 2 47678 38252
0 38254 5 1 1 38253
0 38255 7 1 2 67591 67680
0 38256 5 1 1 38255
0 38257 7 1 2 53724 67678
0 38258 5 1 1 38257
0 38259 7 1 2 38256 38258
0 38260 7 1 2 38254 38259
0 38261 5 1 1 38260
0 38262 7 1 2 54284 38261
0 38263 5 1 1 38262
0 38264 7 1 2 63770 67333
0 38265 7 1 2 62452 38264
0 38266 5 1 1 38265
0 38267 7 1 2 38263 38266
0 38268 5 1 1 38267
0 38269 7 1 2 46317 38268
0 38270 5 1 1 38269
0 38271 7 1 2 46535 61891
0 38272 7 1 2 63975 38271
0 38273 7 1 2 67532 38272
0 38274 7 1 2 61399 38273
0 38275 5 1 1 38274
0 38276 7 1 2 38270 38275
0 38277 5 1 1 38276
0 38278 7 1 2 42895 38277
0 38279 5 1 1 38278
0 38280 7 3 2 43284 64603
0 38281 7 1 2 61193 62751
0 38282 7 1 2 67681 38281
0 38283 5 1 1 38282
0 38284 7 2 2 59036 51494
0 38285 7 1 2 67633 67684
0 38286 7 1 2 46936 38285
0 38287 5 1 1 38286
0 38288 7 1 2 38283 38287
0 38289 5 1 1 38288
0 38290 7 1 2 46697 38289
0 38291 5 1 1 38290
0 38292 7 1 2 38279 38291
0 38293 5 1 1 38292
0 38294 7 1 2 54198 38293
0 38295 5 1 1 38294
0 38296 7 1 2 38245 38295
0 38297 5 1 1 38296
0 38298 7 1 2 42202 38297
0 38299 5 1 1 38298
0 38300 7 1 2 65559 66367
0 38301 5 1 1 38300
0 38302 7 1 2 47363 62603
0 38303 7 1 2 66588 38302
0 38304 5 1 1 38303
0 38305 7 1 2 38301 38304
0 38306 5 1 1 38305
0 38307 7 1 2 44981 38306
0 38308 5 1 1 38307
0 38309 7 1 2 57760 64751
0 38310 5 1 1 38309
0 38311 7 1 2 38308 38310
0 38312 5 1 1 38311
0 38313 7 1 2 47679 38312
0 38314 5 1 1 38313
0 38315 7 1 2 47747 49123
0 38316 7 1 2 60766 38315
0 38317 7 1 2 66589 38316
0 38318 5 1 1 38317
0 38319 7 1 2 38314 38318
0 38320 5 1 1 38319
0 38321 7 1 2 43808 38320
0 38322 5 1 1 38321
0 38323 7 1 2 43464 67553
0 38324 5 1 1 38323
0 38325 7 1 2 48147 38231
0 38326 5 1 1 38325
0 38327 7 1 2 54019 38326
0 38328 5 1 1 38327
0 38329 7 1 2 38324 38328
0 38330 5 1 1 38329
0 38331 7 1 2 49902 38330
0 38332 5 1 1 38331
0 38333 7 1 2 62477 60786
0 38334 5 1 1 38333
0 38335 7 1 2 47680 48145
0 38336 7 1 2 38334 38335
0 38337 5 1 1 38336
0 38338 7 1 2 38332 38337
0 38339 5 1 1 38338
0 38340 7 1 2 57419 38339
0 38341 5 1 1 38340
0 38342 7 3 2 52611 51226
0 38343 5 1 1 67686
0 38344 7 1 2 43465 67687
0 38345 5 1 1 38344
0 38346 7 1 2 62190 57906
0 38347 5 1 1 38346
0 38348 7 1 2 38345 38347
0 38349 5 1 1 38348
0 38350 7 1 2 66537 59819
0 38351 5 1 1 38350
0 38352 7 2 2 61604 58310
0 38353 5 1 1 67689
0 38354 7 1 2 44566 67690
0 38355 5 1 1 38354
0 38356 7 1 2 38351 38355
0 38357 5 1 1 38356
0 38358 7 1 2 38349 38357
0 38359 5 1 1 38358
0 38360 7 1 2 59820 62201
0 38361 5 1 1 38360
0 38362 7 1 2 38361 38353
0 38363 5 1 1 38362
0 38364 7 1 2 66221 57907
0 38365 5 1 1 38364
0 38366 7 1 2 48619 67688
0 38367 5 1 1 38366
0 38368 7 1 2 38365 38367
0 38369 5 1 1 38368
0 38370 7 1 2 38363 38369
0 38371 5 1 1 38370
0 38372 7 1 2 61135 57908
0 38373 5 1 1 38372
0 38374 7 1 2 38343 38373
0 38375 5 1 1 38374
0 38376 7 1 2 59821 67549
0 38377 5 1 1 38376
0 38378 7 1 2 38377 10219
0 38379 5 1 1 38378
0 38380 7 1 2 49903 38379
0 38381 7 1 2 38375 38380
0 38382 5 1 1 38381
0 38383 7 1 2 38371 38382
0 38384 7 1 2 38359 38383
0 38385 7 1 2 38341 38384
0 38386 5 1 1 38385
0 38387 7 1 2 42003 38386
0 38388 5 1 1 38387
0 38389 7 1 2 38322 38388
0 38390 5 1 1 38389
0 38391 7 1 2 67637 38390
0 38392 5 1 1 38391
0 38393 7 1 2 58675 61194
0 38394 7 1 2 59914 50740
0 38395 7 1 2 38393 38394
0 38396 7 1 2 52764 67362
0 38397 7 1 2 38395 38396
0 38398 5 1 1 38397
0 38399 7 1 2 38392 38398
0 38400 7 1 2 38299 38399
0 38401 5 1 1 38400
0 38402 7 1 2 40696 38401
0 38403 5 1 1 38402
0 38404 7 1 2 63771 63425
0 38405 7 2 2 67608 38404
0 38406 5 1 1 67691
0 38407 7 1 2 45537 67692
0 38408 5 1 1 38407
0 38409 7 1 2 48134 65584
0 38410 5 1 1 38409
0 38411 7 1 2 38410 55360
0 38412 5 1 1 38411
0 38413 7 1 2 65991 38412
0 38414 5 1 1 38413
0 38415 7 1 2 64513 52502
0 38416 7 1 2 56947 38415
0 38417 5 1 1 38416
0 38418 7 1 2 38414 38417
0 38419 5 1 1 38418
0 38420 7 1 2 49234 38419
0 38421 5 1 1 38420
0 38422 7 1 2 45538 67604
0 38423 5 1 1 38422
0 38424 7 1 2 55780 56135
0 38425 7 1 2 60767 38424
0 38426 5 1 1 38425
0 38427 7 1 2 38423 38426
0 38428 5 1 1 38427
0 38429 7 1 2 65591 38428
0 38430 5 1 1 38429
0 38431 7 1 2 57315 56638
0 38432 7 1 2 64011 38431
0 38433 5 1 1 38432
0 38434 7 1 2 38430 38433
0 38435 7 1 2 38421 38434
0 38436 5 1 1 38435
0 38437 7 1 2 67638 38436
0 38438 5 1 1 38437
0 38439 7 1 2 38408 38438
0 38440 5 1 1 38439
0 38441 7 1 2 47505 38440
0 38442 5 1 1 38441
0 38443 7 1 2 51227 60661
0 38444 5 1 1 38443
0 38445 7 1 2 57689 51403
0 38446 7 1 2 56228 38445
0 38447 5 1 1 38446
0 38448 7 1 2 38444 38447
0 38449 5 1 1 38448
0 38450 7 1 2 40895 38449
0 38451 5 1 1 38450
0 38452 7 1 2 53218 57035
0 38453 7 1 2 56453 38452
0 38454 5 1 1 38453
0 38455 7 1 2 38451 38454
0 38456 5 1 1 38455
0 38457 7 1 2 43048 38456
0 38458 5 1 1 38457
0 38459 7 1 2 55402 64635
0 38460 5 1 1 38459
0 38461 7 1 2 38458 38460
0 38462 5 1 1 38461
0 38463 7 1 2 40697 38462
0 38464 5 1 1 38463
0 38465 7 1 2 49235 66590
0 38466 5 1 1 38465
0 38467 7 1 2 65560 64021
0 38468 5 1 1 38467
0 38469 7 1 2 38466 38468
0 38470 5 1 1 38469
0 38471 7 1 2 56371 54689
0 38472 7 1 2 38470 38471
0 38473 5 1 1 38472
0 38474 7 1 2 38464 38473
0 38475 5 1 1 38474
0 38476 7 1 2 46536 57667
0 38477 7 1 2 47302 62243
0 38478 7 1 2 38476 38477
0 38479 7 1 2 38475 38478
0 38480 5 1 1 38479
0 38481 7 1 2 38442 38480
0 38482 5 1 1 38481
0 38483 7 1 2 45358 38482
0 38484 5 1 1 38483
0 38485 7 1 2 60583 63959
0 38486 5 1 1 38485
0 38487 7 1 2 54199 57343
0 38488 5 1 1 38487
0 38489 7 1 2 38486 38488
0 38490 5 1 1 38489
0 38491 7 1 2 65585 38490
0 38492 5 1 1 38491
0 38493 7 1 2 37447 38492
0 38494 5 1 1 38493
0 38495 7 1 2 54571 67639
0 38496 7 1 2 38494 38495
0 38497 5 1 1 38496
0 38498 7 1 2 38484 38497
0 38499 5 1 1 38498
0 38500 7 1 2 47827 38499
0 38501 5 1 1 38500
0 38502 7 1 2 40698 67666
0 38503 5 1 1 38502
0 38504 7 1 2 66133 67668
0 38505 7 1 2 62862 38504
0 38506 5 1 1 38505
0 38507 7 1 2 38503 38506
0 38508 5 1 1 38507
0 38509 7 1 2 67156 38508
0 38510 5 1 1 38509
0 38511 7 1 2 45138 58687
0 38512 7 1 2 62194 38511
0 38513 7 1 2 65595 38512
0 38514 7 1 2 67652 38513
0 38515 5 1 1 38514
0 38516 7 1 2 38510 38515
0 38517 5 1 1 38516
0 38518 7 1 2 48285 38517
0 38519 5 1 1 38518
0 38520 7 5 2 54285 56358
0 38521 7 1 2 67693 61627
0 38522 5 1 1 38521
0 38523 7 1 2 54992 57165
0 38524 5 1 1 38523
0 38525 7 1 2 38522 38524
0 38526 5 1 1 38525
0 38527 7 1 2 42203 38526
0 38528 5 1 1 38527
0 38529 7 1 2 66542 62427
0 38530 5 1 1 38529
0 38531 7 1 2 38528 38530
0 38532 5 1 1 38531
0 38533 7 1 2 49904 38532
0 38534 5 1 1 38533
0 38535 7 1 2 54993 67497
0 38536 7 1 2 62422 38535
0 38537 5 1 1 38536
0 38538 7 1 2 54286 67122
0 38539 7 1 2 66833 38538
0 38540 5 1 1 38539
0 38541 7 1 2 38537 38540
0 38542 7 1 2 38534 38541
0 38543 5 1 1 38542
0 38544 7 1 2 67640 38543
0 38545 5 1 1 38544
0 38546 7 2 2 52191 51495
0 38547 7 1 2 57072 67698
0 38548 5 1 1 38547
0 38549 7 1 2 57964 61195
0 38550 7 1 2 66910 38549
0 38551 5 1 1 38550
0 38552 7 1 2 38548 38551
0 38553 5 1 1 38552
0 38554 7 1 2 47681 38553
0 38555 5 1 1 38554
0 38556 7 2 2 57020 51438
0 38557 7 2 2 66540 67700
0 38558 7 1 2 51793 67702
0 38559 5 1 1 38558
0 38560 7 1 2 38555 38559
0 38561 5 1 1 38560
0 38562 7 1 2 67641 38561
0 38563 5 1 1 38562
0 38564 7 1 2 59208 52195
0 38565 7 1 2 67090 67439
0 38566 7 1 2 38564 38565
0 38567 5 1 1 38566
0 38568 7 1 2 38563 38567
0 38569 5 1 1 38568
0 38570 7 1 2 47364 38569
0 38571 5 1 1 38570
0 38572 7 1 2 67649 67699
0 38573 5 1 1 38572
0 38574 7 1 2 43809 50460
0 38575 5 1 1 38574
0 38576 7 1 2 51386 38575
0 38577 5 1 1 38576
0 38578 7 1 2 67642 67694
0 38579 7 1 2 38577 38578
0 38580 5 1 1 38579
0 38581 7 1 2 38573 38580
0 38582 5 1 1 38581
0 38583 7 1 2 54200 38582
0 38584 5 1 1 38583
0 38585 7 1 2 41769 64387
0 38586 7 1 2 52196 38585
0 38587 7 1 2 67658 56912
0 38588 7 1 2 38586 38587
0 38589 5 1 1 38588
0 38590 7 1 2 38584 38589
0 38591 5 1 1 38590
0 38592 7 1 2 47682 38591
0 38593 5 1 1 38592
0 38594 7 1 2 52612 59188
0 38595 7 1 2 62335 38594
0 38596 7 1 2 66538 67363
0 38597 7 1 2 38595 38596
0 38598 5 1 1 38597
0 38599 7 1 2 38593 38598
0 38600 7 1 2 38571 38599
0 38601 7 1 2 38545 38600
0 38602 5 1 1 38601
0 38603 7 1 2 40699 38602
0 38604 5 1 1 38603
0 38605 7 1 2 66134 62305
0 38606 7 1 2 67634 38605
0 38607 7 1 2 67703 38606
0 38608 5 1 1 38607
0 38609 7 1 2 38604 38608
0 38610 5 1 1 38609
0 38611 7 1 2 52946 38610
0 38612 5 1 1 38611
0 38613 7 1 2 38519 38612
0 38614 7 1 2 38501 38613
0 38615 7 1 2 54201 60436
0 38616 5 1 1 38615
0 38617 7 1 2 65874 38616
0 38618 5 1 1 38617
0 38619 7 1 2 38618 59163
0 38620 5 1 1 38619
0 38621 7 1 2 62468 55699
0 38622 7 1 2 49253 38621
0 38623 5 1 1 38622
0 38624 7 1 2 38620 38623
0 38625 5 1 1 38624
0 38626 7 1 2 67650 38625
0 38627 5 1 1 38626
0 38628 7 1 2 49254 67662
0 38629 7 1 2 67294 38628
0 38630 5 1 1 38629
0 38631 7 1 2 38627 38630
0 38632 5 1 1 38631
0 38633 7 1 2 46318 38632
0 38634 5 1 1 38633
0 38635 7 1 2 54202 58442
0 38636 5 1 1 38635
0 38637 7 1 2 65875 38636
0 38638 5 1 1 38637
0 38639 7 1 2 49905 38638
0 38640 5 1 1 38639
0 38641 7 1 2 54203 50308
0 38642 5 1 1 38641
0 38643 7 1 2 43810 58449
0 38644 5 1 1 38643
0 38645 7 1 2 51387 38644
0 38646 5 1 1 38645
0 38647 7 1 2 54107 38646
0 38648 5 1 1 38647
0 38649 7 1 2 60632 38648
0 38650 5 1 1 38649
0 38651 7 1 2 47683 38650
0 38652 5 1 1 38651
0 38653 7 1 2 38642 38652
0 38654 7 1 2 38640 38653
0 38655 5 1 1 38654
0 38656 7 1 2 46537 63317
0 38657 7 1 2 63087 38656
0 38658 7 1 2 38655 38657
0 38659 5 1 1 38658
0 38660 7 1 2 38634 38659
0 38661 5 1 1 38660
0 38662 7 1 2 44835 38661
0 38663 5 1 1 38662
0 38664 7 1 2 50187 51491
0 38665 7 1 2 65681 38664
0 38666 7 1 2 67670 38665
0 38667 5 1 1 38666
0 38668 7 1 2 38663 38667
0 38669 5 1 1 38668
0 38670 7 1 2 54830 38669
0 38671 5 1 1 38670
0 38672 7 1 2 57840 48286
0 38673 5 2 1 38672
0 38674 7 1 2 48245 64078
0 38675 5 2 1 38674
0 38676 7 1 2 48196 67706
0 38677 5 1 1 38676
0 38678 7 1 2 54020 38677
0 38679 5 1 1 38678
0 38680 7 1 2 67704 38679
0 38681 5 1 1 38680
0 38682 7 1 2 40896 38681
0 38683 5 1 1 38682
0 38684 7 1 2 30039 67582
0 38685 5 1 1 38684
0 38686 7 1 2 38683 38685
0 38687 5 1 1 38686
0 38688 7 1 2 49621 38687
0 38689 5 1 1 38688
0 38690 7 1 2 40129 64639
0 38691 5 1 1 38690
0 38692 7 1 2 60213 49989
0 38693 7 1 2 58644 38692
0 38694 5 1 1 38693
0 38695 7 1 2 37697 38694
0 38696 7 1 2 38691 38695
0 38697 5 1 1 38696
0 38698 7 1 2 42896 38697
0 38699 5 1 1 38698
0 38700 7 1 2 57084 57843
0 38701 5 1 1 38700
0 38702 7 1 2 48135 49236
0 38703 7 1 2 38701 38702
0 38704 5 1 1 38703
0 38705 7 1 2 38699 38704
0 38706 5 1 1 38705
0 38707 7 1 2 48527 38706
0 38708 5 1 1 38707
0 38709 7 1 2 38689 38708
0 38710 5 1 1 38709
0 38711 7 1 2 42728 38710
0 38712 5 1 1 38711
0 38713 7 1 2 57087 48287
0 38714 5 1 1 38713
0 38715 7 1 2 66469 38714
0 38716 5 1 1 38715
0 38717 7 1 2 44151 38716
0 38718 5 1 1 38717
0 38719 7 1 2 63845 48446
0 38720 7 1 2 67551 38719
0 38721 5 1 1 38720
0 38722 7 1 2 38718 38721
0 38723 5 1 1 38722
0 38724 7 1 2 65586 38723
0 38725 5 1 1 38724
0 38726 7 1 2 49622 67580
0 38727 5 1 1 38726
0 38728 7 1 2 67585 57697
0 38729 5 1 1 38728
0 38730 7 1 2 67110 38729
0 38731 5 1 1 38730
0 38732 7 1 2 54204 38731
0 38733 5 1 1 38732
0 38734 7 1 2 38727 38733
0 38735 5 1 1 38734
0 38736 7 1 2 42729 38735
0 38737 5 1 1 38736
0 38738 7 1 2 38725 38737
0 38739 5 1 1 38738
0 38740 7 1 2 46769 38739
0 38741 5 1 1 38740
0 38742 7 1 2 63450 67707
0 38743 5 1 1 38742
0 38744 7 1 2 54021 38743
0 38745 5 1 1 38744
0 38746 7 1 2 67705 38745
0 38747 5 1 1 38746
0 38748 7 1 2 44152 38747
0 38749 5 1 1 38748
0 38750 7 1 2 54022 52716
0 38751 5 1 1 38750
0 38752 7 1 2 67601 38751
0 38753 5 1 1 38752
0 38754 7 1 2 61967 38753
0 38755 5 1 1 38754
0 38756 7 1 2 38749 38755
0 38757 5 1 1 38756
0 38758 7 1 2 65544 38757
0 38759 5 1 1 38758
0 38760 7 1 2 38741 38759
0 38761 7 1 2 38712 38760
0 38762 5 1 1 38761
0 38763 7 1 2 67643 38762
0 38764 5 1 1 38763
0 38765 7 1 2 38406 38764
0 38766 5 1 1 38765
0 38767 7 1 2 45539 50215
0 38768 7 1 2 38766 38767
0 38769 5 1 1 38768
0 38770 7 1 2 38671 38769
0 38771 7 1 2 38614 38770
0 38772 7 1 2 38403 38771
0 38773 7 1 2 38205 38772
0 38774 5 1 1 38773
0 38775 7 1 2 46600 38774
0 38776 5 1 1 38775
0 38777 7 1 2 60060 67276
0 38778 7 1 2 62115 38777
0 38779 5 1 1 38778
0 38780 7 1 2 61595 38779
0 38781 5 1 1 38780
0 38782 7 1 2 47748 38781
0 38783 5 1 1 38782
0 38784 7 1 2 41282 61641
0 38785 5 1 1 38784
0 38786 7 1 2 61596 38785
0 38787 5 1 1 38786
0 38788 7 1 2 43811 38787
0 38789 5 1 1 38788
0 38790 7 1 2 38783 38789
0 38791 5 1 1 38790
0 38792 7 1 2 47365 38791
0 38793 5 1 1 38792
0 38794 7 1 2 50216 55921
0 38795 7 1 2 61232 38794
0 38796 5 1 1 38795
0 38797 7 1 2 54205 38796
0 38798 5 1 1 38797
0 38799 7 1 2 37499 38798
0 38800 5 1 1 38799
0 38801 7 1 2 59493 38800
0 38802 5 1 1 38801
0 38803 7 1 2 53932 62248
0 38804 7 1 2 67528 38803
0 38805 5 1 1 38804
0 38806 7 1 2 38802 38805
0 38807 7 1 2 38793 38806
0 38808 5 1 1 38807
0 38809 7 1 2 67695 38808
0 38810 5 1 1 38809
0 38811 7 1 2 67120 61271
0 38812 5 1 1 38811
0 38813 7 1 2 38812 62047
0 38814 5 1 1 38813
0 38815 7 1 2 60035 67624
0 38816 5 1 1 38815
0 38817 7 1 2 40532 38816
0 38818 5 1 1 38817
0 38819 7 1 2 62042 38818
0 38820 5 1 1 38819
0 38821 7 1 2 49157 48797
0 38822 7 1 2 38820 38821
0 38823 5 1 1 38822
0 38824 7 1 2 38814 38823
0 38825 5 1 1 38824
0 38826 7 1 2 37075 60787
0 38827 5 1 1 38826
0 38828 7 1 2 45359 38827
0 38829 5 1 1 38828
0 38830 7 1 2 41283 62684
0 38831 5 1 1 38830
0 38832 7 1 2 48384 57073
0 38833 5 1 1 38832
0 38834 7 1 2 66730 38833
0 38835 5 1 1 38834
0 38836 7 1 2 44567 38835
0 38837 5 1 1 38836
0 38838 7 1 2 38831 38837
0 38839 7 1 2 38829 38838
0 38840 5 1 1 38839
0 38841 7 1 2 43812 38840
0 38842 5 1 1 38841
0 38843 7 1 2 62502 67557
0 38844 5 1 1 38843
0 38845 7 1 2 37123 38844
0 38846 7 1 2 38842 38845
0 38847 5 1 1 38846
0 38848 7 1 2 60314 38847
0 38849 5 1 1 38848
0 38850 7 1 2 38825 38849
0 38851 5 1 1 38850
0 38852 7 3 2 52613 51492
0 38853 7 1 2 38851 67708
0 38854 5 1 1 38853
0 38855 7 1 2 38810 38854
0 38856 5 1 1 38855
0 38857 7 1 2 42204 38856
0 38858 5 1 1 38857
0 38859 7 1 2 60519 59916
0 38860 7 1 2 63704 38859
0 38861 5 2 1 38860
0 38862 7 1 2 66225 58808
0 38863 7 1 2 61556 38862
0 38864 5 1 1 38863
0 38865 7 1 2 67711 38864
0 38866 5 1 1 38865
0 38867 7 1 2 43466 38866
0 38868 5 1 1 38867
0 38869 7 2 2 58676 67696
0 38870 7 1 2 46854 64592
0 38871 7 1 2 67713 38870
0 38872 5 1 1 38871
0 38873 7 1 2 38868 38872
0 38874 5 1 1 38873
0 38875 7 1 2 47684 38874
0 38876 5 1 1 38875
0 38877 7 1 2 58715 64593
0 38878 7 1 2 67714 38877
0 38879 5 1 1 38878
0 38880 7 1 2 38876 38879
0 38881 5 1 1 38880
0 38882 7 1 2 43813 38881
0 38883 5 1 1 38882
0 38884 7 1 2 46319 60100
0 38885 7 1 2 53091 49257
0 38886 7 1 2 38884 38885
0 38887 7 1 2 61622 61613
0 38888 7 1 2 38886 38887
0 38889 5 1 1 38888
0 38890 7 1 2 38883 38889
0 38891 7 1 2 38858 38890
0 38892 5 1 1 38891
0 38893 7 1 2 67380 38892
0 38894 5 1 1 38893
0 38895 7 1 2 63501 58338
0 38896 7 1 2 64420 38895
0 38897 7 1 2 67441 38896
0 38898 5 1 1 38897
0 38899 7 1 2 38894 38898
0 38900 5 1 1 38899
0 38901 7 1 2 40700 38900
0 38902 5 1 1 38901
0 38903 7 1 2 46954 54108
0 38904 5 1 1 38903
0 38905 7 1 2 54030 38904
0 38906 5 1 1 38905
0 38907 7 1 2 47506 38906
0 38908 5 1 1 38907
0 38909 7 1 2 61649 57769
0 38910 5 1 1 38909
0 38911 7 1 2 62007 38910
0 38912 7 1 2 38908 38911
0 38913 5 1 1 38912
0 38914 7 1 2 59390 67685
0 38915 7 1 2 38913 38914
0 38916 5 1 1 38915
0 38917 7 1 2 67712 38916
0 38918 5 1 1 38917
0 38919 7 1 2 44375 66135
0 38920 7 1 2 67576 38919
0 38921 7 1 2 38918 38920
0 38922 5 1 1 38921
0 38923 7 1 2 38902 38922
0 38924 5 1 1 38923
0 38925 7 1 2 52947 38924
0 38926 5 1 1 38925
0 38927 7 1 2 38776 38926
0 38928 7 1 2 63912 67572
0 38929 5 2 1 38928
0 38930 7 1 2 52503 67346
0 38931 5 1 1 38930
0 38932 7 1 2 42205 60796
0 38933 5 1 1 38932
0 38934 7 1 2 38931 38933
0 38935 5 1 1 38934
0 38936 7 1 2 46698 38935
0 38937 5 1 1 38936
0 38938 7 1 2 55842 56530
0 38939 5 1 1 38938
0 38940 7 1 2 38937 38939
0 38941 5 1 1 38940
0 38942 7 1 2 43979 38941
0 38943 5 1 1 38942
0 38944 7 1 2 67715 38943
0 38945 5 1 1 38944
0 38946 7 1 2 44836 38945
0 38947 5 1 1 38946
0 38948 7 1 2 55262 55843
0 38949 7 1 2 52146 38948
0 38950 5 2 1 38949
0 38951 7 1 2 38947 67717
0 38952 5 1 1 38951
0 38953 7 1 2 44153 38952
0 38954 5 1 1 38953
0 38955 7 1 2 44837 47961
0 38956 7 1 2 62910 38955
0 38957 7 1 2 60891 38956
0 38958 5 2 1 38957
0 38959 7 1 2 38954 67719
0 38960 5 1 1 38959
0 38961 7 1 2 60187 67682
0 38962 7 1 2 38960 38961
0 38963 5 1 1 38962
0 38964 7 4 2 48948 67655
0 38965 7 1 2 66552 51794
0 38966 5 1 1 38965
0 38967 7 1 2 50098 59885
0 38968 7 1 2 67431 38967
0 38969 5 1 1 38968
0 38970 7 1 2 38966 38969
0 38971 5 1 1 38970
0 38972 7 1 2 46320 38971
0 38973 5 1 1 38972
0 38974 7 2 2 67347 64005
0 38975 7 1 2 51463 67725
0 38976 5 1 1 38975
0 38977 7 1 2 38973 38976
0 38978 5 1 1 38977
0 38979 7 1 2 42897 38978
0 38980 5 1 1 38979
0 38981 7 1 2 59999 33309
0 38982 5 1 1 38981
0 38983 7 1 2 51077 38982
0 38984 5 1 1 38983
0 38985 7 1 2 55918 57431
0 38986 5 1 1 38985
0 38987 7 1 2 38984 38986
0 38988 5 1 1 38987
0 38989 7 1 2 47366 38988
0 38990 5 1 1 38989
0 38991 7 1 2 64022 58117
0 38992 5 1 1 38991
0 38993 7 1 2 61968 56084
0 38994 5 1 1 38993
0 38995 7 1 2 38992 38994
0 38996 5 1 1 38995
0 38997 7 1 2 47685 38996
0 38998 5 1 1 38997
0 38999 7 1 2 49906 63646
0 39000 5 1 1 38999
0 39001 7 1 2 50062 66252
0 39002 5 1 1 39001
0 39003 7 1 2 39000 39002
0 39004 5 1 1 39003
0 39005 7 1 2 42206 39004
0 39006 5 1 1 39005
0 39007 7 1 2 38998 39006
0 39008 7 1 2 38990 39007
0 39009 5 1 1 39008
0 39010 7 1 2 49967 39009
0 39011 5 1 1 39010
0 39012 7 1 2 38980 39011
0 39013 5 1 1 39012
0 39014 7 1 2 67721 39013
0 39015 5 1 1 39014
0 39016 7 1 2 48308 67340
0 39017 5 1 1 39016
0 39018 7 1 2 46178 60052
0 39019 7 1 2 58868 39018
0 39020 5 1 1 39019
0 39021 7 1 2 39017 39020
0 39022 5 1 1 39021
0 39023 7 1 2 62154 67364
0 39024 7 1 2 39022 39023
0 39025 5 1 1 39024
0 39026 7 1 2 39015 39025
0 39027 5 1 1 39026
0 39028 7 1 2 54375 39027
0 39029 5 1 1 39028
0 39030 7 1 2 47303 65572
0 39031 5 1 1 39030
0 39032 7 1 2 54335 47367
0 39033 5 1 1 39032
0 39034 7 1 2 47507 39033
0 39035 7 1 2 65575 39034
0 39036 5 1 1 39035
0 39037 7 1 2 39031 39036
0 39038 5 1 1 39037
0 39039 7 1 2 49237 39038
0 39040 5 1 1 39039
0 39041 7 1 2 64190 57715
0 39042 5 1 1 39041
0 39043 7 1 2 39040 39042
0 39044 5 1 1 39043
0 39045 7 1 2 51126 39044
0 39046 5 1 1 39045
0 39047 7 1 2 40701 55661
0 39048 5 1 1 39047
0 39049 7 1 2 45360 65573
0 39050 5 1 1 39049
0 39051 7 1 2 39048 39050
0 39052 5 1 1 39051
0 39053 7 1 2 49238 39052
0 39054 5 1 1 39053
0 39055 7 1 2 39054 64452
0 39056 5 1 1 39055
0 39057 7 1 2 50217 39056
0 39058 5 1 1 39057
0 39059 7 1 2 39046 39058
0 39060 5 1 1 39059
0 39061 7 1 2 58612 39060
0 39062 5 1 1 39061
0 39063 7 3 2 66939 57909
0 39064 7 1 2 47164 67727
0 39065 5 1 1 39064
0 39066 7 2 2 52614 57720
0 39067 5 1 1 67730
0 39068 7 1 2 46724 67731
0 39069 5 1 1 39068
0 39070 7 1 2 39065 39069
0 39071 5 1 1 39070
0 39072 7 1 2 43467 39071
0 39073 5 1 1 39072
0 39074 7 1 2 65419 67728
0 39075 5 1 1 39074
0 39076 7 1 2 39073 39075
0 39077 5 1 1 39076
0 39078 7 1 2 47686 39077
0 39079 5 1 1 39078
0 39080 7 1 2 47368 67729
0 39081 5 1 1 39080
0 39082 7 1 2 39067 39081
0 39083 5 1 1 39082
0 39084 7 1 2 55919 39083
0 39085 5 1 1 39084
0 39086 7 1 2 39079 39085
0 39087 7 1 2 39062 39086
0 39088 5 1 1 39087
0 39089 7 1 2 46179 39088
0 39090 5 1 1 39089
0 39091 7 1 2 41542 67726
0 39092 5 1 1 39091
0 39093 7 1 2 44838 51280
0 39094 7 1 2 67295 39093
0 39095 5 1 1 39094
0 39096 7 1 2 39092 39095
0 39097 5 1 1 39096
0 39098 7 1 2 40897 39097
0 39099 5 1 1 39098
0 39100 7 1 2 48606 57239
0 39101 7 1 2 67296 39100
0 39102 5 1 1 39101
0 39103 7 1 2 39099 39102
0 39104 5 1 1 39103
0 39105 7 1 2 43980 39104
0 39106 5 1 1 39105
0 39107 7 1 2 51281 56966
0 39108 7 1 2 67297 39107
0 39109 5 1 1 39108
0 39110 7 1 2 39106 39109
0 39111 5 1 1 39110
0 39112 7 1 2 55263 39111
0 39113 5 1 1 39112
0 39114 7 1 2 39090 39113
0 39115 5 1 1 39114
0 39116 7 1 2 67722 39115
0 39117 5 1 1 39116
0 39118 7 1 2 67323 67709
0 39119 5 1 1 39118
0 39120 7 1 2 49907 67697
0 39121 5 1 1 39120
0 39122 7 1 2 39119 39121
0 39123 5 1 1 39122
0 39124 7 1 2 67723 39123
0 39125 5 1 1 39124
0 39126 7 2 2 60188 67334
0 39127 7 1 2 67710 67732
0 39128 7 1 2 61786 39127
0 39129 5 1 1 39128
0 39130 7 1 2 39125 39129
0 39131 5 1 1 39130
0 39132 7 1 2 42207 39131
0 39133 5 1 1 39132
0 39134 7 1 2 52615 54883
0 39135 7 1 2 67365 39134
0 39136 7 1 2 62717 39135
0 39137 5 1 1 39136
0 39138 7 1 2 39133 39137
0 39139 5 1 1 39138
0 39140 7 1 2 40702 39139
0 39141 5 1 1 39140
0 39142 7 2 2 67139 67432
0 39143 7 1 2 49271 66911
0 39144 7 1 2 67656 39143
0 39145 7 1 2 67734 39144
0 39146 5 1 1 39145
0 39147 7 1 2 39141 39146
0 39148 5 1 1 39147
0 39149 7 1 2 52948 39148
0 39150 5 1 1 39149
0 39151 7 1 2 49908 48288
0 39152 5 1 1 39151
0 39153 7 1 2 51646 60429
0 39154 5 1 1 39153
0 39155 7 1 2 39152 39154
0 39156 5 1 1 39155
0 39157 7 1 2 50960 39156
0 39158 5 1 1 39157
0 39159 7 1 2 42898 49137
0 39160 7 1 2 67735 39159
0 39161 5 1 1 39160
0 39162 7 1 2 39158 39161
0 39163 5 1 1 39162
0 39164 7 1 2 67724 39163
0 39165 5 1 1 39164
0 39166 7 1 2 40703 48289
0 39167 7 1 2 67733 39166
0 39168 7 1 2 67341 39167
0 39169 5 1 1 39168
0 39170 7 1 2 39165 39169
0 39171 5 1 1 39170
0 39172 7 1 2 67157 39171
0 39173 5 1 1 39172
0 39174 7 1 2 39150 39173
0 39175 7 1 2 39117 39174
0 39176 7 1 2 39029 39175
0 39177 7 1 2 38963 39176
0 39178 5 1 1 39177
0 39179 7 1 2 46601 39178
0 39180 5 1 1 39179
0 39181 7 1 2 57604 67412
0 39182 5 1 1 39181
0 39183 7 1 2 57544 52301
0 39184 5 1 1 39183
0 39185 7 1 2 39182 39184
0 39186 5 1 1 39185
0 39187 7 1 2 61677 39186
0 39188 5 1 1 39187
0 39189 7 1 2 40533 47207
0 39190 5 1 1 39189
0 39191 7 1 2 58296 39190
0 39192 5 1 1 39191
0 39193 7 1 2 40306 39192
0 39194 5 1 1 39193
0 39195 7 1 2 40534 58384
0 39196 5 1 1 39195
0 39197 7 1 2 39194 39196
0 39198 5 2 1 39197
0 39199 7 1 2 58647 62945
0 39200 7 1 2 67736 39199
0 39201 5 1 1 39200
0 39202 7 1 2 39188 39201
0 39203 5 1 1 39202
0 39204 7 1 2 44982 39203
0 39205 5 1 1 39204
0 39206 7 1 2 58437 61750
0 39207 5 1 1 39206
0 39208 7 1 2 33526 39207
0 39209 5 1 1 39208
0 39210 7 1 2 47828 39209
0 39211 5 1 1 39210
0 39212 7 1 2 65066 58450
0 39213 5 1 1 39212
0 39214 7 1 2 61751 39213
0 39215 5 1 1 39214
0 39216 7 1 2 39211 39215
0 39217 5 1 1 39216
0 39218 7 1 2 40535 39217
0 39219 5 1 1 39218
0 39220 7 3 2 45065 57219
0 39221 7 1 2 50447 67738
0 39222 7 1 2 65858 39221
0 39223 5 1 1 39222
0 39224 7 1 2 39219 39223
0 39225 5 1 1 39224
0 39226 7 1 2 52616 47234
0 39227 7 1 2 39225 39226
0 39228 5 1 1 39227
0 39229 7 1 2 39205 39228
0 39230 5 1 1 39229
0 39231 7 1 2 40898 39230
0 39232 5 1 1 39231
0 39233 7 1 2 54476 67737
0 39234 5 1 1 39233
0 39235 7 1 2 54049 47249
0 39236 5 1 1 39235
0 39237 7 1 2 36224 39236
0 39238 5 1 1 39237
0 39239 7 1 2 53725 39238
0 39240 5 1 1 39239
0 39241 7 1 2 54706 47255
0 39242 5 1 1 39241
0 39243 7 1 2 43814 67398
0 39244 5 1 1 39243
0 39245 7 1 2 39242 39244
0 39246 7 1 2 39240 39245
0 39247 5 1 1 39246
0 39248 7 1 2 54507 39247
0 39249 5 1 1 39248
0 39250 7 1 2 39234 39249
0 39251 5 1 1 39250
0 39252 7 1 2 61752 39251
0 39253 5 1 1 39252
0 39254 7 1 2 53933 54477
0 39255 7 1 2 67429 39254
0 39256 5 1 1 39255
0 39257 7 1 2 39253 39256
0 39258 5 1 1 39257
0 39259 7 1 2 48290 39258
0 39260 5 1 1 39259
0 39261 7 1 2 44568 53569
0 39262 5 1 1 39261
0 39263 7 1 2 56316 39262
0 39264 5 1 1 39263
0 39265 7 1 2 43815 39264
0 39266 5 1 1 39265
0 39267 7 1 2 51708 54707
0 39268 5 1 1 39267
0 39269 7 1 2 39266 39268
0 39270 5 1 1 39269
0 39271 7 1 2 47235 61753
0 39272 7 1 2 39270 39271
0 39273 5 1 1 39272
0 39274 7 1 2 44569 63585
0 39275 5 1 1 39274
0 39276 7 2 2 57220 62360
0 39277 5 2 1 67741
0 39278 7 1 2 61689 67743
0 39279 5 2 1 39278
0 39280 7 4 2 59978 62698
0 39281 5 1 1 67747
0 39282 7 1 2 40307 39281
0 39283 5 1 1 39282
0 39284 7 1 2 67745 39283
0 39285 5 1 1 39284
0 39286 7 1 2 39275 39285
0 39287 5 1 1 39286
0 39288 7 1 2 42208 39287
0 39289 5 1 1 39288
0 39290 7 1 2 50706 67742
0 39291 5 1 1 39290
0 39292 7 1 2 61678 51101
0 39293 5 1 1 39292
0 39294 7 1 2 39291 39293
0 39295 5 1 1 39294
0 39296 7 1 2 47369 39295
0 39297 5 2 1 39296
0 39298 7 1 2 61679 58316
0 39299 5 1 1 39298
0 39300 7 1 2 67751 39299
0 39301 7 1 2 39289 39300
0 39302 5 1 1 39301
0 39303 7 1 2 43816 39302
0 39304 5 1 1 39303
0 39305 7 1 2 64880 61754
0 39306 5 1 1 39305
0 39307 7 1 2 61690 39306
0 39308 5 1 1 39307
0 39309 7 1 2 39308 51267
0 39310 5 2 1 39309
0 39311 7 1 2 51712 51806
0 39312 5 1 1 39311
0 39313 7 1 2 67748 39312
0 39314 5 1 1 39313
0 39315 7 1 2 67753 39314
0 39316 7 1 2 39304 39315
0 39317 7 1 2 39273 39316
0 39318 5 1 1 39317
0 39319 7 1 2 42730 67583
0 39320 7 1 2 39318 39319
0 39321 5 1 1 39320
0 39322 7 1 2 39260 39321
0 39323 7 1 2 39232 39322
0 39324 5 1 1 39323
0 39325 7 1 2 58063 39324
0 39326 5 1 1 39325
0 39327 7 2 2 50633 54482
0 39328 7 1 2 40130 67755
0 39329 5 1 1 39328
0 39330 7 1 2 45540 57445
0 39331 5 1 1 39330
0 39332 7 1 2 39329 39331
0 39333 5 1 1 39332
0 39334 7 1 2 47829 39333
0 39335 5 1 1 39334
0 39336 7 1 2 56198 67756
0 39337 5 1 1 39336
0 39338 7 1 2 39335 39337
0 39339 5 1 1 39338
0 39340 7 1 2 61680 39339
0 39341 5 1 1 39340
0 39342 7 1 2 57394 64486
0 39343 5 1 1 39342
0 39344 7 1 2 66883 39343
0 39345 5 1 1 39344
0 39346 7 1 2 47830 47169
0 39347 7 1 2 39345 39346
0 39348 5 1 1 39347
0 39349 7 1 2 49131 66889
0 39350 5 1 1 39349
0 39351 7 1 2 66884 39350
0 39352 5 1 1 39351
0 39353 7 1 2 47687 9802
0 39354 5 1 1 39353
0 39355 7 1 2 39352 39354
0 39356 5 1 1 39355
0 39357 7 1 2 45541 57295
0 39358 7 1 2 57520 39357
0 39359 7 1 2 533 39358
0 39360 5 1 1 39359
0 39361 7 1 2 39356 39360
0 39362 7 1 2 39348 39361
0 39363 7 1 2 39341 39362
0 39364 5 1 1 39363
0 39365 7 1 2 40536 39364
0 39366 5 1 1 39365
0 39367 7 1 2 46770 66881
0 39368 5 1 1 39367
0 39369 7 1 2 57765 51475
0 39370 7 1 2 66890 39369
0 39371 5 1 1 39370
0 39372 7 1 2 39368 39371
0 39373 5 1 1 39372
0 39374 7 1 2 40131 39373
0 39375 5 1 1 39374
0 39376 7 1 2 57870 57969
0 39377 7 1 2 51448 39376
0 39378 5 1 1 39377
0 39379 7 1 2 39375 39378
0 39380 5 1 1 39379
0 39381 7 1 2 58244 39380
0 39382 5 1 1 39381
0 39383 7 1 2 39366 39382
0 39384 5 1 1 39383
0 39385 7 1 2 52949 39384
0 39386 5 1 1 39385
0 39387 7 1 2 42004 67744
0 39388 5 1 1 39387
0 39389 7 1 2 67746 64501
0 39390 7 1 2 39388 39389
0 39391 5 1 1 39390
0 39392 7 1 2 57280 51341
0 39393 7 1 2 56129 39392
0 39394 5 1 1 39393
0 39395 7 1 2 39391 39394
0 39396 5 1 1 39395
0 39397 7 1 2 57446 39396
0 39398 5 1 1 39397
0 39399 7 1 2 45361 66898
0 39400 5 1 1 39399
0 39401 7 3 2 63541 63710
0 39402 7 1 2 63489 58956
0 39403 7 1 2 67757 39402
0 39404 5 1 1 39403
0 39405 7 1 2 39400 39404
0 39406 5 1 1 39405
0 39407 7 1 2 47137 39406
0 39408 5 1 1 39407
0 39409 7 1 2 44839 52777
0 39410 7 1 2 55563 39409
0 39411 7 1 2 67758 39410
0 39412 5 1 1 39411
0 39413 7 1 2 39408 39412
0 39414 7 1 2 39398 39413
0 39415 5 1 1 39414
0 39416 7 1 2 40537 39415
0 39417 5 1 1 39416
0 39418 7 1 2 53335 51098
0 39419 7 1 2 52717 39418
0 39420 7 1 2 63440 39419
0 39421 5 1 1 39420
0 39422 7 1 2 39417 39421
0 39423 5 1 1 39422
0 39424 7 1 2 47508 39423
0 39425 5 1 1 39424
0 39426 7 1 2 47304 66903
0 39427 5 1 1 39426
0 39428 7 1 2 63778 66463
0 39429 7 1 2 52839 39428
0 39430 5 1 1 39429
0 39431 7 1 2 39427 39430
0 39432 5 1 1 39431
0 39433 7 1 2 50218 39432
0 39434 5 1 1 39433
0 39435 7 1 2 62525 63542
0 39436 7 1 2 67701 39435
0 39437 5 1 1 39436
0 39438 7 1 2 57775 63071
0 39439 7 1 2 63441 39438
0 39440 5 1 1 39439
0 39441 7 1 2 39437 39440
0 39442 5 1 1 39441
0 39443 7 1 2 51127 39442
0 39444 5 1 1 39443
0 39445 7 1 2 60198 63428
0 39446 5 1 1 39445
0 39447 7 1 2 39444 39446
0 39448 5 1 1 39447
0 39449 7 1 2 47236 39448
0 39450 5 1 1 39449
0 39451 7 1 2 39434 39450
0 39452 5 1 1 39451
0 39453 7 1 2 45542 39452
0 39454 5 1 1 39453
0 39455 7 1 2 50110 50644
0 39456 7 1 2 63421 39455
0 39457 7 1 2 57155 39456
0 39458 7 1 2 62485 39457
0 39459 5 1 1 39458
0 39460 7 1 2 40308 66896
0 39461 7 1 2 64749 39460
0 39462 5 1 1 39461
0 39463 7 1 2 39459 39462
0 39464 5 1 1 39463
0 39465 7 1 2 40538 39464
0 39466 5 1 1 39465
0 39467 7 1 2 42731 39466
0 39468 7 1 2 39454 39467
0 39469 7 1 2 39425 39468
0 39470 7 1 2 39386 39469
0 39471 5 1 1 39470
0 39472 7 2 2 57296 57521
0 39473 7 1 2 50883 67760
0 39474 5 1 1 39473
0 39475 7 1 2 66885 39474
0 39476 5 1 1 39475
0 39477 7 1 2 47688 39476
0 39478 5 1 1 39477
0 39479 7 2 2 57395 51631
0 39480 7 1 2 53325 62429
0 39481 7 1 2 67762 39480
0 39482 5 1 1 39481
0 39483 7 1 2 66886 39482
0 39484 5 1 1 39483
0 39485 7 1 2 42209 39484
0 39486 5 1 1 39485
0 39487 7 1 2 39478 39486
0 39488 5 1 1 39487
0 39489 7 1 2 43817 39488
0 39490 5 1 1 39489
0 39491 7 1 2 64625 66972
0 39492 7 1 2 67763 39491
0 39493 5 1 1 39492
0 39494 7 1 2 66887 39493
0 39495 5 1 1 39494
0 39496 7 1 2 54758 39495
0 39497 5 1 1 39496
0 39498 7 1 2 39490 39497
0 39499 5 1 1 39498
0 39500 7 1 2 47370 39499
0 39501 5 1 1 39500
0 39502 7 1 2 53345 57108
0 39503 7 2 2 60520 39502
0 39504 7 1 2 43611 67764
0 39505 5 1 1 39504
0 39506 7 1 2 60982 62430
0 39507 7 1 2 66891 39506
0 39508 5 1 1 39507
0 39509 7 1 2 39505 39508
0 39510 5 1 1 39509
0 39511 7 1 2 47438 39510
0 39512 5 1 1 39511
0 39513 7 1 2 65995 56484
0 39514 7 1 2 67487 39513
0 39515 5 1 1 39514
0 39516 7 1 2 39512 39515
0 39517 5 1 1 39516
0 39518 7 1 2 47060 39517
0 39519 5 1 1 39518
0 39520 7 1 2 67399 67761
0 39521 5 1 1 39520
0 39522 7 1 2 56051 57970
0 39523 7 1 2 58510 39522
0 39524 5 1 1 39523
0 39525 7 1 2 39521 39524
0 39526 5 1 1 39525
0 39527 7 1 2 43818 39526
0 39528 5 1 1 39527
0 39529 7 1 2 49695 67765
0 39530 5 1 1 39529
0 39531 7 1 2 63232 62431
0 39532 7 1 2 66892 39531
0 39533 5 1 1 39532
0 39534 7 1 2 39530 39533
0 39535 7 1 2 39528 39534
0 39536 5 1 1 39535
0 39537 7 1 2 47156 39536
0 39538 5 1 1 39537
0 39539 7 1 2 39519 39538
0 39540 7 1 2 39501 39539
0 39541 5 1 1 39540
0 39542 7 1 2 52950 39541
0 39543 5 1 1 39542
0 39544 7 2 2 61755 64166
0 39545 7 2 2 42210 67766
0 39546 7 1 2 66738 49260
0 39547 5 1 1 39546
0 39548 7 1 2 47439 47237
0 39549 5 2 1 39548
0 39550 7 1 2 39547 67770
0 39551 5 1 1 39550
0 39552 7 1 2 45362 39551
0 39553 5 1 1 39552
0 39554 7 1 2 50772 66817
0 39555 5 1 1 39554
0 39556 7 1 2 49781 47238
0 39557 5 1 1 39556
0 39558 7 1 2 46944 57113
0 39559 5 1 1 39558
0 39560 7 1 2 39557 39559
0 39561 5 1 1 39560
0 39562 7 1 2 44570 39561
0 39563 5 1 1 39562
0 39564 7 1 2 39555 39563
0 39565 7 1 2 39553 39564
0 39566 5 1 1 39565
0 39567 7 1 2 67768 39566
0 39568 5 1 1 39567
0 39569 7 1 2 42211 66899
0 39570 5 1 1 39569
0 39571 7 1 2 65153 51439
0 39572 7 1 2 47865 39571
0 39573 7 1 2 67759 39572
0 39574 5 1 1 39573
0 39575 7 1 2 39570 39574
0 39576 5 1 1 39575
0 39577 7 1 2 47689 39576
0 39578 5 1 1 39577
0 39579 7 2 2 60157 57447
0 39580 7 3 2 43278 67772
0 39581 7 1 2 47863 49287
0 39582 5 1 1 39581
0 39583 7 1 2 67774 39582
0 39584 5 1 1 39583
0 39585 7 1 2 39578 39584
0 39586 7 1 2 39568 39585
0 39587 5 1 1 39586
0 39588 7 1 2 43819 39587
0 39589 5 1 1 39588
0 39590 7 1 2 44454 52746
0 39591 5 1 1 39590
0 39592 7 1 2 7615 39591
0 39593 5 1 1 39592
0 39594 7 1 2 47690 39593
0 39595 5 1 1 39594
0 39596 7 1 2 49909 52704
0 39597 5 1 1 39596
0 39598 7 1 2 39595 39597
0 39599 5 1 1 39598
0 39600 7 1 2 67775 39599
0 39601 5 1 1 39600
0 39602 7 1 2 67518 58949
0 39603 7 1 2 63429 39602
0 39604 5 1 1 39603
0 39605 7 1 2 39601 39604
0 39606 5 1 1 39605
0 39607 7 1 2 49724 39606
0 39608 5 1 1 39607
0 39609 7 1 2 67435 63430
0 39610 5 1 1 39609
0 39611 7 1 2 67437 67773
0 39612 5 1 1 39611
0 39613 7 1 2 39610 39612
0 39614 5 1 1 39613
0 39615 7 1 2 67502 39614
0 39616 5 1 1 39615
0 39617 7 1 2 47157 54050
0 39618 7 1 2 62458 39617
0 39619 7 1 2 67767 39618
0 39620 5 1 1 39619
0 39621 7 1 2 36945 67776
0 39622 5 1 1 39621
0 39623 7 1 2 39620 39622
0 39624 7 1 2 39616 39623
0 39625 5 1 1 39624
0 39626 7 1 2 47869 39625
0 39627 5 1 1 39626
0 39628 7 1 2 67559 67769
0 39629 5 1 1 39628
0 39630 7 1 2 60594 53336
0 39631 7 1 2 63437 39630
0 39632 5 1 1 39631
0 39633 7 1 2 39629 39632
0 39634 5 1 1 39633
0 39635 7 1 2 47749 47866
0 39636 7 1 2 39634 39635
0 39637 5 1 1 39636
0 39638 7 1 2 46004 39637
0 39639 7 1 2 39627 39638
0 39640 7 1 2 39608 39639
0 39641 7 1 2 39589 39640
0 39642 7 1 2 39543 39641
0 39643 5 1 1 39642
0 39644 7 1 2 39471 39643
0 39645 5 1 1 39644
0 39646 7 1 2 40539 46864
0 39647 5 1 1 39646
0 39648 7 1 2 43612 39647
0 39649 5 1 1 39648
0 39650 7 1 2 46912 63610
0 39651 7 1 2 39649 39650
0 39652 5 1 1 39651
0 39653 7 1 2 63522 52780
0 39654 5 1 1 39653
0 39655 7 1 2 63621 63716
0 39656 5 1 1 39655
0 39657 7 1 2 49868 61756
0 39658 5 1 1 39657
0 39659 7 1 2 39656 39658
0 39660 5 1 1 39659
0 39661 7 1 2 46771 39660
0 39662 5 1 1 39661
0 39663 7 1 2 39654 39662
0 39664 7 1 2 39652 39663
0 39665 5 1 1 39664
0 39666 7 1 2 45543 39665
0 39667 5 1 1 39666
0 39668 7 1 2 47509 61681
0 39669 5 1 1 39668
0 39670 7 1 2 57770 67739
0 39671 5 1 1 39670
0 39672 7 1 2 39669 39671
0 39673 5 1 1 39672
0 39674 7 1 2 47831 39673
0 39675 5 1 1 39674
0 39676 7 1 2 62208 67740
0 39677 5 1 1 39676
0 39678 7 1 2 39675 39677
0 39679 5 1 1 39678
0 39680 7 1 2 45363 39679
0 39681 5 1 1 39680
0 39682 7 1 2 47510 61757
0 39683 5 1 1 39682
0 39684 7 1 2 61691 39683
0 39685 5 1 1 39684
0 39686 7 1 2 47603 39685
0 39687 5 1 1 39686
0 39688 7 1 2 39681 39687
0 39689 5 1 1 39688
0 39690 7 1 2 40540 39689
0 39691 5 1 1 39690
0 39692 7 1 2 42732 39691
0 39693 7 1 2 39667 39692
0 39694 5 1 1 39693
0 39695 7 1 2 59245 65863
0 39696 5 1 1 39695
0 39697 7 1 2 43613 67749
0 39698 5 1 1 39697
0 39699 7 1 2 39696 39698
0 39700 5 1 1 39699
0 39701 7 1 2 47440 39700
0 39702 5 1 1 39701
0 39703 7 1 2 52340 56055
0 39704 7 1 2 62107 39703
0 39705 5 1 1 39704
0 39706 7 1 2 39702 39705
0 39707 5 1 1 39706
0 39708 7 1 2 47061 39707
0 39709 5 1 1 39708
0 39710 7 1 2 61758 67400
0 39711 5 1 1 39710
0 39712 7 1 2 47105 61682
0 39713 5 1 1 39712
0 39714 7 1 2 43165 53726
0 39715 7 1 2 62946 54213
0 39716 7 1 2 39714 39715
0 39717 5 1 1 39716
0 39718 7 1 2 39713 39717
0 39719 7 1 2 39711 39718
0 39720 7 1 2 67752 39719
0 39721 5 1 1 39720
0 39722 7 1 2 43820 39721
0 39723 5 1 1 39722
0 39724 7 1 2 49696 67750
0 39725 5 1 1 39724
0 39726 7 1 2 47441 67483
0 39727 7 1 2 62947 39726
0 39728 5 1 1 39727
0 39729 7 1 2 39725 39728
0 39730 5 1 1 39729
0 39731 7 1 2 47158 39730
0 39732 5 1 1 39731
0 39733 7 1 2 46005 67754
0 39734 7 1 2 39732 39733
0 39735 7 1 2 39723 39734
0 39736 7 1 2 39709 39735
0 39737 5 1 1 39736
0 39738 7 1 2 57105 39737
0 39739 7 1 2 39694 39738
0 39740 5 1 1 39739
0 39741 7 1 2 39645 39740
0 39742 7 1 2 39326 39741
0 39743 5 1 1 39742
0 39744 7 1 2 67381 39743
0 39745 5 1 1 39744
0 39746 7 1 2 65288 67610
0 39747 7 1 2 51694 39746
0 39748 7 1 2 67538 39747
0 39749 5 1 1 39748
0 39750 7 1 2 39745 39749
0 39751 7 1 2 39180 39750
0 39752 5 1 1 39751
0 39753 7 1 2 55134 39752
0 39754 5 1 1 39753
0 39755 7 1 2 57990 63067
0 39756 7 1 2 67185 39755
0 39757 5 1 1 39756
0 39758 7 1 2 50839 65912
0 39759 7 1 2 67187 39758
0 39760 5 1 1 39759
0 39761 7 1 2 39757 39760
0 39762 5 1 1 39761
0 39763 7 1 2 40541 39762
0 39764 5 1 1 39763
0 39765 7 1 2 59408 59025
0 39766 7 1 2 65774 39765
0 39767 7 1 2 67477 39766
0 39768 5 1 1 39767
0 39769 7 1 2 39764 39768
0 39770 5 1 1 39769
0 39771 7 1 2 43981 39770
0 39772 5 1 1 39771
0 39773 7 1 2 52617 62010
0 39774 7 1 2 63191 39773
0 39775 7 1 2 52302 39774
0 39776 5 1 1 39775
0 39777 7 1 2 39772 39776
0 39778 5 1 1 39777
0 39779 7 1 2 41543 39778
0 39780 5 1 1 39779
0 39781 7 1 2 63920 51782
0 39782 5 1 1 39781
0 39783 7 1 2 54831 67543
0 39784 5 1 1 39783
0 39785 7 1 2 63496 63921
0 39786 5 1 1 39785
0 39787 7 1 2 39784 39786
0 39788 5 1 1 39787
0 39789 7 1 2 42212 39788
0 39790 5 1 1 39789
0 39791 7 1 2 60437 63922
0 39792 5 1 1 39791
0 39793 7 1 2 39790 39792
0 39794 5 1 1 39793
0 39795 7 1 2 43821 39794
0 39796 5 1 1 39795
0 39797 7 1 2 39782 39796
0 39798 5 1 1 39797
0 39799 7 1 2 50787 39798
0 39800 5 1 1 39799
0 39801 7 1 2 39780 39800
0 39802 5 1 1 39801
0 39803 7 1 2 44983 39802
0 39804 5 1 1 39803
0 39805 7 1 2 56004 59339
0 39806 7 1 2 67522 39805
0 39807 5 1 1 39806
0 39808 7 1 2 39804 39807
0 39809 5 1 1 39808
0 39810 7 1 2 40899 39809
0 39811 5 1 1 39810
0 39812 7 1 2 66591 51006
0 39813 5 1 1 39812
0 39814 7 1 2 52147 55203
0 39815 5 1 1 39814
0 39816 7 1 2 39813 39815
0 39817 5 1 1 39816
0 39818 7 1 2 59785 39817
0 39819 5 1 1 39818
0 39820 7 1 2 50376 58821
0 39821 7 1 2 67272 39820
0 39822 5 1 1 39821
0 39823 7 1 2 39819 39822
0 39824 5 1 1 39823
0 39825 7 1 2 54659 39824
0 39826 5 1 1 39825
0 39827 7 1 2 56005 56620
0 39828 5 1 1 39827
0 39829 7 1 2 65561 50099
0 39830 5 1 1 39829
0 39831 7 1 2 39828 39830
0 39832 5 1 1 39831
0 39833 7 1 2 67541 39832
0 39834 5 1 1 39833
0 39835 7 1 2 58064 50389
0 39836 7 1 2 58496 39835
0 39837 5 1 1 39836
0 39838 7 1 2 39834 39837
0 39839 5 1 1 39838
0 39840 7 1 2 46321 39839
0 39841 5 1 1 39840
0 39842 7 1 2 48528 50390
0 39843 7 1 2 62936 39842
0 39844 5 1 1 39843
0 39845 7 1 2 39841 39844
0 39846 5 1 1 39845
0 39847 7 1 2 43614 39846
0 39848 5 1 1 39847
0 39849 7 1 2 40704 66592
0 39850 5 1 1 39849
0 39851 7 1 2 58004 55204
0 39852 5 1 1 39851
0 39853 7 1 2 39850 39852
0 39854 5 2 1 39853
0 39855 7 1 2 63372 67777
0 39856 5 1 1 39855
0 39857 7 1 2 39848 39856
0 39858 5 1 1 39857
0 39859 7 1 2 54046 39858
0 39860 5 1 1 39859
0 39861 7 1 2 39826 39860
0 39862 5 1 1 39861
0 39863 7 1 2 41284 39862
0 39864 5 1 1 39863
0 39865 7 1 2 43822 65054
0 39866 5 1 1 39865
0 39867 7 1 2 67597 39866
0 39868 5 1 1 39867
0 39869 7 1 2 67778 39868
0 39870 5 1 1 39869
0 39871 7 1 2 46006 48246
0 39872 7 1 2 67391 39871
0 39873 7 1 2 66969 39872
0 39874 5 1 1 39873
0 39875 7 1 2 39870 39874
0 39876 5 1 1 39875
0 39877 7 1 2 41688 39876
0 39878 5 1 1 39877
0 39879 7 1 2 60983 67672
0 39880 7 1 2 66970 39879
0 39881 5 1 1 39880
0 39882 7 1 2 39878 39881
0 39883 5 1 1 39882
0 39884 7 1 2 47106 39883
0 39885 5 1 1 39884
0 39886 7 1 2 39864 39885
0 39887 5 1 1 39886
0 39888 7 1 2 39887 61948
0 39889 5 1 1 39888
0 39890 7 1 2 39811 39889
0 39891 5 1 1 39890
0 39892 7 1 2 67382 39891
0 39893 5 1 1 39892
0 39894 7 1 2 46699 60438
0 39895 5 1 1 39894
0 39896 7 1 2 67771 39895
0 39897 5 1 1 39896
0 39898 7 1 2 66201 39897
0 39899 5 1 1 39898
0 39900 7 1 2 67716 39899
0 39901 5 1 1 39900
0 39902 7 1 2 44840 39901
0 39903 5 1 1 39902
0 39904 7 1 2 67718 39903
0 39905 5 1 1 39904
0 39906 7 1 2 44154 39905
0 39907 5 1 1 39906
0 39908 7 1 2 67720 39907
0 39909 5 1 1 39908
0 39910 7 1 2 64421 67683
0 39911 7 1 2 39909 39910
0 39912 5 1 1 39911
0 39913 7 1 2 39893 39912
0 39914 5 1 1 39913
0 39915 7 1 2 54206 39914
0 39916 5 1 1 39915
0 39917 7 1 2 39754 39916
0 39918 7 1 2 38927 39917
0 39919 7 1 2 38078 39918
0 39920 7 1 2 37042 39919
0 39921 5 1 1 39920
0 39922 7 1 2 66819 39921
0 39923 5 1 1 39922
0 39924 7 1 2 35523 39923
0 39925 7 1 2 22685 39924
3 79999 5 0 1 39925
