1 0 0 2 0
2 64 1 0
2 65 1 0
1 1 0 2 0
2 66 1 1
2 67 1 1
1 2 0 2 0
2 68 1 2
2 69 1 2
1 3 0 2 0
2 70 1 3
2 71 1 3
1 4 0 2 0
2 72 1 4
2 73 1 4
1 5 0 2 0
2 74 1 5
2 75 1 5
1 6 0 2 0
2 76 1 6
2 77 1 6
1 7 0 2 0
2 78 1 7
2 79 1 7
1 8 0 2 0
2 80 1 8
2 81 1 8
1 9 0 2 0
2 82 1 9
2 83 1 9
1 10 0 2 0
2 84 1 10
2 85 1 10
1 11 0 2 0
2 86 1 11
2 87 1 11
1 12 0 2 0
2 88 1 12
2 89 1 12
1 13 0 2 0
2 90 1 13
2 91 1 13
1 14 0 2 0
2 92 1 14
2 93 1 14
1 15 0 2 0
2 94 1 15
2 95 1 15
1 16 0 2 0
2 96 1 16
2 165 1 16
1 17 0 2 0
2 176 1 17
2 189 1 17
1 18 0 2 0
2 206 1 18
2 221 1 18
1 19 0 2 0
2 240 1 19
2 257 1 19
1 20 0 2 0
2 276 1 20
2 295 1 20
1 21 0 2 0
2 314 1 21
2 331 1 21
1 22 0 2 0
2 348 1 22
2 368 1 22
1 23 0 2 0
2 389 1 23
2 409 1 23
1 24 0 2 0
2 433 1 24
2 453 1 24
1 25 0 2 0
2 475 1 25
2 493 1 25
1 26 0 2 0
2 520 1 26
2 544 1 26
1 27 0 2 0
2 567 1 27
2 591 1 27
1 28 0 2 0
2 614 1 28
2 638 1 28
1 29 0 2 0
2 664 1 29
2 688 1 29
1 30 0 2 0
2 709 1 30
2 733 1 30
1 31 0 2 0
2 754 1 31
2 778 1 31
1 32 0 2 0
2 800 1 32
2 808 1 32
1 33 0 2 0
2 809 1 33
2 810 1 33
1 34 0 2 0
2 811 1 34
2 812 1 34
1 35 0 2 0
2 813 1 35
2 814 1 35
1 36 0 2 0
2 815 1 36
2 816 1 36
1 37 0 2 0
2 817 1 37
2 818 1 37
1 38 0 2 0
2 819 1 38
2 820 1 38
1 39 0 2 0
2 821 1 39
2 822 1 39
1 40 0 2 0
2 823 1 40
2 824 1 40
1 41 0 2 0
2 825 1 41
2 826 1 41
1 42 0 2 0
2 827 1 42
2 828 1 42
1 43 0 2 0
2 829 1 43
2 830 1 43
1 44 0 2 0
2 831 1 44
2 832 1 44
1 45 0 2 0
2 833 1 45
2 834 1 45
1 46 0 2 0
2 835 1 46
2 836 1 46
1 47 0 2 0
2 837 1 47
2 838 1 47
1 48 0 2 0
2 839 1 48
2 840 1 48
1 49 0 2 0
2 841 1 49
2 842 1 49
1 50 0 2 0
2 843 1 50
2 844 1 50
1 51 0 2 0
2 845 1 51
2 846 1 51
1 52 0 2 0
2 847 1 52
2 848 1 52
1 53 0 2 0
2 849 1 53
2 850 1 53
1 54 0 2 0
2 851 1 54
2 852 1 54
1 55 0 2 0
2 853 1 55
2 854 1 55
1 56 0 2 0
2 855 1 56
2 856 1 56
1 57 0 2 0
2 857 1 57
2 858 1 57
1 58 0 2 0
2 859 1 58
2 860 1 58
1 59 0 2 0
2 861 1 59
2 862 1 59
1 60 0 2 0
2 863 1 60
2 864 1 60
1 61 0 2 0
2 865 1 61
2 866 1 61
1 62 0 2 0
2 867 1 62
2 868 1 62
1 63 0 2 0
2 869 1 63
2 870 1 63
2 871 1 161
2 872 1 161
2 873 1 162
2 874 1 162
2 875 1 167
2 876 1 167
2 877 1 167
2 878 1 170
2 879 1 170
2 880 1 173
2 881 1 173
2 882 1 173
2 883 1 177
2 884 1 177
2 885 1 180
2 886 1 180
2 887 1 182
2 888 1 182
2 889 1 183
2 890 1 183
2 891 1 193
2 892 1 193
2 893 1 193
2 894 1 194
2 895 1 194
2 896 1 195
2 897 1 195
2 898 1 196
2 899 1 196
2 900 1 198
2 901 1 198
2 902 1 199
2 903 1 199
2 904 1 199
2 905 1 208
2 906 1 208
2 907 1 208
2 908 1 210
2 909 1 210
2 910 1 211
2 911 1 211
2 912 1 211
2 913 1 215
2 914 1 215
2 915 1 218
2 916 1 218
2 917 1 222
2 918 1 222
2 919 1 223
2 920 1 223
2 921 1 225
2 922 1 225
2 923 1 226
2 924 1 226
2 925 1 226
2 926 1 234
2 927 1 234
2 928 1 235
2 929 1 235
2 930 1 241
2 931 1 241
2 932 1 242
2 933 1 242
2 934 1 244
2 935 1 244
2 936 1 245
2 937 1 245
2 938 1 245
2 939 1 245
2 940 1 250
2 941 1 250
2 942 1 250
2 943 1 258
2 944 1 258
2 945 1 259
2 946 1 259
2 947 1 261
2 948 1 261
2 949 1 262
2 950 1 262
2 951 1 262
2 952 1 262
2 953 1 270
2 954 1 270
2 955 1 271
2 956 1 271
2 957 1 278
2 958 1 278
2 959 1 278
2 960 1 280
2 961 1 280
2 962 1 281
2 963 1 281
2 964 1 281
2 965 1 289
2 966 1 289
2 967 1 292
2 968 1 292
2 969 1 297
2 970 1 297
2 971 1 297
2 972 1 299
2 973 1 299
2 974 1 299
2 975 1 299
2 976 1 300
2 977 1 300
2 978 1 308
2 979 1 308
2 980 1 308
2 981 1 311
2 982 1 311
2 983 1 316
2 984 1 316
2 985 1 316
2 986 1 318
2 987 1 318
2 988 1 319
2 989 1 319
2 990 1 319
2 991 1 324
2 992 1 324
2 993 1 324
2 994 1 332
2 995 1 332
2 996 1 333
2 997 1 333
2 998 1 335
2 999 1 335
2 1000 1 336
2 1001 1 336
2 1002 1 336
2 1003 1 336
2 1004 1 341
2 1005 1 341
2 1006 1 341
2 1007 1 350
2 1008 1 350
2 1009 1 350
2 1010 1 352
2 1011 1 352
2 1012 1 353
2 1013 1 353
2 1014 1 353
2 1015 1 358
2 1016 1 358
2 1017 1 359
2 1018 1 359
2 1019 1 362
2 1020 1 362
2 1021 1 363
2 1022 1 363
2 1023 1 370
2 1024 1 370
2 1025 1 370
2 1026 1 372
2 1027 1 372
2 1028 1 373
2 1029 1 373
2 1030 1 373
2 1031 1 383
2 1032 1 383
2 1033 1 386
2 1034 1 386
2 1035 1 391
2 1036 1 391
2 1037 1 391
2 1038 1 393
2 1039 1 393
2 1040 1 394
2 1041 1 394
2 1042 1 394
2 1043 1 394
2 1044 1 396
2 1045 1 396
2 1046 1 396
2 1047 1 402
2 1048 1 402
2 1049 1 403
2 1050 1 403
2 1051 1 404
2 1052 1 404
2 1053 1 404
2 1054 1 421
2 1055 1 421
2 1056 1 421
2 1057 1 424
2 1058 1 424
2 1059 1 424
2 1060 1 426
2 1061 1 426
2 1062 1 426
2 1063 1 427
2 1064 1 427
2 1065 1 427
2 1066 1 435
2 1067 1 435
2 1068 1 435
2 1069 1 437
2 1070 1 437
2 1071 1 438
2 1072 1 438
2 1073 1 438
2 1074 1 438
2 1075 1 440
2 1076 1 440
2 1077 1 446
2 1078 1 446
2 1079 1 447
2 1080 1 447
2 1081 1 449
2 1082 1 449
2 1083 1 454
2 1084 1 454
2 1085 1 455
2 1086 1 455
2 1087 1 455
2 1088 1 457
2 1089 1 457
2 1090 1 457
2 1091 1 457
2 1092 1 458
2 1093 1 458
2 1094 1 458
2 1095 1 462
2 1096 1 462
2 1097 1 468
2 1098 1 468
2 1099 1 469
2 1100 1 469
2 1101 1 470
2 1102 1 470
2 1103 1 477
2 1104 1 477
2 1105 1 477
2 1106 1 479
2 1107 1 479
2 1108 1 480
2 1109 1 480
2 1110 1 480
2 1111 1 487
2 1112 1 487
2 1113 1 489
2 1114 1 489
2 1115 1 494
2 1116 1 494
2 1117 1 495
2 1118 1 495
2 1119 1 497
2 1120 1 497
2 1121 1 498
2 1122 1 498
2 1123 1 498
2 1124 1 498
2 1125 1 502
2 1126 1 502
2 1127 1 514
2 1128 1 514
2 1129 1 515
2 1130 1 515
2 1131 1 522
2 1132 1 522
2 1133 1 522
2 1134 1 524
2 1135 1 524
2 1136 1 525
2 1137 1 525
2 1138 1 525
2 1139 1 525
2 1140 1 527
2 1141 1 527
2 1142 1 527
2 1143 1 528
2 1144 1 528
2 1145 1 535
2 1146 1 535
2 1147 1 536
2 1148 1 536
2 1149 1 538
2 1150 1 538
2 1151 1 540
2 1152 1 540
2 1153 1 546
2 1154 1 546
2 1155 1 546
2 1156 1 548
2 1157 1 548
2 1158 1 549
2 1159 1 549
2 1160 1 549
2 1161 1 549
2 1162 1 561
2 1163 1 561
2 1164 1 562
2 1165 1 562
2 1166 1 569
2 1167 1 569
2 1168 1 569
2 1169 1 569
2 1170 1 571
2 1171 1 571
2 1172 1 571
2 1173 1 572
2 1174 1 572
2 1175 1 572
2 1176 1 572
2 1177 1 574
2 1178 1 574
2 1179 1 574
2 1180 1 575
2 1181 1 575
2 1182 1 582
2 1183 1 582
2 1184 1 583
2 1185 1 583
2 1186 1 585
2 1187 1 585
2 1188 1 586
2 1189 1 586
2 1190 1 592
2 1191 1 592
2 1192 1 593
2 1193 1 593
2 1194 1 595
2 1195 1 595
2 1196 1 596
2 1197 1 596
2 1198 1 596
2 1199 1 596
2 1200 1 608
2 1201 1 608
2 1202 1 609
2 1203 1 609
2 1204 1 616
2 1205 1 616
2 1206 1 616
2 1207 1 619
2 1208 1 619
2 1209 1 619
2 1210 1 619
2 1211 1 619
2 1212 1 619
2 1213 1 621
2 1214 1 621
2 1215 1 621
2 1216 1 622
2 1217 1 622
2 1218 1 629
2 1219 1 629
2 1220 1 632
2 1221 1 632
2 1222 1 633
2 1223 1 633
2 1224 1 640
2 1225 1 640
2 1226 1 640
2 1227 1 642
2 1228 1 642
2 1229 1 642
2 1230 1 643
2 1231 1 643
2 1232 1 643
2 1233 1 648
2 1234 1 648
2 1235 1 655
2 1236 1 655
2 1237 1 658
2 1238 1 658
2 1239 1 661
2 1240 1 661
2 1241 1 665
2 1242 1 665
2 1243 1 665
2 1244 1 671
2 1245 1 671
2 1246 1 673
2 1247 1 673
2 1248 1 676
2 1249 1 676
2 1250 1 677
2 1251 1 677
2 1252 1 679
2 1253 1 679
2 1254 1 679
2 1255 1 681
2 1256 1 681
2 1257 1 682
2 1258 1 682
2 1259 1 682
2 1260 1 690
2 1261 1 690
2 1262 1 690
2 1263 1 692
2 1264 1 692
2 1265 1 693
2 1266 1 693
2 1267 1 693
2 1268 1 703
2 1269 1 703
2 1270 1 706
2 1271 1 706
2 1272 1 711
2 1273 1 711
2 1274 1 711
2 1275 1 713
2 1276 1 713
2 1277 1 714
2 1278 1 714
2 1279 1 714
2 1280 1 716
2 1281 1 716
2 1282 1 716
2 1283 1 716
2 1284 1 725
2 1285 1 725
2 1286 1 725
2 1287 1 727
2 1288 1 727
2 1289 1 728
2 1290 1 728
2 1291 1 735
2 1292 1 735
2 1293 1 737
2 1294 1 737
2 1295 1 738
2 1296 1 738
2 1297 1 738
2 1298 1 748
2 1299 1 748
2 1300 1 759
2 1301 1 759
2 1302 1 765
2 1303 1 765
2 1304 1 766
2 1305 1 766
2 1306 1 769
2 1307 1 769
2 1308 1 771
2 1309 1 771
2 1310 1 772
2 1311 1 772
2 1312 1 772
2 1313 1 781
2 1314 1 781
2 1315 1 787
2 1316 1 787
2 1317 1 788
2 1318 1 788
2 1319 1 791
2 1320 1 791
2 1321 1 793
2 1322 1 793
2 1323 1 794
2 1324 1 794
0 97 5 1 1 64
0 98 5 1 1 66
0 99 5 1 1 68
0 100 5 1 1 70
0 101 5 1 1 72
0 102 5 1 1 74
0 103 5 1 1 76
0 104 5 1 1 78
0 105 5 1 1 80
0 106 5 1 1 82
0 107 5 1 1 84
0 108 5 1 1 86
0 109 5 1 1 88
0 110 5 1 1 90
0 111 5 1 1 92
0 112 5 1 1 94
0 113 5 1 1 96
0 114 5 1 1 176
0 115 5 1 1 206
0 116 5 1 1 240
0 117 5 1 1 276
0 118 5 1 1 314
0 119 5 1 1 348
0 120 5 1 1 389
0 121 5 1 1 433
0 122 5 1 1 475
0 123 5 1 1 520
0 124 5 1 1 567
0 125 5 1 1 614
0 126 5 1 1 664
0 127 5 1 1 709
0 128 5 1 1 754
0 129 5 1 1 800
0 130 5 1 1 809
0 131 5 1 1 811
0 132 5 1 1 813
0 133 5 1 1 815
0 134 5 1 1 817
0 135 5 1 1 819
0 136 5 1 1 821
0 137 5 1 1 823
0 138 5 1 1 825
0 139 5 1 1 827
0 140 5 1 1 829
0 141 5 1 1 831
0 142 5 1 1 833
0 143 5 1 1 835
0 144 5 1 1 837
0 145 5 1 1 839
0 146 5 1 1 841
0 147 5 1 1 843
0 148 5 1 1 845
0 149 5 1 1 847
0 150 5 1 1 849
0 151 5 1 1 851
0 152 5 1 1 853
0 153 5 1 1 855
0 154 5 1 1 857
0 155 5 1 1 859
0 156 5 1 1 861
0 157 5 1 1 863
0 158 5 1 1 865
0 159 5 1 1 867
0 160 5 1 1 869
0 161 7 2 2 65 808
0 162 5 2 1 871
0 163 7 1 2 97 129
0 164 5 1 1 163
3 1667 7 0 2 873 164
0 166 7 1 2 67 810
0 167 5 3 1 166
0 168 7 1 2 98 130
0 169 5 1 1 168
0 170 7 2 2 875 169
0 171 5 1 1 878
0 172 7 1 2 872 879
0 173 5 3 1 172
0 174 7 1 2 874 171
0 175 5 1 1 174
3 1668 7 0 2 880 175
0 177 7 2 2 876 881
0 178 5 1 1 883
0 179 7 1 2 99 131
0 180 5 2 1 179
0 181 7 1 2 69 812
0 182 5 2 1 181
0 183 7 2 2 885 887
0 184 5 1 1 889
0 185 7 1 2 178 890
0 186 5 1 1 185
0 187 7 1 2 884 184
0 188 5 1 1 187
3 1669 7 0 2 186 188
0 190 7 1 2 877 888
0 191 7 1 2 882 190
0 192 5 1 1 191
0 193 7 3 2 886 192
0 194 5 2 1 891
0 195 7 2 2 71 814
0 196 5 2 1 896
0 197 7 1 2 100 132
0 198 5 2 1 197
0 199 7 3 2 898 900
0 200 5 1 1 902
0 201 7 1 2 892 200
0 202 5 1 1 201
0 203 7 1 2 894 903
0 204 5 1 1 203
0 205 7 1 2 202 204
3 1670 5 0 1 205
0 207 7 1 2 73 816
0 208 5 3 1 207
0 209 7 1 2 101 133
0 210 5 2 1 209
0 211 7 3 2 905 908
0 212 5 1 1 910
0 213 7 1 2 895 899
0 214 5 1 1 213
0 215 7 2 2 901 214
0 216 5 1 1 913
0 217 7 1 2 911 914
0 218 5 2 1 217
0 219 7 1 2 212 216
0 220 5 1 1 219
3 1671 7 0 2 915 220
0 222 7 2 2 75 818
0 223 5 2 1 917
0 224 7 1 2 102 134
0 225 5 2 1 224
0 226 7 3 2 919 921
0 227 5 1 1 923
0 228 7 1 2 904 912
0 229 7 1 2 893 228
0 230 5 1 1 229
0 231 7 1 2 897 909
0 232 5 1 1 231
0 233 7 1 2 906 232
0 234 7 2 2 230 233
0 235 5 2 1 926
0 236 7 1 2 924 928
0 237 5 1 1 236
0 238 7 1 2 227 927
0 239 5 1 1 238
3 1672 7 0 2 237 239
0 241 7 2 2 77 820
0 242 5 2 1 930
0 243 7 1 2 103 135
0 244 5 2 1 243
0 245 7 4 2 932 934
0 246 5 1 1 936
0 247 7 1 2 907 920
0 248 7 1 2 916 247
0 249 5 1 1 248
0 250 7 3 2 922 249
0 251 5 1 1 940
0 252 7 1 2 937 251
0 253 5 1 1 252
0 254 7 1 2 246 941
0 255 5 1 1 254
0 256 7 1 2 253 255
3 1673 5 0 1 256
0 258 7 2 2 79 822
0 259 5 2 1 943
0 260 7 1 2 104 136
0 261 5 2 1 260
0 262 7 4 2 945 947
0 263 5 1 1 949
0 264 7 1 2 925 938
0 265 7 1 2 929 264
0 266 5 1 1 265
0 267 7 1 2 918 935
0 268 5 1 1 267
0 269 7 1 2 933 268
0 270 7 2 2 266 269
0 271 5 2 1 953
0 272 7 1 2 950 955
0 273 5 1 1 272
0 274 7 1 2 263 954
0 275 5 1 1 274
3 1674 7 0 2 273 275
0 277 7 1 2 81 824
0 278 5 3 1 277
0 279 7 1 2 105 137
0 280 5 2 1 279
0 281 7 3 2 957 960
0 282 5 1 1 962
0 283 7 1 2 939 951
0 284 7 1 2 942 283
0 285 5 1 1 284
0 286 7 1 2 931 948
0 287 5 1 1 286
0 288 7 1 2 946 287
0 289 7 2 2 285 288
0 290 5 1 1 965
0 291 7 1 2 963 290
0 292 5 2 1 291
0 293 7 1 2 282 966
0 294 5 1 1 293
3 1675 7 0 2 967 294
0 296 7 1 2 106 138
0 297 5 3 1 296
0 298 7 1 2 83 826
0 299 5 4 1 298
0 300 7 2 2 969 972
0 301 5 1 1 976
0 302 7 1 2 952 964
0 303 7 1 2 956 302
0 304 5 1 1 303
0 305 7 1 2 944 961
0 306 5 1 1 305
0 307 7 1 2 958 306
0 308 7 3 2 304 307
0 309 5 1 1 978
0 310 7 1 2 977 309
0 311 5 2 1 310
0 312 7 1 2 301 979
0 313 5 1 1 312
3 1676 7 0 2 981 313
0 315 7 1 2 85 828
0 316 5 3 1 315
0 317 7 1 2 107 139
0 318 5 2 1 317
0 319 7 3 2 983 986
0 320 5 1 1 988
0 321 7 1 2 959 973
0 322 7 1 2 968 321
0 323 5 1 1 322
0 324 7 3 2 970 323
0 325 5 1 1 991
0 326 7 1 2 989 325
0 327 5 1 1 326
0 328 7 1 2 320 992
0 329 5 1 1 328
0 330 7 1 2 327 329
3 1677 5 0 1 330
0 332 7 2 2 87 830
0 333 5 2 1 994
0 334 7 1 2 108 140
0 335 5 2 1 334
0 336 7 4 2 996 998
0 337 5 1 1 1000
0 338 7 1 2 974 984
0 339 7 1 2 982 338
0 340 5 1 1 339
0 341 7 3 2 987 340
0 342 5 1 1 1004
0 343 7 1 2 1001 342
0 344 5 1 1 343
0 345 7 1 2 337 1005
0 346 5 1 1 345
0 347 7 1 2 344 346
3 1678 5 0 1 347
0 349 7 1 2 89 832
0 350 5 3 1 349
0 351 7 1 2 109 141
0 352 5 2 1 351
0 353 7 3 2 1007 1010
0 354 5 1 1 1012
0 355 7 1 2 985 997
0 356 5 1 1 355
0 357 7 1 2 999 356
0 358 5 2 1 357
0 359 7 2 2 990 1002
0 360 7 1 2 993 1017
0 361 5 1 1 360
0 362 7 2 2 1015 361
0 363 5 2 1 1019
0 364 7 1 2 1013 1021
0 365 5 1 1 364
0 366 7 1 2 354 1020
0 367 5 1 1 366
3 1679 7 0 2 365 367
0 369 7 1 2 91 834
0 370 5 3 1 369
0 371 7 1 2 110 142
0 372 5 2 1 371
0 373 7 3 2 1023 1026
0 374 5 1 1 1028
0 375 7 1 2 975 980
0 376 5 1 1 375
0 377 7 1 2 971 1018
0 378 7 1 2 376 377
0 379 5 1 1 378
0 380 7 1 2 1008 1016
0 381 7 1 2 379 380
0 382 5 1 1 381
0 383 7 2 2 1011 382
0 384 5 1 1 1031
0 385 7 1 2 1029 1032
0 386 5 2 1 385
0 387 7 1 2 374 384
0 388 5 1 1 387
3 1680 7 0 2 1033 388
0 390 7 1 2 93 836
0 391 5 3 1 390
0 392 7 1 2 111 143
0 393 5 2 1 392
0 394 7 4 2 1035 1038
0 395 5 1 1 1040
0 396 7 3 2 1014 1030
0 397 7 1 2 1022 1044
0 398 5 1 1 397
0 399 7 1 2 1009 1024
0 400 5 1 1 399
0 401 7 1 2 1027 400
0 402 5 2 1 401
0 403 7 2 2 398 1047
0 404 5 3 1 1049
0 405 7 1 2 1041 1051
0 406 5 1 1 405
0 407 7 1 2 395 1050
0 408 5 1 1 407
3 1681 7 0 2 406 408
0 410 7 1 2 1003 1042
0 411 7 1 2 1045 410
0 412 7 1 2 1006 411
0 413 5 1 1 412
0 414 7 1 2 995 1046
0 415 5 1 1 414
0 416 7 1 2 1036 1048
0 417 7 1 2 415 416
0 418 5 1 1 417
0 419 7 1 2 1039 418
0 420 5 1 1 419
0 421 7 3 2 413 420
0 422 5 1 1 1054
0 423 7 1 2 95 838
0 424 5 3 1 423
0 425 7 1 2 112 144
0 426 5 3 1 425
0 427 7 3 2 1057 1060
0 428 5 1 1 1063
0 429 7 1 2 422 1064
0 430 5 1 1 429
0 431 7 1 2 1055 428
0 432 5 1 1 431
3 1682 7 0 2 430 432
0 434 7 1 2 165 840
0 435 5 3 1 434
0 436 7 1 2 113 145
0 437 5 2 1 436
0 438 7 4 2 1066 1069
0 439 5 1 1 1071
0 440 7 2 2 1043 1065
0 441 7 1 2 1052 1075
0 442 5 1 1 441
0 443 7 1 2 1037 1058
0 444 5 1 1 443
0 445 7 1 2 1061 444
0 446 5 2 1 445
0 447 7 2 2 442 1077
0 448 5 1 1 1079
0 449 7 2 2 1072 448
0 450 5 1 1 1081
0 451 7 1 2 439 1080
0 452 5 1 1 451
3 1683 7 0 2 450 452
0 454 7 2 2 189 842
0 455 5 3 1 1083
0 456 7 1 2 114 146
0 457 5 4 1 456
0 458 7 3 2 1085 1088
0 459 5 1 1 1092
0 460 7 1 2 1025 1034
0 461 5 1 1 460
0 462 7 2 2 1073 1076
0 463 7 1 2 461 1095
0 464 5 1 1 463
0 465 7 1 2 1067 1078
0 466 5 1 1 465
0 467 7 1 2 1070 466
0 468 5 2 1 467
0 469 7 2 2 464 1097
0 470 5 2 1 1099
0 471 7 1 2 1093 1101
0 472 5 1 1 471
0 473 7 1 2 459 1100
0 474 5 1 1 473
3 1684 7 0 2 472 474
0 476 7 1 2 221 844
0 477 5 3 1 476
0 478 7 1 2 115 147
0 479 5 2 1 478
0 480 7 3 2 1103 1106
0 481 5 1 1 1108
0 482 7 1 2 1053 1096
0 483 5 1 1 482
0 484 7 1 2 1086 1098
0 485 7 1 2 483 484
0 486 5 1 1 485
0 487 7 2 2 1089 486
0 488 5 1 1 1111
0 489 7 2 2 1109 1112
0 490 5 1 1 1113
0 491 7 1 2 481 488
0 492 5 1 1 491
3 1685 7 0 2 490 492
0 494 7 2 2 257 846
0 495 5 2 1 1115
0 496 7 1 2 116 148
0 497 5 2 1 496
0 498 7 4 2 1117 1119
0 499 5 1 1 1121
0 500 7 1 2 1068 1087
0 501 5 1 1 500
0 502 7 2 2 1090 501
0 503 5 1 1 1125
0 504 7 1 2 1056 1059
0 505 5 1 1 504
0 506 7 1 2 1062 1091
0 507 7 1 2 1074 506
0 508 7 1 2 505 507
0 509 5 1 1 508
0 510 7 1 2 503 509
0 511 5 1 1 510
0 512 7 1 2 1107 511
0 513 5 1 1 512
0 514 7 2 2 1104 513
0 515 5 2 1 1127
0 516 7 1 2 1122 1129
0 517 5 1 1 516
0 518 7 1 2 499 1128
0 519 5 1 1 518
3 1686 7 0 2 517 519
0 521 7 1 2 295 848
0 522 5 3 1 521
0 523 7 1 2 117 149
0 524 5 2 1 523
0 525 7 4 2 1131 1134
0 526 5 1 1 1136
0 527 7 3 2 1110 1123
0 528 7 2 2 1094 1140
0 529 7 1 2 1082 1143
0 530 5 1 1 529
0 531 7 1 2 1126 1141
0 532 5 1 1 531
0 533 7 1 2 1105 1118
0 534 5 1 1 533
0 535 7 2 2 1120 534
0 536 5 2 1 1145
0 537 7 1 2 532 1147
0 538 7 2 2 530 537
0 539 5 1 1 1149
0 540 7 2 2 1137 539
0 541 5 1 1 1151
0 542 7 1 2 526 1150
0 543 5 1 1 542
3 1687 7 0 2 541 543
0 545 7 1 2 331 850
0 546 5 3 1 545
0 547 7 1 2 118 150
0 548 5 2 1 547
0 549 7 4 2 1153 1156
0 550 5 1 1 1158
0 551 7 1 2 1084 1142
0 552 5 1 1 551
0 553 7 1 2 1132 1148
0 554 7 1 2 552 553
0 555 5 1 1 554
0 556 7 1 2 1135 555
0 557 5 1 1 556
0 558 7 1 2 1138 1144
0 559 7 1 2 1102 558
0 560 5 1 1 559
0 561 7 2 2 557 560
0 562 5 2 1 1162
0 563 7 1 2 1159 1164
0 564 5 1 1 563
0 565 7 1 2 550 1163
0 566 5 1 1 565
3 1688 7 0 2 564 566
0 568 7 1 2 368 852
0 569 5 4 1 568
0 570 7 1 2 119 151
0 571 5 3 1 570
0 572 7 4 2 1166 1170
0 573 5 1 1 1173
0 574 7 3 2 1139 1160
0 575 7 2 2 1124 1177
0 576 7 1 2 1114 1180
0 577 5 1 1 576
0 578 7 1 2 1146 1178
0 579 5 1 1 578
0 580 7 1 2 1133 1154
0 581 5 1 1 580
0 582 7 2 2 1157 581
0 583 5 2 1 1182
0 584 7 1 2 579 1184
0 585 7 2 2 577 584
0 586 5 2 1 1186
0 587 7 1 2 1174 1188
0 588 5 1 1 587
0 589 7 1 2 573 1187
0 590 5 1 1 589
3 1689 7 0 2 588 590
0 592 7 2 2 409 854
0 593 5 2 1 1190
0 594 7 1 2 120 152
0 595 5 2 1 594
0 596 7 4 2 1192 1194
0 597 5 1 1 1196
0 598 7 1 2 1175 1181
0 599 7 1 2 1130 598
0 600 5 1 1 599
0 601 7 1 2 1116 1179
0 602 5 1 1 601
0 603 7 1 2 1167 1185
0 604 7 1 2 602 603
0 605 5 1 1 604
0 606 7 1 2 1171 605
0 607 5 1 1 606
0 608 7 2 2 600 607
0 609 5 2 1 1200
0 610 7 1 2 1197 1202
0 611 5 1 1 610
0 612 7 1 2 597 1201
0 613 5 1 1 612
3 1690 7 0 2 611 613
0 615 7 1 2 453 856
0 616 5 3 1 615
0 617 7 1 2 121 153
0 618 5 1 1 617
0 619 7 6 2 1204 618
0 620 5 1 1 1207
0 621 7 3 2 1176 1198
0 622 7 2 2 1161 1213
0 623 7 1 2 1152 1216
0 624 5 1 1 623
0 625 7 1 2 1183 1214
0 626 5 1 1 625
0 627 7 1 2 1168 1193
0 628 5 1 1 627
0 629 7 2 2 1195 628
0 630 5 1 1 1218
0 631 7 1 2 626 630
0 632 7 2 2 624 631
0 633 5 2 1 1220
0 634 7 1 2 1208 1222
0 635 5 1 1 634
0 636 7 1 2 620 1221
0 637 5 1 1 636
3 1691 7 0 2 635 637
0 639 7 1 2 493 858
0 640 5 3 1 639
0 641 7 1 2 122 154
0 642 5 3 1 641
0 643 7 3 2 1224 1227
0 644 5 1 1 1230
0 645 7 1 2 1209 1217
0 646 7 1 2 1165 645
0 647 5 1 1 646
0 648 7 2 2 1199 1210
0 649 7 1 2 1155 1169
0 650 5 1 1 649
0 651 7 1 2 1172 650
0 652 7 1 2 1233 651
0 653 5 1 1 652
0 654 7 1 2 1191 1211
0 655 5 2 1 654
0 656 7 1 2 1205 1235
0 657 7 1 2 653 656
0 658 7 2 2 647 657
0 659 5 1 1 1237
0 660 7 1 2 1231 659
0 661 5 2 1 660
0 662 7 1 2 644 1238
0 663 5 1 1 662
3 1692 7 0 2 1239 663
0 665 7 3 2 1212 1232
0 666 7 1 2 1215 1241
0 667 7 1 2 1189 666
0 668 5 1 1 667
0 669 7 1 2 1219 1242
0 670 5 1 1 669
0 671 7 2 2 1206 1225
0 672 5 1 1 1244
0 673 7 2 2 1228 672
0 674 5 1 1 1246
0 675 7 1 2 670 674
0 676 7 2 2 668 675
0 677 5 2 1 1248
0 678 7 1 2 544 860
0 679 5 3 1 678
0 680 7 1 2 123 155
0 681 5 2 1 680
0 682 7 3 2 1252 1255
0 683 5 1 1 1257
0 684 7 1 2 1250 1258
0 685 5 1 1 684
0 686 7 1 2 1249 683
0 687 5 1 1 686
3 1693 7 0 2 685 687
0 689 7 1 2 591 862
0 690 5 3 1 689
0 691 7 1 2 124 156
0 692 5 2 1 691
0 693 7 3 2 1260 1263
0 694 5 1 1 1265
0 695 7 1 2 1203 1234
0 696 5 1 1 695
0 697 7 1 2 1236 1245
0 698 7 1 2 696 697
0 699 5 1 1 698
0 700 7 1 2 1229 1256
0 701 7 1 2 699 700
0 702 5 1 1 701
0 703 7 2 2 1253 702
0 704 5 1 1 1268
0 705 7 1 2 1266 704
0 706 5 2 1 705
0 707 7 1 2 694 1269
0 708 5 1 1 707
3 1694 7 0 2 1270 708
0 710 7 1 2 638 864
0 711 5 3 1 710
0 712 7 1 2 125 157
0 713 5 2 1 712
0 714 7 3 2 1272 1275
0 715 5 1 1 1277
0 716 7 4 2 1259 1267
0 717 7 1 2 1243 1280
0 718 7 1 2 1223 717
0 719 5 1 1 718
0 720 7 1 2 1247 1281
0 721 5 1 1 720
0 722 7 1 2 1254 1261
0 723 5 1 1 722
0 724 7 1 2 1264 723
0 725 5 3 1 724
0 726 7 1 2 721 1284
0 727 7 2 2 719 726
0 728 5 2 1 1287
0 729 7 1 2 1278 1289
0 730 5 1 1 729
0 731 7 1 2 715 1288
0 732 5 1 1 731
3 1695 7 0 2 730 732
0 734 7 1 2 688 866
0 735 5 2 1 734
0 736 7 1 2 126 158
0 737 5 2 1 736
0 738 7 3 2 1291 1293
0 739 5 1 1 1295
0 740 7 1 2 1226 1240
0 741 5 1 1 740
0 742 7 1 2 1282 741
0 743 5 1 1 742
0 744 7 1 2 1285 743
0 745 5 1 1 744
0 746 7 1 2 1276 745
0 747 5 1 1 746
0 748 7 2 2 1273 747
0 749 5 1 1 1298
0 750 7 1 2 1296 749
0 751 5 1 1 750
0 752 7 1 2 739 1299
0 753 5 1 1 752
3 1696 7 0 2 751 753
0 755 7 1 2 1251 1283
0 756 5 1 1 755
0 757 7 1 2 1286 756
0 758 5 1 1 757
0 759 7 2 2 1279 1297
0 760 7 1 2 758 1300
0 761 5 1 1 760
0 762 7 1 2 1274 1292
0 763 5 1 1 762
0 764 7 1 2 1294 763
0 765 5 2 1 764
0 766 7 2 2 761 1302
0 767 5 1 1 1304
0 768 7 1 2 733 868
0 769 5 2 1 768
0 770 7 1 2 127 159
0 771 5 2 1 770
0 772 7 3 2 1306 1308
0 773 5 1 1 1310
0 774 7 1 2 767 1311
0 775 5 1 1 774
0 776 7 1 2 1305 773
0 777 5 1 1 776
3 1697 7 0 2 775 777
0 779 7 1 2 1262 1271
0 780 5 1 1 779
0 781 7 2 2 1301 1312
0 782 7 1 2 780 1313
0 783 5 1 1 782
0 784 7 1 2 1303 1307
0 785 5 1 1 784
0 786 7 1 2 1309 785
0 787 5 2 1 786
0 788 7 2 2 783 1315
0 789 5 1 1 1317
0 790 7 1 2 778 870
0 791 5 2 1 790
0 792 7 1 2 128 160
0 793 5 2 1 792
0 794 7 2 2 1319 1321
0 795 5 1 1 1323
0 796 7 1 2 789 1324
0 797 5 1 1 796
0 798 7 1 2 1318 795
0 799 5 1 1 798
3 1698 7 0 2 797 799
0 801 7 1 2 1290 1314
0 802 5 1 1 801
0 803 7 1 2 1316 802
0 804 5 1 1 803
0 805 7 1 2 1322 804
0 806 5 1 1 805
0 807 7 1 2 1320 806
3 1699 5 0 1 807
