1 0 0 8 0
2 32 1 0
2 1258 1 0
2 1259 1 0
2 1260 1 0
2 1261 1 0
2 1262 1 0
2 1263 1 0
2 1264 1 0
1 1 0 8 0
2 1265 1 1
2 1266 1 1
2 1267 1 1
2 1268 1 1
2 1269 1 1
2 1270 1 1
2 1271 1 1
2 1272 1 1
1 2 0 8 0
2 1273 1 2
2 1274 1 2
2 1275 1 2
2 1276 1 2
2 1277 1 2
2 1278 1 2
2 1279 1 2
2 1280 1 2
1 3 0 9 0
2 1281 1 3
2 1282 1 3
2 1283 1 3
2 1284 1 3
2 1285 1 3
2 1286 1 3
2 1287 1 3
2 1288 1 3
2 1289 1 3
1 4 0 8 0
2 1290 1 4
2 1291 1 4
2 1292 1 4
2 1293 1 4
2 1294 1 4
2 1295 1 4
2 1296 1 4
2 1297 1 4
1 5 0 9 0
2 1298 1 5
2 1299 1 5
2 1300 1 5
2 1301 1 5
2 1302 1 5
2 1303 1 5
2 1304 1 5
2 1305 1 5
2 1306 1 5
1 6 0 8 0
2 1307 1 6
2 1308 1 6
2 1309 1 6
2 1310 1 6
2 1311 1 6
2 1312 1 6
2 1313 1 6
2 1314 1 6
1 7 0 8 0
2 1315 1 7
2 1316 1 7
2 1317 1 7
2 1318 1 7
2 1319 1 7
2 1320 1 7
2 1321 1 7
2 1322 1 7
1 8 0 8 0
2 1323 1 8
2 1324 1 8
2 1325 1 8
2 1326 1 8
2 1327 1 8
2 1328 1 8
2 1329 1 8
2 1330 1 8
1 9 0 8 0
2 1331 1 9
2 1332 1 9
2 1333 1 9
2 1334 1 9
2 1335 1 9
2 1336 1 9
2 1337 1 9
2 1338 1 9
1 10 0 9 0
2 1339 1 10
2 1340 1 10
2 1341 1 10
2 1342 1 10
2 1343 1 10
2 1344 1 10
2 1345 1 10
2 1346 1 10
2 1347 1 10
1 11 0 8 0
2 1348 1 11
2 1349 1 11
2 1350 1 11
2 1351 1 11
2 1352 1 11
2 1353 1 11
2 1354 1 11
2 1355 1 11
1 12 0 8 0
2 1356 1 12
2 1357 1 12
2 1358 1 12
2 1359 1 12
2 1360 1 12
2 1361 1 12
2 1362 1 12
2 1363 1 12
1 13 0 8 0
2 1364 1 13
2 1365 1 13
2 1366 1 13
2 1367 1 13
2 1368 1 13
2 1369 1 13
2 1370 1 13
2 1371 1 13
1 14 0 8 0
2 1372 1 14
2 1373 1 14
2 1374 1 14
2 1375 1 14
2 1376 1 14
2 1377 1 14
2 1378 1 14
2 1379 1 14
1 15 0 8 0
2 1380 1 15
2 1381 1 15
2 1382 1 15
2 1383 1 15
2 1384 1 15
2 1385 1 15
2 1386 1 15
2 1387 1 15
1 16 0 2 0
2 1388 1 16
2 1389 1 16
1 17 0 2 0
2 1390 1 17
2 1391 1 17
1 18 0 2 0
2 1392 1 18
2 1393 1 18
1 19 0 2 0
2 1394 1 19
2 1395 1 19
1 20 0 2 0
2 1396 1 20
2 1397 1 20
1 21 0 2 0
2 1398 1 21
2 1399 1 21
1 22 0 2 0
2 1400 1 22
2 1401 1 22
1 23 0 2 0
2 1402 1 23
2 1403 1 23
1 24 0 2 0
2 1404 1 24
2 1405 1 24
1 25 0 2 0
2 1406 1 25
2 1407 1 25
1 26 0 2 0
2 1408 1 26
2 1409 1 26
1 27 0 2 0
2 1410 1 27
2 1411 1 27
1 28 0 2 0
2 1412 1 28
2 1413 1 28
1 29 0 2 0
2 1414 1 29
2 1415 1 29
1 30 0 2 0
2 1416 1 30
2 1417 1 30
1 31 0 2 0
2 1418 1 31
2 1419 1 31
2 1420 1 49
2 1421 1 49
2 1422 1 51
2 1423 1 51
2 1424 1 53
2 1425 1 53
2 1426 1 55
2 1427 1 55
2 1428 1 58
2 1429 1 58
2 1430 1 61
2 1431 1 61
2 1432 1 64
2 1433 1 64
2 1434 1 67
2 1435 1 67
2 1436 1 70
2 1437 1 70
2 1438 1 71
2 1439 1 71
2 1440 1 75
2 1441 1 75
2 1442 1 78
2 1443 1 78
2 1444 1 79
2 1445 1 79
2 1446 1 81
2 1447 1 81
2 1448 1 83
2 1449 1 83
2 1450 1 85
2 1451 1 85
2 1452 1 87
2 1453 1 87
2 1454 1 89
2 1455 1 89
2 1456 1 92
2 1457 1 92
2 1458 1 95
2 1459 1 95
2 1460 1 98
2 1461 1 98
2 1462 1 101
2 1463 1 101
2 1464 1 104
2 1465 1 104
2 1466 1 107
2 1467 1 107
2 1468 1 110
2 1469 1 110
2 1470 1 113
2 1471 1 113
2 1472 1 116
2 1473 1 116
2 1474 1 117
2 1475 1 117
2 1476 1 119
2 1477 1 119
2 1478 1 121
2 1479 1 121
2 1480 1 123
2 1481 1 123
2 1482 1 124
2 1483 1 124
2 1484 1 125
2 1485 1 125
2 1486 1 126
2 1487 1 126
2 1488 1 128
2 1489 1 128
2 1490 1 129
2 1491 1 129
2 1492 1 133
2 1493 1 133
2 1494 1 136
2 1495 1 136
2 1496 1 137
2 1497 1 137
2 1498 1 141
2 1499 1 141
2 1500 1 144
2 1501 1 144
2 1502 1 145
2 1503 1 145
2 1504 1 149
2 1505 1 149
2 1506 1 152
2 1507 1 152
2 1508 1 153
2 1509 1 153
2 1510 1 157
2 1511 1 157
2 1512 1 160
2 1513 1 160
2 1514 1 161
2 1515 1 161
2 1516 1 165
2 1517 1 165
2 1518 1 168
2 1519 1 168
2 1520 1 169
2 1521 1 169
2 1522 1 173
2 1523 1 173
2 1524 1 176
2 1525 1 176
2 1526 1 177
2 1527 1 177
2 1528 1 179
2 1529 1 179
2 1530 1 181
2 1531 1 181
2 1532 1 183
2 1533 1 183
2 1534 1 184
2 1535 1 184
2 1536 1 185
2 1537 1 185
2 1538 1 187
2 1539 1 187
2 1540 1 190
2 1541 1 190
2 1542 1 193
2 1543 1 193
2 1544 1 196
2 1545 1 196
2 1546 1 199
2 1547 1 199
2 1548 1 202
2 1549 1 202
2 1550 1 205
2 1551 1 205
2 1552 1 208
2 1553 1 208
2 1554 1 211
2 1555 1 211
2 1556 1 214
2 1557 1 214
2 1558 1 215
2 1559 1 215
2 1560 1 217
2 1561 1 217
2 1562 1 220
2 1563 1 220
2 1564 1 223
2 1565 1 223
2 1566 1 227
2 1567 1 227
2 1568 1 230
2 1569 1 230
2 1570 1 231
2 1571 1 231
2 1572 1 235
2 1573 1 235
2 1574 1 238
2 1575 1 238
2 1576 1 239
2 1577 1 239
2 1578 1 241
2 1579 1 241
2 1580 1 244
2 1581 1 244
2 1582 1 245
2 1583 1 245
2 1584 1 247
2 1585 1 247
2 1586 1 253
2 1587 1 253
2 1588 1 256
2 1589 1 256
2 1590 1 259
2 1591 1 259
2 1592 1 262
2 1593 1 262
2 1594 1 265
2 1595 1 265
2 1596 1 269
2 1597 1 269
2 1598 1 272
2 1599 1 272
2 1600 1 273
2 1601 1 273
2 1602 1 277
2 1603 1 277
2 1604 1 280
2 1605 1 280
2 1606 1 281
2 1607 1 281
2 1608 1 283
2 1609 1 283
2 1610 1 286
2 1611 1 286
2 1612 1 289
2 1613 1 289
2 1614 1 293
2 1615 1 293
2 1616 1 296
2 1617 1 296
2 1618 1 297
2 1619 1 297
2 1620 1 301
2 1621 1 301
2 1622 1 304
2 1623 1 304
2 1624 1 305
2 1625 1 305
2 1626 1 309
2 1627 1 309
2 1628 1 312
2 1629 1 312
2 1630 1 313
2 1631 1 313
2 1632 1 317
2 1633 1 317
2 1634 1 320
2 1635 1 320
2 1636 1 321
2 1637 1 321
2 1638 1 325
2 1639 1 325
2 1640 1 328
2 1641 1 328
2 1642 1 329
2 1643 1 329
2 1644 1 331
2 1645 1 331
2 1646 1 334
2 1647 1 334
2 1648 1 335
2 1649 1 335
2 1650 1 339
2 1651 1 339
2 1652 1 342
2 1653 1 342
2 1654 1 343
2 1655 1 343
2 1656 1 345
2 1657 1 345
2 1658 1 347
2 1659 1 347
2 1660 1 350
2 1661 1 350
2 1662 1 351
2 1663 1 351
2 1664 1 353
2 1665 1 353
2 1666 1 355
2 1667 1 355
2 1668 1 357
2 1669 1 357
2 1670 1 358
2 1671 1 358
2 1672 1 359
2 1673 1 359
2 1674 1 360
2 1675 1 360
2 1676 1 361
2 1677 1 361
2 1678 1 362
2 1679 1 362
2 1680 1 363
2 1681 1 363
2 1682 1 364
2 1683 1 364
2 1684 1 365
2 1685 1 365
2 1686 1 368
2 1687 1 368
2 1688 1 371
2 1689 1 371
2 1690 1 375
2 1691 1 375
2 1692 1 378
2 1693 1 378
2 1694 1 381
2 1695 1 381
2 1696 1 385
2 1697 1 385
2 1698 1 388
2 1699 1 388
2 1700 1 389
2 1701 1 389
2 1702 1 392
2 1703 1 392
2 1704 1 393
2 1705 1 393
2 1706 1 397
2 1707 1 397
2 1708 1 400
2 1709 1 400
2 1710 1 401
2 1711 1 401
2 1712 1 405
2 1713 1 405
2 1714 1 408
2 1715 1 408
2 1716 1 409
2 1717 1 409
2 1718 1 413
2 1719 1 413
2 1720 1 416
2 1721 1 416
2 1722 1 419
2 1723 1 419
2 1724 1 423
2 1725 1 423
2 1726 1 426
2 1727 1 426
2 1728 1 429
2 1729 1 429
2 1730 1 433
2 1731 1 433
2 1732 1 436
2 1733 1 436
2 1734 1 437
2 1735 1 437
2 1736 1 439
2 1737 1 439
2 1738 1 442
2 1739 1 442
2 1740 1 443
2 1741 1 443
2 1742 1 447
2 1743 1 447
2 1744 1 450
2 1745 1 450
2 1746 1 451
2 1747 1 451
2 1748 1 455
2 1749 1 455
2 1750 1 458
2 1751 1 458
2 1752 1 459
2 1753 1 459
2 1754 1 463
2 1755 1 463
2 1756 1 466
2 1757 1 466
2 1758 1 467
2 1759 1 467
2 1760 1 471
2 1761 1 471
2 1762 1 474
2 1763 1 474
2 1764 1 475
2 1765 1 475
2 1766 1 479
2 1767 1 479
2 1768 1 482
2 1769 1 482
2 1770 1 483
2 1771 1 483
2 1772 1 485
2 1773 1 485
2 1774 1 491
2 1775 1 491
2 1776 1 494
2 1777 1 494
2 1778 1 497
2 1779 1 497
2 1780 1 500
2 1781 1 500
2 1782 1 503
2 1783 1 503
2 1784 1 507
2 1785 1 507
2 1786 1 510
2 1787 1 510
2 1788 1 511
2 1789 1 511
2 1790 1 515
2 1791 1 515
2 1792 1 518
2 1793 1 518
2 1794 1 519
2 1795 1 519
2 1796 1 523
2 1797 1 523
2 1798 1 526
2 1799 1 526
2 1800 1 527
2 1801 1 527
2 1802 1 531
2 1803 1 531
2 1804 1 534
2 1805 1 534
2 1806 1 535
2 1807 1 535
2 1808 1 539
2 1809 1 539
2 1810 1 542
2 1811 1 542
2 1812 1 543
2 1813 1 543
2 1814 1 547
2 1815 1 547
2 1816 1 550
2 1817 1 550
2 1818 1 551
2 1819 1 551
2 1820 1 555
2 1821 1 555
2 1822 1 558
2 1823 1 558
2 1824 1 559
2 1825 1 559
2 1826 1 561
2 1827 1 561
2 1828 1 564
2 1829 1 564
2 1830 1 567
2 1831 1 567
2 1832 1 571
2 1833 1 571
2 1834 1 574
2 1835 1 574
2 1836 1 575
2 1837 1 575
2 1838 1 579
2 1839 1 579
2 1840 1 582
2 1841 1 582
2 1842 1 583
2 1843 1 583
2 1844 1 587
2 1845 1 587
2 1846 1 590
2 1847 1 590
2 1848 1 591
2 1849 1 591
2 1850 1 595
2 1851 1 595
2 1852 1 598
2 1853 1 598
2 1854 1 599
2 1855 1 599
2 1856 1 605
2 1857 1 605
2 1858 1 608
2 1859 1 608
2 1860 1 609
2 1861 1 609
2 1862 1 613
2 1863 1 613
2 1864 1 616
2 1865 1 616
2 1866 1 617
2 1867 1 617
2 1868 1 621
2 1869 1 621
2 1870 1 624
2 1871 1 624
2 1872 1 625
2 1873 1 625
2 1874 1 629
2 1875 1 629
2 1876 1 632
2 1877 1 632
2 1878 1 633
2 1879 1 633
2 1880 1 635
2 1881 1 635
2 1882 1 638
2 1883 1 638
2 1884 1 641
2 1885 1 641
2 1886 1 645
2 1887 1 645
2 1888 1 648
2 1889 1 648
2 1890 1 649
2 1891 1 649
2 1892 1 653
2 1893 1 653
2 1894 1 656
2 1895 1 656
2 1896 1 659
2 1897 1 659
2 1898 1 661
2 1899 1 661
2 1900 1 663
2 1901 1 663
2 1902 1 665
2 1903 1 665
2 1904 1 667
2 1905 1 667
2 1906 1 669
2 1907 1 669
2 1908 1 671
2 1909 1 671
2 1910 1 672
2 1911 1 672
2 1912 1 673
2 1913 1 673
2 1914 1 673
2 1915 1 676
2 1916 1 676
2 1917 1 679
2 1918 1 679
2 1919 1 687
2 1920 1 687
2 1921 1 690
2 1922 1 690
2 1923 1 691
2 1924 1 691
2 1925 1 695
2 1926 1 695
2 1927 1 698
2 1928 1 698
2 1929 1 701
2 1930 1 701
2 1931 1 703
2 1932 1 703
2 1933 1 705
2 1934 1 705
2 1935 1 707
2 1936 1 707
2 1937 1 708
2 1938 1 708
2 1939 1 710
2 1940 1 710
2 1941 1 711
2 1942 1 711
2 1943 1 715
2 1944 1 715
2 1945 1 718
2 1946 1 718
2 1947 1 719
2 1948 1 719
2 1949 1 723
2 1950 1 723
2 1951 1 726
2 1952 1 726
2 1953 1 727
2 1954 1 727
2 1955 1 731
2 1956 1 731
2 1957 1 734
2 1958 1 734
2 1959 1 735
2 1960 1 735
2 1961 1 739
2 1962 1 739
2 1963 1 742
2 1964 1 742
2 1965 1 743
2 1966 1 743
2 1967 1 747
2 1968 1 747
2 1969 1 750
2 1970 1 750
2 1971 1 751
2 1972 1 751
2 1973 1 755
2 1974 1 755
2 1975 1 758
2 1976 1 758
2 1977 1 759
2 1978 1 759
2 1979 1 763
2 1980 1 763
2 1981 1 766
2 1982 1 766
2 1983 1 767
2 1984 1 767
2 1985 1 771
2 1986 1 771
2 1987 1 774
2 1988 1 774
2 1989 1 775
2 1990 1 775
2 1991 1 779
2 1992 1 779
2 1993 1 782
2 1994 1 782
2 1995 1 783
2 1996 1 783
2 1997 1 787
2 1998 1 787
2 1999 1 790
2 2000 1 790
2 2001 1 791
2 2002 1 791
2 2003 1 793
2 2004 1 793
2 2005 1 795
2 2006 1 795
2 2007 1 797
2 2008 1 797
2 2009 1 799
2 2010 1 799
2 2011 1 805
2 2012 1 805
2 2013 1 808
2 2014 1 808
2 2015 1 808
2 2016 1 811
2 2017 1 811
2 2018 1 814
2 2019 1 814
2 2020 1 817
2 2021 1 817
2 2022 1 820
2 2023 1 820
2 2024 1 823
2 2025 1 823
2 2026 1 826
2 2027 1 826
2 2028 1 826
2 2029 1 828
2 2030 1 828
2 2031 1 828
2 2032 1 831
2 2033 1 831
2 2034 1 834
2 2035 1 834
2 2036 1 834
2 2037 1 836
2 2038 1 836
2 2039 1 836
2 2040 1 839
2 2041 1 839
2 2042 1 842
2 2043 1 842
2 2044 1 842
2 2045 1 844
2 2046 1 844
2 2047 1 844
2 2048 1 847
2 2049 1 847
2 2050 1 850
2 2051 1 850
2 2052 1 850
2 2053 1 850
2 2054 1 852
2 2055 1 852
2 2056 1 852
2 2057 1 855
2 2058 1 855
2 2059 1 858
2 2060 1 858
2 2061 1 858
2 2062 1 858
2 2063 1 860
2 2064 1 860
2 2065 1 860
2 2066 1 863
2 2067 1 863
2 2068 1 866
2 2069 1 866
2 2070 1 866
2 2071 1 866
2 2072 1 868
2 2073 1 868
2 2074 1 868
2 2075 1 871
2 2076 1 871
2 2077 1 874
2 2078 1 874
2 2079 1 874
2 2080 1 874
2 2081 1 876
2 2082 1 876
2 2083 1 876
2 2084 1 879
2 2085 1 879
2 2086 1 882
2 2087 1 882
2 2088 1 882
2 2089 1 884
2 2090 1 884
2 2091 1 884
2 2092 1 887
2 2093 1 887
2 2094 1 890
2 2095 1 890
2 2096 1 890
2 2097 1 890
2 2098 1 892
2 2099 1 892
2 2100 1 892
2 2101 1 895
2 2102 1 895
2 2103 1 898
2 2104 1 898
2 2105 1 898
2 2106 1 898
2 2107 1 900
2 2108 1 900
2 2109 1 900
2 2110 1 903
2 2111 1 903
2 2112 1 906
2 2113 1 906
2 2114 1 906
2 2115 1 908
2 2116 1 908
2 2117 1 908
2 2118 1 911
2 2119 1 911
2 2120 1 914
2 2121 1 914
2 2122 1 914
2 2123 1 914
2 2124 1 916
2 2125 1 916
2 2126 1 916
2 2127 1 919
2 2128 1 919
2 2129 1 922
2 2130 1 922
2 2131 1 924
2 2132 1 924
2 2133 1 925
2 2134 1 925
2 2135 1 931
2 2136 1 931
2 2137 1 932
2 2138 1 932
2 2139 1 935
2 2140 1 935
2 2141 1 936
2 2142 1 936
2 2143 1 939
2 2144 1 939
2 2145 1 940
2 2146 1 940
2 2147 1 943
2 2148 1 943
2 2149 1 948
2 2150 1 948
2 2151 1 951
2 2152 1 951
2 2153 1 952
2 2154 1 952
2 2155 1 955
2 2156 1 955
2 2157 1 956
2 2158 1 956
2 2159 1 959
2 2160 1 959
2 2161 1 960
2 2162 1 960
2 2163 1 963
2 2164 1 963
2 2165 1 964
2 2166 1 964
2 2167 1 967
2 2168 1 967
2 2169 1 968
2 2170 1 968
2 2171 1 971
2 2172 1 971
2 2173 1 972
2 2174 1 972
2 2175 1 975
2 2176 1 975
2 2177 1 976
2 2178 1 976
2 2179 1 979
2 2180 1 979
2 2181 1 981
2 2182 1 981
2 2183 1 983
2 2184 1 983
2 2185 1 988
2 2186 1 988
2 2187 1 991
2 2188 1 991
2 2189 1 994
2 2190 1 994
2 2191 1 997
2 2192 1 997
2 2193 1 999
2 2194 1 999
2 2195 1 1000
2 2196 1 1000
2 2197 1 1002
2 2198 1 1002
2 2199 1 1002
2 2200 1 1002
2 2201 1 1004
2 2202 1 1004
2 2203 1 1007
2 2204 1 1007
2 2205 1 1009
2 2206 1 1009
2 2207 1 1010
2 2208 1 1010
2 2209 1 1011
2 2210 1 1011
2 2211 1 1022
2 2212 1 1022
2 2213 1 1022
2 2214 1 1026
2 2215 1 1026
2 2216 1 1031
2 2217 1 1031
2 2218 1 1034
2 2219 1 1034
2 2220 1 1036
2 2221 1 1036
2 2222 1 1038
2 2223 1 1038
2 2224 1 1039
2 2225 1 1039
2 2226 1 1042
2 2227 1 1042
2 2228 1 1043
2 2229 1 1043
2 2230 1 1046
2 2231 1 1046
2 2232 1 1049
2 2233 1 1049
2 2234 1 1053
2 2235 1 1053
2 2236 1 1063
2 2237 1 1063
2 2238 1 1066
2 2239 1 1066
2 2240 1 1067
2 2241 1 1067
2 2242 1 1070
2 2243 1 1070
2 2244 1 1071
2 2245 1 1071
2 2246 1 1074
2 2247 1 1074
2 2248 1 1077
2 2249 1 1077
2 2250 1 1081
2 2251 1 1081
2 2252 1 1083
2 2253 1 1083
2 2254 1 1083
2 2255 1 1084
2 2256 1 1084
2 2257 1 1091
2 2258 1 1091
2 2259 1 1091
2 2260 1 1092
2 2261 1 1092
2 2262 1 1097
2 2263 1 1097
2 2264 1 1097
2 2265 1 1098
2 2266 1 1098
2 2267 1 1103
2 2268 1 1103
2 2269 1 1104
2 2270 1 1104
2 2271 1 1109
2 2272 1 1109
2 2273 1 1109
2 2274 1 1115
2 2275 1 1115
2 2276 1 1115
2 2277 1 1121
2 2278 1 1121
2 2279 1 1122
2 2280 1 1122
2 2281 1 1129
2 2282 1 1129
2 2283 1 1129
2 2284 1 1130
2 2285 1 1130
2 2286 1 1135
2 2287 1 1135
2 2288 1 1136
2 2289 1 1136
2 2290 1 1139
2 2291 1 1139
2 2292 1 1140
2 2293 1 1140
2 2294 1 1145
2 2295 1 1145
2 2296 1 1145
2 2297 1 1146
2 2298 1 1146
2 2299 1 1150
2 2300 1 1150
2 2301 1 1152
2 2302 1 1152
0 33 5 1 1 1388
0 34 5 1 1 1390
0 35 5 1 1 1392
0 36 5 1 1 1394
0 37 5 1 1 1396
0 38 5 1 1 1398
0 39 5 1 1 1400
0 40 5 1 1 1402
0 41 5 1 1 1404
0 42 5 1 1 1406
0 43 5 1 1 1408
0 44 5 1 1 1410
0 45 5 1 1 1412
0 46 5 1 1 1414
0 47 5 1 1 1416
0 48 5 1 1 1418
0 49 7 2 2 1290 1372
0 50 5 1 1 1420
0 51 7 2 2 1307 1356
0 52 5 1 1 1422
0 53 7 2 2 1281 1380
0 54 5 1 1 1424
0 55 7 2 2 1315 1348
0 56 5 1 1 1426
0 57 7 1 2 1425 1427
0 58 5 2 1 57
0 59 7 1 2 54 56
0 60 5 1 1 59
0 61 7 2 2 1428 60
0 62 5 1 1 1430
0 63 7 1 2 1423 1431
0 64 5 2 1 63
0 65 7 1 2 52 62
0 66 5 1 1 65
0 67 7 2 2 1432 66
0 68 5 1 1 1434
0 69 7 1 2 1421 1435
0 70 5 2 1 69
0 71 7 2 2 1298 1364
0 72 5 1 1 1438
0 73 7 1 2 50 68
0 74 5 1 1 73
0 75 7 2 2 1436 74
0 76 5 1 1 1440
0 77 7 1 2 1439 1441
0 78 5 2 1 77
0 79 7 2 2 1437 1442
0 80 5 1 1 1444
0 81 7 2 2 1429 1433
0 82 5 1 1 1446
0 83 7 2 2 1299 1373
0 84 5 1 1 1448
0 85 7 2 2 1308 1365
0 86 5 1 1 1450
0 87 7 2 2 1291 1381
0 88 5 1 1 1452
0 89 7 2 2 1316 1357
0 90 5 1 1 1454
0 91 7 1 2 1453 1455
0 92 5 2 1 91
0 93 7 1 2 88 90
0 94 5 1 1 93
0 95 7 2 2 1456 94
0 96 5 1 1 1458
0 97 7 1 2 1451 1459
0 98 5 2 1 97
0 99 7 1 2 86 96
0 100 5 1 1 99
0 101 7 2 2 1460 100
0 102 5 1 1 1462
0 103 7 1 2 1449 1463
0 104 5 2 1 103
0 105 7 1 2 84 102
0 106 5 1 1 105
0 107 7 2 2 1464 106
0 108 5 1 1 1466
0 109 7 1 2 82 1467
0 110 5 2 1 109
0 111 7 1 2 1447 108
0 112 5 1 1 111
0 113 7 2 2 1468 112
0 114 5 1 1 1470
0 115 7 1 2 80 1471
0 116 5 2 1 115
0 117 7 2 2 1273 1382
0 118 5 1 1 1474
0 119 7 2 2 1317 1323
0 120 5 1 1 1476
0 121 7 2 2 1309 1331
0 122 5 1 1 1478
0 123 7 2 2 1477 1479
0 124 5 2 1 1480
0 125 7 2 2 1339 1481
0 126 5 2 1 1484
0 127 7 1 2 1475 1485
0 128 5 2 1 127
0 129 7 2 2 1318 1340
0 130 5 1 1 1490
0 131 7 1 2 118 1486
0 132 5 1 1 131
0 133 7 2 2 1488 132
0 134 5 1 1 1492
0 135 7 1 2 1491 1493
0 136 5 2 1 135
0 137 7 2 2 1489 1494
0 138 5 1 1 1496
0 139 7 1 2 72 76
0 140 5 1 1 139
0 141 7 2 2 1443 140
0 142 5 1 1 1498
0 143 7 1 2 138 1499
0 144 5 2 1 143
0 145 7 2 2 1300 1358
0 146 5 1 1 1502
0 147 7 1 2 130 134
0 148 5 1 1 147
0 149 7 2 2 1495 148
0 150 5 1 1 1504
0 151 7 1 2 1503 1505
0 152 5 2 1 151
0 153 7 2 2 1310 1349
0 154 5 1 1 1508
0 155 7 1 2 146 150
0 156 5 1 1 155
0 157 7 2 2 1506 156
0 158 5 1 1 1510
0 159 7 1 2 1509 1511
0 160 5 2 1 159
0 161 7 2 2 1507 1512
0 162 5 1 1 1514
0 163 7 1 2 1497 142
0 164 5 1 1 163
0 165 7 2 2 1500 164
0 166 5 1 1 1516
0 167 7 1 2 162 1517
0 168 5 2 1 167
0 169 7 2 2 1501 1518
0 170 5 1 1 1520
0 171 7 1 2 1445 114
0 172 5 1 1 171
0 173 7 2 2 1472 172
0 174 5 1 1 1522
0 175 7 1 2 170 1523
0 176 5 2 1 175
0 177 7 2 2 1473 1524
0 178 5 1 1 1526
0 179 7 2 2 1465 1469
0 180 5 1 1 1528
0 181 7 2 2 1457 1461
0 182 5 1 1 1530
0 183 7 2 2 1311 1374
0 184 5 2 1 1532
0 185 7 2 2 1301 1383
0 186 5 1 1 1536
0 187 7 2 2 1319 1366
0 188 5 1 1 1538
0 189 7 1 2 1537 1539
0 190 5 2 1 189
0 191 7 1 2 186 188
0 192 5 1 1 191
0 193 7 2 2 1540 192
0 194 5 1 1 1542
0 195 7 1 2 1533 1543
0 196 5 2 1 195
0 197 7 1 2 1534 194
0 198 5 1 1 197
0 199 7 2 2 1544 198
0 200 5 1 1 1546
0 201 7 1 2 182 1547
0 202 5 2 1 201
0 203 7 1 2 1531 200
0 204 5 1 1 203
0 205 7 2 2 1548 204
0 206 5 1 1 1550
0 207 7 1 2 180 1551
0 208 5 2 1 207
0 209 7 1 2 1529 206
0 210 5 1 1 209
0 211 7 2 2 1552 210
0 212 5 1 1 1554
0 213 7 1 2 178 1555
0 214 5 2 1 213
0 215 7 2 2 1282 1375
0 216 5 1 1 1558
0 217 7 2 2 1292 1367
0 218 5 1 1 1560
0 219 7 1 2 1559 1561
0 220 5 2 1 219
0 221 7 1 2 154 158
0 222 5 1 1 221
0 223 7 2 2 1513 222
0 224 5 1 1 1564
0 225 7 1 2 216 218
0 226 5 1 1 225
0 227 7 2 2 1562 226
0 228 5 1 1 1566
0 229 7 1 2 1565 1567
0 230 5 2 1 229
0 231 7 2 2 1563 1568
0 232 5 1 1 1570
0 233 7 1 2 1515 166
0 234 5 1 1 233
0 235 7 2 2 1519 234
0 236 5 1 1 1572
0 237 7 1 2 232 1573
0 238 5 2 1 237
0 239 7 2 2 1302 1350
0 240 5 1 1 1576
0 241 7 2 2 1274 1376
0 242 5 1 1 1578
0 243 7 1 2 1577 1579
0 244 5 2 1 243
0 245 7 2 2 1265 1384
0 246 5 1 1 1582
0 247 7 2 2 1293 1359
0 248 5 1 1 1584
0 249 7 1 2 1312 1341
0 250 5 1 1 249
0 251 7 1 2 1482 250
0 252 5 1 1 251
0 253 7 2 2 1487 252
0 254 5 1 1 1586
0 255 7 1 2 1585 1587
0 256 5 2 1 255
0 257 7 1 2 248 254
0 258 5 1 1 257
0 259 7 2 2 1588 258
0 260 5 1 1 1590
0 261 7 1 2 1583 1591
0 262 5 2 1 261
0 263 7 1 2 246 260
0 264 5 1 1 263
0 265 7 2 2 1592 264
0 266 5 1 1 1594
0 267 7 1 2 240 242
0 268 5 1 1 267
0 269 7 2 2 1580 268
0 270 5 1 1 1596
0 271 7 1 2 1595 1597
0 272 5 2 1 271
0 273 7 2 2 1581 1598
0 274 5 1 1 1600
0 275 7 1 2 224 228
0 276 5 1 1 275
0 277 7 2 2 1569 276
0 278 5 1 1 1602
0 279 7 1 2 274 1603
0 280 5 2 1 279
0 281 7 2 2 1320 1332
0 282 5 1 1 1606
0 283 7 2 2 1283 1368
0 284 5 1 1 1608
0 285 7 1 2 1607 1609
0 286 5 2 1 285
0 287 7 1 2 266 270
0 288 5 1 1 287
0 289 7 2 2 1599 288
0 290 5 1 1 1612
0 291 7 1 2 282 284
0 292 5 1 1 291
0 293 7 2 2 1610 292
0 294 5 1 1 1614
0 295 7 1 2 1613 1615
0 296 5 2 1 295
0 297 7 2 2 1611 1616
0 298 5 1 1 1618
0 299 7 1 2 1601 278
0 300 5 1 1 299
0 301 7 2 2 1604 300
0 302 5 1 1 1620
0 303 7 1 2 298 1621
0 304 5 2 1 303
0 305 7 2 2 1605 1622
0 306 5 1 1 1624
0 307 7 1 2 1571 236
0 308 5 1 1 307
0 309 7 2 2 1574 308
0 310 5 1 1 1626
0 311 7 1 2 306 1627
0 312 5 2 1 311
0 313 7 2 2 1575 1628
0 314 5 1 1 1630
0 315 7 1 2 1521 174
0 316 5 1 1 315
0 317 7 2 2 1525 316
0 318 5 1 1 1632
0 319 7 1 2 314 1633
0 320 5 2 1 319
0 321 7 2 2 1589 1593
0 322 5 1 1 1636
0 323 7 1 2 1619 302
0 324 5 1 1 323
0 325 7 2 2 1623 324
0 326 5 1 1 1638
0 327 7 1 2 322 1639
0 328 5 2 1 327
0 329 7 2 2 1303 1342
0 330 5 1 1 1642
0 331 7 2 2 1294 1351
0 332 5 1 1 1644
0 333 7 1 2 1643 1645
0 334 5 2 1 333
0 335 7 2 2 1266 1377
0 336 5 1 1 1648
0 337 7 1 2 330 332
0 338 5 1 1 337
0 339 7 2 2 1646 338
0 340 5 1 1 1650
0 341 7 1 2 1649 1651
0 342 5 2 1 341
0 343 7 2 2 1647 1652
0 344 5 1 1 1654
0 345 7 2 2 1275 1369
0 346 5 1 1 1656
0 347 7 2 2 32 1385
0 348 5 1 1 1658
0 349 7 1 2 1657 1659
0 350 5 2 1 349
0 351 7 2 2 1295 1333
0 352 5 1 1 1662
0 353 7 2 2 1258 1352
0 354 5 1 1 1664
0 355 7 2 2 1276 1334
0 356 5 1 1 1666
0 357 7 2 2 1665 1667
0 358 5 2 1 1668
0 359 7 2 2 1284 1669
0 360 5 2 1 1672
0 361 7 2 2 1663 1673
0 362 5 2 1 1676
0 363 7 2 2 1304 1677
0 364 5 2 1 1680
0 365 7 2 2 1285 1360
0 366 5 1 1 1684
0 367 7 1 2 1681 1685
0 368 5 2 1 367
0 369 7 1 2 1682 366
0 370 5 1 1 369
0 371 7 2 2 1686 370
0 372 5 1 1 1688
0 373 7 1 2 120 122
0 374 5 1 1 373
0 375 7 2 2 1483 374
0 376 5 1 1 1690
0 377 7 1 2 1689 1691
0 378 5 2 1 377
0 379 7 1 2 372 376
0 380 5 1 1 379
0 381 7 2 2 1692 380
0 382 5 1 1 1694
0 383 7 1 2 346 348
0 384 5 1 1 383
0 385 7 2 2 1660 384
0 386 5 1 1 1696
0 387 7 1 2 1695 1697
0 388 5 2 1 387
0 389 7 2 2 1661 1698
0 390 5 1 1 1700
0 391 7 1 2 344 390
0 392 5 2 1 391
0 393 7 2 2 1687 1693
0 394 5 1 1 1704
0 395 7 1 2 1655 1701
0 396 5 1 1 395
0 397 7 2 2 1702 396
0 398 5 1 1 1706
0 399 7 1 2 394 1707
0 400 5 2 1 399
0 401 7 2 2 1703 1708
0 402 5 1 1 1710
0 403 7 1 2 1637 326
0 404 5 1 1 403
0 405 7 2 2 1640 404
0 406 5 1 1 1712
0 407 7 1 2 402 1713
0 408 5 2 1 407
0 409 7 2 2 1641 1714
0 410 5 1 1 1716
0 411 7 1 2 1625 310
0 412 5 1 1 411
0 413 7 2 2 1629 412
0 414 5 1 1 1718
0 415 7 1 2 410 1719
0 416 5 2 1 415
0 417 7 1 2 290 294
0 418 5 1 1 417
0 419 7 2 2 1617 418
0 420 5 1 1 1722
0 421 7 1 2 1705 398
0 422 5 1 1 421
0 423 7 2 2 1709 422
0 424 5 1 1 1724
0 425 7 1 2 1723 1725
0 426 5 2 1 425
0 427 7 1 2 336 340
0 428 5 1 1 427
0 429 7 2 2 1653 428
0 430 5 1 1 1728
0 431 7 1 2 382 386
0 432 5 1 1 431
0 433 7 2 2 1699 432
0 434 5 1 1 1730
0 435 7 1 2 1729 1731
0 436 5 2 1 435
0 437 7 2 2 1286 1353
0 438 5 1 1 1734
0 439 7 2 2 1277 1361
0 440 5 1 1 1736
0 441 7 1 2 1735 1737
0 442 5 2 1 441
0 443 7 2 2 1267 1370
0 444 5 1 1 1740
0 445 7 1 2 438 440
0 446 5 1 1 445
0 447 7 2 2 1738 446
0 448 5 1 1 1742
0 449 7 1 2 1741 1743
0 450 5 2 1 449
0 451 7 2 2 1739 1744
0 452 5 1 1 1746
0 453 7 1 2 430 434
0 454 5 1 1 453
0 455 7 2 2 1732 454
0 456 5 1 1 1748
0 457 7 1 2 452 1749
0 458 5 2 1 457
0 459 7 2 2 1733 1750
0 460 5 1 1 1752
0 461 7 1 2 420 424
0 462 5 1 1 461
0 463 7 2 2 1726 462
0 464 5 1 1 1754
0 465 7 1 2 460 1755
0 466 5 2 1 465
0 467 7 2 2 1727 1756
0 468 5 1 1 1758
0 469 7 1 2 1711 406
0 470 5 1 1 469
0 471 7 2 2 1715 470
0 472 5 1 1 1760
0 473 7 1 2 468 1761
0 474 5 2 1 473
0 475 7 2 2 1259 1378
0 476 5 1 1 1764
0 477 7 1 2 444 448
0 478 5 1 1 477
0 479 7 2 2 1745 478
0 480 5 1 1 1766
0 481 7 1 2 1765 1767
0 482 5 2 1 481
0 483 7 2 2 1313 1324
0 484 5 1 1 1770
0 485 7 2 2 1296 1343
0 486 5 1 1 1772
0 487 7 1 2 1305 1335
0 488 5 1 1 487
0 489 7 1 2 1678 488
0 490 5 1 1 489
0 491 7 2 2 1683 490
0 492 5 1 1 1774
0 493 7 1 2 1773 1775
0 494 5 2 1 493
0 495 7 1 2 486 492
0 496 5 1 1 495
0 497 7 2 2 1776 496
0 498 5 1 1 1778
0 499 7 1 2 1771 1779
0 500 5 2 1 499
0 501 7 1 2 484 498
0 502 5 1 1 501
0 503 7 2 2 1780 502
0 504 5 1 1 1782
0 505 7 1 2 476 480
0 506 5 1 1 505
0 507 7 2 2 1768 506
0 508 5 1 1 1784
0 509 7 1 2 1783 1785
0 510 5 2 1 509
0 511 7 2 2 1769 1786
0 512 5 1 1 1788
0 513 7 1 2 1747 456
0 514 5 1 1 513
0 515 7 2 2 1751 514
0 516 5 1 1 1790
0 517 7 1 2 512 1791
0 518 5 2 1 517
0 519 7 2 2 1777 1781
0 520 5 1 1 1794
0 521 7 1 2 1789 516
0 522 5 1 1 521
0 523 7 2 2 1792 522
0 524 5 1 1 1796
0 525 7 1 2 520 1797
0 526 5 2 1 525
0 527 7 2 2 1793 1798
0 528 5 1 1 1800
0 529 7 1 2 1753 464
0 530 5 1 1 529
0 531 7 2 2 1757 530
0 532 5 1 1 1802
0 533 7 1 2 528 1803
0 534 5 2 1 533
0 535 7 2 2 1287 1344
0 536 5 1 1 1806
0 537 7 1 2 352 1674
0 538 5 1 1 537
0 539 7 2 2 1679 538
0 540 5 1 1 1808
0 541 7 1 2 1807 1809
0 542 5 2 1 541
0 543 7 2 2 1306 1325
0 544 5 1 1 1812
0 545 7 1 2 536 540
0 546 5 1 1 545
0 547 7 2 2 1810 546
0 548 5 1 1 1814
0 549 7 1 2 1813 1815
0 550 5 2 1 549
0 551 7 2 2 1811 1816
0 552 5 1 1 1818
0 553 7 1 2 504 508
0 554 5 1 1 553
0 555 7 2 2 1787 554
0 556 5 1 1 1820
0 557 7 1 2 552 1821
0 558 5 2 1 557
0 559 7 2 2 1278 1354
0 560 5 1 1 1824
0 561 7 2 2 1260 1371
0 562 5 1 1 1826
0 563 7 1 2 1825 1827
0 564 5 2 1 563
0 565 7 1 2 544 548
0 566 5 1 1 565
0 567 7 2 2 1817 566
0 568 5 1 1 1830
0 569 7 1 2 560 562
0 570 5 1 1 569
0 571 7 2 2 1828 570
0 572 5 1 1 1832
0 573 7 1 2 1831 1833
0 574 5 2 1 573
0 575 7 2 2 1829 1834
0 576 5 1 1 1836
0 577 7 1 2 1819 556
0 578 5 1 1 577
0 579 7 2 2 1822 578
0 580 5 1 1 1838
0 581 7 1 2 576 1839
0 582 5 2 1 581
0 583 7 2 2 1823 1840
0 584 5 1 1 1842
0 585 7 1 2 1795 524
0 586 5 1 1 585
0 587 7 2 2 1799 586
0 588 5 1 1 1844
0 589 7 1 2 584 1845
0 590 5 2 1 589
0 591 7 2 2 1268 1362
0 592 5 1 1 1848
0 593 7 1 2 568 572
0 594 5 1 1 593
0 595 7 2 2 1835 594
0 596 5 1 1 1850
0 597 7 1 2 1849 1851
0 598 5 2 1 597
0 599 7 2 2 1279 1345
0 600 5 1 1 1854
0 601 7 1 2 1288 1336
0 602 5 1 1 601
0 603 7 1 2 1670 602
0 604 5 1 1 603
0 605 7 2 2 1675 604
0 606 5 1 1 1856
0 607 7 1 2 1855 1857
0 608 5 2 1 607
0 609 7 2 2 1297 1326
0 610 5 1 1 1860
0 611 7 1 2 600 606
0 612 5 1 1 611
0 613 7 2 2 1858 612
0 614 5 1 1 1862
0 615 7 1 2 1861 1863
0 616 5 2 1 615
0 617 7 2 2 1859 1864
0 618 5 1 1 1866
0 619 7 1 2 592 596
0 620 5 1 1 619
0 621 7 2 2 1852 620
0 622 5 1 1 1868
0 623 7 1 2 618 1869
0 624 5 2 1 623
0 625 7 2 2 1853 1870
0 626 5 1 1 1872
0 627 7 1 2 1837 580
0 628 5 1 1 627
0 629 7 2 2 1841 628
0 630 5 1 1 1874
0 631 7 1 2 626 1875
0 632 5 2 1 631
0 633 7 2 2 1261 1363
0 634 5 1 1 1878
0 635 7 2 2 1269 1355
0 636 5 1 1 1880
0 637 7 1 2 1879 1881
0 638 5 2 1 637
0 639 7 1 2 610 614
0 640 5 1 1 639
0 641 7 2 2 1865 640
0 642 5 1 1 1884
0 643 7 1 2 634 636
0 644 5 1 1 643
0 645 7 2 2 1882 644
0 646 5 1 1 1886
0 647 7 1 2 1885 1887
0 648 5 2 1 647
0 649 7 2 2 1883 1888
0 650 5 1 1 1890
0 651 7 1 2 1867 622
0 652 5 1 1 651
0 653 7 2 2 1871 652
0 654 5 1 1 1892
0 655 7 1 2 650 1893
0 656 5 2 1 655
0 657 7 1 2 642 646
0 658 5 1 1 657
0 659 7 2 2 1889 658
0 660 5 1 1 1896
0 661 7 2 2 1270 1346
0 662 5 1 1 1898
0 663 7 2 2 1289 1327
0 664 5 1 1 1900
0 665 7 2 2 1899 1901
0 666 5 1 1 1902
0 667 7 2 2 1271 1337
0 668 5 1 1 1904
0 669 7 2 2 1262 1347
0 670 5 1 1 1906
0 671 7 2 2 1905 1907
0 672 5 2 1 1908
0 673 7 3 2 666 1910
0 674 5 1 1 1912
0 675 7 1 2 1897 674
0 676 5 2 1 675
0 677 7 1 2 354 356
0 678 5 1 1 677
0 679 7 2 2 1671 678
0 680 5 1 1 1917
0 681 7 1 2 662 664
0 682 5 1 1 681
0 683 7 1 2 1913 682
0 684 5 1 1 683
0 685 7 1 2 1903 1909
0 686 5 1 1 685
0 687 7 2 2 684 686
0 688 5 1 1 1919
0 689 7 1 2 1918 688
0 690 5 2 1 689
0 691 7 2 2 1280 1328
0 692 5 1 1 1923
0 693 7 1 2 668 670
0 694 5 1 1 693
0 695 7 2 2 1911 694
0 696 5 1 1 1925
0 697 7 1 2 1924 1926
0 698 5 2 1 697
0 699 7 1 2 692 696
0 700 5 1 1 699
0 701 7 2 2 1927 700
0 702 5 1 1 1929
0 703 7 2 2 1263 1338
0 704 5 1 1 1931
0 705 7 2 2 1272 1329
0 706 5 1 1 1933
0 707 7 2 2 1932 1934
0 708 5 2 1 1935
0 709 7 1 2 1930 1936
0 710 5 2 1 709
0 711 7 2 2 1928 1939
0 712 5 1 1 1941
0 713 7 1 2 680 1920
0 714 5 1 1 713
0 715 7 2 2 1921 714
0 716 5 1 1 1943
0 717 7 1 2 712 1944
0 718 5 2 1 717
0 719 7 2 2 1922 1945
0 720 5 1 1 1947
0 721 7 1 2 660 1914
0 722 5 1 1 721
0 723 7 2 2 1915 722
0 724 5 1 1 1949
0 725 7 1 2 720 1950
0 726 5 2 1 725
0 727 7 2 2 1916 1951
0 728 5 1 1 1953
0 729 7 1 2 1891 654
0 730 5 1 1 729
0 731 7 2 2 1894 730
0 732 5 1 1 1955
0 733 7 1 2 728 1956
0 734 5 2 1 733
0 735 7 2 2 1895 1957
0 736 5 1 1 1959
0 737 7 1 2 1873 630
0 738 5 1 1 737
0 739 7 2 2 1876 738
0 740 5 1 1 1961
0 741 7 1 2 736 1962
0 742 5 2 1 741
0 743 7 2 2 1877 1963
0 744 5 1 1 1965
0 745 7 1 2 1843 588
0 746 5 1 1 745
0 747 7 2 2 1846 746
0 748 5 1 1 1967
0 749 7 1 2 744 1968
0 750 5 2 1 749
0 751 7 2 2 1847 1969
0 752 5 1 1 1971
0 753 7 1 2 1801 532
0 754 5 1 1 753
0 755 7 2 2 1804 754
0 756 5 1 1 1973
0 757 7 1 2 752 1974
0 758 5 2 1 757
0 759 7 2 2 1805 1975
0 760 5 1 1 1977
0 761 7 1 2 1759 472
0 762 5 1 1 761
0 763 7 2 2 1762 762
0 764 5 1 1 1979
0 765 7 1 2 760 1980
0 766 5 2 1 765
0 767 7 2 2 1763 1981
0 768 5 1 1 1983
0 769 7 1 2 1717 414
0 770 5 1 1 769
0 771 7 2 2 1720 770
0 772 5 1 1 1985
0 773 7 1 2 768 1986
0 774 5 2 1 773
0 775 7 2 2 1721 1987
0 776 5 1 1 1989
0 777 7 1 2 1631 318
0 778 5 1 1 777
0 779 7 2 2 1634 778
0 780 5 1 1 1991
0 781 7 1 2 776 1992
0 782 5 2 1 781
0 783 7 2 2 1635 1993
0 784 5 1 1 1995
0 785 7 1 2 1527 212
0 786 5 1 1 785
0 787 7 2 2 1556 786
0 788 5 1 1 1997
0 789 7 1 2 784 1998
0 790 5 2 1 789
0 791 7 2 2 1557 1999
0 792 5 1 1 2001
0 793 7 2 2 1549 1553
0 794 5 1 1 2003
0 795 7 2 2 1541 1545
0 796 5 1 1 2005
0 797 7 2 2 1314 1386
0 798 5 1 1 2007
0 799 7 2 2 1321 1379
0 800 5 1 1 2009
0 801 7 1 2 798 2010
0 802 5 1 1 801
0 803 7 1 2 2008 800
0 804 5 1 1 803
0 805 7 2 2 802 804
0 806 5 1 1 2011
0 807 7 1 2 796 806
0 808 5 3 1 807
0 809 7 1 2 2006 2012
0 810 5 1 1 809
0 811 7 2 2 2013 810
0 812 5 1 1 2016
0 813 7 1 2 794 2017
0 814 5 2 1 813
0 815 7 1 2 2004 812
0 816 5 1 1 815
0 817 7 2 2 2018 816
0 818 5 1 1 2020
0 819 7 1 2 792 2021
0 820 5 2 1 819
0 821 7 1 2 2002 818
0 822 5 1 1 821
0 823 7 2 2 2022 822
0 824 5 1 1 2024
0 825 7 1 2 1415 824
0 826 5 3 1 825
0 827 7 1 2 46 2025
0 828 5 3 1 827
0 829 7 1 2 1996 788
0 830 5 1 1 829
0 831 7 2 2 2000 830
0 832 5 1 1 2032
0 833 7 1 2 1413 832
0 834 5 3 1 833
0 835 7 1 2 45 2033
0 836 5 3 1 835
0 837 7 1 2 1990 780
0 838 5 1 1 837
0 839 7 2 2 1994 838
0 840 5 1 1 2040
0 841 7 1 2 1411 840
0 842 5 3 1 841
0 843 7 1 2 44 2041
0 844 5 3 1 843
0 845 7 1 2 1984 772
0 846 5 1 1 845
0 847 7 2 2 1988 846
0 848 5 1 1 2048
0 849 7 1 2 1409 848
0 850 5 4 1 849
0 851 7 1 2 43 2049
0 852 5 3 1 851
0 853 7 1 2 1978 764
0 854 5 1 1 853
0 855 7 2 2 1982 854
0 856 5 1 1 2057
0 857 7 1 2 1407 856
0 858 5 4 1 857
0 859 7 1 2 42 2058
0 860 5 3 1 859
0 861 7 1 2 1972 756
0 862 5 1 1 861
0 863 7 2 2 1976 862
0 864 5 1 1 2066
0 865 7 1 2 1405 864
0 866 5 4 1 865
0 867 7 1 2 41 2067
0 868 5 3 1 867
0 869 7 1 2 1966 748
0 870 5 1 1 869
0 871 7 2 2 1970 870
0 872 5 1 1 2075
0 873 7 1 2 1403 872
0 874 5 4 1 873
0 875 7 1 2 40 2076
0 876 5 3 1 875
0 877 7 1 2 1960 740
0 878 5 1 1 877
0 879 7 2 2 1964 878
0 880 5 1 1 2084
0 881 7 1 2 1401 880
0 882 5 3 1 881
0 883 7 1 2 39 2085
0 884 5 3 1 883
0 885 7 1 2 1954 732
0 886 5 1 1 885
0 887 7 2 2 1958 886
0 888 5 1 1 2092
0 889 7 1 2 1399 888
0 890 5 4 1 889
0 891 7 1 2 38 2093
0 892 5 3 1 891
0 893 7 1 2 1948 724
0 894 5 1 1 893
0 895 7 2 2 1952 894
0 896 5 1 1 2101
0 897 7 1 2 1397 896
0 898 5 4 1 897
0 899 7 1 2 37 2102
0 900 5 3 1 899
0 901 7 1 2 1942 716
0 902 5 1 1 901
0 903 7 2 2 1946 902
0 904 5 1 1 2110
0 905 7 1 2 1395 904
0 906 5 3 1 905
0 907 7 1 2 36 2111
0 908 5 3 1 907
0 909 7 1 2 702 1937
0 910 5 1 1 909
0 911 7 2 2 1940 910
0 912 5 1 1 2118
0 913 7 1 2 1393 912
0 914 5 4 1 913
0 915 7 1 2 35 2119
0 916 5 3 1 915
0 917 7 1 2 704 706
0 918 5 1 1 917
0 919 7 2 2 1938 918
0 920 5 1 1 2127
0 921 7 1 2 1391 920
0 922 5 2 1 921
0 923 7 1 2 34 2128
0 924 5 2 1 923
0 925 7 2 2 1264 1330
0 926 5 1 1 2133
0 927 7 1 2 33 2134
0 928 5 1 1 927
0 929 7 1 2 2131 928
0 930 5 1 1 929
0 931 7 2 2 2129 930
0 932 5 2 1 2135
0 933 7 1 2 2124 2137
0 934 5 1 1 933
0 935 7 2 2 2120 934
0 936 5 2 1 2139
0 937 7 1 2 2115 2141
0 938 5 1 1 937
0 939 7 2 2 2112 938
0 940 5 2 1 2143
0 941 7 1 2 2107 2145
0 942 5 1 1 941
0 943 7 2 2 2103 942
0 944 5 1 1 2147
0 945 7 1 2 2098 944
0 946 5 1 1 945
0 947 7 1 2 2094 946
0 948 5 2 1 947
0 949 7 1 2 2089 2149
0 950 5 1 1 949
0 951 7 2 2 2086 950
0 952 5 2 1 2151
0 953 7 1 2 2081 2153
0 954 5 1 1 953
0 955 7 2 2 2077 954
0 956 5 2 1 2155
0 957 7 1 2 2072 2157
0 958 5 1 1 957
0 959 7 2 2 2068 958
0 960 5 2 1 2159
0 961 7 1 2 2063 2161
0 962 5 1 1 961
0 963 7 2 2 2059 962
0 964 5 2 1 2163
0 965 7 1 2 2054 2165
0 966 5 1 1 965
0 967 7 2 2 2050 966
0 968 5 2 1 2167
0 969 7 1 2 2045 2169
0 970 5 1 1 969
0 971 7 2 2 2042 970
0 972 5 2 1 2171
0 973 7 1 2 2037 2173
0 974 5 1 1 973
0 975 7 2 2 2034 974
0 976 5 2 1 2175
0 977 7 1 2 2029 2177
0 978 5 1 1 977
0 979 7 2 2 2026 978
0 980 5 1 1 2179
0 981 7 2 2 2019 2023
0 982 5 1 1 2181
0 983 7 2 2 1322 1387
0 984 5 1 1 2183
0 985 7 1 2 1535 2014
0 986 5 1 1 985
0 987 7 1 2 2184 986
0 988 5 2 1 987
0 989 7 1 2 984 2015
0 990 5 1 1 989
0 991 7 2 2 2185 990
0 992 5 1 1 2187
0 993 7 1 2 982 2188
0 994 5 2 1 993
0 995 7 1 2 2182 992
0 996 5 1 1 995
0 997 7 2 2 2189 996
0 998 5 1 1 2191
0 999 7 2 2 47 2192
0 1000 5 2 1 2193
0 1001 7 1 2 1417 998
0 1002 5 4 1 1001
0 1003 7 1 2 2195 2197
0 1004 5 2 1 1003
0 1005 7 1 2 980 2201
0 1006 5 1 1 1005
0 1007 7 2 2 2186 2190
0 1008 5 1 1 2203
0 1009 7 2 2 1419 2204
0 1010 5 2 1 2205
0 1011 7 2 2 2198 2180
0 1012 5 1 1 2209
0 1013 7 1 2 2207 1012
0 1014 7 1 2 1006 1013
0 1015 5 1 1 1014
0 1016 7 1 2 2194 2206
0 1017 7 1 2 2210 1016
0 1018 5 1 1 1017
0 1019 7 1 2 1015 1018
0 1020 5 1 1 1019
0 1021 7 1 2 48 1008
0 1022 5 3 1 1021
0 1023 7 1 2 1389 926
0 1024 5 1 1 1023
0 1025 7 1 2 2130 1024
0 1026 5 2 1 1025
0 1027 7 1 2 2132 2214
0 1028 7 1 2 2125 1027
0 1029 5 1 1 1028
0 1030 7 1 2 2121 1029
0 1031 5 2 1 1030
0 1032 7 1 2 2116 2216
0 1033 5 1 1 1032
0 1034 7 2 2 2113 1033
0 1035 5 1 1 2218
0 1036 7 2 2 2108 1035
0 1037 5 1 1 2220
0 1038 7 2 2 2104 1037
0 1039 5 2 1 2222
0 1040 7 1 2 2099 2224
0 1041 5 1 1 1040
0 1042 7 2 2 2095 1041
0 1043 5 2 1 2226
0 1044 7 1 2 2090 2228
0 1045 5 1 1 1044
0 1046 7 2 2 2087 1045
0 1047 5 1 1 2230
0 1048 7 1 2 2082 1047
0 1049 5 2 1 1048
0 1050 7 1 2 2078 2232
0 1051 5 1 1 1050
0 1052 7 1 2 2073 1051
0 1053 5 2 1 1052
0 1054 7 1 2 2069 2234
0 1055 5 1 1 1054
0 1056 7 1 2 2064 1055
0 1057 5 1 1 1056
0 1058 7 1 2 2060 1057
0 1059 5 1 1 1058
0 1060 7 1 2 2055 1059
0 1061 5 1 1 1060
0 1062 7 1 2 2051 1061
0 1063 5 2 1 1062
0 1064 7 1 2 2046 2236
0 1065 5 1 1 1064
0 1066 7 2 2 2043 1065
0 1067 5 2 1 2238
0 1068 7 1 2 2038 2240
0 1069 5 1 1 1068
0 1070 7 2 2 2035 1069
0 1071 5 2 1 2242
0 1072 7 1 2 2030 2244
0 1073 5 1 1 1072
0 1074 7 2 2 2027 1073
0 1075 5 1 1 2246
0 1076 7 1 2 2196 1075
0 1077 5 2 1 1076
0 1078 7 1 2 2199 2208
0 1079 7 1 2 2248 1078
0 1080 5 1 1 1079
0 1081 7 2 2 2211 1080
0 1082 5 1 1 2250
0 1083 7 3 2 2028 2031
0 1084 5 2 1 2252
0 1085 7 1 2 2176 2255
0 1086 5 1 1 1085
0 1087 7 1 2 2178 2253
0 1088 5 1 1 1087
0 1089 7 1 2 1086 1088
0 1090 5 1 1 1089
0 1091 7 3 2 2036 2039
0 1092 5 2 1 2257
0 1093 7 1 2 2172 2258
0 1094 5 1 1 1093
0 1095 7 1 2 2174 2260
0 1096 5 1 1 1095
0 1097 7 3 2 2044 2047
0 1098 5 2 1 2262
0 1099 7 1 2 2168 2263
0 1100 5 1 1 1099
0 1101 7 1 2 2170 2265
0 1102 5 1 1 1101
0 1103 7 2 2 2052 2056
0 1104 5 2 1 2267
0 1105 7 1 2 2166 2269
0 1106 5 1 1 1105
0 1107 7 1 2 2164 2268
0 1108 5 1 1 1107
0 1109 7 3 2 2061 2065
0 1110 5 1 1 2271
0 1111 7 1 2 2160 2272
0 1112 5 1 1 1111
0 1113 7 1 2 2162 1110
0 1114 5 1 1 1113
0 1115 7 3 2 2070 2074
0 1116 5 1 1 2274
0 1117 7 1 2 2158 1116
0 1118 5 1 1 1117
0 1119 7 1 2 2156 2275
0 1120 5 1 1 1119
0 1121 7 2 2 2079 2083
0 1122 5 2 1 2277
0 1123 7 1 2 2152 2279
0 1124 5 1 1 1123
0 1125 7 1 2 2154 2278
0 1126 5 1 1 1125
0 1127 7 1 2 1124 1126
0 1128 5 1 1 1127
0 1129 7 3 2 2088 2091
0 1130 5 2 1 2281
0 1131 7 1 2 2096 2284
0 1132 5 1 1 1131
0 1133 7 1 2 2150 2282
0 1134 5 1 1 1133
0 1135 7 2 2 2097 2100
0 1136 5 2 1 2286
0 1137 7 1 2 2148 2288
0 1138 5 1 1 1137
0 1139 7 2 2 2105 2109
0 1140 5 2 1 2290
0 1141 7 1 2 2144 2291
0 1142 5 1 1 1141
0 1143 7 1 2 2146 2292
0 1144 5 1 1 1143
0 1145 7 3 2 2114 2117
0 1146 5 2 1 2294
0 1147 7 1 2 2140 2295
0 1148 5 1 1 1147
0 1149 7 1 2 2122 2126
0 1150 5 2 1 1149
0 1151 7 1 2 2136 2299
0 1152 5 2 1 1151
0 1153 7 1 2 2215 2300
0 1154 5 1 1 1153
0 1155 7 1 2 2138 1154
0 1156 5 1 1 1155
0 1157 7 1 2 2301 1156
0 1158 5 1 1 1157
0 1159 7 1 2 2142 2297
0 1160 5 1 1 1159
0 1161 7 1 2 1158 1160
0 1162 7 1 2 1148 1161
0 1163 7 1 2 1144 1162
0 1164 7 1 2 1142 1163
0 1165 5 1 1 1164
0 1166 7 1 2 1138 1165
0 1167 7 1 2 1134 1166
0 1168 7 1 2 1132 1167
0 1169 5 1 1 1168
0 1170 7 1 2 1128 1169
0 1171 7 1 2 1120 1170
0 1172 7 1 2 1118 1171
0 1173 7 1 2 1114 1172
0 1174 7 1 2 1112 1173
0 1175 7 1 2 1108 1174
0 1176 7 1 2 1106 1175
0 1177 7 1 2 1102 1176
0 1178 7 1 2 1100 1177
0 1179 7 1 2 1096 1178
0 1180 7 1 2 1094 1179
0 1181 7 1 2 2212 1180
0 1182 7 1 2 1090 1181
0 1183 7 1 2 2251 1182
0 1184 7 1 2 1020 1183
0 1185 5 1 1 1184
0 1186 7 1 2 2213 2249
0 1187 5 1 1 1186
0 1188 7 1 2 2200 1187
0 1189 5 1 1 1188
0 1190 7 1 2 2247 2202
0 1191 5 1 1 1190
0 1192 7 1 2 2245 2256
0 1193 5 1 1 1192
0 1194 7 1 2 2243 2254
0 1195 5 1 1 1194
0 1196 7 1 2 1193 1195
0 1197 5 1 1 1196
0 1198 7 1 2 2241 2259
0 1199 5 1 1 1198
0 1200 7 1 2 2239 2261
0 1201 5 1 1 1200
0 1202 7 1 2 2053 2266
0 1203 5 1 1 1202
0 1204 7 1 2 2237 2264
0 1205 5 1 1 1204
0 1206 7 1 2 2062 2270
0 1207 5 1 1 1206
0 1208 7 1 2 2235 2273
0 1209 5 1 1 1208
0 1210 7 1 2 2071 1209
0 1211 5 1 1 1210
0 1212 7 1 2 2233 2276
0 1213 5 1 1 1212
0 1214 7 1 2 2080 1213
0 1215 5 1 1 1214
0 1216 7 1 2 2231 2280
0 1217 5 1 1 1216
0 1218 7 1 2 2227 2283
0 1219 5 1 1 1218
0 1220 7 1 2 2229 2285
0 1221 5 1 1 1220
0 1222 7 1 2 2223 2287
0 1223 5 1 1 1222
0 1224 7 1 2 2106 2221
0 1225 5 1 1 1224
0 1226 7 1 2 2219 2293
0 1227 5 1 1 1226
0 1228 7 1 2 2123 2298
0 1229 5 1 1 1228
0 1230 7 1 2 2217 2296
0 1231 5 1 1 1230
0 1232 7 1 2 2302 1231
0 1233 7 1 2 1229 1232
0 1234 7 1 2 1227 1233
0 1235 7 1 2 1225 1234
0 1236 5 1 1 1235
0 1237 7 1 2 2225 2289
0 1238 5 1 1 1237
0 1239 7 1 2 1236 1238
0 1240 7 1 2 1223 1239
0 1241 7 1 2 1221 1240
0 1242 7 1 2 1219 1241
0 1243 5 1 1 1242
0 1244 7 1 2 1217 1243
0 1245 7 1 2 1215 1244
0 1246 7 1 2 1211 1245
0 1247 7 1 2 1207 1246
0 1248 7 1 2 1205 1247
0 1249 7 1 2 1203 1248
0 1250 7 1 2 1201 1249
0 1251 7 1 2 1199 1250
0 1252 7 1 2 1197 1251
0 1253 7 1 2 1191 1252
0 1254 7 1 2 1082 1253
0 1255 7 1 2 1189 1254
0 1256 5 1 1 1255
0 1257 7 1 2 1185 1256
3 4299 5 0 1 1257
