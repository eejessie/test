1 0 0 3 0
2 20 1 0
2 21 1 0
2 324 1 0
1 1 0 2 0
2 325 1 1
2 326 1 1
1 2 0 2 0
2 327 1 2
2 328 1 2
1 3 0 7 0
2 329 1 3
2 330 1 3
2 331 1 3
2 332 1 3
2 333 1 3
2 334 1 3
2 335 1 3
1 4 0 6 0
2 336 1 4
2 337 1 4
2 338 1 4
2 339 1 4
2 340 1 4
2 341 1 4
1 5 0 6 0
2 342 1 5
2 343 1 5
2 344 1 5
2 345 1 5
2 346 1 5
2 347 1 5
1 6 0 2 0
2 348 1 6
2 349 1 6
1 7 0 2 0
2 350 1 7
2 351 1 7
1 8 0 2 0
2 352 1 8
2 353 1 8
1 9 0 3 0
2 354 1 9
2 355 1 9
2 356 1 9
1 10 0 4 0
2 357 1 10
2 358 1 10
2 359 1 10
2 360 1 10
1 11 0 4 0
2 361 1 11
2 362 1 11
2 363 1 11
2 364 1 11
1 12 0 2 0
2 365 1 12
2 366 1 12
1 13 0 0 0
1 14 0 0 0
1 15 0 0 0
1 16 0 3 0
2 367 1 16
2 368 1 16
2 369 1 16
1 17 0 4 0
2 370 1 17
2 371 1 17
2 372 1 17
2 373 1 17
1 18 0 4 0
2 374 1 18
2 375 1 18
2 376 1 18
2 377 1 18
1 19 0 3 0
2 378 1 19
2 379 1 19
2 380 1 19
2 381 1 22
2 382 1 22
2 383 1 25
2 384 1 25
2 385 1 25
2 386 1 25
2 387 1 25
2 388 1 26
2 389 1 26
2 390 1 26
2 391 1 26
2 392 1 26
2 393 1 27
2 394 1 27
2 395 1 27
2 396 1 27
2 397 1 28
2 398 1 28
2 399 1 31
2 400 1 31
2 401 1 31
2 402 1 32
2 403 1 32
2 404 1 32
2 405 1 33
2 406 1 33
2 407 1 33
2 408 1 35
2 409 1 35
2 410 1 36
2 411 1 36
2 412 1 36
2 413 1 36
2 414 1 37
2 415 1 37
2 416 1 37
2 417 1 38
2 418 1 38
2 419 1 38
2 420 1 40
2 421 1 40
2 422 1 42
2 423 1 42
2 424 1 44
2 425 1 44
2 426 1 44
2 427 1 44
2 428 1 45
2 429 1 45
2 430 1 45
2 431 1 47
2 432 1 47
2 433 1 47
2 434 1 49
2 435 1 49
2 436 1 51
2 437 1 51
2 438 1 54
2 439 1 54
2 440 1 56
2 441 1 56
2 442 1 56
2 443 1 57
2 444 1 57
2 445 1 58
2 446 1 58
2 447 1 60
2 448 1 60
2 449 1 60
2 450 1 69
2 451 1 69
2 452 1 69
2 453 1 69
2 454 1 69
2 455 1 69
2 456 1 72
2 457 1 72
2 458 1 75
2 459 1 75
2 460 1 79
2 461 1 79
2 462 1 79
2 463 1 79
2 464 1 79
2 465 1 80
2 466 1 80
2 467 1 80
2 468 1 82
2 469 1 82
2 470 1 85
2 471 1 85
2 472 1 85
2 473 1 87
2 474 1 87
2 475 1 99
2 476 1 99
2 477 1 102
2 478 1 102
2 479 1 103
2 480 1 103
2 481 1 105
2 482 1 105
2 483 1 105
2 484 1 108
2 485 1 108
2 486 1 110
2 487 1 110
2 488 1 110
2 489 1 114
2 490 1 114
2 491 1 118
2 492 1 118
2 493 1 118
2 494 1 118
2 495 1 127
2 496 1 127
2 497 1 140
2 498 1 140
2 499 1 156
2 500 1 156
2 501 1 157
2 502 1 157
2 503 1 159
2 504 1 159
2 505 1 163
2 506 1 163
2 507 1 165
2 508 1 165
2 509 1 167
2 510 1 167
2 511 1 179
2 512 1 179
2 513 1 180
2 514 1 180
2 515 1 181
2 516 1 181
2 517 1 181
2 518 1 182
2 519 1 182
2 520 1 188
2 521 1 188
2 522 1 190
2 523 1 190
2 524 1 192
2 525 1 192
2 526 1 194
2 527 1 194
2 528 1 205
2 529 1 205
2 530 1 215
2 531 1 215
2 532 1 216
2 533 1 216
2 534 1 217
2 535 1 217
2 536 1 218
2 537 1 218
2 538 1 219
2 539 1 219
2 540 1 224
2 541 1 224
2 542 1 228
2 543 1 228
2 544 1 238
2 545 1 238
2 546 1 247
2 547 1 247
2 548 1 258
2 549 1 258
2 550 1 282
2 551 1 282
0 22 5 2 1 20
0 23 5 1 1 325
0 24 5 1 1 327
0 25 5 5 1 329
0 26 5 5 1 336
0 27 5 4 1 342
0 28 5 2 1 348
0 29 5 1 1 350
0 30 5 1 1 352
0 31 5 3 1 354
0 32 5 3 1 357
0 33 5 3 1 361
0 34 5 1 1 365
0 35 5 2 1 367
0 36 5 4 1 370
0 37 5 3 1 374
0 38 5 3 1 378
0 39 7 1 2 402 410
0 40 5 2 1 39
0 41 7 1 2 358 371
0 42 5 2 1 41
0 43 7 1 2 420 422
0 44 5 4 1 43
0 45 7 3 2 21 349
0 46 5 1 1 428
0 47 7 3 2 343 379
0 48 5 1 1 431
0 49 7 2 2 330 337
0 50 5 1 1 434
0 51 7 2 2 432 435
0 52 7 1 2 429 436
0 53 5 1 1 52
0 54 7 2 2 381 397
0 55 5 1 1 438
0 56 7 3 2 393 417
0 57 5 2 1 440
0 58 7 2 2 383 388
0 59 5 1 1 445
0 60 7 3 2 441 446
0 61 7 1 2 439 447
0 62 5 1 1 61
0 63 7 1 2 53 62
0 64 5 1 1 63
0 65 7 1 2 362 414
0 66 5 1 1 65
0 67 7 1 2 405 375
0 68 5 1 1 67
0 69 7 6 2 66 68
0 70 7 1 2 64 450
0 71 5 1 1 70
0 72 7 2 2 415 380
0 73 7 1 2 363 456
0 74 5 1 1 73
0 75 7 2 2 376 418
0 76 7 1 2 406 458
0 77 5 1 1 76
0 78 7 1 2 74 77
0 79 5 5 1 78
0 80 7 3 2 338 394
0 81 5 1 1 465
0 82 7 2 2 331 466
0 83 7 1 2 430 468
0 84 5 1 1 83
0 85 7 3 2 389 344
0 86 5 1 1 470
0 87 7 2 2 382 384
0 88 5 1 1 473
0 89 7 1 2 398 474
0 90 7 1 2 471 89
0 91 5 1 1 90
0 92 7 1 2 84 91
0 93 5 1 1 92
0 94 7 1 2 460 93
0 95 5 1 1 94
0 96 7 1 2 71 95
0 97 5 1 1 96
0 98 7 1 2 24 30
0 99 5 2 1 98
0 100 7 1 2 23 29
0 101 5 1 1 100
0 102 7 2 2 475 101
0 103 5 2 1 477
0 104 7 1 2 328 353
0 105 5 3 1 104
0 106 7 1 2 326 351
0 107 5 1 1 106
0 108 7 2 2 481 107
0 109 5 1 1 484
0 110 7 3 2 478 485
0 111 7 1 2 97 486
0 112 5 1 1 111
0 113 7 1 2 385 482
0 114 7 2 2 479 113
0 115 5 1 1 489
0 116 7 1 2 472 490
0 117 5 1 1 116
0 118 7 4 2 476 109
0 119 7 1 2 469 491
0 120 5 1 1 119
0 121 7 1 2 117 120
0 122 5 1 1 121
0 123 7 1 2 461 122
0 124 5 1 1 123
0 125 7 1 2 437 492
0 126 5 1 1 125
0 127 7 2 2 480 483
0 128 7 1 2 448 495
0 129 5 1 1 128
0 130 7 1 2 126 129
0 131 5 1 1 130
0 132 7 1 2 451 131
0 133 5 1 1 132
0 134 7 1 2 124 133
0 135 7 1 2 112 134
0 136 5 1 1 135
0 137 7 1 2 424 136
0 138 5 1 1 137
0 139 7 1 2 345 411
0 140 5 2 1 139
0 141 7 1 2 443 497
0 142 5 1 1 141
0 143 7 1 2 359 419
0 144 5 1 1 143
0 145 7 1 2 421 144
0 146 7 1 2 452 145
0 147 7 1 2 142 146
0 148 5 1 1 147
0 149 7 1 2 395 403
0 150 5 1 1 149
0 151 7 1 2 423 498
0 152 7 1 2 150 151
0 153 7 1 2 462 152
0 154 5 1 1 153
0 155 7 1 2 148 154
0 156 5 2 1 155
0 157 7 2 2 50 59
0 158 5 1 1 501
0 159 7 2 2 499 502
0 160 5 1 1 503
0 161 7 1 2 324 332
0 162 5 1 1 161
0 163 7 2 2 88 162
0 164 5 1 1 505
0 165 7 2 2 46 55
0 166 5 1 1 507
0 167 7 2 2 487 166
0 168 7 1 2 164 509
0 169 5 1 1 168
0 170 7 1 2 333 493
0 171 5 1 1 170
0 172 7 1 2 115 171
0 173 7 1 2 169 172
0 174 5 1 1 173
0 175 7 1 2 504 174
0 176 5 1 1 175
0 177 7 1 2 138 176
0 178 5 1 1 177
0 179 7 2 2 399 368
0 180 5 2 1 511
0 181 7 3 2 355 408
0 182 5 2 1 515
0 183 7 1 2 513 518
0 184 7 1 2 178 183
0 185 5 1 1 184
0 186 7 1 2 386 400
0 187 5 1 1 186
0 188 7 2 2 334 356
0 189 5 1 1 520
0 190 7 2 2 187 189
0 191 5 1 1 522
0 192 7 2 2 81 86
0 193 5 1 1 524
0 194 7 2 2 463 193
0 195 5 1 1 526
0 196 7 1 2 425 158
0 197 7 1 2 527 196
0 198 5 1 1 197
0 199 7 1 2 160 198
0 200 5 1 1 199
0 201 7 1 2 191 200
0 202 5 1 1 201
0 203 7 1 2 401 449
0 204 5 1 1 203
0 205 7 2 2 339 433
0 206 7 1 2 521 528
0 207 5 1 1 206
0 208 7 1 2 204 207
0 209 5 1 1 208
0 210 7 1 2 426 453
0 211 7 1 2 209 210
0 212 5 1 1 211
0 213 7 1 2 202 212
0 214 5 1 1 213
0 215 7 2 2 488 508
0 216 7 2 2 366 409
0 217 5 2 1 532
0 218 7 2 2 34 369
0 219 5 2 1 536
0 220 7 1 2 534 538
0 221 7 1 2 530 220
0 222 7 1 2 214 221
0 223 5 1 1 222
0 224 7 2 2 412 533
0 225 5 1 1 540
0 226 7 1 2 457 541
0 227 5 1 1 226
0 228 7 2 2 372 537
0 229 5 1 1 542
0 230 7 1 2 459 543
0 231 5 1 1 230
0 232 7 1 2 227 231
0 233 5 1 1 232
0 234 7 1 2 396 407
0 235 5 1 1 234
0 236 7 1 2 346 364
0 237 5 1 1 236
0 238 7 2 2 235 237
0 239 5 1 1 544
0 240 7 1 2 233 545
0 241 5 1 1 240
0 242 7 1 2 416 229
0 243 5 1 1 242
0 244 7 1 2 377 225
0 245 5 1 1 244
0 246 7 1 2 48 444
0 247 5 2 1 246
0 248 7 1 2 239 546
0 249 7 1 2 245 248
0 250 7 1 2 243 249
0 251 5 1 1 250
0 252 7 1 2 241 251
0 253 5 1 1 252
0 254 7 1 2 390 404
0 255 5 1 1 254
0 256 7 1 2 340 360
0 257 5 1 1 256
0 258 7 2 2 255 257
0 259 5 1 1 548
0 260 7 1 2 253 549
0 261 5 1 1 260
0 262 7 1 2 454 547
0 263 7 1 2 525 262
0 264 5 1 1 263
0 265 7 1 2 195 264
0 266 5 1 1 265
0 267 7 1 2 413 539
0 268 5 1 1 267
0 269 7 1 2 373 535
0 270 5 1 1 269
0 271 7 1 2 259 270
0 272 7 1 2 268 271
0 273 7 1 2 266 272
0 274 5 1 1 273
0 275 7 1 2 261 274
0 276 5 1 1 275
0 277 7 1 2 523 531
0 278 7 1 2 276 277
0 279 5 1 1 278
0 280 7 1 2 467 516
0 281 5 1 1 280
0 282 7 2 2 391 512
0 283 7 1 2 347 550
0 284 5 1 1 283
0 285 7 1 2 281 284
0 286 5 1 1 285
0 287 7 1 2 464 286
0 288 5 1 1 287
0 289 7 1 2 442 551
0 290 5 1 1 289
0 291 7 1 2 517 529
0 292 5 1 1 291
0 293 7 1 2 290 292
0 294 5 1 1 293
0 295 7 1 2 455 294
0 296 5 1 1 295
0 297 7 1 2 288 296
0 298 5 1 1 297
0 299 7 1 2 427 298
0 300 5 1 1 299
0 301 7 1 2 392 519
0 302 5 1 1 301
0 303 7 1 2 341 514
0 304 5 1 1 303
0 305 7 1 2 302 304
0 306 7 1 2 500 305
0 307 5 1 1 306
0 308 7 1 2 300 307
0 309 5 1 1 308
0 310 7 1 2 506 510
0 311 5 1 1 310
0 312 7 1 2 335 496
0 313 5 1 1 312
0 314 7 1 2 387 494
0 315 5 1 1 314
0 316 7 1 2 313 315
0 317 7 1 2 311 316
0 318 5 1 1 317
0 319 7 1 2 309 318
0 320 5 1 1 319
0 321 7 1 2 279 320
0 322 7 1 2 223 321
0 323 7 1 2 185 322
3 699 5 0 1 323
