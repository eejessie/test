1 0 0 2 0
2 49 1 0
2 1418 1 0
1 1 0 2 0
2 1419 1 1
2 1420 1 1
1 2 0 2 0
2 1421 1 2
2 1422 1 2
1 3 0 2 0
2 1423 1 3
2 1424 1 3
1 4 0 2 0
2 1425 1 4
2 1426 1 4
1 5 0 2 0
2 1427 1 5
2 1428 1 5
1 6 0 2 0
2 1429 1 6
2 1430 1 6
1 7 0 2 0
2 1431 1 7
2 1432 1 7
1 8 0 2 0
2 1433 1 8
2 1434 1 8
1 9 0 2 0
2 1435 1 9
2 1436 1 9
1 10 0 2 0
2 1437 1 10
2 1438 1 10
1 11 0 2 0
2 1439 1 11
2 1440 1 11
1 12 0 2 0
2 1441 1 12
2 1442 1 12
1 13 0 2 0
2 1443 1 13
2 1444 1 13
1 14 0 2 0
2 1445 1 14
2 1446 1 14
1 15 0 2 0
2 1447 1 15
2 1448 1 15
1 16 0 2 0
2 1449 1 16
2 1450 1 16
1 17 0 2 0
2 1451 1 17
2 1452 1 17
1 18 0 2 0
2 1453 1 18
2 1454 1 18
1 19 0 2 0
2 1455 1 19
2 1456 1 19
1 20 0 2 0
2 1457 1 20
2 1458 1 20
1 21 0 2 0
2 1459 1 21
2 1460 1 21
1 22 0 2 0
2 1461 1 22
2 1462 1 22
1 23 0 2 0
2 1463 1 23
2 1464 1 23
1 24 0 2 0
2 1465 1 24
2 1466 1 24
1 25 0 2 0
2 1467 1 25
2 1468 1 25
1 26 0 2 0
2 1469 1 26
2 1470 1 26
1 27 0 2 0
2 1471 1 27
2 1472 1 27
1 28 0 2 0
2 1473 1 28
2 1474 1 28
1 29 0 2 0
2 1475 1 29
2 1476 1 29
1 30 0 2 0
2 1477 1 30
2 1478 1 30
1 31 0 2 0
2 1479 1 31
2 1480 1 31
1 32 0 2 0
2 1481 1 32
2 1482 1 32
1 33 0 2 0
2 1483 1 33
2 1484 1 33
1 34 0 2 0
2 1485 1 34
2 1486 1 34
1 35 0 2 0
2 1487 1 35
2 1488 1 35
1 36 0 2 0
2 1489 1 36
2 1490 1 36
1 37 0 2 0
2 1491 1 37
2 1492 1 37
1 38 0 2 0
2 1493 1 38
2 1494 1 38
1 39 0 2 0
2 1495 1 39
2 1496 1 39
1 40 0 2 0
2 1497 1 40
2 1498 1 40
1 41 0 2 0
2 1499 1 41
2 1500 1 41
1 42 0 2 0
2 1501 1 42
2 1502 1 42
1 43 0 2 0
2 1503 1 43
2 1504 1 43
1 44 0 2 0
2 1505 1 44
2 1506 1 44
1 45 0 2 0
2 1507 1 45
2 1508 1 45
1 46 0 2 0
2 1509 1 46
2 1510 1 46
1 47 0 2 0
2 1511 1 47
2 1512 1 47
1 48 0 2 0
2 1513 1 48
2 1514 1 48
2 1515 1 68
2 1516 1 68
2 1517 1 69
2 1518 1 69
2 1519 1 70
2 1520 1 70
2 1521 1 71
2 1522 1 71
2 1523 1 72
2 1524 1 72
2 1525 1 73
2 1526 1 73
2 1527 1 74
2 1528 1 74
2 1529 1 75
2 1530 1 75
2 1531 1 76
2 1532 1 76
2 1533 1 77
2 1534 1 77
2 1535 1 78
2 1536 1 78
2 1537 1 79
2 1538 1 79
2 1539 1 80
2 1540 1 80
2 1541 1 83
2 1542 1 83
2 1543 1 100
2 1544 1 100
2 1545 1 102
2 1546 1 102
2 1547 1 104
2 1548 1 104
2 1549 1 105
2 1550 1 105
2 1551 1 106
2 1552 1 106
2 1553 1 106
2 1554 1 109
2 1555 1 109
2 1556 1 112
2 1557 1 112
2 1558 1 114
2 1559 1 114
2 1560 1 117
2 1561 1 117
2 1562 1 120
2 1563 1 120
2 1564 1 122
2 1565 1 122
2 1566 1 125
2 1567 1 125
2 1568 1 128
2 1569 1 128
2 1570 1 130
2 1571 1 130
2 1572 1 133
2 1573 1 133
2 1574 1 136
2 1575 1 136
2 1576 1 138
2 1577 1 138
2 1578 1 141
2 1579 1 141
2 1580 1 144
2 1581 1 144
2 1582 1 146
2 1583 1 146
2 1584 1 149
2 1585 1 149
2 1586 1 152
2 1587 1 152
2 1588 1 154
2 1589 1 154
2 1590 1 157
2 1591 1 157
2 1592 1 160
2 1593 1 160
2 1594 1 162
2 1595 1 162
2 1596 1 165
2 1597 1 165
2 1598 1 168
2 1599 1 168
2 1600 1 170
2 1601 1 170
2 1602 1 173
2 1603 1 173
2 1604 1 176
2 1605 1 176
2 1606 1 178
2 1607 1 178
2 1608 1 181
2 1609 1 181
2 1610 1 184
2 1611 1 184
2 1612 1 186
2 1613 1 186
2 1614 1 189
2 1615 1 189
2 1616 1 192
2 1617 1 192
2 1618 1 194
2 1619 1 194
2 1620 1 197
2 1621 1 197
2 1622 1 200
2 1623 1 200
2 1624 1 202
2 1625 1 202
2 1626 1 205
2 1627 1 205
2 1628 1 208
2 1629 1 208
2 1630 1 210
2 1631 1 210
2 1632 1 213
2 1633 1 213
2 1634 1 214
2 1635 1 214
2 1636 1 216
2 1637 1 216
2 1638 1 219
2 1639 1 219
2 1640 1 219
2 1641 1 219
2 1642 1 220
2 1643 1 220
2 1644 1 220
2 1645 1 221
2 1646 1 221
2 1647 1 227
2 1648 1 227
2 1649 1 227
2 1650 1 227
2 1651 1 230
2 1652 1 230
2 1653 1 230
2 1654 1 232
2 1655 1 232
2 1656 1 232
2 1657 1 233
2 1658 1 233
2 1659 1 233
2 1660 1 234
2 1661 1 234
2 1662 1 235
2 1663 1 235
2 1664 1 241
2 1665 1 241
2 1666 1 241
2 1667 1 241
2 1668 1 242
2 1669 1 242
2 1670 1 242
2 1671 1 244
2 1672 1 244
2 1673 1 244
2 1674 1 246
2 1675 1 246
2 1676 1 246
2 1677 1 247
2 1678 1 247
2 1679 1 253
2 1680 1 253
2 1681 1 253
2 1682 1 253
2 1683 1 254
2 1684 1 254
2 1685 1 254
2 1686 1 256
2 1687 1 256
2 1688 1 256
2 1689 1 258
2 1690 1 258
2 1691 1 258
2 1692 1 259
2 1693 1 259
2 1694 1 265
2 1695 1 265
2 1696 1 265
2 1697 1 265
2 1698 1 266
2 1699 1 266
2 1700 1 266
2 1701 1 268
2 1702 1 268
2 1703 1 268
2 1704 1 270
2 1705 1 270
2 1706 1 270
2 1707 1 271
2 1708 1 271
2 1709 1 277
2 1710 1 277
2 1711 1 277
2 1712 1 277
2 1713 1 278
2 1714 1 278
2 1715 1 278
2 1716 1 280
2 1717 1 280
2 1718 1 280
2 1719 1 282
2 1720 1 282
2 1721 1 282
2 1722 1 283
2 1723 1 283
2 1724 1 289
2 1725 1 289
2 1726 1 289
2 1727 1 289
2 1728 1 290
2 1729 1 290
2 1730 1 290
2 1731 1 292
2 1732 1 292
2 1733 1 292
2 1734 1 294
2 1735 1 294
2 1736 1 294
2 1737 1 295
2 1738 1 295
2 1739 1 301
2 1740 1 301
2 1741 1 302
2 1742 1 302
2 1743 1 302
2 1744 1 304
2 1745 1 304
2 1746 1 304
2 1747 1 306
2 1748 1 306
2 1749 1 306
2 1750 1 307
2 1751 1 307
2 1752 1 313
2 1753 1 313
2 1754 1 313
2 1755 1 313
2 1756 1 314
2 1757 1 314
2 1758 1 314
2 1759 1 316
2 1760 1 316
2 1761 1 316
2 1762 1 318
2 1763 1 318
2 1764 1 318
2 1765 1 319
2 1766 1 319
2 1767 1 325
2 1768 1 325
2 1769 1 326
2 1770 1 326
2 1771 1 326
2 1772 1 328
2 1773 1 328
2 1774 1 328
2 1775 1 330
2 1776 1 330
2 1777 1 330
2 1778 1 331
2 1779 1 331
2 1780 1 337
2 1781 1 337
2 1782 1 337
2 1783 1 337
2 1784 1 338
2 1785 1 338
2 1786 1 338
2 1787 1 340
2 1788 1 340
2 1789 1 340
2 1790 1 342
2 1791 1 342
2 1792 1 342
2 1793 1 343
2 1794 1 343
2 1795 1 349
2 1796 1 349
2 1797 1 349
2 1798 1 349
2 1799 1 350
2 1800 1 350
2 1801 1 350
2 1802 1 352
2 1803 1 352
2 1804 1 352
2 1805 1 354
2 1806 1 354
2 1807 1 354
2 1808 1 355
2 1809 1 355
2 1810 1 361
2 1811 1 361
2 1812 1 361
2 1813 1 361
2 1814 1 362
2 1815 1 362
2 1816 1 364
2 1817 1 364
2 1818 1 364
2 1819 1 366
2 1820 1 366
2 1821 1 366
2 1822 1 367
2 1823 1 367
2 1824 1 373
2 1825 1 373
2 1826 1 373
2 1827 1 376
2 1828 1 376
2 1829 1 376
2 1830 1 378
2 1831 1 378
2 1832 1 378
2 1833 1 381
2 1834 1 381
2 1835 1 383
2 1836 1 383
2 1837 1 383
2 1838 1 384
2 1839 1 384
2 1840 1 387
2 1841 1 387
2 1842 1 388
2 1843 1 388
2 1844 1 391
2 1845 1 391
2 1846 1 392
2 1847 1 392
2 1848 1 395
2 1849 1 395
2 1850 1 396
2 1851 1 396
2 1852 1 399
2 1853 1 399
2 1854 1 400
2 1855 1 400
2 1856 1 403
2 1857 1 403
2 1858 1 404
2 1859 1 404
2 1860 1 407
2 1861 1 407
2 1862 1 408
2 1863 1 408
2 1864 1 411
2 1865 1 411
2 1866 1 412
2 1867 1 412
2 1868 1 415
2 1869 1 415
2 1870 1 416
2 1871 1 416
2 1872 1 419
2 1873 1 419
2 1874 1 420
2 1875 1 420
2 1876 1 423
2 1877 1 423
2 1878 1 424
2 1879 1 424
2 1880 1 427
2 1881 1 427
2 1882 1 428
2 1883 1 428
2 1884 1 431
2 1885 1 431
2 1886 1 432
2 1887 1 432
2 1888 1 437
2 1889 1 437
2 1890 1 437
2 1891 1 438
2 1892 1 438
2 1893 1 439
2 1894 1 439
2 1895 1 445
2 1896 1 445
2 1897 1 445
2 1898 1 445
2 1899 1 446
2 1900 1 446
2 1901 1 446
2 1902 1 448
2 1903 1 448
2 1904 1 448
2 1905 1 449
2 1906 1 449
2 1907 1 450
2 1908 1 450
2 1909 1 450
2 1910 1 451
2 1911 1 451
2 1912 1 451
2 1913 1 452
2 1914 1 452
2 1915 1 453
2 1916 1 453
2 1917 1 459
2 1918 1 459
2 1919 1 459
2 1920 1 459
2 1921 1 460
2 1922 1 460
2 1923 1 460
2 1924 1 462
2 1925 1 462
2 1926 1 462
2 1927 1 464
2 1928 1 464
2 1929 1 464
2 1930 1 467
2 1931 1 467
2 1932 1 468
2 1933 1 468
2 1934 1 471
2 1935 1 471
2 1936 1 472
2 1937 1 472
2 1938 1 477
2 1939 1 477
2 1940 1 478
2 1941 1 478
2 1942 1 480
2 1943 1 480
2 1944 1 481
2 1945 1 481
2 1946 1 481
2 1947 1 482
2 1948 1 482
2 1949 1 487
2 1950 1 487
2 1951 1 487
2 1952 1 488
2 1953 1 488
2 1954 1 489
2 1955 1 489
2 1956 1 489
2 1957 1 490
2 1958 1 490
2 1959 1 495
2 1960 1 495
2 1961 1 495
2 1962 1 496
2 1963 1 496
2 1964 1 498
2 1965 1 498
2 1966 1 499
2 1967 1 499
2 1968 1 499
2 1969 1 500
2 1970 1 500
2 1971 1 505
2 1972 1 505
2 1973 1 505
2 1974 1 506
2 1975 1 506
2 1976 1 508
2 1977 1 508
2 1978 1 509
2 1979 1 509
2 1980 1 509
2 1981 1 510
2 1982 1 510
2 1983 1 515
2 1984 1 515
2 1985 1 515
2 1986 1 516
2 1987 1 516
2 1988 1 518
2 1989 1 518
2 1990 1 519
2 1991 1 519
2 1992 1 519
2 1993 1 520
2 1994 1 520
2 1995 1 525
2 1996 1 525
2 1997 1 525
2 1998 1 526
2 1999 1 526
2 2000 1 528
2 2001 1 528
2 2002 1 529
2 2003 1 529
2 2004 1 529
2 2005 1 530
2 2006 1 530
2 2007 1 535
2 2008 1 535
2 2009 1 535
2 2010 1 536
2 2011 1 536
2 2012 1 538
2 2013 1 538
2 2014 1 539
2 2015 1 539
2 2016 1 539
2 2017 1 540
2 2018 1 540
2 2019 1 545
2 2020 1 545
2 2021 1 545
2 2022 1 546
2 2023 1 546
2 2024 1 548
2 2025 1 548
2 2026 1 549
2 2027 1 549
2 2028 1 549
2 2029 1 550
2 2030 1 550
2 2031 1 555
2 2032 1 555
2 2033 1 555
2 2034 1 556
2 2035 1 556
2 2036 1 558
2 2037 1 558
2 2038 1 559
2 2039 1 559
2 2040 1 559
2 2041 1 560
2 2042 1 560
2 2043 1 565
2 2044 1 565
2 2045 1 565
2 2046 1 566
2 2047 1 566
2 2048 1 568
2 2049 1 568
2 2050 1 569
2 2051 1 569
2 2052 1 569
2 2053 1 570
2 2054 1 570
2 2055 1 575
2 2056 1 575
2 2057 1 575
2 2058 1 576
2 2059 1 576
2 2060 1 578
2 2061 1 578
2 2062 1 579
2 2063 1 579
2 2064 1 579
2 2065 1 580
2 2066 1 580
2 2067 1 585
2 2068 1 585
2 2069 1 585
2 2070 1 586
2 2071 1 586
2 2072 1 588
2 2073 1 588
2 2074 1 589
2 2075 1 589
2 2076 1 589
2 2077 1 590
2 2078 1 590
2 2079 1 595
2 2080 1 595
2 2081 1 595
2 2082 1 596
2 2083 1 596
2 2084 1 598
2 2085 1 598
2 2086 1 599
2 2087 1 599
2 2088 1 599
2 2089 1 600
2 2090 1 600
2 2091 1 605
2 2092 1 605
2 2093 1 606
2 2094 1 606
2 2095 1 608
2 2096 1 608
2 2097 1 609
2 2098 1 609
2 2099 1 609
2 2100 1 610
2 2101 1 610
2 2102 1 610
2 2103 1 610
2 2104 1 611
2 2105 1 611
2 2106 1 611
2 2107 1 612
2 2108 1 612
2 2109 1 613
2 2110 1 613
2 2111 1 614
2 2112 1 614
2 2113 1 617
2 2114 1 617
2 2115 1 620
2 2116 1 620
2 2117 1 621
2 2118 1 621
2 2119 1 625
2 2120 1 625
2 2121 1 628
2 2122 1 628
2 2123 1 629
2 2124 1 629
2 2125 1 633
2 2126 1 633
2 2127 1 636
2 2128 1 636
2 2129 1 637
2 2130 1 637
2 2131 1 641
2 2132 1 641
2 2133 1 644
2 2134 1 644
2 2135 1 645
2 2136 1 645
2 2137 1 649
2 2138 1 649
2 2139 1 652
2 2140 1 652
2 2141 1 653
2 2142 1 653
2 2143 1 657
2 2144 1 657
2 2145 1 660
2 2146 1 660
2 2147 1 661
2 2148 1 661
2 2149 1 665
2 2150 1 665
2 2151 1 668
2 2152 1 668
2 2153 1 669
2 2154 1 669
2 2155 1 673
2 2156 1 673
2 2157 1 676
2 2158 1 676
2 2159 1 677
2 2160 1 677
2 2161 1 681
2 2162 1 681
2 2163 1 684
2 2164 1 684
2 2165 1 685
2 2166 1 685
2 2167 1 689
2 2168 1 689
2 2169 1 692
2 2170 1 692
2 2171 1 693
2 2172 1 693
2 2173 1 697
2 2174 1 697
2 2175 1 700
2 2176 1 700
2 2177 1 701
2 2178 1 701
2 2179 1 705
2 2180 1 705
2 2181 1 708
2 2182 1 708
2 2183 1 709
2 2184 1 709
2 2185 1 713
2 2186 1 713
2 2187 1 716
2 2188 1 716
2 2189 1 717
2 2190 1 717
2 2191 1 720
2 2192 1 720
2 2193 1 720
2 2194 1 722
2 2195 1 722
2 2196 1 722
2 2197 1 723
2 2198 1 723
2 2199 1 723
2 2200 1 724
2 2201 1 724
2 2202 1 727
2 2203 1 727
2 2204 1 733
2 2205 1 733
2 2206 1 733
2 2207 1 739
2 2208 1 739
2 2209 1 742
2 2210 1 742
2 2211 1 745
2 2212 1 745
2 2213 1 751
2 2214 1 751
2 2215 1 759
2 2216 1 759
2 2217 1 767
2 2218 1 767
2 2219 1 775
2 2220 1 775
2 2221 1 781
2 2222 1 781
2 2223 1 789
2 2224 1 789
2 2225 1 793
2 2226 1 793
2 2227 1 801
2 2228 1 801
2 2229 1 805
2 2230 1 805
2 2231 1 813
2 2232 1 813
2 2233 1 829
2 2234 1 829
2 2235 1 844
2 2236 1 844
2 2237 1 856
2 2238 1 856
2 2239 1 877
2 2240 1 877
2 2241 1 888
2 2242 1 888
2 2243 1 896
2 2244 1 896
2 2245 1 904
2 2246 1 904
2 2247 1 936
2 2248 1 936
2 2249 1 936
2 2250 1 937
2 2251 1 937
2 2252 1 937
2 2253 1 940
2 2254 1 940
2 2255 1 941
2 2256 1 941
2 2257 1 944
2 2258 1 944
2 2259 1 945
2 2260 1 945
2 2261 1 948
2 2262 1 948
2 2263 1 949
2 2264 1 949
2 2265 1 952
2 2266 1 952
2 2267 1 953
2 2268 1 953
2 2269 1 956
2 2270 1 956
2 2271 1 957
2 2272 1 957
2 2273 1 960
2 2274 1 960
2 2275 1 961
2 2276 1 961
2 2277 1 964
2 2278 1 964
2 2279 1 965
2 2280 1 965
2 2281 1 968
2 2282 1 968
2 2283 1 969
2 2284 1 969
2 2285 1 972
2 2286 1 972
2 2287 1 973
2 2288 1 973
2 2289 1 976
2 2290 1 976
2 2291 1 977
2 2292 1 977
2 2293 1 980
2 2294 1 980
2 2295 1 981
2 2296 1 981
2 2297 1 984
2 2298 1 984
2 2299 1 985
2 2300 1 985
2 2301 1 988
2 2302 1 988
2 2303 1 989
2 2304 1 989
2 2305 1 992
2 2306 1 992
2 2307 1 993
2 2308 1 993
2 2309 1 996
2 2310 1 996
2 2311 1 997
2 2312 1 997
2 2313 1 1004
2 2314 1 1004
2 2315 1 1004
2 2316 1 1005
2 2317 1 1005
2 2318 1 1010
2 2319 1 1010
2 2320 1 1011
2 2321 1 1011
2 2322 1 1013
2 2323 1 1013
2 2324 1 1018
2 2325 1 1018
2 2326 1 1018
2 2327 1 1019
2 2328 1 1019
2 2329 1 1024
2 2330 1 1024
2 2331 1 1024
2 2332 1 1025
2 2333 1 1025
2 2334 1 1027
2 2335 1 1027
2 2336 1 1032
2 2337 1 1032
2 2338 1 1032
2 2339 1 1033
2 2340 1 1033
2 2341 1 1035
2 2342 1 1035
2 2343 1 1040
2 2344 1 1040
2 2345 1 1040
2 2346 1 1041
2 2347 1 1041
2 2348 1 1043
2 2349 1 1043
2 2350 1 1048
2 2351 1 1048
2 2352 1 1048
2 2353 1 1049
2 2354 1 1049
2 2355 1 1051
2 2356 1 1051
2 2357 1 1056
2 2358 1 1056
2 2359 1 1056
2 2360 1 1057
2 2361 1 1057
2 2362 1 1059
2 2363 1 1059
2 2364 1 1064
2 2365 1 1064
2 2366 1 1064
2 2367 1 1065
2 2368 1 1065
2 2369 1 1067
2 2370 1 1067
2 2371 1 1072
2 2372 1 1072
2 2373 1 1072
2 2374 1 1073
2 2375 1 1073
2 2376 1 1075
2 2377 1 1075
2 2378 1 1080
2 2379 1 1080
2 2380 1 1080
2 2381 1 1081
2 2382 1 1081
2 2383 1 1083
2 2384 1 1083
2 2385 1 1088
2 2386 1 1088
2 2387 1 1088
2 2388 1 1089
2 2389 1 1089
2 2390 1 1091
2 2391 1 1091
2 2392 1 1096
2 2393 1 1096
2 2394 1 1096
2 2395 1 1097
2 2396 1 1097
2 2397 1 1099
2 2398 1 1099
2 2399 1 1104
2 2400 1 1104
2 2401 1 1104
2 2402 1 1105
2 2403 1 1105
2 2404 1 1107
2 2405 1 1107
2 2406 1 1112
2 2407 1 1112
2 2408 1 1115
2 2409 1 1115
2 2410 1 1116
2 2411 1 1116
2 2412 1 1117
2 2413 1 1117
2 2414 1 1120
2 2415 1 1120
2 2416 1 1123
2 2417 1 1123
2 2418 1 1124
2 2419 1 1124
2 2420 1 1128
2 2421 1 1128
2 2422 1 1131
2 2423 1 1131
2 2424 1 1132
2 2425 1 1132
2 2426 1 1136
2 2427 1 1136
2 2428 1 1139
2 2429 1 1139
2 2430 1 1140
2 2431 1 1140
2 2432 1 1144
2 2433 1 1144
2 2434 1 1147
2 2435 1 1147
2 2436 1 1148
2 2437 1 1148
2 2438 1 1152
2 2439 1 1152
2 2440 1 1155
2 2441 1 1155
2 2442 1 1156
2 2443 1 1156
2 2444 1 1160
2 2445 1 1160
2 2446 1 1163
2 2447 1 1163
2 2448 1 1164
2 2449 1 1164
2 2450 1 1168
2 2451 1 1168
2 2452 1 1171
2 2453 1 1171
2 2454 1 1172
2 2455 1 1172
2 2456 1 1176
2 2457 1 1176
2 2458 1 1179
2 2459 1 1179
2 2460 1 1180
2 2461 1 1180
2 2462 1 1184
2 2463 1 1184
2 2464 1 1187
2 2465 1 1187
2 2466 1 1188
2 2467 1 1188
2 2468 1 1192
2 2469 1 1192
2 2470 1 1195
2 2471 1 1195
2 2472 1 1196
2 2473 1 1196
2 2474 1 1200
2 2475 1 1200
2 2476 1 1203
2 2477 1 1203
2 2478 1 1204
2 2479 1 1204
2 2480 1 1208
2 2481 1 1208
2 2482 1 1211
2 2483 1 1211
2 2484 1 1212
2 2485 1 1212
2 2486 1 1216
2 2487 1 1216
2 2488 1 1219
2 2489 1 1219
2 2490 1 1220
2 2491 1 1220
2 2492 1 1226
2 2493 1 1226
2 2494 1 1227
2 2495 1 1227
2 2496 1 1232
2 2497 1 1232
2 2498 1 1235
2 2499 1 1235
2 2500 1 1238
2 2501 1 1238
2 2502 1 1244
2 2503 1 1244
2 2504 1 1252
2 2505 1 1252
2 2506 1 1260
2 2507 1 1260
2 2508 1 1268
2 2509 1 1268
2 2510 1 1274
2 2511 1 1274
2 2512 1 1282
2 2513 1 1282
2 2514 1 1286
2 2515 1 1286
2 2516 1 1294
2 2517 1 1294
2 2518 1 1298
2 2519 1 1298
2 2520 1 1306
2 2521 1 1306
2 2522 1 1314
2 2523 1 1314
2 2524 1 1329
2 2525 1 1329
2 2526 1 1341
2 2527 1 1341
2 2528 1 1362
2 2529 1 1362
2 2530 1 1373
2 2531 1 1373
2 2532 1 1381
2 2533 1 1381
2 2534 1 1389
2 2535 1 1389
0 50 5 1 1 49
0 51 5 1 1 1419
0 52 5 1 1 1421
0 53 5 1 1 1423
0 54 5 1 1 1425
0 55 5 1 1 1427
0 56 5 1 1 1429
0 57 5 1 1 1431
0 58 5 1 1 1433
0 59 5 1 1 1435
0 60 5 1 1 1437
0 61 5 1 1 1439
0 62 5 1 1 1441
0 63 5 1 1 1443
0 64 5 1 1 1445
0 65 5 1 1 1447
0 66 5 1 1 1449
0 67 5 1 1 1451
0 68 5 2 1 1453
0 69 5 2 1 1455
0 70 5 2 1 1457
0 71 5 2 1 1459
0 72 5 2 1 1461
0 73 5 2 1 1463
0 74 5 2 1 1465
0 75 5 2 1 1467
0 76 5 2 1 1469
0 77 5 2 1 1471
0 78 5 2 1 1473
0 79 5 2 1 1475
0 80 5 2 1 1477
0 81 5 1 1 1479
0 82 5 1 1 1481
0 83 5 2 1 1483
0 84 5 1 1 1485
0 85 5 1 1 1487
0 86 5 1 1 1489
0 87 5 1 1 1491
0 88 5 1 1 1493
0 89 5 1 1 1495
0 90 5 1 1 1497
0 91 5 1 1 1499
0 92 5 1 1 1501
0 93 5 1 1 1503
0 94 5 1 1 1505
0 95 5 1 1 1507
0 96 5 1 1 1509
0 97 5 1 1 1511
0 98 5 1 1 1513
0 99 7 1 2 65 81
0 100 5 2 1 99
0 101 7 1 2 51 67
0 102 5 2 1 101
0 103 7 1 2 1420 1452
0 104 5 2 1 103
0 105 7 2 2 1418 1450
0 106 5 3 1 1549
0 107 7 1 2 1547 1551
0 108 5 1 1 107
0 109 7 2 2 1545 108
0 110 5 1 1 1554
0 111 7 1 2 52 110
0 112 5 2 1 111
0 113 7 1 2 1422 1555
0 114 5 2 1 113
0 115 7 1 2 1515 1558
0 116 5 1 1 115
0 117 7 2 2 1556 116
0 118 5 1 1 1560
0 119 7 1 2 53 118
0 120 5 2 1 119
0 121 7 1 2 1424 1561
0 122 5 2 1 121
0 123 7 1 2 1517 1564
0 124 5 1 1 123
0 125 7 2 2 1562 124
0 126 5 1 1 1566
0 127 7 1 2 54 126
0 128 5 2 1 127
0 129 7 1 2 1426 1567
0 130 5 2 1 129
0 131 7 1 2 1519 1570
0 132 5 1 1 131
0 133 7 2 2 1568 132
0 134 5 1 1 1572
0 135 7 1 2 55 134
0 136 5 2 1 135
0 137 7 1 2 1428 1573
0 138 5 2 1 137
0 139 7 1 2 1521 1576
0 140 5 1 1 139
0 141 7 2 2 1574 140
0 142 5 1 1 1578
0 143 7 1 2 56 142
0 144 5 2 1 143
0 145 7 1 2 1430 1579
0 146 5 2 1 145
0 147 7 1 2 1523 1582
0 148 5 1 1 147
0 149 7 2 2 1580 148
0 150 5 1 1 1584
0 151 7 1 2 57 150
0 152 5 2 1 151
0 153 7 1 2 1432 1585
0 154 5 2 1 153
0 155 7 1 2 1525 1588
0 156 5 1 1 155
0 157 7 2 2 1586 156
0 158 5 1 1 1590
0 159 7 1 2 58 158
0 160 5 2 1 159
0 161 7 1 2 1434 1591
0 162 5 2 1 161
0 163 7 1 2 1527 1594
0 164 5 1 1 163
0 165 7 2 2 1592 164
0 166 5 1 1 1596
0 167 7 1 2 59 166
0 168 5 2 1 167
0 169 7 1 2 1436 1597
0 170 5 2 1 169
0 171 7 1 2 1529 1600
0 172 5 1 1 171
0 173 7 2 2 1598 172
0 174 5 1 1 1602
0 175 7 1 2 60 174
0 176 5 2 1 175
0 177 7 1 2 1438 1603
0 178 5 2 1 177
0 179 7 1 2 1531 1606
0 180 5 1 1 179
0 181 7 2 2 1604 180
0 182 5 1 1 1608
0 183 7 1 2 61 182
0 184 5 2 1 183
0 185 7 1 2 1440 1609
0 186 5 2 1 185
0 187 7 1 2 1533 1612
0 188 5 1 1 187
0 189 7 2 2 1610 188
0 190 5 1 1 1614
0 191 7 1 2 62 190
0 192 5 2 1 191
0 193 7 1 2 1442 1615
0 194 5 2 1 193
0 195 7 1 2 1535 1618
0 196 5 1 1 195
0 197 7 2 2 1616 196
0 198 5 1 1 1620
0 199 7 1 2 63 198
0 200 5 2 1 199
0 201 7 1 2 1444 1621
0 202 5 2 1 201
0 203 7 1 2 1537 1624
0 204 5 1 1 203
0 205 7 2 2 1622 204
0 206 5 1 1 1626
0 207 7 1 2 64 206
0 208 5 2 1 207
0 209 7 1 2 1446 1627
0 210 5 2 1 209
0 211 7 1 2 1539 1630
0 212 5 1 1 211
0 213 7 2 2 1628 212
0 214 5 2 1 1632
0 215 7 1 2 1448 1480
0 216 5 2 1 215
0 217 7 1 2 1634 1636
0 218 5 1 1 217
0 219 7 4 2 1543 218
0 220 5 3 1 1638
0 221 7 2 2 1623 1625
0 222 5 1 1 1645
0 223 7 1 2 1476 1646
0 224 5 1 1 223
0 225 7 1 2 1538 222
0 226 5 1 1 225
0 227 7 4 2 224 226
0 228 5 1 1 1647
0 229 7 1 2 1508 228
0 230 5 3 1 229
0 231 7 1 2 95 1648
0 232 5 3 1 231
0 233 7 3 2 1651 1654
0 234 5 2 1 1657
0 235 7 2 2 1617 1619
0 236 5 1 1 1662
0 237 7 1 2 1474 1663
0 238 5 1 1 237
0 239 7 1 2 1536 236
0 240 5 1 1 239
0 241 7 4 2 238 240
0 242 5 3 1 1664
0 243 7 1 2 94 1665
0 244 5 3 1 243
0 245 7 1 2 1506 1668
0 246 5 3 1 245
0 247 7 2 2 1611 1613
0 248 5 1 1 1677
0 249 7 1 2 1472 1678
0 250 5 1 1 249
0 251 7 1 2 1534 248
0 252 5 1 1 251
0 253 7 4 2 250 252
0 254 5 3 1 1679
0 255 7 1 2 93 1680
0 256 5 3 1 255
0 257 7 1 2 1504 1683
0 258 5 3 1 257
0 259 7 2 2 1605 1607
0 260 5 1 1 1692
0 261 7 1 2 1470 1693
0 262 5 1 1 261
0 263 7 1 2 1532 260
0 264 5 1 1 263
0 265 7 4 2 262 264
0 266 5 3 1 1694
0 267 7 1 2 92 1695
0 268 5 3 1 267
0 269 7 1 2 1502 1698
0 270 5 3 1 269
0 271 7 2 2 1599 1601
0 272 5 1 1 1707
0 273 7 1 2 1468 1708
0 274 5 1 1 273
0 275 7 1 2 1530 272
0 276 5 1 1 275
0 277 7 4 2 274 276
0 278 5 3 1 1709
0 279 7 1 2 91 1710
0 280 5 3 1 279
0 281 7 1 2 1500 1713
0 282 5 3 1 281
0 283 7 2 2 1593 1595
0 284 5 1 1 1722
0 285 7 1 2 1466 1723
0 286 5 1 1 285
0 287 7 1 2 1528 284
0 288 5 1 1 287
0 289 7 4 2 286 288
0 290 5 3 1 1724
0 291 7 1 2 90 1725
0 292 5 3 1 291
0 293 7 1 2 1498 1728
0 294 5 3 1 293
0 295 7 2 2 1587 1589
0 296 5 1 1 1737
0 297 7 1 2 1464 1738
0 298 5 1 1 297
0 299 7 1 2 1526 296
0 300 5 1 1 299
0 301 7 2 2 298 300
0 302 5 3 1 1739
0 303 7 1 2 89 1740
0 304 5 3 1 303
0 305 7 1 2 1496 1741
0 306 5 3 1 305
0 307 7 2 2 1581 1583
0 308 5 1 1 1750
0 309 7 1 2 1462 1751
0 310 5 1 1 309
0 311 7 1 2 1524 308
0 312 5 1 1 311
0 313 7 4 2 310 312
0 314 5 3 1 1752
0 315 7 1 2 88 1753
0 316 5 3 1 315
0 317 7 1 2 1494 1756
0 318 5 3 1 317
0 319 7 2 2 1575 1577
0 320 5 1 1 1765
0 321 7 1 2 1460 1766
0 322 5 1 1 321
0 323 7 1 2 1522 320
0 324 5 1 1 323
0 325 7 2 2 322 324
0 326 5 3 1 1767
0 327 7 1 2 87 1768
0 328 5 3 1 327
0 329 7 1 2 1492 1769
0 330 5 3 1 329
0 331 7 2 2 1569 1571
0 332 5 1 1 1778
0 333 7 1 2 1458 1779
0 334 5 1 1 333
0 335 7 1 2 1520 332
0 336 5 1 1 335
0 337 7 4 2 334 336
0 338 5 3 1 1780
0 339 7 1 2 86 1781
0 340 5 3 1 339
0 341 7 1 2 1490 1784
0 342 5 3 1 341
0 343 7 2 2 1563 1565
0 344 5 1 1 1793
0 345 7 1 2 1456 1794
0 346 5 1 1 345
0 347 7 1 2 1518 344
0 348 5 1 1 347
0 349 7 4 2 346 348
0 350 5 3 1 1795
0 351 7 1 2 85 1796
0 352 5 3 1 351
0 353 7 1 2 1488 1799
0 354 5 3 1 353
0 355 7 2 2 1557 1559
0 356 5 1 1 1808
0 357 7 1 2 1454 1809
0 358 5 1 1 357
0 359 7 1 2 1516 356
0 360 5 1 1 359
0 361 7 4 2 358 360
0 362 5 2 1 1810
0 363 7 1 2 84 1811
0 364 5 3 1 363
0 365 7 1 2 1486 1814
0 366 5 3 1 365
0 367 7 2 2 1546 1548
0 368 5 1 1 1822
0 369 7 1 2 1550 368
0 370 5 1 1 369
0 371 7 1 2 1552 1823
0 372 5 1 1 371
0 373 7 3 2 370 372
0 374 5 1 1 1824
0 375 7 1 2 1541 374
0 376 5 3 1 375
0 377 7 1 2 1484 1825
0 378 5 3 1 377
0 379 7 1 2 50 66
0 380 5 1 1 379
0 381 7 2 2 1553 380
0 382 5 1 1 1833
0 383 7 3 2 82 1834
0 384 5 2 1 1835
0 385 7 1 2 1830 1836
0 386 5 1 1 385
0 387 7 2 2 1827 386
0 388 5 2 1 1840
0 389 7 1 2 1819 1842
0 390 5 1 1 389
0 391 7 2 2 1816 390
0 392 5 2 1 1844
0 393 7 1 2 1805 1846
0 394 5 1 1 393
0 395 7 2 2 1802 394
0 396 5 2 1 1848
0 397 7 1 2 1790 1850
0 398 5 1 1 397
0 399 7 2 2 1787 398
0 400 5 2 1 1852
0 401 7 1 2 1775 1854
0 402 5 1 1 401
0 403 7 2 2 1772 402
0 404 5 2 1 1856
0 405 7 1 2 1762 1858
0 406 5 1 1 405
0 407 7 2 2 1759 406
0 408 5 2 1 1860
0 409 7 1 2 1747 1862
0 410 5 1 1 409
0 411 7 2 2 1744 410
0 412 5 2 1 1864
0 413 7 1 2 1734 1866
0 414 5 1 1 413
0 415 7 2 2 1731 414
0 416 5 2 1 1868
0 417 7 1 2 1719 1870
0 418 5 1 1 417
0 419 7 2 2 1716 418
0 420 5 2 1 1872
0 421 7 1 2 1704 1874
0 422 5 1 1 421
0 423 7 2 2 1701 422
0 424 5 2 1 1876
0 425 7 1 2 1689 1878
0 426 5 1 1 425
0 427 7 2 2 1686 426
0 428 5 2 1 1880
0 429 7 1 2 1674 1882
0 430 5 1 1 429
0 431 7 2 2 1671 430
0 432 5 2 1 1884
0 433 7 1 2 1658 1885
0 434 5 1 1 433
0 435 7 1 2 1660 1886
0 436 5 1 1 435
0 437 7 3 2 434 436
0 438 5 2 1 1888
0 439 7 2 2 1544 1637
0 440 5 1 1 1893
0 441 7 1 2 1633 440
0 442 5 1 1 441
0 443 7 1 2 1635 1894
0 444 5 1 1 443
0 445 7 4 2 442 444
0 446 5 3 1 1895
0 447 7 1 2 1512 1896
0 448 5 3 1 447
0 449 7 2 2 97 1899
0 450 5 3 1 1905
0 451 7 3 2 1902 1907
0 452 5 2 1 1910
0 453 7 2 2 1629 1631
0 454 5 1 1 1915
0 455 7 1 2 1478 454
0 456 5 1 1 455
0 457 7 1 2 1540 1916
0 458 5 1 1 457
0 459 7 4 2 456 458
0 460 5 3 1 1917
0 461 7 1 2 96 1921
0 462 5 3 1 461
0 463 7 1 2 1510 1918
0 464 5 3 1 463
0 465 7 1 2 1652 1887
0 466 5 1 1 465
0 467 7 2 2 1655 466
0 468 5 2 1 1930
0 469 7 1 2 1927 1932
0 470 5 1 1 469
0 471 7 2 2 1924 470
0 472 5 2 1 1934
0 473 7 1 2 1911 1935
0 474 5 1 1 473
0 475 7 1 2 1913 1936
0 476 5 1 1 475
0 477 7 2 2 474 476
0 478 5 2 1 1938
0 479 7 1 2 1889 1939
0 480 5 2 1 479
0 481 7 3 2 1672 1675
0 482 5 2 1 1944
0 483 7 1 2 1881 1947
0 484 5 1 1 483
0 485 7 1 2 1883 1945
0 486 5 1 1 485
0 487 7 3 2 484 486
0 488 5 2 1 1949
0 489 7 3 2 1925 1928
0 490 5 2 1 1954
0 491 7 1 2 1931 1955
0 492 5 1 1 491
0 493 7 1 2 1933 1957
0 494 5 1 1 493
0 495 7 3 2 492 494
0 496 5 2 1 1959
0 497 7 1 2 1952 1960
0 498 5 2 1 497
0 499 7 3 2 1687 1690
0 500 5 2 1 1966
0 501 7 1 2 1877 1969
0 502 5 1 1 501
0 503 7 1 2 1879 1967
0 504 5 1 1 503
0 505 7 3 2 502 504
0 506 5 2 1 1971
0 507 7 1 2 1890 1974
0 508 5 2 1 507
0 509 7 3 2 1702 1705
0 510 5 2 1 1978
0 511 7 1 2 1873 1981
0 512 5 1 1 511
0 513 7 1 2 1875 1979
0 514 5 1 1 513
0 515 7 3 2 512 514
0 516 5 2 1 1983
0 517 7 1 2 1953 1986
0 518 5 2 1 517
0 519 7 3 2 1717 1720
0 520 5 2 1 1990
0 521 7 1 2 1869 1993
0 522 5 1 1 521
0 523 7 1 2 1871 1991
0 524 5 1 1 523
0 525 7 3 2 522 524
0 526 5 2 1 1995
0 527 7 1 2 1975 1998
0 528 5 2 1 527
0 529 7 3 2 1732 1735
0 530 5 2 1 2002
0 531 7 1 2 1865 2005
0 532 5 1 1 531
0 533 7 1 2 1867 2003
0 534 5 1 1 533
0 535 7 3 2 532 534
0 536 5 2 1 2007
0 537 7 1 2 1987 2010
0 538 5 2 1 537
0 539 7 3 2 1745 1748
0 540 5 2 1 2014
0 541 7 1 2 1861 2017
0 542 5 1 1 541
0 543 7 1 2 1863 2015
0 544 5 1 1 543
0 545 7 3 2 542 544
0 546 5 2 1 2019
0 547 7 1 2 1999 2022
0 548 5 2 1 547
0 549 7 3 2 1760 1763
0 550 5 2 1 2026
0 551 7 1 2 1857 2029
0 552 5 1 1 551
0 553 7 1 2 1859 2027
0 554 5 1 1 553
0 555 7 3 2 552 554
0 556 5 2 1 2031
0 557 7 1 2 2011 2034
0 558 5 2 1 557
0 559 7 3 2 1773 1776
0 560 5 2 1 2038
0 561 7 1 2 1853 2041
0 562 5 1 1 561
0 563 7 1 2 1855 2039
0 564 5 1 1 563
0 565 7 3 2 562 564
0 566 5 2 1 2043
0 567 7 1 2 2023 2046
0 568 5 2 1 567
0 569 7 3 2 1788 1791
0 570 5 2 1 2050
0 571 7 1 2 1849 2053
0 572 5 1 1 571
0 573 7 1 2 1851 2051
0 574 5 1 1 573
0 575 7 3 2 572 574
0 576 5 2 1 2055
0 577 7 1 2 2035 2058
0 578 5 2 1 577
0 579 7 3 2 1803 1806
0 580 5 2 1 2062
0 581 7 1 2 1845 2065
0 582 5 1 1 581
0 583 7 1 2 1847 2063
0 584 5 1 1 583
0 585 7 3 2 582 584
0 586 5 2 1 2067
0 587 7 1 2 2047 2070
0 588 5 2 1 587
0 589 7 3 2 1817 1820
0 590 5 2 1 2074
0 591 7 1 2 1841 2077
0 592 5 1 1 591
0 593 7 1 2 1843 2075
0 594 5 1 1 593
0 595 7 3 2 592 594
0 596 5 2 1 2079
0 597 7 1 2 2059 2082
0 598 5 2 1 597
0 599 7 3 2 1828 1831
0 600 5 2 1 2086
0 601 7 1 2 1838 2087
0 602 5 1 1 601
0 603 7 1 2 1837 2089
0 604 5 1 1 603
0 605 7 2 2 602 604
0 606 5 2 1 2091
0 607 7 1 2 2071 2092
0 608 5 2 1 607
0 609 7 3 2 1482 382
0 610 5 4 1 2097
0 611 7 3 2 1839 2100
0 612 5 2 1 2104
0 613 7 2 2 2083 2107
0 614 5 2 1 2109
0 615 7 1 2 2068 2093
0 616 5 1 1 615
0 617 7 2 2 2095 616
0 618 5 1 1 2113
0 619 7 1 2 2110 2114
0 620 5 2 1 619
0 621 7 2 2 2096 2115
0 622 5 1 1 2117
0 623 7 1 2 2056 2080
0 624 5 1 1 623
0 625 7 2 2 2084 624
0 626 5 1 1 2119
0 627 7 1 2 622 2120
0 628 5 2 1 627
0 629 7 2 2 2085 2121
0 630 5 1 1 2123
0 631 7 1 2 2044 2069
0 632 5 1 1 631
0 633 7 2 2 2072 632
0 634 5 1 1 2125
0 635 7 1 2 630 2126
0 636 5 2 1 635
0 637 7 2 2 2073 2127
0 638 5 1 1 2129
0 639 7 1 2 2032 2057
0 640 5 1 1 639
0 641 7 2 2 2060 640
0 642 5 1 1 2131
0 643 7 1 2 638 2132
0 644 5 2 1 643
0 645 7 2 2 2061 2133
0 646 5 1 1 2135
0 647 7 1 2 2020 2045
0 648 5 1 1 647
0 649 7 2 2 2048 648
0 650 5 1 1 2137
0 651 7 1 2 646 2138
0 652 5 2 1 651
0 653 7 2 2 2049 2139
0 654 5 1 1 2141
0 655 7 1 2 2008 2033
0 656 5 1 1 655
0 657 7 2 2 2036 656
0 658 5 1 1 2143
0 659 7 1 2 654 2144
0 660 5 2 1 659
0 661 7 2 2 2037 2145
0 662 5 1 1 2147
0 663 7 1 2 1996 2021
0 664 5 1 1 663
0 665 7 2 2 2024 664
0 666 5 1 1 2149
0 667 7 1 2 662 2150
0 668 5 2 1 667
0 669 7 2 2 2025 2151
0 670 5 1 1 2153
0 671 7 1 2 1984 2009
0 672 5 1 1 671
0 673 7 2 2 2012 672
0 674 5 1 1 2155
0 675 7 1 2 670 2156
0 676 5 2 1 675
0 677 7 2 2 2013 2157
0 678 5 1 1 2159
0 679 7 1 2 1972 1997
0 680 5 1 1 679
0 681 7 2 2 2000 680
0 682 5 1 1 2161
0 683 7 1 2 678 2162
0 684 5 2 1 683
0 685 7 2 2 2001 2163
0 686 5 1 1 2165
0 687 7 1 2 1950 1985
0 688 5 1 1 687
0 689 7 2 2 1988 688
0 690 5 1 1 2167
0 691 7 1 2 686 2168
0 692 5 2 1 691
0 693 7 2 2 1989 2169
0 694 5 1 1 2171
0 695 7 1 2 1891 1973
0 696 5 1 1 695
0 697 7 2 2 1976 696
0 698 5 1 1 2173
0 699 7 1 2 694 2174
0 700 5 2 1 699
0 701 7 2 2 1977 2175
0 702 5 1 1 2177
0 703 7 1 2 1951 1962
0 704 5 1 1 703
0 705 7 2 2 1964 704
0 706 5 1 1 2179
0 707 7 1 2 702 2180
0 708 5 2 1 707
0 709 7 2 2 1965 2181
0 710 5 1 1 2183
0 711 7 1 2 1892 1940
0 712 5 1 1 711
0 713 7 2 2 1942 712
0 714 5 1 1 2185
0 715 7 1 2 710 2186
0 716 5 2 1 715
0 717 7 2 2 1943 2187
0 718 5 1 1 2189
0 719 7 1 2 1514 1642
0 720 5 3 1 719
0 721 7 1 2 98 1639
0 722 5 3 1 721
0 723 7 3 2 2191 2194
0 724 5 2 1 2197
0 725 7 1 2 1903 1937
0 726 5 1 1 725
0 727 7 2 2 1908 726
0 728 5 1 1 2202
0 729 7 1 2 2198 728
0 730 5 1 1 729
0 731 7 1 2 2200 2203
0 732 5 1 1 731
0 733 7 3 2 730 732
0 734 5 1 1 2204
0 735 7 1 2 1961 2205
0 736 5 1 1 735
0 737 7 1 2 1963 734
0 738 5 1 1 737
0 739 7 2 2 736 738
0 740 5 1 1 2207
0 741 7 1 2 718 740
0 742 5 2 1 741
0 743 7 1 2 2190 2208
0 744 5 1 1 743
0 745 7 2 2 2209 744
0 746 5 1 1 2211
0 747 7 1 2 1640 746
0 748 5 1 1 747
0 749 7 1 2 2184 714
0 750 5 1 1 749
0 751 7 2 2 2188 750
0 752 5 1 1 2213
0 753 7 1 2 1897 2214
0 754 5 1 1 753
0 755 7 1 2 1900 752
0 756 5 1 1 755
0 757 7 1 2 2172 698
0 758 5 1 1 757
0 759 7 2 2 2176 758
0 760 5 1 1 2215
0 761 7 1 2 2166 690
0 762 5 1 1 761
0 763 7 1 2 2170 762
0 764 5 1 1 763
0 765 7 1 2 2154 674
0 766 5 1 1 765
0 767 7 2 2 2158 766
0 768 5 1 1 2217
0 769 7 1 2 1696 768
0 770 5 1 1 769
0 771 7 1 2 1699 2218
0 772 5 1 1 771
0 773 7 1 2 2148 666
0 774 5 1 1 773
0 775 7 2 2 2152 774
0 776 5 1 1 2219
0 777 7 1 2 1714 2220
0 778 5 1 1 777
0 779 7 1 2 2142 658
0 780 5 1 1 779
0 781 7 2 2 2146 780
0 782 5 1 1 2221
0 783 7 1 2 1729 2222
0 784 5 1 1 783
0 785 7 1 2 1726 782
0 786 5 1 1 785
0 787 7 1 2 2136 650
0 788 5 1 1 787
0 789 7 2 2 2140 788
0 790 5 1 1 2223
0 791 7 1 2 2130 642
0 792 5 1 1 791
0 793 7 2 2 2134 792
0 794 5 1 1 2225
0 795 7 1 2 1757 2226
0 796 5 1 1 795
0 797 7 1 2 1754 794
0 798 5 1 1 797
0 799 7 1 2 2124 634
0 800 5 1 1 799
0 801 7 2 2 2128 800
0 802 5 1 1 2227
0 803 7 1 2 2118 626
0 804 5 1 1 803
0 805 7 2 2 2122 804
0 806 5 1 1 2229
0 807 7 1 2 1785 2230
0 808 5 1 1 807
0 809 7 1 2 1782 806
0 810 5 1 1 809
0 811 7 1 2 2081 2105
0 812 5 1 1 811
0 813 7 2 2 2111 812
0 814 5 1 1 2231
0 815 7 1 2 1815 2232
0 816 5 1 1 815
0 817 7 1 2 1812 814
0 818 5 1 1 817
0 819 7 1 2 1542 2098
0 820 5 1 1 819
0 821 7 1 2 2094 2101
0 822 5 1 1 821
0 823 7 1 2 1826 822
0 824 5 1 1 823
0 825 7 1 2 820 824
0 826 5 1 1 825
0 827 7 1 2 818 826
0 828 5 1 1 827
0 829 7 2 2 816 828
0 830 5 1 1 2233
0 831 7 1 2 1797 2234
0 832 5 1 1 831
0 833 7 1 2 2112 618
0 834 5 1 1 833
0 835 7 1 2 2116 834
0 836 7 1 2 832 835
0 837 5 1 1 836
0 838 7 1 2 1800 830
0 839 5 1 1 838
0 840 7 1 2 837 839
0 841 5 1 1 840
0 842 7 1 2 810 841
0 843 5 1 1 842
0 844 7 2 2 808 843
0 845 5 1 1 2235
0 846 7 1 2 2228 845
0 847 5 1 1 846
0 848 7 1 2 802 2236
0 849 5 1 1 848
0 850 7 1 2 1770 849
0 851 5 1 1 850
0 852 7 1 2 847 851
0 853 5 1 1 852
0 854 7 1 2 798 853
0 855 5 1 1 854
0 856 7 2 2 796 855
0 857 5 1 1 2237
0 858 7 1 2 2224 857
0 859 5 1 1 858
0 860 7 1 2 790 2238
0 861 5 1 1 860
0 862 7 1 2 1742 861
0 863 5 1 1 862
0 864 7 1 2 859 863
0 865 5 1 1 864
0 866 7 1 2 786 865
0 867 5 1 1 866
0 868 7 1 2 784 867
0 869 7 1 2 778 868
0 870 5 1 1 869
0 871 7 1 2 1711 776
0 872 5 1 1 871
0 873 7 1 2 870 872
0 874 5 1 1 873
0 875 7 1 2 772 874
0 876 5 1 1 875
0 877 7 2 2 770 876
0 878 5 1 1 2239
0 879 7 1 2 1684 2240
0 880 5 1 1 879
0 881 7 1 2 1681 878
0 882 5 1 1 881
0 883 7 1 2 2160 682
0 884 5 1 1 883
0 885 7 1 2 2164 884
0 886 7 1 2 882 885
0 887 5 1 1 886
0 888 7 2 2 880 887
0 889 5 1 1 2241
0 890 7 1 2 1669 889
0 891 5 1 1 890
0 892 7 1 2 764 891
0 893 5 1 1 892
0 894 7 1 2 1666 2242
0 895 5 1 1 894
0 896 7 2 2 893 895
0 897 5 1 1 2243
0 898 7 1 2 2216 2244
0 899 5 1 1 898
0 900 7 1 2 1649 899
0 901 5 1 1 900
0 902 7 1 2 760 897
0 903 5 1 1 902
0 904 7 2 2 901 903
0 905 5 1 1 2245
0 906 7 1 2 1919 2246
0 907 5 1 1 906
0 908 7 1 2 1922 905
0 909 5 1 1 908
0 910 7 1 2 2178 706
0 911 5 1 1 910
0 912 7 1 2 2182 911
0 913 7 1 2 909 912
0 914 5 1 1 913
0 915 7 1 2 907 914
0 916 5 1 1 915
0 917 7 1 2 756 916
0 918 5 1 1 917
0 919 7 1 2 754 918
0 920 5 1 1 919
0 921 7 1 2 748 920
0 922 5 1 1 921
0 923 7 1 2 1643 2212
0 924 5 1 1 923
0 925 7 1 2 1906 2192
0 926 5 1 1 925
0 927 7 1 2 2195 926
0 928 7 1 2 1941 927
0 929 7 1 2 2206 928
0 930 7 1 2 2210 929
0 931 7 1 2 924 930
0 932 7 1 2 922 931
0 933 5 1 1 932
0 934 7 1 2 1832 2102
0 935 5 1 1 934
0 936 7 3 2 1829 935
0 937 5 3 1 2247
0 938 7 1 2 1821 2250
0 939 5 1 1 938
0 940 7 2 2 1818 939
0 941 5 2 1 2253
0 942 7 1 2 1807 2255
0 943 5 1 1 942
0 944 7 2 2 1804 943
0 945 5 2 1 2257
0 946 7 1 2 1792 2259
0 947 5 1 1 946
0 948 7 2 2 1789 947
0 949 5 2 1 2261
0 950 7 1 2 1777 2263
0 951 5 1 1 950
0 952 7 2 2 1774 951
0 953 5 2 1 2265
0 954 7 1 2 1764 2267
0 955 5 1 1 954
0 956 7 2 2 1761 955
0 957 5 2 1 2269
0 958 7 1 2 1749 2271
0 959 5 1 1 958
0 960 7 2 2 1746 959
0 961 5 2 1 2273
0 962 7 1 2 1736 2275
0 963 5 1 1 962
0 964 7 2 2 1733 963
0 965 5 2 1 2277
0 966 7 1 2 1721 2279
0 967 5 1 1 966
0 968 7 2 2 1718 967
0 969 5 2 1 2281
0 970 7 1 2 1706 2283
0 971 5 1 1 970
0 972 7 2 2 1703 971
0 973 5 2 1 2285
0 974 7 1 2 1691 2287
0 975 5 1 1 974
0 976 7 2 2 1688 975
0 977 5 2 1 2289
0 978 7 1 2 1676 2291
0 979 5 1 1 978
0 980 7 2 2 1673 979
0 981 5 2 1 2293
0 982 7 1 2 1653 2295
0 983 5 1 1 982
0 984 7 2 2 1656 983
0 985 5 2 1 2297
0 986 7 1 2 1929 2299
0 987 5 1 1 986
0 988 7 2 2 1926 987
0 989 5 2 1 2301
0 990 7 1 2 1904 2303
0 991 5 1 1 990
0 992 7 2 2 1909 991
0 993 5 2 1 2305
0 994 7 1 2 2193 2307
0 995 5 1 1 994
0 996 7 2 2 2196 995
0 997 5 2 1 2309
0 998 7 1 2 933 2310
0 999 5 1 1 998
0 1000 7 1 2 1661 2294
0 1001 5 1 1 1000
0 1002 7 1 2 1659 2296
0 1003 5 1 1 1002
0 1004 7 3 2 1001 1003
0 1005 5 2 1 2313
0 1006 7 1 2 1914 2302
0 1007 5 1 1 1006
0 1008 7 1 2 1912 2304
0 1009 5 1 1 1008
0 1010 7 2 2 1007 1009
0 1011 5 2 1 2318
0 1012 7 1 2 2314 2319
0 1013 5 2 1 1012
0 1014 7 1 2 1956 2298
0 1015 5 1 1 1014
0 1016 7 1 2 1958 2300
0 1017 5 1 1 1016
0 1018 7 3 2 1015 1017
0 1019 5 2 1 2324
0 1020 7 1 2 1948 2290
0 1021 5 1 1 1020
0 1022 7 1 2 1946 2292
0 1023 5 1 1 1022
0 1024 7 3 2 1021 1023
0 1025 5 2 1 2329
0 1026 7 1 2 2327 2330
0 1027 5 2 1 1026
0 1028 7 1 2 1970 2286
0 1029 5 1 1 1028
0 1030 7 1 2 1968 2288
0 1031 5 1 1 1030
0 1032 7 3 2 1029 1031
0 1033 5 2 1 2336
0 1034 7 1 2 2315 2337
0 1035 5 2 1 1034
0 1036 7 1 2 1982 2282
0 1037 5 1 1 1036
0 1038 7 1 2 1980 2284
0 1039 5 1 1 1038
0 1040 7 3 2 1037 1039
0 1041 5 2 1 2343
0 1042 7 1 2 2331 2344
0 1043 5 2 1 1042
0 1044 7 1 2 1994 2278
0 1045 5 1 1 1044
0 1046 7 1 2 1992 2280
0 1047 5 1 1 1046
0 1048 7 3 2 1045 1047
0 1049 5 2 1 2350
0 1050 7 1 2 2338 2351
0 1051 5 2 1 1050
0 1052 7 1 2 2006 2274
0 1053 5 1 1 1052
0 1054 7 1 2 2004 2276
0 1055 5 1 1 1054
0 1056 7 3 2 1053 1055
0 1057 5 2 1 2357
0 1058 7 1 2 2345 2358
0 1059 5 2 1 1058
0 1060 7 1 2 2018 2270
0 1061 5 1 1 1060
0 1062 7 1 2 2016 2272
0 1063 5 1 1 1062
0 1064 7 3 2 1061 1063
0 1065 5 2 1 2364
0 1066 7 1 2 2352 2365
0 1067 5 2 1 1066
0 1068 7 1 2 2030 2266
0 1069 5 1 1 1068
0 1070 7 1 2 2028 2268
0 1071 5 1 1 1070
0 1072 7 3 2 1069 1071
0 1073 5 2 1 2371
0 1074 7 1 2 2359 2372
0 1075 5 2 1 1074
0 1076 7 1 2 2042 2262
0 1077 5 1 1 1076
0 1078 7 1 2 2040 2264
0 1079 5 1 1 1078
0 1080 7 3 2 1077 1079
0 1081 5 2 1 2378
0 1082 7 1 2 2366 2379
0 1083 5 2 1 1082
0 1084 7 1 2 2054 2258
0 1085 5 1 1 1084
0 1086 7 1 2 2052 2260
0 1087 5 1 1 1086
0 1088 7 3 2 1085 1087
0 1089 5 2 1 2385
0 1090 7 1 2 2373 2386
0 1091 5 2 1 1090
0 1092 7 1 2 2066 2254
0 1093 5 1 1 1092
0 1094 7 1 2 2064 2256
0 1095 5 1 1 1094
0 1096 7 3 2 1093 1095
0 1097 5 2 1 2392
0 1098 7 1 2 2380 2393
0 1099 5 2 1 1098
0 1100 7 1 2 2078 2248
0 1101 5 1 1 1100
0 1102 7 1 2 2076 2251
0 1103 5 1 1 1102
0 1104 7 3 2 1101 1103
0 1105 5 2 1 2399
0 1106 7 1 2 2387 2400
0 1107 5 2 1 1106
0 1108 7 1 2 2088 2103
0 1109 5 1 1 1108
0 1110 7 1 2 2090 2099
0 1111 5 1 1 1110
0 1112 7 2 2 1109 1111
0 1113 5 1 1 2406
0 1114 7 1 2 2394 2407
0 1115 5 2 1 1114
0 1116 7 2 2 2108 2401
0 1117 5 2 1 2410
0 1118 7 1 2 2395 1113
0 1119 5 1 1 1118
0 1120 7 2 2 2408 1119
0 1121 5 1 1 2414
0 1122 7 1 2 2411 2415
0 1123 5 2 1 1122
0 1124 7 2 2 2409 2416
0 1125 5 1 1 2418
0 1126 7 1 2 2388 2402
0 1127 5 1 1 1126
0 1128 7 2 2 2404 1127
0 1129 5 1 1 2420
0 1130 7 1 2 1125 2421
0 1131 5 2 1 1130
0 1132 7 2 2 2405 2422
0 1133 5 1 1 2424
0 1134 7 1 2 2381 2396
0 1135 5 1 1 1134
0 1136 7 2 2 2397 1135
0 1137 5 1 1 2426
0 1138 7 1 2 1133 2427
0 1139 5 2 1 1138
0 1140 7 2 2 2398 2428
0 1141 5 1 1 2430
0 1142 7 1 2 2374 2389
0 1143 5 1 1 1142
0 1144 7 2 2 2390 1143
0 1145 5 1 1 2432
0 1146 7 1 2 1141 2433
0 1147 5 2 1 1146
0 1148 7 2 2 2391 2434
0 1149 5 1 1 2436
0 1150 7 1 2 2367 2382
0 1151 5 1 1 1150
0 1152 7 2 2 2383 1151
0 1153 5 1 1 2438
0 1154 7 1 2 1149 2439
0 1155 5 2 1 1154
0 1156 7 2 2 2384 2440
0 1157 5 1 1 2442
0 1158 7 1 2 2360 2375
0 1159 5 1 1 1158
0 1160 7 2 2 2376 1159
0 1161 5 1 1 2444
0 1162 7 1 2 1157 2445
0 1163 5 2 1 1162
0 1164 7 2 2 2377 2446
0 1165 5 1 1 2448
0 1166 7 1 2 2353 2368
0 1167 5 1 1 1166
0 1168 7 2 2 2369 1167
0 1169 5 1 1 2450
0 1170 7 1 2 1165 2451
0 1171 5 2 1 1170
0 1172 7 2 2 2370 2452
0 1173 5 1 1 2454
0 1174 7 1 2 2346 2361
0 1175 5 1 1 1174
0 1176 7 2 2 2362 1175
0 1177 5 1 1 2456
0 1178 7 1 2 1173 2457
0 1179 5 2 1 1178
0 1180 7 2 2 2363 2458
0 1181 5 1 1 2460
0 1182 7 1 2 2339 2354
0 1183 5 1 1 1182
0 1184 7 2 2 2355 1183
0 1185 5 1 1 2462
0 1186 7 1 2 1181 2463
0 1187 5 2 1 1186
0 1188 7 2 2 2356 2464
0 1189 5 1 1 2466
0 1190 7 1 2 2332 2347
0 1191 5 1 1 1190
0 1192 7 2 2 2348 1191
0 1193 5 1 1 2468
0 1194 7 1 2 1189 2469
0 1195 5 2 1 1194
0 1196 7 2 2 2349 2470
0 1197 5 1 1 2472
0 1198 7 1 2 2316 2340
0 1199 5 1 1 1198
0 1200 7 2 2 2341 1199
0 1201 5 1 1 2474
0 1202 7 1 2 1197 2475
0 1203 5 2 1 1202
0 1204 7 2 2 2342 2476
0 1205 5 1 1 2478
0 1206 7 1 2 2325 2333
0 1207 5 1 1 1206
0 1208 7 2 2 2334 1207
0 1209 5 1 1 2480
0 1210 7 1 2 1205 2481
0 1211 5 2 1 1210
0 1212 7 2 2 2335 2482
0 1213 5 1 1 2484
0 1214 7 1 2 2317 2320
0 1215 5 1 1 1214
0 1216 7 2 2 2322 1215
0 1217 5 1 1 2486
0 1218 7 1 2 1213 2487
0 1219 5 2 1 1218
0 1220 7 2 2 2323 2488
0 1221 5 1 1 2490
0 1222 7 1 2 2199 2308
0 1223 5 1 1 1222
0 1224 7 1 2 2201 2306
0 1225 5 1 1 1224
0 1226 7 2 2 1223 1225
0 1227 5 2 1 2492
0 1228 7 1 2 2326 2493
0 1229 5 1 1 1228
0 1230 7 1 2 2328 2494
0 1231 5 1 1 1230
0 1232 7 2 2 1229 1231
0 1233 5 1 1 2496
0 1234 7 1 2 1221 1233
0 1235 5 2 1 1234
0 1236 7 1 2 2491 2497
0 1237 5 1 1 1236
0 1238 7 2 2 2498 1237
0 1239 5 1 1 2500
0 1240 7 1 2 1641 1239
0 1241 5 1 1 1240
0 1242 7 1 2 2485 1217
0 1243 5 1 1 1242
0 1244 7 2 2 2489 1243
0 1245 5 1 1 2502
0 1246 7 1 2 1898 2503
0 1247 5 1 1 1246
0 1248 7 1 2 1901 1245
0 1249 5 1 1 1248
0 1250 7 1 2 2473 1201
0 1251 5 1 1 1250
0 1252 7 2 2 2477 1251
0 1253 5 1 1 2504
0 1254 7 1 2 2467 1193
0 1255 5 1 1 1254
0 1256 7 1 2 2471 1255
0 1257 5 1 1 1256
0 1258 7 1 2 2455 1177
0 1259 5 1 1 1258
0 1260 7 2 2 2459 1259
0 1261 5 1 1 2506
0 1262 7 1 2 1697 1261
0 1263 5 1 1 1262
0 1264 7 1 2 1700 2507
0 1265 5 1 1 1264
0 1266 7 1 2 2449 1169
0 1267 5 1 1 1266
0 1268 7 2 2 2453 1267
0 1269 5 1 1 2508
0 1270 7 1 2 1715 2509
0 1271 5 1 1 1270
0 1272 7 1 2 2443 1161
0 1273 5 1 1 1272
0 1274 7 2 2 2447 1273
0 1275 5 1 1 2510
0 1276 7 1 2 1730 2511
0 1277 5 1 1 1276
0 1278 7 1 2 1727 1275
0 1279 5 1 1 1278
0 1280 7 1 2 2437 1153
0 1281 5 1 1 1280
0 1282 7 2 2 2441 1281
0 1283 5 1 1 2512
0 1284 7 1 2 2431 1145
0 1285 5 1 1 1284
0 1286 7 2 2 2435 1285
0 1287 5 1 1 2514
0 1288 7 1 2 1758 2515
0 1289 5 1 1 1288
0 1290 7 1 2 1755 1287
0 1291 5 1 1 1290
0 1292 7 1 2 2425 1137
0 1293 5 1 1 1292
0 1294 7 2 2 2429 1293
0 1295 5 1 1 2516
0 1296 7 1 2 2419 1129
0 1297 5 1 1 1296
0 1298 7 2 2 2423 1297
0 1299 5 1 1 2518
0 1300 7 1 2 1786 2519
0 1301 5 1 1 1300
0 1302 7 1 2 1783 1299
0 1303 5 1 1 1302
0 1304 7 1 2 2106 2403
0 1305 5 1 1 1304
0 1306 7 2 2 2412 1305
0 1307 5 1 1 2520
0 1308 7 1 2 2249 2521
0 1309 5 1 1 1308
0 1310 7 1 2 1813 1309
0 1311 5 1 1 1310
0 1312 7 1 2 2252 1307
0 1313 5 1 1 1312
0 1314 7 2 2 1311 1313
0 1315 5 1 1 2522
0 1316 7 1 2 1798 1315
0 1317 5 1 1 1316
0 1318 7 1 2 2413 1121
0 1319 5 1 1 1318
0 1320 7 1 2 2417 1319
0 1321 7 1 2 1317 1320
0 1322 5 1 1 1321
0 1323 7 1 2 1801 2523
0 1324 5 1 1 1323
0 1325 7 1 2 1322 1324
0 1326 5 1 1 1325
0 1327 7 1 2 1303 1326
0 1328 5 1 1 1327
0 1329 7 2 2 1301 1328
0 1330 5 1 1 2524
0 1331 7 1 2 2517 1330
0 1332 5 1 1 1331
0 1333 7 1 2 1295 2525
0 1334 5 1 1 1333
0 1335 7 1 2 1771 1334
0 1336 5 1 1 1335
0 1337 7 1 2 1332 1336
0 1338 5 1 1 1337
0 1339 7 1 2 1291 1338
0 1340 5 1 1 1339
0 1341 7 2 2 1289 1340
0 1342 5 1 1 2526
0 1343 7 1 2 2513 1342
0 1344 5 1 1 1343
0 1345 7 1 2 1283 2527
0 1346 5 1 1 1345
0 1347 7 1 2 1743 1346
0 1348 5 1 1 1347
0 1349 7 1 2 1344 1348
0 1350 5 1 1 1349
0 1351 7 1 2 1279 1350
0 1352 5 1 1 1351
0 1353 7 1 2 1277 1352
0 1354 7 1 2 1271 1353
0 1355 5 1 1 1354
0 1356 7 1 2 1712 1269
0 1357 5 1 1 1356
0 1358 7 1 2 1355 1357
0 1359 5 1 1 1358
0 1360 7 1 2 1265 1359
0 1361 5 1 1 1360
0 1362 7 2 2 1263 1361
0 1363 5 1 1 2528
0 1364 7 1 2 1685 2529
0 1365 5 1 1 1364
0 1366 7 1 2 1682 1363
0 1367 5 1 1 1366
0 1368 7 1 2 2461 1185
0 1369 5 1 1 1368
0 1370 7 1 2 2465 1369
0 1371 7 1 2 1367 1370
0 1372 5 1 1 1371
0 1373 7 2 2 1365 1372
0 1374 5 1 1 2530
0 1375 7 1 2 1670 1374
0 1376 5 1 1 1375
0 1377 7 1 2 1257 1376
0 1378 5 1 1 1377
0 1379 7 1 2 1667 2531
0 1380 5 1 1 1379
0 1381 7 2 2 1378 1380
0 1382 5 1 1 2532
0 1383 7 1 2 2505 2533
0 1384 5 1 1 1383
0 1385 7 1 2 1650 1384
0 1386 5 1 1 1385
0 1387 7 1 2 1253 1382
0 1388 5 1 1 1387
0 1389 7 2 2 1386 1388
0 1390 5 1 1 2534
0 1391 7 1 2 1920 2535
0 1392 5 1 1 1391
0 1393 7 1 2 1923 1390
0 1394 5 1 1 1393
0 1395 7 1 2 2479 1209
0 1396 5 1 1 1395
0 1397 7 1 2 2483 1396
0 1398 7 1 2 1394 1397
0 1399 5 1 1 1398
0 1400 7 1 2 1392 1399
0 1401 5 1 1 1400
0 1402 7 1 2 1249 1401
0 1403 5 1 1 1402
0 1404 7 1 2 1247 1403
0 1405 5 1 1 1404
0 1406 7 1 2 1241 1405
0 1407 5 1 1 1406
0 1408 7 1 2 1644 2501
0 1409 5 1 1 1408
0 1410 7 1 2 2311 2321
0 1411 7 1 2 2495 1410
0 1412 7 1 2 2499 1411
0 1413 7 1 2 1409 1412
0 1414 7 1 2 1407 1413
0 1415 5 1 1 1414
0 1416 7 1 2 2312 1415
0 1417 5 1 1 1416
3 3499 7 0 2 999 1417
