1 0 0 2 0
2 49 1 0
2 1656 1 0
1 1 0 2 0
2 1657 1 1
2 1658 1 1
1 2 0 2 0
2 1659 1 2
2 1660 1 2
1 3 0 2 0
2 1661 1 3
2 1662 1 3
1 4 0 2 0
2 1663 1 4
2 1664 1 4
1 5 0 2 0
2 1665 1 5
2 1666 1 5
1 6 0 2 0
2 1667 1 6
2 1668 1 6
1 7 0 2 0
2 1669 1 7
2 1670 1 7
1 8 0 2 0
2 1671 1 8
2 1672 1 8
1 9 0 2 0
2 1673 1 9
2 1674 1 9
1 10 0 2 0
2 1675 1 10
2 1676 1 10
1 11 0 2 0
2 1677 1 11
2 1678 1 11
1 12 0 2 0
2 1679 1 12
2 1680 1 12
1 13 0 2 0
2 1681 1 13
2 1682 1 13
1 14 0 2 0
2 1683 1 14
2 1684 1 14
1 15 0 2 0
2 1685 1 15
2 1686 1 15
1 16 0 2 0
2 1687 1 16
2 1688 1 16
1 17 0 2 0
2 1689 1 17
2 1690 1 17
1 18 0 2 0
2 1691 1 18
2 1692 1 18
1 19 0 2 0
2 1693 1 19
2 1694 1 19
1 20 0 2 0
2 1695 1 20
2 1696 1 20
1 21 0 2 0
2 1697 1 21
2 1698 1 21
1 22 0 2 0
2 1699 1 22
2 1700 1 22
1 23 0 2 0
2 1701 1 23
2 1702 1 23
1 24 0 2 0
2 1703 1 24
2 1704 1 24
1 25 0 2 0
2 1705 1 25
2 1706 1 25
1 26 0 2 0
2 1707 1 26
2 1708 1 26
1 27 0 2 0
2 1709 1 27
2 1710 1 27
1 28 0 2 0
2 1711 1 28
2 1712 1 28
1 29 0 2 0
2 1713 1 29
2 1714 1 29
1 30 0 2 0
2 1715 1 30
2 1716 1 30
1 31 0 2 0
2 1717 1 31
2 1718 1 31
1 32 0 2 0
2 1719 1 32
2 1720 1 32
1 33 0 2 0
2 1721 1 33
2 1722 1 33
1 34 0 2 0
2 1723 1 34
2 1724 1 34
1 35 0 2 0
2 1725 1 35
2 1726 1 35
1 36 0 2 0
2 1727 1 36
2 1728 1 36
1 37 0 2 0
2 1729 1 37
2 1730 1 37
1 38 0 2 0
2 1731 1 38
2 1732 1 38
1 39 0 2 0
2 1733 1 39
2 1734 1 39
1 40 0 2 0
2 1735 1 40
2 1736 1 40
1 41 0 2 0
2 1737 1 41
2 1738 1 41
1 42 0 2 0
2 1739 1 42
2 1740 1 42
1 43 0 2 0
2 1741 1 43
2 1742 1 43
1 44 0 2 0
2 1743 1 44
2 1744 1 44
1 45 0 2 0
2 1745 1 45
2 1746 1 45
1 46 0 2 0
2 1747 1 46
2 1748 1 46
1 47 0 2 0
2 1749 1 47
2 1750 1 47
1 48 0 2 0
2 1751 1 48
2 1752 1 48
2 1753 1 69
2 1754 1 69
2 1755 1 70
2 1756 1 70
2 1757 1 71
2 1758 1 71
2 1759 1 72
2 1760 1 72
2 1761 1 73
2 1762 1 73
2 1763 1 74
2 1764 1 74
2 1765 1 75
2 1766 1 75
2 1767 1 76
2 1768 1 76
2 1769 1 77
2 1770 1 77
2 1771 1 78
2 1772 1 78
2 1773 1 79
2 1774 1 79
2 1775 1 80
2 1776 1 80
2 1777 1 81
2 1778 1 81
2 1779 1 100
2 1780 1 100
2 1781 1 102
2 1782 1 102
2 1783 1 104
2 1784 1 104
2 1785 1 106
2 1786 1 106
2 1787 1 107
2 1788 1 107
2 1789 1 108
2 1790 1 108
2 1791 1 108
2 1792 1 111
2 1793 1 111
2 1794 1 112
2 1795 1 112
2 1796 1 115
2 1797 1 115
2 1798 1 118
2 1799 1 118
2 1800 1 120
2 1801 1 120
2 1802 1 123
2 1803 1 123
2 1804 1 126
2 1805 1 126
2 1806 1 128
2 1807 1 128
2 1808 1 131
2 1809 1 131
2 1810 1 134
2 1811 1 134
2 1812 1 136
2 1813 1 136
2 1814 1 139
2 1815 1 139
2 1816 1 142
2 1817 1 142
2 1818 1 144
2 1819 1 144
2 1820 1 147
2 1821 1 147
2 1822 1 150
2 1823 1 150
2 1824 1 152
2 1825 1 152
2 1826 1 155
2 1827 1 155
2 1828 1 158
2 1829 1 158
2 1830 1 160
2 1831 1 160
2 1832 1 163
2 1833 1 163
2 1834 1 166
2 1835 1 166
2 1836 1 168
2 1837 1 168
2 1838 1 171
2 1839 1 171
2 1840 1 174
2 1841 1 174
2 1842 1 176
2 1843 1 176
2 1844 1 179
2 1845 1 179
2 1846 1 182
2 1847 1 182
2 1848 1 184
2 1849 1 184
2 1850 1 187
2 1851 1 187
2 1852 1 190
2 1853 1 190
2 1854 1 192
2 1855 1 192
2 1856 1 195
2 1857 1 195
2 1858 1 198
2 1859 1 198
2 1860 1 200
2 1861 1 200
2 1862 1 203
2 1863 1 203
2 1864 1 206
2 1865 1 206
2 1866 1 208
2 1867 1 208
2 1868 1 209
2 1869 1 209
2 1870 1 215
2 1871 1 215
2 1872 1 215
2 1873 1 215
2 1874 1 216
2 1875 1 216
2 1876 1 216
2 1877 1 218
2 1878 1 218
2 1879 1 218
2 1880 1 220
2 1881 1 220
2 1882 1 220
2 1883 1 221
2 1884 1 221
2 1885 1 221
2 1886 1 222
2 1887 1 222
2 1888 1 223
2 1889 1 223
2 1890 1 229
2 1891 1 229
2 1892 1 229
2 1893 1 229
2 1894 1 230
2 1895 1 230
2 1896 1 230
2 1897 1 232
2 1898 1 232
2 1899 1 232
2 1900 1 234
2 1901 1 234
2 1902 1 234
2 1903 1 235
2 1904 1 235
2 1905 1 241
2 1906 1 241
2 1907 1 241
2 1908 1 241
2 1909 1 242
2 1910 1 242
2 1911 1 242
2 1912 1 244
2 1913 1 244
2 1914 1 244
2 1915 1 246
2 1916 1 246
2 1917 1 246
2 1918 1 247
2 1919 1 247
2 1920 1 253
2 1921 1 253
2 1922 1 254
2 1923 1 254
2 1924 1 254
2 1925 1 256
2 1926 1 256
2 1927 1 256
2 1928 1 258
2 1929 1 258
2 1930 1 258
2 1931 1 259
2 1932 1 259
2 1933 1 265
2 1934 1 265
2 1935 1 265
2 1936 1 265
2 1937 1 266
2 1938 1 266
2 1939 1 266
2 1940 1 268
2 1941 1 268
2 1942 1 268
2 1943 1 270
2 1944 1 270
2 1945 1 270
2 1946 1 271
2 1947 1 271
2 1948 1 277
2 1949 1 277
2 1950 1 278
2 1951 1 278
2 1952 1 278
2 1953 1 280
2 1954 1 280
2 1955 1 280
2 1956 1 282
2 1957 1 282
2 1958 1 282
2 1959 1 283
2 1960 1 283
2 1961 1 289
2 1962 1 289
2 1963 1 289
2 1964 1 289
2 1965 1 290
2 1966 1 290
2 1967 1 290
2 1968 1 292
2 1969 1 292
2 1970 1 292
2 1971 1 294
2 1972 1 294
2 1973 1 294
2 1974 1 295
2 1975 1 295
2 1976 1 301
2 1977 1 301
2 1978 1 301
2 1979 1 301
2 1980 1 302
2 1981 1 302
2 1982 1 302
2 1983 1 304
2 1984 1 304
2 1985 1 304
2 1986 1 306
2 1987 1 306
2 1988 1 306
2 1989 1 307
2 1990 1 307
2 1991 1 313
2 1992 1 313
2 1993 1 313
2 1994 1 313
2 1995 1 314
2 1996 1 314
2 1997 1 314
2 1998 1 316
2 1999 1 316
2 2000 1 316
2 2001 1 318
2 2002 1 318
2 2003 1 318
2 2004 1 319
2 2005 1 319
2 2006 1 325
2 2007 1 325
2 2008 1 325
2 2009 1 325
2 2010 1 326
2 2011 1 326
2 2012 1 326
2 2013 1 328
2 2014 1 328
2 2015 1 328
2 2016 1 330
2 2017 1 330
2 2018 1 330
2 2019 1 331
2 2020 1 331
2 2021 1 337
2 2022 1 337
2 2023 1 337
2 2024 1 338
2 2025 1 338
2 2026 1 340
2 2027 1 340
2 2028 1 340
2 2029 1 342
2 2030 1 342
2 2031 1 342
2 2032 1 343
2 2033 1 343
2 2034 1 349
2 2035 1 349
2 2036 1 350
2 2037 1 350
2 2038 1 352
2 2039 1 352
2 2040 1 352
2 2041 1 354
2 2042 1 354
2 2043 1 354
2 2044 1 355
2 2045 1 355
2 2046 1 361
2 2047 1 361
2 2048 1 364
2 2049 1 364
2 2050 1 364
2 2051 1 366
2 2052 1 366
2 2053 1 366
2 2054 1 367
2 2055 1 367
2 2056 1 373
2 2057 1 373
2 2058 1 376
2 2059 1 376
2 2060 1 376
2 2061 1 378
2 2062 1 378
2 2063 1 378
2 2064 1 381
2 2065 1 381
2 2066 1 383
2 2067 1 383
2 2068 1 383
2 2069 1 384
2 2070 1 384
2 2071 1 387
2 2072 1 387
2 2073 1 388
2 2074 1 388
2 2075 1 391
2 2076 1 391
2 2077 1 392
2 2078 1 392
2 2079 1 395
2 2080 1 395
2 2081 1 396
2 2082 1 396
2 2083 1 399
2 2084 1 399
2 2085 1 400
2 2086 1 400
2 2087 1 403
2 2088 1 403
2 2089 1 404
2 2090 1 404
2 2091 1 407
2 2092 1 407
2 2093 1 408
2 2094 1 408
2 2095 1 411
2 2096 1 411
2 2097 1 412
2 2098 1 412
2 2099 1 415
2 2100 1 415
2 2101 1 416
2 2102 1 416
2 2103 1 419
2 2104 1 419
2 2105 1 420
2 2106 1 420
2 2107 1 423
2 2108 1 423
2 2109 1 424
2 2110 1 424
2 2111 1 427
2 2112 1 427
2 2113 1 428
2 2114 1 428
2 2115 1 431
2 2116 1 431
2 2117 1 432
2 2118 1 432
2 2119 1 435
2 2120 1 435
2 2121 1 436
2 2122 1 436
2 2123 1 441
2 2124 1 441
2 2125 1 441
2 2126 1 441
2 2127 1 442
2 2128 1 442
2 2129 1 442
2 2130 1 445
2 2131 1 445
2 2132 1 448
2 2133 1 448
2 2134 1 450
2 2135 1 450
2 2136 1 453
2 2137 1 453
2 2138 1 453
2 2139 1 453
2 2140 1 454
2 2141 1 454
2 2142 1 454
2 2143 1 456
2 2144 1 456
2 2145 1 456
2 2146 1 456
2 2147 1 458
2 2148 1 458
2 2149 1 458
2 2150 1 458
2 2151 1 459
2 2152 1 459
2 2153 1 465
2 2154 1 465
2 2155 1 465
2 2156 1 465
2 2157 1 466
2 2158 1 466
2 2159 1 466
2 2160 1 468
2 2161 1 468
2 2162 1 468
2 2163 1 470
2 2164 1 470
2 2165 1 470
2 2166 1 473
2 2167 1 473
2 2168 1 474
2 2169 1 474
2 2170 1 477
2 2171 1 477
2 2172 1 477
2 2173 1 478
2 2174 1 478
2 2175 1 478
2 2176 1 481
2 2177 1 481
2 2178 1 481
2 2179 1 481
2 2180 1 482
2 2181 1 482
2 2182 1 483
2 2183 1 483
2 2184 1 483
2 2185 1 484
2 2186 1 484
2 2187 1 489
2 2188 1 489
2 2189 1 489
2 2190 1 490
2 2191 1 490
2 2192 1 490
2 2193 1 495
2 2194 1 495
2 2195 1 499
2 2196 1 499
2 2197 1 499
2 2198 1 500
2 2199 1 500
2 2200 1 505
2 2201 1 505
2 2202 1 505
2 2203 1 505
2 2204 1 506
2 2205 1 506
2 2206 1 506
2 2207 1 511
2 2208 1 511
2 2209 1 513
2 2210 1 513
2 2211 1 513
2 2212 1 514
2 2213 1 514
2 2214 1 519
2 2215 1 519
2 2216 1 519
2 2217 1 519
2 2218 1 520
2 2219 1 520
2 2220 1 520
2 2221 1 522
2 2222 1 522
2 2223 1 535
2 2224 1 535
2 2225 1 535
2 2226 1 536
2 2227 1 536
2 2228 1 541
2 2229 1 541
2 2230 1 541
2 2231 1 541
2 2232 1 542
2 2233 1 542
2 2234 1 542
2 2235 1 544
2 2236 1 544
2 2237 1 547
2 2238 1 547
2 2239 1 549
2 2240 1 549
2 2241 1 549
2 2242 1 550
2 2243 1 550
2 2244 1 555
2 2245 1 555
2 2246 1 555
2 2247 1 555
2 2248 1 556
2 2249 1 556
2 2250 1 556
2 2251 1 558
2 2252 1 558
2 2253 1 559
2 2254 1 559
2 2255 1 561
2 2256 1 561
2 2257 1 561
2 2258 1 562
2 2259 1 562
2 2260 1 567
2 2261 1 567
2 2262 1 567
2 2263 1 567
2 2264 1 568
2 2265 1 568
2 2266 1 568
2 2267 1 570
2 2268 1 570
2 2269 1 573
2 2270 1 573
2 2271 1 576
2 2272 1 576
2 2273 1 579
2 2274 1 579
2 2275 1 582
2 2276 1 582
2 2277 1 583
2 2278 1 583
2 2279 1 583
2 2280 1 584
2 2281 1 584
2 2282 1 589
2 2283 1 589
2 2284 1 589
2 2285 1 589
2 2286 1 590
2 2287 1 590
2 2288 1 590
2 2289 1 591
2 2290 1 591
2 2291 1 591
2 2292 1 592
2 2293 1 592
2 2294 1 597
2 2295 1 597
2 2296 1 597
2 2297 1 597
2 2298 1 598
2 2299 1 598
2 2300 1 598
2 2301 1 600
2 2302 1 600
2 2303 1 603
2 2304 1 603
2 2305 1 606
2 2306 1 606
2 2307 1 607
2 2308 1 607
2 2309 1 611
2 2310 1 611
2 2311 1 614
2 2312 1 614
2 2313 1 615
2 2314 1 615
2 2315 1 615
2 2316 1 616
2 2317 1 616
2 2318 1 621
2 2319 1 621
2 2320 1 621
2 2321 1 621
2 2322 1 622
2 2323 1 622
2 2324 1 622
2 2325 1 624
2 2326 1 624
2 2327 1 627
2 2328 1 627
2 2329 1 630
2 2330 1 630
2 2331 1 631
2 2332 1 631
2 2333 1 635
2 2334 1 635
2 2335 1 638
2 2336 1 638
2 2337 1 639
2 2338 1 639
2 2339 1 639
2 2340 1 640
2 2341 1 640
2 2342 1 645
2 2343 1 645
2 2344 1 645
2 2345 1 645
2 2346 1 646
2 2347 1 646
2 2348 1 646
2 2349 1 648
2 2350 1 648
2 2351 1 651
2 2352 1 651
2 2353 1 654
2 2354 1 654
2 2355 1 655
2 2356 1 655
2 2357 1 659
2 2358 1 659
2 2359 1 662
2 2360 1 662
2 2361 1 663
2 2362 1 663
2 2363 1 663
2 2364 1 664
2 2365 1 664
2 2366 1 669
2 2367 1 669
2 2368 1 669
2 2369 1 669
2 2370 1 669
2 2371 1 670
2 2372 1 670
2 2373 1 670
2 2374 1 672
2 2375 1 672
2 2376 1 675
2 2377 1 675
2 2378 1 678
2 2379 1 678
2 2380 1 679
2 2381 1 679
2 2382 1 683
2 2383 1 683
2 2384 1 686
2 2385 1 686
2 2386 1 687
2 2387 1 687
2 2388 1 687
2 2389 1 688
2 2390 1 688
2 2391 1 693
2 2392 1 693
2 2393 1 693
2 2394 1 693
2 2395 1 694
2 2396 1 694
2 2397 1 694
2 2398 1 696
2 2399 1 696
2 2400 1 699
2 2401 1 699
2 2402 1 702
2 2403 1 702
2 2404 1 703
2 2405 1 703
2 2406 1 707
2 2407 1 707
2 2408 1 710
2 2409 1 710
2 2410 1 711
2 2411 1 711
2 2412 1 711
2 2413 1 712
2 2414 1 712
2 2415 1 717
2 2416 1 717
2 2417 1 717
2 2418 1 717
2 2419 1 718
2 2420 1 718
2 2421 1 720
2 2422 1 720
2 2423 1 723
2 2424 1 723
2 2425 1 726
2 2426 1 726
2 2427 1 727
2 2428 1 727
2 2429 1 731
2 2430 1 731
2 2431 1 734
2 2432 1 734
2 2433 1 735
2 2434 1 735
2 2435 1 736
2 2436 1 736
2 2437 1 739
2 2438 1 739
2 2439 1 742
2 2440 1 742
2 2441 1 745
2 2442 1 745
2 2443 1 747
2 2444 1 747
2 2445 1 748
2 2446 1 748
2 2447 1 748
2 2448 1 749
2 2449 1 749
2 2450 1 749
2 2451 1 750
2 2452 1 750
2 2453 1 750
2 2454 1 750
2 2455 1 750
2 2456 1 753
2 2457 1 753
2 2458 1 754
2 2459 1 754
2 2460 1 757
2 2461 1 757
2 2462 1 760
2 2463 1 760
2 2464 1 761
2 2465 1 761
2 2466 1 765
2 2467 1 765
2 2468 1 768
2 2469 1 768
2 2470 1 769
2 2471 1 769
2 2472 1 773
2 2473 1 773
2 2474 1 776
2 2475 1 776
2 2476 1 777
2 2477 1 777
2 2478 1 781
2 2479 1 781
2 2480 1 784
2 2481 1 784
2 2482 1 785
2 2483 1 785
2 2484 1 789
2 2485 1 789
2 2486 1 792
2 2487 1 792
2 2488 1 793
2 2489 1 793
2 2490 1 797
2 2491 1 797
2 2492 1 800
2 2493 1 800
2 2494 1 801
2 2495 1 801
2 2496 1 805
2 2497 1 805
2 2498 1 808
2 2499 1 808
2 2500 1 809
2 2501 1 809
2 2502 1 813
2 2503 1 813
2 2504 1 816
2 2505 1 816
2 2506 1 817
2 2507 1 817
2 2508 1 819
2 2509 1 819
2 2510 1 821
2 2511 1 821
2 2512 1 821
2 2513 1 822
2 2514 1 822
2 2515 1 827
2 2516 1 827
2 2517 1 827
2 2518 1 830
2 2519 1 830
2 2520 1 833
2 2521 1 833
2 2522 1 836
2 2523 1 836
2 2524 1 839
2 2525 1 839
2 2526 1 842
2 2527 1 842
2 2528 1 845
2 2529 1 845
2 2530 1 848
2 2531 1 848
2 2532 1 851
2 2533 1 851
2 2534 1 857
2 2535 1 857
2 2536 1 863
2 2537 1 863
2 2538 1 871
2 2539 1 871
2 2540 1 879
2 2541 1 879
2 2542 1 883
2 2543 1 883
2 2544 1 891
2 2545 1 891
2 2546 1 895
2 2547 1 895
2 2548 1 901
2 2549 1 901
2 2550 1 902
2 2551 1 902
2 2552 1 907
2 2553 1 907
2 2554 1 915
2 2555 1 915
2 2556 1 925
2 2557 1 925
2 2558 1 928
2 2559 1 928
2 2560 1 930
2 2561 1 930
2 2562 1 948
2 2563 1 948
2 2564 1 960
2 2565 1 960
2 2566 1 975
2 2567 1 975
2 2568 1 996
2 2569 1 996
2 2570 1 1002
2 2571 1 1002
2 2572 1 1005
2 2573 1 1005
2 2574 1 1008
2 2575 1 1008
2 2576 1 1011
2 2577 1 1011
2 2578 1 1016
2 2579 1 1016
2 2580 1 1016
2 2581 1 1017
2 2582 1 1017
2 2583 1 1022
2 2584 1 1022
2 2585 1 1022
2 2586 1 1025
2 2587 1 1025
2 2588 1 1050
2 2589 1 1050
2 2590 1 1051
2 2591 1 1051
2 2592 1 1054
2 2593 1 1054
2 2594 1 1055
2 2595 1 1055
2 2596 1 1058
2 2597 1 1058
2 2598 1 1059
2 2599 1 1059
2 2600 1 1062
2 2601 1 1062
2 2602 1 1063
2 2603 1 1063
2 2604 1 1066
2 2605 1 1066
2 2606 1 1067
2 2607 1 1067
2 2608 1 1070
2 2609 1 1070
2 2610 1 1071
2 2611 1 1071
2 2612 1 1074
2 2613 1 1074
2 2614 1 1075
2 2615 1 1075
2 2616 1 1078
2 2617 1 1078
2 2618 1 1079
2 2619 1 1079
2 2620 1 1082
2 2621 1 1082
2 2622 1 1083
2 2623 1 1083
2 2624 1 1086
2 2625 1 1086
2 2626 1 1087
2 2627 1 1087
2 2628 1 1090
2 2629 1 1090
2 2630 1 1091
2 2631 1 1091
2 2632 1 1094
2 2633 1 1094
2 2634 1 1095
2 2635 1 1095
2 2636 1 1098
2 2637 1 1098
2 2638 1 1099
2 2639 1 1099
2 2640 1 1102
2 2641 1 1102
2 2642 1 1103
2 2643 1 1103
2 2644 1 1106
2 2645 1 1106
2 2646 1 1107
2 2647 1 1107
2 2648 1 1110
2 2649 1 1110
2 2650 1 1110
2 2651 1 1110
2 2652 1 1111
2 2653 1 1111
2 2654 1 1123
2 2655 1 1123
2 2656 1 1123
2 2657 1 1123
2 2658 1 1124
2 2659 1 1124
2 2660 1 1124
2 2661 1 1129
2 2662 1 1129
2 2663 1 1131
2 2664 1 1131
2 2665 1 1135
2 2666 1 1135
2 2667 1 1135
2 2668 1 1136
2 2669 1 1136
2 2670 1 1147
2 2671 1 1147
2 2672 1 1147
2 2673 1 1147
2 2674 1 1148
2 2675 1 1148
2 2676 1 1148
2 2677 1 1148
2 2678 1 1150
2 2679 1 1150
2 2680 1 1153
2 2681 1 1153
2 2682 1 1159
2 2683 1 1159
2 2684 1 1159
2 2685 1 1160
2 2686 1 1160
2 2687 1 1160
2 2688 1 1167
2 2689 1 1167
2 2690 1 1167
2 2691 1 1168
2 2692 1 1168
2 2693 1 1168
2 2694 1 1168
2 2695 1 1173
2 2696 1 1173
2 2697 1 1178
2 2698 1 1178
2 2699 1 1196
2 2700 1 1196
2 2701 1 1196
2 2702 1 1196
2 2703 1 1197
2 2704 1 1197
2 2705 1 1197
2 2706 1 1202
2 2707 1 1202
2 2708 1 1202
2 2709 1 1203
2 2710 1 1203
2 2711 1 1203
2 2712 1 1205
2 2713 1 1205
2 2714 1 1208
2 2715 1 1208
2 2716 1 1214
2 2717 1 1214
2 2718 1 1214
2 2719 1 1214
2 2720 1 1215
2 2721 1 1215
2 2722 1 1215
2 2723 1 1217
2 2724 1 1217
2 2725 1 1218
2 2726 1 1218
2 2727 1 1224
2 2728 1 1224
2 2729 1 1224
2 2730 1 1224
2 2731 1 1225
2 2732 1 1225
2 2733 1 1225
2 2734 1 1227
2 2735 1 1227
2 2736 1 1230
2 2737 1 1230
2 2738 1 1233
2 2739 1 1233
2 2740 1 1236
2 2741 1 1236
2 2742 1 1239
2 2743 1 1239
2 2744 1 1244
2 2745 1 1244
2 2746 1 1244
2 2747 1 1244
2 2748 1 1245
2 2749 1 1245
2 2750 1 1245
2 2751 1 1250
2 2752 1 1250
2 2753 1 1250
2 2754 1 1250
2 2755 1 1251
2 2756 1 1251
2 2757 1 1251
2 2758 1 1253
2 2759 1 1253
2 2760 1 1256
2 2761 1 1256
2 2762 1 1259
2 2763 1 1259
2 2764 1 1260
2 2765 1 1260
2 2766 1 1264
2 2767 1 1264
2 2768 1 1267
2 2769 1 1267
2 2770 1 1272
2 2771 1 1272
2 2772 1 1272
2 2773 1 1272
2 2774 1 1273
2 2775 1 1273
2 2776 1 1273
2 2777 1 1275
2 2778 1 1275
2 2779 1 1278
2 2780 1 1278
2 2781 1 1281
2 2782 1 1281
2 2783 1 1282
2 2784 1 1282
2 2785 1 1286
2 2786 1 1286
2 2787 1 1289
2 2788 1 1289
2 2789 1 1294
2 2790 1 1294
2 2791 1 1294
2 2792 1 1294
2 2793 1 1295
2 2794 1 1295
2 2795 1 1295
2 2796 1 1297
2 2797 1 1297
2 2798 1 1300
2 2799 1 1300
2 2800 1 1303
2 2801 1 1303
2 2802 1 1304
2 2803 1 1304
2 2804 1 1308
2 2805 1 1308
2 2806 1 1311
2 2807 1 1311
2 2808 1 1316
2 2809 1 1316
2 2810 1 1316
2 2811 1 1316
2 2812 1 1317
2 2813 1 1317
2 2814 1 1317
2 2815 1 1317
2 2816 1 1319
2 2817 1 1319
2 2818 1 1322
2 2819 1 1322
2 2820 1 1325
2 2821 1 1325
2 2822 1 1326
2 2823 1 1326
2 2824 1 1330
2 2825 1 1330
2 2826 1 1333
2 2827 1 1333
2 2828 1 1338
2 2829 1 1338
2 2830 1 1338
2 2831 1 1338
2 2832 1 1339
2 2833 1 1339
2 2834 1 1341
2 2835 1 1341
2 2836 1 1344
2 2837 1 1344
2 2838 1 1347
2 2839 1 1347
2 2840 1 1348
2 2841 1 1348
2 2842 1 1352
2 2843 1 1352
2 2844 1 1355
2 2845 1 1355
2 2846 1 1360
2 2847 1 1360
2 2848 1 1360
2 2849 1 1361
2 2850 1 1361
2 2851 1 1361
2 2852 1 1363
2 2853 1 1363
2 2854 1 1366
2 2855 1 1366
2 2856 1 1369
2 2857 1 1369
2 2858 1 1370
2 2859 1 1370
2 2860 1 1374
2 2861 1 1374
2 2862 1 1377
2 2863 1 1377
2 2864 1 1378
2 2865 1 1378
2 2866 1 1379
2 2867 1 1379
2 2868 1 1382
2 2869 1 1382
2 2870 1 1385
2 2871 1 1385
2 2872 1 1388
2 2873 1 1388
2 2874 1 1392
2 2875 1 1392
2 2876 1 1393
2 2877 1 1393
2 2878 1 1396
2 2879 1 1396
2 2880 1 1399
2 2881 1 1399
2 2882 1 1400
2 2883 1 1400
2 2884 1 1404
2 2885 1 1404
2 2886 1 1407
2 2887 1 1407
2 2888 1 1408
2 2889 1 1408
2 2890 1 1412
2 2891 1 1412
2 2892 1 1415
2 2893 1 1415
2 2894 1 1416
2 2895 1 1416
2 2896 1 1420
2 2897 1 1420
2 2898 1 1423
2 2899 1 1423
2 2900 1 1424
2 2901 1 1424
2 2902 1 1428
2 2903 1 1428
2 2904 1 1431
2 2905 1 1431
2 2906 1 1432
2 2907 1 1432
2 2908 1 1436
2 2909 1 1436
2 2910 1 1439
2 2911 1 1439
2 2912 1 1440
2 2913 1 1440
2 2914 1 1444
2 2915 1 1444
2 2916 1 1447
2 2917 1 1447
2 2918 1 1448
2 2919 1 1448
2 2920 1 1452
2 2921 1 1452
2 2922 1 1455
2 2923 1 1455
2 2924 1 1456
2 2925 1 1456
2 2926 1 1458
2 2927 1 1458
2 2928 1 1461
2 2929 1 1461
2 2930 1 1464
2 2931 1 1464
2 2932 1 1467
2 2933 1 1467
2 2934 1 1470
2 2935 1 1470
2 2936 1 1473
2 2937 1 1473
2 2938 1 1476
2 2939 1 1476
2 2940 1 1479
2 2941 1 1479
2 2942 1 1482
2 2943 1 1482
2 2944 1 1488
2 2945 1 1488
2 2946 1 1494
2 2947 1 1494
2 2948 1 1502
2 2949 1 1502
2 2950 1 1510
2 2951 1 1510
2 2952 1 1514
2 2953 1 1514
2 2954 1 1522
2 2955 1 1522
2 2956 1 1526
2 2957 1 1526
2 2958 1 1532
2 2959 1 1532
2 2960 1 1533
2 2961 1 1533
2 2962 1 1538
2 2963 1 1538
2 2964 1 1546
2 2965 1 1546
2 2966 1 1554
2 2967 1 1554
2 2968 1 1574
2 2969 1 1574
2 2970 1 1586
2 2971 1 1586
2 2972 1 1601
2 2973 1 1601
2 2974 1 1625
2 2975 1 1625
2 2976 1 1628
2 2977 1 1628
2 2978 1 1631
2 2979 1 1631
0 50 5 1 1 49
0 51 5 1 1 1657
0 52 5 1 1 1659
0 53 5 1 1 1661
0 54 5 1 1 1663
0 55 5 1 1 1665
0 56 5 1 1 1667
0 57 5 1 1 1669
0 58 5 1 1 1671
0 59 5 1 1 1673
0 60 5 1 1 1675
0 61 5 1 1 1677
0 62 5 1 1 1679
0 63 5 1 1 1681
0 64 5 1 1 1683
0 65 5 1 1 1685
0 66 5 1 1 1687
0 67 5 1 1 1689
0 68 5 1 1 1691
0 69 5 2 1 1693
0 70 5 2 1 1695
0 71 5 2 1 1697
0 72 5 2 1 1699
0 73 5 2 1 1701
0 74 5 2 1 1703
0 75 5 2 1 1705
0 76 5 2 1 1707
0 77 5 2 1 1709
0 78 5 2 1 1711
0 79 5 2 1 1713
0 80 5 2 1 1715
0 81 5 2 1 1717
0 82 5 1 1 1719
0 83 5 1 1 1721
0 84 5 1 1 1723
0 85 5 1 1 1725
0 86 5 1 1 1727
0 87 5 1 1 1729
0 88 5 1 1 1731
0 89 5 1 1 1733
0 90 5 1 1 1735
0 91 5 1 1 1737
0 92 5 1 1 1739
0 93 5 1 1 1741
0 94 5 1 1 1743
0 95 5 1 1 1745
0 96 5 1 1 1747
0 97 5 1 1 1749
0 98 5 1 1 1751
0 99 7 1 2 52 68
0 100 5 2 1 99
0 101 7 1 2 1660 1692
0 102 5 2 1 101
0 103 7 1 2 51 67
0 104 5 2 1 103
0 105 7 1 2 1658 1690
0 106 5 2 1 105
0 107 7 2 2 1656 1688
0 108 5 3 1 1787
0 109 7 1 2 1785 1789
0 110 5 1 1 109
0 111 7 2 2 1783 110
0 112 5 2 1 1792
0 113 7 1 2 1781 1794
0 114 5 1 1 113
0 115 7 2 2 1779 114
0 116 5 1 1 1796
0 117 7 1 2 53 116
0 118 5 2 1 117
0 119 7 1 2 1662 1797
0 120 5 2 1 119
0 121 7 1 2 1753 1800
0 122 5 1 1 121
0 123 7 2 2 1798 122
0 124 5 1 1 1802
0 125 7 1 2 54 124
0 126 5 2 1 125
0 127 7 1 2 1664 1803
0 128 5 2 1 127
0 129 7 1 2 1755 1806
0 130 5 1 1 129
0 131 7 2 2 1804 130
0 132 5 1 1 1808
0 133 7 1 2 55 132
0 134 5 2 1 133
0 135 7 1 2 1666 1809
0 136 5 2 1 135
0 137 7 1 2 1757 1812
0 138 5 1 1 137
0 139 7 2 2 1810 138
0 140 5 1 1 1814
0 141 7 1 2 56 140
0 142 5 2 1 141
0 143 7 1 2 1668 1815
0 144 5 2 1 143
0 145 7 1 2 1759 1818
0 146 5 1 1 145
0 147 7 2 2 1816 146
0 148 5 1 1 1820
0 149 7 1 2 57 148
0 150 5 2 1 149
0 151 7 1 2 1670 1821
0 152 5 2 1 151
0 153 7 1 2 1761 1824
0 154 5 1 1 153
0 155 7 2 2 1822 154
0 156 5 1 1 1826
0 157 7 1 2 58 156
0 158 5 2 1 157
0 159 7 1 2 1672 1827
0 160 5 2 1 159
0 161 7 1 2 1763 1830
0 162 5 1 1 161
0 163 7 2 2 1828 162
0 164 5 1 1 1832
0 165 7 1 2 59 164
0 166 5 2 1 165
0 167 7 1 2 1674 1833
0 168 5 2 1 167
0 169 7 1 2 1765 1836
0 170 5 1 1 169
0 171 7 2 2 1834 170
0 172 5 1 1 1838
0 173 7 1 2 60 172
0 174 5 2 1 173
0 175 7 1 2 1676 1839
0 176 5 2 1 175
0 177 7 1 2 1767 1842
0 178 5 1 1 177
0 179 7 2 2 1840 178
0 180 5 1 1 1844
0 181 7 1 2 61 180
0 182 5 2 1 181
0 183 7 1 2 1678 1845
0 184 5 2 1 183
0 185 7 1 2 1769 1848
0 186 5 1 1 185
0 187 7 2 2 1846 186
0 188 5 1 1 1850
0 189 7 1 2 62 188
0 190 5 2 1 189
0 191 7 1 2 1680 1851
0 192 5 2 1 191
0 193 7 1 2 1771 1854
0 194 5 1 1 193
0 195 7 2 2 1852 194
0 196 5 1 1 1856
0 197 7 1 2 63 196
0 198 5 2 1 197
0 199 7 1 2 1682 1857
0 200 5 2 1 199
0 201 7 1 2 1773 1860
0 202 5 1 1 201
0 203 7 2 2 1858 202
0 204 5 1 1 1862
0 205 7 1 2 64 204
0 206 5 2 1 205
0 207 7 1 2 1684 1863
0 208 5 2 1 207
0 209 7 2 2 1864 1866
0 210 5 1 1 1868
0 211 7 1 2 1716 1869
0 212 5 1 1 211
0 213 7 1 2 1775 210
0 214 5 1 1 213
0 215 7 4 2 212 214
0 216 5 3 1 1870
0 217 7 1 2 96 1871
0 218 5 3 1 217
0 219 7 1 2 1748 1874
0 220 5 3 1 219
0 221 7 3 2 1877 1880
0 222 5 2 1 1883
0 223 7 2 2 1859 1861
0 224 5 1 1 1888
0 225 7 1 2 1714 1889
0 226 5 1 1 225
0 227 7 1 2 1774 224
0 228 5 1 1 227
0 229 7 4 2 226 228
0 230 5 3 1 1890
0 231 7 1 2 95 1891
0 232 5 3 1 231
0 233 7 1 2 1746 1894
0 234 5 3 1 233
0 235 7 2 2 1853 1855
0 236 5 1 1 1903
0 237 7 1 2 1712 1904
0 238 5 1 1 237
0 239 7 1 2 1772 236
0 240 5 1 1 239
0 241 7 4 2 238 240
0 242 5 3 1 1905
0 243 7 1 2 94 1906
0 244 5 3 1 243
0 245 7 1 2 1744 1909
0 246 5 3 1 245
0 247 7 2 2 1847 1849
0 248 5 1 1 1918
0 249 7 1 2 1710 1919
0 250 5 1 1 249
0 251 7 1 2 1770 248
0 252 5 1 1 251
0 253 7 2 2 250 252
0 254 5 3 1 1920
0 255 7 1 2 93 1921
0 256 5 3 1 255
0 257 7 1 2 1742 1922
0 258 5 3 1 257
0 259 7 2 2 1841 1843
0 260 5 1 1 1931
0 261 7 1 2 1708 1932
0 262 5 1 1 261
0 263 7 1 2 1768 260
0 264 5 1 1 263
0 265 7 4 2 262 264
0 266 5 3 1 1933
0 267 7 1 2 92 1934
0 268 5 3 1 267
0 269 7 1 2 1740 1937
0 270 5 3 1 269
0 271 7 2 2 1835 1837
0 272 5 1 1 1946
0 273 7 1 2 1706 1947
0 274 5 1 1 273
0 275 7 1 2 1766 272
0 276 5 1 1 275
0 277 7 2 2 274 276
0 278 5 3 1 1948
0 279 7 1 2 91 1949
0 280 5 3 1 279
0 281 7 1 2 1738 1950
0 282 5 3 1 281
0 283 7 2 2 1829 1831
0 284 5 1 1 1959
0 285 7 1 2 1704 1960
0 286 5 1 1 285
0 287 7 1 2 1764 284
0 288 5 1 1 287
0 289 7 4 2 286 288
0 290 5 3 1 1961
0 291 7 1 2 90 1962
0 292 5 3 1 291
0 293 7 1 2 1736 1965
0 294 5 3 1 293
0 295 7 2 2 1823 1825
0 296 5 1 1 1974
0 297 7 1 2 1702 1975
0 298 5 1 1 297
0 299 7 1 2 1762 296
0 300 5 1 1 299
0 301 7 4 2 298 300
0 302 5 3 1 1976
0 303 7 1 2 89 1977
0 304 5 3 1 303
0 305 7 1 2 1734 1980
0 306 5 3 1 305
0 307 7 2 2 1817 1819
0 308 5 1 1 1989
0 309 7 1 2 1700 1990
0 310 5 1 1 309
0 311 7 1 2 1760 308
0 312 5 1 1 311
0 313 7 4 2 310 312
0 314 5 3 1 1991
0 315 7 1 2 88 1992
0 316 5 3 1 315
0 317 7 1 2 1732 1995
0 318 5 3 1 317
0 319 7 2 2 1811 1813
0 320 5 1 1 2004
0 321 7 1 2 1698 2005
0 322 5 1 1 321
0 323 7 1 2 1758 320
0 324 5 1 1 323
0 325 7 4 2 322 324
0 326 5 3 1 2006
0 327 7 1 2 87 2007
0 328 5 3 1 327
0 329 7 1 2 1730 2010
0 330 5 3 1 329
0 331 7 2 2 1805 1807
0 332 5 1 1 2019
0 333 7 1 2 1696 2020
0 334 5 1 1 333
0 335 7 1 2 1756 332
0 336 5 1 1 335
0 337 7 3 2 334 336
0 338 5 2 1 2021
0 339 7 1 2 86 2022
0 340 5 3 1 339
0 341 7 1 2 1728 2024
0 342 5 3 1 341
0 343 7 2 2 1799 1801
0 344 5 1 1 2032
0 345 7 1 2 1694 2033
0 346 5 1 1 345
0 347 7 1 2 1754 344
0 348 5 1 1 347
0 349 7 2 2 346 348
0 350 5 2 1 2034
0 351 7 1 2 85 2035
0 352 5 3 1 351
0 353 7 1 2 1726 2036
0 354 5 3 1 353
0 355 7 2 2 1780 1782
0 356 5 1 1 2044
0 357 7 1 2 1793 356
0 358 5 1 1 357
0 359 7 1 2 1795 2045
0 360 5 1 1 359
0 361 7 2 2 358 360
0 362 5 1 1 2046
0 363 7 1 2 84 362
0 364 5 3 1 363
0 365 7 1 2 1724 2047
0 366 5 3 1 365
0 367 7 2 2 1784 1786
0 368 5 1 1 2054
0 369 7 1 2 1788 368
0 370 5 1 1 369
0 371 7 1 2 1790 2055
0 372 5 1 1 371
0 373 7 2 2 370 372
0 374 5 1 1 2056
0 375 7 1 2 83 374
0 376 5 3 1 375
0 377 7 1 2 1722 2057
0 378 5 3 1 377
0 379 7 1 2 50 66
0 380 5 1 1 379
0 381 7 2 2 1791 380
0 382 5 1 1 2064
0 383 7 3 2 82 2065
0 384 5 2 1 2066
0 385 7 1 2 2061 2067
0 386 5 1 1 385
0 387 7 2 2 2058 386
0 388 5 2 1 2071
0 389 7 1 2 2051 2073
0 390 5 1 1 389
0 391 7 2 2 2048 390
0 392 5 2 1 2075
0 393 7 1 2 2041 2077
0 394 5 1 1 393
0 395 7 2 2 2038 394
0 396 5 2 1 2079
0 397 7 1 2 2029 2081
0 398 5 1 1 397
0 399 7 2 2 2026 398
0 400 5 2 1 2083
0 401 7 1 2 2016 2085
0 402 5 1 1 401
0 403 7 2 2 2013 402
0 404 5 2 1 2087
0 405 7 1 2 2001 2089
0 406 5 1 1 405
0 407 7 2 2 1998 406
0 408 5 2 1 2091
0 409 7 1 2 1986 2093
0 410 5 1 1 409
0 411 7 2 2 1983 410
0 412 5 2 1 2095
0 413 7 1 2 1971 2097
0 414 5 1 1 413
0 415 7 2 2 1968 414
0 416 5 2 1 2099
0 417 7 1 2 1956 2101
0 418 5 1 1 417
0 419 7 2 2 1953 418
0 420 5 2 1 2103
0 421 7 1 2 1943 2105
0 422 5 1 1 421
0 423 7 2 2 1940 422
0 424 5 2 1 2107
0 425 7 1 2 1928 2109
0 426 5 1 1 425
0 427 7 2 2 1925 426
0 428 5 2 1 2111
0 429 7 1 2 1915 2113
0 430 5 1 1 429
0 431 7 2 2 1912 430
0 432 5 2 1 2115
0 433 7 1 2 1900 2117
0 434 5 1 1 433
0 435 7 2 2 1897 434
0 436 5 2 1 2119
0 437 7 1 2 1884 2120
0 438 5 1 1 437
0 439 7 1 2 1886 2121
0 440 5 1 1 439
0 441 7 4 2 438 440
0 442 5 3 1 2123
0 443 7 1 2 1776 1867
0 444 5 1 1 443
0 445 7 2 2 1865 444
0 446 5 1 1 2130
0 447 7 1 2 65 446
0 448 5 2 1 447
0 449 7 1 2 1686 2131
0 450 5 2 1 449
0 451 7 1 2 1777 2134
0 452 5 1 1 451
0 453 7 4 2 2132 452
0 454 5 3 1 2136
0 455 7 1 2 98 2137
0 456 5 4 1 455
0 457 7 1 2 1752 2140
0 458 5 4 1 457
0 459 7 2 2 2133 2135
0 460 5 1 1 2151
0 461 7 1 2 1718 460
0 462 5 1 1 461
0 463 7 1 2 1778 2152
0 464 5 1 1 463
0 465 7 4 2 462 464
0 466 5 3 1 2153
0 467 7 1 2 97 2157
0 468 5 3 1 467
0 469 7 1 2 1750 2154
0 470 5 3 1 469
0 471 7 1 2 1881 2122
0 472 5 1 1 471
0 473 7 2 2 1878 472
0 474 5 2 1 2166
0 475 7 1 2 2163 2168
0 476 5 1 1 475
0 477 7 3 2 2160 476
0 478 5 3 1 2170
0 479 7 1 2 2147 2173
0 480 5 1 1 479
0 481 7 4 2 2143 480
0 482 5 2 1 2176
0 483 7 3 2 2161 2164
0 484 5 2 1 2182
0 485 7 1 2 2167 2183
0 486 5 1 1 485
0 487 7 1 2 2169 2185
0 488 5 1 1 487
0 489 7 3 2 486 488
0 490 5 3 1 2187
0 491 7 1 2 2180 2188
0 492 5 1 1 491
0 493 7 1 2 2177 2190
0 494 5 1 1 493
0 495 7 2 2 492 494
0 496 5 1 1 2193
0 497 7 1 2 2124 2194
0 498 5 1 1 497
0 499 7 3 2 1926 1929
0 500 5 2 1 2195
0 501 7 1 2 2108 2198
0 502 5 1 1 501
0 503 7 1 2 2110 2196
0 504 5 1 1 503
0 505 7 4 2 502 504
0 506 5 3 1 2200
0 507 7 1 2 2191 2204
0 508 5 1 1 507
0 509 7 1 2 2189 2201
0 510 5 1 1 509
0 511 7 2 2 508 510
0 512 5 1 1 2207
0 513 7 3 2 1913 1916
0 514 5 2 1 2209
0 515 7 1 2 2112 2212
0 516 5 1 1 515
0 517 7 1 2 2114 2210
0 518 5 1 1 517
0 519 7 4 2 516 518
0 520 5 3 1 2214
0 521 7 1 2 512 2218
0 522 5 2 1 521
0 523 7 1 2 2208 2215
0 524 5 1 1 523
0 525 7 1 2 2221 524
0 526 5 1 1 525
0 527 7 1 2 498 526
0 528 7 1 2 2144 2174
0 529 5 1 1 528
0 530 7 1 2 2148 2171
0 531 5 1 1 530
0 532 7 1 2 529 531
0 533 7 1 2 496 532
0 534 5 1 1 533
0 535 7 3 2 1984 1987
0 536 5 2 1 2223
0 537 7 1 2 2092 2226
0 538 5 1 1 537
0 539 7 1 2 2094 2224
0 540 5 1 1 539
0 541 7 4 2 538 540
0 542 5 3 1 2228
0 543 7 1 2 2205 2232
0 544 5 2 1 543
0 545 7 1 2 2202 2229
0 546 5 1 1 545
0 547 7 2 2 2235 546
0 548 5 1 1 2237
0 549 7 3 2 1969 1972
0 550 5 2 1 2239
0 551 7 1 2 2096 2242
0 552 5 1 1 551
0 553 7 1 2 2098 2240
0 554 5 1 1 553
0 555 7 4 2 552 554
0 556 5 3 1 2244
0 557 7 1 2 2238 2248
0 558 5 2 1 557
0 559 7 2 2 2236 2251
0 560 5 1 1 2253
0 561 7 3 2 1954 1957
0 562 5 2 1 2255
0 563 7 1 2 2100 2258
0 564 5 1 1 563
0 565 7 1 2 2102 2256
0 566 5 1 1 565
0 567 7 4 2 564 566
0 568 5 3 1 2260
0 569 7 1 2 2219 2249
0 570 5 2 1 569
0 571 7 1 2 2216 2245
0 572 5 1 1 571
0 573 7 2 2 2267 572
0 574 5 1 1 2269
0 575 7 1 2 2264 2270
0 576 5 2 1 575
0 577 7 1 2 2261 574
0 578 5 1 1 577
0 579 7 2 2 2271 578
0 580 5 1 1 2273
0 581 7 1 2 560 2274
0 582 5 2 1 581
0 583 7 3 2 1941 1944
0 584 5 2 1 2277
0 585 7 1 2 2104 2280
0 586 5 1 1 585
0 587 7 1 2 2106 2278
0 588 5 1 1 587
0 589 7 4 2 586 588
0 590 5 3 1 2282
0 591 7 3 2 1999 2002
0 592 5 2 1 2289
0 593 7 1 2 2088 2292
0 594 5 1 1 593
0 595 7 1 2 2090 2290
0 596 5 1 1 595
0 597 7 4 2 594 596
0 598 5 3 1 2294
0 599 7 1 2 2286 2298
0 600 5 2 1 599
0 601 7 1 2 2283 2295
0 602 5 1 1 601
0 603 7 2 2 2301 602
0 604 5 1 1 2303
0 605 7 1 2 2304 2233
0 606 5 2 1 605
0 607 7 2 2 2302 2305
0 608 5 1 1 2307
0 609 7 1 2 548 2246
0 610 5 1 1 609
0 611 7 2 2 2252 610
0 612 5 1 1 2309
0 613 7 1 2 608 2310
0 614 5 2 1 613
0 615 7 3 2 2014 2017
0 616 5 2 1 2313
0 617 7 1 2 2084 2316
0 618 5 1 1 617
0 619 7 1 2 2086 2314
0 620 5 1 1 619
0 621 7 4 2 618 620
0 622 5 3 1 2318
0 623 7 1 2 2265 2322
0 624 5 2 1 623
0 625 7 1 2 2262 2319
0 626 5 1 1 625
0 627 7 2 2 2325 626
0 628 5 1 1 2327
0 629 7 1 2 2299 2328
0 630 5 2 1 629
0 631 7 2 2 2326 2329
0 632 5 1 1 2331
0 633 7 1 2 604 2230
0 634 5 1 1 633
0 635 7 2 2 2306 634
0 636 5 1 1 2333
0 637 7 1 2 632 2334
0 638 5 2 1 637
0 639 7 3 2 2027 2030
0 640 5 2 1 2337
0 641 7 1 2 2080 2340
0 642 5 1 1 641
0 643 7 1 2 2082 2338
0 644 5 1 1 643
0 645 7 4 2 642 644
0 646 5 3 1 2342
0 647 7 1 2 2250 2346
0 648 5 2 1 647
0 649 7 1 2 2247 2343
0 650 5 1 1 649
0 651 7 2 2 2349 650
0 652 5 1 1 2351
0 653 7 1 2 2323 2352
0 654 5 2 1 653
0 655 7 2 2 2350 2353
0 656 5 1 1 2355
0 657 7 1 2 2296 628
0 658 5 1 1 657
0 659 7 2 2 2330 658
0 660 5 1 1 2357
0 661 7 1 2 656 2358
0 662 5 2 1 661
0 663 7 3 2 2039 2042
0 664 5 2 1 2361
0 665 7 1 2 2076 2364
0 666 5 1 1 665
0 667 7 1 2 2078 2362
0 668 5 1 1 667
0 669 7 5 2 666 668
0 670 5 3 1 2366
0 671 7 1 2 2234 2371
0 672 5 2 1 671
0 673 7 1 2 2231 2367
0 674 5 1 1 673
0 675 7 2 2 2374 674
0 676 5 1 1 2376
0 677 7 1 2 2347 2377
0 678 5 2 1 677
0 679 7 2 2 2375 2378
0 680 5 1 1 2380
0 681 7 1 2 2320 652
0 682 5 1 1 681
0 683 7 2 2 2354 682
0 684 5 1 1 2382
0 685 7 1 2 680 2383
0 686 5 2 1 685
0 687 7 3 2 2049 2052
0 688 5 2 1 2386
0 689 7 1 2 2072 2389
0 690 5 1 1 689
0 691 7 1 2 2074 2387
0 692 5 1 1 691
0 693 7 4 2 690 692
0 694 5 3 1 2391
0 695 7 1 2 2300 2395
0 696 5 2 1 695
0 697 7 1 2 2297 2392
0 698 5 1 1 697
0 699 7 2 2 2398 698
0 700 5 1 1 2400
0 701 7 1 2 2372 2401
0 702 5 2 1 701
0 703 7 2 2 2399 2402
0 704 5 1 1 2404
0 705 7 1 2 2344 676
0 706 5 1 1 705
0 707 7 2 2 2379 706
0 708 5 1 1 2406
0 709 7 1 2 704 2407
0 710 5 2 1 709
0 711 7 3 2 2059 2062
0 712 5 2 1 2410
0 713 7 1 2 2068 2411
0 714 5 1 1 713
0 715 7 1 2 2069 2413
0 716 5 1 1 715
0 717 7 4 2 714 716
0 718 5 2 1 2415
0 719 7 1 2 2324 2419
0 720 5 2 1 719
0 721 7 1 2 2321 2416
0 722 5 1 1 721
0 723 7 2 2 2421 722
0 724 5 1 1 2423
0 725 7 1 2 2396 2424
0 726 5 2 1 725
0 727 7 2 2 2422 2425
0 728 5 1 1 2427
0 729 7 1 2 2368 700
0 730 5 1 1 729
0 731 7 2 2 2403 730
0 732 5 1 1 2429
0 733 7 1 2 728 2430
0 734 5 2 1 733
0 735 7 2 2 2348 2420
0 736 5 2 1 2433
0 737 7 1 2 2393 724
0 738 5 1 1 737
0 739 7 2 2 2426 738
0 740 5 1 1 2437
0 741 7 1 2 2434 2438
0 742 5 2 1 741
0 743 7 1 2 2435 740
0 744 5 1 1 743
0 745 7 2 2 2439 744
0 746 5 1 1 2441
0 747 7 2 2 1720 382
0 748 5 3 1 2443
0 749 7 3 2 2070 2445
0 750 5 5 1 2448
0 751 7 1 2 2345 2417
0 752 5 1 1 751
0 753 7 2 2 2436 752
0 754 5 2 1 2456
0 755 7 1 2 2369 2458
0 756 5 1 1 755
0 757 7 2 2 2451 756
0 758 5 1 1 2460
0 759 7 1 2 2442 2461
0 760 5 2 1 759
0 761 7 2 2 2440 2462
0 762 5 1 1 2464
0 763 7 1 2 2428 732
0 764 5 1 1 763
0 765 7 2 2 2431 764
0 766 5 1 1 2466
0 767 7 1 2 762 2467
0 768 5 2 1 767
0 769 7 2 2 2432 2468
0 770 5 1 1 2470
0 771 7 1 2 2405 708
0 772 5 1 1 771
0 773 7 2 2 2408 772
0 774 5 1 1 2472
0 775 7 1 2 770 2473
0 776 5 2 1 775
0 777 7 2 2 2409 2474
0 778 5 1 1 2476
0 779 7 1 2 2381 684
0 780 5 1 1 779
0 781 7 2 2 2384 780
0 782 5 1 1 2478
0 783 7 1 2 778 2479
0 784 5 2 1 783
0 785 7 2 2 2385 2480
0 786 5 1 1 2482
0 787 7 1 2 2356 660
0 788 5 1 1 787
0 789 7 2 2 2359 788
0 790 5 1 1 2484
0 791 7 1 2 786 2485
0 792 5 2 1 791
0 793 7 2 2 2360 2486
0 794 5 1 1 2488
0 795 7 1 2 2332 636
0 796 5 1 1 795
0 797 7 2 2 2335 796
0 798 5 1 1 2490
0 799 7 1 2 794 2491
0 800 5 2 1 799
0 801 7 2 2 2336 2492
0 802 5 1 1 2494
0 803 7 1 2 2308 612
0 804 5 1 1 803
0 805 7 2 2 2311 804
0 806 5 1 1 2496
0 807 7 1 2 802 2497
0 808 5 2 1 807
0 809 7 2 2 2312 2498
0 810 5 1 1 2500
0 811 7 1 2 2254 580
0 812 5 1 1 811
0 813 7 2 2 2275 812
0 814 5 1 1 2502
0 815 7 1 2 810 2503
0 816 5 2 1 815
0 817 7 2 2 2276 2504
0 818 5 1 1 2506
0 819 7 2 2 2268 2272
0 820 5 1 1 2508
0 821 7 3 2 1898 1901
0 822 5 2 1 2510
0 823 7 1 2 2116 2513
0 824 5 1 1 823
0 825 7 1 2 2118 2511
0 826 5 1 1 825
0 827 7 3 2 824 826
0 828 5 1 1 2515
0 829 7 1 2 2266 828
0 830 5 2 1 829
0 831 7 1 2 2263 2516
0 832 5 1 1 831
0 833 7 2 2 2518 832
0 834 5 1 1 2520
0 835 7 1 2 2287 2521
0 836 5 2 1 835
0 837 7 1 2 2284 834
0 838 5 1 1 837
0 839 7 2 2 2522 838
0 840 5 1 1 2524
0 841 7 1 2 820 2525
0 842 5 2 1 841
0 843 7 1 2 2509 840
0 844 5 1 1 843
0 845 7 2 2 2526 844
0 846 5 1 1 2528
0 847 7 1 2 818 2529
0 848 5 2 1 847
0 849 7 1 2 2507 846
0 850 5 1 1 849
0 851 7 2 2 2530 850
0 852 5 1 1 2532
0 853 7 1 2 2138 852
0 854 5 1 1 853
0 855 7 1 2 2501 814
0 856 5 1 1 855
0 857 7 2 2 2505 856
0 858 5 1 1 2534
0 859 7 1 2 2155 2535
0 860 5 1 1 859
0 861 7 1 2 2489 798
0 862 5 1 1 861
0 863 7 2 2 2493 862
0 864 5 1 1 2536
0 865 7 1 2 1892 864
0 866 5 1 1 865
0 867 7 1 2 1895 2537
0 868 5 1 1 867
0 869 7 1 2 2483 790
0 870 5 1 1 869
0 871 7 2 2 2487 870
0 872 5 1 1 2538
0 873 7 1 2 1907 872
0 874 5 1 1 873
0 875 7 1 2 1910 2539
0 876 5 1 1 875
0 877 7 1 2 2477 782
0 878 5 1 1 877
0 879 7 2 2 2481 878
0 880 5 1 1 2540
0 881 7 1 2 2471 774
0 882 5 1 1 881
0 883 7 2 2 2475 882
0 884 5 1 1 2542
0 885 7 1 2 1938 2543
0 886 5 1 1 885
0 887 7 1 2 1935 884
0 888 5 1 1 887
0 889 7 1 2 2465 766
0 890 5 1 1 889
0 891 7 2 2 2469 890
0 892 5 1 1 2544
0 893 7 1 2 746 758
0 894 5 1 1 893
0 895 7 2 2 2463 894
0 896 5 1 1 2546
0 897 7 1 2 1966 2547
0 898 5 1 1 897
0 899 7 1 2 1963 896
0 900 5 1 1 899
0 901 7 2 2 2370 2452
0 902 5 2 1 2548
0 903 7 1 2 2457 2550
0 904 5 1 1 903
0 905 7 1 2 2459 2549
0 906 5 1 1 905
0 907 7 2 2 904 906
0 908 5 1 1 2552
0 909 7 1 2 1981 908
0 910 5 1 1 909
0 911 7 1 2 1978 2553
0 912 5 1 1 911
0 913 7 1 2 2373 2449
0 914 5 1 1 913
0 915 7 2 2 2551 914
0 916 5 1 1 2554
0 917 7 1 2 1996 916
0 918 5 1 1 917
0 919 7 1 2 1993 2555
0 920 5 1 1 919
0 921 7 1 2 2011 2397
0 922 5 1 1 921
0 923 7 1 2 2008 2394
0 924 5 1 1 923
0 925 7 2 2 2037 2453
0 926 5 1 1 2556
0 927 7 1 2 2023 926
0 928 5 2 1 927
0 929 7 1 2 2025 2557
0 930 5 2 1 929
0 931 7 1 2 2418 2560
0 932 5 1 1 931
0 933 7 1 2 2558 932
0 934 7 1 2 924 933
0 935 5 1 1 934
0 936 7 1 2 922 935
0 937 5 1 1 936
0 938 7 1 2 920 937
0 939 5 1 1 938
0 940 7 1 2 918 939
0 941 5 1 1 940
0 942 7 1 2 912 941
0 943 5 1 1 942
0 944 7 1 2 910 943
0 945 5 1 1 944
0 946 7 1 2 900 945
0 947 5 1 1 946
0 948 7 2 2 898 947
0 949 5 1 1 2562
0 950 7 1 2 2545 949
0 951 5 1 1 950
0 952 7 1 2 892 2563
0 953 5 1 1 952
0 954 7 1 2 1951 953
0 955 5 1 1 954
0 956 7 1 2 951 955
0 957 5 1 1 956
0 958 7 1 2 888 957
0 959 5 1 1 958
0 960 7 2 2 886 959
0 961 5 1 1 2564
0 962 7 1 2 2541 961
0 963 5 1 1 962
0 964 7 1 2 880 2565
0 965 5 1 1 964
0 966 7 1 2 1923 965
0 967 5 1 1 966
0 968 7 1 2 963 967
0 969 7 1 2 876 968
0 970 5 1 1 969
0 971 7 1 2 874 970
0 972 5 1 1 971
0 973 7 1 2 868 972
0 974 5 1 1 973
0 975 7 2 2 866 974
0 976 5 1 1 2566
0 977 7 1 2 1875 2567
0 978 5 1 1 977
0 979 7 1 2 1872 976
0 980 5 1 1 979
0 981 7 1 2 2495 806
0 982 5 1 1 981
0 983 7 1 2 2499 982
0 984 7 1 2 980 983
0 985 5 1 1 984
0 986 7 1 2 978 985
0 987 7 1 2 860 986
0 988 5 1 1 987
0 989 7 1 2 2158 858
0 990 5 1 1 989
0 991 7 1 2 988 990
0 992 7 1 2 854 991
0 993 5 1 1 992
0 994 7 1 2 534 993
0 995 7 1 2 527 994
0 996 7 2 2 2519 2523
0 997 5 1 1 2568
0 998 7 1 2 2127 2288
0 999 5 1 1 998
0 1000 7 1 2 2125 2285
0 1001 5 1 1 1000
0 1002 7 2 2 999 1001
0 1003 5 1 1 2570
0 1004 7 1 2 2206 1003
0 1005 5 2 1 1004
0 1006 7 1 2 2203 2571
0 1007 5 1 1 1006
0 1008 7 2 2 2572 1007
0 1009 5 1 1 2574
0 1010 7 1 2 997 2575
0 1011 5 2 1 1010
0 1012 7 1 2 2569 1009
0 1013 5 1 1 1012
0 1014 7 1 2 2576 1013
0 1015 5 1 1 1014
0 1016 7 3 2 2145 2149
0 1017 5 2 1 2578
0 1018 7 1 2 2172 2581
0 1019 5 1 1 1018
0 1020 7 1 2 2175 2579
0 1021 5 1 1 1020
0 1022 7 3 2 1019 1021
0 1023 5 1 1 2583
0 1024 7 1 2 2220 1023
0 1025 5 2 1 1024
0 1026 7 1 2 2217 2584
0 1027 5 1 1 1026
0 1028 7 1 2 2586 1027
0 1029 5 1 1 1028
0 1030 7 1 2 1015 1029
0 1031 7 1 2 2141 2533
0 1032 5 1 1 1031
0 1033 7 1 2 2126 2181
0 1034 5 1 1 1033
0 1035 7 1 2 2128 2178
0 1036 5 1 1 1035
0 1037 7 1 2 1034 1036
0 1038 5 1 1 1037
0 1039 7 1 2 1032 1038
0 1040 7 1 2 1030 1039
0 1041 7 1 2 2129 2517
0 1042 7 1 2 2527 1041
0 1043 7 1 2 2192 1042
0 1044 7 1 2 2573 1043
0 1045 7 1 2 2577 1044
0 1046 7 1 2 2587 1045
0 1047 7 1 2 2179 2531
0 1048 7 1 2 2063 2446
0 1049 5 1 1 1048
0 1050 7 2 2 2060 1049
0 1051 5 2 1 2588
0 1052 7 1 2 2053 2590
0 1053 5 1 1 1052
0 1054 7 2 2 2050 1053
0 1055 5 2 1 2592
0 1056 7 1 2 2043 2594
0 1057 5 1 1 1056
0 1058 7 2 2 2040 1057
0 1059 5 2 1 2596
0 1060 7 1 2 2031 2598
0 1061 5 1 1 1060
0 1062 7 2 2 2028 1061
0 1063 5 2 1 2600
0 1064 7 1 2 2018 2602
0 1065 5 1 1 1064
0 1066 7 2 2 2015 1065
0 1067 5 2 1 2604
0 1068 7 1 2 2003 2606
0 1069 5 1 1 1068
0 1070 7 2 2 2000 1069
0 1071 5 2 1 2608
0 1072 7 1 2 1988 2610
0 1073 5 1 1 1072
0 1074 7 2 2 1985 1073
0 1075 5 2 1 2612
0 1076 7 1 2 1973 2614
0 1077 5 1 1 1076
0 1078 7 2 2 1970 1077
0 1079 5 2 1 2616
0 1080 7 1 2 1958 2618
0 1081 5 1 1 1080
0 1082 7 2 2 1955 1081
0 1083 5 2 1 2620
0 1084 7 1 2 1945 2622
0 1085 5 1 1 1084
0 1086 7 2 2 1942 1085
0 1087 5 2 1 2624
0 1088 7 1 2 1930 2626
0 1089 5 1 1 1088
0 1090 7 2 2 1927 1089
0 1091 5 2 1 2628
0 1092 7 1 2 1917 2630
0 1093 5 1 1 1092
0 1094 7 2 2 1914 1093
0 1095 5 2 1 2632
0 1096 7 1 2 1902 2634
0 1097 5 1 1 1096
0 1098 7 2 2 1899 1097
0 1099 5 2 1 2636
0 1100 7 1 2 1882 2638
0 1101 5 1 1 1100
0 1102 7 2 2 1879 1101
0 1103 5 2 1 2640
0 1104 7 1 2 2165 2642
0 1105 5 1 1 1104
0 1106 7 2 2 2162 1105
0 1107 5 2 1 2644
0 1108 7 1 2 2150 2646
0 1109 5 1 1 1108
0 1110 7 4 2 2146 1109
0 1111 5 2 1 2648
0 1112 7 1 2 2585 2649
0 1113 7 1 2 1047 1112
0 1114 7 1 2 2222 1113
0 1115 7 1 2 1046 1114
0 1116 7 1 2 1040 1115
0 1117 7 1 2 995 1116
0 1118 5 1 1 1117
0 1119 7 1 2 2580 2647
0 1120 5 1 1 1119
0 1121 7 1 2 2582 2645
0 1122 5 1 1 1121
0 1123 7 4 2 1120 1122
0 1124 5 3 1 2654
0 1125 7 1 2 2184 2641
0 1126 5 1 1 1125
0 1127 7 1 2 2186 2643
0 1128 5 1 1 1127
0 1129 7 2 2 1126 1128
0 1130 5 1 1 2661
0 1131 7 2 2 2652 2662
0 1132 5 1 1 2663
0 1133 7 1 2 2650 1130
0 1134 5 1 1 1133
0 1135 7 3 2 1132 1134
0 1136 5 2 1 2665
0 1137 7 1 2 2658 2668
0 1138 5 1 1 1137
0 1139 7 1 2 2655 2666
0 1140 5 1 1 1139
0 1141 7 1 2 1138 1140
0 1142 5 1 1 1141
0 1143 7 1 2 1887 2637
0 1144 5 1 1 1143
0 1145 7 1 2 1885 2639
0 1146 5 1 1 1145
0 1147 7 4 2 1144 1146
0 1148 5 4 1 2670
0 1149 7 1 2 2651 2671
0 1150 5 2 1 1149
0 1151 7 1 2 2653 2674
0 1152 5 1 1 1151
0 1153 7 2 2 2678 1152
0 1154 5 1 1 2680
0 1155 7 1 2 2514 2633
0 1156 5 1 1 1155
0 1157 7 1 2 2512 2635
0 1158 5 1 1 1157
0 1159 7 3 2 1156 1158
0 1160 5 3 1 2682
0 1161 7 1 2 1154 2685
0 1162 5 1 1 1161
0 1163 7 1 2 2213 2629
0 1164 5 1 1 1163
0 1165 7 1 2 2211 2631
0 1166 5 1 1 1165
0 1167 7 3 2 1164 1166
0 1168 5 4 1 2688
0 1169 7 1 2 2656 2691
0 1170 5 1 1 1169
0 1171 7 1 2 2659 2689
0 1172 5 1 1 1171
0 1173 7 2 2 1170 1172
0 1174 5 1 1 2695
0 1175 7 1 2 1162 2696
0 1176 5 1 1 1175
0 1177 7 1 2 2681 2683
0 1178 5 2 1 1177
0 1179 7 1 2 1174 2697
0 1180 5 1 1 1179
0 1181 7 1 2 1176 1180
0 1182 7 1 2 1142 1181
0 1183 7 1 2 2679 2698
0 1184 5 1 1 1183
0 1185 7 1 2 2675 2669
0 1186 5 1 1 1185
0 1187 7 1 2 2672 2667
0 1188 5 1 1 1187
0 1189 7 1 2 1186 1188
0 1190 7 1 2 1184 1189
0 1191 5 1 1 1190
0 1192 7 1 2 2227 2609
0 1193 5 1 1 1192
0 1194 7 1 2 2225 2611
0 1195 5 1 1 1194
0 1196 7 4 2 1193 1195
0 1197 5 3 1 2699
0 1198 7 1 2 2199 2625
0 1199 5 1 1 1198
0 1200 7 1 2 2197 2627
0 1201 5 1 1 1200
0 1202 7 3 2 1199 1201
0 1203 5 3 1 2706
0 1204 7 1 2 2700 2707
0 1205 5 2 1 1204
0 1206 7 1 2 2703 2709
0 1207 5 1 1 1206
0 1208 7 2 2 2712 1207
0 1209 5 1 1 2714
0 1210 7 1 2 2243 2613
0 1211 5 1 1 1210
0 1212 7 1 2 2241 2615
0 1213 5 1 1 1212
0 1214 7 4 2 1211 1213
0 1215 5 3 1 2716
0 1216 7 1 2 2715 2717
0 1217 5 2 1 1216
0 1218 7 2 2 2713 2723
0 1219 5 1 1 2725
0 1220 7 1 2 2259 2617
0 1221 5 1 1 1220
0 1222 7 1 2 2257 2619
0 1223 5 1 1 1222
0 1224 7 4 2 1221 1223
0 1225 5 3 1 2727
0 1226 7 1 2 2690 2718
0 1227 5 2 1 1226
0 1228 7 1 2 2692 2720
0 1229 5 1 1 1228
0 1230 7 2 2 2734 1229
0 1231 5 1 1 2736
0 1232 7 1 2 2728 2737
0 1233 5 2 1 1232
0 1234 7 1 2 2731 1231
0 1235 5 1 1 1234
0 1236 7 2 2 2738 1235
0 1237 5 1 1 2740
0 1238 7 1 2 1219 2741
0 1239 5 2 1 1238
0 1240 7 1 2 2281 2621
0 1241 5 1 1 1240
0 1242 7 1 2 2279 2623
0 1243 5 1 1 1242
0 1244 7 4 2 1241 1243
0 1245 5 3 1 2744
0 1246 7 1 2 2293 2605
0 1247 5 1 1 1246
0 1248 7 1 2 2291 2607
0 1249 5 1 1 1248
0 1250 7 4 2 1247 1249
0 1251 5 3 1 2751
0 1252 7 1 2 2745 2752
0 1253 5 2 1 1252
0 1254 7 1 2 2748 2755
0 1255 5 1 1 1254
0 1256 7 2 2 2758 1255
0 1257 5 1 1 2760
0 1258 7 1 2 2761 2701
0 1259 5 2 1 1258
0 1260 7 2 2 2759 2762
0 1261 5 1 1 2764
0 1262 7 1 2 1209 2721
0 1263 5 1 1 1262
0 1264 7 2 2 2724 1263
0 1265 5 1 1 2766
0 1266 7 1 2 1261 2767
0 1267 5 2 1 1266
0 1268 7 1 2 2317 2601
0 1269 5 1 1 1268
0 1270 7 1 2 2315 2603
0 1271 5 1 1 1270
0 1272 7 4 2 1269 1271
0 1273 5 3 1 2770
0 1274 7 1 2 2729 2771
0 1275 5 2 1 1274
0 1276 7 1 2 2732 2774
0 1277 5 1 1 1276
0 1278 7 2 2 2777 1277
0 1279 5 1 1 2779
0 1280 7 1 2 2753 2780
0 1281 5 2 1 1280
0 1282 7 2 2 2778 2781
0 1283 5 1 1 2783
0 1284 7 1 2 1257 2704
0 1285 5 1 1 1284
0 1286 7 2 2 2763 1285
0 1287 5 1 1 2785
0 1288 7 1 2 1283 2786
0 1289 5 2 1 1288
0 1290 7 1 2 2341 2597
0 1291 5 1 1 1290
0 1292 7 1 2 2339 2599
0 1293 5 1 1 1292
0 1294 7 4 2 1291 1293
0 1295 5 3 1 2789
0 1296 7 1 2 2719 2790
0 1297 5 2 1 1296
0 1298 7 1 2 2722 2793
0 1299 5 1 1 1298
0 1300 7 2 2 2796 1299
0 1301 5 1 1 2798
0 1302 7 1 2 2772 2799
0 1303 5 2 1 1302
0 1304 7 2 2 2797 2800
0 1305 5 1 1 2802
0 1306 7 1 2 2756 1279
0 1307 5 1 1 1306
0 1308 7 2 2 2782 1307
0 1309 5 1 1 2804
0 1310 7 1 2 1305 2805
0 1311 5 2 1 1310
0 1312 7 1 2 2365 2593
0 1313 5 1 1 1312
0 1314 7 1 2 2363 2595
0 1315 5 1 1 1314
0 1316 7 4 2 1313 1315
0 1317 5 4 1 2808
0 1318 7 1 2 2702 2809
0 1319 5 2 1 1318
0 1320 7 1 2 2705 2812
0 1321 5 1 1 1320
0 1322 7 2 2 2816 1321
0 1323 5 1 1 2818
0 1324 7 1 2 2791 2819
0 1325 5 2 1 1324
0 1326 7 2 2 2817 2820
0 1327 5 1 1 2822
0 1328 7 1 2 2775 1301
0 1329 5 1 1 1328
0 1330 7 2 2 2801 1329
0 1331 5 1 1 2824
0 1332 7 1 2 1327 2825
0 1333 5 2 1 1332
0 1334 7 1 2 2388 2591
0 1335 5 1 1 1334
0 1336 7 1 2 2390 2589
0 1337 5 1 1 1336
0 1338 7 4 2 1335 1337
0 1339 5 2 1 2828
0 1340 7 1 2 2754 2829
0 1341 5 2 1 1340
0 1342 7 1 2 2757 2832
0 1343 5 1 1 1342
0 1344 7 2 2 2834 1343
0 1345 5 1 1 2836
0 1346 7 1 2 2810 2837
0 1347 5 2 1 1346
0 1348 7 2 2 2835 2838
0 1349 5 1 1 2840
0 1350 7 1 2 2794 1323
0 1351 5 1 1 1350
0 1352 7 2 2 2821 1351
0 1353 5 1 1 2842
0 1354 7 1 2 1349 2843
0 1355 5 2 1 1354
0 1356 7 1 2 2412 2447
0 1357 5 1 1 1356
0 1358 7 1 2 2414 2444
0 1359 5 1 1 1358
0 1360 7 3 2 1357 1359
0 1361 5 3 1 2846
0 1362 7 1 2 2773 2847
0 1363 5 2 1 1362
0 1364 7 1 2 2776 2849
0 1365 5 1 1 1364
0 1366 7 2 2 2852 1365
0 1367 5 1 1 2854
0 1368 7 1 2 2830 2855
0 1369 5 2 1 1368
0 1370 7 2 2 2853 2856
0 1371 5 1 1 2858
0 1372 7 1 2 2813 1345
0 1373 5 1 1 1372
0 1374 7 2 2 2839 1373
0 1375 5 1 1 2860
0 1376 7 1 2 1371 2861
0 1377 5 2 1 1376
0 1378 7 2 2 2792 2848
0 1379 5 2 1 2864
0 1380 7 1 2 2833 1367
0 1381 5 1 1 1380
0 1382 7 2 2 2857 1381
0 1383 5 1 1 2868
0 1384 7 1 2 2865 2869
0 1385 5 2 1 1384
0 1386 7 1 2 2866 1383
0 1387 5 1 1 1386
0 1388 7 2 2 2870 1387
0 1389 5 1 1 2872
0 1390 7 1 2 2795 2850
0 1391 5 1 1 1390
0 1392 7 2 2 2867 1391
0 1393 5 2 1 2874
0 1394 7 1 2 2814 2876
0 1395 5 1 1 1394
0 1396 7 2 2 2454 1395
0 1397 5 1 1 2878
0 1398 7 1 2 2873 2879
0 1399 5 2 1 1398
0 1400 7 2 2 2871 2880
0 1401 5 1 1 2882
0 1402 7 1 2 2859 1375
0 1403 5 1 1 1402
0 1404 7 2 2 2862 1403
0 1405 5 1 1 2884
0 1406 7 1 2 1401 2885
0 1407 5 2 1 1406
0 1408 7 2 2 2863 2886
0 1409 5 1 1 2888
0 1410 7 1 2 2841 1353
0 1411 5 1 1 1410
0 1412 7 2 2 2844 1411
0 1413 5 1 1 2890
0 1414 7 1 2 1409 2891
0 1415 5 2 1 1414
0 1416 7 2 2 2845 2892
0 1417 5 1 1 2894
0 1418 7 1 2 2823 1331
0 1419 5 1 1 1418
0 1420 7 2 2 2826 1419
0 1421 5 1 1 2896
0 1422 7 1 2 1417 2897
0 1423 5 2 1 1422
0 1424 7 2 2 2827 2898
0 1425 5 1 1 2900
0 1426 7 1 2 2803 1309
0 1427 5 1 1 1426
0 1428 7 2 2 2806 1427
0 1429 5 1 1 2902
0 1430 7 1 2 1425 2903
0 1431 5 2 1 1430
0 1432 7 2 2 2807 2904
0 1433 5 1 1 2906
0 1434 7 1 2 2784 1287
0 1435 5 1 1 1434
0 1436 7 2 2 2787 1435
0 1437 5 1 1 2908
0 1438 7 1 2 1433 2909
0 1439 5 2 1 1438
0 1440 7 2 2 2788 2910
0 1441 5 1 1 2912
0 1442 7 1 2 2765 1265
0 1443 5 1 1 1442
0 1444 7 2 2 2768 1443
0 1445 5 1 1 2914
0 1446 7 1 2 1441 2915
0 1447 5 2 1 1446
0 1448 7 2 2 2769 2916
0 1449 5 1 1 2918
0 1450 7 1 2 2726 1237
0 1451 5 1 1 1450
0 1452 7 2 2 2742 1451
0 1453 5 1 1 2920
0 1454 7 1 2 1449 2921
0 1455 5 2 1 1454
0 1456 7 2 2 2743 2922
0 1457 5 1 1 2924
0 1458 7 2 2 2735 2739
0 1459 5 1 1 2926
0 1460 7 1 2 2684 2730
0 1461 5 2 1 1460
0 1462 7 1 2 2686 2733
0 1463 5 1 1 1462
0 1464 7 2 2 2928 1463
0 1465 5 1 1 2930
0 1466 7 1 2 2746 2931
0 1467 5 2 1 1466
0 1468 7 1 2 2749 1465
0 1469 5 1 1 1468
0 1470 7 2 2 2932 1469
0 1471 5 1 1 2934
0 1472 7 1 2 1459 2935
0 1473 5 2 1 1472
0 1474 7 1 2 2927 1471
0 1475 5 1 1 1474
0 1476 7 2 2 2936 1475
0 1477 5 1 1 2938
0 1478 7 1 2 1457 2939
0 1479 5 2 1 1478
0 1480 7 1 2 2925 1477
0 1481 5 1 1 1480
0 1482 7 2 2 2940 1481
0 1483 5 1 1 2942
0 1484 7 1 2 2139 1483
0 1485 5 1 1 1484
0 1486 7 1 2 2919 1453
0 1487 5 1 1 1486
0 1488 7 2 2 2923 1487
0 1489 5 1 1 2944
0 1490 7 1 2 2156 2945
0 1491 5 1 1 1490
0 1492 7 1 2 2907 1437
0 1493 5 1 1 1492
0 1494 7 2 2 2911 1493
0 1495 5 1 1 2946
0 1496 7 1 2 1893 1495
0 1497 5 1 1 1496
0 1498 7 1 2 1896 2947
0 1499 5 1 1 1498
0 1500 7 1 2 2901 1429
0 1501 5 1 1 1500
0 1502 7 2 2 2905 1501
0 1503 5 1 1 2948
0 1504 7 1 2 1908 1503
0 1505 5 1 1 1504
0 1506 7 1 2 1911 2949
0 1507 5 1 1 1506
0 1508 7 1 2 2895 1421
0 1509 5 1 1 1508
0 1510 7 2 2 2899 1509
0 1511 5 1 1 2950
0 1512 7 1 2 2889 1413
0 1513 5 1 1 1512
0 1514 7 2 2 2893 1513
0 1515 5 1 1 2952
0 1516 7 1 2 1939 2953
0 1517 5 1 1 1516
0 1518 7 1 2 1936 1515
0 1519 5 1 1 1518
0 1520 7 1 2 2883 1405
0 1521 5 1 1 1520
0 1522 7 2 2 2887 1521
0 1523 5 1 1 2954
0 1524 7 1 2 1389 1397
0 1525 5 1 1 1524
0 1526 7 2 2 2881 1525
0 1527 5 1 1 2956
0 1528 7 1 2 1967 2957
0 1529 5 1 1 1528
0 1530 7 1 2 1964 1527
0 1531 5 1 1 1530
0 1532 7 2 2 2455 2815
0 1533 5 2 1 2958
0 1534 7 1 2 2875 2960
0 1535 5 1 1 1534
0 1536 7 1 2 2877 2959
0 1537 5 1 1 1536
0 1538 7 2 2 1535 1537
0 1539 5 1 1 2962
0 1540 7 1 2 1982 1539
0 1541 5 1 1 1540
0 1542 7 1 2 1979 2963
0 1543 5 1 1 1542
0 1544 7 1 2 2450 2811
0 1545 5 1 1 1544
0 1546 7 2 2 2961 1545
0 1547 5 1 1 2964
0 1548 7 1 2 1997 1547
0 1549 5 1 1 1548
0 1550 7 1 2 1994 2965
0 1551 5 1 1 1550
0 1552 7 1 2 2561 2851
0 1553 5 1 1 1552
0 1554 7 2 2 2559 1553
0 1555 5 1 1 2966
0 1556 7 1 2 2009 1555
0 1557 5 1 1 1556
0 1558 7 1 2 2831 1557
0 1559 5 1 1 1558
0 1560 7 1 2 2012 2967
0 1561 5 1 1 1560
0 1562 7 1 2 1559 1561
0 1563 5 1 1 1562
0 1564 7 1 2 1551 1563
0 1565 5 1 1 1564
0 1566 7 1 2 1549 1565
0 1567 5 1 1 1566
0 1568 7 1 2 1543 1567
0 1569 5 1 1 1568
0 1570 7 1 2 1541 1569
0 1571 5 1 1 1570
0 1572 7 1 2 1531 1571
0 1573 5 1 1 1572
0 1574 7 2 2 1529 1573
0 1575 5 1 1 2968
0 1576 7 1 2 2955 1575
0 1577 5 1 1 1576
0 1578 7 1 2 1523 2969
0 1579 5 1 1 1578
0 1580 7 1 2 1952 1579
0 1581 5 1 1 1580
0 1582 7 1 2 1577 1581
0 1583 5 1 1 1582
0 1584 7 1 2 1519 1583
0 1585 5 1 1 1584
0 1586 7 2 2 1517 1585
0 1587 5 1 1 2970
0 1588 7 1 2 2951 1587
0 1589 5 1 1 1588
0 1590 7 1 2 1511 2971
0 1591 5 1 1 1590
0 1592 7 1 2 1924 1591
0 1593 5 1 1 1592
0 1594 7 1 2 1589 1593
0 1595 7 1 2 1507 1594
0 1596 5 1 1 1595
0 1597 7 1 2 1505 1596
0 1598 5 1 1 1597
0 1599 7 1 2 1499 1598
0 1600 5 1 1 1599
0 1601 7 2 2 1497 1600
0 1602 5 1 1 2972
0 1603 7 1 2 1876 2973
0 1604 5 1 1 1603
0 1605 7 1 2 1873 1602
0 1606 5 1 1 1605
0 1607 7 1 2 2913 1445
0 1608 5 1 1 1607
0 1609 7 1 2 2917 1608
0 1610 7 1 2 1606 1609
0 1611 5 1 1 1610
0 1612 7 1 2 1604 1611
0 1613 7 1 2 1491 1612
0 1614 5 1 1 1613
0 1615 7 1 2 2159 1489
0 1616 5 1 1 1615
0 1617 7 1 2 1614 1616
0 1618 7 1 2 1485 1617
0 1619 5 1 1 1618
0 1620 7 1 2 2687 2693
0 1621 5 1 1 1620
0 1622 7 1 2 2657 1621
0 1623 5 1 1 1622
0 1624 7 1 2 2673 2747
0 1625 5 2 1 1624
0 1626 7 1 2 2676 2750
0 1627 5 1 1 1626
0 1628 7 2 2 2974 1627
0 1629 5 1 1 2976
0 1630 7 1 2 2708 2977
0 1631 5 2 1 1630
0 1632 7 1 2 2694 2710
0 1633 7 1 2 2929 1632
0 1634 7 1 2 2677 1633
0 1635 7 1 2 2933 1634
0 1636 7 1 2 2975 1635
0 1637 7 1 2 2937 1636
0 1638 7 1 2 2978 1637
0 1639 7 1 2 2664 1638
0 1640 7 1 2 1623 1639
0 1641 7 1 2 2142 2943
0 1642 5 1 1 1641
0 1643 7 1 2 2711 1629
0 1644 5 1 1 1643
0 1645 7 1 2 2979 1644
0 1646 5 1 1 1645
0 1647 7 1 2 2660 2941
0 1648 7 1 2 1646 1647
0 1649 7 1 2 1642 1648
0 1650 7 1 2 1640 1649
0 1651 7 1 2 1619 1650
0 1652 7 1 2 1191 1651
0 1653 7 1 2 1182 1652
0 1654 5 1 1 1653
0 1655 7 1 2 1118 1654
3 3499 5 0 1 1655
