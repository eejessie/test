1 0 0 2 0
2 32 1 0
2 33 1 0
1 1 0 2 0
2 34 1 1
2 35 1 1
1 2 0 2 0
2 36 1 2
2 37 1 2
1 3 0 2 0
2 38 1 3
2 39 1 3
1 4 0 2 0
2 40 1 4
2 41 1 4
1 5 0 2 0
2 42 1 5
2 43 1 5
1 6 0 2 0
2 44 1 6
2 45 1 6
1 7 0 2 0
2 46 1 7
2 47 1 7
1 8 0 2 0
2 48 1 8
2 85 1 8
1 9 0 2 0
2 96 1 9
2 109 1 9
1 10 0 2 0
2 126 1 10
2 146 1 10
1 11 0 2 0
2 166 1 11
2 189 1 11
1 12 0 2 0
2 213 1 12
2 238 1 12
1 13 0 2 0
2 263 1 13
2 288 1 13
1 14 0 2 0
2 313 1 14
2 341 1 14
1 15 0 2 0
2 369 1 15
2 397 1 15
1 16 0 2 0
2 424 1 16
2 442 1 16
1 17 0 2 0
2 443 1 17
2 444 1 17
1 18 0 2 0
2 445 1 18
2 446 1 18
1 19 0 2 0
2 447 1 19
2 448 1 19
1 20 0 2 0
2 449 1 20
2 450 1 20
1 21 0 2 0
2 451 1 21
2 452 1 21
1 22 0 2 0
2 453 1 22
2 454 1 22
1 23 0 2 0
2 455 1 23
2 456 1 23
1 24 0 2 0
2 457 1 24
2 458 1 24
1 25 0 2 0
2 459 1 25
2 460 1 25
1 26 0 2 0
2 461 1 26
2 462 1 26
1 27 0 2 0
2 463 1 27
2 464 1 27
1 28 0 2 0
2 465 1 28
2 466 1 28
1 29 0 2 0
2 467 1 29
2 468 1 29
1 30 0 2 0
2 469 1 30
2 470 1 30
1 31 0 2 0
2 471 1 31
2 472 1 31
2 473 1 81
2 474 1 81
2 475 1 82
2 476 1 82
2 477 1 87
2 478 1 87
2 479 1 87
2 480 1 90
2 481 1 90
2 482 1 93
2 483 1 93
2 484 1 93
2 485 1 97
2 486 1 97
2 487 1 98
2 488 1 98
2 489 1 100
2 490 1 100
2 491 1 100
2 492 1 102
2 493 1 102
2 494 1 103
2 495 1 103
2 496 1 103
2 497 1 111
2 498 1 111
2 499 1 111
2 500 1 113
2 501 1 113
2 502 1 114
2 503 1 114
2 504 1 114
2 505 1 114
2 506 1 119
2 507 1 119
2 508 1 119
2 509 1 119
2 510 1 128
2 511 1 128
2 512 1 132
2 513 1 132
2 514 1 134
2 515 1 134
2 516 1 135
2 517 1 135
2 518 1 137
2 519 1 137
2 520 1 137
2 521 1 139
2 522 1 139
2 523 1 140
2 524 1 140
2 525 1 140
2 526 1 140
2 527 1 148
2 528 1 148
2 529 1 148
2 530 1 150
2 531 1 150
2 532 1 151
2 533 1 151
2 534 1 151
2 535 1 151
2 536 1 153
2 537 1 153
2 538 1 158
2 539 1 158
2 540 1 160
2 541 1 160
2 542 1 161
2 543 1 161
2 544 1 161
2 545 1 167
2 546 1 167
2 547 1 167
2 548 1 174
2 549 1 174
2 550 1 177
2 551 1 177
2 552 1 178
2 553 1 178
2 554 1 178
2 555 1 180
2 556 1 180
2 557 1 180
2 558 1 182
2 559 1 182
2 560 1 183
2 561 1 183
2 562 1 183
2 563 1 183
2 564 1 190
2 565 1 190
2 566 1 190
2 567 1 198
2 568 1 198
2 569 1 201
2 570 1 201
2 571 1 202
2 572 1 202
2 573 1 202
2 574 1 204
2 575 1 204
2 576 1 204
2 577 1 206
2 578 1 206
2 579 1 207
2 580 1 207
2 581 1 207
2 582 1 207
2 583 1 214
2 584 1 214
2 585 1 214
2 586 1 219
2 587 1 219
2 588 1 221
2 589 1 221
2 590 1 224
2 591 1 224
2 592 1 226
2 593 1 226
2 594 1 227
2 595 1 227
2 596 1 229
2 597 1 229
2 598 1 229
2 599 1 231
2 600 1 231
2 601 1 232
2 602 1 232
2 603 1 232
2 604 1 232
2 605 1 239
2 606 1 239
2 607 1 239
2 608 1 244
2 609 1 244
2 610 1 246
2 611 1 246
2 612 1 248
2 613 1 248
2 614 1 251
2 615 1 251
2 616 1 254
2 617 1 254
2 618 1 254
2 619 1 256
2 620 1 256
2 621 1 257
2 622 1 257
2 623 1 257
2 624 1 257
2 625 1 264
2 626 1 264
2 627 1 264
2 628 1 269
2 629 1 269
2 630 1 271
2 631 1 271
2 632 1 273
2 633 1 273
2 634 1 276
2 635 1 276
2 636 1 279
2 637 1 279
2 638 1 279
2 639 1 281
2 640 1 281
2 641 1 282
2 642 1 282
2 643 1 282
2 644 1 282
2 645 1 289
2 646 1 289
2 647 1 289
2 648 1 294
2 649 1 294
2 650 1 296
2 651 1 296
2 652 1 298
2 653 1 298
2 654 1 301
2 655 1 301
2 656 1 304
2 657 1 304
2 658 1 304
2 659 1 306
2 660 1 306
2 661 1 307
2 662 1 307
2 663 1 307
2 664 1 307
2 665 1 314
2 666 1 314
2 667 1 314
2 668 1 315
2 669 1 315
2 670 1 315
2 671 1 322
2 672 1 322
2 673 1 324
2 674 1 324
2 675 1 329
2 676 1 329
2 677 1 332
2 678 1 332
2 679 1 332
2 680 1 334
2 681 1 334
2 682 1 335
2 683 1 335
2 684 1 335
2 685 1 335
2 686 1 342
2 687 1 342
2 688 1 342
2 689 1 343
2 690 1 343
2 691 1 353
2 692 1 353
2 693 1 357
2 694 1 357
2 695 1 359
2 696 1 359
2 697 1 360
2 698 1 360
2 699 1 362
2 700 1 362
2 701 1 363
2 702 1 363
2 703 1 363
2 704 1 363
2 705 1 370
2 706 1 370
2 707 1 370
2 708 1 370
2 709 1 371
2 710 1 371
2 711 1 382
2 712 1 382
2 713 1 385
2 714 1 385
2 715 1 388
2 716 1 388
2 717 1 388
2 718 1 390
2 719 1 390
2 720 1 390
2 721 1 391
2 722 1 391
2 723 1 391
2 724 1 391
2 725 1 398
2 726 1 398
2 727 1 399
2 728 1 399
2 729 1 412
2 730 1 412
2 731 1 415
2 732 1 415
2 733 1 417
2 734 1 417
2 735 1 418
2 736 1 418
2 737 1 418
0 49 5 1 1 32
0 50 5 1 1 34
0 51 5 1 1 36
0 52 5 1 1 38
0 53 5 1 1 40
0 54 5 1 1 42
0 55 5 1 1 44
0 56 5 1 1 46
0 57 5 1 1 48
0 58 5 1 1 96
0 59 5 1 1 126
0 60 5 1 1 166
0 61 5 1 1 213
0 62 5 1 1 263
0 63 5 1 1 313
0 64 5 1 1 369
0 65 5 1 1 424
0 66 5 1 1 443
0 67 5 1 1 445
0 68 5 1 1 447
0 69 5 1 1 449
0 70 5 1 1 451
0 71 5 1 1 453
0 72 5 1 1 455
0 73 5 1 1 457
0 74 5 1 1 459
0 75 5 1 1 461
0 76 5 1 1 463
0 77 5 1 1 465
0 78 5 1 1 467
0 79 5 1 1 469
0 80 5 1 1 471
0 81 7 2 2 33 442
0 82 5 2 1 473
0 83 7 1 2 49 65
0 84 5 1 1 83
3 883 7 0 2 475 84
0 86 7 1 2 35 444
0 87 5 3 1 86
0 88 7 1 2 50 66
0 89 5 1 1 88
0 90 7 2 2 477 89
0 91 5 1 1 480
0 92 7 1 2 474 481
0 93 5 3 1 92
0 94 7 1 2 476 91
0 95 5 1 1 94
3 884 7 0 2 482 95
0 97 7 2 2 478 483
0 98 5 2 1 485
0 99 7 1 2 37 446
0 100 5 3 1 99
0 101 7 1 2 51 67
0 102 5 2 1 101
0 103 7 3 2 489 492
0 104 5 1 1 494
0 105 7 1 2 486 104
0 106 5 1 1 105
0 107 7 1 2 487 495
0 108 5 1 1 107
3 885 7 0 2 106 108
0 110 7 1 2 39 448
0 111 5 3 1 110
0 112 7 1 2 52 68
0 113 5 2 1 112
0 114 7 4 2 497 500
0 115 5 1 1 502
0 116 7 1 2 479 490
0 117 7 1 2 484 116
0 118 5 1 1 117
0 119 7 4 2 493 118
0 120 5 1 1 506
0 121 7 1 2 503 120
0 122 5 1 1 121
0 123 7 1 2 115 507
0 124 5 1 1 123
0 125 7 1 2 122 124
3 886 5 0 1 125
0 127 7 1 2 496 504
0 128 7 2 2 488 127
0 129 5 1 1 510
0 130 7 1 2 491 498
0 131 5 1 1 130
0 132 7 2 2 501 131
0 133 5 1 1 512
0 134 7 2 2 129 133
0 135 5 2 1 514
0 136 7 1 2 41 450
0 137 5 3 1 136
0 138 7 1 2 53 69
0 139 5 2 1 138
0 140 7 4 2 518 521
0 141 5 1 1 523
0 142 7 1 2 516 524
0 143 5 1 1 142
0 144 7 1 2 515 141
0 145 5 1 1 144
3 887 7 0 2 143 145
0 147 7 1 2 43 452
0 148 5 3 1 147
0 149 7 1 2 54 70
0 150 5 2 1 149
0 151 7 4 2 527 530
0 152 5 1 1 532
0 153 7 2 2 505 525
0 154 7 1 2 508 536
0 155 5 1 1 154
0 156 7 1 2 499 519
0 157 5 1 1 156
0 158 7 2 2 522 157
0 159 5 1 1 538
0 160 7 2 2 155 159
0 161 5 3 1 540
0 162 7 1 2 533 542
0 163 5 1 1 162
0 164 7 1 2 152 541
0 165 5 1 1 164
3 888 7 0 2 163 165
0 167 7 3 2 526 534
0 168 7 1 2 511 545
0 169 5 1 1 168
0 170 7 1 2 513 546
0 171 5 1 1 170
0 172 7 1 2 520 528
0 173 5 1 1 172
0 174 7 2 2 531 173
0 175 5 1 1 548
0 176 7 1 2 171 175
0 177 7 2 2 169 176
0 178 5 3 1 550
0 179 7 1 2 45 454
0 180 5 3 1 179
0 181 7 1 2 55 71
0 182 5 2 1 181
0 183 7 4 2 555 558
0 184 5 1 1 560
0 185 7 1 2 552 561
0 186 5 1 1 185
0 187 7 1 2 551 184
0 188 5 1 1 187
3 889 7 0 2 186 188
0 190 7 3 2 535 562
0 191 7 1 2 537 564
0 192 7 1 2 509 191
0 193 5 1 1 192
0 194 7 1 2 539 565
0 195 5 1 1 194
0 196 7 1 2 529 556
0 197 5 1 1 196
0 198 7 2 2 559 197
0 199 5 1 1 567
0 200 7 1 2 195 199
0 201 7 2 2 193 200
0 202 5 3 1 569
0 203 7 1 2 47 456
0 204 5 3 1 203
0 205 7 1 2 56 72
0 206 5 2 1 205
0 207 7 4 2 574 577
0 208 5 1 1 579
0 209 7 1 2 571 580
0 210 5 1 1 209
0 211 7 1 2 570 208
0 212 5 1 1 211
3 890 7 0 2 210 212
0 214 7 3 2 563 581
0 215 7 1 2 549 583
0 216 5 1 1 215
0 217 7 1 2 557 575
0 218 5 1 1 217
0 219 7 2 2 578 218
0 220 5 1 1 586
0 221 7 2 2 216 220
0 222 5 1 1 588
0 223 7 1 2 547 584
0 224 7 2 2 517 223
0 225 5 1 1 590
0 226 7 2 2 589 225
0 227 5 2 1 592
0 228 7 1 2 85 458
0 229 5 3 1 228
0 230 7 1 2 57 73
0 231 5 2 1 230
0 232 7 4 2 596 599
0 233 5 1 1 601
0 234 7 1 2 594 602
0 235 5 1 1 234
0 236 7 1 2 593 233
0 237 5 1 1 236
3 891 7 0 2 235 237
0 239 7 3 2 582 603
0 240 7 1 2 568 605
0 241 5 1 1 240
0 242 7 1 2 576 597
0 243 5 1 1 242
0 244 7 2 2 600 243
0 245 5 1 1 608
0 246 7 2 2 241 245
0 247 5 1 1 610
0 248 7 2 2 566 606
0 249 7 1 2 543 612
0 250 5 1 1 249
0 251 7 2 2 611 250
0 252 5 1 1 614
0 253 7 1 2 109 460
0 254 5 3 1 253
0 255 7 1 2 58 74
0 256 5 2 1 255
0 257 7 4 2 616 619
0 258 5 1 1 621
0 259 7 1 2 252 622
0 260 5 1 1 259
0 261 7 1 2 615 258
0 262 5 1 1 261
3 892 7 0 2 260 262
0 264 7 3 2 604 623
0 265 7 1 2 587 625
0 266 5 1 1 265
0 267 7 1 2 598 617
0 268 5 1 1 267
0 269 7 2 2 620 268
0 270 5 1 1 628
0 271 7 2 2 266 270
0 272 5 1 1 630
0 273 7 2 2 585 626
0 274 7 1 2 553 632
0 275 5 1 1 274
0 276 7 2 2 631 275
0 277 5 1 1 634
0 278 7 1 2 146 462
0 279 5 3 1 278
0 280 7 1 2 59 75
0 281 5 2 1 280
0 282 7 4 2 636 639
0 283 5 1 1 641
0 284 7 1 2 277 642
0 285 5 1 1 284
0 286 7 1 2 635 283
0 287 5 1 1 286
3 893 7 0 2 285 287
0 289 7 3 2 624 643
0 290 7 1 2 609 645
0 291 5 1 1 290
0 292 7 1 2 618 637
0 293 5 1 1 292
0 294 7 2 2 640 293
0 295 5 1 1 648
0 296 7 2 2 291 295
0 297 5 1 1 650
0 298 7 2 2 607 646
0 299 7 1 2 572 652
0 300 5 1 1 299
0 301 7 2 2 651 300
0 302 5 1 1 654
0 303 7 1 2 189 464
0 304 5 3 1 303
0 305 7 1 2 60 76
0 306 5 2 1 305
0 307 7 4 2 656 659
0 308 5 1 1 661
0 309 7 1 2 302 662
0 310 5 1 1 309
0 311 7 1 2 655 308
0 312 5 1 1 311
3 894 7 0 2 310 312
0 314 7 3 2 644 663
0 315 7 3 2 627 665
0 316 7 1 2 591 668
0 317 5 1 1 316
0 318 7 1 2 629 666
0 319 5 1 1 318
0 320 7 1 2 638 657
0 321 5 1 1 320
0 322 7 2 2 660 321
0 323 5 1 1 671
0 324 7 2 2 319 323
0 325 5 1 1 673
0 326 7 1 2 222 669
0 327 5 1 1 326
0 328 7 1 2 674 327
0 329 7 2 2 317 328
0 330 5 1 1 675
0 331 7 1 2 238 466
0 332 5 3 1 331
0 333 7 1 2 61 77
0 334 5 2 1 333
0 335 7 4 2 677 680
0 336 5 1 1 682
0 337 7 1 2 330 683
0 338 5 1 1 337
0 339 7 1 2 676 336
0 340 5 1 1 339
3 895 7 0 2 338 340
0 342 7 3 2 664 684
0 343 7 2 2 647 686
0 344 7 1 2 613 689
0 345 7 1 2 544 344
0 346 5 1 1 345
0 347 7 1 2 247 690
0 348 5 1 1 347
0 349 7 1 2 649 687
0 350 5 1 1 349
0 351 7 1 2 658 678
0 352 5 1 1 351
0 353 7 2 2 681 352
0 354 5 1 1 691
0 355 7 1 2 350 354
0 356 7 1 2 348 355
0 357 7 2 2 346 356
0 358 5 1 1 693
0 359 7 2 2 288 468
0 360 5 2 1 695
0 361 7 1 2 62 78
0 362 5 2 1 361
0 363 7 4 2 697 699
0 364 5 1 1 701
0 365 7 1 2 358 702
0 366 5 1 1 365
0 367 7 1 2 694 364
0 368 5 1 1 367
3 896 7 0 2 366 368
0 370 7 4 2 685 703
0 371 7 2 2 667 705
0 372 7 1 2 633 709
0 373 7 1 2 554 372
0 374 5 1 1 373
0 375 7 1 2 272 710
0 376 5 1 1 375
0 377 7 1 2 672 706
0 378 5 1 1 377
0 379 7 1 2 679 698
0 380 5 1 1 379
0 381 7 1 2 700 380
0 382 5 2 1 381
0 383 7 1 2 378 711
0 384 7 1 2 376 383
0 385 7 2 2 374 384
0 386 5 1 1 713
0 387 7 1 2 341 470
0 388 5 3 1 387
0 389 7 1 2 63 79
0 390 5 3 1 389
0 391 7 4 2 715 718
0 392 5 1 1 721
0 393 7 1 2 386 722
0 394 5 1 1 393
0 395 7 1 2 714 392
0 396 5 1 1 395
3 897 7 0 2 394 396
0 398 7 2 2 704 723
0 399 7 2 2 688 725
0 400 7 1 2 653 727
0 401 7 1 2 573 400
0 402 5 1 1 401
0 403 7 1 2 297 728
0 404 5 1 1 403
0 405 7 1 2 692 726
0 406 5 1 1 405
0 407 7 1 2 696 719
0 408 5 1 1 407
0 409 7 1 2 716 408
0 410 7 1 2 406 409
0 411 7 1 2 404 410
0 412 7 2 2 402 411
0 413 5 1 1 729
0 414 7 1 2 397 472
0 415 5 2 1 414
0 416 7 1 2 64 80
0 417 5 2 1 416
0 418 7 3 2 731 733
0 419 5 1 1 735
0 420 7 1 2 413 736
0 421 5 1 1 420
0 422 7 1 2 730 419
0 423 5 1 1 422
3 898 7 0 2 421 423
0 425 7 1 2 325 707
0 426 5 1 1 425
0 427 7 1 2 712 426
0 428 5 1 1 427
0 429 7 1 2 720 428
0 430 5 1 1 429
0 431 7 1 2 717 732
0 432 7 1 2 430 431
0 433 5 1 1 432
0 434 7 1 2 734 433
0 435 5 1 1 434
0 436 7 1 2 724 737
0 437 7 1 2 708 436
0 438 7 1 2 670 437
0 439 7 1 2 595 438
0 440 5 1 1 439
0 441 7 1 2 435 440
3 899 5 0 1 441
