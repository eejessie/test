1 0 0 150 0
2 25 1 0
2 26 1 0
2 41958 1 0
2 41959 1 0
2 41960 1 0
2 41961 1 0
2 41962 1 0
2 41963 1 0
2 41964 1 0
2 41965 1 0
2 41966 1 0
2 41967 1 0
2 41968 1 0
2 41969 1 0
2 41970 1 0
2 41971 1 0
2 41972 1 0
2 41973 1 0
2 41974 1 0
2 41975 1 0
2 41976 1 0
2 41977 1 0
2 41978 1 0
2 41979 1 0
2 41980 1 0
2 41981 1 0
2 41982 1 0
2 41983 1 0
2 41984 1 0
2 41985 1 0
2 41986 1 0
2 41987 1 0
2 41988 1 0
2 41989 1 0
2 41990 1 0
2 41991 1 0
2 41992 1 0
2 41993 1 0
2 41994 1 0
2 41995 1 0
2 41996 1 0
2 41997 1 0
2 41998 1 0
2 41999 1 0
2 42000 1 0
2 42001 1 0
2 42002 1 0
2 42003 1 0
2 42004 1 0
2 42005 1 0
2 42006 1 0
2 42007 1 0
2 42008 1 0
2 42009 1 0
2 42010 1 0
2 42011 1 0
2 42012 1 0
2 42013 1 0
2 42014 1 0
2 42015 1 0
2 42016 1 0
2 42017 1 0
2 42018 1 0
2 42019 1 0
2 42020 1 0
2 42021 1 0
2 42022 1 0
2 42023 1 0
2 42024 1 0
2 42025 1 0
2 42026 1 0
2 42027 1 0
2 42028 1 0
2 42029 1 0
2 42030 1 0
2 42031 1 0
2 42032 1 0
2 42033 1 0
2 42034 1 0
2 42035 1 0
2 42036 1 0
2 42037 1 0
2 42038 1 0
2 42039 1 0
2 42040 1 0
2 42041 1 0
2 42042 1 0
2 42043 1 0
2 42044 1 0
2 42045 1 0
2 42046 1 0
2 42047 1 0
2 42048 1 0
2 42049 1 0
2 42050 1 0
2 42051 1 0
2 42052 1 0
2 42053 1 0
2 42054 1 0
2 42055 1 0
2 42056 1 0
2 42057 1 0
2 42058 1 0
2 42059 1 0
2 42060 1 0
2 42061 1 0
2 42062 1 0
2 42063 1 0
2 42064 1 0
2 42065 1 0
2 42066 1 0
2 42067 1 0
2 42068 1 0
2 42069 1 0
2 42070 1 0
2 42071 1 0
2 42072 1 0
2 42073 1 0
2 42074 1 0
2 42075 1 0
2 42076 1 0
2 42077 1 0
2 42078 1 0
2 42079 1 0
2 42080 1 0
2 42081 1 0
2 42082 1 0
2 42083 1 0
2 42084 1 0
2 42085 1 0
2 42086 1 0
2 42087 1 0
2 42088 1 0
2 42089 1 0
2 42090 1 0
2 42091 1 0
2 42092 1 0
2 42093 1 0
2 42094 1 0
2 42095 1 0
2 42096 1 0
2 42097 1 0
2 42098 1 0
2 42099 1 0
2 42100 1 0
2 42101 1 0
2 42102 1 0
2 42103 1 0
2 42104 1 0
2 42105 1 0
1 1 0 146 0
2 42106 1 1
2 42107 1 1
2 42108 1 1
2 42109 1 1
2 42110 1 1
2 42111 1 1
2 42112 1 1
2 42113 1 1
2 42114 1 1
2 42115 1 1
2 42116 1 1
2 42117 1 1
2 42118 1 1
2 42119 1 1
2 42120 1 1
2 42121 1 1
2 42122 1 1
2 42123 1 1
2 42124 1 1
2 42125 1 1
2 42126 1 1
2 42127 1 1
2 42128 1 1
2 42129 1 1
2 42130 1 1
2 42131 1 1
2 42132 1 1
2 42133 1 1
2 42134 1 1
2 42135 1 1
2 42136 1 1
2 42137 1 1
2 42138 1 1
2 42139 1 1
2 42140 1 1
2 42141 1 1
2 42142 1 1
2 42143 1 1
2 42144 1 1
2 42145 1 1
2 42146 1 1
2 42147 1 1
2 42148 1 1
2 42149 1 1
2 42150 1 1
2 42151 1 1
2 42152 1 1
2 42153 1 1
2 42154 1 1
2 42155 1 1
2 42156 1 1
2 42157 1 1
2 42158 1 1
2 42159 1 1
2 42160 1 1
2 42161 1 1
2 42162 1 1
2 42163 1 1
2 42164 1 1
2 42165 1 1
2 42166 1 1
2 42167 1 1
2 42168 1 1
2 42169 1 1
2 42170 1 1
2 42171 1 1
2 42172 1 1
2 42173 1 1
2 42174 1 1
2 42175 1 1
2 42176 1 1
2 42177 1 1
2 42178 1 1
2 42179 1 1
2 42180 1 1
2 42181 1 1
2 42182 1 1
2 42183 1 1
2 42184 1 1
2 42185 1 1
2 42186 1 1
2 42187 1 1
2 42188 1 1
2 42189 1 1
2 42190 1 1
2 42191 1 1
2 42192 1 1
2 42193 1 1
2 42194 1 1
2 42195 1 1
2 42196 1 1
2 42197 1 1
2 42198 1 1
2 42199 1 1
2 42200 1 1
2 42201 1 1
2 42202 1 1
2 42203 1 1
2 42204 1 1
2 42205 1 1
2 42206 1 1
2 42207 1 1
2 42208 1 1
2 42209 1 1
2 42210 1 1
2 42211 1 1
2 42212 1 1
2 42213 1 1
2 42214 1 1
2 42215 1 1
2 42216 1 1
2 42217 1 1
2 42218 1 1
2 42219 1 1
2 42220 1 1
2 42221 1 1
2 42222 1 1
2 42223 1 1
2 42224 1 1
2 42225 1 1
2 42226 1 1
2 42227 1 1
2 42228 1 1
2 42229 1 1
2 42230 1 1
2 42231 1 1
2 42232 1 1
2 42233 1 1
2 42234 1 1
2 42235 1 1
2 42236 1 1
2 42237 1 1
2 42238 1 1
2 42239 1 1
2 42240 1 1
2 42241 1 1
2 42242 1 1
2 42243 1 1
2 42244 1 1
2 42245 1 1
2 42246 1 1
2 42247 1 1
2 42248 1 1
2 42249 1 1
2 42250 1 1
2 42251 1 1
1 2 0 109 0
2 42252 1 2
2 42253 1 2
2 42254 1 2
2 42255 1 2
2 42256 1 2
2 42257 1 2
2 42258 1 2
2 42259 1 2
2 42260 1 2
2 42261 1 2
2 42262 1 2
2 42263 1 2
2 42264 1 2
2 42265 1 2
2 42266 1 2
2 42267 1 2
2 42268 1 2
2 42269 1 2
2 42270 1 2
2 42271 1 2
2 42272 1 2
2 42273 1 2
2 42274 1 2
2 42275 1 2
2 42276 1 2
2 42277 1 2
2 42278 1 2
2 42279 1 2
2 42280 1 2
2 42281 1 2
2 42282 1 2
2 42283 1 2
2 42284 1 2
2 42285 1 2
2 42286 1 2
2 42287 1 2
2 42288 1 2
2 42289 1 2
2 42290 1 2
2 42291 1 2
2 42292 1 2
2 42293 1 2
2 42294 1 2
2 42295 1 2
2 42296 1 2
2 42297 1 2
2 42298 1 2
2 42299 1 2
2 42300 1 2
2 42301 1 2
2 42302 1 2
2 42303 1 2
2 42304 1 2
2 42305 1 2
2 42306 1 2
2 42307 1 2
2 42308 1 2
2 42309 1 2
2 42310 1 2
2 42311 1 2
2 42312 1 2
2 42313 1 2
2 42314 1 2
2 42315 1 2
2 42316 1 2
2 42317 1 2
2 42318 1 2
2 42319 1 2
2 42320 1 2
2 42321 1 2
2 42322 1 2
2 42323 1 2
2 42324 1 2
2 42325 1 2
2 42326 1 2
2 42327 1 2
2 42328 1 2
2 42329 1 2
2 42330 1 2
2 42331 1 2
2 42332 1 2
2 42333 1 2
2 42334 1 2
2 42335 1 2
2 42336 1 2
2 42337 1 2
2 42338 1 2
2 42339 1 2
2 42340 1 2
2 42341 1 2
2 42342 1 2
2 42343 1 2
2 42344 1 2
2 42345 1 2
2 42346 1 2
2 42347 1 2
2 42348 1 2
2 42349 1 2
2 42350 1 2
2 42351 1 2
2 42352 1 2
2 42353 1 2
2 42354 1 2
2 42355 1 2
2 42356 1 2
2 42357 1 2
2 42358 1 2
2 42359 1 2
2 42360 1 2
1 3 0 49 0
2 42361 1 3
2 42362 1 3
2 42363 1 3
2 42364 1 3
2 42365 1 3
2 42366 1 3
2 42367 1 3
2 42368 1 3
2 42369 1 3
2 42370 1 3
2 42371 1 3
2 42372 1 3
2 42373 1 3
2 42374 1 3
2 42375 1 3
2 42376 1 3
2 42377 1 3
2 42378 1 3
2 42379 1 3
2 42380 1 3
2 42381 1 3
2 42382 1 3
2 42383 1 3
2 42384 1 3
2 42385 1 3
2 42386 1 3
2 42387 1 3
2 42388 1 3
2 42389 1 3
2 42390 1 3
2 42391 1 3
2 42392 1 3
2 42393 1 3
2 42394 1 3
2 42395 1 3
2 42396 1 3
2 42397 1 3
2 42398 1 3
2 42399 1 3
2 42400 1 3
2 42401 1 3
2 42402 1 3
2 42403 1 3
2 42404 1 3
2 42405 1 3
2 42406 1 3
2 42407 1 3
2 42408 1 3
2 42409 1 3
1 4 0 230 0
2 42410 1 4
2 42411 1 4
2 42412 1 4
2 42413 1 4
2 42414 1 4
2 42415 1 4
2 42416 1 4
2 42417 1 4
2 42418 1 4
2 42419 1 4
2 42420 1 4
2 42421 1 4
2 42422 1 4
2 42423 1 4
2 42424 1 4
2 42425 1 4
2 42426 1 4
2 42427 1 4
2 42428 1 4
2 42429 1 4
2 42430 1 4
2 42431 1 4
2 42432 1 4
2 42433 1 4
2 42434 1 4
2 42435 1 4
2 42436 1 4
2 42437 1 4
2 42438 1 4
2 42439 1 4
2 42440 1 4
2 42441 1 4
2 42442 1 4
2 42443 1 4
2 42444 1 4
2 42445 1 4
2 42446 1 4
2 42447 1 4
2 42448 1 4
2 42449 1 4
2 42450 1 4
2 42451 1 4
2 42452 1 4
2 42453 1 4
2 42454 1 4
2 42455 1 4
2 42456 1 4
2 42457 1 4
2 42458 1 4
2 42459 1 4
2 42460 1 4
2 42461 1 4
2 42462 1 4
2 42463 1 4
2 42464 1 4
2 42465 1 4
2 42466 1 4
2 42467 1 4
2 42468 1 4
2 42469 1 4
2 42470 1 4
2 42471 1 4
2 42472 1 4
2 42473 1 4
2 42474 1 4
2 42475 1 4
2 42476 1 4
2 42477 1 4
2 42478 1 4
2 42479 1 4
2 42480 1 4
2 42481 1 4
2 42482 1 4
2 42483 1 4
2 42484 1 4
2 42485 1 4
2 42486 1 4
2 42487 1 4
2 42488 1 4
2 42489 1 4
2 42490 1 4
2 42491 1 4
2 42492 1 4
2 42493 1 4
2 42494 1 4
2 42495 1 4
2 42496 1 4
2 42497 1 4
2 42498 1 4
2 42499 1 4
2 42500 1 4
2 42501 1 4
2 42502 1 4
2 42503 1 4
2 42504 1 4
2 42505 1 4
2 42506 1 4
2 42507 1 4
2 42508 1 4
2 42509 1 4
2 42510 1 4
2 42511 1 4
2 42512 1 4
2 42513 1 4
2 42514 1 4
2 42515 1 4
2 42516 1 4
2 42517 1 4
2 42518 1 4
2 42519 1 4
2 42520 1 4
2 42521 1 4
2 42522 1 4
2 42523 1 4
2 42524 1 4
2 42525 1 4
2 42526 1 4
2 42527 1 4
2 42528 1 4
2 42529 1 4
2 42530 1 4
2 42531 1 4
2 42532 1 4
2 42533 1 4
2 42534 1 4
2 42535 1 4
2 42536 1 4
2 42537 1 4
2 42538 1 4
2 42539 1 4
2 42540 1 4
2 42541 1 4
2 42542 1 4
2 42543 1 4
2 42544 1 4
2 42545 1 4
2 42546 1 4
2 42547 1 4
2 42548 1 4
2 42549 1 4
2 42550 1 4
2 42551 1 4
2 42552 1 4
2 42553 1 4
2 42554 1 4
2 42555 1 4
2 42556 1 4
2 42557 1 4
2 42558 1 4
2 42559 1 4
2 42560 1 4
2 42561 1 4
2 42562 1 4
2 42563 1 4
2 42564 1 4
2 42565 1 4
2 42566 1 4
2 42567 1 4
2 42568 1 4
2 42569 1 4
2 42570 1 4
2 42571 1 4
2 42572 1 4
2 42573 1 4
2 42574 1 4
2 42575 1 4
2 42576 1 4
2 42577 1 4
2 42578 1 4
2 42579 1 4
2 42580 1 4
2 42581 1 4
2 42582 1 4
2 42583 1 4
2 42584 1 4
2 42585 1 4
2 42586 1 4
2 42587 1 4
2 42588 1 4
2 42589 1 4
2 42590 1 4
2 42591 1 4
2 42592 1 4
2 42593 1 4
2 42594 1 4
2 42595 1 4
2 42596 1 4
2 42597 1 4
2 42598 1 4
2 42599 1 4
2 42600 1 4
2 42601 1 4
2 42602 1 4
2 42603 1 4
2 42604 1 4
2 42605 1 4
2 42606 1 4
2 42607 1 4
2 42608 1 4
2 42609 1 4
2 42610 1 4
2 42611 1 4
2 42612 1 4
2 42613 1 4
2 42614 1 4
2 42615 1 4
2 42616 1 4
2 42617 1 4
2 42618 1 4
2 42619 1 4
2 42620 1 4
2 42621 1 4
2 42622 1 4
2 42623 1 4
2 42624 1 4
2 42625 1 4
2 42626 1 4
2 42627 1 4
2 42628 1 4
2 42629 1 4
2 42630 1 4
2 42631 1 4
2 42632 1 4
2 42633 1 4
2 42634 1 4
2 42635 1 4
2 42636 1 4
2 42637 1 4
2 42638 1 4
2 42639 1 4
1 5 0 295 0
2 42640 1 5
2 42641 1 5
2 42642 1 5
2 42643 1 5
2 42644 1 5
2 42645 1 5
2 42646 1 5
2 42647 1 5
2 42648 1 5
2 42649 1 5
2 42650 1 5
2 42651 1 5
2 42652 1 5
2 42653 1 5
2 42654 1 5
2 42655 1 5
2 42656 1 5
2 42657 1 5
2 42658 1 5
2 42659 1 5
2 42660 1 5
2 42661 1 5
2 42662 1 5
2 42663 1 5
2 42664 1 5
2 42665 1 5
2 42666 1 5
2 42667 1 5
2 42668 1 5
2 42669 1 5
2 42670 1 5
2 42671 1 5
2 42672 1 5
2 42673 1 5
2 42674 1 5
2 42675 1 5
2 42676 1 5
2 42677 1 5
2 42678 1 5
2 42679 1 5
2 42680 1 5
2 42681 1 5
2 42682 1 5
2 42683 1 5
2 42684 1 5
2 42685 1 5
2 42686 1 5
2 42687 1 5
2 42688 1 5
2 42689 1 5
2 42690 1 5
2 42691 1 5
2 42692 1 5
2 42693 1 5
2 42694 1 5
2 42695 1 5
2 42696 1 5
2 42697 1 5
2 42698 1 5
2 42699 1 5
2 42700 1 5
2 42701 1 5
2 42702 1 5
2 42703 1 5
2 42704 1 5
2 42705 1 5
2 42706 1 5
2 42707 1 5
2 42708 1 5
2 42709 1 5
2 42710 1 5
2 42711 1 5
2 42712 1 5
2 42713 1 5
2 42714 1 5
2 42715 1 5
2 42716 1 5
2 42717 1 5
2 42718 1 5
2 42719 1 5
2 42720 1 5
2 42721 1 5
2 42722 1 5
2 42723 1 5
2 42724 1 5
2 42725 1 5
2 42726 1 5
2 42727 1 5
2 42728 1 5
2 42729 1 5
2 42730 1 5
2 42731 1 5
2 42732 1 5
2 42733 1 5
2 42734 1 5
2 42735 1 5
2 42736 1 5
2 42737 1 5
2 42738 1 5
2 42739 1 5
2 42740 1 5
2 42741 1 5
2 42742 1 5
2 42743 1 5
2 42744 1 5
2 42745 1 5
2 42746 1 5
2 42747 1 5
2 42748 1 5
2 42749 1 5
2 42750 1 5
2 42751 1 5
2 42752 1 5
2 42753 1 5
2 42754 1 5
2 42755 1 5
2 42756 1 5
2 42757 1 5
2 42758 1 5
2 42759 1 5
2 42760 1 5
2 42761 1 5
2 42762 1 5
2 42763 1 5
2 42764 1 5
2 42765 1 5
2 42766 1 5
2 42767 1 5
2 42768 1 5
2 42769 1 5
2 42770 1 5
2 42771 1 5
2 42772 1 5
2 42773 1 5
2 42774 1 5
2 42775 1 5
2 42776 1 5
2 42777 1 5
2 42778 1 5
2 42779 1 5
2 42780 1 5
2 42781 1 5
2 42782 1 5
2 42783 1 5
2 42784 1 5
2 42785 1 5
2 42786 1 5
2 42787 1 5
2 42788 1 5
2 42789 1 5
2 42790 1 5
2 42791 1 5
2 42792 1 5
2 42793 1 5
2 42794 1 5
2 42795 1 5
2 42796 1 5
2 42797 1 5
2 42798 1 5
2 42799 1 5
2 42800 1 5
2 42801 1 5
2 42802 1 5
2 42803 1 5
2 42804 1 5
2 42805 1 5
2 42806 1 5
2 42807 1 5
2 42808 1 5
2 42809 1 5
2 42810 1 5
2 42811 1 5
2 42812 1 5
2 42813 1 5
2 42814 1 5
2 42815 1 5
2 42816 1 5
2 42817 1 5
2 42818 1 5
2 42819 1 5
2 42820 1 5
2 42821 1 5
2 42822 1 5
2 42823 1 5
2 42824 1 5
2 42825 1 5
2 42826 1 5
2 42827 1 5
2 42828 1 5
2 42829 1 5
2 42830 1 5
2 42831 1 5
2 42832 1 5
2 42833 1 5
2 42834 1 5
2 42835 1 5
2 42836 1 5
2 42837 1 5
2 42838 1 5
2 42839 1 5
2 42840 1 5
2 42841 1 5
2 42842 1 5
2 42843 1 5
2 42844 1 5
2 42845 1 5
2 42846 1 5
2 42847 1 5
2 42848 1 5
2 42849 1 5
2 42850 1 5
2 42851 1 5
2 42852 1 5
2 42853 1 5
2 42854 1 5
2 42855 1 5
2 42856 1 5
2 42857 1 5
2 42858 1 5
2 42859 1 5
2 42860 1 5
2 42861 1 5
2 42862 1 5
2 42863 1 5
2 42864 1 5
2 42865 1 5
2 42866 1 5
2 42867 1 5
2 42868 1 5
2 42869 1 5
2 42870 1 5
2 42871 1 5
2 42872 1 5
2 42873 1 5
2 42874 1 5
2 42875 1 5
2 42876 1 5
2 42877 1 5
2 42878 1 5
2 42879 1 5
2 42880 1 5
2 42881 1 5
2 42882 1 5
2 42883 1 5
2 42884 1 5
2 42885 1 5
2 42886 1 5
2 42887 1 5
2 42888 1 5
2 42889 1 5
2 42890 1 5
2 42891 1 5
2 42892 1 5
2 42893 1 5
2 42894 1 5
2 42895 1 5
2 42896 1 5
2 42897 1 5
2 42898 1 5
2 42899 1 5
2 42900 1 5
2 42901 1 5
2 42902 1 5
2 42903 1 5
2 42904 1 5
2 42905 1 5
2 42906 1 5
2 42907 1 5
2 42908 1 5
2 42909 1 5
2 42910 1 5
2 42911 1 5
2 42912 1 5
2 42913 1 5
2 42914 1 5
2 42915 1 5
2 42916 1 5
2 42917 1 5
2 42918 1 5
2 42919 1 5
2 42920 1 5
2 42921 1 5
2 42922 1 5
2 42923 1 5
2 42924 1 5
2 42925 1 5
2 42926 1 5
2 42927 1 5
2 42928 1 5
2 42929 1 5
2 42930 1 5
2 42931 1 5
2 42932 1 5
2 42933 1 5
2 42934 1 5
1 6 0 249 0
2 42935 1 6
2 42936 1 6
2 42937 1 6
2 42938 1 6
2 42939 1 6
2 42940 1 6
2 42941 1 6
2 42942 1 6
2 42943 1 6
2 42944 1 6
2 42945 1 6
2 42946 1 6
2 42947 1 6
2 42948 1 6
2 42949 1 6
2 42950 1 6
2 42951 1 6
2 42952 1 6
2 42953 1 6
2 42954 1 6
2 42955 1 6
2 42956 1 6
2 42957 1 6
2 42958 1 6
2 42959 1 6
2 42960 1 6
2 42961 1 6
2 42962 1 6
2 42963 1 6
2 42964 1 6
2 42965 1 6
2 42966 1 6
2 42967 1 6
2 42968 1 6
2 42969 1 6
2 42970 1 6
2 42971 1 6
2 42972 1 6
2 42973 1 6
2 42974 1 6
2 42975 1 6
2 42976 1 6
2 42977 1 6
2 42978 1 6
2 42979 1 6
2 42980 1 6
2 42981 1 6
2 42982 1 6
2 42983 1 6
2 42984 1 6
2 42985 1 6
2 42986 1 6
2 42987 1 6
2 42988 1 6
2 42989 1 6
2 42990 1 6
2 42991 1 6
2 42992 1 6
2 42993 1 6
2 42994 1 6
2 42995 1 6
2 42996 1 6
2 42997 1 6
2 42998 1 6
2 42999 1 6
2 43000 1 6
2 43001 1 6
2 43002 1 6
2 43003 1 6
2 43004 1 6
2 43005 1 6
2 43006 1 6
2 43007 1 6
2 43008 1 6
2 43009 1 6
2 43010 1 6
2 43011 1 6
2 43012 1 6
2 43013 1 6
2 43014 1 6
2 43015 1 6
2 43016 1 6
2 43017 1 6
2 43018 1 6
2 43019 1 6
2 43020 1 6
2 43021 1 6
2 43022 1 6
2 43023 1 6
2 43024 1 6
2 43025 1 6
2 43026 1 6
2 43027 1 6
2 43028 1 6
2 43029 1 6
2 43030 1 6
2 43031 1 6
2 43032 1 6
2 43033 1 6
2 43034 1 6
2 43035 1 6
2 43036 1 6
2 43037 1 6
2 43038 1 6
2 43039 1 6
2 43040 1 6
2 43041 1 6
2 43042 1 6
2 43043 1 6
2 43044 1 6
2 43045 1 6
2 43046 1 6
2 43047 1 6
2 43048 1 6
2 43049 1 6
2 43050 1 6
2 43051 1 6
2 43052 1 6
2 43053 1 6
2 43054 1 6
2 43055 1 6
2 43056 1 6
2 43057 1 6
2 43058 1 6
2 43059 1 6
2 43060 1 6
2 43061 1 6
2 43062 1 6
2 43063 1 6
2 43064 1 6
2 43065 1 6
2 43066 1 6
2 43067 1 6
2 43068 1 6
2 43069 1 6
2 43070 1 6
2 43071 1 6
2 43072 1 6
2 43073 1 6
2 43074 1 6
2 43075 1 6
2 43076 1 6
2 43077 1 6
2 43078 1 6
2 43079 1 6
2 43080 1 6
2 43081 1 6
2 43082 1 6
2 43083 1 6
2 43084 1 6
2 43085 1 6
2 43086 1 6
2 43087 1 6
2 43088 1 6
2 43089 1 6
2 43090 1 6
2 43091 1 6
2 43092 1 6
2 43093 1 6
2 43094 1 6
2 43095 1 6
2 43096 1 6
2 43097 1 6
2 43098 1 6
2 43099 1 6
2 43100 1 6
2 43101 1 6
2 43102 1 6
2 43103 1 6
2 43104 1 6
2 43105 1 6
2 43106 1 6
2 43107 1 6
2 43108 1 6
2 43109 1 6
2 43110 1 6
2 43111 1 6
2 43112 1 6
2 43113 1 6
2 43114 1 6
2 43115 1 6
2 43116 1 6
2 43117 1 6
2 43118 1 6
2 43119 1 6
2 43120 1 6
2 43121 1 6
2 43122 1 6
2 43123 1 6
2 43124 1 6
2 43125 1 6
2 43126 1 6
2 43127 1 6
2 43128 1 6
2 43129 1 6
2 43130 1 6
2 43131 1 6
2 43132 1 6
2 43133 1 6
2 43134 1 6
2 43135 1 6
2 43136 1 6
2 43137 1 6
2 43138 1 6
2 43139 1 6
2 43140 1 6
2 43141 1 6
2 43142 1 6
2 43143 1 6
2 43144 1 6
2 43145 1 6
2 43146 1 6
2 43147 1 6
2 43148 1 6
2 43149 1 6
2 43150 1 6
2 43151 1 6
2 43152 1 6
2 43153 1 6
2 43154 1 6
2 43155 1 6
2 43156 1 6
2 43157 1 6
2 43158 1 6
2 43159 1 6
2 43160 1 6
2 43161 1 6
2 43162 1 6
2 43163 1 6
2 43164 1 6
2 43165 1 6
2 43166 1 6
2 43167 1 6
2 43168 1 6
2 43169 1 6
2 43170 1 6
2 43171 1 6
2 43172 1 6
2 43173 1 6
2 43174 1 6
2 43175 1 6
2 43176 1 6
2 43177 1 6
2 43178 1 6
2 43179 1 6
2 43180 1 6
2 43181 1 6
2 43182 1 6
2 43183 1 6
1 7 0 225 0
2 43184 1 7
2 43185 1 7
2 43186 1 7
2 43187 1 7
2 43188 1 7
2 43189 1 7
2 43190 1 7
2 43191 1 7
2 43192 1 7
2 43193 1 7
2 43194 1 7
2 43195 1 7
2 43196 1 7
2 43197 1 7
2 43198 1 7
2 43199 1 7
2 43200 1 7
2 43201 1 7
2 43202 1 7
2 43203 1 7
2 43204 1 7
2 43205 1 7
2 43206 1 7
2 43207 1 7
2 43208 1 7
2 43209 1 7
2 43210 1 7
2 43211 1 7
2 43212 1 7
2 43213 1 7
2 43214 1 7
2 43215 1 7
2 43216 1 7
2 43217 1 7
2 43218 1 7
2 43219 1 7
2 43220 1 7
2 43221 1 7
2 43222 1 7
2 43223 1 7
2 43224 1 7
2 43225 1 7
2 43226 1 7
2 43227 1 7
2 43228 1 7
2 43229 1 7
2 43230 1 7
2 43231 1 7
2 43232 1 7
2 43233 1 7
2 43234 1 7
2 43235 1 7
2 43236 1 7
2 43237 1 7
2 43238 1 7
2 43239 1 7
2 43240 1 7
2 43241 1 7
2 43242 1 7
2 43243 1 7
2 43244 1 7
2 43245 1 7
2 43246 1 7
2 43247 1 7
2 43248 1 7
2 43249 1 7
2 43250 1 7
2 43251 1 7
2 43252 1 7
2 43253 1 7
2 43254 1 7
2 43255 1 7
2 43256 1 7
2 43257 1 7
2 43258 1 7
2 43259 1 7
2 43260 1 7
2 43261 1 7
2 43262 1 7
2 43263 1 7
2 43264 1 7
2 43265 1 7
2 43266 1 7
2 43267 1 7
2 43268 1 7
2 43269 1 7
2 43270 1 7
2 43271 1 7
2 43272 1 7
2 43273 1 7
2 43274 1 7
2 43275 1 7
2 43276 1 7
2 43277 1 7
2 43278 1 7
2 43279 1 7
2 43280 1 7
2 43281 1 7
2 43282 1 7
2 43283 1 7
2 43284 1 7
2 43285 1 7
2 43286 1 7
2 43287 1 7
2 43288 1 7
2 43289 1 7
2 43290 1 7
2 43291 1 7
2 43292 1 7
2 43293 1 7
2 43294 1 7
2 43295 1 7
2 43296 1 7
2 43297 1 7
2 43298 1 7
2 43299 1 7
2 43300 1 7
2 43301 1 7
2 43302 1 7
2 43303 1 7
2 43304 1 7
2 43305 1 7
2 43306 1 7
2 43307 1 7
2 43308 1 7
2 43309 1 7
2 43310 1 7
2 43311 1 7
2 43312 1 7
2 43313 1 7
2 43314 1 7
2 43315 1 7
2 43316 1 7
2 43317 1 7
2 43318 1 7
2 43319 1 7
2 43320 1 7
2 43321 1 7
2 43322 1 7
2 43323 1 7
2 43324 1 7
2 43325 1 7
2 43326 1 7
2 43327 1 7
2 43328 1 7
2 43329 1 7
2 43330 1 7
2 43331 1 7
2 43332 1 7
2 43333 1 7
2 43334 1 7
2 43335 1 7
2 43336 1 7
2 43337 1 7
2 43338 1 7
2 43339 1 7
2 43340 1 7
2 43341 1 7
2 43342 1 7
2 43343 1 7
2 43344 1 7
2 43345 1 7
2 43346 1 7
2 43347 1 7
2 43348 1 7
2 43349 1 7
2 43350 1 7
2 43351 1 7
2 43352 1 7
2 43353 1 7
2 43354 1 7
2 43355 1 7
2 43356 1 7
2 43357 1 7
2 43358 1 7
2 43359 1 7
2 43360 1 7
2 43361 1 7
2 43362 1 7
2 43363 1 7
2 43364 1 7
2 43365 1 7
2 43366 1 7
2 43367 1 7
2 43368 1 7
2 43369 1 7
2 43370 1 7
2 43371 1 7
2 43372 1 7
2 43373 1 7
2 43374 1 7
2 43375 1 7
2 43376 1 7
2 43377 1 7
2 43378 1 7
2 43379 1 7
2 43380 1 7
2 43381 1 7
2 43382 1 7
2 43383 1 7
2 43384 1 7
2 43385 1 7
2 43386 1 7
2 43387 1 7
2 43388 1 7
2 43389 1 7
2 43390 1 7
2 43391 1 7
2 43392 1 7
2 43393 1 7
2 43394 1 7
2 43395 1 7
2 43396 1 7
2 43397 1 7
2 43398 1 7
2 43399 1 7
2 43400 1 7
2 43401 1 7
2 43402 1 7
2 43403 1 7
2 43404 1 7
2 43405 1 7
2 43406 1 7
2 43407 1 7
2 43408 1 7
1 8 0 78 0
2 43409 1 8
2 43410 1 8
2 43411 1 8
2 43412 1 8
2 43413 1 8
2 43414 1 8
2 43415 1 8
2 43416 1 8
2 43417 1 8
2 43418 1 8
2 43419 1 8
2 43420 1 8
2 43421 1 8
2 43422 1 8
2 43423 1 8
2 43424 1 8
2 43425 1 8
2 43426 1 8
2 43427 1 8
2 43428 1 8
2 43429 1 8
2 43430 1 8
2 43431 1 8
2 43432 1 8
2 43433 1 8
2 43434 1 8
2 43435 1 8
2 43436 1 8
2 43437 1 8
2 43438 1 8
2 43439 1 8
2 43440 1 8
2 43441 1 8
2 43442 1 8
2 43443 1 8
2 43444 1 8
2 43445 1 8
2 43446 1 8
2 43447 1 8
2 43448 1 8
2 43449 1 8
2 43450 1 8
2 43451 1 8
2 43452 1 8
2 43453 1 8
2 43454 1 8
2 43455 1 8
2 43456 1 8
2 43457 1 8
2 43458 1 8
2 43459 1 8
2 43460 1 8
2 43461 1 8
2 43462 1 8
2 43463 1 8
2 43464 1 8
2 43465 1 8
2 43466 1 8
2 43467 1 8
2 43468 1 8
2 43469 1 8
2 43470 1 8
2 43471 1 8
2 43472 1 8
2 43473 1 8
2 43474 1 8
2 43475 1 8
2 43476 1 8
2 43477 1 8
2 43478 1 8
2 43479 1 8
2 43480 1 8
2 43481 1 8
2 43482 1 8
2 43483 1 8
2 43484 1 8
2 43485 1 8
2 43486 1 8
1 9 0 80 0
2 43487 1 9
2 43488 1 9
2 43489 1 9
2 43490 1 9
2 43491 1 9
2 43492 1 9
2 43493 1 9
2 43494 1 9
2 43495 1 9
2 43496 1 9
2 43497 1 9
2 43498 1 9
2 43499 1 9
2 43500 1 9
2 43501 1 9
2 43502 1 9
2 43503 1 9
2 43504 1 9
2 43505 1 9
2 43506 1 9
2 43507 1 9
2 43508 1 9
2 43509 1 9
2 43510 1 9
2 43511 1 9
2 43512 1 9
2 43513 1 9
2 43514 1 9
2 43515 1 9
2 43516 1 9
2 43517 1 9
2 43518 1 9
2 43519 1 9
2 43520 1 9
2 43521 1 9
2 43522 1 9
2 43523 1 9
2 43524 1 9
2 43525 1 9
2 43526 1 9
2 43527 1 9
2 43528 1 9
2 43529 1 9
2 43530 1 9
2 43531 1 9
2 43532 1 9
2 43533 1 9
2 43534 1 9
2 43535 1 9
2 43536 1 9
2 43537 1 9
2 43538 1 9
2 43539 1 9
2 43540 1 9
2 43541 1 9
2 43542 1 9
2 43543 1 9
2 43544 1 9
2 43545 1 9
2 43546 1 9
2 43547 1 9
2 43548 1 9
2 43549 1 9
2 43550 1 9
2 43551 1 9
2 43552 1 9
2 43553 1 9
2 43554 1 9
2 43555 1 9
2 43556 1 9
2 43557 1 9
2 43558 1 9
2 43559 1 9
2 43560 1 9
2 43561 1 9
2 43562 1 9
2 43563 1 9
2 43564 1 9
2 43565 1 9
2 43566 1 9
1 10 0 40 0
2 43567 1 10
2 43568 1 10
2 43569 1 10
2 43570 1 10
2 43571 1 10
2 43572 1 10
2 43573 1 10
2 43574 1 10
2 43575 1 10
2 43576 1 10
2 43577 1 10
2 43578 1 10
2 43579 1 10
2 43580 1 10
2 43581 1 10
2 43582 1 10
2 43583 1 10
2 43584 1 10
2 43585 1 10
2 43586 1 10
2 43587 1 10
2 43588 1 10
2 43589 1 10
2 43590 1 10
2 43591 1 10
2 43592 1 10
2 43593 1 10
2 43594 1 10
2 43595 1 10
2 43596 1 10
2 43597 1 10
2 43598 1 10
2 43599 1 10
2 43600 1 10
2 43601 1 10
2 43602 1 10
2 43603 1 10
2 43604 1 10
2 43605 1 10
2 43606 1 10
1 11 0 41 0
2 43607 1 11
2 43608 1 11
2 43609 1 11
2 43610 1 11
2 43611 1 11
2 43612 1 11
2 43613 1 11
2 43614 1 11
2 43615 1 11
2 43616 1 11
2 43617 1 11
2 43618 1 11
2 43619 1 11
2 43620 1 11
2 43621 1 11
2 43622 1 11
2 43623 1 11
2 43624 1 11
2 43625 1 11
2 43626 1 11
2 43627 1 11
2 43628 1 11
2 43629 1 11
2 43630 1 11
2 43631 1 11
2 43632 1 11
2 43633 1 11
2 43634 1 11
2 43635 1 11
2 43636 1 11
2 43637 1 11
2 43638 1 11
2 43639 1 11
2 43640 1 11
2 43641 1 11
2 43642 1 11
2 43643 1 11
2 43644 1 11
2 43645 1 11
2 43646 1 11
2 43647 1 11
1 12 0 135 0
2 43648 1 12
2 43649 1 12
2 43650 1 12
2 43651 1 12
2 43652 1 12
2 43653 1 12
2 43654 1 12
2 43655 1 12
2 43656 1 12
2 43657 1 12
2 43658 1 12
2 43659 1 12
2 43660 1 12
2 43661 1 12
2 43662 1 12
2 43663 1 12
2 43664 1 12
2 43665 1 12
2 43666 1 12
2 43667 1 12
2 43668 1 12
2 43669 1 12
2 43670 1 12
2 43671 1 12
2 43672 1 12
2 43673 1 12
2 43674 1 12
2 43675 1 12
2 43676 1 12
2 43677 1 12
2 43678 1 12
2 43679 1 12
2 43680 1 12
2 43681 1 12
2 43682 1 12
2 43683 1 12
2 43684 1 12
2 43685 1 12
2 43686 1 12
2 43687 1 12
2 43688 1 12
2 43689 1 12
2 43690 1 12
2 43691 1 12
2 43692 1 12
2 43693 1 12
2 43694 1 12
2 43695 1 12
2 43696 1 12
2 43697 1 12
2 43698 1 12
2 43699 1 12
2 43700 1 12
2 43701 1 12
2 43702 1 12
2 43703 1 12
2 43704 1 12
2 43705 1 12
2 43706 1 12
2 43707 1 12
2 43708 1 12
2 43709 1 12
2 43710 1 12
2 43711 1 12
2 43712 1 12
2 43713 1 12
2 43714 1 12
2 43715 1 12
2 43716 1 12
2 43717 1 12
2 43718 1 12
2 43719 1 12
2 43720 1 12
2 43721 1 12
2 43722 1 12
2 43723 1 12
2 43724 1 12
2 43725 1 12
2 43726 1 12
2 43727 1 12
2 43728 1 12
2 43729 1 12
2 43730 1 12
2 43731 1 12
2 43732 1 12
2 43733 1 12
2 43734 1 12
2 43735 1 12
2 43736 1 12
2 43737 1 12
2 43738 1 12
2 43739 1 12
2 43740 1 12
2 43741 1 12
2 43742 1 12
2 43743 1 12
2 43744 1 12
2 43745 1 12
2 43746 1 12
2 43747 1 12
2 43748 1 12
2 43749 1 12
2 43750 1 12
2 43751 1 12
2 43752 1 12
2 43753 1 12
2 43754 1 12
2 43755 1 12
2 43756 1 12
2 43757 1 12
2 43758 1 12
2 43759 1 12
2 43760 1 12
2 43761 1 12
2 43762 1 12
2 43763 1 12
2 43764 1 12
2 43765 1 12
2 43766 1 12
2 43767 1 12
2 43768 1 12
2 43769 1 12
2 43770 1 12
2 43771 1 12
2 43772 1 12
2 43773 1 12
2 43774 1 12
2 43775 1 12
2 43776 1 12
2 43777 1 12
2 43778 1 12
2 43779 1 12
2 43780 1 12
2 43781 1 12
2 43782 1 12
1 13 0 169 0
2 43783 1 13
2 43784 1 13
2 43785 1 13
2 43786 1 13
2 43787 1 13
2 43788 1 13
2 43789 1 13
2 43790 1 13
2 43791 1 13
2 43792 1 13
2 43793 1 13
2 43794 1 13
2 43795 1 13
2 43796 1 13
2 43797 1 13
2 43798 1 13
2 43799 1 13
2 43800 1 13
2 43801 1 13
2 43802 1 13
2 43803 1 13
2 43804 1 13
2 43805 1 13
2 43806 1 13
2 43807 1 13
2 43808 1 13
2 43809 1 13
2 43810 1 13
2 43811 1 13
2 43812 1 13
2 43813 1 13
2 43814 1 13
2 43815 1 13
2 43816 1 13
2 43817 1 13
2 43818 1 13
2 43819 1 13
2 43820 1 13
2 43821 1 13
2 43822 1 13
2 43823 1 13
2 43824 1 13
2 43825 1 13
2 43826 1 13
2 43827 1 13
2 43828 1 13
2 43829 1 13
2 43830 1 13
2 43831 1 13
2 43832 1 13
2 43833 1 13
2 43834 1 13
2 43835 1 13
2 43836 1 13
2 43837 1 13
2 43838 1 13
2 43839 1 13
2 43840 1 13
2 43841 1 13
2 43842 1 13
2 43843 1 13
2 43844 1 13
2 43845 1 13
2 43846 1 13
2 43847 1 13
2 43848 1 13
2 43849 1 13
2 43850 1 13
2 43851 1 13
2 43852 1 13
2 43853 1 13
2 43854 1 13
2 43855 1 13
2 43856 1 13
2 43857 1 13
2 43858 1 13
2 43859 1 13
2 43860 1 13
2 43861 1 13
2 43862 1 13
2 43863 1 13
2 43864 1 13
2 43865 1 13
2 43866 1 13
2 43867 1 13
2 43868 1 13
2 43869 1 13
2 43870 1 13
2 43871 1 13
2 43872 1 13
2 43873 1 13
2 43874 1 13
2 43875 1 13
2 43876 1 13
2 43877 1 13
2 43878 1 13
2 43879 1 13
2 43880 1 13
2 43881 1 13
2 43882 1 13
2 43883 1 13
2 43884 1 13
2 43885 1 13
2 43886 1 13
2 43887 1 13
2 43888 1 13
2 43889 1 13
2 43890 1 13
2 43891 1 13
2 43892 1 13
2 43893 1 13
2 43894 1 13
2 43895 1 13
2 43896 1 13
2 43897 1 13
2 43898 1 13
2 43899 1 13
2 43900 1 13
2 43901 1 13
2 43902 1 13
2 43903 1 13
2 43904 1 13
2 43905 1 13
2 43906 1 13
2 43907 1 13
2 43908 1 13
2 43909 1 13
2 43910 1 13
2 43911 1 13
2 43912 1 13
2 43913 1 13
2 43914 1 13
2 43915 1 13
2 43916 1 13
2 43917 1 13
2 43918 1 13
2 43919 1 13
2 43920 1 13
2 43921 1 13
2 43922 1 13
2 43923 1 13
2 43924 1 13
2 43925 1 13
2 43926 1 13
2 43927 1 13
2 43928 1 13
2 43929 1 13
2 43930 1 13
2 43931 1 13
2 43932 1 13
2 43933 1 13
2 43934 1 13
2 43935 1 13
2 43936 1 13
2 43937 1 13
2 43938 1 13
2 43939 1 13
2 43940 1 13
2 43941 1 13
2 43942 1 13
2 43943 1 13
2 43944 1 13
2 43945 1 13
2 43946 1 13
2 43947 1 13
2 43948 1 13
2 43949 1 13
2 43950 1 13
2 43951 1 13
1 14 0 177 0
2 43952 1 14
2 43953 1 14
2 43954 1 14
2 43955 1 14
2 43956 1 14
2 43957 1 14
2 43958 1 14
2 43959 1 14
2 43960 1 14
2 43961 1 14
2 43962 1 14
2 43963 1 14
2 43964 1 14
2 43965 1 14
2 43966 1 14
2 43967 1 14
2 43968 1 14
2 43969 1 14
2 43970 1 14
2 43971 1 14
2 43972 1 14
2 43973 1 14
2 43974 1 14
2 43975 1 14
2 43976 1 14
2 43977 1 14
2 43978 1 14
2 43979 1 14
2 43980 1 14
2 43981 1 14
2 43982 1 14
2 43983 1 14
2 43984 1 14
2 43985 1 14
2 43986 1 14
2 43987 1 14
2 43988 1 14
2 43989 1 14
2 43990 1 14
2 43991 1 14
2 43992 1 14
2 43993 1 14
2 43994 1 14
2 43995 1 14
2 43996 1 14
2 43997 1 14
2 43998 1 14
2 43999 1 14
2 44000 1 14
2 44001 1 14
2 44002 1 14
2 44003 1 14
2 44004 1 14
2 44005 1 14
2 44006 1 14
2 44007 1 14
2 44008 1 14
2 44009 1 14
2 44010 1 14
2 44011 1 14
2 44012 1 14
2 44013 1 14
2 44014 1 14
2 44015 1 14
2 44016 1 14
2 44017 1 14
2 44018 1 14
2 44019 1 14
2 44020 1 14
2 44021 1 14
2 44022 1 14
2 44023 1 14
2 44024 1 14
2 44025 1 14
2 44026 1 14
2 44027 1 14
2 44028 1 14
2 44029 1 14
2 44030 1 14
2 44031 1 14
2 44032 1 14
2 44033 1 14
2 44034 1 14
2 44035 1 14
2 44036 1 14
2 44037 1 14
2 44038 1 14
2 44039 1 14
2 44040 1 14
2 44041 1 14
2 44042 1 14
2 44043 1 14
2 44044 1 14
2 44045 1 14
2 44046 1 14
2 44047 1 14
2 44048 1 14
2 44049 1 14
2 44050 1 14
2 44051 1 14
2 44052 1 14
2 44053 1 14
2 44054 1 14
2 44055 1 14
2 44056 1 14
2 44057 1 14
2 44058 1 14
2 44059 1 14
2 44060 1 14
2 44061 1 14
2 44062 1 14
2 44063 1 14
2 44064 1 14
2 44065 1 14
2 44066 1 14
2 44067 1 14
2 44068 1 14
2 44069 1 14
2 44070 1 14
2 44071 1 14
2 44072 1 14
2 44073 1 14
2 44074 1 14
2 44075 1 14
2 44076 1 14
2 44077 1 14
2 44078 1 14
2 44079 1 14
2 44080 1 14
2 44081 1 14
2 44082 1 14
2 44083 1 14
2 44084 1 14
2 44085 1 14
2 44086 1 14
2 44087 1 14
2 44088 1 14
2 44089 1 14
2 44090 1 14
2 44091 1 14
2 44092 1 14
2 44093 1 14
2 44094 1 14
2 44095 1 14
2 44096 1 14
2 44097 1 14
2 44098 1 14
2 44099 1 14
2 44100 1 14
2 44101 1 14
2 44102 1 14
2 44103 1 14
2 44104 1 14
2 44105 1 14
2 44106 1 14
2 44107 1 14
2 44108 1 14
2 44109 1 14
2 44110 1 14
2 44111 1 14
2 44112 1 14
2 44113 1 14
2 44114 1 14
2 44115 1 14
2 44116 1 14
2 44117 1 14
2 44118 1 14
2 44119 1 14
2 44120 1 14
2 44121 1 14
2 44122 1 14
2 44123 1 14
2 44124 1 14
2 44125 1 14
2 44126 1 14
2 44127 1 14
2 44128 1 14
1 15 0 148 0
2 44129 1 15
2 44130 1 15
2 44131 1 15
2 44132 1 15
2 44133 1 15
2 44134 1 15
2 44135 1 15
2 44136 1 15
2 44137 1 15
2 44138 1 15
2 44139 1 15
2 44140 1 15
2 44141 1 15
2 44142 1 15
2 44143 1 15
2 44144 1 15
2 44145 1 15
2 44146 1 15
2 44147 1 15
2 44148 1 15
2 44149 1 15
2 44150 1 15
2 44151 1 15
2 44152 1 15
2 44153 1 15
2 44154 1 15
2 44155 1 15
2 44156 1 15
2 44157 1 15
2 44158 1 15
2 44159 1 15
2 44160 1 15
2 44161 1 15
2 44162 1 15
2 44163 1 15
2 44164 1 15
2 44165 1 15
2 44166 1 15
2 44167 1 15
2 44168 1 15
2 44169 1 15
2 44170 1 15
2 44171 1 15
2 44172 1 15
2 44173 1 15
2 44174 1 15
2 44175 1 15
2 44176 1 15
2 44177 1 15
2 44178 1 15
2 44179 1 15
2 44180 1 15
2 44181 1 15
2 44182 1 15
2 44183 1 15
2 44184 1 15
2 44185 1 15
2 44186 1 15
2 44187 1 15
2 44188 1 15
2 44189 1 15
2 44190 1 15
2 44191 1 15
2 44192 1 15
2 44193 1 15
2 44194 1 15
2 44195 1 15
2 44196 1 15
2 44197 1 15
2 44198 1 15
2 44199 1 15
2 44200 1 15
2 44201 1 15
2 44202 1 15
2 44203 1 15
2 44204 1 15
2 44205 1 15
2 44206 1 15
2 44207 1 15
2 44208 1 15
2 44209 1 15
2 44210 1 15
2 44211 1 15
2 44212 1 15
2 44213 1 15
2 44214 1 15
2 44215 1 15
2 44216 1 15
2 44217 1 15
2 44218 1 15
2 44219 1 15
2 44220 1 15
2 44221 1 15
2 44222 1 15
2 44223 1 15
2 44224 1 15
2 44225 1 15
2 44226 1 15
2 44227 1 15
2 44228 1 15
2 44229 1 15
2 44230 1 15
2 44231 1 15
2 44232 1 15
2 44233 1 15
2 44234 1 15
2 44235 1 15
2 44236 1 15
2 44237 1 15
2 44238 1 15
2 44239 1 15
2 44240 1 15
2 44241 1 15
2 44242 1 15
2 44243 1 15
2 44244 1 15
2 44245 1 15
2 44246 1 15
2 44247 1 15
2 44248 1 15
2 44249 1 15
2 44250 1 15
2 44251 1 15
2 44252 1 15
2 44253 1 15
2 44254 1 15
2 44255 1 15
2 44256 1 15
2 44257 1 15
2 44258 1 15
2 44259 1 15
2 44260 1 15
2 44261 1 15
2 44262 1 15
2 44263 1 15
2 44264 1 15
2 44265 1 15
2 44266 1 15
2 44267 1 15
2 44268 1 15
2 44269 1 15
2 44270 1 15
2 44271 1 15
2 44272 1 15
2 44273 1 15
2 44274 1 15
2 44275 1 15
2 44276 1 15
1 16 0 95 0
2 44277 1 16
2 44278 1 16
2 44279 1 16
2 44280 1 16
2 44281 1 16
2 44282 1 16
2 44283 1 16
2 44284 1 16
2 44285 1 16
2 44286 1 16
2 44287 1 16
2 44288 1 16
2 44289 1 16
2 44290 1 16
2 44291 1 16
2 44292 1 16
2 44293 1 16
2 44294 1 16
2 44295 1 16
2 44296 1 16
2 44297 1 16
2 44298 1 16
2 44299 1 16
2 44300 1 16
2 44301 1 16
2 44302 1 16
2 44303 1 16
2 44304 1 16
2 44305 1 16
2 44306 1 16
2 44307 1 16
2 44308 1 16
2 44309 1 16
2 44310 1 16
2 44311 1 16
2 44312 1 16
2 44313 1 16
2 44314 1 16
2 44315 1 16
2 44316 1 16
2 44317 1 16
2 44318 1 16
2 44319 1 16
2 44320 1 16
2 44321 1 16
2 44322 1 16
2 44323 1 16
2 44324 1 16
2 44325 1 16
2 44326 1 16
2 44327 1 16
2 44328 1 16
2 44329 1 16
2 44330 1 16
2 44331 1 16
2 44332 1 16
2 44333 1 16
2 44334 1 16
2 44335 1 16
2 44336 1 16
2 44337 1 16
2 44338 1 16
2 44339 1 16
2 44340 1 16
2 44341 1 16
2 44342 1 16
2 44343 1 16
2 44344 1 16
2 44345 1 16
2 44346 1 16
2 44347 1 16
2 44348 1 16
2 44349 1 16
2 44350 1 16
2 44351 1 16
2 44352 1 16
2 44353 1 16
2 44354 1 16
2 44355 1 16
2 44356 1 16
2 44357 1 16
2 44358 1 16
2 44359 1 16
2 44360 1 16
2 44361 1 16
2 44362 1 16
2 44363 1 16
2 44364 1 16
2 44365 1 16
2 44366 1 16
2 44367 1 16
2 44368 1 16
2 44369 1 16
2 44370 1 16
2 44371 1 16
1 17 0 136 0
2 44372 1 17
2 44373 1 17
2 44374 1 17
2 44375 1 17
2 44376 1 17
2 44377 1 17
2 44378 1 17
2 44379 1 17
2 44380 1 17
2 44381 1 17
2 44382 1 17
2 44383 1 17
2 44384 1 17
2 44385 1 17
2 44386 1 17
2 44387 1 17
2 44388 1 17
2 44389 1 17
2 44390 1 17
2 44391 1 17
2 44392 1 17
2 44393 1 17
2 44394 1 17
2 44395 1 17
2 44396 1 17
2 44397 1 17
2 44398 1 17
2 44399 1 17
2 44400 1 17
2 44401 1 17
2 44402 1 17
2 44403 1 17
2 44404 1 17
2 44405 1 17
2 44406 1 17
2 44407 1 17
2 44408 1 17
2 44409 1 17
2 44410 1 17
2 44411 1 17
2 44412 1 17
2 44413 1 17
2 44414 1 17
2 44415 1 17
2 44416 1 17
2 44417 1 17
2 44418 1 17
2 44419 1 17
2 44420 1 17
2 44421 1 17
2 44422 1 17
2 44423 1 17
2 44424 1 17
2 44425 1 17
2 44426 1 17
2 44427 1 17
2 44428 1 17
2 44429 1 17
2 44430 1 17
2 44431 1 17
2 44432 1 17
2 44433 1 17
2 44434 1 17
2 44435 1 17
2 44436 1 17
2 44437 1 17
2 44438 1 17
2 44439 1 17
2 44440 1 17
2 44441 1 17
2 44442 1 17
2 44443 1 17
2 44444 1 17
2 44445 1 17
2 44446 1 17
2 44447 1 17
2 44448 1 17
2 44449 1 17
2 44450 1 17
2 44451 1 17
2 44452 1 17
2 44453 1 17
2 44454 1 17
2 44455 1 17
2 44456 1 17
2 44457 1 17
2 44458 1 17
2 44459 1 17
2 44460 1 17
2 44461 1 17
2 44462 1 17
2 44463 1 17
2 44464 1 17
2 44465 1 17
2 44466 1 17
2 44467 1 17
2 44468 1 17
2 44469 1 17
2 44470 1 17
2 44471 1 17
2 44472 1 17
2 44473 1 17
2 44474 1 17
2 44475 1 17
2 44476 1 17
2 44477 1 17
2 44478 1 17
2 44479 1 17
2 44480 1 17
2 44481 1 17
2 44482 1 17
2 44483 1 17
2 44484 1 17
2 44485 1 17
2 44486 1 17
2 44487 1 17
2 44488 1 17
2 44489 1 17
2 44490 1 17
2 44491 1 17
2 44492 1 17
2 44493 1 17
2 44494 1 17
2 44495 1 17
2 44496 1 17
2 44497 1 17
2 44498 1 17
2 44499 1 17
2 44500 1 17
2 44501 1 17
2 44502 1 17
2 44503 1 17
2 44504 1 17
2 44505 1 17
2 44506 1 17
2 44507 1 17
1 18 0 96 0
2 44508 1 18
2 44509 1 18
2 44510 1 18
2 44511 1 18
2 44512 1 18
2 44513 1 18
2 44514 1 18
2 44515 1 18
2 44516 1 18
2 44517 1 18
2 44518 1 18
2 44519 1 18
2 44520 1 18
2 44521 1 18
2 44522 1 18
2 44523 1 18
2 44524 1 18
2 44525 1 18
2 44526 1 18
2 44527 1 18
2 44528 1 18
2 44529 1 18
2 44530 1 18
2 44531 1 18
2 44532 1 18
2 44533 1 18
2 44534 1 18
2 44535 1 18
2 44536 1 18
2 44537 1 18
2 44538 1 18
2 44539 1 18
2 44540 1 18
2 44541 1 18
2 44542 1 18
2 44543 1 18
2 44544 1 18
2 44545 1 18
2 44546 1 18
2 44547 1 18
2 44548 1 18
2 44549 1 18
2 44550 1 18
2 44551 1 18
2 44552 1 18
2 44553 1 18
2 44554 1 18
2 44555 1 18
2 44556 1 18
2 44557 1 18
2 44558 1 18
2 44559 1 18
2 44560 1 18
2 44561 1 18
2 44562 1 18
2 44563 1 18
2 44564 1 18
2 44565 1 18
2 44566 1 18
2 44567 1 18
2 44568 1 18
2 44569 1 18
2 44570 1 18
2 44571 1 18
2 44572 1 18
2 44573 1 18
2 44574 1 18
2 44575 1 18
2 44576 1 18
2 44577 1 18
2 44578 1 18
2 44579 1 18
2 44580 1 18
2 44581 1 18
2 44582 1 18
2 44583 1 18
2 44584 1 18
2 44585 1 18
2 44586 1 18
2 44587 1 18
2 44588 1 18
2 44589 1 18
2 44590 1 18
2 44591 1 18
2 44592 1 18
2 44593 1 18
2 44594 1 18
2 44595 1 18
2 44596 1 18
2 44597 1 18
2 44598 1 18
2 44599 1 18
2 44600 1 18
2 44601 1 18
2 44602 1 18
2 44603 1 18
1 19 0 96 0
2 44604 1 19
2 44605 1 19
2 44606 1 19
2 44607 1 19
2 44608 1 19
2 44609 1 19
2 44610 1 19
2 44611 1 19
2 44612 1 19
2 44613 1 19
2 44614 1 19
2 44615 1 19
2 44616 1 19
2 44617 1 19
2 44618 1 19
2 44619 1 19
2 44620 1 19
2 44621 1 19
2 44622 1 19
2 44623 1 19
2 44624 1 19
2 44625 1 19
2 44626 1 19
2 44627 1 19
2 44628 1 19
2 44629 1 19
2 44630 1 19
2 44631 1 19
2 44632 1 19
2 44633 1 19
2 44634 1 19
2 44635 1 19
2 44636 1 19
2 44637 1 19
2 44638 1 19
2 44639 1 19
2 44640 1 19
2 44641 1 19
2 44642 1 19
2 44643 1 19
2 44644 1 19
2 44645 1 19
2 44646 1 19
2 44647 1 19
2 44648 1 19
2 44649 1 19
2 44650 1 19
2 44651 1 19
2 44652 1 19
2 44653 1 19
2 44654 1 19
2 44655 1 19
2 44656 1 19
2 44657 1 19
2 44658 1 19
2 44659 1 19
2 44660 1 19
2 44661 1 19
2 44662 1 19
2 44663 1 19
2 44664 1 19
2 44665 1 19
2 44666 1 19
2 44667 1 19
2 44668 1 19
2 44669 1 19
2 44670 1 19
2 44671 1 19
2 44672 1 19
2 44673 1 19
2 44674 1 19
2 44675 1 19
2 44676 1 19
2 44677 1 19
2 44678 1 19
2 44679 1 19
2 44680 1 19
2 44681 1 19
2 44682 1 19
2 44683 1 19
2 44684 1 19
2 44685 1 19
2 44686 1 19
2 44687 1 19
2 44688 1 19
2 44689 1 19
2 44690 1 19
2 44691 1 19
2 44692 1 19
2 44693 1 19
2 44694 1 19
2 44695 1 19
2 44696 1 19
2 44697 1 19
2 44698 1 19
2 44699 1 19
1 20 0 139 0
2 44700 1 20
2 44701 1 20
2 44702 1 20
2 44703 1 20
2 44704 1 20
2 44705 1 20
2 44706 1 20
2 44707 1 20
2 44708 1 20
2 44709 1 20
2 44710 1 20
2 44711 1 20
2 44712 1 20
2 44713 1 20
2 44714 1 20
2 44715 1 20
2 44716 1 20
2 44717 1 20
2 44718 1 20
2 44719 1 20
2 44720 1 20
2 44721 1 20
2 44722 1 20
2 44723 1 20
2 44724 1 20
2 44725 1 20
2 44726 1 20
2 44727 1 20
2 44728 1 20
2 44729 1 20
2 44730 1 20
2 44731 1 20
2 44732 1 20
2 44733 1 20
2 44734 1 20
2 44735 1 20
2 44736 1 20
2 44737 1 20
2 44738 1 20
2 44739 1 20
2 44740 1 20
2 44741 1 20
2 44742 1 20
2 44743 1 20
2 44744 1 20
2 44745 1 20
2 44746 1 20
2 44747 1 20
2 44748 1 20
2 44749 1 20
2 44750 1 20
2 44751 1 20
2 44752 1 20
2 44753 1 20
2 44754 1 20
2 44755 1 20
2 44756 1 20
2 44757 1 20
2 44758 1 20
2 44759 1 20
2 44760 1 20
2 44761 1 20
2 44762 1 20
2 44763 1 20
2 44764 1 20
2 44765 1 20
2 44766 1 20
2 44767 1 20
2 44768 1 20
2 44769 1 20
2 44770 1 20
2 44771 1 20
2 44772 1 20
2 44773 1 20
2 44774 1 20
2 44775 1 20
2 44776 1 20
2 44777 1 20
2 44778 1 20
2 44779 1 20
2 44780 1 20
2 44781 1 20
2 44782 1 20
2 44783 1 20
2 44784 1 20
2 44785 1 20
2 44786 1 20
2 44787 1 20
2 44788 1 20
2 44789 1 20
2 44790 1 20
2 44791 1 20
2 44792 1 20
2 44793 1 20
2 44794 1 20
2 44795 1 20
2 44796 1 20
2 44797 1 20
2 44798 1 20
2 44799 1 20
2 44800 1 20
2 44801 1 20
2 44802 1 20
2 44803 1 20
2 44804 1 20
2 44805 1 20
2 44806 1 20
2 44807 1 20
2 44808 1 20
2 44809 1 20
2 44810 1 20
2 44811 1 20
2 44812 1 20
2 44813 1 20
2 44814 1 20
2 44815 1 20
2 44816 1 20
2 44817 1 20
2 44818 1 20
2 44819 1 20
2 44820 1 20
2 44821 1 20
2 44822 1 20
2 44823 1 20
2 44824 1 20
2 44825 1 20
2 44826 1 20
2 44827 1 20
2 44828 1 20
2 44829 1 20
2 44830 1 20
2 44831 1 20
2 44832 1 20
2 44833 1 20
2 44834 1 20
2 44835 1 20
2 44836 1 20
2 44837 1 20
2 44838 1 20
1 21 0 154 0
2 44839 1 21
2 44840 1 21
2 44841 1 21
2 44842 1 21
2 44843 1 21
2 44844 1 21
2 44845 1 21
2 44846 1 21
2 44847 1 21
2 44848 1 21
2 44849 1 21
2 44850 1 21
2 44851 1 21
2 44852 1 21
2 44853 1 21
2 44854 1 21
2 44855 1 21
2 44856 1 21
2 44857 1 21
2 44858 1 21
2 44859 1 21
2 44860 1 21
2 44861 1 21
2 44862 1 21
2 44863 1 21
2 44864 1 21
2 44865 1 21
2 44866 1 21
2 44867 1 21
2 44868 1 21
2 44869 1 21
2 44870 1 21
2 44871 1 21
2 44872 1 21
2 44873 1 21
2 44874 1 21
2 44875 1 21
2 44876 1 21
2 44877 1 21
2 44878 1 21
2 44879 1 21
2 44880 1 21
2 44881 1 21
2 44882 1 21
2 44883 1 21
2 44884 1 21
2 44885 1 21
2 44886 1 21
2 44887 1 21
2 44888 1 21
2 44889 1 21
2 44890 1 21
2 44891 1 21
2 44892 1 21
2 44893 1 21
2 44894 1 21
2 44895 1 21
2 44896 1 21
2 44897 1 21
2 44898 1 21
2 44899 1 21
2 44900 1 21
2 44901 1 21
2 44902 1 21
2 44903 1 21
2 44904 1 21
2 44905 1 21
2 44906 1 21
2 44907 1 21
2 44908 1 21
2 44909 1 21
2 44910 1 21
2 44911 1 21
2 44912 1 21
2 44913 1 21
2 44914 1 21
2 44915 1 21
2 44916 1 21
2 44917 1 21
2 44918 1 21
2 44919 1 21
2 44920 1 21
2 44921 1 21
2 44922 1 21
2 44923 1 21
2 44924 1 21
2 44925 1 21
2 44926 1 21
2 44927 1 21
2 44928 1 21
2 44929 1 21
2 44930 1 21
2 44931 1 21
2 44932 1 21
2 44933 1 21
2 44934 1 21
2 44935 1 21
2 44936 1 21
2 44937 1 21
2 44938 1 21
2 44939 1 21
2 44940 1 21
2 44941 1 21
2 44942 1 21
2 44943 1 21
2 44944 1 21
2 44945 1 21
2 44946 1 21
2 44947 1 21
2 44948 1 21
2 44949 1 21
2 44950 1 21
2 44951 1 21
2 44952 1 21
2 44953 1 21
2 44954 1 21
2 44955 1 21
2 44956 1 21
2 44957 1 21
2 44958 1 21
2 44959 1 21
2 44960 1 21
2 44961 1 21
2 44962 1 21
2 44963 1 21
2 44964 1 21
2 44965 1 21
2 44966 1 21
2 44967 1 21
2 44968 1 21
2 44969 1 21
2 44970 1 21
2 44971 1 21
2 44972 1 21
2 44973 1 21
2 44974 1 21
2 44975 1 21
2 44976 1 21
2 44977 1 21
2 44978 1 21
2 44979 1 21
2 44980 1 21
2 44981 1 21
2 44982 1 21
2 44983 1 21
2 44984 1 21
2 44985 1 21
2 44986 1 21
2 44987 1 21
2 44988 1 21
2 44989 1 21
2 44990 1 21
2 44991 1 21
2 44992 1 21
1 22 0 138 0
2 44993 1 22
2 44994 1 22
2 44995 1 22
2 44996 1 22
2 44997 1 22
2 44998 1 22
2 44999 1 22
2 45000 1 22
2 45001 1 22
2 45002 1 22
2 45003 1 22
2 45004 1 22
2 45005 1 22
2 45006 1 22
2 45007 1 22
2 45008 1 22
2 45009 1 22
2 45010 1 22
2 45011 1 22
2 45012 1 22
2 45013 1 22
2 45014 1 22
2 45015 1 22
2 45016 1 22
2 45017 1 22
2 45018 1 22
2 45019 1 22
2 45020 1 22
2 45021 1 22
2 45022 1 22
2 45023 1 22
2 45024 1 22
2 45025 1 22
2 45026 1 22
2 45027 1 22
2 45028 1 22
2 45029 1 22
2 45030 1 22
2 45031 1 22
2 45032 1 22
2 45033 1 22
2 45034 1 22
2 45035 1 22
2 45036 1 22
2 45037 1 22
2 45038 1 22
2 45039 1 22
2 45040 1 22
2 45041 1 22
2 45042 1 22
2 45043 1 22
2 45044 1 22
2 45045 1 22
2 45046 1 22
2 45047 1 22
2 45048 1 22
2 45049 1 22
2 45050 1 22
2 45051 1 22
2 45052 1 22
2 45053 1 22
2 45054 1 22
2 45055 1 22
2 45056 1 22
2 45057 1 22
2 45058 1 22
2 45059 1 22
2 45060 1 22
2 45061 1 22
2 45062 1 22
2 45063 1 22
2 45064 1 22
2 45065 1 22
2 45066 1 22
2 45067 1 22
2 45068 1 22
2 45069 1 22
2 45070 1 22
2 45071 1 22
2 45072 1 22
2 45073 1 22
2 45074 1 22
2 45075 1 22
2 45076 1 22
2 45077 1 22
2 45078 1 22
2 45079 1 22
2 45080 1 22
2 45081 1 22
2 45082 1 22
2 45083 1 22
2 45084 1 22
2 45085 1 22
2 45086 1 22
2 45087 1 22
2 45088 1 22
2 45089 1 22
2 45090 1 22
2 45091 1 22
2 45092 1 22
2 45093 1 22
2 45094 1 22
2 45095 1 22
2 45096 1 22
2 45097 1 22
2 45098 1 22
2 45099 1 22
2 45100 1 22
2 45101 1 22
2 45102 1 22
2 45103 1 22
2 45104 1 22
2 45105 1 22
2 45106 1 22
2 45107 1 22
2 45108 1 22
2 45109 1 22
2 45110 1 22
2 45111 1 22
2 45112 1 22
2 45113 1 22
2 45114 1 22
2 45115 1 22
2 45116 1 22
2 45117 1 22
2 45118 1 22
2 45119 1 22
2 45120 1 22
2 45121 1 22
2 45122 1 22
2 45123 1 22
2 45124 1 22
2 45125 1 22
2 45126 1 22
2 45127 1 22
2 45128 1 22
2 45129 1 22
2 45130 1 22
1 23 0 209 0
2 45131 1 23
2 45132 1 23
2 45133 1 23
2 45134 1 23
2 45135 1 23
2 45136 1 23
2 45137 1 23
2 45138 1 23
2 45139 1 23
2 45140 1 23
2 45141 1 23
2 45142 1 23
2 45143 1 23
2 45144 1 23
2 45145 1 23
2 45146 1 23
2 45147 1 23
2 45148 1 23
2 45149 1 23
2 45150 1 23
2 45151 1 23
2 45152 1 23
2 45153 1 23
2 45154 1 23
2 45155 1 23
2 45156 1 23
2 45157 1 23
2 45158 1 23
2 45159 1 23
2 45160 1 23
2 45161 1 23
2 45162 1 23
2 45163 1 23
2 45164 1 23
2 45165 1 23
2 45166 1 23
2 45167 1 23
2 45168 1 23
2 45169 1 23
2 45170 1 23
2 45171 1 23
2 45172 1 23
2 45173 1 23
2 45174 1 23
2 45175 1 23
2 45176 1 23
2 45177 1 23
2 45178 1 23
2 45179 1 23
2 45180 1 23
2 45181 1 23
2 45182 1 23
2 45183 1 23
2 45184 1 23
2 45185 1 23
2 45186 1 23
2 45187 1 23
2 45188 1 23
2 45189 1 23
2 45190 1 23
2 45191 1 23
2 45192 1 23
2 45193 1 23
2 45194 1 23
2 45195 1 23
2 45196 1 23
2 45197 1 23
2 45198 1 23
2 45199 1 23
2 45200 1 23
2 45201 1 23
2 45202 1 23
2 45203 1 23
2 45204 1 23
2 45205 1 23
2 45206 1 23
2 45207 1 23
2 45208 1 23
2 45209 1 23
2 45210 1 23
2 45211 1 23
2 45212 1 23
2 45213 1 23
2 45214 1 23
2 45215 1 23
2 45216 1 23
2 45217 1 23
2 45218 1 23
2 45219 1 23
2 45220 1 23
2 45221 1 23
2 45222 1 23
2 45223 1 23
2 45224 1 23
2 45225 1 23
2 45226 1 23
2 45227 1 23
2 45228 1 23
2 45229 1 23
2 45230 1 23
2 45231 1 23
2 45232 1 23
2 45233 1 23
2 45234 1 23
2 45235 1 23
2 45236 1 23
2 45237 1 23
2 45238 1 23
2 45239 1 23
2 45240 1 23
2 45241 1 23
2 45242 1 23
2 45243 1 23
2 45244 1 23
2 45245 1 23
2 45246 1 23
2 45247 1 23
2 45248 1 23
2 45249 1 23
2 45250 1 23
2 45251 1 23
2 45252 1 23
2 45253 1 23
2 45254 1 23
2 45255 1 23
2 45256 1 23
2 45257 1 23
2 45258 1 23
2 45259 1 23
2 45260 1 23
2 45261 1 23
2 45262 1 23
2 45263 1 23
2 45264 1 23
2 45265 1 23
2 45266 1 23
2 45267 1 23
2 45268 1 23
2 45269 1 23
2 45270 1 23
2 45271 1 23
2 45272 1 23
2 45273 1 23
2 45274 1 23
2 45275 1 23
2 45276 1 23
2 45277 1 23
2 45278 1 23
2 45279 1 23
2 45280 1 23
2 45281 1 23
2 45282 1 23
2 45283 1 23
2 45284 1 23
2 45285 1 23
2 45286 1 23
2 45287 1 23
2 45288 1 23
2 45289 1 23
2 45290 1 23
2 45291 1 23
2 45292 1 23
2 45293 1 23
2 45294 1 23
2 45295 1 23
2 45296 1 23
2 45297 1 23
2 45298 1 23
2 45299 1 23
2 45300 1 23
2 45301 1 23
2 45302 1 23
2 45303 1 23
2 45304 1 23
2 45305 1 23
2 45306 1 23
2 45307 1 23
2 45308 1 23
2 45309 1 23
2 45310 1 23
2 45311 1 23
2 45312 1 23
2 45313 1 23
2 45314 1 23
2 45315 1 23
2 45316 1 23
2 45317 1 23
2 45318 1 23
2 45319 1 23
2 45320 1 23
2 45321 1 23
2 45322 1 23
2 45323 1 23
2 45324 1 23
2 45325 1 23
2 45326 1 23
2 45327 1 23
2 45328 1 23
2 45329 1 23
2 45330 1 23
2 45331 1 23
2 45332 1 23
2 45333 1 23
2 45334 1 23
2 45335 1 23
2 45336 1 23
2 45337 1 23
2 45338 1 23
2 45339 1 23
1 24 0 166 0
2 45340 1 24
2 45341 1 24
2 45342 1 24
2 45343 1 24
2 45344 1 24
2 45345 1 24
2 45346 1 24
2 45347 1 24
2 45348 1 24
2 45349 1 24
2 45350 1 24
2 45351 1 24
2 45352 1 24
2 45353 1 24
2 45354 1 24
2 45355 1 24
2 45356 1 24
2 45357 1 24
2 45358 1 24
2 45359 1 24
2 45360 1 24
2 45361 1 24
2 45362 1 24
2 45363 1 24
2 45364 1 24
2 45365 1 24
2 45366 1 24
2 45367 1 24
2 45368 1 24
2 45369 1 24
2 45370 1 24
2 45371 1 24
2 45372 1 24
2 45373 1 24
2 45374 1 24
2 45375 1 24
2 45376 1 24
2 45377 1 24
2 45378 1 24
2 45379 1 24
2 45380 1 24
2 45381 1 24
2 45382 1 24
2 45383 1 24
2 45384 1 24
2 45385 1 24
2 45386 1 24
2 45387 1 24
2 45388 1 24
2 45389 1 24
2 45390 1 24
2 45391 1 24
2 45392 1 24
2 45393 1 24
2 45394 1 24
2 45395 1 24
2 45396 1 24
2 45397 1 24
2 45398 1 24
2 45399 1 24
2 45400 1 24
2 45401 1 24
2 45402 1 24
2 45403 1 24
2 45404 1 24
2 45405 1 24
2 45406 1 24
2 45407 1 24
2 45408 1 24
2 45409 1 24
2 45410 1 24
2 45411 1 24
2 45412 1 24
2 45413 1 24
2 45414 1 24
2 45415 1 24
2 45416 1 24
2 45417 1 24
2 45418 1 24
2 45419 1 24
2 45420 1 24
2 45421 1 24
2 45422 1 24
2 45423 1 24
2 45424 1 24
2 45425 1 24
2 45426 1 24
2 45427 1 24
2 45428 1 24
2 45429 1 24
2 45430 1 24
2 45431 1 24
2 45432 1 24
2 45433 1 24
2 45434 1 24
2 45435 1 24
2 45436 1 24
2 45437 1 24
2 45438 1 24
2 45439 1 24
2 45440 1 24
2 45441 1 24
2 45442 1 24
2 45443 1 24
2 45444 1 24
2 45445 1 24
2 45446 1 24
2 45447 1 24
2 45448 1 24
2 45449 1 24
2 45450 1 24
2 45451 1 24
2 45452 1 24
2 45453 1 24
2 45454 1 24
2 45455 1 24
2 45456 1 24
2 45457 1 24
2 45458 1 24
2 45459 1 24
2 45460 1 24
2 45461 1 24
2 45462 1 24
2 45463 1 24
2 45464 1 24
2 45465 1 24
2 45466 1 24
2 45467 1 24
2 45468 1 24
2 45469 1 24
2 45470 1 24
2 45471 1 24
2 45472 1 24
2 45473 1 24
2 45474 1 24
2 45475 1 24
2 45476 1 24
2 45477 1 24
2 45478 1 24
2 45479 1 24
2 45480 1 24
2 45481 1 24
2 45482 1 24
2 45483 1 24
2 45484 1 24
2 45485 1 24
2 45486 1 24
2 45487 1 24
2 45488 1 24
2 45489 1 24
2 45490 1 24
2 45491 1 24
2 45492 1 24
2 45493 1 24
2 45494 1 24
2 45495 1 24
2 45496 1 24
2 45497 1 24
2 45498 1 24
2 45499 1 24
2 45500 1 24
2 45501 1 24
2 45502 1 24
2 45503 1 24
2 45504 1 24
2 45505 1 24
2 45506 1 27
2 45507 1 27
2 45508 1 27
2 45509 1 27
2 45510 1 27
2 45511 1 27
2 45512 1 27
2 45513 1 27
2 45514 1 27
2 45515 1 27
2 45516 1 27
2 45517 1 27
2 45518 1 27
2 45519 1 27
2 45520 1 27
2 45521 1 27
2 45522 1 27
2 45523 1 27
2 45524 1 27
2 45525 1 27
2 45526 1 27
2 45527 1 27
2 45528 1 27
2 45529 1 27
2 45530 1 27
2 45531 1 27
2 45532 1 27
2 45533 1 27
2 45534 1 27
2 45535 1 27
2 45536 1 27
2 45537 1 27
2 45538 1 27
2 45539 1 27
2 45540 1 27
2 45541 1 27
2 45542 1 27
2 45543 1 27
2 45544 1 27
2 45545 1 27
2 45546 1 27
2 45547 1 27
2 45548 1 27
2 45549 1 27
2 45550 1 27
2 45551 1 27
2 45552 1 27
2 45553 1 27
2 45554 1 27
2 45555 1 27
2 45556 1 27
2 45557 1 27
2 45558 1 27
2 45559 1 27
2 45560 1 27
2 45561 1 27
2 45562 1 27
2 45563 1 27
2 45564 1 27
2 45565 1 27
2 45566 1 27
2 45567 1 27
2 45568 1 27
2 45569 1 27
2 45570 1 27
2 45571 1 27
2 45572 1 27
2 45573 1 27
2 45574 1 27
2 45575 1 27
2 45576 1 27
2 45577 1 27
2 45578 1 27
2 45579 1 27
2 45580 1 27
2 45581 1 27
2 45582 1 27
2 45583 1 27
2 45584 1 27
2 45585 1 27
2 45586 1 27
2 45587 1 27
2 45588 1 27
2 45589 1 27
2 45590 1 27
2 45591 1 27
2 45592 1 27
2 45593 1 27
2 45594 1 27
2 45595 1 27
2 45596 1 27
2 45597 1 27
2 45598 1 27
2 45599 1 27
2 45600 1 27
2 45601 1 27
2 45602 1 27
2 45603 1 27
2 45604 1 27
2 45605 1 27
2 45606 1 27
2 45607 1 27
2 45608 1 27
2 45609 1 27
2 45610 1 27
2 45611 1 27
2 45612 1 27
2 45613 1 27
2 45614 1 27
2 45615 1 27
2 45616 1 27
2 45617 1 27
2 45618 1 27
2 45619 1 27
2 45620 1 27
2 45621 1 27
2 45622 1 27
2 45623 1 27
2 45624 1 27
2 45625 1 27
2 45626 1 27
2 45627 1 27
2 45628 1 27
2 45629 1 27
2 45630 1 27
2 45631 1 27
2 45632 1 27
2 45633 1 27
2 45634 1 27
2 45635 1 27
2 45636 1 27
2 45637 1 27
2 45638 1 27
2 45639 1 27
2 45640 1 27
2 45641 1 27
2 45642 1 27
2 45643 1 27
2 45644 1 27
2 45645 1 27
2 45646 1 27
2 45647 1 27
2 45648 1 27
2 45649 1 27
2 45650 1 27
2 45651 1 27
2 45652 1 27
2 45653 1 27
2 45654 1 27
2 45655 1 27
2 45656 1 27
2 45657 1 27
2 45658 1 27
2 45659 1 27
2 45660 1 28
2 45661 1 28
2 45662 1 28
2 45663 1 28
2 45664 1 28
2 45665 1 28
2 45666 1 28
2 45667 1 28
2 45668 1 28
2 45669 1 28
2 45670 1 28
2 45671 1 28
2 45672 1 28
2 45673 1 28
2 45674 1 28
2 45675 1 28
2 45676 1 28
2 45677 1 28
2 45678 1 28
2 45679 1 28
2 45680 1 28
2 45681 1 28
2 45682 1 28
2 45683 1 28
2 45684 1 28
2 45685 1 28
2 45686 1 28
2 45687 1 28
2 45688 1 28
2 45689 1 28
2 45690 1 28
2 45691 1 28
2 45692 1 28
2 45693 1 28
2 45694 1 28
2 45695 1 28
2 45696 1 28
2 45697 1 28
2 45698 1 28
2 45699 1 28
2 45700 1 28
2 45701 1 28
2 45702 1 28
2 45703 1 28
2 45704 1 28
2 45705 1 28
2 45706 1 28
2 45707 1 28
2 45708 1 28
2 45709 1 28
2 45710 1 28
2 45711 1 28
2 45712 1 28
2 45713 1 28
2 45714 1 28
2 45715 1 28
2 45716 1 28
2 45717 1 28
2 45718 1 28
2 45719 1 28
2 45720 1 28
2 45721 1 28
2 45722 1 28
2 45723 1 28
2 45724 1 28
2 45725 1 28
2 45726 1 28
2 45727 1 28
2 45728 1 28
2 45729 1 28
2 45730 1 28
2 45731 1 28
2 45732 1 28
2 45733 1 28
2 45734 1 28
2 45735 1 28
2 45736 1 28
2 45737 1 28
2 45738 1 28
2 45739 1 28
2 45740 1 28
2 45741 1 28
2 45742 1 28
2 45743 1 28
2 45744 1 28
2 45745 1 28
2 45746 1 28
2 45747 1 28
2 45748 1 28
2 45749 1 28
2 45750 1 28
2 45751 1 28
2 45752 1 28
2 45753 1 28
2 45754 1 28
2 45755 1 28
2 45756 1 28
2 45757 1 28
2 45758 1 28
2 45759 1 28
2 45760 1 28
2 45761 1 28
2 45762 1 28
2 45763 1 28
2 45764 1 28
2 45765 1 28
2 45766 1 28
2 45767 1 28
2 45768 1 28
2 45769 1 28
2 45770 1 28
2 45771 1 28
2 45772 1 28
2 45773 1 28
2 45774 1 28
2 45775 1 28
2 45776 1 28
2 45777 1 28
2 45778 1 28
2 45779 1 28
2 45780 1 28
2 45781 1 28
2 45782 1 29
2 45783 1 29
2 45784 1 29
2 45785 1 29
2 45786 1 29
2 45787 1 29
2 45788 1 29
2 45789 1 29
2 45790 1 29
2 45791 1 29
2 45792 1 29
2 45793 1 29
2 45794 1 29
2 45795 1 29
2 45796 1 29
2 45797 1 29
2 45798 1 29
2 45799 1 29
2 45800 1 29
2 45801 1 29
2 45802 1 29
2 45803 1 29
2 45804 1 29
2 45805 1 29
2 45806 1 29
2 45807 1 29
2 45808 1 29
2 45809 1 29
2 45810 1 29
2 45811 1 29
2 45812 1 29
2 45813 1 29
2 45814 1 29
2 45815 1 29
2 45816 1 29
2 45817 1 29
2 45818 1 29
2 45819 1 29
2 45820 1 29
2 45821 1 29
2 45822 1 29
2 45823 1 29
2 45824 1 29
2 45825 1 29
2 45826 1 29
2 45827 1 29
2 45828 1 29
2 45829 1 29
2 45830 1 29
2 45831 1 29
2 45832 1 29
2 45833 1 29
2 45834 1 29
2 45835 1 29
2 45836 1 29
2 45837 1 29
2 45838 1 29
2 45839 1 29
2 45840 1 29
2 45841 1 29
2 45842 1 29
2 45843 1 29
2 45844 1 29
2 45845 1 29
2 45846 1 29
2 45847 1 29
2 45848 1 29
2 45849 1 29
2 45850 1 29
2 45851 1 29
2 45852 1 29
2 45853 1 29
2 45854 1 29
2 45855 1 29
2 45856 1 29
2 45857 1 29
2 45858 1 29
2 45859 1 29
2 45860 1 29
2 45861 1 29
2 45862 1 29
2 45863 1 29
2 45864 1 29
2 45865 1 29
2 45866 1 29
2 45867 1 29
2 45868 1 29
2 45869 1 29
2 45870 1 29
2 45871 1 29
2 45872 1 29
2 45873 1 29
2 45874 1 29
2 45875 1 29
2 45876 1 29
2 45877 1 29
2 45878 1 29
2 45879 1 30
2 45880 1 30
2 45881 1 30
2 45882 1 30
2 45883 1 30
2 45884 1 30
2 45885 1 30
2 45886 1 30
2 45887 1 30
2 45888 1 30
2 45889 1 30
2 45890 1 30
2 45891 1 30
2 45892 1 30
2 45893 1 30
2 45894 1 30
2 45895 1 30
2 45896 1 30
2 45897 1 30
2 45898 1 30
2 45899 1 30
2 45900 1 30
2 45901 1 30
2 45902 1 30
2 45903 1 30
2 45904 1 30
2 45905 1 30
2 45906 1 30
2 45907 1 30
2 45908 1 30
2 45909 1 30
2 45910 1 30
2 45911 1 30
2 45912 1 30
2 45913 1 30
2 45914 1 30
2 45915 1 30
2 45916 1 30
2 45917 1 30
2 45918 1 30
2 45919 1 30
2 45920 1 30
2 45921 1 30
2 45922 1 31
2 45923 1 31
2 45924 1 31
2 45925 1 31
2 45926 1 31
2 45927 1 31
2 45928 1 31
2 45929 1 31
2 45930 1 31
2 45931 1 31
2 45932 1 31
2 45933 1 31
2 45934 1 31
2 45935 1 31
2 45936 1 31
2 45937 1 31
2 45938 1 31
2 45939 1 31
2 45940 1 31
2 45941 1 31
2 45942 1 31
2 45943 1 31
2 45944 1 31
2 45945 1 31
2 45946 1 31
2 45947 1 31
2 45948 1 31
2 45949 1 31
2 45950 1 31
2 45951 1 31
2 45952 1 31
2 45953 1 31
2 45954 1 31
2 45955 1 31
2 45956 1 31
2 45957 1 31
2 45958 1 31
2 45959 1 31
2 45960 1 31
2 45961 1 31
2 45962 1 31
2 45963 1 31
2 45964 1 31
2 45965 1 31
2 45966 1 31
2 45967 1 31
2 45968 1 31
2 45969 1 31
2 45970 1 31
2 45971 1 31
2 45972 1 31
2 45973 1 31
2 45974 1 31
2 45975 1 31
2 45976 1 31
2 45977 1 31
2 45978 1 31
2 45979 1 31
2 45980 1 31
2 45981 1 31
2 45982 1 31
2 45983 1 31
2 45984 1 31
2 45985 1 31
2 45986 1 31
2 45987 1 31
2 45988 1 31
2 45989 1 31
2 45990 1 31
2 45991 1 31
2 45992 1 31
2 45993 1 31
2 45994 1 31
2 45995 1 31
2 45996 1 31
2 45997 1 31
2 45998 1 31
2 45999 1 31
2 46000 1 31
2 46001 1 31
2 46002 1 31
2 46003 1 31
2 46004 1 31
2 46005 1 31
2 46006 1 31
2 46007 1 31
2 46008 1 31
2 46009 1 31
2 46010 1 31
2 46011 1 31
2 46012 1 31
2 46013 1 31
2 46014 1 31
2 46015 1 31
2 46016 1 31
2 46017 1 31
2 46018 1 31
2 46019 1 31
2 46020 1 31
2 46021 1 31
2 46022 1 31
2 46023 1 31
2 46024 1 31
2 46025 1 31
2 46026 1 31
2 46027 1 31
2 46028 1 31
2 46029 1 31
2 46030 1 31
2 46031 1 31
2 46032 1 31
2 46033 1 31
2 46034 1 31
2 46035 1 31
2 46036 1 31
2 46037 1 31
2 46038 1 31
2 46039 1 31
2 46040 1 31
2 46041 1 31
2 46042 1 31
2 46043 1 31
2 46044 1 31
2 46045 1 31
2 46046 1 31
2 46047 1 31
2 46048 1 31
2 46049 1 31
2 46050 1 31
2 46051 1 31
2 46052 1 31
2 46053 1 31
2 46054 1 31
2 46055 1 31
2 46056 1 31
2 46057 1 31
2 46058 1 31
2 46059 1 31
2 46060 1 31
2 46061 1 31
2 46062 1 31
2 46063 1 31
2 46064 1 31
2 46065 1 31
2 46066 1 31
2 46067 1 31
2 46068 1 31
2 46069 1 31
2 46070 1 31
2 46071 1 31
2 46072 1 31
2 46073 1 31
2 46074 1 31
2 46075 1 31
2 46076 1 31
2 46077 1 31
2 46078 1 31
2 46079 1 31
2 46080 1 31
2 46081 1 31
2 46082 1 31
2 46083 1 31
2 46084 1 31
2 46085 1 31
2 46086 1 31
2 46087 1 31
2 46088 1 31
2 46089 1 31
2 46090 1 31
2 46091 1 31
2 46092 1 31
2 46093 1 31
2 46094 1 31
2 46095 1 31
2 46096 1 31
2 46097 1 31
2 46098 1 31
2 46099 1 31
2 46100 1 31
2 46101 1 31
2 46102 1 31
2 46103 1 31
2 46104 1 31
2 46105 1 31
2 46106 1 32
2 46107 1 32
2 46108 1 32
2 46109 1 32
2 46110 1 32
2 46111 1 32
2 46112 1 32
2 46113 1 32
2 46114 1 32
2 46115 1 32
2 46116 1 32
2 46117 1 32
2 46118 1 32
2 46119 1 32
2 46120 1 32
2 46121 1 32
2 46122 1 32
2 46123 1 32
2 46124 1 32
2 46125 1 32
2 46126 1 32
2 46127 1 32
2 46128 1 32
2 46129 1 32
2 46130 1 32
2 46131 1 32
2 46132 1 32
2 46133 1 32
2 46134 1 32
2 46135 1 32
2 46136 1 32
2 46137 1 32
2 46138 1 32
2 46139 1 32
2 46140 1 32
2 46141 1 32
2 46142 1 32
2 46143 1 32
2 46144 1 32
2 46145 1 32
2 46146 1 32
2 46147 1 32
2 46148 1 32
2 46149 1 32
2 46150 1 32
2 46151 1 32
2 46152 1 32
2 46153 1 32
2 46154 1 32
2 46155 1 32
2 46156 1 32
2 46157 1 32
2 46158 1 32
2 46159 1 32
2 46160 1 32
2 46161 1 32
2 46162 1 32
2 46163 1 32
2 46164 1 32
2 46165 1 32
2 46166 1 32
2 46167 1 32
2 46168 1 32
2 46169 1 32
2 46170 1 32
2 46171 1 32
2 46172 1 32
2 46173 1 32
2 46174 1 32
2 46175 1 32
2 46176 1 32
2 46177 1 32
2 46178 1 32
2 46179 1 32
2 46180 1 32
2 46181 1 32
2 46182 1 32
2 46183 1 32
2 46184 1 32
2 46185 1 32
2 46186 1 32
2 46187 1 32
2 46188 1 32
2 46189 1 32
2 46190 1 32
2 46191 1 32
2 46192 1 32
2 46193 1 32
2 46194 1 32
2 46195 1 32
2 46196 1 32
2 46197 1 32
2 46198 1 32
2 46199 1 32
2 46200 1 32
2 46201 1 32
2 46202 1 32
2 46203 1 32
2 46204 1 32
2 46205 1 32
2 46206 1 32
2 46207 1 32
2 46208 1 32
2 46209 1 32
2 46210 1 32
2 46211 1 32
2 46212 1 32
2 46213 1 32
2 46214 1 32
2 46215 1 32
2 46216 1 32
2 46217 1 32
2 46218 1 32
2 46219 1 32
2 46220 1 32
2 46221 1 32
2 46222 1 32
2 46223 1 32
2 46224 1 32
2 46225 1 32
2 46226 1 32
2 46227 1 32
2 46228 1 32
2 46229 1 32
2 46230 1 32
2 46231 1 32
2 46232 1 32
2 46233 1 32
2 46234 1 32
2 46235 1 32
2 46236 1 32
2 46237 1 32
2 46238 1 32
2 46239 1 32
2 46240 1 32
2 46241 1 32
2 46242 1 32
2 46243 1 32
2 46244 1 32
2 46245 1 32
2 46246 1 32
2 46247 1 32
2 46248 1 32
2 46249 1 32
2 46250 1 32
2 46251 1 32
2 46252 1 32
2 46253 1 32
2 46254 1 32
2 46255 1 32
2 46256 1 32
2 46257 1 32
2 46258 1 32
2 46259 1 32
2 46260 1 32
2 46261 1 32
2 46262 1 32
2 46263 1 32
2 46264 1 32
2 46265 1 32
2 46266 1 32
2 46267 1 32
2 46268 1 32
2 46269 1 32
2 46270 1 32
2 46271 1 32
2 46272 1 32
2 46273 1 32
2 46274 1 32
2 46275 1 32
2 46276 1 32
2 46277 1 32
2 46278 1 32
2 46279 1 32
2 46280 1 32
2 46281 1 32
2 46282 1 32
2 46283 1 32
2 46284 1 32
2 46285 1 32
2 46286 1 32
2 46287 1 32
2 46288 1 32
2 46289 1 32
2 46290 1 32
2 46291 1 32
2 46292 1 32
2 46293 1 32
2 46294 1 32
2 46295 1 32
2 46296 1 32
2 46297 1 32
2 46298 1 32
2 46299 1 32
2 46300 1 32
2 46301 1 32
2 46302 1 32
2 46303 1 32
2 46304 1 32
2 46305 1 32
2 46306 1 32
2 46307 1 32
2 46308 1 32
2 46309 1 32
2 46310 1 32
2 46311 1 32
2 46312 1 32
2 46313 1 32
2 46314 1 32
2 46315 1 32
2 46316 1 32
2 46317 1 32
2 46318 1 32
2 46319 1 32
2 46320 1 32
2 46321 1 32
2 46322 1 32
2 46323 1 32
2 46324 1 32
2 46325 1 32
2 46326 1 32
2 46327 1 32
2 46328 1 32
2 46329 1 32
2 46330 1 32
2 46331 1 32
2 46332 1 32
2 46333 1 32
2 46334 1 32
2 46335 1 32
2 46336 1 32
2 46337 1 32
2 46338 1 32
2 46339 1 32
2 46340 1 32
2 46341 1 32
2 46342 1 32
2 46343 1 32
2 46344 1 32
2 46345 1 32
2 46346 1 32
2 46347 1 32
2 46348 1 32
2 46349 1 32
2 46350 1 32
2 46351 1 32
2 46352 1 32
2 46353 1 32
2 46354 1 32
2 46355 1 32
2 46356 1 32
2 46357 1 32
2 46358 1 32
2 46359 1 32
2 46360 1 32
2 46361 1 32
2 46362 1 32
2 46363 1 32
2 46364 1 33
2 46365 1 33
2 46366 1 33
2 46367 1 33
2 46368 1 33
2 46369 1 33
2 46370 1 33
2 46371 1 33
2 46372 1 33
2 46373 1 33
2 46374 1 33
2 46375 1 33
2 46376 1 33
2 46377 1 33
2 46378 1 33
2 46379 1 33
2 46380 1 33
2 46381 1 33
2 46382 1 33
2 46383 1 33
2 46384 1 33
2 46385 1 33
2 46386 1 33
2 46387 1 33
2 46388 1 33
2 46389 1 33
2 46390 1 33
2 46391 1 33
2 46392 1 33
2 46393 1 33
2 46394 1 33
2 46395 1 33
2 46396 1 33
2 46397 1 33
2 46398 1 33
2 46399 1 33
2 46400 1 33
2 46401 1 33
2 46402 1 33
2 46403 1 33
2 46404 1 33
2 46405 1 33
2 46406 1 33
2 46407 1 33
2 46408 1 33
2 46409 1 33
2 46410 1 33
2 46411 1 33
2 46412 1 33
2 46413 1 33
2 46414 1 33
2 46415 1 33
2 46416 1 33
2 46417 1 33
2 46418 1 33
2 46419 1 33
2 46420 1 33
2 46421 1 33
2 46422 1 33
2 46423 1 33
2 46424 1 33
2 46425 1 33
2 46426 1 33
2 46427 1 33
2 46428 1 33
2 46429 1 33
2 46430 1 33
2 46431 1 33
2 46432 1 33
2 46433 1 33
2 46434 1 33
2 46435 1 33
2 46436 1 33
2 46437 1 33
2 46438 1 33
2 46439 1 33
2 46440 1 33
2 46441 1 33
2 46442 1 33
2 46443 1 33
2 46444 1 33
2 46445 1 33
2 46446 1 33
2 46447 1 33
2 46448 1 33
2 46449 1 33
2 46450 1 33
2 46451 1 33
2 46452 1 33
2 46453 1 33
2 46454 1 33
2 46455 1 33
2 46456 1 33
2 46457 1 33
2 46458 1 33
2 46459 1 33
2 46460 1 33
2 46461 1 33
2 46462 1 33
2 46463 1 33
2 46464 1 33
2 46465 1 33
2 46466 1 33
2 46467 1 33
2 46468 1 33
2 46469 1 33
2 46470 1 33
2 46471 1 33
2 46472 1 33
2 46473 1 33
2 46474 1 33
2 46475 1 33
2 46476 1 33
2 46477 1 33
2 46478 1 33
2 46479 1 33
2 46480 1 33
2 46481 1 33
2 46482 1 33
2 46483 1 33
2 46484 1 33
2 46485 1 33
2 46486 1 33
2 46487 1 33
2 46488 1 33
2 46489 1 33
2 46490 1 33
2 46491 1 33
2 46492 1 33
2 46493 1 33
2 46494 1 33
2 46495 1 33
2 46496 1 33
2 46497 1 33
2 46498 1 33
2 46499 1 33
2 46500 1 33
2 46501 1 33
2 46502 1 33
2 46503 1 33
2 46504 1 33
2 46505 1 33
2 46506 1 33
2 46507 1 33
2 46508 1 33
2 46509 1 33
2 46510 1 33
2 46511 1 33
2 46512 1 33
2 46513 1 33
2 46514 1 33
2 46515 1 33
2 46516 1 33
2 46517 1 33
2 46518 1 33
2 46519 1 33
2 46520 1 33
2 46521 1 33
2 46522 1 33
2 46523 1 33
2 46524 1 33
2 46525 1 33
2 46526 1 33
2 46527 1 33
2 46528 1 33
2 46529 1 33
2 46530 1 33
2 46531 1 33
2 46532 1 33
2 46533 1 33
2 46534 1 33
2 46535 1 33
2 46536 1 33
2 46537 1 33
2 46538 1 33
2 46539 1 33
2 46540 1 33
2 46541 1 33
2 46542 1 33
2 46543 1 33
2 46544 1 33
2 46545 1 33
2 46546 1 33
2 46547 1 33
2 46548 1 33
2 46549 1 33
2 46550 1 33
2 46551 1 33
2 46552 1 33
2 46553 1 33
2 46554 1 33
2 46555 1 33
2 46556 1 33
2 46557 1 33
2 46558 1 33
2 46559 1 33
2 46560 1 33
2 46561 1 33
2 46562 1 33
2 46563 1 33
2 46564 1 33
2 46565 1 33
2 46566 1 33
2 46567 1 33
2 46568 1 33
2 46569 1 33
2 46570 1 33
2 46571 1 33
2 46572 1 33
2 46573 1 33
2 46574 1 33
2 46575 1 33
2 46576 1 33
2 46577 1 34
2 46578 1 34
2 46579 1 34
2 46580 1 34
2 46581 1 34
2 46582 1 34
2 46583 1 34
2 46584 1 34
2 46585 1 34
2 46586 1 34
2 46587 1 34
2 46588 1 34
2 46589 1 34
2 46590 1 34
2 46591 1 34
2 46592 1 34
2 46593 1 34
2 46594 1 34
2 46595 1 34
2 46596 1 34
2 46597 1 34
2 46598 1 34
2 46599 1 34
2 46600 1 34
2 46601 1 34
2 46602 1 34
2 46603 1 34
2 46604 1 34
2 46605 1 34
2 46606 1 34
2 46607 1 34
2 46608 1 34
2 46609 1 34
2 46610 1 34
2 46611 1 34
2 46612 1 34
2 46613 1 34
2 46614 1 34
2 46615 1 34
2 46616 1 34
2 46617 1 34
2 46618 1 34
2 46619 1 34
2 46620 1 34
2 46621 1 34
2 46622 1 34
2 46623 1 34
2 46624 1 34
2 46625 1 34
2 46626 1 34
2 46627 1 34
2 46628 1 34
2 46629 1 34
2 46630 1 34
2 46631 1 34
2 46632 1 34
2 46633 1 34
2 46634 1 34
2 46635 1 34
2 46636 1 34
2 46637 1 34
2 46638 1 34
2 46639 1 34
2 46640 1 34
2 46641 1 34
2 46642 1 34
2 46643 1 34
2 46644 1 34
2 46645 1 34
2 46646 1 34
2 46647 1 34
2 46648 1 34
2 46649 1 34
2 46650 1 34
2 46651 1 34
2 46652 1 34
2 46653 1 34
2 46654 1 34
2 46655 1 34
2 46656 1 34
2 46657 1 34
2 46658 1 34
2 46659 1 34
2 46660 1 34
2 46661 1 34
2 46662 1 34
2 46663 1 34
2 46664 1 34
2 46665 1 34
2 46666 1 34
2 46667 1 34
2 46668 1 34
2 46669 1 34
2 46670 1 34
2 46671 1 34
2 46672 1 34
2 46673 1 34
2 46674 1 34
2 46675 1 34
2 46676 1 34
2 46677 1 34
2 46678 1 34
2 46679 1 34
2 46680 1 34
2 46681 1 34
2 46682 1 34
2 46683 1 34
2 46684 1 34
2 46685 1 34
2 46686 1 34
2 46687 1 34
2 46688 1 34
2 46689 1 34
2 46690 1 34
2 46691 1 34
2 46692 1 34
2 46693 1 34
2 46694 1 34
2 46695 1 34
2 46696 1 34
2 46697 1 34
2 46698 1 34
2 46699 1 34
2 46700 1 34
2 46701 1 34
2 46702 1 34
2 46703 1 34
2 46704 1 34
2 46705 1 34
2 46706 1 34
2 46707 1 34
2 46708 1 34
2 46709 1 34
2 46710 1 34
2 46711 1 34
2 46712 1 34
2 46713 1 34
2 46714 1 34
2 46715 1 34
2 46716 1 34
2 46717 1 34
2 46718 1 34
2 46719 1 34
2 46720 1 34
2 46721 1 34
2 46722 1 34
2 46723 1 34
2 46724 1 34
2 46725 1 34
2 46726 1 34
2 46727 1 34
2 46728 1 34
2 46729 1 34
2 46730 1 34
2 46731 1 34
2 46732 1 34
2 46733 1 34
2 46734 1 34
2 46735 1 34
2 46736 1 34
2 46737 1 34
2 46738 1 34
2 46739 1 34
2 46740 1 34
2 46741 1 34
2 46742 1 34
2 46743 1 34
2 46744 1 34
2 46745 1 34
2 46746 1 34
2 46747 1 34
2 46748 1 34
2 46749 1 34
2 46750 1 34
2 46751 1 34
2 46752 1 34
2 46753 1 34
2 46754 1 34
2 46755 1 34
2 46756 1 34
2 46757 1 34
2 46758 1 34
2 46759 1 34
2 46760 1 34
2 46761 1 34
2 46762 1 34
2 46763 1 34
2 46764 1 34
2 46765 1 34
2 46766 1 34
2 46767 1 34
2 46768 1 34
2 46769 1 34
2 46770 1 34
2 46771 1 34
2 46772 1 34
2 46773 1 34
2 46774 1 34
2 46775 1 34
2 46776 1 34
2 46777 1 34
2 46778 1 34
2 46779 1 34
2 46780 1 34
2 46781 1 35
2 46782 1 35
2 46783 1 35
2 46784 1 35
2 46785 1 35
2 46786 1 35
2 46787 1 35
2 46788 1 35
2 46789 1 35
2 46790 1 35
2 46791 1 35
2 46792 1 35
2 46793 1 35
2 46794 1 35
2 46795 1 35
2 46796 1 35
2 46797 1 35
2 46798 1 35
2 46799 1 35
2 46800 1 35
2 46801 1 35
2 46802 1 35
2 46803 1 35
2 46804 1 35
2 46805 1 35
2 46806 1 35
2 46807 1 35
2 46808 1 35
2 46809 1 35
2 46810 1 35
2 46811 1 35
2 46812 1 35
2 46813 1 35
2 46814 1 35
2 46815 1 35
2 46816 1 35
2 46817 1 35
2 46818 1 35
2 46819 1 35
2 46820 1 35
2 46821 1 35
2 46822 1 35
2 46823 1 35
2 46824 1 35
2 46825 1 35
2 46826 1 35
2 46827 1 35
2 46828 1 35
2 46829 1 35
2 46830 1 35
2 46831 1 35
2 46832 1 35
2 46833 1 35
2 46834 1 35
2 46835 1 35
2 46836 1 35
2 46837 1 35
2 46838 1 35
2 46839 1 35
2 46840 1 35
2 46841 1 35
2 46842 1 35
2 46843 1 35
2 46844 1 35
2 46845 1 35
2 46846 1 35
2 46847 1 35
2 46848 1 35
2 46849 1 35
2 46850 1 35
2 46851 1 35
2 46852 1 35
2 46853 1 35
2 46854 1 35
2 46855 1 35
2 46856 1 35
2 46857 1 35
2 46858 1 35
2 46859 1 35
2 46860 1 35
2 46861 1 35
2 46862 1 35
2 46863 1 35
2 46864 1 35
2 46865 1 35
2 46866 1 35
2 46867 1 35
2 46868 1 35
2 46869 1 35
2 46870 1 36
2 46871 1 36
2 46872 1 36
2 46873 1 36
2 46874 1 36
2 46875 1 36
2 46876 1 36
2 46877 1 36
2 46878 1 36
2 46879 1 36
2 46880 1 36
2 46881 1 36
2 46882 1 36
2 46883 1 36
2 46884 1 36
2 46885 1 36
2 46886 1 36
2 46887 1 36
2 46888 1 36
2 46889 1 36
2 46890 1 36
2 46891 1 36
2 46892 1 36
2 46893 1 36
2 46894 1 36
2 46895 1 36
2 46896 1 36
2 46897 1 36
2 46898 1 36
2 46899 1 36
2 46900 1 36
2 46901 1 36
2 46902 1 36
2 46903 1 36
2 46904 1 36
2 46905 1 36
2 46906 1 36
2 46907 1 36
2 46908 1 36
2 46909 1 36
2 46910 1 36
2 46911 1 36
2 46912 1 36
2 46913 1 36
2 46914 1 36
2 46915 1 36
2 46916 1 36
2 46917 1 36
2 46918 1 36
2 46919 1 36
2 46920 1 36
2 46921 1 36
2 46922 1 36
2 46923 1 36
2 46924 1 36
2 46925 1 36
2 46926 1 36
2 46927 1 36
2 46928 1 36
2 46929 1 36
2 46930 1 36
2 46931 1 36
2 46932 1 36
2 46933 1 36
2 46934 1 36
2 46935 1 36
2 46936 1 36
2 46937 1 36
2 46938 1 36
2 46939 1 36
2 46940 1 36
2 46941 1 36
2 46942 1 36
2 46943 1 36
2 46944 1 36
2 46945 1 36
2 46946 1 36
2 46947 1 36
2 46948 1 36
2 46949 1 36
2 46950 1 37
2 46951 1 37
2 46952 1 37
2 46953 1 37
2 46954 1 37
2 46955 1 37
2 46956 1 37
2 46957 1 37
2 46958 1 37
2 46959 1 37
2 46960 1 37
2 46961 1 37
2 46962 1 37
2 46963 1 37
2 46964 1 37
2 46965 1 37
2 46966 1 37
2 46967 1 37
2 46968 1 37
2 46969 1 37
2 46970 1 37
2 46971 1 37
2 46972 1 37
2 46973 1 37
2 46974 1 37
2 46975 1 37
2 46976 1 37
2 46977 1 37
2 46978 1 37
2 46979 1 37
2 46980 1 37
2 46981 1 37
2 46982 1 37
2 46983 1 37
2 46984 1 37
2 46985 1 37
2 46986 1 37
2 46987 1 37
2 46988 1 37
2 46989 1 37
2 46990 1 37
2 46991 1 37
2 46992 1 37
2 46993 1 37
2 46994 1 37
2 46995 1 37
2 46996 1 38
2 46997 1 38
2 46998 1 38
2 46999 1 38
2 47000 1 38
2 47001 1 38
2 47002 1 38
2 47003 1 38
2 47004 1 38
2 47005 1 38
2 47006 1 38
2 47007 1 38
2 47008 1 38
2 47009 1 38
2 47010 1 38
2 47011 1 38
2 47012 1 38
2 47013 1 38
2 47014 1 38
2 47015 1 38
2 47016 1 38
2 47017 1 38
2 47018 1 38
2 47019 1 38
2 47020 1 38
2 47021 1 38
2 47022 1 38
2 47023 1 38
2 47024 1 38
2 47025 1 38
2 47026 1 38
2 47027 1 38
2 47028 1 38
2 47029 1 38
2 47030 1 38
2 47031 1 38
2 47032 1 38
2 47033 1 39
2 47034 1 39
2 47035 1 39
2 47036 1 39
2 47037 1 39
2 47038 1 39
2 47039 1 39
2 47040 1 39
2 47041 1 39
2 47042 1 39
2 47043 1 39
2 47044 1 39
2 47045 1 39
2 47046 1 39
2 47047 1 39
2 47048 1 39
2 47049 1 39
2 47050 1 39
2 47051 1 39
2 47052 1 39
2 47053 1 39
2 47054 1 39
2 47055 1 39
2 47056 1 39
2 47057 1 39
2 47058 1 39
2 47059 1 39
2 47060 1 39
2 47061 1 39
2 47062 1 39
2 47063 1 39
2 47064 1 39
2 47065 1 39
2 47066 1 39
2 47067 1 39
2 47068 1 39
2 47069 1 39
2 47070 1 39
2 47071 1 39
2 47072 1 39
2 47073 1 39
2 47074 1 39
2 47075 1 39
2 47076 1 39
2 47077 1 39
2 47078 1 39
2 47079 1 39
2 47080 1 39
2 47081 1 39
2 47082 1 39
2 47083 1 39
2 47084 1 39
2 47085 1 39
2 47086 1 39
2 47087 1 39
2 47088 1 39
2 47089 1 39
2 47090 1 39
2 47091 1 39
2 47092 1 39
2 47093 1 39
2 47094 1 39
2 47095 1 39
2 47096 1 39
2 47097 1 39
2 47098 1 39
2 47099 1 39
2 47100 1 39
2 47101 1 39
2 47102 1 39
2 47103 1 39
2 47104 1 39
2 47105 1 39
2 47106 1 39
2 47107 1 39
2 47108 1 39
2 47109 1 39
2 47110 1 39
2 47111 1 39
2 47112 1 39
2 47113 1 39
2 47114 1 39
2 47115 1 39
2 47116 1 39
2 47117 1 39
2 47118 1 39
2 47119 1 39
2 47120 1 39
2 47121 1 39
2 47122 1 39
2 47123 1 39
2 47124 1 39
2 47125 1 39
2 47126 1 39
2 47127 1 39
2 47128 1 39
2 47129 1 39
2 47130 1 39
2 47131 1 39
2 47132 1 39
2 47133 1 39
2 47134 1 39
2 47135 1 39
2 47136 1 39
2 47137 1 39
2 47138 1 39
2 47139 1 39
2 47140 1 39
2 47141 1 39
2 47142 1 39
2 47143 1 39
2 47144 1 39
2 47145 1 39
2 47146 1 39
2 47147 1 39
2 47148 1 39
2 47149 1 39
2 47150 1 39
2 47151 1 39
2 47152 1 39
2 47153 1 39
2 47154 1 39
2 47155 1 39
2 47156 1 39
2 47157 1 39
2 47158 1 40
2 47159 1 40
2 47160 1 40
2 47161 1 40
2 47162 1 40
2 47163 1 40
2 47164 1 40
2 47165 1 40
2 47166 1 40
2 47167 1 40
2 47168 1 40
2 47169 1 40
2 47170 1 40
2 47171 1 40
2 47172 1 40
2 47173 1 40
2 47174 1 40
2 47175 1 40
2 47176 1 40
2 47177 1 40
2 47178 1 40
2 47179 1 40
2 47180 1 40
2 47181 1 40
2 47182 1 40
2 47183 1 40
2 47184 1 40
2 47185 1 40
2 47186 1 40
2 47187 1 40
2 47188 1 40
2 47189 1 40
2 47190 1 40
2 47191 1 40
2 47192 1 40
2 47193 1 40
2 47194 1 40
2 47195 1 40
2 47196 1 40
2 47197 1 40
2 47198 1 40
2 47199 1 40
2 47200 1 40
2 47201 1 40
2 47202 1 40
2 47203 1 40
2 47204 1 40
2 47205 1 40
2 47206 1 40
2 47207 1 40
2 47208 1 40
2 47209 1 40
2 47210 1 40
2 47211 1 40
2 47212 1 40
2 47213 1 40
2 47214 1 40
2 47215 1 40
2 47216 1 40
2 47217 1 40
2 47218 1 40
2 47219 1 40
2 47220 1 40
2 47221 1 40
2 47222 1 40
2 47223 1 40
2 47224 1 40
2 47225 1 40
2 47226 1 40
2 47227 1 40
2 47228 1 40
2 47229 1 40
2 47230 1 40
2 47231 1 40
2 47232 1 40
2 47233 1 40
2 47234 1 40
2 47235 1 40
2 47236 1 40
2 47237 1 40
2 47238 1 40
2 47239 1 40
2 47240 1 40
2 47241 1 40
2 47242 1 40
2 47243 1 40
2 47244 1 40
2 47245 1 40
2 47246 1 40
2 47247 1 40
2 47248 1 40
2 47249 1 40
2 47250 1 40
2 47251 1 40
2 47252 1 40
2 47253 1 40
2 47254 1 40
2 47255 1 40
2 47256 1 40
2 47257 1 40
2 47258 1 40
2 47259 1 40
2 47260 1 40
2 47261 1 40
2 47262 1 40
2 47263 1 40
2 47264 1 40
2 47265 1 40
2 47266 1 40
2 47267 1 40
2 47268 1 40
2 47269 1 40
2 47270 1 40
2 47271 1 40
2 47272 1 40
2 47273 1 40
2 47274 1 40
2 47275 1 40
2 47276 1 40
2 47277 1 40
2 47278 1 40
2 47279 1 40
2 47280 1 40
2 47281 1 40
2 47282 1 40
2 47283 1 40
2 47284 1 40
2 47285 1 40
2 47286 1 40
2 47287 1 40
2 47288 1 40
2 47289 1 40
2 47290 1 40
2 47291 1 40
2 47292 1 40
2 47293 1 40
2 47294 1 40
2 47295 1 40
2 47296 1 40
2 47297 1 40
2 47298 1 40
2 47299 1 40
2 47300 1 40
2 47301 1 40
2 47302 1 40
2 47303 1 40
2 47304 1 40
2 47305 1 40
2 47306 1 40
2 47307 1 40
2 47308 1 40
2 47309 1 40
2 47310 1 40
2 47311 1 40
2 47312 1 40
2 47313 1 40
2 47314 1 40
2 47315 1 40
2 47316 1 40
2 47317 1 40
2 47318 1 40
2 47319 1 40
2 47320 1 40
2 47321 1 40
2 47322 1 40
2 47323 1 40
2 47324 1 40
2 47325 1 40
2 47326 1 40
2 47327 1 40
2 47328 1 40
2 47329 1 40
2 47330 1 41
2 47331 1 41
2 47332 1 41
2 47333 1 41
2 47334 1 41
2 47335 1 41
2 47336 1 41
2 47337 1 41
2 47338 1 41
2 47339 1 41
2 47340 1 41
2 47341 1 41
2 47342 1 41
2 47343 1 41
2 47344 1 41
2 47345 1 41
2 47346 1 41
2 47347 1 41
2 47348 1 41
2 47349 1 41
2 47350 1 41
2 47351 1 41
2 47352 1 41
2 47353 1 41
2 47354 1 41
2 47355 1 41
2 47356 1 41
2 47357 1 41
2 47358 1 41
2 47359 1 41
2 47360 1 41
2 47361 1 41
2 47362 1 41
2 47363 1 41
2 47364 1 41
2 47365 1 41
2 47366 1 41
2 47367 1 41
2 47368 1 41
2 47369 1 41
2 47370 1 41
2 47371 1 41
2 47372 1 41
2 47373 1 41
2 47374 1 41
2 47375 1 41
2 47376 1 41
2 47377 1 41
2 47378 1 41
2 47379 1 41
2 47380 1 41
2 47381 1 41
2 47382 1 41
2 47383 1 41
2 47384 1 41
2 47385 1 41
2 47386 1 41
2 47387 1 41
2 47388 1 41
2 47389 1 41
2 47390 1 41
2 47391 1 41
2 47392 1 41
2 47393 1 41
2 47394 1 41
2 47395 1 41
2 47396 1 41
2 47397 1 41
2 47398 1 41
2 47399 1 41
2 47400 1 41
2 47401 1 41
2 47402 1 41
2 47403 1 41
2 47404 1 41
2 47405 1 41
2 47406 1 41
2 47407 1 41
2 47408 1 41
2 47409 1 41
2 47410 1 41
2 47411 1 41
2 47412 1 41
2 47413 1 41
2 47414 1 41
2 47415 1 41
2 47416 1 41
2 47417 1 41
2 47418 1 41
2 47419 1 41
2 47420 1 41
2 47421 1 41
2 47422 1 41
2 47423 1 41
2 47424 1 41
2 47425 1 41
2 47426 1 41
2 47427 1 41
2 47428 1 41
2 47429 1 41
2 47430 1 41
2 47431 1 41
2 47432 1 41
2 47433 1 41
2 47434 1 41
2 47435 1 41
2 47436 1 41
2 47437 1 41
2 47438 1 41
2 47439 1 41
2 47440 1 41
2 47441 1 41
2 47442 1 41
2 47443 1 41
2 47444 1 41
2 47445 1 41
2 47446 1 41
2 47447 1 41
2 47448 1 41
2 47449 1 41
2 47450 1 41
2 47451 1 41
2 47452 1 41
2 47453 1 41
2 47454 1 41
2 47455 1 41
2 47456 1 41
2 47457 1 41
2 47458 1 41
2 47459 1 41
2 47460 1 41
2 47461 1 41
2 47462 1 41
2 47463 1 41
2 47464 1 41
2 47465 1 41
2 47466 1 41
2 47467 1 41
2 47468 1 41
2 47469 1 41
2 47470 1 41
2 47471 1 41
2 47472 1 41
2 47473 1 41
2 47474 1 41
2 47475 1 41
2 47476 1 42
2 47477 1 42
2 47478 1 42
2 47479 1 42
2 47480 1 42
2 47481 1 42
2 47482 1 42
2 47483 1 42
2 47484 1 42
2 47485 1 42
2 47486 1 42
2 47487 1 42
2 47488 1 42
2 47489 1 42
2 47490 1 42
2 47491 1 42
2 47492 1 42
2 47493 1 42
2 47494 1 42
2 47495 1 42
2 47496 1 42
2 47497 1 42
2 47498 1 42
2 47499 1 42
2 47500 1 42
2 47501 1 42
2 47502 1 42
2 47503 1 42
2 47504 1 42
2 47505 1 42
2 47506 1 42
2 47507 1 42
2 47508 1 42
2 47509 1 42
2 47510 1 42
2 47511 1 42
2 47512 1 42
2 47513 1 42
2 47514 1 42
2 47515 1 42
2 47516 1 42
2 47517 1 42
2 47518 1 42
2 47519 1 42
2 47520 1 42
2 47521 1 42
2 47522 1 42
2 47523 1 42
2 47524 1 42
2 47525 1 42
2 47526 1 42
2 47527 1 42
2 47528 1 42
2 47529 1 42
2 47530 1 42
2 47531 1 42
2 47532 1 42
2 47533 1 42
2 47534 1 42
2 47535 1 42
2 47536 1 42
2 47537 1 42
2 47538 1 42
2 47539 1 42
2 47540 1 42
2 47541 1 42
2 47542 1 42
2 47543 1 42
2 47544 1 42
2 47545 1 42
2 47546 1 42
2 47547 1 42
2 47548 1 42
2 47549 1 42
2 47550 1 42
2 47551 1 42
2 47552 1 42
2 47553 1 42
2 47554 1 42
2 47555 1 42
2 47556 1 42
2 47557 1 42
2 47558 1 42
2 47559 1 42
2 47560 1 42
2 47561 1 42
2 47562 1 42
2 47563 1 42
2 47564 1 42
2 47565 1 42
2 47566 1 42
2 47567 1 42
2 47568 1 42
2 47569 1 42
2 47570 1 42
2 47571 1 42
2 47572 1 42
2 47573 1 42
2 47574 1 42
2 47575 1 42
2 47576 1 42
2 47577 1 42
2 47578 1 42
2 47579 1 42
2 47580 1 42
2 47581 1 42
2 47582 1 42
2 47583 1 42
2 47584 1 42
2 47585 1 42
2 47586 1 42
2 47587 1 42
2 47588 1 42
2 47589 1 42
2 47590 1 42
2 47591 1 42
2 47592 1 42
2 47593 1 42
2 47594 1 42
2 47595 1 43
2 47596 1 43
2 47597 1 43
2 47598 1 43
2 47599 1 43
2 47600 1 43
2 47601 1 43
2 47602 1 43
2 47603 1 43
2 47604 1 43
2 47605 1 43
2 47606 1 43
2 47607 1 43
2 47608 1 43
2 47609 1 43
2 47610 1 43
2 47611 1 43
2 47612 1 43
2 47613 1 43
2 47614 1 43
2 47615 1 43
2 47616 1 43
2 47617 1 43
2 47618 1 43
2 47619 1 43
2 47620 1 43
2 47621 1 43
2 47622 1 43
2 47623 1 43
2 47624 1 43
2 47625 1 43
2 47626 1 43
2 47627 1 43
2 47628 1 43
2 47629 1 43
2 47630 1 43
2 47631 1 43
2 47632 1 43
2 47633 1 43
2 47634 1 43
2 47635 1 43
2 47636 1 43
2 47637 1 43
2 47638 1 43
2 47639 1 43
2 47640 1 43
2 47641 1 43
2 47642 1 43
2 47643 1 43
2 47644 1 43
2 47645 1 43
2 47646 1 43
2 47647 1 43
2 47648 1 43
2 47649 1 43
2 47650 1 43
2 47651 1 43
2 47652 1 43
2 47653 1 43
2 47654 1 43
2 47655 1 43
2 47656 1 43
2 47657 1 43
2 47658 1 43
2 47659 1 43
2 47660 1 43
2 47661 1 43
2 47662 1 43
2 47663 1 43
2 47664 1 43
2 47665 1 43
2 47666 1 43
2 47667 1 43
2 47668 1 43
2 47669 1 43
2 47670 1 43
2 47671 1 43
2 47672 1 43
2 47673 1 43
2 47674 1 43
2 47675 1 43
2 47676 1 43
2 47677 1 43
2 47678 1 43
2 47679 1 43
2 47680 1 43
2 47681 1 43
2 47682 1 43
2 47683 1 43
2 47684 1 43
2 47685 1 43
2 47686 1 43
2 47687 1 43
2 47688 1 43
2 47689 1 43
2 47690 1 43
2 47691 1 43
2 47692 1 43
2 47693 1 43
2 47694 1 43
2 47695 1 43
2 47696 1 43
2 47697 1 43
2 47698 1 43
2 47699 1 43
2 47700 1 43
2 47701 1 43
2 47702 1 44
2 47703 1 44
2 47704 1 44
2 47705 1 44
2 47706 1 44
2 47707 1 44
2 47708 1 44
2 47709 1 44
2 47710 1 44
2 47711 1 44
2 47712 1 44
2 47713 1 44
2 47714 1 44
2 47715 1 44
2 47716 1 44
2 47717 1 44
2 47718 1 44
2 47719 1 44
2 47720 1 44
2 47721 1 44
2 47722 1 44
2 47723 1 44
2 47724 1 44
2 47725 1 44
2 47726 1 44
2 47727 1 44
2 47728 1 44
2 47729 1 44
2 47730 1 44
2 47731 1 44
2 47732 1 44
2 47733 1 44
2 47734 1 44
2 47735 1 44
2 47736 1 44
2 47737 1 44
2 47738 1 44
2 47739 1 44
2 47740 1 44
2 47741 1 44
2 47742 1 44
2 47743 1 44
2 47744 1 44
2 47745 1 44
2 47746 1 44
2 47747 1 44
2 47748 1 44
2 47749 1 44
2 47750 1 44
2 47751 1 44
2 47752 1 44
2 47753 1 44
2 47754 1 44
2 47755 1 44
2 47756 1 44
2 47757 1 44
2 47758 1 44
2 47759 1 44
2 47760 1 44
2 47761 1 44
2 47762 1 44
2 47763 1 44
2 47764 1 44
2 47765 1 44
2 47766 1 44
2 47767 1 44
2 47768 1 44
2 47769 1 44
2 47770 1 44
2 47771 1 44
2 47772 1 44
2 47773 1 44
2 47774 1 44
2 47775 1 44
2 47776 1 44
2 47777 1 44
2 47778 1 44
2 47779 1 44
2 47780 1 44
2 47781 1 44
2 47782 1 44
2 47783 1 44
2 47784 1 44
2 47785 1 44
2 47786 1 44
2 47787 1 44
2 47788 1 44
2 47789 1 44
2 47790 1 44
2 47791 1 44
2 47792 1 44
2 47793 1 44
2 47794 1 44
2 47795 1 44
2 47796 1 44
2 47797 1 44
2 47798 1 44
2 47799 1 44
2 47800 1 44
2 47801 1 44
2 47802 1 44
2 47803 1 44
2 47804 1 44
2 47805 1 44
2 47806 1 44
2 47807 1 44
2 47808 1 44
2 47809 1 44
2 47810 1 44
2 47811 1 44
2 47812 1 44
2 47813 1 44
2 47814 1 44
2 47815 1 44
2 47816 1 44
2 47817 1 44
2 47818 1 44
2 47819 1 44
2 47820 1 44
2 47821 1 44
2 47822 1 44
2 47823 1 44
2 47824 1 44
2 47825 1 44
2 47826 1 44
2 47827 1 44
2 47828 1 44
2 47829 1 44
2 47830 1 44
2 47831 1 45
2 47832 1 45
2 47833 1 45
2 47834 1 45
2 47835 1 45
2 47836 1 45
2 47837 1 45
2 47838 1 45
2 47839 1 45
2 47840 1 45
2 47841 1 45
2 47842 1 45
2 47843 1 45
2 47844 1 45
2 47845 1 45
2 47846 1 45
2 47847 1 45
2 47848 1 45
2 47849 1 45
2 47850 1 45
2 47851 1 45
2 47852 1 45
2 47853 1 45
2 47854 1 45
2 47855 1 45
2 47856 1 45
2 47857 1 45
2 47858 1 45
2 47859 1 45
2 47860 1 45
2 47861 1 45
2 47862 1 45
2 47863 1 45
2 47864 1 45
2 47865 1 45
2 47866 1 45
2 47867 1 45
2 47868 1 45
2 47869 1 45
2 47870 1 45
2 47871 1 45
2 47872 1 45
2 47873 1 45
2 47874 1 45
2 47875 1 45
2 47876 1 45
2 47877 1 45
2 47878 1 45
2 47879 1 45
2 47880 1 45
2 47881 1 45
2 47882 1 45
2 47883 1 45
2 47884 1 45
2 47885 1 45
2 47886 1 45
2 47887 1 45
2 47888 1 45
2 47889 1 45
2 47890 1 45
2 47891 1 45
2 47892 1 45
2 47893 1 45
2 47894 1 45
2 47895 1 45
2 47896 1 45
2 47897 1 45
2 47898 1 45
2 47899 1 45
2 47900 1 45
2 47901 1 45
2 47902 1 45
2 47903 1 45
2 47904 1 45
2 47905 1 45
2 47906 1 45
2 47907 1 45
2 47908 1 45
2 47909 1 45
2 47910 1 45
2 47911 1 45
2 47912 1 45
2 47913 1 45
2 47914 1 45
2 47915 1 45
2 47916 1 45
2 47917 1 45
2 47918 1 45
2 47919 1 45
2 47920 1 45
2 47921 1 45
2 47922 1 45
2 47923 1 45
2 47924 1 45
2 47925 1 45
2 47926 1 45
2 47927 1 45
2 47928 1 45
2 47929 1 46
2 47930 1 46
2 47931 1 46
2 47932 1 46
2 47933 1 46
2 47934 1 46
2 47935 1 46
2 47936 1 46
2 47937 1 46
2 47938 1 46
2 47939 1 46
2 47940 1 46
2 47941 1 46
2 47942 1 46
2 47943 1 46
2 47944 1 46
2 47945 1 46
2 47946 1 46
2 47947 1 46
2 47948 1 46
2 47949 1 46
2 47950 1 46
2 47951 1 46
2 47952 1 46
2 47953 1 46
2 47954 1 46
2 47955 1 46
2 47956 1 46
2 47957 1 46
2 47958 1 46
2 47959 1 46
2 47960 1 46
2 47961 1 46
2 47962 1 46
2 47963 1 46
2 47964 1 46
2 47965 1 46
2 47966 1 46
2 47967 1 46
2 47968 1 46
2 47969 1 46
2 47970 1 46
2 47971 1 46
2 47972 1 46
2 47973 1 46
2 47974 1 46
2 47975 1 46
2 47976 1 46
2 47977 1 46
2 47978 1 46
2 47979 1 46
2 47980 1 46
2 47981 1 46
2 47982 1 46
2 47983 1 46
2 47984 1 46
2 47985 1 46
2 47986 1 46
2 47987 1 46
2 47988 1 46
2 47989 1 46
2 47990 1 46
2 47991 1 46
2 47992 1 46
2 47993 1 46
2 47994 1 46
2 47995 1 46
2 47996 1 46
2 47997 1 46
2 47998 1 46
2 47999 1 46
2 48000 1 46
2 48001 1 46
2 48002 1 46
2 48003 1 46
2 48004 1 46
2 48005 1 46
2 48006 1 46
2 48007 1 46
2 48008 1 46
2 48009 1 46
2 48010 1 46
2 48011 1 46
2 48012 1 46
2 48013 1 46
2 48014 1 46
2 48015 1 46
2 48016 1 46
2 48017 1 46
2 48018 1 46
2 48019 1 46
2 48020 1 46
2 48021 1 46
2 48022 1 46
2 48023 1 46
2 48024 1 46
2 48025 1 46
2 48026 1 46
2 48027 1 46
2 48028 1 46
2 48029 1 46
2 48030 1 46
2 48031 1 46
2 48032 1 46
2 48033 1 46
2 48034 1 46
2 48035 1 46
2 48036 1 46
2 48037 1 46
2 48038 1 46
2 48039 1 46
2 48040 1 46
2 48041 1 47
2 48042 1 47
2 48043 1 47
2 48044 1 47
2 48045 1 47
2 48046 1 47
2 48047 1 47
2 48048 1 47
2 48049 1 47
2 48050 1 47
2 48051 1 47
2 48052 1 47
2 48053 1 47
2 48054 1 47
2 48055 1 47
2 48056 1 47
2 48057 1 47
2 48058 1 47
2 48059 1 47
2 48060 1 47
2 48061 1 47
2 48062 1 47
2 48063 1 47
2 48064 1 47
2 48065 1 47
2 48066 1 47
2 48067 1 47
2 48068 1 47
2 48069 1 47
2 48070 1 47
2 48071 1 47
2 48072 1 47
2 48073 1 47
2 48074 1 47
2 48075 1 47
2 48076 1 47
2 48077 1 47
2 48078 1 47
2 48079 1 47
2 48080 1 47
2 48081 1 47
2 48082 1 47
2 48083 1 47
2 48084 1 47
2 48085 1 47
2 48086 1 47
2 48087 1 47
2 48088 1 47
2 48089 1 47
2 48090 1 47
2 48091 1 47
2 48092 1 47
2 48093 1 47
2 48094 1 47
2 48095 1 47
2 48096 1 47
2 48097 1 47
2 48098 1 47
2 48099 1 47
2 48100 1 47
2 48101 1 47
2 48102 1 47
2 48103 1 47
2 48104 1 47
2 48105 1 47
2 48106 1 47
2 48107 1 47
2 48108 1 47
2 48109 1 47
2 48110 1 47
2 48111 1 47
2 48112 1 47
2 48113 1 47
2 48114 1 47
2 48115 1 47
2 48116 1 47
2 48117 1 47
2 48118 1 47
2 48119 1 47
2 48120 1 47
2 48121 1 47
2 48122 1 47
2 48123 1 47
2 48124 1 47
2 48125 1 47
2 48126 1 47
2 48127 1 47
2 48128 1 47
2 48129 1 47
2 48130 1 47
2 48131 1 47
2 48132 1 47
2 48133 1 47
2 48134 1 47
2 48135 1 47
2 48136 1 47
2 48137 1 47
2 48138 1 47
2 48139 1 47
2 48140 1 47
2 48141 1 47
2 48142 1 47
2 48143 1 47
2 48144 1 47
2 48145 1 47
2 48146 1 47
2 48147 1 47
2 48148 1 47
2 48149 1 47
2 48150 1 47
2 48151 1 47
2 48152 1 47
2 48153 1 47
2 48154 1 47
2 48155 1 47
2 48156 1 47
2 48157 1 47
2 48158 1 47
2 48159 1 47
2 48160 1 47
2 48161 1 47
2 48162 1 47
2 48163 1 47
2 48164 1 47
2 48165 1 47
2 48166 1 47
2 48167 1 47
2 48168 1 48
2 48169 1 48
2 48170 1 48
2 48171 1 48
2 48172 1 48
2 48173 1 48
2 48174 1 48
2 48175 1 48
2 48176 1 48
2 48177 1 48
2 48178 1 48
2 48179 1 48
2 48180 1 48
2 48181 1 48
2 48182 1 48
2 48183 1 48
2 48184 1 48
2 48185 1 48
2 48186 1 48
2 48187 1 48
2 48188 1 48
2 48189 1 48
2 48190 1 48
2 48191 1 48
2 48192 1 48
2 48193 1 48
2 48194 1 48
2 48195 1 48
2 48196 1 48
2 48197 1 48
2 48198 1 48
2 48199 1 48
2 48200 1 48
2 48201 1 48
2 48202 1 48
2 48203 1 48
2 48204 1 48
2 48205 1 48
2 48206 1 48
2 48207 1 48
2 48208 1 48
2 48209 1 48
2 48210 1 48
2 48211 1 48
2 48212 1 48
2 48213 1 48
2 48214 1 48
2 48215 1 48
2 48216 1 48
2 48217 1 48
2 48218 1 48
2 48219 1 48
2 48220 1 48
2 48221 1 48
2 48222 1 48
2 48223 1 48
2 48224 1 48
2 48225 1 48
2 48226 1 48
2 48227 1 48
2 48228 1 48
2 48229 1 48
2 48230 1 48
2 48231 1 48
2 48232 1 48
2 48233 1 48
2 48234 1 48
2 48235 1 48
2 48236 1 48
2 48237 1 48
2 48238 1 48
2 48239 1 48
2 48240 1 48
2 48241 1 48
2 48242 1 48
2 48243 1 48
2 48244 1 48
2 48245 1 48
2 48246 1 48
2 48247 1 48
2 48248 1 48
2 48249 1 48
2 48250 1 48
2 48251 1 48
2 48252 1 48
2 48253 1 48
2 48254 1 48
2 48255 1 48
2 48256 1 48
2 48257 1 48
2 48258 1 48
2 48259 1 48
2 48260 1 48
2 48261 1 48
2 48262 1 48
2 48263 1 48
2 48264 1 48
2 48265 1 48
2 48266 1 48
2 48267 1 48
2 48268 1 48
2 48269 1 48
2 48270 1 48
2 48271 1 48
2 48272 1 48
2 48273 1 48
2 48274 1 48
2 48275 1 48
2 48276 1 48
2 48277 1 48
2 48278 1 48
2 48279 1 48
2 48280 1 48
2 48281 1 48
2 48282 1 48
2 48283 1 48
2 48284 1 48
2 48285 1 48
2 48286 1 48
2 48287 1 48
2 48288 1 48
2 48289 1 48
2 48290 1 48
2 48291 1 48
2 48292 1 48
2 48293 1 48
2 48294 1 48
2 48295 1 48
2 48296 1 48
2 48297 1 48
2 48298 1 48
2 48299 1 48
2 48300 1 48
2 48301 1 48
2 48302 1 48
2 48303 1 48
2 48304 1 48
2 48305 1 48
2 48306 1 48
2 48307 1 48
2 48308 1 48
2 48309 1 48
2 48310 1 48
2 48311 1 48
2 48312 1 48
2 48313 1 48
2 48314 1 48
2 48315 1 48
2 48316 1 48
2 48317 1 48
2 48318 1 48
2 48319 1 48
2 48320 1 48
2 48321 1 48
2 48322 1 48
2 48323 1 48
2 48324 1 48
2 48325 1 48
2 48326 1 48
2 48327 1 48
2 48328 1 48
2 48329 1 49
2 48330 1 49
2 48331 1 49
2 48332 1 49
2 48333 1 49
2 48334 1 49
2 48335 1 49
2 48336 1 49
2 48337 1 49
2 48338 1 49
2 48339 1 49
2 48340 1 49
2 48341 1 49
2 48342 1 49
2 48343 1 49
2 48344 1 49
2 48345 1 49
2 48346 1 49
2 48347 1 49
2 48348 1 49
2 48349 1 49
2 48350 1 49
2 48351 1 49
2 48352 1 49
2 48353 1 49
2 48354 1 49
2 48355 1 49
2 48356 1 49
2 48357 1 49
2 48358 1 49
2 48359 1 49
2 48360 1 49
2 48361 1 49
2 48362 1 49
2 48363 1 49
2 48364 1 49
2 48365 1 49
2 48366 1 49
2 48367 1 49
2 48368 1 49
2 48369 1 49
2 48370 1 49
2 48371 1 49
2 48372 1 49
2 48373 1 49
2 48374 1 49
2 48375 1 49
2 48376 1 49
2 48377 1 49
2 48378 1 49
2 48379 1 49
2 48380 1 49
2 48381 1 49
2 48382 1 49
2 48383 1 49
2 48384 1 49
2 48385 1 49
2 48386 1 49
2 48387 1 49
2 48388 1 49
2 48389 1 49
2 48390 1 49
2 48391 1 49
2 48392 1 49
2 48393 1 49
2 48394 1 49
2 48395 1 49
2 48396 1 49
2 48397 1 49
2 48398 1 49
2 48399 1 49
2 48400 1 49
2 48401 1 49
2 48402 1 49
2 48403 1 49
2 48404 1 49
2 48405 1 49
2 48406 1 49
2 48407 1 49
2 48408 1 49
2 48409 1 49
2 48410 1 49
2 48411 1 49
2 48412 1 49
2 48413 1 49
2 48414 1 49
2 48415 1 49
2 48416 1 49
2 48417 1 49
2 48418 1 49
2 48419 1 49
2 48420 1 49
2 48421 1 49
2 48422 1 49
2 48423 1 49
2 48424 1 49
2 48425 1 49
2 48426 1 49
2 48427 1 49
2 48428 1 49
2 48429 1 49
2 48430 1 49
2 48431 1 49
2 48432 1 49
2 48433 1 49
2 48434 1 49
2 48435 1 49
2 48436 1 49
2 48437 1 49
2 48438 1 49
2 48439 1 49
2 48440 1 49
2 48441 1 49
2 48442 1 49
2 48443 1 49
2 48444 1 49
2 48445 1 49
2 48446 1 49
2 48447 1 49
2 48448 1 49
2 48449 1 49
2 48450 1 49
2 48451 1 49
2 48452 1 49
2 48453 1 49
2 48454 1 49
2 48455 1 49
2 48456 1 49
2 48457 1 49
2 48458 1 49
2 48459 1 49
2 48460 1 49
2 48461 1 49
2 48462 1 49
2 48463 1 49
2 48464 1 49
2 48465 1 49
2 48466 1 49
2 48467 1 49
2 48468 1 49
2 48469 1 49
2 48470 1 49
2 48471 1 49
2 48472 1 49
2 48473 1 49
2 48474 1 49
2 48475 1 49
2 48476 1 49
2 48477 1 49
2 48478 1 49
2 48479 1 49
2 48480 1 49
2 48481 1 49
2 48482 1 49
2 48483 1 49
2 48484 1 49
2 48485 1 49
2 48486 1 49
2 48487 1 49
2 48488 1 49
2 48489 1 50
2 48490 1 50
2 48491 1 50
2 48492 1 50
2 48493 1 50
2 48494 1 50
2 48495 1 50
2 48496 1 50
2 48497 1 50
2 48498 1 50
2 48499 1 50
2 48500 1 50
2 48501 1 50
2 48502 1 50
2 48503 1 50
2 48504 1 50
2 48505 1 50
2 48506 1 50
2 48507 1 50
2 48508 1 50
2 48509 1 50
2 48510 1 50
2 48511 1 50
2 48512 1 50
2 48513 1 50
2 48514 1 50
2 48515 1 50
2 48516 1 50
2 48517 1 50
2 48518 1 50
2 48519 1 50
2 48520 1 50
2 48521 1 50
2 48522 1 50
2 48523 1 50
2 48524 1 50
2 48525 1 50
2 48526 1 50
2 48527 1 50
2 48528 1 50
2 48529 1 50
2 48530 1 50
2 48531 1 50
2 48532 1 50
2 48533 1 50
2 48534 1 50
2 48535 1 50
2 48536 1 50
2 48537 1 50
2 48538 1 50
2 48539 1 50
2 48540 1 50
2 48541 1 50
2 48542 1 50
2 48543 1 50
2 48544 1 50
2 48545 1 50
2 48546 1 50
2 48547 1 50
2 48548 1 50
2 48549 1 50
2 48550 1 50
2 48551 1 50
2 48552 1 50
2 48553 1 50
2 48554 1 50
2 48555 1 50
2 48556 1 50
2 48557 1 50
2 48558 1 50
2 48559 1 50
2 48560 1 50
2 48561 1 50
2 48562 1 50
2 48563 1 50
2 48564 1 50
2 48565 1 50
2 48566 1 50
2 48567 1 50
2 48568 1 50
2 48569 1 50
2 48570 1 50
2 48571 1 50
2 48572 1 50
2 48573 1 50
2 48574 1 50
2 48575 1 50
2 48576 1 50
2 48577 1 50
2 48578 1 50
2 48579 1 50
2 48580 1 50
2 48581 1 50
2 48582 1 50
2 48583 1 50
2 48584 1 50
2 48585 1 50
2 48586 1 50
2 48587 1 50
2 48588 1 50
2 48589 1 50
2 48590 1 50
2 48591 1 50
2 48592 1 50
2 48593 1 50
2 48594 1 50
2 48595 1 50
2 48596 1 50
2 48597 1 50
2 48598 1 50
2 48599 1 50
2 48600 1 50
2 48601 1 50
2 48602 1 50
2 48603 1 50
2 48604 1 50
2 48605 1 50
2 48606 1 50
2 48607 1 50
2 48608 1 50
2 48609 1 50
2 48610 1 50
2 48611 1 50
2 48612 1 50
2 48613 1 50
2 48614 1 50
2 48615 1 50
2 48616 1 50
2 48617 1 50
2 48618 1 50
2 48619 1 50
2 48620 1 50
2 48621 1 50
2 48622 1 50
2 48623 1 50
2 48624 1 50
2 48625 1 50
2 48626 1 50
2 48627 1 50
2 48628 1 50
2 48629 1 50
2 48630 1 50
2 48631 1 50
2 48632 1 50
2 48633 1 50
2 48634 1 50
2 48635 1 50
2 48636 1 50
2 48637 1 50
2 48638 1 50
2 48639 1 50
2 48640 1 50
2 48641 1 50
2 48642 1 50
2 48643 1 50
2 48644 1 50
2 48645 1 50
2 48646 1 50
2 48647 1 50
2 48648 1 50
2 48649 1 50
2 48650 1 50
2 48651 1 50
2 48652 1 50
2 48653 1 50
2 48654 1 50
2 48655 1 50
2 48656 1 50
2 48657 1 50
2 48658 1 50
2 48659 1 50
2 48660 1 50
2 48661 1 50
2 48662 1 50
2 48663 1 50
2 48664 1 50
2 48665 1 50
2 48666 1 50
2 48667 1 50
2 48668 1 50
2 48669 1 50
2 48670 1 50
2 48671 1 50
2 48672 1 50
2 48673 1 50
2 48674 1 50
2 48675 1 50
2 48676 1 50
2 48677 1 50
2 48678 1 50
2 48679 1 50
2 48680 1 50
2 48681 1 50
2 48682 1 50
2 48683 1 50
2 48684 1 50
2 48685 1 50
2 48686 1 50
2 48687 1 50
2 48688 1 50
2 48689 1 50
2 48690 1 50
2 48691 1 50
2 48692 1 50
2 48693 1 50
2 48694 1 50
2 48695 1 50
2 48696 1 50
2 48697 1 50
2 48698 1 50
2 48699 1 50
2 48700 1 50
2 48701 1 50
2 48702 1 50
2 48703 1 50
2 48704 1 50
2 48705 1 50
2 48706 1 50
2 48707 1 50
2 48708 1 50
2 48709 1 50
2 48710 1 50
2 48711 1 50
2 48712 1 50
2 48713 1 50
2 48714 1 50
2 48715 1 51
2 48716 1 51
2 48717 1 51
2 48718 1 51
2 48719 1 51
2 48720 1 51
2 48721 1 51
2 48722 1 51
2 48723 1 51
2 48724 1 51
2 48725 1 51
2 48726 1 51
2 48727 1 51
2 48728 1 51
2 48729 1 51
2 48730 1 51
2 48731 1 51
2 48732 1 51
2 48733 1 51
2 48734 1 51
2 48735 1 51
2 48736 1 51
2 48737 1 51
2 48738 1 51
2 48739 1 51
2 48740 1 51
2 48741 1 51
2 48742 1 51
2 48743 1 51
2 48744 1 51
2 48745 1 51
2 48746 1 51
2 48747 1 51
2 48748 1 51
2 48749 1 51
2 48750 1 51
2 48751 1 51
2 48752 1 51
2 48753 1 51
2 48754 1 51
2 48755 1 51
2 48756 1 51
2 48757 1 51
2 48758 1 51
2 48759 1 51
2 48760 1 51
2 48761 1 51
2 48762 1 51
2 48763 1 51
2 48764 1 51
2 48765 1 51
2 48766 1 51
2 48767 1 51
2 48768 1 51
2 48769 1 51
2 48770 1 51
2 48771 1 51
2 48772 1 51
2 48773 1 51
2 48774 1 51
2 48775 1 51
2 48776 1 51
2 48777 1 51
2 48778 1 51
2 48779 1 51
2 48780 1 51
2 48781 1 51
2 48782 1 51
2 48783 1 51
2 48784 1 51
2 48785 1 51
2 48786 1 51
2 48787 1 51
2 48788 1 51
2 48789 1 51
2 48790 1 51
2 48791 1 51
2 48792 1 51
2 48793 1 51
2 48794 1 51
2 48795 1 51
2 48796 1 51
2 48797 1 51
2 48798 1 51
2 48799 1 51
2 48800 1 51
2 48801 1 51
2 48802 1 51
2 48803 1 51
2 48804 1 51
2 48805 1 51
2 48806 1 51
2 48807 1 51
2 48808 1 51
2 48809 1 51
2 48810 1 51
2 48811 1 51
2 48812 1 51
2 48813 1 51
2 48814 1 51
2 48815 1 51
2 48816 1 51
2 48817 1 51
2 48818 1 51
2 48819 1 51
2 48820 1 51
2 48821 1 51
2 48822 1 51
2 48823 1 51
2 48824 1 51
2 48825 1 51
2 48826 1 51
2 48827 1 51
2 48828 1 51
2 48829 1 51
2 48830 1 51
2 48831 1 51
2 48832 1 51
2 48833 1 51
2 48834 1 51
2 48835 1 51
2 48836 1 51
2 48837 1 51
2 48838 1 51
2 48839 1 51
2 48840 1 51
2 48841 1 51
2 48842 1 51
2 48843 1 51
2 48844 1 51
2 48845 1 51
2 48846 1 51
2 48847 1 51
2 48848 1 51
2 48849 1 51
2 48850 1 51
2 48851 1 51
2 48852 1 51
2 48853 1 51
2 48854 1 51
2 48855 1 51
2 48856 1 51
2 48857 1 51
2 48858 1 51
2 48859 1 51
2 48860 1 51
2 48861 1 52
2 48862 1 52
2 48863 1 52
2 48864 1 52
2 48865 1 54
2 48866 1 54
2 48867 1 54
2 48868 1 55
2 48869 1 55
2 48870 1 56
2 48871 1 56
2 48872 1 57
2 48873 1 57
2 48874 1 57
2 48875 1 57
2 48876 1 57
2 48877 1 57
2 48878 1 57
2 48879 1 57
2 48880 1 57
2 48881 1 57
2 48882 1 57
2 48883 1 57
2 48884 1 58
2 48885 1 58
2 48886 1 58
2 48887 1 58
2 48888 1 58
2 48889 1 58
2 48890 1 58
2 48891 1 58
2 48892 1 58
2 48893 1 58
2 48894 1 58
2 48895 1 58
2 48896 1 58
2 48897 1 58
2 48898 1 58
2 48899 1 58
2 48900 1 58
2 48901 1 58
2 48902 1 58
2 48903 1 58
2 48904 1 58
2 48905 1 58
2 48906 1 58
2 48907 1 58
2 48908 1 58
2 48909 1 58
2 48910 1 58
2 48911 1 58
2 48912 1 58
2 48913 1 58
2 48914 1 58
2 48915 1 58
2 48916 1 59
2 48917 1 59
2 48918 1 59
2 48919 1 60
2 48920 1 60
2 48921 1 60
2 48922 1 60
2 48923 1 60
2 48924 1 60
2 48925 1 60
2 48926 1 61
2 48927 1 61
2 48928 1 61
2 48929 1 61
2 48930 1 61
2 48931 1 61
2 48932 1 61
2 48933 1 61
2 48934 1 61
2 48935 1 61
2 48936 1 61
2 48937 1 61
2 48938 1 61
2 48939 1 61
2 48940 1 61
2 48941 1 61
2 48942 1 61
2 48943 1 61
2 48944 1 61
2 48945 1 61
2 48946 1 61
2 48947 1 61
2 48948 1 61
2 48949 1 61
2 48950 1 61
2 48951 1 62
2 48952 1 62
2 48953 1 62
2 48954 1 62
2 48955 1 62
2 48956 1 62
2 48957 1 62
2 48958 1 62
2 48959 1 62
2 48960 1 62
2 48961 1 62
2 48962 1 62
2 48963 1 62
2 48964 1 62
2 48965 1 62
2 48966 1 62
2 48967 1 62
2 48968 1 62
2 48969 1 62
2 48970 1 62
2 48971 1 62
2 48972 1 62
2 48973 1 63
2 48974 1 63
2 48975 1 63
2 48976 1 63
2 48977 1 63
2 48978 1 63
2 48979 1 63
2 48980 1 63
2 48981 1 63
2 48982 1 64
2 48983 1 64
2 48984 1 64
2 48985 1 67
2 48986 1 67
2 48987 1 67
2 48988 1 67
2 48989 1 67
2 48990 1 67
2 48991 1 67
2 48992 1 67
2 48993 1 67
2 48994 1 67
2 48995 1 67
2 48996 1 67
2 48997 1 67
2 48998 1 67
2 48999 1 67
2 49000 1 67
2 49001 1 67
2 49002 1 67
2 49003 1 67
2 49004 1 67
2 49005 1 67
2 49006 1 67
2 49007 1 67
2 49008 1 67
2 49009 1 67
2 49010 1 67
2 49011 1 69
2 49012 1 69
2 49013 1 69
2 49014 1 69
2 49015 1 70
2 49016 1 70
2 49017 1 73
2 49018 1 73
2 49019 1 73
2 49020 1 73
2 49021 1 73
2 49022 1 73
2 49023 1 73
2 49024 1 73
2 49025 1 73
2 49026 1 73
2 49027 1 73
2 49028 1 73
2 49029 1 73
2 49030 1 73
2 49031 1 73
2 49032 1 73
2 49033 1 73
2 49034 1 73
2 49035 1 73
2 49036 1 73
2 49037 1 73
2 49038 1 73
2 49039 1 73
2 49040 1 73
2 49041 1 73
2 49042 1 73
2 49043 1 73
2 49044 1 73
2 49045 1 73
2 49046 1 73
2 49047 1 73
2 49048 1 73
2 49049 1 73
2 49050 1 73
2 49051 1 73
2 49052 1 73
2 49053 1 73
2 49054 1 73
2 49055 1 73
2 49056 1 73
2 49057 1 73
2 49058 1 73
2 49059 1 73
2 49060 1 73
2 49061 1 73
2 49062 1 74
2 49063 1 74
2 49064 1 74
2 49065 1 74
2 49066 1 74
2 49067 1 74
2 49068 1 74
2 49069 1 74
2 49070 1 74
2 49071 1 74
2 49072 1 74
2 49073 1 74
2 49074 1 74
2 49075 1 74
2 49076 1 74
2 49077 1 74
2 49078 1 74
2 49079 1 74
2 49080 1 74
2 49081 1 74
2 49082 1 74
2 49083 1 74
2 49084 1 74
2 49085 1 74
2 49086 1 74
2 49087 1 74
2 49088 1 74
2 49089 1 74
2 49090 1 74
2 49091 1 74
2 49092 1 74
2 49093 1 74
2 49094 1 74
2 49095 1 74
2 49096 1 74
2 49097 1 74
2 49098 1 74
2 49099 1 74
2 49100 1 74
2 49101 1 75
2 49102 1 75
2 49103 1 75
2 49104 1 75
2 49105 1 75
2 49106 1 76
2 49107 1 76
2 49108 1 76
2 49109 1 76
2 49110 1 76
2 49111 1 76
2 49112 1 76
2 49113 1 76
2 49114 1 78
2 49115 1 78
2 49116 1 86
2 49117 1 86
2 49118 1 86
2 49119 1 86
2 49120 1 86
2 49121 1 86
2 49122 1 86
2 49123 1 86
2 49124 1 86
2 49125 1 86
2 49126 1 87
2 49127 1 87
2 49128 1 88
2 49129 1 88
2 49130 1 88
2 49131 1 88
2 49132 1 88
2 49133 1 88
2 49134 1 88
2 49135 1 88
2 49136 1 88
2 49137 1 88
2 49138 1 88
2 49139 1 88
2 49140 1 88
2 49141 1 88
2 49142 1 88
2 49143 1 88
2 49144 1 88
2 49145 1 88
2 49146 1 88
2 49147 1 88
2 49148 1 88
2 49149 1 88
2 49150 1 88
2 49151 1 88
2 49152 1 88
2 49153 1 88
2 49154 1 88
2 49155 1 88
2 49156 1 88
2 49157 1 88
2 49158 1 88
2 49159 1 88
2 49160 1 88
2 49161 1 88
2 49162 1 88
2 49163 1 88
2 49164 1 88
2 49165 1 88
2 49166 1 88
2 49167 1 88
2 49168 1 88
2 49169 1 88
2 49170 1 88
2 49171 1 88
2 49172 1 88
2 49173 1 88
2 49174 1 88
2 49175 1 88
2 49176 1 88
2 49177 1 88
2 49178 1 88
2 49179 1 88
2 49180 1 88
2 49181 1 88
2 49182 1 88
2 49183 1 88
2 49184 1 89
2 49185 1 89
2 49186 1 89
2 49187 1 89
2 49188 1 89
2 49189 1 89
2 49190 1 89
2 49191 1 89
2 49192 1 89
2 49193 1 89
2 49194 1 89
2 49195 1 89
2 49196 1 89
2 49197 1 89
2 49198 1 89
2 49199 1 89
2 49200 1 89
2 49201 1 89
2 49202 1 89
2 49203 1 89
2 49204 1 89
2 49205 1 89
2 49206 1 89
2 49207 1 89
2 49208 1 89
2 49209 1 89
2 49210 1 89
2 49211 1 89
2 49212 1 89
2 49213 1 89
2 49214 1 89
2 49215 1 89
2 49216 1 89
2 49217 1 89
2 49218 1 89
2 49219 1 89
2 49220 1 89
2 49221 1 89
2 49222 1 89
2 49223 1 89
2 49224 1 89
2 49225 1 89
2 49226 1 89
2 49227 1 89
2 49228 1 89
2 49229 1 89
2 49230 1 89
2 49231 1 89
2 49232 1 89
2 49233 1 89
2 49234 1 89
2 49235 1 89
2 49236 1 89
2 49237 1 89
2 49238 1 89
2 49239 1 89
2 49240 1 89
2 49241 1 89
2 49242 1 89
2 49243 1 89
2 49244 1 90
2 49245 1 90
2 49246 1 91
2 49247 1 91
2 49248 1 91
2 49249 1 92
2 49250 1 92
2 49251 1 92
2 49252 1 93
2 49253 1 93
2 49254 1 95
2 49255 1 95
2 49256 1 100
2 49257 1 100
2 49258 1 100
2 49259 1 100
2 49260 1 100
2 49261 1 100
2 49262 1 100
2 49263 1 100
2 49264 1 100
2 49265 1 100
2 49266 1 100
2 49267 1 100
2 49268 1 100
2 49269 1 100
2 49270 1 100
2 49271 1 100
2 49272 1 100
2 49273 1 100
2 49274 1 100
2 49275 1 100
2 49276 1 100
2 49277 1 100
2 49278 1 100
2 49279 1 100
2 49280 1 100
2 49281 1 100
2 49282 1 100
2 49283 1 100
2 49284 1 100
2 49285 1 100
2 49286 1 100
2 49287 1 100
2 49288 1 100
2 49289 1 100
2 49290 1 100
2 49291 1 100
2 49292 1 100
2 49293 1 100
2 49294 1 100
2 49295 1 100
2 49296 1 100
2 49297 1 100
2 49298 1 100
2 49299 1 100
2 49300 1 100
2 49301 1 100
2 49302 1 100
2 49303 1 100
2 49304 1 100
2 49305 1 100
2 49306 1 100
2 49307 1 100
2 49308 1 100
2 49309 1 100
2 49310 1 100
2 49311 1 100
2 49312 1 100
2 49313 1 101
2 49314 1 101
2 49315 1 101
2 49316 1 101
2 49317 1 101
2 49318 1 101
2 49319 1 101
2 49320 1 101
2 49321 1 101
2 49322 1 101
2 49323 1 101
2 49324 1 101
2 49325 1 101
2 49326 1 101
2 49327 1 101
2 49328 1 101
2 49329 1 101
2 49330 1 101
2 49331 1 101
2 49332 1 101
2 49333 1 101
2 49334 1 101
2 49335 1 101
2 49336 1 101
2 49337 1 101
2 49338 1 101
2 49339 1 101
2 49340 1 101
2 49341 1 101
2 49342 1 101
2 49343 1 101
2 49344 1 101
2 49345 1 101
2 49346 1 101
2 49347 1 101
2 49348 1 101
2 49349 1 101
2 49350 1 101
2 49351 1 101
2 49352 1 101
2 49353 1 101
2 49354 1 101
2 49355 1 101
2 49356 1 101
2 49357 1 101
2 49358 1 101
2 49359 1 101
2 49360 1 101
2 49361 1 101
2 49362 1 101
2 49363 1 101
2 49364 1 101
2 49365 1 101
2 49366 1 101
2 49367 1 101
2 49368 1 101
2 49369 1 101
2 49370 1 101
2 49371 1 102
2 49372 1 102
2 49373 1 102
2 49374 1 102
2 49375 1 102
2 49376 1 102
2 49377 1 102
2 49378 1 102
2 49379 1 102
2 49380 1 102
2 49381 1 102
2 49382 1 102
2 49383 1 102
2 49384 1 102
2 49385 1 102
2 49386 1 102
2 49387 1 102
2 49388 1 102
2 49389 1 102
2 49390 1 102
2 49391 1 102
2 49392 1 102
2 49393 1 103
2 49394 1 103
2 49395 1 103
2 49396 1 104
2 49397 1 104
2 49398 1 104
2 49399 1 104
2 49400 1 104
2 49401 1 105
2 49402 1 105
2 49403 1 105
2 49404 1 105
2 49405 1 105
2 49406 1 105
2 49407 1 106
2 49408 1 106
2 49409 1 114
2 49410 1 114
2 49411 1 114
2 49412 1 115
2 49413 1 115
2 49414 1 116
2 49415 1 116
2 49416 1 116
2 49417 1 116
2 49418 1 116
2 49419 1 116
2 49420 1 116
2 49421 1 116
2 49422 1 116
2 49423 1 116
2 49424 1 116
2 49425 1 116
2 49426 1 116
2 49427 1 116
2 49428 1 118
2 49429 1 118
2 49430 1 118
2 49431 1 118
2 49432 1 124
2 49433 1 124
2 49434 1 124
2 49435 1 124
2 49436 1 124
2 49437 1 124
2 49438 1 124
2 49439 1 124
2 49440 1 124
2 49441 1 124
2 49442 1 124
2 49443 1 124
2 49444 1 124
2 49445 1 126
2 49446 1 126
2 49447 1 126
2 49448 1 126
2 49449 1 126
2 49450 1 126
2 49451 1 126
2 49452 1 126
2 49453 1 127
2 49454 1 127
2 49455 1 127
2 49456 1 127
2 49457 1 127
2 49458 1 128
2 49459 1 128
2 49460 1 130
2 49461 1 130
2 49462 1 130
2 49463 1 137
2 49464 1 137
2 49465 1 137
2 49466 1 137
2 49467 1 138
2 49468 1 138
2 49469 1 139
2 49470 1 139
2 49471 1 139
2 49472 1 139
2 49473 1 139
2 49474 1 139
2 49475 1 139
2 49476 1 140
2 49477 1 140
2 49478 1 141
2 49479 1 141
2 49480 1 141
2 49481 1 141
2 49482 1 141
2 49483 1 141
2 49484 1 141
2 49485 1 141
2 49486 1 141
2 49487 1 141
2 49488 1 141
2 49489 1 142
2 49490 1 142
2 49491 1 142
2 49492 1 144
2 49493 1 144
2 49494 1 147
2 49495 1 147
2 49496 1 147
2 49497 1 147
2 49498 1 147
2 49499 1 147
2 49500 1 147
2 49501 1 147
2 49502 1 150
2 49503 1 150
2 49504 1 150
2 49505 1 150
2 49506 1 150
2 49507 1 150
2 49508 1 150
2 49509 1 150
2 49510 1 150
2 49511 1 150
2 49512 1 150
2 49513 1 150
2 49514 1 150
2 49515 1 150
2 49516 1 150
2 49517 1 150
2 49518 1 150
2 49519 1 150
2 49520 1 150
2 49521 1 151
2 49522 1 151
2 49523 1 151
2 49524 1 151
2 49525 1 151
2 49526 1 151
2 49527 1 152
2 49528 1 152
2 49529 1 152
2 49530 1 152
2 49531 1 153
2 49532 1 153
2 49533 1 156
2 49534 1 156
2 49535 1 156
2 49536 1 156
2 49537 1 156
2 49538 1 156
2 49539 1 156
2 49540 1 156
2 49541 1 156
2 49542 1 156
2 49543 1 156
2 49544 1 156
2 49545 1 156
2 49546 1 157
2 49547 1 157
2 49548 1 157
2 49549 1 157
2 49550 1 157
2 49551 1 157
2 49552 1 157
2 49553 1 157
2 49554 1 157
2 49555 1 157
2 49556 1 166
2 49557 1 166
2 49558 1 166
2 49559 1 166
2 49560 1 166
2 49561 1 166
2 49562 1 166
2 49563 1 166
2 49564 1 166
2 49565 1 166
2 49566 1 166
2 49567 1 166
2 49568 1 166
2 49569 1 166
2 49570 1 166
2 49571 1 166
2 49572 1 166
2 49573 1 166
2 49574 1 166
2 49575 1 166
2 49576 1 166
2 49577 1 168
2 49578 1 168
2 49579 1 168
2 49580 1 169
2 49581 1 169
2 49582 1 169
2 49583 1 169
2 49584 1 169
2 49585 1 169
2 49586 1 169
2 49587 1 169
2 49588 1 178
2 49589 1 178
2 49590 1 178
2 49591 1 178
2 49592 1 178
2 49593 1 178
2 49594 1 179
2 49595 1 179
2 49596 1 179
2 49597 1 180
2 49598 1 180
2 49599 1 180
2 49600 1 180
2 49601 1 180
2 49602 1 180
2 49603 1 180
2 49604 1 184
2 49605 1 184
2 49606 1 184
2 49607 1 184
2 49608 1 184
2 49609 1 184
2 49610 1 184
2 49611 1 184
2 49612 1 184
2 49613 1 184
2 49614 1 184
2 49615 1 184
2 49616 1 184
2 49617 1 184
2 49618 1 184
2 49619 1 184
2 49620 1 184
2 49621 1 184
2 49622 1 184
2 49623 1 184
2 49624 1 184
2 49625 1 185
2 49626 1 185
2 49627 1 185
2 49628 1 185
2 49629 1 185
2 49630 1 185
2 49631 1 185
2 49632 1 185
2 49633 1 185
2 49634 1 187
2 49635 1 187
2 49636 1 187
2 49637 1 188
2 49638 1 188
2 49639 1 188
2 49640 1 188
2 49641 1 188
2 49642 1 188
2 49643 1 188
2 49644 1 188
2 49645 1 188
2 49646 1 188
2 49647 1 188
2 49648 1 188
2 49649 1 188
2 49650 1 188
2 49651 1 188
2 49652 1 188
2 49653 1 188
2 49654 1 188
2 49655 1 188
2 49656 1 188
2 49657 1 188
2 49658 1 188
2 49659 1 188
2 49660 1 188
2 49661 1 188
2 49662 1 188
2 49663 1 188
2 49664 1 189
2 49665 1 189
2 49666 1 190
2 49667 1 190
2 49668 1 190
2 49669 1 190
2 49670 1 190
2 49671 1 190
2 49672 1 190
2 49673 1 190
2 49674 1 190
2 49675 1 190
2 49676 1 190
2 49677 1 190
2 49678 1 190
2 49679 1 190
2 49680 1 190
2 49681 1 190
2 49682 1 190
2 49683 1 190
2 49684 1 190
2 49685 1 190
2 49686 1 190
2 49687 1 190
2 49688 1 190
2 49689 1 190
2 49690 1 190
2 49691 1 190
2 49692 1 190
2 49693 1 190
2 49694 1 190
2 49695 1 190
2 49696 1 190
2 49697 1 190
2 49698 1 190
2 49699 1 190
2 49700 1 190
2 49701 1 190
2 49702 1 190
2 49703 1 190
2 49704 1 190
2 49705 1 190
2 49706 1 190
2 49707 1 190
2 49708 1 190
2 49709 1 190
2 49710 1 190
2 49711 1 190
2 49712 1 190
2 49713 1 190
2 49714 1 190
2 49715 1 190
2 49716 1 190
2 49717 1 190
2 49718 1 190
2 49719 1 190
2 49720 1 191
2 49721 1 191
2 49722 1 191
2 49723 1 191
2 49724 1 191
2 49725 1 191
2 49726 1 191
2 49727 1 191
2 49728 1 191
2 49729 1 191
2 49730 1 191
2 49731 1 191
2 49732 1 191
2 49733 1 191
2 49734 1 191
2 49735 1 191
2 49736 1 191
2 49737 1 191
2 49738 1 191
2 49739 1 191
2 49740 1 191
2 49741 1 191
2 49742 1 191
2 49743 1 191
2 49744 1 191
2 49745 1 191
2 49746 1 191
2 49747 1 191
2 49748 1 191
2 49749 1 191
2 49750 1 191
2 49751 1 191
2 49752 1 191
2 49753 1 191
2 49754 1 191
2 49755 1 191
2 49756 1 191
2 49757 1 191
2 49758 1 191
2 49759 1 191
2 49760 1 191
2 49761 1 191
2 49762 1 191
2 49763 1 191
2 49764 1 191
2 49765 1 191
2 49766 1 191
2 49767 1 191
2 49768 1 191
2 49769 1 191
2 49770 1 191
2 49771 1 191
2 49772 1 191
2 49773 1 191
2 49774 1 192
2 49775 1 192
2 49776 1 192
2 49777 1 192
2 49778 1 192
2 49779 1 192
2 49780 1 192
2 49781 1 192
2 49782 1 192
2 49783 1 192
2 49784 1 193
2 49785 1 193
2 49786 1 193
2 49787 1 193
2 49788 1 193
2 49789 1 193
2 49790 1 193
2 49791 1 193
2 49792 1 201
2 49793 1 201
2 49794 1 201
2 49795 1 201
2 49796 1 201
2 49797 1 201
2 49798 1 201
2 49799 1 201
2 49800 1 201
2 49801 1 201
2 49802 1 204
2 49803 1 204
2 49804 1 204
2 49805 1 204
2 49806 1 204
2 49807 1 204
2 49808 1 204
2 49809 1 204
2 49810 1 204
2 49811 1 205
2 49812 1 205
2 49813 1 205
2 49814 1 205
2 49815 1 205
2 49816 1 205
2 49817 1 205
2 49818 1 205
2 49819 1 205
2 49820 1 205
2 49821 1 205
2 49822 1 205
2 49823 1 205
2 49824 1 205
2 49825 1 205
2 49826 1 205
2 49827 1 205
2 49828 1 205
2 49829 1 208
2 49830 1 208
2 49831 1 210
2 49832 1 210
2 49833 1 210
2 49834 1 210
2 49835 1 210
2 49836 1 210
2 49837 1 211
2 49838 1 211
2 49839 1 211
2 49840 1 211
2 49841 1 211
2 49842 1 211
2 49843 1 211
2 49844 1 211
2 49845 1 212
2 49846 1 212
2 49847 1 220
2 49848 1 220
2 49849 1 220
2 49850 1 220
2 49851 1 220
2 49852 1 220
2 49853 1 220
2 49854 1 220
2 49855 1 220
2 49856 1 220
2 49857 1 220
2 49858 1 220
2 49859 1 220
2 49860 1 220
2 49861 1 220
2 49862 1 220
2 49863 1 221
2 49864 1 221
2 49865 1 221
2 49866 1 221
2 49867 1 222
2 49868 1 222
2 49869 1 222
2 49870 1 222
2 49871 1 223
2 49872 1 223
2 49873 1 223
2 49874 1 223
2 49875 1 223
2 49876 1 223
2 49877 1 223
2 49878 1 223
2 49879 1 223
2 49880 1 223
2 49881 1 223
2 49882 1 223
2 49883 1 224
2 49884 1 224
2 49885 1 225
2 49886 1 225
2 49887 1 225
2 49888 1 225
2 49889 1 225
2 49890 1 227
2 49891 1 227
2 49892 1 227
2 49893 1 227
2 49894 1 227
2 49895 1 227
2 49896 1 227
2 49897 1 227
2 49898 1 227
2 49899 1 227
2 49900 1 228
2 49901 1 228
2 49902 1 228
2 49903 1 237
2 49904 1 237
2 49905 1 237
2 49906 1 237
2 49907 1 237
2 49908 1 237
2 49909 1 237
2 49910 1 237
2 49911 1 237
2 49912 1 237
2 49913 1 237
2 49914 1 237
2 49915 1 237
2 49916 1 237
2 49917 1 237
2 49918 1 237
2 49919 1 237
2 49920 1 237
2 49921 1 237
2 49922 1 237
2 49923 1 237
2 49924 1 238
2 49925 1 238
2 49926 1 239
2 49927 1 239
2 49928 1 242
2 49929 1 242
2 49930 1 242
2 49931 1 242
2 49932 1 242
2 49933 1 242
2 49934 1 242
2 49935 1 242
2 49936 1 242
2 49937 1 242
2 49938 1 242
2 49939 1 242
2 49940 1 242
2 49941 1 242
2 49942 1 242
2 49943 1 242
2 49944 1 242
2 49945 1 242
2 49946 1 242
2 49947 1 242
2 49948 1 242
2 49949 1 242
2 49950 1 242
2 49951 1 242
2 49952 1 242
2 49953 1 242
2 49954 1 242
2 49955 1 242
2 49956 1 242
2 49957 1 242
2 49958 1 242
2 49959 1 242
2 49960 1 242
2 49961 1 242
2 49962 1 242
2 49963 1 242
2 49964 1 242
2 49965 1 242
2 49966 1 242
2 49967 1 242
2 49968 1 242
2 49969 1 242
2 49970 1 242
2 49971 1 242
2 49972 1 242
2 49973 1 242
2 49974 1 242
2 49975 1 242
2 49976 1 242
2 49977 1 242
2 49978 1 242
2 49979 1 242
2 49980 1 242
2 49981 1 242
2 49982 1 242
2 49983 1 242
2 49984 1 242
2 49985 1 242
2 49986 1 242
2 49987 1 242
2 49988 1 242
2 49989 1 242
2 49990 1 242
2 49991 1 242
2 49992 1 242
2 49993 1 242
2 49994 1 242
2 49995 1 242
2 49996 1 242
2 49997 1 242
2 49998 1 242
2 49999 1 242
2 50000 1 242
2 50001 1 242
2 50002 1 242
2 50003 1 242
2 50004 1 242
2 50005 1 242
2 50006 1 242
2 50007 1 242
2 50008 1 242
2 50009 1 242
2 50010 1 242
2 50011 1 242
2 50012 1 242
2 50013 1 242
2 50014 1 242
2 50015 1 242
2 50016 1 242
2 50017 1 242
2 50018 1 242
2 50019 1 242
2 50020 1 242
2 50021 1 242
2 50022 1 242
2 50023 1 242
2 50024 1 242
2 50025 1 242
2 50026 1 242
2 50027 1 242
2 50028 1 242
2 50029 1 242
2 50030 1 242
2 50031 1 242
2 50032 1 242
2 50033 1 243
2 50034 1 243
2 50035 1 243
2 50036 1 243
2 50037 1 243
2 50038 1 243
2 50039 1 243
2 50040 1 243
2 50041 1 243
2 50042 1 243
2 50043 1 243
2 50044 1 243
2 50045 1 243
2 50046 1 243
2 50047 1 243
2 50048 1 243
2 50049 1 243
2 50050 1 243
2 50051 1 243
2 50052 1 243
2 50053 1 243
2 50054 1 243
2 50055 1 243
2 50056 1 243
2 50057 1 243
2 50058 1 243
2 50059 1 243
2 50060 1 243
2 50061 1 243
2 50062 1 243
2 50063 1 243
2 50064 1 243
2 50065 1 243
2 50066 1 243
2 50067 1 243
2 50068 1 243
2 50069 1 243
2 50070 1 243
2 50071 1 243
2 50072 1 243
2 50073 1 243
2 50074 1 243
2 50075 1 243
2 50076 1 243
2 50077 1 243
2 50078 1 243
2 50079 1 243
2 50080 1 243
2 50081 1 243
2 50082 1 243
2 50083 1 243
2 50084 1 243
2 50085 1 243
2 50086 1 243
2 50087 1 243
2 50088 1 243
2 50089 1 243
2 50090 1 243
2 50091 1 243
2 50092 1 243
2 50093 1 243
2 50094 1 243
2 50095 1 243
2 50096 1 243
2 50097 1 243
2 50098 1 243
2 50099 1 243
2 50100 1 243
2 50101 1 243
2 50102 1 243
2 50103 1 243
2 50104 1 243
2 50105 1 243
2 50106 1 243
2 50107 1 243
2 50108 1 243
2 50109 1 243
2 50110 1 243
2 50111 1 243
2 50112 1 243
2 50113 1 243
2 50114 1 243
2 50115 1 243
2 50116 1 243
2 50117 1 243
2 50118 1 243
2 50119 1 243
2 50120 1 243
2 50121 1 244
2 50122 1 244
2 50123 1 244
2 50124 1 245
2 50125 1 245
2 50126 1 245
2 50127 1 245
2 50128 1 245
2 50129 1 245
2 50130 1 245
2 50131 1 245
2 50132 1 245
2 50133 1 245
2 50134 1 245
2 50135 1 246
2 50136 1 246
2 50137 1 246
2 50138 1 254
2 50139 1 254
2 50140 1 254
2 50141 1 254
2 50142 1 254
2 50143 1 254
2 50144 1 255
2 50145 1 255
2 50146 1 255
2 50147 1 255
2 50148 1 256
2 50149 1 256
2 50150 1 256
2 50151 1 256
2 50152 1 256
2 50153 1 256
2 50154 1 256
2 50155 1 256
2 50156 1 256
2 50157 1 256
2 50158 1 256
2 50159 1 256
2 50160 1 256
2 50161 1 256
2 50162 1 256
2 50163 1 256
2 50164 1 256
2 50165 1 256
2 50166 1 256
2 50167 1 256
2 50168 1 256
2 50169 1 258
2 50170 1 258
2 50171 1 260
2 50172 1 260
2 50173 1 260
2 50174 1 260
2 50175 1 260
2 50176 1 260
2 50177 1 261
2 50178 1 261
2 50179 1 261
2 50180 1 261
2 50181 1 262
2 50182 1 262
2 50183 1 262
2 50184 1 262
2 50185 1 262
2 50186 1 262
2 50187 1 262
2 50188 1 263
2 50189 1 263
2 50190 1 263
2 50191 1 264
2 50192 1 264
2 50193 1 264
2 50194 1 264
2 50195 1 264
2 50196 1 264
2 50197 1 264
2 50198 1 265
2 50199 1 265
2 50200 1 275
2 50201 1 275
2 50202 1 275
2 50203 1 275
2 50204 1 275
2 50205 1 275
2 50206 1 275
2 50207 1 275
2 50208 1 275
2 50209 1 283
2 50210 1 283
2 50211 1 283
2 50212 1 283
2 50213 1 283
2 50214 1 283
2 50215 1 283
2 50216 1 284
2 50217 1 284
2 50218 1 284
2 50219 1 284
2 50220 1 284
2 50221 1 284
2 50222 1 284
2 50223 1 284
2 50224 1 284
2 50225 1 284
2 50226 1 284
2 50227 1 284
2 50228 1 284
2 50229 1 284
2 50230 1 284
2 50231 1 284
2 50232 1 284
2 50233 1 285
2 50234 1 285
2 50235 1 285
2 50236 1 286
2 50237 1 286
2 50238 1 286
2 50239 1 286
2 50240 1 286
2 50241 1 286
2 50242 1 287
2 50243 1 287
2 50244 1 287
2 50245 1 287
2 50246 1 288
2 50247 1 288
2 50248 1 288
2 50249 1 288
2 50250 1 288
2 50251 1 288
2 50252 1 288
2 50253 1 289
2 50254 1 289
2 50255 1 291
2 50256 1 291
2 50257 1 291
2 50258 1 291
2 50259 1 291
2 50260 1 291
2 50261 1 291
2 50262 1 291
2 50263 1 291
2 50264 1 292
2 50265 1 292
2 50266 1 292
2 50267 1 292
2 50268 1 292
2 50269 1 292
2 50270 1 292
2 50271 1 295
2 50272 1 295
2 50273 1 295
2 50274 1 295
2 50275 1 295
2 50276 1 295
2 50277 1 295
2 50278 1 295
2 50279 1 296
2 50280 1 296
2 50281 1 296
2 50282 1 296
2 50283 1 297
2 50284 1 297
2 50285 1 297
2 50286 1 297
2 50287 1 297
2 50288 1 297
2 50289 1 299
2 50290 1 299
2 50291 1 304
2 50292 1 304
2 50293 1 307
2 50294 1 307
2 50295 1 307
2 50296 1 307
2 50297 1 307
2 50298 1 308
2 50299 1 308
2 50300 1 309
2 50301 1 309
2 50302 1 310
2 50303 1 310
2 50304 1 310
2 50305 1 310
2 50306 1 310
2 50307 1 311
2 50308 1 311
2 50309 1 313
2 50310 1 313
2 50311 1 318
2 50312 1 318
2 50313 1 318
2 50314 1 329
2 50315 1 329
2 50316 1 329
2 50317 1 330
2 50318 1 330
2 50319 1 330
2 50320 1 330
2 50321 1 330
2 50322 1 330
2 50323 1 330
2 50324 1 331
2 50325 1 331
2 50326 1 334
2 50327 1 334
2 50328 1 334
2 50329 1 334
2 50330 1 334
2 50331 1 334
2 50332 1 334
2 50333 1 334
2 50334 1 334
2 50335 1 334
2 50336 1 334
2 50337 1 335
2 50338 1 335
2 50339 1 336
2 50340 1 336
2 50341 1 336
2 50342 1 337
2 50343 1 337
2 50344 1 349
2 50345 1 349
2 50346 1 349
2 50347 1 349
2 50348 1 349
2 50349 1 349
2 50350 1 349
2 50351 1 349
2 50352 1 349
2 50353 1 349
2 50354 1 349
2 50355 1 349
2 50356 1 349
2 50357 1 349
2 50358 1 349
2 50359 1 349
2 50360 1 349
2 50361 1 349
2 50362 1 349
2 50363 1 349
2 50364 1 349
2 50365 1 349
2 50366 1 349
2 50367 1 349
2 50368 1 349
2 50369 1 349
2 50370 1 349
2 50371 1 349
2 50372 1 349
2 50373 1 349
2 50374 1 350
2 50375 1 350
2 50376 1 350
2 50377 1 350
2 50378 1 350
2 50379 1 350
2 50380 1 350
2 50381 1 350
2 50382 1 350
2 50383 1 351
2 50384 1 351
2 50385 1 359
2 50386 1 359
2 50387 1 361
2 50388 1 361
2 50389 1 361
2 50390 1 366
2 50391 1 366
2 50392 1 366
2 50393 1 366
2 50394 1 366
2 50395 1 366
2 50396 1 366
2 50397 1 366
2 50398 1 366
2 50399 1 366
2 50400 1 366
2 50401 1 366
2 50402 1 366
2 50403 1 366
2 50404 1 366
2 50405 1 366
2 50406 1 366
2 50407 1 366
2 50408 1 366
2 50409 1 366
2 50410 1 366
2 50411 1 366
2 50412 1 366
2 50413 1 366
2 50414 1 366
2 50415 1 366
2 50416 1 366
2 50417 1 366
2 50418 1 366
2 50419 1 366
2 50420 1 366
2 50421 1 366
2 50422 1 366
2 50423 1 366
2 50424 1 366
2 50425 1 366
2 50426 1 366
2 50427 1 366
2 50428 1 366
2 50429 1 366
2 50430 1 366
2 50431 1 366
2 50432 1 366
2 50433 1 366
2 50434 1 366
2 50435 1 366
2 50436 1 366
2 50437 1 366
2 50438 1 366
2 50439 1 366
2 50440 1 366
2 50441 1 366
2 50442 1 366
2 50443 1 366
2 50444 1 366
2 50445 1 367
2 50446 1 367
2 50447 1 367
2 50448 1 367
2 50449 1 367
2 50450 1 367
2 50451 1 367
2 50452 1 367
2 50453 1 367
2 50454 1 367
2 50455 1 367
2 50456 1 367
2 50457 1 367
2 50458 1 367
2 50459 1 367
2 50460 1 367
2 50461 1 367
2 50462 1 367
2 50463 1 367
2 50464 1 367
2 50465 1 367
2 50466 1 367
2 50467 1 367
2 50468 1 367
2 50469 1 367
2 50470 1 367
2 50471 1 367
2 50472 1 367
2 50473 1 367
2 50474 1 367
2 50475 1 367
2 50476 1 367
2 50477 1 367
2 50478 1 367
2 50479 1 367
2 50480 1 367
2 50481 1 367
2 50482 1 368
2 50483 1 368
2 50484 1 368
2 50485 1 368
2 50486 1 369
2 50487 1 369
2 50488 1 369
2 50489 1 369
2 50490 1 369
2 50491 1 369
2 50492 1 369
2 50493 1 369
2 50494 1 369
2 50495 1 369
2 50496 1 369
2 50497 1 369
2 50498 1 369
2 50499 1 369
2 50500 1 369
2 50501 1 369
2 50502 1 369
2 50503 1 369
2 50504 1 369
2 50505 1 369
2 50506 1 369
2 50507 1 369
2 50508 1 369
2 50509 1 369
2 50510 1 369
2 50511 1 369
2 50512 1 371
2 50513 1 371
2 50514 1 371
2 50515 1 371
2 50516 1 371
2 50517 1 375
2 50518 1 375
2 50519 1 375
2 50520 1 375
2 50521 1 375
2 50522 1 375
2 50523 1 377
2 50524 1 377
2 50525 1 378
2 50526 1 378
2 50527 1 379
2 50528 1 379
2 50529 1 379
2 50530 1 379
2 50531 1 379
2 50532 1 379
2 50533 1 379
2 50534 1 379
2 50535 1 379
2 50536 1 379
2 50537 1 379
2 50538 1 379
2 50539 1 379
2 50540 1 379
2 50541 1 379
2 50542 1 379
2 50543 1 379
2 50544 1 379
2 50545 1 379
2 50546 1 379
2 50547 1 379
2 50548 1 379
2 50549 1 379
2 50550 1 379
2 50551 1 379
2 50552 1 379
2 50553 1 379
2 50554 1 379
2 50555 1 379
2 50556 1 379
2 50557 1 379
2 50558 1 379
2 50559 1 379
2 50560 1 379
2 50561 1 379
2 50562 1 379
2 50563 1 379
2 50564 1 379
2 50565 1 379
2 50566 1 379
2 50567 1 379
2 50568 1 379
2 50569 1 379
2 50570 1 379
2 50571 1 379
2 50572 1 379
2 50573 1 379
2 50574 1 379
2 50575 1 379
2 50576 1 379
2 50577 1 379
2 50578 1 379
2 50579 1 379
2 50580 1 379
2 50581 1 379
2 50582 1 379
2 50583 1 380
2 50584 1 380
2 50585 1 380
2 50586 1 380
2 50587 1 380
2 50588 1 380
2 50589 1 380
2 50590 1 380
2 50591 1 380
2 50592 1 380
2 50593 1 380
2 50594 1 380
2 50595 1 380
2 50596 1 380
2 50597 1 380
2 50598 1 380
2 50599 1 380
2 50600 1 380
2 50601 1 380
2 50602 1 380
2 50603 1 380
2 50604 1 380
2 50605 1 380
2 50606 1 380
2 50607 1 380
2 50608 1 380
2 50609 1 380
2 50610 1 380
2 50611 1 380
2 50612 1 380
2 50613 1 380
2 50614 1 380
2 50615 1 380
2 50616 1 380
2 50617 1 380
2 50618 1 380
2 50619 1 380
2 50620 1 380
2 50621 1 380
2 50622 1 380
2 50623 1 380
2 50624 1 380
2 50625 1 381
2 50626 1 381
2 50627 1 381
2 50628 1 381
2 50629 1 381
2 50630 1 381
2 50631 1 381
2 50632 1 381
2 50633 1 381
2 50634 1 382
2 50635 1 382
2 50636 1 382
2 50637 1 382
2 50638 1 382
2 50639 1 382
2 50640 1 386
2 50641 1 386
2 50642 1 387
2 50643 1 387
2 50644 1 387
2 50645 1 387
2 50646 1 387
2 50647 1 387
2 50648 1 387
2 50649 1 387
2 50650 1 387
2 50651 1 387
2 50652 1 387
2 50653 1 387
2 50654 1 387
2 50655 1 387
2 50656 1 387
2 50657 1 387
2 50658 1 387
2 50659 1 387
2 50660 1 387
2 50661 1 387
2 50662 1 387
2 50663 1 387
2 50664 1 387
2 50665 1 387
2 50666 1 387
2 50667 1 388
2 50668 1 388
2 50669 1 388
2 50670 1 388
2 50671 1 388
2 50672 1 388
2 50673 1 388
2 50674 1 388
2 50675 1 388
2 50676 1 389
2 50677 1 389
2 50678 1 389
2 50679 1 389
2 50680 1 390
2 50681 1 390
2 50682 1 390
2 50683 1 391
2 50684 1 391
2 50685 1 400
2 50686 1 400
2 50687 1 401
2 50688 1 401
2 50689 1 410
2 50690 1 410
2 50691 1 411
2 50692 1 411
2 50693 1 411
2 50694 1 415
2 50695 1 415
2 50696 1 415
2 50697 1 415
2 50698 1 415
2 50699 1 415
2 50700 1 415
2 50701 1 416
2 50702 1 416
2 50703 1 416
2 50704 1 423
2 50705 1 423
2 50706 1 423
2 50707 1 424
2 50708 1 424
2 50709 1 424
2 50710 1 432
2 50711 1 432
2 50712 1 433
2 50713 1 433
2 50714 1 433
2 50715 1 433
2 50716 1 433
2 50717 1 434
2 50718 1 434
2 50719 1 434
2 50720 1 434
2 50721 1 434
2 50722 1 434
2 50723 1 444
2 50724 1 444
2 50725 1 444
2 50726 1 444
2 50727 1 444
2 50728 1 444
2 50729 1 444
2 50730 1 444
2 50731 1 444
2 50732 1 444
2 50733 1 444
2 50734 1 444
2 50735 1 444
2 50736 1 444
2 50737 1 444
2 50738 1 444
2 50739 1 444
2 50740 1 444
2 50741 1 444
2 50742 1 444
2 50743 1 444
2 50744 1 444
2 50745 1 444
2 50746 1 444
2 50747 1 444
2 50748 1 444
2 50749 1 444
2 50750 1 444
2 50751 1 444
2 50752 1 444
2 50753 1 444
2 50754 1 444
2 50755 1 444
2 50756 1 444
2 50757 1 444
2 50758 1 444
2 50759 1 444
2 50760 1 444
2 50761 1 444
2 50762 1 444
2 50763 1 444
2 50764 1 444
2 50765 1 444
2 50766 1 444
2 50767 1 444
2 50768 1 444
2 50769 1 444
2 50770 1 444
2 50771 1 444
2 50772 1 444
2 50773 1 444
2 50774 1 444
2 50775 1 444
2 50776 1 444
2 50777 1 444
2 50778 1 444
2 50779 1 444
2 50780 1 444
2 50781 1 444
2 50782 1 444
2 50783 1 444
2 50784 1 444
2 50785 1 444
2 50786 1 444
2 50787 1 444
2 50788 1 444
2 50789 1 444
2 50790 1 444
2 50791 1 444
2 50792 1 444
2 50793 1 444
2 50794 1 444
2 50795 1 444
2 50796 1 444
2 50797 1 444
2 50798 1 444
2 50799 1 444
2 50800 1 444
2 50801 1 444
2 50802 1 444
2 50803 1 444
2 50804 1 444
2 50805 1 444
2 50806 1 444
2 50807 1 444
2 50808 1 444
2 50809 1 444
2 50810 1 445
2 50811 1 445
2 50812 1 445
2 50813 1 445
2 50814 1 445
2 50815 1 445
2 50816 1 445
2 50817 1 445
2 50818 1 445
2 50819 1 445
2 50820 1 445
2 50821 1 445
2 50822 1 445
2 50823 1 445
2 50824 1 445
2 50825 1 445
2 50826 1 445
2 50827 1 445
2 50828 1 445
2 50829 1 445
2 50830 1 445
2 50831 1 445
2 50832 1 445
2 50833 1 445
2 50834 1 445
2 50835 1 445
2 50836 1 445
2 50837 1 445
2 50838 1 445
2 50839 1 445
2 50840 1 445
2 50841 1 445
2 50842 1 445
2 50843 1 445
2 50844 1 445
2 50845 1 445
2 50846 1 445
2 50847 1 445
2 50848 1 445
2 50849 1 445
2 50850 1 445
2 50851 1 445
2 50852 1 445
2 50853 1 445
2 50854 1 445
2 50855 1 445
2 50856 1 445
2 50857 1 445
2 50858 1 445
2 50859 1 445
2 50860 1 445
2 50861 1 445
2 50862 1 445
2 50863 1 445
2 50864 1 445
2 50865 1 445
2 50866 1 445
2 50867 1 445
2 50868 1 445
2 50869 1 445
2 50870 1 445
2 50871 1 445
2 50872 1 445
2 50873 1 445
2 50874 1 445
2 50875 1 445
2 50876 1 445
2 50877 1 445
2 50878 1 445
2 50879 1 445
2 50880 1 445
2 50881 1 445
2 50882 1 445
2 50883 1 445
2 50884 1 445
2 50885 1 445
2 50886 1 445
2 50887 1 445
2 50888 1 446
2 50889 1 446
2 50890 1 446
2 50891 1 447
2 50892 1 447
2 50893 1 447
2 50894 1 447
2 50895 1 447
2 50896 1 449
2 50897 1 449
2 50898 1 449
2 50899 1 449
2 50900 1 449
2 50901 1 452
2 50902 1 452
2 50903 1 452
2 50904 1 452
2 50905 1 452
2 50906 1 452
2 50907 1 452
2 50908 1 452
2 50909 1 453
2 50910 1 453
2 50911 1 453
2 50912 1 453
2 50913 1 453
2 50914 1 453
2 50915 1 453
2 50916 1 453
2 50917 1 453
2 50918 1 453
2 50919 1 453
2 50920 1 453
2 50921 1 453
2 50922 1 454
2 50923 1 454
2 50924 1 454
2 50925 1 461
2 50926 1 461
2 50927 1 461
2 50928 1 461
2 50929 1 461
2 50930 1 461
2 50931 1 461
2 50932 1 461
2 50933 1 461
2 50934 1 461
2 50935 1 461
2 50936 1 461
2 50937 1 461
2 50938 1 461
2 50939 1 461
2 50940 1 461
2 50941 1 461
2 50942 1 461
2 50943 1 461
2 50944 1 461
2 50945 1 461
2 50946 1 461
2 50947 1 461
2 50948 1 461
2 50949 1 461
2 50950 1 461
2 50951 1 461
2 50952 1 461
2 50953 1 461
2 50954 1 461
2 50955 1 461
2 50956 1 461
2 50957 1 461
2 50958 1 461
2 50959 1 461
2 50960 1 461
2 50961 1 461
2 50962 1 461
2 50963 1 461
2 50964 1 461
2 50965 1 461
2 50966 1 461
2 50967 1 461
2 50968 1 462
2 50969 1 462
2 50970 1 462
2 50971 1 462
2 50972 1 462
2 50973 1 462
2 50974 1 462
2 50975 1 462
2 50976 1 462
2 50977 1 462
2 50978 1 462
2 50979 1 462
2 50980 1 462
2 50981 1 462
2 50982 1 462
2 50983 1 462
2 50984 1 462
2 50985 1 462
2 50986 1 462
2 50987 1 462
2 50988 1 462
2 50989 1 462
2 50990 1 462
2 50991 1 462
2 50992 1 462
2 50993 1 462
2 50994 1 462
2 50995 1 462
2 50996 1 462
2 50997 1 462
2 50998 1 462
2 50999 1 462
2 51000 1 462
2 51001 1 462
2 51002 1 462
2 51003 1 462
2 51004 1 462
2 51005 1 462
2 51006 1 462
2 51007 1 462
2 51008 1 462
2 51009 1 462
2 51010 1 462
2 51011 1 462
2 51012 1 462
2 51013 1 462
2 51014 1 462
2 51015 1 462
2 51016 1 462
2 51017 1 462
2 51018 1 462
2 51019 1 462
2 51020 1 462
2 51021 1 462
2 51022 1 462
2 51023 1 462
2 51024 1 462
2 51025 1 462
2 51026 1 462
2 51027 1 462
2 51028 1 462
2 51029 1 462
2 51030 1 462
2 51031 1 462
2 51032 1 462
2 51033 1 462
2 51034 1 462
2 51035 1 462
2 51036 1 462
2 51037 1 462
2 51038 1 462
2 51039 1 462
2 51040 1 462
2 51041 1 462
2 51042 1 462
2 51043 1 462
2 51044 1 462
2 51045 1 463
2 51046 1 463
2 51047 1 471
2 51048 1 471
2 51049 1 471
2 51050 1 471
2 51051 1 471
2 51052 1 471
2 51053 1 472
2 51054 1 472
2 51055 1 473
2 51056 1 473
2 51057 1 473
2 51058 1 473
2 51059 1 473
2 51060 1 473
2 51061 1 473
2 51062 1 473
2 51063 1 473
2 51064 1 474
2 51065 1 474
2 51066 1 474
2 51067 1 474
2 51068 1 474
2 51069 1 475
2 51070 1 475
2 51071 1 478
2 51072 1 478
2 51073 1 479
2 51074 1 479
2 51075 1 479
2 51076 1 479
2 51077 1 479
2 51078 1 479
2 51079 1 479
2 51080 1 479
2 51081 1 479
2 51082 1 479
2 51083 1 479
2 51084 1 479
2 51085 1 479
2 51086 1 479
2 51087 1 479
2 51088 1 479
2 51089 1 479
2 51090 1 479
2 51091 1 479
2 51092 1 479
2 51093 1 482
2 51094 1 482
2 51095 1 482
2 51096 1 482
2 51097 1 482
2 51098 1 482
2 51099 1 482
2 51100 1 482
2 51101 1 482
2 51102 1 482
2 51103 1 482
2 51104 1 482
2 51105 1 482
2 51106 1 483
2 51107 1 483
2 51108 1 483
2 51109 1 484
2 51110 1 484
2 51111 1 501
2 51112 1 501
2 51113 1 501
2 51114 1 501
2 51115 1 501
2 51116 1 501
2 51117 1 501
2 51118 1 501
2 51119 1 501
2 51120 1 501
2 51121 1 501
2 51122 1 501
2 51123 1 501
2 51124 1 501
2 51125 1 501
2 51126 1 501
2 51127 1 501
2 51128 1 501
2 51129 1 501
2 51130 1 501
2 51131 1 501
2 51132 1 501
2 51133 1 501
2 51134 1 501
2 51135 1 501
2 51136 1 501
2 51137 1 501
2 51138 1 501
2 51139 1 501
2 51140 1 501
2 51141 1 501
2 51142 1 501
2 51143 1 501
2 51144 1 501
2 51145 1 501
2 51146 1 501
2 51147 1 501
2 51148 1 501
2 51149 1 501
2 51150 1 501
2 51151 1 501
2 51152 1 501
2 51153 1 501
2 51154 1 501
2 51155 1 501
2 51156 1 501
2 51157 1 501
2 51158 1 501
2 51159 1 501
2 51160 1 501
2 51161 1 501
2 51162 1 502
2 51163 1 502
2 51164 1 502
2 51165 1 502
2 51166 1 502
2 51167 1 502
2 51168 1 502
2 51169 1 502
2 51170 1 502
2 51171 1 502
2 51172 1 502
2 51173 1 502
2 51174 1 502
2 51175 1 502
2 51176 1 502
2 51177 1 502
2 51178 1 502
2 51179 1 502
2 51180 1 502
2 51181 1 502
2 51182 1 502
2 51183 1 502
2 51184 1 502
2 51185 1 502
2 51186 1 502
2 51187 1 502
2 51188 1 502
2 51189 1 502
2 51190 1 502
2 51191 1 502
2 51192 1 503
2 51193 1 503
2 51194 1 503
2 51195 1 503
2 51196 1 504
2 51197 1 504
2 51198 1 504
2 51199 1 504
2 51200 1 504
2 51201 1 504
2 51202 1 504
2 51203 1 504
2 51204 1 504
2 51205 1 505
2 51206 1 505
2 51207 1 505
2 51208 1 505
2 51209 1 505
2 51210 1 505
2 51211 1 505
2 51212 1 505
2 51213 1 505
2 51214 1 505
2 51215 1 506
2 51216 1 506
2 51217 1 506
2 51218 1 506
2 51219 1 506
2 51220 1 506
2 51221 1 506
2 51222 1 506
2 51223 1 506
2 51224 1 506
2 51225 1 506
2 51226 1 506
2 51227 1 506
2 51228 1 506
2 51229 1 506
2 51230 1 506
2 51231 1 506
2 51232 1 506
2 51233 1 506
2 51234 1 506
2 51235 1 506
2 51236 1 506
2 51237 1 506
2 51238 1 506
2 51239 1 506
2 51240 1 506
2 51241 1 506
2 51242 1 507
2 51243 1 507
2 51244 1 507
2 51245 1 507
2 51246 1 507
2 51247 1 507
2 51248 1 507
2 51249 1 507
2 51250 1 507
2 51251 1 507
2 51252 1 507
2 51253 1 507
2 51254 1 507
2 51255 1 507
2 51256 1 507
2 51257 1 507
2 51258 1 508
2 51259 1 508
2 51260 1 508
2 51261 1 511
2 51262 1 511
2 51263 1 511
2 51264 1 511
2 51265 1 511
2 51266 1 511
2 51267 1 511
2 51268 1 511
2 51269 1 511
2 51270 1 511
2 51271 1 511
2 51272 1 511
2 51273 1 511
2 51274 1 512
2 51275 1 512
2 51276 1 512
2 51277 1 512
2 51278 1 512
2 51279 1 512
2 51280 1 512
2 51281 1 512
2 51282 1 512
2 51283 1 512
2 51284 1 512
2 51285 1 512
2 51286 1 512
2 51287 1 512
2 51288 1 512
2 51289 1 512
2 51290 1 512
2 51291 1 512
2 51292 1 512
2 51293 1 513
2 51294 1 513
2 51295 1 514
2 51296 1 514
2 51297 1 514
2 51298 1 514
2 51299 1 514
2 51300 1 514
2 51301 1 514
2 51302 1 514
2 51303 1 514
2 51304 1 514
2 51305 1 514
2 51306 1 517
2 51307 1 517
2 51308 1 517
2 51309 1 517
2 51310 1 517
2 51311 1 517
2 51312 1 517
2 51313 1 517
2 51314 1 517
2 51315 1 517
2 51316 1 517
2 51317 1 517
2 51318 1 517
2 51319 1 517
2 51320 1 517
2 51321 1 517
2 51322 1 517
2 51323 1 517
2 51324 1 518
2 51325 1 518
2 51326 1 519
2 51327 1 519
2 51328 1 519
2 51329 1 519
2 51330 1 519
2 51331 1 519
2 51332 1 519
2 51333 1 519
2 51334 1 519
2 51335 1 519
2 51336 1 519
2 51337 1 519
2 51338 1 519
2 51339 1 519
2 51340 1 519
2 51341 1 519
2 51342 1 519
2 51343 1 519
2 51344 1 519
2 51345 1 519
2 51346 1 519
2 51347 1 519
2 51348 1 519
2 51349 1 519
2 51350 1 519
2 51351 1 520
2 51352 1 520
2 51353 1 521
2 51354 1 521
2 51355 1 521
2 51356 1 521
2 51357 1 521
2 51358 1 528
2 51359 1 528
2 51360 1 528
2 51361 1 528
2 51362 1 528
2 51363 1 528
2 51364 1 528
2 51365 1 528
2 51366 1 528
2 51367 1 528
2 51368 1 529
2 51369 1 529
2 51370 1 529
2 51371 1 529
2 51372 1 530
2 51373 1 530
2 51374 1 530
2 51375 1 530
2 51376 1 530
2 51377 1 530
2 51378 1 530
2 51379 1 530
2 51380 1 530
2 51381 1 530
2 51382 1 530
2 51383 1 531
2 51384 1 531
2 51385 1 531
2 51386 1 531
2 51387 1 531
2 51388 1 531
2 51389 1 531
2 51390 1 539
2 51391 1 539
2 51392 1 539
2 51393 1 539
2 51394 1 539
2 51395 1 539
2 51396 1 539
2 51397 1 539
2 51398 1 539
2 51399 1 539
2 51400 1 539
2 51401 1 539
2 51402 1 539
2 51403 1 539
2 51404 1 539
2 51405 1 539
2 51406 1 539
2 51407 1 539
2 51408 1 539
2 51409 1 539
2 51410 1 539
2 51411 1 539
2 51412 1 539
2 51413 1 540
2 51414 1 540
2 51415 1 540
2 51416 1 540
2 51417 1 541
2 51418 1 541
2 51419 1 542
2 51420 1 542
2 51421 1 542
2 51422 1 545
2 51423 1 545
2 51424 1 545
2 51425 1 545
2 51426 1 545
2 51427 1 546
2 51428 1 546
2 51429 1 546
2 51430 1 546
2 51431 1 546
2 51432 1 546
2 51433 1 546
2 51434 1 546
2 51435 1 546
2 51436 1 546
2 51437 1 546
2 51438 1 546
2 51439 1 546
2 51440 1 546
2 51441 1 546
2 51442 1 546
2 51443 1 546
2 51444 1 546
2 51445 1 546
2 51446 1 546
2 51447 1 546
2 51448 1 547
2 51449 1 547
2 51450 1 548
2 51451 1 548
2 51452 1 548
2 51453 1 548
2 51454 1 548
2 51455 1 560
2 51456 1 560
2 51457 1 560
2 51458 1 560
2 51459 1 560
2 51460 1 561
2 51461 1 561
2 51462 1 561
2 51463 1 561
2 51464 1 561
2 51465 1 561
2 51466 1 561
2 51467 1 561
2 51468 1 561
2 51469 1 561
2 51470 1 562
2 51471 1 562
2 51472 1 562
2 51473 1 562
2 51474 1 562
2 51475 1 562
2 51476 1 562
2 51477 1 562
2 51478 1 562
2 51479 1 562
2 51480 1 562
2 51481 1 563
2 51482 1 563
2 51483 1 563
2 51484 1 565
2 51485 1 565
2 51486 1 568
2 51487 1 568
2 51488 1 569
2 51489 1 569
2 51490 1 572
2 51491 1 572
2 51492 1 572
2 51493 1 576
2 51494 1 576
2 51495 1 576
2 51496 1 576
2 51497 1 576
2 51498 1 576
2 51499 1 576
2 51500 1 576
2 51501 1 576
2 51502 1 576
2 51503 1 576
2 51504 1 576
2 51505 1 576
2 51506 1 576
2 51507 1 576
2 51508 1 576
2 51509 1 576
2 51510 1 576
2 51511 1 578
2 51512 1 578
2 51513 1 584
2 51514 1 584
2 51515 1 584
2 51516 1 585
2 51517 1 585
2 51518 1 585
2 51519 1 585
2 51520 1 586
2 51521 1 586
2 51522 1 586
2 51523 1 586
2 51524 1 586
2 51525 1 586
2 51526 1 586
2 51527 1 586
2 51528 1 586
2 51529 1 586
2 51530 1 586
2 51531 1 586
2 51532 1 586
2 51533 1 586
2 51534 1 587
2 51535 1 587
2 51536 1 588
2 51537 1 588
2 51538 1 588
2 51539 1 588
2 51540 1 589
2 51541 1 589
2 51542 1 589
2 51543 1 589
2 51544 1 595
2 51545 1 595
2 51546 1 595
2 51547 1 595
2 51548 1 595
2 51549 1 595
2 51550 1 595
2 51551 1 600
2 51552 1 600
2 51553 1 601
2 51554 1 601
2 51555 1 601
2 51556 1 601
2 51557 1 601
2 51558 1 601
2 51559 1 601
2 51560 1 601
2 51561 1 601
2 51562 1 601
2 51563 1 601
2 51564 1 601
2 51565 1 601
2 51566 1 601
2 51567 1 601
2 51568 1 601
2 51569 1 601
2 51570 1 601
2 51571 1 601
2 51572 1 601
2 51573 1 601
2 51574 1 609
2 51575 1 609
2 51576 1 610
2 51577 1 610
2 51578 1 610
2 51579 1 610
2 51580 1 610
2 51581 1 610
2 51582 1 610
2 51583 1 610
2 51584 1 610
2 51585 1 610
2 51586 1 610
2 51587 1 610
2 51588 1 610
2 51589 1 610
2 51590 1 610
2 51591 1 610
2 51592 1 610
2 51593 1 610
2 51594 1 610
2 51595 1 610
2 51596 1 610
2 51597 1 610
2 51598 1 610
2 51599 1 610
2 51600 1 610
2 51601 1 610
2 51602 1 610
2 51603 1 610
2 51604 1 610
2 51605 1 610
2 51606 1 610
2 51607 1 610
2 51608 1 610
2 51609 1 610
2 51610 1 610
2 51611 1 610
2 51612 1 610
2 51613 1 610
2 51614 1 610
2 51615 1 610
2 51616 1 610
2 51617 1 610
2 51618 1 610
2 51619 1 610
2 51620 1 610
2 51621 1 610
2 51622 1 610
2 51623 1 610
2 51624 1 610
2 51625 1 610
2 51626 1 611
2 51627 1 611
2 51628 1 611
2 51629 1 611
2 51630 1 611
2 51631 1 611
2 51632 1 611
2 51633 1 612
2 51634 1 612
2 51635 1 612
2 51636 1 612
2 51637 1 613
2 51638 1 613
2 51639 1 613
2 51640 1 613
2 51641 1 615
2 51642 1 615
2 51643 1 615
2 51644 1 615
2 51645 1 615
2 51646 1 623
2 51647 1 623
2 51648 1 623
2 51649 1 624
2 51650 1 624
2 51651 1 624
2 51652 1 631
2 51653 1 631
2 51654 1 631
2 51655 1 631
2 51656 1 631
2 51657 1 631
2 51658 1 631
2 51659 1 631
2 51660 1 631
2 51661 1 631
2 51662 1 631
2 51663 1 631
2 51664 1 631
2 51665 1 631
2 51666 1 631
2 51667 1 631
2 51668 1 631
2 51669 1 631
2 51670 1 631
2 51671 1 631
2 51672 1 631
2 51673 1 631
2 51674 1 631
2 51675 1 631
2 51676 1 631
2 51677 1 631
2 51678 1 631
2 51679 1 631
2 51680 1 631
2 51681 1 631
2 51682 1 631
2 51683 1 631
2 51684 1 631
2 51685 1 631
2 51686 1 631
2 51687 1 631
2 51688 1 631
2 51689 1 631
2 51690 1 631
2 51691 1 631
2 51692 1 631
2 51693 1 631
2 51694 1 633
2 51695 1 633
2 51696 1 633
2 51697 1 641
2 51698 1 641
2 51699 1 643
2 51700 1 643
2 51701 1 643
2 51702 1 643
2 51703 1 643
2 51704 1 643
2 51705 1 643
2 51706 1 643
2 51707 1 643
2 51708 1 643
2 51709 1 643
2 51710 1 643
2 51711 1 643
2 51712 1 644
2 51713 1 644
2 51714 1 644
2 51715 1 644
2 51716 1 644
2 51717 1 644
2 51718 1 644
2 51719 1 645
2 51720 1 645
2 51721 1 645
2 51722 1 645
2 51723 1 645
2 51724 1 645
2 51725 1 645
2 51726 1 645
2 51727 1 645
2 51728 1 645
2 51729 1 645
2 51730 1 645
2 51731 1 645
2 51732 1 645
2 51733 1 645
2 51734 1 645
2 51735 1 645
2 51736 1 645
2 51737 1 645
2 51738 1 646
2 51739 1 646
2 51740 1 646
2 51741 1 646
2 51742 1 646
2 51743 1 646
2 51744 1 646
2 51745 1 646
2 51746 1 646
2 51747 1 646
2 51748 1 646
2 51749 1 646
2 51750 1 646
2 51751 1 646
2 51752 1 646
2 51753 1 646
2 51754 1 646
2 51755 1 646
2 51756 1 646
2 51757 1 646
2 51758 1 646
2 51759 1 646
2 51760 1 646
2 51761 1 646
2 51762 1 646
2 51763 1 646
2 51764 1 646
2 51765 1 646
2 51766 1 646
2 51767 1 646
2 51768 1 646
2 51769 1 646
2 51770 1 646
2 51771 1 646
2 51772 1 646
2 51773 1 646
2 51774 1 646
2 51775 1 646
2 51776 1 647
2 51777 1 647
2 51778 1 647
2 51779 1 647
2 51780 1 648
2 51781 1 648
2 51782 1 654
2 51783 1 654
2 51784 1 654
2 51785 1 654
2 51786 1 655
2 51787 1 655
2 51788 1 655
2 51789 1 655
2 51790 1 655
2 51791 1 655
2 51792 1 655
2 51793 1 655
2 51794 1 655
2 51795 1 655
2 51796 1 655
2 51797 1 655
2 51798 1 655
2 51799 1 655
2 51800 1 655
2 51801 1 655
2 51802 1 655
2 51803 1 655
2 51804 1 655
2 51805 1 655
2 51806 1 655
2 51807 1 655
2 51808 1 655
2 51809 1 656
2 51810 1 656
2 51811 1 657
2 51812 1 657
2 51813 1 667
2 51814 1 667
2 51815 1 667
2 51816 1 667
2 51817 1 667
2 51818 1 667
2 51819 1 667
2 51820 1 667
2 51821 1 667
2 51822 1 668
2 51823 1 668
2 51824 1 668
2 51825 1 668
2 51826 1 668
2 51827 1 668
2 51828 1 669
2 51829 1 669
2 51830 1 670
2 51831 1 670
2 51832 1 670
2 51833 1 670
2 51834 1 670
2 51835 1 671
2 51836 1 671
2 51837 1 671
2 51838 1 671
2 51839 1 671
2 51840 1 671
2 51841 1 671
2 51842 1 671
2 51843 1 671
2 51844 1 671
2 51845 1 671
2 51846 1 680
2 51847 1 680
2 51848 1 680
2 51849 1 680
2 51850 1 680
2 51851 1 680
2 51852 1 680
2 51853 1 680
2 51854 1 680
2 51855 1 680
2 51856 1 680
2 51857 1 680
2 51858 1 680
2 51859 1 680
2 51860 1 680
2 51861 1 680
2 51862 1 680
2 51863 1 680
2 51864 1 680
2 51865 1 680
2 51866 1 683
2 51867 1 683
2 51868 1 683
2 51869 1 683
2 51870 1 684
2 51871 1 684
2 51872 1 684
2 51873 1 684
2 51874 1 685
2 51875 1 685
2 51876 1 685
2 51877 1 685
2 51878 1 685
2 51879 1 685
2 51880 1 686
2 51881 1 686
2 51882 1 686
2 51883 1 694
2 51884 1 694
2 51885 1 694
2 51886 1 694
2 51887 1 694
2 51888 1 694
2 51889 1 694
2 51890 1 694
2 51891 1 694
2 51892 1 694
2 51893 1 695
2 51894 1 695
2 51895 1 695
2 51896 1 695
2 51897 1 695
2 51898 1 695
2 51899 1 695
2 51900 1 695
2 51901 1 695
2 51902 1 695
2 51903 1 695
2 51904 1 695
2 51905 1 695
2 51906 1 695
2 51907 1 695
2 51908 1 695
2 51909 1 695
2 51910 1 695
2 51911 1 695
2 51912 1 695
2 51913 1 695
2 51914 1 695
2 51915 1 695
2 51916 1 695
2 51917 1 695
2 51918 1 695
2 51919 1 695
2 51920 1 695
2 51921 1 695
2 51922 1 695
2 51923 1 695
2 51924 1 695
2 51925 1 695
2 51926 1 695
2 51927 1 695
2 51928 1 695
2 51929 1 695
2 51930 1 695
2 51931 1 695
2 51932 1 695
2 51933 1 695
2 51934 1 695
2 51935 1 695
2 51936 1 695
2 51937 1 695
2 51938 1 695
2 51939 1 695
2 51940 1 695
2 51941 1 695
2 51942 1 695
2 51943 1 695
2 51944 1 695
2 51945 1 695
2 51946 1 695
2 51947 1 695
2 51948 1 695
2 51949 1 695
2 51950 1 695
2 51951 1 695
2 51952 1 695
2 51953 1 695
2 51954 1 695
2 51955 1 705
2 51956 1 705
2 51957 1 705
2 51958 1 705
2 51959 1 705
2 51960 1 705
2 51961 1 705
2 51962 1 705
2 51963 1 705
2 51964 1 705
2 51965 1 705
2 51966 1 705
2 51967 1 705
2 51968 1 705
2 51969 1 705
2 51970 1 705
2 51971 1 705
2 51972 1 705
2 51973 1 705
2 51974 1 705
2 51975 1 705
2 51976 1 705
2 51977 1 705
2 51978 1 705
2 51979 1 705
2 51980 1 705
2 51981 1 705
2 51982 1 705
2 51983 1 705
2 51984 1 705
2 51985 1 706
2 51986 1 706
2 51987 1 706
2 51988 1 706
2 51989 1 706
2 51990 1 706
2 51991 1 706
2 51992 1 706
2 51993 1 706
2 51994 1 706
2 51995 1 706
2 51996 1 706
2 51997 1 706
2 51998 1 706
2 51999 1 706
2 52000 1 706
2 52001 1 706
2 52002 1 706
2 52003 1 706
2 52004 1 706
2 52005 1 706
2 52006 1 706
2 52007 1 706
2 52008 1 706
2 52009 1 707
2 52010 1 707
2 52011 1 707
2 52012 1 707
2 52013 1 707
2 52014 1 707
2 52015 1 707
2 52016 1 707
2 52017 1 707
2 52018 1 707
2 52019 1 707
2 52020 1 707
2 52021 1 707
2 52022 1 707
2 52023 1 707
2 52024 1 707
2 52025 1 707
2 52026 1 707
2 52027 1 707
2 52028 1 707
2 52029 1 707
2 52030 1 707
2 52031 1 707
2 52032 1 707
2 52033 1 707
2 52034 1 707
2 52035 1 707
2 52036 1 707
2 52037 1 707
2 52038 1 707
2 52039 1 707
2 52040 1 707
2 52041 1 707
2 52042 1 707
2 52043 1 707
2 52044 1 707
2 52045 1 707
2 52046 1 707
2 52047 1 707
2 52048 1 707
2 52049 1 708
2 52050 1 708
2 52051 1 708
2 52052 1 708
2 52053 1 708
2 52054 1 708
2 52055 1 708
2 52056 1 708
2 52057 1 708
2 52058 1 708
2 52059 1 708
2 52060 1 708
2 52061 1 708
2 52062 1 708
2 52063 1 708
2 52064 1 708
2 52065 1 708
2 52066 1 708
2 52067 1 708
2 52068 1 708
2 52069 1 709
2 52070 1 709
2 52071 1 709
2 52072 1 709
2 52073 1 709
2 52074 1 709
2 52075 1 709
2 52076 1 709
2 52077 1 709
2 52078 1 709
2 52079 1 709
2 52080 1 709
2 52081 1 709
2 52082 1 710
2 52083 1 710
2 52084 1 710
2 52085 1 710
2 52086 1 710
2 52087 1 711
2 52088 1 711
2 52089 1 711
2 52090 1 711
2 52091 1 711
2 52092 1 711
2 52093 1 711
2 52094 1 711
2 52095 1 711
2 52096 1 711
2 52097 1 711
2 52098 1 711
2 52099 1 711
2 52100 1 711
2 52101 1 711
2 52102 1 711
2 52103 1 711
2 52104 1 711
2 52105 1 711
2 52106 1 711
2 52107 1 711
2 52108 1 712
2 52109 1 712
2 52110 1 714
2 52111 1 714
2 52112 1 714
2 52113 1 715
2 52114 1 715
2 52115 1 715
2 52116 1 715
2 52117 1 716
2 52118 1 716
2 52119 1 716
2 52120 1 716
2 52121 1 716
2 52122 1 716
2 52123 1 716
2 52124 1 717
2 52125 1 717
2 52126 1 717
2 52127 1 717
2 52128 1 718
2 52129 1 718
2 52130 1 718
2 52131 1 718
2 52132 1 718
2 52133 1 718
2 52134 1 718
2 52135 1 718
2 52136 1 718
2 52137 1 718
2 52138 1 718
2 52139 1 718
2 52140 1 721
2 52141 1 721
2 52142 1 722
2 52143 1 722
2 52144 1 722
2 52145 1 722
2 52146 1 722
2 52147 1 722
2 52148 1 722
2 52149 1 722
2 52150 1 725
2 52151 1 725
2 52152 1 725
2 52153 1 725
2 52154 1 725
2 52155 1 725
2 52156 1 725
2 52157 1 725
2 52158 1 725
2 52159 1 725
2 52160 1 725
2 52161 1 725
2 52162 1 725
2 52163 1 725
2 52164 1 725
2 52165 1 725
2 52166 1 725
2 52167 1 725
2 52168 1 725
2 52169 1 725
2 52170 1 725
2 52171 1 725
2 52172 1 725
2 52173 1 726
2 52174 1 726
2 52175 1 728
2 52176 1 728
2 52177 1 728
2 52178 1 728
2 52179 1 728
2 52180 1 728
2 52181 1 728
2 52182 1 729
2 52183 1 729
2 52184 1 729
2 52185 1 729
2 52186 1 729
2 52187 1 729
2 52188 1 729
2 52189 1 730
2 52190 1 730
2 52191 1 730
2 52192 1 730
2 52193 1 730
2 52194 1 730
2 52195 1 731
2 52196 1 731
2 52197 1 731
2 52198 1 731
2 52199 1 732
2 52200 1 732
2 52201 1 732
2 52202 1 733
2 52203 1 733
2 52204 1 736
2 52205 1 736
2 52206 1 736
2 52207 1 744
2 52208 1 744
2 52209 1 744
2 52210 1 745
2 52211 1 745
2 52212 1 745
2 52213 1 745
2 52214 1 745
2 52215 1 745
2 52216 1 746
2 52217 1 746
2 52218 1 747
2 52219 1 747
2 52220 1 747
2 52221 1 747
2 52222 1 747
2 52223 1 747
2 52224 1 747
2 52225 1 747
2 52226 1 747
2 52227 1 750
2 52228 1 750
2 52229 1 750
2 52230 1 751
2 52231 1 751
2 52232 1 751
2 52233 1 751
2 52234 1 751
2 52235 1 751
2 52236 1 751
2 52237 1 751
2 52238 1 751
2 52239 1 751
2 52240 1 751
2 52241 1 751
2 52242 1 751
2 52243 1 754
2 52244 1 754
2 52245 1 754
2 52246 1 754
2 52247 1 754
2 52248 1 755
2 52249 1 755
2 52250 1 755
2 52251 1 755
2 52252 1 755
2 52253 1 755
2 52254 1 755
2 52255 1 764
2 52256 1 764
2 52257 1 765
2 52258 1 765
2 52259 1 765
2 52260 1 765
2 52261 1 765
2 52262 1 765
2 52263 1 779
2 52264 1 779
2 52265 1 779
2 52266 1 779
2 52267 1 779
2 52268 1 779
2 52269 1 779
2 52270 1 779
2 52271 1 779
2 52272 1 779
2 52273 1 780
2 52274 1 780
2 52275 1 780
2 52276 1 780
2 52277 1 780
2 52278 1 780
2 52279 1 780
2 52280 1 780
2 52281 1 780
2 52282 1 780
2 52283 1 782
2 52284 1 782
2 52285 1 782
2 52286 1 782
2 52287 1 782
2 52288 1 783
2 52289 1 783
2 52290 1 792
2 52291 1 792
2 52292 1 792
2 52293 1 792
2 52294 1 792
2 52295 1 792
2 52296 1 792
2 52297 1 792
2 52298 1 792
2 52299 1 792
2 52300 1 792
2 52301 1 792
2 52302 1 792
2 52303 1 792
2 52304 1 792
2 52305 1 793
2 52306 1 793
2 52307 1 793
2 52308 1 793
2 52309 1 793
2 52310 1 794
2 52311 1 794
2 52312 1 794
2 52313 1 794
2 52314 1 794
2 52315 1 794
2 52316 1 794
2 52317 1 794
2 52318 1 794
2 52319 1 794
2 52320 1 794
2 52321 1 794
2 52322 1 794
2 52323 1 794
2 52324 1 794
2 52325 1 795
2 52326 1 795
2 52327 1 795
2 52328 1 795
2 52329 1 795
2 52330 1 795
2 52331 1 795
2 52332 1 795
2 52333 1 795
2 52334 1 795
2 52335 1 795
2 52336 1 796
2 52337 1 796
2 52338 1 796
2 52339 1 797
2 52340 1 797
2 52341 1 798
2 52342 1 798
2 52343 1 798
2 52344 1 798
2 52345 1 799
2 52346 1 799
2 52347 1 799
2 52348 1 799
2 52349 1 801
2 52350 1 801
2 52351 1 802
2 52352 1 802
2 52353 1 802
2 52354 1 802
2 52355 1 802
2 52356 1 803
2 52357 1 803
2 52358 1 803
2 52359 1 803
2 52360 1 803
2 52361 1 803
2 52362 1 803
2 52363 1 803
2 52364 1 805
2 52365 1 805
2 52366 1 805
2 52367 1 806
2 52368 1 806
2 52369 1 806
2 52370 1 806
2 52371 1 806
2 52372 1 806
2 52373 1 806
2 52374 1 806
2 52375 1 806
2 52376 1 806
2 52377 1 806
2 52378 1 806
2 52379 1 806
2 52380 1 806
2 52381 1 806
2 52382 1 806
2 52383 1 806
2 52384 1 806
2 52385 1 806
2 52386 1 806
2 52387 1 806
2 52388 1 806
2 52389 1 806
2 52390 1 806
2 52391 1 806
2 52392 1 806
2 52393 1 806
2 52394 1 806
2 52395 1 806
2 52396 1 807
2 52397 1 807
2 52398 1 807
2 52399 1 807
2 52400 1 807
2 52401 1 807
2 52402 1 808
2 52403 1 808
2 52404 1 808
2 52405 1 808
2 52406 1 808
2 52407 1 808
2 52408 1 808
2 52409 1 809
2 52410 1 809
2 52411 1 809
2 52412 1 814
2 52413 1 814
2 52414 1 823
2 52415 1 823
2 52416 1 823
2 52417 1 824
2 52418 1 824
2 52419 1 824
2 52420 1 826
2 52421 1 826
2 52422 1 826
2 52423 1 831
2 52424 1 831
2 52425 1 831
2 52426 1 835
2 52427 1 835
2 52428 1 835
2 52429 1 835
2 52430 1 837
2 52431 1 837
2 52432 1 837
2 52433 1 837
2 52434 1 837
2 52435 1 837
2 52436 1 837
2 52437 1 840
2 52438 1 840
2 52439 1 841
2 52440 1 841
2 52441 1 841
2 52442 1 842
2 52443 1 842
2 52444 1 849
2 52445 1 849
2 52446 1 849
2 52447 1 849
2 52448 1 849
2 52449 1 849
2 52450 1 849
2 52451 1 849
2 52452 1 849
2 52453 1 849
2 52454 1 849
2 52455 1 849
2 52456 1 849
2 52457 1 849
2 52458 1 850
2 52459 1 850
2 52460 1 852
2 52461 1 852
2 52462 1 852
2 52463 1 852
2 52464 1 852
2 52465 1 855
2 52466 1 855
2 52467 1 855
2 52468 1 855
2 52469 1 856
2 52470 1 856
2 52471 1 863
2 52472 1 863
2 52473 1 863
2 52474 1 863
2 52475 1 863
2 52476 1 863
2 52477 1 863
2 52478 1 863
2 52479 1 863
2 52480 1 863
2 52481 1 863
2 52482 1 863
2 52483 1 863
2 52484 1 863
2 52485 1 863
2 52486 1 863
2 52487 1 863
2 52488 1 863
2 52489 1 863
2 52490 1 863
2 52491 1 863
2 52492 1 864
2 52493 1 864
2 52494 1 864
2 52495 1 865
2 52496 1 865
2 52497 1 865
2 52498 1 865
2 52499 1 865
2 52500 1 865
2 52501 1 865
2 52502 1 865
2 52503 1 865
2 52504 1 865
2 52505 1 865
2 52506 1 865
2 52507 1 865
2 52508 1 865
2 52509 1 865
2 52510 1 865
2 52511 1 865
2 52512 1 866
2 52513 1 866
2 52514 1 866
2 52515 1 873
2 52516 1 873
2 52517 1 873
2 52518 1 873
2 52519 1 873
2 52520 1 873
2 52521 1 875
2 52522 1 875
2 52523 1 875
2 52524 1 901
2 52525 1 901
2 52526 1 901
2 52527 1 901
2 52528 1 902
2 52529 1 902
2 52530 1 902
2 52531 1 902
2 52532 1 905
2 52533 1 905
2 52534 1 905
2 52535 1 905
2 52536 1 905
2 52537 1 906
2 52538 1 906
2 52539 1 906
2 52540 1 907
2 52541 1 907
2 52542 1 907
2 52543 1 907
2 52544 1 909
2 52545 1 909
2 52546 1 909
2 52547 1 910
2 52548 1 910
2 52549 1 916
2 52550 1 916
2 52551 1 916
2 52552 1 916
2 52553 1 916
2 52554 1 918
2 52555 1 918
2 52556 1 919
2 52557 1 919
2 52558 1 923
2 52559 1 923
2 52560 1 923
2 52561 1 923
2 52562 1 923
2 52563 1 923
2 52564 1 923
2 52565 1 923
2 52566 1 923
2 52567 1 925
2 52568 1 925
2 52569 1 925
2 52570 1 925
2 52571 1 925
2 52572 1 925
2 52573 1 925
2 52574 1 925
2 52575 1 925
2 52576 1 925
2 52577 1 925
2 52578 1 925
2 52579 1 925
2 52580 1 925
2 52581 1 925
2 52582 1 925
2 52583 1 925
2 52584 1 925
2 52585 1 925
2 52586 1 925
2 52587 1 925
2 52588 1 925
2 52589 1 925
2 52590 1 925
2 52591 1 925
2 52592 1 925
2 52593 1 925
2 52594 1 925
2 52595 1 925
2 52596 1 925
2 52597 1 925
2 52598 1 925
2 52599 1 925
2 52600 1 925
2 52601 1 925
2 52602 1 926
2 52603 1 926
2 52604 1 926
2 52605 1 926
2 52606 1 926
2 52607 1 926
2 52608 1 926
2 52609 1 926
2 52610 1 926
2 52611 1 926
2 52612 1 926
2 52613 1 926
2 52614 1 926
2 52615 1 926
2 52616 1 926
2 52617 1 926
2 52618 1 926
2 52619 1 926
2 52620 1 926
2 52621 1 926
2 52622 1 926
2 52623 1 926
2 52624 1 926
2 52625 1 926
2 52626 1 926
2 52627 1 926
2 52628 1 926
2 52629 1 926
2 52630 1 926
2 52631 1 926
2 52632 1 926
2 52633 1 926
2 52634 1 926
2 52635 1 926
2 52636 1 926
2 52637 1 926
2 52638 1 926
2 52639 1 926
2 52640 1 926
2 52641 1 926
2 52642 1 926
2 52643 1 926
2 52644 1 926
2 52645 1 926
2 52646 1 926
2 52647 1 926
2 52648 1 926
2 52649 1 926
2 52650 1 926
2 52651 1 926
2 52652 1 926
2 52653 1 926
2 52654 1 926
2 52655 1 926
2 52656 1 927
2 52657 1 927
2 52658 1 928
2 52659 1 928
2 52660 1 928
2 52661 1 928
2 52662 1 928
2 52663 1 928
2 52664 1 928
2 52665 1 928
2 52666 1 928
2 52667 1 928
2 52668 1 928
2 52669 1 929
2 52670 1 929
2 52671 1 929
2 52672 1 930
2 52673 1 930
2 52674 1 930
2 52675 1 930
2 52676 1 930
2 52677 1 930
2 52678 1 931
2 52679 1 931
2 52680 1 932
2 52681 1 932
2 52682 1 932
2 52683 1 932
2 52684 1 933
2 52685 1 933
2 52686 1 933
2 52687 1 933
2 52688 1 933
2 52689 1 933
2 52690 1 934
2 52691 1 934
2 52692 1 934
2 52693 1 934
2 52694 1 935
2 52695 1 935
2 52696 1 935
2 52697 1 939
2 52698 1 939
2 52699 1 939
2 52700 1 939
2 52701 1 939
2 52702 1 940
2 52703 1 940
2 52704 1 942
2 52705 1 942
2 52706 1 942
2 52707 1 942
2 52708 1 942
2 52709 1 943
2 52710 1 943
2 52711 1 943
2 52712 1 943
2 52713 1 943
2 52714 1 944
2 52715 1 944
2 52716 1 944
2 52717 1 944
2 52718 1 944
2 52719 1 944
2 52720 1 944
2 52721 1 944
2 52722 1 944
2 52723 1 946
2 52724 1 946
2 52725 1 948
2 52726 1 948
2 52727 1 950
2 52728 1 950
2 52729 1 950
2 52730 1 950
2 52731 1 950
2 52732 1 950
2 52733 1 952
2 52734 1 952
2 52735 1 964
2 52736 1 964
2 52737 1 964
2 52738 1 966
2 52739 1 966
2 52740 1 966
2 52741 1 966
2 52742 1 966
2 52743 1 966
2 52744 1 966
2 52745 1 966
2 52746 1 966
2 52747 1 966
2 52748 1 966
2 52749 1 966
2 52750 1 966
2 52751 1 966
2 52752 1 966
2 52753 1 966
2 52754 1 966
2 52755 1 966
2 52756 1 967
2 52757 1 967
2 52758 1 967
2 52759 1 967
2 52760 1 968
2 52761 1 968
2 52762 1 968
2 52763 1 971
2 52764 1 971
2 52765 1 971
2 52766 1 971
2 52767 1 971
2 52768 1 971
2 52769 1 971
2 52770 1 971
2 52771 1 971
2 52772 1 972
2 52773 1 972
2 52774 1 985
2 52775 1 985
2 52776 1 985
2 52777 1 985
2 52778 1 985
2 52779 1 985
2 52780 1 985
2 52781 1 985
2 52782 1 985
2 52783 1 985
2 52784 1 985
2 52785 1 985
2 52786 1 985
2 52787 1 985
2 52788 1 985
2 52789 1 985
2 52790 1 985
2 52791 1 985
2 52792 1 985
2 52793 1 985
2 52794 1 985
2 52795 1 986
2 52796 1 986
2 52797 1 986
2 52798 1 987
2 52799 1 987
2 52800 1 987
2 52801 1 988
2 52802 1 988
2 52803 1 988
2 52804 1 988
2 52805 1 988
2 52806 1 988
2 52807 1 988
2 52808 1 988
2 52809 1 988
2 52810 1 989
2 52811 1 989
2 52812 1 990
2 52813 1 990
2 52814 1 990
2 52815 1 990
2 52816 1 991
2 52817 1 991
2 52818 1 991
2 52819 1 991
2 52820 1 992
2 52821 1 992
2 52822 1 993
2 52823 1 993
2 52824 1 994
2 52825 1 994
2 52826 1 995
2 52827 1 995
2 52828 1 998
2 52829 1 998
2 52830 1 998
2 52831 1 998
2 52832 1 998
2 52833 1 998
2 52834 1 999
2 52835 1 999
2 52836 1 999
2 52837 1 1000
2 52838 1 1000
2 52839 1 1000
2 52840 1 1000
2 52841 1 1000
2 52842 1 1000
2 52843 1 1000
2 52844 1 1000
2 52845 1 1000
2 52846 1 1000
2 52847 1 1000
2 52848 1 1000
2 52849 1 1000
2 52850 1 1000
2 52851 1 1000
2 52852 1 1000
2 52853 1 1000
2 52854 1 1000
2 52855 1 1000
2 52856 1 1001
2 52857 1 1001
2 52858 1 1001
2 52859 1 1002
2 52860 1 1002
2 52861 1 1002
2 52862 1 1003
2 52863 1 1003
2 52864 1 1004
2 52865 1 1004
2 52866 1 1013
2 52867 1 1013
2 52868 1 1013
2 52869 1 1013
2 52870 1 1013
2 52871 1 1013
2 52872 1 1013
2 52873 1 1013
2 52874 1 1013
2 52875 1 1013
2 52876 1 1013
2 52877 1 1014
2 52878 1 1014
2 52879 1 1015
2 52880 1 1015
2 52881 1 1016
2 52882 1 1016
2 52883 1 1029
2 52884 1 1029
2 52885 1 1029
2 52886 1 1030
2 52887 1 1030
2 52888 1 1030
2 52889 1 1030
2 52890 1 1030
2 52891 1 1030
2 52892 1 1030
2 52893 1 1030
2 52894 1 1030
2 52895 1 1030
2 52896 1 1030
2 52897 1 1030
2 52898 1 1030
2 52899 1 1030
2 52900 1 1030
2 52901 1 1030
2 52902 1 1030
2 52903 1 1030
2 52904 1 1030
2 52905 1 1030
2 52906 1 1030
2 52907 1 1030
2 52908 1 1030
2 52909 1 1030
2 52910 1 1032
2 52911 1 1032
2 52912 1 1032
2 52913 1 1033
2 52914 1 1033
2 52915 1 1033
2 52916 1 1033
2 52917 1 1033
2 52918 1 1033
2 52919 1 1033
2 52920 1 1033
2 52921 1 1033
2 52922 1 1033
2 52923 1 1033
2 52924 1 1034
2 52925 1 1034
2 52926 1 1034
2 52927 1 1034
2 52928 1 1034
2 52929 1 1034
2 52930 1 1041
2 52931 1 1041
2 52932 1 1041
2 52933 1 1041
2 52934 1 1041
2 52935 1 1041
2 52936 1 1041
2 52937 1 1041
2 52938 1 1041
2 52939 1 1042
2 52940 1 1042
2 52941 1 1042
2 52942 1 1042
2 52943 1 1042
2 52944 1 1042
2 52945 1 1044
2 52946 1 1044
2 52947 1 1052
2 52948 1 1052
2 52949 1 1052
2 52950 1 1052
2 52951 1 1052
2 52952 1 1052
2 52953 1 1052
2 52954 1 1052
2 52955 1 1052
2 52956 1 1052
2 52957 1 1052
2 52958 1 1052
2 52959 1 1052
2 52960 1 1052
2 52961 1 1052
2 52962 1 1052
2 52963 1 1052
2 52964 1 1052
2 52965 1 1052
2 52966 1 1054
2 52967 1 1054
2 52968 1 1054
2 52969 1 1054
2 52970 1 1054
2 52971 1 1054
2 52972 1 1054
2 52973 1 1055
2 52974 1 1055
2 52975 1 1056
2 52976 1 1056
2 52977 1 1056
2 52978 1 1056
2 52979 1 1056
2 52980 1 1056
2 52981 1 1056
2 52982 1 1056
2 52983 1 1056
2 52984 1 1057
2 52985 1 1057
2 52986 1 1058
2 52987 1 1058
2 52988 1 1059
2 52989 1 1059
2 52990 1 1060
2 52991 1 1060
2 52992 1 1060
2 52993 1 1060
2 52994 1 1060
2 52995 1 1062
2 52996 1 1062
2 52997 1 1062
2 52998 1 1062
2 52999 1 1062
2 53000 1 1062
2 53001 1 1062
2 53002 1 1062
2 53003 1 1062
2 53004 1 1064
2 53005 1 1064
2 53006 1 1064
2 53007 1 1064
2 53008 1 1064
2 53009 1 1066
2 53010 1 1066
2 53011 1 1066
2 53012 1 1066
2 53013 1 1067
2 53014 1 1067
2 53015 1 1067
2 53016 1 1067
2 53017 1 1067
2 53018 1 1083
2 53019 1 1083
2 53020 1 1083
2 53021 1 1083
2 53022 1 1083
2 53023 1 1083
2 53024 1 1084
2 53025 1 1084
2 53026 1 1084
2 53027 1 1084
2 53028 1 1084
2 53029 1 1084
2 53030 1 1084
2 53031 1 1084
2 53032 1 1084
2 53033 1 1084
2 53034 1 1084
2 53035 1 1084
2 53036 1 1084
2 53037 1 1084
2 53038 1 1084
2 53039 1 1084
2 53040 1 1084
2 53041 1 1086
2 53042 1 1086
2 53043 1 1086
2 53044 1 1086
2 53045 1 1086
2 53046 1 1086
2 53047 1 1086
2 53048 1 1086
2 53049 1 1086
2 53050 1 1087
2 53051 1 1087
2 53052 1 1095
2 53053 1 1095
2 53054 1 1095
2 53055 1 1095
2 53056 1 1095
2 53057 1 1095
2 53058 1 1095
2 53059 1 1095
2 53060 1 1096
2 53061 1 1096
2 53062 1 1096
2 53063 1 1096
2 53064 1 1096
2 53065 1 1097
2 53066 1 1097
2 53067 1 1097
2 53068 1 1097
2 53069 1 1097
2 53070 1 1097
2 53071 1 1097
2 53072 1 1097
2 53073 1 1097
2 53074 1 1098
2 53075 1 1098
2 53076 1 1098
2 53077 1 1098
2 53078 1 1100
2 53079 1 1100
2 53080 1 1100
2 53081 1 1115
2 53082 1 1115
2 53083 1 1115
2 53084 1 1115
2 53085 1 1115
2 53086 1 1115
2 53087 1 1115
2 53088 1 1115
2 53089 1 1115
2 53090 1 1115
2 53091 1 1116
2 53092 1 1116
2 53093 1 1117
2 53094 1 1117
2 53095 1 1117
2 53096 1 1117
2 53097 1 1117
2 53098 1 1117
2 53099 1 1125
2 53100 1 1125
2 53101 1 1137
2 53102 1 1137
2 53103 1 1137
2 53104 1 1137
2 53105 1 1137
2 53106 1 1137
2 53107 1 1137
2 53108 1 1137
2 53109 1 1137
2 53110 1 1137
2 53111 1 1137
2 53112 1 1137
2 53113 1 1137
2 53114 1 1137
2 53115 1 1137
2 53116 1 1137
2 53117 1 1137
2 53118 1 1137
2 53119 1 1137
2 53120 1 1137
2 53121 1 1137
2 53122 1 1137
2 53123 1 1137
2 53124 1 1137
2 53125 1 1137
2 53126 1 1137
2 53127 1 1137
2 53128 1 1137
2 53129 1 1138
2 53130 1 1138
2 53131 1 1138
2 53132 1 1138
2 53133 1 1138
2 53134 1 1138
2 53135 1 1138
2 53136 1 1138
2 53137 1 1138
2 53138 1 1138
2 53139 1 1138
2 53140 1 1138
2 53141 1 1138
2 53142 1 1138
2 53143 1 1138
2 53144 1 1138
2 53145 1 1138
2 53146 1 1138
2 53147 1 1138
2 53148 1 1138
2 53149 1 1139
2 53150 1 1139
2 53151 1 1139
2 53152 1 1139
2 53153 1 1141
2 53154 1 1141
2 53155 1 1141
2 53156 1 1142
2 53157 1 1142
2 53158 1 1142
2 53159 1 1142
2 53160 1 1142
2 53161 1 1142
2 53162 1 1142
2 53163 1 1142
2 53164 1 1142
2 53165 1 1142
2 53166 1 1142
2 53167 1 1142
2 53168 1 1142
2 53169 1 1142
2 53170 1 1142
2 53171 1 1142
2 53172 1 1142
2 53173 1 1144
2 53174 1 1144
2 53175 1 1144
2 53176 1 1144
2 53177 1 1144
2 53178 1 1144
2 53179 1 1151
2 53180 1 1151
2 53181 1 1151
2 53182 1 1151
2 53183 1 1151
2 53184 1 1151
2 53185 1 1151
2 53186 1 1151
2 53187 1 1151
2 53188 1 1151
2 53189 1 1151
2 53190 1 1153
2 53191 1 1153
2 53192 1 1153
2 53193 1 1153
2 53194 1 1153
2 53195 1 1153
2 53196 1 1153
2 53197 1 1153
2 53198 1 1153
2 53199 1 1153
2 53200 1 1153
2 53201 1 1153
2 53202 1 1153
2 53203 1 1153
2 53204 1 1153
2 53205 1 1153
2 53206 1 1153
2 53207 1 1153
2 53208 1 1153
2 53209 1 1155
2 53210 1 1155
2 53211 1 1155
2 53212 1 1155
2 53213 1 1155
2 53214 1 1155
2 53215 1 1155
2 53216 1 1155
2 53217 1 1155
2 53218 1 1156
2 53219 1 1156
2 53220 1 1156
2 53221 1 1156
2 53222 1 1156
2 53223 1 1156
2 53224 1 1156
2 53225 1 1156
2 53226 1 1156
2 53227 1 1156
2 53228 1 1156
2 53229 1 1156
2 53230 1 1156
2 53231 1 1156
2 53232 1 1156
2 53233 1 1156
2 53234 1 1156
2 53235 1 1156
2 53236 1 1156
2 53237 1 1156
2 53238 1 1156
2 53239 1 1156
2 53240 1 1156
2 53241 1 1156
2 53242 1 1156
2 53243 1 1156
2 53244 1 1156
2 53245 1 1156
2 53246 1 1156
2 53247 1 1156
2 53248 1 1156
2 53249 1 1156
2 53250 1 1156
2 53251 1 1156
2 53252 1 1156
2 53253 1 1156
2 53254 1 1156
2 53255 1 1156
2 53256 1 1156
2 53257 1 1156
2 53258 1 1156
2 53259 1 1156
2 53260 1 1156
2 53261 1 1156
2 53262 1 1156
2 53263 1 1156
2 53264 1 1156
2 53265 1 1156
2 53266 1 1156
2 53267 1 1156
2 53268 1 1156
2 53269 1 1156
2 53270 1 1156
2 53271 1 1156
2 53272 1 1156
2 53273 1 1156
2 53274 1 1156
2 53275 1 1156
2 53276 1 1156
2 53277 1 1156
2 53278 1 1156
2 53279 1 1156
2 53280 1 1156
2 53281 1 1156
2 53282 1 1156
2 53283 1 1156
2 53284 1 1156
2 53285 1 1156
2 53286 1 1156
2 53287 1 1156
2 53288 1 1156
2 53289 1 1156
2 53290 1 1156
2 53291 1 1156
2 53292 1 1156
2 53293 1 1156
2 53294 1 1156
2 53295 1 1156
2 53296 1 1156
2 53297 1 1156
2 53298 1 1156
2 53299 1 1157
2 53300 1 1157
2 53301 1 1157
2 53302 1 1157
2 53303 1 1157
2 53304 1 1157
2 53305 1 1157
2 53306 1 1157
2 53307 1 1157
2 53308 1 1157
2 53309 1 1157
2 53310 1 1157
2 53311 1 1157
2 53312 1 1157
2 53313 1 1157
2 53314 1 1157
2 53315 1 1158
2 53316 1 1158
2 53317 1 1158
2 53318 1 1163
2 53319 1 1163
2 53320 1 1171
2 53321 1 1171
2 53322 1 1172
2 53323 1 1172
2 53324 1 1172
2 53325 1 1179
2 53326 1 1179
2 53327 1 1179
2 53328 1 1179
2 53329 1 1179
2 53330 1 1180
2 53331 1 1180
2 53332 1 1180
2 53333 1 1189
2 53334 1 1189
2 53335 1 1189
2 53336 1 1189
2 53337 1 1189
2 53338 1 1189
2 53339 1 1189
2 53340 1 1189
2 53341 1 1189
2 53342 1 1189
2 53343 1 1190
2 53344 1 1190
2 53345 1 1190
2 53346 1 1190
2 53347 1 1190
2 53348 1 1190
2 53349 1 1190
2 53350 1 1190
2 53351 1 1193
2 53352 1 1193
2 53353 1 1193
2 53354 1 1193
2 53355 1 1193
2 53356 1 1193
2 53357 1 1193
2 53358 1 1193
2 53359 1 1193
2 53360 1 1193
2 53361 1 1193
2 53362 1 1193
2 53363 1 1193
2 53364 1 1193
2 53365 1 1193
2 53366 1 1193
2 53367 1 1193
2 53368 1 1193
2 53369 1 1194
2 53370 1 1194
2 53371 1 1196
2 53372 1 1196
2 53373 1 1199
2 53374 1 1199
2 53375 1 1199
2 53376 1 1200
2 53377 1 1200
2 53378 1 1200
2 53379 1 1200
2 53380 1 1200
2 53381 1 1200
2 53382 1 1201
2 53383 1 1201
2 53384 1 1202
2 53385 1 1202
2 53386 1 1203
2 53387 1 1203
2 53388 1 1203
2 53389 1 1203
2 53390 1 1203
2 53391 1 1203
2 53392 1 1206
2 53393 1 1206
2 53394 1 1206
2 53395 1 1206
2 53396 1 1206
2 53397 1 1206
2 53398 1 1206
2 53399 1 1206
2 53400 1 1206
2 53401 1 1206
2 53402 1 1215
2 53403 1 1215
2 53404 1 1216
2 53405 1 1216
2 53406 1 1219
2 53407 1 1219
2 53408 1 1219
2 53409 1 1219
2 53410 1 1219
2 53411 1 1219
2 53412 1 1220
2 53413 1 1220
2 53414 1 1220
2 53415 1 1220
2 53416 1 1220
2 53417 1 1220
2 53418 1 1220
2 53419 1 1220
2 53420 1 1220
2 53421 1 1220
2 53422 1 1220
2 53423 1 1220
2 53424 1 1220
2 53425 1 1220
2 53426 1 1220
2 53427 1 1220
2 53428 1 1220
2 53429 1 1220
2 53430 1 1220
2 53431 1 1220
2 53432 1 1220
2 53433 1 1220
2 53434 1 1220
2 53435 1 1220
2 53436 1 1220
2 53437 1 1229
2 53438 1 1229
2 53439 1 1229
2 53440 1 1229
2 53441 1 1229
2 53442 1 1229
2 53443 1 1229
2 53444 1 1230
2 53445 1 1230
2 53446 1 1230
2 53447 1 1230
2 53448 1 1232
2 53449 1 1232
2 53450 1 1232
2 53451 1 1234
2 53452 1 1234
2 53453 1 1237
2 53454 1 1237
2 53455 1 1237
2 53456 1 1238
2 53457 1 1238
2 53458 1 1238
2 53459 1 1239
2 53460 1 1239
2 53461 1 1239
2 53462 1 1239
2 53463 1 1239
2 53464 1 1239
2 53465 1 1239
2 53466 1 1239
2 53467 1 1239
2 53468 1 1239
2 53469 1 1239
2 53470 1 1241
2 53471 1 1241
2 53472 1 1256
2 53473 1 1256
2 53474 1 1256
2 53475 1 1256
2 53476 1 1256
2 53477 1 1256
2 53478 1 1256
2 53479 1 1256
2 53480 1 1257
2 53481 1 1257
2 53482 1 1257
2 53483 1 1259
2 53484 1 1259
2 53485 1 1259
2 53486 1 1260
2 53487 1 1260
2 53488 1 1262
2 53489 1 1262
2 53490 1 1264
2 53491 1 1264
2 53492 1 1271
2 53493 1 1271
2 53494 1 1271
2 53495 1 1271
2 53496 1 1272
2 53497 1 1272
2 53498 1 1272
2 53499 1 1272
2 53500 1 1273
2 53501 1 1273
2 53502 1 1284
2 53503 1 1284
2 53504 1 1284
2 53505 1 1284
2 53506 1 1284
2 53507 1 1285
2 53508 1 1285
2 53509 1 1286
2 53510 1 1286
2 53511 1 1299
2 53512 1 1299
2 53513 1 1299
2 53514 1 1299
2 53515 1 1300
2 53516 1 1300
2 53517 1 1310
2 53518 1 1310
2 53519 1 1310
2 53520 1 1310
2 53521 1 1310
2 53522 1 1310
2 53523 1 1310
2 53524 1 1310
2 53525 1 1310
2 53526 1 1310
2 53527 1 1310
2 53528 1 1310
2 53529 1 1311
2 53530 1 1311
2 53531 1 1311
2 53532 1 1311
2 53533 1 1311
2 53534 1 1312
2 53535 1 1312
2 53536 1 1312
2 53537 1 1313
2 53538 1 1313
2 53539 1 1313
2 53540 1 1313
2 53541 1 1313
2 53542 1 1313
2 53543 1 1313
2 53544 1 1315
2 53545 1 1315
2 53546 1 1315
2 53547 1 1315
2 53548 1 1315
2 53549 1 1315
2 53550 1 1315
2 53551 1 1321
2 53552 1 1321
2 53553 1 1321
2 53554 1 1321
2 53555 1 1322
2 53556 1 1322
2 53557 1 1322
2 53558 1 1322
2 53559 1 1322
2 53560 1 1322
2 53561 1 1322
2 53562 1 1324
2 53563 1 1324
2 53564 1 1324
2 53565 1 1324
2 53566 1 1325
2 53567 1 1325
2 53568 1 1325
2 53569 1 1325
2 53570 1 1325
2 53571 1 1325
2 53572 1 1325
2 53573 1 1325
2 53574 1 1325
2 53575 1 1325
2 53576 1 1325
2 53577 1 1325
2 53578 1 1325
2 53579 1 1325
2 53580 1 1325
2 53581 1 1325
2 53582 1 1325
2 53583 1 1325
2 53584 1 1325
2 53585 1 1325
2 53586 1 1325
2 53587 1 1325
2 53588 1 1325
2 53589 1 1325
2 53590 1 1325
2 53591 1 1325
2 53592 1 1325
2 53593 1 1325
2 53594 1 1325
2 53595 1 1325
2 53596 1 1325
2 53597 1 1325
2 53598 1 1325
2 53599 1 1325
2 53600 1 1325
2 53601 1 1325
2 53602 1 1325
2 53603 1 1325
2 53604 1 1325
2 53605 1 1325
2 53606 1 1325
2 53607 1 1325
2 53608 1 1325
2 53609 1 1325
2 53610 1 1325
2 53611 1 1325
2 53612 1 1325
2 53613 1 1325
2 53614 1 1325
2 53615 1 1325
2 53616 1 1325
2 53617 1 1325
2 53618 1 1325
2 53619 1 1325
2 53620 1 1325
2 53621 1 1325
2 53622 1 1326
2 53623 1 1326
2 53624 1 1336
2 53625 1 1336
2 53626 1 1336
2 53627 1 1336
2 53628 1 1336
2 53629 1 1336
2 53630 1 1336
2 53631 1 1336
2 53632 1 1336
2 53633 1 1336
2 53634 1 1336
2 53635 1 1336
2 53636 1 1336
2 53637 1 1337
2 53638 1 1337
2 53639 1 1337
2 53640 1 1337
2 53641 1 1339
2 53642 1 1339
2 53643 1 1339
2 53644 1 1339
2 53645 1 1339
2 53646 1 1339
2 53647 1 1339
2 53648 1 1339
2 53649 1 1339
2 53650 1 1339
2 53651 1 1339
2 53652 1 1339
2 53653 1 1339
2 53654 1 1339
2 53655 1 1339
2 53656 1 1339
2 53657 1 1339
2 53658 1 1339
2 53659 1 1339
2 53660 1 1339
2 53661 1 1340
2 53662 1 1340
2 53663 1 1343
2 53664 1 1343
2 53665 1 1343
2 53666 1 1343
2 53667 1 1343
2 53668 1 1343
2 53669 1 1343
2 53670 1 1343
2 53671 1 1343
2 53672 1 1343
2 53673 1 1343
2 53674 1 1343
2 53675 1 1343
2 53676 1 1343
2 53677 1 1343
2 53678 1 1343
2 53679 1 1343
2 53680 1 1343
2 53681 1 1346
2 53682 1 1346
2 53683 1 1346
2 53684 1 1346
2 53685 1 1346
2 53686 1 1346
2 53687 1 1346
2 53688 1 1346
2 53689 1 1346
2 53690 1 1347
2 53691 1 1347
2 53692 1 1347
2 53693 1 1347
2 53694 1 1347
2 53695 1 1348
2 53696 1 1348
2 53697 1 1348
2 53698 1 1351
2 53699 1 1351
2 53700 1 1351
2 53701 1 1351
2 53702 1 1351
2 53703 1 1351
2 53704 1 1351
2 53705 1 1351
2 53706 1 1351
2 53707 1 1351
2 53708 1 1351
2 53709 1 1351
2 53710 1 1351
2 53711 1 1351
2 53712 1 1351
2 53713 1 1351
2 53714 1 1351
2 53715 1 1352
2 53716 1 1352
2 53717 1 1352
2 53718 1 1352
2 53719 1 1352
2 53720 1 1352
2 53721 1 1352
2 53722 1 1353
2 53723 1 1353
2 53724 1 1353
2 53725 1 1353
2 53726 1 1353
2 53727 1 1353
2 53728 1 1353
2 53729 1 1353
2 53730 1 1353
2 53731 1 1353
2 53732 1 1353
2 53733 1 1353
2 53734 1 1356
2 53735 1 1356
2 53736 1 1356
2 53737 1 1356
2 53738 1 1356
2 53739 1 1356
2 53740 1 1356
2 53741 1 1356
2 53742 1 1356
2 53743 1 1356
2 53744 1 1356
2 53745 1 1356
2 53746 1 1356
2 53747 1 1356
2 53748 1 1357
2 53749 1 1357
2 53750 1 1357
2 53751 1 1357
2 53752 1 1357
2 53753 1 1357
2 53754 1 1357
2 53755 1 1357
2 53756 1 1357
2 53757 1 1357
2 53758 1 1357
2 53759 1 1357
2 53760 1 1358
2 53761 1 1358
2 53762 1 1358
2 53763 1 1358
2 53764 1 1358
2 53765 1 1359
2 53766 1 1359
2 53767 1 1359
2 53768 1 1359
2 53769 1 1359
2 53770 1 1359
2 53771 1 1363
2 53772 1 1363
2 53773 1 1363
2 53774 1 1363
2 53775 1 1363
2 53776 1 1363
2 53777 1 1363
2 53778 1 1364
2 53779 1 1364
2 53780 1 1364
2 53781 1 1372
2 53782 1 1372
2 53783 1 1372
2 53784 1 1372
2 53785 1 1372
2 53786 1 1380
2 53787 1 1380
2 53788 1 1381
2 53789 1 1381
2 53790 1 1381
2 53791 1 1382
2 53792 1 1382
2 53793 1 1382
2 53794 1 1382
2 53795 1 1382
2 53796 1 1382
2 53797 1 1382
2 53798 1 1382
2 53799 1 1389
2 53800 1 1389
2 53801 1 1389
2 53802 1 1389
2 53803 1 1389
2 53804 1 1389
2 53805 1 1389
2 53806 1 1389
2 53807 1 1389
2 53808 1 1389
2 53809 1 1389
2 53810 1 1389
2 53811 1 1389
2 53812 1 1389
2 53813 1 1391
2 53814 1 1391
2 53815 1 1391
2 53816 1 1392
2 53817 1 1392
2 53818 1 1393
2 53819 1 1393
2 53820 1 1394
2 53821 1 1394
2 53822 1 1394
2 53823 1 1394
2 53824 1 1394
2 53825 1 1394
2 53826 1 1394
2 53827 1 1397
2 53828 1 1397
2 53829 1 1397
2 53830 1 1397
2 53831 1 1400
2 53832 1 1400
2 53833 1 1400
2 53834 1 1400
2 53835 1 1400
2 53836 1 1400
2 53837 1 1400
2 53838 1 1403
2 53839 1 1403
2 53840 1 1403
2 53841 1 1405
2 53842 1 1405
2 53843 1 1406
2 53844 1 1406
2 53845 1 1417
2 53846 1 1417
2 53847 1 1417
2 53848 1 1417
2 53849 1 1417
2 53850 1 1417
2 53851 1 1417
2 53852 1 1417
2 53853 1 1417
2 53854 1 1417
2 53855 1 1417
2 53856 1 1417
2 53857 1 1417
2 53858 1 1417
2 53859 1 1417
2 53860 1 1417
2 53861 1 1417
2 53862 1 1417
2 53863 1 1419
2 53864 1 1419
2 53865 1 1419
2 53866 1 1419
2 53867 1 1422
2 53868 1 1422
2 53869 1 1423
2 53870 1 1423
2 53871 1 1431
2 53872 1 1431
2 53873 1 1431
2 53874 1 1431
2 53875 1 1432
2 53876 1 1432
2 53877 1 1434
2 53878 1 1434
2 53879 1 1435
2 53880 1 1435
2 53881 1 1440
2 53882 1 1440
2 53883 1 1440
2 53884 1 1440
2 53885 1 1440
2 53886 1 1440
2 53887 1 1440
2 53888 1 1440
2 53889 1 1440
2 53890 1 1440
2 53891 1 1441
2 53892 1 1441
2 53893 1 1450
2 53894 1 1450
2 53895 1 1450
2 53896 1 1452
2 53897 1 1452
2 53898 1 1452
2 53899 1 1452
2 53900 1 1452
2 53901 1 1452
2 53902 1 1452
2 53903 1 1455
2 53904 1 1455
2 53905 1 1455
2 53906 1 1455
2 53907 1 1455
2 53908 1 1455
2 53909 1 1455
2 53910 1 1455
2 53911 1 1455
2 53912 1 1455
2 53913 1 1455
2 53914 1 1455
2 53915 1 1455
2 53916 1 1455
2 53917 1 1455
2 53918 1 1455
2 53919 1 1455
2 53920 1 1455
2 53921 1 1455
2 53922 1 1455
2 53923 1 1456
2 53924 1 1456
2 53925 1 1456
2 53926 1 1456
2 53927 1 1458
2 53928 1 1458
2 53929 1 1459
2 53930 1 1459
2 53931 1 1459
2 53932 1 1459
2 53933 1 1459
2 53934 1 1459
2 53935 1 1459
2 53936 1 1459
2 53937 1 1459
2 53938 1 1459
2 53939 1 1459
2 53940 1 1459
2 53941 1 1459
2 53942 1 1460
2 53943 1 1460
2 53944 1 1460
2 53945 1 1460
2 53946 1 1460
2 53947 1 1460
2 53948 1 1460
2 53949 1 1461
2 53950 1 1461
2 53951 1 1461
2 53952 1 1461
2 53953 1 1462
2 53954 1 1462
2 53955 1 1466
2 53956 1 1466
2 53957 1 1466
2 53958 1 1467
2 53959 1 1467
2 53960 1 1468
2 53961 1 1468
2 53962 1 1468
2 53963 1 1468
2 53964 1 1468
2 53965 1 1468
2 53966 1 1468
2 53967 1 1468
2 53968 1 1468
2 53969 1 1468
2 53970 1 1468
2 53971 1 1468
2 53972 1 1468
2 53973 1 1469
2 53974 1 1469
2 53975 1 1469
2 53976 1 1478
2 53977 1 1478
2 53978 1 1481
2 53979 1 1481
2 53980 1 1487
2 53981 1 1487
2 53982 1 1487
2 53983 1 1487
2 53984 1 1487
2 53985 1 1487
2 53986 1 1487
2 53987 1 1487
2 53988 1 1489
2 53989 1 1489
2 53990 1 1489
2 53991 1 1489
2 53992 1 1489
2 53993 1 1489
2 53994 1 1489
2 53995 1 1489
2 53996 1 1489
2 53997 1 1489
2 53998 1 1489
2 53999 1 1489
2 54000 1 1489
2 54001 1 1489
2 54002 1 1489
2 54003 1 1489
2 54004 1 1489
2 54005 1 1489
2 54006 1 1489
2 54007 1 1491
2 54008 1 1491
2 54009 1 1501
2 54010 1 1501
2 54011 1 1501
2 54012 1 1504
2 54013 1 1504
2 54014 1 1504
2 54015 1 1504
2 54016 1 1504
2 54017 1 1504
2 54018 1 1504
2 54019 1 1504
2 54020 1 1504
2 54021 1 1504
2 54022 1 1504
2 54023 1 1504
2 54024 1 1504
2 54025 1 1505
2 54026 1 1505
2 54027 1 1505
2 54028 1 1505
2 54029 1 1505
2 54030 1 1505
2 54031 1 1505
2 54032 1 1505
2 54033 1 1505
2 54034 1 1505
2 54035 1 1505
2 54036 1 1505
2 54037 1 1505
2 54038 1 1505
2 54039 1 1505
2 54040 1 1505
2 54041 1 1505
2 54042 1 1510
2 54043 1 1510
2 54044 1 1510
2 54045 1 1512
2 54046 1 1512
2 54047 1 1513
2 54048 1 1513
2 54049 1 1516
2 54050 1 1516
2 54051 1 1516
2 54052 1 1516
2 54053 1 1516
2 54054 1 1516
2 54055 1 1516
2 54056 1 1516
2 54057 1 1516
2 54058 1 1516
2 54059 1 1516
2 54060 1 1516
2 54061 1 1516
2 54062 1 1516
2 54063 1 1516
2 54064 1 1516
2 54065 1 1516
2 54066 1 1516
2 54067 1 1517
2 54068 1 1517
2 54069 1 1517
2 54070 1 1527
2 54071 1 1527
2 54072 1 1527
2 54073 1 1527
2 54074 1 1527
2 54075 1 1527
2 54076 1 1527
2 54077 1 1527
2 54078 1 1527
2 54079 1 1529
2 54080 1 1529
2 54081 1 1529
2 54082 1 1529
2 54083 1 1529
2 54084 1 1529
2 54085 1 1529
2 54086 1 1529
2 54087 1 1530
2 54088 1 1530
2 54089 1 1530
2 54090 1 1530
2 54091 1 1530
2 54092 1 1530
2 54093 1 1530
2 54094 1 1530
2 54095 1 1530
2 54096 1 1530
2 54097 1 1530
2 54098 1 1530
2 54099 1 1530
2 54100 1 1530
2 54101 1 1530
2 54102 1 1531
2 54103 1 1531
2 54104 1 1531
2 54105 1 1540
2 54106 1 1540
2 54107 1 1540
2 54108 1 1540
2 54109 1 1540
2 54110 1 1545
2 54111 1 1545
2 54112 1 1546
2 54113 1 1546
2 54114 1 1546
2 54115 1 1546
2 54116 1 1546
2 54117 1 1546
2 54118 1 1554
2 54119 1 1554
2 54120 1 1554
2 54121 1 1555
2 54122 1 1555
2 54123 1 1555
2 54124 1 1556
2 54125 1 1556
2 54126 1 1556
2 54127 1 1569
2 54128 1 1569
2 54129 1 1569
2 54130 1 1569
2 54131 1 1572
2 54132 1 1572
2 54133 1 1572
2 54134 1 1572
2 54135 1 1572
2 54136 1 1572
2 54137 1 1572
2 54138 1 1572
2 54139 1 1572
2 54140 1 1573
2 54141 1 1573
2 54142 1 1581
2 54143 1 1581
2 54144 1 1582
2 54145 1 1582
2 54146 1 1582
2 54147 1 1582
2 54148 1 1584
2 54149 1 1584
2 54150 1 1589
2 54151 1 1589
2 54152 1 1589
2 54153 1 1589
2 54154 1 1589
2 54155 1 1589
2 54156 1 1589
2 54157 1 1589
2 54158 1 1589
2 54159 1 1589
2 54160 1 1589
2 54161 1 1589
2 54162 1 1589
2 54163 1 1589
2 54164 1 1589
2 54165 1 1589
2 54166 1 1591
2 54167 1 1591
2 54168 1 1591
2 54169 1 1593
2 54170 1 1593
2 54171 1 1609
2 54172 1 1609
2 54173 1 1609
2 54174 1 1609
2 54175 1 1609
2 54176 1 1609
2 54177 1 1612
2 54178 1 1612
2 54179 1 1613
2 54180 1 1613
2 54181 1 1613
2 54182 1 1613
2 54183 1 1613
2 54184 1 1613
2 54185 1 1613
2 54186 1 1613
2 54187 1 1613
2 54188 1 1615
2 54189 1 1615
2 54190 1 1620
2 54191 1 1620
2 54192 1 1620
2 54193 1 1621
2 54194 1 1621
2 54195 1 1623
2 54196 1 1623
2 54197 1 1623
2 54198 1 1624
2 54199 1 1624
2 54200 1 1624
2 54201 1 1626
2 54202 1 1626
2 54203 1 1626
2 54204 1 1626
2 54205 1 1626
2 54206 1 1626
2 54207 1 1626
2 54208 1 1626
2 54209 1 1626
2 54210 1 1626
2 54211 1 1626
2 54212 1 1626
2 54213 1 1626
2 54214 1 1626
2 54215 1 1626
2 54216 1 1626
2 54217 1 1626
2 54218 1 1626
2 54219 1 1626
2 54220 1 1626
2 54221 1 1626
2 54222 1 1626
2 54223 1 1626
2 54224 1 1626
2 54225 1 1626
2 54226 1 1626
2 54227 1 1627
2 54228 1 1627
2 54229 1 1627
2 54230 1 1627
2 54231 1 1627
2 54232 1 1627
2 54233 1 1627
2 54234 1 1627
2 54235 1 1627
2 54236 1 1627
2 54237 1 1627
2 54238 1 1627
2 54239 1 1627
2 54240 1 1628
2 54241 1 1628
2 54242 1 1628
2 54243 1 1628
2 54244 1 1628
2 54245 1 1628
2 54246 1 1628
2 54247 1 1628
2 54248 1 1628
2 54249 1 1628
2 54250 1 1633
2 54251 1 1633
2 54252 1 1633
2 54253 1 1634
2 54254 1 1634
2 54255 1 1634
2 54256 1 1634
2 54257 1 1634
2 54258 1 1634
2 54259 1 1634
2 54260 1 1634
2 54261 1 1634
2 54262 1 1634
2 54263 1 1634
2 54264 1 1634
2 54265 1 1634
2 54266 1 1634
2 54267 1 1634
2 54268 1 1634
2 54269 1 1634
2 54270 1 1634
2 54271 1 1634
2 54272 1 1634
2 54273 1 1634
2 54274 1 1634
2 54275 1 1634
2 54276 1 1634
2 54277 1 1634
2 54278 1 1634
2 54279 1 1634
2 54280 1 1634
2 54281 1 1634
2 54282 1 1634
2 54283 1 1634
2 54284 1 1634
2 54285 1 1634
2 54286 1 1634
2 54287 1 1634
2 54288 1 1634
2 54289 1 1634
2 54290 1 1635
2 54291 1 1635
2 54292 1 1635
2 54293 1 1635
2 54294 1 1635
2 54295 1 1648
2 54296 1 1648
2 54297 1 1648
2 54298 1 1648
2 54299 1 1649
2 54300 1 1649
2 54301 1 1649
2 54302 1 1650
2 54303 1 1650
2 54304 1 1650
2 54305 1 1650
2 54306 1 1650
2 54307 1 1650
2 54308 1 1650
2 54309 1 1650
2 54310 1 1650
2 54311 1 1650
2 54312 1 1650
2 54313 1 1650
2 54314 1 1650
2 54315 1 1650
2 54316 1 1650
2 54317 1 1650
2 54318 1 1658
2 54319 1 1658
2 54320 1 1658
2 54321 1 1658
2 54322 1 1671
2 54323 1 1671
2 54324 1 1671
2 54325 1 1671
2 54326 1 1671
2 54327 1 1671
2 54328 1 1671
2 54329 1 1671
2 54330 1 1671
2 54331 1 1673
2 54332 1 1673
2 54333 1 1676
2 54334 1 1676
2 54335 1 1678
2 54336 1 1678
2 54337 1 1678
2 54338 1 1678
2 54339 1 1678
2 54340 1 1678
2 54341 1 1679
2 54342 1 1679
2 54343 1 1686
2 54344 1 1686
2 54345 1 1686
2 54346 1 1687
2 54347 1 1687
2 54348 1 1687
2 54349 1 1687
2 54350 1 1687
2 54351 1 1687
2 54352 1 1695
2 54353 1 1695
2 54354 1 1697
2 54355 1 1697
2 54356 1 1697
2 54357 1 1697
2 54358 1 1697
2 54359 1 1698
2 54360 1 1698
2 54361 1 1698
2 54362 1 1698
2 54363 1 1701
2 54364 1 1701
2 54365 1 1706
2 54366 1 1706
2 54367 1 1706
2 54368 1 1706
2 54369 1 1706
2 54370 1 1706
2 54371 1 1706
2 54372 1 1706
2 54373 1 1706
2 54374 1 1706
2 54375 1 1706
2 54376 1 1706
2 54377 1 1706
2 54378 1 1706
2 54379 1 1706
2 54380 1 1706
2 54381 1 1706
2 54382 1 1706
2 54383 1 1706
2 54384 1 1706
2 54385 1 1706
2 54386 1 1706
2 54387 1 1706
2 54388 1 1706
2 54389 1 1706
2 54390 1 1706
2 54391 1 1706
2 54392 1 1706
2 54393 1 1706
2 54394 1 1708
2 54395 1 1708
2 54396 1 1708
2 54397 1 1708
2 54398 1 1708
2 54399 1 1718
2 54400 1 1718
2 54401 1 1718
2 54402 1 1718
2 54403 1 1721
2 54404 1 1721
2 54405 1 1721
2 54406 1 1722
2 54407 1 1722
2 54408 1 1722
2 54409 1 1734
2 54410 1 1734
2 54411 1 1734
2 54412 1 1734
2 54413 1 1734
2 54414 1 1734
2 54415 1 1734
2 54416 1 1734
2 54417 1 1734
2 54418 1 1735
2 54419 1 1735
2 54420 1 1735
2 54421 1 1735
2 54422 1 1735
2 54423 1 1735
2 54424 1 1735
2 54425 1 1735
2 54426 1 1735
2 54427 1 1735
2 54428 1 1735
2 54429 1 1735
2 54430 1 1737
2 54431 1 1737
2 54432 1 1737
2 54433 1 1737
2 54434 1 1737
2 54435 1 1737
2 54436 1 1737
2 54437 1 1738
2 54438 1 1738
2 54439 1 1738
2 54440 1 1738
2 54441 1 1738
2 54442 1 1738
2 54443 1 1738
2 54444 1 1738
2 54445 1 1740
2 54446 1 1740
2 54447 1 1741
2 54448 1 1741
2 54449 1 1741
2 54450 1 1741
2 54451 1 1741
2 54452 1 1741
2 54453 1 1741
2 54454 1 1742
2 54455 1 1742
2 54456 1 1742
2 54457 1 1749
2 54458 1 1749
2 54459 1 1749
2 54460 1 1749
2 54461 1 1749
2 54462 1 1749
2 54463 1 1749
2 54464 1 1749
2 54465 1 1749
2 54466 1 1749
2 54467 1 1750
2 54468 1 1750
2 54469 1 1750
2 54470 1 1750
2 54471 1 1752
2 54472 1 1752
2 54473 1 1755
2 54474 1 1755
2 54475 1 1763
2 54476 1 1763
2 54477 1 1763
2 54478 1 1763
2 54479 1 1763
2 54480 1 1763
2 54481 1 1763
2 54482 1 1763
2 54483 1 1763
2 54484 1 1763
2 54485 1 1763
2 54486 1 1765
2 54487 1 1765
2 54488 1 1765
2 54489 1 1766
2 54490 1 1766
2 54491 1 1771
2 54492 1 1771
2 54493 1 1775
2 54494 1 1775
2 54495 1 1775
2 54496 1 1775
2 54497 1 1775
2 54498 1 1775
2 54499 1 1775
2 54500 1 1775
2 54501 1 1775
2 54502 1 1775
2 54503 1 1775
2 54504 1 1775
2 54505 1 1775
2 54506 1 1775
2 54507 1 1775
2 54508 1 1775
2 54509 1 1775
2 54510 1 1775
2 54511 1 1775
2 54512 1 1776
2 54513 1 1776
2 54514 1 1776
2 54515 1 1776
2 54516 1 1776
2 54517 1 1776
2 54518 1 1776
2 54519 1 1777
2 54520 1 1777
2 54521 1 1791
2 54522 1 1791
2 54523 1 1791
2 54524 1 1791
2 54525 1 1791
2 54526 1 1793
2 54527 1 1793
2 54528 1 1793
2 54529 1 1793
2 54530 1 1793
2 54531 1 1793
2 54532 1 1793
2 54533 1 1793
2 54534 1 1793
2 54535 1 1793
2 54536 1 1793
2 54537 1 1793
2 54538 1 1795
2 54539 1 1795
2 54540 1 1795
2 54541 1 1796
2 54542 1 1796
2 54543 1 1796
2 54544 1 1799
2 54545 1 1799
2 54546 1 1799
2 54547 1 1799
2 54548 1 1799
2 54549 1 1800
2 54550 1 1800
2 54551 1 1803
2 54552 1 1803
2 54553 1 1803
2 54554 1 1803
2 54555 1 1803
2 54556 1 1805
2 54557 1 1805
2 54558 1 1805
2 54559 1 1808
2 54560 1 1808
2 54561 1 1808
2 54562 1 1808
2 54563 1 1808
2 54564 1 1808
2 54565 1 1808
2 54566 1 1808
2 54567 1 1808
2 54568 1 1808
2 54569 1 1809
2 54570 1 1809
2 54571 1 1809
2 54572 1 1809
2 54573 1 1809
2 54574 1 1809
2 54575 1 1809
2 54576 1 1809
2 54577 1 1810
2 54578 1 1810
2 54579 1 1818
2 54580 1 1818
2 54581 1 1834
2 54582 1 1834
2 54583 1 1839
2 54584 1 1839
2 54585 1 1839
2 54586 1 1842
2 54587 1 1842
2 54588 1 1842
2 54589 1 1842
2 54590 1 1843
2 54591 1 1843
2 54592 1 1843
2 54593 1 1843
2 54594 1 1843
2 54595 1 1850
2 54596 1 1850
2 54597 1 1850
2 54598 1 1850
2 54599 1 1850
2 54600 1 1850
2 54601 1 1850
2 54602 1 1850
2 54603 1 1850
2 54604 1 1859
2 54605 1 1859
2 54606 1 1859
2 54607 1 1860
2 54608 1 1860
2 54609 1 1860
2 54610 1 1862
2 54611 1 1862
2 54612 1 1862
2 54613 1 1862
2 54614 1 1862
2 54615 1 1862
2 54616 1 1862
2 54617 1 1873
2 54618 1 1873
2 54619 1 1873
2 54620 1 1873
2 54621 1 1873
2 54622 1 1873
2 54623 1 1873
2 54624 1 1873
2 54625 1 1873
2 54626 1 1873
2 54627 1 1873
2 54628 1 1884
2 54629 1 1884
2 54630 1 1891
2 54631 1 1891
2 54632 1 1891
2 54633 1 1893
2 54634 1 1893
2 54635 1 1900
2 54636 1 1900
2 54637 1 1900
2 54638 1 1900
2 54639 1 1901
2 54640 1 1901
2 54641 1 1902
2 54642 1 1902
2 54643 1 1902
2 54644 1 1902
2 54645 1 1902
2 54646 1 1902
2 54647 1 1902
2 54648 1 1904
2 54649 1 1904
2 54650 1 1905
2 54651 1 1905
2 54652 1 1905
2 54653 1 1909
2 54654 1 1909
2 54655 1 1909
2 54656 1 1909
2 54657 1 1909
2 54658 1 1909
2 54659 1 1909
2 54660 1 1910
2 54661 1 1910
2 54662 1 1910
2 54663 1 1911
2 54664 1 1911
2 54665 1 1911
2 54666 1 1911
2 54667 1 1911
2 54668 1 1935
2 54669 1 1935
2 54670 1 1936
2 54671 1 1936
2 54672 1 1938
2 54673 1 1938
2 54674 1 1941
2 54675 1 1941
2 54676 1 1941
2 54677 1 1941
2 54678 1 1941
2 54679 1 1941
2 54680 1 1941
2 54681 1 1942
2 54682 1 1942
2 54683 1 1943
2 54684 1 1943
2 54685 1 1943
2 54686 1 1949
2 54687 1 1949
2 54688 1 1949
2 54689 1 1953
2 54690 1 1953
2 54691 1 1955
2 54692 1 1955
2 54693 1 1962
2 54694 1 1962
2 54695 1 1962
2 54696 1 1962
2 54697 1 1962
2 54698 1 1962
2 54699 1 1962
2 54700 1 1962
2 54701 1 1962
2 54702 1 1962
2 54703 1 1963
2 54704 1 1963
2 54705 1 1963
2 54706 1 1963
2 54707 1 1971
2 54708 1 1971
2 54709 1 1972
2 54710 1 1972
2 54711 1 1973
2 54712 1 1973
2 54713 1 1973
2 54714 1 1973
2 54715 1 1973
2 54716 1 1973
2 54717 1 1973
2 54718 1 1974
2 54719 1 1974
2 54720 1 1977
2 54721 1 1977
2 54722 1 1977
2 54723 1 1977
2 54724 1 1977
2 54725 1 1977
2 54726 1 1977
2 54727 1 1977
2 54728 1 1977
2 54729 1 1977
2 54730 1 1977
2 54731 1 1978
2 54732 1 1978
2 54733 1 1978
2 54734 1 1978
2 54735 1 1978
2 54736 1 1978
2 54737 1 1979
2 54738 1 1979
2 54739 1 1985
2 54740 1 1985
2 54741 1 1985
2 54742 1 1985
2 54743 1 1985
2 54744 1 1985
2 54745 1 1985
2 54746 1 1985
2 54747 1 1985
2 54748 1 1985
2 54749 1 1987
2 54750 1 1987
2 54751 1 1988
2 54752 1 1988
2 54753 1 1988
2 54754 1 1988
2 54755 1 1988
2 54756 1 1988
2 54757 1 1988
2 54758 1 1988
2 54759 1 1988
2 54760 1 1988
2 54761 1 1988
2 54762 1 1988
2 54763 1 1988
2 54764 1 1988
2 54765 1 1988
2 54766 1 1988
2 54767 1 1988
2 54768 1 1988
2 54769 1 1988
2 54770 1 1988
2 54771 1 1988
2 54772 1 1988
2 54773 1 1988
2 54774 1 1988
2 54775 1 1988
2 54776 1 1988
2 54777 1 1988
2 54778 1 1988
2 54779 1 1988
2 54780 1 1988
2 54781 1 1988
2 54782 1 1988
2 54783 1 1988
2 54784 1 1988
2 54785 1 1988
2 54786 1 1988
2 54787 1 1988
2 54788 1 1988
2 54789 1 1988
2 54790 1 1988
2 54791 1 1988
2 54792 1 1988
2 54793 1 1988
2 54794 1 1988
2 54795 1 1988
2 54796 1 1988
2 54797 1 1988
2 54798 1 1988
2 54799 1 1988
2 54800 1 1988
2 54801 1 1988
2 54802 1 1988
2 54803 1 1988
2 54804 1 1988
2 54805 1 1988
2 54806 1 1988
2 54807 1 1988
2 54808 1 1988
2 54809 1 1988
2 54810 1 1988
2 54811 1 1988
2 54812 1 1988
2 54813 1 1988
2 54814 1 1988
2 54815 1 1988
2 54816 1 1988
2 54817 1 1989
2 54818 1 1989
2 54819 1 1989
2 54820 1 2001
2 54821 1 2001
2 54822 1 2004
2 54823 1 2004
2 54824 1 2004
2 54825 1 2004
2 54826 1 2004
2 54827 1 2004
2 54828 1 2004
2 54829 1 2004
2 54830 1 2004
2 54831 1 2004
2 54832 1 2004
2 54833 1 2004
2 54834 1 2004
2 54835 1 2004
2 54836 1 2013
2 54837 1 2013
2 54838 1 2013
2 54839 1 2013
2 54840 1 2013
2 54841 1 2013
2 54842 1 2013
2 54843 1 2013
2 54844 1 2013
2 54845 1 2013
2 54846 1 2013
2 54847 1 2013
2 54848 1 2013
2 54849 1 2013
2 54850 1 2013
2 54851 1 2013
2 54852 1 2013
2 54853 1 2013
2 54854 1 2013
2 54855 1 2013
2 54856 1 2015
2 54857 1 2015
2 54858 1 2015
2 54859 1 2022
2 54860 1 2022
2 54861 1 2022
2 54862 1 2022
2 54863 1 2022
2 54864 1 2023
2 54865 1 2023
2 54866 1 2023
2 54867 1 2023
2 54868 1 2023
2 54869 1 2025
2 54870 1 2025
2 54871 1 2025
2 54872 1 2025
2 54873 1 2025
2 54874 1 2025
2 54875 1 2025
2 54876 1 2025
2 54877 1 2028
2 54878 1 2028
2 54879 1 2028
2 54880 1 2028
2 54881 1 2029
2 54882 1 2029
2 54883 1 2029
2 54884 1 2040
2 54885 1 2040
2 54886 1 2043
2 54887 1 2043
2 54888 1 2043
2 54889 1 2043
2 54890 1 2044
2 54891 1 2044
2 54892 1 2044
2 54893 1 2044
2 54894 1 2044
2 54895 1 2044
2 54896 1 2044
2 54897 1 2044
2 54898 1 2044
2 54899 1 2044
2 54900 1 2044
2 54901 1 2044
2 54902 1 2044
2 54903 1 2045
2 54904 1 2045
2 54905 1 2045
2 54906 1 2045
2 54907 1 2045
2 54908 1 2045
2 54909 1 2045
2 54910 1 2058
2 54911 1 2058
2 54912 1 2058
2 54913 1 2058
2 54914 1 2058
2 54915 1 2058
2 54916 1 2058
2 54917 1 2058
2 54918 1 2058
2 54919 1 2063
2 54920 1 2063
2 54921 1 2063
2 54922 1 2063
2 54923 1 2066
2 54924 1 2066
2 54925 1 2066
2 54926 1 2066
2 54927 1 2066
2 54928 1 2066
2 54929 1 2066
2 54930 1 2066
2 54931 1 2066
2 54932 1 2066
2 54933 1 2066
2 54934 1 2066
2 54935 1 2066
2 54936 1 2066
2 54937 1 2066
2 54938 1 2066
2 54939 1 2066
2 54940 1 2066
2 54941 1 2066
2 54942 1 2067
2 54943 1 2067
2 54944 1 2067
2 54945 1 2067
2 54946 1 2067
2 54947 1 2067
2 54948 1 2067
2 54949 1 2067
2 54950 1 2067
2 54951 1 2067
2 54952 1 2067
2 54953 1 2067
2 54954 1 2067
2 54955 1 2067
2 54956 1 2067
2 54957 1 2067
2 54958 1 2067
2 54959 1 2067
2 54960 1 2067
2 54961 1 2067
2 54962 1 2067
2 54963 1 2067
2 54964 1 2067
2 54965 1 2067
2 54966 1 2067
2 54967 1 2067
2 54968 1 2067
2 54969 1 2067
2 54970 1 2067
2 54971 1 2067
2 54972 1 2067
2 54973 1 2067
2 54974 1 2067
2 54975 1 2067
2 54976 1 2067
2 54977 1 2067
2 54978 1 2067
2 54979 1 2067
2 54980 1 2067
2 54981 1 2067
2 54982 1 2068
2 54983 1 2068
2 54984 1 2068
2 54985 1 2068
2 54986 1 2068
2 54987 1 2068
2 54988 1 2068
2 54989 1 2068
2 54990 1 2068
2 54991 1 2069
2 54992 1 2069
2 54993 1 2069
2 54994 1 2070
2 54995 1 2070
2 54996 1 2076
2 54997 1 2076
2 54998 1 2083
2 54999 1 2083
2 55000 1 2083
2 55001 1 2083
2 55002 1 2083
2 55003 1 2083
2 55004 1 2083
2 55005 1 2083
2 55006 1 2083
2 55007 1 2084
2 55008 1 2084
2 55009 1 2084
2 55010 1 2091
2 55011 1 2091
2 55012 1 2091
2 55013 1 2091
2 55014 1 2100
2 55015 1 2100
2 55016 1 2100
2 55017 1 2100
2 55018 1 2100
2 55019 1 2100
2 55020 1 2102
2 55021 1 2102
2 55022 1 2102
2 55023 1 2102
2 55024 1 2102
2 55025 1 2102
2 55026 1 2103
2 55027 1 2103
2 55028 1 2103
2 55029 1 2105
2 55030 1 2105
2 55031 1 2105
2 55032 1 2114
2 55033 1 2114
2 55034 1 2114
2 55035 1 2114
2 55036 1 2114
2 55037 1 2114
2 55038 1 2114
2 55039 1 2114
2 55040 1 2126
2 55041 1 2126
2 55042 1 2126
2 55043 1 2126
2 55044 1 2126
2 55045 1 2139
2 55046 1 2139
2 55047 1 2139
2 55048 1 2142
2 55049 1 2142
2 55050 1 2143
2 55051 1 2143
2 55052 1 2154
2 55053 1 2154
2 55054 1 2154
2 55055 1 2154
2 55056 1 2154
2 55057 1 2160
2 55058 1 2160
2 55059 1 2160
2 55060 1 2160
2 55061 1 2161
2 55062 1 2161
2 55063 1 2162
2 55064 1 2162
2 55065 1 2162
2 55066 1 2162
2 55067 1 2162
2 55068 1 2162
2 55069 1 2162
2 55070 1 2162
2 55071 1 2162
2 55072 1 2162
2 55073 1 2163
2 55074 1 2163
2 55075 1 2163
2 55076 1 2165
2 55077 1 2165
2 55078 1 2165
2 55079 1 2165
2 55080 1 2165
2 55081 1 2165
2 55082 1 2166
2 55083 1 2166
2 55084 1 2168
2 55085 1 2168
2 55086 1 2168
2 55087 1 2171
2 55088 1 2171
2 55089 1 2171
2 55090 1 2178
2 55091 1 2178
2 55092 1 2181
2 55093 1 2181
2 55094 1 2181
2 55095 1 2181
2 55096 1 2181
2 55097 1 2181
2 55098 1 2181
2 55099 1 2181
2 55100 1 2181
2 55101 1 2181
2 55102 1 2181
2 55103 1 2181
2 55104 1 2181
2 55105 1 2181
2 55106 1 2181
2 55107 1 2181
2 55108 1 2181
2 55109 1 2181
2 55110 1 2183
2 55111 1 2183
2 55112 1 2183
2 55113 1 2183
2 55114 1 2185
2 55115 1 2185
2 55116 1 2186
2 55117 1 2186
2 55118 1 2201
2 55119 1 2201
2 55120 1 2201
2 55121 1 2201
2 55122 1 2202
2 55123 1 2202
2 55124 1 2202
2 55125 1 2204
2 55126 1 2204
2 55127 1 2204
2 55128 1 2204
2 55129 1 2204
2 55130 1 2204
2 55131 1 2204
2 55132 1 2205
2 55133 1 2205
2 55134 1 2205
2 55135 1 2210
2 55136 1 2210
2 55137 1 2210
2 55138 1 2210
2 55139 1 2210
2 55140 1 2210
2 55141 1 2210
2 55142 1 2210
2 55143 1 2211
2 55144 1 2211
2 55145 1 2211
2 55146 1 2211
2 55147 1 2211
2 55148 1 2211
2 55149 1 2211
2 55150 1 2211
2 55151 1 2211
2 55152 1 2211
2 55153 1 2211
2 55154 1 2212
2 55155 1 2212
2 55156 1 2212
2 55157 1 2212
2 55158 1 2212
2 55159 1 2212
2 55160 1 2212
2 55161 1 2212
2 55162 1 2212
2 55163 1 2212
2 55164 1 2213
2 55165 1 2213
2 55166 1 2213
2 55167 1 2213
2 55168 1 2213
2 55169 1 2222
2 55170 1 2222
2 55171 1 2222
2 55172 1 2222
2 55173 1 2223
2 55174 1 2223
2 55175 1 2224
2 55176 1 2224
2 55177 1 2225
2 55178 1 2225
2 55179 1 2226
2 55180 1 2226
2 55181 1 2226
2 55182 1 2226
2 55183 1 2226
2 55184 1 2226
2 55185 1 2226
2 55186 1 2226
2 55187 1 2226
2 55188 1 2226
2 55189 1 2226
2 55190 1 2226
2 55191 1 2226
2 55192 1 2226
2 55193 1 2226
2 55194 1 2226
2 55195 1 2230
2 55196 1 2230
2 55197 1 2230
2 55198 1 2230
2 55199 1 2230
2 55200 1 2230
2 55201 1 2230
2 55202 1 2230
2 55203 1 2230
2 55204 1 2231
2 55205 1 2231
2 55206 1 2232
2 55207 1 2232
2 55208 1 2232
2 55209 1 2237
2 55210 1 2237
2 55211 1 2238
2 55212 1 2238
2 55213 1 2239
2 55214 1 2239
2 55215 1 2239
2 55216 1 2239
2 55217 1 2239
2 55218 1 2239
2 55219 1 2239
2 55220 1 2239
2 55221 1 2239
2 55222 1 2239
2 55223 1 2239
2 55224 1 2239
2 55225 1 2248
2 55226 1 2248
2 55227 1 2248
2 55228 1 2248
2 55229 1 2248
2 55230 1 2248
2 55231 1 2248
2 55232 1 2248
2 55233 1 2248
2 55234 1 2248
2 55235 1 2252
2 55236 1 2252
2 55237 1 2256
2 55238 1 2256
2 55239 1 2256
2 55240 1 2256
2 55241 1 2268
2 55242 1 2268
2 55243 1 2280
2 55244 1 2280
2 55245 1 2285
2 55246 1 2285
2 55247 1 2287
2 55248 1 2287
2 55249 1 2287
2 55250 1 2287
2 55251 1 2287
2 55252 1 2287
2 55253 1 2288
2 55254 1 2288
2 55255 1 2288
2 55256 1 2289
2 55257 1 2289
2 55258 1 2289
2 55259 1 2289
2 55260 1 2296
2 55261 1 2296
2 55262 1 2296
2 55263 1 2296
2 55264 1 2296
2 55265 1 2296
2 55266 1 2298
2 55267 1 2298
2 55268 1 2298
2 55269 1 2298
2 55270 1 2298
2 55271 1 2314
2 55272 1 2314
2 55273 1 2314
2 55274 1 2315
2 55275 1 2315
2 55276 1 2315
2 55277 1 2315
2 55278 1 2315
2 55279 1 2315
2 55280 1 2316
2 55281 1 2316
2 55282 1 2316
2 55283 1 2329
2 55284 1 2329
2 55285 1 2329
2 55286 1 2329
2 55287 1 2329
2 55288 1 2329
2 55289 1 2329
2 55290 1 2329
2 55291 1 2329
2 55292 1 2341
2 55293 1 2341
2 55294 1 2342
2 55295 1 2342
2 55296 1 2342
2 55297 1 2342
2 55298 1 2342
2 55299 1 2343
2 55300 1 2343
2 55301 1 2344
2 55302 1 2344
2 55303 1 2344
2 55304 1 2344
2 55305 1 2345
2 55306 1 2345
2 55307 1 2351
2 55308 1 2351
2 55309 1 2357
2 55310 1 2357
2 55311 1 2357
2 55312 1 2365
2 55313 1 2365
2 55314 1 2365
2 55315 1 2365
2 55316 1 2365
2 55317 1 2365
2 55318 1 2365
2 55319 1 2366
2 55320 1 2366
2 55321 1 2366
2 55322 1 2366
2 55323 1 2366
2 55324 1 2366
2 55325 1 2366
2 55326 1 2366
2 55327 1 2366
2 55328 1 2366
2 55329 1 2366
2 55330 1 2370
2 55331 1 2370
2 55332 1 2375
2 55333 1 2375
2 55334 1 2375
2 55335 1 2383
2 55336 1 2383
2 55337 1 2394
2 55338 1 2394
2 55339 1 2394
2 55340 1 2394
2 55341 1 2394
2 55342 1 2394
2 55343 1 2394
2 55344 1 2394
2 55345 1 2394
2 55346 1 2395
2 55347 1 2395
2 55348 1 2395
2 55349 1 2397
2 55350 1 2397
2 55351 1 2398
2 55352 1 2398
2 55353 1 2401
2 55354 1 2401
2 55355 1 2401
2 55356 1 2404
2 55357 1 2404
2 55358 1 2413
2 55359 1 2413
2 55360 1 2413
2 55361 1 2413
2 55362 1 2414
2 55363 1 2414
2 55364 1 2414
2 55365 1 2415
2 55366 1 2415
2 55367 1 2416
2 55368 1 2416
2 55369 1 2440
2 55370 1 2440
2 55371 1 2440
2 55372 1 2440
2 55373 1 2440
2 55374 1 2440
2 55375 1 2440
2 55376 1 2440
2 55377 1 2440
2 55378 1 2440
2 55379 1 2440
2 55380 1 2440
2 55381 1 2440
2 55382 1 2440
2 55383 1 2440
2 55384 1 2440
2 55385 1 2440
2 55386 1 2440
2 55387 1 2440
2 55388 1 2440
2 55389 1 2440
2 55390 1 2445
2 55391 1 2445
2 55392 1 2445
2 55393 1 2446
2 55394 1 2446
2 55395 1 2454
2 55396 1 2454
2 55397 1 2454
2 55398 1 2454
2 55399 1 2454
2 55400 1 2454
2 55401 1 2454
2 55402 1 2454
2 55403 1 2454
2 55404 1 2455
2 55405 1 2455
2 55406 1 2470
2 55407 1 2470
2 55408 1 2470
2 55409 1 2470
2 55410 1 2470
2 55411 1 2470
2 55412 1 2470
2 55413 1 2470
2 55414 1 2471
2 55415 1 2471
2 55416 1 2472
2 55417 1 2472
2 55418 1 2472
2 55419 1 2472
2 55420 1 2472
2 55421 1 2472
2 55422 1 2472
2 55423 1 2472
2 55424 1 2472
2 55425 1 2472
2 55426 1 2472
2 55427 1 2472
2 55428 1 2472
2 55429 1 2472
2 55430 1 2472
2 55431 1 2473
2 55432 1 2473
2 55433 1 2473
2 55434 1 2473
2 55435 1 2482
2 55436 1 2482
2 55437 1 2482
2 55438 1 2482
2 55439 1 2482
2 55440 1 2483
2 55441 1 2483
2 55442 1 2483
2 55443 1 2483
2 55444 1 2483
2 55445 1 2483
2 55446 1 2483
2 55447 1 2484
2 55448 1 2484
2 55449 1 2484
2 55450 1 2485
2 55451 1 2485
2 55452 1 2490
2 55453 1 2490
2 55454 1 2490
2 55455 1 2490
2 55456 1 2490
2 55457 1 2490
2 55458 1 2490
2 55459 1 2490
2 55460 1 2490
2 55461 1 2490
2 55462 1 2490
2 55463 1 2490
2 55464 1 2490
2 55465 1 2490
2 55466 1 2491
2 55467 1 2491
2 55468 1 2491
2 55469 1 2492
2 55470 1 2492
2 55471 1 2492
2 55472 1 2492
2 55473 1 2492
2 55474 1 2492
2 55475 1 2492
2 55476 1 2492
2 55477 1 2492
2 55478 1 2492
2 55479 1 2492
2 55480 1 2493
2 55481 1 2493
2 55482 1 2494
2 55483 1 2494
2 55484 1 2494
2 55485 1 2494
2 55486 1 2495
2 55487 1 2495
2 55488 1 2495
2 55489 1 2495
2 55490 1 2495
2 55491 1 2495
2 55492 1 2495
2 55493 1 2495
2 55494 1 2495
2 55495 1 2495
2 55496 1 2504
2 55497 1 2504
2 55498 1 2504
2 55499 1 2504
2 55500 1 2504
2 55501 1 2504
2 55502 1 2504
2 55503 1 2505
2 55504 1 2505
2 55505 1 2507
2 55506 1 2507
2 55507 1 2507
2 55508 1 2507
2 55509 1 2534
2 55510 1 2534
2 55511 1 2535
2 55512 1 2535
2 55513 1 2535
2 55514 1 2535
2 55515 1 2536
2 55516 1 2536
2 55517 1 2537
2 55518 1 2537
2 55519 1 2537
2 55520 1 2537
2 55521 1 2537
2 55522 1 2537
2 55523 1 2537
2 55524 1 2537
2 55525 1 2537
2 55526 1 2537
2 55527 1 2537
2 55528 1 2537
2 55529 1 2538
2 55530 1 2538
2 55531 1 2539
2 55532 1 2539
2 55533 1 2539
2 55534 1 2539
2 55535 1 2539
2 55536 1 2559
2 55537 1 2559
2 55538 1 2560
2 55539 1 2560
2 55540 1 2560
2 55541 1 2560
2 55542 1 2561
2 55543 1 2561
2 55544 1 2561
2 55545 1 2561
2 55546 1 2562
2 55547 1 2562
2 55548 1 2562
2 55549 1 2563
2 55550 1 2563
2 55551 1 2563
2 55552 1 2563
2 55553 1 2564
2 55554 1 2564
2 55555 1 2564
2 55556 1 2564
2 55557 1 2564
2 55558 1 2564
2 55559 1 2564
2 55560 1 2564
2 55561 1 2564
2 55562 1 2564
2 55563 1 2564
2 55564 1 2564
2 55565 1 2564
2 55566 1 2564
2 55567 1 2564
2 55568 1 2564
2 55569 1 2564
2 55570 1 2564
2 55571 1 2564
2 55572 1 2564
2 55573 1 2564
2 55574 1 2564
2 55575 1 2564
2 55576 1 2564
2 55577 1 2564
2 55578 1 2564
2 55579 1 2564
2 55580 1 2564
2 55581 1 2564
2 55582 1 2564
2 55583 1 2564
2 55584 1 2564
2 55585 1 2564
2 55586 1 2564
2 55587 1 2564
2 55588 1 2564
2 55589 1 2564
2 55590 1 2564
2 55591 1 2564
2 55592 1 2564
2 55593 1 2564
2 55594 1 2564
2 55595 1 2564
2 55596 1 2564
2 55597 1 2565
2 55598 1 2565
2 55599 1 2565
2 55600 1 2565
2 55601 1 2565
2 55602 1 2565
2 55603 1 2565
2 55604 1 2565
2 55605 1 2565
2 55606 1 2565
2 55607 1 2565
2 55608 1 2565
2 55609 1 2565
2 55610 1 2565
2 55611 1 2565
2 55612 1 2565
2 55613 1 2565
2 55614 1 2565
2 55615 1 2565
2 55616 1 2565
2 55617 1 2565
2 55618 1 2565
2 55619 1 2565
2 55620 1 2565
2 55621 1 2565
2 55622 1 2565
2 55623 1 2565
2 55624 1 2565
2 55625 1 2565
2 55626 1 2565
2 55627 1 2565
2 55628 1 2565
2 55629 1 2565
2 55630 1 2565
2 55631 1 2565
2 55632 1 2565
2 55633 1 2565
2 55634 1 2565
2 55635 1 2569
2 55636 1 2569
2 55637 1 2570
2 55638 1 2570
2 55639 1 2570
2 55640 1 2570
2 55641 1 2570
2 55642 1 2570
2 55643 1 2579
2 55644 1 2579
2 55645 1 2579
2 55646 1 2579
2 55647 1 2579
2 55648 1 2579
2 55649 1 2581
2 55650 1 2581
2 55651 1 2581
2 55652 1 2581
2 55653 1 2581
2 55654 1 2581
2 55655 1 2581
2 55656 1 2581
2 55657 1 2581
2 55658 1 2581
2 55659 1 2581
2 55660 1 2581
2 55661 1 2589
2 55662 1 2589
2 55663 1 2590
2 55664 1 2590
2 55665 1 2590
2 55666 1 2590
2 55667 1 2590
2 55668 1 2590
2 55669 1 2598
2 55670 1 2598
2 55671 1 2598
2 55672 1 2598
2 55673 1 2598
2 55674 1 2598
2 55675 1 2598
2 55676 1 2599
2 55677 1 2599
2 55678 1 2599
2 55679 1 2599
2 55680 1 2599
2 55681 1 2600
2 55682 1 2600
2 55683 1 2602
2 55684 1 2602
2 55685 1 2602
2 55686 1 2603
2 55687 1 2603
2 55688 1 2607
2 55689 1 2607
2 55690 1 2608
2 55691 1 2608
2 55692 1 2608
2 55693 1 2608
2 55694 1 2608
2 55695 1 2610
2 55696 1 2610
2 55697 1 2610
2 55698 1 2611
2 55699 1 2611
2 55700 1 2615
2 55701 1 2615
2 55702 1 2616
2 55703 1 2616
2 55704 1 2617
2 55705 1 2617
2 55706 1 2617
2 55707 1 2617
2 55708 1 2617
2 55709 1 2617
2 55710 1 2617
2 55711 1 2617
2 55712 1 2617
2 55713 1 2617
2 55714 1 2617
2 55715 1 2617
2 55716 1 2618
2 55717 1 2618
2 55718 1 2618
2 55719 1 2618
2 55720 1 2618
2 55721 1 2619
2 55722 1 2619
2 55723 1 2619
2 55724 1 2619
2 55725 1 2619
2 55726 1 2619
2 55727 1 2619
2 55728 1 2619
2 55729 1 2620
2 55730 1 2620
2 55731 1 2620
2 55732 1 2620
2 55733 1 2620
2 55734 1 2620
2 55735 1 2620
2 55736 1 2621
2 55737 1 2621
2 55738 1 2624
2 55739 1 2624
2 55740 1 2624
2 55741 1 2632
2 55742 1 2632
2 55743 1 2632
2 55744 1 2632
2 55745 1 2632
2 55746 1 2632
2 55747 1 2645
2 55748 1 2645
2 55749 1 2645
2 55750 1 2645
2 55751 1 2645
2 55752 1 2645
2 55753 1 2645
2 55754 1 2645
2 55755 1 2645
2 55756 1 2645
2 55757 1 2645
2 55758 1 2645
2 55759 1 2645
2 55760 1 2645
2 55761 1 2645
2 55762 1 2645
2 55763 1 2645
2 55764 1 2645
2 55765 1 2645
2 55766 1 2645
2 55767 1 2645
2 55768 1 2645
2 55769 1 2645
2 55770 1 2647
2 55771 1 2647
2 55772 1 2647
2 55773 1 2647
2 55774 1 2647
2 55775 1 2647
2 55776 1 2647
2 55777 1 2647
2 55778 1 2647
2 55779 1 2647
2 55780 1 2647
2 55781 1 2647
2 55782 1 2647
2 55783 1 2647
2 55784 1 2647
2 55785 1 2647
2 55786 1 2647
2 55787 1 2647
2 55788 1 2648
2 55789 1 2648
2 55790 1 2648
2 55791 1 2651
2 55792 1 2651
2 55793 1 2651
2 55794 1 2651
2 55795 1 2651
2 55796 1 2651
2 55797 1 2651
2 55798 1 2651
2 55799 1 2651
2 55800 1 2651
2 55801 1 2651
2 55802 1 2651
2 55803 1 2651
2 55804 1 2651
2 55805 1 2651
2 55806 1 2651
2 55807 1 2652
2 55808 1 2652
2 55809 1 2652
2 55810 1 2653
2 55811 1 2653
2 55812 1 2653
2 55813 1 2653
2 55814 1 2653
2 55815 1 2653
2 55816 1 2653
2 55817 1 2653
2 55818 1 2653
2 55819 1 2653
2 55820 1 2653
2 55821 1 2653
2 55822 1 2653
2 55823 1 2653
2 55824 1 2653
2 55825 1 2653
2 55826 1 2654
2 55827 1 2654
2 55828 1 2654
2 55829 1 2654
2 55830 1 2654
2 55831 1 2654
2 55832 1 2654
2 55833 1 2656
2 55834 1 2656
2 55835 1 2656
2 55836 1 2662
2 55837 1 2662
2 55838 1 2663
2 55839 1 2663
2 55840 1 2663
2 55841 1 2663
2 55842 1 2663
2 55843 1 2663
2 55844 1 2663
2 55845 1 2663
2 55846 1 2663
2 55847 1 2663
2 55848 1 2663
2 55849 1 2663
2 55850 1 2663
2 55851 1 2663
2 55852 1 2663
2 55853 1 2663
2 55854 1 2664
2 55855 1 2664
2 55856 1 2664
2 55857 1 2664
2 55858 1 2664
2 55859 1 2664
2 55860 1 2664
2 55861 1 2664
2 55862 1 2664
2 55863 1 2664
2 55864 1 2664
2 55865 1 2664
2 55866 1 2678
2 55867 1 2678
2 55868 1 2678
2 55869 1 2678
2 55870 1 2678
2 55871 1 2686
2 55872 1 2686
2 55873 1 2686
2 55874 1 2686
2 55875 1 2686
2 55876 1 2686
2 55877 1 2686
2 55878 1 2686
2 55879 1 2686
2 55880 1 2686
2 55881 1 2686
2 55882 1 2686
2 55883 1 2686
2 55884 1 2686
2 55885 1 2686
2 55886 1 2686
2 55887 1 2686
2 55888 1 2686
2 55889 1 2686
2 55890 1 2686
2 55891 1 2686
2 55892 1 2686
2 55893 1 2686
2 55894 1 2686
2 55895 1 2686
2 55896 1 2686
2 55897 1 2686
2 55898 1 2686
2 55899 1 2686
2 55900 1 2686
2 55901 1 2686
2 55902 1 2686
2 55903 1 2686
2 55904 1 2686
2 55905 1 2686
2 55906 1 2686
2 55907 1 2686
2 55908 1 2686
2 55909 1 2686
2 55910 1 2686
2 55911 1 2686
2 55912 1 2686
2 55913 1 2686
2 55914 1 2686
2 55915 1 2686
2 55916 1 2686
2 55917 1 2686
2 55918 1 2686
2 55919 1 2686
2 55920 1 2686
2 55921 1 2686
2 55922 1 2686
2 55923 1 2686
2 55924 1 2687
2 55925 1 2687
2 55926 1 2687
2 55927 1 2687
2 55928 1 2687
2 55929 1 2687
2 55930 1 2687
2 55931 1 2688
2 55932 1 2688
2 55933 1 2688
2 55934 1 2704
2 55935 1 2704
2 55936 1 2712
2 55937 1 2712
2 55938 1 2713
2 55939 1 2713
2 55940 1 2715
2 55941 1 2715
2 55942 1 2733
2 55943 1 2733
2 55944 1 2734
2 55945 1 2734
2 55946 1 2734
2 55947 1 2734
2 55948 1 2734
2 55949 1 2736
2 55950 1 2736
2 55951 1 2737
2 55952 1 2737
2 55953 1 2737
2 55954 1 2737
2 55955 1 2737
2 55956 1 2737
2 55957 1 2737
2 55958 1 2737
2 55959 1 2737
2 55960 1 2737
2 55961 1 2737
2 55962 1 2737
2 55963 1 2737
2 55964 1 2737
2 55965 1 2737
2 55966 1 2737
2 55967 1 2737
2 55968 1 2737
2 55969 1 2745
2 55970 1 2745
2 55971 1 2745
2 55972 1 2745
2 55973 1 2745
2 55974 1 2745
2 55975 1 2745
2 55976 1 2745
2 55977 1 2752
2 55978 1 2752
2 55979 1 2755
2 55980 1 2755
2 55981 1 2759
2 55982 1 2759
2 55983 1 2761
2 55984 1 2761
2 55985 1 2767
2 55986 1 2767
2 55987 1 2767
2 55988 1 2767
2 55989 1 2767
2 55990 1 2767
2 55991 1 2767
2 55992 1 2767
2 55993 1 2767
2 55994 1 2767
2 55995 1 2767
2 55996 1 2767
2 55997 1 2770
2 55998 1 2770
2 55999 1 2778
2 56000 1 2778
2 56001 1 2778
2 56002 1 2778
2 56003 1 2779
2 56004 1 2779
2 56005 1 2779
2 56006 1 2793
2 56007 1 2793
2 56008 1 2804
2 56009 1 2804
2 56010 1 2805
2 56011 1 2805
2 56012 1 2805
2 56013 1 2805
2 56014 1 2805
2 56015 1 2805
2 56016 1 2805
2 56017 1 2805
2 56018 1 2805
2 56019 1 2805
2 56020 1 2805
2 56021 1 2805
2 56022 1 2805
2 56023 1 2805
2 56024 1 2806
2 56025 1 2806
2 56026 1 2806
2 56027 1 2808
2 56028 1 2808
2 56029 1 2819
2 56030 1 2819
2 56031 1 2819
2 56032 1 2819
2 56033 1 2819
2 56034 1 2819
2 56035 1 2819
2 56036 1 2820
2 56037 1 2820
2 56038 1 2820
2 56039 1 2820
2 56040 1 2820
2 56041 1 2820
2 56042 1 2820
2 56043 1 2820
2 56044 1 2821
2 56045 1 2821
2 56046 1 2826
2 56047 1 2826
2 56048 1 2827
2 56049 1 2827
2 56050 1 2827
2 56051 1 2834
2 56052 1 2834
2 56053 1 2835
2 56054 1 2835
2 56055 1 2835
2 56056 1 2836
2 56057 1 2836
2 56058 1 2836
2 56059 1 2845
2 56060 1 2845
2 56061 1 2845
2 56062 1 2845
2 56063 1 2845
2 56064 1 2845
2 56065 1 2847
2 56066 1 2847
2 56067 1 2859
2 56068 1 2859
2 56069 1 2859
2 56070 1 2859
2 56071 1 2866
2 56072 1 2866
2 56073 1 2866
2 56074 1 2866
2 56075 1 2866
2 56076 1 2866
2 56077 1 2866
2 56078 1 2866
2 56079 1 2867
2 56080 1 2867
2 56081 1 2868
2 56082 1 2868
2 56083 1 2868
2 56084 1 2869
2 56085 1 2869
2 56086 1 2869
2 56087 1 2869
2 56088 1 2869
2 56089 1 2882
2 56090 1 2882
2 56091 1 2885
2 56092 1 2885
2 56093 1 2885
2 56094 1 2885
2 56095 1 2885
2 56096 1 2885
2 56097 1 2886
2 56098 1 2886
2 56099 1 2886
2 56100 1 2894
2 56101 1 2894
2 56102 1 2894
2 56103 1 2894
2 56104 1 2894
2 56105 1 2894
2 56106 1 2894
2 56107 1 2894
2 56108 1 2894
2 56109 1 2894
2 56110 1 2896
2 56111 1 2896
2 56112 1 2896
2 56113 1 2899
2 56114 1 2899
2 56115 1 2899
2 56116 1 2899
2 56117 1 2900
2 56118 1 2900
2 56119 1 2900
2 56120 1 2900
2 56121 1 2900
2 56122 1 2900
2 56123 1 2900
2 56124 1 2900
2 56125 1 2900
2 56126 1 2900
2 56127 1 2900
2 56128 1 2908
2 56129 1 2908
2 56130 1 2911
2 56131 1 2911
2 56132 1 2911
2 56133 1 2911
2 56134 1 2911
2 56135 1 2911
2 56136 1 2911
2 56137 1 2912
2 56138 1 2912
2 56139 1 2912
2 56140 1 2913
2 56141 1 2913
2 56142 1 2913
2 56143 1 2913
2 56144 1 2913
2 56145 1 2913
2 56146 1 2914
2 56147 1 2914
2 56148 1 2925
2 56149 1 2925
2 56150 1 2925
2 56151 1 2926
2 56152 1 2926
2 56153 1 2943
2 56154 1 2943
2 56155 1 2943
2 56156 1 2955
2 56157 1 2955
2 56158 1 2955
2 56159 1 2955
2 56160 1 2955
2 56161 1 2955
2 56162 1 2955
2 56163 1 2955
2 56164 1 2956
2 56165 1 2956
2 56166 1 2956
2 56167 1 2956
2 56168 1 2963
2 56169 1 2963
2 56170 1 2964
2 56171 1 2964
2 56172 1 2965
2 56173 1 2965
2 56174 1 2965
2 56175 1 2968
2 56176 1 2968
2 56177 1 2968
2 56178 1 2968
2 56179 1 2968
2 56180 1 2968
2 56181 1 2969
2 56182 1 2969
2 56183 1 2969
2 56184 1 2969
2 56185 1 2969
2 56186 1 2969
2 56187 1 2969
2 56188 1 2969
2 56189 1 2969
2 56190 1 2969
2 56191 1 2969
2 56192 1 2969
2 56193 1 2969
2 56194 1 2970
2 56195 1 2970
2 56196 1 2970
2 56197 1 2972
2 56198 1 2972
2 56199 1 2972
2 56200 1 2972
2 56201 1 2972
2 56202 1 2973
2 56203 1 2973
2 56204 1 2973
2 56205 1 2981
2 56206 1 2981
2 56207 1 2981
2 56208 1 2981
2 56209 1 2981
2 56210 1 2981
2 56211 1 2981
2 56212 1 2981
2 56213 1 2981
2 56214 1 2981
2 56215 1 2981
2 56216 1 2981
2 56217 1 2981
2 56218 1 2981
2 56219 1 2981
2 56220 1 2981
2 56221 1 2981
2 56222 1 2981
2 56223 1 2981
2 56224 1 2981
2 56225 1 2981
2 56226 1 2983
2 56227 1 2983
2 56228 1 2983
2 56229 1 2983
2 56230 1 2983
2 56231 1 2983
2 56232 1 2983
2 56233 1 2983
2 56234 1 2983
2 56235 1 2983
2 56236 1 2983
2 56237 1 2983
2 56238 1 2983
2 56239 1 2983
2 56240 1 2983
2 56241 1 2983
2 56242 1 2983
2 56243 1 2983
2 56244 1 2984
2 56245 1 2984
2 56246 1 2984
2 56247 1 2985
2 56248 1 2985
2 56249 1 2985
2 56250 1 2985
2 56251 1 2985
2 56252 1 2985
2 56253 1 2985
2 56254 1 2985
2 56255 1 2986
2 56256 1 2986
2 56257 1 2987
2 56258 1 2987
2 56259 1 2987
2 56260 1 2987
2 56261 1 2987
2 56262 1 2987
2 56263 1 2987
2 56264 1 2987
2 56265 1 2987
2 56266 1 2987
2 56267 1 2987
2 56268 1 2996
2 56269 1 2996
2 56270 1 2996
2 56271 1 2996
2 56272 1 3000
2 56273 1 3000
2 56274 1 3000
2 56275 1 3000
2 56276 1 3000
2 56277 1 3000
2 56278 1 3000
2 56279 1 3000
2 56280 1 3000
2 56281 1 3000
2 56282 1 3000
2 56283 1 3000
2 56284 1 3000
2 56285 1 3000
2 56286 1 3000
2 56287 1 3000
2 56288 1 3000
2 56289 1 3001
2 56290 1 3001
2 56291 1 3001
2 56292 1 3001
2 56293 1 3001
2 56294 1 3001
2 56295 1 3009
2 56296 1 3009
2 56297 1 3011
2 56298 1 3011
2 56299 1 3011
2 56300 1 3011
2 56301 1 3013
2 56302 1 3013
2 56303 1 3013
2 56304 1 3013
2 56305 1 3042
2 56306 1 3042
2 56307 1 3042
2 56308 1 3042
2 56309 1 3042
2 56310 1 3042
2 56311 1 3042
2 56312 1 3043
2 56313 1 3043
2 56314 1 3044
2 56315 1 3044
2 56316 1 3045
2 56317 1 3045
2 56318 1 3045
2 56319 1 3052
2 56320 1 3052
2 56321 1 3052
2 56322 1 3052
2 56323 1 3052
2 56324 1 3052
2 56325 1 3052
2 56326 1 3052
2 56327 1 3054
2 56328 1 3054
2 56329 1 3055
2 56330 1 3055
2 56331 1 3055
2 56332 1 3060
2 56333 1 3060
2 56334 1 3060
2 56335 1 3071
2 56336 1 3071
2 56337 1 3071
2 56338 1 3071
2 56339 1 3071
2 56340 1 3071
2 56341 1 3071
2 56342 1 3072
2 56343 1 3072
2 56344 1 3078
2 56345 1 3078
2 56346 1 3078
2 56347 1 3078
2 56348 1 3078
2 56349 1 3078
2 56350 1 3078
2 56351 1 3078
2 56352 1 3078
2 56353 1 3078
2 56354 1 3078
2 56355 1 3078
2 56356 1 3078
2 56357 1 3078
2 56358 1 3078
2 56359 1 3078
2 56360 1 3078
2 56361 1 3079
2 56362 1 3079
2 56363 1 3084
2 56364 1 3084
2 56365 1 3086
2 56366 1 3086
2 56367 1 3086
2 56368 1 3086
2 56369 1 3086
2 56370 1 3087
2 56371 1 3087
2 56372 1 3090
2 56373 1 3090
2 56374 1 3090
2 56375 1 3090
2 56376 1 3090
2 56377 1 3090
2 56378 1 3113
2 56379 1 3113
2 56380 1 3114
2 56381 1 3114
2 56382 1 3127
2 56383 1 3127
2 56384 1 3132
2 56385 1 3132
2 56386 1 3135
2 56387 1 3135
2 56388 1 3141
2 56389 1 3141
2 56390 1 3141
2 56391 1 3141
2 56392 1 3141
2 56393 1 3141
2 56394 1 3141
2 56395 1 3141
2 56396 1 3141
2 56397 1 3142
2 56398 1 3142
2 56399 1 3142
2 56400 1 3142
2 56401 1 3144
2 56402 1 3144
2 56403 1 3146
2 56404 1 3146
2 56405 1 3146
2 56406 1 3146
2 56407 1 3146
2 56408 1 3157
2 56409 1 3157
2 56410 1 3157
2 56411 1 3158
2 56412 1 3158
2 56413 1 3162
2 56414 1 3162
2 56415 1 3162
2 56416 1 3162
2 56417 1 3162
2 56418 1 3162
2 56419 1 3162
2 56420 1 3162
2 56421 1 3162
2 56422 1 3162
2 56423 1 3162
2 56424 1 3162
2 56425 1 3162
2 56426 1 3162
2 56427 1 3162
2 56428 1 3162
2 56429 1 3162
2 56430 1 3162
2 56431 1 3162
2 56432 1 3163
2 56433 1 3163
2 56434 1 3163
2 56435 1 3163
2 56436 1 3163
2 56437 1 3164
2 56438 1 3164
2 56439 1 3164
2 56440 1 3164
2 56441 1 3164
2 56442 1 3164
2 56443 1 3165
2 56444 1 3165
2 56445 1 3167
2 56446 1 3167
2 56447 1 3169
2 56448 1 3169
2 56449 1 3169
2 56450 1 3169
2 56451 1 3169
2 56452 1 3184
2 56453 1 3184
2 56454 1 3184
2 56455 1 3184
2 56456 1 3184
2 56457 1 3184
2 56458 1 3184
2 56459 1 3185
2 56460 1 3185
2 56461 1 3185
2 56462 1 3185
2 56463 1 3186
2 56464 1 3186
2 56465 1 3186
2 56466 1 3190
2 56467 1 3190
2 56468 1 3196
2 56469 1 3196
2 56470 1 3203
2 56471 1 3203
2 56472 1 3203
2 56473 1 3204
2 56474 1 3204
2 56475 1 3204
2 56476 1 3204
2 56477 1 3204
2 56478 1 3204
2 56479 1 3204
2 56480 1 3204
2 56481 1 3204
2 56482 1 3207
2 56483 1 3207
2 56484 1 3207
2 56485 1 3208
2 56486 1 3208
2 56487 1 3208
2 56488 1 3208
2 56489 1 3208
2 56490 1 3208
2 56491 1 3208
2 56492 1 3209
2 56493 1 3209
2 56494 1 3210
2 56495 1 3210
2 56496 1 3219
2 56497 1 3219
2 56498 1 3219
2 56499 1 3219
2 56500 1 3219
2 56501 1 3219
2 56502 1 3219
2 56503 1 3223
2 56504 1 3223
2 56505 1 3223
2 56506 1 3223
2 56507 1 3223
2 56508 1 3223
2 56509 1 3223
2 56510 1 3224
2 56511 1 3224
2 56512 1 3224
2 56513 1 3224
2 56514 1 3224
2 56515 1 3225
2 56516 1 3225
2 56517 1 3226
2 56518 1 3226
2 56519 1 3226
2 56520 1 3226
2 56521 1 3226
2 56522 1 3227
2 56523 1 3227
2 56524 1 3227
2 56525 1 3227
2 56526 1 3227
2 56527 1 3227
2 56528 1 3237
2 56529 1 3237
2 56530 1 3240
2 56531 1 3240
2 56532 1 3240
2 56533 1 3240
2 56534 1 3241
2 56535 1 3241
2 56536 1 3249
2 56537 1 3249
2 56538 1 3249
2 56539 1 3250
2 56540 1 3250
2 56541 1 3250
2 56542 1 3258
2 56543 1 3258
2 56544 1 3258
2 56545 1 3266
2 56546 1 3266
2 56547 1 3267
2 56548 1 3267
2 56549 1 3267
2 56550 1 3267
2 56551 1 3267
2 56552 1 3268
2 56553 1 3268
2 56554 1 3268
2 56555 1 3271
2 56556 1 3271
2 56557 1 3271
2 56558 1 3271
2 56559 1 3271
2 56560 1 3312
2 56561 1 3312
2 56562 1 3312
2 56563 1 3312
2 56564 1 3312
2 56565 1 3312
2 56566 1 3322
2 56567 1 3322
2 56568 1 3322
2 56569 1 3322
2 56570 1 3322
2 56571 1 3322
2 56572 1 3330
2 56573 1 3330
2 56574 1 3330
2 56575 1 3333
2 56576 1 3333
2 56577 1 3333
2 56578 1 3334
2 56579 1 3334
2 56580 1 3342
2 56581 1 3342
2 56582 1 3342
2 56583 1 3342
2 56584 1 3342
2 56585 1 3342
2 56586 1 3342
2 56587 1 3342
2 56588 1 3342
2 56589 1 3342
2 56590 1 3342
2 56591 1 3342
2 56592 1 3342
2 56593 1 3343
2 56594 1 3343
2 56595 1 3343
2 56596 1 3345
2 56597 1 3345
2 56598 1 3345
2 56599 1 3346
2 56600 1 3346
2 56601 1 3346
2 56602 1 3358
2 56603 1 3358
2 56604 1 3359
2 56605 1 3359
2 56606 1 3361
2 56607 1 3361
2 56608 1 3361
2 56609 1 3371
2 56610 1 3371
2 56611 1 3371
2 56612 1 3371
2 56613 1 3376
2 56614 1 3376
2 56615 1 3376
2 56616 1 3376
2 56617 1 3385
2 56618 1 3385
2 56619 1 3385
2 56620 1 3385
2 56621 1 3386
2 56622 1 3386
2 56623 1 3388
2 56624 1 3388
2 56625 1 3391
2 56626 1 3391
2 56627 1 3391
2 56628 1 3391
2 56629 1 3393
2 56630 1 3393
2 56631 1 3408
2 56632 1 3408
2 56633 1 3408
2 56634 1 3408
2 56635 1 3408
2 56636 1 3408
2 56637 1 3409
2 56638 1 3409
2 56639 1 3409
2 56640 1 3415
2 56641 1 3415
2 56642 1 3441
2 56643 1 3441
2 56644 1 3441
2 56645 1 3441
2 56646 1 3441
2 56647 1 3441
2 56648 1 3442
2 56649 1 3442
2 56650 1 3442
2 56651 1 3442
2 56652 1 3442
2 56653 1 3442
2 56654 1 3442
2 56655 1 3442
2 56656 1 3442
2 56657 1 3442
2 56658 1 3442
2 56659 1 3442
2 56660 1 3442
2 56661 1 3442
2 56662 1 3442
2 56663 1 3442
2 56664 1 3443
2 56665 1 3443
2 56666 1 3445
2 56667 1 3445
2 56668 1 3445
2 56669 1 3445
2 56670 1 3446
2 56671 1 3446
2 56672 1 3446
2 56673 1 3449
2 56674 1 3449
2 56675 1 3449
2 56676 1 3450
2 56677 1 3450
2 56678 1 3454
2 56679 1 3454
2 56680 1 3455
2 56681 1 3455
2 56682 1 3455
2 56683 1 3456
2 56684 1 3456
2 56685 1 3456
2 56686 1 3456
2 56687 1 3457
2 56688 1 3457
2 56689 1 3457
2 56690 1 3462
2 56691 1 3462
2 56692 1 3463
2 56693 1 3463
2 56694 1 3471
2 56695 1 3471
2 56696 1 3471
2 56697 1 3471
2 56698 1 3471
2 56699 1 3478
2 56700 1 3478
2 56701 1 3478
2 56702 1 3478
2 56703 1 3478
2 56704 1 3478
2 56705 1 3478
2 56706 1 3478
2 56707 1 3479
2 56708 1 3479
2 56709 1 3480
2 56710 1 3480
2 56711 1 3480
2 56712 1 3480
2 56713 1 3480
2 56714 1 3480
2 56715 1 3482
2 56716 1 3482
2 56717 1 3482
2 56718 1 3483
2 56719 1 3483
2 56720 1 3491
2 56721 1 3491
2 56722 1 3491
2 56723 1 3491
2 56724 1 3500
2 56725 1 3500
2 56726 1 3500
2 56727 1 3500
2 56728 1 3500
2 56729 1 3500
2 56730 1 3500
2 56731 1 3500
2 56732 1 3500
2 56733 1 3502
2 56734 1 3502
2 56735 1 3505
2 56736 1 3505
2 56737 1 3505
2 56738 1 3505
2 56739 1 3505
2 56740 1 3505
2 56741 1 3505
2 56742 1 3506
2 56743 1 3506
2 56744 1 3506
2 56745 1 3506
2 56746 1 3506
2 56747 1 3506
2 56748 1 3506
2 56749 1 3506
2 56750 1 3506
2 56751 1 3506
2 56752 1 3506
2 56753 1 3506
2 56754 1 3506
2 56755 1 3506
2 56756 1 3513
2 56757 1 3513
2 56758 1 3513
2 56759 1 3513
2 56760 1 3521
2 56761 1 3521
2 56762 1 3521
2 56763 1 3521
2 56764 1 3524
2 56765 1 3524
2 56766 1 3524
2 56767 1 3524
2 56768 1 3525
2 56769 1 3525
2 56770 1 3525
2 56771 1 3526
2 56772 1 3526
2 56773 1 3534
2 56774 1 3534
2 56775 1 3534
2 56776 1 3534
2 56777 1 3534
2 56778 1 3534
2 56779 1 3534
2 56780 1 3534
2 56781 1 3534
2 56782 1 3534
2 56783 1 3534
2 56784 1 3534
2 56785 1 3534
2 56786 1 3535
2 56787 1 3535
2 56788 1 3535
2 56789 1 3535
2 56790 1 3536
2 56791 1 3536
2 56792 1 3536
2 56793 1 3536
2 56794 1 3536
2 56795 1 3537
2 56796 1 3537
2 56797 1 3537
2 56798 1 3537
2 56799 1 3537
2 56800 1 3537
2 56801 1 3537
2 56802 1 3537
2 56803 1 3539
2 56804 1 3539
2 56805 1 3543
2 56806 1 3543
2 56807 1 3546
2 56808 1 3546
2 56809 1 3551
2 56810 1 3551
2 56811 1 3563
2 56812 1 3563
2 56813 1 3563
2 56814 1 3563
2 56815 1 3563
2 56816 1 3563
2 56817 1 3563
2 56818 1 3563
2 56819 1 3563
2 56820 1 3563
2 56821 1 3563
2 56822 1 3563
2 56823 1 3563
2 56824 1 3563
2 56825 1 3563
2 56826 1 3563
2 56827 1 3563
2 56828 1 3565
2 56829 1 3565
2 56830 1 3565
2 56831 1 3565
2 56832 1 3565
2 56833 1 3566
2 56834 1 3566
2 56835 1 3566
2 56836 1 3575
2 56837 1 3575
2 56838 1 3575
2 56839 1 3576
2 56840 1 3576
2 56841 1 3576
2 56842 1 3576
2 56843 1 3577
2 56844 1 3577
2 56845 1 3578
2 56846 1 3578
2 56847 1 3578
2 56848 1 3579
2 56849 1 3579
2 56850 1 3579
2 56851 1 3579
2 56852 1 3579
2 56853 1 3583
2 56854 1 3583
2 56855 1 3583
2 56856 1 3583
2 56857 1 3585
2 56858 1 3585
2 56859 1 3586
2 56860 1 3586
2 56861 1 3586
2 56862 1 3586
2 56863 1 3596
2 56864 1 3596
2 56865 1 3596
2 56866 1 3596
2 56867 1 3596
2 56868 1 3596
2 56869 1 3596
2 56870 1 3596
2 56871 1 3596
2 56872 1 3596
2 56873 1 3596
2 56874 1 3596
2 56875 1 3596
2 56876 1 3596
2 56877 1 3596
2 56878 1 3596
2 56879 1 3596
2 56880 1 3597
2 56881 1 3597
2 56882 1 3605
2 56883 1 3605
2 56884 1 3605
2 56885 1 3605
2 56886 1 3605
2 56887 1 3605
2 56888 1 3605
2 56889 1 3605
2 56890 1 3605
2 56891 1 3605
2 56892 1 3605
2 56893 1 3606
2 56894 1 3606
2 56895 1 3606
2 56896 1 3606
2 56897 1 3607
2 56898 1 3607
2 56899 1 3607
2 56900 1 3608
2 56901 1 3608
2 56902 1 3608
2 56903 1 3609
2 56904 1 3609
2 56905 1 3609
2 56906 1 3609
2 56907 1 3609
2 56908 1 3609
2 56909 1 3609
2 56910 1 3609
2 56911 1 3610
2 56912 1 3610
2 56913 1 3611
2 56914 1 3611
2 56915 1 3611
2 56916 1 3611
2 56917 1 3611
2 56918 1 3611
2 56919 1 3611
2 56920 1 3611
2 56921 1 3611
2 56922 1 3611
2 56923 1 3611
2 56924 1 3612
2 56925 1 3612
2 56926 1 3612
2 56927 1 3612
2 56928 1 3612
2 56929 1 3613
2 56930 1 3613
2 56931 1 3617
2 56932 1 3617
2 56933 1 3617
2 56934 1 3617
2 56935 1 3620
2 56936 1 3620
2 56937 1 3620
2 56938 1 3620
2 56939 1 3621
2 56940 1 3621
2 56941 1 3621
2 56942 1 3621
2 56943 1 3621
2 56944 1 3622
2 56945 1 3622
2 56946 1 3623
2 56947 1 3623
2 56948 1 3623
2 56949 1 3623
2 56950 1 3623
2 56951 1 3623
2 56952 1 3623
2 56953 1 3623
2 56954 1 3623
2 56955 1 3623
2 56956 1 3623
2 56957 1 3623
2 56958 1 3623
2 56959 1 3623
2 56960 1 3623
2 56961 1 3623
2 56962 1 3624
2 56963 1 3624
2 56964 1 3624
2 56965 1 3624
2 56966 1 3627
2 56967 1 3627
2 56968 1 3627
2 56969 1 3627
2 56970 1 3627
2 56971 1 3627
2 56972 1 3627
2 56973 1 3627
2 56974 1 3627
2 56975 1 3627
2 56976 1 3627
2 56977 1 3634
2 56978 1 3634
2 56979 1 3641
2 56980 1 3641
2 56981 1 3649
2 56982 1 3649
2 56983 1 3649
2 56984 1 3651
2 56985 1 3651
2 56986 1 3652
2 56987 1 3652
2 56988 1 3653
2 56989 1 3653
2 56990 1 3654
2 56991 1 3654
2 56992 1 3654
2 56993 1 3654
2 56994 1 3654
2 56995 1 3654
2 56996 1 3654
2 56997 1 3654
2 56998 1 3667
2 56999 1 3667
2 57000 1 3667
2 57001 1 3674
2 57002 1 3674
2 57003 1 3674
2 57004 1 3674
2 57005 1 3688
2 57006 1 3688
2 57007 1 3688
2 57008 1 3688
2 57009 1 3688
2 57010 1 3688
2 57011 1 3688
2 57012 1 3688
2 57013 1 3688
2 57014 1 3688
2 57015 1 3688
2 57016 1 3688
2 57017 1 3688
2 57018 1 3688
2 57019 1 3688
2 57020 1 3688
2 57021 1 3689
2 57022 1 3689
2 57023 1 3689
2 57024 1 3691
2 57025 1 3691
2 57026 1 3691
2 57027 1 3691
2 57028 1 3691
2 57029 1 3691
2 57030 1 3692
2 57031 1 3692
2 57032 1 3693
2 57033 1 3693
2 57034 1 3693
2 57035 1 3697
2 57036 1 3697
2 57037 1 3697
2 57038 1 3697
2 57039 1 3697
2 57040 1 3697
2 57041 1 3698
2 57042 1 3698
2 57043 1 3698
2 57044 1 3702
2 57045 1 3702
2 57046 1 3710
2 57047 1 3710
2 57048 1 3716
2 57049 1 3716
2 57050 1 3716
2 57051 1 3716
2 57052 1 3716
2 57053 1 3716
2 57054 1 3716
2 57055 1 3716
2 57056 1 3716
2 57057 1 3717
2 57058 1 3717
2 57059 1 3718
2 57060 1 3718
2 57061 1 3721
2 57062 1 3721
2 57063 1 3721
2 57064 1 3722
2 57065 1 3722
2 57066 1 3724
2 57067 1 3724
2 57068 1 3724
2 57069 1 3734
2 57070 1 3734
2 57071 1 3735
2 57072 1 3735
2 57073 1 3735
2 57074 1 3735
2 57075 1 3736
2 57076 1 3736
2 57077 1 3736
2 57078 1 3741
2 57079 1 3741
2 57080 1 3741
2 57081 1 3741
2 57082 1 3741
2 57083 1 3741
2 57084 1 3742
2 57085 1 3742
2 57086 1 3743
2 57087 1 3743
2 57088 1 3743
2 57089 1 3743
2 57090 1 3743
2 57091 1 3743
2 57092 1 3743
2 57093 1 3744
2 57094 1 3744
2 57095 1 3745
2 57096 1 3745
2 57097 1 3745
2 57098 1 3745
2 57099 1 3745
2 57100 1 3745
2 57101 1 3745
2 57102 1 3745
2 57103 1 3745
2 57104 1 3746
2 57105 1 3746
2 57106 1 3747
2 57107 1 3747
2 57108 1 3747
2 57109 1 3747
2 57110 1 3747
2 57111 1 3747
2 57112 1 3747
2 57113 1 3747
2 57114 1 3747
2 57115 1 3754
2 57116 1 3754
2 57117 1 3754
2 57118 1 3754
2 57119 1 3754
2 57120 1 3754
2 57121 1 3755
2 57122 1 3755
2 57123 1 3755
2 57124 1 3755
2 57125 1 3757
2 57126 1 3757
2 57127 1 3757
2 57128 1 3759
2 57129 1 3759
2 57130 1 3764
2 57131 1 3764
2 57132 1 3764
2 57133 1 3764
2 57134 1 3764
2 57135 1 3773
2 57136 1 3773
2 57137 1 3773
2 57138 1 3773
2 57139 1 3773
2 57140 1 3774
2 57141 1 3774
2 57142 1 3774
2 57143 1 3774
2 57144 1 3774
2 57145 1 3775
2 57146 1 3775
2 57147 1 3776
2 57148 1 3776
2 57149 1 3776
2 57150 1 3776
2 57151 1 3776
2 57152 1 3776
2 57153 1 3776
2 57154 1 3778
2 57155 1 3778
2 57156 1 3781
2 57157 1 3781
2 57158 1 3782
2 57159 1 3782
2 57160 1 3784
2 57161 1 3784
2 57162 1 3784
2 57163 1 3784
2 57164 1 3784
2 57165 1 3784
2 57166 1 3784
2 57167 1 3785
2 57168 1 3785
2 57169 1 3792
2 57170 1 3792
2 57171 1 3793
2 57172 1 3793
2 57173 1 3793
2 57174 1 3794
2 57175 1 3794
2 57176 1 3795
2 57177 1 3795
2 57178 1 3795
2 57179 1 3795
2 57180 1 3795
2 57181 1 3795
2 57182 1 3795
2 57183 1 3795
2 57184 1 3795
2 57185 1 3795
2 57186 1 3795
2 57187 1 3795
2 57188 1 3799
2 57189 1 3799
2 57190 1 3800
2 57191 1 3800
2 57192 1 3800
2 57193 1 3800
2 57194 1 3800
2 57195 1 3800
2 57196 1 3800
2 57197 1 3800
2 57198 1 3800
2 57199 1 3800
2 57200 1 3800
2 57201 1 3800
2 57202 1 3800
2 57203 1 3800
2 57204 1 3800
2 57205 1 3803
2 57206 1 3803
2 57207 1 3803
2 57208 1 3803
2 57209 1 3803
2 57210 1 3803
2 57211 1 3803
2 57212 1 3805
2 57213 1 3805
2 57214 1 3805
2 57215 1 3805
2 57216 1 3805
2 57217 1 3813
2 57218 1 3813
2 57219 1 3813
2 57220 1 3813
2 57221 1 3813
2 57222 1 3813
2 57223 1 3813
2 57224 1 3813
2 57225 1 3813
2 57226 1 3813
2 57227 1 3814
2 57228 1 3814
2 57229 1 3815
2 57230 1 3815
2 57231 1 3819
2 57232 1 3819
2 57233 1 3819
2 57234 1 3819
2 57235 1 3819
2 57236 1 3821
2 57237 1 3821
2 57238 1 3822
2 57239 1 3822
2 57240 1 3830
2 57241 1 3830
2 57242 1 3830
2 57243 1 3830
2 57244 1 3830
2 57245 1 3830
2 57246 1 3830
2 57247 1 3830
2 57248 1 3830
2 57249 1 3830
2 57250 1 3830
2 57251 1 3831
2 57252 1 3831
2 57253 1 3831
2 57254 1 3831
2 57255 1 3831
2 57256 1 3832
2 57257 1 3832
2 57258 1 3834
2 57259 1 3834
2 57260 1 3840
2 57261 1 3840
2 57262 1 3840
2 57263 1 3849
2 57264 1 3849
2 57265 1 3849
2 57266 1 3849
2 57267 1 3849
2 57268 1 3852
2 57269 1 3852
2 57270 1 3853
2 57271 1 3853
2 57272 1 3854
2 57273 1 3854
2 57274 1 3854
2 57275 1 3854
2 57276 1 3854
2 57277 1 3855
2 57278 1 3855
2 57279 1 3855
2 57280 1 3855
2 57281 1 3855
2 57282 1 3855
2 57283 1 3869
2 57284 1 3869
2 57285 1 3873
2 57286 1 3873
2 57287 1 3873
2 57288 1 3873
2 57289 1 3873
2 57290 1 3873
2 57291 1 3873
2 57292 1 3873
2 57293 1 3874
2 57294 1 3874
2 57295 1 3876
2 57296 1 3876
2 57297 1 3877
2 57298 1 3877
2 57299 1 3882
2 57300 1 3882
2 57301 1 3882
2 57302 1 3883
2 57303 1 3883
2 57304 1 3893
2 57305 1 3893
2 57306 1 3893
2 57307 1 3893
2 57308 1 3893
2 57309 1 3893
2 57310 1 3893
2 57311 1 3893
2 57312 1 3893
2 57313 1 3893
2 57314 1 3893
2 57315 1 3894
2 57316 1 3894
2 57317 1 3894
2 57318 1 3905
2 57319 1 3905
2 57320 1 3905
2 57321 1 3905
2 57322 1 3905
2 57323 1 3905
2 57324 1 3905
2 57325 1 3905
2 57326 1 3906
2 57327 1 3906
2 57328 1 3906
2 57329 1 3907
2 57330 1 3907
2 57331 1 3907
2 57332 1 3908
2 57333 1 3908
2 57334 1 3908
2 57335 1 3910
2 57336 1 3910
2 57337 1 3911
2 57338 1 3911
2 57339 1 3916
2 57340 1 3916
2 57341 1 3916
2 57342 1 3916
2 57343 1 3916
2 57344 1 3916
2 57345 1 3916
2 57346 1 3916
2 57347 1 3916
2 57348 1 3916
2 57349 1 3916
2 57350 1 3916
2 57351 1 3916
2 57352 1 3916
2 57353 1 3916
2 57354 1 3916
2 57355 1 3916
2 57356 1 3916
2 57357 1 3918
2 57358 1 3918
2 57359 1 3918
2 57360 1 3918
2 57361 1 3918
2 57362 1 3918
2 57363 1 3918
2 57364 1 3918
2 57365 1 3918
2 57366 1 3933
2 57367 1 3933
2 57368 1 3933
2 57369 1 3933
2 57370 1 3933
2 57371 1 3933
2 57372 1 3933
2 57373 1 3933
2 57374 1 3933
2 57375 1 3933
2 57376 1 3933
2 57377 1 3933
2 57378 1 3933
2 57379 1 3933
2 57380 1 3933
2 57381 1 3933
2 57382 1 3933
2 57383 1 3938
2 57384 1 3938
2 57385 1 3939
2 57386 1 3939
2 57387 1 3939
2 57388 1 3953
2 57389 1 3953
2 57390 1 3953
2 57391 1 3953
2 57392 1 3954
2 57393 1 3954
2 57394 1 3954
2 57395 1 3954
2 57396 1 3954
2 57397 1 3954
2 57398 1 3954
2 57399 1 3954
2 57400 1 3954
2 57401 1 3954
2 57402 1 3954
2 57403 1 3954
2 57404 1 3954
2 57405 1 3955
2 57406 1 3955
2 57407 1 3965
2 57408 1 3965
2 57409 1 3966
2 57410 1 3966
2 57411 1 3968
2 57412 1 3968
2 57413 1 3968
2 57414 1 3968
2 57415 1 3968
2 57416 1 3982
2 57417 1 3982
2 57418 1 3982
2 57419 1 3982
2 57420 1 3982
2 57421 1 3982
2 57422 1 3982
2 57423 1 3982
2 57424 1 3982
2 57425 1 3982
2 57426 1 3983
2 57427 1 3983
2 57428 1 3983
2 57429 1 3983
2 57430 1 3986
2 57431 1 3986
2 57432 1 3986
2 57433 1 3986
2 57434 1 3986
2 57435 1 3986
2 57436 1 3986
2 57437 1 3987
2 57438 1 3987
2 57439 1 3994
2 57440 1 3994
2 57441 1 3994
2 57442 1 4001
2 57443 1 4001
2 57444 1 4013
2 57445 1 4013
2 57446 1 4013
2 57447 1 4014
2 57448 1 4014
2 57449 1 4015
2 57450 1 4015
2 57451 1 4015
2 57452 1 4016
2 57453 1 4016
2 57454 1 4018
2 57455 1 4018
2 57456 1 4021
2 57457 1 4021
2 57458 1 4021
2 57459 1 4021
2 57460 1 4021
2 57461 1 4021
2 57462 1 4021
2 57463 1 4021
2 57464 1 4022
2 57465 1 4022
2 57466 1 4033
2 57467 1 4033
2 57468 1 4043
2 57469 1 4043
2 57470 1 4056
2 57471 1 4056
2 57472 1 4059
2 57473 1 4059
2 57474 1 4060
2 57475 1 4060
2 57476 1 4061
2 57477 1 4061
2 57478 1 4061
2 57479 1 4061
2 57480 1 4061
2 57481 1 4070
2 57482 1 4070
2 57483 1 4070
2 57484 1 4070
2 57485 1 4070
2 57486 1 4070
2 57487 1 4071
2 57488 1 4071
2 57489 1 4086
2 57490 1 4086
2 57491 1 4086
2 57492 1 4086
2 57493 1 4086
2 57494 1 4086
2 57495 1 4086
2 57496 1 4086
2 57497 1 4086
2 57498 1 4087
2 57499 1 4087
2 57500 1 4087
2 57501 1 4087
2 57502 1 4087
2 57503 1 4087
2 57504 1 4088
2 57505 1 4088
2 57506 1 4096
2 57507 1 4096
2 57508 1 4096
2 57509 1 4096
2 57510 1 4097
2 57511 1 4097
2 57512 1 4101
2 57513 1 4101
2 57514 1 4101
2 57515 1 4101
2 57516 1 4101
2 57517 1 4101
2 57518 1 4111
2 57519 1 4111
2 57520 1 4112
2 57521 1 4112
2 57522 1 4112
2 57523 1 4112
2 57524 1 4114
2 57525 1 4114
2 57526 1 4114
2 57527 1 4114
2 57528 1 4116
2 57529 1 4116
2 57530 1 4124
2 57531 1 4124
2 57532 1 4124
2 57533 1 4124
2 57534 1 4124
2 57535 1 4124
2 57536 1 4124
2 57537 1 4125
2 57538 1 4125
2 57539 1 4125
2 57540 1 4127
2 57541 1 4127
2 57542 1 4127
2 57543 1 4127
2 57544 1 4129
2 57545 1 4129
2 57546 1 4130
2 57547 1 4130
2 57548 1 4130
2 57549 1 4130
2 57550 1 4130
2 57551 1 4130
2 57552 1 4130
2 57553 1 4130
2 57554 1 4130
2 57555 1 4131
2 57556 1 4131
2 57557 1 4131
2 57558 1 4131
2 57559 1 4131
2 57560 1 4131
2 57561 1 4131
2 57562 1 4131
2 57563 1 4131
2 57564 1 4131
2 57565 1 4131
2 57566 1 4131
2 57567 1 4132
2 57568 1 4132
2 57569 1 4132
2 57570 1 4132
2 57571 1 4137
2 57572 1 4137
2 57573 1 4141
2 57574 1 4141
2 57575 1 4141
2 57576 1 4141
2 57577 1 4141
2 57578 1 4141
2 57579 1 4141
2 57580 1 4141
2 57581 1 4142
2 57582 1 4142
2 57583 1 4143
2 57584 1 4143
2 57585 1 4143
2 57586 1 4147
2 57587 1 4147
2 57588 1 4148
2 57589 1 4148
2 57590 1 4149
2 57591 1 4149
2 57592 1 4149
2 57593 1 4149
2 57594 1 4149
2 57595 1 4149
2 57596 1 4149
2 57597 1 4149
2 57598 1 4149
2 57599 1 4162
2 57600 1 4162
2 57601 1 4162
2 57602 1 4162
2 57603 1 4163
2 57604 1 4163
2 57605 1 4163
2 57606 1 4163
2 57607 1 4163
2 57608 1 4163
2 57609 1 4163
2 57610 1 4163
2 57611 1 4163
2 57612 1 4163
2 57613 1 4163
2 57614 1 4163
2 57615 1 4163
2 57616 1 4163
2 57617 1 4164
2 57618 1 4164
2 57619 1 4164
2 57620 1 4164
2 57621 1 4164
2 57622 1 4165
2 57623 1 4165
2 57624 1 4165
2 57625 1 4165
2 57626 1 4165
2 57627 1 4165
2 57628 1 4165
2 57629 1 4165
2 57630 1 4165
2 57631 1 4165
2 57632 1 4165
2 57633 1 4165
2 57634 1 4165
2 57635 1 4165
2 57636 1 4165
2 57637 1 4165
2 57638 1 4165
2 57639 1 4165
2 57640 1 4165
2 57641 1 4165
2 57642 1 4165
2 57643 1 4165
2 57644 1 4165
2 57645 1 4165
2 57646 1 4165
2 57647 1 4165
2 57648 1 4179
2 57649 1 4179
2 57650 1 4180
2 57651 1 4180
2 57652 1 4180
2 57653 1 4180
2 57654 1 4180
2 57655 1 4180
2 57656 1 4180
2 57657 1 4181
2 57658 1 4181
2 57659 1 4181
2 57660 1 4181
2 57661 1 4181
2 57662 1 4184
2 57663 1 4184
2 57664 1 4199
2 57665 1 4199
2 57666 1 4199
2 57667 1 4199
2 57668 1 4204
2 57669 1 4204
2 57670 1 4213
2 57671 1 4213
2 57672 1 4219
2 57673 1 4219
2 57674 1 4220
2 57675 1 4220
2 57676 1 4227
2 57677 1 4227
2 57678 1 4232
2 57679 1 4232
2 57680 1 4233
2 57681 1 4233
2 57682 1 4233
2 57683 1 4233
2 57684 1 4233
2 57685 1 4233
2 57686 1 4233
2 57687 1 4233
2 57688 1 4242
2 57689 1 4242
2 57690 1 4242
2 57691 1 4243
2 57692 1 4243
2 57693 1 4243
2 57694 1 4246
2 57695 1 4246
2 57696 1 4246
2 57697 1 4246
2 57698 1 4246
2 57699 1 4250
2 57700 1 4250
2 57701 1 4250
2 57702 1 4251
2 57703 1 4251
2 57704 1 4251
2 57705 1 4259
2 57706 1 4259
2 57707 1 4259
2 57708 1 4262
2 57709 1 4262
2 57710 1 4263
2 57711 1 4263
2 57712 1 4263
2 57713 1 4268
2 57714 1 4268
2 57715 1 4268
2 57716 1 4268
2 57717 1 4268
2 57718 1 4277
2 57719 1 4277
2 57720 1 4277
2 57721 1 4277
2 57722 1 4277
2 57723 1 4277
2 57724 1 4278
2 57725 1 4278
2 57726 1 4279
2 57727 1 4279
2 57728 1 4279
2 57729 1 4280
2 57730 1 4280
2 57731 1 4283
2 57732 1 4283
2 57733 1 4284
2 57734 1 4284
2 57735 1 4284
2 57736 1 4284
2 57737 1 4284
2 57738 1 4284
2 57739 1 4293
2 57740 1 4293
2 57741 1 4293
2 57742 1 4293
2 57743 1 4293
2 57744 1 4294
2 57745 1 4294
2 57746 1 4308
2 57747 1 4308
2 57748 1 4308
2 57749 1 4308
2 57750 1 4308
2 57751 1 4308
2 57752 1 4308
2 57753 1 4308
2 57754 1 4310
2 57755 1 4310
2 57756 1 4328
2 57757 1 4328
2 57758 1 4340
2 57759 1 4340
2 57760 1 4340
2 57761 1 4340
2 57762 1 4340
2 57763 1 4340
2 57764 1 4340
2 57765 1 4341
2 57766 1 4341
2 57767 1 4341
2 57768 1 4341
2 57769 1 4341
2 57770 1 4341
2 57771 1 4341
2 57772 1 4350
2 57773 1 4350
2 57774 1 4350
2 57775 1 4350
2 57776 1 4350
2 57777 1 4350
2 57778 1 4351
2 57779 1 4351
2 57780 1 4351
2 57781 1 4351
2 57782 1 4351
2 57783 1 4351
2 57784 1 4351
2 57785 1 4351
2 57786 1 4351
2 57787 1 4351
2 57788 1 4351
2 57789 1 4351
2 57790 1 4351
2 57791 1 4351
2 57792 1 4353
2 57793 1 4353
2 57794 1 4355
2 57795 1 4355
2 57796 1 4358
2 57797 1 4358
2 57798 1 4358
2 57799 1 4358
2 57800 1 4358
2 57801 1 4358
2 57802 1 4361
2 57803 1 4361
2 57804 1 4361
2 57805 1 4370
2 57806 1 4370
2 57807 1 4370
2 57808 1 4382
2 57809 1 4382
2 57810 1 4384
2 57811 1 4384
2 57812 1 4384
2 57813 1 4384
2 57814 1 4384
2 57815 1 4385
2 57816 1 4385
2 57817 1 4385
2 57818 1 4386
2 57819 1 4386
2 57820 1 4388
2 57821 1 4388
2 57822 1 4395
2 57823 1 4395
2 57824 1 4396
2 57825 1 4396
2 57826 1 4397
2 57827 1 4397
2 57828 1 4397
2 57829 1 4398
2 57830 1 4398
2 57831 1 4400
2 57832 1 4400
2 57833 1 4405
2 57834 1 4405
2 57835 1 4405
2 57836 1 4405
2 57837 1 4405
2 57838 1 4405
2 57839 1 4405
2 57840 1 4405
2 57841 1 4405
2 57842 1 4421
2 57843 1 4421
2 57844 1 4431
2 57845 1 4431
2 57846 1 4431
2 57847 1 4431
2 57848 1 4432
2 57849 1 4432
2 57850 1 4438
2 57851 1 4438
2 57852 1 4438
2 57853 1 4438
2 57854 1 4438
2 57855 1 4438
2 57856 1 4438
2 57857 1 4452
2 57858 1 4452
2 57859 1 4458
2 57860 1 4458
2 57861 1 4458
2 57862 1 4459
2 57863 1 4459
2 57864 1 4460
2 57865 1 4460
2 57866 1 4460
2 57867 1 4460
2 57868 1 4460
2 57869 1 4460
2 57870 1 4461
2 57871 1 4461
2 57872 1 4475
2 57873 1 4475
2 57874 1 4475
2 57875 1 4475
2 57876 1 4475
2 57877 1 4475
2 57878 1 4487
2 57879 1 4487
2 57880 1 4489
2 57881 1 4489
2 57882 1 4489
2 57883 1 4489
2 57884 1 4492
2 57885 1 4492
2 57886 1 4492
2 57887 1 4492
2 57888 1 4499
2 57889 1 4499
2 57890 1 4499
2 57891 1 4499
2 57892 1 4499
2 57893 1 4507
2 57894 1 4507
2 57895 1 4508
2 57896 1 4508
2 57897 1 4511
2 57898 1 4511
2 57899 1 4511
2 57900 1 4511
2 57901 1 4511
2 57902 1 4519
2 57903 1 4519
2 57904 1 4531
2 57905 1 4531
2 57906 1 4531
2 57907 1 4531
2 57908 1 4531
2 57909 1 4531
2 57910 1 4531
2 57911 1 4531
2 57912 1 4531
2 57913 1 4531
2 57914 1 4531
2 57915 1 4531
2 57916 1 4531
2 57917 1 4531
2 57918 1 4531
2 57919 1 4531
2 57920 1 4531
2 57921 1 4531
2 57922 1 4531
2 57923 1 4531
2 57924 1 4531
2 57925 1 4531
2 57926 1 4531
2 57927 1 4532
2 57928 1 4532
2 57929 1 4532
2 57930 1 4532
2 57931 1 4537
2 57932 1 4537
2 57933 1 4537
2 57934 1 4541
2 57935 1 4541
2 57936 1 4541
2 57937 1 4541
2 57938 1 4541
2 57939 1 4541
2 57940 1 4541
2 57941 1 4541
2 57942 1 4541
2 57943 1 4541
2 57944 1 4541
2 57945 1 4541
2 57946 1 4541
2 57947 1 4541
2 57948 1 4541
2 57949 1 4541
2 57950 1 4542
2 57951 1 4542
2 57952 1 4542
2 57953 1 4542
2 57954 1 4551
2 57955 1 4551
2 57956 1 4554
2 57957 1 4554
2 57958 1 4575
2 57959 1 4575
2 57960 1 4576
2 57961 1 4576
2 57962 1 4576
2 57963 1 4576
2 57964 1 4580
2 57965 1 4580
2 57966 1 4580
2 57967 1 4580
2 57968 1 4580
2 57969 1 4581
2 57970 1 4581
2 57971 1 4581
2 57972 1 4581
2 57973 1 4582
2 57974 1 4582
2 57975 1 4589
2 57976 1 4589
2 57977 1 4589
2 57978 1 4589
2 57979 1 4589
2 57980 1 4589
2 57981 1 4589
2 57982 1 4589
2 57983 1 4589
2 57984 1 4635
2 57985 1 4635
2 57986 1 4643
2 57987 1 4643
2 57988 1 4643
2 57989 1 4643
2 57990 1 4643
2 57991 1 4643
2 57992 1 4643
2 57993 1 4643
2 57994 1 4643
2 57995 1 4643
2 57996 1 4644
2 57997 1 4644
2 57998 1 4644
2 57999 1 4644
2 58000 1 4644
2 58001 1 4647
2 58002 1 4647
2 58003 1 4647
2 58004 1 4647
2 58005 1 4647
2 58006 1 4655
2 58007 1 4655
2 58008 1 4656
2 58009 1 4656
2 58010 1 4656
2 58011 1 4656
2 58012 1 4656
2 58013 1 4656
2 58014 1 4656
2 58015 1 4670
2 58016 1 4670
2 58017 1 4671
2 58018 1 4671
2 58019 1 4671
2 58020 1 4671
2 58021 1 4671
2 58022 1 4671
2 58023 1 4671
2 58024 1 4671
2 58025 1 4671
2 58026 1 4671
2 58027 1 4673
2 58028 1 4673
2 58029 1 4682
2 58030 1 4682
2 58031 1 4684
2 58032 1 4684
2 58033 1 4695
2 58034 1 4695
2 58035 1 4695
2 58036 1 4696
2 58037 1 4696
2 58038 1 4697
2 58039 1 4697
2 58040 1 4697
2 58041 1 4697
2 58042 1 4697
2 58043 1 4705
2 58044 1 4705
2 58045 1 4724
2 58046 1 4724
2 58047 1 4724
2 58048 1 4724
2 58049 1 4724
2 58050 1 4724
2 58051 1 4724
2 58052 1 4725
2 58053 1 4725
2 58054 1 4728
2 58055 1 4728
2 58056 1 4728
2 58057 1 4731
2 58058 1 4731
2 58059 1 4731
2 58060 1 4731
2 58061 1 4731
2 58062 1 4731
2 58063 1 4731
2 58064 1 4731
2 58065 1 4731
2 58066 1 4731
2 58067 1 4731
2 58068 1 4731
2 58069 1 4731
2 58070 1 4732
2 58071 1 4732
2 58072 1 4732
2 58073 1 4734
2 58074 1 4734
2 58075 1 4734
2 58076 1 4734
2 58077 1 4734
2 58078 1 4734
2 58079 1 4734
2 58080 1 4734
2 58081 1 4734
2 58082 1 4735
2 58083 1 4735
2 58084 1 4735
2 58085 1 4752
2 58086 1 4752
2 58087 1 4752
2 58088 1 4752
2 58089 1 4752
2 58090 1 4752
2 58091 1 4752
2 58092 1 4752
2 58093 1 4754
2 58094 1 4754
2 58095 1 4754
2 58096 1 4754
2 58097 1 4754
2 58098 1 4754
2 58099 1 4754
2 58100 1 4761
2 58101 1 4761
2 58102 1 4761
2 58103 1 4772
2 58104 1 4772
2 58105 1 4772
2 58106 1 4772
2 58107 1 4772
2 58108 1 4772
2 58109 1 4774
2 58110 1 4774
2 58111 1 4774
2 58112 1 4774
2 58113 1 4774
2 58114 1 4774
2 58115 1 4774
2 58116 1 4774
2 58117 1 4776
2 58118 1 4776
2 58119 1 4776
2 58120 1 4776
2 58121 1 4776
2 58122 1 4777
2 58123 1 4777
2 58124 1 4777
2 58125 1 4777
2 58126 1 4777
2 58127 1 4780
2 58128 1 4780
2 58129 1 4780
2 58130 1 4780
2 58131 1 4780
2 58132 1 4780
2 58133 1 4780
2 58134 1 4780
2 58135 1 4780
2 58136 1 4780
2 58137 1 4780
2 58138 1 4780
2 58139 1 4780
2 58140 1 4780
2 58141 1 4780
2 58142 1 4780
2 58143 1 4781
2 58144 1 4781
2 58145 1 4781
2 58146 1 4781
2 58147 1 4782
2 58148 1 4782
2 58149 1 4790
2 58150 1 4790
2 58151 1 4791
2 58152 1 4791
2 58153 1 4800
2 58154 1 4800
2 58155 1 4800
2 58156 1 4800
2 58157 1 4800
2 58158 1 4800
2 58159 1 4800
2 58160 1 4800
2 58161 1 4800
2 58162 1 4800
2 58163 1 4801
2 58164 1 4801
2 58165 1 4810
2 58166 1 4810
2 58167 1 4810
2 58168 1 4810
2 58169 1 4810
2 58170 1 4812
2 58171 1 4812
2 58172 1 4812
2 58173 1 4812
2 58174 1 4812
2 58175 1 4812
2 58176 1 4812
2 58177 1 4812
2 58178 1 4812
2 58179 1 4812
2 58180 1 4812
2 58181 1 4812
2 58182 1 4812
2 58183 1 4812
2 58184 1 4812
2 58185 1 4812
2 58186 1 4812
2 58187 1 4812
2 58188 1 4812
2 58189 1 4812
2 58190 1 4812
2 58191 1 4812
2 58192 1 4812
2 58193 1 4812
2 58194 1 4812
2 58195 1 4812
2 58196 1 4812
2 58197 1 4812
2 58198 1 4812
2 58199 1 4812
2 58200 1 4812
2 58201 1 4812
2 58202 1 4812
2 58203 1 4812
2 58204 1 4812
2 58205 1 4812
2 58206 1 4813
2 58207 1 4813
2 58208 1 4814
2 58209 1 4814
2 58210 1 4821
2 58211 1 4821
2 58212 1 4821
2 58213 1 4826
2 58214 1 4826
2 58215 1 4828
2 58216 1 4828
2 58217 1 4828
2 58218 1 4828
2 58219 1 4828
2 58220 1 4829
2 58221 1 4829
2 58222 1 4838
2 58223 1 4838
2 58224 1 4838
2 58225 1 4838
2 58226 1 4838
2 58227 1 4838
2 58228 1 4838
2 58229 1 4838
2 58230 1 4838
2 58231 1 4838
2 58232 1 4840
2 58233 1 4840
2 58234 1 4841
2 58235 1 4841
2 58236 1 4841
2 58237 1 4841
2 58238 1 4841
2 58239 1 4841
2 58240 1 4841
2 58241 1 4841
2 58242 1 4841
2 58243 1 4841
2 58244 1 4841
2 58245 1 4841
2 58246 1 4841
2 58247 1 4841
2 58248 1 4841
2 58249 1 4841
2 58250 1 4842
2 58251 1 4842
2 58252 1 4842
2 58253 1 4846
2 58254 1 4846
2 58255 1 4846
2 58256 1 4846
2 58257 1 4846
2 58258 1 4846
2 58259 1 4846
2 58260 1 4846
2 58261 1 4846
2 58262 1 4846
2 58263 1 4846
2 58264 1 4846
2 58265 1 4847
2 58266 1 4847
2 58267 1 4848
2 58268 1 4848
2 58269 1 4848
2 58270 1 4848
2 58271 1 4848
2 58272 1 4848
2 58273 1 4849
2 58274 1 4849
2 58275 1 4849
2 58276 1 4849
2 58277 1 4849
2 58278 1 4849
2 58279 1 4849
2 58280 1 4849
2 58281 1 4849
2 58282 1 4849
2 58283 1 4849
2 58284 1 4849
2 58285 1 4849
2 58286 1 4849
2 58287 1 4856
2 58288 1 4856
2 58289 1 4856
2 58290 1 4856
2 58291 1 4856
2 58292 1 4856
2 58293 1 4856
2 58294 1 4856
2 58295 1 4856
2 58296 1 4856
2 58297 1 4857
2 58298 1 4857
2 58299 1 4865
2 58300 1 4865
2 58301 1 4866
2 58302 1 4866
2 58303 1 4866
2 58304 1 4866
2 58305 1 4866
2 58306 1 4866
2 58307 1 4866
2 58308 1 4866
2 58309 1 4866
2 58310 1 4866
2 58311 1 4868
2 58312 1 4868
2 58313 1 4868
2 58314 1 4868
2 58315 1 4869
2 58316 1 4869
2 58317 1 4873
2 58318 1 4873
2 58319 1 4873
2 58320 1 4873
2 58321 1 4886
2 58322 1 4886
2 58323 1 4887
2 58324 1 4887
2 58325 1 4887
2 58326 1 4887
2 58327 1 4896
2 58328 1 4896
2 58329 1 4908
2 58330 1 4908
2 58331 1 4924
2 58332 1 4924
2 58333 1 4935
2 58334 1 4935
2 58335 1 4935
2 58336 1 4935
2 58337 1 4935
2 58338 1 4936
2 58339 1 4936
2 58340 1 4937
2 58341 1 4937
2 58342 1 4937
2 58343 1 4937
2 58344 1 4937
2 58345 1 4937
2 58346 1 4937
2 58347 1 4937
2 58348 1 4937
2 58349 1 4937
2 58350 1 4937
2 58351 1 4938
2 58352 1 4938
2 58353 1 4939
2 58354 1 4939
2 58355 1 4940
2 58356 1 4940
2 58357 1 4940
2 58358 1 4940
2 58359 1 4940
2 58360 1 4940
2 58361 1 4940
2 58362 1 4940
2 58363 1 4940
2 58364 1 4943
2 58365 1 4943
2 58366 1 4943
2 58367 1 4943
2 58368 1 4943
2 58369 1 4943
2 58370 1 4943
2 58371 1 4943
2 58372 1 4943
2 58373 1 4943
2 58374 1 4943
2 58375 1 4943
2 58376 1 4943
2 58377 1 4943
2 58378 1 4943
2 58379 1 4944
2 58380 1 4944
2 58381 1 4944
2 58382 1 4945
2 58383 1 4945
2 58384 1 4945
2 58385 1 4955
2 58386 1 4955
2 58387 1 4955
2 58388 1 4957
2 58389 1 4957
2 58390 1 4961
2 58391 1 4961
2 58392 1 4969
2 58393 1 4969
2 58394 1 4969
2 58395 1 4969
2 58396 1 4969
2 58397 1 4969
2 58398 1 4969
2 58399 1 4969
2 58400 1 4969
2 58401 1 4969
2 58402 1 4987
2 58403 1 4987
2 58404 1 4988
2 58405 1 4988
2 58406 1 4988
2 58407 1 4996
2 58408 1 4996
2 58409 1 4996
2 58410 1 4996
2 58411 1 5010
2 58412 1 5010
2 58413 1 5010
2 58414 1 5010
2 58415 1 5010
2 58416 1 5010
2 58417 1 5010
2 58418 1 5010
2 58419 1 5010
2 58420 1 5010
2 58421 1 5011
2 58422 1 5011
2 58423 1 5011
2 58424 1 5011
2 58425 1 5012
2 58426 1 5012
2 58427 1 5012
2 58428 1 5012
2 58429 1 5020
2 58430 1 5020
2 58431 1 5020
2 58432 1 5020
2 58433 1 5020
2 58434 1 5020
2 58435 1 5020
2 58436 1 5020
2 58437 1 5023
2 58438 1 5023
2 58439 1 5047
2 58440 1 5047
2 58441 1 5047
2 58442 1 5051
2 58443 1 5051
2 58444 1 5051
2 58445 1 5051
2 58446 1 5052
2 58447 1 5052
2 58448 1 5052
2 58449 1 5052
2 58450 1 5052
2 58451 1 5053
2 58452 1 5053
2 58453 1 5068
2 58454 1 5068
2 58455 1 5075
2 58456 1 5075
2 58457 1 5075
2 58458 1 5076
2 58459 1 5076
2 58460 1 5076
2 58461 1 5079
2 58462 1 5079
2 58463 1 5079
2 58464 1 5080
2 58465 1 5080
2 58466 1 5080
2 58467 1 5083
2 58468 1 5083
2 58469 1 5084
2 58470 1 5084
2 58471 1 5085
2 58472 1 5085
2 58473 1 5085
2 58474 1 5086
2 58475 1 5086
2 58476 1 5088
2 58477 1 5088
2 58478 1 5100
2 58479 1 5100
2 58480 1 5100
2 58481 1 5100
2 58482 1 5100
2 58483 1 5101
2 58484 1 5101
2 58485 1 5101
2 58486 1 5102
2 58487 1 5102
2 58488 1 5103
2 58489 1 5103
2 58490 1 5105
2 58491 1 5105
2 58492 1 5105
2 58493 1 5105
2 58494 1 5105
2 58495 1 5105
2 58496 1 5105
2 58497 1 5105
2 58498 1 5105
2 58499 1 5105
2 58500 1 5120
2 58501 1 5120
2 58502 1 5120
2 58503 1 5120
2 58504 1 5121
2 58505 1 5121
2 58506 1 5122
2 58507 1 5122
2 58508 1 5122
2 58509 1 5133
2 58510 1 5133
2 58511 1 5146
2 58512 1 5146
2 58513 1 5147
2 58514 1 5147
2 58515 1 5165
2 58516 1 5165
2 58517 1 5174
2 58518 1 5174
2 58519 1 5174
2 58520 1 5174
2 58521 1 5190
2 58522 1 5190
2 58523 1 5197
2 58524 1 5197
2 58525 1 5198
2 58526 1 5198
2 58527 1 5215
2 58528 1 5215
2 58529 1 5215
2 58530 1 5215
2 58531 1 5215
2 58532 1 5216
2 58533 1 5216
2 58534 1 5233
2 58535 1 5233
2 58536 1 5233
2 58537 1 5234
2 58538 1 5234
2 58539 1 5239
2 58540 1 5239
2 58541 1 5239
2 58542 1 5240
2 58543 1 5240
2 58544 1 5259
2 58545 1 5259
2 58546 1 5259
2 58547 1 5259
2 58548 1 5260
2 58549 1 5260
2 58550 1 5260
2 58551 1 5260
2 58552 1 5260
2 58553 1 5262
2 58554 1 5262
2 58555 1 5262
2 58556 1 5262
2 58557 1 5262
2 58558 1 5262
2 58559 1 5262
2 58560 1 5263
2 58561 1 5263
2 58562 1 5264
2 58563 1 5264
2 58564 1 5264
2 58565 1 5264
2 58566 1 5264
2 58567 1 5264
2 58568 1 5264
2 58569 1 5264
2 58570 1 5264
2 58571 1 5264
2 58572 1 5265
2 58573 1 5265
2 58574 1 5265
2 58575 1 5265
2 58576 1 5265
2 58577 1 5265
2 58578 1 5265
2 58579 1 5265
2 58580 1 5265
2 58581 1 5274
2 58582 1 5274
2 58583 1 5275
2 58584 1 5275
2 58585 1 5275
2 58586 1 5284
2 58587 1 5284
2 58588 1 5284
2 58589 1 5284
2 58590 1 5284
2 58591 1 5284
2 58592 1 5284
2 58593 1 5293
2 58594 1 5293
2 58595 1 5293
2 58596 1 5324
2 58597 1 5324
2 58598 1 5324
2 58599 1 5324
2 58600 1 5324
2 58601 1 5325
2 58602 1 5325
2 58603 1 5326
2 58604 1 5326
2 58605 1 5334
2 58606 1 5334
2 58607 1 5338
2 58608 1 5338
2 58609 1 5338
2 58610 1 5338
2 58611 1 5338
2 58612 1 5338
2 58613 1 5338
2 58614 1 5338
2 58615 1 5340
2 58616 1 5340
2 58617 1 5341
2 58618 1 5341
2 58619 1 5344
2 58620 1 5344
2 58621 1 5345
2 58622 1 5345
2 58623 1 5345
2 58624 1 5352
2 58625 1 5352
2 58626 1 5352
2 58627 1 5352
2 58628 1 5352
2 58629 1 5352
2 58630 1 5356
2 58631 1 5356
2 58632 1 5356
2 58633 1 5356
2 58634 1 5356
2 58635 1 5356
2 58636 1 5356
2 58637 1 5356
2 58638 1 5364
2 58639 1 5364
2 58640 1 5389
2 58641 1 5389
2 58642 1 5389
2 58643 1 5389
2 58644 1 5389
2 58645 1 5402
2 58646 1 5402
2 58647 1 5402
2 58648 1 5404
2 58649 1 5404
2 58650 1 5404
2 58651 1 5405
2 58652 1 5405
2 58653 1 5405
2 58654 1 5406
2 58655 1 5406
2 58656 1 5412
2 58657 1 5412
2 58658 1 5412
2 58659 1 5421
2 58660 1 5421
2 58661 1 5421
2 58662 1 5431
2 58663 1 5431
2 58664 1 5431
2 58665 1 5431
2 58666 1 5431
2 58667 1 5452
2 58668 1 5452
2 58669 1 5453
2 58670 1 5453
2 58671 1 5453
2 58672 1 5453
2 58673 1 5453
2 58674 1 5453
2 58675 1 5454
2 58676 1 5454
2 58677 1 5454
2 58678 1 5457
2 58679 1 5457
2 58680 1 5457
2 58681 1 5458
2 58682 1 5458
2 58683 1 5458
2 58684 1 5458
2 58685 1 5465
2 58686 1 5465
2 58687 1 5465
2 58688 1 5465
2 58689 1 5465
2 58690 1 5465
2 58691 1 5474
2 58692 1 5474
2 58693 1 5474
2 58694 1 5474
2 58695 1 5474
2 58696 1 5475
2 58697 1 5475
2 58698 1 5475
2 58699 1 5476
2 58700 1 5476
2 58701 1 5476
2 58702 1 5477
2 58703 1 5477
2 58704 1 5477
2 58705 1 5478
2 58706 1 5478
2 58707 1 5481
2 58708 1 5481
2 58709 1 5484
2 58710 1 5484
2 58711 1 5484
2 58712 1 5484
2 58713 1 5484
2 58714 1 5484
2 58715 1 5484
2 58716 1 5484
2 58717 1 5484
2 58718 1 5484
2 58719 1 5484
2 58720 1 5484
2 58721 1 5484
2 58722 1 5484
2 58723 1 5484
2 58724 1 5484
2 58725 1 5484
2 58726 1 5484
2 58727 1 5484
2 58728 1 5484
2 58729 1 5491
2 58730 1 5491
2 58731 1 5491
2 58732 1 5491
2 58733 1 5491
2 58734 1 5503
2 58735 1 5503
2 58736 1 5503
2 58737 1 5503
2 58738 1 5503
2 58739 1 5503
2 58740 1 5503
2 58741 1 5503
2 58742 1 5504
2 58743 1 5504
2 58744 1 5506
2 58745 1 5506
2 58746 1 5509
2 58747 1 5509
2 58748 1 5509
2 58749 1 5509
2 58750 1 5509
2 58751 1 5510
2 58752 1 5510
2 58753 1 5510
2 58754 1 5510
2 58755 1 5511
2 58756 1 5511
2 58757 1 5545
2 58758 1 5545
2 58759 1 5549
2 58760 1 5549
2 58761 1 5552
2 58762 1 5552
2 58763 1 5552
2 58764 1 5560
2 58765 1 5560
2 58766 1 5560
2 58767 1 5560
2 58768 1 5560
2 58769 1 5562
2 58770 1 5562
2 58771 1 5563
2 58772 1 5563
2 58773 1 5563
2 58774 1 5563
2 58775 1 5564
2 58776 1 5564
2 58777 1 5569
2 58778 1 5569
2 58779 1 5586
2 58780 1 5586
2 58781 1 5587
2 58782 1 5587
2 58783 1 5595
2 58784 1 5595
2 58785 1 5596
2 58786 1 5596
2 58787 1 5596
2 58788 1 5596
2 58789 1 5596
2 58790 1 5596
2 58791 1 5596
2 58792 1 5596
2 58793 1 5596
2 58794 1 5596
2 58795 1 5597
2 58796 1 5597
2 58797 1 5598
2 58798 1 5598
2 58799 1 5598
2 58800 1 5599
2 58801 1 5599
2 58802 1 5604
2 58803 1 5604
2 58804 1 5604
2 58805 1 5604
2 58806 1 5604
2 58807 1 5605
2 58808 1 5605
2 58809 1 5606
2 58810 1 5606
2 58811 1 5606
2 58812 1 5619
2 58813 1 5619
2 58814 1 5621
2 58815 1 5621
2 58816 1 5621
2 58817 1 5631
2 58818 1 5631
2 58819 1 5637
2 58820 1 5637
2 58821 1 5638
2 58822 1 5638
2 58823 1 5638
2 58824 1 5638
2 58825 1 5640
2 58826 1 5640
2 58827 1 5659
2 58828 1 5659
2 58829 1 5659
2 58830 1 5659
2 58831 1 5660
2 58832 1 5660
2 58833 1 5662
2 58834 1 5662
2 58835 1 5668
2 58836 1 5668
2 58837 1 5672
2 58838 1 5672
2 58839 1 5677
2 58840 1 5677
2 58841 1 5706
2 58842 1 5706
2 58843 1 5706
2 58844 1 5706
2 58845 1 5717
2 58846 1 5717
2 58847 1 5718
2 58848 1 5718
2 58849 1 5727
2 58850 1 5727
2 58851 1 5752
2 58852 1 5752
2 58853 1 5752
2 58854 1 5752
2 58855 1 5759
2 58856 1 5759
2 58857 1 5760
2 58858 1 5760
2 58859 1 5760
2 58860 1 5760
2 58861 1 5766
2 58862 1 5766
2 58863 1 5766
2 58864 1 5766
2 58865 1 5766
2 58866 1 5766
2 58867 1 5779
2 58868 1 5779
2 58869 1 5779
2 58870 1 5779
2 58871 1 5779
2 58872 1 5779
2 58873 1 5779
2 58874 1 5779
2 58875 1 5789
2 58876 1 5789
2 58877 1 5789
2 58878 1 5789
2 58879 1 5789
2 58880 1 5789
2 58881 1 5794
2 58882 1 5794
2 58883 1 5794
2 58884 1 5794
2 58885 1 5796
2 58886 1 5796
2 58887 1 5797
2 58888 1 5797
2 58889 1 5797
2 58890 1 5797
2 58891 1 5797
2 58892 1 5797
2 58893 1 5806
2 58894 1 5806
2 58895 1 5806
2 58896 1 5806
2 58897 1 5806
2 58898 1 5806
2 58899 1 5806
2 58900 1 5806
2 58901 1 5806
2 58902 1 5806
2 58903 1 5806
2 58904 1 5806
2 58905 1 5809
2 58906 1 5809
2 58907 1 5809
2 58908 1 5814
2 58909 1 5814
2 58910 1 5814
2 58911 1 5814
2 58912 1 5815
2 58913 1 5815
2 58914 1 5815
2 58915 1 5819
2 58916 1 5819
2 58917 1 5819
2 58918 1 5819
2 58919 1 5819
2 58920 1 5819
2 58921 1 5819
2 58922 1 5819
2 58923 1 5819
2 58924 1 5819
2 58925 1 5820
2 58926 1 5820
2 58927 1 5828
2 58928 1 5828
2 58929 1 5828
2 58930 1 5828
2 58931 1 5828
2 58932 1 5829
2 58933 1 5829
2 58934 1 5834
2 58935 1 5834
2 58936 1 5858
2 58937 1 5858
2 58938 1 5858
2 58939 1 5858
2 58940 1 5858
2 58941 1 5858
2 58942 1 5858
2 58943 1 5858
2 58944 1 5858
2 58945 1 5858
2 58946 1 5858
2 58947 1 5858
2 58948 1 5858
2 58949 1 5858
2 58950 1 5858
2 58951 1 5858
2 58952 1 5858
2 58953 1 5858
2 58954 1 5858
2 58955 1 5858
2 58956 1 5859
2 58957 1 5859
2 58958 1 5859
2 58959 1 5868
2 58960 1 5868
2 58961 1 5869
2 58962 1 5869
2 58963 1 5870
2 58964 1 5870
2 58965 1 5870
2 58966 1 5879
2 58967 1 5879
2 58968 1 5879
2 58969 1 5879
2 58970 1 5879
2 58971 1 5879
2 58972 1 5879
2 58973 1 5880
2 58974 1 5880
2 58975 1 5888
2 58976 1 5888
2 58977 1 5889
2 58978 1 5889
2 58979 1 5889
2 58980 1 5889
2 58981 1 5889
2 58982 1 5890
2 58983 1 5890
2 58984 1 5902
2 58985 1 5902
2 58986 1 5902
2 58987 1 5902
2 58988 1 5921
2 58989 1 5921
2 58990 1 5929
2 58991 1 5929
2 58992 1 5937
2 58993 1 5937
2 58994 1 5937
2 58995 1 5937
2 58996 1 5937
2 58997 1 5937
2 58998 1 5937
2 58999 1 5937
2 59000 1 5937
2 59001 1 5937
2 59002 1 5938
2 59003 1 5938
2 59004 1 5939
2 59005 1 5939
2 59006 1 5946
2 59007 1 5946
2 59008 1 5946
2 59009 1 5946
2 59010 1 5946
2 59011 1 5946
2 59012 1 5946
2 59013 1 5946
2 59014 1 5946
2 59015 1 5946
2 59016 1 5946
2 59017 1 5946
2 59018 1 5946
2 59019 1 5946
2 59020 1 5946
2 59021 1 5946
2 59022 1 5946
2 59023 1 5947
2 59024 1 5947
2 59025 1 5947
2 59026 1 5983
2 59027 1 5983
2 59028 1 5984
2 59029 1 5984
2 59030 1 5984
2 59031 1 5984
2 59032 1 5984
2 59033 1 5984
2 59034 1 5984
2 59035 1 5984
2 59036 1 5984
2 59037 1 5984
2 59038 1 5984
2 59039 1 5984
2 59040 1 5984
2 59041 1 5984
2 59042 1 5984
2 59043 1 5984
2 59044 1 5985
2 59045 1 5985
2 59046 1 5986
2 59047 1 5986
2 59048 1 5989
2 59049 1 5989
2 59050 1 5989
2 59051 1 5996
2 59052 1 5996
2 59053 1 6003
2 59054 1 6003
2 59055 1 6003
2 59056 1 6006
2 59057 1 6006
2 59058 1 6006
2 59059 1 6006
2 59060 1 6006
2 59061 1 6006
2 59062 1 6006
2 59063 1 6006
2 59064 1 6012
2 59065 1 6012
2 59066 1 6012
2 59067 1 6013
2 59068 1 6013
2 59069 1 6014
2 59070 1 6014
2 59071 1 6037
2 59072 1 6037
2 59073 1 6046
2 59074 1 6046
2 59075 1 6047
2 59076 1 6047
2 59077 1 6047
2 59078 1 6047
2 59079 1 6048
2 59080 1 6048
2 59081 1 6049
2 59082 1 6049
2 59083 1 6049
2 59084 1 6049
2 59085 1 6049
2 59086 1 6049
2 59087 1 6049
2 59088 1 6049
2 59089 1 6049
2 59090 1 6049
2 59091 1 6049
2 59092 1 6050
2 59093 1 6050
2 59094 1 6052
2 59095 1 6052
2 59096 1 6053
2 59097 1 6053
2 59098 1 6053
2 59099 1 6053
2 59100 1 6053
2 59101 1 6053
2 59102 1 6053
2 59103 1 6053
2 59104 1 6053
2 59105 1 6053
2 59106 1 6053
2 59107 1 6053
2 59108 1 6053
2 59109 1 6053
2 59110 1 6053
2 59111 1 6053
2 59112 1 6071
2 59113 1 6071
2 59114 1 6098
2 59115 1 6098
2 59116 1 6098
2 59117 1 6100
2 59118 1 6100
2 59119 1 6109
2 59120 1 6109
2 59121 1 6113
2 59122 1 6113
2 59123 1 6113
2 59124 1 6113
2 59125 1 6113
2 59126 1 6113
2 59127 1 6113
2 59128 1 6113
2 59129 1 6113
2 59130 1 6113
2 59131 1 6121
2 59132 1 6121
2 59133 1 6121
2 59134 1 6121
2 59135 1 6121
2 59136 1 6121
2 59137 1 6121
2 59138 1 6121
2 59139 1 6121
2 59140 1 6121
2 59141 1 6121
2 59142 1 6121
2 59143 1 6121
2 59144 1 6121
2 59145 1 6121
2 59146 1 6121
2 59147 1 6121
2 59148 1 6121
2 59149 1 6121
2 59150 1 6121
2 59151 1 6121
2 59152 1 6121
2 59153 1 6121
2 59154 1 6121
2 59155 1 6121
2 59156 1 6121
2 59157 1 6121
2 59158 1 6121
2 59159 1 6121
2 59160 1 6121
2 59161 1 6121
2 59162 1 6121
2 59163 1 6121
2 59164 1 6121
2 59165 1 6121
2 59166 1 6121
2 59167 1 6121
2 59168 1 6121
2 59169 1 6121
2 59170 1 6121
2 59171 1 6122
2 59172 1 6122
2 59173 1 6122
2 59174 1 6122
2 59175 1 6122
2 59176 1 6124
2 59177 1 6124
2 59178 1 6124
2 59179 1 6124
2 59180 1 6136
2 59181 1 6136
2 59182 1 6137
2 59183 1 6137
2 59184 1 6139
2 59185 1 6139
2 59186 1 6145
2 59187 1 6145
2 59188 1 6145
2 59189 1 6145
2 59190 1 6145
2 59191 1 6145
2 59192 1 6145
2 59193 1 6145
2 59194 1 6145
2 59195 1 6145
2 59196 1 6145
2 59197 1 6145
2 59198 1 6145
2 59199 1 6145
2 59200 1 6145
2 59201 1 6145
2 59202 1 6145
2 59203 1 6145
2 59204 1 6145
2 59205 1 6145
2 59206 1 6145
2 59207 1 6145
2 59208 1 6145
2 59209 1 6145
2 59210 1 6145
2 59211 1 6145
2 59212 1 6145
2 59213 1 6145
2 59214 1 6145
2 59215 1 6153
2 59216 1 6153
2 59217 1 6156
2 59218 1 6156
2 59219 1 6156
2 59220 1 6156
2 59221 1 6156
2 59222 1 6156
2 59223 1 6157
2 59224 1 6157
2 59225 1 6157
2 59226 1 6157
2 59227 1 6157
2 59228 1 6157
2 59229 1 6157
2 59230 1 6157
2 59231 1 6162
2 59232 1 6162
2 59233 1 6165
2 59234 1 6165
2 59235 1 6181
2 59236 1 6181
2 59237 1 6181
2 59238 1 6181
2 59239 1 6181
2 59240 1 6181
2 59241 1 6181
2 59242 1 6181
2 59243 1 6181
2 59244 1 6182
2 59245 1 6182
2 59246 1 6182
2 59247 1 6190
2 59248 1 6190
2 59249 1 6190
2 59250 1 6190
2 59251 1 6190
2 59252 1 6190
2 59253 1 6190
2 59254 1 6190
2 59255 1 6190
2 59256 1 6190
2 59257 1 6190
2 59258 1 6190
2 59259 1 6190
2 59260 1 6190
2 59261 1 6190
2 59262 1 6190
2 59263 1 6190
2 59264 1 6190
2 59265 1 6190
2 59266 1 6190
2 59267 1 6190
2 59268 1 6190
2 59269 1 6190
2 59270 1 6190
2 59271 1 6190
2 59272 1 6190
2 59273 1 6190
2 59274 1 6190
2 59275 1 6190
2 59276 1 6190
2 59277 1 6190
2 59278 1 6190
2 59279 1 6190
2 59280 1 6190
2 59281 1 6190
2 59282 1 6190
2 59283 1 6190
2 59284 1 6190
2 59285 1 6190
2 59286 1 6190
2 59287 1 6190
2 59288 1 6190
2 59289 1 6190
2 59290 1 6190
2 59291 1 6190
2 59292 1 6190
2 59293 1 6190
2 59294 1 6190
2 59295 1 6190
2 59296 1 6190
2 59297 1 6190
2 59298 1 6190
2 59299 1 6190
2 59300 1 6190
2 59301 1 6190
2 59302 1 6190
2 59303 1 6190
2 59304 1 6190
2 59305 1 6190
2 59306 1 6190
2 59307 1 6190
2 59308 1 6190
2 59309 1 6190
2 59310 1 6190
2 59311 1 6190
2 59312 1 6190
2 59313 1 6190
2 59314 1 6190
2 59315 1 6190
2 59316 1 6190
2 59317 1 6190
2 59318 1 6190
2 59319 1 6190
2 59320 1 6190
2 59321 1 6191
2 59322 1 6191
2 59323 1 6191
2 59324 1 6192
2 59325 1 6192
2 59326 1 6192
2 59327 1 6200
2 59328 1 6200
2 59329 1 6200
2 59330 1 6200
2 59331 1 6200
2 59332 1 6200
2 59333 1 6200
2 59334 1 6200
2 59335 1 6201
2 59336 1 6201
2 59337 1 6201
2 59338 1 6201
2 59339 1 6208
2 59340 1 6208
2 59341 1 6208
2 59342 1 6209
2 59343 1 6209
2 59344 1 6212
2 59345 1 6212
2 59346 1 6213
2 59347 1 6213
2 59348 1 6213
2 59349 1 6218
2 59350 1 6218
2 59351 1 6219
2 59352 1 6219
2 59353 1 6219
2 59354 1 6219
2 59355 1 6219
2 59356 1 6219
2 59357 1 6219
2 59358 1 6219
2 59359 1 6219
2 59360 1 6219
2 59361 1 6219
2 59362 1 6219
2 59363 1 6219
2 59364 1 6219
2 59365 1 6219
2 59366 1 6219
2 59367 1 6219
2 59368 1 6219
2 59369 1 6219
2 59370 1 6219
2 59371 1 6219
2 59372 1 6219
2 59373 1 6219
2 59374 1 6219
2 59375 1 6219
2 59376 1 6219
2 59377 1 6219
2 59378 1 6219
2 59379 1 6220
2 59380 1 6220
2 59381 1 6220
2 59382 1 6220
2 59383 1 6220
2 59384 1 6220
2 59385 1 6220
2 59386 1 6220
2 59387 1 6220
2 59388 1 6220
2 59389 1 6220
2 59390 1 6220
2 59391 1 6220
2 59392 1 6220
2 59393 1 6220
2 59394 1 6220
2 59395 1 6220
2 59396 1 6220
2 59397 1 6220
2 59398 1 6220
2 59399 1 6220
2 59400 1 6220
2 59401 1 6220
2 59402 1 6220
2 59403 1 6220
2 59404 1 6220
2 59405 1 6220
2 59406 1 6220
2 59407 1 6220
2 59408 1 6220
2 59409 1 6220
2 59410 1 6220
2 59411 1 6220
2 59412 1 6220
2 59413 1 6220
2 59414 1 6220
2 59415 1 6220
2 59416 1 6223
2 59417 1 6223
2 59418 1 6223
2 59419 1 6224
2 59420 1 6224
2 59421 1 6225
2 59422 1 6225
2 59423 1 6225
2 59424 1 6225
2 59425 1 6225
2 59426 1 6225
2 59427 1 6225
2 59428 1 6225
2 59429 1 6238
2 59430 1 6238
2 59431 1 6239
2 59432 1 6239
2 59433 1 6239
2 59434 1 6249
2 59435 1 6249
2 59436 1 6249
2 59437 1 6265
2 59438 1 6265
2 59439 1 6265
2 59440 1 6265
2 59441 1 6265
2 59442 1 6265
2 59443 1 6265
2 59444 1 6265
2 59445 1 6265
2 59446 1 6265
2 59447 1 6265
2 59448 1 6265
2 59449 1 6266
2 59450 1 6266
2 59451 1 6274
2 59452 1 6274
2 59453 1 6274
2 59454 1 6274
2 59455 1 6274
2 59456 1 6275
2 59457 1 6275
2 59458 1 6276
2 59459 1 6276
2 59460 1 6276
2 59461 1 6276
2 59462 1 6277
2 59463 1 6277
2 59464 1 6277
2 59465 1 6277
2 59466 1 6277
2 59467 1 6277
2 59468 1 6277
2 59469 1 6282
2 59470 1 6282
2 59471 1 6285
2 59472 1 6285
2 59473 1 6285
2 59474 1 6285
2 59475 1 6285
2 59476 1 6285
2 59477 1 6285
2 59478 1 6285
2 59479 1 6285
2 59480 1 6285
2 59481 1 6285
2 59482 1 6285
2 59483 1 6285
2 59484 1 6285
2 59485 1 6285
2 59486 1 6285
2 59487 1 6285
2 59488 1 6286
2 59489 1 6286
2 59490 1 6286
2 59491 1 6286
2 59492 1 6286
2 59493 1 6286
2 59494 1 6286
2 59495 1 6286
2 59496 1 6286
2 59497 1 6286
2 59498 1 6286
2 59499 1 6286
2 59500 1 6286
2 59501 1 6287
2 59502 1 6287
2 59503 1 6288
2 59504 1 6288
2 59505 1 6288
2 59506 1 6291
2 59507 1 6291
2 59508 1 6291
2 59509 1 6294
2 59510 1 6294
2 59511 1 6303
2 59512 1 6303
2 59513 1 6306
2 59514 1 6306
2 59515 1 6306
2 59516 1 6306
2 59517 1 6306
2 59518 1 6306
2 59519 1 6306
2 59520 1 6306
2 59521 1 6306
2 59522 1 6306
2 59523 1 6306
2 59524 1 6306
2 59525 1 6306
2 59526 1 6306
2 59527 1 6307
2 59528 1 6307
2 59529 1 6307
2 59530 1 6307
2 59531 1 6307
2 59532 1 6307
2 59533 1 6307
2 59534 1 6307
2 59535 1 6307
2 59536 1 6307
2 59537 1 6307
2 59538 1 6307
2 59539 1 6307
2 59540 1 6307
2 59541 1 6307
2 59542 1 6307
2 59543 1 6307
2 59544 1 6307
2 59545 1 6307
2 59546 1 6307
2 59547 1 6307
2 59548 1 6307
2 59549 1 6308
2 59550 1 6308
2 59551 1 6308
2 59552 1 6308
2 59553 1 6308
2 59554 1 6316
2 59555 1 6316
2 59556 1 6316
2 59557 1 6316
2 59558 1 6316
2 59559 1 6317
2 59560 1 6317
2 59561 1 6325
2 59562 1 6325
2 59563 1 6325
2 59564 1 6325
2 59565 1 6325
2 59566 1 6325
2 59567 1 6325
2 59568 1 6325
2 59569 1 6325
2 59570 1 6325
2 59571 1 6325
2 59572 1 6325
2 59573 1 6325
2 59574 1 6325
2 59575 1 6325
2 59576 1 6325
2 59577 1 6325
2 59578 1 6325
2 59579 1 6325
2 59580 1 6326
2 59581 1 6326
2 59582 1 6326
2 59583 1 6326
2 59584 1 6334
2 59585 1 6334
2 59586 1 6334
2 59587 1 6336
2 59588 1 6336
2 59589 1 6337
2 59590 1 6337
2 59591 1 6337
2 59592 1 6337
2 59593 1 6337
2 59594 1 6344
2 59595 1 6344
2 59596 1 6344
2 59597 1 6345
2 59598 1 6345
2 59599 1 6345
2 59600 1 6345
2 59601 1 6345
2 59602 1 6345
2 59603 1 6345
2 59604 1 6345
2 59605 1 6345
2 59606 1 6345
2 59607 1 6345
2 59608 1 6345
2 59609 1 6345
2 59610 1 6346
2 59611 1 6346
2 59612 1 6346
2 59613 1 6346
2 59614 1 6346
2 59615 1 6346
2 59616 1 6346
2 59617 1 6346
2 59618 1 6361
2 59619 1 6361
2 59620 1 6361
2 59621 1 6361
2 59622 1 6362
2 59623 1 6362
2 59624 1 6363
2 59625 1 6363
2 59626 1 6363
2 59627 1 6363
2 59628 1 6363
2 59629 1 6364
2 59630 1 6364
2 59631 1 6364
2 59632 1 6365
2 59633 1 6365
2 59634 1 6370
2 59635 1 6370
2 59636 1 6370
2 59637 1 6370
2 59638 1 6370
2 59639 1 6370
2 59640 1 6370
2 59641 1 6371
2 59642 1 6371
2 59643 1 6371
2 59644 1 6371
2 59645 1 6372
2 59646 1 6372
2 59647 1 6372
2 59648 1 6372
2 59649 1 6375
2 59650 1 6375
2 59651 1 6386
2 59652 1 6386
2 59653 1 6387
2 59654 1 6387
2 59655 1 6395
2 59656 1 6395
2 59657 1 6395
2 59658 1 6395
2 59659 1 6395
2 59660 1 6399
2 59661 1 6399
2 59662 1 6399
2 59663 1 6399
2 59664 1 6399
2 59665 1 6399
2 59666 1 6399
2 59667 1 6399
2 59668 1 6421
2 59669 1 6421
2 59670 1 6421
2 59671 1 6421
2 59672 1 6422
2 59673 1 6422
2 59674 1 6422
2 59675 1 6422
2 59676 1 6422
2 59677 1 6422
2 59678 1 6422
2 59679 1 6422
2 59680 1 6422
2 59681 1 6422
2 59682 1 6422
2 59683 1 6422
2 59684 1 6422
2 59685 1 6422
2 59686 1 6424
2 59687 1 6424
2 59688 1 6424
2 59689 1 6424
2 59690 1 6425
2 59691 1 6425
2 59692 1 6425
2 59693 1 6425
2 59694 1 6425
2 59695 1 6425
2 59696 1 6425
2 59697 1 6426
2 59698 1 6426
2 59699 1 6427
2 59700 1 6427
2 59701 1 6427
2 59702 1 6427
2 59703 1 6442
2 59704 1 6442
2 59705 1 6442
2 59706 1 6442
2 59707 1 6442
2 59708 1 6444
2 59709 1 6444
2 59710 1 6462
2 59711 1 6462
2 59712 1 6462
2 59713 1 6462
2 59714 1 6462
2 59715 1 6462
2 59716 1 6462
2 59717 1 6462
2 59718 1 6462
2 59719 1 6462
2 59720 1 6467
2 59721 1 6467
2 59722 1 6467
2 59723 1 6470
2 59724 1 6470
2 59725 1 6470
2 59726 1 6474
2 59727 1 6474
2 59728 1 6477
2 59729 1 6477
2 59730 1 6477
2 59731 1 6477
2 59732 1 6477
2 59733 1 6477
2 59734 1 6477
2 59735 1 6477
2 59736 1 6484
2 59737 1 6484
2 59738 1 6485
2 59739 1 6485
2 59740 1 6485
2 59741 1 6485
2 59742 1 6486
2 59743 1 6486
2 59744 1 6486
2 59745 1 6494
2 59746 1 6494
2 59747 1 6494
2 59748 1 6494
2 59749 1 6494
2 59750 1 6494
2 59751 1 6494
2 59752 1 6494
2 59753 1 6495
2 59754 1 6495
2 59755 1 6498
2 59756 1 6498
2 59757 1 6498
2 59758 1 6498
2 59759 1 6498
2 59760 1 6498
2 59761 1 6498
2 59762 1 6513
2 59763 1 6513
2 59764 1 6520
2 59765 1 6520
2 59766 1 6520
2 59767 1 6520
2 59768 1 6520
2 59769 1 6527
2 59770 1 6527
2 59771 1 6527
2 59772 1 6529
2 59773 1 6529
2 59774 1 6529
2 59775 1 6542
2 59776 1 6542
2 59777 1 6542
2 59778 1 6542
2 59779 1 6542
2 59780 1 6542
2 59781 1 6542
2 59782 1 6542
2 59783 1 6542
2 59784 1 6542
2 59785 1 6542
2 59786 1 6542
2 59787 1 6542
2 59788 1 6542
2 59789 1 6542
2 59790 1 6542
2 59791 1 6542
2 59792 1 6542
2 59793 1 6542
2 59794 1 6542
2 59795 1 6542
2 59796 1 6542
2 59797 1 6542
2 59798 1 6542
2 59799 1 6542
2 59800 1 6544
2 59801 1 6544
2 59802 1 6544
2 59803 1 6544
2 59804 1 6545
2 59805 1 6545
2 59806 1 6549
2 59807 1 6549
2 59808 1 6549
2 59809 1 6549
2 59810 1 6550
2 59811 1 6550
2 59812 1 6550
2 59813 1 6551
2 59814 1 6551
2 59815 1 6551
2 59816 1 6556
2 59817 1 6556
2 59818 1 6556
2 59819 1 6556
2 59820 1 6557
2 59821 1 6557
2 59822 1 6557
2 59823 1 6557
2 59824 1 6560
2 59825 1 6560
2 59826 1 6560
2 59827 1 6560
2 59828 1 6560
2 59829 1 6560
2 59830 1 6560
2 59831 1 6560
2 59832 1 6560
2 59833 1 6560
2 59834 1 6560
2 59835 1 6560
2 59836 1 6560
2 59837 1 6560
2 59838 1 6560
2 59839 1 6560
2 59840 1 6560
2 59841 1 6560
2 59842 1 6560
2 59843 1 6560
2 59844 1 6560
2 59845 1 6560
2 59846 1 6560
2 59847 1 6560
2 59848 1 6560
2 59849 1 6560
2 59850 1 6560
2 59851 1 6560
2 59852 1 6560
2 59853 1 6560
2 59854 1 6560
2 59855 1 6560
2 59856 1 6560
2 59857 1 6560
2 59858 1 6560
2 59859 1 6560
2 59860 1 6560
2 59861 1 6560
2 59862 1 6560
2 59863 1 6560
2 59864 1 6560
2 59865 1 6560
2 59866 1 6560
2 59867 1 6560
2 59868 1 6561
2 59869 1 6561
2 59870 1 6562
2 59871 1 6562
2 59872 1 6572
2 59873 1 6572
2 59874 1 6573
2 59875 1 6573
2 59876 1 6573
2 59877 1 6573
2 59878 1 6573
2 59879 1 6573
2 59880 1 6573
2 59881 1 6573
2 59882 1 6573
2 59883 1 6573
2 59884 1 6573
2 59885 1 6573
2 59886 1 6573
2 59887 1 6573
2 59888 1 6573
2 59889 1 6573
2 59890 1 6577
2 59891 1 6577
2 59892 1 6577
2 59893 1 6577
2 59894 1 6577
2 59895 1 6579
2 59896 1 6579
2 59897 1 6580
2 59898 1 6580
2 59899 1 6580
2 59900 1 6580
2 59901 1 6581
2 59902 1 6581
2 59903 1 6584
2 59904 1 6584
2 59905 1 6584
2 59906 1 6584
2 59907 1 6584
2 59908 1 6584
2 59909 1 6584
2 59910 1 6584
2 59911 1 6584
2 59912 1 6584
2 59913 1 6584
2 59914 1 6584
2 59915 1 6584
2 59916 1 6584
2 59917 1 6584
2 59918 1 6584
2 59919 1 6584
2 59920 1 6584
2 59921 1 6584
2 59922 1 6584
2 59923 1 6584
2 59924 1 6584
2 59925 1 6585
2 59926 1 6585
2 59927 1 6588
2 59928 1 6588
2 59929 1 6588
2 59930 1 6588
2 59931 1 6590
2 59932 1 6590
2 59933 1 6611
2 59934 1 6611
2 59935 1 6611
2 59936 1 6616
2 59937 1 6616
2 59938 1 6616
2 59939 1 6616
2 59940 1 6616
2 59941 1 6617
2 59942 1 6617
2 59943 1 6617
2 59944 1 6617
2 59945 1 6618
2 59946 1 6618
2 59947 1 6618
2 59948 1 6618
2 59949 1 6618
2 59950 1 6618
2 59951 1 6618
2 59952 1 6618
2 59953 1 6626
2 59954 1 6626
2 59955 1 6626
2 59956 1 6626
2 59957 1 6626
2 59958 1 6643
2 59959 1 6643
2 59960 1 6643
2 59961 1 6643
2 59962 1 6643
2 59963 1 6643
2 59964 1 6643
2 59965 1 6643
2 59966 1 6643
2 59967 1 6643
2 59968 1 6644
2 59969 1 6644
2 59970 1 6644
2 59971 1 6644
2 59972 1 6644
2 59973 1 6644
2 59974 1 6646
2 59975 1 6646
2 59976 1 6647
2 59977 1 6647
2 59978 1 6665
2 59979 1 6665
2 59980 1 6665
2 59981 1 6665
2 59982 1 6665
2 59983 1 6665
2 59984 1 6665
2 59985 1 6665
2 59986 1 6666
2 59987 1 6666
2 59988 1 6666
2 59989 1 6666
2 59990 1 6666
2 59991 1 6666
2 59992 1 6667
2 59993 1 6667
2 59994 1 6667
2 59995 1 6675
2 59996 1 6675
2 59997 1 6675
2 59998 1 6675
2 59999 1 6675
2 60000 1 6675
2 60001 1 6675
2 60002 1 6675
2 60003 1 6675
2 60004 1 6675
2 60005 1 6675
2 60006 1 6675
2 60007 1 6675
2 60008 1 6676
2 60009 1 6676
2 60010 1 6676
2 60011 1 6677
2 60012 1 6677
2 60013 1 6684
2 60014 1 6684
2 60015 1 6684
2 60016 1 6684
2 60017 1 6690
2 60018 1 6690
2 60019 1 6690
2 60020 1 6690
2 60021 1 6690
2 60022 1 6690
2 60023 1 6690
2 60024 1 6690
2 60025 1 6690
2 60026 1 6690
2 60027 1 6690
2 60028 1 6692
2 60029 1 6692
2 60030 1 6692
2 60031 1 6693
2 60032 1 6693
2 60033 1 6702
2 60034 1 6702
2 60035 1 6702
2 60036 1 6702
2 60037 1 6702
2 60038 1 6702
2 60039 1 6702
2 60040 1 6702
2 60041 1 6702
2 60042 1 6702
2 60043 1 6703
2 60044 1 6703
2 60045 1 6703
2 60046 1 6708
2 60047 1 6708
2 60048 1 6708
2 60049 1 6708
2 60050 1 6708
2 60051 1 6708
2 60052 1 6709
2 60053 1 6709
2 60054 1 6710
2 60055 1 6710
2 60056 1 6710
2 60057 1 6710
2 60058 1 6723
2 60059 1 6723
2 60060 1 6723
2 60061 1 6736
2 60062 1 6736
2 60063 1 6736
2 60064 1 6737
2 60065 1 6737
2 60066 1 6745
2 60067 1 6745
2 60068 1 6746
2 60069 1 6746
2 60070 1 6747
2 60071 1 6747
2 60072 1 6749
2 60073 1 6749
2 60074 1 6758
2 60075 1 6758
2 60076 1 6766
2 60077 1 6766
2 60078 1 6766
2 60079 1 6766
2 60080 1 6766
2 60081 1 6767
2 60082 1 6767
2 60083 1 6768
2 60084 1 6768
2 60085 1 6772
2 60086 1 6772
2 60087 1 6772
2 60088 1 6772
2 60089 1 6772
2 60090 1 6772
2 60091 1 6772
2 60092 1 6774
2 60093 1 6774
2 60094 1 6782
2 60095 1 6782
2 60096 1 6784
2 60097 1 6784
2 60098 1 6784
2 60099 1 6787
2 60100 1 6787
2 60101 1 6787
2 60102 1 6787
2 60103 1 6787
2 60104 1 6787
2 60105 1 6788
2 60106 1 6788
2 60107 1 6788
2 60108 1 6788
2 60109 1 6795
2 60110 1 6795
2 60111 1 6795
2 60112 1 6795
2 60113 1 6795
2 60114 1 6795
2 60115 1 6795
2 60116 1 6796
2 60117 1 6796
2 60118 1 6797
2 60119 1 6797
2 60120 1 6797
2 60121 1 6797
2 60122 1 6807
2 60123 1 6807
2 60124 1 6814
2 60125 1 6814
2 60126 1 6814
2 60127 1 6814
2 60128 1 6818
2 60129 1 6818
2 60130 1 6818
2 60131 1 6818
2 60132 1 6818
2 60133 1 6819
2 60134 1 6819
2 60135 1 6819
2 60136 1 6819
2 60137 1 6819
2 60138 1 6819
2 60139 1 6819
2 60140 1 6820
2 60141 1 6820
2 60142 1 6820
2 60143 1 6820
2 60144 1 6821
2 60145 1 6821
2 60146 1 6822
2 60147 1 6822
2 60148 1 6822
2 60149 1 6836
2 60150 1 6836
2 60151 1 6836
2 60152 1 6836
2 60153 1 6842
2 60154 1 6842
2 60155 1 6842
2 60156 1 6842
2 60157 1 6842
2 60158 1 6842
2 60159 1 6842
2 60160 1 6842
2 60161 1 6850
2 60162 1 6850
2 60163 1 6851
2 60164 1 6851
2 60165 1 6851
2 60166 1 6854
2 60167 1 6854
2 60168 1 6854
2 60169 1 6855
2 60170 1 6855
2 60171 1 6864
2 60172 1 6864
2 60173 1 6869
2 60174 1 6869
2 60175 1 6869
2 60176 1 6869
2 60177 1 6869
2 60178 1 6869
2 60179 1 6869
2 60180 1 6869
2 60181 1 6869
2 60182 1 6869
2 60183 1 6869
2 60184 1 6869
2 60185 1 6869
2 60186 1 6869
2 60187 1 6869
2 60188 1 6869
2 60189 1 6870
2 60190 1 6870
2 60191 1 6870
2 60192 1 6886
2 60193 1 6886
2 60194 1 6886
2 60195 1 6888
2 60196 1 6888
2 60197 1 6888
2 60198 1 6888
2 60199 1 6897
2 60200 1 6897
2 60201 1 6898
2 60202 1 6898
2 60203 1 6898
2 60204 1 6899
2 60205 1 6899
2 60206 1 6899
2 60207 1 6899
2 60208 1 6900
2 60209 1 6900
2 60210 1 6900
2 60211 1 6901
2 60212 1 6901
2 60213 1 6901
2 60214 1 6901
2 60215 1 6902
2 60216 1 6902
2 60217 1 6902
2 60218 1 6902
2 60219 1 6902
2 60220 1 6903
2 60221 1 6903
2 60222 1 6903
2 60223 1 6906
2 60224 1 6906
2 60225 1 6913
2 60226 1 6913
2 60227 1 6913
2 60228 1 6913
2 60229 1 6913
2 60230 1 6913
2 60231 1 6913
2 60232 1 6913
2 60233 1 6913
2 60234 1 6913
2 60235 1 6913
2 60236 1 6913
2 60237 1 6914
2 60238 1 6914
2 60239 1 6927
2 60240 1 6927
2 60241 1 6948
2 60242 1 6948
2 60243 1 6948
2 60244 1 6950
2 60245 1 6950
2 60246 1 6950
2 60247 1 6950
2 60248 1 6959
2 60249 1 6959
2 60250 1 6959
2 60251 1 6971
2 60252 1 6971
2 60253 1 6971
2 60254 1 6971
2 60255 1 6987
2 60256 1 6987
2 60257 1 7007
2 60258 1 7007
2 60259 1 7007
2 60260 1 7007
2 60261 1 7007
2 60262 1 7007
2 60263 1 7027
2 60264 1 7027
2 60265 1 7027
2 60266 1 7027
2 60267 1 7027
2 60268 1 7027
2 60269 1 7027
2 60270 1 7028
2 60271 1 7028
2 60272 1 7028
2 60273 1 7028
2 60274 1 7028
2 60275 1 7028
2 60276 1 7028
2 60277 1 7028
2 60278 1 7028
2 60279 1 7028
2 60280 1 7028
2 60281 1 7028
2 60282 1 7028
2 60283 1 7028
2 60284 1 7028
2 60285 1 7028
2 60286 1 7028
2 60287 1 7028
2 60288 1 7028
2 60289 1 7028
2 60290 1 7028
2 60291 1 7028
2 60292 1 7028
2 60293 1 7028
2 60294 1 7028
2 60295 1 7028
2 60296 1 7028
2 60297 1 7028
2 60298 1 7028
2 60299 1 7036
2 60300 1 7036
2 60301 1 7036
2 60302 1 7036
2 60303 1 7036
2 60304 1 7036
2 60305 1 7036
2 60306 1 7036
2 60307 1 7036
2 60308 1 7036
2 60309 1 7036
2 60310 1 7036
2 60311 1 7036
2 60312 1 7036
2 60313 1 7036
2 60314 1 7037
2 60315 1 7037
2 60316 1 7038
2 60317 1 7038
2 60318 1 7038
2 60319 1 7038
2 60320 1 7038
2 60321 1 7038
2 60322 1 7038
2 60323 1 7038
2 60324 1 7038
2 60325 1 7038
2 60326 1 7040
2 60327 1 7040
2 60328 1 7040
2 60329 1 7040
2 60330 1 7040
2 60331 1 7040
2 60332 1 7040
2 60333 1 7040
2 60334 1 7040
2 60335 1 7040
2 60336 1 7040
2 60337 1 7040
2 60338 1 7040
2 60339 1 7040
2 60340 1 7040
2 60341 1 7043
2 60342 1 7043
2 60343 1 7043
2 60344 1 7043
2 60345 1 7043
2 60346 1 7043
2 60347 1 7043
2 60348 1 7043
2 60349 1 7043
2 60350 1 7043
2 60351 1 7043
2 60352 1 7043
2 60353 1 7043
2 60354 1 7043
2 60355 1 7043
2 60356 1 7043
2 60357 1 7043
2 60358 1 7043
2 60359 1 7043
2 60360 1 7043
2 60361 1 7043
2 60362 1 7043
2 60363 1 7043
2 60364 1 7043
2 60365 1 7043
2 60366 1 7043
2 60367 1 7043
2 60368 1 7043
2 60369 1 7043
2 60370 1 7043
2 60371 1 7043
2 60372 1 7043
2 60373 1 7043
2 60374 1 7043
2 60375 1 7043
2 60376 1 7043
2 60377 1 7043
2 60378 1 7043
2 60379 1 7043
2 60380 1 7043
2 60381 1 7043
2 60382 1 7043
2 60383 1 7043
2 60384 1 7043
2 60385 1 7043
2 60386 1 7043
2 60387 1 7043
2 60388 1 7043
2 60389 1 7043
2 60390 1 7043
2 60391 1 7043
2 60392 1 7043
2 60393 1 7043
2 60394 1 7043
2 60395 1 7043
2 60396 1 7043
2 60397 1 7043
2 60398 1 7043
2 60399 1 7043
2 60400 1 7043
2 60401 1 7043
2 60402 1 7043
2 60403 1 7043
2 60404 1 7043
2 60405 1 7043
2 60406 1 7043
2 60407 1 7043
2 60408 1 7043
2 60409 1 7043
2 60410 1 7043
2 60411 1 7051
2 60412 1 7051
2 60413 1 7051
2 60414 1 7051
2 60415 1 7051
2 60416 1 7051
2 60417 1 7051
2 60418 1 7051
2 60419 1 7052
2 60420 1 7052
2 60421 1 7052
2 60422 1 7052
2 60423 1 7052
2 60424 1 7052
2 60425 1 7052
2 60426 1 7052
2 60427 1 7054
2 60428 1 7054
2 60429 1 7062
2 60430 1 7062
2 60431 1 7062
2 60432 1 7062
2 60433 1 7063
2 60434 1 7063
2 60435 1 7063
2 60436 1 7063
2 60437 1 7072
2 60438 1 7072
2 60439 1 7072
2 60440 1 7074
2 60441 1 7074
2 60442 1 7075
2 60443 1 7075
2 60444 1 7075
2 60445 1 7075
2 60446 1 7075
2 60447 1 7075
2 60448 1 7075
2 60449 1 7075
2 60450 1 7075
2 60451 1 7075
2 60452 1 7075
2 60453 1 7075
2 60454 1 7075
2 60455 1 7075
2 60456 1 7075
2 60457 1 7075
2 60458 1 7075
2 60459 1 7075
2 60460 1 7075
2 60461 1 7075
2 60462 1 7075
2 60463 1 7075
2 60464 1 7075
2 60465 1 7075
2 60466 1 7075
2 60467 1 7075
2 60468 1 7075
2 60469 1 7075
2 60470 1 7075
2 60471 1 7075
2 60472 1 7075
2 60473 1 7075
2 60474 1 7075
2 60475 1 7075
2 60476 1 7075
2 60477 1 7075
2 60478 1 7075
2 60479 1 7075
2 60480 1 7075
2 60481 1 7075
2 60482 1 7075
2 60483 1 7083
2 60484 1 7083
2 60485 1 7085
2 60486 1 7085
2 60487 1 7085
2 60488 1 7085
2 60489 1 7086
2 60490 1 7086
2 60491 1 7086
2 60492 1 7086
2 60493 1 7094
2 60494 1 7094
2 60495 1 7094
2 60496 1 7094
2 60497 1 7094
2 60498 1 7094
2 60499 1 7094
2 60500 1 7095
2 60501 1 7095
2 60502 1 7095
2 60503 1 7095
2 60504 1 7095
2 60505 1 7096
2 60506 1 7096
2 60507 1 7103
2 60508 1 7103
2 60509 1 7103
2 60510 1 7103
2 60511 1 7103
2 60512 1 7103
2 60513 1 7110
2 60514 1 7110
2 60515 1 7118
2 60516 1 7118
2 60517 1 7118
2 60518 1 7118
2 60519 1 7118
2 60520 1 7118
2 60521 1 7118
2 60522 1 7118
2 60523 1 7119
2 60524 1 7119
2 60525 1 7119
2 60526 1 7119
2 60527 1 7119
2 60528 1 7119
2 60529 1 7119
2 60530 1 7119
2 60531 1 7119
2 60532 1 7119
2 60533 1 7119
2 60534 1 7119
2 60535 1 7119
2 60536 1 7119
2 60537 1 7119
2 60538 1 7119
2 60539 1 7119
2 60540 1 7119
2 60541 1 7119
2 60542 1 7119
2 60543 1 7119
2 60544 1 7119
2 60545 1 7119
2 60546 1 7119
2 60547 1 7119
2 60548 1 7119
2 60549 1 7119
2 60550 1 7119
2 60551 1 7119
2 60552 1 7119
2 60553 1 7119
2 60554 1 7128
2 60555 1 7128
2 60556 1 7136
2 60557 1 7136
2 60558 1 7136
2 60559 1 7136
2 60560 1 7136
2 60561 1 7136
2 60562 1 7136
2 60563 1 7136
2 60564 1 7136
2 60565 1 7136
2 60566 1 7136
2 60567 1 7136
2 60568 1 7136
2 60569 1 7136
2 60570 1 7136
2 60571 1 7136
2 60572 1 7136
2 60573 1 7136
2 60574 1 7136
2 60575 1 7136
2 60576 1 7138
2 60577 1 7138
2 60578 1 7138
2 60579 1 7138
2 60580 1 7138
2 60581 1 7139
2 60582 1 7139
2 60583 1 7142
2 60584 1 7142
2 60585 1 7142
2 60586 1 7145
2 60587 1 7145
2 60588 1 7145
2 60589 1 7147
2 60590 1 7147
2 60591 1 7153
2 60592 1 7153
2 60593 1 7153
2 60594 1 7153
2 60595 1 7161
2 60596 1 7161
2 60597 1 7162
2 60598 1 7162
2 60599 1 7162
2 60600 1 7162
2 60601 1 7163
2 60602 1 7163
2 60603 1 7164
2 60604 1 7164
2 60605 1 7169
2 60606 1 7169
2 60607 1 7169
2 60608 1 7169
2 60609 1 7170
2 60610 1 7170
2 60611 1 7170
2 60612 1 7170
2 60613 1 7170
2 60614 1 7170
2 60615 1 7170
2 60616 1 7170
2 60617 1 7170
2 60618 1 7187
2 60619 1 7187
2 60620 1 7187
2 60621 1 7187
2 60622 1 7187
2 60623 1 7187
2 60624 1 7187
2 60625 1 7187
2 60626 1 7187
2 60627 1 7187
2 60628 1 7187
2 60629 1 7187
2 60630 1 7187
2 60631 1 7187
2 60632 1 7187
2 60633 1 7187
2 60634 1 7187
2 60635 1 7187
2 60636 1 7187
2 60637 1 7187
2 60638 1 7187
2 60639 1 7187
2 60640 1 7187
2 60641 1 7187
2 60642 1 7187
2 60643 1 7187
2 60644 1 7187
2 60645 1 7187
2 60646 1 7187
2 60647 1 7187
2 60648 1 7187
2 60649 1 7187
2 60650 1 7187
2 60651 1 7187
2 60652 1 7187
2 60653 1 7187
2 60654 1 7187
2 60655 1 7187
2 60656 1 7188
2 60657 1 7188
2 60658 1 7188
2 60659 1 7188
2 60660 1 7188
2 60661 1 7188
2 60662 1 7188
2 60663 1 7189
2 60664 1 7189
2 60665 1 7189
2 60666 1 7200
2 60667 1 7200
2 60668 1 7200
2 60669 1 7200
2 60670 1 7200
2 60671 1 7200
2 60672 1 7200
2 60673 1 7200
2 60674 1 7200
2 60675 1 7200
2 60676 1 7200
2 60677 1 7200
2 60678 1 7200
2 60679 1 7200
2 60680 1 7200
2 60681 1 7200
2 60682 1 7201
2 60683 1 7201
2 60684 1 7201
2 60685 1 7201
2 60686 1 7202
2 60687 1 7202
2 60688 1 7202
2 60689 1 7202
2 60690 1 7203
2 60691 1 7203
2 60692 1 7210
2 60693 1 7210
2 60694 1 7210
2 60695 1 7211
2 60696 1 7211
2 60697 1 7212
2 60698 1 7212
2 60699 1 7225
2 60700 1 7225
2 60701 1 7225
2 60702 1 7225
2 60703 1 7225
2 60704 1 7225
2 60705 1 7225
2 60706 1 7225
2 60707 1 7226
2 60708 1 7226
2 60709 1 7226
2 60710 1 7228
2 60711 1 7228
2 60712 1 7228
2 60713 1 7228
2 60714 1 7228
2 60715 1 7228
2 60716 1 7228
2 60717 1 7229
2 60718 1 7229
2 60719 1 7229
2 60720 1 7229
2 60721 1 7229
2 60722 1 7229
2 60723 1 7230
2 60724 1 7230
2 60725 1 7232
2 60726 1 7232
2 60727 1 7232
2 60728 1 7232
2 60729 1 7233
2 60730 1 7233
2 60731 1 7237
2 60732 1 7237
2 60733 1 7238
2 60734 1 7238
2 60735 1 7257
2 60736 1 7257
2 60737 1 7257
2 60738 1 7257
2 60739 1 7257
2 60740 1 7257
2 60741 1 7257
2 60742 1 7257
2 60743 1 7257
2 60744 1 7257
2 60745 1 7258
2 60746 1 7258
2 60747 1 7258
2 60748 1 7258
2 60749 1 7258
2 60750 1 7258
2 60751 1 7258
2 60752 1 7258
2 60753 1 7258
2 60754 1 7258
2 60755 1 7259
2 60756 1 7259
2 60757 1 7259
2 60758 1 7260
2 60759 1 7260
2 60760 1 7260
2 60761 1 7260
2 60762 1 7260
2 60763 1 7260
2 60764 1 7260
2 60765 1 7262
2 60766 1 7262
2 60767 1 7262
2 60768 1 7262
2 60769 1 7263
2 60770 1 7263
2 60771 1 7277
2 60772 1 7277
2 60773 1 7278
2 60774 1 7278
2 60775 1 7278
2 60776 1 7278
2 60777 1 7278
2 60778 1 7278
2 60779 1 7279
2 60780 1 7279
2 60781 1 7287
2 60782 1 7287
2 60783 1 7287
2 60784 1 7290
2 60785 1 7290
2 60786 1 7290
2 60787 1 7290
2 60788 1 7290
2 60789 1 7291
2 60790 1 7291
2 60791 1 7291
2 60792 1 7291
2 60793 1 7291
2 60794 1 7291
2 60795 1 7291
2 60796 1 7291
2 60797 1 7291
2 60798 1 7292
2 60799 1 7292
2 60800 1 7292
2 60801 1 7293
2 60802 1 7293
2 60803 1 7293
2 60804 1 7293
2 60805 1 7293
2 60806 1 7293
2 60807 1 7300
2 60808 1 7300
2 60809 1 7300
2 60810 1 7300
2 60811 1 7300
2 60812 1 7300
2 60813 1 7301
2 60814 1 7301
2 60815 1 7303
2 60816 1 7303
2 60817 1 7303
2 60818 1 7303
2 60819 1 7303
2 60820 1 7303
2 60821 1 7303
2 60822 1 7303
2 60823 1 7303
2 60824 1 7320
2 60825 1 7320
2 60826 1 7330
2 60827 1 7330
2 60828 1 7331
2 60829 1 7331
2 60830 1 7331
2 60831 1 7332
2 60832 1 7332
2 60833 1 7333
2 60834 1 7333
2 60835 1 7333
2 60836 1 7338
2 60837 1 7338
2 60838 1 7352
2 60839 1 7352
2 60840 1 7352
2 60841 1 7353
2 60842 1 7353
2 60843 1 7353
2 60844 1 7353
2 60845 1 7354
2 60846 1 7354
2 60847 1 7354
2 60848 1 7358
2 60849 1 7358
2 60850 1 7358
2 60851 1 7359
2 60852 1 7359
2 60853 1 7359
2 60854 1 7366
2 60855 1 7366
2 60856 1 7366
2 60857 1 7366
2 60858 1 7379
2 60859 1 7379
2 60860 1 7379
2 60861 1 7379
2 60862 1 7380
2 60863 1 7380
2 60864 1 7392
2 60865 1 7392
2 60866 1 7393
2 60867 1 7393
2 60868 1 7393
2 60869 1 7405
2 60870 1 7405
2 60871 1 7410
2 60872 1 7410
2 60873 1 7411
2 60874 1 7411
2 60875 1 7411
2 60876 1 7419
2 60877 1 7419
2 60878 1 7419
2 60879 1 7426
2 60880 1 7426
2 60881 1 7427
2 60882 1 7427
2 60883 1 7428
2 60884 1 7428
2 60885 1 7428
2 60886 1 7437
2 60887 1 7437
2 60888 1 7437
2 60889 1 7437
2 60890 1 7437
2 60891 1 7437
2 60892 1 7437
2 60893 1 7437
2 60894 1 7438
2 60895 1 7438
2 60896 1 7438
2 60897 1 7438
2 60898 1 7438
2 60899 1 7438
2 60900 1 7438
2 60901 1 7439
2 60902 1 7439
2 60903 1 7441
2 60904 1 7441
2 60905 1 7444
2 60906 1 7444
2 60907 1 7444
2 60908 1 7444
2 60909 1 7444
2 60910 1 7444
2 60911 1 7460
2 60912 1 7460
2 60913 1 7460
2 60914 1 7460
2 60915 1 7460
2 60916 1 7460
2 60917 1 7460
2 60918 1 7460
2 60919 1 7461
2 60920 1 7461
2 60921 1 7462
2 60922 1 7462
2 60923 1 7462
2 60924 1 7462
2 60925 1 7462
2 60926 1 7462
2 60927 1 7462
2 60928 1 7462
2 60929 1 7462
2 60930 1 7462
2 60931 1 7478
2 60932 1 7478
2 60933 1 7478
2 60934 1 7478
2 60935 1 7478
2 60936 1 7478
2 60937 1 7479
2 60938 1 7479
2 60939 1 7479
2 60940 1 7480
2 60941 1 7480
2 60942 1 7480
2 60943 1 7483
2 60944 1 7483
2 60945 1 7484
2 60946 1 7484
2 60947 1 7484
2 60948 1 7484
2 60949 1 7484
2 60950 1 7485
2 60951 1 7485
2 60952 1 7486
2 60953 1 7486
2 60954 1 7486
2 60955 1 7486
2 60956 1 7486
2 60957 1 7487
2 60958 1 7487
2 60959 1 7487
2 60960 1 7487
2 60961 1 7487
2 60962 1 7487
2 60963 1 7491
2 60964 1 7491
2 60965 1 7491
2 60966 1 7491
2 60967 1 7491
2 60968 1 7491
2 60969 1 7501
2 60970 1 7501
2 60971 1 7501
2 60972 1 7501
2 60973 1 7501
2 60974 1 7501
2 60975 1 7501
2 60976 1 7501
2 60977 1 7501
2 60978 1 7501
2 60979 1 7501
2 60980 1 7501
2 60981 1 7501
2 60982 1 7501
2 60983 1 7501
2 60984 1 7501
2 60985 1 7501
2 60986 1 7501
2 60987 1 7501
2 60988 1 7501
2 60989 1 7501
2 60990 1 7501
2 60991 1 7501
2 60992 1 7501
2 60993 1 7501
2 60994 1 7502
2 60995 1 7502
2 60996 1 7502
2 60997 1 7502
2 60998 1 7502
2 60999 1 7502
2 61000 1 7505
2 61001 1 7505
2 61002 1 7505
2 61003 1 7505
2 61004 1 7507
2 61005 1 7507
2 61006 1 7507
2 61007 1 7507
2 61008 1 7507
2 61009 1 7507
2 61010 1 7507
2 61011 1 7508
2 61012 1 7508
2 61013 1 7509
2 61014 1 7509
2 61015 1 7509
2 61016 1 7509
2 61017 1 7509
2 61018 1 7509
2 61019 1 7509
2 61020 1 7509
2 61021 1 7509
2 61022 1 7509
2 61023 1 7509
2 61024 1 7509
2 61025 1 7509
2 61026 1 7509
2 61027 1 7509
2 61028 1 7509
2 61029 1 7509
2 61030 1 7509
2 61031 1 7510
2 61032 1 7510
2 61033 1 7510
2 61034 1 7518
2 61035 1 7518
2 61036 1 7518
2 61037 1 7518
2 61038 1 7518
2 61039 1 7519
2 61040 1 7519
2 61041 1 7519
2 61042 1 7519
2 61043 1 7519
2 61044 1 7519
2 61045 1 7519
2 61046 1 7519
2 61047 1 7519
2 61048 1 7519
2 61049 1 7519
2 61050 1 7519
2 61051 1 7519
2 61052 1 7519
2 61053 1 7519
2 61054 1 7519
2 61055 1 7519
2 61056 1 7519
2 61057 1 7519
2 61058 1 7519
2 61059 1 7521
2 61060 1 7521
2 61061 1 7521
2 61062 1 7521
2 61063 1 7521
2 61064 1 7522
2 61065 1 7522
2 61066 1 7522
2 61067 1 7528
2 61068 1 7528
2 61069 1 7528
2 61070 1 7528
2 61071 1 7528
2 61072 1 7529
2 61073 1 7529
2 61074 1 7529
2 61075 1 7530
2 61076 1 7530
2 61077 1 7535
2 61078 1 7535
2 61079 1 7535
2 61080 1 7535
2 61081 1 7535
2 61082 1 7535
2 61083 1 7535
2 61084 1 7535
2 61085 1 7535
2 61086 1 7535
2 61087 1 7536
2 61088 1 7536
2 61089 1 7536
2 61090 1 7536
2 61091 1 7540
2 61092 1 7540
2 61093 1 7540
2 61094 1 7540
2 61095 1 7540
2 61096 1 7540
2 61097 1 7540
2 61098 1 7540
2 61099 1 7540
2 61100 1 7541
2 61101 1 7541
2 61102 1 7541
2 61103 1 7541
2 61104 1 7550
2 61105 1 7550
2 61106 1 7550
2 61107 1 7550
2 61108 1 7559
2 61109 1 7559
2 61110 1 7559
2 61111 1 7559
2 61112 1 7559
2 61113 1 7559
2 61114 1 7575
2 61115 1 7575
2 61116 1 7599
2 61117 1 7599
2 61118 1 7599
2 61119 1 7599
2 61120 1 7599
2 61121 1 7599
2 61122 1 7599
2 61123 1 7599
2 61124 1 7599
2 61125 1 7599
2 61126 1 7599
2 61127 1 7599
2 61128 1 7599
2 61129 1 7599
2 61130 1 7599
2 61131 1 7599
2 61132 1 7599
2 61133 1 7599
2 61134 1 7599
2 61135 1 7599
2 61136 1 7599
2 61137 1 7599
2 61138 1 7599
2 61139 1 7599
2 61140 1 7599
2 61141 1 7599
2 61142 1 7599
2 61143 1 7599
2 61144 1 7599
2 61145 1 7599
2 61146 1 7599
2 61147 1 7599
2 61148 1 7599
2 61149 1 7599
2 61150 1 7599
2 61151 1 7599
2 61152 1 7599
2 61153 1 7599
2 61154 1 7599
2 61155 1 7599
2 61156 1 7599
2 61157 1 7599
2 61158 1 7599
2 61159 1 7599
2 61160 1 7599
2 61161 1 7599
2 61162 1 7599
2 61163 1 7599
2 61164 1 7599
2 61165 1 7599
2 61166 1 7599
2 61167 1 7599
2 61168 1 7599
2 61169 1 7599
2 61170 1 7599
2 61171 1 7599
2 61172 1 7599
2 61173 1 7599
2 61174 1 7599
2 61175 1 7600
2 61176 1 7600
2 61177 1 7601
2 61178 1 7601
2 61179 1 7601
2 61180 1 7601
2 61181 1 7601
2 61182 1 7601
2 61183 1 7601
2 61184 1 7601
2 61185 1 7601
2 61186 1 7601
2 61187 1 7601
2 61188 1 7601
2 61189 1 7601
2 61190 1 7601
2 61191 1 7601
2 61192 1 7601
2 61193 1 7601
2 61194 1 7601
2 61195 1 7601
2 61196 1 7601
2 61197 1 7601
2 61198 1 7601
2 61199 1 7601
2 61200 1 7612
2 61201 1 7612
2 61202 1 7613
2 61203 1 7613
2 61204 1 7613
2 61205 1 7613
2 61206 1 7613
2 61207 1 7613
2 61208 1 7613
2 61209 1 7621
2 61210 1 7621
2 61211 1 7626
2 61212 1 7626
2 61213 1 7627
2 61214 1 7627
2 61215 1 7627
2 61216 1 7628
2 61217 1 7628
2 61218 1 7628
2 61219 1 7628
2 61220 1 7630
2 61221 1 7630
2 61222 1 7633
2 61223 1 7633
2 61224 1 7633
2 61225 1 7637
2 61226 1 7637
2 61227 1 7637
2 61228 1 7640
2 61229 1 7640
2 61230 1 7640
2 61231 1 7640
2 61232 1 7640
2 61233 1 7640
2 61234 1 7640
2 61235 1 7640
2 61236 1 7641
2 61237 1 7641
2 61238 1 7648
2 61239 1 7648
2 61240 1 7648
2 61241 1 7650
2 61242 1 7650
2 61243 1 7651
2 61244 1 7651
2 61245 1 7651
2 61246 1 7651
2 61247 1 7651
2 61248 1 7653
2 61249 1 7653
2 61250 1 7662
2 61251 1 7662
2 61252 1 7662
2 61253 1 7662
2 61254 1 7662
2 61255 1 7662
2 61256 1 7670
2 61257 1 7670
2 61258 1 7670
2 61259 1 7670
2 61260 1 7671
2 61261 1 7671
2 61262 1 7671
2 61263 1 7671
2 61264 1 7671
2 61265 1 7671
2 61266 1 7671
2 61267 1 7671
2 61268 1 7671
2 61269 1 7671
2 61270 1 7671
2 61271 1 7671
2 61272 1 7671
2 61273 1 7671
2 61274 1 7671
2 61275 1 7671
2 61276 1 7671
2 61277 1 7671
2 61278 1 7672
2 61279 1 7672
2 61280 1 7672
2 61281 1 7672
2 61282 1 7677
2 61283 1 7677
2 61284 1 7678
2 61285 1 7678
2 61286 1 7678
2 61287 1 7679
2 61288 1 7679
2 61289 1 7679
2 61290 1 7679
2 61291 1 7679
2 61292 1 7679
2 61293 1 7679
2 61294 1 7694
2 61295 1 7694
2 61296 1 7717
2 61297 1 7717
2 61298 1 7718
2 61299 1 7718
2 61300 1 7718
2 61301 1 7719
2 61302 1 7719
2 61303 1 7719
2 61304 1 7719
2 61305 1 7719
2 61306 1 7719
2 61307 1 7723
2 61308 1 7723
2 61309 1 7723
2 61310 1 7723
2 61311 1 7723
2 61312 1 7723
2 61313 1 7723
2 61314 1 7723
2 61315 1 7723
2 61316 1 7723
2 61317 1 7723
2 61318 1 7723
2 61319 1 7723
2 61320 1 7723
2 61321 1 7725
2 61322 1 7725
2 61323 1 7725
2 61324 1 7725
2 61325 1 7725
2 61326 1 7725
2 61327 1 7729
2 61328 1 7729
2 61329 1 7732
2 61330 1 7732
2 61331 1 7732
2 61332 1 7736
2 61333 1 7736
2 61334 1 7736
2 61335 1 7736
2 61336 1 7736
2 61337 1 7745
2 61338 1 7745
2 61339 1 7745
2 61340 1 7745
2 61341 1 7745
2 61342 1 7745
2 61343 1 7745
2 61344 1 7745
2 61345 1 7745
2 61346 1 7745
2 61347 1 7745
2 61348 1 7745
2 61349 1 7745
2 61350 1 7745
2 61351 1 7745
2 61352 1 7745
2 61353 1 7746
2 61354 1 7746
2 61355 1 7746
2 61356 1 7747
2 61357 1 7747
2 61358 1 7747
2 61359 1 7747
2 61360 1 7747
2 61361 1 7747
2 61362 1 7756
2 61363 1 7756
2 61364 1 7764
2 61365 1 7764
2 61366 1 7764
2 61367 1 7765
2 61368 1 7765
2 61369 1 7765
2 61370 1 7765
2 61371 1 7765
2 61372 1 7765
2 61373 1 7765
2 61374 1 7765
2 61375 1 7765
2 61376 1 7765
2 61377 1 7765
2 61378 1 7765
2 61379 1 7765
2 61380 1 7765
2 61381 1 7765
2 61382 1 7765
2 61383 1 7765
2 61384 1 7768
2 61385 1 7768
2 61386 1 7772
2 61387 1 7772
2 61388 1 7772
2 61389 1 7786
2 61390 1 7786
2 61391 1 7786
2 61392 1 7786
2 61393 1 7786
2 61394 1 7786
2 61395 1 7786
2 61396 1 7786
2 61397 1 7786
2 61398 1 7787
2 61399 1 7787
2 61400 1 7787
2 61401 1 7787
2 61402 1 7790
2 61403 1 7790
2 61404 1 7790
2 61405 1 7790
2 61406 1 7790
2 61407 1 7793
2 61408 1 7793
2 61409 1 7793
2 61410 1 7793
2 61411 1 7794
2 61412 1 7794
2 61413 1 7819
2 61414 1 7819
2 61415 1 7819
2 61416 1 7819
2 61417 1 7819
2 61418 1 7820
2 61419 1 7820
2 61420 1 7820
2 61421 1 7820
2 61422 1 7834
2 61423 1 7834
2 61424 1 7834
2 61425 1 7835
2 61426 1 7835
2 61427 1 7840
2 61428 1 7840
2 61429 1 7840
2 61430 1 7840
2 61431 1 7840
2 61432 1 7840
2 61433 1 7840
2 61434 1 7840
2 61435 1 7840
2 61436 1 7840
2 61437 1 7840
2 61438 1 7840
2 61439 1 7840
2 61440 1 7840
2 61441 1 7840
2 61442 1 7840
2 61443 1 7841
2 61444 1 7841
2 61445 1 7841
2 61446 1 7845
2 61447 1 7845
2 61448 1 7845
2 61449 1 7845
2 61450 1 7845
2 61451 1 7845
2 61452 1 7845
2 61453 1 7845
2 61454 1 7845
2 61455 1 7845
2 61456 1 7845
2 61457 1 7845
2 61458 1 7845
2 61459 1 7846
2 61460 1 7846
2 61461 1 7846
2 61462 1 7846
2 61463 1 7846
2 61464 1 7846
2 61465 1 7846
2 61466 1 7846
2 61467 1 7846
2 61468 1 7846
2 61469 1 7847
2 61470 1 7847
2 61471 1 7856
2 61472 1 7856
2 61473 1 7857
2 61474 1 7857
2 61475 1 7865
2 61476 1 7865
2 61477 1 7865
2 61478 1 7866
2 61479 1 7866
2 61480 1 7866
2 61481 1 7866
2 61482 1 7877
2 61483 1 7877
2 61484 1 7877
2 61485 1 7877
2 61486 1 7877
2 61487 1 7877
2 61488 1 7885
2 61489 1 7885
2 61490 1 7885
2 61491 1 7886
2 61492 1 7886
2 61493 1 7902
2 61494 1 7902
2 61495 1 7902
2 61496 1 7904
2 61497 1 7904
2 61498 1 7906
2 61499 1 7906
2 61500 1 7906
2 61501 1 7912
2 61502 1 7912
2 61503 1 7912
2 61504 1 7917
2 61505 1 7917
2 61506 1 7917
2 61507 1 7917
2 61508 1 7917
2 61509 1 7917
2 61510 1 7918
2 61511 1 7918
2 61512 1 7918
2 61513 1 7918
2 61514 1 7918
2 61515 1 7918
2 61516 1 7918
2 61517 1 7918
2 61518 1 7918
2 61519 1 7918
2 61520 1 7918
2 61521 1 7919
2 61522 1 7919
2 61523 1 7919
2 61524 1 7919
2 61525 1 7919
2 61526 1 7919
2 61527 1 7919
2 61528 1 7919
2 61529 1 7919
2 61530 1 7919
2 61531 1 7919
2 61532 1 7919
2 61533 1 7929
2 61534 1 7929
2 61535 1 7930
2 61536 1 7930
2 61537 1 7931
2 61538 1 7931
2 61539 1 7932
2 61540 1 7932
2 61541 1 7934
2 61542 1 7934
2 61543 1 7935
2 61544 1 7935
2 61545 1 7938
2 61546 1 7938
2 61547 1 7938
2 61548 1 7958
2 61549 1 7958
2 61550 1 7959
2 61551 1 7959
2 61552 1 7962
2 61553 1 7962
2 61554 1 7962
2 61555 1 7963
2 61556 1 7963
2 61557 1 7963
2 61558 1 7963
2 61559 1 7963
2 61560 1 7963
2 61561 1 7963
2 61562 1 7963
2 61563 1 7971
2 61564 1 7971
2 61565 1 7971
2 61566 1 7971
2 61567 1 7971
2 61568 1 7971
2 61569 1 7972
2 61570 1 7972
2 61571 1 7973
2 61572 1 7973
2 61573 1 7981
2 61574 1 7981
2 61575 1 7996
2 61576 1 7996
2 61577 1 7997
2 61578 1 7997
2 61579 1 7997
2 61580 1 7997
2 61581 1 7997
2 61582 1 7997
2 61583 1 7997
2 61584 1 7997
2 61585 1 7997
2 61586 1 8005
2 61587 1 8005
2 61588 1 8005
2 61589 1 8006
2 61590 1 8006
2 61591 1 8007
2 61592 1 8007
2 61593 1 8007
2 61594 1 8007
2 61595 1 8007
2 61596 1 8007
2 61597 1 8007
2 61598 1 8007
2 61599 1 8007
2 61600 1 8018
2 61601 1 8018
2 61602 1 8023
2 61603 1 8023
2 61604 1 8023
2 61605 1 8023
2 61606 1 8024
2 61607 1 8024
2 61608 1 8024
2 61609 1 8036
2 61610 1 8036
2 61611 1 8036
2 61612 1 8036
2 61613 1 8036
2 61614 1 8044
2 61615 1 8044
2 61616 1 8045
2 61617 1 8045
2 61618 1 8046
2 61619 1 8046
2 61620 1 8055
2 61621 1 8055
2 61622 1 8063
2 61623 1 8063
2 61624 1 8063
2 61625 1 8063
2 61626 1 8071
2 61627 1 8071
2 61628 1 8071
2 61629 1 8072
2 61630 1 8072
2 61631 1 8072
2 61632 1 8072
2 61633 1 8072
2 61634 1 8072
2 61635 1 8072
2 61636 1 8072
2 61637 1 8072
2 61638 1 8072
2 61639 1 8075
2 61640 1 8075
2 61641 1 8075
2 61642 1 8075
2 61643 1 8075
2 61644 1 8075
2 61645 1 8075
2 61646 1 8075
2 61647 1 8075
2 61648 1 8075
2 61649 1 8075
2 61650 1 8075
2 61651 1 8075
2 61652 1 8075
2 61653 1 8075
2 61654 1 8075
2 61655 1 8075
2 61656 1 8075
2 61657 1 8075
2 61658 1 8075
2 61659 1 8075
2 61660 1 8075
2 61661 1 8077
2 61662 1 8077
2 61663 1 8077
2 61664 1 8077
2 61665 1 8077
2 61666 1 8077
2 61667 1 8085
2 61668 1 8085
2 61669 1 8086
2 61670 1 8086
2 61671 1 8087
2 61672 1 8087
2 61673 1 8087
2 61674 1 8087
2 61675 1 8087
2 61676 1 8096
2 61677 1 8096
2 61678 1 8113
2 61679 1 8113
2 61680 1 8113
2 61681 1 8114
2 61682 1 8114
2 61683 1 8116
2 61684 1 8116
2 61685 1 8121
2 61686 1 8121
2 61687 1 8121
2 61688 1 8121
2 61689 1 8122
2 61690 1 8122
2 61691 1 8122
2 61692 1 8123
2 61693 1 8123
2 61694 1 8123
2 61695 1 8123
2 61696 1 8123
2 61697 1 8123
2 61698 1 8128
2 61699 1 8128
2 61700 1 8131
2 61701 1 8131
2 61702 1 8131
2 61703 1 8132
2 61704 1 8132
2 61705 1 8132
2 61706 1 8132
2 61707 1 8132
2 61708 1 8133
2 61709 1 8133
2 61710 1 8134
2 61711 1 8134
2 61712 1 8143
2 61713 1 8143
2 61714 1 8144
2 61715 1 8144
2 61716 1 8144
2 61717 1 8144
2 61718 1 8145
2 61719 1 8145
2 61720 1 8145
2 61721 1 8159
2 61722 1 8159
2 61723 1 8159
2 61724 1 8162
2 61725 1 8162
2 61726 1 8162
2 61727 1 8162
2 61728 1 8162
2 61729 1 8162
2 61730 1 8162
2 61731 1 8169
2 61732 1 8169
2 61733 1 8170
2 61734 1 8170
2 61735 1 8170
2 61736 1 8170
2 61737 1 8194
2 61738 1 8194
2 61739 1 8194
2 61740 1 8194
2 61741 1 8194
2 61742 1 8194
2 61743 1 8194
2 61744 1 8194
2 61745 1 8195
2 61746 1 8195
2 61747 1 8195
2 61748 1 8195
2 61749 1 8195
2 61750 1 8195
2 61751 1 8195
2 61752 1 8196
2 61753 1 8196
2 61754 1 8198
2 61755 1 8198
2 61756 1 8198
2 61757 1 8206
2 61758 1 8206
2 61759 1 8214
2 61760 1 8214
2 61761 1 8221
2 61762 1 8221
2 61763 1 8221
2 61764 1 8222
2 61765 1 8222
2 61766 1 8222
2 61767 1 8222
2 61768 1 8222
2 61769 1 8222
2 61770 1 8222
2 61771 1 8223
2 61772 1 8223
2 61773 1 8224
2 61774 1 8224
2 61775 1 8224
2 61776 1 8228
2 61777 1 8228
2 61778 1 8228
2 61779 1 8236
2 61780 1 8236
2 61781 1 8237
2 61782 1 8237
2 61783 1 8237
2 61784 1 8237
2 61785 1 8237
2 61786 1 8237
2 61787 1 8244
2 61788 1 8244
2 61789 1 8244
2 61790 1 8245
2 61791 1 8245
2 61792 1 8245
2 61793 1 8245
2 61794 1 8257
2 61795 1 8257
2 61796 1 8257
2 61797 1 8261
2 61798 1 8261
2 61799 1 8261
2 61800 1 8262
2 61801 1 8262
2 61802 1 8262
2 61803 1 8262
2 61804 1 8263
2 61805 1 8263
2 61806 1 8263
2 61807 1 8263
2 61808 1 8271
2 61809 1 8271
2 61810 1 8272
2 61811 1 8272
2 61812 1 8273
2 61813 1 8273
2 61814 1 8281
2 61815 1 8281
2 61816 1 8281
2 61817 1 8281
2 61818 1 8286
2 61819 1 8286
2 61820 1 8286
2 61821 1 8286
2 61822 1 8286
2 61823 1 8286
2 61824 1 8286
2 61825 1 8286
2 61826 1 8286
2 61827 1 8286
2 61828 1 8287
2 61829 1 8287
2 61830 1 8301
2 61831 1 8301
2 61832 1 8301
2 61833 1 8301
2 61834 1 8303
2 61835 1 8303
2 61836 1 8303
2 61837 1 8303
2 61838 1 8303
2 61839 1 8303
2 61840 1 8303
2 61841 1 8304
2 61842 1 8304
2 61843 1 8306
2 61844 1 8306
2 61845 1 8307
2 61846 1 8307
2 61847 1 8308
2 61848 1 8308
2 61849 1 8321
2 61850 1 8321
2 61851 1 8321
2 61852 1 8321
2 61853 1 8321
2 61854 1 8321
2 61855 1 8321
2 61856 1 8321
2 61857 1 8321
2 61858 1 8321
2 61859 1 8322
2 61860 1 8322
2 61861 1 8322
2 61862 1 8322
2 61863 1 8323
2 61864 1 8323
2 61865 1 8328
2 61866 1 8328
2 61867 1 8328
2 61868 1 8328
2 61869 1 8336
2 61870 1 8336
2 61871 1 8336
2 61872 1 8336
2 61873 1 8339
2 61874 1 8339
2 61875 1 8339
2 61876 1 8339
2 61877 1 8339
2 61878 1 8339
2 61879 1 8339
2 61880 1 8340
2 61881 1 8340
2 61882 1 8340
2 61883 1 8340
2 61884 1 8340
2 61885 1 8340
2 61886 1 8340
2 61887 1 8355
2 61888 1 8355
2 61889 1 8355
2 61890 1 8355
2 61891 1 8359
2 61892 1 8359
2 61893 1 8360
2 61894 1 8360
2 61895 1 8360
2 61896 1 8368
2 61897 1 8368
2 61898 1 8368
2 61899 1 8373
2 61900 1 8373
2 61901 1 8376
2 61902 1 8376
2 61903 1 8377
2 61904 1 8377
2 61905 1 8386
2 61906 1 8386
2 61907 1 8397
2 61908 1 8397
2 61909 1 8407
2 61910 1 8407
2 61911 1 8407
2 61912 1 8413
2 61913 1 8413
2 61914 1 8428
2 61915 1 8428
2 61916 1 8428
2 61917 1 8428
2 61918 1 8428
2 61919 1 8430
2 61920 1 8430
2 61921 1 8448
2 61922 1 8448
2 61923 1 8448
2 61924 1 8448
2 61925 1 8452
2 61926 1 8452
2 61927 1 8452
2 61928 1 8452
2 61929 1 8452
2 61930 1 8453
2 61931 1 8453
2 61932 1 8453
2 61933 1 8453
2 61934 1 8472
2 61935 1 8472
2 61936 1 8473
2 61937 1 8473
2 61938 1 8474
2 61939 1 8474
2 61940 1 8474
2 61941 1 8497
2 61942 1 8497
2 61943 1 8498
2 61944 1 8498
2 61945 1 8500
2 61946 1 8500
2 61947 1 8502
2 61948 1 8502
2 61949 1 8505
2 61950 1 8505
2 61951 1 8505
2 61952 1 8505
2 61953 1 8505
2 61954 1 8506
2 61955 1 8506
2 61956 1 8508
2 61957 1 8508
2 61958 1 8520
2 61959 1 8520
2 61960 1 8520
2 61961 1 8521
2 61962 1 8521
2 61963 1 8524
2 61964 1 8524
2 61965 1 8524
2 61966 1 8526
2 61967 1 8526
2 61968 1 8526
2 61969 1 8529
2 61970 1 8529
2 61971 1 8536
2 61972 1 8536
2 61973 1 8537
2 61974 1 8537
2 61975 1 8537
2 61976 1 8537
2 61977 1 8546
2 61978 1 8546
2 61979 1 8547
2 61980 1 8547
2 61981 1 8555
2 61982 1 8555
2 61983 1 8556
2 61984 1 8556
2 61985 1 8557
2 61986 1 8557
2 61987 1 8567
2 61988 1 8567
2 61989 1 8567
2 61990 1 8567
2 61991 1 8567
2 61992 1 8567
2 61993 1 8568
2 61994 1 8568
2 61995 1 8571
2 61996 1 8571
2 61997 1 8572
2 61998 1 8572
2 61999 1 8572
2 62000 1 8575
2 62001 1 8575
2 62002 1 8575
2 62003 1 8576
2 62004 1 8576
2 62005 1 8579
2 62006 1 8579
2 62007 1 8589
2 62008 1 8589
2 62009 1 8589
2 62010 1 8589
2 62011 1 8589
2 62012 1 8589
2 62013 1 8589
2 62014 1 8592
2 62015 1 8592
2 62016 1 8592
2 62017 1 8593
2 62018 1 8593
2 62019 1 8604
2 62020 1 8604
2 62021 1 8613
2 62022 1 8613
2 62023 1 8613
2 62024 1 8613
2 62025 1 8627
2 62026 1 8627
2 62027 1 8630
2 62028 1 8630
2 62029 1 8632
2 62030 1 8632
2 62031 1 8637
2 62032 1 8637
2 62033 1 8654
2 62034 1 8654
2 62035 1 8657
2 62036 1 8657
2 62037 1 8657
2 62038 1 8657
2 62039 1 8657
2 62040 1 8660
2 62041 1 8660
2 62042 1 8671
2 62043 1 8671
2 62044 1 8671
2 62045 1 8682
2 62046 1 8682
2 62047 1 8682
2 62048 1 8709
2 62049 1 8709
2 62050 1 8723
2 62051 1 8723
2 62052 1 8728
2 62053 1 8728
2 62054 1 8732
2 62055 1 8732
2 62056 1 8732
2 62057 1 8736
2 62058 1 8736
2 62059 1 8737
2 62060 1 8737
2 62061 1 8738
2 62062 1 8738
2 62063 1 8739
2 62064 1 8739
2 62065 1 8747
2 62066 1 8747
2 62067 1 8747
2 62068 1 8747
2 62069 1 8747
2 62070 1 8748
2 62071 1 8748
2 62072 1 8748
2 62073 1 8748
2 62074 1 8749
2 62075 1 8749
2 62076 1 8750
2 62077 1 8750
2 62078 1 8750
2 62079 1 8758
2 62080 1 8758
2 62081 1 8758
2 62082 1 8762
2 62083 1 8762
2 62084 1 8762
2 62085 1 8762
2 62086 1 8762
2 62087 1 8762
2 62088 1 8762
2 62089 1 8762
2 62090 1 8762
2 62091 1 8762
2 62092 1 8762
2 62093 1 8776
2 62094 1 8776
2 62095 1 8776
2 62096 1 8776
2 62097 1 8776
2 62098 1 8777
2 62099 1 8777
2 62100 1 8780
2 62101 1 8780
2 62102 1 8784
2 62103 1 8784
2 62104 1 8784
2 62105 1 8784
2 62106 1 8786
2 62107 1 8786
2 62108 1 8800
2 62109 1 8800
2 62110 1 8800
2 62111 1 8800
2 62112 1 8801
2 62113 1 8801
2 62114 1 8808
2 62115 1 8808
2 62116 1 8808
2 62117 1 8809
2 62118 1 8809
2 62119 1 8816
2 62120 1 8816
2 62121 1 8818
2 62122 1 8818
2 62123 1 8842
2 62124 1 8842
2 62125 1 8842
2 62126 1 8842
2 62127 1 8842
2 62128 1 8842
2 62129 1 8842
2 62130 1 8842
2 62131 1 8842
2 62132 1 8842
2 62133 1 8842
2 62134 1 8842
2 62135 1 8842
2 62136 1 8842
2 62137 1 8842
2 62138 1 8842
2 62139 1 8843
2 62140 1 8843
2 62141 1 8843
2 62142 1 8847
2 62143 1 8847
2 62144 1 8854
2 62145 1 8854
2 62146 1 8864
2 62147 1 8864
2 62148 1 8875
2 62149 1 8875
2 62150 1 8875
2 62151 1 8897
2 62152 1 8897
2 62153 1 8908
2 62154 1 8908
2 62155 1 8908
2 62156 1 8908
2 62157 1 8922
2 62158 1 8922
2 62159 1 8931
2 62160 1 8931
2 62161 1 8931
2 62162 1 8931
2 62163 1 8931
2 62164 1 8931
2 62165 1 8931
2 62166 1 8944
2 62167 1 8944
2 62168 1 8944
2 62169 1 8949
2 62170 1 8949
2 62171 1 8949
2 62172 1 8962
2 62173 1 8962
2 62174 1 8962
2 62175 1 8964
2 62176 1 8964
2 62177 1 8965
2 62178 1 8965
2 62179 1 8965
2 62180 1 8965
2 62181 1 8992
2 62182 1 8992
2 62183 1 8992
2 62184 1 8992
2 62185 1 8992
2 62186 1 8993
2 62187 1 8993
2 62188 1 9017
2 62189 1 9017
2 62190 1 9017
2 62191 1 9017
2 62192 1 9018
2 62193 1 9018
2 62194 1 9034
2 62195 1 9034
2 62196 1 9034
2 62197 1 9034
2 62198 1 9034
2 62199 1 9034
2 62200 1 9034
2 62201 1 9034
2 62202 1 9034
2 62203 1 9034
2 62204 1 9034
2 62205 1 9035
2 62206 1 9035
2 62207 1 9035
2 62208 1 9035
2 62209 1 9037
2 62210 1 9037
2 62211 1 9053
2 62212 1 9053
2 62213 1 9054
2 62214 1 9054
2 62215 1 9054
2 62216 1 9054
2 62217 1 9057
2 62218 1 9057
2 62219 1 9062
2 62220 1 9062
2 62221 1 9062
2 62222 1 9063
2 62223 1 9063
2 62224 1 9071
2 62225 1 9071
2 62226 1 9072
2 62227 1 9072
2 62228 1 9072
2 62229 1 9075
2 62230 1 9075
2 62231 1 9080
2 62232 1 9080
2 62233 1 9080
2 62234 1 9080
2 62235 1 9080
2 62236 1 9080
2 62237 1 9107
2 62238 1 9107
2 62239 1 9111
2 62240 1 9111
2 62241 1 9111
2 62242 1 9111
2 62243 1 9111
2 62244 1 9113
2 62245 1 9113
2 62246 1 9113
2 62247 1 9129
2 62248 1 9129
2 62249 1 9136
2 62250 1 9136
2 62251 1 9138
2 62252 1 9138
2 62253 1 9139
2 62254 1 9139
2 62255 1 9140
2 62256 1 9140
2 62257 1 9141
2 62258 1 9141
2 62259 1 9141
2 62260 1 9159
2 62261 1 9159
2 62262 1 9159
2 62263 1 9160
2 62264 1 9160
2 62265 1 9172
2 62266 1 9172
2 62267 1 9175
2 62268 1 9175
2 62269 1 9175
2 62270 1 9176
2 62271 1 9176
2 62272 1 9176
2 62273 1 9176
2 62274 1 9176
2 62275 1 9176
2 62276 1 9176
2 62277 1 9176
2 62278 1 9176
2 62279 1 9177
2 62280 1 9177
2 62281 1 9177
2 62282 1 9177
2 62283 1 9177
2 62284 1 9181
2 62285 1 9181
2 62286 1 9182
2 62287 1 9182
2 62288 1 9183
2 62289 1 9183
2 62290 1 9183
2 62291 1 9183
2 62292 1 9183
2 62293 1 9183
2 62294 1 9206
2 62295 1 9206
2 62296 1 9215
2 62297 1 9215
2 62298 1 9222
2 62299 1 9222
2 62300 1 9222
2 62301 1 9222
2 62302 1 9223
2 62303 1 9223
2 62304 1 9223
2 62305 1 9224
2 62306 1 9224
2 62307 1 9225
2 62308 1 9225
2 62309 1 9225
2 62310 1 9225
2 62311 1 9227
2 62312 1 9227
2 62313 1 9234
2 62314 1 9234
2 62315 1 9245
2 62316 1 9245
2 62317 1 9246
2 62318 1 9246
2 62319 1 9250
2 62320 1 9250
2 62321 1 9250
2 62322 1 9250
2 62323 1 9255
2 62324 1 9255
2 62325 1 9261
2 62326 1 9261
2 62327 1 9262
2 62328 1 9262
2 62329 1 9262
2 62330 1 9262
2 62331 1 9264
2 62332 1 9264
2 62333 1 9264
2 62334 1 9264
2 62335 1 9264
2 62336 1 9265
2 62337 1 9265
2 62338 1 9265
2 62339 1 9265
2 62340 1 9265
2 62341 1 9266
2 62342 1 9266
2 62343 1 9267
2 62344 1 9267
2 62345 1 9271
2 62346 1 9271
2 62347 1 9271
2 62348 1 9271
2 62349 1 9272
2 62350 1 9272
2 62351 1 9276
2 62352 1 9276
2 62353 1 9276
2 62354 1 9288
2 62355 1 9288
2 62356 1 9288
2 62357 1 9289
2 62358 1 9289
2 62359 1 9289
2 62360 1 9289
2 62361 1 9297
2 62362 1 9297
2 62363 1 9297
2 62364 1 9297
2 62365 1 9297
2 62366 1 9297
2 62367 1 9297
2 62368 1 9297
2 62369 1 9298
2 62370 1 9298
2 62371 1 9299
2 62372 1 9299
2 62373 1 9301
2 62374 1 9301
2 62375 1 9317
2 62376 1 9317
2 62377 1 9317
2 62378 1 9319
2 62379 1 9319
2 62380 1 9333
2 62381 1 9333
2 62382 1 9336
2 62383 1 9336
2 62384 1 9338
2 62385 1 9338
2 62386 1 9340
2 62387 1 9340
2 62388 1 9340
2 62389 1 9343
2 62390 1 9343
2 62391 1 9344
2 62392 1 9344
2 62393 1 9346
2 62394 1 9346
2 62395 1 9349
2 62396 1 9349
2 62397 1 9349
2 62398 1 9349
2 62399 1 9349
2 62400 1 9349
2 62401 1 9351
2 62402 1 9351
2 62403 1 9351
2 62404 1 9351
2 62405 1 9351
2 62406 1 9356
2 62407 1 9356
2 62408 1 9359
2 62409 1 9359
2 62410 1 9364
2 62411 1 9364
2 62412 1 9364
2 62413 1 9364
2 62414 1 9364
2 62415 1 9365
2 62416 1 9365
2 62417 1 9365
2 62418 1 9366
2 62419 1 9366
2 62420 1 9366
2 62421 1 9367
2 62422 1 9367
2 62423 1 9372
2 62424 1 9372
2 62425 1 9374
2 62426 1 9374
2 62427 1 9374
2 62428 1 9399
2 62429 1 9399
2 62430 1 9401
2 62431 1 9401
2 62432 1 9407
2 62433 1 9407
2 62434 1 9407
2 62435 1 9409
2 62436 1 9409
2 62437 1 9410
2 62438 1 9410
2 62439 1 9419
2 62440 1 9419
2 62441 1 9419
2 62442 1 9420
2 62443 1 9420
2 62444 1 9420
2 62445 1 9421
2 62446 1 9421
2 62447 1 9430
2 62448 1 9430
2 62449 1 9439
2 62450 1 9439
2 62451 1 9450
2 62452 1 9450
2 62453 1 9450
2 62454 1 9466
2 62455 1 9466
2 62456 1 9470
2 62457 1 9470
2 62458 1 9471
2 62459 1 9471
2 62460 1 9471
2 62461 1 9471
2 62462 1 9479
2 62463 1 9479
2 62464 1 9480
2 62465 1 9480
2 62466 1 9480
2 62467 1 9494
2 62468 1 9494
2 62469 1 9494
2 62470 1 9494
2 62471 1 9494
2 62472 1 9494
2 62473 1 9502
2 62474 1 9502
2 62475 1 9518
2 62476 1 9518
2 62477 1 9518
2 62478 1 9518
2 62479 1 9518
2 62480 1 9518
2 62481 1 9527
2 62482 1 9527
2 62483 1 9527
2 62484 1 9527
2 62485 1 9527
2 62486 1 9527
2 62487 1 9527
2 62488 1 9527
2 62489 1 9527
2 62490 1 9527
2 62491 1 9527
2 62492 1 9527
2 62493 1 9527
2 62494 1 9527
2 62495 1 9527
2 62496 1 9527
2 62497 1 9527
2 62498 1 9527
2 62499 1 9527
2 62500 1 9527
2 62501 1 9527
2 62502 1 9527
2 62503 1 9527
2 62504 1 9527
2 62505 1 9527
2 62506 1 9527
2 62507 1 9527
2 62508 1 9527
2 62509 1 9527
2 62510 1 9527
2 62511 1 9527
2 62512 1 9527
2 62513 1 9527
2 62514 1 9527
2 62515 1 9527
2 62516 1 9527
2 62517 1 9527
2 62518 1 9527
2 62519 1 9527
2 62520 1 9527
2 62521 1 9527
2 62522 1 9527
2 62523 1 9527
2 62524 1 9527
2 62525 1 9527
2 62526 1 9527
2 62527 1 9527
2 62528 1 9527
2 62529 1 9527
2 62530 1 9527
2 62531 1 9527
2 62532 1 9527
2 62533 1 9527
2 62534 1 9527
2 62535 1 9527
2 62536 1 9527
2 62537 1 9527
2 62538 1 9527
2 62539 1 9527
2 62540 1 9527
2 62541 1 9527
2 62542 1 9527
2 62543 1 9527
2 62544 1 9527
2 62545 1 9527
2 62546 1 9527
2 62547 1 9527
2 62548 1 9527
2 62549 1 9527
2 62550 1 9528
2 62551 1 9528
2 62552 1 9528
2 62553 1 9531
2 62554 1 9531
2 62555 1 9544
2 62556 1 9544
2 62557 1 9552
2 62558 1 9552
2 62559 1 9560
2 62560 1 9560
2 62561 1 9561
2 62562 1 9561
2 62563 1 9561
2 62564 1 9561
2 62565 1 9604
2 62566 1 9604
2 62567 1 9604
2 62568 1 9604
2 62569 1 9604
2 62570 1 9604
2 62571 1 9612
2 62572 1 9612
2 62573 1 9620
2 62574 1 9620
2 62575 1 9623
2 62576 1 9623
2 62577 1 9623
2 62578 1 9627
2 62579 1 9627
2 62580 1 9627
2 62581 1 9639
2 62582 1 9639
2 62583 1 9639
2 62584 1 9645
2 62585 1 9645
2 62586 1 9645
2 62587 1 9645
2 62588 1 9645
2 62589 1 9645
2 62590 1 9645
2 62591 1 9645
2 62592 1 9645
2 62593 1 9645
2 62594 1 9646
2 62595 1 9646
2 62596 1 9655
2 62597 1 9655
2 62598 1 9656
2 62599 1 9656
2 62600 1 9656
2 62601 1 9656
2 62602 1 9661
2 62603 1 9661
2 62604 1 9666
2 62605 1 9666
2 62606 1 9672
2 62607 1 9672
2 62608 1 9672
2 62609 1 9673
2 62610 1 9673
2 62611 1 9676
2 62612 1 9676
2 62613 1 9677
2 62614 1 9677
2 62615 1 9692
2 62616 1 9692
2 62617 1 9693
2 62618 1 9693
2 62619 1 9696
2 62620 1 9696
2 62621 1 9696
2 62622 1 9696
2 62623 1 9696
2 62624 1 9697
2 62625 1 9697
2 62626 1 9714
2 62627 1 9714
2 62628 1 9724
2 62629 1 9724
2 62630 1 9724
2 62631 1 9724
2 62632 1 9724
2 62633 1 9731
2 62634 1 9731
2 62635 1 9761
2 62636 1 9761
2 62637 1 9761
2 62638 1 9761
2 62639 1 9762
2 62640 1 9762
2 62641 1 9778
2 62642 1 9778
2 62643 1 9779
2 62644 1 9779
2 62645 1 9779
2 62646 1 9779
2 62647 1 9779
2 62648 1 9789
2 62649 1 9789
2 62650 1 9789
2 62651 1 9789
2 62652 1 9789
2 62653 1 9793
2 62654 1 9793
2 62655 1 9793
2 62656 1 9793
2 62657 1 9793
2 62658 1 9793
2 62659 1 9793
2 62660 1 9793
2 62661 1 9796
2 62662 1 9796
2 62663 1 9797
2 62664 1 9797
2 62665 1 9814
2 62666 1 9814
2 62667 1 9814
2 62668 1 9814
2 62669 1 9814
2 62670 1 9814
2 62671 1 9815
2 62672 1 9815
2 62673 1 9817
2 62674 1 9817
2 62675 1 9817
2 62676 1 9817
2 62677 1 9817
2 62678 1 9817
2 62679 1 9817
2 62680 1 9817
2 62681 1 9821
2 62682 1 9821
2 62683 1 9821
2 62684 1 9821
2 62685 1 9821
2 62686 1 9821
2 62687 1 9821
2 62688 1 9821
2 62689 1 9821
2 62690 1 9821
2 62691 1 9821
2 62692 1 9821
2 62693 1 9821
2 62694 1 9821
2 62695 1 9824
2 62696 1 9824
2 62697 1 9824
2 62698 1 9824
2 62699 1 9824
2 62700 1 9825
2 62701 1 9825
2 62702 1 9825
2 62703 1 9825
2 62704 1 9825
2 62705 1 9825
2 62706 1 9825
2 62707 1 9825
2 62708 1 9825
2 62709 1 9825
2 62710 1 9825
2 62711 1 9825
2 62712 1 9825
2 62713 1 9825
2 62714 1 9825
2 62715 1 9825
2 62716 1 9825
2 62717 1 9827
2 62718 1 9827
2 62719 1 9827
2 62720 1 9827
2 62721 1 9827
2 62722 1 9827
2 62723 1 9828
2 62724 1 9828
2 62725 1 9828
2 62726 1 9828
2 62727 1 9828
2 62728 1 9828
2 62729 1 9828
2 62730 1 9828
2 62731 1 9828
2 62732 1 9828
2 62733 1 9828
2 62734 1 9828
2 62735 1 9828
2 62736 1 9828
2 62737 1 9828
2 62738 1 9828
2 62739 1 9828
2 62740 1 9828
2 62741 1 9828
2 62742 1 9829
2 62743 1 9829
2 62744 1 9829
2 62745 1 9829
2 62746 1 9829
2 62747 1 9829
2 62748 1 9829
2 62749 1 9830
2 62750 1 9830
2 62751 1 9830
2 62752 1 9830
2 62753 1 9830
2 62754 1 9830
2 62755 1 9830
2 62756 1 9830
2 62757 1 9830
2 62758 1 9831
2 62759 1 9831
2 62760 1 9832
2 62761 1 9832
2 62762 1 9834
2 62763 1 9834
2 62764 1 9834
2 62765 1 9834
2 62766 1 9834
2 62767 1 9841
2 62768 1 9841
2 62769 1 9842
2 62770 1 9842
2 62771 1 9842
2 62772 1 9843
2 62773 1 9843
2 62774 1 9849
2 62775 1 9849
2 62776 1 9849
2 62777 1 9851
2 62778 1 9851
2 62779 1 9851
2 62780 1 9851
2 62781 1 9852
2 62782 1 9852
2 62783 1 9853
2 62784 1 9853
2 62785 1 9855
2 62786 1 9855
2 62787 1 9856
2 62788 1 9856
2 62789 1 9857
2 62790 1 9857
2 62791 1 9859
2 62792 1 9859
2 62793 1 9859
2 62794 1 9859
2 62795 1 9887
2 62796 1 9887
2 62797 1 9887
2 62798 1 9887
2 62799 1 9887
2 62800 1 9887
2 62801 1 9887
2 62802 1 9888
2 62803 1 9888
2 62804 1 9889
2 62805 1 9889
2 62806 1 9893
2 62807 1 9893
2 62808 1 9893
2 62809 1 9911
2 62810 1 9911
2 62811 1 9911
2 62812 1 9911
2 62813 1 9911
2 62814 1 9914
2 62815 1 9914
2 62816 1 9914
2 62817 1 9914
2 62818 1 9914
2 62819 1 9914
2 62820 1 9914
2 62821 1 9915
2 62822 1 9915
2 62823 1 9925
2 62824 1 9925
2 62825 1 9925
2 62826 1 9925
2 62827 1 9944
2 62828 1 9944
2 62829 1 9963
2 62830 1 9963
2 62831 1 9975
2 62832 1 9975
2 62833 1 9975
2 62834 1 9975
2 62835 1 9975
2 62836 1 9975
2 62837 1 9975
2 62838 1 9975
2 62839 1 9977
2 62840 1 9977
2 62841 1 9977
2 62842 1 9982
2 62843 1 9982
2 62844 1 9982
2 62845 1 9982
2 62846 1 9982
2 62847 1 9982
2 62848 1 9982
2 62849 1 9983
2 62850 1 9983
2 62851 1 9983
2 62852 1 9983
2 62853 1 9983
2 62854 1 9983
2 62855 1 9983
2 62856 1 9983
2 62857 1 10002
2 62858 1 10002
2 62859 1 10002
2 62860 1 10002
2 62861 1 10004
2 62862 1 10004
2 62863 1 10007
2 62864 1 10007
2 62865 1 10007
2 62866 1 10007
2 62867 1 10007
2 62868 1 10008
2 62869 1 10008
2 62870 1 10008
2 62871 1 10008
2 62872 1 10008
2 62873 1 10008
2 62874 1 10022
2 62875 1 10022
2 62876 1 10034
2 62877 1 10034
2 62878 1 10042
2 62879 1 10042
2 62880 1 10042
2 62881 1 10042
2 62882 1 10042
2 62883 1 10042
2 62884 1 10042
2 62885 1 10042
2 62886 1 10042
2 62887 1 10042
2 62888 1 10042
2 62889 1 10044
2 62890 1 10044
2 62891 1 10047
2 62892 1 10047
2 62893 1 10048
2 62894 1 10048
2 62895 1 10070
2 62896 1 10070
2 62897 1 10070
2 62898 1 10076
2 62899 1 10076
2 62900 1 10076
2 62901 1 10126
2 62902 1 10126
2 62903 1 10126
2 62904 1 10126
2 62905 1 10127
2 62906 1 10127
2 62907 1 10127
2 62908 1 10127
2 62909 1 10129
2 62910 1 10129
2 62911 1 10129
2 62912 1 10129
2 62913 1 10129
2 62914 1 10129
2 62915 1 10129
2 62916 1 10129
2 62917 1 10129
2 62918 1 10129
2 62919 1 10129
2 62920 1 10129
2 62921 1 10129
2 62922 1 10129
2 62923 1 10129
2 62924 1 10129
2 62925 1 10129
2 62926 1 10129
2 62927 1 10129
2 62928 1 10129
2 62929 1 10131
2 62930 1 10131
2 62931 1 10132
2 62932 1 10132
2 62933 1 10132
2 62934 1 10132
2 62935 1 10132
2 62936 1 10133
2 62937 1 10133
2 62938 1 10148
2 62939 1 10148
2 62940 1 10148
2 62941 1 10148
2 62942 1 10151
2 62943 1 10151
2 62944 1 10151
2 62945 1 10151
2 62946 1 10152
2 62947 1 10152
2 62948 1 10153
2 62949 1 10153
2 62950 1 10154
2 62951 1 10154
2 62952 1 10162
2 62953 1 10162
2 62954 1 10164
2 62955 1 10164
2 62956 1 10164
2 62957 1 10165
2 62958 1 10165
2 62959 1 10165
2 62960 1 10165
2 62961 1 10168
2 62962 1 10168
2 62963 1 10168
2 62964 1 10169
2 62965 1 10169
2 62966 1 10170
2 62967 1 10170
2 62968 1 10181
2 62969 1 10181
2 62970 1 10181
2 62971 1 10181
2 62972 1 10184
2 62973 1 10184
2 62974 1 10184
2 62975 1 10184
2 62976 1 10184
2 62977 1 10185
2 62978 1 10185
2 62979 1 10185
2 62980 1 10194
2 62981 1 10194
2 62982 1 10201
2 62983 1 10201
2 62984 1 10203
2 62985 1 10203
2 62986 1 10203
2 62987 1 10203
2 62988 1 10203
2 62989 1 10203
2 62990 1 10203
2 62991 1 10203
2 62992 1 10207
2 62993 1 10207
2 62994 1 10207
2 62995 1 10207
2 62996 1 10207
2 62997 1 10207
2 62998 1 10207
2 62999 1 10207
2 63000 1 10207
2 63001 1 10207
2 63002 1 10207
2 63003 1 10207
2 63004 1 10217
2 63005 1 10217
2 63006 1 10217
2 63007 1 10217
2 63008 1 10217
2 63009 1 10217
2 63010 1 10225
2 63011 1 10225
2 63012 1 10232
2 63013 1 10232
2 63014 1 10234
2 63015 1 10234
2 63016 1 10234
2 63017 1 10234
2 63018 1 10234
2 63019 1 10234
2 63020 1 10234
2 63021 1 10234
2 63022 1 10234
2 63023 1 10234
2 63024 1 10234
2 63025 1 10234
2 63026 1 10234
2 63027 1 10234
2 63028 1 10234
2 63029 1 10234
2 63030 1 10234
2 63031 1 10234
2 63032 1 10235
2 63033 1 10235
2 63034 1 10235
2 63035 1 10235
2 63036 1 10235
2 63037 1 10238
2 63038 1 10238
2 63039 1 10238
2 63040 1 10238
2 63041 1 10239
2 63042 1 10239
2 63043 1 10239
2 63044 1 10239
2 63045 1 10239
2 63046 1 10239
2 63047 1 10239
2 63048 1 10239
2 63049 1 10239
2 63050 1 10239
2 63051 1 10239
2 63052 1 10239
2 63053 1 10239
2 63054 1 10240
2 63055 1 10240
2 63056 1 10240
2 63057 1 10265
2 63058 1 10265
2 63059 1 10282
2 63060 1 10282
2 63061 1 10282
2 63062 1 10282
2 63063 1 10282
2 63064 1 10282
2 63065 1 10282
2 63066 1 10282
2 63067 1 10282
2 63068 1 10282
2 63069 1 10282
2 63070 1 10282
2 63071 1 10282
2 63072 1 10282
2 63073 1 10282
2 63074 1 10282
2 63075 1 10282
2 63076 1 10282
2 63077 1 10282
2 63078 1 10283
2 63079 1 10283
2 63080 1 10284
2 63081 1 10284
2 63082 1 10284
2 63083 1 10284
2 63084 1 10284
2 63085 1 10284
2 63086 1 10298
2 63087 1 10298
2 63088 1 10298
2 63089 1 10298
2 63090 1 10298
2 63091 1 10298
2 63092 1 10298
2 63093 1 10298
2 63094 1 10298
2 63095 1 10298
2 63096 1 10298
2 63097 1 10299
2 63098 1 10299
2 63099 1 10299
2 63100 1 10306
2 63101 1 10306
2 63102 1 10306
2 63103 1 10306
2 63104 1 10306
2 63105 1 10307
2 63106 1 10307
2 63107 1 10308
2 63108 1 10308
2 63109 1 10309
2 63110 1 10309
2 63111 1 10309
2 63112 1 10309
2 63113 1 10309
2 63114 1 10309
2 63115 1 10309
2 63116 1 10309
2 63117 1 10309
2 63118 1 10309
2 63119 1 10309
2 63120 1 10309
2 63121 1 10309
2 63122 1 10309
2 63123 1 10309
2 63124 1 10309
2 63125 1 10309
2 63126 1 10309
2 63127 1 10310
2 63128 1 10310
2 63129 1 10323
2 63130 1 10323
2 63131 1 10323
2 63132 1 10323
2 63133 1 10323
2 63134 1 10323
2 63135 1 10323
2 63136 1 10323
2 63137 1 10324
2 63138 1 10324
2 63139 1 10325
2 63140 1 10325
2 63141 1 10325
2 63142 1 10347
2 63143 1 10347
2 63144 1 10348
2 63145 1 10348
2 63146 1 10348
2 63147 1 10348
2 63148 1 10349
2 63149 1 10349
2 63150 1 10382
2 63151 1 10382
2 63152 1 10382
2 63153 1 10382
2 63154 1 10382
2 63155 1 10382
2 63156 1 10382
2 63157 1 10382
2 63158 1 10382
2 63159 1 10384
2 63160 1 10384
2 63161 1 10401
2 63162 1 10401
2 63163 1 10417
2 63164 1 10417
2 63165 1 10417
2 63166 1 10425
2 63167 1 10425
2 63168 1 10425
2 63169 1 10429
2 63170 1 10429
2 63171 1 10429
2 63172 1 10433
2 63173 1 10433
2 63174 1 10433
2 63175 1 10433
2 63176 1 10433
2 63177 1 10433
2 63178 1 10434
2 63179 1 10434
2 63180 1 10434
2 63181 1 10434
2 63182 1 10505
2 63183 1 10505
2 63184 1 10505
2 63185 1 10518
2 63186 1 10518
2 63187 1 10518
2 63188 1 10518
2 63189 1 10518
2 63190 1 10518
2 63191 1 10518
2 63192 1 10518
2 63193 1 10518
2 63194 1 10518
2 63195 1 10518
2 63196 1 10518
2 63197 1 10518
2 63198 1 10519
2 63199 1 10519
2 63200 1 10536
2 63201 1 10536
2 63202 1 10536
2 63203 1 10538
2 63204 1 10538
2 63205 1 10539
2 63206 1 10539
2 63207 1 10543
2 63208 1 10543
2 63209 1 10544
2 63210 1 10544
2 63211 1 10544
2 63212 1 10544
2 63213 1 10544
2 63214 1 10544
2 63215 1 10544
2 63216 1 10544
2 63217 1 10544
2 63218 1 10552
2 63219 1 10552
2 63220 1 10552
2 63221 1 10552
2 63222 1 10552
2 63223 1 10552
2 63224 1 10552
2 63225 1 10554
2 63226 1 10554
2 63227 1 10554
2 63228 1 10554
2 63229 1 10554
2 63230 1 10554
2 63231 1 10554
2 63232 1 10554
2 63233 1 10555
2 63234 1 10555
2 63235 1 10556
2 63236 1 10556
2 63237 1 10556
2 63238 1 10556
2 63239 1 10556
2 63240 1 10559
2 63241 1 10559
2 63242 1 10575
2 63243 1 10575
2 63244 1 10575
2 63245 1 10575
2 63246 1 10576
2 63247 1 10576
2 63248 1 10576
2 63249 1 10576
2 63250 1 10576
2 63251 1 10576
2 63252 1 10576
2 63253 1 10577
2 63254 1 10577
2 63255 1 10578
2 63256 1 10578
2 63257 1 10582
2 63258 1 10582
2 63259 1 10582
2 63260 1 10582
2 63261 1 10582
2 63262 1 10582
2 63263 1 10588
2 63264 1 10588
2 63265 1 10597
2 63266 1 10597
2 63267 1 10597
2 63268 1 10602
2 63269 1 10602
2 63270 1 10603
2 63271 1 10603
2 63272 1 10604
2 63273 1 10604
2 63274 1 10618
2 63275 1 10618
2 63276 1 10618
2 63277 1 10619
2 63278 1 10619
2 63279 1 10619
2 63280 1 10619
2 63281 1 10619
2 63282 1 10619
2 63283 1 10619
2 63284 1 10622
2 63285 1 10622
2 63286 1 10622
2 63287 1 10622
2 63288 1 10631
2 63289 1 10631
2 63290 1 10631
2 63291 1 10631
2 63292 1 10631
2 63293 1 10631
2 63294 1 10631
2 63295 1 10631
2 63296 1 10631
2 63297 1 10631
2 63298 1 10631
2 63299 1 10631
2 63300 1 10631
2 63301 1 10632
2 63302 1 10632
2 63303 1 10632
2 63304 1 10632
2 63305 1 10634
2 63306 1 10634
2 63307 1 10635
2 63308 1 10635
2 63309 1 10635
2 63310 1 10635
2 63311 1 10635
2 63312 1 10635
2 63313 1 10635
2 63314 1 10635
2 63315 1 10635
2 63316 1 10639
2 63317 1 10639
2 63318 1 10641
2 63319 1 10641
2 63320 1 10641
2 63321 1 10641
2 63322 1 10641
2 63323 1 10642
2 63324 1 10642
2 63325 1 10643
2 63326 1 10643
2 63327 1 10648
2 63328 1 10648
2 63329 1 10651
2 63330 1 10651
2 63331 1 10651
2 63332 1 10651
2 63333 1 10655
2 63334 1 10655
2 63335 1 10655
2 63336 1 10655
2 63337 1 10655
2 63338 1 10669
2 63339 1 10669
2 63340 1 10669
2 63341 1 10669
2 63342 1 10669
2 63343 1 10669
2 63344 1 10669
2 63345 1 10669
2 63346 1 10669
2 63347 1 10671
2 63348 1 10671
2 63349 1 10671
2 63350 1 10671
2 63351 1 10672
2 63352 1 10672
2 63353 1 10682
2 63354 1 10682
2 63355 1 10682
2 63356 1 10683
2 63357 1 10683
2 63358 1 10683
2 63359 1 10684
2 63360 1 10684
2 63361 1 10698
2 63362 1 10698
2 63363 1 10700
2 63364 1 10700
2 63365 1 10700
2 63366 1 10703
2 63367 1 10703
2 63368 1 10714
2 63369 1 10714
2 63370 1 10714
2 63371 1 10714
2 63372 1 10715
2 63373 1 10715
2 63374 1 10715
2 63375 1 10715
2 63376 1 10715
2 63377 1 10715
2 63378 1 10715
2 63379 1 10715
2 63380 1 10715
2 63381 1 10718
2 63382 1 10718
2 63383 1 10718
2 63384 1 10718
2 63385 1 10719
2 63386 1 10719
2 63387 1 10719
2 63388 1 10719
2 63389 1 10719
2 63390 1 10719
2 63391 1 10719
2 63392 1 10719
2 63393 1 10719
2 63394 1 10720
2 63395 1 10720
2 63396 1 10720
2 63397 1 10720
2 63398 1 10729
2 63399 1 10729
2 63400 1 10729
2 63401 1 10729
2 63402 1 10729
2 63403 1 10729
2 63404 1 10729
2 63405 1 10729
2 63406 1 10730
2 63407 1 10730
2 63408 1 10730
2 63409 1 10730
2 63410 1 10730
2 63411 1 10730
2 63412 1 10730
2 63413 1 10731
2 63414 1 10731
2 63415 1 10732
2 63416 1 10732
2 63417 1 10732
2 63418 1 10732
2 63419 1 10732
2 63420 1 10732
2 63421 1 10732
2 63422 1 10732
2 63423 1 10732
2 63424 1 10732
2 63425 1 10732
2 63426 1 10733
2 63427 1 10733
2 63428 1 10733
2 63429 1 10733
2 63430 1 10747
2 63431 1 10747
2 63432 1 10757
2 63433 1 10757
2 63434 1 10757
2 63435 1 10767
2 63436 1 10767
2 63437 1 10768
2 63438 1 10768
2 63439 1 10771
2 63440 1 10771
2 63441 1 10771
2 63442 1 10771
2 63443 1 10771
2 63444 1 10771
2 63445 1 10772
2 63446 1 10772
2 63447 1 10774
2 63448 1 10774
2 63449 1 10789
2 63450 1 10789
2 63451 1 10789
2 63452 1 10797
2 63453 1 10797
2 63454 1 10797
2 63455 1 10797
2 63456 1 10797
2 63457 1 10797
2 63458 1 10797
2 63459 1 10798
2 63460 1 10798
2 63461 1 10799
2 63462 1 10799
2 63463 1 10799
2 63464 1 10799
2 63465 1 10799
2 63466 1 10807
2 63467 1 10807
2 63468 1 10807
2 63469 1 10807
2 63470 1 10810
2 63471 1 10810
2 63472 1 10811
2 63473 1 10811
2 63474 1 10832
2 63475 1 10832
2 63476 1 10832
2 63477 1 10832
2 63478 1 10832
2 63479 1 10833
2 63480 1 10833
2 63481 1 10839
2 63482 1 10839
2 63483 1 10840
2 63484 1 10840
2 63485 1 10840
2 63486 1 10856
2 63487 1 10856
2 63488 1 10864
2 63489 1 10864
2 63490 1 10877
2 63491 1 10877
2 63492 1 10877
2 63493 1 10877
2 63494 1 10877
2 63495 1 10877
2 63496 1 10877
2 63497 1 10878
2 63498 1 10878
2 63499 1 10878
2 63500 1 10878
2 63501 1 10879
2 63502 1 10879
2 63503 1 10880
2 63504 1 10880
2 63505 1 10882
2 63506 1 10882
2 63507 1 10882
2 63508 1 10884
2 63509 1 10884
2 63510 1 10887
2 63511 1 10887
2 63512 1 10888
2 63513 1 10888
2 63514 1 10888
2 63515 1 10888
2 63516 1 10888
2 63517 1 10889
2 63518 1 10889
2 63519 1 10892
2 63520 1 10892
2 63521 1 10902
2 63522 1 10902
2 63523 1 10904
2 63524 1 10904
2 63525 1 10905
2 63526 1 10905
2 63527 1 10905
2 63528 1 10905
2 63529 1 10906
2 63530 1 10906
2 63531 1 10906
2 63532 1 10926
2 63533 1 10926
2 63534 1 10926
2 63535 1 10929
2 63536 1 10929
2 63537 1 10930
2 63538 1 10930
2 63539 1 10935
2 63540 1 10935
2 63541 1 10935
2 63542 1 10935
2 63543 1 10935
2 63544 1 10935
2 63545 1 10935
2 63546 1 10935
2 63547 1 10935
2 63548 1 10935
2 63549 1 10935
2 63550 1 10943
2 63551 1 10943
2 63552 1 10943
2 63553 1 10943
2 63554 1 10943
2 63555 1 10943
2 63556 1 10943
2 63557 1 10945
2 63558 1 10945
2 63559 1 10946
2 63560 1 10946
2 63561 1 10949
2 63562 1 10949
2 63563 1 10954
2 63564 1 10954
2 63565 1 10965
2 63566 1 10965
2 63567 1 10965
2 63568 1 10965
2 63569 1 10965
2 63570 1 10965
2 63571 1 10966
2 63572 1 10966
2 63573 1 10966
2 63574 1 10966
2 63575 1 10966
2 63576 1 10966
2 63577 1 10966
2 63578 1 10970
2 63579 1 10970
2 63580 1 10970
2 63581 1 10980
2 63582 1 10980
2 63583 1 10990
2 63584 1 10990
2 63585 1 10994
2 63586 1 10994
2 63587 1 10997
2 63588 1 10997
2 63589 1 11000
2 63590 1 11000
2 63591 1 11000
2 63592 1 11000
2 63593 1 11000
2 63594 1 11000
2 63595 1 11007
2 63596 1 11007
2 63597 1 11008
2 63598 1 11008
2 63599 1 11008
2 63600 1 11008
2 63601 1 11010
2 63602 1 11010
2 63603 1 11010
2 63604 1 11010
2 63605 1 11010
2 63606 1 11010
2 63607 1 11010
2 63608 1 11010
2 63609 1 11010
2 63610 1 11010
2 63611 1 11010
2 63612 1 11010
2 63613 1 11010
2 63614 1 11010
2 63615 1 11010
2 63616 1 11010
2 63617 1 11010
2 63618 1 11010
2 63619 1 11010
2 63620 1 11022
2 63621 1 11022
2 63622 1 11023
2 63623 1 11023
2 63624 1 11024
2 63625 1 11024
2 63626 1 11024
2 63627 1 11024
2 63628 1 11027
2 63629 1 11027
2 63630 1 11041
2 63631 1 11041
2 63632 1 11041
2 63633 1 11042
2 63634 1 11042
2 63635 1 11042
2 63636 1 11042
2 63637 1 11049
2 63638 1 11049
2 63639 1 11049
2 63640 1 11051
2 63641 1 11051
2 63642 1 11066
2 63643 1 11066
2 63644 1 11067
2 63645 1 11067
2 63646 1 11076
2 63647 1 11076
2 63648 1 11077
2 63649 1 11077
2 63650 1 11077
2 63651 1 11077
2 63652 1 11077
2 63653 1 11077
2 63654 1 11077
2 63655 1 11077
2 63656 1 11078
2 63657 1 11078
2 63658 1 11079
2 63659 1 11079
2 63660 1 11094
2 63661 1 11094
2 63662 1 11094
2 63663 1 11094
2 63664 1 11094
2 63665 1 11094
2 63666 1 11094
2 63667 1 11095
2 63668 1 11095
2 63669 1 11096
2 63670 1 11096
2 63671 1 11102
2 63672 1 11102
2 63673 1 11102
2 63674 1 11102
2 63675 1 11102
2 63676 1 11114
2 63677 1 11114
2 63678 1 11114
2 63679 1 11115
2 63680 1 11115
2 63681 1 11115
2 63682 1 11117
2 63683 1 11117
2 63684 1 11117
2 63685 1 11117
2 63686 1 11117
2 63687 1 11117
2 63688 1 11117
2 63689 1 11117
2 63690 1 11117
2 63691 1 11118
2 63692 1 11118
2 63693 1 11118
2 63694 1 11118
2 63695 1 11118
2 63696 1 11118
2 63697 1 11118
2 63698 1 11128
2 63699 1 11128
2 63700 1 11128
2 63701 1 11128
2 63702 1 11128
2 63703 1 11128
2 63704 1 11128
2 63705 1 11128
2 63706 1 11128
2 63707 1 11128
2 63708 1 11128
2 63709 1 11131
2 63710 1 11131
2 63711 1 11131
2 63712 1 11131
2 63713 1 11135
2 63714 1 11135
2 63715 1 11135
2 63716 1 11135
2 63717 1 11138
2 63718 1 11138
2 63719 1 11138
2 63720 1 11160
2 63721 1 11160
2 63722 1 11160
2 63723 1 11160
2 63724 1 11160
2 63725 1 11187
2 63726 1 11187
2 63727 1 11187
2 63728 1 11187
2 63729 1 11187
2 63730 1 11187
2 63731 1 11187
2 63732 1 11187
2 63733 1 11187
2 63734 1 11187
2 63735 1 11187
2 63736 1 11187
2 63737 1 11187
2 63738 1 11187
2 63739 1 11187
2 63740 1 11187
2 63741 1 11187
2 63742 1 11187
2 63743 1 11187
2 63744 1 11187
2 63745 1 11187
2 63746 1 11187
2 63747 1 11189
2 63748 1 11189
2 63749 1 11191
2 63750 1 11191
2 63751 1 11191
2 63752 1 11191
2 63753 1 11191
2 63754 1 11191
2 63755 1 11191
2 63756 1 11191
2 63757 1 11192
2 63758 1 11192
2 63759 1 11192
2 63760 1 11192
2 63761 1 11192
2 63762 1 11193
2 63763 1 11193
2 63764 1 11204
2 63765 1 11204
2 63766 1 11204
2 63767 1 11204
2 63768 1 11204
2 63769 1 11204
2 63770 1 11206
2 63771 1 11206
2 63772 1 11208
2 63773 1 11208
2 63774 1 11216
2 63775 1 11216
2 63776 1 11218
2 63777 1 11218
2 63778 1 11218
2 63779 1 11226
2 63780 1 11226
2 63781 1 11226
2 63782 1 11235
2 63783 1 11235
2 63784 1 11235
2 63785 1 11235
2 63786 1 11235
2 63787 1 11235
2 63788 1 11236
2 63789 1 11236
2 63790 1 11236
2 63791 1 11243
2 63792 1 11243
2 63793 1 11245
2 63794 1 11245
2 63795 1 11245
2 63796 1 11245
2 63797 1 11245
2 63798 1 11245
2 63799 1 11245
2 63800 1 11245
2 63801 1 11245
2 63802 1 11245
2 63803 1 11245
2 63804 1 11245
2 63805 1 11245
2 63806 1 11246
2 63807 1 11246
2 63808 1 11246
2 63809 1 11246
2 63810 1 11246
2 63811 1 11247
2 63812 1 11247
2 63813 1 11255
2 63814 1 11255
2 63815 1 11255
2 63816 1 11255
2 63817 1 11255
2 63818 1 11256
2 63819 1 11256
2 63820 1 11264
2 63821 1 11264
2 63822 1 11264
2 63823 1 11269
2 63824 1 11269
2 63825 1 11273
2 63826 1 11273
2 63827 1 11273
2 63828 1 11273
2 63829 1 11273
2 63830 1 11273
2 63831 1 11273
2 63832 1 11273
2 63833 1 11273
2 63834 1 11273
2 63835 1 11273
2 63836 1 11273
2 63837 1 11273
2 63838 1 11273
2 63839 1 11286
2 63840 1 11286
2 63841 1 11287
2 63842 1 11287
2 63843 1 11287
2 63844 1 11288
2 63845 1 11288
2 63846 1 11296
2 63847 1 11296
2 63848 1 11297
2 63849 1 11297
2 63850 1 11297
2 63851 1 11300
2 63852 1 11300
2 63853 1 11300
2 63854 1 11300
2 63855 1 11300
2 63856 1 11300
2 63857 1 11300
2 63858 1 11300
2 63859 1 11302
2 63860 1 11302
2 63861 1 11302
2 63862 1 11304
2 63863 1 11304
2 63864 1 11323
2 63865 1 11323
2 63866 1 11323
2 63867 1 11324
2 63868 1 11324
2 63869 1 11325
2 63870 1 11325
2 63871 1 11343
2 63872 1 11343
2 63873 1 11343
2 63874 1 11345
2 63875 1 11345
2 63876 1 11350
2 63877 1 11350
2 63878 1 11366
2 63879 1 11366
2 63880 1 11380
2 63881 1 11380
2 63882 1 11381
2 63883 1 11381
2 63884 1 11381
2 63885 1 11389
2 63886 1 11389
2 63887 1 11406
2 63888 1 11406
2 63889 1 11428
2 63890 1 11428
2 63891 1 11428
2 63892 1 11430
2 63893 1 11430
2 63894 1 11431
2 63895 1 11431
2 63896 1 11431
2 63897 1 11431
2 63898 1 11431
2 63899 1 11431
2 63900 1 11432
2 63901 1 11432
2 63902 1 11440
2 63903 1 11440
2 63904 1 11440
2 63905 1 11449
2 63906 1 11449
2 63907 1 11450
2 63908 1 11450
2 63909 1 11450
2 63910 1 11450
2 63911 1 11451
2 63912 1 11451
2 63913 1 11453
2 63914 1 11453
2 63915 1 11453
2 63916 1 11453
2 63917 1 11453
2 63918 1 11453
2 63919 1 11453
2 63920 1 11461
2 63921 1 11461
2 63922 1 11473
2 63923 1 11473
2 63924 1 11474
2 63925 1 11474
2 63926 1 11474
2 63927 1 11475
2 63928 1 11475
2 63929 1 11483
2 63930 1 11483
2 63931 1 11501
2 63932 1 11501
2 63933 1 11501
2 63934 1 11501
2 63935 1 11501
2 63936 1 11501
2 63937 1 11501
2 63938 1 11501
2 63939 1 11501
2 63940 1 11501
2 63941 1 11501
2 63942 1 11501
2 63943 1 11501
2 63944 1 11501
2 63945 1 11501
2 63946 1 11501
2 63947 1 11501
2 63948 1 11501
2 63949 1 11501
2 63950 1 11501
2 63951 1 11501
2 63952 1 11510
2 63953 1 11510
2 63954 1 11510
2 63955 1 11510
2 63956 1 11510
2 63957 1 11510
2 63958 1 11510
2 63959 1 11511
2 63960 1 11511
2 63961 1 11511
2 63962 1 11512
2 63963 1 11512
2 63964 1 11513
2 63965 1 11513
2 63966 1 11520
2 63967 1 11520
2 63968 1 11520
2 63969 1 11521
2 63970 1 11521
2 63971 1 11521
2 63972 1 11521
2 63973 1 11530
2 63974 1 11530
2 63975 1 11538
2 63976 1 11538
2 63977 1 11538
2 63978 1 11538
2 63979 1 11538
2 63980 1 11541
2 63981 1 11541
2 63982 1 11550
2 63983 1 11550
2 63984 1 11550
2 63985 1 11553
2 63986 1 11553
2 63987 1 11564
2 63988 1 11564
2 63989 1 11585
2 63990 1 11585
2 63991 1 11585
2 63992 1 11585
2 63993 1 11585
2 63994 1 11585
2 63995 1 11585
2 63996 1 11585
2 63997 1 11585
2 63998 1 11585
2 63999 1 11585
2 64000 1 11585
2 64001 1 11585
2 64002 1 11585
2 64003 1 11585
2 64004 1 11585
2 64005 1 11585
2 64006 1 11585
2 64007 1 11585
2 64008 1 11586
2 64009 1 11586
2 64010 1 11586
2 64011 1 11586
2 64012 1 11596
2 64013 1 11596
2 64014 1 11596
2 64015 1 11596
2 64016 1 11597
2 64017 1 11597
2 64018 1 11611
2 64019 1 11611
2 64020 1 11611
2 64021 1 11611
2 64022 1 11611
2 64023 1 11611
2 64024 1 11611
2 64025 1 11611
2 64026 1 11611
2 64027 1 11611
2 64028 1 11611
2 64029 1 11611
2 64030 1 11611
2 64031 1 11611
2 64032 1 11620
2 64033 1 11620
2 64034 1 11620
2 64035 1 11621
2 64036 1 11621
2 64037 1 11621
2 64038 1 11621
2 64039 1 11623
2 64040 1 11623
2 64041 1 11624
2 64042 1 11624
2 64043 1 11640
2 64044 1 11640
2 64045 1 11640
2 64046 1 11641
2 64047 1 11641
2 64048 1 11641
2 64049 1 11641
2 64050 1 11641
2 64051 1 11641
2 64052 1 11641
2 64053 1 11641
2 64054 1 11649
2 64055 1 11649
2 64056 1 11649
2 64057 1 11665
2 64058 1 11665
2 64059 1 11665
2 64060 1 11667
2 64061 1 11667
2 64062 1 11672
2 64063 1 11672
2 64064 1 11679
2 64065 1 11679
2 64066 1 11679
2 64067 1 11679
2 64068 1 11680
2 64069 1 11680
2 64070 1 11680
2 64071 1 11680
2 64072 1 11700
2 64073 1 11700
2 64074 1 11700
2 64075 1 11700
2 64076 1 11700
2 64077 1 11700
2 64078 1 11700
2 64079 1 11700
2 64080 1 11700
2 64081 1 11700
2 64082 1 11700
2 64083 1 11702
2 64084 1 11702
2 64085 1 11704
2 64086 1 11704
2 64087 1 11708
2 64088 1 11708
2 64089 1 11708
2 64090 1 11709
2 64091 1 11709
2 64092 1 11709
2 64093 1 11709
2 64094 1 11709
2 64095 1 11709
2 64096 1 11719
2 64097 1 11719
2 64098 1 11719
2 64099 1 11719
2 64100 1 11719
2 64101 1 11719
2 64102 1 11719
2 64103 1 11719
2 64104 1 11719
2 64105 1 11719
2 64106 1 11719
2 64107 1 11724
2 64108 1 11724
2 64109 1 11724
2 64110 1 11724
2 64111 1 11724
2 64112 1 11724
2 64113 1 11724
2 64114 1 11724
2 64115 1 11724
2 64116 1 11724
2 64117 1 11724
2 64118 1 11724
2 64119 1 11724
2 64120 1 11724
2 64121 1 11724
2 64122 1 11724
2 64123 1 11724
2 64124 1 11724
2 64125 1 11727
2 64126 1 11727
2 64127 1 11727
2 64128 1 11728
2 64129 1 11728
2 64130 1 11736
2 64131 1 11736
2 64132 1 11736
2 64133 1 11736
2 64134 1 11748
2 64135 1 11748
2 64136 1 11752
2 64137 1 11752
2 64138 1 11761
2 64139 1 11761
2 64140 1 11761
2 64141 1 11763
2 64142 1 11763
2 64143 1 11763
2 64144 1 11763
2 64145 1 11764
2 64146 1 11764
2 64147 1 11774
2 64148 1 11774
2 64149 1 11775
2 64150 1 11775
2 64151 1 11786
2 64152 1 11786
2 64153 1 11799
2 64154 1 11799
2 64155 1 11814
2 64156 1 11814
2 64157 1 11815
2 64158 1 11815
2 64159 1 11837
2 64160 1 11837
2 64161 1 11849
2 64162 1 11849
2 64163 1 11864
2 64164 1 11864
2 64165 1 11892
2 64166 1 11892
2 64167 1 11892
2 64168 1 11899
2 64169 1 11899
2 64170 1 11926
2 64171 1 11926
2 64172 1 11931
2 64173 1 11931
2 64174 1 11932
2 64175 1 11932
2 64176 1 11933
2 64177 1 11933
2 64178 1 11945
2 64179 1 11945
2 64180 1 11946
2 64181 1 11946
2 64182 1 11951
2 64183 1 11951
2 64184 1 11963
2 64185 1 11963
2 64186 1 11972
2 64187 1 11972
2 64188 1 11984
2 64189 1 11984
2 64190 1 12037
2 64191 1 12037
2 64192 1 12038
2 64193 1 12038
2 64194 1 12038
2 64195 1 12038
2 64196 1 12038
2 64197 1 12038
2 64198 1 12038
2 64199 1 12038
2 64200 1 12038
2 64201 1 12041
2 64202 1 12041
2 64203 1 12042
2 64204 1 12042
2 64205 1 12064
2 64206 1 12064
2 64207 1 12071
2 64208 1 12071
2 64209 1 12071
2 64210 1 12071
2 64211 1 12071
2 64212 1 12071
2 64213 1 12071
2 64214 1 12083
2 64215 1 12083
2 64216 1 12086
2 64217 1 12086
2 64218 1 12110
2 64219 1 12110
2 64220 1 12123
2 64221 1 12123
2 64222 1 12137
2 64223 1 12137
2 64224 1 12141
2 64225 1 12141
2 64226 1 12151
2 64227 1 12151
2 64228 1 12151
2 64229 1 12151
2 64230 1 12151
2 64231 1 12167
2 64232 1 12167
2 64233 1 12167
2 64234 1 12167
2 64235 1 12167
2 64236 1 12170
2 64237 1 12170
2 64238 1 12170
2 64239 1 12170
2 64240 1 12170
2 64241 1 12170
2 64242 1 12171
2 64243 1 12171
2 64244 1 12173
2 64245 1 12173
2 64246 1 12187
2 64247 1 12187
2 64248 1 12187
2 64249 1 12187
2 64250 1 12193
2 64251 1 12193
2 64252 1 12213
2 64253 1 12213
2 64254 1 12220
2 64255 1 12220
2 64256 1 12221
2 64257 1 12221
2 64258 1 12238
2 64259 1 12238
2 64260 1 12238
2 64261 1 12238
2 64262 1 12238
2 64263 1 12246
2 64264 1 12246
2 64265 1 12246
2 64266 1 12246
2 64267 1 12250
2 64268 1 12250
2 64269 1 12256
2 64270 1 12256
2 64271 1 12293
2 64272 1 12293
2 64273 1 12294
2 64274 1 12294
2 64275 1 12295
2 64276 1 12295
2 64277 1 12295
2 64278 1 12295
2 64279 1 12325
2 64280 1 12325
2 64281 1 12345
2 64282 1 12345
2 64283 1 12345
2 64284 1 12361
2 64285 1 12361
2 64286 1 12361
2 64287 1 12372
2 64288 1 12372
2 64289 1 12372
2 64290 1 12372
2 64291 1 12384
2 64292 1 12384
2 64293 1 12388
2 64294 1 12388
2 64295 1 12443
2 64296 1 12443
2 64297 1 12443
2 64298 1 12444
2 64299 1 12444
2 64300 1 12444
2 64301 1 12444
2 64302 1 12444
2 64303 1 12444
2 64304 1 12444
2 64305 1 12444
2 64306 1 12444
2 64307 1 12444
2 64308 1 12444
2 64309 1 12444
2 64310 1 12444
2 64311 1 12444
2 64312 1 12446
2 64313 1 12446
2 64314 1 12447
2 64315 1 12447
2 64316 1 12447
2 64317 1 12447
2 64318 1 12447
2 64319 1 12453
2 64320 1 12453
2 64321 1 12467
2 64322 1 12467
2 64323 1 12478
2 64324 1 12478
2 64325 1 12478
2 64326 1 12521
2 64327 1 12521
2 64328 1 12521
2 64329 1 12521
2 64330 1 12521
2 64331 1 12530
2 64332 1 12530
2 64333 1 12530
2 64334 1 12531
2 64335 1 12531
2 64336 1 12531
2 64337 1 12531
2 64338 1 12549
2 64339 1 12549
2 64340 1 12549
2 64341 1 12552
2 64342 1 12552
2 64343 1 12570
2 64344 1 12570
2 64345 1 12570
2 64346 1 12584
2 64347 1 12584
2 64348 1 12584
2 64349 1 12606
2 64350 1 12606
2 64351 1 12607
2 64352 1 12607
2 64353 1 12607
2 64354 1 12607
2 64355 1 12607
2 64356 1 12608
2 64357 1 12608
2 64358 1 12616
2 64359 1 12616
2 64360 1 12616
2 64361 1 12636
2 64362 1 12636
2 64363 1 12636
2 64364 1 12637
2 64365 1 12637
2 64366 1 12637
2 64367 1 12637
2 64368 1 12637
2 64369 1 12637
2 64370 1 12637
2 64371 1 12637
2 64372 1 12637
2 64373 1 12650
2 64374 1 12650
2 64375 1 12650
2 64376 1 12650
2 64377 1 12651
2 64378 1 12651
2 64379 1 12664
2 64380 1 12664
2 64381 1 12665
2 64382 1 12665
2 64383 1 12665
2 64384 1 12665
2 64385 1 12668
2 64386 1 12668
2 64387 1 12669
2 64388 1 12669
2 64389 1 12669
2 64390 1 12669
2 64391 1 12669
2 64392 1 12684
2 64393 1 12684
2 64394 1 12684
2 64395 1 12684
2 64396 1 12684
2 64397 1 12684
2 64398 1 12684
2 64399 1 12684
2 64400 1 12684
2 64401 1 12684
2 64402 1 12684
2 64403 1 12684
2 64404 1 12684
2 64405 1 12685
2 64406 1 12685
2 64407 1 12686
2 64408 1 12686
2 64409 1 12686
2 64410 1 12701
2 64411 1 12701
2 64412 1 12702
2 64413 1 12702
2 64414 1 12710
2 64415 1 12710
2 64416 1 12718
2 64417 1 12718
2 64418 1 12718
2 64419 1 12718
2 64420 1 12720
2 64421 1 12720
2 64422 1 12720
2 64423 1 12720
2 64424 1 12720
2 64425 1 12720
2 64426 1 12794
2 64427 1 12794
2 64428 1 12794
2 64429 1 12794
2 64430 1 12794
2 64431 1 12794
2 64432 1 12794
2 64433 1 12794
2 64434 1 12794
2 64435 1 12794
2 64436 1 12812
2 64437 1 12812
2 64438 1 12812
2 64439 1 12812
2 64440 1 12812
2 64441 1 12820
2 64442 1 12820
2 64443 1 12820
2 64444 1 12820
2 64445 1 12820
2 64446 1 12820
2 64447 1 12820
2 64448 1 12823
2 64449 1 12823
2 64450 1 12852
2 64451 1 12852
2 64452 1 12852
2 64453 1 12852
2 64454 1 12861
2 64455 1 12861
2 64456 1 12861
2 64457 1 12870
2 64458 1 12870
2 64459 1 12870
2 64460 1 12870
2 64461 1 12870
2 64462 1 12870
2 64463 1 12870
2 64464 1 12870
2 64465 1 12870
2 64466 1 12870
2 64467 1 12870
2 64468 1 12870
2 64469 1 12870
2 64470 1 12871
2 64471 1 12871
2 64472 1 12889
2 64473 1 12889
2 64474 1 12889
2 64475 1 12900
2 64476 1 12900
2 64477 1 12904
2 64478 1 12904
2 64479 1 12905
2 64480 1 12905
2 64481 1 12913
2 64482 1 12913
2 64483 1 12930
2 64484 1 12930
2 64485 1 12930
2 64486 1 12945
2 64487 1 12945
2 64488 1 12945
2 64489 1 12945
2 64490 1 12945
2 64491 1 12945
2 64492 1 12946
2 64493 1 12946
2 64494 1 12947
2 64495 1 12947
2 64496 1 12947
2 64497 1 12947
2 64498 1 12948
2 64499 1 12948
2 64500 1 12948
2 64501 1 12948
2 64502 1 12948
2 64503 1 12948
2 64504 1 12948
2 64505 1 12948
2 64506 1 12972
2 64507 1 12972
2 64508 1 12972
2 64509 1 12972
2 64510 1 12986
2 64511 1 12986
2 64512 1 12994
2 64513 1 12994
2 64514 1 13015
2 64515 1 13015
2 64516 1 13033
2 64517 1 13033
2 64518 1 13033
2 64519 1 13034
2 64520 1 13034
2 64521 1 13045
2 64522 1 13045
2 64523 1 13045
2 64524 1 13045
2 64525 1 13045
2 64526 1 13045
2 64527 1 13045
2 64528 1 13045
2 64529 1 13045
2 64530 1 13045
2 64531 1 13045
2 64532 1 13045
2 64533 1 13046
2 64534 1 13046
2 64535 1 13047
2 64536 1 13047
2 64537 1 13050
2 64538 1 13050
2 64539 1 13050
2 64540 1 13050
2 64541 1 13050
2 64542 1 13050
2 64543 1 13051
2 64544 1 13051
2 64545 1 13051
2 64546 1 13065
2 64547 1 13065
2 64548 1 13066
2 64549 1 13066
2 64550 1 13066
2 64551 1 13066
2 64552 1 13066
2 64553 1 13066
2 64554 1 13066
2 64555 1 13066
2 64556 1 13066
2 64557 1 13066
2 64558 1 13066
2 64559 1 13067
2 64560 1 13067
2 64561 1 13067
2 64562 1 13068
2 64563 1 13068
2 64564 1 13069
2 64565 1 13069
2 64566 1 13069
2 64567 1 13069
2 64568 1 13070
2 64569 1 13070
2 64570 1 13074
2 64571 1 13074
2 64572 1 13083
2 64573 1 13083
2 64574 1 13084
2 64575 1 13084
2 64576 1 13084
2 64577 1 13084
2 64578 1 13084
2 64579 1 13102
2 64580 1 13102
2 64581 1 13120
2 64582 1 13120
2 64583 1 13128
2 64584 1 13128
2 64585 1 13132
2 64586 1 13132
2 64587 1 13132
2 64588 1 13132
2 64589 1 13132
2 64590 1 13132
2 64591 1 13134
2 64592 1 13134
2 64593 1 13135
2 64594 1 13135
2 64595 1 13151
2 64596 1 13151
2 64597 1 13151
2 64598 1 13151
2 64599 1 13151
2 64600 1 13151
2 64601 1 13151
2 64602 1 13152
2 64603 1 13152
2 64604 1 13159
2 64605 1 13159
2 64606 1 13159
2 64607 1 13159
2 64608 1 13171
2 64609 1 13171
2 64610 1 13182
2 64611 1 13182
2 64612 1 13183
2 64613 1 13183
2 64614 1 13184
2 64615 1 13184
2 64616 1 13184
2 64617 1 13184
2 64618 1 13184
2 64619 1 13184
2 64620 1 13184
2 64621 1 13184
2 64622 1 13184
2 64623 1 13184
2 64624 1 13184
2 64625 1 13184
2 64626 1 13218
2 64627 1 13218
2 64628 1 13235
2 64629 1 13235
2 64630 1 13238
2 64631 1 13238
2 64632 1 13239
2 64633 1 13239
2 64634 1 13239
2 64635 1 13243
2 64636 1 13243
2 64637 1 13243
2 64638 1 13243
2 64639 1 13252
2 64640 1 13252
2 64641 1 13253
2 64642 1 13253
2 64643 1 13255
2 64644 1 13255
2 64645 1 13255
2 64646 1 13255
2 64647 1 13255
2 64648 1 13255
2 64649 1 13255
2 64650 1 13256
2 64651 1 13256
2 64652 1 13263
2 64653 1 13263
2 64654 1 13263
2 64655 1 13263
2 64656 1 13265
2 64657 1 13265
2 64658 1 13265
2 64659 1 13283
2 64660 1 13283
2 64661 1 13283
2 64662 1 13284
2 64663 1 13284
2 64664 1 13284
2 64665 1 13284
2 64666 1 13284
2 64667 1 13302
2 64668 1 13302
2 64669 1 13302
2 64670 1 13302
2 64671 1 13302
2 64672 1 13354
2 64673 1 13354
2 64674 1 13354
2 64675 1 13354
2 64676 1 13407
2 64677 1 13407
2 64678 1 13421
2 64679 1 13421
2 64680 1 13421
2 64681 1 13421
2 64682 1 13421
2 64683 1 13421
2 64684 1 13421
2 64685 1 13421
2 64686 1 13421
2 64687 1 13421
2 64688 1 13421
2 64689 1 13421
2 64690 1 13421
2 64691 1 13421
2 64692 1 13421
2 64693 1 13421
2 64694 1 13421
2 64695 1 13421
2 64696 1 13421
2 64697 1 13421
2 64698 1 13422
2 64699 1 13422
2 64700 1 13422
2 64701 1 13422
2 64702 1 13441
2 64703 1 13441
2 64704 1 13442
2 64705 1 13442
2 64706 1 13481
2 64707 1 13481
2 64708 1 13481
2 64709 1 13489
2 64710 1 13489
2 64711 1 13497
2 64712 1 13497
2 64713 1 13497
2 64714 1 13497
2 64715 1 13497
2 64716 1 13497
2 64717 1 13497
2 64718 1 13497
2 64719 1 13497
2 64720 1 13497
2 64721 1 13497
2 64722 1 13497
2 64723 1 13497
2 64724 1 13516
2 64725 1 13516
2 64726 1 13516
2 64727 1 13516
2 64728 1 13516
2 64729 1 13516
2 64730 1 13516
2 64731 1 13539
2 64732 1 13539
2 64733 1 13555
2 64734 1 13555
2 64735 1 13556
2 64736 1 13556
2 64737 1 13559
2 64738 1 13559
2 64739 1 13559
2 64740 1 13559
2 64741 1 13559
2 64742 1 13584
2 64743 1 13584
2 64744 1 13584
2 64745 1 13599
2 64746 1 13599
2 64747 1 13611
2 64748 1 13611
2 64749 1 13611
2 64750 1 13611
2 64751 1 13611
2 64752 1 13611
2 64753 1 13611
2 64754 1 13611
2 64755 1 13611
2 64756 1 13611
2 64757 1 13611
2 64758 1 13611
2 64759 1 13611
2 64760 1 13611
2 64761 1 13612
2 64762 1 13612
2 64763 1 13612
2 64764 1 13612
2 64765 1 13612
2 64766 1 13612
2 64767 1 13617
2 64768 1 13617
2 64769 1 13643
2 64770 1 13643
2 64771 1 13643
2 64772 1 13652
2 64773 1 13652
2 64774 1 13652
2 64775 1 13652
2 64776 1 13653
2 64777 1 13653
2 64778 1 13677
2 64779 1 13677
2 64780 1 13677
2 64781 1 13697
2 64782 1 13697
2 64783 1 13720
2 64784 1 13720
2 64785 1 13735
2 64786 1 13735
2 64787 1 13742
2 64788 1 13742
2 64789 1 13742
2 64790 1 13743
2 64791 1 13743
2 64792 1 13746
2 64793 1 13746
2 64794 1 13747
2 64795 1 13747
2 64796 1 13749
2 64797 1 13749
2 64798 1 13753
2 64799 1 13753
2 64800 1 13764
2 64801 1 13764
2 64802 1 13779
2 64803 1 13779
2 64804 1 13798
2 64805 1 13798
2 64806 1 13803
2 64807 1 13803
2 64808 1 13810
2 64809 1 13810
2 64810 1 13820
2 64811 1 13820
2 64812 1 13820
2 64813 1 13830
2 64814 1 13830
2 64815 1 13846
2 64816 1 13846
2 64817 1 13846
2 64818 1 13846
2 64819 1 13846
2 64820 1 13846
2 64821 1 13846
2 64822 1 13846
2 64823 1 13861
2 64824 1 13861
2 64825 1 13873
2 64826 1 13873
2 64827 1 13883
2 64828 1 13883
2 64829 1 13902
2 64830 1 13902
2 64831 1 13919
2 64832 1 13919
2 64833 1 13923
2 64834 1 13923
2 64835 1 13923
2 64836 1 13957
2 64837 1 13957
2 64838 1 13957
2 64839 1 13958
2 64840 1 13958
2 64841 1 13963
2 64842 1 13963
2 64843 1 13969
2 64844 1 13969
2 64845 1 13972
2 64846 1 13972
2 64847 1 13972
2 64848 1 13973
2 64849 1 13973
2 64850 1 13974
2 64851 1 13974
2 64852 1 13990
2 64853 1 13990
2 64854 1 13995
2 64855 1 13995
2 64856 1 13995
2 64857 1 13995
2 64858 1 14003
2 64859 1 14003
2 64860 1 14003
2 64861 1 14025
2 64862 1 14025
2 64863 1 14054
2 64864 1 14054
2 64865 1 14076
2 64866 1 14076
2 64867 1 14076
2 64868 1 14076
2 64869 1 14094
2 64870 1 14094
2 64871 1 14098
2 64872 1 14098
2 64873 1 14104
2 64874 1 14104
2 64875 1 14117
2 64876 1 14117
2 64877 1 14117
2 64878 1 14118
2 64879 1 14118
2 64880 1 14118
2 64881 1 14118
2 64882 1 14118
2 64883 1 14118
2 64884 1 14118
2 64885 1 14132
2 64886 1 14132
2 64887 1 14133
2 64888 1 14133
2 64889 1 14151
2 64890 1 14151
2 64891 1 14154
2 64892 1 14154
2 64893 1 14166
2 64894 1 14166
2 64895 1 14166
2 64896 1 14169
2 64897 1 14169
2 64898 1 14177
2 64899 1 14177
2 64900 1 14177
2 64901 1 14178
2 64902 1 14178
2 64903 1 14178
2 64904 1 14179
2 64905 1 14179
2 64906 1 14179
2 64907 1 14179
2 64908 1 14190
2 64909 1 14190
2 64910 1 14190
2 64911 1 14190
2 64912 1 14209
2 64913 1 14209
2 64914 1 14209
2 64915 1 14209
2 64916 1 14209
2 64917 1 14209
2 64918 1 14210
2 64919 1 14210
2 64920 1 14219
2 64921 1 14219
2 64922 1 14219
2 64923 1 14219
2 64924 1 14219
2 64925 1 14227
2 64926 1 14227
2 64927 1 14231
2 64928 1 14231
2 64929 1 14233
2 64930 1 14233
2 64931 1 14233
2 64932 1 14254
2 64933 1 14254
2 64934 1 14257
2 64935 1 14257
2 64936 1 14257
2 64937 1 14257
2 64938 1 14257
2 64939 1 14257
2 64940 1 14257
2 64941 1 14257
2 64942 1 14257
2 64943 1 14257
2 64944 1 14257
2 64945 1 14257
2 64946 1 14257
2 64947 1 14258
2 64948 1 14258
2 64949 1 14258
2 64950 1 14258
2 64951 1 14258
2 64952 1 14258
2 64953 1 14272
2 64954 1 14272
2 64955 1 14275
2 64956 1 14275
2 64957 1 14275
2 64958 1 14275
2 64959 1 14275
2 64960 1 14275
2 64961 1 14275
2 64962 1 14276
2 64963 1 14276
2 64964 1 14277
2 64965 1 14277
2 64966 1 14282
2 64967 1 14282
2 64968 1 14285
2 64969 1 14285
2 64970 1 14285
2 64971 1 14286
2 64972 1 14286
2 64973 1 14286
2 64974 1 14286
2 64975 1 14287
2 64976 1 14287
2 64977 1 14287
2 64978 1 14287
2 64979 1 14287
2 64980 1 14287
2 64981 1 14287
2 64982 1 14289
2 64983 1 14289
2 64984 1 14296
2 64985 1 14296
2 64986 1 14296
2 64987 1 14296
2 64988 1 14296
2 64989 1 14297
2 64990 1 14297
2 64991 1 14298
2 64992 1 14298
2 64993 1 14309
2 64994 1 14309
2 64995 1 14309
2 64996 1 14309
2 64997 1 14309
2 64998 1 14309
2 64999 1 14309
2 65000 1 14313
2 65001 1 14313
2 65002 1 14322
2 65003 1 14322
2 65004 1 14326
2 65005 1 14326
2 65006 1 14326
2 65007 1 14327
2 65008 1 14327
2 65009 1 14327
2 65010 1 14328
2 65011 1 14328
2 65012 1 14330
2 65013 1 14330
2 65014 1 14330
2 65015 1 14330
2 65016 1 14330
2 65017 1 14330
2 65018 1 14342
2 65019 1 14342
2 65020 1 14345
2 65021 1 14345
2 65022 1 14345
2 65023 1 14345
2 65024 1 14345
2 65025 1 14345
2 65026 1 14345
2 65027 1 14345
2 65028 1 14346
2 65029 1 14346
2 65030 1 14346
2 65031 1 14354
2 65032 1 14354
2 65033 1 14354
2 65034 1 14366
2 65035 1 14366
2 65036 1 14417
2 65037 1 14417
2 65038 1 14417
2 65039 1 14421
2 65040 1 14421
2 65041 1 14421
2 65042 1 14422
2 65043 1 14422
2 65044 1 14440
2 65045 1 14440
2 65046 1 14440
2 65047 1 14440
2 65048 1 14440
2 65049 1 14440
2 65050 1 14440
2 65051 1 14441
2 65052 1 14441
2 65053 1 14443
2 65054 1 14443
2 65055 1 14443
2 65056 1 14466
2 65057 1 14466
2 65058 1 14480
2 65059 1 14480
2 65060 1 14492
2 65061 1 14492
2 65062 1 14527
2 65063 1 14527
2 65064 1 14527
2 65065 1 14527
2 65066 1 14527
2 65067 1 14528
2 65068 1 14528
2 65069 1 14528
2 65070 1 14528
2 65071 1 14540
2 65072 1 14540
2 65073 1 14540
2 65074 1 14543
2 65075 1 14543
2 65076 1 14543
2 65077 1 14543
2 65078 1 14543
2 65079 1 14543
2 65080 1 14543
2 65081 1 14543
2 65082 1 14543
2 65083 1 14543
2 65084 1 14544
2 65085 1 14544
2 65086 1 14546
2 65087 1 14546
2 65088 1 14579
2 65089 1 14579
2 65090 1 14628
2 65091 1 14628
2 65092 1 14637
2 65093 1 14637
2 65094 1 14670
2 65095 1 14670
2 65096 1 14671
2 65097 1 14671
2 65098 1 14698
2 65099 1 14698
2 65100 1 14715
2 65101 1 14715
2 65102 1 14758
2 65103 1 14758
2 65104 1 14813
2 65105 1 14813
2 65106 1 14816
2 65107 1 14816
2 65108 1 14842
2 65109 1 14842
2 65110 1 14847
2 65111 1 14847
2 65112 1 14861
2 65113 1 14861
2 65114 1 14862
2 65115 1 14862
2 65116 1 14862
2 65117 1 14871
2 65118 1 14871
2 65119 1 14871
2 65120 1 14871
2 65121 1 14883
2 65122 1 14883
2 65123 1 14897
2 65124 1 14897
2 65125 1 14897
2 65126 1 14897
2 65127 1 14897
2 65128 1 14901
2 65129 1 14901
2 65130 1 14901
2 65131 1 14925
2 65132 1 14925
2 65133 1 14925
2 65134 1 14933
2 65135 1 14933
2 65136 1 14952
2 65137 1 14952
2 65138 1 14954
2 65139 1 14954
2 65140 1 14957
2 65141 1 14957
2 65142 1 14962
2 65143 1 14962
2 65144 1 14976
2 65145 1 14976
2 65146 1 14984
2 65147 1 14984
2 65148 1 15016
2 65149 1 15016
2 65150 1 15037
2 65151 1 15037
2 65152 1 15037
2 65153 1 15046
2 65154 1 15046
2 65155 1 15054
2 65156 1 15054
2 65157 1 15056
2 65158 1 15056
2 65159 1 15056
2 65160 1 15056
2 65161 1 15056
2 65162 1 15059
2 65163 1 15059
2 65164 1 15059
2 65165 1 15059
2 65166 1 15059
2 65167 1 15063
2 65168 1 15063
2 65169 1 15064
2 65170 1 15064
2 65171 1 15087
2 65172 1 15087
2 65173 1 15087
2 65174 1 15087
2 65175 1 15087
2 65176 1 15087
2 65177 1 15087
2 65178 1 15087
2 65179 1 15087
2 65180 1 15088
2 65181 1 15088
2 65182 1 15095
2 65183 1 15095
2 65184 1 15095
2 65185 1 15143
2 65186 1 15143
2 65187 1 15144
2 65188 1 15144
2 65189 1 15151
2 65190 1 15151
2 65191 1 15183
2 65192 1 15183
2 65193 1 15184
2 65194 1 15184
2 65195 1 15185
2 65196 1 15185
2 65197 1 15185
2 65198 1 15195
2 65199 1 15195
2 65200 1 15200
2 65201 1 15200
2 65202 1 15200
2 65203 1 15203
2 65204 1 15203
2 65205 1 15208
2 65206 1 15208
2 65207 1 15228
2 65208 1 15228
2 65209 1 15228
2 65210 1 15263
2 65211 1 15263
2 65212 1 15285
2 65213 1 15285
2 65214 1 15285
2 65215 1 15285
2 65216 1 15285
2 65217 1 15302
2 65218 1 15302
2 65219 1 15310
2 65220 1 15310
2 65221 1 15310
2 65222 1 15310
2 65223 1 15313
2 65224 1 15313
2 65225 1 15313
2 65226 1 15314
2 65227 1 15314
2 65228 1 15320
2 65229 1 15320
2 65230 1 15321
2 65231 1 15321
2 65232 1 15332
2 65233 1 15332
2 65234 1 15345
2 65235 1 15345
2 65236 1 15346
2 65237 1 15346
2 65238 1 15348
2 65239 1 15348
2 65240 1 15379
2 65241 1 15379
2 65242 1 15428
2 65243 1 15428
2 65244 1 15443
2 65245 1 15443
2 65246 1 15461
2 65247 1 15461
2 65248 1 15461
2 65249 1 15461
2 65250 1 15461
2 65251 1 15461
2 65252 1 15463
2 65253 1 15463
2 65254 1 15463
2 65255 1 15463
2 65256 1 15465
2 65257 1 15465
2 65258 1 15467
2 65259 1 15467
2 65260 1 15473
2 65261 1 15473
2 65262 1 15473
2 65263 1 15473
2 65264 1 15473
2 65265 1 15475
2 65266 1 15475
2 65267 1 15482
2 65268 1 15482
2 65269 1 15499
2 65270 1 15499
2 65271 1 15500
2 65272 1 15500
2 65273 1 15501
2 65274 1 15501
2 65275 1 15502
2 65276 1 15502
2 65277 1 15537
2 65278 1 15537
2 65279 1 15537
2 65280 1 15537
2 65281 1 15550
2 65282 1 15550
2 65283 1 15554
2 65284 1 15554
2 65285 1 15568
2 65286 1 15568
2 65287 1 15568
2 65288 1 15570
2 65289 1 15570
2 65290 1 15570
2 65291 1 15570
2 65292 1 15570
2 65293 1 15570
2 65294 1 15578
2 65295 1 15578
2 65296 1 15578
2 65297 1 15578
2 65298 1 15580
2 65299 1 15580
2 65300 1 15580
2 65301 1 15580
2 65302 1 15580
2 65303 1 15580
2 65304 1 15580
2 65305 1 15580
2 65306 1 15600
2 65307 1 15600
2 65308 1 15601
2 65309 1 15601
2 65310 1 15613
2 65311 1 15613
2 65312 1 15620
2 65313 1 15620
2 65314 1 15632
2 65315 1 15632
2 65316 1 15632
2 65317 1 15632
2 65318 1 15632
2 65319 1 15670
2 65320 1 15670
2 65321 1 15686
2 65322 1 15686
2 65323 1 15692
2 65324 1 15692
2 65325 1 15693
2 65326 1 15693
2 65327 1 15696
2 65328 1 15696
2 65329 1 15696
2 65330 1 15729
2 65331 1 15729
2 65332 1 15735
2 65333 1 15735
2 65334 1 15735
2 65335 1 15735
2 65336 1 15738
2 65337 1 15738
2 65338 1 15738
2 65339 1 15738
2 65340 1 15738
2 65341 1 15738
2 65342 1 15739
2 65343 1 15739
2 65344 1 15741
2 65345 1 15741
2 65346 1 15741
2 65347 1 15741
2 65348 1 15798
2 65349 1 15798
2 65350 1 15799
2 65351 1 15799
2 65352 1 15844
2 65353 1 15844
2 65354 1 15844
2 65355 1 15850
2 65356 1 15850
2 65357 1 15850
2 65358 1 15857
2 65359 1 15857
2 65360 1 15858
2 65361 1 15858
2 65362 1 15858
2 65363 1 15858
2 65364 1 15858
2 65365 1 15858
2 65366 1 15887
2 65367 1 15887
2 65368 1 15887
2 65369 1 15888
2 65370 1 15888
2 65371 1 15917
2 65372 1 15917
2 65373 1 15917
2 65374 1 15917
2 65375 1 15933
2 65376 1 15933
2 65377 1 15946
2 65378 1 15946
2 65379 1 15991
2 65380 1 15991
2 65381 1 16084
2 65382 1 16084
2 65383 1 16084
2 65384 1 16085
2 65385 1 16085
2 65386 1 16098
2 65387 1 16098
2 65388 1 16098
2 65389 1 16101
2 65390 1 16101
2 65391 1 16132
2 65392 1 16132
2 65393 1 16141
2 65394 1 16141
2 65395 1 16164
2 65396 1 16164
2 65397 1 16164
2 65398 1 16175
2 65399 1 16175
2 65400 1 16175
2 65401 1 16176
2 65402 1 16176
2 65403 1 16184
2 65404 1 16184
2 65405 1 16199
2 65406 1 16199
2 65407 1 16206
2 65408 1 16206
2 65409 1 16206
2 65410 1 16206
2 65411 1 16238
2 65412 1 16238
2 65413 1 16255
2 65414 1 16255
2 65415 1 16258
2 65416 1 16258
2 65417 1 16259
2 65418 1 16259
2 65419 1 16259
2 65420 1 16277
2 65421 1 16277
2 65422 1 16277
2 65423 1 16297
2 65424 1 16297
2 65425 1 16297
2 65426 1 16297
2 65427 1 16297
2 65428 1 16297
2 65429 1 16298
2 65430 1 16298
2 65431 1 16303
2 65432 1 16303
2 65433 1 16303
2 65434 1 16303
2 65435 1 16319
2 65436 1 16319
2 65437 1 16327
2 65438 1 16327
2 65439 1 16366
2 65440 1 16366
2 65441 1 16393
2 65442 1 16393
2 65443 1 16394
2 65444 1 16394
2 65445 1 16395
2 65446 1 16395
2 65447 1 16395
2 65448 1 16397
2 65449 1 16397
2 65450 1 16397
2 65451 1 16397
2 65452 1 16400
2 65453 1 16400
2 65454 1 16401
2 65455 1 16401
2 65456 1 16404
2 65457 1 16404
2 65458 1 16404
2 65459 1 16405
2 65460 1 16405
2 65461 1 16405
2 65462 1 16406
2 65463 1 16406
2 65464 1 16406
2 65465 1 16421
2 65466 1 16421
2 65467 1 16422
2 65468 1 16422
2 65469 1 16422
2 65470 1 16422
2 65471 1 16422
2 65472 1 16422
2 65473 1 16424
2 65474 1 16424
2 65475 1 16442
2 65476 1 16442
2 65477 1 16443
2 65478 1 16443
2 65479 1 16480
2 65480 1 16480
2 65481 1 16480
2 65482 1 16480
2 65483 1 16483
2 65484 1 16483
2 65485 1 16486
2 65486 1 16486
2 65487 1 16486
2 65488 1 16486
2 65489 1 16486
2 65490 1 16486
2 65491 1 16487
2 65492 1 16487
2 65493 1 16491
2 65494 1 16491
2 65495 1 16491
2 65496 1 16491
2 65497 1 16491
2 65498 1 16492
2 65499 1 16492
2 65500 1 16492
2 65501 1 16492
2 65502 1 16526
2 65503 1 16526
2 65504 1 16527
2 65505 1 16527
2 65506 1 16528
2 65507 1 16528
2 65508 1 16529
2 65509 1 16529
2 65510 1 16553
2 65511 1 16553
2 65512 1 16553
2 65513 1 16553
2 65514 1 16592
2 65515 1 16592
2 65516 1 16592
2 65517 1 16592
2 65518 1 16609
2 65519 1 16609
2 65520 1 16609
2 65521 1 16612
2 65522 1 16612
2 65523 1 16612
2 65524 1 16614
2 65525 1 16614
2 65526 1 16614
2 65527 1 16617
2 65528 1 16617
2 65529 1 16617
2 65530 1 16617
2 65531 1 16617
2 65532 1 16617
2 65533 1 16620
2 65534 1 16620
2 65535 1 16621
2 65536 1 16621
2 65537 1 16621
2 65538 1 16621
2 65539 1 16621
2 65540 1 16621
2 65541 1 16621
2 65542 1 16621
2 65543 1 16621
2 65544 1 16621
2 65545 1 16621
2 65546 1 16621
2 65547 1 16629
2 65548 1 16629
2 65549 1 16630
2 65550 1 16630
2 65551 1 16630
2 65552 1 16647
2 65553 1 16647
2 65554 1 16674
2 65555 1 16674
2 65556 1 16677
2 65557 1 16677
2 65558 1 16678
2 65559 1 16678
2 65560 1 16678
2 65561 1 16684
2 65562 1 16684
2 65563 1 16690
2 65564 1 16690
2 65565 1 16690
2 65566 1 16691
2 65567 1 16691
2 65568 1 16706
2 65569 1 16706
2 65570 1 16709
2 65571 1 16709
2 65572 1 16709
2 65573 1 16709
2 65574 1 16709
2 65575 1 16709
2 65576 1 16710
2 65577 1 16710
2 65578 1 16710
2 65579 1 16710
2 65580 1 16736
2 65581 1 16736
2 65582 1 16736
2 65583 1 16739
2 65584 1 16739
2 65585 1 16739
2 65586 1 16739
2 65587 1 16739
2 65588 1 16739
2 65589 1 16739
2 65590 1 16769
2 65591 1 16769
2 65592 1 16802
2 65593 1 16802
2 65594 1 16808
2 65595 1 16808
2 65596 1 16813
2 65597 1 16813
2 65598 1 16829
2 65599 1 16829
2 65600 1 16843
2 65601 1 16843
2 65602 1 16844
2 65603 1 16844
2 65604 1 16849
2 65605 1 16849
2 65606 1 16849
2 65607 1 16852
2 65608 1 16852
2 65609 1 16857
2 65610 1 16857
2 65611 1 16857
2 65612 1 16857
2 65613 1 16857
2 65614 1 16858
2 65615 1 16858
2 65616 1 16858
2 65617 1 16859
2 65618 1 16859
2 65619 1 16859
2 65620 1 16859
2 65621 1 16859
2 65622 1 16859
2 65623 1 16859
2 65624 1 16859
2 65625 1 16859
2 65626 1 16860
2 65627 1 16860
2 65628 1 16893
2 65629 1 16893
2 65630 1 16893
2 65631 1 16894
2 65632 1 16894
2 65633 1 16897
2 65634 1 16897
2 65635 1 16910
2 65636 1 16910
2 65637 1 16911
2 65638 1 16911
2 65639 1 16911
2 65640 1 16922
2 65641 1 16922
2 65642 1 16922
2 65643 1 16922
2 65644 1 16923
2 65645 1 16923
2 65646 1 16923
2 65647 1 16923
2 65648 1 16923
2 65649 1 16931
2 65650 1 16931
2 65651 1 16954
2 65652 1 16954
2 65653 1 16954
2 65654 1 16963
2 65655 1 16963
2 65656 1 16978
2 65657 1 16978
2 65658 1 16978
2 65659 1 16998
2 65660 1 16998
2 65661 1 16998
2 65662 1 16998
2 65663 1 16998
2 65664 1 16998
2 65665 1 16998
2 65666 1 16999
2 65667 1 16999
2 65668 1 16999
2 65669 1 16999
2 65670 1 17014
2 65671 1 17014
2 65672 1 17014
2 65673 1 17017
2 65674 1 17017
2 65675 1 17017
2 65676 1 17017
2 65677 1 17017
2 65678 1 17018
2 65679 1 17018
2 65680 1 17018
2 65681 1 17018
2 65682 1 17018
2 65683 1 17018
2 65684 1 17018
2 65685 1 17018
2 65686 1 17018
2 65687 1 17018
2 65688 1 17018
2 65689 1 17018
2 65690 1 17018
2 65691 1 17018
2 65692 1 17018
2 65693 1 17018
2 65694 1 17018
2 65695 1 17018
2 65696 1 17018
2 65697 1 17018
2 65698 1 17018
2 65699 1 17018
2 65700 1 17018
2 65701 1 17018
2 65702 1 17018
2 65703 1 17018
2 65704 1 17018
2 65705 1 17018
2 65706 1 17018
2 65707 1 17018
2 65708 1 17018
2 65709 1 17018
2 65710 1 17018
2 65711 1 17018
2 65712 1 17018
2 65713 1 17018
2 65714 1 17018
2 65715 1 17018
2 65716 1 17018
2 65717 1 17018
2 65718 1 17018
2 65719 1 17018
2 65720 1 17018
2 65721 1 17018
2 65722 1 17018
2 65723 1 17018
2 65724 1 17018
2 65725 1 17018
2 65726 1 17018
2 65727 1 17018
2 65728 1 17018
2 65729 1 17018
2 65730 1 17018
2 65731 1 17018
2 65732 1 17018
2 65733 1 17018
2 65734 1 17018
2 65735 1 17018
2 65736 1 17018
2 65737 1 17018
2 65738 1 17018
2 65739 1 17018
2 65740 1 17018
2 65741 1 17018
2 65742 1 17018
2 65743 1 17018
2 65744 1 17018
2 65745 1 17018
2 65746 1 17018
2 65747 1 17018
2 65748 1 17018
2 65749 1 17018
2 65750 1 17018
2 65751 1 17018
2 65752 1 17018
2 65753 1 17018
2 65754 1 17018
2 65755 1 17018
2 65756 1 17018
2 65757 1 17018
2 65758 1 17018
2 65759 1 17018
2 65760 1 17018
2 65761 1 17018
2 65762 1 17018
2 65763 1 17018
2 65764 1 17018
2 65765 1 17018
2 65766 1 17018
2 65767 1 17018
2 65768 1 17018
2 65769 1 17018
2 65770 1 17018
2 65771 1 17018
2 65772 1 17018
2 65773 1 17018
2 65774 1 17018
2 65775 1 17018
2 65776 1 17018
2 65777 1 17018
2 65778 1 17018
2 65779 1 17018
2 65780 1 17018
2 65781 1 17018
2 65782 1 17018
2 65783 1 17018
2 65784 1 17018
2 65785 1 17019
2 65786 1 17019
2 65787 1 17019
2 65788 1 17019
2 65789 1 17019
2 65790 1 17019
2 65791 1 17019
2 65792 1 17019
2 65793 1 17022
2 65794 1 17022
2 65795 1 17026
2 65796 1 17026
2 65797 1 17029
2 65798 1 17029
2 65799 1 17029
2 65800 1 17030
2 65801 1 17030
2 65802 1 17030
2 65803 1 17030
2 65804 1 17030
2 65805 1 17033
2 65806 1 17033
2 65807 1 17033
2 65808 1 17033
2 65809 1 17033
2 65810 1 17033
2 65811 1 17033
2 65812 1 17036
2 65813 1 17036
2 65814 1 17036
2 65815 1 17036
2 65816 1 17037
2 65817 1 17037
2 65818 1 17038
2 65819 1 17038
2 65820 1 17038
2 65821 1 17038
2 65822 1 17039
2 65823 1 17039
2 65824 1 17041
2 65825 1 17041
2 65826 1 17049
2 65827 1 17049
2 65828 1 17049
2 65829 1 17049
2 65830 1 17049
2 65831 1 17049
2 65832 1 17049
2 65833 1 17049
2 65834 1 17049
2 65835 1 17049
2 65836 1 17049
2 65837 1 17049
2 65838 1 17050
2 65839 1 17050
2 65840 1 17050
2 65841 1 17054
2 65842 1 17054
2 65843 1 17057
2 65844 1 17057
2 65845 1 17057
2 65846 1 17069
2 65847 1 17069
2 65848 1 17077
2 65849 1 17077
2 65850 1 17077
2 65851 1 17077
2 65852 1 17077
2 65853 1 17077
2 65854 1 17077
2 65855 1 17077
2 65856 1 17077
2 65857 1 17077
2 65858 1 17077
2 65859 1 17077
2 65860 1 17077
2 65861 1 17077
2 65862 1 17077
2 65863 1 17078
2 65864 1 17078
2 65865 1 17078
2 65866 1 17078
2 65867 1 17080
2 65868 1 17080
2 65869 1 17080
2 65870 1 17080
2 65871 1 17081
2 65872 1 17081
2 65873 1 17081
2 65874 1 17088
2 65875 1 17088
2 65876 1 17088
2 65877 1 17088
2 65878 1 17089
2 65879 1 17089
2 65880 1 17089
2 65881 1 17089
2 65882 1 17089
2 65883 1 17090
2 65884 1 17090
2 65885 1 17090
2 65886 1 17098
2 65887 1 17098
2 65888 1 17098
2 65889 1 17099
2 65890 1 17099
2 65891 1 17099
2 65892 1 17099
2 65893 1 17099
2 65894 1 17099
2 65895 1 17099
2 65896 1 17099
2 65897 1 17099
2 65898 1 17099
2 65899 1 17099
2 65900 1 17099
2 65901 1 17099
2 65902 1 17099
2 65903 1 17099
2 65904 1 17099
2 65905 1 17099
2 65906 1 17099
2 65907 1 17099
2 65908 1 17099
2 65909 1 17099
2 65910 1 17099
2 65911 1 17099
2 65912 1 17099
2 65913 1 17099
2 65914 1 17099
2 65915 1 17099
2 65916 1 17099
2 65917 1 17099
2 65918 1 17099
2 65919 1 17099
2 65920 1 17099
2 65921 1 17099
2 65922 1 17099
2 65923 1 17099
2 65924 1 17099
2 65925 1 17099
2 65926 1 17099
2 65927 1 17099
2 65928 1 17099
2 65929 1 17099
2 65930 1 17099
2 65931 1 17099
2 65932 1 17099
2 65933 1 17099
2 65934 1 17099
2 65935 1 17099
2 65936 1 17099
2 65937 1 17099
2 65938 1 17099
2 65939 1 17099
2 65940 1 17099
2 65941 1 17099
2 65942 1 17099
2 65943 1 17099
2 65944 1 17099
2 65945 1 17099
2 65946 1 17099
2 65947 1 17099
2 65948 1 17099
2 65949 1 17099
2 65950 1 17099
2 65951 1 17099
2 65952 1 17099
2 65953 1 17099
2 65954 1 17099
2 65955 1 17099
2 65956 1 17099
2 65957 1 17099
2 65958 1 17099
2 65959 1 17099
2 65960 1 17099
2 65961 1 17099
2 65962 1 17099
2 65963 1 17099
2 65964 1 17099
2 65965 1 17099
2 65966 1 17099
2 65967 1 17099
2 65968 1 17099
2 65969 1 17099
2 65970 1 17099
2 65971 1 17099
2 65972 1 17099
2 65973 1 17099
2 65974 1 17099
2 65975 1 17099
2 65976 1 17099
2 65977 1 17099
2 65978 1 17099
2 65979 1 17099
2 65980 1 17099
2 65981 1 17099
2 65982 1 17099
2 65983 1 17099
2 65984 1 17099
2 65985 1 17099
2 65986 1 17102
2 65987 1 17102
2 65988 1 17102
2 65989 1 17102
2 65990 1 17102
2 65991 1 17102
2 65992 1 17102
2 65993 1 17102
2 65994 1 17102
2 65995 1 17102
2 65996 1 17102
2 65997 1 17102
2 65998 1 17102
2 65999 1 17102
2 66000 1 17102
2 66001 1 17102
2 66002 1 17102
2 66003 1 17102
2 66004 1 17102
2 66005 1 17102
2 66006 1 17102
2 66007 1 17102
2 66008 1 17102
2 66009 1 17102
2 66010 1 17102
2 66011 1 17102
2 66012 1 17102
2 66013 1 17102
2 66014 1 17102
2 66015 1 17102
2 66016 1 17102
2 66017 1 17102
2 66018 1 17102
2 66019 1 17102
2 66020 1 17102
2 66021 1 17102
2 66022 1 17102
2 66023 1 17102
2 66024 1 17102
2 66025 1 17102
2 66026 1 17102
2 66027 1 17102
2 66028 1 17102
2 66029 1 17102
2 66030 1 17102
2 66031 1 17102
2 66032 1 17111
2 66033 1 17111
2 66034 1 17111
2 66035 1 17111
2 66036 1 17111
2 66037 1 17111
2 66038 1 17111
2 66039 1 17111
2 66040 1 17111
2 66041 1 17111
2 66042 1 17111
2 66043 1 17111
2 66044 1 17112
2 66045 1 17112
2 66046 1 17112
2 66047 1 17113
2 66048 1 17113
2 66049 1 17113
2 66050 1 17113
2 66051 1 17113
2 66052 1 17113
2 66053 1 17113
2 66054 1 17113
2 66055 1 17113
2 66056 1 17113
2 66057 1 17113
2 66058 1 17113
2 66059 1 17113
2 66060 1 17113
2 66061 1 17113
2 66062 1 17113
2 66063 1 17113
2 66064 1 17113
2 66065 1 17113
2 66066 1 17113
2 66067 1 17113
2 66068 1 17113
2 66069 1 17113
2 66070 1 17113
2 66071 1 17113
2 66072 1 17113
2 66073 1 17113
2 66074 1 17113
2 66075 1 17122
2 66076 1 17122
2 66077 1 17125
2 66078 1 17125
2 66079 1 17125
2 66080 1 17126
2 66081 1 17126
2 66082 1 17142
2 66083 1 17142
2 66084 1 17142
2 66085 1 17142
2 66086 1 17142
2 66087 1 17143
2 66088 1 17143
2 66089 1 17145
2 66090 1 17145
2 66091 1 17145
2 66092 1 17145
2 66093 1 17145
2 66094 1 17145
2 66095 1 17145
2 66096 1 17148
2 66097 1 17148
2 66098 1 17164
2 66099 1 17164
2 66100 1 17164
2 66101 1 17164
2 66102 1 17167
2 66103 1 17167
2 66104 1 17167
2 66105 1 17167
2 66106 1 17175
2 66107 1 17175
2 66108 1 17175
2 66109 1 17175
2 66110 1 17175
2 66111 1 17176
2 66112 1 17176
2 66113 1 17179
2 66114 1 17179
2 66115 1 17188
2 66116 1 17188
2 66117 1 17190
2 66118 1 17190
2 66119 1 17190
2 66120 1 17190
2 66121 1 17205
2 66122 1 17205
2 66123 1 17205
2 66124 1 17222
2 66125 1 17222
2 66126 1 17222
2 66127 1 17222
2 66128 1 17222
2 66129 1 17222
2 66130 1 17222
2 66131 1 17222
2 66132 1 17222
2 66133 1 17222
2 66134 1 17222
2 66135 1 17222
2 66136 1 17222
2 66137 1 17222
2 66138 1 17222
2 66139 1 17222
2 66140 1 17222
2 66141 1 17222
2 66142 1 17222
2 66143 1 17222
2 66144 1 17222
2 66145 1 17222
2 66146 1 17222
2 66147 1 17222
2 66148 1 17223
2 66149 1 17223
2 66150 1 17224
2 66151 1 17224
2 66152 1 17224
2 66153 1 17224
2 66154 1 17224
2 66155 1 17224
2 66156 1 17224
2 66157 1 17224
2 66158 1 17224
2 66159 1 17224
2 66160 1 17224
2 66161 1 17224
2 66162 1 17224
2 66163 1 17225
2 66164 1 17225
2 66165 1 17225
2 66166 1 17225
2 66167 1 17225
2 66168 1 17225
2 66169 1 17225
2 66170 1 17225
2 66171 1 17225
2 66172 1 17225
2 66173 1 17225
2 66174 1 17225
2 66175 1 17225
2 66176 1 17226
2 66177 1 17226
2 66178 1 17226
2 66179 1 17226
2 66180 1 17228
2 66181 1 17228
2 66182 1 17228
2 66183 1 17228
2 66184 1 17228
2 66185 1 17229
2 66186 1 17229
2 66187 1 17229
2 66188 1 17229
2 66189 1 17229
2 66190 1 17229
2 66191 1 17229
2 66192 1 17229
2 66193 1 17229
2 66194 1 17229
2 66195 1 17229
2 66196 1 17229
2 66197 1 17229
2 66198 1 17229
2 66199 1 17233
2 66200 1 17233
2 66201 1 17233
2 66202 1 17233
2 66203 1 17233
2 66204 1 17233
2 66205 1 17233
2 66206 1 17233
2 66207 1 17233
2 66208 1 17233
2 66209 1 17233
2 66210 1 17233
2 66211 1 17233
2 66212 1 17236
2 66213 1 17236
2 66214 1 17236
2 66215 1 17236
2 66216 1 17236
2 66217 1 17236
2 66218 1 17237
2 66219 1 17237
2 66220 1 17237
2 66221 1 17237
2 66222 1 17237
2 66223 1 17237
2 66224 1 17238
2 66225 1 17238
2 66226 1 17238
2 66227 1 17241
2 66228 1 17241
2 66229 1 17241
2 66230 1 17241
2 66231 1 17241
2 66232 1 17241
2 66233 1 17241
2 66234 1 17241
2 66235 1 17244
2 66236 1 17244
2 66237 1 17244
2 66238 1 17244
2 66239 1 17244
2 66240 1 17244
2 66241 1 17244
2 66242 1 17245
2 66243 1 17245
2 66244 1 17245
2 66245 1 17245
2 66246 1 17245
2 66247 1 17247
2 66248 1 17247
2 66249 1 17247
2 66250 1 17247
2 66251 1 17247
2 66252 1 17247
2 66253 1 17247
2 66254 1 17248
2 66255 1 17248
2 66256 1 17251
2 66257 1 17251
2 66258 1 17251
2 66259 1 17251
2 66260 1 17251
2 66261 1 17251
2 66262 1 17251
2 66263 1 17251
2 66264 1 17251
2 66265 1 17251
2 66266 1 17251
2 66267 1 17251
2 66268 1 17251
2 66269 1 17251
2 66270 1 17251
2 66271 1 17251
2 66272 1 17251
2 66273 1 17251
2 66274 1 17251
2 66275 1 17251
2 66276 1 17251
2 66277 1 17251
2 66278 1 17251
2 66279 1 17251
2 66280 1 17251
2 66281 1 17251
2 66282 1 17251
2 66283 1 17251
2 66284 1 17251
2 66285 1 17251
2 66286 1 17251
2 66287 1 17252
2 66288 1 17252
2 66289 1 17258
2 66290 1 17258
2 66291 1 17258
2 66292 1 17258
2 66293 1 17259
2 66294 1 17259
2 66295 1 17259
2 66296 1 17259
2 66297 1 17260
2 66298 1 17260
2 66299 1 17263
2 66300 1 17263
2 66301 1 17263
2 66302 1 17263
2 66303 1 17263
2 66304 1 17263
2 66305 1 17263
2 66306 1 17263
2 66307 1 17263
2 66308 1 17263
2 66309 1 17263
2 66310 1 17263
2 66311 1 17268
2 66312 1 17268
2 66313 1 17271
2 66314 1 17271
2 66315 1 17271
2 66316 1 17271
2 66317 1 17271
2 66318 1 17271
2 66319 1 17271
2 66320 1 17275
2 66321 1 17275
2 66322 1 17275
2 66323 1 17275
2 66324 1 17287
2 66325 1 17287
2 66326 1 17287
2 66327 1 17288
2 66328 1 17288
2 66329 1 17292
2 66330 1 17292
2 66331 1 17304
2 66332 1 17304
2 66333 1 17304
2 66334 1 17304
2 66335 1 17304
2 66336 1 17304
2 66337 1 17304
2 66338 1 17305
2 66339 1 17305
2 66340 1 17305
2 66341 1 17305
2 66342 1 17305
2 66343 1 17305
2 66344 1 17305
2 66345 1 17305
2 66346 1 17305
2 66347 1 17305
2 66348 1 17307
2 66349 1 17307
2 66350 1 17307
2 66351 1 17310
2 66352 1 17310
2 66353 1 17311
2 66354 1 17311
2 66355 1 17311
2 66356 1 17311
2 66357 1 17311
2 66358 1 17311
2 66359 1 17311
2 66360 1 17311
2 66361 1 17311
2 66362 1 17311
2 66363 1 17311
2 66364 1 17311
2 66365 1 17319
2 66366 1 17319
2 66367 1 17320
2 66368 1 17320
2 66369 1 17320
2 66370 1 17320
2 66371 1 17320
2 66372 1 17323
2 66373 1 17323
2 66374 1 17323
2 66375 1 17323
2 66376 1 17323
2 66377 1 17323
2 66378 1 17323
2 66379 1 17323
2 66380 1 17323
2 66381 1 17323
2 66382 1 17323
2 66383 1 17323
2 66384 1 17323
2 66385 1 17323
2 66386 1 17323
2 66387 1 17323
2 66388 1 17323
2 66389 1 17323
2 66390 1 17323
2 66391 1 17331
2 66392 1 17331
2 66393 1 17331
2 66394 1 17331
2 66395 1 17331
2 66396 1 17332
2 66397 1 17332
2 66398 1 17332
2 66399 1 17339
2 66400 1 17339
2 66401 1 17340
2 66402 1 17340
2 66403 1 17340
2 66404 1 17348
2 66405 1 17348
2 66406 1 17348
2 66407 1 17348
2 66408 1 17349
2 66409 1 17349
2 66410 1 17349
2 66411 1 17349
2 66412 1 17349
2 66413 1 17349
2 66414 1 17352
2 66415 1 17352
2 66416 1 17352
2 66417 1 17380
2 66418 1 17380
2 66419 1 17380
2 66420 1 17380
2 66421 1 17381
2 66422 1 17381
2 66423 1 17381
2 66424 1 17391
2 66425 1 17391
2 66426 1 17391
2 66427 1 17391
2 66428 1 17414
2 66429 1 17414
2 66430 1 17414
2 66431 1 17414
2 66432 1 17424
2 66433 1 17424
2 66434 1 17424
2 66435 1 17429
2 66436 1 17429
2 66437 1 17430
2 66438 1 17430
2 66439 1 17430
2 66440 1 17430
2 66441 1 17430
2 66442 1 17431
2 66443 1 17431
2 66444 1 17431
2 66445 1 17431
2 66446 1 17455
2 66447 1 17455
2 66448 1 17455
2 66449 1 17455
2 66450 1 17455
2 66451 1 17458
2 66452 1 17458
2 66453 1 17458
2 66454 1 17458
2 66455 1 17468
2 66456 1 17468
2 66457 1 17477
2 66458 1 17477
2 66459 1 17483
2 66460 1 17483
2 66461 1 17483
2 66462 1 17483
2 66463 1 17483
2 66464 1 17483
2 66465 1 17483
2 66466 1 17485
2 66467 1 17485
2 66468 1 17489
2 66469 1 17489
2 66470 1 17489
2 66471 1 17489
2 66472 1 17489
2 66473 1 17489
2 66474 1 17489
2 66475 1 17489
2 66476 1 17489
2 66477 1 17504
2 66478 1 17504
2 66479 1 17504
2 66480 1 17504
2 66481 1 17504
2 66482 1 17504
2 66483 1 17504
2 66484 1 17504
2 66485 1 17504
2 66486 1 17504
2 66487 1 17504
2 66488 1 17504
2 66489 1 17504
2 66490 1 17504
2 66491 1 17504
2 66492 1 17505
2 66493 1 17505
2 66494 1 17505
2 66495 1 17505
2 66496 1 17513
2 66497 1 17513
2 66498 1 17513
2 66499 1 17513
2 66500 1 17513
2 66501 1 17513
2 66502 1 17513
2 66503 1 17513
2 66504 1 17513
2 66505 1 17513
2 66506 1 17513
2 66507 1 17513
2 66508 1 17513
2 66509 1 17513
2 66510 1 17513
2 66511 1 17513
2 66512 1 17513
2 66513 1 17513
2 66514 1 17517
2 66515 1 17517
2 66516 1 17517
2 66517 1 17517
2 66518 1 17517
2 66519 1 17517
2 66520 1 17517
2 66521 1 17517
2 66522 1 17517
2 66523 1 17517
2 66524 1 17517
2 66525 1 17517
2 66526 1 17518
2 66527 1 17518
2 66528 1 17518
2 66529 1 17525
2 66530 1 17525
2 66531 1 17525
2 66532 1 17525
2 66533 1 17525
2 66534 1 17532
2 66535 1 17532
2 66536 1 17532
2 66537 1 17533
2 66538 1 17533
2 66539 1 17533
2 66540 1 17533
2 66541 1 17533
2 66542 1 17533
2 66543 1 17533
2 66544 1 17533
2 66545 1 17533
2 66546 1 17533
2 66547 1 17533
2 66548 1 17533
2 66549 1 17533
2 66550 1 17533
2 66551 1 17533
2 66552 1 17533
2 66553 1 17533
2 66554 1 17533
2 66555 1 17533
2 66556 1 17533
2 66557 1 17533
2 66558 1 17533
2 66559 1 17533
2 66560 1 17533
2 66561 1 17533
2 66562 1 17533
2 66563 1 17533
2 66564 1 17533
2 66565 1 17533
2 66566 1 17534
2 66567 1 17534
2 66568 1 17535
2 66569 1 17535
2 66570 1 17535
2 66571 1 17535
2 66572 1 17535
2 66573 1 17535
2 66574 1 17535
2 66575 1 17535
2 66576 1 17535
2 66577 1 17535
2 66578 1 17535
2 66579 1 17536
2 66580 1 17536
2 66581 1 17538
2 66582 1 17538
2 66583 1 17539
2 66584 1 17539
2 66585 1 17539
2 66586 1 17539
2 66587 1 17546
2 66588 1 17546
2 66589 1 17546
2 66590 1 17546
2 66591 1 17546
2 66592 1 17546
2 66593 1 17546
2 66594 1 17546
2 66595 1 17569
2 66596 1 17569
2 66597 1 17570
2 66598 1 17570
2 66599 1 17570
2 66600 1 17571
2 66601 1 17571
2 66602 1 17571
2 66603 1 17579
2 66604 1 17579
2 66605 1 17579
2 66606 1 17579
2 66607 1 17579
2 66608 1 17579
2 66609 1 17581
2 66610 1 17581
2 66611 1 17581
2 66612 1 17581
2 66613 1 17582
2 66614 1 17582
2 66615 1 17582
2 66616 1 17587
2 66617 1 17587
2 66618 1 17589
2 66619 1 17589
2 66620 1 17589
2 66621 1 17590
2 66622 1 17590
2 66623 1 17598
2 66624 1 17598
2 66625 1 17604
2 66626 1 17604
2 66627 1 17608
2 66628 1 17608
2 66629 1 17608
2 66630 1 17608
2 66631 1 17608
2 66632 1 17608
2 66633 1 17608
2 66634 1 17608
2 66635 1 17608
2 66636 1 17608
2 66637 1 17608
2 66638 1 17611
2 66639 1 17611
2 66640 1 17611
2 66641 1 17611
2 66642 1 17612
2 66643 1 17612
2 66644 1 17612
2 66645 1 17613
2 66646 1 17613
2 66647 1 17613
2 66648 1 17613
2 66649 1 17613
2 66650 1 17613
2 66651 1 17613
2 66652 1 17613
2 66653 1 17613
2 66654 1 17614
2 66655 1 17614
2 66656 1 17624
2 66657 1 17624
2 66658 1 17642
2 66659 1 17642
2 66660 1 17642
2 66661 1 17642
2 66662 1 17642
2 66663 1 17654
2 66664 1 17654
2 66665 1 17654
2 66666 1 17682
2 66667 1 17682
2 66668 1 17692
2 66669 1 17692
2 66670 1 17700
2 66671 1 17700
2 66672 1 17700
2 66673 1 17705
2 66674 1 17705
2 66675 1 17705
2 66676 1 17718
2 66677 1 17718
2 66678 1 17718
2 66679 1 17718
2 66680 1 17718
2 66681 1 17718
2 66682 1 17729
2 66683 1 17729
2 66684 1 17729
2 66685 1 17729
2 66686 1 17729
2 66687 1 17741
2 66688 1 17741
2 66689 1 17741
2 66690 1 17741
2 66691 1 17742
2 66692 1 17742
2 66693 1 17750
2 66694 1 17750
2 66695 1 17750
2 66696 1 17752
2 66697 1 17752
2 66698 1 17752
2 66699 1 17752
2 66700 1 17752
2 66701 1 17752
2 66702 1 17752
2 66703 1 17755
2 66704 1 17755
2 66705 1 17767
2 66706 1 17767
2 66707 1 17767
2 66708 1 17768
2 66709 1 17768
2 66710 1 17769
2 66711 1 17769
2 66712 1 17769
2 66713 1 17769
2 66714 1 17780
2 66715 1 17780
2 66716 1 17780
2 66717 1 17780
2 66718 1 17781
2 66719 1 17781
2 66720 1 17782
2 66721 1 17782
2 66722 1 17782
2 66723 1 17782
2 66724 1 17782
2 66725 1 17782
2 66726 1 17782
2 66727 1 17796
2 66728 1 17796
2 66729 1 17796
2 66730 1 17796
2 66731 1 17796
2 66732 1 17796
2 66733 1 17796
2 66734 1 17796
2 66735 1 17796
2 66736 1 17796
2 66737 1 17797
2 66738 1 17797
2 66739 1 17804
2 66740 1 17804
2 66741 1 17804
2 66742 1 17805
2 66743 1 17805
2 66744 1 17806
2 66745 1 17806
2 66746 1 17807
2 66747 1 17807
2 66748 1 17807
2 66749 1 17807
2 66750 1 17813
2 66751 1 17813
2 66752 1 17813
2 66753 1 17813
2 66754 1 17813
2 66755 1 17814
2 66756 1 17814
2 66757 1 17817
2 66758 1 17817
2 66759 1 17817
2 66760 1 17818
2 66761 1 17818
2 66762 1 17818
2 66763 1 17830
2 66764 1 17830
2 66765 1 17831
2 66766 1 17831
2 66767 1 17832
2 66768 1 17832
2 66769 1 17832
2 66770 1 17832
2 66771 1 17833
2 66772 1 17833
2 66773 1 17835
2 66774 1 17835
2 66775 1 17835
2 66776 1 17835
2 66777 1 17840
2 66778 1 17840
2 66779 1 17845
2 66780 1 17845
2 66781 1 17846
2 66782 1 17846
2 66783 1 17846
2 66784 1 17846
2 66785 1 17850
2 66786 1 17850
2 66787 1 17850
2 66788 1 17850
2 66789 1 17850
2 66790 1 17850
2 66791 1 17850
2 66792 1 17850
2 66793 1 17850
2 66794 1 17850
2 66795 1 17850
2 66796 1 17867
2 66797 1 17867
2 66798 1 17872
2 66799 1 17872
2 66800 1 17903
2 66801 1 17903
2 66802 1 17903
2 66803 1 17903
2 66804 1 17904
2 66805 1 17904
2 66806 1 17904
2 66807 1 17904
2 66808 1 17907
2 66809 1 17907
2 66810 1 17914
2 66811 1 17914
2 66812 1 17916
2 66813 1 17916
2 66814 1 17916
2 66815 1 17916
2 66816 1 17916
2 66817 1 17917
2 66818 1 17917
2 66819 1 17917
2 66820 1 17917
2 66821 1 17918
2 66822 1 17918
2 66823 1 17918
2 66824 1 17918
2 66825 1 17918
2 66826 1 17918
2 66827 1 17918
2 66828 1 17918
2 66829 1 17918
2 66830 1 17918
2 66831 1 17918
2 66832 1 17918
2 66833 1 17921
2 66834 1 17921
2 66835 1 17921
2 66836 1 17922
2 66837 1 17922
2 66838 1 17922
2 66839 1 17922
2 66840 1 17922
2 66841 1 17922
2 66842 1 17922
2 66843 1 17922
2 66844 1 17922
2 66845 1 17924
2 66846 1 17924
2 66847 1 17929
2 66848 1 17929
2 66849 1 17932
2 66850 1 17932
2 66851 1 17932
2 66852 1 17938
2 66853 1 17938
2 66854 1 17938
2 66855 1 17938
2 66856 1 17938
2 66857 1 17939
2 66858 1 17939
2 66859 1 17939
2 66860 1 17941
2 66861 1 17941
2 66862 1 17941
2 66863 1 17944
2 66864 1 17944
2 66865 1 17946
2 66866 1 17946
2 66867 1 17946
2 66868 1 17946
2 66869 1 17946
2 66870 1 17946
2 66871 1 17947
2 66872 1 17947
2 66873 1 17947
2 66874 1 17947
2 66875 1 17948
2 66876 1 17948
2 66877 1 17949
2 66878 1 17949
2 66879 1 17949
2 66880 1 17949
2 66881 1 17949
2 66882 1 17949
2 66883 1 17949
2 66884 1 17952
2 66885 1 17952
2 66886 1 17952
2 66887 1 17952
2 66888 1 17952
2 66889 1 17952
2 66890 1 17952
2 66891 1 17952
2 66892 1 17952
2 66893 1 17952
2 66894 1 17955
2 66895 1 17955
2 66896 1 17956
2 66897 1 17956
2 66898 1 17956
2 66899 1 17956
2 66900 1 17956
2 66901 1 17960
2 66902 1 17960
2 66903 1 17977
2 66904 1 17977
2 66905 1 17977
2 66906 1 17977
2 66907 1 17979
2 66908 1 17979
2 66909 1 17979
2 66910 1 17979
2 66911 1 17979
2 66912 1 17979
2 66913 1 17980
2 66914 1 17980
2 66915 1 17980
2 66916 1 17980
2 66917 1 17980
2 66918 1 17980
2 66919 1 17980
2 66920 1 17980
2 66921 1 17980
2 66922 1 17980
2 66923 1 17980
2 66924 1 17980
2 66925 1 17983
2 66926 1 17983
2 66927 1 18001
2 66928 1 18001
2 66929 1 18007
2 66930 1 18007
2 66931 1 18007
2 66932 1 18008
2 66933 1 18008
2 66934 1 18022
2 66935 1 18022
2 66936 1 18030
2 66937 1 18030
2 66938 1 18030
2 66939 1 18030
2 66940 1 18030
2 66941 1 18030
2 66942 1 18031
2 66943 1 18031
2 66944 1 18031
2 66945 1 18033
2 66946 1 18033
2 66947 1 18033
2 66948 1 18033
2 66949 1 18033
2 66950 1 18033
2 66951 1 18033
2 66952 1 18034
2 66953 1 18034
2 66954 1 18034
2 66955 1 18034
2 66956 1 18035
2 66957 1 18035
2 66958 1 18035
2 66959 1 18035
2 66960 1 18047
2 66961 1 18047
2 66962 1 18051
2 66963 1 18051
2 66964 1 18051
2 66965 1 18051
2 66966 1 18051
2 66967 1 18054
2 66968 1 18054
2 66969 1 18059
2 66970 1 18059
2 66971 1 18059
2 66972 1 18059
2 66973 1 18059
2 66974 1 18059
2 66975 1 18060
2 66976 1 18060
2 66977 1 18061
2 66978 1 18061
2 66979 1 18061
2 66980 1 18062
2 66981 1 18062
2 66982 1 18062
2 66983 1 18064
2 66984 1 18064
2 66985 1 18064
2 66986 1 18067
2 66987 1 18067
2 66988 1 18067
2 66989 1 18067
2 66990 1 18067
2 66991 1 18068
2 66992 1 18068
2 66993 1 18076
2 66994 1 18076
2 66995 1 18086
2 66996 1 18086
2 66997 1 18086
2 66998 1 18121
2 66999 1 18121
2 67000 1 18121
2 67001 1 18131
2 67002 1 18131
2 67003 1 18132
2 67004 1 18132
2 67005 1 18132
2 67006 1 18148
2 67007 1 18148
2 67008 1 18153
2 67009 1 18153
2 67010 1 18153
2 67011 1 18153
2 67012 1 18153
2 67013 1 18153
2 67014 1 18153
2 67015 1 18153
2 67016 1 18153
2 67017 1 18153
2 67018 1 18153
2 67019 1 18153
2 67020 1 18153
2 67021 1 18153
2 67022 1 18153
2 67023 1 18153
2 67024 1 18153
2 67025 1 18153
2 67026 1 18153
2 67027 1 18153
2 67028 1 18153
2 67029 1 18153
2 67030 1 18153
2 67031 1 18153
2 67032 1 18153
2 67033 1 18153
2 67034 1 18153
2 67035 1 18153
2 67036 1 18153
2 67037 1 18153
2 67038 1 18158
2 67039 1 18158
2 67040 1 18158
2 67041 1 18158
2 67042 1 18162
2 67043 1 18162
2 67044 1 18162
2 67045 1 18162
2 67046 1 18162
2 67047 1 18162
2 67048 1 18162
2 67049 1 18162
2 67050 1 18162
2 67051 1 18162
2 67052 1 18162
2 67053 1 18162
2 67054 1 18162
2 67055 1 18162
2 67056 1 18171
2 67057 1 18171
2 67058 1 18171
2 67059 1 18176
2 67060 1 18176
2 67061 1 18198
2 67062 1 18198
2 67063 1 18199
2 67064 1 18199
2 67065 1 18204
2 67066 1 18204
2 67067 1 18204
2 67068 1 18204
2 67069 1 18207
2 67070 1 18207
2 67071 1 18207
2 67072 1 18207
2 67073 1 18207
2 67074 1 18207
2 67075 1 18207
2 67076 1 18209
2 67077 1 18209
2 67078 1 18223
2 67079 1 18223
2 67080 1 18223
2 67081 1 18223
2 67082 1 18223
2 67083 1 18226
2 67084 1 18226
2 67085 1 18226
2 67086 1 18226
2 67087 1 18227
2 67088 1 18227
2 67089 1 18227
2 67090 1 18227
2 67091 1 18227
2 67092 1 18227
2 67093 1 18227
2 67094 1 18227
2 67095 1 18227
2 67096 1 18227
2 67097 1 18227
2 67098 1 18227
2 67099 1 18234
2 67100 1 18234
2 67101 1 18234
2 67102 1 18244
2 67103 1 18244
2 67104 1 18252
2 67105 1 18252
2 67106 1 18262
2 67107 1 18262
2 67108 1 18262
2 67109 1 18272
2 67110 1 18272
2 67111 1 18272
2 67112 1 18283
2 67113 1 18283
2 67114 1 18283
2 67115 1 18284
2 67116 1 18284
2 67117 1 18284
2 67118 1 18284
2 67119 1 18284
2 67120 1 18284
2 67121 1 18284
2 67122 1 18284
2 67123 1 18284
2 67124 1 18284
2 67125 1 18284
2 67126 1 18285
2 67127 1 18285
2 67128 1 18285
2 67129 1 18294
2 67130 1 18294
2 67131 1 18294
2 67132 1 18294
2 67133 1 18294
2 67134 1 18294
2 67135 1 18294
2 67136 1 18302
2 67137 1 18302
2 67138 1 18302
2 67139 1 18317
2 67140 1 18317
2 67141 1 18325
2 67142 1 18325
2 67143 1 18325
2 67144 1 18325
2 67145 1 18326
2 67146 1 18326
2 67147 1 18343
2 67148 1 18343
2 67149 1 18343
2 67150 1 18344
2 67151 1 18344
2 67152 1 18345
2 67153 1 18345
2 67154 1 18365
2 67155 1 18365
2 67156 1 18365
2 67157 1 18365
2 67158 1 18365
2 67159 1 18365
2 67160 1 18373
2 67161 1 18373
2 67162 1 18373
2 67163 1 18373
2 67164 1 18373
2 67165 1 18373
2 67166 1 18373
2 67167 1 18373
2 67168 1 18373
2 67169 1 18373
2 67170 1 18373
2 67171 1 18373
2 67172 1 18373
2 67173 1 18373
2 67174 1 18379
2 67175 1 18379
2 67176 1 18379
2 67177 1 18391
2 67178 1 18391
2 67179 1 18391
2 67180 1 18391
2 67181 1 18392
2 67182 1 18392
2 67183 1 18392
2 67184 1 18392
2 67185 1 18392
2 67186 1 18392
2 67187 1 18392
2 67188 1 18392
2 67189 1 18392
2 67190 1 18408
2 67191 1 18408
2 67192 1 18408
2 67193 1 18408
2 67194 1 18408
2 67195 1 18411
2 67196 1 18411
2 67197 1 18411
2 67198 1 18411
2 67199 1 18419
2 67200 1 18419
2 67201 1 18426
2 67202 1 18426
2 67203 1 18426
2 67204 1 18433
2 67205 1 18433
2 67206 1 18433
2 67207 1 18434
2 67208 1 18434
2 67209 1 18434
2 67210 1 18434
2 67211 1 18440
2 67212 1 18440
2 67213 1 18440
2 67214 1 18441
2 67215 1 18441
2 67216 1 18442
2 67217 1 18442
2 67218 1 18443
2 67219 1 18443
2 67220 1 18443
2 67221 1 18443
2 67222 1 18443
2 67223 1 18443
2 67224 1 18443
2 67225 1 18443
2 67226 1 18443
2 67227 1 18446
2 67228 1 18446
2 67229 1 18447
2 67230 1 18447
2 67231 1 18468
2 67232 1 18468
2 67233 1 18468
2 67234 1 18468
2 67235 1 18469
2 67236 1 18469
2 67237 1 18476
2 67238 1 18476
2 67239 1 18477
2 67240 1 18477
2 67241 1 18477
2 67242 1 18477
2 67243 1 18477
2 67244 1 18490
2 67245 1 18490
2 67246 1 18490
2 67247 1 18490
2 67248 1 18492
2 67249 1 18492
2 67250 1 18492
2 67251 1 18519
2 67252 1 18519
2 67253 1 18519
2 67254 1 18519
2 67255 1 18520
2 67256 1 18520
2 67257 1 18527
2 67258 1 18527
2 67259 1 18527
2 67260 1 18529
2 67261 1 18529
2 67262 1 18538
2 67263 1 18538
2 67264 1 18538
2 67265 1 18539
2 67266 1 18539
2 67267 1 18539
2 67268 1 18539
2 67269 1 18548
2 67270 1 18548
2 67271 1 18548
2 67272 1 18562
2 67273 1 18562
2 67274 1 18571
2 67275 1 18571
2 67276 1 18571
2 67277 1 18591
2 67278 1 18591
2 67279 1 18650
2 67280 1 18650
2 67281 1 18650
2 67282 1 18650
2 67283 1 18650
2 67284 1 18650
2 67285 1 18650
2 67286 1 18650
2 67287 1 18650
2 67288 1 18652
2 67289 1 18652
2 67290 1 18652
2 67291 1 18652
2 67292 1 18653
2 67293 1 18653
2 67294 1 18655
2 67295 1 18655
2 67296 1 18655
2 67297 1 18655
2 67298 1 18655
2 67299 1 18655
2 67300 1 18655
2 67301 1 18655
2 67302 1 18660
2 67303 1 18660
2 67304 1 18664
2 67305 1 18664
2 67306 1 18664
2 67307 1 18676
2 67308 1 18676
2 67309 1 18676
2 67310 1 18677
2 67311 1 18677
2 67312 1 18687
2 67313 1 18687
2 67314 1 18695
2 67315 1 18695
2 67316 1 18695
2 67317 1 18695
2 67318 1 18695
2 67319 1 18695
2 67320 1 18698
2 67321 1 18698
2 67322 1 18699
2 67323 1 18699
2 67324 1 18699
2 67325 1 18699
2 67326 1 18699
2 67327 1 18704
2 67328 1 18704
2 67329 1 18714
2 67330 1 18714
2 67331 1 18715
2 67332 1 18715
2 67333 1 18720
2 67334 1 18720
2 67335 1 18721
2 67336 1 18721
2 67337 1 18729
2 67338 1 18729
2 67339 1 18729
2 67340 1 18732
2 67341 1 18732
2 67342 1 18736
2 67343 1 18736
2 67344 1 18736
2 67345 1 18736
2 67346 1 18736
2 67347 1 18736
2 67348 1 18736
2 67349 1 18736
2 67350 1 18736
2 67351 1 18736
2 67352 1 18736
2 67353 1 18736
2 67354 1 18736
2 67355 1 18737
2 67356 1 18737
2 67357 1 18747
2 67358 1 18747
2 67359 1 18747
2 67360 1 18747
2 67361 1 18747
2 67362 1 18747
2 67363 1 18748
2 67364 1 18748
2 67365 1 18748
2 67366 1 18749
2 67367 1 18749
2 67368 1 18749
2 67369 1 18749
2 67370 1 18749
2 67371 1 18749
2 67372 1 18750
2 67373 1 18750
2 67374 1 18756
2 67375 1 18756
2 67376 1 18756
2 67377 1 18756
2 67378 1 18756
2 67379 1 18756
2 67380 1 18764
2 67381 1 18764
2 67382 1 18764
2 67383 1 18764
2 67384 1 18770
2 67385 1 18770
2 67386 1 18770
2 67387 1 18770
2 67388 1 18770
2 67389 1 18770
2 67390 1 18770
2 67391 1 18770
2 67392 1 18770
2 67393 1 18772
2 67394 1 18772
2 67395 1 18781
2 67396 1 18781
2 67397 1 18784
2 67398 1 18784
2 67399 1 18784
2 67400 1 18797
2 67401 1 18797
2 67402 1 18797
2 67403 1 18797
2 67404 1 18797
2 67405 1 18797
2 67406 1 18797
2 67407 1 18803
2 67408 1 18803
2 67409 1 18803
2 67410 1 18803
2 67411 1 18803
2 67412 1 18803
2 67413 1 18804
2 67414 1 18804
2 67415 1 18806
2 67416 1 18806
2 67417 1 18806
2 67418 1 18806
2 67419 1 18806
2 67420 1 18806
2 67421 1 18806
2 67422 1 18807
2 67423 1 18807
2 67424 1 18808
2 67425 1 18808
2 67426 1 18811
2 67427 1 18811
2 67428 1 18811
2 67429 1 18812
2 67430 1 18812
2 67431 1 18821
2 67432 1 18821
2 67433 1 18822
2 67434 1 18822
2 67435 1 18822
2 67436 1 18822
2 67437 1 18824
2 67438 1 18824
2 67439 1 18827
2 67440 1 18827
2 67441 1 18828
2 67442 1 18828
2 67443 1 18828
2 67444 1 18832
2 67445 1 18832
2 67446 1 18832
2 67447 1 18833
2 67448 1 18833
2 67449 1 18833
2 67450 1 18833
2 67451 1 18833
2 67452 1 18833
2 67453 1 18834
2 67454 1 18834
2 67455 1 18836
2 67456 1 18836
2 67457 1 18836
2 67458 1 18840
2 67459 1 18840
2 67460 1 18841
2 67461 1 18841
2 67462 1 18841
2 67463 1 18842
2 67464 1 18842
2 67465 1 18842
2 67466 1 18842
2 67467 1 18842
2 67468 1 18853
2 67469 1 18853
2 67470 1 18855
2 67471 1 18855
2 67472 1 18855
2 67473 1 18855
2 67474 1 18855
2 67475 1 18859
2 67476 1 18859
2 67477 1 18859
2 67478 1 18859
2 67479 1 18859
2 67480 1 18860
2 67481 1 18860
2 67482 1 18860
2 67483 1 18860
2 67484 1 18860
2 67485 1 18862
2 67486 1 18862
2 67487 1 18866
2 67488 1 18866
2 67489 1 18875
2 67490 1 18875
2 67491 1 18914
2 67492 1 18914
2 67493 1 18914
2 67494 1 18914
2 67495 1 18914
2 67496 1 18914
2 67497 1 18914
2 67498 1 18915
2 67499 1 18915
2 67500 1 18916
2 67501 1 18916
2 67502 1 18935
2 67503 1 18935
2 67504 1 18935
2 67505 1 18936
2 67506 1 18936
2 67507 1 18936
2 67508 1 18936
2 67509 1 18937
2 67510 1 18937
2 67511 1 18945
2 67512 1 18945
2 67513 1 18945
2 67514 1 18966
2 67515 1 18966
2 67516 1 18978
2 67517 1 18978
2 67518 1 18978
2 67519 1 18987
2 67520 1 18987
2 67521 1 18988
2 67522 1 18988
2 67523 1 18988
2 67524 1 18988
2 67525 1 18988
2 67526 1 18989
2 67527 1 18989
2 67528 1 18998
2 67529 1 18998
2 67530 1 19008
2 67531 1 19008
2 67532 1 19008
2 67533 1 19008
2 67534 1 19010
2 67535 1 19010
2 67536 1 19010
2 67537 1 19010
2 67538 1 19010
2 67539 1 19012
2 67540 1 19012
2 67541 1 19012
2 67542 1 19012
2 67543 1 19012
2 67544 1 19013
2 67545 1 19013
2 67546 1 19013
2 67547 1 19013
2 67548 1 19015
2 67549 1 19015
2 67550 1 19015
2 67551 1 19015
2 67552 1 19015
2 67553 1 19015
2 67554 1 19015
2 67555 1 19015
2 67556 1 19015
2 67557 1 19015
2 67558 1 19016
2 67559 1 19016
2 67560 1 19016
2 67561 1 19016
2 67562 1 19016
2 67563 1 19016
2 67564 1 19016
2 67565 1 19016
2 67566 1 19016
2 67567 1 19017
2 67568 1 19017
2 67569 1 19017
2 67570 1 19028
2 67571 1 19028
2 67572 1 19032
2 67573 1 19032
2 67574 1 19032
2 67575 1 19032
2 67576 1 19032
2 67577 1 19039
2 67578 1 19039
2 67579 1 19040
2 67580 1 19040
2 67581 1 19040
2 67582 1 19054
2 67583 1 19054
2 67584 1 19055
2 67585 1 19055
2 67586 1 19055
2 67587 1 19055
2 67588 1 19056
2 67589 1 19056
2 67590 1 19056
2 67591 1 19057
2 67592 1 19057
2 67593 1 19057
2 67594 1 19057
2 67595 1 19057
2 67596 1 19057
2 67597 1 19057
2 67598 1 19057
2 67599 1 19057
2 67600 1 19060
2 67601 1 19060
2 67602 1 19060
2 67603 1 19060
2 67604 1 19060
2 67605 1 19060
2 67606 1 19060
2 67607 1 19060
2 67608 1 19060
2 67609 1 19060
2 67610 1 19060
2 67611 1 19070
2 67612 1 19070
2 67613 1 19071
2 67614 1 19071
2 67615 1 19071
2 67616 1 19071
2 67617 1 19086
2 67618 1 19086
2 67619 1 19086
2 67620 1 19086
2 67621 1 19086
2 67622 1 19087
2 67623 1 19087
2 67624 1 19089
2 67625 1 19089
2 67626 1 19102
2 67627 1 19102
2 67628 1 19108
2 67629 1 19108
2 67630 1 19124
2 67631 1 19124
2 67632 1 19124
2 67633 1 19142
2 67634 1 19142
2 67635 1 19144
2 67636 1 19144
2 67637 1 19144
2 67638 1 19145
2 67639 1 19145
2 67640 1 19150
2 67641 1 19150
2 67642 1 19153
2 67643 1 19153
2 67644 1 19161
2 67645 1 19161
2 67646 1 19162
2 67647 1 19162
2 67648 1 19170
2 67649 1 19170
2 67650 1 19170
2 67651 1 19170
2 67652 1 19181
2 67653 1 19181
2 67654 1 19191
2 67655 1 19191
2 67656 1 19210
2 67657 1 19210
2 67658 1 19219
2 67659 1 19219
2 67660 1 19227
2 67661 1 19227
2 67662 1 19235
2 67663 1 19235
2 67664 1 19235
2 67665 1 19243
2 67666 1 19243
2 67667 1 19245
2 67668 1 19245
2 67669 1 19245
2 67670 1 19253
2 67671 1 19253
2 67672 1 19253
2 67673 1 19266
2 67674 1 19266
2 67675 1 19276
2 67676 1 19276
2 67677 1 19276
2 67678 1 19276
2 67679 1 19278
2 67680 1 19278
2 67681 1 19278
2 67682 1 19278
2 67683 1 19279
2 67684 1 19279
2 67685 1 19279
2 67686 1 19283
2 67687 1 19283
2 67688 1 19284
2 67689 1 19284
2 67690 1 19308
2 67691 1 19308
2 67692 1 19313
2 67693 1 19313
2 67694 1 19313
2 67695 1 19313
2 67696 1 19313
2 67697 1 19313
2 67698 1 19313
2 67699 1 19313
2 67700 1 19313
2 67701 1 19314
2 67702 1 19314
2 67703 1 19314
2 67704 1 19325
2 67705 1 19325
2 67706 1 19325
2 67707 1 19325
2 67708 1 19325
2 67709 1 19325
2 67710 1 19325
2 67711 1 19325
2 67712 1 19325
2 67713 1 19325
2 67714 1 19328
2 67715 1 19328
2 67716 1 19345
2 67717 1 19345
2 67718 1 19345
2 67719 1 19345
2 67720 1 19348
2 67721 1 19348
2 67722 1 19352
2 67723 1 19352
2 67724 1 19352
2 67725 1 19352
2 67726 1 19353
2 67727 1 19353
2 67728 1 19360
2 67729 1 19360
2 67730 1 19362
2 67731 1 19362
2 67732 1 19369
2 67733 1 19369
2 67734 1 19387
2 67735 1 19387
2 67736 1 19388
2 67737 1 19388
2 67738 1 19389
2 67739 1 19389
2 67740 1 19399
2 67741 1 19399
2 67742 1 19400
2 67743 1 19400
2 67744 1 19401
2 67745 1 19401
2 67746 1 19401
2 67747 1 19401
2 67748 1 19401
2 67749 1 19401
2 67750 1 19405
2 67751 1 19405
2 67752 1 19430
2 67753 1 19430
2 67754 1 19430
2 67755 1 19431
2 67756 1 19431
2 67757 1 19442
2 67758 1 19442
2 67759 1 19454
2 67760 1 19454
2 67761 1 19454
2 67762 1 19463
2 67763 1 19463
2 67764 1 19463
2 67765 1 19463
2 67766 1 19464
2 67767 1 19464
2 67768 1 19480
2 67769 1 19480
2 67770 1 19490
2 67771 1 19490
2 67772 1 19490
2 67773 1 19490
2 67774 1 19491
2 67775 1 19491
2 67776 1 19505
2 67777 1 19505
2 67778 1 19508
2 67779 1 19508
2 67780 1 19509
2 67781 1 19509
2 67782 1 19509
2 67783 1 19509
2 67784 1 19509
2 67785 1 19509
2 67786 1 19513
2 67787 1 19513
2 67788 1 19513
2 67789 1 19520
2 67790 1 19520
2 67791 1 19520
2 67792 1 19524
2 67793 1 19524
2 67794 1 19525
2 67795 1 19525
2 67796 1 19541
2 67797 1 19541
2 67798 1 19541
2 67799 1 19556
2 67800 1 19556
2 67801 1 19557
2 67802 1 19557
2 67803 1 19565
2 67804 1 19565
2 67805 1 19565
2 67806 1 19566
2 67807 1 19566
2 67808 1 19566
2 67809 1 19566
2 67810 1 19566
2 67811 1 19566
2 67812 1 19566
2 67813 1 19566
2 67814 1 19566
2 67815 1 19566
2 67816 1 19579
2 67817 1 19579
2 67818 1 19579
2 67819 1 19580
2 67820 1 19580
2 67821 1 19580
2 67822 1 19584
2 67823 1 19584
2 67824 1 19592
2 67825 1 19592
2 67826 1 19593
2 67827 1 19593
2 67828 1 19610
2 67829 1 19610
2 67830 1 19627
2 67831 1 19627
2 67832 1 19634
2 67833 1 19634
2 67834 1 19635
2 67835 1 19635
2 67836 1 19640
2 67837 1 19640
2 67838 1 19641
2 67839 1 19641
2 67840 1 19641
2 67841 1 19641
2 67842 1 19642
2 67843 1 19642
2 67844 1 19642
2 67845 1 19642
2 67846 1 19654
2 67847 1 19654
2 67848 1 19654
2 67849 1 19654
2 67850 1 19654
2 67851 1 19666
2 67852 1 19666
2 67853 1 19669
2 67854 1 19669
2 67855 1 19669
2 67856 1 19669
2 67857 1 19678
2 67858 1 19678
2 67859 1 19679
2 67860 1 19679
2 67861 1 19679
2 67862 1 19680
2 67863 1 19680
2 67864 1 19684
2 67865 1 19684
2 67866 1 19686
2 67867 1 19686
2 67868 1 19687
2 67869 1 19687
2 67870 1 19696
2 67871 1 19696
2 67872 1 19706
2 67873 1 19706
2 67874 1 19737
2 67875 1 19737
2 67876 1 19737
2 67877 1 19740
2 67878 1 19740
2 67879 1 19740
2 67880 1 19740
2 67881 1 19752
2 67882 1 19752
2 67883 1 19752
2 67884 1 19753
2 67885 1 19753
2 67886 1 19771
2 67887 1 19771
2 67888 1 19779
2 67889 1 19779
2 67890 1 19779
2 67891 1 19779
2 67892 1 19779
2 67893 1 19780
2 67894 1 19780
2 67895 1 19780
2 67896 1 19780
2 67897 1 19780
2 67898 1 19780
2 67899 1 19780
2 67900 1 19789
2 67901 1 19789
2 67902 1 19790
2 67903 1 19790
2 67904 1 19819
2 67905 1 19819
2 67906 1 19820
2 67907 1 19820
2 67908 1 19827
2 67909 1 19827
2 67910 1 19839
2 67911 1 19839
2 67912 1 19849
2 67913 1 19849
2 67914 1 19850
2 67915 1 19850
2 67916 1 19850
2 67917 1 19850
2 67918 1 19851
2 67919 1 19851
2 67920 1 19851
2 67921 1 19861
2 67922 1 19861
2 67923 1 19870
2 67924 1 19870
2 67925 1 19897
2 67926 1 19897
2 67927 1 19898
2 67928 1 19898
2 67929 1 19918
2 67930 1 19918
2 67931 1 19920
2 67932 1 19920
2 67933 1 19934
2 67934 1 19934
2 67935 1 19934
2 67936 1 19935
2 67937 1 19935
2 67938 1 19935
2 67939 1 19936
2 67940 1 19936
2 67941 1 19936
2 67942 1 19937
2 67943 1 19937
2 67944 1 19937
2 67945 1 19941
2 67946 1 19941
2 67947 1 19941
2 67948 1 19959
2 67949 1 19959
2 67950 1 19959
2 67951 1 19959
2 67952 1 19961
2 67953 1 19961
2 67954 1 19976
2 67955 1 19976
2 67956 1 19984
2 67957 1 19984
2 67958 1 19984
2 67959 1 19984
2 67960 1 19985
2 67961 1 19985
2 67962 1 19985
2 67963 1 19986
2 67964 1 19986
2 67965 1 19986
2 67966 1 19986
2 67967 1 19988
2 67968 1 19988
2 67969 1 19999
2 67970 1 19999
2 67971 1 19999
2 67972 1 19999
2 67973 1 19999
2 67974 1 20000
2 67975 1 20000
2 67976 1 20013
2 67977 1 20013
2 67978 1 20025
2 67979 1 20025
2 67980 1 20025
2 67981 1 20025
2 67982 1 20056
2 67983 1 20056
2 67984 1 20056
2 67985 1 20056
2 67986 1 20056
2 67987 1 20074
2 67988 1 20074
2 67989 1 20077
2 67990 1 20077
2 67991 1 20077
2 67992 1 20086
2 67993 1 20086
2 67994 1 20093
2 67995 1 20093
2 67996 1 20093
2 67997 1 20093
2 67998 1 20112
2 67999 1 20112
2 68000 1 20117
2 68001 1 20117
2 68002 1 20120
2 68003 1 20120
2 68004 1 20163
2 68005 1 20163
2 68006 1 20163
2 68007 1 20240
2 68008 1 20240
2 68009 1 20241
2 68010 1 20241
2 68011 1 20248
2 68012 1 20248
2 68013 1 20256
2 68014 1 20256
2 68015 1 20259
2 68016 1 20259
2 68017 1 20274
2 68018 1 20274
2 68019 1 20274
2 68020 1 20275
2 68021 1 20275
2 68022 1 20276
2 68023 1 20276
2 68024 1 20287
2 68025 1 20287
2 68026 1 20287
2 68027 1 20296
2 68028 1 20296
2 68029 1 20324
2 68030 1 20324
2 68031 1 20332
2 68032 1 20332
2 68033 1 20346
2 68034 1 20346
2 68035 1 20372
2 68036 1 20372
2 68037 1 20376
2 68038 1 20376
2 68039 1 20411
2 68040 1 20411
2 68041 1 20429
2 68042 1 20429
2 68043 1 20429
2 68044 1 20430
2 68045 1 20430
2 68046 1 20430
2 68047 1 20430
2 68048 1 20430
2 68049 1 20450
2 68050 1 20450
2 68051 1 20457
2 68052 1 20457
2 68053 1 20458
2 68054 1 20458
2 68055 1 20472
2 68056 1 20472
2 68057 1 20488
2 68058 1 20488
2 68059 1 20488
2 68060 1 20489
2 68061 1 20489
2 68062 1 20494
2 68063 1 20494
2 68064 1 20509
2 68065 1 20509
2 68066 1 20509
2 68067 1 20512
2 68068 1 20512
2 68069 1 20512
2 68070 1 20513
2 68071 1 20513
2 68072 1 20524
2 68073 1 20524
2 68074 1 20555
2 68075 1 20555
2 68076 1 20558
2 68077 1 20558
2 68078 1 20558
2 68079 1 20572
2 68080 1 20572
2 68081 1 20573
2 68082 1 20573
2 68083 1 20573
2 68084 1 20579
2 68085 1 20579
2 68086 1 20579
2 68087 1 20579
2 68088 1 20579
2 68089 1 20580
2 68090 1 20580
2 68091 1 20588
2 68092 1 20588
2 68093 1 20588
2 68094 1 20588
2 68095 1 20588
2 68096 1 20588
2 68097 1 20603
2 68098 1 20603
2 68099 1 20603
2 68100 1 20610
2 68101 1 20610
2 68102 1 20648
2 68103 1 20648
2 68104 1 20649
2 68105 1 20649
2 68106 1 20652
2 68107 1 20652
2 68108 1 20658
2 68109 1 20658
2 68110 1 20658
2 68111 1 20658
2 68112 1 20658
2 68113 1 20658
2 68114 1 20658
2 68115 1 20658
2 68116 1 20658
2 68117 1 20659
2 68118 1 20659
2 68119 1 20659
2 68120 1 20670
2 68121 1 20670
2 68122 1 20670
2 68123 1 20670
2 68124 1 20686
2 68125 1 20686
2 68126 1 20687
2 68127 1 20687
2 68128 1 20699
2 68129 1 20699
2 68130 1 20708
2 68131 1 20708
2 68132 1 20710
2 68133 1 20710
2 68134 1 20710
2 68135 1 20710
2 68136 1 20710
2 68137 1 20710
2 68138 1 20711
2 68139 1 20711
2 68140 1 20725
2 68141 1 20725
2 68142 1 20732
2 68143 1 20732
2 68144 1 20732
2 68145 1 20744
2 68146 1 20744
2 68147 1 20744
2 68148 1 20746
2 68149 1 20746
2 68150 1 20746
2 68151 1 20746
2 68152 1 20746
2 68153 1 20765
2 68154 1 20765
2 68155 1 20767
2 68156 1 20767
2 68157 1 20769
2 68158 1 20769
2 68159 1 20770
2 68160 1 20770
2 68161 1 20770
2 68162 1 20770
2 68163 1 20770
2 68164 1 20770
2 68165 1 20770
2 68166 1 20770
2 68167 1 20771
2 68168 1 20771
2 68169 1 20786
2 68170 1 20786
2 68171 1 20786
2 68172 1 20786
2 68173 1 20786
2 68174 1 20786
2 68175 1 20786
2 68176 1 20786
2 68177 1 20786
2 68178 1 20786
2 68179 1 20786
2 68180 1 20786
2 68181 1 20786
2 68182 1 20786
2 68183 1 20786
2 68184 1 20790
2 68185 1 20790
2 68186 1 20794
2 68187 1 20794
2 68188 1 20794
2 68189 1 20803
2 68190 1 20803
2 68191 1 20827
2 68192 1 20827
2 68193 1 20828
2 68194 1 20828
2 68195 1 20828
2 68196 1 20837
2 68197 1 20837
2 68198 1 20837
2 68199 1 20839
2 68200 1 20839
2 68201 1 20840
2 68202 1 20840
2 68203 1 20855
2 68204 1 20855
2 68205 1 20857
2 68206 1 20857
2 68207 1 20859
2 68208 1 20859
2 68209 1 20859
2 68210 1 20859
2 68211 1 20859
2 68212 1 20873
2 68213 1 20873
2 68214 1 20873
2 68215 1 20874
2 68216 1 20874
2 68217 1 20874
2 68218 1 20885
2 68219 1 20885
2 68220 1 20885
2 68221 1 20905
2 68222 1 20905
2 68223 1 20917
2 68224 1 20917
2 68225 1 20934
2 68226 1 20934
2 68227 1 20969
2 68228 1 20969
2 68229 1 20984
2 68230 1 20984
2 68231 1 20993
2 68232 1 20993
2 68233 1 21017
2 68234 1 21017
2 68235 1 21017
2 68236 1 21018
2 68237 1 21018
2 68238 1 21018
2 68239 1 21018
2 68240 1 21018
2 68241 1 21018
2 68242 1 21020
2 68243 1 21020
2 68244 1 21020
2 68245 1 21020
2 68246 1 21021
2 68247 1 21021
2 68248 1 21021
2 68249 1 21036
2 68250 1 21036
2 68251 1 21045
2 68252 1 21045
2 68253 1 21059
2 68254 1 21059
2 68255 1 21059
2 68256 1 21086
2 68257 1 21086
2 68258 1 21104
2 68259 1 21104
2 68260 1 21107
2 68261 1 21107
2 68262 1 21121
2 68263 1 21121
2 68264 1 21129
2 68265 1 21129
2 68266 1 21138
2 68267 1 21138
2 68268 1 21145
2 68269 1 21145
2 68270 1 21166
2 68271 1 21166
2 68272 1 21182
2 68273 1 21182
2 68274 1 21182
2 68275 1 21182
2 68276 1 21182
2 68277 1 21182
2 68278 1 21182
2 68279 1 21183
2 68280 1 21183
2 68281 1 21199
2 68282 1 21199
2 68283 1 21199
2 68284 1 21208
2 68285 1 21208
2 68286 1 21209
2 68287 1 21209
2 68288 1 21218
2 68289 1 21218
2 68290 1 21219
2 68291 1 21219
2 68292 1 21237
2 68293 1 21237
2 68294 1 21286
2 68295 1 21286
2 68296 1 21286
2 68297 1 21290
2 68298 1 21290
2 68299 1 21290
2 68300 1 21303
2 68301 1 21303
2 68302 1 21311
2 68303 1 21311
2 68304 1 21341
2 68305 1 21341
2 68306 1 21341
2 68307 1 21343
2 68308 1 21343
2 68309 1 21344
2 68310 1 21344
2 68311 1 21373
2 68312 1 21373
2 68313 1 21373
2 68314 1 21376
2 68315 1 21376
2 68316 1 21376
2 68317 1 21376
2 68318 1 21376
2 68319 1 21376
2 68320 1 21376
2 68321 1 21376
2 68322 1 21376
2 68323 1 21389
2 68324 1 21389
2 68325 1 21390
2 68326 1 21390
2 68327 1 21400
2 68328 1 21400
2 68329 1 21400
2 68330 1 21401
2 68331 1 21401
2 68332 1 21401
2 68333 1 21401
2 68334 1 21411
2 68335 1 21411
2 68336 1 21418
2 68337 1 21418
2 68338 1 21418
2 68339 1 21418
2 68340 1 21419
2 68341 1 21419
2 68342 1 21447
2 68343 1 21447
2 68344 1 21455
2 68345 1 21455
2 68346 1 21464
2 68347 1 21464
2 68348 1 21464
2 68349 1 21465
2 68350 1 21465
2 68351 1 21465
2 68352 1 21465
2 68353 1 21465
2 68354 1 21469
2 68355 1 21469
2 68356 1 21484
2 68357 1 21484
2 68358 1 21484
2 68359 1 21504
2 68360 1 21504
2 68361 1 21504
2 68362 1 21504
2 68363 1 21504
2 68364 1 21504
2 68365 1 21504
2 68366 1 21504
2 68367 1 21504
2 68368 1 21504
2 68369 1 21504
2 68370 1 21504
2 68371 1 21515
2 68372 1 21515
2 68373 1 21523
2 68374 1 21523
2 68375 1 21550
2 68376 1 21550
2 68377 1 21561
2 68378 1 21561
2 68379 1 21561
2 68380 1 21561
2 68381 1 21561
2 68382 1 21562
2 68383 1 21562
2 68384 1 21562
2 68385 1 21591
2 68386 1 21591
2 68387 1 21619
2 68388 1 21619
2 68389 1 21620
2 68390 1 21620
2 68391 1 21620
2 68392 1 21620
2 68393 1 21663
2 68394 1 21663
2 68395 1 21682
2 68396 1 21682
2 68397 1 21682
2 68398 1 21682
2 68399 1 21682
2 68400 1 21682
2 68401 1 21682
2 68402 1 21682
2 68403 1 21717
2 68404 1 21717
2 68405 1 21719
2 68406 1 21719
2 68407 1 21719
2 68408 1 21719
2 68409 1 21721
2 68410 1 21721
2 68411 1 21725
2 68412 1 21725
2 68413 1 21728
2 68414 1 21728
2 68415 1 21767
2 68416 1 21767
2 68417 1 21767
2 68418 1 21767
2 68419 1 21767
2 68420 1 21767
2 68421 1 21767
2 68422 1 21798
2 68423 1 21798
2 68424 1 21807
2 68425 1 21807
2 68426 1 21807
2 68427 1 21829
2 68428 1 21829
2 68429 1 21834
2 68430 1 21834
2 68431 1 21855
2 68432 1 21855
2 68433 1 21858
2 68434 1 21858
2 68435 1 21859
2 68436 1 21859
2 68437 1 21875
2 68438 1 21875
2 68439 1 21882
2 68440 1 21882
2 68441 1 21889
2 68442 1 21889
2 68443 1 21889
2 68444 1 21889
2 68445 1 21889
2 68446 1 21889
2 68447 1 21889
2 68448 1 21889
2 68449 1 21889
2 68450 1 21912
2 68451 1 21912
2 68452 1 21912
2 68453 1 21922
2 68454 1 21922
2 68455 1 21922
2 68456 1 21922
2 68457 1 21922
2 68458 1 21922
2 68459 1 21939
2 68460 1 21939
2 68461 1 21939
2 68462 1 21989
2 68463 1 21989
2 68464 1 22009
2 68465 1 22009
2 68466 1 22009
2 68467 1 22015
2 68468 1 22015
2 68469 1 22028
2 68470 1 22028
2 68471 1 22036
2 68472 1 22036
2 68473 1 22036
2 68474 1 22046
2 68475 1 22046
2 68476 1 22046
2 68477 1 22046
2 68478 1 22046
2 68479 1 22047
2 68480 1 22047
2 68481 1 22055
2 68482 1 22055
2 68483 1 22056
2 68484 1 22056
2 68485 1 22070
2 68486 1 22070
2 68487 1 22082
2 68488 1 22082
2 68489 1 22083
2 68490 1 22083
2 68491 1 22098
2 68492 1 22098
2 68493 1 22120
2 68494 1 22120
2 68495 1 22120
2 68496 1 22120
2 68497 1 22120
2 68498 1 22120
2 68499 1 22124
2 68500 1 22124
2 68501 1 22132
2 68502 1 22132
2 68503 1 22133
2 68504 1 22133
2 68505 1 22146
2 68506 1 22146
2 68507 1 22165
2 68508 1 22165
2 68509 1 22165
2 68510 1 22165
2 68511 1 22166
2 68512 1 22166
2 68513 1 22169
2 68514 1 22169
2 68515 1 22178
2 68516 1 22178
2 68517 1 22182
2 68518 1 22182
2 68519 1 22193
2 68520 1 22193
2 68521 1 22202
2 68522 1 22202
2 68523 1 22202
2 68524 1 22202
2 68525 1 22219
2 68526 1 22219
2 68527 1 22219
2 68528 1 22219
2 68529 1 22219
2 68530 1 22253
2 68531 1 22253
2 68532 1 22253
2 68533 1 22253
2 68534 1 22253
2 68535 1 22261
2 68536 1 22261
2 68537 1 22269
2 68538 1 22269
2 68539 1 22279
2 68540 1 22279
2 68541 1 22287
2 68542 1 22287
2 68543 1 22287
2 68544 1 22337
2 68545 1 22337
2 68546 1 22337
2 68547 1 22337
2 68548 1 22337
2 68549 1 22337
2 68550 1 22337
2 68551 1 22338
2 68552 1 22338
2 68553 1 22338
2 68554 1 22340
2 68555 1 22340
2 68556 1 22340
2 68557 1 22348
2 68558 1 22348
2 68559 1 22350
2 68560 1 22350
2 68561 1 22358
2 68562 1 22358
2 68563 1 22377
2 68564 1 22377
2 68565 1 22377
2 68566 1 22377
2 68567 1 22384
2 68568 1 22384
2 68569 1 22392
2 68570 1 22392
2 68571 1 22404
2 68572 1 22404
2 68573 1 22410
2 68574 1 22410
2 68575 1 22417
2 68576 1 22417
2 68577 1 22434
2 68578 1 22434
2 68579 1 22434
2 68580 1 22442
2 68581 1 22442
2 68582 1 22454
2 68583 1 22454
2 68584 1 22454
2 68585 1 22454
2 68586 1 22464
2 68587 1 22464
2 68588 1 22465
2 68589 1 22465
2 68590 1 22465
2 68591 1 22472
2 68592 1 22472
2 68593 1 22472
2 68594 1 22472
2 68595 1 22473
2 68596 1 22473
2 68597 1 22473
2 68598 1 22480
2 68599 1 22480
2 68600 1 22481
2 68601 1 22481
2 68602 1 22495
2 68603 1 22495
2 68604 1 22501
2 68605 1 22501
2 68606 1 22511
2 68607 1 22511
2 68608 1 22511
2 68609 1 22518
2 68610 1 22518
2 68611 1 22527
2 68612 1 22527
2 68613 1 22534
2 68614 1 22534
2 68615 1 22548
2 68616 1 22548
2 68617 1 22548
2 68618 1 22550
2 68619 1 22550
2 68620 1 22551
2 68621 1 22551
2 68622 1 22551
2 68623 1 22557
2 68624 1 22557
2 68625 1 22561
2 68626 1 22561
2 68627 1 22562
2 68628 1 22562
2 68629 1 22562
2 68630 1 22569
2 68631 1 22569
2 68632 1 22570
2 68633 1 22570
2 68634 1 22570
2 68635 1 22574
2 68636 1 22574
2 68637 1 22577
2 68638 1 22577
2 68639 1 22584
2 68640 1 22584
2 68641 1 22584
2 68642 1 22584
2 68643 1 22584
2 68644 1 22584
2 68645 1 22584
2 68646 1 22584
2 68647 1 22585
2 68648 1 22585
2 68649 1 22585
2 68650 1 22586
2 68651 1 22586
2 68652 1 22587
2 68653 1 22587
2 68654 1 22603
2 68655 1 22603
2 68656 1 22603
2 68657 1 22603
2 68658 1 22604
2 68659 1 22604
2 68660 1 22616
2 68661 1 22616
2 68662 1 22670
2 68663 1 22670
2 68664 1 22670
2 68665 1 22702
2 68666 1 22702
2 68667 1 22702
2 68668 1 22716
2 68669 1 22716
2 68670 1 22717
2 68671 1 22717
2 68672 1 22718
2 68673 1 22718
2 68674 1 22718
2 68675 1 22718
2 68676 1 22732
2 68677 1 22732
2 68678 1 22739
2 68679 1 22739
2 68680 1 22739
2 68681 1 22739
2 68682 1 22739
2 68683 1 22741
2 68684 1 22741
2 68685 1 22742
2 68686 1 22742
2 68687 1 22779
2 68688 1 22779
2 68689 1 22779
2 68690 1 22779
2 68691 1 22779
2 68692 1 22795
2 68693 1 22795
2 68694 1 22797
2 68695 1 22797
2 68696 1 22798
2 68697 1 22798
2 68698 1 22798
2 68699 1 22798
2 68700 1 22798
2 68701 1 22808
2 68702 1 22808
2 68703 1 22808
2 68704 1 22810
2 68705 1 22810
2 68706 1 22813
2 68707 1 22813
2 68708 1 22813
2 68709 1 22813
2 68710 1 22813
2 68711 1 22841
2 68712 1 22841
2 68713 1 22849
2 68714 1 22849
2 68715 1 22849
2 68716 1 22849
2 68717 1 22849
2 68718 1 22849
2 68719 1 22849
2 68720 1 22851
2 68721 1 22851
2 68722 1 22871
2 68723 1 22871
2 68724 1 22871
2 68725 1 22871
2 68726 1 22871
2 68727 1 22896
2 68728 1 22896
2 68729 1 22896
2 68730 1 22897
2 68731 1 22897
2 68732 1 22897
2 68733 1 22900
2 68734 1 22900
2 68735 1 22900
2 68736 1 22913
2 68737 1 22913
2 68738 1 22915
2 68739 1 22915
2 68740 1 22915
2 68741 1 22917
2 68742 1 22917
2 68743 1 22923
2 68744 1 22923
2 68745 1 22935
2 68746 1 22935
2 68747 1 22942
2 68748 1 22942
2 68749 1 22947
2 68750 1 22947
2 68751 1 22954
2 68752 1 22954
2 68753 1 22954
2 68754 1 22958
2 68755 1 22958
2 68756 1 22976
2 68757 1 22976
2 68758 1 22987
2 68759 1 22987
2 68760 1 22987
2 68761 1 22987
2 68762 1 23004
2 68763 1 23004
2 68764 1 23013
2 68765 1 23013
2 68766 1 23015
2 68767 1 23015
2 68768 1 23024
2 68769 1 23024
2 68770 1 23025
2 68771 1 23025
2 68772 1 23025
2 68773 1 23028
2 68774 1 23028
2 68775 1 23037
2 68776 1 23037
2 68777 1 23037
2 68778 1 23037
2 68779 1 23038
2 68780 1 23038
2 68781 1 23038
2 68782 1 23038
2 68783 1 23038
2 68784 1 23042
2 68785 1 23042
2 68786 1 23055
2 68787 1 23055
2 68788 1 23076
2 68789 1 23076
2 68790 1 23098
2 68791 1 23098
2 68792 1 23106
2 68793 1 23106
2 68794 1 23106
2 68795 1 23106
2 68796 1 23117
2 68797 1 23117
2 68798 1 23119
2 68799 1 23119
2 68800 1 23127
2 68801 1 23127
2 68802 1 23130
2 68803 1 23130
2 68804 1 23142
2 68805 1 23142
2 68806 1 23143
2 68807 1 23143
2 68808 1 23145
2 68809 1 23145
2 68810 1 23150
2 68811 1 23150
2 68812 1 23153
2 68813 1 23153
2 68814 1 23156
2 68815 1 23156
2 68816 1 23156
2 68817 1 23156
2 68818 1 23156
2 68819 1 23156
2 68820 1 23158
2 68821 1 23158
2 68822 1 23163
2 68823 1 23163
2 68824 1 23164
2 68825 1 23164
2 68826 1 23164
2 68827 1 23164
2 68828 1 23164
2 68829 1 23175
2 68830 1 23175
2 68831 1 23185
2 68832 1 23185
2 68833 1 23189
2 68834 1 23189
2 68835 1 23192
2 68836 1 23192
2 68837 1 23200
2 68838 1 23200
2 68839 1 23205
2 68840 1 23205
2 68841 1 23231
2 68842 1 23231
2 68843 1 23242
2 68844 1 23242
2 68845 1 23242
2 68846 1 23242
2 68847 1 23253
2 68848 1 23253
2 68849 1 23253
2 68850 1 23253
2 68851 1 23253
2 68852 1 23253
2 68853 1 23254
2 68854 1 23254
2 68855 1 23259
2 68856 1 23259
2 68857 1 23259
2 68858 1 23259
2 68859 1 23271
2 68860 1 23271
2 68861 1 23271
2 68862 1 23275
2 68863 1 23275
2 68864 1 23278
2 68865 1 23278
2 68866 1 23278
2 68867 1 23280
2 68868 1 23280
2 68869 1 23291
2 68870 1 23291
2 68871 1 23332
2 68872 1 23332
2 68873 1 23341
2 68874 1 23341
2 68875 1 23341
2 68876 1 23356
2 68877 1 23356
2 68878 1 23356
2 68879 1 23357
2 68880 1 23357
2 68881 1 23357
2 68882 1 23365
2 68883 1 23365
2 68884 1 23369
2 68885 1 23369
2 68886 1 23390
2 68887 1 23390
2 68888 1 23390
2 68889 1 23390
2 68890 1 23390
2 68891 1 23410
2 68892 1 23410
2 68893 1 23410
2 68894 1 23410
2 68895 1 23410
2 68896 1 23410
2 68897 1 23437
2 68898 1 23437
2 68899 1 23442
2 68900 1 23442
2 68901 1 23451
2 68902 1 23451
2 68903 1 23469
2 68904 1 23469
2 68905 1 23469
2 68906 1 23480
2 68907 1 23480
2 68908 1 23486
2 68909 1 23486
2 68910 1 23493
2 68911 1 23493
2 68912 1 23498
2 68913 1 23498
2 68914 1 23537
2 68915 1 23537
2 68916 1 23537
2 68917 1 23537
2 68918 1 23545
2 68919 1 23545
2 68920 1 23545
2 68921 1 23545
2 68922 1 23562
2 68923 1 23562
2 68924 1 23579
2 68925 1 23579
2 68926 1 23611
2 68927 1 23611
2 68928 1 23626
2 68929 1 23626
2 68930 1 23649
2 68931 1 23649
2 68932 1 23649
2 68933 1 23661
2 68934 1 23661
2 68935 1 23661
2 68936 1 23661
2 68937 1 23661
2 68938 1 23661
2 68939 1 23662
2 68940 1 23662
2 68941 1 23666
2 68942 1 23666
2 68943 1 23666
2 68944 1 23674
2 68945 1 23674
2 68946 1 23674
2 68947 1 23674
2 68948 1 23675
2 68949 1 23675
2 68950 1 23675
2 68951 1 23675
2 68952 1 23675
2 68953 1 23676
2 68954 1 23676
2 68955 1 23678
2 68956 1 23678
2 68957 1 23703
2 68958 1 23703
2 68959 1 23703
2 68960 1 23703
2 68961 1 23704
2 68962 1 23704
2 68963 1 23704
2 68964 1 23705
2 68965 1 23705
2 68966 1 23721
2 68967 1 23721
2 68968 1 23722
2 68969 1 23722
2 68970 1 23728
2 68971 1 23728
2 68972 1 23734
2 68973 1 23734
2 68974 1 23734
2 68975 1 23738
2 68976 1 23738
2 68977 1 23738
2 68978 1 23738
2 68979 1 23757
2 68980 1 23757
2 68981 1 23757
2 68982 1 23757
2 68983 1 23757
2 68984 1 23757
2 68985 1 23758
2 68986 1 23758
2 68987 1 23758
2 68988 1 23761
2 68989 1 23761
2 68990 1 23761
2 68991 1 23761
2 68992 1 23761
2 68993 1 23761
2 68994 1 23761
2 68995 1 23762
2 68996 1 23762
2 68997 1 23764
2 68998 1 23764
2 68999 1 23776
2 69000 1 23776
2 69001 1 23794
2 69002 1 23794
2 69003 1 23794
2 69004 1 23794
2 69005 1 23794
2 69006 1 23794
2 69007 1 23794
2 69008 1 23795
2 69009 1 23795
2 69010 1 23798
2 69011 1 23798
2 69012 1 23805
2 69013 1 23805
2 69014 1 23805
2 69015 1 23815
2 69016 1 23815
2 69017 1 23839
2 69018 1 23839
2 69019 1 23847
2 69020 1 23847
2 69021 1 23847
2 69022 1 23847
2 69023 1 23855
2 69024 1 23855
2 69025 1 23861
2 69026 1 23861
2 69027 1 23876
2 69028 1 23876
2 69029 1 23876
2 69030 1 23877
2 69031 1 23877
2 69032 1 23885
2 69033 1 23885
2 69034 1 23885
2 69035 1 23885
2 69036 1 23940
2 69037 1 23940
2 69038 1 23940
2 69039 1 24026
2 69040 1 24026
2 69041 1 24031
2 69042 1 24031
2 69043 1 24038
2 69044 1 24038
2 69045 1 24049
2 69046 1 24049
2 69047 1 24049
2 69048 1 24106
2 69049 1 24106
2 69050 1 24118
2 69051 1 24118
2 69052 1 24119
2 69053 1 24119
2 69054 1 24160
2 69055 1 24160
2 69056 1 24173
2 69057 1 24173
2 69058 1 24180
2 69059 1 24180
2 69060 1 24180
2 69061 1 24180
2 69062 1 24181
2 69063 1 24181
2 69064 1 24213
2 69065 1 24213
2 69066 1 24213
2 69067 1 24253
2 69068 1 24253
2 69069 1 24262
2 69070 1 24262
2 69071 1 24262
2 69072 1 24262
2 69073 1 24262
2 69074 1 24262
2 69075 1 24262
2 69076 1 24262
2 69077 1 24263
2 69078 1 24263
2 69079 1 24264
2 69080 1 24264
2 69081 1 24264
2 69082 1 24264
2 69083 1 24277
2 69084 1 24277
2 69085 1 24277
2 69086 1 24277
2 69087 1 24286
2 69088 1 24286
2 69089 1 24286
2 69090 1 24286
2 69091 1 24294
2 69092 1 24294
2 69093 1 24295
2 69094 1 24295
2 69095 1 24295
2 69096 1 24304
2 69097 1 24304
2 69098 1 24312
2 69099 1 24312
2 69100 1 24312
2 69101 1 24321
2 69102 1 24321
2 69103 1 24340
2 69104 1 24340
2 69105 1 24340
2 69106 1 24340
2 69107 1 24341
2 69108 1 24341
2 69109 1 24342
2 69110 1 24342
2 69111 1 24343
2 69112 1 24343
2 69113 1 24349
2 69114 1 24349
2 69115 1 24358
2 69116 1 24358
2 69117 1 24358
2 69118 1 24393
2 69119 1 24393
2 69120 1 24393
2 69121 1 24406
2 69122 1 24406
2 69123 1 24406
2 69124 1 24415
2 69125 1 24415
2 69126 1 24438
2 69127 1 24438
2 69128 1 24450
2 69129 1 24450
2 69130 1 24450
2 69131 1 24450
2 69132 1 24451
2 69133 1 24451
2 69134 1 24451
2 69135 1 24451
2 69136 1 24454
2 69137 1 24454
2 69138 1 24467
2 69139 1 24467
2 69140 1 24485
2 69141 1 24485
2 69142 1 24486
2 69143 1 24486
2 69144 1 24486
2 69145 1 24495
2 69146 1 24495
2 69147 1 24495
2 69148 1 24495
2 69149 1 24499
2 69150 1 24499
2 69151 1 24500
2 69152 1 24500
2 69153 1 24500
2 69154 1 24504
2 69155 1 24504
2 69156 1 24519
2 69157 1 24519
2 69158 1 24546
2 69159 1 24546
2 69160 1 24546
2 69161 1 24546
2 69162 1 24553
2 69163 1 24553
2 69164 1 24562
2 69165 1 24562
2 69166 1 24562
2 69167 1 24567
2 69168 1 24567
2 69169 1 24570
2 69170 1 24570
2 69171 1 24571
2 69172 1 24571
2 69173 1 24593
2 69174 1 24593
2 69175 1 24593
2 69176 1 24608
2 69177 1 24608
2 69178 1 24608
2 69179 1 24621
2 69180 1 24621
2 69181 1 24635
2 69182 1 24635
2 69183 1 24647
2 69184 1 24647
2 69185 1 24647
2 69186 1 24654
2 69187 1 24654
2 69188 1 24674
2 69189 1 24674
2 69190 1 24674
2 69191 1 24677
2 69192 1 24677
2 69193 1 24680
2 69194 1 24680
2 69195 1 24681
2 69196 1 24681
2 69197 1 24687
2 69198 1 24687
2 69199 1 24687
2 69200 1 24687
2 69201 1 24719
2 69202 1 24719
2 69203 1 24719
2 69204 1 24719
2 69205 1 24733
2 69206 1 24733
2 69207 1 24733
2 69208 1 24733
2 69209 1 24733
2 69210 1 24733
2 69211 1 24733
2 69212 1 24733
2 69213 1 24733
2 69214 1 24733
2 69215 1 24742
2 69216 1 24742
2 69217 1 24742
2 69218 1 24742
2 69219 1 24742
2 69220 1 24750
2 69221 1 24750
2 69222 1 24751
2 69223 1 24751
2 69224 1 24792
2 69225 1 24792
2 69226 1 24792
2 69227 1 24792
2 69228 1 24801
2 69229 1 24801
2 69230 1 24806
2 69231 1 24806
2 69232 1 24806
2 69233 1 24807
2 69234 1 24807
2 69235 1 24807
2 69236 1 24807
2 69237 1 24818
2 69238 1 24818
2 69239 1 24818
2 69240 1 24818
2 69241 1 24818
2 69242 1 24827
2 69243 1 24827
2 69244 1 24837
2 69245 1 24837
2 69246 1 24847
2 69247 1 24847
2 69248 1 24869
2 69249 1 24869
2 69250 1 24869
2 69251 1 24869
2 69252 1 24869
2 69253 1 24869
2 69254 1 24869
2 69255 1 24869
2 69256 1 24870
2 69257 1 24870
2 69258 1 24876
2 69259 1 24876
2 69260 1 24878
2 69261 1 24878
2 69262 1 24878
2 69263 1 24885
2 69264 1 24885
2 69265 1 24885
2 69266 1 24885
2 69267 1 24886
2 69268 1 24886
2 69269 1 24886
2 69270 1 24899
2 69271 1 24899
2 69272 1 24899
2 69273 1 24899
2 69274 1 24900
2 69275 1 24900
2 69276 1 24901
2 69277 1 24901
2 69278 1 24916
2 69279 1 24916
2 69280 1 24916
2 69281 1 24916
2 69282 1 24917
2 69283 1 24917
2 69284 1 24917
2 69285 1 24917
2 69286 1 24922
2 69287 1 24922
2 69288 1 24925
2 69289 1 24925
2 69290 1 24926
2 69291 1 24926
2 69292 1 24933
2 69293 1 24933
2 69294 1 24933
2 69295 1 24939
2 69296 1 24939
2 69297 1 24948
2 69298 1 24948
2 69299 1 24975
2 69300 1 24975
2 69301 1 24976
2 69302 1 24976
2 69303 1 24976
2 69304 1 24985
2 69305 1 24985
2 69306 1 24986
2 69307 1 24986
2 69308 1 24986
2 69309 1 24986
2 69310 1 24995
2 69311 1 24995
2 69312 1 25020
2 69313 1 25020
2 69314 1 25020
2 69315 1 25023
2 69316 1 25023
2 69317 1 25023
2 69318 1 25023
2 69319 1 25023
2 69320 1 25024
2 69321 1 25024
2 69322 1 25024
2 69323 1 25024
2 69324 1 25025
2 69325 1 25025
2 69326 1 25025
2 69327 1 25026
2 69328 1 25026
2 69329 1 25041
2 69330 1 25041
2 69331 1 25042
2 69332 1 25042
2 69333 1 25077
2 69334 1 25077
2 69335 1 25082
2 69336 1 25082
2 69337 1 25082
2 69338 1 25082
2 69339 1 25082
2 69340 1 25082
2 69341 1 25082
2 69342 1 25082
2 69343 1 25082
2 69344 1 25082
2 69345 1 25089
2 69346 1 25089
2 69347 1 25089
2 69348 1 25098
2 69349 1 25098
2 69350 1 25107
2 69351 1 25107
2 69352 1 25114
2 69353 1 25114
2 69354 1 25114
2 69355 1 25114
2 69356 1 25115
2 69357 1 25115
2 69358 1 25115
2 69359 1 25116
2 69360 1 25116
2 69361 1 25127
2 69362 1 25127
2 69363 1 25159
2 69364 1 25159
2 69365 1 25162
2 69366 1 25162
2 69367 1 25176
2 69368 1 25176
2 69369 1 25176
2 69370 1 25185
2 69371 1 25185
2 69372 1 25185
2 69373 1 25185
2 69374 1 25189
2 69375 1 25189
2 69376 1 25196
2 69377 1 25196
2 69378 1 25206
2 69379 1 25206
2 69380 1 25211
2 69381 1 25211
2 69382 1 25214
2 69383 1 25214
2 69384 1 25215
2 69385 1 25215
2 69386 1 25230
2 69387 1 25230
2 69388 1 25258
2 69389 1 25258
2 69390 1 25261
2 69391 1 25261
2 69392 1 25269
2 69393 1 25269
2 69394 1 25269
2 69395 1 25270
2 69396 1 25270
2 69397 1 25270
2 69398 1 25272
2 69399 1 25272
2 69400 1 25283
2 69401 1 25283
2 69402 1 25283
2 69403 1 25288
2 69404 1 25288
2 69405 1 25291
2 69406 1 25291
2 69407 1 25294
2 69408 1 25294
2 69409 1 25294
2 69410 1 25294
2 69411 1 25294
2 69412 1 25300
2 69413 1 25300
2 69414 1 25301
2 69415 1 25301
2 69416 1 25357
2 69417 1 25357
2 69418 1 25357
2 69419 1 25357
2 69420 1 25357
2 69421 1 25357
2 69422 1 25357
2 69423 1 25358
2 69424 1 25358
2 69425 1 25363
2 69426 1 25363
2 69427 1 25363
2 69428 1 25368
2 69429 1 25368
2 69430 1 25368
2 69431 1 25368
2 69432 1 25368
2 69433 1 25368
2 69434 1 25379
2 69435 1 25379
2 69436 1 25379
2 69437 1 25380
2 69438 1 25380
2 69439 1 25380
2 69440 1 25380
2 69441 1 25388
2 69442 1 25388
2 69443 1 25391
2 69444 1 25391
2 69445 1 25398
2 69446 1 25398
2 69447 1 25412
2 69448 1 25412
2 69449 1 25412
2 69450 1 25413
2 69451 1 25413
2 69452 1 25414
2 69453 1 25414
2 69454 1 25414
2 69455 1 25414
2 69456 1 25414
2 69457 1 25414
2 69458 1 25414
2 69459 1 25443
2 69460 1 25443
2 69461 1 25450
2 69462 1 25450
2 69463 1 25460
2 69464 1 25460
2 69465 1 25472
2 69466 1 25472
2 69467 1 25474
2 69468 1 25474
2 69469 1 25482
2 69470 1 25482
2 69471 1 25486
2 69472 1 25486
2 69473 1 25502
2 69474 1 25502
2 69475 1 25502
2 69476 1 25510
2 69477 1 25510
2 69478 1 25534
2 69479 1 25534
2 69480 1 25542
2 69481 1 25542
2 69482 1 25542
2 69483 1 25542
2 69484 1 25543
2 69485 1 25543
2 69486 1 25557
2 69487 1 25557
2 69488 1 25558
2 69489 1 25558
2 69490 1 25563
2 69491 1 25563
2 69492 1 25566
2 69493 1 25566
2 69494 1 25590
2 69495 1 25590
2 69496 1 25612
2 69497 1 25612
2 69498 1 25612
2 69499 1 25636
2 69500 1 25636
2 69501 1 25644
2 69502 1 25644
2 69503 1 25647
2 69504 1 25647
2 69505 1 25653
2 69506 1 25653
2 69507 1 25653
2 69508 1 25678
2 69509 1 25678
2 69510 1 25686
2 69511 1 25686
2 69512 1 25686
2 69513 1 25702
2 69514 1 25702
2 69515 1 25739
2 69516 1 25739
2 69517 1 25752
2 69518 1 25752
2 69519 1 25752
2 69520 1 25761
2 69521 1 25761
2 69522 1 25762
2 69523 1 25762
2 69524 1 25774
2 69525 1 25774
2 69526 1 25798
2 69527 1 25798
2 69528 1 25798
2 69529 1 25817
2 69530 1 25817
2 69531 1 25833
2 69532 1 25833
2 69533 1 25833
2 69534 1 25834
2 69535 1 25834
2 69536 1 25834
2 69537 1 25834
2 69538 1 25888
2 69539 1 25888
2 69540 1 25888
2 69541 1 25888
2 69542 1 25889
2 69543 1 25889
2 69544 1 25889
2 69545 1 25889
2 69546 1 25904
2 69547 1 25904
2 69548 1 25908
2 69549 1 25908
2 69550 1 25908
2 69551 1 25927
2 69552 1 25927
2 69553 1 25927
2 69554 1 25952
2 69555 1 25952
2 69556 1 25952
2 69557 1 25952
2 69558 1 25952
2 69559 1 25952
2 69560 1 25952
2 69561 1 25952
2 69562 1 25952
2 69563 1 25952
2 69564 1 25952
2 69565 1 25952
2 69566 1 25953
2 69567 1 25953
2 69568 1 25953
2 69569 1 25954
2 69570 1 25954
2 69571 1 25955
2 69572 1 25955
2 69573 1 25964
2 69574 1 25964
2 69575 1 25968
2 69576 1 25968
2 69577 1 25968
2 69578 1 25969
2 69579 1 25969
2 69580 1 25982
2 69581 1 25982
2 69582 1 25998
2 69583 1 25998
2 69584 1 26025
2 69585 1 26025
2 69586 1 26053
2 69587 1 26053
2 69588 1 26073
2 69589 1 26073
2 69590 1 26073
2 69591 1 26075
2 69592 1 26075
2 69593 1 26092
2 69594 1 26092
2 69595 1 26103
2 69596 1 26103
2 69597 1 26103
2 69598 1 26103
2 69599 1 26112
2 69600 1 26112
2 69601 1 26182
2 69602 1 26182
2 69603 1 26185
2 69604 1 26185
2 69605 1 26185
2 69606 1 26185
2 69607 1 26185
2 69608 1 26197
2 69609 1 26197
2 69610 1 26199
2 69611 1 26199
2 69612 1 26291
2 69613 1 26291
2 69614 1 26300
2 69615 1 26300
2 69616 1 26307
2 69617 1 26307
2 69618 1 26332
2 69619 1 26332
2 69620 1 26375
2 69621 1 26375
2 69622 1 26410
2 69623 1 26410
2 69624 1 26413
2 69625 1 26413
2 69626 1 26462
2 69627 1 26462
2 69628 1 26465
2 69629 1 26465
2 69630 1 26466
2 69631 1 26466
2 69632 1 26467
2 69633 1 26467
2 69634 1 26468
2 69635 1 26468
2 69636 1 26469
2 69637 1 26469
2 69638 1 26477
2 69639 1 26477
2 69640 1 26486
2 69641 1 26486
2 69642 1 26489
2 69643 1 26489
2 69644 1 26489
2 69645 1 26490
2 69646 1 26490
2 69647 1 26498
2 69648 1 26498
2 69649 1 26502
2 69650 1 26502
2 69651 1 26528
2 69652 1 26528
2 69653 1 26535
2 69654 1 26535
2 69655 1 26535
2 69656 1 26542
2 69657 1 26542
2 69658 1 26551
2 69659 1 26551
2 69660 1 26553
2 69661 1 26553
2 69662 1 26566
2 69663 1 26566
2 69664 1 26567
2 69665 1 26567
2 69666 1 26569
2 69667 1 26569
2 69668 1 26573
2 69669 1 26573
2 69670 1 26599
2 69671 1 26599
2 69672 1 26601
2 69673 1 26601
2 69674 1 26609
2 69675 1 26609
2 69676 1 26624
2 69677 1 26624
2 69678 1 26677
2 69679 1 26677
2 69680 1 26682
2 69681 1 26682
2 69682 1 26712
2 69683 1 26712
2 69684 1 26721
2 69685 1 26721
2 69686 1 26729
2 69687 1 26729
2 69688 1 26729
2 69689 1 26746
2 69690 1 26746
2 69691 1 26769
2 69692 1 26769
2 69693 1 26802
2 69694 1 26802
2 69695 1 26846
2 69696 1 26846
2 69697 1 26846
2 69698 1 26891
2 69699 1 26891
2 69700 1 26894
2 69701 1 26894
2 69702 1 26907
2 69703 1 26907
2 69704 1 26907
2 69705 1 26907
2 69706 1 26907
2 69707 1 26925
2 69708 1 26925
2 69709 1 26949
2 69710 1 26949
2 69711 1 26950
2 69712 1 26950
2 69713 1 26973
2 69714 1 26973
2 69715 1 26974
2 69716 1 26974
2 69717 1 26975
2 69718 1 26975
2 69719 1 26979
2 69720 1 26979
2 69721 1 26988
2 69722 1 26988
2 69723 1 26988
2 69724 1 26988
2 69725 1 26990
2 69726 1 26990
2 69727 1 26994
2 69728 1 26994
2 69729 1 26999
2 69730 1 26999
2 69731 1 27013
2 69732 1 27013
2 69733 1 27040
2 69734 1 27040
2 69735 1 27043
2 69736 1 27043
2 69737 1 27044
2 69738 1 27044
2 69739 1 27062
2 69740 1 27062
2 69741 1 27076
2 69742 1 27076
2 69743 1 27076
2 69744 1 27077
2 69745 1 27077
2 69746 1 27106
2 69747 1 27106
2 69748 1 27119
2 69749 1 27119
2 69750 1 27119
2 69751 1 27120
2 69752 1 27120
2 69753 1 27124
2 69754 1 27124
2 69755 1 27138
2 69756 1 27138
2 69757 1 27138
2 69758 1 27146
2 69759 1 27146
2 69760 1 27165
2 69761 1 27165
2 69762 1 27165
2 69763 1 27176
2 69764 1 27176
2 69765 1 27176
2 69766 1 27179
2 69767 1 27179
2 69768 1 27179
2 69769 1 27185
2 69770 1 27185
2 69771 1 27202
2 69772 1 27202
2 69773 1 27202
2 69774 1 27202
2 69775 1 27202
2 69776 1 27241
2 69777 1 27241
2 69778 1 27253
2 69779 1 27253
2 69780 1 27254
2 69781 1 27254
2 69782 1 27254
2 69783 1 27256
2 69784 1 27256
2 69785 1 27259
2 69786 1 27259
2 69787 1 27259
2 69788 1 27259
2 69789 1 27276
2 69790 1 27276
2 69791 1 27278
2 69792 1 27278
2 69793 1 27286
2 69794 1 27286
2 69795 1 27294
2 69796 1 27294
2 69797 1 27312
2 69798 1 27312
2 69799 1 27313
2 69800 1 27313
2 69801 1 27324
2 69802 1 27324
2 69803 1 27332
2 69804 1 27332
2 69805 1 27351
2 69806 1 27351
2 69807 1 27396
2 69808 1 27396
2 69809 1 27410
2 69810 1 27410
2 69811 1 27418
2 69812 1 27418
2 69813 1 27419
2 69814 1 27419
2 69815 1 27437
2 69816 1 27437
2 69817 1 27437
2 69818 1 27453
2 69819 1 27453
2 69820 1 27453
2 69821 1 27461
2 69822 1 27461
2 69823 1 27465
2 69824 1 27465
2 69825 1 27495
2 69826 1 27495
2 69827 1 27501
2 69828 1 27501
2 69829 1 27501
2 69830 1 27501
2 69831 1 27501
2 69832 1 27504
2 69833 1 27504
2 69834 1 27525
2 69835 1 27525
2 69836 1 27527
2 69837 1 27527
2 69838 1 27537
2 69839 1 27537
2 69840 1 27549
2 69841 1 27549
2 69842 1 27549
2 69843 1 27564
2 69844 1 27564
2 69845 1 27591
2 69846 1 27591
2 69847 1 27606
2 69848 1 27606
2 69849 1 27622
2 69850 1 27622
2 69851 1 27651
2 69852 1 27651
2 69853 1 27651
2 69854 1 27652
2 69855 1 27652
2 69856 1 27652
2 69857 1 27652
2 69858 1 27661
2 69859 1 27661
2 69860 1 27692
2 69861 1 27692
2 69862 1 27692
2 69863 1 27708
2 69864 1 27708
2 69865 1 27708
2 69866 1 27715
2 69867 1 27715
2 69868 1 27732
2 69869 1 27732
2 69870 1 27732
2 69871 1 27732
2 69872 1 27733
2 69873 1 27733
2 69874 1 27748
2 69875 1 27748
2 69876 1 27769
2 69877 1 27769
2 69878 1 27789
2 69879 1 27789
2 69880 1 27845
2 69881 1 27845
2 69882 1 27901
2 69883 1 27901
2 69884 1 27901
2 69885 1 27901
2 69886 1 27904
2 69887 1 27904
2 69888 1 27920
2 69889 1 27920
2 69890 1 27920
2 69891 1 27922
2 69892 1 27922
2 69893 1 27922
2 69894 1 27922
2 69895 1 27922
2 69896 1 27995
2 69897 1 27995
2 69898 1 27995
2 69899 1 28023
2 69900 1 28023
2 69901 1 28024
2 69902 1 28024
2 69903 1 28043
2 69904 1 28043
2 69905 1 28043
2 69906 1 28056
2 69907 1 28056
2 69908 1 28077
2 69909 1 28077
2 69910 1 28085
2 69911 1 28085
2 69912 1 28097
2 69913 1 28097
2 69914 1 28106
2 69915 1 28106
2 69916 1 28108
2 69917 1 28108
2 69918 1 28109
2 69919 1 28109
2 69920 1 28109
2 69921 1 28110
2 69922 1 28110
2 69923 1 28116
2 69924 1 28116
2 69925 1 28125
2 69926 1 28125
2 69927 1 28126
2 69928 1 28126
2 69929 1 28141
2 69930 1 28141
2 69931 1 28144
2 69932 1 28144
2 69933 1 28162
2 69934 1 28162
2 69935 1 28164
2 69936 1 28164
2 69937 1 28164
2 69938 1 28166
2 69939 1 28166
2 69940 1 28167
2 69941 1 28167
2 69942 1 28170
2 69943 1 28170
2 69944 1 28173
2 69945 1 28173
2 69946 1 28197
2 69947 1 28197
2 69948 1 28201
2 69949 1 28201
2 69950 1 28214
2 69951 1 28214
2 69952 1 28223
2 69953 1 28223
2 69954 1 28230
2 69955 1 28230
2 69956 1 28234
2 69957 1 28234
2 69958 1 28239
2 69959 1 28239
2 69960 1 28246
2 69961 1 28246
2 69962 1 28253
2 69963 1 28253
2 69964 1 28261
2 69965 1 28261
2 69966 1 28300
2 69967 1 28300
2 69968 1 28301
2 69969 1 28301
2 69970 1 28303
2 69971 1 28303
2 69972 1 28304
2 69973 1 28304
2 69974 1 28307
2 69975 1 28307
2 69976 1 28315
2 69977 1 28315
2 69978 1 28315
2 69979 1 28336
2 69980 1 28336
2 69981 1 28336
2 69982 1 28336
2 69983 1 28338
2 69984 1 28338
2 69985 1 28369
2 69986 1 28369
2 69987 1 28374
2 69988 1 28374
2 69989 1 28381
2 69990 1 28381
2 69991 1 28384
2 69992 1 28384
2 69993 1 28384
2 69994 1 28385
2 69995 1 28385
2 69996 1 28388
2 69997 1 28388
2 69998 1 28389
2 69999 1 28389
2 70000 1 28389
2 70001 1 28401
2 70002 1 28401
2 70003 1 28401
2 70004 1 28410
2 70005 1 28410
2 70006 1 28410
2 70007 1 28419
2 70008 1 28419
2 70009 1 28419
2 70010 1 28426
2 70011 1 28426
2 70012 1 28455
2 70013 1 28455
2 70014 1 28456
2 70015 1 28456
2 70016 1 28456
2 70017 1 28469
2 70018 1 28469
2 70019 1 28469
2 70020 1 28470
2 70021 1 28470
2 70022 1 28470
2 70023 1 28470
2 70024 1 28475
2 70025 1 28475
2 70026 1 28475
2 70027 1 28475
2 70028 1 28475
2 70029 1 28484
2 70030 1 28484
2 70031 1 28491
2 70032 1 28491
2 70033 1 28500
2 70034 1 28500
2 70035 1 28509
2 70036 1 28509
2 70037 1 28521
2 70038 1 28521
2 70039 1 28521
2 70040 1 28521
2 70041 1 28521
2 70042 1 28523
2 70043 1 28523
2 70044 1 28523
2 70045 1 28575
2 70046 1 28575
2 70047 1 28576
2 70048 1 28576
2 70049 1 28576
2 70050 1 28576
2 70051 1 28576
2 70052 1 28577
2 70053 1 28577
2 70054 1 28580
2 70055 1 28580
2 70056 1 28598
2 70057 1 28598
2 70058 1 28598
2 70059 1 28598
2 70060 1 28598
2 70061 1 28598
2 70062 1 28601
2 70063 1 28601
2 70064 1 28602
2 70065 1 28602
2 70066 1 28610
2 70067 1 28610
2 70068 1 28619
2 70069 1 28619
2 70070 1 28630
2 70071 1 28630
2 70072 1 28630
2 70073 1 28631
2 70074 1 28631
2 70075 1 28634
2 70076 1 28634
2 70077 1 28634
2 70078 1 28634
2 70079 1 28634
2 70080 1 28640
2 70081 1 28640
2 70082 1 28640
2 70083 1 28644
2 70084 1 28644
2 70085 1 28655
2 70086 1 28655
2 70087 1 28672
2 70088 1 28672
2 70089 1 28675
2 70090 1 28675
2 70091 1 28681
2 70092 1 28681
2 70093 1 28692
2 70094 1 28692
2 70095 1 28694
2 70096 1 28694
2 70097 1 28706
2 70098 1 28706
2 70099 1 28709
2 70100 1 28709
2 70101 1 28733
2 70102 1 28733
2 70103 1 28733
2 70104 1 28741
2 70105 1 28741
2 70106 1 28742
2 70107 1 28742
2 70108 1 28748
2 70109 1 28748
2 70110 1 28748
2 70111 1 28748
2 70112 1 28748
2 70113 1 28748
2 70114 1 28748
2 70115 1 28748
2 70116 1 28748
2 70117 1 28768
2 70118 1 28768
2 70119 1 28768
2 70120 1 28777
2 70121 1 28777
2 70122 1 28777
2 70123 1 28777
2 70124 1 28777
2 70125 1 28777
2 70126 1 28778
2 70127 1 28778
2 70128 1 28789
2 70129 1 28789
2 70130 1 28789
2 70131 1 28789
2 70132 1 28790
2 70133 1 28790
2 70134 1 28800
2 70135 1 28800
2 70136 1 28812
2 70137 1 28812
2 70138 1 28812
2 70139 1 28812
2 70140 1 28812
2 70141 1 28821
2 70142 1 28821
2 70143 1 28821
2 70144 1 28822
2 70145 1 28822
2 70146 1 28834
2 70147 1 28834
2 70148 1 28835
2 70149 1 28835
2 70150 1 28850
2 70151 1 28850
2 70152 1 28852
2 70153 1 28852
2 70154 1 28859
2 70155 1 28859
2 70156 1 28873
2 70157 1 28873
2 70158 1 28873
2 70159 1 28887
2 70160 1 28887
2 70161 1 28899
2 70162 1 28899
2 70163 1 28899
2 70164 1 28899
2 70165 1 28961
2 70166 1 28961
2 70167 1 28961
2 70168 1 28980
2 70169 1 28980
2 70170 1 28991
2 70171 1 28991
2 70172 1 28991
2 70173 1 28991
2 70174 1 28991
2 70175 1 28991
2 70176 1 28992
2 70177 1 28992
2 70178 1 28993
2 70179 1 28993
2 70180 1 29024
2 70181 1 29024
2 70182 1 29024
2 70183 1 29042
2 70184 1 29042
2 70185 1 29051
2 70186 1 29051
2 70187 1 29068
2 70188 1 29068
2 70189 1 29069
2 70190 1 29069
2 70191 1 29139
2 70192 1 29139
2 70193 1 29139
2 70194 1 29141
2 70195 1 29141
2 70196 1 29141
2 70197 1 29141
2 70198 1 29142
2 70199 1 29142
2 70200 1 29147
2 70201 1 29147
2 70202 1 29150
2 70203 1 29150
2 70204 1 29153
2 70205 1 29153
2 70206 1 29153
2 70207 1 29153
2 70208 1 29154
2 70209 1 29154
2 70210 1 29181
2 70211 1 29181
2 70212 1 29188
2 70213 1 29188
2 70214 1 29189
2 70215 1 29189
2 70216 1 29190
2 70217 1 29190
2 70218 1 29195
2 70219 1 29195
2 70220 1 29197
2 70221 1 29197
2 70222 1 29198
2 70223 1 29198
2 70224 1 29207
2 70225 1 29207
2 70226 1 29207
2 70227 1 29207
2 70228 1 29208
2 70229 1 29208
2 70230 1 29225
2 70231 1 29225
2 70232 1 29225
2 70233 1 29225
2 70234 1 29233
2 70235 1 29233
2 70236 1 29242
2 70237 1 29242
2 70238 1 29242
2 70239 1 29277
2 70240 1 29277
2 70241 1 29277
2 70242 1 29280
2 70243 1 29280
2 70244 1 29280
2 70245 1 29280
2 70246 1 29280
2 70247 1 29315
2 70248 1 29315
2 70249 1 29315
2 70250 1 29331
2 70251 1 29331
2 70252 1 29335
2 70253 1 29335
2 70254 1 29338
2 70255 1 29338
2 70256 1 29348
2 70257 1 29348
2 70258 1 29368
2 70259 1 29368
2 70260 1 29378
2 70261 1 29378
2 70262 1 29380
2 70263 1 29380
2 70264 1 29418
2 70265 1 29418
2 70266 1 29428
2 70267 1 29428
2 70268 1 29429
2 70269 1 29429
2 70270 1 29437
2 70271 1 29437
2 70272 1 29437
2 70273 1 29437
2 70274 1 29437
2 70275 1 29437
2 70276 1 29458
2 70277 1 29458
2 70278 1 29458
2 70279 1 29458
2 70280 1 29458
2 70281 1 29468
2 70282 1 29468
2 70283 1 29471
2 70284 1 29471
2 70285 1 29471
2 70286 1 29471
2 70287 1 29471
2 70288 1 29471
2 70289 1 29471
2 70290 1 29471
2 70291 1 29471
2 70292 1 29471
2 70293 1 29471
2 70294 1 29471
2 70295 1 29471
2 70296 1 29471
2 70297 1 29471
2 70298 1 29471
2 70299 1 29471
2 70300 1 29471
2 70301 1 29481
2 70302 1 29481
2 70303 1 29499
2 70304 1 29499
2 70305 1 29499
2 70306 1 29500
2 70307 1 29500
2 70308 1 29507
2 70309 1 29507
2 70310 1 29507
2 70311 1 29507
2 70312 1 29507
2 70313 1 29508
2 70314 1 29508
2 70315 1 29547
2 70316 1 29547
2 70317 1 29547
2 70318 1 29553
2 70319 1 29553
2 70320 1 29577
2 70321 1 29577
2 70322 1 29594
2 70323 1 29594
2 70324 1 29595
2 70325 1 29595
2 70326 1 29618
2 70327 1 29618
2 70328 1 29642
2 70329 1 29642
2 70330 1 29645
2 70331 1 29645
2 70332 1 29645
2 70333 1 29679
2 70334 1 29679
2 70335 1 29679
2 70336 1 29679
2 70337 1 29716
2 70338 1 29716
2 70339 1 29719
2 70340 1 29719
2 70341 1 29720
2 70342 1 29720
2 70343 1 29761
2 70344 1 29761
2 70345 1 29776
2 70346 1 29776
2 70347 1 29779
2 70348 1 29779
2 70349 1 29793
2 70350 1 29793
2 70351 1 29808
2 70352 1 29808
2 70353 1 29808
2 70354 1 29842
2 70355 1 29842
2 70356 1 29843
2 70357 1 29843
2 70358 1 29872
2 70359 1 29872
2 70360 1 29885
2 70361 1 29885
2 70362 1 29888
2 70363 1 29888
2 70364 1 29888
2 70365 1 29888
2 70366 1 29888
2 70367 1 29915
2 70368 1 29915
2 70369 1 29915
2 70370 1 29915
2 70371 1 29941
2 70372 1 29941
2 70373 1 29942
2 70374 1 29942
2 70375 1 29945
2 70376 1 29945
2 70377 1 29962
2 70378 1 29962
2 70379 1 29971
2 70380 1 29971
2 70381 1 29977
2 70382 1 29977
2 70383 1 29978
2 70384 1 29978
2 70385 1 29981
2 70386 1 29981
2 70387 1 29995
2 70388 1 29995
2 70389 1 30015
2 70390 1 30015
2 70391 1 30020
2 70392 1 30020
2 70393 1 30031
2 70394 1 30031
2 70395 1 30032
2 70396 1 30032
2 70397 1 30036
2 70398 1 30036
2 70399 1 30047
2 70400 1 30047
2 70401 1 30048
2 70402 1 30048
2 70403 1 30064
2 70404 1 30064
2 70405 1 30068
2 70406 1 30068
2 70407 1 30073
2 70408 1 30073
2 70409 1 30081
2 70410 1 30081
2 70411 1 30091
2 70412 1 30091
2 70413 1 30102
2 70414 1 30102
2 70415 1 30114
2 70416 1 30114
2 70417 1 30128
2 70418 1 30128
2 70419 1 30128
2 70420 1 30128
2 70421 1 30129
2 70422 1 30129
2 70423 1 30129
2 70424 1 30130
2 70425 1 30130
2 70426 1 30132
2 70427 1 30132
2 70428 1 30132
2 70429 1 30152
2 70430 1 30152
2 70431 1 30167
2 70432 1 30167
2 70433 1 30186
2 70434 1 30186
2 70435 1 30191
2 70436 1 30191
2 70437 1 30201
2 70438 1 30201
2 70439 1 30202
2 70440 1 30202
2 70441 1 30210
2 70442 1 30210
2 70443 1 30213
2 70444 1 30213
2 70445 1 30228
2 70446 1 30228
2 70447 1 30228
2 70448 1 30228
2 70449 1 30232
2 70450 1 30232
2 70451 1 30235
2 70452 1 30235
2 70453 1 30236
2 70454 1 30236
2 70455 1 30236
2 70456 1 30244
2 70457 1 30244
2 70458 1 30244
2 70459 1 30249
2 70460 1 30249
2 70461 1 30268
2 70462 1 30268
2 70463 1 30269
2 70464 1 30269
2 70465 1 30290
2 70466 1 30290
2 70467 1 30326
2 70468 1 30326
2 70469 1 30328
2 70470 1 30328
2 70471 1 30328
2 70472 1 30331
2 70473 1 30331
2 70474 1 30340
2 70475 1 30340
2 70476 1 30341
2 70477 1 30341
2 70478 1 30365
2 70479 1 30365
2 70480 1 30368
2 70481 1 30368
2 70482 1 30379
2 70483 1 30379
2 70484 1 30379
2 70485 1 30403
2 70486 1 30403
2 70487 1 30403
2 70488 1 30403
2 70489 1 30403
2 70490 1 30403
2 70491 1 30403
2 70492 1 30403
2 70493 1 30403
2 70494 1 30403
2 70495 1 30403
2 70496 1 30403
2 70497 1 30403
2 70498 1 30403
2 70499 1 30403
2 70500 1 30403
2 70501 1 30403
2 70502 1 30403
2 70503 1 30403
2 70504 1 30403
2 70505 1 30403
2 70506 1 30403
2 70507 1 30403
2 70508 1 30403
2 70509 1 30403
2 70510 1 30403
2 70511 1 30403
2 70512 1 30403
2 70513 1 30403
2 70514 1 30403
2 70515 1 30403
2 70516 1 30403
2 70517 1 30403
2 70518 1 30403
2 70519 1 30406
2 70520 1 30406
2 70521 1 30406
2 70522 1 30421
2 70523 1 30421
2 70524 1 30430
2 70525 1 30430
2 70526 1 30440
2 70527 1 30440
2 70528 1 30441
2 70529 1 30441
2 70530 1 30441
2 70531 1 30443
2 70532 1 30443
2 70533 1 30447
2 70534 1 30447
2 70535 1 30448
2 70536 1 30448
2 70537 1 30448
2 70538 1 30454
2 70539 1 30454
2 70540 1 30457
2 70541 1 30457
2 70542 1 30457
2 70543 1 30469
2 70544 1 30469
2 70545 1 30470
2 70546 1 30470
2 70547 1 30471
2 70548 1 30471
2 70549 1 30471
2 70550 1 30471
2 70551 1 30471
2 70552 1 30471
2 70553 1 30472
2 70554 1 30472
2 70555 1 30521
2 70556 1 30521
2 70557 1 30522
2 70558 1 30522
2 70559 1 30522
2 70560 1 30522
2 70561 1 30523
2 70562 1 30523
2 70563 1 30540
2 70564 1 30540
2 70565 1 30556
2 70566 1 30556
2 70567 1 30574
2 70568 1 30574
2 70569 1 30579
2 70570 1 30579
2 70571 1 30583
2 70572 1 30583
2 70573 1 30618
2 70574 1 30618
2 70575 1 30621
2 70576 1 30621
2 70577 1 30621
2 70578 1 30621
2 70579 1 30637
2 70580 1 30637
2 70581 1 30647
2 70582 1 30647
2 70583 1 30661
2 70584 1 30661
2 70585 1 30669
2 70586 1 30669
2 70587 1 30669
2 70588 1 30689
2 70589 1 30689
2 70590 1 30701
2 70591 1 30701
2 70592 1 30734
2 70593 1 30734
2 70594 1 30752
2 70595 1 30752
2 70596 1 30762
2 70597 1 30762
2 70598 1 30772
2 70599 1 30772
2 70600 1 30786
2 70601 1 30786
2 70602 1 30800
2 70603 1 30800
2 70604 1 30805
2 70605 1 30805
2 70606 1 30805
2 70607 1 30805
2 70608 1 30805
2 70609 1 30828
2 70610 1 30828
2 70611 1 30829
2 70612 1 30829
2 70613 1 30836
2 70614 1 30836
2 70615 1 30866
2 70616 1 30866
2 70617 1 30868
2 70618 1 30868
2 70619 1 30868
2 70620 1 30900
2 70621 1 30900
2 70622 1 30901
2 70623 1 30901
2 70624 1 30901
2 70625 1 30901
2 70626 1 30957
2 70627 1 30957
2 70628 1 30958
2 70629 1 30958
2 70630 1 31004
2 70631 1 31004
2 70632 1 31018
2 70633 1 31018
2 70634 1 31026
2 70635 1 31026
2 70636 1 31066
2 70637 1 31066
2 70638 1 31066
2 70639 1 31067
2 70640 1 31067
2 70641 1 31080
2 70642 1 31080
2 70643 1 31092
2 70644 1 31092
2 70645 1 31097
2 70646 1 31097
2 70647 1 31101
2 70648 1 31101
2 70649 1 31107
2 70650 1 31107
2 70651 1 31120
2 70652 1 31120
2 70653 1 31128
2 70654 1 31128
2 70655 1 31157
2 70656 1 31157
2 70657 1 31158
2 70658 1 31158
2 70659 1 31166
2 70660 1 31166
2 70661 1 31166
2 70662 1 31171
2 70663 1 31171
2 70664 1 31178
2 70665 1 31178
2 70666 1 31193
2 70667 1 31193
2 70668 1 31196
2 70669 1 31196
2 70670 1 31223
2 70671 1 31223
2 70672 1 31235
2 70673 1 31235
2 70674 1 31255
2 70675 1 31255
2 70676 1 31270
2 70677 1 31270
2 70678 1 31270
2 70679 1 31270
2 70680 1 31272
2 70681 1 31272
2 70682 1 31276
2 70683 1 31276
2 70684 1 31282
2 70685 1 31282
2 70686 1 31305
2 70687 1 31305
2 70688 1 31305
2 70689 1 31305
2 70690 1 31312
2 70691 1 31312
2 70692 1 31312
2 70693 1 31320
2 70694 1 31320
2 70695 1 31320
2 70696 1 31322
2 70697 1 31322
2 70698 1 31341
2 70699 1 31341
2 70700 1 31362
2 70701 1 31362
2 70702 1 31375
2 70703 1 31375
2 70704 1 31377
2 70705 1 31377
2 70706 1 31388
2 70707 1 31388
2 70708 1 31389
2 70709 1 31389
2 70710 1 31392
2 70711 1 31392
2 70712 1 31396
2 70713 1 31396
2 70714 1 31433
2 70715 1 31433
2 70716 1 31441
2 70717 1 31441
2 70718 1 31442
2 70719 1 31442
2 70720 1 31442
2 70721 1 31467
2 70722 1 31467
2 70723 1 31476
2 70724 1 31476
2 70725 1 31477
2 70726 1 31477
2 70727 1 31522
2 70728 1 31522
2 70729 1 31527
2 70730 1 31527
2 70731 1 31527
2 70732 1 31527
2 70733 1 31527
2 70734 1 31527
2 70735 1 31527
2 70736 1 31527
2 70737 1 31553
2 70738 1 31553
2 70739 1 31605
2 70740 1 31605
2 70741 1 31614
2 70742 1 31614
2 70743 1 31614
2 70744 1 31614
2 70745 1 31614
2 70746 1 31614
2 70747 1 31615
2 70748 1 31615
2 70749 1 31615
2 70750 1 31615
2 70751 1 31625
2 70752 1 31625
2 70753 1 31625
2 70754 1 31629
2 70755 1 31629
2 70756 1 31629
2 70757 1 31641
2 70758 1 31641
2 70759 1 31648
2 70760 1 31648
2 70761 1 31669
2 70762 1 31669
2 70763 1 31670
2 70764 1 31670
2 70765 1 31682
2 70766 1 31682
2 70767 1 31682
2 70768 1 31683
2 70769 1 31683
2 70770 1 31703
2 70771 1 31703
2 70772 1 31716
2 70773 1 31716
2 70774 1 31735
2 70775 1 31735
2 70776 1 31736
2 70777 1 31736
2 70778 1 31741
2 70779 1 31741
2 70780 1 31741
2 70781 1 31741
2 70782 1 31741
2 70783 1 31741
2 70784 1 31763
2 70785 1 31763
2 70786 1 31763
2 70787 1 31764
2 70788 1 31764
2 70789 1 31764
2 70790 1 31802
2 70791 1 31802
2 70792 1 31811
2 70793 1 31811
2 70794 1 31811
2 70795 1 31819
2 70796 1 31819
2 70797 1 31819
2 70798 1 31819
2 70799 1 31820
2 70800 1 31820
2 70801 1 31820
2 70802 1 31820
2 70803 1 31820
2 70804 1 31843
2 70805 1 31843
2 70806 1 31875
2 70807 1 31875
2 70808 1 31875
2 70809 1 31878
2 70810 1 31878
2 70811 1 31887
2 70812 1 31887
2 70813 1 31892
2 70814 1 31892
2 70815 1 31893
2 70816 1 31893
2 70817 1 31893
2 70818 1 31895
2 70819 1 31895
2 70820 1 31904
2 70821 1 31904
2 70822 1 31905
2 70823 1 31905
2 70824 1 31927
2 70825 1 31927
2 70826 1 31944
2 70827 1 31944
2 70828 1 31947
2 70829 1 31947
2 70830 1 31951
2 70831 1 31951
2 70832 1 31981
2 70833 1 31981
2 70834 1 31984
2 70835 1 31984
2 70836 1 31992
2 70837 1 31992
2 70838 1 32004
2 70839 1 32004
2 70840 1 32004
2 70841 1 32040
2 70842 1 32040
2 70843 1 32040
2 70844 1 32042
2 70845 1 32042
2 70846 1 32042
2 70847 1 32045
2 70848 1 32045
2 70849 1 32046
2 70850 1 32046
2 70851 1 32060
2 70852 1 32060
2 70853 1 32067
2 70854 1 32067
2 70855 1 32076
2 70856 1 32076
2 70857 1 32077
2 70858 1 32077
2 70859 1 32079
2 70860 1 32079
2 70861 1 32107
2 70862 1 32107
2 70863 1 32107
2 70864 1 32119
2 70865 1 32119
2 70866 1 32120
2 70867 1 32120
2 70868 1 32136
2 70869 1 32136
2 70870 1 32140
2 70871 1 32140
2 70872 1 32140
2 70873 1 32149
2 70874 1 32149
2 70875 1 32156
2 70876 1 32156
2 70877 1 32165
2 70878 1 32165
2 70879 1 32166
2 70880 1 32166
2 70881 1 32167
2 70882 1 32167
2 70883 1 32172
2 70884 1 32172
2 70885 1 32172
2 70886 1 32180
2 70887 1 32180
2 70888 1 32189
2 70889 1 32189
2 70890 1 32192
2 70891 1 32192
2 70892 1 32219
2 70893 1 32219
2 70894 1 32219
2 70895 1 32232
2 70896 1 32232
2 70897 1 32251
2 70898 1 32251
2 70899 1 32259
2 70900 1 32259
2 70901 1 32279
2 70902 1 32279
2 70903 1 32279
2 70904 1 32338
2 70905 1 32338
2 70906 1 32398
2 70907 1 32398
2 70908 1 32398
2 70909 1 32458
2 70910 1 32458
2 70911 1 32460
2 70912 1 32460
2 70913 1 32471
2 70914 1 32471
2 70915 1 32540
2 70916 1 32540
2 70917 1 32549
2 70918 1 32549
2 70919 1 32549
2 70920 1 32549
2 70921 1 32549
2 70922 1 32570
2 70923 1 32570
2 70924 1 32581
2 70925 1 32581
2 70926 1 32581
2 70927 1 32582
2 70928 1 32582
2 70929 1 32627
2 70930 1 32627
2 70931 1 32649
2 70932 1 32649
2 70933 1 32652
2 70934 1 32652
2 70935 1 32653
2 70936 1 32653
2 70937 1 32682
2 70938 1 32682
2 70939 1 32699
2 70940 1 32699
2 70941 1 32733
2 70942 1 32733
2 70943 1 32744
2 70944 1 32744
2 70945 1 32779
2 70946 1 32779
2 70947 1 32779
2 70948 1 32779
2 70949 1 32779
2 70950 1 32786
2 70951 1 32786
2 70952 1 32796
2 70953 1 32796
2 70954 1 32797
2 70955 1 32797
2 70956 1 32814
2 70957 1 32814
2 70958 1 32854
2 70959 1 32854
2 70960 1 32868
2 70961 1 32868
2 70962 1 32877
2 70963 1 32877
2 70964 1 32885
2 70965 1 32885
2 70966 1 32885
2 70967 1 32888
2 70968 1 32888
2 70969 1 32895
2 70970 1 32895
2 70971 1 32914
2 70972 1 32914
2 70973 1 32937
2 70974 1 32937
2 70975 1 32980
2 70976 1 32980
2 70977 1 32980
2 70978 1 32980
2 70979 1 32998
2 70980 1 32998
2 70981 1 32998
2 70982 1 33043
2 70983 1 33043
2 70984 1 33067
2 70985 1 33067
2 70986 1 33077
2 70987 1 33077
2 70988 1 33102
2 70989 1 33102
2 70990 1 33116
2 70991 1 33116
2 70992 1 33117
2 70993 1 33117
2 70994 1 33140
2 70995 1 33140
2 70996 1 33140
2 70997 1 33140
2 70998 1 33163
2 70999 1 33163
2 71000 1 33179
2 71001 1 33179
2 71002 1 33184
2 71003 1 33184
2 71004 1 33225
2 71005 1 33225
2 71006 1 33226
2 71007 1 33226
2 71008 1 33263
2 71009 1 33263
2 71010 1 33287
2 71011 1 33287
2 71012 1 33315
2 71013 1 33315
2 71014 1 33325
2 71015 1 33325
2 71016 1 33344
2 71017 1 33344
2 71018 1 33345
2 71019 1 33345
2 71020 1 33367
2 71021 1 33367
2 71022 1 33445
2 71023 1 33445
2 71024 1 33445
2 71025 1 33454
2 71026 1 33454
2 71027 1 33464
2 71028 1 33464
2 71029 1 33464
2 71030 1 33474
2 71031 1 33474
2 71032 1 33474
2 71033 1 33474
2 71034 1 33475
2 71035 1 33475
2 71036 1 33492
2 71037 1 33492
2 71038 1 33532
2 71039 1 33532
2 71040 1 33574
2 71041 1 33574
2 71042 1 33594
2 71043 1 33594
2 71044 1 33594
2 71045 1 33594
2 71046 1 33600
2 71047 1 33600
2 71048 1 33600
2 71049 1 33623
2 71050 1 33623
2 71051 1 33632
2 71052 1 33632
2 71053 1 33650
2 71054 1 33650
2 71055 1 33666
2 71056 1 33666
2 71057 1 33666
2 71058 1 33684
2 71059 1 33684
2 71060 1 33711
2 71061 1 33711
2 71062 1 33720
2 71063 1 33720
2 71064 1 33768
2 71065 1 33768
2 71066 1 33771
2 71067 1 33771
2 71068 1 33771
2 71069 1 33771
2 71070 1 33773
2 71071 1 33773
2 71072 1 33786
2 71073 1 33786
2 71074 1 33813
2 71075 1 33813
2 71076 1 33825
2 71077 1 33825
2 71078 1 33834
2 71079 1 33834
2 71080 1 33837
2 71081 1 33837
2 71082 1 33839
2 71083 1 33839
2 71084 1 33867
2 71085 1 33867
2 71086 1 33873
2 71087 1 33873
2 71088 1 33873
2 71089 1 33892
2 71090 1 33892
2 71091 1 33892
2 71092 1 33922
2 71093 1 33922
2 71094 1 33925
2 71095 1 33925
2 71096 1 33925
2 71097 1 33975
2 71098 1 33975
2 71099 1 33999
2 71100 1 33999
2 71101 1 34006
2 71102 1 34006
2 71103 1 34120
2 71104 1 34120
2 71105 1 34120
2 71106 1 34132
2 71107 1 34132
2 71108 1 34178
2 71109 1 34178
2 71110 1 34191
2 71111 1 34191
2 71112 1 34241
2 71113 1 34241
2 71114 1 34245
2 71115 1 34245
2 71116 1 34253
2 71117 1 34253
2 71118 1 34253
2 71119 1 34256
2 71120 1 34256
2 71121 1 34259
2 71122 1 34259
2 71123 1 34316
2 71124 1 34316
2 71125 1 34325
2 71126 1 34325
2 71127 1 34372
2 71128 1 34372
2 71129 1 34410
2 71130 1 34410
2 71131 1 34494
2 71132 1 34494
2 71133 1 34508
2 71134 1 34508
2 71135 1 34508
2 71136 1 34589
2 71137 1 34589
2 71138 1 34721
2 71139 1 34721
2 71140 1 34750
2 71141 1 34750
2 71142 1 34751
2 71143 1 34751
2 71144 1 34803
2 71145 1 34803
2 71146 1 34844
2 71147 1 34844
2 71148 1 34857
2 71149 1 34857
2 71150 1 34857
2 71151 1 34863
2 71152 1 34863
2 71153 1 34870
2 71154 1 34870
2 71155 1 34870
2 71156 1 34870
2 71157 1 34899
2 71158 1 34899
2 71159 1 34935
2 71160 1 34935
2 71161 1 34943
2 71162 1 34943
2 71163 1 34956
2 71164 1 34956
2 71165 1 34977
2 71166 1 34977
2 71167 1 34995
2 71168 1 34995
2 71169 1 35014
2 71170 1 35014
2 71171 1 35047
2 71172 1 35047
2 71173 1 35047
2 71174 1 35059
2 71175 1 35059
2 71176 1 35059
2 71177 1 35062
2 71178 1 35062
2 71179 1 35077
2 71180 1 35077
2 71181 1 35129
2 71182 1 35129
2 71183 1 35136
2 71184 1 35136
2 71185 1 35139
2 71186 1 35139
2 71187 1 35139
2 71188 1 35158
2 71189 1 35158
2 71190 1 35164
2 71191 1 35164
2 71192 1 35164
2 71193 1 35164
2 71194 1 35165
2 71195 1 35165
2 71196 1 35172
2 71197 1 35172
2 71198 1 35183
2 71199 1 35183
2 71200 1 35189
2 71201 1 35189
2 71202 1 35208
2 71203 1 35208
2 71204 1 35210
2 71205 1 35210
2 71206 1 35239
2 71207 1 35239
2 71208 1 35261
2 71209 1 35261
2 71210 1 35261
2 71211 1 35267
2 71212 1 35267
2 71213 1 35278
2 71214 1 35278
2 71215 1 35295
2 71216 1 35295
2 71217 1 35307
2 71218 1 35307
2 71219 1 35315
2 71220 1 35315
2 71221 1 35365
2 71222 1 35365
2 71223 1 35373
2 71224 1 35373
2 71225 1 35377
2 71226 1 35377
2 71227 1 35386
2 71228 1 35386
2 71229 1 35431
2 71230 1 35431
2 71231 1 35433
2 71232 1 35433
2 71233 1 35452
2 71234 1 35452
2 71235 1 35459
2 71236 1 35459
2 71237 1 35502
2 71238 1 35502
2 71239 1 35507
2 71240 1 35507
2 71241 1 35507
2 71242 1 35548
2 71243 1 35548
2 71244 1 35552
2 71245 1 35552
2 71246 1 35578
2 71247 1 35578
2 71248 1 35578
2 71249 1 35584
2 71250 1 35584
2 71251 1 35585
2 71252 1 35585
2 71253 1 35601
2 71254 1 35601
2 71255 1 35622
2 71256 1 35622
2 71257 1 35638
2 71258 1 35638
2 71259 1 35638
2 71260 1 35640
2 71261 1 35640
2 71262 1 35641
2 71263 1 35641
2 71264 1 35660
2 71265 1 35660
2 71266 1 35667
2 71267 1 35667
2 71268 1 35675
2 71269 1 35675
2 71270 1 35692
2 71271 1 35692
2 71272 1 35693
2 71273 1 35693
2 71274 1 35703
2 71275 1 35703
2 71276 1 35708
2 71277 1 35708
2 71278 1 35715
2 71279 1 35715
2 71280 1 35722
2 71281 1 35722
2 71282 1 35748
2 71283 1 35748
2 71284 1 35751
2 71285 1 35751
2 71286 1 35817
2 71287 1 35817
2 71288 1 35850
2 71289 1 35850
2 71290 1 35850
2 71291 1 35850
2 71292 1 35852
2 71293 1 35852
2 71294 1 35855
2 71295 1 35855
2 71296 1 35900
2 71297 1 35900
2 71298 1 35900
2 71299 1 35900
2 71300 1 35905
2 71301 1 35905
2 71302 1 35910
2 71303 1 35910
2 71304 1 35932
2 71305 1 35932
2 71306 1 35933
2 71307 1 35933
2 71308 1 35998
2 71309 1 35998
2 71310 1 36001
2 71311 1 36001
2 71312 1 36002
2 71313 1 36002
2 71314 1 36033
2 71315 1 36033
2 71316 1 36033
2 71317 1 36051
2 71318 1 36051
2 71319 1 36052
2 71320 1 36052
2 71321 1 36055
2 71322 1 36055
2 71323 1 36055
2 71324 1 36077
2 71325 1 36077
2 71326 1 36077
2 71327 1 36078
2 71328 1 36078
2 71329 1 36082
2 71330 1 36082
2 71331 1 36086
2 71332 1 36086
2 71333 1 36086
2 71334 1 36088
2 71335 1 36088
2 71336 1 36101
2 71337 1 36101
2 71338 1 36113
2 71339 1 36113
2 71340 1 36113
2 71341 1 36123
2 71342 1 36123
2 71343 1 36123
2 71344 1 36139
2 71345 1 36139
2 71346 1 36142
2 71347 1 36142
2 71348 1 36174
2 71349 1 36174
2 71350 1 36183
2 71351 1 36183
2 71352 1 36183
2 71353 1 36204
2 71354 1 36204
2 71355 1 36229
2 71356 1 36229
2 71357 1 36279
2 71358 1 36279
2 71359 1 36281
2 71360 1 36281
2 71361 1 36344
2 71362 1 36344
2 71363 1 36352
2 71364 1 36352
2 71365 1 36356
2 71366 1 36356
2 71367 1 36396
2 71368 1 36396
2 71369 1 36404
2 71370 1 36404
2 71371 1 36405
2 71372 1 36405
2 71373 1 36482
2 71374 1 36482
2 71375 1 36484
2 71376 1 36484
2 71377 1 36484
2 71378 1 36525
2 71379 1 36525
2 71380 1 36534
2 71381 1 36534
2 71382 1 36546
2 71383 1 36546
2 71384 1 36548
2 71385 1 36548
2 71386 1 36552
2 71387 1 36552
2 71388 1 36562
2 71389 1 36562
2 71390 1 36566
2 71391 1 36566
2 71392 1 36569
2 71393 1 36569
2 71394 1 36581
2 71395 1 36581
2 71396 1 36582
2 71397 1 36582
2 71398 1 36582
2 71399 1 36591
2 71400 1 36591
2 71401 1 36591
2 71402 1 36621
2 71403 1 36621
2 71404 1 36625
2 71405 1 36625
2 71406 1 36626
2 71407 1 36626
2 71408 1 36627
2 71409 1 36627
2 71410 1 36654
2 71411 1 36654
2 71412 1 36662
2 71413 1 36662
2 71414 1 36665
2 71415 1 36665
2 71416 1 36673
2 71417 1 36673
2 71418 1 36710
2 71419 1 36710
2 71420 1 36723
2 71421 1 36723
2 71422 1 36723
2 71423 1 36737
2 71424 1 36737
2 71425 1 36737
2 71426 1 36737
2 71427 1 36742
2 71428 1 36742
2 71429 1 36751
2 71430 1 36751
2 71431 1 36765
2 71432 1 36765
2 71433 1 36765
2 71434 1 36767
2 71435 1 36767
2 71436 1 36821
2 71437 1 36821
2 71438 1 36822
2 71439 1 36822
2 71440 1 36873
2 71441 1 36873
2 71442 1 36908
2 71443 1 36908
2 71444 1 36917
2 71445 1 36917
2 71446 1 36948
2 71447 1 36948
2 71448 1 36948
2 71449 1 36949
2 71450 1 36949
2 71451 1 36960
2 71452 1 36960
2 71453 1 37102
2 71454 1 37102
2 71455 1 37108
2 71456 1 37108
2 71457 1 37115
2 71458 1 37115
2 71459 1 37148
2 71460 1 37148
2 71461 1 37148
2 71462 1 37194
2 71463 1 37194
2 71464 1 37213
2 71465 1 37213
2 71466 1 37213
2 71467 1 37219
2 71468 1 37219
2 71469 1 37230
2 71470 1 37230
2 71471 1 37261
2 71472 1 37261
2 71473 1 37262
2 71474 1 37262
2 71475 1 37270
2 71476 1 37270
2 71477 1 37312
2 71478 1 37312
2 71479 1 37325
2 71480 1 37325
2 71481 1 37396
2 71482 1 37396
2 71483 1 37436
2 71484 1 37436
2 71485 1 37455
2 71486 1 37455
2 71487 1 37493
2 71488 1 37493
2 71489 1 37496
2 71490 1 37496
2 71491 1 37575
2 71492 1 37575
2 71493 1 37594
2 71494 1 37594
2 71495 1 37595
2 71496 1 37595
2 71497 1 37615
2 71498 1 37615
2 71499 1 37640
2 71500 1 37640
2 71501 1 37676
2 71502 1 37676
2 71503 1 37677
2 71504 1 37677
2 71505 1 37717
2 71506 1 37717
2 71507 1 37762
2 71508 1 37762
2 71509 1 37778
2 71510 1 37778
2 71511 1 37809
2 71512 1 37809
2 71513 1 37818
2 71514 1 37818
2 71515 1 37834
2 71516 1 37834
2 71517 1 37846
2 71518 1 37846
2 71519 1 37899
2 71520 1 37899
2 71521 1 37934
2 71522 1 37934
2 71523 1 37938
2 71524 1 37938
2 71525 1 37978
2 71526 1 37978
2 71527 1 37979
2 71528 1 37979
2 71529 1 37979
2 71530 1 37989
2 71531 1 37989
2 71532 1 37989
2 71533 1 37989
2 71534 1 38015
2 71535 1 38015
2 71536 1 38076
2 71537 1 38076
2 71538 1 38086
2 71539 1 38086
2 71540 1 38089
2 71541 1 38089
2 71542 1 38136
2 71543 1 38136
2 71544 1 38137
2 71545 1 38137
2 71546 1 38145
2 71547 1 38145
2 71548 1 38185
2 71549 1 38185
2 71550 1 38216
2 71551 1 38216
2 71552 1 38235
2 71553 1 38235
2 71554 1 38269
2 71555 1 38269
2 71556 1 38282
2 71557 1 38282
2 71558 1 38332
2 71559 1 38332
2 71560 1 38347
2 71561 1 38347
2 71562 1 38366
2 71563 1 38366
2 71564 1 38367
2 71565 1 38367
2 71566 1 38393
2 71567 1 38393
2 71568 1 38423
2 71569 1 38423
2 71570 1 38437
2 71571 1 38437
2 71572 1 38569
2 71573 1 38569
2 71574 1 38572
2 71575 1 38572
2 71576 1 38580
2 71577 1 38580
2 71578 1 38588
2 71579 1 38588
2 71580 1 38592
2 71581 1 38592
2 71582 1 38592
2 71583 1 38592
2 71584 1 38592
2 71585 1 38592
2 71586 1 38592
2 71587 1 38620
2 71588 1 38620
2 71589 1 38634
2 71590 1 38634
2 71591 1 38634
2 71592 1 38634
2 71593 1 38656
2 71594 1 38656
2 71595 1 38657
2 71596 1 38657
2 71597 1 38711
2 71598 1 38711
2 71599 1 38732
2 71600 1 38732
2 71601 1 38814
2 71602 1 38814
2 71603 1 38818
2 71604 1 38818
2 71605 1 38847
2 71606 1 38847
2 71607 1 38861
2 71608 1 38861
2 71609 1 38868
2 71610 1 38868
2 71611 1 38895
2 71612 1 38895
2 71613 1 38925
2 71614 1 38925
2 71615 1 39005
2 71616 1 39005
2 71617 1 39006
2 71618 1 39006
2 71619 1 39034
2 71620 1 39034
2 71621 1 39083
2 71622 1 39083
2 71623 1 39146
2 71624 1 39146
2 71625 1 39159
2 71626 1 39159
2 71627 1 39167
2 71628 1 39167
2 71629 1 39167
2 71630 1 39205
2 71631 1 39205
2 71632 1 39205
2 71633 1 39277
2 71634 1 39277
2 71635 1 39336
2 71636 1 39336
2 71637 1 39397
2 71638 1 39397
2 71639 1 39440
2 71640 1 39440
2 71641 1 39584
2 71642 1 39584
2 71643 1 39638
2 71644 1 39638
2 71645 1 39724
2 71646 1 39724
2 71647 1 39751
2 71648 1 39751
2 71649 1 39800
2 71650 1 39800
2 71651 1 39876
2 71652 1 39876
2 71653 1 39907
2 71654 1 39907
2 71655 1 39925
2 71656 1 39925
2 71657 1 39926
2 71658 1 39926
2 71659 1 39926
2 71660 1 39939
2 71661 1 39939
2 71662 1 40018
2 71663 1 40018
2 71664 1 40068
2 71665 1 40068
2 71666 1 40089
2 71667 1 40089
2 71668 1 40089
2 71669 1 40089
2 71670 1 40089
2 71671 1 40333
2 71672 1 40333
2 71673 1 40419
2 71674 1 40419
2 71675 1 40420
2 71676 1 40420
2 71677 1 40424
2 71678 1 40424
2 71679 1 40428
2 71680 1 40428
2 71681 1 40466
2 71682 1 40466
2 71683 1 40473
2 71684 1 40473
2 71685 1 40476
2 71686 1 40476
2 71687 1 40603
2 71688 1 40603
2 71689 1 40617
2 71690 1 40617
2 71691 1 40631
2 71692 1 40631
2 71693 1 40674
2 71694 1 40674
2 71695 1 40675
2 71696 1 40675
2 71697 1 40686
2 71698 1 40686
2 71699 1 40725
2 71700 1 40725
2 71701 1 40779
2 71702 1 40779
2 71703 1 40786
2 71704 1 40786
2 71705 1 40807
2 71706 1 40807
2 71707 1 40820
2 71708 1 40820
2 71709 1 41044
2 71710 1 41044
2 71711 1 41059
2 71712 1 41059
2 71713 1 41086
2 71714 1 41086
2 71715 1 41089
2 71716 1 41089
2 71717 1 41097
2 71718 1 41097
2 71719 1 41132
2 71720 1 41132
2 71721 1 41133
2 71722 1 41133
2 71723 1 41135
2 71724 1 41135
2 71725 1 41142
2 71726 1 41142
2 71727 1 41143
2 71728 1 41143
2 71729 1 41143
2 71730 1 41175
2 71731 1 41175
2 71732 1 41235
2 71733 1 41235
2 71734 1 41246
2 71735 1 41246
2 71736 1 41246
2 71737 1 41277
2 71738 1 41277
2 71739 1 41334
2 71740 1 41334
2 71741 1 41469
2 71742 1 41469
2 71743 1 41529
2 71744 1 41529
2 71745 1 41557
2 71746 1 41557
2 71747 1 41561
2 71748 1 41561
2 71749 1 41572
2 71750 1 41572
2 71751 1 41637
2 71752 1 41637
2 71753 1 41694
2 71754 1 41694
2 71755 1 41747
2 71756 1 41747
0 27 5 154 1 25
0 28 5 122 1 42106
0 29 5 97 1 42252
0 30 5 43 1 42361
0 31 5 184 1 42410
0 32 5 258 1 42640
0 33 5 213 1 42935
0 34 5 204 1 43184
0 35 5 89 1 43409
0 36 5 80 1 43487
0 37 5 46 1 43567
0 38 5 37 1 43607
0 39 5 125 1 43648
0 40 5 172 1 43783
0 41 5 146 1 43952
0 42 5 119 1 44129
0 43 5 107 1 44277
0 44 5 129 1 44372
0 45 5 98 1 44508
0 46 5 112 1 44604
0 47 5 127 1 44700
0 48 5 161 1 44839
0 49 5 160 1 44993
0 50 5 226 1 45131
0 51 5 146 1 45340
0 52 7 4 2 42362 46996
0 53 5 1 1 48861
0 54 7 3 2 45879 43608
0 55 5 2 1 48865
0 56 7 2 2 53 48868
0 57 5 12 1 48870
0 58 7 32 2 26 43410
0 59 5 3 1 48884
0 60 7 7 2 44373 48885
0 61 7 25 2 44509 47929
0 62 7 22 2 45132 45341
0 63 5 9 1 48951
0 64 7 3 2 46364 43953
0 65 7 1 2 48952 48982
0 66 5 1 1 65
0 67 7 26 2 48489 45342
0 68 5 1 1 48985
0 69 7 4 2 44130 48986
0 70 5 2 1 49011
0 71 7 1 2 46365 49015
0 72 5 1 1 71
0 73 7 45 2 44131 48715
0 74 5 39 1 49017
0 75 7 5 2 45133 49062
0 76 5 8 1 49101
0 77 7 1 2 42936 49106
0 78 5 2 1 77
0 79 7 1 2 47330 49114
0 80 7 1 2 72 79
0 81 5 1 1 80
0 82 7 1 2 66 81
0 83 5 1 1 82
0 84 7 1 2 43185 83
0 85 5 1 1 84
0 86 7 10 2 46577 43954
0 87 5 2 1 49116
0 88 7 56 2 47476 45343
0 89 5 60 1 49128
0 90 7 2 2 49117 49129
0 91 5 3 1 49244
0 92 7 3 2 48490 49245
0 93 5 2 1 49249
0 94 7 1 2 46366 49250
0 95 5 2 1 94
0 96 7 1 2 85 49254
0 97 5 1 1 96
0 98 7 1 2 44994 97
0 99 5 1 1 98
0 100 7 57 2 46367 47331
0 101 5 58 1 49256
0 102 7 22 2 48329 45134
0 103 5 3 1 49371
0 104 7 5 2 49130 49372
0 105 5 6 1 49396
0 106 7 2 2 46578 49397
0 107 5 1 1 49407
0 108 7 1 2 49257 49408
0 109 5 1 1 108
0 110 7 1 2 99 109
0 111 5 1 1 110
0 112 7 1 2 48168 111
0 113 5 1 1 112
0 114 7 3 2 42937 45344
0 115 5 2 1 49409
0 116 7 14 2 44995 48716
0 117 5 1 1 49414
0 118 7 4 2 44132 49415
0 119 5 1 1 49428
0 120 7 1 2 49412 119
0 121 5 1 1 120
0 122 7 1 2 42411 121
0 123 5 1 1 122
0 124 7 13 2 43955 48330
0 125 5 1 1 49432
0 126 7 8 2 48491 49433
0 127 7 5 2 46368 49018
0 128 5 2 1 49453
0 129 7 1 2 49413 49458
0 130 5 3 1 129
0 131 7 1 2 49445 49460
0 132 5 1 1 131
0 133 7 1 2 123 132
0 134 5 1 1 133
0 135 7 1 2 43186 134
0 136 5 1 1 135
0 137 7 4 2 42412 49313
0 138 5 2 1 49463
0 139 7 7 2 42938 48331
0 140 5 2 1 49469
0 141 7 11 2 43956 48717
0 142 5 3 1 49478
0 143 7 1 2 49470 49479
0 144 5 2 1 143
0 145 7 1 2 49467 49492
0 146 5 1 1 145
0 147 7 8 2 46579 48492
0 148 7 1 2 146 49494
0 149 5 1 1 148
0 150 7 19 2 42939 48718
0 151 5 6 1 49502
0 152 7 4 2 46580 49503
0 153 5 2 1 49527
0 154 7 1 2 44996 49531
0 155 5 1 1 154
0 156 7 13 2 43187 49019
0 157 5 10 1 49533
0 158 7 1 2 42413 49546
0 159 7 1 2 155 158
0 160 5 1 1 159
0 161 7 1 2 149 160
0 162 7 1 2 136 161
0 163 5 1 1 162
0 164 7 1 2 44840 163
0 165 5 1 1 164
0 166 7 21 2 44997 45135
0 167 5 1 1 49556
0 168 7 3 2 49131 49557
0 169 7 8 2 42414 42940
0 170 7 1 2 49118 49580
0 171 7 1 2 49577 170
0 172 5 1 1 171
0 173 7 1 2 165 172
0 174 7 1 2 113 173
0 175 5 1 1 174
0 176 7 1 2 43649 175
0 177 5 1 1 176
0 178 7 6 2 46581 48719
0 179 5 3 1 49588
0 180 7 7 2 42941 44841
0 181 5 1 1 49597
0 182 7 1 2 49446 49598
0 183 5 1 1 182
0 184 7 21 2 44133 48493
0 185 5 9 1 49604
0 186 7 1 2 47332 49625
0 187 5 3 1 186
0 188 7 27 2 48169 44998
0 189 5 2 1 49637
0 190 7 54 2 43957 48494
0 191 5 54 1 49666
0 192 7 10 2 46369 49720
0 193 5 8 1 49774
0 194 7 1 2 49638 49775
0 195 7 1 2 49634 194
0 196 5 1 1 195
0 197 7 1 2 183 196
0 198 5 1 1 197
0 199 7 1 2 49589 198
0 200 5 1 1 199
0 201 7 10 2 44842 48495
0 202 7 1 2 49434 49792
0 203 5 1 1 202
0 204 7 9 2 47333 44999
0 205 7 18 2 48170 45136
0 206 5 1 1 49811
0 207 7 1 2 49802 49812
0 208 5 2 1 207
0 209 7 1 2 203 49829
0 210 5 6 1 209
0 211 7 8 2 43188 45345
0 212 5 2 1 49837
0 213 7 1 2 42942 49838
0 214 7 1 2 49831 213
0 215 5 1 1 214
0 216 7 1 2 200 215
0 217 5 1 1 216
0 218 7 1 2 42415 217
0 219 5 1 1 218
0 220 7 16 2 48332 48496
0 221 5 4 1 49847
0 222 7 4 2 48171 49848
0 223 7 12 2 43958 44134
0 224 5 2 1 49871
0 225 7 5 2 42943 49872
0 226 5 1 1 49885
0 227 7 10 2 45922 43189
0 228 7 3 2 47033 49890
0 229 7 1 2 49886 49900
0 230 7 1 2 49867 229
0 231 5 1 1 230
0 232 7 1 2 219 231
0 233 7 1 2 177 232
0 234 5 1 1 233
0 235 7 1 2 48041 234
0 236 5 1 1 235
0 237 7 21 2 46370 46582
0 238 5 2 1 49903
0 239 7 2 2 48042 49558
0 240 7 1 2 49904 49926
0 241 5 1 1 240
0 242 7 105 2 43190 44135
0 243 5 88 1 49928
0 244 7 3 2 46371 50033
0 245 5 11 1 50121
0 246 7 3 2 44701 49849
0 247 7 1 2 42416 50135
0 248 7 1 2 50124 247
0 249 5 1 1 248
0 250 7 1 2 241 249
0 251 5 1 1 250
0 252 7 1 2 43959 251
0 253 5 1 1 252
0 254 7 6 2 47334 48043
0 255 7 4 2 45000 50138
0 256 7 21 2 42944 46583
0 257 5 1 1 50148
0 258 7 2 2 45137 50149
0 259 5 1 1 50169
0 260 7 6 2 46372 44136
0 261 5 4 1 50171
0 262 7 7 2 46584 45138
0 263 5 3 1 50181
0 264 7 7 2 43191 48497
0 265 5 2 1 50191
0 266 7 1 2 50188 50198
0 267 7 1 2 50172 266
0 268 5 1 1 267
0 269 7 1 2 259 268
0 270 5 1 1 269
0 271 7 1 2 50144 270
0 272 5 1 1 271
0 273 7 1 2 253 272
0 274 5 1 1 273
0 275 7 9 2 48172 48720
0 276 7 1 2 43650 50200
0 277 7 1 2 274 276
0 278 5 1 1 277
0 279 7 1 2 236 278
0 280 5 1 1 279
0 281 7 1 2 48926 280
0 282 5 1 1 281
0 283 7 7 2 47034 45346
0 284 7 17 2 45001 48498
0 285 5 3 1 50216
0 286 7 6 2 43960 50217
0 287 5 4 1 50236
0 288 7 7 2 47335 49373
0 289 5 2 1 50246
0 290 7 1 2 50242 50253
0 291 5 9 1 290
0 292 7 7 2 47477 49905
0 293 7 1 2 50255 50264
0 294 5 1 1 293
0 295 7 8 2 43192 45139
0 296 5 4 1 50271
0 297 7 6 2 42945 44137
0 298 5 1 1 50283
0 299 7 2 2 50272 50284
0 300 5 1 1 50289
0 301 7 1 2 49803 50290
0 302 5 1 1 301
0 303 7 1 2 294 302
0 304 5 2 1 303
0 305 7 1 2 50209 50291
0 306 5 1 1 305
0 307 7 5 2 47035 44138
0 308 7 2 2 43193 50293
0 309 5 2 1 50298
0 310 7 5 2 46373 49132
0 311 5 2 1 50302
0 312 7 1 2 49119 50303
0 313 5 2 1 312
0 314 7 1 2 50300 50309
0 315 5 1 1 314
0 316 7 1 2 48499 315
0 317 5 1 1 316
0 318 7 3 2 47336 48953
0 319 5 1 1 50311
0 320 7 1 2 43651 319
0 321 5 1 1 320
0 322 7 1 2 49314 49929
0 323 7 1 2 321 322
0 324 5 1 1 323
0 325 7 1 2 317 324
0 326 5 1 1 325
0 327 7 1 2 45002 326
0 328 5 1 1 327
0 329 7 3 2 45003 49721
0 330 5 7 1 50314
0 331 7 2 2 47036 50034
0 332 7 1 2 50317 50324
0 333 5 1 1 332
0 334 7 11 2 47337 45347
0 335 5 2 1 50326
0 336 7 3 2 50265 50327
0 337 5 2 1 50339
0 338 7 1 2 43652 50342
0 339 5 1 1 338
0 340 7 1 2 49374 339
0 341 5 1 1 340
0 342 7 1 2 333 341
0 343 7 1 2 328 342
0 344 5 1 1 343
0 345 7 1 2 45923 344
0 346 5 1 1 345
0 347 7 1 2 306 346
0 348 5 1 1 347
0 349 7 30 2 47831 44605
0 350 7 9 2 44702 44843
0 351 7 2 2 50344 50374
0 352 7 1 2 348 50383
0 353 5 1 1 352
0 354 7 1 2 282 353
0 355 5 1 1 354
0 356 7 1 2 42641 355
0 357 5 1 1 356
0 358 7 1 2 49393 50243
0 359 5 2 1 358
0 360 7 1 2 42946 50385
0 361 5 3 1 360
0 362 7 1 2 49521 49850
0 363 5 1 1 362
0 364 7 1 2 50387 363
0 365 5 1 1 364
0 366 7 55 2 45924 47037
0 367 5 37 1 50390
0 368 7 4 2 47832 50391
0 369 7 26 2 44606 44703
0 370 5 1 1 50486
0 371 7 5 2 50482 50487
0 372 5 1 1 50512
0 373 7 1 2 365 50513
0 374 5 1 1 373
0 375 7 6 2 48333 49722
0 376 5 1 1 50517
0 377 7 2 2 50244 376
0 378 5 2 1 50523
0 379 7 56 2 47338 45140
0 380 5 42 1 50527
0 381 7 9 2 42947 50583
0 382 5 6 1 50625
0 383 7 1 2 49863 50626
0 384 5 1 1 383
0 385 7 1 2 50524 384
0 386 5 2 1 385
0 387 7 25 2 47930 48044
0 388 7 9 2 43653 44510
0 389 7 4 2 50642 50667
0 390 7 3 2 42417 48721
0 391 5 2 1 50680
0 392 7 1 2 50676 50681
0 393 7 1 2 50640 392
0 394 5 1 1 393
0 395 7 1 2 374 394
0 396 5 1 1 395
0 397 7 1 2 44139 396
0 398 5 1 1 397
0 399 7 1 2 43654 50318
0 400 7 2 2 44511 49581
0 401 7 2 2 45348 50643
0 402 7 1 2 50685 50687
0 403 7 1 2 399 402
0 404 5 1 1 403
0 405 7 1 2 398 404
0 406 5 1 1 405
0 407 7 1 2 43194 406
0 408 5 1 1 407
0 409 7 1 2 45004 49522
0 410 5 2 1 409
0 411 7 3 2 42418 50677
0 412 5 1 1 50691
0 413 7 1 2 50689 50692
0 414 5 1 1 413
0 415 7 7 2 44704 48334
0 416 7 3 2 44607 50694
0 417 7 1 2 50701 50483
0 418 5 1 1 417
0 419 7 1 2 414 418
0 420 5 1 1 419
0 421 7 1 2 46585 420
0 422 5 1 1 421
0 423 7 3 2 45925 50345
0 424 7 3 2 47038 47478
0 425 7 1 2 50695 50707
0 426 7 1 2 50704 425
0 427 5 1 1 426
0 428 7 1 2 422 427
0 429 5 1 1 428
0 430 7 1 2 49667 429
0 431 5 1 1 430
0 432 7 2 2 42419 50150
0 433 7 5 2 48722 50644
0 434 7 6 2 43655 48335
0 435 7 1 2 44512 50717
0 436 7 1 2 50712 435
0 437 7 1 2 50710 436
0 438 5 1 1 437
0 439 7 1 2 431 438
0 440 7 1 2 408 439
0 441 5 1 1 440
0 442 7 1 2 44844 441
0 443 5 1 1 442
0 444 7 87 2 46586 47479
0 445 5 78 1 50723
0 446 7 3 2 43961 50810
0 447 5 5 1 50888
0 448 7 1 2 412 372
0 449 5 5 1 448
0 450 7 1 2 50891 50896
0 451 5 1 1 450
0 452 7 8 2 44705 50346
0 453 7 13 2 45926 46374
0 454 7 3 2 47039 50909
0 455 7 1 2 50901 50922
0 456 5 1 1 455
0 457 7 1 2 451 456
0 458 5 1 1 457
0 459 7 1 2 45141 458
0 460 5 1 1 459
0 461 7 43 2 42948 43962
0 462 5 77 1 50925
0 463 7 2 2 50724 50968
0 464 5 1 1 51045
0 465 7 1 2 50514 51046
0 466 5 1 1 465
0 467 7 1 2 460 466
0 468 5 1 1 467
0 469 7 1 2 45349 468
0 470 5 1 1 469
0 471 7 6 2 44706 45142
0 472 7 2 2 50347 51047
0 473 7 9 2 46375 47040
0 474 7 5 2 45927 47339
0 475 7 2 2 51055 51064
0 476 7 1 2 51053 51069
0 477 5 1 1 476
0 478 7 2 2 49784 50584
0 479 5 20 1 51071
0 480 7 1 2 50515 51073
0 481 5 1 1 480
0 482 7 13 2 46376 43656
0 483 7 3 2 42420 51093
0 484 7 2 2 48927 50139
0 485 7 1 2 51106 51109
0 486 5 1 1 485
0 487 7 1 2 481 486
0 488 5 1 1 487
0 489 7 1 2 50035 488
0 490 5 1 1 489
0 491 7 1 2 477 490
0 492 7 1 2 470 491
0 493 5 1 1 492
0 494 7 1 2 49639 493
0 495 5 1 1 494
0 496 7 1 2 443 495
0 497 7 1 2 357 496
0 498 5 1 1 497
0 499 7 1 2 43488 498
0 500 5 1 1 499
0 501 7 51 2 42421 43657
0 502 5 30 1 51111
0 503 7 4 2 46587 49063
0 504 5 9 1 51192
0 505 7 10 2 49184 51196
0 506 5 27 1 51205
0 507 7 16 2 48045 44845
0 508 7 3 2 51215 51242
0 509 7 1 2 51112 51258
0 510 5 1 1 509
0 511 7 13 2 48173 48336
0 512 7 19 2 44707 51113
0 513 5 2 1 51274
0 514 7 11 2 48046 50392
0 515 5 1 1 51295
0 516 7 1 2 51293 515
0 517 5 18 1 516
0 518 7 2 2 51261 51306
0 519 7 25 2 42949 43195
0 520 5 2 1 51326
0 521 7 5 2 44140 51327
0 522 7 1 2 51324 51353
0 523 5 1 1 522
0 524 7 1 2 510 523
0 525 5 1 1 524
0 526 7 1 2 48500 525
0 527 5 1 1 526
0 528 7 10 2 43196 43658
0 529 7 4 2 42422 51358
0 530 7 11 2 44846 45143
0 531 7 7 2 44141 48047
0 532 7 1 2 51372 51383
0 533 7 1 2 51368 532
0 534 5 1 1 533
0 535 7 1 2 527 534
0 536 5 1 1 535
0 537 7 1 2 43963 536
0 538 5 1 1 537
0 539 7 23 2 42950 45144
0 540 5 4 1 51390
0 541 7 2 2 50233 51413
0 542 5 3 1 51417
0 543 7 1 2 49930 51419
0 544 5 1 1 543
0 545 7 5 2 48501 49185
0 546 5 21 1 51422
0 547 7 2 2 51197 51423
0 548 5 5 1 51448
0 549 7 1 2 48337 51450
0 550 5 1 1 549
0 551 7 1 2 544 550
0 552 5 1 1 551
0 553 7 1 2 51114 51243
0 554 7 1 2 552 553
0 555 5 1 1 554
0 556 7 1 2 538 555
0 557 5 1 1 556
0 558 7 1 2 42642 557
0 559 5 1 1 558
0 560 7 5 2 46377 50528
0 561 5 10 1 51455
0 562 7 11 2 49723 50634
0 563 5 3 1 51470
0 564 7 1 2 50036 51471
0 565 5 2 1 564
0 566 7 1 2 51460 51484
0 567 5 1 1 566
0 568 7 2 2 45005 567
0 569 7 2 2 48723 51461
0 570 7 1 2 50811 51488
0 571 5 1 1 570
0 572 7 3 2 51486 571
0 573 5 1 1 51490
0 574 7 1 2 48174 573
0 575 5 1 1 574
0 576 7 18 2 46378 48502
0 577 5 1 1 51493
0 578 7 2 2 48338 51494
0 579 5 1 1 51511
0 580 7 1 2 50388 579
0 581 5 1 1 580
0 582 7 1 2 49931 581
0 583 5 1 1 582
0 584 7 3 2 43197 49186
0 585 5 4 1 51513
0 586 7 14 2 49064 51516
0 587 5 2 1 51520
0 588 7 4 2 48503 51521
0 589 5 4 1 51536
0 590 7 1 2 49435 51537
0 591 5 1 1 590
0 592 7 1 2 44847 591
0 593 7 1 2 583 592
0 594 5 1 1 593
0 595 7 7 2 48048 51115
0 596 7 1 2 594 51544
0 597 7 1 2 575 596
0 598 5 1 1 597
0 599 7 1 2 559 598
0 600 5 2 1 599
0 601 7 21 2 47833 47931
0 602 7 1 2 46870 51553
0 603 7 1 2 51551 602
0 604 5 1 1 603
0 605 7 1 2 500 604
0 606 5 1 1 605
0 607 7 1 2 42107 606
0 608 5 1 1 607
0 609 7 2 2 47932 51116
0 610 7 50 2 43489 44513
0 611 5 7 1 51576
0 612 7 4 2 44848 45350
0 613 7 4 2 48049 51633
0 614 5 1 1 51637
0 615 7 5 2 44142 44708
0 616 7 1 2 49504 51262
0 617 7 1 2 51641 616
0 618 5 1 1 617
0 619 7 1 2 614 618
0 620 5 1 1 619
0 621 7 1 2 43198 620
0 622 5 1 1 621
0 623 7 3 2 46588 48050
0 624 7 3 2 48724 51646
0 625 7 1 2 44849 51649
0 626 5 1 1 625
0 627 7 1 2 622 626
0 628 5 1 1 627
0 629 7 1 2 51577 628
0 630 5 1 1 629
0 631 7 42 2 46871 47834
0 632 5 1 1 51652
0 633 7 3 2 42951 51653
0 634 5 1 1 51694
0 635 7 1 2 51259 51695
0 636 5 1 1 635
0 637 7 1 2 630 636
0 638 5 1 1 637
0 639 7 1 2 42643 638
0 640 5 1 1 639
0 641 7 2 2 46589 51578
0 642 5 1 1 51697
0 643 7 13 2 48725 50812
0 644 5 7 1 51699
0 645 7 19 2 50037 51712
0 646 5 38 1 51719
0 647 7 4 2 47835 51720
0 648 7 2 2 46872 51776
0 649 5 1 1 51780
0 650 7 1 2 642 649
0 651 5 1 1 650
0 652 7 1 2 42952 651
0 653 5 1 1 652
0 654 7 4 2 49594 49845
0 655 5 23 1 51782
0 656 7 2 2 51579 51786
0 657 5 2 1 51809
0 658 7 1 2 653 51811
0 659 5 1 1 658
0 660 7 1 2 48339 51244
0 661 7 1 2 659 660
0 662 5 1 1 661
0 663 7 1 2 640 662
0 664 5 1 1 663
0 665 7 1 2 42108 664
0 666 5 1 1 665
0 667 7 9 2 45660 42953
0 668 7 6 2 47836 51813
0 669 5 2 1 51822
0 670 7 5 2 46106 45006
0 671 5 11 1 51830
0 672 7 1 2 43490 51835
0 673 7 1 2 51823 672
0 674 7 1 2 51260 673
0 675 5 1 1 674
0 676 7 1 2 666 675
0 677 5 1 1 676
0 678 7 1 2 51574 677
0 679 5 1 1 678
0 680 7 20 2 42109 47837
0 681 7 1 2 50393 51836
0 682 7 1 2 51846 681
0 683 7 4 2 43491 44608
0 684 7 4 2 50375 51866
0 685 7 6 2 42954 50038
0 686 5 3 1 51874
0 687 7 1 2 51870 51875
0 688 7 1 2 682 687
0 689 5 1 1 688
0 690 7 1 2 679 689
0 691 5 1 1 690
0 692 7 1 2 50585 691
0 693 5 1 1 692
0 694 7 10 2 43492 47933
0 695 7 62 2 45661 47838
0 696 5 1 1 51893
0 697 7 1 2 51883 51894
0 698 7 1 2 51552 697
0 699 5 1 1 698
0 700 7 1 2 693 699
0 701 7 1 2 608 700
0 702 5 1 1 701
0 703 7 1 2 43784 702
0 704 5 1 1 703
0 705 7 30 2 42644 43785
0 706 5 24 1 51955
0 707 7 40 2 46107 47158
0 708 5 20 1 52009
0 709 7 13 2 45145 50969
0 710 5 5 1 52069
0 711 7 21 2 49315 52082
0 712 7 2 2 52049 52087
0 713 5 1 1 52108
0 714 7 3 2 51985 713
0 715 5 4 1 52110
0 716 7 7 2 48051 48340
0 717 7 4 2 47934 52117
0 718 7 12 2 43659 48175
0 719 7 1 2 52124 52128
0 720 7 1 2 51216 719
0 721 7 2 2 52111 720
0 722 7 8 2 42423 46873
0 723 7 1 2 52140 52142
0 724 5 1 1 723
0 725 7 23 2 44709 48176
0 726 7 2 2 48341 51986
0 727 5 1 1 52173
0 728 7 7 2 47480 45146
0 729 5 7 1 52175
0 730 7 6 2 46590 52176
0 731 5 4 1 52189
0 732 7 3 2 464 52083
0 733 5 2 1 52199
0 734 7 1 2 52195 52200
0 735 5 1 1 734
0 736 7 3 2 45351 735
0 737 5 1 1 52204
0 738 7 1 2 46108 52205
0 739 5 1 1 738
0 740 7 1 2 51485 739
0 741 5 1 1 740
0 742 7 1 2 52174 741
0 743 5 1 1 742
0 744 7 3 2 48342 49316
0 745 5 6 1 52207
0 746 7 2 2 46109 52210
0 747 7 9 2 48504 49932
0 748 7 1 2 52216 52218
0 749 5 1 1 748
0 750 7 3 2 43786 49317
0 751 5 13 1 52227
0 752 7 1 2 48343 52202
0 753 5 1 1 752
0 754 7 5 2 43199 49605
0 755 5 7 1 52243
0 756 7 1 2 49258 52244
0 757 5 1 1 756
0 758 7 1 2 753 757
0 759 5 1 1 758
0 760 7 1 2 47159 759
0 761 5 1 1 760
0 762 7 1 2 49375 50725
0 763 5 1 1 762
0 764 7 2 2 49933 50218
0 765 5 6 1 52255
0 766 7 1 2 763 52257
0 767 7 1 2 761 766
0 768 5 1 1 767
0 769 7 1 2 52230 768
0 770 5 1 1 769
0 771 7 1 2 749 770
0 772 5 1 1 771
0 773 7 1 2 45352 772
0 774 5 1 1 773
0 775 7 1 2 743 774
0 776 5 1 1 775
0 777 7 1 2 52150 776
0 778 5 1 1 777
0 779 7 10 2 48052 45147
0 780 7 10 2 45007 45353
0 781 5 1 1 52273
0 782 7 5 2 44850 52274
0 783 7 2 2 52263 52283
0 784 7 1 2 49259 50726
0 785 7 1 2 51987 784
0 786 7 1 2 52288 785
0 787 5 1 1 786
0 788 7 1 2 778 787
0 789 5 1 1 788
0 790 7 1 2 50394 789
0 791 5 1 1 790
0 792 7 15 2 48726 49934
0 793 5 5 1 52290
0 794 7 15 2 46591 49133
0 795 5 11 1 52310
0 796 7 3 2 48505 52325
0 797 5 2 1 52336
0 798 7 4 2 52305 52339
0 799 5 4 1 52341
0 800 7 1 2 45008 52342
0 801 5 2 1 800
0 802 7 5 2 47481 48954
0 803 5 8 1 52351
0 804 7 1 2 48344 52356
0 805 5 3 1 804
0 806 7 29 2 48506 48727
0 807 5 6 1 52367
0 808 7 7 2 44143 52368
0 809 5 3 1 52402
0 810 7 1 2 45009 52409
0 811 5 1 1 810
0 812 7 1 2 43200 811
0 813 5 1 1 812
0 814 7 2 2 52364 813
0 815 7 1 2 47340 52412
0 816 5 1 1 815
0 817 7 1 2 52349 816
0 818 5 1 1 817
0 819 7 1 2 46379 818
0 820 5 1 1 819
0 821 7 1 2 47341 52343
0 822 5 1 1 821
0 823 7 3 2 49134 50182
0 824 5 3 1 52414
0 825 7 1 2 822 52417
0 826 5 3 1 825
0 827 7 1 2 45010 52420
0 828 5 1 1 827
0 829 7 1 2 820 828
0 830 5 1 1 829
0 831 7 3 2 50395 51245
0 832 5 1 1 52423
0 833 7 1 2 830 52424
0 834 5 1 1 833
0 835 7 4 2 47041 48345
0 836 5 1 1 52426
0 837 7 7 2 45928 48177
0 838 5 1 1 52430
0 839 7 1 2 52427 52431
0 840 5 2 1 839
0 841 7 3 2 45011 51472
0 842 7 2 2 44851 52439
0 843 7 1 2 51117 52442
0 844 5 1 1 843
0 845 7 1 2 52437 844
0 846 5 1 1 845
0 847 7 1 2 50039 846
0 848 5 1 1 847
0 849 7 14 2 44852 45012
0 850 7 2 2 42424 52444
0 851 5 1 1 52458
0 852 7 5 2 50529 51094
0 853 7 1 2 52459 52460
0 854 5 1 1 853
0 855 7 4 2 47042 48178
0 856 5 2 1 52465
0 857 7 1 2 49436 49599
0 858 5 1 1 857
0 859 7 1 2 52469 858
0 860 5 1 1 859
0 861 7 1 2 45929 860
0 862 5 1 1 861
0 863 7 21 2 44853 48346
0 864 5 3 1 52471
0 865 7 17 2 42955 47043
0 866 7 3 2 43964 52495
0 867 7 1 2 52472 52512
0 868 5 1 1 867
0 869 7 1 2 862 868
0 870 5 1 1 869
0 871 7 1 2 52219 870
0 872 5 1 1 871
0 873 7 6 2 47044 44854
0 874 5 1 1 52515
0 875 7 3 2 42425 52129
0 876 5 1 1 52521
0 877 7 1 2 874 876
0 878 7 1 2 50292 877
0 879 5 1 1 878
0 880 7 1 2 872 879
0 881 5 1 1 880
0 882 7 1 2 45354 881
0 883 5 1 1 882
0 884 7 1 2 854 883
0 885 7 1 2 848 884
0 886 5 1 1 885
0 887 7 1 2 44710 886
0 888 5 1 1 887
0 889 7 1 2 834 888
0 890 5 1 1 889
0 891 7 1 2 52010 890
0 892 5 1 1 891
0 893 7 1 2 791 892
0 894 5 1 1 893
0 895 7 1 2 51867 894
0 896 5 1 1 895
0 897 7 1 2 724 896
0 898 5 1 1 897
0 899 7 1 2 42110 898
0 900 5 1 1 899
0 901 7 4 2 45662 42426
0 902 7 4 2 43493 52524
0 903 7 1 2 52528 52141
0 904 5 1 1 903
0 905 7 5 2 43660 47935
0 906 7 3 2 48053 52532
0 907 7 4 2 52143 52537
0 908 5 1 1 52540
0 909 7 3 2 43494 50488
0 910 7 2 2 50396 52544
0 911 5 1 1 52547
0 912 7 1 2 908 911
0 913 5 1 1 912
0 914 7 1 2 42111 913
0 915 5 1 1 914
0 916 7 5 2 45663 43495
0 917 5 1 1 52549
0 918 7 2 2 42427 52550
0 919 7 2 2 52538 52554
0 920 5 1 1 52556
0 921 7 1 2 915 920
0 922 5 1 1 921
0 923 7 9 2 48179 48507
0 924 5 1 1 52558
0 925 7 35 2 47160 45013
0 926 5 54 1 52567
0 927 7 2 2 47161 50970
0 928 5 11 1 52656
0 929 7 3 2 45014 50971
0 930 5 6 1 52669
0 931 7 2 2 52658 52672
0 932 5 4 1 52678
0 933 7 6 2 52602 52679
0 934 5 4 1 52684
0 935 7 3 2 46380 52568
0 936 5 1 1 52694
0 937 7 1 2 42645 936
0 938 5 1 1 937
0 939 7 5 2 52690 938
0 940 7 2 2 52559 52697
0 941 5 1 1 52702
0 942 7 5 2 43965 44855
0 943 7 5 2 42956 48508
0 944 5 9 1 52709
0 945 7 1 2 45015 52714
0 946 5 2 1 945
0 947 7 1 2 42646 49864
0 948 7 2 2 52723 947
0 949 5 1 1 52725
0 950 7 6 2 47162 48347
0 951 5 1 1 52727
0 952 7 2 2 42957 52728
0 953 5 1 1 52733
0 954 7 1 2 48509 52734
0 955 5 1 1 954
0 956 7 1 2 949 955
0 957 5 1 1 956
0 958 7 1 2 52704 957
0 959 5 1 1 958
0 960 7 1 2 941 959
0 961 5 1 1 960
0 962 7 1 2 49935 961
0 963 5 1 1 962
0 964 7 3 2 46110 52231
0 965 5 1 1 52735
0 966 7 18 2 47163 47342
0 967 5 4 1 52738
0 968 7 3 2 46381 52739
0 969 5 1 1 52760
0 970 7 1 2 965 969
0 971 5 9 1 970
0 972 7 2 2 48348 52763
0 973 5 1 1 52772
0 974 7 1 2 49813 52773
0 975 5 1 1 974
0 976 7 1 2 963 975
0 977 5 1 1 976
0 978 7 1 2 922 977
0 979 5 1 1 978
0 980 7 1 2 904 979
0 981 7 1 2 900 980
0 982 5 1 1 981
0 983 7 1 2 47839 982
0 984 5 1 1 983
0 985 7 21 2 42112 43496
0 986 5 3 1 52774
0 987 7 3 2 48054 48928
0 988 7 9 2 44144 45148
0 989 5 2 1 52801
0 990 7 4 2 43201 52802
0 991 5 4 1 52812
0 992 7 2 2 48510 50040
0 993 5 2 1 52820
0 994 7 2 2 52816 52822
0 995 5 2 1 52824
0 996 7 1 2 52208 52826
0 997 5 1 1 996
0 998 7 6 2 43966 45355
0 999 5 3 1 52828
0 1000 7 19 2 45149 48728
0 1001 5 3 1 52837
0 1002 7 3 2 44145 52838
0 1003 5 2 1 52859
0 1004 7 2 2 52834 52862
0 1005 5 1 1 52864
0 1006 7 1 2 47482 52369
0 1007 5 1 1 1006
0 1008 7 1 2 49016 1007
0 1009 7 1 2 52865 1008
0 1010 5 1 1 1009
0 1011 7 1 2 43202 1010
0 1012 5 1 1 1011
0 1013 7 11 2 48349 45356
0 1014 5 2 1 52866
0 1015 7 2 2 45357 49724
0 1016 5 2 1 52879
0 1017 7 1 2 46592 49785
0 1018 7 1 2 52881 1017
0 1019 5 1 1 1018
0 1020 7 1 2 52877 1019
0 1021 7 1 2 1012 1020
0 1022 5 1 1 1021
0 1023 7 1 2 43787 1022
0 1024 5 1 1 1023
0 1025 7 1 2 997 1024
0 1026 5 1 1 1025
0 1027 7 1 2 42647 1026
0 1028 5 1 1 1027
0 1029 7 3 2 51414 577
0 1030 5 24 1 52883
0 1031 7 1 2 49936 52886
0 1032 5 3 1 1031
0 1033 7 11 2 48511 49318
0 1034 5 6 1 52913
0 1035 7 1 2 50041 52914
0 1036 5 1 1 1035
0 1037 7 1 2 52910 1036
0 1038 5 1 1 1037
0 1039 7 1 2 43788 1038
0 1040 5 1 1 1039
0 1041 7 9 2 47164 43967
0 1042 7 6 2 42958 52930
0 1043 5 1 1 52939
0 1044 7 2 2 49606 52940
0 1045 5 1 1 52945
0 1046 7 1 2 43203 52946
0 1047 5 1 1 1046
0 1048 7 1 2 1040 1047
0 1049 5 1 1 1048
0 1050 7 1 2 48350 1049
0 1051 5 1 1 1050
0 1052 7 19 2 43789 43968
0 1053 5 1 1 52947
0 1054 7 7 2 42959 52948
0 1055 5 2 1 52966
0 1056 7 9 2 46382 47165
0 1057 5 2 1 52975
0 1058 7 2 2 42648 52984
0 1059 5 2 1 52986
0 1060 7 5 2 52973 52988
0 1061 5 1 1 52990
0 1062 7 9 2 52756 1061
0 1063 5 1 1 52995
0 1064 7 5 2 48351 50042
0 1065 5 1 1 53004
0 1066 7 4 2 49416 49937
0 1067 5 5 1 53009
0 1068 7 1 2 1065 53013
0 1069 5 1 1 1068
0 1070 7 1 2 52996 1069
0 1071 5 1 1 1070
0 1072 7 1 2 1051 1071
0 1073 7 1 2 1028 1072
0 1074 5 1 1 1073
0 1075 7 1 2 52798 1074
0 1076 5 1 1 1075
0 1077 7 1 2 50902 52011
0 1078 7 1 2 51487 1077
0 1079 5 1 1 1078
0 1080 7 1 2 48180 1079
0 1081 7 1 2 1076 1080
0 1082 5 1 1 1081
0 1083 7 6 2 42649 50586
0 1084 5 17 1 53018
0 1085 7 1 2 49786 53019
0 1086 5 9 1 1085
0 1087 7 2 2 48352 53041
0 1088 5 1 1 53050
0 1089 7 1 2 45016 52088
0 1090 5 1 1 1089
0 1091 7 1 2 1088 1090
0 1092 5 1 1 1091
0 1093 7 1 2 47166 1092
0 1094 5 1 1 1093
0 1095 7 8 2 43790 45017
0 1096 5 5 1 53052
0 1097 7 9 2 46111 48353
0 1098 5 4 1 53065
0 1099 7 1 2 53060 53074
0 1100 5 3 1 1099
0 1101 7 1 2 51074 53078
0 1102 5 1 1 1101
0 1103 7 1 2 1094 1102
0 1104 5 1 1 1103
0 1105 7 1 2 50043 1104
0 1106 5 1 1 1105
0 1107 7 1 2 49376 52232
0 1108 5 1 1 1107
0 1109 7 1 2 52220 52691
0 1110 5 1 1 1109
0 1111 7 1 2 1108 1110
0 1112 5 1 1 1111
0 1113 7 1 2 46112 1112
0 1114 5 1 1 1113
0 1115 7 10 2 46383 43791
0 1116 5 2 1 53081
0 1117 7 6 2 47343 49559
0 1118 5 1 1 53093
0 1119 7 1 2 53082 53094
0 1120 5 1 1 1119
0 1121 7 1 2 46384 50254
0 1122 7 1 2 52258 1121
0 1123 5 1 1 1122
0 1124 7 1 2 49560 49938
0 1125 5 2 1 1124
0 1126 7 1 2 42960 53099
0 1127 5 1 1 1126
0 1128 7 1 2 47167 1127
0 1129 7 1 2 1123 1128
0 1130 5 1 1 1129
0 1131 7 1 2 1120 1130
0 1132 7 1 2 1114 1131
0 1133 7 1 2 1106 1132
0 1134 5 1 1 1133
0 1135 7 1 2 50903 1134
0 1136 5 1 1 1135
0 1137 7 28 2 43792 48354
0 1138 5 20 1 53101
0 1139 7 4 2 49020 49668
0 1140 5 1 1 53149
0 1141 7 3 2 53102 53150
0 1142 7 17 2 42650 43204
0 1143 5 1 1 53156
0 1144 7 6 2 44514 50645
0 1145 7 1 2 53157 53173
0 1146 7 1 2 53153 1145
0 1147 5 1 1 1146
0 1148 7 1 2 44856 1147
0 1149 7 1 2 1136 1148
0 1150 5 1 1 1149
0 1151 7 11 2 45930 43661
0 1152 5 1 1 53179
0 1153 7 19 2 42428 47045
0 1154 5 1 1 53190
0 1155 7 9 2 1152 1154
0 1156 5 81 1 53209
0 1157 7 16 2 45664 46874
0 1158 5 3 1 53299
0 1159 7 1 2 53218 53315
0 1160 7 1 2 1150 1159
0 1161 7 1 2 1082 1160
0 1162 5 1 1 1161
0 1163 7 2 2 47168 48987
0 1164 5 1 1 53318
0 1165 7 1 2 48729 1063
0 1166 5 1 1 1165
0 1167 7 1 2 1164 1166
0 1168 5 1 1 1167
0 1169 7 1 2 49939 1168
0 1170 5 1 1 1169
0 1171 7 2 2 50151 52177
0 1172 5 3 1 53320
0 1173 7 1 2 52829 53321
0 1174 5 1 1 1173
0 1175 7 1 2 1170 1174
0 1176 5 1 1 1175
0 1177 7 1 2 45018 1176
0 1178 5 1 1 1177
0 1179 7 5 2 46385 51988
0 1180 5 3 1 53325
0 1181 7 1 2 53005 53326
0 1182 5 1 1 1181
0 1183 7 1 2 49534 52012
0 1184 5 1 1 1183
0 1185 7 1 2 1182 1184
0 1186 5 1 1 1185
0 1187 7 1 2 49725 1186
0 1188 5 1 1 1187
0 1189 7 10 2 43205 48730
0 1190 5 8 1 53333
0 1191 7 1 2 48355 53343
0 1192 5 1 1 1191
0 1193 7 18 2 46386 43206
0 1194 5 2 1 53351
0 1195 7 1 2 49021 53352
0 1196 5 2 1 1195
0 1197 7 1 2 1192 53371
0 1198 5 1 1 1197
0 1199 7 3 2 43793 50587
0 1200 5 6 1 53373
0 1201 7 2 2 53024 53376
0 1202 5 2 1 53382
0 1203 7 6 2 51989 53383
0 1204 7 1 2 1198 53386
0 1205 5 1 1 1204
0 1206 7 10 2 47169 47483
0 1207 5 1 1 53392
0 1208 7 1 2 53066 53393
0 1209 5 1 1 1208
0 1210 7 1 2 48181 1209
0 1211 7 1 2 1205 1210
0 1212 7 1 2 1188 1211
0 1213 7 1 2 1178 1212
0 1214 5 1 1 1213
0 1215 7 2 2 52291 53129
0 1216 5 2 1 53402
0 1217 7 1 2 49319 53403
0 1218 5 1 1 1217
0 1219 7 6 2 46113 50972
0 1220 5 25 1 53406
0 1221 7 1 2 51787 52673
0 1222 7 1 2 53412 1221
0 1223 5 1 1 1222
0 1224 7 1 2 1218 1223
0 1225 5 1 1 1224
0 1226 7 1 2 48512 51837
0 1227 7 1 2 1225 1226
0 1228 5 1 1 1227
0 1229 7 7 2 46593 48356
0 1230 5 4 1 53437
0 1231 7 1 2 49022 50273
0 1232 5 3 1 1231
0 1233 7 1 2 53444 53448
0 1234 5 2 1 1233
0 1235 7 1 2 42651 53451
0 1236 5 1 1 1235
0 1237 7 3 2 45150 49940
0 1238 5 3 1 53453
0 1239 7 11 2 48357 48731
0 1240 7 1 2 53454 53459
0 1241 5 2 1 1240
0 1242 7 1 2 1236 53470
0 1243 5 1 1 1242
0 1244 7 1 2 50926 1243
0 1245 5 1 1 1244
0 1246 7 1 2 44857 1245
0 1247 7 1 2 1228 1246
0 1248 5 1 1 1247
0 1249 7 1 2 50693 1248
0 1250 7 1 2 1214 1249
0 1251 5 1 1 1250
0 1252 7 1 2 1162 1251
0 1253 5 1 1 1252
0 1254 7 1 2 52775 1253
0 1255 5 1 1 1254
0 1256 7 8 2 43794 48513
0 1257 5 3 1 53472
0 1258 7 1 2 47170 49726
0 1259 5 3 1 1258
0 1260 7 2 2 44146 53483
0 1261 5 1 1 53486
0 1262 7 2 2 53480 53487
0 1263 7 1 2 43207 53488
0 1264 5 2 1 1263
0 1265 7 1 2 43795 51538
0 1266 5 1 1 1265
0 1267 7 1 2 53490 1266
0 1268 5 1 1 1267
0 1269 7 1 2 42961 1268
0 1270 5 1 1 1269
0 1271 7 4 2 46387 49941
0 1272 5 4 1 53492
0 1273 7 2 2 43969 51721
0 1274 5 1 1 53500
0 1275 7 1 2 53496 1274
0 1276 5 1 1 1275
0 1277 7 1 2 53473 1276
0 1278 5 1 1 1277
0 1279 7 1 2 1270 1278
0 1280 5 1 1 1279
0 1281 7 1 2 48358 1280
0 1282 5 1 1 1281
0 1283 7 1 2 52211 52233
0 1284 5 5 1 1283
0 1285 7 2 2 51540 53456
0 1286 5 2 1 53507
0 1287 7 1 2 53502 53509
0 1288 5 1 1 1287
0 1289 7 1 2 50927 51722
0 1290 5 1 1 1289
0 1291 7 1 2 49394 1290
0 1292 5 1 1 1291
0 1293 7 1 2 43796 1292
0 1294 5 1 1 1293
0 1295 7 1 2 1288 1294
0 1296 5 1 1 1295
0 1297 7 1 2 42652 1296
0 1298 5 1 1 1297
0 1299 7 4 2 48359 51723
0 1300 5 2 1 53511
0 1301 7 1 2 52259 53515
0 1302 5 1 1 1301
0 1303 7 1 2 52997 1302
0 1304 5 1 1 1303
0 1305 7 1 2 1298 1304
0 1306 7 1 2 1282 1305
0 1307 5 1 1 1306
0 1308 7 1 2 48182 1307
0 1309 5 1 1 1308
0 1310 7 12 2 42962 43797
0 1311 5 5 1 53517
0 1312 7 3 2 53158 53518
0 1313 7 7 2 44147 48360
0 1314 5 1 1 53537
0 1315 7 7 2 44858 49669
0 1316 7 1 2 53538 53544
0 1317 7 1 2 53534 1316
0 1318 5 1 1 1317
0 1319 7 1 2 1309 1318
0 1320 5 1 1 1319
0 1321 7 4 2 48055 51554
0 1322 7 7 2 42113 46875
0 1323 5 1 1 53555
0 1324 7 4 2 917 1323
0 1325 5 56 1 53562
0 1326 7 2 2 53219 53566
0 1327 7 1 2 53551 53622
0 1328 7 1 2 1320 1327
0 1329 5 1 1 1328
0 1330 7 1 2 1255 1329
0 1331 7 1 2 984 1330
0 1332 7 1 2 704 1331
0 1333 5 1 1 1332
0 1334 7 1 2 48919 1333
0 1335 5 1 1 1334
0 1336 7 13 2 46781 43497
0 1337 7 4 2 42114 53624
0 1338 5 1 1 53637
0 1339 7 20 2 43411 46876
0 1340 7 2 2 45665 53641
0 1341 5 1 1 53661
0 1342 7 1 2 1338 1341
0 1343 5 18 1 1342
0 1344 7 1 2 41958 53663
0 1345 5 1 1 1344
0 1346 7 9 2 42115 43412
0 1347 7 5 2 45506 43498
0 1348 7 3 2 53681 53690
0 1349 5 1 1 53695
0 1350 7 1 2 1345 1349
0 1351 5 17 1 1350
0 1352 7 7 2 46114 49727
0 1353 5 12 1 53715
0 1354 7 1 2 45019 53716
0 1355 5 1 1 1354
0 1356 7 14 2 46388 45358
0 1357 5 12 1 53734
0 1358 7 5 2 48361 50588
0 1359 5 6 1 53760
0 1360 7 1 2 53748 53765
0 1361 7 1 2 1355 1360
0 1362 5 1 1 1361
0 1363 7 7 2 42653 48362
0 1364 5 3 1 53771
0 1365 7 1 2 50589 53778
0 1366 7 1 2 50690 1365
0 1367 5 1 1 1366
0 1368 7 1 2 1362 1367
0 1369 5 1 1 1368
0 1370 7 1 2 44859 1369
0 1371 5 1 1 1370
0 1372 7 5 2 46115 49640
0 1373 5 1 1 53781
0 1374 7 1 2 51473 53782
0 1375 5 1 1 1374
0 1376 7 1 2 1371 1375
0 1377 5 1 1 1376
0 1378 7 1 2 47484 1377
0 1379 5 1 1 1378
0 1380 7 2 2 48183 52275
0 1381 7 3 2 50635 53717
0 1382 5 8 1 53788
0 1383 7 1 2 53786 53789
0 1384 5 1 1 1383
0 1385 7 1 2 1379 1384
0 1386 5 1 1 1385
0 1387 7 1 2 46594 1386
0 1388 5 1 1 1387
0 1389 7 14 2 46116 48184
0 1390 5 1 1 53799
0 1391 7 3 2 47344 51427
0 1392 5 2 1 53813
0 1393 7 2 2 52357 53816
0 1394 5 7 1 53818
0 1395 7 1 2 46389 53820
0 1396 5 1 1 1395
0 1397 7 4 2 49135 50530
0 1398 5 1 1 53827
0 1399 7 1 2 1396 1398
0 1400 5 7 1 1399
0 1401 7 1 2 53800 53831
0 1402 5 1 1 1401
0 1403 7 3 2 50285 53334
0 1404 5 1 1 53838
0 1405 7 2 2 45151 53839
0 1406 5 2 1 53841
0 1407 7 1 2 44860 53842
0 1408 5 1 1 1407
0 1409 7 1 2 1402 1408
0 1410 5 1 1 1409
0 1411 7 1 2 45020 1410
0 1412 5 1 1 1411
0 1413 7 1 2 1388 1412
0 1414 5 1 1 1413
0 1415 7 1 2 53220 1414
0 1416 5 1 1 1415
0 1417 7 18 2 42429 46117
0 1418 5 1 1 53845
0 1419 7 4 2 43662 53846
0 1420 7 1 2 51491 53863
0 1421 5 1 1 1420
0 1422 7 2 2 52370 53413
0 1423 7 2 2 48363 50397
0 1424 7 1 2 49942 53869
0 1425 7 1 2 53867 1424
0 1426 5 1 1 1425
0 1427 7 1 2 1421 1426
0 1428 5 1 1 1427
0 1429 7 1 2 44861 1428
0 1430 5 1 1 1429
0 1431 7 4 2 46118 50590
0 1432 5 2 1 53871
0 1433 7 1 2 48364 53872
0 1434 5 2 1 1433
0 1435 7 2 2 51838 53766
0 1436 7 1 2 53749 53879
0 1437 5 1 1 1436
0 1438 7 1 2 53877 1437
0 1439 5 1 1 1438
0 1440 7 10 2 48185 50398
0 1441 5 2 1 53881
0 1442 7 1 2 50727 53882
0 1443 7 1 2 1439 1442
0 1444 5 1 1 1443
0 1445 7 1 2 1430 1444
0 1446 7 1 2 1416 1445
0 1447 5 1 1 1446
0 1448 7 1 2 47171 1447
0 1449 5 1 1 1448
0 1450 7 3 2 42430 52516
0 1451 5 1 1 53893
0 1452 7 7 2 43663 44862
0 1453 5 1 1 53896
0 1454 7 1 2 52470 1453
0 1455 5 20 1 1454
0 1456 7 4 2 45931 53903
0 1457 5 1 1 53923
0 1458 7 2 2 1451 1457
0 1459 5 13 1 53927
0 1460 7 7 2 47172 45152
0 1461 5 4 1 53942
0 1462 7 2 2 49776 53949
0 1463 5 1 1 53953
0 1464 7 1 2 53067 53954
0 1465 5 1 1 1464
0 1466 7 3 2 46119 53735
0 1467 5 2 1 53955
0 1468 7 13 2 43798 47345
0 1469 7 3 2 49561 53960
0 1470 5 1 1 53973
0 1471 7 1 2 53958 53974
0 1472 5 1 1 1471
0 1473 7 1 2 1465 1472
0 1474 5 1 1 1473
0 1475 7 1 2 53929 1474
0 1476 5 1 1 1475
0 1477 7 1 2 52396 53779
0 1478 5 2 1 1477
0 1479 7 1 2 49320 53976
0 1480 5 1 1 1479
0 1481 7 2 2 48973 52674
0 1482 5 1 1 53978
0 1483 7 1 2 53414 53979
0 1484 5 1 1 1483
0 1485 7 1 2 1480 1484
0 1486 5 1 1 1485
0 1487 7 8 2 45932 44863
0 1488 5 1 1 53980
0 1489 7 19 2 47046 43799
0 1490 5 1 1 53988
0 1491 7 2 2 51839 53989
0 1492 5 1 1 54007
0 1493 7 1 2 53981 54008
0 1494 7 1 2 1486 1493
0 1495 5 1 1 1494
0 1496 7 1 2 1476 1495
0 1497 5 1 1 1496
0 1498 7 1 2 50728 1497
0 1499 5 1 1 1498
0 1500 7 1 2 45021 52998
0 1501 5 3 1 1500
0 1502 7 1 2 48514 54009
0 1503 5 1 1 1502
0 1504 7 13 2 42654 49321
0 1505 5 17 1 54012
0 1506 7 1 2 49476 54025
0 1507 5 1 1 1506
0 1508 7 1 2 43800 1507
0 1509 5 1 1 1508
0 1510 7 3 2 42655 49437
0 1511 5 1 1 54042
0 1512 7 2 2 1509 1511
0 1513 5 2 1 54045
0 1514 7 1 2 45153 54046
0 1515 5 1 1 1514
0 1516 7 18 2 44864 48732
0 1517 7 3 2 49891 50294
0 1518 7 1 2 54049 54067
0 1519 7 1 2 1515 1518
0 1520 7 1 2 1503 1519
0 1521 5 1 1 1520
0 1522 7 1 2 1499 1521
0 1523 7 1 2 1449 1522
0 1524 5 1 1 1523
0 1525 7 1 2 44711 1524
0 1526 5 1 1 1525
0 1527 7 9 2 47173 44865
0 1528 5 1 1 54070
0 1529 7 8 2 45933 48056
0 1530 7 15 2 46120 47047
0 1531 7 3 2 54079 54087
0 1532 5 1 1 54102
0 1533 7 1 2 54071 54103
0 1534 7 1 2 51492 1533
0 1535 5 1 1 1534
0 1536 7 1 2 1526 1535
0 1537 5 1 1 1536
0 1538 7 1 2 50348 1537
0 1539 5 1 1 1538
0 1540 7 5 2 47174 50591
0 1541 5 1 1 54105
0 1542 7 1 2 1463 1541
0 1543 5 1 1 1542
0 1544 7 1 2 46121 1543
0 1545 5 2 1 1544
0 1546 7 6 2 45154 52740
0 1547 7 1 2 53750 54112
0 1548 5 1 1 1547
0 1549 7 1 2 51118 1548
0 1550 7 1 2 54110 1549
0 1551 5 1 1 1550
0 1552 7 1 2 48974 52999
0 1553 5 1 1 1552
0 1554 7 3 2 45155 51990
0 1555 5 3 1 54118
0 1556 7 3 2 45359 51991
0 1557 5 1 1 54124
0 1558 7 1 2 49322 52050
0 1559 7 1 2 1557 1558
0 1560 7 1 2 54121 1559
0 1561 5 1 1 1560
0 1562 7 1 2 51162 1561
0 1563 7 1 2 1553 1562
0 1564 5 1 1 1563
0 1565 7 1 2 48365 50445
0 1566 7 1 2 1564 1565
0 1567 7 1 2 1551 1566
0 1568 5 1 1 1567
0 1569 7 4 2 48733 53221
0 1570 7 1 2 50627 54127
0 1571 5 1 1 1570
0 1572 7 9 2 43664 47346
0 1573 7 2 2 49562 54131
0 1574 5 1 1 54140
0 1575 7 1 2 42431 54141
0 1576 5 1 1 1575
0 1577 7 1 2 1571 1576
0 1578 5 1 1 1577
0 1579 7 1 2 51956 1578
0 1580 5 1 1 1579
0 1581 7 2 2 43665 52569
0 1582 5 4 1 54142
0 1583 7 1 2 49670 53990
0 1584 5 2 1 1583
0 1585 7 1 2 54144 54148
0 1586 5 1 1 1585
0 1587 7 1 2 42432 1586
0 1588 5 1 1 1587
0 1589 7 16 2 43666 43801
0 1590 5 1 1 54150
0 1591 7 3 2 45934 49671
0 1592 7 1 2 54151 54166
0 1593 5 2 1 1592
0 1594 7 1 2 1588 54169
0 1595 5 1 1 1594
0 1596 7 1 2 42656 1595
0 1597 5 1 1 1596
0 1598 7 1 2 51119 53975
0 1599 5 1 1 1598
0 1600 7 1 2 1597 1599
0 1601 5 1 1 1600
0 1602 7 1 2 53751 1601
0 1603 5 1 1 1602
0 1604 7 1 2 1580 1603
0 1605 7 1 2 1568 1604
0 1606 5 1 1 1605
0 1607 7 1 2 50729 1606
0 1608 5 1 1 1607
0 1609 7 6 2 43802 53222
0 1610 7 1 2 49471 54171
0 1611 5 1 1 1610
0 1612 7 2 2 49323 53223
0 1613 7 9 2 42657 52603
0 1614 5 1 1 54179
0 1615 7 2 2 54177 54180
0 1616 5 1 1 54188
0 1617 7 1 2 45156 1616
0 1618 7 1 2 1611 1617
0 1619 5 1 1 1618
0 1620 7 3 2 45935 53103
0 1621 5 2 1 54190
0 1622 7 1 2 53210 54193
0 1623 5 3 1 1622
0 1624 7 3 2 48366 53224
0 1625 5 1 1 54198
0 1626 7 26 2 42658 42963
0 1627 5 13 1 54201
0 1628 7 10 2 43970 54202
0 1629 5 1 1 54240
0 1630 7 1 2 1625 54241
0 1631 7 1 2 54195 1630
0 1632 5 1 1 1631
0 1633 7 3 2 951 53061
0 1634 5 37 1 54250
0 1635 7 5 2 53225 54253
0 1636 5 1 1 54290
0 1637 7 1 2 53415 54291
0 1638 5 1 1 1637
0 1639 7 1 2 48515 1638
0 1640 7 1 2 1632 1639
0 1641 5 1 1 1640
0 1642 7 1 2 52292 1641
0 1643 7 1 2 1619 1642
0 1644 5 1 1 1643
0 1645 7 1 2 48186 1644
0 1646 7 1 2 1608 1645
0 1647 5 1 1 1646
0 1648 7 4 2 48975 50730
0 1649 5 3 1 54295
0 1650 7 16 2 42659 43971
0 1651 5 1 1 54302
0 1652 7 1 2 54296 54303
0 1653 5 1 1 1652
0 1654 7 1 2 53471 1653
0 1655 5 1 1 1654
0 1656 7 1 2 42964 1655
0 1657 5 1 1 1656
0 1658 7 4 2 44148 53159
0 1659 7 1 2 52839 54318
0 1660 5 1 1 1659
0 1661 7 1 2 50731 51840
0 1662 7 1 2 53977 1661
0 1663 5 1 1 1662
0 1664 7 1 2 1660 1663
0 1665 7 1 2 1657 1664
0 1666 5 1 1 1665
0 1667 7 1 2 52228 1666
0 1668 5 1 1 1667
0 1669 7 1 2 52293 54254
0 1670 5 1 1 1669
0 1671 7 9 2 43803 47485
0 1672 7 1 2 53438 54322
0 1673 5 2 1 1672
0 1674 7 1 2 1670 54331
0 1675 5 1 1 1674
0 1676 7 2 2 53416 1675
0 1677 5 1 1 54333
0 1678 7 6 2 46595 54323
0 1679 5 2 1 54335
0 1680 7 1 2 53460 54336
0 1681 5 1 1 1680
0 1682 7 1 2 45157 1681
0 1683 5 1 1 1682
0 1684 7 1 2 54334 1683
0 1685 5 1 1 1684
0 1686 7 3 2 49873 53335
0 1687 5 6 1 54343
0 1688 7 1 2 52726 54344
0 1689 5 1 1 1688
0 1690 7 1 2 1685 1689
0 1691 7 1 2 1668 1690
0 1692 5 1 1 1691
0 1693 7 1 2 43667 1692
0 1694 5 1 1 1693
0 1695 7 2 2 43208 53991
0 1696 5 1 1 54352
0 1697 7 5 2 50286 54304
0 1698 7 4 2 48367 52371
0 1699 7 1 2 54354 54359
0 1700 7 1 2 54353 1699
0 1701 5 2 1 1700
0 1702 7 1 2 1694 54363
0 1703 5 1 1 1702
0 1704 7 1 2 42433 1703
0 1705 5 1 1 1704
0 1706 7 29 2 45936 42660
0 1707 5 1 1 54365
0 1708 7 5 2 42965 54366
0 1709 7 1 2 51359 54394
0 1710 7 1 2 53154 1709
0 1711 5 1 1 1710
0 1712 7 1 2 44866 1711
0 1713 7 1 2 1705 1712
0 1714 5 1 1 1713
0 1715 7 1 2 48057 1714
0 1716 7 1 2 1647 1715
0 1717 5 1 1 1716
0 1718 7 4 2 42434 54203
0 1719 7 1 2 43209 54152
0 1720 7 1 2 54399 1719
0 1721 7 3 2 52560 53461
0 1722 7 3 2 43972 51642
0 1723 7 1 2 54403 54406
0 1724 7 1 2 1720 1723
0 1725 5 1 1 1724
0 1726 7 1 2 1717 1725
0 1727 5 1 1 1726
0 1728 7 1 2 48929 1727
0 1729 5 1 1 1728
0 1730 7 1 2 1539 1729
0 1731 5 1 1 1730
0 1732 7 1 2 53698 1731
0 1733 5 1 1 1732
0 1734 7 9 2 43413 47048
0 1735 7 12 2 44515 44712
0 1736 5 1 1 54418
0 1737 7 7 2 44609 44867
0 1738 7 8 2 54419 54430
0 1739 7 1 2 54409 54437
0 1740 5 2 1 1739
0 1741 7 7 2 46782 47840
0 1742 7 3 2 50713 54447
0 1743 7 1 2 52130 54454
0 1744 5 1 1 1743
0 1745 7 1 2 54445 1744
0 1746 5 1 1 1745
0 1747 7 1 2 42435 1746
0 1748 5 1 1 1747
0 1749 7 10 2 43414 44516
0 1750 7 4 2 50489 54457
0 1751 7 1 2 53924 54467
0 1752 5 2 1 1751
0 1753 7 1 2 1748 54471
0 1754 5 1 1 1753
0 1755 7 2 2 41959 1754
0 1756 5 1 1 54473
0 1757 7 1 2 54446 54472
0 1758 5 1 1 1757
0 1759 7 1 2 54474 1758
0 1760 5 1 1 1759
0 1761 7 1 2 43973 1760
0 1762 5 1 1 1761
0 1763 7 11 2 45507 43415
0 1764 5 1 1 54475
0 1765 7 3 2 51555 54476
0 1766 7 2 2 48734 54486
0 1767 7 1 2 48187 51545
0 1768 7 1 2 54489 1767
0 1769 5 1 1 1768
0 1770 7 1 2 1756 1769
0 1771 5 2 1 1770
0 1772 7 1 2 46390 54491
0 1773 7 1 2 1762 1772
0 1774 5 1 1 1773
0 1775 7 19 2 44517 44610
0 1776 7 7 2 44713 54493
0 1777 7 2 2 48886 54512
0 1778 7 1 2 47347 54519
0 1779 7 1 2 53930 1778
0 1780 5 1 1 1779
0 1781 7 1 2 1774 1780
0 1782 5 1 1 1781
0 1783 7 1 2 53130 1782
0 1784 5 1 1 1783
0 1785 7 1 2 52570 54492
0 1786 5 1 1 1785
0 1787 7 1 2 1784 1786
0 1788 5 1 1 1787
0 1789 7 1 2 46122 1788
0 1790 5 1 1 1789
0 1791 7 5 2 48368 52151
0 1792 5 1 1 54521
0 1793 7 12 2 42661 43668
0 1794 5 1 1 54526
0 1795 7 3 2 49582 54527
0 1796 7 3 2 52949 54538
0 1797 7 1 2 54522 54541
0 1798 5 1 1 1797
0 1799 7 5 2 42662 53104
0 1800 5 2 1 54544
0 1801 7 1 2 53931 54545
0 1802 5 1 1 1801
0 1803 7 5 2 45937 52131
0 1804 5 1 1 54551
0 1805 7 3 2 42436 53904
0 1806 5 1 1 54556
0 1807 7 1 2 1804 1806
0 1808 5 10 1 1807
0 1809 7 8 2 46123 52571
0 1810 5 2 1 54569
0 1811 7 1 2 53131 54577
0 1812 7 1 2 54559 1811
0 1813 5 1 1 1812
0 1814 7 1 2 1802 1813
0 1815 5 1 1 1814
0 1816 7 1 2 50928 1815
0 1817 5 1 1 1816
0 1818 7 2 2 49641 51957
0 1819 5 1 1 54579
0 1820 7 1 2 53180 54580
0 1821 5 1 1 1820
0 1822 7 1 2 42663 53053
0 1823 7 1 2 54557 1822
0 1824 5 1 1 1823
0 1825 7 1 2 1821 1824
0 1826 7 1 2 1817 1825
0 1827 5 1 1 1826
0 1828 7 1 2 48058 1827
0 1829 5 1 1 1828
0 1830 7 1 2 1798 1829
0 1831 5 1 1 1830
0 1832 7 1 2 54490 1831
0 1833 5 1 1 1832
0 1834 7 2 2 48369 52659
0 1835 5 1 1 54581
0 1836 7 1 2 53529 54582
0 1837 5 1 1 1836
0 1838 7 1 2 54010 1837
0 1839 5 3 1 1838
0 1840 7 1 2 44868 54583
0 1841 5 1 1 1840
0 1842 7 4 2 47175 49642
0 1843 5 5 1 54586
0 1844 7 1 2 46391 54587
0 1845 5 1 1 1844
0 1846 7 1 2 1841 1845
0 1847 5 1 1 1846
0 1848 7 1 2 47049 1847
0 1849 5 1 1 1848
0 1850 7 9 2 47176 52445
0 1851 7 1 2 51095 54595
0 1852 5 1 1 1851
0 1853 7 1 2 1849 1852
0 1854 5 1 1 1853
0 1855 7 1 2 54468 1854
0 1856 5 1 1 1855
0 1857 7 1 2 48188 54255
0 1858 5 1 1 1857
0 1859 7 3 2 43804 52473
0 1860 5 3 1 54604
0 1861 7 1 2 49664 54607
0 1862 5 7 1 1861
0 1863 7 1 2 42664 54610
0 1864 5 1 1 1863
0 1865 7 1 2 1858 1864
0 1866 5 1 1 1865
0 1867 7 1 2 50929 1866
0 1868 5 1 1 1867
0 1869 7 1 2 1819 1868
0 1870 5 1 1 1869
0 1871 7 1 2 43669 1870
0 1872 5 1 1 1871
0 1873 7 11 2 43805 48189
0 1874 7 1 2 52496 54617
0 1875 7 1 2 54043 1874
0 1876 5 1 1 1875
0 1877 7 1 2 1872 1876
0 1878 5 1 1 1877
0 1879 7 1 2 54455 1878
0 1880 5 1 1 1879
0 1881 7 1 2 45938 1880
0 1882 7 1 2 1856 1881
0 1883 5 1 1 1882
0 1884 7 2 2 43974 49472
0 1885 7 1 2 47177 54628
0 1886 5 1 1 1885
0 1887 7 1 2 54011 1886
0 1888 5 1 1 1887
0 1889 7 1 2 53905 1888
0 1890 5 1 1 1889
0 1891 7 3 2 42665 52474
0 1892 5 1 1 54630
0 1893 7 2 2 52497 52950
0 1894 7 1 2 54631 54633
0 1895 5 1 1 1894
0 1896 7 1 2 1890 1895
0 1897 5 1 1 1896
0 1898 7 1 2 54456 1897
0 1899 5 1 1 1898
0 1900 7 4 2 48190 53462
0 1901 7 2 2 54204 54635
0 1902 7 7 2 43975 47936
0 1903 5 1 1 54641
0 1904 7 2 2 47841 54642
0 1905 7 3 2 46783 54153
0 1906 7 1 2 54648 54650
0 1907 7 1 2 54639 1906
0 1908 5 1 1 1907
0 1909 7 7 2 47050 44518
0 1910 7 3 2 44869 54653
0 1911 7 5 2 43416 44611
0 1912 5 1 1 54663
0 1913 7 1 2 52695 54664
0 1914 7 1 2 54660 1913
0 1915 5 1 1 1914
0 1916 7 1 2 1908 1915
0 1917 5 1 1 1916
0 1918 7 1 2 44714 1917
0 1919 5 1 1 1918
0 1920 7 1 2 42437 1919
0 1921 7 1 2 1899 1920
0 1922 5 1 1 1921
0 1923 7 1 2 41960 1922
0 1924 7 1 2 1883 1923
0 1925 5 1 1 1924
0 1926 7 1 2 1833 1925
0 1927 7 1 2 1790 1926
0 1928 5 1 1 1927
0 1929 7 1 2 48516 1928
0 1930 5 1 1 1929
0 1931 7 1 2 1492 54145
0 1932 5 1 1 1931
0 1933 7 1 2 45939 1932
0 1934 5 1 1 1933
0 1935 7 2 2 52572 53191
0 1936 5 2 1 54668
0 1937 7 1 2 1934 54670
0 1938 5 2 1 1937
0 1939 7 1 2 42966 54672
0 1940 5 1 1 1939
0 1941 7 7 2 43976 52604
0 1942 5 2 1 54674
0 1943 7 3 2 54367 54675
0 1944 5 1 1 54683
0 1945 7 1 2 47051 54684
0 1946 5 1 1 1945
0 1947 7 1 2 1940 1946
0 1948 5 1 1 1947
0 1949 7 3 2 45158 48887
0 1950 7 1 2 54438 54686
0 1951 7 1 2 1948 1950
0 1952 5 1 1 1951
0 1953 7 2 2 43977 45022
0 1954 7 1 2 43806 54689
0 1955 5 2 1 1954
0 1956 7 1 2 42967 54256
0 1957 5 1 1 1956
0 1958 7 1 2 54691 1957
0 1959 5 1 1 1958
0 1960 7 1 2 42666 1959
0 1961 5 1 1 1960
0 1962 7 10 2 47348 48370
0 1963 7 4 2 43807 54693
0 1964 5 1 1 54703
0 1965 7 1 2 51391 54704
0 1966 5 1 1 1965
0 1967 7 1 2 1961 1966
0 1968 5 1 1 1967
0 1969 7 1 2 54560 1968
0 1970 5 1 1 1969
0 1971 7 2 2 42968 50531
0 1972 5 2 1 54707
0 1973 7 7 2 46124 43978
0 1974 5 2 1 54711
0 1975 7 1 2 54709 54718
0 1976 5 1 1 1975
0 1977 7 11 2 47178 48191
0 1978 7 6 2 45023 54720
0 1979 5 2 1 54731
0 1980 7 1 2 51120 54732
0 1981 7 1 2 1976 1980
0 1982 5 1 1 1981
0 1983 7 1 2 1970 1982
0 1984 5 1 1 1983
0 1985 7 10 2 41961 46784
0 1986 5 1 1 54739
0 1987 7 2 2 1764 1986
0 1988 5 66 1 54749
0 1989 7 3 2 48735 54751
0 1990 7 1 2 53552 54817
0 1991 7 1 2 1984 1990
0 1992 5 1 1 1991
0 1993 7 1 2 1952 1992
0 1994 7 1 2 1930 1993
0 1995 5 1 1 1994
0 1996 7 1 2 44149 1995
0 1997 5 1 1 1996
0 1998 7 1 2 49804 53083
0 1999 5 1 1 1998
0 2000 7 1 2 973 1999
0 2001 5 2 1 2000
0 2002 7 1 2 48192 54820
0 2003 5 1 1 2002
0 2004 7 14 2 42667 44870
0 2005 7 1 2 52974 1835
0 2006 5 1 1 2005
0 2007 7 1 2 54822 2006
0 2008 5 1 1 2007
0 2009 7 1 2 2003 2008
0 2010 5 1 1 2009
0 2011 7 1 2 43670 2010
0 2012 5 1 1 2011
0 2013 7 20 2 42668 47052
0 2014 5 1 1 54836
0 2015 7 3 2 48193 54837
0 2016 7 1 2 52685 54856
0 2017 5 1 1 2016
0 2018 7 1 2 2012 2017
0 2019 5 1 1 2018
0 2020 7 1 2 45159 2019
0 2021 5 1 1 2020
0 2022 7 5 2 46392 49672
0 2023 5 5 1 54859
0 2024 7 1 2 54608 54590
0 2025 5 8 1 2024
0 2026 7 1 2 43671 54869
0 2027 5 1 1 2026
0 2028 7 4 2 47053 53105
0 2029 5 3 1 54877
0 2030 7 1 2 48194 54878
0 2031 5 1 1 2030
0 2032 7 1 2 2027 2031
0 2033 5 1 1 2032
0 2034 7 1 2 54860 2033
0 2035 5 1 1 2034
0 2036 7 1 2 2021 2035
0 2037 5 1 1 2036
0 2038 7 1 2 42438 2037
0 2039 5 1 1 2038
0 2040 7 2 2 48371 53084
0 2041 5 1 1 54884
0 2042 7 1 2 49673 54885
0 2043 5 4 1 2042
0 2044 7 13 2 42669 45160
0 2045 5 7 1 54890
0 2046 7 1 2 52686 54891
0 2047 5 1 1 2046
0 2048 7 1 2 54886 2047
0 2049 5 1 1 2048
0 2050 7 1 2 54552 2049
0 2051 5 1 1 2050
0 2052 7 1 2 2039 2051
0 2053 5 1 1 2052
0 2054 7 1 2 45360 2053
0 2055 5 1 1 2054
0 2056 7 1 2 51958 53906
0 2057 5 1 1 2056
0 2058 7 9 2 48195 52013
0 2059 5 1 1 54910
0 2060 7 1 2 43672 54911
0 2061 5 1 1 2060
0 2062 7 1 2 2057 2061
0 2063 5 4 1 2062
0 2064 7 1 2 47349 54919
0 2065 5 1 1 2064
0 2066 7 19 2 43673 47179
0 2067 7 40 2 46125 46393
0 2068 5 9 1 54942
0 2069 7 3 2 54923 54943
0 2070 7 2 2 48196 54991
0 2071 5 1 1 54994
0 2072 7 1 2 2065 2071
0 2073 5 1 1 2072
0 2074 7 1 2 48372 2073
0 2075 5 1 1 2074
0 2076 7 2 2 51831 54618
0 2077 7 1 2 51096 54996
0 2078 5 1 1 2077
0 2079 7 1 2 2075 2078
0 2080 5 1 1 2079
0 2081 7 1 2 42439 2080
0 2082 5 1 1 2081
0 2083 7 9 2 42670 47350
0 2084 5 3 1 54998
0 2085 7 1 2 52132 54999
0 2086 7 1 2 54191 2085
0 2087 5 1 1 2086
0 2088 7 1 2 2082 2087
0 2089 7 1 2 2055 2088
0 2090 5 1 1 2089
0 2091 7 4 2 47842 54752
0 2092 7 1 2 50646 52397
0 2093 7 1 2 55010 2092
0 2094 7 1 2 2090 2093
0 2095 5 1 1 2094
0 2096 7 1 2 1997 2095
0 2097 5 1 1 2096
0 2098 7 1 2 43210 2097
0 2099 5 1 1 2098
0 2100 7 6 2 45940 48373
0 2101 5 1 1 55014
0 2102 7 6 2 42440 52573
0 2103 5 3 1 55020
0 2104 7 1 2 2101 55026
0 2105 5 3 1 2104
0 2106 7 1 2 46126 55029
0 2107 5 1 1 2106
0 2108 7 1 2 45941 54257
0 2109 5 1 1 2108
0 2110 7 1 2 2107 2109
0 2111 5 1 1 2110
0 2112 7 1 2 49260 2111
0 2113 5 1 1 2112
0 2114 7 8 2 45942 47180
0 2115 5 1 1 55032
0 2116 7 1 2 53068 55033
0 2117 5 1 1 2116
0 2118 7 1 2 2113 2117
0 2119 5 1 1 2118
0 2120 7 1 2 53907 2119
0 2121 5 1 1 2120
0 2122 7 1 2 53894 54821
0 2123 5 1 1 2122
0 2124 7 1 2 49805 54995
0 2125 5 1 1 2124
0 2126 7 5 2 43808 54838
0 2127 7 1 2 52475 55040
0 2128 5 1 1 2127
0 2129 7 1 2 2125 2128
0 2130 5 1 1 2129
0 2131 7 1 2 45943 2130
0 2132 5 1 1 2131
0 2133 7 1 2 2123 2132
0 2134 7 1 2 2121 2133
0 2135 5 1 1 2134
0 2136 7 1 2 45161 2135
0 2137 5 1 1 2136
0 2138 7 1 2 836 54146
0 2139 5 3 1 2138
0 2140 7 1 2 46127 55045
0 2141 5 1 1 2140
0 2142 7 2 2 47054 54258
0 2143 5 2 1 55048
0 2144 7 1 2 2141 55050
0 2145 5 1 1 2144
0 2146 7 1 2 45944 2145
0 2147 5 1 1 2146
0 2148 7 1 2 53192 54570
0 2149 5 1 1 2148
0 2150 7 1 2 2147 2149
0 2151 5 1 1 2150
0 2152 7 1 2 51075 2151
0 2153 5 1 1 2152
0 2154 7 5 2 50399 52014
0 2155 7 1 2 48374 55052
0 2156 5 1 1 2155
0 2157 7 1 2 48197 2156
0 2158 7 1 2 2153 2157
0 2159 5 1 1 2158
0 2160 7 4 2 42671 53992
0 2161 5 2 1 55057
0 2162 7 10 2 46128 54924
0 2163 5 3 1 55063
0 2164 7 1 2 55061 55073
0 2165 5 6 1 2164
0 2166 7 2 2 45945 55076
0 2167 5 1 1 55082
0 2168 7 3 2 52015 53193
0 2169 5 1 1 55084
0 2170 7 1 2 2167 2169
0 2171 5 3 1 2170
0 2172 7 1 2 48375 55087
0 2173 5 1 1 2172
0 2174 7 1 2 44871 2173
0 2175 7 1 2 52089 54673
0 2176 5 1 1 2175
0 2177 7 1 2 727 53062
0 2178 5 2 1 2177
0 2179 7 1 2 53226 55090
0 2180 5 1 1 2179
0 2181 7 18 2 46129 43674
0 2182 5 1 1 55092
0 2183 7 4 2 52574 55093
0 2184 5 1 1 55110
0 2185 7 2 2 42441 55111
0 2186 5 2 1 55114
0 2187 7 1 2 2180 55116
0 2188 5 1 1 2187
0 2189 7 1 2 51076 2188
0 2190 5 1 1 2189
0 2191 7 1 2 2176 2190
0 2192 7 1 2 2174 2191
0 2193 5 1 1 2192
0 2194 7 1 2 51217 2193
0 2195 7 1 2 2159 2194
0 2196 5 1 1 2195
0 2197 7 1 2 2137 2196
0 2198 5 1 1 2197
0 2199 7 1 2 54520 2198
0 2200 5 1 1 2199
0 2201 7 4 2 47937 54448
0 2202 7 3 2 48736 52605
0 2203 5 1 1 55122
0 2204 7 7 2 42672 50930
0 2205 5 3 1 55125
0 2206 7 1 2 55123 55126
0 2207 7 1 2 54561 2206
0 2208 5 1 1 2207
0 2209 7 1 2 48198 52867
0 2210 7 8 2 43675 47486
0 2211 7 11 2 42442 46394
0 2212 7 10 2 46130 43809
0 2213 5 5 1 55154
0 2214 7 1 2 55143 55155
0 2215 7 1 2 55135 2214
0 2216 7 1 2 2209 2215
0 2217 5 1 1 2216
0 2218 7 1 2 2208 2217
0 2219 5 1 1 2218
0 2220 7 1 2 55118 2219
0 2221 5 1 1 2220
0 2222 7 4 2 47181 44612
0 2223 7 2 2 52517 55169
0 2224 7 2 2 43417 55173
0 2225 7 2 2 44519 49065
0 2226 7 16 2 45946 46131
0 2227 7 1 2 55177 55179
0 2228 7 1 2 55175 2227
0 2229 5 1 1 2228
0 2230 7 9 2 46395 48737
0 2231 5 2 1 55195
0 2232 7 3 2 45361 54982
0 2233 5 1 1 55206
0 2234 7 1 2 47487 55207
0 2235 5 1 1 2234
0 2236 7 1 2 55204 2235
0 2237 5 2 1 2236
0 2238 7 2 2 51121 54449
0 2239 7 12 2 47938 48199
0 2240 7 1 2 43810 55213
0 2241 7 1 2 55211 2240
0 2242 7 1 2 55209 2241
0 2243 5 1 1 2242
0 2244 7 1 2 2229 2243
0 2245 5 1 1 2244
0 2246 7 1 2 45024 2245
0 2247 5 1 1 2246
0 2248 7 10 2 42969 47182
0 2249 5 1 1 55225
0 2250 7 1 2 49136 55226
0 2251 5 1 1 2250
0 2252 7 2 2 51992 55196
0 2253 5 1 1 55235
0 2254 7 1 2 2251 2253
0 2255 5 1 1 2254
0 2256 7 4 2 47939 51263
0 2257 7 1 2 55212 55237
0 2258 7 1 2 2255 2257
0 2259 5 1 1 2258
0 2260 7 1 2 2247 2259
0 2261 5 1 1 2260
0 2262 7 1 2 47351 2261
0 2263 5 1 1 2262
0 2264 7 1 2 2221 2263
0 2265 5 1 1 2264
0 2266 7 1 2 45162 2265
0 2267 5 1 1 2266
0 2268 7 2 2 42970 50319
0 2269 5 1 1 55241
0 2270 7 1 2 53767 2269
0 2271 5 1 1 2270
0 2272 7 1 2 42673 2271
0 2273 5 1 1 2272
0 2274 7 1 2 42971 49447
0 2275 5 1 1 2274
0 2276 7 1 2 2273 2275
0 2277 5 1 1 2276
0 2278 7 1 2 49137 2277
0 2279 5 1 1 2278
0 2280 7 2 2 49480 51495
0 2281 7 1 2 48376 55243
0 2282 5 1 1 2281
0 2283 7 1 2 2279 2282
0 2284 5 1 1 2283
0 2285 7 2 2 43811 2284
0 2286 5 1 1 55245
0 2287 7 6 2 47488 52868
0 2288 5 3 1 55247
0 2289 7 4 2 52710 54305
0 2290 5 1 1 55256
0 2291 7 1 2 55248 55257
0 2292 5 1 1 2291
0 2293 7 1 2 51163 2292
0 2294 7 1 2 2286 2293
0 2295 5 1 1 2294
0 2296 7 6 2 48200 50446
0 2297 5 1 1 55260
0 2298 7 5 2 42674 45025
0 2299 5 1 1 55266
0 2300 7 1 2 42972 55267
0 2301 5 1 1 2300
0 2302 7 1 2 53878 2301
0 2303 5 1 1 2302
0 2304 7 1 2 49138 2303
0 2305 5 1 1 2304
0 2306 7 1 2 53780 55197
0 2307 7 1 2 50320 2306
0 2308 5 1 1 2307
0 2309 7 1 2 2305 2308
0 2310 5 1 1 2309
0 2311 7 1 2 47183 2310
0 2312 5 1 1 2311
0 2313 7 1 2 43812 49417
0 2314 5 3 1 2313
0 2315 7 6 2 47352 49139
0 2316 5 3 1 55274
0 2317 7 1 2 49851 55275
0 2318 5 1 1 2317
0 2319 7 1 2 55271 2318
0 2320 5 1 1 2319
0 2321 7 1 2 54944 2320
0 2322 5 1 1 2321
0 2323 7 1 2 51122 2322
0 2324 7 1 2 2312 2323
0 2325 5 1 1 2324
0 2326 7 1 2 55261 2325
0 2327 7 1 2 2295 2326
0 2328 5 1 1 2327
0 2329 7 9 2 44872 51123
0 2330 5 1 1 55283
0 2331 7 1 2 55246 55284
0 2332 5 1 1 2331
0 2333 7 1 2 2328 2332
0 2334 5 1 1 2333
0 2335 7 1 2 55119 2334
0 2336 5 1 1 2335
0 2337 7 1 2 2267 2336
0 2338 5 1 1 2337
0 2339 7 1 2 41962 2338
0 2340 5 1 1 2339
0 2341 7 2 2 47489 48988
0 2342 5 5 1 55292
0 2343 7 2 2 52856 55294
0 2344 5 4 1 55299
0 2345 7 2 2 43979 55301
0 2346 5 1 1 55305
0 2347 7 1 2 55253 2346
0 2348 5 1 1 2347
0 2349 7 1 2 43813 2348
0 2350 5 1 1 2349
0 2351 7 2 2 49438 52840
0 2352 5 1 1 55307
0 2353 7 1 2 2350 2352
0 2354 5 1 1 2353
0 2355 7 1 2 42973 2354
0 2356 5 1 1 2355
0 2357 7 3 2 52869 54324
0 2358 5 1 1 55309
0 2359 7 1 2 50592 55310
0 2360 5 1 1 2359
0 2361 7 1 2 2356 2360
0 2362 5 1 1 2361
0 2363 7 1 2 42675 2362
0 2364 5 1 1 2363
0 2365 7 7 2 42974 49187
0 2366 5 11 1 55312
0 2367 7 1 2 49674 53106
0 2368 7 1 2 53752 2367
0 2369 7 1 2 55319 2368
0 2370 5 2 1 2369
0 2371 7 1 2 2364 55330
0 2372 5 1 1 2371
0 2373 7 1 2 55285 2372
0 2374 5 1 1 2373
0 2375 7 3 2 42975 53943
0 2376 5 1 1 55332
0 2377 7 1 2 47353 55333
0 2378 5 1 1 2377
0 2379 7 1 2 48377 2378
0 2380 7 1 2 54111 2379
0 2381 5 1 1 2380
0 2382 7 1 2 52987 53377
0 2383 5 2 1 2382
0 2384 7 1 2 51392 53961
0 2385 5 1 1 2384
0 2386 7 1 2 45026 2385
0 2387 7 1 2 55335 2386
0 2388 5 1 1 2387
0 2389 7 1 2 49140 2388
0 2390 7 1 2 2381 2389
0 2391 5 1 1 2390
0 2392 7 1 2 53025 54259
0 2393 5 1 1 2392
0 2394 7 9 2 46132 47354
0 2395 7 3 2 48378 55337
0 2396 5 1 1 55346
0 2397 7 2 2 48517 52931
0 2398 5 2 1 55349
0 2399 7 1 2 2396 55351
0 2400 5 1 1 2399
0 2401 7 3 2 49865 2400
0 2402 5 1 1 55353
0 2403 7 1 2 2393 2402
0 2404 5 2 1 2403
0 2405 7 1 2 55198 55356
0 2406 5 1 1 2405
0 2407 7 1 2 2391 2406
0 2408 5 1 1 2407
0 2409 7 1 2 42443 2408
0 2410 5 1 1 2409
0 2411 7 1 2 53211 2410
0 2412 5 1 1 2411
0 2413 7 4 2 45163 49261
0 2414 5 3 1 55358
0 2415 7 2 2 43814 55362
0 2416 5 2 1 55365
0 2417 7 1 2 55249 55366
0 2418 5 1 1 2417
0 2419 7 1 2 50931 52606
0 2420 7 1 2 55302 2419
0 2421 5 1 1 2420
0 2422 7 1 2 2418 2421
0 2423 5 1 1 2422
0 2424 7 1 2 42676 2423
0 2425 5 1 1 2424
0 2426 7 1 2 51164 55331
0 2427 7 1 2 2425 2426
0 2428 5 1 1 2427
0 2429 7 1 2 48201 2428
0 2430 7 1 2 2412 2429
0 2431 5 1 1 2430
0 2432 7 1 2 2374 2431
0 2433 5 1 1 2432
0 2434 7 1 2 54487 2433
0 2435 5 1 1 2434
0 2436 7 1 2 2340 2435
0 2437 5 1 1 2436
0 2438 7 1 2 46596 2437
0 2439 5 1 1 2438
0 2440 7 21 2 42677 46597
0 2441 7 1 2 51556 55369
0 2442 7 1 2 54636 2441
0 2443 7 1 2 54651 2442
0 2444 5 1 1 2443
0 2445 7 3 2 45027 51218
0 2446 7 2 2 44520 54945
0 2447 7 1 2 55176 55393
0 2448 7 1 2 55390 2447
0 2449 5 1 1 2448
0 2450 7 1 2 2444 2449
0 2451 5 1 1 2450
0 2452 7 1 2 45947 2451
0 2453 5 1 1 2452
0 2454 7 9 2 42444 46785
0 2455 7 2 2 48738 55395
0 2456 7 1 2 51557 53439
0 2457 7 1 2 55404 2456
0 2458 7 1 2 54920 2457
0 2459 5 1 1 2458
0 2460 7 1 2 2453 2459
0 2461 5 1 1 2460
0 2462 7 1 2 41963 2461
0 2463 5 1 1 2462
0 2464 7 1 2 42445 54921
0 2465 5 1 1 2464
0 2466 7 1 2 51959 54553
0 2467 5 1 1 2466
0 2468 7 1 2 2465 2467
0 2469 5 1 1 2468
0 2470 7 8 2 46598 43418
0 2471 7 2 2 45508 55406
0 2472 7 15 2 47843 48739
0 2473 7 4 2 47940 48379
0 2474 7 1 2 55416 55431
0 2475 7 1 2 55414 2474
0 2476 7 1 2 2469 2475
0 2477 5 1 1 2476
0 2478 7 1 2 2463 2477
0 2479 5 1 1 2478
0 2480 7 1 2 49728 2479
0 2481 5 1 1 2480
0 2482 7 5 2 43419 47355
0 2483 7 7 2 44613 45164
0 2484 7 3 2 44521 55440
0 2485 7 2 2 55435 55447
0 2486 7 1 2 54072 54088
0 2487 7 1 2 55320 2486
0 2488 7 1 2 55450 2487
0 2489 5 1 1 2488
0 2490 7 14 2 42678 46786
0 2491 7 3 2 54154 55452
0 2492 7 11 2 48740 49324
0 2493 5 2 1 55469
0 2494 7 4 2 47844 48202
0 2495 7 10 2 47941 48518
0 2496 7 1 2 55482 55486
0 2497 7 1 2 55470 2496
0 2498 7 1 2 55466 2497
0 2499 5 1 1 2498
0 2500 7 1 2 2489 2499
0 2501 5 1 1 2500
0 2502 7 1 2 45948 2501
0 2503 5 1 1 2502
0 2504 7 7 2 43980 48203
0 2505 7 2 2 55064 55496
0 2506 5 1 1 55503
0 2507 7 4 2 49325 51960
0 2508 5 1 1 55505
0 2509 7 1 2 53908 55506
0 2510 5 1 1 2509
0 2511 7 1 2 2506 2510
0 2512 5 1 1 2511
0 2513 7 1 2 47845 55487
0 2514 7 1 2 55405 2513
0 2515 7 1 2 2512 2514
0 2516 5 1 1 2515
0 2517 7 1 2 2503 2516
0 2518 5 1 1 2517
0 2519 7 1 2 41964 2518
0 2520 5 1 1 2519
0 2521 7 1 2 54562 55507
0 2522 5 1 1 2521
0 2523 7 1 2 42446 55504
0 2524 5 1 1 2523
0 2525 7 1 2 2522 2524
0 2526 5 1 1 2525
0 2527 7 1 2 52372 54488
0 2528 7 1 2 2526 2527
0 2529 5 1 1 2528
0 2530 7 1 2 2520 2529
0 2531 5 1 1 2530
0 2532 7 1 2 45028 2531
0 2533 5 1 1 2532
0 2534 7 2 2 54563 54818
0 2535 7 4 2 47846 48380
0 2536 7 2 2 48519 55511
0 2537 7 12 2 42679 47184
0 2538 5 2 1 55517
0 2539 7 5 2 42976 47942
0 2540 7 1 2 55518 55531
0 2541 7 1 2 55515 2540
0 2542 7 1 2 55509 2541
0 2543 5 1 1 2542
0 2544 7 1 2 2533 2543
0 2545 7 1 2 2481 2544
0 2546 7 1 2 2439 2545
0 2547 5 1 1 2546
0 2548 7 1 2 48059 2547
0 2549 5 1 1 2548
0 2550 7 1 2 2200 2549
0 2551 7 1 2 2099 2550
0 2552 5 1 1 2551
0 2553 7 1 2 53567 2552
0 2554 5 1 1 2553
0 2555 7 1 2 1733 2554
0 2556 5 1 1 2555
0 2557 7 1 2 47702 2556
0 2558 5 1 1 2557
0 2559 7 2 2 46599 44150
0 2560 5 4 1 55536
0 2561 7 4 2 43211 47490
0 2562 5 3 1 55542
0 2563 7 4 2 55538 55546
0 2564 5 44 1 55549
0 2565 7 38 2 46787 47703
0 2566 5 1 1 55597
0 2567 7 1 2 51654 54922
0 2568 5 1 1 2567
0 2569 7 2 2 48204 50668
0 2570 7 6 2 46396 43499
0 2571 7 1 2 54125 55637
0 2572 7 1 2 55635 2571
0 2573 5 1 1 2572
0 2574 7 1 2 2568 2573
0 2575 5 1 1 2574
0 2576 7 1 2 48381 2575
0 2577 5 1 1 2576
0 2578 7 1 2 51580 53085
0 2579 7 6 2 43676 45029
0 2580 5 1 1 55643
0 2581 7 12 2 48205 45362
0 2582 7 1 2 55644 55649
0 2583 7 1 2 2578 2582
0 2584 5 1 1 2583
0 2585 7 1 2 2577 2584
0 2586 5 1 1 2585
0 2587 7 1 2 42447 2586
0 2588 5 1 1 2587
0 2589 7 2 2 54619 55512
0 2590 7 6 2 46877 43677
0 2591 7 1 2 54368 55663
0 2592 7 1 2 55661 2591
0 2593 5 1 1 2592
0 2594 7 1 2 2588 2593
0 2595 5 1 1 2594
0 2596 7 1 2 49729 2595
0 2597 5 1 1 2596
0 2598 7 7 2 43981 47847
0 2599 7 5 2 46397 46878
0 2600 7 2 2 55669 55676
0 2601 5 1 1 55681
0 2602 7 3 2 43815 49852
0 2603 5 2 1 55683
0 2604 7 1 2 47055 55684
0 2605 7 1 2 55682 2604
0 2606 5 1 1 2605
0 2607 7 2 2 47185 49675
0 2608 5 5 1 55688
0 2609 7 1 2 55164 55690
0 2610 5 3 1 2609
0 2611 7 2 2 45030 55695
0 2612 5 1 1 55698
0 2613 7 1 2 48382 53387
0 2614 5 1 1 2613
0 2615 7 2 2 2612 2614
0 2616 5 2 1 55700
0 2617 7 12 2 44522 45363
0 2618 7 5 2 43500 55704
0 2619 5 8 1 55716
0 2620 7 7 2 46398 47848
0 2621 7 2 2 46879 55729
0 2622 5 1 1 55736
0 2623 7 1 2 55721 2622
0 2624 5 3 1 2623
0 2625 7 1 2 43678 55738
0 2626 7 1 2 55702 2625
0 2627 5 1 1 2626
0 2628 7 1 2 2606 2627
0 2629 5 1 1 2628
0 2630 7 1 2 42448 2629
0 2631 5 1 1 2630
0 2632 7 6 2 46880 43816
0 2633 7 1 2 48983 53181
0 2634 7 1 2 55741 2633
0 2635 7 1 2 55516 2634
0 2636 5 1 1 2635
0 2637 7 1 2 2631 2636
0 2638 5 1 1 2637
0 2639 7 1 2 48206 2638
0 2640 5 1 1 2639
0 2641 7 1 2 2597 2640
0 2642 5 1 1 2641
0 2643 7 1 2 55598 2642
0 2644 5 1 1 2643
0 2645 7 23 2 43420 43501
0 2646 5 1 1 55747
0 2647 7 18 2 44374 44523
0 2648 7 3 2 48520 55770
0 2649 7 1 2 55748 55788
0 2650 5 1 1 2649
0 2651 7 16 2 46788 46881
0 2652 7 3 2 42977 55791
0 2653 7 16 2 47849 45165
0 2654 7 7 2 43982 47704
0 2655 7 1 2 55810 55826
0 2656 7 3 2 55807 2655
0 2657 5 1 1 55833
0 2658 7 1 2 2650 2657
0 2659 5 1 1 2658
0 2660 7 1 2 42680 2659
0 2661 5 1 1 2660
0 2662 7 2 2 44524 49676
0 2663 7 16 2 43502 44375
0 2664 7 12 2 42978 43421
0 2665 7 1 2 55838 55854
0 2666 7 1 2 55836 2665
0 2667 5 1 1 2666
0 2668 7 1 2 2661 2667
0 2669 5 1 1 2668
0 2670 7 1 2 53897 2669
0 2671 5 1 1 2670
0 2672 7 1 2 54857 55834
0 2673 5 1 1 2672
0 2674 7 1 2 2671 2673
0 2675 5 1 1 2674
0 2676 7 1 2 42449 2675
0 2677 5 1 1 2676
0 2678 7 5 2 43679 54369
0 2679 7 1 2 48207 55866
0 2680 7 1 2 55835 2679
0 2681 5 1 1 2680
0 2682 7 1 2 2677 2681
0 2683 5 1 1 2682
0 2684 7 1 2 52607 2683
0 2685 5 1 1 2684
0 2686 7 53 2 43422 44376
0 2687 5 7 1 55871
0 2688 7 3 2 51581 55872
0 2689 7 1 2 181 49665
0 2690 5 1 1 2689
0 2691 7 1 2 50447 51418
0 2692 7 1 2 2690 2691
0 2693 5 1 1 2692
0 2694 7 1 2 2330 2693
0 2695 5 1 1 2694
0 2696 7 1 2 43983 2695
0 2697 5 1 1 2696
0 2698 7 1 2 42979 54564
0 2699 5 1 1 2698
0 2700 7 1 2 2697 2699
0 2701 5 1 1 2700
0 2702 7 1 2 42681 2701
0 2703 5 1 1 2702
0 2704 7 2 2 51124 51462
0 2705 5 1 1 55934
0 2706 7 1 2 52476 55935
0 2707 5 1 1 2706
0 2708 7 1 2 2703 2707
0 2709 5 1 1 2708
0 2710 7 1 2 43817 2709
0 2711 5 1 1 2710
0 2712 7 2 2 49600 54306
0 2713 5 2 1 55936
0 2714 7 1 2 49418 54721
0 2715 5 2 1 2714
0 2716 7 1 2 55938 55940
0 2717 5 1 1 2716
0 2718 7 1 2 48521 51125
0 2719 7 1 2 2717 2718
0 2720 5 1 1 2719
0 2721 7 1 2 2711 2720
0 2722 5 1 1 2721
0 2723 7 1 2 55931 2722
0 2724 5 1 1 2723
0 2725 7 1 2 2685 2724
0 2726 7 1 2 2644 2725
0 2727 5 1 1 2726
0 2728 7 1 2 50647 2727
0 2729 5 1 1 2728
0 2730 7 1 2 49777 55091
0 2731 5 1 1 2730
0 2732 7 1 2 55701 2731
0 2733 5 2 1 2732
0 2734 7 5 2 45364 50490
0 2735 7 1 2 53932 55944
0 2736 7 2 2 55942 2735
0 2737 7 18 2 43503 47850
0 2738 7 1 2 55599 55951
0 2739 7 1 2 55949 2738
0 2740 5 1 1 2739
0 2741 7 1 2 2729 2740
0 2742 5 1 1 2741
0 2743 7 1 2 42116 2742
0 2744 5 1 1 2743
0 2745 7 8 2 45666 47705
0 2746 7 1 2 53642 55950
0 2747 5 1 1 2746
0 2748 7 1 2 45166 52687
0 2749 5 1 1 2748
0 2750 7 1 2 1964 2749
0 2751 5 1 1 2750
0 2752 7 2 2 42682 2751
0 2753 5 1 1 55977
0 2754 7 1 2 54887 2753
0 2755 5 2 1 2754
0 2756 7 1 2 53182 55979
0 2757 5 1 1 2756
0 2758 7 1 2 52660 54839
0 2759 5 2 1 2758
0 2760 7 1 2 43680 52764
0 2761 5 2 1 2760
0 2762 7 1 2 55981 55983
0 2763 5 1 1 2762
0 2764 7 1 2 45167 2763
0 2765 5 1 1 2764
0 2766 7 1 2 54864 55007
0 2767 5 12 1 2766
0 2768 7 1 2 53993 55985
0 2769 5 1 1 2768
0 2770 7 2 2 2765 2769
0 2771 5 1 1 55997
0 2772 7 1 2 50973 55065
0 2773 5 1 1 2772
0 2774 7 1 2 55998 2773
0 2775 5 1 1 2774
0 2776 7 1 2 48383 2775
0 2777 5 1 1 2776
0 2778 7 4 2 43984 45168
0 2779 7 3 2 42980 55999
0 2780 7 1 2 55058 56003
0 2781 5 1 1 2780
0 2782 7 1 2 51097 55699
0 2783 5 1 1 2782
0 2784 7 1 2 2781 2783
0 2785 7 1 2 2777 2784
0 2786 5 1 1 2785
0 2787 7 1 2 42450 2786
0 2788 5 1 1 2787
0 2789 7 1 2 2757 2788
0 2790 5 1 1 2789
0 2791 7 1 2 48208 2790
0 2792 5 1 1 2791
0 2793 7 2 2 55286 55978
0 2794 5 1 1 56006
0 2795 7 1 2 2792 2794
0 2796 5 1 1 2795
0 2797 7 1 2 50648 53625
0 2798 7 1 2 2796 2797
0 2799 5 1 1 2798
0 2800 7 1 2 2747 2799
0 2801 5 1 1 2800
0 2802 7 1 2 47851 2801
0 2803 5 1 1 2802
0 2804 7 2 2 43423 52144
0 2805 7 14 2 48060 45365
0 2806 7 3 2 47943 56010
0 2807 7 1 2 55636 56024
0 2808 7 2 2 55943 2807
0 2809 7 1 2 56008 56027
0 2810 5 1 1 2809
0 2811 7 1 2 2803 2810
0 2812 5 1 1 2811
0 2813 7 1 2 55969 2812
0 2814 5 1 1 2813
0 2815 7 1 2 2744 2814
0 2816 5 1 1 2815
0 2817 7 1 2 41965 2816
0 2818 5 1 1 2817
0 2819 7 7 2 47706 54477
0 2820 7 8 2 42117 42451
0 2821 7 2 2 43504 56036
0 2822 7 1 2 56028 56044
0 2823 5 1 1 2822
0 2824 7 1 2 46399 52541
0 2825 5 1 1 2824
0 2826 7 2 2 45949 43505
0 2827 7 3 2 47056 56046
0 2828 7 1 2 55945 56048
0 2829 5 1 1 2828
0 2830 7 1 2 2825 2829
0 2831 5 1 1 2830
0 2832 7 1 2 42118 2831
0 2833 5 1 1 2832
0 2834 7 2 2 50649 55144
0 2835 7 3 2 43506 43681
0 2836 7 3 2 45667 56053
0 2837 7 1 2 56051 56056
0 2838 5 1 1 2837
0 2839 7 1 2 2833 2838
0 2840 5 1 1 2839
0 2841 7 1 2 55703 2840
0 2842 5 1 1 2841
0 2843 7 1 2 47186 52542
0 2844 5 1 1 2843
0 2845 7 6 2 43507 47057
0 2846 7 1 2 50910 56059
0 2847 7 2 2 55946 2846
0 2848 5 1 1 56065
0 2849 7 1 2 2844 2848
0 2850 5 1 1 2849
0 2851 7 1 2 42119 2850
0 2852 5 1 1 2851
0 2853 7 1 2 47187 52557
0 2854 5 1 1 2853
0 2855 7 1 2 2852 2854
0 2856 5 1 1 2855
0 2857 7 1 2 46133 2856
0 2858 5 1 1 2857
0 2859 7 4 2 42120 47188
0 2860 7 1 2 56066 56067
0 2861 5 1 1 2860
0 2862 7 1 2 2858 2861
0 2863 5 1 1 2862
0 2864 7 1 2 48384 2863
0 2865 5 1 1 2864
0 2866 7 8 2 42121 45950
0 2867 7 2 2 56060 56071
0 2868 7 3 2 44715 52276
0 2869 7 5 2 43818 44614
0 2870 7 1 2 46400 56084
0 2871 7 1 2 56081 2870
0 2872 7 1 2 56079 2871
0 2873 5 1 1 2872
0 2874 7 1 2 2865 2873
0 2875 5 1 1 2874
0 2876 7 1 2 49730 2875
0 2877 5 1 1 2876
0 2878 7 1 2 2842 2877
0 2879 5 1 1 2878
0 2880 7 1 2 48209 2879
0 2881 5 1 1 2880
0 2882 7 2 2 45366 52765
0 2883 7 1 2 51871 56089
0 2884 5 1 1 2883
0 2885 7 6 2 48061 48210
0 2886 7 3 2 47944 56091
0 2887 7 1 2 55742 56097
0 2888 7 1 2 55986 2887
0 2889 5 1 1 2888
0 2890 7 1 2 2884 2889
0 2891 5 1 1 2890
0 2892 7 1 2 48385 2891
0 2893 5 1 1 2892
0 2894 7 10 2 45367 50974
0 2895 5 1 1 56100
0 2896 7 3 2 51993 56101
0 2897 7 1 2 51872 56110
0 2898 5 1 1 2897
0 2899 7 4 2 48211 50650
0 2900 7 11 2 42683 46882
0 2901 7 1 2 52661 56117
0 2902 7 1 2 56113 2901
0 2903 5 1 1 2902
0 2904 7 1 2 2898 2903
0 2905 5 1 1 2904
0 2906 7 1 2 48386 2905
0 2907 5 1 1 2906
0 2908 7 2 2 51873 52277
0 2909 7 1 2 46401 56128
0 2910 5 1 1 2909
0 2911 7 7 2 42981 46883
0 2912 7 3 2 42684 56130
0 2913 7 6 2 43985 48062
0 2914 7 2 2 55214 56140
0 2915 7 1 2 56137 56146
0 2916 5 1 1 2915
0 2917 7 1 2 2910 2916
0 2918 5 1 1 2917
0 2919 7 1 2 43819 2918
0 2920 5 1 1 2919
0 2921 7 1 2 2907 2920
0 2922 5 1 1 2921
0 2923 7 1 2 45169 2922
0 2924 5 1 1 2923
0 2925 7 3 2 43820 54026
0 2926 5 2 1 56148
0 2927 7 1 2 55691 56151
0 2928 5 1 1 2927
0 2929 7 1 2 56129 2928
0 2930 5 1 1 2929
0 2931 7 1 2 2924 2930
0 2932 7 1 2 2893 2931
0 2933 5 1 1 2932
0 2934 7 1 2 42122 2933
0 2935 5 1 1 2934
0 2936 7 1 2 52551 56114
0 2937 7 1 2 55980 2936
0 2938 5 1 1 2937
0 2939 7 1 2 2935 2938
0 2940 5 1 1 2939
0 2941 7 1 2 53227 2940
0 2942 5 1 1 2941
0 2943 7 3 2 50651 53568
0 2944 7 1 2 56007 56153
0 2945 5 1 1 2944
0 2946 7 1 2 2942 2945
0 2947 7 1 2 2881 2946
0 2948 5 1 1 2947
0 2949 7 1 2 47852 2948
0 2950 5 1 1 2949
0 2951 7 1 2 2823 2950
0 2952 5 1 1 2951
0 2953 7 1 2 56029 2952
0 2954 5 1 1 2953
0 2955 7 8 2 48063 51264
0 2956 7 4 2 48930 56156
0 2957 5 1 1 56164
0 2958 7 1 2 49677 56165
0 2959 5 1 1 2958
0 2960 7 1 2 50384 53095
0 2961 5 1 1 2960
0 2962 7 1 2 2959 2961
0 2963 5 2 1 2962
0 2964 7 2 2 45368 53228
0 2965 7 3 2 47707 53699
0 2966 7 1 2 56170 56172
0 2967 5 1 1 2966
0 2968 7 6 2 41966 42982
0 2969 7 13 2 44377 48741
0 2970 7 3 2 56175 56181
0 2971 5 1 1 56194
0 2972 7 5 2 42123 42685
0 2973 7 3 2 43424 56061
0 2974 7 1 2 56197 56202
0 2975 7 1 2 56195 2974
0 2976 5 1 1 2975
0 2977 7 1 2 2967 2976
0 2978 5 1 1 2977
0 2979 7 1 2 43821 2978
0 2980 5 1 1 2979
0 2981 7 21 2 46134 42983
0 2982 5 1 1 56205
0 2983 7 18 2 41967 42124
0 2984 7 3 2 56206 56226
0 2985 7 8 2 43508 47189
0 2986 7 2 2 55873 56247
0 2987 7 11 2 48742 50448
0 2988 5 1 1 56257
0 2989 7 1 2 56255 56258
0 2990 7 1 2 56244 2989
0 2991 5 1 1 2990
0 2992 7 1 2 2980 2991
0 2993 5 1 1 2992
0 2994 7 1 2 56168 2993
0 2995 5 1 1 2994
0 2996 7 4 2 43822 47708
0 2997 7 1 2 45369 50897
0 2998 7 1 2 53700 2997
0 2999 5 1 1 2998
0 3000 7 17 2 53569 54753
0 3001 7 6 2 43682 47853
0 3002 7 1 2 56052 56289
0 3003 7 1 2 56272 3002
0 3004 5 1 1 3003
0 3005 7 1 2 2999 3004
0 3006 5 1 1 3005
0 3007 7 1 2 56268 3006
0 3008 5 1 1 3007
0 3009 7 2 2 47190 56062
0 3010 7 1 2 56245 56295
0 3011 7 4 2 43425 56182
0 3012 5 1 1 56297
0 3013 7 4 2 47854 50491
0 3014 7 1 2 56298 56301
0 3015 7 1 2 3010 3014
0 3016 5 1 1 3015
0 3017 7 1 2 3008 3016
0 3018 5 1 1 3017
0 3019 7 1 2 49832 3018
0 3020 5 1 1 3019
0 3021 7 1 2 2995 3020
0 3022 7 1 2 2954 3021
0 3023 7 1 2 2818 3022
0 3024 5 1 1 3023
0 3025 7 1 2 55553 3024
0 3026 5 1 1 3025
0 3027 7 1 2 43683 52703
0 3028 5 1 1 3027
0 3029 7 1 2 43823 53545
0 3030 5 1 1 3029
0 3031 7 1 2 206 3030
0 3032 5 1 1 3031
0 3033 7 1 2 52498 53772
0 3034 7 1 2 3032 3033
0 3035 5 1 1 3034
0 3036 7 1 2 3028 3035
0 3037 5 1 1 3036
0 3038 7 1 2 42452 3037
0 3039 5 1 1 3038
0 3040 7 1 2 43824 50386
0 3041 5 1 1 3040
0 3042 7 7 2 47191 48522
0 3043 5 2 1 56305
0 3044 7 2 2 49439 56306
0 3045 5 3 1 56314
0 3046 7 1 2 3041 56316
0 3047 5 1 1 3046
0 3048 7 1 2 42984 3047
0 3049 5 1 1 3048
0 3050 7 1 2 50219 52662
0 3051 5 1 1 3050
0 3052 7 8 2 45170 52608
0 3053 5 1 1 56319
0 3054 7 2 2 49326 56320
0 3055 5 3 1 56327
0 3056 7 1 2 3051 56329
0 3057 5 1 1 3056
0 3058 7 1 2 42686 3057
0 3059 5 1 1 3058
0 3060 7 3 2 51496 53107
0 3061 5 1 1 56332
0 3062 7 1 2 3059 3061
0 3063 7 1 2 3049 3062
0 3064 5 1 1 3063
0 3065 7 1 2 54554 3064
0 3066 5 1 1 3065
0 3067 7 1 2 3039 3066
0 3068 5 1 1 3067
0 3069 7 1 2 48064 3068
0 3070 5 1 1 3069
0 3071 7 7 2 42687 53519
0 3072 7 2 2 51126 56335
0 3073 7 1 2 50136 55497
0 3074 7 1 2 56342 3073
0 3075 5 1 1 3074
0 3076 7 1 2 3070 3075
0 3077 5 1 1 3076
0 3078 7 17 2 47945 48743
0 3079 7 2 2 55952 56344
0 3080 7 1 2 3077 56361
0 3081 5 1 1 3080
0 3082 7 1 2 44378 3081
0 3083 5 1 1 3082
0 3084 7 2 2 45951 54584
0 3085 5 1 1 56363
0 3086 7 5 2 42453 45031
0 3087 5 2 1 56365
0 3088 7 1 2 52991 56366
0 3089 5 1 1 3088
0 3090 7 6 2 42454 52016
0 3091 5 1 1 56372
0 3092 7 1 2 50975 56373
0 3093 5 1 1 3092
0 3094 7 1 2 48523 3093
0 3095 7 1 2 3089 3094
0 3096 7 1 2 3085 3095
0 3097 5 1 1 3096
0 3098 7 1 2 45952 54047
0 3099 5 1 1 3098
0 3100 7 1 2 55227 56367
0 3101 5 1 1 3100
0 3102 7 1 2 45171 3101
0 3103 7 1 2 3099 3102
0 3104 5 1 1 3103
0 3105 7 1 2 47058 3104
0 3106 7 1 2 3097 3105
0 3107 5 1 1 3106
0 3108 7 1 2 45953 55645
0 3109 7 1 2 55334 3108
0 3110 5 1 1 3109
0 3111 7 1 2 3107 3110
0 3112 5 1 1 3111
0 3113 7 2 2 44873 51582
0 3114 7 2 2 48744 50492
0 3115 7 1 2 56378 56380
0 3116 7 1 2 3112 3115
0 3117 5 1 1 3116
0 3118 7 1 2 43825 50641
0 3119 5 1 1 3118
0 3120 7 1 2 42985 53481
0 3121 7 1 2 53761 3120
0 3122 5 1 1 3121
0 3123 7 1 2 3119 3122
0 3124 5 1 1 3123
0 3125 7 1 2 42688 3124
0 3126 5 1 1 3125
0 3127 7 2 2 54888 3126
0 3128 5 1 1 56382
0 3129 7 1 2 45954 56383
0 3130 5 1 1 3129
0 3131 7 1 2 50525 52017
0 3132 5 2 1 3131
0 3133 7 1 2 46402 55357
0 3134 5 1 1 3133
0 3135 7 2 2 56384 3134
0 3136 5 1 1 56386
0 3137 7 1 2 42455 56387
0 3138 5 1 1 3137
0 3139 7 1 2 52133 53174
0 3140 5 1 1 3139
0 3141 7 9 2 47855 44874
0 3142 7 4 2 47059 50493
0 3143 7 1 2 56388 56397
0 3144 5 2 1 3143
0 3145 7 1 2 3140 56401
0 3146 5 5 1 3145
0 3147 7 1 2 46884 56403
0 3148 7 1 2 3138 3147
0 3149 7 1 2 3130 3148
0 3150 5 1 1 3149
0 3151 7 1 2 47709 3150
0 3152 7 1 2 3117 3151
0 3153 5 1 1 3152
0 3154 7 1 2 45668 3153
0 3155 7 1 2 3083 3154
0 3156 5 1 1 3155
0 3157 7 3 2 47060 47710
0 3158 7 2 2 54439 56408
0 3159 5 1 1 56411
0 3160 7 1 2 52698 56412
0 3161 5 1 1 3160
0 3162 7 19 2 44379 47856
0 3163 7 5 2 47946 56413
0 3164 7 6 2 43684 52152
0 3165 5 2 1 56437
0 3166 7 1 2 47061 51246
0 3167 5 2 1 3166
0 3168 7 1 2 56443 56445
0 3169 5 5 1 3168
0 3170 7 1 2 50932 54546
0 3171 7 1 2 56447 3170
0 3172 5 1 1 3171
0 3173 7 1 2 48065 52134
0 3174 7 1 2 52699 3173
0 3175 5 1 1 3174
0 3176 7 1 2 3172 3175
0 3177 5 1 1 3176
0 3178 7 1 2 56432 3177
0 3179 5 1 1 3178
0 3180 7 1 2 3161 3179
0 3181 5 1 1 3180
0 3182 7 1 2 42456 3181
0 3183 5 1 1 3182
0 3184 7 7 2 43685 44380
0 3185 7 4 2 47857 48066
0 3186 7 3 2 55215 56459
0 3187 7 1 2 56452 56463
0 3188 5 1 1 3187
0 3189 7 1 2 3159 3188
0 3190 5 2 1 3189
0 3191 7 1 2 56466 56364
0 3192 5 1 1 3191
0 3193 7 1 2 48524 3192
0 3194 7 1 2 3183 3193
0 3195 5 1 1 3194
0 3196 7 2 2 45955 53520
0 3197 7 1 2 51841 56468
0 3198 5 1 1 3197
0 3199 7 1 2 1944 3198
0 3200 5 1 1 3199
0 3201 7 1 2 56467 3200
0 3202 5 1 1 3201
0 3203 7 3 2 42689 56414
0 3204 7 9 2 52118 55216
0 3205 7 1 2 56470 56473
0 3206 5 1 1 3205
0 3207 7 3 2 47711 44716
0 3208 7 7 2 54494 56482
0 3209 7 2 2 54596 56485
0 3210 5 2 1 56492
0 3211 7 1 2 3206 56494
0 3212 5 1 1 3211
0 3213 7 1 2 42986 53229
0 3214 7 1 2 3212 3213
0 3215 5 1 1 3214
0 3216 7 1 2 45172 3215
0 3217 7 1 2 3202 3216
0 3218 5 1 1 3217
0 3219 7 7 2 46885 48745
0 3220 7 1 2 3218 56496
0 3221 7 1 2 3195 3220
0 3222 5 1 1 3221
0 3223 7 7 2 43986 49853
0 3224 7 5 2 42457 43826
0 3225 7 2 2 56503 56510
0 3226 7 5 2 47947 55771
0 3227 7 6 2 42690 43509
0 3228 7 1 2 42987 56522
0 3229 7 1 2 56438 3228
0 3230 7 1 2 56517 3229
0 3231 7 1 2 56515 3230
0 3232 5 1 1 3231
0 3233 7 1 2 3222 3232
0 3234 5 1 1 3233
0 3235 7 1 2 42125 3234
0 3236 5 1 1 3235
0 3237 7 2 2 45956 53570
0 3238 7 1 2 52700 56486
0 3239 5 1 1 3238
0 3240 7 4 2 43827 54205
0 3241 7 2 2 43987 56415
0 3242 7 1 2 52125 56534
0 3243 7 1 2 56530 3242
0 3244 5 1 1 3243
0 3245 7 1 2 3239 3244
0 3246 5 1 1 3245
0 3247 7 1 2 56528 3246
0 3248 5 1 1 3247
0 3249 7 3 2 42458 44381
0 3250 7 3 2 53571 56536
0 3251 7 1 2 53553 56539
0 3252 7 1 2 54585 3251
0 3253 5 1 1 3252
0 3254 7 1 2 3248 3253
0 3255 5 1 1 3254
0 3256 7 1 2 48525 3255
0 3257 5 1 1 3256
0 3258 7 3 2 51558 52264
0 3259 7 1 2 56540 56542
0 3260 7 1 2 54048 3259
0 3261 5 1 1 3260
0 3262 7 1 2 3257 3261
0 3263 5 1 1 3262
0 3264 7 1 2 48746 3263
0 3265 5 1 1 3264
0 3266 7 2 2 47712 53300
0 3267 7 5 2 42459 50652
0 3268 7 3 2 44525 56547
0 3269 7 1 2 56552 3128
0 3270 5 1 1 3269
0 3271 7 5 2 45957 50904
0 3272 7 1 2 56555 3136
0 3273 5 1 1 3272
0 3274 7 1 2 3270 3273
0 3275 5 1 1 3274
0 3276 7 1 2 56545 3275
0 3277 5 1 1 3276
0 3278 7 1 2 3265 3277
0 3279 5 1 1 3278
0 3280 7 1 2 53909 3279
0 3281 5 1 1 3280
0 3282 7 1 2 3236 3281
0 3283 7 1 2 3156 3282
0 3284 5 1 1 3283
0 3285 7 1 2 41968 3284
0 3286 5 1 1 3285
0 3287 7 1 2 54750 3286
0 3288 5 1 1 3287
0 3289 7 1 2 51420 54676
0 3290 5 1 1 3289
0 3291 7 1 2 43828 50518
0 3292 5 1 1 3291
0 3293 7 1 2 3290 3292
0 3294 5 1 1 3293
0 3295 7 1 2 42691 3294
0 3296 5 1 1 3295
0 3297 7 1 2 54889 3296
0 3298 5 1 1 3297
0 3299 7 1 2 3298 56553
0 3300 5 1 1 3299
0 3301 7 1 2 46403 55354
0 3302 5 1 1 3301
0 3303 7 1 2 56385 3302
0 3304 5 1 1 3303
0 3305 7 1 2 3304 56556
0 3306 5 1 1 3305
0 3307 7 1 2 3300 3306
0 3308 5 1 1 3307
0 3309 7 1 2 43510 3308
0 3310 5 1 1 3309
0 3311 7 1 2 50653 52145
0 3312 7 6 2 47858 48526
0 3313 7 1 2 53054 54307
0 3314 7 1 2 56560 3313
0 3315 7 1 2 3311 3314
0 3316 5 1 1 3315
0 3317 7 1 2 3310 3316
0 3318 5 1 1 3317
0 3319 7 1 2 42126 3318
0 3320 5 1 1 3319
0 3321 7 1 2 50237 51961
0 3322 7 6 2 47859 50654
0 3323 7 1 2 52529 56566
0 3324 7 1 2 3321 3323
0 3325 5 1 1 3324
0 3326 7 1 2 3320 3325
0 3327 5 1 1 3326
0 3328 7 1 2 53910 3327
0 3329 5 1 1 3328
0 3330 7 3 2 43511 56404
0 3331 7 1 2 53026 55145
0 3332 5 1 1 3331
0 3333 7 3 2 42692 52711
0 3334 5 2 1 56575
0 3335 7 1 2 45958 56576
0 3336 5 1 1 3335
0 3337 7 1 2 3332 3336
0 3338 5 1 1 3337
0 3339 7 1 2 56572 3338
0 3340 5 1 1 3339
0 3341 7 1 2 51626 632
0 3342 5 13 1 3341
0 3343 7 3 2 48527 56580
0 3344 5 1 1 56593
0 3345 7 3 2 42693 48067
0 3346 7 3 2 42460 56596
0 3347 7 1 2 55532 56599
0 3348 7 1 2 56594 3347
0 3349 5 1 1 3348
0 3350 7 1 2 50494 50911
0 3351 7 1 2 55953 3350
0 3352 7 1 2 53027 3351
0 3353 5 1 1 3352
0 3354 7 1 2 3349 3353
0 3355 5 1 1 3354
0 3356 7 1 2 53911 3355
0 3357 5 1 1 3356
0 3358 7 2 2 48068 52561
0 3359 7 2 2 53183 56602
0 3360 5 1 1 56604
0 3361 7 3 2 42694 51655
0 3362 5 1 1 56606
0 3363 7 1 2 55533 56607
0 3364 7 1 2 56605 3363
0 3365 5 1 1 3364
0 3366 7 1 2 3357 3365
0 3367 7 1 2 3340 3366
0 3368 5 1 1 3367
0 3369 7 1 2 42127 3368
0 3370 5 1 1 3369
0 3371 7 4 2 48069 48528
0 3372 7 1 2 54558 56609
0 3373 5 1 1 3372
0 3374 7 1 2 3360 3373
0 3375 5 1 1 3374
0 3376 7 4 2 47948 55954
0 3377 7 1 2 45669 54206
0 3378 7 1 2 56613 3377
0 3379 7 1 2 3375 3378
0 3380 5 1 1 3379
0 3381 7 1 2 3370 3380
0 3382 5 1 1 3381
0 3383 7 1 2 54260 3382
0 3384 5 1 1 3383
0 3385 7 4 2 45959 51962
0 3386 5 2 1 56617
0 3387 7 1 2 3091 56621
0 3388 5 2 1 3387
0 3389 7 1 2 50526 56573
0 3390 5 1 1 3389
0 3391 7 4 2 48212 50220
0 3392 7 1 2 48070 54649
0 3393 7 2 2 56625 3392
0 3394 7 1 2 55664 56629
0 3395 5 1 1 3394
0 3396 7 1 2 3390 3395
0 3397 5 1 1 3396
0 3398 7 1 2 42128 3397
0 3399 5 1 1 3398
0 3400 7 1 2 56057 56630
0 3401 5 1 1 3400
0 3402 7 1 2 3399 3401
0 3403 5 1 1 3402
0 3404 7 1 2 56623 3403
0 3405 5 1 1 3404
0 3406 7 1 2 42461 55355
0 3407 5 1 1 3406
0 3408 7 6 2 45960 43829
0 3409 7 3 2 49448 56631
0 3410 5 1 1 56637
0 3411 7 1 2 3407 3410
0 3412 5 1 1 3411
0 3413 7 1 2 46404 3412
0 3414 5 1 1 3413
0 3415 7 2 2 42988 54685
0 3416 5 1 1 56640
0 3417 7 1 2 45173 56641
0 3418 5 1 1 3417
0 3419 7 1 2 3414 3418
0 3420 5 1 1 3419
0 3421 7 1 2 42129 56574
0 3422 7 1 2 3420 3421
0 3423 5 1 1 3422
0 3424 7 1 2 3405 3423
0 3425 7 1 2 3384 3424
0 3426 7 1 2 3329 3425
0 3427 5 1 1 3426
0 3428 7 1 2 47713 3427
0 3429 5 1 1 3428
0 3430 7 1 2 48916 3429
0 3431 5 1 1 3430
0 3432 7 1 2 50813 3431
0 3433 7 1 2 3288 3432
0 3434 5 1 1 3433
0 3435 7 1 2 3026 3434
0 3436 7 1 2 2558 3435
0 3437 7 1 2 1335 3436
0 3438 5 1 1 3437
0 3439 7 1 2 44278 3438
0 3440 5 1 1 3439
0 3441 7 6 2 48529 50814
0 3442 5 16 1 56642
0 3443 7 2 2 50892 56648
0 3444 5 1 1 56664
0 3445 7 4 2 49731 56665
0 3446 5 3 1 56666
0 3447 7 1 2 50044 52880
0 3448 5 1 1 3447
0 3449 7 3 2 56670 3448
0 3450 7 2 2 45032 56673
0 3451 5 1 1 56676
0 3452 7 1 2 49401 3451
0 3453 5 1 1 3452
0 3454 7 2 2 48213 3453
0 3455 7 3 2 43830 50655
0 3456 7 4 2 54528 56680
0 3457 7 3 2 46886 56683
0 3458 7 1 2 56678 56687
0 3459 5 1 1 3458
0 3460 7 1 2 53801 54106
0 3461 5 1 1 3460
0 3462 7 2 2 49732 51994
0 3463 5 2 1 56690
0 3464 7 1 2 52051 54050
0 3465 7 1 2 56692 3464
0 3466 5 1 1 3465
0 3467 7 1 2 3461 3466
0 3468 5 1 1 3467
0 3469 7 1 2 44151 3468
0 3470 5 1 1 3469
0 3471 7 5 2 48530 54823
0 3472 7 1 2 43831 56694
0 3473 5 1 1 3472
0 3474 7 1 2 3470 3473
0 3475 5 1 1 3474
0 3476 7 1 2 43212 3475
0 3477 5 1 1 3476
0 3478 7 8 2 47356 47491
0 3479 5 2 1 56699
0 3480 7 6 2 46600 56700
0 3481 5 1 1 56709
0 3482 7 3 2 45174 55650
0 3483 7 2 2 56710 56715
0 3484 5 1 1 56718
0 3485 7 1 2 49188 56695
0 3486 5 1 1 3485
0 3487 7 1 2 3484 3486
0 3488 5 1 1 3487
0 3489 7 1 2 43832 3488
0 3490 5 1 1 3489
0 3491 7 4 2 48531 54712
0 3492 5 1 1 56720
0 3493 7 1 2 54722 56721
0 3494 5 1 1 3493
0 3495 7 1 2 3490 3494
0 3496 7 1 2 3477 3495
0 3497 5 1 1 3496
0 3498 7 1 2 45033 3497
0 3499 5 1 1 3498
0 3500 7 9 2 42695 48532
0 3501 5 1 1 56724
0 3502 7 2 2 54051 56725
0 3503 7 1 2 50815 56733
0 3504 5 1 1 3503
0 3505 7 7 2 45175 50045
0 3506 5 14 1 56735
0 3507 7 1 2 53802 56736
0 3508 5 1 1 3507
0 3509 7 1 2 3504 3508
0 3510 5 1 1 3509
0 3511 7 1 2 47192 3510
0 3512 5 1 1 3511
0 3513 7 4 2 45176 55554
0 3514 7 1 2 49481 54824
0 3515 7 1 2 56756 3514
0 3516 5 1 1 3515
0 3517 7 1 2 3512 3516
0 3518 5 1 1 3517
0 3519 7 1 2 48387 3518
0 3520 5 1 1 3519
0 3521 7 4 2 45177 49189
0 3522 5 1 1 56760
0 3523 7 1 2 55295 3522
0 3524 5 4 1 3523
0 3525 7 3 2 44875 56764
0 3526 7 2 2 52951 55370
0 3527 7 1 2 56768 56771
0 3528 5 1 1 3527
0 3529 7 1 2 3520 3528
0 3530 7 1 2 3499 3529
0 3531 5 1 1 3530
0 3532 7 1 2 47062 3531
0 3533 5 1 1 3532
0 3534 7 13 2 46601 43833
0 3535 7 4 2 49141 56773
0 3536 5 5 1 56786
0 3537 7 8 2 47193 44152
0 3538 5 1 1 56795
0 3539 7 2 2 48747 56796
0 3540 7 1 2 43213 56803
0 3541 5 1 1 3540
0 3542 7 1 2 56790 3541
0 3543 5 2 1 3542
0 3544 7 1 2 50532 56805
0 3545 5 1 1 3544
0 3546 7 2 2 47194 53722
0 3547 5 1 1 56807
0 3548 7 1 2 52311 56808
0 3549 5 1 1 3548
0 3550 7 1 2 3545 3549
0 3551 5 2 1 3550
0 3552 7 1 2 44876 55646
0 3553 7 1 2 56809 3552
0 3554 5 1 1 3553
0 3555 7 1 2 3533 3554
0 3556 5 1 1 3555
0 3557 7 1 2 52545 3556
0 3558 5 1 1 3557
0 3559 7 1 2 3459 3558
0 3560 5 1 1 3559
0 3561 7 1 2 44526 3560
0 3562 5 1 1 3561
0 3563 7 17 2 47063 47195
0 3564 5 1 1 56811
0 3565 7 5 2 46135 56812
0 3566 7 3 2 50905 56828
0 3567 5 1 1 56833
0 3568 7 1 2 46887 56834
0 3569 7 1 2 56679 3568
0 3570 5 1 1 3569
0 3571 7 1 2 3562 3570
0 3572 5 1 1 3571
0 3573 7 1 2 43426 3572
0 3574 5 1 1 3573
0 3575 7 3 2 47357 50046
0 3576 5 4 1 56836
0 3577 7 2 2 50593 56742
0 3578 7 3 2 56839 56843
0 3579 5 5 1 56845
0 3580 7 1 2 45034 56848
0 3581 5 1 1 3580
0 3582 7 1 2 48388 52196
0 3583 5 4 1 3582
0 3584 7 1 2 50201 56853
0 3585 7 2 2 3581 3584
0 3586 7 4 2 42696 47860
0 3587 7 1 2 48071 51884
0 3588 7 1 2 56859 3587
0 3589 7 1 2 54652 3588
0 3590 7 1 2 56857 3589
0 3591 5 1 1 3590
0 3592 7 1 2 3574 3591
0 3593 5 1 1 3592
0 3594 7 1 2 44382 3593
0 3595 5 1 1 3594
0 3596 7 17 2 46136 46789
0 3597 7 2 2 56296 56863
0 3598 7 1 2 56487 56880
0 3599 7 1 2 56858 3598
0 3600 5 1 1 3599
0 3601 7 1 2 3595 3600
0 3602 5 1 1 3601
0 3603 7 1 2 42989 3602
0 3604 5 1 1 3603
0 3605 7 11 2 43988 47492
0 3606 5 4 1 56882
0 3607 7 3 2 46602 56883
0 3608 5 3 1 56897
0 3609 7 8 2 47861 55839
0 3610 5 2 1 56903
0 3611 7 11 2 46888 47714
0 3612 7 5 2 44527 56913
0 3613 5 2 1 56924
0 3614 7 1 2 45370 56925
0 3615 5 1 1 3614
0 3616 7 1 2 56911 3615
0 3617 5 4 1 3616
0 3618 7 1 2 56684 56931
0 3619 5 1 1 3618
0 3620 7 4 2 47196 47715
0 3621 7 5 2 50495 54089
0 3622 7 2 2 56935 56939
0 3623 7 16 2 47862 45371
0 3624 7 4 2 46889 56946
0 3625 5 1 1 56962
0 3626 7 1 2 51627 3625
0 3627 5 11 1 3626
0 3628 7 1 2 56944 56966
0 3629 5 1 1 3628
0 3630 7 1 2 3619 3629
0 3631 5 1 1 3630
0 3632 7 1 2 56898 3631
0 3633 5 1 1 3632
0 3634 7 2 2 47358 51656
0 3635 7 1 2 48748 56977
0 3636 5 1 1 3635
0 3637 7 1 2 55722 3636
0 3638 5 1 1 3637
0 3639 7 1 2 56945 3638
0 3640 5 1 1 3639
0 3641 7 2 2 55840 56685
0 3642 5 1 1 56979
0 3643 7 1 2 56947 56980
0 3644 5 1 1 3643
0 3645 7 1 2 3640 3644
0 3646 5 1 1 3645
0 3647 7 1 2 55555 3646
0 3648 5 1 1 3647
0 3649 7 3 2 45372 52741
0 3650 5 1 1 56981
0 3651 7 2 2 56398 56982
0 3652 7 2 2 46137 44153
0 3653 5 2 1 56986
0 3654 7 8 2 43214 47863
0 3655 7 1 2 56914 56990
0 3656 7 1 2 56987 3655
0 3657 7 1 2 56984 3656
0 3658 5 1 1 3657
0 3659 7 1 2 3648 3658
0 3660 7 1 2 3633 3659
0 3661 5 1 1 3660
0 3662 7 1 2 46790 3661
0 3663 5 1 1 3662
0 3664 7 1 2 53394 56967
0 3665 5 1 1 3664
0 3666 7 1 2 43834 55280
0 3667 5 3 1 3666
0 3668 7 1 2 51698 56998
0 3669 5 1 1 3668
0 3670 7 1 2 3665 3669
0 3671 5 1 1 3670
0 3672 7 1 2 56940 3671
0 3673 5 1 1 3672
0 3674 7 4 2 42697 45373
0 3675 5 1 1 57001
0 3676 7 1 2 55136 55743
0 3677 7 1 2 57002 3676
0 3678 7 1 2 53175 3677
0 3679 5 1 1 3678
0 3680 7 1 2 3673 3679
0 3681 5 1 1 3680
0 3682 7 1 2 55874 3681
0 3683 5 1 1 3682
0 3684 7 1 2 3663 3683
0 3685 5 1 1 3684
0 3686 7 1 2 48533 3685
0 3687 5 1 1 3686
0 3688 7 16 2 46138 46603
0 3689 7 3 2 50496 57005
0 3690 7 1 2 56761 57021
0 3691 7 6 2 47716 47864
0 3692 7 2 2 43989 57024
0 3693 7 3 2 46791 56813
0 3694 7 1 2 57030 57032
0 3695 7 1 2 3690 3694
0 3696 5 1 1 3695
0 3697 7 6 2 42698 54155
0 3698 7 3 2 52799 57035
0 3699 5 1 1 57041
0 3700 7 1 2 3567 3699
0 3701 5 1 1 3700
0 3702 7 2 2 51738 3701
0 3703 7 1 2 49733 55875
0 3704 7 1 2 57044 3703
0 3705 5 1 1 3704
0 3706 7 1 2 3696 3705
0 3707 5 1 1 3706
0 3708 7 1 2 46890 3707
0 3709 5 1 1 3708
0 3710 7 2 2 49943 53378
0 3711 5 1 1 57046
0 3712 7 1 2 48749 53484
0 3713 5 1 1 3712
0 3714 7 1 2 57047 3713
0 3715 5 1 1 3714
0 3716 7 9 2 43835 45374
0 3717 7 2 2 52190 57048
0 3718 5 2 1 57057
0 3719 7 1 2 3715 57059
0 3720 5 1 1 3719
0 3721 7 3 2 46139 43512
0 3722 7 2 2 44383 50497
0 3723 7 1 2 47064 54458
0 3724 7 3 2 57064 3723
0 3725 7 1 2 57061 57066
0 3726 7 1 2 3720 3725
0 3727 5 1 1 3726
0 3728 7 1 2 3709 3727
0 3729 7 1 2 3687 3728
0 3730 5 1 1 3729
0 3731 7 1 2 48214 3730
0 3732 5 1 1 3731
0 3733 7 1 2 49839 52803
0 3734 5 2 1 3733
0 3735 7 4 2 48750 56757
0 3736 5 3 1 57071
0 3737 7 1 2 57069 57075
0 3738 5 1 1 3737
0 3739 7 1 2 47197 3738
0 3740 5 1 1 3739
0 3741 7 6 2 46140 45375
0 3742 5 2 1 57078
0 3743 7 7 2 47493 48534
0 3744 7 2 2 46604 57086
0 3745 5 9 1 57093
0 3746 7 2 2 52817 57095
0 3747 5 9 1 57104
0 3748 7 1 2 57079 57106
0 3749 5 1 1 3748
0 3750 7 1 2 3740 3749
0 3751 5 1 1 3750
0 3752 7 1 2 47359 3751
0 3753 5 1 1 3752
0 3754 7 6 2 43215 56797
0 3755 5 4 1 57115
0 3756 7 1 2 52178 56774
0 3757 5 3 1 3756
0 3758 7 1 2 57121 57125
0 3759 5 2 1 3758
0 3760 7 1 2 57080 57128
0 3761 5 1 1 3760
0 3762 7 1 2 3753 3761
0 3763 5 1 1 3762
0 3764 7 5 2 43427 43686
0 3765 7 1 2 55841 57130
0 3766 7 1 2 54440 3765
0 3767 7 1 2 3763 3766
0 3768 5 1 1 3767
0 3769 7 1 2 3732 3768
0 3770 5 1 1 3769
0 3771 7 1 2 48389 3770
0 3772 5 1 1 3771
0 3773 7 5 2 44615 45035
0 3774 7 5 2 43836 45178
0 3775 5 2 1 57140
0 3776 7 7 2 47360 48751
0 3777 5 1 1 57147
0 3778 7 2 2 49607 57148
0 3779 5 1 1 57154
0 3780 7 1 2 57145 3779
0 3781 5 2 1 3780
0 3782 7 2 2 43216 57156
0 3783 5 1 1 57158
0 3784 7 7 2 46605 49190
0 3785 5 2 1 57160
0 3786 7 1 2 43837 57161
0 3787 5 1 1 3786
0 3788 7 1 2 3783 3787
0 3789 5 1 1 3788
0 3790 7 1 2 46141 3789
0 3791 5 1 1 3790
0 3792 7 2 2 43838 50533
0 3793 5 3 1 57169
0 3794 7 2 2 55692 57171
0 3795 5 12 1 57174
0 3796 7 1 2 57162 57176
0 3797 5 1 1 3796
0 3798 7 1 2 3791 3797
0 3799 5 2 1 3798
0 3800 7 15 2 43687 44717
0 3801 7 1 2 57188 57190
0 3802 5 1 1 3801
0 3803 7 7 2 46606 47065
0 3804 5 1 1 57205
0 3805 7 5 2 48072 52018
0 3806 7 1 2 57206 57212
0 3807 7 1 2 53821 3806
0 3808 5 1 1 3807
0 3809 7 1 2 3802 3808
0 3810 5 1 1 3809
0 3811 7 1 2 51583 3810
0 3812 5 1 1 3811
0 3813 7 10 2 47066 48073
0 3814 7 2 2 52019 57217
0 3815 5 2 1 57227
0 3816 7 1 2 44718 57036
0 3817 5 1 1 3816
0 3818 7 1 2 57229 3817
0 3819 5 5 1 3818
0 3820 7 1 2 45376 55811
0 3821 7 2 2 57231 3820
0 3822 7 2 2 46891 47494
0 3823 7 1 2 47361 57238
0 3824 7 1 2 57236 3823
0 3825 5 1 1 3824
0 3826 7 1 2 3812 3825
0 3827 5 1 1 3826
0 3828 7 1 2 44877 3827
0 3829 5 1 1 3828
0 3830 7 11 2 43217 47067
0 3831 7 5 2 43839 44154
0 3832 7 2 2 57240 57251
0 3833 5 1 1 57256
0 3834 7 2 2 43688 56667
0 3835 5 1 1 57258
0 3836 7 1 2 47198 57259
0 3837 5 1 1 3836
0 3838 7 1 2 3833 3837
0 3839 5 1 1 3838
0 3840 7 3 2 48215 54420
0 3841 7 1 2 45377 57062
0 3842 7 1 2 57260 3841
0 3843 7 1 2 3839 3842
0 3844 5 1 1 3843
0 3845 7 1 2 3829 3844
0 3846 5 1 1 3845
0 3847 7 1 2 55876 3846
0 3848 5 1 1 3847
0 3849 7 5 2 46607 51657
0 3850 5 1 1 57263
0 3851 7 1 2 51628 3850
0 3852 5 2 1 3851
0 3853 7 2 2 47717 48955
0 3854 7 5 2 46792 47495
0 3855 7 6 2 47362 44878
0 3856 7 1 2 57272 57277
0 3857 7 1 2 57270 3856
0 3858 7 1 2 57268 3857
0 3859 7 1 2 57232 3858
0 3860 5 1 1 3859
0 3861 7 1 2 3848 3860
0 3862 5 1 1 3861
0 3863 7 1 2 57135 3862
0 3864 5 1 1 3863
0 3865 7 1 2 3772 3864
0 3866 5 1 1 3865
0 3867 7 1 2 46405 3866
0 3868 5 1 1 3867
0 3869 7 2 2 42699 51700
0 3870 5 1 1 57283
0 3871 7 1 2 52705 57284
0 3872 5 1 1 3871
0 3873 7 8 2 47496 48216
0 3874 7 2 2 45378 57285
0 3875 5 1 1 57293
0 3876 7 2 2 57006 57294
0 3877 5 2 1 57295
0 3878 7 1 2 3872 57297
0 3879 5 1 1 3878
0 3880 7 1 2 48535 3879
0 3881 5 1 1 3880
0 3882 7 3 2 48217 49734
0 3883 7 2 2 49944 57081
0 3884 5 1 1 57302
0 3885 7 1 2 57299 57303
0 3886 5 1 1 3885
0 3887 7 1 2 3881 3886
0 3888 5 1 1 3887
0 3889 7 1 2 47199 3888
0 3890 5 1 1 3889
0 3891 7 1 2 47363 57296
0 3892 5 1 1 3891
0 3893 7 11 2 48752 55556
0 3894 5 3 1 57304
0 3895 7 1 2 54825 57305
0 3896 5 1 1 3895
0 3897 7 1 2 3892 3896
0 3898 5 1 1 3897
0 3899 7 1 2 57141 3898
0 3900 5 1 1 3899
0 3901 7 1 2 3890 3900
0 3902 5 1 1 3901
0 3903 7 1 2 48390 3902
0 3904 5 1 1 3903
0 3905 7 8 2 47364 44155
0 3906 5 3 1 57318
0 3907 7 3 2 43218 57319
0 3908 5 3 1 57329
0 3909 7 1 2 57096 57332
0 3910 5 2 1 3909
0 3911 7 2 2 45379 57335
0 3912 7 1 2 55156 57337
0 3913 5 1 1 3912
0 3914 7 1 2 55519 57306
0 3915 5 1 1 3914
0 3916 7 18 2 46142 43219
0 3917 5 1 1 57339
0 3918 7 9 2 44156 57340
0 3919 5 1 1 57357
0 3920 7 1 2 57049 57358
0 3921 5 1 1 3920
0 3922 7 1 2 3915 3921
0 3923 5 1 1 3922
0 3924 7 1 2 45179 3923
0 3925 5 1 1 3924
0 3926 7 1 2 3913 3925
0 3927 5 1 1 3926
0 3928 7 1 2 49643 3927
0 3929 5 1 1 3928
0 3930 7 1 2 47068 3929
0 3931 7 1 2 3904 3930
0 3932 5 1 1 3931
0 3933 7 17 2 45380 50732
0 3934 7 1 2 49854 57366
0 3935 5 1 1 3934
0 3936 7 1 2 117 52878
0 3937 5 1 1 3936
0 3938 7 2 2 68 52857
0 3939 5 3 1 57383
0 3940 7 1 2 49945 57384
0 3941 7 1 2 3937 3940
0 3942 5 1 1 3941
0 3943 7 1 2 3935 3942
0 3944 5 1 1 3943
0 3945 7 1 2 44879 3944
0 3946 5 1 1 3945
0 3947 7 1 2 45036 56719
0 3948 5 1 1 3947
0 3949 7 1 2 3946 3948
0 3950 5 1 1 3949
0 3951 7 1 2 52020 3950
0 3952 5 1 1 3951
0 3953 7 4 2 45381 52179
0 3954 7 13 2 43840 44880
0 3955 7 2 2 55371 57392
0 3956 7 1 2 49806 57405
0 3957 7 1 2 57388 3956
0 3958 5 1 1 3957
0 3959 7 1 2 43689 3958
0 3960 7 1 2 3952 3959
0 3961 5 1 1 3960
0 3962 7 1 2 44719 3961
0 3963 7 1 2 3932 3962
0 3964 5 1 1 3963
0 3965 7 2 2 50534 57218
0 3966 7 2 2 47200 57407
0 3967 5 1 1 57409
0 3968 7 5 2 47497 57007
0 3969 7 1 2 52284 57411
0 3970 7 1 2 57410 3969
0 3971 5 1 1 3970
0 3972 7 1 2 3964 3971
0 3973 5 1 1 3972
0 3974 7 1 2 44528 54665
0 3975 7 1 2 55842 3974
0 3976 7 1 2 3973 3975
0 3977 5 1 1 3976
0 3978 7 1 2 45670 3977
0 3979 7 1 2 3868 3978
0 3980 7 1 2 3604 3979
0 3981 5 1 1 3980
0 3982 7 10 2 46892 44529
0 3983 7 4 2 50733 56011
0 3984 7 1 2 56814 57426
0 3985 5 1 1 3984
0 3986 7 7 2 44720 48753
0 3987 7 2 2 49608 57430
0 3988 7 1 2 51360 57437
0 3989 5 1 1 3988
0 3990 7 1 2 3985 3989
0 3991 5 1 1 3990
0 3992 7 1 2 54946 3991
0 3993 5 1 1 3992
0 3994 7 3 2 43841 57191
0 3995 7 1 2 49191 57439
0 3996 5 1 1 3995
0 3997 7 1 2 57230 3996
0 3998 5 1 1 3997
0 3999 7 1 2 49906 3998
0 4000 5 1 1 3999
0 4001 7 2 2 42990 51361
0 4002 7 1 2 56798 57431
0 4003 7 1 2 57442 4002
0 4004 5 1 1 4003
0 4005 7 1 2 4000 4004
0 4006 5 1 1 4005
0 4007 7 1 2 45180 4006
0 4008 5 1 1 4007
0 4009 7 1 2 3993 4008
0 4010 5 1 1 4009
0 4011 7 1 2 55877 4010
0 4012 5 1 1 4011
0 4013 7 3 2 46406 55600
0 4014 5 2 1 57444
0 4015 7 3 2 46608 55878
0 4016 5 2 1 57449
0 4017 7 1 2 57447 57452
0 4018 5 2 1 4017
0 4019 7 1 2 57233 57454
0 4020 5 1 1 4019
0 4021 7 8 2 46609 44384
0 4022 7 2 2 55855 57456
0 4023 7 1 2 57440 57464
0 4024 5 1 1 4023
0 4025 7 1 2 4020 4024
0 4026 5 1 1 4025
0 4027 7 1 2 52352 4026
0 4028 5 1 1 4027
0 4029 7 1 2 4012 4028
0 4030 5 1 1 4029
0 4031 7 1 2 47365 4030
0 4032 5 1 1 4031
0 4033 7 2 2 55696 57192
0 4034 7 1 2 49192 57466
0 4035 5 1 1 4034
0 4036 7 1 2 49142 52265
0 4037 7 1 2 56829 4036
0 4038 5 1 1 4037
0 4039 7 1 2 4035 4038
0 4040 5 1 1 4039
0 4041 7 1 2 46610 4040
0 4042 5 1 1 4041
0 4043 7 2 2 46143 51362
0 4044 7 1 2 43842 51048
0 4045 7 1 2 57468 4044
0 4046 5 1 1 4045
0 4047 7 1 2 4042 4046
0 4048 5 1 1 4047
0 4049 7 1 2 46407 4048
0 4050 5 1 1 4049
0 4051 7 1 2 48754 57257
0 4052 5 1 1 4051
0 4053 7 1 2 54925 57367
0 4054 5 1 1 4053
0 4055 7 1 2 4052 4054
0 4056 5 2 1 4055
0 4057 7 1 2 53723 57470
0 4058 5 1 1 4057
0 4059 7 2 2 48536 54840
0 4060 7 2 2 43843 52326
0 4061 5 5 1 57474
0 4062 7 1 2 54346 57476
0 4063 5 1 1 4062
0 4064 7 1 2 57472 4063
0 4065 5 1 1 4064
0 4066 7 1 2 4058 4065
0 4067 5 1 1 4066
0 4068 7 1 2 42991 4067
0 4069 5 1 1 4068
0 4070 7 6 2 49609 53336
0 4071 5 2 1 57481
0 4072 7 1 2 55066 57482
0 4073 5 1 1 4072
0 4074 7 1 2 4069 4073
0 4075 5 1 1 4074
0 4076 7 1 2 44721 4075
0 4077 5 1 1 4076
0 4078 7 1 2 4050 4077
0 4079 5 1 1 4078
0 4080 7 1 2 55879 4079
0 4081 5 1 1 4080
0 4082 7 1 2 4032 4081
0 4083 5 1 1 4082
0 4084 7 1 2 57416 4083
0 4085 5 1 1 4084
0 4086 7 9 2 43513 47498
0 4087 7 6 2 46793 44385
0 4088 7 2 2 49262 57498
0 4089 7 1 2 57489 57504
0 4090 7 1 2 57237 4089
0 4091 5 1 1 4090
0 4092 7 1 2 4085 4091
0 4093 5 1 1 4092
0 4094 7 1 2 44881 4093
0 4095 5 1 1 4094
0 4096 7 4 2 43428 57417
0 4097 5 2 1 57506
0 4098 7 1 2 42700 57507
0 4099 7 1 2 56758 4098
0 4100 5 1 1 4099
0 4101 7 6 2 46794 55955
0 4102 5 1 1 57512
0 4103 7 1 2 56207 57513
0 4104 7 1 2 3444 4103
0 4105 5 1 1 4104
0 4106 7 1 2 4100 4105
0 4107 5 1 1 4106
0 4108 7 1 2 48755 4107
0 4109 5 1 1 4108
0 4110 7 1 2 57510 4102
0 4111 5 2 1 4110
0 4112 7 4 2 42992 56840
0 4113 5 1 1 57520
0 4114 7 4 2 56844 57521
0 4115 5 1 1 57524
0 4116 7 2 2 46144 57525
0 4117 5 1 1 57528
0 4118 7 1 2 57518 57529
0 4119 5 1 1 4118
0 4120 7 1 2 4109 4119
0 4121 5 1 1 4120
0 4122 7 1 2 56815 4121
0 4123 5 1 1 4122
0 4124 7 7 2 46145 48537
0 4125 5 3 1 57530
0 4126 7 1 2 54710 57537
0 4127 5 4 1 4126
0 4128 7 1 2 50734 57540
0 4129 5 2 1 4128
0 4130 7 9 2 43990 52712
0 4131 5 12 1 57546
0 4132 7 4 2 49946 57555
0 4133 5 1 1 57567
0 4134 7 1 2 46146 57568
0 4135 5 1 1 4134
0 4136 7 1 2 57544 4135
0 4137 5 2 1 4136
0 4138 7 1 2 53994 57508
0 4139 7 1 2 57571 4138
0 4140 5 1 1 4139
0 4141 7 8 2 46611 47366
0 4142 5 2 1 57573
0 4143 7 3 2 52180 57574
0 4144 5 1 1 57583
0 4145 7 1 2 46408 56668
0 4146 5 1 1 4145
0 4147 7 2 2 4144 4146
0 4148 5 2 1 57586
0 4149 7 9 2 46147 46893
0 4150 7 1 2 54459 54926
0 4151 7 1 2 57590 4150
0 4152 7 1 2 57588 4151
0 4153 5 1 1 4152
0 4154 7 1 2 4140 4153
0 4155 5 1 1 4154
0 4156 7 1 2 45382 4155
0 4157 5 1 1 4156
0 4158 7 1 2 4123 4157
0 4159 5 1 1 4158
0 4160 7 1 2 44386 4159
0 4161 5 1 1 4160
0 4162 7 4 2 48756 56846
0 4163 7 14 2 42993 46795
0 4164 7 5 2 57591 57603
0 4165 7 26 2 47718 44530
0 4166 7 1 2 56816 57622
0 4167 7 1 2 57617 4166
0 4168 7 1 2 57599 4167
0 4169 5 1 1 4168
0 4170 7 1 2 4161 4169
0 4171 5 1 1 4170
0 4172 7 1 2 52153 4171
0 4173 5 1 1 4172
0 4174 7 1 2 4095 4173
0 4175 5 1 1 4174
0 4176 7 1 2 45037 4175
0 4177 5 1 1 4176
0 4178 7 1 2 2566 55924
0 4179 5 2 1 4178
0 4180 7 7 2 47499 48757
0 4181 5 5 1 57650
0 4182 7 1 2 47719 57657
0 4183 5 1 1 4182
0 4184 7 2 2 57648 4183
0 4185 7 1 2 51393 57662
0 4186 5 1 1 4185
0 4187 7 1 2 55321 55880
0 4188 5 1 1 4187
0 4189 7 1 2 56884 57445
0 4190 5 1 1 4189
0 4191 7 1 2 4188 4190
0 4192 5 1 1 4191
0 4193 7 1 2 48538 4192
0 4194 5 1 1 4193
0 4195 7 1 2 4186 4194
0 4196 5 1 1 4195
0 4197 7 1 2 46612 4196
0 4198 5 1 1 4197
0 4199 7 4 2 47500 52887
0 4200 5 1 1 57664
0 4201 7 1 2 48758 49787
0 4202 5 1 1 4201
0 4203 7 1 2 57569 4202
0 4204 5 2 1 4203
0 4205 7 1 2 4200 57668
0 4206 5 1 1 4205
0 4207 7 1 2 55881 4206
0 4208 5 1 1 4207
0 4209 7 1 2 4198 4208
0 4210 5 1 1 4209
0 4211 7 1 2 47201 4210
0 4212 5 1 1 4211
0 4213 7 2 2 49947 51456
0 4214 5 1 1 57670
0 4215 7 1 2 50735 53950
0 4216 7 1 2 51077 4215
0 4217 5 1 1 4216
0 4218 7 1 2 4214 4217
0 4219 5 2 1 4218
0 4220 7 2 2 45383 57672
0 4221 7 1 2 55882 57674
0 4222 5 1 1 4221
0 4223 7 1 2 4212 4222
0 4224 5 1 1 4223
0 4225 7 1 2 52466 4224
0 4226 5 1 1 4225
0 4227 7 2 2 52234 57107
0 4228 5 1 1 57676
0 4229 7 1 2 46409 57129
0 4230 5 1 1 4229
0 4231 7 1 2 4228 4230
0 4232 5 2 1 4231
0 4233 7 8 2 44387 44882
0 4234 7 1 2 45384 57131
0 4235 7 1 2 57680 4234
0 4236 7 1 2 57678 4235
0 4237 5 1 1 4236
0 4238 7 1 2 4226 4237
0 4239 5 1 1 4238
0 4240 7 1 2 46148 4239
0 4241 5 1 1 4240
0 4242 7 3 2 49263 54927
0 4243 5 3 1 57688
0 4244 7 1 2 55982 57691
0 4245 5 1 1 4244
0 4246 7 5 2 44883 52841
0 4247 7 1 2 55883 57694
0 4248 7 1 2 4245 4247
0 4249 5 1 1 4248
0 4250 7 3 2 51056 56864
0 4251 7 3 2 47720 48218
0 4252 7 1 2 53319 57702
0 4253 7 1 2 57699 4252
0 4254 5 1 1 4253
0 4255 7 1 2 4249 4254
0 4256 5 1 1 4255
0 4257 7 1 2 55557 4256
0 4258 5 1 1 4257
0 4259 7 3 2 50816 55471
0 4260 7 1 2 57473 57705
0 4261 5 1 1 4260
0 4262 7 2 2 43690 53353
0 4263 7 3 2 48956 57320
0 4264 7 1 2 57708 57710
0 4265 5 1 1 4264
0 4266 7 1 2 4261 4265
0 4267 5 1 1 4266
0 4268 7 5 2 43429 47202
0 4269 7 1 2 57681 57713
0 4270 7 1 2 4267 4269
0 4271 5 1 1 4270
0 4272 7 1 2 4258 4271
0 4273 7 1 2 4241 4272
0 4274 5 1 1 4273
0 4275 7 1 2 57418 4274
0 4276 5 1 1 4275
0 4277 7 6 2 49735 51739
0 4278 7 2 2 46410 57718
0 4279 5 3 1 57724
0 4280 7 2 2 45385 57665
0 4281 5 1 1 57729
0 4282 7 1 2 57726 4281
0 4283 5 2 1 4282
0 4284 7 6 2 44388 48219
0 4285 7 1 2 47865 57733
0 4286 7 1 2 56881 4285
0 4287 7 1 2 57731 4286
0 4288 5 1 1 4287
0 4289 7 1 2 4276 4288
0 4290 5 1 1 4289
0 4291 7 1 2 48391 4290
0 4292 5 1 1 4291
0 4293 7 5 2 50933 51963
0 4294 5 2 1 57739
0 4295 7 1 2 46894 54654
0 4296 7 1 2 57450 4295
0 4297 7 1 2 57740 4296
0 4298 7 1 2 56769 4297
0 4299 5 1 1 4298
0 4300 7 1 2 4292 4299
0 4301 5 1 1 4300
0 4302 7 1 2 44722 4301
0 4303 5 1 1 4302
0 4304 7 1 2 4177 4303
0 4305 5 1 1 4304
0 4306 7 1 2 44616 4305
0 4307 5 1 1 4306
0 4308 7 8 2 46613 47866
0 4309 7 1 2 56497 57746
0 4310 5 2 1 4309
0 4311 7 1 2 55723 57754
0 4312 5 1 1 4311
0 4313 7 1 2 51394 4312
0 4314 5 1 1 4313
0 4315 7 1 2 51658 53344
0 4316 7 1 2 57581 4315
0 4317 5 1 1 4316
0 4318 7 1 2 55724 4317
0 4319 5 1 1 4318
0 4320 7 1 2 51497 4319
0 4321 5 1 1 4320
0 4322 7 1 2 4314 4321
0 4323 5 1 1 4322
0 4324 7 1 2 47501 4323
0 4325 5 1 1 4324
0 4326 7 1 2 51584 57719
0 4327 5 1 1 4326
0 4328 7 2 2 48539 56963
0 4329 5 1 1 57756
0 4330 7 1 2 55537 57757
0 4331 5 1 1 4330
0 4332 7 1 2 4327 4331
0 4333 5 1 1 4332
0 4334 7 1 2 46411 4333
0 4335 5 1 1 4334
0 4336 7 1 2 4325 4335
0 4337 5 1 1 4336
0 4338 7 1 2 48392 4337
0 4339 5 1 1 4338
0 4340 7 7 2 42994 45038
0 4341 7 7 2 44157 47867
0 4342 7 1 2 56498 57765
0 4343 5 1 1 4342
0 4344 7 1 2 49193 51585
0 4345 5 1 1 4344
0 4346 7 1 2 4343 4345
0 4347 5 1 1 4346
0 4348 7 1 2 43220 4347
0 4349 5 1 1 4348
0 4350 7 6 2 43514 44158
0 4351 7 14 2 44531 48759
0 4352 7 1 2 57772 57778
0 4353 5 2 1 4352
0 4354 7 1 2 4349 57792
0 4355 5 2 1 4354
0 4356 7 1 2 50594 57794
0 4357 5 1 1 4356
0 4358 7 6 2 46895 55417
0 4359 5 1 1 57796
0 4360 7 1 2 51629 4359
0 4361 5 3 1 4360
0 4362 7 1 2 49678 57802
0 4363 5 1 1 4362
0 4364 7 1 2 4357 4363
0 4365 5 1 1 4364
0 4366 7 1 2 57758 4365
0 4367 5 1 1 4366
0 4368 7 1 2 4339 4367
0 4369 5 1 1 4368
0 4370 7 3 2 44389 48074
0 4371 7 1 2 55217 57805
0 4372 7 1 2 55467 4371
0 4373 7 1 2 4369 4372
0 4374 5 1 1 4373
0 4375 7 1 2 42130 4374
0 4376 7 1 2 4307 4375
0 4377 5 1 1 4376
0 4378 7 1 2 3981 4377
0 4379 5 1 1 4378
0 4380 7 1 2 45961 4379
0 4381 5 1 1 4380
0 4382 7 2 2 44390 53664
0 4383 7 1 2 42995 50817
0 4384 5 5 1 4383
0 4385 7 3 2 50893 57810
0 4386 5 2 1 57815
0 4387 7 1 2 56307 57818
0 4388 5 2 1 4387
0 4389 7 1 2 50047 56004
0 4390 5 1 1 4389
0 4391 7 1 2 57820 4390
0 4392 5 1 1 4391
0 4393 7 1 2 42701 4392
0 4394 5 1 1 4393
0 4395 7 2 2 50048 53417
0 4396 5 2 1 57822
0 4397 7 3 2 49948 50976
0 4398 5 2 1 57826
0 4399 7 1 2 49327 57827
0 4400 5 2 1 4399
0 4401 7 1 2 57824 57831
0 4402 5 1 1 4401
0 4403 7 1 2 45181 4402
0 4404 5 1 1 4403
0 4405 7 9 2 49328 50977
0 4406 5 1 1 57833
0 4407 7 1 2 48540 55558
0 4408 7 1 2 57834 4407
0 4409 5 1 1 4408
0 4410 7 1 2 4404 4409
0 4411 5 1 1 4410
0 4412 7 1 2 43844 4411
0 4413 5 1 1 4412
0 4414 7 1 2 4394 4413
0 4415 5 1 1 4414
0 4416 7 1 2 48760 4415
0 4417 5 1 1 4416
0 4418 7 1 2 48976 52229
0 4419 5 1 1 4418
0 4420 7 1 2 47203 52924
0 4421 5 2 1 4420
0 4422 7 1 2 54319 57842
0 4423 7 1 2 4419 4422
0 4424 5 1 1 4423
0 4425 7 1 2 4417 4424
0 4426 5 1 1 4425
0 4427 7 1 2 50678 4426
0 4428 5 1 1 4427
0 4429 7 1 2 56835 57725
0 4430 5 1 1 4429
0 4431 7 4 2 43845 44532
0 4432 7 2 2 47949 57844
0 4433 7 1 2 48075 50049
0 4434 7 1 2 54529 4433
0 4435 7 1 2 57848 4434
0 4436 5 1 1 4435
0 4437 7 1 2 49143 50349
0 4438 7 7 2 47069 44723
0 4439 5 1 1 57850
0 4440 7 1 2 52021 57851
0 4441 7 1 2 4437 4440
0 4442 5 1 1 4441
0 4443 7 1 2 4436 4442
0 4444 5 1 1 4443
0 4445 7 1 2 52888 4444
0 4446 5 1 1 4445
0 4447 7 1 2 4430 4446
0 4448 7 1 2 4428 4447
0 4449 5 1 1 4448
0 4450 7 1 2 48393 4449
0 4451 5 1 1 4450
0 4452 7 2 2 45039 56743
0 4453 5 1 1 57857
0 4454 7 1 2 57076 4453
0 4455 5 1 1 4454
0 4456 7 1 2 57042 4455
0 4457 5 1 1 4456
0 4458 7 3 2 49102 51517
0 4459 5 2 1 57859
0 4460 7 6 2 47204 47868
0 4461 7 2 2 56941 57864
0 4462 7 1 2 45040 57870
0 4463 7 1 2 57862 4462
0 4464 5 1 1 4463
0 4465 7 1 2 4457 4464
0 4466 5 1 1 4465
0 4467 7 1 2 43991 4466
0 4468 5 1 1 4467
0 4469 7 1 2 50221 57045
0 4470 5 1 1 4469
0 4471 7 1 2 4468 4470
0 4472 5 1 1 4471
0 4473 7 1 2 42996 4472
0 4474 5 1 1 4473
0 4475 7 6 2 43992 44533
0 4476 7 1 2 42702 55647
0 4477 7 1 2 57872 4476
0 4478 7 1 2 56681 4477
0 4479 7 1 2 51449 4478
0 4480 5 1 1 4479
0 4481 7 1 2 4474 4480
0 4482 7 1 2 4451 4481
0 4483 5 1 1 4482
0 4484 7 1 2 57808 4483
0 4485 5 1 1 4484
0 4486 7 1 2 43993 52345
0 4487 5 2 1 4486
0 4488 7 1 2 57487 57878
0 4489 5 4 1 4488
0 4490 7 1 2 55884 57880
0 4491 5 1 1 4490
0 4492 7 4 2 47721 57604
0 4493 7 1 2 57600 57884
0 4494 5 1 1 4493
0 4495 7 1 2 4491 4494
0 4496 5 1 1 4495
0 4497 7 1 2 52022 4496
0 4498 5 1 1 4497
0 4499 7 5 2 42997 55885
0 4500 7 1 2 56810 57888
0 4501 5 1 1 4500
0 4502 7 1 2 4498 4501
0 4503 5 1 1 4502
0 4504 7 1 2 50498 54655
0 4505 7 1 2 4503 4504
0 4506 5 1 1 4505
0 4507 7 2 2 46412 54460
0 4508 7 2 2 57065 57893
0 4509 7 1 2 47070 57189
0 4510 5 1 1 4509
0 4511 7 5 2 46614 47205
0 4512 7 1 2 55094 57897
0 4513 7 1 2 53822 4512
0 4514 5 1 1 4513
0 4515 7 1 2 4510 4514
0 4516 5 1 1 4515
0 4517 7 1 2 57895 4516
0 4518 5 1 1 4517
0 4519 7 2 2 50656 54450
0 4520 7 1 2 56453 56336
0 4521 7 1 2 57902 4520
0 4522 7 1 2 57601 4521
0 4523 5 1 1 4522
0 4524 7 1 2 4518 4523
0 4525 7 1 2 4506 4524
0 4526 5 1 1 4525
0 4527 7 1 2 45041 4526
0 4528 5 1 1 4527
0 4529 7 1 2 56488 56830
0 4530 5 1 1 4529
0 4531 7 23 2 44391 47950
0 4532 7 4 2 56460 57904
0 4533 7 1 2 57037 57927
0 4534 5 1 1 4533
0 4535 7 1 2 4530 4534
0 4536 5 1 1 4535
0 4537 7 3 2 46796 48989
0 4538 7 1 2 4536 57931
0 4539 5 1 1 4538
0 4540 7 1 2 50535 54410
0 4541 7 16 2 44617 48761
0 4542 7 4 2 47206 44392
0 4543 7 1 2 54421 57950
0 4544 7 1 2 57934 4543
0 4545 7 1 2 4540 4544
0 4546 5 1 1 4545
0 4547 7 1 2 4539 4546
0 4548 5 1 1 4547
0 4549 7 1 2 55559 4548
0 4550 5 1 1 4549
0 4551 7 2 2 49736 50736
0 4552 5 1 1 57954
0 4553 7 1 2 53951 57955
0 4554 5 2 1 4553
0 4555 7 1 2 3711 57956
0 4556 5 1 1 4555
0 4557 7 1 2 45386 4556
0 4558 5 1 1 4557
0 4559 7 1 2 47207 52827
0 4560 5 1 1 4559
0 4561 7 1 2 4558 4560
0 4562 5 1 1 4561
0 4563 7 1 2 46149 4562
0 4564 5 1 1 4563
0 4565 7 1 2 53455 56983
0 4566 5 1 1 4565
0 4567 7 1 2 4564 4566
0 4568 5 1 1 4567
0 4569 7 1 2 57067 4568
0 4570 5 1 1 4569
0 4571 7 1 2 4550 4570
0 4572 5 1 1 4571
0 4573 7 1 2 46413 4572
0 4574 5 1 1 4573
0 4575 7 2 2 55468 56567
0 4576 7 4 2 47502 44393
0 4577 7 1 2 49528 57960
0 4578 7 1 2 57958 4577
0 4579 5 1 1 4578
0 4580 7 5 2 47503 47722
0 4581 7 4 2 46797 57964
0 4582 7 2 2 49529 57969
0 4583 5 1 1 57973
0 4584 7 1 2 50125 55886
0 4585 7 1 2 54347 4584
0 4586 5 1 1 4585
0 4587 7 1 2 4583 4586
0 4588 5 1 1 4587
0 4589 7 9 2 47208 44724
0 4590 7 1 2 54090 54495
0 4591 7 1 2 57975 4590
0 4592 7 1 2 4588 4591
0 4593 5 1 1 4592
0 4594 7 1 2 4579 4593
0 4595 5 1 1 4594
0 4596 7 1 2 45182 4595
0 4597 5 1 1 4596
0 4598 7 1 2 52023 57068
0 4599 7 1 2 57338 4598
0 4600 5 1 1 4599
0 4601 7 1 2 4597 4600
0 4602 7 1 2 4574 4601
0 4603 5 1 1 4602
0 4604 7 1 2 48394 4603
0 4605 5 1 1 4604
0 4606 7 1 2 52024 57241
0 4607 7 1 2 57155 4606
0 4608 7 1 2 57896 4607
0 4609 5 1 1 4608
0 4610 7 1 2 4605 4609
0 4611 7 1 2 4528 4610
0 4612 5 1 1 4611
0 4613 7 1 2 53572 4612
0 4614 5 1 1 4613
0 4615 7 1 2 4485 4614
0 4616 5 1 1 4615
0 4617 7 1 2 44884 4616
0 4618 5 1 1 4617
0 4619 7 1 2 42703 56837
0 4620 5 1 1 4619
0 4621 7 1 2 49246 4620
0 4622 5 1 1 4621
0 4623 7 1 2 46414 4622
0 4624 5 1 1 4623
0 4625 7 1 2 3884 4624
0 4626 5 1 1 4625
0 4627 7 1 2 43846 4626
0 4628 5 1 1 4627
0 4629 7 1 2 52941 57307
0 4630 5 1 1 4629
0 4631 7 1 2 4628 4630
0 4632 5 1 1 4631
0 4633 7 1 2 50679 4632
0 4634 5 1 1 4633
0 4635 7 2 2 47504 54947
0 4636 7 1 2 47869 57984
0 4637 7 1 2 56985 4636
0 4638 5 1 1 4637
0 4639 7 1 2 4634 4638
0 4640 5 1 1 4639
0 4641 7 1 2 53665 4640
0 4642 5 1 1 4641
0 4643 7 10 2 45387 50050
0 4644 5 5 1 57986
0 4645 7 1 2 57987 57959
0 4646 5 1 1 4645
0 4647 7 5 2 47209 44534
0 4648 7 1 2 54411 58001
0 4649 7 1 2 57022 4648
0 4650 5 1 1 4649
0 4651 7 1 2 4646 4650
0 4652 5 1 1 4651
0 4653 7 1 2 49264 4652
0 4654 5 1 1 4653
0 4655 7 2 2 50499 56831
0 4656 7 7 2 47505 44535
0 4657 7 1 2 45388 55407
0 4658 7 1 2 58008 4657
0 4659 7 1 2 58006 4658
0 4660 5 1 1 4659
0 4661 7 1 2 4654 4660
0 4662 5 1 1 4661
0 4663 7 1 2 50978 53573
0 4664 7 1 2 4662 4663
0 4665 5 1 1 4664
0 4666 7 1 2 4642 4665
0 4667 5 1 1 4666
0 4668 7 1 2 44394 4667
0 4669 5 1 1 4668
0 4670 7 2 2 53574 57623
0 4671 7 10 2 44618 45389
0 4672 5 1 1 58017
0 4673 7 2 2 57700 58018
0 4674 7 1 2 56838 57976
0 4675 7 1 2 58027 4674
0 4676 7 1 2 58015 4675
0 4677 5 1 1 4676
0 4678 7 1 2 4669 4677
0 4679 5 1 1 4678
0 4680 7 1 2 45183 4679
0 4681 5 1 1 4680
0 4682 7 2 2 43847 47951
0 4683 7 1 2 56141 58029
0 4684 7 2 2 51701 4683
0 4685 7 1 2 56138 58031
0 4686 5 1 1 4685
0 4687 7 1 2 54948 56248
0 4688 7 1 2 55947 4687
0 4689 7 1 2 56711 4688
0 4690 5 1 1 4689
0 4691 7 1 2 4686 4690
0 4692 5 1 1 4691
0 4693 7 1 2 45671 4692
0 4694 5 1 1 4693
0 4695 7 3 2 46150 49907
0 4696 7 2 2 53556 58033
0 4697 7 5 2 47210 56701
0 4698 7 1 2 55948 58038
0 4699 7 1 2 58036 4698
0 4700 5 1 1 4699
0 4701 7 1 2 4694 4700
0 4702 5 1 1 4701
0 4703 7 1 2 43430 4702
0 4704 5 1 1 4703
0 4705 7 2 2 52776 54207
0 4706 7 1 2 46798 58043
0 4707 7 1 2 58032 4706
0 4708 5 1 1 4707
0 4709 7 1 2 4704 4708
0 4710 5 1 1 4709
0 4711 7 1 2 44395 54656
0 4712 7 1 2 4710 4711
0 4713 5 1 1 4712
0 4714 7 1 2 4681 4713
0 4715 5 1 1 4714
0 4716 7 1 2 49644 4715
0 4717 5 1 1 4716
0 4718 7 1 2 42462 4717
0 4719 7 1 2 4618 4718
0 4720 5 1 1 4719
0 4721 7 1 2 45509 4720
0 4722 7 1 2 4381 4721
0 4723 5 1 1 4722
0 4724 7 7 2 44536 53575
0 4725 7 2 2 46615 55601
0 4726 5 1 1 58052
0 4727 7 1 2 55925 4726
0 4728 5 3 1 4727
0 4729 7 1 2 57228 58054
0 4730 5 1 1 4729
0 4731 7 13 2 43221 43431
0 4732 7 3 2 44396 58057
0 4733 5 1 1 58070
0 4734 7 9 2 46616 46799
0 4735 7 3 2 47723 58073
0 4736 7 1 2 42704 58082
0 4737 5 1 1 4736
0 4738 7 1 2 4733 4737
0 4739 5 1 1 4738
0 4740 7 1 2 57441 4739
0 4741 5 1 1 4740
0 4742 7 1 2 4730 4741
0 4743 5 1 1 4742
0 4744 7 1 2 50536 4743
0 4745 5 1 1 4744
0 4746 7 1 2 57467 58071
0 4747 5 1 1 4746
0 4748 7 1 2 4745 4747
0 4749 5 1 1 4748
0 4750 7 1 2 45510 4749
0 4751 5 1 1 4750
0 4752 7 8 2 44397 54740
0 4753 5 1 1 58085
0 4754 7 7 2 43222 44725
0 4755 7 1 2 54156 58093
0 4756 5 1 1 4755
0 4757 7 1 2 3967 4756
0 4758 5 1 1 4757
0 4759 7 1 2 46151 4758
0 4760 5 1 1 4759
0 4761 7 3 2 43223 57177
0 4762 7 1 2 57193 58100
0 4763 5 1 1 4762
0 4764 7 1 2 4760 4763
0 4765 5 1 1 4764
0 4766 7 1 2 58086 4765
0 4767 5 1 1 4766
0 4768 7 1 2 4751 4767
0 4769 5 1 1 4768
0 4770 7 1 2 58045 4769
0 4771 5 1 1 4770
0 4772 7 6 2 45511 53666
0 4773 5 1 1 58103
0 4774 7 8 2 45672 46800
0 4775 5 1 1 58109
0 4776 7 5 2 41969 46896
0 4777 7 5 2 58110 58117
0 4778 5 1 1 58122
0 4779 7 1 2 4773 4778
0 4780 5 16 1 4779
0 4781 7 4 2 44398 58127
0 4782 7 2 2 55812 57575
0 4783 7 1 2 57234 58147
0 4784 7 1 2 58143 4783
0 4785 5 1 1 4784
0 4786 7 1 2 4771 4785
0 4787 5 1 1 4786
0 4788 7 1 2 45962 4787
0 4789 5 1 1 4788
0 4790 7 2 2 50537 54928
0 4791 5 2 1 58149
0 4792 7 1 2 1696 58151
0 4793 5 1 1 4792
0 4794 7 1 2 46152 4793
0 4795 5 1 1 4794
0 4796 7 1 2 57178 57242
0 4797 5 1 1 4796
0 4798 7 1 2 4795 4797
0 4799 5 1 1 4798
0 4800 7 10 2 44399 54754
0 4801 7 2 2 53576 54422
0 4802 7 1 2 42463 58163
0 4803 7 1 2 58153 4802
0 4804 7 1 2 4799 4803
0 4805 5 1 1 4804
0 4806 7 1 2 4789 4805
0 4807 5 1 1 4806
0 4808 7 1 2 44885 4807
0 4809 5 1 1 4808
0 4810 7 5 2 54755 57419
0 4811 5 1 1 58165
0 4812 7 36 2 45512 46801
0 4813 5 2 1 58170
0 4814 7 2 2 55956 58171
0 4815 7 1 2 46617 58208
0 4816 5 1 1 4815
0 4817 7 1 2 4811 4816
0 4818 5 1 1 4817
0 4819 7 1 2 42131 4818
0 4820 5 1 1 4819
0 4821 7 3 2 45673 54756
0 4822 7 1 2 57269 58210
0 4823 5 1 1 4822
0 4824 7 1 2 4820 4823
0 4825 5 1 1 4824
0 4826 7 2 2 53194 54912
0 4827 5 1 1 58213
0 4828 7 5 2 44400 44726
0 4829 7 2 2 45184 58215
0 4830 7 1 2 47367 58220
0 4831 7 1 2 58214 4830
0 4832 7 1 2 4825 4831
0 4833 5 1 1 4832
0 4834 7 1 2 4809 4833
0 4835 5 1 1 4834
0 4836 7 1 2 45042 4835
0 4837 5 1 1 4836
0 4838 7 10 2 42464 44886
0 4839 5 1 1 58222
0 4840 7 2 2 838 4839
0 4841 5 16 1 58232
0 4842 7 3 2 58128 58234
0 4843 7 1 2 48541 57457
0 4844 7 1 2 58250 4843
0 4845 5 1 1 4844
0 4846 7 12 2 45513 45963
0 4847 7 2 2 55970 58253
0 4848 7 6 2 46897 43994
0 4849 7 14 2 43224 46802
0 4850 7 1 2 49814 58273
0 4851 7 1 2 58267 4850
0 4852 7 1 2 58265 4851
0 4853 5 1 1 4852
0 4854 7 1 2 4845 4853
0 4855 5 1 1 4854
0 4856 7 10 2 47870 44727
0 4857 7 2 2 52729 58287
0 4858 7 1 2 54091 58297
0 4859 7 1 2 4855 4858
0 4860 5 1 1 4859
0 4861 7 1 2 4837 4860
0 4862 5 1 1 4861
0 4863 7 1 2 46415 4862
0 4864 5 1 1 4863
0 4865 7 2 2 44537 56273
0 4866 7 10 2 43225 43848
0 4867 5 1 1 58301
0 4868 7 4 2 44887 58302
0 4869 7 2 2 43995 54370
0 4870 7 1 2 58311 58315
0 4871 7 1 2 58299 4870
0 4872 5 1 1 4871
0 4873 7 4 2 47211 57008
0 4874 7 1 2 55513 58317
0 4875 7 1 2 58251 4874
0 4876 5 1 1 4875
0 4877 7 1 2 4872 4876
0 4878 5 1 1 4877
0 4879 7 1 2 52499 58221
0 4880 7 1 2 4878 4879
0 4881 5 1 1 4880
0 4882 7 1 2 4864 4881
0 4883 5 1 1 4882
0 4884 7 1 2 44619 4883
0 4885 5 1 1 4884
0 4886 7 2 2 52889 58129
0 4887 7 4 2 54371 56775
0 4888 7 1 2 56454 58323
0 4889 7 1 2 56166 4888
0 4890 7 1 2 58321 4889
0 4891 5 1 1 4890
0 4892 7 1 2 4885 4891
0 4893 5 1 1 4892
0 4894 7 1 2 49066 4893
0 4895 5 1 1 4894
0 4896 7 2 2 48220 55338
0 4897 5 1 1 58327
0 4898 7 1 2 46416 57116
0 4899 5 1 1 4898
0 4900 7 1 2 57060 4899
0 4901 5 1 1 4900
0 4902 7 1 2 58328 4901
0 4903 5 1 1 4902
0 4904 7 1 2 52663 56759
0 4905 5 1 1 4904
0 4906 7 1 2 57821 4905
0 4907 5 1 1 4906
0 4908 7 2 2 48762 4907
0 4909 5 1 1 58329
0 4910 7 1 2 54826 58330
0 4911 5 1 1 4910
0 4912 7 1 2 4903 4911
0 4913 5 1 1 4912
0 4914 7 1 2 47071 4913
0 4915 5 1 1 4914
0 4916 7 1 2 46153 57679
0 4917 5 1 1 4916
0 4918 7 1 2 47212 57671
0 4919 5 1 1 4918
0 4920 7 1 2 4917 4919
0 4921 5 1 1 4920
0 4922 7 1 2 45390 4921
0 4923 5 1 1 4922
0 4924 7 2 2 52742 57072
0 4925 7 1 2 46417 58331
0 4926 5 1 1 4925
0 4927 7 1 2 4923 4926
0 4928 5 1 1 4927
0 4929 7 1 2 53898 4928
0 4930 5 1 1 4929
0 4931 7 1 2 4915 4930
0 4932 5 1 1 4931
0 4933 7 1 2 45964 4932
0 4934 5 1 1 4933
0 4935 7 5 2 46154 49949
0 4936 5 2 1 58333
0 4937 7 11 2 44159 45391
0 4938 5 2 1 58340
0 4939 7 2 2 57658 58351
0 4940 5 9 1 58353
0 4941 7 1 2 43226 58354
0 4942 5 1 1 4941
0 4943 7 15 2 51198 4942
0 4944 7 3 2 46418 58364
0 4945 5 3 1 58379
0 4946 7 1 2 58338 58382
0 4947 5 1 1 4946
0 4948 7 1 2 53895 54113
0 4949 7 1 2 4947 4948
0 4950 5 1 1 4949
0 4951 7 1 2 4934 4950
0 4952 5 1 1 4951
0 4953 7 1 2 48395 4952
0 4954 5 1 1 4953
0 4955 7 3 2 43996 50183
0 4956 5 1 1 58385
0 4957 7 2 2 53521 54372
0 4958 5 1 1 58388
0 4959 7 1 2 58386 58389
0 4960 5 1 1 4959
0 4961 7 2 2 56308 57149
0 4962 7 1 2 53354 53847
0 4963 7 1 2 58390 4962
0 4964 5 1 1 4963
0 4965 7 1 2 4960 4964
0 4966 5 1 1 4965
0 4967 7 1 2 44160 4966
0 4968 5 1 1 4967
0 4969 7 10 2 45965 46618
0 4970 7 1 2 56337 58392
0 4971 7 1 2 55306 4970
0 4972 5 1 1 4971
0 4973 7 1 2 4968 4972
0 4974 5 1 1 4973
0 4975 7 1 2 52518 4974
0 4976 5 1 1 4975
0 4977 7 1 2 4954 4976
0 4978 5 1 1 4977
0 4979 7 1 2 4978 58164
0 4980 5 1 1 4979
0 4981 7 1 2 52154 53230
0 4982 5 1 1 4981
0 4983 7 1 2 832 4982
0 4984 5 1 1 4983
0 4985 7 1 2 52025 4984
0 4986 5 1 1 4985
0 4987 7 2 2 44888 53184
0 4988 7 3 2 43849 44728
0 4989 7 1 2 54983 58404
0 4990 7 1 2 58402 4989
0 4991 5 1 1 4990
0 4992 7 1 2 4986 4991
0 4993 5 1 1 4992
0 4994 7 1 2 50737 4993
0 4995 5 1 1 4994
0 4996 7 4 2 45966 54949
0 4997 7 1 2 52155 54929
0 4998 7 1 2 58407 4997
0 4999 5 1 1 4998
0 5000 7 1 2 4995 4999
0 5001 5 1 1 5000
0 5002 7 1 2 58046 5001
0 5003 5 1 1 5002
0 5004 7 1 2 53982 57235
0 5005 5 1 1 5004
0 5006 7 1 2 52156 55085
0 5007 5 1 1 5006
0 5008 7 1 2 5005 5007
0 5009 5 1 1 5008
0 5010 7 10 2 46419 47506
0 5011 5 4 1 58411
0 5012 7 4 2 46898 51895
0 5013 7 1 2 58412 58425
0 5014 7 1 2 5009 5013
0 5015 5 1 1 5014
0 5016 7 1 2 5003 5015
0 5017 5 1 1 5016
0 5018 7 1 2 50312 5017
0 5019 5 1 1 5018
0 5020 7 8 2 42465 46619
0 5021 7 1 2 58039 58429
0 5022 5 1 1 5021
0 5023 7 2 2 49892 57252
0 5024 5 1 1 58437
0 5025 7 1 2 5022 5024
0 5026 5 1 1 5025
0 5027 7 1 2 46420 5026
0 5028 5 1 1 5027
0 5029 7 1 2 56632 57336
0 5030 5 1 1 5029
0 5031 7 1 2 5028 5030
0 5032 5 1 1 5031
0 5033 7 1 2 45392 5032
0 5034 5 1 1 5033
0 5035 7 1 2 55034 57526
0 5036 5 1 1 5035
0 5037 7 1 2 5034 5036
0 5038 5 1 1 5037
0 5039 7 1 2 48221 5038
0 5040 5 1 1 5039
0 5041 7 1 2 43850 49908
0 5042 5 1 1 5041
0 5043 7 1 2 55352 5042
0 5044 5 1 1 5043
0 5045 7 1 2 49194 5044
0 5046 5 1 1 5045
0 5047 7 3 2 46421 57321
0 5048 5 1 1 58439
0 5049 7 1 2 52373 58440
0 5050 5 1 1 5049
0 5051 7 4 2 47368 49067
0 5052 5 5 1 58442
0 5053 7 2 2 49107 58446
0 5054 7 1 2 54107 58451
0 5055 5 1 1 5054
0 5056 7 1 2 5050 5055
0 5057 5 1 1 5056
0 5058 7 1 2 43227 5057
0 5059 5 1 1 5058
0 5060 7 1 2 5046 5059
0 5061 5 1 1 5060
0 5062 7 1 2 58223 5061
0 5063 5 1 1 5062
0 5064 7 1 2 5040 5063
0 5065 5 1 1 5064
0 5066 7 1 2 46155 5065
0 5067 5 1 1 5066
0 5068 7 2 2 42466 49909
0 5069 7 1 2 52932 58453
0 5070 5 1 1 5069
0 5071 7 1 2 4958 5070
0 5072 5 1 1 5071
0 5073 7 1 2 49195 5072
0 5074 5 1 1 5073
0 5075 7 3 2 43997 49144
0 5076 7 3 2 42467 57898
0 5077 7 1 2 58455 58458
0 5078 5 1 1 5077
0 5079 7 3 2 48763 49874
0 5080 5 3 1 58461
0 5081 7 1 2 47213 58464
0 5082 5 1 1 5081
0 5083 7 2 2 43228 5082
0 5084 5 2 1 58467
0 5085 7 3 2 45967 52052
0 5086 5 2 1 58471
0 5087 7 1 2 46156 58465
0 5088 5 2 1 5087
0 5089 7 1 2 58472 58476
0 5090 7 1 2 58468 5089
0 5091 5 1 1 5090
0 5092 7 1 2 5078 5091
0 5093 5 1 1 5092
0 5094 7 1 2 42998 5093
0 5095 5 1 1 5094
0 5096 7 1 2 5074 5095
0 5097 5 1 1 5096
0 5098 7 1 2 48542 5097
0 5099 5 1 1 5098
0 5100 7 5 2 44161 49893
0 5101 7 3 2 43851 48764
0 5102 5 2 1 58483
0 5103 7 2 2 58478 58484
0 5104 5 1 1 58488
0 5105 7 10 2 42468 47214
0 5106 7 1 2 57368 58490
0 5107 5 1 1 5106
0 5108 7 1 2 5104 5107
0 5109 5 1 1 5108
0 5110 7 1 2 54208 5109
0 5111 5 1 1 5110
0 5112 7 1 2 5099 5111
0 5113 5 1 1 5112
0 5114 7 1 2 44889 5113
0 5115 5 1 1 5114
0 5116 7 1 2 5067 5115
0 5117 5 1 1 5116
0 5118 7 1 2 47072 5117
0 5119 5 1 1 5118
0 5120 7 4 2 47215 49145
0 5121 5 2 1 58500
0 5122 7 3 2 42999 53724
0 5123 5 1 1 58506
0 5124 7 1 2 58501 58507
0 5125 5 1 1 5124
0 5126 7 1 2 46422 49196
0 5127 7 1 2 55697 5126
0 5128 5 1 1 5127
0 5129 7 1 2 5125 5128
0 5130 5 1 1 5129
0 5131 7 1 2 46620 5130
0 5132 5 1 1 5131
0 5133 7 2 2 52403 57341
0 5134 5 1 1 58509
0 5135 7 1 2 52235 58510
0 5136 5 1 1 5135
0 5137 7 1 2 5132 5136
0 5138 5 1 1 5137
0 5139 7 1 2 58403 5138
0 5140 5 1 1 5139
0 5141 7 1 2 5119 5140
0 5142 5 1 1 5141
0 5143 7 1 2 44729 5142
0 5144 5 1 1 5143
0 5145 7 1 2 53848 54930
0 5146 5 2 1 5145
0 5147 7 2 2 49197 53231
0 5148 7 1 2 43852 58513
0 5149 5 1 1 5148
0 5150 7 1 2 58511 5149
0 5151 5 1 1 5150
0 5152 7 1 2 44890 5151
0 5153 5 1 1 5152
0 5154 7 1 2 5153 4827
0 5155 5 1 1 5154
0 5156 7 1 2 49910 5155
0 5157 5 1 1 5156
0 5158 7 1 2 49601 57117
0 5159 7 1 2 54128 5158
0 5160 5 1 1 5159
0 5161 7 1 2 5157 5160
0 5162 5 1 1 5161
0 5163 7 1 2 44730 5162
0 5164 5 1 1 5163
0 5165 7 2 2 50912 57219
0 5166 5 1 1 58515
0 5167 7 1 2 54073 57009
0 5168 7 1 2 58516 5167
0 5169 5 1 1 5168
0 5170 7 1 2 5164 5169
0 5171 5 1 1 5170
0 5172 7 1 2 47369 5171
0 5173 5 1 1 5172
0 5174 7 4 2 45968 49950
0 5175 5 1 1 58517
0 5176 7 1 2 57050 58518
0 5177 5 1 1 5176
0 5178 7 1 2 50304 58459
0 5179 5 1 1 5178
0 5180 7 1 2 5177 5179
0 5181 5 1 1 5180
0 5182 7 1 2 48222 5181
0 5183 5 1 1 5182
0 5184 7 1 2 55146 58312
0 5185 5 1 1 5184
0 5186 7 1 2 5183 5185
0 5187 5 1 1 5186
0 5188 7 1 2 46157 5187
0 5189 5 1 1 5188
0 5190 7 2 2 54373 54723
0 5191 7 1 2 57308 58521
0 5192 5 1 1 5191
0 5193 7 1 2 5189 5192
0 5194 5 1 1 5193
0 5195 7 1 2 44731 5194
0 5196 5 1 1 5195
0 5197 7 2 2 50738 52026
0 5198 7 2 2 50913 58523
0 5199 7 1 2 51638 58525
0 5200 5 1 1 5199
0 5201 7 1 2 5196 5200
0 5202 5 1 1 5201
0 5203 7 1 2 47073 5202
0 5204 5 1 1 5203
0 5205 7 1 2 50914 53899
0 5206 7 1 2 57342 58405
0 5207 7 1 2 5205 5206
0 5208 5 1 1 5207
0 5209 7 1 2 5204 5208
0 5210 7 1 2 5173 5209
0 5211 5 1 1 5210
0 5212 7 1 2 45185 5211
0 5213 5 1 1 5212
0 5214 7 1 2 56012 58040
0 5215 7 5 2 46423 57207
0 5216 7 2 2 44891 55180
0 5217 7 1 2 58527 58532
0 5218 7 1 2 5214 5217
0 5219 5 1 1 5218
0 5220 7 1 2 5213 5219
0 5221 7 1 2 5144 5220
0 5222 5 1 1 5221
0 5223 7 1 2 58047 5222
0 5224 5 1 1 5223
0 5225 7 1 2 5019 5224
0 5226 5 1 1 5225
0 5227 7 1 2 45043 5226
0 5228 5 1 1 5227
0 5229 7 1 2 4980 5228
0 5230 5 1 1 5229
0 5231 7 1 2 44620 5230
0 5232 5 1 1 5231
0 5233 7 3 2 43998 56744
0 5234 5 2 1 58534
0 5235 7 1 2 51451 58537
0 5236 5 1 1 5235
0 5237 7 1 2 57759 5236
0 5238 5 1 1 5237
0 5239 7 3 2 43229 53539
0 5240 5 2 1 58539
0 5241 7 1 2 49265 58540
0 5242 5 1 1 5241
0 5243 7 1 2 5238 5242
0 5244 5 1 1 5243
0 5245 7 1 2 57043 5244
0 5246 5 1 1 5245
0 5247 7 1 2 48396 57732
0 5248 5 1 1 5247
0 5249 7 1 2 43000 56677
0 5250 5 1 1 5249
0 5251 7 1 2 5248 5250
0 5252 5 1 1 5251
0 5253 7 1 2 57871 5252
0 5254 5 1 1 5253
0 5255 7 1 2 5246 5254
0 5256 5 1 1 5255
0 5257 7 1 2 53301 5256
0 5258 5 1 1 5257
0 5259 7 4 2 50051 52890
0 5260 5 5 1 58544
0 5261 7 1 2 48990 50739
0 5262 5 7 1 5261
0 5263 7 2 2 58548 58553
0 5264 7 10 2 46424 45186
0 5265 5 9 1 58562
0 5266 7 1 2 48765 58572
0 5267 5 1 1 5266
0 5268 7 1 2 57570 5267
0 5269 5 1 1 5268
0 5270 7 1 2 58560 5269
0 5271 5 1 1 5270
0 5272 7 1 2 47216 5271
0 5273 5 1 1 5272
0 5274 7 2 2 49951 50538
0 5275 5 3 1 58581
0 5276 7 1 2 57957 58583
0 5277 5 1 1 5276
0 5278 7 1 2 53736 5277
0 5279 5 1 1 5278
0 5280 7 1 2 5273 5279
0 5281 5 1 1 5280
0 5282 7 1 2 52428 5281
0 5283 5 1 1 5282
0 5284 7 7 2 49146 49911
0 5285 5 1 1 58586
0 5286 7 1 2 50315 54931
0 5287 7 1 2 58587 5286
0 5288 5 1 1 5287
0 5289 7 1 2 5283 5288
0 5290 5 1 1 5289
0 5291 7 1 2 46158 5290
0 5292 5 1 1 5291
0 5293 7 3 2 45393 52500
0 5294 5 1 1 58593
0 5295 7 1 2 53096 54337
0 5296 7 1 2 58594 5295
0 5297 5 1 1 5296
0 5298 7 1 2 5292 5297
0 5299 5 1 1 5298
0 5300 7 1 2 53316 54513
0 5301 7 1 2 5299 5300
0 5302 5 1 1 5301
0 5303 7 1 2 5258 5302
0 5304 5 1 1 5303
0 5305 7 1 2 52795 58235
0 5306 7 1 2 5304 5305
0 5307 5 1 1 5306
0 5308 7 1 2 57070 58549
0 5309 5 1 1 5308
0 5310 7 1 2 43853 5309
0 5311 5 1 1 5310
0 5312 7 1 2 52915 57118
0 5313 5 1 1 5312
0 5314 7 1 2 5311 5313
0 5315 5 1 1 5314
0 5316 7 1 2 48397 5315
0 5317 5 1 1 5316
0 5318 7 1 2 52256 52952
0 5319 5 1 1 5318
0 5320 7 1 2 5317 5319
0 5321 5 1 1 5320
0 5322 7 1 2 44892 5321
0 5323 5 1 1 5322
0 5324 7 5 2 46425 53962
0 5325 5 2 1 58596
0 5326 7 2 2 49645 56737
0 5327 5 1 1 58603
0 5328 7 1 2 58597 58604
0 5329 5 1 1 5328
0 5330 7 1 2 5323 5329
0 5331 5 1 1 5330
0 5332 7 1 2 42469 5331
0 5333 5 1 1 5332
0 5334 7 2 2 51428 56745
0 5335 5 1 1 58605
0 5336 7 1 2 46426 58606
0 5337 5 1 1 5336
0 5338 7 8 2 43001 47507
0 5339 5 1 1 58607
0 5340 7 2 2 48957 58608
0 5341 5 2 1 58615
0 5342 7 1 2 5337 58617
0 5343 5 1 1 5342
0 5344 7 2 2 54620 55015
0 5345 5 3 1 58619
0 5346 7 1 2 5343 58620
0 5347 5 1 1 5346
0 5348 7 1 2 5333 5347
0 5349 5 1 1 5348
0 5350 7 1 2 43691 5349
0 5351 5 1 1 5350
0 5352 7 6 2 45969 43999
0 5353 7 1 2 43854 49646
0 5354 7 1 2 58624 5353
0 5355 5 1 1 5354
0 5356 7 8 2 44893 49855
0 5357 5 1 1 58630
0 5358 7 1 2 58491 58631
0 5359 5 1 1 5358
0 5360 7 1 2 5355 5359
0 5361 5 1 1 5360
0 5362 7 1 2 43002 5361
0 5363 5 1 1 5362
0 5364 7 2 2 45970 53086
0 5365 7 1 2 48223 50519
0 5366 7 1 2 58638 5365
0 5367 5 1 1 5366
0 5368 7 1 2 42470 53546
0 5369 7 1 2 54261 5368
0 5370 5 1 1 5369
0 5371 7 1 2 5367 5370
0 5372 7 1 2 5363 5371
0 5373 5 1 1 5372
0 5374 7 1 2 43692 5373
0 5375 5 1 1 5374
0 5376 7 1 2 42471 49647
0 5377 7 1 2 54634 5376
0 5378 5 1 1 5377
0 5379 7 1 2 5375 5378
0 5380 5 1 1 5379
0 5381 7 1 2 50818 5380
0 5382 5 1 1 5381
0 5383 7 1 2 52967 55560
0 5384 5 1 1 5383
0 5385 7 1 2 52664 53006
0 5386 5 1 1 5385
0 5387 7 1 2 5384 5386
0 5388 5 1 1 5387
0 5389 7 5 2 42472 45187
0 5390 5 1 1 58640
0 5391 7 1 2 53900 58641
0 5392 7 1 2 5388 5391
0 5393 5 1 1 5392
0 5394 7 1 2 5382 5393
0 5395 5 1 1 5394
0 5396 7 1 2 48766 5395
0 5397 5 1 1 5396
0 5398 7 1 2 5351 5397
0 5399 5 1 1 5398
0 5400 7 1 2 42705 5399
0 5401 5 1 1 5400
0 5402 7 3 2 52575 55498
0 5403 5 1 1 58645
0 5404 7 3 2 45188 58646
0 5405 5 3 1 58648
0 5406 7 2 2 53963 58632
0 5407 5 1 1 58654
0 5408 7 1 2 58651 5407
0 5409 5 1 1 5408
0 5410 7 1 2 43003 5409
0 5411 5 1 1 5410
0 5412 7 3 2 53087 58633
0 5413 5 1 1 58656
0 5414 7 1 2 44000 58657
0 5415 5 1 1 5414
0 5416 7 1 2 5411 5415
0 5417 5 1 1 5416
0 5418 7 1 2 55561 5417
0 5419 5 1 1 5418
0 5420 7 1 2 44001 51876
0 5421 5 3 1 5420
0 5422 7 1 2 57832 58659
0 5423 5 1 1 5422
0 5424 7 1 2 51373 53108
0 5425 7 1 2 5423 5424
0 5426 5 1 1 5425
0 5427 7 1 2 5419 5426
0 5428 5 1 1 5427
0 5429 7 1 2 48767 5428
0 5430 5 1 1 5429
0 5431 7 5 2 49912 56885
0 5432 5 1 1 58662
0 5433 7 1 2 3919 5432
0 5434 5 1 1 5433
0 5435 7 1 2 53055 56716
0 5436 7 1 2 5434 5435
0 5437 5 1 1 5436
0 5438 7 1 2 5430 5437
0 5439 5 1 1 5438
0 5440 7 1 2 51127 5439
0 5441 5 1 1 5440
0 5442 7 1 2 5401 5441
0 5443 5 1 1 5442
0 5444 7 1 2 53302 53176
0 5445 7 1 2 5443 5444
0 5446 5 1 1 5445
0 5447 7 1 2 5307 5446
0 5448 7 1 2 5232 5447
0 5449 5 1 1 5448
0 5450 7 1 2 58087 5449
0 5451 5 1 1 5450
0 5452 7 2 2 48224 56548
0 5453 7 6 2 47871 53577
0 5454 7 3 2 49068 56707
0 5455 7 1 2 58669 58675
0 5456 5 1 1 5455
0 5457 7 3 2 42132 55178
0 5458 5 4 1 58678
0 5459 7 1 2 43515 58679
0 5460 5 1 1 5459
0 5461 7 1 2 5456 5460
0 5462 5 1 1 5461
0 5463 7 1 2 44401 5462
0 5464 5 1 1 5463
0 5465 7 6 2 45674 57624
0 5466 5 1 1 58685
0 5467 7 1 2 46899 58686
0 5468 7 1 2 58456 5467
0 5469 5 1 1 5468
0 5470 7 1 2 5464 5469
0 5471 5 1 1 5470
0 5472 7 1 2 58667 5471
0 5473 5 1 1 5472
0 5474 7 5 2 50500 53983
0 5475 7 3 2 43516 56416
0 5476 5 3 1 58696
0 5477 7 3 2 46900 44162
0 5478 7 2 2 57625 58702
0 5479 5 1 1 58705
0 5480 7 1 2 58699 5479
0 5481 5 2 1 5480
0 5482 7 1 2 42133 58707
0 5483 5 1 1 5482
0 5484 7 20 2 44538 55971
0 5485 7 1 2 57773 58709
0 5486 5 1 1 5485
0 5487 7 1 2 5483 5486
0 5488 5 1 1 5487
0 5489 7 1 2 45394 5488
0 5490 5 1 1 5489
0 5491 7 5 2 42134 56417
0 5492 5 1 1 58729
0 5493 7 1 2 57490 58730
0 5494 5 1 1 5493
0 5495 7 1 2 5490 5494
0 5496 5 1 1 5495
0 5497 7 1 2 58691 5496
0 5498 5 1 1 5497
0 5499 7 1 2 5473 5498
0 5500 5 1 1 5499
0 5501 7 1 2 46621 5500
0 5502 5 1 1 5501
0 5503 7 8 2 44539 48225
0 5504 7 2 2 56549 58734
0 5505 5 1 1 58742
0 5506 7 2 2 50376 50705
0 5507 5 1 1 58744
0 5508 7 1 2 5505 5507
0 5509 5 5 1 5508
0 5510 7 4 2 44402 52777
0 5511 7 2 2 58746 58751
0 5512 5 1 1 58755
0 5513 7 1 2 53984 56489
0 5514 5 1 1 5513
0 5515 7 1 2 56418 58668
0 5516 5 1 1 5515
0 5517 7 1 2 5514 5516
0 5518 5 1 1 5517
0 5519 7 1 2 43230 53578
0 5520 7 1 2 5518 5519
0 5521 5 1 1 5520
0 5522 7 1 2 5512 5521
0 5523 5 1 1 5522
0 5524 7 1 2 49147 5523
0 5525 5 1 1 5524
0 5526 7 1 2 5502 5525
0 5527 5 1 1 5526
0 5528 7 1 2 48543 5527
0 5529 5 1 1 5528
0 5530 7 1 2 57720 58756
0 5531 5 1 1 5530
0 5532 7 1 2 5529 5531
0 5533 5 1 1 5532
0 5534 7 1 2 46803 5533
0 5535 5 1 1 5534
0 5536 7 1 2 56968 58692
0 5537 5 1 1 5536
0 5538 7 1 2 55651 57420
0 5539 7 1 2 56550 5538
0 5540 5 1 1 5539
0 5541 7 1 2 5537 5540
0 5542 5 1 1 5541
0 5543 7 1 2 45675 5542
0 5544 5 1 1 5543
0 5545 7 2 2 45971 53557
0 5546 7 1 2 54441 58757
0 5547 5 1 1 5546
0 5548 7 1 2 5544 5547
0 5549 5 2 1 5548
0 5550 7 1 2 50052 58759
0 5551 5 1 1 5550
0 5552 7 3 2 46901 58747
0 5553 7 1 2 45676 50740
0 5554 7 1 2 58761 5553
0 5555 5 1 1 5554
0 5556 7 1 2 5551 5555
0 5557 5 1 1 5556
0 5558 7 1 2 48544 5557
0 5559 5 1 1 5558
0 5560 7 5 2 46902 49952
0 5561 5 1 1 58764
0 5562 7 2 2 56072 58765
0 5563 7 4 2 44540 50501
0 5564 7 2 2 51374 58771
0 5565 7 1 2 58769 58775
0 5566 5 1 1 5565
0 5567 7 1 2 57721 58762
0 5568 5 1 1 5567
0 5569 7 2 2 43517 58479
0 5570 7 1 2 58777 58776
0 5571 5 1 1 5570
0 5572 7 1 2 5568 5571
0 5573 5 1 1 5572
0 5574 7 1 2 45677 5573
0 5575 5 1 1 5574
0 5576 7 1 2 5566 5575
0 5577 7 1 2 5559 5576
0 5578 5 1 1 5577
0 5579 7 1 2 55887 5578
0 5580 5 1 1 5579
0 5581 7 1 2 5535 5580
0 5582 5 1 1 5581
0 5583 7 1 2 46427 5582
0 5584 5 1 1 5583
0 5585 7 1 2 56098 58430
0 5586 7 2 2 44403 54451
0 5587 7 2 2 52842 58609
0 5588 5 1 1 58781
0 5589 7 1 2 58779 58782
0 5590 7 1 2 5585 5589
0 5591 5 1 1 5590
0 5592 7 1 2 51880 57333
0 5593 5 1 1 5592
0 5594 7 1 2 45189 5593
0 5595 5 2 1 5594
0 5596 7 10 2 43231 47370
0 5597 5 2 1 58785
0 5598 7 3 2 58341 58786
0 5599 5 2 1 58797
0 5600 7 1 2 58783 58800
0 5601 5 1 1 5600
0 5602 7 1 2 55888 5601
0 5603 5 1 1 5602
0 5604 7 5 2 43004 52843
0 5605 5 2 1 58802
0 5606 7 3 2 57965 58074
0 5607 5 1 1 58809
0 5608 7 1 2 58803 58810
0 5609 5 1 1 5608
0 5610 7 1 2 5603 5609
0 5611 5 1 1 5610
0 5612 7 1 2 53985 58772
0 5613 7 1 2 5611 5612
0 5614 5 1 1 5613
0 5615 7 1 2 5591 5614
0 5616 5 1 1 5615
0 5617 7 1 2 53579 5616
0 5618 5 1 1 5617
0 5619 7 2 2 53667 58748
0 5620 5 1 1 58812
0 5621 7 3 2 44404 51724
0 5622 7 1 2 51395 58814
0 5623 7 1 2 58813 5622
0 5624 5 1 1 5623
0 5625 7 1 2 5618 5624
0 5626 7 1 2 5584 5625
0 5627 5 1 1 5626
0 5628 7 1 2 45514 5627
0 5629 5 1 1 5628
0 5630 7 1 2 46622 57666
0 5631 5 2 1 5630
0 5632 7 1 2 57727 58817
0 5633 5 1 1 5632
0 5634 7 1 2 58763 5633
0 5635 5 1 1 5634
0 5636 7 1 2 48545 50337
0 5637 5 2 1 5636
0 5638 7 4 2 44894 50979
0 5639 7 1 2 54514 58821
0 5640 7 2 2 58819 5639
0 5641 7 1 2 58778 58825
0 5642 5 1 1 5641
0 5643 7 1 2 5635 5642
0 5644 5 1 1 5643
0 5645 7 1 2 45678 5644
0 5646 5 1 1 5645
0 5647 7 1 2 58826 58770
0 5648 5 1 1 5647
0 5649 7 1 2 58760 58545
0 5650 5 1 1 5649
0 5651 7 1 2 5648 5650
0 5652 7 1 2 5646 5651
0 5653 5 1 1 5652
0 5654 7 1 2 58088 5653
0 5655 5 1 1 5654
0 5656 7 1 2 48398 5655
0 5657 7 1 2 5629 5656
0 5658 5 1 1 5657
0 5659 7 4 2 48768 53580
0 5660 7 2 2 55218 58827
0 5661 7 1 2 55396 56461
0 5662 7 2 2 58831 5661
0 5663 5 1 1 58833
0 5664 7 1 2 5620 5663
0 5665 5 1 1 5664
0 5666 7 1 2 44405 5665
0 5667 5 1 1 5666
0 5668 7 2 2 57626 57935
0 5669 7 1 2 46804 50377
0 5670 7 1 2 58835 5669
0 5671 7 1 2 56529 5670
0 5672 5 2 1 5671
0 5673 7 1 2 5667 58837
0 5674 5 1 1 5673
0 5675 7 1 2 44163 5674
0 5676 5 1 1 5675
0 5677 7 2 2 48769 53668
0 5678 7 1 2 56419 58693
0 5679 7 1 2 58839 5678
0 5680 5 1 1 5679
0 5681 7 1 2 5676 5680
0 5682 5 1 1 5681
0 5683 7 1 2 45515 5682
0 5684 5 1 1 5683
0 5685 7 1 2 44164 58749
0 5686 5 1 1 5685
0 5687 7 1 2 48770 58745
0 5688 5 1 1 5687
0 5689 7 1 2 5686 5688
0 5690 5 1 1 5689
0 5691 7 1 2 44406 58123
0 5692 7 1 2 5690 5691
0 5693 5 1 1 5692
0 5694 7 1 2 5684 5693
0 5695 5 1 1 5694
0 5696 7 1 2 43232 5695
0 5697 5 1 1 5696
0 5698 7 1 2 44002 58750
0 5699 5 1 1 5698
0 5700 7 1 2 51702 58743
0 5701 5 1 1 5700
0 5702 7 1 2 5699 5701
0 5703 5 1 1 5702
0 5704 7 1 2 58144 5703
0 5705 5 1 1 5704
0 5706 7 4 2 45516 44003
0 5707 7 1 2 44407 58834
0 5708 5 1 1 5707
0 5709 7 1 2 58838 5708
0 5710 5 1 1 5709
0 5711 7 1 2 58841 5710
0 5712 5 1 1 5711
0 5713 7 1 2 5705 5712
0 5714 5 1 1 5713
0 5715 7 1 2 48546 5714
0 5716 5 1 1 5715
0 5717 7 2 2 48771 58130
0 5718 7 2 2 44408 57766
0 5719 7 1 2 58694 58847
0 5720 7 1 2 58845 5719
0 5721 5 1 1 5720
0 5722 7 1 2 5716 5721
0 5723 7 1 2 5697 5722
0 5724 5 1 1 5723
0 5725 7 1 2 50628 5724
0 5726 5 1 1 5725
0 5727 7 2 2 49266 50053
0 5728 7 1 2 49815 58849
0 5729 5 1 1 5728
0 5730 7 1 2 52346 52706
0 5731 5 1 1 5730
0 5732 7 1 2 5729 5731
0 5733 5 1 1 5732
0 5734 7 1 2 45972 5733
0 5735 5 1 1 5734
0 5736 7 1 2 57278 58642
0 5737 7 1 2 52312 5736
0 5738 5 1 1 5737
0 5739 7 1 2 5735 5738
0 5740 5 1 1 5739
0 5741 7 1 2 58300 5740
0 5742 5 1 1 5741
0 5743 7 1 2 51777 55359
0 5744 7 1 2 58252 5743
0 5745 5 1 1 5744
0 5746 7 1 2 5742 5745
0 5747 5 1 1 5746
0 5748 7 1 2 44409 5747
0 5749 5 1 1 5748
0 5750 7 1 2 57988 58236
0 5751 5 1 1 5750
0 5752 7 4 2 44895 50741
0 5753 7 1 2 42473 58851
0 5754 5 1 1 5753
0 5755 7 1 2 5751 5754
0 5756 5 1 1 5755
0 5757 7 1 2 58048 5756
0 5758 5 1 1 5757
0 5759 7 2 2 51634 52525
0 5760 7 4 2 50742 51659
0 5761 5 1 1 58857
0 5762 7 1 2 58855 58858
0 5763 5 1 1 5762
0 5764 7 1 2 5758 5763
0 5765 5 1 1 5764
0 5766 7 6 2 47724 58172
0 5767 7 1 2 55360 58861
0 5768 7 1 2 5765 5767
0 5769 5 1 1 5768
0 5770 7 1 2 5749 5769
0 5771 5 1 1 5770
0 5772 7 1 2 50502 5771
0 5773 5 1 1 5772
0 5774 7 1 2 45044 5773
0 5775 7 1 2 5726 5774
0 5776 5 1 1 5775
0 5777 7 1 2 5658 5776
0 5778 5 1 1 5777
0 5779 7 8 2 47371 44410
0 5780 7 1 2 50915 58867
0 5781 7 1 2 54442 5780
0 5782 7 1 2 57483 5781
0 5783 7 1 2 56274 5782
0 5784 5 1 1 5783
0 5785 7 1 2 5778 5784
0 5786 5 1 1 5785
0 5787 7 1 2 55077 5786
0 5788 5 1 1 5787
0 5789 7 6 2 45973 56399
0 5790 5 1 1 58875
0 5791 7 1 2 53581 58876
0 5792 7 1 2 58365 5791
0 5793 5 1 1 5792
0 5794 7 4 2 43693 44165
0 5795 5 1 1 58881
0 5796 7 2 2 43233 58882
0 5797 7 6 2 45679 47952
0 5798 7 1 2 52146 56013
0 5799 7 1 2 58887 5798
0 5800 7 1 2 58885 5799
0 5801 5 1 1 5800
0 5802 7 1 2 5793 5801
0 5803 5 1 1 5802
0 5804 7 1 2 58089 5803
0 5805 5 1 1 5804
0 5806 7 12 2 42706 47508
0 5807 5 1 1 58893
0 5808 7 1 2 58053 58894
0 5809 5 3 1 5808
0 5810 7 1 2 55889 58366
0 5811 5 1 1 5810
0 5812 7 1 2 58905 5811
0 5813 5 1 1 5812
0 5814 7 4 2 46903 44621
0 5815 7 3 2 44732 58908
0 5816 7 1 2 50400 58912
0 5817 7 1 2 5813 5816
0 5818 5 1 1 5817
0 5819 7 10 2 44166 44411
0 5820 7 2 2 43234 58915
0 5821 7 1 2 55397 56054
0 5822 7 1 2 50688 5821
0 5823 7 1 2 58925 5822
0 5824 5 1 1 5823
0 5825 7 1 2 42135 5824
0 5826 7 1 2 5818 5825
0 5827 5 1 1 5826
0 5828 7 5 2 58058 58916
0 5829 5 2 1 58927
0 5830 7 1 2 58906 58932
0 5831 5 1 1 5830
0 5832 7 1 2 52543 5831
0 5833 5 1 1 5832
0 5834 7 2 2 49894 55749
0 5835 7 1 2 56400 58917
0 5836 7 1 2 58934 5835
0 5837 5 1 1 5836
0 5838 7 1 2 5833 5837
0 5839 5 1 1 5838
0 5840 7 1 2 45395 5839
0 5841 5 1 1 5840
0 5842 7 1 2 55562 56299
0 5843 5 1 1 5842
0 5844 7 1 2 58907 5843
0 5845 5 1 1 5844
0 5846 7 1 2 52548 5845
0 5847 5 1 1 5846
0 5848 7 1 2 45680 5847
0 5849 7 1 2 5841 5848
0 5850 5 1 1 5849
0 5851 7 1 2 45517 5850
0 5852 7 1 2 5827 5851
0 5853 5 1 1 5852
0 5854 7 1 2 5805 5853
0 5855 5 1 1 5854
0 5856 7 1 2 43855 5855
0 5857 5 1 1 5856
0 5858 7 20 2 47725 44622
0 5859 7 3 2 44733 58936
0 5860 7 1 2 58173 58524
0 5861 7 1 2 58956 5860
0 5862 7 1 2 53623 5861
0 5863 5 1 1 5862
0 5864 7 1 2 5857 5863
0 5865 5 1 1 5864
0 5866 7 1 2 46428 5865
0 5867 5 1 1 5866
0 5868 7 2 2 45396 58131
0 5869 7 2 2 55137 58431
0 5870 7 3 2 44412 50657
0 5871 7 1 2 53522 58963
0 5872 7 1 2 58961 5871
0 5873 7 1 2 58959 5872
0 5874 5 1 1 5873
0 5875 7 1 2 5867 5874
0 5876 5 1 1 5875
0 5877 7 1 2 44541 5876
0 5878 5 1 1 5877
0 5879 7 7 2 47217 45397
0 5880 5 2 1 58966
0 5881 7 1 2 56915 58967
0 5882 7 1 2 56942 5881
0 5883 5 1 1 5882
0 5884 7 1 2 3642 5883
0 5885 5 1 1 5884
0 5886 7 1 2 42474 5885
0 5887 5 1 1 5886
0 5888 7 2 2 45398 55078
0 5889 7 5 2 45974 47726
0 5890 7 2 2 58913 58977
0 5891 7 1 2 58975 58982
0 5892 5 1 1 5891
0 5893 7 1 2 5887 5892
0 5894 5 1 1 5893
0 5895 7 1 2 45681 5894
0 5896 5 1 1 5895
0 5897 7 1 2 44413 56037
0 5898 7 1 2 56688 5897
0 5899 5 1 1 5898
0 5900 7 1 2 5896 5899
0 5901 5 1 1 5900
0 5902 7 4 2 45518 47509
0 5903 7 1 2 55730 58075
0 5904 7 1 2 58984 5903
0 5905 7 1 2 5901 5904
0 5906 5 1 1 5905
0 5907 7 1 2 5878 5906
0 5908 5 1 1 5907
0 5909 7 1 2 49833 5908
0 5910 5 1 1 5909
0 5911 7 1 2 56131 56686
0 5912 5 1 1 5911
0 5913 7 1 2 46159 55170
0 5914 7 1 2 56063 57432
0 5915 7 1 2 5913 5914
0 5916 5 1 1 5915
0 5917 7 1 2 5912 5916
0 5918 5 1 1 5917
0 5919 7 1 2 42475 5918
0 5920 5 1 1 5919
0 5921 7 2 2 52546 55083
0 5922 5 1 1 58988
0 5923 7 1 2 48772 58989
0 5924 5 1 1 5923
0 5925 7 1 2 5920 5924
0 5926 5 1 1 5925
0 5927 7 1 2 42136 5926
0 5928 5 1 1 5927
0 5929 7 2 2 52526 54209
0 5930 7 1 2 56055 56682
0 5931 7 1 2 58990 5930
0 5932 5 1 1 5931
0 5933 7 1 2 5928 5932
0 5934 5 1 1 5933
0 5935 7 1 2 46805 5934
0 5936 5 1 1 5935
0 5937 7 10 2 45682 43432
0 5938 7 2 2 55088 58914
0 5939 7 2 2 48773 59002
0 5940 7 1 2 58992 59004
0 5941 5 1 1 5940
0 5942 7 1 2 5936 5941
0 5943 5 1 1 5942
0 5944 7 1 2 45519 5943
0 5945 5 1 1 5944
0 5946 7 17 2 41970 45683
0 5947 7 3 2 46806 59006
0 5948 7 1 2 59005 59023
0 5949 5 1 1 5948
0 5950 7 1 2 5945 5949
0 5951 5 1 1 5950
0 5952 7 1 2 50819 5951
0 5953 5 1 1 5952
0 5954 7 1 2 56249 56943
0 5955 5 1 1 5954
0 5956 7 1 2 48774 56689
0 5957 5 1 1 5956
0 5958 7 1 2 5955 5957
0 5959 5 1 1 5958
0 5960 7 1 2 42476 5959
0 5961 5 1 1 5960
0 5962 7 1 2 5922 5961
0 5963 5 1 1 5962
0 5964 7 1 2 42137 5963
0 5965 5 1 1 5964
0 5966 7 1 2 50714 52530
0 5967 7 1 2 57038 5966
0 5968 5 1 1 5967
0 5969 7 1 2 5965 5968
0 5970 5 1 1 5969
0 5971 7 1 2 58174 5970
0 5972 5 1 1 5971
0 5973 7 1 2 58211 59003
0 5974 5 1 1 5973
0 5975 7 1 2 5972 5974
0 5976 5 1 1 5975
0 5977 7 1 2 49953 5976
0 5978 5 1 1 5977
0 5979 7 1 2 5953 5978
0 5980 5 1 1 5979
0 5981 7 1 2 56389 5980
0 5982 5 1 1 5981
0 5983 7 2 2 49547 57811
0 5984 5 16 1 59026
0 5985 7 2 2 56154 59028
0 5986 7 2 2 58175 59044
0 5987 7 1 2 57039 59046
0 5988 5 1 1 5987
0 5989 7 3 2 51740 58132
0 5990 7 1 2 58007 59048
0 5991 5 1 1 5990
0 5992 7 1 2 5988 5991
0 5993 5 1 1 5992
0 5994 7 1 2 45975 5993
0 5995 5 1 1 5994
0 5996 7 2 2 42477 55079
0 5997 5 1 1 59051
0 5998 7 1 2 59052 59047
0 5999 5 1 1 5998
0 6000 7 1 2 47872 5999
0 6001 7 1 2 5995 6000
0 6002 5 1 1 6001
0 6003 7 3 2 54374 54157
0 6004 5 1 1 59053
0 6005 7 1 2 5997 6004
0 6006 5 8 1 6005
0 6007 7 1 2 50658 59056
0 6008 7 1 2 59049 6007
0 6009 5 1 1 6008
0 6010 7 1 2 47218 56275
0 6011 7 1 2 58877 6010
0 6012 7 3 2 43005 49148
0 6013 5 2 1 59064
0 6014 7 2 2 49459 59067
0 6015 5 1 1 59069
0 6016 7 1 2 46623 59070
0 6017 5 1 1 6016
0 6018 7 1 2 46429 58355
0 6019 5 1 1 6018
0 6020 7 1 2 43235 56988
0 6021 7 1 2 6019 6020
0 6022 5 1 1 6021
0 6023 7 1 2 6017 6022
0 6024 7 1 2 6011 6023
0 6025 5 1 1 6024
0 6026 7 1 2 44542 6025
0 6027 7 1 2 6009 6026
0 6028 5 1 1 6027
0 6029 7 1 2 48226 6028
0 6030 7 1 2 6002 6029
0 6031 5 1 1 6030
0 6032 7 1 2 5982 6031
0 6033 5 1 1 6032
0 6034 7 1 2 44414 6033
0 6035 5 1 1 6034
0 6036 7 1 2 55035 58773
0 6037 7 2 2 59029 6036
0 6038 7 1 2 57063 59071
0 6039 5 1 1 6038
0 6040 7 1 2 51964 56554
0 6041 5 1 1 6040
0 6042 7 1 2 52027 56557
0 6043 5 1 1 6042
0 6044 7 1 2 6041 6043
0 6045 5 1 1 6044
0 6046 7 2 2 43236 49069
0 6047 5 4 1 59073
0 6048 7 2 2 57167 59075
0 6049 5 11 1 59079
0 6050 7 2 2 43006 59081
0 6051 5 1 1 59092
0 6052 7 2 2 53372 6051
0 6053 5 16 1 59094
0 6054 7 1 2 46904 59096
0 6055 7 1 2 6045 6054
0 6056 5 1 1 6055
0 6057 7 1 2 6039 6056
0 6058 5 1 1 6057
0 6059 7 1 2 45684 6058
0 6060 5 1 1 6059
0 6061 7 1 2 46160 53558
0 6062 7 1 2 59072 6061
0 6063 5 1 1 6062
0 6064 7 1 2 6060 6063
0 6065 5 1 1 6064
0 6066 7 1 2 53912 6065
0 6067 5 1 1 6066
0 6068 7 1 2 53303 56405
0 6069 7 1 2 59097 6068
0 6070 5 1 1 6069
0 6071 7 2 2 54431 57852
0 6072 7 1 2 58049 59112
0 6073 7 1 2 59030 6072
0 6074 5 1 1 6073
0 6075 7 1 2 6070 6074
0 6076 5 1 1 6075
0 6077 7 1 2 56624 6076
0 6078 5 1 1 6077
0 6079 7 1 2 6067 6078
0 6080 5 1 1 6079
0 6081 7 1 2 58862 6080
0 6082 5 1 1 6081
0 6083 7 1 2 6035 6082
0 6084 5 1 1 6083
0 6085 7 1 2 50256 6084
0 6086 5 1 1 6085
0 6087 7 1 2 5910 6086
0 6088 7 1 2 5788 6087
0 6089 7 1 2 5451 6088
0 6090 7 1 2 4895 6089
0 6091 7 1 2 4723 6090
0 6092 5 1 1 6091
0 6093 7 1 2 47595 6092
0 6094 5 1 1 6093
0 6095 7 1 2 50595 51725
0 6096 5 1 1 6095
0 6097 7 1 2 51199 56762
0 6098 5 3 1 6097
0 6099 7 1 2 6096 59114
0 6100 5 2 1 6099
0 6101 7 1 2 55890 59117
0 6102 5 1 1 6101
0 6103 7 1 2 49251 55602
0 6104 5 1 1 6103
0 6105 7 1 2 6102 6104
0 6106 5 1 1 6105
0 6107 7 1 2 58670 6106
0 6108 5 1 1 6107
0 6109 7 2 2 46624 52358
0 6110 5 1 1 59119
0 6111 7 1 2 59076 6110
0 6112 5 1 1 6111
0 6113 7 10 2 43518 53682
0 6114 7 1 2 55772 59121
0 6115 7 1 2 6112 6114
0 6116 5 1 1 6115
0 6117 7 1 2 6108 6116
0 6118 5 1 1 6117
0 6119 7 1 2 44279 6118
0 6120 5 1 1 6119
0 6121 7 40 2 47596 44415
0 6122 7 5 2 44167 59131
0 6123 7 1 2 48958 57421
0 6124 7 4 2 45685 44004
0 6125 7 1 2 58274 59176
0 6126 7 1 2 6123 6125
0 6127 7 1 2 59171 6126
0 6128 5 1 1 6127
0 6129 7 1 2 6120 6128
0 6130 5 1 1 6129
0 6131 7 1 2 50659 51128
0 6132 7 1 2 6130 6131
0 6133 5 1 1 6132
0 6134 7 1 2 58016 59118
0 6135 5 1 1 6134
0 6136 7 2 2 44005 50054
0 6137 5 2 1 59180
0 6138 7 1 2 52825 59182
0 6139 5 2 1 6138
0 6140 7 1 2 51847 55843
0 6141 7 1 2 59184 6140
0 6142 5 1 1 6141
0 6143 7 1 2 6135 6142
0 6144 5 1 1 6143
0 6145 7 29 2 43433 44280
0 6146 7 1 2 58878 59186
0 6147 7 1 2 6144 6146
0 6148 5 1 1 6147
0 6149 7 1 2 6133 6148
0 6150 5 1 1 6149
0 6151 7 1 2 43007 6150
0 6152 5 1 1 6151
0 6153 7 2 2 42478 56455
0 6154 7 1 2 53554 59215
0 6155 5 1 1 6154
0 6156 7 6 2 44734 50401
0 6157 7 8 2 47727 54496
0 6158 7 1 2 59217 59223
0 6159 5 1 1 6158
0 6160 7 1 2 6155 6159
0 6161 5 1 1 6160
0 6162 7 2 2 53582 6161
0 6163 7 1 2 45399 59231
0 6164 5 1 1 6163
0 6165 7 2 2 50503 56420
0 6166 7 1 2 56080 59233
0 6167 5 1 1 6166
0 6168 7 1 2 6164 6167
0 6169 5 1 1 6168
0 6170 7 1 2 47510 6169
0 6171 5 1 1 6170
0 6172 7 1 2 52778 57458
0 6173 7 1 2 50898 6172
0 6174 5 1 1 6173
0 6175 7 1 2 6171 6174
0 6176 5 1 1 6175
0 6177 7 1 2 48547 6176
0 6178 5 1 1 6177
0 6179 7 1 2 49495 59232
0 6180 5 1 1 6179
0 6181 7 9 2 43237 43519
0 6182 7 3 2 42138 59235
0 6183 7 1 2 53177 59216
0 6184 7 1 2 59244 6183
0 6185 5 1 1 6184
0 6186 7 1 2 6180 6185
0 6187 5 1 1 6186
0 6188 7 1 2 49070 6187
0 6189 5 1 1 6188
0 6190 7 74 2 42139 44543
0 6191 5 3 1 59247
0 6192 7 3 2 55844 59248
0 6193 7 1 2 49198 58432
0 6194 7 1 2 52539 6193
0 6195 7 1 2 59324 6194
0 6196 5 1 1 6195
0 6197 7 1 2 6189 6196
0 6198 7 1 2 6178 6197
0 6199 5 1 1 6198
0 6200 7 8 2 44006 44281
0 6201 7 4 2 43434 59327
0 6202 7 1 2 6199 59335
0 6203 5 1 1 6202
0 6204 7 1 2 6152 6203
0 6205 5 1 1 6204
0 6206 7 1 2 41971 6205
0 6207 5 1 1 6206
0 6208 7 3 2 44007 52374
0 6209 5 2 1 59339
0 6210 7 1 2 50629 52882
0 6211 5 1 1 6210
0 6212 7 2 2 59342 6211
0 6213 5 3 1 59344
0 6214 7 1 2 50743 59346
0 6215 5 1 1 6214
0 6216 7 1 2 53843 6215
0 6217 5 1 1 6216
0 6218 7 2 2 50899 6217
0 6219 7 28 2 41972 44282
0 6220 7 37 2 47728 59351
0 6221 7 1 2 59349 59379
0 6222 5 1 1 6221
0 6223 7 3 2 45520 48959
0 6224 7 2 2 51328 59416
0 6225 7 8 2 47597 55773
0 6226 7 1 2 51129 51384
0 6227 7 1 2 54643 6226
0 6228 7 1 2 59421 6227
0 6229 7 1 2 59419 6228
0 6230 5 1 1 6229
0 6231 7 1 2 6222 6230
0 6232 5 1 1 6231
0 6233 7 1 2 53669 6232
0 6234 5 1 1 6233
0 6235 7 1 2 43520 59350
0 6236 5 1 1 6235
0 6237 7 1 2 43008 58859
0 6238 7 2 2 48991 50660
0 6239 7 3 2 44008 51130
0 6240 7 1 2 59429 59431
0 6241 7 1 2 6237 6240
0 6242 5 1 1 6241
0 6243 7 1 2 6236 6242
0 6244 5 1 1 6243
0 6245 7 1 2 42140 6244
0 6246 5 1 1 6245
0 6247 7 1 2 43009 55670
0 6248 7 1 2 52531 6247
0 6249 7 3 2 46625 55138
0 6250 7 1 2 59430 59434
0 6251 7 1 2 6248 6250
0 6252 5 1 1 6251
0 6253 7 1 2 6246 6252
0 6254 5 1 1 6253
0 6255 7 1 2 44283 56030
0 6256 7 1 2 6254 6255
0 6257 5 1 1 6256
0 6258 7 1 2 6234 6257
0 6259 7 1 2 6207 6258
0 6260 5 1 1 6259
0 6261 7 1 2 54591 1892
0 6262 5 1 1 6261
0 6263 7 1 2 6260 6262
0 6264 5 1 1 6263
0 6265 7 12 2 47598 58133
0 6266 7 2 2 49548 49737
0 6267 5 1 1 59449
0 6268 7 1 2 43010 6267
0 6269 5 1 1 6268
0 6270 7 1 2 54348 6269
0 6271 5 1 1 6270
0 6272 7 1 2 59437 6271
0 6273 5 1 1 6272
0 6274 7 5 2 43435 44168
0 6275 7 2 2 59236 59451
0 6276 7 4 2 56227 59456
0 6277 7 7 2 44284 48775
0 6278 7 1 2 59458 59462
0 6279 5 1 1 6278
0 6280 7 1 2 6273 6279
0 6281 5 1 1 6280
0 6282 7 2 2 42479 52477
0 6283 7 1 2 6281 59469
0 6284 5 1 1 6283
0 6285 7 17 2 46807 47599
0 6286 7 13 2 53304 59471
0 6287 7 2 2 47372 51741
0 6288 5 3 1 59501
0 6289 7 1 2 46430 59502
0 6290 5 1 1 6289
0 6291 7 3 2 45190 49329
0 6292 5 1 1 59506
0 6293 7 1 2 48548 56102
0 6294 5 2 1 6293
0 6295 7 1 2 6292 59509
0 6296 5 1 1 6295
0 6297 7 1 2 50055 6296
0 6298 5 1 1 6297
0 6299 7 1 2 52203 56746
0 6300 5 1 1 6299
0 6301 7 1 2 6298 6300
0 6302 7 1 2 6290 6301
0 6303 5 2 1 6302
0 6304 7 1 2 59488 59511
0 6305 5 1 1 6304
0 6306 7 14 2 43521 44285
0 6307 7 22 2 53683 59513
0 6308 5 5 1 59527
0 6309 7 1 2 52306 59528
0 6310 5 1 1 6309
0 6311 7 1 2 6305 6310
0 6312 5 1 1 6311
0 6313 7 1 2 42480 6312
0 6314 5 1 1 6313
0 6315 7 1 2 43011 57385
0 6316 7 5 2 42141 44009
0 6317 7 2 2 44286 59554
0 6318 7 1 2 59457 59559
0 6319 7 1 2 6315 6318
0 6320 5 1 1 6319
0 6321 7 1 2 6314 6320
0 6322 5 1 1 6321
0 6323 7 1 2 41973 6322
0 6324 5 1 1 6323
0 6325 7 19 2 45521 47600
0 6326 7 4 2 53670 59561
0 6327 5 1 1 59580
0 6328 7 1 2 42481 59581
0 6329 7 1 2 59512 6328
0 6330 5 1 1 6329
0 6331 7 1 2 45045 6330
0 6332 7 1 2 6324 6331
0 6333 5 1 1 6332
0 6334 7 3 2 47373 57860
0 6335 7 1 2 55147 59584
0 6336 5 2 1 6335
0 6337 7 5 2 45976 43012
0 6338 7 1 2 56674 59589
0 6339 5 1 1 6338
0 6340 7 1 2 59587 6339
0 6341 5 1 1 6340
0 6342 7 1 2 59438 6341
0 6343 5 1 1 6342
0 6344 7 3 2 41974 53684
0 6345 7 13 2 44169 44287
0 6346 7 8 2 48549 59597
0 6347 7 1 2 43522 49895
0 6348 7 1 2 59610 6347
0 6349 7 1 2 59594 6348
0 6350 5 1 1 6349
0 6351 7 1 2 48399 6350
0 6352 7 1 2 6343 6351
0 6353 5 1 1 6352
0 6354 7 1 2 48227 6353
0 6355 7 1 2 6333 6354
0 6356 5 1 1 6355
0 6357 7 1 2 6284 6356
0 6358 5 1 1 6357
0 6359 7 1 2 50661 6358
0 6360 5 1 1 6359
0 6361 7 4 2 48776 49738
0 6362 5 2 1 59618
0 6363 7 5 2 45400 50596
0 6364 7 3 2 47511 59624
0 6365 5 2 1 59629
0 6366 7 1 2 59622 59632
0 6367 5 1 1 6366
0 6368 7 1 2 46626 6367
0 6369 5 1 1 6368
0 6370 7 7 2 48777 50597
0 6371 5 4 1 59634
0 6372 7 4 2 43238 49739
0 6373 5 1 1 59645
0 6374 7 1 2 59641 59646
0 6375 5 2 1 6374
0 6376 7 1 2 6369 59649
0 6377 5 1 1 6376
0 6378 7 1 2 45046 6377
0 6379 5 1 1 6378
0 6380 7 1 2 55205 55254
0 6381 5 1 1 6380
0 6382 7 1 2 45191 57576
0 6383 7 1 2 6381 6382
0 6384 5 1 1 6383
0 6385 7 1 2 6379 6384
0 6386 5 2 1 6385
0 6387 7 2 2 47601 56276
0 6388 7 1 2 58695 59653
0 6389 7 1 2 59651 6388
0 6390 5 1 1 6389
0 6391 7 1 2 6360 6390
0 6392 5 1 1 6391
0 6393 7 1 2 43694 6392
0 6394 5 1 1 6393
0 6395 7 5 2 44896 50504
0 6396 7 1 2 56277 59655
0 6397 7 1 2 59652 6396
0 6398 5 1 1 6397
0 6399 7 8 2 45522 43013
0 6400 7 1 2 53638 59660
0 6401 5 1 1 6400
0 6402 7 1 2 56132 58212
0 6403 5 1 1 6402
0 6404 7 1 2 6401 6403
0 6405 5 1 1 6404
0 6406 7 1 2 56474 56675
0 6407 7 1 2 6405 6406
0 6408 5 1 1 6407
0 6409 7 1 2 6398 6408
0 6410 5 1 1 6409
0 6411 7 1 2 47602 6410
0 6412 5 1 1 6411
0 6413 7 1 2 44288 50662
0 6414 7 1 2 49868 6413
0 6415 7 1 2 59459 6414
0 6416 5 1 1 6415
0 6417 7 1 2 6412 6416
0 6418 5 1 1 6417
0 6419 7 1 2 47074 6418
0 6420 5 1 1 6419
0 6421 7 4 2 48076 49648
0 6422 7 14 2 44289 47953
0 6423 7 1 2 59668 59672
0 6424 7 4 2 42142 51329
0 6425 7 7 2 41975 55750
0 6426 7 2 2 49610 52830
0 6427 5 4 1 59697
0 6428 7 1 2 59690 59698
0 6429 7 1 2 59686 6428
0 6430 7 1 2 6423 6429
0 6431 5 1 1 6430
0 6432 7 1 2 6420 6431
0 6433 5 1 1 6432
0 6434 7 1 2 42482 6433
0 6435 5 1 1 6434
0 6436 7 1 2 52478 56847
0 6437 5 1 1 6436
0 6438 7 1 2 5327 6437
0 6439 5 1 1 6438
0 6440 7 1 2 43014 6439
0 6441 5 1 1 6440
0 6442 7 5 2 46431 48228
0 6443 7 1 2 49679 49954
0 6444 5 2 1 6443
0 6445 7 1 2 57858 59708
0 6446 5 1 1 6445
0 6447 7 1 2 50056 50247
0 6448 5 1 1 6447
0 6449 7 1 2 6446 6448
0 6450 5 1 1 6449
0 6451 7 1 2 59703 6450
0 6452 5 1 1 6451
0 6453 7 1 2 6441 6452
0 6454 5 1 1 6453
0 6455 7 1 2 58879 59654
0 6456 7 1 2 6454 6455
0 6457 5 1 1 6456
0 6458 7 1 2 44544 6457
0 6459 7 1 2 6435 6458
0 6460 7 1 2 6394 6459
0 6461 5 1 1 6460
0 6462 7 10 2 44897 53232
0 6463 5 1 1 59710
0 6464 7 1 2 53891 6463
0 6465 5 1 1 6464
0 6466 7 1 2 51713 58546
0 6467 5 3 1 6466
0 6468 7 1 2 57728 59720
0 6469 5 1 1 6468
0 6470 7 3 2 47603 55792
0 6471 7 1 2 59007 59723
0 6472 5 1 1 6471
0 6473 7 1 2 6327 6472
0 6474 5 2 1 6473
0 6475 7 1 2 6469 59726
0 6476 5 1 1 6475
0 6477 7 8 2 59122 59352
0 6478 7 1 2 52248 59728
0 6479 5 1 1 6478
0 6480 7 1 2 6476 6479
0 6481 5 1 1 6480
0 6482 7 1 2 45047 6481
0 6483 5 1 1 6482
0 6484 7 2 2 51219 58134
0 6485 7 4 2 47374 47604
0 6486 7 3 2 49377 59738
0 6487 7 1 2 46432 59742
0 6488 7 1 2 59736 6487
0 6489 5 1 1 6488
0 6490 7 1 2 6483 6489
0 6491 5 1 1 6490
0 6492 7 1 2 6465 6491
0 6493 5 1 1 6492
0 6494 7 8 2 47605 50402
0 6495 7 2 2 53762 59745
0 6496 7 1 2 58104 59753
0 6497 5 1 1 6496
0 6498 7 7 2 46905 58111
0 6499 7 1 2 59754 59755
0 6500 5 1 1 6499
0 6501 7 1 2 45401 59529
0 6502 7 1 2 50257 6501
0 6503 5 1 1 6502
0 6504 7 1 2 6500 6503
0 6505 5 1 1 6504
0 6506 7 1 2 41976 51165
0 6507 7 1 2 6505 6506
0 6508 5 1 1 6507
0 6509 7 1 2 6497 6508
0 6510 5 1 1 6509
0 6511 7 1 2 44170 6510
0 6512 5 1 1 6511
0 6513 7 2 2 53870 59439
0 6514 7 1 2 59635 59762
0 6515 5 1 1 6514
0 6516 7 1 2 6512 6515
0 6517 5 1 1 6516
0 6518 7 1 2 43239 6517
0 6519 5 1 1 6518
0 6520 7 5 2 50598 58452
0 6521 7 1 2 59763 59764
0 6522 5 1 1 6521
0 6523 7 1 2 6519 6522
0 6524 5 1 1 6523
0 6525 7 1 2 43015 6524
0 6526 5 1 1 6525
0 6527 7 3 2 58059 59353
0 6528 5 1 1 59769
0 6529 7 3 2 45977 49611
0 6530 7 1 2 52429 52779
0 6531 7 1 2 59772 6530
0 6532 7 1 2 59770 6531
0 6533 5 1 1 6532
0 6534 7 1 2 6526 6533
0 6535 5 1 1 6534
0 6536 7 1 2 44898 6535
0 6537 5 1 1 6536
0 6538 7 1 2 6493 6537
0 6539 5 1 1 6538
0 6540 7 1 2 50505 6539
0 6541 5 1 1 6540
0 6542 7 25 2 47606 58176
0 6543 7 1 2 54865 58807
0 6544 5 4 1 6543
0 6545 7 2 2 50744 59800
0 6546 5 1 1 59804
0 6547 7 1 2 59775 59805
0 6548 5 1 1 6547
0 6549 7 4 2 44290 45192
0 6550 7 3 2 48888 59806
0 6551 5 3 1 59810
0 6552 7 1 2 6548 59813
0 6553 5 1 1 6552
0 6554 7 1 2 45048 6553
0 6555 5 1 1 6554
0 6556 7 4 2 46433 47607
0 6557 7 4 2 58177 59816
0 6558 7 1 2 50248 59820
0 6559 5 1 1 6558
0 6560 7 44 2 44291 48889
0 6561 5 2 1 59824
0 6562 7 2 2 45049 59825
0 6563 5 1 1 59870
0 6564 7 1 2 6559 6563
0 6565 5 1 1 6564
0 6566 7 1 2 51220 6565
0 6567 5 1 1 6566
0 6568 7 1 2 6555 6567
0 6569 5 1 1 6568
0 6570 7 1 2 51131 6569
0 6571 5 1 1 6570
0 6572 7 2 2 58275 59661
0 6573 7 16 2 44010 47608
0 6574 7 1 2 49023 59874
0 6575 7 1 2 59872 6574
0 6576 5 1 1 6575
0 6577 7 5 2 45523 43240
0 6578 7 1 2 49071 50980
0 6579 5 2 1 6578
0 6580 7 4 2 49330 59895
0 6581 7 2 2 59472 59897
0 6582 7 1 2 59890 59901
0 6583 5 1 1 6582
0 6584 7 22 2 41977 59187
0 6585 5 2 1 59903
0 6586 7 1 2 49024 59904
0 6587 5 1 1 6586
0 6588 7 4 2 46808 59662
0 6589 7 1 2 59875 59927
0 6590 5 2 1 6589
0 6591 7 1 2 6528 59931
0 6592 5 1 1 6591
0 6593 7 1 2 49199 6592
0 6594 5 1 1 6593
0 6595 7 1 2 6587 6594
0 6596 7 1 2 6583 6595
0 6597 5 1 1 6596
0 6598 7 1 2 48550 6597
0 6599 5 1 1 6598
0 6600 7 1 2 6576 6599
0 6601 5 1 1 6600
0 6602 7 1 2 54199 6601
0 6603 5 1 1 6602
0 6604 7 1 2 6571 6603
0 6605 5 1 1 6604
0 6606 7 1 2 48229 6605
0 6607 5 1 1 6606
0 6608 7 1 2 57522 59776
0 6609 5 1 1 6608
0 6610 7 1 2 50820 59905
0 6611 5 3 1 6610
0 6612 7 1 2 6609 59933
0 6613 5 1 1 6612
0 6614 7 1 2 48551 6613
0 6615 5 1 1 6614
0 6616 7 5 2 46809 44011
0 6617 7 4 2 45524 59936
0 6618 7 8 2 43241 47609
0 6619 7 1 2 50287 59945
0 6620 7 1 2 59941 6619
0 6621 5 1 1 6620
0 6622 7 1 2 6615 6621
0 6623 5 1 1 6622
0 6624 7 1 2 48778 6623
0 6625 5 1 1 6624
0 6626 7 5 2 41978 58060
0 6627 7 1 2 59611 59953
0 6628 5 1 1 6627
0 6629 7 1 2 6625 6628
0 6630 5 1 1 6629
0 6631 7 1 2 50718 58224
0 6632 7 1 2 6630 6631
0 6633 5 1 1 6632
0 6634 7 1 2 6607 6633
0 6635 5 1 1 6634
0 6636 7 1 2 56155 6635
0 6637 5 1 1 6636
0 6638 7 1 2 47873 6637
0 6639 7 1 2 6541 6638
0 6640 5 1 1 6639
0 6641 7 1 2 6461 6640
0 6642 5 1 1 6641
0 6643 7 10 2 46434 43436
0 6644 7 6 2 45402 51166
0 6645 5 1 1 59968
0 6646 7 2 2 59958 59969
0 6647 7 2 2 50745 52780
0 6648 7 1 2 44292 59976
0 6649 7 1 2 59974 6648
0 6650 5 1 1 6649
0 6651 7 1 2 59746 59756
0 6652 7 1 2 51206 6651
0 6653 5 1 1 6652
0 6654 7 1 2 6650 6653
0 6655 5 1 1 6654
0 6656 7 1 2 41979 6655
0 6657 5 1 1 6656
0 6658 7 1 2 51742 59747
0 6659 7 1 2 58105 6658
0 6660 5 1 1 6659
0 6661 7 1 2 6657 6660
0 6662 5 1 1 6661
0 6663 7 1 2 50506 6662
0 6664 5 1 1 6663
0 6665 7 8 2 46810 43695
0 6666 7 6 2 45525 42483
0 6667 7 3 2 47610 59986
0 6668 7 1 2 59978 59992
0 6669 7 1 2 59045 6668
0 6670 5 1 1 6669
0 6671 7 1 2 6664 6670
0 6672 5 1 1 6671
0 6673 7 1 2 47874 6672
0 6674 5 1 1 6673
0 6675 7 13 2 47611 44545
0 6676 7 3 2 50507 59995
0 6677 7 2 2 56278 60008
0 6678 7 1 2 54068 60011
0 6679 5 1 1 6678
0 6680 7 1 2 6674 6679
0 6681 5 1 1 6680
0 6682 7 1 2 49834 6681
0 6683 5 1 1 6682
0 6684 7 4 2 53233 54757
0 6685 7 1 2 50321 55363
0 6686 5 1 1 6685
0 6687 7 1 2 54443 6686
0 6688 7 1 2 60013 6687
0 6689 5 1 1 6688
0 6690 7 11 2 46435 46811
0 6691 7 1 2 56464 60017
0 6692 7 3 2 45050 48992
0 6693 7 2 2 45526 51132
0 6694 7 1 2 60028 60031
0 6695 7 1 2 6691 6694
0 6696 5 1 1 6695
0 6697 7 1 2 6689 6696
0 6698 5 1 1 6697
0 6699 7 1 2 47612 53583
0 6700 7 1 2 6698 6699
0 6701 5 1 1 6700
0 6702 7 10 2 44546 48077
0 6703 7 3 2 55219 60033
0 6704 7 1 2 50449 60043
0 6705 5 1 1 6704
0 6706 7 1 2 56402 6705
0 6707 5 1 1 6706
0 6708 7 6 2 41980 43523
0 6709 7 2 2 48779 60046
0 6710 7 4 2 44293 53685
0 6711 7 1 2 43016 60054
0 6712 7 1 2 60052 6711
0 6713 7 1 2 50258 6712
0 6714 7 1 2 6707 6713
0 6715 5 1 1 6714
0 6716 7 1 2 6701 6715
0 6717 5 1 1 6716
0 6718 7 1 2 55563 6717
0 6719 5 1 1 6718
0 6720 7 1 2 51207 53234
0 6721 7 1 2 59440 6720
0 6722 5 1 1 6721
0 6723 7 3 2 50746 51098
0 6724 7 1 2 45403 60058
0 6725 7 1 2 59729 6724
0 6726 5 1 1 6725
0 6727 7 1 2 6722 6726
0 6728 5 1 1 6727
0 6729 7 1 2 56169 6728
0 6730 5 1 1 6729
0 6731 7 1 2 44416 6730
0 6732 7 1 2 6719 6731
0 6733 7 1 2 6683 6732
0 6734 7 1 2 6642 6733
0 6735 5 1 1 6734
0 6736 7 3 2 46812 59996
0 6737 7 2 2 59113 60061
0 6738 7 1 2 52375 58625
0 6739 7 1 2 50126 6738
0 6740 5 1 1 6739
0 6741 7 1 2 59588 6740
0 6742 5 1 1 6741
0 6743 7 1 2 48400 6742
0 6744 5 1 1 6743
0 6745 7 2 2 48993 58413
0 6746 5 2 1 60066
0 6747 7 2 2 49025 50539
0 6748 5 1 1 60070
0 6749 7 2 2 60068 6748
0 6750 7 1 2 43242 60072
0 6751 5 1 1 6750
0 6752 7 1 2 51498 58676
0 6753 5 1 1 6752
0 6754 7 1 2 46627 5588
0 6755 7 1 2 6753 6754
0 6756 5 1 1 6755
0 6757 7 1 2 45051 6756
0 6758 7 2 2 6751 6757
0 6759 5 1 1 60074
0 6760 7 1 2 42484 60075
0 6761 5 1 1 6760
0 6762 7 1 2 6744 6761
0 6763 5 1 1 6762
0 6764 7 1 2 60064 6763
0 6765 5 1 1 6764
0 6766 7 5 2 47375 44623
0 6767 7 2 2 60076 60062
0 6768 7 2 2 44735 49563
0 6769 7 1 2 60083 59590
0 6770 7 1 2 60081 6769
0 6771 5 1 1 6770
0 6772 7 7 2 42485 48401
0 6773 5 1 1 60085
0 6774 7 2 2 48552 60086
0 6775 7 1 2 56568 59336
0 6776 7 1 2 60092 6775
0 6777 5 1 1 6776
0 6778 7 1 2 6771 6777
0 6779 5 1 1 6778
0 6780 7 1 2 53913 6779
0 6781 5 1 1 6780
0 6782 7 2 2 49680 55016
0 6783 5 1 1 60094
0 6784 7 3 2 52501 59473
0 6785 7 1 2 54444 60096
0 6786 5 1 1 6785
0 6787 7 6 2 43696 44294
0 6788 7 4 2 43437 60099
0 6789 7 1 2 56465 60105
0 6790 5 1 1 6789
0 6791 7 1 2 6786 6790
0 6792 5 1 1 6791
0 6793 7 1 2 60095 6792
0 6794 5 1 1 6793
0 6795 7 7 2 44736 52446
0 6796 7 2 2 54497 60109
0 6797 7 4 2 47075 59739
0 6798 7 1 2 51396 55398
0 6799 7 1 2 60118 6798
0 6800 7 1 2 60116 6799
0 6801 5 1 1 6800
0 6802 7 1 2 6794 6801
0 6803 7 1 2 6781 6802
0 6804 5 1 1 6803
0 6805 7 1 2 50821 6804
0 6806 5 1 1 6805
0 6807 7 2 2 56569 59188
0 6808 7 1 2 54565 60122
0 6809 5 1 1 6808
0 6810 7 1 2 59591 60065
0 6811 5 1 1 6810
0 6812 7 1 2 6809 6811
0 6813 5 1 1 6812
0 6814 7 4 2 49955 53463
0 6815 5 1 1 60124
0 6816 7 1 2 6813 60125
0 6817 5 1 1 6816
0 6818 7 5 2 47512 44295
0 6819 7 7 2 46628 43697
0 6820 7 4 2 42486 60133
0 6821 7 2 2 60128 60140
0 6822 7 3 2 43438 48230
0 6823 7 1 2 52278 60146
0 6824 7 1 2 56570 6823
0 6825 7 1 2 60144 6824
0 6826 5 1 1 6825
0 6827 7 1 2 6817 6826
0 6828 5 1 1 6827
0 6829 7 1 2 50599 6828
0 6830 5 1 1 6829
0 6831 7 1 2 6806 6830
0 6832 7 1 2 6765 6831
0 6833 7 1 2 49482 60093
0 6834 7 1 2 60123 6833
0 6835 5 1 1 6834
0 6836 7 4 2 54694 58563
0 6837 5 1 1 60149
0 6838 7 1 2 51726 60150
0 6839 5 1 1 6838
0 6840 7 1 2 6759 6839
0 6841 5 1 1 6840
0 6842 7 8 2 45978 46813
0 6843 7 1 2 60153 60009
0 6844 7 1 2 6841 6843
0 6845 5 1 1 6844
0 6846 7 1 2 6835 6845
0 6847 5 1 1 6846
0 6848 7 1 2 53914 6847
0 6849 5 1 1 6848
0 6850 7 2 2 47376 50274
0 6851 5 3 1 60161
0 6852 7 1 2 52327 59450
0 6853 5 1 1 6852
0 6854 7 3 2 60163 6853
0 6855 5 2 1 60166
0 6856 7 1 2 45052 60169
0 6857 5 1 1 6856
0 6858 7 1 2 53440 53828
0 6859 5 1 1 6858
0 6860 7 1 2 6857 6859
0 6861 5 1 1 6860
0 6862 7 1 2 42487 6861
0 6863 5 1 1 6862
0 6864 7 2 2 48553 55017
0 6865 7 1 2 49483 60171
0 6866 5 1 1 6865
0 6867 7 1 2 6863 6866
0 6868 5 1 1 6867
0 6869 7 16 2 44296 47875
0 6870 7 3 2 57132 60173
0 6871 7 1 2 56115 60189
0 6872 7 1 2 6868 6871
0 6873 5 1 1 6872
0 6874 7 1 2 6849 6873
0 6875 7 1 2 6832 6874
0 6876 5 1 1 6875
0 6877 7 1 2 53584 6876
0 6878 5 1 1 6877
0 6879 7 1 2 42488 56406
0 6880 5 1 1 6879
0 6881 7 1 2 53915 56558
0 6882 5 1 1 6881
0 6883 7 1 2 6880 6882
0 6884 5 1 1 6883
0 6885 7 1 2 49535 50540
0 6886 5 3 1 6885
0 6887 7 1 2 49252 60192
0 6888 5 4 1 6887
0 6889 7 1 2 46436 60195
0 6890 5 1 1 6889
0 6891 7 1 2 54708 59082
0 6892 5 1 1 6891
0 6893 7 1 2 6890 6892
0 6894 5 1 1 6893
0 6895 7 1 2 59489 6894
0 6896 5 1 1 6895
0 6897 7 2 2 50600 50747
0 6898 5 3 1 60199
0 6899 7 4 2 47377 50822
0 6900 5 3 1 60204
0 6901 7 4 2 45193 50823
0 6902 5 5 1 60211
0 6903 7 3 2 60208 60215
0 6904 5 1 1 60220
0 6905 7 1 2 60201 60221
0 6906 5 2 1 6905
0 6907 7 1 2 60223 59530
0 6908 5 1 1 6907
0 6909 7 1 2 6896 6908
0 6910 5 1 1 6909
0 6911 7 1 2 45053 6910
0 6912 5 1 1 6911
0 6913 7 12 2 47613 45404
0 6914 7 2 2 55677 58112
0 6915 7 1 2 60225 60237
0 6916 5 1 1 6915
0 6917 7 1 2 59549 6916
0 6918 5 1 1 6917
0 6919 7 1 2 48402 57584
0 6920 7 1 2 6918 6919
0 6921 5 1 1 6920
0 6922 7 1 2 6912 6921
0 6923 5 1 1 6922
0 6924 7 1 2 6884 6923
0 6925 5 1 1 6924
0 6926 7 1 2 50824 59531
0 6927 5 2 1 6926
0 6928 7 1 2 59098 59490
0 6929 5 1 1 6928
0 6930 7 1 2 60239 6929
0 6931 5 1 1 6930
0 6932 7 1 2 52800 54566
0 6933 5 1 1 6932
0 6934 7 1 2 44899 50516
0 6935 5 1 1 6934
0 6936 7 1 2 6933 6935
0 6937 5 1 1 6936
0 6938 7 1 2 56504 6937
0 6939 7 1 2 6931 6938
0 6940 5 1 1 6939
0 6941 7 1 2 6925 6940
0 6942 7 1 2 6878 6941
0 6943 5 1 1 6942
0 6944 7 1 2 45527 6943
0 6945 5 1 1 6944
0 6946 7 1 2 54567 57881
0 6947 5 1 1 6946
0 6948 7 3 2 49149 60134
0 6949 5 1 1 60241
0 6950 7 4 2 47378 48231
0 6951 7 1 2 58643 60244
0 6952 7 1 2 60242 6951
0 6953 5 1 1 6952
0 6954 7 1 2 6947 6953
0 6955 5 1 1 6954
0 6956 7 1 2 48403 6955
0 6957 5 1 1 6956
0 6958 7 1 2 50601 57369
0 6959 5 3 1 6958
0 6960 7 1 2 60167 60248
0 6961 5 1 1 6960
0 6962 7 1 2 45054 52522
0 6963 7 1 2 6961 6962
0 6964 5 1 1 6963
0 6965 7 1 2 6957 6964
0 6966 5 1 1 6965
0 6967 7 1 2 57903 6966
0 6968 5 1 1 6967
0 6969 7 1 2 45055 51452
0 6970 5 1 1 6969
0 6971 7 4 2 45979 52519
0 6972 5 1 1 60251
0 6973 7 1 2 6970 6972
0 6974 5 1 1 6973
0 6975 7 1 2 51208 60172
0 6976 5 1 1 6975
0 6977 7 1 2 53928 6976
0 6978 5 1 1 6977
0 6979 7 1 2 54469 6978
0 6980 7 1 2 6974 6979
0 6981 5 1 1 6980
0 6982 7 1 2 6968 6981
0 6983 5 1 1 6982
0 6984 7 1 2 53585 6983
0 6985 5 1 1 6984
0 6986 7 1 2 50748 1118
0 6987 7 2 2 53768 6986
0 6988 5 1 1 60255
0 6989 7 1 2 42489 60256
0 6990 5 1 1 6989
0 6991 7 1 2 49740 56368
0 6992 5 1 1 6991
0 6993 7 1 2 6783 6992
0 6994 5 1 1 6993
0 6995 7 1 2 50825 6994
0 6996 5 1 1 6995
0 6997 7 1 2 6990 6996
0 6998 5 1 1 6997
0 6999 7 1 2 56407 6998
0 7000 5 1 1 6999
0 7001 7 1 2 50316 50826
0 7002 5 1 1 7001
0 7003 7 1 2 6988 7002
0 7004 5 1 1 7003
0 7005 7 1 2 56559 7004
0 7006 5 1 1 7005
0 7007 7 6 2 44547 48554
0 7008 7 1 2 48404 60257
0 7009 7 1 2 50889 7008
0 7010 7 1 2 56551 7009
0 7011 5 1 1 7010
0 7012 7 1 2 7006 7011
0 7013 5 1 1 7012
0 7014 7 1 2 53916 7013
0 7015 5 1 1 7014
0 7016 7 1 2 7000 7015
0 7017 5 1 1 7016
0 7018 7 1 2 53671 7017
0 7019 5 1 1 7018
0 7020 7 1 2 6985 7019
0 7021 5 1 1 7020
0 7022 7 1 2 59354 7021
0 7023 5 1 1 7022
0 7024 7 1 2 47729 7023
0 7025 7 1 2 6945 7024
0 7026 5 1 1 7025
0 7027 7 7 2 55165 55529
0 7028 5 29 1 60263
0 7029 7 1 2 7026 60270
0 7030 7 1 2 6735 7029
0 7031 5 1 1 7030
0 7032 7 1 2 6264 7031
0 7033 7 1 2 6094 7032
0 7034 7 1 2 3440 7033
0 7035 5 1 1 7034
0 7036 7 15 2 45782 46950
0 7037 5 2 1 60299
0 7038 7 10 2 42253 43568
0 7039 5 1 1 60316
0 7040 7 15 2 60314 7039
0 7041 7 1 2 7035 60326
0 7042 5 1 1 7041
0 7043 7 70 2 44624 48078
0 7044 5 1 1 60341
0 7045 7 1 2 46161 57309
0 7046 5 1 1 7045
0 7047 7 1 2 50301 7046
0 7048 5 1 1 7047
0 7049 7 1 2 55891 7048
0 7050 5 1 1 7049
0 7051 7 8 2 47730 48780
0 7052 7 8 2 46814 44171
0 7053 5 1 1 60419
0 7054 7 2 2 60411 60420
0 7055 5 1 1 60427
0 7056 7 1 2 57243 60428
0 7057 5 1 1 7056
0 7058 7 1 2 7050 7057
0 7059 5 1 1 7058
0 7060 7 1 2 44012 7059
0 7061 5 1 1 7060
0 7062 7 4 2 46815 47076
0 7063 7 4 2 42707 47731
0 7064 7 1 2 60429 60433
0 7065 7 1 2 52328 7064
0 7066 5 1 1 7065
0 7067 7 1 2 7061 7066
0 7068 5 1 1 7067
0 7069 7 1 2 41981 7068
0 7070 5 1 1 7069
0 7071 7 1 2 42708 52329
0 7072 5 3 1 7071
0 7073 7 1 2 54349 60437
0 7074 5 2 1 7073
0 7075 7 41 2 45528 47732
0 7076 7 1 2 54412 60442
0 7077 7 1 2 60440 7076
0 7078 5 1 1 7077
0 7079 7 1 2 7070 7078
0 7080 5 1 1 7079
0 7081 7 1 2 44297 7080
0 7082 5 1 1 7081
0 7083 7 2 2 47379 51522
0 7084 5 1 1 60483
0 7085 7 4 2 42709 44417
0 7086 7 4 2 59562 60485
0 7087 7 1 2 60430 60489
0 7088 7 1 2 7084 7087
0 7089 5 1 1 7088
0 7090 7 1 2 7082 7089
0 7091 5 1 1 7090
0 7092 7 1 2 51848 7091
0 7093 5 1 1 7092
0 7094 7 7 2 42710 47614
0 7095 7 5 2 41982 57499
0 7096 5 2 1 60500
0 7097 7 1 2 45529 57649
0 7098 5 1 1 7097
0 7099 7 1 2 60505 7098
0 7100 5 1 1 7099
0 7101 7 1 2 44013 7100
0 7102 5 1 1 7101
0 7103 7 6 2 47733 59891
0 7104 7 1 2 60421 60507
0 7105 5 1 1 7104
0 7106 7 1 2 7102 7105
0 7107 5 1 1 7106
0 7108 7 1 2 60493 7107
0 7109 5 1 1 7108
0 7110 7 2 2 55453 59132
0 7111 5 1 1 60513
0 7112 7 1 2 47734 59337
0 7113 5 1 1 7112
0 7114 7 1 2 7111 7113
0 7115 5 1 1 7114
0 7116 7 1 2 41983 7115
0 7117 5 1 1 7116
0 7118 7 8 2 42711 43439
0 7119 7 31 2 44418 59563
0 7120 7 1 2 60515 60523
0 7121 5 1 1 7120
0 7122 7 1 2 7117 7121
0 7123 5 1 1 7122
0 7124 7 1 2 51743 7123
0 7125 5 1 1 7124
0 7126 7 1 2 7109 7125
0 7127 5 1 1 7126
0 7128 7 2 2 45686 47077
0 7129 7 1 2 44548 60554
0 7130 7 1 2 7127 7129
0 7131 5 1 1 7130
0 7132 7 1 2 7093 7131
0 7133 5 1 1 7132
0 7134 7 1 2 43017 7133
0 7135 5 1 1 7134
0 7136 7 20 2 45687 44549
0 7137 5 1 1 60556
0 7138 7 5 2 43440 47735
0 7139 7 2 2 60557 60576
0 7140 7 1 2 48781 60581
0 7141 5 1 1 7140
0 7142 7 3 2 46816 60412
0 7143 5 1 1 60583
0 7144 7 1 2 55926 7143
0 7145 5 3 1 7144
0 7146 7 1 2 42143 56991
0 7147 7 2 2 60586 7146
0 7148 5 1 1 60589
0 7149 7 1 2 7141 7148
0 7150 5 1 1 7149
0 7151 7 1 2 44298 7150
0 7152 5 1 1 7151
0 7153 7 4 2 45688 59133
0 7154 7 1 2 57779 59937
0 7155 7 1 2 60591 7154
0 7156 5 1 1 7155
0 7157 7 1 2 41984 7156
0 7158 7 1 2 7152 7157
0 7159 5 1 1 7158
0 7160 7 1 2 59134 59938
0 7161 5 2 1 7160
0 7162 7 4 2 43243 44299
0 7163 7 2 2 60597 60577
0 7164 5 2 1 60601
0 7165 7 1 2 60595 60603
0 7166 5 1 1 7165
0 7167 7 1 2 51849 7166
0 7168 5 1 1 7167
0 7169 7 4 2 43441 44014
0 7170 7 9 2 59135 60558
0 7171 5 1 1 60609
0 7172 7 1 2 60605 60610
0 7173 5 1 1 7172
0 7174 7 1 2 7168 7173
0 7175 5 1 1 7174
0 7176 7 1 2 48782 7175
0 7177 5 1 1 7176
0 7178 7 1 2 58276 59876
0 7179 7 1 2 58687 7178
0 7180 5 1 1 7179
0 7181 7 1 2 45530 7180
0 7182 7 1 2 7177 7181
0 7183 5 1 1 7182
0 7184 7 1 2 44172 7183
0 7185 7 1 2 7159 7184
0 7186 5 1 1 7185
0 7187 7 38 2 44300 47736
0 7188 7 7 2 43442 60618
0 7189 5 3 1 60656
0 7190 7 1 2 60663 60596
0 7191 5 1 1 7190
0 7192 7 1 2 41985 7191
0 7193 5 1 1 7192
0 7194 7 1 2 60524 60606
0 7195 5 1 1 7194
0 7196 7 1 2 7193 7195
0 7197 5 1 1 7196
0 7198 7 1 2 60559 7197
0 7199 5 1 1 7198
0 7200 7 16 2 42144 46817
0 7201 7 4 2 45531 60666
0 7202 7 4 2 47615 56421
0 7203 7 2 2 60682 60686
0 7204 7 1 2 44015 60690
0 7205 5 1 1 7204
0 7206 7 1 2 7199 7205
0 7207 5 1 1 7206
0 7208 7 1 2 51514 7207
0 7209 5 1 1 7208
0 7210 7 3 2 54758 60619
0 7211 7 2 2 52330 60692
0 7212 5 2 1 60695
0 7213 7 1 2 42145 55671
0 7214 7 1 2 60696 7213
0 7215 5 1 1 7214
0 7216 7 1 2 7209 7215
0 7217 7 1 2 7186 7216
0 7218 5 1 1 7217
0 7219 7 1 2 54841 7218
0 7220 5 1 1 7219
0 7221 7 1 2 7135 7220
0 7222 5 1 1 7221
0 7223 7 1 2 42490 7222
0 7224 5 1 1 7223
0 7225 7 8 2 43018 49026
0 7226 5 3 1 60699
0 7227 7 1 2 46162 60707
0 7228 5 7 1 7227
0 7229 7 6 2 47513 53737
0 7230 5 2 1 60717
0 7231 7 1 2 42712 60723
0 7232 5 4 1 7231
0 7233 7 2 2 60710 60725
0 7234 7 1 2 46629 60729
0 7235 5 1 1 7234
0 7236 7 1 2 45980 44173
0 7237 5 2 1 7236
0 7238 7 2 2 46163 58356
0 7239 5 1 1 60733
0 7240 7 1 2 60731 7239
0 7241 5 1 1 7240
0 7242 7 1 2 51330 7241
0 7243 5 1 1 7242
0 7244 7 1 2 7235 7243
0 7245 5 1 1 7244
0 7246 7 1 2 55892 7245
0 7247 5 1 1 7246
0 7248 7 1 2 1404 60438
0 7249 5 1 1 7248
0 7250 7 1 2 45981 55603
0 7251 7 1 2 7249 7250
0 7252 5 1 1 7251
0 7253 7 1 2 7247 7252
0 7254 5 1 1 7253
0 7255 7 1 2 44016 7254
0 7256 5 1 1 7255
0 7257 7 10 2 46630 45405
0 7258 5 10 1 60735
0 7259 7 3 2 43019 60745
0 7260 5 7 1 60755
0 7261 7 1 2 46437 53345
0 7262 5 4 1 7261
0 7263 7 2 2 44174 60765
0 7264 5 1 1 60769
0 7265 7 1 2 60758 7264
0 7266 5 1 1 7265
0 7267 7 1 2 55604 7266
0 7268 5 1 1 7267
0 7269 7 1 2 58933 7268
0 7270 5 1 1 7269
0 7271 7 1 2 54375 7270
0 7272 5 1 1 7271
0 7273 7 1 2 7256 7272
0 7274 5 1 1 7273
0 7275 7 1 2 51850 7274
0 7276 5 1 1 7275
0 7277 7 2 2 51744 53418
0 7278 7 6 2 45689 54461
0 7279 5 2 1 60773
0 7280 7 1 2 58978 60774
0 7281 7 1 2 60771 7280
0 7282 5 1 1 7281
0 7283 7 1 2 7276 7282
0 7284 5 1 1 7283
0 7285 7 1 2 44301 7284
0 7286 5 1 1 7285
0 7287 7 3 2 49331 51745
0 7288 5 1 1 60781
0 7289 7 1 2 50981 7288
0 7290 5 5 1 7289
0 7291 7 9 2 45690 45982
0 7292 7 3 2 55454 60789
0 7293 7 6 2 44550 59136
0 7294 7 1 2 60798 60801
0 7295 7 1 2 60784 7294
0 7296 5 1 1 7295
0 7297 7 1 2 41986 7296
0 7298 7 1 2 7286 7297
0 7299 5 1 1 7298
0 7300 7 6 2 43244 49875
0 7301 5 2 1 60807
0 7302 7 1 2 4113 60813
0 7303 5 9 1 7302
0 7304 7 1 2 54376 60815
0 7305 5 1 1 7304
0 7306 7 1 2 42491 57010
0 7307 7 1 2 58443 7306
0 7308 5 1 1 7307
0 7309 7 1 2 7305 7308
0 7310 5 1 1 7309
0 7311 7 1 2 55605 7310
0 7312 5 1 1 7311
0 7313 7 1 2 54377 55893
0 7314 7 1 2 60785 7313
0 7315 5 1 1 7314
0 7316 7 1 2 7312 7315
0 7317 5 1 1 7316
0 7318 7 1 2 60560 7317
0 7319 5 1 1 7318
0 7320 7 2 2 46818 56073
0 7321 7 1 2 56471 60824
0 7322 7 1 2 60786 7321
0 7323 5 1 1 7322
0 7324 7 1 2 7319 7323
0 7325 5 1 1 7324
0 7326 7 1 2 47616 7325
0 7327 5 1 1 7326
0 7328 7 1 2 43020 60441
0 7329 5 1 1 7328
0 7330 7 2 2 44017 52331
0 7331 5 3 1 60826
0 7332 7 2 2 52307 60828
0 7333 5 3 1 60831
0 7334 7 1 2 42713 60833
0 7335 5 1 1 7334
0 7336 7 1 2 7329 7335
0 7337 5 1 1 7336
0 7338 7 2 2 56074 60174
0 7339 7 1 2 60578 60836
0 7340 7 1 2 7337 7339
0 7341 5 1 1 7340
0 7342 7 1 2 45532 7341
0 7343 7 1 2 7327 7342
0 7344 5 1 1 7343
0 7345 7 1 2 43698 7344
0 7346 7 1 2 7299 7345
0 7347 5 1 1 7346
0 7348 7 1 2 7224 7347
0 7349 5 1 1 7348
0 7350 7 1 2 48555 7349
0 7351 5 1 1 7350
0 7352 7 3 2 44018 54842
0 7353 7 4 2 44419 51746
0 7354 7 3 2 51851 60841
0 7355 5 1 1 60845
0 7356 7 1 2 60838 60846
0 7357 5 1 1 7356
0 7358 7 3 2 50541 55095
0 7359 5 3 1 60848
0 7360 7 1 2 49027 60839
0 7361 5 1 1 7360
0 7362 7 1 2 60851 7361
0 7363 5 1 1 7362
0 7364 7 1 2 43245 7363
0 7365 5 1 1 7364
0 7366 7 4 2 45194 55096
0 7367 7 1 2 49883 55547
0 7368 7 1 2 55281 7367
0 7369 7 1 2 60854 7368
0 7370 5 1 1 7369
0 7371 7 1 2 7365 7370
0 7372 5 1 1 7371
0 7373 7 1 2 58710 7372
0 7374 5 1 1 7373
0 7375 7 1 2 7357 7374
0 7376 5 1 1 7375
0 7377 7 1 2 42492 7376
0 7378 5 1 1 7377
0 7379 7 4 2 47737 57780
0 7380 7 2 2 45691 49956
0 7381 7 1 2 60858 60862
0 7382 5 1 1 7381
0 7383 7 1 2 7355 7382
0 7384 5 1 1 7383
0 7385 7 1 2 54530 58626
0 7386 7 1 2 7384 7385
0 7387 5 1 1 7386
0 7388 7 1 2 7378 7387
0 7389 5 1 1 7388
0 7390 7 1 2 46819 7389
0 7391 5 1 1 7390
0 7392 7 2 2 53235 55774
0 7393 7 3 2 42714 58061
0 7394 7 1 2 45692 49876
0 7395 7 1 2 60866 7394
0 7396 7 1 2 60864 7395
0 7397 5 1 1 7396
0 7398 7 1 2 7391 7397
0 7399 5 1 1 7398
0 7400 7 1 2 43021 7399
0 7401 5 1 1 7400
0 7402 7 1 2 49778 60847
0 7403 5 1 1 7402
0 7404 7 1 2 46631 58357
0 7405 5 2 1 7404
0 7406 7 1 2 50177 60869
0 7407 5 1 1 7406
0 7408 7 1 2 44019 7407
0 7409 5 1 1 7408
0 7410 7 2 2 49028 58787
0 7411 5 3 1 60871
0 7412 7 1 2 7409 60873
0 7413 5 1 1 7412
0 7414 7 1 2 45195 58711
0 7415 7 1 2 7413 7414
0 7416 5 1 1 7415
0 7417 7 1 2 7403 7416
0 7418 5 1 1 7417
0 7419 7 3 2 53849 59979
0 7420 7 1 2 7418 60876
0 7421 5 1 1 7420
0 7422 7 1 2 7401 7421
0 7423 5 1 1 7422
0 7424 7 1 2 47617 7423
0 7425 5 1 1 7424
0 7426 7 2 2 53236 60579
0 7427 7 2 2 56198 59598
0 7428 7 3 2 43246 49332
0 7429 7 1 2 55418 60883
0 7430 7 1 2 60881 7429
0 7431 7 1 2 60879 7430
0 7432 5 1 1 7431
0 7433 7 1 2 7425 7432
0 7434 5 1 1 7433
0 7435 7 1 2 45533 7434
0 7436 5 1 1 7435
0 7437 7 8 2 47876 60667
0 7438 7 7 2 42715 44175
0 7439 7 2 2 55472 60894
0 7440 5 1 1 60901
0 7441 7 2 2 60886 60902
0 7442 7 1 2 57244 60903
0 7443 5 1 1 7442
0 7444 7 6 2 45196 54027
0 7445 5 1 1 60905
0 7446 7 1 2 50669 58993
0 7447 7 1 2 60906 7446
0 7448 5 1 1 7447
0 7449 7 1 2 7443 7448
0 7450 5 1 1 7449
0 7451 7 1 2 42493 7450
0 7452 5 1 1 7451
0 7453 7 1 2 45983 51363
0 7454 7 1 2 60904 7453
0 7455 5 1 1 7454
0 7456 7 1 2 7452 7455
0 7457 5 1 1 7456
0 7458 7 1 2 60620 7457
0 7459 5 1 1 7458
0 7460 7 8 2 45693 42716
0 7461 7 2 2 51331 60911
0 7462 7 10 2 44176 47618
0 7463 7 1 2 59939 60921
0 7464 7 1 2 60919 7463
0 7465 7 1 2 60865 7464
0 7466 5 1 1 7465
0 7467 7 1 2 7459 7466
0 7468 5 1 1 7467
0 7469 7 1 2 41987 7468
0 7470 5 1 1 7469
0 7471 7 1 2 7436 7470
0 7472 7 1 2 7351 7471
0 7473 5 1 1 7472
0 7474 7 1 2 60342 7473
0 7475 5 1 1 7474
0 7476 7 1 2 42717 49788
0 7477 5 1 1 7476
0 7478 7 6 2 48890 60621
0 7479 7 3 2 60561 60931
0 7480 5 3 1 60937
0 7481 7 1 2 7477 60938
0 7482 5 1 1 7481
0 7483 7 2 2 42718 50542
0 7484 5 5 1 60943
0 7485 7 2 2 57538 60945
0 7486 5 5 1 60950
0 7487 7 6 2 45694 46438
0 7488 7 1 2 57627 60957
0 7489 7 1 2 60952 7488
0 7490 5 1 1 7489
0 7491 7 6 2 42146 46164
0 7492 7 1 2 56422 60963
0 7493 7 1 2 52891 7492
0 7494 5 1 1 7493
0 7495 7 1 2 7490 7494
0 7496 5 1 1 7495
0 7497 7 1 2 59777 7496
0 7498 5 1 1 7497
0 7499 7 1 2 7482 7498
0 7500 5 1 1 7499
0 7501 7 25 2 51133 60343
0 7502 5 6 1 60969
0 7503 7 1 2 7500 60970
0 7504 5 1 1 7503
0 7505 7 4 2 44020 59137
0 7506 7 1 2 56865 61000
0 7507 7 7 2 47954 45197
0 7508 7 2 2 58288 61004
0 7509 7 18 2 45534 42147
0 7510 7 3 2 50403 61013
0 7511 7 1 2 61011 61031
0 7512 7 1 2 7506 7511
0 7513 5 1 1 7512
0 7514 7 1 2 7504 7513
0 7515 5 1 1 7514
0 7516 7 1 2 51221 7515
0 7517 5 1 1 7516
0 7518 7 5 2 42148 44420
0 7519 7 20 2 47877 61034
0 7520 5 1 1 61039
0 7521 7 5 2 45406 55564
0 7522 5 3 1 61059
0 7523 7 1 2 60209 61064
0 7524 5 1 1 7523
0 7525 7 1 2 46439 7524
0 7526 5 1 1 7525
0 7527 7 1 2 43247 49150
0 7528 5 5 1 7527
0 7529 7 3 2 60870 61067
0 7530 5 2 1 61072
0 7531 7 1 2 47380 61075
0 7532 5 1 1 7531
0 7533 7 1 2 7526 7532
0 7534 5 1 1 7533
0 7535 7 10 2 45535 46165
0 7536 7 4 2 48556 59474
0 7537 7 1 2 61077 61087
0 7538 7 1 2 7534 7537
0 7539 5 1 1 7538
0 7540 7 9 2 46166 47619
0 7541 7 4 2 58178 61091
0 7542 7 1 2 57835 61100
0 7543 5 1 1 7542
0 7544 7 1 2 56103 59826
0 7545 5 1 1 7544
0 7546 7 1 2 7543 7545
0 7547 5 1 1 7546
0 7548 7 1 2 56649 7547
0 7549 5 1 1 7548
0 7550 7 4 2 46632 48891
0 7551 7 1 2 48960 60129
0 7552 7 1 2 61104 7551
0 7553 5 1 1 7552
0 7554 7 1 2 7549 7553
0 7555 7 1 2 7539 7554
0 7556 5 1 1 7555
0 7557 7 1 2 61040 7556
0 7558 5 1 1 7557
0 7559 7 6 2 45407 49681
0 7560 5 1 1 61108
0 7561 7 1 2 59821 61109
0 7562 5 1 1 7561
0 7563 7 1 2 50602 59906
0 7564 5 1 1 7563
0 7565 7 1 2 7562 7564
0 7566 5 1 1 7565
0 7567 7 1 2 47514 7566
0 7568 5 1 1 7567
0 7569 7 1 2 58342 59907
0 7570 5 1 1 7569
0 7571 7 1 2 7568 7570
0 7572 5 1 1 7571
0 7573 7 1 2 46633 7572
0 7574 5 1 1 7573
0 7575 7 2 2 50827 57556
0 7576 5 1 1 61114
0 7577 7 1 2 61068 7576
0 7578 5 1 1 7577
0 7579 7 1 2 59827 7578
0 7580 5 1 1 7579
0 7581 7 1 2 7574 7580
0 7582 5 1 1 7581
0 7583 7 1 2 46167 7582
0 7584 5 1 1 7583
0 7585 7 1 2 49779 61060
0 7586 5 1 1 7585
0 7587 7 1 2 52191 55000
0 7588 5 1 1 7587
0 7589 7 1 2 7586 7588
0 7590 5 1 1 7589
0 7591 7 1 2 59828 7590
0 7592 5 1 1 7591
0 7593 7 1 2 7584 7592
0 7594 5 1 1 7593
0 7595 7 1 2 58712 7594
0 7596 5 1 1 7595
0 7597 7 1 2 7558 7596
0 7598 5 1 1 7597
0 7599 7 59 2 47955 44737
0 7600 5 2 1 61116
0 7601 7 23 2 50404 61117
0 7602 5 1 1 61177
0 7603 7 1 2 7598 61178
0 7604 5 1 1 7603
0 7605 7 1 2 7517 7604
0 7606 7 1 2 7475 7605
0 7607 5 1 1 7606
0 7608 7 1 2 43856 7607
0 7609 5 1 1 7608
0 7610 7 1 2 53346 61041
0 7611 5 1 1 7610
0 7612 7 2 2 44551 50338
0 7613 7 7 2 45695 46634
0 7614 7 1 2 47738 61202
0 7615 7 1 2 61200 7614
0 7616 5 1 1 7615
0 7617 7 1 2 7611 7616
0 7618 5 1 1 7617
0 7619 7 1 2 43022 7618
0 7620 5 1 1 7619
0 7621 7 2 2 45696 49120
0 7622 7 1 2 60859 61209
0 7623 5 1 1 7622
0 7624 7 1 2 7620 7623
0 7625 5 1 1 7624
0 7626 7 2 2 55455 59987
0 7627 7 3 2 43699 44625
0 7628 7 4 2 48079 61213
0 7629 7 1 2 47620 61216
0 7630 7 2 2 61211 7629
0 7631 7 1 2 7625 61220
0 7632 5 1 1 7631
0 7633 7 3 2 51852 60622
0 7634 5 1 1 61222
0 7635 7 1 2 7171 7634
0 7636 5 1 1 7635
0 7637 7 3 2 54759 7636
0 7638 7 1 2 60759 61225
0 7639 5 1 1 7638
0 7640 7 8 2 45536 46440
0 7641 7 2 2 59138 61228
0 7642 7 1 2 60887 61236
0 7643 5 1 1 7642
0 7644 7 1 2 60940 7643
0 7645 5 1 1 7644
0 7646 7 1 2 53347 7645
0 7647 5 1 1 7646
0 7648 7 3 2 48920 51853
0 7649 7 1 2 44302 61238
0 7650 5 2 1 7649
0 7651 7 5 2 45408 49913
0 7652 5 1 1 61243
0 7653 7 2 2 58688 59778
0 7654 7 1 2 61244 61248
0 7655 5 1 1 7654
0 7656 7 1 2 61241 7655
0 7657 7 1 2 7647 7656
0 7658 7 1 2 7639 7657
0 7659 5 1 1 7658
0 7660 7 1 2 50450 7659
0 7661 5 1 1 7660
0 7662 7 6 2 47078 47878
0 7663 7 1 2 56183 61250
0 7664 7 1 2 59687 7663
0 7665 7 1 2 59908 7664
0 7666 5 1 1 7665
0 7667 7 1 2 46168 7666
0 7668 7 1 2 7661 7667
0 7669 5 1 1 7668
0 7670 7 4 2 43023 58277
0 7671 7 18 2 45537 45697
0 7672 7 4 2 47621 61260
0 7673 7 1 2 54657 58979
0 7674 7 1 2 61278 7673
0 7675 7 1 2 61256 7674
0 7676 5 1 1 7675
0 7677 7 2 2 49914 56228
0 7678 7 3 2 43443 56948
0 7679 7 7 2 44303 44421
0 7680 7 1 2 61284 61287
0 7681 7 1 2 61282 7680
0 7682 5 1 1 7681
0 7683 7 1 2 42719 7682
0 7684 7 1 2 7676 7683
0 7685 5 1 1 7684
0 7686 7 1 2 47381 51167
0 7687 7 1 2 7685 7686
0 7688 7 1 2 7669 7687
0 7689 5 1 1 7688
0 7690 7 1 2 60736 61226
0 7691 5 1 1 7690
0 7692 7 1 2 61242 7691
0 7693 5 1 1 7692
0 7694 7 2 2 53237 54950
0 7695 7 1 2 7693 61294
0 7696 5 1 1 7695
0 7697 7 1 2 60939 61295
0 7698 5 1 1 7697
0 7699 7 1 2 47079 47622
0 7700 7 1 2 54378 7699
0 7701 7 1 2 59942 7700
0 7702 7 1 2 61042 7701
0 7703 5 1 1 7702
0 7704 7 1 2 7698 7703
0 7705 5 1 1 7704
0 7706 7 1 2 53348 7705
0 7707 5 1 1 7706
0 7708 7 1 2 7696 7707
0 7709 7 1 2 7689 7708
0 7710 5 1 1 7709
0 7711 7 1 2 61118 7710
0 7712 5 1 1 7711
0 7713 7 1 2 7632 7712
0 7714 5 1 1 7713
0 7715 7 1 2 47515 7714
0 7716 5 1 1 7715
0 7717 7 2 2 47080 59877
0 7718 7 3 2 54379 58179
0 7719 7 6 2 44422 45409
0 7720 7 1 2 61298 61301
0 7721 7 1 2 61296 7720
0 7722 5 1 1 7721
0 7723 7 14 2 47739 59189
0 7724 5 1 1 61307
0 7725 7 6 2 44423 59475
0 7726 7 1 2 45410 61321
0 7727 5 1 1 7726
0 7728 7 1 2 7724 7727
0 7729 5 2 1 7728
0 7730 7 1 2 45538 61327
0 7731 5 1 1 7730
0 7732 7 3 2 55606 59355
0 7733 5 1 1 61329
0 7734 7 1 2 7731 7733
0 7735 5 1 1 7734
0 7736 7 5 2 46169 53238
0 7737 7 1 2 49267 61332
0 7738 7 1 2 7735 7737
0 7739 5 1 1 7738
0 7740 7 1 2 7722 7739
0 7741 5 1 1 7740
0 7742 7 1 2 61119 7741
0 7743 5 1 1 7742
0 7744 7 1 2 56014 59928
0 7745 7 16 2 42494 42720
0 7746 7 3 2 43700 61337
0 7747 7 6 2 44626 59139
0 7748 7 1 2 61353 61356
0 7749 7 1 2 7744 7748
0 7750 5 1 1 7749
0 7751 7 1 2 7743 7750
0 7752 5 1 1 7751
0 7753 7 1 2 46635 7752
0 7754 5 1 1 7753
0 7755 7 1 2 53239 58868
0 7756 7 2 2 54951 61120
0 7757 7 1 2 59909 61362
0 7758 7 1 2 7755 7757
0 7759 5 1 1 7758
0 7760 7 1 2 7754 7759
0 7761 5 1 1 7760
0 7762 7 1 2 51854 7761
0 7763 5 1 1 7762
0 7764 7 3 2 60994 7602
0 7765 5 17 1 61364
0 7766 7 1 2 51332 60995
0 7767 5 1 1 7766
0 7768 7 2 2 47382 60766
0 7769 7 1 2 7767 61384
0 7770 7 1 2 61367 7769
0 7771 5 1 1 7770
0 7772 7 3 2 44021 44627
0 7773 7 1 2 51546 61386
0 7774 7 1 2 60760 7773
0 7775 5 1 1 7774
0 7776 7 1 2 7771 7775
0 7777 5 1 1 7776
0 7778 7 1 2 59779 7777
0 7779 5 1 1 7778
0 7780 7 1 2 59910 61179
0 7781 5 1 1 7780
0 7782 7 1 2 7779 7781
0 7783 5 1 1 7782
0 7784 7 1 2 42721 7783
0 7785 5 1 1 7784
0 7786 7 9 2 47081 61121
0 7787 7 4 2 49896 61389
0 7788 5 1 1 61398
0 7789 7 1 2 60996 7788
0 7790 5 5 1 7789
0 7791 7 1 2 48783 61402
0 7792 5 1 1 7791
0 7793 7 4 2 43248 44628
0 7794 7 2 2 51547 61407
0 7795 5 1 1 61411
0 7796 7 1 2 7792 7795
0 7797 5 1 1 7796
0 7798 7 1 2 55856 59356
0 7799 7 1 2 7797 7798
0 7800 5 1 1 7799
0 7801 7 1 2 7785 7800
0 7802 5 1 1 7801
0 7803 7 1 2 58713 7802
0 7804 5 1 1 7803
0 7805 7 1 2 45411 53369
0 7806 5 1 1 7805
0 7807 7 1 2 50982 7806
0 7808 7 1 2 61221 7807
0 7809 5 1 1 7808
0 7810 7 1 2 49484 58528
0 7811 5 1 1 7810
0 7812 7 1 2 3804 6645
0 7813 5 1 1 7812
0 7814 7 1 2 47383 60756
0 7815 7 1 2 7813 7814
0 7816 5 1 1 7815
0 7817 7 1 2 7811 7816
0 7818 5 1 1 7817
0 7819 7 5 2 46170 47956
0 7820 7 4 2 44738 61413
0 7821 7 1 2 59829 61418
0 7822 7 1 2 7818 7821
0 7823 5 1 1 7822
0 7824 7 1 2 7809 7823
0 7825 5 1 1 7824
0 7826 7 1 2 61043 7825
0 7827 5 1 1 7826
0 7828 7 1 2 7804 7827
0 7829 5 1 1 7828
0 7830 7 1 2 44177 7829
0 7831 5 1 1 7830
0 7832 7 1 2 49505 60971
0 7833 5 1 1 7832
0 7834 7 3 2 54380 61390
0 7835 5 2 1 61422
0 7836 7 1 2 7833 61425
0 7837 5 1 1 7836
0 7838 7 1 2 59830 7837
0 7839 5 1 1 7838
0 7840 7 16 2 47957 45412
0 7841 7 3 2 59218 61427
0 7842 5 1 1 61443
0 7843 7 1 2 60997 7842
0 7844 5 1 1 7843
0 7845 7 13 2 45539 42722
0 7846 7 10 2 43024 47384
0 7847 7 2 2 59476 61459
0 7848 7 1 2 61446 61469
0 7849 7 1 2 7844 7848
0 7850 5 1 1 7849
0 7851 7 1 2 7839 7850
0 7852 5 1 1 7851
0 7853 7 1 2 43249 7852
0 7854 5 1 1 7853
0 7855 7 1 2 45540 54381
0 7856 7 2 2 60119 7855
0 7857 7 2 2 49506 58076
0 7858 7 1 2 61122 61473
0 7859 7 1 2 61471 7858
0 7860 5 1 1 7859
0 7861 7 1 2 7854 7860
0 7862 5 1 1 7861
0 7863 7 1 2 47740 7862
0 7864 5 1 1 7863
0 7865 7 3 2 59140 61123
0 7866 7 4 2 49268 57011
0 7867 7 1 2 61475 61478
0 7868 7 1 2 60014 7867
0 7869 5 1 1 7868
0 7870 7 1 2 7864 7869
0 7871 5 1 1 7870
0 7872 7 1 2 60562 7871
0 7873 5 1 1 7872
0 7874 7 1 2 48080 57500
0 7875 7 1 2 59946 61014
0 7876 7 1 2 7874 7875
0 7877 7 6 2 47879 57936
0 7878 5 1 1 61482
0 7879 7 1 2 61354 61483
0 7880 7 1 2 7876 7879
0 7881 5 1 1 7880
0 7882 7 1 2 45413 58714
0 7883 5 1 1 7882
0 7884 7 1 2 7520 7883
0 7885 5 3 1 7884
0 7886 7 2 2 44739 59673
0 7887 7 1 2 61105 61491
0 7888 7 1 2 61333 7887
0 7889 7 1 2 61488 7888
0 7890 5 1 1 7889
0 7891 7 1 2 7881 7890
0 7892 5 1 1 7891
0 7893 7 1 2 50983 7892
0 7894 5 1 1 7893
0 7895 7 1 2 7873 7894
0 7896 7 1 2 7831 7895
0 7897 7 1 2 7763 7896
0 7898 7 1 2 7716 7897
0 7899 5 1 1 7898
0 7900 7 1 2 45198 7899
0 7901 5 1 1 7900
0 7902 7 3 2 59780 60972
0 7903 7 1 2 44022 50127
0 7904 5 2 1 7903
0 7905 7 1 2 51200 55313
0 7906 5 3 1 7905
0 7907 7 1 2 61496 61498
0 7908 5 1 1 7907
0 7909 7 1 2 46171 7908
0 7910 5 1 1 7909
0 7911 7 1 2 55372 58414
0 7912 5 3 1 7911
0 7913 7 1 2 7910 61501
0 7914 5 1 1 7913
0 7915 7 1 2 61493 7914
0 7916 5 1 1 7915
0 7917 7 6 2 47082 47958
0 7918 7 11 2 44740 61504
0 7919 7 12 2 46172 49269
0 7920 5 1 1 61521
0 7921 7 1 2 49590 61522
0 7922 5 1 1 7921
0 7923 7 1 2 45414 58480
0 7924 5 1 1 7923
0 7925 7 1 2 7922 7924
0 7926 5 1 1 7925
0 7927 7 1 2 59831 7926
0 7928 5 1 1 7927
0 7929 7 2 2 42723 49270
0 7930 5 2 1 61533
0 7931 7 2 2 46173 50934
0 7932 5 2 1 61537
0 7933 7 1 2 61535 61539
0 7934 5 2 1 7933
0 7935 7 2 2 50828 61541
0 7936 5 1 1 61543
0 7937 7 1 2 46174 60816
0 7938 5 3 1 7937
0 7939 7 1 2 50749 55001
0 7940 5 1 1 7939
0 7941 7 1 2 61545 7940
0 7942 5 1 1 7941
0 7943 7 1 2 48784 7942
0 7944 5 1 1 7943
0 7945 7 1 2 7936 7944
0 7946 5 1 1 7945
0 7947 7 1 2 60154 59564
0 7948 7 1 2 7946 7947
0 7949 5 1 1 7948
0 7950 7 1 2 7928 7949
0 7951 5 1 1 7950
0 7952 7 1 2 61510 7951
0 7953 5 1 1 7952
0 7954 7 1 2 7916 7953
0 7955 5 1 1 7954
0 7956 7 1 2 48557 7955
0 7957 5 1 1 7956
0 7958 7 2 2 47623 56104
0 7959 7 2 2 61391 61548
0 7960 7 1 2 61299 61550
0 7961 5 1 1 7960
0 7962 7 3 2 48892 51134
0 7963 7 8 2 44304 48081
0 7964 7 1 2 57937 61555
0 7965 7 1 2 61552 7964
0 7966 5 1 1 7965
0 7967 7 1 2 7961 7966
0 7968 5 1 1 7967
0 7969 7 1 2 48558 7968
0 7970 5 1 1 7969
0 7971 7 6 2 44305 44629
0 7972 7 2 2 48082 61563
0 7973 7 2 2 55473 61553
0 7974 7 1 2 61569 61571
0 7975 5 1 1 7974
0 7976 7 1 2 7970 7975
0 7977 5 1 1 7976
0 7978 7 1 2 55565 7977
0 7979 5 1 1 7978
0 7980 7 1 2 53493 55002
0 7981 5 2 1 7980
0 7982 7 1 2 48785 61544
0 7983 5 1 1 7982
0 7984 7 1 2 61573 7983
0 7985 5 1 1 7984
0 7986 7 1 2 61494 7985
0 7987 5 1 1 7986
0 7988 7 1 2 7979 7987
0 7989 7 1 2 7957 7988
0 7990 5 1 1 7989
0 7991 7 1 2 61044 7990
0 7992 5 1 1 7991
0 7993 7 1 2 47083 57836
0 7994 7 1 2 60514 7993
0 7995 5 1 1 7994
0 7996 7 2 2 54132 59190
0 7997 7 9 2 47741 45415
0 7998 7 1 2 54952 61577
0 7999 7 1 2 61575 7998
0 8000 5 1 1 7999
0 8001 7 1 2 7995 8000
0 8002 5 1 1 8001
0 8003 7 1 2 51855 8002
0 8004 5 1 1 8003
0 8005 7 3 2 44424 55705
0 8006 7 2 2 43701 55436
0 8007 7 9 2 45698 47624
0 8008 7 1 2 54953 61591
0 8009 7 1 2 61589 8008
0 8010 7 1 2 61586 8009
0 8011 5 1 1 8010
0 8012 7 1 2 8004 8011
0 8013 5 1 1 8012
0 8014 7 1 2 45541 8013
0 8015 5 1 1 8014
0 8016 7 1 2 60563 61328
0 8017 5 1 1 8016
0 8018 7 2 2 44306 61578
0 8019 7 1 2 60888 61600
0 8020 5 1 1 8019
0 8021 7 1 2 8017 8020
0 8022 5 1 1 8021
0 8023 7 4 2 41988 46441
0 8024 7 3 2 47385 61602
0 8025 7 1 2 55097 61606
0 8026 7 1 2 8022 8025
0 8027 5 1 1 8026
0 8028 7 1 2 8015 8027
0 8029 5 1 1 8028
0 8030 7 1 2 45984 8029
0 8031 5 1 1 8030
0 8032 7 1 2 45416 61227
0 8033 5 1 1 8032
0 8034 7 1 2 60941 8033
0 8035 5 1 1 8034
0 8036 7 5 2 47386 54954
0 8037 7 1 2 53195 61609
0 8038 7 1 2 8035 8037
0 8039 5 1 1 8038
0 8040 7 1 2 8031 8039
0 8041 5 1 1 8040
0 8042 7 1 2 61124 8041
0 8043 5 1 1 8042
0 8044 7 2 2 59008 60516
0 8045 7 2 2 51135 60623
0 8046 7 2 2 44552 60344
0 8047 7 1 2 61616 61618
0 8048 7 1 2 61614 8047
0 8049 5 1 1 8048
0 8050 7 1 2 8043 8049
0 8051 5 1 1 8050
0 8052 7 1 2 56650 8051
0 8053 5 1 1 8052
0 8054 7 1 2 5466 5492
0 8055 5 2 1 8054
0 8056 7 1 2 61088 61229
0 8057 7 1 2 61620 8056
0 8058 5 1 1 8057
0 8059 7 1 2 60942 8058
0 8060 5 1 1 8059
0 8061 7 1 2 42724 8060
0 8062 5 1 1 8061
0 8063 7 4 2 59009 60624
0 8064 7 1 2 50630 54462
0 8065 7 1 2 61622 8064
0 8066 5 1 1 8065
0 8067 7 1 2 8062 8066
0 8068 5 1 1 8067
0 8069 7 1 2 61217 8068
0 8070 5 1 1 8069
0 8071 7 3 2 46442 54413
0 8072 7 10 2 45699 46175
0 8073 7 1 2 47387 61629
0 8074 7 1 2 61626 8073
0 8075 7 22 2 41989 60625
0 8076 5 1 1 61639
0 8077 7 6 2 44741 48931
0 8078 7 1 2 61640 61661
0 8079 7 1 2 8074 8078
0 8080 5 1 1 8079
0 8081 7 1 2 8070 8080
0 8082 5 1 1 8081
0 8083 7 1 2 45417 8082
0 8084 5 1 1 8083
0 8085 7 2 2 41990 60964
0 8086 7 2 2 61627 61667
0 8087 7 5 2 44742 51559
0 8088 7 1 2 47388 61288
0 8089 7 1 2 61671 8088
0 8090 7 1 2 61669 8089
0 8091 5 1 1 8090
0 8092 7 1 2 8084 8091
0 8093 5 1 1 8092
0 8094 7 1 2 42495 8093
0 8095 5 1 1 8094
0 8096 7 2 2 41991 61125
0 8097 7 1 2 58408 61676
0 8098 7 1 2 61576 8097
0 8099 7 1 2 61489 8098
0 8100 5 1 1 8099
0 8101 7 1 2 8095 8100
0 8102 5 1 1 8101
0 8103 7 1 2 50057 8102
0 8104 5 1 1 8103
0 8105 7 1 2 58421 58447
0 8106 5 1 1 8105
0 8107 7 1 2 55373 8106
0 8108 5 1 1 8107
0 8109 7 1 2 61546 8108
0 8110 5 1 1 8109
0 8111 7 1 2 48559 8110
0 8112 5 1 1 8111
0 8113 7 3 2 49029 57343
0 8114 5 2 1 61678
0 8115 7 1 2 50935 61679
0 8116 5 2 1 8115
0 8117 7 1 2 8112 61683
0 8118 5 1 1 8117
0 8119 7 1 2 61495 8118
0 8120 5 1 1 8119
0 8121 7 4 2 44023 49507
0 8122 5 3 1 61685
0 8123 7 6 2 47389 53738
0 8124 5 1 1 61692
0 8125 7 1 2 42725 8124
0 8126 5 1 1 8125
0 8127 7 1 2 61689 8126
0 8128 5 2 1 8127
0 8129 7 1 2 61180 61698
0 8130 5 1 1 8129
0 8131 7 3 2 48083 61387
0 8132 7 5 2 43025 43702
0 8133 5 2 1 61703
0 8134 7 2 2 42496 61704
0 8135 7 1 2 61700 61710
0 8136 5 1 1 8135
0 8137 7 1 2 8130 8136
0 8138 5 1 1 8137
0 8139 7 1 2 50750 8138
0 8140 5 1 1 8139
0 8141 7 1 2 48786 54227
0 8142 7 1 2 60973 8141
0 8143 5 2 1 8142
0 8144 7 4 2 45985 54092
0 8145 7 3 2 44743 54644
0 8146 7 1 2 61714 61718
0 8147 5 1 1 8146
0 8148 7 1 2 61712 8147
0 8149 5 1 1 8148
0 8150 7 1 2 48560 8149
0 8151 5 1 1 8150
0 8152 7 1 2 47390 61423
0 8153 5 1 1 8152
0 8154 7 1 2 8151 8153
0 8155 5 1 1 8154
0 8156 7 1 2 50829 8155
0 8157 5 1 1 8156
0 8158 7 1 2 46176 49523
0 8159 5 3 1 8158
0 8160 7 1 2 61181 61721
0 8161 5 1 1 8160
0 8162 7 7 2 43703 60345
0 8163 7 1 2 49583 61724
0 8164 5 1 1 8163
0 8165 7 1 2 8161 8164
0 8166 5 1 1 8165
0 8167 7 1 2 50751 8166
0 8168 5 1 1 8167
0 8169 7 2 2 48084 54228
0 8170 7 4 2 44178 44630
0 8171 7 1 2 51369 61733
0 8172 7 1 2 61731 8171
0 8173 5 1 1 8172
0 8174 7 1 2 8168 8173
0 8175 5 1 1 8174
0 8176 7 1 2 48561 8175
0 8177 5 1 1 8176
0 8178 7 1 2 8157 8177
0 8179 7 1 2 8140 8178
0 8180 5 1 1 8179
0 8181 7 1 2 59832 8180
0 8182 5 1 1 8181
0 8183 7 1 2 8120 8182
0 8184 5 1 1 8183
0 8185 7 1 2 58715 8184
0 8186 5 1 1 8185
0 8187 7 1 2 8104 8186
0 8188 7 1 2 8053 8187
0 8189 7 1 2 7992 8188
0 8190 7 1 2 7901 8189
0 8191 5 1 1 8190
0 8192 7 1 2 47219 8191
0 8193 5 1 1 8192
0 8194 7 8 2 47625 48787
0 8195 7 7 2 58180 61737
0 8196 7 2 2 56208 61745
0 8197 5 1 1 61752
0 8198 7 3 2 47516 53753
0 8199 5 1 1 61754
0 8200 7 1 2 59833 61755
0 8201 5 1 1 8200
0 8202 7 1 2 8197 8201
0 8203 5 1 1 8202
0 8204 7 1 2 46636 8203
0 8205 5 1 1 8204
0 8206 7 2 2 61078 61738
0 8207 7 1 2 53355 60422
0 8208 7 1 2 61757 8207
0 8209 5 1 1 8208
0 8210 7 1 2 8205 8209
0 8211 5 1 1 8210
0 8212 7 1 2 61182 8211
0 8213 5 1 1 8212
0 8214 7 2 2 59834 60346
0 8215 7 1 2 58962 61759
0 8216 5 1 1 8215
0 8217 7 1 2 8213 8216
0 8218 5 1 1 8217
0 8219 7 1 2 58716 8218
0 8220 5 1 1 8219
0 8221 7 3 2 47880 59191
0 8222 7 7 2 44425 56229
0 8223 7 2 2 61761 61764
0 8224 7 3 2 42726 51333
0 8225 7 1 2 58883 60347
0 8226 7 1 2 61773 8225
0 8227 5 1 1 8226
0 8228 7 3 2 46443 51168
0 8229 7 1 2 50752 61419
0 8230 7 1 2 61776 8229
0 8231 5 1 1 8230
0 8232 7 1 2 8227 8231
0 8233 5 1 1 8232
0 8234 7 1 2 61771 8233
0 8235 5 1 1 8234
0 8236 7 2 2 58181 59748
0 8237 7 6 2 46177 51334
0 8238 5 1 1 61781
0 8239 7 1 2 61502 8238
0 8240 5 1 1 8239
0 8241 7 1 2 61126 8240
0 8242 7 1 2 61779 8241
0 8243 5 1 1 8242
0 8244 7 3 2 43444 51136
0 8245 7 4 2 50058 60348
0 8246 7 1 2 59357 61790
0 8247 7 1 2 61787 8246
0 8248 5 1 1 8247
0 8249 7 1 2 8243 8248
0 8250 5 1 1 8249
0 8251 7 1 2 58717 8250
0 8252 5 1 1 8251
0 8253 7 1 2 8235 8252
0 8254 5 1 1 8253
0 8255 7 1 2 45418 8254
0 8256 5 1 1 8255
0 8257 7 3 2 56259 60349
0 8258 7 1 2 54210 58731
0 8259 7 1 2 61794 8258
0 8260 5 1 1 8259
0 8261 7 3 2 47959 57628
0 8262 7 4 2 44744 45419
0 8263 7 4 2 45986 61800
0 8264 7 1 2 60555 61804
0 8265 7 1 2 61797 8264
0 8266 5 1 1 8265
0 8267 7 1 2 8260 8266
0 8268 5 1 1 8267
0 8269 7 1 2 59835 8268
0 8270 5 1 1 8269
0 8271 7 2 2 46178 60097
0 8272 7 2 2 45542 60790
0 8273 7 2 2 57629 61127
0 8274 7 1 2 61810 61812
0 8275 7 1 2 61808 8274
0 8276 5 1 1 8275
0 8277 7 1 2 8270 8276
0 8278 5 1 1 8277
0 8279 7 1 2 55566 8278
0 8280 5 1 1 8279
0 8281 7 4 2 44553 59010
0 8282 7 1 2 59959 60626
0 8283 7 1 2 61183 8282
0 8284 7 1 2 61814 8283
0 8285 5 1 1 8284
0 8286 7 10 2 46179 48788
0 8287 5 2 1 61818
0 8288 7 1 2 60974 61819
0 8289 7 1 2 60691 8288
0 8290 5 1 1 8289
0 8291 7 1 2 8285 8290
0 8292 5 1 1 8291
0 8293 7 1 2 50830 8292
0 8294 5 1 1 8293
0 8295 7 1 2 8280 8294
0 8296 7 1 2 8256 8295
0 8297 7 1 2 8220 8296
0 8298 5 1 1 8297
0 8299 7 1 2 57179 8298
0 8300 5 1 1 8299
0 8301 7 4 2 44307 48562
0 8302 7 1 2 46444 50831
0 8303 5 7 1 8302
0 8304 7 2 2 60210 61834
0 8305 5 1 1 61841
0 8306 7 2 2 57996 8305
0 8307 7 2 2 44554 61843
0 8308 7 2 2 53850 57133
0 8309 7 1 2 47742 59011
0 8310 7 1 2 61847 8309
0 8311 7 1 2 61845 8310
0 8312 5 1 1 8311
0 8313 7 1 2 44179 60590
0 8314 5 1 1 8313
0 8315 7 1 2 51747 60582
0 8316 5 1 1 8315
0 8317 7 1 2 8314 8316
0 8318 5 1 1 8317
0 8319 7 1 2 41992 8318
0 8320 5 1 1 8319
0 8321 7 10 2 42149 43250
0 8322 7 4 2 54478 61849
0 8323 7 2 2 60413 61859
0 8324 7 1 2 57767 61863
0 8325 5 1 1 8324
0 8326 7 1 2 8320 8325
0 8327 5 1 1 8326
0 8328 7 4 2 50936 53240
0 8329 7 1 2 42727 61865
0 8330 7 1 2 8327 8329
0 8331 5 1 1 8330
0 8332 7 1 2 8312 8331
0 8333 5 1 1 8332
0 8334 7 1 2 60350 8333
0 8335 5 1 1 8334
0 8336 7 4 2 41993 43251
0 8337 7 1 2 50210 59452
0 8338 7 1 2 61869 8337
0 8339 7 7 2 45987 47960
0 8340 7 7 2 44745 61873
0 8341 7 1 2 54028 61045
0 8342 7 1 2 61880 8341
0 8343 7 1 2 8338 8342
0 8344 5 1 1 8343
0 8345 7 1 2 8335 8344
0 8346 5 1 1 8345
0 8347 7 1 2 61830 8346
0 8348 5 1 1 8347
0 8349 7 1 2 8300 8348
0 8350 7 1 2 8193 8349
0 8351 7 1 2 7609 8350
0 8352 5 1 1 8351
0 8353 7 1 2 45056 8352
0 8354 5 1 1 8353
0 8355 7 4 2 59141 60018
0 8356 7 1 2 60271 61887
0 8357 5 1 1 8356
0 8358 7 1 2 2249 60264
0 8359 5 2 1 8358
0 8360 7 3 2 45420 61308
0 8361 5 1 1 61893
0 8362 7 1 2 61891 61894
0 8363 5 1 1 8362
0 8364 7 1 2 8357 8363
0 8365 5 1 1 8364
0 8366 7 1 2 47517 8365
0 8367 5 1 1 8366
0 8368 7 3 2 49200 60627
0 8369 7 1 2 51995 59960
0 8370 7 1 2 61896 8369
0 8371 5 1 1 8370
0 8372 7 1 2 8367 8371
0 8373 5 2 1 8372
0 8374 7 1 2 45199 61899
0 8375 5 1 1 8374
0 8376 7 2 2 48994 54955
0 8377 7 2 2 43445 47518
0 8378 7 1 2 60628 61903
0 8379 7 1 2 61901 8378
0 8380 5 1 1 8379
0 8381 7 1 2 8375 8380
0 8382 5 1 1 8381
0 8383 7 1 2 47391 8382
0 8384 5 1 1 8383
0 8385 7 1 2 43857 52359
0 8386 5 2 1 8385
0 8387 7 1 2 54956 58504
0 8388 7 1 2 60657 8387
0 8389 7 1 2 61905 8388
0 8390 5 1 1 8389
0 8391 7 1 2 8384 8390
0 8392 5 1 1 8391
0 8393 7 1 2 43704 8392
0 8394 5 1 1 8393
0 8395 7 1 2 53091 54903
0 8396 5 1 1 8395
0 8397 7 2 2 58573 8396
0 8398 7 1 2 49201 61907
0 8399 5 1 1 8398
0 8400 7 1 2 48995 52053
0 8401 7 1 2 58610 8400
0 8402 5 1 1 8401
0 8403 7 1 2 8399 8402
0 8404 5 1 1 8403
0 8405 7 1 2 44024 8404
0 8406 5 1 1 8405
0 8407 7 3 2 43858 49151
0 8408 5 1 1 61909
0 8409 7 1 2 54211 61910
0 8410 5 1 1 8409
0 8411 7 1 2 8406 8410
0 8412 5 1 1 8411
0 8413 7 2 2 60629 8412
0 8414 7 1 2 54414 61912
0 8415 5 1 1 8414
0 8416 7 1 2 8394 8415
0 8417 5 1 1 8416
0 8418 7 1 2 42497 8417
0 8419 5 1 1 8418
0 8420 7 1 2 52892 61322
0 8421 5 1 1 8420
0 8422 7 1 2 59625 60658
0 8423 5 1 1 8422
0 8424 7 1 2 8421 8423
0 8425 5 1 1 8424
0 8426 7 1 2 47519 8425
0 8427 5 1 1 8426
0 8428 7 5 2 44180 49741
0 8429 5 1 1 61914
0 8430 7 2 2 59623 8429
0 8431 5 1 1 61919
0 8432 7 1 2 61309 8431
0 8433 5 1 1 8432
0 8434 7 1 2 8427 8433
0 8435 5 1 1 8434
0 8436 7 1 2 59057 8435
0 8437 5 1 1 8436
0 8438 7 1 2 45988 57134
0 8439 7 1 2 61913 8438
0 8440 5 1 1 8439
0 8441 7 1 2 8437 8440
0 8442 7 1 2 8419 8441
0 8443 5 1 1 8442
0 8444 7 1 2 60351 8443
0 8445 5 1 1 8444
0 8446 7 1 2 47392 61900
0 8447 5 1 1 8446
0 8448 7 4 2 46820 47220
0 8449 7 1 2 49508 59142
0 8450 7 1 2 61921 8449
0 8451 5 1 1 8450
0 8452 7 5 2 46445 44308
0 8453 7 4 2 43446 61925
0 8454 7 1 2 45421 56269
0 8455 7 1 2 61930 8454
0 8456 5 1 1 8455
0 8457 7 1 2 8451 8456
0 8458 5 1 1 8457
0 8459 7 1 2 47520 8458
0 8460 5 1 1 8459
0 8461 7 1 2 57714 61897
0 8462 5 1 1 8461
0 8463 7 1 2 8460 8462
0 8464 5 1 1 8463
0 8465 7 1 2 46180 8464
0 8466 5 1 1 8465
0 8467 7 1 2 8447 8466
0 8468 5 1 1 8467
0 8469 7 1 2 45200 8468
0 8470 5 1 1 8469
0 8471 7 1 2 57087 61693
0 8472 5 2 1 8471
0 8473 7 2 2 44025 55314
0 8474 5 3 1 61936
0 8475 7 1 2 47221 52360
0 8476 7 1 2 61938 8475
0 8477 5 1 1 8476
0 8478 7 1 2 61934 8477
0 8479 5 1 1 8478
0 8480 7 1 2 61310 8479
0 8481 5 1 1 8480
0 8482 7 1 2 47222 49012
0 8483 7 1 2 61888 8482
0 8484 5 1 1 8483
0 8485 7 1 2 8481 8484
0 8486 5 1 1 8485
0 8487 7 1 2 46181 8486
0 8488 5 1 1 8487
0 8489 7 1 2 8470 8488
0 8490 5 1 1 8489
0 8491 7 1 2 61184 8490
0 8492 5 1 1 8491
0 8493 7 1 2 8445 8492
0 8494 5 1 1 8493
0 8495 7 1 2 46637 8494
0 8496 5 1 1 8495
0 8497 7 2 2 57605 59143
0 8498 5 2 1 61941
0 8499 7 1 2 59192 60414
0 8500 5 2 1 8499
0 8501 7 1 2 61943 61945
0 8502 5 2 1 8501
0 8503 7 1 2 50603 61947
0 8504 5 1 1 8503
0 8505 7 5 2 44426 48563
0 8506 7 2 2 59878 61949
0 8507 7 1 2 46821 61954
0 8508 5 2 1 8507
0 8509 7 1 2 8504 61956
0 8510 5 1 1 8509
0 8511 7 1 2 46182 8510
0 8512 5 1 1 8511
0 8513 7 1 2 55437 60630
0 8514 7 1 2 58804 8513
0 8515 5 1 1 8514
0 8516 7 1 2 8512 8515
0 8517 5 1 1 8516
0 8518 7 1 2 43859 8517
0 8519 5 1 1 8518
0 8520 7 3 2 43860 50984
0 8521 7 2 2 52925 61958
0 8522 5 1 1 61961
0 8523 7 1 2 49789 54108
0 8524 5 3 1 8523
0 8525 7 1 2 8522 61963
0 8526 5 3 1 8525
0 8527 7 1 2 61323 61966
0 8528 5 1 1 8527
0 8529 7 2 2 57715 60631
0 8530 7 1 2 51489 61969
0 8531 5 1 1 8530
0 8532 7 1 2 8528 8531
0 8533 5 1 1 8532
0 8534 7 1 2 42728 8533
0 8535 5 1 1 8534
0 8536 7 2 2 48564 59463
0 8537 7 4 2 43026 60607
0 8538 7 1 2 56936 61973
0 8539 7 1 2 61971 8538
0 8540 5 1 1 8539
0 8541 7 1 2 8535 8540
0 8542 7 1 2 8519 8541
0 8543 5 1 1 8542
0 8544 7 1 2 43705 8543
0 8545 5 1 1 8544
0 8546 7 2 2 47743 52376
0 8547 7 2 2 51965 52502
0 8548 7 1 2 59338 61979
0 8549 7 1 2 61977 8548
0 8550 5 1 1 8549
0 8551 7 1 2 8545 8550
0 8552 5 1 1 8551
0 8553 7 1 2 60352 8552
0 8554 5 1 1 8553
0 8555 7 2 2 52743 52844
0 8556 7 2 2 57853 61981
0 8557 7 2 2 46822 57905
0 8558 7 1 2 61092 61985
0 8559 7 1 2 61983 8558
0 8560 5 1 1 8559
0 8561 7 1 2 8554 8560
0 8562 5 1 1 8561
0 8563 7 1 2 44181 8562
0 8564 5 1 1 8563
0 8565 7 1 2 44026 61908
0 8566 5 1 1 8565
0 8567 7 6 2 42729 49742
0 8568 5 2 1 61987
0 8569 7 1 2 43861 61988
0 8570 5 1 1 8569
0 8571 7 2 2 8566 8570
0 8572 5 3 1 61995
0 8573 7 1 2 61218 61997
0 8574 5 1 1 8573
0 8575 7 3 2 55367 57557
0 8576 5 2 1 62000
0 8577 7 1 2 46183 62001
0 8578 5 1 1 8577
0 8579 7 2 2 50543 52976
0 8580 5 1 1 62005
0 8581 7 1 2 8578 8580
0 8582 5 1 1 8581
0 8583 7 1 2 61511 8582
0 8584 5 1 1 8583
0 8585 7 1 2 8574 8584
0 8586 5 1 1 8585
0 8587 7 1 2 49072 8586
0 8588 5 1 1 8587
0 8589 7 7 2 54158 60353
0 8590 7 1 2 55003 62007
0 8591 5 1 1 8590
0 8592 7 3 2 52028 61128
0 8593 7 2 2 50985 62014
0 8594 7 1 2 47084 62017
0 8595 5 1 1 8594
0 8596 7 1 2 8591 8595
0 8597 5 1 1 8596
0 8598 7 1 2 45201 8597
0 8599 5 1 1 8598
0 8600 7 1 2 8588 8599
0 8601 5 1 1 8600
0 8602 7 1 2 61311 8601
0 8603 5 1 1 8602
0 8604 7 2 2 48996 61476
0 8605 7 1 2 53395 57701
0 8606 7 1 2 62019 8605
0 8607 5 1 1 8606
0 8608 7 1 2 8603 8607
0 8609 7 1 2 8564 8608
0 8610 5 1 1 8609
0 8611 7 1 2 45989 8610
0 8612 5 1 1 8611
0 8613 7 4 2 42498 44631
0 8614 7 1 2 50604 61324
0 8615 5 1 1 8614
0 8616 7 1 2 61946 8615
0 8617 5 1 1 8616
0 8618 7 1 2 43027 8617
0 8619 5 1 1 8618
0 8620 7 1 2 59636 61312
0 8621 5 1 1 8620
0 8622 7 1 2 61957 8621
0 8623 7 1 2 8619 8622
0 8624 5 1 1 8623
0 8625 7 1 2 56799 8624
0 8626 5 1 1 8625
0 8627 7 2 2 49103 60632
0 8628 7 1 2 61974 62025
0 8629 5 1 1 8628
0 8630 7 2 2 59172 60019
0 8631 5 1 1 62027
0 8632 7 2 2 49073 61313
0 8633 5 1 1 62029
0 8634 7 1 2 8631 8633
0 8635 5 1 1 8634
0 8636 7 1 2 49743 8635
0 8637 5 2 1 8636
0 8638 7 1 2 46823 59173
0 8639 5 1 1 8638
0 8640 7 1 2 60664 8639
0 8641 5 1 1 8640
0 8642 7 1 2 50544 8641
0 8643 5 1 1 8642
0 8644 7 1 2 62031 8643
0 8645 5 1 1 8644
0 8646 7 1 2 43862 8645
0 8647 5 1 1 8646
0 8648 7 1 2 8629 8647
0 8649 7 1 2 8626 8648
0 8650 5 1 1 8649
0 8651 7 1 2 42730 8650
0 8652 5 1 1 8651
0 8653 7 1 2 44427 56866
0 8654 7 2 2 60922 8653
0 8655 7 1 2 52090 62033
0 8656 5 1 1 8655
0 8657 7 5 2 53028 55364
0 8658 5 1 1 62035
0 8659 7 1 2 49030 62036
0 8660 5 2 1 8659
0 8661 7 1 2 49074 54861
0 8662 5 1 1 8661
0 8663 7 1 2 62040 8662
0 8664 5 1 1 8663
0 8665 7 1 2 60659 8664
0 8666 5 1 1 8665
0 8667 7 1 2 8656 8666
0 8668 5 1 1 8667
0 8669 7 1 2 43863 8668
0 8670 5 1 1 8669
0 8671 7 3 2 44027 59599
0 8672 7 1 2 43447 55228
0 8673 7 1 2 61978 8672
0 8674 7 1 2 62042 8673
0 8675 5 1 1 8674
0 8676 7 1 2 47085 8675
0 8677 7 1 2 8670 8676
0 8678 7 1 2 8652 8677
0 8679 5 1 1 8678
0 8680 7 1 2 50986 61314
0 8681 5 1 1 8680
0 8682 7 3 2 46824 60923
0 8683 7 1 2 58869 62045
0 8684 5 1 1 8683
0 8685 7 1 2 8681 8684
0 8686 5 1 1 8685
0 8687 7 1 2 45202 8686
0 8688 5 1 1 8687
0 8689 7 1 2 46446 62030
0 8690 5 1 1 8689
0 8691 7 1 2 62032 8690
0 8692 7 1 2 8688 8691
0 8693 5 1 1 8692
0 8694 7 1 2 52029 8693
0 8695 5 1 1 8694
0 8696 7 1 2 47393 59961
0 8697 7 1 2 62026 8696
0 8698 5 1 1 8697
0 8699 7 1 2 8695 8698
0 8700 5 1 1 8699
0 8701 7 1 2 51996 8700
0 8702 5 1 1 8701
0 8703 7 1 2 43706 8702
0 8704 5 1 1 8703
0 8705 7 1 2 48085 8704
0 8706 7 1 2 8679 8705
0 8707 5 1 1 8706
0 8708 7 1 2 54212 57438
0 8709 7 2 2 43707 52953
0 8710 7 1 2 60660 62048
0 8711 7 1 2 8708 8710
0 8712 5 1 1 8711
0 8713 7 1 2 8707 8712
0 8714 5 1 1 8713
0 8715 7 1 2 62021 8714
0 8716 5 1 1 8715
0 8717 7 1 2 8612 8716
0 8718 5 1 1 8717
0 8719 7 1 2 43252 8718
0 8720 5 1 1 8719
0 8721 7 1 2 51078 59058
0 8722 5 1 1 8721
0 8723 7 2 2 53241 60272
0 8724 7 1 2 52091 62050
0 8725 5 1 1 8724
0 8726 7 1 2 8722 8725
0 8727 5 1 1 8726
0 8728 7 2 2 56184 59477
0 8729 5 1 1 62052
0 8730 7 1 2 8727 62053
0 8731 5 1 1 8730
0 8732 7 3 2 44028 60273
0 8733 5 1 1 62054
0 8734 7 1 2 51997 54213
0 8735 5 1 1 8734
0 8736 7 2 2 8733 8735
0 8737 5 2 1 62057
0 8738 7 2 2 48565 62059
0 8739 5 2 1 62061
0 8740 7 1 2 53242 61315
0 8741 7 1 2 62062 8740
0 8742 5 1 1 8741
0 8743 7 1 2 8731 8742
0 8744 5 1 1 8743
0 8745 7 1 2 60354 8744
0 8746 5 1 1 8745
0 8747 7 5 2 47394 47961
0 8748 7 4 2 51049 62065
0 8749 7 2 2 59144 62070
0 8750 7 3 2 52030 52503
0 8751 7 1 2 60155 62076
0 8752 7 1 2 62074 8751
0 8753 5 1 1 8752
0 8754 7 1 2 8746 8753
0 8755 5 1 1 8754
0 8756 7 1 2 50832 8755
0 8757 5 1 1 8756
0 8758 7 3 2 48566 60355
0 8759 7 1 2 44029 61948
0 8760 7 1 2 62051 8759
0 8761 5 1 1 8760
0 8762 7 11 2 42731 53243
0 8763 7 1 2 49509 61970
0 8764 7 1 2 62082 8763
0 8765 5 1 1 8764
0 8766 7 1 2 8761 8765
0 8767 5 1 1 8766
0 8768 7 1 2 62079 8767
0 8769 5 1 1 8768
0 8770 7 1 2 8757 8769
0 8771 7 1 2 8720 8770
0 8772 7 1 2 8496 8771
0 8773 5 1 1 8772
0 8774 7 1 2 45543 8773
0 8775 5 1 1 8774
0 8776 7 5 2 49271 52031
0 8777 7 2 2 49152 57208
0 8778 7 1 2 62093 62098
0 8779 5 1 1 8778
0 8780 7 2 2 49272 56817
0 8781 5 1 1 62100
0 8782 7 1 2 49333 57475
0 8783 5 1 1 8782
0 8784 7 4 2 47395 52977
0 8785 7 1 2 57370 62102
0 8786 5 2 1 8785
0 8787 7 1 2 43708 62106
0 8788 5 1 1 8787
0 8789 7 1 2 46184 8788
0 8790 7 1 2 8783 8789
0 8791 5 1 1 8790
0 8792 7 1 2 8781 8791
0 8793 5 1 1 8792
0 8794 7 1 2 45990 8793
0 8795 5 1 1 8794
0 8796 7 1 2 8779 8795
0 8797 5 1 1 8796
0 8798 7 1 2 61129 8797
0 8799 5 1 1 8798
0 8800 7 4 2 42499 51998
0 8801 5 2 1 62108
0 8802 7 1 2 55374 61911
0 8803 5 1 1 8802
0 8804 7 1 2 62112 8803
0 8805 5 1 1 8804
0 8806 7 1 2 46447 8805
0 8807 5 1 1 8806
0 8808 7 3 2 43028 58367
0 8809 5 2 1 62114
0 8810 7 1 2 60274 62115
0 8811 5 1 1 8810
0 8812 7 1 2 8807 8811
0 8813 5 1 1 8812
0 8814 7 1 2 43709 8813
0 8815 5 1 1 8814
0 8816 7 2 2 49510 55567
0 8817 5 1 1 62119
0 8818 7 2 2 42500 62120
0 8819 7 1 2 60275 62121
0 8820 5 1 1 8819
0 8821 7 1 2 8815 8820
0 8822 5 1 1 8821
0 8823 7 1 2 47396 8822
0 8824 5 1 1 8823
0 8825 7 1 2 53530 54029
0 8826 5 1 1 8825
0 8827 7 1 2 49957 8826
0 8828 5 1 1 8827
0 8829 7 1 2 51999 8828
0 8830 5 1 1 8829
0 8831 7 1 2 53244 8830
0 8832 5 1 1 8831
0 8833 7 1 2 58512 8832
0 8834 7 1 2 8824 8833
0 8835 5 1 1 8834
0 8836 7 1 2 60356 8835
0 8837 5 1 1 8836
0 8838 7 1 2 8799 8837
0 8839 5 1 1 8838
0 8840 7 1 2 45203 8839
0 8841 5 1 1 8840
0 8842 7 16 2 44632 48567
0 8843 7 3 2 51169 51966
0 8844 5 1 1 62139
0 8845 7 1 2 2988 62140
0 8846 5 1 1 8845
0 8847 7 2 2 55098 58968
0 8848 5 1 1 62142
0 8849 7 1 2 8846 8848
0 8850 5 1 1 8849
0 8851 7 1 2 50937 8850
0 8852 5 1 1 8851
0 8853 7 1 2 47223 53419
0 8854 5 2 1 8853
0 8855 7 1 2 53092 55166
0 8856 7 1 2 62144 8855
0 8857 5 1 1 8856
0 8858 7 1 2 53245 8857
0 8859 5 1 1 8858
0 8860 7 1 2 8852 8859
0 8861 5 1 1 8860
0 8862 7 1 2 44182 8861
0 8863 5 1 1 8862
0 8864 7 2 2 49485 58611
0 8865 7 1 2 50451 52032
0 8866 5 1 1 8865
0 8867 7 1 2 55062 8866
0 8868 5 1 1 8867
0 8869 7 1 2 62146 8868
0 8870 5 1 1 8869
0 8871 7 1 2 8863 8870
0 8872 5 1 1 8871
0 8873 7 1 2 43253 8872
0 8874 5 1 1 8873
0 8875 7 3 2 44183 56260
0 8876 7 1 2 55229 62148
0 8877 5 1 1 8876
0 8878 7 1 2 54159 60718
0 8879 5 1 1 8878
0 8880 7 1 2 46185 8879
0 8881 7 1 2 8877 8880
0 8882 5 1 1 8881
0 8883 7 1 2 53995 60700
0 8884 5 1 1 8883
0 8885 7 1 2 54932 60719
0 8886 5 1 1 8885
0 8887 7 1 2 42732 8886
0 8888 7 1 2 8884 8887
0 8889 5 1 1 8888
0 8890 7 1 2 49121 8889
0 8891 7 1 2 8882 8890
0 8892 5 1 1 8891
0 8893 7 1 2 8874 8892
0 8894 5 1 1 8893
0 8895 7 1 2 48086 8894
0 8896 5 1 1 8895
0 8897 7 2 2 44184 57433
0 8898 7 1 2 54542 62151
0 8899 5 1 1 8898
0 8900 7 1 2 8896 8899
0 8901 5 1 1 8900
0 8902 7 1 2 62123 8901
0 8903 5 1 1 8902
0 8904 7 1 2 8841 8903
0 8905 5 1 1 8904
0 8906 7 1 2 55894 8905
0 8907 5 1 1 8906
0 8908 7 4 2 45991 47521
0 8909 7 1 2 61505 62153
0 8910 7 1 2 62006 8909
0 8911 5 1 1 8910
0 8912 7 1 2 49612 57938
0 8913 7 1 2 54543 8912
0 8914 5 1 1 8913
0 8915 7 1 2 8911 8914
0 8916 5 1 1 8915
0 8917 7 1 2 44746 8916
0 8918 5 1 1 8917
0 8919 7 1 2 49075 61996
0 8920 5 1 1 8919
0 8921 7 1 2 43029 57180
0 8922 5 2 1 8921
0 8923 7 1 2 48568 55157
0 8924 5 1 1 8923
0 8925 7 1 2 49031 8924
0 8926 7 1 2 62058 8925
0 8927 7 1 2 62157 8926
0 8928 5 1 1 8927
0 8929 7 1 2 8920 8928
0 8930 5 1 1 8929
0 8931 7 7 2 47224 48789
0 8932 5 1 1 62159
0 8933 7 1 2 49613 62160
0 8934 5 1 1 8933
0 8935 7 1 2 57172 8934
0 8936 5 1 1 8935
0 8937 7 1 2 42733 8936
0 8938 5 1 1 8937
0 8939 7 1 2 62063 8938
0 8940 7 1 2 8930 8939
0 8941 5 1 1 8940
0 8942 7 1 2 53246 8941
0 8943 5 1 1 8942
0 8944 7 3 2 47397 54933
0 8945 5 1 1 62166
0 8946 7 1 2 49104 55148
0 8947 7 1 2 62167 8946
0 8948 5 1 1 8947
0 8949 7 3 2 52504 54382
0 8950 7 1 2 52404 52954
0 8951 7 1 2 62169 8950
0 8952 5 1 1 8951
0 8953 7 1 2 8948 8952
0 8954 7 1 2 8943 8953
0 8955 5 1 1 8954
0 8956 7 1 2 60357 8955
0 8957 5 1 1 8956
0 8958 7 1 2 8918 8957
0 8959 5 1 1 8958
0 8960 7 1 2 43254 8959
0 8961 5 1 1 8960
0 8962 7 3 2 53875 60946
0 8963 5 1 1 62172
0 8964 7 2 2 2982 62173
0 8965 5 4 1 62175
0 8966 7 1 2 47225 62177
0 8967 5 1 1 8966
0 8968 7 1 2 48569 61523
0 8969 5 1 1 8968
0 8970 7 1 2 8967 8969
0 8971 5 1 1 8970
0 8972 7 1 2 42501 8971
0 8973 5 1 1 8972
0 8974 7 1 2 53212 8973
0 8975 5 1 1 8974
0 8976 7 1 2 42734 62003
0 8977 5 1 1 8976
0 8978 7 1 2 43864 57547
0 8979 5 1 1 8978
0 8980 7 1 2 51170 8979
0 8981 7 1 2 8977 8980
0 8982 5 1 1 8981
0 8983 7 1 2 52313 60358
0 8984 7 1 2 8982 8983
0 8985 7 1 2 8975 8984
0 8986 5 1 1 8985
0 8987 7 1 2 8961 8986
0 8988 5 1 1 8987
0 8989 7 1 2 55607 8988
0 8990 5 1 1 8989
0 8991 7 1 2 42735 49924
0 8992 5 5 1 8991
0 8993 7 2 2 49682 62181
0 8994 7 1 2 43865 62186
0 8995 5 1 1 8994
0 8996 7 1 2 56312 4956
0 8997 5 1 1 8996
0 8998 7 1 2 43030 8997
0 8999 5 1 1 8998
0 9000 7 1 2 49744 56776
0 9001 5 1 1 9000
0 9002 7 1 2 55693 9001
0 9003 7 1 2 8999 9002
0 9004 5 1 1 9003
0 9005 7 1 2 42736 9004
0 9006 5 1 1 9005
0 9007 7 1 2 8995 9006
0 9008 5 1 1 9007
0 9009 7 1 2 53247 9008
0 9010 5 1 1 9009
0 9011 7 1 2 58454 58150
0 9012 5 1 1 9011
0 9013 7 1 2 9010 9012
0 9014 5 1 1 9013
0 9015 7 1 2 60359 9014
0 9016 5 1 1 9015
0 9017 7 4 2 52744 61392
0 9018 7 2 2 50184 50916
0 9019 7 1 2 62188 62192
0 9020 5 1 1 9019
0 9021 7 1 2 9016 9020
0 9022 5 1 1 9021
0 9023 7 1 2 55608 9022
0 9024 5 1 1 9023
0 9025 7 1 2 49683 50508
0 9026 7 1 2 55895 58303
0 9027 7 1 2 9025 9026
0 9028 7 1 2 54539 9027
0 9029 5 1 1 9028
0 9030 7 1 2 9024 9029
0 9031 5 1 1 9030
0 9032 7 1 2 49202 9031
0 9033 5 1 1 9032
0 9034 7 11 2 43255 47226
0 9035 5 4 1 62194
0 9036 7 1 2 56791 62205
0 9037 5 2 1 9036
0 9038 7 1 2 60975 62209
0 9039 5 1 1 9038
0 9040 7 1 2 47227 61399
0 9041 5 1 1 9040
0 9042 7 1 2 9039 9041
0 9043 5 1 1 9042
0 9044 7 1 2 55609 9043
0 9045 5 1 1 9044
0 9046 7 1 2 54415 57906
0 9047 7 1 2 61805 9046
0 9048 5 1 1 9047
0 9049 7 1 2 9045 9048
0 9050 5 1 1 9049
0 9051 7 1 2 45204 9050
0 9052 5 1 1 9051
0 9053 7 2 2 54416 58393
0 9054 7 4 2 44428 61130
0 9055 7 1 2 49153 62213
0 9056 7 1 2 62211 9055
0 9057 5 2 1 9056
0 9058 7 1 2 9052 62217
0 9059 5 1 1 9058
0 9060 7 1 2 46186 9059
0 9061 5 1 1 9060
0 9062 7 3 2 45205 61428
0 9063 7 2 2 57854 62219
0 9064 7 1 2 55036 55896
0 9065 7 1 2 62222 9064
0 9066 5 1 1 9065
0 9067 7 1 2 9061 9066
0 9068 5 1 1 9067
0 9069 7 1 2 50987 9068
0 9070 5 1 1 9069
0 9071 7 2 2 55548 57168
0 9072 5 3 1 62224
0 9073 7 1 2 61368 62226
0 9074 5 1 1 9073
0 9075 7 2 2 44633 56015
0 9076 7 1 2 51370 62229
0 9077 5 1 1 9076
0 9078 7 1 2 9074 9077
0 9079 5 1 1 9078
0 9080 7 6 2 47744 56867
0 9081 7 1 2 9079 62231
0 9082 5 1 1 9081
0 9083 7 1 2 62218 9082
0 9084 5 1 1 9083
0 9085 7 1 2 62002 9084
0 9086 5 1 1 9085
0 9087 7 1 2 9070 9086
0 9088 7 1 2 9033 9087
0 9089 7 1 2 8990 9088
0 9090 7 1 2 8907 9089
0 9091 5 1 1 9090
0 9092 7 1 2 59358 9091
0 9093 5 1 1 9092
0 9094 7 1 2 8775 9093
0 9095 5 1 1 9094
0 9096 7 1 2 51856 9095
0 9097 5 1 1 9096
0 9098 7 1 2 61369 62103
0 9099 5 1 1 9098
0 9100 7 1 2 52092 60360
0 9101 7 1 2 54172 9100
0 9102 5 1 1 9101
0 9103 7 1 2 9099 9102
0 9104 5 1 1 9103
0 9105 7 1 2 49958 9104
0 9106 5 1 1 9105
0 9107 7 2 2 45422 57677
0 9108 5 1 1 62237
0 9109 7 1 2 61370 62238
0 9110 5 1 1 9109
0 9111 7 5 2 48570 53248
0 9112 5 1 1 62239
0 9113 7 3 2 53523 61701
0 9114 7 1 2 62240 62244
0 9115 5 1 1 9114
0 9116 7 1 2 9110 9115
0 9117 7 1 2 9106 9116
0 9118 5 1 1 9117
0 9119 7 1 2 58154 9118
0 9120 5 1 1 9119
0 9121 7 1 2 57837 60976
0 9122 5 1 1 9121
0 9123 7 1 2 50923 61719
0 9124 5 1 1 9123
0 9125 7 1 2 9122 9124
0 9126 5 1 1 9125
0 9127 7 1 2 56309 9126
0 9128 5 1 1 9127
0 9129 7 2 2 50917 53996
0 9130 7 1 2 62071 62247
0 9131 5 1 1 9130
0 9132 7 1 2 9128 9131
0 9133 5 1 1 9132
0 9134 7 1 2 47522 9133
0 9135 5 1 1 9134
0 9136 7 2 2 43031 56708
0 9137 5 1 1 62249
0 9138 7 2 2 49884 9137
0 9139 5 2 1 62251
0 9140 7 2 2 45206 62253
0 9141 7 3 2 51548 55171
0 9142 7 1 2 62255 62257
0 9143 5 1 1 9142
0 9144 7 1 2 9135 9143
0 9145 5 1 1 9144
0 9146 7 1 2 45423 9145
0 9147 5 1 1 9146
0 9148 7 1 2 44185 51499
0 9149 5 1 1 9148
0 9150 7 1 2 58808 9149
0 9151 5 1 1 9150
0 9152 7 1 2 52745 60977
0 9153 7 1 2 9151 9152
0 9154 5 1 1 9153
0 9155 7 1 2 9147 9154
0 9156 5 1 1 9155
0 9157 7 1 2 46638 9156
0 9158 5 1 1 9157
0 9159 7 3 2 49684 60361
0 9160 7 2 2 56511 62260
0 9161 7 1 2 47086 62263
0 9162 5 1 1 9161
0 9163 7 1 2 49685 62008
0 9164 5 1 1 9163
0 9165 7 1 2 45207 62189
0 9166 5 1 1 9165
0 9167 7 1 2 9164 9166
0 9168 5 1 1 9167
0 9169 7 1 2 45992 9168
0 9170 5 1 1 9169
0 9171 7 1 2 9162 9170
0 9172 5 2 1 9171
0 9173 7 1 2 59099 62265
0 9174 5 1 1 9173
0 9175 7 3 2 46448 49076
0 9176 5 9 1 62267
0 9177 7 5 2 60708 62270
0 9178 5 1 1 62279
0 9179 7 1 2 47398 9178
0 9180 5 1 1 9179
0 9181 7 2 2 45208 60362
0 9182 7 2 2 44030 49203
0 9183 5 6 1 62286
0 9184 7 1 2 51364 58492
0 9185 7 1 2 62288 9184
0 9186 7 1 2 62284 9185
0 9187 7 1 2 9180 9186
0 9188 5 1 1 9187
0 9189 7 1 2 9174 9188
0 9190 7 1 2 9158 9189
0 9191 5 1 1 9190
0 9192 7 1 2 58863 9191
0 9193 5 1 1 9192
0 9194 7 1 2 9120 9193
0 9195 5 1 1 9194
0 9196 7 1 2 46187 9195
0 9197 5 1 1 9196
0 9198 7 1 2 45209 59059
0 9199 5 1 1 9198
0 9200 7 1 2 42502 62143
0 9201 5 1 1 9200
0 9202 7 1 2 9199 9201
0 9203 5 1 1 9202
0 9204 7 1 2 60363 9203
0 9205 5 1 1 9204
0 9206 7 2 2 47962 54093
0 9207 7 1 2 45993 52398
0 9208 7 1 2 57977 9207
0 9209 7 1 2 62294 9208
0 9210 5 1 1 9209
0 9211 7 1 2 9205 9210
0 9212 5 1 1 9211
0 9213 7 1 2 49959 9212
0 9214 5 1 1 9213
0 9215 7 2 2 46188 61371
0 9216 7 1 2 57058 62296
0 9217 5 1 1 9216
0 9218 7 1 2 9214 9217
0 9219 5 1 1 9218
0 9220 7 1 2 50988 9219
0 9221 5 1 1 9220
0 9222 7 4 2 58612 60737
0 9223 5 3 1 62298
0 9224 7 2 2 58383 62302
0 9225 5 4 1 62305
0 9226 7 1 2 54149 58152
0 9227 5 2 1 9226
0 9228 7 1 2 42503 62311
0 9229 5 1 1 9228
0 9230 7 1 2 54170 9229
0 9231 5 1 1 9230
0 9232 7 1 2 60364 9231
0 9233 5 1 1 9232
0 9234 7 2 2 50545 61393
0 9235 7 1 2 55037 62313
0 9236 5 1 1 9235
0 9237 7 1 2 9233 9236
0 9238 5 1 1 9237
0 9239 7 1 2 62307 9238
0 9240 5 1 1 9239
0 9241 7 1 2 58601 61964
0 9242 5 1 1 9241
0 9243 7 1 2 49960 9242
0 9244 5 1 1 9243
0 9245 7 2 2 49686 55230
0 9246 5 2 1 62315
0 9247 7 1 2 9244 62317
0 9248 7 1 2 4909 9247
0 9249 5 1 1 9248
0 9250 7 4 2 53249 60365
0 9251 5 1 1 62319
0 9252 7 1 2 42737 62320
0 9253 7 1 2 9249 9252
0 9254 5 1 1 9253
0 9255 7 2 2 9240 9254
0 9256 5 1 1 62323
0 9257 7 1 2 9221 62324
0 9258 5 1 1 9257
0 9259 7 1 2 58155 9258
0 9260 5 1 1 9259
0 9261 7 2 2 47963 51050
0 9262 7 4 2 45994 56818
0 9263 5 1 1 62327
0 9264 7 5 2 46639 49273
0 9265 7 5 2 47523 62331
0 9266 7 2 2 62328 62336
0 9267 7 2 2 62325 62341
0 9268 5 1 1 62343
0 9269 7 1 2 45424 62344
0 9270 5 1 1 9269
0 9271 7 4 2 46449 56702
0 9272 5 2 1 62345
0 9273 7 1 2 48571 57659
0 9274 7 1 2 62349 9273
0 9275 7 1 2 62252 9274
0 9276 5 3 1 9275
0 9277 7 1 2 45425 62256
0 9278 5 1 1 9277
0 9279 7 1 2 62351 9278
0 9280 5 1 1 9279
0 9281 7 1 2 43866 9280
0 9282 5 1 1 9281
0 9283 7 1 2 1045 9282
0 9284 5 1 1 9283
0 9285 7 1 2 46640 9284
0 9286 5 1 1 9285
0 9287 7 1 2 257 53497
0 9288 5 3 1 9287
0 9289 7 4 2 48790 62354
0 9290 5 1 1 62357
0 9291 7 1 2 43032 59074
0 9292 5 1 1 9291
0 9293 7 1 2 9290 9292
0 9294 5 1 1 9293
0 9295 7 1 2 57181 9294
0 9296 5 1 1 9295
0 9297 7 8 2 43256 44031
0 9298 5 2 1 62361
0 9299 7 2 2 57051 62362
0 9300 7 1 2 52181 62371
0 9301 5 2 1 9300
0 9302 7 1 2 9296 62373
0 9303 7 1 2 9286 9302
0 9304 5 1 1 9303
0 9305 7 1 2 62321 9304
0 9306 5 1 1 9305
0 9307 7 1 2 9270 9306
0 9308 5 1 1 9307
0 9309 7 1 2 42738 58864
0 9310 7 1 2 9308 9309
0 9311 5 1 1 9310
0 9312 7 1 2 9260 9311
0 9313 7 1 2 9197 9312
0 9314 5 1 1 9313
0 9315 7 1 2 47626 9314
0 9316 5 1 1 9315
0 9317 7 3 2 47524 52845
0 9318 5 1 1 62375
0 9319 7 2 2 44186 53739
0 9320 5 1 1 62378
0 9321 7 1 2 9318 9320
0 9322 5 1 1 9321
0 9323 7 1 2 46641 9322
0 9324 5 1 1 9323
0 9325 7 1 2 52810 61069
0 9326 5 1 1 9325
0 9327 7 1 2 46450 9326
0 9328 5 1 1 9327
0 9329 7 1 2 9324 9328
0 9330 5 1 1 9329
0 9331 7 1 2 62190 9330
0 9332 5 1 1 9331
0 9333 7 2 2 49614 57245
0 9334 5 1 1 62380
0 9335 7 1 2 57741 62381
0 9336 5 2 1 9335
0 9337 7 1 2 43033 56747
0 9338 5 2 1 9337
0 9339 7 1 2 58538 62384
0 9340 5 3 1 9339
0 9341 7 1 2 56651 62386
0 9342 5 1 1 9341
0 9343 7 2 2 50152 56886
0 9344 5 2 1 62389
0 9345 7 1 2 9342 62391
0 9346 5 2 1 9345
0 9347 7 1 2 42739 62393
0 9348 5 1 1 9347
0 9349 7 6 2 48791 50989
0 9350 5 1 1 62395
0 9351 7 5 2 50833 62396
0 9352 5 1 1 62401
0 9353 7 1 2 49334 62402
0 9354 5 1 1 9353
0 9355 7 1 2 42740 56652
0 9356 5 2 1 9355
0 9357 7 1 2 49790 60200
0 9358 5 1 1 9357
0 9359 7 2 2 62406 9358
0 9360 7 1 2 43867 52911
0 9361 7 1 2 62408 9360
0 9362 7 1 2 9354 9361
0 9363 5 1 1 9362
0 9364 7 5 2 44032 49615
0 9365 5 3 1 62410
0 9366 7 3 2 42741 48792
0 9367 5 2 1 62418
0 9368 7 1 2 62415 62421
0 9369 5 1 1 9368
0 9370 7 1 2 43034 9369
0 9371 5 1 1 9370
0 9372 7 2 2 45426 49626
0 9373 5 1 1 62423
0 9374 7 3 2 49635 9373
0 9375 7 1 2 42742 62425
0 9376 5 1 1 9375
0 9377 7 1 2 9371 9376
0 9378 5 1 1 9377
0 9379 7 1 2 43257 9378
0 9380 5 1 1 9379
0 9381 7 1 2 47228 7440
0 9382 7 1 2 9380 9381
0 9383 5 1 1 9382
0 9384 7 1 2 9363 9383
0 9385 5 1 1 9384
0 9386 7 1 2 9348 9385
0 9387 5 1 1 9386
0 9388 7 1 2 43710 9387
0 9389 5 1 1 9388
0 9390 7 1 2 62382 9389
0 9391 5 1 1 9390
0 9392 7 1 2 60366 9391
0 9393 5 1 1 9392
0 9394 7 1 2 9332 9393
0 9395 5 1 1 9394
0 9396 7 1 2 45995 9395
0 9397 5 1 1 9396
0 9398 7 1 2 44747 53474
0 9399 7 2 2 62287 9398
0 9400 7 1 2 43035 51201
0 9401 7 2 2 62428 9400
0 9402 7 1 2 54531 62430
0 9403 5 1 1 9402
0 9404 7 1 2 43258 62426
0 9405 5 1 1 9404
0 9406 7 1 2 58466 9405
0 9407 5 3 1 9406
0 9408 7 1 2 53997 62432
0 9409 5 2 1 9408
0 9410 7 2 2 43711 56653
0 9411 7 1 2 52746 62437
0 9412 5 1 1 9411
0 9413 7 1 2 62435 9412
0 9414 5 1 1 9413
0 9415 7 1 2 46451 9414
0 9416 5 1 1 9415
0 9417 7 1 2 47229 62433
0 9418 5 1 1 9417
0 9419 7 3 2 50834 62161
0 9420 5 3 1 62439
0 9421 7 2 2 53457 60202
0 9422 7 1 2 62442 62445
0 9423 5 1 1 9422
0 9424 7 1 2 43036 9423
0 9425 5 1 1 9424
0 9426 7 1 2 50753 53485
0 9427 5 1 1 9426
0 9428 7 1 2 47230 60814
0 9429 5 1 1 9428
0 9430 7 2 2 45210 9429
0 9431 5 1 1 62447
0 9432 7 1 2 9427 9431
0 9433 7 1 2 9425 9432
0 9434 7 1 2 9418 9433
0 9435 5 1 1 9434
0 9436 7 1 2 42743 9435
0 9437 5 1 1 9436
0 9438 7 1 2 50835 57150
0 9439 5 2 1 9438
0 9440 7 1 2 62446 62449
0 9441 5 1 1 9440
0 9442 7 1 2 43868 9441
0 9443 5 1 1 9442
0 9444 7 1 2 52245 52933
0 9445 5 1 1 9444
0 9446 7 1 2 9443 9445
0 9447 5 1 1 9446
0 9448 7 1 2 43037 9447
0 9449 5 1 1 9448
0 9450 7 3 2 46642 52955
0 9451 7 1 2 57088 62451
0 9452 5 1 1 9451
0 9453 7 1 2 9449 9452
0 9454 7 1 2 9437 9453
0 9455 5 1 1 9454
0 9456 7 1 2 47087 9455
0 9457 5 1 1 9456
0 9458 7 1 2 9416 9457
0 9459 5 1 1 9458
0 9460 7 1 2 48087 9459
0 9461 5 1 1 9460
0 9462 7 1 2 9403 9461
0 9463 5 1 1 9462
0 9464 7 1 2 62022 9463
0 9465 5 1 1 9464
0 9466 7 2 2 9397 9465
0 9467 5 1 1 62454
0 9468 7 1 2 54173 62434
0 9469 5 1 1 9468
0 9470 7 2 2 43712 52236
0 9471 7 4 2 42504 56654
0 9472 5 1 1 62458
0 9473 7 1 2 62456 62459
0 9474 5 1 1 9473
0 9475 7 1 2 9469 9474
0 9476 5 1 1 9475
0 9477 7 1 2 60367 9476
0 9478 5 1 1 9477
0 9479 7 2 2 48572 60746
0 9480 5 3 1 62462
0 9481 7 1 2 44187 62464
0 9482 5 1 1 9481
0 9483 7 1 2 61070 9482
0 9484 5 1 1 9483
0 9485 7 1 2 52237 61185
0 9486 7 1 2 9484 9485
0 9487 5 1 1 9486
0 9488 7 1 2 9478 9487
0 9489 5 1 1 9488
0 9490 7 1 2 46189 9489
0 9491 5 1 1 9490
0 9492 7 1 2 55568 61444
0 9493 5 1 1 9492
0 9494 7 6 2 47525 44634
0 9495 7 1 2 48088 62467
0 9496 7 1 2 60141 9495
0 9497 5 1 1 9496
0 9498 7 1 2 9493 9497
0 9499 5 1 1 9498
0 9500 7 1 2 54119 9499
0 9501 5 1 1 9500
0 9502 7 2 2 46190 56800
0 9503 7 1 2 61186 62473
0 9504 5 1 1 9503
0 9505 7 1 2 9501 9504
0 9506 5 1 1 9505
0 9507 7 1 2 50990 9506
0 9508 5 1 1 9507
0 9509 7 1 2 9491 9508
0 9510 7 1 2 62455 9509
0 9511 5 1 1 9510
0 9512 7 1 2 60932 9511
0 9513 5 1 1 9512
0 9514 7 1 2 9316 9513
0 9515 5 1 1 9514
0 9516 7 1 2 60564 9515
0 9517 5 1 1 9516
0 9518 7 6 2 44429 56176
0 9519 7 1 2 59060 60368
0 9520 5 1 1 9519
0 9521 7 1 2 55053 61131
0 9522 5 1 1 9521
0 9523 7 1 2 9520 9522
0 9524 5 1 1 9523
0 9525 7 1 2 62475 9524
0 9526 5 1 1 9525
0 9527 7 69 2 41994 44430
0 9528 5 3 1 62481
0 9529 7 1 2 61372 62482
0 9530 5 1 1 9529
0 9531 7 2 2 56016 58937
0 9532 7 1 2 60032 62553
0 9533 5 1 1 9532
0 9534 7 1 2 9530 9533
0 9535 5 1 1 9534
0 9536 7 1 2 49274 60276
0 9537 7 1 2 9535 9536
0 9538 5 1 1 9537
0 9539 7 1 2 9526 9538
0 9540 5 1 1 9539
0 9541 7 1 2 46825 9540
0 9542 5 1 1 9541
0 9543 7 1 2 45544 62214
0 9544 7 2 2 46191 55857
0 9545 7 1 2 62329 62555
0 9546 7 1 2 9543 9545
0 9547 5 1 1 9546
0 9548 7 1 2 9542 9547
0 9549 5 1 1 9548
0 9550 7 1 2 47627 9549
0 9551 5 1 1 9550
0 9552 7 2 2 60369 60633
0 9553 7 1 2 61554 62557
0 9554 7 1 2 56111 9553
0 9555 5 1 1 9554
0 9556 7 1 2 9551 9555
0 9557 5 1 1 9556
0 9558 7 1 2 45211 9557
0 9559 5 1 1 9558
0 9560 7 2 2 55181 59145
0 9561 7 4 2 48573 61132
0 9562 7 1 2 57033 62561
0 9563 7 1 2 62559 9562
0 9564 5 1 1 9563
0 9565 7 1 2 51137 55438
0 9566 7 1 2 54126 9565
0 9567 7 1 2 62558 9566
0 9568 5 1 1 9567
0 9569 7 1 2 9564 9568
0 9570 5 1 1 9569
0 9571 7 1 2 46452 9570
0 9572 5 1 1 9571
0 9573 7 1 2 61895 62322
0 9574 7 1 2 52109 9573
0 9575 5 1 1 9574
0 9576 7 1 2 9572 9575
0 9577 5 1 1 9576
0 9578 7 1 2 41995 9577
0 9579 5 1 1 9578
0 9580 7 1 2 48574 52033
0 9581 7 1 2 58254 9580
0 9582 7 1 2 61477 61628
0 9583 7 1 2 9581 9582
0 9584 5 1 1 9583
0 9585 7 1 2 9579 9584
0 9586 7 1 2 9559 9585
0 9587 5 1 1 9586
0 9588 7 1 2 60565 9587
0 9589 5 1 1 9588
0 9590 7 1 2 52112 61365
0 9591 5 1 1 9590
0 9592 7 1 2 52113 9251
0 9593 5 1 1 9592
0 9594 7 1 2 61772 9593
0 9595 7 1 2 9591 9594
0 9596 5 1 1 9595
0 9597 7 1 2 9589 9596
0 9598 5 1 1 9597
0 9599 7 1 2 50059 9598
0 9600 5 1 1 9599
0 9601 7 1 2 56949 60668
0 9602 5 1 1 9601
0 9603 7 1 2 60779 9602
0 9604 5 6 1 9603
0 9605 7 1 2 57126 62206
0 9606 5 1 1 9605
0 9607 7 1 2 50991 9606
0 9608 5 1 1 9607
0 9609 7 1 2 47231 56899
0 9610 5 1 1 9609
0 9611 7 1 2 50279 57097
0 9612 5 2 1 9611
0 9613 7 1 2 52238 62571
0 9614 5 1 1 9613
0 9615 7 1 2 9610 9614
0 9616 7 1 2 9608 9615
0 9617 5 1 1 9616
0 9618 7 1 2 46192 9617
0 9619 5 1 1 9618
0 9620 7 2 2 46643 54957
0 9621 5 1 1 62573
0 9622 7 1 2 51351 55539
0 9623 7 3 2 9621 9622
0 9624 7 1 2 54114 62575
0 9625 5 1 1 9624
0 9626 7 1 2 9619 9625
0 9627 5 3 1 9626
0 9628 7 1 2 61641 61512
0 9629 7 1 2 62578 9628
0 9630 5 1 1 9629
0 9631 7 1 2 52893 62009
0 9632 5 1 1 9631
0 9633 7 1 2 58564 62191
0 9634 5 1 1 9633
0 9635 7 1 2 9632 9634
0 9636 5 1 1 9635
0 9637 7 1 2 42744 9636
0 9638 5 1 1 9637
0 9639 7 3 2 46193 53088
0 9640 5 1 1 62581
0 9641 7 1 2 62582 62314
0 9642 5 1 1 9641
0 9643 7 1 2 9638 9642
0 9644 5 1 1 9643
0 9645 7 10 2 45545 59146
0 9646 7 2 2 50060 62584
0 9647 7 1 2 9644 62594
0 9648 5 1 1 9647
0 9649 7 1 2 9630 9648
0 9650 5 1 1 9649
0 9651 7 1 2 45996 9650
0 9652 5 1 1 9651
0 9653 7 1 2 52894 55080
0 9654 5 1 1 9653
0 9655 7 2 2 45212 60277
0 9656 7 4 2 47399 51099
0 9657 7 1 2 62596 62598
0 9658 5 1 1 9657
0 9659 7 1 2 9654 9658
0 9660 5 1 1 9659
0 9661 7 2 2 59147 59988
0 9662 7 1 2 61791 62602
0 9663 7 1 2 9660 9662
0 9664 5 1 1 9663
0 9665 7 1 2 9652 9664
0 9666 5 2 1 9665
0 9667 7 1 2 62565 62604
0 9668 5 1 1 9667
0 9669 7 1 2 48575 61889
0 9670 5 1 1 9669
0 9671 7 1 2 8361 9670
0 9672 5 3 1 9671
0 9673 7 2 2 59061 61792
0 9674 7 1 2 61815 62609
0 9675 5 1 1 9674
0 9676 7 2 2 57012 61032
0 9677 7 2 2 47232 56887
0 9678 7 1 2 61672 62613
0 9679 7 1 2 62611 9678
0 9680 5 1 1 9679
0 9681 7 1 2 9675 9680
0 9682 5 1 1 9681
0 9683 7 1 2 62606 9682
0 9684 5 1 1 9683
0 9685 7 1 2 9668 9684
0 9686 7 1 2 9600 9685
0 9687 7 1 2 9517 9686
0 9688 7 1 2 9097 9687
0 9689 5 1 1 9688
0 9690 7 1 2 48405 9689
0 9691 5 1 1 9690
0 9692 7 2 2 48576 61373
0 9693 7 2 2 49032 62615
0 9694 7 1 2 62094 62617
0 9695 5 1 1 9694
0 9696 7 5 2 45213 53250
0 9697 7 2 2 42745 49077
0 9698 5 1 1 62624
0 9699 7 1 2 62245 62625
0 9700 7 1 2 62619 9699
0 9701 5 1 1 9700
0 9702 7 1 2 9695 9701
0 9703 5 1 1 9702
0 9704 7 1 2 43259 9703
0 9705 5 1 1 9704
0 9706 7 1 2 46644 56765
0 9707 7 1 2 62083 62246
0 9708 7 1 2 9706 9707
0 9709 5 1 1 9708
0 9710 7 1 2 9705 9709
0 9711 5 1 1 9710
0 9712 7 1 2 61223 9711
0 9713 5 1 1 9712
0 9714 7 2 2 53524 60370
0 9715 7 1 2 59177 59422
0 9716 7 1 2 62626 9715
0 9717 7 1 2 62084 9716
0 9718 7 1 2 57073 9717
0 9719 5 1 1 9718
0 9720 7 1 2 9713 9719
0 9721 5 1 1 9720
0 9722 7 1 2 54760 9721
0 9723 5 1 1 9722
0 9724 7 5 2 51967 60371
0 9725 7 1 2 50061 61490
0 9726 5 1 1 9725
0 9727 7 1 2 50754 58718
0 9728 5 1 1 9727
0 9729 7 1 2 9726 9728
0 9730 5 1 1 9729
0 9731 7 2 2 53251 9730
0 9732 7 1 2 44033 62633
0 9733 5 1 1 9732
0 9734 7 1 2 49961 61046
0 9735 5 1 1 9734
0 9736 7 1 2 51209 58719
0 9737 5 1 1 9736
0 9738 7 1 2 9735 9737
0 9739 5 1 1 9738
0 9740 7 1 2 62620 9739
0 9741 5 1 1 9740
0 9742 7 1 2 9733 9741
0 9743 5 1 1 9742
0 9744 7 1 2 43038 9743
0 9745 5 1 1 9744
0 9746 7 1 2 60808 61621
0 9747 7 1 2 62621 9746
0 9748 5 1 1 9747
0 9749 7 1 2 9745 9748
0 9750 5 1 1 9749
0 9751 7 1 2 62628 9750
0 9752 5 1 1 9751
0 9753 7 1 2 58689 60978
0 9754 5 1 1 9753
0 9755 7 1 2 61047 61374
0 9756 5 1 1 9755
0 9757 7 1 2 9754 9756
0 9758 5 1 1 9757
0 9759 7 1 2 50992 9758
0 9760 5 1 1 9759
0 9761 7 4 2 47088 56075
0 9762 7 2 2 58289 61429
0 9763 7 1 2 44431 62639
0 9764 7 1 2 62635 9763
0 9765 5 1 1 9764
0 9766 7 1 2 9760 9765
0 9767 5 1 1 9766
0 9768 7 1 2 47233 9767
0 9769 5 1 1 9768
0 9770 7 1 2 56423 61133
0 9771 7 1 2 61694 9770
0 9772 7 1 2 62636 9771
0 9773 5 1 1 9772
0 9774 7 1 2 9769 9773
0 9775 5 1 1 9774
0 9776 7 1 2 49962 9775
0 9777 5 1 1 9776
0 9778 7 2 2 57630 60372
0 9779 7 5 2 42505 54934
0 9780 5 1 1 62643
0 9781 7 1 2 45700 62644
0 9782 7 1 2 62641 9781
0 9783 7 1 2 62403 9782
0 9784 5 1 1 9783
0 9785 7 1 2 9777 9784
0 9786 5 1 1 9785
0 9787 7 1 2 46194 9786
0 9788 5 1 1 9787
0 9789 7 5 2 48089 56085
0 9790 7 1 2 54013 62648
0 9791 7 1 2 62634 9790
0 9792 5 1 1 9791
0 9793 7 8 2 42150 46453
0 9794 7 1 2 45997 62653
0 9795 7 1 2 62640 9794
0 9796 7 2 2 43260 56819
0 9797 7 2 2 47400 58918
0 9798 7 1 2 62661 62663
0 9799 7 1 2 9795 9798
0 9800 5 1 1 9799
0 9801 7 1 2 9792 9800
0 9802 7 1 2 9788 9801
0 9803 5 1 1 9802
0 9804 7 1 2 48577 9803
0 9805 5 1 1 9804
0 9806 7 1 2 9752 9805
0 9807 5 1 1 9806
0 9808 7 1 2 59836 9807
0 9809 5 1 1 9808
0 9810 7 1 2 9723 9809
0 9811 7 1 2 9691 9810
0 9812 7 1 2 8354 9811
0 9813 5 1 1 9812
0 9814 7 6 2 46906 43569
0 9815 7 2 2 42254 62665
0 9816 5 1 1 62671
0 9817 7 8 2 43524 46951
0 9818 7 1 2 45783 62673
0 9819 5 1 1 9818
0 9820 7 1 2 9816 9819
0 9821 5 14 1 9820
0 9822 7 1 2 9813 62681
0 9823 5 1 1 9822
0 9824 7 5 2 42255 44309
0 9825 7 17 2 43525 43570
0 9826 5 1 1 62700
0 9827 7 6 2 43448 62701
0 9828 7 19 2 62695 62717
0 9829 5 7 1 62723
0 9830 7 9 2 45701 56950
0 9831 5 2 1 62749
0 9832 7 2 2 47526 62750
0 9833 5 1 1 62760
0 9834 7 5 2 46454 44555
0 9835 7 1 2 42151 62762
0 9836 5 1 1 9835
0 9837 7 1 2 9833 9836
0 9838 5 1 1 9837
0 9839 7 1 2 56633 9838
0 9840 5 1 1 9839
0 9841 7 2 2 45702 55731
0 9842 5 3 1 62767
0 9843 7 2 2 49154 59249
0 9844 5 1 1 62772
0 9845 7 1 2 62769 9844
0 9846 5 1 1 9845
0 9847 7 1 2 42506 9846
0 9848 5 1 1 9847
0 9849 7 3 2 49204 59250
0 9850 5 1 1 62774
0 9851 7 4 2 45703 57768
0 9852 7 2 2 48793 62777
0 9853 5 2 1 62781
0 9854 7 1 2 9850 62783
0 9855 5 2 1 9854
0 9856 7 2 2 43039 62785
0 9857 5 2 1 62787
0 9858 7 1 2 696 59321
0 9859 5 4 1 9858
0 9860 7 1 2 42507 62791
0 9861 5 1 1 9860
0 9862 7 1 2 62789 9861
0 9863 5 1 1 9862
0 9864 7 1 2 47401 9863
0 9865 5 1 1 9864
0 9866 7 1 2 9848 9865
0 9867 5 1 1 9866
0 9868 7 1 2 52034 9867
0 9869 5 1 1 9868
0 9870 7 1 2 9840 9869
0 9871 5 1 1 9870
0 9872 7 1 2 47089 9871
0 9873 5 1 1 9872
0 9874 7 1 2 59251 62289
0 9875 5 1 1 9874
0 9876 7 1 2 50993 51896
0 9877 5 1 1 9876
0 9878 7 1 2 9875 9877
0 9879 5 1 1 9878
0 9880 7 1 2 55038 55099
0 9881 7 1 2 9879 9880
0 9882 5 1 1 9881
0 9883 7 1 2 9873 9882
0 9884 5 1 1 9883
0 9885 7 1 2 61134 9884
0 9886 5 1 1 9885
0 9887 7 7 2 48794 61135
0 9888 7 2 2 57769 61630
0 9889 7 2 2 46455 56820
0 9890 7 1 2 62802 62804
0 9891 7 1 2 62795 9890
0 9892 5 1 1 9891
0 9893 7 3 2 48090 58009
0 9894 7 1 2 42152 58019
0 9895 7 1 2 61711 9894
0 9896 7 1 2 62806 9895
0 9897 5 1 1 9896
0 9898 7 1 2 9892 9897
0 9899 5 1 1 9898
0 9900 7 1 2 44034 9899
0 9901 5 1 1 9900
0 9902 7 1 2 50452 55004
0 9903 7 1 2 62627 9902
0 9904 7 1 2 62786 9903
0 9905 5 1 1 9904
0 9906 7 1 2 9901 9905
0 9907 7 1 2 9886 9906
0 9908 5 1 1 9907
0 9909 7 1 2 46645 9908
0 9910 5 1 1 9909
0 9911 7 5 2 44188 51171
0 9912 7 1 2 51814 56951
0 9913 5 1 1 9912
0 9914 7 7 2 42153 57781
0 9915 5 2 1 62814
0 9916 7 1 2 46456 62815
0 9917 5 1 1 9916
0 9918 7 1 2 9913 9917
0 9919 5 1 1 9918
0 9920 7 1 2 62809 9919
0 9921 5 1 1 9920
0 9922 7 1 2 51897 57651
0 9923 5 1 1 9922
0 9924 7 1 2 58681 9923
0 9925 5 4 1 9924
0 9926 7 1 2 52505 62823
0 9927 5 1 1 9926
0 9928 7 1 2 9921 9927
0 9929 5 1 1 9928
0 9930 7 1 2 43261 9929
0 9931 5 1 1 9930
0 9932 7 1 2 298 51898
0 9933 5 1 1 9932
0 9934 7 1 2 58682 9933
0 9935 5 1 1 9934
0 9936 7 1 2 53252 9935
0 9937 5 1 1 9936
0 9938 7 1 2 9931 9937
0 9939 5 1 1 9938
0 9940 7 1 2 52035 9939
0 9941 5 1 1 9940
0 9942 7 1 2 51899 57052
0 9943 5 1 1 9942
0 9944 7 2 2 53356 59252
0 9945 7 1 2 49033 62827
0 9946 5 1 1 9945
0 9947 7 1 2 9943 9946
0 9948 5 1 1 9947
0 9949 7 1 2 50405 9948
0 9950 5 1 1 9949
0 9951 7 1 2 9941 9950
0 9952 5 1 1 9951
0 9953 7 1 2 61136 9952
0 9954 5 1 1 9953
0 9955 7 1 2 50453 62824
0 9956 5 1 1 9955
0 9957 7 1 2 58884 62751
0 9958 5 1 1 9957
0 9959 7 1 2 9956 9958
0 9960 5 1 1 9959
0 9961 7 1 2 43040 9960
0 9962 5 1 1 9961
0 9963 7 2 2 42154 50670
0 9964 7 1 2 49454 62829
0 9965 5 1 1 9964
0 9966 7 1 2 9962 9965
0 9967 5 1 1 9966
0 9968 7 1 2 53160 62649
0 9969 7 1 2 9967 9968
0 9970 5 1 1 9969
0 9971 7 1 2 9954 9970
0 9972 5 1 1 9971
0 9973 7 1 2 47402 9972
0 9974 5 1 1 9973
0 9975 7 8 2 46457 47964
0 9976 5 1 1 62831
0 9977 7 3 2 44748 62832
0 9978 7 1 2 58683 62758
0 9979 5 1 1 9978
0 9980 7 1 2 53998 9979
0 9981 5 1 1 9980
0 9982 7 7 2 47527 47881
0 9983 7 8 2 45704 62842
0 9984 5 1 1 62849
0 9985 7 1 2 55067 62850
0 9986 5 1 1 9985
0 9987 7 1 2 9981 9986
0 9988 5 1 1 9987
0 9989 7 1 2 45998 9988
0 9990 5 1 1 9989
0 9991 7 1 2 55086 62851
0 9992 5 1 1 9991
0 9993 7 1 2 9990 9992
0 9994 5 1 1 9993
0 9995 7 1 2 62839 9994
0 9996 5 1 1 9995
0 9997 7 1 2 9974 9996
0 9998 7 1 2 9910 9997
0 9999 5 1 1 9998
0 10000 7 1 2 45214 9999
0 10001 5 1 1 10000
0 10002 7 4 2 44035 52054
0 10003 7 1 2 51828 62821
0 10004 5 2 1 10003
0 10005 7 1 2 62857 62861
0 10006 5 1 1 10005
0 10007 7 5 2 43869 47882
0 10008 7 6 2 45705 62863
0 10009 7 1 2 42746 62868
0 10010 5 1 1 10009
0 10011 7 1 2 10006 10010
0 10012 5 1 1 10011
0 10013 7 1 2 48578 10012
0 10014 5 1 1 10013
0 10015 7 1 2 51968 62816
0 10016 5 1 1 10015
0 10017 7 1 2 10014 10016
0 10018 5 1 1 10017
0 10019 7 1 2 49963 60373
0 10020 7 1 2 10018 10019
0 10021 5 1 1 10020
0 10022 7 2 2 46646 62773
0 10023 5 1 1 62874
0 10024 7 1 2 62770 10023
0 10025 5 1 1 10024
0 10026 7 1 2 50062 52747
0 10027 7 1 2 61420 10026
0 10028 7 1 2 10025 10027
0 10029 5 1 1 10028
0 10030 7 1 2 10021 10029
0 10031 5 1 1 10030
0 10032 7 1 2 53253 10031
0 10033 5 1 1 10032
0 10034 7 2 2 57865 61631
0 10035 5 1 1 62876
0 10036 7 1 2 48795 62877
0 10037 5 1 1 10036
0 10038 7 1 2 45999 62775
0 10039 5 1 1 10038
0 10040 7 1 2 10037 10039
0 10041 5 1 1 10040
0 10042 7 11 2 47403 48579
0 10043 5 1 1 62878
0 10044 7 2 2 61513 62879
0 10045 7 1 2 10041 62889
0 10046 5 1 1 10045
0 10047 7 2 2 49687 52036
0 10048 5 2 1 62891
0 10049 7 1 2 1490 62893
0 10050 5 1 1 10049
0 10051 7 1 2 46000 10050
0 10052 5 1 1 10051
0 10053 7 1 2 54094 55689
0 10054 5 1 1 10053
0 10055 7 1 2 10052 10054
0 10056 5 1 1 10055
0 10057 7 1 2 61137 10056
0 10058 5 1 1 10057
0 10059 7 1 2 57040 62261
0 10060 5 1 1 10059
0 10061 7 1 2 10058 10060
0 10062 5 1 1 10061
0 10063 7 1 2 49155 62792
0 10064 7 1 2 10062 10063
0 10065 5 1 1 10064
0 10066 7 1 2 10046 10065
0 10067 5 1 1 10066
0 10068 7 1 2 46458 10067
0 10069 5 1 1 10068
0 10070 7 3 2 43041 59253
0 10071 5 1 1 62895
0 10072 7 1 2 62784 10071
0 10073 5 1 1 10072
0 10074 7 1 2 48580 10073
0 10075 5 1 1 10074
0 10076 7 3 2 45706 55419
0 10077 5 1 1 62898
0 10078 7 1 2 49877 62899
0 10079 5 1 1 10078
0 10080 7 1 2 62790 10079
0 10081 7 1 2 10075 10080
0 10082 5 1 1 10081
0 10083 7 1 2 62258 10082
0 10084 5 1 1 10083
0 10085 7 1 2 53964 62852
0 10086 7 1 2 61445 10085
0 10087 5 1 1 10086
0 10088 7 1 2 46647 10087
0 10089 7 1 2 10084 10088
0 10090 7 1 2 10069 10089
0 10091 5 1 1 10090
0 10092 7 1 2 43042 62825
0 10093 5 1 1 10092
0 10094 7 1 2 59637 62853
0 10095 5 1 1 10094
0 10096 7 1 2 10093 10095
0 10097 5 1 1 10096
0 10098 7 1 2 62259 10097
0 10099 5 1 1 10098
0 10100 7 1 2 55236 59254
0 10101 5 1 1 10100
0 10102 7 1 2 48997 51900
0 10103 7 1 2 2508 10102
0 10104 5 1 1 10103
0 10105 7 1 2 10101 10104
0 10106 5 1 1 10105
0 10107 7 1 2 44189 10106
0 10108 5 1 1 10107
0 10109 7 1 2 59255 62880
0 10110 7 1 2 62268 10109
0 10111 5 1 1 10110
0 10112 7 1 2 10108 10111
0 10113 5 1 1 10112
0 10114 7 1 2 61187 10113
0 10115 5 1 1 10114
0 10116 7 1 2 43262 10115
0 10117 7 1 2 10099 10116
0 10118 5 1 1 10117
0 10119 7 1 2 10091 10118
0 10120 5 1 1 10119
0 10121 7 1 2 10033 10120
0 10122 7 1 2 10001 10121
0 10123 5 1 1 10122
0 10124 7 1 2 62724 10123
0 10125 5 1 1 10124
0 10126 7 4 2 46826 46952
0 10127 7 4 2 45784 46907
0 10128 7 1 2 47628 62905
0 10129 7 20 2 62901 10128
0 10130 7 1 2 56748 59256
0 10131 5 2 1 10130
0 10132 7 5 2 45707 56561
0 10133 5 2 1 62931
0 10134 7 1 2 62929 62936
0 10135 5 1 1 10134
0 10136 7 1 2 50938 10135
0 10137 5 1 1 10136
0 10138 7 1 2 52916 62793
0 10139 5 1 1 10138
0 10140 7 1 2 44036 51824
0 10141 5 1 1 10140
0 10142 7 1 2 10139 10141
0 10143 5 1 1 10142
0 10144 7 1 2 51748 10143
0 10145 5 1 1 10144
0 10146 7 1 2 10137 10145
0 10147 5 1 1 10146
0 10148 7 4 2 53254 62629
0 10149 7 1 2 10147 62938
0 10150 5 1 1 10149
0 10151 7 4 2 48581 60787
0 10152 5 2 1 62942
0 10153 7 2 2 43043 49486
0 10154 5 2 1 62948
0 10155 7 1 2 50836 62949
0 10156 5 1 1 10155
0 10157 7 1 2 62946 10156
0 10158 5 1 1 10157
0 10159 7 1 2 60979 10158
0 10160 5 1 1 10159
0 10161 7 1 2 43044 60834
0 10162 5 2 1 10161
0 10163 7 1 2 54350 62952
0 10164 5 3 1 10163
0 10165 7 4 2 48582 50406
0 10166 7 1 2 62954 62957
0 10167 5 1 1 10166
0 10168 7 3 2 51727 53255
0 10169 7 2 2 55361 62961
0 10170 5 2 1 62964
0 10171 7 1 2 10167 62966
0 10172 5 1 1 10171
0 10173 7 1 2 61138 10172
0 10174 5 1 1 10173
0 10175 7 1 2 10160 10174
0 10176 5 1 1 10175
0 10177 7 1 2 51901 10176
0 10178 5 1 1 10177
0 10179 7 1 2 46459 52421
0 10180 5 1 1 10179
0 10181 7 4 2 57389 57577
0 10182 5 1 1 62968
0 10183 7 1 2 10180 10182
0 10184 5 5 1 10183
0 10185 7 3 2 53256 61139
0 10186 7 1 2 59257 62977
0 10187 7 1 2 62972 10186
0 10188 5 1 1 10187
0 10189 7 1 2 10178 10188
0 10190 5 1 1 10189
0 10191 7 1 2 52037 10190
0 10192 5 1 1 10191
0 10193 7 1 2 10150 10192
0 10194 5 2 1 10193
0 10195 7 1 2 62909 62980
0 10196 5 1 1 10195
0 10197 7 1 2 10125 10196
0 10198 5 1 1 10197
0 10199 7 1 2 41996 10198
0 10200 5 1 1 10199
0 10201 7 2 2 53626 60317
0 10202 5 1 1 62982
0 10203 7 8 2 46953 62906
0 10204 7 1 2 43449 62984
0 10205 5 1 1 10204
0 10206 7 1 2 10202 10205
0 10207 5 12 1 10206
0 10208 7 1 2 59565 62992
0 10209 7 1 2 62981 10208
0 10210 5 1 1 10209
0 10211 7 1 2 10200 10210
0 10212 5 1 1 10211
0 10213 7 1 2 44432 10212
0 10214 5 1 1 10213
0 10215 7 1 2 52332 62725
0 10216 5 1 1 10215
0 10217 7 6 2 55793 60300
0 10218 7 1 2 59879 63004
0 10219 7 1 2 58368 10218
0 10220 5 1 1 10219
0 10221 7 1 2 10216 10220
0 10222 5 1 1 10221
0 10223 7 1 2 45546 10222
0 10224 5 1 1 10223
0 10225 7 2 2 59359 62993
0 10226 7 1 2 52333 63010
0 10227 5 1 1 10226
0 10228 7 1 2 10224 10227
0 10229 5 1 1 10228
0 10230 7 1 2 43045 10229
0 10231 5 1 1 10230
0 10232 7 2 2 41997 62994
0 10233 5 1 1 63012
0 10234 7 18 2 45547 42256
0 10235 7 5 2 62718 63014
0 10236 5 1 1 63032
0 10237 7 1 2 10233 10236
0 10238 5 4 1 10237
0 10239 7 13 2 44310 63037
0 10240 5 3 1 63041
0 10241 7 1 2 60835 63042
0 10242 5 1 1 10241
0 10243 7 1 2 10231 10242
0 10244 5 1 1 10243
0 10245 7 1 2 51902 10244
0 10246 5 1 1 10245
0 10247 7 1 2 60817 62910
0 10248 5 1 1 10247
0 10249 7 1 2 51749 62726
0 10250 5 1 1 10249
0 10251 7 1 2 10248 10250
0 10252 5 1 1 10251
0 10253 7 1 2 45548 10252
0 10254 5 1 1 10253
0 10255 7 1 2 51750 63011
0 10256 5 1 1 10255
0 10257 7 1 2 10254 10256
0 10258 5 1 1 10257
0 10259 7 1 2 59258 10258
0 10260 5 1 1 10259
0 10261 7 1 2 10246 10260
0 10262 5 1 1 10261
0 10263 7 1 2 51969 10262
0 10264 5 1 1 10263
0 10265 7 2 2 51202 62776
0 10266 5 1 1 63057
0 10267 7 1 2 43263 62782
0 10268 5 1 1 10267
0 10269 7 1 2 10266 10268
0 10270 5 1 1 10269
0 10271 7 1 2 43046 62858
0 10272 7 1 2 10270 10271
0 10273 7 1 2 63043 10272
0 10274 5 1 1 10273
0 10275 7 1 2 10264 10274
0 10276 5 1 1 10275
0 10277 7 1 2 48583 10276
0 10278 5 1 1 10277
0 10279 7 1 2 49335 51903
0 10280 7 1 2 63044 10279
0 10281 5 1 1 10280
0 10282 7 19 2 46908 46954
0 10283 7 2 2 61015 63059
0 10284 7 6 2 45785 44037
0 10285 7 1 2 57606 59997
0 10286 7 1 2 63080 10285
0 10287 7 1 2 63078 10286
0 10288 5 1 1 10287
0 10289 7 1 2 10281 10288
0 10290 5 1 1 10289
0 10291 7 1 2 49536 51970
0 10292 7 1 2 10290 10291
0 10293 5 1 1 10292
0 10294 7 1 2 10278 10293
0 10295 5 1 1 10294
0 10296 7 1 2 60374 10295
0 10297 5 1 1 10296
0 10298 7 11 2 47629 45215
0 10299 7 3 2 45549 63086
0 10300 7 1 2 63005 63097
0 10301 5 1 1 10300
0 10302 7 1 2 63054 10301
0 10303 5 1 1 10302
0 10304 7 1 2 51904 10303
0 10305 5 1 1 10304
0 10306 7 5 2 44556 45216
0 10307 7 2 2 47630 63100
0 10308 7 2 2 63060 63105
0 10309 7 18 2 45550 45786
0 10310 7 2 2 60669 63109
0 10311 7 1 2 63107 63127
0 10312 5 1 1 10311
0 10313 7 1 2 10305 10312
0 10314 5 1 1 10313
0 10315 7 1 2 45427 10314
0 10316 5 1 1 10315
0 10317 7 1 2 59259 63045
0 10318 5 1 1 10317
0 10319 7 1 2 10316 10318
0 10320 5 1 1 10319
0 10321 7 1 2 47528 10320
0 10322 5 1 1 10321
0 10323 7 8 2 42155 55706
0 10324 5 2 1 63129
0 10325 7 3 2 45217 51905
0 10326 5 1 1 63139
0 10327 7 1 2 63137 10326
0 10328 5 1 1 10327
0 10329 7 1 2 63046 10328
0 10330 5 1 1 10329
0 10331 7 1 2 10322 10330
0 10332 5 1 1 10331
0 10333 7 1 2 46648 10332
0 10334 5 1 1 10333
0 10335 7 1 2 51429 59260
0 10336 5 1 1 10335
0 10337 7 1 2 49105 51906
0 10338 5 1 1 10337
0 10339 7 1 2 10336 10338
0 10340 5 1 1 10339
0 10341 7 1 2 63047 10340
0 10342 5 1 1 10341
0 10343 7 1 2 10334 10342
0 10344 5 1 1 10343
0 10345 7 1 2 49275 10344
0 10346 5 1 1 10345
0 10347 7 2 2 51518 58680
0 10348 5 4 1 63142
0 10349 7 2 2 50755 62752
0 10350 5 1 1 63148
0 10351 7 1 2 63144 10350
0 10352 5 1 1 10351
0 10353 7 1 2 59807 10352
0 10354 7 1 2 63038 10353
0 10355 5 1 1 10354
0 10356 7 1 2 10346 10355
0 10357 5 1 1 10356
0 10358 7 1 2 62018 10357
0 10359 5 1 1 10358
0 10360 7 1 2 10297 10359
0 10361 5 1 1 10360
0 10362 7 1 2 53257 10361
0 10363 5 1 1 10362
0 10364 7 1 2 54229 59219
0 10365 5 1 1 10364
0 10366 7 1 2 57209 61806
0 10367 5 1 1 10366
0 10368 7 1 2 10365 10367
0 10369 5 1 1 10368
0 10370 7 1 2 54645 10369
0 10371 5 1 1 10370
0 10372 7 1 2 61713 10371
0 10373 5 1 1 10372
0 10374 7 1 2 48584 10373
0 10375 5 1 1 10374
0 10376 7 1 2 58805 61403
0 10377 5 1 1 10376
0 10378 7 1 2 10375 10377
0 10379 5 1 1 10378
0 10380 7 1 2 47234 10379
0 10381 5 1 1 10380
0 10382 7 9 2 48091 48796
0 10383 5 1 1 63150
0 10384 7 2 2 62124 63151
0 10385 7 1 2 42508 55100
0 10386 7 1 2 63159 10385
0 10387 5 1 1 10386
0 10388 7 1 2 46001 56777
0 10389 7 1 2 62223 10388
0 10390 5 1 1 10389
0 10391 7 1 2 10387 10390
0 10392 5 1 1 10391
0 10393 7 1 2 50994 10392
0 10394 5 1 1 10393
0 10395 7 1 2 46195 60761
0 10396 5 1 1 10395
0 10397 7 1 2 49276 62465
0 10398 5 1 1 10397
0 10399 7 1 2 10396 10398
0 10400 5 1 1 10399
0 10401 7 2 2 56634 61514
0 10402 7 1 2 10400 63161
0 10403 5 1 1 10402
0 10404 7 1 2 10394 10403
0 10405 7 1 2 10381 10404
0 10406 5 1 1 10405
0 10407 7 1 2 63048 10406
0 10408 5 1 1 10407
0 10409 7 1 2 52926 61690
0 10410 5 1 1 10409
0 10411 7 1 2 60980 10410
0 10412 5 1 1 10411
0 10413 7 1 2 55244 61188
0 10414 5 1 1 10413
0 10415 7 1 2 10412 10414
0 10416 5 1 1 10415
0 10417 7 3 2 45551 62911
0 10418 7 1 2 47235 57344
0 10419 7 1 2 63163 10418
0 10420 7 1 2 10416 10419
0 10421 5 1 1 10420
0 10422 7 1 2 44190 10421
0 10423 7 1 2 10408 10422
0 10424 5 1 1 10423
0 10425 7 3 2 44311 49745
0 10426 7 1 2 61404 63166
0 10427 7 1 2 63039 10426
0 10428 5 1 1 10427
0 10429 7 3 2 58394 61394
0 10430 5 1 1 63169
0 10431 7 1 2 60998 10430
0 10432 5 1 1 10431
0 10433 7 6 2 47631 63061
0 10434 7 4 2 46827 63110
0 10435 7 1 2 60944 63178
0 10436 7 1 2 63172 10435
0 10437 7 1 2 10432 10436
0 10438 5 1 1 10437
0 10439 7 1 2 10428 10438
0 10440 5 1 1 10439
0 10441 7 1 2 46460 10440
0 10442 5 1 1 10441
0 10443 7 1 2 50546 61405
0 10444 5 1 1 10443
0 10445 7 1 2 49901 61421
0 10446 5 1 1 10445
0 10447 7 1 2 10444 10446
0 10448 5 1 1 10447
0 10449 7 1 2 63049 10448
0 10450 5 1 1 10449
0 10451 7 1 2 43870 10450
0 10452 7 1 2 10442 10451
0 10453 5 1 1 10452
0 10454 7 1 2 52093 60981
0 10455 5 1 1 10454
0 10456 7 1 2 58094 61506
0 10457 7 1 2 54167 10456
0 10458 5 1 1 10457
0 10459 7 1 2 10455 10458
0 10460 5 1 1 10459
0 10461 7 1 2 63050 10460
0 10462 5 1 1 10461
0 10463 7 1 2 47236 10462
0 10464 5 1 1 10463
0 10465 7 1 2 45428 10464
0 10466 7 1 2 10453 10465
0 10467 5 1 1 10466
0 10468 7 1 2 3547 57173
0 10469 5 1 1 10468
0 10470 7 1 2 53754 10469
0 10471 5 1 1 10470
0 10472 7 1 2 49511 54109
0 10473 5 1 1 10472
0 10474 7 1 2 53965 54892
0 10475 5 1 1 10474
0 10476 7 1 2 10473 10475
0 10477 7 1 2 10471 10476
0 10478 5 1 1 10477
0 10479 7 1 2 63170 10478
0 10480 7 1 2 63051 10479
0 10481 5 1 1 10480
0 10482 7 1 2 47529 10481
0 10483 7 1 2 10467 10482
0 10484 5 1 1 10483
0 10485 7 1 2 10424 10484
0 10486 5 1 1 10485
0 10487 7 1 2 58268 59566
0 10488 7 1 2 60301 61922
0 10489 7 1 2 10487 10488
0 10490 7 1 2 50153 57531
0 10491 7 1 2 61189 10490
0 10492 7 1 2 10489 10491
0 10493 5 1 1 10492
0 10494 7 1 2 48585 52992
0 10495 5 1 1 10494
0 10496 7 1 2 2376 10495
0 10497 5 1 1 10496
0 10498 7 1 2 61412 10497
0 10499 7 1 2 63052 10498
0 10500 5 1 1 10499
0 10501 7 1 2 10493 10500
0 10502 5 1 1 10501
0 10503 7 1 2 49205 10502
0 10504 5 1 1 10503
0 10505 7 3 2 58433 61725
0 10506 5 1 1 63182
0 10507 7 1 2 51457 51971
0 10508 7 1 2 63183 10507
0 10509 5 1 1 10508
0 10510 7 1 2 55182 57246
0 10511 7 1 2 52942 10510
0 10512 7 1 2 62562 10511
0 10513 5 1 1 10512
0 10514 7 1 2 10509 10513
0 10515 5 1 1 10514
0 10516 7 1 2 62912 10515
0 10517 5 1 1 10516
0 10518 7 13 2 44312 55751
0 10519 7 2 2 60318 63185
0 10520 7 1 2 63184 63198
0 10521 7 1 2 61967 10520
0 10522 5 1 1 10521
0 10523 7 1 2 10517 10522
0 10524 5 1 1 10523
0 10525 7 1 2 45552 10524
0 10526 5 1 1 10525
0 10527 7 1 2 60142 61570
0 10528 7 1 2 61968 10527
0 10529 7 1 2 63013 10528
0 10530 5 1 1 10529
0 10531 7 1 2 10526 10530
0 10532 5 1 1 10531
0 10533 7 1 2 49078 10532
0 10534 5 1 1 10533
0 10535 7 1 2 55167 57175
0 10536 5 3 1 10535
0 10537 7 1 2 46461 63200
0 10538 5 2 1 10537
0 10539 7 2 2 63203 62894
0 10540 5 1 1 63205
0 10541 7 1 2 61400 10540
0 10542 5 1 1 10541
0 10543 7 2 2 54133 55149
0 10544 7 9 2 43871 48092
0 10545 7 1 2 55441 63209
0 10546 7 1 2 63207 10545
0 10547 5 1 1 10546
0 10548 7 1 2 10542 10547
0 10549 5 1 1 10548
0 10550 7 1 2 63053 10549
0 10551 5 1 1 10550
0 10552 7 7 2 45787 43047
0 10553 7 1 2 58182 63218
0 10554 7 8 2 46955 44635
0 10555 5 2 1 63225
0 10556 7 5 2 42509 47632
0 10557 7 1 2 63226 63235
0 10558 7 1 2 10553 10557
0 10559 7 2 2 46196 52934
0 10560 7 1 2 55665 56610
0 10561 7 1 2 63240 10560
0 10562 7 1 2 10558 10561
0 10563 5 1 1 10562
0 10564 7 1 2 10551 10563
0 10565 7 1 2 10534 10564
0 10566 7 1 2 10504 10565
0 10567 7 1 2 10486 10566
0 10568 5 1 1 10567
0 10569 7 1 2 59261 10568
0 10570 5 1 1 10569
0 10571 7 1 2 10363 10570
0 10572 5 1 1 10571
0 10573 7 1 2 47745 10572
0 10574 5 1 1 10573
0 10575 7 4 2 48093 62023
0 10576 7 7 2 42257 43048
0 10577 7 2 2 59954 63246
0 10578 7 2 2 59328 62702
0 10579 7 1 2 61950 63255
0 10580 7 1 2 63253 10579
0 10581 5 1 1 10580
0 10582 7 6 2 48586 50995
0 10583 5 1 1 63257
0 10584 7 1 2 63164 63258
0 10585 5 1 1 10584
0 10586 7 1 2 63055 10585
0 10587 5 1 1 10586
0 10588 7 2 2 43713 47746
0 10589 7 1 2 46649 63263
0 10590 7 1 2 10587 10589
0 10591 5 1 1 10590
0 10592 7 1 2 10581 10591
0 10593 5 1 1 10592
0 10594 7 1 2 49079 10593
0 10595 5 1 1 10594
0 10596 7 1 2 44038 50307
0 10597 5 3 1 10596
0 10598 7 1 2 49524 63265
0 10599 5 1 1 10598
0 10600 7 1 2 51193 10599
0 10601 5 1 1 10600
0 10602 7 2 2 47404 59031
0 10603 5 2 1 63268
0 10604 7 2 2 44039 50173
0 10605 5 1 1 63272
0 10606 7 1 2 45218 10605
0 10607 7 1 2 63270 10606
0 10608 7 1 2 10601 10607
0 10609 5 1 1 10608
0 10610 7 1 2 52715 63165
0 10611 7 1 2 10609 10610
0 10612 5 1 1 10611
0 10613 7 1 2 63056 10612
0 10614 5 1 1 10613
0 10615 7 1 2 51430 63264
0 10616 7 1 2 10614 10615
0 10617 5 1 1 10616
0 10618 7 3 2 44040 44433
0 10619 7 7 2 43571 44313
0 10620 7 1 2 63274 63277
0 10621 7 1 2 51424 10620
0 10622 7 4 2 42258 50154
0 10623 7 1 2 59691 63284
0 10624 7 1 2 10621 10623
0 10625 5 1 1 10624
0 10626 7 1 2 10617 10625
0 10627 7 1 2 10595 10626
0 10628 5 1 1 10627
0 10629 7 1 2 63242 10628
0 10630 5 1 1 10629
0 10631 7 13 2 45788 46002
0 10632 7 4 2 45553 63288
0 10633 7 1 2 56483 61005
0 10634 7 2 2 63301 10633
0 10635 7 9 2 46828 63062
0 10636 7 1 2 60120 63307
0 10637 7 1 2 63305 10636
0 10638 5 1 1 10637
0 10639 7 2 2 43714 62703
0 10640 7 1 2 62080 63316
0 10641 7 5 2 42259 43450
0 10642 7 2 2 41998 63318
0 10643 7 2 2 44041 61289
0 10644 7 1 2 63323 63325
0 10645 7 1 2 10640 10644
0 10646 5 1 1 10645
0 10647 7 1 2 10638 10646
0 10648 5 2 1 10647
0 10649 7 1 2 59100 63327
0 10650 5 1 1 10649
0 10651 7 4 2 47747 50407
0 10652 7 1 2 62983 63329
0 10653 5 1 1 10652
0 10654 7 1 2 46909 56409
0 10655 7 5 2 46003 43451
0 10656 7 1 2 60302 63333
0 10657 7 1 2 10654 10656
0 10658 5 1 1 10657
0 10659 7 1 2 10653 10658
0 10660 5 1 1 10659
0 10661 7 1 2 41999 10660
0 10662 5 1 1 10661
0 10663 7 1 2 63033 63330
0 10664 5 1 1 10663
0 10665 7 1 2 10662 10664
0 10666 5 1 1 10665
0 10667 7 1 2 60224 10666
0 10668 5 1 1 10667
0 10669 7 9 2 42260 43526
0 10670 5 1 1 63338
0 10671 7 4 2 43572 63339
0 10672 7 2 2 47405 62483
0 10673 5 1 1 63351
0 10674 7 1 2 52192 63352
0 10675 7 1 2 63347 10674
0 10676 7 1 2 59975 10675
0 10677 5 1 1 10676
0 10678 7 1 2 10668 10677
0 10679 5 1 1 10678
0 10680 7 1 2 44314 10679
0 10681 5 1 1 10680
0 10682 7 3 2 48998 56888
0 10683 5 3 1 63353
0 10684 7 2 2 55610 63354
0 10685 7 1 2 58529 63173
0 10686 7 1 2 63302 10685
0 10687 7 1 2 63359 10686
0 10688 5 1 1 10687
0 10689 7 1 2 10681 10688
0 10690 5 1 1 10689
0 10691 7 1 2 61140 10690
0 10692 5 1 1 10691
0 10693 7 1 2 10650 10692
0 10694 7 1 2 10630 10693
0 10695 5 1 1 10694
0 10696 7 1 2 59262 10695
0 10697 5 1 1 10696
0 10698 7 2 2 45554 62995
0 10699 5 1 1 63361
0 10700 7 3 2 54741 62985
0 10701 5 1 1 63363
0 10702 7 1 2 10699 10701
0 10703 5 2 1 10702
0 10704 7 1 2 50211 58395
0 10705 7 1 2 59880 10704
0 10706 5 1 1 10705
0 10707 7 1 2 49336 59749
0 10708 7 1 2 61939 10707
0 10709 5 1 1 10708
0 10710 7 1 2 10706 10709
0 10711 5 1 1 10710
0 10712 7 1 2 63366 10711
0 10713 5 1 1 10712
0 10714 7 4 2 47633 63367
0 10715 7 9 2 47090 44042
0 10716 7 1 2 63368 63372
0 10717 5 1 1 10716
0 10718 7 4 2 43573 45429
0 10719 7 9 2 42261 46462
0 10720 7 4 2 47406 44315
0 10721 7 1 2 63385 63394
0 10722 7 1 2 63381 10721
0 10723 7 1 2 59692 10722
0 10724 5 1 1 10723
0 10725 7 1 2 10717 10724
0 10726 5 1 1 10725
0 10727 7 1 2 46004 10726
0 10728 5 1 1 10727
0 10729 7 8 2 42000 42262
0 10730 7 7 2 44316 63398
0 10731 7 2 2 47407 63406
0 10732 7 11 2 43452 43574
0 10733 7 4 2 55638 63415
0 10734 7 1 2 50212 63426
0 10735 7 1 2 63413 10734
0 10736 5 1 1 10735
0 10737 7 1 2 10728 10736
0 10738 5 1 1 10737
0 10739 7 1 2 50756 10738
0 10740 5 1 1 10739
0 10741 7 1 2 10713 10740
0 10742 5 1 1 10741
0 10743 7 1 2 61141 10742
0 10744 5 1 1 10743
0 10745 7 1 2 51714 51877
0 10746 5 1 1 10745
0 10747 7 2 2 9352 10746
0 10748 7 1 2 53498 63430
0 10749 5 1 1 10748
0 10750 7 1 2 60982 10749
0 10751 7 1 2 63369 10750
0 10752 5 1 1 10751
0 10753 7 1 2 10744 10752
0 10754 5 1 1 10753
0 10755 7 1 2 45219 10754
0 10756 5 1 1 10755
0 10757 7 3 2 51751 60375
0 10758 7 1 2 63208 63432
0 10759 5 1 1 10758
0 10760 7 1 2 47530 57838
0 10761 7 1 2 63171 10760
0 10762 5 1 1 10761
0 10763 7 1 2 10759 10762
0 10764 5 1 1 10763
0 10765 7 1 2 63370 10764
0 10766 5 1 1 10765
0 10767 7 2 2 46910 60156
0 10768 7 2 2 60303 63435
0 10769 7 1 2 61551 63437
0 10770 5 1 1 10769
0 10771 7 6 2 63340 63416
0 10772 7 2 2 43049 63439
0 10773 7 1 2 59329 61795
0 10774 7 2 2 63445 10773
0 10775 5 1 1 63447
0 10776 7 1 2 10770 10775
0 10777 5 1 1 10776
0 10778 7 1 2 42001 10777
0 10779 5 1 1 10778
0 10780 7 1 2 61190 61549
0 10781 7 1 2 63362 10780
0 10782 5 1 1 10781
0 10783 7 1 2 10779 10782
0 10784 5 1 1 10783
0 10785 7 1 2 55569 10784
0 10786 5 1 1 10785
0 10787 7 1 2 51222 60983
0 10788 5 1 1 10787
0 10789 7 3 2 44749 50837
0 10790 7 1 2 51065 61507
0 10791 7 1 2 63449 10790
0 10792 5 1 1 10791
0 10793 7 1 2 10788 10792
0 10794 5 1 1 10793
0 10795 7 1 2 46463 10794
0 10796 5 1 1 10795
0 10797 7 7 2 46650 47965
0 10798 7 2 2 62154 63452
0 10799 7 5 2 47091 47408
0 10800 7 1 2 57434 63461
0 10801 7 1 2 63459 10800
0 10802 5 1 1 10801
0 10803 7 1 2 10796 10802
0 10804 5 1 1 10803
0 10805 7 1 2 63371 10804
0 10806 5 1 1 10805
0 10807 7 4 2 42002 43715
0 10808 7 1 2 51385 52831
0 10809 7 1 2 63466 10808
0 10810 7 2 2 59237 63417
0 10811 7 2 2 61564 63247
0 10812 7 1 2 63470 63472
0 10813 7 1 2 10809 10812
0 10814 5 1 1 10813
0 10815 7 1 2 10806 10814
0 10816 7 1 2 10786 10815
0 10817 5 1 1 10816
0 10818 7 1 2 48587 10817
0 10819 5 1 1 10818
0 10820 7 1 2 10766 10819
0 10821 7 1 2 10756 10820
0 10822 5 1 1 10821
0 10823 7 1 2 44434 51907
0 10824 7 1 2 10822 10823
0 10825 5 1 1 10824
0 10826 7 1 2 10697 10825
0 10827 5 1 1 10826
0 10828 7 1 2 60278 10827
0 10829 5 1 1 10828
0 10830 7 1 2 54230 62484
0 10831 5 1 1 10830
0 10832 7 5 2 47748 61079
0 10833 7 2 2 48797 63474
0 10834 5 1 1 63479
0 10835 7 1 2 10831 10834
0 10836 5 1 1 10835
0 10837 7 1 2 44191 10836
0 10838 5 1 1 10837
0 10839 7 2 2 42747 53755
0 10840 5 3 1 63481
0 10841 7 1 2 44043 60443
0 10842 7 1 2 63483 10841
0 10843 5 1 1 10842
0 10844 7 1 2 10838 10843
0 10845 5 1 1 10844
0 10846 7 1 2 43264 10845
0 10847 5 1 1 10846
0 10848 7 1 2 51881 56893
0 10849 5 1 1 10848
0 10850 7 1 2 62485 10849
0 10851 5 1 1 10850
0 10852 7 1 2 10847 10851
0 10853 5 1 1 10852
0 10854 7 1 2 47237 10853
0 10855 5 1 1 10854
0 10856 7 2 2 49964 62486
0 10857 5 1 1 63486
0 10858 7 1 2 54958 63487
0 10859 5 1 1 10858
0 10860 7 1 2 55199 60444
0 10861 5 1 1 10860
0 10862 7 1 2 62550 10861
0 10863 5 1 1 10862
0 10864 7 2 2 57322 57345
0 10865 5 1 1 63488
0 10866 7 1 2 47238 49122
0 10867 5 1 1 10866
0 10868 7 1 2 10865 10867
0 10869 5 1 1 10868
0 10870 7 1 2 10863 10869
0 10871 5 1 1 10870
0 10872 7 1 2 10859 10871
0 10873 7 1 2 10855 10872
0 10874 5 1 1 10873
0 10875 7 1 2 48588 10874
0 10876 5 1 1 10875
0 10877 7 7 2 43050 49965
0 10878 5 4 1 63490
0 10879 7 2 2 46197 63497
0 10880 5 2 1 63501
0 10881 7 1 2 45220 63503
0 10882 5 3 1 10881
0 10883 7 1 2 57825 63505
0 10884 5 2 1 10883
0 10885 7 1 2 62487 63508
0 10886 5 1 1 10885
0 10887 7 2 2 49156 55375
0 10888 5 5 1 63510
0 10889 7 2 2 46198 49206
0 10890 5 1 1 63517
0 10891 7 1 2 62303 10890
0 10892 5 2 1 10891
0 10893 7 1 2 44044 63519
0 10894 5 1 1 10893
0 10895 7 1 2 63512 10894
0 10896 5 1 1 10895
0 10897 7 1 2 48589 10896
0 10898 5 1 1 10897
0 10899 7 1 2 60193 63513
0 10900 5 1 1 10899
0 10901 7 1 2 43051 10900
0 10902 5 2 1 10901
0 10903 7 1 2 46199 54351
0 10904 5 2 1 10903
0 10905 7 4 2 43265 50547
0 10906 5 3 1 63525
0 10907 7 1 2 42748 49247
0 10908 7 1 2 63529 10907
0 10909 5 1 1 10908
0 10910 7 1 2 63523 10909
0 10911 5 1 1 10910
0 10912 7 1 2 63521 10911
0 10913 7 1 2 10898 10912
0 10914 5 1 1 10913
0 10915 7 1 2 60445 10914
0 10916 5 1 1 10915
0 10917 7 1 2 10886 10916
0 10918 5 1 1 10917
0 10919 7 1 2 47239 10918
0 10920 5 1 1 10919
0 10921 7 1 2 10876 10920
0 10922 5 1 1 10921
0 10923 7 1 2 51908 10922
0 10924 5 1 1 10923
0 10925 7 1 2 42749 49549
0 10926 5 3 1 10925
0 10927 7 1 2 50605 51788
0 10928 5 1 1 10927
0 10929 7 2 2 46651 49688
0 10930 5 2 1 63535
0 10931 7 1 2 61681 63537
0 10932 7 1 2 10928 10931
0 10933 7 1 2 63532 10932
0 10934 5 1 1 10933
0 10935 7 11 2 55775 56230
0 10936 7 1 2 47240 63539
0 10937 7 1 2 10934 10936
0 10938 5 1 1 10937
0 10939 7 1 2 10924 10938
0 10940 5 1 1 10939
0 10941 7 1 2 62727 10940
0 10942 5 1 1 10941
0 10943 7 7 2 44317 57025
0 10944 7 1 2 60164 60249
0 10945 5 2 1 10944
0 10946 7 2 2 63550 63557
0 10947 7 1 2 59012 63559
0 10948 5 1 1 10947
0 10949 7 2 2 49966 51909
0 10950 5 1 1 63561
0 10951 7 1 2 50548 63562
0 10952 5 1 1 10951
0 10953 7 1 2 58784 58554
0 10954 5 2 1 10953
0 10955 7 1 2 59263 63563
0 10956 5 1 1 10955
0 10957 7 1 2 10952 10956
0 10958 5 1 1 10957
0 10959 7 1 2 60525 10958
0 10960 5 1 1 10959
0 10961 7 1 2 10948 10960
0 10962 5 1 1 10961
0 10963 7 1 2 46200 10962
0 10964 5 1 1 10963
0 10965 7 6 2 47883 60634
0 10966 7 7 2 59013 63565
0 10967 5 1 1 63571
0 10968 7 1 2 54984 63572
0 10969 5 1 1 10968
0 10970 7 3 2 60802 61016
0 10971 7 1 2 43052 63578
0 10972 5 1 1 10971
0 10973 7 1 2 10969 10972
0 10974 5 1 1 10973
0 10975 7 1 2 62969 10974
0 10976 5 1 1 10975
0 10977 7 1 2 43872 10976
0 10978 7 1 2 10964 10977
0 10979 5 1 1 10978
0 10980 7 2 2 42750 56749
0 10981 5 1 1 63581
0 10982 7 1 2 46201 56849
0 10983 5 1 1 10982
0 10984 7 1 2 10981 10983
0 10985 5 1 1 10984
0 10986 7 1 2 49253 10985
0 10987 5 1 1 10986
0 10988 7 1 2 43053 10987
0 10989 5 1 1 10988
0 10990 7 2 2 49967 53725
0 10991 7 1 2 53029 63583
0 10992 5 1 1 10991
0 10993 7 1 2 10989 10992
0 10994 5 2 1 10993
0 10995 7 1 2 63579 63585
0 10996 5 1 1 10995
0 10997 7 2 2 59360 60415
0 10998 7 1 2 62037 63587
0 10999 5 1 1 10998
0 11000 7 6 2 53030 53420
0 11001 7 1 2 62585 63589
0 11002 5 1 1 11001
0 11003 7 1 2 10999 11002
0 11004 5 1 1 11003
0 11005 7 1 2 44192 11004
0 11006 5 1 1 11005
0 11007 7 2 2 46202 49689
0 11008 5 4 1 63595
0 11009 7 1 2 60947 63597
0 11010 5 19 1 11009
0 11011 7 1 2 61642 63601
0 11012 5 1 1 11011
0 11013 7 1 2 11006 11012
0 11014 5 1 1 11013
0 11015 7 1 2 43266 11014
0 11016 5 1 1 11015
0 11017 7 1 2 48590 63520
0 11018 5 1 1 11017
0 11019 7 1 2 11018 63514
0 11020 5 1 1 11019
0 11021 7 1 2 44045 11020
0 11022 5 2 1 11021
0 11023 7 2 2 49157 58574
0 11024 5 4 1 63622
0 11025 7 1 2 55376 63623
0 11026 5 1 1 11025
0 11027 7 2 2 63620 11026
0 11028 5 1 1 63628
0 11029 7 1 2 59380 11028
0 11030 5 1 1 11029
0 11031 7 1 2 11016 11030
0 11032 5 1 1 11031
0 11033 7 1 2 51910 11032
0 11034 5 1 1 11033
0 11035 7 1 2 47241 11034
0 11036 7 1 2 10996 11035
0 11037 5 1 1 11036
0 11038 7 1 2 10979 11037
0 11039 5 1 1 11038
0 11040 7 1 2 51789 63573
0 11041 5 3 1 11040
0 11042 7 4 2 45555 59174
0 11043 7 1 2 62828 63633
0 11044 5 1 1 11043
0 11045 7 1 2 63630 11044
0 11046 5 1 1 11045
0 11047 7 1 2 60279 11046
0 11048 5 1 1 11047
0 11049 7 3 2 63130 63634
0 11050 5 1 1 63637
0 11051 7 2 2 43267 63638
0 11052 5 1 1 63640
0 11053 7 1 2 55158 63641
0 11054 5 1 1 11053
0 11055 7 1 2 11048 11054
0 11056 5 1 1 11055
0 11057 7 1 2 49746 11056
0 11058 5 1 1 11057
0 11059 7 1 2 63631 11052
0 11060 5 1 1 11059
0 11061 7 1 2 63201 11060
0 11062 5 1 1 11061
0 11063 7 1 2 57346 61643
0 11064 7 1 2 57157 11063
0 11065 5 1 1 11064
0 11066 7 2 2 44435 57861
0 11067 7 2 2 47634 61447
0 11068 7 1 2 53966 63644
0 11069 7 1 2 63642 11068
0 11070 5 1 1 11069
0 11071 7 1 2 11065 11070
0 11072 5 1 1 11071
0 11073 7 1 2 51911 11072
0 11074 5 1 1 11073
0 11075 7 1 2 60265 60948
0 11076 5 2 1 11075
0 11077 7 8 2 44557 50063
0 11078 7 2 2 42156 63648
0 11079 5 2 1 63656
0 11080 7 1 2 54122 60526
0 11081 7 1 2 63657 11080
0 11082 7 1 2 63646 11081
0 11083 5 1 1 11082
0 11084 7 1 2 11074 11083
0 11085 7 1 2 11062 11084
0 11086 5 1 1 11085
0 11087 7 1 2 46464 11086
0 11088 5 1 1 11087
0 11089 7 1 2 11058 11088
0 11090 7 1 2 11039 11089
0 11091 5 1 1 11090
0 11092 7 1 2 62996 11091
0 11093 5 1 1 11092
0 11094 7 7 2 47242 47635
0 11095 7 2 2 63006 63660
0 11096 7 2 2 52221 63540
0 11097 5 1 1 63669
0 11098 7 1 2 62930 10950
0 11099 5 1 1 11098
0 11100 7 1 2 62488 11099
0 11101 5 1 1 11100
0 11102 7 5 2 57026 61261
0 11103 7 1 2 45430 52246
0 11104 7 1 2 63671 11103
0 11105 5 1 1 11104
0 11106 7 1 2 11101 11105
0 11107 5 1 1 11106
0 11108 7 1 2 43054 11107
0 11109 5 1 1 11108
0 11110 7 1 2 11097 11109
0 11111 5 1 1 11110
0 11112 7 1 2 46203 11111
0 11113 5 1 1 11112
0 11114 7 3 2 43055 50757
0 11115 5 3 1 63676
0 11116 7 1 2 53499 63679
0 11117 5 9 1 11116
0 11118 7 7 2 45431 63682
0 11119 7 1 2 60258 61765
0 11120 7 1 2 63691 11119
0 11121 5 1 1 11120
0 11122 7 1 2 11113 11121
0 11123 5 1 1 11122
0 11124 7 1 2 44046 11123
0 11125 5 1 1 11124
0 11126 7 1 2 56209 63670
0 11127 5 1 1 11126
0 11128 7 11 2 45556 61579
0 11129 5 1 1 63698
0 11130 7 1 2 50758 54862
0 11131 5 4 1 11130
0 11132 7 1 2 52813 61460
0 11133 5 1 1 11132
0 11134 7 1 2 63709 11133
0 11135 5 4 1 11134
0 11136 7 1 2 63699 63713
0 11137 5 1 1 11136
0 11138 7 3 2 42003 58919
0 11139 7 1 2 63526 63717
0 11140 5 1 1 11139
0 11141 7 1 2 11137 11140
0 11142 5 1 1 11141
0 11143 7 1 2 51912 11142
0 11144 5 1 1 11143
0 11145 7 1 2 58550 58584
0 11146 5 1 1 11145
0 11147 7 1 2 63541 11146
0 11148 5 1 1 11147
0 11149 7 1 2 11144 11148
0 11150 5 1 1 11149
0 11151 7 1 2 42751 11150
0 11152 5 1 1 11151
0 11153 7 1 2 11127 11152
0 11154 7 1 2 11125 11153
0 11155 5 1 1 11154
0 11156 7 1 2 63667 11155
0 11157 5 1 1 11156
0 11158 7 1 2 51790 63475
0 11159 5 1 1 11158
0 11160 7 5 2 50064 62489
0 11161 5 1 1 63720
0 11162 7 1 2 46465 63721
0 11163 5 1 1 11162
0 11164 7 1 2 11159 11163
0 11165 5 1 1 11164
0 11166 7 1 2 43873 11165
0 11167 5 1 1 11166
0 11168 7 1 2 56937 61448
0 11169 7 1 2 51791 11168
0 11170 5 1 1 11169
0 11171 7 1 2 11167 11170
0 11172 5 1 1 11171
0 11173 7 1 2 51913 11172
0 11174 5 1 1 11173
0 11175 7 1 2 52000 52294
0 11176 5 1 1 11175
0 11177 7 1 2 56792 11176
0 11178 5 1 1 11177
0 11179 7 1 2 63542 11178
0 11180 5 1 1 11179
0 11181 7 1 2 11174 11180
0 11182 5 1 1 11181
0 11183 7 1 2 62728 11182
0 11184 5 1 1 11183
0 11185 7 1 2 46956 49525
0 11186 7 1 2 52055 11185
0 11187 7 22 2 42157 45789
0 11188 5 1 1 63725
0 11189 7 2 2 61870 63726
0 11190 7 1 2 52989 63747
0 11191 7 8 2 46911 47636
0 11192 7 5 2 44558 63749
0 11193 7 2 2 44436 60423
0 11194 7 1 2 63757 63762
0 11195 7 1 2 11190 11194
0 11196 7 1 2 11186 11195
0 11197 5 1 1 11196
0 11198 7 1 2 11184 11197
0 11199 5 1 1 11198
0 11200 7 1 2 49747 11199
0 11201 5 1 1 11200
0 11202 7 1 2 63167 63440
0 11203 5 1 1 11202
0 11204 7 6 2 45790 46829
0 11205 7 1 2 51397 63764
0 11206 7 2 2 63750 11205
0 11207 7 1 2 46957 48798
0 11208 7 2 2 63770 11207
0 11209 5 1 1 63772
0 11210 7 1 2 47409 63773
0 11211 5 1 1 11210
0 11212 7 1 2 11203 11211
0 11213 5 1 1 11212
0 11214 7 1 2 63672 11213
0 11215 5 1 1 11214
0 11216 7 2 2 53559 60304
0 11217 5 1 1 63774
0 11218 7 3 2 54742 63775
0 11219 7 1 2 52846 60803
0 11220 7 1 2 63776 11219
0 11221 5 1 1 11220
0 11222 7 1 2 11215 11221
0 11223 5 1 1 11222
0 11224 7 1 2 42752 11223
0 11225 5 1 1 11224
0 11226 7 3 2 55776 62704
0 11227 7 1 2 50606 62696
0 11228 7 1 2 59595 11227
0 11229 7 1 2 63779 11228
0 11230 5 1 1 11229
0 11231 7 1 2 11225 11230
0 11232 5 1 1 11231
0 11233 7 1 2 47243 11232
0 11234 5 1 1 11233
0 11235 7 6 2 44437 57782
0 11236 7 3 2 47637 53627
0 11237 7 1 2 63782 63788
0 11238 5 1 1 11237
0 11239 7 1 2 53643 63551
0 11240 5 1 1 11239
0 11241 7 1 2 11238 11240
0 11242 5 1 1 11241
0 11243 7 2 2 60319 61017
0 11244 5 1 1 63791
0 11245 7 13 2 45708 45791
0 11246 7 5 2 42004 46958
0 11247 7 2 2 63793 63806
0 11248 5 1 1 63811
0 11249 7 1 2 11244 11248
0 11250 5 1 1 11249
0 11251 7 1 2 11242 11250
0 11252 5 1 1 11251
0 11253 7 1 2 63751 63783
0 11254 5 1 1 11253
0 11255 7 5 2 55957 60635
0 11256 5 2 1 63813
0 11257 7 1 2 11254 63818
0 11258 5 1 1 11257
0 11259 7 1 2 45709 60320
0 11260 5 1 1 11259
0 11261 7 1 2 42158 60305
0 11262 5 1 1 11261
0 11263 7 1 2 11260 11262
0 11264 5 3 1 11263
0 11265 7 1 2 54761 63820
0 11266 7 1 2 11258 11265
0 11267 5 1 1 11266
0 11268 7 1 2 46959 61279
0 11269 7 2 2 45792 55752
0 11270 7 1 2 63823 63784
0 11271 7 1 2 11268 11270
0 11272 5 1 1 11271
0 11273 7 14 2 42263 46830
0 11274 5 1 1 63825
0 11275 7 1 2 56231 62666
0 11276 7 1 2 63826 11275
0 11277 7 1 2 63566 11276
0 11278 5 1 1 11277
0 11279 7 1 2 11272 11278
0 11280 7 1 2 11267 11279
0 11281 7 1 2 11252 11280
0 11282 5 1 1 11281
0 11283 7 1 2 46466 11282
0 11284 5 1 1 11283
0 11285 7 1 2 46204 57607
0 11286 7 2 2 63174 11285
0 11287 7 3 2 47749 55420
0 11288 7 2 2 61262 63841
0 11289 7 1 2 45793 63844
0 11290 7 1 2 63839 11289
0 11291 5 1 1 11290
0 11292 7 1 2 11284 11291
0 11293 5 1 1 11292
0 11294 7 1 2 57182 11293
0 11295 5 1 1 11294
0 11296 7 2 2 59148 60912
0 11297 7 3 2 52847 58002
0 11298 7 1 2 63846 63848
0 11299 5 1 1 11298
0 11300 7 8 2 42159 63567
0 11301 7 1 2 49748 60280
0 11302 5 3 1 11301
0 11303 7 1 2 9640 63859
0 11304 5 2 1 11303
0 11305 7 1 2 63851 63862
0 11306 5 1 1 11305
0 11307 7 1 2 11299 11306
0 11308 5 1 1 11307
0 11309 7 1 2 54762 62682
0 11310 7 1 2 11308 11309
0 11311 5 1 1 11310
0 11312 7 1 2 63574 63863
0 11313 5 1 1 11312
0 11314 7 1 2 56199 60527
0 11315 7 1 2 63849 11314
0 11316 5 1 1 11315
0 11317 7 1 2 11313 11316
0 11318 5 1 1 11317
0 11319 7 1 2 62997 11318
0 11320 5 1 1 11319
0 11321 7 1 2 55159 62705
0 11322 7 1 2 63568 11321
0 11323 7 3 2 58994 63015
0 11324 7 2 2 43056 49690
0 11325 5 2 1 63867
0 11326 7 1 2 63864 63869
0 11327 7 1 2 11322 11326
0 11328 5 1 1 11327
0 11329 7 1 2 11320 11328
0 11330 7 1 2 11311 11329
0 11331 7 1 2 11295 11330
0 11332 7 1 2 11234 11331
0 11333 5 1 1 11332
0 11334 7 1 2 55570 11333
0 11335 5 1 1 11334
0 11336 7 1 2 11201 11335
0 11337 7 1 2 11157 11336
0 11338 7 1 2 11093 11337
0 11339 7 1 2 10942 11338
0 11340 7 1 2 60611 63586
0 11341 5 1 1 11340
0 11342 7 1 2 50549 60711
0 11343 5 3 1 11342
0 11344 7 1 2 46205 59765
0 11345 5 2 1 11344
0 11346 7 1 2 63871 63874
0 11347 5 1 1 11346
0 11348 7 1 2 43268 11347
0 11349 5 1 1 11348
0 11350 7 2 2 63629 11349
0 11351 5 1 1 63876
0 11352 7 1 2 63852 11351
0 11353 5 1 1 11352
0 11354 7 1 2 11341 11353
0 11355 5 1 1 11354
0 11356 7 1 2 47244 11355
0 11357 5 1 1 11356
0 11358 7 1 2 42160 63560
0 11359 5 1 1 11358
0 11360 7 1 2 60612 63564
0 11361 5 1 1 11360
0 11362 7 1 2 11359 11361
0 11363 5 1 1 11362
0 11364 7 1 2 46206 11363
0 11365 5 1 1 11364
0 11366 7 2 2 51815 59423
0 11367 5 1 1 63878
0 11368 7 1 2 42161 54985
0 11369 7 1 2 63552 11368
0 11370 5 1 1 11369
0 11371 7 1 2 11367 11370
0 11372 5 1 1 11371
0 11373 7 1 2 62970 11372
0 11374 5 1 1 11373
0 11375 7 1 2 11365 11374
0 11376 5 1 1 11375
0 11377 7 1 2 43874 11376
0 11378 5 1 1 11377
0 11379 7 1 2 51792 61224
0 11380 5 2 1 11379
0 11381 7 3 2 45710 53357
0 11382 7 1 2 55777 60924
0 11383 7 1 2 63882 11382
0 11384 5 1 1 11383
0 11385 7 1 2 63880 11384
0 11386 5 1 1 11385
0 11387 7 1 2 60281 11386
0 11388 5 1 1 11387
0 11389 7 2 2 60925 61587
0 11390 7 1 2 58304 61632
0 11391 7 1 2 63885 11390
0 11392 5 1 1 11391
0 11393 7 1 2 11388 11392
0 11394 5 1 1 11393
0 11395 7 1 2 49749 11394
0 11396 5 1 1 11395
0 11397 7 1 2 57159 63853
0 11398 5 1 1 11397
0 11399 7 1 2 53475 60592
0 11400 7 1 2 63649 11399
0 11401 5 1 1 11400
0 11402 7 1 2 11398 11401
0 11403 5 1 1 11402
0 11404 7 1 2 46207 11403
0 11405 5 1 1 11404
0 11406 7 2 2 55707 59149
0 11407 7 1 2 60863 63887
0 11408 5 1 1 11407
0 11409 7 1 2 63881 11408
0 11410 5 1 1 11409
0 11411 7 1 2 63202 11410
0 11412 5 1 1 11411
0 11413 7 1 2 53379 53952
0 11414 7 1 2 63650 63847
0 11415 7 1 2 11413 11414
0 11416 5 1 1 11415
0 11417 7 1 2 11412 11416
0 11418 7 1 2 11405 11417
0 11419 5 1 1 11418
0 11420 7 1 2 46467 11419
0 11421 5 1 1 11420
0 11422 7 1 2 11396 11421
0 11423 7 1 2 11378 11422
0 11424 7 1 2 11357 11423
0 11425 5 1 1 11424
0 11426 7 1 2 54763 11425
0 11427 5 1 1 11426
0 11428 7 3 2 42005 47245
0 11429 7 1 2 59193 63889
0 11430 5 2 1 11429
0 11431 7 6 2 47531 47638
0 11432 7 2 2 46652 63894
0 11433 7 1 2 58183 58598
0 11434 7 1 2 63900 11433
0 11435 5 1 1 11434
0 11436 7 1 2 63892 11435
0 11437 5 1 1 11436
0 11438 7 1 2 42753 11437
0 11439 5 1 1 11438
0 11440 7 3 2 54030 59911
0 11441 5 1 1 63902
0 11442 7 1 2 43875 63903
0 11443 5 1 1 11442
0 11444 7 1 2 11439 11443
0 11445 5 1 1 11444
0 11446 7 1 2 45221 11445
0 11447 5 1 1 11446
0 11448 7 1 2 59781 63590
0 11449 5 2 1 11448
0 11450 7 4 2 48591 54231
0 11451 5 2 1 63907
0 11452 7 1 2 51415 63911
0 11453 5 7 1 11452
0 11454 7 1 2 59837 63913
0 11455 5 1 1 11454
0 11456 7 1 2 63905 11455
0 11457 5 1 1 11456
0 11458 7 1 2 47246 11457
0 11459 5 1 1 11458
0 11460 7 1 2 59838 63259
0 11461 5 2 1 11460
0 11462 7 1 2 53967 58184
0 11463 7 1 2 63087 11462
0 11464 5 1 1 11463
0 11465 7 1 2 63920 11464
0 11466 5 1 1 11465
0 11467 7 1 2 46208 11466
0 11468 5 1 1 11467
0 11469 7 1 2 11459 11468
0 11470 5 1 1 11469
0 11471 7 1 2 49968 11470
0 11472 5 1 1 11471
0 11473 7 2 2 46831 43876
0 11474 7 3 2 61230 63922
0 11475 7 2 2 50550 60226
0 11476 7 1 2 63924 63927
0 11477 5 1 1 11476
0 11478 7 1 2 11477 63893
0 11479 5 1 1 11478
0 11480 7 1 2 42754 11479
0 11481 5 1 1 11480
0 11482 7 1 2 43877 53042
0 11483 5 2 1 11482
0 11484 7 1 2 61965 63929
0 11485 5 1 1 11484
0 11486 7 1 2 59839 11485
0 11487 5 1 1 11486
0 11488 7 1 2 11481 11487
0 11489 5 1 1 11488
0 11490 7 1 2 50065 11489
0 11491 5 1 1 11490
0 11492 7 1 2 11472 11491
0 11493 7 1 2 11447 11492
0 11494 5 1 1 11493
0 11495 7 1 2 61048 11494
0 11496 5 1 1 11495
0 11497 7 1 2 11427 11496
0 11498 5 1 1 11497
0 11499 7 1 2 62683 11498
0 11500 5 1 1 11499
0 11501 7 21 2 42755 46468
0 11502 7 1 2 51914 63931
0 11503 5 1 1 11502
0 11504 7 1 2 45432 62896
0 11505 5 1 1 11504
0 11506 7 1 2 11503 11505
0 11507 5 1 1 11506
0 11508 7 1 2 62490 11507
0 11509 5 1 1 11508
0 11510 7 7 2 46469 47750
0 11511 7 3 2 45557 63952
0 11512 7 2 2 56952 60913
0 11513 5 2 1 63962
0 11514 7 1 2 63959 63963
0 11515 5 1 1 11514
0 11516 7 1 2 11509 11515
0 11517 5 1 1 11516
0 11518 7 1 2 62913 11517
0 11519 5 1 1 11518
0 11520 7 3 2 43527 47751
0 11521 7 4 2 63278 63966
0 11522 7 1 2 54986 56953
0 11523 7 1 2 63865 11522
0 11524 7 1 2 63969 11523
0 11525 5 1 1 11524
0 11526 7 1 2 11519 11525
0 11527 5 1 1 11526
0 11528 7 1 2 47532 11527
0 11529 5 1 1 11528
0 11530 7 2 2 46470 62729
0 11531 5 1 1 63973
0 11532 7 1 2 63974 63845
0 11533 5 1 1 11532
0 11534 7 1 2 11529 11533
0 11535 5 1 1 11534
0 11536 7 1 2 46653 11535
0 11537 5 1 1 11536
0 11538 7 5 2 45433 49969
0 11539 5 1 1 63975
0 11540 7 1 2 5807 11539
0 11541 5 2 1 11540
0 11542 7 1 2 59264 63980
0 11543 5 1 1 11542
0 11544 7 1 2 42756 62761
0 11545 5 1 1 11544
0 11546 7 1 2 11543 11545
0 11547 5 1 1 11546
0 11548 7 1 2 62914 11547
0 11549 5 1 1 11548
0 11550 7 3 2 45711 62706
0 11551 7 1 2 60175 63319
0 11552 7 1 2 63982 11551
0 11553 5 2 1 11552
0 11554 7 1 2 11549 63985
0 11555 5 1 1 11554
0 11556 7 1 2 46471 11555
0 11557 5 1 1 11556
0 11558 7 1 2 62915 63932
0 11559 5 1 1 11558
0 11560 7 1 2 62742 11559
0 11561 5 1 1 11560
0 11562 7 1 2 59265 11561
0 11563 5 1 1 11562
0 11564 7 2 2 63933 63765
0 11565 7 1 2 60227 63063
0 11566 7 1 2 63987 11565
0 11567 5 1 1 11566
0 11568 7 1 2 62743 11567
0 11569 5 1 1 11568
0 11570 7 1 2 51915 11569
0 11571 5 1 1 11570
0 11572 7 1 2 11563 11571
0 11573 5 1 1 11572
0 11574 7 1 2 46654 11573
0 11575 5 1 1 11574
0 11576 7 1 2 58684 9984
0 11577 5 1 1 11576
0 11578 7 1 2 62730 11577
0 11579 5 1 1 11578
0 11580 7 1 2 11575 11579
0 11581 7 1 2 11557 11580
0 11582 5 1 1 11581
0 11583 7 1 2 62491 11582
0 11584 5 1 1 11583
0 11585 7 19 2 45712 42264
0 11586 7 4 2 58062 63989
0 11587 7 1 2 56954 61231
0 11588 7 1 2 63970 11587
0 11589 7 1 2 64008 11588
0 11590 5 1 1 11589
0 11591 7 1 2 11584 11590
0 11592 7 1 2 11537 11591
0 11593 5 1 1 11592
0 11594 7 1 2 50551 11593
0 11595 5 1 1 11594
0 11596 7 4 2 46960 47410
0 11597 7 2 2 44193 64012
0 11598 7 1 2 64016 63771
0 11599 5 1 1 11598
0 11600 7 1 2 11531 11599
0 11601 5 1 1 11600
0 11602 7 1 2 11601 63673
0 11603 5 1 1 11602
0 11604 7 1 2 50174 60804
0 11605 7 1 2 63777 11604
0 11606 5 1 1 11605
0 11607 7 1 2 11603 11606
0 11608 5 1 1 11607
0 11609 7 1 2 43269 11608
0 11610 5 1 1 11609
0 11611 7 14 2 45794 46655
0 11612 7 1 2 48592 57273
0 11613 7 1 2 64018 11612
0 11614 7 1 2 63175 11613
0 11615 5 1 1 11614
0 11616 7 1 2 62744 11615
0 11617 5 1 1 11616
0 11618 7 1 2 63543 11617
0 11619 5 1 1 11618
0 11620 7 3 2 47533 63279
0 11621 7 4 2 45558 63990
0 11622 7 1 2 64032 64035
0 11623 7 2 2 46656 55753
0 11624 7 2 2 47752 56562
0 11625 7 1 2 64039 64041
0 11626 7 1 2 11622 11625
0 11627 5 1 1 11626
0 11628 7 1 2 11619 11627
0 11629 7 1 2 11610 11628
0 11630 5 1 1 11629
0 11631 7 1 2 45434 11630
0 11632 5 1 1 11631
0 11633 7 1 2 57608 63727
0 11634 7 1 2 63108 11633
0 11635 5 1 1 11634
0 11636 7 1 2 63986 11635
0 11637 5 1 1 11636
0 11638 7 1 2 50066 11637
0 11639 5 1 1 11638
0 11640 7 3 2 58703 59478
0 11641 7 8 2 45795 43270
0 11642 7 1 2 64013 64046
0 11643 7 1 2 64043 11642
0 11644 5 1 1 11643
0 11645 7 1 2 62745 11644
0 11646 5 1 1 11645
0 11647 7 1 2 51916 11646
0 11648 5 1 1 11647
0 11649 7 3 2 45796 59266
0 11650 7 1 2 55794 59947
0 11651 7 1 2 64017 11650
0 11652 7 1 2 64054 11651
0 11653 5 1 1 11652
0 11654 7 1 2 11648 11653
0 11655 5 1 1 11654
0 11656 7 1 2 45222 11655
0 11657 5 1 1 11656
0 11658 7 1 2 11639 11657
0 11659 5 1 1 11658
0 11660 7 1 2 62492 11659
0 11661 5 1 1 11660
0 11662 7 1 2 51500 62916
0 11663 5 1 1 11662
0 11664 7 1 2 62746 11663
0 11665 5 3 1 11664
0 11666 7 1 2 61766 63651
0 11667 5 2 1 11666
0 11668 7 1 2 61210 62843
0 11669 7 1 2 63700 11668
0 11670 5 1 1 11669
0 11671 7 1 2 64060 11670
0 11672 5 2 1 11671
0 11673 7 1 2 64057 64062
0 11674 5 1 1 11673
0 11675 7 1 2 43057 63530
0 11676 5 1 1 11675
0 11677 7 1 2 60176 63441
0 11678 7 1 2 49595 50280
0 11679 5 4 1 11678
0 11680 7 4 2 47753 61263
0 11681 7 1 2 64064 64068
0 11682 7 1 2 11677 11681
0 11683 7 1 2 11676 11682
0 11684 5 1 1 11683
0 11685 7 1 2 11674 11684
0 11686 7 1 2 11661 11685
0 11687 7 1 2 11632 11686
0 11688 5 1 1 11687
0 11689 7 1 2 46209 11688
0 11690 5 1 1 11689
0 11691 7 1 2 11595 11690
0 11692 5 1 1 11691
0 11693 7 1 2 43878 11692
0 11694 5 1 1 11693
0 11695 7 1 2 11500 11694
0 11696 7 1 2 11339 11695
0 11697 5 1 1 11696
0 11698 7 1 2 61375 11697
0 11699 5 1 1 11698
0 11700 7 11 2 47639 47754
0 11701 7 1 2 55322 64072
0 11702 7 2 2 50671 60376
0 11703 7 1 2 60282 64083
0 11704 7 2 2 11701 11703
0 11705 7 1 2 55399 61264
0 11706 7 1 2 64085 11705
0 11707 5 1 1 11706
0 11708 7 3 2 51560 57435
0 11709 7 6 2 47247 44318
0 11710 7 1 2 57961 64090
0 11711 7 1 2 64087 11710
0 11712 7 1 2 61670 11711
0 11713 5 1 1 11712
0 11714 7 1 2 11707 11713
0 11715 5 1 1 11714
0 11716 7 1 2 62684 11715
0 11717 5 1 1 11716
0 11718 7 1 2 46961 55795
0 11719 7 11 2 45797 42510
0 11720 7 1 2 61018 64096
0 11721 7 1 2 11718 11720
0 11722 7 1 2 64086 11721
0 11723 5 1 1 11722
0 11724 7 18 2 42265 46210
0 11725 7 1 2 50708 64091
0 11726 7 1 2 64107 11725
0 11727 7 3 2 56424 59014
0 11728 5 2 1 64125
0 11729 7 1 2 62796 63427
0 11730 7 1 2 64126 11729
0 11731 7 1 2 11726 11730
0 11732 5 1 1 11731
0 11733 7 1 2 11723 11732
0 11734 7 1 2 11717 11733
0 11735 5 1 1 11734
0 11736 7 4 2 49750 50607
0 11737 7 1 2 50189 64130
0 11738 7 1 2 11735 11737
0 11739 5 1 1 11738
0 11740 7 1 2 11699 11739
0 11741 7 1 2 10829 11740
0 11742 7 1 2 10574 11741
0 11743 7 1 2 10214 11742
0 11744 5 1 1 11743
0 11745 7 1 2 45057 11744
0 11746 5 1 1 11745
0 11747 7 1 2 57098 59503
0 11748 5 2 1 11747
0 11749 7 1 2 54532 62650
0 11750 7 1 2 64134 11749
0 11751 5 1 1 11750
0 11752 7 2 2 56821 56889
0 11753 7 1 2 57013 62563
0 11754 7 1 2 64136 11753
0 11755 5 1 1 11754
0 11756 7 1 2 11751 11755
0 11757 5 1 1 11756
0 11758 7 1 2 46472 11757
0 11759 5 1 1 11758
0 11760 7 1 2 46657 57652
0 11761 5 3 1 11760
0 11762 7 1 2 57326 64138
0 11763 5 4 1 11762
0 11764 7 2 2 52038 61395
0 11765 5 1 1 64145
0 11766 7 1 2 64141 64146
0 11767 5 1 1 11766
0 11768 7 1 2 59435 62630
0 11769 5 1 1 11768
0 11770 7 1 2 11767 11769
0 11771 5 1 1 11770
0 11772 7 1 2 45223 11771
0 11773 5 1 1 11772
0 11774 7 2 2 50608 60283
0 11775 5 2 1 64147
0 11776 7 1 2 51752 61726
0 11777 7 1 2 64148 11776
0 11778 5 1 1 11777
0 11779 7 1 2 11773 11778
0 11780 5 1 1 11779
0 11781 7 1 2 43058 11780
0 11782 5 1 1 11781
0 11783 7 1 2 51365 51425
0 11784 7 1 2 61702 11783
0 11785 5 1 1 11784
0 11786 7 2 2 58415 63453
0 11787 7 1 2 51051 63462
0 11788 7 1 2 64151 11787
0 11789 5 1 1 11788
0 11790 7 1 2 11785 11789
0 11791 5 1 1 11790
0 11792 7 1 2 60284 11791
0 11793 5 1 1 11792
0 11794 7 1 2 11782 11793
0 11795 7 1 2 11759 11794
0 11796 5 1 1 11795
0 11797 7 1 2 60528 11796
0 11798 5 1 1 11797
0 11799 7 2 2 52766 61515
0 11800 5 1 1 64153
0 11801 7 1 2 54533 60377
0 11802 7 1 2 52665 11801
0 11803 5 1 1 11802
0 11804 7 1 2 11800 11803
0 11805 5 1 1 11804
0 11806 7 1 2 45224 11805
0 11807 5 1 1 11806
0 11808 7 1 2 55987 62010
0 11809 5 1 1 11808
0 11810 7 1 2 11807 11809
0 11811 5 1 1 11810
0 11812 7 1 2 46658 11811
0 11813 5 1 1 11812
0 11814 7 2 2 54031 57558
0 11815 5 2 1 64155
0 11816 7 1 2 47248 64156
0 11817 5 1 1 11816
0 11818 7 1 2 43879 8658
0 11819 5 1 1 11818
0 11820 7 1 2 49970 11819
0 11821 7 1 2 11817 11820
0 11822 5 1 1 11821
0 11823 7 1 2 62064 11822
0 11824 5 1 1 11823
0 11825 7 1 2 43716 11824
0 11826 5 1 1 11825
0 11827 7 1 2 62383 11826
0 11828 5 1 1 11827
0 11829 7 1 2 60378 11828
0 11830 5 1 1 11829
0 11831 7 1 2 11813 11830
0 11832 5 1 1 11831
0 11833 7 1 2 48799 11832
0 11834 5 1 1 11833
0 11835 7 1 2 50838 60285
0 11836 5 1 1 11835
0 11837 7 2 2 43880 53358
0 11838 5 1 1 64159
0 11839 7 1 2 52056 63677
0 11840 5 1 1 11839
0 11841 7 1 2 11838 11840
0 11842 5 1 1 11841
0 11843 7 1 2 45435 11842
0 11844 5 1 1 11843
0 11845 7 1 2 11836 11844
0 11846 5 1 1 11845
0 11847 7 1 2 48593 11846
0 11848 5 1 1 11847
0 11849 7 2 2 45225 51335
0 11850 5 1 1 64161
0 11851 7 1 2 54341 11850
0 11852 5 1 1 11851
0 11853 7 1 2 57003 11852
0 11854 5 1 1 11853
0 11855 7 1 2 11848 11854
0 11856 5 1 1 11855
0 11857 7 1 2 44047 11856
0 11858 5 1 1 11857
0 11859 7 1 2 58555 59650
0 11860 5 1 1 11859
0 11861 7 1 2 43881 11860
0 11862 5 1 1 11861
0 11863 7 1 2 47249 49627
0 11864 5 2 1 11863
0 11865 7 1 2 43059 64163
0 11866 7 1 2 57477 11865
0 11867 5 1 1 11866
0 11868 7 1 2 11862 11867
0 11869 5 1 1 11868
0 11870 7 1 2 42757 11869
0 11871 5 1 1 11870
0 11872 7 1 2 11858 11871
0 11873 5 1 1 11872
0 11874 7 1 2 61219 11873
0 11875 5 1 1 11874
0 11876 7 1 2 11834 11875
0 11877 5 1 1 11876
0 11878 7 1 2 59381 11877
0 11879 5 1 1 11878
0 11880 7 1 2 11798 11879
0 11881 5 1 1 11880
0 11882 7 1 2 46005 11881
0 11883 5 1 1 11882
0 11884 7 1 2 42511 2771
0 11885 5 1 1 11884
0 11886 7 1 2 53185 61998
0 11887 5 1 1 11886
0 11888 7 1 2 11885 11887
0 11889 5 1 1 11888
0 11890 7 1 2 60379 11889
0 11891 5 1 1 11890
0 11892 7 3 2 59220 61006
0 11893 7 1 2 52767 64165
0 11894 5 1 1 11893
0 11895 7 1 2 11891 11894
0 11896 5 1 1 11895
0 11897 7 1 2 59382 11896
0 11898 5 1 1 11897
0 11899 7 2 2 45559 55183
0 11900 7 1 2 62805 64168
0 11901 7 1 2 62020 11900
0 11902 5 1 1 11901
0 11903 7 1 2 11898 11902
0 11904 5 1 1 11903
0 11905 7 1 2 55571 11904
0 11906 5 1 1 11905
0 11907 7 1 2 62662 64169
0 11908 7 1 2 62075 11907
0 11909 5 1 1 11908
0 11910 7 1 2 47250 53161
0 11911 7 1 2 59383 11910
0 11912 5 1 1 11911
0 11913 7 1 2 62055 62586
0 11914 5 1 1 11913
0 11915 7 1 2 11912 11914
0 11916 5 1 1 11915
0 11917 7 1 2 60380 62241
0 11918 7 1 2 11916 11917
0 11919 5 1 1 11918
0 11920 7 1 2 11909 11919
0 11921 5 1 1 11920
0 11922 7 1 2 62271 11921
0 11923 5 1 1 11922
0 11924 7 1 2 60907 63588
0 11925 5 1 1 11924
0 11926 7 2 2 59361 61580
0 11927 7 1 2 62178 64170
0 11928 5 1 1 11927
0 11929 7 1 2 60953 61237
0 11930 5 1 1 11929
0 11931 7 2 2 44438 45226
0 11932 7 2 2 47640 64172
0 11933 7 2 2 45560 56210
0 11934 7 1 2 64174 64176
0 11935 5 1 1 11934
0 11936 7 1 2 11930 11935
0 11937 7 1 2 11928 11936
0 11938 5 1 1 11937
0 11939 7 1 2 47534 11938
0 11940 5 1 1 11939
0 11941 7 1 2 11925 11940
0 11942 5 1 1 11941
0 11943 7 1 2 46659 11942
0 11944 5 1 1 11943
0 11945 7 2 2 49277 61080
0 11946 7 2 2 56185 60926
0 11947 7 1 2 64178 64180
0 11948 5 1 1 11947
0 11949 7 1 2 60908 64171
0 11950 5 1 1 11949
0 11951 7 2 2 49207 59150
0 11952 7 1 2 64179 64182
0 11953 5 1 1 11952
0 11954 7 1 2 11950 11953
0 11955 5 1 1 11954
0 11956 7 1 2 43271 11955
0 11957 5 1 1 11956
0 11958 7 1 2 11948 11957
0 11959 7 1 2 11944 11958
0 11960 5 1 1 11959
0 11961 7 1 2 47251 11960
0 11962 5 1 1 11961
0 11963 7 2 2 45561 54325
0 11964 7 1 2 64184 64175
0 11965 5 1 1 11964
0 11966 7 1 2 55303 59384
0 11967 5 1 1 11966
0 11968 7 1 2 11965 11967
0 11969 5 1 1 11968
0 11970 7 1 2 46660 11969
0 11971 5 1 1 11970
0 11972 7 2 2 42006 60598
0 11973 7 1 2 57271 64186
0 11974 5 1 1 11973
0 11975 7 1 2 11971 11974
0 11976 5 1 1 11975
0 11977 7 1 2 61524 11976
0 11978 5 1 1 11977
0 11979 7 1 2 43717 11978
0 11980 7 1 2 11962 11979
0 11981 5 1 1 11980
0 11982 7 1 2 49208 62060
0 11983 5 1 1 11982
0 11984 7 2 2 45436 53000
0 11985 7 1 2 50759 64188
0 11986 5 1 1 11985
0 11987 7 1 2 11983 11986
0 11988 5 1 1 11987
0 11989 7 1 2 48594 11988
0 11990 5 1 1 11989
0 11991 7 1 2 53380 54032
0 11992 5 1 1 11991
0 11993 7 1 2 49034 52001
0 11994 7 1 2 11992 11993
0 11995 5 1 1 11994
0 11996 7 1 2 57183 60712
0 11997 5 1 1 11996
0 11998 7 1 2 49691 55160
0 11999 5 1 1 11998
0 12000 7 1 2 11997 11999
0 12001 7 1 2 11995 12000
0 12002 5 1 1 12001
0 12003 7 1 2 43272 12002
0 12004 5 1 1 12003
0 12005 7 1 2 51793 61999
0 12006 5 1 1 12005
0 12007 7 1 2 54014 56787
0 12008 5 1 1 12007
0 12009 7 1 2 12006 12008
0 12010 7 1 2 12004 12009
0 12011 7 1 2 11990 12010
0 12012 5 1 1 12011
0 12013 7 1 2 59385 12012
0 12014 5 1 1 12013
0 12015 7 1 2 46473 64135
0 12016 5 1 1 12015
0 12017 7 1 2 51972 53322
0 12018 7 1 2 12016 12017
0 12019 5 1 1 12018
0 12020 7 1 2 51515 52094
0 12021 5 1 1 12020
0 12022 7 1 2 50609 60701
0 12023 5 1 1 12022
0 12024 7 1 2 52002 12023
0 12025 7 1 2 12021 12024
0 12026 5 1 1 12025
0 12027 7 1 2 52057 60529
0 12028 7 1 2 12026 12027
0 12029 7 1 2 12019 12028
0 12030 5 1 1 12029
0 12031 7 1 2 47092 12030
0 12032 7 1 2 12014 12031
0 12033 5 1 1 12032
0 12034 7 1 2 48094 12033
0 12035 7 1 2 11981 12034
0 12036 5 1 1 12035
0 12037 7 2 2 42007 44750
0 12038 7 9 2 47755 48595
0 12039 7 1 2 49512 64192
0 12040 7 1 2 64190 12039
0 12041 7 2 2 42758 62363
0 12042 7 2 2 54160 59600
0 12043 7 1 2 64201 64203
0 12044 7 1 2 12040 12043
0 12045 5 1 1 12044
0 12046 7 1 2 12036 12045
0 12047 5 1 1 12046
0 12048 7 1 2 62024 12047
0 12049 5 1 1 12048
0 12050 7 1 2 11923 12049
0 12051 7 1 2 11906 12050
0 12052 7 1 2 11883 12051
0 12053 5 1 1 12052
0 12054 7 1 2 51917 12053
0 12055 5 1 1 12054
0 12056 7 1 2 59386 9467
0 12057 5 1 1 12056
0 12058 7 1 2 56655 62457
0 12059 5 1 1 12058
0 12060 7 1 2 62436 12059
0 12061 5 1 1 12060
0 12062 7 1 2 59387 12061
0 12063 5 1 1 12062
0 12064 7 2 2 58441 62195
0 12065 5 1 1 64205
0 12066 7 1 2 9108 12065
0 12067 5 1 1 12066
0 12068 7 1 2 43718 12067
0 12069 5 1 1 12068
0 12070 7 1 2 4115 59709
0 12071 5 7 1 12070
0 12072 7 1 2 53999 64207
0 12073 5 1 1 12072
0 12074 7 1 2 12069 12073
0 12075 5 1 1 12074
0 12076 7 1 2 60530 12075
0 12077 5 1 1 12076
0 12078 7 1 2 12063 12077
0 12079 5 1 1 12078
0 12080 7 1 2 42512 12079
0 12081 5 1 1 12080
0 12082 7 1 2 52249 62385
0 12083 5 2 1 12082
0 12084 7 1 2 60531 64214
0 12085 5 1 1 12084
0 12086 7 2 2 50839 61644
0 12087 5 1 1 64216
0 12088 7 1 2 48800 64217
0 12089 5 1 1 12088
0 12090 7 1 2 12085 12089
0 12091 5 1 1 12090
0 12092 7 1 2 44048 12091
0 12093 5 1 1 12092
0 12094 7 1 2 59151 59663
0 12095 5 1 1 12094
0 12096 7 1 2 8076 12095
0 12097 5 1 1 12096
0 12098 7 1 2 52222 12097
0 12099 5 1 1 12098
0 12100 7 1 2 12093 12099
0 12101 5 1 1 12100
0 12102 7 1 2 46006 54161
0 12103 7 1 2 12101 12102
0 12104 5 1 1 12103
0 12105 7 1 2 12081 12104
0 12106 5 1 1 12105
0 12107 7 1 2 60381 12106
0 12108 5 1 1 12107
0 12109 7 1 2 55572 59388
0 12110 5 2 1 12109
0 12111 7 1 2 57108 60532
0 12112 5 1 1 12111
0 12113 7 1 2 64218 12112
0 12114 5 1 1 12113
0 12115 7 1 2 45437 12114
0 12116 5 1 1 12115
0 12117 7 1 2 52804 59389
0 12118 5 1 1 12117
0 12119 7 1 2 12116 12118
0 12120 5 1 1 12119
0 12121 7 1 2 52239 12120
0 12122 5 1 1 12121
0 12123 7 2 2 61232 62196
0 12124 7 1 2 58870 60927
0 12125 7 1 2 64220 12124
0 12126 5 1 1 12125
0 12127 7 1 2 12122 12126
0 12128 5 1 1 12127
0 12129 7 1 2 61191 12128
0 12130 5 1 1 12129
0 12131 7 1 2 12108 12130
0 12132 5 1 1 12131
0 12133 7 1 2 46211 12132
0 12134 5 1 1 12133
0 12135 7 1 2 60533 9256
0 12136 5 1 1 12135
0 12137 7 2 2 47093 52114
0 12138 5 1 1 64222
0 12139 7 1 2 55984 12138
0 12140 5 1 1 12139
0 12141 7 2 2 42513 59390
0 12142 7 1 2 12140 64224
0 12143 5 1 1 12142
0 12144 7 1 2 53186 61645
0 12145 7 1 2 52115 12144
0 12146 5 1 1 12145
0 12147 7 1 2 12143 12146
0 12148 5 1 1 12147
0 12149 7 1 2 62230 12148
0 12150 5 1 1 12149
0 12151 7 5 2 52895 62587
0 12152 5 1 1 64226
0 12153 7 1 2 56832 61881
0 12154 7 1 2 64227 12153
0 12155 5 1 1 12154
0 12156 7 1 2 12150 12155
0 12157 5 1 1 12156
0 12158 7 1 2 50067 12157
0 12159 5 1 1 12158
0 12160 7 1 2 12136 12159
0 12161 7 1 2 12134 12160
0 12162 7 1 2 12057 12161
0 12163 5 1 1 12162
0 12164 7 1 2 59267 12163
0 12165 5 1 1 12164
0 12166 7 1 2 59322 62759
0 12167 5 5 1 12166
0 12168 7 1 2 62605 64231
0 12169 5 1 1 12168
0 12170 7 6 2 44194 44559
0 12171 7 2 2 61850 64236
0 12172 5 1 1 64242
0 12173 7 2 2 47884 51753
0 12174 7 1 2 45713 64244
0 12175 5 1 1 12174
0 12176 7 1 2 12172 12175
0 12177 5 1 1 12176
0 12178 7 1 2 59062 12177
0 12179 5 1 1 12178
0 12180 7 1 2 53851 54162
0 12181 7 1 2 62875 12180
0 12182 5 1 1 12181
0 12183 7 1 2 12179 12182
0 12184 5 1 1 12183
0 12185 7 1 2 60534 12184
0 12186 5 1 1 12185
0 12187 7 4 2 47885 61633
0 12188 5 1 1 64246
0 12189 7 1 2 62210 64247
0 12190 5 1 1 12189
0 12191 7 1 2 63145 12190
0 12192 5 1 1 12191
0 12193 7 2 2 60636 63467
0 12194 7 1 2 62109 64250
0 12195 7 1 2 12192 12194
0 12196 5 1 1 12195
0 12197 7 1 2 12186 12196
0 12198 5 1 1 12197
0 12199 7 1 2 60382 12198
0 12200 5 1 1 12199
0 12201 7 1 2 54338 60535
0 12202 5 1 1 12201
0 12203 7 1 2 64219 12202
0 12204 5 1 1 12203
0 12205 7 1 2 45438 12204
0 12206 5 1 1 12205
0 12207 7 1 2 62197 63635
0 12208 5 1 1 12207
0 12209 7 1 2 12206 12208
0 12210 5 1 1 12209
0 12211 7 1 2 46212 12210
0 12212 5 1 1 12211
0 12213 7 2 2 60637 61061
0 12214 7 1 2 63890 64252
0 12215 5 1 1 12214
0 12216 7 1 2 12212 12215
0 12217 5 1 1 12216
0 12218 7 1 2 59268 12217
0 12219 5 1 1 12218
0 12220 7 2 2 57347 59015
0 12221 7 2 2 57866 60638
0 12222 7 1 2 64254 64256
0 12223 5 1 1 12222
0 12224 7 1 2 12219 12223
0 12225 5 1 1 12224
0 12226 7 1 2 61192 12225
0 12227 5 1 1 12226
0 12228 7 1 2 12200 12227
0 12229 5 1 1 12228
0 12230 7 1 2 45227 12229
0 12231 5 1 1 12230
0 12232 7 1 2 61623 62844
0 12233 5 1 1 12232
0 12234 7 1 2 11050 12233
0 12235 5 1 1 12234
0 12236 7 1 2 43273 12235
0 12237 5 1 1 12236
0 12238 7 5 2 46661 51918
0 12239 7 1 2 49209 61646
0 12240 7 1 2 64258 12239
0 12241 5 1 1 12240
0 12242 7 1 2 12237 12241
0 12243 5 1 1 12242
0 12244 7 1 2 61376 12243
0 12245 5 1 1 12244
0 12246 7 4 2 42162 64237
0 12247 5 1 1 64263
0 12248 7 1 2 61193 64264
0 12249 5 1 1 12248
0 12250 7 2 2 50350 56017
0 12251 7 1 2 45714 51371
0 12252 7 1 2 64267 12251
0 12253 5 1 1 12252
0 12254 7 1 2 12249 12253
0 12255 5 1 1 12254
0 12256 7 2 2 60639 12255
0 12257 7 1 2 42008 64269
0 12258 5 1 1 12257
0 12259 7 1 2 12245 12258
0 12260 5 1 1 12259
0 12261 7 1 2 52039 12260
0 12262 5 1 1 12261
0 12263 7 1 2 12231 12262
0 12264 5 1 1 12263
0 12265 7 1 2 50996 12264
0 12266 5 1 1 12265
0 12267 7 1 2 12169 12266
0 12268 7 1 2 12165 12267
0 12269 7 1 2 12055 12268
0 12270 5 1 1 12269
0 12271 7 1 2 48406 12270
0 12272 5 1 1 12271
0 12273 7 1 2 55550 63632
0 12274 5 1 1 12273
0 12275 7 1 2 62588 62817
0 12276 5 1 1 12275
0 12277 7 1 2 10967 12276
0 12278 5 1 1 12277
0 12279 7 1 2 45228 12278
0 12280 7 1 2 12274 12279
0 12281 5 1 1 12280
0 12282 7 1 2 48596 63149
0 12283 5 1 1 12282
0 12284 7 1 2 63146 12283
0 12285 5 1 1 12284
0 12286 7 1 2 59391 12285
0 12287 5 1 1 12286
0 12288 7 1 2 12281 12287
0 12289 5 1 1 12288
0 12290 7 1 2 44049 12289
0 12291 5 1 1 12290
0 12292 7 1 2 51541 59115
0 12293 5 2 1 12292
0 12294 7 2 2 44560 60640
0 12295 7 4 2 56232 64273
0 12296 7 1 2 64271 64275
0 12297 5 1 1 12296
0 12298 7 1 2 12291 12297
0 12299 5 1 1 12298
0 12300 7 1 2 43060 12299
0 12301 5 1 1 12300
0 12302 7 1 2 44050 64276
0 12303 7 1 2 53510 12302
0 12304 5 1 1 12303
0 12305 7 1 2 12301 12304
0 12306 5 1 1 12305
0 12307 7 1 2 51973 53258
0 12308 7 1 2 12306 12307
0 12309 5 1 1 12308
0 12310 7 1 2 60872 62768
0 12311 5 1 1 12310
0 12312 7 1 2 42163 61846
0 12313 5 1 1 12312
0 12314 7 1 2 12311 12313
0 12315 5 1 1 12314
0 12316 7 1 2 57532 58493
0 12317 7 1 2 64251 12316
0 12318 7 1 2 12315 12317
0 12319 5 1 1 12318
0 12320 7 1 2 12309 12319
0 12321 5 1 1 12320
0 12322 7 1 2 60383 12321
0 12323 5 1 1 12322
0 12324 7 1 2 55339 59773
0 12325 7 2 2 52978 57247
0 12326 7 1 2 62797 64279
0 12327 7 1 2 12324 12326
0 12328 7 1 2 63575 12327
0 12329 5 1 1 12328
0 12330 7 1 2 12323 12329
0 12331 7 1 2 12272 12330
0 12332 5 1 1 12331
0 12333 7 1 2 62998 12332
0 12334 5 1 1 12333
0 12335 7 1 2 52250 52768
0 12336 5 1 1 12335
0 12337 7 1 2 55340 57371
0 12338 5 1 1 12337
0 12339 7 1 2 12336 12338
0 12340 5 1 1 12339
0 12341 7 1 2 61194 12340
0 12342 5 1 1 12341
0 12343 7 1 2 61338 62431
0 12344 5 1 1 12343
0 12345 7 3 2 45439 60286
0 12346 5 1 1 64281
0 12347 7 1 2 47411 64282
0 12348 5 1 1 12347
0 12349 7 1 2 58474 12348
0 12350 5 1 1 12349
0 12351 7 1 2 45229 12350
0 12352 5 1 1 12351
0 12353 7 1 2 42514 57084
0 12354 5 1 1 12353
0 12355 7 1 2 55350 12354
0 12356 5 1 1 12355
0 12357 7 1 2 49971 12356
0 12358 7 1 2 12352 12357
0 12359 5 1 1 12358
0 12360 7 1 2 50610 58473
0 12361 5 3 1 12360
0 12362 7 1 2 50068 64284
0 12363 5 1 1 12362
0 12364 7 1 2 43061 12363
0 12365 7 1 2 12359 12364
0 12366 5 1 1 12365
0 12367 7 1 2 56894 57122
0 12368 5 1 1 12367
0 12369 7 1 2 42759 12368
0 12370 5 1 1 12369
0 12371 7 1 2 49972 54232
0 12372 5 4 1 12371
0 12373 7 1 2 56895 64287
0 12374 5 1 1 12373
0 12375 7 1 2 43882 12374
0 12376 5 1 1 12375
0 12377 7 1 2 12370 12376
0 12378 5 1 1 12377
0 12379 7 1 2 48597 12378
0 12380 5 1 1 12379
0 12381 7 1 2 42760 62448
0 12382 5 1 1 12381
0 12383 7 1 2 12380 12382
0 12384 5 2 1 12383
0 12385 7 1 2 46007 64291
0 12386 5 1 1 12385
0 12387 7 1 2 46213 53944
0 12388 5 2 1 12387
0 12389 7 1 2 53327 56850
0 12390 5 1 1 12389
0 12391 7 1 2 64293 12390
0 12392 5 1 1 12391
0 12393 7 1 2 42515 12392
0 12394 5 1 1 12393
0 12395 7 1 2 12386 12394
0 12396 7 1 2 12366 12395
0 12397 5 1 1 12396
0 12398 7 1 2 48095 12397
0 12399 5 1 1 12398
0 12400 7 1 2 12344 12399
0 12401 5 1 1 12400
0 12402 7 1 2 43719 12401
0 12403 5 1 1 12402
0 12404 7 1 2 50069 53374
0 12405 5 1 1 12404
0 12406 7 1 2 53491 12405
0 12407 5 1 1 12406
0 12408 7 1 2 53196 12407
0 12409 5 1 1 12408
0 12410 7 1 2 42516 59185
0 12411 5 1 1 12410
0 12412 7 1 2 50683 52956
0 12413 7 1 2 52223 12412
0 12414 5 1 1 12413
0 12415 7 1 2 12411 12414
0 12416 5 1 1 12415
0 12417 7 1 2 47094 12416
0 12418 5 1 1 12417
0 12419 7 1 2 58438 61110
0 12420 5 1 1 12419
0 12421 7 1 2 12418 12420
0 12422 5 1 1 12421
0 12423 7 1 2 42761 12422
0 12424 5 1 1 12423
0 12425 7 1 2 12409 12424
0 12426 5 1 1 12425
0 12427 7 1 2 43062 12426
0 12428 5 1 1 12427
0 12429 7 1 2 53197 64292
0 12430 5 1 1 12429
0 12431 7 1 2 12428 12430
0 12432 5 1 1 12431
0 12433 7 1 2 48096 12432
0 12434 5 1 1 12433
0 12435 7 1 2 12403 12434
0 12436 5 1 1 12435
0 12437 7 1 2 44636 12436
0 12438 5 1 1 12437
0 12439 7 1 2 12342 12438
0 12440 5 1 1 12439
0 12441 7 1 2 62731 12440
0 12442 5 1 1 12441
0 12443 7 3 2 55184 55796
0 12444 7 14 2 45798 46474
0 12445 7 1 2 63661 64298
0 12446 7 2 2 64295 12445
0 12447 7 5 2 46962 44751
0 12448 7 1 2 61430 64314
0 12449 7 1 2 64312 12448
0 12450 5 1 1 12449
0 12451 7 1 2 43453 57939
0 12452 7 1 2 63210 12451
0 12453 7 2 2 42266 54214
0 12454 7 1 2 63256 64319
0 12455 7 1 2 12452 12454
0 12456 5 1 1 12455
0 12457 7 1 2 12450 12456
0 12458 5 1 1 12457
0 12459 7 1 2 47095 12458
0 12460 5 1 1 12459
0 12461 7 1 2 52040 63448
0 12462 5 1 1 12461
0 12463 7 1 2 12460 12462
0 12464 5 1 1 12463
0 12465 7 1 2 48598 12464
0 12466 5 1 1 12465
0 12467 7 2 2 43575 47412
0 12468 7 1 2 52266 55754
0 12469 7 1 2 64321 12468
0 12470 7 1 2 56261 60287
0 12471 7 1 2 63473 12470
0 12472 7 1 2 12469 12471
0 12473 5 1 1 12472
0 12474 7 1 2 12466 12473
0 12475 5 1 1 12474
0 12476 7 1 2 55573 12475
0 12477 5 1 1 12476
0 12478 7 3 2 52084 57706
0 12479 5 1 1 64323
0 12480 7 1 2 62011 64324
0 12481 5 1 1 12480
0 12482 7 1 2 46475 57184
0 12483 5 1 1 12482
0 12484 7 1 2 47252 58806
0 12485 5 1 1 12484
0 12486 7 1 2 12483 12485
0 12487 5 1 1 12486
0 12488 7 1 2 50760 12487
0 12489 5 1 1 12488
0 12490 7 1 2 54115 59032
0 12491 5 1 1 12490
0 12492 7 1 2 12489 12491
0 12493 5 1 1 12492
0 12494 7 1 2 61516 12493
0 12495 5 1 1 12494
0 12496 7 1 2 12481 12495
0 12497 5 1 1 12496
0 12498 7 1 2 46008 12497
0 12499 5 1 1 12498
0 12500 7 1 2 49278 62440
0 12501 5 1 1 12500
0 12502 7 1 2 47253 52884
0 12503 5 1 1 12502
0 12504 7 1 2 50761 55368
0 12505 7 1 2 12503 12504
0 12506 5 1 1 12505
0 12507 7 1 2 12501 12506
0 12508 5 1 1 12507
0 12509 7 1 2 43720 12508
0 12510 5 1 1 12509
0 12511 7 1 2 54000 64325
0 12512 5 1 1 12511
0 12513 7 1 2 12510 12512
0 12514 5 1 1 12513
0 12515 7 1 2 63243 12514
0 12516 5 1 1 12515
0 12517 7 1 2 46214 12516
0 12518 7 1 2 12499 12517
0 12519 5 1 1 12518
0 12520 7 1 2 1043 58602
0 12521 5 5 1 12520
0 12522 7 1 2 51703 64326
0 12523 5 1 1 12522
0 12524 7 1 2 52896 54339
0 12525 5 1 1 12524
0 12526 7 1 2 12523 12525
0 12527 5 1 1 12526
0 12528 7 1 2 53259 12527
0 12529 5 1 1 12528
0 12530 7 3 2 49279 58494
0 12531 7 4 2 50185 55139
0 12532 7 1 2 64331 64334
0 12533 5 1 1 12532
0 12534 7 1 2 12529 12533
0 12535 5 1 1 12534
0 12536 7 1 2 60384 12535
0 12537 5 1 1 12536
0 12538 7 1 2 42762 9268
0 12539 7 1 2 12537 12538
0 12540 5 1 1 12539
0 12541 7 1 2 62917 12540
0 12542 7 1 2 12519 12541
0 12543 5 1 1 12542
0 12544 7 1 2 12477 12543
0 12545 7 1 2 12442 12544
0 12546 5 1 1 12545
0 12547 7 1 2 62493 12546
0 12548 5 1 1 12547
0 12549 7 3 2 61565 63442
0 12550 7 1 2 45230 59080
0 12551 5 1 1 12550
0 12552 7 2 2 52340 12551
0 12553 7 1 2 44051 64341
0 12554 5 1 1 12553
0 12555 7 1 2 47254 52347
0 12556 5 1 1 12555
0 12557 7 1 2 12554 12556
0 12558 5 1 1 12557
0 12559 7 1 2 42763 12558
0 12560 5 1 1 12559
0 12561 7 1 2 49537 57185
0 12562 5 1 1 12561
0 12563 7 1 2 55293 62452
0 12564 5 1 1 12563
0 12565 7 1 2 12562 12564
0 12566 7 1 2 12560 12565
0 12567 5 1 1 12566
0 12568 7 1 2 43721 12567
0 12569 5 1 1 12568
0 12570 7 3 2 49487 52224
0 12571 5 1 1 64343
0 12572 7 1 2 47096 64344
0 12573 5 1 1 12572
0 12574 7 1 2 6949 12573
0 12575 5 1 1 12574
0 12576 7 1 2 51974 12575
0 12577 5 1 1 12576
0 12578 7 1 2 46009 12577
0 12579 7 1 2 12569 12578
0 12580 5 1 1 12579
0 12581 7 1 2 53726 56806
0 12582 5 1 1 12581
0 12583 7 1 2 50328 50762
0 12584 5 3 1 12583
0 12585 7 1 2 56726 64346
0 12586 7 1 2 57478 12585
0 12587 5 1 1 12586
0 12588 7 1 2 12582 12587
0 12589 5 1 1 12588
0 12590 7 1 2 47097 12589
0 12591 5 1 1 12590
0 12592 7 1 2 47413 57471
0 12593 5 1 1 12592
0 12594 7 1 2 59083 60840
0 12595 5 1 1 12594
0 12596 7 1 2 12593 12595
0 12597 5 1 1 12596
0 12598 7 1 2 45231 12597
0 12599 5 1 1 12598
0 12600 7 1 2 42517 12599
0 12601 7 1 2 12591 12600
0 12602 5 1 1 12601
0 12603 7 1 2 48097 12602
0 12604 7 1 2 12580 12603
0 12605 5 1 1 12604
0 12606 7 2 2 58462 61339
0 12607 7 5 2 44752 48599
0 12608 7 2 2 51366 64351
0 12609 7 1 2 43883 64356
0 12610 7 1 2 64349 12609
0 12611 5 1 1 12610
0 12612 7 1 2 12605 12611
0 12613 5 1 1 12612
0 12614 7 1 2 64338 12613
0 12615 5 1 1 12614
0 12616 7 3 2 56693 63647
0 12617 7 1 2 53260 64358
0 12618 5 1 1 12617
0 12619 7 1 2 58495 60849
0 12620 5 1 1 12619
0 12621 7 1 2 12618 12620
0 12622 5 1 1 12621
0 12623 7 1 2 60385 12622
0 12624 5 1 1 12623
0 12625 7 1 2 55054 62072
0 12626 5 1 1 12625
0 12627 7 1 2 12624 12626
0 12628 5 1 1 12627
0 12629 7 1 2 58369 62918
0 12630 7 1 2 12628 12629
0 12631 5 1 1 12630
0 12632 7 1 2 12615 12631
0 12633 5 1 1 12632
0 12634 7 1 2 43063 12633
0 12635 5 1 1 12634
0 12636 7 3 2 54866 61993
0 12637 5 9 1 64361
0 12638 7 1 2 59084 64364
0 12639 5 1 1 12638
0 12640 7 1 2 58556 60165
0 12641 5 1 1 12640
0 12642 7 1 2 42764 12641
0 12643 5 1 1 12642
0 12644 7 1 2 12639 12643
0 12645 5 1 1 12644
0 12646 7 1 2 54174 12645
0 12647 5 1 1 12646
0 12648 7 1 2 52736 64342
0 12649 5 1 1 12648
0 12650 7 4 2 46476 59085
0 12651 5 2 1 64373
0 12652 7 1 2 63515 64377
0 12653 5 1 1 12652
0 12654 7 1 2 54116 12653
0 12655 5 1 1 12654
0 12656 7 1 2 12649 12655
0 12657 5 1 1 12656
0 12658 7 1 2 51138 12657
0 12659 5 1 1 12658
0 12660 7 1 2 12647 12659
0 12661 5 1 1 12660
0 12662 7 1 2 62732 12661
0 12663 5 1 1 12662
0 12664 7 2 2 48961 54134
0 12665 7 4 2 46963 47535
0 12666 7 1 2 47641 64381
0 12667 7 1 2 64379 12666
0 12668 7 2 2 45799 55150
0 12669 7 5 2 46662 55797
0 12670 7 1 2 64385 64387
0 12671 7 1 2 12667 12670
0 12672 5 1 1 12671
0 12673 7 1 2 53261 62733
0 12674 7 1 2 57882 12673
0 12675 5 1 1 12674
0 12676 7 1 2 12672 12675
0 12677 5 1 1 12676
0 12678 7 1 2 60288 12677
0 12679 5 1 1 12678
0 12680 7 1 2 12663 12679
0 12681 5 1 1 12680
0 12682 7 1 2 60386 12681
0 12683 5 1 1 12682
0 12684 7 13 2 42267 46010
0 12685 7 2 2 45232 64392
0 12686 7 3 2 59514 63418
0 12687 7 1 2 64405 64407
0 12688 7 1 2 62227 12687
0 12689 7 1 2 64154 12688
0 12690 5 1 1 12689
0 12691 7 1 2 12683 12690
0 12692 7 1 2 12635 12691
0 12693 5 1 1 12692
0 12694 7 1 2 60446 12693
0 12695 5 1 1 12694
0 12696 7 1 2 12548 12695
0 12697 5 1 1 12696
0 12698 7 1 2 51919 12697
0 12699 5 1 1 12698
0 12700 7 1 2 49973 63914
0 12701 5 2 1 12700
0 12702 7 2 2 62409 64410
0 12703 5 1 1 64412
0 12704 7 1 2 55132 57707
0 12705 5 1 1 12704
0 12706 7 1 2 64413 12705
0 12707 5 1 1 12706
0 12708 7 1 2 43722 12707
0 12709 5 1 1 12708
0 12710 7 2 2 51336 54843
0 12711 5 1 1 64414
0 12712 7 1 2 62411 64415
0 12713 5 1 1 12712
0 12714 7 1 2 12709 12713
0 12715 5 1 1 12714
0 12716 7 1 2 54080 12715
0 12717 5 1 1 12716
0 12718 7 4 2 48098 63463
0 12719 5 1 1 64416
0 12720 7 6 2 48600 54308
0 12721 5 1 1 64420
0 12722 7 1 2 57194 64421
0 12723 5 1 1 12722
0 12724 7 1 2 12719 12723
0 12725 5 1 1 12724
0 12726 7 1 2 43064 12725
0 12727 5 1 1 12726
0 12728 7 1 2 61732 63373
0 12729 5 1 1 12728
0 12730 7 1 2 12727 12729
0 12731 5 1 1 12730
0 12732 7 1 2 51704 12731
0 12733 5 1 1 12732
0 12734 7 1 2 57220 12703
0 12735 5 1 1 12734
0 12736 7 1 2 54355 64357
0 12737 5 1 1 12736
0 12738 7 1 2 12735 12737
0 12739 7 1 2 12733 12738
0 12740 5 1 1 12739
0 12741 7 1 2 42518 12740
0 12742 5 1 1 12741
0 12743 7 1 2 12717 12742
0 12744 5 1 1 12743
0 12745 7 1 2 43884 12744
0 12746 5 1 1 12745
0 12747 7 1 2 57105 62443
0 12748 5 1 1 12747
0 12749 7 1 2 49337 12748
0 12750 5 1 1 12749
0 12751 7 1 2 48601 57119
0 12752 5 1 1 12751
0 12753 7 1 2 62392 12752
0 12754 7 1 2 12750 12753
0 12755 5 1 1 12754
0 12756 7 1 2 62085 12755
0 12757 5 1 1 12756
0 12758 7 1 2 52935 63491
0 12759 7 1 2 62242 12758
0 12760 5 1 1 12759
0 12761 7 1 2 12757 12760
0 12762 5 1 1 12761
0 12763 7 1 2 48099 12762
0 12764 5 1 1 12763
0 12765 7 1 2 12746 12764
0 12766 5 1 1 12765
0 12767 7 1 2 44637 12766
0 12768 5 1 1 12767
0 12769 7 1 2 61984 63460
0 12770 5 1 1 12769
0 12771 7 1 2 44195 64166
0 12772 5 1 1 12771
0 12773 7 1 2 61727 62460
0 12774 5 1 1 12773
0 12775 7 1 2 12772 12774
0 12776 5 1 1 12775
0 12777 7 1 2 52769 12776
0 12778 5 1 1 12777
0 12779 7 1 2 12770 12778
0 12780 7 1 2 12768 12779
0 12781 5 1 1 12780
0 12782 7 1 2 62734 12781
0 12783 5 1 1 12782
0 12784 7 1 2 48962 62250
0 12785 5 1 1 12784
0 12786 7 1 2 62352 12785
0 12787 5 1 1 12786
0 12788 7 1 2 46663 12787
0 12789 5 1 1 12788
0 12790 7 1 2 56703 64162
0 12791 5 1 1 12790
0 12792 7 1 2 12789 12791
0 12793 5 1 1 12792
0 12794 7 10 2 47642 44638
0 12795 7 1 2 48100 64426
0 12796 7 1 2 63007 12795
0 12797 7 1 2 59063 12796
0 12798 7 1 2 12793 12797
0 12799 5 1 1 12798
0 12800 7 1 2 12783 12799
0 12801 5 1 1 12800
0 12802 7 1 2 60447 12801
0 12803 5 1 1 12802
0 12804 7 1 2 49974 52770
0 12805 5 1 1 12804
0 12806 7 1 2 50155 58041
0 12807 5 1 1 12806
0 12808 7 1 2 12805 12807
0 12809 5 1 1 12808
0 12810 7 1 2 45233 12809
0 12811 5 1 1 12810
0 12812 7 5 2 48602 50763
0 12813 5 1 1 64436
0 12814 7 1 2 52041 64437
0 12815 5 1 1 12814
0 12816 7 1 2 12811 12815
0 12817 5 1 1 12816
0 12818 7 1 2 62919 12817
0 12819 5 1 1 12818
0 12820 7 7 2 46215 43454
0 12821 7 1 2 64092 64441
0 12822 7 1 2 63348 12821
0 12823 5 2 1 12822
0 12824 7 1 2 12819 64448
0 12825 5 1 1 12824
0 12826 7 1 2 61377 12825
0 12827 5 1 1 12826
0 12828 7 1 2 46216 50199
0 12829 5 1 1 12828
0 12830 7 1 2 62735 12829
0 12831 5 1 1 12830
0 12832 7 1 2 43274 62736
0 12833 5 1 1 12832
0 12834 7 1 2 61089 62986
0 12835 7 1 2 63683 12834
0 12836 5 1 1 12835
0 12837 7 1 2 12833 12836
0 12838 5 1 1 12837
0 12839 7 1 2 44052 12838
0 12840 5 1 1 12839
0 12841 7 1 2 12831 12840
0 12842 5 1 1 12841
0 12843 7 1 2 43885 12842
0 12844 5 1 1 12843
0 12845 7 1 2 53020 60599
0 12846 7 1 2 63443 12845
0 12847 5 1 1 12846
0 12848 7 1 2 12844 12847
0 12849 5 1 1 12848
0 12850 7 1 2 53262 12849
0 12851 5 1 1 12850
0 12852 7 4 2 43723 45234
0 12853 7 1 2 50894 64450
0 12854 5 1 1 12853
0 12855 7 1 2 43065 58101
0 12856 5 1 1 12855
0 12857 7 1 2 12854 12856
0 12858 5 1 1 12857
0 12859 7 1 2 46217 12858
0 12860 5 1 1 12859
0 12861 7 3 2 54893 61461
0 12862 7 1 2 43275 64454
0 12863 5 1 1 12862
0 12864 7 1 2 3835 12863
0 12865 5 1 1 12864
0 12866 7 1 2 47255 12865
0 12867 5 1 1 12866
0 12868 7 1 2 12860 12867
0 12869 5 1 1 12868
0 12870 7 13 2 42268 42519
0 12871 7 2 2 59515 64457
0 12872 7 1 2 63419 64470
0 12873 7 1 2 12869 12872
0 12874 5 1 1 12873
0 12875 7 1 2 12851 12874
0 12876 5 1 1 12875
0 12877 7 1 2 60387 12876
0 12878 5 1 1 12877
0 12879 7 1 2 12827 12878
0 12880 5 1 1 12879
0 12881 7 1 2 45440 12880
0 12882 5 1 1 12881
0 12883 7 1 2 54540 62429
0 12884 5 1 1 12883
0 12885 7 1 2 53263 53384
0 12886 5 1 1 12885
0 12887 7 1 2 55694 60266
0 12888 5 1 1 12887
0 12889 7 3 2 64149 12888
0 12890 7 1 2 49584 64472
0 12891 5 1 1 12890
0 12892 7 1 2 12886 12891
0 12893 5 1 1 12892
0 12894 7 1 2 51650 12893
0 12895 5 1 1 12894
0 12896 7 1 2 12884 12895
0 12897 5 1 1 12896
0 12898 7 1 2 64339 12897
0 12899 5 1 1 12898
0 12900 7 2 2 61142 63464
0 12901 7 1 2 46964 64475
0 12902 7 1 2 64313 12901
0 12903 5 1 1 12902
0 12904 7 2 2 44753 52095
0 12905 7 2 2 51139 51975
0 12906 7 1 2 64477 64479
0 12907 5 1 1 12906
0 12908 7 1 2 60267 61994
0 12909 7 1 2 63598 12908
0 12910 5 1 1 12909
0 12911 7 1 2 53264 12910
0 12912 5 1 1 12911
0 12913 7 2 2 48603 54383
0 12914 7 1 2 52957 61708
0 12915 7 1 2 64481 12914
0 12916 5 1 1 12915
0 12917 7 1 2 12912 12916
0 12918 5 1 1 12917
0 12919 7 1 2 48101 12918
0 12920 5 1 1 12919
0 12921 7 1 2 12907 12920
0 12922 5 1 1 12921
0 12923 7 1 2 48801 64340
0 12924 7 1 2 12922 12923
0 12925 5 1 1 12924
0 12926 7 1 2 12903 12925
0 12927 5 1 1 12926
0 12928 7 1 2 44196 12927
0 12929 5 1 1 12928
0 12930 7 3 2 44319 44754
0 12931 7 1 2 61340 62125
0 12932 7 1 2 64483 12931
0 12933 7 1 2 62049 12932
0 12934 7 1 2 63446 12933
0 12935 5 1 1 12934
0 12936 7 1 2 12929 12935
0 12937 5 1 1 12936
0 12938 7 1 2 43276 12937
0 12939 5 1 1 12938
0 12940 7 1 2 12899 12939
0 12941 7 1 2 12882 12940
0 12942 5 1 1 12941
0 12943 7 1 2 62494 12942
0 12944 5 1 1 12943
0 12945 7 6 2 45800 50408
0 12946 7 2 2 46965 64486
0 12947 7 4 2 42009 57907
0 12948 7 8 2 47643 44755
0 12949 7 1 2 53945 64498
0 12950 7 1 2 57618 12949
0 12951 7 1 2 64494 12950
0 12952 7 1 2 64492 12951
0 12953 5 1 1 12952
0 12954 7 1 2 52003 62737
0 12955 5 1 1 12954
0 12956 7 1 2 62597 62920
0 12957 5 1 1 12956
0 12958 7 1 2 12955 12957
0 12959 5 1 1 12958
0 12960 7 1 2 49280 12959
0 12961 5 1 1 12960
0 12962 7 1 2 64449 12961
0 12963 5 1 1 12962
0 12964 7 1 2 43724 12963
0 12965 5 1 1 12964
0 12966 7 1 2 63199 64223
0 12967 5 1 1 12966
0 12968 7 1 2 12965 12967
0 12969 5 1 1 12968
0 12970 7 1 2 42520 12969
0 12971 5 1 1 12970
0 12972 7 4 2 43576 43725
0 12973 7 1 2 64393 64506
0 12974 7 1 2 63186 12973
0 12975 7 1 2 52116 12974
0 12976 5 1 1 12975
0 12977 7 1 2 12971 12976
0 12978 5 1 1 12977
0 12979 7 1 2 60388 63701
0 12980 7 1 2 12978 12979
0 12981 5 1 1 12980
0 12982 7 1 2 12953 12981
0 12983 5 1 1 12982
0 12984 7 1 2 50070 12983
0 12985 5 1 1 12984
0 12986 7 2 2 56186 61603
0 12987 5 1 1 64510
0 12988 7 1 2 43066 63476
0 12989 5 1 1 12988
0 12990 7 1 2 12987 12989
0 12991 5 1 1 12990
0 12992 7 1 2 62266 12991
0 12993 5 1 1 12992
0 12994 7 2 2 48802 62495
0 12995 7 1 2 52666 64512
0 12996 5 1 1 12995
0 12997 7 1 2 52958 63702
0 12998 5 1 1 12997
0 12999 7 1 2 12996 12998
0 13000 5 1 1 12999
0 13001 7 1 2 62086 13000
0 13002 5 1 1 13001
0 13003 7 1 2 54713 63703
0 13004 5 1 1 13003
0 13005 7 1 2 47414 64511
0 13006 5 1 1 13005
0 13007 7 1 2 13004 13006
0 13008 5 1 1 13007
0 13009 7 1 2 62645 13008
0 13010 5 1 1 13009
0 13011 7 1 2 13002 13010
0 13012 5 1 1 13011
0 13013 7 1 2 45235 13012
0 13014 5 1 1 13013
0 13015 7 2 2 61449 64193
0 13016 7 1 2 53265 52943
0 13017 7 1 2 64514 13016
0 13018 5 1 1 13017
0 13019 7 1 2 13014 13018
0 13020 5 1 1 13019
0 13021 7 1 2 60389 13020
0 13022 5 1 1 13021
0 13023 7 1 2 12993 13022
0 13024 5 1 1 13023
0 13025 7 1 2 62921 13024
0 13026 5 1 1 13025
0 13027 7 1 2 43067 64473
0 13028 5 1 1 13027
0 13029 7 1 2 64285 13028
0 13030 5 1 1 13029
0 13031 7 1 2 50454 13030
0 13032 5 1 1 13031
0 13033 7 3 2 42521 50611
0 13034 5 2 1 64516
0 13035 7 1 2 52058 64517
0 13036 5 1 1 13035
0 13037 7 1 2 49692 56338
0 13038 5 1 1 13037
0 13039 7 1 2 13036 13038
0 13040 5 1 1 13039
0 13041 7 1 2 47098 13040
0 13042 5 1 1 13041
0 13043 7 1 2 13032 13042
0 13044 5 1 1 13043
0 13045 7 12 2 44439 44639
0 13046 7 2 2 48102 64521
0 13047 7 2 2 42010 64533
0 13048 7 1 2 13044 64535
0 13049 5 1 1 13048
0 13050 7 6 2 47756 47966
0 13051 7 3 2 44756 64537
0 13052 7 1 2 47099 58255
0 13053 7 1 2 64543 13052
0 13054 7 1 2 56090 13053
0 13055 5 1 1 13054
0 13056 7 1 2 13049 13055
0 13057 5 1 1 13056
0 13058 7 1 2 62738 13057
0 13059 5 1 1 13058
0 13060 7 1 2 13026 13059
0 13061 5 1 1 13060
0 13062 7 1 2 55574 13061
0 13063 5 1 1 13062
0 13064 7 1 2 50178 51783
0 13065 5 2 1 13064
0 13066 7 11 2 60767 64546
0 13067 7 3 2 43577 44440
0 13068 7 2 2 59516 64559
0 13069 7 4 2 42011 42765
0 13070 7 2 2 63320 64564
0 13071 7 1 2 64562 64568
0 13072 5 1 1 13071
0 13073 7 1 2 63111 64073
0 13074 7 2 2 63308 13073
0 13075 7 1 2 53852 64570
0 13076 5 1 1 13075
0 13077 7 1 2 13072 13076
0 13078 5 1 1 13077
0 13079 7 1 2 62312 13078
0 13080 5 1 1 13079
0 13081 7 1 2 62087 64571
0 13082 5 1 1 13081
0 13083 7 2 2 59194 64108
0 13084 7 5 2 43528 64560
0 13085 7 1 2 63468 64574
0 13086 7 1 2 64572 13085
0 13087 5 1 1 13086
0 13088 7 1 2 13082 13087
0 13089 5 1 1 13088
0 13090 7 1 2 57186 13089
0 13091 5 1 1 13090
0 13092 7 1 2 54163 55611
0 13093 7 1 2 63176 13092
0 13094 7 1 2 63303 63596
0 13095 7 1 2 13093 13094
0 13096 5 1 1 13095
0 13097 7 1 2 13091 13096
0 13098 7 1 2 13080 13097
0 13099 5 1 1 13098
0 13100 7 1 2 60390 13099
0 13101 5 1 1 13100
0 13102 7 2 2 63465 63662
0 13103 7 1 2 56868 63064
0 13104 7 1 2 64579 13103
0 13105 7 1 2 63306 13104
0 13106 5 1 1 13105
0 13107 7 1 2 13101 13106
0 13108 5 1 1 13107
0 13109 7 1 2 64548 13108
0 13110 5 1 1 13109
0 13111 7 1 2 13063 13110
0 13112 7 1 2 12985 13111
0 13113 7 1 2 12944 13112
0 13114 7 1 2 12803 13113
0 13115 5 1 1 13114
0 13116 7 1 2 59269 13115
0 13117 5 1 1 13116
0 13118 7 1 2 58588 63328
0 13119 5 1 1 13118
0 13120 7 2 2 53266 64208
0 13121 7 1 2 62922 64536
0 13122 7 1 2 64581 13121
0 13123 5 1 1 13122
0 13124 7 1 2 13119 13123
0 13125 5 1 1 13124
0 13126 7 1 2 60289 13125
0 13127 5 1 1 13126
0 13128 7 2 2 51474 58334
0 13129 5 1 1 64583
0 13130 7 1 2 58496 64584
0 13131 5 1 1 13130
0 13132 7 6 2 44197 59647
0 13133 5 1 1 64585
0 13134 7 2 2 50636 64586
0 13135 5 2 1 64591
0 13136 7 1 2 62444 64593
0 13137 5 1 1 13136
0 13138 7 1 2 54384 57843
0 13139 7 1 2 13137 13138
0 13140 5 1 1 13139
0 13141 7 1 2 13131 13140
0 13142 5 1 1 13141
0 13143 7 1 2 62923 13142
0 13144 5 1 1 13143
0 13145 7 1 2 51976 60720
0 13146 5 1 1 13145
0 13147 7 1 2 62113 13146
0 13148 5 1 1 13147
0 13149 7 1 2 50552 13148
0 13150 5 1 1 13149
0 13151 7 7 2 46011 48604
0 13152 5 2 1 64595
0 13153 7 1 2 62859 64596
0 13154 5 1 1 13153
0 13155 7 1 2 13150 13154
0 13156 5 1 1 13155
0 13157 7 1 2 46664 13156
0 13158 5 1 1 13157
0 13159 7 4 2 42522 47415
0 13160 7 1 2 47536 64604
0 13161 7 1 2 54120 13160
0 13162 5 1 1 13161
0 13163 7 1 2 13158 13162
0 13164 5 1 1 13163
0 13165 7 1 2 62739 13164
0 13166 5 1 1 13165
0 13167 7 1 2 13144 13166
0 13168 5 1 1 13167
0 13169 7 1 2 43726 13168
0 13170 5 1 1 13169
0 13171 7 2 2 55408 59517
0 13172 7 1 2 60321 62860
0 13173 7 1 2 64608 13172
0 13174 5 1 1 13173
0 13175 7 1 2 51705 54015
0 13176 7 1 2 63668 13175
0 13177 5 1 1 13176
0 13178 7 1 2 13174 13177
0 13179 5 1 1 13178
0 13180 7 1 2 48605 13179
0 13181 5 1 1 13180
0 13182 7 2 2 51079 60928
0 13183 7 2 2 43886 63065
0 13184 7 12 2 45801 42766
0 13185 7 1 2 58278 64614
0 13186 7 1 2 64612 13185
0 13187 7 1 2 64610 13186
0 13188 5 1 1 13187
0 13189 7 1 2 13181 13188
0 13190 5 1 1 13189
0 13191 7 1 2 53198 13190
0 13192 5 1 1 13191
0 13193 7 1 2 13170 13192
0 13194 5 1 1 13193
0 13195 7 1 2 60391 13194
0 13196 5 1 1 13195
0 13197 7 1 2 52004 52308
0 13198 7 1 2 62953 13197
0 13199 5 1 1 13198
0 13200 7 1 2 50343 13199
0 13201 5 1 1 13200
0 13202 7 1 2 46012 13201
0 13203 5 1 1 13202
0 13204 7 1 2 58502 61479
0 13205 5 1 1 13204
0 13206 7 1 2 13203 13205
0 13207 5 1 1 13206
0 13208 7 1 2 47100 13207
0 13209 5 1 1 13208
0 13210 7 1 2 50329 58526
0 13211 5 1 1 13210
0 13212 7 1 2 13209 13211
0 13213 5 1 1 13212
0 13214 7 1 2 45236 13213
0 13215 5 1 1 13214
0 13216 7 1 2 52757 53330
0 13217 5 1 1 13216
0 13218 7 2 2 47101 49158
0 13219 7 1 2 58396 64626
0 13220 7 1 2 13217 13219
0 13221 5 1 1 13220
0 13222 7 1 2 13215 13221
0 13223 5 1 1 13222
0 13224 7 1 2 61492 63444
0 13225 7 1 2 13223 13224
0 13226 5 1 1 13225
0 13227 7 1 2 13196 13226
0 13228 5 1 1 13227
0 13229 7 1 2 62496 13228
0 13230 5 1 1 13229
0 13231 7 1 2 13127 13230
0 13232 5 1 1 13231
0 13233 7 1 2 62794 13232
0 13234 5 1 1 13233
0 13235 7 2 2 43887 63807
0 13236 7 1 2 47537 64019
0 13237 7 1 2 64628 13236
0 13238 7 2 2 46218 55798
0 13239 7 3 2 47644 61302
0 13240 7 1 2 64630 64632
0 13241 7 1 2 13237 13240
0 13242 5 1 1 13241
0 13243 7 4 2 47757 63016
0 13244 7 1 2 52005 64408
0 13245 7 1 2 64635 13244
0 13246 7 1 2 51223 13245
0 13247 5 1 1 13246
0 13248 7 1 2 13242 13247
0 13249 5 1 1 13248
0 13250 7 1 2 62830 13249
0 13251 5 1 1 13250
0 13252 7 2 2 51706 59152
0 13253 7 2 2 63364 64639
0 13254 5 1 1 64641
0 13255 7 7 2 42269 43277
0 13256 7 2 2 54479 64643
0 13257 7 1 2 63971 64650
0 13258 5 1 1 13257
0 13259 7 1 2 13254 13258
0 13260 5 1 1 13259
0 13261 7 1 2 47256 13260
0 13262 5 1 1 13261
0 13263 7 4 2 46665 43578
0 13264 7 1 2 61601 64652
0 13265 7 3 2 42270 55755
0 13266 7 1 2 64656 64185
0 13267 7 1 2 13264 13266
0 13268 5 1 1 13267
0 13269 7 1 2 13262 13268
0 13270 5 1 1 13269
0 13271 7 1 2 55101 13270
0 13272 5 1 1 13271
0 13273 7 1 2 55059 64642
0 13274 5 1 1 13273
0 13275 7 1 2 13272 13274
0 13276 5 1 1 13275
0 13277 7 1 2 51920 13276
0 13278 5 1 1 13277
0 13279 7 1 2 13251 13278
0 13280 5 1 1 13279
0 13281 7 1 2 42523 13280
0 13282 5 1 1 13281
0 13283 7 3 2 54385 55799
0 13284 7 5 2 45802 43727
0 13285 7 1 2 51921 64662
0 13286 7 1 2 64629 13285
0 13287 7 1 2 64659 13286
0 13288 7 1 2 64640 13287
0 13289 5 1 1 13288
0 13290 7 1 2 13282 13289
0 13291 5 1 1 13290
0 13292 7 1 2 60392 13291
0 13293 5 1 1 13292
0 13294 7 1 2 52042 63471
0 13295 7 1 2 63553 64036
0 13296 7 1 2 13294 13295
0 13297 5 1 1 13296
0 13298 7 1 2 63034 64253
0 13299 5 1 1 13298
0 13300 7 1 2 56793 57123
0 13301 5 1 1 13300
0 13302 7 5 2 46219 62497
0 13303 7 1 2 62924 64667
0 13304 7 1 2 13301 13303
0 13305 5 1 1 13304
0 13306 7 1 2 13299 13305
0 13307 5 1 1 13306
0 13308 7 1 2 52006 59270
0 13309 7 1 2 13307 13308
0 13310 5 1 1 13309
0 13311 7 1 2 13297 13310
0 13312 5 1 1 13311
0 13313 7 1 2 61195 13312
0 13314 5 1 1 13313
0 13315 7 1 2 13293 13314
0 13316 5 1 1 13315
0 13317 7 1 2 45237 13316
0 13318 5 1 1 13317
0 13319 7 1 2 63886 63778
0 13320 5 1 1 13319
0 13321 7 1 2 63674 64033
0 13322 7 1 2 64657 13321
0 13323 5 1 1 13322
0 13324 7 1 2 13320 13323
0 13325 5 1 1 13324
0 13326 7 1 2 43278 13325
0 13327 5 1 1 13326
0 13328 7 1 2 55958 64653
0 13329 7 1 2 61898 13328
0 13330 7 1 2 63866 13329
0 13331 5 1 1 13330
0 13332 7 1 2 13327 13331
0 13333 5 1 1 13332
0 13334 7 1 2 61378 13333
0 13335 5 1 1 13334
0 13336 7 1 2 63035 64270
0 13337 5 1 1 13336
0 13338 7 1 2 13335 13337
0 13339 5 1 1 13338
0 13340 7 1 2 52043 13339
0 13341 5 1 1 13340
0 13342 7 1 2 13318 13341
0 13343 5 1 1 13342
0 13344 7 1 2 50997 13343
0 13345 5 1 1 13344
0 13346 7 1 2 61705 62651
0 13347 5 1 1 13346
0 13348 7 1 2 61517 62104
0 13349 5 1 1 13348
0 13350 7 1 2 13347 13349
0 13351 5 1 1 13350
0 13352 7 1 2 42767 13351
0 13353 5 1 1 13352
0 13354 7 4 2 46220 51057
0 13355 7 1 2 53968 61143
0 13356 7 1 2 64672 13355
0 13357 5 1 1 13356
0 13358 7 1 2 13353 13357
0 13359 5 1 1 13358
0 13360 7 1 2 62925 63722
0 13361 7 1 2 13359 13360
0 13362 5 1 1 13361
0 13363 7 1 2 52748 62576
0 13364 5 1 1 13363
0 13365 7 1 2 54342 58795
0 13366 5 1 1 13365
0 13367 7 1 2 46477 13366
0 13368 5 1 1 13367
0 13369 7 1 2 47416 54340
0 13370 5 1 1 13369
0 13371 7 1 2 62207 13370
0 13372 7 1 2 13368 13371
0 13373 5 1 1 13372
0 13374 7 1 2 46221 13373
0 13375 5 1 1 13374
0 13376 7 1 2 13364 13375
0 13377 5 1 1 13376
0 13378 7 1 2 61518 64409
0 13379 7 1 2 64636 13378
0 13380 7 1 2 13377 13379
0 13381 5 1 1 13380
0 13382 7 1 2 13362 13381
0 13383 5 1 1 13382
0 13384 7 1 2 45238 13383
0 13385 5 1 1 13384
0 13386 7 1 2 58796 12813
0 13387 5 1 1 13386
0 13388 7 1 2 47257 13387
0 13389 5 1 1 13388
0 13390 7 1 2 48606 56712
0 13391 5 1 1 13390
0 13392 7 1 2 62208 13391
0 13393 5 1 1 13392
0 13394 7 1 2 46478 13393
0 13395 5 1 1 13394
0 13396 7 1 2 13389 13395
0 13397 5 1 1 13396
0 13398 7 1 2 44320 54095
0 13399 7 1 2 64544 13398
0 13400 7 1 2 63036 13399
0 13401 7 1 2 13397 13400
0 13402 5 1 1 13401
0 13403 7 1 2 13385 13402
0 13404 5 1 1 13403
0 13405 7 1 2 46013 13404
0 13406 5 1 1 13405
0 13407 7 2 2 43068 54001
0 13408 5 1 1 64676
0 13409 7 1 2 57692 13408
0 13410 5 1 1 13409
0 13411 7 1 2 42768 13410
0 13412 5 1 1 13411
0 13413 7 1 2 43728 52985
0 13414 7 1 2 52737 13413
0 13415 5 1 1 13414
0 13416 7 1 2 13412 13415
0 13417 5 1 1 13416
0 13418 7 1 2 44640 50071
0 13419 7 1 2 52267 63236
0 13420 7 1 2 13418 13419
0 13421 7 20 2 42012 45803
0 13422 7 4 2 44441 64678
0 13423 7 1 2 63309 64698
0 13424 7 1 2 13420 13423
0 13425 7 1 2 13417 13424
0 13426 5 1 1 13425
0 13427 7 1 2 13406 13426
0 13428 5 1 1 13427
0 13429 7 1 2 64232 13428
0 13430 5 1 1 13429
0 13431 7 1 2 56999 63544
0 13432 5 1 1 13431
0 13433 7 1 2 51922 55827
0 13434 7 1 2 58985 58969
0 13435 7 1 2 13433 13434
0 13436 5 1 1 13435
0 13437 7 1 2 13432 13436
0 13438 5 1 1 13437
0 13439 7 1 2 46666 13438
0 13440 5 1 1 13439
0 13441 7 2 2 47538 55778
0 13442 7 2 2 42164 63891
0 13443 7 1 2 64702 64704
0 13444 5 1 1 13443
0 13445 7 1 2 13440 13444
0 13446 5 1 1 13445
0 13447 7 1 2 62297 13446
0 13448 5 1 1 13447
0 13449 7 1 2 62939 64063
0 13450 5 1 1 13449
0 13451 7 1 2 13448 13450
0 13452 5 1 1 13451
0 13453 7 1 2 64058 13452
0 13454 5 1 1 13453
0 13455 7 1 2 62610 64127
0 13456 5 1 1 13455
0 13457 7 1 2 61813 62614
0 13458 7 1 2 62612 13457
0 13459 5 1 1 13458
0 13460 7 1 2 13456 13459
0 13461 5 1 1 13460
0 13462 7 1 2 48803 62747
0 13463 5 1 1 13462
0 13464 7 1 2 64059 13463
0 13465 7 1 2 13461 13464
0 13466 5 1 1 13465
0 13467 7 1 2 13454 13466
0 13468 7 1 2 13430 13467
0 13469 7 1 2 13345 13468
0 13470 7 1 2 13234 13469
0 13471 7 1 2 13117 13470
0 13472 7 1 2 12699 13471
0 13473 5 1 1 13472
0 13474 7 1 2 48407 13473
0 13475 5 1 1 13474
0 13476 7 1 2 62748 11209
0 13477 5 1 1 13476
0 13478 7 1 2 63545 13477
0 13479 5 1 1 13478
0 13480 7 1 2 45562 63140
0 13481 7 3 2 42271 55858
0 13482 7 1 2 63972 64706
0 13483 7 1 2 13480 13482
0 13484 5 1 1 13483
0 13485 7 1 2 13479 13484
0 13486 5 1 1 13485
0 13487 7 1 2 44053 13486
0 13488 5 1 1 13487
0 13489 7 2 2 56233 64658
0 13490 7 1 2 55789 63280
0 13491 7 1 2 64709 13490
0 13492 5 1 1 13491
0 13493 7 1 2 13488 13492
0 13494 5 1 1 13493
0 13495 7 1 2 62940 13494
0 13496 5 1 1 13495
0 13497 7 13 2 42272 44561
0 13498 7 1 2 48893 56076
0 13499 7 1 2 64711 13498
0 13500 7 1 2 53328 64563
0 13501 7 1 2 13499 13500
0 13502 7 1 2 62890 13501
0 13503 5 1 1 13502
0 13504 7 1 2 13496 13503
0 13505 5 1 1 13504
0 13506 7 1 2 55575 13505
0 13507 5 1 1 13506
0 13508 7 1 2 51501 55068
0 13509 5 1 1 13508
0 13510 7 1 2 55041 59507
0 13511 5 1 1 13510
0 13512 7 1 2 13509 13511
0 13513 5 1 1 13512
0 13514 7 1 2 51923 13513
0 13515 5 1 1 13514
0 13516 7 7 2 46222 45239
0 13517 5 1 1 64724
0 13518 7 1 2 54935 64725
0 13519 7 1 2 62818 13518
0 13520 5 1 1 13519
0 13521 7 1 2 13515 13520
0 13522 5 1 1 13521
0 13523 7 1 2 44198 13522
0 13524 5 1 1 13523
0 13525 7 1 2 53021 54002
0 13526 7 1 2 63131 13525
0 13527 5 1 1 13526
0 13528 7 1 2 13524 13527
0 13529 5 1 1 13528
0 13530 7 1 2 43279 13529
0 13531 5 1 1 13530
0 13532 7 1 2 42165 61201
0 13533 5 1 1 13532
0 13534 7 1 2 51829 13533
0 13535 5 1 1 13534
0 13536 7 1 2 46667 13535
0 13537 5 1 1 13536
0 13538 7 1 2 49338 62854
0 13539 5 2 1 13538
0 13540 7 1 2 13537 64731
0 13541 5 1 1 13540
0 13542 7 1 2 48607 13541
0 13543 5 1 1 13542
0 13544 7 1 2 51825 59181
0 13545 5 1 1 13544
0 13546 7 1 2 13543 13545
0 13547 5 1 1 13546
0 13548 7 1 2 55042 13547
0 13549 5 1 1 13548
0 13550 7 1 2 13531 13549
0 13551 5 1 1 13550
0 13552 7 1 2 42524 13551
0 13553 5 1 1 13552
0 13554 7 1 2 62822 62937
0 13555 5 2 1 13554
0 13556 7 2 2 47258 57323
0 13557 7 1 2 57469 64735
0 13558 5 1 1 13557
0 13559 7 5 2 42769 56778
0 13560 5 1 1 64737
0 13561 7 1 2 63374 64738
0 13562 5 1 1 13561
0 13563 7 1 2 13558 13562
0 13564 5 1 1 13563
0 13565 7 1 2 42525 13564
0 13566 5 1 1 13565
0 13567 7 1 2 53187 56772
0 13568 5 1 1 13567
0 13569 7 1 2 13566 13568
0 13570 5 1 1 13569
0 13571 7 1 2 64733 13570
0 13572 5 1 1 13571
0 13573 7 1 2 43280 56896
0 13574 5 1 1 13573
0 13575 7 1 2 50631 13574
0 13576 5 1 1 13575
0 13577 7 1 2 49628 62387
0 13578 5 1 1 13577
0 13579 7 1 2 13576 13578
0 13580 5 1 1 13579
0 13581 7 1 2 51924 13580
0 13582 5 1 1 13581
0 13583 7 1 2 43281 50612
0 13584 5 3 1 13583
0 13585 7 1 2 58820 64742
0 13586 5 1 1 13585
0 13587 7 1 2 53349 59271
0 13588 7 1 2 13586 13587
0 13589 5 1 1 13588
0 13590 7 1 2 13582 13589
0 13591 5 1 1 13590
0 13592 7 1 2 59054 13591
0 13593 5 1 1 13592
0 13594 7 1 2 13572 13593
0 13595 7 1 2 13553 13594
0 13596 5 1 1 13595
0 13597 7 1 2 60393 13596
0 13598 5 1 1 13597
0 13599 7 2 2 56801 57348
0 13600 7 1 2 64734 64745
0 13601 5 1 1 13600
0 13602 7 1 2 48999 62778
0 13603 5 1 1 13602
0 13604 7 1 2 52399 59272
0 13605 7 1 2 49108 13604
0 13606 5 1 1 13605
0 13607 7 1 2 13603 13606
0 13608 5 1 1 13607
0 13609 7 1 2 43282 13608
0 13610 5 1 1 13609
0 13611 7 14 2 42166 46668
0 13612 7 6 2 44562 64747
0 13613 7 1 2 52377 64761
0 13614 5 1 1 13613
0 13615 7 1 2 13610 13614
0 13616 5 1 1 13615
0 13617 7 2 2 47417 52007
0 13618 5 1 1 64767
0 13619 7 1 2 13616 64768
0 13620 5 1 1 13619
0 13621 7 1 2 13601 13620
0 13622 5 1 1 13621
0 13623 7 1 2 46479 13622
0 13624 5 1 1 13623
0 13625 7 1 2 49489 62932
0 13626 5 1 1 13625
0 13627 7 1 2 59273 59619
0 13628 5 1 1 13627
0 13629 7 1 2 13626 13628
0 13630 5 1 1 13629
0 13631 7 1 2 64746 13630
0 13632 5 1 1 13631
0 13633 7 1 2 13624 13632
0 13634 5 1 1 13633
0 13635 7 1 2 61196 13634
0 13636 5 1 1 13635
0 13637 7 1 2 13598 13636
0 13638 5 1 1 13637
0 13639 7 1 2 62498 13638
0 13640 5 1 1 13639
0 13641 7 1 2 57742 62099
0 13642 5 1 1 13641
0 13643 7 3 2 49035 51367
0 13644 7 1 2 62095 64769
0 13645 5 1 1 13644
0 13646 7 1 2 13642 13645
0 13647 5 1 1 13646
0 13648 7 1 2 51925 13647
0 13649 5 1 1 13648
0 13650 7 1 2 55069 61844
0 13651 5 1 1 13650
0 13652 7 4 2 49339 51224
0 13653 5 2 1 64772
0 13654 7 1 2 55043 64773
0 13655 5 1 1 13654
0 13656 7 1 2 13651 13655
0 13657 5 1 1 13656
0 13658 7 1 2 59274 13657
0 13659 5 1 1 13658
0 13660 7 1 2 13649 13659
0 13661 5 1 1 13660
0 13662 7 1 2 42526 13661
0 13663 5 1 1 13662
0 13664 7 1 2 59275 64774
0 13665 5 1 1 13664
0 13666 7 1 2 62390 62753
0 13667 5 1 1 13666
0 13668 7 1 2 13665 13667
0 13669 5 1 1 13668
0 13670 7 1 2 59055 13669
0 13671 5 1 1 13670
0 13672 7 1 2 13663 13671
0 13673 5 1 1 13672
0 13674 7 1 2 60394 13673
0 13675 5 1 1 13674
0 13676 7 1 2 49902 64088
0 13677 7 3 2 46480 61634
0 13678 7 1 2 64736 64778
0 13679 7 1 2 13676 13678
0 13680 5 1 1 13679
0 13681 7 1 2 13675 13680
0 13682 5 1 1 13681
0 13683 7 1 2 48608 13682
0 13684 5 1 1 13683
0 13685 7 1 2 51794 63141
0 13686 5 1 1 13685
0 13687 7 1 2 63147 13686
0 13688 5 1 1 13687
0 13689 7 1 2 44054 13688
0 13690 5 1 1 13689
0 13691 7 1 2 45240 63058
0 13692 5 1 1 13691
0 13693 7 1 2 13690 13692
0 13694 5 1 1 13693
0 13695 7 1 2 43069 13694
0 13696 5 1 1 13695
0 13697 7 2 2 42167 57873
0 13698 7 1 2 52814 64781
0 13699 5 1 1 13698
0 13700 7 1 2 13696 13699
0 13701 5 1 1 13700
0 13702 7 1 2 62941 13701
0 13703 5 1 1 13702
0 13704 7 1 2 13684 13703
0 13705 5 1 1 13704
0 13706 7 1 2 60448 13705
0 13707 5 1 1 13706
0 13708 7 1 2 13640 13707
0 13709 5 1 1 13708
0 13710 7 1 2 62740 13709
0 13711 5 1 1 13710
0 13712 7 1 2 13507 13711
0 13713 7 1 2 13475 13712
0 13714 7 1 2 12334 13713
0 13715 7 1 2 11746 13714
0 13716 7 1 2 9823 13715
0 13717 5 1 1 13716
0 13718 7 1 2 48232 13717
0 13719 5 1 1 13718
0 13720 7 2 2 57743 63160
0 13721 7 1 2 43283 60889
0 13722 5 1 1 13721
0 13723 7 1 2 60780 13722
0 13724 5 1 1 13723
0 13725 7 1 2 64783 13724
0 13726 5 1 1 13725
0 13727 7 1 2 53388 60762
0 13728 5 1 1 13727
0 13729 7 1 2 52059 7652
0 13730 5 1 1 13729
0 13731 7 1 2 56691 13730
0 13732 5 1 1 13731
0 13733 7 1 2 13728 13732
0 13734 5 1 1 13733
0 13735 7 2 2 61662 13734
0 13736 7 1 2 58995 64785
0 13737 5 1 1 13736
0 13738 7 1 2 13726 13737
0 13739 5 1 1 13738
0 13740 7 1 2 53540 13739
0 13741 5 1 1 13740
0 13742 7 3 2 46223 47886
0 13743 7 2 2 60670 64787
0 13744 5 1 1 64790
0 13745 7 1 2 52070 64791
0 13746 5 2 1 13745
0 13747 7 2 2 45441 60775
0 13748 5 1 1 64794
0 13749 7 2 2 46481 64795
0 13750 5 1 1 64796
0 13751 7 1 2 13744 13750
0 13752 5 1 1 13751
0 13753 7 2 2 49751 13752
0 13754 5 1 1 64798
0 13755 7 1 2 47539 64799
0 13756 5 1 1 13755
0 13757 7 1 2 64792 13756
0 13758 5 1 1 13757
0 13759 7 1 2 47259 13758
0 13760 5 1 1 13759
0 13761 7 1 2 46482 60890
0 13762 5 1 1 13761
0 13763 7 1 2 13748 13762
0 13764 5 2 1 13763
0 13765 7 1 2 53389 64800
0 13766 5 1 1 13765
0 13767 7 1 2 53718 64797
0 13768 5 1 1 13767
0 13769 7 1 2 13766 13768
0 13770 5 1 1 13769
0 13771 7 1 2 47540 13770
0 13772 5 1 1 13771
0 13773 7 1 2 13760 13772
0 13774 5 1 1 13773
0 13775 7 1 2 43284 13774
0 13776 5 1 1 13775
0 13777 7 1 2 62566 62579
0 13778 5 1 1 13777
0 13779 7 2 2 50764 58996
0 13780 7 1 2 47418 63850
0 13781 7 1 2 64802 13780
0 13782 5 1 1 13781
0 13783 7 1 2 48408 13782
0 13784 7 1 2 13778 13783
0 13785 7 1 2 13776 13784
0 13786 5 1 1 13785
0 13787 7 1 2 53031 64801
0 13788 5 1 1 13787
0 13789 7 1 2 13754 13788
0 13790 5 1 1 13789
0 13791 7 1 2 47541 13790
0 13792 5 1 1 13791
0 13793 7 1 2 64793 13792
0 13794 5 1 1 13793
0 13795 7 1 2 43888 13794
0 13796 5 1 1 13795
0 13797 7 1 2 42770 49210
0 13798 5 2 1 13797
0 13799 7 1 2 60776 64804
0 13800 5 1 1 13799
0 13801 7 1 2 42771 58422
0 13802 5 1 1 13801
0 13803 7 2 2 47887 13802
0 13804 7 1 2 60671 64806
0 13805 5 1 1 13804
0 13806 7 1 2 13800 13805
0 13807 5 1 1 13806
0 13808 7 1 2 49693 13807
0 13809 5 1 1 13808
0 13810 7 2 2 45715 55859
0 13811 7 1 2 63101 64808
0 13812 5 1 1 13811
0 13813 7 1 2 60891 62038
0 13814 5 1 1 13813
0 13815 7 1 2 13812 13814
0 13816 5 1 1 13815
0 13817 7 1 2 49036 13816
0 13818 5 1 1 13817
0 13819 7 1 2 49636 52182
0 13820 5 3 1 13819
0 13821 7 1 2 56860 60672
0 13822 7 1 2 64810 13821
0 13823 5 1 1 13822
0 13824 7 1 2 13818 13823
0 13825 7 1 2 13809 13824
0 13826 5 1 1 13825
0 13827 7 1 2 47260 13826
0 13828 5 1 1 13827
0 13829 7 1 2 47888 52378
0 13830 7 2 2 57324 13829
0 13831 7 1 2 56869 62654
0 13832 7 1 2 64813 13831
0 13833 5 1 1 13832
0 13834 7 1 2 13828 13833
0 13835 7 1 2 13796 13834
0 13836 5 1 1 13835
0 13837 7 1 2 43285 13836
0 13838 5 1 1 13837
0 13839 7 1 2 53791 57653
0 13840 5 1 1 13839
0 13841 7 1 2 47261 59699
0 13842 7 1 2 13840 13841
0 13843 5 1 1 13842
0 13844 7 1 2 53043 58343
0 13845 5 1 1 13844
0 13846 7 8 2 47419 52848
0 13847 5 1 1 64815
0 13848 7 1 2 47542 64816
0 13849 5 1 1 13848
0 13850 7 1 2 43889 13849
0 13851 7 1 2 13845 13850
0 13852 5 1 1 13851
0 13853 7 1 2 46669 13852
0 13854 7 1 2 13843 13853
0 13855 5 1 1 13854
0 13856 7 1 2 63206 63860
0 13857 5 1 1 13856
0 13858 7 1 2 44199 13857
0 13859 5 1 1 13858
0 13860 7 1 2 13855 13859
0 13861 5 2 1 13860
0 13862 7 1 2 60777 64823
0 13863 5 1 1 13862
0 13864 7 1 2 63204 63861
0 13865 5 1 1 13864
0 13866 7 1 2 43286 13865
0 13867 5 1 1 13866
0 13868 7 1 2 55336 64150
0 13869 7 1 2 62158 13868
0 13870 5 1 1 13869
0 13871 7 1 2 50765 13870
0 13872 5 1 1 13871
0 13873 7 2 2 13867 13872
0 13874 5 1 1 64825
0 13875 7 1 2 62567 13874
0 13876 5 1 1 13875
0 13877 7 1 2 45058 13876
0 13878 7 1 2 13863 13877
0 13879 7 1 2 13838 13878
0 13880 5 1 1 13879
0 13881 7 1 2 13786 13880
0 13882 5 1 1 13881
0 13883 7 2 2 42168 52379
0 13884 7 1 2 47889 56870
0 13885 7 1 2 64827 13884
0 13886 7 1 2 64206 13885
0 13887 5 1 1 13886
0 13888 7 1 2 13882 13887
0 13889 5 1 1 13888
0 13890 7 1 2 61144 13889
0 13891 5 1 1 13890
0 13892 7 1 2 13741 13891
0 13893 5 1 1 13892
0 13894 7 1 2 53267 13893
0 13895 5 1 1 13894
0 13896 7 1 2 61197 62572
0 13897 5 1 1 13896
0 13898 7 1 2 10506 13897
0 13899 5 1 1 13898
0 13900 7 1 2 50939 13899
0 13901 5 1 1 13900
0 13902 7 2 2 43729 49464
0 13903 7 1 2 55576 62081
0 13904 7 1 2 64829 13903
0 13905 5 1 1 13904
0 13906 7 1 2 13901 13905
0 13907 5 1 1 13906
0 13908 7 1 2 45442 13907
0 13909 5 1 1 13908
0 13910 7 1 2 44200 60999
0 13911 5 1 1 13910
0 13912 7 1 2 56005 13911
0 13913 7 1 2 61406 13912
0 13914 5 1 1 13913
0 13915 7 1 2 13909 13914
0 13916 5 1 1 13915
0 13917 7 1 2 51977 13916
0 13918 5 1 1 13917
0 13919 7 2 2 42772 64167
0 13920 5 1 1 64831
0 13921 7 1 2 44055 64832
0 13922 5 1 1 13921
0 13923 7 3 2 42527 54164
0 13924 5 1 1 64833
0 13925 7 1 2 60395 62881
0 13926 7 1 2 64834 13925
0 13927 5 1 1 13926
0 13928 7 1 2 13922 13927
0 13929 5 1 1 13928
0 13930 7 1 2 43070 13929
0 13931 5 1 1 13930
0 13932 7 1 2 55988 61379
0 13933 5 1 1 13932
0 13934 7 1 2 13920 13933
0 13935 5 1 1 13934
0 13936 7 1 2 43890 13935
0 13937 5 1 1 13936
0 13938 7 1 2 13931 13937
0 13939 5 1 1 13938
0 13940 7 1 2 49080 13939
0 13941 5 1 1 13940
0 13942 7 1 2 49037 54714
0 13943 5 1 1 13942
0 13944 7 1 2 43891 13943
0 13945 7 1 2 63872 13944
0 13946 5 1 1 13945
0 13947 7 1 2 49038 64157
0 13948 5 1 1 13947
0 13949 7 1 2 47262 56578
0 13950 7 1 2 13948 13949
0 13951 5 1 1 13950
0 13952 7 1 2 61198 13951
0 13953 7 1 2 13946 13952
0 13954 5 1 1 13953
0 13955 7 1 2 60290 62616
0 13956 5 1 1 13955
0 13957 7 3 2 43071 44641
0 13958 7 2 2 45241 64836
0 13959 7 1 2 51549 52060
0 13960 7 1 2 64839 13959
0 13961 5 1 1 13960
0 13962 7 1 2 13956 13961
0 13963 5 2 1 13962
0 13964 7 1 2 58448 64841
0 13965 5 1 1 13964
0 13966 7 1 2 43072 56310
0 13967 5 1 1 13966
0 13968 7 1 2 57146 13967
0 13969 5 2 1 13968
0 13970 7 1 2 58477 64843
0 13971 5 1 1 13970
0 13972 7 3 2 42773 56000
0 13973 5 2 1 64845
0 13974 7 2 2 51502 53969
0 13975 5 1 1 64850
0 13976 7 1 2 64848 13975
0 13977 5 1 1 13976
0 13978 7 1 2 49039 13977
0 13979 5 1 1 13978
0 13980 7 1 2 13971 13979
0 13981 5 1 1 13980
0 13982 7 1 2 60984 13981
0 13983 5 1 1 13982
0 13984 7 1 2 13965 13983
0 13985 7 1 2 13954 13984
0 13986 7 1 2 13941 13985
0 13987 5 1 1 13986
0 13988 7 1 2 43287 13987
0 13989 5 1 1 13988
0 13990 7 2 2 52183 60738
0 13991 5 1 1 64852
0 13992 7 1 2 53421 64853
0 13993 5 1 1 13992
0 13994 7 1 2 46224 52716
0 13995 5 4 1 13994
0 13996 7 1 2 47420 64854
0 13997 5 1 1 13996
0 13998 7 1 2 54867 13997
0 13999 5 1 1 13998
0 14000 7 1 2 46670 13999
0 14001 5 1 1 14000
0 14002 7 1 2 51416 57539
0 14003 5 3 1 14002
0 14004 7 1 2 44056 64858
0 14005 5 1 1 14004
0 14006 7 1 2 54904 14005
0 14007 7 1 2 14001 14006
0 14008 5 1 1 14007
0 14009 7 1 2 48804 14008
0 14010 5 1 1 14009
0 14011 7 1 2 13993 14010
0 14012 5 1 1 14011
0 14013 7 1 2 43892 14012
0 14014 5 1 1 14013
0 14015 7 1 2 52858 13991
0 14016 5 1 1 14015
0 14017 7 1 2 54242 14016
0 14018 5 1 1 14017
0 14019 7 1 2 14014 14018
0 14020 5 1 1 14019
0 14021 7 1 2 60985 14020
0 14022 5 1 1 14021
0 14023 7 1 2 49629 52008
0 14024 5 1 1 14023
0 14025 7 2 2 52061 14024
0 14026 7 1 2 60739 64861
0 14027 5 1 1 14026
0 14028 7 1 2 56727 62162
0 14029 5 1 1 14028
0 14030 7 1 2 14027 14029
0 14031 5 1 1 14030
0 14032 7 1 2 60986 14031
0 14033 5 1 1 14032
0 14034 7 1 2 56788 61424
0 14035 5 1 1 14034
0 14036 7 1 2 14033 14035
0 14037 5 1 1 14036
0 14038 7 1 2 49340 14037
0 14039 5 1 1 14038
0 14040 7 1 2 61199 64438
0 14041 7 1 2 64189 14040
0 14042 5 1 1 14041
0 14043 7 1 2 48409 14042
0 14044 7 1 2 14039 14043
0 14045 7 1 2 14022 14044
0 14046 7 1 2 13989 14045
0 14047 5 1 1 14046
0 14048 7 1 2 52380 52667
0 14049 5 1 1 14048
0 14050 7 1 2 52240 14049
0 14051 5 1 1 14050
0 14052 7 1 2 60987 14051
0 14053 5 1 1 14052
0 14054 7 2 2 48805 50409
0 14055 7 1 2 61145 64863
0 14056 7 1 2 62004 14055
0 14057 5 1 1 14056
0 14058 7 1 2 14053 14057
0 14059 5 1 1 14058
0 14060 7 1 2 44201 14059
0 14061 5 1 1 14060
0 14062 7 1 2 52917 63162
0 14063 5 1 1 14062
0 14064 7 1 2 14061 14063
0 14065 5 1 1 14064
0 14066 7 1 2 42774 14065
0 14067 5 1 1 14066
0 14068 7 1 2 52968 62618
0 14069 5 1 1 14068
0 14070 7 1 2 14067 14069
0 14071 5 1 1 14070
0 14072 7 1 2 43288 14071
0 14073 5 1 1 14072
0 14074 7 1 2 62015 62973
0 14075 5 1 1 14074
0 14076 7 4 2 48806 52918
0 14077 5 1 1 64865
0 14078 7 1 2 62631 64866
0 14079 5 1 1 14078
0 14080 7 1 2 14075 14079
0 14081 5 1 1 14080
0 14082 7 1 2 51140 14081
0 14083 5 1 1 14082
0 14084 7 1 2 50663 55055
0 14085 7 1 2 62974 14084
0 14086 5 1 1 14085
0 14087 7 1 2 45059 14086
0 14088 7 1 2 14083 14087
0 14089 7 1 2 14073 14088
0 14090 5 1 1 14089
0 14091 7 1 2 14047 14090
0 14092 5 1 1 14091
0 14093 7 1 2 13918 14092
0 14094 5 2 1 14093
0 14095 7 1 2 60892 64869
0 14096 5 1 1 14095
0 14097 7 1 2 49040 54233
0 14098 5 2 1 14097
0 14099 7 1 2 64776 64871
0 14100 5 1 1 14099
0 14101 7 1 2 48609 14100
0 14102 5 1 1 14101
0 14103 7 1 2 49041 51398
0 14104 5 2 1 14103
0 14105 7 1 2 14102 64873
0 14106 5 1 1 14105
0 14107 7 1 2 53109 14106
0 14108 5 1 1 14107
0 14109 7 1 2 51542 52863
0 14110 5 1 1 14109
0 14111 7 1 2 53503 14110
0 14112 5 1 1 14111
0 14113 7 1 2 45242 53110
0 14114 5 1 1 14113
0 14115 7 1 2 51225 52609
0 14116 5 1 1 14115
0 14117 7 3 2 49419 49616
0 14118 5 7 1 64875
0 14119 7 1 2 14116 64878
0 14120 5 1 1 14119
0 14121 7 1 2 50940 14120
0 14122 5 1 1 14121
0 14123 7 1 2 14114 14122
0 14124 7 1 2 14112 14123
0 14125 5 1 1 14124
0 14126 7 1 2 42775 14125
0 14127 5 1 1 14126
0 14128 7 1 2 53516 64879
0 14129 5 1 1 14128
0 14130 7 1 2 43893 14129
0 14131 5 1 1 14130
0 14132 7 2 2 47263 53464
0 14133 5 2 1 64885
0 14134 7 1 2 49617 64886
0 14135 5 1 1 14134
0 14136 7 1 2 14131 14135
0 14137 7 1 2 14127 14136
0 14138 5 1 1 14137
0 14139 7 1 2 53422 14138
0 14140 5 1 1 14139
0 14141 7 1 2 14108 14140
0 14142 5 1 1 14141
0 14143 7 1 2 60988 14142
0 14144 5 1 1 14143
0 14145 7 1 2 55268 60702
0 14146 5 1 1 14145
0 14147 7 1 2 2358 14146
0 14148 5 1 1 14147
0 14149 7 1 2 43289 14148
0 14150 5 1 1 14149
0 14151 7 2 2 53756 58895
0 14152 7 1 2 52610 64889
0 14153 5 1 1 14152
0 14154 7 2 2 48410 49211
0 14155 5 1 1 64891
0 14156 7 1 2 43894 64892
0 14157 5 1 1 14156
0 14158 7 1 2 14153 14157
0 14159 5 1 1 14158
0 14160 7 1 2 51194 14159
0 14161 5 1 1 14160
0 14162 7 1 2 14150 14161
0 14163 5 1 1 14162
0 14164 7 1 2 44057 14163
0 14165 5 1 1 14164
0 14166 7 3 2 48411 52959
0 14167 7 1 2 54234 64893
0 14168 5 1 1 14167
0 14169 7 2 2 49341 54262
0 14170 7 1 2 42776 64896
0 14171 5 1 1 14170
0 14172 7 1 2 14168 14171
0 14173 5 1 1 14172
0 14174 7 1 2 50840 14173
0 14175 5 1 1 14174
0 14176 7 1 2 53132 1614
0 14177 5 3 1 14176
0 14178 7 3 2 49591 58613
0 14179 5 4 1 64901
0 14180 7 1 2 64898 64902
0 14181 5 1 1 14180
0 14182 7 1 2 1677 14181
0 14183 7 1 2 14175 14182
0 14184 7 1 2 14165 14183
0 14185 5 1 1 14184
0 14186 7 1 2 48610 14185
0 14187 5 1 1 14186
0 14188 7 1 2 45060 62950
0 14189 5 1 1 14188
0 14190 7 4 2 45443 49281
0 14191 5 1 1 64908
0 14192 7 1 2 43895 14191
0 14193 7 1 2 14189 14192
0 14194 5 1 1 14193
0 14195 7 1 2 49493 14194
0 14196 5 1 1 14195
0 14197 7 1 2 42777 14196
0 14198 5 1 1 14197
0 14199 7 1 2 53111 61686
0 14200 5 1 1 14199
0 14201 7 1 2 14198 14200
0 14202 5 1 1 14201
0 14203 7 1 2 50766 14202
0 14204 5 1 1 14203
0 14205 7 1 2 14187 14204
0 14206 5 1 1 14205
0 14207 7 1 2 59221 14206
0 14208 5 1 1 14207
0 14209 7 6 2 47264 48103
0 14210 7 2 2 54959 64912
0 14211 7 1 2 55391 64918
0 14212 5 1 1 14211
0 14213 7 1 2 54547 63450
0 14214 5 1 1 14213
0 14215 7 1 2 14212 14214
0 14216 5 1 1 14215
0 14217 7 1 2 50410 14216
0 14218 5 1 1 14217
0 14219 7 5 2 42528 44757
0 14220 7 1 2 54992 64920
0 14221 7 1 2 55392 14220
0 14222 5 1 1 14221
0 14223 7 1 2 14218 14222
0 14224 5 1 1 14223
0 14225 7 1 2 49752 14224
0 14226 5 1 1 14225
0 14227 7 2 2 49042 49473
0 14228 7 1 2 58305 64925
0 14229 5 1 1 14228
0 14230 7 1 2 59896 60884
0 14231 5 2 1 14230
0 14232 7 1 2 226 64927
0 14233 5 3 1 14232
0 14234 7 1 2 54181 64929
0 14235 5 1 1 14234
0 14236 7 1 2 14229 14235
0 14237 5 1 1 14236
0 14238 7 1 2 59222 14237
0 14239 5 1 1 14238
0 14240 7 1 2 52576 55341
0 14241 7 1 2 51307 14240
0 14242 7 1 2 61499 14241
0 14243 5 1 1 14242
0 14244 7 1 2 14239 14243
0 14245 5 1 1 14244
0 14246 7 1 2 45243 14245
0 14247 5 1 1 14246
0 14248 7 1 2 14226 14247
0 14249 7 1 2 14208 14248
0 14250 5 1 1 14249
0 14251 7 1 2 47967 14250
0 14252 5 1 1 14251
0 14253 7 1 2 14144 14252
0 14254 5 2 1 14253
0 14255 7 1 2 60778 64932
0 14256 5 1 1 14255
0 14257 7 13 2 53032 5123
0 14258 5 6 1 64934
0 14259 7 1 2 53441 64935
0 14260 5 1 1 14259
0 14261 7 1 2 50238 62182
0 14262 5 1 1 14261
0 14263 7 1 2 14260 14262
0 14264 5 1 1 14263
0 14265 7 1 2 47265 14264
0 14266 5 1 1 14265
0 14267 7 1 2 50249 58034
0 14268 5 1 1 14267
0 14269 7 1 2 14266 14268
0 14270 5 1 1 14269
0 14271 7 1 2 61146 61251
0 14272 7 2 2 14270 14271
0 14273 7 1 2 60673 64953
0 14274 5 1 1 14273
0 14275 7 7 2 45716 43290
0 14276 5 2 1 64955
0 14277 7 2 2 43455 64956
0 14278 7 1 2 48412 63908
0 14279 5 1 1 14278
0 14280 7 1 2 50389 14279
0 14281 5 1 1 14280
0 14282 7 2 2 64084 14281
0 14283 7 1 2 64964 64966
0 14284 5 1 1 14283
0 14285 7 3 2 46832 64748
0 14286 7 4 2 47968 64936
0 14287 7 7 2 44758 45061
0 14288 7 1 2 61252 64975
0 14289 7 2 2 64971 14288
0 14290 7 1 2 64968 64982
0 14291 5 1 1 14290
0 14292 7 1 2 14284 14291
0 14293 5 1 1 14292
0 14294 7 1 2 43896 14293
0 14295 5 1 1 14294
0 14296 7 5 2 48104 54498
0 14297 7 2 2 56505 64984
0 14298 7 2 2 45717 51337
0 14299 7 1 2 43730 57716
0 14300 7 1 2 64991 14299
0 14301 7 1 2 64989 14300
0 14302 5 1 1 14301
0 14303 7 1 2 14295 14302
0 14304 7 1 2 14274 14303
0 14305 5 1 1 14304
0 14306 7 1 2 42529 14305
0 14307 5 1 1 14306
0 14308 7 1 2 54147 54881
0 14309 5 7 1 14308
0 14310 7 1 2 62187 64993
0 14311 5 1 1 14310
0 14312 7 1 2 55347 58565
0 14313 5 2 1 14312
0 14314 7 1 2 54263 64937
0 14315 5 1 1 14314
0 14316 7 1 2 65000 14315
0 14317 5 1 1 14316
0 14318 7 1 2 60135 14317
0 14319 5 1 1 14318
0 14320 7 1 2 14311 14319
0 14321 5 1 1 14320
0 14322 7 2 2 61673 14321
0 14323 7 1 2 60825 65002
0 14324 5 1 1 14323
0 14325 7 1 2 50455 52611
0 14326 5 3 1 14325
0 14327 7 3 2 54196 65004
0 14328 7 2 2 49753 65007
0 14329 5 1 1 65010
0 14330 7 6 2 43073 63375
0 14331 7 1 2 46014 56321
0 14332 7 1 2 65012 14331
0 14333 5 1 1 14332
0 14334 7 1 2 14329 14333
0 14335 5 1 1 14334
0 14336 7 1 2 46671 14335
0 14337 5 1 1 14336
0 14338 7 1 2 62958 64897
0 14339 5 1 1 14338
0 14340 7 1 2 14337 14339
0 14341 5 1 1 14340
0 14342 7 2 2 61674 14341
0 14343 7 1 2 60674 65018
0 14344 5 1 1 14343
0 14345 7 8 2 48611 53133
0 14346 7 3 2 50998 52577
0 14347 5 1 1 65028
0 14348 7 1 2 65020 14347
0 14349 5 1 1 14348
0 14350 7 1 2 56330 14349
0 14351 5 1 1 14350
0 14352 7 1 2 43731 14351
0 14353 5 1 1 14352
0 14354 7 3 2 52506 53476
0 14355 5 1 1 65031
0 14356 7 1 2 49440 65032
0 14357 5 1 1 14356
0 14358 7 1 2 14353 14357
0 14359 5 1 1 14358
0 14360 7 1 2 42530 14359
0 14361 5 1 1 14360
0 14362 7 1 2 56638 61706
0 14363 5 1 1 14362
0 14364 7 1 2 14361 14363
0 14365 5 1 1 14364
0 14366 7 2 2 64985 14365
0 14367 7 1 2 64965 65034
0 14368 5 1 1 14367
0 14369 7 1 2 14344 14368
0 14370 5 1 1 14369
0 14371 7 1 2 42778 14370
0 14372 5 1 1 14371
0 14373 7 1 2 14324 14372
0 14374 7 1 2 14307 14373
0 14375 5 1 1 14374
0 14376 7 1 2 49212 14375
0 14377 5 1 1 14376
0 14378 7 1 2 14256 14377
0 14379 7 1 2 14096 14378
0 14380 7 1 2 13895 14379
0 14381 5 1 1 14380
0 14382 7 1 2 47758 14381
0 14383 5 1 1 14382
0 14384 7 1 2 50072 52096
0 14385 5 1 1 14384
0 14386 7 1 2 52912 14385
0 14387 5 1 1 14386
0 14388 7 1 2 46015 14387
0 14389 5 1 1 14388
0 14390 7 1 2 42531 63498
0 14391 5 1 1 14390
0 14392 7 1 2 62117 14391
0 14393 5 1 1 14392
0 14394 7 1 2 45244 14393
0 14395 5 1 1 14394
0 14396 7 1 2 42532 50122
0 14397 5 1 1 14396
0 14398 7 1 2 14395 14397
0 14399 5 1 1 14398
0 14400 7 1 2 47421 14399
0 14401 5 1 1 14400
0 14402 7 1 2 50310 5175
0 14403 5 1 1 14402
0 14404 7 1 2 48612 14403
0 14405 5 1 1 14404
0 14406 7 1 2 55151 56738
0 14407 5 1 1 14406
0 14408 7 1 2 14405 14407
0 14409 7 1 2 14401 14408
0 14410 5 1 1 14409
0 14411 7 1 2 46225 14410
0 14412 5 1 1 14411
0 14413 7 1 2 14389 14412
0 14414 5 1 1 14413
0 14415 7 1 2 45062 14414
0 14416 5 1 1 14415
0 14417 7 3 2 52251 54033
0 14418 5 1 1 65036
0 14419 7 1 2 48413 65037
0 14420 5 1 1 14419
0 14421 7 3 2 49618 57349
0 14422 5 2 1 65039
0 14423 7 1 2 45245 53007
0 14424 5 1 1 14423
0 14425 7 1 2 65042 14424
0 14426 5 1 1 14425
0 14427 7 1 2 50999 14426
0 14428 5 1 1 14427
0 14429 7 1 2 14420 14428
0 14430 5 1 1 14429
0 14431 7 1 2 46016 14430
0 14432 5 1 1 14431
0 14433 7 1 2 49398 61480
0 14434 5 1 1 14433
0 14435 7 1 2 14432 14434
0 14436 7 1 2 14416 14435
0 14437 5 1 1 14436
0 14438 7 1 2 47266 14437
0 14439 5 1 1 14438
0 14440 7 7 2 45063 48963
0 14441 7 2 2 56779 65044
0 14442 5 1 1 65051
0 14443 7 3 2 54960 56704
0 14444 7 1 2 65052 65053
0 14445 5 1 1 14444
0 14446 7 1 2 53079 56739
0 14447 5 1 1 14446
0 14448 7 1 2 50222 58335
0 14449 5 1 1 14448
0 14450 7 1 2 14447 14449
0 14451 5 1 1 14450
0 14452 7 1 2 51000 14451
0 14453 5 1 1 14452
0 14454 7 1 2 52212 53080
0 14455 7 1 2 65038 14454
0 14456 5 1 1 14455
0 14457 7 1 2 14453 14456
0 14458 5 1 1 14457
0 14459 7 1 2 46017 14458
0 14460 5 1 1 14459
0 14461 7 1 2 14445 14460
0 14462 7 1 2 14439 14461
0 14463 5 1 1 14462
0 14464 7 1 2 61147 14463
0 14465 5 1 1 14464
0 14466 7 2 2 52823 57315
0 14467 5 1 1 65056
0 14468 7 1 2 44058 14467
0 14469 5 1 1 14468
0 14470 7 1 2 57316 64288
0 14471 5 1 1 14470
0 14472 7 1 2 48613 14471
0 14473 5 1 1 14472
0 14474 7 1 2 14469 14473
0 14475 5 1 1 14474
0 14476 7 1 2 48414 14475
0 14477 5 1 1 14476
0 14478 7 1 2 51523 53769
0 14479 5 1 1 14478
0 14480 7 2 2 49856 49975
0 14481 5 1 1 65058
0 14482 7 1 2 55242 14481
0 14483 7 1 2 14479 14482
0 14484 5 1 1 14483
0 14485 7 1 2 14477 14484
0 14486 5 1 1 14485
0 14487 7 1 2 43897 14486
0 14488 5 1 1 14487
0 14489 7 1 2 55551 3538
0 14490 5 1 1 14489
0 14491 7 1 2 48415 57997
0 14492 7 2 2 14490 14491
0 14493 5 1 1 65060
0 14494 7 1 2 57548 65061
0 14495 5 1 1 14494
0 14496 7 1 2 14488 14495
0 14497 5 1 1 14496
0 14498 7 1 2 63244 14497
0 14499 5 1 1 14498
0 14500 7 1 2 51203 52668
0 14501 7 1 2 58542 61071
0 14502 7 1 2 14500 14501
0 14503 5 1 1 14502
0 14504 7 1 2 14493 14503
0 14505 5 1 1 14504
0 14506 7 1 2 48614 14505
0 14507 5 1 1 14506
0 14508 7 1 2 53458 58660
0 14509 7 1 2 65057 14508
0 14510 5 1 1 14509
0 14511 7 1 2 53504 14510
0 14512 5 1 1 14511
0 14513 7 1 2 14507 14512
0 14514 5 1 1 14513
0 14515 7 1 2 42533 14514
0 14516 5 1 1 14515
0 14517 7 1 2 55552 60732
0 14518 5 1 1 14517
0 14519 7 1 2 53112 57998
0 14520 7 1 2 63868 14519
0 14521 7 1 2 14518 14520
0 14522 5 1 1 14521
0 14523 7 1 2 14516 14522
0 14524 5 1 1 14523
0 14525 7 1 2 60396 14524
0 14526 5 1 1 14525
0 14527 7 5 2 53525 62364
0 14528 7 4 2 44202 60397
0 14529 7 1 2 49857 65067
0 14530 7 1 2 65062 14529
0 14531 5 1 1 14530
0 14532 7 1 2 47969 53396
0 14533 7 1 2 60084 14532
0 14534 7 1 2 62332 14533
0 14535 5 1 1 14534
0 14536 7 1 2 14531 14535
0 14537 5 1 1 14536
0 14538 7 1 2 45444 14537
0 14539 5 1 1 14538
0 14540 7 3 2 47970 64976
0 14541 7 1 2 55039 65071
0 14542 5 1 1 14541
0 14543 7 10 2 44642 48416
0 14544 7 2 2 43898 65074
0 14545 7 1 2 42534 48105
0 14546 7 2 2 65084 14545
0 14547 5 1 1 65086
0 14548 7 1 2 14542 14547
0 14549 5 1 1 14548
0 14550 7 1 2 52252 14549
0 14551 5 1 1 14550
0 14552 7 1 2 14539 14551
0 14553 7 1 2 14526 14552
0 14554 5 1 1 14553
0 14555 7 1 2 42779 14554
0 14556 5 1 1 14555
0 14557 7 1 2 14499 14556
0 14558 7 1 2 14465 14557
0 14559 5 1 1 14558
0 14560 7 1 2 43732 14559
0 14561 5 1 1 14560
0 14562 7 1 2 60291 62147
0 14563 5 1 1 14562
0 14564 7 1 2 58475 12346
0 14565 5 1 1 14564
0 14566 7 1 2 50941 14565
0 14567 5 1 1 14566
0 14568 7 1 2 42535 52993
0 14569 5 1 1 14568
0 14570 7 1 2 56622 14569
0 14571 7 1 2 14567 14570
0 14572 5 1 1 14571
0 14573 7 1 2 44203 14572
0 14574 5 1 1 14573
0 14575 7 1 2 14563 14574
0 14576 5 1 1 14575
0 14577 7 1 2 43291 14576
0 14578 5 1 1 14577
0 14579 7 2 2 54309 60703
0 14580 5 1 1 65088
0 14581 7 1 2 49468 14580
0 14582 5 1 1 14581
0 14583 7 1 2 47267 14582
0 14584 5 1 1 14583
0 14585 7 1 2 52960 60730
0 14586 5 1 1 14585
0 14587 7 1 2 14584 14586
0 14588 5 1 1 14587
0 14589 7 1 2 46672 14588
0 14590 5 1 1 14589
0 14591 7 1 2 49465 53397
0 14592 5 1 1 14591
0 14593 7 1 2 14590 14592
0 14594 7 1 2 14578 14593
0 14595 5 1 1 14594
0 14596 7 1 2 48615 14595
0 14597 5 1 1 14596
0 14598 7 1 2 62145 63930
0 14599 5 1 1 14598
0 14600 7 1 2 50073 14599
0 14601 5 1 1 14600
0 14602 7 1 2 47268 63504
0 14603 5 1 1 14602
0 14604 7 1 2 56152 14603
0 14605 5 1 1 14604
0 14606 7 1 2 45246 14605
0 14607 5 1 1 14606
0 14608 7 1 2 14601 14607
0 14609 5 1 1 14608
0 14610 7 1 2 42536 14609
0 14611 5 1 1 14610
0 14612 7 1 2 50553 56339
0 14613 7 1 2 58370 14612
0 14614 5 1 1 14613
0 14615 7 1 2 14611 14614
0 14616 7 1 2 14597 14615
0 14617 5 1 1 14616
0 14618 7 1 2 47102 14617
0 14619 5 1 1 14618
0 14620 7 1 2 42537 58332
0 14621 5 1 1 14620
0 14622 7 1 2 59774 62372
0 14623 5 1 1 14622
0 14624 7 1 2 14621 14623
0 14625 5 1 1 14624
0 14626 7 1 2 46226 14625
0 14627 5 1 1 14626
0 14628 7 2 2 46018 58344
0 14629 5 1 1 65090
0 14630 7 1 2 42780 65091
0 14631 7 1 2 58102 14630
0 14632 5 1 1 14631
0 14633 7 1 2 14627 14632
0 14634 5 1 1 14633
0 14635 7 1 2 43074 14634
0 14636 5 1 1 14635
0 14637 7 2 2 49159 54863
0 14638 7 1 2 58324 65092
0 14639 5 1 1 14638
0 14640 7 1 2 14636 14639
0 14641 7 1 2 14619 14640
0 14642 5 1 1 14641
0 14643 7 1 2 44759 14642
0 14644 5 1 1 14643
0 14645 7 1 2 47269 52422
0 14646 5 1 1 14645
0 14647 7 1 2 57578 61906
0 14648 5 1 1 14647
0 14649 7 1 2 47270 52410
0 14650 7 1 2 57879 14649
0 14651 5 1 1 14650
0 14652 7 1 2 14648 14651
0 14653 5 1 1 14652
0 14654 7 1 2 46483 14653
0 14655 5 1 1 14654
0 14656 7 1 2 14646 14655
0 14657 5 1 1 14656
0 14658 7 1 2 46227 14657
0 14659 5 1 1 14658
0 14660 7 1 2 52979 62971
0 14661 5 1 1 14660
0 14662 7 1 2 14659 14661
0 14663 5 1 1 14662
0 14664 7 1 2 51296 14663
0 14665 5 1 1 14664
0 14666 7 1 2 14644 14665
0 14667 5 1 1 14666
0 14668 7 1 2 45064 14667
0 14669 5 1 1 14668
0 14670 7 2 2 51882 59183
0 14671 5 2 1 65094
0 14672 7 1 2 56618 65096
0 14673 5 1 1 14672
0 14674 7 1 2 56374 57828
0 14675 5 1 1 14674
0 14676 7 1 2 14673 14675
0 14677 5 1 1 14676
0 14678 7 1 2 48616 14677
0 14679 5 1 1 14678
0 14680 7 1 2 49976 59508
0 14681 5 1 1 14680
0 14682 7 1 2 58661 14681
0 14683 5 1 1 14682
0 14684 7 1 2 56619 14683
0 14685 5 1 1 14684
0 14686 7 1 2 14679 14685
0 14687 5 1 1 14686
0 14688 7 1 2 57855 14687
0 14689 5 1 1 14688
0 14690 7 1 2 14669 14689
0 14691 5 1 1 14690
0 14692 7 1 2 47971 14691
0 14693 5 1 1 14692
0 14694 7 1 2 50456 3650
0 14695 5 1 1 14694
0 14696 7 1 2 62810 14695
0 14697 5 1 1 14696
0 14698 7 2 2 47103 52749
0 14699 7 1 2 57654 65098
0 14700 5 1 1 14699
0 14701 7 1 2 14697 14700
0 14702 5 1 1 14701
0 14703 7 1 2 62326 14702
0 14704 5 1 1 14703
0 14705 7 1 2 49213 5795
0 14706 7 1 2 62264 14705
0 14707 5 1 1 14706
0 14708 7 1 2 14704 14707
0 14709 5 1 1 14708
0 14710 7 1 2 42781 14709
0 14711 5 1 1 14710
0 14712 7 1 2 50411 53489
0 14713 5 1 1 14712
0 14714 7 1 2 43733 14629
0 14715 5 2 1 14714
0 14716 7 1 2 57187 60734
0 14717 7 1 2 65100 14716
0 14718 5 1 1 14717
0 14719 7 1 2 14713 14718
0 14720 5 1 1 14719
0 14721 7 1 2 61148 14720
0 14722 5 1 1 14721
0 14723 7 1 2 14711 14722
0 14724 5 1 1 14723
0 14725 7 1 2 43292 14724
0 14726 5 1 1 14725
0 14727 7 1 2 49043 64474
0 14728 5 1 1 14727
0 14729 7 1 2 64286 14728
0 14730 5 1 1 14729
0 14731 7 1 2 46673 14730
0 14732 5 1 1 14731
0 14733 7 1 2 53385 62155
0 14734 5 1 1 14733
0 14735 7 1 2 14732 14734
0 14736 5 1 1 14735
0 14737 7 1 2 61519 14736
0 14738 5 1 1 14737
0 14739 7 1 2 52381 61341
0 14740 7 1 2 62453 14739
0 14741 7 1 2 65068 14740
0 14742 5 1 1 14741
0 14743 7 1 2 14738 14742
0 14744 7 1 2 14726 14743
0 14745 5 1 1 14744
0 14746 7 1 2 43075 14745
0 14747 5 1 1 14746
0 14748 7 1 2 49160 64359
0 14749 5 1 1 14748
0 14750 7 1 2 49754 62110
0 14751 5 1 1 14750
0 14752 7 1 2 14749 14751
0 14753 5 1 1 14752
0 14754 7 1 2 46674 14753
0 14755 5 1 1 14754
0 14756 7 1 2 62111 64811
0 14757 5 1 1 14756
0 14758 7 2 2 52247 56635
0 14759 5 1 1 65102
0 14760 7 1 2 14757 14759
0 14761 7 1 2 14755 14760
0 14762 5 1 1 14761
0 14763 7 1 2 46484 14762
0 14764 5 1 1 14763
0 14765 7 1 2 50074 53390
0 14766 5 1 1 14765
0 14767 7 1 2 64294 14766
0 14768 5 1 1 14767
0 14769 7 1 2 42538 14768
0 14770 5 1 1 14769
0 14771 7 1 2 47271 56851
0 14772 5 1 1 14771
0 14773 7 1 2 53477 56841
0 14774 5 1 1 14773
0 14775 7 1 2 46228 14774
0 14776 5 1 1 14775
0 14777 7 1 2 50192 58485
0 14778 7 1 2 60895 14777
0 14779 5 1 1 14778
0 14780 7 1 2 46019 14779
0 14781 7 1 2 14776 14780
0 14782 7 1 2 14772 14781
0 14783 5 1 1 14782
0 14784 7 1 2 14770 14783
0 14785 7 1 2 14764 14784
0 14786 5 1 1 14785
0 14787 7 1 2 47104 14786
0 14788 5 1 1 14787
0 14789 7 1 2 50918 57372
0 14790 7 1 2 64360 14789
0 14791 5 1 1 14790
0 14792 7 1 2 14788 14791
0 14793 5 1 1 14792
0 14794 7 1 2 61149 14793
0 14795 5 1 1 14794
0 14796 7 1 2 14747 14795
0 14797 5 1 1 14796
0 14798 7 1 2 48417 14797
0 14799 5 1 1 14798
0 14800 7 1 2 14693 14799
0 14801 7 1 2 14561 14800
0 14802 5 1 1 14801
0 14803 7 1 2 51857 55897
0 14804 7 1 2 14802 14803
0 14805 5 1 1 14804
0 14806 7 1 2 14383 14805
0 14807 5 1 1 14806
0 14808 7 1 2 42013 14807
0 14809 5 1 1 14808
0 14810 7 1 2 60740 62254
0 14811 5 1 1 14810
0 14812 7 1 2 49596 59077
0 14813 5 2 1 14812
0 14814 7 1 2 57839 65104
0 14815 5 1 1 14814
0 14816 7 2 2 49455 58788
0 14817 5 1 1 65106
0 14818 7 1 2 14815 14817
0 14819 7 1 2 14811 14818
0 14820 5 1 1 14819
0 14821 7 1 2 48617 14820
0 14822 5 1 1 14821
0 14823 7 1 2 44204 50156
0 14824 7 1 2 52832 14823
0 14825 5 1 1 14824
0 14826 7 1 2 14822 14825
0 14827 5 1 1 14826
0 14828 7 1 2 48418 14827
0 14829 5 1 1 14828
0 14830 7 1 2 50239 53840
0 14831 5 1 1 14830
0 14832 7 1 2 14829 14831
0 14833 5 1 1 14832
0 14834 7 1 2 43899 14833
0 14835 5 1 1 14834
0 14836 7 1 2 48419 60741
0 14837 5 1 1 14836
0 14838 7 1 2 53014 14837
0 14839 5 1 1 14838
0 14840 7 1 2 43076 14839
0 14841 5 1 1 14840
0 14842 7 2 2 46675 52612
0 14843 5 1 1 65108
0 14844 7 1 2 44205 14843
0 14845 5 1 1 14844
0 14846 7 1 2 47543 4867
0 14847 5 2 1 14846
0 14848 7 1 2 45445 65110
0 14849 7 1 2 14845 14848
0 14850 5 1 1 14849
0 14851 7 1 2 48618 55272
0 14852 7 1 2 14850 14851
0 14853 7 1 2 14841 14852
0 14854 5 1 1 14853
0 14855 7 1 2 45247 53531
0 14856 7 1 2 6815 14855
0 14857 5 1 1 14856
0 14858 7 1 2 14854 14857
0 14859 5 1 1 14858
0 14860 7 1 2 47272 1314
0 14861 5 2 1 14860
0 14862 7 3 2 46485 53134
0 14863 5 1 1 65114
0 14864 7 1 2 60742 14863
0 14865 7 1 2 65112 14864
0 14866 5 1 1 14865
0 14867 7 1 2 14859 14866
0 14868 5 1 1 14867
0 14869 7 1 2 44059 14868
0 14870 5 1 1 14869
0 14871 7 4 2 44206 45065
0 14872 5 1 1 65117
0 14873 7 1 2 55296 14872
0 14874 5 1 1 14873
0 14875 7 1 2 43077 14874
0 14876 5 1 1 14875
0 14877 7 1 2 48420 58444
0 14878 5 1 1 14877
0 14879 7 1 2 43293 14878
0 14880 7 1 2 14876 14879
0 14881 5 1 1 14880
0 14882 7 1 2 48421 58575
0 14883 5 2 1 14882
0 14884 7 1 2 44207 52724
0 14885 5 1 1 14884
0 14886 7 1 2 65121 14885
0 14887 5 1 1 14886
0 14888 7 1 2 45446 14887
0 14889 5 1 1 14888
0 14890 7 1 2 47422 53465
0 14891 5 1 1 14890
0 14892 7 1 2 46676 14891
0 14893 7 1 2 14889 14892
0 14894 5 1 1 14893
0 14895 7 1 2 14881 14894
0 14896 5 1 1 14895
0 14897 7 5 2 45066 52382
0 14898 7 1 2 50128 65123
0 14899 5 1 1 14898
0 14900 7 1 2 62365 65118
0 14901 5 3 1 14900
0 14902 7 1 2 14899 65128
0 14903 7 1 2 14896 14902
0 14904 5 1 1 14903
0 14905 7 1 2 43900 14904
0 14906 5 1 1 14905
0 14907 7 1 2 49000 50157
0 14908 7 1 2 53541 14907
0 14909 5 1 1 14908
0 14910 7 1 2 14906 14909
0 14911 7 1 2 14870 14910
0 14912 5 1 1 14911
0 14913 7 1 2 42782 14912
0 14914 5 1 1 14913
0 14915 7 1 2 14835 14914
0 14916 5 1 1 14915
0 14917 7 1 2 43734 14916
0 14918 5 1 1 14917
0 14919 7 1 2 54364 14918
0 14920 5 1 1 14919
0 14921 7 1 2 60398 14920
0 14922 5 1 1 14921
0 14923 7 1 2 55112 62975
0 14924 5 1 1 14923
0 14925 7 3 2 53946 57760
0 14926 5 1 1 65131
0 14927 7 1 2 54961 65021
0 14928 5 1 1 14927
0 14929 7 1 2 14926 14928
0 14930 5 1 1 14929
0 14931 7 1 2 49044 14930
0 14932 5 1 1 14931
0 14933 7 2 2 49564 55520
0 14934 5 1 1 65134
0 14935 7 1 2 14932 14934
0 14936 5 1 1 14935
0 14937 7 1 2 47423 14936
0 14938 5 1 1 14937
0 14939 7 1 2 52578 64365
0 14940 5 1 1 14939
0 14941 7 1 2 65001 14940
0 14942 5 1 1 14941
0 14943 7 1 2 49081 14942
0 14944 5 1 1 14943
0 14945 7 1 2 49429 63241
0 14946 5 1 1 14945
0 14947 7 1 2 43294 14946
0 14948 7 1 2 14944 14947
0 14949 7 1 2 14938 14948
0 14950 5 1 1 14949
0 14951 7 1 2 49214 64366
0 14952 5 2 1 14951
0 14953 7 1 2 49161 64947
0 14954 5 2 1 14953
0 14955 7 1 2 65136 65138
0 14956 5 1 1 14955
0 14957 7 2 2 45067 14956
0 14958 5 1 1 65140
0 14959 7 1 2 47273 65141
0 14960 5 1 1 14959
0 14961 7 1 2 55323 58505
0 14962 7 2 2 63266 14961
0 14963 7 1 2 45248 65142
0 14964 5 1 1 14963
0 14965 7 1 2 61935 14964
0 14966 5 1 1 14965
0 14967 7 1 2 53069 14966
0 14968 5 1 1 14967
0 14969 7 1 2 46677 14968
0 14970 7 1 2 14960 14969
0 14971 5 1 1 14970
0 14972 7 1 2 14950 14971
0 14973 5 1 1 14972
0 14974 7 1 2 62892 65119
0 14975 5 1 1 14974
0 14976 7 2 2 43295 52071
0 14977 5 1 1 65144
0 14978 7 1 2 60250 14977
0 14979 5 1 1 14978
0 14980 7 1 2 46229 14979
0 14981 5 1 1 14980
0 14982 7 1 2 59086 64938
0 14983 5 1 1 14982
0 14984 7 2 2 54987 57373
0 14985 5 1 1 65146
0 14986 7 1 2 50554 65147
0 14987 5 1 1 14986
0 14988 7 1 2 14983 14987
0 14989 7 1 2 14981 14988
0 14990 5 1 1 14989
0 14991 7 1 2 54264 14990
0 14992 5 1 1 14991
0 14993 7 1 2 14975 14992
0 14994 7 1 2 14973 14993
0 14995 5 1 1 14994
0 14996 7 1 2 47105 14995
0 14997 5 1 1 14996
0 14998 7 1 2 14924 14997
0 14999 5 1 1 14998
0 15000 7 1 2 61150 14999
0 15001 5 1 1 15000
0 15002 7 1 2 14922 15001
0 15003 5 1 1 15002
0 15004 7 1 2 42539 15003
0 15005 5 1 1 15004
0 15006 7 1 2 43901 53880
0 15007 5 1 1 15006
0 15008 7 1 2 42783 53135
0 15009 7 1 2 50322 15008
0 15010 5 1 1 15009
0 15011 7 1 2 15007 15010
0 15012 5 1 1 15011
0 15013 7 1 2 47106 15012
0 15014 5 1 1 15013
0 15015 7 1 2 49565 62168
0 15016 5 2 1 15015
0 15017 7 1 2 15014 65148
0 15018 5 1 1 15017
0 15019 7 1 2 43078 15018
0 15020 5 1 1 15019
0 15021 7 1 2 54310 55049
0 15022 5 1 1 15021
0 15023 7 1 2 44060 64994
0 15024 5 1 1 15023
0 15025 7 1 2 51503 53136
0 15026 7 1 2 54135 15025
0 15027 5 1 1 15026
0 15028 7 1 2 15024 15027
0 15029 5 1 1 15028
0 15030 7 1 2 46230 15029
0 15031 5 1 1 15030
0 15032 7 1 2 15022 15031
0 15033 7 1 2 15020 15032
0 15034 5 1 1 15033
0 15035 7 1 2 49045 15034
0 15036 5 1 1 15035
0 15037 7 3 2 54265 55102
0 15038 5 1 1 65150
0 15039 7 1 2 46486 65151
0 15040 5 1 1 15039
0 15041 7 1 2 44061 15040
0 15042 5 1 1 15041
0 15043 7 1 2 42784 64995
0 15044 5 1 1 15043
0 15045 7 1 2 15044 15038
0 15046 5 2 1 15045
0 15047 7 1 2 45249 65153
0 15048 7 1 2 15042 15047
0 15049 5 1 1 15048
0 15050 7 1 2 15036 15049
0 15051 5 1 1 15050
0 15052 7 1 2 43296 15051
0 15053 5 1 1 15052
0 15054 7 2 2 42785 54266
0 15055 5 1 1 65155
0 15056 7 5 2 46231 53113
0 15057 5 1 1 65157
0 15058 7 1 2 15055 15057
0 15059 5 5 1 15058
0 15060 7 1 2 47107 65162
0 15061 5 1 1 15060
0 15062 7 1 2 2184 15061
0 15063 5 2 1 15062
0 15064 7 2 2 44062 65167
0 15065 5 1 1 65169
0 15066 7 1 2 52507 65156
0 15067 5 1 1 15066
0 15068 7 1 2 15065 15067
0 15069 5 1 1 15068
0 15070 7 1 2 49619 15069
0 15071 5 1 1 15070
0 15072 7 1 2 15053 15071
0 15073 5 1 1 15072
0 15074 7 1 2 44760 15073
0 15075 5 1 1 15074
0 15076 7 1 2 49162 62176
0 15077 5 1 1 15076
0 15078 7 1 2 49215 64948
0 15079 5 1 1 15078
0 15080 7 1 2 48422 15079
0 15081 7 1 2 15077 15080
0 15082 5 1 1 15081
0 15083 7 1 2 14958 15082
0 15084 5 1 1 15083
0 15085 7 1 2 57195 15084
0 15086 5 1 1 15085
0 15087 7 9 2 48106 45068
0 15088 7 2 2 54096 65171
0 15089 7 1 2 53832 65180
0 15090 5 1 1 15089
0 15091 7 1 2 15086 15090
0 15092 5 1 1 15091
0 15093 7 1 2 47274 15092
0 15094 5 1 1 15093
0 15095 7 3 2 43735 52613
0 15096 5 1 1 65182
0 15097 7 1 2 52217 65183
0 15098 5 1 1 15097
0 15099 7 1 2 52688 54844
0 15100 5 1 1 15099
0 15101 7 1 2 15098 15100
0 15102 5 1 1 15101
0 15103 7 1 2 56766 15102
0 15104 5 1 1 15103
0 15105 7 1 2 51463 53423
0 15106 5 1 1 15105
0 15107 7 1 2 49216 15106
0 15108 5 1 1 15107
0 15109 7 1 2 49163 1651
0 15110 7 1 2 10043 15109
0 15111 7 1 2 7920 15110
0 15112 5 1 1 15111
0 15113 7 1 2 15108 15112
0 15114 5 1 1 15113
0 15115 7 1 2 55648 15114
0 15116 5 1 1 15115
0 15117 7 1 2 47108 64158
0 15118 5 1 1 15117
0 15119 7 1 2 52072 55103
0 15120 5 1 1 15119
0 15121 7 1 2 49164 15120
0 15122 7 1 2 15118 15121
0 15123 5 1 1 15122
0 15124 7 1 2 47109 55989
0 15125 5 1 1 15124
0 15126 7 1 2 49217 15125
0 15127 5 1 1 15126
0 15128 7 1 2 48423 15127
0 15129 7 1 2 15123 15128
0 15130 5 1 1 15129
0 15131 7 1 2 15116 15130
0 15132 5 1 1 15131
0 15133 7 1 2 43902 15132
0 15134 5 1 1 15133
0 15135 7 1 2 15104 15134
0 15136 5 1 1 15135
0 15137 7 1 2 44761 15136
0 15138 5 1 1 15137
0 15139 7 1 2 15094 15138
0 15140 5 1 1 15139
0 15141 7 1 2 46678 15140
0 15142 5 1 1 15141
0 15143 7 2 2 49282 52268
0 15144 7 2 2 54571 65185
0 15145 5 1 1 65187
0 15146 7 1 2 47110 65188
0 15147 5 1 1 15146
0 15148 7 1 2 54034 54267
0 15149 5 1 1 15148
0 15150 7 1 2 54695 54962
0 15151 5 2 1 15150
0 15152 7 1 2 15149 65189
0 15153 5 1 1 15152
0 15154 7 1 2 43736 15153
0 15155 5 1 1 15154
0 15156 7 1 2 47111 52692
0 15157 5 1 1 15156
0 15158 7 1 2 42786 15096
0 15159 7 1 2 15157 15158
0 15160 5 1 1 15159
0 15161 7 1 2 15155 15160
0 15162 5 1 1 15161
0 15163 7 1 2 45250 15162
0 15164 5 1 1 15163
0 15165 7 1 2 55990 64996
0 15166 5 1 1 15165
0 15167 7 1 2 51001 65152
0 15168 5 1 1 15167
0 15169 7 1 2 15166 15168
0 15170 7 1 2 15164 15169
0 15171 5 1 1 15170
0 15172 7 1 2 58095 15171
0 15173 5 1 1 15172
0 15174 7 1 2 15147 15173
0 15175 5 1 1 15174
0 15176 7 1 2 49082 15175
0 15177 5 1 1 15176
0 15178 7 1 2 15142 15177
0 15179 7 1 2 15075 15178
0 15180 5 1 1 15179
0 15181 7 1 2 47972 15180
0 15182 5 1 1 15181
0 15183 7 2 2 53114 61728
0 15184 5 2 1 65191
0 15185 7 3 2 51338 54311
0 15186 7 1 2 52405 65195
0 15187 7 1 2 65192 15186
0 15188 5 1 1 15187
0 15189 7 1 2 15182 15188
0 15190 5 1 1 15189
0 15191 7 1 2 46020 15190
0 15192 5 1 1 15191
0 15193 7 1 2 48424 64842
0 15194 5 1 1 15193
0 15195 7 2 2 50223 61151
0 15196 7 1 2 55089 65198
0 15197 5 1 1 15196
0 15198 7 1 2 15194 15197
0 15199 5 1 1 15198
0 15200 7 3 2 44063 60747
0 15201 5 1 1 65200
0 15202 7 1 2 52309 15201
0 15203 5 2 1 15202
0 15204 7 1 2 15199 65203
0 15205 5 1 1 15204
0 15206 7 1 2 60989 64844
0 15207 5 1 1 15206
0 15208 7 2 2 46021 52508
0 15209 7 1 2 55488 57978
0 15210 7 1 2 65205 15209
0 15211 5 1 1 15210
0 15212 7 1 2 15207 15211
0 15213 5 1 1 15212
0 15214 7 1 2 48425 15213
0 15215 5 1 1 15214
0 15216 7 1 2 46022 64677
0 15217 7 1 2 65199 15216
0 15218 5 1 1 15217
0 15219 7 1 2 15215 15218
0 15220 5 1 1 15219
0 15221 7 1 2 60748 63524
0 15222 7 1 2 15220 15221
0 15223 5 1 1 15222
0 15224 7 1 2 15205 15223
0 15225 7 1 2 15192 15224
0 15226 7 1 2 15005 15225
0 15227 5 1 1 15226
0 15228 7 3 2 43456 61019
0 15229 7 1 2 57027 65207
0 15230 7 1 2 15227 15229
0 15231 5 1 1 15230
0 15232 7 1 2 14809 15231
0 15233 5 1 1 15232
0 15234 7 1 2 62685 15233
0 15235 5 1 1 15234
0 15236 7 1 2 42540 52701
0 15237 5 1 1 15236
0 15238 7 1 2 52833 55521
0 15239 7 1 2 57761 15238
0 15240 5 1 1 15239
0 15241 7 1 2 15237 15240
0 15242 5 1 1 15241
0 15243 7 1 2 47112 15242
0 15244 5 1 1 15243
0 15245 7 1 2 43737 52994
0 15246 5 1 1 15245
0 15247 7 1 2 43738 58973
0 15248 5 1 1 15247
0 15249 7 1 2 54243 15248
0 15250 5 1 1 15249
0 15251 7 1 2 15246 15250
0 15252 5 1 1 15251
0 15253 7 1 2 45069 15252
0 15254 5 1 1 15253
0 15255 7 1 2 54882 55074
0 15256 5 1 1 15255
0 15257 7 1 2 46487 15256
0 15258 5 1 1 15257
0 15259 7 1 2 54883 8945
0 15260 5 1 1 15259
0 15261 7 1 2 46232 15260
0 15262 5 1 1 15261
0 15263 7 2 2 52870 54003
0 15264 5 1 1 65210
0 15265 7 1 2 15262 15264
0 15266 7 1 2 15258 15265
0 15267 7 1 2 15254 15266
0 15268 5 1 1 15267
0 15269 7 1 2 46023 15268
0 15270 5 1 1 15269
0 15271 7 1 2 15244 15270
0 15272 5 1 1 15271
0 15273 7 1 2 44208 15272
0 15274 5 1 1 15273
0 15275 7 1 2 50457 57085
0 15276 5 1 1 15275
0 15277 7 1 2 62811 15276
0 15278 5 1 1 15277
0 15279 7 1 2 54097 57655
0 15280 5 1 1 15279
0 15281 7 1 2 15278 15280
0 15282 5 1 1 15281
0 15283 7 1 2 50942 15282
0 15284 5 1 1 15283
0 15285 7 5 2 47113 54386
0 15286 7 1 2 44209 65212
0 15287 5 1 1 15286
0 15288 7 1 2 15284 15287
0 15289 5 1 1 15288
0 15290 7 1 2 54268 15289
0 15291 5 1 1 15290
0 15292 7 1 2 49513 55269
0 15293 7 1 2 64137 15292
0 15294 5 1 1 15293
0 15295 7 1 2 15291 15294
0 15296 7 1 2 15274 15295
0 15297 5 1 1 15296
0 15298 7 1 2 43297 15297
0 15299 5 1 1 15298
0 15300 7 1 2 55250 62583
0 15301 5 1 1 15300
0 15302 7 2 2 49420 55231
0 15303 5 1 1 65217
0 15304 7 1 2 60896 65218
0 15305 5 1 1 15304
0 15306 7 1 2 15301 15305
0 15307 5 1 1 15306
0 15308 7 1 2 47114 15307
0 15309 5 1 1 15308
0 15310 7 4 2 42787 51172
0 15311 7 1 2 50305 65219
0 15312 5 1 1 15311
0 15313 7 3 2 47115 49046
0 15314 7 2 2 56211 65223
0 15315 5 1 1 65226
0 15316 7 1 2 15312 15315
0 15317 5 1 1 15316
0 15318 7 1 2 54269 15317
0 15319 5 1 1 15318
0 15320 7 2 2 54251 3564
0 15321 7 2 2 49165 54963
0 15322 5 1 1 65230
0 15323 7 1 2 6773 65231
0 15324 7 1 2 65228 15323
0 15325 5 1 1 15324
0 15326 7 1 2 15319 15325
0 15327 7 1 2 15309 15326
0 15328 5 1 1 15327
0 15329 7 1 2 49123 15328
0 15330 5 1 1 15329
0 15331 7 1 2 46024 64899
0 15332 5 2 1 15331
0 15333 7 1 2 53213 65232
0 15334 5 1 1 15333
0 15335 7 1 2 65005 65097
0 15336 7 1 2 15334 15335
0 15337 5 1 1 15336
0 15338 7 1 2 15330 15337
0 15339 7 1 2 15299 15338
0 15340 5 1 1 15339
0 15341 7 1 2 51926 15340
0 15342 5 1 1 15341
0 15343 7 1 2 46233 54270
0 15344 5 1 1 15343
0 15345 7 2 2 42788 52579
0 15346 5 2 1 65234
0 15347 7 1 2 15344 65236
0 15348 5 2 1 15347
0 15349 7 1 2 50943 65238
0 15350 5 1 1 15349
0 15351 7 1 2 55027 65233
0 15352 7 1 2 15350 15351
0 15353 5 1 1 15352
0 15354 7 1 2 47116 15353
0 15355 5 1 1 15354
0 15356 7 1 2 46025 54143
0 15357 5 1 1 15356
0 15358 7 1 2 15355 15357
0 15359 5 1 1 15358
0 15360 7 1 2 59087 15359
0 15361 5 1 1 15360
0 15362 7 1 2 51058 65239
0 15363 5 1 1 15362
0 15364 7 1 2 53075 2014
0 15365 7 1 2 60268 15364
0 15366 5 1 1 15365
0 15367 7 1 2 47275 1794
0 15368 5 1 1 15367
0 15369 7 1 2 48426 15368
0 15370 5 1 1 15369
0 15371 7 1 2 46026 61709
0 15372 7 1 2 15370 15371
0 15373 7 1 2 15366 15372
0 15374 5 1 1 15373
0 15375 7 1 2 15363 15374
0 15376 5 1 1 15375
0 15377 7 1 2 52295 15376
0 15378 5 1 1 15377
0 15379 7 2 2 54271 60721
0 15380 7 1 2 51173 65240
0 15381 5 1 1 15380
0 15382 7 1 2 50412 52614
0 15383 5 1 1 15382
0 15384 7 1 2 15381 15383
0 15385 5 1 1 15384
0 15386 7 1 2 42789 15385
0 15387 5 1 1 15386
0 15388 7 1 2 42541 15322
0 15389 5 1 1 15388
0 15390 7 1 2 64997 15389
0 15391 5 1 1 15390
0 15392 7 1 2 55311 58409
0 15393 5 1 1 15392
0 15394 7 1 2 54671 15393
0 15395 7 1 2 15391 15394
0 15396 7 1 2 15387 15395
0 15397 5 1 1 15396
0 15398 7 1 2 46679 15397
0 15399 5 1 1 15398
0 15400 7 1 2 15378 15399
0 15401 5 1 1 15400
0 15402 7 1 2 44064 15401
0 15403 5 1 1 15402
0 15404 7 1 2 15361 15403
0 15405 5 1 1 15404
0 15406 7 1 2 59276 15405
0 15407 5 1 1 15406
0 15408 7 1 2 15342 15407
0 15409 5 1 1 15408
0 15410 7 1 2 61152 15409
0 15411 5 1 1 15410
0 15412 7 1 2 42542 54235
0 15413 5 1 1 15412
0 15414 7 1 2 45447 55127
0 15415 5 1 1 15414
0 15416 7 1 2 15413 15415
0 15417 5 1 1 15416
0 15418 7 1 2 51927 15417
0 15419 5 1 1 15418
0 15420 7 1 2 44065 63934
0 15421 7 1 2 62819 15420
0 15422 5 1 1 15421
0 15423 7 1 2 15419 15422
0 15424 5 1 1 15423
0 15425 7 1 2 44210 15424
0 15426 5 1 1 15425
0 15427 7 1 2 46027 55133
0 15428 5 2 1 15427
0 15429 7 1 2 62826 65242
0 15430 5 1 1 15429
0 15431 7 1 2 15426 15430
0 15432 5 1 1 15431
0 15433 7 1 2 43298 15432
0 15434 5 1 1 15433
0 15435 7 1 2 51928 58449
0 15436 5 1 1 15435
0 15437 7 1 2 12247 15436
0 15438 5 1 1 15437
0 15439 7 1 2 46680 15438
0 15440 5 1 1 15439
0 15441 7 1 2 49342 64762
0 15442 5 1 1 15441
0 15443 7 2 2 64732 15442
0 15444 5 1 1 65244
0 15445 7 1 2 15440 65245
0 15446 5 1 1 15445
0 15447 7 1 2 42543 15446
0 15448 5 1 1 15447
0 15449 7 1 2 44066 55377
0 15450 7 1 2 62788 15449
0 15451 5 1 1 15450
0 15452 7 1 2 15448 15451
0 15453 7 1 2 15434 15452
0 15454 5 1 1 15453
0 15455 7 1 2 48427 15454
0 15456 5 1 1 15455
0 15457 7 1 2 45070 49977
0 15458 5 1 1 15457
0 15459 7 1 2 49126 15458
0 15460 5 1 1 15459
0 15461 7 6 2 42790 51929
0 15462 5 1 1 65246
0 15463 7 4 2 42169 43079
0 15464 7 1 2 57783 65252
0 15465 5 2 1 15464
0 15466 7 1 2 15462 65256
0 15467 5 2 1 15466
0 15468 7 1 2 15460 65258
0 15469 5 1 1 15468
0 15470 7 1 2 42791 15444
0 15471 5 1 1 15470
0 15472 7 1 2 59323 10077
0 15473 5 5 1 15472
0 15474 7 1 2 55577 65260
0 15475 5 2 1 15474
0 15476 7 1 2 43299 63132
0 15477 5 1 1 15476
0 15478 7 1 2 65265 15477
0 15479 7 1 2 15471 15478
0 15480 5 1 1 15479
0 15481 7 1 2 53424 15480
0 15482 5 2 1 15481
0 15483 7 1 2 15469 65267
0 15484 5 1 1 15483
0 15485 7 1 2 42544 15484
0 15486 5 1 1 15485
0 15487 7 1 2 15456 15486
0 15488 5 1 1 15487
0 15489 7 1 2 43903 15488
0 15490 5 1 1 15489
0 15491 7 1 2 49127 57124
0 15492 5 1 1 15491
0 15493 7 1 2 65259 15492
0 15494 5 1 1 15493
0 15495 7 1 2 65268 15494
0 15496 5 1 1 15495
0 15497 7 1 2 48428 15496
0 15498 5 1 1 15497
0 15499 7 2 2 51795 59277
0 15500 5 2 1 65269
0 15501 7 2 2 65266 65271
0 15502 5 2 1 65273
0 15503 7 1 2 44067 65275
0 15504 5 1 1 15503
0 15505 7 1 2 53010 59278
0 15506 5 1 1 15505
0 15507 7 1 2 15504 15506
0 15508 5 1 1 15507
0 15509 7 1 2 54215 15508
0 15510 5 1 1 15509
0 15511 7 1 2 15498 15510
0 15512 5 1 1 15511
0 15513 7 1 2 42545 15512
0 15514 5 1 1 15513
0 15515 7 1 2 15490 15514
0 15516 5 1 1 15515
0 15517 7 1 2 43739 15516
0 15518 5 1 1 15517
0 15519 7 1 2 53445 65129
0 15520 5 1 1 15519
0 15521 7 1 2 52062 15520
0 15522 5 1 1 15521
0 15523 7 1 2 52936 58541
0 15524 5 1 1 15523
0 15525 7 1 2 13560 15524
0 15526 7 1 2 15522 15525
0 15527 5 1 1 15526
0 15528 7 1 2 51141 15527
0 15529 5 1 1 15528
0 15530 7 1 2 49978 54044
0 15531 7 1 2 54175 15530
0 15532 5 1 1 15531
0 15533 7 1 2 15529 15532
0 15534 5 1 1 15533
0 15535 7 1 2 62862 15534
0 15536 5 1 1 15535
0 15537 7 4 2 54216 56512
0 15538 7 1 2 49441 65277
0 15539 7 1 2 65276 15538
0 15540 5 1 1 15539
0 15541 7 1 2 15536 15540
0 15542 7 1 2 15518 15541
0 15543 5 1 1 15542
0 15544 7 1 2 60399 15543
0 15545 5 1 1 15544
0 15546 7 1 2 15411 15545
0 15547 5 1 1 15546
0 15548 7 1 2 48619 15547
0 15549 5 1 1 15548
0 15550 7 2 2 45071 51174
0 15551 5 1 1 65281
0 15552 7 1 2 53214 55028
0 15553 5 1 1 15552
0 15554 7 2 2 15551 15553
0 15555 7 1 2 49550 65283
0 15556 5 1 1 15555
0 15557 7 1 2 54252 1590
0 15558 7 1 2 9263 15557
0 15559 7 1 2 59093 15558
0 15560 5 1 1 15559
0 15561 7 1 2 15556 15560
0 15562 5 1 1 15561
0 15563 7 1 2 45251 15562
0 15564 5 1 1 15563
0 15565 7 1 2 55021 60243
0 15566 5 1 1 15565
0 15567 7 1 2 50767 52871
0 15568 5 3 1 15567
0 15569 7 1 2 53404 65285
0 15570 5 6 1 15569
0 15571 7 1 2 53268 65288
0 15572 5 1 1 15571
0 15573 7 1 2 15566 15572
0 15574 7 1 2 15564 15573
0 15575 5 1 1 15574
0 15576 7 1 2 46234 15575
0 15577 5 1 1 15576
0 15578 7 4 2 13924 65229
0 15579 7 1 2 61682 63516
0 15580 5 8 1 15579
0 15581 7 1 2 58566 65298
0 15582 7 1 2 65294 15581
0 15583 5 1 1 15582
0 15584 7 1 2 15577 15583
0 15585 5 1 1 15584
0 15586 7 1 2 44762 15585
0 15587 5 1 1 15586
0 15588 7 1 2 46488 52413
0 15589 5 1 1 15588
0 15590 7 1 2 52350 15589
0 15591 5 1 1 15590
0 15592 7 1 2 47276 15591
0 15593 5 1 1 15592
0 15594 7 1 2 50266 65045
0 15595 5 1 1 15594
0 15596 7 1 2 15593 15595
0 15597 5 1 1 15596
0 15598 7 1 2 46235 15597
0 15599 5 1 1 15598
0 15600 7 2 2 46489 57899
0 15601 7 2 2 49578 65306
0 15602 5 1 1 65308
0 15603 7 1 2 15599 15602
0 15604 5 1 1 15603
0 15605 7 1 2 51297 15604
0 15606 5 1 1 15605
0 15607 7 1 2 15587 15606
0 15608 5 1 1 15607
0 15609 7 1 2 47424 15608
0 15610 5 1 1 15609
0 15611 7 1 2 51059 53115
0 15612 5 1 1 15611
0 15613 7 2 2 46236 49566
0 15614 7 1 2 43740 65310
0 15615 5 1 1 15614
0 15616 7 1 2 15612 15615
0 15617 5 1 1 15616
0 15618 7 1 2 52296 15617
0 15619 5 1 1 15618
0 15620 7 2 2 52365 52615
0 15621 7 1 2 46237 60136
0 15622 7 1 2 65312 15621
0 15623 5 1 1 15622
0 15624 7 1 2 15619 15623
0 15625 5 1 1 15624
0 15626 7 1 2 44763 15625
0 15627 5 1 1 15626
0 15628 7 1 2 46490 52344
0 15629 5 1 1 15628
0 15630 7 1 2 52418 15629
0 15631 5 1 1 15630
0 15632 7 5 2 45072 64913
0 15633 7 1 2 54098 65314
0 15634 7 1 2 15631 15633
0 15635 5 1 1 15634
0 15636 7 1 2 15627 15635
0 15637 5 1 1 15636
0 15638 7 1 2 46028 15637
0 15639 5 1 1 15638
0 15640 7 1 2 47117 65313
0 15641 5 1 1 15640
0 15642 7 1 2 49579 54936
0 15643 5 1 1 15642
0 15644 7 1 2 15641 15643
0 15645 5 1 1 15644
0 15646 7 1 2 46681 15645
0 15647 5 1 1 15646
0 15648 7 1 2 45252 49421
0 15649 7 1 2 50299 15648
0 15650 5 1 1 15649
0 15651 7 1 2 15647 15650
0 15652 5 1 1 15651
0 15653 7 1 2 44764 53853
0 15654 7 1 2 15652 15653
0 15655 5 1 1 15654
0 15656 7 1 2 15639 15655
0 15657 7 1 2 15610 15656
0 15658 5 1 1 15657
0 15659 7 1 2 47973 15658
0 15660 5 1 1 15659
0 15661 7 1 2 55200 62812
0 15662 5 1 1 15661
0 15663 7 1 2 5294 15662
0 15664 5 1 1 15663
0 15665 7 1 2 43300 15664
0 15666 5 1 1 15665
0 15667 7 1 2 52509 57163
0 15668 5 1 1 15667
0 15669 7 1 2 15666 15668
0 15670 5 2 1 15669
0 15671 7 1 2 42792 65319
0 15672 5 1 1 15671
0 15673 7 1 2 53956 60137
0 15674 5 1 1 15673
0 15675 7 1 2 12711 15674
0 15676 5 1 1 15675
0 15677 7 1 2 47544 15676
0 15678 5 1 1 15677
0 15679 7 1 2 49551 53269
0 15680 5 1 1 15679
0 15681 7 1 2 15678 15680
0 15682 7 1 2 15672 15681
0 15683 5 1 1 15682
0 15684 7 1 2 45253 15683
0 15685 5 1 1 15684
0 15686 7 2 2 53270 57374
0 15687 5 1 1 65321
0 15688 7 1 2 15685 15687
0 15689 5 1 1 15688
0 15690 7 1 2 47425 15689
0 15691 5 1 1 15690
0 15692 7 2 2 53162 65224
0 15693 5 2 1 65323
0 15694 7 1 2 46029 65324
0 15695 5 1 1 15694
0 15696 7 3 2 46238 49083
0 15697 5 1 1 65327
0 15698 7 1 2 52419 15697
0 15699 5 1 1 15698
0 15700 7 1 2 53271 15699
0 15701 5 1 1 15700
0 15702 7 1 2 15695 15701
0 15703 7 1 2 15691 15702
0 15704 5 1 1 15703
0 15705 7 1 2 61153 15704
0 15706 5 1 1 15705
0 15707 7 1 2 44643 56600
0 15708 7 1 2 64770 15707
0 15709 5 1 1 15708
0 15710 7 1 2 15706 15709
0 15711 5 1 1 15710
0 15712 7 1 2 54272 15711
0 15713 5 1 1 15712
0 15714 7 1 2 55128 61729
0 15715 5 1 1 15714
0 15716 7 1 2 11765 15715
0 15717 5 1 1 15716
0 15718 7 1 2 42546 15717
0 15719 5 1 1 15718
0 15720 7 1 2 55070 61882
0 15721 5 1 1 15720
0 15722 7 1 2 15719 15721
0 15723 5 1 1 15722
0 15724 7 1 2 53452 15723
0 15725 5 1 1 15724
0 15726 7 1 2 56822 65072
0 15727 5 1 1 15726
0 15728 7 1 2 65193 15727
0 15729 5 2 1 15728
0 15730 7 1 2 42547 65330
0 15731 5 1 1 15730
0 15732 7 1 2 61883 64998
0 15733 5 1 1 15732
0 15734 7 1 2 15731 15733
0 15735 5 4 1 15734
0 15736 7 1 2 49552 60827
0 15737 5 1 1 15736
0 15738 7 6 2 42793 49694
0 15739 5 2 1 65336
0 15740 7 1 2 49538 65342
0 15741 5 4 1 15740
0 15742 7 1 2 63533 65344
0 15743 7 1 2 15737 15742
0 15744 5 1 1 15743
0 15745 7 1 2 65332 15744
0 15746 5 1 1 15745
0 15747 7 1 2 49553 61707
0 15748 7 1 2 64347 15747
0 15749 7 1 2 65087 15748
0 15750 5 1 1 15749
0 15751 7 1 2 15746 15750
0 15752 7 1 2 15725 15751
0 15753 7 1 2 15713 15752
0 15754 7 1 2 15660 15753
0 15755 5 1 1 15754
0 15756 7 1 2 59279 15755
0 15757 5 1 1 15756
0 15758 7 1 2 50275 62779
0 15759 5 1 1 15758
0 15760 7 1 2 65274 15759
0 15761 5 1 1 15760
0 15762 7 1 2 60990 15761
0 15763 5 1 1 15762
0 15764 7 1 2 50075 51826
0 15765 7 1 2 61380 15764
0 15766 5 1 1 15765
0 15767 7 1 2 61663 62637
0 15768 7 1 2 59088 15767
0 15769 5 1 1 15768
0 15770 7 1 2 15766 15769
0 15771 5 1 1 15770
0 15772 7 1 2 44068 15771
0 15773 5 1 1 15772
0 15774 7 1 2 51930 52805
0 15775 7 1 2 61401 15774
0 15776 5 1 1 15775
0 15777 7 1 2 15773 15776
0 15778 7 1 2 15763 15777
0 15779 5 1 1 15778
0 15780 7 1 2 54016 15779
0 15781 5 1 1 15780
0 15782 7 1 2 52860 57874
0 15783 7 1 2 59688 60991
0 15784 7 1 2 15782 15783
0 15785 5 1 1 15784
0 15786 7 1 2 15781 15785
0 15787 5 1 1 15786
0 15788 7 1 2 52616 15787
0 15789 5 1 1 15788
0 15790 7 1 2 63492 65220
0 15791 5 1 1 15790
0 15792 7 1 2 51100 57412
0 15793 5 1 1 15792
0 15794 7 1 2 15791 15793
0 15795 5 1 1 15794
0 15796 7 1 2 54273 15795
0 15797 5 1 1 15796
0 15798 7 2 2 49979 56212
0 15799 5 2 1 65348
0 15800 7 1 2 61503 65350
0 15801 5 1 1 15800
0 15802 7 1 2 65295 15801
0 15803 5 1 1 15802
0 15804 7 1 2 15797 15803
0 15805 5 1 1 15804
0 15806 7 1 2 45448 15805
0 15807 5 1 1 15806
0 15808 7 1 2 54292 63499
0 15809 5 1 1 15808
0 15810 7 1 2 15807 15809
0 15811 5 1 1 15810
0 15812 7 1 2 47426 15811
0 15813 5 1 1 15812
0 15814 7 1 2 42794 50129
0 15815 5 1 1 15814
0 15816 7 1 2 54293 15815
0 15817 5 1 1 15816
0 15818 7 1 2 61497 63502
0 15819 7 1 2 65284 15818
0 15820 5 1 1 15819
0 15821 7 1 2 15817 15820
0 15822 7 1 2 15813 15821
0 15823 5 1 1 15822
0 15824 7 1 2 44765 15823
0 15825 5 1 1 15824
0 15826 7 1 2 47277 60832
0 15827 5 1 1 15826
0 15828 7 1 2 46491 57000
0 15829 7 1 2 58469 15828
0 15830 5 1 1 15829
0 15831 7 1 2 15827 15830
0 15832 5 1 1 15831
0 15833 7 1 2 46239 15832
0 15834 5 1 1 15833
0 15835 7 1 2 62107 15834
0 15836 5 1 1 15835
0 15837 7 1 2 50413 65172
0 15838 7 1 2 15836 15837
0 15839 5 1 1 15838
0 15840 7 1 2 15825 15839
0 15841 5 1 1 15840
0 15842 7 1 2 45254 15841
0 15843 5 1 1 15842
0 15844 7 3 2 48107 52617
0 15845 5 1 1 65352
0 15846 7 1 2 49283 2580
0 15847 7 1 2 4439 15846
0 15848 7 1 2 15845 15847
0 15849 5 1 1 15848
0 15850 7 3 2 44766 54274
0 15851 7 1 2 43741 65355
0 15852 5 1 1 15851
0 15853 7 1 2 15849 15852
0 15854 5 1 1 15853
0 15855 7 1 2 50076 15854
0 15856 5 1 1 15855
0 15857 7 2 2 51002 57816
0 15858 7 6 2 47278 65173
0 15859 7 1 2 50213 65360
0 15860 7 1 2 65358 15859
0 15861 5 1 1 15860
0 15862 7 1 2 15856 15861
0 15863 5 1 1 15862
0 15864 7 1 2 46030 15863
0 15865 5 1 1 15864
0 15866 7 1 2 49284 55046
0 15867 5 1 1 15866
0 15868 7 1 2 55051 15867
0 15869 5 1 1 15868
0 15870 7 1 2 50077 64921
0 15871 7 1 2 15869 15870
0 15872 5 1 1 15871
0 15873 7 1 2 15865 15872
0 15874 5 1 1 15873
0 15875 7 1 2 46240 15874
0 15876 5 1 1 15875
0 15877 7 1 2 53272 58850
0 15878 7 1 2 65356 15877
0 15879 5 1 1 15878
0 15880 7 1 2 15876 15879
0 15881 7 1 2 15843 15880
0 15882 5 1 1 15881
0 15883 7 1 2 47974 15882
0 15884 5 1 1 15883
0 15885 7 1 2 63509 65333
0 15886 5 1 1 15885
0 15887 7 3 2 44767 52750
0 15888 7 2 2 51832 65366
0 15889 7 1 2 61007 65369
0 15890 5 1 1 15889
0 15891 7 1 2 65194 15890
0 15892 5 1 1 15891
0 15893 7 1 2 42548 15892
0 15894 5 1 1 15893
0 15895 7 1 2 62073 65168
0 15896 5 1 1 15895
0 15897 7 1 2 15894 15896
0 15898 5 1 1 15897
0 15899 7 1 2 43080 15898
0 15900 5 1 1 15899
0 15901 7 1 2 56142 65075
0 15902 7 1 2 64835 15901
0 15903 5 1 1 15902
0 15904 7 1 2 15900 15903
0 15905 5 1 1 15904
0 15906 7 1 2 57310 15905
0 15907 5 1 1 15906
0 15908 7 1 2 15886 15907
0 15909 7 1 2 15884 15908
0 15910 5 1 1 15909
0 15911 7 1 2 51931 15910
0 15912 5 1 1 15911
0 15913 7 1 2 15789 15912
0 15914 7 1 2 15757 15913
0 15915 7 1 2 15549 15914
0 15916 5 1 1 15915
0 15917 7 4 2 55845 60322
0 15918 7 1 2 48894 65371
0 15919 7 1 2 15916 15918
0 15920 5 1 1 15919
0 15921 7 1 2 42170 64786
0 15922 5 1 1 15921
0 15923 7 1 2 47890 64962
0 15924 5 1 1 15923
0 15925 7 1 2 7137 15924
0 15926 7 1 2 64784 15925
0 15927 5 1 1 15926
0 15928 7 1 2 15922 15927
0 15929 5 1 1 15928
0 15930 7 1 2 44211 15929
0 15931 5 1 1 15930
0 15932 7 1 2 63138 62771
0 15933 5 2 1 15932
0 15934 7 1 2 53391 65375
0 15935 5 1 1 15934
0 15936 7 1 2 53329 63133
0 15937 5 1 1 15936
0 15938 7 1 2 10035 15937
0 15939 5 1 1 15938
0 15940 7 1 2 49755 15939
0 15941 5 1 1 15940
0 15942 7 1 2 15935 15941
0 15943 5 1 1 15942
0 15944 7 1 2 47545 15943
0 15945 5 1 1 15944
0 15946 7 2 2 52073 64248
0 15947 5 1 1 65377
0 15948 7 1 2 47279 65378
0 15949 5 1 1 15948
0 15950 7 1 2 15945 15949
0 15951 5 1 1 15950
0 15952 7 1 2 43301 15951
0 15953 5 1 1 15952
0 15954 7 1 2 62580 64233
0 15955 5 1 1 15954
0 15956 7 1 2 47546 61982
0 15957 7 1 2 64763 15956
0 15958 5 1 1 15957
0 15959 7 1 2 15955 15958
0 15960 7 1 2 15953 15959
0 15961 5 1 1 15960
0 15962 7 1 2 61154 15961
0 15963 5 1 1 15962
0 15964 7 1 2 15931 15963
0 15965 5 1 1 15964
0 15966 7 1 2 48429 15965
0 15967 5 1 1 15966
0 15968 7 1 2 51932 62039
0 15969 5 1 1 15968
0 15970 7 1 2 45255 62897
0 15971 5 1 1 15970
0 15972 7 1 2 15969 15971
0 15973 5 1 1 15972
0 15974 7 1 2 49047 15973
0 15975 5 1 1 15974
0 15976 7 1 2 59280 64805
0 15977 5 1 1 15976
0 15978 7 1 2 45718 64807
0 15979 5 1 1 15978
0 15980 7 1 2 15977 15979
0 15981 5 1 1 15980
0 15982 7 1 2 49695 15981
0 15983 5 1 1 15982
0 15984 7 1 2 64812 65247
0 15985 5 1 1 15984
0 15986 7 1 2 15983 15985
0 15987 7 1 2 15975 15986
0 15988 5 1 1 15987
0 15989 7 1 2 47280 15988
0 15990 5 1 1 15989
0 15991 7 2 2 55708 62655
0 15992 5 1 1 65379
0 15993 7 1 2 12188 15992
0 15994 5 1 1 15993
0 15995 7 1 2 49756 15994
0 15996 5 1 1 15995
0 15997 7 1 2 53033 65376
0 15998 5 1 1 15997
0 15999 7 1 2 15996 15998
0 16000 5 1 1 15999
0 16001 7 1 2 47547 16000
0 16002 5 1 1 16001
0 16003 7 1 2 15947 16002
0 16004 5 1 1 16003
0 16005 7 1 2 43904 16004
0 16006 5 1 1 16005
0 16007 7 1 2 51504 57151
0 16008 7 1 2 62803 16007
0 16009 5 1 1 16008
0 16010 7 1 2 16006 16009
0 16011 7 1 2 15990 16010
0 16012 5 1 1 16011
0 16013 7 1 2 43302 16012
0 16014 5 1 1 16013
0 16015 7 1 2 59281 64824
0 16016 5 1 1 16015
0 16017 7 1 2 64826 16016
0 16018 5 1 1 16017
0 16019 7 1 2 64234 16018
0 16020 5 1 1 16019
0 16021 7 1 2 16014 16020
0 16022 5 1 1 16021
0 16023 7 1 2 45073 16022
0 16024 5 1 1 16023
0 16025 7 1 2 62198 64779
0 16026 7 1 2 64814 16025
0 16027 5 1 1 16026
0 16028 7 1 2 16024 16027
0 16029 5 1 1 16028
0 16030 7 1 2 61155 16029
0 16031 5 1 1 16030
0 16032 7 1 2 15967 16031
0 16033 5 1 1 16032
0 16034 7 1 2 53273 16033
0 16035 5 1 1 16034
0 16036 7 1 2 51933 64870
0 16037 5 1 1 16036
0 16038 7 1 2 59282 64933
0 16039 5 1 1 16038
0 16040 7 1 2 45719 64954
0 16041 5 1 1 16040
0 16042 7 1 2 54937 59689
0 16043 7 1 2 64990 16042
0 16044 5 1 1 16043
0 16045 7 1 2 61851 64967
0 16046 5 1 1 16045
0 16047 7 1 2 61203 64983
0 16048 5 1 1 16047
0 16049 7 1 2 16046 16048
0 16050 5 1 1 16049
0 16051 7 1 2 43905 16050
0 16052 5 1 1 16051
0 16053 7 1 2 16044 16052
0 16054 7 1 2 16041 16053
0 16055 5 1 1 16054
0 16056 7 1 2 42549 16055
0 16057 5 1 1 16056
0 16058 7 1 2 60791 65003
0 16059 5 1 1 16058
0 16060 7 1 2 45720 65019
0 16061 5 1 1 16060
0 16062 7 1 2 61852 65035
0 16063 5 1 1 16062
0 16064 7 1 2 16061 16063
0 16065 5 1 1 16064
0 16066 7 1 2 42795 16065
0 16067 5 1 1 16066
0 16068 7 1 2 16059 16067
0 16069 7 1 2 16057 16068
0 16070 5 1 1 16069
0 16071 7 1 2 49218 16070
0 16072 5 1 1 16071
0 16073 7 1 2 16039 16072
0 16074 7 1 2 16037 16073
0 16075 7 1 2 16035 16074
0 16076 5 1 1 16075
0 16077 7 1 2 47759 63040
0 16078 7 1 2 16076 16077
0 16079 5 1 1 16078
0 16080 7 1 2 44321 16079
0 16081 7 1 2 15920 16080
0 16082 7 1 2 15235 16081
0 16083 5 1 1 16082
0 16084 7 3 2 45074 50555
0 16085 7 2 2 58970 65381
0 16086 7 1 2 61363 65384
0 16087 5 1 1 16086
0 16088 7 1 2 53773 62652
0 16089 7 1 2 59801 16088
0 16090 5 1 1 16089
0 16091 7 1 2 16087 16090
0 16092 5 1 1 16091
0 16093 7 1 2 50768 16092
0 16094 5 1 1 16093
0 16095 7 1 2 43906 50259
0 16096 5 1 1 16095
0 16097 7 1 2 56317 16096
0 16098 5 3 1 16097
0 16099 7 1 2 42796 65386
0 16100 5 1 1 16099
0 16101 7 2 2 49449 55161
0 16102 5 1 1 65389
0 16103 7 1 2 16100 16102
0 16104 5 1 1 16103
0 16105 7 1 2 59033 16104
0 16106 5 1 1 16105
0 16107 7 1 2 48807 57527
0 16108 7 1 2 65163 16107
0 16109 5 1 1 16108
0 16110 7 1 2 16106 16109
0 16111 5 1 1 16110
0 16112 7 1 2 60400 16111
0 16113 5 1 1 16112
0 16114 7 1 2 16094 16113
0 16115 5 1 1 16114
0 16116 7 1 2 43742 16115
0 16117 5 1 1 16116
0 16118 7 1 2 55522 58589
0 16119 5 1 1 16118
0 16120 7 1 2 47281 64549
0 16121 5 1 1 16120
0 16122 7 1 2 54326 61245
0 16123 5 1 1 16122
0 16124 7 1 2 16121 16123
0 16125 5 1 1 16124
0 16126 7 1 2 46241 16125
0 16127 5 1 1 16126
0 16128 7 1 2 16119 16127
0 16129 5 1 1 16128
0 16130 7 1 2 50260 16129
0 16131 5 1 1 16130
0 16132 7 2 2 49166 56506
0 16133 7 1 2 52980 57014
0 16134 7 1 2 65391 16133
0 16135 5 1 1 16134
0 16136 7 1 2 60292 64550
0 16137 5 1 1 16136
0 16138 7 1 2 50306 64739
0 16139 5 1 1 16138
0 16140 7 1 2 16137 16139
0 16141 5 2 1 16140
0 16142 7 1 2 65382 65393
0 16143 5 1 1 16142
0 16144 7 1 2 16135 16143
0 16145 7 1 2 16131 16144
0 16146 5 1 1 16145
0 16147 7 1 2 61520 16146
0 16148 5 1 1 16147
0 16149 7 1 2 16117 16148
0 16150 5 1 1 16149
0 16151 7 1 2 42550 16150
0 16152 5 1 1 16151
0 16153 7 1 2 55081 64551
0 16154 5 1 1 16153
0 16155 7 1 2 60059 64283
0 16156 5 1 1 16155
0 16157 7 1 2 16154 16156
0 16158 5 1 1 16157
0 16159 7 1 2 50261 16158
0 16160 5 1 1 16159
0 16161 7 1 2 47118 56507
0 16162 5 1 1 16161
0 16163 7 1 2 1574 16162
0 16164 5 3 1 16163
0 16165 7 1 2 65394 65395
0 16166 5 1 1 16165
0 16167 7 1 2 54938 58035
0 16168 7 1 2 65392 16167
0 16169 5 1 1 16168
0 16170 7 1 2 16166 16169
0 16171 7 1 2 16160 16170
0 16172 5 1 1 16171
0 16173 7 1 2 44768 16172
0 16174 5 1 1 16173
0 16175 7 3 2 61525 65361
0 16176 5 2 1 65398
0 16177 7 1 2 47119 52415
0 16178 7 1 2 65399 16177
0 16179 5 1 1 16178
0 16180 7 1 2 16174 16179
0 16181 5 1 1 16180
0 16182 7 1 2 61874 16181
0 16183 5 1 1 16182
0 16184 7 2 2 16152 16183
0 16185 5 1 1 65403
0 16186 7 1 2 64476 65132
0 16187 5 1 1 16186
0 16188 7 1 2 49858 53740
0 16189 7 1 2 62012 16188
0 16190 5 1 1 16189
0 16191 7 1 2 16187 16190
0 16192 5 1 1 16191
0 16193 7 1 2 42551 16192
0 16194 5 1 1 16193
0 16195 7 1 2 47120 65387
0 16196 5 1 1 16195
0 16197 7 1 2 65149 16196
0 16198 5 1 1 16197
0 16199 7 2 2 59592 61156
0 16200 7 1 2 16198 65405
0 16201 5 1 1 16200
0 16202 7 1 2 16194 16201
0 16203 5 1 1 16202
0 16204 7 1 2 42797 16203
0 16205 5 1 1 16204
0 16206 7 4 2 47282 50262
0 16207 5 1 1 65407
0 16208 7 1 2 1470 16207
0 16209 5 1 1 16208
0 16210 7 1 2 53274 16209
0 16211 5 1 1 16210
0 16212 7 1 2 47121 56639
0 16213 5 1 1 16212
0 16214 7 1 2 16211 16213
0 16215 5 1 1 16214
0 16216 7 1 2 56213 61157
0 16217 7 1 2 16215 16216
0 16218 5 1 1 16217
0 16219 7 1 2 16205 16218
0 16220 5 1 1 16219
0 16221 7 1 2 55578 16220
0 16222 5 1 1 16221
0 16223 7 1 2 65404 16222
0 16224 5 1 1 16223
0 16225 7 1 2 58720 16224
0 16226 5 1 1 16225
0 16227 7 1 2 42798 65331
0 16228 5 1 1 16227
0 16229 7 1 2 62295 65357
0 16230 5 1 1 16229
0 16231 7 1 2 16228 16230
0 16232 5 1 1 16231
0 16233 7 1 2 42552 16232
0 16234 5 1 1 16233
0 16235 7 1 2 61884 65154
0 16236 5 1 1 16235
0 16237 7 1 2 16234 16236
0 16238 5 2 1 16237
0 16239 7 1 2 52897 65411
0 16240 5 1 1 16239
0 16241 7 1 2 53275 65164
0 16242 5 1 1 16241
0 16243 7 1 2 55117 16242
0 16244 5 1 1 16243
0 16245 7 1 2 44769 16244
0 16246 5 1 1 16245
0 16247 7 1 2 61715 65362
0 16248 5 1 1 16247
0 16249 7 1 2 16246 16248
0 16250 5 1 1 16249
0 16251 7 1 2 50556 62833
0 16252 7 1 2 16250 16251
0 16253 5 1 1 16252
0 16254 7 1 2 16240 16253
0 16255 5 2 1 16254
0 16256 7 1 2 51226 65413
0 16257 5 1 1 16256
0 16258 7 2 2 50637 61989
0 16259 5 3 1 65415
0 16260 7 1 2 65334 65416
0 16261 5 1 1 16260
0 16262 7 1 2 61381 64422
0 16263 5 1 1 16262
0 16264 7 1 2 53276 53719
0 16265 7 1 2 62840 16264
0 16266 5 1 1 16265
0 16267 7 1 2 16263 16266
0 16268 5 1 1 16267
0 16269 7 1 2 54275 16268
0 16270 5 1 1 16269
0 16271 7 1 2 16261 16270
0 16272 5 1 1 16271
0 16273 7 1 2 51754 16272
0 16274 5 1 1 16273
0 16275 7 1 2 61382 65165
0 16276 5 1 1 16275
0 16277 7 3 2 45075 53277
0 16278 7 1 2 62016 65420
0 16279 5 1 1 16278
0 16280 7 1 2 16276 16279
0 16281 5 1 1 16280
0 16282 7 1 2 50632 51755
0 16283 5 1 1 16282
0 16284 7 1 2 57559 16283
0 16285 5 1 1 16284
0 16286 7 1 2 16281 16285
0 16287 5 1 1 16286
0 16288 7 1 2 16274 16287
0 16289 7 1 2 16257 16288
0 16290 5 1 1 16289
0 16291 7 1 2 61049 16290
0 16292 5 1 1 16291
0 16293 7 1 2 16226 16292
0 16294 5 1 1 16293
0 16295 7 1 2 62686 16294
0 16296 5 1 1 16295
0 16297 7 6 2 45804 47760
0 16298 7 2 2 63066 65423
0 16299 7 1 2 16185 65429
0 16300 5 1 1 16299
0 16301 7 1 2 56187 63349
0 16302 5 1 1 16301
0 16303 7 4 2 43081 47761
0 16304 7 1 2 47427 65431
0 16305 7 1 2 62987 16304
0 16306 5 1 1 16305
0 16307 7 1 2 16302 16306
0 16308 5 1 1 16307
0 16309 7 1 2 65008 16308
0 16310 5 1 1 16309
0 16311 7 1 2 55124 64394
0 16312 7 1 2 64575 65013
0 16313 7 1 2 16311 16312
0 16314 5 1 1 16313
0 16315 7 1 2 16310 16314
0 16316 5 1 1 16315
0 16317 7 1 2 61158 16316
0 16318 5 1 1 16317
0 16319 7 2 2 60992 65372
0 16320 7 1 2 48808 65435
0 16321 7 1 2 52689 16320
0 16322 5 1 1 16321
0 16323 7 1 2 16318 16322
0 16324 5 1 1 16323
0 16325 7 1 2 42799 16324
0 16326 5 1 1 16325
0 16327 7 2 2 45805 64538
0 16328 7 1 2 57592 61462
0 16329 7 1 2 64315 16328
0 16330 7 1 2 65437 16329
0 16331 7 1 2 54294 16330
0 16332 5 1 1 16331
0 16333 7 1 2 16326 16332
0 16334 5 1 1 16333
0 16335 7 1 2 45256 16334
0 16336 5 1 1 16335
0 16337 7 1 2 45076 61720
0 16338 7 1 2 62077 16337
0 16339 5 1 1 16338
0 16340 7 1 2 52872 63935
0 16341 7 1 2 62013 16340
0 16342 5 1 1 16341
0 16343 7 1 2 16339 16342
0 16344 5 1 1 16343
0 16345 7 1 2 42553 16344
0 16346 5 1 1 16345
0 16347 7 1 2 65170 65406
0 16348 5 1 1 16347
0 16349 7 1 2 16346 16348
0 16350 5 1 1 16349
0 16351 7 1 2 62988 64194
0 16352 7 1 2 16350 16351
0 16353 5 1 1 16352
0 16354 7 1 2 16336 16353
0 16355 5 1 1 16354
0 16356 7 1 2 55579 16355
0 16357 5 1 1 16356
0 16358 7 1 2 62646 64977
0 16359 5 1 1 16358
0 16360 7 1 2 50414 65363
0 16361 5 1 1 16360
0 16362 7 1 2 16359 16361
0 16363 5 1 1 16362
0 16364 7 1 2 62976 16363
0 16365 5 1 1 16364
0 16366 7 2 2 50078 60829
0 16367 7 1 2 43907 65439
0 16368 5 1 1 16367
0 16369 7 1 2 58801 16368
0 16370 5 1 1 16369
0 16371 7 1 2 45257 16370
0 16372 5 1 1 16371
0 16373 7 1 2 50330 64439
0 16374 5 1 1 16373
0 16375 7 1 2 16372 16374
0 16376 5 1 1 16375
0 16377 7 1 2 46492 16376
0 16378 5 1 1 16377
0 16379 7 1 2 52314 57170
0 16380 5 1 1 16379
0 16381 7 1 2 16378 16380
0 16382 5 1 1 16381
0 16383 7 1 2 50696 53278
0 16384 7 1 2 16382 16383
0 16385 5 1 1 16384
0 16386 7 1 2 16365 16385
0 16387 5 1 1 16386
0 16388 7 1 2 61414 16387
0 16389 5 1 1 16388
0 16390 7 1 2 61342 61730
0 16391 5 1 1 16390
0 16392 7 1 2 61426 16391
0 16393 5 2 1 16392
0 16394 7 2 2 49980 50944
0 16395 5 3 1 65443
0 16396 7 1 2 62947 65445
0 16397 5 4 1 16396
0 16398 7 1 2 65441 65448
0 16399 5 1 1 16398
0 16400 7 2 2 42800 58576
0 16401 5 2 1 65452
0 16402 7 1 2 52885 55008
0 16403 5 1 1 16402
0 16404 7 3 2 65454 16403
0 16405 7 3 2 50079 65456
0 16406 5 3 1 65459
0 16407 7 1 2 57669 58557
0 16408 5 1 1 16407
0 16409 7 1 2 46242 16408
0 16410 5 1 1 16409
0 16411 7 1 2 65462 16410
0 16412 5 1 1 16411
0 16413 7 1 2 62978 16412
0 16414 5 1 1 16413
0 16415 7 1 2 16399 16414
0 16416 5 1 1 16415
0 16417 7 1 2 54276 16416
0 16418 5 1 1 16417
0 16419 7 1 2 42801 64592
0 16420 5 1 1 16419
0 16421 7 2 2 42802 50080
0 16422 5 6 1 65465
0 16423 7 1 2 52898 65466
0 16424 5 2 1 16423
0 16425 7 1 2 4117 65473
0 16426 7 1 2 16420 16425
0 16427 5 1 1 16426
0 16428 7 1 2 65335 16427
0 16429 5 1 1 16428
0 16430 7 1 2 16418 16429
0 16431 7 1 2 16389 16430
0 16432 5 1 1 16431
0 16433 7 1 2 65373 16432
0 16434 5 1 1 16433
0 16435 7 1 2 16357 16434
0 16436 7 1 2 16300 16435
0 16437 5 1 1 16436
0 16438 7 1 2 59283 16437
0 16439 5 1 1 16438
0 16440 7 1 2 62962 64726
0 16441 5 1 1 16440
0 16442 7 2 2 49696 54845
0 16443 5 2 1 65475
0 16444 7 1 2 46031 65476
0 16445 5 1 1 16444
0 16446 7 1 2 16441 16445
0 16447 5 1 1 16446
0 16448 7 1 2 54277 16447
0 16449 5 1 1 16448
0 16450 7 1 2 51524 54894
0 16451 5 1 1 16450
0 16452 7 1 2 3492 16451
0 16453 5 1 1 16452
0 16454 7 1 2 65009 16453
0 16455 5 1 1 16454
0 16456 7 1 2 16449 16455
0 16457 5 1 1 16456
0 16458 7 1 2 43082 16457
0 16459 5 1 1 16458
0 16460 7 1 2 53763 62170
0 16461 5 1 1 16460
0 16462 7 1 2 54988 8963
0 16463 7 1 2 65421 16462
0 16464 5 1 1 16463
0 16465 7 1 2 16461 16464
0 16466 5 1 1 16465
0 16467 7 1 2 47283 16466
0 16468 5 1 1 16467
0 16469 7 1 2 53076 2299
0 16470 5 1 1 16469
0 16471 7 1 2 53375 65206
0 16472 7 1 2 16470 16471
0 16473 5 1 1 16472
0 16474 7 1 2 16468 16473
0 16475 5 1 1 16474
0 16476 7 1 2 51756 16475
0 16477 5 1 1 16476
0 16478 7 1 2 16459 16477
0 16479 5 1 1 16478
0 16480 7 4 2 44770 65374
0 16481 7 1 2 16479 65479
0 16482 5 1 1 16481
0 16483 7 2 2 54200 65480
0 16484 7 1 2 51757 65483
0 16485 5 1 1 16484
0 16486 7 6 2 44442 50081
0 16487 7 2 2 63350 65485
0 16488 5 1 1 65491
0 16489 7 1 2 51715 65492
0 16490 5 1 1 16489
0 16491 7 5 2 47762 63067
0 16492 7 4 2 45806 47548
0 16493 7 1 2 60743 65498
0 16494 7 1 2 65493 16493
0 16495 5 1 1 16494
0 16496 7 1 2 16490 16495
0 16497 5 1 1 16496
0 16498 7 1 2 49567 51308
0 16499 7 1 2 16497 16498
0 16500 5 1 1 16499
0 16501 7 1 2 16485 16500
0 16502 5 1 1 16501
0 16503 7 1 2 47428 16502
0 16504 5 1 1 16503
0 16505 7 1 2 64272 65484
0 16506 5 1 1 16505
0 16507 7 1 2 16504 16506
0 16508 5 1 1 16507
0 16509 7 1 2 47284 16508
0 16510 5 1 1 16509
0 16511 7 1 2 57722 65422
0 16512 5 1 1 16511
0 16513 7 1 2 167 53770
0 16514 7 1 2 62963 16513
0 16515 5 1 1 16514
0 16516 7 1 2 16512 16515
0 16517 5 1 1 16516
0 16518 7 1 2 43908 65481
0 16519 7 1 2 16517 16518
0 16520 5 1 1 16519
0 16521 7 1 2 46243 16520
0 16522 7 1 2 16510 16521
0 16523 5 1 1 16522
0 16524 7 1 2 1636 9112
0 16525 5 1 1 16524
0 16526 7 2 2 48620 52618
0 16527 5 2 1 65502
0 16528 7 2 2 54681 65504
0 16529 5 2 1 65506
0 16530 7 1 2 16525 65507
0 16531 5 1 1 16530
0 16532 7 1 2 54879 64597
0 16533 5 1 1 16532
0 16534 7 1 2 16531 16533
0 16535 5 1 1 16534
0 16536 7 1 2 51227 16535
0 16537 5 1 1 16536
0 16538 7 1 2 51758 65011
0 16539 5 1 1 16538
0 16540 7 1 2 16537 16539
0 16541 5 1 1 16540
0 16542 7 1 2 65482 16541
0 16543 5 1 1 16542
0 16544 7 1 2 42803 16543
0 16545 5 1 1 16544
0 16546 7 1 2 46493 16545
0 16547 7 1 2 16523 16546
0 16548 5 1 1 16547
0 16549 7 1 2 16482 16548
0 16550 5 1 1 16549
0 16551 7 1 2 47975 16550
0 16552 5 1 1 16551
0 16553 7 4 2 45807 54964
0 16554 7 1 2 65494 65510
0 16555 7 1 2 65322 16554
0 16556 5 1 1 16555
0 16557 7 1 2 54387 56064
0 16558 7 1 2 60323 16557
0 16559 7 1 2 60842 16558
0 16560 5 1 1 16559
0 16561 7 1 2 16556 16560
0 16562 5 1 1 16561
0 16563 7 1 2 61159 16562
0 16564 5 1 1 16563
0 16565 7 1 2 54534 64458
0 16566 7 1 2 64576 16565
0 16567 7 1 2 63433 16566
0 16568 5 1 1 16567
0 16569 7 1 2 16564 16568
0 16570 5 1 1 16569
0 16571 7 1 2 65388 16570
0 16572 5 1 1 16571
0 16573 7 1 2 48430 57863
0 16574 5 1 1 16573
0 16575 7 1 2 43909 50323
0 16576 7 1 2 16574 16575
0 16577 5 1 1 16576
0 16578 7 1 2 56318 16577
0 16579 5 1 1 16578
0 16580 7 1 2 43083 16579
0 16581 5 1 1 16580
0 16582 7 1 2 51525 56333
0 16583 5 1 1 16582
0 16584 7 1 2 16581 16583
0 16585 5 1 1 16584
0 16586 7 1 2 42804 16585
0 16587 5 1 1 16586
0 16588 7 1 2 43084 65390
0 16589 5 1 1 16588
0 16590 7 1 2 50633 65166
0 16591 5 1 1 16590
0 16592 7 4 2 42805 53089
0 16593 7 1 2 50520 65514
0 16594 5 1 1 16593
0 16595 7 1 2 16591 16594
0 16596 5 1 1 16595
0 16597 7 1 2 51759 16596
0 16598 5 1 1 16597
0 16599 7 1 2 16589 16598
0 16600 7 1 2 16587 16599
0 16601 5 1 1 16600
0 16602 7 1 2 65436 16601
0 16603 5 1 1 16602
0 16604 7 1 2 16572 16603
0 16605 7 1 2 16552 16604
0 16606 5 1 1 16605
0 16607 7 1 2 51934 16606
0 16608 5 1 1 16607
0 16609 7 3 2 46244 44443
0 16610 7 1 2 42171 62687
0 16611 5 1 1 16610
0 16612 7 3 2 45721 43579
0 16613 5 1 1 65521
0 16614 7 3 2 63341 65522
0 16615 5 1 1 65524
0 16616 7 1 2 16611 16615
0 16617 5 6 1 16616
0 16618 7 1 2 64245 65527
0 16619 5 1 1 16618
0 16620 7 2 2 44563 62707
0 16621 7 12 2 42172 42273
0 16622 7 1 2 49981 65535
0 16623 7 1 2 65533 16622
0 16624 5 1 1 16623
0 16625 7 1 2 16619 16624
0 16626 5 1 1 16625
0 16627 7 1 2 65518 16626
0 16628 5 1 1 16627
0 16629 7 2 2 47891 63794
0 16630 7 3 2 65495 65547
0 16631 7 1 2 63936 65549
0 16632 5 1 1 16631
0 16633 7 1 2 42173 63248
0 16634 7 1 2 63780 16633
0 16635 5 1 1 16634
0 16636 7 1 2 16632 16635
0 16637 5 1 1 16636
0 16638 7 1 2 57375 16637
0 16639 5 1 1 16638
0 16640 7 1 2 16628 16639
0 16641 5 1 1 16640
0 16642 7 1 2 50719 62262
0 16643 5 1 1 16642
0 16644 7 1 2 53097 61396
0 16645 5 1 1 16644
0 16646 7 1 2 16643 16645
0 16647 5 2 1 16646
0 16648 7 1 2 43910 65552
0 16649 5 1 1 16648
0 16650 7 1 2 61397 65408
0 16651 5 1 1 16650
0 16652 7 1 2 16649 16651
0 16653 5 1 1 16652
0 16654 7 1 2 42554 16653
0 16655 5 1 1 16654
0 16656 7 1 2 43911 65396
0 16657 5 1 1 16656
0 16658 7 1 2 43743 65409
0 16659 5 1 1 16658
0 16660 7 1 2 16657 16659
0 16661 5 1 1 16660
0 16662 7 1 2 61885 16661
0 16663 5 1 1 16662
0 16664 7 1 2 16655 16663
0 16665 5 1 1 16664
0 16666 7 1 2 16641 16665
0 16667 5 1 1 16666
0 16668 7 1 2 16608 16667
0 16669 7 1 2 16439 16668
0 16670 7 1 2 16296 16669
0 16671 5 1 1 16670
0 16672 7 1 2 58185 16671
0 16673 5 1 1 16672
0 16674 7 2 2 62989 64249
0 16675 7 1 2 52085 60782
0 16676 5 1 1 16675
0 16677 7 2 2 57560 16676
0 16678 5 3 1 65556
0 16679 7 1 2 46032 65557
0 16680 5 1 1 16679
0 16681 7 1 2 49285 52193
0 16682 5 1 1 16681
0 16683 7 1 2 42555 16682
0 16684 5 2 1 16683
0 16685 7 1 2 64999 65561
0 16686 7 1 2 16680 16685
0 16687 5 1 1 16686
0 16688 7 1 2 54669 65558
0 16689 5 1 1 16688
0 16690 7 3 2 54327 58397
0 16691 7 2 2 49378 65563
0 16692 5 1 1 65566
0 16693 7 1 2 62599 65567
0 16694 5 1 1 16693
0 16695 7 1 2 16689 16694
0 16696 7 1 2 16687 16695
0 16697 5 1 1 16696
0 16698 7 1 2 44771 16697
0 16699 5 1 1 16698
0 16700 7 1 2 49927 62342
0 16701 5 1 1 16700
0 16702 7 1 2 16699 16701
0 16703 5 1 1 16702
0 16704 7 1 2 65554 16703
0 16705 5 1 1 16704
0 16706 7 2 2 45722 62688
0 16707 5 1 1 65568
0 16708 7 1 2 11217 16707
0 16709 5 6 1 16708
0 16710 7 4 2 44564 65570
0 16711 7 1 2 53199 57675
0 16712 5 1 1 16711
0 16713 7 1 2 47122 64209
0 16714 5 1 1 16713
0 16715 7 1 2 56105 64335
0 16716 5 1 1 16715
0 16717 7 1 2 16714 16716
0 16718 5 1 1 16717
0 16719 7 1 2 43912 16718
0 16720 5 1 1 16719
0 16721 7 1 2 43744 64909
0 16722 7 1 2 57109 16721
0 16723 5 1 1 16722
0 16724 7 1 2 16720 16723
0 16725 5 1 1 16724
0 16726 7 1 2 46033 16725
0 16727 5 1 1 16726
0 16728 7 1 2 16712 16727
0 16729 5 1 1 16728
0 16730 7 1 2 53070 16729
0 16731 5 1 1 16730
0 16732 7 1 2 54572 64582
0 16733 5 1 1 16732
0 16734 7 1 2 52693 53215
0 16735 5 1 1 16734
0 16736 7 3 2 42806 57074
0 16737 7 1 2 16735 65580
0 16738 5 1 1 16737
0 16739 7 7 2 48621 50945
0 16740 7 1 2 57376 65583
0 16741 7 1 2 54197 16740
0 16742 5 1 1 16741
0 16743 7 1 2 16738 16742
0 16744 5 1 1 16743
0 16745 7 1 2 65006 16744
0 16746 5 1 1 16745
0 16747 7 1 2 16733 16746
0 16748 7 1 2 16731 16747
0 16749 5 1 1 16748
0 16750 7 1 2 44772 16749
0 16751 5 1 1 16750
0 16752 7 1 2 45449 54573
0 16753 7 1 2 51309 16752
0 16754 7 1 2 57589 16753
0 16755 5 1 1 16754
0 16756 7 1 2 16751 16755
0 16757 5 1 1 16756
0 16758 7 1 2 65576 16757
0 16759 5 1 1 16758
0 16760 7 1 2 16705 16759
0 16761 5 1 1 16760
0 16762 7 1 2 47976 16761
0 16763 5 1 1 16762
0 16764 7 1 2 52675 65581
0 16765 5 1 1 16764
0 16766 7 1 2 46245 64210
0 16767 5 1 1 16766
0 16768 7 1 2 52315 57549
0 16769 5 2 1 16768
0 16770 7 1 2 16767 65590
0 16771 5 1 1 16770
0 16772 7 1 2 48431 16771
0 16773 5 1 1 16772
0 16774 7 1 2 16765 16773
0 16775 5 1 1 16774
0 16776 7 1 2 43913 16775
0 16777 5 1 1 16776
0 16778 7 1 2 54629 65582
0 16779 5 1 1 16778
0 16780 7 1 2 16777 16779
0 16781 5 1 1 16780
0 16782 7 1 2 65577 16781
0 16783 5 1 1 16782
0 16784 7 1 2 53116 65555
0 16785 7 1 2 65559 16784
0 16786 5 1 1 16785
0 16787 7 1 2 16783 16786
0 16788 5 1 1 16787
0 16789 7 1 2 60993 16788
0 16790 5 1 1 16789
0 16791 7 1 2 56750 65578
0 16792 5 1 1 16791
0 16793 7 1 2 62990 62933
0 16794 5 1 1 16793
0 16795 7 1 2 16792 16794
0 16796 5 1 1 16795
0 16797 7 1 2 50946 16796
0 16798 5 1 1 16797
0 16799 7 1 2 56581 60306
0 16800 5 1 1 16799
0 16801 7 1 2 62667 64712
0 16802 5 2 1 16801
0 16803 7 1 2 16800 65592
0 16804 5 1 1 16803
0 16805 7 1 2 45723 16804
0 16806 5 1 1 16805
0 16807 7 1 2 63068 64055
0 16808 5 2 1 16807
0 16809 7 1 2 16806 65594
0 16810 5 1 1 16809
0 16811 7 1 2 52919 16810
0 16812 5 1 1 16811
0 16813 7 2 2 44069 51660
0 16814 5 1 1 65596
0 16815 7 1 2 51816 60307
0 16816 7 1 2 65597 16815
0 16817 5 1 1 16816
0 16818 7 1 2 16812 16817
0 16819 5 1 1 16818
0 16820 7 1 2 51760 16819
0 16821 5 1 1 16820
0 16822 7 1 2 16798 16821
0 16823 5 1 1 16822
0 16824 7 1 2 16823 65442
0 16825 5 1 1 16824
0 16826 7 1 2 55709 57572
0 16827 7 1 2 65571 16826
0 16828 5 1 1 16827
0 16829 7 2 2 55732 56118
0 16830 5 1 1 65598
0 16831 7 1 2 64014 63795
0 16832 7 1 2 52194 16831
0 16833 7 1 2 65599 16832
0 16834 5 1 1 16833
0 16835 7 1 2 16828 16834
0 16836 5 1 1 16835
0 16837 7 1 2 62979 16836
0 16838 5 1 1 16837
0 16839 7 1 2 16825 16838
0 16840 5 1 1 16839
0 16841 7 1 2 54278 16840
0 16842 5 1 1 16841
0 16843 7 2 2 51475 51761
0 16844 5 2 1 65600
0 16845 7 1 2 58818 65602
0 16846 5 1 1 16845
0 16847 7 1 2 51661 16846
0 16848 5 1 1 16847
0 16849 7 3 2 49982 51586
0 16850 5 1 1 65604
0 16851 7 1 2 51080 65605
0 16852 5 2 1 16851
0 16853 7 1 2 16848 65607
0 16854 5 1 1 16853
0 16855 7 1 2 60308 16854
0 16856 5 1 1 16855
0 16857 7 5 2 44565 51081
0 16858 7 3 2 44212 65609
0 16859 7 9 2 42274 46912
0 16860 7 2 2 43303 65617
0 16861 7 1 2 43580 65626
0 16862 7 1 2 65614 16861
0 16863 5 1 1 16862
0 16864 7 1 2 16856 16863
0 16865 5 1 1 16864
0 16866 7 1 2 45724 16865
0 16867 5 1 1 16866
0 16868 7 1 2 61853 62991
0 16869 7 1 2 65615 16868
0 16870 5 1 1 16869
0 16871 7 1 2 16867 16870
0 16872 5 1 1 16871
0 16873 7 1 2 65412 16872
0 16874 5 1 1 16873
0 16875 7 1 2 56969 60309
0 16876 5 1 1 16875
0 16877 7 1 2 65593 16876
0 16878 5 1 1 16877
0 16879 7 1 2 45725 16878
0 16880 5 1 1 16879
0 16881 7 1 2 65595 16880
0 16882 5 1 1 16881
0 16883 7 1 2 50082 16882
0 16884 7 1 2 65414 16883
0 16885 5 1 1 16884
0 16886 7 1 2 16874 16885
0 16887 7 1 2 16842 16886
0 16888 7 1 2 16790 16887
0 16889 7 1 2 16763 16888
0 16890 5 1 1 16889
0 16891 7 1 2 58156 16890
0 16892 5 1 1 16891
0 16893 7 3 2 47285 53279
0 16894 7 2 2 55779 59962
0 16895 7 1 2 43529 65631
0 16896 5 1 1 16895
0 16897 7 2 2 51696 56871
0 16898 7 1 2 47763 65633
0 16899 5 1 1 16898
0 16900 7 1 2 16896 16899
0 16901 5 1 1 16900
0 16902 7 1 2 60310 16901
0 16903 5 1 1 16902
0 16904 7 1 2 62672 65632
0 16905 5 1 1 16904
0 16906 7 1 2 16903 16905
0 16907 5 1 1 16906
0 16908 7 1 2 65628 16907
0 16909 5 1 1 16908
0 16910 7 2 2 42807 57609
0 16911 7 3 2 51662 56270
0 16912 7 1 2 65635 65637
0 16913 7 1 2 64493 16912
0 16914 5 1 1 16913
0 16915 7 1 2 16909 16914
0 16916 5 1 1 16915
0 16917 7 1 2 61160 16916
0 16918 5 1 1 16917
0 16919 7 1 2 46966 54165
0 16920 7 1 2 60434 64097
0 16921 7 1 2 16919 16920
0 16922 7 4 2 46913 57610
0 16923 7 5 2 48108 50351
0 16924 7 1 2 65640 65644
0 16925 7 1 2 16921 16924
0 16926 5 1 1 16925
0 16927 7 1 2 16918 16926
0 16928 5 1 1 16927
0 16929 7 1 2 45726 16928
0 16930 5 1 1 16929
0 16931 7 2 2 46494 65629
0 16932 7 1 2 61035 61664
0 16933 7 1 2 62999 16932
0 16934 7 1 2 65649 16933
0 16935 5 1 1 16934
0 16936 7 1 2 16930 16935
0 16937 5 1 1 16936
0 16938 7 1 2 45563 16937
0 16939 5 1 1 16938
0 16940 7 1 2 58090 61665
0 16941 7 1 2 65650 16940
0 16942 7 1 2 65572 16941
0 16943 5 1 1 16942
0 16944 7 1 2 16939 16943
0 16945 5 1 1 16944
0 16946 7 1 2 50263 16945
0 16947 5 1 1 16946
0 16948 7 1 2 42556 65553
0 16949 5 1 1 16948
0 16950 7 1 2 61886 65397
0 16951 5 1 1 16950
0 16952 7 1 2 16949 16951
0 16953 5 1 1 16952
0 16954 7 3 2 44444 62763
0 16955 7 1 2 42174 63000
0 16956 5 1 1 16955
0 16957 7 1 2 58997 62689
0 16958 5 1 1 16957
0 16959 7 1 2 16956 16958
0 16960 5 1 1 16959
0 16961 7 1 2 65651 16960
0 16962 5 1 1 16961
0 16963 7 2 2 47764 51817
0 16964 7 1 2 63008 64788
0 16965 7 1 2 65654 16964
0 16966 5 1 1 16965
0 16967 7 1 2 16962 16966
0 16968 5 1 1 16967
0 16969 7 1 2 43914 16968
0 16970 5 1 1 16969
0 16971 7 1 2 55456 55232
0 16972 7 1 2 65550 16971
0 16973 5 1 1 16972
0 16974 7 1 2 16970 16973
0 16975 5 1 1 16974
0 16976 7 1 2 45564 16975
0 16977 5 1 1 16976
0 16978 7 3 2 46833 44566
0 16979 7 1 2 53090 62499
0 16980 7 1 2 65656 16979
0 16981 7 1 2 65573 16980
0 16982 5 1 1 16981
0 16983 7 1 2 16977 16982
0 16984 5 1 1 16983
0 16985 7 1 2 16953 16984
0 16986 5 1 1 16985
0 16987 7 1 2 16947 16986
0 16988 5 1 1 16987
0 16989 7 1 2 58371 16988
0 16990 5 1 1 16989
0 16991 7 1 2 47645 16990
0 16992 7 1 2 16892 16991
0 16993 7 1 2 16673 16992
0 16994 5 1 1 16993
0 16995 7 1 2 44900 16994
0 16996 7 1 2 16083 16995
0 16997 5 1 1 16996
0 16998 7 7 2 59195 62500
0 16999 7 4 2 42275 61343
0 17000 7 1 2 64986 65666
0 17001 7 1 2 65659 17000
0 17002 7 1 2 45077 52961
0 17003 7 1 2 64749 17002
0 17004 7 1 2 58616 63317
0 17005 7 1 2 17003 17004
0 17006 7 1 2 17001 17005
0 17007 5 1 1 17006
0 17008 7 1 2 16997 17007
0 17009 7 1 2 13719 17008
0 17010 7 1 2 7042 17009
0 17011 5 1 1 17010
0 17012 7 1 2 48872 17011
0 17013 5 1 1 17012
0 17014 7 3 2 46997 44773
0 17015 5 1 1 65670
0 17016 7 1 2 50179 64139
0 17017 5 5 1 17016
0 17018 7 107 2 42276 44644
0 17019 5 8 1 65678
0 17020 7 1 2 65673 65679
0 17021 5 1 1 17020
0 17022 7 2 2 56345 64020
0 17023 5 1 1 65793
0 17024 7 1 2 46495 65794
0 17025 5 1 1 17024
0 17026 7 2 2 17021 17025
0 17027 5 1 1 65795
0 17028 7 1 2 53370 63680
0 17029 5 3 1 17028
0 17030 7 5 2 45808 61431
0 17031 5 1 1 65800
0 17032 7 1 2 65785 17031
0 17033 5 7 1 17032
0 17034 7 1 2 65797 65805
0 17035 5 1 1 17034
0 17036 7 4 2 47977 64299
0 17037 5 2 1 65812
0 17038 7 4 2 42277 58020
0 17039 5 2 1 65818
0 17040 7 1 2 65816 65822
0 17041 5 2 1 17040
0 17042 7 1 2 55580 65824
0 17043 5 1 1 17042
0 17044 7 1 2 17035 17043
0 17045 7 1 2 65796 17044
0 17046 5 1 1 17045
0 17047 7 1 2 55612 17046
0 17048 5 1 1 17047
0 17049 7 12 2 45809 43457
0 17050 7 3 2 47978 65486
0 17051 7 1 2 65826 65838
0 17052 5 1 1 17051
0 17053 7 1 2 17048 17052
0 17054 5 2 1 17053
0 17055 7 1 2 65671 65841
0 17056 5 1 1 17055
0 17057 7 3 2 43609 44445
0 17058 7 1 2 65827 65843
0 17059 7 1 2 61793 17058
0 17060 5 1 1 17059
0 17061 7 1 2 17056 17060
0 17062 5 1 1 17061
0 17063 7 1 2 45565 17062
0 17064 5 1 1 17063
0 17065 7 1 2 43610 7044
0 17066 5 1 1 17065
0 17067 7 1 2 46998 61175
0 17068 5 1 1 17067
0 17069 7 2 2 17066 17068
0 17070 7 1 2 63766 63723
0 17071 7 1 2 65846 17070
0 17072 5 1 1 17071
0 17073 7 1 2 17064 17072
0 17074 5 1 1 17073
0 17075 7 1 2 42363 17074
0 17076 5 1 1 17075
0 17077 7 15 2 45880 46999
0 17078 7 4 2 42278 65848
0 17079 5 1 1 65863
0 17080 7 4 2 50083 54764
0 17081 7 3 2 64534 65867
0 17082 7 1 2 65864 65871
0 17083 5 1 1 17082
0 17084 7 1 2 17076 17083
0 17085 5 1 1 17084
0 17086 7 1 2 46967 17085
0 17087 5 1 1 17086
0 17088 7 4 2 45881 43581
0 17089 7 5 2 47000 65874
0 17090 7 3 2 45810 65878
0 17091 7 1 2 65872 65883
0 17092 5 1 1 17091
0 17093 7 1 2 17087 17092
0 17094 5 1 1 17093
0 17095 7 1 2 46246 17094
0 17096 5 1 1 17095
0 17097 7 1 2 54765 58216
0 17098 7 3 2 46968 48862
0 17099 7 97 2 45811 47979
0 17100 5 1 1 65889
0 17101 7 1 2 65786 17100
0 17102 5 46 1 17101
0 17103 7 1 2 58590 65986
0 17104 7 1 2 65886 17103
0 17105 7 1 2 17097 17104
0 17106 5 1 1 17105
0 17107 7 1 2 17096 17106
0 17108 5 1 1 17107
0 17109 7 1 2 42175 17108
0 17110 5 1 1 17109
0 17111 7 12 2 42364 46247
0 17112 7 3 2 45727 66032
0 17113 7 28 2 43582 43611
0 17114 7 1 2 42279 66047
0 17115 7 1 2 66044 17114
0 17116 7 1 2 65873 17115
0 17117 5 1 1 17116
0 17118 7 1 2 17110 17117
0 17119 5 1 1 17118
0 17120 7 1 2 47646 17119
0 17121 5 1 1 17120
0 17122 7 2 2 47001 47549
0 17123 7 1 2 63808 66075
0 17124 7 1 2 60661 17123
0 17125 7 3 2 42365 49915
0 17126 7 2 2 61161 63728
0 17127 7 1 2 66077 66080
0 17128 7 1 2 17124 17127
0 17129 5 1 1 17128
0 17130 7 1 2 44567 17129
0 17131 7 1 2 17121 17130
0 17132 5 1 1 17131
0 17133 7 1 2 51228 58157
0 17134 5 1 1 17133
0 17135 7 1 2 50769 57611
0 17136 7 1 2 63704 17135
0 17137 5 1 1 17136
0 17138 7 1 2 17134 17137
0 17139 5 1 1 17138
0 17140 7 1 2 65987 17139
0 17141 5 1 1 17140
0 17142 7 5 2 45812 56346
0 17143 5 2 1 66082
0 17144 7 1 2 65787 66087
0 17145 5 7 1 17144
0 17146 7 1 2 55581 66089
0 17147 5 1 1 17146
0 17148 7 2 2 47980 64047
0 17149 5 1 1 66096
0 17150 7 1 2 58345 66097
0 17151 5 1 1 17150
0 17152 7 1 2 51796 65680
0 17153 5 1 1 17152
0 17154 7 1 2 17151 17153
0 17155 7 1 2 17147 17154
0 17156 5 1 1 17155
0 17157 7 1 2 58186 63953
0 17158 7 1 2 17156 17157
0 17159 5 1 1 17158
0 17160 7 1 2 17141 17159
0 17161 5 1 1 17160
0 17162 7 1 2 48863 17161
0 17163 5 1 1 17162
0 17164 7 4 2 47981 64021
0 17165 7 1 2 55898 66098
0 17166 5 1 1 17165
0 17167 7 4 2 42280 47765
0 17168 7 1 2 60020 61408
0 17169 7 1 2 66102 17168
0 17170 5 1 1 17169
0 17171 7 1 2 17166 17170
0 17172 5 1 1 17171
0 17173 7 1 2 49084 17172
0 17174 5 1 1 17173
0 17175 7 5 2 44645 49219
0 17176 7 2 2 63386 66106
0 17177 7 1 2 58083 66111
0 17178 5 1 1 17177
0 17179 7 2 2 44446 61432
0 17180 7 1 2 47550 65828
0 17181 7 1 2 66113 17180
0 17182 5 1 1 17181
0 17183 7 1 2 17178 17182
0 17184 7 1 2 17174 17183
0 17185 5 1 1 17184
0 17186 7 1 2 45566 17185
0 17187 5 1 1 17186
0 17188 7 2 2 61433 65499
0 17189 5 1 1 66115
0 17190 7 4 2 47982 49085
0 17191 7 1 2 64022 66117
0 17192 5 1 1 17191
0 17193 7 1 2 17189 17192
0 17194 5 1 1 17193
0 17195 7 1 2 60501 17194
0 17196 5 1 1 17195
0 17197 7 1 2 17187 17196
0 17198 5 1 1 17197
0 17199 7 1 2 48866 17198
0 17200 5 1 1 17199
0 17201 7 1 2 17163 17200
0 17202 5 1 1 17201
0 17203 7 1 2 46969 17202
0 17204 5 1 1 17203
0 17205 7 3 2 44646 65424
0 17206 7 1 2 43583 58187
0 17207 7 1 2 48873 17206
0 17208 7 1 2 66121 17207
0 17209 7 1 2 64374 17208
0 17210 5 1 1 17209
0 17211 7 1 2 17204 17210
0 17212 5 1 1 17211
0 17213 7 1 2 45728 17212
0 17214 5 1 1 17213
0 17215 7 1 2 48874 61986
0 17216 7 1 2 63792 17215
0 17217 7 1 2 51229 17216
0 17218 5 1 1 17217
0 17219 7 1 2 44774 17218
0 17220 7 1 2 17214 17219
0 17221 5 1 1 17220
0 17222 7 24 2 46970 47002
0 17223 5 2 1 66124
0 17224 7 13 2 45729 45882
0 17225 7 13 2 66125 66150
0 17226 7 4 2 43458 66163
0 17227 5 1 1 66176
0 17228 7 5 2 42366 43584
0 17229 7 14 2 43612 66180
0 17230 7 1 2 60675 66185
0 17231 5 1 1 17230
0 17232 7 1 2 17227 17231
0 17233 5 13 1 17232
0 17234 7 1 2 45567 66199
0 17235 5 1 1 17234
0 17236 7 6 2 47003 62902
0 17237 7 6 2 66151 66212
0 17238 7 3 2 42014 66218
0 17239 5 1 1 66224
0 17240 7 1 2 17235 17239
0 17241 5 8 1 17240
0 17242 7 1 2 45813 66227
0 17243 5 1 1 17242
0 17244 7 7 2 43585 47004
0 17245 7 5 2 45883 66235
0 17246 5 1 1 66242
0 17247 7 7 2 46971 43613
0 17248 7 2 2 42367 66247
0 17249 5 1 1 66254
0 17250 7 1 2 17246 17249
0 17251 5 31 1 17250
0 17252 7 2 2 42281 66256
0 17253 5 1 1 66287
0 17254 7 1 2 60683 66288
0 17255 5 1 1 17254
0 17256 7 1 2 17243 17255
0 17257 5 1 1 17256
0 17258 7 4 2 50770 53757
0 17259 5 4 1 66289
0 17260 7 2 2 61065 66293
0 17261 5 1 1 66297
0 17262 7 1 2 61835 66298
0 17263 5 12 1 17262
0 17264 7 1 2 57908 66299
0 17265 7 1 2 17257 17264
0 17266 5 1 1 17265
0 17267 7 1 2 58938 61265
0 17268 7 2 2 58372 17267
0 17269 7 1 2 45814 66257
0 17270 5 1 1 17269
0 17271 7 7 2 42282 45884
0 17272 7 1 2 66126 66313
0 17273 5 1 1 17272
0 17274 7 1 2 17270 17273
0 17275 5 4 1 17274
0 17276 7 1 2 60021 66320
0 17277 7 1 2 66311 17276
0 17278 5 1 1 17277
0 17279 7 1 2 48109 17278
0 17280 7 1 2 17266 17279
0 17281 5 1 1 17280
0 17282 7 1 2 61093 17281
0 17283 7 1 2 17221 17282
0 17284 5 1 1 17283
0 17285 7 1 2 65801 65887
0 17286 5 1 1 17285
0 17287 7 3 2 44647 60327
0 17288 7 2 2 48875 66324
0 17289 5 1 1 66327
0 17290 7 1 2 17286 17289
0 17291 5 1 1 17290
0 17292 7 2 2 49916 61904
0 17293 7 1 2 44775 61624
0 17294 7 1 2 66329 17293
0 17295 7 1 2 17291 17294
0 17296 5 1 1 17295
0 17297 7 1 2 47892 17296
0 17298 7 1 2 17284 17297
0 17299 5 1 1 17298
0 17300 7 1 2 17132 17299
0 17301 5 1 1 17300
0 17302 7 1 2 46914 17301
0 17303 5 1 1 17302
0 17304 7 7 2 45815 45885
0 17305 7 10 2 66127 66331
0 17306 5 1 1 66338
0 17307 7 3 2 51561 66300
0 17308 7 1 2 66339 66348
0 17309 5 1 1 17308
0 17310 7 2 2 50084 65988
0 17311 7 12 2 42368 66048
0 17312 7 1 2 44568 66353
0 17313 7 1 2 66351 17312
0 17314 5 1 1 17313
0 17315 7 1 2 17309 17314
0 17316 5 1 1 17315
0 17317 7 1 2 60684 17316
0 17318 5 1 1 17317
0 17319 7 2 2 44569 66128
0 17320 7 5 2 45886 43459
0 17321 7 1 2 66365 66367
0 17322 5 1 1 17321
0 17323 7 19 2 42369 43614
0 17324 7 1 2 54452 63382
0 17325 7 1 2 66372 17324
0 17326 5 1 1 17325
0 17327 7 1 2 17322 17326
0 17328 5 1 1 17327
0 17329 7 1 2 45568 17328
0 17330 5 1 1 17329
0 17331 7 5 2 42015 45887
0 17332 7 3 2 46834 66391
0 17333 7 1 2 66366 66396
0 17334 5 1 1 17333
0 17335 7 1 2 17330 17334
0 17336 5 1 1 17335
0 17337 7 1 2 50085 17336
0 17338 5 1 1 17337
0 17339 7 2 2 58077 66049
0 17340 7 3 2 45569 42370
0 17341 7 1 2 62845 66401
0 17342 7 1 2 66399 17341
0 17343 5 1 1 17342
0 17344 7 1 2 17338 17343
0 17345 5 1 1 17344
0 17346 7 1 2 65681 17345
0 17347 5 1 1 17346
0 17348 7 4 2 45816 44570
0 17349 7 6 2 44648 66404
0 17350 7 1 2 65868 66408
0 17351 5 1 1 17350
0 17352 7 3 2 46835 63017
0 17353 7 1 2 66349 66414
0 17354 5 1 1 17353
0 17355 7 1 2 17351 17354
0 17356 5 1 1 17355
0 17357 7 1 2 66258 17356
0 17358 5 1 1 17357
0 17359 7 1 2 63179 66354
0 17360 7 1 2 66350 17359
0 17361 5 1 1 17360
0 17362 7 1 2 17358 17361
0 17363 7 1 2 17347 17362
0 17364 5 1 1 17363
0 17365 7 1 2 45730 17364
0 17366 5 1 1 17365
0 17367 7 1 2 17318 17366
0 17368 5 1 1 17367
0 17369 7 1 2 48110 17368
0 17370 5 1 1 17369
0 17371 7 1 2 48876 58188
0 17372 7 1 2 61675 17371
0 17373 7 1 2 51230 63821
0 17374 7 1 2 17372 17373
0 17375 5 1 1 17374
0 17376 7 1 2 17370 17375
0 17377 5 1 1 17376
0 17378 7 1 2 46248 17377
0 17379 5 1 1 17378
0 17380 7 4 2 45450 65989
0 17381 7 3 2 42371 46496
0 17382 7 1 2 61020 66421
0 17383 7 1 2 62807 17382
0 17384 7 1 2 66400 17383
0 17385 7 1 2 66417 17384
0 17386 5 1 1 17385
0 17387 7 1 2 17379 17386
0 17388 5 1 1 17387
0 17389 7 1 2 59153 17388
0 17390 5 1 1 17389
0 17391 7 4 2 65890 66186
0 17392 7 1 2 60034 66424
0 17393 5 1 1 17392
0 17394 7 1 2 58290 66328
0 17395 5 1 1 17394
0 17396 7 1 2 17393 17395
0 17397 5 1 1 17396
0 17398 7 1 2 42176 17397
0 17399 5 1 1 17398
0 17400 7 1 2 48111 62754
0 17401 7 1 2 66425 17400
0 17402 5 1 1 17401
0 17403 7 1 2 17399 17402
0 17404 5 1 1 17403
0 17405 7 1 2 50267 60693
0 17406 7 1 2 17404 17405
0 17407 5 1 1 17406
0 17408 7 1 2 43530 17407
0 17409 7 1 2 17390 17408
0 17410 5 1 1 17409
0 17411 7 1 2 44901 17410
0 17412 7 1 2 17303 17411
0 17413 5 1 1 17412
0 17414 7 4 2 42372 44902
0 17415 7 1 2 63342 65839
0 17416 5 1 1 17415
0 17417 7 1 2 58939 62907
0 17418 7 1 2 66301 17417
0 17419 5 1 1 17418
0 17420 7 1 2 17416 17419
0 17421 5 1 1 17420
0 17422 7 1 2 42177 17421
0 17423 5 1 1 17422
0 17424 7 3 2 45817 51868
0 17425 5 1 1 66432
0 17426 7 1 2 66302 66433
0 17427 5 1 1 17426
0 17428 7 1 2 51784 5339
0 17429 5 2 1 17428
0 17430 7 5 2 46915 47983
0 17431 7 4 2 42283 66437
0 17432 5 1 1 66442
0 17433 7 1 2 60763 66443
0 17434 7 1 2 66435 17433
0 17435 5 1 1 17434
0 17436 7 1 2 62834 65618
0 17437 7 1 2 55582 17436
0 17438 5 1 1 17437
0 17439 7 1 2 17435 17438
0 17440 7 1 2 17427 17439
0 17441 5 1 1 17440
0 17442 7 1 2 55972 17441
0 17443 5 1 1 17442
0 17444 7 1 2 17423 17443
0 17445 5 1 1 17444
0 17446 7 1 2 46249 17445
0 17447 5 1 1 17446
0 17448 7 1 2 59977 63387
0 17449 7 1 2 66114 17448
0 17450 5 1 1 17449
0 17451 7 1 2 17447 17450
0 17452 5 1 1 17451
0 17453 7 1 2 66428 17452
0 17454 5 1 1 17453
0 17455 7 5 2 43304 47766
0 17456 7 1 2 55220 56119
0 17457 7 1 2 66446 17456
0 17458 7 4 2 45731 66314
0 17459 7 1 2 60704 66451
0 17460 7 1 2 17457 17459
0 17461 5 1 1 17460
0 17462 7 1 2 17454 17461
0 17463 5 1 1 17462
0 17464 7 1 2 46836 17463
0 17465 5 1 1 17464
0 17466 7 1 2 60726 66444
0 17467 5 1 1 17466
0 17468 7 2 2 57491 64300
0 17469 7 1 2 58021 66455
0 17470 5 1 1 17469
0 17471 7 1 2 17467 17470
0 17472 5 1 1 17471
0 17473 7 1 2 45732 17472
0 17474 5 1 1 17473
0 17475 7 1 2 42178 53741
0 17476 7 1 2 62468 62908
0 17477 7 2 2 17475 17476
0 17478 5 1 1 66457
0 17479 7 1 2 17474 17478
0 17480 5 1 1 17479
0 17481 7 1 2 46682 17480
0 17482 5 1 1 17481
0 17483 7 7 2 42284 47551
0 17484 7 1 2 57593 58888
0 17485 7 2 2 66459 17484
0 17486 5 1 1 66466
0 17487 7 1 2 17482 17486
0 17488 5 1 1 17487
0 17489 7 9 2 42373 43460
0 17490 7 1 2 57682 66468
0 17491 7 1 2 17488 17490
0 17492 5 1 1 17491
0 17493 7 1 2 17465 17492
0 17494 5 1 1 17493
0 17495 7 1 2 44571 17494
0 17496 5 1 1 17495
0 17497 7 1 2 51231 57809
0 17498 5 1 1 17497
0 17499 7 1 2 55800 55973
0 17500 7 1 2 62299 17499
0 17501 5 1 1 17500
0 17502 7 1 2 17498 17501
0 17503 5 1 1 17502
0 17504 7 15 2 45818 46250
0 17505 7 4 2 50352 66477
0 17506 7 1 2 66429 66492
0 17507 7 1 2 17503 17506
0 17508 5 1 1 17507
0 17509 7 1 2 17496 17508
0 17510 5 1 1 17509
0 17511 7 1 2 45570 17510
0 17512 5 1 1 17511
0 17513 7 18 2 45819 50353
0 17514 5 1 1 66496
0 17515 7 1 2 65328 66497
0 17516 5 1 1 17515
0 17517 7 12 2 42285 48932
0 17518 5 3 1 66514
0 17519 7 1 2 60727 66515
0 17520 5 1 1 17519
0 17521 7 1 2 17516 17520
0 17522 5 1 1 17521
0 17523 7 1 2 46916 17522
0 17524 5 1 1 17523
0 17525 7 5 2 44572 58022
0 17526 7 1 2 66456 66529
0 17527 5 1 1 17526
0 17528 7 1 2 17524 17527
0 17529 5 1 1 17528
0 17530 7 1 2 46683 17529
0 17531 5 1 1 17530
0 17532 7 3 2 47552 57594
0 17533 7 29 2 47984 64713
0 17534 5 2 1 66537
0 17535 7 11 2 45820 47893
0 17536 7 2 2 58023 66568
0 17537 5 1 1 66579
0 17538 7 2 2 66566 17537
0 17539 5 4 1 66581
0 17540 7 1 2 66534 66583
0 17541 5 1 1 17540
0 17542 7 1 2 17531 17541
0 17543 5 1 1 17542
0 17544 7 1 2 45733 17543
0 17545 5 1 1 17544
0 17546 7 8 2 46684 44573
0 17547 7 1 2 66458 66587
0 17548 5 1 1 17547
0 17549 7 1 2 17545 17548
0 17550 5 1 1 17549
0 17551 7 1 2 60502 66430
0 17552 7 1 2 17550 17551
0 17553 5 1 1 17552
0 17554 7 1 2 17512 17553
0 17555 5 1 1 17554
0 17556 7 1 2 47647 17555
0 17557 5 1 1 17556
0 17558 7 1 2 42179 56970
0 17559 5 1 1 17558
0 17560 7 1 2 43531 62755
0 17561 5 1 1 17560
0 17562 7 1 2 17559 17561
0 17563 5 1 1 17562
0 17564 7 1 2 54766 17563
0 17565 5 1 1 17564
0 17566 7 1 2 53644 61816
0 17567 5 1 1 17566
0 17568 7 1 2 17565 17567
0 17569 5 2 1 17568
0 17570 7 3 2 42286 50771
0 17571 7 3 2 47767 44903
0 17572 7 1 2 59674 66600
0 17573 7 1 2 66422 17572
0 17574 7 1 2 66597 17573
0 17575 7 1 2 66595 17574
0 17576 5 1 1 17575
0 17577 7 1 2 17557 17576
0 17578 5 1 1 17577
0 17579 7 6 2 43586 48112
0 17580 5 1 1 66603
0 17581 7 4 2 43615 44776
0 17582 5 3 1 66609
0 17583 7 1 2 66613 66148
0 17584 7 1 2 17580 17583
0 17585 7 1 2 17578 17584
0 17586 5 1 1 17585
0 17587 7 2 2 43616 48113
0 17588 5 1 1 66616
0 17589 7 3 2 17015 17588
0 17590 7 2 2 58050 66303
0 17591 5 1 1 66621
0 17592 7 1 2 58426 62300
0 17593 5 1 1 17592
0 17594 7 1 2 17591 17593
0 17595 5 1 1 17594
0 17596 7 1 2 47768 17595
0 17597 5 1 1 17596
0 17598 7 2 2 51728 61050
0 17599 5 1 1 66623
0 17600 7 1 2 43532 66624
0 17601 5 1 1 17600
0 17602 7 1 2 17597 17601
0 17603 5 1 1 17602
0 17604 7 2 2 45888 46251
0 17605 7 1 2 54432 66625
0 17606 7 1 2 17603 17605
0 17607 5 1 1 17606
0 17608 7 11 2 44213 47985
0 17609 7 1 2 58735 60416
0 17610 7 1 2 66627 17609
0 17611 7 4 2 42374 42808
0 17612 7 3 2 45734 66638
0 17613 7 9 2 43305 46917
0 17614 7 2 2 43085 66645
0 17615 7 1 2 66642 66654
0 17616 7 1 2 17610 17615
0 17617 5 1 1 17616
0 17618 7 1 2 17607 17617
0 17619 5 1 1 17618
0 17620 7 1 2 58189 17619
0 17621 5 1 1 17620
0 17622 7 1 2 51663 65329
0 17623 5 1 1 17622
0 17624 7 2 2 51587 53742
0 17625 5 1 1 66656
0 17626 7 1 2 47553 66657
0 17627 5 1 1 17626
0 17628 7 1 2 17623 17627
0 17629 5 1 1 17628
0 17630 7 1 2 45735 17629
0 17631 5 1 1 17630
0 17632 7 1 2 57239 65380
0 17633 5 1 1 17632
0 17634 7 1 2 17631 17633
0 17635 5 1 1 17634
0 17636 7 1 2 46685 17635
0 17637 5 1 1 17636
0 17638 7 1 2 62756 66535
0 17639 5 1 1 17638
0 17640 7 1 2 17637 17639
0 17641 5 1 1 17640
0 17642 7 5 2 45889 44649
0 17643 7 1 2 57683 66658
0 17644 7 1 2 54767 17643
0 17645 7 1 2 17641 17644
0 17646 5 1 1 17645
0 17647 7 1 2 17621 17646
0 17648 5 1 1 17647
0 17649 7 1 2 60328 17648
0 17650 5 1 1 17649
0 17651 7 1 2 62308 65551
0 17652 5 1 1 17651
0 17653 7 1 2 62304 64378
0 17654 5 3 1 17653
0 17655 7 1 2 65430 66663
0 17656 5 1 1 17655
0 17657 7 1 2 16488 17656
0 17658 5 1 1 17657
0 17659 7 1 2 42180 17658
0 17660 5 1 1 17659
0 17661 7 1 2 47769 65569
0 17662 7 1 2 66664 17661
0 17663 5 1 1 17662
0 17664 7 1 2 17660 17663
0 17665 5 1 1 17664
0 17666 7 1 2 44574 17665
0 17667 5 1 1 17666
0 17668 7 1 2 17652 17667
0 17669 5 1 1 17668
0 17670 7 1 2 58190 17669
0 17671 5 1 1 17670
0 17672 7 1 2 58206 65487
0 17673 7 1 2 65579 17672
0 17674 5 1 1 17673
0 17675 7 1 2 17671 17674
0 17676 5 1 1 17675
0 17677 7 1 2 46252 48917
0 17678 7 1 2 17676 17677
0 17679 5 1 1 17678
0 17680 7 1 2 54768 65574
0 17681 5 1 1 17680
0 17682 7 2 2 62708 65536
0 17683 7 1 2 58191 66666
0 17684 5 1 1 17683
0 17685 7 1 2 17681 17684
0 17686 5 1 1 17685
0 17687 7 1 2 57377 65652
0 17688 7 1 2 17686 17687
0 17689 5 1 1 17688
0 17690 7 1 2 17679 17689
0 17691 5 1 1 17690
0 17692 7 2 2 45890 47986
0 17693 7 1 2 44904 66668
0 17694 7 1 2 17691 17693
0 17695 5 1 1 17694
0 17696 7 1 2 17650 17695
0 17697 5 1 1 17696
0 17698 7 1 2 47648 17697
0 17699 5 1 1 17698
0 17700 7 3 2 42287 61021
0 17701 7 1 2 63420 66670
0 17702 5 1 1 17701
0 17703 7 1 2 60315 11274
0 17704 5 1 1 17703
0 17705 7 3 2 42181 46972
0 17706 5 1 1 66673
0 17707 7 1 2 42016 4775
0 17708 7 1 2 17706 17707
0 17709 7 1 2 17704 17708
0 17710 5 1 1 17709
0 17711 7 1 2 17702 17710
0 17712 5 1 1 17711
0 17713 7 1 2 56971 17712
0 17714 5 1 1 17713
0 17715 7 1 2 53628 56955
0 17716 5 1 1 17715
0 17717 7 1 2 57511 17716
0 17718 5 6 1 17717
0 17719 7 1 2 42017 66676
0 17720 5 1 1 17719
0 17721 7 1 2 53691 61285
0 17722 5 1 1 17721
0 17723 7 1 2 17720 17722
0 17724 5 1 1 17723
0 17725 7 1 2 63822 17724
0 17726 5 1 1 17725
0 17727 7 1 2 17714 17726
0 17728 5 1 1 17727
0 17729 7 5 2 45891 47770
0 17730 7 1 2 47987 61926
0 17731 7 1 2 66682 17730
0 17732 7 1 2 58852 17731
0 17733 7 1 2 17728 17732
0 17734 5 1 1 17733
0 17735 7 1 2 17699 17734
0 17736 5 1 1 17735
0 17737 7 1 2 66618 17736
0 17738 5 1 1 17737
0 17739 7 1 2 46253 65842
0 17740 5 1 1 17739
0 17741 7 4 2 44447 65990
0 17742 7 2 2 55409 60722
0 17743 7 1 2 66687 66691
0 17744 5 1 1 17743
0 17745 7 1 2 17740 17744
0 17746 5 1 1 17745
0 17747 7 1 2 45571 17746
0 17748 5 1 1 17747
0 17749 7 1 2 46254 50086
0 17750 5 3 1 17749
0 17751 7 1 2 5285 66693
0 17752 5 7 1 17751
0 17753 7 1 2 65891 66696
0 17754 5 1 1 17753
0 17755 7 2 2 53743 65682
0 17756 5 1 1 66703
0 17757 7 1 2 50772 66704
0 17758 5 1 1 17757
0 17759 7 1 2 17754 17758
0 17760 5 1 1 17759
0 17761 7 1 2 58091 17760
0 17762 5 1 1 17761
0 17763 7 1 2 17748 17762
0 17764 5 1 1 17763
0 17765 7 1 2 60566 17764
0 17766 5 1 1 17765
0 17767 7 3 2 44448 50354
0 17768 7 2 2 51526 66705
0 17769 7 4 2 45572 56872
0 17770 7 1 2 65537 66710
0 17771 7 1 2 66708 17770
0 17772 5 1 1 17771
0 17773 7 1 2 17766 17772
0 17774 5 1 1 17773
0 17775 7 1 2 66431 17774
0 17776 5 1 1 17775
0 17777 7 1 2 46837 57703
0 17778 7 1 2 57784 66628
0 17779 7 1 2 17777 17778
0 17780 7 4 2 45892 42809
0 17781 7 2 2 51339 66714
0 17782 7 7 2 45573 63796
0 17783 7 1 2 66718 66720
0 17784 7 1 2 17779 17783
0 17785 5 1 1 17784
0 17786 7 1 2 17776 17785
0 17787 5 1 1 17786
0 17788 7 1 2 47649 17787
0 17789 5 1 1 17788
0 17790 7 1 2 42018 62568
0 17791 5 1 1 17790
0 17792 7 1 2 61022 61286
0 17793 5 1 1 17792
0 17794 7 1 2 17791 17793
0 17795 5 1 1 17794
0 17796 7 10 2 45821 42375
0 17797 7 2 2 59675 66727
0 17798 7 1 2 58853 63954
0 17799 7 1 2 66737 17798
0 17800 7 1 2 17795 17799
0 17801 5 1 1 17800
0 17802 7 1 2 17789 17801
0 17803 5 1 1 17802
0 17804 7 3 2 46973 48114
0 17805 5 2 1 66739
0 17806 7 2 2 9826 66742
0 17807 7 4 2 46918 47005
0 17808 5 1 1 66746
0 17809 7 1 2 66614 17808
0 17810 7 1 2 66744 17809
0 17811 7 1 2 17803 17810
0 17812 5 1 1 17811
0 17813 7 5 2 43086 44777
0 17814 7 2 2 60897 66750
0 17815 7 1 2 50202 61023
0 17816 7 1 2 66755 17815
0 17817 7 3 2 48933 64074
0 17818 7 3 2 43306 55801
0 17819 7 1 2 66757 66760
0 17820 7 1 2 66340 17819
0 17821 7 1 2 17816 17820
0 17822 5 1 1 17821
0 17823 7 1 2 17812 17822
0 17824 7 1 2 17738 17823
0 17825 7 1 2 17586 17824
0 17826 7 1 2 17413 17825
0 17827 5 1 1 17826
0 17828 7 1 2 54279 17827
0 17829 5 1 1 17828
0 17830 7 2 2 50697 54621
0 17831 5 2 1 66763
0 17832 7 4 2 54074 65174
0 17833 5 2 1 66767
0 17834 7 1 2 66765 66771
0 17835 5 4 1 17834
0 17836 7 1 2 50773 66498
0 17837 5 1 1 17836
0 17838 7 1 2 66582 17837
0 17839 5 1 1 17838
0 17840 7 2 2 65488 17839
0 17841 7 1 2 58124 66777
0 17842 5 1 1 17841
0 17843 7 1 2 53639 66778
0 17844 5 1 1 17843
0 17845 7 2 2 47988 49220
0 17846 7 4 2 44575 63388
0 17847 7 1 2 66779 66781
0 17848 5 1 1 17847
0 17849 7 1 2 17514 66526
0 17850 5 11 1 17849
0 17851 7 1 2 59065 66785
0 17852 5 1 1 17851
0 17853 7 1 2 17848 17852
0 17854 5 1 1 17853
0 17855 7 1 2 55613 17854
0 17856 5 1 1 17855
0 17857 7 1 2 49086 66499
0 17858 5 1 1 17857
0 17859 7 1 2 66527 17858
0 17860 5 1 1 17859
0 17861 7 1 2 55899 17860
0 17862 5 1 1 17861
0 17863 7 1 2 17856 17862
0 17864 5 1 1 17863
0 17865 7 1 2 46686 17864
0 17866 5 1 1 17865
0 17867 7 2 2 43307 55614
0 17868 5 1 1 66796
0 17869 7 1 2 62269 66516
0 17870 7 1 2 66797 17869
0 17871 5 1 1 17870
0 17872 7 2 2 43461 57962
0 17873 5 1 1 66798
0 17874 7 1 2 66584 66799
0 17875 5 1 1 17874
0 17876 7 1 2 17871 17875
0 17877 7 1 2 17866 17876
0 17878 5 1 1 17877
0 17879 7 1 2 53305 17878
0 17880 5 1 1 17879
0 17881 7 1 2 17844 17880
0 17882 5 1 1 17881
0 17883 7 1 2 45574 17882
0 17884 5 1 1 17883
0 17885 7 1 2 17842 17884
0 17886 5 1 1 17885
0 17887 7 1 2 42810 17886
0 17888 5 1 1 17887
0 17889 7 1 2 58145 58373
0 17890 5 1 1 17889
0 17891 7 1 2 58766 58113
0 17892 7 1 2 63480 17891
0 17893 5 1 1 17892
0 17894 7 1 2 17890 17893
0 17895 5 1 1 17894
0 17896 7 1 2 43087 66517
0 17897 7 1 2 17895 17896
0 17898 5 1 1 17897
0 17899 7 1 2 17888 17898
0 17900 5 1 1 17899
0 17901 7 1 2 47650 17900
0 17902 5 1 1 17901
0 17903 7 4 2 45822 44449
0 17904 7 4 2 50355 66800
0 17905 7 1 2 59460 66804
0 17906 5 1 1 17905
0 17907 7 2 2 56173 59034
0 17908 5 1 1 66808
0 17909 7 1 2 66538 66809
0 17910 5 1 1 17909
0 17911 7 1 2 17906 17910
0 17912 5 1 1 17911
0 17913 7 1 2 44322 17912
0 17914 5 2 1 17913
0 17915 7 1 2 62118 65467
0 17916 5 5 1 17915
0 17917 7 4 2 54499 59154
0 17918 7 12 2 45823 66817
0 17919 7 1 2 66812 66821
0 17920 5 1 1 17919
0 17921 7 3 2 47989 60177
0 17922 7 9 2 66103 66833
0 17923 7 1 2 59101 66836
0 17924 5 2 1 17923
0 17925 7 1 2 17920 66845
0 17926 5 1 1 17925
0 17927 7 1 2 54769 17926
0 17928 5 1 1 17927
0 17929 7 2 2 58986 60228
0 17930 7 1 2 55457 66847
0 17931 5 1 1 17930
0 17932 7 3 2 44214 59840
0 17933 5 1 1 66849
0 17934 7 1 2 17931 17933
0 17935 5 1 1 17934
0 17936 7 1 2 43308 17935
0 17937 5 1 1 17936
0 17938 7 5 2 55458 59567
0 17939 7 3 2 46687 66852
0 17940 7 1 2 58352 8199
0 17941 5 3 1 17940
0 17942 7 1 2 66857 66860
0 17943 5 1 1 17942
0 17944 7 2 2 17937 17943
0 17945 5 1 1 66863
0 17946 7 6 2 42288 47894
0 17947 7 4 2 57909 66865
0 17948 5 2 1 66871
0 17949 7 7 2 58940 66405
0 17950 5 1 1 66877
0 17951 7 1 2 66875 17950
0 17952 5 10 1 17951
0 17953 7 1 2 17945 66884
0 17954 5 1 1 17953
0 17955 7 2 2 58192 63937
0 17956 7 5 2 47651 66894
0 17957 5 1 1 66896
0 17958 7 1 2 66897 66885
0 17959 5 1 1 17958
0 17960 7 2 2 59196 64679
0 17961 7 1 2 58836 66901
0 17962 5 1 1 17961
0 17963 7 1 2 17959 17962
0 17964 5 1 1 17963
0 17965 7 1 2 50841 17964
0 17966 5 1 1 17965
0 17967 7 1 2 17954 17966
0 17968 7 1 2 17928 17967
0 17969 5 1 1 17968
0 17970 7 1 2 53586 17969
0 17971 5 1 1 17970
0 17972 7 1 2 66810 17971
0 17973 7 1 2 17902 17972
0 17974 5 1 1 17973
0 17975 7 1 2 66259 17974
0 17976 5 1 1 17975
0 17977 7 4 2 45893 46919
0 17978 5 1 1 66903
0 17979 7 6 2 66213 66904
0 17980 7 12 2 47652 66907
0 17981 7 1 2 59284 65798
0 17982 5 1 1 17981
0 17983 7 2 2 51935 63684
0 17984 5 1 1 66925
0 17985 7 1 2 17982 17984
0 17986 5 1 1 17985
0 17987 7 1 2 45451 17986
0 17988 5 1 1 17987
0 17989 7 1 2 55201 64764
0 17990 5 1 1 17989
0 17991 7 1 2 17988 17990
0 17992 5 1 1 17991
0 17993 7 1 2 42811 17992
0 17994 5 1 1 17993
0 17995 7 1 2 62820 65349
0 17996 5 1 1 17995
0 17997 7 1 2 17994 17996
0 17998 5 1 1 17997
0 17999 7 1 2 66913 17998
0 18000 5 1 1 17999
0 18001 7 2 2 52297 59285
0 18002 5 1 1 66927
0 18003 7 1 2 51936 64552
0 18004 5 1 1 18003
0 18005 7 1 2 18002 18004
0 18006 5 1 1 18005
0 18007 7 3 2 43533 66050
0 18008 7 2 2 42376 59197
0 18009 7 1 2 66929 66932
0 18010 7 1 2 18006 18009
0 18011 5 1 1 18010
0 18012 7 1 2 18000 18011
0 18013 5 1 1 18012
0 18014 7 1 2 60449 18013
0 18015 5 1 1 18014
0 18016 7 1 2 51937 66290
0 18017 5 1 1 18016
0 18018 7 1 2 63658 18017
0 18019 5 1 1 18018
0 18020 7 1 2 42812 18019
0 18021 5 1 1 18020
0 18022 7 2 2 49840 50288
0 18023 5 1 1 66934
0 18024 7 1 2 59286 66935
0 18025 5 1 1 18024
0 18026 7 1 2 18021 18025
0 18027 5 1 1 18026
0 18028 7 1 2 66914 18027
0 18029 5 1 1 18028
0 18030 7 6 2 45736 42377
0 18031 7 3 2 66051 66936
0 18032 5 1 1 66942
0 18033 7 7 2 55959 59198
0 18034 5 4 1 66945
0 18035 7 4 2 66943 66946
0 18036 5 1 1 66956
0 18037 7 1 2 49983 66957
0 18038 5 1 1 18037
0 18039 7 1 2 18029 18038
0 18040 5 1 1 18039
0 18041 7 1 2 62501 18040
0 18042 5 1 1 18041
0 18043 7 1 2 18015 18042
0 18044 5 1 1 18043
0 18045 7 1 2 65892 18044
0 18046 5 1 1 18045
0 18047 7 2 2 60613 66813
0 18048 5 1 1 66960
0 18049 7 1 2 65991 66961
0 18050 5 1 1 18049
0 18051 7 5 2 60178 64539
0 18052 7 1 2 63729 66962
0 18053 7 1 2 59102 18052
0 18054 5 2 1 18053
0 18055 7 1 2 18050 66967
0 18056 5 1 1 18055
0 18057 7 1 2 54770 18056
0 18058 5 1 1 18057
0 18059 7 6 2 42289 57940
0 18060 5 2 1 66969
0 18061 7 3 2 43088 65893
0 18062 5 3 1 66977
0 18063 7 1 2 66975 66980
0 18064 5 3 1 18063
0 18065 7 1 2 59841 66983
0 18066 5 1 1 18065
0 18067 7 5 2 42290 42813
0 18068 7 2 2 45575 66986
0 18069 7 1 2 60022 64427
0 18070 7 1 2 66991 18069
0 18071 5 1 1 18070
0 18072 7 1 2 18066 18071
0 18073 5 1 1 18072
0 18074 7 1 2 58721 18073
0 18075 5 1 1 18074
0 18076 7 2 2 57910 66569
0 18077 7 1 2 56200 59822
0 18078 7 1 2 66993 18077
0 18079 5 1 1 18078
0 18080 7 1 2 18075 18079
0 18081 5 1 1 18080
0 18082 7 1 2 50842 18081
0 18083 5 1 1 18082
0 18084 7 1 2 18058 18083
0 18085 7 1 2 58024 66460
0 18086 5 3 1 18085
0 18087 7 1 2 64301 66118
0 18088 5 1 1 18087
0 18089 7 1 2 66995 18088
0 18090 5 1 1 18089
0 18091 7 1 2 66853 18090
0 18092 5 1 1 18091
0 18093 7 1 2 61753 65894
0 18094 5 1 1 18093
0 18095 7 1 2 59842 66090
0 18096 5 1 1 18095
0 18097 7 1 2 18094 18096
0 18098 5 1 1 18097
0 18099 7 1 2 44215 18098
0 18100 5 1 1 18099
0 18101 7 1 2 18092 18100
0 18102 5 1 1 18101
0 18103 7 1 2 43309 18102
0 18104 5 1 1 18103
0 18105 7 1 2 45824 49514
0 18106 5 1 1 18105
0 18107 7 1 2 60724 65992
0 18108 7 1 2 18106 18107
0 18109 7 1 2 44216 4672
0 18110 7 1 2 9976 18109
0 18111 5 1 1 18110
0 18112 7 1 2 66858 18111
0 18113 7 1 2 18108 18112
0 18114 5 1 1 18113
0 18115 7 1 2 18104 18114
0 18116 5 1 1 18115
0 18117 7 1 2 58722 18116
0 18118 5 1 1 18117
0 18119 7 1 2 65993 66850
0 18120 5 1 1 18119
0 18121 7 3 2 61434 63112
0 18122 7 1 2 58896 59479
0 18123 7 1 2 66998 18122
0 18124 5 1 1 18123
0 18125 7 1 2 18120 18124
0 18126 5 1 1 18125
0 18127 7 1 2 43310 18126
0 18128 5 1 1 18127
0 18129 7 1 2 65895 66861
0 18130 5 1 1 18129
0 18131 7 2 2 49087 65683
0 18132 5 3 1 67001
0 18133 7 1 2 18130 67003
0 18134 5 1 1 18133
0 18135 7 1 2 46688 18134
0 18136 5 1 1 18135
0 18137 7 1 2 66996 18136
0 18138 5 1 1 18137
0 18139 7 1 2 66854 18138
0 18140 5 1 1 18139
0 18141 7 1 2 18128 18140
0 18142 5 1 1 18141
0 18143 7 1 2 61051 18142
0 18144 5 1 1 18143
0 18145 7 1 2 18118 18144
0 18146 7 1 2 18084 18145
0 18147 5 1 1 18146
0 18148 7 2 2 62674 65849
0 18149 5 1 1 67006
0 18150 7 1 2 46920 66355
0 18151 5 1 1 18150
0 18152 7 1 2 18149 18151
0 18153 5 30 1 18152
0 18154 7 1 2 18147 67008
0 18155 5 1 1 18154
0 18156 7 1 2 53629 66187
0 18157 5 1 1 18156
0 18158 7 4 2 46921 66129
0 18159 7 1 2 66368 67038
0 18160 5 1 1 18159
0 18161 7 1 2 18157 18160
0 18162 5 14 1 18161
0 18163 7 1 2 49461 63576
0 18164 5 1 1 18163
0 18165 7 1 2 43089 63639
0 18166 5 1 1 18165
0 18167 7 1 2 18164 18166
0 18168 5 1 1 18167
0 18169 7 1 2 43311 18168
0 18170 5 1 1 18169
0 18171 7 3 2 42019 60179
0 18172 7 1 2 65655 67056
0 18173 5 1 1 18172
0 18174 7 1 2 63964 65257
0 18175 5 1 1 18174
0 18176 7 2 2 44450 18175
0 18177 7 1 2 59568 67059
0 18178 5 1 1 18177
0 18179 7 1 2 18173 18178
0 18180 5 1 1 18179
0 18181 7 1 2 55583 18180
0 18182 5 1 1 18181
0 18183 7 1 2 58614 64259
0 18184 5 1 1 18183
0 18185 7 1 2 63659 18184
0 18186 5 1 1 18185
0 18187 7 1 2 60490 18186
0 18188 5 1 1 18187
0 18189 7 1 2 49515 57747
0 18190 7 1 2 61625 18189
0 18191 5 1 1 18190
0 18192 7 1 2 18188 18191
0 18193 7 1 2 18182 18192
0 18194 7 1 2 18170 18193
0 18195 5 1 1 18194
0 18196 7 1 2 65896 18195
0 18197 5 1 1 18196
0 18198 7 2 2 59287 66814
0 18199 5 2 1 67061
0 18200 7 1 2 57989 65248
0 18201 5 1 1 18200
0 18202 7 1 2 67063 18201
0 18203 5 1 1 18202
0 18204 7 4 2 61357 63018
0 18205 7 1 2 18203 67065
0 18206 5 1 1 18205
0 18207 7 7 2 47554 55378
0 18208 5 1 1 67069
0 18209 7 2 2 60687 61266
0 18210 7 1 2 67070 67076
0 18211 5 1 1 18210
0 18212 7 1 2 61647 64243
0 18213 5 1 1 18212
0 18214 7 1 2 18211 18213
0 18215 5 1 1 18214
0 18216 7 1 2 66091 18215
0 18217 5 1 1 18216
0 18218 7 1 2 18206 18217
0 18219 7 1 2 18197 18218
0 18220 5 1 1 18219
0 18221 7 1 2 67042 18220
0 18222 5 1 1 18221
0 18223 7 5 2 59288 60450
0 18224 7 1 2 63938 66915
0 18225 5 1 1 18224
0 18226 7 4 2 42378 55756
0 18227 7 12 2 66052 67083
0 18228 7 1 2 59464 67087
0 18229 5 1 1 18228
0 18230 7 1 2 18225 18229
0 18231 5 1 1 18230
0 18232 7 1 2 65684 18231
0 18233 5 1 1 18232
0 18234 7 3 2 55860 62709
0 18235 7 1 2 43617 66738
0 18236 7 1 2 67099 18235
0 18237 5 1 1 18236
0 18238 7 1 2 18233 18237
0 18239 5 1 1 18238
0 18240 7 1 2 67078 18239
0 18241 5 1 1 18240
0 18242 7 1 2 64277 66984
0 18243 5 1 1 18242
0 18244 7 2 2 47653 60914
0 18245 7 1 2 61233 67102
0 18246 7 1 2 66994 18245
0 18247 5 1 1 18246
0 18248 7 1 2 18243 18247
0 18249 5 1 1 18248
0 18250 7 1 2 67043 18249
0 18251 5 1 1 18250
0 18252 7 2 2 63797 64495
0 18253 7 1 2 55733 60494
0 18254 7 1 2 66908 18253
0 18255 7 1 2 67104 18254
0 18256 5 1 1 18255
0 18257 7 1 2 18251 18256
0 18258 7 1 2 18241 18257
0 18259 5 1 1 18258
0 18260 7 1 2 50843 18259
0 18261 5 1 1 18260
0 18262 7 3 2 60451 65261
0 18263 5 1 1 67106
0 18264 7 1 2 63939 67107
0 18265 5 1 1 18264
0 18266 7 1 2 42020 67060
0 18267 5 1 1 18266
0 18268 7 1 2 18265 18267
0 18269 5 1 1 18268
0 18270 7 1 2 65897 18269
0 18271 5 1 1 18270
0 18272 7 3 2 59289 65685
0 18273 7 1 2 42814 63705
0 18274 5 1 1 18273
0 18275 7 1 2 2971 18274
0 18276 5 1 1 18275
0 18277 7 1 2 67109 18276
0 18278 5 1 1 18277
0 18279 7 1 2 18271 18278
0 18280 5 1 1 18279
0 18281 7 1 2 18280 66916
0 18282 5 1 1 18281
0 18283 7 3 2 42379 55861
0 18284 7 11 2 43618 62710
0 18285 7 3 2 67112 67115
0 18286 7 1 2 66721 66963
0 18287 7 1 2 67126 18286
0 18288 5 1 1 18287
0 18289 7 1 2 18282 18288
0 18290 5 1 1 18289
0 18291 7 1 2 55584 18290
0 18292 5 1 1 18291
0 18293 7 1 2 45894 63134
0 18294 7 7 2 47654 66130
0 18295 7 1 2 65641 67129
0 18296 7 1 2 18293 18295
0 18297 5 1 1 18296
0 18298 7 1 2 18036 18297
0 18299 5 1 1 18298
0 18300 7 1 2 62502 18299
0 18301 5 1 1 18300
0 18302 7 3 2 61024 66356
0 18303 5 1 1 67136
0 18304 7 1 2 57631 63187
0 18305 7 1 2 67137 18304
0 18306 5 1 1 18305
0 18307 7 1 2 18301 18306
0 18308 5 1 1 18307
0 18309 7 1 2 49984 18308
0 18310 5 1 1 18309
0 18311 7 1 2 60452 63678
0 18312 5 1 1 18311
0 18313 7 1 2 11161 18312
0 18314 5 1 1 18313
0 18315 7 1 2 64235 18314
0 18316 5 1 1 18315
0 18317 7 2 2 48809 67079
0 18318 5 1 1 67139
0 18319 7 1 2 64128 18318
0 18320 5 1 1 18319
0 18321 7 1 2 50774 18320
0 18322 5 1 1 18321
0 18323 7 1 2 18316 18322
0 18324 5 1 1 18323
0 18325 7 4 2 62903 66747
0 18326 7 2 2 66715 67141
0 18327 7 1 2 47655 67145
0 18328 7 1 2 18324 18327
0 18329 5 1 1 18328
0 18330 7 1 2 18310 18329
0 18331 5 1 1 18330
0 18332 7 1 2 65686 18331
0 18333 5 1 1 18332
0 18334 7 1 2 18292 18333
0 18335 7 1 2 18261 18334
0 18336 7 1 2 18222 18335
0 18337 7 1 2 18155 18336
0 18338 7 1 2 18046 18337
0 18339 7 1 2 17976 18338
0 18340 5 1 1 18339
0 18341 7 1 2 66773 18340
0 18342 5 1 1 18341
0 18343 7 3 2 44650 57028
0 18344 7 2 2 43534 48432
0 18345 7 2 2 60055 67150
0 18346 7 1 2 62272 67152
0 18347 5 1 1 18346
0 18348 7 1 2 49430 55808
0 18349 7 1 2 67103 18348
0 18350 5 1 1 18349
0 18351 7 1 2 18347 18350
0 18352 5 1 1 18351
0 18353 7 1 2 48233 58406
0 18354 7 1 2 18352 18353
0 18355 5 1 1 18354
0 18356 7 1 2 54827 63663
0 18357 7 1 2 65175 18356
0 18358 7 1 2 58358 60238
0 18359 7 1 2 18357 18358
0 18360 5 1 1 18359
0 18361 7 1 2 18355 18360
0 18362 5 1 1 18361
0 18363 7 1 2 45576 18362
0 18364 5 1 1 18363
0 18365 7 6 2 53672 59362
0 18366 7 1 2 62273 66764
0 18367 7 1 2 67154 18366
0 18368 5 1 1 18367
0 18369 7 1 2 18364 18368
0 18370 5 1 1 18369
0 18371 7 1 2 43312 18370
0 18372 5 1 1 18371
0 18373 7 14 2 44323 53701
0 18374 7 1 2 53526 54523
0 18375 7 1 2 67160 18374
0 18376 5 1 1 18375
0 18377 7 1 2 56120 61267
0 18378 7 1 2 61739 18377
0 18379 7 3 2 46497 58078
0 18380 7 1 2 67174 66768
0 18381 7 1 2 18378 18380
0 18382 5 1 1 18381
0 18383 7 1 2 18376 18382
0 18384 5 1 1 18383
0 18385 7 1 2 44217 18384
0 18386 5 1 1 18385
0 18387 7 1 2 18372 18386
0 18388 5 1 1 18387
0 18389 7 1 2 66321 18388
0 18390 5 1 1 18389
0 18391 7 4 2 44324 66053
0 18392 7 9 2 42291 42380
0 18393 7 1 2 43915 67181
0 18394 7 1 2 54524 18393
0 18395 7 1 2 67177 18394
0 18396 7 1 2 56279 59035
0 18397 7 1 2 18395 18396
0 18398 5 1 1 18397
0 18399 7 1 2 18390 18398
0 18400 5 1 1 18399
0 18401 7 1 2 67147 18400
0 18402 5 1 1 18401
0 18403 7 1 2 43090 65299
0 18404 5 1 1 18403
0 18405 7 1 2 42815 64375
0 18406 5 1 1 18405
0 18407 7 1 2 18404 18406
0 18408 5 5 1 18407
0 18409 7 1 2 55615 67190
0 18410 5 1 1 18409
0 18411 7 4 2 42816 55900
0 18412 5 1 1 67195
0 18413 7 1 2 51729 67196
0 18414 5 1 1 18413
0 18415 7 1 2 18410 18414
0 18416 5 1 1 18415
0 18417 7 1 2 53306 18416
0 18418 5 1 1 18417
0 18419 7 2 2 56523 60676
0 18420 7 1 2 58815 67199
0 18421 5 1 1 18420
0 18422 7 1 2 18418 18421
0 18423 5 1 1 18422
0 18424 7 1 2 45577 18423
0 18425 5 1 1 18424
0 18426 7 3 2 53307 55459
0 18427 7 1 2 42021 67201
0 18428 7 1 2 58816 18427
0 18429 5 1 1 18428
0 18430 7 1 2 47656 18429
0 18431 7 1 2 18425 18430
0 18432 5 1 1 18431
0 18433 7 3 2 42022 49985
0 18434 7 4 2 52781 55901
0 18435 7 1 2 67204 67207
0 18436 5 1 1 18435
0 18437 7 1 2 44325 18436
0 18438 7 1 2 17908 18437
0 18439 5 1 1 18438
0 18440 7 3 2 45078 54075
0 18441 7 2 2 50906 67211
0 18442 5 2 1 67214
0 18443 7 9 2 48433 56092
0 18444 7 1 2 57849 67218
0 18445 5 1 1 18444
0 18446 7 2 2 67216 18445
0 18447 5 2 1 67227
0 18448 7 1 2 18439 67229
0 18449 7 1 2 18432 18448
0 18450 5 1 1 18449
0 18451 7 1 2 45079 59095
0 18452 5 1 1 18451
0 18453 7 1 2 48434 66694
0 18454 5 1 1 18453
0 18455 7 1 2 58003 59155
0 18456 7 1 2 59656 18455
0 18457 7 1 2 18454 18456
0 18458 7 1 2 18452 18457
0 18459 5 1 1 18458
0 18460 7 1 2 56271 60180
0 18461 7 1 2 56475 18460
0 18462 7 1 2 59103 18461
0 18463 5 1 1 18462
0 18464 7 1 2 18459 18463
0 18465 5 1 1 18464
0 18466 7 1 2 56280 18465
0 18467 5 1 1 18466
0 18468 7 4 2 48895 59465
0 18469 5 2 1 67231
0 18470 7 1 2 17957 67235
0 18471 5 1 1 18470
0 18472 7 1 2 50844 18471
0 18473 5 1 1 18472
0 18474 7 1 2 66864 18473
0 18475 5 1 1 18474
0 18476 7 2 2 53587 18475
0 18477 7 5 2 43916 51265
0 18478 5 1 1 67239
0 18479 7 1 2 57928 67240
0 18480 5 1 1 18479
0 18481 7 1 2 56495 18480
0 18482 5 1 1 18481
0 18483 7 1 2 67237 18482
0 18484 5 1 1 18483
0 18485 7 1 2 18467 18484
0 18486 7 1 2 18450 18485
0 18487 5 1 1 18486
0 18488 7 1 2 60329 18487
0 18489 5 1 1 18488
0 18490 7 4 2 52447 61162
0 18491 7 1 2 59036 59912
0 18492 5 3 1 18491
0 18493 7 1 2 55324 58423
0 18494 7 1 2 66859 18493
0 18495 5 1 1 18494
0 18496 7 1 2 67248 18495
0 18497 5 1 1 18496
0 18498 7 1 2 67244 18497
0 18499 5 1 1 18498
0 18500 7 1 2 58193 59948
0 18501 7 1 2 65069 18500
0 18502 7 1 2 54640 18501
0 18503 5 1 1 18502
0 18504 7 1 2 18499 18503
0 18505 5 1 1 18504
0 18506 7 1 2 47286 18505
0 18507 5 1 1 18506
0 18508 7 1 2 3870 58543
0 18509 5 1 1 18508
0 18510 7 1 2 54622 61760
0 18511 7 1 2 18509 18510
0 18512 5 1 1 18511
0 18513 7 1 2 18507 18512
0 18514 5 1 1 18513
0 18515 7 1 2 65575 18514
0 18516 5 1 1 18515
0 18517 7 1 2 50203 62632
0 18518 5 1 1 18517
0 18519 7 4 2 47287 67245
0 18520 5 2 1 67251
0 18521 7 1 2 43091 67252
0 18522 5 1 1 18521
0 18523 7 1 2 18518 18522
0 18524 5 1 1 18523
0 18525 7 1 2 50845 18524
0 18526 5 1 1 18525
0 18527 7 3 2 54623 65076
0 18528 7 1 2 48115 67257
0 18529 5 2 1 18528
0 18530 7 1 2 54597 62798
0 18531 5 1 1 18530
0 18532 7 1 2 67260 18531
0 18533 5 1 1 18532
0 18534 7 1 2 49986 18533
0 18535 5 1 1 18534
0 18536 7 1 2 18526 18535
0 18537 5 1 1 18536
0 18538 7 3 2 54771 65538
0 18539 7 4 2 44326 62711
0 18540 7 1 2 67262 67265
0 18541 7 1 2 18537 18540
0 18542 5 1 1 18541
0 18543 7 1 2 18516 18542
0 18544 5 1 1 18543
0 18545 7 1 2 57632 18544
0 18546 5 1 1 18545
0 18547 7 1 2 67255 67261
0 18548 5 3 1 18547
0 18549 7 1 2 51778 60915
0 18550 5 1 1 18549
0 18551 7 1 2 67064 18550
0 18552 5 1 1 18551
0 18553 7 1 2 62926 18552
0 18554 5 1 1 18553
0 18555 7 1 2 57770 64009
0 18556 7 1 2 67266 18555
0 18557 5 1 1 18556
0 18558 7 1 2 18554 18557
0 18559 5 1 1 18558
0 18560 7 1 2 62503 18559
0 18561 5 1 1 18560
0 18562 7 2 2 59104 63854
0 18563 5 1 1 67272
0 18564 7 1 2 18048 18563
0 18565 5 1 1 18564
0 18566 7 1 2 54772 18565
0 18567 5 1 1 18566
0 18568 7 1 2 59601 61239
0 18569 5 1 1 18568
0 18570 7 1 2 42817 62274
0 18571 5 3 1 18570
0 18572 7 1 2 60713 61249
0 18573 7 1 2 67274 18572
0 18574 5 1 1 18573
0 18575 7 1 2 18569 18574
0 18576 5 1 1 18575
0 18577 7 1 2 43313 18576
0 18578 5 1 1 18577
0 18579 7 1 2 46689 60958
0 18580 7 1 2 60860 18579
0 18581 5 1 1 18580
0 18582 7 1 2 17599 18581
0 18583 5 1 1 18582
0 18584 7 1 2 66855 18583
0 18585 5 1 1 18584
0 18586 7 1 2 18578 18585
0 18587 7 1 2 18567 18586
0 18588 5 1 1 18587
0 18589 7 1 2 62690 18588
0 18590 5 1 1 18589
0 18591 7 2 2 51730 60491
0 18592 5 1 1 67277
0 18593 7 1 2 59105 59392
0 18594 5 1 1 18593
0 18595 7 1 2 18592 18594
0 18596 5 1 1 18595
0 18597 7 1 2 51938 18596
0 18598 5 1 1 18597
0 18599 7 1 2 62589 67062
0 18600 5 1 1 18599
0 18601 7 1 2 18598 18600
0 18602 5 1 1 18601
0 18603 7 1 2 63001 18602
0 18604 5 1 1 18603
0 18605 7 1 2 46255 66928
0 18606 5 1 1 18605
0 18607 7 1 2 62757 67071
0 18608 5 1 1 18607
0 18609 7 1 2 18606 18608
0 18610 5 1 1 18609
0 18611 7 1 2 43092 18610
0 18612 5 1 1 18611
0 18613 7 1 2 55543 65262
0 18614 5 1 1 18613
0 18615 7 1 2 51797 62780
0 18616 5 1 1 18615
0 18617 7 1 2 65272 18616
0 18618 7 1 2 18614 18617
0 18619 5 1 1 18618
0 18620 7 1 2 63940 18619
0 18621 5 1 1 18620
0 18622 7 1 2 18612 18621
0 18623 5 1 1 18622
0 18624 7 1 2 62927 18623
0 18625 5 1 1 18624
0 18626 7 1 2 61762 65525
0 18627 7 1 2 59106 18626
0 18628 5 1 1 18627
0 18629 7 1 2 18625 18628
0 18630 5 1 1 18629
0 18631 7 1 2 60453 18630
0 18632 5 1 1 18631
0 18633 7 1 2 18604 18632
0 18634 7 1 2 18590 18633
0 18635 7 1 2 18561 18634
0 18636 5 1 1 18635
0 18637 7 1 2 67269 18636
0 18638 5 1 1 18637
0 18639 7 1 2 18546 18638
0 18640 7 1 2 18489 18639
0 18641 5 1 1 18640
0 18642 7 1 2 48877 18641
0 18643 5 1 1 18642
0 18644 7 1 2 18402 18643
0 18645 7 1 2 18342 18644
0 18646 7 1 2 17829 18645
0 18647 5 1 1 18646
0 18648 7 1 2 53280 18647
0 18649 5 1 1 18648
0 18650 7 9 2 47006 47123
0 18651 5 1 1 67279
0 18652 7 4 2 60157 63069
0 18653 7 2 2 67280 67288
0 18654 7 1 2 61836 66294
0 18655 5 8 1 18654
0 18656 7 1 2 63477 64499
0 18657 7 1 2 67294 18656
0 18658 7 1 2 67292 18657
0 18659 5 1 1 18658
0 18660 7 2 2 10383 66619
0 18661 7 1 2 50775 63482
0 18662 7 1 2 67302 18661
0 18663 5 1 1 18662
0 18664 7 3 2 47007 44218
0 18665 7 1 2 63152 67304
0 18666 7 1 2 61782 18665
0 18667 5 1 1 18666
0 18668 7 1 2 18663 18667
0 18669 5 1 1 18668
0 18670 7 1 2 50458 18669
0 18671 5 1 1 18670
0 18672 7 1 2 43314 67303
0 18673 5 1 1 18672
0 18674 7 1 2 47008 51651
0 18675 5 1 1 18674
0 18676 7 3 2 43619 44219
0 18677 7 2 2 44778 67307
0 18678 5 1 1 67310
0 18679 7 1 2 18675 18678
0 18680 7 1 2 18673 18679
0 18681 5 1 1 18680
0 18682 7 1 2 43745 63941
0 18683 7 1 2 18681 18682
0 18684 5 1 1 18683
0 18685 7 1 2 18671 18684
0 18686 5 1 1 18685
0 18687 7 2 2 55757 59363
0 18688 7 1 2 64561 67312
0 18689 7 1 2 18686 18688
0 18690 5 1 1 18689
0 18691 7 1 2 18659 18690
0 18692 5 1 1 18691
0 18693 7 1 2 42381 18692
0 18694 5 1 1 18693
0 18695 7 6 2 46498 51798
0 18696 5 1 1 67314
0 18697 7 1 2 54535 67315
0 18698 5 2 1 18697
0 18699 7 5 2 43093 50459
0 18700 7 1 2 65300 67322
0 18701 5 1 1 18700
0 18702 7 1 2 67320 18701
0 18703 5 1 1 18702
0 18704 7 2 2 55902 67116
0 18705 7 1 2 61556 66392
0 18706 7 1 2 67327 18705
0 18707 7 1 2 18703 18706
0 18708 5 1 1 18707
0 18709 7 1 2 18694 18708
0 18710 5 1 1 18709
0 18711 7 1 2 48234 18710
0 18712 5 1 1 18711
0 18713 7 1 2 43315 65227
0 18714 5 2 1 18713
0 18715 7 2 2 42818 67316
0 18716 7 1 2 51175 67331
0 18717 5 1 1 18716
0 18718 7 1 2 67329 18717
0 18719 5 1 1 18718
0 18720 7 2 2 44905 61557
0 18721 7 2 2 62504 67088
0 18722 7 1 2 67333 67335
0 18723 7 1 2 18719 18722
0 18724 5 1 1 18723
0 18725 7 1 2 18712 18724
0 18726 5 1 1 18725
0 18727 7 1 2 42182 18726
0 18728 5 1 1 18727
0 18729 7 3 2 51142 66054
0 18730 7 1 2 46922 67337
0 18731 5 1 1 18730
0 18732 7 2 2 50415 66131
0 18733 7 1 2 43535 67340
0 18734 5 1 1 18733
0 18735 7 1 2 18731 18734
0 18736 5 13 1 18735
0 18737 7 2 2 48235 58194
0 18738 7 1 2 56484 61592
0 18739 7 1 2 66033 18738
0 18740 7 1 2 67355 18739
0 18741 7 1 2 67295 18740
0 18742 7 1 2 67342 18741
0 18743 5 1 1 18742
0 18744 7 1 2 44576 18743
0 18745 7 1 2 18728 18744
0 18746 5 1 1 18745
0 18747 7 6 2 42382 44779
0 18748 5 3 1 67357
0 18749 7 6 2 55758 66055
0 18750 7 2 2 60145 67366
0 18751 5 1 1 67372
0 18752 7 1 2 59704 67373
0 18753 5 1 1 18752
0 18754 7 1 2 51340 54052
0 18755 7 1 2 60929 18754
0 18756 7 6 2 46974 67281
0 18757 7 1 2 64660 67374
0 18758 7 1 2 18755 18757
0 18759 5 1 1 18758
0 18760 7 1 2 18753 18759
0 18761 5 1 1 18760
0 18762 7 1 2 67358 18761
0 18763 5 1 1 18762
0 18764 7 4 2 62046 66646
0 18765 7 1 2 61716 66132
0 18766 7 1 2 67380 18765
0 18767 5 1 1 18766
0 18768 7 1 2 18751 18767
0 18769 5 1 1 18768
0 18770 7 9 2 45895 48116
0 18771 5 1 1 67384
0 18772 7 2 2 46499 67385
0 18773 5 1 1 67393
0 18774 7 1 2 55652 67394
0 18775 7 1 2 18769 18774
0 18776 5 1 1 18775
0 18777 7 1 2 18763 18776
0 18778 5 1 1 18777
0 18779 7 1 2 45737 18778
0 18780 5 1 1 18779
0 18781 7 2 2 45896 56018
0 18782 5 1 1 67395
0 18783 7 1 2 67363 18782
0 18784 5 3 1 18783
0 18785 7 1 2 44327 57286
0 18786 7 1 2 59963 64750
0 18787 7 1 2 18785 18786
0 18788 7 1 2 67397 18787
0 18789 7 1 2 67343 18788
0 18790 5 1 1 18789
0 18791 7 1 2 18780 18790
0 18792 5 1 1 18791
0 18793 7 1 2 45578 18792
0 18794 5 1 1 18793
0 18795 7 1 2 42183 67344
0 18796 5 1 1 18795
0 18797 7 7 2 43620 43746
0 18798 5 1 1 67400
0 18799 7 1 2 43587 67401
0 18800 7 1 2 52555 18799
0 18801 5 1 1 18800
0 18802 7 1 2 18796 18801
0 18803 5 6 1 18802
0 18804 7 2 2 46838 67407
0 18805 5 1 1 67413
0 18806 7 7 2 47009 63070
0 18807 7 2 2 60792 67415
0 18808 7 2 2 54417 67422
0 18809 5 1 1 67424
0 18810 7 1 2 18805 18809
0 18811 5 3 1 18810
0 18812 7 2 2 59364 67426
0 18813 7 1 2 49917 57287
0 18814 7 1 2 67398 18813
0 18815 7 1 2 67429 18814
0 18816 5 1 1 18815
0 18817 7 1 2 18794 18816
0 18818 5 1 1 18817
0 18819 7 1 2 47771 18818
0 18820 5 1 1 18819
0 18821 7 2 2 67364 18771
0 18822 5 4 1 67431
0 18823 7 1 2 66745 17978
0 18824 7 2 2 67432 18823
0 18825 7 1 2 42184 67437
0 18826 5 1 1 18825
0 18827 7 2 2 42383 43536
0 18828 7 3 2 45738 67439
0 18829 7 1 2 66604 67441
0 18830 5 1 1 18829
0 18831 7 1 2 18826 18830
0 18832 5 3 1 18831
0 18833 7 6 2 44906 51176
0 18834 7 2 2 43621 67447
0 18835 5 1 1 67453
0 18836 7 3 2 47010 48236
0 18837 7 1 2 43747 67455
0 18838 5 1 1 18837
0 18839 7 1 2 18835 18838
0 18840 5 2 1 18839
0 18841 7 3 2 63685 67458
0 18842 7 5 2 59365 60517
0 18843 7 1 2 61303 67463
0 18844 7 1 2 67460 18843
0 18845 7 1 2 67444 18844
0 18846 5 1 1 18845
0 18847 7 1 2 47895 18846
0 18848 7 1 2 18820 18847
0 18849 5 1 1 18848
0 18850 7 1 2 44651 18849
0 18851 7 1 2 18746 18850
0 18852 5 1 1 18851
0 18853 7 2 2 44780 65875
0 18854 5 1 1 67468
0 18855 7 5 2 42384 46975
0 18856 7 1 2 48117 67470
0 18857 5 1 1 18856
0 18858 7 1 2 18854 18857
0 18859 5 5 1 18858
0 18860 7 5 2 43622 47124
0 18861 5 1 1 67480
0 18862 7 2 2 44907 67481
0 18863 5 1 1 67485
0 18864 7 1 2 67475 67486
0 18865 5 1 1 18864
0 18866 7 2 2 44781 55262
0 18867 5 1 1 67487
0 18868 7 1 2 65879 67488
0 18869 5 1 1 18868
0 18870 7 1 2 18865 18869
0 18871 5 1 1 18870
0 18872 7 1 2 65301 18871
0 18873 5 1 1 18872
0 18874 7 1 2 47011 55140
0 18875 7 2 2 56019 18874
0 18876 7 1 2 55379 67489
0 18877 5 1 1 18876
0 18878 7 1 2 56262 57350
0 18879 7 1 2 67311 18878
0 18880 5 1 1 18879
0 18881 7 1 2 18877 18880
0 18882 5 1 1 18881
0 18883 7 1 2 48237 67471
0 18884 7 1 2 18882 18883
0 18885 5 1 1 18884
0 18886 7 1 2 18873 18885
0 18887 5 1 1 18886
0 18888 7 1 2 43094 18887
0 18889 5 1 1 18888
0 18890 7 1 2 67448 67476
0 18891 5 1 1 18890
0 18892 7 1 2 56439 67472
0 18893 5 1 1 18892
0 18894 7 1 2 18891 18893
0 18895 5 1 1 18894
0 18896 7 1 2 43623 18895
0 18897 5 1 1 18896
0 18898 7 1 2 56440 66243
0 18899 5 1 1 18898
0 18900 7 1 2 18897 18899
0 18901 5 1 1 18900
0 18902 7 1 2 67332 18901
0 18903 5 1 1 18902
0 18904 7 1 2 18889 18903
0 18905 5 1 1 18904
0 18906 7 1 2 51588 18905
0 18907 5 1 1 18906
0 18908 7 1 2 52135 66260
0 18909 5 1 1 18908
0 18910 7 1 2 65876 67454
0 18911 5 1 1 18910
0 18912 7 1 2 18909 18911
0 18913 5 1 1 18912
0 18914 7 7 2 56956 63686
0 18915 7 2 2 44782 67491
0 18916 7 2 2 18913 67498
0 18917 7 1 2 56121 67500
0 18918 5 1 1 18917
0 18919 7 1 2 18907 18918
0 18920 5 1 1 18919
0 18921 7 1 2 42185 18920
0 18922 5 1 1 18921
0 18923 7 1 2 45739 56524
0 18924 7 1 2 67501 18923
0 18925 5 1 1 18924
0 18926 7 1 2 18922 18925
0 18927 5 1 1 18926
0 18928 7 1 2 48921 59676
0 18929 7 1 2 18927 18928
0 18930 5 1 1 18929
0 18931 7 1 2 18852 18930
0 18932 5 1 1 18931
0 18933 7 1 2 42292 18932
0 18934 5 1 1 18933
0 18935 7 3 2 43462 66056
0 18936 7 4 2 59518 67502
0 18937 7 2 2 43095 61680
0 18938 5 1 1 67509
0 18939 7 1 2 50460 67510
0 18940 5 1 1 18939
0 18941 7 1 2 67321 18940
0 18942 5 1 1 18941
0 18943 7 1 2 67505 18942
0 18944 5 1 1 18943
0 18945 7 3 2 47657 67293
0 18946 7 1 2 66697 67511
0 18947 5 1 1 18946
0 18948 7 1 2 18944 18947
0 18949 5 1 1 18948
0 18950 7 1 2 44783 18949
0 18951 5 1 1 18950
0 18952 7 1 2 47012 54217
0 18953 7 1 2 60100 18952
0 18954 7 1 2 57427 62719
0 18955 7 1 2 18953 18954
0 18956 5 1 1 18955
0 18957 7 1 2 18951 18956
0 18958 5 1 1 18957
0 18959 7 1 2 48238 18958
0 18960 5 1 1 18959
0 18961 7 1 2 51177 67317
0 18962 5 1 1 18961
0 18963 7 1 2 50158 64627
0 18964 5 1 1 18963
0 18965 7 1 2 18962 18964
0 18966 5 2 1 18965
0 18967 7 1 2 42819 67514
0 18968 5 1 1 18967
0 18969 7 1 2 67330 18968
0 18970 5 1 1 18969
0 18971 7 1 2 67367 67334
0 18972 7 1 2 18970 18971
0 18973 5 1 1 18972
0 18974 7 1 2 18960 18973
0 18975 5 1 1 18974
0 18976 7 1 2 42186 18975
0 18977 5 1 1 18976
0 18978 7 3 2 48239 66698
0 18979 7 1 2 58114 64500
0 18980 7 1 2 67345 18979
0 18981 7 1 2 67516 18980
0 18982 5 1 1 18981
0 18983 7 1 2 18977 18982
0 18984 5 1 1 18983
0 18985 7 1 2 44577 18984
0 18986 5 1 1 18985
0 18987 7 2 2 42820 53588
0 18988 7 5 2 43624 44328
0 18989 7 2 2 64507 67521
0 18990 7 1 2 60147 67526
0 18991 7 1 2 67519 18990
0 18992 7 1 2 67499 18991
0 18993 5 1 1 18992
0 18994 7 1 2 18986 18993
0 18995 5 1 1 18994
0 18996 7 1 2 47990 18995
0 18997 5 1 1 18996
0 18998 7 2 2 46976 44329
0 18999 7 1 2 42821 67528
0 19000 7 1 2 59123 18999
0 19001 7 1 2 64268 19000
0 19002 7 1 2 67461 19001
0 19003 5 1 1 19002
0 19004 7 1 2 18997 19003
0 19005 5 1 1 19004
0 19006 7 1 2 42385 19005
0 19007 5 1 1 19006
0 19008 7 4 2 59519 60518
0 19009 7 1 2 56957 67530
0 19010 7 5 2 46977 47991
0 19011 5 1 1 67534
0 19012 7 5 2 43588 44652
0 19013 5 4 1 67539
0 19014 7 1 2 19011 67544
0 19015 5 10 1 19014
0 19016 7 9 2 42187 45897
0 19017 7 3 2 44784 67558
0 19018 7 1 2 67548 67567
0 19019 7 1 2 19009 19018
0 19020 7 1 2 67462 19019
0 19021 5 1 1 19020
0 19022 7 1 2 19007 19021
0 19023 5 1 1 19022
0 19024 7 1 2 42023 19023
0 19025 5 1 1 19024
0 19026 7 1 2 53645 67341
0 19027 5 1 1 19026
0 19028 7 2 2 51143 67117
0 19029 7 1 2 46839 67570
0 19030 5 1 1 19029
0 19031 7 1 2 19027 19030
0 19032 5 5 1 19031
0 19033 7 1 2 42188 67572
0 19034 5 1 1 19033
0 19035 7 1 2 58998 67346
0 19036 5 1 1 19035
0 19037 7 1 2 19034 19036
0 19038 5 1 1 19037
0 19039 7 2 2 44785 66699
0 19040 7 3 2 42386 47992
0 19041 7 1 2 58736 59569
0 19042 7 1 2 67579 19041
0 19043 7 1 2 67577 19042
0 19044 7 1 2 19038 19043
0 19045 5 1 1 19044
0 19046 7 1 2 19025 19045
0 19047 5 1 1 19046
0 19048 7 1 2 66801 19047
0 19049 5 1 1 19048
0 19050 7 1 2 18934 19049
0 19051 5 1 1 19050
0 19052 7 1 2 54280 19051
0 19053 5 1 1 19052
0 19054 7 2 2 48240 60641
0 19055 7 4 2 42387 60401
0 19056 5 3 1 67584
0 19057 7 9 2 45898 61163
0 19058 5 1 1 67591
0 19059 7 1 2 67588 19058
0 19060 5 11 1 19059
0 19061 7 1 2 65241 67600
0 19062 5 1 1 19061
0 19063 7 1 2 52580 55315
0 19064 7 1 2 67585 19063
0 19065 5 1 1 19064
0 19066 7 1 2 19062 19065
0 19067 5 1 1 19066
0 19068 7 1 2 46690 19067
0 19069 5 1 1 19068
0 19070 7 2 2 62280 65176
0 19071 7 4 2 42388 44653
0 19072 7 1 2 62199 67613
0 19073 7 1 2 67611 19072
0 19074 5 1 1 19073
0 19075 7 1 2 19069 19074
0 19076 5 1 1 19075
0 19077 7 1 2 54773 65528
0 19078 5 1 1 19077
0 19079 7 1 2 58999 63071
0 19080 7 1 2 64680 19079
0 19081 5 1 1 19080
0 19082 7 1 2 19078 19081
0 19083 5 1 1 19082
0 19084 7 1 2 19076 19083
0 19085 5 1 1 19084
0 19086 7 5 2 45899 43537
0 19087 7 2 2 50509 67617
0 19088 5 1 1 67622
0 19089 7 2 2 42389 66438
0 19090 7 1 2 56020 67624
0 19091 5 1 1 19090
0 19092 7 1 2 19088 19091
0 19093 5 1 1 19092
0 19094 7 1 2 42189 19093
0 19095 5 1 1 19094
0 19096 7 1 2 56025 67442
0 19097 5 1 1 19096
0 19098 7 1 2 19095 19097
0 19099 5 1 1 19098
0 19100 7 1 2 54774 19099
0 19101 5 1 1 19100
0 19102 7 2 2 42024 66152
0 19103 7 1 2 50510 53646
0 19104 7 1 2 67626 19103
0 19105 5 1 1 19104
0 19106 7 1 2 19101 19105
0 19107 5 1 1 19106
0 19108 7 2 2 50268 54281
0 19109 7 1 2 60330 67628
0 19110 7 1 2 19107 19109
0 19111 5 1 1 19110
0 19112 7 1 2 19085 19111
0 19113 5 1 1 19112
0 19114 7 1 2 47896 19113
0 19115 5 1 1 19114
0 19116 7 1 2 42293 67477
0 19117 5 1 1 19116
0 19118 7 1 2 66728 66605
0 19119 5 1 1 19118
0 19120 7 1 2 19117 19119
0 19121 5 1 1 19120
0 19122 7 1 2 53702 19121
0 19123 5 1 1 19122
0 19124 7 3 2 43463 64681
0 19125 7 1 2 45900 64316
0 19126 7 1 2 53589 19125
0 19127 7 1 2 67630 19126
0 19128 5 1 1 19127
0 19129 7 1 2 19123 19128
0 19130 5 1 1 19129
0 19131 7 1 2 48934 67629
0 19132 7 1 2 19130 19131
0 19133 5 1 1 19132
0 19134 7 1 2 19115 19133
0 19135 5 1 1 19134
0 19136 7 1 2 67582 19135
0 19137 5 1 1 19136
0 19138 7 1 2 54053 54320
0 19139 5 1 1 19138
0 19140 7 1 2 57298 19139
0 19141 5 1 1 19140
0 19142 7 2 2 43096 19141
0 19143 5 1 1 67633
0 19144 7 3 2 48118 67580
0 19145 7 2 2 44578 67635
0 19146 5 1 1 67638
0 19147 7 1 2 58291 66659
0 19148 5 1 1 19147
0 19149 7 1 2 19146 19148
0 19150 5 2 1 19149
0 19151 7 1 2 67634 67640
0 19152 5 1 1 19151
0 19153 7 2 2 53803 64376
0 19154 5 1 1 67642
0 19155 7 1 2 67639 67643
0 19156 5 1 1 19155
0 19157 7 1 2 19152 19156
0 19158 5 1 1 19157
0 19159 7 1 2 55616 19158
0 19160 5 1 1 19159
0 19161 7 2 2 48241 51232
0 19162 7 2 2 65519 67644
0 19163 7 1 2 50907 66369
0 19164 7 1 2 67646 19163
0 19165 5 1 1 19164
0 19166 7 1 2 19160 19165
0 19167 5 1 1 19166
0 19168 7 1 2 46923 19167
0 19169 5 1 1 19168
0 19170 7 4 2 64522 67517
0 19171 7 1 2 45901 54423
0 19172 7 1 2 55759 19171
0 19173 7 1 2 67648 19172
0 19174 5 1 1 19173
0 19175 7 1 2 19169 19174
0 19176 5 1 1 19175
0 19177 7 1 2 45740 19176
0 19178 5 1 1 19177
0 19179 7 1 2 50087 66677
0 19180 5 1 1 19179
0 19181 7 2 2 50776 57514
0 19182 5 1 1 67652
0 19183 7 1 2 19180 19182
0 19184 5 1 1 19183
0 19185 7 1 2 46256 19184
0 19186 5 1 1 19185
0 19187 7 1 2 57422 66692
0 19188 5 1 1 19187
0 19189 7 1 2 19186 19188
0 19190 5 1 1 19189
0 19191 7 2 2 48242 19190
0 19192 7 1 2 64523 67568
0 19193 7 1 2 67654 19192
0 19194 5 1 1 19193
0 19195 7 1 2 19178 19194
0 19196 5 1 1 19195
0 19197 7 1 2 60331 19196
0 19198 5 1 1 19197
0 19199 7 1 2 51939 67601
0 19200 7 1 2 62309 19199
0 19201 5 1 1 19200
0 19202 7 1 2 61666 67559
0 19203 7 1 2 66665 19202
0 19204 5 1 1 19203
0 19205 7 1 2 19201 19204
0 19206 5 1 1 19205
0 19207 7 1 2 53804 19206
0 19208 5 1 1 19207
0 19209 7 1 2 54054 61774
0 19210 7 2 2 44220 48935
0 19211 7 1 2 67569 67656
0 19212 7 1 2 19209 19211
0 19213 5 1 1 19212
0 19214 7 1 2 19208 19213
0 19215 5 1 1 19214
0 19216 7 1 2 47772 63009
0 19217 7 1 2 19215 19216
0 19218 5 1 1 19217
0 19219 7 2 2 51779 60402
0 19220 7 1 2 66045 67658
0 19221 5 1 1 19220
0 19222 7 1 2 59290 66700
0 19223 7 1 2 67602 19222
0 19224 5 1 1 19223
0 19225 7 1 2 19221 19224
0 19226 5 1 1 19225
0 19227 7 2 2 57734 19226
0 19228 7 1 2 63002 67660
0 19229 5 1 1 19228
0 19230 7 1 2 19218 19229
0 19231 7 1 2 19198 19230
0 19232 5 1 1 19231
0 19233 7 1 2 54282 19232
0 19234 5 1 1 19233
0 19235 7 3 2 42390 44451
0 19236 7 1 2 56571 67662
0 19237 5 1 1 19236
0 19238 7 1 2 54515 66683
0 19239 5 1 1 19238
0 19240 7 1 2 19237 19239
0 19241 5 1 1 19240
0 19242 7 1 2 53590 60332
0 19243 7 2 2 19241 19242
0 19244 5 1 1 67665
0 19245 7 3 2 47897 63991
0 19246 7 1 2 64577 67592
0 19247 7 1 2 67667 19246
0 19248 5 1 1 19247
0 19249 7 1 2 19244 19248
0 19250 5 1 1 19249
0 19251 7 1 2 54913 19250
0 19252 5 1 1 19251
0 19253 7 3 2 54433 57633
0 19254 7 1 2 63211 66643
0 19255 7 1 2 67670 19254
0 19256 5 1 1 19255
0 19257 7 1 2 51858 53805
0 19258 7 1 2 57951 19257
0 19259 7 1 2 67593 19258
0 19260 5 1 1 19259
0 19261 7 1 2 19256 19260
0 19262 5 1 1 19261
0 19263 7 1 2 62691 19262
0 19264 5 1 1 19263
0 19265 7 1 2 42822 63072
0 19266 7 2 2 67671 19265
0 19267 7 1 2 42391 63212
0 19268 7 1 2 63730 19267
0 19269 7 1 2 67673 19268
0 19270 5 1 1 19269
0 19271 7 1 2 19264 19270
0 19272 7 1 2 19252 19271
0 19273 5 1 1 19272
0 19274 7 1 2 66304 19273
0 19275 5 1 1 19274
0 19276 7 4 2 42392 47288
0 19277 7 1 2 58690 67675
0 19278 7 4 2 46257 53359
0 19279 7 3 2 48243 60403
0 19280 7 1 2 67679 67683
0 19281 7 1 2 19277 19280
0 19282 5 1 1 19281
0 19283 7 2 2 57911 67560
0 19284 7 2 2 44786 67686
0 19285 7 1 2 56390 64740
0 19286 7 1 2 67688 19285
0 19287 5 1 1 19286
0 19288 7 1 2 19282 19287
0 19289 5 1 1 19288
0 19290 7 1 2 49088 19289
0 19291 5 1 1 19290
0 19292 7 1 2 48810 56093
0 19293 7 1 2 59224 19292
0 19294 7 1 2 65307 66046
0 19295 7 1 2 19293 19294
0 19296 5 1 1 19295
0 19297 7 1 2 57393 56958
0 19298 7 1 2 58897 19297
0 19299 7 1 2 67689 19298
0 19300 5 1 1 19299
0 19301 7 1 2 19296 19300
0 19302 7 1 2 19291 19301
0 19303 5 1 1 19302
0 19304 7 1 2 62692 19303
0 19305 5 1 1 19304
0 19306 7 1 2 62200 62656
0 19307 7 1 2 67473 19306
0 19308 7 2 2 56916 66478
0 19309 7 1 2 58737 60404
0 19310 7 1 2 67690 19309
0 19311 7 1 2 19307 19310
0 19312 5 1 1 19311
0 19313 7 9 2 43589 47993
0 19314 5 3 1 67692
0 19315 7 1 2 50378 67693
0 19316 7 1 2 58697 19315
0 19317 7 1 2 64741 66452
0 19318 7 1 2 19316 19317
0 19319 5 1 1 19318
0 19320 7 1 2 19312 19319
0 19321 5 1 1 19320
0 19322 7 1 2 49089 19321
0 19323 5 1 1 19322
0 19324 7 1 2 51885 57394
0 19325 7 10 2 42823 44787
0 19326 7 1 2 63383 67704
0 19327 7 1 2 19324 19326
0 19328 7 2 2 47555 56425
0 19329 7 1 2 66453 67714
0 19330 7 1 2 19327 19329
0 19331 5 1 1 19330
0 19332 7 1 2 50204 52044
0 19333 7 1 2 63073 63731
0 19334 7 1 2 19332 19333
0 19335 7 1 2 62642 66078
0 19336 7 1 2 19334 19335
0 19337 5 1 1 19336
0 19338 7 1 2 19331 19337
0 19339 7 1 2 19323 19338
0 19340 7 1 2 19305 19339
0 19341 7 1 2 19275 19340
0 19342 5 1 1 19341
0 19343 7 1 2 48435 19342
0 19344 5 1 1 19343
0 19345 7 4 2 45080 52157
0 19346 7 1 2 44654 65638
0 19347 7 1 2 67716 19346
0 19348 7 2 2 59089 19347
0 19349 7 1 2 54965 66153
0 19350 7 1 2 67720 19349
0 19351 5 1 1 19350
0 19352 7 4 2 44908 51978
0 19353 5 2 1 67722
0 19354 7 1 2 45452 54914
0 19355 5 1 1 19354
0 19356 7 1 2 67726 19355
0 19357 5 1 1 19356
0 19358 7 1 2 50088 19357
0 19359 5 1 1 19358
0 19360 7 2 2 57288 58318
0 19361 5 1 1 67728
0 19362 7 2 2 43097 58306
0 19363 7 1 2 44221 51635
0 19364 7 1 2 67730 19363
0 19365 5 1 1 19364
0 19366 7 1 2 19361 19365
0 19367 7 1 2 19359 19366
0 19368 5 1 1 19367
0 19369 7 2 2 52119 19368
0 19370 7 1 2 59325 67581
0 19371 7 1 2 67732 19370
0 19372 5 1 1 19371
0 19373 7 1 2 19351 19372
0 19374 5 1 1 19373
0 19375 7 1 2 60333 19374
0 19376 5 1 1 19375
0 19377 7 1 2 54997 66305
0 19378 7 1 2 67666 19377
0 19379 5 1 1 19378
0 19380 7 1 2 19376 19379
0 19381 7 1 2 19344 19380
0 19382 5 1 1 19381
0 19383 7 1 2 46840 19382
0 19384 5 1 1 19383
0 19385 7 1 2 47289 52158
0 19386 7 1 2 55432 56426
0 19387 7 2 2 19385 19386
0 19388 7 2 2 63074 64442
0 19389 7 2 2 45741 66332
0 19390 7 1 2 67736 67738
0 19391 7 1 2 67734 19390
0 19392 7 1 2 66306 19391
0 19393 5 1 1 19392
0 19394 7 1 2 19384 19393
0 19395 7 1 2 19234 19394
0 19396 5 1 1 19395
0 19397 7 1 2 45579 19396
0 19398 5 1 1 19397
0 19399 7 2 2 44579 60334
0 19400 7 2 2 49987 51869
0 19401 7 6 2 45902 43098
0 19402 7 1 2 64978 67744
0 19403 7 1 2 67742 19402
0 19404 5 1 1 19403
0 19405 7 2 2 48119 66439
0 19406 7 1 2 53008 66034
0 19407 7 1 2 67750 19406
0 19408 5 1 1 19407
0 19409 7 1 2 19404 19408
0 19410 5 1 1 19409
0 19411 7 1 2 45742 19410
0 19412 5 1 1 19411
0 19413 7 1 2 64979 66660
0 19414 7 1 2 65253 19413
0 19415 7 1 2 58767 19414
0 19416 5 1 1 19415
0 19417 7 1 2 19412 19416
0 19418 5 1 1 19417
0 19419 7 1 2 45453 19418
0 19420 5 1 1 19419
0 19421 7 1 2 46691 66937
0 19422 7 1 2 52126 19421
0 19423 7 1 2 66536 19422
0 19424 5 1 1 19423
0 19425 7 1 2 19420 19424
0 19426 5 1 1 19425
0 19427 7 1 2 54724 19426
0 19428 5 1 1 19427
0 19429 7 1 2 65468 18023
0 19430 5 3 1 19429
0 19431 7 2 2 45743 52479
0 19432 7 1 2 63213 67625
0 19433 7 1 2 67755 19432
0 19434 7 1 2 67752 19433
0 19435 5 1 1 19434
0 19436 7 1 2 19428 19435
0 19437 5 1 1 19436
0 19438 7 1 2 67740 19437
0 19439 5 1 1 19438
0 19440 7 1 2 54828 61164
0 19441 7 1 2 66570 19440
0 19442 7 2 2 53512 19441
0 19443 7 1 2 64613 66154
0 19444 7 1 2 67757 19443
0 19445 5 1 1 19444
0 19446 7 1 2 19439 19445
0 19447 5 1 1 19446
0 19448 7 1 2 58158 19447
0 19449 5 1 1 19448
0 19450 7 1 2 58159 67603
0 19451 7 1 2 67518 19450
0 19452 5 1 1 19451
0 19453 7 1 2 19143 19154
0 19454 5 3 1 19453
0 19455 7 1 2 45580 55617
0 19456 7 1 2 67594 19455
0 19457 7 1 2 67759 19456
0 19458 5 1 1 19457
0 19459 7 1 2 19452 19458
0 19460 5 1 1 19459
0 19461 7 1 2 60567 19460
0 19462 5 1 1 19461
0 19463 7 4 2 42393 46841
0 19464 7 2 2 61025 67762
0 19465 7 1 2 65645 67766
0 19466 7 1 2 67647 19465
0 19467 5 1 1 19466
0 19468 7 1 2 19462 19467
0 19469 5 1 1 19468
0 19470 7 1 2 62693 19469
0 19471 5 1 1 19470
0 19472 7 1 2 63365 67661
0 19473 5 1 1 19472
0 19474 7 1 2 58051 66701
0 19475 5 1 1 19474
0 19476 7 1 2 51781 61635
0 19477 5 1 1 19476
0 19478 7 1 2 19475 19477
0 19479 5 1 1 19478
0 19480 7 2 2 48244 19479
0 19481 7 1 2 58217 66397
0 19482 7 1 2 66325 19481
0 19483 7 1 2 67768 19482
0 19484 5 1 1 19483
0 19485 7 1 2 19473 19484
0 19486 7 1 2 19471 19485
0 19487 5 1 1 19486
0 19488 7 1 2 54283 19487
0 19489 5 1 1 19488
0 19490 7 4 2 45903 46842
0 19491 7 2 2 57595 67770
0 19492 7 1 2 63812 67774
0 19493 7 1 2 67735 19492
0 19494 7 1 2 66307 19493
0 19495 5 1 1 19494
0 19496 7 1 2 19489 19495
0 19497 7 1 2 19449 19496
0 19498 7 1 2 19398 19497
0 19499 5 1 1 19498
0 19500 7 1 2 47658 19499
0 19501 5 1 1 19500
0 19502 7 1 2 19137 19501
0 19503 5 1 1 19502
0 19504 7 1 2 18651 18798
0 19505 7 2 2 53216 19504
0 19506 7 1 2 19503 67776
0 19507 5 1 1 19506
0 19508 7 2 2 57845 59156
0 19509 7 6 2 44909 52873
0 19510 7 1 2 51818 67780
0 19511 7 1 2 67778 19510
0 19512 5 1 1 19511
0 19513 7 3 2 48245 49422
0 19514 5 1 1 67786
0 19515 7 1 2 62657 64257
0 19516 7 1 2 67787 19515
0 19517 5 1 1 19516
0 19518 7 1 2 19512 19517
0 19519 5 1 1 19518
0 19520 7 3 2 42294 44222
0 19521 7 1 2 61409 67789
0 19522 7 1 2 19519 19521
0 19523 5 1 1 19522
0 19524 7 2 2 61593 65898
0 19525 7 2 2 55780 67792
0 19526 7 1 2 54915 67794
0 19527 7 1 2 53513 19526
0 19528 5 1 1 19527
0 19529 7 1 2 19523 19528
0 19530 5 1 1 19529
0 19531 7 1 2 67386 19530
0 19532 5 1 1 19531
0 19533 7 1 2 67676 67717
0 19534 7 1 2 67753 19533
0 19535 7 1 2 67795 19534
0 19536 5 1 1 19535
0 19537 7 1 2 19532 19536
0 19538 5 1 1 19537
0 19539 7 1 2 54775 19538
0 19540 5 1 1 19539
0 19541 7 3 2 45081 67296
0 19542 7 1 2 55523 55974
0 19543 7 1 2 67182 19542
0 19544 7 1 2 54516 19543
0 19545 5 1 1 19544
0 19546 7 1 2 63214 66479
0 19547 7 1 2 67561 19546
0 19548 7 1 2 56433 19547
0 19549 5 1 1 19548
0 19550 7 1 2 19545 19549
0 19551 5 1 1 19550
0 19552 7 1 2 67796 19551
0 19553 5 1 1 19552
0 19554 7 1 2 45904 53398
0 19555 7 1 2 67680 19554
0 19556 7 2 2 45744 66104
0 19557 7 2 2 60035 65077
0 19558 7 1 2 67799 67801
0 19559 7 1 2 19555 19558
0 19560 5 1 1 19559
0 19561 7 1 2 19553 19560
0 19562 5 1 1 19561
0 19563 7 1 2 48246 19562
0 19564 5 1 1 19563
0 19565 7 3 2 43917 44452
0 19566 7 10 2 42190 42394
0 19567 5 1 1 67806
0 19568 7 1 2 67803 67807
0 19569 7 1 2 67758 19568
0 19570 5 1 1 19569
0 19571 7 1 2 19564 19570
0 19572 5 1 1 19571
0 19573 7 1 2 59782 19572
0 19574 5 1 1 19573
0 19575 7 1 2 19540 19574
0 19576 5 1 1 19575
0 19577 7 1 2 67347 19576
0 19578 5 1 1 19577
0 19579 7 3 2 59570 67804
0 19580 7 3 2 49649 51562
0 19581 7 1 2 45825 64780
0 19582 7 1 2 67819 19581
0 19583 5 1 1 19582
0 19584 7 2 2 64837 67790
0 19585 7 1 2 59291 67781
0 19586 7 1 2 67822 19585
0 19587 5 1 1 19586
0 19588 7 1 2 19583 19587
0 19589 5 1 1 19588
0 19590 7 1 2 67816 19589
0 19591 5 1 1 19590
0 19592 7 2 2 42295 63577
0 19593 7 2 2 49650 55172
0 19594 7 1 2 49456 67826
0 19595 7 1 2 67824 19594
0 19596 5 1 1 19595
0 19597 7 1 2 19591 19596
0 19598 5 1 1 19597
0 19599 7 1 2 43316 19598
0 19600 5 1 1 19599
0 19601 7 1 2 52730 63143
0 19602 5 1 1 19601
0 19603 7 1 2 50180 66295
0 19604 5 1 1 19603
0 19605 7 1 2 45082 62869
0 19606 7 1 2 19604 19605
0 19607 5 1 1 19606
0 19608 7 1 2 19602 19607
0 19609 5 1 1 19608
0 19610 7 2 2 48247 57912
0 19611 7 1 2 59571 66480
0 19612 7 1 2 67828 19611
0 19613 7 1 2 19609 19612
0 19614 5 1 1 19613
0 19615 7 1 2 19600 19614
0 19616 5 1 1 19615
0 19617 7 1 2 67387 19616
0 19618 5 1 1 19617
0 19619 7 1 2 62870 67782
0 19620 5 1 1 19619
0 19621 7 1 2 54588 59292
0 19622 5 1 1 19621
0 19623 7 1 2 19620 19622
0 19624 5 1 1 19623
0 19625 7 1 2 50089 19624
0 19626 5 1 1 19625
0 19627 7 2 2 54328 57748
0 19628 7 1 2 67756 67830
0 19629 5 1 1 19628
0 19630 7 1 2 19626 19629
0 19631 5 1 1 19630
0 19632 7 1 2 42824 19631
0 19633 5 1 1 19632
0 19634 7 2 2 49651 58971
0 19635 7 2 2 51341 67832
0 19636 7 1 2 64265 67834
0 19637 5 1 1 19636
0 19638 7 1 2 19633 19637
0 19639 5 1 1 19638
0 19640 7 2 2 44788 19639
0 19641 7 4 2 47994 66802
0 19642 7 4 2 59572 67838
0 19643 7 1 2 42395 67842
0 19644 7 1 2 67836 19643
0 19645 5 1 1 19644
0 19646 7 1 2 19618 19645
0 19647 5 1 1 19646
0 19648 7 1 2 67573 19647
0 19649 5 1 1 19648
0 19650 7 1 2 19578 19649
0 19651 7 1 2 19507 19650
0 19652 7 1 2 51247 55113
0 19653 5 1 1 19652
0 19654 7 5 2 48120 52448
0 19655 5 1 1 67846
0 19656 7 1 2 65221 67847
0 19657 5 1 1 19656
0 19658 7 1 2 53071 56441
0 19659 5 1 1 19658
0 19660 7 1 2 19657 19659
0 19661 5 1 1 19660
0 19662 7 1 2 43918 19661
0 19663 5 1 1 19662
0 19664 7 1 2 19653 19663
0 19665 5 1 1 19664
0 19666 7 2 2 43625 19665
0 19667 7 1 2 51664 67851
0 19668 5 1 1 19667
0 19669 7 4 2 47013 43919
0 19670 7 1 2 51589 55104
0 19671 7 1 2 67853 19670
0 19672 7 1 2 56157 19671
0 19673 5 1 1 19672
0 19674 7 1 2 19668 19673
0 19675 5 1 1 19674
0 19676 7 1 2 63687 19675
0 19677 5 1 1 19676
0 19678 7 2 2 50777 57762
0 19679 7 3 2 46258 43626
0 19680 7 2 2 43748 67859
0 19681 7 1 2 54076 67862
0 19682 5 1 1 19681
0 19683 7 1 2 42557 1390
0 19684 7 2 2 47014 44910
0 19685 5 1 1 67864
0 19686 7 2 2 43627 43920
0 19687 5 2 1 67866
0 19688 7 1 2 55530 67868
0 19689 7 1 2 19685 19688
0 19690 7 1 2 19683 19689
0 19691 5 1 1 19690
0 19692 7 1 2 19682 19691
0 19693 5 1 1 19692
0 19694 7 1 2 67857 19693
0 19695 5 1 1 19694
0 19696 7 2 2 53360 54939
0 19697 7 1 2 44223 53774
0 19698 7 1 2 67456 19697
0 19699 7 1 2 67870 19698
0 19700 5 1 1 19699
0 19701 7 1 2 19695 19700
0 19702 5 1 1 19701
0 19703 7 1 2 48121 19702
0 19704 5 1 1 19703
0 19705 7 1 2 47556 66610
0 19706 7 2 2 50711 19705
0 19707 5 1 1 67872
0 19708 7 1 2 51266 60293
0 19709 7 1 2 67873 19708
0 19710 5 1 1 19709
0 19711 7 1 2 19704 19710
0 19712 5 1 1 19711
0 19713 7 1 2 51590 19712
0 19714 5 1 1 19713
0 19715 7 1 2 19677 19714
0 19716 5 1 1 19715
0 19717 7 1 2 42191 19716
0 19718 5 1 1 19717
0 19719 7 1 2 43538 66926
0 19720 7 1 2 67852 19719
0 19721 5 1 1 19720
0 19722 7 1 2 19718 19721
0 19723 5 1 1 19722
0 19724 7 1 2 43590 19723
0 19725 5 1 1 19724
0 19726 7 1 2 50379 51178
0 19727 7 1 2 51859 55524
0 19728 7 1 2 66133 67151
0 19729 7 1 2 19727 19728
0 19730 7 1 2 19726 19729
0 19731 7 1 2 63688 19730
0 19732 5 1 1 19731
0 19733 7 1 2 19725 19732
0 19734 5 1 1 19733
0 19735 7 1 2 45454 19734
0 19736 5 1 1 19735
0 19737 7 3 2 51248 53117
0 19738 7 1 2 47015 67874
0 19739 5 1 1 19738
0 19740 7 4 2 43628 47290
0 19741 7 1 2 44789 49652
0 19742 7 1 2 67877 19741
0 19743 5 1 1 19742
0 19744 7 1 2 19739 19743
0 19745 5 1 1 19744
0 19746 7 1 2 50461 19745
0 19747 5 1 1 19746
0 19748 7 1 2 66774 67482
0 19749 5 1 1 19748
0 19750 7 1 2 19747 19749
0 19751 5 1 1 19750
0 19752 7 3 2 44224 57785
0 19753 7 2 2 43317 43591
0 19754 7 1 2 58044 67884
0 19755 7 1 2 67881 19754
0 19756 7 1 2 19751 19755
0 19757 5 1 1 19756
0 19758 7 1 2 19736 19757
0 19759 5 1 1 19758
0 19760 7 1 2 59199 19759
0 19761 5 1 1 19760
0 19762 7 1 2 67512 67837
0 19763 5 1 1 19762
0 19764 7 1 2 42396 19763
0 19765 7 1 2 19761 19764
0 19766 5 1 1 19765
0 19767 7 1 2 57196 67153
0 19768 7 1 2 63692 19767
0 19769 5 1 1 19768
0 19770 7 1 2 47659 53308
0 19771 7 2 2 57221 19770
0 19772 7 1 2 60158 67886
0 19773 7 1 2 67797 19772
0 19774 5 1 1 19773
0 19775 7 1 2 19769 19774
0 19776 5 1 1 19775
0 19777 7 1 2 62864 19776
0 19778 5 1 1 19777
0 19779 7 5 2 46034 57222
0 19780 7 7 2 55802 59998
0 19781 7 1 2 56068 67893
0 19782 7 1 2 67888 19781
0 19783 7 1 2 53514 19782
0 19784 5 1 1 19783
0 19785 7 1 2 19778 19784
0 19786 5 1 1 19785
0 19787 7 1 2 66134 19786
0 19788 5 1 1 19787
0 19789 7 2 2 52874 60036
0 19790 7 2 2 67368 67900
0 19791 7 1 2 42192 53361
0 19792 7 1 2 64204 19791
0 19793 7 1 2 67902 19792
0 19794 5 1 1 19793
0 19795 7 1 2 19788 19794
0 19796 5 1 1 19795
0 19797 7 1 2 46259 19796
0 19798 5 1 1 19797
0 19799 7 1 2 60882 67871
0 19800 7 1 2 67903 19799
0 19801 5 1 1 19800
0 19802 7 1 2 19798 19801
0 19803 5 1 1 19802
0 19804 7 1 2 48248 19803
0 19805 5 1 1 19804
0 19806 7 1 2 60101 64443
0 19807 7 1 2 66248 19806
0 19808 7 1 2 51860 56250
0 19809 7 1 2 60110 19808
0 19810 7 1 2 19807 19809
0 19811 7 1 2 63693 19810
0 19812 5 1 1 19811
0 19813 7 1 2 45905 19812
0 19814 7 1 2 19805 19813
0 19815 5 1 1 19814
0 19816 7 1 2 47995 19815
0 19817 7 1 2 19766 19816
0 19818 5 1 1 19817
0 19819 7 2 2 60965 63188
0 19820 7 2 2 43629 52449
0 19821 5 1 1 67906
0 19822 7 1 2 18478 19821
0 19823 5 1 1 19822
0 19824 7 1 2 56290 67869
0 19825 7 1 2 19823 19824
0 19826 7 1 2 67904 19825
0 19827 7 2 2 44655 67478
0 19828 7 1 2 63694 67908
0 19829 7 1 2 19826 19828
0 19830 5 1 1 19829
0 19831 7 1 2 19818 19830
0 19832 5 1 1 19831
0 19833 7 1 2 64699 19832
0 19834 5 1 1 19833
0 19835 7 1 2 51819 67183
0 19836 7 1 2 67375 19835
0 19837 7 1 2 58983 19836
0 19838 5 1 1 19837
0 19839 7 2 2 58964 66333
0 19840 7 1 2 48811 67910
0 19841 7 1 2 67408 19840
0 19842 5 1 1 19841
0 19843 7 1 2 19838 19842
0 19844 5 1 1 19843
0 19845 7 1 2 50846 19844
0 19846 5 1 1 19845
0 19847 7 1 2 46924 50295
0 19848 7 1 2 65672 19847
0 19849 7 2 2 46978 58941
0 19850 7 4 2 45745 67184
0 19851 7 3 2 46035 53337
0 19852 5 1 1 67918
0 19853 7 1 2 67914 67919
0 19854 7 1 2 67912 19853
0 19855 7 1 2 19848 19854
0 19856 5 1 1 19855
0 19857 7 1 2 48871 67589
0 19858 5 1 1 19857
0 19859 7 1 2 48878 61176
0 19860 5 1 1 19859
0 19861 7 2 2 19858 19860
0 19862 7 1 2 65529 67921
0 19863 5 1 1 19862
0 19864 7 1 2 45906 52782
0 19865 7 1 2 66611 19864
0 19866 7 1 2 66326 19865
0 19867 5 1 1 19866
0 19868 7 1 2 19863 19867
0 19869 5 1 1 19868
0 19870 7 2 2 59970 63689
0 19871 5 1 1 67923
0 19872 7 1 2 65520 67924
0 19873 7 1 2 19869 19872
0 19874 5 1 1 19873
0 19875 7 1 2 19856 19874
0 19876 7 1 2 19846 19875
0 19877 5 1 1 19876
0 19878 7 1 2 47898 19877
0 19879 5 1 1 19878
0 19880 7 1 2 67515 67860
0 19881 5 1 1 19880
0 19882 7 1 2 47016 61775
0 19883 7 1 2 62149 19882
0 19884 5 1 1 19883
0 19885 7 1 2 19881 19884
0 19886 5 1 1 19885
0 19887 7 1 2 67604 19886
0 19888 5 1 1 19887
0 19889 7 1 2 66719 67308
0 19890 7 1 2 61796 19889
0 19891 5 1 1 19890
0 19892 7 1 2 19888 19891
0 19893 5 1 1 19892
0 19894 7 1 2 43592 19893
0 19895 5 1 1 19894
0 19896 7 1 2 47557 67483
0 19897 7 2 2 56026 19896
0 19898 7 2 2 57015 67474
0 19899 7 1 2 43099 67927
0 19900 7 1 2 67925 19899
0 19901 5 1 1 19900
0 19902 7 1 2 19895 19901
0 19903 5 1 1 19902
0 19904 7 1 2 42296 19903
0 19905 5 1 1 19904
0 19906 7 1 2 56214 64023
0 19907 7 1 2 66181 19906
0 19908 7 1 2 67926 19907
0 19909 5 1 1 19908
0 19910 7 1 2 19905 19909
0 19911 5 1 1 19910
0 19912 7 1 2 59326 19911
0 19913 5 1 1 19912
0 19914 7 1 2 19879 19913
0 19915 5 1 1 19914
0 19916 7 1 2 43464 19915
0 19917 5 1 1 19916
0 19918 7 2 2 58292 58942
0 19919 7 1 2 67185 67929
0 19920 7 2 2 59037 19919
0 19921 7 1 2 67414 67931
0 19922 5 1 1 19921
0 19923 7 1 2 19917 19922
0 19924 5 1 1 19923
0 19925 7 1 2 42025 19924
0 19926 5 1 1 19925
0 19927 7 1 2 54480 67932
0 19928 7 1 2 67409 19927
0 19929 5 1 1 19928
0 19930 7 1 2 19926 19929
0 19931 5 1 1 19930
0 19932 7 1 2 44330 19931
0 19933 5 1 1 19932
0 19934 7 3 2 47660 47899
0 19935 7 3 2 55846 66057
0 19936 7 3 2 43749 64098
0 19937 7 3 2 47996 50847
0 19938 7 1 2 67939 67942
0 19939 7 1 2 67936 19938
0 19940 5 1 1 19939
0 19941 7 3 2 50416 65687
0 19942 7 1 2 58346 66447
0 19943 7 1 2 67416 19942
0 19944 7 1 2 67945 19943
0 19945 5 1 1 19944
0 19946 7 1 2 19940 19945
0 19947 5 1 1 19946
0 19948 7 1 2 67388 19947
0 19949 5 1 1 19948
0 19950 7 1 2 46925 66105
0 19951 7 1 2 51799 19950
0 19952 7 1 2 65888 19951
0 19953 7 1 2 58880 19952
0 19954 5 1 1 19953
0 19955 7 1 2 19949 19954
0 19956 5 1 1 19955
0 19957 7 1 2 45746 19956
0 19958 5 1 1 19957
0 19959 7 4 2 45826 48122
0 19960 5 1 1 67948
0 19961 7 2 2 67949 67687
0 19962 7 1 2 50848 67952
0 19963 7 1 2 67348 19962
0 19964 5 1 1 19963
0 19965 7 1 2 19958 19964
0 19966 5 1 1 19965
0 19967 7 1 2 46500 19966
0 19968 5 1 1 19967
0 19969 7 1 2 66291 67911
0 19970 7 1 2 67410 19969
0 19971 5 1 1 19970
0 19972 7 1 2 19968 19971
0 19973 5 1 1 19972
0 19974 7 1 2 46843 19973
0 19975 5 1 1 19974
0 19976 7 2 2 58965 67297
0 19977 7 1 2 66334 67425
0 19978 7 1 2 67954 19977
0 19979 5 1 1 19978
0 19980 7 1 2 19975 19979
0 19981 5 1 1 19980
0 19982 7 1 2 45581 19981
0 19983 5 1 1 19982
0 19984 7 4 2 46926 47125
0 19985 7 3 2 66135 67956
0 19986 7 4 2 42026 46036
0 19987 7 1 2 58115 67963
0 19988 7 2 2 67960 19987
0 19989 5 1 1 67967
0 19990 7 1 2 66335 67968
0 19991 7 1 2 67955 19990
0 19992 5 1 1 19991
0 19993 7 1 2 19983 19992
0 19994 5 1 1 19993
0 19995 7 1 2 42825 19994
0 19996 5 1 1 19995
0 19997 7 1 2 64109 66938
0 19998 7 1 2 56381 19997
0 19999 7 5 2 44225 47773
0 20000 7 2 2 58256 67969
0 20001 7 1 2 61257 67961
0 20002 7 1 2 67974 20001
0 20003 7 1 2 19998 20002
0 20004 5 1 1 20003
0 20005 7 1 2 19996 20004
0 20006 5 1 1 20005
0 20007 7 1 2 67933 20006
0 20008 5 1 1 20007
0 20009 7 1 2 67238 67636
0 20010 5 1 1 20009
0 20011 7 1 2 59737 60495
0 20012 5 1 1 20011
0 20013 7 2 2 49988 59730
0 20014 5 1 1 67976
0 20015 7 1 2 20012 20014
0 20016 5 1 1 20015
0 20017 7 1 2 44790 66661
0 20018 7 1 2 20016 20017
0 20019 5 1 1 20018
0 20020 7 1 2 20010 20019
0 20021 5 1 1 20020
0 20022 7 1 2 47900 20021
0 20023 5 1 1 20022
0 20024 7 1 2 8817 65469
0 20025 5 4 1 20024
0 20026 7 1 2 45907 60012
0 20027 7 1 2 67978 20026
0 20028 5 1 1 20027
0 20029 7 1 2 44453 20028
0 20030 7 1 2 20023 20029
0 20031 5 1 1 20030
0 20032 7 1 2 59491 67191
0 20033 5 1 1 20032
0 20034 7 1 2 59038 59532
0 20035 5 1 1 20034
0 20036 7 1 2 20033 20035
0 20037 5 1 1 20036
0 20038 7 1 2 45582 20037
0 20039 5 1 1 20038
0 20040 7 1 2 59039 67155
0 20041 5 1 1 20040
0 20042 7 1 2 20039 20041
0 20043 5 1 1 20042
0 20044 7 1 2 67641 20043
0 20045 5 1 1 20044
0 20046 7 1 2 54470 66393
0 20047 7 1 2 51534 20046
0 20048 5 1 1 20047
0 20049 7 1 2 55011 67637
0 20050 7 1 2 59107 20049
0 20051 5 1 1 20050
0 20052 7 1 2 20048 20051
0 20053 5 1 1 20052
0 20054 7 1 2 44331 20053
0 20055 5 1 1 20054
0 20056 7 5 2 45583 45908
0 20057 7 1 2 55460 67982
0 20058 7 1 2 60010 20057
0 20059 7 1 2 66308 20058
0 20060 5 1 1 20059
0 20061 7 1 2 20055 20060
0 20062 5 1 1 20061
0 20063 7 1 2 53591 20062
0 20064 5 1 1 20063
0 20065 7 1 2 47774 20064
0 20066 7 1 2 20045 20065
0 20067 5 1 1 20066
0 20068 7 1 2 60335 20067
0 20069 7 1 2 20031 20068
0 20070 5 1 1 20069
0 20071 7 1 2 59783 67192
0 20072 5 1 1 20071
0 20073 7 1 2 67249 20072
0 20074 5 2 1 20073
0 20075 7 1 2 67595 67987
0 20076 5 1 1 20075
0 20077 7 3 2 59366 66469
0 20078 7 1 2 63434 67989
0 20079 5 1 1 20078
0 20080 7 1 2 20076 20079
0 20081 5 1 1 20080
0 20082 7 1 2 58723 20081
0 20083 5 1 1 20082
0 20084 7 1 2 67273 67596
0 20085 5 1 1 20084
0 20086 7 2 2 66815 67605
0 20087 7 1 2 60614 67992
0 20088 5 1 1 20087
0 20089 7 1 2 20085 20088
0 20090 5 1 1 20089
0 20091 7 1 2 54776 20090
0 20092 5 1 1 20091
0 20093 7 4 2 59200 67205
0 20094 5 1 1 67994
0 20095 7 1 2 67606 67995
0 20096 5 1 1 20095
0 20097 7 1 2 60405 67763
0 20098 7 1 2 63645 20097
0 20099 7 1 2 51731 20098
0 20100 5 1 1 20099
0 20101 7 1 2 20096 20100
0 20102 5 1 1 20101
0 20103 7 1 2 61052 20102
0 20104 5 1 1 20103
0 20105 7 1 2 20092 20104
0 20106 7 1 2 20083 20105
0 20107 5 1 1 20106
0 20108 7 1 2 62694 20107
0 20109 5 1 1 20108
0 20110 7 1 2 60536 67993
0 20111 5 1 1 20110
0 20112 7 2 2 61165 67745
0 20113 5 1 1 67998
0 20114 7 1 2 63153 67614
0 20115 5 1 1 20114
0 20116 7 1 2 20113 20115
0 20117 5 2 1 20116
0 20118 7 1 2 50849 68000
0 20119 5 1 1 20118
0 20120 7 2 2 48812 67597
0 20121 5 1 1 68002
0 20122 7 1 2 67590 20121
0 20123 5 1 1 20122
0 20124 7 1 2 49989 20123
0 20125 5 1 1 20124
0 20126 7 1 2 20119 20125
0 20127 5 1 1 20126
0 20128 7 1 2 59393 20127
0 20129 5 1 1 20128
0 20130 7 1 2 20111 20129
0 20131 5 1 1 20130
0 20132 7 1 2 59293 20131
0 20133 5 1 1 20132
0 20134 7 1 2 67278 67586
0 20135 5 1 1 20134
0 20136 7 1 2 61648 67598
0 20137 7 1 2 59108 20136
0 20138 5 1 1 20137
0 20139 7 1 2 20135 20138
0 20140 5 1 1 20139
0 20141 7 1 2 51940 20140
0 20142 5 1 1 20141
0 20143 7 1 2 20133 20142
0 20144 5 1 1 20143
0 20145 7 1 2 63003 20144
0 20146 5 1 1 20145
0 20147 7 1 2 62275 67599
0 20148 5 1 1 20147
0 20149 7 1 2 49221 67587
0 20150 5 1 1 20149
0 20151 7 1 2 20148 20150
0 20152 5 1 1 20151
0 20153 7 1 2 67080 20152
0 20154 5 1 1 20153
0 20155 7 1 2 62505 67607
0 20156 5 1 1 20155
0 20157 7 1 2 63960 68003
0 20158 5 1 1 20157
0 20159 7 1 2 20156 20158
0 20160 5 1 1 20159
0 20161 7 1 2 44226 20160
0 20162 5 1 1 20161
0 20163 7 3 2 47775 67983
0 20164 7 1 2 66751 66119
0 20165 7 1 2 68004 20164
0 20166 5 1 1 20165
0 20167 7 1 2 20162 20166
0 20168 5 1 1 20167
0 20169 7 1 2 51941 20168
0 20170 5 1 1 20169
0 20171 7 1 2 20154 20170
0 20172 5 1 1 20171
0 20173 7 1 2 43318 20172
0 20174 5 1 1 20173
0 20175 7 1 2 59294 68001
0 20176 5 1 1 20175
0 20177 7 1 2 64260 67999
0 20178 5 1 1 20177
0 20179 7 1 2 20176 20178
0 20180 5 1 1 20179
0 20181 7 1 2 44227 20180
0 20182 5 1 1 20181
0 20183 7 1 2 50159 66155
0 20184 7 1 2 64089 20183
0 20185 5 1 1 20184
0 20186 7 1 2 20182 20185
0 20187 5 1 1 20186
0 20188 7 1 2 60454 20187
0 20189 5 1 1 20188
0 20190 7 1 2 20174 20189
0 20191 5 1 1 20190
0 20192 7 1 2 62741 20191
0 20193 5 1 1 20192
0 20194 7 1 2 63961 65249
0 20195 5 1 1 20194
0 20196 7 1 2 43100 63546
0 20197 5 1 1 20196
0 20198 7 1 2 20195 20197
0 20199 5 1 1 20198
0 20200 7 1 2 58374 20199
0 20201 5 1 1 20200
0 20202 7 1 2 50160 62855
0 20203 7 1 2 63706 20202
0 20204 5 1 1 20203
0 20205 7 1 2 64061 20204
0 20206 5 1 1 20205
0 20207 7 1 2 42826 20206
0 20208 5 1 1 20207
0 20209 7 1 2 20201 20208
0 20210 5 1 1 20209
0 20211 7 1 2 67608 20210
0 20212 5 1 1 20211
0 20213 7 1 2 59295 67984
0 20214 7 1 2 64545 20213
0 20215 7 1 2 67193 20214
0 20216 5 1 1 20215
0 20217 7 1 2 62506 66644
0 20218 7 1 2 67659 20217
0 20219 5 1 1 20218
0 20220 7 1 2 20216 20219
0 20221 7 1 2 20212 20220
0 20222 5 1 1 20221
0 20223 7 1 2 62928 20222
0 20224 5 1 1 20223
0 20225 7 1 2 20193 20224
0 20226 7 1 2 20146 20225
0 20227 7 1 2 20109 20226
0 20228 7 1 2 20070 20227
0 20229 5 1 1 20228
0 20230 7 1 2 67777 20229
0 20231 5 1 1 20230
0 20232 7 1 2 20008 20231
0 20233 7 1 2 19933 20232
0 20234 5 1 1 20233
0 20235 7 1 2 54870 20234
0 20236 5 1 1 20235
0 20237 7 1 2 19834 20236
0 20238 7 1 2 19651 20237
0 20239 7 1 2 19053 20238
0 20240 7 2 2 48123 48879
0 20241 7 2 2 49167 57016
0 20242 7 1 2 50462 68009
0 20243 5 1 1 20242
0 20244 7 1 2 65325 20243
0 20245 5 1 1 20244
0 20246 7 1 2 68007 20245
0 20247 5 1 1 20246
0 20248 7 2 2 66612 66035
0 20249 7 1 2 50463 50778
0 20250 7 1 2 68011 20249
0 20251 5 1 1 20250
0 20252 7 1 2 20247 20251
0 20253 5 1 1 20252
0 20254 7 1 2 43101 20253
0 20255 5 1 1 20254
0 20256 7 2 2 52334 57812
0 20257 7 1 2 43750 68013
0 20258 5 1 1 20257
0 20259 7 2 2 47558 50682
0 20260 5 1 1 68015
0 20261 7 1 2 46692 68016
0 20262 5 1 1 20261
0 20263 7 1 2 20258 20262
0 20264 5 1 1 20263
0 20265 7 1 2 68012 20264
0 20266 5 1 1 20265
0 20267 7 1 2 20255 20266
0 20268 5 1 1 20267
0 20269 7 1 2 48896 67805
0 20270 7 1 2 67267 20269
0 20271 7 1 2 20268 20270
0 20272 5 1 1 20271
0 20273 7 1 2 62156 63478
0 20274 7 3 2 55678 58279
0 20275 7 2 2 56823 66136
0 20276 7 2 2 47661 67389
0 20277 7 1 2 68020 68022
0 20278 7 1 2 68017 20277
0 20279 7 1 2 20273 20278
0 20280 5 1 1 20279
0 20281 7 1 2 20272 20280
0 20282 5 1 1 20281
0 20283 7 1 2 48436 20282
0 20284 5 1 1 20283
0 20285 7 1 2 64075 64317
0 20286 7 1 2 66402 20285
0 20287 7 3 2 47017 56824
0 20288 7 1 2 64661 68024
0 20289 7 1 2 20286 20288
0 20290 7 1 2 67798 20289
0 20291 5 1 1 20290
0 20292 7 1 2 20284 20291
0 20293 5 1 1 20292
0 20294 7 1 2 44656 20293
0 20295 5 1 1 20294
0 20296 7 2 2 52316 53854
0 20297 5 1 1 68027
0 20298 7 1 2 65326 20297
0 20299 5 1 1 20298
0 20300 7 1 2 66261 20299
0 20301 5 1 1 20300
0 20302 7 1 2 52317 55105
0 20303 7 1 2 66244 20302
0 20304 5 1 1 20303
0 20305 7 1 2 20301 20304
0 20306 5 1 1 20305
0 20307 7 1 2 44791 20306
0 20308 5 1 1 20307
0 20309 7 1 2 67490 67928
0 20310 5 1 1 20309
0 20311 7 1 2 20308 20310
0 20312 5 1 1 20311
0 20313 7 1 2 43102 20312
0 20314 5 1 1 20313
0 20315 7 1 2 46260 58347
0 20316 7 1 2 66740 20315
0 20317 7 1 2 48880 57709
0 20318 7 1 2 20316 20317
0 20319 5 1 1 20318
0 20320 7 1 2 20314 20319
0 20321 5 1 1 20320
0 20322 7 1 2 43921 20321
0 20323 5 1 1 20322
0 20324 7 2 2 43319 47018
0 20325 7 1 2 51101 51386
0 20326 7 1 2 68029 20325
0 20327 5 1 1 20326
0 20328 7 1 2 19707 20327
0 20329 5 1 1 20328
0 20330 7 1 2 42397 20329
0 20331 5 1 1 20330
0 20332 7 2 2 45909 67402
0 20333 7 1 2 51387 53362
0 20334 7 1 2 68031 20333
0 20335 5 1 1 20334
0 20336 7 1 2 20331 20335
0 20337 5 1 1 20336
0 20338 7 1 2 46979 47291
0 20339 7 1 2 57004 20338
0 20340 7 1 2 20337 20339
0 20341 5 1 1 20340
0 20342 7 1 2 20323 20341
0 20343 5 1 1 20342
0 20344 7 1 2 48437 20343
0 20345 5 1 1 20344
0 20346 7 2 2 53338 67878
0 20347 7 1 2 50464 51643
0 20348 7 1 2 68033 20347
0 20349 5 1 1 20348
0 20350 7 1 2 42558 67854
0 20351 7 1 2 57428 20350
0 20352 5 1 1 20351
0 20353 7 1 2 20349 20352
0 20354 5 1 1 20353
0 20355 7 1 2 46980 57763
0 20356 7 1 2 66639 20355
0 20357 7 1 2 20354 20356
0 20358 5 1 1 20357
0 20359 7 1 2 20345 20358
0 20360 5 1 1 20359
0 20361 7 1 2 63189 64496
0 20362 7 1 2 20360 20361
0 20363 5 1 1 20362
0 20364 7 1 2 20295 20363
0 20365 5 1 1 20364
0 20366 7 1 2 44580 20365
0 20367 5 1 1 20366
0 20368 7 1 2 42398 370
0 20369 7 1 2 66743 67701
0 20370 7 1 2 20368 20369
0 20371 7 1 2 66620 20370
0 20372 5 2 1 20371
0 20373 7 1 2 61166 66245
0 20374 5 1 1 20373
0 20375 7 1 2 68035 20374
0 20376 5 2 1 20375
0 20377 7 1 2 46927 68037
0 20378 5 1 1 20377
0 20379 7 1 2 66137 67623
0 20380 5 1 1 20379
0 20381 7 1 2 20378 20380
0 20382 5 1 1 20381
0 20383 7 1 2 50720 55162
0 20384 7 1 2 65660 20383
0 20385 7 1 2 67492 20384
0 20386 7 1 2 20382 20385
0 20387 5 1 1 20386
0 20388 7 1 2 20367 20387
0 20389 5 1 1 20388
0 20390 7 1 2 42193 20389
0 20391 5 1 1 20390
0 20392 7 1 2 45910 49423
0 20393 7 1 2 66058 67970
0 20394 7 1 2 20392 20393
0 20395 7 1 2 63245 64221
0 20396 7 1 2 20394 20395
0 20397 5 1 1 20396
0 20398 7 1 2 62507 65158
0 20399 7 1 2 63695 20398
0 20400 7 1 2 68038 20399
0 20401 5 1 1 20400
0 20402 7 1 2 20397 20401
0 20403 5 1 1 20402
0 20404 7 1 2 52552 60190
0 20405 7 1 2 20403 20404
0 20406 5 1 1 20405
0 20407 7 1 2 20391 20406
0 20408 5 1 1 20407
0 20409 7 1 2 48249 20408
0 20410 5 1 1 20409
0 20411 7 2 2 52318 54574
0 20412 7 1 2 43630 68039
0 20413 5 1 1 20412
0 20414 7 1 2 47019 52298
0 20415 7 1 2 54548 20414
0 20416 5 1 1 20415
0 20417 7 1 2 20413 20416
0 20418 5 1 1 20417
0 20419 7 1 2 50465 20418
0 20420 5 1 1 20419
0 20421 7 1 2 50296 55270
0 20422 7 1 2 68034 20421
0 20423 5 1 1 20422
0 20424 7 1 2 20420 20423
0 20425 5 1 1 20424
0 20426 7 1 2 51591 20425
0 20427 5 1 1 20426
0 20428 7 1 2 55075 8844
0 20429 5 3 1 20428
0 20430 7 5 2 47559 52279
0 20431 5 1 1 68044
0 20432 7 1 2 43631 57264
0 20433 7 1 2 68045 20432
0 20434 7 1 2 68041 20433
0 20435 5 1 1 20434
0 20436 7 1 2 20427 20435
0 20437 5 1 1 20436
0 20438 7 1 2 66741 20437
0 20439 5 1 1 20438
0 20440 7 1 2 56122 64654
0 20441 7 1 2 66076 20440
0 20442 7 1 2 58298 59971
0 20443 7 1 2 20441 20442
0 20444 5 1 1 20443
0 20445 7 1 2 20439 20444
0 20446 5 1 1 20445
0 20447 7 1 2 42399 20446
0 20448 5 1 1 20447
0 20449 7 1 2 46928 56291
0 20450 5 2 1 20449
0 20451 7 1 2 50466 51592
0 20452 5 1 1 20451
0 20453 7 1 2 68049 20452
0 20454 5 1 1 20453
0 20455 7 1 2 68010 20454
0 20456 5 1 1 20455
0 20457 7 2 2 42827 59238
0 20458 7 2 2 67882 68051
0 20459 5 1 1 68053
0 20460 7 1 2 47126 68054
0 20461 5 1 1 20460
0 20462 7 1 2 20456 20461
0 20463 5 1 1 20462
0 20464 7 1 2 45083 67879
0 20465 7 1 2 67469 20464
0 20466 7 1 2 20463 20465
0 20467 5 1 1 20466
0 20468 7 1 2 20448 20467
0 20469 5 1 1 20468
0 20470 7 1 2 43103 20469
0 20471 5 1 1 20470
0 20472 7 2 2 65177 66249
0 20473 7 1 2 43922 68055
0 20474 5 1 1 20473
0 20475 7 1 2 48438 57979
0 20476 7 1 2 66236 20475
0 20477 5 1 1 20476
0 20478 7 1 2 20474 20477
0 20479 5 1 1 20478
0 20480 7 1 2 65222 20479
0 20481 5 1 1 20480
0 20482 7 1 2 55071 68056
0 20483 5 1 1 20482
0 20484 7 1 2 20481 20483
0 20485 5 1 1 20484
0 20486 7 1 2 42400 20485
0 20487 5 1 1 20486
0 20488 7 3 2 45911 43751
0 20489 7 2 2 66059 68057
0 20490 7 1 2 51833 57980
0 20491 7 1 2 68060 20490
0 20492 5 1 1 20491
0 20493 7 1 2 20487 20492
0 20494 5 2 1 20493
0 20495 7 1 2 55737 63976
0 20496 7 1 2 68062 20495
0 20497 5 1 1 20496
0 20498 7 1 2 20471 20497
0 20499 5 1 1 20498
0 20500 7 1 2 42194 20499
0 20501 5 1 1 20500
0 20502 7 1 2 52553 67493
0 20503 7 1 2 68063 20502
0 20504 5 1 1 20503
0 20505 7 1 2 20501 20504
0 20506 5 1 1 20505
0 20507 7 1 2 47997 20506
0 20508 5 1 1 20507
0 20509 7 3 2 43632 44657
0 20510 7 1 2 67445 67494
0 20511 5 1 1 20510
0 20512 7 3 2 60037 67808
0 20513 7 2 2 46501 55544
0 20514 5 1 1 68070
0 20515 7 1 2 62712 68071
0 20516 7 1 2 68067 20515
0 20517 5 1 1 20516
0 20518 7 1 2 20511 20517
0 20519 5 1 1 20518
0 20520 7 1 2 55106 20519
0 20521 5 1 1 20520
0 20522 7 1 2 51342 51593
0 20523 7 1 2 66606 20522
0 20524 7 2 2 42195 66640
0 20525 7 1 2 65225 68072
0 20526 7 1 2 20523 20525
0 20527 5 1 1 20526
0 20528 7 1 2 20521 20527
0 20529 5 1 1 20528
0 20530 7 1 2 47292 20529
0 20531 5 1 1 20530
0 20532 7 1 2 59239 62658
0 20533 7 1 2 66182 20532
0 20534 7 1 2 62141 62808
0 20535 7 1 2 20533 20534
0 20536 5 1 1 20535
0 20537 7 1 2 20531 20536
0 20538 5 1 1 20537
0 20539 7 1 2 45084 20538
0 20540 5 1 1 20539
0 20541 7 1 2 47127 50161
0 20542 7 1 2 53399 62713
0 20543 7 1 2 20541 20542
0 20544 7 1 2 68073 67901
0 20545 7 1 2 20543 20544
0 20546 5 1 1 20545
0 20547 7 1 2 20540 20546
0 20548 5 1 1 20547
0 20549 7 1 2 68064 20548
0 20550 5 1 1 20549
0 20551 7 1 2 20508 20550
0 20552 5 1 1 20551
0 20553 7 1 2 59201 20552
0 20554 5 1 1 20553
0 20555 7 2 2 67417 67562
0 20556 5 1 1 68074
0 20557 7 1 2 59593 64987
0 20558 7 3 2 58280 60930
0 20559 7 1 2 65211 68076
0 20560 7 1 2 20557 20559
0 20561 7 1 2 68075 20560
0 20562 5 1 1 20561
0 20563 7 1 2 20554 20562
0 20564 5 1 1 20563
0 20565 7 1 2 44911 62508
0 20566 7 1 2 20564 20565
0 20567 5 1 1 20566
0 20568 7 1 2 20410 20567
0 20569 5 1 1 20568
0 20570 7 1 2 42297 20569
0 20571 5 1 1 20570
0 20572 7 2 2 60106 67118
0 20573 7 3 2 42196 67186
0 20574 7 1 2 54424 65078
0 20575 7 1 2 68081 20574
0 20576 7 1 2 68079 20575
0 20577 5 1 1 20576
0 20578 7 1 2 65178 67289
0 20579 7 5 2 63798 65850
0 20580 7 2 2 61508 67934
0 20581 7 1 2 68084 68089
0 20582 7 1 2 20578 20581
0 20583 5 1 1 20582
0 20584 7 1 2 20577 20583
0 20585 5 1 1 20584
0 20586 7 1 2 45455 20585
0 20587 5 1 1 20586
0 20588 7 6 2 43539 43633
0 20589 5 1 1 68091
0 20590 7 1 2 45912 60038
0 20591 7 1 2 68092 20590
0 20592 5 1 1 20591
0 20593 7 1 2 51630 66615
0 20594 5 1 1 20593
0 20595 7 1 2 42401 1736
0 20596 7 1 2 20589 20595
0 20597 7 1 2 20594 20596
0 20598 5 1 1 20597
0 20599 7 1 2 20592 20598
0 20600 5 1 1 20599
0 20601 7 1 2 47998 20600
0 20602 5 1 1 20601
0 20603 7 3 2 47020 67618
0 20604 7 1 2 56302 68097
0 20605 5 1 1 20604
0 20606 7 1 2 20602 20605
0 20607 5 1 1 20606
0 20608 7 1 2 42197 20607
0 20609 5 1 1 20608
0 20610 7 2 2 43634 47901
0 20611 7 1 2 61167 68100
0 20612 7 1 2 67443 20611
0 20613 5 1 1 20612
0 20614 7 1 2 20609 20613
0 20615 5 1 1 20614
0 20616 7 1 2 60336 20615
0 20617 5 1 1 20616
0 20618 7 1 2 47021 47902
0 20619 7 1 2 67609 20618
0 20620 7 1 2 65530 20619
0 20621 5 1 1 20620
0 20622 7 1 2 20617 20621
0 20623 5 1 1 20622
0 20624 7 1 2 56263 20623
0 20625 5 1 1 20624
0 20626 7 1 2 65847 65877
0 20627 5 1 1 20626
0 20628 7 1 2 68036 20627
0 20629 5 1 1 20628
0 20630 7 1 2 42298 20629
0 20631 5 1 1 20630
0 20632 7 1 2 44792 66426
0 20633 5 1 1 20632
0 20634 7 1 2 20631 20633
0 20635 5 1 1 20634
0 20636 7 1 2 50672 52783
0 20637 7 1 2 20635 20636
0 20638 5 1 1 20637
0 20639 7 1 2 20625 20638
0 20640 5 1 1 20639
0 20641 7 1 2 48439 61931
0 20642 7 1 2 20640 20641
0 20643 5 1 1 20642
0 20644 7 1 2 20587 20643
0 20645 5 1 1 20644
0 20646 7 1 2 48250 20645
0 20647 5 1 1 20646
0 20648 7 2 2 55421 65531
0 20649 7 2 2 48881 57856
0 20650 7 1 2 68102 68104
0 20651 5 1 1 20650
0 20652 7 2 2 51594 67809
0 20653 7 1 2 60337 66617
0 20654 7 1 2 68106 20653
0 20655 5 1 1 20654
0 20656 7 1 2 20651 20655
0 20657 5 1 1 20656
0 20658 7 9 2 47999 44912
0 20659 7 3 2 48440 68108
0 20660 7 1 2 59202 61777
0 20661 7 1 2 68117 20660
0 20662 7 1 2 20657 20661
0 20663 5 1 1 20662
0 20664 7 1 2 20647 20663
0 20665 5 1 1 20664
0 20666 7 1 2 43923 20665
0 20667 5 1 1 20666
0 20668 7 1 2 64714 68061
0 20669 5 1 1 20668
0 20670 7 4 2 50467 55422
0 20671 7 1 2 48882 60311
0 20672 7 1 2 68120 20671
0 20673 5 1 1 20672
0 20674 7 1 2 20669 20673
0 20675 5 1 1 20674
0 20676 7 1 2 44913 20675
0 20677 5 1 1 20676
0 20678 7 1 2 48864 51179
0 20679 7 1 2 58738 60324
0 20680 7 1 2 20678 20679
0 20681 5 1 1 20680
0 20682 7 1 2 20677 20681
0 20683 5 1 1 20682
0 20684 7 1 2 48000 20683
0 20685 5 1 1 20684
0 20686 7 2 2 56264 60338
0 20687 7 2 2 47903 54434
0 20688 7 1 2 48867 68126
0 20689 7 1 2 68124 20688
0 20690 5 1 1 20689
0 20691 7 1 2 20685 20690
0 20692 5 1 1 20691
0 20693 7 1 2 44793 20692
0 20694 5 1 1 20693
0 20695 7 1 2 46981 66539
0 20696 5 1 1 20695
0 20697 7 1 2 7878 67702
0 20698 5 1 1 20697
0 20699 7 2 2 43593 47904
0 20700 5 1 1 68128
0 20701 7 1 2 45827 20700
0 20702 7 1 2 20698 20701
0 20703 5 1 1 20702
0 20704 7 1 2 20696 20703
0 20705 5 1 1 20704
0 20706 7 1 2 43752 20705
0 20707 5 1 1 20706
0 20708 7 2 2 42559 46982
0 20709 5 1 1 68130
0 20710 7 6 2 57941 66571
0 20711 5 2 1 68132
0 20712 7 1 2 68131 68133
0 20713 5 1 1 20712
0 20714 7 1 2 20707 20713
0 20715 5 1 1 20714
0 20716 7 1 2 51249 66373
0 20717 7 1 2 20715 20716
0 20718 5 1 1 20717
0 20719 7 1 2 20694 20718
0 20720 5 1 1 20719
0 20721 7 1 2 43540 20720
0 20722 5 1 1 20721
0 20723 7 1 2 50468 54055
0 20724 7 1 2 68129 20723
0 20725 7 2 2 67922 20724
0 20726 7 1 2 65619 68140
0 20727 5 1 1 20726
0 20728 7 1 2 20722 20727
0 20729 5 1 1 20728
0 20730 7 1 2 42198 20729
0 20731 5 1 1 20730
0 20732 7 3 2 43541 63992
0 20733 7 1 2 68141 68142
0 20734 5 1 1 20733
0 20735 7 1 2 20731 20734
0 20736 5 1 1 20735
0 20737 7 1 2 52581 61932
0 20738 7 1 2 20736 20737
0 20739 5 1 1 20738
0 20740 7 1 2 20667 20739
0 20741 5 1 1 20740
0 20742 7 1 2 46261 20741
0 20743 5 1 1 20742
0 20744 7 3 2 48124 67449
0 20745 5 1 1 68145
0 20746 7 5 2 42299 54500
0 20747 7 1 2 66357 68148
0 20748 7 1 2 68146 20747
0 20749 5 1 1 20748
0 20750 7 1 2 58293 66341
0 20751 5 1 1 20750
0 20752 7 1 2 68008 67741
0 20753 5 1 1 20752
0 20754 7 1 2 20751 20753
0 20755 5 1 1 20754
0 20756 7 1 2 55263 56347
0 20757 7 1 2 20755 20756
0 20758 5 1 1 20757
0 20759 7 1 2 20749 20758
0 20760 5 1 1 20759
0 20761 7 1 2 42199 20760
0 20762 5 1 1 20761
0 20763 7 1 2 53563 20762
0 20764 5 1 1 20763
0 20765 7 2 2 45828 66374
0 20766 5 1 1 68153
0 20767 7 2 2 43594 68154
0 20768 5 1 1 68155
0 20769 7 2 2 17253 20768
0 20770 5 8 1 68157
0 20771 7 2 2 48251 61168
0 20772 7 1 2 68121 68167
0 20773 7 1 2 68159 20772
0 20774 5 1 1 20773
0 20775 7 1 2 52796 20774
0 20776 5 1 1 20775
0 20777 7 1 2 52731 59203
0 20778 7 1 2 63942 20777
0 20779 7 1 2 20776 20778
0 20780 7 1 2 20764 20779
0 20781 5 1 1 20780
0 20782 7 1 2 20743 20781
0 20783 5 1 1 20782
0 20784 7 1 2 62509 20783
0 20785 5 1 1 20784
0 20786 7 15 2 67178 67084
0 20787 7 1 2 63154 64668
0 20788 7 1 2 68169 20787
0 20789 5 1 1 20788
0 20790 7 2 2 45913 63155
0 20791 5 1 1 68184
0 20792 7 1 2 67365 20791
0 20793 5 1 1 20792
0 20794 7 3 2 47022 47662
0 20795 7 1 2 61300 68186
0 20796 7 1 2 65496 20795
0 20797 7 1 2 20793 20796
0 20798 5 1 1 20797
0 20799 7 1 2 20789 20798
0 20800 5 1 1 20799
0 20801 7 1 2 45747 20800
0 20802 5 1 1 20801
0 20803 7 2 2 61036 67861
0 20804 7 1 2 67232 68189
0 20805 7 1 2 67438 20804
0 20806 5 1 1 20805
0 20807 7 1 2 20802 20806
0 20808 5 1 1 20807
0 20809 7 1 2 47905 20808
0 20810 5 1 1 20809
0 20811 7 1 2 64669 68068
0 20812 7 1 2 67506 20811
0 20813 5 1 1 20812
0 20814 7 1 2 20810 20813
0 20815 5 1 1 20814
0 20816 7 1 2 44658 20815
0 20817 5 1 1 20816
0 20818 7 1 2 46262 55781
0 20819 7 1 2 67563 20818
0 20820 7 1 2 61677 20819
0 20821 7 1 2 67507 20820
0 20822 5 1 1 20821
0 20823 7 1 2 20817 20822
0 20824 5 1 1 20823
0 20825 7 1 2 47128 20824
0 20826 5 1 1 20825
0 20827 7 2 2 56234 67369
0 20828 7 3 2 44581 61290
0 20829 7 1 2 55185 68193
0 20830 7 1 2 67610 20829
0 20831 7 1 2 68191 20830
0 20832 5 1 1 20831
0 20833 7 1 2 20826 20832
0 20834 5 1 1 20833
0 20835 7 1 2 42300 20834
0 20836 5 1 1 20835
0 20837 7 3 2 58752 59843
0 20838 5 1 1 68196
0 20839 7 2 2 50356 68197
0 20840 7 2 2 48813 67484
0 20841 7 1 2 66481 68201
0 20842 7 1 2 67479 20841
0 20843 7 1 2 68199 20842
0 20844 5 1 1 20843
0 20845 7 1 2 20836 20844
0 20846 5 1 1 20845
0 20847 7 1 2 46502 20846
0 20848 5 1 1 20847
0 20849 7 1 2 65250 67396
0 20850 5 1 1 20849
0 20851 7 1 2 49516 54425
0 20852 7 1 2 67810 20851
0 20853 5 1 1 20852
0 20854 7 1 2 20850 20853
0 20855 5 2 1 20854
0 20856 7 1 2 63809 67282
0 20857 7 2 2 63436 20856
0 20858 5 1 1 68205
0 20859 7 5 2 47663 48001
0 20860 7 1 2 66803 68207
0 20861 7 1 2 68206 20860
0 20862 7 1 2 68203 20861
0 20863 5 1 1 20862
0 20864 7 1 2 20848 20863
0 20865 5 1 1 20864
0 20866 7 1 2 54871 20865
0 20867 5 1 1 20866
0 20868 7 1 2 46983 54658
0 20869 7 1 2 59573 20868
0 20870 7 1 2 61807 62232
0 20871 7 1 2 20869 20870
0 20872 5 1 1 20871
0 20873 7 3 2 48897 60486
0 20874 7 3 2 61927 68212
0 20875 7 1 2 66607 68122
0 20876 7 1 2 68215 20875
0 20877 5 1 1 20876
0 20878 7 1 2 20872 20877
0 20879 5 1 1 20878
0 20880 7 1 2 67811 20879
0 20881 5 1 1 20880
0 20882 7 1 2 46984 54453
0 20883 7 1 2 61740 63955
0 20884 7 1 2 20882 20883
0 20885 7 3 2 45584 66156
0 20886 7 1 2 54104 68218
0 20887 7 1 2 20884 20886
0 20888 5 1 1 20887
0 20889 7 1 2 20881 20888
0 20890 5 1 1 20889
0 20891 7 1 2 46929 20890
0 20892 5 1 1 20891
0 20893 7 1 2 66608 66939
0 20894 5 1 1 20893
0 20895 7 1 2 64318 67564
0 20896 5 1 1 20895
0 20897 7 1 2 20894 20896
0 20898 5 1 1 20897
0 20899 7 1 2 68123 20898
0 20900 5 1 1 20899
0 20901 7 1 2 64508 68069
0 20902 5 1 1 20901
0 20903 7 1 2 20900 20902
0 20904 5 1 1 20903
0 20905 7 2 2 44454 61604
0 20906 7 1 2 67531 68221
0 20907 7 1 2 20904 20906
0 20908 5 1 1 20907
0 20909 7 1 2 20892 20908
0 20910 5 1 1 20909
0 20911 7 1 2 47023 20910
0 20912 5 1 1 20911
0 20913 7 1 2 42402 61801
0 20914 5 1 1 20913
0 20915 7 1 2 18773 20914
0 20916 5 1 1 20915
0 20917 7 2 2 60519 67403
0 20918 7 1 2 56235 62714
0 20919 7 1 2 68194 20918
0 20920 7 1 2 68223 20919
0 20921 7 1 2 20916 20920
0 20922 5 1 1 20921
0 20923 7 1 2 20912 20922
0 20924 5 1 1 20923
0 20925 7 1 2 48252 20924
0 20926 5 1 1 20925
0 20927 7 1 2 56391 68202
0 20928 7 1 2 68216 20927
0 20929 7 1 2 67446 20928
0 20930 5 1 1 20929
0 20931 7 1 2 44659 20930
0 20932 7 1 2 20926 20931
0 20933 5 1 1 20932
0 20934 7 2 2 66250 68107
0 20935 7 1 2 52136 68225
0 20936 5 1 1 20935
0 20937 7 1 2 59296 67619
0 20938 7 1 2 67459 20937
0 20939 5 1 1 20938
0 20940 7 1 2 44914 61253
0 20941 7 1 2 48883 20940
0 20942 7 1 2 58828 20941
0 20943 5 1 1 20942
0 20944 7 1 2 20939 20943
0 20945 5 1 1 20944
0 20946 7 1 2 43595 20945
0 20947 5 1 1 20946
0 20948 7 1 2 20936 20947
0 20949 5 1 1 20948
0 20950 7 1 2 44794 20949
0 20951 5 1 1 20950
0 20952 7 1 2 68147 68226
0 20953 5 1 1 20952
0 20954 7 1 2 20951 20953
0 20955 5 1 1 20954
0 20956 7 1 2 68217 20955
0 20957 5 1 1 20956
0 20958 7 1 2 48002 20957
0 20959 5 1 1 20958
0 20960 7 1 2 42301 20959
0 20961 7 1 2 20933 20960
0 20962 5 1 1 20961
0 20963 7 1 2 47024 55264
0 20964 5 1 1 20963
0 20965 7 1 2 18863 20964
0 20966 5 1 1 20965
0 20967 7 1 2 67909 20966
0 20968 5 1 1 20967
0 20969 7 2 2 46985 68109
0 20970 7 1 2 68105 68227
0 20971 5 1 1 20970
0 20972 7 1 2 20968 20971
0 20973 5 1 1 20972
0 20974 7 1 2 55423 20973
0 20975 5 1 1 20974
0 20976 7 1 2 56444 20745
0 20977 5 1 1 20976
0 20978 7 1 2 48936 66188
0 20979 7 1 2 20977 20978
0 20980 5 1 1 20979
0 20981 7 1 2 20975 20980
0 20982 5 1 1 20981
0 20983 7 1 2 56525 62659
0 20984 7 2 2 64682 20983
0 20985 7 1 2 44455 59204
0 20986 7 1 2 68229 20985
0 20987 7 1 2 20982 20986
0 20988 5 1 1 20987
0 20989 7 1 2 20962 20988
0 20990 5 1 1 20989
0 20991 7 1 2 54284 20990
0 20992 5 1 1 20991
0 20993 7 2 2 63664 67283
0 20994 7 1 2 53466 66036
0 20995 7 1 2 62841 20994
0 20996 7 1 2 68231 20995
0 20997 7 1 2 63438 20996
0 20998 5 1 1 20997
0 20999 7 1 2 55233 67390
0 21000 7 1 2 63190 20999
0 21001 7 1 2 67338 21000
0 21002 5 1 1 21001
0 21003 7 1 2 61094 67359
0 21004 7 1 2 67284 21003
0 21005 7 1 2 58639 63310
0 21006 7 1 2 21004 21005
0 21007 5 1 1 21006
0 21008 7 1 2 21002 21007
0 21009 5 1 1 21008
0 21010 7 1 2 45085 65688
0 21011 7 1 2 21009 21010
0 21012 5 1 1 21011
0 21013 7 1 2 20998 21012
0 21014 5 1 1 21013
0 21015 7 1 2 51942 21014
0 21016 5 1 1 21015
0 21017 7 3 2 44660 66987
0 21018 7 6 2 59297 68233
0 21019 7 1 2 61802 63311
0 21020 7 4 2 42403 46037
0 21021 7 3 2 45086 68242
0 21022 7 1 2 68232 68246
0 21023 7 1 2 21019 21022
0 21024 7 1 2 68236 21023
0 21025 5 1 1 21024
0 21026 7 1 2 21016 21025
0 21027 5 1 1 21026
0 21028 7 1 2 48253 60455
0 21029 7 1 2 21027 21028
0 21030 5 1 1 21029
0 21031 7 1 2 60615 66729
0 21032 7 1 2 62799 21031
0 21033 7 1 2 54872 21032
0 21034 5 1 1 21033
0 21035 7 1 2 56069 59669
0 21036 7 2 2 45914 65689
0 21037 7 1 2 63554 68249
0 21038 7 1 2 21035 21037
0 21039 5 1 1 21038
0 21040 7 1 2 21034 21039
0 21041 5 1 1 21040
0 21042 7 1 2 43104 54777
0 21043 7 1 2 21041 21042
0 21044 5 1 1 21043
0 21045 7 2 2 52159 63993
0 21046 7 1 2 52045 57634
0 21047 7 1 2 67615 21046
0 21048 7 1 2 68251 21047
0 21049 5 1 1 21048
0 21050 7 1 2 54829 62865
0 21051 7 1 2 67953 21050
0 21052 5 1 1 21051
0 21053 7 1 2 21049 21052
0 21054 5 1 1 21053
0 21055 7 1 2 48441 21054
0 21056 5 1 1 21055
0 21057 7 1 2 56490 67915
0 21058 5 1 1 21057
0 21059 7 3 2 42200 66336
0 21060 7 1 2 57929 68253
0 21061 5 1 1 21060
0 21062 7 1 2 21058 21061
0 21063 5 1 1 21062
0 21064 7 1 2 49653 60294
0 21065 7 1 2 21063 21064
0 21066 5 1 1 21065
0 21067 7 1 2 21056 21066
0 21068 5 1 1 21067
0 21069 7 1 2 58195 60229
0 21070 7 1 2 21068 21069
0 21071 5 1 1 21070
0 21072 7 1 2 21044 21071
0 21073 5 1 1 21072
0 21074 7 1 2 67349 21073
0 21075 5 1 1 21074
0 21076 7 1 2 54873 68204
0 21077 5 1 1 21076
0 21078 7 1 2 63215 64789
0 21079 7 1 2 66157 21078
0 21080 7 1 2 53787 21079
0 21081 5 1 1 21080
0 21082 7 1 2 21077 21081
0 21083 5 1 1 21082
0 21084 7 1 2 67843 21083
0 21085 5 1 1 21084
0 21086 7 2 2 54589 60406
0 21087 7 1 2 68256 67746
0 21088 7 1 2 67825 21087
0 21089 5 1 1 21088
0 21090 7 1 2 21085 21089
0 21091 5 1 1 21090
0 21092 7 1 2 67574 21091
0 21093 5 1 1 21092
0 21094 7 1 2 21075 21093
0 21095 7 1 2 21030 21094
0 21096 7 1 2 20992 21095
0 21097 7 1 2 20867 21096
0 21098 7 1 2 20785 21097
0 21099 5 1 1 21098
0 21100 7 1 2 55585 21099
0 21101 5 1 1 21100
0 21102 7 1 2 20571 21101
0 21103 7 1 2 20239 21102
0 21104 7 2 2 50090 54426
0 21105 7 1 2 67440 68258
0 21106 5 1 1 21105
0 21107 7 2 2 56462 66309
0 21108 7 1 2 66905 68260
0 21109 5 1 1 21108
0 21110 7 1 2 21106 21109
0 21111 5 1 1 21110
0 21112 7 1 2 42201 21111
0 21113 5 1 1 21112
0 21114 7 1 2 45748 67620
0 21115 7 1 2 68261 21114
0 21116 5 1 1 21115
0 21117 7 1 2 21113 21116
0 21118 5 1 1 21117
0 21119 7 1 2 46844 21118
0 21120 5 1 1 21119
0 21121 7 2 2 42404 53647
0 21122 7 1 2 45749 68259
0 21123 7 1 2 68262 21122
0 21124 5 1 1 21123
0 21125 7 1 2 21120 21124
0 21126 5 1 1 21125
0 21127 7 1 2 46263 21126
0 21128 5 1 1 21127
0 21129 7 2 2 45456 53673
0 21130 7 1 2 42405 54427
0 21131 7 1 2 50269 21130
0 21132 7 1 2 68264 21131
0 21133 5 1 1 21132
0 21134 7 1 2 21128 21133
0 21135 5 1 1 21134
0 21136 7 1 2 45585 21135
0 21137 5 1 1 21136
0 21138 7 2 2 58118 65657
0 21139 5 1 1 68266
0 21140 7 1 2 66940 68267
0 21141 7 1 2 67578 21140
0 21142 5 1 1 21141
0 21143 7 1 2 21137 21142
0 21144 5 1 1 21143
0 21145 7 2 2 42302 44456
0 21146 7 1 2 48003 68268
0 21147 7 1 2 21144 21146
0 21148 5 1 1 21147
0 21149 7 1 2 66622 67360
0 21150 5 1 1 21149
0 21151 7 1 2 58427 67391
0 21152 7 1 2 58380 21151
0 21153 5 1 1 21152
0 21154 7 1 2 21150 21153
0 21155 5 1 1 21154
0 21156 7 1 2 56873 58943
0 21157 7 1 2 63113 21156
0 21158 7 1 2 21155 21157
0 21159 5 1 1 21158
0 21160 7 1 2 21148 21159
0 21161 5 1 1 21160
0 21162 7 1 2 48254 21161
0 21163 5 1 1 21162
0 21164 7 1 2 66540 67760
0 21165 5 1 1 21164
0 21166 7 2 2 44661 66482
0 21167 7 1 2 50162 57289
0 21168 7 1 2 56959 21167
0 21169 7 1 2 68270 21168
0 21170 5 1 1 21169
0 21171 7 1 2 21165 21170
0 21172 5 1 1 21171
0 21173 7 1 2 55618 21172
0 21174 5 1 1 21173
0 21175 7 1 2 55903 66493
0 21176 7 1 2 67645 21175
0 21177 5 1 1 21176
0 21178 7 1 2 21174 21177
0 21179 5 1 1 21178
0 21180 7 1 2 46930 21179
0 21181 5 1 1 21180
0 21182 7 7 2 44662 48255
0 21183 7 2 2 45829 68272
0 21184 7 1 2 55932 68279
0 21185 7 1 2 66702 21184
0 21186 5 1 1 21185
0 21187 7 1 2 21181 21186
0 21188 5 1 1 21187
0 21189 7 1 2 45750 21188
0 21190 5 1 1 21189
0 21191 7 1 2 63732 64524
0 21192 7 1 2 67655 21191
0 21193 5 1 1 21192
0 21194 7 1 2 21190 21193
0 21195 5 1 1 21194
0 21196 7 1 2 45586 21195
0 21197 5 1 1 21196
0 21198 7 1 2 46845 64683
0 21199 7 3 2 64525 21198
0 21200 7 1 2 67769 68281
0 21201 5 1 1 21200
0 21202 7 1 2 21197 21201
0 21203 5 1 1 21202
0 21204 7 1 2 67433 21203
0 21205 5 1 1 21204
0 21206 7 1 2 54056 58704
0 21207 7 1 2 67930 21206
0 21208 7 2 2 61268 66730
0 21209 7 2 2 53163 57612
0 21210 7 1 2 68284 68286
0 21211 7 1 2 21207 21210
0 21212 5 1 1 21211
0 21213 7 1 2 21205 21212
0 21214 7 1 2 21163 21213
0 21215 5 1 1 21214
0 21216 7 1 2 54285 21215
0 21217 5 1 1 21216
0 21218 7 2 2 44457 45087
0 21219 7 2 2 51644 68288
0 21220 7 1 2 67113 68290
0 21221 5 1 1 21220
0 21222 7 1 2 52120 66626
0 21223 7 1 2 57446 21222
0 21224 5 1 1 21223
0 21225 7 1 2 21221 21224
0 21226 5 1 1 21225
0 21227 7 1 2 45587 21226
0 21228 5 1 1 21227
0 21229 7 1 2 56177 67764
0 21230 7 1 2 68291 21229
0 21231 5 1 1 21230
0 21232 7 1 2 21228 21231
0 21233 5 1 1 21232
0 21234 7 1 2 45457 21233
0 21235 5 1 1 21234
0 21236 7 1 2 46846 52121
0 21237 7 2 2 68005 21236
0 21238 7 1 2 57985 68292
0 21239 5 1 1 21238
0 21240 7 1 2 21235 21239
0 21241 5 1 1 21240
0 21242 7 1 2 54725 21241
0 21243 5 1 1 21242
0 21244 7 1 2 55325 55461
0 21245 7 1 2 67875 68006
0 21246 7 1 2 21244 21245
0 21247 5 1 1 21246
0 21248 7 1 2 21243 21247
0 21249 5 1 1 21248
0 21250 7 1 2 43320 21249
0 21251 5 1 1 21250
0 21252 7 1 2 50205 58319
0 21253 5 1 1 21252
0 21254 7 1 2 57395 60898
0 21255 5 1 1 21254
0 21256 7 1 2 21253 21255
0 21257 5 1 1 21256
0 21258 7 1 2 46503 21257
0 21259 5 1 1 21258
0 21260 7 1 2 57406 66862
0 21261 5 1 1 21260
0 21262 7 1 2 21259 21261
0 21263 5 1 1 21262
0 21264 7 1 2 68293 21263
0 21265 5 1 1 21264
0 21266 7 1 2 21251 21265
0 21267 5 1 1 21266
0 21268 7 1 2 66409 21267
0 21269 5 1 1 21268
0 21270 7 1 2 54916 66310
0 21271 5 1 1 21270
0 21272 7 1 2 51233 67723
0 21273 5 1 1 21272
0 21274 7 1 2 21271 21273
0 21275 5 1 1 21274
0 21276 7 1 2 48442 57501
0 21277 7 1 2 61169 66403
0 21278 7 1 2 66866 21277
0 21279 7 1 2 21276 21278
0 21280 7 1 2 21275 21279
0 21281 5 1 1 21280
0 21282 7 1 2 21269 21281
0 21283 5 1 1 21282
0 21284 7 1 2 53592 21283
0 21285 5 1 1 21284
0 21286 7 3 2 46264 60023
0 21287 7 1 2 68285 68294
0 21288 7 1 2 67721 21287
0 21289 5 1 1 21288
0 21290 7 3 2 48004 58135
0 21291 7 1 2 55782 66315
0 21292 7 1 2 68297 21291
0 21293 7 1 2 67733 21292
0 21294 5 1 1 21293
0 21295 7 1 2 21289 21294
0 21296 7 1 2 21285 21295
0 21297 7 1 2 21217 21296
0 21298 5 1 1 21297
0 21299 7 1 2 47664 21298
0 21300 5 1 1 21299
0 21301 7 1 2 66541 67194
0 21302 5 1 1 21301
0 21303 7 2 2 58898 66572
0 21304 7 1 2 50163 58025
0 21305 7 1 2 68300 21304
0 21306 5 1 1 21305
0 21307 7 1 2 21302 21306
0 21308 5 1 1 21307
0 21309 7 1 2 55619 21308
0 21310 5 1 1 21309
0 21311 7 2 2 51527 66805
0 21312 7 1 2 60520 68302
0 21313 5 1 1 21312
0 21314 7 1 2 21310 21313
0 21315 5 1 1 21314
0 21316 7 1 2 53309 21315
0 21317 5 1 1 21316
0 21318 7 1 2 67200 68303
0 21319 5 1 1 21318
0 21320 7 1 2 21317 21319
0 21321 5 1 1 21320
0 21322 7 1 2 45588 21321
0 21323 5 1 1 21322
0 21324 7 1 2 58125 64615
0 21325 7 1 2 66709 21324
0 21326 5 1 1 21325
0 21327 7 1 2 21323 21326
0 21328 5 1 1 21327
0 21329 7 1 2 47665 21328
0 21330 5 1 1 21329
0 21331 7 1 2 42303 63652
0 21332 7 1 2 64497 21331
0 21333 5 1 1 21332
0 21334 7 1 2 63114 67148
0 21335 7 1 2 67318 21334
0 21336 5 1 1 21335
0 21337 7 1 2 21333 21336
0 21338 5 1 1 21337
0 21339 7 1 2 42828 21338
0 21340 5 1 1 21339
0 21341 7 3 2 61435 64715
0 21342 5 1 1 68304
0 21343 7 2 2 62510 68305
0 21344 5 2 1 68307
0 21345 7 1 2 45589 63842
0 21346 7 1 2 68271 21345
0 21347 5 1 1 21346
0 21348 7 1 2 68309 21347
0 21349 5 1 1 21348
0 21350 7 1 2 63493 21349
0 21351 5 1 1 21350
0 21352 7 1 2 21340 21351
0 21353 5 1 1 21352
0 21354 7 1 2 53310 21353
0 21355 5 1 1 21354
0 21356 7 1 2 45751 55739
0 21357 5 1 1 21356
0 21358 7 1 2 53560 55710
0 21359 5 1 1 21358
0 21360 7 1 2 21357 21359
0 21361 5 1 1 21360
0 21362 7 1 2 61450 66122
0 21363 7 1 2 21361 21362
0 21364 5 1 1 21363
0 21365 7 1 2 51820 63399
0 21366 7 1 2 66440 21365
0 21367 7 1 2 63785 21366
0 21368 5 1 1 21367
0 21369 7 1 2 21364 21368
0 21370 5 1 1 21369
0 21371 7 1 2 55586 21370
0 21372 5 1 1 21371
0 21373 7 3 2 61026 64024
0 21374 7 1 2 46931 68311
0 21375 5 1 1 21374
0 21376 7 9 2 46693 43542
0 21377 7 1 2 66722 68314
0 21378 5 1 1 21377
0 21379 7 1 2 21375 21378
0 21380 5 1 1 21379
0 21381 7 1 2 59225 64890
0 21382 7 1 2 21380 21381
0 21383 5 1 1 21382
0 21384 7 1 2 21372 21383
0 21385 7 1 2 21355 21384
0 21386 5 1 1 21385
0 21387 7 1 2 59480 21386
0 21388 5 1 1 21387
0 21389 7 2 2 45830 49990
0 21390 7 2 2 61649 68323
0 21391 7 1 2 61484 68325
0 21392 5 1 1 21391
0 21393 7 1 2 60537 66542
0 21394 7 1 2 66816 21393
0 21395 5 1 1 21394
0 21396 7 1 2 21392 21395
0 21397 5 1 1 21396
0 21398 7 1 2 53674 21397
0 21399 5 1 1 21398
0 21400 7 3 2 44228 57942
0 21401 7 4 2 43321 55760
0 21402 7 1 2 63115 68330
0 21403 7 1 2 68327 21402
0 21404 7 1 2 63855 21403
0 21405 5 1 1 21404
0 21406 7 1 2 21399 21405
0 21407 7 1 2 21388 21406
0 21408 5 1 1 21407
0 21409 7 1 2 67361 21408
0 21410 5 1 1 21409
0 21411 7 2 2 66818 67979
0 21412 7 1 2 45831 68334
0 21413 5 1 1 21412
0 21414 7 1 2 66846 21413
0 21415 5 1 1 21414
0 21416 7 1 2 54778 21415
0 21417 5 1 1 21416
0 21418 7 4 2 44458 51563
0 21419 7 2 2 64644 68336
0 21420 5 1 1 68340
0 21421 7 1 2 44229 68341
0 21422 5 1 1 21421
0 21423 7 1 2 51762 66878
0 21424 5 1 1 21423
0 21425 7 1 2 21422 21424
0 21426 5 1 1 21425
0 21427 7 1 2 59844 21426
0 21428 5 1 1 21427
0 21429 7 1 2 21417 21428
0 21430 5 1 1 21429
0 21431 7 1 2 53593 21430
0 21432 5 1 1 21431
0 21433 7 1 2 66811 21432
0 21434 7 1 2 21410 21433
0 21435 7 1 2 21330 21434
0 21436 5 1 1 21435
0 21437 7 1 2 67434 21436
0 21438 5 1 1 21437
0 21439 7 1 2 56491 66731
0 21440 5 1 1 21439
0 21441 7 1 2 57930 66316
0 21442 5 1 1 21441
0 21443 7 1 2 21440 21442
0 21444 5 1 1 21443
0 21445 7 1 2 66898 21444
0 21446 5 1 1 21445
0 21447 7 2 2 48898 62697
0 21448 7 1 2 56434 68185
0 21449 7 1 2 68342 21448
0 21450 5 1 1 21449
0 21451 7 1 2 21446 21450
0 21452 5 1 1 21451
0 21453 7 1 2 53594 21452
0 21454 5 1 1 21453
0 21455 7 2 2 50511 60181
0 21456 7 1 2 65432 66732
0 21457 7 1 2 68344 21456
0 21458 7 1 2 53703 21457
0 21459 5 1 1 21458
0 21460 7 1 2 21454 21459
0 21461 5 1 1 21460
0 21462 7 1 2 50850 21461
0 21463 5 1 1 21462
0 21464 7 3 2 44459 53595
0 21465 7 5 2 51564 63827
0 21466 7 1 2 42829 55587
0 21467 7 1 2 68349 21466
0 21468 5 1 1 21467
0 21469 7 2 2 51343 54501
0 21470 7 1 2 45832 59453
0 21471 7 1 2 68354 21470
0 21472 5 1 1 21471
0 21473 7 1 2 21468 21472
0 21474 5 1 1 21473
0 21475 7 1 2 45590 21474
0 21476 5 1 1 21475
0 21477 7 1 2 60424 64684
0 21478 7 1 2 68355 21477
0 21479 5 1 1 21478
0 21480 7 1 2 21476 21479
0 21481 5 1 1 21480
0 21482 7 1 2 45458 21481
0 21483 5 1 1 21482
0 21484 7 3 2 61451 63828
0 21485 7 1 2 51565 66292
0 21486 7 1 2 68356 21485
0 21487 5 1 1 21486
0 21488 7 1 2 21483 21487
0 21489 5 1 1 21488
0 21490 7 1 2 68346 21489
0 21491 5 1 1 21490
0 21492 7 1 2 51665 63988
0 21493 7 1 2 66312 21492
0 21494 5 1 1 21493
0 21495 7 1 2 21491 21494
0 21496 5 1 1 21495
0 21497 7 1 2 68023 21496
0 21498 5 1 1 21497
0 21499 7 1 2 21463 21498
0 21500 7 1 2 21438 21499
0 21501 5 1 1 21500
0 21502 7 1 2 54874 21501
0 21503 5 1 1 21502
0 21504 7 12 2 44663 66573
0 21505 7 1 2 54286 58416
0 21506 7 1 2 67399 21505
0 21507 5 1 1 21506
0 21508 7 1 2 49222 67747
0 21509 7 1 2 65364 21508
0 21510 5 1 1 21509
0 21511 7 1 2 21507 21510
0 21512 5 1 1 21511
0 21513 7 1 2 46694 21512
0 21514 5 1 1 21513
0 21515 7 2 2 45915 43322
0 21516 7 1 2 47293 68371
0 21517 7 1 2 67612 21516
0 21518 5 1 1 21517
0 21519 7 1 2 21514 21518
0 21520 5 1 1 21519
0 21521 7 1 2 68359 21520
0 21522 5 1 1 21521
0 21523 7 2 2 54287 67435
0 21524 7 1 2 64716 64152
0 21525 7 1 2 68373 21524
0 21526 5 1 1 21525
0 21527 7 1 2 21522 21526
0 21528 5 1 1 21527
0 21529 7 1 2 53704 21528
0 21530 5 1 1 21529
0 21531 7 1 2 62835 66867
0 21532 7 1 2 52319 21531
0 21533 7 1 2 56281 21532
0 21534 7 1 2 68374 21533
0 21535 5 1 1 21534
0 21536 7 1 2 21530 21535
0 21537 5 1 1 21536
0 21538 7 1 2 67583 21537
0 21539 5 1 1 21538
0 21540 7 1 2 21503 21539
0 21541 7 1 2 21300 21540
0 21542 5 1 1 21541
0 21543 7 1 2 50469 20709
0 21544 5 1 1 21543
0 21545 7 1 2 66149 18861
0 21546 7 1 2 21544 21545
0 21547 7 1 2 21542 21546
0 21548 5 1 1 21547
0 21549 7 1 2 50673 53118
0 21550 7 2 2 63428 21549
0 21551 7 1 2 68190 68375
0 21552 5 1 1 21551
0 21553 7 1 2 47776 57764
0 21554 7 1 2 57867 21553
0 21555 7 1 2 67427 21554
0 21556 5 1 1 21555
0 21557 7 1 2 21552 21556
0 21558 5 1 1 21557
0 21559 7 1 2 45916 21558
0 21560 5 1 1 21559
0 21561 7 5 2 47025 44460
0 21562 7 3 2 42202 66037
0 21563 7 1 2 68377 68382
0 21564 7 1 2 68376 21563
0 21565 5 1 1 21564
0 21566 7 1 2 21560 21565
0 21567 5 1 1 21566
0 21568 7 1 2 48256 21567
0 21569 5 1 1 21568
0 21570 7 1 2 56456 58004
0 21571 7 1 2 63429 21570
0 21572 7 1 2 67907 68383
0 21573 7 1 2 21571 21572
0 21574 5 1 1 21573
0 21575 7 1 2 21569 21574
0 21576 5 1 1 21575
0 21577 7 1 2 42027 21576
0 21578 5 1 1 21577
0 21579 7 1 2 43465 52582
0 21580 7 1 2 55483 65433
0 21581 7 1 2 67985 21580
0 21582 7 1 2 21579 21581
0 21583 7 1 2 67411 21582
0 21584 5 1 1 21583
0 21585 7 1 2 21578 21584
0 21586 5 1 1 21585
0 21587 7 1 2 44664 21586
0 21588 5 1 1 21587
0 21589 7 1 2 44915 51886
0 21590 7 1 2 66251 21589
0 21591 7 2 2 59964 66038
0 21592 7 1 2 63547 68385
0 21593 7 1 2 21590 21592
0 21594 7 1 2 65296 21593
0 21595 5 1 1 21594
0 21596 7 1 2 21588 21595
0 21597 5 1 1 21596
0 21598 7 1 2 48125 21597
0 21599 5 1 1 21598
0 21600 7 1 2 65282 67677
0 21601 5 1 1 21600
0 21602 7 1 2 53119 68058
0 21603 5 1 1 21602
0 21604 7 1 2 21601 21603
0 21605 5 1 1 21604
0 21606 7 1 2 67457 21605
0 21607 5 1 1 21606
0 21608 7 1 2 54598 68032
0 21609 5 1 1 21608
0 21610 7 1 2 21607 21609
0 21611 5 1 1 21610
0 21612 7 1 2 43596 21611
0 21613 5 1 1 21612
0 21614 7 1 2 50721 54624
0 21615 7 1 2 66255 21614
0 21616 5 1 1 21615
0 21617 7 1 2 21613 21616
0 21618 5 1 1 21617
0 21619 7 2 2 48937 58218
0 21620 7 4 2 48899 52784
0 21621 7 1 2 54966 68389
0 21622 7 1 2 68387 21621
0 21623 7 1 2 21618 21622
0 21624 5 1 1 21623
0 21625 7 1 2 21599 21624
0 21626 5 1 1 21625
0 21627 7 1 2 42304 21626
0 21628 5 1 1 21627
0 21629 7 1 2 43753 66775
0 21630 5 1 1 21629
0 21631 7 1 2 51180 67876
0 21632 5 1 1 21631
0 21633 7 1 2 21630 21632
0 21634 5 1 1 21633
0 21635 7 1 2 64302 66039
0 21636 7 1 2 56518 21635
0 21637 7 1 2 68192 21636
0 21638 7 1 2 21634 21637
0 21639 5 1 1 21638
0 21640 7 1 2 21628 21639
0 21641 5 1 1 21640
0 21642 7 1 2 44332 21641
0 21643 5 1 1 21642
0 21644 7 1 2 54004 58294
0 21645 7 1 2 67418 21644
0 21646 7 1 2 68247 21645
0 21647 5 1 1 21646
0 21648 7 1 2 48443 58005
0 21649 7 1 2 67392 21648
0 21650 7 1 2 67350 21649
0 21651 5 1 1 21650
0 21652 7 1 2 21647 21651
0 21653 5 1 1 21652
0 21654 7 1 2 45752 21653
0 21655 5 1 1 21654
0 21656 7 1 2 55018 60039
0 21657 7 1 2 63075 67565
0 21658 7 1 2 21656 21657
0 21659 7 1 2 68025 21658
0 21660 5 1 1 21659
0 21661 7 1 2 21655 21660
0 21662 5 1 1 21661
0 21663 7 2 2 54967 64076
0 21664 7 1 2 65690 67356
0 21665 7 1 2 68393 21664
0 21666 7 1 2 21662 21665
0 21667 5 1 1 21666
0 21668 7 1 2 21643 21667
0 21669 5 1 1 21668
0 21670 7 1 2 51800 21669
0 21671 5 1 1 21670
0 21672 7 1 2 61809 67423
0 21673 5 1 1 21672
0 21674 7 1 2 61933 67412
0 21675 5 1 1 21674
0 21676 7 1 2 21673 21675
0 21677 5 1 1 21676
0 21678 7 1 2 65899 21677
0 21679 5 1 1 21678
0 21680 7 1 2 46847 51821
0 21681 7 1 2 59750 21680
0 21682 7 8 2 44665 64110
0 21683 7 1 2 67039 68395
0 21684 7 1 2 21681 21683
0 21685 5 1 1 21684
0 21686 7 1 2 21679 21685
0 21687 5 1 1 21686
0 21688 7 1 2 45591 21687
0 21689 5 1 1 21688
0 21690 7 1 2 65813 67430
0 21691 5 1 1 21690
0 21692 7 1 2 21689 21691
0 21693 5 1 1 21692
0 21694 7 1 2 47777 21693
0 21695 5 1 1 21694
0 21696 7 1 2 61566 62476
0 21697 7 1 2 68224 21696
0 21698 7 1 2 65532 21697
0 21699 5 1 1 21698
0 21700 7 1 2 21695 21699
0 21701 5 1 1 21700
0 21702 7 1 2 45459 21701
0 21703 5 1 1 21702
0 21704 7 1 2 45592 67428
0 21705 5 1 1 21704
0 21706 7 1 2 19989 21705
0 21707 5 1 1 21706
0 21708 7 1 2 61358 64111
0 21709 7 1 2 21707 21708
0 21710 5 1 1 21709
0 21711 7 1 2 21703 21710
0 21712 5 1 1 21711
0 21713 7 1 2 47560 21712
0 21714 5 1 1 21713
0 21715 7 1 2 61095 64395
0 21716 7 1 2 67376 21715
0 21717 7 2 2 58960 21716
0 21718 5 1 1 68403
0 21719 7 4 2 53596 60325
0 21720 7 1 2 45593 60230
0 21721 7 2 2 60877 21720
0 21722 5 1 1 68409
0 21723 7 1 2 68405 68410
0 21724 5 1 1 21723
0 21725 7 2 2 43466 46986
0 21726 7 1 2 68230 68411
0 21727 5 1 1 21726
0 21728 7 2 2 48900 63943
0 21729 7 1 2 68406 68413
0 21730 5 1 1 21729
0 21731 7 1 2 21727 21730
0 21732 5 1 1 21731
0 21733 7 1 2 44333 62150
0 21734 7 1 2 21732 21733
0 21735 5 1 1 21734
0 21736 7 1 2 21724 21735
0 21737 5 1 1 21736
0 21738 7 1 2 43635 21737
0 21739 5 1 1 21738
0 21740 7 1 2 21718 21739
0 21741 5 1 1 21740
0 21742 7 1 2 64526 21741
0 21743 5 1 1 21742
0 21744 7 1 2 21714 21743
0 21745 5 1 1 21744
0 21746 7 1 2 46695 21745
0 21747 5 1 1 21746
0 21748 7 1 2 46504 50470
0 21749 7 1 2 53164 21748
0 21750 7 1 2 67233 21749
0 21751 5 1 1 21750
0 21752 7 1 2 21722 21751
0 21753 5 1 1 21752
0 21754 7 1 2 47561 21753
0 21755 5 1 1 21754
0 21756 7 1 2 53744 58886
0 21757 7 1 2 67464 21756
0 21758 5 1 1 21757
0 21759 7 1 2 21755 21758
0 21760 5 1 1 21759
0 21761 7 1 2 68407 21760
0 21762 5 1 1 21761
0 21763 7 1 2 43754 58359
0 21764 5 1 1 21763
0 21765 7 1 2 20260 21764
0 21766 5 1 1 21765
0 21767 7 7 2 45833 43543
0 21768 7 1 2 61854 67529
0 21769 7 1 2 68415 21768
0 21770 7 1 2 68414 21769
0 21771 7 1 2 21766 21770
0 21772 5 1 1 21771
0 21773 7 1 2 21762 21772
0 21774 5 1 1 21773
0 21775 7 1 2 43636 21774
0 21776 5 1 1 21775
0 21777 7 1 2 47562 68404
0 21778 5 1 1 21777
0 21779 7 1 2 21776 21778
0 21780 5 1 1 21779
0 21781 7 1 2 64527 21780
0 21782 5 1 1 21781
0 21783 7 1 2 60793 67285
0 21784 7 1 2 62047 21783
0 21785 7 1 2 65497 66999
0 21786 7 1 2 67681 21785
0 21787 7 1 2 21784 21786
0 21788 5 1 1 21787
0 21789 7 1 2 21782 21788
0 21790 7 1 2 21747 21789
0 21791 5 1 1 21790
0 21792 7 1 2 48257 21791
0 21793 5 1 1 21792
0 21794 7 1 2 51060 57311
0 21795 5 1 1 21794
0 21796 7 1 2 19871 21795
0 21797 5 1 1 21796
0 21798 7 2 2 60339 21797
0 21799 7 1 2 54435 56236
0 21800 7 1 2 68378 21799
0 21801 7 1 2 67532 21800
0 21802 7 1 2 68422 21801
0 21803 5 1 1 21802
0 21804 7 1 2 47906 21803
0 21805 7 1 2 21793 21804
0 21806 5 1 1 21805
0 21807 7 3 2 42560 57290
0 21808 7 1 2 65425 67404
0 21809 7 1 2 54779 21808
0 21810 7 1 2 68424 21809
0 21811 5 1 1 21810
0 21812 7 1 2 49223 68379
0 21813 7 1 2 64569 21812
0 21814 7 1 2 67450 21813
0 21815 5 1 1 21814
0 21816 7 1 2 21811 21815
0 21817 5 1 1 21816
0 21818 7 1 2 46696 21817
0 21819 5 1 1 21818
0 21820 7 1 2 42305 49090
0 21821 7 1 2 68030 21820
0 21822 7 1 2 67451 68213
0 21823 7 1 2 21821 21822
0 21824 5 1 1 21823
0 21825 7 1 2 21819 21824
0 21826 5 1 1 21825
0 21827 7 1 2 46505 21826
0 21828 5 1 1 21827
0 21829 7 2 2 45834 55380
0 21830 7 1 2 43637 49168
0 21831 7 1 2 52137 21830
0 21832 7 1 2 68427 21831
0 21833 5 1 1 21832
0 21834 7 2 2 42306 47129
0 21835 7 1 2 67865 68429
0 21836 7 1 2 65302 21835
0 21837 5 1 1 21836
0 21838 7 1 2 21833 21837
0 21839 5 1 1 21838
0 21840 7 1 2 55862 62511
0 21841 7 1 2 21839 21840
0 21842 5 1 1 21841
0 21843 7 1 2 21828 21842
0 21844 5 1 1 21843
0 21845 7 1 2 59677 21844
0 21846 5 1 1 21845
0 21847 7 1 2 64459 67405
0 21848 7 1 2 59784 21847
0 21849 7 1 2 67649 21848
0 21850 5 1 1 21849
0 21851 7 1 2 21846 21850
0 21852 5 1 1 21851
0 21853 7 1 2 43597 21852
0 21854 5 1 1 21853
0 21855 7 2 2 50164 55653
0 21856 7 1 2 64382 67406
0 21857 7 1 2 68431 21856
0 21858 7 2 2 42028 66988
0 21859 7 2 2 55904 59678
0 21860 7 1 2 68433 68435
0 21861 7 1 2 21857 21860
0 21862 5 1 1 21861
0 21863 7 1 2 21854 21862
0 21864 5 1 1 21863
0 21865 7 1 2 52785 21864
0 21866 5 1 1 21865
0 21867 7 1 2 45753 67351
0 21868 5 1 1 21867
0 21869 7 1 2 58758 67377
0 21870 5 1 1 21869
0 21871 7 1 2 21868 21870
0 21872 5 1 1 21871
0 21873 7 1 2 63321 67650
0 21874 5 1 1 21873
0 21875 7 2 2 63767 64540
0 21876 7 1 2 67761 68437
0 21877 5 1 1 21876
0 21878 7 1 2 21874 21877
0 21879 5 1 1 21878
0 21880 7 1 2 45594 21879
0 21881 5 1 1 21880
0 21882 7 2 2 42307 54743
0 21883 7 1 2 67651 68439
0 21884 5 1 1 21883
0 21885 7 1 2 21881 21884
0 21886 5 1 1 21885
0 21887 7 1 2 47666 21886
0 21888 5 1 1 21887
0 21889 7 9 2 59394 65900
0 21890 7 1 2 48258 66330
0 21891 7 1 2 68441 21890
0 21892 5 1 1 21891
0 21893 7 1 2 21888 21892
0 21894 5 1 1 21893
0 21895 7 1 2 21872 21894
0 21896 5 1 1 21895
0 21897 7 1 2 44582 21896
0 21898 7 1 2 21866 21897
0 21899 5 1 1 21898
0 21900 7 1 2 54288 21899
0 21901 7 1 2 21806 21900
0 21902 5 1 1 21901
0 21903 7 1 2 66237 68040
0 21904 5 1 1 21903
0 21905 7 1 2 51979 66252
0 21906 7 1 2 60126 21905
0 21907 5 1 1 21906
0 21908 7 1 2 21904 21907
0 21909 5 1 1 21908
0 21910 7 1 2 42308 21909
0 21911 5 1 1 21910
0 21912 7 3 2 44230 53467
0 21913 5 1 1 68450
0 21914 7 1 2 58307 64616
0 21915 7 1 2 66060 21914
0 21916 7 1 2 68451 21915
0 21917 5 1 1 21916
0 21918 7 1 2 21911 21917
0 21919 5 1 1 21918
0 21920 7 1 2 50471 21919
0 21921 5 1 1 21920
0 21922 7 6 2 42309 47294
0 21923 7 1 2 54846 66238
0 21924 7 1 2 68453 21923
0 21925 7 1 2 53011 21924
0 21926 5 1 1 21925
0 21927 7 1 2 21921 21926
0 21928 5 1 1 21927
0 21929 7 1 2 43105 21928
0 21930 5 1 1 21929
0 21931 7 1 2 64112 66239
0 21932 7 1 2 67319 21931
0 21933 7 1 2 65297 21932
0 21934 5 1 1 21933
0 21935 7 1 2 21930 21934
0 21936 5 1 1 21935
0 21937 7 1 2 44583 21936
0 21938 5 1 1 21937
0 21939 7 3 2 47026 45088
0 21940 7 1 2 60312 68459
0 21941 7 1 2 68042 21940
0 21942 7 1 2 67495 21941
0 21943 5 1 1 21942
0 21944 7 1 2 21938 21943
0 21945 5 1 1 21944
0 21946 7 1 2 44916 21945
0 21947 5 1 1 21946
0 21948 7 1 2 51842 58010
0 21949 7 1 2 67867 21948
0 21950 7 1 2 2182 56370
0 21951 5 1 1 21950
0 21952 7 1 2 60340 68432
0 21953 7 1 2 21951 21952
0 21954 7 1 2 21949 21953
0 21955 5 1 1 21954
0 21956 7 1 2 21947 21955
0 21957 5 1 1 21956
0 21958 7 1 2 48005 21957
0 21959 5 1 1 21958
0 21960 7 1 2 66253 67241
0 21961 5 1 1 21960
0 21962 7 1 2 66240 67212
0 21963 5 1 1 21962
0 21964 7 1 2 21961 21963
0 21965 5 1 1 21964
0 21966 7 1 2 45835 21965
0 21967 5 1 1 21966
0 21968 7 1 2 52450 66138
0 21969 7 1 2 68454 21968
0 21970 5 1 1 21969
0 21971 7 1 2 21967 21970
0 21972 5 1 1 21971
0 21973 7 1 2 46265 61214
0 21974 7 1 2 67496 21973
0 21975 7 1 2 21972 21974
0 21976 5 1 1 21975
0 21977 7 1 2 21959 21976
0 21978 5 1 1 21977
0 21979 7 1 2 43544 21978
0 21980 5 1 1 21979
0 21981 7 1 2 67258 67863
0 21982 5 1 1 21981
0 21983 7 1 2 68110 68460
0 21984 7 1 2 68043 21983
0 21985 5 1 1 21984
0 21986 7 1 2 21982 21985
0 21987 5 1 1 21986
0 21988 7 1 2 43598 67497
0 21989 7 2 2 21987 21988
0 21990 7 1 2 65620 68462
0 21991 5 1 1 21990
0 21992 7 1 2 21980 21991
0 21993 5 1 1 21992
0 21994 7 1 2 42203 21993
0 21995 5 1 1 21994
0 21996 7 1 2 68143 68463
0 21997 5 1 1 21996
0 21998 7 1 2 21995 21997
0 21999 5 1 1 21998
0 22000 7 1 2 65661 21999
0 22001 5 1 1 22000
0 22002 7 1 2 48901 56215
0 22003 7 1 2 61304 22002
0 22004 7 1 2 66598 67268
0 22005 7 1 2 22003 22004
0 22006 5 1 1 22005
0 22007 7 1 2 59090 66899
0 22008 5 1 1 22007
0 22009 7 3 2 59481 59664
0 22010 7 1 2 65303 68464
0 22011 5 1 1 22010
0 22012 7 1 2 67250 22011
0 22013 7 1 2 22008 22012
0 22014 5 1 1 22013
0 22015 7 2 2 56917 63289
0 22016 7 1 2 46987 68467
0 22017 7 1 2 22014 22016
0 22018 5 1 1 22017
0 22019 7 1 2 22006 22018
0 22020 5 1 1 22019
0 22021 7 1 2 48006 22020
0 22022 5 1 1 22021
0 22023 7 1 2 61325 67980
0 22024 5 1 1 22023
0 22025 7 1 2 51535 61316
0 22026 5 1 1 22025
0 22027 7 1 2 22024 22026
0 22028 5 2 1 22027
0 22029 7 1 2 42029 68469
0 22030 5 1 1 22029
0 22031 7 1 2 55905 59574
0 22032 7 1 2 67981 22031
0 22033 5 1 1 22032
0 22034 7 1 2 22030 22033
0 22035 5 1 1 22034
0 22036 7 3 2 44666 63076
0 22037 7 1 2 64396 68471
0 22038 7 1 2 22035 22037
0 22039 5 1 1 22038
0 22040 7 1 2 22022 22039
0 22041 5 1 1 22040
0 22042 7 1 2 67286 22041
0 22043 5 1 1 22042
0 22044 7 1 2 65691 68470
0 22045 5 1 1 22044
0 22046 7 5 2 48007 60642
0 22047 7 2 2 65829 68474
0 22048 7 1 2 59040 68479
0 22049 5 1 1 22048
0 22050 7 1 2 22045 22049
0 22051 5 1 1 22050
0 22052 7 1 2 45595 22051
0 22053 5 1 1 22052
0 22054 7 1 2 49991 66092
0 22055 5 2 1 22054
0 22056 7 2 2 50851 66985
0 22057 5 1 1 68483
0 22058 7 1 2 68481 22057
0 22059 5 1 1 22058
0 22060 7 1 2 61330 22059
0 22061 5 1 1 22060
0 22062 7 1 2 22053 22061
0 22063 5 1 1 22062
0 22064 7 1 2 67571 22063
0 22065 5 1 1 22064
0 22066 7 1 2 22043 22065
0 22067 5 1 1 22066
0 22068 7 1 2 44584 22067
0 22069 5 1 1 22068
0 22070 7 2 2 44667 60182
0 22071 7 1 2 60047 64444
0 22072 7 1 2 68380 22071
0 22073 7 1 2 68485 22072
0 22074 7 1 2 68423 22073
0 22075 5 1 1 22074
0 22076 7 1 2 22069 22075
0 22077 5 1 1 22076
0 22078 7 1 2 42204 22077
0 22079 5 1 1 22078
0 22080 7 1 2 65901 67988
0 22081 5 1 1 22080
0 22082 7 2 2 51763 65692
0 22083 5 2 1 68487
0 22084 7 1 2 59845 68488
0 22085 5 1 1 22084
0 22086 7 1 2 22081 22085
0 22087 5 1 1 22086
0 22088 7 1 2 58724 22087
0 22089 5 1 1 22088
0 22090 7 1 2 63994 68335
0 22091 5 1 1 22090
0 22092 7 1 2 66968 22091
0 22093 5 1 1 22092
0 22094 7 1 2 54780 22093
0 22095 5 1 1 22094
0 22096 7 1 2 65994 67996
0 22097 5 1 1 22096
0 22098 7 2 2 64428 68357
0 22099 7 1 2 51528 68491
0 22100 5 1 1 22099
0 22101 7 1 2 22097 22100
0 22102 5 1 1 22101
0 22103 7 1 2 61053 22102
0 22104 5 1 1 22103
0 22105 7 1 2 22095 22104
0 22106 7 1 2 22089 22105
0 22107 5 1 1 22106
0 22108 7 1 2 67352 22107
0 22109 5 1 1 22108
0 22110 7 1 2 51144 67508
0 22111 7 1 2 59109 22110
0 22112 5 1 1 22111
0 22113 7 1 2 42830 67513
0 22114 7 1 2 62310 22113
0 22115 5 1 1 22114
0 22116 7 1 2 22112 22115
0 22117 5 1 1 22116
0 22118 7 1 2 65902 22117
0 22119 5 1 1 22118
0 22120 7 6 2 46697 46932
0 22121 5 1 1 68493
0 22122 7 1 2 63829 68494
0 22123 7 1 2 54395 22122
0 22124 7 2 2 60231 62469
0 22125 7 1 2 67378 68499
0 22126 7 1 2 22123 22125
0 22127 5 1 1 22126
0 22128 7 1 2 22119 22127
0 22129 5 1 1 22128
0 22130 7 1 2 60456 22129
0 22131 5 1 1 22130
0 22132 7 2 2 51519 67002
0 22133 5 2 1 68501
0 22134 7 1 2 60492 68502
0 22135 5 1 1 22134
0 22136 7 1 2 59110 68442
0 22137 5 1 1 22136
0 22138 7 1 2 22135 22137
0 22139 5 1 1 22138
0 22140 7 1 2 67575 22139
0 22141 5 1 1 22140
0 22142 7 1 2 59602 65995
0 22143 7 1 2 67339 68331
0 22144 7 1 2 22142 22143
0 22145 5 1 1 22144
0 22146 7 2 2 55462 64397
0 22147 7 1 2 64429 67962
0 22148 7 1 2 68505 22147
0 22149 7 1 2 51529 22148
0 22150 5 1 1 22149
0 22151 7 1 2 22145 22150
0 22152 5 1 1 22151
0 22153 7 1 2 62512 22152
0 22154 5 1 1 22153
0 22155 7 1 2 22141 22154
0 22156 7 1 2 22131 22155
0 22157 5 1 1 22156
0 22158 7 1 2 51943 22157
0 22159 5 1 1 22158
0 22160 7 1 2 22109 22159
0 22161 7 1 2 22079 22160
0 22162 5 1 1 22161
0 22163 7 1 2 54875 22162
0 22164 5 1 1 22163
0 22165 7 4 2 55484 57913
0 22166 7 2 2 52046 68507
0 22167 7 1 2 63733 68511
0 22168 5 1 1 22167
0 22169 7 2 2 42310 43924
0 22170 7 1 2 60916 68513
0 22171 7 1 2 67672 22170
0 22172 5 1 1 22171
0 22173 7 1 2 22168 22172
0 22174 5 1 1 22173
0 22175 7 1 2 67353 22174
0 22176 5 1 1 22175
0 22177 7 1 2 55072 67119
0 22178 7 2 2 45754 64099
0 22179 7 1 2 68508 68515
0 22180 7 1 2 22177 22179
0 22181 5 1 1 22180
0 22182 7 2 2 46038 65539
0 22183 7 1 2 47027 54005
0 22184 7 1 2 68517 22183
0 22185 7 1 2 67674 22184
0 22186 5 1 1 22185
0 22187 7 1 2 22181 22186
0 22188 7 1 2 22176 22187
0 22189 5 1 1 22188
0 22190 7 1 2 46848 22189
0 22191 5 1 1 22190
0 22192 7 1 2 68026 67737
0 22193 7 2 2 45755 63290
0 22194 7 1 2 68509 68519
0 22195 7 1 2 22192 22194
0 22196 5 1 1 22195
0 22197 7 1 2 22191 22196
0 22198 5 1 1 22197
0 22199 7 1 2 45596 22198
0 22200 5 1 1 22199
0 22201 7 1 2 64296 68021
0 22202 7 4 2 42030 63799
0 22203 7 1 2 68510 68521
0 22204 7 1 2 22201 22203
0 22205 5 1 1 22204
0 22206 7 1 2 22200 22205
0 22207 5 1 1 22206
0 22208 7 1 2 60232 22207
0 22209 5 1 1 22208
0 22210 7 1 2 55265 68065
0 22211 7 1 2 68103 22210
0 22212 5 1 1 22211
0 22213 7 1 2 47028 48938
0 22214 7 1 2 66667 22213
0 22215 7 1 2 67452 22214
0 22216 5 1 1 22215
0 22217 7 1 2 22212 22216
0 22218 5 1 1 22217
0 22219 7 5 2 43467 61605
0 22220 7 1 2 55163 61291
0 22221 7 1 2 68525 22220
0 22222 7 1 2 22218 22221
0 22223 5 1 1 22222
0 22224 7 1 2 22209 22223
0 22225 5 1 1 22224
0 22226 7 1 2 48444 22225
0 22227 5 1 1 22226
0 22228 7 1 2 54625 60417
0 22229 7 1 2 66723 22228
0 22230 7 1 2 67290 68090
0 22231 7 1 2 22229 22230
0 22232 5 1 1 22231
0 22233 7 1 2 50357 68125
0 22234 5 1 1 22233
0 22235 7 1 2 64509 66518
0 22236 5 1 1 22235
0 22237 7 1 2 22234 22236
0 22238 5 1 1 22237
0 22239 7 1 2 54077 68198
0 22240 7 1 2 22238 22239
0 22241 5 1 1 22240
0 22242 7 1 2 22232 22241
0 22243 5 1 1 22242
0 22244 7 1 2 54968 68461
0 22245 7 1 2 22243 22244
0 22246 5 1 1 22245
0 22247 7 1 2 22227 22246
0 22248 5 1 1 22247
0 22249 7 1 2 55588 22248
0 22250 5 1 1 22249
0 22251 7 1 2 65869 67839
0 22252 5 1 1 22251
0 22253 7 5 2 58944 63019
0 22254 7 1 2 46849 68530
0 22255 7 1 2 67298 22254
0 22256 5 1 1 22255
0 22257 7 1 2 22252 22256
0 22258 5 1 1 22257
0 22259 7 1 2 42831 22258
0 22260 5 1 1 22259
0 22261 7 2 2 45460 54781
0 22262 7 1 2 58926 66978
0 22263 7 1 2 68535 22262
0 22264 5 1 1 22263
0 22265 7 1 2 22260 22264
0 22266 5 1 1 22265
0 22267 7 1 2 54605 22266
0 22268 5 1 1 22267
0 22269 7 2 2 44668 49654
0 22270 7 1 2 58920 62201
0 22271 7 1 2 63249 22270
0 22272 7 1 2 68537 22271
0 22273 7 1 2 68536 22272
0 22274 5 1 1 22273
0 22275 7 1 2 22268 22274
0 22276 5 1 1 22275
0 22277 7 1 2 60568 22276
0 22278 5 1 1 22277
0 22279 7 2 2 48445 67299
0 22280 7 1 2 63128 68512
0 22281 7 1 2 68539 22280
0 22282 5 1 1 22281
0 22283 7 1 2 22278 22282
0 22284 5 1 1 22283
0 22285 7 1 2 67354 22284
0 22286 5 1 1 22285
0 22287 7 3 2 44231 54502
0 22288 7 1 2 65540 68541
0 22289 7 1 2 67835 22288
0 22290 5 1 1 22289
0 22291 7 1 2 57396 59298
0 22292 7 1 2 67754 22291
0 22293 5 1 1 22292
0 22294 7 1 2 51944 54917
0 22295 7 1 2 67300 22294
0 22296 5 1 1 22295
0 22297 7 1 2 22293 22296
0 22298 5 1 1 22297
0 22299 7 1 2 48446 65903
0 22300 7 1 2 22298 22299
0 22301 5 1 1 22300
0 22302 7 1 2 22290 22301
0 22303 5 1 1 22302
0 22304 7 1 2 45597 67576
0 22305 5 1 1 22304
0 22306 7 1 2 20858 22305
0 22307 5 1 1 22306
0 22308 7 1 2 44461 22307
0 22309 7 1 2 22303 22308
0 22310 5 1 1 22309
0 22311 7 1 2 58945 67855
0 22312 7 1 2 54661 22311
0 22313 7 1 2 63079 68506
0 22314 7 1 2 22312 22313
0 22315 7 1 2 68540 22314
0 22316 5 1 1 22315
0 22317 7 1 2 22310 22316
0 22318 7 1 2 22286 22317
0 22319 5 1 1 22318
0 22320 7 1 2 47667 22319
0 22321 5 1 1 22320
0 22322 7 1 2 22250 22321
0 22323 7 1 2 22164 22322
0 22324 7 1 2 22001 22323
0 22325 7 1 2 21902 22324
0 22326 5 1 1 22325
0 22327 7 1 2 67436 22326
0 22328 5 1 1 22327
0 22329 7 1 2 21671 22328
0 22330 7 1 2 21548 22329
0 22331 7 1 2 21103 22330
0 22332 7 1 2 18649 22331
0 22333 5 1 1 22332
0 22334 7 1 2 64131 22333
0 22335 5 1 1 22334
0 22336 7 1 2 52492 54592
0 22337 5 7 1 22336
0 22338 7 3 2 49286 68544
0 22339 7 1 2 51431 68551
0 22340 5 3 1 22339
0 22341 7 1 2 53400 67783
0 22342 5 1 1 22341
0 22343 7 1 2 68554 22342
0 22344 5 1 1 22343
0 22345 7 1 2 46266 22344
0 22346 5 1 1 22345
0 22347 7 1 2 52751 58417
0 22348 7 2 2 67784 22347
0 22349 5 1 1 68557
0 22350 7 2 2 22346 22349
0 22351 7 1 2 49620 54057
0 22352 5 1 1 22351
0 22353 7 1 2 49655 52353
0 22354 5 1 1 22353
0 22355 7 1 2 22352 22354
0 22356 5 1 1 22355
0 22357 7 1 2 47295 22356
0 22358 5 2 1 22357
0 22359 7 1 2 49402 52260
0 22360 5 1 1 22359
0 22361 7 1 2 44917 22360
0 22362 5 1 1 22361
0 22363 7 1 2 68561 22362
0 22364 5 1 1 22363
0 22365 7 1 2 46267 22364
0 22366 5 1 1 22365
0 22367 7 1 2 49399 54078
0 22368 5 1 1 22367
0 22369 7 1 2 22366 22368
0 22370 5 1 1 22369
0 22371 7 1 2 51003 22370
0 22372 5 1 1 22371
0 22373 7 1 2 68559 22372
0 22374 5 1 1 22373
0 22375 7 1 2 46039 22374
0 22376 5 1 1 22375
0 22377 7 4 2 50557 54969
0 22378 7 1 2 52451 2115
0 22379 7 1 2 68563 22378
0 22380 7 1 2 57479 22379
0 22381 5 1 1 22380
0 22382 7 1 2 22376 22381
0 22383 5 1 1 22382
0 22384 7 2 2 61558 22383
0 22385 7 1 2 48902 68567
0 22386 5 1 1 22385
0 22387 7 1 2 62882 68014
0 22388 5 1 1 22387
0 22389 7 1 2 52201 52361
0 22390 5 1 1 22389
0 22391 7 1 2 49343 22390
0 22392 5 2 1 22391
0 22393 7 1 2 22388 68569
0 22394 5 1 1 22393
0 22395 7 1 2 60295 22394
0 22396 5 1 1 22395
0 22397 7 1 2 52806 53970
0 22398 5 1 1 22397
0 22399 7 1 2 62318 22398
0 22400 5 1 1 22399
0 22401 7 1 2 57351 22400
0 22402 5 1 1 22401
0 22403 7 1 2 22396 22402
0 22404 5 2 1 22403
0 22405 7 1 2 59785 68571
0 22406 5 1 1 22405
0 22407 7 1 2 42832 58974
0 22408 5 1 1 22407
0 22409 7 1 2 49490 59612
0 22410 7 2 2 22408 22409
0 22411 7 1 2 59955 68573
0 22412 5 1 1 22411
0 22413 7 1 2 22406 22412
0 22414 5 1 1 22413
0 22415 7 1 2 45089 22414
0 22416 5 1 1 22415
0 22417 7 2 2 52849 59786
0 22418 7 1 2 54696 68575
0 22419 5 1 1 22418
0 22420 7 1 2 63921 22419
0 22421 5 1 1 22420
0 22422 7 1 2 44232 22421
0 22423 5 1 1 22422
0 22424 7 1 2 59743 59929
0 22425 5 1 1 22424
0 22426 7 1 2 22423 22425
0 22427 5 1 1 22426
0 22428 7 1 2 43323 22427
0 22429 5 1 1 22428
0 22430 7 1 2 51399 64142
0 22431 5 1 1 22430
0 22432 7 1 2 63710 22431
0 22433 5 1 1 22432
0 22434 7 3 2 48447 22433
0 22435 5 1 1 68577
0 22436 7 1 2 59787 68578
0 22437 5 1 1 22436
0 22438 7 1 2 22429 22437
0 22439 5 1 1 22438
0 22440 7 1 2 47296 22439
0 22441 5 1 1 22440
0 22442 7 2 2 49379 63395
0 22443 7 1 2 68526 68580
0 22444 5 1 1 22443
0 22445 7 1 2 22441 22444
0 22446 5 1 1 22445
0 22447 7 1 2 46268 22446
0 22448 5 1 1 22447
0 22449 7 1 2 22416 22448
0 22450 5 1 1 22449
0 22451 7 1 2 42561 22450
0 22452 5 1 1 22451
0 22453 7 1 2 53063 64887
0 22454 5 4 1 22453
0 22455 7 1 2 68465 68582
0 22456 5 1 1 22455
0 22457 7 1 2 52383 59871
0 22458 5 1 1 22457
0 22459 7 1 2 22456 22458
0 22460 5 1 1 22459
0 22461 7 1 2 42833 22460
0 22462 5 1 1 22461
0 22463 7 1 2 953 55273
0 22464 5 2 1 22463
0 22465 7 3 2 48622 68586
0 22466 7 1 2 59913 68588
0 22467 5 1 1 22466
0 22468 7 1 2 22462 22467
0 22469 5 1 1 22468
0 22470 7 1 2 46040 22469
0 22471 5 1 1 22470
0 22472 7 4 2 45090 60296
0 22473 7 3 2 61972 68591
0 22474 7 1 2 68527 68595
0 22475 5 1 1 22474
0 22476 7 1 2 22471 22475
0 22477 5 1 1 22476
0 22478 7 1 2 44070 22477
0 22479 5 1 1 22478
0 22480 7 2 2 43468 56178
0 22481 7 2 2 47429 68596
0 22482 7 1 2 68598 68600
0 22483 5 1 1 22482
0 22484 7 1 2 22479 22483
0 22485 5 1 1 22484
0 22486 7 1 2 49992 22485
0 22487 5 1 1 22486
0 22488 7 1 2 48259 22487
0 22489 7 1 2 22452 22488
0 22490 5 1 1 22489
0 22491 7 1 2 45091 55129
0 22492 5 1 1 22491
0 22493 7 1 2 2041 22492
0 22494 5 1 1 22493
0 22495 7 2 2 61831 22494
0 22496 7 1 2 59956 68602
0 22497 5 1 1 22496
0 22498 7 1 2 61540 65417
0 22499 5 1 1 22498
0 22500 7 1 2 53120 61741
0 22501 7 2 2 22499 22500
0 22502 7 1 2 58196 68604
0 22503 5 1 1 22502
0 22504 7 1 2 22497 22503
0 22505 5 1 1 22504
0 22506 7 1 2 44233 22505
0 22507 5 1 1 22506
0 22508 7 1 2 48964 58899
0 22509 5 1 1 22508
0 22510 7 1 2 45258 53350
0 22511 5 3 1 22510
0 22512 7 1 2 54715 68606
0 22513 5 1 1 22512
0 22514 7 1 2 22509 22513
0 22515 5 1 1 22514
0 22516 7 1 2 43106 22515
0 22517 5 1 1 22516
0 22518 7 2 2 52850 58789
0 22519 5 1 1 68609
0 22520 7 1 2 60069 22519
0 22521 5 1 1 22520
0 22522 7 1 2 42834 22521
0 22523 5 1 1 22522
0 22524 7 1 2 22517 22523
0 22525 5 1 1 22524
0 22526 7 1 2 47668 53121
0 22527 7 2 2 22525 22526
0 22528 7 1 2 58197 68611
0 22529 5 1 1 22528
0 22530 7 1 2 22507 22529
0 22531 5 1 1 22530
0 22532 7 1 2 42562 22531
0 22533 5 1 1 22532
0 22534 7 2 2 53775 64598
0 22535 7 1 2 52969 68613
0 22536 7 1 2 67997 22535
0 22537 5 1 1 22536
0 22538 7 1 2 44918 22537
0 22539 7 1 2 22533 22538
0 22540 5 1 1 22539
0 22541 7 1 2 44795 22540
0 22542 7 1 2 22490 22541
0 22543 5 1 1 22542
0 22544 7 1 2 22386 22543
0 22545 5 1 1 22544
0 22546 7 1 2 48008 22545
0 22547 5 1 1 22546
0 22548 7 3 2 43469 43925
0 22549 7 1 2 54637 68615
0 22550 7 2 2 65584 22549
0 22551 7 3 2 42031 61344
0 22552 7 1 2 51388 61567
0 22553 7 1 2 68620 22552
0 22554 7 1 2 68618 22553
0 22555 5 1 1 22554
0 22556 7 1 2 22547 22555
0 22557 5 2 1 22556
0 22558 7 1 2 45836 68623
0 22559 5 1 1 22558
0 22560 7 1 2 1792 66772
0 22561 5 2 1 22560
0 22562 7 3 2 42563 68625
0 22563 5 1 1 68627
0 22564 7 1 2 54081 68545
0 22565 5 1 1 22564
0 22566 7 1 2 22563 22565
0 22567 5 1 1 22566
0 22568 7 1 2 68564 22567
0 22569 5 2 1 22568
0 22570 7 3 2 52680 53806
0 22571 5 1 1 68632
0 22572 7 1 2 42564 68633
0 22573 5 1 1 22572
0 22574 7 2 2 46041 54611
0 22575 5 1 1 68635
0 22576 7 1 2 851 22575
0 22577 5 2 1 22576
0 22578 7 1 2 54244 68637
0 22579 5 1 1 22578
0 22580 7 1 2 22573 22579
0 22581 5 1 1 22580
0 22582 7 1 2 44796 22581
0 22583 5 1 1 22582
0 22584 7 8 2 46269 48126
0 22585 7 3 2 53137 58822
0 22586 7 2 2 68639 68647
0 22587 5 2 1 68650
0 22588 7 1 2 46042 68651
0 22589 5 1 1 22588
0 22590 7 1 2 22583 22589
0 22591 5 1 1 22590
0 22592 7 1 2 52225 22591
0 22593 5 1 1 22592
0 22594 7 1 2 68630 22593
0 22595 5 1 1 22594
0 22596 7 1 2 59914 65693
0 22597 7 1 2 22595 22596
0 22598 5 1 1 22597
0 22599 7 1 2 22559 22598
0 22600 5 1 1 22599
0 22601 7 1 2 42205 22600
0 22602 5 1 1 22601
0 22603 7 4 2 54360 56094
0 22604 7 2 2 59016 64460
0 22605 7 1 2 59679 68616
0 22606 7 1 2 54356 22605
0 22607 7 1 2 68658 22606
0 22608 7 1 2 68654 22607
0 22609 5 1 1 22608
0 22610 7 1 2 22602 22609
0 22611 5 1 1 22610
0 22612 7 1 2 67009 22611
0 22613 5 1 1 22612
0 22614 7 1 2 67089 68568
0 22615 5 1 1 22614
0 22616 7 2 2 66189 68332
0 22617 7 1 2 68574 68660
0 22618 5 1 1 22617
0 22619 7 1 2 66917 68572
0 22620 5 1 1 22619
0 22621 7 1 2 22618 22620
0 22622 5 1 1 22621
0 22623 7 1 2 45092 22622
0 22624 5 1 1 22623
0 22625 7 1 2 50250 51344
0 22626 5 1 1 22625
0 22627 7 1 2 22435 22626
0 22628 5 1 1 22627
0 22629 7 1 2 66918 22628
0 22630 5 1 1 22629
0 22631 7 1 2 63260 68170
0 22632 5 1 1 22631
0 22633 7 1 2 48814 59744
0 22634 7 1 2 66909 22633
0 22635 5 1 1 22634
0 22636 7 1 2 22632 22635
0 22637 5 1 1 22636
0 22638 7 1 2 49993 22637
0 22639 5 1 1 22638
0 22640 7 1 2 22630 22639
0 22641 5 1 1 22640
0 22642 7 1 2 47297 22641
0 22643 5 1 1 22642
0 22644 7 1 2 60151 68171
0 22645 5 1 1 22644
0 22646 7 1 2 22643 22645
0 22647 5 1 1 22646
0 22648 7 1 2 46270 22647
0 22649 5 1 1 22648
0 22650 7 1 2 22624 22649
0 22651 5 1 1 22650
0 22652 7 1 2 42565 22651
0 22653 5 1 1 22652
0 22654 7 1 2 65124 68172
0 22655 5 1 1 22654
0 22656 7 1 2 47669 67748
0 22657 7 1 2 67142 22656
0 22658 7 1 2 68583 22657
0 22659 5 1 1 22658
0 22660 7 1 2 22655 22659
0 22661 5 1 1 22660
0 22662 7 1 2 42835 22661
0 22663 5 1 1 22662
0 22664 7 1 2 68173 68589
0 22665 5 1 1 22664
0 22666 7 1 2 22663 22665
0 22667 5 1 1 22666
0 22668 7 1 2 46043 22667
0 22669 5 1 1 22668
0 22670 7 3 2 66470 66061
0 22671 7 1 2 55639 68662
0 22672 7 1 2 68597 22671
0 22673 5 1 1 22672
0 22674 7 1 2 22669 22673
0 22675 5 1 1 22674
0 22676 7 1 2 44071 22675
0 22677 5 1 1 22676
0 22678 7 1 2 67127 68601
0 22679 5 1 1 22678
0 22680 7 1 2 22677 22679
0 22681 5 1 1 22680
0 22682 7 1 2 49994 22681
0 22683 5 1 1 22682
0 22684 7 1 2 48260 22683
0 22685 7 1 2 22653 22684
0 22686 5 1 1 22685
0 22687 7 1 2 68603 68661
0 22688 5 1 1 22687
0 22689 7 1 2 66910 68605
0 22690 5 1 1 22689
0 22691 7 1 2 22688 22690
0 22692 5 1 1 22691
0 22693 7 1 2 44234 22692
0 22694 5 1 1 22693
0 22695 7 1 2 66911 68612
0 22696 5 1 1 22695
0 22697 7 1 2 22694 22696
0 22698 5 1 1 22697
0 22699 7 1 2 42566 22698
0 22700 5 1 1 22699
0 22701 7 1 2 65063 67085
0 22702 7 3 2 59603 66062
0 22703 7 1 2 68614 68665
0 22704 7 1 2 22701 22703
0 22705 5 1 1 22704
0 22706 7 1 2 44919 22705
0 22707 7 1 2 22700 22706
0 22708 5 1 1 22707
0 22709 7 1 2 44797 22708
0 22710 7 1 2 22686 22709
0 22711 5 1 1 22710
0 22712 7 1 2 22615 22711
0 22713 5 1 1 22712
0 22714 7 1 2 68522 22713
0 22715 5 1 1 22714
0 22716 7 2 2 49585 52562
0 22717 7 2 2 51980 68668
0 22718 7 4 2 42032 65541
0 22719 7 1 2 53542 59330
0 22720 7 1 2 63156 22719
0 22721 7 1 2 68672 22720
0 22722 7 1 2 68670 22721
0 22723 5 1 1 22722
0 22724 7 1 2 50224 58599
0 22725 5 1 1 22724
0 22726 7 1 2 43107 65410
0 22727 5 1 1 22726
0 22728 7 1 2 22725 22727
0 22729 5 1 1 22728
0 22730 7 1 2 46271 22729
0 22731 5 1 1 22730
0 22732 7 2 2 49287 55525
0 22733 7 1 2 50225 68676
0 22734 5 1 1 22733
0 22735 7 1 2 22731 22734
0 22736 5 1 1 22735
0 22737 7 1 2 42567 22736
0 22738 5 1 1 22737
0 22739 7 5 2 50947 54388
0 22740 5 1 1 68678
0 22741 7 2 2 50558 53855
0 22742 5 2 1 68683
0 22743 7 1 2 22740 68685
0 22744 5 1 1 22743
0 22745 7 1 2 44235 68584
0 22746 7 1 2 22744 22745
0 22747 5 1 1 22746
0 22748 7 1 2 22738 22747
0 22749 5 1 1 22748
0 22750 7 1 2 43324 22749
0 22751 5 1 1 22750
0 22752 7 1 2 62883 65674
0 22753 5 1 1 22752
0 22754 7 1 2 68570 22753
0 22755 5 1 1 22754
0 22756 7 1 2 68592 22755
0 22757 5 1 1 22756
0 22758 7 1 2 52047 68579
0 22759 5 1 1 22758
0 22760 7 1 2 22757 22759
0 22761 5 1 1 22760
0 22762 7 1 2 42568 22761
0 22763 5 1 1 22762
0 22764 7 1 2 22751 22763
0 22765 5 1 1 22764
0 22766 7 1 2 48261 22765
0 22767 5 1 1 22766
0 22768 7 1 2 50852 63591
0 22769 5 1 1 22768
0 22770 7 1 2 61915 63944
0 22771 5 1 1 22770
0 22772 7 1 2 22769 22771
0 22773 5 1 1 22772
0 22774 7 1 2 48815 22773
0 22775 5 1 1 22774
0 22776 7 1 2 42836 57730
0 22777 5 1 1 22776
0 22778 7 1 2 49697 56216
0 22779 5 5 1 22778
0 22780 7 1 2 22777 68687
0 22781 7 1 2 22775 22780
0 22782 5 1 1 22781
0 22783 7 1 2 57397 60087
0 22784 7 1 2 22782 22783
0 22785 5 1 1 22784
0 22786 7 1 2 22767 22785
0 22787 5 1 1 22786
0 22788 7 1 2 64501 66724
0 22789 7 1 2 22787 22788
0 22790 5 1 1 22789
0 22791 7 1 2 22723 22790
0 22792 5 1 1 22791
0 22793 7 1 2 67044 22792
0 22794 5 1 1 22793
0 22795 7 2 2 56513 66375
0 22796 7 1 2 54218 68692
0 22797 7 2 2 68655 22796
0 22798 7 5 2 45598 65542
0 22799 7 1 2 62043 62720
0 22800 7 1 2 68696 22799
0 22801 7 1 2 68694 22800
0 22802 5 1 1 22801
0 22803 7 1 2 22794 22802
0 22804 7 1 2 22715 22803
0 22805 5 1 1 22804
0 22806 7 1 2 48009 22805
0 22807 5 1 1 22806
0 22808 7 3 2 46044 51250
0 22809 5 1 1 68701
0 22810 7 2 2 42569 52160
0 22811 5 1 1 68704
0 22812 7 1 2 22809 22811
0 22813 5 5 1 22812
0 22814 7 1 2 52681 65040
0 22815 7 1 2 68706 22814
0 22816 5 1 1 22815
0 22817 7 1 2 68631 22816
0 22818 5 1 1 22817
0 22819 7 1 2 42311 22818
0 22820 5 1 1 22819
0 22821 7 1 2 60111 64645
0 22822 5 1 1 22821
0 22823 7 1 2 50206 53122
0 22824 7 1 2 67950 22823
0 22825 5 1 1 22824
0 22826 7 1 2 22822 22825
0 22827 5 1 1 22826
0 22828 7 1 2 42570 22827
0 22829 5 1 1 22828
0 22830 7 1 2 42312 58096
0 22831 7 1 2 68636 22830
0 22832 5 1 1 22831
0 22833 7 1 2 22829 22832
0 22834 5 1 1 22833
0 22835 7 1 2 54219 62412
0 22836 7 1 2 22834 22835
0 22837 5 1 1 22836
0 22838 7 1 2 22820 22837
0 22839 5 1 1 22838
0 22840 7 1 2 59017 66183
0 22841 7 2 2 63191 22840
0 22842 7 1 2 68066 68711
0 22843 7 1 2 22839 22842
0 22844 5 1 1 22843
0 22845 7 1 2 44462 22844
0 22846 7 1 2 22807 22845
0 22847 7 1 2 22613 22846
0 22848 5 1 1 22847
0 22849 7 7 2 52619 58237
0 22850 5 1 1 68713
0 22851 7 2 2 50948 68714
0 22852 5 1 1 68720
0 22853 7 1 2 58621 22852
0 22854 5 1 1 22853
0 22855 7 1 2 45259 22854
0 22856 5 1 1 22855
0 22857 7 1 2 51066 67242
0 22858 5 1 1 22857
0 22859 7 1 2 22856 22858
0 22860 5 1 1 22859
0 22861 7 1 2 50853 22860
0 22862 5 1 1 22861
0 22863 7 1 2 49431 50193
0 22864 5 1 1 22863
0 22865 7 1 2 52620 54297
0 22866 5 1 1 22865
0 22867 7 1 2 22864 22866
0 22868 5 1 1 22867
0 22869 7 1 2 58238 22868
0 22870 5 1 1 22869
0 22871 7 5 2 44920 53468
0 22872 5 1 1 68722
0 22873 7 1 2 65103 68723
0 22874 5 1 1 22873
0 22875 7 1 2 22870 22874
0 22876 5 1 1 22875
0 22877 7 1 2 50949 22876
0 22878 5 1 1 22877
0 22879 7 1 2 48977 51267
0 22880 7 1 2 65564 22879
0 22881 5 1 1 22880
0 22882 7 1 2 22878 22881
0 22883 7 1 2 22862 22882
0 22884 5 1 1 22883
0 22885 7 1 2 42837 22884
0 22886 5 1 1 22885
0 22887 7 1 2 43108 58489
0 22888 5 1 1 22887
0 22889 7 1 2 49288 50854
0 22890 7 1 2 53856 22889
0 22891 5 1 1 22890
0 22892 7 1 2 22888 22891
0 22893 5 1 1 22892
0 22894 7 1 2 45260 22893
0 22895 5 1 1 22894
0 22896 7 3 2 44072 48978
0 22897 5 3 1 68727
0 22898 7 1 2 56469 68728
0 22899 5 1 1 22898
0 22900 7 3 2 42571 54970
0 22901 7 1 2 62884 68733
0 22902 5 1 1 22901
0 22903 7 1 2 22899 22902
0 22904 5 1 1 22903
0 22905 7 1 2 50779 22904
0 22906 5 1 1 22905
0 22907 7 1 2 22895 22906
0 22908 5 1 1 22907
0 22909 7 1 2 51268 22908
0 22910 5 1 1 22909
0 22911 7 1 2 22886 22910
0 22912 5 1 1 22911
0 22913 7 2 2 44798 22912
0 22914 5 1 1 68736
0 22915 7 3 2 52184 62466
0 22916 5 1 1 68738
0 22917 7 2 2 46506 68739
0 22918 5 1 1 68741
0 22919 7 1 2 53323 22918
0 22920 5 1 1 22919
0 22921 7 1 2 47430 22920
0 22922 5 1 1 22921
0 22923 7 2 2 45261 56890
0 22924 5 1 1 68743
0 22925 7 1 2 61828 22924
0 22926 5 1 1 22925
0 22927 7 1 2 46507 22926
0 22928 5 1 1 22927
0 22929 7 1 2 45461 53873
0 22930 5 1 1 22929
0 22931 7 1 2 22928 22930
0 22932 5 1 1 22931
0 22933 7 1 2 46698 22932
0 22934 5 1 1 22933
0 22935 7 2 2 45262 61820
0 22936 5 1 1 68745
0 22937 7 1 2 22934 22936
0 22938 7 1 2 22922 22937
0 22939 5 1 1 22938
0 22940 7 1 2 48448 22939
0 22941 5 1 1 22940
0 22942 7 2 2 53425 56656
0 22943 5 1 1 68747
0 22944 7 1 2 45093 68748
0 22945 5 1 1 22944
0 22946 7 1 2 49621 53363
0 22947 5 2 1 22946
0 22948 7 1 2 53446 68749
0 22949 5 1 1 22948
0 22950 7 1 2 61821 22949
0 22951 5 1 1 22950
0 22952 7 1 2 42838 56854
0 22953 5 1 1 22952
0 22954 7 3 2 43109 50226
0 22955 5 1 1 68751
0 22956 7 1 2 50855 68752
0 22957 5 1 1 22956
0 22958 7 2 2 22953 22957
0 22959 7 1 2 22951 68754
0 22960 5 1 1 22959
0 22961 7 1 2 47431 22960
0 22962 5 1 1 22961
0 22963 7 1 2 22945 22962
0 22964 7 1 2 22941 22963
0 22965 5 1 1 22964
0 22966 7 1 2 47298 22965
0 22967 5 1 1 22966
0 22968 7 1 2 54697 68742
0 22969 5 1 1 22968
0 22970 7 1 2 56855 61959
0 22971 5 1 1 22970
0 22972 7 1 2 22969 22971
0 22973 5 1 1 22972
0 22974 7 1 2 46272 22973
0 22975 5 1 1 22974
0 22976 7 2 2 48965 52670
0 22977 7 1 2 54329 68756
0 22978 5 1 1 22977
0 22979 7 1 2 22975 22978
0 22980 7 1 2 22967 22979
0 22981 5 1 1 22980
0 22982 7 1 2 44921 22981
0 22983 5 1 1 22982
0 22984 7 1 2 43325 52732
0 22985 5 1 1 22984
0 22986 7 1 2 53064 22985
0 22987 5 4 1 22986
0 22988 7 1 2 54035 68758
0 22989 5 1 1 22988
0 22990 7 1 2 54698 67682
0 22991 5 1 1 22990
0 22992 7 1 2 22989 22991
0 22993 5 1 1 22992
0 22994 7 1 2 44922 22993
0 22995 5 1 1 22994
0 22996 7 1 2 45094 54918
0 22997 7 1 2 62333 22996
0 22998 5 1 1 22997
0 22999 7 1 2 22995 22998
0 23000 5 1 1 22999
0 23001 7 1 2 51432 23000
0 23002 5 1 1 23001
0 23003 7 1 2 45462 52074
0 23004 7 2 2 67729 23003
0 23005 5 1 1 68762
0 23006 7 1 2 45095 68763
0 23007 5 1 1 23006
0 23008 7 1 2 23002 23007
0 23009 7 1 2 22983 23008
0 23010 5 1 1 23009
0 23011 7 1 2 46045 23010
0 23012 5 1 1 23011
0 23013 7 2 2 54971 58497
0 23014 7 1 2 51433 57279
0 23015 7 2 2 68764 23014
0 23016 5 1 1 68766
0 23017 7 1 2 45096 68767
0 23018 5 1 1 23017
0 23019 7 1 2 23012 23018
0 23020 5 1 1 23019
0 23021 7 1 2 48127 23020
0 23022 5 1 1 23021
0 23023 7 1 2 22914 23022
0 23024 5 2 1 23023
0 23025 7 3 2 44669 68768
0 23026 7 1 2 59018 68770
0 23027 5 1 1 23026
0 23028 7 2 2 53151 56476
0 23029 7 1 2 45599 56038
0 23030 7 1 2 53535 23029
0 23031 7 1 2 68773 23030
0 23032 5 1 1 23031
0 23033 7 1 2 23027 23032
0 23034 5 1 1 23033
0 23035 7 1 2 67045 23034
0 23036 5 1 1 23035
0 23037 7 4 2 54782 67010
0 23038 7 5 2 42206 44670
0 23039 5 1 1 68779
0 23040 7 1 2 68769 68780
0 23041 5 1 1 23040
0 23042 7 2 2 52406 56477
0 23043 7 1 2 45756 62366
0 23044 7 1 2 65278 23043
0 23045 7 1 2 68784 23044
0 23046 5 1 1 23045
0 23047 7 1 2 23041 23046
0 23048 5 1 1 23047
0 23049 7 1 2 68775 23048
0 23050 5 1 1 23049
0 23051 7 1 2 54312 56039
0 23052 7 1 2 66629 66394
0 23053 7 1 2 67856 23052
0 23054 7 1 2 23051 23053
0 23055 7 2 2 51345 63312
0 23056 7 1 2 68656 68786
0 23057 7 1 2 23054 23056
0 23058 5 1 1 23057
0 23059 7 1 2 61269 67090
0 23060 7 1 2 68771 23059
0 23061 5 1 1 23060
0 23062 7 1 2 23058 23061
0 23063 7 1 2 23050 23062
0 23064 7 1 2 23036 23063
0 23065 5 1 1 23064
0 23066 7 1 2 44334 23065
0 23067 5 1 1 23066
0 23068 7 1 2 49001 64332
0 23069 5 1 1 23068
0 23070 7 1 2 46046 57142
0 23071 7 1 2 61687 23070
0 23072 5 1 1 23071
0 23073 7 1 2 46273 23072
0 23074 7 1 2 23069 23073
0 23075 5 1 1 23074
0 23076 7 2 2 46047 57386
0 23077 5 1 1 68788
0 23078 7 1 2 64327 68789
0 23079 5 1 1 23078
0 23080 7 1 2 42839 23079
0 23081 5 1 1 23080
0 23082 7 1 2 48449 23081
0 23083 7 1 2 23075 23082
0 23084 5 1 1 23083
0 23085 7 1 2 49424 54168
0 23086 7 1 2 65515 23085
0 23087 5 1 1 23086
0 23088 7 1 2 23084 23087
0 23089 5 1 1 23088
0 23090 7 1 2 52161 23089
0 23091 5 1 1 23090
0 23092 7 1 2 52752 54396
0 23093 7 1 2 52289 23092
0 23094 5 1 1 23093
0 23095 7 1 2 23091 23094
0 23096 5 1 1 23095
0 23097 7 1 2 61280 61734
0 23098 7 2 2 23096 23097
0 23099 7 1 2 67143 68372
0 23100 7 1 2 68790 23099
0 23101 5 1 1 23100
0 23102 7 1 2 23067 23101
0 23103 5 1 1 23102
0 23104 7 1 2 42313 23103
0 23105 5 1 1 23104
0 23106 7 4 2 54313 66752
0 23107 7 1 2 65503 68792
0 23108 5 1 1 23107
0 23109 7 1 2 65401 23108
0 23110 5 1 1 23109
0 23111 7 1 2 49169 23110
0 23112 5 1 1 23111
0 23113 7 1 2 15145 23112
0 23114 5 1 1 23113
0 23115 7 1 2 46699 23114
0 23116 5 1 1 23115
0 23117 7 2 2 64352 65089
0 23118 5 1 1 68796
0 23119 7 2 2 43326 68797
0 23120 5 1 1 68798
0 23121 7 1 2 45097 68799
0 23122 5 1 1 23121
0 23123 7 1 2 23116 23122
0 23124 5 1 1 23123
0 23125 7 1 2 58239 23124
0 23126 5 1 1 23125
0 23127 7 2 2 61526 68707
0 23128 7 1 2 65289 68800
0 23129 5 1 1 23128
0 23130 7 2 2 46048 53536
0 23131 7 1 2 54407 68724
0 23132 7 1 2 68802 23131
0 23133 5 1 1 23132
0 23134 7 1 2 23129 23133
0 23135 5 1 1 23134
0 23136 7 1 2 48623 23135
0 23137 5 1 1 23136
0 23138 7 1 2 23126 23137
0 23139 5 1 1 23138
0 23140 7 1 2 48010 23139
0 23141 5 1 1 23140
0 23142 7 2 2 43327 52962
0 23143 7 2 2 54400 68804
0 23144 7 1 2 49869 65070
0 23145 7 2 2 68806 23144
0 23146 5 1 1 68808
0 23147 7 1 2 48816 68809
0 23148 5 1 1 23147
0 23149 7 1 2 23141 23148
0 23150 5 2 1 23149
0 23151 7 1 2 42207 67011
0 23152 5 1 1 23151
0 23153 7 2 2 67120 66941
0 23154 5 1 1 68812
0 23155 7 1 2 23152 23154
0 23156 5 6 1 23155
0 23157 7 1 2 54783 68814
0 23158 5 2 1 23157
0 23159 7 1 2 59019 66370
0 23160 7 1 2 67419 23159
0 23161 5 1 1 23160
0 23162 7 1 2 68820 23161
0 23163 5 2 1 23162
0 23164 7 5 2 44335 68822
0 23165 7 1 2 45837 68824
0 23166 7 1 2 68810 23165
0 23167 5 1 1 23166
0 23168 7 1 2 47778 23167
0 23169 7 1 2 23105 23168
0 23170 5 1 1 23169
0 23171 7 1 2 22848 23170
0 23172 5 1 1 23171
0 23173 7 1 2 47907 23172
0 23174 5 1 1 23173
0 23175 7 2 2 44923 52299
0 23176 5 1 1 68829
0 23177 7 1 2 56780 68046
0 23178 5 1 1 23177
0 23179 7 1 2 23176 23178
0 23180 5 1 1 23179
0 23181 7 1 2 42840 23180
0 23182 5 1 1 23181
0 23183 7 1 2 52621 68830
0 23184 5 1 1 23183
0 23185 7 2 2 49656 52320
0 23186 5 1 1 68831
0 23187 7 1 2 23184 23186
0 23188 7 1 2 23182 23187
0 23189 5 2 1 23188
0 23190 7 1 2 55906 68833
0 23191 5 1 1 23190
0 23192 7 2 2 50856 52622
0 23193 7 1 2 55463 66601
0 23194 7 1 2 68835 23193
0 23195 5 1 1 23194
0 23196 7 1 2 23191 23195
0 23197 5 1 1 23196
0 23198 7 1 2 45263 23197
0 23199 5 1 1 23198
0 23200 7 2 2 48450 52063
0 23201 5 1 1 68837
0 23202 7 1 2 55907 68838
0 23203 5 1 1 23202
0 23204 7 1 2 2203 65505
0 23205 5 2 1 23204
0 23206 7 1 2 55620 58900
0 23207 7 1 2 68839 23206
0 23208 5 1 1 23207
0 23209 7 1 2 23203 23208
0 23210 5 1 1 23209
0 23211 7 1 2 46700 23210
0 23212 5 1 1 23211
0 23213 7 1 2 49425 56728
0 23214 7 1 2 60425 66448
0 23215 7 1 2 23213 23214
0 23216 5 1 1 23215
0 23217 7 1 2 23212 23216
0 23218 5 1 1 23217
0 23219 7 1 2 44924 23218
0 23220 5 1 1 23219
0 23221 7 1 2 23199 23220
0 23222 5 1 1 23221
0 23223 7 1 2 61170 23222
0 23224 5 1 1 23223
0 23225 7 1 2 49109 55908
0 23226 5 1 1 23225
0 23227 7 1 2 60426 64195
0 23228 5 1 1 23227
0 23229 7 1 2 23226 23228
0 23230 5 1 1 23229
0 23231 7 2 2 53165 56086
0 23232 7 1 2 67219 68841
0 23233 7 1 2 23230 23232
0 23234 5 1 1 23233
0 23235 7 1 2 23224 23234
0 23236 5 1 1 23235
0 23237 7 1 2 50950 23236
0 23238 5 1 1 23237
0 23239 7 1 2 46701 68626
0 23240 7 1 2 53823 23239
0 23241 5 1 1 23240
0 23242 7 4 2 48817 53138
0 23243 7 1 2 52162 68843
0 23244 7 1 2 64587 23243
0 23245 5 1 1 23244
0 23246 7 1 2 23241 23245
0 23247 5 1 1 23246
0 23248 7 1 2 55909 23247
0 23249 5 1 1 23248
0 23250 7 1 2 51434 66769
0 23251 5 1 1 23250
0 23252 7 1 2 57099 60216
0 23253 5 6 1 23252
0 23254 7 2 2 48451 68847
0 23255 7 1 2 52163 68853
0 23256 5 1 1 23255
0 23257 7 1 2 23251 23256
0 23258 5 1 1 23257
0 23259 7 4 2 47432 47779
0 23260 7 1 2 60024 68855
0 23261 7 1 2 23258 23260
0 23262 5 1 1 23261
0 23263 7 1 2 23249 23262
0 23264 5 1 1 23263
0 23265 7 1 2 61415 23264
0 23266 5 1 1 23265
0 23267 7 1 2 23238 23266
0 23268 5 1 1 23267
0 23269 7 1 2 42572 23268
0 23270 5 1 1 23269
0 23271 7 3 2 48452 51435
0 23272 7 1 2 46702 68859
0 23273 5 1 1 23272
0 23274 7 1 2 53405 23273
0 23275 5 2 1 23274
0 23276 7 1 2 44925 68862
0 23277 5 1 1 23276
0 23278 7 3 2 45098 51436
0 23279 5 1 1 68864
0 23280 7 2 2 54726 68865
0 23281 5 1 1 68867
0 23282 7 1 2 46703 68868
0 23283 5 1 1 23282
0 23284 7 1 2 23277 23283
0 23285 5 1 1 23284
0 23286 7 1 2 47433 23285
0 23287 5 1 1 23286
0 23288 7 1 2 44926 65290
0 23289 5 1 1 23288
0 23290 7 1 2 47299 68832
0 23291 5 2 1 23290
0 23292 7 1 2 23289 68869
0 23293 5 1 1 23292
0 23294 7 1 2 45264 23293
0 23295 5 1 1 23294
0 23296 7 1 2 23287 23295
0 23297 5 1 1 23296
0 23298 7 1 2 55910 23297
0 23299 5 1 1 23298
0 23300 7 1 2 52480 57970
0 23301 5 1 1 23300
0 23302 7 1 2 52583 56300
0 23303 5 1 1 23302
0 23304 7 1 2 23301 23303
0 23305 5 1 1 23304
0 23306 7 1 2 49496 23305
0 23307 5 1 1 23306
0 23308 7 1 2 52481 60212
0 23309 5 1 1 23308
0 23310 7 1 2 23281 23309
0 23311 5 1 1 23310
0 23312 7 1 2 55621 23311
0 23313 5 1 1 23312
0 23314 7 1 2 23307 23313
0 23315 5 1 1 23314
0 23316 7 1 2 49289 23315
0 23317 5 1 1 23316
0 23318 7 1 2 23299 23317
0 23319 5 1 1 23318
0 23320 7 1 2 68640 23319
0 23321 5 1 1 23320
0 23322 7 1 2 7053 65109
0 23323 5 1 1 23322
0 23324 7 1 2 53015 23323
0 23325 5 1 1 23324
0 23326 7 1 2 48262 23325
0 23327 5 1 1 23326
0 23328 7 1 2 57398 60127
0 23329 5 1 1 23328
0 23330 7 1 2 23327 23329
0 23331 5 1 1 23330
0 23332 7 2 2 43110 55622
0 23333 5 1 1 68871
0 23334 7 1 2 55927 23333
0 23335 5 1 1 23334
0 23336 7 1 2 48624 23335
0 23337 7 1 2 23331 23336
0 23338 5 1 1 23337
0 23339 7 1 2 60217 64140
0 23340 5 1 1 23339
0 23341 7 3 2 48263 52623
0 23342 7 1 2 68873 68872
0 23343 7 1 2 23340 23342
0 23344 5 1 1 23343
0 23345 7 1 2 23338 23344
0 23346 5 1 1 23345
0 23347 7 1 2 44799 54314
0 23348 7 1 2 23346 23347
0 23349 5 1 1 23348
0 23350 7 1 2 23321 23349
0 23351 5 1 1 23350
0 23352 7 1 2 61875 23351
0 23353 5 1 1 23352
0 23354 7 1 2 23270 23353
0 23355 5 1 1 23354
0 23356 7 3 2 66184 68093
0 23357 7 3 2 63734 68876
0 23358 7 1 2 23355 68879
0 23359 5 1 1 23358
0 23360 7 1 2 46508 57413
0 23361 5 1 1 23360
0 23362 7 1 2 42573 23361
0 23363 5 1 1 23362
0 23364 7 1 2 54666 67362
0 23365 7 2 2 67937 23364
0 23366 7 1 2 23363 68882
0 23367 5 1 1 23366
0 23368 7 1 2 55928 17868
0 23369 5 2 1 23368
0 23370 7 1 2 49586 60899
0 23371 7 1 2 50715 23370
0 23372 7 1 2 68884 23371
0 23373 7 1 2 67012 23372
0 23374 5 1 1 23373
0 23375 7 1 2 23367 23374
0 23376 5 1 1 23375
0 23377 7 1 2 48625 23376
0 23378 5 1 1 23377
0 23379 7 1 2 64528 68243
0 23380 7 1 2 63451 23379
0 23381 7 1 2 67370 23380
0 23382 5 1 1 23381
0 23383 7 1 2 23378 23382
0 23384 5 1 1 23383
0 23385 7 1 2 44073 23384
0 23386 5 1 1 23385
0 23387 7 1 2 42841 65562
0 23388 5 1 1 23387
0 23389 7 1 2 57334 63681
0 23390 5 5 1 23389
0 23391 7 1 2 68746 68886
0 23392 5 1 1 23391
0 23393 7 1 2 50559 56217
0 23394 5 1 1 23393
0 23395 7 1 2 64602 23394
0 23396 5 1 1 23395
0 23397 7 1 2 50857 23396
0 23398 5 1 1 23397
0 23399 7 1 2 23392 23398
0 23400 7 1 2 23388 23399
0 23401 5 1 1 23400
0 23402 7 1 2 68883 23401
0 23403 5 1 1 23402
0 23404 7 1 2 23386 23403
0 23405 5 1 1 23404
0 23406 7 1 2 42208 23405
0 23407 5 1 1 23406
0 23408 7 1 2 68877 68885
0 23409 5 1 1 23408
0 23410 7 6 2 66684 67040
0 23411 7 1 2 58063 68891
0 23412 5 1 1 23411
0 23413 7 1 2 23409 23412
0 23414 5 1 1 23413
0 23415 7 1 2 50716 58991
0 23416 7 1 2 62413 23415
0 23417 7 1 2 23414 23416
0 23418 5 1 1 23417
0 23419 7 1 2 23407 23418
0 23420 5 1 1 23419
0 23421 7 1 2 67243 23420
0 23422 5 1 1 23421
0 23423 7 1 2 57451 65365
0 23424 5 1 1 23423
0 23425 7 1 2 44800 57885
0 23426 7 1 2 53155 23425
0 23427 5 1 1 23426
0 23428 7 1 2 23424 23427
0 23429 5 1 1 23428
0 23430 7 1 2 42842 23429
0 23431 5 1 1 23430
0 23432 7 1 2 53016 65286
0 23433 5 1 1 23432
0 23434 7 1 2 49757 23433
0 23435 5 1 1 23434
0 23436 7 1 2 49380 57579
0 23437 5 2 1 23436
0 23438 7 1 2 23435 68897
0 23439 5 1 1 23438
0 23440 7 1 2 46274 23439
0 23441 5 1 1 23440
0 23442 7 2 2 14442 23441
0 23443 7 1 2 46704 68729
0 23444 5 1 1 23443
0 23445 7 1 2 65345 23444
0 23446 5 1 1 23445
0 23447 7 1 2 45099 23446
0 23448 5 1 1 23447
0 23449 7 1 2 61822 64588
0 23450 5 1 1 23449
0 23451 7 2 2 107 23450
0 23452 7 1 2 23448 68901
0 23453 5 1 1 23452
0 23454 7 1 2 47300 23453
0 23455 5 1 1 23454
0 23456 7 1 2 68899 23455
0 23457 5 1 1 23456
0 23458 7 1 2 55911 23457
0 23459 5 1 1 23458
0 23460 7 1 2 49048 65022
0 23461 5 1 1 23460
0 23462 7 1 2 49403 23461
0 23463 5 1 1 23462
0 23464 7 1 2 51004 23463
0 23465 5 1 1 23464
0 23466 7 1 2 49290 68860
0 23467 5 1 1 23466
0 23468 7 1 2 23465 23467
0 23469 5 3 1 23468
0 23470 7 1 2 62233 68903
0 23471 5 1 1 23470
0 23472 7 1 2 23459 23471
0 23473 5 1 1 23472
0 23474 7 1 2 48128 23473
0 23475 5 1 1 23474
0 23476 7 1 2 23431 23475
0 23477 5 1 1 23476
0 23478 7 1 2 46049 23477
0 23479 5 1 1 23478
0 23480 7 2 2 42574 51437
0 23481 7 1 2 68730 68906
0 23482 5 1 1 23481
0 23483 7 1 2 49491 51400
0 23484 7 1 2 55282 23483
0 23485 5 1 1 23484
0 23486 7 2 2 62353 23485
0 23487 5 1 1 68908
0 23488 7 1 2 23482 68909
0 23489 5 1 1 23488
0 23490 7 1 2 45100 23489
0 23491 5 1 1 23490
0 23492 7 1 2 51458 55251
0 23493 5 2 1 23492
0 23494 7 1 2 23491 68910
0 23495 5 1 1 23494
0 23496 7 1 2 46705 23495
0 23497 5 1 1 23496
0 23498 7 2 2 45265 65107
0 23499 5 1 1 68912
0 23500 7 1 2 45101 68913
0 23501 5 1 1 23500
0 23502 7 1 2 23497 23501
0 23503 5 1 1 23502
0 23504 7 1 2 57213 23503
0 23505 5 1 1 23504
0 23506 7 1 2 43926 49110
0 23507 5 1 1 23506
0 23508 7 1 2 21913 23507
0 23509 5 1 1 23508
0 23510 7 1 2 43328 23509
0 23511 5 1 1 23510
0 23512 7 1 2 49866 23511
0 23513 5 1 1 23512
0 23514 7 1 2 53426 23513
0 23515 5 1 1 23514
0 23516 7 1 2 49111 53166
0 23517 5 1 1 23516
0 23518 7 1 2 23201 23517
0 23519 5 1 1 23518
0 23520 7 1 2 50951 23519
0 23521 5 1 1 23520
0 23522 7 1 2 55686 23521
0 23523 7 1 2 23515 23522
0 23524 5 1 1 23523
0 23525 7 1 2 42575 23524
0 23526 5 1 1 23525
0 23527 7 1 2 56508 56340
0 23528 5 1 1 23527
0 23529 7 1 2 23526 23528
0 23530 5 1 1 23529
0 23531 7 1 2 44801 23530
0 23532 5 1 1 23531
0 23533 7 1 2 23505 23532
0 23534 5 1 1 23533
0 23535 7 1 2 55912 23534
0 23536 5 1 1 23535
0 23537 7 4 2 52624 68793
0 23538 5 1 1 68914
0 23539 7 1 2 52440 57214
0 23540 5 1 1 23539
0 23541 7 1 2 23538 23540
0 23542 5 1 1 23541
0 23543 7 1 2 49170 23542
0 23544 5 1 1 23543
0 23545 7 4 2 46275 52269
0 23546 7 1 2 52761 68918
0 23547 5 1 1 23546
0 23548 7 1 2 23118 23547
0 23549 5 1 1 23548
0 23550 7 1 2 45102 23549
0 23551 5 1 1 23550
0 23552 7 1 2 23544 23551
0 23553 5 1 1 23552
0 23554 7 1 2 42576 55623
0 23555 7 1 2 23553 23554
0 23556 5 1 1 23555
0 23557 7 1 2 23536 23556
0 23558 7 1 2 23479 23557
0 23559 5 1 1 23558
0 23560 7 1 2 44927 23559
0 23561 5 1 1 23560
0 23562 7 2 2 44463 68617
0 23563 7 1 2 52197 68922
0 23564 5 1 1 23563
0 23565 7 1 2 8408 64880
0 23566 5 1 1 23565
0 23567 7 1 2 57886 23566
0 23568 5 1 1 23567
0 23569 7 1 2 23564 23568
0 23570 5 1 1 23569
0 23571 7 1 2 44074 23570
0 23572 5 1 1 23571
0 23573 7 1 2 56643 68923
0 23574 5 1 1 23573
0 23575 7 1 2 23572 23574
0 23576 5 1 1 23575
0 23577 7 1 2 67705 23576
0 23578 5 1 1 23577
0 23579 7 2 2 53829 55624
0 23580 5 1 1 68924
0 23581 7 1 2 53824 57455
0 23582 5 1 1 23581
0 23583 7 1 2 23580 23582
0 23584 5 1 1 23583
0 23585 7 1 2 52584 68641
0 23586 7 1 2 23584 23585
0 23587 5 1 1 23586
0 23588 7 1 2 23578 23587
0 23589 5 1 1 23588
0 23590 7 1 2 46050 23589
0 23591 5 1 1 23590
0 23592 7 1 2 53857 53833
0 23593 5 1 1 23592
0 23594 7 1 2 54397 58457
0 23595 5 1 1 23594
0 23596 7 1 2 23593 23595
0 23597 5 1 1 23596
0 23598 7 1 2 55625 23597
0 23599 5 1 1 23598
0 23600 7 1 2 1418 56669
0 23601 5 1 1 23600
0 23602 7 1 2 1707 56671
0 23603 5 1 1 23602
0 23604 7 1 2 55913 23603
0 23605 7 1 2 23601 23604
0 23606 5 1 1 23605
0 23607 7 1 2 23599 23606
0 23608 5 1 1 23607
0 23609 7 1 2 48453 23608
0 23610 5 1 1 23609
0 23611 7 2 2 56874 67971
0 23612 7 1 2 62397 68926
0 23613 5 1 1 23612
0 23614 7 1 2 47301 58072
0 23615 5 1 1 23614
0 23616 7 1 2 23613 23615
0 23617 5 1 1 23616
0 23618 7 1 2 48626 23617
0 23619 5 1 1 23618
0 23620 7 1 2 57465 68744
0 23621 5 1 1 23620
0 23622 7 1 2 23619 23621
0 23623 5 1 1 23622
0 23624 7 1 2 42577 23623
0 23625 5 1 1 23624
0 23626 7 2 2 53167 55863
0 23627 7 1 2 52937 61951
0 23628 7 1 2 68928 23627
0 23629 5 1 1 23628
0 23630 7 1 2 23625 23629
0 23631 5 1 1 23630
0 23632 7 1 2 45103 23631
0 23633 5 1 1 23632
0 23634 7 1 2 51005 52384
0 23635 7 1 2 58498 23634
0 23636 7 1 2 68927 23635
0 23637 5 1 1 23636
0 23638 7 1 2 23633 23637
0 23639 7 1 2 23610 23638
0 23640 5 1 1 23639
0 23641 7 1 2 44802 23640
0 23642 5 1 1 23641
0 23643 7 1 2 23591 23642
0 23644 5 1 1 23643
0 23645 7 1 2 48264 23644
0 23646 5 1 1 23645
0 23647 7 1 2 23561 23646
0 23648 5 1 1 23647
0 23649 7 3 2 44671 52786
0 23650 7 1 2 66358 68930
0 23651 7 1 2 23648 23650
0 23652 5 1 1 23651
0 23653 7 1 2 23422 23652
0 23654 5 1 1 23653
0 23655 7 1 2 42314 23654
0 23656 5 1 1 23655
0 23657 7 1 2 23359 23656
0 23658 5 1 1 23657
0 23659 7 1 2 44336 23658
0 23660 5 1 1 23659
0 23661 7 6 2 48454 57110
0 23662 7 2 2 57082 68933
0 23663 5 1 1 68939
0 23664 7 1 2 65996 68940
0 23665 5 1 1 23664
0 23666 7 3 2 42315 53168
0 23667 7 1 2 56802 57136
0 23668 7 1 2 68941 23667
0 23669 5 1 1 23668
0 23670 7 1 2 23665 23669
0 23671 5 1 1 23670
0 23672 7 1 2 48265 23671
0 23673 5 1 1 23672
0 23674 7 4 2 44928 52385
0 23675 7 5 2 44672 64646
0 23676 5 2 1 68948
0 23677 7 1 2 44236 51981
0 23678 7 2 2 68949 23677
0 23679 7 1 2 68944 68955
0 23680 5 1 1 23679
0 23681 7 1 2 23673 23680
0 23682 5 1 1 23681
0 23683 7 1 2 46509 23682
0 23684 5 1 1 23683
0 23685 7 1 2 67785 68956
0 23686 5 1 1 23685
0 23687 7 1 2 23684 23686
0 23688 5 1 1 23687
0 23689 7 1 2 47434 23688
0 23690 5 1 1 23689
0 23691 7 1 2 52064 53012
0 23692 5 1 1 23691
0 23693 7 1 2 54182 57480
0 23694 5 1 1 23693
0 23695 7 1 2 23692 23694
0 23696 5 1 1 23695
0 23697 7 1 2 44929 23696
0 23698 5 1 1 23697
0 23699 7 1 2 68870 23698
0 23700 5 1 1 23699
0 23701 7 1 2 48627 23700
0 23702 5 1 1 23701
0 23703 7 4 2 44237 44930
0 23704 7 3 2 48455 68957
0 23705 7 2 2 53169 68961
0 23706 5 1 1 68964
0 23707 7 1 2 47302 68965
0 23708 5 1 1 23707
0 23709 7 1 2 23702 23708
0 23710 5 1 1 23709
0 23711 7 1 2 61388 63250
0 23712 7 1 2 23710 23711
0 23713 5 1 1 23712
0 23714 7 1 2 23690 23713
0 23715 5 1 1 23714
0 23716 7 1 2 55400 59157
0 23717 7 1 2 23715 23716
0 23718 5 1 1 23717
0 23719 7 1 2 53807 68904
0 23720 5 1 1 23719
0 23721 7 2 2 49171 52625
0 23722 5 2 1 68966
0 23723 7 1 2 64881 68968
0 23724 5 1 1 23723
0 23725 7 1 2 55937 23724
0 23726 5 1 1 23725
0 23727 7 1 2 23720 23726
0 23728 5 2 1 23727
0 23729 7 1 2 65694 68970
0 23730 5 1 1 23729
0 23731 7 1 2 44931 52626
0 23732 7 1 2 55130 23731
0 23733 5 1 1 23732
0 23734 7 3 2 46276 51269
0 23735 7 1 2 49291 68972
0 23736 5 1 1 23735
0 23737 7 1 2 23733 23736
0 23738 5 4 1 23737
0 23739 7 1 2 68848 68975
0 23740 5 1 1 23739
0 23741 7 1 2 50780 52627
0 23742 5 1 1 23741
0 23743 7 1 2 52261 23742
0 23744 5 1 1 23743
0 23745 7 1 2 54058 54245
0 23746 7 1 2 23744 23745
0 23747 5 1 1 23746
0 23748 7 1 2 23740 23747
0 23749 5 1 1 23748
0 23750 7 1 2 65904 23749
0 23751 5 1 1 23750
0 23752 7 1 2 23730 23751
0 23753 5 1 1 23752
0 23754 7 1 2 42578 23753
0 23755 5 1 1 23754
0 23756 7 1 2 65788 17149
0 23757 5 6 1 23756
0 23758 7 3 2 52386 68979
0 23759 7 1 2 54612 68985
0 23760 5 1 1 23759
0 23761 7 7 2 45838 61008
0 23762 7 2 2 52628 68988
0 23763 5 1 1 68995
0 23764 7 2 2 48266 68996
0 23765 5 1 1 68997
0 23766 7 1 2 23760 23765
0 23767 5 1 1 23766
0 23768 7 1 2 44238 23767
0 23769 5 1 1 23768
0 23770 7 1 2 50281 54299
0 23771 5 1 1 23770
0 23772 7 1 2 65905 23771
0 23773 5 1 1 23772
0 23774 7 1 2 66997 23773
0 23775 5 1 1 23774
0 23776 7 2 2 52629 23775
0 23777 5 1 1 68999
0 23778 7 1 2 48267 69000
0 23779 5 1 1 23778
0 23780 7 1 2 23769 23779
0 23781 5 1 1 23780
0 23782 7 1 2 68679 23781
0 23783 5 1 1 23782
0 23784 7 1 2 23755 23783
0 23785 5 1 1 23784
0 23786 7 1 2 61317 23785
0 23787 5 1 1 23786
0 23788 7 1 2 44803 23787
0 23789 7 1 2 23718 23788
0 23790 5 1 1 23789
0 23791 7 1 2 45757 67013
0 23792 5 1 1 23791
0 23793 7 1 2 20556 23792
0 23794 5 7 1 23793
0 23795 7 2 2 44673 49878
0 23796 7 1 2 68671 69008
0 23797 5 1 1 23796
0 23798 7 2 2 55186 68111
0 23799 7 1 2 51459 69010
0 23800 5 1 1 23799
0 23801 7 1 2 23797 23800
0 23802 5 1 1 23801
0 23803 7 1 2 43329 23802
0 23804 5 1 1 23803
0 23805 7 3 2 50919 55342
0 23806 7 1 2 52185 68112
0 23807 7 1 2 56657 23806
0 23808 7 1 2 69012 23807
0 23809 5 1 1 23808
0 23810 7 1 2 23804 23809
0 23811 5 1 1 23810
0 23812 7 1 2 48456 23811
0 23813 5 1 1 23812
0 23814 7 1 2 51438 54972
0 23815 7 2 2 52585 62066
0 23816 7 1 2 58240 69015
0 23817 7 1 2 23814 23816
0 23818 5 1 1 23817
0 23819 7 1 2 23813 23818
0 23820 5 1 1 23819
0 23821 7 1 2 45839 23820
0 23822 5 1 1 23821
0 23823 7 1 2 52493 58233
0 23824 5 1 1 23823
0 23825 7 1 2 22850 23824
0 23826 7 1 2 53834 23825
0 23827 5 1 1 23826
0 23828 7 1 2 49049 64599
0 23829 7 1 2 68648 23828
0 23830 5 1 1 23829
0 23831 7 1 2 23827 23830
0 23832 5 1 1 23831
0 23833 7 1 2 68396 23832
0 23834 5 1 1 23833
0 23835 7 1 2 23822 23834
0 23836 5 1 1 23835
0 23837 7 1 2 61318 23836
0 23838 5 1 1 23837
0 23839 7 2 2 52586 62461
0 23840 5 1 1 69017
0 23841 7 1 2 46051 68934
0 23842 5 1 1 23841
0 23843 7 1 2 23840 23842
0 23844 5 1 1 23843
0 23845 7 1 2 44932 23844
0 23846 5 1 1 23845
0 23847 7 4 2 46052 49816
0 23848 5 1 1 69019
0 23849 7 1 2 52587 69020
0 23850 5 1 1 23849
0 23851 7 1 2 23846 23850
0 23852 5 1 1 23851
0 23853 7 1 2 65997 23852
0 23854 5 1 1 23853
0 23855 7 2 2 66599 67827
0 23856 5 1 1 69023
0 23857 7 1 2 46053 69024
0 23858 5 1 1 23857
0 23859 7 1 2 23854 23858
0 23860 5 1 1 23859
0 23861 7 2 2 50331 59158
0 23862 7 1 2 68295 69025
0 23863 7 1 2 23860 23862
0 23864 5 1 1 23863
0 23865 7 1 2 48129 23864
0 23866 7 1 2 23838 23865
0 23867 5 1 1 23866
0 23868 7 1 2 69001 23867
0 23869 7 1 2 23790 23868
0 23870 5 1 1 23869
0 23871 7 1 2 42033 23870
0 23872 7 1 2 23660 23871
0 23873 5 1 1 23872
0 23874 7 1 2 65695 68905
0 23875 5 1 1 23874
0 23876 7 3 2 45840 47435
0 23877 7 2 2 62836 69027
0 23878 5 1 1 69030
0 23879 7 1 2 68854 69031
0 23880 5 1 1 23879
0 23881 7 1 2 23875 23880
0 23882 5 1 1 23881
0 23883 7 1 2 68708 23882
0 23884 5 1 1 23883
0 23885 7 4 2 44674 48966
0 23886 7 1 2 66461 69032
0 23887 5 1 1 23886
0 23888 7 1 2 46510 65998
0 23889 7 1 2 53814 23888
0 23890 5 1 1 23889
0 23891 7 1 2 23887 23890
0 23892 5 1 1 23891
0 23893 7 1 2 51006 58241
0 23894 7 1 2 65315 23893
0 23895 7 1 2 23892 23894
0 23896 5 1 1 23895
0 23897 7 1 2 23884 23896
0 23898 5 1 1 23897
0 23899 7 1 2 46277 23898
0 23900 5 1 1 23899
0 23901 7 1 2 45104 68986
0 23902 5 1 1 23901
0 23903 7 1 2 23763 23902
0 23904 5 1 1 23903
0 23905 7 1 2 44239 23904
0 23906 5 1 1 23905
0 23907 7 1 2 23777 23906
0 23908 5 1 1 23907
0 23909 7 1 2 58242 23908
0 23910 5 1 1 23909
0 23911 7 1 2 56636 68962
0 23912 7 1 2 68987 23911
0 23913 5 1 1 23912
0 23914 7 1 2 23910 23913
0 23915 5 1 1 23914
0 23916 7 1 2 44804 23915
0 23917 5 1 1 23916
0 23918 7 1 2 54626 60407
0 23919 7 1 2 64100 23918
0 23920 7 1 2 65059 23919
0 23921 5 1 1 23920
0 23922 7 1 2 23917 23921
0 23923 5 1 1 23922
0 23924 7 1 2 54246 23923
0 23925 5 1 1 23924
0 23926 7 1 2 23900 23925
0 23927 5 1 1 23926
0 23928 7 1 2 43545 23927
0 23929 5 1 1 23928
0 23930 7 1 2 53527 66647
0 23931 7 1 2 65667 23930
0 23932 7 1 2 68774 23931
0 23933 5 1 1 23932
0 23934 7 1 2 23929 23933
0 23935 5 1 1 23934
0 23936 7 1 2 66190 23935
0 23937 5 1 1 23936
0 23938 7 1 2 45917 66630
0 23939 7 1 2 65064 23938
0 23940 7 3 2 43546 66139
0 23941 7 1 2 65668 69036
0 23942 7 1 2 23939 23941
0 23943 7 1 2 68657 23942
0 23944 5 1 1 23943
0 23945 7 1 2 23937 23944
0 23946 5 1 1 23945
0 23947 7 1 2 42209 23946
0 23948 5 1 1 23947
0 23949 7 1 2 62367 66631
0 23950 7 1 2 65526 23949
0 23951 7 1 2 68695 23950
0 23952 5 1 1 23951
0 23953 7 1 2 23948 23952
0 23954 5 1 1 23953
0 23955 7 1 2 61319 23954
0 23956 5 1 1 23955
0 23957 7 1 2 53776 66753
0 23958 7 1 2 58535 23957
0 23959 5 1 1 23958
0 23960 7 1 2 50145 53957
0 23961 7 1 2 56658 23960
0 23962 5 1 1 23961
0 23963 7 1 2 23959 23962
0 23964 5 1 1 23963
0 23965 7 1 2 47303 23964
0 23966 5 1 1 23965
0 23967 7 1 2 53017 56794
0 23968 5 1 1 23967
0 23969 7 1 2 50952 23968
0 23970 5 1 1 23969
0 23971 7 1 2 49539 58600
0 23972 5 1 1 23971
0 23973 7 1 2 23970 23972
0 23974 5 1 1 23973
0 23975 7 1 2 48628 23974
0 23976 5 1 1 23975
0 23977 7 1 2 53123 58798
0 23978 5 1 1 23977
0 23979 7 1 2 23976 23978
0 23980 5 1 1 23979
0 23981 7 1 2 42843 23980
0 23982 5 1 1 23981
0 23983 7 1 2 64876 65065
0 23984 5 1 1 23983
0 23985 7 1 2 23982 23984
0 23986 5 1 1 23985
0 23987 7 1 2 44805 23986
0 23988 5 1 1 23987
0 23989 7 1 2 23966 23988
0 23990 5 1 1 23989
0 23991 7 1 2 44933 23990
0 23992 5 1 1 23991
0 23993 7 1 2 49995 65235
0 23994 5 1 1 23993
0 23995 7 1 2 23663 23994
0 23996 5 1 1 23995
0 23997 7 1 2 49292 23996
0 23998 5 1 1 23997
0 23999 7 1 2 49002 52938
0 24000 7 1 2 67858 23999
0 24001 5 1 1 24000
0 24002 7 1 2 23998 24001
0 24003 5 1 1 24002
0 24004 7 1 2 52164 24003
0 24005 5 1 1 24004
0 24006 7 1 2 23992 24005
0 24007 5 1 1 24006
0 24008 7 1 2 42579 24007
0 24009 5 1 1 24008
0 24010 7 1 2 54593 5357
0 24011 5 1 1 24010
0 24012 7 1 2 50781 24011
0 24013 5 1 1 24012
0 24014 7 1 2 43330 68963
0 24015 5 1 1 24014
0 24016 7 1 2 54737 24015
0 24017 5 1 1 24016
0 24018 7 1 2 45266 24017
0 24019 5 1 1 24018
0 24020 7 1 2 24013 24019
0 24021 5 1 1 24020
0 24022 7 1 2 56021 69013
0 24023 7 1 2 24021 24022
0 24024 5 1 1 24023
0 24025 7 1 2 24009 24024
0 24026 5 2 1 24025
0 24027 7 1 2 65696 69039
0 24028 5 1 1 24027
0 24029 7 1 2 68935 68709
0 24030 5 1 1 24029
0 24031 7 2 2 56659 58225
0 24032 5 1 1 69041
0 24033 7 1 2 23848 24032
0 24034 5 1 1 24033
0 24035 7 1 2 65316 24034
0 24036 5 1 1 24035
0 24037 7 1 2 24030 24036
0 24038 5 2 1 24037
0 24039 7 1 2 61527 65802
0 24040 7 1 2 69043 24039
0 24041 5 1 1 24040
0 24042 7 1 2 24028 24041
0 24043 5 1 1 24042
0 24044 7 1 2 42210 67046
0 24045 5 1 1 24044
0 24046 7 1 2 59000 67014
0 24047 5 1 1 24046
0 24048 7 1 2 24045 24047
0 24049 5 3 1 24048
0 24050 7 1 2 59159 69045
0 24051 7 1 2 24043 24050
0 24052 5 1 1 24051
0 24053 7 1 2 45600 24052
0 24054 7 1 2 23956 24053
0 24055 5 1 1 24054
0 24056 7 1 2 23873 24055
0 24057 5 1 1 24056
0 24058 7 1 2 44585 24057
0 24059 5 1 1 24058
0 24060 7 1 2 43755 24059
0 24061 7 1 2 23174 24060
0 24062 5 1 1 24061
0 24063 7 1 2 42844 52362
0 24064 5 1 1 24063
0 24065 7 1 2 61960 24064
0 24066 5 1 1 24065
0 24067 7 1 2 43111 56644
0 24068 5 1 1 24067
0 24069 7 1 2 46278 24068
0 24070 5 1 1 24069
0 24071 7 1 2 47436 24070
0 24072 5 1 1 24071
0 24073 7 1 2 22943 24072
0 24074 5 1 1 24073
0 24075 7 1 2 47304 24074
0 24076 5 1 1 24075
0 24077 7 1 2 24066 24076
0 24078 5 1 1 24077
0 24079 7 1 2 44934 24078
0 24080 5 1 1 24079
0 24081 7 1 2 54727 61481
0 24082 5 1 1 24081
0 24083 7 1 2 44935 56149
0 24084 5 1 1 24083
0 24085 7 1 2 24082 24084
0 24086 5 1 1 24085
0 24087 7 1 2 51439 24086
0 24088 5 1 1 24087
0 24089 7 1 2 24088 23005
0 24090 7 1 2 24080 24089
0 24091 5 1 1 24090
0 24092 7 1 2 46054 24091
0 24093 5 1 1 24092
0 24094 7 1 2 23016 24093
0 24095 5 1 1 24094
0 24096 7 1 2 45105 24095
0 24097 5 1 1 24096
0 24098 7 1 2 54036 59626
0 24099 5 1 1 24098
0 24100 7 1 2 48818 53407
0 24101 5 1 1 24100
0 24102 7 1 2 24099 24101
0 24103 5 1 1 24102
0 24104 7 1 2 46706 24103
0 24105 5 1 1 24104
0 24106 7 2 2 49344 50782
0 24107 7 1 2 51007 69048
0 24108 5 1 1 24107
0 24109 7 1 2 5048 61829
0 24110 7 1 2 24108 24109
0 24111 5 1 1 24110
0 24112 7 1 2 45267 24111
0 24113 5 1 1 24112
0 24114 7 1 2 24105 24113
0 24115 5 1 1 24114
0 24116 7 1 2 47305 24115
0 24117 5 1 1 24116
0 24118 7 2 2 43331 51440
0 24119 5 2 1 69050
0 24120 7 1 2 52771 69051
0 24121 5 1 1 24120
0 24122 7 1 2 61610 68740
0 24123 5 1 1 24122
0 24124 7 1 2 24121 24123
0 24125 7 1 2 24117 24124
0 24126 5 1 1 24125
0 24127 7 1 2 48457 24126
0 24128 5 1 1 24127
0 24129 7 1 2 54117 67072
0 24130 5 1 1 24129
0 24131 7 1 2 53494 58391
0 24132 5 1 1 24131
0 24133 7 1 2 57127 24132
0 24134 5 1 1 24133
0 24135 7 1 2 53408 24134
0 24136 5 1 1 24135
0 24137 7 1 2 24130 24136
0 24138 7 1 2 24128 24137
0 24139 5 1 1 24138
0 24140 7 1 2 53986 24139
0 24141 5 1 1 24140
0 24142 7 1 2 24097 24141
0 24143 5 1 1 24142
0 24144 7 1 2 68931 24143
0 24145 5 1 1 24144
0 24146 7 1 2 49996 56509
0 24147 7 1 2 65279 24146
0 24148 7 1 2 58832 24147
0 24149 5 1 1 24148
0 24150 7 1 2 24145 24149
0 24151 5 1 1 24150
0 24152 7 1 2 48130 24151
0 24153 5 1 1 24152
0 24154 7 1 2 68932 68737
0 24155 5 1 1 24154
0 24156 7 1 2 24153 24155
0 24157 5 1 1 24156
0 24158 7 1 2 54784 24157
0 24159 5 1 1 24158
0 24160 7 2 2 53648 59020
0 24161 7 1 2 68772 69054
0 24162 5 1 1 24161
0 24163 7 1 2 24159 24162
0 24164 5 1 1 24163
0 24165 7 1 2 44337 24164
0 24166 5 1 1 24165
0 24167 7 1 2 66761 68791
0 24168 5 1 1 24167
0 24169 7 1 2 24166 24168
0 24170 5 1 1 24169
0 24171 7 1 2 45841 24170
0 24172 5 1 1 24171
0 24173 7 2 2 56282 62698
0 24174 7 1 2 68811 69056
0 24175 5 1 1 24174
0 24176 7 1 2 24172 24175
0 24177 5 1 1 24176
0 24178 7 1 2 47908 24177
0 24179 5 1 1 24178
0 24180 7 4 2 44338 44586
0 24181 7 2 2 61528 64914
0 24182 7 1 2 51441 69062
0 24183 5 1 1 24182
0 24184 7 1 2 23120 24183
0 24185 5 1 1 24184
0 24186 7 1 2 45106 24185
0 24187 5 1 1 24186
0 24188 7 1 2 54300 60218
0 24189 5 1 1 24188
0 24190 7 1 2 68915 24189
0 24191 5 1 1 24190
0 24192 7 1 2 24187 24191
0 24193 5 1 1 24192
0 24194 7 1 2 58243 24193
0 24195 5 1 1 24194
0 24196 7 1 2 68849 68801
0 24197 5 1 1 24196
0 24198 7 1 2 54408 68945
0 24199 7 1 2 68803 24198
0 24200 5 1 1 24199
0 24201 7 1 2 24197 24200
0 24202 5 1 1 24201
0 24203 7 1 2 48458 24202
0 24204 5 1 1 24203
0 24205 7 1 2 24195 24204
0 24206 5 1 1 24205
0 24207 7 1 2 48011 24206
0 24208 5 1 1 24207
0 24209 7 1 2 24208 23146
0 24210 5 1 1 24209
0 24211 7 1 2 42316 24210
0 24212 5 1 1 24211
0 24213 7 3 2 45842 61345
0 24214 7 1 2 65066 69064
0 24215 7 1 2 68785 24214
0 24216 5 1 1 24215
0 24217 7 1 2 24212 24216
0 24218 5 1 1 24217
0 24219 7 1 2 53705 24218
0 24220 5 1 1 24219
0 24221 7 1 2 52407 52482
0 24222 5 1 1 24221
0 24223 7 1 2 3875 24222
0 24224 5 1 1 24223
0 24225 7 1 2 43927 24224
0 24226 5 1 1 24225
0 24227 7 1 2 55255 64882
0 24228 5 1 1 24227
0 24229 7 1 2 48268 24228
0 24230 5 1 1 24229
0 24231 7 1 2 24226 24230
0 24232 5 1 1 24231
0 24233 7 1 2 68794 24232
0 24234 5 1 1 24233
0 24235 7 1 2 49404 64883
0 24236 5 1 1 24235
0 24237 7 1 2 44936 24236
0 24238 5 1 1 24237
0 24239 7 1 2 68562 24238
0 24240 5 1 1 24239
0 24241 7 1 2 51008 24240
0 24242 5 1 1 24241
0 24243 7 1 2 68555 24242
0 24244 5 1 1 24243
0 24245 7 1 2 68642 24244
0 24246 5 1 1 24245
0 24247 7 1 2 24234 24246
0 24248 5 1 1 24247
0 24249 7 1 2 46055 24248
0 24250 5 1 1 24249
0 24251 7 1 2 44806 68971
0 24252 5 1 1 24251
0 24253 7 2 2 52452 53835
0 24254 7 1 2 57215 69067
0 24255 5 1 1 24254
0 24256 7 1 2 24252 24255
0 24257 5 1 1 24256
0 24258 7 1 2 42580 24257
0 24259 5 1 1 24258
0 24260 7 1 2 24250 24259
0 24261 5 1 1 24260
0 24262 7 8 2 45843 44675
0 24263 5 2 1 69069
0 24264 7 4 2 53597 69070
0 24265 7 1 2 48903 69079
0 24266 7 1 2 24261 24265
0 24267 5 1 1 24266
0 24268 7 1 2 24220 24267
0 24269 5 1 1 24268
0 24270 7 1 2 69058 24269
0 24271 5 1 1 24270
0 24272 7 1 2 47780 24271
0 24273 7 1 2 24179 24272
0 24274 5 1 1 24273
0 24275 7 1 2 42317 68624
0 24276 5 1 1 24275
0 24277 7 4 2 45844 66632
0 24278 7 1 2 56601 59367
0 24279 7 1 2 69083 24278
0 24280 7 1 2 68619 24279
0 24281 5 1 1 24280
0 24282 7 1 2 24276 24281
0 24283 5 1 1 24282
0 24284 7 1 2 47909 24283
0 24285 5 1 1 24284
0 24286 7 4 2 64430 66406
0 24287 7 1 2 54785 69087
0 24288 7 1 2 69040 24287
0 24289 5 1 1 24288
0 24290 7 1 2 24285 24289
0 24291 5 1 1 24290
0 24292 7 1 2 53598 24291
0 24293 5 1 1 24292
0 24294 7 2 2 49003 60959
0 24295 7 3 2 57274 63752
0 24296 7 1 2 69091 69093
0 24297 5 1 1 24296
0 24298 7 1 2 51442 59533
0 24299 5 1 1 24298
0 24300 7 1 2 24297 24299
0 24301 5 1 1 24300
0 24302 7 1 2 46707 24301
0 24303 5 1 1 24302
0 24304 7 2 2 45758 48967
0 24305 7 1 2 46511 69096
0 24306 7 1 2 67381 24305
0 24307 5 1 1 24306
0 24308 7 1 2 24303 24307
0 24309 5 1 1 24308
0 24310 7 1 2 48459 24309
0 24311 5 1 1 24310
0 24312 7 3 2 43470 59520
0 24313 7 1 2 44240 61855
0 24314 7 1 2 68844 24313
0 24315 7 1 2 69098 24314
0 24316 5 1 1 24315
0 24317 7 1 2 24311 24316
0 24318 5 1 1 24317
0 24319 7 1 2 47437 24318
0 24320 5 1 1 24319
0 24321 7 2 2 59124 59808
0 24322 7 1 2 65291 69101
0 24323 5 1 1 24322
0 24324 7 1 2 24320 24323
0 24325 5 1 1 24324
0 24326 7 1 2 66543 24325
0 24327 5 1 1 24326
0 24328 7 1 2 52226 52682
0 24329 5 1 1 24328
0 24330 7 1 2 6837 24329
0 24331 5 1 1 24330
0 24332 7 1 2 45845 59125
0 24333 7 1 2 68486 24332
0 24334 7 1 2 24331 24333
0 24335 5 1 1 24334
0 24336 7 1 2 24327 24335
0 24337 5 1 1 24336
0 24338 7 1 2 68710 24337
0 24339 5 1 1 24338
0 24340 7 4 2 42318 46708
0 24341 7 2 2 48939 69103
0 24342 5 2 1 69107
0 24343 7 2 2 50358 64303
0 24344 5 1 1 69111
0 24345 7 1 2 69109 24344
0 24346 5 1 1 24345
0 24347 7 1 2 59534 24346
0 24348 5 1 1 24347
0 24349 7 2 2 47670 61436
0 24350 7 1 2 59757 66782
0 24351 7 1 2 69113 24350
0 24352 5 1 1 24351
0 24353 7 1 2 24348 24352
0 24354 5 1 1 24353
0 24355 7 1 2 50560 24354
0 24356 5 1 1 24355
0 24357 7 1 2 49172 63168
0 24358 7 3 2 48940 65543
0 24359 7 1 2 64040 69115
0 24360 7 1 2 24357 24359
0 24361 5 1 1 24360
0 24362 7 1 2 24356 24361
0 24363 5 1 1 24362
0 24364 7 1 2 58244 24363
0 24365 5 1 1 24364
0 24366 7 1 2 58856 69094
0 24367 5 1 1 24366
0 24368 7 1 2 59521 63334
0 24369 7 1 2 64828 24368
0 24370 5 1 1 24369
0 24371 7 1 2 24367 24370
0 24372 5 1 1 24371
0 24373 7 1 2 62334 66544
0 24374 7 1 2 24372 24373
0 24375 5 1 1 24374
0 24376 7 1 2 24365 24375
0 24377 5 1 1 24376
0 24378 7 1 2 65317 24377
0 24379 5 1 1 24378
0 24380 7 1 2 24339 24379
0 24381 5 1 1 24380
0 24382 7 1 2 46279 24381
0 24383 5 1 1 24382
0 24384 7 1 2 45268 68834
0 24385 5 1 1 24384
0 24386 7 1 2 44937 52065
0 24387 7 1 2 53442 24386
0 24388 5 1 1 24387
0 24389 7 1 2 24385 24388
0 24390 5 1 1 24389
0 24391 7 1 2 49587 24390
0 24392 5 1 1 24391
0 24393 7 3 2 46709 68874
0 24394 5 1 1 69118
0 24395 7 1 2 52300 54613
0 24396 5 1 1 24395
0 24397 7 1 2 24394 24396
0 24398 5 1 1 24397
0 24399 7 1 2 64482 24398
0 24400 5 1 1 24399
0 24401 7 1 2 24392 24400
0 24402 5 1 1 24401
0 24403 7 1 2 61171 24402
0 24404 5 1 1 24403
0 24405 7 1 2 49112 67220
0 24406 7 3 2 44676 61346
0 24407 7 1 2 67731 69121
0 24408 7 1 2 24405 24407
0 24409 5 1 1 24408
0 24410 7 1 2 24404 24409
0 24411 5 1 1 24410
0 24412 7 1 2 42319 24411
0 24413 5 1 1 24412
0 24414 7 1 2 54361 57253
0 24415 7 2 2 54220 64101
0 24416 7 1 2 56099 69124
0 24417 7 1 2 24414 24416
0 24418 5 1 1 24417
0 24419 7 1 2 24413 24418
0 24420 5 1 1 24419
0 24421 7 1 2 44587 24420
0 24422 5 1 1 24421
0 24423 7 1 2 48629 51346
0 24424 7 1 2 61735 66574
0 24425 7 1 2 67706 24424
0 24426 7 1 2 24423 24425
0 24427 7 1 2 68638 24426
0 24428 5 1 1 24427
0 24429 7 1 2 24422 24428
0 24430 5 1 1 24429
0 24431 7 1 2 59126 59331
0 24432 7 1 2 24430 24431
0 24433 5 1 1 24432
0 24434 7 1 2 24383 24433
0 24435 5 1 1 24434
0 24436 7 1 2 42034 24435
0 24437 5 1 1 24436
0 24438 7 2 2 48941 64113
0 24439 7 1 2 64910 69126
0 24440 7 1 2 59582 24439
0 24441 7 1 2 69044 24440
0 24442 5 1 1 24441
0 24443 7 1 2 44464 24442
0 24444 7 1 2 24437 24443
0 24445 7 1 2 24293 24444
0 24446 5 1 1 24445
0 24447 7 1 2 43756 24446
0 24448 7 1 2 24274 24447
0 24449 5 1 1 24448
0 24450 7 4 2 46710 54786
0 24451 7 4 2 44938 50140
0 24452 7 1 2 58410 69132
0 24453 5 1 1 24452
0 24454 7 2 2 55343 59705
0 24455 5 1 1 69136
0 24456 7 1 2 42581 55939
0 24457 7 1 2 24455 24456
0 24458 5 1 1 24457
0 24459 7 1 2 44807 1488
0 24460 7 1 2 65243 24459
0 24461 7 1 2 24458 24460
0 24462 5 1 1 24461
0 24463 7 1 2 24453 24462
0 24464 5 1 1 24463
0 24465 7 1 2 48460 24464
0 24466 5 1 1 24465
0 24467 7 2 2 44075 44808
0 24468 7 1 2 56531 69138
0 24469 7 1 2 58245 24468
0 24470 5 1 1 24469
0 24471 7 1 2 24466 24470
0 24472 5 1 1 24471
0 24473 7 1 2 66837 24472
0 24474 5 1 1 24473
0 24475 7 1 2 52970 59424
0 24476 7 1 2 59657 69065
0 24477 7 1 2 24475 24476
0 24478 5 1 1 24477
0 24479 7 1 2 24474 24478
0 24480 5 1 1 24479
0 24481 7 1 2 69128 24480
0 24482 5 1 1 24481
0 24483 7 1 2 47671 58219
0 24484 7 1 2 64461 24483
0 24485 7 2 2 58308 63945
0 24486 7 3 2 45601 52483
0 24487 7 1 2 55120 69142
0 24488 7 1 2 69140 24487
0 24489 7 1 2 24484 24488
0 24490 5 1 1 24489
0 24491 7 1 2 24482 24490
0 24492 5 1 1 24491
0 24493 7 1 2 45269 24492
0 24494 5 1 1 24493
0 24495 7 4 2 44588 62126
0 24496 7 1 2 52453 54247
0 24497 5 1 1 24496
0 24498 7 1 2 22571 24497
0 24499 5 2 1 24498
0 24500 7 3 2 69145 69149
0 24501 7 1 2 60602 64685
0 24502 7 1 2 69151 24501
0 24503 5 1 1 24502
0 24504 7 2 2 52484 58790
0 24505 5 1 1 69154
0 24506 7 1 2 65516 69155
0 24507 5 1 1 24506
0 24508 7 1 2 53783 62316
0 24509 5 1 1 24508
0 24510 7 1 2 24507 24509
0 24511 5 1 1 24510
0 24512 7 1 2 60538 68350
0 24513 7 1 2 24511 24512
0 24514 5 1 1 24513
0 24515 7 1 2 24503 24514
0 24516 5 1 1 24515
0 24517 7 1 2 44809 24516
0 24518 5 1 1 24517
0 24519 7 2 2 56603 64894
0 24520 7 1 2 54221 61871
0 24521 7 1 2 61763 24520
0 24522 7 1 2 66688 24521
0 24523 7 1 2 69156 24522
0 24524 5 1 1 24523
0 24525 7 1 2 24518 24524
0 24526 5 1 1 24525
0 24527 7 1 2 42582 24526
0 24528 5 1 1 24527
0 24529 7 1 2 53139 66879
0 24530 5 1 1 24529
0 24531 7 1 2 68455 68337
0 24532 5 1 1 24531
0 24533 7 1 2 24530 24532
0 24534 5 1 1 24533
0 24535 7 1 2 48131 53409
0 24536 7 1 2 24534 24535
0 24537 5 1 1 24536
0 24538 7 1 2 57635 64617
0 24539 7 1 2 50702 24538
0 24540 7 1 2 52971 24539
0 24541 5 1 1 24540
0 24542 7 1 2 24537 24541
0 24543 5 1 1 24542
0 24544 7 1 2 44939 24543
0 24545 5 1 1 24544
0 24546 7 4 2 43112 64618
0 24547 7 1 2 57875 58946
0 24548 7 1 2 67718 24547
0 24549 7 1 2 69158 24548
0 24550 5 1 1 24549
0 24551 7 1 2 24545 24550
0 24552 5 1 1 24551
0 24553 7 2 2 58064 67964
0 24554 7 1 2 61832 69162
0 24555 7 1 2 24552 24554
0 24556 5 1 1 24555
0 24557 7 1 2 24528 24556
0 24558 7 1 2 24494 24557
0 24559 5 1 1 24558
0 24560 7 1 2 53599 24559
0 24561 5 1 1 24560
0 24562 7 3 2 63407 67208
0 24563 7 1 2 48942 52630
0 24564 7 1 2 69164 24563
0 24565 5 1 1 24564
0 24566 7 1 2 46512 49381
0 24567 5 2 1 24566
0 24568 7 1 2 22955 69167
0 24569 5 1 1 24568
0 24570 7 2 2 44677 24569
0 24571 7 2 2 47910 64077
0 24572 7 1 2 43928 63116
0 24573 7 1 2 59758 24572
0 24574 7 1 2 69171 24573
0 24575 7 1 2 69169 24574
0 24576 5 1 1 24575
0 24577 7 1 2 24565 24576
0 24578 5 1 1 24577
0 24579 7 1 2 54389 24578
0 24580 5 1 1 24579
0 24581 7 1 2 52147 52981
0 24582 7 1 2 56875 64078
0 24583 7 1 2 24581 24582
0 24584 7 1 2 49382 50359
0 24585 7 1 2 66725 24584
0 24586 7 1 2 24583 24585
0 24587 5 1 1 24586
0 24588 7 1 2 24580 24587
0 24589 5 1 1 24588
0 24590 7 1 2 48269 24589
0 24591 5 1 1 24590
0 24592 7 1 2 49793 54578
0 24593 7 3 2 53686 56179
0 24594 7 1 2 56519 64471
0 24595 7 1 2 69173 24594
0 24596 7 1 2 24592 24595
0 24597 5 1 1 24596
0 24598 7 1 2 24591 24597
0 24599 5 1 1 24598
0 24600 7 1 2 44076 24599
0 24601 5 1 1 24600
0 24602 7 1 2 49383 60794
0 24603 7 1 2 63117 68273
0 24604 7 1 2 24602 24603
0 24605 7 1 2 61470 65639
0 24606 7 1 2 24604 24605
0 24607 5 1 1 24606
0 24608 7 3 2 44589 55489
0 24609 7 1 2 68715 69176
0 24610 7 1 2 69165 24609
0 24611 5 1 1 24610
0 24612 7 1 2 24607 24611
0 24613 5 1 1 24612
0 24614 7 1 2 42845 24613
0 24615 5 1 1 24614
0 24616 7 1 2 24601 24615
0 24617 5 1 1 24616
0 24618 7 1 2 46711 44810
0 24619 7 1 2 24617 24618
0 24620 5 1 1 24619
0 24621 7 2 2 59299 68980
0 24622 5 1 1 69179
0 24623 7 1 2 61347 62477
0 24624 7 1 2 63192 24623
0 24625 7 1 2 69157 24624
0 24626 7 1 2 69180 24625
0 24627 5 1 1 24626
0 24628 7 1 2 24620 24627
0 24629 7 1 2 24561 24628
0 24630 5 1 1 24629
0 24631 7 1 2 43757 24630
0 24632 5 1 1 24631
0 24633 7 1 2 55761 61559
0 24634 7 1 2 64398 24633
0 24635 7 2 2 57017 62837
0 24636 7 1 2 63548 69181
0 24637 7 1 2 24634 24636
0 24638 7 1 2 58649 24637
0 24639 5 1 1 24638
0 24640 7 1 2 24632 24639
0 24641 5 1 1 24640
0 24642 7 1 2 49224 24641
0 24643 5 1 1 24642
0 24644 7 1 2 51639 58627
0 24645 5 1 1 24644
0 24646 7 1 2 52835 3777
0 24647 5 3 1 24646
0 24648 7 1 2 68705 69183
0 24649 5 1 1 24648
0 24650 7 1 2 24645 24649
0 24651 5 1 1 24650
0 24652 7 1 2 57533 24651
0 24653 5 1 1 24652
0 24654 7 2 2 48968 55005
0 24655 7 1 2 68702 69186
0 24656 5 1 1 24655
0 24657 7 1 2 24653 24656
0 24658 5 1 1 24657
0 24659 7 1 2 43929 24658
0 24660 5 1 1 24659
0 24661 7 1 2 52563 58499
0 24662 7 1 2 67707 24661
0 24663 7 1 2 69184 24662
0 24664 5 1 1 24663
0 24665 7 1 2 24660 24664
0 24666 5 1 1 24665
0 24667 7 1 2 51354 24666
0 24668 5 1 1 24667
0 24669 7 1 2 44940 56143
0 24670 7 1 2 58325 24669
0 24671 7 1 2 60067 24670
0 24672 5 1 1 24671
0 24673 7 1 2 24668 24672
0 24674 5 3 1 24673
0 24675 7 1 2 58671 69188
0 24676 5 1 1 24675
0 24677 7 2 2 53364 56251
0 24678 7 1 2 47438 55654
0 24679 7 1 2 64238 24678
0 24680 7 2 2 69191 24679
0 24681 7 2 2 42211 55187
0 24682 7 1 2 56611 69195
0 24683 7 1 2 69193 24682
0 24684 5 1 1 24683
0 24685 7 1 2 24676 24684
0 24686 5 1 1 24685
0 24687 7 4 2 57914 68343
0 24688 7 1 2 45107 69197
0 24689 7 1 2 24686 24688
0 24690 5 1 1 24689
0 24691 7 1 2 24643 24690
0 24692 7 1 2 24449 24691
0 24693 5 1 1 24692
0 24694 7 1 2 66262 24693
0 24695 5 1 1 24694
0 24696 7 1 2 50613 64926
0 24697 5 1 1 24696
0 24698 7 1 2 49450 62276
0 24699 5 1 1 24698
0 24700 7 1 2 64519 24699
0 24701 7 1 2 24697 24700
0 24702 5 1 1 24701
0 24703 7 1 2 43930 24702
0 24704 5 1 1 24703
0 24705 7 1 2 42583 53764
0 24706 5 1 1 24705
0 24707 7 1 2 24704 24706
0 24708 5 1 1 24707
0 24709 7 1 2 43332 24708
0 24710 5 1 1 24709
0 24711 7 1 2 49698 55316
0 24712 5 1 1 24711
0 24713 7 1 2 46056 24712
0 24714 5 1 1 24713
0 24715 7 1 2 53124 24714
0 24716 5 1 1 24715
0 24717 7 1 2 24710 24716
0 24718 5 1 1 24717
0 24719 7 4 2 42320 43638
0 24720 5 1 1 69201
0 24721 7 1 2 67616 69202
0 24722 7 1 2 24718 24721
0 24723 5 1 1 24722
0 24724 7 1 2 54194 56371
0 24725 5 1 1 24724
0 24726 7 1 2 64345 24725
0 24727 5 1 1 24726
0 24728 7 1 2 52631 58434
0 24729 5 1 1 24728
0 24730 7 1 2 24727 24729
0 24731 5 1 1 24730
0 24732 7 1 2 17079 20766
0 24733 5 10 1 24732
0 24734 7 1 2 48012 69205
0 24735 7 1 2 53819 24734
0 24736 7 1 2 24731 24735
0 24737 5 1 1 24736
0 24738 7 1 2 24723 24737
0 24739 5 1 1 24738
0 24740 7 1 2 42846 24739
0 24741 5 1 1 24740
0 24742 7 5 2 48461 65697
0 24743 7 1 2 68693 69215
0 24744 7 1 2 56672 24743
0 24745 5 1 1 24744
0 24746 7 1 2 24741 24745
0 24747 5 1 1 24746
0 24748 7 1 2 48270 24747
0 24749 5 1 1 24748
0 24750 7 2 2 49859 58309
0 24751 7 2 2 69206 69220
0 24752 7 1 2 64350 69222
0 24753 5 1 1 24752
0 24754 7 1 2 45108 53825
0 24755 5 1 1 24754
0 24756 7 1 2 44077 23279
0 24757 5 1 1 24756
0 24758 7 1 2 46513 52366
0 24759 7 1 2 24757 24758
0 24760 5 1 1 24759
0 24761 7 1 2 24755 24760
0 24762 5 1 1 24761
0 24763 7 1 2 47306 24762
0 24764 5 1 1 24763
0 24765 7 1 2 62346 65046
0 24766 5 1 1 24765
0 24767 7 1 2 24764 24766
0 24768 5 1 1 24767
0 24769 7 1 2 46712 24768
0 24770 5 1 1 24769
0 24771 7 1 2 52982 53098
0 24772 5 1 1 24771
0 24773 7 1 2 24770 24772
0 24774 5 1 1 24773
0 24775 7 1 2 46280 24774
0 24776 5 1 1 24775
0 24777 7 1 2 47439 65309
0 24778 5 1 1 24777
0 24779 7 1 2 24776 24778
0 24780 5 1 1 24779
0 24781 7 1 2 64399 66376
0 24782 7 1 2 24780 24781
0 24783 5 1 1 24782
0 24784 7 1 2 24753 24783
0 24785 5 1 1 24784
0 24786 7 1 2 68113 24785
0 24787 5 1 1 24786
0 24788 7 1 2 24749 24787
0 24789 5 1 1 24788
0 24790 7 1 2 63193 24789
0 24791 5 1 1 24790
0 24792 7 4 2 53836 54599
0 24793 7 1 2 55188 64431
0 24794 7 1 2 64388 24793
0 24795 7 1 2 69207 24794
0 24796 7 1 2 69224 24795
0 24797 5 1 1 24796
0 24798 7 1 2 43599 24797
0 24799 7 1 2 24791 24798
0 24800 5 1 1 24799
0 24801 7 2 2 44678 63665
0 24802 7 1 2 64297 69228
0 24803 7 1 2 69068 24802
0 24804 5 1 1 24803
0 24805 7 1 2 52632 59638
0 24806 7 3 2 48271 61348
0 24807 7 4 2 55762 59680
0 24808 7 1 2 69230 69233
0 24809 7 1 2 24805 24808
0 24810 5 1 1 24809
0 24811 7 1 2 24804 24810
0 24812 5 1 1 24811
0 24813 7 1 2 46713 24812
0 24814 5 1 1 24813
0 24815 7 1 2 42584 54614
0 24816 5 1 1 24815
0 24817 7 1 2 58622 24816
0 24818 5 5 1 24817
0 24819 7 1 2 49540 65337
0 24820 7 1 2 69234 24819
0 24821 7 1 2 69237 24820
0 24822 5 1 1 24821
0 24823 7 1 2 24814 24822
0 24824 5 1 1 24823
0 24825 7 1 2 66377 24824
0 24826 5 1 1 24825
0 24827 7 2 2 68208 69225
0 24828 7 1 2 47029 58398
0 24829 7 1 2 67775 24828
0 24830 7 1 2 69242 24829
0 24831 5 1 1 24830
0 24832 7 1 2 24826 24831
0 24833 5 1 1 24832
0 24834 7 1 2 42321 24833
0 24835 5 1 1 24834
0 24836 7 1 2 43639 63291
0 24837 7 2 2 66040 24836
0 24838 7 1 2 64389 69244
0 24839 7 1 2 69243 24838
0 24840 5 1 1 24839
0 24841 7 1 2 46988 24840
0 24842 7 1 2 24835 24841
0 24843 5 1 1 24842
0 24844 7 1 2 42212 24843
0 24845 7 1 2 24800 24844
0 24846 5 1 1 24845
0 24847 7 2 2 47672 69226
0 24848 7 1 2 67549 69208
0 24849 5 1 1 24848
0 24850 7 1 2 48013 65884
0 24851 5 1 1 24850
0 24852 7 1 2 24849 24851
0 24853 5 1 1 24852
0 24854 7 1 2 53630 24853
0 24855 5 1 1 24854
0 24856 7 1 2 65830 65851
0 24857 7 1 2 68472 24856
0 24858 5 1 1 24857
0 24859 7 1 2 24855 24858
0 24860 5 1 1 24859
0 24861 7 1 2 55189 61204
0 24862 7 1 2 24860 24861
0 24863 7 1 2 69246 24862
0 24864 5 1 1 24863
0 24865 7 1 2 24846 24864
0 24866 5 1 1 24865
0 24867 7 1 2 42035 24866
0 24868 5 1 1 24867
0 24869 7 8 2 43547 67694
0 24870 7 2 2 47030 69248
0 24871 7 1 2 67739 69256
0 24872 5 1 1 24871
0 24873 7 1 2 43640 68082
0 24874 7 1 2 68473 24873
0 24875 5 1 1 24874
0 24876 7 2 2 24872 24875
0 24877 5 1 1 69258
0 24878 7 3 2 53600 69209
0 24879 7 1 2 67550 69260
0 24880 5 1 1 24879
0 24881 7 1 2 69259 24880
0 24882 5 1 1 24881
0 24883 7 1 2 43471 24882
0 24884 5 1 1 24883
0 24885 7 4 2 43641 67187
0 24886 7 3 2 60677 69263
0 24887 5 1 1 69267
0 24888 7 1 2 69249 69268
0 24889 5 1 1 24888
0 24890 7 1 2 24884 24889
0 24891 5 1 1 24890
0 24892 7 1 2 57018 58257
0 24893 7 1 2 69247 24892
0 24894 7 1 2 24891 24893
0 24895 5 1 1 24894
0 24896 7 1 2 44465 24895
0 24897 7 1 2 24868 24896
0 24898 5 1 1 24897
0 24899 7 4 2 52787 54787
0 24900 7 2 2 46714 67535
0 24901 5 2 1 69274
0 24902 7 1 2 48819 69276
0 24903 5 1 1 24902
0 24904 7 1 2 45463 67545
0 24905 5 1 1 24904
0 24906 7 1 2 66378 24905
0 24907 7 1 2 24903 24906
0 24908 5 1 1 24907
0 24909 7 1 2 49592 65852
0 24910 7 1 2 67695 24909
0 24911 5 1 1 24910
0 24912 7 1 2 24908 24911
0 24913 5 1 1 24912
0 24914 7 1 2 42322 24913
0 24915 5 1 1 24914
0 24916 7 4 2 42406 46715
0 24917 7 4 2 66063 69278
0 24918 7 1 2 66083 69282
0 24919 5 1 1 24918
0 24920 7 1 2 24915 24919
0 24921 5 1 1 24920
0 24922 7 2 2 52633 24921
0 24923 7 1 2 50614 69286
0 24924 5 1 1 24923
0 24925 7 2 2 52634 68160
0 24926 7 2 2 49497 54646
0 24927 7 1 2 69288 69290
0 24928 5 1 1 24927
0 24929 7 1 2 24924 24928
0 24930 5 1 1 24929
0 24931 7 1 2 68425 24930
0 24932 5 1 1 24931
0 24933 7 3 2 44241 56348
0 24934 7 1 2 46989 69292
0 24935 5 1 1 24934
0 24936 7 1 2 43600 66107
0 24937 5 1 1 24936
0 24938 7 1 2 24935 24937
0 24939 5 2 1 24938
0 24940 7 1 2 66379 69295
0 24941 5 1 1 24940
0 24942 7 1 2 65880 69293
0 24943 5 1 1 24942
0 24944 7 1 2 24941 24943
0 24945 5 1 1 24944
0 24946 7 1 2 43333 24945
0 24947 5 1 1 24946
0 24948 7 2 2 49050 67540
0 24949 5 1 1 69297
0 24950 7 1 2 66380 69298
0 24951 5 1 1 24950
0 24952 7 1 2 24947 24951
0 24953 5 1 1 24952
0 24954 7 1 2 42323 24953
0 24955 5 1 1 24954
0 24956 7 1 2 49541 66427
0 24957 5 1 1 24956
0 24958 7 1 2 24955 24957
0 24959 5 1 1 24958
0 24960 7 1 2 49699 69238
0 24961 7 1 2 24959 24960
0 24962 5 1 1 24961
0 24963 7 1 2 24932 24962
0 24964 5 1 1 24963
0 24965 7 1 2 43113 24964
0 24966 5 1 1 24965
0 24967 7 1 2 49700 68426
0 24968 7 1 2 69287 24967
0 24969 5 1 1 24968
0 24970 7 1 2 24966 24969
0 24971 5 1 1 24970
0 24972 7 1 2 42847 24971
0 24973 5 1 1 24972
0 24974 7 1 2 51636 58042
0 24975 7 2 2 43642 67696
0 24976 7 3 2 42324 54973
0 24977 7 1 2 68248 69301
0 24978 7 1 2 69299 24977
0 24979 7 1 2 24974 24978
0 24980 5 1 1 24979
0 24981 7 1 2 24973 24980
0 24982 5 1 1 24981
0 24983 7 1 2 69270 24982
0 24984 5 1 1 24983
0 24985 7 2 2 42407 46933
0 24986 7 4 2 43643 69304
0 24987 7 1 2 69306 69294
0 24988 5 1 1 24987
0 24989 7 1 2 66108 68098
0 24990 5 1 1 24989
0 24991 7 1 2 24988 24990
0 24992 5 1 1 24991
0 24993 7 1 2 45846 24992
0 24994 5 1 1 24993
0 24995 7 2 2 56349 67305
0 24996 7 1 2 46934 66317
0 24997 7 1 2 69310 24996
0 24998 5 1 1 24997
0 24999 7 1 2 24994 24998
0 25000 5 1 1 24999
0 25001 7 1 2 43601 25000
0 25002 5 1 1 25001
0 25003 7 1 2 60313 67621
0 25004 7 1 2 69311 25003
0 25005 5 1 1 25004
0 25006 7 1 2 25002 25005
0 25007 5 1 1 25006
0 25008 7 1 2 43334 25007
0 25009 5 1 1 25008
0 25010 7 1 2 65881 68416
0 25011 7 1 2 68328 25010
0 25012 5 1 1 25011
0 25013 7 1 2 25009 25012
0 25014 5 1 1 25013
0 25015 7 1 2 56577 59178
0 25016 7 1 2 69239 25015
0 25017 7 1 2 25014 25016
0 25018 5 1 1 25017
0 25019 7 1 2 55190 57280
0 25020 7 3 2 52696 25019
0 25021 7 1 2 24877 69312
0 25022 5 1 1 25021
0 25023 7 5 2 52097 52635
0 25024 7 4 2 48272 69315
0 25025 7 3 2 69122 69320
0 25026 7 2 2 45847 68099
0 25027 5 1 1 69327
0 25028 7 1 2 65523 69328
0 25029 7 1 2 69324 25028
0 25030 5 1 1 25029
0 25031 7 1 2 25022 25030
0 25032 5 1 1 25031
0 25033 7 1 2 45464 25032
0 25034 5 1 1 25033
0 25035 7 1 2 45848 67015
0 25036 5 1 1 25035
0 25037 7 1 2 65621 65882
0 25038 5 1 1 25037
0 25039 7 1 2 25036 25038
0 25040 5 1 1 25039
0 25041 7 2 2 52527 52636
0 25042 7 2 2 48014 55381
0 25043 7 1 2 48273 69331
0 25044 7 1 2 69329 25043
0 25045 7 1 2 59347 25044
0 25046 7 1 2 25040 25045
0 25047 5 1 1 25046
0 25048 7 1 2 25034 25047
0 25049 5 1 1 25048
0 25050 7 1 2 47563 25049
0 25051 5 1 1 25050
0 25052 7 1 2 67551 69313
0 25053 5 1 1 25052
0 25054 7 1 2 46990 69325
0 25055 5 1 1 25054
0 25056 7 1 2 25053 25055
0 25057 5 1 1 25056
0 25058 7 1 2 49173 25057
0 25059 5 1 1 25058
0 25060 7 1 2 55258 63227
0 25061 7 1 2 51764 25060
0 25062 7 1 2 69240 25061
0 25063 5 1 1 25062
0 25064 7 1 2 25059 25063
0 25065 5 1 1 25064
0 25066 7 1 2 69261 25065
0 25067 5 1 1 25066
0 25068 7 1 2 25051 25067
0 25069 7 1 2 25018 25068
0 25070 5 1 1 25069
0 25071 7 1 2 48904 25070
0 25072 5 1 1 25071
0 25073 7 1 2 24984 25072
0 25074 5 1 1 25073
0 25075 7 1 2 44339 25074
0 25076 5 1 1 25075
0 25077 7 2 2 42036 67047
0 25078 5 1 1 69333
0 25079 7 1 2 53692 68663
0 25080 5 1 1 25079
0 25081 7 1 2 25078 25080
0 25082 5 10 1 25081
0 25083 7 1 2 42213 69335
0 25084 5 1 1 25083
0 25085 7 1 2 59693 66164
0 25086 5 1 1 25085
0 25087 7 1 2 25084 25086
0 25088 5 1 1 25087
0 25089 7 3 2 51204 66109
0 25090 7 1 2 25088 69345
0 25091 5 1 1 25090
0 25092 7 1 2 66263 69271
0 25093 5 1 1 25092
0 25094 7 1 2 63421 66748
0 25095 7 1 2 67627 25094
0 25096 5 1 1 25095
0 25097 7 1 2 25093 25096
0 25098 5 2 1 25097
0 25099 7 1 2 53339 66633
0 25100 7 1 2 69348 25099
0 25101 5 1 1 25100
0 25102 7 1 2 25091 25101
0 25103 5 1 1 25102
0 25104 7 1 2 53505 25103
0 25105 5 1 1 25104
0 25106 7 1 2 44078 55534
0 25107 7 2 2 68836 25106
0 25108 7 1 2 69350 69349
0 25109 5 1 1 25108
0 25110 7 1 2 25105 25109
0 25111 5 1 1 25110
0 25112 7 1 2 69231 25111
0 25113 5 1 1 25112
0 25114 7 4 2 55326 63267
0 25115 7 3 2 53987 54575
0 25116 7 2 2 69352 69356
0 25117 7 1 2 44679 66674
0 25118 7 1 2 69307 25117
0 25119 5 1 1 25118
0 25120 7 1 2 53601 65853
0 25121 7 1 2 67552 25120
0 25122 5 1 1 25121
0 25123 7 1 2 25119 25122
0 25124 5 1 1 25123
0 25125 7 1 2 48905 25124
0 25126 5 1 1 25125
0 25127 7 2 2 43644 67812
0 25128 7 1 2 54788 69250
0 25129 7 1 2 69361 25128
0 25130 5 1 1 25129
0 25131 7 1 2 25126 25130
0 25132 5 1 1 25131
0 25133 7 1 2 69359 25132
0 25134 5 1 1 25133
0 25135 7 1 2 25113 25134
0 25136 5 1 1 25135
0 25137 7 1 2 44340 25136
0 25138 5 1 1 25137
0 25139 7 1 2 46850 58258
0 25140 7 1 2 66675 25139
0 25141 7 1 2 52285 65054
0 25142 7 1 2 69308 69229
0 25143 7 1 2 25141 25142
0 25144 7 1 2 25140 25143
0 25145 5 1 1 25144
0 25146 7 1 2 42325 25145
0 25147 7 1 2 25138 25146
0 25148 5 1 1 25147
0 25149 7 1 2 63194 67697
0 25150 5 1 1 25149
0 25151 7 1 2 63313 68500
0 25152 5 1 1 25151
0 25153 7 1 2 25150 25152
0 25154 5 1 1 25153
0 25155 7 1 2 42037 25154
0 25156 5 1 1 25155
0 25157 7 1 2 58079 69251
0 25158 5 1 1 25157
0 25159 7 2 2 53649 63228
0 25160 5 1 1 69363
0 25161 7 1 2 25158 25160
0 25162 5 2 1 25161
0 25163 7 1 2 66848 69365
0 25164 5 1 1 25163
0 25165 7 1 2 25156 25164
0 25166 5 1 1 25165
0 25167 7 1 2 47440 25166
0 25168 5 1 1 25167
0 25169 7 1 2 49174 59915
0 25170 7 1 2 69252 25169
0 25171 5 1 1 25170
0 25172 7 1 2 25168 25171
0 25173 5 1 1 25172
0 25174 7 1 2 46514 25173
0 25175 5 1 1 25174
0 25176 7 3 2 47564 61437
0 25177 7 1 2 48906 62715
0 25178 7 1 2 63396 25177
0 25179 7 1 2 69367 25178
0 25180 5 1 1 25179
0 25181 7 1 2 25175 25180
0 25182 5 1 1 25181
0 25183 7 1 2 69357 25182
0 25184 5 1 1 25183
0 25185 7 4 2 44341 48274
0 25186 7 1 2 43335 69296
0 25187 5 1 1 25186
0 25188 7 1 2 25187 24949
0 25189 5 2 1 25188
0 25190 7 1 2 53506 69374
0 25191 5 1 1 25190
0 25192 7 1 2 46991 69351
0 25193 5 1 1 25192
0 25194 7 1 2 25191 25193
0 25195 5 1 1 25194
0 25196 7 2 2 69370 25195
0 25197 7 1 2 55763 68621
0 25198 7 1 2 69376 25197
0 25199 5 1 1 25198
0 25200 7 1 2 25184 25199
0 25201 5 1 1 25200
0 25202 7 1 2 65854 25201
0 25203 5 1 1 25202
0 25204 7 1 2 67553 69360
0 25205 5 1 1 25204
0 25206 7 2 2 52637 69232
0 25207 7 1 2 63229 69378
0 25208 7 1 2 60783 25207
0 25209 5 1 1 25208
0 25210 7 1 2 25205 25209
0 25211 5 2 1 25210
0 25212 7 1 2 43548 69380
0 25213 5 1 1 25212
0 25214 7 2 2 64930 68875
0 25215 7 2 2 46935 61349
0 25216 7 1 2 67698 69384
0 25217 7 1 2 69382 25216
0 25218 5 1 1 25217
0 25219 7 1 2 25213 25218
0 25220 5 1 1 25219
0 25221 7 1 2 43645 67990
0 25222 7 1 2 25220 25221
0 25223 5 1 1 25222
0 25224 7 1 2 25203 25223
0 25225 5 1 1 25224
0 25226 7 1 2 45759 25225
0 25227 5 1 1 25226
0 25228 7 1 2 53650 69381
0 25229 5 1 1 25228
0 25230 7 2 2 69253 69383
0 25231 7 1 2 42848 55401
0 25232 7 1 2 69386 25231
0 25233 5 1 1 25232
0 25234 7 1 2 25229 25233
0 25235 5 1 1 25234
0 25236 7 1 2 42038 25235
0 25237 5 1 1 25236
0 25238 7 1 2 59989 60521
0 25239 7 1 2 69387 25238
0 25240 5 1 1 25239
0 25241 7 1 2 25237 25240
0 25242 5 1 1 25241
0 25243 7 1 2 44342 69362
0 25244 7 1 2 25242 25243
0 25245 5 1 1 25244
0 25246 7 1 2 45849 25245
0 25247 7 1 2 25227 25246
0 25248 5 1 1 25247
0 25249 7 1 2 45270 25248
0 25250 7 1 2 25148 25249
0 25251 5 1 1 25250
0 25252 7 1 2 47781 25251
0 25253 7 1 2 25076 25252
0 25254 5 1 1 25253
0 25255 7 1 2 24898 25254
0 25256 5 1 1 25255
0 25257 7 1 2 67546 69277
0 25258 5 2 1 25257
0 25259 7 1 2 58259 61923
0 25260 7 1 2 64079 25259
0 25261 7 2 2 51375 52280
0 25262 7 1 2 65055 69390
0 25263 7 1 2 25260 25262
0 25264 7 1 2 69262 25263
0 25265 5 1 1 25264
0 25266 7 1 2 44079 52186
0 25267 5 1 1 25266
0 25268 7 1 2 49630 25267
0 25269 5 3 1 25268
0 25270 7 3 2 62699 66381
0 25271 7 1 2 69392 69395
0 25272 7 2 2 48922 52788
0 25273 7 1 2 69398 69379
0 25274 7 1 2 25271 25273
0 25275 5 1 1 25274
0 25276 7 1 2 25265 25275
0 25277 5 1 1 25276
0 25278 7 1 2 69388 25277
0 25279 5 1 1 25278
0 25280 7 1 2 11188 24720
0 25281 5 1 1 25280
0 25282 7 1 2 48869 19567
0 25283 7 3 2 25281 25282
0 25284 7 1 2 42585 58119
0 25285 7 1 2 60522 25284
0 25286 7 1 2 69377 25285
0 25287 5 1 1 25286
0 25288 7 2 2 55327 62290
0 25289 5 1 1 69403
0 25290 7 1 2 46936 67703
0 25291 5 2 1 25290
0 25292 7 1 2 43549 63233
0 25293 5 1 1 25292
0 25294 7 5 2 69405 25293
0 25295 7 1 2 59846 69407
0 25296 7 1 2 69404 25295
0 25297 5 1 1 25296
0 25298 7 1 2 63234 22121
0 25299 5 1 1 25298
0 25300 7 2 2 69406 25299
0 25301 7 2 2 49175 49293
0 25302 7 1 2 59788 69414
0 25303 7 1 2 69412 25302
0 25304 5 1 1 25303
0 25305 7 1 2 25297 25304
0 25306 5 1 1 25305
0 25307 7 1 2 51009 69358
0 25308 7 1 2 25306 25307
0 25309 5 1 1 25308
0 25310 7 1 2 25287 25309
0 25311 5 1 1 25310
0 25312 7 1 2 45271 25311
0 25313 5 1 1 25312
0 25314 7 1 2 69408 69314
0 25315 5 1 1 25314
0 25316 7 1 2 62668 69326
0 25317 5 1 1 25316
0 25318 7 1 2 25315 25317
0 25319 5 1 1 25318
0 25320 7 1 2 45465 25319
0 25321 5 1 1 25320
0 25322 7 1 2 67536 69385
0 25323 7 1 2 69119 25322
0 25324 7 1 2 59348 25323
0 25325 5 1 1 25324
0 25326 7 1 2 25321 25325
0 25327 5 1 1 25326
0 25328 7 1 2 47565 25327
0 25329 5 1 1 25328
0 25330 7 1 2 56123 57550
0 25331 7 1 2 69241 25330
0 25332 7 1 2 69375 25331
0 25333 5 1 1 25332
0 25334 7 1 2 25329 25333
0 25335 5 1 1 25334
0 25336 7 1 2 59847 25335
0 25337 5 1 1 25336
0 25338 7 1 2 25313 25337
0 25339 5 1 1 25338
0 25340 7 1 2 47782 25339
0 25341 5 1 1 25340
0 25342 7 1 2 62560 69129
0 25343 7 1 2 69409 25342
0 25344 7 1 2 69227 25343
0 25345 5 1 1 25344
0 25346 7 1 2 25341 25345
0 25347 5 1 1 25346
0 25348 7 1 2 69400 25347
0 25349 5 1 1 25348
0 25350 7 1 2 25279 25349
0 25351 7 1 2 25256 25350
0 25352 5 1 1 25351
0 25353 7 1 2 44811 25352
0 25354 5 1 1 25353
0 25355 7 1 2 42039 69046
0 25356 5 1 1 25355
0 25357 7 7 2 67503 67813
0 25358 7 2 2 45602 69416
0 25359 5 1 1 69423
0 25360 7 1 2 43550 69424
0 25361 5 1 1 25360
0 25362 7 1 2 25356 25361
0 25363 5 3 1 25362
0 25364 7 1 2 43931 66099
0 25365 5 1 1 25364
0 25366 7 1 2 65823 25365
0 25367 5 1 1 25366
0 25368 7 6 2 47783 45272
0 25369 7 1 2 25367 69428
0 25370 7 1 2 69425 25369
0 25371 5 1 1 25370
0 25372 7 1 2 66418 69283
0 25373 7 1 2 69399 25372
0 25374 5 1 1 25373
0 25375 7 1 2 25371 25374
0 25376 5 1 1 25375
0 25377 7 1 2 47566 25376
0 25378 5 1 1 25377
0 25379 7 3 2 67328 69279
0 25380 7 4 2 45273 65999
0 25381 7 1 2 56237 69437
0 25382 7 1 2 69434 25381
0 25383 5 1 1 25382
0 25384 7 1 2 25378 25383
0 25385 5 1 1 25384
0 25386 7 1 2 48462 25385
0 25387 5 1 1 25386
0 25388 7 2 2 44242 68845
0 25389 7 1 2 64196 69002
0 25390 5 1 1 25389
0 25391 7 2 2 55847 66191
0 25392 7 1 2 61856 69443
0 25393 5 1 1 25392
0 25394 7 1 2 25390 25393
0 25395 5 1 1 25394
0 25396 7 1 2 43472 25395
0 25397 5 1 1 25396
0 25398 7 2 2 53640 66192
0 25399 7 1 2 64197 69445
0 25400 5 1 1 25399
0 25401 7 1 2 25397 25400
0 25402 5 1 1 25401
0 25403 7 1 2 65698 25402
0 25404 5 1 1 25403
0 25405 7 1 2 57915 58065
0 25406 7 1 2 68880 25405
0 25407 5 1 1 25406
0 25408 7 1 2 25404 25407
0 25409 5 1 1 25408
0 25410 7 1 2 42040 25409
0 25411 5 1 1 25410
0 25412 7 3 2 63967 66064
0 25413 7 2 2 61027 66471
0 25414 7 7 2 42326 62127
0 25415 7 1 2 69450 69452
0 25416 7 1 2 69447 25415
0 25417 5 1 1 25416
0 25418 7 1 2 25411 25417
0 25419 5 1 1 25418
0 25420 7 1 2 69441 25419
0 25421 5 1 1 25420
0 25422 7 1 2 25387 25421
0 25423 5 1 1 25422
0 25424 7 1 2 46057 25423
0 25425 5 1 1 25424
0 25426 7 1 2 53401 58947
0 25427 7 1 2 64462 25426
0 25428 7 1 2 65047 25427
0 25429 7 1 2 69426 25428
0 25430 5 1 1 25429
0 25431 7 1 2 25425 25430
0 25432 5 1 1 25431
0 25433 7 1 2 51010 25432
0 25434 5 1 1 25433
0 25435 7 1 2 63956 69047
0 25436 5 1 1 25435
0 25437 7 1 2 67209 69284
0 25438 5 1 1 25437
0 25439 7 1 2 25436 25438
0 25440 5 1 1 25439
0 25441 7 1 2 42041 25440
0 25442 5 1 1 25441
0 25443 7 2 2 61028 63957
0 25444 7 1 2 67091 69459
0 25445 5 1 1 25444
0 25446 7 1 2 25442 25445
0 25447 5 1 1 25446
0 25448 7 1 2 53815 25447
0 25449 5 1 1 25448
0 25450 7 2 2 62513 69417
0 25451 7 1 2 43551 52416
0 25452 7 1 2 69461 25451
0 25453 5 1 1 25452
0 25454 7 1 2 25449 25453
0 25455 5 1 1 25454
0 25456 7 1 2 56369 25455
0 25457 5 1 1 25456
0 25458 7 1 2 52807 56188
0 25459 7 1 2 67965 25458
0 25460 7 2 2 61857 66472
0 25461 7 1 2 67121 69463
0 25462 7 1 2 25459 25461
0 25463 5 1 1 25462
0 25464 7 1 2 25457 25463
0 25465 5 1 1 25464
0 25466 7 1 2 47307 25465
0 25467 5 1 1 25466
0 25468 7 1 2 52213 52301
0 25469 5 1 1 25468
0 25470 7 1 2 65287 25469
0 25471 5 1 1 25470
0 25472 7 2 2 44466 66065
0 25473 7 1 2 68244 68390
0 25474 7 2 2 69465 25473
0 25475 7 1 2 45274 69467
0 25476 7 1 2 25471 25475
0 25477 5 1 1 25476
0 25478 7 1 2 25467 25477
0 25479 5 1 1 25478
0 25480 7 1 2 66000 25479
0 25481 5 1 1 25480
0 25482 7 2 2 64383 66749
0 25483 7 1 2 53443 66685
0 25484 7 1 2 69469 25483
0 25485 5 1 1 25484
0 25486 7 2 2 62716 67309
0 25487 7 1 2 49841 67663
0 25488 7 1 2 69471 25487
0 25489 5 1 1 25488
0 25490 7 1 2 25485 25489
0 25491 5 1 1 25490
0 25492 7 1 2 46058 25491
0 25493 5 1 1 25492
0 25494 7 1 2 52588 58921
0 25495 7 1 2 51801 25494
0 25496 7 1 2 68878 25495
0 25497 5 1 1 25496
0 25498 7 1 2 25493 25497
0 25499 5 1 1 25498
0 25500 7 1 2 48630 25499
0 25501 5 1 1 25500
0 25502 7 3 2 46059 68892
0 25503 7 1 2 48463 60213
0 25504 7 1 2 69473 25503
0 25505 5 1 1 25504
0 25506 7 1 2 25501 25505
0 25507 5 1 1 25506
0 25508 7 1 2 42214 25507
0 25509 5 1 1 25508
0 25510 7 2 2 55019 68850
0 25511 5 1 1 69476
0 25512 7 1 2 55975 67016
0 25513 7 1 2 69477 25512
0 25514 5 1 1 25513
0 25515 7 1 2 25509 25514
0 25516 5 1 1 25515
0 25517 7 1 2 65906 25516
0 25518 5 1 1 25517
0 25519 7 1 2 58948 64400
0 25520 7 1 2 68861 25519
0 25521 7 1 2 69003 25520
0 25522 5 1 1 25521
0 25523 7 1 2 25518 25522
0 25524 5 1 1 25523
0 25525 7 1 2 43473 25524
0 25526 5 1 1 25525
0 25527 7 1 2 51443 65699
0 25528 5 1 1 25527
0 25529 7 1 2 65907 68851
0 25530 5 1 1 25529
0 25531 7 1 2 25528 25530
0 25532 5 1 1 25531
0 25533 7 1 2 48464 69448
0 25534 7 2 2 25532 25533
0 25535 7 1 2 56077 67765
0 25536 7 1 2 69478 25535
0 25537 5 1 1 25536
0 25538 7 1 2 25526 25537
0 25539 5 1 1 25538
0 25540 7 1 2 42042 25539
0 25541 5 1 1 25540
0 25542 7 4 2 42215 66473
0 25543 7 2 2 58260 69480
0 25544 7 1 2 69479 69484
0 25545 5 1 1 25544
0 25546 7 1 2 25541 25545
0 25547 5 1 1 25546
0 25548 7 1 2 49294 25547
0 25549 5 1 1 25548
0 25550 7 1 2 25481 25549
0 25551 7 1 2 25434 25550
0 25552 5 1 1 25551
0 25553 7 1 2 46281 25552
0 25554 5 1 1 25553
0 25555 7 1 2 52589 56001
0 25556 7 1 2 65844 25555
0 25557 7 2 2 56238 66733
0 25558 7 2 2 54974 55410
0 25559 7 1 2 69254 69488
0 25560 7 1 2 69486 25559
0 25561 7 1 2 25556 25560
0 25562 5 1 1 25561
0 25563 7 2 2 53140 57352
0 25564 7 1 2 68893 69490
0 25565 5 1 1 25564
0 25566 7 2 2 42408 68315
0 25567 7 1 2 58871 66066
0 25568 7 1 2 69492 25567
0 25569 5 1 1 25568
0 25570 7 1 2 25565 25569
0 25571 5 1 1 25570
0 25572 7 1 2 42216 54549
0 25573 7 1 2 25571 25572
0 25574 5 1 1 25573
0 25575 7 1 2 53141 61636
0 25576 7 1 2 66449 25575
0 25577 7 1 2 67017 25576
0 25578 5 1 1 25577
0 25579 7 1 2 25574 25578
0 25580 5 1 1 25579
0 25581 7 1 2 46515 25580
0 25582 5 1 1 25581
0 25583 7 1 2 68856 69491
0 25584 7 1 2 69004 25583
0 25585 5 1 1 25584
0 25586 7 1 2 25582 25585
0 25587 5 1 1 25586
0 25588 7 1 2 43474 25587
0 25589 5 1 1 25588
0 25590 7 2 2 52683 69449
0 25591 7 1 2 58281 68384
0 25592 7 1 2 69494 25591
0 25593 5 1 1 25592
0 25594 7 1 2 25589 25593
0 25595 5 1 1 25594
0 25596 7 1 2 42043 25595
0 25597 5 1 1 25596
0 25598 7 1 2 61860 66041
0 25599 7 1 2 69495 25598
0 25600 5 1 1 25599
0 25601 7 1 2 25597 25600
0 25602 5 1 1 25601
0 25603 7 1 2 62128 64401
0 25604 7 1 2 25602 25603
0 25605 5 1 1 25604
0 25606 7 1 2 25562 25605
0 25607 5 1 1 25606
0 25608 7 1 2 49225 25607
0 25609 5 1 1 25608
0 25610 7 1 2 65292 69438
0 25611 5 1 1 25610
0 25612 7 3 2 64048 66634
0 25613 5 1 1 69496
0 25614 7 1 2 45466 65023
0 25615 7 1 2 69497 25614
0 25616 5 1 1 25615
0 25617 7 1 2 25611 25616
0 25618 5 1 1 25617
0 25619 7 1 2 49295 25618
0 25620 5 1 1 25619
0 25621 7 1 2 50194 58360
0 25622 5 1 1 25621
0 25623 7 1 2 49532 25622
0 25624 5 1 1 25623
0 25625 7 1 2 52590 65908
0 25626 7 1 2 25624 25625
0 25627 5 1 1 25626
0 25628 7 1 2 25620 25627
0 25629 5 1 1 25628
0 25630 7 1 2 69468 25629
0 25631 5 1 1 25630
0 25632 7 1 2 48275 25631
0 25633 7 1 2 25609 25632
0 25634 7 1 2 25554 25633
0 25635 5 1 1 25634
0 25636 7 2 2 43114 57900
0 25637 5 1 1 69499
0 25638 7 1 2 19852 25637
0 25639 5 1 1 25638
0 25640 7 1 2 44080 25639
0 25641 5 1 1 25640
0 25642 7 1 2 57582 8932
0 25643 5 1 1 25642
0 25644 7 2 2 47308 62369
0 25645 5 1 1 69501
0 25646 7 1 2 46516 25645
0 25647 7 2 2 25643 25646
0 25648 5 1 1 69503
0 25649 7 1 2 25641 25648
0 25650 5 1 1 25649
0 25651 7 1 2 45109 25650
0 25652 5 1 1 25651
0 25653 7 3 2 46060 52638
0 25654 7 1 2 46716 69505
0 25655 5 1 1 25654
0 25656 7 1 2 25652 25655
0 25657 5 1 1 25656
0 25658 7 1 2 48631 25657
0 25659 5 1 1 25658
0 25660 7 1 2 46061 49442
0 25661 5 1 1 25660
0 25662 7 1 2 781 52758
0 25663 5 1 1 25662
0 25664 7 1 2 51401 52639
0 25665 7 1 2 25663 25664
0 25666 5 1 1 25665
0 25667 7 1 2 25661 25666
0 25668 5 1 1 25667
0 25669 7 1 2 46717 25668
0 25670 5 1 1 25669
0 25671 7 1 2 25659 25670
0 25672 5 1 1 25671
0 25673 7 1 2 69444 25672
0 25674 5 1 1 25673
0 25675 7 1 2 45110 57551
0 25676 5 1 1 25675
0 25677 7 1 2 56331 25676
0 25678 5 2 1 25677
0 25679 7 1 2 60749 69474
0 25680 7 1 2 69508 25679
0 25681 5 1 1 25680
0 25682 7 1 2 25674 25681
0 25683 5 1 1 25682
0 25684 7 1 2 44243 25683
0 25685 5 1 1 25684
0 25686 7 3 2 67938 69280
0 25687 7 1 2 48979 69510
0 25688 5 1 1 25687
0 25689 7 1 2 51444 68607
0 25690 7 1 2 68894 25689
0 25691 5 1 1 25690
0 25692 7 1 2 25688 25691
0 25693 5 1 1 25692
0 25694 7 1 2 44081 25693
0 25695 5 1 1 25694
0 25696 7 1 2 52387 69511
0 25697 5 1 1 25696
0 25698 7 1 2 25695 25697
0 25699 5 1 1 25698
0 25700 7 1 2 69506 25699
0 25701 5 1 1 25700
0 25702 7 2 2 47567 50615
0 25703 5 1 1 69513
0 25704 7 1 2 52640 69514
0 25705 7 1 2 69475 25704
0 25706 5 1 1 25705
0 25707 7 1 2 53056 57327
0 25708 7 1 2 64132 25707
0 25709 7 1 2 69512 25708
0 25710 5 1 1 25709
0 25711 7 1 2 45467 25710
0 25712 7 1 2 25706 25711
0 25713 5 1 1 25712
0 25714 7 1 2 50245 3053
0 25715 5 1 1 25714
0 25716 7 1 2 49897 68895
0 25717 7 1 2 25715 25716
0 25718 5 1 1 25717
0 25719 7 1 2 57952 66067
0 25720 7 1 2 50240 25719
0 25721 7 1 2 69493 25720
0 25722 5 1 1 25721
0 25723 7 1 2 48820 25722
0 25724 7 1 2 25718 25723
0 25725 5 1 1 25724
0 25726 7 1 2 43115 25725
0 25727 7 1 2 25713 25726
0 25728 5 1 1 25727
0 25729 7 1 2 25701 25728
0 25730 7 1 2 25685 25729
0 25731 5 1 1 25730
0 25732 7 1 2 42327 25731
0 25733 5 1 1 25732
0 25734 7 1 2 51765 69509
0 25735 5 1 1 25734
0 25736 7 1 2 49176 69316
0 25737 5 1 1 25736
0 25738 7 1 2 25735 25737
0 25739 5 2 1 25738
0 25740 7 1 2 66264 68468
0 25741 7 1 2 69515 25740
0 25742 5 1 1 25741
0 25743 7 1 2 25733 25742
0 25744 5 1 1 25743
0 25745 7 1 2 42217 25744
0 25746 5 1 1 25745
0 25747 7 1 2 42328 67018
0 25748 5 1 1 25747
0 25749 7 1 2 66265 68417
0 25750 5 1 1 25749
0 25751 7 1 2 25748 25750
0 25752 5 3 1 25751
0 25753 7 1 2 47784 60795
0 25754 7 1 2 69517 25753
0 25755 7 1 2 69516 25754
0 25756 5 1 1 25755
0 25757 7 1 2 25746 25756
0 25758 5 1 1 25757
0 25759 7 1 2 42849 25758
0 25760 5 1 1 25759
0 25761 7 2 2 51766 65024
0 25762 5 2 1 69520
0 25763 7 1 2 48465 53826
0 25764 5 1 1 25763
0 25765 7 1 2 69522 25764
0 25766 5 1 1 25765
0 25767 7 1 2 46517 25766
0 25768 5 1 1 25767
0 25769 7 1 2 49405 69523
0 25770 5 1 1 25769
0 25771 7 1 2 47441 25770
0 25772 5 1 1 25771
0 25773 7 1 2 25768 25772
0 25774 5 2 1 25773
0 25775 7 1 2 64114 68896
0 25776 5 1 1 25775
0 25777 7 1 2 66266 67691
0 25778 5 1 1 25777
0 25779 7 1 2 25776 25778
0 25780 5 1 1 25779
0 25781 7 1 2 69524 25780
0 25782 5 1 1 25781
0 25783 7 1 2 46282 51445
0 25784 7 1 2 68731 25783
0 25785 5 1 1 25784
0 25786 7 1 2 46718 25785
0 25787 5 1 1 25786
0 25788 7 1 2 65346 25787
0 25789 5 1 1 25788
0 25790 7 1 2 45111 25789
0 25791 5 1 1 25790
0 25792 7 1 2 68902 25791
0 25793 5 1 1 25792
0 25794 7 1 2 47309 25793
0 25795 5 1 1 25794
0 25796 7 1 2 68900 25795
0 25797 5 1 1 25796
0 25798 7 3 2 63343 66193
0 25799 7 1 2 44467 69526
0 25800 7 1 2 25797 25799
0 25801 5 1 1 25800
0 25802 7 1 2 25782 25801
0 25803 5 1 1 25802
0 25804 7 1 2 42218 25803
0 25805 5 1 1 25804
0 25806 7 1 2 47785 61637
0 25807 7 1 2 69518 25806
0 25808 7 1 2 69525 25807
0 25809 5 1 1 25808
0 25810 7 1 2 25805 25809
0 25811 5 1 1 25810
0 25812 7 1 2 42586 25811
0 25813 5 1 1 25812
0 25814 7 1 2 44680 25813
0 25815 7 1 2 25760 25814
0 25816 5 1 1 25815
0 25817 7 2 2 60088 61529
0 25818 5 1 1 69529
0 25819 7 1 2 3416 25818
0 25820 5 1 1 25819
0 25821 7 1 2 68852 25820
0 25822 5 1 1 25821
0 25823 7 1 2 52641 62394
0 25824 5 1 1 25823
0 25825 7 1 2 50241 63494
0 25826 5 1 1 25825
0 25827 7 1 2 25824 25826
0 25828 5 1 1 25827
0 25829 7 1 2 46062 62419
0 25830 7 1 2 25828 25829
0 25831 5 1 1 25830
0 25832 7 1 2 25822 25831
0 25833 5 3 1 25832
0 25834 7 4 2 63077 65855
0 25835 7 1 2 65426 69534
0 25836 7 1 2 69531 25835
0 25837 5 1 1 25836
0 25838 7 1 2 49758 65293
0 25839 5 1 1 25838
0 25840 7 1 2 68898 25839
0 25841 5 1 1 25840
0 25842 7 1 2 42587 25841
0 25843 5 1 1 25842
0 25844 7 1 2 49517 56781
0 25845 7 1 2 50251 25844
0 25846 5 1 1 25845
0 25847 7 1 2 25843 25846
0 25848 5 1 1 25847
0 25849 7 1 2 46283 25848
0 25850 5 1 1 25849
0 25851 7 1 2 64202 64877
0 25852 5 1 1 25851
0 25853 7 1 2 52187 54183
0 25854 5 1 1 25853
0 25855 7 1 2 62424 25854
0 25856 5 1 1 25855
0 25857 7 1 2 46719 53817
0 25858 7 1 2 64900 25857
0 25859 7 1 2 25856 25858
0 25860 5 1 1 25859
0 25861 7 1 2 25852 25860
0 25862 5 1 1 25861
0 25863 7 1 2 46063 25862
0 25864 5 1 1 25863
0 25865 7 1 2 25850 25864
0 25866 5 1 1 25865
0 25867 7 1 2 55848 68161
0 25868 7 1 2 25866 25867
0 25869 5 1 1 25868
0 25870 7 1 2 25837 25869
0 25871 5 1 1 25870
0 25872 7 1 2 42219 25871
0 25873 5 1 1 25872
0 25874 7 1 2 46937 68158
0 25875 5 1 1 25874
0 25876 7 1 2 43552 17306
0 25877 5 1 1 25876
0 25878 7 1 2 55976 25877
0 25879 7 1 2 25875 25878
0 25880 7 1 2 69532 25879
0 25881 5 1 1 25880
0 25882 7 1 2 48015 25881
0 25883 7 1 2 25873 25882
0 25884 5 1 1 25883
0 25885 7 1 2 48907 25884
0 25886 7 1 2 25816 25885
0 25887 5 1 1 25886
0 25888 7 4 2 42588 51011
0 25889 7 4 2 46284 69538
0 25890 7 1 2 53142 69542
0 25891 5 1 1 25890
0 25892 7 1 2 54398 54690
0 25893 5 1 1 25892
0 25894 7 1 2 25891 25893
0 25895 5 1 1 25894
0 25896 7 1 2 48632 25895
0 25897 5 1 1 25896
0 25898 7 1 2 54390 56328
0 25899 5 1 1 25898
0 25900 7 1 2 25897 25899
0 25901 5 1 1 25900
0 25902 7 1 2 51767 25901
0 25903 5 1 1 25902
0 25904 7 2 2 49177 51072
0 25905 5 1 1 69546
0 25906 7 1 2 56620 69547
0 25907 5 1 1 25906
0 25908 7 3 2 52927 69543
0 25909 5 1 1 69548
0 25910 7 1 2 52098 54391
0 25911 5 1 1 25910
0 25912 7 1 2 25909 25911
0 25913 5 1 1 25912
0 25914 7 1 2 49178 25913
0 25915 5 1 1 25914
0 25916 7 1 2 46518 68684
0 25917 5 1 1 25916
0 25918 7 1 2 25915 25917
0 25919 5 1 1 25918
0 25920 7 1 2 48466 25919
0 25921 5 1 1 25920
0 25922 7 1 2 25907 25921
0 25923 7 1 2 25903 25922
0 25924 5 1 1 25923
0 25925 7 1 2 67541 25924
0 25926 5 1 1 25925
0 25927 7 3 2 48016 69533
0 25928 7 1 2 46992 69551
0 25929 5 1 1 25928
0 25930 7 1 2 25926 25929
0 25931 5 1 1 25930
0 25932 7 1 2 66382 25931
0 25933 5 1 1 25932
0 25934 7 1 2 66246 69552
0 25935 5 1 1 25934
0 25936 7 1 2 25933 25935
0 25937 5 1 1 25936
0 25938 7 1 2 42329 25937
0 25939 5 1 1 25938
0 25940 7 1 2 68156 69553
0 25941 5 1 1 25940
0 25942 7 1 2 25939 25941
0 25943 5 1 1 25942
0 25944 7 1 2 47786 69272
0 25945 7 1 2 25943 25944
0 25946 5 1 1 25945
0 25947 7 1 2 44941 25946
0 25948 7 1 2 25887 25947
0 25949 5 1 1 25948
0 25950 7 1 2 25635 25949
0 25951 5 1 1 25950
0 25952 7 12 2 42330 48017
0 25953 5 3 1 69554
0 25954 7 2 2 58753 69555
0 25955 7 2 2 46064 69569
0 25956 7 1 2 15303 68911
0 25957 5 1 1 25956
0 25958 7 1 2 46720 25957
0 25959 5 1 1 25958
0 25960 7 1 2 47442 57387
0 25961 7 1 2 65115 25960
0 25962 5 1 1 25961
0 25963 7 1 2 49004 52591
0 25964 5 2 1 25963
0 25965 7 1 2 44244 69573
0 25966 7 1 2 25962 25965
0 25967 5 1 1 25966
0 25968 7 3 2 50227 62163
0 25969 5 2 1 69575
0 25970 7 1 2 47568 69578
0 25971 5 1 1 25970
0 25972 7 1 2 43336 25971
0 25973 7 1 2 25967 25972
0 25974 5 1 1 25973
0 25975 7 1 2 25959 25974
0 25976 5 1 1 25975
0 25977 7 1 2 69571 25976
0 25978 5 1 1 25977
0 25979 7 1 2 52592 68907
0 25980 5 1 1 25979
0 25981 7 1 2 25511 25980
0 25982 5 2 1 25981
0 25983 7 1 2 56546 69580
0 25984 5 1 1 25983
0 25985 7 1 2 43337 69574
0 25986 7 1 2 23077 25985
0 25987 5 1 1 25986
0 25988 7 1 2 46721 69579
0 25989 5 1 1 25988
0 25990 7 1 2 57774 61037
0 25991 7 1 2 25989 25990
0 25992 7 1 2 25987 25991
0 25993 5 1 1 25992
0 25994 7 1 2 25984 25993
0 25995 5 1 1 25994
0 25996 7 1 2 47443 25995
0 25997 5 1 1 25996
0 25998 7 2 2 45112 56252
0 25999 7 1 2 63275 64751
0 26000 7 1 2 56763 25999
0 26001 7 1 2 69582 26000
0 26002 5 1 1 26001
0 26003 7 1 2 25997 26002
0 26004 5 1 1 26003
0 26005 7 1 2 69556 26004
0 26006 5 1 1 26005
0 26007 7 1 2 51446 68857
0 26008 7 1 2 55030 26007
0 26009 7 1 2 69080 26008
0 26010 5 1 1 26009
0 26011 7 1 2 26006 26010
0 26012 5 1 1 26011
0 26013 7 1 2 46519 26012
0 26014 5 1 1 26013
0 26015 7 1 2 68863 69572
0 26016 5 1 1 26015
0 26017 7 1 2 46065 69521
0 26018 5 1 1 26017
0 26019 7 1 2 55031 57390
0 26020 5 1 1 26019
0 26021 7 1 2 26018 26020
0 26022 5 1 1 26021
0 26023 7 1 2 69081 26022
0 26024 5 1 1 26023
0 26025 7 2 2 45760 58399
0 26026 7 1 2 48018 49384
0 26027 7 1 2 55744 66462
0 26028 7 1 2 26026 26027
0 26029 7 1 2 69584 26028
0 26030 5 1 1 26029
0 26031 7 1 2 26024 26030
0 26032 5 1 1 26031
0 26033 7 1 2 47787 26032
0 26034 5 1 1 26033
0 26035 7 1 2 26016 26034
0 26036 5 1 1 26035
0 26037 7 1 2 51012 26036
0 26038 5 1 1 26037
0 26039 7 1 2 55022 62291
0 26040 5 1 1 26039
0 26041 7 1 2 46066 55252
0 26042 5 1 1 26041
0 26043 7 1 2 26040 26042
0 26044 5 1 1 26043
0 26045 7 1 2 46722 26044
0 26046 5 1 1 26045
0 26047 7 1 2 49898 69442
0 26048 5 1 1 26047
0 26049 7 1 2 26046 26048
0 26050 5 1 1 26049
0 26051 7 1 2 45275 26050
0 26052 5 1 1 26051
0 26053 7 2 2 49179 49807
0 26054 7 1 2 58460 69586
0 26055 5 1 1 26054
0 26056 7 1 2 26052 26055
0 26057 5 1 1 26056
0 26058 7 1 2 69570 26057
0 26059 5 1 1 26058
0 26060 7 1 2 26038 26059
0 26061 7 1 2 26014 26060
0 26062 5 1 1 26061
0 26063 7 1 2 46285 26062
0 26064 5 1 1 26063
0 26065 7 1 2 25978 26064
0 26066 5 1 1 26065
0 26067 7 1 2 43475 26066
0 26068 5 1 1 26067
0 26069 7 1 2 49296 69581
0 26070 5 1 1 26069
0 26071 7 1 2 16692 26070
0 26072 5 1 1 26071
0 26073 7 3 2 47788 51013
0 26074 7 1 2 51887 69588
0 26075 7 2 2 26072 26074
0 26076 7 1 2 60966 63830
0 26077 7 1 2 69591 26076
0 26078 5 1 1 26077
0 26079 7 1 2 26068 26078
0 26080 5 1 1 26079
0 26081 7 1 2 42044 26080
0 26082 5 1 1 26081
0 26083 7 1 2 64445 66671
0 26084 7 1 2 69592 26083
0 26085 5 1 1 26084
0 26086 7 1 2 26082 26085
0 26087 5 1 1 26086
0 26088 7 1 2 48276 26087
0 26089 5 1 1 26088
0 26090 7 1 2 51888 58872
0 26091 7 1 2 69576 26090
0 26092 7 2 2 56040 63400
0 26093 7 1 2 69593 69489
0 26094 7 1 2 26091 26093
0 26095 5 1 1 26094
0 26096 7 1 2 26089 26095
0 26097 5 1 1 26096
0 26098 7 1 2 66267 26097
0 26099 5 1 1 26098
0 26100 7 1 2 49297 57916
0 26101 7 1 2 67814 26100
0 26102 7 1 2 56375 65125
0 26103 7 4 2 55411 64686
0 26104 7 1 2 67122 69595
0 26105 7 1 2 26102 26104
0 26106 7 1 2 26101 26105
0 26107 5 1 1 26106
0 26108 7 1 2 44343 26107
0 26109 7 1 2 26099 26108
0 26110 7 1 2 25951 26109
0 26111 5 1 1 26110
0 26112 7 2 2 51014 55480
0 26113 5 1 1 69599
0 26114 7 1 2 50186 26113
0 26115 5 1 1 26114
0 26116 7 1 2 59510 26115
0 26117 5 1 1 26116
0 26118 7 1 2 47569 26117
0 26119 5 1 1 26118
0 26120 7 1 2 50858 57840
0 26121 5 1 1 26120
0 26122 7 1 2 45276 60874
0 26123 7 1 2 26121 26122
0 26124 5 1 1 26123
0 26125 7 1 2 52928 26124
0 26126 5 1 1 26125
0 26127 7 1 2 26119 26126
0 26128 5 1 1 26127
0 26129 7 1 2 49657 26128
0 26130 5 1 1 26129
0 26131 7 1 2 58634 62955
0 26132 5 1 1 26131
0 26133 7 1 2 26130 26132
0 26134 5 1 1 26133
0 26135 7 1 2 43932 26134
0 26136 5 1 1 26135
0 26137 7 1 2 46723 23487
0 26138 5 1 1 26137
0 26139 7 1 2 23499 26138
0 26140 5 1 1 26139
0 26141 7 1 2 48467 26140
0 26142 5 1 1 26141
0 26143 7 1 2 50228 60818
0 26144 5 1 1 26143
0 26145 7 1 2 26142 26144
0 26146 5 1 1 26145
0 26147 7 1 2 54728 26146
0 26148 5 1 1 26147
0 26149 7 1 2 26136 26148
0 26150 5 1 1 26149
0 26151 7 1 2 46286 26150
0 26152 5 1 1 26151
0 26153 7 1 2 49835 56782
0 26154 5 1 1 26153
0 26155 7 1 2 54729 60029
0 26156 5 1 1 26155
0 26157 7 1 2 26154 26156
0 26158 5 1 1 26157
0 26159 7 1 2 47570 26158
0 26160 5 1 1 26159
0 26161 7 1 2 54733 56900
0 26162 7 1 2 64133 26161
0 26163 5 1 1 26162
0 26164 7 1 2 26160 26163
0 26165 5 1 1 26164
0 26166 7 1 2 46520 26165
0 26167 5 1 1 26166
0 26168 7 1 2 53758 58387
0 26169 5 1 1 26168
0 26170 7 1 2 45468 62885
0 26171 5 1 1 26170
0 26172 7 1 2 26169 26171
0 26173 5 1 1 26172
0 26174 7 1 2 52593 57291
0 26175 7 1 2 26173 26174
0 26176 5 1 1 26175
0 26177 7 1 2 26167 26176
0 26178 5 1 1 26177
0 26179 7 1 2 42850 26178
0 26180 5 1 1 26179
0 26181 7 1 2 26152 26180
0 26182 5 2 1 26181
0 26183 7 1 2 69082 69601
0 26184 5 1 1 26183
0 26185 7 5 2 48277 49385
0 26186 5 1 1 69603
0 26187 7 1 2 57053 62335
0 26188 7 1 2 69604 26187
0 26189 7 1 2 66467 26188
0 26190 5 1 1 26189
0 26191 7 1 2 26184 26190
0 26192 5 1 1 26191
0 26193 7 1 2 66268 26192
0 26194 5 1 1 26193
0 26195 7 1 2 65700 69602
0 26196 5 1 1 26195
0 26197 7 2 2 53745 57414
0 26198 5 1 1 69608
0 26199 7 2 2 49817 65909
0 26200 7 1 2 54705 69610
0 26201 7 1 2 69609 26200
0 26202 5 1 1 26201
0 26203 7 1 2 26196 26202
0 26204 5 1 1 26203
0 26205 7 1 2 69005 26204
0 26206 5 1 1 26205
0 26207 7 1 2 26194 26206
0 26208 5 1 1 26207
0 26209 7 1 2 58198 58980
0 26210 7 1 2 26208 26209
0 26211 5 1 1 26210
0 26212 7 1 2 56751 69042
0 26213 5 1 1 26212
0 26214 7 1 2 54330 69021
0 26215 5 1 1 26214
0 26216 7 1 2 26213 26215
0 26217 5 1 1 26216
0 26218 7 1 2 50332 26217
0 26219 5 1 1 26218
0 26220 7 1 2 62441 69022
0 26221 5 1 1 26220
0 26222 7 1 2 26219 26221
0 26223 5 1 1 26222
0 26224 7 1 2 46521 26223
0 26225 5 1 1 26224
0 26226 7 1 2 54730 57391
0 26227 5 1 1 26226
0 26228 7 1 2 49542 57399
0 26229 5 1 1 26228
0 26230 7 1 2 26227 26229
0 26231 5 1 1 26230
0 26232 7 1 2 43116 26231
0 26233 5 1 1 26232
0 26234 7 1 2 49879 58313
0 26235 5 1 1 26234
0 26236 7 1 2 49818 50859
0 26237 7 1 2 52753 26236
0 26238 5 1 1 26237
0 26239 7 1 2 26235 26238
0 26240 5 1 1 26239
0 26241 7 1 2 48821 26240
0 26242 5 1 1 26241
0 26243 7 1 2 26233 26242
0 26244 5 1 1 26243
0 26245 7 1 2 46067 26244
0 26246 5 1 1 26245
0 26247 7 1 2 26225 26246
0 26248 5 1 1 26247
0 26249 7 1 2 48468 26248
0 26250 5 1 1 26249
0 26251 7 1 2 47571 62886
0 26252 5 1 1 26251
0 26253 7 1 2 52818 26252
0 26254 5 1 1 26253
0 26255 7 1 2 57054 26254
0 26256 5 1 1 26255
0 26257 7 1 2 51210 52920
0 26258 5 1 1 26257
0 26259 7 1 2 65446 26258
0 26260 5 1 1 26259
0 26261 7 1 2 47310 26260
0 26262 5 1 1 26261
0 26263 7 1 2 26256 26262
0 26264 5 1 1 26263
0 26265 7 1 2 46068 26264
0 26266 5 1 1 26265
0 26267 7 1 2 48969 64333
0 26268 5 1 1 26267
0 26269 7 1 2 26266 26268
0 26270 5 1 1 26269
0 26271 7 1 2 49658 26270
0 26272 5 1 1 26271
0 26273 7 1 2 26250 26272
0 26274 5 1 1 26273
0 26275 7 1 2 42331 68298
0 26276 7 1 2 26274 26275
0 26277 5 1 1 26276
0 26278 7 1 2 58246 68936
0 26279 5 1 1 26278
0 26280 7 1 2 48278 69018
0 26281 5 1 1 26280
0 26282 7 1 2 26279 26281
0 26283 5 1 1 26282
0 26284 7 1 2 49298 26283
0 26285 5 1 1 26284
0 26286 7 1 2 51015 65565
0 26287 7 1 2 69605 26286
0 26288 5 1 1 26287
0 26289 7 1 2 26285 26288
0 26290 5 1 1 26289
0 26291 7 2 2 56283 69071
0 26292 7 1 2 45469 69612
0 26293 7 1 2 26290 26292
0 26294 5 1 1 26293
0 26295 7 1 2 26277 26294
0 26296 5 1 1 26295
0 26297 7 1 2 66269 26296
0 26298 5 1 1 26297
0 26299 7 1 2 54789 69006
0 26300 5 2 1 26299
0 26301 7 1 2 67123 67767
0 26302 5 1 1 26301
0 26303 7 1 2 69614 26302
0 26304 5 1 1 26303
0 26305 7 1 2 51426 54734
0 26306 5 1 1 26305
0 26307 7 2 2 43933 53469
0 26308 5 1 1 69616
0 26309 7 1 2 68958 69617
0 26310 5 1 1 26309
0 26311 7 1 2 26306 26310
0 26312 5 1 1 26311
0 26313 7 1 2 43338 26312
0 26314 5 1 1 26313
0 26315 7 1 2 56626 56804
0 26316 5 1 1 26315
0 26317 7 1 2 26314 26316
0 26318 5 1 1 26317
0 26319 7 1 2 49345 26318
0 26320 5 1 1 26319
0 26321 7 1 2 49406 65130
0 26322 5 1 1 26321
0 26323 7 1 2 43117 26322
0 26324 5 1 1 26323
0 26325 7 1 2 49386 62404
0 26326 5 1 1 26325
0 26327 7 1 2 26324 26326
0 26328 5 1 1 26327
0 26329 7 1 2 47311 26328
0 26330 5 1 1 26329
0 26331 7 1 2 50234 69168
0 26332 5 2 1 26331
0 26333 7 1 2 56705 69618
0 26334 5 1 1 26333
0 26335 7 1 2 53100 26334
0 26336 5 1 1 26335
0 26337 7 1 2 57055 26336
0 26338 5 1 1 26337
0 26339 7 1 2 26330 26338
0 26340 5 1 1 26339
0 26341 7 1 2 48279 26340
0 26342 5 1 1 26341
0 26343 7 1 2 26320 26342
0 26344 5 1 1 26343
0 26345 7 1 2 65910 26344
0 26346 5 1 1 26345
0 26347 7 1 2 55655 69216
0 26348 7 1 2 57673 26347
0 26349 5 1 1 26348
0 26350 7 1 2 26346 26349
0 26351 5 1 1 26350
0 26352 7 1 2 46069 26351
0 26353 5 1 1 26352
0 26354 7 1 2 49819 52594
0 26355 5 1 1 26354
0 26356 7 1 2 44942 68937
0 26357 5 1 1 26356
0 26358 7 1 2 26355 26357
0 26359 5 1 1 26358
0 26360 7 1 2 66001 26359
0 26361 5 1 1 26360
0 26362 7 1 2 23856 26361
0 26363 5 1 1 26362
0 26364 7 1 2 42589 61695
0 26365 7 1 2 26363 26364
0 26366 5 1 1 26365
0 26367 7 1 2 26353 26366
0 26368 5 1 1 26367
0 26369 7 1 2 26304 26368
0 26370 5 1 1 26369
0 26371 7 1 2 26298 26370
0 26372 5 1 1 26371
0 26373 7 1 2 46287 26372
0 26374 5 1 1 26373
0 26375 7 2 2 49602 60809
0 26376 5 1 1 69620
0 26377 7 1 2 52762 57292
0 26378 5 1 1 26377
0 26379 7 1 2 26376 26378
0 26380 5 1 1 26379
0 26381 7 1 2 53777 26380
0 26382 5 1 1 26381
0 26383 7 1 2 49659 62202
0 26384 7 1 2 49887 26383
0 26385 5 1 1 26384
0 26386 7 1 2 26382 26385
0 26387 5 1 1 26386
0 26388 7 1 2 45277 26387
0 26389 5 1 1 26388
0 26390 7 1 2 49836 63690
0 26391 5 1 1 26390
0 26392 7 1 2 49660 58663
0 26393 5 1 1 26392
0 26394 7 1 2 23706 26393
0 26395 5 1 1 26394
0 26396 7 1 2 45278 26395
0 26397 5 1 1 26396
0 26398 7 1 2 26391 26397
0 26399 5 1 1 26398
0 26400 7 1 2 43934 26399
0 26401 5 1 1 26400
0 26402 7 1 2 52564 58901
0 26403 7 1 2 65029 26402
0 26404 5 1 1 26403
0 26405 7 1 2 26401 26404
0 26406 7 1 2 26389 26405
0 26407 5 1 1 26406
0 26408 7 1 2 45470 26407
0 26409 5 1 1 26408
0 26410 7 2 2 48822 57841
0 26411 7 1 2 54606 69622
0 26412 5 1 1 26411
0 26413 7 2 2 48280 52671
0 26414 7 1 2 55526 69624
0 26415 5 1 1 26414
0 26416 7 1 2 26412 26415
0 26417 5 1 1 26416
0 26418 7 1 2 45279 26417
0 26419 5 1 1 26418
0 26420 7 1 2 54692 64888
0 26421 5 1 1 26420
0 26422 7 1 2 43118 26421
0 26423 5 1 1 26422
0 26424 7 1 2 49443 62164
0 26425 5 1 1 26424
0 26426 7 1 2 26423 26425
0 26427 5 1 1 26426
0 26428 7 1 2 54830 26427
0 26429 5 1 1 26428
0 26430 7 1 2 26419 26429
0 26431 5 1 1 26430
0 26432 7 1 2 49997 26431
0 26433 5 1 1 26432
0 26434 7 1 2 50860 67788
0 26435 7 1 2 68677 26434
0 26436 5 1 1 26435
0 26437 7 1 2 26433 26436
0 26438 7 1 2 26409 26437
0 26439 5 1 1 26438
0 26440 7 1 2 56284 66342
0 26441 5 1 1 26440
0 26442 7 1 2 58136 68162
0 26443 5 1 1 26442
0 26444 7 1 2 26441 26443
0 26445 5 1 1 26444
0 26446 7 1 2 61876 26445
0 26447 7 1 2 26439 26446
0 26448 5 1 1 26447
0 26449 7 1 2 26374 26448
0 26450 5 1 1 26449
0 26451 7 1 2 44468 26450
0 26452 5 1 1 26451
0 26453 7 1 2 47673 26452
0 26454 7 1 2 26211 26453
0 26455 5 1 1 26454
0 26456 7 1 2 48132 26455
0 26457 7 1 2 26111 26456
0 26458 5 1 1 26457
0 26459 7 1 2 44590 26458
0 26460 7 1 2 25354 26459
0 26461 5 1 1 26460
0 26462 7 2 2 59205 68815
0 26463 7 1 2 67848 69626
0 26464 5 1 1 26463
0 26465 7 2 2 45761 66214
0 26466 7 2 2 66716 69628
0 26467 7 2 2 66648 69630
0 26468 7 2 2 44245 64502
0 26469 7 2 2 54638 69634
0 26470 7 1 2 69632 69636
0 26471 5 1 1 26470
0 26472 7 1 2 26464 26471
0 26473 5 1 1 26472
0 26474 7 1 2 45280 26473
0 26475 5 1 1 26474
0 26476 7 1 2 49005 51270
0 26477 7 2 2 69635 26476
0 26478 7 1 2 69633 69638
0 26479 5 1 1 26478
0 26480 7 1 2 26475 26479
0 26481 5 1 1 26480
0 26482 7 1 2 45603 26481
0 26483 5 1 1 26482
0 26484 7 1 2 46851 68816
0 26485 5 1 1 26484
0 26486 7 2 2 46938 66177
0 26487 5 1 1 69640
0 26488 7 1 2 26485 26487
0 26489 5 3 1 26488
0 26490 7 2 2 49568 51251
0 26491 7 1 2 59368 69645
0 26492 7 1 2 69642 26491
0 26493 5 1 1 26492
0 26494 7 1 2 26483 26493
0 26495 5 1 1 26494
0 26496 7 1 2 64328 26495
0 26497 5 1 1 26496
0 26498 7 2 2 48469 53528
0 26499 7 1 2 44082 54298
0 26500 5 1 1 26499
0 26501 7 1 2 53449 26500
0 26502 5 2 1 26501
0 26503 7 1 2 68825 69649
0 26504 5 1 1 26503
0 26505 7 1 2 50276 58842
0 26506 7 1 2 61823 26505
0 26507 7 1 2 64044 66165
0 26508 7 1 2 26506 26507
0 26509 5 1 1 26508
0 26510 7 1 2 26504 26509
0 26511 5 1 1 26510
0 26512 7 1 2 69647 26511
0 26513 5 1 1 26512
0 26514 7 1 2 49395 64884
0 26515 5 1 1 26514
0 26516 7 1 2 43339 26515
0 26517 5 1 1 26516
0 26518 7 1 2 52811 54301
0 26519 5 1 1 26518
0 26520 7 1 2 48470 26519
0 26521 5 1 1 26520
0 26522 7 1 2 26517 26521
0 26523 5 1 1 26522
0 26524 7 1 2 50953 26523
0 26525 5 1 1 26524
0 26526 7 1 2 55474 68938
0 26527 5 1 1 26526
0 26528 7 2 2 26525 26527
0 26529 5 1 1 69651
0 26530 7 1 2 68826 26529
0 26531 5 1 1 26530
0 26532 7 1 2 52214 1482
0 26533 7 1 2 14077 26532
0 26534 5 1 1 26533
0 26535 7 3 2 60130 26534
0 26536 7 1 2 69643 69653
0 26537 5 1 1 26536
0 26538 7 1 2 42045 26537
0 26539 5 1 1 26538
0 26540 7 1 2 45762 67092
0 26541 5 1 1 26540
0 26542 7 2 2 53687 67019
0 26543 5 1 1 69656
0 26544 7 1 2 26541 26543
0 26545 5 1 1 26544
0 26546 7 1 2 69654 26545
0 26547 5 1 1 26546
0 26548 7 1 2 50235 4406
0 26549 5 1 1 26548
0 26550 7 1 2 52676 10583
0 26551 7 2 2 26549 26550
0 26552 7 1 2 47674 49226
0 26553 7 2 2 69658 26552
0 26554 7 1 2 45763 66912
0 26555 7 1 2 69660 26554
0 26556 5 1 1 26555
0 26557 7 1 2 45604 26556
0 26558 7 1 2 26547 26557
0 26559 5 1 1 26558
0 26560 7 1 2 46724 26559
0 26561 7 1 2 26539 26560
0 26562 5 1 1 26561
0 26563 7 1 2 42046 69641
0 26564 5 1 1 26563
0 26565 7 1 2 68821 26564
0 26566 5 2 1 26565
0 26567 7 2 2 49346 53340
0 26568 5 1 1 69664
0 26569 7 2 2 52808 69665
0 26570 5 1 1 69666
0 26571 7 1 2 69662 69667
0 26572 5 1 1 26571
0 26573 7 2 2 52677 6904
0 26574 5 1 1 69668
0 26575 7 1 2 68823 69669
0 26576 5 1 1 26575
0 26577 7 1 2 26572 26576
0 26578 5 1 1 26577
0 26579 7 1 2 44344 26578
0 26580 5 1 1 26579
0 26581 7 1 2 45113 59575
0 26582 7 1 2 53152 26581
0 26583 7 1 2 66166 68018
0 26584 7 1 2 26582 26583
0 26585 5 1 1 26584
0 26586 7 1 2 26580 26585
0 26587 7 1 2 26562 26586
0 26588 5 1 1 26587
0 26589 7 1 2 43935 26588
0 26590 5 1 1 26589
0 26591 7 1 2 26531 26590
0 26592 5 1 1 26591
0 26593 7 1 2 42851 26592
0 26594 5 1 1 26593
0 26595 7 1 2 26513 26594
0 26596 5 1 1 26595
0 26597 7 1 2 44812 26596
0 26598 5 1 1 26597
0 26599 7 2 2 46725 61560
0 26600 7 1 2 54576 69670
0 26601 7 2 2 53837 26600
0 26602 7 1 2 69663 69672
0 26603 5 1 1 26602
0 26604 7 1 2 48281 26603
0 26605 7 1 2 26598 26604
0 26606 5 1 1 26605
0 26607 7 1 2 69052 22916
0 26608 5 1 1 26607
0 26609 7 2 2 46522 26608
0 26610 5 1 1 69674
0 26611 7 1 2 53324 26610
0 26612 5 1 1 26611
0 26613 7 1 2 48471 26612
0 26614 5 1 1 26613
0 26615 7 1 2 68755 26614
0 26616 5 1 1 26615
0 26617 7 1 2 47444 26616
0 26618 5 1 1 26617
0 26619 7 1 2 49387 58664
0 26620 5 1 1 26619
0 26621 7 1 2 52819 56901
0 26622 5 1 1 26621
0 26623 7 1 2 43119 26622
0 26624 5 2 1 26623
0 26625 7 1 2 45281 60810
0 26626 5 1 1 26625
0 26627 7 1 2 62407 26626
0 26628 7 1 2 69676 26627
0 26629 5 1 1 26628
0 26630 7 1 2 45114 26629
0 26631 5 1 1 26630
0 26632 7 1 2 26620 26631
0 26633 7 1 2 26618 26632
0 26634 5 1 1 26633
0 26635 7 1 2 47312 26634
0 26636 5 1 1 26635
0 26637 7 1 2 46726 59627
0 26638 5 1 1 26637
0 26639 7 1 2 69053 26638
0 26640 5 1 1 26639
0 26641 7 1 2 48472 26640
0 26642 5 1 1 26641
0 26643 7 1 2 51505 57330
0 26644 5 1 1 26643
0 26645 7 1 2 53447 26644
0 26646 5 1 1 26645
0 26647 7 1 2 62398 26646
0 26648 5 1 1 26647
0 26649 7 1 2 26642 26648
0 26650 5 1 1 26649
0 26651 7 1 2 47313 26650
0 26652 5 1 1 26651
0 26653 7 1 2 54699 69675
0 26654 5 1 1 26653
0 26655 7 1 2 51016 56856
0 26656 5 1 1 26655
0 26657 7 1 2 20431 26656
0 26658 5 1 1 26657
0 26659 7 1 2 43936 26658
0 26660 5 1 1 26659
0 26661 7 1 2 26654 26660
0 26662 7 1 2 26652 26661
0 26663 5 1 1 26662
0 26664 7 1 2 46288 26663
0 26665 5 1 1 26664
0 26666 7 1 2 61962 68047
0 26667 5 1 1 26666
0 26668 7 1 2 26665 26667
0 26669 7 1 2 26636 26668
0 26670 5 1 1 26669
0 26671 7 1 2 48133 26670
0 26672 5 1 1 26671
0 26673 7 1 2 54362 66756
0 26674 7 1 2 68805 26673
0 26675 5 1 1 26674
0 26676 7 1 2 26672 26675
0 26677 5 2 1 26676
0 26678 7 1 2 68827 69678
0 26679 5 1 1 26678
0 26680 7 1 2 60900 64915
0 26681 7 1 2 65856 26680
0 26682 7 2 2 59740 61270
0 26683 7 1 2 65048 69680
0 26684 7 1 2 26681 26683
0 26685 7 1 2 68787 26684
0 26686 5 1 1 26685
0 26687 7 1 2 44943 26686
0 26688 7 1 2 26679 26687
0 26689 5 1 1 26688
0 26690 7 1 2 26606 26689
0 26691 5 1 1 26690
0 26692 7 1 2 26497 26691
0 26693 5 1 1 26692
0 26694 7 1 2 65701 26693
0 26695 5 1 1 26694
0 26696 7 1 2 56767 68916
0 26697 5 1 1 26696
0 26698 7 1 2 69063 68866
0 26699 5 1 1 26698
0 26700 7 1 2 26697 26699
0 26701 5 1 1 26700
0 26702 7 1 2 48282 26701
0 26703 5 1 1 26702
0 26704 7 1 2 52122 61530
0 26705 7 1 2 56770 26704
0 26706 5 1 1 26705
0 26707 7 1 2 26703 26706
0 26708 5 1 1 26707
0 26709 7 1 2 46727 26708
0 26710 5 1 1 26709
0 26711 7 1 2 54615 68795
0 26712 5 2 1 26711
0 26713 7 1 2 53143 54975
0 26714 7 1 2 69133 26713
0 26715 5 1 1 26714
0 26716 7 1 2 69682 26715
0 26717 5 1 1 26716
0 26718 7 1 2 57484 26717
0 26719 5 1 1 26718
0 26720 7 1 2 26710 26719
0 26721 5 2 1 26720
0 26722 7 1 2 65911 68828
0 26723 7 1 2 69684 26722
0 26724 5 1 1 26723
0 26725 7 1 2 26695 26724
0 26726 5 1 1 26725
0 26727 7 1 2 47789 26726
0 26728 5 1 1 26727
0 26729 7 3 2 53602 69557
0 26730 7 1 2 62474 68946
0 26731 5 1 1 26730
0 26732 7 1 2 42852 1528
0 26733 5 1 1 26732
0 26734 7 1 2 52354 26733
0 26735 7 1 2 68546 26734
0 26736 5 1 1 26735
0 26737 7 1 2 26731 26736
0 26738 5 1 1 26737
0 26739 7 1 2 51017 26738
0 26740 5 1 1 26739
0 26741 7 1 2 68560 26740
0 26742 5 1 1 26741
0 26743 7 1 2 48134 26742
0 26744 5 1 1 26743
0 26745 7 1 2 49603 53125
0 26746 5 2 1 26745
0 26747 7 1 2 19514 69689
0 26748 5 1 1 26747
0 26749 7 1 2 42853 26748
0 26750 5 1 1 26749
0 26751 7 1 2 48283 68587
0 26752 5 1 1 26751
0 26753 7 1 2 26750 26752
0 26754 5 1 1 26753
0 26755 7 1 2 69139 26754
0 26756 5 1 1 26755
0 26757 7 1 2 68652 26756
0 26758 5 1 1 26757
0 26759 7 1 2 44246 26758
0 26760 5 1 1 26759
0 26761 7 1 2 51252 52048
0 26762 7 1 2 62399 26761
0 26763 5 1 1 26762
0 26764 7 1 2 26760 26763
0 26765 5 1 1 26764
0 26766 7 1 2 48633 26765
0 26767 5 1 1 26766
0 26768 7 1 2 52165 54017
0 26769 7 2 2 56322 26768
0 26770 5 1 1 69691
0 26771 7 1 2 44247 69692
0 26772 5 1 1 26771
0 26773 7 1 2 26767 26772
0 26774 5 1 1 26773
0 26775 7 1 2 43340 26774
0 26776 5 1 1 26775
0 26777 7 1 2 26744 26776
0 26778 5 1 1 26777
0 26779 7 1 2 69686 26778
0 26780 5 1 1 26779
0 26781 7 1 2 68653 69683
0 26782 5 1 1 26781
0 26783 7 1 2 48634 26782
0 26784 5 1 1 26783
0 26785 7 1 2 26770 26784
0 26786 5 1 1 26785
0 26787 7 1 2 49998 26786
0 26788 5 1 1 26787
0 26789 7 1 2 68552 68919
0 26790 5 1 1 26789
0 26791 7 1 2 26788 26790
0 26792 5 1 1 26791
0 26793 7 1 2 42220 66434
0 26794 7 1 2 26792 26793
0 26795 5 1 1 26794
0 26796 7 1 2 26780 26795
0 26797 5 1 1 26796
0 26798 7 1 2 65662 26797
0 26799 5 1 1 26798
0 26800 7 1 2 67161 67849
0 26801 5 1 1 26800
0 26802 7 2 2 59892 67202
0 26803 7 1 2 69637 69693
0 26804 5 1 1 26803
0 26805 7 1 2 26801 26804
0 26806 5 1 1 26805
0 26807 7 1 2 45282 26806
0 26808 5 1 1 26807
0 26809 7 1 2 69639 69694
0 26810 5 1 1 26809
0 26811 7 1 2 26808 26810
0 26812 5 1 1 26811
0 26813 7 1 2 64329 26812
0 26814 5 1 1 26813
0 26815 7 1 2 67162 69679
0 26816 5 1 1 26815
0 26817 7 1 2 49808 60917
0 26818 7 1 2 64916 26817
0 26819 7 1 2 64045 26818
0 26820 7 1 2 59420 26819
0 26821 5 1 1 26820
0 26822 7 1 2 44944 26821
0 26823 7 1 2 26816 26822
0 26824 5 1 1 26823
0 26825 7 1 2 67163 69650
0 26826 5 1 1 26825
0 26827 7 1 2 50277 57596
0 26828 7 1 2 58199 61594
0 26829 7 1 2 26827 26828
0 26830 7 1 2 58463 26829
0 26831 5 1 1 26830
0 26832 7 1 2 26826 26831
0 26833 5 1 1 26832
0 26834 7 1 2 69648 26833
0 26835 5 1 1 26834
0 26836 7 1 2 26570 26574
0 26837 5 1 1 26836
0 26838 7 1 2 43937 26837
0 26839 5 1 1 26838
0 26840 7 1 2 69652 26839
0 26841 5 1 1 26840
0 26842 7 1 2 67164 26841
0 26843 5 1 1 26842
0 26844 7 1 2 53706 69655
0 26845 5 1 1 26844
0 26846 7 3 2 55803 61271
0 26847 7 1 2 69661 69695
0 26848 5 1 1 26847
0 26849 7 1 2 26845 26848
0 26850 5 1 1 26849
0 26851 7 1 2 46728 26850
0 26852 5 1 1 26851
0 26853 7 1 2 59949 63273
0 26854 7 1 2 65126 69696
0 26855 7 1 2 26853 26854
0 26856 5 1 1 26855
0 26857 7 1 2 26852 26856
0 26858 5 1 1 26857
0 26859 7 1 2 43938 26858
0 26860 5 1 1 26859
0 26861 7 1 2 26843 26860
0 26862 5 1 1 26861
0 26863 7 1 2 42854 26862
0 26864 5 1 1 26863
0 26865 7 1 2 26835 26864
0 26866 5 1 1 26865
0 26867 7 1 2 44813 26866
0 26868 5 1 1 26867
0 26869 7 1 2 53707 69673
0 26870 5 1 1 26869
0 26871 7 1 2 48284 26870
0 26872 7 1 2 26868 26871
0 26873 5 1 1 26872
0 26874 7 1 2 26824 26873
0 26875 5 1 1 26874
0 26876 7 1 2 26814 26875
0 26877 5 1 1 26876
0 26878 7 1 2 69072 26877
0 26879 5 1 1 26878
0 26880 7 1 2 48019 69057
0 26881 7 1 2 69685 26880
0 26882 5 1 1 26881
0 26883 7 1 2 26879 26882
0 26884 5 1 1 26883
0 26885 7 1 2 47790 26884
0 26886 5 1 1 26885
0 26887 7 1 2 26799 26886
0 26888 5 1 1 26887
0 26889 7 1 2 66270 26888
0 26890 5 1 1 26889
0 26891 7 2 2 49999 66002
0 26892 7 1 2 53144 69698
0 26893 5 1 1 26892
0 26894 7 2 2 50861 66084
0 26895 7 1 2 47314 69700
0 26896 5 1 1 26895
0 26897 7 1 2 26893 26896
0 26898 5 1 1 26897
0 26899 7 1 2 48635 26898
0 26900 5 1 1 26899
0 26901 7 1 2 49400 65912
0 26902 5 1 1 26901
0 26903 7 1 2 26900 26902
0 26904 5 1 1 26903
0 26905 7 1 2 58823 26904
0 26906 5 1 1 26905
0 26907 7 5 2 42332 55442
0 26908 5 1 1 69702
0 26909 7 1 2 68553 69703
0 26910 5 1 1 26909
0 26911 7 1 2 52485 58503
0 26912 5 1 1 26911
0 26913 7 1 2 68556 26912
0 26914 5 1 1 26913
0 26915 7 1 2 65913 26914
0 26916 5 1 1 26915
0 26917 7 1 2 26910 26916
0 26918 7 1 2 26906 26917
0 26919 5 1 1 26918
0 26920 7 1 2 46289 26919
0 26921 5 1 1 26920
0 26922 7 1 2 65914 68558
0 26923 5 1 1 26922
0 26924 7 1 2 52494 1373
0 26925 5 2 1 26924
0 26926 7 1 2 51018 53947
0 26927 7 1 2 66116 26926
0 26928 7 1 2 69707 26927
0 26929 5 1 1 26928
0 26930 7 1 2 26923 26929
0 26931 7 1 2 26921 26930
0 26932 5 1 1 26931
0 26933 7 1 2 48135 26932
0 26934 5 1 1 26933
0 26935 7 1 2 125 52241
0 26936 5 1 1 26935
0 26937 7 1 2 49820 26936
0 26938 5 1 1 26937
0 26939 7 1 2 49451 57400
0 26940 5 1 1 26939
0 26941 7 1 2 26186 26940
0 26942 5 1 1 26941
0 26943 7 1 2 43120 26942
0 26944 5 1 1 26943
0 26945 7 1 2 26938 26944
0 26946 5 1 1 26945
0 26947 7 1 2 66003 26946
0 26948 5 1 1 26947
0 26949 7 2 2 42333 64838
0 26950 5 2 1 69709
0 26951 7 1 2 66088 69711
0 26952 5 1 1 26951
0 26953 7 1 2 44083 56627
0 26954 7 1 2 26952 26953
0 26955 5 1 1 26954
0 26956 7 1 2 26948 26955
0 26957 5 1 1 26956
0 26958 7 1 2 42855 26957
0 26959 5 1 1 26958
0 26960 7 1 2 55221 63081
0 26961 7 1 2 68590 26960
0 26962 5 1 1 26961
0 26963 7 1 2 26959 26962
0 26964 5 1 1 26963
0 26965 7 1 2 44814 50000
0 26966 7 1 2 26964 26965
0 26967 5 1 1 26966
0 26968 7 1 2 26934 26967
0 26969 5 1 1 26968
0 26970 7 1 2 62514 69627
0 26971 7 1 2 26969 26970
0 26972 5 1 1 26971
0 26973 7 2 2 45283 53708
0 26974 7 2 2 60643 66483
0 26975 7 2 2 44681 51253
0 26976 7 1 2 69715 69717
0 26977 7 1 2 69713 26976
0 26978 5 1 1 26977
0 26979 7 2 2 61001 63495
0 26980 7 1 2 53603 68168
0 26981 7 1 2 68358 26980
0 26982 7 1 2 69719 26981
0 26983 5 1 1 26982
0 26984 7 1 2 26978 26983
0 26985 5 1 1 26984
0 26986 7 1 2 66271 26985
0 26987 5 1 1 26986
0 26988 7 4 2 47791 48136
0 26989 7 1 2 44682 51376
0 26990 7 2 2 69721 26989
0 26991 7 1 2 64573 69725
0 26992 5 1 1 26991
0 26993 7 1 2 55499 59175
0 26994 7 2 2 61172 64619
0 26995 7 1 2 61258 69727
0 26996 7 1 2 26993 26995
0 26997 5 1 1 26996
0 26998 7 1 2 26992 26997
0 26999 5 2 1 26998
0 27000 7 1 2 45605 69729
0 27001 5 1 1 27000
0 27002 7 1 2 56876 63408
0 27003 7 1 2 69726 27002
0 27004 5 1 1 27003
0 27005 7 1 2 27001 27004
0 27006 5 1 1 27005
0 27007 7 1 2 68817 27006
0 27008 5 1 1 27007
0 27009 7 1 2 42047 69730
0 27010 5 1 1 27009
0 27011 7 1 2 54481 57917
0 27012 7 1 2 64620 27011
0 27013 7 2 2 47675 49880
0 27014 7 1 2 51347 52166
0 27015 7 1 2 69731 27014
0 27016 7 1 2 27012 27015
0 27017 5 1 1 27016
0 27018 7 1 2 27010 27017
0 27019 5 1 1 27018
0 27020 7 1 2 66158 67420
0 27021 7 1 2 27019 27020
0 27022 5 1 1 27021
0 27023 7 1 2 27008 27022
0 27024 7 1 2 26987 27023
0 27025 5 1 1 27024
0 27026 7 1 2 68585 27025
0 27027 5 1 1 27026
0 27028 7 1 2 42590 27027
0 27029 7 1 2 26972 27028
0 27030 7 1 2 26890 27029
0 27031 7 1 2 26728 27030
0 27032 5 1 1 27031
0 27033 7 1 2 63389 65370
0 27034 5 1 1 27033
0 27035 7 1 2 49701 65353
0 27036 7 1 2 69159 27035
0 27037 5 1 1 27036
0 27038 7 1 2 27034 27037
0 27039 5 1 1 27038
0 27040 7 2 2 48020 27039
0 27041 7 1 2 64969 69733
0 27042 5 1 1 27041
0 27043 7 2 2 57137 65367
0 27044 7 2 2 46290 59965
0 27045 7 1 2 63800 69737
0 27046 7 1 2 69735 27045
0 27047 5 1 1 27046
0 27048 7 1 2 27042 27047
0 27049 5 1 1 27048
0 27050 7 1 2 47572 27049
0 27051 5 1 1 27050
0 27052 7 1 2 52188 53001
0 27053 5 1 1 27052
0 27054 7 1 2 49347 64862
0 27055 5 1 1 27054
0 27056 7 1 2 27053 27055
0 27057 5 1 1 27056
0 27058 7 1 2 48473 27057
0 27059 5 1 1 27058
0 27060 7 1 2 57744 27059
0 27061 5 1 1 27060
0 27062 7 2 2 60408 27061
0 27063 7 1 2 63831 64752
0 27064 7 1 2 69739 27063
0 27065 5 1 1 27064
0 27066 7 1 2 27051 27065
0 27067 5 1 1 27066
0 27068 7 1 2 42048 27067
0 27069 5 1 1 27068
0 27070 7 1 2 53381 1261
0 27071 5 1 1 27070
0 27072 7 1 2 69217 27071
0 27073 5 1 1 27072
0 27074 7 1 2 64164 69218
0 27075 5 1 1 27074
0 27076 7 3 2 47573 48021
0 27077 7 2 2 45850 69741
0 27078 5 1 1 69744
0 27079 7 1 2 65789 27078
0 27080 5 1 1 27079
0 27081 7 1 2 1207 65702
0 27082 5 1 1 27081
0 27083 7 1 2 45284 27082
0 27084 5 1 1 27083
0 27085 7 1 2 54677 27084
0 27086 7 1 2 27080 27085
0 27087 5 1 1 27086
0 27088 7 1 2 27075 27087
0 27089 5 1 1 27088
0 27090 7 1 2 43121 27089
0 27091 5 1 1 27090
0 27092 7 1 2 27073 27091
0 27093 5 1 1 27092
0 27094 7 1 2 42856 27093
0 27095 5 1 1 27094
0 27096 7 1 2 46523 62416
0 27097 5 1 1 27096
0 27098 7 1 2 53126 65703
0 27099 7 1 2 69393 27098
0 27100 7 1 2 27097 27099
0 27101 5 1 1 27100
0 27102 7 1 2 27095 27101
0 27103 5 1 1 27102
0 27104 7 1 2 48137 27103
0 27105 5 1 1 27104
0 27106 7 2 2 47315 64115
0 27107 7 1 2 62347 65073
0 27108 7 1 2 69746 27107
0 27109 5 1 1 27108
0 27110 7 1 2 27105 27109
0 27111 5 1 1 27110
0 27112 7 1 2 54482 64753
0 27113 7 1 2 27111 27112
0 27114 5 1 1 27113
0 27115 7 1 2 27069 27114
0 27116 5 1 1 27115
0 27117 7 1 2 45471 27116
0 27118 5 1 1 27117
0 27119 7 3 2 47316 49860
0 27120 5 2 1 69748
0 27121 7 1 2 45115 57254
0 27122 5 1 1 27121
0 27123 7 1 2 69751 27122
0 27124 5 2 1 27123
0 27125 7 1 2 54018 69753
0 27126 5 1 1 27125
0 27127 7 1 2 64851 68452
0 27128 5 1 1 27127
0 27129 7 1 2 27126 27128
0 27130 5 1 1 27129
0 27131 7 1 2 43341 27130
0 27132 5 1 1 27131
0 27133 7 1 2 53478 54700
0 27134 7 1 2 49530 27133
0 27135 5 1 1 27134
0 27136 7 1 2 27132 27135
0 27137 5 1 1 27136
0 27138 7 3 2 60409 27137
0 27139 7 1 2 67263 69755
0 27140 5 1 1 27139
0 27141 7 1 2 27118 27140
0 27142 5 1 1 27141
0 27143 7 1 2 44945 27142
0 27144 5 1 1 27143
0 27145 7 1 2 46524 49498
0 27146 5 2 1 27145
0 27147 7 1 2 46291 68608
0 27148 5 1 1 27147
0 27149 7 1 2 69758 27148
0 27150 5 1 1 27149
0 27151 7 1 2 44248 27150
0 27152 5 1 1 27151
0 27153 7 1 2 57378 64855
0 27154 5 1 1 27153
0 27155 7 1 2 27152 27154
0 27156 5 1 1 27155
0 27157 7 1 2 44084 27156
0 27158 5 1 1 27157
0 27159 7 1 2 57328 63624
0 27160 5 1 1 27159
0 27161 7 1 2 55382 27160
0 27162 5 1 1 27161
0 27163 7 1 2 27158 27162
0 27164 5 1 1 27163
0 27165 7 3 2 68257 27164
0 27166 7 1 2 67264 69760
0 27167 5 1 1 27166
0 27168 7 1 2 27144 27167
0 27169 5 1 1 27168
0 27170 7 1 2 67020 27169
0 27171 5 1 1 27170
0 27172 7 1 2 45851 69761
0 27173 5 1 1 27172
0 27174 7 1 2 45852 69756
0 27175 5 1 1 27174
0 27176 7 3 2 45853 63454
0 27177 5 1 1 69763
0 27178 7 1 2 65790 27177
0 27179 5 3 1 27178
0 27180 7 1 2 47574 44815
0 27181 7 1 2 45116 27180
0 27182 7 1 2 62096 27181
0 27183 7 1 2 69766 27182
0 27184 5 1 1 27183
0 27185 7 2 2 46729 69740
0 27186 7 1 2 45854 69769
0 27187 5 1 1 27186
0 27188 7 1 2 27184 27187
0 27189 5 1 1 27188
0 27190 7 1 2 45472 27189
0 27191 5 1 1 27190
0 27192 7 1 2 27175 27191
0 27193 5 1 1 27192
0 27194 7 1 2 44946 27193
0 27195 5 1 1 27194
0 27196 7 1 2 27173 27195
0 27197 5 1 1 27196
0 27198 7 1 2 53709 27197
0 27199 5 1 1 27198
0 27200 7 1 2 56022 58902
0 27201 7 1 2 53547 27200
0 27202 7 5 2 48022 52642
0 27203 7 1 2 63285 69771
0 27204 7 1 2 27201 27203
0 27205 7 1 2 56285 27204
0 27206 5 1 1 27205
0 27207 7 1 2 27199 27206
0 27208 5 1 1 27207
0 27209 7 1 2 66272 27208
0 27210 5 1 1 27209
0 27211 7 1 2 61205 69734
0 27212 5 1 1 27211
0 27213 7 1 2 60967 64304
0 27214 7 1 2 69736 27213
0 27215 5 1 1 27214
0 27216 7 1 2 27212 27215
0 27217 5 1 1 27216
0 27218 7 1 2 47575 27217
0 27219 5 1 1 27218
0 27220 7 1 2 63995 69770
0 27221 5 1 1 27220
0 27222 7 1 2 27219 27221
0 27223 5 1 1 27222
0 27224 7 1 2 45473 27223
0 27225 5 1 1 27224
0 27226 7 1 2 63996 69757
0 27227 5 1 1 27226
0 27228 7 1 2 27225 27227
0 27229 5 1 1 27228
0 27230 7 1 2 44947 27229
0 27231 5 1 1 27230
0 27232 7 1 2 63997 69762
0 27233 5 1 1 27232
0 27234 7 1 2 27231 27233
0 27235 5 1 1 27234
0 27236 7 1 2 69336 27235
0 27237 5 1 1 27236
0 27238 7 1 2 66766 19655
0 27239 5 1 1 27238
0 27240 7 1 2 54248 27239
0 27241 5 2 1 27240
0 27242 7 1 2 60245 68643
0 27243 7 1 2 65116 27242
0 27244 5 1 1 27243
0 27245 7 1 2 69776 27244
0 27246 5 1 1 27245
0 27247 7 1 2 52302 27246
0 27248 5 1 1 27247
0 27249 7 1 2 46292 67221
0 27250 7 1 2 50340 27249
0 27251 5 1 1 27250
0 27252 7 1 2 27248 27251
0 27253 5 2 1 27252
0 27254 7 3 2 53604 67699
0 27255 5 1 1 69780
0 27256 7 2 2 62675 68781
0 27257 5 1 1 69783
0 27258 7 1 2 27255 27257
0 27259 5 4 1 27258
0 27260 7 1 2 54790 69785
0 27261 5 1 1 27260
0 27262 7 1 2 63230 69055
0 27263 5 1 1 27262
0 27264 7 1 2 27261 27263
0 27265 5 1 1 27264
0 27266 7 1 2 48636 69210
0 27267 7 1 2 27265 27266
0 27268 7 1 2 69778 27267
0 27269 5 1 1 27268
0 27270 7 1 2 27237 27269
0 27271 7 1 2 27210 27270
0 27272 7 1 2 27171 27271
0 27273 5 1 1 27272
0 27274 7 1 2 47792 27273
0 27275 5 1 1 27274
0 27276 7 2 2 44469 52875
0 27277 7 1 2 55439 57492
0 27278 7 2 2 61283 27277
0 27279 7 1 2 69789 69791
0 27280 5 1 1 27279
0 27281 7 1 2 42857 57164
0 27282 5 1 1 27281
0 27283 7 1 2 58791 60714
0 27284 5 1 1 27283
0 27285 7 1 2 27282 27284
0 27286 5 2 1 27285
0 27287 7 1 2 52595 69793
0 27288 7 1 2 56174 27287
0 27289 5 1 1 27288
0 27290 7 1 2 27280 27289
0 27291 5 1 1 27290
0 27292 7 1 2 66322 27291
0 27293 5 1 1 27292
0 27294 7 2 2 56713 68528
0 27295 7 1 2 69790 69795
0 27296 5 1 1 27295
0 27297 7 1 2 45117 56938
0 27298 7 1 2 54791 27297
0 27299 7 1 2 69794 27298
0 27300 5 1 1 27299
0 27301 7 1 2 27296 27300
0 27302 5 1 1 27301
0 27303 7 1 2 66383 68408
0 27304 7 1 2 27302 27303
0 27305 5 1 1 27304
0 27306 7 1 2 27293 27305
0 27307 5 1 1 27306
0 27308 7 1 2 67684 27307
0 27309 5 1 1 27308
0 27310 7 1 2 52215 53532
0 27311 5 1 1 27310
0 27312 7 2 2 51389 27311
0 27313 7 2 2 53170 69797
0 27314 7 1 2 65857 69799
0 27315 5 1 1 27314
0 27316 7 1 2 66423 67880
0 27317 7 1 2 56082 27316
0 27318 7 1 2 56714 27317
0 27319 5 1 1 27318
0 27320 7 1 2 27315 27319
0 27321 5 1 1 27320
0 27322 7 1 2 45855 27321
0 27323 5 1 1 27322
0 27324 7 2 2 57981 69587
0 27325 7 1 2 49918 65865
0 27326 7 1 2 69801 27325
0 27327 5 1 1 27326
0 27328 7 1 2 27323 27327
0 27329 5 1 1 27328
0 27330 7 1 2 43553 27329
0 27331 5 1 1 27330
0 27332 7 2 2 43646 69798
0 27333 7 1 2 68942 69305
0 27334 7 1 2 69803 27333
0 27335 5 1 1 27334
0 27336 7 1 2 27331 27335
0 27337 5 1 1 27336
0 27338 7 1 2 42221 27337
0 27339 5 1 1 27338
0 27340 7 1 2 68052 67916
0 27341 7 1 2 69804 27340
0 27342 5 1 1 27341
0 27343 7 1 2 27339 27342
0 27344 5 1 1 27343
0 27345 7 1 2 67554 27344
0 27346 5 1 1 27345
0 27347 7 1 2 52963 63735
0 27348 7 1 2 67743 27347
0 27349 5 1 1 27348
0 27350 7 1 2 49477 54682
0 27351 5 2 1 27350
0 27352 7 1 2 51707 69687
0 27353 7 1 2 69805 27352
0 27354 5 1 1 27353
0 27355 7 1 2 27349 27354
0 27356 5 1 1 27355
0 27357 7 1 2 66273 27356
0 27358 5 1 1 27357
0 27359 7 1 2 69701 69806
0 27360 5 1 1 27359
0 27361 7 1 2 42334 58310
0 27362 7 1 2 69009 27361
0 27363 5 1 1 27362
0 27364 7 1 2 27360 27363
0 27365 5 1 1 27364
0 27366 7 1 2 68818 27365
0 27367 5 1 1 27366
0 27368 7 1 2 27358 27367
0 27369 5 1 1 27368
0 27370 7 1 2 56597 27369
0 27371 5 1 1 27370
0 27372 7 1 2 69211 69800
0 27373 5 1 1 27372
0 27374 7 1 2 66079 69203
0 27375 7 1 2 69802 27374
0 27376 5 1 1 27375
0 27377 7 1 2 27373 27376
0 27378 5 1 1 27377
0 27379 7 1 2 69786 27378
0 27380 5 1 1 27379
0 27381 7 1 2 47317 56083
0 27382 7 1 2 68254 27381
0 27383 7 1 2 62337 69257
0 27384 7 1 2 27382 27383
0 27385 5 1 1 27384
0 27386 7 1 2 27380 27385
0 27387 7 1 2 27371 27386
0 27388 7 1 2 27346 27387
0 27389 5 1 1 27388
0 27390 7 1 2 44470 27389
0 27391 5 1 1 27390
0 27392 7 1 2 48474 65204
0 27393 5 1 1 27392
0 27394 7 1 2 1053 27393
0 27395 5 1 1 27394
0 27396 7 2 2 44683 27395
0 27397 7 1 2 66274 69807
0 27398 5 1 1 27397
0 27399 7 1 2 46993 52643
0 27400 7 1 2 54647 65858
0 27401 7 1 2 27399 27400
0 27402 7 1 2 57165 27401
0 27403 5 1 1 27402
0 27404 7 1 2 27398 27403
0 27405 5 1 1 27404
0 27406 7 1 2 43122 27405
0 27407 5 1 1 27406
0 27408 7 1 2 58470 58486
0 27409 5 1 1 27408
0 27410 7 2 2 65079 27409
0 27411 7 1 2 66275 69809
0 27412 5 1 1 27411
0 27413 7 1 2 27407 27412
0 27414 5 1 1 27413
0 27415 7 1 2 42858 27414
0 27416 5 1 1 27415
0 27417 7 1 2 61691 64928
0 27418 5 2 1 27417
0 27419 7 2 2 65085 69811
0 27420 7 1 2 66276 69813
0 27421 5 1 1 27420
0 27422 7 1 2 27416 27421
0 27423 5 1 1 27422
0 27424 7 1 2 45856 27423
0 27425 5 1 1 27424
0 27426 7 1 2 52066 69812
0 27427 5 1 1 27426
0 27428 7 1 2 51982 60750
0 27429 5 1 1 27428
0 27430 7 1 2 27427 27429
0 27431 5 1 1 27430
0 27432 7 1 2 48475 27431
0 27433 5 1 1 27432
0 27434 7 1 2 57745 27433
0 27435 5 1 1 27434
0 27436 7 1 2 47031 63231
0 27437 7 3 2 66318 27436
0 27438 7 1 2 27435 69815
0 27439 5 1 1 27438
0 27440 7 1 2 27425 27439
0 27441 5 1 1 27440
0 27442 7 1 2 53311 69722
0 27443 7 1 2 27441 27442
0 27444 5 1 1 27443
0 27445 7 1 2 48908 27444
0 27446 7 1 2 27391 27445
0 27447 5 1 1 27446
0 27448 7 1 2 42222 69519
0 27449 5 1 1 27448
0 27450 7 1 2 66194 68144
0 27451 5 1 1 27450
0 27452 7 1 2 27449 27451
0 27453 5 3 1 27452
0 27454 7 1 2 69814 69818
0 27455 5 1 1 27454
0 27456 7 1 2 69810 69819
0 27457 5 1 1 27456
0 27458 7 1 2 69808 69820
0 27459 5 1 1 27458
0 27460 7 1 2 53605 68163
0 27461 5 2 1 27460
0 27462 7 1 2 68255 69037
0 27463 5 1 1 27462
0 27464 7 1 2 69821 27463
0 27465 5 2 1 27464
0 27466 7 1 2 49227 63455
0 27467 7 1 2 54678 27466
0 27468 7 1 2 69823 27467
0 27469 5 1 1 27468
0 27470 7 1 2 27459 27469
0 27471 5 1 1 27470
0 27472 7 1 2 43123 27471
0 27473 5 1 1 27472
0 27474 7 1 2 27457 27473
0 27475 5 1 1 27474
0 27476 7 1 2 42859 27475
0 27477 5 1 1 27476
0 27478 7 1 2 27455 27477
0 27479 5 1 1 27478
0 27480 7 1 2 69723 27479
0 27481 5 1 1 27480
0 27482 7 1 2 48918 27481
0 27483 5 1 1 27482
0 27484 7 1 2 44948 58207
0 27485 7 1 2 27483 27484
0 27486 7 1 2 27447 27485
0 27487 5 1 1 27486
0 27488 7 1 2 27309 27487
0 27489 5 1 1 27488
0 27490 7 1 2 45285 27489
0 27491 5 1 1 27490
0 27492 7 1 2 42335 69309
0 27493 5 1 1 27492
0 27494 7 1 2 25027 27493
0 27495 5 2 1 27494
0 27496 7 1 2 42223 69825
0 27497 5 1 1 27496
0 27498 7 1 2 68094 67917
0 27499 5 1 1 27498
0 27500 7 1 2 27497 27499
0 27501 5 5 1 27500
0 27502 7 1 2 54792 69827
0 27503 5 1 1 27502
0 27504 7 2 2 47032 53651
0 27505 7 1 2 64687 66159
0 27506 7 1 2 69832 27505
0 27507 5 1 1 27506
0 27508 7 1 2 27503 27507
0 27509 5 1 1 27508
0 27510 7 1 2 47793 69779
0 27511 7 1 2 27509 27510
0 27512 5 1 1 27511
0 27513 7 1 2 48138 68634
0 27514 5 1 1 27513
0 27515 7 1 2 69777 27514
0 27516 5 1 1 27515
0 27517 7 1 2 42049 58928
0 27518 7 1 2 69828 27517
0 27519 7 1 2 27516 27518
0 27520 5 1 1 27519
0 27521 7 1 2 27512 27520
0 27522 5 1 1 27521
0 27523 7 1 2 48637 27522
0 27524 5 1 1 27523
0 27525 7 2 2 46730 69353
0 27526 5 1 1 69834
0 27527 7 2 2 50380 69212
0 27528 7 1 2 51834 56239
0 27529 7 1 2 56256 27528
0 27530 7 1 2 69836 27529
0 27531 7 1 2 69835 27530
0 27532 5 1 1 27531
0 27533 7 1 2 27524 27532
0 27534 5 1 1 27533
0 27535 7 1 2 67555 27534
0 27536 5 1 1 27535
0 27537 7 2 2 52876 62470
0 27538 7 1 2 64655 69838
0 27539 5 1 1 27538
0 27540 7 1 2 56645 67537
0 27541 7 1 2 68846 27540
0 27542 5 1 1 27541
0 27543 7 1 2 27539 27542
0 27544 5 1 1 27543
0 27545 7 1 2 51019 27544
0 27546 5 1 1 27545
0 27547 7 1 2 43939 52209
0 27548 5 1 1 27547
0 27549 7 3 2 44249 62129
0 27550 7 1 2 67885 69840
0 27551 7 1 2 27548 27550
0 27552 5 1 1 27551
0 27553 7 1 2 54701 62838
0 27554 7 1 2 64384 27553
0 27555 5 1 1 27554
0 27556 7 1 2 27552 27555
0 27557 5 1 1 27556
0 27558 7 1 2 45474 27557
0 27559 5 1 1 27558
0 27560 7 1 2 27546 27559
0 27561 5 1 1 27560
0 27562 7 1 2 46293 27561
0 27563 5 1 1 27562
0 27564 7 2 2 58348 62130
0 27565 7 1 2 53145 53365
0 27566 7 1 2 64322 27565
0 27567 7 1 2 69843 27566
0 27568 5 1 1 27567
0 27569 7 1 2 27563 27568
0 27570 5 1 1 27569
0 27571 7 1 2 48285 27570
0 27572 5 1 1 27571
0 27573 7 1 2 51708 56315
0 27574 5 1 1 27573
0 27575 7 1 2 54184 59630
0 27576 5 1 1 27575
0 27577 7 1 2 27574 27576
0 27578 5 1 1 27577
0 27579 7 1 2 43124 27578
0 27580 5 1 1 27579
0 27581 7 1 2 64423 68967
0 27582 5 1 1 27581
0 27583 7 1 2 27580 27582
0 27584 5 1 1 27583
0 27585 7 1 2 68228 27584
0 27586 5 1 1 27585
0 27587 7 1 2 27572 27586
0 27588 5 1 1 27587
0 27589 7 1 2 69829 27588
0 27590 5 1 1 27589
0 27591 7 2 2 50001 69784
0 27592 5 1 1 69845
0 27593 7 1 2 51768 69781
0 27594 5 1 1 27593
0 27595 7 1 2 27592 27594
0 27596 5 1 1 27595
0 27597 7 1 2 65025 27596
0 27598 5 1 1 27597
0 27599 7 1 2 62676 64754
0 27600 7 1 2 69839 27599
0 27601 5 1 1 27600
0 27602 7 1 2 27598 27601
0 27603 5 1 1 27602
0 27604 7 1 2 51020 27603
0 27605 5 1 1 27604
0 27606 7 2 2 47576 55433
0 27607 7 1 2 62669 69847
0 27608 5 1 1 27607
0 27609 7 1 2 43342 62677
0 27610 7 1 2 69841 27609
0 27611 5 1 1 27610
0 27612 7 1 2 27608 27611
0 27613 5 1 1 27612
0 27614 7 1 2 42224 27613
0 27615 5 1 1 27614
0 27616 7 1 2 63983 69848
0 27617 5 1 1 27616
0 27618 7 1 2 27615 27617
0 27619 5 1 1 27618
0 27620 7 1 2 49299 27619
0 27621 5 1 1 27620
0 27622 7 2 2 61858 62678
0 27623 7 1 2 53146 69842
0 27624 7 1 2 69849 27623
0 27625 5 1 1 27624
0 27626 7 1 2 27621 27625
0 27627 5 1 1 27626
0 27628 7 1 2 45475 27627
0 27629 5 1 1 27628
0 27630 7 1 2 27605 27629
0 27631 5 1 1 27630
0 27632 7 1 2 46294 27631
0 27633 5 1 1 27632
0 27634 7 1 2 64911 65026
0 27635 7 1 2 69846 27634
0 27636 5 1 1 27635
0 27637 7 1 2 48286 27636
0 27638 7 1 2 27633 27637
0 27639 5 1 1 27638
0 27640 7 1 2 52262 68969
0 27641 5 1 1 27640
0 27642 7 1 2 69782 27641
0 27643 5 1 1 27642
0 27644 7 1 2 62131 65120
0 27645 7 1 2 69850 27644
0 27646 5 1 1 27645
0 27647 7 1 2 27643 27646
0 27648 5 1 1 27647
0 27649 7 1 2 50954 27648
0 27650 5 1 1 27649
0 27651 7 3 2 52644 53606
0 27652 7 4 2 48023 49348
0 27653 7 1 2 57089 63384
0 27654 7 1 2 69854 27653
0 27655 7 1 2 69851 27654
0 27656 5 1 1 27655
0 27657 7 1 2 27650 27656
0 27658 5 1 1 27657
0 27659 7 1 2 42860 27658
0 27660 5 1 1 27659
0 27661 7 2 2 48638 55434
0 27662 7 1 2 43602 55234
0 27663 7 1 2 50890 27662
0 27664 7 1 2 69858 27663
0 27665 7 1 2 58829 27664
0 27666 5 1 1 27665
0 27667 7 1 2 44949 27666
0 27668 7 1 2 27660 27667
0 27669 5 1 1 27668
0 27670 7 1 2 69213 27669
0 27671 7 1 2 27639 27670
0 27672 5 1 1 27671
0 27673 7 1 2 27590 27672
0 27674 5 1 1 27673
0 27675 7 1 2 48139 27674
0 27676 5 1 1 27675
0 27677 7 1 2 52167 54357
0 27678 7 1 2 69787 27677
0 27679 7 1 2 69223 27678
0 27680 5 1 1 27679
0 27681 7 1 2 69264 69410
0 27682 5 1 1 27681
0 27683 7 1 2 51889 65885
0 27684 5 1 1 27683
0 27685 7 1 2 27682 27684
0 27686 5 1 1 27685
0 27687 7 1 2 42225 27686
0 27688 5 1 1 27687
0 27689 7 1 2 58889 69527
0 27690 5 1 1 27689
0 27691 7 1 2 27688 27690
0 27692 5 3 1 27691
0 27693 7 1 2 58320 60112
0 27694 7 1 2 69354 27693
0 27695 7 1 2 69860 27694
0 27696 5 1 1 27695
0 27697 7 1 2 27680 27696
0 27698 7 1 2 27676 27697
0 27699 5 1 1 27698
0 27700 7 1 2 48923 27699
0 27701 5 1 1 27700
0 27702 7 1 2 27536 27701
0 27703 7 1 2 27491 27702
0 27704 7 1 2 27275 27703
0 27705 5 1 1 27704
0 27706 7 1 2 44345 27705
0 27707 5 1 1 27706
0 27708 7 3 2 59724 64069
0 27709 7 1 2 55276 69863
0 27710 5 1 1 27709
0 27711 7 1 2 20838 27710
0 27712 5 1 1 27711
0 27713 7 1 2 46731 27712
0 27714 5 1 1 27713
0 27715 7 2 2 47577 60233
0 27716 7 1 2 59759 69866
0 27717 5 1 1 27716
0 27718 7 1 2 59550 27717
0 27719 5 1 1 27718
0 27720 7 1 2 42050 27719
0 27721 5 1 1 27720
0 27722 7 1 2 58106 69867
0 27723 5 1 1 27722
0 27724 7 1 2 27721 27723
0 27725 5 1 1 27724
0 27726 7 1 2 58873 27725
0 27727 5 1 1 27726
0 27728 7 1 2 27714 27727
0 27729 5 1 1 27728
0 27730 7 1 2 46525 27729
0 27731 5 1 1 27730
0 27732 7 4 2 61767 63195
0 27733 7 2 2 46732 69868
0 27734 7 1 2 62292 69872
0 27735 5 1 1 27734
0 27736 7 1 2 27731 27735
0 27737 5 1 1 27736
0 27738 7 1 2 45118 27737
0 27739 5 1 1 27738
0 27740 7 1 2 44346 61305
0 27741 7 1 2 69792 27740
0 27742 5 1 1 27741
0 27743 7 1 2 27739 27742
0 27744 5 1 1 27743
0 27745 7 1 2 47318 27744
0 27746 5 1 1 27745
0 27747 7 1 2 57459 59694
0 27748 7 2 2 62660 63397
0 27749 7 1 2 68048 69874
0 27750 7 1 2 27747 27749
0 27751 5 1 1 27750
0 27752 7 1 2 27746 27751
0 27753 5 1 1 27752
0 27754 7 1 2 69837 27753
0 27755 5 1 1 27754
0 27756 7 1 2 55914 61607
0 27757 5 1 1 27756
0 27758 7 1 2 47794 69130
0 27759 7 1 2 65143 27758
0 27760 5 1 1 27759
0 27761 7 1 2 27757 27760
0 27762 5 1 1 27761
0 27763 7 1 2 44347 27762
0 27764 5 1 1 27763
0 27765 7 1 2 56706 63925
0 27766 7 1 2 64633 27765
0 27767 5 1 1 27766
0 27768 7 1 2 27764 27767
0 27769 5 2 1 27768
0 27770 7 1 2 69830 69876
0 27771 5 1 1 27770
0 27772 7 1 2 57166 60933
0 27773 5 1 1 27772
0 27774 7 1 2 45606 58055
0 27775 5 1 1 27774
0 27776 7 1 2 60506 27775
0 27777 5 1 1 27776
0 27778 7 1 2 57056 63895
0 27779 7 1 2 27777 27778
0 27780 5 1 1 27779
0 27781 7 1 2 27773 27780
0 27782 5 1 1 27781
0 27783 7 1 2 49300 27782
0 27784 5 1 1 27783
0 27785 7 1 2 56789 60934
0 27786 5 1 1 27785
0 27787 7 1 2 27784 27786
0 27788 5 1 1 27787
0 27789 7 2 2 51021 27788
0 27790 7 1 2 46939 68085
0 27791 7 1 2 69878 27790
0 27792 5 1 1 27791
0 27793 7 1 2 27771 27792
0 27794 5 1 1 27793
0 27795 7 1 2 67222 27794
0 27796 5 1 1 27795
0 27797 7 1 2 27755 27796
0 27798 5 1 1 27797
0 27799 7 1 2 67556 27798
0 27800 5 1 1 27799
0 27801 7 1 2 58056 68086
0 27802 5 1 1 27801
0 27803 7 1 2 44471 69269
0 27804 5 1 1 27803
0 27805 7 1 2 27802 27804
0 27806 5 1 1 27805
0 27807 7 1 2 45607 27806
0 27808 5 1 1 27807
0 27809 7 1 2 67771 68381
0 27810 7 1 2 68523 27809
0 27811 5 1 1 27810
0 27812 7 1 2 27808 27811
0 27813 5 1 1 27812
0 27814 7 1 2 69411 27813
0 27815 5 1 1 27814
0 27816 7 1 2 67913 68495
0 27817 5 1 1 27816
0 27818 7 1 2 48024 64578
0 27819 5 1 1 27818
0 27820 7 1 2 27817 27819
0 27821 5 1 1 27820
0 27822 7 1 2 46852 27821
0 27823 5 1 1 27822
0 27824 7 1 2 44472 69364
0 27825 5 1 1 27824
0 27826 7 1 2 27823 27825
0 27827 5 1 1 27826
0 27828 7 1 2 45608 27827
0 27829 5 1 1 27828
0 27830 7 1 2 57502 58909
0 27831 7 1 2 63810 27830
0 27832 5 1 1 27831
0 27833 7 1 2 27829 27832
0 27834 5 1 1 27833
0 27835 7 1 2 69401 27834
0 27836 5 1 1 27835
0 27837 7 1 2 27815 27836
0 27838 5 1 1 27837
0 27839 7 1 2 47676 57982
0 27840 7 1 2 52286 27839
0 27841 7 1 2 62348 27840
0 27842 7 1 2 27838 27841
0 27843 5 1 1 27842
0 27844 7 1 2 27800 27843
0 27845 7 2 2 68529 69861
0 27846 7 1 2 57460 69880
0 27847 5 1 1 27846
0 27848 7 1 2 43476 68087
0 27849 5 1 1 27848
0 27850 7 1 2 24887 27849
0 27851 5 1 1 27850
0 27852 7 1 2 42051 27851
0 27853 5 1 1 27852
0 27854 7 1 2 69204 69451
0 27855 5 1 1 27854
0 27856 7 1 2 27853 27855
0 27857 5 1 1 27856
0 27858 7 1 2 27857 69413
0 27859 5 1 1 27858
0 27860 7 1 2 42052 69366
0 27861 5 1 1 27860
0 27862 7 1 2 55415 69255
0 27863 5 1 1 27862
0 27864 7 1 2 27861 27863
0 27865 5 1 1 27864
0 27866 7 1 2 27865 69402
0 27867 5 1 1 27866
0 27868 7 1 2 27859 27867
0 27869 5 1 1 27868
0 27870 7 1 2 47795 45119
0 27871 7 1 2 27869 27870
0 27872 5 1 1 27871
0 27873 7 1 2 27847 27872
0 27874 5 1 1 27873
0 27875 7 1 2 55277 27874
0 27876 5 1 1 27875
0 27877 7 1 2 68289 69881
0 27878 5 1 1 27877
0 27879 7 1 2 27876 27878
0 27880 5 1 1 27879
0 27881 7 1 2 69502 27880
0 27882 5 1 1 27881
0 27883 7 1 2 44473 52281
0 27884 7 1 2 69796 27883
0 27885 7 1 2 69862 27884
0 27886 5 1 1 27885
0 27887 7 1 2 27882 27886
0 27888 5 1 1 27887
0 27889 7 1 2 50381 27888
0 27890 5 1 1 27889
0 27891 7 1 2 58949 60960
0 27892 7 1 2 68412 27891
0 27893 5 1 1 27892
0 27894 7 1 2 55929 57448
0 27895 5 1 1 27894
0 27896 7 1 2 64755 67700
0 27897 7 1 2 27895 27896
0 27898 5 1 1 27897
0 27899 7 1 2 27893 27898
0 27900 5 1 1 27899
0 27901 7 4 2 52454 57983
0 27902 7 1 2 27900 69882
0 27903 5 1 1 27902
0 27904 7 2 2 55915 67542
0 27905 7 1 2 56158 64756
0 27906 7 1 2 69886 27905
0 27907 5 1 1 27906
0 27908 7 1 2 27903 27907
0 27909 5 1 1 27908
0 27910 7 1 2 42053 27909
0 27911 5 1 1 27910
0 27912 7 1 2 46733 63422
0 27913 7 1 2 69460 27912
0 27914 7 1 2 67253 27913
0 27915 5 1 1 27914
0 27916 7 1 2 27911 27915
0 27917 5 1 1 27916
0 27918 7 1 2 69826 27917
0 27919 5 1 1 27918
0 27920 7 3 2 52123 68274
0 27921 5 1 1 69888
0 27922 7 5 2 42054 63998
0 27923 7 1 2 69889 69891
0 27924 7 1 2 69435 27923
0 27925 5 1 1 27924
0 27926 7 1 2 66337 69833
0 27927 5 1 1 27926
0 27928 7 1 2 53631 69265
0 27929 5 1 1 27928
0 27930 7 1 2 27927 27929
0 27931 5 1 1 27930
0 27932 7 1 2 42055 27931
0 27933 5 1 1 27932
0 27934 7 1 2 54483 67188
0 27935 7 1 2 68095 27934
0 27936 5 1 1 27935
0 27937 7 1 2 27933 27936
0 27938 5 1 1 27937
0 27939 7 1 2 63958 64963
0 27940 7 1 2 27938 27939
0 27941 5 1 1 27940
0 27942 7 1 2 48909 68096
0 27943 7 1 2 67664 69104
0 27944 7 1 2 27942 27943
0 27945 5 1 1 27944
0 27946 7 1 2 27941 27945
0 27947 5 1 1 27946
0 27948 7 1 2 16613 23039
0 27949 5 1 1 27948
0 27950 7 1 2 67547 69883
0 27951 7 1 2 27949 27950
0 27952 7 1 2 27947 27951
0 27953 5 1 1 27952
0 27954 7 1 2 27925 27953
0 27955 7 1 2 27919 27954
0 27956 5 1 1 27955
0 27957 7 1 2 62293 27956
0 27958 5 1 1 27957
0 27959 7 1 2 49919 67543
0 27960 5 1 1 27959
0 27961 7 1 2 46994 69368
0 27962 5 1 1 27961
0 27963 7 1 2 27960 27962
0 27964 5 1 1 27963
0 27965 7 1 2 48924 51022
0 27966 7 1 2 56159 27965
0 27967 7 1 2 27964 27966
0 27968 7 1 2 69831 27967
0 27969 5 1 1 27968
0 27970 7 1 2 27958 27969
0 27971 7 1 2 27890 27970
0 27972 5 1 1 27971
0 27973 7 1 2 44348 27972
0 27974 5 1 1 27973
0 27975 7 1 2 53312 69879
0 27976 5 1 1 27975
0 27977 7 1 2 61940 69873
0 27978 5 1 1 27977
0 27979 7 1 2 27976 27978
0 27980 5 1 1 27979
0 27981 7 1 2 63232 27980
0 27982 5 1 1 27981
0 27983 7 1 2 69788 69877
0 27984 5 1 1 27983
0 27985 7 1 2 48910 51023
0 27986 7 1 2 61438 27985
0 27987 7 1 2 64034 27986
0 27988 7 1 2 68347 27987
0 27989 5 1 1 27988
0 27990 7 1 2 27984 27989
0 27991 7 1 2 27982 27990
0 27992 5 1 1 27991
0 27993 7 1 2 67223 27992
0 27994 5 1 1 27993
0 27995 7 3 2 47796 67165
0 27996 7 1 2 69884 69389
0 27997 7 1 2 69355 27996
0 27998 7 1 2 69896 27997
0 27999 5 1 1 27998
0 28000 7 1 2 27994 27999
0 28001 5 1 1 28000
0 28002 7 1 2 69214 28001
0 28003 5 1 1 28002
0 28004 7 1 2 27974 28003
0 28005 7 1 2 27844 28004
0 28006 5 1 1 28005
0 28007 7 1 2 64727 28006
0 28008 5 1 1 28007
0 28009 7 1 2 46070 28008
0 28010 7 1 2 27707 28009
0 28011 5 1 1 28010
0 28012 7 1 2 27032 28011
0 28013 5 1 1 28012
0 28014 7 1 2 63736 67007
0 28015 5 1 1 28014
0 28016 7 1 2 69822 28015
0 28017 5 1 1 28016
0 28018 7 1 2 42861 63714
0 28019 5 1 1 28018
0 28020 7 1 2 61783 62414
0 28021 5 1 1 28020
0 28022 7 1 2 28019 28021
0 28023 5 2 1 28022
0 28024 7 2 2 51254 52282
0 28025 7 1 2 58030 65663
0 28026 7 1 2 69901 28025
0 28027 7 1 2 69899 28026
0 28028 7 1 2 28017 28027
0 28029 5 1 1 28028
0 28030 7 1 2 47911 28029
0 28031 7 1 2 28013 28030
0 28032 5 1 1 28031
0 28033 7 1 2 47130 28032
0 28034 7 1 2 26461 28033
0 28035 5 1 1 28034
0 28036 7 1 2 45476 60811
0 28037 5 1 1 28036
0 28038 7 1 2 65470 28037
0 28039 5 1 1 28038
0 28040 7 1 2 46526 28039
0 28041 5 1 1 28040
0 28042 7 1 2 50955 57379
0 28043 5 3 1 28042
0 28044 7 1 2 28041 69903
0 28045 5 1 1 28044
0 28046 7 1 2 48639 28045
0 28047 5 1 1 28046
0 28048 7 1 2 51878 54895
0 28049 5 1 1 28048
0 28050 7 1 2 28047 28049
0 28051 5 1 1 28050
0 28052 7 1 2 66545 28051
0 28053 5 1 1 28052
0 28054 7 1 2 52929 62405
0 28055 5 1 1 28054
0 28056 7 2 2 59721 28055
0 28057 5 1 1 69906
0 28058 7 1 2 42862 69907
0 28059 5 1 1 28058
0 28060 7 1 2 46295 12479
0 28061 5 1 1 28060
0 28062 7 1 2 68360 28061
0 28063 7 1 2 28059 28062
0 28064 5 1 1 28063
0 28065 7 1 2 28053 28064
0 28066 5 1 1 28065
0 28067 7 1 2 59441 28066
0 28068 5 1 1 28067
0 28069 7 1 2 61638 67382
0 28070 5 1 1 28069
0 28071 7 1 2 64757 69099
0 28072 5 1 1 28071
0 28073 7 1 2 28070 28072
0 28074 5 1 1 28073
0 28075 7 1 2 42056 28074
0 28076 5 1 1 28075
0 28077 7 2 2 50002 61081
0 28078 7 1 2 47677 69908
0 28079 7 1 2 53675 28078
0 28080 5 1 1 28079
0 28081 7 1 2 28076 28080
0 28082 5 1 1 28081
0 28083 7 1 2 52921 28082
0 28084 5 1 1 28083
0 28085 7 2 2 50091 59916
0 28086 5 1 1 69910
0 28087 7 1 2 52789 69911
0 28088 5 1 1 28087
0 28089 7 1 2 43343 64611
0 28090 7 1 2 58137 28089
0 28091 5 1 1 28090
0 28092 7 1 2 28088 28091
0 28093 5 1 1 28092
0 28094 7 1 2 42863 28093
0 28095 5 1 1 28094
0 28096 7 1 2 56218 60812
0 28097 5 2 1 28096
0 28098 7 1 2 68688 69912
0 28099 5 1 1 28098
0 28100 7 1 2 59442 28099
0 28101 5 1 1 28100
0 28102 7 1 2 44474 28101
0 28103 7 1 2 28095 28102
0 28104 7 1 2 28084 28103
0 28105 5 1 1 28104
0 28106 7 2 2 66786 28105
0 28107 5 1 1 69914
0 28108 7 2 2 56350 64717
0 28109 5 3 1 69916
0 28110 7 2 2 62132 66575
0 28111 5 1 1 69921
0 28112 7 1 2 69918 28111
0 28113 5 1 1 28112
0 28114 7 1 2 46296 28113
0 28115 5 1 1 28114
0 28116 7 2 2 44684 52899
0 28117 7 1 2 66576 69923
0 28118 5 1 1 28117
0 28119 7 1 2 59620 66546
0 28120 5 1 1 28119
0 28121 7 1 2 28118 28120
0 28122 7 1 2 28115 28121
0 28123 5 1 1 28122
0 28124 7 1 2 50003 28123
0 28125 5 2 1 28124
0 28126 7 2 2 50360 63082
0 28127 5 1 1 69927
0 28128 7 1 2 69919 28127
0 28129 5 1 1 28128
0 28130 7 1 2 43125 28129
0 28131 5 1 1 28130
0 28132 7 1 2 59639 66547
0 28133 5 1 1 28132
0 28134 7 1 2 28131 28133
0 28135 5 1 1 28134
0 28136 7 1 2 46734 28135
0 28137 5 1 1 28136
0 28138 7 1 2 43344 51464
0 28139 7 1 2 68306 28138
0 28140 5 1 1 28139
0 28141 7 2 2 55813 69073
0 28142 5 1 1 69929
0 28143 7 1 2 21342 28142
0 28144 5 2 1 28143
0 28145 7 1 2 42864 69931
0 28146 5 1 1 28145
0 28147 7 1 2 50361 65500
0 28148 7 1 2 51481 28147
0 28149 5 1 1 28148
0 28150 7 1 2 28146 28149
0 28151 7 1 2 28140 28150
0 28152 7 1 2 28137 28151
0 28153 7 1 2 69925 28152
0 28154 5 1 1 28153
0 28155 7 1 2 59731 28154
0 28156 5 1 1 28155
0 28157 7 1 2 28107 28156
0 28158 7 1 2 28068 28157
0 28159 5 1 1 28158
0 28160 7 1 2 44475 28159
0 28161 5 1 1 28160
0 28162 7 2 2 46297 50862
0 28163 5 1 1 69933
0 28164 7 3 2 61837 28163
0 28165 5 1 1 69935
0 28166 7 2 2 66296 69936
0 28167 5 2 1 69938
0 28168 7 1 2 59535 69940
0 28169 5 1 1 28168
0 28170 7 2 2 46298 64553
0 28171 5 1 1 69942
0 28172 7 1 2 59492 69943
0 28173 5 2 1 28172
0 28174 7 1 2 28169 69944
0 28175 5 1 1 28174
0 28176 7 1 2 45609 28175
0 28177 5 1 1 28176
0 28178 7 1 2 67156 69941
0 28179 5 1 1 28178
0 28180 7 1 2 28177 28179
0 28181 5 1 1 28180
0 28182 7 1 2 48640 28181
0 28183 5 1 1 28182
0 28184 7 1 2 64903 67166
0 28185 5 1 1 28184
0 28186 7 1 2 28183 28185
0 28187 5 1 1 28186
0 28188 7 1 2 44085 28187
0 28189 5 1 1 28188
0 28190 7 1 2 50561 64554
0 28191 5 1 1 28190
0 28192 7 1 2 49255 28191
0 28193 5 1 1 28192
0 28194 7 1 2 59493 28193
0 28195 5 1 1 28194
0 28196 7 1 2 50333 58567
0 28197 5 2 1 28196
0 28198 7 1 2 50783 69946
0 28199 5 1 1 28198
0 28200 7 1 2 60222 28199
0 28201 5 2 1 28200
0 28202 7 1 2 59536 69948
0 28203 5 1 1 28202
0 28204 7 1 2 28195 28203
0 28205 5 1 1 28204
0 28206 7 1 2 45610 28205
0 28207 5 1 1 28206
0 28208 7 1 2 67157 69949
0 28209 5 1 1 28208
0 28210 7 1 2 28207 28209
0 28211 5 1 1 28210
0 28212 7 1 2 42865 28211
0 28213 5 1 1 28212
0 28214 7 2 2 49518 57111
0 28215 5 1 1 69950
0 28216 7 1 2 67167 69951
0 28217 5 1 1 28216
0 28218 7 1 2 28213 28217
0 28219 7 1 2 28189 28218
0 28220 5 1 1 28219
0 28221 7 1 2 69915 28220
0 28222 5 1 1 28221
0 28223 7 2 2 47678 67073
0 28224 7 1 2 59943 69952
0 28225 5 1 1 28224
0 28226 7 1 2 20094 28225
0 28227 5 1 1 28226
0 28228 7 1 2 46527 28227
0 28229 5 1 1 28228
0 28230 7 2 2 46299 56842
0 28231 7 1 2 61746 69954
0 28232 5 1 1 28231
0 28233 7 1 2 51732 59917
0 28234 5 2 1 28233
0 28235 7 1 2 28232 69956
0 28236 5 1 1 28235
0 28237 7 1 2 43126 28236
0 28238 5 1 1 28237
0 28239 7 2 2 44086 61747
0 28240 5 1 1 69958
0 28241 7 1 2 59925 28240
0 28242 5 1 1 28241
0 28243 7 1 2 57359 28242
0 28244 5 1 1 28243
0 28245 7 1 2 53501 59918
0 28246 5 2 1 28245
0 28247 7 1 2 28244 69960
0 28248 7 1 2 28238 28247
0 28249 7 1 2 28229 28248
0 28250 5 1 1 28249
0 28251 7 1 2 48641 28250
0 28252 5 1 1 28251
0 28253 7 2 2 59789 63602
0 28254 5 1 1 69962
0 28255 7 1 2 52851 59848
0 28256 5 1 1 28255
0 28257 7 1 2 28254 28256
0 28258 5 1 1 28257
0 28259 7 1 2 43127 28258
0 28260 5 1 1 28259
0 28261 7 2 2 59466 63909
0 28262 7 1 2 48911 69964
0 28263 5 1 1 28262
0 28264 7 1 2 28260 28263
0 28265 5 1 1 28264
0 28266 7 1 2 50863 28265
0 28267 5 1 1 28266
0 28268 7 1 2 61748 68887
0 28269 5 1 1 28268
0 28270 7 1 2 59868 28269
0 28271 5 1 1 28270
0 28272 7 1 2 45286 28271
0 28273 5 1 1 28272
0 28274 7 1 2 69957 28273
0 28275 5 1 1 28274
0 28276 7 1 2 42866 28275
0 28277 5 1 1 28276
0 28278 7 1 2 54716 61749
0 28279 5 1 1 28278
0 28280 7 1 2 59814 28279
0 28281 5 1 1 28280
0 28282 7 1 2 50004 28281
0 28283 5 1 1 28282
0 28284 7 1 2 69961 28283
0 28285 5 1 1 28284
0 28286 7 1 2 43128 28285
0 28287 5 1 1 28286
0 28288 7 1 2 28277 28287
0 28289 7 1 2 28267 28288
0 28290 7 1 2 28252 28289
0 28291 5 1 1 28290
0 28292 7 1 2 66880 28291
0 28293 5 1 1 28292
0 28294 7 1 2 59919 64859
0 28295 5 1 1 28294
0 28296 7 1 2 63906 28295
0 28297 5 1 1 28296
0 28298 7 1 2 50005 28297
0 28299 5 1 1 28298
0 28300 7 2 2 50092 53727
0 28301 5 2 1 69966
0 28302 7 1 2 50616 51879
0 28303 5 2 1 28302
0 28304 7 2 2 54905 69970
0 28305 5 1 1 69972
0 28306 7 1 2 69968 69973
0 28307 5 2 1 28306
0 28308 7 1 2 59920 69974
0 28309 5 1 1 28308
0 28310 7 1 2 28299 28309
0 28311 5 1 1 28310
0 28312 7 1 2 66872 28311
0 28313 5 1 1 28312
0 28314 7 1 2 48823 57561
0 28315 5 3 1 28314
0 28316 7 1 2 63625 69976
0 28317 5 1 1 28316
0 28318 7 1 2 55383 28317
0 28319 5 1 1 28318
0 28320 7 1 2 63621 28319
0 28321 5 1 1 28320
0 28322 7 1 2 66838 28321
0 28323 5 1 1 28322
0 28324 7 1 2 49702 63484
0 28325 5 1 1 28324
0 28326 7 1 2 59642 61990
0 28327 5 1 1 28326
0 28328 7 1 2 28325 28327
0 28329 7 1 2 62041 28328
0 28330 5 1 1 28329
0 28331 7 1 2 66839 28330
0 28332 5 1 1 28331
0 28333 7 1 2 42867 52075
0 28334 5 1 1 28333
0 28335 7 1 2 49791 53874
0 28336 5 4 1 28335
0 28337 7 1 2 48984 49006
0 28338 5 2 1 28337
0 28339 7 1 2 69979 69983
0 28340 7 1 2 28334 28339
0 28341 5 1 1 28340
0 28342 7 1 2 44250 66822
0 28343 7 1 2 28341 28342
0 28344 5 1 1 28343
0 28345 7 1 2 28332 28344
0 28346 5 1 1 28345
0 28347 7 1 2 43345 28346
0 28348 5 1 1 28347
0 28349 7 1 2 65474 68689
0 28350 5 1 1 28349
0 28351 7 1 2 66823 28350
0 28352 5 1 1 28351
0 28353 7 1 2 28348 28352
0 28354 7 1 2 28323 28353
0 28355 5 1 1 28354
0 28356 7 1 2 54793 28355
0 28357 5 1 1 28356
0 28358 7 1 2 28313 28357
0 28359 7 1 2 28293 28358
0 28360 5 1 1 28359
0 28361 7 1 2 53607 28360
0 28362 5 1 1 28361
0 28363 7 1 2 28222 28362
0 28364 7 1 2 28161 28363
0 28365 5 1 1 28364
0 28366 7 1 2 42591 28365
0 28367 5 1 1 28366
0 28368 7 1 2 59206 65444
0 28369 7 2 2 49007 51566
0 28370 7 1 2 68434 69985
0 28371 7 1 2 28368 28370
0 28372 7 1 2 68348 28371
0 28373 5 1 1 28372
0 28374 7 2 2 50362 63219
0 28375 5 1 1 69987
0 28376 7 1 2 58349 69988
0 28377 5 1 1 28376
0 28378 7 1 2 49462 66548
0 28379 5 1 1 28378
0 28380 7 1 2 28377 28379
0 28381 5 2 1 28380
0 28382 7 1 2 43346 69989
0 28383 5 1 1 28382
0 28384 7 3 2 44591 56351
0 28385 7 2 2 63286 69991
0 28386 5 1 1 69994
0 28387 7 1 2 28383 28386
0 28388 5 2 1 28387
0 28389 7 3 2 48642 56240
0 28390 7 1 2 42868 55764
0 28391 7 1 2 63326 28390
0 28392 7 1 2 69998 28391
0 28393 7 1 2 69996 28392
0 28394 5 1 1 28393
0 28395 7 1 2 28373 28394
0 28396 7 1 2 28367 28395
0 28397 5 1 1 28396
0 28398 7 1 2 43758 28397
0 28399 5 1 1 28398
0 28400 7 1 2 57552 64463
0 28401 7 3 2 42057 56201
0 28402 7 1 2 68436 70001
0 28403 7 1 2 28400 28402
0 28404 7 1 2 51810 28403
0 28405 5 1 1 28404
0 28406 7 1 2 28399 28405
0 28407 5 1 1 28406
0 28408 7 1 2 44816 28407
0 28409 5 1 1 28408
0 28410 7 3 2 59665 59760
0 28411 7 1 2 61096 70004
0 28412 5 1 1 28411
0 28413 7 1 2 45477 67168
0 28414 5 1 1 28413
0 28415 7 1 2 28412 28414
0 28416 5 1 1 28415
0 28417 7 1 2 49703 28416
0 28418 5 1 1 28417
0 28419 7 3 2 55804 61281
0 28420 7 1 2 64455 70007
0 28421 5 1 1 28420
0 28422 7 1 2 28418 28421
0 28423 5 1 1 28422
0 28424 7 1 2 51275 28423
0 28425 5 1 1 28424
0 28426 7 2 2 48824 63603
0 28427 7 1 2 57613 58261
0 28428 7 1 2 67887 28427
0 28429 7 1 2 70010 28428
0 28430 5 1 1 28429
0 28431 7 1 2 28425 28430
0 28432 5 1 1 28431
0 28433 7 1 2 66123 28432
0 28434 5 1 1 28433
0 28435 7 1 2 61572 64484
0 28436 5 1 1 28435
0 28437 7 1 2 49008 51298
0 28438 7 1 2 66900 28437
0 28439 5 1 1 28438
0 28440 7 1 2 28436 28439
0 28441 5 1 1 28440
0 28442 7 1 2 69688 28441
0 28443 5 1 1 28442
0 28444 7 1 2 64424 67323
0 28445 5 1 1 28444
0 28446 7 1 2 2705 28445
0 28447 5 1 1 28446
0 28448 7 1 2 44817 28447
0 28449 5 1 1 28448
0 28450 7 1 2 46300 51402
0 28451 7 1 2 64417 28450
0 28452 5 1 1 28451
0 28453 7 1 2 28449 28452
0 28454 5 1 1 28453
0 28455 7 2 2 45857 59522
0 28456 7 3 2 59596 70012
0 28457 7 1 2 57943 70014
0 28458 7 1 2 28454 28457
0 28459 5 1 1 28458
0 28460 7 1 2 28443 28459
0 28461 5 1 1 28460
0 28462 7 1 2 44476 28461
0 28463 5 1 1 28462
0 28464 7 1 2 28434 28463
0 28465 5 1 1 28464
0 28466 7 1 2 47912 28465
0 28467 5 1 1 28466
0 28468 7 1 2 53608 55626
0 28469 7 3 2 63118 63946
0 28470 7 4 2 44685 49009
0 28471 7 1 2 70017 70020
0 28472 7 1 2 28468 28471
0 28473 5 1 1 28472
0 28474 7 1 2 54868 54906
0 28475 5 5 1 28474
0 28476 7 1 2 56352 68269
0 28477 7 1 2 70024 28476
0 28478 7 1 2 58138 28477
0 28479 5 1 1 28478
0 28480 7 1 2 28473 28479
0 28481 5 1 1 28480
0 28482 7 1 2 47679 28481
0 28483 5 1 1 28482
0 28484 7 2 2 48025 51465
0 28485 7 1 2 69166 70029
0 28486 5 1 1 28485
0 28487 7 1 2 28483 28486
0 28488 5 1 1 28487
0 28489 7 1 2 43759 28488
0 28490 5 1 1 28489
0 28491 7 2 2 66989 69174
0 28492 7 1 2 51890 59332
0 28493 7 1 2 61952 28492
0 28494 7 1 2 70031 28493
0 28495 5 1 1 28494
0 28496 7 1 2 28490 28495
0 28497 5 1 1 28496
0 28498 7 1 2 42592 28497
0 28499 5 1 1 28498
0 28500 7 2 2 43554 61292
0 28501 7 1 2 49704 52533
0 28502 7 1 2 70033 28501
0 28503 7 1 2 70032 28502
0 28504 5 1 1 28503
0 28505 7 1 2 28499 28504
0 28506 5 1 1 28505
0 28507 7 1 2 54428 28506
0 28508 5 1 1 28507
0 28509 7 2 2 42336 64541
0 28510 7 1 2 64367 66947
0 28511 5 1 1 28510
0 28512 7 1 2 59999 65642
0 28513 7 1 2 63604 28512
0 28514 5 1 1 28513
0 28515 7 1 2 28511 28514
0 28516 5 1 1 28515
0 28517 7 1 2 45764 28516
0 28518 5 1 1 28517
0 28519 7 1 2 51666 64368
0 28520 5 1 1 28519
0 28521 7 5 2 48643 51595
0 28522 5 1 1 70037
0 28523 7 3 2 45478 70038
0 28524 5 1 1 70042
0 28525 7 1 2 44087 70043
0 28526 5 1 1 28525
0 28527 7 1 2 28520 28526
0 28528 5 1 1 28527
0 28529 7 1 2 60056 28528
0 28530 5 1 1 28529
0 28531 7 1 2 28518 28530
0 28532 5 1 1 28531
0 28533 7 1 2 45611 28532
0 28534 5 1 1 28533
0 28535 7 1 2 58672 64369
0 28536 5 1 1 28535
0 28537 7 1 2 59555 70044
0 28538 5 1 1 28537
0 28539 7 1 2 28536 28538
0 28540 5 1 1 28539
0 28541 7 1 2 46853 28540
0 28542 5 1 1 28541
0 28543 7 1 2 53652 60569
0 28544 7 1 2 61111 28543
0 28545 5 1 1 28544
0 28546 7 1 2 28542 28545
0 28547 5 1 1 28546
0 28548 7 1 2 59369 28547
0 28549 5 1 1 28548
0 28550 7 1 2 28534 28549
0 28551 5 1 1 28550
0 28552 7 1 2 70035 28551
0 28553 5 1 1 28552
0 28554 7 1 2 54794 58830
0 28555 7 1 2 66824 70025
0 28556 7 1 2 28554 28555
0 28557 5 1 1 28556
0 28558 7 1 2 28553 28557
0 28559 5 1 1 28558
0 28560 7 1 2 51310 28559
0 28561 5 1 1 28560
0 28562 7 1 2 28508 28561
0 28563 7 1 2 28467 28562
0 28564 5 1 1 28563
0 28565 7 1 2 55589 28564
0 28566 5 1 1 28565
0 28567 7 1 2 51802 64370
0 28568 5 1 1 28567
0 28569 7 1 2 63877 28568
0 28570 5 1 1 28569
0 28571 7 1 2 63322 66834
0 28572 7 1 2 28570 28571
0 28573 5 1 1 28572
0 28574 7 1 2 63271 64904
0 28575 5 2 1 28574
0 28576 7 5 2 45287 70045
0 28577 5 2 1 70047
0 28578 7 1 2 42869 70048
0 28579 5 1 1 28578
0 28580 7 2 2 61684 28579
0 28581 5 1 1 70054
0 28582 7 1 2 60063 69074
0 28583 7 1 2 28581 28582
0 28584 5 1 1 28583
0 28585 7 1 2 28573 28584
0 28586 5 1 1 28585
0 28587 7 1 2 47131 28586
0 28588 5 1 1 28587
0 28589 7 1 2 58011 59482
0 28590 7 1 2 64663 28589
0 28591 7 1 2 61611 69033
0 28592 7 1 2 28590 28591
0 28593 5 1 1 28592
0 28594 7 1 2 28588 28593
0 28595 5 1 1 28594
0 28596 7 1 2 46071 28595
0 28597 5 1 1 28596
0 28598 7 6 2 46854 45288
0 28599 7 1 2 50214 54503
0 28600 7 1 2 70056 28599
0 28601 7 2 2 47445 63896
0 28602 7 2 2 53858 64305
0 28603 7 1 2 70062 70064
0 28604 7 1 2 28600 28603
0 28605 5 1 1 28604
0 28606 7 1 2 28597 28605
0 28607 5 1 1 28606
0 28608 7 1 2 45612 28607
0 28609 5 1 1 28608
0 28610 7 2 2 50417 59370
0 28611 7 1 2 45479 55991
0 28612 5 1 1 28611
0 28613 7 1 2 63875 28612
0 28614 5 1 1 28613
0 28615 7 1 2 43347 28614
0 28616 5 1 1 28615
0 28617 7 1 2 49705 63518
0 28618 5 1 1 28617
0 28619 7 2 2 48825 55992
0 28620 5 1 1 70068
0 28621 7 1 2 65139 28620
0 28622 5 1 1 28621
0 28623 7 1 2 46735 28622
0 28624 5 1 1 28623
0 28625 7 1 2 28618 28624
0 28626 7 1 2 28616 28625
0 28627 5 1 1 28626
0 28628 7 1 2 68351 28627
0 28629 5 1 1 28628
0 28630 7 3 2 42337 58282
0 28631 7 2 2 47446 51567
0 28632 7 1 2 70070 70073
0 28633 5 1 1 28632
0 28634 7 5 2 54504 65831
0 28635 5 1 1 70075
0 28636 7 1 2 28633 28635
0 28637 5 1 1 28636
0 28638 7 1 2 60715 28637
0 28639 5 1 1 28638
0 28640 7 3 2 48026 51803
0 28641 7 1 2 56861 63832
0 28642 7 1 2 70080 28641
0 28643 5 1 1 28642
0 28644 7 2 2 43348 63220
0 28645 7 1 2 54463 66110
0 28646 7 1 2 70083 28645
0 28647 5 1 1 28646
0 28648 7 1 2 28643 28647
0 28649 7 1 2 28639 28648
0 28650 5 1 1 28649
0 28651 7 1 2 45289 28650
0 28652 5 1 1 28651
0 28653 7 1 2 49180 53792
0 28654 5 1 1 28653
0 28655 7 2 2 57999 28165
0 28656 7 1 2 48644 70085
0 28657 5 1 1 28656
0 28658 7 1 2 28654 28657
0 28659 5 1 1 28658
0 28660 7 1 2 70076 28659
0 28661 5 1 1 28660
0 28662 7 1 2 28652 28661
0 28663 7 1 2 28629 28662
0 28664 5 1 1 28663
0 28665 7 1 2 70066 28664
0 28666 5 1 1 28665
0 28667 7 1 2 47797 28666
0 28668 7 1 2 28609 28667
0 28669 5 1 1 28668
0 28670 7 1 2 52900 54847
0 28671 5 1 1 28670
0 28672 7 2 2 43760 68565
0 28673 5 1 1 70087
0 28674 7 1 2 28671 28673
0 28675 5 2 1 28674
0 28676 7 1 2 46072 70089
0 28677 5 1 1 28676
0 28678 7 1 2 53200 68566
0 28679 5 1 1 28678
0 28680 7 1 2 28677 28679
0 28681 5 2 1 28680
0 28682 7 1 2 65870 70091
0 28683 5 1 1 28682
0 28684 7 1 2 55009 7560
0 28685 5 1 1 28684
0 28686 7 1 2 46528 28685
0 28687 5 1 1 28686
0 28688 7 1 2 69980 28687
0 28689 5 1 1 28688
0 28690 7 1 2 50006 28689
0 28691 5 1 1 28690
0 28692 7 2 2 50956 60439
0 28693 5 1 1 70093
0 28694 7 2 2 48645 70094
0 28695 5 1 1 70095
0 28696 7 1 2 28691 28695
0 28697 5 1 1 28696
0 28698 7 1 2 50418 54795
0 28699 7 1 2 28697 28698
0 28700 5 1 1 28699
0 28701 7 1 2 28683 28700
0 28702 5 1 1 28701
0 28703 7 1 2 66410 28702
0 28704 5 1 1 28703
0 28705 7 1 2 51061 58644
0 28706 7 2 2 55278 28705
0 28707 5 1 1 70097
0 28708 7 1 2 46301 70098
0 28709 5 2 1 28708
0 28710 7 1 2 45480 70088
0 28711 5 1 1 28710
0 28712 7 1 2 42870 57210
0 28713 7 1 2 59802 28712
0 28714 5 1 1 28713
0 28715 7 1 2 28711 28714
0 28716 5 1 1 28715
0 28717 7 1 2 47578 28716
0 28718 5 1 1 28717
0 28719 7 1 2 59041 63605
0 28720 5 1 1 28719
0 28721 7 1 2 56219 57602
0 28722 5 1 1 28721
0 28723 7 1 2 28720 28722
0 28724 5 1 1 28723
0 28725 7 1 2 47132 28724
0 28726 5 1 1 28725
0 28727 7 1 2 28718 28726
0 28728 5 1 1 28727
0 28729 7 1 2 46073 28728
0 28730 5 1 1 28729
0 28731 7 1 2 70099 28730
0 28732 5 1 1 28731
0 28733 7 3 2 51568 66415
0 28734 7 1 2 28732 70101
0 28735 5 1 1 28734
0 28736 7 1 2 28704 28735
0 28737 5 1 1 28736
0 28738 7 1 2 47680 28737
0 28739 5 1 1 28738
0 28740 7 1 2 51709 63915
0 28741 5 2 1 28740
0 28742 7 2 2 64411 70104
0 28743 7 1 2 42871 51447
0 28744 5 1 1 28743
0 28745 7 1 2 25905 28744
0 28746 7 1 2 70106 28745
0 28747 5 1 1 28746
0 28748 7 9 2 48027 66868
0 28749 7 1 2 50419 59849
0 28750 7 1 2 70108 28749
0 28751 7 1 2 28747 28750
0 28752 5 1 1 28751
0 28753 7 1 2 44477 28752
0 28754 7 1 2 28739 28753
0 28755 5 1 1 28754
0 28756 7 1 2 53609 28755
0 28757 7 1 2 28669 28756
0 28758 5 1 1 28757
0 28759 7 1 2 46736 53793
0 28760 7 1 2 58673 28759
0 28761 5 1 1 28760
0 28762 7 1 2 56526 59300
0 28763 5 1 1 28762
0 28764 7 1 2 28761 28763
0 28765 5 1 1 28764
0 28766 7 1 2 69198 28765
0 28767 5 1 1 28766
0 28768 7 3 2 60644 61872
0 28769 7 1 2 55993 70117
0 28770 5 1 1 28769
0 28771 7 1 2 55384 64228
0 28772 5 1 1 28771
0 28773 7 1 2 28770 28772
0 28774 5 1 1 28773
0 28775 7 1 2 53676 28774
0 28776 5 1 1 28775
0 28777 7 6 2 43555 47447
0 28778 7 2 2 60645 70120
0 28779 7 1 2 61861 70126
0 28780 5 1 1 28779
0 28781 7 1 2 61595 62515
0 28782 7 1 2 52901 28781
0 28783 7 1 2 64390 28782
0 28784 5 1 1 28783
0 28785 7 1 2 28780 28784
0 28786 5 1 1 28785
0 28787 7 1 2 42872 28786
0 28788 5 1 1 28787
0 28789 7 4 2 43556 44088
0 28790 7 2 2 64198 70128
0 28791 7 1 2 61862 61928
0 28792 7 1 2 70132 28791
0 28793 5 1 1 28792
0 28794 7 1 2 28788 28793
0 28795 7 1 2 28776 28794
0 28796 5 1 1 28795
0 28797 7 1 2 47913 28796
0 28798 5 1 1 28797
0 28799 7 1 2 53610 69059
0 28800 7 2 2 61106 28799
0 28801 7 1 2 47798 53794
0 28802 7 1 2 70134 28801
0 28803 5 1 1 28802
0 28804 7 1 2 28798 28803
0 28805 5 1 1 28804
0 28806 7 1 2 69075 28805
0 28807 5 1 1 28806
0 28808 7 1 2 28767 28807
0 28809 5 1 1 28808
0 28810 7 1 2 47133 28809
0 28811 5 1 1 28810
0 28812 7 5 2 47448 63088
0 28813 7 1 2 53611 66886
0 28814 5 1 1 28813
0 28815 7 1 2 58754 66500
0 28816 5 1 1 28815
0 28817 7 1 2 28814 28816
0 28818 5 1 1 28817
0 28819 7 1 2 46855 28818
0 28820 5 1 1 28819
0 28821 7 3 2 43477 63801
0 28822 7 2 2 58910 70141
0 28823 5 1 1 70144
0 28824 7 1 2 56427 70145
0 28825 5 1 1 28824
0 28826 7 1 2 28820 28825
0 28827 5 1 1 28826
0 28828 7 1 2 45613 28827
0 28829 5 1 1 28828
0 28830 7 1 2 58428 68282
0 28831 5 1 1 28830
0 28832 7 1 2 28829 28831
0 28833 5 1 1 28832
0 28834 7 2 2 70136 28833
0 28835 7 2 2 54976 60138
0 28836 7 1 2 70146 70148
0 28837 5 1 1 28836
0 28838 7 1 2 28811 28837
0 28839 5 1 1 28838
0 28840 7 1 2 46074 28839
0 28841 5 1 1 28840
0 28842 7 1 2 57211 68734
0 28843 7 1 2 70147 28842
0 28844 5 1 1 28843
0 28845 7 1 2 28841 28844
0 28846 5 1 1 28845
0 28847 7 1 2 49091 28846
0 28848 5 1 1 28847
0 28849 7 1 2 63606 69869
0 28850 5 2 1 28849
0 28851 7 1 2 60852 65477
0 28852 5 2 1 28851
0 28853 7 1 2 69864 70152
0 28854 5 1 1 28853
0 28855 7 1 2 70150 28854
0 28856 5 1 1 28855
0 28857 7 1 2 57380 28856
0 28858 5 1 1 28857
0 28859 7 2 2 58922 59443
0 28860 7 1 2 54848 58792
0 28861 7 1 2 70154 28860
0 28862 5 1 1 28861
0 28863 7 1 2 28858 28862
0 28864 5 1 1 28863
0 28865 7 1 2 46529 28864
0 28866 5 1 1 28865
0 28867 7 1 2 43349 62234
0 28868 5 1 1 28867
0 28869 7 1 2 57453 28868
0 28870 5 1 1 28869
0 28871 7 1 2 52790 28870
0 28872 5 1 1 28871
0 28873 7 3 2 45765 57353
0 28874 7 1 2 46940 60580
0 28875 7 1 2 70156 28874
0 28876 5 1 1 28875
0 28877 7 1 2 28872 28876
0 28878 5 1 1 28877
0 28879 7 1 2 44349 28878
0 28880 5 1 1 28879
0 28881 7 1 2 57619 60593
0 28882 5 1 1 28881
0 28883 7 1 2 28880 28882
0 28884 5 1 1 28883
0 28885 7 1 2 49706 28884
0 28886 5 1 1 28885
0 28887 7 2 2 55849 59207
0 28888 7 1 2 42226 55385
0 28889 7 1 2 70159 28888
0 28890 5 1 1 28889
0 28891 7 1 2 28886 28890
0 28892 5 1 1 28891
0 28893 7 1 2 42058 28892
0 28894 5 1 1 28893
0 28895 7 1 2 60604 61944
0 28896 5 1 1 28895
0 28897 7 1 2 52791 28896
0 28898 5 1 1 28897
0 28899 7 4 2 46941 59160
0 28900 7 1 2 64809 70161
0 28901 5 1 1 28900
0 28902 7 1 2 28898 28901
0 28903 5 1 1 28902
0 28904 7 1 2 49707 61082
0 28905 7 1 2 28903 28904
0 28906 5 1 1 28905
0 28907 7 1 2 28894 28906
0 28908 5 1 1 28907
0 28909 7 1 2 47134 28908
0 28910 5 1 1 28909
0 28911 7 1 2 28866 28910
0 28912 5 1 1 28911
0 28913 7 1 2 46075 28912
0 28914 5 1 1 28913
0 28915 7 1 2 56918 58116
0 28916 7 1 2 61083 63089
0 28917 7 1 2 64605 28916
0 28918 7 1 2 28915 28917
0 28919 5 1 1 28918
0 28920 7 1 2 70151 28919
0 28921 5 1 1 28920
0 28922 7 1 2 50709 61246
0 28923 7 1 2 28921 28922
0 28924 5 1 1 28923
0 28925 7 1 2 28914 28924
0 28926 5 1 1 28925
0 28927 7 1 2 66787 28926
0 28928 5 1 1 28927
0 28929 7 1 2 49181 70090
0 28930 5 1 1 28929
0 28931 7 1 2 61536 69981
0 28932 5 1 1 28931
0 28933 7 1 2 51710 28932
0 28934 5 1 1 28933
0 28935 7 1 2 51482 57360
0 28936 5 1 1 28935
0 28937 7 1 2 28934 28936
0 28938 5 1 1 28937
0 28939 7 1 2 47135 28938
0 28940 5 1 1 28939
0 28941 7 1 2 28930 28940
0 28942 5 1 1 28941
0 28943 7 1 2 46076 28942
0 28944 5 1 1 28943
0 28945 7 1 2 70100 28944
0 28946 5 1 1 28945
0 28947 7 1 2 59444 28946
0 28948 5 1 1 28947
0 28949 7 1 2 43129 52400
0 28950 5 1 1 28949
0 28951 7 1 2 63912 28950
0 28952 5 1 1 28951
0 28953 7 1 2 50007 28952
0 28954 5 1 1 28953
0 28955 7 1 2 49631 53728
0 28956 5 1 1 28955
0 28957 7 1 2 28954 28956
0 28958 5 1 1 28957
0 28959 7 1 2 47136 28958
0 28960 5 1 1 28959
0 28961 7 3 2 50334 51403
0 28962 5 1 1 70165
0 28963 7 1 2 57361 70166
0 28964 5 1 1 28963
0 28965 7 1 2 28960 28964
0 28966 5 1 1 28965
0 28967 7 1 2 46077 28966
0 28968 5 1 1 28967
0 28969 7 1 2 56220 57248
0 28970 7 1 2 57711 28969
0 28971 5 1 1 28970
0 28972 7 1 2 28968 28971
0 28973 5 1 1 28972
0 28974 7 1 2 59732 28973
0 28975 5 1 1 28974
0 28976 7 1 2 28948 28975
0 28977 5 1 1 28976
0 28978 7 1 2 68361 28977
0 28979 5 1 1 28978
0 28980 7 2 2 47681 54896
0 28981 7 1 2 66549 70168
0 28982 7 1 2 58139 28981
0 28983 5 1 1 28982
0 28984 7 1 2 50363 50617
0 28985 7 1 2 70015 28984
0 28986 5 1 1 28985
0 28987 7 1 2 28983 28986
0 28988 5 1 1 28987
0 28989 7 1 2 52510 28988
0 28990 5 1 1 28989
0 28991 7 6 2 47449 44592
0 28992 7 2 2 63090 70170
0 28993 7 2 2 68299 70176
0 28994 7 1 2 51102 64116
0 28995 7 1 2 70178 28994
0 28996 5 1 1 28995
0 28997 7 1 2 28990 28996
0 28998 5 1 1 28997
0 28999 7 1 2 46078 28998
0 29000 5 1 1 28999
0 29001 7 1 2 64673 64464
0 29002 7 1 2 70179 29001
0 29003 5 1 1 29002
0 29004 7 1 2 29000 29003
0 29005 5 1 1 29004
0 29006 7 1 2 50093 29005
0 29007 5 1 1 29006
0 29008 7 1 2 47137 48970
0 29009 7 1 2 61463 29008
0 29010 5 1 1 29009
0 29011 7 1 2 50472 51466
0 29012 5 1 1 29011
0 29013 7 1 2 49051 51181
0 29014 7 1 2 29012 29013
0 29015 5 1 1 29014
0 29016 7 1 2 29010 29015
0 29017 5 1 1 29016
0 29018 7 1 2 46302 29017
0 29019 5 1 1 29018
0 29020 7 1 2 50420 1005
0 29021 5 1 1 29020
0 29022 7 1 2 29019 29021
0 29023 5 1 1 29022
0 29024 7 3 2 44593 59681
0 29025 7 1 2 64647 68391
0 29026 7 1 2 70180 29025
0 29027 7 1 2 29023 29026
0 29028 5 1 1 29027
0 29029 7 1 2 29007 29028
0 29030 7 1 2 28979 29029
0 29031 5 1 1 29030
0 29032 7 1 2 44478 29031
0 29033 5 1 1 29032
0 29034 7 1 2 54849 58481
0 29035 5 1 1 29034
0 29036 7 1 2 52321 61334
0 29037 5 1 1 29036
0 29038 7 1 2 29035 29037
0 29039 5 1 1 29038
0 29040 7 1 2 69613 29039
0 29041 5 1 1 29040
0 29042 7 2 2 57019 66463
0 29043 7 1 2 53281 61439
0 29044 7 1 2 70183 29043
0 29045 7 1 2 58140 29044
0 29046 5 1 1 29045
0 29047 7 1 2 29041 29046
0 29048 5 1 1 29047
0 29049 7 1 2 44594 29048
0 29050 5 1 1 29049
0 29051 7 2 2 54850 63292
0 29052 7 1 2 50364 70185
0 29053 7 1 2 59050 29052
0 29054 5 1 1 29053
0 29055 7 1 2 29050 29054
0 29056 5 1 1 29055
0 29057 7 1 2 59161 29056
0 29058 5 1 1 29057
0 29059 7 1 2 53282 68475
0 29060 7 1 2 70184 29059
0 29061 7 1 2 66596 29060
0 29062 5 1 1 29061
0 29063 7 1 2 29058 29062
0 29064 5 1 1 29063
0 29065 7 1 2 45290 29064
0 29066 5 1 1 29065
0 29067 7 1 2 58935 68673
0 29068 7 2 2 47138 59604
0 29069 7 2 2 57786 57918
0 29070 7 1 2 70187 70189
0 29071 7 1 2 29067 29070
0 29072 5 1 1 29071
0 29073 7 1 2 29066 29072
0 29074 5 1 1 29073
0 29075 7 1 2 51024 29074
0 29076 5 1 1 29075
0 29077 7 1 2 44089 62183
0 29078 5 1 1 29077
0 29079 7 1 2 58339 29078
0 29080 5 1 1 29079
0 29081 7 1 2 68134 29080
0 29082 5 1 1 29081
0 29083 7 1 2 56989 61838
0 29084 5 1 1 29083
0 29085 7 1 2 44090 29084
0 29086 5 1 1 29085
0 29087 7 1 2 53410 55481
0 29088 5 1 1 29087
0 29089 7 1 2 50784 29088
0 29090 5 1 1 29089
0 29091 7 1 2 29086 29090
0 29092 5 1 1 29091
0 29093 7 1 2 66550 29092
0 29094 5 1 1 29093
0 29095 7 1 2 29082 29094
0 29096 5 1 1 29095
0 29097 7 1 2 48646 29096
0 29098 5 1 1 29097
0 29099 7 1 2 50785 61699
0 29100 5 1 1 29099
0 29101 7 1 2 50864 61991
0 29102 5 1 1 29101
0 29103 7 1 2 53844 29102
0 29104 7 1 2 29100 29103
0 29105 5 1 1 29104
0 29106 7 1 2 66551 29105
0 29107 5 1 1 29106
0 29108 7 1 2 55424 60077
0 29109 7 1 2 68428 29108
0 29110 5 1 1 29109
0 29111 7 1 2 29107 29110
0 29112 7 1 2 29098 29111
0 29113 5 1 1 29112
0 29114 7 1 2 67169 29113
0 29115 5 1 1 29114
0 29116 7 1 2 53313 69963
0 29117 7 1 2 69997 29116
0 29118 5 1 1 29117
0 29119 7 1 2 29115 29118
0 29120 5 1 1 29119
0 29121 7 1 2 63331 29120
0 29122 5 1 1 29121
0 29123 7 1 2 29076 29122
0 29124 7 1 2 29033 29123
0 29125 7 1 2 28928 29124
0 29126 7 1 2 28848 29125
0 29127 7 1 2 28758 29126
0 29128 5 1 1 29127
0 29129 7 1 2 48140 29128
0 29130 5 1 1 29129
0 29131 7 1 2 28566 29130
0 29132 7 1 2 28409 29131
0 29133 5 1 1 29132
0 29134 7 1 2 66277 29133
0 29135 5 1 1 29134
0 29136 7 1 2 64025 69369
0 29137 5 1 1 29136
0 29138 7 1 2 68503 29137
0 29139 5 3 1 29138
0 29140 7 1 2 61531 68059
0 29141 7 4 2 61272 66140
0 29142 7 2 2 46856 69429
0 29143 7 1 2 70194 70198
0 29144 7 1 2 29140 29143
0 29145 7 1 2 70191 29144
0 29146 5 1 1 29145
0 29147 7 2 2 47139 65704
0 29148 7 1 2 61574 65591
0 29149 5 1 1 29148
0 29150 7 2 2 70200 29149
0 29151 5 1 1 70202
0 29152 7 1 2 62350 27526
0 29153 5 4 1 29152
0 29154 7 2 2 55107 70204
0 29155 7 1 2 69439 70208
0 29156 5 1 1 29155
0 29157 7 1 2 29151 29156
0 29158 5 1 1 29157
0 29159 7 1 2 44479 66228
0 29160 7 1 2 29158 29159
0 29161 5 1 1 29160
0 29162 7 1 2 29146 29161
0 29163 5 1 1 29162
0 29164 7 1 2 54082 29163
0 29165 5 1 1 29164
0 29166 7 1 2 57317 57829
0 29167 5 1 1 29166
0 29168 7 1 2 54897 29167
0 29169 5 1 1 29168
0 29170 7 1 2 44091 58375
0 29171 5 1 1 29170
0 29172 7 1 2 65471 29171
0 29173 5 1 1 29172
0 29174 7 1 2 46530 29173
0 29175 5 1 1 29174
0 29176 7 1 2 61547 69904
0 29177 7 1 2 29175 29176
0 29178 5 1 1 29177
0 29179 7 1 2 48647 29178
0 29180 5 1 1 29179
0 29181 7 2 2 69913 29180
0 29182 5 1 1 70210
0 29183 7 1 2 29169 70211
0 29184 5 1 1 29183
0 29185 7 1 2 66200 67840
0 29186 7 1 2 29184 29185
0 29187 5 1 1 29186
0 29188 7 2 2 51733 3481
0 29189 7 2 2 63947 70212
0 29190 5 2 1 70214
0 29191 7 1 2 46303 62956
0 29192 5 1 1 29191
0 29193 7 1 2 70216 29192
0 29194 5 1 1 29193
0 29195 7 2 2 48648 29194
0 29196 5 1 1 70218
0 29197 7 2 2 63833 66167
0 29198 7 2 2 58950 70220
0 29199 7 1 2 70219 70222
0 29200 5 1 1 29199
0 29201 7 1 2 29187 29200
0 29202 5 1 1 29201
0 29203 7 1 2 57197 29202
0 29204 5 1 1 29203
0 29205 7 1 2 45481 70223
0 29206 5 1 1 29205
0 29207 7 4 2 44480 66201
0 29208 7 2 2 66004 70224
0 29209 5 1 1 70228
0 29210 7 1 2 29206 29209
0 29211 5 1 1 29210
0 29212 7 1 2 50094 29211
0 29213 5 1 1 29212
0 29214 7 1 2 58811 66168
0 29215 7 1 2 65806 29214
0 29216 5 1 1 29215
0 29217 7 1 2 29213 29216
0 29218 5 1 1 29217
0 29219 7 1 2 49301 29218
0 29220 5 1 1 29219
0 29221 7 1 2 57381 70229
0 29222 5 1 1 29221
0 29223 7 1 2 29220 29222
0 29224 5 1 1 29223
0 29225 7 4 2 47140 51025
0 29226 7 1 2 68920 70230
0 29227 7 1 2 29224 29226
0 29228 5 1 1 29227
0 29229 7 1 2 29204 29228
0 29230 5 1 1 29229
0 29231 7 1 2 45614 29230
0 29232 5 1 1 29231
0 29233 7 2 2 44481 66225
0 29234 7 1 2 54099 57429
0 29235 5 1 1 29234
0 29236 7 1 2 54321 57198
0 29237 5 1 1 29236
0 29238 7 1 2 29235 29237
0 29239 5 1 1 29238
0 29240 7 1 2 51026 29239
0 29241 5 1 1 29240
0 29242 7 3 2 44818 54536
0 29243 7 1 2 57312 70236
0 29244 5 1 1 29243
0 29245 7 1 2 50095 54977
0 29246 7 1 2 64418 29245
0 29247 5 1 1 29246
0 29248 7 1 2 29244 29247
0 29249 7 1 2 29241 29248
0 29250 5 1 1 29249
0 29251 7 1 2 65915 29250
0 29252 5 1 1 29251
0 29253 7 1 2 57223 68397
0 29254 7 1 2 70205 29253
0 29255 5 1 1 29254
0 29256 7 1 2 29252 29255
0 29257 5 1 1 29256
0 29258 7 1 2 45291 29257
0 29259 5 1 1 29258
0 29260 7 1 2 57199 65916
0 29261 7 1 2 29182 29260
0 29262 5 1 1 29261
0 29263 7 1 2 29259 29262
0 29264 5 1 1 29263
0 29265 7 1 2 70234 29264
0 29266 5 1 1 29265
0 29267 7 1 2 29232 29266
0 29268 5 1 1 29267
0 29269 7 1 2 42593 29268
0 29270 5 1 1 29269
0 29271 7 1 2 29165 29270
0 29272 5 1 1 29271
0 29273 7 1 2 47682 29272
0 29274 5 1 1 29273
0 29275 7 1 2 46304 57817
0 29276 5 1 1 29275
0 29277 7 3 2 44482 69418
0 29278 7 1 2 29276 70239
0 29279 5 1 1 29278
0 29280 7 5 2 66068 67815
0 29281 7 1 2 48649 62235
0 29282 5 1 1 29281
0 29283 7 1 2 3012 29282
0 29284 5 1 1 29283
0 29285 7 1 2 70242 29284
0 29286 5 1 1 29285
0 29287 7 1 2 64446 64199
0 29288 7 1 2 66169 29287
0 29289 5 1 1 29288
0 29290 7 1 2 29286 29289
0 29291 5 1 1 29290
0 29292 7 1 2 50008 29291
0 29293 5 1 1 29292
0 29294 7 1 2 29279 29293
0 29295 5 1 1 29294
0 29296 7 1 2 65705 29295
0 29297 5 1 1 29296
0 29298 7 1 2 46737 62427
0 29299 5 1 1 29298
0 29300 7 1 2 51804 58577
0 29301 5 1 1 29300
0 29302 7 1 2 49925 57090
0 29303 5 1 1 29302
0 29304 7 1 2 29301 29303
0 29305 7 1 2 29299 29304
0 29306 5 1 1 29305
0 29307 7 1 2 65917 69466
0 29308 7 1 2 69481 29307
0 29309 7 1 2 29306 29308
0 29310 5 1 1 29309
0 29311 7 1 2 29297 29310
0 29312 5 1 1 29311
0 29313 7 1 2 42594 29312
0 29314 5 1 1 29313
0 29315 7 3 2 48650 65918
0 29316 5 1 1 70247
0 29317 7 1 2 59111 70248
0 29318 5 1 1 29317
0 29319 7 1 2 49543 69710
0 29320 5 1 1 29319
0 29321 7 1 2 29318 29320
0 29322 5 1 1 29321
0 29323 7 1 2 59556 66359
0 29324 7 1 2 67197 29323
0 29325 7 1 2 29322 29324
0 29326 5 1 1 29325
0 29327 7 1 2 29314 29326
0 29328 5 1 1 29327
0 29329 7 1 2 43761 29328
0 29330 5 1 1 29329
0 29331 7 2 2 49554 52337
0 29332 7 1 2 65919 70250
0 29333 5 1 1 29332
0 29334 7 1 2 49544 65706
0 29335 5 2 1 29334
0 29336 7 1 2 29333 70252
0 29337 5 1 1 29336
0 29338 7 2 2 54401 69419
0 29339 7 1 2 63276 70254
0 29340 7 1 2 29337 29339
0 29341 5 1 1 29340
0 29342 7 1 2 29330 29341
0 29343 5 1 1 29342
0 29344 7 1 2 42059 29343
0 29345 5 1 1 29344
0 29346 7 1 2 58951 63423
0 29347 7 1 2 65041 29346
0 29348 7 2 2 51145 66384
0 29349 7 1 2 68697 70256
0 29350 7 1 2 29347 29349
0 29351 5 1 1 29350
0 29352 7 1 2 44819 29351
0 29353 7 1 2 29345 29352
0 29354 5 1 1 29353
0 29355 7 1 2 60159 70243
0 29356 5 1 1 29355
0 29357 7 1 2 63335 66170
0 29358 5 1 1 29357
0 29359 7 1 2 29356 29358
0 29360 5 1 1 29359
0 29361 7 1 2 42060 29360
0 29362 5 1 1 29361
0 29363 7 1 2 66069 69485
0 29364 5 1 1 29363
0 29365 7 1 2 29362 29364
0 29366 5 1 1 29365
0 29367 7 1 2 50786 53795
0 29368 5 2 1 29367
0 29369 7 1 2 300 70258
0 29370 5 1 1 29369
0 29371 7 1 2 47799 29370
0 29372 7 1 2 29366 29371
0 29373 5 1 1 29372
0 29374 7 1 2 46305 60196
0 29375 5 1 1 29374
0 29376 7 1 2 50562 63511
0 29377 5 1 1 29376
0 29378 7 2 2 29375 29377
0 29379 5 1 1 70260
0 29380 7 2 2 46531 29379
0 29381 5 1 1 70262
0 29382 7 1 2 49052 3501
0 29383 5 1 1 29382
0 29384 7 1 2 25703 29383
0 29385 5 1 1 29384
0 29386 7 1 2 43350 29385
0 29387 5 1 1 29386
0 29388 7 1 2 46738 69394
0 29389 5 1 1 29388
0 29390 7 1 2 63534 29389
0 29391 7 1 2 29387 29390
0 29392 5 1 1 29391
0 29393 7 1 2 46079 29392
0 29394 5 1 1 29393
0 29395 7 1 2 51467 51805
0 29396 7 1 2 60949 64520
0 29397 7 1 2 29395 29396
0 29398 5 1 1 29397
0 29399 7 1 2 29394 29398
0 29400 7 1 2 29381 29399
0 29401 5 1 1 29400
0 29402 7 1 2 69462 29401
0 29403 5 1 1 29402
0 29404 7 1 2 29373 29403
0 29405 5 1 1 29404
0 29406 7 1 2 65707 29405
0 29407 5 1 1 29406
0 29408 7 1 2 57354 70167
0 29409 5 1 1 29408
0 29410 7 1 2 46080 49545
0 29411 5 1 1 29410
0 29412 7 1 2 70261 29411
0 29413 5 1 1 29412
0 29414 7 1 2 46532 29413
0 29415 5 1 1 29414
0 29416 7 1 2 29409 29415
0 29417 5 1 1 29416
0 29418 7 2 2 63424 66734
0 29419 7 1 2 43647 48028
0 29420 7 1 2 61768 29419
0 29421 7 1 2 70264 29420
0 29422 7 1 2 29417 29421
0 29423 5 1 1 29422
0 29424 7 1 2 29407 29423
0 29425 5 1 1 29424
0 29426 7 1 2 47141 29425
0 29427 5 1 1 29426
0 29428 7 2 2 50421 66385
0 29429 7 2 2 43603 70266
0 29430 7 1 2 56241 58929
0 29431 7 1 2 66970 29430
0 29432 7 1 2 70268 29431
0 29433 5 1 1 29432
0 29434 7 1 2 42061 66202
0 29435 5 1 1 29434
0 29436 7 1 2 25359 29435
0 29437 5 6 1 29436
0 29438 7 1 2 57415 65438
0 29439 7 1 2 62622 29438
0 29440 7 1 2 70270 29439
0 29441 5 1 1 29440
0 29442 7 1 2 29433 29441
0 29443 5 1 1 29442
0 29444 7 1 2 51027 29443
0 29445 5 1 1 29444
0 29446 7 1 2 61769 68245
0 29447 7 1 2 66005 67504
0 29448 7 1 2 29446 29447
0 29449 7 1 2 70263 29448
0 29450 5 1 1 29449
0 29451 7 1 2 48141 29450
0 29452 7 1 2 29445 29451
0 29453 7 1 2 29427 29452
0 29454 5 1 1 29453
0 29455 7 1 2 44350 29454
0 29456 7 1 2 29354 29455
0 29457 5 1 1 29456
0 29458 7 5 2 44351 70271
0 29459 7 1 2 50787 61722
0 29460 5 1 1 29459
0 29461 7 1 2 48651 17261
0 29462 5 1 1 29461
0 29463 7 1 2 29460 29462
0 29464 5 1 1 29463
0 29465 7 1 2 70276 29464
0 29466 5 1 1 29465
0 29467 7 1 2 53746 67074
0 29468 5 2 1 29467
0 29469 7 1 2 28171 70281
0 29470 5 1 1 29469
0 29471 7 18 2 59483 66171
0 29472 7 1 2 45615 48652
0 29473 7 1 2 70283 29472
0 29474 7 1 2 29470 29473
0 29475 5 1 1 29474
0 29476 7 1 2 29466 29475
0 29477 5 1 1 29476
0 29478 7 1 2 65920 29477
0 29479 5 1 1 29478
0 29480 7 1 2 61784 66215
0 29481 7 2 2 44251 61742
0 29482 7 1 2 68219 70301
0 29483 7 1 2 29480 29482
0 29484 5 1 1 29483
0 29485 7 1 2 57990 58578
0 29486 7 1 2 70277 29485
0 29487 5 1 1 29486
0 29488 7 1 2 29484 29487
0 29489 5 1 1 29488
0 29490 7 1 2 65708 29489
0 29491 5 1 1 29490
0 29492 7 1 2 29479 29491
0 29493 5 1 1 29492
0 29494 7 1 2 44092 29493
0 29495 5 1 1 29494
0 29496 7 1 2 63916 66971
0 29497 5 1 1 29496
0 29498 7 1 2 63599 64362
0 29499 5 3 1 29498
0 29500 7 2 2 48029 70303
0 29501 7 1 2 45858 70306
0 29502 5 1 1 29501
0 29503 7 1 2 29497 29502
0 29504 5 1 1 29503
0 29505 7 1 2 70278 29504
0 29506 5 1 1 29505
0 29507 7 5 2 62904 65859
0 29508 7 2 2 54222 70308
0 29509 7 1 2 60078 63091
0 29510 7 1 2 64037 29509
0 29511 7 1 2 70313 29510
0 29512 5 1 1 29511
0 29513 7 1 2 29506 29512
0 29514 5 1 1 29513
0 29515 7 1 2 50865 29514
0 29516 5 1 1 29515
0 29517 7 1 2 49519 68989
0 29518 5 1 1 29517
0 29519 7 1 2 46533 69453
0 29520 5 1 1 29519
0 29521 7 1 2 29518 29520
0 29522 5 1 1 29521
0 29523 7 1 2 50009 29522
0 29524 5 1 1 29523
0 29525 7 1 2 58579 64026
0 29526 7 1 2 69742 29525
0 29527 5 1 1 29526
0 29528 7 1 2 26908 29527
0 29529 5 1 1 29528
0 29530 7 1 2 42873 29529
0 29531 5 1 1 29530
0 29532 7 1 2 57991 65709
0 29533 5 1 1 29532
0 29534 7 1 2 57656 66100
0 29535 5 1 1 29534
0 29536 7 1 2 29533 29535
0 29537 7 1 2 29531 29536
0 29538 5 1 1 29537
0 29539 7 1 2 64856 29538
0 29540 5 1 1 29539
0 29541 7 1 2 29524 29540
0 29542 5 1 1 29541
0 29543 7 1 2 70279 29542
0 29544 5 1 1 29543
0 29545 7 1 2 65710 68888
0 29546 5 1 1 29545
0 29547 7 3 2 45859 62067
0 29548 7 1 2 62355 70315
0 29549 5 1 1 29548
0 29550 7 1 2 29546 29549
0 29551 5 1 1 29550
0 29552 7 1 2 48826 29551
0 29553 5 2 1 29552
0 29554 7 1 2 43351 61464
0 29555 7 1 2 65803 29554
0 29556 5 1 1 29555
0 29557 7 1 2 70318 29556
0 29558 5 1 1 29557
0 29559 7 1 2 61273 70169
0 29560 7 1 2 70309 29559
0 29561 7 1 2 29558 29560
0 29562 5 1 1 29561
0 29563 7 1 2 29544 29562
0 29564 7 1 2 29516 29563
0 29565 7 1 2 29495 29564
0 29566 5 1 1 29565
0 29567 7 1 2 47800 29566
0 29568 5 1 1 29567
0 29569 7 1 2 49053 12721
0 29570 5 1 1 29569
0 29571 7 1 2 43352 52836
0 29572 7 1 2 9698 29571
0 29573 7 1 2 29570 29572
0 29574 5 1 1 29573
0 29575 7 1 2 46739 53720
0 29576 5 1 1 29575
0 29577 7 2 2 48030 67522
0 29578 7 1 2 56242 70265
0 29579 7 1 2 70320 29578
0 29580 7 1 2 29576 29579
0 29581 7 1 2 29574 29580
0 29582 5 1 1 29581
0 29583 7 1 2 52076 65711
0 29584 5 1 1 29583
0 29585 7 1 2 23878 29584
0 29586 5 1 1 29585
0 29587 7 1 2 44252 29586
0 29588 5 1 1 29587
0 29589 7 1 2 62376 65712
0 29590 5 1 1 29589
0 29591 7 1 2 29588 29590
0 29592 5 1 1 29591
0 29593 7 1 2 43353 29592
0 29594 5 2 1 29593
0 29595 7 2 2 52902 65713
0 29596 5 1 1 70324
0 29597 7 1 2 43130 68990
0 29598 5 1 1 29597
0 29599 7 1 2 29596 29598
0 29600 5 1 1 29599
0 29601 7 1 2 50096 29600
0 29602 5 1 1 29601
0 29603 7 1 2 70322 29602
0 29604 5 1 1 29603
0 29605 7 1 2 42874 29604
0 29606 5 1 1 29605
0 29607 7 1 2 46306 64215
0 29608 5 1 1 29607
0 29609 7 1 2 48653 58381
0 29610 5 1 1 29609
0 29611 7 1 2 29608 29610
0 29612 5 1 1 29611
0 29613 7 1 2 44093 29612
0 29614 5 1 1 29613
0 29615 7 1 2 52861 55386
0 29616 5 1 1 29615
0 29617 7 1 2 52713 58336
0 29618 5 2 1 29617
0 29619 7 1 2 29616 70326
0 29620 7 1 2 29614 29619
0 29621 5 1 1 29620
0 29622 7 1 2 65714 29621
0 29623 5 1 1 29622
0 29624 7 1 2 29606 29623
0 29625 5 1 1 29624
0 29626 7 1 2 47683 66229
0 29627 7 1 2 29625 29626
0 29628 5 1 1 29627
0 29629 7 1 2 29582 29628
0 29630 5 1 1 29629
0 29631 7 1 2 44483 29630
0 29632 5 1 1 29631
0 29633 7 1 2 29568 29632
0 29634 5 1 1 29633
0 29635 7 1 2 51311 29634
0 29636 5 1 1 29635
0 29637 7 1 2 29457 29636
0 29638 7 1 2 29274 29637
0 29639 5 1 1 29638
0 29640 7 1 2 51596 29639
0 29641 5 1 1 29640
0 29642 7 2 2 66141 67566
0 29643 5 1 1 70328
0 29644 7 1 2 18032 29643
0 29645 5 3 1 29644
0 29646 7 1 2 46081 70203
0 29647 5 1 1 29646
0 29648 7 1 2 61335 69440
0 29649 7 1 2 70206 29648
0 29650 5 1 1 29649
0 29651 7 1 2 29647 29650
0 29652 5 1 1 29651
0 29653 7 1 2 58166 29652
0 29654 5 1 1 29653
0 29655 7 1 2 64211 64864
0 29656 5 1 1 29655
0 29657 7 1 2 62967 29656
0 29658 5 1 1 29657
0 29659 7 1 2 46307 29658
0 29660 5 1 1 29659
0 29661 7 1 2 60194 6546
0 29662 5 1 1 29661
0 29663 7 1 2 65213 29662
0 29664 5 1 1 29663
0 29665 7 1 2 29660 29664
0 29666 5 1 1 29665
0 29667 7 1 2 65921 29666
0 29668 5 1 1 29667
0 29669 7 1 2 62965 68398
0 29670 5 1 1 29669
0 29671 7 1 2 29668 29670
0 29672 5 1 1 29671
0 29673 7 1 2 58209 29672
0 29674 5 1 1 29673
0 29675 7 1 2 29654 29674
0 29676 5 1 1 29675
0 29677 7 1 2 48142 29676
0 29678 5 1 1 29677
0 29679 7 4 2 61173 67940
0 29680 5 1 1 70333
0 29681 7 1 2 45616 57519
0 29682 5 1 1 29681
0 29683 7 1 2 21139 29682
0 29684 5 1 1 29683
0 29685 7 1 2 63592 29684
0 29686 5 1 1 29685
0 29687 7 1 2 52922 63485
0 29688 5 1 1 29687
0 29689 7 1 2 42875 58568
0 29690 5 1 1 29689
0 29691 7 1 2 29688 29690
0 29692 5 1 1 29691
0 29693 7 1 2 58167 29692
0 29694 5 1 1 29693
0 29695 7 1 2 29686 29694
0 29696 5 1 1 29695
0 29697 7 1 2 50010 29696
0 29698 5 1 1 29697
0 29699 7 1 2 42876 50123
0 29700 5 1 1 29699
0 29701 7 1 2 69905 29700
0 29702 5 1 1 29701
0 29703 7 1 2 48654 58168
0 29704 7 1 2 29702 29703
0 29705 5 1 1 29704
0 29706 7 1 2 29698 29705
0 29707 5 1 1 29706
0 29708 7 1 2 70334 29707
0 29709 5 1 1 29708
0 29710 7 1 2 29678 29709
0 29711 5 1 1 29710
0 29712 7 1 2 47684 29711
0 29713 5 1 1 29712
0 29714 7 1 2 46308 63715
0 29715 5 1 1 29714
0 29716 7 2 2 49302 58903
0 29717 7 1 2 50187 70337
0 29718 5 1 1 29717
0 29719 7 2 2 29715 29718
0 29720 5 2 1 70339
0 29721 7 1 2 9334 70340
0 29722 5 1 1 29721
0 29723 7 1 2 65715 29722
0 29724 5 1 1 29723
0 29725 7 1 2 50325 65922
0 29726 7 1 2 53796 29725
0 29727 5 1 1 29726
0 29728 7 1 2 29724 29727
0 29729 5 1 1 29728
0 29730 7 1 2 46082 29729
0 29731 5 1 1 29730
0 29732 7 1 2 70201 70341
0 29733 5 1 1 29732
0 29734 7 1 2 29731 29733
0 29735 5 1 1 29734
0 29736 7 1 2 45482 29735
0 29737 5 1 1 29736
0 29738 7 1 2 68750 70259
0 29739 5 1 1 29738
0 29740 7 1 2 61509 63293
0 29741 7 1 2 29739 29740
0 29742 5 1 1 29741
0 29743 7 1 2 29737 29742
0 29744 5 1 1 29743
0 29745 7 1 2 48143 29744
0 29746 5 1 1 29745
0 29747 7 1 2 42595 50097
0 29748 5 1 1 29747
0 29749 7 1 2 49013 53171
0 29750 5 1 1 29749
0 29751 7 1 2 29748 29750
0 29752 5 1 1 29751
0 29753 7 1 2 65923 29752
0 29754 5 1 1 29753
0 29755 7 1 2 68943 69844
0 29756 5 1 1 29755
0 29757 7 1 2 29754 29756
0 29758 5 1 1 29757
0 29759 7 1 2 44094 29758
0 29760 5 1 1 29759
0 29761 7 2 2 48031 64102
0 29762 7 1 2 52821 70343
0 29763 5 1 1 29762
0 29764 7 1 2 29760 29763
0 29765 5 1 1 29764
0 29766 7 1 2 43131 29765
0 29767 5 1 1 29766
0 29768 7 1 2 69967 70344
0 29769 5 1 1 29768
0 29770 7 1 2 29767 29769
0 29771 5 1 1 29770
0 29772 7 1 2 57200 29771
0 29773 5 1 1 29772
0 29774 7 1 2 29746 29773
0 29775 5 1 1 29774
0 29776 7 2 2 55960 59850
0 29777 7 1 2 29775 70345
0 29778 5 1 1 29777
0 29779 7 2 2 45483 61090
0 29780 7 1 2 61877 70018
0 29781 7 1 2 70347 29780
0 29782 5 1 1 29781
0 29783 7 1 2 45292 57944
0 29784 7 1 2 62556 29783
0 29785 7 1 2 63414 29784
0 29786 5 1 1 29785
0 29787 7 1 2 29782 29786
0 29788 5 1 1 29787
0 29789 7 1 2 57224 29788
0 29790 5 1 1 29789
0 29791 7 1 2 51182 1629
0 29792 5 1 1 29791
0 29793 7 2 2 50473 29792
0 29794 7 1 2 69454 70349
0 29795 5 1 1 29794
0 29796 7 1 2 64830 66006
0 29797 5 1 1 29796
0 29798 7 1 2 29795 29797
0 29799 5 1 1 29798
0 29800 7 1 2 57436 59851
0 29801 7 1 2 29799 29800
0 29802 5 1 1 29801
0 29803 7 1 2 29790 29802
0 29804 5 1 1 29803
0 29805 7 1 2 55961 29804
0 29806 5 1 1 29805
0 29807 7 1 2 54796 64103
0 29808 7 3 2 55666 60000
0 29809 7 1 2 62800 70351
0 29810 7 1 2 29807 29809
0 29811 7 1 2 70026 29810
0 29812 5 1 1 29811
0 29813 7 1 2 29806 29812
0 29814 5 1 1 29813
0 29815 7 1 2 55590 29814
0 29816 5 1 1 29815
0 29817 7 1 2 29778 29816
0 29818 7 1 2 29713 29817
0 29819 5 1 1 29818
0 29820 7 1 2 44484 29819
0 29821 5 1 1 29820
0 29822 7 1 2 62281 70199
0 29823 5 1 1 29822
0 29824 7 1 2 58923 59966
0 29825 5 1 1 29824
0 29826 7 1 2 29823 29825
0 29827 5 1 1 29826
0 29828 7 1 2 65924 29827
0 29829 5 1 1 29828
0 29830 7 1 2 55627 62277
0 29831 5 1 1 29830
0 29832 7 1 2 44485 59454
0 29833 5 1 1 29832
0 29834 7 1 2 29831 29833
0 29835 5 1 1 29834
0 29836 7 1 2 69704 29835
0 29837 5 1 1 29836
0 29838 7 1 2 29829 29837
0 29839 5 1 1 29838
0 29840 7 1 2 43354 29839
0 29841 5 1 1 29840
0 29842 7 2 2 42338 61736
0 29843 5 2 1 70354
0 29844 7 1 2 64027 66780
0 29845 5 1 1 29844
0 29846 7 1 2 70356 29845
0 29847 5 1 1 29846
0 29848 7 1 2 65434 70057
0 29849 7 1 2 29847 29848
0 29850 5 1 1 29849
0 29851 7 1 2 29841 29850
0 29852 5 1 1 29851
0 29853 7 1 2 47450 29852
0 29854 5 1 1 29853
0 29855 7 1 2 57974 65716
0 29856 5 1 1 29855
0 29857 7 1 2 66981 68489
0 29858 5 1 1 29857
0 29859 7 1 2 55916 63500
0 29860 7 1 2 29858 29859
0 29861 5 1 1 29860
0 29862 7 1 2 29856 29861
0 29863 5 1 1 29862
0 29864 7 1 2 45293 29863
0 29865 5 1 1 29864
0 29866 7 1 2 29854 29865
0 29867 5 1 1 29866
0 29868 7 1 2 63758 29867
0 29869 5 1 1 29868
0 29870 7 1 2 61326 66112
0 29871 5 1 1 29870
0 29872 7 2 2 49092 68476
0 29873 7 1 2 65832 70358
0 29874 5 1 1 29873
0 29875 7 1 2 29871 29874
0 29876 5 1 1 29875
0 29877 7 1 2 43355 29876
0 29878 5 1 1 29877
0 29879 7 1 2 62028 66972
0 29880 5 1 1 29879
0 29881 7 1 2 29878 29880
0 29882 5 1 1 29881
0 29883 7 1 2 49759 29882
0 29884 5 1 1 29883
0 29885 7 2 2 51211 61359
0 29886 7 1 2 63834 70360
0 29887 5 1 1 29886
0 29888 7 5 2 43356 65925
0 29889 7 1 2 60662 70362
0 29890 5 1 1 29889
0 29891 7 1 2 29887 29890
0 29892 5 1 1 29891
0 29893 7 1 2 50563 29892
0 29894 5 1 1 29893
0 29895 7 1 2 61920 63626
0 29896 5 1 1 29895
0 29897 7 1 2 68480 29896
0 29898 5 1 1 29897
0 29899 7 1 2 61360 63835
0 29900 7 1 2 57667 29899
0 29901 5 1 1 29900
0 29902 7 1 2 29898 29901
0 29903 5 1 1 29902
0 29904 7 1 2 46740 29903
0 29905 5 1 1 29904
0 29906 7 1 2 29894 29905
0 29907 7 1 2 29884 29906
0 29908 5 1 1 29907
0 29909 7 1 2 55962 29908
0 29910 5 1 1 29909
0 29911 7 1 2 29869 29910
0 29912 5 1 1 29911
0 29913 7 1 2 45617 29912
0 29914 5 1 1 29913
0 29915 7 4 2 55783 63753
0 29916 7 1 2 68329 69105
0 29917 5 1 1 29916
0 29918 7 1 2 43132 66352
0 29919 5 1 1 29918
0 29920 7 1 2 29917 29919
0 29921 5 1 1 29920
0 29922 7 1 2 45294 29921
0 29923 5 1 1 29922
0 29924 7 1 2 70323 29923
0 29925 5 1 1 29924
0 29926 7 1 2 70367 29925
0 29927 5 1 1 29926
0 29928 7 1 2 62225 63531
0 29929 5 1 1 29928
0 29930 7 1 2 49760 68418
0 29931 7 1 2 66964 29930
0 29932 7 1 2 29929 29931
0 29933 5 1 1 29932
0 29934 7 1 2 29927 29933
0 29935 5 1 1 29934
0 29936 7 1 2 46857 29935
0 29937 5 1 1 29936
0 29938 7 1 2 58708 65926
0 29939 5 1 1 29938
0 29940 7 1 2 56912 56929
0 29941 5 2 1 29940
0 29942 7 2 2 65717 70371
0 29943 5 1 1 70373
0 29944 7 1 2 29939 29943
0 29945 5 2 1 29944
0 29946 7 1 2 45295 70375
0 29947 5 1 1 29946
0 29948 7 1 2 64143 65927
0 29949 5 1 1 29948
0 29950 7 1 2 68504 29949
0 29951 5 1 1 29950
0 29952 7 1 2 56926 29951
0 29953 5 1 1 29952
0 29954 7 1 2 29947 29953
0 29955 5 1 1 29954
0 29956 7 1 2 59208 29955
0 29957 5 1 1 29956
0 29958 7 1 2 29937 29957
0 29959 5 1 1 29958
0 29960 7 1 2 42062 29959
0 29961 5 1 1 29960
0 29962 7 2 2 50788 51468
0 29963 5 1 1 70377
0 29964 7 1 2 6373 29963
0 29965 5 1 1 29964
0 29966 7 1 2 68443 29965
0 29967 5 1 1 29966
0 29968 7 1 2 62595 70325
0 29969 5 1 1 29968
0 29970 7 1 2 29967 29969
0 29971 5 2 1 29970
0 29972 7 1 2 66678 70379
0 29973 5 1 1 29972
0 29974 7 1 2 51506 67894
0 29975 5 1 1 29974
0 29976 7 1 2 66952 29975
0 29977 5 2 1 29976
0 29978 7 2 2 49124 57966
0 29979 7 1 2 67000 70383
0 29980 5 1 1 29979
0 29981 7 2 2 44686 63401
0 29982 7 1 2 65489 70385
0 29983 5 1 1 29982
0 29984 7 1 2 29980 29983
0 29985 5 1 1 29984
0 29986 7 1 2 70381 29985
0 29987 5 1 1 29986
0 29988 7 1 2 29973 29987
0 29989 7 1 2 29961 29988
0 29990 7 1 2 29914 29989
0 29991 5 1 1 29990
0 29992 7 1 2 42877 29991
0 29993 5 1 1 29992
0 29994 7 1 2 49228 62184
0 29995 5 2 1 29994
0 29996 7 1 2 43357 67275
0 29997 5 1 1 29996
0 29998 7 1 2 70387 29997
0 29999 5 1 1 29998
0 30000 7 1 2 63814 29999
0 30001 5 1 1 30000
0 30002 7 1 2 57597 59425
0 30003 5 1 1 30002
0 30004 7 1 2 52322 63815
0 30005 5 1 1 30004
0 30006 7 1 2 30003 30005
0 30007 5 1 1 30006
0 30008 7 1 2 43133 30007
0 30009 5 1 1 30008
0 30010 7 1 2 30001 30009
0 30011 5 1 1 30010
0 30012 7 1 2 65928 30011
0 30013 5 1 1 30012
0 30014 7 1 2 46309 50130
0 30015 5 2 1 30014
0 30016 7 1 2 58384 70389
0 30017 5 1 1 30016
0 30018 7 1 2 30017 70368
0 30019 5 1 1 30018
0 30020 7 2 2 46310 59240
0 30021 7 1 2 63555 70391
0 30022 5 1 1 30021
0 30023 7 1 2 30019 30022
0 30024 5 1 1 30023
0 30025 7 1 2 65718 30024
0 30026 5 1 1 30025
0 30027 7 1 2 30013 30026
0 30028 5 1 1 30027
0 30029 7 1 2 48655 30028
0 30030 5 1 1 30029
0 30031 7 2 2 47801 51569
0 30032 7 2 2 70013 70393
0 30033 5 1 1 70395
0 30034 7 1 2 48827 70396
0 30035 5 1 1 30034
0 30036 7 2 2 43134 70162
0 30037 7 1 2 68149 70397
0 30038 5 1 1 30037
0 30039 7 1 2 30035 30038
0 30040 5 1 1 30039
0 30041 7 1 2 57362 30040
0 30042 5 1 1 30041
0 30043 7 1 2 30030 30042
0 30044 5 1 1 30043
0 30045 7 1 2 44095 30044
0 30046 5 1 1 30045
0 30047 7 2 2 56353 57541
0 30048 7 2 2 63569 70399
0 30049 7 1 2 68419 70401
0 30050 5 1 1 30049
0 30051 7 1 2 60259 68399
0 30052 7 1 2 70398 30051
0 30053 5 1 1 30052
0 30054 7 1 2 30050 30053
0 30055 5 1 1 30054
0 30056 7 1 2 50011 30055
0 30057 5 1 1 30056
0 30058 7 1 2 30046 30057
0 30059 5 1 1 30058
0 30060 7 1 2 54797 30059
0 30061 5 1 1 30060
0 30062 7 1 2 50098 56932
0 30063 5 1 1 30062
0 30064 7 2 2 47579 57636
0 30065 7 1 2 68496 70403
0 30066 5 1 1 30065
0 30067 7 1 2 30063 30066
0 30068 5 2 1 30067
0 30069 7 1 2 44096 70405
0 30070 5 1 1 30069
0 30071 7 1 2 50099 56930
0 30072 5 1 1 30071
0 30073 7 2 2 51769 30072
0 30074 7 1 2 54236 70372
0 30075 7 1 2 70407 30074
0 30076 5 1 1 30075
0 30077 7 1 2 30070 30076
0 30078 5 1 1 30077
0 30079 7 1 2 59852 30078
0 30080 5 1 1 30079
0 30081 7 2 2 59881 66711
0 30082 7 1 2 55963 70409
0 30083 7 1 2 60843 30082
0 30084 5 1 1 30083
0 30085 7 1 2 30080 30084
0 30086 5 1 1 30085
0 30087 7 1 2 65719 30086
0 30088 5 1 1 30087
0 30089 7 1 2 58848 70392
0 30090 5 1 1 30089
0 30091 7 2 2 57637 58269
0 30092 5 1 1 70411
0 30093 7 1 2 61073 69937
0 30094 5 1 1 30093
0 30095 7 1 2 70412 30094
0 30096 5 1 1 30095
0 30097 7 1 2 30090 30096
0 30098 5 1 1 30097
0 30099 7 1 2 59853 30098
0 30100 5 1 1 30099
0 30101 7 1 2 59882 60508
0 30102 7 2 2 55679 56877
0 30103 7 1 2 67883 70413
0 30104 7 1 2 30101 30103
0 30105 5 1 1 30104
0 30106 7 1 2 30100 30105
0 30107 5 1 1 30106
0 30108 7 1 2 65929 30107
0 30109 5 1 1 30108
0 30110 7 1 2 30088 30109
0 30111 5 1 1 30110
0 30112 7 1 2 48656 30111
0 30113 5 1 1 30112
0 30114 7 2 2 47685 51212
0 30115 7 1 2 66712 70415
0 30116 5 1 1 30115
0 30117 7 1 2 28086 30116
0 30118 5 1 1 30117
0 30119 7 1 2 56904 30118
0 30120 5 1 1 30119
0 30121 7 1 2 57423 60935
0 30122 7 1 2 51530 30121
0 30123 5 1 1 30122
0 30124 7 1 2 30120 30123
0 30125 5 1 1 30124
0 30126 7 1 2 65720 30125
0 30127 5 1 1 30126
0 30128 7 4 2 42063 64028
0 30129 7 3 2 60646 70417
0 30130 7 2 2 48032 70421
0 30131 5 1 1 70424
0 30132 7 3 2 47580 57787
0 30133 7 1 2 53653 70426
0 30134 7 1 2 70425 30133
0 30135 5 1 1 30134
0 30136 7 1 2 30127 30135
0 30137 5 1 1 30136
0 30138 7 1 2 50618 30137
0 30139 5 1 1 30138
0 30140 7 1 2 70251 70410
0 30141 5 1 1 30140
0 30142 7 1 2 47581 63536
0 30143 5 1 1 30142
0 30144 7 1 2 53450 30143
0 30145 5 1 1 30144
0 30146 7 1 2 59854 30145
0 30147 5 1 1 30146
0 30148 7 1 2 30141 30147
0 30149 5 1 1 30148
0 30150 7 1 2 65930 30149
0 30151 5 1 1 30150
0 30152 7 2 2 49881 58283
0 30153 7 1 2 61758 70429
0 30154 5 1 1 30153
0 30155 7 1 2 51770 59811
0 30156 5 1 1 30155
0 30157 7 1 2 30154 30156
0 30158 5 1 1 30157
0 30159 7 1 2 65721 30158
0 30160 5 1 1 30159
0 30161 7 1 2 30151 30160
0 30162 5 1 1 30161
0 30163 7 1 2 56927 30162
0 30164 5 1 1 30163
0 30165 7 1 2 59812 69699
0 30166 5 1 1 30165
0 30167 7 2 2 58200 64117
0 30168 7 1 2 59883 62133
0 30169 7 1 2 70431 30168
0 30170 5 1 1 30169
0 30171 7 1 2 30166 30170
0 30172 5 1 1 30171
0 30173 7 1 2 56905 30172
0 30174 5 1 1 30173
0 30175 7 1 2 30164 30174
0 30176 7 1 2 30139 30175
0 30177 5 1 1 30176
0 30178 7 1 2 43135 30177
0 30179 5 1 1 30178
0 30180 7 1 2 30113 30179
0 30181 7 1 2 30061 30180
0 30182 7 1 2 29993 30181
0 30183 5 1 1 30182
0 30184 7 1 2 51312 30183
0 30185 5 1 1 30184
0 30186 7 2 2 48144 63607
0 30187 7 1 2 57919 63294
0 30188 7 1 2 60098 30187
0 30189 7 1 2 70433 30188
0 30190 5 1 1 30189
0 30191 7 2 2 58957 64371
0 30192 7 1 2 60107 64465
0 30193 7 1 2 70435 30192
0 30194 5 1 1 30193
0 30195 7 1 2 30190 30194
0 30196 5 1 1 30195
0 30197 7 1 2 55964 30196
0 30198 5 1 1 30197
0 30199 7 1 2 53859 64353
0 30200 7 1 2 68150 30199
0 30201 7 2 2 44097 64080
0 30202 7 2 2 55667 57614
0 30203 7 1 2 70437 70439
0 30204 7 1 2 30200 30203
0 30205 5 1 1 30204
0 30206 7 1 2 30198 30205
0 30207 5 1 1 30206
0 30208 7 1 2 45618 30207
0 30209 5 1 1 30208
0 30210 7 2 2 59980 64466
0 30211 7 1 2 70436 70441
0 30212 5 1 1 30211
0 30213 7 2 2 50422 63157
0 30214 5 1 1 70443
0 30215 7 1 2 57920 65833
0 30216 7 1 2 70444 30215
0 30217 7 1 2 63917 30216
0 30218 5 1 1 30217
0 30219 7 1 2 30212 30218
0 30220 5 1 1 30219
0 30221 7 1 2 55965 59371
0 30222 7 1 2 30220 30221
0 30223 5 1 1 30222
0 30224 7 1 2 30209 30223
0 30225 5 1 1 30224
0 30226 7 1 2 50866 30225
0 30227 5 1 1 30226
0 30228 7 4 2 51276 65722
0 30229 7 1 2 42878 69947
0 30230 5 1 1 30229
0 30231 7 1 2 59345 30230
0 30232 5 2 1 30231
0 30233 7 1 2 70445 70449
0 30234 5 1 1 30233
0 30235 7 2 2 51028 53283
0 30236 7 3 2 61416 67951
0 30237 7 1 2 48971 70453
0 30238 7 1 2 70451 30237
0 30239 5 1 1 30238
0 30240 7 1 2 30234 30239
0 30241 5 1 1 30240
0 30242 7 1 2 47582 30241
0 30243 5 1 1 30242
0 30244 7 3 2 51146 51645
0 30245 5 1 1 70456
0 30246 7 1 2 61112 70457
0 30247 5 1 1 30246
0 30248 7 1 2 51299 70069
0 30249 5 2 1 30248
0 30250 7 1 2 30247 70459
0 30251 5 1 1 30250
0 30252 7 1 2 65723 30251
0 30253 5 1 1 30252
0 30254 7 1 2 30243 30253
0 30255 5 1 1 30254
0 30256 7 1 2 54798 55966
0 30257 7 1 2 30255 30256
0 30258 5 1 1 30257
0 30259 7 1 2 58012 66484
0 30260 7 1 2 54687 30259
0 30261 7 1 2 67751 30260
0 30262 7 1 2 70452 30261
0 30263 5 1 1 30262
0 30264 7 1 2 30258 30263
0 30265 5 1 1 30264
0 30266 7 1 2 46741 30265
0 30267 5 1 1 30266
0 30268 7 2 2 63356 64874
0 30269 5 2 1 70461
0 30270 7 1 2 51277 70463
0 30271 5 1 1 30270
0 30272 7 1 2 49093 55994
0 30273 5 1 1 30272
0 30274 7 1 2 49622 61824
0 30275 5 1 1 30274
0 30276 7 1 2 30273 30275
0 30277 5 1 1 30276
0 30278 7 1 2 67889 30277
0 30279 5 1 1 30278
0 30280 7 1 2 30271 30279
0 30281 5 1 1 30280
0 30282 7 1 2 43358 30281
0 30283 5 1 1 30282
0 30284 7 1 2 30214 30245
0 30285 5 1 1 30284
0 30286 7 1 2 56722 30285
0 30287 5 1 1 30286
0 30288 7 1 2 30283 30287
0 30289 5 1 1 30288
0 30290 7 2 2 55967 65724
0 30291 7 1 2 54799 70465
0 30292 7 1 2 30289 30291
0 30293 5 1 1 30292
0 30294 7 1 2 30267 30293
0 30295 5 1 1 30294
0 30296 7 1 2 44352 30295
0 30297 5 1 1 30296
0 30298 7 1 2 52388 70446
0 30299 7 1 2 60819 30298
0 30300 5 1 1 30299
0 30301 7 1 2 53284 65186
0 30302 7 1 2 70192 30301
0 30303 5 1 1 30302
0 30304 7 1 2 30300 30303
0 30305 5 1 1 30304
0 30306 7 1 2 46311 30305
0 30307 5 1 1 30306
0 30308 7 1 2 48657 70447
0 30309 7 1 2 70215 30308
0 30310 5 1 1 30309
0 30311 7 1 2 30307 30310
0 30312 5 1 1 30311
0 30313 7 1 2 58201 63759
0 30314 7 1 2 30312 30313
0 30315 5 1 1 30314
0 30316 7 1 2 30297 30315
0 30317 5 1 1 30316
0 30318 7 1 2 47802 30317
0 30319 5 1 1 30318
0 30320 7 1 2 30227 30319
0 30321 7 1 2 30185 30320
0 30322 7 1 2 29821 30321
0 30323 5 1 1 30322
0 30324 7 1 2 70330 30323
0 30325 5 1 1 30324
0 30326 7 2 2 56243 66474
0 30327 7 1 2 63281 65845
0 30328 7 3 2 70467 30327
0 30329 7 1 2 49349 70469
0 30330 5 1 1 30329
0 30331 7 2 2 63608 64081
0 30332 7 1 2 61274 67749
0 30333 7 1 2 66216 30332
0 30334 7 1 2 70472 30333
0 30335 5 1 1 30334
0 30336 7 1 2 30330 30335
0 30337 5 1 1 30336
0 30338 7 1 2 51278 30337
0 30339 5 1 1 30338
0 30340 7 2 2 47686 67379
0 30341 7 2 2 45918 46083
0 30342 7 1 2 57615 70476
0 30343 7 1 2 64070 30342
0 30344 7 1 2 70474 30343
0 30345 7 1 2 70434 30344
0 30346 5 1 1 30345
0 30347 7 1 2 30339 30346
0 30348 5 1 1 30347
0 30349 7 1 2 65931 30348
0 30350 5 1 1 30349
0 30351 7 1 2 56246 57408
0 30352 7 1 2 69887 69396
0 30353 7 1 2 30351 30352
0 30354 5 1 1 30353
0 30355 7 1 2 30350 30354
0 30356 5 1 1 30355
0 30357 7 1 2 55591 30356
0 30358 5 1 1 30357
0 30359 7 1 2 51279 69049
0 30360 5 1 1 30359
0 30361 7 1 2 51300 57363
0 30362 5 1 1 30361
0 30363 7 1 2 30360 30362
0 30364 5 1 1 30363
0 30365 7 2 2 65725 30364
0 30366 7 1 2 61650 70478
0 30367 5 1 1 30366
0 30368 7 2 2 61084 63221
0 30369 7 1 2 57806 61878
0 30370 7 1 2 61297 30369
0 30371 7 1 2 70480 30370
0 30372 5 1 1 30371
0 30373 7 1 2 30367 30372
0 30374 5 1 1 30373
0 30375 7 1 2 66203 30374
0 30376 5 1 1 30375
0 30377 7 1 2 59021 61417
0 30378 7 1 2 61942 30377
0 30379 7 3 2 54083 63376
0 30380 7 1 2 66343 70482
0 30381 7 1 2 30378 30380
0 30382 5 1 1 30381
0 30383 7 1 2 61320 67138
0 30384 7 1 2 70479 30383
0 30385 5 1 1 30384
0 30386 7 1 2 30382 30385
0 30387 7 1 2 30376 30386
0 30388 5 1 1 30387
0 30389 7 1 2 48658 30388
0 30390 5 1 1 30389
0 30391 7 1 2 18208 69677
0 30392 5 1 1 30391
0 30393 7 1 2 60102 64467
0 30394 7 1 2 58958 30393
0 30395 7 1 2 30392 30394
0 30396 7 1 2 70272 30395
0 30397 5 1 1 30396
0 30398 7 1 2 30390 30397
0 30399 7 1 2 30358 30398
0 30400 5 1 1 30399
0 30401 7 1 2 57803 30400
0 30402 5 1 1 30401
0 30403 7 34 2 59209 70244
0 30404 7 1 2 64860 70485
0 30405 5 1 1 30404
0 30406 7 3 2 61596 70310
0 30407 7 1 2 63593 70519
0 30408 5 1 1 30407
0 30409 7 1 2 30405 30408
0 30410 5 1 1 30409
0 30411 7 1 2 50012 30410
0 30412 5 1 1 30411
0 30413 7 1 2 69975 70486
0 30414 5 1 1 30413
0 30415 7 1 2 30412 30414
0 30416 5 1 1 30415
0 30417 7 1 2 42596 30416
0 30418 5 1 1 30417
0 30419 7 1 2 43136 58066
0 30420 7 1 2 49014 30419
0 30421 7 2 2 66641 66070
0 30422 7 1 2 59560 70522
0 30423 7 1 2 30420 30422
0 30424 5 1 1 30423
0 30425 7 1 2 30418 30424
0 30426 5 1 1 30425
0 30427 7 1 2 57201 30426
0 30428 5 1 1 30427
0 30429 7 1 2 53285 70137
0 30430 7 2 2 66219 30429
0 30431 7 1 2 54978 70524
0 30432 5 1 1 30431
0 30433 7 1 2 50423 53797
0 30434 7 1 2 70487 30433
0 30435 5 1 1 30434
0 30436 7 1 2 30432 30435
0 30437 5 1 1 30436
0 30438 7 1 2 51234 30437
0 30439 5 1 1 30438
0 30440 7 2 2 49882 66142
0 30441 7 3 2 61259 66160
0 30442 7 1 2 48828 61097
0 30443 7 2 2 70528 30442
0 30444 7 1 2 70526 70531
0 30445 5 1 1 30444
0 30446 7 1 2 68666 69464
0 30447 5 2 1 30446
0 30448 7 3 2 55464 66161
0 30449 7 1 2 61743 66143
0 30450 7 1 2 70535 30449
0 30451 5 1 1 30450
0 30452 7 1 2 50789 30451
0 30453 5 1 1 30452
0 30454 7 2 2 59467 66071
0 30455 7 1 2 69482 70538
0 30456 5 1 1 30455
0 30457 7 3 2 64015 68187
0 30458 7 1 2 70536 70540
0 30459 5 1 1 30458
0 30460 7 1 2 50867 30459
0 30461 7 1 2 30456 30460
0 30462 5 1 1 30461
0 30463 7 1 2 30453 30462
0 30464 5 1 1 30463
0 30465 7 1 2 70533 30464
0 30466 5 1 1 30465
0 30467 7 1 2 43137 30466
0 30468 5 1 1 30467
0 30469 7 2 2 43604 67523
0 30470 7 2 2 69483 70543
0 30471 5 6 1 70545
0 30472 7 2 2 48829 57325
0 30473 7 1 2 59950 70553
0 30474 7 1 2 66220 30473
0 30475 5 1 1 30474
0 30476 7 1 2 70547 30475
0 30477 5 1 1 30476
0 30478 7 1 2 42879 30477
0 30479 5 1 1 30478
0 30480 7 1 2 45296 30479
0 30481 7 1 2 30468 30480
0 30482 5 1 1 30481
0 30483 7 1 2 46312 64931
0 30484 5 1 1 30483
0 30485 7 1 2 70217 30484
0 30486 5 1 1 30485
0 30487 7 1 2 70284 30486
0 30488 5 1 1 30487
0 30489 7 1 2 70086 70488
0 30490 5 1 1 30489
0 30491 7 1 2 48659 30490
0 30492 7 1 2 30488 30491
0 30493 5 1 1 30492
0 30494 7 1 2 30482 30493
0 30495 5 1 1 30494
0 30496 7 1 2 30445 30495
0 30497 5 1 1 30496
0 30498 7 1 2 50424 30497
0 30499 5 1 1 30498
0 30500 7 1 2 30439 30499
0 30501 5 1 1 30500
0 30502 7 1 2 48145 30501
0 30503 5 1 1 30502
0 30504 7 1 2 30428 30503
0 30505 5 1 1 30504
0 30506 7 1 2 65932 30505
0 30507 5 1 1 30506
0 30508 7 1 2 45484 52903
0 30509 7 1 2 70285 30508
0 30510 5 1 1 30509
0 30511 7 1 2 70548 30510
0 30512 5 1 1 30511
0 30513 7 1 2 42880 30512
0 30514 5 1 1 30513
0 30515 7 1 2 52099 70489
0 30516 5 1 1 30515
0 30517 7 1 2 30514 30516
0 30518 5 1 1 30517
0 30519 7 1 2 50100 30518
0 30520 5 1 1 30519
0 30521 7 2 2 65418 69982
0 30522 5 4 1 70555
0 30523 7 2 2 50868 70557
0 30524 7 1 2 70286 70561
0 30525 5 1 1 30524
0 30526 7 1 2 51469 55592
0 30527 7 1 2 70490 30526
0 30528 5 1 1 30527
0 30529 7 1 2 30525 30528
0 30530 5 1 1 30529
0 30531 7 1 2 48830 30530
0 30532 5 1 1 30531
0 30533 7 1 2 50013 70558
0 30534 5 1 1 30533
0 30535 7 1 2 68690 30534
0 30536 5 1 1 30535
0 30537 7 1 2 70287 30536
0 30538 5 1 1 30537
0 30539 7 1 2 67075 70520
0 30540 5 2 1 30539
0 30541 7 1 2 70534 70563
0 30542 5 1 1 30541
0 30543 7 1 2 52904 30542
0 30544 5 1 1 30543
0 30545 7 1 2 54907 65043
0 30546 5 1 1 30545
0 30547 7 1 2 70491 30546
0 30548 5 1 1 30547
0 30549 7 1 2 30544 30548
0 30550 7 1 2 30538 30549
0 30551 7 1 2 30532 30550
0 30552 7 1 2 30520 30551
0 30553 5 1 1 30552
0 30554 7 1 2 42597 30553
0 30555 5 1 1 30554
0 30556 7 2 2 48660 58376
0 30557 7 1 2 54249 70492
0 30558 7 1 2 70565 30557
0 30559 5 1 1 30558
0 30560 7 1 2 30555 30559
0 30561 5 1 1 30560
0 30562 7 1 2 43762 30561
0 30563 5 1 1 30562
0 30564 7 1 2 44353 49708
0 30565 7 1 2 57313 30564
0 30566 7 1 2 70255 30565
0 30567 5 1 1 30566
0 30568 7 1 2 44820 30567
0 30569 7 1 2 30563 30568
0 30570 5 1 1 30569
0 30571 7 1 2 51183 70342
0 30572 5 1 1 30571
0 30573 7 1 2 50014 62959
0 30574 5 2 1 30573
0 30575 7 1 2 30572 70567
0 30576 5 1 1 30575
0 30577 7 1 2 45485 30576
0 30578 5 1 1 30577
0 30579 7 2 2 69969 69971
0 30580 5 1 1 70569
0 30581 7 1 2 50015 63910
0 30582 5 1 1 30581
0 30583 7 2 2 63506 30582
0 30584 5 1 1 70571
0 30585 7 1 2 70570 70572
0 30586 5 1 1 30585
0 30587 7 1 2 50425 30586
0 30588 5 1 1 30587
0 30589 7 1 2 30578 30588
0 30590 5 1 1 30589
0 30591 7 1 2 70493 30590
0 30592 5 1 1 30591
0 30593 7 1 2 51235 70092
0 30594 5 1 1 30593
0 30595 7 1 2 58000 70562
0 30596 5 1 1 30595
0 30597 7 1 2 68691 30596
0 30598 5 1 1 30597
0 30599 7 1 2 50426 30598
0 30600 5 1 1 30599
0 30601 7 1 2 30594 30600
0 30602 5 1 1 30601
0 30603 7 1 2 70288 30602
0 30604 5 1 1 30603
0 30605 7 1 2 48146 30604
0 30606 7 1 2 30592 30605
0 30607 5 1 1 30606
0 30608 7 1 2 65726 30607
0 30609 7 1 2 30570 30608
0 30610 5 1 1 30609
0 30611 7 1 2 30507 30610
0 30612 5 1 1 30611
0 30613 7 1 2 62516 30612
0 30614 5 1 1 30613
0 30615 7 1 2 55995 65105
0 30616 5 1 1 30615
0 30617 7 1 2 49709 61825
0 30618 5 2 1 30617
0 30619 7 1 2 30616 70573
0 30620 5 1 1 30619
0 30621 7 4 2 61651 65727
0 30622 7 1 2 30620 70575
0 30623 5 1 1 30622
0 30624 7 1 2 51507 70213
0 30625 5 1 1 30624
0 30626 7 1 2 70052 30625
0 30627 5 1 1 30626
0 30628 7 1 2 42881 30627
0 30629 5 1 1 30628
0 30630 7 1 2 43359 59766
0 30631 5 1 1 30630
0 30632 7 1 2 62417 30631
0 30633 5 1 1 30632
0 30634 7 1 2 56221 30633
0 30635 5 1 1 30634
0 30636 7 1 2 57364 59340
0 30637 5 2 1 30636
0 30638 7 1 2 30635 70579
0 30639 7 1 2 30629 30638
0 30640 5 1 1 30639
0 30641 7 1 2 67844 30640
0 30642 5 1 1 30641
0 30643 7 1 2 30623 30642
0 30644 5 1 1 30643
0 30645 7 1 2 50427 30644
0 30646 5 1 1 30645
0 30647 7 2 2 56106 61652
0 30648 5 1 1 70581
0 30649 7 1 2 49303 62590
0 30650 5 1 1 30649
0 30651 7 1 2 30648 30650
0 30652 5 1 1 30651
0 30653 7 1 2 47583 30652
0 30654 5 1 1 30653
0 30655 7 1 2 61234 69026
0 30656 5 1 1 30655
0 30657 7 1 2 30654 30656
0 30658 5 1 1 30657
0 30659 7 1 2 65933 30658
0 30660 5 1 1 30659
0 30661 7 2 2 45619 63390
0 30662 7 1 2 58445 61361
0 30663 7 1 2 70583 30662
0 30664 5 1 1 30663
0 30665 7 1 2 30660 30664
0 30666 5 1 1 30665
0 30667 7 1 2 46742 30666
0 30668 5 1 1 30667
0 30669 7 3 2 59576 66689
0 30670 7 1 2 69415 70585
0 30671 5 1 1 30670
0 30672 7 1 2 30668 30671
0 30673 5 1 1 30672
0 30674 7 1 2 45297 61336
0 30675 7 1 2 30673 30674
0 30676 5 1 1 30675
0 30677 7 1 2 30646 30676
0 30678 5 1 1 30677
0 30679 7 1 2 48147 30678
0 30680 5 1 1 30679
0 30681 7 1 2 66007 70118
0 30682 5 1 1 30681
0 30683 7 1 2 49054 67066
0 30684 5 1 1 30683
0 30685 7 1 2 30682 30684
0 30686 5 1 1 30685
0 30687 7 1 2 48661 30686
0 30688 5 1 1 30687
0 30689 7 2 2 45620 63251
0 30690 7 1 2 70361 70588
0 30691 5 1 1 30690
0 30692 7 1 2 56354 68326
0 30693 5 1 1 30692
0 30694 7 1 2 30691 30693
0 30695 7 1 2 30688 30694
0 30696 5 1 1 30695
0 30697 7 1 2 46313 30696
0 30698 5 1 1 30697
0 30699 7 1 2 62185 68444
0 30700 5 1 1 30699
0 30701 7 2 2 60539 68400
0 30702 5 1 1 70590
0 30703 7 1 2 43360 70591
0 30704 5 1 1 30703
0 30705 7 1 2 30700 30704
0 30706 5 1 1 30705
0 30707 7 1 2 49229 30706
0 30708 5 1 1 30707
0 30709 7 1 2 57382 68445
0 30710 5 1 1 30709
0 30711 7 1 2 30702 30710
0 30712 5 1 1 30711
0 30713 7 1 2 43138 30712
0 30714 5 1 1 30713
0 30715 7 1 2 53366 64688
0 30716 7 1 2 70359 30715
0 30717 5 1 1 30716
0 30718 7 1 2 30714 30717
0 30719 7 1 2 30708 30718
0 30720 5 1 1 30719
0 30721 7 1 2 48662 30720
0 30722 5 1 1 30721
0 30723 7 1 2 30698 30722
0 30724 5 1 1 30723
0 30725 7 1 2 44098 30724
0 30726 5 1 1 30725
0 30727 7 1 2 59951 64529
0 30728 7 1 2 70584 30727
0 30729 5 1 1 30728
0 30730 7 1 2 30131 30729
0 30731 5 1 1 30730
0 30732 7 1 2 49761 30731
0 30733 5 1 1 30732
0 30734 7 2 2 55443 59162
0 30735 7 1 2 58793 63020
0 30736 7 1 2 70592 30735
0 30737 5 1 1 30736
0 30738 7 1 2 49230 30737
0 30739 7 1 2 30733 30738
0 30740 5 1 1 30739
0 30741 7 1 2 64229 65728
0 30742 5 1 1 30741
0 30743 7 1 2 70030 70422
0 30744 5 1 1 30743
0 30745 7 1 2 49182 30744
0 30746 7 1 2 30742 30745
0 30747 5 1 1 30746
0 30748 7 1 2 30740 30747
0 30749 5 1 1 30748
0 30750 7 1 2 59648 68446
0 30751 5 1 1 30750
0 30752 7 2 2 46743 63021
0 30753 7 1 2 59163 70594
0 30754 7 1 2 69924 30753
0 30755 5 1 1 30754
0 30756 7 1 2 30751 30755
0 30757 5 1 1 30756
0 30758 7 1 2 49094 30757
0 30759 5 1 1 30758
0 30760 7 1 2 63527 68447
0 30761 5 1 1 30760
0 30762 7 2 2 51476 66973
0 30763 5 1 1 70596
0 30764 7 1 2 63636 70597
0 30765 5 1 1 30764
0 30766 7 1 2 30761 30765
0 30767 7 1 2 30759 30766
0 30768 7 1 2 30749 30767
0 30769 5 1 1 30768
0 30770 7 1 2 42882 30769
0 30771 5 1 1 30770
0 30772 7 2 2 57921 63119
0 30773 7 1 2 59952 70598
0 30774 7 1 2 63594 30773
0 30775 5 1 1 30774
0 30776 7 1 2 60757 65338
0 30777 5 1 1 30776
0 30778 7 1 2 53729 70576
0 30779 7 1 2 30777 30778
0 30780 5 1 1 30779
0 30781 7 1 2 30775 30780
0 30782 5 1 1 30781
0 30783 7 1 2 44253 30782
0 30784 5 1 1 30783
0 30785 7 1 2 47584 64949
0 30786 5 2 1 30785
0 30787 7 1 2 46744 70600
0 30788 5 1 1 30787
0 30789 7 1 2 43361 63357
0 30790 7 1 2 64363 30789
0 30791 5 1 1 30790
0 30792 7 1 2 70577 30791
0 30793 7 1 2 30788 30792
0 30794 5 1 1 30793
0 30795 7 1 2 30784 30794
0 30796 5 1 1 30795
0 30797 7 1 2 51280 30796
0 30798 5 1 1 30797
0 30799 7 1 2 59666 62134
0 30800 7 2 2 64118 30799
0 30801 7 1 2 64181 70602
0 30802 5 1 1 30801
0 30803 7 1 2 64183 70603
0 30804 5 1 1 30803
0 30805 7 5 2 60647 64689
0 30806 7 1 2 44254 70604
0 30807 7 1 2 70400 30806
0 30808 5 1 1 30807
0 30809 7 1 2 30804 30808
0 30810 5 1 1 30809
0 30811 7 1 2 43362 30810
0 30812 5 1 1 30811
0 30813 7 1 2 30802 30812
0 30814 7 1 2 30798 30813
0 30815 7 1 2 30771 30814
0 30816 7 1 2 30726 30815
0 30817 5 1 1 30816
0 30818 7 1 2 51313 30817
0 30819 5 1 1 30818
0 30820 7 1 2 30680 30819
0 30821 5 1 1 30820
0 30822 7 1 2 66204 30821
0 30823 5 1 1 30822
0 30824 7 1 2 52408 65014
0 30825 5 1 1 30824
0 30826 7 1 2 52355 62600
0 30827 5 1 1 30826
0 30828 7 2 2 30825 30827
0 30829 5 2 1 70609
0 30830 7 1 2 46084 70611
0 30831 5 1 1 30830
0 30832 7 1 2 28707 30831
0 30833 5 1 1 30832
0 30834 7 1 2 48148 30833
0 30835 5 1 1 30834
0 30836 7 2 2 49231 51281
0 30837 5 1 1 70613
0 30838 7 1 2 57553 70614
0 30839 5 1 1 30838
0 30840 7 1 2 30835 30839
0 30841 5 1 1 30840
0 30842 7 1 2 46314 30841
0 30843 5 1 1 30842
0 30844 7 1 2 49055 51301
0 30845 5 1 1 30844
0 30846 7 1 2 30837 30845
0 30847 5 1 1 30846
0 30848 7 1 2 64456 30847
0 30849 5 1 1 30848
0 30850 7 1 2 30843 30849
0 30851 5 1 1 30850
0 30852 7 1 2 70289 30851
0 30853 5 1 1 30852
0 30854 7 1 2 59700 70601
0 30855 5 1 1 30854
0 30856 7 1 2 51282 30855
0 30857 5 1 1 30856
0 30858 7 1 2 70460 30857
0 30859 5 1 1 30858
0 30860 7 1 2 70494 30859
0 30861 5 1 1 30860
0 30862 7 1 2 30853 30861
0 30863 5 1 1 30862
0 30864 7 1 2 65729 30863
0 30865 5 1 1 30864
0 30866 7 2 2 51029 70495
0 30867 5 1 1 70615
0 30868 7 3 2 60025 66162
0 30869 7 1 2 70541 70617
0 30870 5 1 1 30869
0 30871 7 1 2 30867 30870
0 30872 5 1 1 30871
0 30873 7 1 2 68921 69745
0 30874 7 1 2 56171 30873
0 30875 7 1 2 30872 30874
0 30876 5 1 1 30875
0 30877 7 1 2 30865 30876
0 30878 5 1 1 30877
0 30879 7 1 2 46745 30878
0 30880 5 1 1 30879
0 30881 7 1 2 60170 70496
0 30882 5 1 1 30881
0 30883 7 1 2 57712 67130
0 30884 7 1 2 70529 30883
0 30885 5 1 1 30884
0 30886 7 1 2 30882 30885
0 30887 5 1 1 30886
0 30888 7 1 2 42883 30887
0 30889 5 1 1 30888
0 30890 7 1 2 48663 65304
0 30891 5 1 1 30890
0 30892 7 1 2 63522 30891
0 30893 5 1 1 30892
0 30894 7 1 2 70497 30893
0 30895 5 1 1 30894
0 30896 7 1 2 30889 30895
0 30897 5 1 1 30896
0 30898 7 1 2 65934 30897
0 30899 5 1 1 30898
0 30900 7 2 2 63737 66933
0 30901 7 4 2 69300 70620
0 30902 7 1 2 65305 70622
0 30903 5 1 1 30902
0 30904 7 1 2 20514 70388
0 30905 5 1 1 30904
0 30906 7 1 2 70498 30905
0 30907 5 1 1 30906
0 30908 7 1 2 65799 70499
0 30909 5 1 1 30908
0 30910 7 1 2 51355 61098
0 30911 7 1 2 66221 30910
0 30912 5 1 1 30911
0 30913 7 1 2 30909 30912
0 30914 5 1 1 30913
0 30915 7 1 2 45486 30914
0 30916 5 1 1 30915
0 30917 7 1 2 30907 30916
0 30918 5 1 1 30917
0 30919 7 1 2 65935 30918
0 30920 5 1 1 30919
0 30921 7 1 2 61247 63897
0 30922 7 1 2 69631 30921
0 30923 5 1 1 30922
0 30924 7 1 2 57355 70500
0 30925 5 1 1 30924
0 30926 7 1 2 30923 30925
0 30927 7 1 2 30920 30926
0 30928 5 1 1 30927
0 30929 7 1 2 48664 66008
0 30930 7 1 2 30928 30929
0 30931 5 1 1 30930
0 30932 7 1 2 30903 30931
0 30933 5 1 1 30932
0 30934 7 1 2 44099 30933
0 30935 5 1 1 30934
0 30936 7 1 2 30899 30935
0 30937 5 1 1 30936
0 30938 7 1 2 51314 30937
0 30939 5 1 1 30938
0 30940 7 1 2 54908 63358
0 30941 5 1 1 30940
0 30942 7 1 2 51283 30941
0 30943 5 1 1 30942
0 30944 7 1 2 49056 51294
0 30945 5 1 1 30944
0 30946 7 1 2 51315 55996
0 30947 7 1 2 30945 30946
0 30948 5 1 1 30947
0 30949 7 1 2 30943 30948
0 30950 5 1 1 30949
0 30951 7 1 2 70501 30950
0 30952 5 1 1 30951
0 30953 7 1 2 51107 62152
0 30954 5 1 1 30953
0 30955 7 1 2 51316 58361
0 30956 5 1 1 30955
0 30957 7 2 2 51147 61803
0 30958 5 2 1 70626
0 30959 7 1 2 30956 70628
0 30960 5 1 1 30959
0 30961 7 1 2 43139 30960
0 30962 5 1 1 30961
0 30963 7 1 2 30954 30962
0 30964 5 1 1 30963
0 30965 7 1 2 63609 70290
0 30966 7 1 2 30964 30965
0 30967 5 1 1 30966
0 30968 7 1 2 30952 30967
0 30969 5 1 1 30968
0 30970 7 1 2 43363 30969
0 30971 5 1 1 30970
0 30972 7 1 2 70304 70458
0 30973 5 1 1 30972
0 30974 7 1 2 49710 63158
0 30975 7 1 2 61717 30974
0 30976 5 1 1 30975
0 30977 7 1 2 30973 30976
0 30978 5 1 1 30977
0 30979 7 1 2 70502 30978
0 30980 5 1 1 30979
0 30981 7 1 2 30971 30980
0 30982 5 1 1 30981
0 30983 7 1 2 65730 30982
0 30984 5 1 1 30983
0 30985 7 1 2 30939 30984
0 30986 7 1 2 30880 30985
0 30987 5 1 1 30986
0 30988 7 1 2 60457 30987
0 30989 5 1 1 30988
0 30990 7 1 2 30823 30989
0 30991 7 1 2 30614 30990
0 30992 5 1 1 30991
0 30993 7 1 2 51667 30992
0 30994 5 1 1 30993
0 30995 7 1 2 30402 30994
0 30996 7 1 2 30325 30995
0 30997 7 1 2 29641 30996
0 30998 7 1 2 29135 30997
0 30999 5 1 1 30998
0 31000 7 1 2 54876 30999
0 31001 5 1 1 31000
0 31002 7 1 2 54940 70582
0 31003 5 1 1 31002
0 31004 7 2 2 47142 49350
0 31005 7 1 2 67817 70630
0 31006 5 1 1 31005
0 31007 7 1 2 31003 31006
0 31008 5 1 1 31007
0 31009 7 1 2 46085 31008
0 31010 5 1 1 31009
0 31011 7 1 2 58972 70231
0 31012 7 1 2 64225 31011
0 31013 5 1 1 31012
0 31014 7 1 2 31010 31013
0 31015 5 1 1 31014
0 31016 7 1 2 48287 31015
0 31017 5 1 1 31016
0 31018 7 2 2 45487 58824
0 31019 7 1 2 59395 62647
0 31020 7 1 2 70632 31019
0 31021 5 1 1 31020
0 31022 7 1 2 31017 31021
0 31023 5 1 1 31022
0 31024 7 1 2 66552 31023
0 31025 5 1 1 31024
0 31026 7 2 2 50365 51148
0 31027 7 1 2 47319 70605
0 31028 7 1 2 70634 31027
0 31029 7 1 2 70633 31028
0 31030 5 1 1 31029
0 31031 7 1 2 31025 31030
0 31032 5 1 1 31031
0 31033 7 1 2 46315 31032
0 31034 5 1 1 31033
0 31035 7 1 2 52759 55222
0 31036 7 1 2 63022 31035
0 31037 7 1 2 52242 59426
0 31038 7 1 2 65214 31037
0 31039 7 1 2 31036 31038
0 31040 5 1 1 31039
0 31041 7 1 2 31034 31040
0 31042 5 1 1 31041
0 31043 7 1 2 45120 31042
0 31044 5 1 1 31043
0 31045 7 1 2 47143 53002
0 31046 5 1 1 31045
0 31047 7 1 2 57693 31046
0 31048 5 1 1 31047
0 31049 7 1 2 46086 31048
0 31050 5 1 1 31049
0 31051 7 1 2 53201 62105
0 31052 5 1 1 31051
0 31053 7 1 2 31050 31052
0 31054 5 1 1 31053
0 31055 7 1 2 48831 59164
0 31056 7 1 2 66519 31055
0 31057 7 1 2 69143 31056
0 31058 7 1 2 31054 31057
0 31059 5 1 1 31058
0 31060 7 1 2 31044 31059
0 31061 5 1 1 31060
0 31062 7 1 2 45298 31061
0 31063 5 1 1 31062
0 31064 7 1 2 59165 62764
0 31065 7 1 2 55060 31064
0 31066 7 3 2 45621 64402
0 31067 7 2 2 52486 55490
0 31068 7 1 2 70636 70639
0 31069 7 1 2 31065 31068
0 31070 5 1 1 31069
0 31071 7 1 2 31063 31070
0 31072 5 1 1 31071
0 31073 7 1 2 53677 31072
0 31074 5 1 1 31073
0 31075 7 1 2 51082 55108
0 31076 5 1 1 31075
0 31077 7 1 2 52100 54851
0 31078 5 1 1 31077
0 31079 7 1 2 31076 31078
0 31080 5 2 1 31079
0 31081 7 1 2 48476 70641
0 31082 5 1 1 31081
0 31083 7 1 2 51483 55044
0 31084 5 1 1 31083
0 31085 7 1 2 31082 31084
0 31086 5 1 1 31085
0 31087 7 1 2 46087 31086
0 31088 5 1 1 31087
0 31089 7 1 2 55047 69549
0 31090 5 1 1 31089
0 31091 7 1 2 31088 31090
0 31092 5 2 1 31091
0 31093 7 1 2 44950 70643
0 31094 5 1 1 31093
0 31095 7 1 2 52441 65630
0 31096 5 1 1 31095
0 31097 7 2 2 48477 51070
0 31098 5 1 1 70645
0 31099 7 1 2 31096 31098
0 31100 5 1 1 31099
0 31101 7 2 2 53808 31100
0 31102 5 1 1 70647
0 31103 7 1 2 31094 31102
0 31104 5 1 1 31103
0 31105 7 1 2 68362 31104
0 31106 5 1 1 31105
0 31107 7 2 2 64403 64674
0 31108 7 1 2 55238 70171
0 31109 7 1 2 70649 31108
0 31110 5 1 1 31109
0 31111 7 1 2 31106 31110
0 31112 5 1 1 31111
0 31113 7 1 2 59537 31112
0 31114 5 1 1 31113
0 31115 7 1 2 49474 54059
0 31116 5 1 1 31115
0 31117 7 1 2 54738 31116
0 31118 5 1 1 31117
0 31119 7 1 2 54315 31118
0 31120 5 2 1 31119
0 31121 7 1 2 49809 59706
0 31122 5 1 1 31121
0 31123 7 1 2 22872 31122
0 31124 5 1 1 31123
0 31125 7 1 2 42884 31124
0 31126 5 1 1 31125
0 31127 7 1 2 49351 53784
0 31128 5 2 1 31127
0 31129 7 1 2 52487 61688
0 31130 5 1 1 31129
0 31131 7 1 2 70653 31130
0 31132 7 1 2 31126 31131
0 31133 5 1 1 31132
0 31134 7 1 2 43940 31133
0 31135 5 1 1 31134
0 31136 7 1 2 70651 31135
0 31137 5 1 1 31136
0 31138 7 1 2 45299 31137
0 31139 5 1 1 31138
0 31140 7 1 2 54831 56334
0 31141 5 1 1 31140
0 31142 7 1 2 31139 31141
0 31143 5 1 1 31142
0 31144 7 1 2 47144 31143
0 31145 5 1 1 31144
0 31146 7 1 2 52488 52852
0 31147 7 1 2 57689 31146
0 31148 5 1 1 31147
0 31149 7 1 2 31145 31148
0 31150 5 1 1 31149
0 31151 7 1 2 46088 31150
0 31152 5 1 1 31151
0 31153 7 1 2 57695 60089
0 31154 7 1 2 62101 31153
0 31155 5 1 1 31154
0 31156 7 1 2 31152 31155
0 31157 5 2 1 31156
0 31158 7 2 2 48033 63999
0 31159 7 1 2 67895 70657
0 31160 7 1 2 70655 31159
0 31161 5 1 1 31160
0 31162 7 1 2 31114 31161
0 31163 5 1 1 31162
0 31164 7 1 2 62517 31163
0 31165 5 1 1 31164
0 31166 7 3 2 53917 66553
0 31167 5 1 1 70659
0 31168 7 1 2 53901 66501
0 31169 5 1 1 31168
0 31170 7 1 2 31167 31169
0 31171 5 2 1 31170
0 31172 7 1 2 42598 70662
0 31173 5 1 1 31172
0 31174 7 1 2 54555 66520
0 31175 5 1 1 31174
0 31176 7 1 2 31173 31175
0 31177 5 1 1 31176
0 31178 7 2 2 47320 60648
0 31179 7 1 2 59127 61085
0 31180 7 1 2 70664 31179
0 31181 7 1 2 68757 31180
0 31182 7 1 2 31177 31181
0 31183 5 1 1 31182
0 31184 7 1 2 31165 31183
0 31185 7 1 2 31074 31184
0 31186 5 1 1 31185
0 31187 7 1 2 48149 31186
0 31188 5 1 1 31187
0 31189 7 1 2 56457 67465
0 31190 7 1 2 70109 31189
0 31191 7 1 2 64478 31190
0 31192 5 1 1 31191
0 31193 7 2 2 46858 61581
0 31194 5 1 1 70666
0 31195 7 1 2 55930 31194
0 31196 5 2 1 31195
0 31197 7 1 2 45622 70668
0 31198 5 1 1 31197
0 31199 7 1 2 4753 31198
0 31200 5 1 1 31199
0 31201 7 1 2 51062 66485
0 31202 7 1 2 67802 31201
0 31203 7 1 2 70138 31202
0 31204 7 1 2 31200 31203
0 31205 5 1 1 31204
0 31206 7 1 2 31192 31205
0 31207 5 1 1 31206
0 31208 7 1 2 46089 31207
0 31209 5 1 1 31208
0 31210 7 1 2 49466 54852
0 31211 5 1 1 31210
0 31212 7 1 2 45121 56265
0 31213 7 1 2 61542 31212
0 31214 5 1 1 31213
0 31215 7 1 2 31211 31214
0 31216 5 1 1 31215
0 31217 7 1 2 48665 31216
0 31218 5 1 1 31217
0 31219 7 1 2 61350 65015
0 31220 5 1 1 31219
0 31221 7 1 2 31218 31220
0 31222 5 1 1 31221
0 31223 7 2 2 58295 69199
0 31224 7 1 2 31222 70670
0 31225 5 1 1 31224
0 31226 7 1 2 31209 31225
0 31227 5 1 1 31226
0 31228 7 1 2 43941 31227
0 31229 5 1 1 31228
0 31230 7 1 2 42599 70642
0 31231 5 1 1 31230
0 31232 7 1 2 52101 55867
0 31233 5 1 1 31232
0 31234 7 1 2 31231 31233
0 31235 5 2 1 31234
0 31236 7 1 2 48478 70672
0 31237 5 1 1 31236
0 31238 7 1 2 69577 70350
0 31239 5 1 1 31238
0 31240 7 1 2 31237 31239
0 31241 5 1 1 31240
0 31242 7 1 2 70671 31241
0 31243 5 1 1 31242
0 31244 7 1 2 31229 31243
0 31245 5 1 1 31244
0 31246 7 1 2 48288 31245
0 31247 5 1 1 31246
0 31248 7 1 2 52102 55168
0 31249 5 1 1 31248
0 31250 7 1 2 47321 51184
0 31251 5 1 1 31250
0 31252 7 1 2 52067 53217
0 31253 5 1 1 31252
0 31254 7 1 2 31251 31253
0 31255 7 2 2 31249 31254
0 31256 7 1 2 65179 70674
0 31257 5 1 1 31256
0 31258 7 1 2 42600 70237
0 31259 7 1 2 69317 31258
0 31260 5 1 1 31259
0 31261 7 1 2 31257 31260
0 31262 5 1 1 31261
0 31263 7 1 2 56392 69200
0 31264 7 1 2 31262 31263
0 31265 5 1 1 31264
0 31266 7 1 2 31247 31265
0 31267 5 1 1 31266
0 31268 7 1 2 53612 31267
0 31269 5 1 1 31268
0 31270 7 4 2 44951 52103
0 31271 7 1 2 42885 70676
0 31272 5 2 1 31271
0 31273 7 1 2 51477 53809
0 31274 5 1 1 31273
0 31275 7 1 2 70680 31274
0 31276 5 2 1 31275
0 31277 7 1 2 48479 70682
0 31278 5 1 1 31277
0 31279 7 1 2 51983 70677
0 31280 5 1 1 31279
0 31281 7 1 2 31278 31280
0 31282 5 2 1 31281
0 31283 7 1 2 43763 70684
0 31284 5 1 1 31283
0 31285 7 1 2 54853 69321
0 31286 5 1 1 31285
0 31287 7 1 2 31284 31286
0 31288 5 1 1 31287
0 31289 7 1 2 42601 31288
0 31290 5 1 1 31289
0 31291 7 1 2 55868 69322
0 31292 5 1 1 31291
0 31293 7 1 2 31290 31292
0 31294 5 1 1 31293
0 31295 7 1 2 59234 70016
0 31296 7 1 2 31294 31295
0 31297 5 1 1 31296
0 31298 7 1 2 31269 31297
0 31299 7 1 2 31188 31298
0 31300 5 1 1 31299
0 31301 7 1 2 66278 31300
0 31302 5 1 1 31301
0 31303 7 1 2 68401 68547
0 31304 5 1 1 31303
0 31305 7 4 2 45122 65936
0 31306 7 1 2 57401 70686
0 31307 5 1 1 31306
0 31308 7 1 2 31304 31307
0 31309 5 1 1 31308
0 31310 7 1 2 61054 31309
0 31311 5 1 1 31310
0 31312 7 3 2 46316 63802
0 31313 7 1 2 61798 67833
0 31314 7 1 2 70690 31313
0 31315 5 1 1 31314
0 31316 7 1 2 31311 31315
0 31317 5 1 1 31316
0 31318 7 1 2 53286 31317
0 31319 5 1 1 31318
0 31320 7 3 2 51861 66690
0 31321 5 1 1 70693
0 31322 7 2 2 48943 61582
0 31323 7 1 2 63803 70696
0 31324 5 1 1 31323
0 31325 7 1 2 31321 31324
0 31326 5 1 1 31325
0 31327 7 1 2 44952 55115
0 31328 7 1 2 31326 31327
0 31329 5 1 1 31328
0 31330 7 1 2 31319 31329
0 31331 5 1 1 31330
0 31332 7 1 2 48150 31331
0 31333 5 1 1 31332
0 31334 7 1 2 53864 54525
0 31335 7 1 2 70694 31334
0 31336 5 1 1 31335
0 31337 7 1 2 31333 31336
0 31338 5 1 1 31337
0 31339 7 1 2 43478 31338
0 31340 5 1 1 31339
0 31341 7 2 2 67149 69902
0 31342 7 1 2 59981 65544
0 31343 7 1 2 56376 31342
0 31344 7 1 2 70698 31343
0 31345 5 1 1 31344
0 31346 7 1 2 31340 31345
0 31347 5 1 1 31346
0 31348 7 1 2 42064 31347
0 31349 5 1 1 31348
0 31350 7 1 2 61029 68456
0 31351 7 1 2 61848 31350
0 31352 7 1 2 70699 31351
0 31353 5 1 1 31352
0 31354 7 1 2 31349 31353
0 31355 5 1 1 31354
0 31356 7 1 2 52077 31355
0 31357 5 1 1 31356
0 31358 7 1 2 54189 66009
0 31359 5 1 1 31358
0 31360 7 1 2 49352 60269
0 31361 5 1 1 31360
0 31362 7 2 2 53331 13618
0 31363 5 1 1 70700
0 31364 7 1 2 50474 70701
0 31365 7 1 2 31361 31364
0 31366 5 1 1 31365
0 31367 7 1 2 9780 31366
0 31368 5 1 1 31367
0 31369 7 1 2 49426 65937
0 31370 7 1 2 31368 31369
0 31371 5 1 1 31370
0 31372 7 1 2 31359 31371
0 31373 5 1 1 31372
0 31374 7 1 2 48666 31373
0 31375 5 2 1 31374
0 31376 7 1 2 54185 61866
0 31377 5 2 1 31376
0 31378 7 1 2 43764 69530
0 31379 5 1 1 31378
0 31380 7 1 2 70704 31379
0 31381 5 1 1 31380
0 31382 7 1 2 66010 31381
0 31383 5 1 1 31382
0 31384 7 1 2 70702 31383
0 31385 5 1 1 31384
0 31386 7 1 2 48289 31385
0 31387 5 1 1 31386
0 31388 7 2 2 52104 66011
0 31389 7 2 2 44953 54186
0 31390 7 1 2 51149 70708
0 31391 7 1 2 70706 31390
0 31392 5 2 1 31391
0 31393 7 1 2 44821 70710
0 31394 7 1 2 31387 31393
0 31395 5 1 1 31394
0 31396 7 2 2 52645 70678
0 31397 7 1 2 65215 70712
0 31398 5 1 1 31397
0 31399 7 1 2 53287 68548
0 31400 5 1 1 31399
0 31401 7 1 2 53902 55023
0 31402 5 1 1 31401
0 31403 7 1 2 52438 31402
0 31404 7 1 2 31400 31403
0 31405 5 1 1 31404
0 31406 7 1 2 61612 31405
0 31407 5 1 1 31406
0 31408 7 1 2 31398 31407
0 31409 5 1 1 31408
0 31410 7 1 2 65731 31409
0 31411 5 1 1 31410
0 31412 7 1 2 54136 68765
0 31413 5 1 1 31412
0 31414 7 1 2 54037 54176
0 31415 5 1 1 31414
0 31416 7 1 2 31413 31415
0 31417 5 1 1 31416
0 31418 7 1 2 52455 65938
0 31419 7 1 2 31417 31418
0 31420 5 1 1 31419
0 31421 7 1 2 48151 31420
0 31422 7 1 2 31411 31421
0 31423 5 1 1 31422
0 31424 7 1 2 61240 31423
0 31425 7 1 2 31395 31424
0 31426 5 1 1 31425
0 31427 7 1 2 31357 31426
0 31428 5 1 1 31427
0 31429 7 1 2 44354 31428
0 31430 5 1 1 31429
0 31431 7 1 2 65939 70656
0 31432 5 1 1 31431
0 31433 7 2 2 49821 54702
0 31434 7 1 2 56087 70714
0 31435 7 1 2 70650 31434
0 31436 5 1 1 31435
0 31437 7 1 2 31432 31436
0 31438 5 1 1 31437
0 31439 7 1 2 58160 31438
0 31440 5 1 1 31439
0 31441 7 2 2 54192 63023
0 31442 7 3 2 60246 69430
0 31443 7 1 2 58028 70718
0 31444 7 1 2 70716 31443
0 31445 5 1 1 31444
0 31446 7 1 2 31440 31445
0 31447 5 1 1 31446
0 31448 7 1 2 60040 61597
0 31449 7 1 2 31447 31448
0 31450 5 1 1 31449
0 31451 7 1 2 31430 31450
0 31452 5 1 1 31451
0 31453 7 1 2 67021 31452
0 31454 5 1 1 31453
0 31455 7 1 2 52287 60103
0 31456 7 1 2 67093 31455
0 31457 5 1 1 31456
0 31458 7 1 2 51271 65860
0 31459 7 1 2 59751 31458
0 31460 7 1 2 63314 31459
0 31461 5 1 1 31460
0 31462 7 1 2 31457 31461
0 31463 5 1 1 31462
0 31464 7 1 2 68402 31463
0 31465 5 1 1 31464
0 31466 7 1 2 54854 70477
0 31467 7 2 2 67144 31466
0 31468 7 1 2 45860 49661
0 31469 7 1 2 68209 31468
0 31470 7 1 2 70721 31469
0 31471 5 1 1 31470
0 31472 7 1 2 31465 31471
0 31473 5 1 1 31472
0 31474 7 1 2 43942 31473
0 31475 5 1 1 31474
0 31476 7 2 2 63768 66906
0 31477 7 2 2 63666 66144
0 31478 7 1 2 68118 70725
0 31479 7 1 2 70723 31478
0 31480 7 1 2 54129 31479
0 31481 5 1 1 31480
0 31482 7 1 2 31475 31481
0 31483 5 1 1 31482
0 31484 7 1 2 45300 31483
0 31485 5 1 1 31484
0 31486 7 1 2 45861 68973
0 31487 7 1 2 69235 31486
0 31488 7 1 2 70269 31487
0 31489 5 1 1 31488
0 31490 7 1 2 31485 31489
0 31491 5 1 1 31490
0 31492 7 1 2 42065 31491
0 31493 5 1 1 31492
0 31494 7 1 2 54941 68725
0 31495 5 1 1 31494
0 31496 7 1 2 53057 54858
0 31497 5 1 1 31496
0 31498 7 1 2 31495 31497
0 31499 5 1 1 31498
0 31500 7 1 2 65940 31499
0 31501 5 1 1 31500
0 31502 7 1 2 42339 54100
0 31503 7 1 2 67259 31502
0 31504 5 1 1 31503
0 31505 7 1 2 31501 31504
0 31506 5 1 1 31505
0 31507 7 1 2 46090 31506
0 31508 5 1 1 31507
0 31509 7 1 2 52489 56355
0 31510 7 1 2 56825 64104
0 31511 7 1 2 31509 31510
0 31512 5 1 1 31511
0 31513 7 1 2 31508 31512
0 31514 5 1 1 31513
0 31515 7 1 2 63098 67048
0 31516 7 1 2 31514 31515
0 31517 5 1 1 31516
0 31518 7 1 2 31493 31517
0 31519 5 1 1 31518
0 31520 7 1 2 47451 31519
0 31521 5 1 1 31520
0 31522 7 2 2 45623 67049
0 31523 5 1 1 70727
0 31524 7 1 2 66398 67421
0 31525 5 1 1 31524
0 31526 7 1 2 31523 31525
0 31527 5 8 1 31526
0 31528 7 1 2 49794 53127
0 31529 7 1 2 68210 31528
0 31530 7 1 2 70186 31529
0 31531 7 1 2 70729 31530
0 31532 5 1 1 31531
0 31533 7 1 2 31521 31532
0 31534 5 1 1 31533
0 31535 7 1 2 46534 31534
0 31536 5 1 1 31535
0 31537 7 1 2 53427 68726
0 31538 5 1 1 31537
0 31539 7 1 2 70654 31538
0 31540 5 1 1 31539
0 31541 7 1 2 43943 31540
0 31542 5 1 1 31541
0 31543 7 1 2 70652 31542
0 31544 5 1 1 31543
0 31545 7 1 2 59752 68991
0 31546 7 1 2 70730 31545
0 31547 7 1 2 31544 31546
0 31548 5 1 1 31547
0 31549 7 1 2 31536 31548
0 31550 5 1 1 31549
0 31551 7 1 2 59301 31550
0 31552 5 1 1 31551
0 31553 7 2 2 68101 68712
0 31554 7 1 2 65732 70644
0 31555 5 1 1 31554
0 31556 7 1 2 70687 70675
0 31557 5 1 1 31556
0 31558 7 1 2 31555 31557
0 31559 5 1 1 31558
0 31560 7 1 2 44954 31559
0 31561 5 1 1 31560
0 31562 7 1 2 65733 70648
0 31563 5 1 1 31562
0 31564 7 1 2 31561 31563
0 31565 5 1 1 31564
0 31566 7 1 2 70737 31565
0 31567 5 1 1 31566
0 31568 7 1 2 48152 31567
0 31569 7 1 2 31552 31568
0 31570 5 1 1 31569
0 31571 7 1 2 50722 69550
0 31572 5 1 1 31571
0 31573 7 1 2 31572 70705
0 31574 5 1 1 31573
0 31575 7 1 2 66012 31574
0 31576 5 1 1 31575
0 31577 7 1 2 70703 31576
0 31578 5 1 1 31577
0 31579 7 1 2 48290 31578
0 31580 5 1 1 31579
0 31581 7 1 2 31580 70711
0 31582 5 1 1 31581
0 31583 7 1 2 70738 31582
0 31584 5 1 1 31583
0 31585 7 1 2 44822 31584
0 31586 5 1 1 31585
0 31587 7 1 2 44486 31586
0 31588 7 1 2 31570 31587
0 31589 5 1 1 31588
0 31590 7 1 2 52596 59682
0 31591 7 1 2 64664 31590
0 31592 7 1 2 69337 31591
0 31593 5 1 1 31592
0 31594 7 1 2 59577 67287
0 31595 7 1 2 54706 31594
0 31596 7 1 2 63315 68250
0 31597 7 1 2 31595 31596
0 31598 5 1 1 31597
0 31599 7 1 2 31593 31598
0 31600 5 1 1 31599
0 31601 7 1 2 45301 63135
0 31602 7 1 2 31600 31601
0 31603 5 1 1 31602
0 31604 7 1 2 55514 64580
0 31605 7 2 2 48832 55491
0 31606 7 1 2 66344 69697
0 31607 7 1 2 70739 31606
0 31608 7 1 2 31604 31607
0 31609 5 1 1 31608
0 31610 7 1 2 31603 31609
0 31611 5 1 1 31610
0 31612 7 1 2 46091 31611
0 31613 5 1 1 31612
0 31614 7 6 2 59302 65941
0 31615 5 4 1 70741
0 31616 7 1 2 53202 64093
0 31617 7 1 2 65049 31616
0 31618 7 1 2 70742 31617
0 31619 7 1 2 69338 31618
0 31620 5 1 1 31619
0 31621 7 1 2 31613 31620
0 31622 5 1 1 31621
0 31623 7 1 2 48291 31622
0 31624 5 1 1 31623
0 31625 7 3 2 42340 50366
0 31626 7 1 2 45766 70751
0 31627 5 1 1 31626
0 31628 7 1 2 70747 31627
0 31629 5 3 1 31628
0 31630 7 1 2 51150 64094
0 31631 7 1 2 69391 31630
0 31632 7 1 2 70754 31631
0 31633 7 1 2 69339 31632
0 31634 5 1 1 31633
0 31635 7 1 2 31624 31634
0 31636 5 1 1 31635
0 31637 7 1 2 46535 31636
0 31638 5 1 1 31637
0 31639 7 1 2 43765 64000
0 31640 7 1 2 68127 31639
0 31641 5 2 1 31640
0 31642 7 1 2 53918 70743
0 31643 5 1 1 31642
0 31644 7 1 2 70757 31643
0 31645 5 1 1 31644
0 31646 7 1 2 42602 31645
0 31647 5 1 1 31646
0 31648 7 2 2 42227 63295
0 31649 7 1 2 52534 58739
0 31650 7 1 2 70759 31649
0 31651 5 1 1 31650
0 31652 7 1 2 31647 31651
0 31653 5 1 1 31652
0 31654 7 1 2 44355 65385
0 31655 7 1 2 69340 31654
0 31656 7 1 2 31653 31655
0 31657 5 1 1 31656
0 31658 7 1 2 31638 31657
0 31659 5 1 1 31658
0 31660 7 1 2 47803 68644
0 31661 7 1 2 31659 31660
0 31662 5 1 1 31661
0 31663 7 1 2 31589 31662
0 31664 7 1 2 31454 31663
0 31665 7 1 2 31302 31664
0 31666 5 1 1 31665
0 31667 7 1 2 50101 31666
0 31668 5 1 1 31667
0 31669 7 2 2 50141 52511
0 31670 7 2 2 46092 60001
0 31671 7 1 2 49861 70763
0 31672 7 1 2 70731 31671
0 31673 5 1 1 31672
0 31674 7 1 2 45123 55814
0 31675 7 1 2 67466 31674
0 31676 7 1 2 67022 31675
0 31677 5 1 1 31676
0 31678 7 1 2 31673 31677
0 31679 5 1 1 31678
0 31680 7 1 2 70761 31679
0 31681 5 1 1 31680
0 31682 7 3 2 42066 42603
0 31683 7 2 2 64354 70765
0 31684 7 1 2 51843 60191
0 31685 7 1 2 70768 31684
0 31686 7 1 2 67023 31685
0 31687 5 1 1 31686
0 31688 7 1 2 31681 31687
0 31689 5 1 1 31688
0 31690 7 1 2 43944 31689
0 31691 5 1 1 31690
0 31692 7 1 2 53533 65122
0 31693 5 1 1 31692
0 31694 7 1 2 58296 60108
0 31695 7 1 2 68622 31694
0 31696 7 1 2 31693 31695
0 31697 7 1 2 67024 31696
0 31698 5 1 1 31697
0 31699 7 1 2 31691 31698
0 31700 5 1 1 31699
0 31701 7 1 2 65942 31700
0 31702 5 1 1 31701
0 31703 7 2 2 52646 65453
0 31704 5 1 1 70770
0 31705 7 1 2 61788 63402
0 31706 7 1 2 68345 31705
0 31707 7 1 2 70771 31706
0 31708 7 1 2 67025 31707
0 31709 5 1 1 31708
0 31710 7 1 2 31702 31709
0 31711 5 1 1 31710
0 31712 7 1 2 48833 31711
0 31713 5 1 1 31712
0 31714 7 1 2 53178 66735
0 31715 7 1 2 66930 68581
0 31716 7 2 2 46317 54006
0 31717 7 1 2 68599 70772
0 31718 7 1 2 31715 31717
0 31719 7 1 2 31714 31718
0 31720 5 1 1 31719
0 31721 7 1 2 31713 31720
0 31722 5 1 1 31721
0 31723 7 1 2 44955 31722
0 31724 5 1 1 31723
0 31725 7 1 2 48944 64095
0 31726 7 1 2 64690 31725
0 31727 7 1 2 59670 67100
0 31728 7 1 2 70267 31727
0 31729 7 1 2 31726 31728
0 31730 5 1 1 31729
0 31731 7 1 2 31724 31730
0 31732 5 1 1 31731
0 31733 7 1 2 44487 31732
0 31734 5 1 1 31733
0 31735 7 2 2 47914 67026
0 31736 7 2 2 48153 67946
0 31737 5 1 1 70776
0 31738 7 1 2 54800 61583
0 31739 7 1 2 70777 31738
0 31740 5 1 1 31739
0 31741 7 6 2 57922 64691
0 31742 7 1 2 50698 55864
0 31743 7 1 2 56266 31742
0 31744 7 1 2 70778 31743
0 31745 5 1 1 31744
0 31746 7 1 2 31740 31745
0 31747 5 1 1 31746
0 31748 7 1 2 42886 31747
0 31749 5 1 1 31748
0 31750 7 1 2 51284 66013
0 31751 5 1 1 31750
0 31752 7 1 2 65181 65943
0 31753 5 1 1 31752
0 31754 7 1 2 31751 31753
0 31755 5 1 1 31754
0 31756 7 1 2 43479 56196
0 31757 7 1 2 31755 31756
0 31758 5 1 1 31757
0 31759 7 1 2 31749 31758
0 31760 5 1 1 31759
0 31761 7 1 2 43945 31760
0 31762 5 1 1 31761
0 31763 7 3 2 48834 66014
0 31764 7 3 2 56537 63469
0 31765 7 1 2 44823 51844
0 31766 7 1 2 55865 31765
0 31767 7 1 2 70787 31766
0 31768 7 1 2 70784 31767
0 31769 5 1 1 31768
0 31770 7 1 2 31762 31769
0 31771 5 1 1 31770
0 31772 7 1 2 48667 31771
0 31773 5 1 1 31772
0 31774 7 1 2 52647 66015
0 31775 7 1 2 70238 31774
0 31776 5 1 1 31775
0 31777 7 1 2 49569 52983
0 31778 7 1 2 70454 31777
0 31779 5 1 1 31778
0 31780 7 1 2 31776 31779
0 31781 5 1 1 31780
0 31782 7 1 2 42604 31781
0 31783 5 1 1 31782
0 31784 7 1 2 52270 54993
0 31785 7 1 2 70688 31784
0 31786 5 1 1 31785
0 31787 7 1 2 31783 31786
0 31788 5 1 1 31787
0 31789 7 1 2 48912 56189
0 31790 7 1 2 31788 31789
0 31791 5 1 1 31790
0 31792 7 1 2 31773 31791
0 31793 5 1 1 31792
0 31794 7 1 2 44956 31793
0 31795 5 1 1 31794
0 31796 7 1 2 49570 65517
0 31797 5 1 1 31796
0 31798 7 1 2 56222 69749
0 31799 5 1 1 31798
0 31800 7 1 2 31797 31799
0 31801 5 1 1 31800
0 31802 7 2 2 50475 31801
0 31803 7 1 2 57735 62801
0 31804 7 1 2 67631 31803
0 31805 7 1 2 70790 31804
0 31806 5 1 1 31805
0 31807 7 1 2 31795 31806
0 31808 5 1 1 31807
0 31809 7 1 2 70774 31808
0 31810 5 1 1 31809
0 31811 7 3 2 48034 63296
0 31812 7 1 2 54880 70792
0 31813 5 1 1 31812
0 31814 7 1 2 49571 65734
0 31815 7 1 2 58976 31814
0 31816 5 1 1 31815
0 31817 7 1 2 31813 31816
0 31818 5 1 1 31817
0 31819 7 4 2 59695 66195
0 31820 7 5 2 44595 44957
0 31821 7 1 2 57807 70799
0 31822 7 1 2 70795 31821
0 31823 7 1 2 31818 31822
0 31824 5 1 1 31823
0 31825 7 1 2 31810 31824
0 31826 5 1 1 31825
0 31827 7 1 2 44356 31826
0 31828 5 1 1 31827
0 31829 7 1 2 57225 67772
0 31830 7 1 2 58522 31829
0 31831 7 1 2 65050 67041
0 31832 7 1 2 68531 31831
0 31833 7 1 2 31830 31832
0 31834 5 1 1 31833
0 31835 7 1 2 55223 65318
0 31836 5 1 1 31835
0 31837 7 1 2 50664 67724
0 31838 5 1 1 31837
0 31839 7 1 2 31836 31838
0 31840 5 1 1 31839
0 31841 7 1 2 64487 31840
0 31842 5 1 1 31841
0 31843 7 2 2 57202 60090
0 31844 5 1 1 70804
0 31845 7 1 2 65735 70805
0 31846 5 1 1 31845
0 31847 7 1 2 29680 31737
0 31848 5 1 1 31847
0 31849 7 1 2 52648 31848
0 31850 5 1 1 31849
0 31851 7 1 2 31846 31850
0 31852 5 1 1 31851
0 31853 7 1 2 54832 31852
0 31854 5 1 1 31853
0 31855 7 1 2 31842 31854
0 31856 5 1 1 31855
0 31857 7 1 2 51404 31856
0 31858 5 1 1 31857
0 31859 7 1 2 50665 64488
0 31860 7 1 2 58658 31859
0 31861 5 1 1 31860
0 31862 7 1 2 31858 31861
0 31863 5 1 1 31862
0 31864 7 1 2 56190 70732
0 31865 7 1 2 31863 31864
0 31866 5 1 1 31865
0 31867 7 1 2 31834 31866
0 31868 5 1 1 31867
0 31869 7 1 2 60002 31868
0 31870 5 1 1 31869
0 31871 7 1 2 31828 31870
0 31872 5 1 1 31871
0 31873 7 1 2 44100 31872
0 31874 5 1 1 31873
0 31875 7 3 2 51083 51272
0 31876 7 1 2 44824 53865
0 31877 7 1 2 70806 31876
0 31878 5 2 1 31877
0 31879 7 1 2 49795 63216
0 31880 7 1 2 62171 31879
0 31881 5 1 1 31880
0 31882 7 1 2 70809 31881
0 31883 5 1 1 31882
0 31884 7 1 2 60694 65736
0 31885 7 1 2 31883 31884
0 31886 5 1 1 31885
0 31887 7 2 2 46318 53971
0 31888 5 1 1 70811
0 31889 7 1 2 51030 55527
0 31890 5 1 1 31889
0 31891 7 1 2 31888 31890
0 31892 5 2 1 31891
0 31893 7 3 2 56628 70813
0 31894 5 1 1 70815
0 31895 7 2 2 45862 51151
0 31896 7 1 2 59790 62215
0 31897 7 1 2 70818 31896
0 31898 7 1 2 70816 31897
0 31899 5 1 1 31898
0 31900 7 1 2 31886 31899
0 31901 5 1 1 31900
0 31902 7 1 2 70775 31901
0 31903 5 1 1 31902
0 31904 7 2 2 44596 48480
0 31905 7 2 2 51317 69341
0 31906 7 1 2 49762 55224
0 31907 7 1 2 69716 31906
0 31908 7 1 2 70822 31907
0 31909 5 1 1 31908
0 31910 7 1 2 45624 51255
0 31911 7 1 2 64082 31910
0 31912 7 1 2 70722 31911
0 31913 5 1 1 31912
0 31914 7 1 2 57736 64191
0 31915 7 1 2 66042 31914
0 31916 7 1 2 68080 31915
0 31917 5 1 1 31916
0 31918 7 1 2 31913 31917
0 31919 5 1 1 31918
0 31920 7 1 2 43946 69455
0 31921 7 1 2 31919 31920
0 31922 5 1 1 31921
0 31923 7 1 2 31909 31922
0 31924 5 1 1 31923
0 31925 7 1 2 46536 31924
0 31926 5 1 1 31925
0 31927 7 2 2 59683 66486
0 31928 7 1 2 70719 70824
0 31929 7 1 2 70823 31928
0 31930 5 1 1 31929
0 31931 7 1 2 31926 31930
0 31932 5 1 1 31931
0 31933 7 1 2 70820 31932
0 31934 5 1 1 31933
0 31935 7 1 2 31903 31934
0 31936 5 1 1 31935
0 31937 7 1 2 45488 31936
0 31938 5 1 1 31937
0 31939 7 1 2 31874 31938
0 31940 7 1 2 31734 31939
0 31941 5 1 1 31940
0 31942 7 1 2 42228 31941
0 31943 5 1 1 31942
0 31944 7 2 2 44825 55500
0 31945 7 1 2 70791 70826
0 31946 5 1 1 31945
0 31947 7 2 2 45124 68645
0 31948 7 1 2 65033 70828
0 31949 5 1 1 31948
0 31950 7 1 2 49572 64919
0 31951 5 2 1 31950
0 31952 7 1 2 50137 56341
0 31953 5 1 1 31952
0 31954 7 1 2 70830 31953
0 31955 5 1 1 31954
0 31956 7 1 2 50476 31955
0 31957 5 1 1 31956
0 31958 7 1 2 31949 31957
0 31959 5 1 1 31958
0 31960 7 1 2 44101 31959
0 31961 5 1 1 31960
0 31962 7 1 2 52597 56579
0 31963 5 1 1 31962
0 31964 7 1 2 44102 64857
0 31965 7 1 2 31963 31964
0 31966 5 1 1 31965
0 31967 7 1 2 55687 31704
0 31968 7 1 2 31966 31967
0 31969 5 1 1 31968
0 31970 7 1 2 51285 31969
0 31971 5 1 1 31970
0 31972 7 1 2 48154 61980
0 31973 7 1 2 65383 31972
0 31974 5 1 1 31973
0 31975 7 1 2 31971 31974
0 31976 7 1 2 31961 31975
0 31977 5 1 1 31976
0 31978 7 1 2 44958 31977
0 31979 5 1 1 31978
0 31980 7 1 2 31946 31979
0 31981 5 2 1 31980
0 31982 7 1 2 67234 70832
0 31983 5 1 1 31982
0 31984 7 2 2 45489 70817
0 31985 7 1 2 51286 59791
0 31986 7 1 2 70834 31985
0 31987 5 1 1 31986
0 31988 7 1 2 31983 31987
0 31989 5 1 1 31988
0 31990 7 1 2 51668 31989
0 31991 5 1 1 31990
0 31992 7 2 2 45302 52490
0 31993 7 1 2 70812 70836
0 31994 5 1 1 31993
0 31995 7 1 2 52432 52598
0 31996 5 1 1 31995
0 31997 7 1 2 31994 31996
0 31998 5 1 1 31997
0 31999 7 1 2 59855 31998
0 32000 5 1 1 31999
0 32001 7 1 2 48481 62887
0 32002 5 1 1 32001
0 32003 7 1 2 64849 32002
0 32004 5 3 1 32003
0 32005 7 1 2 57402 70838
0 32006 5 1 1 32005
0 32007 7 1 2 58652 32006
0 32008 5 1 1 32007
0 32009 7 1 2 46093 61750
0 32010 7 1 2 32008 32009
0 32011 5 1 1 32010
0 32012 7 1 2 32000 32011
0 32013 5 1 1 32012
0 32014 7 1 2 57226 32013
0 32015 5 1 1 32014
0 32016 7 1 2 54060 64451
0 32017 7 1 2 64503 32016
0 32018 7 1 2 54679 61212
0 32019 7 1 2 32017 32018
0 32020 5 1 1 32019
0 32021 7 1 2 32015 32020
0 32022 5 1 1 32021
0 32023 7 1 2 43140 32022
0 32024 5 1 1 32023
0 32025 7 1 2 52389 59823
0 32026 5 1 1 32025
0 32027 7 1 2 59869 32026
0 32028 5 1 1 32027
0 32029 7 1 2 52425 64895
0 32030 7 1 2 32028 32029
0 32031 5 1 1 32030
0 32032 7 1 2 32024 32031
0 32033 5 1 1 32032
0 32034 7 1 2 51597 32033
0 32035 5 1 1 32034
0 32036 7 1 2 31991 32035
0 32037 5 1 1 32036
0 32038 7 1 2 69558 32037
0 32039 5 1 1 32038
0 32040 7 3 2 50428 60041
0 32041 7 1 2 45303 59884
0 32042 7 3 2 70841 32041
0 32043 7 1 2 55805 70844
0 32044 5 1 1 32043
0 32045 7 2 2 42605 55765
0 32046 7 2 2 57203 60183
0 32047 7 1 2 70847 70849
0 32048 5 1 1 32047
0 32049 7 1 2 32044 32048
0 32050 5 1 1 32049
0 32051 7 1 2 42067 32050
0 32052 5 1 1 32051
0 32053 7 1 2 45625 53654
0 32054 7 1 2 70845 32053
0 32055 5 1 1 32054
0 32056 7 1 2 32052 32055
0 32057 5 1 1 32056
0 32058 7 1 2 43141 32057
0 32059 5 1 1 32058
0 32060 7 2 2 64518 70850
0 32061 7 1 2 59696 70851
0 32062 5 1 1 32061
0 32063 7 1 2 32059 32062
0 32064 5 1 1 32063
0 32065 7 1 2 42887 32064
0 32066 5 1 1 32065
0 32067 7 2 2 43142 55766
0 32068 7 1 2 56292 59333
0 32069 7 1 2 70853 32068
0 32070 7 1 2 70769 32069
0 32071 5 1 1 32070
0 32072 7 1 2 32066 32071
0 32073 5 1 1 32072
0 32074 7 1 2 52649 32073
0 32075 5 1 1 32074
0 32076 7 2 2 51287 55131
0 32077 7 2 2 44357 56563
0 32078 7 1 2 55767 70857
0 32079 5 2 1 32078
0 32080 7 1 2 63754 70058
0 32081 7 1 2 70821 32080
0 32082 5 1 1 32081
0 32083 7 1 2 70859 32082
0 32084 5 1 1 32083
0 32085 7 1 2 42068 32084
0 32086 5 1 1 32085
0 32087 7 1 2 48482 57509
0 32088 7 1 2 63099 32087
0 32089 5 1 1 32088
0 32090 7 1 2 32086 32089
0 32091 5 1 1 32090
0 32092 7 1 2 70855 32091
0 32093 5 1 1 32092
0 32094 7 1 2 32075 32093
0 32095 5 1 1 32094
0 32096 7 1 2 54061 69076
0 32097 7 1 2 32095 32096
0 32098 5 1 1 32097
0 32099 7 1 2 32039 32098
0 32100 5 1 1 32099
0 32101 7 1 2 44488 32100
0 32102 5 1 1 32101
0 32103 7 1 2 55508 56612
0 32104 7 1 2 60252 32103
0 32105 5 1 1 32104
0 32106 7 1 2 70810 32105
0 32107 5 3 1 32106
0 32108 7 1 2 68363 70861
0 32109 5 1 1 32108
0 32110 7 1 2 51318 69127
0 32111 7 1 2 70807 32110
0 32112 5 1 1 32111
0 32113 7 1 2 32109 32112
0 32114 5 1 1 32113
0 32115 7 1 2 54801 59523
0 32116 7 1 2 32114 32115
0 32117 5 1 1 32116
0 32118 7 1 2 58653 5413
0 32119 5 2 1 32118
0 32120 7 2 2 60431 63755
0 32121 7 1 2 54392 63120
0 32122 7 1 2 64988 32121
0 32123 7 1 2 70866 32122
0 32124 7 1 2 70864 32123
0 32125 5 1 1 32124
0 32126 7 1 2 32117 32125
0 32127 5 1 1 32126
0 32128 7 1 2 61584 32127
0 32129 5 1 1 32128
0 32130 7 1 2 32102 32129
0 32131 5 1 1 32130
0 32132 7 1 2 42229 32131
0 32133 5 1 1 32132
0 32134 7 1 2 48835 52565
0 32135 7 1 2 64504 32134
0 32136 7 2 2 64330 32135
0 32137 7 1 2 67203 70868
0 32138 5 1 1 32137
0 32139 7 1 2 51377 61561
0 32140 7 3 2 56112 32139
0 32141 7 1 2 59128 70870
0 32142 5 1 1 32141
0 32143 7 1 2 32138 32142
0 32144 5 1 1 32143
0 32145 7 1 2 45626 32144
0 32146 5 1 1 32145
0 32147 7 1 2 51378 56023
0 32148 7 1 2 59372 32147
0 32149 7 2 2 31363 32148
0 32150 7 1 2 53678 70873
0 32151 5 1 1 32150
0 32152 7 1 2 32146 32151
0 32153 5 1 1 32152
0 32154 7 1 2 68364 32153
0 32155 5 1 1 32154
0 32156 7 2 2 51640 65610
0 32157 7 1 2 46319 69559
0 32158 7 1 2 70875 32157
0 32159 7 1 2 67170 32158
0 32160 5 1 1 32159
0 32161 7 1 2 32155 32160
0 32162 5 1 1 32161
0 32163 7 1 2 47804 32162
0 32164 5 1 1 32163
0 32165 7 2 2 55784 59885
0 32166 7 2 2 52168 52853
0 32167 7 2 2 70877 70879
0 32168 7 1 2 53564 69566
0 32169 5 1 1 32168
0 32170 7 1 2 53317 69077
0 32171 5 1 1 32170
0 32172 7 3 2 32169 32171
0 32173 7 1 2 54802 70883
0 32174 5 1 1 32173
0 32175 7 1 2 46859 51891
0 32176 7 1 2 68698 32175
0 32177 5 1 1 32176
0 32178 7 1 2 32174 32177
0 32179 5 1 1 32178
0 32180 7 2 2 70881 32179
0 32181 7 1 2 54223 70886
0 32182 5 1 1 32181
0 32183 7 1 2 32164 32182
0 32184 5 1 1 32183
0 32185 7 1 2 48483 32184
0 32186 5 1 1 32185
0 32187 7 1 2 56532 70887
0 32188 5 1 1 32187
0 32189 7 2 2 47687 44959
0 32190 7 1 2 47322 69431
0 32191 7 1 2 70888 32190
0 32192 7 2 2 55465 56133
0 32193 7 1 2 61485 66726
0 32194 7 1 2 70890 32193
0 32195 7 1 2 32191 32194
0 32196 5 1 1 32195
0 32197 7 1 2 54062 57143
0 32198 7 1 2 59727 32197
0 32199 5 1 1 32198
0 32200 7 1 2 43557 61833
0 32201 7 1 2 64447 32200
0 32202 7 1 2 64705 32201
0 32203 5 1 1 32202
0 32204 7 1 2 32199 32203
0 32205 5 1 1 32204
0 32206 7 1 2 57923 66783
0 32207 7 1 2 32205 32206
0 32208 5 1 1 32207
0 32209 7 1 2 32196 32208
0 32210 5 1 1 32209
0 32211 7 1 2 50146 32210
0 32212 5 1 1 32211
0 32213 7 1 2 32188 32212
0 32214 7 1 2 32186 32213
0 32215 5 1 1 32214
0 32216 7 1 2 53288 32215
0 32217 5 1 1 32216
0 32218 7 1 2 17425 17432
0 32219 5 3 1 32218
0 32220 7 1 2 48484 70892
0 32221 5 1 1 32220
0 32222 7 1 2 55745 69560
0 32223 5 1 1 32222
0 32224 7 1 2 32221 32223
0 32225 5 1 1 32224
0 32226 7 1 2 57889 70800
0 32227 7 1 2 64846 32226
0 32228 7 1 2 32225 32227
0 32229 5 1 1 32228
0 32230 7 1 2 58911 61924
0 32231 7 1 2 49870 32230
0 32232 7 2 2 47452 57029
0 32233 7 1 2 65511 70895
0 32234 7 1 2 32231 32233
0 32235 5 1 1 32234
0 32236 7 1 2 32229 32235
0 32237 5 1 1 32236
0 32238 7 1 2 48836 32237
0 32239 5 1 1 32238
0 32240 7 1 2 55850 68352
0 32241 7 1 2 70835 32240
0 32242 5 1 1 32241
0 32243 7 1 2 32239 32242
0 32244 5 1 1 32243
0 32245 7 1 2 51288 32244
0 32246 5 1 1 32245
0 32247 7 1 2 63968 64306
0 32248 7 1 2 65080 32247
0 32249 7 1 2 57932 32248
0 32250 5 1 1 32249
0 32251 7 2 2 45304 56191
0 32252 7 1 2 61975 70897
0 32253 7 1 2 70893 32252
0 32254 5 1 1 32253
0 32255 7 1 2 32250 32254
0 32256 5 1 1 32255
0 32257 7 1 2 42888 32256
0 32258 5 1 1 32257
0 32259 7 2 2 42341 53655
0 32260 7 1 2 49862 57924
0 32261 7 1 2 70899 32260
0 32262 7 1 2 69623 32261
0 32263 5 1 1 32262
0 32264 7 1 2 32258 32263
0 32265 5 1 1 32264
0 32266 7 1 2 43947 32265
0 32267 5 1 1 32266
0 32268 7 1 2 64530 64621
0 32269 7 1 2 55308 32268
0 32270 7 1 2 70854 32269
0 32271 5 1 1 32270
0 32272 7 1 2 32267 32271
0 32273 5 1 1 32272
0 32274 7 1 2 44960 32273
0 32275 5 1 1 32274
0 32276 7 1 2 56499 57925
0 32277 7 1 2 64707 32276
0 32278 5 1 1 32277
0 32279 7 3 2 47805 58026
0 32280 7 1 2 53632 64622
0 32281 7 1 2 70901 32280
0 32282 5 1 1 32281
0 32283 7 1 2 32278 32282
0 32284 5 1 1 32283
0 32285 7 1 2 58650 32284
0 32286 5 1 1 32285
0 32287 7 1 2 32275 32286
0 32288 5 1 1 32287
0 32289 7 1 2 70842 32288
0 32290 5 1 1 32289
0 32291 7 1 2 32246 32290
0 32292 5 1 1 32291
0 32293 7 1 2 45627 32292
0 32294 5 1 1 32293
0 32295 7 1 2 64922 64847
0 32296 7 1 2 65184 32295
0 32297 5 1 1 32296
0 32298 7 1 2 43948 67890
0 32299 7 1 2 70839 32298
0 32300 5 1 1 32299
0 32301 7 1 2 32297 32300
0 32302 5 1 1 32301
0 32303 7 1 2 43143 32302
0 32304 5 1 1 32303
0 32305 7 1 2 48155 49452
0 32306 7 1 2 62248 32305
0 32307 5 1 1 32306
0 32308 7 1 2 32304 32307
0 32309 5 1 1 32308
0 32310 7 1 2 66445 32309
0 32311 5 1 1 32310
0 32312 7 1 2 50429 65354
0 32313 5 1 1 32312
0 32314 7 1 2 31844 32313
0 32315 5 1 1 32314
0 32316 7 1 2 56527 63083
0 32317 7 1 2 64840 32316
0 32318 7 1 2 32315 32317
0 32319 5 1 1 32318
0 32320 7 1 2 32311 32319
0 32321 5 1 1 32320
0 32322 7 1 2 44961 32321
0 32323 5 1 1 32322
0 32324 7 1 2 64404 67957
0 32325 7 1 2 56147 32324
0 32326 7 1 2 65133 32325
0 32327 5 1 1 32326
0 32328 7 1 2 32323 32327
0 32329 5 1 1 32328
0 32330 7 1 2 54744 63786
0 32331 7 1 2 32329 32330
0 32332 5 1 1 32331
0 32333 7 1 2 32294 32332
0 32334 5 1 1 32333
0 32335 7 1 2 47688 32334
0 32336 5 1 1 32335
0 32337 7 1 2 55656 57638
0 32338 7 2 2 51478 32337
0 32339 7 1 2 57598 70904
0 32340 5 1 1 32339
0 32341 7 1 2 53482 64939
0 32342 5 1 1 32341
0 32343 7 1 2 54063 56906
0 32344 7 1 2 32342 32343
0 32345 5 1 1 32344
0 32346 7 1 2 32340 32345
0 32347 5 1 1 32346
0 32348 7 1 2 51152 32347
0 32349 5 1 1 32348
0 32350 7 1 2 2059 67727
0 32351 5 1 1 32350
0 32352 7 1 2 56907 59341
0 32353 7 1 2 67324 32352
0 32354 7 1 2 32351 32353
0 32355 5 1 1 32354
0 32356 7 1 2 32349 32355
0 32357 5 1 1 32356
0 32358 7 1 2 44826 32357
0 32359 5 1 1 32358
0 32360 7 1 2 48156 55191
0 32361 7 1 2 67958 32360
0 32362 7 1 2 70905 32361
0 32363 5 1 1 32362
0 32364 7 1 2 32359 32363
0 32365 5 1 1 32364
0 32366 7 1 2 48485 32365
0 32367 5 1 1 32366
0 32368 7 1 2 52068 57204
0 32369 7 1 2 53332 32368
0 32370 7 1 2 54123 32369
0 32371 5 1 1 32370
0 32372 7 1 2 70831 32371
0 32373 5 1 1 32372
0 32374 7 1 2 42606 32373
0 32375 5 1 1 32374
0 32376 7 1 2 51103 53948
0 32377 5 1 1 32376
0 32378 7 1 2 14355 32377
0 32379 5 1 1 32378
0 32380 7 1 2 70829 32379
0 32381 5 1 1 32380
0 32382 7 1 2 32375 32381
0 32383 5 1 1 32382
0 32384 7 1 2 44103 32383
0 32385 5 1 1 32384
0 32386 7 1 2 51289 58580
0 32387 5 1 1 32386
0 32388 7 1 2 49573 70762
0 32389 5 1 1 32388
0 32390 7 1 2 32387 32389
0 32391 5 1 1 32390
0 32392 7 1 2 51984 32391
0 32393 5 1 1 32392
0 32394 7 1 2 32385 32393
0 32395 5 1 1 32394
0 32396 7 1 2 44962 32395
0 32397 5 1 1 32396
0 32398 7 3 2 45305 50477
0 32399 7 1 2 52964 63948
0 32400 7 1 2 67719 32399
0 32401 7 1 2 70906 32400
0 32402 5 1 1 32401
0 32403 7 1 2 32397 32402
0 32404 5 1 1 32403
0 32405 7 1 2 55425 55851
0 32406 7 1 2 32404 32405
0 32407 5 1 1 32406
0 32408 7 1 2 32367 32407
0 32409 5 1 1 32408
0 32410 7 1 2 69561 32409
0 32411 5 1 1 32410
0 32412 7 1 2 56919 66580
0 32413 7 1 2 70862 32412
0 32414 5 1 1 32413
0 32415 7 1 2 32411 32414
0 32416 5 1 1 32415
0 32417 7 1 2 59856 32416
0 32418 5 1 1 32417
0 32419 7 1 2 32336 32418
0 32420 5 1 1 32419
0 32421 7 1 2 45767 32420
0 32422 5 1 1 32421
0 32423 7 1 2 32217 32422
0 32424 7 1 2 32133 32423
0 32425 5 1 1 32424
0 32426 7 1 2 66279 32425
0 32427 5 1 1 32426
0 32428 7 1 2 67146 70869
0 32429 5 1 1 32428
0 32430 7 1 2 67094 70871
0 32431 5 1 1 32430
0 32432 7 1 2 32429 32431
0 32433 5 1 1 32432
0 32434 7 1 2 45768 32433
0 32435 5 1 1 32434
0 32436 7 1 2 69657 70872
0 32437 5 1 1 32436
0 32438 7 1 2 32435 32437
0 32439 5 1 1 32438
0 32440 7 1 2 45628 32439
0 32441 5 1 1 32440
0 32442 7 1 2 69644 70874
0 32443 5 1 1 32442
0 32444 7 1 2 32441 32443
0 32445 5 1 1 32444
0 32446 7 1 2 70752 32445
0 32447 5 1 1 32446
0 32448 7 1 2 70876 70825
0 32449 7 1 2 69427 32448
0 32450 5 1 1 32449
0 32451 7 1 2 32447 32450
0 32452 5 1 1 32451
0 32453 7 1 2 47806 32452
0 32454 5 1 1 32453
0 32455 7 1 2 45629 69446
0 32456 5 1 1 32455
0 32457 7 1 2 69615 32456
0 32458 5 2 1 32457
0 32459 7 1 2 66016 70882
0 32460 7 2 2 70909 32459
0 32461 7 1 2 54224 70911
0 32462 5 1 1 32461
0 32463 7 1 2 32454 32462
0 32464 5 1 1 32463
0 32465 7 1 2 48486 32464
0 32466 5 1 1 32465
0 32467 7 1 2 56533 70912
0 32468 5 1 1 32467
0 32469 7 1 2 55492 67524
0 32470 7 1 2 63781 32469
0 32471 7 2 2 42069 63738
0 32472 7 1 2 68386 70913
0 32473 7 1 2 32470 32472
0 32474 5 1 1 32473
0 32475 7 1 2 57696 61275
0 32476 7 1 2 69172 70891
0 32477 7 1 2 32475 32476
0 32478 7 1 2 69816 32477
0 32479 5 1 1 32478
0 32480 7 1 2 32474 32479
0 32481 5 1 1 32480
0 32482 7 1 2 47323 32481
0 32483 5 1 1 32482
0 32484 7 1 2 57697 65814
0 32485 7 1 2 67779 32484
0 32486 7 1 2 70910 32485
0 32487 5 1 1 32486
0 32488 7 1 2 32483 32487
0 32489 5 1 1 32488
0 32490 7 1 2 50147 32489
0 32491 5 1 1 32490
0 32492 7 1 2 32468 32491
0 32493 7 1 2 32466 32492
0 32494 5 1 1 32493
0 32495 7 1 2 53289 32494
0 32496 5 1 1 32495
0 32497 7 1 2 68776 70846
0 32498 5 1 1 32497
0 32499 7 1 2 42409 51290
0 32500 7 1 2 67057 67371
0 32501 7 1 2 32499 32500
0 32502 5 1 1 32501
0 32503 7 1 2 32498 32502
0 32504 5 1 1 32503
0 32505 7 1 2 43144 32504
0 32506 5 1 1 32505
0 32507 7 1 2 70852 70796
0 32508 5 1 1 32507
0 32509 7 1 2 32506 32508
0 32510 5 1 1 32509
0 32511 7 1 2 42889 32510
0 32512 5 1 1 32511
0 32513 7 1 2 44827 49711
0 32514 7 1 2 67101 32513
0 32515 7 1 2 67058 70257
0 32516 7 1 2 32514 32515
0 32517 5 1 1 32516
0 32518 7 1 2 32512 32517
0 32519 5 1 1 32518
0 32520 7 1 2 52650 32519
0 32521 5 1 1 32520
0 32522 7 1 2 70858 70797
0 32523 5 1 1 32522
0 32524 7 1 2 49388 60003
0 32525 7 1 2 68777 32524
0 32526 5 1 1 32525
0 32527 7 1 2 32523 32526
0 32528 5 1 1 32527
0 32529 7 1 2 70856 32528
0 32530 5 1 1 32529
0 32531 7 1 2 32521 32530
0 32532 5 1 1 32531
0 32533 7 1 2 54064 65737
0 32534 7 1 2 32532 32533
0 32535 5 1 1 32534
0 32536 7 1 2 55485 60030
0 32537 7 1 2 70814 32536
0 32538 7 1 2 70733 32537
0 32539 5 1 1 32538
0 32540 7 2 2 57788 68778
0 32541 7 1 2 51405 52707
0 32542 7 1 2 54187 32541
0 32543 7 1 2 70915 32542
0 32544 5 1 1 32543
0 32545 7 1 2 32539 32544
0 32546 5 1 1 32545
0 32547 7 1 2 51291 32546
0 32548 5 1 1 32547
0 32549 7 5 2 48292 49574
0 32550 7 1 2 52944 70917
0 32551 5 1 1 32550
0 32552 7 1 2 43145 70840
0 32553 5 1 1 32552
0 32554 7 1 2 44104 51512
0 32555 5 1 1 32554
0 32556 7 1 2 32553 32555
0 32557 5 1 1 32556
0 32558 7 1 2 57403 32557
0 32559 5 1 1 32558
0 32560 7 1 2 32551 32559
0 32561 5 1 1 32560
0 32562 7 1 2 67891 70916
0 32563 7 1 2 32561 32562
0 32564 5 1 1 32563
0 32565 7 1 2 32548 32564
0 32566 5 1 1 32565
0 32567 7 1 2 47689 32566
0 32568 5 1 1 32567
0 32569 7 1 2 60184 63425
0 32570 7 2 2 66386 32569
0 32571 7 1 2 60053 70922
0 32572 7 1 2 70833 32571
0 32573 5 1 1 32572
0 32574 7 1 2 32568 32573
0 32575 5 1 1 32574
0 32576 7 1 2 65944 32575
0 32577 5 1 1 32576
0 32578 7 1 2 44489 32577
0 32579 7 1 2 32535 32578
0 32580 5 1 1 32579
0 32581 7 3 2 48035 66487
0 32582 5 2 1 70924
0 32583 7 1 2 59857 70925
0 32584 7 1 2 51319 32583
0 32585 7 1 2 70808 32584
0 32586 5 1 1 32585
0 32587 7 1 2 51302 68492
0 32588 7 1 2 70865 32587
0 32589 5 1 1 32588
0 32590 7 1 2 32586 32589
0 32591 5 1 1 32590
0 32592 7 1 2 44597 67027
0 32593 7 1 2 32591 32592
0 32594 5 1 1 32593
0 32595 7 1 2 61568 66869
0 32596 7 1 2 69342 32595
0 32597 7 1 2 70863 32596
0 32598 5 1 1 32597
0 32599 7 1 2 32594 32598
0 32600 5 1 1 32599
0 32601 7 1 2 45490 32600
0 32602 5 1 1 32601
0 32603 7 1 2 62888 70448
0 32604 5 1 1 32603
0 32605 7 1 2 68992 70483
0 32606 5 1 1 32605
0 32607 7 1 2 32604 32606
0 32608 5 1 1 32607
0 32609 7 1 2 51273 55426
0 32610 7 1 2 67986 32609
0 32611 7 1 2 70414 70726
0 32612 7 1 2 32610 32611
0 32613 7 1 2 32608 32612
0 32614 5 1 1 32613
0 32615 7 1 2 47807 32614
0 32616 7 1 2 32602 32615
0 32617 5 1 1 32616
0 32618 7 1 2 45769 32617
0 32619 7 1 2 32580 32618
0 32620 5 1 1 32619
0 32621 7 1 2 32496 32620
0 32622 7 1 2 32427 32621
0 32623 7 1 2 31943 32622
0 32624 5 1 1 32623
0 32625 7 1 2 55593 32624
0 32626 5 1 1 32625
0 32627 7 2 2 51570 63739
0 32628 7 1 2 60152 70929
0 32629 7 1 2 69131 32628
0 32630 5 1 1 32629
0 32631 7 1 2 53147 64001
0 32632 7 1 2 59957 32631
0 32633 7 1 2 69146 32632
0 32634 5 1 1 32633
0 32635 7 1 2 32630 32634
0 32636 5 1 1 32635
0 32637 7 1 2 69589 32636
0 32638 5 1 1 32637
0 32639 7 1 2 56435 57717
0 32640 7 1 2 63261 63748
0 32641 7 1 2 32639 32640
0 32642 5 1 1 32641
0 32643 7 1 2 32638 32642
0 32644 5 1 1 32643
0 32645 7 1 2 58533 32644
0 32646 5 1 1 32645
0 32647 7 1 2 42230 66788
0 32648 5 1 1 32647
0 32649 7 2 2 58890 66870
0 32650 5 1 1 70931
0 32651 7 1 2 32648 32650
0 32652 5 2 1 32651
0 32653 7 2 2 48293 62518
0 32654 7 1 2 68929 70935
0 32655 7 1 2 56516 32654
0 32656 7 1 2 70933 32655
0 32657 5 1 1 32656
0 32658 7 1 2 32646 32657
0 32659 5 1 1 32658
0 32660 7 1 2 67028 32659
0 32661 5 1 1 32660
0 32662 7 1 2 55192 59226
0 32663 7 1 2 68649 32662
0 32664 5 1 1 32663
0 32665 7 1 2 42607 52972
0 32666 7 1 2 55239 56472
0 32667 7 1 2 32665 32666
0 32668 5 1 1 32667
0 32669 7 1 2 32664 32668
0 32670 5 1 1 32669
0 32671 7 1 2 50195 65545
0 32672 7 1 2 32670 32671
0 32673 5 1 1 32672
0 32674 7 1 2 68520 69182
0 32675 7 1 2 70837 70896
0 32676 7 1 2 32674 32675
0 32677 5 1 1 32676
0 32678 7 1 2 32673 32677
0 32679 5 1 1 32678
0 32680 7 1 2 69343 32679
0 32681 5 1 1 32680
0 32682 7 2 2 42342 58400
0 32683 7 1 2 54600 70937
0 32684 5 1 1 32683
0 32685 7 1 2 49444 54627
0 32686 7 1 2 69125 32685
0 32687 5 1 1 32686
0 32688 7 1 2 32684 32687
0 32689 5 1 1 32688
0 32690 7 1 2 68782 32689
0 32691 5 1 1 32690
0 32692 7 1 2 55240 64002
0 32693 7 1 2 68807 32692
0 32694 5 1 1 32693
0 32695 7 1 2 32691 32694
0 32696 5 1 1 32695
0 32697 7 1 2 44598 32696
0 32698 5 1 1 32697
0 32699 7 2 2 51945 64049
0 32700 7 1 2 52657 69011
0 32701 5 1 1 32700
0 32702 7 1 2 55501 65081
0 32703 7 1 2 65280 32702
0 32704 5 1 1 32703
0 32705 7 1 2 32701 32704
0 32706 5 1 1 32705
0 32707 7 1 2 70939 32706
0 32708 5 1 1 32707
0 32709 7 1 2 32698 32708
0 32710 5 1 1 32709
0 32711 7 1 2 61953 70798
0 32712 7 1 2 32710 32711
0 32713 5 1 1 32712
0 32714 7 1 2 32681 32713
0 32715 7 1 2 32661 32714
0 32716 5 1 1 32715
0 32717 7 1 2 61562 32716
0 32718 5 1 1 32717
0 32719 7 1 2 60509 69150
0 32720 5 1 1 32719
0 32721 7 1 2 44963 53003
0 32722 5 1 1 32721
0 32723 7 1 2 54594 32722
0 32724 5 1 1 32723
0 32725 7 1 2 62519 32724
0 32726 5 1 1 32725
0 32727 7 1 2 32720 32726
0 32728 5 1 1 32727
0 32729 7 1 2 65738 32728
0 32730 5 1 1 32729
0 32731 7 1 2 52599 55134
0 32732 5 1 1 32731
0 32733 7 2 2 57461 64692
0 32734 7 1 2 53428 68114
0 32735 7 1 2 70941 32734
0 32736 7 1 2 32732 32735
0 32737 5 1 1 32736
0 32738 7 1 2 32730 32737
0 32739 5 1 1 32738
0 32740 7 1 2 42608 32739
0 32741 5 1 1 32740
0 32742 7 1 2 69772 70942
0 32743 5 1 1 32742
0 32744 7 2 2 55828 63024
0 32745 7 1 2 51348 57138
0 32746 7 1 2 70943 32745
0 32747 5 1 1 32746
0 32748 7 1 2 32743 32747
0 32749 5 1 1 32748
0 32750 7 1 2 48294 32749
0 32751 5 1 1 32750
0 32752 7 1 2 51349 57404
0 32753 7 1 2 65082 32752
0 32754 7 1 2 70944 32753
0 32755 5 1 1 32754
0 32756 7 1 2 32751 32755
0 32757 5 1 1 32756
0 32758 7 1 2 46094 32757
0 32759 5 1 1 32758
0 32760 7 1 2 44105 68457
0 32761 7 1 2 62478 32760
0 32762 7 1 2 68538 32761
0 32763 5 1 1 32762
0 32764 7 1 2 32759 32763
0 32765 5 1 1 32764
0 32766 7 1 2 42890 32765
0 32767 5 1 1 32766
0 32768 7 1 2 32741 32767
0 32769 5 1 1 32768
0 32770 7 1 2 48668 32769
0 32771 5 1 1 32770
0 32772 7 1 2 58316 70779
0 32773 7 1 2 69120 32772
0 32774 5 1 1 32773
0 32775 7 1 2 32771 32774
0 32776 5 1 1 32775
0 32777 7 1 2 59303 32776
0 32778 5 1 1 32777
0 32779 7 5 2 47915 61009
0 32780 7 1 2 60091 69137
0 32781 5 1 1 32780
0 32782 7 1 2 42891 68721
0 32783 5 1 1 32782
0 32784 7 1 2 32781 32783
0 32785 5 1 1 32784
0 32786 7 2 2 70945 32785
0 32787 7 1 2 64029 64071
0 32788 7 1 2 70950 32787
0 32789 5 1 1 32788
0 32790 7 1 2 32778 32789
0 32791 5 1 1 32790
0 32792 7 1 2 68174 32791
0 32793 5 1 1 32792
0 32794 7 1 2 64010 69152
0 32795 5 1 1 32794
0 32796 7 2 2 68976 70946
0 32797 7 2 2 63769 64758
0 32798 7 1 2 70952 70954
0 32799 5 1 1 32798
0 32800 7 1 2 32795 32799
0 32801 5 1 1 32800
0 32802 7 1 2 42609 32801
0 32803 5 1 1 32802
0 32804 7 1 2 55815 69773
0 32805 7 1 2 70955 32804
0 32806 5 1 1 32805
0 32807 7 1 2 50229 54505
0 32808 7 1 2 64011 32807
0 32809 5 1 1 32808
0 32810 7 1 2 32806 32809
0 32811 5 1 1 32810
0 32812 7 1 2 48295 32811
0 32813 5 1 1 32812
0 32814 7 2 2 43364 64003
0 32815 7 1 2 54464 56088
0 32816 7 1 2 58635 32815
0 32817 7 1 2 70956 32816
0 32818 5 1 1 32817
0 32819 7 1 2 32813 32818
0 32820 5 1 1 32819
0 32821 7 1 2 68680 32820
0 32822 5 1 1 32821
0 32823 7 1 2 32803 32822
0 32824 5 1 1 32823
0 32825 7 1 2 42070 32824
0 32826 5 1 1 32825
0 32827 7 1 2 43480 68312
0 32828 7 1 2 70951 32827
0 32829 5 1 1 32828
0 32830 7 1 2 32826 32829
0 32831 5 1 1 32830
0 32832 7 1 2 60649 32831
0 32833 5 1 1 32832
0 32834 7 1 2 53367 63740
0 32835 7 1 2 50521 32834
0 32836 7 1 2 55121 32835
0 32837 5 1 1 32836
0 32838 7 1 2 50165 60570
0 32839 7 1 2 60608 32838
0 32840 7 1 2 69705 32839
0 32841 5 1 1 32840
0 32842 7 1 2 32837 32841
0 32843 5 1 1 32842
0 32844 7 1 2 45630 32843
0 32845 5 1 1 32844
0 32846 7 1 2 50166 59179
0 32847 7 1 2 55448 32846
0 32848 7 1 2 68440 32847
0 32849 5 1 1 32848
0 32850 7 1 2 32845 32849
0 32851 5 1 1 32850
0 32852 7 1 2 67725 32851
0 32853 5 1 1 32852
0 32854 7 2 2 56311 67820
0 32855 7 1 2 56223 59557
0 32856 7 1 2 63180 32855
0 32857 7 1 2 70958 32856
0 32858 5 1 1 32857
0 32859 7 1 2 32853 32858
0 32860 5 1 1 32859
0 32861 7 1 2 42610 59166
0 32862 7 1 2 32860 32861
0 32863 5 1 1 32862
0 32864 7 1 2 32833 32863
0 32865 5 1 1 32864
0 32866 7 1 2 67029 32865
0 32867 5 1 1 32866
0 32868 7 2 2 70959 70691
0 32869 5 1 1 70960
0 32870 7 1 2 51379 56783
0 32871 7 1 2 68237 32870
0 32872 5 1 1 32871
0 32873 7 1 2 32869 32872
0 32874 5 1 1 32873
0 32875 7 1 2 50957 32874
0 32876 5 1 1 32875
0 32877 7 2 2 50522 68115
0 32878 7 1 2 65548 69141
0 32879 7 1 2 70962 32878
0 32880 5 1 1 32879
0 32881 7 1 2 32876 32880
0 32882 5 1 1 32881
0 32883 7 1 2 62603 32882
0 32884 5 1 1 32883
0 32885 7 3 2 45770 64030
0 32886 7 1 2 70953 70964
0 32887 5 1 1 32886
0 32888 7 2 2 43365 65546
0 32889 7 1 2 69153 70967
0 32890 5 1 1 32889
0 32891 7 1 2 32887 32890
0 32892 5 1 1 32891
0 32893 7 1 2 42611 32892
0 32894 5 1 1 32893
0 32895 7 2 2 69147 70968
0 32896 7 1 2 54616 70969
0 32897 5 1 1 32896
0 32898 7 1 2 64261 68998
0 32899 5 1 1 32898
0 32900 7 1 2 32897 32899
0 32901 5 1 1 32900
0 32902 7 1 2 68681 32901
0 32903 5 1 1 32902
0 32904 7 1 2 32894 32903
0 32905 5 1 1 32904
0 32906 7 1 2 59396 32905
0 32907 5 1 1 32906
0 32908 7 1 2 32884 32907
0 32909 5 1 1 32908
0 32910 7 1 2 67050 32909
0 32911 5 1 1 32910
0 32912 7 1 2 68753 70780
0 32913 5 1 1 32912
0 32914 7 2 2 49920 63025
0 32915 7 1 2 49389 58952
0 32916 7 1 2 70971 32915
0 32917 5 1 1 32916
0 32918 7 1 2 32913 32917
0 32919 5 1 1 32918
0 32920 7 1 2 56377 32919
0 32921 5 1 1 32920
0 32922 7 1 2 58326 64637
0 32923 7 1 2 69170 32922
0 32924 5 1 1 32923
0 32925 7 1 2 32921 32924
0 32926 5 1 1 32925
0 32927 7 1 2 44106 32926
0 32928 5 1 1 32927
0 32929 7 1 2 55006 58953
0 32930 7 1 2 50170 32929
0 32931 7 1 2 70717 32930
0 32932 5 1 1 32931
0 32933 7 1 2 32928 32932
0 32934 5 1 1 32933
0 32935 7 1 2 48296 32934
0 32936 5 1 1 32935
0 32937 7 2 2 62520 69066
0 32938 7 1 2 64160 70963
0 32939 7 1 2 70973 32938
0 32940 5 1 1 32939
0 32941 7 1 2 32936 32940
0 32942 5 1 1 32941
0 32943 7 1 2 51946 32942
0 32944 5 1 1 32943
0 32945 7 1 2 50167 56002
0 32946 7 1 2 57684 57846
0 32947 7 1 2 32945 32946
0 32948 7 1 2 69123 68674
0 32949 7 1 2 32947 32948
0 32950 5 1 1 32949
0 32951 7 1 2 32944 32950
0 32952 5 1 1 32951
0 32953 7 1 2 66919 32952
0 32954 5 1 1 32953
0 32955 7 1 2 32911 32954
0 32956 7 1 2 32867 32955
0 32957 7 1 2 32793 32956
0 32958 5 1 1 32957
0 32959 7 1 2 44828 32958
0 32960 5 1 1 32959
0 32961 7 1 2 32718 32960
0 32962 5 1 1 32961
0 32963 7 1 2 43766 32962
0 32964 5 1 1 32963
0 32965 7 1 2 62193 70455
0 32966 5 1 1 32965
0 32967 7 1 2 62135 66754
0 32968 7 1 2 65669 32967
0 32969 5 1 1 32968
0 32970 7 1 2 32966 32969
0 32971 5 1 1 32970
0 32972 7 1 2 51598 58647
0 32973 7 1 2 70470 32972
0 32974 7 1 2 32971 32973
0 32975 5 1 1 32974
0 32976 7 1 2 32964 32975
0 32977 5 1 1 32976
0 32978 7 1 2 49232 32977
0 32979 5 1 1 32978
0 32980 7 4 2 51599 65739
0 32981 5 1 1 70975
0 32982 7 1 2 49623 69504
0 32983 5 1 1 32982
0 32984 7 1 2 62374 32983
0 32985 5 1 1 32984
0 32986 7 1 2 54393 32985
0 32987 5 1 1 32986
0 32988 7 1 2 47453 55300
0 32989 5 1 1 32988
0 32990 7 1 2 53860 68732
0 32991 7 1 2 69500 32990
0 32992 7 1 2 32989 32991
0 32993 5 1 1 32992
0 32994 7 1 2 32987 32993
0 32995 5 1 1 32994
0 32996 7 1 2 70976 32995
0 32997 5 1 1 32996
0 32998 7 3 2 45491 51571
0 32999 7 1 2 55746 63297
0 33000 7 1 2 70979 32999
0 33001 7 1 2 69900 33000
0 33002 5 1 1 33001
0 33003 7 1 2 32997 33002
0 33004 5 1 1 33003
0 33005 7 1 2 44964 33004
0 33006 5 1 1 33005
0 33007 7 1 2 55193 70249
0 33008 7 1 2 69194 33007
0 33009 5 1 1 33008
0 33010 7 1 2 33006 33009
0 33011 5 1 1 33010
0 33012 7 1 2 48157 33011
0 33013 5 1 1 33012
0 33014 7 1 2 54316 56253
0 33015 7 1 2 68151 33014
0 33016 5 1 1 33015
0 33017 7 1 2 51669 60297
0 33018 7 1 2 69084 69185
0 33019 7 1 2 33017 33018
0 33020 5 1 1 33019
0 33021 7 1 2 33016 33020
0 33022 5 1 1 33021
0 33023 7 1 2 58097 68669
0 33024 7 1 2 33022 33023
0 33025 5 1 1 33024
0 33026 7 1 2 33013 33025
0 33027 5 1 1 33026
0 33028 7 1 2 66196 33027
0 33029 5 1 1 33028
0 33030 7 1 2 56614 66345
0 33031 7 1 2 69189 33030
0 33032 5 1 1 33031
0 33033 7 1 2 33029 33032
0 33034 5 1 1 33033
0 33035 7 1 2 45125 33034
0 33036 5 1 1 33035
0 33037 7 1 2 53810 70049
0 33038 5 1 1 33037
0 33039 7 1 2 50958 56696
0 33040 5 1 1 33039
0 33041 7 1 2 33038 33040
0 33042 5 1 1 33041
0 33043 7 2 2 42612 66931
0 33044 7 1 2 57847 67189
0 33045 7 1 2 50703 33044
0 33046 7 1 2 70982 33045
0 33047 7 1 2 33042 33046
0 33048 5 1 1 33047
0 33049 7 1 2 33036 33048
0 33050 5 1 1 33049
0 33051 7 1 2 42231 33050
0 33052 5 1 1 33051
0 33053 7 1 2 47916 70689
0 33054 7 1 2 68813 33053
0 33055 7 1 2 69190 33054
0 33056 5 1 1 33055
0 33057 7 1 2 33052 33056
0 33058 5 1 1 33057
0 33059 7 1 2 65664 33058
0 33060 5 1 1 33059
0 33061 7 1 2 32979 33060
0 33062 7 1 2 32626 33061
0 33063 7 1 2 31668 33062
0 33064 7 1 2 52271 56393
0 33065 7 1 2 58266 33064
0 33066 5 1 1 33065
0 33067 7 2 2 44490 62420
0 33068 7 1 2 57261 69999
0 33069 7 1 2 70984 33068
0 33070 5 1 1 33069
0 33071 7 1 2 33066 33070
0 33072 5 1 1 33071
0 33073 7 1 2 52600 33072
0 33074 5 1 1 33073
0 33075 7 1 2 55816 69330
0 33076 5 1 1 33075
0 33077 7 2 2 42232 60260
0 33078 7 1 2 50684 53148
0 33079 5 1 1 33078
0 33080 7 1 2 70986 33079
0 33081 5 1 1 33080
0 33082 7 1 2 33076 33081
0 33083 5 1 1 33082
0 33084 7 1 2 62521 33083
0 33085 5 1 1 33084
0 33086 7 1 2 42613 56323
0 33087 7 1 2 67108 33086
0 33088 5 1 1 33087
0 33089 7 1 2 33085 33088
0 33090 5 1 1 33089
0 33091 7 1 2 44965 33090
0 33092 5 1 1 33091
0 33093 7 1 2 64129 18263
0 33094 5 1 1 33093
0 33095 7 1 2 49822 69507
0 33096 7 1 2 33094 33095
0 33097 5 1 1 33096
0 33098 7 1 2 33092 33097
0 33099 5 1 1 33098
0 33100 7 1 2 42892 33099
0 33101 5 1 1 33100
0 33102 7 2 2 56538 70801
0 33103 7 1 2 45126 58487
0 33104 5 1 1 33103
0 33105 7 1 2 70000 33104
0 33106 7 1 2 70988 33105
0 33107 5 1 1 33106
0 33108 7 1 2 33101 33107
0 33109 5 1 1 33108
0 33110 7 1 2 44829 33109
0 33111 5 1 1 33110
0 33112 7 1 2 33074 33111
0 33113 5 1 1 33112
0 33114 7 1 2 44255 33113
0 33115 5 1 1 33114
0 33116 7 2 2 48837 68716
0 33117 7 2 2 45306 70990
0 33118 7 1 2 60458 70992
0 33119 5 1 1 33118
0 33120 7 1 2 59470 62522
0 33121 5 1 1 33120
0 33122 7 1 2 33119 33121
0 33123 5 1 1 33122
0 33124 7 1 2 59304 67708
0 33125 7 1 2 33123 33124
0 33126 5 1 1 33125
0 33127 7 1 2 33115 33126
0 33128 5 1 1 33127
0 33129 7 1 2 42343 33128
0 33130 5 1 1 33129
0 33131 7 1 2 44256 59305
0 33132 7 1 2 63217 33131
0 33133 7 1 2 54404 33132
0 33134 7 1 2 70974 33133
0 33135 5 1 1 33134
0 33136 7 1 2 33130 33135
0 33137 5 1 1 33136
0 33138 7 1 2 43366 33137
0 33139 5 1 1 33138
0 33140 7 4 2 42344 44830
0 33141 5 1 1 70994
0 33142 7 1 2 46746 62377
0 33143 5 1 1 33142
0 33144 7 1 2 56313 33143
0 33145 5 1 1 33144
0 33146 7 1 2 49662 33145
0 33147 5 1 1 33146
0 33148 7 1 2 43949 48980
0 33149 5 1 1 33148
0 33150 7 1 2 14155 33149
0 33151 5 1 1 33150
0 33152 7 1 2 42893 33151
0 33153 5 1 1 33152
0 33154 7 1 2 26308 33153
0 33155 5 1 1 33154
0 33156 7 1 2 44966 33155
0 33157 5 1 1 33156
0 33158 7 1 2 33147 33157
0 33159 5 1 1 33158
0 33160 7 1 2 62523 33159
0 33161 5 1 1 33160
0 33162 7 1 2 49632 57660
0 33163 7 2 2 68840 33162
0 33164 7 1 2 61452 66602
0 33165 7 1 2 70998 33164
0 33166 5 1 1 33165
0 33167 7 1 2 33161 33166
0 33168 5 1 1 33167
0 33169 7 1 2 42614 33168
0 33170 5 1 1 33169
0 33171 7 1 2 48297 58262
0 33172 7 1 2 60435 33171
0 33173 7 1 2 70999 33172
0 33174 5 1 1 33173
0 33175 7 1 2 33170 33174
0 33176 5 1 1 33175
0 33177 7 1 2 59306 33176
0 33178 5 1 1 33177
0 33179 7 2 2 48669 68717
0 33180 7 1 2 48838 71000
0 33181 5 1 1 33180
0 33182 7 1 2 58623 33181
0 33183 5 1 1 33182
0 33184 7 2 2 45771 55387
0 33185 7 1 2 60459 62846
0 33186 7 1 2 71002 33185
0 33187 7 1 2 33183 33186
0 33188 5 1 1 33187
0 33189 7 1 2 33178 33188
0 33190 5 1 1 33189
0 33191 7 1 2 70995 33190
0 33192 5 1 1 33191
0 33193 7 1 2 33139 33192
0 33194 5 1 1 33193
0 33195 7 1 2 44687 33194
0 33196 5 1 1 33195
0 33197 7 1 2 57112 67140
0 33198 5 1 1 33197
0 33199 7 1 2 55817 64957
0 33200 7 1 2 63718 33199
0 33201 5 1 1 33200
0 33202 7 1 2 33198 33201
0 33203 5 1 1 33202
0 33204 7 1 2 58247 33203
0 33205 5 1 1 33204
0 33206 7 1 2 58226 63549
0 33207 7 1 2 59120 33206
0 33208 5 1 1 33207
0 33209 7 1 2 33205 33208
0 33210 5 1 1 33209
0 33211 7 1 2 52651 33210
0 33212 5 1 1 33211
0 33213 7 1 2 42233 65127
0 33214 7 1 2 67206 70989
0 33215 7 1 2 33213 33214
0 33216 5 1 1 33215
0 33217 7 1 2 33212 33216
0 33218 5 1 1 33217
0 33219 7 1 2 69728 33218
0 33220 5 1 1 33219
0 33221 7 1 2 33196 33220
0 33222 5 1 1 33221
0 33223 7 1 2 68175 33222
0 33224 5 1 1 33223
0 33225 7 2 2 44831 65945
0 33226 7 2 2 56324 67467
0 33227 5 1 1 71006
0 33228 7 1 2 55685 61101
0 33229 5 1 1 33228
0 33230 7 1 2 33227 33229
0 33231 5 1 1 33230
0 33232 7 1 2 44967 33231
0 33233 5 1 1 33232
0 33234 7 1 2 52390 54735
0 33235 7 1 2 61102 33234
0 33236 5 1 1 33235
0 33237 7 1 2 33233 33236
0 33238 5 1 1 33237
0 33239 7 1 2 42615 33238
0 33240 5 1 1 33239
0 33241 7 1 2 52433 71007
0 33242 5 1 1 33241
0 33243 7 1 2 33240 33242
0 33244 5 1 1 33243
0 33245 7 1 2 44257 33244
0 33246 5 1 1 33245
0 33247 7 1 2 61826 63923
0 33248 7 1 2 58636 33247
0 33249 7 1 2 59993 33248
0 33250 5 1 1 33249
0 33251 7 1 2 33246 33250
0 33252 5 1 1 33251
0 33253 7 1 2 61055 33252
0 33254 5 1 1 33253
0 33255 7 1 2 67972 69060
0 33256 7 1 2 61615 33255
0 33257 7 1 2 70993 33256
0 33258 5 1 1 33257
0 33259 7 1 2 33254 33258
0 33260 5 1 1 33259
0 33261 7 1 2 43367 33260
0 33262 5 1 1 33261
0 33263 7 2 2 64565 68718
0 33264 7 1 2 64274 64803
0 33265 7 1 2 71008 33264
0 33266 5 1 1 33265
0 33267 7 1 2 56041 62866
0 33268 7 1 2 69144 33267
0 33269 7 1 2 62034 33268
0 33270 5 1 1 33269
0 33271 7 1 2 33266 33270
0 33272 5 1 1 33271
0 33273 7 1 2 52391 33272
0 33274 5 1 1 33273
0 33275 7 1 2 33262 33274
0 33276 5 1 1 33275
0 33277 7 1 2 71004 33276
0 33278 5 1 1 33277
0 33279 7 1 2 43368 69754
0 33280 5 1 1 33279
0 33281 7 1 2 65027 65113
0 33282 5 1 1 33281
0 33283 7 1 2 33280 33282
0 33284 5 1 1 33283
0 33285 7 1 2 60616 33284
0 33286 5 1 1 33285
0 33287 7 2 2 52652 57113
0 33288 7 1 2 63856 71010
0 33289 5 1 1 33288
0 33290 7 1 2 33286 33289
0 33291 5 1 1 33290
0 33292 7 1 2 48839 33291
0 33293 5 1 1 33292
0 33294 7 1 2 55790 61598
0 33295 7 1 2 65111 33294
0 33296 7 1 2 68759 33295
0 33297 5 1 1 33296
0 33298 7 1 2 33293 33297
0 33299 5 1 1 33298
0 33300 7 1 2 58227 33299
0 33301 5 1 1 33300
0 33302 7 1 2 48840 71011
0 33303 5 1 1 33302
0 33304 7 1 2 54332 33303
0 33305 5 1 1 33304
0 33306 7 1 2 57704 60837
0 33307 7 1 2 33305 33306
0 33308 5 1 1 33307
0 33309 7 1 2 33301 33308
0 33310 5 1 1 33309
0 33311 7 1 2 67709 33310
0 33312 5 1 1 33311
0 33313 7 1 2 56394 59605
0 33314 7 1 2 64917 33313
0 33315 7 2 2 42234 49575
0 33316 7 1 2 47808 49899
0 33317 7 1 2 71012 33316
0 33318 7 1 2 33314 33317
0 33319 5 1 1 33318
0 33320 7 1 2 33312 33319
0 33321 5 1 1 33320
0 33322 7 1 2 54803 33321
0 33323 5 1 1 33322
0 33324 7 1 2 55297 59116
0 33325 5 2 1 33324
0 33326 7 1 2 58725 71014
0 33327 5 1 1 33326
0 33328 7 1 2 52815 58732
0 33329 5 1 1 33328
0 33330 7 1 2 33327 33329
0 33331 5 1 1 33330
0 33332 7 1 2 59858 67710
0 33333 7 1 2 68719 33332
0 33334 7 1 2 33331 33333
0 33335 5 1 1 33334
0 33336 7 1 2 33323 33335
0 33337 5 1 1 33336
0 33338 7 1 2 65740 33337
0 33339 5 1 1 33338
0 33340 7 1 2 33278 33339
0 33341 5 1 1 33340
0 33342 7 1 2 67030 33341
0 33343 5 1 1 33342
0 33344 7 2 2 43369 53058
0 33345 5 2 1 71016
0 33346 7 1 2 69752 71018
0 33347 5 1 1 33346
0 33348 7 1 2 68238 33347
0 33349 5 1 1 33348
0 33350 7 1 2 62871 66488
0 33351 7 1 2 69859 33350
0 33352 5 1 1 33351
0 33353 7 1 2 33349 33352
0 33354 5 1 1 33353
0 33355 7 1 2 44968 33354
0 33356 5 1 1 33355
0 33357 7 1 2 43370 70961
0 33358 5 1 1 33357
0 33359 7 1 2 33356 33358
0 33360 5 1 1 33359
0 33361 7 1 2 60540 33360
0 33362 5 1 1 33361
0 33363 7 1 2 64958 70753
0 33364 5 1 1 33363
0 33365 7 1 2 24622 33364
0 33366 5 1 1 33365
0 33367 7 2 2 56325 33366
0 33368 7 1 2 54833 61653
0 33369 7 1 2 71020 33368
0 33370 5 1 1 33369
0 33371 7 1 2 33362 33370
0 33372 5 1 1 33371
0 33373 7 1 2 42616 33372
0 33374 5 1 1 33373
0 33375 7 1 2 60436 67966
0 33376 7 1 2 69371 33375
0 33377 7 1 2 71021 33376
0 33378 5 1 1 33377
0 33379 7 1 2 33374 33378
0 33380 5 1 1 33379
0 33381 7 1 2 44258 33380
0 33382 5 1 1 33381
0 33383 7 1 2 60650 64440
0 33384 7 1 2 70755 33383
0 33385 7 1 2 71009 33384
0 33386 5 1 1 33385
0 33387 7 1 2 33382 33386
0 33388 5 1 1 33387
0 33389 7 1 2 48841 33388
0 33390 5 1 1 33389
0 33391 7 1 2 60541 69750
0 33392 5 1 1 33391
0 33393 7 1 2 56326 59397
0 33394 5 1 1 33393
0 33395 7 1 2 33392 33394
0 33396 5 1 1 33395
0 33397 7 1 2 43371 33396
0 33398 5 1 1 33397
0 33399 7 1 2 50230 67818
0 33400 5 1 1 33399
0 33401 7 1 2 33398 33400
0 33402 5 1 1 33401
0 33403 7 1 2 58228 33402
0 33404 5 1 1 33403
0 33405 7 1 2 49823 52653
0 33406 7 1 2 58981 33405
0 33407 7 1 2 64187 33406
0 33408 5 1 1 33407
0 33409 7 1 2 33404 33408
0 33410 5 1 1 33409
0 33411 7 1 2 68239 33410
0 33412 5 1 1 33411
0 33413 7 1 2 56514 63121
0 33414 7 1 2 60688 33413
0 33415 7 1 2 70157 70640
0 33416 7 1 2 33414 33415
0 33417 5 1 1 33416
0 33418 7 1 2 33412 33417
0 33419 5 1 1 33418
0 33420 7 1 2 49233 33419
0 33421 5 1 1 33420
0 33422 7 1 2 42617 50231
0 33423 7 1 2 58314 33422
0 33424 7 1 2 63580 33423
0 33425 5 1 1 33424
0 33426 7 1 2 55662 69585
0 33427 5 1 1 33426
0 33428 7 1 2 63136 71001
0 33429 5 1 1 33428
0 33430 7 1 2 33427 33429
0 33431 5 1 1 33430
0 33432 7 1 2 57967 59373
0 33433 7 1 2 33431 33432
0 33434 5 1 1 33433
0 33435 7 1 2 33425 33434
0 33436 5 1 1 33435
0 33437 7 1 2 68234 33436
0 33438 5 1 1 33437
0 33439 7 1 2 33421 33438
0 33440 7 1 2 33390 33439
0 33441 5 1 1 33440
0 33442 7 1 2 44832 33441
0 33443 5 1 1 33442
0 33444 7 1 2 58482 65646
0 33445 7 3 2 44969 49576
0 33446 7 1 2 69892 70665
0 33447 7 1 2 71022 33446
0 33448 7 1 2 33444 33447
0 33449 5 1 1 33448
0 33450 7 1 2 33443 33449
0 33451 5 1 1 33450
0 33452 7 1 2 67051 33451
0 33453 5 1 1 33452
0 33454 7 2 2 52792 66588
0 33455 5 1 1 71025
0 33456 7 1 2 58229 69562
0 33457 7 1 2 52363 33456
0 33458 7 1 2 71026 33457
0 33459 5 1 1 33458
0 33460 7 1 2 53565 69078
0 33461 5 1 1 33460
0 33462 7 1 2 52797 69567
0 33463 5 1 1 33462
0 33464 7 3 2 33461 33463
0 33465 7 1 2 52809 56992
0 33466 7 1 2 58248 33465
0 33467 7 1 2 71027 33466
0 33468 5 1 1 33467
0 33469 7 1 2 33459 33468
0 33470 5 1 1 33469
0 33471 7 1 2 52654 33470
0 33472 5 1 1 33471
0 33473 7 1 2 52392 65606
0 33474 7 4 2 42235 64468
0 33475 7 2 2 45127 68116
0 33476 7 1 2 71030 71034
0 33477 7 1 2 33473 33476
0 33478 5 1 1 33477
0 33479 7 1 2 33472 33478
0 33480 5 1 1 33479
0 33481 7 1 2 44833 33480
0 33482 5 1 1 33481
0 33483 7 1 2 57255 59241
0 33484 7 1 2 54405 33483
0 33485 7 1 2 61619 71031
0 33486 7 1 2 33484 33485
0 33487 5 1 1 33486
0 33488 7 1 2 33482 33487
0 33489 5 1 1 33488
0 33490 7 1 2 68214 33489
0 33491 5 1 1 33490
0 33492 7 2 2 48298 63298
0 33493 7 1 2 65083 67831
0 33494 7 1 2 71036 33493
0 33495 5 1 1 33494
0 33496 7 1 2 57114 66789
0 33497 7 1 2 70991 33496
0 33498 5 1 1 33497
0 33499 7 1 2 33495 33498
0 33500 5 1 1 33499
0 33501 7 1 2 67711 33500
0 33502 5 1 1 33501
0 33503 7 1 2 45863 50706
0 33504 7 1 2 57120 69646
0 33505 7 1 2 33503 33504
0 33506 5 1 1 33505
0 33507 7 1 2 33502 33506
0 33508 5 1 1 33507
0 33509 7 1 2 53710 33508
0 33510 5 1 1 33509
0 33511 7 1 2 64566 65834
0 33512 7 1 2 54517 33511
0 33513 7 1 2 58249 33512
0 33514 7 1 2 69852 33513
0 33515 7 1 2 71015 33514
0 33516 5 1 1 33515
0 33517 7 1 2 33510 33516
0 33518 5 1 1 33517
0 33519 7 1 2 47809 33518
0 33520 5 1 1 33519
0 33521 7 1 2 33491 33520
0 33522 5 1 1 33521
0 33523 7 1 2 44358 33522
0 33524 5 1 1 33523
0 33525 7 1 2 51771 65159
0 33526 7 1 2 70102 33525
0 33527 5 1 1 33526
0 33528 7 1 2 49234 68760
0 33529 5 1 1 33528
0 33530 7 1 2 53543 62165
0 33531 5 1 1 33530
0 33532 7 2 2 71019 33531
0 33533 5 1 1 71038
0 33534 7 1 2 33529 71039
0 33535 5 1 1 33534
0 33536 7 1 2 54506 64623
0 33537 7 1 2 54804 33536
0 33538 7 1 2 33535 33537
0 33539 5 1 1 33538
0 33540 7 1 2 33527 33539
0 33541 5 1 1 33540
0 33542 7 1 2 48670 33541
0 33543 5 1 1 33542
0 33544 7 1 2 64624 68542
0 33545 7 1 2 71017 33544
0 33546 7 1 2 54819 33545
0 33547 5 1 1 33546
0 33548 7 1 2 33543 33547
0 33549 5 1 1 33548
0 33550 7 1 2 44970 33549
0 33551 5 1 1 33550
0 33552 7 1 2 57485 58202
0 33553 7 1 2 67821 69747
0 33554 7 1 2 33552 33553
0 33555 5 1 1 33554
0 33556 7 1 2 33551 33555
0 33557 5 1 1 33556
0 33558 7 1 2 56541 64505
0 33559 7 1 2 33557 33558
0 33560 5 1 1 33559
0 33561 7 1 2 33524 33560
0 33562 5 1 1 33561
0 33563 7 1 2 66280 33562
0 33564 5 1 1 33563
0 33565 7 1 2 68240 68761
0 33566 5 1 1 33565
0 33567 7 1 2 48036 65160
0 33568 7 1 2 70940 33567
0 33569 5 1 1 33568
0 33570 7 1 2 33566 33569
0 33571 5 1 1 33570
0 33572 7 1 2 49235 33571
0 33573 5 1 1 33572
0 33574 7 2 2 55427 66635
0 33575 7 1 2 63804 65161
0 33576 7 1 2 71040 33575
0 33577 5 1 1 33576
0 33578 7 1 2 68241 33533
0 33579 5 1 1 33578
0 33580 7 1 2 33577 33579
0 33581 7 1 2 33573 33580
0 33582 5 1 1 33581
0 33583 7 1 2 48671 33582
0 33584 5 1 1 33583
0 33585 7 1 2 42345 49427
0 33586 7 1 2 64266 33585
0 33587 7 1 2 68842 33586
0 33588 5 1 1 33587
0 33589 7 1 2 33584 33588
0 33590 5 1 1 33589
0 33591 7 1 2 44971 33590
0 33592 5 1 1 33591
0 33593 7 1 2 47324 53785
0 33594 7 4 2 58891 66577
0 33595 7 1 2 57486 71042
0 33596 7 1 2 33593 33595
0 33597 5 1 1 33596
0 33598 7 1 2 33592 33597
0 33599 5 1 1 33598
0 33600 7 3 2 63177 65861
0 33601 7 1 2 60503 64923
0 33602 7 1 2 71046 33601
0 33603 7 1 2 33599 33602
0 33604 5 1 1 33603
0 33605 7 1 2 33564 33604
0 33606 7 1 2 33453 33605
0 33607 7 1 2 33343 33606
0 33608 7 1 2 33224 33607
0 33609 5 1 1 33608
0 33610 7 1 2 43767 33609
0 33611 5 1 1 33610
0 33612 7 1 2 60744 64728
0 33613 7 1 2 66770 33612
0 33614 5 1 1 33613
0 33615 7 1 2 54609 55941
0 33616 5 1 1 33615
0 33617 7 1 2 56729 58098
0 33618 7 1 2 33616 33617
0 33619 5 1 1 33618
0 33620 7 1 2 33614 33619
0 33621 5 1 1 33620
0 33622 7 1 2 67991 69472
0 33623 7 2 2 44491 54507
0 33624 7 1 2 71032 71049
0 33625 7 1 2 33622 33624
0 33626 7 1 2 33621 33625
0 33627 5 1 1 33626
0 33628 7 1 2 33611 33627
0 33629 5 1 1 33628
0 33630 7 1 2 49353 33629
0 33631 5 1 1 33630
0 33632 7 2 2 49236 55917
0 33633 5 1 1 71051
0 33634 7 1 2 61465 71052
0 33635 5 1 1 33634
0 33636 7 1 2 57971 69539
0 33637 5 1 1 33636
0 33638 7 1 2 33635 33637
0 33639 5 1 1 33638
0 33640 7 1 2 51600 33639
0 33641 5 1 1 33640
0 33642 7 1 2 55402 56920
0 33643 7 1 2 62847 33642
0 33644 7 1 2 56107 33643
0 33645 5 1 1 33644
0 33646 7 1 2 33641 33645
0 33647 5 1 1 33646
0 33648 7 1 2 46747 33647
0 33649 5 1 1 33648
0 33650 7 2 2 55852 58067
0 33651 7 1 2 70172 71053
0 33652 7 1 2 62282 33651
0 33653 5 1 1 33652
0 33654 7 1 2 33649 33653
0 33655 5 1 1 33654
0 33656 7 1 2 43768 33655
0 33657 5 1 1 33656
0 33658 7 1 2 55918 70121
0 33659 7 1 2 50686 33658
0 33660 7 1 2 59091 33659
0 33661 5 1 1 33660
0 33662 7 1 2 33657 33661
0 33663 5 1 1 33662
0 33664 7 1 2 66197 33663
0 33665 5 1 1 33664
0 33666 7 3 2 45919 42618
0 33667 7 1 2 66145 71055
0 33668 7 1 2 59436 33667
0 33669 7 1 2 69590 33668
0 33670 7 1 2 66679 33669
0 33671 5 1 1 33670
0 33672 7 1 2 33665 33671
0 33673 5 1 1 33672
0 33674 7 1 2 45307 33673
0 33675 5 1 1 33674
0 33676 7 1 2 46537 50674
0 33677 7 1 2 63355 33676
0 33678 7 1 2 69436 33677
0 33679 5 1 1 33678
0 33680 7 1 2 33675 33679
0 33681 5 1 1 33680
0 33682 7 1 2 46320 33681
0 33683 5 1 1 33682
0 33684 7 2 2 46538 60139
0 33685 7 1 2 50313 71058
0 33686 5 1 1 33685
0 33687 7 1 2 50196 65016
0 33688 5 1 1 33687
0 33689 7 1 2 33686 33688
0 33690 5 1 1 33689
0 33691 7 1 2 47585 33690
0 33692 5 1 1 33691
0 33693 7 1 2 49712 65320
0 33694 5 1 1 33693
0 33695 7 1 2 33692 33694
0 33696 5 1 1 33695
0 33697 7 1 2 55933 70523
0 33698 7 1 2 33696 33697
0 33699 5 1 1 33698
0 33700 7 1 2 33683 33699
0 33701 5 1 1 33700
0 33702 7 1 2 42236 33701
0 33703 5 1 1 33702
0 33704 7 1 2 66680 66198
0 33705 5 1 1 33704
0 33706 7 1 2 66146 66371
0 33707 7 1 2 56972 33706
0 33708 5 1 1 33707
0 33709 7 1 2 33705 33708
0 33710 5 1 1 33709
0 33711 7 2 2 61206 69544
0 33712 7 1 2 55141 69432
0 33713 7 1 2 71060 33712
0 33714 7 1 2 33710 33713
0 33715 5 1 1 33714
0 33716 7 1 2 33703 33715
0 33717 5 1 1 33716
0 33718 7 1 2 65946 33717
0 33719 5 1 1 33718
0 33720 7 2 2 47917 57968
0 33721 7 1 2 56878 69540
0 33722 7 1 2 71062 33721
0 33723 7 1 2 67031 33722
0 33724 5 1 1 33723
0 33725 7 1 2 50335 60487
0 33726 7 1 2 62765 33725
0 33727 7 1 2 67095 33726
0 33728 5 1 1 33727
0 33729 7 1 2 33724 33728
0 33730 5 1 1 33729
0 33731 7 1 2 46748 33730
0 33732 5 1 1 33731
0 33733 7 1 2 61588 70338
0 33734 7 1 2 67096 33733
0 33735 5 1 1 33734
0 33736 7 1 2 33732 33735
0 33737 5 1 1 33736
0 33738 7 1 2 42237 33737
0 33739 5 1 1 33738
0 33740 7 1 2 67052 71063
0 33741 7 1 2 71061 33740
0 33742 5 1 1 33741
0 33743 7 1 2 33739 33742
0 33744 5 1 1 33743
0 33745 7 1 2 64452 65741
0 33746 7 1 2 33744 33745
0 33747 5 1 1 33746
0 33748 7 1 2 33719 33747
0 33749 5 1 1 33748
0 33750 7 1 2 42071 33749
0 33751 5 1 1 33750
0 33752 7 1 2 48945 68881
0 33753 5 1 1 33752
0 33754 7 1 2 47918 65807
0 33755 7 1 2 68819 33754
0 33756 5 1 1 33755
0 33757 7 1 2 33753 33756
0 33758 5 1 1 33757
0 33759 7 1 2 56031 64336
0 33760 7 1 2 69545 33759
0 33761 7 1 2 33758 33760
0 33762 5 1 1 33761
0 33763 7 1 2 33751 33762
0 33764 5 1 1 33763
0 33765 7 1 2 44359 33764
0 33766 5 1 1 33765
0 33767 7 1 2 65791 65817
0 33768 5 2 1 33767
0 33769 7 1 2 60770 71064
0 33770 5 1 1 33769
0 33771 7 4 2 45864 50168
0 33772 7 1 2 56356 71066
0 33773 5 2 1 33772
0 33774 7 1 2 33770 71070
0 33775 5 1 1 33774
0 33776 7 1 2 47454 33775
0 33777 5 1 1 33776
0 33778 7 1 2 48842 62471
0 33779 7 1 2 63287 33778
0 33780 5 1 1 33779
0 33781 7 1 2 33777 33780
0 33782 5 1 1 33781
0 33783 7 1 2 45308 33782
0 33784 5 1 1 33783
0 33785 7 1 2 51406 70316
0 33786 5 2 1 33785
0 33787 7 1 2 63391 70021
0 33788 5 1 1 33787
0 33789 7 1 2 71072 33788
0 33790 5 1 1 33789
0 33791 7 1 2 55594 33790
0 33792 5 1 1 33791
0 33793 7 1 2 43146 60162
0 33794 5 1 1 33793
0 33795 7 1 2 63711 33794
0 33796 5 1 1 33795
0 33797 7 1 2 65808 33796
0 33798 5 1 1 33797
0 33799 7 1 2 33792 33798
0 33800 7 1 2 33784 33799
0 33801 5 1 1 33800
0 33802 7 1 2 58726 33801
0 33803 5 1 1 33802
0 33804 7 1 2 61062 65947
0 33805 5 1 1 33804
0 33806 7 1 2 62472 69106
0 33807 5 1 1 33806
0 33808 7 1 2 33805 33807
0 33809 5 1 1 33808
0 33810 7 1 2 48672 33809
0 33811 5 1 1 33810
0 33812 7 1 2 57723 65742
0 33813 5 2 1 33812
0 33814 7 1 2 33811 71074
0 33815 5 1 1 33814
0 33816 7 1 2 46539 33815
0 33817 5 1 1 33816
0 33818 7 1 2 66093 68889
0 33819 5 1 1 33818
0 33820 7 1 2 47455 68484
0 33821 5 1 1 33820
0 33822 7 1 2 33819 33821
0 33823 5 1 1 33822
0 33824 7 1 2 45309 33823
0 33825 5 2 1 33824
0 33826 7 1 2 33817 71076
0 33827 5 1 1 33826
0 33828 7 1 2 61056 33827
0 33829 5 1 1 33828
0 33830 7 1 2 33803 33829
0 33831 5 1 1 33830
0 33832 7 1 2 45631 33831
0 33833 5 1 1 33832
0 33834 7 2 2 57077 64594
0 33835 5 1 1 71078
0 33836 7 1 2 66017 33835
0 33837 5 2 1 33836
0 33838 7 1 2 55493 64307
0 33839 5 2 1 33838
0 33840 7 1 2 51407 66018
0 33841 5 1 1 33840
0 33842 7 1 2 71082 33841
0 33843 5 1 1 33842
0 33844 7 1 2 50102 33843
0 33845 5 1 1 33844
0 33846 7 1 2 71080 33845
0 33847 5 1 1 33846
0 33848 7 1 2 55785 59022
0 33849 7 1 2 33847 33848
0 33850 5 1 1 33849
0 33851 7 1 2 33833 33850
0 33852 5 1 1 33851
0 33853 7 1 2 46860 33852
0 33854 5 1 1 33853
0 33855 7 1 2 58547 65948
0 33856 5 1 1 33855
0 33857 7 1 2 71081 33856
0 33858 5 1 1 33857
0 33859 7 1 2 43481 55786
0 33860 7 1 2 61276 33859
0 33861 7 1 2 33858 33860
0 33862 5 1 1 33861
0 33863 7 1 2 33854 33862
0 33864 5 1 1 33863
0 33865 7 1 2 47690 33864
0 33866 5 1 1 33865
0 33867 7 2 2 52253 58733
0 33868 5 1 1 71084
0 33869 7 1 2 56660 58727
0 33870 5 1 1 33869
0 33871 7 1 2 33868 33870
0 33872 5 1 1 33871
0 33873 7 3 2 54667 63403
0 33874 7 1 2 33872 71086
0 33875 5 1 1 33874
0 33876 7 1 2 48913 71085
0 33877 5 1 1 33876
0 33878 7 1 2 49842 54484
0 33879 5 1 1 33878
0 33880 7 1 2 54805 62228
0 33881 5 1 1 33880
0 33882 7 1 2 33879 33881
0 33883 5 1 1 33882
0 33884 7 1 2 51862 33883
0 33885 5 1 1 33884
0 33886 7 1 2 59455 61817
0 33887 5 1 1 33886
0 33888 7 1 2 33885 33887
0 33889 5 1 1 33888
0 33890 7 1 2 49763 33889
0 33891 5 1 1 33890
0 33892 7 3 2 45772 55412
0 33893 7 1 2 70427 71089
0 33894 5 1 1 33893
0 33895 7 1 2 60893 63528
0 33896 5 1 1 33895
0 33897 7 1 2 33894 33896
0 33898 5 1 1 33897
0 33899 7 1 2 42072 33898
0 33900 5 1 1 33899
0 33901 7 1 2 46749 63627
0 33902 5 1 1 33901
0 33903 7 1 2 47919 64743
0 33904 7 1 2 65208 33903
0 33905 7 1 2 33902 33904
0 33906 5 1 1 33905
0 33907 7 1 2 33900 33906
0 33908 7 1 2 33891 33907
0 33909 5 1 1 33908
0 33910 7 1 2 47810 33909
0 33911 5 1 1 33910
0 33912 7 1 2 33877 33911
0 33913 5 1 1 33912
0 33914 7 1 2 65949 33913
0 33915 5 1 1 33914
0 33916 7 1 2 33875 33915
0 33917 5 1 1 33916
0 33918 7 1 2 44360 33917
0 33919 5 1 1 33918
0 33920 7 1 2 62569 70380
0 33921 5 1 1 33920
0 33922 7 2 2 55672 69743
0 33923 7 1 2 68313 71092
0 33924 5 1 1 33923
0 33925 7 3 2 44688 63653
0 33926 7 1 2 69893 71094
0 33927 5 1 1 33926
0 33928 7 1 2 33924 33927
0 33929 5 1 1 33928
0 33930 7 1 2 62607 33929
0 33931 5 1 1 33930
0 33932 7 1 2 33921 33931
0 33933 7 1 2 33919 33932
0 33934 7 1 2 33866 33933
0 33935 5 1 1 33934
0 33936 7 1 2 42894 33935
0 33937 5 1 1 33936
0 33938 7 1 2 64289 65095
0 33939 5 1 1 33938
0 33940 7 1 2 48673 33939
0 33941 5 1 1 33940
0 33942 7 1 2 52254 57523
0 33943 5 1 1 33942
0 33944 7 1 2 33941 33943
0 33945 5 1 1 33944
0 33946 7 1 2 70695 33945
0 33947 5 1 1 33946
0 33948 7 1 2 52086 64775
0 33949 5 1 1 33948
0 33950 7 1 2 70107 33949
0 33951 5 1 1 33950
0 33952 7 1 2 65743 33951
0 33953 5 1 1 33952
0 33954 7 1 2 61066 69939
0 33955 5 1 1 33954
0 33956 7 1 2 48674 33955
0 33957 5 1 1 33956
0 33958 7 1 2 64905 33957
0 33959 5 1 1 33958
0 33960 7 1 2 44107 33959
0 33961 5 1 1 33960
0 33962 7 1 2 28215 33961
0 33963 5 1 1 33962
0 33964 7 1 2 65950 33963
0 33965 5 1 1 33964
0 33966 7 1 2 33953 33965
0 33967 5 1 1 33966
0 33968 7 1 2 58728 33967
0 33969 5 1 1 33968
0 33970 7 1 2 33947 33969
0 33971 5 1 1 33970
0 33972 7 1 2 59859 33971
0 33973 5 1 1 33972
0 33974 7 1 2 62306 70390
0 33975 5 2 1 33974
0 33976 7 1 2 60617 71097
0 33977 5 1 1 33976
0 33978 7 1 2 63857 69934
0 33979 5 1 1 33978
0 33980 7 1 2 33977 33979
0 33981 5 1 1 33980
0 33982 7 1 2 49713 33981
0 33983 5 1 1 33982
0 33984 7 1 2 50619 57365
0 33985 7 1 2 63879 33984
0 33986 5 1 1 33985
0 33987 7 1 2 33983 33986
0 33988 5 1 1 33987
0 33989 7 1 2 66019 33988
0 33990 5 1 1 33989
0 33991 7 1 2 61074 61839
0 33992 5 1 1 33991
0 33993 7 1 2 44108 33992
0 33994 5 1 1 33993
0 33995 7 1 2 64906 33994
0 33996 5 1 1 33995
0 33997 7 1 2 69456 33996
0 33998 5 1 1 33997
0 33999 7 2 2 46321 56752
0 34000 5 1 1 71099
0 34001 7 1 2 69759 34000
0 34002 5 1 1 34001
0 34003 7 1 2 48843 34002
0 34004 5 1 1 34003
0 34005 7 1 2 55540 59078
0 34006 5 2 1 34005
0 34007 7 1 2 51508 71101
0 34008 5 1 1 34007
0 34009 7 1 2 34004 34008
0 34010 5 1 1 34009
0 34011 7 1 2 44109 34010
0 34012 5 1 1 34011
0 34013 7 1 2 43147 60197
0 34014 5 1 1 34013
0 34015 7 1 2 5134 34014
0 34016 7 1 2 34012 34015
0 34017 5 1 1 34016
0 34018 7 1 2 65951 34017
0 34019 5 1 1 34018
0 34020 7 1 2 33998 34019
0 34021 5 1 1 34020
0 34022 7 1 2 63858 34021
0 34023 5 1 1 34022
0 34024 7 1 2 33990 34023
0 34025 5 1 1 34024
0 34026 7 1 2 54806 34025
0 34027 5 1 1 34026
0 34028 7 1 2 68953 29316
0 34029 5 1 1 34028
0 34030 7 1 2 61057 34029
0 34031 5 1 1 34030
0 34032 7 1 2 60571 64200
0 34033 7 1 2 69767 34032
0 34034 5 1 1 34033
0 34035 7 1 2 34031 34034
0 34036 5 1 1 34035
0 34037 7 1 2 50959 34036
0 34038 5 1 1 34037
0 34039 7 1 2 56428 64648
0 34040 7 1 2 68783 34039
0 34041 7 1 2 52923 34040
0 34042 5 1 1 34041
0 34043 7 1 2 34038 34042
0 34044 5 1 1 34043
0 34045 7 1 2 49237 34044
0 34046 5 1 1 34045
0 34047 7 1 2 59227 70957
0 34048 5 1 1 34047
0 34049 7 1 2 61058 68981
0 34050 5 1 1 34049
0 34051 7 1 2 34048 34050
0 34052 5 1 1 34051
0 34053 7 1 2 49115 52411
0 34054 5 1 1 34053
0 34055 7 1 2 44110 34054
0 34056 5 1 1 34055
0 34057 7 1 2 48675 60705
0 34058 5 1 1 34057
0 34059 7 1 2 34056 34058
0 34060 5 1 1 34059
0 34061 7 1 2 34052 34060
0 34062 5 1 1 34061
0 34063 7 1 2 47811 63084
0 34064 7 1 2 64959 34063
0 34065 7 1 2 69177 34064
0 34066 7 1 2 62283 34065
0 34067 5 1 1 34066
0 34068 7 1 2 34062 34067
0 34069 7 1 2 34046 34068
0 34070 5 1 1 34069
0 34071 7 1 2 61103 34070
0 34072 5 1 1 34071
0 34073 7 1 2 34027 34072
0 34074 7 1 2 33973 34073
0 34075 7 1 2 33937 34074
0 34076 5 1 1 34075
0 34077 7 1 2 67032 34076
0 34078 5 1 1 34077
0 34079 7 1 2 70055 29196
0 34080 5 1 1 34079
0 34081 7 1 2 59792 34080
0 34082 5 1 1 34081
0 34083 7 1 2 59860 30584
0 34084 5 1 1 34083
0 34085 7 1 2 34082 34084
0 34086 5 1 1 34085
0 34087 7 1 2 66887 34086
0 34088 5 1 1 34087
0 34089 7 1 2 6015 66825
0 34090 5 1 1 34089
0 34091 7 1 2 50308 55328
0 34092 7 1 2 66840 34091
0 34093 5 1 1 34092
0 34094 7 1 2 34090 34093
0 34095 5 1 1 34094
0 34096 7 1 2 46750 34095
0 34097 5 1 1 34096
0 34098 7 1 2 58362 66826
0 34099 5 1 1 34098
0 34100 7 1 2 49095 66841
0 34101 5 1 1 34100
0 34102 7 1 2 34099 34101
0 34103 5 1 1 34102
0 34104 7 1 2 53368 34103
0 34105 5 1 1 34104
0 34106 7 1 2 34097 34105
0 34107 5 1 1 34106
0 34108 7 1 2 48676 34107
0 34109 5 1 1 34108
0 34110 7 1 2 50869 66842
0 34111 5 1 1 34110
0 34112 7 1 2 66819 68324
0 34113 5 1 1 34112
0 34114 7 1 2 34111 34113
0 34115 5 1 1 34114
0 34116 7 1 2 48677 34115
0 34117 5 1 1 34116
0 34118 7 1 2 48844 66843
0 34119 5 1 1 34118
0 34120 7 3 2 63222 66820
0 34121 5 1 1 71103
0 34122 7 1 2 34119 34121
0 34123 7 1 2 34117 34122
0 34124 5 1 1 34123
0 34125 7 1 2 71100 34124
0 34126 5 1 1 34125
0 34127 7 1 2 34109 34126
0 34128 5 1 1 34127
0 34129 7 1 2 44111 34128
0 34130 5 1 1 34129
0 34131 7 1 2 58551 71079
0 34132 5 2 1 34131
0 34133 7 1 2 66827 71106
0 34134 5 1 1 34133
0 34135 7 1 2 45492 70378
0 34136 5 1 1 34135
0 34137 7 1 2 60168 34136
0 34138 5 1 1 34137
0 34139 7 1 2 66844 34138
0 34140 5 1 1 34139
0 34141 7 1 2 34134 34140
0 34142 5 1 1 34141
0 34143 7 1 2 42895 34142
0 34144 5 1 1 34143
0 34145 7 1 2 42346 70402
0 34146 5 1 1 34145
0 34147 7 1 2 57534 71104
0 34148 5 1 1 34147
0 34149 7 1 2 34146 34148
0 34150 5 1 1 34149
0 34151 7 1 2 50016 34150
0 34152 5 1 1 34151
0 34153 7 1 2 34144 34152
0 34154 7 1 2 34130 34153
0 34155 5 1 1 34154
0 34156 7 1 2 54807 34155
0 34157 5 1 1 34156
0 34158 7 1 2 51734 53798
0 34159 5 1 1 34158
0 34160 7 1 2 70105 34159
0 34161 5 1 1 34160
0 34162 7 1 2 66881 34161
0 34163 5 1 1 34162
0 34164 7 1 2 66873 30580
0 34165 5 1 1 34164
0 34166 7 1 2 34163 34165
0 34167 5 1 1 34166
0 34168 7 1 2 59861 34167
0 34169 5 1 1 34168
0 34170 7 1 2 34157 34169
0 34171 7 1 2 34088 34170
0 34172 5 1 1 34171
0 34173 7 1 2 53613 34172
0 34174 5 1 1 34173
0 34175 7 1 2 68135 70559
0 34176 5 1 1 34175
0 34177 7 1 2 69984 70556
0 34178 5 2 1 34177
0 34179 7 1 2 43372 71108
0 34180 5 1 1 34179
0 34181 7 1 2 49593 70027
0 34182 5 1 1 34181
0 34183 7 1 2 34180 34182
0 34184 5 1 1 34183
0 34185 7 1 2 66554 34184
0 34186 5 1 1 34185
0 34187 7 1 2 34176 34186
0 34188 5 1 1 34187
0 34189 7 1 2 44259 34188
0 34190 5 1 1 34189
0 34191 7 2 2 53429 68365
0 34192 7 1 2 60728 71110
0 34193 5 1 1 34192
0 34194 7 1 2 49488 55545
0 34195 5 1 1 34194
0 34196 7 1 2 65472 34195
0 34197 5 1 1 34196
0 34198 7 1 2 46540 34197
0 34199 5 1 1 34198
0 34200 7 1 2 28693 34199
0 34201 5 1 1 34200
0 34202 7 1 2 66555 34201
0 34203 5 1 1 34202
0 34204 7 1 2 34193 34203
0 34205 5 1 1 34204
0 34206 7 1 2 48678 34205
0 34207 5 1 1 34206
0 34208 7 1 2 59066 66502
0 34209 5 1 1 34208
0 34210 7 1 2 50103 60768
0 34211 7 1 2 66556 34210
0 34212 5 1 1 34211
0 34213 7 1 2 34209 34212
0 34214 5 1 1 34213
0 34215 7 1 2 54898 34214
0 34216 5 1 1 34215
0 34217 7 1 2 34207 34216
0 34218 7 1 2 34190 34217
0 34219 5 1 1 34218
0 34220 7 1 2 59445 34219
0 34221 5 1 1 34220
0 34222 7 1 2 50104 68366
0 34223 5 1 1 34222
0 34224 7 1 2 69110 34223
0 34225 5 1 1 34224
0 34226 7 1 2 53730 34225
0 34227 5 1 1 34226
0 34228 7 1 2 68367 28305
0 34229 5 1 1 34228
0 34230 7 1 2 34227 34229
0 34231 7 1 2 69926 34230
0 34232 5 1 1 34231
0 34233 7 1 2 59733 34232
0 34234 5 1 1 34233
0 34235 7 1 2 44492 34234
0 34236 7 1 2 34221 34235
0 34237 5 1 1 34236
0 34238 7 1 2 47586 70450
0 34239 5 1 1 34238
0 34240 7 1 2 59701 34239
0 34241 5 2 1 34240
0 34242 7 1 2 46751 71112
0 34243 5 1 1 34242
0 34244 7 1 2 43373 70464
0 34245 5 2 1 34244
0 34246 7 1 2 34243 71114
0 34247 5 1 1 34246
0 34248 7 1 2 66557 34247
0 34249 5 1 1 34248
0 34250 7 1 2 44112 61076
0 34251 5 1 1 34250
0 34252 7 1 2 64907 34251
0 34253 5 3 1 34252
0 34254 7 1 2 69922 71116
0 34255 5 1 1 34254
0 34256 7 2 2 49714 54237
0 34257 7 1 2 66790 71119
0 34258 5 1 1 34257
0 34259 7 2 2 48946 61992
0 34260 7 1 2 42347 71121
0 34261 5 1 1 34260
0 34262 7 1 2 34258 34261
0 34263 5 1 1 34262
0 34264 7 1 2 50870 34263
0 34265 5 1 1 34264
0 34266 7 1 2 34255 34265
0 34267 7 1 2 34249 34266
0 34268 5 1 1 34267
0 34269 7 1 2 67171 34268
0 34270 5 1 1 34269
0 34271 7 1 2 42896 60198
0 34272 5 1 1 34271
0 34273 7 1 2 70580 34272
0 34274 5 1 1 34273
0 34275 7 1 2 66558 34274
0 34276 5 1 1 34275
0 34277 7 1 2 49125 68301
0 34278 7 1 2 70022 34277
0 34279 5 1 1 34278
0 34280 7 1 2 34276 34279
0 34281 5 1 1 34280
0 34282 7 1 2 46541 34281
0 34283 5 1 1 34282
0 34284 7 1 2 61538 66503
0 34285 7 1 2 70566 34284
0 34286 5 1 1 34285
0 34287 7 1 2 34283 34286
0 34288 5 1 1 34287
0 34289 7 1 2 70008 34288
0 34290 5 1 1 34289
0 34291 7 1 2 47812 34290
0 34292 7 1 2 34270 34291
0 34293 5 1 1 34292
0 34294 7 1 2 34237 34293
0 34295 5 1 1 34294
0 34296 7 1 2 64609 69116
0 34297 5 1 1 34296
0 34298 7 1 2 45773 59725
0 34299 7 1 2 61785 66504
0 34300 7 1 2 34298 34299
0 34301 5 1 1 34300
0 34302 7 1 2 34297 34301
0 34303 5 1 1 34302
0 34304 7 1 2 42073 34303
0 34305 5 1 1 34304
0 34306 7 1 2 56993 64432
0 34307 7 1 2 70481 34306
0 34308 7 1 2 53679 34307
0 34309 5 1 1 34308
0 34310 7 1 2 34305 34309
0 34311 5 1 1 34310
0 34312 7 1 2 50620 34311
0 34313 5 1 1 34312
0 34314 7 1 2 63600 65419
0 34315 5 1 1 34314
0 34316 7 2 2 44689 67935
0 34317 7 1 2 64050 71123
0 34318 7 1 2 34315 34317
0 34319 7 1 2 58141 34318
0 34320 5 1 1 34319
0 34321 7 1 2 34313 34320
0 34322 5 1 1 34321
0 34323 7 1 2 44493 34322
0 34324 5 1 1 34323
0 34325 7 2 2 56134 61599
0 34326 7 1 2 58865 71125
0 34327 7 1 2 69108 34326
0 34328 7 1 2 63610 34327
0 34329 5 1 1 34328
0 34330 7 1 2 34324 34329
0 34331 5 1 1 34330
0 34332 7 1 2 49238 34331
0 34333 5 1 1 34332
0 34334 7 1 2 50621 69870
0 34335 5 1 1 34334
0 34336 7 1 2 70005 70473
0 34337 5 1 1 34336
0 34338 7 1 2 34335 34337
0 34339 5 1 1 34338
0 34340 7 1 2 43374 34339
0 34341 5 1 1 34340
0 34342 7 1 2 70160 70002
0 34343 5 1 1 34342
0 34344 7 1 2 34341 34343
0 34345 5 1 1 34344
0 34346 7 1 2 66559 34345
0 34347 5 1 1 34346
0 34348 7 1 2 57462 64625
0 34349 7 1 2 71124 34348
0 34350 7 1 2 58322 34349
0 34351 5 1 1 34350
0 34352 7 1 2 34347 34351
0 34353 5 1 1 34352
0 34354 7 1 2 49096 34353
0 34355 5 1 1 34354
0 34356 7 1 2 34333 34355
0 34357 7 1 2 34295 34356
0 34358 7 1 2 34174 34357
0 34359 5 1 1 34358
0 34360 7 1 2 66281 34359
0 34361 5 1 1 34360
0 34362 7 1 2 66101 71113
0 34363 5 1 1 34362
0 34364 7 1 2 49354 51195
0 34365 5 1 1 34364
0 34366 7 1 2 59068 64872
0 34367 7 1 2 34365 34366
0 34368 5 1 1 34367
0 34369 7 1 2 48679 34368
0 34370 5 1 1 34369
0 34371 7 1 2 51716 57823
0 34372 5 2 1 34371
0 34373 7 1 2 54909 71127
0 34374 7 1 2 34370 34373
0 34375 5 1 1 34374
0 34376 7 1 2 65744 34375
0 34377 5 1 1 34376
0 34378 7 1 2 70462 34377
0 34379 5 1 1 34378
0 34380 7 1 2 68982 34379
0 34381 5 1 1 34380
0 34382 7 1 2 34363 34381
0 34383 5 1 1 34382
0 34384 7 1 2 59398 34383
0 34385 5 1 1 34384
0 34386 7 1 2 48680 71098
0 34387 5 1 1 34386
0 34388 7 1 2 65351 34387
0 34389 5 1 1 34388
0 34390 7 1 2 44113 34389
0 34391 5 1 1 34390
0 34392 7 1 2 42897 71107
0 34393 5 1 1 34392
0 34394 7 1 2 70327 34393
0 34395 7 1 2 34391 34394
0 34396 5 1 1 34395
0 34397 7 1 2 70586 34396
0 34398 5 1 1 34397
0 34399 7 1 2 34385 34398
0 34400 5 1 1 34399
0 34401 7 1 2 59307 34400
0 34402 5 1 1 34401
0 34403 7 1 2 69457 71117
0 34404 5 1 1 34403
0 34405 7 1 2 49097 64372
0 34406 5 1 1 34405
0 34407 7 1 2 63873 34406
0 34408 5 1 1 34407
0 34409 7 1 2 43375 34408
0 34410 5 2 1 34409
0 34411 7 1 2 52323 64950
0 34412 5 1 1 34411
0 34413 7 1 2 57356 59767
0 34414 5 1 1 34413
0 34415 7 1 2 34412 34414
0 34416 7 1 2 71129 34415
0 34417 5 1 1 34416
0 34418 7 1 2 65952 34417
0 34419 5 1 1 34418
0 34420 7 1 2 34404 34419
0 34421 5 1 1 34420
0 34422 7 1 2 59399 34421
0 34423 5 1 1 34422
0 34424 7 1 2 58677 65953
0 34425 5 1 1 34424
0 34426 7 1 2 67004 34425
0 34427 5 1 1 34426
0 34428 7 1 2 51509 34427
0 34429 5 1 1 34428
0 34430 7 1 2 47587 66085
0 34431 5 1 1 34430
0 34432 7 1 2 67005 34431
0 34433 5 1 1 34432
0 34434 7 1 2 51408 34433
0 34435 5 1 1 34434
0 34436 7 1 2 34429 34435
0 34437 5 1 1 34436
0 34438 7 1 2 55388 34437
0 34439 5 1 1 34438
0 34440 7 1 2 55202 61916
0 34441 5 1 1 34440
0 34442 7 1 2 58618 34441
0 34443 5 1 1 34442
0 34444 7 1 2 65745 34443
0 34445 5 1 1 34444
0 34446 7 1 2 42898 60073
0 34447 7 1 2 34445 34446
0 34448 5 1 1 34447
0 34449 7 1 2 43148 59768
0 34450 5 1 1 34449
0 34451 7 1 2 46322 1140
0 34452 7 1 2 34450 34451
0 34453 5 1 1 34452
0 34454 7 1 2 68983 34453
0 34455 7 1 2 34448 34454
0 34456 5 1 1 34455
0 34457 7 1 2 34439 34456
0 34458 5 1 1 34457
0 34459 7 1 2 60542 34458
0 34460 5 1 1 34459
0 34461 7 1 2 34423 34460
0 34462 5 1 1 34461
0 34463 7 1 2 51947 34462
0 34464 5 1 1 34463
0 34465 7 1 2 63918 64278
0 34466 5 1 1 34465
0 34467 7 1 2 67077 70560
0 34468 5 1 1 34467
0 34469 7 1 2 34466 34468
0 34470 5 1 1 34469
0 34471 7 1 2 68950 34470
0 34472 5 1 1 34471
0 34473 7 1 2 61955 64177
0 34474 5 1 1 34473
0 34475 7 1 2 1143 59400
0 34476 7 1 2 70305 34475
0 34477 5 1 1 34476
0 34478 7 1 2 34474 34477
0 34479 5 1 1 34478
0 34480 7 1 2 71043 34479
0 34481 5 1 1 34480
0 34482 7 1 2 34472 34481
0 34483 5 1 1 34482
0 34484 7 1 2 49239 34483
0 34485 5 1 1 34484
0 34486 7 1 2 70756 71120
0 34487 5 1 1 34486
0 34488 7 1 2 63741 71122
0 34489 5 1 1 34488
0 34490 7 1 2 34487 34489
0 34491 5 1 1 34490
0 34492 7 1 2 59401 34491
0 34493 5 1 1 34492
0 34494 7 2 2 56429 61010
0 34495 7 1 2 69160 69681
0 34496 7 1 2 71131 34495
0 34497 5 1 1 34496
0 34498 7 1 2 34493 34497
0 34499 5 1 1 34498
0 34500 7 1 2 50871 34499
0 34501 5 1 1 34500
0 34502 7 1 2 34485 34501
0 34503 7 1 2 34464 34502
0 34504 7 1 2 34402 34503
0 34505 5 1 1 34504
0 34506 7 1 2 67053 34505
0 34507 5 1 1 34506
0 34508 7 3 2 51948 66020
0 34509 5 1 1 71133
0 34510 7 1 2 46323 62116
0 34511 5 1 1 34510
0 34512 7 1 2 70282 34511
0 34513 5 1 1 34512
0 34514 7 1 2 71134 34513
0 34515 5 1 1 34514
0 34516 7 1 2 66120 70084
0 34517 5 1 1 34516
0 34518 7 1 2 48845 50131
0 34519 7 1 2 71065 34518
0 34520 5 1 1 34519
0 34521 7 1 2 34517 34520
0 34522 5 1 1 34521
0 34523 7 1 2 46324 34522
0 34524 5 1 1 34523
0 34525 7 1 2 55317 70926
0 34526 5 1 1 34525
0 34527 7 1 2 42899 58418
0 34528 7 1 2 65809 34527
0 34529 5 1 1 34528
0 34530 7 1 2 34526 34529
0 34531 5 1 1 34530
0 34532 7 1 2 46752 34531
0 34533 5 1 1 34532
0 34534 7 1 2 34524 34533
0 34535 5 1 1 34534
0 34536 7 1 2 59308 34535
0 34537 5 1 1 34536
0 34538 7 1 2 34515 34537
0 34539 5 1 1 34538
0 34540 7 1 2 44114 34539
0 34541 5 1 1 34540
0 34542 7 1 2 61063 63949
0 34543 5 1 1 34542
0 34544 7 1 2 18938 34543
0 34545 5 1 1 34544
0 34546 7 1 2 67110 34545
0 34547 5 1 1 34546
0 34548 7 1 2 34541 34547
0 34549 5 1 1 34548
0 34550 7 1 2 48681 34549
0 34551 5 1 1 34550
0 34552 7 1 2 55535 69028
0 34553 7 1 2 71102 34552
0 34554 5 1 1 34553
0 34555 7 1 2 70319 34554
0 34556 5 1 1 34555
0 34557 7 1 2 59309 34556
0 34558 5 1 1 34557
0 34559 7 1 2 61466 71044
0 34560 7 1 2 58377 34559
0 34561 5 1 1 34560
0 34562 7 1 2 34558 34561
0 34563 5 1 1 34562
0 34564 7 1 2 54899 34563
0 34565 5 1 1 34564
0 34566 7 1 2 57945 64119
0 34567 7 1 2 51356 34566
0 34568 7 1 2 64782 34567
0 34569 5 1 1 34568
0 34570 7 1 2 34565 34569
0 34571 7 1 2 34551 34570
0 34572 5 1 1 34571
0 34573 7 1 2 66920 34572
0 34574 5 1 1 34573
0 34575 7 1 2 52854 68176
0 34576 5 1 1 34575
0 34577 7 1 2 63611 66921
0 34578 5 1 1 34577
0 34579 7 1 2 34576 34578
0 34580 5 1 1 34579
0 34581 7 1 2 43149 34580
0 34582 5 1 1 34581
0 34583 7 1 2 67097 69965
0 34584 5 1 1 34583
0 34585 7 1 2 34582 34584
0 34586 5 1 1 34585
0 34587 7 1 2 65746 34586
0 34588 5 1 1 34587
0 34589 7 2 2 55768 66736
0 34590 7 1 2 67179 71136
0 34591 7 1 2 70307 34590
0 34592 5 1 1 34591
0 34593 7 1 2 34588 34592
0 34594 5 1 1 34593
0 34595 7 1 2 59310 34594
0 34596 5 1 1 34595
0 34597 7 1 2 54238 65747
0 34598 5 1 1 34597
0 34599 7 1 2 70927 34598
0 34600 5 1 1 34599
0 34601 7 1 2 59334 62934
0 34602 7 1 2 67098 34601
0 34603 7 1 2 34600 34602
0 34604 5 1 1 34603
0 34605 7 1 2 34596 34604
0 34606 5 1 1 34605
0 34607 7 1 2 50872 34606
0 34608 5 1 1 34607
0 34609 7 1 2 62935 71118
0 34610 5 1 1 34609
0 34611 7 1 2 64290 64777
0 34612 5 1 1 34611
0 34613 7 1 2 48682 34612
0 34614 5 1 1 34613
0 34615 7 1 2 63507 71128
0 34616 7 1 2 34614 34615
0 34617 5 1 1 34616
0 34618 7 1 2 59311 34617
0 34619 5 1 1 34618
0 34620 7 1 2 34610 34619
0 34621 5 1 1 34620
0 34622 7 1 2 65748 34621
0 34623 5 1 1 34622
0 34624 7 1 2 49183 58508
0 34625 5 1 1 34624
0 34626 7 1 2 65137 34625
0 34627 5 1 1 34626
0 34628 7 1 2 46753 34627
0 34629 5 1 1 34628
0 34630 7 1 2 70574 71130
0 34631 7 1 2 34629 34630
0 34632 5 1 1 34631
0 34633 7 1 2 51949 34632
0 34634 5 1 1 34633
0 34635 7 1 2 59312 61723
0 34636 5 1 1 34635
0 34637 7 1 2 63965 34636
0 34638 5 1 1 34637
0 34639 7 1 2 50790 34638
0 34640 5 1 1 34639
0 34641 7 1 2 58337 62900
0 34642 5 1 1 34641
0 34643 7 1 2 34640 34642
0 34644 5 1 1 34643
0 34645 7 1 2 50622 34644
0 34646 5 1 1 34645
0 34647 7 1 2 53731 61756
0 34648 5 1 1 34647
0 34649 7 1 2 59702 34648
0 34650 5 1 1 34649
0 34651 7 1 2 46754 34650
0 34652 5 1 1 34651
0 34653 7 1 2 71115 34652
0 34654 5 1 1 34653
0 34655 7 1 2 59313 34654
0 34656 5 1 1 34655
0 34657 7 1 2 34646 34656
0 34658 7 1 2 34634 34657
0 34659 5 1 1 34658
0 34660 7 1 2 65954 34659
0 34661 5 1 1 34660
0 34662 7 1 2 34623 34661
0 34663 5 1 1 34662
0 34664 7 1 2 68177 34663
0 34665 5 1 1 34664
0 34666 7 1 2 34608 34665
0 34667 7 1 2 34574 34666
0 34668 5 1 1 34667
0 34669 7 1 2 60460 34668
0 34670 5 1 1 34669
0 34671 7 1 2 45865 1903
0 34672 5 1 1 34671
0 34673 7 1 2 57094 69568
0 34674 7 1 2 34672 34673
0 34675 5 1 1 34674
0 34676 7 1 2 71075 34675
0 34677 5 1 1 34676
0 34678 7 1 2 46542 34677
0 34679 5 1 1 34678
0 34680 7 1 2 71077 34679
0 34681 5 1 1 34680
0 34682 7 1 2 42900 34681
0 34683 5 1 1 34682
0 34684 7 1 2 66982 68954
0 34685 5 1 1 34684
0 34686 7 1 2 49240 34685
0 34687 5 1 1 34686
0 34688 7 1 2 62278 68984
0 34689 5 1 1 34688
0 34690 7 1 2 34687 34689
0 34691 5 1 1 34690
0 34692 7 1 2 56723 34691
0 34693 5 1 1 34692
0 34694 7 1 2 34683 34693
0 34695 5 1 1 34694
0 34696 7 1 2 51670 70291
0 34697 7 1 2 34695 34696
0 34698 5 1 1 34697
0 34699 7 1 2 43605 50623
0 34700 7 1 2 70321 34699
0 34701 7 1 2 71137 34700
0 34702 5 1 1 34701
0 34703 7 1 2 70028 70785
0 34704 7 1 2 66922 34703
0 34705 5 1 1 34704
0 34706 7 1 2 34702 34705
0 34707 5 1 1 34706
0 34708 7 1 2 59314 34707
0 34709 5 1 1 34708
0 34710 7 1 2 51510 60918
0 34711 7 1 2 67131 34710
0 34712 7 1 2 70980 70724
0 34713 7 1 2 34711 34712
0 34714 5 1 1 34713
0 34715 7 1 2 34709 34714
0 34716 5 1 1 34715
0 34717 7 1 2 55595 34716
0 34718 5 1 1 34717
0 34719 7 1 2 65270 68178
0 34720 5 1 1 34719
0 34721 7 2 2 46942 57771
0 34722 5 1 1 71138
0 34723 7 1 2 66147 71139
0 34724 7 1 2 70532 34723
0 34725 5 1 1 34724
0 34726 7 1 2 34720 34725
0 34727 5 1 1 34726
0 34728 7 1 2 65955 34727
0 34729 5 1 1 34728
0 34730 7 1 2 65862 67668
0 34731 7 1 2 63840 34730
0 34732 7 1 2 69346 34731
0 34733 5 1 1 34732
0 34734 7 1 2 34729 34733
0 34735 5 1 1 34734
0 34736 7 1 2 50624 34735
0 34737 5 1 1 34736
0 34738 7 1 2 3675 63538
0 34739 7 1 2 65347 34738
0 34740 5 1 1 34739
0 34741 7 1 2 68179 70744
0 34742 7 1 2 34740 34741
0 34743 5 1 1 34742
0 34744 7 1 2 34737 34743
0 34745 7 1 2 34718 34744
0 34746 7 1 2 70748 34509
0 34747 5 1 1 34746
0 34748 7 1 2 68180 34747
0 34749 5 1 1 34748
0 34750 7 2 2 59315 66021
0 34751 5 2 1 71140
0 34752 7 1 2 51950 65819
0 34753 5 1 1 34752
0 34754 7 1 2 71142 34753
0 34755 5 1 1 34754
0 34756 7 1 2 52905 66923
0 34757 7 1 2 34755 34756
0 34758 5 1 1 34757
0 34759 7 1 2 34749 34758
0 34760 5 1 1 34759
0 34761 7 1 2 42901 34760
0 34762 5 1 1 34761
0 34763 7 1 2 66958 70707
0 34764 5 1 1 34763
0 34765 7 1 2 34762 34764
0 34766 5 1 1 34765
0 34767 7 1 2 50105 34766
0 34768 5 1 1 34767
0 34769 7 1 2 63919 66959
0 34770 5 1 1 34769
0 34771 7 1 2 67896 70329
0 34772 7 1 2 71109 34771
0 34773 5 1 1 34772
0 34774 7 1 2 34770 34773
0 34775 5 1 1 34774
0 34776 7 1 2 50017 34775
0 34777 5 1 1 34776
0 34778 7 1 2 60004 60678
0 34779 7 1 2 69535 34778
0 34780 7 1 2 70096 34779
0 34781 5 1 1 34780
0 34782 7 1 2 55818 66944
0 34783 7 1 2 67533 34782
0 34784 5 1 1 34783
0 34785 7 1 2 34781 34784
0 34786 7 1 2 34777 34785
0 34787 5 1 1 34786
0 34788 7 1 2 66022 34787
0 34789 5 1 1 34788
0 34790 7 1 2 34768 34789
0 34791 7 1 2 34745 34790
0 34792 7 1 2 34698 34791
0 34793 5 1 1 34792
0 34794 7 1 2 62524 34793
0 34795 5 1 1 34794
0 34796 7 1 2 34670 34795
0 34797 7 1 2 34507 34796
0 34798 7 1 2 34361 34797
0 34799 7 1 2 34078 34798
0 34800 5 1 1 34799
0 34801 7 1 2 53290 34800
0 34802 5 1 1 34801
0 34803 7 2 2 44361 67128
0 34804 7 1 2 58378 71144
0 34805 5 1 1 34804
0 34806 7 1 2 42619 60026
0 34807 7 1 2 51236 34806
0 34808 7 1 2 71047 34807
0 34809 5 1 1 34808
0 34810 7 1 2 34805 34809
0 34811 5 1 1 34810
0 34812 7 1 2 43769 34811
0 34813 5 1 1 34812
0 34814 7 1 2 62122 68181
0 34815 5 1 1 34814
0 34816 7 1 2 34813 34815
0 34817 5 1 1 34816
0 34818 7 1 2 50564 34817
0 34819 5 1 1 34818
0 34820 7 1 2 49715 60104
0 34821 7 1 2 66387 34820
0 34822 7 1 2 58591 62721
0 34823 7 1 2 34821 34822
0 34824 5 1 1 34823
0 34825 7 1 2 34819 34824
0 34826 5 1 1 34825
0 34827 7 1 2 46325 34826
0 34828 5 1 1 34827
0 34829 7 1 2 46755 70612
0 34830 5 1 1 34829
0 34831 7 1 2 43376 57554
0 34832 7 1 2 58363 34831
0 34833 7 1 2 65101 34832
0 34834 5 1 1 34833
0 34835 7 1 2 34830 34834
0 34836 5 1 1 34835
0 34837 7 1 2 42902 68182
0 34838 7 1 2 34836 34837
0 34839 5 1 1 34838
0 34840 7 1 2 34828 34839
0 34841 5 1 1 34840
0 34842 7 1 2 42074 34841
0 34843 5 1 1 34842
0 34844 7 2 2 53861 61235
0 34845 7 1 2 54137 63092
0 34846 7 1 2 71146 34845
0 34847 7 1 2 51237 34846
0 34848 7 1 2 67054 34847
0 34849 5 1 1 34848
0 34850 7 1 2 34843 34849
0 34851 5 1 1 34850
0 34852 7 1 2 51951 34851
0 34853 5 1 1 34852
0 34854 7 1 2 55344 70907
0 34855 5 1 1 34854
0 34856 7 1 2 65478 34855
0 34857 5 3 1 34856
0 34858 7 1 2 57314 71148
0 34859 5 1 1 34858
0 34860 7 1 2 51185 65339
0 34861 5 1 1 34860
0 34862 7 1 2 60853 34861
0 34863 5 2 1 34862
0 34864 7 1 2 63977 71151
0 34865 5 1 1 34864
0 34866 7 1 2 34859 34865
0 34867 5 1 1 34866
0 34868 7 1 2 43150 34867
0 34869 5 1 1 34868
0 34870 7 4 2 45493 63612
0 34871 7 1 2 60060 71153
0 34872 5 1 1 34871
0 34873 7 1 2 34869 34872
0 34874 5 1 1 34873
0 34875 7 1 2 51863 59210
0 34876 7 1 2 34874 34875
0 34877 5 1 1 34876
0 34878 7 1 2 60572 63237
0 34879 7 1 2 70059 34878
0 34880 7 1 2 70209 34879
0 34881 5 1 1 34880
0 34882 7 1 2 34877 34881
0 34883 5 1 1 34882
0 34884 7 1 2 42075 34883
0 34885 5 1 1 34884
0 34886 7 1 2 50106 62570
0 34887 5 1 1 34886
0 34888 7 1 2 62848 64970
0 34889 5 1 1 34888
0 34890 7 1 2 34887 34889
0 34891 5 1 1 34890
0 34892 7 1 2 49304 34891
0 34893 5 1 1 34892
0 34894 7 1 2 47588 55711
0 34895 7 1 2 71090 34894
0 34896 5 1 1 34895
0 34897 7 1 2 34893 34896
0 34898 5 1 1 34897
0 34899 7 2 2 59994 60855
0 34900 7 1 2 51031 71157
0 34901 7 1 2 34898 34900
0 34902 5 1 1 34901
0 34903 7 1 2 34885 34902
0 34904 5 1 1 34903
0 34905 7 1 2 67033 34904
0 34906 5 1 1 34905
0 34907 7 1 2 56042 60005
0 34908 7 1 2 60856 34907
0 34909 7 1 2 70207 34908
0 34910 7 1 2 70734 34909
0 34911 5 1 1 34910
0 34912 7 1 2 34906 34911
0 34913 7 1 2 34853 34912
0 34914 5 1 1 34913
0 34915 7 1 2 44494 34914
0 34916 5 1 1 34915
0 34917 7 1 2 56293 71056
0 34918 7 1 2 53830 34917
0 34919 7 1 2 64391 68394
0 34920 7 1 2 70195 34919
0 34921 7 1 2 34918 34920
0 34922 5 1 1 34921
0 34923 7 1 2 34916 34922
0 34924 5 1 1 34923
0 34925 7 1 2 66023 34924
0 34926 5 1 1 34925
0 34927 7 1 2 55640 57789
0 34928 5 1 1 34927
0 34929 7 1 2 43151 56964
0 34930 5 1 1 34929
0 34931 7 1 2 34928 34930
0 34932 5 1 1 34931
0 34933 7 1 2 69563 34932
0 34934 5 1 1 34933
0 34935 7 2 2 49410 66505
0 34936 5 1 1 71159
0 34937 7 1 2 43558 71160
0 34938 5 1 1 34937
0 34939 7 1 2 34934 34938
0 34940 5 1 1 34939
0 34941 7 1 2 42238 34940
0 34942 5 1 1 34941
0 34943 7 2 2 45774 61440
0 34944 7 1 2 55968 63252
0 34945 7 1 2 71161 34944
0 34946 5 1 1 34945
0 34947 7 1 2 34942 34946
0 34948 5 1 1 34947
0 34949 7 1 2 44260 71152
0 34950 7 1 2 34948 34949
0 34951 5 1 1 34950
0 34952 7 1 2 57493 68136
0 34953 5 1 1 34952
0 34954 7 1 2 47920 57661
0 34955 5 1 1 34954
0 34956 7 2 2 56582 34955
0 34957 7 1 2 49098 69564
0 34958 7 1 2 71163 34957
0 34959 5 1 1 34958
0 34960 7 1 2 34953 34959
0 34961 5 1 1 34960
0 34962 7 1 2 42239 34961
0 34963 5 1 1 34962
0 34964 7 1 2 56357 63344
0 34965 7 1 2 62856 34964
0 34966 5 1 1 34965
0 34967 7 1 2 34963 34966
0 34968 5 1 1 34967
0 34969 7 1 2 43152 71149
0 34970 7 1 2 34968 34969
0 34971 5 1 1 34970
0 34972 7 1 2 43377 34971
0 34973 7 1 2 34951 34972
0 34974 5 1 1 34973
0 34975 7 1 2 60071 67325
0 34976 5 1 1 34975
0 34977 7 2 2 43770 58419
0 34978 7 1 2 61113 71165
0 34979 5 1 1 34978
0 34980 7 1 2 46326 34979
0 34981 7 1 2 34976 34980
0 34982 5 1 1 34981
0 34983 7 1 2 42903 70610
0 34984 5 1 1 34983
0 34985 7 1 2 47921 71028
0 34986 7 1 2 34984 34985
0 34987 7 1 2 34982 34986
0 34988 5 1 1 34987
0 34989 7 1 2 71154 71166
0 34990 5 1 1 34989
0 34991 7 1 2 55318 71150
0 34992 5 1 1 34991
0 34993 7 1 2 34990 34992
0 34994 5 1 1 34993
0 34995 7 2 2 52793 66521
0 34996 7 1 2 34994 71167
0 34997 5 1 1 34996
0 34998 7 1 2 46756 34997
0 34999 7 1 2 34988 34998
0 35000 5 1 1 34999
0 35001 7 1 2 59211 35000
0 35002 7 1 2 34974 35001
0 35003 5 1 1 35002
0 35004 7 1 2 60830 63654
0 35005 7 1 2 70884 35004
0 35006 5 1 1 35005
0 35007 7 1 2 53314 66506
0 35008 7 1 2 60484 35007
0 35009 5 1 1 35008
0 35010 7 1 2 35006 35009
0 35011 5 1 1 35010
0 35012 7 1 2 46543 35011
0 35013 5 1 1 35012
0 35014 7 2 2 55279 66589
0 35015 5 1 1 71169
0 35016 7 1 2 70885 71170
0 35017 5 1 1 35016
0 35018 7 1 2 35013 35017
0 35019 5 1 1 35018
0 35020 7 1 2 60878 63093
0 35021 7 1 2 35019 35020
0 35022 5 1 1 35021
0 35023 7 1 2 35003 35022
0 35024 5 1 1 35023
0 35025 7 1 2 42076 35024
0 35026 5 1 1 35025
0 35027 7 1 2 62766 65440
0 35028 5 1 1 35027
0 35029 7 1 2 35015 35028
0 35030 5 1 1 35029
0 35031 7 1 2 59001 70894
0 35032 5 1 1 35031
0 35033 7 1 2 1912 10670
0 35034 5 1 1 35033
0 35035 7 1 2 42240 2646
0 35036 7 1 2 65792 35035
0 35037 7 1 2 35034 35036
0 35038 5 1 1 35037
0 35039 7 1 2 35032 35038
0 35040 5 1 1 35039
0 35041 7 1 2 35030 35040
0 35042 5 1 1 35041
0 35043 7 1 2 46861 71029
0 35044 5 1 1 35043
0 35045 7 1 2 28823 35044
0 35046 5 1 1 35045
0 35047 7 3 2 47922 49305
0 35048 7 1 2 51238 71171
0 35049 7 1 2 35046 35048
0 35050 5 1 1 35049
0 35051 7 1 2 35042 35050
0 35052 5 1 1 35051
0 35053 7 1 2 71158 35052
0 35054 5 1 1 35053
0 35055 7 1 2 35026 35054
0 35056 5 1 1 35055
0 35057 7 1 2 44495 35056
0 35058 5 1 1 35057
0 35059 7 3 2 45632 64308
0 35060 7 1 2 60082 71174
0 35061 5 1 1 35060
0 35062 7 2 2 54808 70110
0 35063 7 1 2 44362 56108
0 35064 7 1 2 71177 35063
0 35065 5 1 1 35064
0 35066 7 1 2 35061 35065
0 35067 5 1 1 35066
0 35068 7 1 2 47589 35067
0 35069 5 1 1 35068
0 35070 7 1 2 58203 61696
0 35071 7 1 2 69088 35070
0 35072 5 1 1 35071
0 35073 7 1 2 35069 35072
0 35074 5 1 1 35073
0 35075 7 1 2 46757 35074
0 35076 5 1 1 35075
0 35077 7 2 2 57275 59741
0 35078 7 1 2 66530 71175
0 35079 7 1 2 71179 35078
0 35080 5 1 1 35079
0 35081 7 1 2 35076 35080
0 35082 5 1 1 35081
0 35083 7 1 2 53614 35082
0 35084 5 1 1 35083
0 35085 7 1 2 51032 67172
0 35086 5 1 1 35085
0 35087 7 1 2 61697 70009
0 35088 5 1 1 35087
0 35089 7 1 2 35086 35088
0 35090 5 1 1 35089
0 35091 7 1 2 50791 66791
0 35092 7 1 2 35090 35091
0 35093 5 1 1 35092
0 35094 7 1 2 35084 35093
0 35095 5 1 1 35094
0 35096 7 1 2 53866 69433
0 35097 7 1 2 35095 35096
0 35098 5 1 1 35097
0 35099 7 1 2 35058 35098
0 35100 5 1 1 35099
0 35101 7 1 2 66282 35100
0 35102 5 1 1 35101
0 35103 7 1 2 57639 59982
0 35104 7 1 2 70139 35103
0 35105 7 1 2 71147 35104
0 35106 7 1 2 70193 35105
0 35107 7 1 2 69007 35106
0 35108 5 1 1 35107
0 35109 7 1 2 35102 35108
0 35110 7 1 2 34926 35109
0 35111 7 1 2 34802 35110
0 35112 7 1 2 33766 35111
0 35113 5 1 1 35112
0 35114 7 1 2 66776 35113
0 35115 5 1 1 35114
0 35116 7 1 2 33631 35115
0 35117 7 1 2 33063 35116
0 35118 7 1 2 31001 35117
0 35119 7 1 2 47145 65449
0 35120 5 1 1 35119
0 35121 7 1 2 50107 52461
0 35122 5 1 1 35121
0 35123 7 1 2 35120 35122
0 35124 5 1 1 35123
0 35125 7 1 2 42904 35124
0 35126 5 1 1 35125
0 35127 7 1 2 51033 52401
0 35128 5 1 1 35127
0 35129 7 2 2 48981 35128
0 35130 5 1 1 71181
0 35131 7 1 2 49355 71182
0 35132 5 1 1 35131
0 35133 7 1 2 50018 35132
0 35134 5 1 1 35133
0 35135 7 1 2 58561 35134
0 35136 5 2 1 35135
0 35137 7 1 2 46327 71183
0 35138 5 1 1 35137
0 35139 7 3 2 50565 63696
0 35140 5 1 1 71185
0 35141 7 1 2 35138 35140
0 35142 5 1 1 35141
0 35143 7 1 2 43771 35142
0 35144 5 1 1 35143
0 35145 7 1 2 35126 35144
0 35146 5 1 1 35145
0 35147 7 1 2 42620 35146
0 35148 5 1 1 35147
0 35149 7 1 2 55869 65450
0 35150 5 1 1 35149
0 35151 7 1 2 35148 35150
0 35152 5 1 1 35151
0 35153 7 1 2 70369 35152
0 35154 5 1 1 35153
0 35155 7 1 2 44115 60716
0 35156 5 1 1 35155
0 35157 7 1 2 67276 35156
0 35158 5 2 1 35157
0 35159 7 1 2 43378 71188
0 35160 5 1 1 35159
0 35161 7 1 2 44261 54019
0 35162 5 1 1 35161
0 35163 7 1 2 35160 35162
0 35164 5 4 1 35163
0 35165 7 2 2 62243 71190
0 35166 7 1 2 63816 71194
0 35167 5 1 1 35166
0 35168 7 1 2 35154 35167
0 35169 5 1 1 35168
0 35170 7 1 2 48299 35169
0 35171 5 1 1 35170
0 35172 7 2 2 48683 55287
0 35173 7 1 2 63817 71196
0 35174 7 1 2 71191 35173
0 35175 5 1 1 35174
0 35176 7 1 2 35171 35175
0 35177 5 1 1 35176
0 35178 7 1 2 54809 35177
0 35179 5 1 1 35178
0 35180 7 1 2 54020 59793
0 35181 5 1 1 35180
0 35182 7 1 2 53430 59862
0 35183 5 2 1 35182
0 35184 7 1 2 35181 71198
0 35185 5 1 1 35184
0 35186 7 1 2 44262 35185
0 35187 5 1 1 35186
0 35188 7 1 2 54021 61751
0 35189 5 2 1 35188
0 35190 7 1 2 35187 71200
0 35191 5 1 1 35190
0 35192 7 1 2 43379 35191
0 35193 5 1 1 35192
0 35194 7 1 2 59902 61453
0 35195 5 1 1 35194
0 35196 7 1 2 35193 35195
0 35197 5 1 1 35196
0 35198 7 1 2 48684 35197
0 35199 5 1 1 35198
0 35200 7 1 2 54317 59930
0 35201 7 1 2 70416 35200
0 35202 5 1 1 35201
0 35203 7 1 2 44972 35202
0 35204 7 1 2 35199 35203
0 35205 5 1 1 35204
0 35206 7 1 2 63928 66895
0 35207 5 1 1 35206
0 35208 7 2 2 42077 53044
0 35209 7 1 2 59212 71202
0 35210 5 2 1 35209
0 35211 7 1 2 35207 71204
0 35212 5 1 1 35211
0 35213 7 1 2 50108 35212
0 35214 5 1 1 35213
0 35215 7 1 2 49921 61454
0 35216 7 1 2 71180 35215
0 35217 5 1 1 35216
0 35218 7 1 2 11441 35217
0 35219 5 1 1 35218
0 35220 7 1 2 45310 35219
0 35221 5 1 1 35220
0 35222 7 1 2 48300 35221
0 35223 7 1 2 35214 35222
0 35224 5 1 1 35223
0 35225 7 1 2 42621 35224
0 35226 7 1 2 35205 35225
0 35227 5 1 1 35226
0 35228 7 1 2 64603 28962
0 35229 5 1 1 35228
0 35230 7 1 2 42905 35229
0 35231 5 1 1 35230
0 35232 7 1 2 57083 65585
0 35233 5 1 1 35232
0 35234 7 1 2 35231 35233
0 35235 5 1 1 35234
0 35236 7 1 2 50019 35235
0 35237 5 1 1 35236
0 35238 7 1 2 58592 65340
0 35239 5 2 1 35238
0 35240 7 1 2 35237 71206
0 35241 5 1 1 35240
0 35242 7 1 2 48914 69372
0 35243 7 1 2 35241 35242
0 35244 5 1 1 35243
0 35245 7 1 2 35227 35244
0 35246 5 1 1 35245
0 35247 7 1 2 43772 35246
0 35248 5 1 1 35247
0 35249 7 1 2 52566 70766
0 35250 7 1 2 60867 35249
0 35251 7 1 2 70188 35250
0 35252 5 1 1 35251
0 35253 7 1 2 35248 35252
0 35254 5 1 1 35253
0 35255 7 1 2 56908 35254
0 35256 5 1 1 35255
0 35257 7 1 2 35179 35256
0 35258 5 1 1 35257
0 35259 7 1 2 66024 35258
0 35260 5 1 1 35259
0 35261 7 3 2 48301 53291
0 35262 7 1 2 57640 66649
0 35263 5 1 1 35262
0 35264 7 1 2 58700 35263
0 35265 5 1 1 35264
0 35266 7 1 2 65749 35265
0 35267 5 2 1 35266
0 35268 7 1 2 55680 57641
0 35269 5 1 1 35268
0 35270 7 1 2 58701 35269
0 35271 5 1 1 35270
0 35272 7 1 2 70363 35271
0 35273 5 1 1 35272
0 35274 7 1 2 71211 35273
0 35275 5 1 1 35274
0 35276 7 1 2 44263 35275
0 35277 5 1 1 35276
0 35278 7 2 2 48947 56921
0 35279 7 1 2 71067 71213
0 35280 5 1 1 35279
0 35281 7 1 2 35277 35280
0 35282 5 1 1 35281
0 35283 7 1 2 44116 59484
0 35284 7 1 2 35282 35283
0 35285 5 1 1 35284
0 35286 7 1 2 49356 63824
0 35287 7 1 2 66965 35286
0 35288 5 1 1 35287
0 35289 7 1 2 35285 35288
0 35290 5 1 1 35289
0 35291 7 1 2 45633 35290
0 35292 5 1 1 35291
0 35293 7 1 2 68543 70900
0 35294 5 1 1 35293
0 35295 7 2 2 45866 69855
0 35296 5 1 1 71215
0 35297 7 1 2 57515 71216
0 35298 5 1 1 35297
0 35299 7 1 2 35294 35298
0 35300 5 1 1 35299
0 35301 7 1 2 59402 35300
0 35302 5 1 1 35301
0 35303 7 1 2 35292 35302
0 35304 5 1 1 35303
0 35305 7 1 2 48846 35304
0 35306 5 1 1 35305
0 35307 7 2 2 55853 56994
0 35308 5 1 1 71217
0 35309 7 1 2 65956 71218
0 35310 5 1 1 35309
0 35311 7 1 2 71212 35310
0 35312 5 1 1 35311
0 35313 7 1 2 68466 35312
0 35314 5 1 1 35313
0 35315 7 2 2 58068 64693
0 35316 7 1 2 56922 70181
0 35317 7 1 2 71219 35316
0 35318 5 1 1 35317
0 35319 7 1 2 35314 35318
0 35320 5 1 1 35319
0 35321 7 1 2 58450 35320
0 35322 5 1 1 35321
0 35323 7 1 2 58843 58284
0 35324 7 1 2 60234 35323
0 35325 5 1 1 35324
0 35326 7 1 2 59934 35325
0 35327 5 1 1 35326
0 35328 7 1 2 43153 35327
0 35329 5 1 1 35328
0 35330 7 1 2 44117 66851
0 35331 5 1 1 35330
0 35332 7 1 2 35329 35331
0 35333 5 1 1 35332
0 35334 7 1 2 45867 71214
0 35335 7 1 2 35333 35334
0 35336 5 1 1 35335
0 35337 7 1 2 35322 35336
0 35338 7 1 2 35306 35337
0 35339 5 1 1 35338
0 35340 7 1 2 48685 35339
0 35341 5 1 1 35340
0 35342 7 1 2 30092 35308
0 35343 5 1 1 35342
0 35344 7 1 2 43154 35343
0 35345 5 1 1 35344
0 35346 7 1 2 56909 62368
0 35347 5 1 1 35346
0 35348 7 1 2 35345 35347
0 35349 5 1 1 35348
0 35350 7 1 2 59794 35349
0 35351 5 1 1 35350
0 35352 7 1 2 56928 59771
0 35353 5 1 1 35352
0 35354 7 1 2 35351 35353
0 35355 5 1 1 35354
0 35356 7 1 2 48686 35355
0 35357 5 1 1 35356
0 35358 7 1 2 58698 59886
0 35359 7 1 2 59873 35358
0 35360 5 1 1 35359
0 35361 7 1 2 35357 35360
0 35362 5 1 1 35361
0 35363 7 1 2 65750 35362
0 35364 5 1 1 35363
0 35365 7 2 2 50960 63789
0 35366 7 1 2 56564 70599
0 35367 7 1 2 71221 35366
0 35368 5 1 1 35367
0 35369 7 1 2 35364 35368
0 35370 5 1 1 35369
0 35371 7 1 2 49241 35370
0 35372 5 1 1 35371
0 35373 7 2 2 54810 69856
0 35374 7 1 2 60185 68420
0 35375 7 1 2 71223 35374
0 35376 5 1 1 35375
0 35377 7 2 2 57616 58270
0 35378 7 1 2 45634 64433
0 35379 7 1 2 64718 35378
0 35380 7 1 2 71225 35379
0 35381 5 1 1 35380
0 35382 7 1 2 35376 35381
0 35383 5 1 1 35382
0 35384 7 1 2 66450 35383
0 35385 5 1 1 35384
0 35386 7 2 2 63026 66706
0 35387 7 1 2 71222 71227
0 35388 5 1 1 35387
0 35389 7 1 2 35385 35388
0 35390 5 1 1 35389
0 35391 7 1 2 49057 35390
0 35392 5 1 1 35391
0 35393 7 1 2 35372 35392
0 35394 7 1 2 35341 35393
0 35395 5 1 1 35394
0 35396 7 1 2 42906 35395
0 35397 5 1 1 35396
0 35398 7 1 2 70408 70374
0 35399 5 1 1 35398
0 35400 7 1 2 56358 64051
0 35401 7 1 2 58706 35400
0 35402 5 1 1 35401
0 35403 7 1 2 35399 35402
0 35404 5 1 1 35403
0 35405 7 1 2 59921 65586
0 35406 7 1 2 35404 35405
0 35407 5 1 1 35406
0 35408 7 1 2 35397 35407
0 35409 5 1 1 35408
0 35410 7 1 2 71208 35409
0 35411 5 1 1 35410
0 35412 7 1 2 43155 64144
0 35413 5 1 1 35412
0 35414 7 1 2 60875 35413
0 35415 5 1 1 35414
0 35416 7 1 2 59795 35415
0 35417 5 1 1 35416
0 35418 7 1 2 59926 35417
0 35419 5 1 1 35418
0 35420 7 1 2 46328 35419
0 35421 5 1 1 35420
0 35422 7 1 2 59863 65359
0 35423 5 1 1 35422
0 35424 7 1 2 35421 35423
0 35425 5 1 1 35424
0 35426 7 1 2 45311 35425
0 35427 5 1 1 35426
0 35428 7 1 2 50792 63904
0 35429 5 1 1 35428
0 35430 7 1 2 46862 61455
0 35431 7 2 2 70140 35430
0 35432 5 1 1 71229
0 35433 7 2 2 46544 71230
0 35434 5 1 1 71231
0 35435 7 1 2 71205 35434
0 35436 5 1 1 35435
0 35437 7 1 2 57992 35436
0 35438 5 1 1 35437
0 35439 7 1 2 35429 35438
0 35440 7 1 2 35427 35439
0 35441 5 1 1 35440
0 35442 7 1 2 65751 35441
0 35443 5 1 1 35442
0 35444 7 1 2 62356 68576
0 35445 5 1 1 35444
0 35446 7 1 2 59935 35445
0 35447 5 1 1 35446
0 35448 7 1 2 47456 35447
0 35449 5 1 1 35448
0 35450 7 1 2 60203 60219
0 35451 7 1 2 61840 35450
0 35452 5 2 1 35451
0 35453 7 1 2 59922 71233
0 35454 5 1 1 35453
0 35455 7 1 2 35449 35454
0 35456 5 1 1 35455
0 35457 7 1 2 46329 35456
0 35458 5 1 1 35457
0 35459 7 2 2 50566 59923
0 35460 7 1 2 57813 26198
0 35461 7 1 2 71235 35460
0 35462 5 1 1 35461
0 35463 7 1 2 35458 35462
0 35464 5 1 1 35463
0 35465 7 1 2 65957 35464
0 35466 5 1 1 35465
0 35467 7 1 2 35443 35466
0 35468 5 1 1 35467
0 35469 7 1 2 57424 35468
0 35470 5 1 1 35469
0 35471 7 1 2 54989 66948
0 35472 5 1 1 35471
0 35473 7 1 2 56124 60006
0 35474 7 1 2 60027 35473
0 35475 5 1 1 35474
0 35476 7 1 2 35472 35475
0 35477 5 1 1 35476
0 35478 7 1 2 50567 35477
0 35479 5 1 1 35478
0 35480 7 1 2 44118 70382
0 35481 5 1 1 35480
0 35482 7 1 2 70860 35481
0 35483 5 1 1 35482
0 35484 7 1 2 46330 35483
0 35485 5 1 1 35484
0 35486 7 1 2 35479 35485
0 35487 5 1 1 35486
0 35488 7 1 2 50793 35487
0 35489 5 1 1 35488
0 35490 7 1 2 64940 66949
0 35491 5 1 1 35490
0 35492 7 1 2 57620 70177
0 35493 5 1 1 35492
0 35494 7 1 2 35491 35493
0 35495 5 1 1 35494
0 35496 7 1 2 43380 35495
0 35497 5 1 1 35496
0 35498 7 1 2 35489 35497
0 35499 5 1 1 35498
0 35500 7 1 2 45635 35499
0 35501 5 1 1 35500
0 35502 7 2 2 43381 64941
0 35503 5 1 1 71237
0 35504 7 1 2 50794 62179
0 35505 5 1 1 35504
0 35506 7 1 2 35503 35505
0 35507 5 3 1 35506
0 35508 7 1 2 47923 54745
0 35509 7 1 2 59524 35508
0 35510 7 1 2 71239 35509
0 35511 5 1 1 35510
0 35512 7 1 2 35501 35511
0 35513 5 1 1 35512
0 35514 7 1 2 65810 35513
0 35515 5 1 1 35514
0 35516 7 1 2 50568 17027
0 35517 5 1 1 35516
0 35518 7 1 2 17023 70357
0 35519 5 1 1 35518
0 35520 7 1 2 57562 35519
0 35521 5 1 1 35520
0 35522 7 1 2 52078 70364
0 35523 5 1 1 35522
0 35524 7 1 2 35521 35523
0 35525 5 1 1 35524
0 35526 7 1 2 46331 35525
0 35527 5 1 1 35526
0 35528 7 1 2 35517 35527
0 35529 5 1 1 35528
0 35530 7 1 2 55012 59525
0 35531 7 1 2 35529 35530
0 35532 5 1 1 35531
0 35533 7 1 2 35515 35532
0 35534 7 1 2 35470 35533
0 35535 5 1 1 35534
0 35536 7 1 2 47813 35535
0 35537 5 1 1 35536
0 35538 7 1 2 59722 65603
0 35539 5 1 1 35538
0 35540 7 1 2 56910 64434
0 35541 7 1 2 70432 35540
0 35542 7 1 2 35539 35541
0 35543 5 1 1 35542
0 35544 7 1 2 48302 35543
0 35545 7 1 2 35537 35544
0 35546 5 1 1 35545
0 35547 7 1 2 55809 63027
0 35548 7 2 2 44599 57946
0 35549 7 1 2 70438 71242
0 35550 7 1 2 35547 35549
0 35551 5 1 1 35550
0 35552 7 2 2 58271 59427
0 35553 5 1 1 71244
0 35554 7 1 2 43156 71245
0 35555 5 1 1 35554
0 35556 7 1 2 49357 59526
0 35557 7 1 2 63843 35556
0 35558 5 1 1 35557
0 35559 7 1 2 35555 35558
0 35560 5 1 1 35559
0 35561 7 1 2 54811 65958
0 35562 7 1 2 35560 35561
0 35563 5 1 1 35562
0 35564 7 1 2 35551 35563
0 35565 5 1 1 35564
0 35566 7 1 2 56753 35565
0 35567 5 1 1 35566
0 35568 7 1 2 60651 71087
0 35569 5 1 1 35568
0 35570 7 1 2 45868 59167
0 35571 7 1 2 71224 35570
0 35572 5 1 1 35571
0 35573 7 1 2 35569 35572
0 35574 5 1 1 35573
0 35575 7 1 2 51772 35574
0 35576 5 1 1 35575
0 35577 7 1 2 50873 65752
0 35578 5 3 1 35577
0 35579 7 1 2 45869 70081
0 35580 5 1 1 35579
0 35581 7 1 2 71246 35580
0 35582 5 1 1 35581
0 35583 7 1 2 43157 35582
0 35584 5 2 1 35583
0 35585 7 2 2 49457 70365
0 35586 5 1 1 71251
0 35587 7 1 2 71249 35586
0 35588 5 1 1 35587
0 35589 7 1 2 44119 59796
0 35590 7 1 2 35588 35589
0 35591 5 1 1 35590
0 35592 7 1 2 66902 67943
0 35593 5 1 1 35592
0 35594 7 1 2 45636 66974
0 35595 7 1 2 68077 35594
0 35596 5 1 1 35595
0 35597 7 1 2 35593 35596
0 35598 5 1 1 35597
0 35599 7 1 2 49358 35598
0 35600 5 1 1 35599
0 35601 7 2 2 59468 66636
0 35602 7 1 2 71220 71253
0 35603 5 1 1 35602
0 35604 7 1 2 35600 35603
0 35605 7 1 2 35591 35604
0 35606 5 1 1 35605
0 35607 7 1 2 47814 35606
0 35608 5 1 1 35607
0 35609 7 1 2 35576 35608
0 35610 5 1 1 35609
0 35611 7 1 2 46943 60261
0 35612 7 1 2 35610 35611
0 35613 5 1 1 35612
0 35614 7 1 2 35567 35613
0 35615 5 1 1 35614
0 35616 7 1 2 42907 35615
0 35617 5 1 1 35616
0 35618 7 1 2 49058 70366
0 35619 5 1 1 35618
0 35620 7 1 2 68490 35619
0 35621 5 1 1 35620
0 35622 7 2 2 48687 35621
0 35623 7 1 2 56135 57876
0 35624 7 1 2 60936 35623
0 35625 7 1 2 71255 35624
0 35626 5 1 1 35625
0 35627 7 1 2 44973 35626
0 35628 7 1 2 35617 35627
0 35629 5 1 1 35628
0 35630 7 1 2 51153 35629
0 35631 7 1 2 35546 35630
0 35632 5 1 1 35631
0 35633 7 1 2 35411 35632
0 35634 7 1 2 35260 35633
0 35635 5 1 1 35634
0 35636 7 1 2 70331 35635
0 35637 5 1 1 35636
0 35638 7 3 2 53633 57642
0 35639 5 1 1 71257
0 35640 7 2 2 53656 56430
0 35641 5 2 1 71260
0 35642 7 1 2 35639 71262
0 35643 5 1 1 35642
0 35644 7 1 2 65753 35643
0 35645 5 1 1 35644
0 35646 7 1 2 56583 60584
0 35647 5 1 1 35646
0 35648 7 1 2 71263 35647
0 35649 5 1 1 35648
0 35650 7 1 2 65959 35649
0 35651 5 1 1 35650
0 35652 7 1 2 35645 35651
0 35653 5 1 1 35652
0 35654 7 1 2 70245 35653
0 35655 5 1 1 35654
0 35656 7 1 2 56584 66086
0 35657 5 1 1 35656
0 35658 7 1 2 32981 35657
0 35659 5 1 1 35658
0 35660 7 2 2 47815 35659
0 35661 7 1 2 66178 71264
0 35662 5 1 1 35661
0 35663 7 1 2 35655 35662
0 35664 5 1 1 35663
0 35665 7 1 2 42078 35664
0 35666 5 1 1 35665
0 35667 7 2 2 65209 66360
0 35668 7 1 2 71265 71266
0 35669 5 1 1 35668
0 35670 7 1 2 35666 35669
0 35671 5 1 1 35670
0 35672 7 1 2 44120 35671
0 35673 5 1 1 35672
0 35674 7 1 2 62525 67086
0 35675 7 2 2 63742 66072
0 35676 7 1 2 69992 71268
0 35677 7 1 2 35674 35676
0 35678 5 1 1 35677
0 35679 7 1 2 35673 35678
0 35680 5 1 1 35679
0 35681 7 1 2 43382 35680
0 35682 5 1 1 35681
0 35683 7 1 2 48847 55829
0 35684 7 1 2 70977 35683
0 35685 7 1 2 70273 35684
0 35686 5 1 1 35685
0 35687 7 1 2 35682 35686
0 35688 5 1 1 35687
0 35689 7 1 2 43158 35688
0 35690 5 1 1 35689
0 35691 7 1 2 59242 66475
0 35692 7 2 2 70914 35691
0 35693 7 2 2 44121 48948
0 35694 7 1 2 56192 66073
0 35695 7 1 2 71272 35694
0 35696 7 1 2 71270 35695
0 35697 5 1 1 35696
0 35698 7 1 2 35690 35697
0 35699 5 1 1 35698
0 35700 7 1 2 59613 35699
0 35701 5 1 1 35700
0 35702 7 1 2 49520 61002
0 35703 7 2 2 66230 35702
0 35704 5 1 1 71274
0 35705 7 1 2 42079 66172
0 35706 5 1 1 35705
0 35707 7 1 2 18303 35706
0 35708 5 2 1 35707
0 35709 7 1 2 60665 8729
0 35710 5 1 1 35709
0 35711 7 1 2 71276 35710
0 35712 5 1 1 35711
0 35713 7 1 2 61331 70246
0 35714 5 1 1 35713
0 35715 7 2 2 45637 56193
0 35716 7 1 2 47691 71278
0 35717 7 1 2 66179 35716
0 35718 5 1 1 35717
0 35719 7 1 2 35714 35718
0 35720 7 1 2 35712 35719
0 35721 5 1 1 35720
0 35722 7 2 2 49359 35721
0 35723 7 1 2 48688 71280
0 35724 5 1 1 35723
0 35725 7 1 2 35704 35724
0 35726 5 1 1 35725
0 35727 7 1 2 43383 35726
0 35728 5 1 1 35727
0 35729 7 1 2 44264 71275
0 35730 5 1 1 35729
0 35731 7 1 2 47816 25289
0 35732 7 1 2 70280 35731
0 35733 5 1 1 35732
0 35734 7 1 2 59168 59898
0 35735 7 1 2 66231 35734
0 35736 5 1 1 35735
0 35737 7 1 2 35733 35736
0 35738 5 1 1 35737
0 35739 7 1 2 48689 35738
0 35740 5 1 1 35739
0 35741 7 1 2 35730 35740
0 35742 7 1 2 35728 35741
0 35743 5 1 1 35742
0 35744 7 1 2 51671 35743
0 35745 5 1 1 35744
0 35746 7 1 2 51601 70240
0 35747 5 1 1 35746
0 35748 7 2 2 49360 51672
0 35749 5 1 1 71282
0 35750 7 1 2 3344 35749
0 35751 5 2 1 35750
0 35752 7 1 2 47817 66205
0 35753 7 1 2 71284 35752
0 35754 5 1 1 35753
0 35755 7 1 2 35747 35754
0 35756 5 1 1 35755
0 35757 7 1 2 48848 35756
0 35758 5 1 1 35757
0 35759 7 1 2 46944 56565
0 35760 7 1 2 70241 35759
0 35761 5 1 1 35760
0 35762 7 1 2 35758 35761
0 35763 5 1 1 35762
0 35764 7 1 2 42080 35763
0 35765 5 1 1 35764
0 35766 7 1 2 60418 71267
0 35767 7 1 2 71285 35766
0 35768 5 1 1 35767
0 35769 7 1 2 35765 35768
0 35770 5 1 1 35769
0 35771 7 1 2 44363 35770
0 35772 5 1 1 35771
0 35773 7 1 2 51673 59169
0 35774 7 1 2 52105 35773
0 35775 7 1 2 66232 35774
0 35776 5 1 1 35775
0 35777 7 1 2 35772 35776
0 35778 5 1 1 35777
0 35779 7 1 2 50020 35778
0 35780 5 1 1 35779
0 35781 7 1 2 35745 35780
0 35782 5 1 1 35781
0 35783 7 1 2 65960 35782
0 35784 5 1 1 35783
0 35785 7 1 2 57503 57797
0 35786 7 1 2 71277 35785
0 35787 5 1 1 35786
0 35788 7 1 2 48690 71258
0 35789 5 1 1 35788
0 35790 7 1 2 48849 71261
0 35791 5 1 1 35790
0 35792 7 1 2 35789 35791
0 35793 5 1 1 35792
0 35794 7 1 2 45920 70196
0 35795 7 1 2 35793 35794
0 35796 5 1 1 35795
0 35797 7 1 2 35787 35796
0 35798 5 1 1 35797
0 35799 7 1 2 50874 35798
0 35800 5 1 1 35799
0 35801 7 1 2 4329 57793
0 35802 5 1 1 35801
0 35803 7 1 2 43384 35802
0 35804 5 1 1 35803
0 35805 7 1 2 51602 52393
0 35806 5 1 1 35805
0 35807 7 1 2 35804 35806
0 35808 5 1 1 35807
0 35809 7 1 2 60461 66222
0 35810 7 1 2 35808 35809
0 35811 5 1 1 35810
0 35812 7 1 2 35800 35811
0 35813 5 1 1 35812
0 35814 7 1 2 44122 35813
0 35815 5 1 1 35814
0 35816 7 1 2 48691 60861
0 35817 7 2 2 68220 35816
0 35818 7 1 2 58285 62679
0 35819 7 1 2 67306 35818
0 35820 7 1 2 71286 35819
0 35821 5 1 1 35820
0 35822 7 1 2 35815 35821
0 35823 5 1 1 35822
0 35824 7 1 2 43159 35823
0 35825 5 1 1 35824
0 35826 7 1 2 69038 70430
0 35827 7 1 2 71287 35826
0 35828 5 1 1 35827
0 35829 7 1 2 35825 35828
0 35830 5 1 1 35829
0 35831 7 1 2 47692 35830
0 35832 5 1 1 35831
0 35833 7 1 2 53688 56995
0 35834 7 1 2 62526 62670
0 35835 7 1 2 66388 35834
0 35836 7 1 2 35833 35835
0 35837 5 1 1 35836
0 35838 7 1 2 43559 57643
0 35839 7 1 2 60751 35838
0 35840 7 1 2 70274 35839
0 35841 5 1 1 35840
0 35842 7 1 2 35837 35841
0 35843 5 1 1 35842
0 35844 7 1 2 59614 35843
0 35845 5 1 1 35844
0 35846 7 1 2 35832 35845
0 35847 5 1 1 35846
0 35848 7 1 2 65754 35847
0 35849 5 1 1 35848
0 35850 7 4 2 51892 66407
0 35851 5 1 1 71288
0 35852 7 2 2 50367 65622
0 35853 5 1 1 71292
0 35854 7 1 2 35851 35853
0 35855 5 2 1 35854
0 35856 7 1 2 50875 71281
0 35857 5 1 1 35856
0 35858 7 1 2 50132 70225
0 35859 5 1 1 35858
0 35860 7 1 2 66686 69629
0 35861 7 1 2 62358 35860
0 35862 5 1 1 35861
0 35863 7 1 2 35859 35862
0 35864 5 1 1 35863
0 35865 7 1 2 44123 35864
0 35866 5 1 1 35865
0 35867 7 1 2 63496 70226
0 35868 5 1 1 35867
0 35869 7 1 2 35866 35868
0 35870 5 1 1 35869
0 35871 7 1 2 45638 35870
0 35872 5 1 1 35871
0 35873 7 1 2 60820 70235
0 35874 5 1 1 35873
0 35875 7 1 2 35872 35874
0 35876 5 1 1 35875
0 35877 7 1 2 47693 35876
0 35878 5 1 1 35877
0 35879 7 1 2 35857 35878
0 35880 5 1 1 35879
0 35881 7 1 2 48692 35880
0 35882 5 1 1 35881
0 35883 7 1 2 66233 69720
0 35884 5 1 1 35883
0 35885 7 1 2 35882 35884
0 35886 5 1 1 35885
0 35887 7 1 2 71294 35886
0 35888 5 1 1 35887
0 35889 7 1 2 35849 35888
0 35890 7 1 2 35784 35889
0 35891 5 1 1 35890
0 35892 7 1 2 42908 35891
0 35893 5 1 1 35892
0 35894 7 1 2 35701 35893
0 35895 5 1 1 35894
0 35896 7 1 2 55288 35895
0 35897 5 1 1 35896
0 35898 7 1 2 44690 53689
0 35899 7 1 2 63282 35898
0 35900 7 4 2 69266 35899
0 35901 5 1 1 71296
0 35902 7 1 2 48850 53431
0 35903 7 1 2 71297 35902
0 35904 5 1 1 35903
0 35905 7 2 2 63085 66173
0 35906 7 1 2 65636 69114
0 35907 7 1 2 71300 35906
0 35908 5 1 1 35907
0 35909 7 1 2 35904 35908
0 35910 5 2 1 35909
0 35911 7 1 2 64600 71302
0 35912 5 1 1 35911
0 35913 7 1 2 64606 67538
0 35914 7 1 2 70060 35913
0 35915 7 1 2 49411 61099
0 35916 7 1 2 68088 35915
0 35917 7 1 2 35914 35916
0 35918 5 1 1 35917
0 35919 7 1 2 35912 35918
0 35920 5 1 1 35919
0 35921 7 1 2 43385 35920
0 35922 5 1 1 35921
0 35923 7 1 2 42622 60909
0 35924 7 1 2 71298 35923
0 35925 5 1 1 35924
0 35926 7 1 2 35922 35925
0 35927 5 1 1 35926
0 35928 7 1 2 60462 35927
0 35929 5 1 1 35928
0 35930 7 1 2 70503 71155
0 35931 5 1 1 35930
0 35932 7 2 2 45921 60799
0 35933 7 2 2 52394 67132
0 35934 7 1 2 71304 71306
0 35935 5 1 1 35934
0 35936 7 1 2 35931 35935
0 35937 5 1 1 35936
0 35938 7 1 2 43386 35937
0 35939 5 1 1 35938
0 35940 7 1 2 49716 67133
0 35941 7 1 2 71305 35940
0 35942 5 1 1 35941
0 35943 7 1 2 35939 35942
0 35944 5 1 1 35943
0 35945 7 1 2 43160 35944
0 35946 5 1 1 35945
0 35947 7 1 2 44124 58286
0 35948 7 1 2 60796 66717
0 35949 7 1 2 35947 35948
0 35950 7 1 2 71307 35949
0 35951 5 1 1 35950
0 35952 7 1 2 35946 35951
0 35953 5 1 1 35952
0 35954 7 1 2 70781 35953
0 35955 5 1 1 35954
0 35956 7 1 2 35929 35955
0 35957 5 1 1 35956
0 35958 7 1 2 43773 35957
0 35959 5 1 1 35958
0 35960 7 1 2 56032 57947
0 35961 7 1 2 67180 68083
0 35962 7 1 2 35960 35961
0 35963 5 1 1 35962
0 35964 7 1 2 50961 63707
0 35965 5 1 1 35964
0 35966 7 1 2 55475 62527
0 35967 5 1 1 35966
0 35968 7 1 2 35965 35967
0 35969 5 1 1 35968
0 35970 7 1 2 67793 70311
0 35971 7 1 2 35969 35970
0 35972 5 1 1 35971
0 35973 7 1 2 35963 35972
0 35974 5 1 1 35973
0 35975 7 1 2 42909 35974
0 35976 5 1 1 35975
0 35977 7 1 2 44691 55830
0 35978 7 1 2 66672 35977
0 35979 7 1 2 67114 70539
0 35980 7 1 2 35978 35979
0 35981 5 1 1 35980
0 35982 7 1 2 35976 35981
0 35983 5 1 1 35982
0 35984 7 1 2 43387 35983
0 35985 5 1 1 35984
0 35986 7 1 2 59887 67105
0 35987 7 1 2 70314 35986
0 35988 5 1 1 35987
0 35989 7 1 2 35985 35988
0 35990 5 1 1 35989
0 35991 7 1 2 48693 53203
0 35992 7 1 2 35990 35991
0 35993 5 1 1 35992
0 35994 7 1 2 35959 35993
0 35995 5 1 1 35994
0 35996 7 1 2 48303 35995
0 35997 5 1 1 35996
0 35998 7 2 2 53432 54568
0 35999 7 1 2 70578 71308
0 36000 5 1 1 35999
0 36001 7 2 2 60496 63122
0 36002 7 2 2 67829 71310
0 36003 7 1 2 54178 71312
0 36004 5 1 1 36003
0 36005 7 1 2 36000 36004
0 36006 5 1 1 36005
0 36007 7 1 2 53341 36006
0 36008 5 1 1 36007
0 36009 7 1 2 61867 71313
0 36010 5 1 1 36009
0 36011 7 1 2 36008 36010
0 36012 5 1 1 36011
0 36013 7 1 2 48694 36012
0 36014 5 1 1 36013
0 36015 7 1 2 63404 68275
0 36016 7 1 2 61617 36015
0 36017 7 1 2 60910 36016
0 36018 5 1 1 36017
0 36019 7 1 2 36014 36018
0 36020 5 1 1 36019
0 36021 7 1 2 66206 36020
0 36022 5 1 1 36021
0 36023 7 1 2 60510 71197
0 36024 7 1 2 71303 36023
0 36025 5 1 1 36024
0 36026 7 1 2 36022 36025
0 36027 7 1 2 35997 36026
0 36028 5 1 1 36027
0 36029 7 1 2 51631 34722
0 36030 5 1 1 36029
0 36031 7 1 2 36028 36030
0 36032 5 1 1 36031
0 36033 7 3 2 48695 51674
0 36034 5 1 1 71314
0 36035 7 1 2 63377 71315
0 36036 5 1 1 36035
0 36037 7 1 2 46332 51603
0 36038 7 1 2 59640 36037
0 36039 5 1 1 36038
0 36040 7 1 2 36036 36039
0 36041 5 1 1 36040
0 36042 7 1 2 62528 36041
0 36043 5 1 1 36042
0 36044 7 1 2 45639 54659
0 36045 7 1 2 70133 36044
0 36046 5 1 1 36045
0 36047 7 1 2 36043 36046
0 36048 5 1 1 36047
0 36049 7 1 2 43388 36048
0 36050 5 1 1 36049
0 36051 7 2 2 57790 70129
0 36052 5 2 1 71317
0 36053 7 1 2 3362 71319
0 36054 5 1 1 36053
0 36055 7 3 2 48696 60463
0 36056 7 1 2 47146 71321
0 36057 7 1 2 36054 36056
0 36058 5 1 1 36057
0 36059 7 1 2 36050 36058
0 36060 5 1 1 36059
0 36061 7 1 2 44265 36060
0 36062 5 1 1 36061
0 36063 7 1 2 42910 52198
0 36064 5 1 1 36063
0 36065 7 1 2 53732 60048
0 36066 7 1 2 63787 36065
0 36067 7 1 2 36064 36066
0 36068 5 1 1 36067
0 36069 7 1 2 36062 36068
0 36070 5 1 1 36069
0 36071 7 1 2 43161 36070
0 36072 5 1 1 36071
0 36073 7 1 2 61456 66650
0 36074 7 1 2 64042 36073
0 36075 7 1 2 70631 36074
0 36076 5 1 1 36075
0 36077 7 3 2 56431 58120
0 36078 5 2 1 71324
0 36079 7 1 2 53693 57644
0 36080 5 1 1 36079
0 36081 7 1 2 71327 36080
0 36082 5 2 1 36081
0 36083 7 1 2 43389 71329
0 36084 5 1 1 36083
0 36085 7 1 2 43560 57791
0 36086 5 3 1 36085
0 36087 7 1 2 16814 71331
0 36088 5 2 1 36087
0 36089 7 1 2 60464 71334
0 36090 5 1 1 36089
0 36091 7 1 2 36084 36090
0 36092 5 1 1 36091
0 36093 7 1 2 50297 56730
0 36094 7 1 2 36092 36093
0 36095 5 1 1 36094
0 36096 7 1 2 36076 36095
0 36097 7 1 2 36072 36096
0 36098 5 1 1 36097
0 36099 7 1 2 42623 36098
0 36100 5 1 1 36099
0 36101 7 2 2 51034 60465
0 36102 5 1 1 71336
0 36103 7 1 2 62551 36102
0 36104 5 1 1 36103
0 36105 7 1 2 42624 36104
0 36106 5 1 1 36105
0 36107 7 1 2 56180 70985
0 36108 5 1 1 36107
0 36109 7 1 2 36106 36108
0 36110 5 1 1 36109
0 36111 7 1 2 51604 36110
0 36112 5 1 1 36111
0 36113 7 3 2 47818 59990
0 36114 7 1 2 53959 56978
0 36115 7 1 2 71338 36114
0 36116 5 1 1 36115
0 36117 7 1 2 36112 36116
0 36118 5 1 1 36117
0 36119 7 1 2 47590 36118
0 36120 5 1 1 36119
0 36121 7 1 2 48851 71328
0 36122 5 1 1 36121
0 36123 7 3 2 71330 36122
0 36124 7 1 2 69541 71341
0 36125 5 1 1 36124
0 36126 7 1 2 36120 36125
0 36127 5 1 1 36126
0 36128 7 1 2 46758 36127
0 36129 5 1 1 36128
0 36130 7 1 2 51035 58987
0 36131 7 1 2 61585 36130
0 36132 5 1 1 36131
0 36133 7 1 2 10673 36132
0 36134 5 1 1 36133
0 36135 7 1 2 51605 36134
0 36136 5 1 1 36135
0 36137 7 1 2 54038 60511
0 36138 5 1 1 36137
0 36139 7 2 2 42081 57963
0 36140 7 1 2 51036 71344
0 36141 5 1 1 36140
0 36142 7 2 2 54039 62529
0 36143 5 1 1 71346
0 36144 7 1 2 36141 36143
0 36145 7 1 2 36138 36144
0 36146 5 1 1 36145
0 36147 7 1 2 51675 36146
0 36148 5 1 1 36147
0 36149 7 1 2 36136 36148
0 36150 5 1 1 36149
0 36151 7 1 2 42625 36150
0 36152 5 1 1 36151
0 36153 7 1 2 36129 36152
0 36154 5 1 1 36153
0 36155 7 1 2 45312 36154
0 36156 5 1 1 36155
0 36157 7 1 2 56902 61842
0 36158 5 1 1 36157
0 36159 7 1 2 51676 36158
0 36160 5 1 1 36159
0 36161 7 1 2 51531 51606
0 36162 5 1 1 36161
0 36163 7 1 2 36160 36162
0 36164 5 1 1 36163
0 36165 7 1 2 60466 36164
0 36166 5 1 1 36165
0 36167 7 1 2 56585 62530
0 36168 7 1 2 5561 36167
0 36169 5 1 1 36168
0 36170 7 1 2 36166 36169
0 36171 5 1 1 36170
0 36172 7 1 2 42626 36171
0 36173 5 1 1 36172
0 36174 7 2 2 51357 62531
0 36175 7 1 2 71318 71348
0 36176 5 1 1 36175
0 36177 7 1 2 36173 36176
0 36178 5 1 1 36177
0 36179 7 1 2 46333 36178
0 36180 5 1 1 36179
0 36181 7 1 2 50876 71283
0 36182 5 1 1 36181
0 36183 7 3 2 43561 64239
0 36184 5 1 1 71350
0 36185 7 1 2 60752 71351
0 36186 5 1 1 36185
0 36187 7 1 2 36182 36186
0 36188 5 1 1 36187
0 36189 7 1 2 60467 36188
0 36190 5 1 1 36189
0 36191 7 1 2 50021 71325
0 36192 5 1 1 36191
0 36193 7 1 2 36190 36192
0 36194 5 1 1 36193
0 36195 7 1 2 46095 36194
0 36196 5 1 1 36195
0 36197 7 1 2 58665 62532
0 36198 7 1 2 56973 36197
0 36199 5 1 1 36198
0 36200 7 1 2 36196 36199
0 36201 5 1 1 36200
0 36202 7 1 2 42911 36201
0 36203 5 1 1 36202
0 36204 7 2 2 50795 60468
0 36205 7 1 2 53862 71353
0 36206 5 1 1 36205
0 36207 7 1 2 58628 71349
0 36208 5 1 1 36207
0 36209 7 1 2 36206 36208
0 36210 5 1 1 36209
0 36211 7 1 2 51677 36210
0 36212 5 1 1 36211
0 36213 7 1 2 64513 69955
0 36214 5 1 1 36213
0 36215 7 1 2 65201 67975
0 36216 5 1 1 36215
0 36217 7 1 2 36214 36216
0 36218 5 1 1 36217
0 36219 7 1 2 43162 51607
0 36220 7 1 2 36218 36219
0 36221 5 1 1 36220
0 36222 7 1 2 36212 36221
0 36223 7 1 2 36203 36222
0 36224 5 1 1 36223
0 36225 7 1 2 48697 36224
0 36226 5 1 1 36225
0 36227 7 1 2 50109 71342
0 36228 5 1 1 36227
0 36229 7 2 2 45640 68316
0 36230 7 1 2 70404 71355
0 36231 5 1 1 36230
0 36232 7 1 2 36228 36231
0 36233 5 1 1 36232
0 36234 7 1 2 46545 36233
0 36235 5 1 1 36234
0 36236 7 1 2 46759 60049
0 36237 7 1 2 64703 36236
0 36238 5 1 1 36237
0 36239 7 1 2 36235 36238
0 36240 5 1 1 36239
0 36241 7 1 2 64607 36240
0 36242 5 1 1 36241
0 36243 7 1 2 36226 36242
0 36244 7 1 2 36180 36243
0 36245 7 1 2 36156 36244
0 36246 5 1 1 36245
0 36247 7 1 2 43774 36246
0 36248 5 1 1 36247
0 36249 7 1 2 36100 36248
0 36250 5 1 1 36249
0 36251 7 1 2 70504 36250
0 36252 5 1 1 36251
0 36253 7 1 2 60857 68890
0 36254 5 1 1 36253
0 36255 7 1 2 54855 64212
0 36256 5 1 1 36255
0 36257 7 1 2 36254 36256
0 36258 5 1 1 36257
0 36259 7 1 2 42627 36258
0 36260 5 1 1 36259
0 36261 7 1 2 55870 64213
0 36262 5 1 1 36261
0 36263 7 1 2 36260 36262
0 36264 5 1 1 36263
0 36265 7 1 2 48852 36264
0 36266 5 1 1 36265
0 36267 7 1 2 52462 61351
0 36268 7 1 2 57993 36267
0 36269 5 1 1 36268
0 36270 7 1 2 36266 36269
0 36271 5 1 1 36270
0 36272 7 1 2 60469 36271
0 36273 5 1 1 36272
0 36274 7 1 2 44266 71238
0 36275 5 1 1 36274
0 36276 7 1 2 57545 36275
0 36277 5 1 1 36276
0 36278 7 1 2 45494 36277
0 36279 5 2 1 36278
0 36280 7 1 2 65463 71357
0 36281 5 2 1 36280
0 36282 7 1 2 70788 71359
0 36283 5 1 1 36282
0 36284 7 1 2 36273 36283
0 36285 5 1 1 36284
0 36286 7 1 2 51608 36285
0 36287 5 1 1 36286
0 36288 7 1 2 51609 60850
0 36289 7 1 2 71339 36288
0 36290 5 1 1 36289
0 36291 7 1 2 57798 62533
0 36292 5 1 1 36291
0 36293 7 1 2 51610 71322
0 36294 5 1 1 36293
0 36295 7 1 2 36292 36294
0 36296 5 1 1 36295
0 36297 7 1 2 44125 62088
0 36298 7 1 2 36296 36297
0 36299 5 1 1 36298
0 36300 7 1 2 36290 36299
0 36301 5 1 1 36300
0 36302 7 1 2 43163 36301
0 36303 5 1 1 36302
0 36304 7 1 2 51678 61827
0 36305 7 1 2 70789 36304
0 36306 7 1 2 51479 36305
0 36307 5 1 1 36306
0 36308 7 1 2 36303 36307
0 36309 5 1 1 36308
0 36310 7 1 2 50877 36309
0 36311 5 1 1 36310
0 36312 7 1 2 51735 62479
0 36313 5 1 1 36312
0 36314 7 1 2 60470 61385
0 36315 7 1 2 64547 36314
0 36316 5 1 1 36315
0 36317 7 1 2 36313 36316
0 36318 5 1 1 36317
0 36319 7 1 2 45313 36318
0 36320 5 1 1 36319
0 36321 7 1 2 51539 68222
0 36322 5 1 1 36321
0 36323 7 1 2 36320 36322
0 36324 5 1 1 36323
0 36325 7 1 2 46334 36324
0 36326 5 1 1 36325
0 36327 7 1 2 42082 61534
0 36328 7 1 2 63643 36327
0 36329 5 1 1 36328
0 36330 7 1 2 36326 36329
0 36331 5 1 1 36330
0 36332 7 1 2 52148 56294
0 36333 7 1 2 36331 36332
0 36334 5 1 1 36333
0 36335 7 1 2 36311 36334
0 36336 7 1 2 36287 36335
0 36337 5 1 1 36336
0 36338 7 1 2 70292 36337
0 36339 5 1 1 36338
0 36340 7 1 2 36252 36339
0 36341 5 1 1 36340
0 36342 7 1 2 65755 36341
0 36343 5 1 1 36342
0 36344 7 2 2 45495 57542
0 36345 7 1 2 50796 71361
0 36346 5 1 1 36345
0 36347 7 1 2 65464 36346
0 36348 5 1 1 36347
0 36349 7 1 2 51154 36348
0 36350 5 1 1 36349
0 36351 7 1 2 62089 64867
0 36352 5 2 1 36351
0 36353 7 1 2 52106 62090
0 36354 5 1 1 36353
0 36355 7 1 2 53034 62422
0 36356 7 2 2 59343 36355
0 36357 5 1 1 71365
0 36358 7 1 2 53721 59643
0 36359 5 1 1 36358
0 36360 7 1 2 43164 36359
0 36361 5 1 1 36360
0 36362 7 1 2 51155 36361
0 36363 7 1 2 71366 36362
0 36364 5 1 1 36363
0 36365 7 1 2 36354 36364
0 36366 5 1 1 36365
0 36367 7 1 2 43390 36366
0 36368 5 1 1 36367
0 36369 7 1 2 71363 36368
0 36370 5 1 1 36369
0 36371 7 1 2 44267 36370
0 36372 5 1 1 36371
0 36373 7 1 2 36350 36372
0 36374 5 1 1 36373
0 36375 7 1 2 62534 36374
0 36376 5 1 1 36375
0 36377 7 1 2 42628 70153
0 36378 5 1 1 36377
0 36379 7 1 2 53188 65341
0 36380 5 1 1 36379
0 36381 7 1 2 36378 36380
0 36382 5 1 1 36381
0 36383 7 1 2 60471 62359
0 36384 7 1 2 36382 36383
0 36385 5 1 1 36384
0 36386 7 1 2 36376 36385
0 36387 5 1 1 36386
0 36388 7 1 2 70293 36387
0 36389 5 1 1 36388
0 36390 7 1 2 54130 63584
0 36391 5 1 1 36390
0 36392 7 1 2 53022 4552
0 36393 5 1 1 36392
0 36394 7 1 2 45496 51156
0 36395 7 1 2 36393 36394
0 36396 5 2 1 36395
0 36397 7 1 2 36391 71367
0 36398 5 1 1 36397
0 36399 7 1 2 62535 36398
0 36400 5 1 1 36399
0 36401 7 1 2 50878 64951
0 36402 5 1 1 36401
0 36403 7 1 2 50569 53759
0 36404 5 2 1 36403
0 36405 7 2 2 62174 71369
0 36406 5 1 1 71371
0 36407 7 1 2 50797 71372
0 36408 5 1 1 36407
0 36409 7 1 2 43775 71340
0 36410 7 1 2 36408 36409
0 36411 7 1 2 36402 36410
0 36412 5 1 1 36411
0 36413 7 1 2 36400 36412
0 36414 5 1 1 36413
0 36415 7 1 2 70505 36414
0 36416 5 1 1 36415
0 36417 7 1 2 36389 36416
0 36418 5 1 1 36417
0 36419 7 1 2 51611 36418
0 36420 5 1 1 36419
0 36421 7 1 2 52513 62463
0 36422 5 1 1 36421
0 36423 7 1 2 51104 59585
0 36424 5 1 1 36423
0 36425 7 1 2 36422 36424
0 36426 5 1 1 36425
0 36427 7 1 2 70294 36426
0 36428 5 1 1 36427
0 36429 7 1 2 57249 59615
0 36430 7 1 2 69420 36429
0 36431 5 1 1 36430
0 36432 7 1 2 36428 36431
0 36433 5 1 1 36432
0 36434 7 1 2 62536 36433
0 36435 5 1 1 36434
0 36436 7 1 2 50336 64337
0 36437 5 1 1 36436
0 36438 7 1 2 47147 55476
0 36439 7 1 2 56754 36438
0 36440 5 1 1 36439
0 36441 7 1 2 36437 36440
0 36442 5 1 1 36441
0 36443 7 1 2 60472 70506
0 36444 7 1 2 36442 36443
0 36445 5 1 1 36444
0 36446 7 1 2 36435 36445
0 36447 5 1 1 36446
0 36448 7 1 2 42629 36447
0 36449 5 1 1 36448
0 36450 7 1 2 55477 60473
0 36451 5 1 1 36450
0 36452 7 1 2 10857 36451
0 36453 5 1 1 36452
0 36454 7 1 2 70507 36453
0 36455 5 1 1 36454
0 36456 7 1 2 43165 66395
0 36457 7 1 2 60594 36456
0 36458 7 1 2 65202 66217
0 36459 7 1 2 36457 36458
0 36460 5 1 1 36459
0 36461 7 1 2 36455 36460
0 36462 5 1 1 36461
0 36463 7 1 2 48698 36462
0 36464 5 1 1 36463
0 36465 7 1 2 49361 59606
0 36466 7 1 2 66361 36465
0 36467 7 1 2 61864 36466
0 36468 5 1 1 36467
0 36469 7 1 2 36464 36468
0 36470 5 1 1 36469
0 36471 7 1 2 53189 36470
0 36472 5 1 1 36471
0 36473 7 1 2 36449 36472
0 36474 5 1 1 36473
0 36475 7 1 2 42912 36474
0 36476 5 1 1 36475
0 36477 7 1 2 59633 69977
0 36478 5 1 1 36477
0 36479 7 1 2 46760 36478
0 36480 5 1 1 36479
0 36481 7 1 2 43391 35130
0 36482 5 2 1 36481
0 36483 7 1 2 36480 71373
0 36484 5 3 1 36483
0 36485 7 1 2 46335 71375
0 36486 5 1 1 36485
0 36487 7 1 2 50570 60764
0 36488 7 1 2 66436 36487
0 36489 5 1 1 36488
0 36490 7 1 2 36486 36489
0 36491 5 1 1 36490
0 36492 7 1 2 60474 36491
0 36493 5 1 1 36492
0 36494 7 1 2 46546 56852
0 36495 5 1 1 36494
0 36496 7 1 2 13517 36495
0 36497 5 1 1 36496
0 36498 7 1 2 62537 36497
0 36499 5 1 1 36498
0 36500 7 1 2 36493 36499
0 36501 5 1 1 36500
0 36502 7 1 2 56043 66476
0 36503 7 1 2 67527 36502
0 36504 7 1 2 36501 36503
0 36505 5 1 1 36504
0 36506 7 1 2 36476 36505
0 36507 5 1 1 36506
0 36508 7 1 2 51679 36507
0 36509 5 1 1 36508
0 36510 7 1 2 36420 36509
0 36511 5 1 1 36510
0 36512 7 1 2 65961 36511
0 36513 5 1 1 36512
0 36514 7 1 2 13129 71358
0 36515 5 1 1 36514
0 36516 7 1 2 51612 36515
0 36517 5 1 1 36516
0 36518 7 1 2 56125 58420
0 36519 7 1 2 58148 36518
0 36520 5 1 1 36519
0 36521 7 1 2 36517 36520
0 36522 5 1 1 36521
0 36523 7 1 2 66025 36522
0 36524 5 1 1 36523
0 36525 7 2 2 50110 71289
0 36526 5 1 1 71378
0 36527 7 1 2 50368 66464
0 36528 7 1 2 68497 36527
0 36529 5 1 1 36528
0 36530 7 1 2 36526 36529
0 36531 5 1 1 36530
0 36532 7 1 2 52906 36531
0 36533 5 1 1 36532
0 36534 7 2 2 50369 65601
0 36535 5 1 1 71380
0 36536 7 1 2 65623 71381
0 36537 5 1 1 36536
0 36538 7 1 2 36533 36537
0 36539 5 1 1 36538
0 36540 7 1 2 46336 36539
0 36541 5 1 1 36540
0 36542 7 1 2 36524 36541
0 36543 5 1 1 36542
0 36544 7 1 2 60543 36543
0 36545 5 1 1 36544
0 36546 7 2 2 68477 71240
0 36547 7 1 2 64694 71382
0 36548 5 2 1 36547
0 36549 7 1 2 60954 65756
0 36550 5 1 1 36549
0 36551 7 1 2 54900 70317
0 36552 5 2 1 36551
0 36553 7 1 2 36550 71386
0 36554 5 1 1 36553
0 36555 7 1 2 46547 36554
0 36556 5 1 1 36555
0 36557 7 1 2 56224 69706
0 36558 5 1 1 36557
0 36559 7 1 2 36556 36558
0 36560 5 1 1 36559
0 36561 7 1 2 47694 65490
0 36562 7 2 2 36560 36561
0 36563 7 1 2 45641 71388
0 36564 5 1 1 36563
0 36565 7 1 2 71384 36564
0 36566 5 2 1 36565
0 36567 7 1 2 56974 71390
0 36568 5 1 1 36567
0 36569 7 2 2 64065 65962
0 36570 5 1 1 71392
0 36571 7 1 2 71247 36570
0 36572 5 1 1 36571
0 36573 7 1 2 51680 36572
0 36574 5 1 1 36573
0 36575 7 1 2 44268 71290
0 36576 5 1 1 36575
0 36577 7 1 2 36574 36576
0 36578 5 1 1 36577
0 36579 7 1 2 46337 36578
0 36580 5 1 1 36579
0 36581 7 2 2 51717 71095
0 36582 7 3 2 63345 71394
0 36583 5 1 1 71396
0 36584 7 1 2 45314 71397
0 36585 5 1 1 36584
0 36586 7 1 2 36580 36585
0 36587 5 1 1 36586
0 36588 7 1 2 51037 36587
0 36589 5 1 1 36588
0 36590 7 1 2 57755 36184
0 36591 5 3 1 36590
0 36592 7 1 2 65963 71399
0 36593 5 1 1 36592
0 36594 7 1 2 51681 68951
0 36595 5 1 1 36594
0 36596 7 1 2 36593 36595
0 36597 5 1 1 36596
0 36598 7 1 2 45315 36597
0 36599 5 1 1 36598
0 36600 7 1 2 36583 36599
0 36601 5 1 1 36600
0 36602 7 1 2 54040 36601
0 36603 5 1 1 36602
0 36604 7 1 2 36406 71293
0 36605 5 1 1 36604
0 36606 7 1 2 64817 71291
0 36607 5 1 1 36606
0 36608 7 1 2 36605 36607
0 36609 5 1 1 36608
0 36610 7 1 2 50798 36609
0 36611 5 1 1 36610
0 36612 7 1 2 36603 36611
0 36613 7 1 2 36589 36612
0 36614 5 1 1 36613
0 36615 7 1 2 59403 36614
0 36616 5 1 1 36615
0 36617 7 1 2 51157 36616
0 36618 7 1 2 36568 36617
0 36619 7 1 2 36545 36618
0 36620 5 1 1 36619
0 36621 7 2 2 54022 60544
0 36622 5 1 1 71402
0 36623 7 1 2 56586 71403
0 36624 5 1 1 36623
0 36625 7 2 2 47819 53433
0 36626 7 2 2 60050 69061
0 36627 7 2 2 71404 71406
0 36628 5 1 1 71408
0 36629 7 1 2 36624 36628
0 36630 5 1 1 36629
0 36631 7 1 2 65757 36630
0 36632 5 1 1 36631
0 36633 7 1 2 61457 68421
0 36634 7 1 2 60805 36633
0 36635 7 1 2 69857 36634
0 36636 5 1 1 36635
0 36637 7 1 2 36632 36636
0 36638 5 1 1 36637
0 36639 7 1 2 44269 36638
0 36640 5 1 1 36639
0 36641 7 1 2 49362 59404
0 36642 5 1 1 36641
0 36643 7 1 2 50962 62591
0 36644 5 1 1 36643
0 36645 7 1 2 36642 36644
0 36646 5 1 1 36645
0 36647 7 1 2 56608 65964
0 36648 7 1 2 36646 36647
0 36649 5 1 1 36648
0 36650 7 1 2 36640 36649
0 36651 5 1 1 36650
0 36652 7 1 2 48699 36651
0 36653 5 1 1 36652
0 36654 7 2 2 54225 69732
0 36655 7 1 2 46945 71228
0 36656 7 1 2 71410 36655
0 36657 5 1 1 36656
0 36658 7 1 2 36653 36657
0 36659 5 1 1 36658
0 36660 7 1 2 60753 36659
0 36661 5 1 1 36660
0 36662 7 2 2 61654 71316
0 36663 7 1 2 49363 71412
0 36664 5 1 1 36663
0 36665 7 2 2 43562 51350
0 36666 7 1 2 45642 70878
0 36667 7 1 2 71414 36666
0 36668 5 1 1 36667
0 36669 7 1 2 36664 36668
0 36670 5 1 1 36669
0 36671 7 1 2 66026 36670
0 36672 5 1 1 36671
0 36673 7 2 2 56500 56996
0 36674 5 1 1 71416
0 36675 7 1 2 28522 36674
0 36676 5 1 1 36675
0 36677 7 1 2 49364 36676
0 36678 5 1 1 36677
0 36679 7 1 2 53342 56595
0 36680 5 1 1 36679
0 36681 7 1 2 36678 36680
0 36682 5 1 1 36681
0 36683 7 1 2 68448 36682
0 36684 5 1 1 36683
0 36685 7 1 2 36672 36684
0 36686 5 1 1 36685
0 36687 7 1 2 44270 36686
0 36688 5 1 1 36687
0 36689 7 1 2 51038 26568
0 36690 5 1 1 36689
0 36691 7 1 2 56587 67067
0 36692 7 1 2 36690 36691
0 36693 5 1 1 36692
0 36694 7 1 2 59405 60885
0 36695 7 1 2 71295 36694
0 36696 5 1 1 36695
0 36697 7 1 2 36693 36696
0 36698 5 1 1 36697
0 36699 7 1 2 48700 36698
0 36700 5 1 1 36699
0 36701 7 1 2 61003 63028
0 36702 7 1 2 61486 66655
0 36703 7 1 2 36701 36702
0 36704 5 1 1 36703
0 36705 7 1 2 36700 36704
0 36706 7 1 2 36688 36705
0 36707 5 1 1 36706
0 36708 7 1 2 42913 36707
0 36709 5 1 1 36708
0 36710 7 2 2 52303 65587
0 36711 5 1 1 71418
0 36712 7 1 2 56588 68449
0 36713 7 1 2 71419 36712
0 36714 5 1 1 36713
0 36715 7 1 2 51186 36714
0 36716 7 1 2 36709 36715
0 36717 7 1 2 36661 36716
0 36718 5 1 1 36717
0 36719 7 1 2 50478 66207
0 36720 7 1 2 36718 36719
0 36721 7 1 2 36620 36720
0 36722 5 1 1 36721
0 36723 7 3 2 65758 70295
0 36724 7 1 2 44271 70673
0 36725 5 1 1 36724
0 36726 7 1 2 71364 36725
0 36727 5 1 1 36726
0 36728 7 1 2 43392 36727
0 36729 5 1 1 36728
0 36730 7 1 2 48701 59899
0 36731 7 1 2 62091 36730
0 36732 5 1 1 36731
0 36733 7 1 2 36729 36732
0 36734 5 1 1 36733
0 36735 7 1 2 71420 36734
0 36736 5 1 1 36735
0 36737 7 4 2 50111 53035
0 36738 7 1 2 42630 71423
0 36739 5 1 1 36738
0 36740 7 1 2 71207 36739
0 36741 5 1 1 36740
0 36742 7 2 2 63743 68664
0 36743 7 1 2 44364 52535
0 36744 7 1 2 71427 36743
0 36745 7 1 2 36741 36744
0 36746 5 1 1 36745
0 36747 7 1 2 36736 36746
0 36748 5 1 1 36747
0 36749 7 1 2 62538 36748
0 36750 5 1 1 36749
0 36751 7 2 2 45643 71428
0 36752 7 1 2 68478 71429
0 36753 7 1 2 71195 36752
0 36754 5 1 1 36753
0 36755 7 1 2 36750 36754
0 36756 5 1 1 36755
0 36757 7 1 2 56589 36756
0 36758 5 1 1 36757
0 36759 7 1 2 59042 65759
0 36760 5 1 1 36759
0 36761 7 1 2 71071 36760
0 36762 5 1 1 36761
0 36763 7 1 2 51613 36762
0 36764 5 1 1 36763
0 36765 7 3 2 56960 66651
0 36766 5 1 1 71431
0 36767 7 2 2 67823 71432
0 36768 5 1 1 71434
0 36769 7 1 2 36764 36768
0 36770 5 1 1 36769
0 36771 7 1 2 70471 36770
0 36772 5 1 1 36771
0 36773 7 1 2 68667 70190
0 36774 7 1 2 71271 36773
0 36775 5 1 1 36774
0 36776 7 1 2 56975 65760
0 36777 5 1 1 36776
0 36778 7 1 2 56590 65804
0 36779 5 1 1 36778
0 36780 7 1 2 36777 36779
0 36781 5 1 1 36780
0 36782 7 1 2 63898 71057
0 36783 7 1 2 58084 36782
0 36784 7 1 2 70197 36783
0 36785 7 1 2 36781 36784
0 36786 5 1 1 36785
0 36787 7 1 2 36775 36786
0 36788 5 1 1 36787
0 36789 7 1 2 46548 36788
0 36790 5 1 1 36789
0 36791 7 1 2 36772 36790
0 36792 5 1 1 36791
0 36793 7 1 2 43776 36792
0 36794 5 1 1 36793
0 36795 7 1 2 70253 71250
0 36796 5 1 1 36795
0 36797 7 1 2 68195 70468
0 36798 7 1 2 70983 36797
0 36799 7 1 2 36796 36798
0 36800 5 1 1 36799
0 36801 7 1 2 36794 36800
0 36802 5 1 1 36801
0 36803 7 1 2 63613 36802
0 36804 5 1 1 36803
0 36805 7 1 2 36758 36804
0 36806 7 1 2 36722 36805
0 36807 7 1 2 36513 36806
0 36808 7 1 2 36343 36807
0 36809 5 1 1 36808
0 36810 7 1 2 48304 36809
0 36811 5 1 1 36810
0 36812 7 1 2 36032 36811
0 36813 7 1 2 35897 36812
0 36814 7 1 2 35637 36813
0 36815 5 1 1 36814
0 36816 7 1 2 44834 36815
0 36817 5 1 1 36816
0 36818 7 1 2 43166 57883
0 36819 5 1 1 36818
0 36820 7 1 2 12571 36819
0 36821 5 2 1 36820
0 36822 7 2 2 44974 71436
0 36823 5 1 1 71438
0 36824 7 1 2 59586 59707
0 36825 5 1 1 36824
0 36826 7 1 2 36823 36825
0 36827 5 1 1 36826
0 36828 7 1 2 51682 36827
0 36829 5 1 1 36828
0 36830 7 1 2 56379 62943
0 36831 5 1 1 36830
0 36832 7 1 2 36829 36831
0 36833 5 1 1 36832
0 36834 7 1 2 60545 36833
0 36835 5 1 1 36834
0 36836 7 1 2 56395 56501
0 36837 7 1 2 59406 36836
0 36838 7 1 2 62388 36837
0 36839 5 1 1 36838
0 36840 7 1 2 36835 36839
0 36841 5 1 1 36840
0 36842 7 1 2 42914 36841
0 36843 5 1 1 36842
0 36844 7 1 2 46549 71400
0 36845 5 1 1 36844
0 36846 7 1 2 68317 70428
0 36847 5 1 1 36846
0 36848 7 1 2 36845 36847
0 36849 5 1 1 36848
0 36850 7 1 2 59374 70720
0 36851 7 1 2 36849 36850
0 36852 5 1 1 36851
0 36853 7 1 2 36843 36852
0 36854 5 1 1 36853
0 36855 7 1 2 65965 36854
0 36856 5 1 1 36855
0 36857 7 1 2 43167 55717
0 36858 5 1 1 36857
0 36859 7 1 2 16830 36858
0 36860 5 1 1 36859
0 36861 7 1 2 60546 36860
0 36862 5 1 1 36861
0 36863 7 1 2 46946 2233
0 36864 5 1 1 36863
0 36865 7 1 2 56591 61655
0 36866 7 1 2 36864 36865
0 36867 5 1 1 36866
0 36868 7 1 2 36862 36867
0 36869 5 1 1 36868
0 36870 7 1 2 47591 36869
0 36871 5 1 1 36870
0 36872 7 1 2 55734 56502
0 36873 5 2 1 36872
0 36874 7 1 2 55725 71440
0 36875 5 1 1 36874
0 36876 7 1 2 59407 36875
0 36877 5 1 1 36876
0 36878 7 1 2 36871 36877
0 36879 5 1 1 36878
0 36880 7 1 2 46761 36879
0 36881 5 1 1 36880
0 36882 7 1 2 51632 36766
0 36883 5 1 1 36882
0 36884 7 1 2 59408 36883
0 36885 5 1 1 36884
0 36886 7 1 2 57775 59893
0 36887 7 1 2 63888 36886
0 36888 5 1 1 36887
0 36889 7 1 2 36885 36888
0 36890 5 1 1 36889
0 36891 7 1 2 46550 36890
0 36892 5 1 1 36891
0 36893 7 1 2 55712 57494
0 36894 7 1 2 61656 36893
0 36895 5 1 1 36894
0 36896 7 1 2 36892 36895
0 36897 7 1 2 36881 36896
0 36898 5 1 1 36897
0 36899 7 1 2 50571 36898
0 36900 5 1 1 36899
0 36901 7 1 2 47820 49780
0 36902 7 1 2 71407 36901
0 36903 7 1 2 51532 36902
0 36904 5 1 1 36903
0 36905 7 1 2 48305 36904
0 36906 7 1 2 36900 36905
0 36907 5 1 1 36906
0 36908 7 2 2 48702 71409
0 36909 5 1 1 71442
0 36910 7 1 2 56139 58844
0 36911 7 1 2 60689 36910
0 36912 5 1 1 36911
0 36913 7 1 2 36909 36912
0 36914 5 1 1 36913
0 36915 7 1 2 50879 36914
0 36916 5 1 1 36915
0 36917 7 2 2 50022 53434
0 36918 5 1 1 71444
0 36919 7 1 2 54041 36918
0 36920 5 1 1 36919
0 36921 7 1 2 71413 36920
0 36922 5 1 1 36921
0 36923 7 1 2 36916 36922
0 36924 5 1 1 36923
0 36925 7 1 2 48853 36924
0 36926 5 1 1 36925
0 36927 7 1 2 50023 71443
0 36928 5 1 1 36927
0 36929 7 1 2 44975 36928
0 36930 7 1 2 36926 36929
0 36931 5 1 1 36930
0 36932 7 1 2 65761 36931
0 36933 7 1 2 36907 36932
0 36934 5 1 1 36933
0 36935 7 1 2 36856 36934
0 36936 5 1 1 36935
0 36937 7 1 2 50430 36936
0 36938 5 1 1 36937
0 36939 7 1 2 53508 59504
0 36940 5 1 1 36939
0 36941 7 1 2 46551 36940
0 36942 5 1 1 36941
0 36943 7 1 2 58585 36942
0 36944 5 1 1 36943
0 36945 7 1 2 65966 36944
0 36946 5 1 1 36945
0 36947 7 1 2 57100 4133
0 36948 5 3 1 36947
0 36949 7 2 2 45497 71446
0 36950 5 1 1 71449
0 36951 7 1 2 65762 71450
0 36952 5 1 1 36951
0 36953 7 1 2 36946 36952
0 36954 5 1 1 36953
0 36955 7 1 2 60547 36954
0 36956 5 1 1 36955
0 36957 7 1 2 51453 65763
0 36958 5 1 1 36957
0 36959 7 1 2 57563 69085
0 36960 5 2 1 36959
0 36961 7 1 2 36958 71451
0 36962 5 1 1 36961
0 36963 7 1 2 59409 36962
0 36964 5 1 1 36963
0 36965 7 1 2 36956 36964
0 36966 5 1 1 36965
0 36967 7 1 2 53883 36966
0 36968 5 1 1 36967
0 36969 7 1 2 51084 69498
0 36970 5 1 1 36969
0 36971 7 1 2 66419 71447
0 36972 5 1 1 36971
0 36973 7 1 2 36970 36972
0 36974 5 1 1 36973
0 36975 7 1 2 60548 36974
0 36976 5 1 1 36975
0 36977 7 1 2 63409 70902
0 36978 5 1 1 36977
0 36979 7 1 2 64230 65967
0 36980 5 1 1 36979
0 36981 7 1 2 36978 36980
0 36982 5 1 1 36981
0 36983 7 1 2 50112 36982
0 36984 5 1 1 36983
0 36985 7 1 2 56661 65764
0 36986 5 1 1 36985
0 36987 7 1 2 71452 36986
0 36988 5 1 1 36987
0 36989 7 1 2 59410 36988
0 36990 5 1 1 36989
0 36991 7 1 2 36984 36990
0 36992 7 1 2 36976 36991
0 36993 5 1 1 36992
0 36994 7 1 2 59711 36993
0 36995 5 1 1 36994
0 36996 7 1 2 36968 36995
0 36997 5 1 1 36996
0 36998 7 1 2 51614 36997
0 36999 5 1 1 36998
0 37000 7 1 2 59411 59628
0 37001 5 1 1 37000
0 37002 7 1 2 12152 37001
0 37003 5 1 1 37002
0 37004 7 1 2 65765 37003
0 37005 5 1 1 37004
0 37006 7 1 2 59803 67845
0 37007 5 1 1 37006
0 37008 7 1 2 37005 37007
0 37009 5 1 1 37008
0 37010 7 1 2 47592 37009
0 37011 5 1 1 37010
0 37012 7 1 2 59412 63870
0 37013 7 1 2 70786 37012
0 37014 5 1 1 37013
0 37015 7 1 2 37011 37014
0 37016 5 1 1 37015
0 37017 7 1 2 46762 37016
0 37018 5 1 1 37017
0 37019 7 1 2 57564 65820
0 37020 5 1 1 37019
0 37021 7 1 2 52079 66027
0 37022 5 1 1 37021
0 37023 7 1 2 37020 37022
0 37024 5 1 1 37023
0 37025 7 1 2 70119 37024
0 37026 5 1 1 37025
0 37027 7 1 2 30763 71073
0 37028 5 1 1 37027
0 37029 7 1 2 50880 37028
0 37030 5 1 1 37029
0 37031 7 1 2 68610 69086
0 37032 5 1 1 37031
0 37033 7 1 2 37030 37032
0 37034 5 1 1 37033
0 37035 7 1 2 60549 37034
0 37036 5 1 1 37035
0 37037 7 1 2 37026 37036
0 37038 7 1 2 37018 37037
0 37039 5 1 1 37038
0 37040 7 1 2 53884 37039
0 37041 5 1 1 37040
0 37042 7 1 2 50881 59621
0 37043 5 1 1 37042
0 37044 7 1 2 57101 37043
0 37045 5 1 1 37044
0 37046 7 1 2 65766 37045
0 37047 5 1 1 37046
0 37048 7 1 2 65501 69291
0 37049 5 1 1 37048
0 37050 7 1 2 37047 37049
0 37051 5 1 1 37050
0 37052 7 1 2 46552 37051
0 37053 5 1 1 37052
0 37054 7 1 2 50799 66094
0 37055 5 1 1 37054
0 37056 7 1 2 60205 65968
0 37057 5 1 1 37056
0 37058 7 1 2 37055 37057
0 37059 5 1 1 37058
0 37060 7 1 2 43168 37059
0 37061 5 1 1 37060
0 37062 7 1 2 25613 71248
0 37063 5 1 1 37062
0 37064 7 1 2 57152 37063
0 37065 5 1 1 37064
0 37066 7 1 2 37061 37065
0 37067 5 1 1 37066
0 37068 7 1 2 45316 37067
0 37069 5 1 1 37068
0 37070 7 1 2 37053 37069
0 37071 5 1 1 37070
0 37072 7 1 2 60550 37071
0 37073 5 1 1 37072
0 37074 7 1 2 50190 50963
0 37075 5 1 1 37074
0 37076 7 1 2 61657 37075
0 37077 7 1 2 71393 37076
0 37078 5 1 1 37077
0 37079 7 1 2 37073 37078
0 37080 5 1 1 37079
0 37081 7 1 2 59712 37080
0 37082 5 1 1 37081
0 37083 7 1 2 37041 37082
0 37084 5 1 1 37083
0 37085 7 1 2 51683 37084
0 37086 5 1 1 37085
0 37087 7 1 2 36999 37086
0 37088 5 1 1 37087
0 37089 7 1 2 46338 37088
0 37090 5 1 1 37089
0 37091 7 1 2 49843 71352
0 37092 5 1 1 37091
0 37093 7 1 2 42915 58860
0 37094 5 1 1 37093
0 37095 7 1 2 37092 37094
0 37096 5 1 1 37095
0 37097 7 1 2 46553 37096
0 37098 5 1 1 37097
0 37099 7 1 2 51615 62301
0 37100 5 1 1 37099
0 37101 7 1 2 37098 37100
0 37102 5 2 1 37101
0 37103 7 1 2 70587 71453
0 37104 5 1 1 37103
0 37105 7 1 2 61500 65767
0 37106 5 1 1 37105
0 37107 7 1 2 65675 65969
0 37108 5 2 1 37107
0 37109 7 1 2 37106 71455
0 37110 5 1 1 37109
0 37111 7 1 2 51616 37110
0 37112 5 1 1 37111
0 37113 7 1 2 49922 65970
0 37114 7 1 2 57799 37113
0 37115 5 2 1 37114
0 37116 7 1 2 37112 71457
0 37117 5 1 1 37116
0 37118 7 1 2 59413 37117
0 37119 5 1 1 37118
0 37120 7 1 2 37104 37119
0 37121 5 1 1 37120
0 37122 7 1 2 50572 37121
0 37123 5 1 1 37122
0 37124 7 1 2 49781 61658
0 37125 7 1 2 71398 37124
0 37126 5 1 1 37125
0 37127 7 1 2 37123 37126
0 37128 5 1 1 37127
0 37129 7 1 2 59713 37128
0 37130 5 1 1 37129
0 37131 7 1 2 37090 37130
0 37132 7 1 2 36938 37131
0 37133 5 1 1 37132
0 37134 7 1 2 66208 37133
0 37135 5 1 1 37134
0 37136 7 1 2 51409 53172
0 37137 5 1 1 37136
0 37138 7 1 2 9472 37137
0 37139 5 1 1 37138
0 37140 7 1 2 45498 37139
0 37141 5 1 1 37140
0 37142 7 1 2 54901 62360
0 37143 5 1 1 37142
0 37144 7 1 2 37141 37143
0 37145 5 1 1 37144
0 37146 7 1 2 51617 37145
0 37147 5 1 1 37146
0 37148 7 3 2 46947 55819
0 37149 5 1 1 71459
0 37150 7 1 2 55152 71460
0 37151 5 1 1 37150
0 37152 7 1 2 37147 37151
0 37153 5 1 1 37152
0 37154 7 1 2 47457 37153
0 37155 5 1 1 37154
0 37156 7 1 2 36034 71332
0 37157 5 1 1 37156
0 37158 7 1 2 42916 37157
0 37159 5 1 1 37158
0 37160 7 1 2 634 71333
0 37161 5 1 1 37160
0 37162 7 1 2 49717 37161
0 37163 5 1 1 37162
0 37164 7 1 2 37159 37163
0 37165 5 1 1 37164
0 37166 7 1 2 58519 37165
0 37167 5 1 1 37166
0 37168 7 1 2 37155 37167
0 37169 5 1 1 37168
0 37170 7 1 2 47148 37169
0 37171 5 1 1 37170
0 37172 7 1 2 68050 20459
0 37173 5 1 1 37172
0 37174 7 1 2 58569 37173
0 37175 5 1 1 37174
0 37176 7 1 2 55718 62438
0 37177 5 1 1 37176
0 37178 7 1 2 37175 37177
0 37179 5 1 1 37178
0 37180 7 1 2 51067 37179
0 37181 5 1 1 37180
0 37182 7 1 2 37171 37181
0 37183 5 1 1 37182
0 37184 7 1 2 70508 37183
0 37185 5 1 1 37184
0 37186 7 1 2 70525 71454
0 37187 5 1 1 37186
0 37188 7 1 2 37185 37187
0 37189 5 1 1 37188
0 37190 7 1 2 44976 37189
0 37191 5 1 1 37190
0 37192 7 1 2 70549 70564
0 37193 5 1 1 37192
0 37194 7 2 2 51063 52434
0 37195 7 1 2 50573 51684
0 37196 7 1 2 71462 37195
0 37197 7 1 2 37193 37196
0 37198 5 1 1 37197
0 37199 7 1 2 37191 37198
0 37200 5 1 1 37199
0 37201 7 1 2 62539 37200
0 37202 5 1 1 37201
0 37203 7 1 2 55478 70509
0 37204 5 1 1 37203
0 37205 7 1 2 60235 70527
0 37206 7 1 2 70530 37205
0 37207 5 1 1 37206
0 37208 7 1 2 37204 37207
0 37209 5 1 1 37208
0 37210 7 1 2 56697 37209
0 37211 5 1 1 37210
0 37212 7 1 2 43482 69875
0 37213 7 3 2 48306 52855
0 37214 7 1 2 69285 71464
0 37215 7 1 2 37212 37214
0 37216 5 1 1 37215
0 37217 7 1 2 37211 37216
0 37218 5 1 1 37217
0 37219 7 2 2 56410 58263
0 37220 7 1 2 51685 71467
0 37221 7 1 2 37218 37220
0 37222 5 1 1 37221
0 37223 7 1 2 37202 37222
0 37224 5 1 1 37223
0 37225 7 1 2 66028 37224
0 37226 5 1 1 37225
0 37227 7 1 2 61917 68952
0 37228 7 1 2 70227 37227
0 37229 5 1 1 37228
0 37230 7 2 2 45870 66174
0 37231 7 1 2 63360 63456
0 37232 7 1 2 71469 37231
0 37233 5 1 1 37232
0 37234 7 1 2 37229 37233
0 37235 5 1 1 37234
0 37236 7 1 2 46339 37235
0 37237 5 1 1 37236
0 37238 7 1 2 68925 69332
0 37239 7 1 2 71470 37238
0 37240 5 1 1 37239
0 37241 7 1 2 37237 37240
0 37242 5 1 1 37241
0 37243 7 1 2 46554 37242
0 37244 5 1 1 37243
0 37245 7 1 2 64120 64531
0 37246 7 1 2 58582 37245
0 37247 7 1 2 66209 37246
0 37248 5 1 1 37247
0 37249 7 1 2 37244 37248
0 37250 5 1 1 37249
0 37251 7 1 2 45644 37250
0 37252 5 1 1 37251
0 37253 7 1 2 63763 64255
0 37254 7 1 2 51085 37253
0 37255 7 1 2 69817 37254
0 37256 5 1 1 37255
0 37257 7 1 2 37252 37256
0 37258 5 1 1 37257
0 37259 7 1 2 47695 37258
0 37260 5 1 1 37259
0 37261 7 2 2 59375 69421
0 37262 7 2 2 44496 65768
0 37263 7 1 2 71424 71473
0 37264 7 1 2 71471 37263
0 37265 5 1 1 37264
0 37266 7 1 2 37260 37265
0 37267 5 1 1 37266
0 37268 7 1 2 53933 37267
0 37269 5 1 1 37268
0 37270 7 2 2 52435 70232
0 37271 7 1 2 45317 71475
0 37272 5 1 1 37271
0 37273 7 1 2 4897 65343
0 37274 5 1 1 37273
0 37275 7 1 2 924 61778
0 37276 7 1 2 37274 37275
0 37277 5 1 1 37276
0 37278 7 1 2 53892 37277
0 37279 5 1 1 37278
0 37280 7 1 2 50800 57565
0 37281 7 1 2 37279 37280
0 37282 5 1 1 37281
0 37283 7 1 2 37272 37282
0 37284 5 1 1 37283
0 37285 7 1 2 45499 37284
0 37286 5 1 1 37285
0 37287 7 1 2 56740 71463
0 37288 5 1 1 37287
0 37289 7 1 2 37286 37288
0 37290 5 1 1 37289
0 37291 7 1 2 71472 37290
0 37292 5 1 1 37291
0 37293 7 1 2 60253 60497
0 37294 7 1 2 66234 37293
0 37295 7 1 2 65451 37294
0 37296 5 1 1 37295
0 37297 7 1 2 37292 37296
0 37298 5 1 1 37297
0 37299 7 1 2 71474 37298
0 37300 5 1 1 37299
0 37301 7 1 2 52520 59684
0 37302 7 1 2 64601 65427
0 37303 7 1 2 37301 37302
0 37304 7 1 2 70275 37303
0 37305 7 1 2 71192 37304
0 37306 5 1 1 37305
0 37307 7 1 2 37300 37306
0 37308 7 1 2 37269 37307
0 37309 5 1 1 37308
0 37310 7 1 2 56592 37309
0 37311 5 1 1 37310
0 37312 7 2 2 42348 56136
0 37313 7 1 2 47924 55444
0 37314 7 1 2 57331 37313
0 37315 7 1 2 71477 37314
0 37316 5 1 1 37315
0 37317 7 1 2 49499 58013
0 37318 7 1 2 70130 37317
0 37319 7 1 2 65815 37318
0 37320 5 1 1 37319
0 37321 7 1 2 37316 37320
0 37322 5 1 1 37321
0 37323 7 1 2 59972 37322
0 37324 5 1 1 37323
0 37325 7 2 2 55445 70173
0 37326 7 1 2 66465 71415
0 37327 7 1 2 71479 37326
0 37328 5 1 1 37327
0 37329 7 1 2 56646 57800
0 37330 7 1 2 70793 37329
0 37331 5 1 1 37330
0 37332 7 1 2 37328 37331
0 37333 5 1 1 37332
0 37334 7 1 2 47149 37333
0 37335 5 1 1 37334
0 37336 7 1 2 37324 37335
0 37337 5 1 1 37336
0 37338 7 1 2 70510 37337
0 37339 5 1 1 37338
0 37340 7 1 2 43169 71335
0 37341 5 1 1 37340
0 37342 7 1 2 71320 37341
0 37343 5 1 1 37342
0 37344 7 1 2 50882 37343
0 37345 5 1 1 37344
0 37346 7 1 2 57804 60821
0 37347 5 1 1 37346
0 37348 7 1 2 37345 37347
0 37349 5 1 1 37348
0 37350 7 1 2 48703 37349
0 37351 5 1 1 37350
0 37352 7 1 2 49888 71417
0 37353 5 1 1 37352
0 37354 7 1 2 37351 37353
0 37355 5 1 1 37354
0 37356 7 1 2 65971 37355
0 37357 5 1 1 37356
0 37358 7 1 2 44692 55673
0 37359 7 1 2 51711 37358
0 37360 7 1 2 71478 37359
0 37361 5 1 1 37360
0 37362 7 1 2 37357 37361
0 37363 5 1 1 37362
0 37364 7 1 2 60797 67773
0 37365 7 1 2 70475 37364
0 37366 7 1 2 37363 37365
0 37367 5 1 1 37366
0 37368 7 1 2 37339 37367
0 37369 5 1 1 37368
0 37370 7 1 2 62540 37369
0 37371 5 1 1 37370
0 37372 7 1 2 49059 70511
0 37373 5 1 1 37372
0 37374 7 1 2 61937 70296
0 37375 5 1 1 37374
0 37376 7 1 2 37373 37375
0 37377 5 1 1 37376
0 37378 7 1 2 65769 37377
0 37379 5 1 1 37378
0 37380 7 1 2 61474 68211
0 37381 7 1 2 71301 37380
0 37382 5 1 1 37381
0 37383 7 1 2 37379 37382
0 37384 5 1 1 37383
0 37385 7 1 2 70039 37384
0 37386 5 1 1 37385
0 37387 7 1 2 49242 71299
0 37388 5 1 1 37387
0 37389 7 1 2 50964 65811
0 37390 7 1 2 70297 37389
0 37391 5 1 1 37390
0 37392 7 1 2 37388 37391
0 37393 5 1 1 37392
0 37394 7 1 2 70040 37393
0 37395 5 1 1 37394
0 37396 7 2 2 68263 70544
0 37397 7 1 2 70930 71481
0 37398 5 1 1 37397
0 37399 7 1 2 70041 71421
0 37400 5 1 1 37399
0 37401 7 1 2 37398 37400
0 37402 5 1 1 37401
0 37403 7 1 2 49365 37402
0 37404 5 1 1 37403
0 37405 7 1 2 51864 69458
0 37406 7 1 2 71482 37405
0 37407 5 1 1 37406
0 37408 7 1 2 69712 71083
0 37409 5 1 1 37408
0 37410 7 1 2 57877 63790
0 37411 7 1 2 66175 37410
0 37412 7 1 2 37409 37411
0 37413 5 1 1 37412
0 37414 7 1 2 37407 37413
0 37415 7 1 2 37404 37414
0 37416 5 1 1 37415
0 37417 7 1 2 49060 37416
0 37418 5 1 1 37417
0 37419 7 1 2 37395 37418
0 37420 5 1 1 37419
0 37421 7 1 2 43393 37420
0 37422 5 1 1 37421
0 37423 7 1 2 37386 37422
0 37424 5 1 1 37423
0 37425 7 1 2 71468 37424
0 37426 5 1 1 37425
0 37427 7 1 2 37371 37426
0 37428 5 1 1 37427
0 37429 7 1 2 42917 37428
0 37430 5 1 1 37429
0 37431 7 1 2 57814 65770
0 37432 5 1 1 37431
0 37433 7 1 2 71456 37432
0 37434 5 1 1 37433
0 37435 7 1 2 51618 37434
0 37436 5 2 1 37435
0 37437 7 1 2 71458 71483
0 37438 5 1 1 37437
0 37439 7 1 2 45318 37438
0 37440 5 1 1 37439
0 37441 7 1 2 50270 70978
0 37442 5 1 1 37441
0 37443 7 1 2 37440 37442
0 37444 5 1 1 37443
0 37445 7 1 2 47458 37444
0 37446 5 1 1 37445
0 37447 7 1 2 57495 58570
0 37448 7 1 2 65771 66590
0 37449 7 1 2 37447 37448
0 37450 5 1 1 37449
0 37451 7 1 2 37446 37450
0 37452 5 1 1 37451
0 37453 7 1 2 60475 37452
0 37454 5 1 1 37453
0 37455 7 2 2 55787 62220
0 37456 7 1 2 57496 70418
0 37457 7 1 2 71485 37456
0 37458 5 1 1 37457
0 37459 7 1 2 37454 37458
0 37460 5 1 1 37459
0 37461 7 1 2 53292 37460
0 37462 5 1 1 37461
0 37463 7 1 2 50431 65588
0 37464 7 1 2 68532 37463
0 37465 7 1 2 57795 37464
0 37466 5 1 1 37465
0 37467 7 1 2 37462 37466
0 37468 5 1 1 37467
0 37469 7 1 2 70512 37468
0 37470 5 1 1 37469
0 37471 7 1 2 37430 37470
0 37472 5 1 1 37471
0 37473 7 1 2 44977 37472
0 37474 5 1 1 37473
0 37475 7 1 2 51686 65821
0 37476 7 1 2 62577 37475
0 37477 5 1 1 37476
0 37478 7 1 2 71484 37477
0 37479 5 1 1 37478
0 37480 7 1 2 70513 37479
0 37481 5 1 1 37480
0 37482 7 1 2 56961 58080
0 37483 7 1 2 63950 64435
0 37484 7 1 2 37482 37483
0 37485 7 1 2 66454 69470
0 37486 7 1 2 37484 37485
0 37487 5 1 1 37486
0 37488 7 1 2 37481 37487
0 37489 5 1 1 37488
0 37490 7 1 2 60476 37489
0 37491 5 1 1 37490
0 37492 7 1 2 55726 5761
0 37493 5 2 1 37492
0 37494 7 1 2 70623 71487
0 37495 5 1 1 37494
0 37496 7 2 2 62680 68188
0 37497 7 1 2 60573 63836
0 37498 7 1 2 66662 37497
0 37499 7 1 2 71489 37498
0 37500 7 1 2 63697 37499
0 37501 5 1 1 37500
0 37502 7 1 2 37495 37501
0 37503 5 1 1 37502
0 37504 7 1 2 62541 37503
0 37505 5 1 1 37504
0 37506 7 1 2 37491 37505
0 37507 5 1 1 37506
0 37508 7 1 2 47459 37507
0 37509 5 1 1 37508
0 37510 7 1 2 46555 71488
0 37511 5 1 1 37510
0 37512 7 1 2 51619 52324
0 37513 5 1 1 37512
0 37514 7 1 2 37511 37513
0 37515 5 1 1 37514
0 37516 7 1 2 70782 37515
0 37517 5 1 1 37516
0 37518 7 1 2 57497 59228
0 37519 7 1 2 70972 37518
0 37520 5 1 1 37519
0 37521 7 1 2 37517 37520
0 37522 5 1 1 37521
0 37523 7 1 2 70514 37522
0 37524 5 1 1 37523
0 37525 7 1 2 37509 37524
0 37526 5 1 1 37525
0 37527 7 1 2 45319 37526
0 37528 5 1 1 37527
0 37529 7 1 2 47460 55740
0 37530 5 1 1 37529
0 37531 7 1 2 17625 37530
0 37532 5 1 1 37531
0 37533 7 1 2 70783 37532
0 37534 5 1 1 37533
0 37535 7 1 2 46556 54508
0 37536 7 1 2 70122 37535
0 37537 7 1 2 64638 37536
0 37538 5 1 1 37537
0 37539 7 1 2 37534 37538
0 37540 5 1 1 37539
0 37541 7 1 2 50801 70515
0 37542 7 1 2 37540 37541
0 37543 5 1 1 37542
0 37544 7 1 2 37528 37543
0 37545 5 1 1 37544
0 37546 7 1 2 53885 37545
0 37547 5 1 1 37546
0 37548 7 1 2 49782 71343
0 37549 5 1 1 37548
0 37550 7 1 2 57645 70123
0 37551 7 1 2 59417 37550
0 37552 5 1 1 37551
0 37553 7 1 2 37549 37552
0 37554 5 1 1 37553
0 37555 7 1 2 65772 37554
0 37556 5 1 1 37555
0 37557 7 1 2 57926 60051
0 37558 7 1 2 63102 69029
0 37559 7 1 2 37557 37558
0 37560 5 1 1 37559
0 37561 7 1 2 37556 37560
0 37562 5 1 1 37561
0 37563 7 1 2 70516 37562
0 37564 5 1 1 37563
0 37565 7 1 2 61277 63951
0 37566 7 1 2 66319 37565
0 37567 7 1 2 69034 70542
0 37568 7 1 2 71259 37567
0 37569 7 1 2 37566 37568
0 37570 5 1 1 37569
0 37571 7 1 2 37564 37570
0 37572 5 1 1 37571
0 37573 7 1 2 59714 37572
0 37574 5 1 1 37573
0 37575 7 2 2 67134 70537
0 37576 7 1 2 45500 68993
0 37577 7 1 2 71491 37576
0 37578 5 1 1 37577
0 37579 7 1 2 35901 37578
0 37580 5 1 1 37579
0 37581 7 1 2 71326 37580
0 37582 5 1 1 37581
0 37583 7 1 2 45320 71492
0 37584 5 1 1 37583
0 37585 7 1 2 70550 37584
0 37586 5 1 1 37585
0 37587 7 1 2 55719 68533
0 37588 7 1 2 37586 37587
0 37589 5 1 1 37588
0 37590 7 1 2 37582 37589
0 37591 5 1 1 37590
0 37592 7 1 2 49306 37591
0 37593 5 1 1 37592
0 37594 7 2 2 59213 66362
0 37595 7 2 2 43563 63103
0 37596 5 1 1 71495
0 37597 7 1 2 68699 70903
0 37598 7 1 2 71496 37597
0 37599 7 1 2 71493 37598
0 37600 5 1 1 37599
0 37601 7 1 2 37593 37600
0 37602 5 1 1 37601
0 37603 7 1 2 71476 37602
0 37604 5 1 1 37603
0 37605 7 1 2 37574 37604
0 37606 5 1 1 37605
0 37607 7 1 2 50113 37606
0 37608 5 1 1 37607
0 37609 7 1 2 66210 71391
0 37610 5 1 1 37609
0 37611 7 1 2 66226 71389
0 37612 5 1 1 37611
0 37613 7 1 2 62180 70624
0 37614 5 1 1 37613
0 37615 7 2 2 44693 63614
0 37616 7 1 2 59817 70221
0 37617 7 1 2 71497 37616
0 37618 5 1 1 37617
0 37619 7 1 2 37614 37618
0 37620 5 1 1 37619
0 37621 7 1 2 50802 37620
0 37622 5 1 1 37621
0 37623 7 1 2 58069 63283
0 37624 7 1 2 63744 66389
0 37625 7 1 2 37623 37624
0 37626 7 1 2 64972 37625
0 37627 5 1 1 37626
0 37628 7 1 2 37622 37627
0 37629 5 1 1 37628
0 37630 7 1 2 60477 37629
0 37631 5 1 1 37630
0 37632 7 1 2 37612 37631
0 37633 7 1 2 37610 37632
0 37634 5 1 1 37633
0 37635 7 1 2 59715 37634
0 37636 5 1 1 37635
0 37637 7 1 2 65460 67068
0 37638 5 1 1 37637
0 37639 7 1 2 71385 37638
0 37640 5 2 1 37639
0 37641 7 1 2 66211 71499
0 37642 5 1 1 37641
0 37643 7 1 2 71430 71383
0 37644 5 1 1 37643
0 37645 7 1 2 53045 70625
0 37646 5 1 1 37645
0 37647 7 1 2 65457 71422
0 37648 5 1 1 37647
0 37649 7 1 2 37646 37648
0 37650 5 1 1 37649
0 37651 7 1 2 63724 37650
0 37652 5 1 1 37651
0 37653 7 1 2 37644 37652
0 37654 7 1 2 37642 37653
0 37655 5 1 1 37654
0 37656 7 1 2 53886 37655
0 37657 5 1 1 37656
0 37658 7 1 2 37636 37657
0 37659 5 1 1 37658
0 37660 7 1 2 56976 37659
0 37661 5 1 1 37660
0 37662 7 1 2 37608 37661
0 37663 7 1 2 37547 37662
0 37664 7 1 2 37474 37663
0 37665 7 1 2 37311 37664
0 37666 7 1 2 37226 37665
0 37667 7 1 2 37135 37666
0 37668 7 1 2 50432 71437
0 37669 5 1 1 37668
0 37670 7 1 2 62338 62623
0 37671 5 1 1 37670
0 37672 7 1 2 37669 37671
0 37673 5 1 1 37672
0 37674 7 1 2 65773 37673
0 37675 5 1 1 37674
0 37676 7 2 2 55494 64555
0 37677 7 2 2 63299 63378
0 37678 7 1 2 71501 71503
0 37679 5 1 1 37678
0 37680 7 1 2 37675 37679
0 37681 5 1 1 37680
0 37682 7 1 2 59797 37681
0 37683 5 1 1 37682
0 37684 7 1 2 66976 35296
0 37685 5 1 1 37684
0 37686 7 1 2 50883 37685
0 37687 5 1 1 37686
0 37688 7 1 2 68482 37687
0 37689 5 1 1 37688
0 37690 7 1 2 59924 62960
0 37691 7 1 2 37689 37690
0 37692 5 1 1 37691
0 37693 7 1 2 37683 37692
0 37694 5 1 1 37693
0 37695 7 1 2 42918 37694
0 37696 5 1 1 37695
0 37697 7 1 2 59376 63336
0 37698 7 1 2 52514 37697
0 37699 7 1 2 71256 37698
0 37700 5 1 1 37699
0 37701 7 1 2 37696 37700
0 37702 5 1 1 37701
0 37703 7 1 2 56923 70802
0 37704 7 1 2 37702 37703
0 37705 5 1 1 37704
0 37706 7 1 2 67715 71356
0 37707 5 1 1 37706
0 37708 7 1 2 62552 11129
0 37709 5 1 1 37708
0 37710 7 1 2 46948 63655
0 37711 7 1 2 37709 37710
0 37712 5 1 1 37711
0 37713 7 1 2 37707 37712
0 37714 5 1 1 37713
0 37715 7 1 2 65774 37714
0 37716 5 1 1 37715
0 37717 7 2 2 48037 50803
0 37718 7 1 2 63123 71505
0 37719 7 1 2 56933 37718
0 37720 5 1 1 37719
0 37721 7 1 2 37716 37720
0 37722 5 1 1 37721
0 37723 7 1 2 42919 37722
0 37724 5 1 1 37723
0 37725 7 1 2 63719 65627
0 37726 7 1 2 66531 37725
0 37727 5 1 1 37726
0 37728 7 1 2 37724 37727
0 37729 5 1 1 37728
0 37730 7 1 2 47696 37729
0 37731 5 1 1 37730
0 37732 7 1 2 56362 70423
0 37733 5 1 1 37732
0 37734 7 1 2 37731 37733
0 37735 5 1 1 37734
0 37736 7 1 2 46557 37735
0 37737 5 1 1 37736
0 37738 7 1 2 62480 65624
0 37739 7 1 2 63901 66532
0 37740 7 1 2 37738 37739
0 37741 5 1 1 37740
0 37742 7 1 2 46863 37741
0 37743 7 1 2 37737 37742
0 37744 5 1 1 37743
0 37745 7 1 2 42083 57425
0 37746 7 1 2 66095 37745
0 37747 5 1 1 37746
0 37748 7 1 2 55208 63124
0 37749 7 1 2 56615 37748
0 37750 5 1 1 37749
0 37751 7 1 2 37747 37750
0 37752 5 1 1 37751
0 37753 7 1 2 60652 37752
0 37754 5 1 1 37753
0 37755 7 1 2 66533 70163
0 37756 7 1 2 70589 37755
0 37757 5 1 1 37756
0 37758 7 1 2 37754 37757
0 37759 5 1 1 37758
0 37760 7 1 2 47593 37759
0 37761 5 1 1 37760
0 37762 7 2 2 56934 70386
0 37763 5 1 1 71507
0 37764 7 1 2 55428 55641
0 37765 7 1 2 63125 64542
0 37766 7 1 2 37764 37765
0 37767 5 1 1 37766
0 37768 7 1 2 37763 37767
0 37769 5 1 1 37768
0 37770 7 1 2 44365 37769
0 37771 5 1 1 37770
0 37772 7 1 2 37761 37771
0 37773 5 1 1 37772
0 37774 7 1 2 46763 37773
0 37775 5 1 1 37774
0 37776 7 1 2 59377 70376
0 37777 5 1 1 37776
0 37778 7 2 2 64240 70164
0 37779 5 1 1 71509
0 37780 7 1 2 65775 71510
0 37781 5 1 1 37780
0 37782 7 1 2 30033 37781
0 37783 5 1 1 37782
0 37784 7 1 2 45501 59894
0 37785 7 1 2 37783 37784
0 37786 5 1 1 37785
0 37787 7 1 2 37777 37786
0 37788 5 1 1 37787
0 37789 7 1 2 46558 37788
0 37790 5 1 1 37789
0 37791 7 1 2 60131 71508
0 37792 5 1 1 37791
0 37793 7 1 2 43483 37792
0 37794 7 1 2 37790 37793
0 37795 7 1 2 37775 37794
0 37796 5 1 1 37795
0 37797 7 1 2 50574 37796
0 37798 7 1 2 37744 37797
0 37799 5 1 1 37798
0 37800 7 1 2 49764 61929
0 37801 7 1 2 71088 37800
0 37802 7 1 2 70406 37801
0 37803 5 1 1 37802
0 37804 7 1 2 37799 37803
0 37805 5 1 1 37804
0 37806 7 1 2 53934 37805
0 37807 5 1 1 37806
0 37808 7 1 2 55657 60186
0 37809 7 2 2 56203 37808
0 37810 5 1 1 71511
0 37811 7 1 2 54834 70061
0 37812 7 1 2 70352 37811
0 37813 5 1 1 37812
0 37814 7 1 2 37810 37813
0 37815 5 1 1 37814
0 37816 7 1 2 46096 37815
0 37817 5 1 1 37816
0 37818 7 2 2 44600 51380
0 37819 7 1 2 61352 70867
0 37820 7 1 2 71513 37819
0 37821 5 1 1 37820
0 37822 7 1 2 37817 37821
0 37823 5 1 1 37822
0 37824 7 1 2 49307 37823
0 37825 5 1 1 37824
0 37826 7 1 2 46097 45321
0 37827 7 1 2 71512 37826
0 37828 5 1 1 37827
0 37829 7 1 2 37825 37828
0 37830 5 1 1 37829
0 37831 7 1 2 42084 51039
0 37832 7 1 2 37830 37831
0 37833 5 1 1 37832
0 37834 7 2 2 53634 55735
0 37835 5 1 1 71515
0 37836 7 1 2 56717 71516
0 37837 7 1 2 61472 37836
0 37838 5 1 1 37837
0 37839 7 1 2 37833 37838
0 37840 5 1 1 37839
0 37841 7 1 2 50114 37840
0 37842 5 1 1 37841
0 37843 7 1 2 66856 71439
0 37844 5 1 1 37843
0 37845 7 1 2 42920 51213
0 37846 5 2 1 37845
0 37847 7 1 2 65447 71517
0 37848 5 1 1 37847
0 37849 7 1 2 49796 37848
0 37850 5 1 1 37849
0 37851 7 1 2 50638 50804
0 37852 7 1 2 57300 37851
0 37853 5 1 1 37852
0 37854 7 1 2 37850 37853
0 37855 5 1 1 37854
0 37856 7 1 2 59864 37855
0 37857 5 1 1 37856
0 37858 7 1 2 37844 37857
0 37859 5 1 1 37858
0 37860 7 1 2 43564 50484
0 37861 7 1 2 37859 37860
0 37862 5 1 1 37861
0 37863 7 1 2 37842 37862
0 37864 5 1 1 37863
0 37865 7 1 2 65972 37864
0 37866 5 1 1 37865
0 37867 7 1 2 61780 65560
0 37868 5 1 1 37867
0 37869 7 1 2 59973 63716
0 37870 5 1 1 37869
0 37871 7 1 2 70568 37870
0 37872 5 1 1 37871
0 37873 7 1 2 59865 37872
0 37874 5 1 1 37873
0 37875 7 1 2 37868 37874
0 37876 5 1 1 37875
0 37877 7 1 2 42921 37876
0 37878 5 1 1 37877
0 37879 7 1 2 59616 65017
0 37880 7 1 2 69163 37879
0 37881 5 1 1 37880
0 37882 7 1 2 37878 37881
0 37883 5 1 1 37882
0 37884 7 1 2 44978 37883
0 37885 5 1 1 37884
0 37886 7 1 2 60148 70067
0 37887 7 1 2 52206 37886
0 37888 5 1 1 37887
0 37889 7 1 2 37885 37888
0 37890 5 1 1 37889
0 37891 7 1 2 70466 37890
0 37892 5 1 1 37891
0 37893 7 1 2 37866 37892
0 37894 5 1 1 37893
0 37895 7 1 2 44497 37894
0 37896 5 1 1 37895
0 37897 7 1 2 53935 71500
0 37898 5 1 1 37897
0 37899 7 2 2 57281 63094
0 37900 7 1 2 53293 70019
0 37901 7 1 2 71519 37900
0 37902 7 1 2 65840 37901
0 37903 5 1 1 37902
0 37904 7 1 2 37898 37903
0 37905 5 1 1 37904
0 37906 7 1 2 66681 37905
0 37907 5 1 1 37906
0 37908 7 1 2 37896 37907
0 37909 7 1 2 37807 37908
0 37910 7 1 2 37705 37909
0 37911 7 1 2 53294 71186
0 37912 5 1 1 37911
0 37913 7 1 2 62944 65216
0 37914 5 1 1 37913
0 37915 7 1 2 37912 37914
0 37916 5 1 1 37915
0 37917 7 1 2 70370 37916
0 37918 5 1 1 37917
0 37919 7 1 2 49366 52348
0 37920 5 1 1 37919
0 37921 7 1 2 57488 37920
0 37922 5 1 1 37921
0 37923 7 1 2 42922 37922
0 37924 5 1 1 37923
0 37925 7 1 2 36711 37924
0 37926 5 1 1 37925
0 37927 7 1 2 56049 63570
0 37928 7 1 2 37926 37927
0 37929 5 1 1 37928
0 37930 7 1 2 37918 37929
0 37931 5 1 1 37930
0 37932 7 1 2 65973 37931
0 37933 5 1 1 37932
0 37934 7 2 2 56126 60806
0 37935 5 1 1 71521
0 37936 7 1 2 60822 71522
0 37937 5 1 1 37936
0 37938 7 2 2 57776 63556
0 37939 5 1 1 71523
0 37940 7 1 2 44126 71524
0 37941 5 1 1 37940
0 37942 7 1 2 37935 37941
0 37943 5 1 1 37942
0 37944 7 1 2 43170 37943
0 37945 5 1 1 37944
0 37946 7 1 2 35553 37939
0 37947 5 1 1 37946
0 37948 7 1 2 42923 37947
0 37949 5 1 1 37948
0 37950 7 1 2 37945 37949
0 37951 5 1 1 37950
0 37952 7 1 2 43394 37951
0 37953 5 1 1 37952
0 37954 7 1 2 63819 37779
0 37955 5 1 1 37954
0 37956 7 1 2 54023 37955
0 37957 5 1 1 37956
0 37958 7 1 2 37953 37957
0 37959 5 1 1 37958
0 37960 7 1 2 48854 37959
0 37961 5 1 1 37960
0 37962 7 1 2 37937 37961
0 37963 5 1 1 37962
0 37964 7 1 2 48704 37963
0 37965 5 1 1 37964
0 37966 7 1 2 54358 66652
0 37967 7 1 2 59428 37966
0 37968 5 1 1 37967
0 37969 7 1 2 37965 37968
0 37970 5 1 1 37969
0 37971 7 1 2 67947 37970
0 37972 5 1 1 37971
0 37973 7 1 2 37933 37972
0 37974 5 1 1 37973
0 37975 7 1 2 44979 37974
0 37976 5 1 1 37975
0 37977 7 1 2 14985 18696
0 37978 5 2 1 37977
0 37979 7 3 2 61254 68276
0 37980 7 1 2 64406 70127
0 37981 7 1 2 71527 37980
0 37982 7 1 2 71525 37981
0 37983 5 1 1 37982
0 37984 7 1 2 37976 37983
0 37985 5 1 1 37984
0 37986 7 1 2 54812 37985
0 37987 5 1 1 37986
0 37988 7 1 2 63712 70053
0 37989 5 4 1 37988
0 37990 7 1 2 57516 71530
0 37991 5 1 1 37990
0 37992 7 1 2 50024 53657
0 37993 7 1 2 65611 37992
0 37994 5 1 1 37993
0 37995 7 1 2 37991 37994
0 37996 5 1 1 37995
0 37997 7 1 2 45645 37996
0 37998 5 1 1 37997
0 37999 7 1 2 54746 66653
0 38000 7 1 2 65616 37999
0 38001 5 1 1 38000
0 38002 7 1 2 37998 38001
0 38003 5 1 1 38002
0 38004 7 1 2 47697 38003
0 38005 5 1 1 38004
0 38006 7 1 2 55820 67313
0 38007 5 1 1 38006
0 38008 7 1 2 38005 38007
0 38009 5 1 1 38008
0 38010 7 1 2 53936 38009
0 38011 5 1 1 38010
0 38012 7 1 2 51736 70346
0 38013 5 1 1 38012
0 38014 7 1 2 51543 62450
0 38015 5 2 1 38014
0 38016 7 1 2 58169 59818
0 38017 7 1 2 71534 38016
0 38018 5 1 1 38017
0 38019 7 1 2 38013 38018
0 38020 5 1 1 38019
0 38021 7 1 2 53887 38020
0 38022 5 1 1 38021
0 38023 7 1 2 58552 36950
0 38024 5 1 1 38023
0 38025 7 1 2 44980 63760
0 38026 7 1 2 60015 38025
0 38027 7 1 2 38024 38026
0 38028 5 1 1 38027
0 38029 7 1 2 38022 38028
0 38030 7 1 2 38011 38029
0 38031 5 1 1 38030
0 38032 7 1 2 65974 38031
0 38033 5 1 1 38032
0 38034 7 1 2 65612 67383
0 38035 5 1 1 38034
0 38036 7 1 2 55821 63196
0 38037 5 1 1 38036
0 38038 7 1 2 52907 67897
0 38039 5 1 1 38038
0 38040 7 1 2 66953 38039
0 38041 5 1 1 38040
0 38042 7 1 2 50115 38041
0 38043 5 1 1 38042
0 38044 7 1 2 38037 38043
0 38045 7 1 2 38035 38044
0 38046 5 1 1 38045
0 38047 7 1 2 53937 38046
0 38048 5 1 1 38047
0 38049 7 1 2 48705 69621
0 38050 5 1 1 38049
0 38051 7 1 2 49824 62339
0 38052 5 1 1 38051
0 38053 7 1 2 38050 38052
0 38054 5 1 1 38053
0 38055 7 1 2 51187 38054
0 38056 5 1 1 38055
0 38057 7 1 2 52463 58854
0 38058 5 1 1 38057
0 38059 7 1 2 38056 38058
0 38060 5 1 1 38059
0 38061 7 1 2 66950 38060
0 38062 5 1 1 38061
0 38063 7 1 2 53938 67898
0 38064 7 1 2 71448 38063
0 38065 5 1 1 38064
0 38066 7 1 2 38062 38065
0 38067 5 1 1 38066
0 38068 7 1 2 45502 38067
0 38069 5 1 1 38068
0 38070 7 1 2 38048 38069
0 38071 5 1 1 38070
0 38072 7 1 2 42085 38071
0 38073 5 1 1 38072
0 38074 7 1 2 51410 67653
0 38075 5 1 1 38074
0 38076 7 2 2 53635 55429
0 38077 7 1 2 50884 71536
0 38078 5 1 1 38077
0 38079 7 1 2 54465 58768
0 38080 5 1 1 38079
0 38081 7 1 2 38078 38080
0 38082 5 1 1 38081
0 38083 7 1 2 51086 38082
0 38084 5 1 1 38083
0 38085 7 1 2 38075 38084
0 38086 7 2 2 47461 55822
0 38087 7 1 2 53636 71538
0 38088 5 1 1 38087
0 38089 7 2 2 53658 55713
0 38090 5 1 1 71540
0 38091 7 1 2 46559 71541
0 38092 5 1 1 38091
0 38093 7 1 2 38088 38092
0 38094 5 1 1 38093
0 38095 7 1 2 50025 38094
0 38096 5 1 1 38095
0 38097 7 1 2 38090 37835
0 38098 5 1 1 38097
0 38099 7 1 2 57102 13133
0 38100 5 1 1 38099
0 38101 7 1 2 38098 38100
0 38102 5 1 1 38101
0 38103 7 1 2 38096 38102
0 38104 7 1 2 38085 38103
0 38105 5 1 1 38104
0 38106 7 1 2 53939 59578
0 38107 7 1 2 38105 38106
0 38108 5 1 1 38107
0 38109 7 1 2 38073 38108
0 38110 5 1 1 38109
0 38111 7 1 2 65776 38110
0 38112 5 1 1 38111
0 38113 7 1 2 44498 38112
0 38114 7 1 2 38033 38113
0 38115 5 1 1 38114
0 38116 7 1 2 57301 61255
0 38117 7 1 2 63197 38116
0 38118 5 1 1 38117
0 38119 7 1 2 63899 70440
0 38120 7 1 2 71514 38119
0 38121 5 1 1 38120
0 38122 7 1 2 38118 38121
0 38123 5 1 1 38122
0 38124 7 1 2 48855 38123
0 38125 5 1 1 38124
0 38126 7 1 2 55430 69373
0 38127 7 1 2 56204 38126
0 38128 5 1 1 38127
0 38129 7 1 2 53548 57276
0 38130 7 1 2 70353 38129
0 38131 5 1 1 38130
0 38132 7 1 2 38128 38131
0 38133 5 1 1 38132
0 38134 7 1 2 46560 38133
0 38135 5 1 1 38134
0 38136 7 2 2 52467 60187
0 38137 7 2 2 55769 71542
0 38138 7 1 2 59631 71544
0 38139 5 1 1 38138
0 38140 7 1 2 38135 38139
0 38141 7 1 2 38125 38140
0 38142 5 1 1 38141
0 38143 7 1 2 46764 38142
0 38144 5 1 1 38143
0 38145 7 2 2 43395 71545
0 38146 7 1 2 56109 71546
0 38147 5 1 1 38146
0 38148 7 1 2 62951 71547
0 38149 5 1 1 38148
0 38150 7 1 2 55668 65658
0 38151 7 1 2 70889 38150
0 38152 7 1 2 63269 38151
0 38153 5 1 1 38152
0 38154 7 1 2 38149 38153
0 38155 5 1 1 38154
0 38156 7 1 2 45322 38155
0 38157 5 1 1 38156
0 38158 7 1 2 38147 38157
0 38159 7 1 2 38144 38158
0 38160 5 1 1 38159
0 38161 7 1 2 46098 38160
0 38162 5 1 1 38161
0 38163 7 1 2 55806 63238
0 38164 7 1 2 54662 38163
0 38165 7 1 2 71531 38164
0 38166 5 1 1 38165
0 38167 7 1 2 38162 38166
0 38168 5 1 1 38167
0 38169 7 1 2 45646 38168
0 38170 5 1 1 38169
0 38171 7 1 2 54747 56047
0 38172 7 1 2 71543 38171
0 38173 7 1 2 71376 38172
0 38174 5 1 1 38173
0 38175 7 1 2 38170 38174
0 38176 5 1 1 38175
0 38177 7 1 2 65777 38176
0 38178 5 1 1 38177
0 38179 7 1 2 63106 65643
0 38180 5 1 1 38179
0 38181 7 1 2 66954 38180
0 38182 5 1 1 38181
0 38183 7 1 2 47462 38182
0 38184 5 1 1 38183
0 38185 7 2 2 47925 52717
0 38186 7 1 2 69100 71548
0 38187 5 1 1 38186
0 38188 7 1 2 38184 38187
0 38189 5 1 1 38188
0 38190 7 1 2 51806 38189
0 38191 5 1 1 38190
0 38192 7 1 2 67899 70554
0 38193 5 1 1 38192
0 38194 7 1 2 66955 38193
0 38195 5 1 1 38194
0 38196 7 1 2 50278 38195
0 38197 5 1 1 38196
0 38198 7 1 2 46765 58014
0 38199 7 1 2 58272 38198
0 38200 7 1 2 70348 38199
0 38201 5 1 1 38200
0 38202 7 1 2 38197 38201
0 38203 5 1 1 38202
0 38204 7 1 2 46561 38203
0 38205 5 1 1 38204
0 38206 7 1 2 63558 66951
0 38207 5 1 1 38206
0 38208 7 1 2 38205 38207
0 38209 7 1 2 38191 38208
0 38210 5 1 1 38209
0 38211 7 1 2 45647 38210
0 38212 5 1 1 38211
0 38213 7 1 2 57517 64066
0 38214 5 1 1 38213
0 38215 7 1 2 53659 64241
0 38216 5 2 1 38215
0 38217 7 1 2 38214 71550
0 38218 5 1 1 38217
0 38219 7 1 2 51040 38218
0 38220 5 1 1 38219
0 38221 7 1 2 46766 71537
0 38222 5 1 1 38221
0 38223 7 1 2 71551 38222
0 38224 5 1 1 38223
0 38225 7 1 2 45323 38224
0 38226 5 1 1 38225
0 38227 7 1 2 38220 38226
0 38228 5 1 1 38227
0 38229 7 1 2 59378 38228
0 38230 5 1 1 38229
0 38231 7 1 2 38212 38230
0 38232 5 1 1 38231
0 38233 7 1 2 65975 38232
0 38234 5 1 1 38233
0 38235 7 2 2 51454 54509
0 38236 7 1 2 53660 63410
0 38237 7 1 2 71552 38236
0 38238 5 1 1 38237
0 38239 7 1 2 38234 38238
0 38240 5 1 1 38239
0 38241 7 1 2 53940 38240
0 38242 5 1 1 38241
0 38243 7 1 2 47821 38242
0 38244 7 1 2 38178 38243
0 38245 5 1 1 38244
0 38246 7 1 2 46340 38245
0 38247 7 1 2 38115 38246
0 38248 5 1 1 38247
0 38249 7 1 2 37987 38248
0 38250 7 1 2 37910 38249
0 38251 5 1 1 38250
0 38252 7 1 2 70332 38251
0 38253 5 1 1 38252
0 38254 7 1 2 55714 57777
0 38255 5 1 1 38254
0 38256 7 1 2 71441 38255
0 38257 5 1 1 38256
0 38258 7 1 2 49765 38257
0 38259 5 1 1 38258
0 38260 7 1 2 50175 55720
0 38261 5 1 1 38260
0 38262 7 1 2 57153 71461
0 38263 5 1 1 38262
0 38264 7 1 2 38261 38263
0 38265 7 1 2 38259 38264
0 38266 5 1 1 38265
0 38267 7 1 2 43396 38266
0 38268 5 1 1 38267
0 38269 7 2 2 50639 61918
0 38270 7 1 2 57801 71554
0 38271 5 1 1 38270
0 38272 7 1 2 51687 52908
0 38273 5 1 1 38272
0 38274 7 1 2 28524 38273
0 38275 5 1 1 38274
0 38276 7 1 2 50805 38275
0 38277 5 1 1 38276
0 38278 7 1 2 38271 38277
0 38279 7 1 2 38268 38278
0 38280 5 1 1 38279
0 38281 7 1 2 65778 38280
0 38282 5 2 1 38281
0 38283 7 1 2 51688 71532
0 38284 5 1 1 38283
0 38285 7 1 2 65608 38284
0 38286 5 1 1 38285
0 38287 7 1 2 65976 38286
0 38288 5 1 1 38287
0 38289 7 1 2 71556 38288
0 38290 5 1 1 38289
0 38291 7 1 2 62542 38290
0 38292 5 1 1 38291
0 38293 7 1 2 50026 56965
0 38294 5 1 1 38293
0 38295 7 1 2 51812 38294
0 38296 5 1 1 38295
0 38297 7 1 2 65977 38296
0 38298 5 1 1 38297
0 38299 7 1 2 70355 71433
0 38300 5 1 1 38299
0 38301 7 1 2 38298 38300
0 38302 5 1 1 38301
0 38303 7 1 2 43171 38302
0 38304 5 1 1 38303
0 38305 7 1 2 51620 71252
0 38306 5 1 1 38305
0 38307 7 1 2 38304 38306
0 38308 5 1 1 38307
0 38309 7 1 2 50575 60478
0 38310 7 1 2 38308 38309
0 38311 5 1 1 38310
0 38312 7 1 2 38292 38311
0 38313 5 1 1 38312
0 38314 7 1 2 70298 38313
0 38315 5 1 1 38314
0 38316 7 1 2 63346 71553
0 38317 5 1 1 38316
0 38318 7 1 2 51689 65145
0 38319 5 1 1 38318
0 38320 7 1 2 57566 71401
0 38321 5 1 1 38320
0 38322 7 1 2 38319 38321
0 38323 5 1 1 38322
0 38324 7 1 2 65978 38323
0 38325 5 1 1 38324
0 38326 7 1 2 38317 38325
0 38327 5 1 1 38326
0 38328 7 1 2 60479 38327
0 38329 5 1 1 38328
0 38330 7 1 2 55727 37149
0 38331 5 1 1 38330
0 38332 7 2 2 66029 38331
0 38333 7 1 2 62543 71558
0 38334 5 1 1 38333
0 38335 7 1 2 38329 38334
0 38336 5 1 1 38335
0 38337 7 1 2 70517 38336
0 38338 5 1 1 38337
0 38339 7 1 2 38315 38338
0 38340 5 1 1 38339
0 38341 7 1 2 46099 38340
0 38342 5 1 1 38341
0 38343 7 1 2 62722 67525
0 38344 7 1 2 69487 38343
0 38345 7 1 2 62340 71486
0 38346 7 1 2 38344 38345
0 38347 5 2 1 38346
0 38348 7 1 2 38342 71560
0 38349 5 1 1 38348
0 38350 7 1 2 53919 38349
0 38351 5 1 1 38350
0 38352 7 1 2 51690 59043
0 38353 5 1 1 38352
0 38354 7 1 2 16850 38353
0 38355 5 1 1 38354
0 38356 7 1 2 47463 38355
0 38357 5 1 1 38356
0 38358 7 1 2 51621 55541
0 38359 7 1 2 58424 38358
0 38360 7 1 2 60709 38359
0 38361 5 1 1 38360
0 38362 7 1 2 38357 38361
0 38363 5 1 1 38362
0 38364 7 1 2 45324 38363
0 38365 5 1 1 38364
0 38366 7 2 2 50027 69600
0 38367 5 2 1 71562
0 38368 7 1 2 51622 71563
0 38369 5 1 1 38368
0 38370 7 1 2 51411 71164
0 38371 5 1 1 38370
0 38372 7 1 2 2601 55728
0 38373 5 1 1 38372
0 38374 7 1 2 57091 38373
0 38375 5 1 1 38374
0 38376 7 1 2 38371 38375
0 38377 5 1 1 38376
0 38378 7 1 2 46767 38377
0 38379 5 1 1 38378
0 38380 7 1 2 38369 38379
0 38381 7 1 2 38365 38380
0 38382 5 1 1 38381
0 38383 7 1 2 65979 38382
0 38384 5 1 1 38383
0 38385 7 1 2 71557 38384
0 38386 5 1 1 38385
0 38387 7 1 2 53204 38386
0 38388 5 1 1 38387
0 38389 7 1 2 57103 57830
0 38390 5 1 1 38389
0 38391 7 1 2 45503 38390
0 38392 5 1 1 38391
0 38393 7 2 2 45325 50133
0 38394 7 1 2 49555 71566
0 38395 5 1 1 38394
0 38396 7 1 2 38392 38395
0 38397 5 1 1 38396
0 38398 7 1 2 51623 61879
0 38399 7 1 2 64665 38398
0 38400 7 1 2 38397 38399
0 38401 5 1 1 38400
0 38402 7 1 2 38388 38401
0 38403 5 1 1 38402
0 38404 7 1 2 70299 38403
0 38405 5 1 1 38404
0 38406 7 1 2 51188 71435
0 38407 5 1 1 38406
0 38408 7 1 2 47150 64556
0 38409 5 1 1 38408
0 38410 7 1 2 50176 67920
0 38411 5 1 1 38410
0 38412 7 1 2 38409 38411
0 38413 5 1 1 38412
0 38414 7 1 2 51624 66030
0 38415 7 1 2 38413 38414
0 38416 5 1 1 38415
0 38417 7 1 2 38407 38416
0 38418 5 1 1 38417
0 38419 7 1 2 49718 38418
0 38420 5 1 1 38419
0 38421 7 1 2 53205 71559
0 38422 5 1 1 38421
0 38423 7 2 2 57749 65625
0 38424 7 1 2 49308 55142
0 38425 7 1 2 69035 38424
0 38426 7 1 2 71568 38425
0 38427 5 1 1 38426
0 38428 7 1 2 38422 38427
0 38429 7 1 2 38420 38428
0 38430 5 1 1 38429
0 38431 7 1 2 70518 38430
0 38432 5 1 1 38431
0 38433 7 1 2 38405 38432
0 38434 5 1 1 38433
0 38435 7 1 2 62544 38434
0 38436 5 1 1 38435
0 38437 7 2 2 63095 64557
0 38438 7 1 2 66223 71570
0 38439 5 1 1 38438
0 38440 7 1 2 44272 70546
0 38441 5 1 1 38440
0 38442 7 1 2 38439 38441
0 38443 5 1 1 38442
0 38444 7 1 2 47464 38443
0 38445 5 1 1 38444
0 38446 7 1 2 52718 59607
0 38447 7 1 2 69422 38446
0 38448 5 1 1 38447
0 38449 7 1 2 38445 38448
0 38450 5 1 1 38449
0 38451 7 1 2 65980 38450
0 38452 5 1 1 38451
0 38453 7 1 2 70046 70300
0 38454 5 1 1 38453
0 38455 7 1 2 70551 38454
0 38456 5 1 1 38455
0 38457 7 1 2 45326 38456
0 38458 5 1 1 38457
0 38459 7 1 2 60057 66363
0 38460 7 1 2 51737 38459
0 38461 5 1 1 38460
0 38462 7 1 2 38458 38461
0 38463 5 1 1 38462
0 38464 7 1 2 65779 38463
0 38465 5 1 1 38464
0 38466 7 1 2 38452 38465
0 38467 5 1 1 38466
0 38468 7 1 2 51625 38467
0 38469 5 1 1 38468
0 38470 7 1 2 65981 70616
0 38471 5 1 1 38470
0 38472 7 1 2 44273 61467
0 38473 7 1 2 66420 38472
0 38474 7 1 2 70521 38473
0 38475 5 1 1 38474
0 38476 7 1 2 38471 38475
0 38477 5 1 1 38476
0 38478 7 1 2 43397 38477
0 38479 5 1 1 38478
0 38480 7 1 2 56359 59214
0 38481 7 1 2 69281 38480
0 38482 7 1 2 71269 38481
0 38483 5 1 1 38482
0 38484 7 1 2 38479 38483
0 38485 5 1 1 38484
0 38486 7 1 2 45327 38485
0 38487 5 1 1 38486
0 38488 7 1 2 63457 66074
0 38489 7 1 2 62400 38488
0 38490 7 1 2 70621 38489
0 38491 5 1 1 38490
0 38492 7 1 2 38487 38491
0 38493 5 1 1 38492
0 38494 7 1 2 51691 38493
0 38495 5 1 1 38494
0 38496 7 1 2 38469 38495
0 38497 5 1 1 38496
0 38498 7 1 2 53206 38497
0 38499 5 1 1 38498
0 38500 7 1 2 56058 65780
0 38501 7 1 2 70312 70764
0 38502 7 1 2 38500 38501
0 38503 7 1 2 70050 38502
0 38504 5 1 1 38503
0 38505 7 1 2 38499 38504
0 38506 5 1 1 38505
0 38507 7 1 2 60480 38506
0 38508 5 1 1 38507
0 38509 7 1 2 38436 38508
0 38510 5 1 1 38509
0 38511 7 1 2 44981 38510
0 38512 5 1 1 38511
0 38513 7 1 2 48706 67135
0 38514 7 1 2 70618 38513
0 38515 5 1 1 38514
0 38516 7 1 2 70552 38515
0 38517 5 1 1 38516
0 38518 7 1 2 59716 62545
0 38519 7 1 2 71379 38518
0 38520 5 1 1 38519
0 38521 7 1 2 50215 51692
0 38522 7 1 2 68277 38521
0 38523 7 1 2 70384 70637
0 38524 7 1 2 38522 38523
0 38525 5 1 1 38524
0 38526 7 1 2 38520 38525
0 38527 5 1 1 38526
0 38528 7 1 2 38517 38527
0 38529 5 1 1 38528
0 38530 7 1 2 56520 64695
0 38531 7 1 2 70619 71490
0 38532 7 1 2 38530 38531
0 38533 7 1 2 71535 38532
0 38534 5 1 1 38533
0 38535 7 1 2 55298 69978
0 38536 5 1 1 38535
0 38537 7 1 2 46768 38536
0 38538 5 1 1 38537
0 38539 7 1 2 71374 38538
0 38540 5 1 1 38539
0 38541 7 1 2 68534 38540
0 38542 5 1 1 38541
0 38543 7 1 2 64700 71506
0 38544 5 1 1 38543
0 38545 7 1 2 38542 38544
0 38546 5 1 1 38545
0 38547 7 1 2 53561 70923
0 38548 7 1 2 38546 38547
0 38549 5 1 1 38548
0 38550 7 1 2 38534 38549
0 38551 5 1 1 38550
0 38552 7 1 2 47151 38551
0 38553 5 1 1 38552
0 38554 7 1 2 71561 38553
0 38555 5 1 1 38554
0 38556 7 1 2 52436 38555
0 38557 5 1 1 38556
0 38558 7 1 2 38529 38557
0 38559 7 1 2 38512 38558
0 38560 7 1 2 38351 38559
0 38561 5 1 1 38560
0 38562 7 1 2 46341 38561
0 38563 5 1 1 38562
0 38564 7 1 2 38253 38563
0 38565 7 1 2 37667 38564
0 38566 5 1 1 38565
0 38567 7 1 2 48158 38566
0 38568 5 1 1 38567
0 38569 7 2 2 55628 65455
0 38570 7 1 2 51320 71572
0 38571 5 1 1 38570
0 38572 7 2 2 48856 70908
0 38573 7 1 2 57890 67712
0 38574 7 1 2 71574 38573
0 38575 5 1 1 38574
0 38576 7 1 2 38571 38575
0 38577 5 1 1 38576
0 38578 7 1 2 48307 38577
0 38579 5 1 1 38578
0 38580 7 2 2 48159 59717
0 38581 7 1 2 71576 71573
0 38582 5 1 1 38581
0 38583 7 1 2 38579 38582
0 38584 5 1 1 38583
0 38585 7 1 2 47465 38584
0 38586 5 1 1 38585
0 38587 7 1 2 42631 56448
0 38588 5 2 1 38587
0 38589 7 1 2 53920 54084
0 38590 5 1 1 38589
0 38591 7 1 2 71578 38590
0 38592 5 7 1 38591
0 38593 7 1 2 52719 62236
0 38594 7 1 2 71580 38593
0 38595 5 1 1 38594
0 38596 7 1 2 38586 38595
0 38597 5 1 1 38596
0 38598 7 1 2 42086 38597
0 38599 5 1 1 38598
0 38600 7 1 2 56033 64942
0 38601 7 1 2 71581 38600
0 38602 5 1 1 38601
0 38603 7 1 2 38599 38602
0 38604 5 1 1 38603
0 38605 7 1 2 44366 38604
0 38606 5 1 1 38605
0 38607 7 1 2 49010 61086
0 38608 7 1 2 61890 38607
0 38609 7 1 2 71582 38608
0 38610 5 1 1 38609
0 38611 7 1 2 38606 38610
0 38612 5 1 1 38611
0 38613 7 1 2 70111 38612
0 38614 5 1 1 38613
0 38615 7 1 2 55919 64818
0 38616 5 1 1 38615
0 38617 7 1 2 57535 70667
0 38618 5 1 1 38617
0 38619 7 1 2 38616 38618
0 38620 5 2 1 38619
0 38621 7 1 2 45648 71587
0 38622 5 1 1 38621
0 38623 7 1 2 58092 64819
0 38624 5 1 1 38623
0 38625 7 1 2 38622 38624
0 38626 5 1 1 38625
0 38627 7 1 2 43777 68703
0 38628 5 1 1 38627
0 38629 7 1 2 71579 38628
0 38630 5 1 1 38629
0 38631 7 1 2 38626 38630
0 38632 5 1 1 38631
0 38633 7 1 2 50207 51303
0 38634 7 4 2 45328 58874
0 38635 7 1 2 54813 71589
0 38636 7 1 2 38633 38635
0 38637 5 1 1 38636
0 38638 7 1 2 38632 38637
0 38639 5 1 1 38638
0 38640 7 1 2 46562 38639
0 38641 5 1 1 38640
0 38642 7 1 2 48160 48972
0 38643 7 1 2 55502 38642
0 38644 7 1 2 63332 66713
0 38645 7 1 2 38643 38644
0 38646 5 1 1 38645
0 38647 7 1 2 38641 38646
0 38648 5 1 1 38647
0 38649 7 1 2 69089 38648
0 38650 5 1 1 38649
0 38651 7 1 2 38614 38650
0 38652 5 1 1 38651
0 38653 7 1 2 53615 38652
0 38654 5 1 1 38653
0 38655 7 1 2 66528 68138
0 38656 5 2 1 38655
0 38657 7 2 2 61811 64631
0 38658 7 1 2 47822 52272
0 38659 7 1 2 60121 38658
0 38660 7 1 2 71595 38659
0 38661 5 1 1 38660
0 38662 7 1 2 64485 70767
0 38663 7 1 2 67210 38662
0 38664 7 1 2 63615 38663
0 38665 5 1 1 38664
0 38666 7 1 2 38661 38665
0 38667 5 1 1 38666
0 38668 7 1 2 48308 38667
0 38669 5 1 1 38668
0 38670 7 1 2 43778 69724
0 38671 7 1 2 71520 38670
0 38672 7 1 2 71596 38671
0 38673 5 1 1 38672
0 38674 7 1 2 38669 38673
0 38675 5 1 1 38674
0 38676 7 1 2 71593 38675
0 38677 5 1 1 38676
0 38678 7 1 2 64425 70663
0 38679 5 1 1 38678
0 38680 7 1 2 49825 54138
0 38681 7 1 2 66494 38680
0 38682 5 1 1 38681
0 38683 7 1 2 38679 38682
0 38684 5 1 1 38683
0 38685 7 1 2 44835 38684
0 38686 5 1 1 38685
0 38687 7 1 2 57698 64419
0 38688 7 1 2 66495 38687
0 38689 5 1 1 38688
0 38690 7 1 2 38686 38689
0 38691 5 1 1 38690
0 38692 7 1 2 42632 38691
0 38693 5 1 1 38692
0 38694 7 1 2 56734 65647
0 38695 7 1 2 71504 38694
0 38696 5 1 1 38695
0 38697 7 1 2 38693 38696
0 38698 5 1 1 38697
0 38699 7 1 2 69865 38698
0 38700 5 1 1 38699
0 38701 7 1 2 38677 38700
0 38702 5 1 1 38701
0 38703 7 1 2 43172 38702
0 38704 5 1 1 38703
0 38705 7 1 2 56009 64004
0 38706 5 1 1 38705
0 38707 7 1 2 56045 63837
0 38708 5 1 1 38707
0 38709 7 1 2 38706 38708
0 38710 5 1 1 38709
0 38711 7 2 2 53046 70697
0 38712 7 1 2 38710 71597
0 38713 5 1 1 38712
0 38714 7 1 2 52794 57891
0 38715 7 1 2 63616 38714
0 38716 7 1 2 71594 38715
0 38717 5 1 1 38716
0 38718 7 1 2 38713 38717
0 38719 5 1 1 38718
0 38720 7 1 2 42087 38719
0 38721 5 1 1 38720
0 38722 7 1 2 68700 70848
0 38723 7 1 2 71598 38722
0 38724 5 1 1 38723
0 38725 7 1 2 38721 38724
0 38726 5 1 1 38725
0 38727 7 1 2 44367 38726
0 38728 5 1 1 38727
0 38729 7 1 2 56731 58629
0 38730 5 1 1 38729
0 38731 7 1 2 68686 38730
0 38732 5 2 1 38731
0 38733 7 1 2 42349 66758
0 38734 7 1 2 70006 38733
0 38735 7 1 2 71599 38734
0 38736 5 1 1 38735
0 38737 7 1 2 38728 38736
0 38738 5 1 1 38737
0 38739 7 1 2 56449 38738
0 38740 5 1 1 38739
0 38741 7 1 2 66489 71528
0 38742 5 1 1 38741
0 38743 7 1 2 53747 70660
0 38744 5 1 1 38743
0 38745 7 1 2 38742 38744
0 38746 5 1 1 38745
0 38747 7 1 2 49766 38746
0 38748 5 1 1 38747
0 38749 7 1 2 64309 71529
0 38750 5 1 1 38749
0 38751 7 1 2 45504 70661
0 38752 5 1 1 38751
0 38753 7 1 2 38750 38752
0 38754 5 1 1 38753
0 38755 7 1 2 53036 38754
0 38756 5 1 1 38755
0 38757 7 1 2 38748 38756
0 38758 5 1 1 38757
0 38759 7 1 2 54085 38758
0 38760 5 1 1 38759
0 38761 7 1 2 53037 56303
0 38762 5 1 1 38761
0 38763 7 1 2 49783 50908
0 38764 5 1 1 38763
0 38765 7 1 2 38762 38764
0 38766 5 1 1 38765
0 38767 7 1 2 55658 67941
0 38768 7 1 2 38766 38767
0 38769 5 1 1 38768
0 38770 7 1 2 38760 38769
0 38771 5 1 1 38770
0 38772 7 1 2 69897 38771
0 38773 5 1 1 38772
0 38774 7 1 2 49309 59983
0 38775 7 1 2 63756 38774
0 38776 7 1 2 68388 68659
0 38777 7 1 2 71465 38776
0 38778 7 1 2 38775 38777
0 38779 5 1 1 38778
0 38780 7 1 2 52169 63239
0 38781 7 1 2 62601 38780
0 38782 7 1 2 66522 70898
0 38783 7 1 2 38781 38782
0 38784 7 1 2 58107 38783
0 38785 5 1 1 38784
0 38786 7 1 2 38779 38785
0 38787 7 1 2 38773 38786
0 38788 7 1 2 38740 38787
0 38789 7 1 2 38704 38788
0 38790 7 1 2 38654 38789
0 38791 5 1 1 38790
0 38792 7 1 2 66283 38791
0 38793 5 1 1 38792
0 38794 7 1 2 46563 70627
0 38795 5 1 1 38794
0 38796 7 1 2 1532 38795
0 38797 5 1 1 38796
0 38798 7 1 2 49767 38797
0 38799 5 1 1 38798
0 38800 7 1 2 5166 70629
0 38801 5 1 1 38800
0 38802 7 1 2 53038 38801
0 38803 5 1 1 38802
0 38804 7 1 2 38799 38803
0 38805 5 1 1 38804
0 38806 7 1 2 65781 38805
0 38807 5 1 1 38806
0 38808 7 1 2 53039 64310
0 38809 5 1 1 38808
0 38810 7 1 2 49768 66490
0 38811 5 1 1 38810
0 38812 7 1 2 38809 38811
0 38813 5 1 1 38812
0 38814 7 2 2 48038 38813
0 38815 7 1 2 51321 71601
0 38816 5 1 1 38815
0 38817 7 1 2 38807 38816
0 38818 5 2 1 38817
0 38819 7 1 2 48309 71603
0 38820 5 1 1 38819
0 38821 7 1 2 71602 71577
0 38822 5 1 1 38821
0 38823 7 1 2 38820 38822
0 38824 5 1 1 38823
0 38825 7 1 2 51952 38824
0 38826 5 1 1 38825
0 38827 7 1 2 61441 64056
0 38828 7 1 2 53047 38827
0 38829 7 1 2 71583 38828
0 38830 5 1 1 38829
0 38831 7 1 2 38826 38830
0 38832 5 1 1 38831
0 38833 7 1 2 53694 71494
0 38834 5 1 1 38833
0 38835 7 1 2 44368 69334
0 38836 5 1 1 38835
0 38837 7 1 2 38834 38836
0 38838 5 1 1 38837
0 38839 7 1 2 38832 38838
0 38840 5 1 1 38839
0 38841 7 1 2 48857 71135
0 38842 5 1 1 38841
0 38843 7 1 2 70749 38842
0 38844 5 1 1 38843
0 38845 7 1 2 53925 38844
0 38846 5 1 1 38845
0 38847 7 2 2 54065 64005
0 38848 7 1 2 50370 53207
0 38849 7 1 2 71605 38848
0 38850 5 1 1 38849
0 38851 7 1 2 38846 38850
0 38852 5 1 1 38851
0 38853 7 1 2 48161 38852
0 38854 5 1 1 38853
0 38855 7 1 2 68252 70635
0 38856 5 1 1 38855
0 38857 7 1 2 38854 38856
0 38858 5 1 1 38857
0 38859 7 1 2 61468 38858
0 38860 5 1 1 38859
0 38861 7 2 2 55659 67111
0 38862 7 1 2 70484 71607
0 38863 5 1 1 38862
0 38864 7 1 2 38860 38863
0 38865 5 1 1 38864
0 38866 7 1 2 45329 38865
0 38867 5 1 1 38866
0 38868 7 2 2 49797 51105
0 38869 5 1 1 71609
0 38870 7 1 2 55715 60410
0 38871 7 1 2 68518 38870
0 38872 7 1 2 71610 38871
0 38873 5 1 1 38872
0 38874 7 1 2 38867 38873
0 38875 5 1 1 38874
0 38876 7 1 2 46342 38875
0 38877 5 1 1 38876
0 38878 7 1 2 65263 66979
0 38879 7 1 2 71600 38878
0 38880 5 1 1 38879
0 38881 7 1 2 55394 70023
0 38882 7 1 2 71033 38881
0 38883 5 1 1 38882
0 38884 7 1 2 38880 38883
0 38885 5 1 1 38884
0 38886 7 1 2 56450 38885
0 38887 5 1 1 38886
0 38888 7 1 2 53921 65982
0 38889 7 1 2 65264 38888
0 38890 5 1 1 38889
0 38891 7 1 2 70758 38890
0 38892 5 1 1 38891
0 38893 7 1 2 64924 38892
0 38894 5 1 1 38893
0 38895 7 2 2 50433 65648
0 38896 7 1 2 71606 71611
0 38897 5 1 1 38896
0 38898 7 1 2 38894 38897
0 38899 5 1 1 38898
0 38900 7 1 2 55259 38899
0 38901 5 1 1 38900
0 38902 7 1 2 38887 38901
0 38903 7 1 2 38877 38902
0 38904 5 1 1 38903
0 38905 7 1 2 58204 71048
0 38906 7 1 2 38904 38905
0 38907 5 1 1 38906
0 38908 7 1 2 38840 38907
0 38909 5 1 1 38908
0 38910 7 1 2 47823 38909
0 38911 5 1 1 38910
0 38912 7 1 2 69986 70692
0 38913 7 1 2 71584 38912
0 38914 5 1 1 38913
0 38915 7 1 2 65782 71585
0 38916 5 1 1 38915
0 38917 7 1 2 48310 70335
0 38918 5 1 1 38917
0 38919 7 1 2 38916 38918
0 38920 5 1 1 38919
0 38921 7 1 2 59316 64820
0 38922 7 1 2 38920 38921
0 38923 5 1 1 38922
0 38924 7 1 2 38914 38923
0 38925 5 2 1 38924
0 38926 7 1 2 66924 71613
0 38927 5 1 1 38926
0 38928 7 1 2 54537 64355
0 38929 7 1 2 68183 38928
0 38930 7 1 2 71608 38929
0 38931 5 1 1 38930
0 38932 7 1 2 38927 38931
0 38933 5 1 1 38932
0 38934 7 1 2 46564 38933
0 38935 5 1 1 38934
0 38936 7 1 2 56446 18867
0 38937 5 1 1 38936
0 38938 7 1 2 57948 67669
0 38939 5 1 1 38938
0 38940 7 1 2 70750 38939
0 38941 5 1 1 38940
0 38942 7 1 2 63617 38941
0 38943 7 1 2 38937 38942
0 38944 5 1 1 38943
0 38945 7 1 2 60247 65251
0 38946 7 1 2 71005 38945
0 38947 7 1 2 71575 38946
0 38948 5 1 1 38947
0 38949 7 1 2 63379 64121
0 38950 7 1 2 69718 38949
0 38951 7 1 2 70987 38950
0 38952 5 1 1 38951
0 38953 7 1 2 38948 38952
0 38954 7 1 2 38944 38953
0 38955 5 1 1 38954
0 38956 7 1 2 71145 38955
0 38957 5 1 1 38956
0 38958 7 1 2 38935 38957
0 38959 5 1 1 38958
0 38960 7 1 2 42088 38959
0 38961 5 1 1 38960
0 38962 7 1 2 59819 70728
0 38963 7 1 2 71614 38962
0 38964 5 1 1 38963
0 38965 7 1 2 38961 38964
0 38966 5 1 1 38965
0 38967 7 1 2 44499 38966
0 38968 5 1 1 38967
0 38969 7 1 2 42350 71498
0 38970 5 1 1 38969
0 38971 7 1 2 71387 38970
0 38972 5 1 1 38971
0 38973 7 1 2 56267 57892
0 38974 7 1 2 38972 38973
0 38975 5 1 1 38974
0 38976 7 1 2 17756 70928
0 38977 5 1 1 38976
0 38978 7 1 2 49769 38977
0 38979 5 1 1 38978
0 38980 7 1 2 53040 65825
0 38981 5 1 1 38980
0 38982 7 1 2 38979 38981
0 38983 5 1 1 38982
0 38984 7 1 2 51158 55629
0 38985 7 1 2 38983 38984
0 38986 5 1 1 38985
0 38987 7 1 2 38975 38986
0 38988 5 1 1 38987
0 38989 7 1 2 44836 38988
0 38990 5 1 1 38989
0 38991 7 1 2 51304 55630
0 38992 7 1 2 66031 38991
0 38993 7 1 2 64943 38992
0 38994 5 1 1 38993
0 38995 7 1 2 38990 38994
0 38996 5 1 1 38995
0 38997 7 1 2 42089 38996
0 38998 5 1 1 38997
0 38999 7 1 2 56034 71604
0 39000 5 1 1 38999
0 39001 7 1 2 38998 39000
0 39002 5 1 1 39001
0 39003 7 1 2 48311 39002
0 39004 5 1 1 39003
0 39005 7 2 2 46864 64105
0 39006 7 2 2 47824 64973
0 39007 7 1 2 71615 71617
0 39008 5 1 1 39007
0 39009 7 1 2 64532 64708
0 39010 7 1 2 70011 39009
0 39011 5 1 1 39010
0 39012 7 1 2 39008 39011
0 39013 5 1 1 39012
0 39014 7 1 2 47152 39013
0 39015 5 1 1 39014
0 39016 7 1 2 59984 63300
0 39017 7 1 2 71618 39016
0 39018 5 1 1 39017
0 39019 7 1 2 39015 39018
0 39020 5 1 1 39019
0 39021 7 1 2 42090 39020
0 39022 5 1 1 39021
0 39023 7 1 2 60880 63126
0 39024 7 1 2 64974 39023
0 39025 5 1 1 39024
0 39026 7 1 2 39022 39025
0 39027 5 1 1 39026
0 39028 7 1 2 51256 39027
0 39029 5 1 1 39028
0 39030 7 1 2 39004 39029
0 39031 5 1 1 39030
0 39032 7 1 2 51865 39031
0 39033 5 1 1 39032
0 39034 7 2 2 57646 65835
0 39035 7 1 2 71162 71619
0 39036 7 1 2 71203 39035
0 39037 7 1 2 71586 39036
0 39038 5 1 1 39037
0 39039 7 1 2 44369 39038
0 39040 7 1 2 39033 39039
0 39041 5 1 1 39040
0 39042 7 1 2 44694 63392
0 39043 7 1 2 71588 39042
0 39044 5 1 1 39043
0 39045 7 1 2 55345 57887
0 39046 7 1 2 68994 39045
0 39047 5 1 1 39046
0 39048 7 1 2 39044 39047
0 39049 5 1 1 39048
0 39050 7 1 2 42633 39049
0 39051 5 1 1 39050
0 39052 7 1 2 45871 55495
0 39053 7 1 2 55631 39052
0 39054 7 1 2 68682 39053
0 39055 5 1 1 39054
0 39056 7 1 2 39051 39055
0 39057 5 1 1 39056
0 39058 7 1 2 60574 39057
0 39059 5 1 1 39058
0 39060 7 1 2 57933 63745
0 39061 7 1 2 68338 68735
0 39062 7 1 2 39060 39061
0 39063 5 1 1 39062
0 39064 7 1 2 39059 39063
0 39065 5 1 1 39064
0 39066 7 1 2 45649 39065
0 39067 5 1 1 39066
0 39068 7 1 2 44695 55403
0 39069 7 1 2 64821 39068
0 39070 7 1 2 65653 69894
0 39071 7 1 2 39069 39070
0 39072 5 1 1 39071
0 39073 7 1 2 39067 39072
0 39074 5 1 1 39073
0 39075 7 1 2 56451 39074
0 39076 5 1 1 39075
0 39077 7 1 2 54402 55831
0 39078 7 1 2 62564 63181
0 39079 7 1 2 39077 39078
0 39080 5 1 1 39079
0 39081 7 1 2 56225 68438
0 39082 5 1 1 39081
0 39083 7 2 2 57949 63393
0 39084 7 1 2 55920 71621
0 39085 5 1 1 39084
0 39086 7 1 2 39082 39085
0 39087 5 1 1 39086
0 39088 7 1 2 45650 39087
0 39089 5 1 1 39088
0 39090 7 1 2 60504 71622
0 39091 5 1 1 39090
0 39092 7 1 2 39089 39091
0 39093 5 1 1 39092
0 39094 7 1 2 50576 54086
0 39095 7 1 2 39093 39094
0 39096 5 1 1 39095
0 39097 7 1 2 39080 39096
0 39098 5 1 1 39097
0 39099 7 1 2 53922 39098
0 39100 5 1 1 39099
0 39101 7 1 2 49826 63380
0 39102 5 1 1 39101
0 39103 7 1 2 38869 39102
0 39104 5 1 1 39103
0 39105 7 1 2 60160 64122
0 39106 7 1 2 62554 39105
0 39107 7 1 2 39104 39106
0 39108 5 1 1 39107
0 39109 7 1 2 61590 62216
0 39110 7 1 2 64386 71466
0 39111 7 1 2 39109 39110
0 39112 5 1 1 39111
0 39113 7 1 2 39108 39112
0 39114 5 1 1 39113
0 39115 7 1 2 45651 39114
0 39116 5 1 1 39115
0 39117 7 1 2 44500 52536
0 39118 7 1 2 61608 39117
0 39119 7 1 2 70880 71616
0 39120 7 1 2 39118 39119
0 39121 5 1 1 39120
0 39122 7 1 2 39116 39121
0 39123 7 1 2 39100 39122
0 39124 5 1 1 39123
0 39125 7 1 2 60575 39124
0 39126 5 1 1 39125
0 39127 7 1 2 45872 50666
0 39128 7 1 2 61030 39127
0 39129 7 1 2 58780 61902
0 39130 7 1 2 39128 39129
0 39131 7 1 2 53926 39130
0 39132 5 1 1 39131
0 39133 7 1 2 47698 39132
0 39134 7 1 2 39126 39133
0 39135 7 1 2 39076 39134
0 39136 5 1 1 39135
0 39137 7 1 2 67034 39136
0 39138 7 1 2 39041 39137
0 39139 5 1 1 39138
0 39140 7 1 2 38968 39139
0 39141 7 1 2 38911 39140
0 39142 7 1 2 38793 39141
0 39143 5 1 1 39142
0 39144 7 1 2 55596 39143
0 39145 5 1 1 39144
0 39146 7 2 2 48312 53208
0 39147 7 1 2 69898 71193
0 39148 5 1 1 39147
0 39149 7 1 2 60498 60788
0 39150 7 1 2 58146 39149
0 39151 5 1 1 39150
0 39152 7 1 2 39148 39151
0 39153 5 1 1 39152
0 39154 7 1 2 48707 39153
0 39155 5 1 1 39154
0 39156 7 1 2 65196 70155
0 39157 5 1 1 39156
0 39158 7 1 2 39155 39157
0 39159 5 2 1 39158
0 39160 7 1 2 71623 71625
0 39161 5 1 1 39160
0 39162 7 1 2 46100 71626
0 39163 5 1 1 39162
0 39164 7 1 2 55413 70034
0 39165 7 1 2 70003 39164
0 39166 7 1 2 65093 39165
0 39167 5 3 1 39166
0 39168 7 1 2 39163 71627
0 39169 5 1 1 39168
0 39170 7 1 2 48313 39169
0 39171 5 1 1 39170
0 39172 7 1 2 59761 71571
0 39173 5 1 1 39172
0 39174 7 1 2 60240 39173
0 39175 5 1 1 39174
0 39176 7 1 2 47466 39175
0 39177 5 1 1 39176
0 39178 7 1 2 59538 71234
0 39179 5 1 1 39178
0 39180 7 1 2 56891 59485
0 39181 7 1 2 68498 39180
0 39182 7 1 2 69092 39181
0 39183 5 1 1 39182
0 39184 7 1 2 39179 39183
0 39185 7 1 2 39177 39184
0 39186 5 1 1 39185
0 39187 7 1 2 46343 39186
0 39188 5 1 1 39187
0 39189 7 1 2 47467 67301
0 39190 7 1 2 69102 39189
0 39191 5 1 1 39190
0 39192 7 1 2 39188 39191
0 39193 5 1 1 39192
0 39194 7 1 2 48314 39193
0 39195 5 1 1 39194
0 39196 7 1 2 53549 64558
0 39197 5 1 1 39196
0 39198 7 1 2 49827 50341
0 39199 5 1 1 39198
0 39200 7 1 2 39197 39199
0 39201 5 1 1 39200
0 39202 7 1 2 59494 39201
0 39203 5 1 1 39202
0 39204 7 1 2 48315 57585
0 39205 5 3 1 39204
0 39206 7 1 2 50895 59027
0 39207 5 1 1 39206
0 39208 7 1 2 49798 39207
0 39209 5 1 1 39208
0 39210 7 1 2 71630 39209
0 39211 5 1 1 39210
0 39212 7 1 2 59539 39211
0 39213 5 1 1 39212
0 39214 7 1 2 39203 39213
0 39215 5 1 1 39214
0 39216 7 1 2 42924 39215
0 39217 5 1 1 39216
0 39218 7 1 2 62044 65254
0 39219 7 1 2 68333 68947
0 39220 7 1 2 39218 39219
0 39221 5 1 1 39220
0 39222 7 1 2 39217 39221
0 39223 7 1 2 39195 39222
0 39224 5 1 1 39223
0 39225 7 1 2 45652 39224
0 39226 5 1 1 39225
0 39227 7 1 2 49799 71189
0 39228 5 1 1 39227
0 39229 7 1 2 48316 64944
0 39230 5 1 1 39229
0 39231 7 1 2 39228 39230
0 39232 5 1 1 39231
0 39233 7 1 2 43398 39232
0 39234 5 1 1 39233
0 39235 7 1 2 44274 64945
0 39236 5 1 1 39235
0 39237 7 1 2 53876 13847
0 39238 5 1 1 39237
0 39239 7 1 2 50806 39238
0 39240 5 1 1 39239
0 39241 7 1 2 39236 39240
0 39242 5 1 1 39241
0 39243 7 1 2 48317 39242
0 39244 5 1 1 39243
0 39245 7 1 2 56732 68959
0 39246 5 1 1 39245
0 39247 7 1 2 71631 39246
0 39248 5 1 1 39247
0 39249 7 1 2 43173 39248
0 39250 5 1 1 39249
0 39251 7 1 2 44275 53550
0 39252 5 1 1 39251
0 39253 7 1 2 71632 39252
0 39254 5 1 1 39253
0 39255 7 1 2 42925 39254
0 39256 5 1 1 39255
0 39257 7 1 2 39250 39256
0 39258 7 1 2 39244 39257
0 39259 7 1 2 39234 39258
0 39260 5 1 1 39259
0 39261 7 1 2 67158 39260
0 39262 5 1 1 39261
0 39263 7 1 2 47825 39262
0 39264 7 1 2 39226 39263
0 39265 5 1 1 39264
0 39266 7 1 2 44276 70683
0 39267 5 1 1 39266
0 39268 7 1 2 54835 64868
0 39269 5 1 1 39268
0 39270 7 1 2 39267 39269
0 39271 5 1 1 39270
0 39272 7 1 2 43399 39271
0 39273 5 1 1 39272
0 39274 7 1 2 56698 59900
0 39275 5 1 1 39274
0 39276 7 1 2 39273 39275
0 39277 5 2 1 39276
0 39278 7 1 2 59495 71633
0 39279 5 1 1 39278
0 39280 7 1 2 48318 59540
0 39281 7 1 2 71425 39280
0 39282 5 1 1 39281
0 39283 7 1 2 39279 39282
0 39284 5 1 1 39283
0 39285 7 1 2 42091 39284
0 39286 5 1 1 39285
0 39287 7 1 2 59583 71634
0 39288 5 1 1 39287
0 39289 7 1 2 44501 39288
0 39290 7 1 2 39286 39289
0 39291 5 1 1 39290
0 39292 7 1 2 42634 39291
0 39293 7 1 2 39265 39292
0 39294 5 1 1 39293
0 39295 7 1 2 39171 39294
0 39296 5 1 1 39295
0 39297 7 1 2 43779 39296
0 39298 5 1 1 39297
0 39299 7 1 2 39161 39298
0 39300 5 1 1 39299
0 39301 7 1 2 66792 39300
0 39302 5 1 1 39301
0 39303 7 1 2 50965 58930
0 39304 5 1 1 39303
0 39305 7 1 2 57972 58435
0 39306 5 1 1 39305
0 39307 7 1 2 39304 39306
0 39308 5 1 1 39307
0 39309 7 1 2 46344 39308
0 39310 5 1 1 39309
0 39311 7 1 2 58666 67198
0 39312 5 1 1 39311
0 39313 7 1 2 39310 39312
0 39314 5 1 1 39313
0 39315 7 1 2 45505 39314
0 39316 5 1 1 39315
0 39317 7 1 2 53435 60585
0 39318 5 1 1 39317
0 39319 7 1 2 18412 39318
0 39320 5 1 1 39319
0 39321 7 1 2 58520 39320
0 39322 5 1 1 39321
0 39323 7 1 2 39316 39322
0 39324 5 1 1 39323
0 39325 7 1 2 70112 39324
0 39326 5 1 1 39325
0 39327 7 1 2 63337 66882
0 39328 7 1 2 60772 39327
0 39329 5 1 1 39328
0 39330 7 1 2 39326 39329
0 39331 5 1 1 39330
0 39332 7 1 2 48319 39331
0 39333 5 1 1 39332
0 39334 7 1 2 69347 71620
0 39335 5 1 1 39334
0 39336 7 2 2 50028 60587
0 39337 7 1 2 70113 71635
0 39338 5 1 1 39337
0 39339 7 1 2 39335 39338
0 39340 5 1 1 39339
0 39341 7 1 2 53436 58230
0 39342 7 1 2 39340 39341
0 39343 5 1 1 39342
0 39344 7 1 2 39333 39343
0 39345 5 1 1 39344
0 39346 7 1 2 43780 39345
0 39347 5 1 1 39346
0 39348 7 1 2 51773 70077
0 39349 5 1 1 39348
0 39350 7 1 2 70071 71041
0 39351 5 1 1 39350
0 39352 7 1 2 39349 39351
0 39353 5 1 1 39352
0 39354 7 1 2 71405 39353
0 39355 5 1 1 39354
0 39356 7 1 2 51572 66990
0 39357 7 1 2 58931 39356
0 39358 5 1 1 39357
0 39359 7 1 2 39355 39358
0 39360 5 1 1 39359
0 39361 7 1 2 71624 39360
0 39362 5 1 1 39361
0 39363 7 1 2 39347 39362
0 39364 5 1 1 39363
0 39365 7 1 2 42092 39364
0 39366 5 1 1 39365
0 39367 7 1 2 52138 68028
0 39368 5 1 1 39367
0 39369 7 1 2 52304 71309
0 39370 5 1 1 39369
0 39371 7 1 2 39368 39370
0 39372 5 1 1 39371
0 39373 7 1 2 56035 70114
0 39374 7 1 2 39372 39373
0 39375 5 1 1 39374
0 39376 7 1 2 39366 39375
0 39377 5 1 1 39376
0 39378 7 1 2 48708 39377
0 39379 5 1 1 39378
0 39380 7 1 2 50577 71526
0 39381 5 1 1 39380
0 39382 7 1 2 50282 51785
0 39383 5 1 1 39382
0 39384 7 1 2 51041 39383
0 39385 5 1 1 39384
0 39386 7 1 2 45330 51807
0 39387 5 1 1 39386
0 39388 7 1 2 49248 39387
0 39389 7 1 2 39385 39388
0 39390 5 1 1 39389
0 39391 7 1 2 46345 39390
0 39392 5 1 1 39391
0 39393 7 1 2 39381 39392
0 39394 5 1 1 39393
0 39395 7 1 2 71178 39394
0 39396 5 1 1 39395
0 39397 7 2 2 50116 53048
0 39398 5 1 1 71637
0 39399 7 1 2 51718 71638
0 39400 5 1 1 39399
0 39401 7 1 2 7445 39400
0 39402 5 1 1 39401
0 39403 7 1 2 54510 67632
0 39404 7 1 2 39402 39403
0 39405 5 1 1 39404
0 39406 7 1 2 39396 39405
0 39407 5 1 1 39406
0 39408 7 1 2 47826 39407
0 39409 5 1 1 39408
0 39410 7 1 2 51042 56741
0 39411 5 1 1 39410
0 39412 7 1 2 14418 39411
0 39413 5 1 1 39412
0 39414 7 1 2 63324 68339
0 39415 7 1 2 39413 39414
0 39416 5 1 1 39415
0 39417 7 1 2 39409 39416
0 39418 5 1 1 39417
0 39419 7 1 2 42635 39418
0 39420 5 1 1 39419
0 39421 7 1 2 56862 62221
0 39422 7 1 2 62664 39421
0 39423 7 1 2 63254 39422
0 39424 5 1 1 39423
0 39425 7 1 2 39420 39424
0 39426 5 1 1 39425
0 39427 7 1 2 52139 39426
0 39428 5 1 1 39427
0 39429 7 1 2 44370 39428
0 39430 7 1 2 39379 39429
0 39431 5 1 1 39430
0 39432 7 1 2 56755 60588
0 39433 5 1 1 39432
0 39434 7 1 2 55632 56647
0 39435 5 1 1 39434
0 39436 7 1 2 39433 39435
0 39437 5 1 1 39436
0 39438 7 1 2 66411 39437
0 39439 5 1 1 39438
0 39440 7 2 2 46865 66874
0 39441 7 1 2 52338 71639
0 39442 5 1 1 39441
0 39443 7 1 2 39439 39442
0 39444 5 1 1 39443
0 39445 7 1 2 61868 39444
0 39446 5 1 1 39445
0 39447 7 1 2 50117 70669
0 39448 5 1 1 39447
0 39449 7 1 2 5607 39448
0 39450 5 1 1 39449
0 39451 7 1 2 66412 39450
0 39452 5 1 1 39451
0 39453 7 1 2 51533 71640
0 39454 5 1 1 39453
0 39455 7 1 2 39452 39454
0 39456 5 1 1 39455
0 39457 7 1 2 42636 52464
0 39458 7 1 2 39456 39457
0 39459 5 1 1 39458
0 39460 7 1 2 39446 39459
0 39461 5 1 1 39460
0 39462 7 1 2 48320 39461
0 39463 5 1 1 39462
0 39464 7 1 2 65428 69148
0 39465 5 1 1 39464
0 39466 7 1 2 21420 39465
0 39467 5 1 1 39466
0 39468 7 1 2 49243 39467
0 39469 5 1 1 39468
0 39470 7 1 2 59229 64052
0 39471 5 1 1 39470
0 39472 7 1 2 66876 39471
0 39473 5 1 1 39472
0 39474 7 1 2 49113 39473
0 39475 5 1 1 39474
0 39476 7 1 2 39469 39475
0 39477 5 1 1 39476
0 39478 7 1 2 43174 59940
0 39479 7 1 2 55289 39478
0 39480 7 1 2 39477 39479
0 39481 5 1 1 39480
0 39482 7 1 2 39463 39481
0 39483 5 1 1 39482
0 39484 7 1 2 42926 39483
0 39485 5 1 1 39484
0 39486 7 1 2 55921 71187
0 39487 5 1 1 39486
0 39488 7 1 2 49526 55922
0 39489 5 1 1 39488
0 39490 7 1 2 44127 39489
0 39491 5 1 1 39490
0 39492 7 1 2 71636 39491
0 39493 5 1 1 39492
0 39494 7 1 2 46769 57663
0 39495 5 1 1 39494
0 39496 7 1 2 55633 60206
0 39497 5 1 1 39496
0 39498 7 1 2 17873 39497
0 39499 7 1 2 39495 39498
0 39500 5 1 1 39499
0 39501 7 1 2 43175 39500
0 39502 5 1 1 39501
0 39503 7 1 2 39493 39502
0 39504 5 1 1 39503
0 39505 7 1 2 45331 39504
0 39506 5 1 1 39505
0 39507 7 1 2 50134 52335
0 39508 5 1 1 39507
0 39509 7 1 2 48709 39508
0 39510 5 1 1 39509
0 39511 7 1 2 71564 39510
0 39512 5 1 1 39511
0 39513 7 1 2 55923 39512
0 39514 5 1 1 39513
0 39515 7 1 2 55832 57092
0 39516 7 1 2 67175 39515
0 39517 5 1 1 39516
0 39518 7 1 2 39514 39517
0 39519 7 1 2 39506 39518
0 39520 5 1 1 39519
0 39521 7 1 2 46346 39520
0 39522 5 1 1 39521
0 39523 7 1 2 39487 39522
0 39524 5 1 1 39523
0 39525 7 1 2 52523 66413
0 39526 7 1 2 39524 39525
0 39527 5 1 1 39526
0 39528 7 1 2 39485 39527
0 39529 5 1 1 39528
0 39530 7 1 2 45653 39529
0 39531 5 1 1 39530
0 39532 7 1 2 58536 62092
0 39533 5 1 1 39532
0 39534 7 1 2 64348 66695
0 39535 5 1 1 39534
0 39536 7 1 2 42637 64453
0 39537 7 1 2 39535 39536
0 39538 5 1 1 39537
0 39539 7 1 2 39533 39538
0 39540 5 1 1 39539
0 39541 7 1 2 43176 39540
0 39542 5 1 1 39541
0 39543 7 1 2 59644 64589
0 39544 5 1 1 39543
0 39545 7 1 2 58558 39544
0 39546 5 1 1 39545
0 39547 7 1 2 46347 39546
0 39548 5 1 1 39547
0 39549 7 1 2 50029 36357
0 39550 5 1 1 39549
0 39551 7 1 2 50118 60951
0 39552 5 1 1 39551
0 39553 7 1 2 46565 39552
0 39554 7 1 2 39550 39553
0 39555 5 1 1 39554
0 39556 7 1 2 39548 39555
0 39557 5 1 1 39556
0 39558 7 1 2 51159 39557
0 39559 5 1 1 39558
0 39560 7 1 2 39542 39559
0 39561 5 1 1 39560
0 39562 7 1 2 58740 68283
0 39563 7 1 2 39561 39562
0 39564 5 1 1 39563
0 39565 7 1 2 47699 39564
0 39566 7 1 2 39531 39565
0 39567 5 1 1 39566
0 39568 7 1 2 53616 39567
0 39569 7 1 2 39431 39568
0 39570 5 1 1 39569
0 39571 7 1 2 49624 59541
0 39572 5 1 1 39571
0 39573 7 1 2 45775 61744
0 39574 7 1 2 71226 39573
0 39575 5 1 1 39574
0 39576 7 1 2 39572 39575
0 39577 5 1 1 39576
0 39578 7 1 2 42093 39577
0 39579 5 1 1 39578
0 39580 7 1 2 59667 59888
0 39581 7 1 2 58840 39580
0 39582 5 1 1 39581
0 39583 7 1 2 39579 39582
0 39584 5 2 1 39583
0 39585 7 1 2 68368 71641
0 39586 5 1 1 39585
0 39587 7 1 2 49061 70182
0 39588 7 1 2 64710 39587
0 39589 5 1 1 39588
0 39590 7 1 2 39586 39589
0 39591 5 1 1 39590
0 39592 7 1 2 43400 39591
0 39593 5 1 1 39592
0 39594 7 1 2 60706 69928
0 39595 7 1 2 59446 39594
0 39596 5 1 1 39595
0 39597 7 1 2 39593 39596
0 39598 5 1 1 39597
0 39599 7 1 2 44502 39598
0 39600 5 1 1 39599
0 39601 7 1 2 59944 63761
0 39602 7 1 2 67800 39601
0 39603 7 1 2 71502 39602
0 39604 5 1 1 39603
0 39605 7 1 2 39600 39604
0 39606 5 1 1 39605
0 39607 7 1 2 42927 39606
0 39608 5 1 1 39607
0 39609 7 1 2 28375 69920
0 39610 5 1 1 39609
0 39611 7 1 2 49719 61293
0 39612 7 1 2 59461 39611
0 39613 7 1 2 39610 39612
0 39614 5 1 1 39613
0 39615 7 1 2 39608 39614
0 39616 5 1 1 39615
0 39617 7 1 2 53295 39616
0 39618 5 1 1 39617
0 39619 7 1 2 51808 67326
0 39620 5 1 1 39619
0 39621 7 1 2 46566 64771
0 39622 5 1 1 39621
0 39623 7 1 2 39620 39622
0 39624 5 1 1 39623
0 39625 7 1 2 63618 39624
0 39626 5 1 1 39625
0 39627 7 1 2 71368 39626
0 39628 5 1 1 39627
0 39629 7 1 2 59734 39628
0 39630 5 1 1 39629
0 39631 7 1 2 51160 59447
0 39632 7 1 2 71360 39631
0 39633 5 1 1 39632
0 39634 7 1 2 39630 39633
0 39635 5 1 1 39634
0 39636 7 1 2 66560 39635
0 39637 5 1 1 39636
0 39638 7 2 2 56127 59486
0 39639 7 1 2 69097 71643
0 39640 5 1 1 39639
0 39641 7 1 2 59551 39640
0 39642 5 1 1 39641
0 39643 7 1 2 42094 39642
0 39644 5 1 1 39643
0 39645 7 1 2 61458 63096
0 39646 7 1 2 68265 39645
0 39647 5 1 1 39646
0 39648 7 1 2 39644 39647
0 39649 5 1 1 39648
0 39650 7 1 2 47468 39649
0 39651 5 1 1 39650
0 39652 7 1 2 59809 68392
0 39653 5 1 1 39652
0 39654 7 1 2 39651 39653
0 39655 5 1 1 39654
0 39656 7 1 2 50119 39655
0 39657 5 1 1 39656
0 39658 7 1 2 69095 71003
0 39659 5 1 1 39658
0 39660 7 1 2 59552 39659
0 39661 5 1 1 39660
0 39662 7 1 2 42095 39661
0 39663 5 1 1 39662
0 39664 7 1 2 58108 69953
0 39665 5 1 1 39664
0 39666 7 1 2 39663 39665
0 39667 5 1 1 39666
0 39668 7 1 2 50578 39667
0 39669 5 1 1 39668
0 39670 7 1 2 39657 39669
0 39671 5 1 1 39670
0 39672 7 1 2 55153 39671
0 39673 5 1 1 39672
0 39674 7 1 2 63978 65589
0 39675 5 1 1 39674
0 39676 7 1 2 5390 39675
0 39677 5 1 1 39676
0 39678 7 1 2 59735 39677
0 39679 5 1 1 39678
0 39680 7 1 2 42638 28057
0 39681 7 1 2 59448 39680
0 39682 5 1 1 39681
0 39683 7 1 2 39679 39682
0 39684 5 1 1 39683
0 39685 7 1 2 46348 39684
0 39686 5 1 1 39685
0 39687 7 1 2 43177 69187
0 39688 7 1 2 67977 39687
0 39689 5 1 1 39688
0 39690 7 1 2 39686 39689
0 39691 7 1 2 39673 39690
0 39692 5 1 1 39691
0 39693 7 1 2 50371 64666
0 39694 7 1 2 39692 39693
0 39695 5 1 1 39694
0 39696 7 1 2 39637 39695
0 39697 5 1 1 39696
0 39698 7 1 2 44503 39697
0 39699 5 1 1 39698
0 39700 7 1 2 39618 39699
0 39701 5 1 1 39700
0 39702 7 1 2 48321 39701
0 39703 5 1 1 39702
0 39704 7 1 2 68078 71279
0 39705 5 1 1 39704
0 39706 7 1 2 60697 39705
0 39707 5 1 1 39706
0 39708 7 1 2 71209 39707
0 39709 5 1 1 39708
0 39710 7 1 2 59798 60844
0 39711 5 1 1 39710
0 39712 7 1 2 60698 39711
0 39713 5 1 1 39712
0 39714 7 1 2 55290 39713
0 39715 5 1 1 39714
0 39716 7 1 2 39709 39715
0 39717 5 1 1 39716
0 39718 7 1 2 70115 39717
0 39719 5 1 1 39718
0 39720 7 1 2 7055 33633
0 39721 5 1 1 39720
0 39722 7 1 2 71210 39721
0 39723 5 1 1 39722
0 39724 7 2 2 42639 59985
0 39725 7 1 2 54066 67973
0 39726 7 1 2 71645 39725
0 39727 5 1 1 39726
0 39728 7 1 2 39723 39727
0 39729 5 1 1 39728
0 39730 7 1 2 45654 39729
0 39731 5 1 1 39730
0 39732 7 1 2 54748 57737
0 39733 7 1 2 58514 39732
0 39734 5 1 1 39733
0 39735 7 1 2 39731 39734
0 39736 5 1 1 39735
0 39737 7 1 2 43401 39736
0 39738 5 1 1 39737
0 39739 7 1 2 50208 58924
0 39740 7 1 2 60016 39739
0 39741 5 1 1 39740
0 39742 7 1 2 39738 39741
0 39743 5 1 1 39742
0 39744 7 1 2 69090 39743
0 39745 5 1 1 39744
0 39746 7 1 2 39719 39745
0 39747 5 1 1 39746
0 39748 7 1 2 48710 39747
0 39749 5 1 1 39748
0 39750 7 1 2 60600 67791
0 39751 7 2 2 70394 39750
0 39752 7 1 2 55510 71647
0 39753 5 1 1 39752
0 39754 7 1 2 39749 39753
0 39755 5 1 1 39754
0 39756 7 1 2 67520 39755
0 39757 5 1 1 39756
0 39758 7 1 2 49800 50675
0 39759 7 1 2 69594 39758
0 39760 7 1 2 71054 71254
0 39761 7 1 2 39759 39760
0 39762 5 1 1 39761
0 39763 7 1 2 39757 39762
0 39764 5 1 1 39763
0 39765 7 1 2 49367 39764
0 39766 5 1 1 39765
0 39767 7 1 2 42928 71642
0 39768 5 1 1 39767
0 39769 7 1 2 59617 70131
0 39770 7 1 2 69175 39769
0 39771 5 1 1 39770
0 39772 7 1 2 39768 39771
0 39773 5 1 1 39772
0 39774 7 1 2 43402 39773
0 39775 5 1 1 39774
0 39776 7 1 2 58846 71411
0 39777 5 1 1 39776
0 39778 7 1 2 39775 39777
0 39779 5 1 1 39778
0 39780 7 1 2 68369 39779
0 39781 5 1 1 39780
0 39782 7 1 2 43565 59608
0 39783 7 1 2 60868 39782
0 39784 7 1 2 68675 69993
0 39785 7 1 2 39783 39784
0 39786 5 1 1 39785
0 39787 7 1 2 39781 39786
0 39788 5 1 1 39787
0 39789 7 1 2 56458 58231
0 39790 7 1 2 39788 39789
0 39791 5 1 1 39790
0 39792 7 1 2 44837 39791
0 39793 7 1 2 39766 39792
0 39794 7 1 2 39703 39793
0 39795 7 1 2 39570 39794
0 39796 7 1 2 39302 39795
0 39797 5 1 1 39796
0 39798 7 1 2 42096 64173
0 39799 7 1 2 63489 39798
0 39800 5 2 1 39799
0 39801 7 1 2 49099 62546
0 39802 5 1 1 39801
0 39803 7 1 2 56892 63708
0 39804 5 1 1 39803
0 39805 7 1 2 39802 39804
0 39806 5 1 1 39805
0 39807 7 1 2 57536 39806
0 39808 5 1 1 39807
0 39809 7 1 2 58904 68858
0 39810 7 1 2 59418 39809
0 39811 5 1 1 39810
0 39812 7 1 2 39808 39811
0 39813 5 1 1 39812
0 39814 7 1 2 46770 39813
0 39815 5 1 1 39814
0 39816 7 1 2 5335 59505
0 39817 5 1 1 39816
0 39818 7 1 2 64670 39817
0 39819 5 1 1 39818
0 39820 7 1 2 39815 39819
0 39821 5 1 1 39820
0 39822 7 1 2 46567 39821
0 39823 5 1 1 39822
0 39824 7 1 2 71649 39823
0 39825 5 1 1 39824
0 39826 7 1 2 48322 39825
0 39827 5 1 1 39826
0 39828 7 1 2 57685 64567
0 39829 7 1 2 62945 39828
0 39830 5 1 1 39829
0 39831 7 1 2 39827 39830
0 39832 5 1 1 39831
0 39833 7 1 2 59496 39832
0 39834 5 1 1 39833
0 39835 7 1 2 737 39398
0 39836 5 1 1 39835
0 39837 7 1 2 70936 39836
0 39838 5 1 1 39837
0 39839 7 1 2 60512 68960
0 39840 7 1 2 53868 39839
0 39841 5 1 1 39840
0 39842 7 1 2 39838 39841
0 39843 5 1 1 39842
0 39844 7 1 2 59542 39843
0 39845 5 1 1 39844
0 39846 7 1 2 50434 71628
0 39847 5 1 1 39846
0 39848 7 1 2 44982 39847
0 39849 5 1 1 39848
0 39850 7 1 2 39845 39849
0 39851 7 1 2 39834 39850
0 39852 5 1 1 39851
0 39853 7 1 2 71156 71354
0 39854 5 1 1 39853
0 39855 7 1 2 64671 64590
0 39856 5 1 1 39855
0 39857 7 1 2 39854 39856
0 39858 5 1 1 39857
0 39859 7 1 2 46568 39858
0 39860 5 1 1 39859
0 39861 7 1 2 39860 71650
0 39862 5 1 1 39861
0 39863 7 1 2 59497 39862
0 39864 5 1 1 39863
0 39865 7 1 2 69871 71426
0 39866 5 1 1 39865
0 39867 7 1 2 50479 39866
0 39868 7 1 2 71629 39867
0 39869 7 1 2 39864 39868
0 39870 5 1 1 39869
0 39871 7 1 2 2297 39870
0 39872 7 1 2 39852 39871
0 39873 5 1 1 39872
0 39874 7 1 2 60132 59967
0 39875 7 1 2 68318 39874
0 39876 7 2 2 61668 39875
0 39877 7 1 2 55660 71590
0 39878 7 1 2 71651 39877
0 39879 5 1 1 39878
0 39880 7 1 2 39873 39879
0 39881 5 1 1 39880
0 39882 7 1 2 51189 39881
0 39883 5 1 1 39882
0 39884 7 1 2 57686 64380
0 39885 7 1 2 71652 39884
0 39886 5 1 1 39885
0 39887 7 1 2 39883 39886
0 39888 5 1 1 39887
0 39889 7 1 2 66793 39888
0 39890 5 1 1 39889
0 39891 7 1 2 58350 66523
0 39892 5 1 1 39891
0 39893 7 1 2 55203 66507
0 39894 5 1 1 39893
0 39895 7 1 2 39892 39894
0 39896 5 1 1 39895
0 39897 7 1 2 49770 39896
0 39898 5 1 1 39897
0 39899 7 1 2 62379 66524
0 39900 5 1 1 39899
0 39901 7 1 2 39898 39900
0 39902 5 1 1 39901
0 39903 7 1 2 62547 39902
0 39904 5 1 1 39903
0 39905 7 1 2 60481 69990
0 39906 5 1 1 39905
0 39907 7 2 2 61487 64701
0 39908 5 1 1 71653
0 39909 7 1 2 39906 39908
0 39910 5 1 1 39909
0 39911 7 1 2 50579 39910
0 39912 5 1 1 39911
0 39913 7 1 2 39904 39912
0 39914 5 1 1 39913
0 39915 7 1 2 43403 39914
0 39916 5 1 1 39915
0 39917 7 1 2 71555 71654
0 39918 5 1 1 39917
0 39919 7 1 2 39916 39918
0 39920 5 1 1 39919
0 39921 7 1 2 59498 39920
0 39922 5 1 1 39921
0 39923 7 1 2 62548 69932
0 39924 5 1 1 39923
0 39925 7 2 2 57647 63029
0 39926 7 3 2 48039 71655
0 39927 7 1 2 61115 71657
0 39928 5 1 1 39927
0 39929 7 1 2 39924 39928
0 39930 5 1 1 39929
0 39931 7 1 2 59543 39930
0 39932 5 1 1 39931
0 39933 7 1 2 39922 39932
0 39934 5 1 1 39933
0 39935 7 1 2 46349 39934
0 39936 5 1 1 39935
0 39937 7 1 2 54719 71370
0 39938 5 1 1 39937
0 39939 7 2 2 60653 39938
0 39940 7 1 2 53696 71660
0 39941 5 1 1 39940
0 39942 7 1 2 57543 59499
0 39943 5 1 1 39942
0 39944 7 1 2 49771 59544
0 39945 5 1 1 39944
0 39946 7 1 2 39943 39945
0 39947 5 1 1 39946
0 39948 7 1 2 42097 61306
0 39949 7 1 2 39947 39948
0 39950 5 1 1 39949
0 39951 7 1 2 39941 39950
0 39952 5 1 1 39951
0 39953 7 1 2 66561 39952
0 39954 5 1 1 39953
0 39955 7 1 2 42351 67081
0 39956 7 1 2 69236 39955
0 39957 5 1 1 39956
0 39958 7 1 2 58121 59487
0 39959 7 1 2 60961 39958
0 39960 7 1 2 66806 39959
0 39961 5 1 1 39960
0 39962 7 1 2 39957 39961
0 39963 5 1 1 39962
0 39964 7 1 2 60955 39963
0 39965 5 1 1 39964
0 39966 7 1 2 68524 70593
0 39967 7 1 2 65634 39966
0 39968 5 1 1 39967
0 39969 7 1 2 39965 39968
0 39970 7 1 2 39954 39969
0 39971 5 1 1 39970
0 39972 7 1 2 47594 39971
0 39973 5 1 1 39972
0 39974 7 1 2 57621 64038
0 39975 7 1 2 64822 66759
0 39976 7 1 2 39974 39975
0 39977 5 1 1 39976
0 39978 7 1 2 49772 64311
0 39979 7 1 2 68200 39978
0 39980 5 1 1 39979
0 39981 7 1 2 39977 39980
0 39982 7 1 2 39973 39981
0 39983 5 1 1 39982
0 39984 7 1 2 46771 39983
0 39985 5 1 1 39984
0 39986 7 1 2 60214 71658
0 39987 5 1 1 39986
0 39988 7 1 2 42098 49633
0 39989 7 1 2 66807 39988
0 39990 5 1 1 39989
0 39991 7 1 2 39987 39990
0 39992 5 1 1 39991
0 39993 7 1 2 47469 39992
0 39994 5 1 1 39993
0 39995 7 1 2 69930 71345
0 39996 5 1 1 39995
0 39997 7 1 2 39994 39996
0 39998 5 1 1 39997
0 39999 7 1 2 46569 39998
0 40000 5 1 1 39999
0 40001 7 1 2 50580 68308
0 40002 5 1 1 40001
0 40003 7 1 2 40000 40002
0 40004 5 1 1 40003
0 40005 7 1 2 59545 40004
0 40006 5 1 1 40005
0 40007 7 1 2 60236 68019
0 40008 7 1 2 67657 69895
0 40009 7 1 2 71591 40008
0 40010 7 1 2 40007 40009
0 40011 5 1 1 40010
0 40012 7 1 2 40006 40011
0 40013 7 1 2 39985 40012
0 40014 7 1 2 39936 40013
0 40015 5 1 1 40014
0 40016 7 1 2 53296 40015
0 40017 5 1 1 40016
0 40018 7 2 2 56360 66784
0 40019 5 1 1 71662
0 40020 7 1 2 34936 40019
0 40021 5 1 1 40020
0 40022 7 1 2 62813 40021
0 40023 5 1 1 40022
0 40024 7 1 2 58595 66562
0 40025 5 1 1 40024
0 40026 7 1 2 40023 40025
0 40027 5 1 1 40026
0 40028 7 1 2 43404 40027
0 40029 5 1 1 40028
0 40030 7 1 2 47153 69995
0 40031 5 1 1 40030
0 40032 7 1 2 40029 40031
0 40033 5 1 1 40032
0 40034 7 1 2 63619 40033
0 40035 5 1 1 40034
0 40036 7 1 2 53733 69917
0 40037 5 1 1 40036
0 40038 7 1 2 48711 71111
0 40039 5 1 1 40038
0 40040 7 1 2 40037 40039
0 40041 5 1 1 40040
0 40042 7 1 2 54069 40041
0 40043 5 1 1 40042
0 40044 7 1 2 40035 40043
0 40045 5 1 1 40044
0 40046 7 1 2 62549 40045
0 40047 5 1 1 40046
0 40048 7 1 2 64719 67944
0 40049 5 1 1 40048
0 40050 7 1 2 68139 40049
0 40051 5 1 1 40050
0 40052 7 1 2 49368 50435
0 40053 7 1 2 64515 40052
0 40054 7 1 2 40051 40053
0 40055 5 1 1 40054
0 40056 7 1 2 40047 40055
0 40057 5 1 1 40056
0 40058 7 1 2 59546 40057
0 40059 5 1 1 40058
0 40060 7 1 2 63979 66508
0 40061 5 1 1 40060
0 40062 7 1 2 64720 70082
0 40063 5 1 1 40062
0 40064 7 1 2 40061 40063
0 40065 5 1 1 40064
0 40066 7 1 2 71323 40065
0 40067 5 1 1 40066
0 40068 7 2 2 51774 66707
0 40069 7 1 2 64696 71664
0 40070 5 1 1 40069
0 40071 7 1 2 40067 40070
0 40072 5 1 1 40071
0 40073 7 1 2 43178 40072
0 40074 5 1 1 40073
0 40075 7 1 2 53495 70740
0 40076 7 1 2 71656 40075
0 40077 5 1 1 40076
0 40078 7 1 2 40074 40077
0 40079 5 1 1 40078
0 40080 7 1 2 59889 67959
0 40081 7 1 2 60800 40080
0 40082 7 1 2 40079 40081
0 40083 5 1 1 40082
0 40084 7 1 2 40059 40083
0 40085 7 1 2 40017 40084
0 40086 5 1 1 40085
0 40087 7 1 2 44983 40086
0 40088 5 1 1 40087
0 40089 7 5 2 60654 70116
0 40090 7 1 2 46772 55304
0 40091 5 1 1 40090
0 40092 7 1 2 50197 2895
0 40093 5 1 1 40092
0 40094 7 1 2 49846 9350
0 40095 5 1 1 40094
0 40096 7 1 2 40093 40095
0 40097 5 1 1 40096
0 40098 7 1 2 40091 40097
0 40099 5 1 1 40098
0 40100 7 1 2 71666 40099
0 40101 5 1 1 40100
0 40102 7 1 2 43179 54345
0 40103 5 1 1 40102
0 40104 7 1 2 71567 40103
0 40105 5 1 1 40104
0 40106 7 1 2 58559 71565
0 40107 7 1 2 40105 40106
0 40108 5 1 1 40107
0 40109 7 1 2 66828 40108
0 40110 5 1 1 40109
0 40111 7 1 2 40101 40110
0 40112 5 1 1 40111
0 40113 7 1 2 54814 40112
0 40114 5 1 1 40113
0 40115 7 1 2 63411 70981
0 40116 5 1 1 40115
0 40117 7 1 2 60007 62136
0 40118 7 1 2 71176 40117
0 40119 5 1 1 40118
0 40120 7 1 2 40116 40119
0 40121 5 1 1 40120
0 40122 7 1 2 50120 40121
0 40123 5 1 1 40122
0 40124 7 1 2 56662 63405
0 40125 7 1 2 66835 40124
0 40126 5 1 1 40125
0 40127 7 1 2 40123 40126
0 40128 5 1 1 40127
0 40129 7 1 2 43484 40128
0 40130 5 1 1 40129
0 40131 7 1 2 59579 68353
0 40132 7 1 2 70051 40131
0 40133 5 1 1 40132
0 40134 7 1 2 40130 40133
0 40135 5 1 1 40134
0 40136 7 1 2 44504 40135
0 40137 5 1 1 40136
0 40138 7 1 2 64697 71096
0 40139 5 1 1 40138
0 40140 7 1 2 70595 71093
0 40141 5 1 1 40140
0 40142 7 1 2 40139 40141
0 40143 5 1 1 40142
0 40144 7 1 2 62608 40143
0 40145 5 1 1 40144
0 40146 7 1 2 56663 70078
0 40147 5 1 1 40146
0 40148 7 1 2 50807 55674
0 40149 7 1 2 61442 63838
0 40150 7 1 2 40148 40149
0 40151 5 1 1 40150
0 40152 7 1 2 40147 40151
0 40153 5 1 1 40152
0 40154 7 1 2 59414 40153
0 40155 5 1 1 40154
0 40156 7 1 2 40145 40155
0 40157 7 1 2 40137 40156
0 40158 7 1 2 40114 40157
0 40159 5 1 1 40158
0 40160 7 1 2 53888 40159
0 40161 5 1 1 40160
0 40162 7 1 2 59799 71533
0 40163 5 1 1 40162
0 40164 7 1 2 59815 40163
0 40165 5 1 1 40164
0 40166 7 1 2 66888 40165
0 40167 5 1 1 40166
0 40168 7 1 2 66829 71184
0 40169 5 1 1 40168
0 40170 7 1 2 71377 71667
0 40171 5 1 1 40170
0 40172 7 1 2 40169 40171
0 40173 5 1 1 40172
0 40174 7 1 2 54815 40173
0 40175 5 1 1 40174
0 40176 7 1 2 61659 65836
0 40177 7 1 2 71395 40176
0 40178 5 1 1 40177
0 40179 7 1 2 40175 40178
0 40180 7 1 2 40167 40179
0 40181 5 1 1 40180
0 40182 7 1 2 59718 40181
0 40183 5 1 1 40182
0 40184 7 1 2 40161 40183
0 40185 5 1 1 40184
0 40186 7 1 2 46350 40185
0 40187 5 1 1 40186
0 40188 7 1 2 48858 71648
0 40189 5 1 1 40188
0 40190 7 1 2 50885 71668
0 40191 5 1 1 40190
0 40192 7 1 2 51775 66830
0 40193 5 1 1 40192
0 40194 7 1 2 40191 40193
0 40195 5 1 1 40194
0 40196 7 1 2 49369 40195
0 40197 5 1 1 40196
0 40198 7 1 2 40189 40197
0 40199 5 1 1 40198
0 40200 7 1 2 48712 40199
0 40201 5 1 1 40200
0 40202 7 1 2 55479 71669
0 40203 5 1 1 40202
0 40204 7 1 2 44128 71105
0 40205 5 1 1 40204
0 40206 7 1 2 40203 40205
0 40207 7 1 2 40201 40206
0 40208 5 1 1 40207
0 40209 7 1 2 63582 40208
0 40210 5 1 1 40209
0 40211 7 1 2 52395 64649
0 40212 7 1 2 49889 40211
0 40213 7 1 2 66966 40212
0 40214 5 1 1 40213
0 40215 7 1 2 40210 40214
0 40216 5 1 1 40215
0 40217 7 1 2 60254 40216
0 40218 5 1 1 40217
0 40219 7 1 2 55210 71670
0 40220 5 1 1 40219
0 40221 7 1 2 54990 55329
0 40222 7 1 2 66831 40221
0 40223 5 1 1 40222
0 40224 7 1 2 40220 40223
0 40225 5 1 1 40224
0 40226 7 1 2 46773 40225
0 40227 5 1 1 40226
0 40228 7 1 2 63981 66832
0 40229 5 1 1 40228
0 40230 7 1 2 49844 60188
0 40231 7 1 2 70036 40230
0 40232 5 1 1 40231
0 40233 7 1 2 40229 40232
0 40234 5 1 1 40233
0 40235 7 1 2 46570 40234
0 40236 5 1 1 40235
0 40237 7 1 2 40227 40236
0 40238 5 1 1 40237
0 40239 7 1 2 50581 53941
0 40240 7 1 2 40238 40239
0 40241 5 1 1 40240
0 40242 7 1 2 40218 40241
0 40243 5 1 1 40242
0 40244 7 1 2 54816 40243
0 40245 5 1 1 40244
0 40246 7 1 2 49773 59866
0 40247 5 1 1 40246
0 40248 7 1 2 35432 40247
0 40249 5 1 1 40248
0 40250 7 1 2 66883 40249
0 40251 5 1 1 40250
0 40252 7 1 2 60499 71592
0 40253 7 1 2 70103 40252
0 40254 5 1 1 40253
0 40255 7 1 2 40251 40254
0 40256 5 1 1 40255
0 40257 7 1 2 51239 40256
0 40258 5 1 1 40257
0 40259 7 1 2 66889 71236
0 40260 5 1 1 40259
0 40261 7 1 2 40258 40260
0 40262 5 1 1 40261
0 40263 7 1 2 46571 40262
0 40264 5 1 1 40263
0 40265 7 1 2 51240 70606
0 40266 7 1 2 55451 40265
0 40267 5 1 1 40266
0 40268 7 1 2 40264 40267
0 40269 5 1 1 40268
0 40270 7 1 2 59719 40269
0 40271 5 1 1 40270
0 40272 7 1 2 57994 71232
0 40273 5 1 1 40272
0 40274 7 1 2 51480 57995
0 40275 5 1 1 40274
0 40276 7 1 2 57587 40275
0 40277 5 1 1 40276
0 40278 7 1 2 59867 40277
0 40279 5 1 1 40278
0 40280 7 1 2 40273 40279
0 40281 5 1 1 40280
0 40282 7 1 2 66890 40281
0 40283 5 1 1 40282
0 40284 7 1 2 67176 66992
0 40285 7 1 2 70063 71132
0 40286 7 1 2 40284 40285
0 40287 5 1 1 40286
0 40288 7 1 2 48323 40287
0 40289 7 1 2 40283 40288
0 40290 5 1 1 40289
0 40291 7 1 2 71199 71201
0 40292 5 1 1 40291
0 40293 7 1 2 50030 40292
0 40294 5 1 1 40293
0 40295 7 1 2 54226 69959
0 40296 5 1 1 40295
0 40297 7 1 2 40294 40296
0 40298 5 1 1 40297
0 40299 7 1 2 66891 40298
0 40300 5 1 1 40299
0 40301 7 1 2 61976 70607
0 40302 7 1 2 71243 40301
0 40303 5 1 1 40302
0 40304 7 1 2 59932 67236
0 40305 5 1 1 40304
0 40306 7 1 2 42929 66892
0 40307 7 1 2 40305 40306
0 40308 5 1 1 40307
0 40309 7 1 2 40303 40308
0 40310 5 1 1 40309
0 40311 7 1 2 50886 40310
0 40312 5 1 1 40311
0 40313 7 1 2 40300 40312
0 40314 5 1 1 40313
0 40315 7 1 2 48713 40314
0 40316 5 1 1 40315
0 40317 7 1 2 58205 65197
0 40318 7 1 2 70302 40317
0 40319 7 1 2 66893 40318
0 40320 5 1 1 40319
0 40321 7 1 2 44984 40320
0 40322 7 1 2 40316 40321
0 40323 5 1 1 40322
0 40324 7 1 2 50436 40323
0 40325 7 1 2 40290 40324
0 40326 5 1 1 40325
0 40327 7 1 2 40271 40326
0 40328 7 1 2 40245 40327
0 40329 7 1 2 40187 40328
0 40330 5 1 1 40329
0 40331 7 1 2 53617 40330
0 40332 5 1 1 40331
0 40333 7 2 2 61799 63412
0 40334 5 1 1 71671
0 40335 7 1 2 62592 69112
0 40336 5 1 1 40335
0 40337 7 1 2 40334 40336
0 40338 5 1 1 40337
0 40339 7 1 2 60956 40338
0 40340 5 1 1 40339
0 40341 7 1 2 60551 71362
0 40342 5 1 1 40341
0 40343 7 1 2 42099 71661
0 40344 5 1 1 40343
0 40345 7 1 2 40342 40344
0 40346 5 1 1 40345
0 40347 7 1 2 66563 40346
0 40348 5 1 1 40347
0 40349 7 1 2 40340 40348
0 40350 5 1 1 40349
0 40351 7 1 2 50808 40350
0 40352 5 1 1 40351
0 40353 7 1 2 45655 50031
0 40354 7 1 2 64634 40353
0 40355 5 1 1 40354
0 40356 7 1 2 12087 40355
0 40357 5 1 1 40356
0 40358 7 1 2 64946 40357
0 40359 5 1 1 40358
0 40360 7 1 2 59170 69909
0 40361 7 1 2 51087 40360
0 40362 5 1 1 40361
0 40363 7 1 2 40359 40362
0 40364 5 1 1 40363
0 40365 7 1 2 66564 40364
0 40366 5 1 1 40365
0 40367 7 1 2 50372 50809
0 40368 7 1 2 51412 40367
0 40369 5 1 1 40368
0 40370 7 1 2 36535 40369
0 40371 5 1 1 40370
0 40372 7 1 2 62593 66491
0 40373 7 1 2 40371 40372
0 40374 5 1 1 40373
0 40375 7 1 2 40366 40374
0 40376 7 1 2 40352 40375
0 40377 5 1 1 40376
0 40378 7 1 2 53297 40377
0 40379 5 1 1 40378
0 40380 7 1 2 50373 54024
0 40381 7 1 2 70608 40380
0 40382 5 1 1 40381
0 40383 7 1 2 61660 71445
0 40384 5 1 1 40383
0 40385 7 1 2 36622 40384
0 40386 5 1 1 40385
0 40387 7 1 2 50887 66794
0 40388 7 1 2 40386 40387
0 40389 5 1 1 40388
0 40390 7 1 2 40382 40389
0 40391 5 1 1 40390
0 40392 7 1 2 48859 40391
0 40393 5 1 1 40392
0 40394 7 1 2 57819 71672
0 40395 5 1 1 40394
0 40396 7 1 2 60552 66795
0 40397 7 1 2 60823 40396
0 40398 5 1 1 40397
0 40399 7 1 2 40395 40398
0 40400 5 1 1 40399
0 40401 7 1 2 42930 40400
0 40402 5 1 1 40401
0 40403 7 1 2 40393 40402
0 40404 5 1 1 40403
0 40405 7 1 2 48714 40404
0 40406 5 1 1 40405
0 40407 7 1 2 50966 71311
0 40408 7 1 2 71665 40407
0 40409 5 1 1 40408
0 40410 7 1 2 40406 40409
0 40411 5 1 1 40410
0 40412 7 1 2 50437 40411
0 40413 5 1 1 40412
0 40414 7 1 2 40379 40413
0 40415 5 1 1 40414
0 40416 7 1 2 44985 40415
0 40417 5 1 1 40416
0 40418 7 1 2 47700 57687
0 40419 7 2 2 65461 40418
0 40420 7 2 2 47154 71673
0 40421 7 1 2 59991 71675
0 40422 5 1 1 40421
0 40423 7 1 2 52468 60655
0 40424 7 2 2 71241 40423
0 40425 5 1 1 71677
0 40426 7 1 2 42100 40425
0 40427 5 1 1 40426
0 40428 7 2 2 43781 71674
0 40429 5 1 1 71679
0 40430 7 1 2 45656 40429
0 40431 5 1 1 40430
0 40432 7 1 2 46101 40431
0 40433 7 1 2 40427 40432
0 40434 5 1 1 40433
0 40435 7 1 2 40422 40434
0 40436 5 1 1 40435
0 40437 7 1 2 66585 40436
0 40438 5 1 1 40437
0 40439 7 1 2 69178 69302
0 40440 5 1 1 40439
0 40441 7 1 2 65458 66509
0 40442 5 1 1 40441
0 40443 7 1 2 40440 40442
0 40444 5 1 1 40443
0 40445 7 1 2 51241 40444
0 40446 5 1 1 40445
0 40447 7 1 2 60207 71663
0 40448 5 1 1 40447
0 40449 7 1 2 50032 66565
0 40450 5 1 1 40449
0 40451 7 1 2 51214 66510
0 40452 5 1 1 40451
0 40453 7 1 2 40450 40452
0 40454 5 1 1 40453
0 40455 7 1 2 51088 40454
0 40456 5 1 1 40455
0 40457 7 1 2 40448 40456
0 40458 5 1 1 40457
0 40459 7 1 2 46351 40458
0 40460 5 1 1 40459
0 40461 7 1 2 40446 40460
0 40462 5 1 1 40461
0 40463 7 1 2 60553 40462
0 40464 5 1 1 40463
0 40465 7 1 2 64721 66637
0 40466 5 2 1 40465
0 40467 7 1 2 64067 66511
0 40468 5 1 1 40467
0 40469 7 1 2 71681 40468
0 40470 5 1 1 40469
0 40471 7 1 2 51043 40470
0 40472 5 1 1 40471
0 40473 7 2 2 46774 68137
0 40474 5 1 1 71683
0 40475 7 1 2 71682 40474
0 40476 5 2 1 40475
0 40477 7 1 2 45332 71685
0 40478 5 1 1 40477
0 40479 7 1 2 40472 40478
0 40480 5 1 1 40479
0 40481 7 1 2 46352 40480
0 40482 5 1 1 40481
0 40483 7 1 2 65676 66525
0 40484 5 1 1 40483
0 40485 7 1 2 46572 71684
0 40486 5 1 1 40485
0 40487 7 1 2 40484 40486
0 40488 5 1 1 40487
0 40489 7 1 2 50582 40488
0 40490 5 1 1 40489
0 40491 7 1 2 40482 40490
0 40492 5 1 1 40491
0 40493 7 1 2 59415 40492
0 40494 5 1 1 40493
0 40495 7 1 2 40464 40494
0 40496 5 1 1 40495
0 40497 7 1 2 53889 40496
0 40498 5 1 1 40497
0 40499 7 1 2 40438 40498
0 40500 7 1 2 40417 40499
0 40501 5 1 1 40500
0 40502 7 1 2 53680 40501
0 40503 5 1 1 40502
0 40504 7 1 2 59547 65677
0 40505 5 1 1 40504
0 40506 7 1 2 69945 40505
0 40507 5 1 1 40506
0 40508 7 1 2 47470 40507
0 40509 5 1 1 40508
0 40510 7 1 2 46353 59609
0 40511 7 1 2 59129 40510
0 40512 5 1 1 40511
0 40513 7 1 2 40509 40512
0 40514 5 1 1 40513
0 40515 7 1 2 71659 40514
0 40516 5 1 1 40515
0 40517 7 1 2 46354 63431
0 40518 5 1 1 40517
0 40519 7 1 2 59500 71518
0 40520 7 1 2 40518 40519
0 40521 5 1 1 40520
0 40522 7 1 2 59553 40521
0 40523 5 1 1 40522
0 40524 7 1 2 71347 40523
0 40525 5 1 1 40524
0 40526 7 1 2 48860 57580
0 40527 5 1 1 40526
0 40528 7 1 2 3917 40527
0 40529 5 1 1 40528
0 40530 7 1 2 46573 40529
0 40531 5 1 1 40530
0 40532 7 1 2 46355 60754
0 40533 7 1 2 62370 40532
0 40534 5 1 1 40533
0 40535 7 1 2 40531 40534
0 40536 5 1 1 40535
0 40537 7 1 2 59548 40536
0 40538 5 1 1 40537
0 40539 7 1 2 56879 58799
0 40540 7 1 2 71126 40539
0 40541 5 1 1 40540
0 40542 7 1 2 40538 40541
0 40543 5 1 1 40542
0 40544 7 1 2 60482 40543
0 40545 5 1 1 40544
0 40546 7 1 2 40525 40545
0 40547 5 1 1 40546
0 40548 7 1 2 68370 40547
0 40549 5 1 1 40548
0 40550 7 1 2 40516 40549
0 40551 5 1 1 40550
0 40552 7 1 2 45333 40551
0 40553 5 1 1 40552
0 40554 7 1 2 71337 71686
0 40555 5 1 1 40554
0 40556 7 1 2 68310 40555
0 40557 5 1 1 40556
0 40558 7 1 2 67905 40557
0 40559 5 1 1 40558
0 40560 7 1 2 40553 40559
0 40561 5 1 1 40560
0 40562 7 1 2 53890 40561
0 40563 5 1 1 40562
0 40564 7 1 2 58126 71680
0 40565 5 1 1 40564
0 40566 7 1 2 53697 71678
0 40567 5 1 1 40566
0 40568 7 1 2 40565 40567
0 40569 5 1 1 40568
0 40570 7 1 2 46102 40569
0 40571 5 1 1 40570
0 40572 7 1 2 52149 59024
0 40573 7 1 2 71676 40572
0 40574 5 1 1 40573
0 40575 7 1 2 40571 40574
0 40576 5 1 1 40575
0 40577 7 1 2 66586 40576
0 40578 5 1 1 40577
0 40579 7 1 2 48162 40578
0 40580 7 1 2 40563 40579
0 40581 7 1 2 40503 40580
0 40582 7 1 2 40332 40581
0 40583 7 1 2 40088 40582
0 40584 7 1 2 39890 40583
0 40585 5 1 1 40584
0 40586 7 1 2 66284 40585
0 40587 7 1 2 39797 40586
0 40588 5 1 1 40587
0 40589 7 1 2 39145 40588
0 40590 7 1 2 38568 40589
0 40591 7 1 2 36817 40590
0 40592 5 1 1 40591
0 40593 7 1 2 54289 40592
0 40594 5 1 1 40593
0 40595 7 1 2 42241 67230
0 40596 5 1 1 40595
0 40597 7 1 2 56478 62872
0 40598 5 1 1 40597
0 40599 7 1 2 40596 40598
0 40600 5 1 1 40599
0 40601 7 1 2 45873 40600
0 40602 5 1 1 40601
0 40603 7 2 2 47926 67270
0 40604 5 1 1 71687
0 40605 7 1 2 64006 71688
0 40606 5 1 1 40605
0 40607 7 1 2 40602 40606
0 40608 5 1 1 40607
0 40609 7 1 2 44505 40608
0 40610 5 1 1 40609
0 40611 7 1 2 56493 63805
0 40612 5 1 1 40611
0 40613 7 1 2 40610 40612
0 40614 5 1 1 40613
0 40615 7 1 2 46775 40614
0 40616 5 1 1 40615
0 40617 7 2 2 57953 60113
0 40618 7 1 2 69117 71689
0 40619 5 1 1 40618
0 40620 7 1 2 40616 40619
0 40621 5 1 1 40620
0 40622 7 1 2 46866 40621
0 40623 5 1 1 40622
0 40624 7 1 2 54511 70142
0 40625 7 1 2 71690 40624
0 40626 5 1 1 40625
0 40627 7 1 2 40623 40626
0 40628 5 1 1 40627
0 40629 7 1 2 49310 40628
0 40630 5 1 1 40629
0 40631 7 2 2 56521 67224
0 40632 7 1 2 57901 60679
0 40633 7 1 2 63223 40632
0 40634 7 1 2 71691 40633
0 40635 5 1 1 40634
0 40636 7 1 2 40630 40635
0 40637 5 1 1 40636
0 40638 7 1 2 50438 40637
0 40639 5 1 1 40638
0 40640 7 1 2 46867 53059
0 40641 7 1 2 63458 40640
0 40642 7 1 2 56442 56535
0 40643 7 1 2 68516 40642
0 40644 7 1 2 40641 40643
0 40645 5 1 1 40644
0 40646 7 1 2 40639 40645
0 40647 5 1 1 40646
0 40648 7 1 2 69536 40647
0 40649 5 1 1 40648
0 40650 7 1 2 45776 67678
0 40651 7 1 2 57505 40650
0 40652 7 1 2 64489 67124
0 40653 7 1 2 40651 40652
0 40654 7 1 2 60117 40653
0 40655 5 1 1 40654
0 40656 7 1 2 42101 40655
0 40657 7 1 2 40649 40656
0 40658 5 1 1 40657
0 40659 7 1 2 46776 66512
0 40660 5 1 1 40659
0 40661 7 1 2 66567 40660
0 40662 5 1 1 40661
0 40663 7 1 2 42242 40662
0 40664 5 1 1 40663
0 40665 7 1 2 57750 70658
0 40666 5 1 1 40665
0 40667 7 1 2 40664 40666
0 40668 5 1 1 40667
0 40669 7 1 2 44506 40668
0 40670 5 1 1 40669
0 40671 7 1 2 59230 70965
0 40672 5 1 1 40671
0 40673 7 1 2 40670 40672
0 40674 5 2 1 40673
0 40675 7 2 2 49311 60114
0 40676 7 1 2 71693 71695
0 40677 5 1 1 40676
0 40678 7 1 2 61038 71068
0 40679 7 1 2 56167 40678
0 40680 5 1 1 40679
0 40681 7 1 2 40677 40680
0 40682 5 1 1 40681
0 40683 7 1 2 43485 40682
0 40684 5 1 1 40683
0 40685 7 1 2 65255 67225
0 40686 7 2 2 55634 58794
0 40687 7 1 2 68152 71697
0 40688 7 1 2 40685 40687
0 40689 5 1 1 40688
0 40690 7 1 2 40684 40689
0 40691 5 1 1 40690
0 40692 7 1 2 50439 40691
0 40693 5 1 1 40692
0 40694 7 1 2 50699 68278
0 40695 7 1 2 57031 40694
0 40696 7 1 2 63883 70442
0 40697 7 1 2 40695 40696
0 40698 5 1 1 40697
0 40699 7 1 2 40693 40698
0 40700 5 1 1 40699
0 40701 7 1 2 69537 40700
0 40702 5 1 1 40701
0 40703 7 1 2 46868 71694
0 40704 5 1 1 40703
0 40705 7 1 2 70143 71050
0 40706 5 1 1 40705
0 40707 7 1 2 40704 40706
0 40708 5 1 1 40707
0 40709 7 1 2 71696 40708
0 40710 5 1 1 40709
0 40711 7 1 2 60680 71069
0 40712 7 1 2 71692 40711
0 40713 5 1 1 40712
0 40714 7 1 2 40710 40713
0 40715 5 1 1 40714
0 40716 7 1 2 56050 66364
0 40717 7 1 2 40715 40716
0 40718 5 1 1 40717
0 40719 7 1 2 40702 40718
0 40720 5 1 1 40719
0 40721 7 1 2 47325 40720
0 40722 5 1 1 40721
0 40723 7 1 2 59432 64980
0 40724 5 1 1 40723
0 40725 7 2 2 48163 70646
0 40726 5 1 1 71699
0 40727 7 1 2 40724 40726
0 40728 5 1 1 40727
0 40729 7 1 2 65983 40728
0 40730 5 1 1 40729
0 40731 7 1 2 50142 50924
0 40732 7 1 2 69219 40731
0 40733 5 1 1 40732
0 40734 7 1 2 40730 40733
0 40735 5 1 1 40734
0 40736 7 1 2 51953 40735
0 40737 5 1 1 40736
0 40738 7 1 2 70745 71700
0 40739 5 1 1 40738
0 40740 7 1 2 40737 40739
0 40741 5 1 1 40740
0 40742 7 1 2 56784 57738
0 40743 7 1 2 67055 40742
0 40744 7 1 2 40741 40743
0 40745 5 1 1 40744
0 40746 7 1 2 45657 40745
0 40747 7 1 2 40722 40746
0 40748 5 1 1 40747
0 40749 7 1 2 46356 40748
0 40750 7 1 2 40658 40749
0 40751 5 1 1 40750
0 40752 7 1 2 52965 64469
0 40753 7 1 2 57443 40752
0 40754 7 1 2 59658 40753
0 40755 5 1 1 40754
0 40756 7 1 2 52127 52754
0 40757 7 1 2 58530 71037
0 40758 7 1 2 40756 40757
0 40759 5 1 1 40758
0 40760 7 1 2 40755 40759
0 40761 5 1 1 40760
0 40762 7 1 2 59317 40761
0 40763 5 1 1 40762
0 40764 7 1 2 5403 69690
0 40765 5 1 1 40764
0 40766 7 1 2 61174 64262
0 40767 7 1 2 70819 40766
0 40768 7 1 2 40765 40767
0 40769 5 1 1 40768
0 40770 7 1 2 40763 40769
0 40771 5 1 1 40770
0 40772 7 1 2 60488 70735
0 40773 7 1 2 40771 40772
0 40774 5 1 1 40773
0 40775 7 1 2 40751 40774
0 40776 5 1 1 40775
0 40777 7 1 2 45334 40776
0 40778 5 1 1 40777
0 40779 7 2 2 50920 54101
0 40780 7 1 2 69016 71701
0 40781 5 1 1 40780
0 40782 7 1 2 50967 61410
0 40783 7 1 2 64480 40782
0 40784 5 1 1 40783
0 40785 7 1 2 40781 40784
0 40786 5 2 1 40785
0 40787 7 1 2 51381 70996
0 40788 7 1 2 71703 40787
0 40789 5 1 1 40788
0 40790 7 1 2 49370 60298
0 40791 5 1 1 40790
0 40792 7 1 2 61892 69606
0 40793 7 1 2 40791 40792
0 40794 5 1 1 40793
0 40795 7 1 2 31894 40794
0 40796 5 1 1 40795
0 40797 7 1 2 47155 51647
0 40798 7 1 2 70794 40797
0 40799 7 1 2 40796 40798
0 40800 5 1 1 40799
0 40801 7 1 2 40789 40800
0 40802 5 1 1 40801
0 40803 7 1 2 45777 40802
0 40804 5 1 1 40803
0 40805 7 1 2 51382 64981
0 40806 7 1 2 64675 40805
0 40807 7 2 2 47326 60079
0 40808 7 1 2 70760 71705
0 40809 7 1 2 40806 40808
0 40810 5 1 1 40809
0 40811 7 1 2 40804 40810
0 40812 5 1 1 40811
0 40813 7 1 2 58161 40812
0 40814 5 1 1 40813
0 40815 7 1 2 64759 65368
0 40816 7 1 2 65512 71023
0 40817 7 1 2 40815 40816
0 40818 5 1 1 40817
0 40819 7 1 2 46777 63262
0 40820 7 2 2 68593 40819
0 40821 5 1 1 71707
0 40822 7 1 2 47327 50252
0 40823 7 1 2 61786 40822
0 40824 5 1 1 40823
0 40825 7 1 2 40821 40824
0 40826 5 1 1 40825
0 40827 7 1 2 56095 64007
0 40828 7 1 2 40826 40827
0 40829 5 1 1 40828
0 40830 7 1 2 40818 40829
0 40831 5 1 1 40830
0 40832 7 1 2 58264 58954
0 40833 7 1 2 60432 40832
0 40834 7 1 2 40831 40833
0 40835 5 1 1 40834
0 40836 7 1 2 40814 40835
0 40837 5 1 1 40836
0 40838 7 1 2 44601 40837
0 40839 5 1 1 40838
0 40840 7 1 2 48324 60681
0 40841 7 1 2 51575 40840
0 40842 7 1 2 62056 40841
0 40843 5 1 1 40842
0 40844 7 1 2 45778 44986
0 40845 7 1 2 60080 40844
0 40846 7 1 2 62330 40845
0 40847 7 1 2 69738 40846
0 40848 5 1 1 40847
0 40849 7 1 2 40843 40848
0 40850 5 1 1 40849
0 40851 7 1 2 45658 40850
0 40852 5 1 1 40851
0 40853 7 1 2 55174 59025
0 40854 7 1 2 69014 40853
0 40855 5 1 1 40854
0 40856 7 1 2 40852 40855
0 40857 5 1 1 40856
0 40858 7 1 2 45128 40857
0 40859 5 1 1 40858
0 40860 7 1 2 60685 68119
0 40861 7 1 2 56343 40860
0 40862 5 1 1 40861
0 40863 7 1 2 40859 40862
0 40864 5 1 1 40863
0 40865 7 1 2 44838 40864
0 40866 5 1 1 40865
0 40867 7 1 2 53972 56479
0 40868 7 1 2 61033 68296
0 40869 7 1 2 40867 40868
0 40870 5 1 1 40869
0 40871 7 1 2 40866 40870
0 40872 5 1 1 40871
0 40873 7 1 2 45874 40872
0 40874 5 1 1 40873
0 40875 7 1 2 61532 62638
0 40876 7 1 2 66416 40875
0 40877 7 1 2 67271 40876
0 40878 5 1 1 40877
0 40879 7 1 2 40874 40878
0 40880 5 1 1 40879
0 40881 7 1 2 45335 40880
0 40882 5 1 1 40881
0 40883 7 1 2 58637 61355
0 40884 7 1 2 63926 66081
0 40885 7 1 2 40883 40884
0 40886 5 1 1 40885
0 40887 7 1 2 40882 40886
0 40888 5 1 1 40887
0 40889 7 1 2 44507 57751
0 40890 7 1 2 40888 40889
0 40891 5 1 1 40890
0 40892 7 1 2 40839 40891
0 40893 5 1 1 40892
0 40894 7 1 2 67035 40893
0 40895 5 1 1 40894
0 40896 7 1 2 67291 67685
0 40897 7 1 2 70233 40896
0 40898 7 1 2 65866 67082
0 40899 7 1 2 68594 40898
0 40900 7 1 2 40897 40899
0 40901 5 1 1 40900
0 40902 7 1 2 56070 70843
0 40903 7 1 2 69625 40902
0 40904 5 1 1 40903
0 40905 7 1 2 44987 50700
0 40906 7 1 2 51108 40905
0 40907 7 1 2 62873 40906
0 40908 5 1 1 40907
0 40909 7 1 2 40904 40908
0 40910 5 1 1 40909
0 40911 7 1 2 42931 40910
0 40912 5 1 1 40911
0 40913 7 1 2 56078 70174
0 40914 7 1 2 59671 40913
0 40915 7 1 2 70773 40914
0 40916 5 1 1 40915
0 40917 7 1 2 40912 40916
0 40918 5 1 1 40917
0 40919 7 1 2 67841 70736
0 40920 7 1 2 40918 40919
0 40921 5 1 1 40920
0 40922 7 1 2 40901 40921
0 40923 5 1 1 40922
0 40924 7 1 2 49500 40923
0 40925 5 1 1 40924
0 40926 7 1 2 45875 71704
0 40927 5 1 1 40926
0 40928 7 1 2 51068 56826
0 40929 7 1 2 57139 40928
0 40930 7 1 2 69303 40929
0 40931 5 1 1 40930
0 40932 7 1 2 40927 40931
0 40933 5 1 1 40932
0 40934 7 1 2 58162 40933
0 40935 5 1 1 40934
0 40936 7 1 2 49810 58955
0 40937 7 1 2 57034 40936
0 40938 7 1 2 62574 70638
0 40939 7 1 2 40937 40938
0 40940 5 1 1 40939
0 40941 7 1 2 40935 40940
0 40942 5 1 1 40941
0 40943 7 1 2 50382 40942
0 40944 5 1 1 40943
0 40945 7 1 2 62078 63304
0 40946 7 1 2 69890 71698
0 40947 7 1 2 40945 40946
0 40948 5 1 1 40947
0 40949 7 1 2 40944 40948
0 40950 5 1 1 40949
0 40951 7 1 2 45336 40950
0 40952 5 1 1 40951
0 40953 7 1 2 58866 67892
0 40954 7 1 2 68280 40953
0 40955 7 1 2 71708 40954
0 40956 5 1 1 40955
0 40957 7 1 2 40952 40956
0 40958 5 1 1 40957
0 40959 7 1 2 44602 40958
0 40960 5 1 1 40959
0 40961 7 1 2 52909 54632
0 40962 5 1 1 40961
0 40963 7 1 2 54717 70918
0 40964 5 1 1 40963
0 40965 7 1 2 40962 40964
0 40966 5 1 1 40965
0 40967 7 1 2 51292 40966
0 40968 5 1 1 40967
0 40969 7 1 2 50143 69607
0 40970 7 1 2 71702 40969
0 40971 5 1 1 40970
0 40972 7 1 2 40968 40971
0 40973 5 1 1 40972
0 40974 7 1 2 43950 40973
0 40975 5 1 1 40974
0 40976 7 1 2 52170 59433
0 40977 7 1 2 65135 40976
0 40978 5 1 1 40977
0 40979 7 1 2 40975 40978
0 40980 5 1 1 40979
0 40981 7 1 2 58081 63030
0 40982 7 1 2 56436 40981
0 40983 7 1 2 40980 40982
0 40984 5 1 1 40983
0 40985 7 1 2 40960 40984
0 40986 5 1 1 40985
0 40987 7 1 2 53618 40986
0 40988 5 1 1 40987
0 40989 7 1 2 47328 49390
0 40990 7 1 2 61215 40989
0 40991 7 1 2 63675 66762
0 40992 7 1 2 70065 70827
0 40993 7 1 2 40991 40992
0 40994 7 1 2 40990 40993
0 40995 5 1 1 40994
0 40996 7 1 2 45876 40604
0 40997 5 1 1 40996
0 40998 7 1 2 42352 67228
0 40999 5 1 1 40998
0 41000 7 1 2 58571 40999
0 41001 7 1 2 40997 41000
0 41002 5 1 1 41001
0 41003 7 1 2 50232 68514
0 41004 7 1 2 60044 41003
0 41005 5 1 1 41004
0 41006 7 1 2 41002 41005
0 41007 5 1 1 41006
0 41008 7 1 2 46357 41007
0 41009 5 1 1 41008
0 41010 7 1 2 55528 64722
0 41011 7 1 2 56116 41010
0 41012 7 1 2 69619 41011
0 41013 5 1 1 41012
0 41014 7 1 2 41009 41013
0 41015 5 1 1 41014
0 41016 7 1 2 47471 41015
0 41017 5 1 1 41016
0 41018 7 1 2 51845 54239
0 41019 7 1 2 68458 41018
0 41020 7 1 2 51421 60045
0 41021 7 1 2 41019 41020
0 41022 5 1 1 41021
0 41023 7 1 2 41017 41022
0 41024 5 1 1 41023
0 41025 7 1 2 50440 57463
0 41026 7 1 2 58142 41025
0 41027 7 1 2 41024 41026
0 41028 5 1 1 41027
0 41029 7 1 2 40995 41028
0 41030 7 1 2 40988 41029
0 41031 5 1 1 41030
0 41032 7 1 2 66285 41031
0 41033 5 1 1 41032
0 41034 7 1 2 40925 41033
0 41035 7 1 2 40895 41034
0 41036 7 1 2 40778 41035
0 41037 5 1 1 41036
0 41038 7 1 2 47701 41037
0 41039 5 1 1 41038
0 41040 7 1 2 52171 64960
0 41041 7 1 2 71644 41040
0 41042 7 1 2 69659 41041
0 41043 5 1 1 41042
0 41044 7 2 2 52456 53049
0 41045 7 1 2 59130 69671
0 41046 7 1 2 71709 41045
0 41047 5 1 1 41046
0 41048 7 1 2 41043 41047
0 41049 5 1 1 41048
0 41050 7 1 2 45659 41049
0 41051 5 1 1 41050
0 41052 7 1 2 51648 67159
0 41053 7 1 2 71710 41052
0 41054 5 1 1 41053
0 41055 7 1 2 41051 41054
0 41056 5 1 1 41055
0 41057 7 1 2 43951 41056
0 41058 5 1 1 41057
0 41059 7 2 2 43405 52491
0 41060 5 1 1 71711
0 41061 7 1 2 49830 41060
0 41062 5 1 1 41061
0 41063 7 1 2 43180 24505
0 41064 5 1 1 41063
0 41065 7 1 2 57216 41064
0 41066 7 1 2 41062 41065
0 41067 7 1 2 67173 41066
0 41068 5 1 1 41067
0 41069 7 1 2 41058 41068
0 41070 5 1 1 41069
0 41071 7 1 2 47927 41070
0 41072 5 1 1 41071
0 41073 7 1 2 67713 69323
0 41074 5 1 1 41073
0 41075 7 1 2 51089 68646
0 41076 7 1 2 68549 41075
0 41077 5 1 1 41076
0 41078 7 1 2 41074 41077
0 41079 5 1 1 41078
0 41080 7 1 2 70135 41079
0 41081 5 1 1 41080
0 41082 7 1 2 41072 41081
0 41083 5 1 1 41082
0 41084 7 1 2 66323 41083
0 41085 5 1 1 41084
0 41086 7 2 2 56286 57868
0 41087 7 1 2 71712 71713
0 41088 5 1 1 41087
0 41089 7 2 2 66591 68550
0 41090 7 1 2 69714 71715
0 41091 5 1 1 41090
0 41092 7 1 2 41088 41091
0 41093 5 1 1 41092
0 41094 7 1 2 46358 41093
0 41095 5 1 1 41094
0 41096 7 1 2 52457 57752
0 41097 7 2 2 56287 41096
0 41098 7 1 2 57144 71717
0 41099 5 1 1 41098
0 41100 7 1 2 41095 41099
0 41101 5 1 1 41100
0 41102 7 1 2 51044 41101
0 41103 5 1 1 41102
0 41104 7 1 2 56150 71718
0 41105 5 1 1 41104
0 41106 7 1 2 53711 71716
0 41107 5 1 1 41106
0 41108 7 1 2 70919 71714
0 41109 5 1 1 41108
0 41110 7 1 2 41107 41109
0 41111 5 1 1 41110
0 41112 7 1 2 61613 41111
0 41113 5 1 1 41112
0 41114 7 1 2 41105 41113
0 41115 7 1 2 41103 41114
0 41116 5 1 1 41115
0 41117 7 1 2 48164 41116
0 41118 5 1 1 41117
0 41119 7 1 2 55389 57262
0 41120 7 1 2 69318 41119
0 41121 7 1 2 53712 41120
0 41122 5 1 1 41121
0 41123 7 1 2 41118 41122
0 41124 5 1 1 41123
0 41125 7 1 2 43606 69397
0 41126 7 1 2 41124 41125
0 41127 5 1 1 41126
0 41128 7 1 2 41085 41127
0 41129 5 1 1 41128
0 41130 7 1 2 44696 41129
0 41131 5 1 1 41130
0 41132 7 2 2 45129 60042
0 41133 7 2 2 52755 71719
0 41134 7 1 2 55642 57020
0 41135 7 2 2 71721 41134
0 41136 5 1 1 71723
0 41137 7 1 2 42243 71724
0 41138 5 1 1 41137
0 41139 7 1 2 43406 68917
0 41140 5 1 1 41139
0 41141 7 1 2 65402 41140
0 41142 5 2 1 41141
0 41143 7 3 2 55823 71725
0 41144 7 1 2 53619 71727
0 41145 5 1 1 41144
0 41146 7 1 2 41138 41145
0 41147 5 1 1 41146
0 41148 7 1 2 54485 41147
0 41149 5 1 1 41148
0 41150 7 1 2 53620 55824
0 41151 5 1 1 41150
0 41152 7 1 2 33455 41151
0 41153 5 1 1 41152
0 41154 7 1 2 46869 41153
0 41155 5 1 1 41154
0 41156 7 1 2 53662 66592
0 41157 5 1 1 41156
0 41158 7 1 2 41155 41157
0 41159 5 1 1 41158
0 41160 7 1 2 65400 41159
0 41161 5 1 1 41160
0 41162 7 1 2 51052 55675
0 41163 7 1 2 68287 41162
0 41164 7 1 2 69853 41163
0 41165 5 1 1 41164
0 41166 7 1 2 41161 41165
0 41167 5 1 1 41166
0 41168 7 1 2 42102 41167
0 41169 5 1 1 41168
0 41170 7 1 2 41149 41169
0 41171 5 1 1 41170
0 41172 7 1 2 48325 41171
0 41173 5 1 1 41172
0 41174 7 1 2 54979 56997
0 41175 7 2 2 69134 41174
0 41176 7 1 2 49391 56288
0 41177 7 1 2 71730 41176
0 41178 5 1 1 41177
0 41179 7 1 2 41173 41178
0 41180 5 1 1 41179
0 41181 7 1 2 68164 41180
0 41182 5 1 1 41181
0 41183 7 1 2 69273 71728
0 41184 5 1 1 41183
0 41185 7 1 2 46949 71729
0 41186 5 1 1 41185
0 41187 7 1 2 41136 41186
0 41188 5 1 1 41187
0 41189 7 1 2 45779 41188
0 41190 5 1 1 41189
0 41191 7 1 2 58037 71722
0 41192 5 1 1 41191
0 41193 7 1 2 41190 41192
0 41194 5 1 1 41193
0 41195 7 1 2 48915 41194
0 41196 5 1 1 41195
0 41197 7 1 2 41184 41196
0 41198 5 1 1 41197
0 41199 7 1 2 48326 41198
0 41200 5 1 1 41199
0 41201 7 1 2 49392 71731
0 41202 7 1 2 53713 41201
0 41203 5 1 1 41202
0 41204 7 1 2 41200 41203
0 41205 5 1 1 41204
0 41206 7 1 2 66346 41205
0 41207 5 1 1 41206
0 41208 7 1 2 41182 41207
0 41209 5 1 1 41208
0 41210 7 1 2 59685 41209
0 41211 5 1 1 41210
0 41212 7 1 2 41131 41211
0 41213 5 1 1 41212
0 41214 7 1 2 47827 41213
0 41215 5 1 1 41214
0 41216 7 1 2 63104 70124
0 41217 7 1 2 67557 41216
0 41218 5 1 1 41217
0 41219 7 1 2 51693 69275
0 41220 7 1 2 51090 41219
0 41221 5 1 1 41220
0 41222 7 1 2 41218 41221
0 41223 5 1 1 41222
0 41224 7 1 2 53811 41223
0 41225 5 1 1 41224
0 41226 7 1 2 46359 64744
0 41227 5 1 1 41226
0 41228 7 1 2 54436 65534
0 41229 7 1 2 41227 41228
0 41230 5 1 1 41229
0 41231 7 1 2 41225 41230
0 41232 5 1 1 41231
0 41233 7 1 2 45130 41232
0 41234 5 1 1 41233
0 41235 7 2 2 46778 66441
0 41236 7 1 2 46995 56396
0 41237 7 1 2 71732 41236
0 41238 7 1 2 53051 41237
0 41239 5 1 1 41238
0 41240 7 1 2 41234 41239
0 41241 5 1 1 41240
0 41242 7 1 2 66390 41241
0 41243 5 1 1 41242
0 41244 7 1 2 52107 53077
0 41245 5 1 1 41244
0 41246 7 3 2 69708 41245
0 41247 7 1 2 57265 71734
0 41248 5 1 1 41247
0 41249 7 1 2 58741 70125
0 41250 7 1 2 65311 41249
0 41251 5 1 1 41250
0 41252 7 1 2 41248 41251
0 41253 5 1 1 41252
0 41254 7 1 2 66669 66241
0 41255 7 1 2 41253 41254
0 41256 5 1 1 41255
0 41257 7 1 2 41243 41256
0 41258 5 1 1 41257
0 41259 7 1 2 42353 41258
0 41260 5 1 1 41259
0 41261 7 1 2 57753 67036
0 41262 7 1 2 71735 41261
0 41263 5 1 1 41262
0 41264 7 1 2 66043 70175
0 41265 7 1 2 67125 41264
0 41266 7 1 2 70920 41265
0 41267 5 1 1 41266
0 41268 7 1 2 41263 41267
0 41269 5 1 1 41268
0 41270 7 1 2 65984 41269
0 41271 5 1 1 41270
0 41272 7 1 2 41260 41271
0 41273 5 1 1 41272
0 41274 7 1 2 42244 41273
0 41275 5 1 1 41274
0 41276 7 1 2 56616 61207
0 41277 7 2 2 68165 41276
0 41278 7 1 2 71736 71737
0 41279 5 1 1 41278
0 41280 7 1 2 41275 41279
0 41281 5 1 1 41280
0 41282 7 1 2 47329 41281
0 41283 5 1 1 41282
0 41284 7 1 2 52720 57266
0 41285 5 1 1 41284
0 41286 7 1 2 37596 41285
0 41287 5 1 1 41286
0 41288 7 1 2 68166 41287
0 41289 5 1 1 41288
0 41290 7 1 2 66347 68319
0 41291 7 1 2 71549 41290
0 41292 5 1 1 41291
0 41293 7 1 2 41289 41292
0 41294 5 1 1 41293
0 41295 7 1 2 48040 41294
0 41296 5 1 1 41295
0 41297 7 1 2 55449 69528
0 41298 5 1 1 41297
0 41299 7 1 2 41296 41298
0 41300 5 1 1 41299
0 41301 7 1 2 42245 41300
0 41302 5 1 1 41301
0 41303 7 1 2 52721 71738
0 41304 5 1 1 41303
0 41305 7 1 2 41302 41304
0 41306 5 1 1 41305
0 41307 7 1 2 47472 41306
0 41308 5 1 1 41307
0 41309 7 1 2 49923 70947
0 41310 7 1 2 69824 41309
0 41311 5 1 1 41310
0 41312 7 1 2 41308 41311
0 41313 5 1 1 41312
0 41314 7 1 2 44988 53072
0 41315 7 1 2 41313 41314
0 41316 5 1 1 41315
0 41317 7 1 2 41283 41316
0 41318 5 1 1 41317
0 41319 7 1 2 48165 41318
0 41320 5 1 1 41319
0 41321 7 1 2 48949 52172
0 41322 7 1 2 53023 41321
0 41323 7 1 2 59245 41322
0 41324 7 1 2 69289 41323
0 41325 5 1 1 41324
0 41326 7 1 2 41320 41325
0 41327 5 1 1 41326
0 41328 7 1 2 65665 41327
0 41329 5 1 1 41328
0 41330 7 1 2 41215 41329
0 41331 5 1 1 41330
0 41332 7 1 2 53298 41331
0 41333 5 1 1 41332
0 41334 7 2 2 64053 71612
0 41335 7 1 2 70715 71739
0 41336 5 1 1 41335
0 41337 7 1 2 42354 50900
0 41338 5 1 1 41337
0 41339 7 1 2 51550 66513
0 41340 5 1 1 41339
0 41341 7 1 2 41338 41340
0 41342 5 1 1 41341
0 41343 7 1 2 46779 41342
0 41344 5 1 1 41343
0 41345 7 1 2 61012 64490
0 41346 5 1 1 41345
0 41347 7 1 2 41344 41346
0 41348 5 1 1 41347
0 41349 7 1 2 47473 41348
0 41350 5 1 1 41349
0 41351 7 1 2 58401 68430
0 41352 7 1 2 51054 41351
0 41353 5 1 1 41352
0 41354 7 1 2 41350 41353
0 41355 5 1 1 41354
0 41356 7 1 2 67213 41355
0 41357 5 1 1 41356
0 41358 7 1 2 41336 41357
0 41359 5 1 1 41358
0 41360 7 1 2 46574 41359
0 41361 5 1 1 41360
0 41362 7 1 2 56304 65099
0 41363 7 1 2 70938 71024
0 41364 7 1 2 41362 41363
0 41365 5 1 1 41364
0 41366 7 1 2 41361 41365
0 41367 5 1 1 41366
0 41368 7 1 2 46360 41367
0 41369 5 1 1 41368
0 41370 7 1 2 43181 58655
0 41371 5 1 1 41370
0 41372 7 1 2 54736 54902
0 41373 5 1 1 41372
0 41374 7 1 2 41371 41373
0 41375 5 1 1 41374
0 41376 7 1 2 71740 41375
0 41377 5 1 1 41376
0 41378 7 1 2 41369 41377
0 41379 5 1 1 41378
0 41380 7 1 2 53714 41379
0 41381 5 1 1 41380
0 41382 7 1 2 46780 70079
0 41383 5 1 1 41382
0 41384 7 1 2 70072 70948
0 41385 5 1 1 41384
0 41386 7 1 2 41383 41385
0 41387 5 1 1 41386
0 41388 7 1 2 42103 41387
0 41389 5 1 1 41388
0 41390 7 1 2 64651 70949
0 41391 5 1 1 41390
0 41392 7 1 2 41389 41391
0 41393 5 1 1 41392
0 41394 7 1 2 68977 41393
0 41395 5 1 1 41394
0 41396 7 1 2 44697 55837
0 41397 7 1 2 69596 41396
0 41398 5 1 1 41397
0 41399 7 1 2 43182 54466
0 41400 7 1 2 62137 41399
0 41401 7 1 2 70419 41400
0 41402 5 1 1 41401
0 41403 7 1 2 41398 41402
0 41404 5 1 1 41403
0 41405 7 1 2 70709 41404
0 41406 5 1 1 41405
0 41407 7 1 2 69597 71480
0 41408 5 1 1 41407
0 41409 7 1 2 55446 57894
0 41410 7 1 2 70420 41409
0 41411 5 1 1 41410
0 41412 7 1 2 41408 41411
0 41413 5 1 1 41412
0 41414 7 1 2 68974 41413
0 41415 5 1 1 41414
0 41416 7 1 2 41406 41415
0 41417 7 1 2 41395 41416
0 41418 5 1 1 41417
0 41419 7 1 2 51322 41418
0 41420 5 1 1 41419
0 41421 7 1 2 56543 71646
0 41422 5 1 1 41421
0 41423 7 1 2 58774 62212
0 41424 5 1 1 41423
0 41425 7 1 2 41422 41424
0 41426 5 1 1 41425
0 41427 7 1 2 42355 41426
0 41428 5 1 1 41427
0 41429 7 1 2 65837 66593
0 41430 7 1 2 61383 41429
0 41431 5 1 1 41430
0 41432 7 1 2 41428 41431
0 41433 5 1 1 41432
0 41434 7 1 2 42104 41433
0 41435 5 1 1 41434
0 41436 7 1 2 56544 63031
0 41437 7 1 2 61789 41436
0 41438 5 1 1 41437
0 41439 7 1 2 41435 41438
0 41440 5 1 1 41439
0 41441 7 1 2 49312 41440
0 41442 5 1 1 41441
0 41443 7 1 2 42356 5790
0 41444 5 1 1 41443
0 41445 7 1 2 45877 61366
0 41446 5 1 1 41445
0 41447 7 1 2 54688 66594
0 41448 7 1 2 41446 41447
0 41449 7 1 2 41444 41448
0 41450 5 1 1 41449
0 41451 7 1 2 41442 41450
0 41452 5 1 1 41451
0 41453 7 1 2 53411 54601
0 41454 7 1 2 41452 41453
0 41455 5 1 1 41454
0 41456 7 1 2 41420 41455
0 41457 5 1 1 41456
0 41458 7 1 2 53621 41457
0 41459 5 1 1 41458
0 41460 7 1 2 41381 41459
0 41461 5 1 1 41460
0 41462 7 1 2 47828 41461
0 41463 5 1 1 41462
0 41464 7 1 2 2957 67217
0 41465 5 1 1 41464
0 41466 7 1 2 42357 41465
0 41467 5 1 1 41466
0 41468 7 1 2 67256 27921
0 41469 5 2 1 41468
0 41470 7 1 2 66578 71741
0 41471 5 1 1 41470
0 41472 7 1 2 41467 41471
0 41473 5 1 1 41472
0 41474 7 1 2 43566 41473
0 41475 5 1 1 41474
0 41476 7 1 2 56480 71569
0 41477 5 1 1 41476
0 41478 7 1 2 41475 41477
0 41479 5 1 1 41478
0 41480 7 1 2 42246 41479
0 41481 5 1 1 41480
0 41482 7 1 2 56160 68320
0 41483 7 1 2 70932 41482
0 41484 5 1 1 41483
0 41485 7 1 2 41481 41484
0 41486 5 1 1 41485
0 41487 7 1 2 52080 41486
0 41488 5 1 1 41487
0 41489 7 1 2 59659 69583
0 41490 5 1 1 41489
0 41491 7 1 2 56161 71733
0 41492 5 1 1 41491
0 41493 7 1 2 41490 41492
0 41494 5 1 1 41493
0 41495 7 1 2 42247 41494
0 41496 5 1 1 41495
0 41497 7 1 2 45780 68321
0 41498 7 1 2 56481 41497
0 41499 5 1 1 41498
0 41500 7 1 2 41496 41499
0 41501 5 1 1 41500
0 41502 7 1 2 42358 41501
0 41503 5 1 1 41502
0 41504 7 1 2 56254 63746
0 41505 7 1 2 67246 41504
0 41506 5 1 1 41505
0 41507 7 1 2 41503 41506
0 41508 5 1 1 41507
0 41509 7 1 2 71172 41508
0 41510 5 1 1 41509
0 41511 7 1 2 41488 41510
0 41512 5 1 1 41511
0 41513 7 1 2 46361 41512
0 41514 5 1 1 41513
0 41515 7 1 2 44603 59243
0 41516 5 1 1 41515
0 41517 7 1 2 43183 57267
0 41518 5 1 1 41517
0 41519 7 1 2 41516 41518
0 41520 5 1 1 41519
0 41521 7 1 2 42248 41520
0 41522 5 1 1 41521
0 41523 7 1 2 51827 68322
0 41524 5 1 1 41523
0 41525 7 1 2 41522 41524
0 41526 5 1 1 41525
0 41527 7 1 2 65508 41526
0 41528 5 1 1 41527
0 41529 7 2 2 49501 54680
0 41530 7 1 2 58674 71743
0 41531 5 1 1 41530
0 41532 7 1 2 41528 41531
0 41533 5 1 1 41532
0 41534 7 1 2 42932 41533
0 41535 5 1 1 41534
0 41536 7 1 2 53128 60262
0 41537 7 1 2 59246 41536
0 41538 5 1 1 41537
0 41539 7 1 2 41535 41538
0 41540 5 1 1 41539
0 41541 7 1 2 51257 69565
0 41542 7 1 2 41540 41541
0 41543 5 1 1 41542
0 41544 7 1 2 41514 41543
0 41545 5 1 1 41544
0 41546 7 1 2 47156 41545
0 41547 5 1 1 41546
0 41548 7 1 2 56096 64123
0 41549 7 1 2 69192 41548
0 41550 7 1 2 71013 71273
0 41551 7 1 2 41549 41550
0 41552 5 1 1 41551
0 41553 7 1 2 41547 41552
0 41554 5 1 1 41553
0 41555 7 1 2 46103 41554
0 41556 5 1 1 41555
0 41557 7 2 2 49663 56144
0 41558 7 1 2 64280 71745
0 41559 5 1 1 41558
0 41560 7 1 2 54139 68628
0 41561 5 2 1 41560
0 41562 7 1 2 41559 71747
0 41563 5 1 1 41562
0 41564 7 1 2 64729 41563
0 41565 5 1 1 41564
0 41566 7 1 2 52655 64952
0 41567 5 1 1 41566
0 41568 7 1 2 2290 41567
0 41569 5 1 1 41568
0 41570 7 1 2 55291 58099
0 41571 7 1 2 41569 41570
0 41572 5 2 1 41571
0 41573 7 1 2 41565 71749
0 41574 5 1 1 41573
0 41575 7 1 2 71168 41574
0 41576 5 1 1 41575
0 41577 7 1 2 41556 41576
0 41578 5 1 1 41577
0 41579 7 1 2 48925 41578
0 41580 5 1 1 41579
0 41581 7 1 2 41463 41580
0 41582 5 1 1 41581
0 41583 7 1 2 66286 41582
0 41584 5 1 1 41583
0 41585 7 1 2 68978 70336
0 41586 5 1 1 41585
0 41587 7 1 2 65190 65237
0 41588 5 1 1 41587
0 41589 7 1 2 65783 41588
0 41590 5 1 1 41589
0 41591 7 1 2 48487 62068
0 41592 7 1 2 65513 41591
0 41593 5 1 1 41592
0 41594 7 1 2 41590 41593
0 41595 5 1 1 41594
0 41596 7 1 2 48327 41595
0 41597 5 1 1 41596
0 41598 7 1 2 52708 69161
0 41599 7 1 2 69774 41598
0 41600 5 1 1 41599
0 41601 7 1 2 41597 41600
0 41602 5 1 1 41601
0 41603 7 1 2 51305 41602
0 41604 5 1 1 41603
0 41605 7 1 2 41586 41604
0 41606 5 1 1 41605
0 41607 7 1 2 43407 41606
0 41608 5 1 1 41607
0 41609 7 1 2 62097 71035
0 41610 7 1 2 50480 19960
0 41611 5 1 1 41610
0 41612 7 1 2 51190 33141
0 41613 5 1 1 41612
0 41614 7 1 2 41611 41613
0 41615 7 1 2 41609 41614
0 41616 5 1 1 41615
0 41617 7 1 2 41608 41616
0 41618 5 1 1 41617
0 41619 7 1 2 45337 41618
0 41620 5 1 1 41619
0 41621 7 1 2 55024 70149
0 41622 5 1 1 41621
0 41623 7 1 2 46104 49475
0 41624 7 1 2 53479 57250
0 41625 7 1 2 41623 41624
0 41626 5 1 1 41625
0 41627 7 1 2 41622 41626
0 41628 5 1 1 41627
0 41629 7 1 2 65784 69135
0 41630 7 1 2 41628 41629
0 41631 5 1 1 41630
0 41632 7 1 2 41620 41631
0 41633 5 1 1 41632
0 41634 7 1 2 55013 41633
0 41635 5 1 1 41634
0 41636 7 1 2 54518 56827
0 41637 7 2 2 52443 41636
0 41638 7 1 2 55194 69598
0 41639 7 1 2 71751 41638
0 41640 5 1 1 41639
0 41641 7 1 2 41635 41640
0 41642 5 1 1 41641
0 41643 7 1 2 42249 41642
0 41644 5 1 1 41643
0 41645 7 1 2 43782 68629
0 41646 5 1 1 41645
0 41647 7 1 2 50441 67226
0 41648 5 1 1 41647
0 41649 7 1 2 41646 41648
0 41650 5 1 1 41649
0 41651 7 1 2 44698 41650
0 41652 5 1 1 41651
0 41653 7 1 2 50442 67254
0 41654 5 1 1 41653
0 41655 7 1 2 41652 41654
0 41656 5 1 1 41655
0 41657 7 1 2 64723 41656
0 41658 5 1 1 41657
0 41659 7 1 2 64491 67215
0 41660 5 1 1 41659
0 41661 7 1 2 41658 41660
0 41662 5 1 1 41661
0 41663 7 1 2 51091 41662
0 41664 5 1 1 41663
0 41665 7 1 2 48950 64106
0 41666 7 1 2 57690 41665
0 41667 7 1 2 67850 41666
0 41668 5 1 1 41667
0 41669 7 1 2 41664 41668
0 41670 5 1 1 41669
0 41671 7 1 2 46362 41670
0 41672 5 1 1 41671
0 41673 7 1 2 68235 70803
0 41674 7 1 2 51323 41673
0 41675 7 1 2 69319 41674
0 41676 5 1 1 41675
0 41677 7 1 2 41672 41676
0 41678 5 1 1 41677
0 41679 7 1 2 42105 71091
0 41680 7 1 2 41678 41679
0 41681 5 1 1 41680
0 41682 7 1 2 41644 41681
0 41683 5 1 1 41682
0 41684 7 1 2 47829 41683
0 41685 5 1 1 41684
0 41686 7 1 2 42359 71742
0 41687 5 1 1 41686
0 41688 7 1 2 56162 69764
0 41689 5 1 1 41688
0 41690 7 1 2 41687 41689
0 41691 5 1 1 41690
0 41692 7 1 2 52081 41691
0 41693 5 1 1 41692
0 41694 7 2 2 46575 62069
0 41695 7 1 2 56163 64031
0 41696 5 1 1 41695
0 41697 7 1 2 54602 70997
0 41698 5 1 1 41697
0 41699 7 1 2 41696 41698
0 41700 5 1 1 41699
0 41701 7 1 2 71753 41700
0 41702 5 1 1 41701
0 41703 7 1 2 41693 41702
0 41704 5 1 1 41703
0 41705 7 1 2 46363 41704
0 41706 5 1 1 41705
0 41707 7 1 2 56598 69765
0 41708 7 1 2 70713 41707
0 41709 5 1 1 41708
0 41710 7 1 2 41706 41709
0 41711 5 1 1 41710
0 41712 7 1 2 43486 50485
0 41713 7 1 2 61770 41712
0 41714 7 1 2 41711 41713
0 41715 5 1 1 41714
0 41716 7 1 2 41685 41715
0 41717 5 1 1 41716
0 41718 7 1 2 67037 41717
0 41719 5 1 1 41718
0 41720 7 1 2 50921 62203
0 41721 7 1 2 71746 41720
0 41722 5 1 1 41721
0 41723 7 1 2 71748 41722
0 41724 5 1 1 41723
0 41725 7 1 2 64730 41724
0 41726 5 1 1 41725
0 41727 7 1 2 71750 41726
0 41728 5 1 1 41727
0 41729 7 1 2 65985 41728
0 41730 5 1 1 41729
0 41731 7 1 2 50481 52601
0 41732 7 1 2 57282 64124
0 41733 7 1 2 41731 41732
0 41734 7 1 2 51191 51352
0 41735 5 1 1 41734
0 41736 7 1 2 62285 41735
0 41737 7 1 2 41733 41736
0 41738 5 1 1 41737
0 41739 7 1 2 41730 41738
0 41740 5 1 1 41739
0 41741 7 1 2 59318 41740
0 41742 5 1 1 41741
0 41743 7 1 2 51954 69768
0 41744 5 1 1 41743
0 41745 7 1 2 71143 41744
0 41746 5 1 1 41745
0 41747 7 2 2 45338 41746
0 41748 5 1 1 71755
0 41749 7 1 2 70074 70966
0 41750 5 1 1 41749
0 41751 7 1 2 41748 41750
0 41752 5 1 1 41751
0 41753 7 1 2 53073 41752
0 41754 5 1 1 41753
0 41755 7 1 2 47474 70970
0 41756 5 1 1 41755
0 41757 7 1 2 41754 41756
0 41758 5 1 1 41757
0 41759 7 1 2 46576 54550
0 41760 7 1 2 41758 41759
0 41761 5 1 1 41760
0 41762 7 1 2 55348 71756
0 41763 5 1 1 41762
0 41764 7 1 2 48328 41763
0 41765 7 1 2 41761 41764
0 41766 5 1 1 41765
0 41767 7 1 2 71045 71744
0 41768 5 1 1 41767
0 41769 7 1 2 43408 71141
0 41770 5 1 1 41769
0 41771 7 1 2 51573 61208
0 41772 7 1 2 63224 41771
0 41773 5 1 1 41772
0 41774 7 1 2 41770 41773
0 41775 5 1 1 41774
0 41776 7 1 2 65509 41775
0 41777 5 1 1 41776
0 41778 7 1 2 41768 41777
0 41779 5 1 1 41778
0 41780 7 1 2 42933 41779
0 41781 5 1 1 41780
0 41782 7 1 2 69221 70746
0 41783 5 1 1 41782
0 41784 7 1 2 44989 41783
0 41785 7 1 2 41781 41784
0 41786 5 1 1 41785
0 41787 7 1 2 48166 41786
0 41788 7 1 2 41766 41787
0 41789 5 1 1 41788
0 41790 7 1 2 53790 69885
0 41791 7 1 2 70934 41790
0 41792 5 1 1 41791
0 41793 7 1 2 41789 41792
0 41794 5 1 1 41793
0 41795 7 1 2 46105 41794
0 41796 5 1 1 41795
0 41797 7 1 2 54980 69611
0 41798 5 1 1 41797
0 41799 7 1 2 44990 62138
0 41800 7 1 2 64320 41799
0 41801 5 1 1 41800
0 41802 7 1 2 41798 41801
0 41803 5 1 1 41802
0 41804 7 1 2 59558 62204
0 41805 7 1 2 71720 41804
0 41806 7 1 2 41803 41805
0 41807 5 1 1 41806
0 41808 7 1 2 41796 41807
0 41809 5 1 1 41808
0 41810 7 1 2 47157 41809
0 41811 5 1 1 41810
0 41812 7 1 2 41742 41811
0 41813 5 1 1 41812
0 41814 7 1 2 67336 41813
0 41815 5 1 1 41814
0 41816 7 1 2 52722 64765
0 41817 5 1 1 41816
0 41818 7 1 2 55825 63884
0 41819 5 1 1 41818
0 41820 7 1 2 41817 41819
0 41821 5 1 1 41820
0 41822 7 1 2 53812 41821
0 41823 5 1 1 41822
0 41824 7 1 2 49801 62867
0 41825 7 1 2 64992 41824
0 41826 5 1 1 41825
0 41827 7 1 2 41823 41826
0 41828 5 1 1 41827
0 41829 7 1 2 47475 41828
0 41830 5 1 1 41829
0 41831 7 1 2 49828 54981
0 41832 5 1 1 41831
0 41833 7 1 2 70681 41832
0 41834 5 1 1 41833
0 41835 7 1 2 64766 41834
0 41836 5 1 1 41835
0 41837 7 1 2 41830 41836
0 41838 5 1 1 41837
0 41839 7 1 2 48488 41838
0 41840 5 1 1 41839
0 41841 7 1 2 56785 59319
0 41842 7 1 2 70679 41841
0 41843 5 1 1 41842
0 41844 7 1 2 57869 64961
0 41845 7 1 2 70921 41844
0 41846 5 1 1 41845
0 41847 7 1 2 41843 41846
0 41848 5 1 1 41847
0 41849 7 1 2 42934 41848
0 41850 5 1 1 41849
0 41851 7 1 2 41840 41850
0 41852 5 1 1 41851
0 41853 7 1 2 50443 41852
0 41854 5 1 1 41853
0 41855 7 1 2 51092 59320
0 41856 5 1 1 41855
0 41857 7 1 2 45781 71173
0 41858 5 1 1 41857
0 41859 7 1 2 41856 41858
0 41860 5 1 1 41859
0 41861 7 1 2 55109 58436
0 41862 7 1 2 54603 41861
0 41863 7 1 2 41860 41862
0 41864 5 1 1 41863
0 41865 7 1 2 41854 41864
0 41866 5 1 1 41865
0 41867 7 1 2 48167 41866
0 41868 5 1 1 41867
0 41869 7 1 2 42250 54429
0 41870 7 1 2 60143 41869
0 41871 7 1 2 70685 41870
0 41872 5 1 1 41871
0 41873 7 1 2 41868 41872
0 41874 5 1 1 41873
0 41875 7 1 2 44699 41874
0 41876 5 1 1 41875
0 41877 7 1 2 60962 71539
0 41878 5 1 1 41877
0 41879 7 1 2 64760 65613
0 41880 5 1 1 41879
0 41881 7 1 2 41878 41880
0 41882 5 1 1 41881
0 41883 7 1 2 55056 67247
0 41884 7 1 2 41882 41883
0 41885 5 1 1 41884
0 41886 7 1 2 42360 41885
0 41887 7 1 2 41876 41886
0 41888 5 1 1 41887
0 41889 7 1 2 56145 60920
0 41890 7 1 2 69775 41889
0 41891 5 1 1 41890
0 41892 7 1 2 42251 57023
0 41893 7 1 2 65030 41892
0 41894 5 1 1 41893
0 41895 7 1 2 41891 41894
0 41896 5 1 1 41895
0 41897 7 1 2 50444 41896
0 41898 5 1 1 41897
0 41899 7 1 2 51161 58892
0 41900 7 1 2 71726 41899
0 41901 5 1 1 41900
0 41902 7 1 2 41898 41901
0 41903 5 1 1 41902
0 41904 7 1 2 44991 41903
0 41905 5 1 1 41904
0 41906 7 1 2 70158 71754
0 41907 7 1 2 51325 41906
0 41908 5 1 1 41907
0 41909 7 1 2 41905 41908
0 41910 5 1 1 41909
0 41911 7 1 2 45339 41910
0 41912 5 1 1 41911
0 41913 7 1 2 58531 60115
0 41914 7 1 2 69196 71706
0 41915 7 1 2 41913 41914
0 41916 5 1 1 41915
0 41917 7 1 2 41912 41916
0 41918 5 1 1 41917
0 41919 7 1 2 47928 41918
0 41920 5 1 1 41919
0 41921 7 1 2 44992 60968
0 41922 7 1 2 51110 41921
0 41923 7 1 2 55025 71059
0 41924 7 1 2 41922 41923
0 41925 5 1 1 41924
0 41926 7 1 2 45878 41925
0 41927 7 1 2 41920 41926
0 41928 5 1 1 41927
0 41929 7 1 2 69344 41928
0 41930 7 1 2 41888 41929
0 41931 5 1 1 41930
0 41932 7 1 2 61107 63984
0 41933 7 1 2 69245 41932
0 41934 7 1 2 71752 41933
0 41935 5 1 1 41934
0 41936 7 1 2 41931 41935
0 41937 5 1 1 41936
0 41938 7 1 2 47830 41937
0 41939 5 1 1 41938
0 41940 7 1 2 41815 41939
0 41941 7 1 2 41719 41940
0 41942 7 1 2 41584 41941
0 41943 5 1 1 41942
0 41944 7 1 2 44371 41943
0 41945 5 1 1 41944
0 41946 7 1 2 41333 41945
0 41947 7 1 2 41039 41946
0 41948 5 1 1 41947
0 41949 7 1 2 49100 41948
0 41950 5 1 1 41949
0 41951 7 1 2 40594 41950
0 41952 7 1 2 35118 41951
0 41953 7 1 2 28035 41952
0 41954 7 1 2 24695 41953
0 41955 7 1 2 24062 41954
0 41956 7 1 2 22335 41955
0 41957 7 1 2 17013 41956
3 89999 5 0 1 41957
