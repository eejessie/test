1 0 0 68 0
2 25 1 0
2 26 1 0
2 22307 1 0
2 22308 1 0
2 22309 1 0
2 22310 1 0
2 22311 1 0
2 22312 1 0
2 22313 1 0
2 22314 1 0
2 22315 1 0
2 22316 1 0
2 22317 1 0
2 22318 1 0
2 22319 1 0
2 22320 1 0
2 22321 1 0
2 22322 1 0
2 22323 1 0
2 22324 1 0
2 22325 1 0
2 22326 1 0
2 22327 1 0
2 22328 1 0
2 22329 1 0
2 22330 1 0
2 22331 1 0
2 22332 1 0
2 22333 1 0
2 22334 1 0
2 22335 1 0
2 22336 1 0
2 22337 1 0
2 22338 1 0
2 22339 1 0
2 22340 1 0
2 22341 1 0
2 22342 1 0
2 22343 1 0
2 22344 1 0
2 22345 1 0
2 22346 1 0
2 22347 1 0
2 22348 1 0
2 22349 1 0
2 22350 1 0
2 22351 1 0
2 22352 1 0
2 22353 1 0
2 22354 1 0
2 22355 1 0
2 22356 1 0
2 22357 1 0
2 22358 1 0
2 22359 1 0
2 22360 1 0
2 22361 1 0
2 22362 1 0
2 22363 1 0
2 22364 1 0
2 22365 1 0
2 22366 1 0
2 22367 1 0
2 22368 1 0
2 22369 1 0
2 22370 1 0
2 22371 1 0
2 22372 1 0
1 1 0 154 0
2 22373 1 1
2 22374 1 1
2 22375 1 1
2 22376 1 1
2 22377 1 1
2 22378 1 1
2 22379 1 1
2 22380 1 1
2 22381 1 1
2 22382 1 1
2 22383 1 1
2 22384 1 1
2 22385 1 1
2 22386 1 1
2 22387 1 1
2 22388 1 1
2 22389 1 1
2 22390 1 1
2 22391 1 1
2 22392 1 1
2 22393 1 1
2 22394 1 1
2 22395 1 1
2 22396 1 1
2 22397 1 1
2 22398 1 1
2 22399 1 1
2 22400 1 1
2 22401 1 1
2 22402 1 1
2 22403 1 1
2 22404 1 1
2 22405 1 1
2 22406 1 1
2 22407 1 1
2 22408 1 1
2 22409 1 1
2 22410 1 1
2 22411 1 1
2 22412 1 1
2 22413 1 1
2 22414 1 1
2 22415 1 1
2 22416 1 1
2 22417 1 1
2 22418 1 1
2 22419 1 1
2 22420 1 1
2 22421 1 1
2 22422 1 1
2 22423 1 1
2 22424 1 1
2 22425 1 1
2 22426 1 1
2 22427 1 1
2 22428 1 1
2 22429 1 1
2 22430 1 1
2 22431 1 1
2 22432 1 1
2 22433 1 1
2 22434 1 1
2 22435 1 1
2 22436 1 1
2 22437 1 1
2 22438 1 1
2 22439 1 1
2 22440 1 1
2 22441 1 1
2 22442 1 1
2 22443 1 1
2 22444 1 1
2 22445 1 1
2 22446 1 1
2 22447 1 1
2 22448 1 1
2 22449 1 1
2 22450 1 1
2 22451 1 1
2 22452 1 1
2 22453 1 1
2 22454 1 1
2 22455 1 1
2 22456 1 1
2 22457 1 1
2 22458 1 1
2 22459 1 1
2 22460 1 1
2 22461 1 1
2 22462 1 1
2 22463 1 1
2 22464 1 1
2 22465 1 1
2 22466 1 1
2 22467 1 1
2 22468 1 1
2 22469 1 1
2 22470 1 1
2 22471 1 1
2 22472 1 1
2 22473 1 1
2 22474 1 1
2 22475 1 1
2 22476 1 1
2 22477 1 1
2 22478 1 1
2 22479 1 1
2 22480 1 1
2 22481 1 1
2 22482 1 1
2 22483 1 1
2 22484 1 1
2 22485 1 1
2 22486 1 1
2 22487 1 1
2 22488 1 1
2 22489 1 1
2 22490 1 1
2 22491 1 1
2 22492 1 1
2 22493 1 1
2 22494 1 1
2 22495 1 1
2 22496 1 1
2 22497 1 1
2 22498 1 1
2 22499 1 1
2 22500 1 1
2 22501 1 1
2 22502 1 1
2 22503 1 1
2 22504 1 1
2 22505 1 1
2 22506 1 1
2 22507 1 1
2 22508 1 1
2 22509 1 1
2 22510 1 1
2 22511 1 1
2 22512 1 1
2 22513 1 1
2 22514 1 1
2 22515 1 1
2 22516 1 1
2 22517 1 1
2 22518 1 1
2 22519 1 1
2 22520 1 1
2 22521 1 1
2 22522 1 1
2 22523 1 1
2 22524 1 1
2 22525 1 1
2 22526 1 1
1 2 0 136 0
2 22527 1 2
2 22528 1 2
2 22529 1 2
2 22530 1 2
2 22531 1 2
2 22532 1 2
2 22533 1 2
2 22534 1 2
2 22535 1 2
2 22536 1 2
2 22537 1 2
2 22538 1 2
2 22539 1 2
2 22540 1 2
2 22541 1 2
2 22542 1 2
2 22543 1 2
2 22544 1 2
2 22545 1 2
2 22546 1 2
2 22547 1 2
2 22548 1 2
2 22549 1 2
2 22550 1 2
2 22551 1 2
2 22552 1 2
2 22553 1 2
2 22554 1 2
2 22555 1 2
2 22556 1 2
2 22557 1 2
2 22558 1 2
2 22559 1 2
2 22560 1 2
2 22561 1 2
2 22562 1 2
2 22563 1 2
2 22564 1 2
2 22565 1 2
2 22566 1 2
2 22567 1 2
2 22568 1 2
2 22569 1 2
2 22570 1 2
2 22571 1 2
2 22572 1 2
2 22573 1 2
2 22574 1 2
2 22575 1 2
2 22576 1 2
2 22577 1 2
2 22578 1 2
2 22579 1 2
2 22580 1 2
2 22581 1 2
2 22582 1 2
2 22583 1 2
2 22584 1 2
2 22585 1 2
2 22586 1 2
2 22587 1 2
2 22588 1 2
2 22589 1 2
2 22590 1 2
2 22591 1 2
2 22592 1 2
2 22593 1 2
2 22594 1 2
2 22595 1 2
2 22596 1 2
2 22597 1 2
2 22598 1 2
2 22599 1 2
2 22600 1 2
2 22601 1 2
2 22602 1 2
2 22603 1 2
2 22604 1 2
2 22605 1 2
2 22606 1 2
2 22607 1 2
2 22608 1 2
2 22609 1 2
2 22610 1 2
2 22611 1 2
2 22612 1 2
2 22613 1 2
2 22614 1 2
2 22615 1 2
2 22616 1 2
2 22617 1 2
2 22618 1 2
2 22619 1 2
2 22620 1 2
2 22621 1 2
2 22622 1 2
2 22623 1 2
2 22624 1 2
2 22625 1 2
2 22626 1 2
2 22627 1 2
2 22628 1 2
2 22629 1 2
2 22630 1 2
2 22631 1 2
2 22632 1 2
2 22633 1 2
2 22634 1 2
2 22635 1 2
2 22636 1 2
2 22637 1 2
2 22638 1 2
2 22639 1 2
2 22640 1 2
2 22641 1 2
2 22642 1 2
2 22643 1 2
2 22644 1 2
2 22645 1 2
2 22646 1 2
2 22647 1 2
2 22648 1 2
2 22649 1 2
2 22650 1 2
2 22651 1 2
2 22652 1 2
2 22653 1 2
2 22654 1 2
2 22655 1 2
2 22656 1 2
2 22657 1 2
2 22658 1 2
2 22659 1 2
2 22660 1 2
2 22661 1 2
2 22662 1 2
1 3 0 113 0
2 22663 1 3
2 22664 1 3
2 22665 1 3
2 22666 1 3
2 22667 1 3
2 22668 1 3
2 22669 1 3
2 22670 1 3
2 22671 1 3
2 22672 1 3
2 22673 1 3
2 22674 1 3
2 22675 1 3
2 22676 1 3
2 22677 1 3
2 22678 1 3
2 22679 1 3
2 22680 1 3
2 22681 1 3
2 22682 1 3
2 22683 1 3
2 22684 1 3
2 22685 1 3
2 22686 1 3
2 22687 1 3
2 22688 1 3
2 22689 1 3
2 22690 1 3
2 22691 1 3
2 22692 1 3
2 22693 1 3
2 22694 1 3
2 22695 1 3
2 22696 1 3
2 22697 1 3
2 22698 1 3
2 22699 1 3
2 22700 1 3
2 22701 1 3
2 22702 1 3
2 22703 1 3
2 22704 1 3
2 22705 1 3
2 22706 1 3
2 22707 1 3
2 22708 1 3
2 22709 1 3
2 22710 1 3
2 22711 1 3
2 22712 1 3
2 22713 1 3
2 22714 1 3
2 22715 1 3
2 22716 1 3
2 22717 1 3
2 22718 1 3
2 22719 1 3
2 22720 1 3
2 22721 1 3
2 22722 1 3
2 22723 1 3
2 22724 1 3
2 22725 1 3
2 22726 1 3
2 22727 1 3
2 22728 1 3
2 22729 1 3
2 22730 1 3
2 22731 1 3
2 22732 1 3
2 22733 1 3
2 22734 1 3
2 22735 1 3
2 22736 1 3
2 22737 1 3
2 22738 1 3
2 22739 1 3
2 22740 1 3
2 22741 1 3
2 22742 1 3
2 22743 1 3
2 22744 1 3
2 22745 1 3
2 22746 1 3
2 22747 1 3
2 22748 1 3
2 22749 1 3
2 22750 1 3
2 22751 1 3
2 22752 1 3
2 22753 1 3
2 22754 1 3
2 22755 1 3
2 22756 1 3
2 22757 1 3
2 22758 1 3
2 22759 1 3
2 22760 1 3
2 22761 1 3
2 22762 1 3
2 22763 1 3
2 22764 1 3
2 22765 1 3
2 22766 1 3
2 22767 1 3
2 22768 1 3
2 22769 1 3
2 22770 1 3
2 22771 1 3
2 22772 1 3
2 22773 1 3
2 22774 1 3
2 22775 1 3
1 4 0 96 0
2 22776 1 4
2 22777 1 4
2 22778 1 4
2 22779 1 4
2 22780 1 4
2 22781 1 4
2 22782 1 4
2 22783 1 4
2 22784 1 4
2 22785 1 4
2 22786 1 4
2 22787 1 4
2 22788 1 4
2 22789 1 4
2 22790 1 4
2 22791 1 4
2 22792 1 4
2 22793 1 4
2 22794 1 4
2 22795 1 4
2 22796 1 4
2 22797 1 4
2 22798 1 4
2 22799 1 4
2 22800 1 4
2 22801 1 4
2 22802 1 4
2 22803 1 4
2 22804 1 4
2 22805 1 4
2 22806 1 4
2 22807 1 4
2 22808 1 4
2 22809 1 4
2 22810 1 4
2 22811 1 4
2 22812 1 4
2 22813 1 4
2 22814 1 4
2 22815 1 4
2 22816 1 4
2 22817 1 4
2 22818 1 4
2 22819 1 4
2 22820 1 4
2 22821 1 4
2 22822 1 4
2 22823 1 4
2 22824 1 4
2 22825 1 4
2 22826 1 4
2 22827 1 4
2 22828 1 4
2 22829 1 4
2 22830 1 4
2 22831 1 4
2 22832 1 4
2 22833 1 4
2 22834 1 4
2 22835 1 4
2 22836 1 4
2 22837 1 4
2 22838 1 4
2 22839 1 4
2 22840 1 4
2 22841 1 4
2 22842 1 4
2 22843 1 4
2 22844 1 4
2 22845 1 4
2 22846 1 4
2 22847 1 4
2 22848 1 4
2 22849 1 4
2 22850 1 4
2 22851 1 4
2 22852 1 4
2 22853 1 4
2 22854 1 4
2 22855 1 4
2 22856 1 4
2 22857 1 4
2 22858 1 4
2 22859 1 4
2 22860 1 4
2 22861 1 4
2 22862 1 4
2 22863 1 4
2 22864 1 4
2 22865 1 4
2 22866 1 4
2 22867 1 4
2 22868 1 4
2 22869 1 4
2 22870 1 4
2 22871 1 4
1 5 0 118 0
2 22872 1 5
2 22873 1 5
2 22874 1 5
2 22875 1 5
2 22876 1 5
2 22877 1 5
2 22878 1 5
2 22879 1 5
2 22880 1 5
2 22881 1 5
2 22882 1 5
2 22883 1 5
2 22884 1 5
2 22885 1 5
2 22886 1 5
2 22887 1 5
2 22888 1 5
2 22889 1 5
2 22890 1 5
2 22891 1 5
2 22892 1 5
2 22893 1 5
2 22894 1 5
2 22895 1 5
2 22896 1 5
2 22897 1 5
2 22898 1 5
2 22899 1 5
2 22900 1 5
2 22901 1 5
2 22902 1 5
2 22903 1 5
2 22904 1 5
2 22905 1 5
2 22906 1 5
2 22907 1 5
2 22908 1 5
2 22909 1 5
2 22910 1 5
2 22911 1 5
2 22912 1 5
2 22913 1 5
2 22914 1 5
2 22915 1 5
2 22916 1 5
2 22917 1 5
2 22918 1 5
2 22919 1 5
2 22920 1 5
2 22921 1 5
2 22922 1 5
2 22923 1 5
2 22924 1 5
2 22925 1 5
2 22926 1 5
2 22927 1 5
2 22928 1 5
2 22929 1 5
2 22930 1 5
2 22931 1 5
2 22932 1 5
2 22933 1 5
2 22934 1 5
2 22935 1 5
2 22936 1 5
2 22937 1 5
2 22938 1 5
2 22939 1 5
2 22940 1 5
2 22941 1 5
2 22942 1 5
2 22943 1 5
2 22944 1 5
2 22945 1 5
2 22946 1 5
2 22947 1 5
2 22948 1 5
2 22949 1 5
2 22950 1 5
2 22951 1 5
2 22952 1 5
2 22953 1 5
2 22954 1 5
2 22955 1 5
2 22956 1 5
2 22957 1 5
2 22958 1 5
2 22959 1 5
2 22960 1 5
2 22961 1 5
2 22962 1 5
2 22963 1 5
2 22964 1 5
2 22965 1 5
2 22966 1 5
2 22967 1 5
2 22968 1 5
2 22969 1 5
2 22970 1 5
2 22971 1 5
2 22972 1 5
2 22973 1 5
2 22974 1 5
2 22975 1 5
2 22976 1 5
2 22977 1 5
2 22978 1 5
2 22979 1 5
2 22980 1 5
2 22981 1 5
2 22982 1 5
2 22983 1 5
2 22984 1 5
2 22985 1 5
2 22986 1 5
2 22987 1 5
2 22988 1 5
2 22989 1 5
1 6 0 66 0
2 22990 1 6
2 22991 1 6
2 22992 1 6
2 22993 1 6
2 22994 1 6
2 22995 1 6
2 22996 1 6
2 22997 1 6
2 22998 1 6
2 22999 1 6
2 23000 1 6
2 23001 1 6
2 23002 1 6
2 23003 1 6
2 23004 1 6
2 23005 1 6
2 23006 1 6
2 23007 1 6
2 23008 1 6
2 23009 1 6
2 23010 1 6
2 23011 1 6
2 23012 1 6
2 23013 1 6
2 23014 1 6
2 23015 1 6
2 23016 1 6
2 23017 1 6
2 23018 1 6
2 23019 1 6
2 23020 1 6
2 23021 1 6
2 23022 1 6
2 23023 1 6
2 23024 1 6
2 23025 1 6
2 23026 1 6
2 23027 1 6
2 23028 1 6
2 23029 1 6
2 23030 1 6
2 23031 1 6
2 23032 1 6
2 23033 1 6
2 23034 1 6
2 23035 1 6
2 23036 1 6
2 23037 1 6
2 23038 1 6
2 23039 1 6
2 23040 1 6
2 23041 1 6
2 23042 1 6
2 23043 1 6
2 23044 1 6
2 23045 1 6
2 23046 1 6
2 23047 1 6
2 23048 1 6
2 23049 1 6
2 23050 1 6
2 23051 1 6
2 23052 1 6
2 23053 1 6
2 23054 1 6
2 23055 1 6
1 7 0 101 0
2 23056 1 7
2 23057 1 7
2 23058 1 7
2 23059 1 7
2 23060 1 7
2 23061 1 7
2 23062 1 7
2 23063 1 7
2 23064 1 7
2 23065 1 7
2 23066 1 7
2 23067 1 7
2 23068 1 7
2 23069 1 7
2 23070 1 7
2 23071 1 7
2 23072 1 7
2 23073 1 7
2 23074 1 7
2 23075 1 7
2 23076 1 7
2 23077 1 7
2 23078 1 7
2 23079 1 7
2 23080 1 7
2 23081 1 7
2 23082 1 7
2 23083 1 7
2 23084 1 7
2 23085 1 7
2 23086 1 7
2 23087 1 7
2 23088 1 7
2 23089 1 7
2 23090 1 7
2 23091 1 7
2 23092 1 7
2 23093 1 7
2 23094 1 7
2 23095 1 7
2 23096 1 7
2 23097 1 7
2 23098 1 7
2 23099 1 7
2 23100 1 7
2 23101 1 7
2 23102 1 7
2 23103 1 7
2 23104 1 7
2 23105 1 7
2 23106 1 7
2 23107 1 7
2 23108 1 7
2 23109 1 7
2 23110 1 7
2 23111 1 7
2 23112 1 7
2 23113 1 7
2 23114 1 7
2 23115 1 7
2 23116 1 7
2 23117 1 7
2 23118 1 7
2 23119 1 7
2 23120 1 7
2 23121 1 7
2 23122 1 7
2 23123 1 7
2 23124 1 7
2 23125 1 7
2 23126 1 7
2 23127 1 7
2 23128 1 7
2 23129 1 7
2 23130 1 7
2 23131 1 7
2 23132 1 7
2 23133 1 7
2 23134 1 7
2 23135 1 7
2 23136 1 7
2 23137 1 7
2 23138 1 7
2 23139 1 7
2 23140 1 7
2 23141 1 7
2 23142 1 7
2 23143 1 7
2 23144 1 7
2 23145 1 7
2 23146 1 7
2 23147 1 7
2 23148 1 7
2 23149 1 7
2 23150 1 7
2 23151 1 7
2 23152 1 7
2 23153 1 7
2 23154 1 7
2 23155 1 7
2 23156 1 7
1 8 0 50 0
2 23157 1 8
2 23158 1 8
2 23159 1 8
2 23160 1 8
2 23161 1 8
2 23162 1 8
2 23163 1 8
2 23164 1 8
2 23165 1 8
2 23166 1 8
2 23167 1 8
2 23168 1 8
2 23169 1 8
2 23170 1 8
2 23171 1 8
2 23172 1 8
2 23173 1 8
2 23174 1 8
2 23175 1 8
2 23176 1 8
2 23177 1 8
2 23178 1 8
2 23179 1 8
2 23180 1 8
2 23181 1 8
2 23182 1 8
2 23183 1 8
2 23184 1 8
2 23185 1 8
2 23186 1 8
2 23187 1 8
2 23188 1 8
2 23189 1 8
2 23190 1 8
2 23191 1 8
2 23192 1 8
2 23193 1 8
2 23194 1 8
2 23195 1 8
2 23196 1 8
2 23197 1 8
2 23198 1 8
2 23199 1 8
2 23200 1 8
2 23201 1 8
2 23202 1 8
2 23203 1 8
2 23204 1 8
2 23205 1 8
2 23206 1 8
1 9 0 82 0
2 23207 1 9
2 23208 1 9
2 23209 1 9
2 23210 1 9
2 23211 1 9
2 23212 1 9
2 23213 1 9
2 23214 1 9
2 23215 1 9
2 23216 1 9
2 23217 1 9
2 23218 1 9
2 23219 1 9
2 23220 1 9
2 23221 1 9
2 23222 1 9
2 23223 1 9
2 23224 1 9
2 23225 1 9
2 23226 1 9
2 23227 1 9
2 23228 1 9
2 23229 1 9
2 23230 1 9
2 23231 1 9
2 23232 1 9
2 23233 1 9
2 23234 1 9
2 23235 1 9
2 23236 1 9
2 23237 1 9
2 23238 1 9
2 23239 1 9
2 23240 1 9
2 23241 1 9
2 23242 1 9
2 23243 1 9
2 23244 1 9
2 23245 1 9
2 23246 1 9
2 23247 1 9
2 23248 1 9
2 23249 1 9
2 23250 1 9
2 23251 1 9
2 23252 1 9
2 23253 1 9
2 23254 1 9
2 23255 1 9
2 23256 1 9
2 23257 1 9
2 23258 1 9
2 23259 1 9
2 23260 1 9
2 23261 1 9
2 23262 1 9
2 23263 1 9
2 23264 1 9
2 23265 1 9
2 23266 1 9
2 23267 1 9
2 23268 1 9
2 23269 1 9
2 23270 1 9
2 23271 1 9
2 23272 1 9
2 23273 1 9
2 23274 1 9
2 23275 1 9
2 23276 1 9
2 23277 1 9
2 23278 1 9
2 23279 1 9
2 23280 1 9
2 23281 1 9
2 23282 1 9
2 23283 1 9
2 23284 1 9
2 23285 1 9
2 23286 1 9
2 23287 1 9
2 23288 1 9
1 10 0 79 0
2 23289 1 10
2 23290 1 10
2 23291 1 10
2 23292 1 10
2 23293 1 10
2 23294 1 10
2 23295 1 10
2 23296 1 10
2 23297 1 10
2 23298 1 10
2 23299 1 10
2 23300 1 10
2 23301 1 10
2 23302 1 10
2 23303 1 10
2 23304 1 10
2 23305 1 10
2 23306 1 10
2 23307 1 10
2 23308 1 10
2 23309 1 10
2 23310 1 10
2 23311 1 10
2 23312 1 10
2 23313 1 10
2 23314 1 10
2 23315 1 10
2 23316 1 10
2 23317 1 10
2 23318 1 10
2 23319 1 10
2 23320 1 10
2 23321 1 10
2 23322 1 10
2 23323 1 10
2 23324 1 10
2 23325 1 10
2 23326 1 10
2 23327 1 10
2 23328 1 10
2 23329 1 10
2 23330 1 10
2 23331 1 10
2 23332 1 10
2 23333 1 10
2 23334 1 10
2 23335 1 10
2 23336 1 10
2 23337 1 10
2 23338 1 10
2 23339 1 10
2 23340 1 10
2 23341 1 10
2 23342 1 10
2 23343 1 10
2 23344 1 10
2 23345 1 10
2 23346 1 10
2 23347 1 10
2 23348 1 10
2 23349 1 10
2 23350 1 10
2 23351 1 10
2 23352 1 10
2 23353 1 10
2 23354 1 10
2 23355 1 10
2 23356 1 10
2 23357 1 10
2 23358 1 10
2 23359 1 10
2 23360 1 10
2 23361 1 10
2 23362 1 10
2 23363 1 10
2 23364 1 10
2 23365 1 10
2 23366 1 10
2 23367 1 10
1 11 0 70 0
2 23368 1 11
2 23369 1 11
2 23370 1 11
2 23371 1 11
2 23372 1 11
2 23373 1 11
2 23374 1 11
2 23375 1 11
2 23376 1 11
2 23377 1 11
2 23378 1 11
2 23379 1 11
2 23380 1 11
2 23381 1 11
2 23382 1 11
2 23383 1 11
2 23384 1 11
2 23385 1 11
2 23386 1 11
2 23387 1 11
2 23388 1 11
2 23389 1 11
2 23390 1 11
2 23391 1 11
2 23392 1 11
2 23393 1 11
2 23394 1 11
2 23395 1 11
2 23396 1 11
2 23397 1 11
2 23398 1 11
2 23399 1 11
2 23400 1 11
2 23401 1 11
2 23402 1 11
2 23403 1 11
2 23404 1 11
2 23405 1 11
2 23406 1 11
2 23407 1 11
2 23408 1 11
2 23409 1 11
2 23410 1 11
2 23411 1 11
2 23412 1 11
2 23413 1 11
2 23414 1 11
2 23415 1 11
2 23416 1 11
2 23417 1 11
2 23418 1 11
2 23419 1 11
2 23420 1 11
2 23421 1 11
2 23422 1 11
2 23423 1 11
2 23424 1 11
2 23425 1 11
2 23426 1 11
2 23427 1 11
2 23428 1 11
2 23429 1 11
2 23430 1 11
2 23431 1 11
2 23432 1 11
2 23433 1 11
2 23434 1 11
2 23435 1 11
2 23436 1 11
2 23437 1 11
1 12 0 52 0
2 23438 1 12
2 23439 1 12
2 23440 1 12
2 23441 1 12
2 23442 1 12
2 23443 1 12
2 23444 1 12
2 23445 1 12
2 23446 1 12
2 23447 1 12
2 23448 1 12
2 23449 1 12
2 23450 1 12
2 23451 1 12
2 23452 1 12
2 23453 1 12
2 23454 1 12
2 23455 1 12
2 23456 1 12
2 23457 1 12
2 23458 1 12
2 23459 1 12
2 23460 1 12
2 23461 1 12
2 23462 1 12
2 23463 1 12
2 23464 1 12
2 23465 1 12
2 23466 1 12
2 23467 1 12
2 23468 1 12
2 23469 1 12
2 23470 1 12
2 23471 1 12
2 23472 1 12
2 23473 1 12
2 23474 1 12
2 23475 1 12
2 23476 1 12
2 23477 1 12
2 23478 1 12
2 23479 1 12
2 23480 1 12
2 23481 1 12
2 23482 1 12
2 23483 1 12
2 23484 1 12
2 23485 1 12
2 23486 1 12
2 23487 1 12
2 23488 1 12
2 23489 1 12
1 13 0 77 0
2 23490 1 13
2 23491 1 13
2 23492 1 13
2 23493 1 13
2 23494 1 13
2 23495 1 13
2 23496 1 13
2 23497 1 13
2 23498 1 13
2 23499 1 13
2 23500 1 13
2 23501 1 13
2 23502 1 13
2 23503 1 13
2 23504 1 13
2 23505 1 13
2 23506 1 13
2 23507 1 13
2 23508 1 13
2 23509 1 13
2 23510 1 13
2 23511 1 13
2 23512 1 13
2 23513 1 13
2 23514 1 13
2 23515 1 13
2 23516 1 13
2 23517 1 13
2 23518 1 13
2 23519 1 13
2 23520 1 13
2 23521 1 13
2 23522 1 13
2 23523 1 13
2 23524 1 13
2 23525 1 13
2 23526 1 13
2 23527 1 13
2 23528 1 13
2 23529 1 13
2 23530 1 13
2 23531 1 13
2 23532 1 13
2 23533 1 13
2 23534 1 13
2 23535 1 13
2 23536 1 13
2 23537 1 13
2 23538 1 13
2 23539 1 13
2 23540 1 13
2 23541 1 13
2 23542 1 13
2 23543 1 13
2 23544 1 13
2 23545 1 13
2 23546 1 13
2 23547 1 13
2 23548 1 13
2 23549 1 13
2 23550 1 13
2 23551 1 13
2 23552 1 13
2 23553 1 13
2 23554 1 13
2 23555 1 13
2 23556 1 13
2 23557 1 13
2 23558 1 13
2 23559 1 13
2 23560 1 13
2 23561 1 13
2 23562 1 13
2 23563 1 13
2 23564 1 13
2 23565 1 13
2 23566 1 13
1 14 0 29 0
2 23567 1 14
2 23568 1 14
2 23569 1 14
2 23570 1 14
2 23571 1 14
2 23572 1 14
2 23573 1 14
2 23574 1 14
2 23575 1 14
2 23576 1 14
2 23577 1 14
2 23578 1 14
2 23579 1 14
2 23580 1 14
2 23581 1 14
2 23582 1 14
2 23583 1 14
2 23584 1 14
2 23585 1 14
2 23586 1 14
2 23587 1 14
2 23588 1 14
2 23589 1 14
2 23590 1 14
2 23591 1 14
2 23592 1 14
2 23593 1 14
2 23594 1 14
2 23595 1 14
1 15 0 49 0
2 23596 1 15
2 23597 1 15
2 23598 1 15
2 23599 1 15
2 23600 1 15
2 23601 1 15
2 23602 1 15
2 23603 1 15
2 23604 1 15
2 23605 1 15
2 23606 1 15
2 23607 1 15
2 23608 1 15
2 23609 1 15
2 23610 1 15
2 23611 1 15
2 23612 1 15
2 23613 1 15
2 23614 1 15
2 23615 1 15
2 23616 1 15
2 23617 1 15
2 23618 1 15
2 23619 1 15
2 23620 1 15
2 23621 1 15
2 23622 1 15
2 23623 1 15
2 23624 1 15
2 23625 1 15
2 23626 1 15
2 23627 1 15
2 23628 1 15
2 23629 1 15
2 23630 1 15
2 23631 1 15
2 23632 1 15
2 23633 1 15
2 23634 1 15
2 23635 1 15
2 23636 1 15
2 23637 1 15
2 23638 1 15
2 23639 1 15
2 23640 1 15
2 23641 1 15
2 23642 1 15
2 23643 1 15
2 23644 1 15
1 16 0 2 0
2 23645 1 16
2 23646 1 16
1 17 0 103 0
2 23647 1 17
2 23648 1 17
2 23649 1 17
2 23650 1 17
2 23651 1 17
2 23652 1 17
2 23653 1 17
2 23654 1 17
2 23655 1 17
2 23656 1 17
2 23657 1 17
2 23658 1 17
2 23659 1 17
2 23660 1 17
2 23661 1 17
2 23662 1 17
2 23663 1 17
2 23664 1 17
2 23665 1 17
2 23666 1 17
2 23667 1 17
2 23668 1 17
2 23669 1 17
2 23670 1 17
2 23671 1 17
2 23672 1 17
2 23673 1 17
2 23674 1 17
2 23675 1 17
2 23676 1 17
2 23677 1 17
2 23678 1 17
2 23679 1 17
2 23680 1 17
2 23681 1 17
2 23682 1 17
2 23683 1 17
2 23684 1 17
2 23685 1 17
2 23686 1 17
2 23687 1 17
2 23688 1 17
2 23689 1 17
2 23690 1 17
2 23691 1 17
2 23692 1 17
2 23693 1 17
2 23694 1 17
2 23695 1 17
2 23696 1 17
2 23697 1 17
2 23698 1 17
2 23699 1 17
2 23700 1 17
2 23701 1 17
2 23702 1 17
2 23703 1 17
2 23704 1 17
2 23705 1 17
2 23706 1 17
2 23707 1 17
2 23708 1 17
2 23709 1 17
2 23710 1 17
2 23711 1 17
2 23712 1 17
2 23713 1 17
2 23714 1 17
2 23715 1 17
2 23716 1 17
2 23717 1 17
2 23718 1 17
2 23719 1 17
2 23720 1 17
2 23721 1 17
2 23722 1 17
2 23723 1 17
2 23724 1 17
2 23725 1 17
2 23726 1 17
2 23727 1 17
2 23728 1 17
2 23729 1 17
2 23730 1 17
2 23731 1 17
2 23732 1 17
2 23733 1 17
2 23734 1 17
2 23735 1 17
2 23736 1 17
2 23737 1 17
2 23738 1 17
2 23739 1 17
2 23740 1 17
2 23741 1 17
2 23742 1 17
2 23743 1 17
2 23744 1 17
2 23745 1 17
2 23746 1 17
2 23747 1 17
2 23748 1 17
2 23749 1 17
1 18 0 110 0
2 23750 1 18
2 23751 1 18
2 23752 1 18
2 23753 1 18
2 23754 1 18
2 23755 1 18
2 23756 1 18
2 23757 1 18
2 23758 1 18
2 23759 1 18
2 23760 1 18
2 23761 1 18
2 23762 1 18
2 23763 1 18
2 23764 1 18
2 23765 1 18
2 23766 1 18
2 23767 1 18
2 23768 1 18
2 23769 1 18
2 23770 1 18
2 23771 1 18
2 23772 1 18
2 23773 1 18
2 23774 1 18
2 23775 1 18
2 23776 1 18
2 23777 1 18
2 23778 1 18
2 23779 1 18
2 23780 1 18
2 23781 1 18
2 23782 1 18
2 23783 1 18
2 23784 1 18
2 23785 1 18
2 23786 1 18
2 23787 1 18
2 23788 1 18
2 23789 1 18
2 23790 1 18
2 23791 1 18
2 23792 1 18
2 23793 1 18
2 23794 1 18
2 23795 1 18
2 23796 1 18
2 23797 1 18
2 23798 1 18
2 23799 1 18
2 23800 1 18
2 23801 1 18
2 23802 1 18
2 23803 1 18
2 23804 1 18
2 23805 1 18
2 23806 1 18
2 23807 1 18
2 23808 1 18
2 23809 1 18
2 23810 1 18
2 23811 1 18
2 23812 1 18
2 23813 1 18
2 23814 1 18
2 23815 1 18
2 23816 1 18
2 23817 1 18
2 23818 1 18
2 23819 1 18
2 23820 1 18
2 23821 1 18
2 23822 1 18
2 23823 1 18
2 23824 1 18
2 23825 1 18
2 23826 1 18
2 23827 1 18
2 23828 1 18
2 23829 1 18
2 23830 1 18
2 23831 1 18
2 23832 1 18
2 23833 1 18
2 23834 1 18
2 23835 1 18
2 23836 1 18
2 23837 1 18
2 23838 1 18
2 23839 1 18
2 23840 1 18
2 23841 1 18
2 23842 1 18
2 23843 1 18
2 23844 1 18
2 23845 1 18
2 23846 1 18
2 23847 1 18
2 23848 1 18
2 23849 1 18
2 23850 1 18
2 23851 1 18
2 23852 1 18
2 23853 1 18
2 23854 1 18
2 23855 1 18
2 23856 1 18
2 23857 1 18
2 23858 1 18
2 23859 1 18
1 19 0 102 0
2 23860 1 19
2 23861 1 19
2 23862 1 19
2 23863 1 19
2 23864 1 19
2 23865 1 19
2 23866 1 19
2 23867 1 19
2 23868 1 19
2 23869 1 19
2 23870 1 19
2 23871 1 19
2 23872 1 19
2 23873 1 19
2 23874 1 19
2 23875 1 19
2 23876 1 19
2 23877 1 19
2 23878 1 19
2 23879 1 19
2 23880 1 19
2 23881 1 19
2 23882 1 19
2 23883 1 19
2 23884 1 19
2 23885 1 19
2 23886 1 19
2 23887 1 19
2 23888 1 19
2 23889 1 19
2 23890 1 19
2 23891 1 19
2 23892 1 19
2 23893 1 19
2 23894 1 19
2 23895 1 19
2 23896 1 19
2 23897 1 19
2 23898 1 19
2 23899 1 19
2 23900 1 19
2 23901 1 19
2 23902 1 19
2 23903 1 19
2 23904 1 19
2 23905 1 19
2 23906 1 19
2 23907 1 19
2 23908 1 19
2 23909 1 19
2 23910 1 19
2 23911 1 19
2 23912 1 19
2 23913 1 19
2 23914 1 19
2 23915 1 19
2 23916 1 19
2 23917 1 19
2 23918 1 19
2 23919 1 19
2 23920 1 19
2 23921 1 19
2 23922 1 19
2 23923 1 19
2 23924 1 19
2 23925 1 19
2 23926 1 19
2 23927 1 19
2 23928 1 19
2 23929 1 19
2 23930 1 19
2 23931 1 19
2 23932 1 19
2 23933 1 19
2 23934 1 19
2 23935 1 19
2 23936 1 19
2 23937 1 19
2 23938 1 19
2 23939 1 19
2 23940 1 19
2 23941 1 19
2 23942 1 19
2 23943 1 19
2 23944 1 19
2 23945 1 19
2 23946 1 19
2 23947 1 19
2 23948 1 19
2 23949 1 19
2 23950 1 19
2 23951 1 19
2 23952 1 19
2 23953 1 19
2 23954 1 19
2 23955 1 19
2 23956 1 19
2 23957 1 19
2 23958 1 19
2 23959 1 19
2 23960 1 19
2 23961 1 19
1 20 0 86 0
2 23962 1 20
2 23963 1 20
2 23964 1 20
2 23965 1 20
2 23966 1 20
2 23967 1 20
2 23968 1 20
2 23969 1 20
2 23970 1 20
2 23971 1 20
2 23972 1 20
2 23973 1 20
2 23974 1 20
2 23975 1 20
2 23976 1 20
2 23977 1 20
2 23978 1 20
2 23979 1 20
2 23980 1 20
2 23981 1 20
2 23982 1 20
2 23983 1 20
2 23984 1 20
2 23985 1 20
2 23986 1 20
2 23987 1 20
2 23988 1 20
2 23989 1 20
2 23990 1 20
2 23991 1 20
2 23992 1 20
2 23993 1 20
2 23994 1 20
2 23995 1 20
2 23996 1 20
2 23997 1 20
2 23998 1 20
2 23999 1 20
2 24000 1 20
2 24001 1 20
2 24002 1 20
2 24003 1 20
2 24004 1 20
2 24005 1 20
2 24006 1 20
2 24007 1 20
2 24008 1 20
2 24009 1 20
2 24010 1 20
2 24011 1 20
2 24012 1 20
2 24013 1 20
2 24014 1 20
2 24015 1 20
2 24016 1 20
2 24017 1 20
2 24018 1 20
2 24019 1 20
2 24020 1 20
2 24021 1 20
2 24022 1 20
2 24023 1 20
2 24024 1 20
2 24025 1 20
2 24026 1 20
2 24027 1 20
2 24028 1 20
2 24029 1 20
2 24030 1 20
2 24031 1 20
2 24032 1 20
2 24033 1 20
2 24034 1 20
2 24035 1 20
2 24036 1 20
2 24037 1 20
2 24038 1 20
2 24039 1 20
2 24040 1 20
2 24041 1 20
2 24042 1 20
2 24043 1 20
2 24044 1 20
2 24045 1 20
2 24046 1 20
2 24047 1 20
1 21 0 92 0
2 24048 1 21
2 24049 1 21
2 24050 1 21
2 24051 1 21
2 24052 1 21
2 24053 1 21
2 24054 1 21
2 24055 1 21
2 24056 1 21
2 24057 1 21
2 24058 1 21
2 24059 1 21
2 24060 1 21
2 24061 1 21
2 24062 1 21
2 24063 1 21
2 24064 1 21
2 24065 1 21
2 24066 1 21
2 24067 1 21
2 24068 1 21
2 24069 1 21
2 24070 1 21
2 24071 1 21
2 24072 1 21
2 24073 1 21
2 24074 1 21
2 24075 1 21
2 24076 1 21
2 24077 1 21
2 24078 1 21
2 24079 1 21
2 24080 1 21
2 24081 1 21
2 24082 1 21
2 24083 1 21
2 24084 1 21
2 24085 1 21
2 24086 1 21
2 24087 1 21
2 24088 1 21
2 24089 1 21
2 24090 1 21
2 24091 1 21
2 24092 1 21
2 24093 1 21
2 24094 1 21
2 24095 1 21
2 24096 1 21
2 24097 1 21
2 24098 1 21
2 24099 1 21
2 24100 1 21
2 24101 1 21
2 24102 1 21
2 24103 1 21
2 24104 1 21
2 24105 1 21
2 24106 1 21
2 24107 1 21
2 24108 1 21
2 24109 1 21
2 24110 1 21
2 24111 1 21
2 24112 1 21
2 24113 1 21
2 24114 1 21
2 24115 1 21
2 24116 1 21
2 24117 1 21
2 24118 1 21
2 24119 1 21
2 24120 1 21
2 24121 1 21
2 24122 1 21
2 24123 1 21
2 24124 1 21
2 24125 1 21
2 24126 1 21
2 24127 1 21
2 24128 1 21
2 24129 1 21
2 24130 1 21
2 24131 1 21
2 24132 1 21
2 24133 1 21
2 24134 1 21
2 24135 1 21
2 24136 1 21
2 24137 1 21
2 24138 1 21
2 24139 1 21
1 22 0 81 0
2 24140 1 22
2 24141 1 22
2 24142 1 22
2 24143 1 22
2 24144 1 22
2 24145 1 22
2 24146 1 22
2 24147 1 22
2 24148 1 22
2 24149 1 22
2 24150 1 22
2 24151 1 22
2 24152 1 22
2 24153 1 22
2 24154 1 22
2 24155 1 22
2 24156 1 22
2 24157 1 22
2 24158 1 22
2 24159 1 22
2 24160 1 22
2 24161 1 22
2 24162 1 22
2 24163 1 22
2 24164 1 22
2 24165 1 22
2 24166 1 22
2 24167 1 22
2 24168 1 22
2 24169 1 22
2 24170 1 22
2 24171 1 22
2 24172 1 22
2 24173 1 22
2 24174 1 22
2 24175 1 22
2 24176 1 22
2 24177 1 22
2 24178 1 22
2 24179 1 22
2 24180 1 22
2 24181 1 22
2 24182 1 22
2 24183 1 22
2 24184 1 22
2 24185 1 22
2 24186 1 22
2 24187 1 22
2 24188 1 22
2 24189 1 22
2 24190 1 22
2 24191 1 22
2 24192 1 22
2 24193 1 22
2 24194 1 22
2 24195 1 22
2 24196 1 22
2 24197 1 22
2 24198 1 22
2 24199 1 22
2 24200 1 22
2 24201 1 22
2 24202 1 22
2 24203 1 22
2 24204 1 22
2 24205 1 22
2 24206 1 22
2 24207 1 22
2 24208 1 22
2 24209 1 22
2 24210 1 22
2 24211 1 22
2 24212 1 22
2 24213 1 22
2 24214 1 22
2 24215 1 22
2 24216 1 22
2 24217 1 22
2 24218 1 22
2 24219 1 22
2 24220 1 22
1 23 0 88 0
2 24221 1 23
2 24222 1 23
2 24223 1 23
2 24224 1 23
2 24225 1 23
2 24226 1 23
2 24227 1 23
2 24228 1 23
2 24229 1 23
2 24230 1 23
2 24231 1 23
2 24232 1 23
2 24233 1 23
2 24234 1 23
2 24235 1 23
2 24236 1 23
2 24237 1 23
2 24238 1 23
2 24239 1 23
2 24240 1 23
2 24241 1 23
2 24242 1 23
2 24243 1 23
2 24244 1 23
2 24245 1 23
2 24246 1 23
2 24247 1 23
2 24248 1 23
2 24249 1 23
2 24250 1 23
2 24251 1 23
2 24252 1 23
2 24253 1 23
2 24254 1 23
2 24255 1 23
2 24256 1 23
2 24257 1 23
2 24258 1 23
2 24259 1 23
2 24260 1 23
2 24261 1 23
2 24262 1 23
2 24263 1 23
2 24264 1 23
2 24265 1 23
2 24266 1 23
2 24267 1 23
2 24268 1 23
2 24269 1 23
2 24270 1 23
2 24271 1 23
2 24272 1 23
2 24273 1 23
2 24274 1 23
2 24275 1 23
2 24276 1 23
2 24277 1 23
2 24278 1 23
2 24279 1 23
2 24280 1 23
2 24281 1 23
2 24282 1 23
2 24283 1 23
2 24284 1 23
2 24285 1 23
2 24286 1 23
2 24287 1 23
2 24288 1 23
2 24289 1 23
2 24290 1 23
2 24291 1 23
2 24292 1 23
2 24293 1 23
2 24294 1 23
2 24295 1 23
2 24296 1 23
2 24297 1 23
2 24298 1 23
2 24299 1 23
2 24300 1 23
2 24301 1 23
2 24302 1 23
2 24303 1 23
2 24304 1 23
2 24305 1 23
2 24306 1 23
2 24307 1 23
2 24308 1 23
1 24 0 31 0
2 24309 1 24
2 24310 1 24
2 24311 1 24
2 24312 1 24
2 24313 1 24
2 24314 1 24
2 24315 1 24
2 24316 1 24
2 24317 1 24
2 24318 1 24
2 24319 1 24
2 24320 1 24
2 24321 1 24
2 24322 1 24
2 24323 1 24
2 24324 1 24
2 24325 1 24
2 24326 1 24
2 24327 1 24
2 24328 1 24
2 24329 1 24
2 24330 1 24
2 24331 1 24
2 24332 1 24
2 24333 1 24
2 24334 1 24
2 24335 1 24
2 24336 1 24
2 24337 1 24
2 24338 1 24
2 24339 1 24
2 24340 1 27
2 24341 1 27
2 24342 1 27
2 24343 1 27
2 24344 1 27
2 24345 1 27
2 24346 1 27
2 24347 1 27
2 24348 1 27
2 24349 1 27
2 24350 1 27
2 24351 1 27
2 24352 1 27
2 24353 1 27
2 24354 1 27
2 24355 1 27
2 24356 1 27
2 24357 1 27
2 24358 1 27
2 24359 1 27
2 24360 1 27
2 24361 1 27
2 24362 1 27
2 24363 1 27
2 24364 1 27
2 24365 1 27
2 24366 1 27
2 24367 1 27
2 24368 1 27
2 24369 1 27
2 24370 1 27
2 24371 1 27
2 24372 1 27
2 24373 1 27
2 24374 1 27
2 24375 1 27
2 24376 1 27
2 24377 1 27
2 24378 1 27
2 24379 1 27
2 24380 1 27
2 24381 1 27
2 24382 1 27
2 24383 1 27
2 24384 1 27
2 24385 1 27
2 24386 1 27
2 24387 1 27
2 24388 1 27
2 24389 1 27
2 24390 1 27
2 24391 1 28
2 24392 1 28
2 24393 1 28
2 24394 1 28
2 24395 1 28
2 24396 1 28
2 24397 1 28
2 24398 1 28
2 24399 1 28
2 24400 1 28
2 24401 1 28
2 24402 1 28
2 24403 1 28
2 24404 1 28
2 24405 1 28
2 24406 1 28
2 24407 1 28
2 24408 1 28
2 24409 1 28
2 24410 1 28
2 24411 1 28
2 24412 1 28
2 24413 1 28
2 24414 1 28
2 24415 1 28
2 24416 1 28
2 24417 1 28
2 24418 1 28
2 24419 1 28
2 24420 1 28
2 24421 1 28
2 24422 1 28
2 24423 1 28
2 24424 1 28
2 24425 1 28
2 24426 1 28
2 24427 1 28
2 24428 1 28
2 24429 1 28
2 24430 1 28
2 24431 1 28
2 24432 1 28
2 24433 1 28
2 24434 1 28
2 24435 1 28
2 24436 1 28
2 24437 1 28
2 24438 1 28
2 24439 1 28
2 24440 1 28
2 24441 1 28
2 24442 1 28
2 24443 1 28
2 24444 1 28
2 24445 1 28
2 24446 1 28
2 24447 1 28
2 24448 1 28
2 24449 1 28
2 24450 1 28
2 24451 1 28
2 24452 1 28
2 24453 1 28
2 24454 1 28
2 24455 1 28
2 24456 1 28
2 24457 1 28
2 24458 1 28
2 24459 1 28
2 24460 1 28
2 24461 1 28
2 24462 1 28
2 24463 1 28
2 24464 1 28
2 24465 1 28
2 24466 1 28
2 24467 1 28
2 24468 1 28
2 24469 1 28
2 24470 1 28
2 24471 1 28
2 24472 1 28
2 24473 1 28
2 24474 1 28
2 24475 1 28
2 24476 1 28
2 24477 1 28
2 24478 1 28
2 24479 1 28
2 24480 1 28
2 24481 1 28
2 24482 1 28
2 24483 1 28
2 24484 1 28
2 24485 1 28
2 24486 1 28
2 24487 1 28
2 24488 1 28
2 24489 1 28
2 24490 1 28
2 24491 1 28
2 24492 1 28
2 24493 1 28
2 24494 1 28
2 24495 1 28
2 24496 1 28
2 24497 1 28
2 24498 1 28
2 24499 1 28
2 24500 1 28
2 24501 1 28
2 24502 1 28
2 24503 1 28
2 24504 1 28
2 24505 1 28
2 24506 1 28
2 24507 1 28
2 24508 1 28
2 24509 1 28
2 24510 1 28
2 24511 1 28
2 24512 1 28
2 24513 1 28
2 24514 1 28
2 24515 1 28
2 24516 1 28
2 24517 1 28
2 24518 1 28
2 24519 1 28
2 24520 1 28
2 24521 1 28
2 24522 1 28
2 24523 1 28
2 24524 1 29
2 24525 1 29
2 24526 1 29
2 24527 1 29
2 24528 1 29
2 24529 1 29
2 24530 1 29
2 24531 1 29
2 24532 1 29
2 24533 1 29
2 24534 1 29
2 24535 1 29
2 24536 1 29
2 24537 1 29
2 24538 1 29
2 24539 1 29
2 24540 1 29
2 24541 1 29
2 24542 1 29
2 24543 1 29
2 24544 1 29
2 24545 1 29
2 24546 1 29
2 24547 1 29
2 24548 1 29
2 24549 1 29
2 24550 1 29
2 24551 1 29
2 24552 1 29
2 24553 1 29
2 24554 1 29
2 24555 1 29
2 24556 1 29
2 24557 1 29
2 24558 1 29
2 24559 1 29
2 24560 1 29
2 24561 1 29
2 24562 1 29
2 24563 1 29
2 24564 1 29
2 24565 1 29
2 24566 1 29
2 24567 1 29
2 24568 1 29
2 24569 1 29
2 24570 1 29
2 24571 1 29
2 24572 1 29
2 24573 1 29
2 24574 1 29
2 24575 1 29
2 24576 1 29
2 24577 1 29
2 24578 1 29
2 24579 1 29
2 24580 1 29
2 24581 1 29
2 24582 1 29
2 24583 1 29
2 24584 1 29
2 24585 1 29
2 24586 1 29
2 24587 1 29
2 24588 1 29
2 24589 1 29
2 24590 1 29
2 24591 1 29
2 24592 1 29
2 24593 1 29
2 24594 1 29
2 24595 1 29
2 24596 1 29
2 24597 1 29
2 24598 1 29
2 24599 1 29
2 24600 1 29
2 24601 1 29
2 24602 1 29
2 24603 1 29
2 24604 1 29
2 24605 1 29
2 24606 1 29
2 24607 1 29
2 24608 1 29
2 24609 1 29
2 24610 1 29
2 24611 1 29
2 24612 1 29
2 24613 1 29
2 24614 1 29
2 24615 1 29
2 24616 1 29
2 24617 1 29
2 24618 1 29
2 24619 1 29
2 24620 1 29
2 24621 1 29
2 24622 1 29
2 24623 1 29
2 24624 1 29
2 24625 1 29
2 24626 1 30
2 24627 1 30
2 24628 1 30
2 24629 1 30
2 24630 1 30
2 24631 1 30
2 24632 1 30
2 24633 1 30
2 24634 1 30
2 24635 1 30
2 24636 1 30
2 24637 1 30
2 24638 1 30
2 24639 1 30
2 24640 1 30
2 24641 1 30
2 24642 1 30
2 24643 1 30
2 24644 1 30
2 24645 1 30
2 24646 1 30
2 24647 1 30
2 24648 1 30
2 24649 1 30
2 24650 1 30
2 24651 1 30
2 24652 1 30
2 24653 1 30
2 24654 1 30
2 24655 1 30
2 24656 1 30
2 24657 1 30
2 24658 1 30
2 24659 1 30
2 24660 1 30
2 24661 1 30
2 24662 1 30
2 24663 1 30
2 24664 1 30
2 24665 1 30
2 24666 1 30
2 24667 1 30
2 24668 1 30
2 24669 1 30
2 24670 1 30
2 24671 1 30
2 24672 1 30
2 24673 1 30
2 24674 1 30
2 24675 1 30
2 24676 1 30
2 24677 1 30
2 24678 1 30
2 24679 1 30
2 24680 1 30
2 24681 1 30
2 24682 1 30
2 24683 1 30
2 24684 1 30
2 24685 1 30
2 24686 1 30
2 24687 1 30
2 24688 1 30
2 24689 1 30
2 24690 1 30
2 24691 1 30
2 24692 1 30
2 24693 1 30
2 24694 1 30
2 24695 1 30
2 24696 1 30
2 24697 1 30
2 24698 1 30
2 24699 1 30
2 24700 1 30
2 24701 1 30
2 24702 1 30
2 24703 1 30
2 24704 1 30
2 24705 1 30
2 24706 1 30
2 24707 1 30
2 24708 1 30
2 24709 1 30
2 24710 1 30
2 24711 1 30
2 24712 1 30
2 24713 1 30
2 24714 1 30
2 24715 1 30
2 24716 1 30
2 24717 1 30
2 24718 1 30
2 24719 1 30
2 24720 1 31
2 24721 1 31
2 24722 1 31
2 24723 1 31
2 24724 1 31
2 24725 1 31
2 24726 1 31
2 24727 1 31
2 24728 1 31
2 24729 1 31
2 24730 1 31
2 24731 1 31
2 24732 1 31
2 24733 1 31
2 24734 1 31
2 24735 1 31
2 24736 1 31
2 24737 1 31
2 24738 1 31
2 24739 1 31
2 24740 1 31
2 24741 1 31
2 24742 1 31
2 24743 1 31
2 24744 1 31
2 24745 1 31
2 24746 1 31
2 24747 1 31
2 24748 1 31
2 24749 1 31
2 24750 1 31
2 24751 1 31
2 24752 1 31
2 24753 1 31
2 24754 1 31
2 24755 1 31
2 24756 1 31
2 24757 1 31
2 24758 1 31
2 24759 1 31
2 24760 1 31
2 24761 1 31
2 24762 1 31
2 24763 1 31
2 24764 1 31
2 24765 1 31
2 24766 1 31
2 24767 1 31
2 24768 1 31
2 24769 1 31
2 24770 1 31
2 24771 1 31
2 24772 1 31
2 24773 1 31
2 24774 1 31
2 24775 1 31
2 24776 1 31
2 24777 1 31
2 24778 1 31
2 24779 1 31
2 24780 1 31
2 24781 1 31
2 24782 1 31
2 24783 1 31
2 24784 1 31
2 24785 1 31
2 24786 1 31
2 24787 1 31
2 24788 1 31
2 24789 1 31
2 24790 1 31
2 24791 1 31
2 24792 1 31
2 24793 1 31
2 24794 1 31
2 24795 1 31
2 24796 1 31
2 24797 1 31
2 24798 1 31
2 24799 1 31
2 24800 1 31
2 24801 1 31
2 24802 1 31
2 24803 1 31
2 24804 1 31
2 24805 1 32
2 24806 1 32
2 24807 1 32
2 24808 1 32
2 24809 1 32
2 24810 1 32
2 24811 1 32
2 24812 1 32
2 24813 1 32
2 24814 1 32
2 24815 1 32
2 24816 1 32
2 24817 1 32
2 24818 1 32
2 24819 1 32
2 24820 1 32
2 24821 1 32
2 24822 1 32
2 24823 1 32
2 24824 1 32
2 24825 1 32
2 24826 1 32
2 24827 1 32
2 24828 1 32
2 24829 1 32
2 24830 1 32
2 24831 1 32
2 24832 1 32
2 24833 1 32
2 24834 1 32
2 24835 1 32
2 24836 1 32
2 24837 1 32
2 24838 1 32
2 24839 1 32
2 24840 1 32
2 24841 1 32
2 24842 1 32
2 24843 1 32
2 24844 1 32
2 24845 1 32
2 24846 1 32
2 24847 1 32
2 24848 1 32
2 24849 1 32
2 24850 1 32
2 24851 1 32
2 24852 1 32
2 24853 1 32
2 24854 1 32
2 24855 1 32
2 24856 1 32
2 24857 1 32
2 24858 1 32
2 24859 1 32
2 24860 1 32
2 24861 1 32
2 24862 1 32
2 24863 1 32
2 24864 1 32
2 24865 1 32
2 24866 1 32
2 24867 1 32
2 24868 1 32
2 24869 1 32
2 24870 1 32
2 24871 1 32
2 24872 1 32
2 24873 1 32
2 24874 1 32
2 24875 1 32
2 24876 1 32
2 24877 1 32
2 24878 1 32
2 24879 1 32
2 24880 1 32
2 24881 1 32
2 24882 1 32
2 24883 1 32
2 24884 1 32
2 24885 1 32
2 24886 1 32
2 24887 1 32
2 24888 1 32
2 24889 1 32
2 24890 1 32
2 24891 1 32
2 24892 1 32
2 24893 1 32
2 24894 1 32
2 24895 1 32
2 24896 1 32
2 24897 1 32
2 24898 1 32
2 24899 1 32
2 24900 1 32
2 24901 1 32
2 24902 1 32
2 24903 1 32
2 24904 1 32
2 24905 1 32
2 24906 1 32
2 24907 1 32
2 24908 1 32
2 24909 1 32
2 24910 1 32
2 24911 1 32
2 24912 1 32
2 24913 1 32
2 24914 1 32
2 24915 1 32
2 24916 1 32
2 24917 1 32
2 24918 1 32
2 24919 1 32
2 24920 1 32
2 24921 1 32
2 24922 1 32
2 24923 1 32
2 24924 1 32
2 24925 1 32
2 24926 1 32
2 24927 1 32
2 24928 1 32
2 24929 1 32
2 24930 1 32
2 24931 1 33
2 24932 1 33
2 24933 1 33
2 24934 1 33
2 24935 1 33
2 24936 1 33
2 24937 1 33
2 24938 1 33
2 24939 1 33
2 24940 1 33
2 24941 1 33
2 24942 1 33
2 24943 1 33
2 24944 1 33
2 24945 1 33
2 24946 1 33
2 24947 1 33
2 24948 1 33
2 24949 1 33
2 24950 1 33
2 24951 1 33
2 24952 1 33
2 24953 1 33
2 24954 1 33
2 24955 1 33
2 24956 1 33
2 24957 1 33
2 24958 1 33
2 24959 1 33
2 24960 1 33
2 24961 1 33
2 24962 1 33
2 24963 1 33
2 24964 1 33
2 24965 1 33
2 24966 1 33
2 24967 1 33
2 24968 1 33
2 24969 1 33
2 24970 1 33
2 24971 1 33
2 24972 1 33
2 24973 1 33
2 24974 1 33
2 24975 1 33
2 24976 1 33
2 24977 1 33
2 24978 1 33
2 24979 1 33
2 24980 1 33
2 24981 1 33
2 24982 1 33
2 24983 1 33
2 24984 1 33
2 24985 1 33
2 24986 1 33
2 24987 1 33
2 24988 1 33
2 24989 1 33
2 24990 1 33
2 24991 1 33
2 24992 1 33
2 24993 1 33
2 24994 1 33
2 24995 1 33
2 24996 1 33
2 24997 1 33
2 24998 1 33
2 24999 1 33
2 25000 1 33
2 25001 1 33
2 25002 1 33
2 25003 1 33
2 25004 1 33
2 25005 1 33
2 25006 1 33
2 25007 1 34
2 25008 1 34
2 25009 1 34
2 25010 1 34
2 25011 1 34
2 25012 1 34
2 25013 1 34
2 25014 1 34
2 25015 1 34
2 25016 1 34
2 25017 1 34
2 25018 1 34
2 25019 1 34
2 25020 1 34
2 25021 1 34
2 25022 1 34
2 25023 1 34
2 25024 1 34
2 25025 1 34
2 25026 1 34
2 25027 1 34
2 25028 1 34
2 25029 1 34
2 25030 1 34
2 25031 1 34
2 25032 1 34
2 25033 1 34
2 25034 1 34
2 25035 1 34
2 25036 1 34
2 25037 1 34
2 25038 1 34
2 25039 1 34
2 25040 1 34
2 25041 1 34
2 25042 1 34
2 25043 1 34
2 25044 1 34
2 25045 1 34
2 25046 1 34
2 25047 1 34
2 25048 1 34
2 25049 1 34
2 25050 1 34
2 25051 1 34
2 25052 1 34
2 25053 1 34
2 25054 1 34
2 25055 1 34
2 25056 1 34
2 25057 1 34
2 25058 1 34
2 25059 1 34
2 25060 1 34
2 25061 1 34
2 25062 1 34
2 25063 1 34
2 25064 1 34
2 25065 1 34
2 25066 1 34
2 25067 1 34
2 25068 1 34
2 25069 1 34
2 25070 1 34
2 25071 1 34
2 25072 1 34
2 25073 1 34
2 25074 1 34
2 25075 1 34
2 25076 1 34
2 25077 1 34
2 25078 1 34
2 25079 1 34
2 25080 1 34
2 25081 1 34
2 25082 1 34
2 25083 1 34
2 25084 1 34
2 25085 1 34
2 25086 1 34
2 25087 1 34
2 25088 1 34
2 25089 1 34
2 25090 1 34
2 25091 1 34
2 25092 1 34
2 25093 1 34
2 25094 1 34
2 25095 1 34
2 25096 1 34
2 25097 1 34
2 25098 1 34
2 25099 1 34
2 25100 1 34
2 25101 1 34
2 25102 1 34
2 25103 1 34
2 25104 1 34
2 25105 1 34
2 25106 1 34
2 25107 1 35
2 25108 1 35
2 25109 1 35
2 25110 1 35
2 25111 1 35
2 25112 1 35
2 25113 1 35
2 25114 1 35
2 25115 1 35
2 25116 1 35
2 25117 1 35
2 25118 1 35
2 25119 1 35
2 25120 1 35
2 25121 1 35
2 25122 1 35
2 25123 1 35
2 25124 1 35
2 25125 1 35
2 25126 1 35
2 25127 1 35
2 25128 1 35
2 25129 1 35
2 25130 1 35
2 25131 1 35
2 25132 1 35
2 25133 1 35
2 25134 1 35
2 25135 1 35
2 25136 1 35
2 25137 1 35
2 25138 1 35
2 25139 1 35
2 25140 1 35
2 25141 1 35
2 25142 1 35
2 25143 1 35
2 25144 1 35
2 25145 1 35
2 25146 1 35
2 25147 1 35
2 25148 1 35
2 25149 1 35
2 25150 1 35
2 25151 1 35
2 25152 1 35
2 25153 1 35
2 25154 1 35
2 25155 1 35
2 25156 1 35
2 25157 1 35
2 25158 1 35
2 25159 1 35
2 25160 1 35
2 25161 1 35
2 25162 1 35
2 25163 1 36
2 25164 1 36
2 25165 1 36
2 25166 1 36
2 25167 1 36
2 25168 1 36
2 25169 1 36
2 25170 1 36
2 25171 1 36
2 25172 1 36
2 25173 1 36
2 25174 1 36
2 25175 1 36
2 25176 1 36
2 25177 1 36
2 25178 1 36
2 25179 1 36
2 25180 1 36
2 25181 1 36
2 25182 1 36
2 25183 1 36
2 25184 1 36
2 25185 1 36
2 25186 1 36
2 25187 1 36
2 25188 1 36
2 25189 1 36
2 25190 1 36
2 25191 1 36
2 25192 1 36
2 25193 1 36
2 25194 1 36
2 25195 1 36
2 25196 1 36
2 25197 1 36
2 25198 1 36
2 25199 1 36
2 25200 1 36
2 25201 1 36
2 25202 1 36
2 25203 1 36
2 25204 1 36
2 25205 1 36
2 25206 1 36
2 25207 1 36
2 25208 1 36
2 25209 1 36
2 25210 1 36
2 25211 1 36
2 25212 1 36
2 25213 1 36
2 25214 1 36
2 25215 1 36
2 25216 1 36
2 25217 1 36
2 25218 1 36
2 25219 1 36
2 25220 1 36
2 25221 1 36
2 25222 1 36
2 25223 1 36
2 25224 1 36
2 25225 1 36
2 25226 1 36
2 25227 1 36
2 25228 1 36
2 25229 1 36
2 25230 1 36
2 25231 1 36
2 25232 1 36
2 25233 1 36
2 25234 1 36
2 25235 1 36
2 25236 1 36
2 25237 1 36
2 25238 1 36
2 25239 1 36
2 25240 1 36
2 25241 1 36
2 25242 1 36
2 25243 1 36
2 25244 1 36
2 25245 1 36
2 25246 1 36
2 25247 1 36
2 25248 1 37
2 25249 1 37
2 25250 1 37
2 25251 1 37
2 25252 1 37
2 25253 1 37
2 25254 1 37
2 25255 1 37
2 25256 1 37
2 25257 1 37
2 25258 1 37
2 25259 1 37
2 25260 1 37
2 25261 1 37
2 25262 1 37
2 25263 1 37
2 25264 1 37
2 25265 1 37
2 25266 1 37
2 25267 1 37
2 25268 1 37
2 25269 1 37
2 25270 1 37
2 25271 1 37
2 25272 1 37
2 25273 1 37
2 25274 1 37
2 25275 1 37
2 25276 1 37
2 25277 1 37
2 25278 1 37
2 25279 1 37
2 25280 1 37
2 25281 1 37
2 25282 1 37
2 25283 1 37
2 25284 1 37
2 25285 1 37
2 25286 1 37
2 25287 1 37
2 25288 1 37
2 25289 1 37
2 25290 1 37
2 25291 1 37
2 25292 1 37
2 25293 1 37
2 25294 1 37
2 25295 1 37
2 25296 1 37
2 25297 1 37
2 25298 1 37
2 25299 1 37
2 25300 1 37
2 25301 1 37
2 25302 1 37
2 25303 1 37
2 25304 1 37
2 25305 1 37
2 25306 1 37
2 25307 1 37
2 25308 1 37
2 25309 1 37
2 25310 1 37
2 25311 1 37
2 25312 1 37
2 25313 1 37
2 25314 1 37
2 25315 1 37
2 25316 1 37
2 25317 1 37
2 25318 1 37
2 25319 1 37
2 25320 1 37
2 25321 1 37
2 25322 1 37
2 25323 1 37
2 25324 1 37
2 25325 1 37
2 25326 1 37
2 25327 1 38
2 25328 1 38
2 25329 1 38
2 25330 1 38
2 25331 1 38
2 25332 1 38
2 25333 1 38
2 25334 1 38
2 25335 1 38
2 25336 1 38
2 25337 1 38
2 25338 1 38
2 25339 1 38
2 25340 1 38
2 25341 1 38
2 25342 1 38
2 25343 1 38
2 25344 1 38
2 25345 1 38
2 25346 1 38
2 25347 1 38
2 25348 1 38
2 25349 1 38
2 25350 1 38
2 25351 1 38
2 25352 1 38
2 25353 1 38
2 25354 1 38
2 25355 1 38
2 25356 1 38
2 25357 1 38
2 25358 1 38
2 25359 1 38
2 25360 1 38
2 25361 1 38
2 25362 1 38
2 25363 1 38
2 25364 1 38
2 25365 1 38
2 25366 1 38
2 25367 1 38
2 25368 1 38
2 25369 1 38
2 25370 1 38
2 25371 1 38
2 25372 1 38
2 25373 1 38
2 25374 1 38
2 25375 1 38
2 25376 1 38
2 25377 1 38
2 25378 1 38
2 25379 1 38
2 25380 1 38
2 25381 1 38
2 25382 1 38
2 25383 1 38
2 25384 1 38
2 25385 1 38
2 25386 1 38
2 25387 1 38
2 25388 1 38
2 25389 1 38
2 25390 1 38
2 25391 1 38
2 25392 1 38
2 25393 1 38
2 25394 1 38
2 25395 1 38
2 25396 1 39
2 25397 1 39
2 25398 1 39
2 25399 1 39
2 25400 1 39
2 25401 1 39
2 25402 1 39
2 25403 1 39
2 25404 1 39
2 25405 1 39
2 25406 1 39
2 25407 1 39
2 25408 1 39
2 25409 1 39
2 25410 1 39
2 25411 1 39
2 25412 1 39
2 25413 1 39
2 25414 1 39
2 25415 1 39
2 25416 1 39
2 25417 1 39
2 25418 1 39
2 25419 1 39
2 25420 1 39
2 25421 1 39
2 25422 1 39
2 25423 1 39
2 25424 1 39
2 25425 1 39
2 25426 1 39
2 25427 1 39
2 25428 1 39
2 25429 1 39
2 25430 1 39
2 25431 1 39
2 25432 1 39
2 25433 1 39
2 25434 1 39
2 25435 1 39
2 25436 1 39
2 25437 1 39
2 25438 1 39
2 25439 1 39
2 25440 1 39
2 25441 1 39
2 25442 1 39
2 25443 1 39
2 25444 1 39
2 25445 1 39
2 25446 1 39
2 25447 1 39
2 25448 1 39
2 25449 1 39
2 25450 1 39
2 25451 1 40
2 25452 1 40
2 25453 1 40
2 25454 1 40
2 25455 1 40
2 25456 1 40
2 25457 1 40
2 25458 1 40
2 25459 1 40
2 25460 1 40
2 25461 1 40
2 25462 1 40
2 25463 1 40
2 25464 1 40
2 25465 1 40
2 25466 1 40
2 25467 1 40
2 25468 1 40
2 25469 1 40
2 25470 1 40
2 25471 1 40
2 25472 1 40
2 25473 1 40
2 25474 1 40
2 25475 1 40
2 25476 1 40
2 25477 1 40
2 25478 1 40
2 25479 1 40
2 25480 1 40
2 25481 1 40
2 25482 1 40
2 25483 1 40
2 25484 1 40
2 25485 1 40
2 25486 1 40
2 25487 1 40
2 25488 1 40
2 25489 1 40
2 25490 1 40
2 25491 1 40
2 25492 1 40
2 25493 1 40
2 25494 1 40
2 25495 1 40
2 25496 1 40
2 25497 1 40
2 25498 1 40
2 25499 1 40
2 25500 1 40
2 25501 1 40
2 25502 1 40
2 25503 1 40
2 25504 1 40
2 25505 1 40
2 25506 1 40
2 25507 1 40
2 25508 1 40
2 25509 1 40
2 25510 1 40
2 25511 1 40
2 25512 1 40
2 25513 1 40
2 25514 1 40
2 25515 1 40
2 25516 1 40
2 25517 1 40
2 25518 1 41
2 25519 1 41
2 25520 1 41
2 25521 1 41
2 25522 1 41
2 25523 1 41
2 25524 1 41
2 25525 1 41
2 25526 1 41
2 25527 1 41
2 25528 1 41
2 25529 1 41
2 25530 1 41
2 25531 1 41
2 25532 1 41
2 25533 1 41
2 25534 1 41
2 25535 1 41
2 25536 1 41
2 25537 1 41
2 25538 1 41
2 25539 1 41
2 25540 1 41
2 25541 1 41
2 25542 1 41
2 25543 1 41
2 25544 1 41
2 25545 1 41
2 25546 1 41
2 25547 1 41
2 25548 1 41
2 25549 1 41
2 25550 1 41
2 25551 1 41
2 25552 1 41
2 25553 1 41
2 25554 1 41
2 25555 1 41
2 25556 1 41
2 25557 1 41
2 25558 1 41
2 25559 1 41
2 25560 1 41
2 25561 1 41
2 25562 1 41
2 25563 1 41
2 25564 1 41
2 25565 1 41
2 25566 1 41
2 25567 1 41
2 25568 1 41
2 25569 1 41
2 25570 1 41
2 25571 1 41
2 25572 1 41
2 25573 1 41
2 25574 1 41
2 25575 1 41
2 25576 1 41
2 25577 1 41
2 25578 1 41
2 25579 1 41
2 25580 1 41
2 25581 1 41
2 25582 1 41
2 25583 1 41
2 25584 1 41
2 25585 1 41
2 25586 1 41
2 25587 1 41
2 25588 1 41
2 25589 1 42
2 25590 1 42
2 25591 1 42
2 25592 1 42
2 25593 1 42
2 25594 1 42
2 25595 1 42
2 25596 1 42
2 25597 1 42
2 25598 1 42
2 25599 1 42
2 25600 1 42
2 25601 1 42
2 25602 1 42
2 25603 1 42
2 25604 1 42
2 25605 1 42
2 25606 1 42
2 25607 1 42
2 25608 1 42
2 25609 1 42
2 25610 1 42
2 25611 1 42
2 25612 1 42
2 25613 1 42
2 25614 1 42
2 25615 1 42
2 25616 1 42
2 25617 1 42
2 25618 1 42
2 25619 1 42
2 25620 1 42
2 25621 1 42
2 25622 1 42
2 25623 1 42
2 25624 1 42
2 25625 1 42
2 25626 1 42
2 25627 1 42
2 25628 1 42
2 25629 1 42
2 25630 1 42
2 25631 1 42
2 25632 1 42
2 25633 1 42
2 25634 1 42
2 25635 1 42
2 25636 1 42
2 25637 1 42
2 25638 1 42
2 25639 1 42
2 25640 1 42
2 25641 1 42
2 25642 1 42
2 25643 1 42
2 25644 1 42
2 25645 1 42
2 25646 1 42
2 25647 1 44
2 25648 1 44
2 25649 1 44
2 25650 1 44
2 25651 1 44
2 25652 1 44
2 25653 1 44
2 25654 1 44
2 25655 1 44
2 25656 1 44
2 25657 1 44
2 25658 1 44
2 25659 1 44
2 25660 1 44
2 25661 1 44
2 25662 1 44
2 25663 1 44
2 25664 1 44
2 25665 1 44
2 25666 1 44
2 25667 1 44
2 25668 1 44
2 25669 1 44
2 25670 1 44
2 25671 1 44
2 25672 1 44
2 25673 1 44
2 25674 1 44
2 25675 1 44
2 25676 1 44
2 25677 1 44
2 25678 1 44
2 25679 1 44
2 25680 1 44
2 25681 1 44
2 25682 1 44
2 25683 1 44
2 25684 1 44
2 25685 1 44
2 25686 1 44
2 25687 1 44
2 25688 1 44
2 25689 1 44
2 25690 1 44
2 25691 1 44
2 25692 1 44
2 25693 1 44
2 25694 1 44
2 25695 1 44
2 25696 1 44
2 25697 1 44
2 25698 1 44
2 25699 1 44
2 25700 1 44
2 25701 1 44
2 25702 1 44
2 25703 1 44
2 25704 1 44
2 25705 1 44
2 25706 1 44
2 25707 1 44
2 25708 1 44
2 25709 1 44
2 25710 1 44
2 25711 1 44
2 25712 1 44
2 25713 1 44
2 25714 1 44
2 25715 1 44
2 25716 1 44
2 25717 1 44
2 25718 1 44
2 25719 1 44
2 25720 1 44
2 25721 1 45
2 25722 1 45
2 25723 1 45
2 25724 1 45
2 25725 1 45
2 25726 1 45
2 25727 1 45
2 25728 1 45
2 25729 1 45
2 25730 1 45
2 25731 1 45
2 25732 1 45
2 25733 1 45
2 25734 1 45
2 25735 1 45
2 25736 1 45
2 25737 1 45
2 25738 1 45
2 25739 1 45
2 25740 1 45
2 25741 1 45
2 25742 1 45
2 25743 1 45
2 25744 1 45
2 25745 1 45
2 25746 1 45
2 25747 1 45
2 25748 1 45
2 25749 1 45
2 25750 1 45
2 25751 1 45
2 25752 1 45
2 25753 1 45
2 25754 1 45
2 25755 1 45
2 25756 1 45
2 25757 1 45
2 25758 1 45
2 25759 1 45
2 25760 1 45
2 25761 1 45
2 25762 1 45
2 25763 1 45
2 25764 1 45
2 25765 1 45
2 25766 1 45
2 25767 1 45
2 25768 1 45
2 25769 1 45
2 25770 1 45
2 25771 1 45
2 25772 1 45
2 25773 1 45
2 25774 1 45
2 25775 1 45
2 25776 1 45
2 25777 1 45
2 25778 1 45
2 25779 1 45
2 25780 1 45
2 25781 1 45
2 25782 1 45
2 25783 1 45
2 25784 1 45
2 25785 1 45
2 25786 1 45
2 25787 1 45
2 25788 1 45
2 25789 1 45
2 25790 1 45
2 25791 1 45
2 25792 1 45
2 25793 1 45
2 25794 1 45
2 25795 1 45
2 25796 1 45
2 25797 1 45
2 25798 1 45
2 25799 1 45
2 25800 1 45
2 25801 1 45
2 25802 1 45
2 25803 1 45
2 25804 1 45
2 25805 1 45
2 25806 1 45
2 25807 1 45
2 25808 1 45
2 25809 1 45
2 25810 1 45
2 25811 1 45
2 25812 1 45
2 25813 1 45
2 25814 1 45
2 25815 1 45
2 25816 1 45
2 25817 1 45
2 25818 1 45
2 25819 1 45
2 25820 1 45
2 25821 1 45
2 25822 1 45
2 25823 1 45
2 25824 1 45
2 25825 1 45
2 25826 1 45
2 25827 1 45
2 25828 1 45
2 25829 1 45
2 25830 1 45
2 25831 1 45
2 25832 1 45
2 25833 1 45
2 25834 1 46
2 25835 1 46
2 25836 1 46
2 25837 1 46
2 25838 1 46
2 25839 1 46
2 25840 1 46
2 25841 1 46
2 25842 1 46
2 25843 1 46
2 25844 1 46
2 25845 1 46
2 25846 1 46
2 25847 1 46
2 25848 1 46
2 25849 1 46
2 25850 1 46
2 25851 1 46
2 25852 1 46
2 25853 1 46
2 25854 1 46
2 25855 1 46
2 25856 1 46
2 25857 1 46
2 25858 1 46
2 25859 1 46
2 25860 1 46
2 25861 1 46
2 25862 1 46
2 25863 1 46
2 25864 1 46
2 25865 1 46
2 25866 1 46
2 25867 1 46
2 25868 1 46
2 25869 1 46
2 25870 1 46
2 25871 1 46
2 25872 1 46
2 25873 1 46
2 25874 1 46
2 25875 1 46
2 25876 1 46
2 25877 1 46
2 25878 1 46
2 25879 1 46
2 25880 1 46
2 25881 1 46
2 25882 1 46
2 25883 1 46
2 25884 1 46
2 25885 1 46
2 25886 1 46
2 25887 1 46
2 25888 1 46
2 25889 1 46
2 25890 1 46
2 25891 1 46
2 25892 1 46
2 25893 1 46
2 25894 1 46
2 25895 1 46
2 25896 1 46
2 25897 1 46
2 25898 1 46
2 25899 1 46
2 25900 1 46
2 25901 1 46
2 25902 1 46
2 25903 1 46
2 25904 1 46
2 25905 1 46
2 25906 1 46
2 25907 1 46
2 25908 1 46
2 25909 1 46
2 25910 1 46
2 25911 1 46
2 25912 1 46
2 25913 1 46
2 25914 1 46
2 25915 1 46
2 25916 1 46
2 25917 1 46
2 25918 1 46
2 25919 1 46
2 25920 1 46
2 25921 1 46
2 25922 1 46
2 25923 1 46
2 25924 1 46
2 25925 1 46
2 25926 1 46
2 25927 1 46
2 25928 1 46
2 25929 1 46
2 25930 1 46
2 25931 1 46
2 25932 1 47
2 25933 1 47
2 25934 1 47
2 25935 1 47
2 25936 1 47
2 25937 1 47
2 25938 1 47
2 25939 1 47
2 25940 1 47
2 25941 1 47
2 25942 1 47
2 25943 1 47
2 25944 1 47
2 25945 1 47
2 25946 1 47
2 25947 1 47
2 25948 1 47
2 25949 1 47
2 25950 1 47
2 25951 1 47
2 25952 1 47
2 25953 1 47
2 25954 1 47
2 25955 1 47
2 25956 1 47
2 25957 1 47
2 25958 1 47
2 25959 1 47
2 25960 1 47
2 25961 1 47
2 25962 1 47
2 25963 1 47
2 25964 1 47
2 25965 1 47
2 25966 1 47
2 25967 1 47
2 25968 1 47
2 25969 1 47
2 25970 1 47
2 25971 1 47
2 25972 1 47
2 25973 1 47
2 25974 1 47
2 25975 1 47
2 25976 1 47
2 25977 1 47
2 25978 1 47
2 25979 1 47
2 25980 1 47
2 25981 1 47
2 25982 1 47
2 25983 1 47
2 25984 1 47
2 25985 1 47
2 25986 1 47
2 25987 1 47
2 25988 1 47
2 25989 1 47
2 25990 1 47
2 25991 1 47
2 25992 1 47
2 25993 1 47
2 25994 1 47
2 25995 1 47
2 25996 1 47
2 25997 1 47
2 25998 1 47
2 25999 1 47
2 26000 1 47
2 26001 1 47
2 26002 1 47
2 26003 1 47
2 26004 1 47
2 26005 1 47
2 26006 1 47
2 26007 1 47
2 26008 1 47
2 26009 1 47
2 26010 1 47
2 26011 1 47
2 26012 1 47
2 26013 1 47
2 26014 1 47
2 26015 1 47
2 26016 1 47
2 26017 1 47
2 26018 1 47
2 26019 1 47
2 26020 1 47
2 26021 1 48
2 26022 1 48
2 26023 1 48
2 26024 1 48
2 26025 1 48
2 26026 1 48
2 26027 1 48
2 26028 1 48
2 26029 1 48
2 26030 1 48
2 26031 1 48
2 26032 1 48
2 26033 1 48
2 26034 1 48
2 26035 1 48
2 26036 1 48
2 26037 1 48
2 26038 1 48
2 26039 1 48
2 26040 1 48
2 26041 1 48
2 26042 1 48
2 26043 1 48
2 26044 1 48
2 26045 1 48
2 26046 1 48
2 26047 1 48
2 26048 1 48
2 26049 1 48
2 26050 1 48
2 26051 1 48
2 26052 1 48
2 26053 1 48
2 26054 1 48
2 26055 1 48
2 26056 1 48
2 26057 1 48
2 26058 1 48
2 26059 1 48
2 26060 1 48
2 26061 1 48
2 26062 1 48
2 26063 1 48
2 26064 1 48
2 26065 1 48
2 26066 1 48
2 26067 1 48
2 26068 1 48
2 26069 1 48
2 26070 1 48
2 26071 1 48
2 26072 1 48
2 26073 1 48
2 26074 1 48
2 26075 1 48
2 26076 1 48
2 26077 1 48
2 26078 1 48
2 26079 1 48
2 26080 1 48
2 26081 1 48
2 26082 1 48
2 26083 1 48
2 26084 1 48
2 26085 1 48
2 26086 1 48
2 26087 1 48
2 26088 1 48
2 26089 1 48
2 26090 1 48
2 26091 1 48
2 26092 1 48
2 26093 1 48
2 26094 1 48
2 26095 1 48
2 26096 1 48
2 26097 1 48
2 26098 1 48
2 26099 1 48
2 26100 1 48
2 26101 1 48
2 26102 1 48
2 26103 1 48
2 26104 1 48
2 26105 1 48
2 26106 1 48
2 26107 1 48
2 26108 1 48
2 26109 1 48
2 26110 1 48
2 26111 1 49
2 26112 1 49
2 26113 1 49
2 26114 1 49
2 26115 1 49
2 26116 1 49
2 26117 1 49
2 26118 1 49
2 26119 1 49
2 26120 1 49
2 26121 1 49
2 26122 1 49
2 26123 1 49
2 26124 1 49
2 26125 1 49
2 26126 1 49
2 26127 1 49
2 26128 1 49
2 26129 1 49
2 26130 1 49
2 26131 1 49
2 26132 1 49
2 26133 1 49
2 26134 1 49
2 26135 1 49
2 26136 1 49
2 26137 1 49
2 26138 1 49
2 26139 1 49
2 26140 1 49
2 26141 1 49
2 26142 1 49
2 26143 1 49
2 26144 1 49
2 26145 1 49
2 26146 1 49
2 26147 1 49
2 26148 1 49
2 26149 1 49
2 26150 1 49
2 26151 1 49
2 26152 1 49
2 26153 1 49
2 26154 1 49
2 26155 1 49
2 26156 1 49
2 26157 1 49
2 26158 1 49
2 26159 1 49
2 26160 1 49
2 26161 1 49
2 26162 1 49
2 26163 1 49
2 26164 1 49
2 26165 1 49
2 26166 1 49
2 26167 1 49
2 26168 1 49
2 26169 1 49
2 26170 1 49
2 26171 1 49
2 26172 1 49
2 26173 1 49
2 26174 1 49
2 26175 1 49
2 26176 1 49
2 26177 1 49
2 26178 1 49
2 26179 1 49
2 26180 1 49
2 26181 1 49
2 26182 1 49
2 26183 1 49
2 26184 1 49
2 26185 1 49
2 26186 1 49
2 26187 1 49
2 26188 1 49
2 26189 1 49
2 26190 1 49
2 26191 1 49
2 26192 1 49
2 26193 1 49
2 26194 1 49
2 26195 1 49
2 26196 1 49
2 26197 1 49
2 26198 1 49
2 26199 1 49
2 26200 1 49
2 26201 1 49
2 26202 1 49
2 26203 1 49
2 26204 1 49
2 26205 1 49
2 26206 1 50
2 26207 1 50
2 26208 1 50
2 26209 1 50
2 26210 1 50
2 26211 1 50
2 26212 1 50
2 26213 1 50
2 26214 1 50
2 26215 1 50
2 26216 1 50
2 26217 1 50
2 26218 1 50
2 26219 1 50
2 26220 1 50
2 26221 1 50
2 26222 1 50
2 26223 1 50
2 26224 1 50
2 26225 1 50
2 26226 1 50
2 26227 1 50
2 26228 1 50
2 26229 1 50
2 26230 1 50
2 26231 1 50
2 26232 1 50
2 26233 1 50
2 26234 1 50
2 26235 1 50
2 26236 1 50
2 26237 1 50
2 26238 1 50
2 26239 1 50
2 26240 1 50
2 26241 1 50
2 26242 1 50
2 26243 1 50
2 26244 1 50
2 26245 1 50
2 26246 1 50
2 26247 1 50
2 26248 1 50
2 26249 1 50
2 26250 1 50
2 26251 1 50
2 26252 1 50
2 26253 1 50
2 26254 1 50
2 26255 1 50
2 26256 1 50
2 26257 1 50
2 26258 1 50
2 26259 1 50
2 26260 1 50
2 26261 1 50
2 26262 1 50
2 26263 1 50
2 26264 1 50
2 26265 1 50
2 26266 1 50
2 26267 1 50
2 26268 1 50
2 26269 1 50
2 26270 1 50
2 26271 1 50
2 26272 1 50
2 26273 1 50
2 26274 1 50
2 26275 1 50
2 26276 1 50
2 26277 1 50
2 26278 1 50
2 26279 1 50
2 26280 1 50
2 26281 1 50
2 26282 1 50
2 26283 1 51
2 26284 1 51
2 26285 1 51
2 26286 1 51
2 26287 1 51
2 26288 1 51
2 26289 1 51
2 26290 1 51
2 26291 1 51
2 26292 1 51
2 26293 1 51
2 26294 1 51
2 26295 1 51
2 26296 1 51
2 26297 1 51
2 26298 1 51
2 26299 1 51
2 26300 1 51
2 26301 1 51
2 26302 1 51
2 26303 1 51
2 26304 1 51
2 26305 1 51
2 26306 1 51
2 26307 1 51
2 26308 1 51
2 26309 1 51
2 26310 1 51
2 26311 1 51
2 26312 1 51
2 26313 1 51
2 26314 1 51
2 26315 1 51
2 26316 1 51
2 26317 1 51
2 26318 1 51
2 26319 1 51
2 26320 1 51
2 26321 1 51
2 26322 1 51
2 26323 1 51
2 26324 1 51
2 26325 1 52
2 26326 1 52
2 26327 1 52
2 26328 1 52
2 26329 1 52
2 26330 1 52
2 26331 1 52
2 26332 1 52
2 26333 1 52
2 26334 1 52
2 26335 1 52
2 26336 1 52
2 26337 1 52
2 26338 1 52
2 26339 1 52
2 26340 1 52
2 26341 1 52
2 26342 1 52
2 26343 1 52
2 26344 1 52
2 26345 1 52
2 26346 1 52
2 26347 1 52
2 26348 1 52
2 26349 1 52
2 26350 1 52
2 26351 1 52
2 26352 1 52
2 26353 1 52
2 26354 1 52
2 26355 1 52
2 26356 1 52
2 26357 1 52
2 26358 1 52
2 26359 1 52
2 26360 1 54
2 26361 1 54
2 26362 1 54
2 26363 1 54
2 26364 1 54
2 26365 1 54
2 26366 1 54
2 26367 1 54
2 26368 1 54
2 26369 1 54
2 26370 1 54
2 26371 1 54
2 26372 1 54
2 26373 1 54
2 26374 1 54
2 26375 1 54
2 26376 1 54
2 26377 1 54
2 26378 1 54
2 26379 1 54
2 26380 1 54
2 26381 1 55
2 26382 1 55
2 26383 1 55
2 26384 1 55
2 26385 1 56
2 26386 1 56
2 26387 1 56
2 26388 1 56
2 26389 1 57
2 26390 1 57
2 26391 1 58
2 26392 1 58
2 26393 1 58
2 26394 1 58
2 26395 1 58
2 26396 1 58
2 26397 1 58
2 26398 1 59
2 26399 1 59
2 26400 1 59
2 26401 1 59
2 26402 1 59
2 26403 1 59
2 26404 1 59
2 26405 1 59
2 26406 1 59
2 26407 1 59
2 26408 1 59
2 26409 1 59
2 26410 1 59
2 26411 1 59
2 26412 1 59
2 26413 1 59
2 26414 1 59
2 26415 1 59
2 26416 1 59
2 26417 1 59
2 26418 1 59
2 26419 1 60
2 26420 1 60
2 26421 1 60
2 26422 1 60
2 26423 1 60
2 26424 1 60
2 26425 1 60
2 26426 1 60
2 26427 1 60
2 26428 1 60
2 26429 1 60
2 26430 1 60
2 26431 1 60
2 26432 1 60
2 26433 1 60
2 26434 1 60
2 26435 1 60
2 26436 1 60
2 26437 1 60
2 26438 1 60
2 26439 1 60
2 26440 1 60
2 26441 1 60
2 26442 1 62
2 26443 1 62
2 26444 1 67
2 26445 1 67
2 26446 1 67
2 26447 1 67
2 26448 1 67
2 26449 1 67
2 26450 1 67
2 26451 1 67
2 26452 1 67
2 26453 1 67
2 26454 1 67
2 26455 1 67
2 26456 1 67
2 26457 1 67
2 26458 1 67
2 26459 1 67
2 26460 1 67
2 26461 1 67
2 26462 1 67
2 26463 1 67
2 26464 1 67
2 26465 1 68
2 26466 1 68
2 26467 1 68
2 26468 1 68
2 26469 1 68
2 26470 1 68
2 26471 1 68
2 26472 1 68
2 26473 1 68
2 26474 1 68
2 26475 1 68
2 26476 1 68
2 26477 1 68
2 26478 1 69
2 26479 1 69
2 26480 1 69
2 26481 1 70
2 26482 1 70
2 26483 1 70
2 26484 1 71
2 26485 1 71
2 26486 1 71
2 26487 1 71
2 26488 1 71
2 26489 1 71
2 26490 1 71
2 26491 1 71
2 26492 1 71
2 26493 1 71
2 26494 1 71
2 26495 1 71
2 26496 1 71
2 26497 1 71
2 26498 1 71
2 26499 1 71
2 26500 1 71
2 26501 1 72
2 26502 1 72
2 26503 1 72
2 26504 1 72
2 26505 1 72
2 26506 1 72
2 26507 1 72
2 26508 1 72
2 26509 1 72
2 26510 1 72
2 26511 1 72
2 26512 1 72
2 26513 1 72
2 26514 1 72
2 26515 1 72
2 26516 1 72
2 26517 1 72
2 26518 1 72
2 26519 1 72
2 26520 1 72
2 26521 1 72
2 26522 1 72
2 26523 1 72
2 26524 1 72
2 26525 1 73
2 26526 1 73
2 26527 1 73
2 26528 1 73
2 26529 1 73
2 26530 1 73
2 26531 1 73
2 26532 1 75
2 26533 1 75
2 26534 1 84
2 26535 1 84
2 26536 1 84
2 26537 1 84
2 26538 1 84
2 26539 1 84
2 26540 1 84
2 26541 1 84
2 26542 1 84
2 26543 1 85
2 26544 1 85
2 26545 1 86
2 26546 1 86
2 26547 1 86
2 26548 1 86
2 26549 1 87
2 26550 1 87
2 26551 1 87
2 26552 1 90
2 26553 1 90
2 26554 1 98
2 26555 1 98
2 26556 1 98
2 26557 1 98
2 26558 1 99
2 26559 1 99
2 26560 1 100
2 26561 1 100
2 26562 1 100
2 26563 1 100
2 26564 1 100
2 26565 1 100
2 26566 1 100
2 26567 1 100
2 26568 1 104
2 26569 1 104
2 26570 1 104
2 26571 1 104
2 26572 1 104
2 26573 1 104
2 26574 1 104
2 26575 1 104
2 26576 1 104
2 26577 1 104
2 26578 1 104
2 26579 1 104
2 26580 1 105
2 26581 1 105
2 26582 1 105
2 26583 1 105
2 26584 1 105
2 26585 1 105
2 26586 1 105
2 26587 1 105
2 26588 1 105
2 26589 1 105
2 26590 1 105
2 26591 1 105
2 26592 1 105
2 26593 1 105
2 26594 1 105
2 26595 1 105
2 26596 1 105
2 26597 1 105
2 26598 1 105
2 26599 1 105
2 26600 1 105
2 26601 1 105
2 26602 1 105
2 26603 1 105
2 26604 1 105
2 26605 1 105
2 26606 1 105
2 26607 1 106
2 26608 1 106
2 26609 1 106
2 26610 1 106
2 26611 1 106
2 26612 1 107
2 26613 1 107
2 26614 1 108
2 26615 1 108
2 26616 1 108
2 26617 1 108
2 26618 1 108
2 26619 1 108
2 26620 1 108
2 26621 1 108
2 26622 1 111
2 26623 1 111
2 26624 1 111
2 26625 1 111
2 26626 1 111
2 26627 1 111
2 26628 1 111
2 26629 1 111
2 26630 1 111
2 26631 1 111
2 26632 1 111
2 26633 1 111
2 26634 1 120
2 26635 1 120
2 26636 1 120
2 26637 1 120
2 26638 1 120
2 26639 1 120
2 26640 1 120
2 26641 1 121
2 26642 1 121
2 26643 1 121
2 26644 1 121
2 26645 1 121
2 26646 1 121
2 26647 1 121
2 26648 1 121
2 26649 1 121
2 26650 1 122
2 26651 1 122
2 26652 1 122
2 26653 1 122
2 26654 1 125
2 26655 1 125
2 26656 1 126
2 26657 1 126
2 26658 1 126
2 26659 1 126
2 26660 1 126
2 26661 1 126
2 26662 1 126
2 26663 1 126
2 26664 1 127
2 26665 1 127
2 26666 1 128
2 26667 1 128
2 26668 1 128
2 26669 1 128
2 26670 1 128
2 26671 1 128
2 26672 1 128
2 26673 1 128
2 26674 1 129
2 26675 1 129
2 26676 1 130
2 26677 1 130
2 26678 1 130
2 26679 1 130
2 26680 1 132
2 26681 1 132
2 26682 1 133
2 26683 1 133
2 26684 1 133
2 26685 1 133
2 26686 1 133
2 26687 1 133
2 26688 1 133
2 26689 1 133
2 26690 1 133
2 26691 1 136
2 26692 1 136
2 26693 1 144
2 26694 1 144
2 26695 1 144
2 26696 1 144
2 26697 1 145
2 26698 1 145
2 26699 1 145
2 26700 1 145
2 26701 1 145
2 26702 1 145
2 26703 1 145
2 26704 1 145
2 26705 1 146
2 26706 1 146
2 26707 1 146
2 26708 1 146
2 26709 1 146
2 26710 1 147
2 26711 1 147
2 26712 1 147
2 26713 1 147
2 26714 1 147
2 26715 1 149
2 26716 1 149
2 26717 1 149
2 26718 1 149
2 26719 1 156
2 26720 1 156
2 26721 1 156
2 26722 1 157
2 26723 1 157
2 26724 1 158
2 26725 1 158
2 26726 1 158
2 26727 1 159
2 26728 1 159
2 26729 1 160
2 26730 1 160
2 26731 1 160
2 26732 1 160
2 26733 1 160
2 26734 1 160
2 26735 1 160
2 26736 1 160
2 26737 1 160
2 26738 1 160
2 26739 1 160
2 26740 1 160
2 26741 1 160
2 26742 1 160
2 26743 1 160
2 26744 1 160
2 26745 1 160
2 26746 1 160
2 26747 1 160
2 26748 1 161
2 26749 1 161
2 26750 1 161
2 26751 1 161
2 26752 1 161
2 26753 1 161
2 26754 1 161
2 26755 1 161
2 26756 1 161
2 26757 1 161
2 26758 1 161
2 26759 1 161
2 26760 1 161
2 26761 1 161
2 26762 1 170
2 26763 1 170
2 26764 1 170
2 26765 1 170
2 26766 1 170
2 26767 1 170
2 26768 1 170
2 26769 1 170
2 26770 1 170
2 26771 1 170
2 26772 1 170
2 26773 1 170
2 26774 1 170
2 26775 1 170
2 26776 1 170
2 26777 1 170
2 26778 1 170
2 26779 1 172
2 26780 1 172
2 26781 1 172
2 26782 1 172
2 26783 1 172
2 26784 1 173
2 26785 1 173
2 26786 1 174
2 26787 1 174
2 26788 1 175
2 26789 1 175
2 26790 1 175
2 26791 1 175
2 26792 1 175
2 26793 1 175
2 26794 1 175
2 26795 1 175
2 26796 1 175
2 26797 1 175
2 26798 1 175
2 26799 1 175
2 26800 1 175
2 26801 1 175
2 26802 1 175
2 26803 1 175
2 26804 1 175
2 26805 1 175
2 26806 1 175
2 26807 1 175
2 26808 1 177
2 26809 1 177
2 26810 1 177
2 26811 1 178
2 26812 1 178
2 26813 1 178
2 26814 1 178
2 26815 1 178
2 26816 1 178
2 26817 1 178
2 26818 1 178
2 26819 1 178
2 26820 1 178
2 26821 1 178
2 26822 1 178
2 26823 1 178
2 26824 1 178
2 26825 1 179
2 26826 1 179
2 26827 1 179
2 26828 1 179
2 26829 1 179
2 26830 1 180
2 26831 1 180
2 26832 1 180
2 26833 1 180
2 26834 1 180
2 26835 1 187
2 26836 1 187
2 26837 1 187
2 26838 1 187
2 26839 1 187
2 26840 1 187
2 26841 1 187
2 26842 1 187
2 26843 1 188
2 26844 1 188
2 26845 1 188
2 26846 1 188
2 26847 1 188
2 26848 1 188
2 26849 1 188
2 26850 1 188
2 26851 1 188
2 26852 1 188
2 26853 1 188
2 26854 1 188
2 26855 1 188
2 26856 1 188
2 26857 1 189
2 26858 1 189
2 26859 1 197
2 26860 1 197
2 26861 1 197
2 26862 1 197
2 26863 1 197
2 26864 1 197
2 26865 1 197
2 26866 1 197
2 26867 1 199
2 26868 1 199
2 26869 1 199
2 26870 1 199
2 26871 1 199
2 26872 1 200
2 26873 1 200
2 26874 1 200
2 26875 1 200
2 26876 1 200
2 26877 1 201
2 26878 1 201
2 26879 1 210
2 26880 1 210
2 26881 1 210
2 26882 1 210
2 26883 1 210
2 26884 1 210
2 26885 1 210
2 26886 1 210
2 26887 1 210
2 26888 1 210
2 26889 1 210
2 26890 1 210
2 26891 1 210
2 26892 1 210
2 26893 1 210
2 26894 1 210
2 26895 1 210
2 26896 1 210
2 26897 1 210
2 26898 1 212
2 26899 1 212
2 26900 1 213
2 26901 1 213
2 26902 1 213
2 26903 1 213
2 26904 1 213
2 26905 1 213
2 26906 1 213
2 26907 1 213
2 26908 1 213
2 26909 1 213
2 26910 1 213
2 26911 1 213
2 26912 1 213
2 26913 1 213
2 26914 1 213
2 26915 1 213
2 26916 1 213
2 26917 1 213
2 26918 1 213
2 26919 1 213
2 26920 1 213
2 26921 1 213
2 26922 1 213
2 26923 1 213
2 26924 1 213
2 26925 1 214
2 26926 1 214
2 26927 1 214
2 26928 1 214
2 26929 1 214
2 26930 1 215
2 26931 1 215
2 26932 1 217
2 26933 1 217
2 26934 1 217
2 26935 1 217
2 26936 1 217
2 26937 1 217
2 26938 1 217
2 26939 1 217
2 26940 1 217
2 26941 1 217
2 26942 1 217
2 26943 1 217
2 26944 1 217
2 26945 1 217
2 26946 1 217
2 26947 1 217
2 26948 1 217
2 26949 1 217
2 26950 1 217
2 26951 1 217
2 26952 1 217
2 26953 1 217
2 26954 1 217
2 26955 1 217
2 26956 1 218
2 26957 1 218
2 26958 1 218
2 26959 1 218
2 26960 1 218
2 26961 1 220
2 26962 1 220
2 26963 1 220
2 26964 1 220
2 26965 1 220
2 26966 1 220
2 26967 1 220
2 26968 1 220
2 26969 1 220
2 26970 1 220
2 26971 1 220
2 26972 1 220
2 26973 1 220
2 26974 1 220
2 26975 1 220
2 26976 1 220
2 26977 1 220
2 26978 1 220
2 26979 1 221
2 26980 1 221
2 26981 1 221
2 26982 1 221
2 26983 1 221
2 26984 1 224
2 26985 1 224
2 26986 1 224
2 26987 1 224
2 26988 1 224
2 26989 1 224
2 26990 1 224
2 26991 1 224
2 26992 1 224
2 26993 1 224
2 26994 1 224
2 26995 1 224
2 26996 1 224
2 26997 1 224
2 26998 1 224
2 26999 1 224
2 27000 1 224
2 27001 1 224
2 27002 1 224
2 27003 1 224
2 27004 1 224
2 27005 1 224
2 27006 1 224
2 27007 1 228
2 27008 1 228
2 27009 1 229
2 27010 1 229
2 27011 1 229
2 27012 1 237
2 27013 1 237
2 27014 1 237
2 27015 1 237
2 27016 1 237
2 27017 1 237
2 27018 1 237
2 27019 1 237
2 27020 1 237
2 27021 1 237
2 27022 1 237
2 27023 1 237
2 27024 1 237
2 27025 1 237
2 27026 1 237
2 27027 1 237
2 27028 1 239
2 27029 1 239
2 27030 1 239
2 27031 1 239
2 27032 1 239
2 27033 1 239
2 27034 1 239
2 27035 1 239
2 27036 1 239
2 27037 1 239
2 27038 1 239
2 27039 1 239
2 27040 1 241
2 27041 1 241
2 27042 1 241
2 27043 1 241
2 27044 1 241
2 27045 1 241
2 27046 1 241
2 27047 1 241
2 27048 1 241
2 27049 1 241
2 27050 1 241
2 27051 1 241
2 27052 1 241
2 27053 1 241
2 27054 1 241
2 27055 1 242
2 27056 1 242
2 27057 1 243
2 27058 1 243
2 27059 1 243
2 27060 1 243
2 27061 1 243
2 27062 1 243
2 27063 1 243
2 27064 1 243
2 27065 1 243
2 27066 1 243
2 27067 1 243
2 27068 1 243
2 27069 1 243
2 27070 1 243
2 27071 1 243
2 27072 1 243
2 27073 1 243
2 27074 1 243
2 27075 1 243
2 27076 1 243
2 27077 1 243
2 27078 1 243
2 27079 1 243
2 27080 1 243
2 27081 1 243
2 27082 1 243
2 27083 1 243
2 27084 1 243
2 27085 1 243
2 27086 1 243
2 27087 1 243
2 27088 1 243
2 27089 1 243
2 27090 1 243
2 27091 1 243
2 27092 1 243
2 27093 1 243
2 27094 1 243
2 27095 1 250
2 27096 1 250
2 27097 1 255
2 27098 1 255
2 27099 1 256
2 27100 1 256
2 27101 1 256
2 27102 1 263
2 27103 1 263
2 27104 1 263
2 27105 1 263
2 27106 1 263
2 27107 1 263
2 27108 1 263
2 27109 1 264
2 27110 1 264
2 27111 1 264
2 27112 1 272
2 27113 1 272
2 27114 1 274
2 27115 1 274
2 27116 1 278
2 27117 1 278
2 27118 1 278
2 27119 1 288
2 27120 1 288
2 27121 1 288
2 27122 1 288
2 27123 1 288
2 27124 1 288
2 27125 1 288
2 27126 1 288
2 27127 1 288
2 27128 1 288
2 27129 1 288
2 27130 1 288
2 27131 1 288
2 27132 1 288
2 27133 1 288
2 27134 1 288
2 27135 1 288
2 27136 1 288
2 27137 1 288
2 27138 1 288
2 27139 1 288
2 27140 1 289
2 27141 1 289
2 27142 1 289
2 27143 1 289
2 27144 1 289
2 27145 1 289
2 27146 1 289
2 27147 1 289
2 27148 1 289
2 27149 1 290
2 27150 1 290
2 27151 1 290
2 27152 1 290
2 27153 1 290
2 27154 1 290
2 27155 1 290
2 27156 1 290
2 27157 1 290
2 27158 1 290
2 27159 1 291
2 27160 1 291
2 27161 1 291
2 27162 1 292
2 27163 1 292
2 27164 1 293
2 27165 1 293
2 27166 1 293
2 27167 1 293
2 27168 1 293
2 27169 1 293
2 27170 1 293
2 27171 1 293
2 27172 1 294
2 27173 1 294
2 27174 1 294
2 27175 1 294
2 27176 1 294
2 27177 1 294
2 27178 1 294
2 27179 1 294
2 27180 1 294
2 27181 1 294
2 27182 1 294
2 27183 1 295
2 27184 1 295
2 27185 1 298
2 27186 1 298
2 27187 1 298
2 27188 1 298
2 27189 1 300
2 27190 1 300
2 27191 1 306
2 27192 1 306
2 27193 1 307
2 27194 1 307
2 27195 1 307
2 27196 1 307
2 27197 1 307
2 27198 1 307
2 27199 1 307
2 27200 1 307
2 27201 1 307
2 27202 1 307
2 27203 1 307
2 27204 1 307
2 27205 1 307
2 27206 1 307
2 27207 1 307
2 27208 1 307
2 27209 1 307
2 27210 1 307
2 27211 1 307
2 27212 1 307
2 27213 1 307
2 27214 1 307
2 27215 1 307
2 27216 1 307
2 27217 1 307
2 27218 1 307
2 27219 1 307
2 27220 1 307
2 27221 1 307
2 27222 1 307
2 27223 1 307
2 27224 1 307
2 27225 1 308
2 27226 1 308
2 27227 1 308
2 27228 1 308
2 27229 1 310
2 27230 1 310
2 27231 1 310
2 27232 1 310
2 27233 1 310
2 27234 1 310
2 27235 1 310
2 27236 1 310
2 27237 1 310
2 27238 1 310
2 27239 1 310
2 27240 1 310
2 27241 1 310
2 27242 1 310
2 27243 1 310
2 27244 1 310
2 27245 1 310
2 27246 1 310
2 27247 1 310
2 27248 1 310
2 27249 1 310
2 27250 1 313
2 27251 1 313
2 27252 1 315
2 27253 1 315
2 27254 1 315
2 27255 1 315
2 27256 1 315
2 27257 1 315
2 27258 1 315
2 27259 1 315
2 27260 1 315
2 27261 1 315
2 27262 1 315
2 27263 1 315
2 27264 1 316
2 27265 1 316
2 27266 1 316
2 27267 1 316
2 27268 1 316
2 27269 1 316
2 27270 1 316
2 27271 1 316
2 27272 1 317
2 27273 1 317
2 27274 1 317
2 27275 1 317
2 27276 1 317
2 27277 1 317
2 27278 1 317
2 27279 1 317
2 27280 1 319
2 27281 1 319
2 27282 1 320
2 27283 1 320
2 27284 1 320
2 27285 1 320
2 27286 1 320
2 27287 1 320
2 27288 1 320
2 27289 1 320
2 27290 1 321
2 27291 1 321
2 27292 1 321
2 27293 1 321
2 27294 1 322
2 27295 1 322
2 27296 1 323
2 27297 1 323
2 27298 1 323
2 27299 1 323
2 27300 1 323
2 27301 1 323
2 27302 1 323
2 27303 1 323
2 27304 1 323
2 27305 1 323
2 27306 1 323
2 27307 1 323
2 27308 1 323
2 27309 1 323
2 27310 1 323
2 27311 1 323
2 27312 1 323
2 27313 1 323
2 27314 1 323
2 27315 1 323
2 27316 1 323
2 27317 1 323
2 27318 1 323
2 27319 1 323
2 27320 1 323
2 27321 1 323
2 27322 1 323
2 27323 1 323
2 27324 1 323
2 27325 1 323
2 27326 1 323
2 27327 1 323
2 27328 1 323
2 27329 1 323
2 27330 1 323
2 27331 1 324
2 27332 1 324
2 27333 1 324
2 27334 1 324
2 27335 1 324
2 27336 1 324
2 27337 1 324
2 27338 1 324
2 27339 1 324
2 27340 1 324
2 27341 1 324
2 27342 1 324
2 27343 1 324
2 27344 1 324
2 27345 1 324
2 27346 1 324
2 27347 1 325
2 27348 1 325
2 27349 1 325
2 27350 1 325
2 27351 1 325
2 27352 1 325
2 27353 1 325
2 27354 1 325
2 27355 1 325
2 27356 1 326
2 27357 1 326
2 27358 1 326
2 27359 1 336
2 27360 1 336
2 27361 1 336
2 27362 1 336
2 27363 1 336
2 27364 1 336
2 27365 1 336
2 27366 1 336
2 27367 1 344
2 27368 1 344
2 27369 1 344
2 27370 1 344
2 27371 1 344
2 27372 1 344
2 27373 1 347
2 27374 1 347
2 27375 1 347
2 27376 1 347
2 27377 1 352
2 27378 1 352
2 27379 1 355
2 27380 1 355
2 27381 1 355
2 27382 1 355
2 27383 1 355
2 27384 1 355
2 27385 1 355
2 27386 1 355
2 27387 1 355
2 27388 1 355
2 27389 1 355
2 27390 1 355
2 27391 1 355
2 27392 1 357
2 27393 1 357
2 27394 1 357
2 27395 1 357
2 27396 1 357
2 27397 1 357
2 27398 1 357
2 27399 1 357
2 27400 1 357
2 27401 1 357
2 27402 1 358
2 27403 1 358
2 27404 1 368
2 27405 1 368
2 27406 1 368
2 27407 1 368
2 27408 1 368
2 27409 1 368
2 27410 1 368
2 27411 1 368
2 27412 1 368
2 27413 1 368
2 27414 1 368
2 27415 1 368
2 27416 1 369
2 27417 1 369
2 27418 1 369
2 27419 1 369
2 27420 1 369
2 27421 1 369
2 27422 1 369
2 27423 1 369
2 27424 1 370
2 27425 1 370
2 27426 1 374
2 27427 1 374
2 27428 1 377
2 27429 1 377
2 27430 1 377
2 27431 1 377
2 27432 1 377
2 27433 1 377
2 27434 1 377
2 27435 1 377
2 27436 1 377
2 27437 1 377
2 27438 1 377
2 27439 1 377
2 27440 1 377
2 27441 1 377
2 27442 1 377
2 27443 1 378
2 27444 1 378
2 27445 1 379
2 27446 1 379
2 27447 1 379
2 27448 1 379
2 27449 1 379
2 27450 1 379
2 27451 1 379
2 27452 1 379
2 27453 1 379
2 27454 1 379
2 27455 1 379
2 27456 1 379
2 27457 1 379
2 27458 1 379
2 27459 1 379
2 27460 1 379
2 27461 1 380
2 27462 1 380
2 27463 1 391
2 27464 1 391
2 27465 1 398
2 27466 1 398
2 27467 1 398
2 27468 1 398
2 27469 1 398
2 27470 1 398
2 27471 1 399
2 27472 1 399
2 27473 1 406
2 27474 1 406
2 27475 1 406
2 27476 1 406
2 27477 1 406
2 27478 1 406
2 27479 1 406
2 27480 1 406
2 27481 1 406
2 27482 1 406
2 27483 1 406
2 27484 1 407
2 27485 1 407
2 27486 1 407
2 27487 1 407
2 27488 1 407
2 27489 1 407
2 27490 1 407
2 27491 1 407
2 27492 1 407
2 27493 1 407
2 27494 1 407
2 27495 1 407
2 27496 1 407
2 27497 1 408
2 27498 1 408
2 27499 1 408
2 27500 1 408
2 27501 1 408
2 27502 1 409
2 27503 1 409
2 27504 1 409
2 27505 1 409
2 27506 1 409
2 27507 1 409
2 27508 1 409
2 27509 1 409
2 27510 1 409
2 27511 1 409
2 27512 1 410
2 27513 1 410
2 27514 1 410
2 27515 1 410
2 27516 1 412
2 27517 1 412
2 27518 1 412
2 27519 1 412
2 27520 1 412
2 27521 1 412
2 27522 1 412
2 27523 1 412
2 27524 1 412
2 27525 1 412
2 27526 1 412
2 27527 1 414
2 27528 1 414
2 27529 1 414
2 27530 1 417
2 27531 1 417
2 27532 1 417
2 27533 1 417
2 27534 1 417
2 27535 1 417
2 27536 1 417
2 27537 1 417
2 27538 1 417
2 27539 1 417
2 27540 1 417
2 27541 1 417
2 27542 1 420
2 27543 1 420
2 27544 1 420
2 27545 1 420
2 27546 1 420
2 27547 1 420
2 27548 1 420
2 27549 1 420
2 27550 1 420
2 27551 1 420
2 27552 1 420
2 27553 1 420
2 27554 1 422
2 27555 1 422
2 27556 1 423
2 27557 1 423
2 27558 1 424
2 27559 1 424
2 27560 1 436
2 27561 1 436
2 27562 1 436
2 27563 1 437
2 27564 1 437
2 27565 1 438
2 27566 1 438
2 27567 1 438
2 27568 1 439
2 27569 1 439
2 27570 1 439
2 27571 1 439
2 27572 1 439
2 27573 1 439
2 27574 1 439
2 27575 1 439
2 27576 1 439
2 27577 1 439
2 27578 1 439
2 27579 1 439
2 27580 1 439
2 27581 1 439
2 27582 1 439
2 27583 1 439
2 27584 1 439
2 27585 1 439
2 27586 1 439
2 27587 1 439
2 27588 1 439
2 27589 1 439
2 27590 1 439
2 27591 1 439
2 27592 1 439
2 27593 1 439
2 27594 1 440
2 27595 1 440
2 27596 1 440
2 27597 1 441
2 27598 1 441
2 27599 1 441
2 27600 1 441
2 27601 1 441
2 27602 1 441
2 27603 1 441
2 27604 1 441
2 27605 1 441
2 27606 1 441
2 27607 1 441
2 27608 1 441
2 27609 1 441
2 27610 1 441
2 27611 1 441
2 27612 1 441
2 27613 1 441
2 27614 1 441
2 27615 1 441
2 27616 1 441
2 27617 1 442
2 27618 1 442
2 27619 1 442
2 27620 1 442
2 27621 1 442
2 27622 1 442
2 27623 1 442
2 27624 1 442
2 27625 1 443
2 27626 1 443
2 27627 1 443
2 27628 1 444
2 27629 1 444
2 27630 1 451
2 27631 1 451
2 27632 1 451
2 27633 1 453
2 27634 1 453
2 27635 1 453
2 27636 1 453
2 27637 1 453
2 27638 1 453
2 27639 1 453
2 27640 1 461
2 27641 1 461
2 27642 1 462
2 27643 1 462
2 27644 1 462
2 27645 1 462
2 27646 1 462
2 27647 1 462
2 27648 1 462
2 27649 1 462
2 27650 1 462
2 27651 1 462
2 27652 1 464
2 27653 1 464
2 27654 1 464
2 27655 1 464
2 27656 1 464
2 27657 1 473
2 27658 1 473
2 27659 1 473
2 27660 1 473
2 27661 1 473
2 27662 1 473
2 27663 1 473
2 27664 1 473
2 27665 1 474
2 27666 1 474
2 27667 1 475
2 27668 1 475
2 27669 1 475
2 27670 1 475
2 27671 1 475
2 27672 1 475
2 27673 1 475
2 27674 1 475
2 27675 1 477
2 27676 1 477
2 27677 1 485
2 27678 1 485
2 27679 1 485
2 27680 1 485
2 27681 1 487
2 27682 1 487
2 27683 1 488
2 27684 1 488
2 27685 1 489
2 27686 1 489
2 27687 1 502
2 27688 1 502
2 27689 1 502
2 27690 1 503
2 27691 1 503
2 27692 1 503
2 27693 1 508
2 27694 1 508
2 27695 1 510
2 27696 1 510
2 27697 1 510
2 27698 1 510
2 27699 1 510
2 27700 1 510
2 27701 1 510
2 27702 1 510
2 27703 1 510
2 27704 1 510
2 27705 1 511
2 27706 1 511
2 27707 1 511
2 27708 1 512
2 27709 1 512
2 27710 1 518
2 27711 1 518
2 27712 1 519
2 27713 1 519
2 27714 1 527
2 27715 1 527
2 27716 1 527
2 27717 1 527
2 27718 1 527
2 27719 1 527
2 27720 1 527
2 27721 1 527
2 27722 1 527
2 27723 1 527
2 27724 1 527
2 27725 1 527
2 27726 1 527
2 27727 1 527
2 27728 1 528
2 27729 1 528
2 27730 1 529
2 27731 1 529
2 27732 1 529
2 27733 1 529
2 27734 1 529
2 27735 1 529
2 27736 1 529
2 27737 1 529
2 27738 1 531
2 27739 1 531
2 27740 1 531
2 27741 1 535
2 27742 1 535
2 27743 1 535
2 27744 1 535
2 27745 1 535
2 27746 1 535
2 27747 1 536
2 27748 1 536
2 27749 1 536
2 27750 1 544
2 27751 1 544
2 27752 1 544
2 27753 1 544
2 27754 1 544
2 27755 1 544
2 27756 1 544
2 27757 1 544
2 27758 1 544
2 27759 1 544
2 27760 1 546
2 27761 1 546
2 27762 1 554
2 27763 1 554
2 27764 1 554
2 27765 1 554
2 27766 1 554
2 27767 1 554
2 27768 1 555
2 27769 1 555
2 27770 1 555
2 27771 1 555
2 27772 1 555
2 27773 1 555
2 27774 1 556
2 27775 1 556
2 27776 1 561
2 27777 1 561
2 27778 1 561
2 27779 1 563
2 27780 1 563
2 27781 1 570
2 27782 1 570
2 27783 1 570
2 27784 1 570
2 27785 1 570
2 27786 1 570
2 27787 1 570
2 27788 1 570
2 27789 1 570
2 27790 1 571
2 27791 1 571
2 27792 1 571
2 27793 1 579
2 27794 1 579
2 27795 1 579
2 27796 1 579
2 27797 1 579
2 27798 1 579
2 27799 1 579
2 27800 1 579
2 27801 1 579
2 27802 1 579
2 27803 1 579
2 27804 1 579
2 27805 1 579
2 27806 1 579
2 27807 1 579
2 27808 1 579
2 27809 1 579
2 27810 1 579
2 27811 1 579
2 27812 1 579
2 27813 1 579
2 27814 1 579
2 27815 1 579
2 27816 1 580
2 27817 1 580
2 27818 1 580
2 27819 1 580
2 27820 1 584
2 27821 1 584
2 27822 1 584
2 27823 1 586
2 27824 1 586
2 27825 1 587
2 27826 1 587
2 27827 1 587
2 27828 1 587
2 27829 1 587
2 27830 1 587
2 27831 1 587
2 27832 1 587
2 27833 1 588
2 27834 1 588
2 27835 1 588
2 27836 1 592
2 27837 1 592
2 27838 1 593
2 27839 1 593
2 27840 1 593
2 27841 1 593
2 27842 1 593
2 27843 1 593
2 27844 1 593
2 27845 1 593
2 27846 1 593
2 27847 1 593
2 27848 1 593
2 27849 1 593
2 27850 1 593
2 27851 1 593
2 27852 1 593
2 27853 1 593
2 27854 1 593
2 27855 1 595
2 27856 1 595
2 27857 1 595
2 27858 1 596
2 27859 1 596
2 27860 1 603
2 27861 1 603
2 27862 1 603
2 27863 1 603
2 27864 1 603
2 27865 1 603
2 27866 1 603
2 27867 1 604
2 27868 1 604
2 27869 1 604
2 27870 1 604
2 27871 1 604
2 27872 1 604
2 27873 1 604
2 27874 1 604
2 27875 1 604
2 27876 1 604
2 27877 1 604
2 27878 1 604
2 27879 1 608
2 27880 1 608
2 27881 1 613
2 27882 1 613
2 27883 1 613
2 27884 1 613
2 27885 1 613
2 27886 1 613
2 27887 1 614
2 27888 1 614
2 27889 1 615
2 27890 1 615
2 27891 1 615
2 27892 1 617
2 27893 1 617
2 27894 1 617
2 27895 1 617
2 27896 1 617
2 27897 1 617
2 27898 1 617
2 27899 1 617
2 27900 1 619
2 27901 1 619
2 27902 1 622
2 27903 1 622
2 27904 1 627
2 27905 1 627
2 27906 1 627
2 27907 1 627
2 27908 1 627
2 27909 1 627
2 27910 1 627
2 27911 1 627
2 27912 1 627
2 27913 1 627
2 27914 1 627
2 27915 1 629
2 27916 1 629
2 27917 1 629
2 27918 1 629
2 27919 1 629
2 27920 1 629
2 27921 1 629
2 27922 1 629
2 27923 1 629
2 27924 1 629
2 27925 1 629
2 27926 1 629
2 27927 1 631
2 27928 1 631
2 27929 1 631
2 27930 1 631
2 27931 1 631
2 27932 1 631
2 27933 1 631
2 27934 1 632
2 27935 1 632
2 27936 1 632
2 27937 1 632
2 27938 1 632
2 27939 1 632
2 27940 1 632
2 27941 1 632
2 27942 1 632
2 27943 1 632
2 27944 1 632
2 27945 1 632
2 27946 1 632
2 27947 1 632
2 27948 1 632
2 27949 1 632
2 27950 1 632
2 27951 1 632
2 27952 1 632
2 27953 1 632
2 27954 1 632
2 27955 1 632
2 27956 1 632
2 27957 1 632
2 27958 1 632
2 27959 1 632
2 27960 1 632
2 27961 1 632
2 27962 1 632
2 27963 1 632
2 27964 1 632
2 27965 1 632
2 27966 1 632
2 27967 1 632
2 27968 1 632
2 27969 1 632
2 27970 1 632
2 27971 1 632
2 27972 1 632
2 27973 1 632
2 27974 1 632
2 27975 1 632
2 27976 1 632
2 27977 1 632
2 27978 1 632
2 27979 1 632
2 27980 1 632
2 27981 1 632
2 27982 1 632
2 27983 1 632
2 27984 1 632
2 27985 1 632
2 27986 1 632
2 27987 1 632
2 27988 1 632
2 27989 1 632
2 27990 1 632
2 27991 1 632
2 27992 1 632
2 27993 1 632
2 27994 1 632
2 27995 1 632
2 27996 1 632
2 27997 1 633
2 27998 1 633
2 27999 1 633
2 28000 1 633
2 28001 1 634
2 28002 1 634
2 28003 1 635
2 28004 1 635
2 28005 1 635
2 28006 1 636
2 28007 1 636
2 28008 1 638
2 28009 1 638
2 28010 1 638
2 28011 1 638
2 28012 1 638
2 28013 1 640
2 28014 1 640
2 28015 1 640
2 28016 1 640
2 28017 1 640
2 28018 1 640
2 28019 1 640
2 28020 1 640
2 28021 1 643
2 28022 1 643
2 28023 1 643
2 28024 1 643
2 28025 1 643
2 28026 1 643
2 28027 1 643
2 28028 1 646
2 28029 1 646
2 28030 1 646
2 28031 1 646
2 28032 1 646
2 28033 1 646
2 28034 1 646
2 28035 1 647
2 28036 1 647
2 28037 1 647
2 28038 1 647
2 28039 1 648
2 28040 1 648
2 28041 1 651
2 28042 1 651
2 28043 1 651
2 28044 1 651
2 28045 1 651
2 28046 1 651
2 28047 1 651
2 28048 1 651
2 28049 1 651
2 28050 1 654
2 28051 1 654
2 28052 1 654
2 28053 1 654
2 28054 1 654
2 28055 1 654
2 28056 1 654
2 28057 1 654
2 28058 1 654
2 28059 1 654
2 28060 1 654
2 28061 1 654
2 28062 1 655
2 28063 1 655
2 28064 1 655
2 28065 1 655
2 28066 1 655
2 28067 1 655
2 28068 1 656
2 28069 1 656
2 28070 1 656
2 28071 1 656
2 28072 1 656
2 28073 1 656
2 28074 1 656
2 28075 1 656
2 28076 1 656
2 28077 1 656
2 28078 1 656
2 28079 1 657
2 28080 1 657
2 28081 1 657
2 28082 1 664
2 28083 1 664
2 28084 1 664
2 28085 1 664
2 28086 1 664
2 28087 1 664
2 28088 1 664
2 28089 1 665
2 28090 1 665
2 28091 1 666
2 28092 1 666
2 28093 1 666
2 28094 1 666
2 28095 1 666
2 28096 1 666
2 28097 1 666
2 28098 1 666
2 28099 1 668
2 28100 1 668
2 28101 1 669
2 28102 1 669
2 28103 1 669
2 28104 1 669
2 28105 1 669
2 28106 1 669
2 28107 1 669
2 28108 1 669
2 28109 1 669
2 28110 1 669
2 28111 1 669
2 28112 1 669
2 28113 1 669
2 28114 1 669
2 28115 1 669
2 28116 1 669
2 28117 1 669
2 28118 1 669
2 28119 1 669
2 28120 1 669
2 28121 1 669
2 28122 1 669
2 28123 1 669
2 28124 1 669
2 28125 1 669
2 28126 1 669
2 28127 1 669
2 28128 1 669
2 28129 1 669
2 28130 1 669
2 28131 1 669
2 28132 1 669
2 28133 1 669
2 28134 1 669
2 28135 1 669
2 28136 1 669
2 28137 1 669
2 28138 1 669
2 28139 1 669
2 28140 1 669
2 28141 1 669
2 28142 1 669
2 28143 1 669
2 28144 1 669
2 28145 1 669
2 28146 1 669
2 28147 1 669
2 28148 1 669
2 28149 1 669
2 28150 1 669
2 28151 1 669
2 28152 1 669
2 28153 1 669
2 28154 1 669
2 28155 1 669
2 28156 1 669
2 28157 1 669
2 28158 1 669
2 28159 1 669
2 28160 1 669
2 28161 1 669
2 28162 1 669
2 28163 1 669
2 28164 1 669
2 28165 1 669
2 28166 1 669
2 28167 1 669
2 28168 1 669
2 28169 1 669
2 28170 1 669
2 28171 1 669
2 28172 1 669
2 28173 1 669
2 28174 1 669
2 28175 1 669
2 28176 1 669
2 28177 1 669
2 28178 1 670
2 28179 1 670
2 28180 1 670
2 28181 1 670
2 28182 1 670
2 28183 1 670
2 28184 1 670
2 28185 1 670
2 28186 1 670
2 28187 1 670
2 28188 1 670
2 28189 1 672
2 28190 1 672
2 28191 1 672
2 28192 1 672
2 28193 1 672
2 28194 1 672
2 28195 1 672
2 28196 1 672
2 28197 1 672
2 28198 1 672
2 28199 1 672
2 28200 1 672
2 28201 1 672
2 28202 1 672
2 28203 1 672
2 28204 1 672
2 28205 1 672
2 28206 1 672
2 28207 1 672
2 28208 1 672
2 28209 1 672
2 28210 1 672
2 28211 1 672
2 28212 1 672
2 28213 1 672
2 28214 1 672
2 28215 1 672
2 28216 1 672
2 28217 1 673
2 28218 1 673
2 28219 1 673
2 28220 1 673
2 28221 1 673
2 28222 1 673
2 28223 1 673
2 28224 1 681
2 28225 1 681
2 28226 1 681
2 28227 1 681
2 28228 1 681
2 28229 1 681
2 28230 1 681
2 28231 1 681
2 28232 1 681
2 28233 1 681
2 28234 1 681
2 28235 1 681
2 28236 1 681
2 28237 1 681
2 28238 1 681
2 28239 1 681
2 28240 1 681
2 28241 1 681
2 28242 1 681
2 28243 1 681
2 28244 1 681
2 28245 1 681
2 28246 1 681
2 28247 1 681
2 28248 1 681
2 28249 1 681
2 28250 1 682
2 28251 1 682
2 28252 1 682
2 28253 1 683
2 28254 1 683
2 28255 1 683
2 28256 1 683
2 28257 1 683
2 28258 1 683
2 28259 1 683
2 28260 1 683
2 28261 1 683
2 28262 1 683
2 28263 1 683
2 28264 1 683
2 28265 1 684
2 28266 1 684
2 28267 1 684
2 28268 1 685
2 28269 1 685
2 28270 1 685
2 28271 1 685
2 28272 1 685
2 28273 1 685
2 28274 1 685
2 28275 1 685
2 28276 1 685
2 28277 1 685
2 28278 1 685
2 28279 1 685
2 28280 1 687
2 28281 1 687
2 28282 1 688
2 28283 1 688
2 28284 1 688
2 28285 1 688
2 28286 1 688
2 28287 1 688
2 28288 1 688
2 28289 1 688
2 28290 1 688
2 28291 1 688
2 28292 1 691
2 28293 1 691
2 28294 1 691
2 28295 1 691
2 28296 1 691
2 28297 1 691
2 28298 1 691
2 28299 1 691
2 28300 1 691
2 28301 1 691
2 28302 1 691
2 28303 1 691
2 28304 1 691
2 28305 1 691
2 28306 1 691
2 28307 1 691
2 28308 1 691
2 28309 1 691
2 28310 1 691
2 28311 1 691
2 28312 1 691
2 28313 1 691
2 28314 1 691
2 28315 1 691
2 28316 1 691
2 28317 1 691
2 28318 1 691
2 28319 1 692
2 28320 1 692
2 28321 1 692
2 28322 1 692
2 28323 1 692
2 28324 1 693
2 28325 1 693
2 28326 1 693
2 28327 1 693
2 28328 1 693
2 28329 1 693
2 28330 1 695
2 28331 1 695
2 28332 1 698
2 28333 1 698
2 28334 1 701
2 28335 1 701
2 28336 1 701
2 28337 1 701
2 28338 1 701
2 28339 1 701
2 28340 1 701
2 28341 1 701
2 28342 1 701
2 28343 1 701
2 28344 1 701
2 28345 1 701
2 28346 1 701
2 28347 1 701
2 28348 1 701
2 28349 1 701
2 28350 1 701
2 28351 1 701
2 28352 1 701
2 28353 1 702
2 28354 1 702
2 28355 1 702
2 28356 1 702
2 28357 1 702
2 28358 1 702
2 28359 1 702
2 28360 1 702
2 28361 1 702
2 28362 1 702
2 28363 1 702
2 28364 1 702
2 28365 1 702
2 28366 1 704
2 28367 1 704
2 28368 1 704
2 28369 1 704
2 28370 1 705
2 28371 1 705
2 28372 1 708
2 28373 1 708
2 28374 1 708
2 28375 1 708
2 28376 1 708
2 28377 1 711
2 28378 1 711
2 28379 1 711
2 28380 1 721
2 28381 1 721
2 28382 1 721
2 28383 1 721
2 28384 1 721
2 28385 1 721
2 28386 1 721
2 28387 1 721
2 28388 1 721
2 28389 1 721
2 28390 1 721
2 28391 1 721
2 28392 1 721
2 28393 1 721
2 28394 1 721
2 28395 1 721
2 28396 1 725
2 28397 1 725
2 28398 1 725
2 28399 1 725
2 28400 1 725
2 28401 1 725
2 28402 1 726
2 28403 1 726
2 28404 1 726
2 28405 1 726
2 28406 1 727
2 28407 1 727
2 28408 1 727
2 28409 1 727
2 28410 1 728
2 28411 1 728
2 28412 1 730
2 28413 1 730
2 28414 1 731
2 28415 1 731
2 28416 1 731
2 28417 1 731
2 28418 1 731
2 28419 1 731
2 28420 1 731
2 28421 1 731
2 28422 1 731
2 28423 1 731
2 28424 1 731
2 28425 1 731
2 28426 1 731
2 28427 1 731
2 28428 1 731
2 28429 1 732
2 28430 1 732
2 28431 1 733
2 28432 1 733
2 28433 1 734
2 28434 1 734
2 28435 1 734
2 28436 1 734
2 28437 1 734
2 28438 1 734
2 28439 1 734
2 28440 1 734
2 28441 1 734
2 28442 1 734
2 28443 1 734
2 28444 1 734
2 28445 1 734
2 28446 1 734
2 28447 1 734
2 28448 1 734
2 28449 1 734
2 28450 1 734
2 28451 1 735
2 28452 1 735
2 28453 1 736
2 28454 1 736
2 28455 1 736
2 28456 1 736
2 28457 1 737
2 28458 1 737
2 28459 1 737
2 28460 1 737
2 28461 1 737
2 28462 1 737
2 28463 1 746
2 28464 1 746
2 28465 1 746
2 28466 1 746
2 28467 1 746
2 28468 1 746
2 28469 1 746
2 28470 1 748
2 28471 1 748
2 28472 1 748
2 28473 1 748
2 28474 1 750
2 28475 1 750
2 28476 1 750
2 28477 1 751
2 28478 1 751
2 28479 1 756
2 28480 1 756
2 28481 1 757
2 28482 1 757
2 28483 1 757
2 28484 1 764
2 28485 1 764
2 28486 1 764
2 28487 1 764
2 28488 1 764
2 28489 1 766
2 28490 1 766
2 28491 1 767
2 28492 1 767
2 28493 1 776
2 28494 1 776
2 28495 1 776
2 28496 1 776
2 28497 1 776
2 28498 1 776
2 28499 1 776
2 28500 1 776
2 28501 1 776
2 28502 1 776
2 28503 1 776
2 28504 1 776
2 28505 1 776
2 28506 1 776
2 28507 1 776
2 28508 1 776
2 28509 1 776
2 28510 1 776
2 28511 1 776
2 28512 1 776
2 28513 1 776
2 28514 1 776
2 28515 1 777
2 28516 1 777
2 28517 1 777
2 28518 1 777
2 28519 1 777
2 28520 1 777
2 28521 1 777
2 28522 1 777
2 28523 1 777
2 28524 1 777
2 28525 1 778
2 28526 1 778
2 28527 1 779
2 28528 1 779
2 28529 1 779
2 28530 1 779
2 28531 1 780
2 28532 1 780
2 28533 1 781
2 28534 1 781
2 28535 1 782
2 28536 1 782
2 28537 1 782
2 28538 1 783
2 28539 1 783
2 28540 1 784
2 28541 1 784
2 28542 1 784
2 28543 1 788
2 28544 1 788
2 28545 1 788
2 28546 1 788
2 28547 1 788
2 28548 1 788
2 28549 1 788
2 28550 1 788
2 28551 1 788
2 28552 1 788
2 28553 1 788
2 28554 1 788
2 28555 1 788
2 28556 1 788
2 28557 1 788
2 28558 1 790
2 28559 1 790
2 28560 1 790
2 28561 1 790
2 28562 1 790
2 28563 1 790
2 28564 1 790
2 28565 1 790
2 28566 1 790
2 28567 1 790
2 28568 1 792
2 28569 1 792
2 28570 1 792
2 28571 1 796
2 28572 1 796
2 28573 1 796
2 28574 1 796
2 28575 1 796
2 28576 1 796
2 28577 1 796
2 28578 1 797
2 28579 1 797
2 28580 1 798
2 28581 1 798
2 28582 1 806
2 28583 1 806
2 28584 1 806
2 28585 1 806
2 28586 1 806
2 28587 1 806
2 28588 1 806
2 28589 1 806
2 28590 1 806
2 28591 1 806
2 28592 1 806
2 28593 1 810
2 28594 1 810
2 28595 1 816
2 28596 1 816
2 28597 1 819
2 28598 1 819
2 28599 1 819
2 28600 1 819
2 28601 1 821
2 28602 1 821
2 28603 1 821
2 28604 1 821
2 28605 1 821
2 28606 1 821
2 28607 1 836
2 28608 1 836
2 28609 1 836
2 28610 1 837
2 28611 1 837
2 28612 1 839
2 28613 1 839
2 28614 1 840
2 28615 1 840
2 28616 1 844
2 28617 1 844
2 28618 1 844
2 28619 1 844
2 28620 1 846
2 28621 1 846
2 28622 1 848
2 28623 1 848
2 28624 1 848
2 28625 1 852
2 28626 1 852
2 28627 1 852
2 28628 1 853
2 28629 1 853
2 28630 1 854
2 28631 1 854
2 28632 1 854
2 28633 1 876
2 28634 1 876
2 28635 1 882
2 28636 1 882
2 28637 1 882
2 28638 1 882
2 28639 1 882
2 28640 1 882
2 28641 1 882
2 28642 1 882
2 28643 1 882
2 28644 1 882
2 28645 1 882
2 28646 1 882
2 28647 1 882
2 28648 1 882
2 28649 1 882
2 28650 1 882
2 28651 1 882
2 28652 1 882
2 28653 1 882
2 28654 1 882
2 28655 1 882
2 28656 1 882
2 28657 1 883
2 28658 1 883
2 28659 1 883
2 28660 1 883
2 28661 1 883
2 28662 1 884
2 28663 1 884
2 28664 1 891
2 28665 1 891
2 28666 1 891
2 28667 1 891
2 28668 1 891
2 28669 1 891
2 28670 1 891
2 28671 1 891
2 28672 1 891
2 28673 1 891
2 28674 1 891
2 28675 1 891
2 28676 1 891
2 28677 1 891
2 28678 1 891
2 28679 1 891
2 28680 1 891
2 28681 1 891
2 28682 1 891
2 28683 1 891
2 28684 1 892
2 28685 1 892
2 28686 1 902
2 28687 1 902
2 28688 1 902
2 28689 1 911
2 28690 1 911
2 28691 1 911
2 28692 1 911
2 28693 1 911
2 28694 1 915
2 28695 1 915
2 28696 1 922
2 28697 1 922
2 28698 1 922
2 28699 1 922
2 28700 1 922
2 28701 1 922
2 28702 1 922
2 28703 1 922
2 28704 1 922
2 28705 1 922
2 28706 1 922
2 28707 1 922
2 28708 1 922
2 28709 1 924
2 28710 1 924
2 28711 1 944
2 28712 1 944
2 28713 1 944
2 28714 1 944
2 28715 1 944
2 28716 1 944
2 28717 1 944
2 28718 1 949
2 28719 1 949
2 28720 1 949
2 28721 1 949
2 28722 1 949
2 28723 1 949
2 28724 1 949
2 28725 1 949
2 28726 1 949
2 28727 1 949
2 28728 1 949
2 28729 1 949
2 28730 1 949
2 28731 1 949
2 28732 1 949
2 28733 1 949
2 28734 1 949
2 28735 1 949
2 28736 1 949
2 28737 1 949
2 28738 1 949
2 28739 1 949
2 28740 1 949
2 28741 1 949
2 28742 1 949
2 28743 1 949
2 28744 1 950
2 28745 1 950
2 28746 1 950
2 28747 1 950
2 28748 1 950
2 28749 1 951
2 28750 1 951
2 28751 1 951
2 28752 1 955
2 28753 1 955
2 28754 1 955
2 28755 1 955
2 28756 1 955
2 28757 1 955
2 28758 1 955
2 28759 1 955
2 28760 1 955
2 28761 1 955
2 28762 1 955
2 28763 1 962
2 28764 1 962
2 28765 1 962
2 28766 1 962
2 28767 1 962
2 28768 1 962
2 28769 1 962
2 28770 1 962
2 28771 1 962
2 28772 1 962
2 28773 1 962
2 28774 1 962
2 28775 1 962
2 28776 1 963
2 28777 1 963
2 28778 1 963
2 28779 1 964
2 28780 1 964
2 28781 1 964
2 28782 1 972
2 28783 1 972
2 28784 1 972
2 28785 1 972
2 28786 1 972
2 28787 1 972
2 28788 1 972
2 28789 1 972
2 28790 1 972
2 28791 1 972
2 28792 1 972
2 28793 1 972
2 28794 1 973
2 28795 1 973
2 28796 1 973
2 28797 1 973
2 28798 1 973
2 28799 1 975
2 28800 1 975
2 28801 1 975
2 28802 1 975
2 28803 1 975
2 28804 1 975
2 28805 1 975
2 28806 1 975
2 28807 1 975
2 28808 1 975
2 28809 1 975
2 28810 1 975
2 28811 1 976
2 28812 1 976
2 28813 1 976
2 28814 1 976
2 28815 1 976
2 28816 1 976
2 28817 1 976
2 28818 1 980
2 28819 1 980
2 28820 1 980
2 28821 1 980
2 28822 1 980
2 28823 1 980
2 28824 1 980
2 28825 1 980
2 28826 1 980
2 28827 1 980
2 28828 1 980
2 28829 1 980
2 28830 1 983
2 28831 1 983
2 28832 1 983
2 28833 1 983
2 28834 1 983
2 28835 1 984
2 28836 1 984
2 28837 1 984
2 28838 1 988
2 28839 1 988
2 28840 1 988
2 28841 1 988
2 28842 1 988
2 28843 1 988
2 28844 1 989
2 28845 1 989
2 28846 1 989
2 28847 1 989
2 28848 1 989
2 28849 1 989
2 28850 1 989
2 28851 1 989
2 28852 1 989
2 28853 1 989
2 28854 1 989
2 28855 1 989
2 28856 1 989
2 28857 1 989
2 28858 1 989
2 28859 1 989
2 28860 1 989
2 28861 1 989
2 28862 1 989
2 28863 1 989
2 28864 1 989
2 28865 1 990
2 28866 1 990
2 28867 1 1005
2 28868 1 1005
2 28869 1 1005
2 28870 1 1005
2 28871 1 1005
2 28872 1 1005
2 28873 1 1005
2 28874 1 1005
2 28875 1 1005
2 28876 1 1005
2 28877 1 1005
2 28878 1 1005
2 28879 1 1005
2 28880 1 1009
2 28881 1 1009
2 28882 1 1012
2 28883 1 1012
2 28884 1 1012
2 28885 1 1012
2 28886 1 1012
2 28887 1 1016
2 28888 1 1016
2 28889 1 1017
2 28890 1 1017
2 28891 1 1017
2 28892 1 1017
2 28893 1 1025
2 28894 1 1025
2 28895 1 1025
2 28896 1 1025
2 28897 1 1025
2 28898 1 1026
2 28899 1 1026
2 28900 1 1028
2 28901 1 1028
2 28902 1 1032
2 28903 1 1032
2 28904 1 1035
2 28905 1 1035
2 28906 1 1038
2 28907 1 1038
2 28908 1 1041
2 28909 1 1041
2 28910 1 1041
2 28911 1 1041
2 28912 1 1043
2 28913 1 1043
2 28914 1 1054
2 28915 1 1054
2 28916 1 1055
2 28917 1 1055
2 28918 1 1062
2 28919 1 1062
2 28920 1 1062
2 28921 1 1062
2 28922 1 1063
2 28923 1 1063
2 28924 1 1063
2 28925 1 1072
2 28926 1 1072
2 28927 1 1072
2 28928 1 1079
2 28929 1 1079
2 28930 1 1079
2 28931 1 1094
2 28932 1 1094
2 28933 1 1094
2 28934 1 1094
2 28935 1 1094
2 28936 1 1094
2 28937 1 1094
2 28938 1 1094
2 28939 1 1094
2 28940 1 1094
2 28941 1 1094
2 28942 1 1094
2 28943 1 1094
2 28944 1 1094
2 28945 1 1094
2 28946 1 1094
2 28947 1 1094
2 28948 1 1094
2 28949 1 1094
2 28950 1 1094
2 28951 1 1094
2 28952 1 1094
2 28953 1 1094
2 28954 1 1094
2 28955 1 1095
2 28956 1 1095
2 28957 1 1095
2 28958 1 1095
2 28959 1 1095
2 28960 1 1095
2 28961 1 1095
2 28962 1 1095
2 28963 1 1108
2 28964 1 1108
2 28965 1 1108
2 28966 1 1108
2 28967 1 1108
2 28968 1 1108
2 28969 1 1108
2 28970 1 1111
2 28971 1 1111
2 28972 1 1111
2 28973 1 1111
2 28974 1 1111
2 28975 1 1111
2 28976 1 1111
2 28977 1 1111
2 28978 1 1111
2 28979 1 1111
2 28980 1 1111
2 28981 1 1111
2 28982 1 1111
2 28983 1 1111
2 28984 1 1111
2 28985 1 1111
2 28986 1 1111
2 28987 1 1111
2 28988 1 1111
2 28989 1 1111
2 28990 1 1111
2 28991 1 1111
2 28992 1 1111
2 28993 1 1111
2 28994 1 1111
2 28995 1 1111
2 28996 1 1111
2 28997 1 1111
2 28998 1 1111
2 28999 1 1111
2 29000 1 1111
2 29001 1 1111
2 29002 1 1111
2 29003 1 1111
2 29004 1 1111
2 29005 1 1111
2 29006 1 1111
2 29007 1 1111
2 29008 1 1111
2 29009 1 1111
2 29010 1 1111
2 29011 1 1111
2 29012 1 1111
2 29013 1 1111
2 29014 1 1111
2 29015 1 1111
2 29016 1 1111
2 29017 1 1111
2 29018 1 1111
2 29019 1 1111
2 29020 1 1111
2 29021 1 1111
2 29022 1 1112
2 29023 1 1112
2 29024 1 1112
2 29025 1 1112
2 29026 1 1112
2 29027 1 1113
2 29028 1 1113
2 29029 1 1113
2 29030 1 1115
2 29031 1 1115
2 29032 1 1115
2 29033 1 1115
2 29034 1 1115
2 29035 1 1115
2 29036 1 1115
2 29037 1 1115
2 29038 1 1115
2 29039 1 1115
2 29040 1 1117
2 29041 1 1117
2 29042 1 1117
2 29043 1 1117
2 29044 1 1117
2 29045 1 1117
2 29046 1 1117
2 29047 1 1123
2 29048 1 1123
2 29049 1 1123
2 29050 1 1123
2 29051 1 1123
2 29052 1 1123
2 29053 1 1123
2 29054 1 1123
2 29055 1 1123
2 29056 1 1123
2 29057 1 1123
2 29058 1 1123
2 29059 1 1123
2 29060 1 1123
2 29061 1 1123
2 29062 1 1123
2 29063 1 1123
2 29064 1 1123
2 29065 1 1124
2 29066 1 1124
2 29067 1 1124
2 29068 1 1124
2 29069 1 1124
2 29070 1 1124
2 29071 1 1124
2 29072 1 1124
2 29073 1 1128
2 29074 1 1128
2 29075 1 1128
2 29076 1 1128
2 29077 1 1128
2 29078 1 1131
2 29079 1 1131
2 29080 1 1131
2 29081 1 1131
2 29082 1 1131
2 29083 1 1131
2 29084 1 1131
2 29085 1 1134
2 29086 1 1134
2 29087 1 1134
2 29088 1 1142
2 29089 1 1142
2 29090 1 1142
2 29091 1 1142
2 29092 1 1143
2 29093 1 1143
2 29094 1 1143
2 29095 1 1143
2 29096 1 1143
2 29097 1 1143
2 29098 1 1143
2 29099 1 1143
2 29100 1 1143
2 29101 1 1143
2 29102 1 1143
2 29103 1 1143
2 29104 1 1143
2 29105 1 1143
2 29106 1 1143
2 29107 1 1143
2 29108 1 1143
2 29109 1 1143
2 29110 1 1143
2 29111 1 1143
2 29112 1 1143
2 29113 1 1143
2 29114 1 1143
2 29115 1 1143
2 29116 1 1143
2 29117 1 1143
2 29118 1 1143
2 29119 1 1143
2 29120 1 1143
2 29121 1 1143
2 29122 1 1143
2 29123 1 1144
2 29124 1 1144
2 29125 1 1146
2 29126 1 1146
2 29127 1 1146
2 29128 1 1146
2 29129 1 1146
2 29130 1 1170
2 29131 1 1170
2 29132 1 1170
2 29133 1 1173
2 29134 1 1173
2 29135 1 1174
2 29136 1 1174
2 29137 1 1174
2 29138 1 1174
2 29139 1 1174
2 29140 1 1178
2 29141 1 1178
2 29142 1 1178
2 29143 1 1178
2 29144 1 1178
2 29145 1 1178
2 29146 1 1178
2 29147 1 1178
2 29148 1 1178
2 29149 1 1178
2 29150 1 1178
2 29151 1 1178
2 29152 1 1178
2 29153 1 1178
2 29154 1 1178
2 29155 1 1178
2 29156 1 1178
2 29157 1 1178
2 29158 1 1178
2 29159 1 1178
2 29160 1 1178
2 29161 1 1178
2 29162 1 1178
2 29163 1 1178
2 29164 1 1178
2 29165 1 1178
2 29166 1 1178
2 29167 1 1178
2 29168 1 1178
2 29169 1 1178
2 29170 1 1178
2 29171 1 1178
2 29172 1 1178
2 29173 1 1178
2 29174 1 1178
2 29175 1 1178
2 29176 1 1179
2 29177 1 1179
2 29178 1 1179
2 29179 1 1179
2 29180 1 1179
2 29181 1 1179
2 29182 1 1179
2 29183 1 1179
2 29184 1 1179
2 29185 1 1179
2 29186 1 1179
2 29187 1 1179
2 29188 1 1179
2 29189 1 1179
2 29190 1 1179
2 29191 1 1179
2 29192 1 1179
2 29193 1 1179
2 29194 1 1181
2 29195 1 1181
2 29196 1 1182
2 29197 1 1182
2 29198 1 1182
2 29199 1 1182
2 29200 1 1182
2 29201 1 1192
2 29202 1 1192
2 29203 1 1192
2 29204 1 1192
2 29205 1 1192
2 29206 1 1194
2 29207 1 1194
2 29208 1 1194
2 29209 1 1194
2 29210 1 1194
2 29211 1 1194
2 29212 1 1194
2 29213 1 1194
2 29214 1 1195
2 29215 1 1195
2 29216 1 1195
2 29217 1 1198
2 29218 1 1198
2 29219 1 1198
2 29220 1 1198
2 29221 1 1198
2 29222 1 1198
2 29223 1 1198
2 29224 1 1198
2 29225 1 1198
2 29226 1 1198
2 29227 1 1198
2 29228 1 1198
2 29229 1 1198
2 29230 1 1198
2 29231 1 1198
2 29232 1 1198
2 29233 1 1198
2 29234 1 1199
2 29235 1 1199
2 29236 1 1199
2 29237 1 1201
2 29238 1 1201
2 29239 1 1201
2 29240 1 1201
2 29241 1 1201
2 29242 1 1201
2 29243 1 1201
2 29244 1 1204
2 29245 1 1204
2 29246 1 1204
2 29247 1 1204
2 29248 1 1204
2 29249 1 1204
2 29250 1 1204
2 29251 1 1204
2 29252 1 1204
2 29253 1 1204
2 29254 1 1204
2 29255 1 1204
2 29256 1 1204
2 29257 1 1204
2 29258 1 1204
2 29259 1 1204
2 29260 1 1204
2 29261 1 1204
2 29262 1 1204
2 29263 1 1204
2 29264 1 1204
2 29265 1 1204
2 29266 1 1204
2 29267 1 1204
2 29268 1 1204
2 29269 1 1205
2 29270 1 1205
2 29271 1 1205
2 29272 1 1205
2 29273 1 1205
2 29274 1 1205
2 29275 1 1205
2 29276 1 1205
2 29277 1 1205
2 29278 1 1205
2 29279 1 1205
2 29280 1 1205
2 29281 1 1205
2 29282 1 1205
2 29283 1 1205
2 29284 1 1205
2 29285 1 1205
2 29286 1 1205
2 29287 1 1206
2 29288 1 1206
2 29289 1 1206
2 29290 1 1206
2 29291 1 1207
2 29292 1 1207
2 29293 1 1208
2 29294 1 1208
2 29295 1 1210
2 29296 1 1210
2 29297 1 1210
2 29298 1 1219
2 29299 1 1219
2 29300 1 1219
2 29301 1 1219
2 29302 1 1219
2 29303 1 1219
2 29304 1 1219
2 29305 1 1219
2 29306 1 1219
2 29307 1 1220
2 29308 1 1220
2 29309 1 1220
2 29310 1 1220
2 29311 1 1221
2 29312 1 1221
2 29313 1 1221
2 29314 1 1221
2 29315 1 1226
2 29316 1 1226
2 29317 1 1226
2 29318 1 1226
2 29319 1 1226
2 29320 1 1227
2 29321 1 1227
2 29322 1 1227
2 29323 1 1227
2 29324 1 1230
2 29325 1 1230
2 29326 1 1230
2 29327 1 1230
2 29328 1 1230
2 29329 1 1230
2 29330 1 1231
2 29331 1 1231
2 29332 1 1243
2 29333 1 1243
2 29334 1 1251
2 29335 1 1251
2 29336 1 1251
2 29337 1 1251
2 29338 1 1251
2 29339 1 1251
2 29340 1 1252
2 29341 1 1252
2 29342 1 1252
2 29343 1 1252
2 29344 1 1252
2 29345 1 1252
2 29346 1 1253
2 29347 1 1253
2 29348 1 1253
2 29349 1 1256
2 29350 1 1256
2 29351 1 1259
2 29352 1 1259
2 29353 1 1259
2 29354 1 1259
2 29355 1 1260
2 29356 1 1260
2 29357 1 1273
2 29358 1 1273
2 29359 1 1284
2 29360 1 1284
2 29361 1 1284
2 29362 1 1284
2 29363 1 1284
2 29364 1 1284
2 29365 1 1284
2 29366 1 1284
2 29367 1 1284
2 29368 1 1284
2 29369 1 1285
2 29370 1 1285
2 29371 1 1285
2 29372 1 1285
2 29373 1 1285
2 29374 1 1285
2 29375 1 1285
2 29376 1 1285
2 29377 1 1286
2 29378 1 1286
2 29379 1 1287
2 29380 1 1287
2 29381 1 1287
2 29382 1 1295
2 29383 1 1295
2 29384 1 1295
2 29385 1 1295
2 29386 1 1295
2 29387 1 1295
2 29388 1 1295
2 29389 1 1295
2 29390 1 1297
2 29391 1 1297
2 29392 1 1298
2 29393 1 1298
2 29394 1 1298
2 29395 1 1298
2 29396 1 1298
2 29397 1 1298
2 29398 1 1298
2 29399 1 1298
2 29400 1 1298
2 29401 1 1298
2 29402 1 1298
2 29403 1 1298
2 29404 1 1298
2 29405 1 1299
2 29406 1 1299
2 29407 1 1301
2 29408 1 1301
2 29409 1 1301
2 29410 1 1301
2 29411 1 1301
2 29412 1 1301
2 29413 1 1301
2 29414 1 1301
2 29415 1 1301
2 29416 1 1301
2 29417 1 1301
2 29418 1 1301
2 29419 1 1301
2 29420 1 1301
2 29421 1 1301
2 29422 1 1301
2 29423 1 1301
2 29424 1 1301
2 29425 1 1301
2 29426 1 1302
2 29427 1 1302
2 29428 1 1302
2 29429 1 1303
2 29430 1 1303
2 29431 1 1305
2 29432 1 1305
2 29433 1 1311
2 29434 1 1311
2 29435 1 1314
2 29436 1 1314
2 29437 1 1314
2 29438 1 1314
2 29439 1 1314
2 29440 1 1314
2 29441 1 1314
2 29442 1 1315
2 29443 1 1315
2 29444 1 1315
2 29445 1 1316
2 29446 1 1316
2 29447 1 1320
2 29448 1 1320
2 29449 1 1320
2 29450 1 1320
2 29451 1 1321
2 29452 1 1321
2 29453 1 1321
2 29454 1 1322
2 29455 1 1322
2 29456 1 1322
2 29457 1 1335
2 29458 1 1335
2 29459 1 1335
2 29460 1 1335
2 29461 1 1335
2 29462 1 1336
2 29463 1 1336
2 29464 1 1336
2 29465 1 1336
2 29466 1 1337
2 29467 1 1337
2 29468 1 1340
2 29469 1 1340
2 29470 1 1340
2 29471 1 1343
2 29472 1 1343
2 29473 1 1343
2 29474 1 1343
2 29475 1 1343
2 29476 1 1343
2 29477 1 1343
2 29478 1 1343
2 29479 1 1343
2 29480 1 1343
2 29481 1 1343
2 29482 1 1343
2 29483 1 1343
2 29484 1 1343
2 29485 1 1343
2 29486 1 1343
2 29487 1 1343
2 29488 1 1343
2 29489 1 1343
2 29490 1 1343
2 29491 1 1343
2 29492 1 1343
2 29493 1 1343
2 29494 1 1343
2 29495 1 1343
2 29496 1 1343
2 29497 1 1343
2 29498 1 1343
2 29499 1 1343
2 29500 1 1344
2 29501 1 1344
2 29502 1 1350
2 29503 1 1350
2 29504 1 1357
2 29505 1 1357
2 29506 1 1357
2 29507 1 1357
2 29508 1 1358
2 29509 1 1358
2 29510 1 1364
2 29511 1 1364
2 29512 1 1364
2 29513 1 1364
2 29514 1 1364
2 29515 1 1364
2 29516 1 1364
2 29517 1 1364
2 29518 1 1364
2 29519 1 1364
2 29520 1 1364
2 29521 1 1364
2 29522 1 1365
2 29523 1 1365
2 29524 1 1365
2 29525 1 1365
2 29526 1 1365
2 29527 1 1365
2 29528 1 1366
2 29529 1 1366
2 29530 1 1368
2 29531 1 1368
2 29532 1 1368
2 29533 1 1368
2 29534 1 1368
2 29535 1 1372
2 29536 1 1372
2 29537 1 1372
2 29538 1 1372
2 29539 1 1372
2 29540 1 1372
2 29541 1 1373
2 29542 1 1373
2 29543 1 1374
2 29544 1 1374
2 29545 1 1374
2 29546 1 1374
2 29547 1 1374
2 29548 1 1374
2 29549 1 1374
2 29550 1 1374
2 29551 1 1374
2 29552 1 1375
2 29553 1 1375
2 29554 1 1375
2 29555 1 1375
2 29556 1 1375
2 29557 1 1375
2 29558 1 1375
2 29559 1 1375
2 29560 1 1375
2 29561 1 1376
2 29562 1 1376
2 29563 1 1376
2 29564 1 1376
2 29565 1 1376
2 29566 1 1377
2 29567 1 1377
2 29568 1 1380
2 29569 1 1380
2 29570 1 1380
2 29571 1 1380
2 29572 1 1383
2 29573 1 1383
2 29574 1 1383
2 29575 1 1383
2 29576 1 1383
2 29577 1 1383
2 29578 1 1383
2 29579 1 1384
2 29580 1 1384
2 29581 1 1384
2 29582 1 1386
2 29583 1 1386
2 29584 1 1386
2 29585 1 1386
2 29586 1 1386
2 29587 1 1386
2 29588 1 1386
2 29589 1 1386
2 29590 1 1386
2 29591 1 1386
2 29592 1 1387
2 29593 1 1387
2 29594 1 1387
2 29595 1 1387
2 29596 1 1387
2 29597 1 1387
2 29598 1 1387
2 29599 1 1387
2 29600 1 1387
2 29601 1 1387
2 29602 1 1387
2 29603 1 1387
2 29604 1 1387
2 29605 1 1387
2 29606 1 1387
2 29607 1 1387
2 29608 1 1387
2 29609 1 1389
2 29610 1 1389
2 29611 1 1393
2 29612 1 1393
2 29613 1 1393
2 29614 1 1393
2 29615 1 1393
2 29616 1 1393
2 29617 1 1393
2 29618 1 1393
2 29619 1 1393
2 29620 1 1393
2 29621 1 1393
2 29622 1 1393
2 29623 1 1393
2 29624 1 1393
2 29625 1 1393
2 29626 1 1393
2 29627 1 1393
2 29628 1 1393
2 29629 1 1395
2 29630 1 1395
2 29631 1 1395
2 29632 1 1395
2 29633 1 1399
2 29634 1 1399
2 29635 1 1399
2 29636 1 1399
2 29637 1 1399
2 29638 1 1399
2 29639 1 1400
2 29640 1 1400
2 29641 1 1400
2 29642 1 1400
2 29643 1 1400
2 29644 1 1402
2 29645 1 1402
2 29646 1 1402
2 29647 1 1421
2 29648 1 1421
2 29649 1 1421
2 29650 1 1421
2 29651 1 1423
2 29652 1 1423
2 29653 1 1423
2 29654 1 1423
2 29655 1 1424
2 29656 1 1424
2 29657 1 1426
2 29658 1 1426
2 29659 1 1426
2 29660 1 1426
2 29661 1 1426
2 29662 1 1426
2 29663 1 1426
2 29664 1 1426
2 29665 1 1426
2 29666 1 1426
2 29667 1 1427
2 29668 1 1427
2 29669 1 1427
2 29670 1 1427
2 29671 1 1427
2 29672 1 1427
2 29673 1 1427
2 29674 1 1427
2 29675 1 1428
2 29676 1 1428
2 29677 1 1429
2 29678 1 1429
2 29679 1 1429
2 29680 1 1429
2 29681 1 1432
2 29682 1 1432
2 29683 1 1435
2 29684 1 1435
2 29685 1 1435
2 29686 1 1435
2 29687 1 1435
2 29688 1 1435
2 29689 1 1435
2 29690 1 1435
2 29691 1 1435
2 29692 1 1435
2 29693 1 1435
2 29694 1 1435
2 29695 1 1437
2 29696 1 1437
2 29697 1 1437
2 29698 1 1437
2 29699 1 1437
2 29700 1 1437
2 29701 1 1437
2 29702 1 1437
2 29703 1 1445
2 29704 1 1445
2 29705 1 1448
2 29706 1 1448
2 29707 1 1448
2 29708 1 1448
2 29709 1 1448
2 29710 1 1455
2 29711 1 1455
2 29712 1 1456
2 29713 1 1456
2 29714 1 1456
2 29715 1 1456
2 29716 1 1457
2 29717 1 1457
2 29718 1 1464
2 29719 1 1464
2 29720 1 1480
2 29721 1 1480
2 29722 1 1480
2 29723 1 1480
2 29724 1 1480
2 29725 1 1488
2 29726 1 1488
2 29727 1 1488
2 29728 1 1488
2 29729 1 1488
2 29730 1 1489
2 29731 1 1489
2 29732 1 1489
2 29733 1 1490
2 29734 1 1490
2 29735 1 1490
2 29736 1 1504
2 29737 1 1504
2 29738 1 1504
2 29739 1 1504
2 29740 1 1505
2 29741 1 1505
2 29742 1 1508
2 29743 1 1508
2 29744 1 1509
2 29745 1 1509
2 29746 1 1509
2 29747 1 1509
2 29748 1 1510
2 29749 1 1510
2 29750 1 1519
2 29751 1 1519
2 29752 1 1519
2 29753 1 1519
2 29754 1 1519
2 29755 1 1519
2 29756 1 1519
2 29757 1 1519
2 29758 1 1519
2 29759 1 1519
2 29760 1 1519
2 29761 1 1519
2 29762 1 1519
2 29763 1 1519
2 29764 1 1519
2 29765 1 1519
2 29766 1 1519
2 29767 1 1519
2 29768 1 1519
2 29769 1 1519
2 29770 1 1519
2 29771 1 1520
2 29772 1 1520
2 29773 1 1520
2 29774 1 1520
2 29775 1 1520
2 29776 1 1520
2 29777 1 1520
2 29778 1 1523
2 29779 1 1523
2 29780 1 1523
2 29781 1 1523
2 29782 1 1523
2 29783 1 1523
2 29784 1 1523
2 29785 1 1523
2 29786 1 1523
2 29787 1 1523
2 29788 1 1524
2 29789 1 1524
2 29790 1 1526
2 29791 1 1526
2 29792 1 1527
2 29793 1 1527
2 29794 1 1528
2 29795 1 1528
2 29796 1 1536
2 29797 1 1536
2 29798 1 1537
2 29799 1 1537
2 29800 1 1537
2 29801 1 1540
2 29802 1 1540
2 29803 1 1540
2 29804 1 1541
2 29805 1 1541
2 29806 1 1541
2 29807 1 1541
2 29808 1 1541
2 29809 1 1550
2 29810 1 1550
2 29811 1 1550
2 29812 1 1550
2 29813 1 1550
2 29814 1 1550
2 29815 1 1550
2 29816 1 1550
2 29817 1 1550
2 29818 1 1552
2 29819 1 1552
2 29820 1 1552
2 29821 1 1552
2 29822 1 1552
2 29823 1 1552
2 29824 1 1552
2 29825 1 1552
2 29826 1 1552
2 29827 1 1552
2 29828 1 1552
2 29829 1 1552
2 29830 1 1552
2 29831 1 1552
2 29832 1 1552
2 29833 1 1552
2 29834 1 1552
2 29835 1 1552
2 29836 1 1552
2 29837 1 1552
2 29838 1 1553
2 29839 1 1553
2 29840 1 1560
2 29841 1 1560
2 29842 1 1561
2 29843 1 1561
2 29844 1 1561
2 29845 1 1570
2 29846 1 1570
2 29847 1 1574
2 29848 1 1574
2 29849 1 1574
2 29850 1 1574
2 29851 1 1574
2 29852 1 1574
2 29853 1 1574
2 29854 1 1577
2 29855 1 1577
2 29856 1 1577
2 29857 1 1585
2 29858 1 1585
2 29859 1 1585
2 29860 1 1585
2 29861 1 1585
2 29862 1 1586
2 29863 1 1586
2 29864 1 1591
2 29865 1 1591
2 29866 1 1591
2 29867 1 1591
2 29868 1 1591
2 29869 1 1591
2 29870 1 1591
2 29871 1 1591
2 29872 1 1591
2 29873 1 1591
2 29874 1 1591
2 29875 1 1591
2 29876 1 1591
2 29877 1 1591
2 29878 1 1591
2 29879 1 1591
2 29880 1 1591
2 29881 1 1591
2 29882 1 1591
2 29883 1 1591
2 29884 1 1599
2 29885 1 1599
2 29886 1 1599
2 29887 1 1599
2 29888 1 1599
2 29889 1 1599
2 29890 1 1599
2 29891 1 1599
2 29892 1 1599
2 29893 1 1599
2 29894 1 1599
2 29895 1 1599
2 29896 1 1599
2 29897 1 1599
2 29898 1 1599
2 29899 1 1599
2 29900 1 1599
2 29901 1 1599
2 29902 1 1599
2 29903 1 1599
2 29904 1 1599
2 29905 1 1600
2 29906 1 1600
2 29907 1 1600
2 29908 1 1601
2 29909 1 1601
2 29910 1 1602
2 29911 1 1602
2 29912 1 1602
2 29913 1 1602
2 29914 1 1605
2 29915 1 1605
2 29916 1 1605
2 29917 1 1620
2 29918 1 1620
2 29919 1 1620
2 29920 1 1620
2 29921 1 1620
2 29922 1 1620
2 29923 1 1621
2 29924 1 1621
2 29925 1 1633
2 29926 1 1633
2 29927 1 1633
2 29928 1 1634
2 29929 1 1634
2 29930 1 1634
2 29931 1 1634
2 29932 1 1634
2 29933 1 1634
2 29934 1 1634
2 29935 1 1635
2 29936 1 1635
2 29937 1 1635
2 29938 1 1635
2 29939 1 1635
2 29940 1 1645
2 29941 1 1645
2 29942 1 1645
2 29943 1 1645
2 29944 1 1646
2 29945 1 1646
2 29946 1 1646
2 29947 1 1646
2 29948 1 1646
2 29949 1 1646
2 29950 1 1646
2 29951 1 1646
2 29952 1 1646
2 29953 1 1646
2 29954 1 1646
2 29955 1 1646
2 29956 1 1646
2 29957 1 1646
2 29958 1 1646
2 29959 1 1646
2 29960 1 1646
2 29961 1 1646
2 29962 1 1646
2 29963 1 1646
2 29964 1 1646
2 29965 1 1647
2 29966 1 1647
2 29967 1 1647
2 29968 1 1647
2 29969 1 1647
2 29970 1 1647
2 29971 1 1647
2 29972 1 1647
2 29973 1 1647
2 29974 1 1647
2 29975 1 1647
2 29976 1 1647
2 29977 1 1647
2 29978 1 1647
2 29979 1 1647
2 29980 1 1647
2 29981 1 1650
2 29982 1 1650
2 29983 1 1650
2 29984 1 1650
2 29985 1 1650
2 29986 1 1650
2 29987 1 1650
2 29988 1 1650
2 29989 1 1654
2 29990 1 1654
2 29991 1 1654
2 29992 1 1658
2 29993 1 1658
2 29994 1 1661
2 29995 1 1661
2 29996 1 1662
2 29997 1 1662
2 29998 1 1662
2 29999 1 1662
2 30000 1 1662
2 30001 1 1674
2 30002 1 1674
2 30003 1 1674
2 30004 1 1674
2 30005 1 1675
2 30006 1 1675
2 30007 1 1676
2 30008 1 1676
2 30009 1 1681
2 30010 1 1681
2 30011 1 1681
2 30012 1 1681
2 30013 1 1682
2 30014 1 1682
2 30015 1 1682
2 30016 1 1692
2 30017 1 1692
2 30018 1 1692
2 30019 1 1693
2 30020 1 1693
2 30021 1 1695
2 30022 1 1695
2 30023 1 1695
2 30024 1 1695
2 30025 1 1695
2 30026 1 1695
2 30027 1 1695
2 30028 1 1695
2 30029 1 1695
2 30030 1 1695
2 30031 1 1695
2 30032 1 1695
2 30033 1 1695
2 30034 1 1695
2 30035 1 1695
2 30036 1 1697
2 30037 1 1697
2 30038 1 1710
2 30039 1 1710
2 30040 1 1710
2 30041 1 1711
2 30042 1 1711
2 30043 1 1711
2 30044 1 1711
2 30045 1 1714
2 30046 1 1714
2 30047 1 1714
2 30048 1 1714
2 30049 1 1714
2 30050 1 1714
2 30051 1 1718
2 30052 1 1718
2 30053 1 1725
2 30054 1 1725
2 30055 1 1725
2 30056 1 1738
2 30057 1 1738
2 30058 1 1738
2 30059 1 1738
2 30060 1 1739
2 30061 1 1739
2 30062 1 1739
2 30063 1 1748
2 30064 1 1748
2 30065 1 1756
2 30066 1 1756
2 30067 1 1757
2 30068 1 1757
2 30069 1 1757
2 30070 1 1757
2 30071 1 1757
2 30072 1 1757
2 30073 1 1757
2 30074 1 1757
2 30075 1 1757
2 30076 1 1757
2 30077 1 1757
2 30078 1 1757
2 30079 1 1758
2 30080 1 1758
2 30081 1 1758
2 30082 1 1758
2 30083 1 1759
2 30084 1 1759
2 30085 1 1760
2 30086 1 1760
2 30087 1 1761
2 30088 1 1761
2 30089 1 1771
2 30090 1 1771
2 30091 1 1771
2 30092 1 1771
2 30093 1 1772
2 30094 1 1772
2 30095 1 1772
2 30096 1 1779
2 30097 1 1779
2 30098 1 1779
2 30099 1 1779
2 30100 1 1779
2 30101 1 1787
2 30102 1 1787
2 30103 1 1793
2 30104 1 1793
2 30105 1 1793
2 30106 1 1796
2 30107 1 1796
2 30108 1 1796
2 30109 1 1796
2 30110 1 1796
2 30111 1 1796
2 30112 1 1796
2 30113 1 1796
2 30114 1 1796
2 30115 1 1796
2 30116 1 1796
2 30117 1 1796
2 30118 1 1796
2 30119 1 1797
2 30120 1 1797
2 30121 1 1798
2 30122 1 1798
2 30123 1 1798
2 30124 1 1799
2 30125 1 1799
2 30126 1 1799
2 30127 1 1807
2 30128 1 1807
2 30129 1 1807
2 30130 1 1807
2 30131 1 1807
2 30132 1 1807
2 30133 1 1807
2 30134 1 1807
2 30135 1 1807
2 30136 1 1807
2 30137 1 1807
2 30138 1 1807
2 30139 1 1807
2 30140 1 1807
2 30141 1 1807
2 30142 1 1808
2 30143 1 1808
2 30144 1 1808
2 30145 1 1809
2 30146 1 1809
2 30147 1 1809
2 30148 1 1809
2 30149 1 1810
2 30150 1 1810
2 30151 1 1811
2 30152 1 1811
2 30153 1 1824
2 30154 1 1824
2 30155 1 1825
2 30156 1 1825
2 30157 1 1828
2 30158 1 1828
2 30159 1 1834
2 30160 1 1834
2 30161 1 1834
2 30162 1 1834
2 30163 1 1834
2 30164 1 1834
2 30165 1 1834
2 30166 1 1834
2 30167 1 1834
2 30168 1 1834
2 30169 1 1834
2 30170 1 1834
2 30171 1 1834
2 30172 1 1834
2 30173 1 1834
2 30174 1 1834
2 30175 1 1834
2 30176 1 1834
2 30177 1 1834
2 30178 1 1834
2 30179 1 1834
2 30180 1 1843
2 30181 1 1843
2 30182 1 1844
2 30183 1 1844
2 30184 1 1844
2 30185 1 1845
2 30186 1 1845
2 30187 1 1869
2 30188 1 1869
2 30189 1 1869
2 30190 1 1869
2 30191 1 1869
2 30192 1 1869
2 30193 1 1869
2 30194 1 1869
2 30195 1 1869
2 30196 1 1869
2 30197 1 1875
2 30198 1 1875
2 30199 1 1875
2 30200 1 1875
2 30201 1 1875
2 30202 1 1879
2 30203 1 1879
2 30204 1 1879
2 30205 1 1879
2 30206 1 1880
2 30207 1 1880
2 30208 1 1880
2 30209 1 1880
2 30210 1 1880
2 30211 1 1880
2 30212 1 1881
2 30213 1 1881
2 30214 1 1881
2 30215 1 1884
2 30216 1 1884
2 30217 1 1884
2 30218 1 1884
2 30219 1 1884
2 30220 1 1885
2 30221 1 1885
2 30222 1 1893
2 30223 1 1893
2 30224 1 1893
2 30225 1 1893
2 30226 1 1893
2 30227 1 1893
2 30228 1 1895
2 30229 1 1895
2 30230 1 1895
2 30231 1 1896
2 30232 1 1896
2 30233 1 1905
2 30234 1 1905
2 30235 1 1916
2 30236 1 1916
2 30237 1 1916
2 30238 1 1916
2 30239 1 1917
2 30240 1 1917
2 30241 1 1920
2 30242 1 1920
2 30243 1 1920
2 30244 1 1927
2 30245 1 1927
2 30246 1 1927
2 30247 1 1927
2 30248 1 1927
2 30249 1 1931
2 30250 1 1931
2 30251 1 1931
2 30252 1 1931
2 30253 1 1931
2 30254 1 1931
2 30255 1 1931
2 30256 1 1931
2 30257 1 1931
2 30258 1 1931
2 30259 1 1931
2 30260 1 1931
2 30261 1 1935
2 30262 1 1935
2 30263 1 1935
2 30264 1 1938
2 30265 1 1938
2 30266 1 1938
2 30267 1 1940
2 30268 1 1940
2 30269 1 1947
2 30270 1 1947
2 30271 1 1947
2 30272 1 1957
2 30273 1 1957
2 30274 1 1957
2 30275 1 1957
2 30276 1 1957
2 30277 1 1957
2 30278 1 1957
2 30279 1 1958
2 30280 1 1958
2 30281 1 1959
2 30282 1 1959
2 30283 1 1970
2 30284 1 1970
2 30285 1 1970
2 30286 1 1970
2 30287 1 1970
2 30288 1 1970
2 30289 1 1970
2 30290 1 1970
2 30291 1 1970
2 30292 1 1971
2 30293 1 1971
2 30294 1 1971
2 30295 1 1975
2 30296 1 1975
2 30297 1 1976
2 30298 1 1976
2 30299 1 1976
2 30300 1 1976
2 30301 1 1976
2 30302 1 1990
2 30303 1 1990
2 30304 1 1990
2 30305 1 1990
2 30306 1 1990
2 30307 1 1990
2 30308 1 1990
2 30309 1 1990
2 30310 1 1998
2 30311 1 1998
2 30312 1 1998
2 30313 1 1998
2 30314 1 1998
2 30315 1 1998
2 30316 1 1998
2 30317 1 1998
2 30318 1 1998
2 30319 1 1998
2 30320 1 1998
2 30321 1 1998
2 30322 1 1998
2 30323 1 1998
2 30324 1 1998
2 30325 1 1998
2 30326 1 1999
2 30327 1 1999
2 30328 1 1999
2 30329 1 1999
2 30330 1 1999
2 30331 1 1999
2 30332 1 1999
2 30333 1 1999
2 30334 1 1999
2 30335 1 1999
2 30336 1 1999
2 30337 1 1999
2 30338 1 1999
2 30339 1 1999
2 30340 1 1999
2 30341 1 1999
2 30342 1 1999
2 30343 1 1999
2 30344 1 1999
2 30345 1 1999
2 30346 1 2000
2 30347 1 2000
2 30348 1 2000
2 30349 1 2000
2 30350 1 2001
2 30351 1 2001
2 30352 1 2001
2 30353 1 2001
2 30354 1 2003
2 30355 1 2003
2 30356 1 2003
2 30357 1 2003
2 30358 1 2003
2 30359 1 2003
2 30360 1 2003
2 30361 1 2003
2 30362 1 2004
2 30363 1 2004
2 30364 1 2014
2 30365 1 2014
2 30366 1 2014
2 30367 1 2014
2 30368 1 2014
2 30369 1 2014
2 30370 1 2014
2 30371 1 2015
2 30372 1 2015
2 30373 1 2015
2 30374 1 2019
2 30375 1 2019
2 30376 1 2019
2 30377 1 2019
2 30378 1 2020
2 30379 1 2020
2 30380 1 2020
2 30381 1 2020
2 30382 1 2020
2 30383 1 2020
2 30384 1 2020
2 30385 1 2020
2 30386 1 2028
2 30387 1 2028
2 30388 1 2028
2 30389 1 2029
2 30390 1 2029
2 30391 1 2029
2 30392 1 2029
2 30393 1 2029
2 30394 1 2037
2 30395 1 2037
2 30396 1 2037
2 30397 1 2037
2 30398 1 2038
2 30399 1 2038
2 30400 1 2039
2 30401 1 2039
2 30402 1 2039
2 30403 1 2039
2 30404 1 2039
2 30405 1 2039
2 30406 1 2039
2 30407 1 2039
2 30408 1 2040
2 30409 1 2040
2 30410 1 2045
2 30411 1 2045
2 30412 1 2046
2 30413 1 2046
2 30414 1 2047
2 30415 1 2047
2 30416 1 2057
2 30417 1 2057
2 30418 1 2057
2 30419 1 2057
2 30420 1 2076
2 30421 1 2076
2 30422 1 2076
2 30423 1 2078
2 30424 1 2078
2 30425 1 2078
2 30426 1 2078
2 30427 1 2079
2 30428 1 2079
2 30429 1 2079
2 30430 1 2079
2 30431 1 2079
2 30432 1 2079
2 30433 1 2079
2 30434 1 2079
2 30435 1 2079
2 30436 1 2079
2 30437 1 2079
2 30438 1 2079
2 30439 1 2089
2 30440 1 2089
2 30441 1 2089
2 30442 1 2089
2 30443 1 2089
2 30444 1 2091
2 30445 1 2091
2 30446 1 2092
2 30447 1 2092
2 30448 1 2092
2 30449 1 2092
2 30450 1 2092
2 30451 1 2092
2 30452 1 2092
2 30453 1 2097
2 30454 1 2097
2 30455 1 2097
2 30456 1 2097
2 30457 1 2097
2 30458 1 2098
2 30459 1 2098
2 30460 1 2098
2 30461 1 2098
2 30462 1 2098
2 30463 1 2098
2 30464 1 2098
2 30465 1 2098
2 30466 1 2098
2 30467 1 2098
2 30468 1 2098
2 30469 1 2098
2 30470 1 2098
2 30471 1 2098
2 30472 1 2098
2 30473 1 2098
2 30474 1 2098
2 30475 1 2107
2 30476 1 2107
2 30477 1 2107
2 30478 1 2107
2 30479 1 2107
2 30480 1 2108
2 30481 1 2108
2 30482 1 2130
2 30483 1 2130
2 30484 1 2131
2 30485 1 2131
2 30486 1 2131
2 30487 1 2140
2 30488 1 2140
2 30489 1 2140
2 30490 1 2140
2 30491 1 2140
2 30492 1 2140
2 30493 1 2140
2 30494 1 2140
2 30495 1 2150
2 30496 1 2150
2 30497 1 2154
2 30498 1 2154
2 30499 1 2154
2 30500 1 2154
2 30501 1 2179
2 30502 1 2179
2 30503 1 2180
2 30504 1 2180
2 30505 1 2180
2 30506 1 2180
2 30507 1 2180
2 30508 1 2180
2 30509 1 2180
2 30510 1 2180
2 30511 1 2180
2 30512 1 2181
2 30513 1 2181
2 30514 1 2182
2 30515 1 2182
2 30516 1 2185
2 30517 1 2185
2 30518 1 2186
2 30519 1 2186
2 30520 1 2186
2 30521 1 2192
2 30522 1 2192
2 30523 1 2199
2 30524 1 2199
2 30525 1 2202
2 30526 1 2202
2 30527 1 2202
2 30528 1 2202
2 30529 1 2203
2 30530 1 2203
2 30531 1 2203
2 30532 1 2203
2 30533 1 2203
2 30534 1 2203
2 30535 1 2205
2 30536 1 2205
2 30537 1 2217
2 30538 1 2217
2 30539 1 2217
2 30540 1 2217
2 30541 1 2217
2 30542 1 2218
2 30543 1 2218
2 30544 1 2218
2 30545 1 2218
2 30546 1 2221
2 30547 1 2221
2 30548 1 2229
2 30549 1 2229
2 30550 1 2229
2 30551 1 2229
2 30552 1 2229
2 30553 1 2229
2 30554 1 2229
2 30555 1 2230
2 30556 1 2230
2 30557 1 2230
2 30558 1 2230
2 30559 1 2231
2 30560 1 2231
2 30561 1 2232
2 30562 1 2232
2 30563 1 2232
2 30564 1 2232
2 30565 1 2233
2 30566 1 2233
2 30567 1 2233
2 30568 1 2233
2 30569 1 2233
2 30570 1 2247
2 30571 1 2247
2 30572 1 2247
2 30573 1 2247
2 30574 1 2247
2 30575 1 2247
2 30576 1 2247
2 30577 1 2247
2 30578 1 2247
2 30579 1 2247
2 30580 1 2248
2 30581 1 2248
2 30582 1 2248
2 30583 1 2248
2 30584 1 2248
2 30585 1 2249
2 30586 1 2249
2 30587 1 2250
2 30588 1 2250
2 30589 1 2250
2 30590 1 2262
2 30591 1 2262
2 30592 1 2262
2 30593 1 2263
2 30594 1 2263
2 30595 1 2267
2 30596 1 2267
2 30597 1 2267
2 30598 1 2267
2 30599 1 2267
2 30600 1 2267
2 30601 1 2267
2 30602 1 2267
2 30603 1 2267
2 30604 1 2273
2 30605 1 2273
2 30606 1 2274
2 30607 1 2274
2 30608 1 2274
2 30609 1 2274
2 30610 1 2274
2 30611 1 2274
2 30612 1 2275
2 30613 1 2275
2 30614 1 2275
2 30615 1 2302
2 30616 1 2302
2 30617 1 2302
2 30618 1 2302
2 30619 1 2302
2 30620 1 2302
2 30621 1 2302
2 30622 1 2302
2 30623 1 2302
2 30624 1 2303
2 30625 1 2303
2 30626 1 2303
2 30627 1 2303
2 30628 1 2306
2 30629 1 2306
2 30630 1 2306
2 30631 1 2306
2 30632 1 2307
2 30633 1 2307
2 30634 1 2307
2 30635 1 2314
2 30636 1 2314
2 30637 1 2314
2 30638 1 2314
2 30639 1 2314
2 30640 1 2314
2 30641 1 2314
2 30642 1 2314
2 30643 1 2314
2 30644 1 2314
2 30645 1 2314
2 30646 1 2314
2 30647 1 2314
2 30648 1 2314
2 30649 1 2314
2 30650 1 2314
2 30651 1 2314
2 30652 1 2314
2 30653 1 2314
2 30654 1 2314
2 30655 1 2314
2 30656 1 2317
2 30657 1 2317
2 30658 1 2328
2 30659 1 2328
2 30660 1 2329
2 30661 1 2329
2 30662 1 2340
2 30663 1 2340
2 30664 1 2340
2 30665 1 2341
2 30666 1 2341
2 30667 1 2342
2 30668 1 2342
2 30669 1 2342
2 30670 1 2342
2 30671 1 2342
2 30672 1 2342
2 30673 1 2342
2 30674 1 2342
2 30675 1 2352
2 30676 1 2352
2 30677 1 2352
2 30678 1 2352
2 30679 1 2352
2 30680 1 2352
2 30681 1 2353
2 30682 1 2353
2 30683 1 2353
2 30684 1 2353
2 30685 1 2353
2 30686 1 2357
2 30687 1 2357
2 30688 1 2357
2 30689 1 2357
2 30690 1 2357
2 30691 1 2357
2 30692 1 2357
2 30693 1 2357
2 30694 1 2357
2 30695 1 2357
2 30696 1 2357
2 30697 1 2357
2 30698 1 2357
2 30699 1 2358
2 30700 1 2358
2 30701 1 2359
2 30702 1 2359
2 30703 1 2368
2 30704 1 2368
2 30705 1 2368
2 30706 1 2368
2 30707 1 2368
2 30708 1 2368
2 30709 1 2368
2 30710 1 2368
2 30711 1 2369
2 30712 1 2369
2 30713 1 2377
2 30714 1 2377
2 30715 1 2391
2 30716 1 2391
2 30717 1 2391
2 30718 1 2391
2 30719 1 2393
2 30720 1 2393
2 30721 1 2396
2 30722 1 2396
2 30723 1 2396
2 30724 1 2397
2 30725 1 2397
2 30726 1 2397
2 30727 1 2397
2 30728 1 2412
2 30729 1 2412
2 30730 1 2412
2 30731 1 2412
2 30732 1 2412
2 30733 1 2412
2 30734 1 2412
2 30735 1 2412
2 30736 1 2412
2 30737 1 2413
2 30738 1 2413
2 30739 1 2413
2 30740 1 2413
2 30741 1 2413
2 30742 1 2428
2 30743 1 2428
2 30744 1 2428
2 30745 1 2428
2 30746 1 2429
2 30747 1 2429
2 30748 1 2432
2 30749 1 2432
2 30750 1 2440
2 30751 1 2440
2 30752 1 2440
2 30753 1 2440
2 30754 1 2440
2 30755 1 2441
2 30756 1 2441
2 30757 1 2449
2 30758 1 2449
2 30759 1 2459
2 30760 1 2459
2 30761 1 2459
2 30762 1 2459
2 30763 1 2459
2 30764 1 2459
2 30765 1 2459
2 30766 1 2479
2 30767 1 2479
2 30768 1 2480
2 30769 1 2480
2 30770 1 2481
2 30771 1 2481
2 30772 1 2481
2 30773 1 2481
2 30774 1 2481
2 30775 1 2481
2 30776 1 2481
2 30777 1 2485
2 30778 1 2485
2 30779 1 2485
2 30780 1 2485
2 30781 1 2485
2 30782 1 2485
2 30783 1 2485
2 30784 1 2486
2 30785 1 2486
2 30786 1 2494
2 30787 1 2494
2 30788 1 2494
2 30789 1 2494
2 30790 1 2494
2 30791 1 2494
2 30792 1 2494
2 30793 1 2494
2 30794 1 2495
2 30795 1 2495
2 30796 1 2495
2 30797 1 2496
2 30798 1 2496
2 30799 1 2496
2 30800 1 2504
2 30801 1 2504
2 30802 1 2504
2 30803 1 2504
2 30804 1 2504
2 30805 1 2504
2 30806 1 2520
2 30807 1 2520
2 30808 1 2520
2 30809 1 2520
2 30810 1 2520
2 30811 1 2523
2 30812 1 2523
2 30813 1 2523
2 30814 1 2526
2 30815 1 2526
2 30816 1 2527
2 30817 1 2527
2 30818 1 2527
2 30819 1 2527
2 30820 1 2527
2 30821 1 2527
2 30822 1 2527
2 30823 1 2527
2 30824 1 2527
2 30825 1 2527
2 30826 1 2527
2 30827 1 2527
2 30828 1 2527
2 30829 1 2531
2 30830 1 2531
2 30831 1 2543
2 30832 1 2543
2 30833 1 2543
2 30834 1 2543
2 30835 1 2543
2 30836 1 2543
2 30837 1 2543
2 30838 1 2543
2 30839 1 2543
2 30840 1 2547
2 30841 1 2547
2 30842 1 2547
2 30843 1 2547
2 30844 1 2557
2 30845 1 2557
2 30846 1 2557
2 30847 1 2557
2 30848 1 2557
2 30849 1 2557
2 30850 1 2557
2 30851 1 2557
2 30852 1 2562
2 30853 1 2562
2 30854 1 2562
2 30855 1 2562
2 30856 1 2562
2 30857 1 2562
2 30858 1 2563
2 30859 1 2563
2 30860 1 2576
2 30861 1 2576
2 30862 1 2576
2 30863 1 2580
2 30864 1 2580
2 30865 1 2583
2 30866 1 2583
2 30867 1 2583
2 30868 1 2583
2 30869 1 2583
2 30870 1 2583
2 30871 1 2583
2 30872 1 2590
2 30873 1 2590
2 30874 1 2597
2 30875 1 2597
2 30876 1 2597
2 30877 1 2598
2 30878 1 2598
2 30879 1 2598
2 30880 1 2598
2 30881 1 2607
2 30882 1 2607
2 30883 1 2617
2 30884 1 2617
2 30885 1 2620
2 30886 1 2620
2 30887 1 2620
2 30888 1 2621
2 30889 1 2621
2 30890 1 2622
2 30891 1 2622
2 30892 1 2624
2 30893 1 2624
2 30894 1 2625
2 30895 1 2625
2 30896 1 2625
2 30897 1 2625
2 30898 1 2625
2 30899 1 2625
2 30900 1 2625
2 30901 1 2625
2 30902 1 2625
2 30903 1 2629
2 30904 1 2629
2 30905 1 2629
2 30906 1 2629
2 30907 1 2629
2 30908 1 2629
2 30909 1 2630
2 30910 1 2630
2 30911 1 2645
2 30912 1 2645
2 30913 1 2646
2 30914 1 2646
2 30915 1 2648
2 30916 1 2648
2 30917 1 2649
2 30918 1 2649
2 30919 1 2651
2 30920 1 2651
2 30921 1 2654
2 30922 1 2654
2 30923 1 2657
2 30924 1 2657
2 30925 1 2657
2 30926 1 2657
2 30927 1 2657
2 30928 1 2664
2 30929 1 2664
2 30930 1 2664
2 30931 1 2672
2 30932 1 2672
2 30933 1 2696
2 30934 1 2696
2 30935 1 2696
2 30936 1 2696
2 30937 1 2696
2 30938 1 2696
2 30939 1 2696
2 30940 1 2696
2 30941 1 2696
2 30942 1 2696
2 30943 1 2696
2 30944 1 2696
2 30945 1 2699
2 30946 1 2699
2 30947 1 2699
2 30948 1 2701
2 30949 1 2701
2 30950 1 2701
2 30951 1 2701
2 30952 1 2701
2 30953 1 2701
2 30954 1 2701
2 30955 1 2707
2 30956 1 2707
2 30957 1 2710
2 30958 1 2710
2 30959 1 2710
2 30960 1 2710
2 30961 1 2710
2 30962 1 2711
2 30963 1 2711
2 30964 1 2713
2 30965 1 2713
2 30966 1 2718
2 30967 1 2718
2 30968 1 2721
2 30969 1 2721
2 30970 1 2735
2 30971 1 2735
2 30972 1 2735
2 30973 1 2735
2 30974 1 2735
2 30975 1 2735
2 30976 1 2735
2 30977 1 2735
2 30978 1 2735
2 30979 1 2735
2 30980 1 2735
2 30981 1 2735
2 30982 1 2735
2 30983 1 2735
2 30984 1 2735
2 30985 1 2735
2 30986 1 2735
2 30987 1 2735
2 30988 1 2736
2 30989 1 2736
2 30990 1 2737
2 30991 1 2737
2 30992 1 2737
2 30993 1 2737
2 30994 1 2737
2 30995 1 2737
2 30996 1 2737
2 30997 1 2737
2 30998 1 2756
2 30999 1 2756
2 31000 1 2756
2 31001 1 2756
2 31002 1 2757
2 31003 1 2757
2 31004 1 2760
2 31005 1 2760
2 31006 1 2760
2 31007 1 2760
2 31008 1 2760
2 31009 1 2760
2 31010 1 2760
2 31011 1 2760
2 31012 1 2760
2 31013 1 2760
2 31014 1 2760
2 31015 1 2760
2 31016 1 2760
2 31017 1 2760
2 31018 1 2760
2 31019 1 2760
2 31020 1 2760
2 31021 1 2760
2 31022 1 2761
2 31023 1 2761
2 31024 1 2766
2 31025 1 2766
2 31026 1 2767
2 31027 1 2767
2 31028 1 2767
2 31029 1 2767
2 31030 1 2767
2 31031 1 2767
2 31032 1 2767
2 31033 1 2767
2 31034 1 2767
2 31035 1 2767
2 31036 1 2767
2 31037 1 2767
2 31038 1 2767
2 31039 1 2767
2 31040 1 2768
2 31041 1 2768
2 31042 1 2785
2 31043 1 2785
2 31044 1 2798
2 31045 1 2798
2 31046 1 2798
2 31047 1 2798
2 31048 1 2799
2 31049 1 2799
2 31050 1 2800
2 31051 1 2800
2 31052 1 2800
2 31053 1 2800
2 31054 1 2800
2 31055 1 2801
2 31056 1 2801
2 31057 1 2801
2 31058 1 2801
2 31059 1 2801
2 31060 1 2815
2 31061 1 2815
2 31062 1 2815
2 31063 1 2816
2 31064 1 2816
2 31065 1 2817
2 31066 1 2817
2 31067 1 2817
2 31068 1 2817
2 31069 1 2818
2 31070 1 2818
2 31071 1 2818
2 31072 1 2840
2 31073 1 2840
2 31074 1 2840
2 31075 1 2840
2 31076 1 2840
2 31077 1 2840
2 31078 1 2843
2 31079 1 2843
2 31080 1 2856
2 31081 1 2856
2 31082 1 2863
2 31083 1 2863
2 31084 1 2870
2 31085 1 2870
2 31086 1 2870
2 31087 1 2870
2 31088 1 2870
2 31089 1 2872
2 31090 1 2872
2 31091 1 2872
2 31092 1 2872
2 31093 1 2872
2 31094 1 2872
2 31095 1 2888
2 31096 1 2888
2 31097 1 2888
2 31098 1 2894
2 31099 1 2894
2 31100 1 2916
2 31101 1 2916
2 31102 1 2916
2 31103 1 2916
2 31104 1 2916
2 31105 1 2916
2 31106 1 2916
2 31107 1 2916
2 31108 1 2917
2 31109 1 2917
2 31110 1 2917
2 31111 1 2917
2 31112 1 2917
2 31113 1 2917
2 31114 1 2917
2 31115 1 2917
2 31116 1 2917
2 31117 1 2917
2 31118 1 2917
2 31119 1 2917
2 31120 1 2917
2 31121 1 2917
2 31122 1 2917
2 31123 1 2917
2 31124 1 2917
2 31125 1 2917
2 31126 1 2917
2 31127 1 2917
2 31128 1 2917
2 31129 1 2917
2 31130 1 2918
2 31131 1 2918
2 31132 1 2918
2 31133 1 2918
2 31134 1 2918
2 31135 1 2918
2 31136 1 2921
2 31137 1 2921
2 31138 1 2922
2 31139 1 2922
2 31140 1 2922
2 31141 1 2922
2 31142 1 2925
2 31143 1 2925
2 31144 1 2925
2 31145 1 2925
2 31146 1 2925
2 31147 1 2936
2 31148 1 2936
2 31149 1 2937
2 31150 1 2937
2 31151 1 2937
2 31152 1 2938
2 31153 1 2938
2 31154 1 2938
2 31155 1 2941
2 31156 1 2941
2 31157 1 2941
2 31158 1 2941
2 31159 1 2941
2 31160 1 2941
2 31161 1 2941
2 31162 1 2941
2 31163 1 2941
2 31164 1 2941
2 31165 1 2941
2 31166 1 2941
2 31167 1 2948
2 31168 1 2948
2 31169 1 2948
2 31170 1 2948
2 31171 1 2952
2 31172 1 2952
2 31173 1 2952
2 31174 1 2952
2 31175 1 2952
2 31176 1 2952
2 31177 1 2952
2 31178 1 2964
2 31179 1 2964
2 31180 1 2973
2 31181 1 2973
2 31182 1 2973
2 31183 1 2974
2 31184 1 2974
2 31185 1 2974
2 31186 1 2974
2 31187 1 2974
2 31188 1 2974
2 31189 1 2974
2 31190 1 2974
2 31191 1 2974
2 31192 1 2974
2 31193 1 2974
2 31194 1 2974
2 31195 1 2974
2 31196 1 2974
2 31197 1 2974
2 31198 1 2974
2 31199 1 2974
2 31200 1 2975
2 31201 1 2975
2 31202 1 2975
2 31203 1 2975
2 31204 1 2975
2 31205 1 2976
2 31206 1 2976
2 31207 1 2976
2 31208 1 2991
2 31209 1 2991
2 31210 1 2991
2 31211 1 3019
2 31212 1 3019
2 31213 1 3019
2 31214 1 3019
2 31215 1 3019
2 31216 1 3019
2 31217 1 3019
2 31218 1 3019
2 31219 1 3019
2 31220 1 3019
2 31221 1 3019
2 31222 1 3019
2 31223 1 3021
2 31224 1 3021
2 31225 1 3022
2 31226 1 3022
2 31227 1 3022
2 31228 1 3022
2 31229 1 3022
2 31230 1 3022
2 31231 1 3022
2 31232 1 3023
2 31233 1 3023
2 31234 1 3023
2 31235 1 3023
2 31236 1 3023
2 31237 1 3023
2 31238 1 3023
2 31239 1 3023
2 31240 1 3023
2 31241 1 3028
2 31242 1 3028
2 31243 1 3036
2 31244 1 3036
2 31245 1 3045
2 31246 1 3045
2 31247 1 3045
2 31248 1 3046
2 31249 1 3046
2 31250 1 3048
2 31251 1 3048
2 31252 1 3048
2 31253 1 3055
2 31254 1 3055
2 31255 1 3055
2 31256 1 3057
2 31257 1 3057
2 31258 1 3058
2 31259 1 3058
2 31260 1 3058
2 31261 1 3066
2 31262 1 3066
2 31263 1 3066
2 31264 1 3066
2 31265 1 3066
2 31266 1 3066
2 31267 1 3067
2 31268 1 3067
2 31269 1 3070
2 31270 1 3070
2 31271 1 3070
2 31272 1 3071
2 31273 1 3071
2 31274 1 3072
2 31275 1 3072
2 31276 1 3072
2 31277 1 3072
2 31278 1 3072
2 31279 1 3072
2 31280 1 3072
2 31281 1 3072
2 31282 1 3073
2 31283 1 3073
2 31284 1 3078
2 31285 1 3078
2 31286 1 3079
2 31287 1 3079
2 31288 1 3081
2 31289 1 3081
2 31290 1 3082
2 31291 1 3082
2 31292 1 3083
2 31293 1 3083
2 31294 1 3083
2 31295 1 3084
2 31296 1 3084
2 31297 1 3108
2 31298 1 3108
2 31299 1 3108
2 31300 1 3108
2 31301 1 3112
2 31302 1 3112
2 31303 1 3112
2 31304 1 3112
2 31305 1 3112
2 31306 1 3113
2 31307 1 3113
2 31308 1 3113
2 31309 1 3113
2 31310 1 3113
2 31311 1 3114
2 31312 1 3114
2 31313 1 3115
2 31314 1 3115
2 31315 1 3123
2 31316 1 3123
2 31317 1 3123
2 31318 1 3123
2 31319 1 3123
2 31320 1 3123
2 31321 1 3123
2 31322 1 3123
2 31323 1 3123
2 31324 1 3123
2 31325 1 3123
2 31326 1 3126
2 31327 1 3126
2 31328 1 3127
2 31329 1 3127
2 31330 1 3127
2 31331 1 3127
2 31332 1 3128
2 31333 1 3128
2 31334 1 3128
2 31335 1 3137
2 31336 1 3137
2 31337 1 3137
2 31338 1 3137
2 31339 1 3137
2 31340 1 3137
2 31341 1 3139
2 31342 1 3139
2 31343 1 3140
2 31344 1 3140
2 31345 1 3140
2 31346 1 3140
2 31347 1 3140
2 31348 1 3140
2 31349 1 3140
2 31350 1 3153
2 31351 1 3153
2 31352 1 3155
2 31353 1 3155
2 31354 1 3155
2 31355 1 3155
2 31356 1 3155
2 31357 1 3155
2 31358 1 3155
2 31359 1 3158
2 31360 1 3158
2 31361 1 3159
2 31362 1 3159
2 31363 1 3159
2 31364 1 3159
2 31365 1 3159
2 31366 1 3163
2 31367 1 3163
2 31368 1 3163
2 31369 1 3163
2 31370 1 3166
2 31371 1 3166
2 31372 1 3167
2 31373 1 3167
2 31374 1 3167
2 31375 1 3167
2 31376 1 3176
2 31377 1 3176
2 31378 1 3176
2 31379 1 3183
2 31380 1 3183
2 31381 1 3199
2 31382 1 3199
2 31383 1 3202
2 31384 1 3202
2 31385 1 3210
2 31386 1 3210
2 31387 1 3210
2 31388 1 3210
2 31389 1 3210
2 31390 1 3212
2 31391 1 3212
2 31392 1 3212
2 31393 1 3220
2 31394 1 3220
2 31395 1 3220
2 31396 1 3220
2 31397 1 3220
2 31398 1 3220
2 31399 1 3221
2 31400 1 3221
2 31401 1 3235
2 31402 1 3235
2 31403 1 3236
2 31404 1 3236
2 31405 1 3236
2 31406 1 3236
2 31407 1 3236
2 31408 1 3236
2 31409 1 3236
2 31410 1 3236
2 31411 1 3239
2 31412 1 3239
2 31413 1 3242
2 31414 1 3242
2 31415 1 3242
2 31416 1 3242
2 31417 1 3243
2 31418 1 3243
2 31419 1 3245
2 31420 1 3245
2 31421 1 3245
2 31422 1 3245
2 31423 1 3245
2 31424 1 3245
2 31425 1 3245
2 31426 1 3245
2 31427 1 3245
2 31428 1 3245
2 31429 1 3245
2 31430 1 3245
2 31431 1 3246
2 31432 1 3246
2 31433 1 3246
2 31434 1 3251
2 31435 1 3251
2 31436 1 3255
2 31437 1 3255
2 31438 1 3256
2 31439 1 3256
2 31440 1 3256
2 31441 1 3256
2 31442 1 3256
2 31443 1 3256
2 31444 1 3256
2 31445 1 3265
2 31446 1 3265
2 31447 1 3265
2 31448 1 3265
2 31449 1 3265
2 31450 1 3266
2 31451 1 3266
2 31452 1 3266
2 31453 1 3266
2 31454 1 3266
2 31455 1 3266
2 31456 1 3266
2 31457 1 3266
2 31458 1 3266
2 31459 1 3266
2 31460 1 3266
2 31461 1 3266
2 31462 1 3266
2 31463 1 3266
2 31464 1 3266
2 31465 1 3266
2 31466 1 3278
2 31467 1 3278
2 31468 1 3278
2 31469 1 3278
2 31470 1 3278
2 31471 1 3278
2 31472 1 3278
2 31473 1 3278
2 31474 1 3278
2 31475 1 3278
2 31476 1 3278
2 31477 1 3278
2 31478 1 3278
2 31479 1 3278
2 31480 1 3278
2 31481 1 3278
2 31482 1 3278
2 31483 1 3278
2 31484 1 3278
2 31485 1 3278
2 31486 1 3278
2 31487 1 3278
2 31488 1 3278
2 31489 1 3280
2 31490 1 3280
2 31491 1 3281
2 31492 1 3281
2 31493 1 3282
2 31494 1 3282
2 31495 1 3282
2 31496 1 3282
2 31497 1 3282
2 31498 1 3282
2 31499 1 3286
2 31500 1 3286
2 31501 1 3292
2 31502 1 3292
2 31503 1 3295
2 31504 1 3295
2 31505 1 3295
2 31506 1 3295
2 31507 1 3295
2 31508 1 3295
2 31509 1 3295
2 31510 1 3295
2 31511 1 3295
2 31512 1 3295
2 31513 1 3295
2 31514 1 3295
2 31515 1 3295
2 31516 1 3295
2 31517 1 3296
2 31518 1 3296
2 31519 1 3296
2 31520 1 3296
2 31521 1 3296
2 31522 1 3297
2 31523 1 3297
2 31524 1 3298
2 31525 1 3298
2 31526 1 3298
2 31527 1 3311
2 31528 1 3311
2 31529 1 3312
2 31530 1 3312
2 31531 1 3323
2 31532 1 3323
2 31533 1 3335
2 31534 1 3335
2 31535 1 3335
2 31536 1 3336
2 31537 1 3336
2 31538 1 3346
2 31539 1 3346
2 31540 1 3346
2 31541 1 3347
2 31542 1 3347
2 31543 1 3347
2 31544 1 3354
2 31545 1 3354
2 31546 1 3356
2 31547 1 3356
2 31548 1 3356
2 31549 1 3356
2 31550 1 3356
2 31551 1 3357
2 31552 1 3357
2 31553 1 3358
2 31554 1 3358
2 31555 1 3358
2 31556 1 3358
2 31557 1 3358
2 31558 1 3367
2 31559 1 3367
2 31560 1 3368
2 31561 1 3368
2 31562 1 3368
2 31563 1 3368
2 31564 1 3368
2 31565 1 3370
2 31566 1 3370
2 31567 1 3373
2 31568 1 3373
2 31569 1 3373
2 31570 1 3373
2 31571 1 3374
2 31572 1 3374
2 31573 1 3375
2 31574 1 3375
2 31575 1 3375
2 31576 1 3383
2 31577 1 3383
2 31578 1 3386
2 31579 1 3386
2 31580 1 3386
2 31581 1 3386
2 31582 1 3392
2 31583 1 3392
2 31584 1 3392
2 31585 1 3392
2 31586 1 3398
2 31587 1 3398
2 31588 1 3398
2 31589 1 3399
2 31590 1 3399
2 31591 1 3399
2 31592 1 3411
2 31593 1 3411
2 31594 1 3411
2 31595 1 3411
2 31596 1 3412
2 31597 1 3412
2 31598 1 3412
2 31599 1 3413
2 31600 1 3413
2 31601 1 3413
2 31602 1 3413
2 31603 1 3413
2 31604 1 3413
2 31605 1 3413
2 31606 1 3413
2 31607 1 3413
2 31608 1 3413
2 31609 1 3413
2 31610 1 3413
2 31611 1 3413
2 31612 1 3414
2 31613 1 3414
2 31614 1 3414
2 31615 1 3414
2 31616 1 3415
2 31617 1 3415
2 31618 1 3415
2 31619 1 3417
2 31620 1 3417
2 31621 1 3417
2 31622 1 3417
2 31623 1 3417
2 31624 1 3417
2 31625 1 3418
2 31626 1 3418
2 31627 1 3418
2 31628 1 3420
2 31629 1 3420
2 31630 1 3420
2 31631 1 3420
2 31632 1 3420
2 31633 1 3420
2 31634 1 3420
2 31635 1 3420
2 31636 1 3420
2 31637 1 3420
2 31638 1 3421
2 31639 1 3421
2 31640 1 3421
2 31641 1 3421
2 31642 1 3426
2 31643 1 3426
2 31644 1 3427
2 31645 1 3427
2 31646 1 3431
2 31647 1 3431
2 31648 1 3431
2 31649 1 3431
2 31650 1 3431
2 31651 1 3431
2 31652 1 3440
2 31653 1 3440
2 31654 1 3440
2 31655 1 3440
2 31656 1 3440
2 31657 1 3440
2 31658 1 3440
2 31659 1 3440
2 31660 1 3440
2 31661 1 3440
2 31662 1 3440
2 31663 1 3440
2 31664 1 3440
2 31665 1 3440
2 31666 1 3440
2 31667 1 3443
2 31668 1 3443
2 31669 1 3443
2 31670 1 3443
2 31671 1 3443
2 31672 1 3443
2 31673 1 3443
2 31674 1 3443
2 31675 1 3443
2 31676 1 3443
2 31677 1 3443
2 31678 1 3443
2 31679 1 3443
2 31680 1 3443
2 31681 1 3443
2 31682 1 3443
2 31683 1 3443
2 31684 1 3443
2 31685 1 3443
2 31686 1 3443
2 31687 1 3443
2 31688 1 3443
2 31689 1 3443
2 31690 1 3443
2 31691 1 3443
2 31692 1 3444
2 31693 1 3444
2 31694 1 3444
2 31695 1 3445
2 31696 1 3445
2 31697 1 3446
2 31698 1 3446
2 31699 1 3446
2 31700 1 3446
2 31701 1 3450
2 31702 1 3450
2 31703 1 3450
2 31704 1 3450
2 31705 1 3450
2 31706 1 3450
2 31707 1 3450
2 31708 1 3451
2 31709 1 3451
2 31710 1 3452
2 31711 1 3452
2 31712 1 3452
2 31713 1 3452
2 31714 1 3452
2 31715 1 3453
2 31716 1 3453
2 31717 1 3453
2 31718 1 3453
2 31719 1 3453
2 31720 1 3453
2 31721 1 3453
2 31722 1 3453
2 31723 1 3455
2 31724 1 3455
2 31725 1 3463
2 31726 1 3463
2 31727 1 3464
2 31728 1 3464
2 31729 1 3470
2 31730 1 3470
2 31731 1 3493
2 31732 1 3493
2 31733 1 3493
2 31734 1 3502
2 31735 1 3502
2 31736 1 3502
2 31737 1 3506
2 31738 1 3506
2 31739 1 3506
2 31740 1 3506
2 31741 1 3507
2 31742 1 3507
2 31743 1 3507
2 31744 1 3507
2 31745 1 3507
2 31746 1 3511
2 31747 1 3511
2 31748 1 3511
2 31749 1 3514
2 31750 1 3514
2 31751 1 3514
2 31752 1 3514
2 31753 1 3515
2 31754 1 3515
2 31755 1 3516
2 31756 1 3516
2 31757 1 3532
2 31758 1 3532
2 31759 1 3533
2 31760 1 3533
2 31761 1 3533
2 31762 1 3541
2 31763 1 3541
2 31764 1 3541
2 31765 1 3543
2 31766 1 3543
2 31767 1 3543
2 31768 1 3543
2 31769 1 3558
2 31770 1 3558
2 31771 1 3558
2 31772 1 3558
2 31773 1 3563
2 31774 1 3563
2 31775 1 3563
2 31776 1 3567
2 31777 1 3567
2 31778 1 3567
2 31779 1 3568
2 31780 1 3568
2 31781 1 3568
2 31782 1 3568
2 31783 1 3568
2 31784 1 3570
2 31785 1 3570
2 31786 1 3585
2 31787 1 3585
2 31788 1 3585
2 31789 1 3595
2 31790 1 3595
2 31791 1 3595
2 31792 1 3595
2 31793 1 3595
2 31794 1 3599
2 31795 1 3599
2 31796 1 3605
2 31797 1 3605
2 31798 1 3605
2 31799 1 3605
2 31800 1 3605
2 31801 1 3605
2 31802 1 3607
2 31803 1 3607
2 31804 1 3615
2 31805 1 3615
2 31806 1 3618
2 31807 1 3618
2 31808 1 3625
2 31809 1 3625
2 31810 1 3625
2 31811 1 3625
2 31812 1 3625
2 31813 1 3636
2 31814 1 3636
2 31815 1 3637
2 31816 1 3637
2 31817 1 3637
2 31818 1 3645
2 31819 1 3645
2 31820 1 3645
2 31821 1 3648
2 31822 1 3648
2 31823 1 3648
2 31824 1 3669
2 31825 1 3669
2 31826 1 3669
2 31827 1 3669
2 31828 1 3685
2 31829 1 3685
2 31830 1 3685
2 31831 1 3685
2 31832 1 3686
2 31833 1 3686
2 31834 1 3686
2 31835 1 3686
2 31836 1 3686
2 31837 1 3691
2 31838 1 3691
2 31839 1 3691
2 31840 1 3691
2 31841 1 3691
2 31842 1 3691
2 31843 1 3692
2 31844 1 3692
2 31845 1 3692
2 31846 1 3692
2 31847 1 3692
2 31848 1 3692
2 31849 1 3692
2 31850 1 3695
2 31851 1 3695
2 31852 1 3695
2 31853 1 3695
2 31854 1 3695
2 31855 1 3695
2 31856 1 3695
2 31857 1 3695
2 31858 1 3695
2 31859 1 3695
2 31860 1 3695
2 31861 1 3697
2 31862 1 3697
2 31863 1 3713
2 31864 1 3713
2 31865 1 3713
2 31866 1 3713
2 31867 1 3713
2 31868 1 3715
2 31869 1 3715
2 31870 1 3716
2 31871 1 3716
2 31872 1 3716
2 31873 1 3716
2 31874 1 3717
2 31875 1 3717
2 31876 1 3722
2 31877 1 3722
2 31878 1 3724
2 31879 1 3724
2 31880 1 3732
2 31881 1 3732
2 31882 1 3732
2 31883 1 3732
2 31884 1 3732
2 31885 1 3732
2 31886 1 3733
2 31887 1 3733
2 31888 1 3734
2 31889 1 3734
2 31890 1 3736
2 31891 1 3736
2 31892 1 3736
2 31893 1 3736
2 31894 1 3736
2 31895 1 3743
2 31896 1 3743
2 31897 1 3743
2 31898 1 3743
2 31899 1 3751
2 31900 1 3751
2 31901 1 3769
2 31902 1 3769
2 31903 1 3780
2 31904 1 3780
2 31905 1 3780
2 31906 1 3780
2 31907 1 3780
2 31908 1 3780
2 31909 1 3780
2 31910 1 3781
2 31911 1 3781
2 31912 1 3794
2 31913 1 3794
2 31914 1 3797
2 31915 1 3797
2 31916 1 3798
2 31917 1 3798
2 31918 1 3798
2 31919 1 3798
2 31920 1 3799
2 31921 1 3799
2 31922 1 3799
2 31923 1 3814
2 31924 1 3814
2 31925 1 3820
2 31926 1 3820
2 31927 1 3821
2 31928 1 3821
2 31929 1 3821
2 31930 1 3821
2 31931 1 3825
2 31932 1 3825
2 31933 1 3832
2 31934 1 3832
2 31935 1 3832
2 31936 1 3844
2 31937 1 3844
2 31938 1 3847
2 31939 1 3847
2 31940 1 3858
2 31941 1 3858
2 31942 1 3858
2 31943 1 3858
2 31944 1 3858
2 31945 1 3858
2 31946 1 3858
2 31947 1 3858
2 31948 1 3858
2 31949 1 3858
2 31950 1 3859
2 31951 1 3859
2 31952 1 3859
2 31953 1 3860
2 31954 1 3860
2 31955 1 3860
2 31956 1 3861
2 31957 1 3861
2 31958 1 3867
2 31959 1 3867
2 31960 1 3868
2 31961 1 3868
2 31962 1 3868
2 31963 1 3869
2 31964 1 3869
2 31965 1 3877
2 31966 1 3877
2 31967 1 3877
2 31968 1 3877
2 31969 1 3877
2 31970 1 3878
2 31971 1 3878
2 31972 1 3878
2 31973 1 3878
2 31974 1 3878
2 31975 1 3878
2 31976 1 3883
2 31977 1 3883
2 31978 1 3883
2 31979 1 3883
2 31980 1 3884
2 31981 1 3884
2 31982 1 3884
2 31983 1 3884
2 31984 1 3899
2 31985 1 3899
2 31986 1 3900
2 31987 1 3900
2 31988 1 3907
2 31989 1 3907
2 31990 1 3921
2 31991 1 3921
2 31992 1 3921
2 31993 1 3921
2 31994 1 3921
2 31995 1 3922
2 31996 1 3922
2 31997 1 3924
2 31998 1 3924
2 31999 1 3925
2 32000 1 3925
2 32001 1 3925
2 32002 1 3925
2 32003 1 3925
2 32004 1 3944
2 32005 1 3944
2 32006 1 3949
2 32007 1 3949
2 32008 1 3952
2 32009 1 3952
2 32010 1 3952
2 32011 1 3952
2 32012 1 3952
2 32013 1 3953
2 32014 1 3953
2 32015 1 3961
2 32016 1 3961
2 32017 1 3961
2 32018 1 3961
2 32019 1 3961
2 32020 1 3961
2 32021 1 3961
2 32022 1 3961
2 32023 1 3961
2 32024 1 3961
2 32025 1 3961
2 32026 1 3961
2 32027 1 3963
2 32028 1 3963
2 32029 1 3963
2 32030 1 3973
2 32031 1 3973
2 32032 1 3983
2 32033 1 3983
2 32034 1 3983
2 32035 1 3983
2 32036 1 3983
2 32037 1 3983
2 32038 1 3983
2 32039 1 3984
2 32040 1 3984
2 32041 1 3985
2 32042 1 3985
2 32043 1 4012
2 32044 1 4012
2 32045 1 4012
2 32046 1 4012
2 32047 1 4012
2 32048 1 4012
2 32049 1 4012
2 32050 1 4012
2 32051 1 4012
2 32052 1 4012
2 32053 1 4012
2 32054 1 4012
2 32055 1 4012
2 32056 1 4012
2 32057 1 4012
2 32058 1 4012
2 32059 1 4012
2 32060 1 4012
2 32061 1 4012
2 32062 1 4012
2 32063 1 4012
2 32064 1 4013
2 32065 1 4013
2 32066 1 4013
2 32067 1 4013
2 32068 1 4014
2 32069 1 4014
2 32070 1 4015
2 32071 1 4015
2 32072 1 4015
2 32073 1 4015
2 32074 1 4015
2 32075 1 4015
2 32076 1 4015
2 32077 1 4015
2 32078 1 4015
2 32079 1 4015
2 32080 1 4015
2 32081 1 4015
2 32082 1 4015
2 32083 1 4015
2 32084 1 4015
2 32085 1 4015
2 32086 1 4015
2 32087 1 4015
2 32088 1 4015
2 32089 1 4015
2 32090 1 4015
2 32091 1 4015
2 32092 1 4015
2 32093 1 4015
2 32094 1 4015
2 32095 1 4015
2 32096 1 4015
2 32097 1 4015
2 32098 1 4015
2 32099 1 4015
2 32100 1 4015
2 32101 1 4015
2 32102 1 4015
2 32103 1 4015
2 32104 1 4015
2 32105 1 4015
2 32106 1 4015
2 32107 1 4015
2 32108 1 4015
2 32109 1 4015
2 32110 1 4015
2 32111 1 4015
2 32112 1 4015
2 32113 1 4015
2 32114 1 4015
2 32115 1 4015
2 32116 1 4015
2 32117 1 4015
2 32118 1 4015
2 32119 1 4015
2 32120 1 4015
2 32121 1 4015
2 32122 1 4015
2 32123 1 4015
2 32124 1 4015
2 32125 1 4015
2 32126 1 4015
2 32127 1 4015
2 32128 1 4015
2 32129 1 4018
2 32130 1 4018
2 32131 1 4030
2 32132 1 4030
2 32133 1 4030
2 32134 1 4032
2 32135 1 4032
2 32136 1 4036
2 32137 1 4036
2 32138 1 4041
2 32139 1 4041
2 32140 1 4045
2 32141 1 4045
2 32142 1 4060
2 32143 1 4060
2 32144 1 4060
2 32145 1 4060
2 32146 1 4060
2 32147 1 4060
2 32148 1 4060
2 32149 1 4069
2 32150 1 4069
2 32151 1 4069
2 32152 1 4069
2 32153 1 4070
2 32154 1 4070
2 32155 1 4079
2 32156 1 4079
2 32157 1 4079
2 32158 1 4079
2 32159 1 4079
2 32160 1 4080
2 32161 1 4080
2 32162 1 4080
2 32163 1 4080
2 32164 1 4080
2 32165 1 4080
2 32166 1 4081
2 32167 1 4081
2 32168 1 4081
2 32169 1 4082
2 32170 1 4082
2 32171 1 4082
2 32172 1 4083
2 32173 1 4083
2 32174 1 4093
2 32175 1 4093
2 32176 1 4093
2 32177 1 4098
2 32178 1 4098
2 32179 1 4101
2 32180 1 4101
2 32181 1 4101
2 32182 1 4102
2 32183 1 4102
2 32184 1 4111
2 32185 1 4111
2 32186 1 4111
2 32187 1 4111
2 32188 1 4111
2 32189 1 4111
2 32190 1 4111
2 32191 1 4111
2 32192 1 4111
2 32193 1 4111
2 32194 1 4111
2 32195 1 4111
2 32196 1 4111
2 32197 1 4115
2 32198 1 4115
2 32199 1 4118
2 32200 1 4118
2 32201 1 4130
2 32202 1 4130
2 32203 1 4130
2 32204 1 4130
2 32205 1 4132
2 32206 1 4132
2 32207 1 4132
2 32208 1 4133
2 32209 1 4133
2 32210 1 4141
2 32211 1 4141
2 32212 1 4141
2 32213 1 4141
2 32214 1 4141
2 32215 1 4142
2 32216 1 4142
2 32217 1 4143
2 32218 1 4143
2 32219 1 4144
2 32220 1 4144
2 32221 1 4144
2 32222 1 4144
2 32223 1 4144
2 32224 1 4154
2 32225 1 4154
2 32226 1 4154
2 32227 1 4154
2 32228 1 4154
2 32229 1 4154
2 32230 1 4154
2 32231 1 4154
2 32232 1 4154
2 32233 1 4154
2 32234 1 4158
2 32235 1 4158
2 32236 1 4158
2 32237 1 4158
2 32238 1 4158
2 32239 1 4158
2 32240 1 4158
2 32241 1 4158
2 32242 1 4158
2 32243 1 4158
2 32244 1 4158
2 32245 1 4158
2 32246 1 4158
2 32247 1 4158
2 32248 1 4158
2 32249 1 4158
2 32250 1 4158
2 32251 1 4158
2 32252 1 4158
2 32253 1 4158
2 32254 1 4158
2 32255 1 4158
2 32256 1 4158
2 32257 1 4158
2 32258 1 4158
2 32259 1 4158
2 32260 1 4159
2 32261 1 4159
2 32262 1 4159
2 32263 1 4170
2 32264 1 4170
2 32265 1 4184
2 32266 1 4184
2 32267 1 4187
2 32268 1 4187
2 32269 1 4187
2 32270 1 4188
2 32271 1 4188
2 32272 1 4195
2 32273 1 4195
2 32274 1 4205
2 32275 1 4205
2 32276 1 4205
2 32277 1 4205
2 32278 1 4208
2 32279 1 4208
2 32280 1 4208
2 32281 1 4209
2 32282 1 4209
2 32283 1 4212
2 32284 1 4212
2 32285 1 4215
2 32286 1 4215
2 32287 1 4215
2 32288 1 4215
2 32289 1 4215
2 32290 1 4215
2 32291 1 4250
2 32292 1 4250
2 32293 1 4250
2 32294 1 4251
2 32295 1 4251
2 32296 1 4261
2 32297 1 4261
2 32298 1 4262
2 32299 1 4262
2 32300 1 4270
2 32301 1 4270
2 32302 1 4271
2 32303 1 4271
2 32304 1 4301
2 32305 1 4301
2 32306 1 4303
2 32307 1 4303
2 32308 1 4304
2 32309 1 4304
2 32310 1 4304
2 32311 1 4304
2 32312 1 4304
2 32313 1 4304
2 32314 1 4304
2 32315 1 4305
2 32316 1 4305
2 32317 1 4315
2 32318 1 4315
2 32319 1 4315
2 32320 1 4315
2 32321 1 4315
2 32322 1 4315
2 32323 1 4316
2 32324 1 4316
2 32325 1 4316
2 32326 1 4316
2 32327 1 4316
2 32328 1 4316
2 32329 1 4316
2 32330 1 4316
2 32331 1 4316
2 32332 1 4316
2 32333 1 4316
2 32334 1 4316
2 32335 1 4316
2 32336 1 4316
2 32337 1 4316
2 32338 1 4317
2 32339 1 4317
2 32340 1 4327
2 32341 1 4327
2 32342 1 4328
2 32343 1 4328
2 32344 1 4328
2 32345 1 4328
2 32346 1 4328
2 32347 1 4328
2 32348 1 4328
2 32349 1 4329
2 32350 1 4329
2 32351 1 4329
2 32352 1 4329
2 32353 1 4341
2 32354 1 4341
2 32355 1 4341
2 32356 1 4341
2 32357 1 4342
2 32358 1 4342
2 32359 1 4342
2 32360 1 4344
2 32361 1 4344
2 32362 1 4344
2 32363 1 4344
2 32364 1 4344
2 32365 1 4359
2 32366 1 4359
2 32367 1 4359
2 32368 1 4359
2 32369 1 4359
2 32370 1 4359
2 32371 1 4364
2 32372 1 4364
2 32373 1 4364
2 32374 1 4365
2 32375 1 4365
2 32376 1 4374
2 32377 1 4374
2 32378 1 4374
2 32379 1 4375
2 32380 1 4375
2 32381 1 4375
2 32382 1 4375
2 32383 1 4375
2 32384 1 4384
2 32385 1 4384
2 32386 1 4384
2 32387 1 4404
2 32388 1 4404
2 32389 1 4404
2 32390 1 4404
2 32391 1 4404
2 32392 1 4404
2 32393 1 4404
2 32394 1 4404
2 32395 1 4406
2 32396 1 4406
2 32397 1 4406
2 32398 1 4406
2 32399 1 4406
2 32400 1 4406
2 32401 1 4406
2 32402 1 4408
2 32403 1 4408
2 32404 1 4415
2 32405 1 4415
2 32406 1 4415
2 32407 1 4415
2 32408 1 4459
2 32409 1 4459
2 32410 1 4459
2 32411 1 4460
2 32412 1 4460
2 32413 1 4460
2 32414 1 4486
2 32415 1 4486
2 32416 1 4486
2 32417 1 4486
2 32418 1 4493
2 32419 1 4493
2 32420 1 4493
2 32421 1 4494
2 32422 1 4494
2 32423 1 4494
2 32424 1 4504
2 32425 1 4504
2 32426 1 4507
2 32427 1 4507
2 32428 1 4526
2 32429 1 4526
2 32430 1 4527
2 32431 1 4527
2 32432 1 4527
2 32433 1 4532
2 32434 1 4532
2 32435 1 4532
2 32436 1 4533
2 32437 1 4533
2 32438 1 4533
2 32439 1 4533
2 32440 1 4533
2 32441 1 4533
2 32442 1 4535
2 32443 1 4535
2 32444 1 4535
2 32445 1 4535
2 32446 1 4535
2 32447 1 4535
2 32448 1 4536
2 32449 1 4536
2 32450 1 4538
2 32451 1 4538
2 32452 1 4538
2 32453 1 4538
2 32454 1 4538
2 32455 1 4538
2 32456 1 4538
2 32457 1 4538
2 32458 1 4538
2 32459 1 4538
2 32460 1 4538
2 32461 1 4538
2 32462 1 4538
2 32463 1 4539
2 32464 1 4539
2 32465 1 4539
2 32466 1 4541
2 32467 1 4541
2 32468 1 4541
2 32469 1 4541
2 32470 1 4541
2 32471 1 4541
2 32472 1 4541
2 32473 1 4541
2 32474 1 4541
2 32475 1 4542
2 32476 1 4542
2 32477 1 4543
2 32478 1 4543
2 32479 1 4546
2 32480 1 4546
2 32481 1 4546
2 32482 1 4546
2 32483 1 4546
2 32484 1 4546
2 32485 1 4546
2 32486 1 4546
2 32487 1 4546
2 32488 1 4546
2 32489 1 4546
2 32490 1 4546
2 32491 1 4546
2 32492 1 4546
2 32493 1 4546
2 32494 1 4549
2 32495 1 4549
2 32496 1 4551
2 32497 1 4551
2 32498 1 4551
2 32499 1 4555
2 32500 1 4555
2 32501 1 4556
2 32502 1 4556
2 32503 1 4556
2 32504 1 4560
2 32505 1 4560
2 32506 1 4561
2 32507 1 4561
2 32508 1 4569
2 32509 1 4569
2 32510 1 4569
2 32511 1 4569
2 32512 1 4569
2 32513 1 4569
2 32514 1 4569
2 32515 1 4569
2 32516 1 4569
2 32517 1 4569
2 32518 1 4569
2 32519 1 4569
2 32520 1 4571
2 32521 1 4571
2 32522 1 4571
2 32523 1 4571
2 32524 1 4571
2 32525 1 4571
2 32526 1 4571
2 32527 1 4571
2 32528 1 4571
2 32529 1 4571
2 32530 1 4571
2 32531 1 4571
2 32532 1 4571
2 32533 1 4571
2 32534 1 4571
2 32535 1 4571
2 32536 1 4573
2 32537 1 4573
2 32538 1 4574
2 32539 1 4574
2 32540 1 4574
2 32541 1 4574
2 32542 1 4574
2 32543 1 4574
2 32544 1 4574
2 32545 1 4574
2 32546 1 4574
2 32547 1 4574
2 32548 1 4574
2 32549 1 4574
2 32550 1 4574
2 32551 1 4574
2 32552 1 4574
2 32553 1 4574
2 32554 1 4574
2 32555 1 4574
2 32556 1 4574
2 32557 1 4574
2 32558 1 4574
2 32559 1 4574
2 32560 1 4574
2 32561 1 4574
2 32562 1 4574
2 32563 1 4574
2 32564 1 4575
2 32565 1 4575
2 32566 1 4575
2 32567 1 4575
2 32568 1 4575
2 32569 1 4577
2 32570 1 4577
2 32571 1 4577
2 32572 1 4577
2 32573 1 4577
2 32574 1 4577
2 32575 1 4577
2 32576 1 4577
2 32577 1 4577
2 32578 1 4577
2 32579 1 4577
2 32580 1 4577
2 32581 1 4577
2 32582 1 4577
2 32583 1 4577
2 32584 1 4577
2 32585 1 4577
2 32586 1 4577
2 32587 1 4577
2 32588 1 4577
2 32589 1 4577
2 32590 1 4577
2 32591 1 4577
2 32592 1 4577
2 32593 1 4577
2 32594 1 4577
2 32595 1 4577
2 32596 1 4577
2 32597 1 4578
2 32598 1 4578
2 32599 1 4578
2 32600 1 4578
2 32601 1 4584
2 32602 1 4584
2 32603 1 4584
2 32604 1 4584
2 32605 1 4584
2 32606 1 4585
2 32607 1 4585
2 32608 1 4585
2 32609 1 4585
2 32610 1 4585
2 32611 1 4585
2 32612 1 4585
2 32613 1 4585
2 32614 1 4585
2 32615 1 4585
2 32616 1 4585
2 32617 1 4585
2 32618 1 4585
2 32619 1 4585
2 32620 1 4585
2 32621 1 4587
2 32622 1 4587
2 32623 1 4587
2 32624 1 4587
2 32625 1 4587
2 32626 1 4587
2 32627 1 4590
2 32628 1 4590
2 32629 1 4590
2 32630 1 4590
2 32631 1 4590
2 32632 1 4590
2 32633 1 4590
2 32634 1 4590
2 32635 1 4590
2 32636 1 4590
2 32637 1 4590
2 32638 1 4590
2 32639 1 4590
2 32640 1 4590
2 32641 1 4590
2 32642 1 4590
2 32643 1 4592
2 32644 1 4592
2 32645 1 4592
2 32646 1 4592
2 32647 1 4592
2 32648 1 4592
2 32649 1 4596
2 32650 1 4596
2 32651 1 4596
2 32652 1 4596
2 32653 1 4596
2 32654 1 4596
2 32655 1 4596
2 32656 1 4596
2 32657 1 4596
2 32658 1 4596
2 32659 1 4596
2 32660 1 4599
2 32661 1 4599
2 32662 1 4599
2 32663 1 4599
2 32664 1 4599
2 32665 1 4600
2 32666 1 4600
2 32667 1 4601
2 32668 1 4601
2 32669 1 4604
2 32670 1 4604
2 32671 1 4614
2 32672 1 4614
2 32673 1 4614
2 32674 1 4617
2 32675 1 4617
2 32676 1 4634
2 32677 1 4634
2 32678 1 4634
2 32679 1 4634
2 32680 1 4641
2 32681 1 4641
2 32682 1 4641
2 32683 1 4641
2 32684 1 4641
2 32685 1 4650
2 32686 1 4650
2 32687 1 4650
2 32688 1 4650
2 32689 1 4650
2 32690 1 4651
2 32691 1 4651
2 32692 1 4656
2 32693 1 4656
2 32694 1 4657
2 32695 1 4657
2 32696 1 4657
2 32697 1 4658
2 32698 1 4658
2 32699 1 4659
2 32700 1 4659
2 32701 1 4659
2 32702 1 4659
2 32703 1 4659
2 32704 1 4668
2 32705 1 4668
2 32706 1 4668
2 32707 1 4668
2 32708 1 4668
2 32709 1 4668
2 32710 1 4669
2 32711 1 4669
2 32712 1 4671
2 32713 1 4671
2 32714 1 4671
2 32715 1 4671
2 32716 1 4671
2 32717 1 4672
2 32718 1 4672
2 32719 1 4672
2 32720 1 4675
2 32721 1 4675
2 32722 1 4675
2 32723 1 4675
2 32724 1 4675
2 32725 1 4675
2 32726 1 4675
2 32727 1 4675
2 32728 1 4675
2 32729 1 4675
2 32730 1 4675
2 32731 1 4675
2 32732 1 4675
2 32733 1 4675
2 32734 1 4675
2 32735 1 4675
2 32736 1 4675
2 32737 1 4675
2 32738 1 4675
2 32739 1 4675
2 32740 1 4675
2 32741 1 4675
2 32742 1 4675
2 32743 1 4676
2 32744 1 4676
2 32745 1 4677
2 32746 1 4677
2 32747 1 4677
2 32748 1 4677
2 32749 1 4680
2 32750 1 4680
2 32751 1 4680
2 32752 1 4680
2 32753 1 4683
2 32754 1 4683
2 32755 1 4683
2 32756 1 4683
2 32757 1 4683
2 32758 1 4683
2 32759 1 4683
2 32760 1 4683
2 32761 1 4683
2 32762 1 4683
2 32763 1 4683
2 32764 1 4683
2 32765 1 4683
2 32766 1 4683
2 32767 1 4685
2 32768 1 4685
2 32769 1 4685
2 32770 1 4685
2 32771 1 4686
2 32772 1 4686
2 32773 1 4686
2 32774 1 4690
2 32775 1 4690
2 32776 1 4690
2 32777 1 4692
2 32778 1 4692
2 32779 1 4692
2 32780 1 4692
2 32781 1 4697
2 32782 1 4697
2 32783 1 4699
2 32784 1 4699
2 32785 1 4702
2 32786 1 4702
2 32787 1 4705
2 32788 1 4705
2 32789 1 4705
2 32790 1 4705
2 32791 1 4705
2 32792 1 4707
2 32793 1 4707
2 32794 1 4707
2 32795 1 4707
2 32796 1 4707
2 32797 1 4707
2 32798 1 4710
2 32799 1 4710
2 32800 1 4710
2 32801 1 4710
2 32802 1 4710
2 32803 1 4710
2 32804 1 4710
2 32805 1 4710
2 32806 1 4710
2 32807 1 4710
2 32808 1 4710
2 32809 1 4710
2 32810 1 4710
2 32811 1 4710
2 32812 1 4711
2 32813 1 4711
2 32814 1 4714
2 32815 1 4714
2 32816 1 4714
2 32817 1 4714
2 32818 1 4715
2 32819 1 4715
2 32820 1 4715
2 32821 1 4715
2 32822 1 4715
2 32823 1 4715
2 32824 1 4716
2 32825 1 4716
2 32826 1 4717
2 32827 1 4717
2 32828 1 4717
2 32829 1 4718
2 32830 1 4718
2 32831 1 4721
2 32832 1 4721
2 32833 1 4721
2 32834 1 4721
2 32835 1 4721
2 32836 1 4721
2 32837 1 4728
2 32838 1 4728
2 32839 1 4736
2 32840 1 4736
2 32841 1 4737
2 32842 1 4737
2 32843 1 4737
2 32844 1 4737
2 32845 1 4751
2 32846 1 4751
2 32847 1 4751
2 32848 1 4751
2 32849 1 4751
2 32850 1 4751
2 32851 1 4751
2 32852 1 4751
2 32853 1 4751
2 32854 1 4757
2 32855 1 4757
2 32856 1 4757
2 32857 1 4761
2 32858 1 4761
2 32859 1 4761
2 32860 1 4761
2 32861 1 4761
2 32862 1 4762
2 32863 1 4762
2 32864 1 4762
2 32865 1 4770
2 32866 1 4770
2 32867 1 4772
2 32868 1 4772
2 32869 1 4772
2 32870 1 4772
2 32871 1 4772
2 32872 1 4774
2 32873 1 4774
2 32874 1 4774
2 32875 1 4774
2 32876 1 4774
2 32877 1 4778
2 32878 1 4778
2 32879 1 4778
2 32880 1 4778
2 32881 1 4778
2 32882 1 4778
2 32883 1 4778
2 32884 1 4779
2 32885 1 4779
2 32886 1 4780
2 32887 1 4780
2 32888 1 4781
2 32889 1 4781
2 32890 1 4781
2 32891 1 4781
2 32892 1 4782
2 32893 1 4782
2 32894 1 4792
2 32895 1 4792
2 32896 1 4792
2 32897 1 4792
2 32898 1 4792
2 32899 1 4792
2 32900 1 4792
2 32901 1 4792
2 32902 1 4792
2 32903 1 4792
2 32904 1 4792
2 32905 1 4794
2 32906 1 4794
2 32907 1 4795
2 32908 1 4795
2 32909 1 4795
2 32910 1 4795
2 32911 1 4799
2 32912 1 4799
2 32913 1 4799
2 32914 1 4799
2 32915 1 4799
2 32916 1 4800
2 32917 1 4800
2 32918 1 4800
2 32919 1 4800
2 32920 1 4800
2 32921 1 4801
2 32922 1 4801
2 32923 1 4802
2 32924 1 4802
2 32925 1 4802
2 32926 1 4802
2 32927 1 4805
2 32928 1 4805
2 32929 1 4805
2 32930 1 4805
2 32931 1 4805
2 32932 1 4805
2 32933 1 4805
2 32934 1 4805
2 32935 1 4805
2 32936 1 4805
2 32937 1 4805
2 32938 1 4805
2 32939 1 4819
2 32940 1 4819
2 32941 1 4819
2 32942 1 4819
2 32943 1 4823
2 32944 1 4823
2 32945 1 4823
2 32946 1 4823
2 32947 1 4826
2 32948 1 4826
2 32949 1 4829
2 32950 1 4829
2 32951 1 4833
2 32952 1 4833
2 32953 1 4833
2 32954 1 4833
2 32955 1 4836
2 32956 1 4836
2 32957 1 4836
2 32958 1 4838
2 32959 1 4838
2 32960 1 4838
2 32961 1 4841
2 32962 1 4841
2 32963 1 4841
2 32964 1 4841
2 32965 1 4841
2 32966 1 4841
2 32967 1 4842
2 32968 1 4842
2 32969 1 4843
2 32970 1 4843
2 32971 1 4843
2 32972 1 4843
2 32973 1 4843
2 32974 1 4852
2 32975 1 4852
2 32976 1 4853
2 32977 1 4853
2 32978 1 4853
2 32979 1 4858
2 32980 1 4858
2 32981 1 4858
2 32982 1 4871
2 32983 1 4871
2 32984 1 4871
2 32985 1 4871
2 32986 1 4871
2 32987 1 4871
2 32988 1 4871
2 32989 1 4871
2 32990 1 4871
2 32991 1 4871
2 32992 1 4871
2 32993 1 4871
2 32994 1 4871
2 32995 1 4871
2 32996 1 4871
2 32997 1 4871
2 32998 1 4871
2 32999 1 4872
2 33000 1 4872
2 33001 1 4872
2 33002 1 4872
2 33003 1 4879
2 33004 1 4879
2 33005 1 4879
2 33006 1 4879
2 33007 1 4879
2 33008 1 4887
2 33009 1 4887
2 33010 1 4887
2 33011 1 4887
2 33012 1 4888
2 33013 1 4888
2 33014 1 4888
2 33015 1 4888
2 33016 1 4889
2 33017 1 4889
2 33018 1 4890
2 33019 1 4890
2 33020 1 4891
2 33021 1 4891
2 33022 1 4902
2 33023 1 4902
2 33024 1 4902
2 33025 1 4905
2 33026 1 4905
2 33027 1 4910
2 33028 1 4910
2 33029 1 4912
2 33030 1 4912
2 33031 1 4912
2 33032 1 4912
2 33033 1 4913
2 33034 1 4913
2 33035 1 4916
2 33036 1 4916
2 33037 1 4916
2 33038 1 4916
2 33039 1 4916
2 33040 1 4919
2 33041 1 4919
2 33042 1 4919
2 33043 1 4919
2 33044 1 4919
2 33045 1 4920
2 33046 1 4920
2 33047 1 4923
2 33048 1 4923
2 33049 1 4923
2 33050 1 4928
2 33051 1 4928
2 33052 1 4939
2 33053 1 4939
2 33054 1 4939
2 33055 1 4939
2 33056 1 4939
2 33057 1 4939
2 33058 1 4939
2 33059 1 4939
2 33060 1 4939
2 33061 1 4939
2 33062 1 4939
2 33063 1 4939
2 33064 1 4939
2 33065 1 4939
2 33066 1 4940
2 33067 1 4940
2 33068 1 4940
2 33069 1 4941
2 33070 1 4941
2 33071 1 4941
2 33072 1 4942
2 33073 1 4942
2 33074 1 4944
2 33075 1 4944
2 33076 1 4944
2 33077 1 4944
2 33078 1 4944
2 33079 1 4944
2 33080 1 4947
2 33081 1 4947
2 33082 1 4948
2 33083 1 4948
2 33084 1 4948
2 33085 1 4948
2 33086 1 4948
2 33087 1 4964
2 33088 1 4964
2 33089 1 4964
2 33090 1 4981
2 33091 1 4981
2 33092 1 4981
2 33093 1 4981
2 33094 1 4981
2 33095 1 4981
2 33096 1 4981
2 33097 1 4982
2 33098 1 4982
2 33099 1 4982
2 33100 1 4982
2 33101 1 4983
2 33102 1 4983
2 33103 1 4983
2 33104 1 4983
2 33105 1 4983
2 33106 1 4983
2 33107 1 4983
2 33108 1 4986
2 33109 1 4986
2 33110 1 4998
2 33111 1 4998
2 33112 1 4998
2 33113 1 4998
2 33114 1 5011
2 33115 1 5011
2 33116 1 5012
2 33117 1 5012
2 33118 1 5012
2 33119 1 5012
2 33120 1 5025
2 33121 1 5025
2 33122 1 5030
2 33123 1 5030
2 33124 1 5030
2 33125 1 5032
2 33126 1 5032
2 33127 1 5035
2 33128 1 5035
2 33129 1 5035
2 33130 1 5035
2 33131 1 5035
2 33132 1 5047
2 33133 1 5047
2 33134 1 5047
2 33135 1 5047
2 33136 1 5047
2 33137 1 5047
2 33138 1 5047
2 33139 1 5049
2 33140 1 5049
2 33141 1 5049
2 33142 1 5049
2 33143 1 5049
2 33144 1 5049
2 33145 1 5049
2 33146 1 5049
2 33147 1 5049
2 33148 1 5049
2 33149 1 5049
2 33150 1 5049
2 33151 1 5049
2 33152 1 5049
2 33153 1 5049
2 33154 1 5053
2 33155 1 5053
2 33156 1 5053
2 33157 1 5056
2 33158 1 5056
2 33159 1 5056
2 33160 1 5056
2 33161 1 5056
2 33162 1 5056
2 33163 1 5056
2 33164 1 5056
2 33165 1 5056
2 33166 1 5057
2 33167 1 5057
2 33168 1 5057
2 33169 1 5057
2 33170 1 5060
2 33171 1 5060
2 33172 1 5063
2 33173 1 5063
2 33174 1 5064
2 33175 1 5064
2 33176 1 5069
2 33177 1 5069
2 33178 1 5076
2 33179 1 5076
2 33180 1 5076
2 33181 1 5076
2 33182 1 5076
2 33183 1 5078
2 33184 1 5078
2 33185 1 5078
2 33186 1 5079
2 33187 1 5079
2 33188 1 5081
2 33189 1 5081
2 33190 1 5081
2 33191 1 5081
2 33192 1 5081
2 33193 1 5085
2 33194 1 5085
2 33195 1 5085
2 33196 1 5105
2 33197 1 5105
2 33198 1 5105
2 33199 1 5106
2 33200 1 5106
2 33201 1 5106
2 33202 1 5106
2 33203 1 5107
2 33204 1 5107
2 33205 1 5115
2 33206 1 5115
2 33207 1 5129
2 33208 1 5129
2 33209 1 5129
2 33210 1 5135
2 33211 1 5135
2 33212 1 5135
2 33213 1 5135
2 33214 1 5135
2 33215 1 5139
2 33216 1 5139
2 33217 1 5142
2 33218 1 5142
2 33219 1 5142
2 33220 1 5160
2 33221 1 5160
2 33222 1 5160
2 33223 1 5160
2 33224 1 5160
2 33225 1 5160
2 33226 1 5160
2 33227 1 5161
2 33228 1 5161
2 33229 1 5175
2 33230 1 5175
2 33231 1 5175
2 33232 1 5176
2 33233 1 5176
2 33234 1 5187
2 33235 1 5187
2 33236 1 5187
2 33237 1 5187
2 33238 1 5187
2 33239 1 5187
2 33240 1 5187
2 33241 1 5187
2 33242 1 5187
2 33243 1 5187
2 33244 1 5187
2 33245 1 5187
2 33246 1 5187
2 33247 1 5190
2 33248 1 5190
2 33249 1 5190
2 33250 1 5214
2 33251 1 5214
2 33252 1 5214
2 33253 1 5214
2 33254 1 5214
2 33255 1 5214
2 33256 1 5218
2 33257 1 5218
2 33258 1 5218
2 33259 1 5225
2 33260 1 5225
2 33261 1 5225
2 33262 1 5230
2 33263 1 5230
2 33264 1 5239
2 33265 1 5239
2 33266 1 5240
2 33267 1 5240
2 33268 1 5251
2 33269 1 5251
2 33270 1 5251
2 33271 1 5256
2 33272 1 5256
2 33273 1 5269
2 33274 1 5269
2 33275 1 5269
2 33276 1 5269
2 33277 1 5269
2 33278 1 5269
2 33279 1 5271
2 33280 1 5271
2 33281 1 5271
2 33282 1 5271
2 33283 1 5275
2 33284 1 5275
2 33285 1 5278
2 33286 1 5278
2 33287 1 5278
2 33288 1 5278
2 33289 1 5278
2 33290 1 5278
2 33291 1 5278
2 33292 1 5279
2 33293 1 5279
2 33294 1 5292
2 33295 1 5292
2 33296 1 5293
2 33297 1 5293
2 33298 1 5293
2 33299 1 5298
2 33300 1 5298
2 33301 1 5299
2 33302 1 5299
2 33303 1 5303
2 33304 1 5303
2 33305 1 5303
2 33306 1 5304
2 33307 1 5304
2 33308 1 5304
2 33309 1 5308
2 33310 1 5308
2 33311 1 5309
2 33312 1 5309
2 33313 1 5342
2 33314 1 5342
2 33315 1 5350
2 33316 1 5350
2 33317 1 5353
2 33318 1 5353
2 33319 1 5356
2 33320 1 5356
2 33321 1 5356
2 33322 1 5356
2 33323 1 5356
2 33324 1 5356
2 33325 1 5356
2 33326 1 5356
2 33327 1 5368
2 33328 1 5368
2 33329 1 5368
2 33330 1 5368
2 33331 1 5368
2 33332 1 5368
2 33333 1 5369
2 33334 1 5369
2 33335 1 5377
2 33336 1 5377
2 33337 1 5377
2 33338 1 5389
2 33339 1 5389
2 33340 1 5389
2 33341 1 5389
2 33342 1 5405
2 33343 1 5405
2 33344 1 5434
2 33345 1 5434
2 33346 1 5434
2 33347 1 5434
2 33348 1 5435
2 33349 1 5435
2 33350 1 5439
2 33351 1 5439
2 33352 1 5467
2 33353 1 5467
2 33354 1 5475
2 33355 1 5475
2 33356 1 5475
2 33357 1 5475
2 33358 1 5475
2 33359 1 5475
2 33360 1 5475
2 33361 1 5475
2 33362 1 5475
2 33363 1 5475
2 33364 1 5475
2 33365 1 5475
2 33366 1 5475
2 33367 1 5476
2 33368 1 5476
2 33369 1 5476
2 33370 1 5479
2 33371 1 5479
2 33372 1 5479
2 33373 1 5479
2 33374 1 5479
2 33375 1 5479
2 33376 1 5479
2 33377 1 5479
2 33378 1 5479
2 33379 1 5487
2 33380 1 5487
2 33381 1 5488
2 33382 1 5488
2 33383 1 5488
2 33384 1 5488
2 33385 1 5496
2 33386 1 5496
2 33387 1 5497
2 33388 1 5497
2 33389 1 5497
2 33390 1 5497
2 33391 1 5555
2 33392 1 5555
2 33393 1 5562
2 33394 1 5562
2 33395 1 5562
2 33396 1 5562
2 33397 1 5562
2 33398 1 5593
2 33399 1 5593
2 33400 1 5593
2 33401 1 5593
2 33402 1 5593
2 33403 1 5593
2 33404 1 5593
2 33405 1 5593
2 33406 1 5593
2 33407 1 5594
2 33408 1 5594
2 33409 1 5594
2 33410 1 5594
2 33411 1 5594
2 33412 1 5594
2 33413 1 5599
2 33414 1 5599
2 33415 1 5599
2 33416 1 5599
2 33417 1 5599
2 33418 1 5599
2 33419 1 5599
2 33420 1 5599
2 33421 1 5599
2 33422 1 5599
2 33423 1 5599
2 33424 1 5599
2 33425 1 5599
2 33426 1 5599
2 33427 1 5600
2 33428 1 5600
2 33429 1 5600
2 33430 1 5600
2 33431 1 5601
2 33432 1 5601
2 33433 1 5609
2 33434 1 5609
2 33435 1 5610
2 33436 1 5610
2 33437 1 5610
2 33438 1 5610
2 33439 1 5618
2 33440 1 5618
2 33441 1 5620
2 33442 1 5620
2 33443 1 5620
2 33444 1 5620
2 33445 1 5620
2 33446 1 5620
2 33447 1 5620
2 33448 1 5620
2 33449 1 5621
2 33450 1 5621
2 33451 1 5621
2 33452 1 5621
2 33453 1 5621
2 33454 1 5621
2 33455 1 5621
2 33456 1 5621
2 33457 1 5621
2 33458 1 5621
2 33459 1 5621
2 33460 1 5631
2 33461 1 5631
2 33462 1 5631
2 33463 1 5631
2 33464 1 5634
2 33465 1 5634
2 33466 1 5634
2 33467 1 5635
2 33468 1 5635
2 33469 1 5635
2 33470 1 5635
2 33471 1 5635
2 33472 1 5635
2 33473 1 5635
2 33474 1 5637
2 33475 1 5637
2 33476 1 5645
2 33477 1 5645
2 33478 1 5645
2 33479 1 5645
2 33480 1 5645
2 33481 1 5645
2 33482 1 5645
2 33483 1 5645
2 33484 1 5648
2 33485 1 5648
2 33486 1 5648
2 33487 1 5648
2 33488 1 5648
2 33489 1 5650
2 33490 1 5650
2 33491 1 5650
2 33492 1 5651
2 33493 1 5651
2 33494 1 5659
2 33495 1 5659
2 33496 1 5659
2 33497 1 5659
2 33498 1 5659
2 33499 1 5659
2 33500 1 5659
2 33501 1 5659
2 33502 1 5660
2 33503 1 5660
2 33504 1 5660
2 33505 1 5661
2 33506 1 5661
2 33507 1 5661
2 33508 1 5661
2 33509 1 5661
2 33510 1 5663
2 33511 1 5663
2 33512 1 5664
2 33513 1 5664
2 33514 1 5664
2 33515 1 5664
2 33516 1 5664
2 33517 1 5664
2 33518 1 5668
2 33519 1 5668
2 33520 1 5675
2 33521 1 5675
2 33522 1 5675
2 33523 1 5675
2 33524 1 5675
2 33525 1 5675
2 33526 1 5684
2 33527 1 5684
2 33528 1 5684
2 33529 1 5684
2 33530 1 5685
2 33531 1 5685
2 33532 1 5685
2 33533 1 5685
2 33534 1 5686
2 33535 1 5686
2 33536 1 5686
2 33537 1 5689
2 33538 1 5689
2 33539 1 5689
2 33540 1 5690
2 33541 1 5690
2 33542 1 5692
2 33543 1 5692
2 33544 1 5695
2 33545 1 5695
2 33546 1 5697
2 33547 1 5697
2 33548 1 5697
2 33549 1 5697
2 33550 1 5697
2 33551 1 5697
2 33552 1 5697
2 33553 1 5697
2 33554 1 5697
2 33555 1 5697
2 33556 1 5697
2 33557 1 5697
2 33558 1 5697
2 33559 1 5697
2 33560 1 5697
2 33561 1 5697
2 33562 1 5697
2 33563 1 5697
2 33564 1 5698
2 33565 1 5698
2 33566 1 5698
2 33567 1 5698
2 33568 1 5698
2 33569 1 5698
2 33570 1 5698
2 33571 1 5698
2 33572 1 5698
2 33573 1 5698
2 33574 1 5698
2 33575 1 5698
2 33576 1 5698
2 33577 1 5698
2 33578 1 5698
2 33579 1 5699
2 33580 1 5699
2 33581 1 5699
2 33582 1 5699
2 33583 1 5699
2 33584 1 5699
2 33585 1 5719
2 33586 1 5719
2 33587 1 5719
2 33588 1 5720
2 33589 1 5720
2 33590 1 5720
2 33591 1 5730
2 33592 1 5730
2 33593 1 5730
2 33594 1 5738
2 33595 1 5738
2 33596 1 5741
2 33597 1 5741
2 33598 1 5741
2 33599 1 5744
2 33600 1 5744
2 33601 1 5744
2 33602 1 5744
2 33603 1 5744
2 33604 1 5744
2 33605 1 5746
2 33606 1 5746
2 33607 1 5749
2 33608 1 5749
2 33609 1 5749
2 33610 1 5756
2 33611 1 5756
2 33612 1 5757
2 33613 1 5757
2 33614 1 5759
2 33615 1 5759
2 33616 1 5759
2 33617 1 5759
2 33618 1 5759
2 33619 1 5759
2 33620 1 5765
2 33621 1 5765
2 33622 1 5766
2 33623 1 5766
2 33624 1 5766
2 33625 1 5766
2 33626 1 5767
2 33627 1 5767
2 33628 1 5767
2 33629 1 5767
2 33630 1 5775
2 33631 1 5775
2 33632 1 5775
2 33633 1 5775
2 33634 1 5775
2 33635 1 5775
2 33636 1 5775
2 33637 1 5775
2 33638 1 5775
2 33639 1 5775
2 33640 1 5775
2 33641 1 5775
2 33642 1 5777
2 33643 1 5777
2 33644 1 5777
2 33645 1 5785
2 33646 1 5785
2 33647 1 5785
2 33648 1 5785
2 33649 1 5785
2 33650 1 5785
2 33651 1 5786
2 33652 1 5786
2 33653 1 5786
2 33654 1 5786
2 33655 1 5786
2 33656 1 5786
2 33657 1 5786
2 33658 1 5786
2 33659 1 5786
2 33660 1 5786
2 33661 1 5786
2 33662 1 5786
2 33663 1 5786
2 33664 1 5786
2 33665 1 5787
2 33666 1 5787
2 33667 1 5787
2 33668 1 5787
2 33669 1 5788
2 33670 1 5788
2 33671 1 5788
2 33672 1 5788
2 33673 1 5788
2 33674 1 5788
2 33675 1 5788
2 33676 1 5788
2 33677 1 5788
2 33678 1 5788
2 33679 1 5788
2 33680 1 5788
2 33681 1 5788
2 33682 1 5788
2 33683 1 5788
2 33684 1 5788
2 33685 1 5788
2 33686 1 5788
2 33687 1 5790
2 33688 1 5790
2 33689 1 5793
2 33690 1 5793
2 33691 1 5793
2 33692 1 5793
2 33693 1 5793
2 33694 1 5793
2 33695 1 5796
2 33696 1 5796
2 33697 1 5796
2 33698 1 5798
2 33699 1 5798
2 33700 1 5798
2 33701 1 5798
2 33702 1 5798
2 33703 1 5798
2 33704 1 5798
2 33705 1 5798
2 33706 1 5798
2 33707 1 5799
2 33708 1 5799
2 33709 1 5807
2 33710 1 5807
2 33711 1 5807
2 33712 1 5807
2 33713 1 5808
2 33714 1 5808
2 33715 1 5808
2 33716 1 5808
2 33717 1 5808
2 33718 1 5810
2 33719 1 5810
2 33720 1 5810
2 33721 1 5810
2 33722 1 5810
2 33723 1 5810
2 33724 1 5810
2 33725 1 5810
2 33726 1 5810
2 33727 1 5811
2 33728 1 5811
2 33729 1 5811
2 33730 1 5811
2 33731 1 5812
2 33732 1 5812
2 33733 1 5820
2 33734 1 5820
2 33735 1 5820
2 33736 1 5820
2 33737 1 5820
2 33738 1 5820
2 33739 1 5820
2 33740 1 5820
2 33741 1 5821
2 33742 1 5821
2 33743 1 5821
2 33744 1 5829
2 33745 1 5829
2 33746 1 5829
2 33747 1 5838
2 33748 1 5838
2 33749 1 5839
2 33750 1 5839
2 33751 1 5846
2 33752 1 5846
2 33753 1 5847
2 33754 1 5847
2 33755 1 5848
2 33756 1 5848
2 33757 1 5849
2 33758 1 5849
2 33759 1 5849
2 33760 1 5849
2 33761 1 5849
2 33762 1 5850
2 33763 1 5850
2 33764 1 5858
2 33765 1 5858
2 33766 1 5859
2 33767 1 5859
2 33768 1 5859
2 33769 1 5859
2 33770 1 5859
2 33771 1 5859
2 33772 1 5863
2 33773 1 5863
2 33774 1 5863
2 33775 1 5863
2 33776 1 5863
2 33777 1 5863
2 33778 1 5865
2 33779 1 5865
2 33780 1 5865
2 33781 1 5865
2 33782 1 5865
2 33783 1 5865
2 33784 1 5865
2 33785 1 5865
2 33786 1 5866
2 33787 1 5866
2 33788 1 5876
2 33789 1 5876
2 33790 1 5876
2 33791 1 5876
2 33792 1 5876
2 33793 1 5876
2 33794 1 5877
2 33795 1 5877
2 33796 1 5877
2 33797 1 5882
2 33798 1 5882
2 33799 1 5882
2 33800 1 5882
2 33801 1 5882
2 33802 1 5882
2 33803 1 5882
2 33804 1 5882
2 33805 1 5882
2 33806 1 5882
2 33807 1 5884
2 33808 1 5884
2 33809 1 5885
2 33810 1 5885
2 33811 1 5891
2 33812 1 5891
2 33813 1 5891
2 33814 1 5891
2 33815 1 5891
2 33816 1 5891
2 33817 1 5891
2 33818 1 5891
2 33819 1 5892
2 33820 1 5892
2 33821 1 5892
2 33822 1 5892
2 33823 1 5892
2 33824 1 5900
2 33825 1 5900
2 33826 1 5900
2 33827 1 5900
2 33828 1 5901
2 33829 1 5901
2 33830 1 5908
2 33831 1 5908
2 33832 1 5909
2 33833 1 5909
2 33834 1 5909
2 33835 1 5909
2 33836 1 5909
2 33837 1 5909
2 33838 1 5910
2 33839 1 5910
2 33840 1 5910
2 33841 1 5911
2 33842 1 5911
2 33843 1 5914
2 33844 1 5914
2 33845 1 5914
2 33846 1 5914
2 33847 1 5914
2 33848 1 5914
2 33849 1 5914
2 33850 1 5914
2 33851 1 5915
2 33852 1 5915
2 33853 1 5915
2 33854 1 5915
2 33855 1 5915
2 33856 1 5917
2 33857 1 5917
2 33858 1 5918
2 33859 1 5918
2 33860 1 5918
2 33861 1 5918
2 33862 1 5918
2 33863 1 5942
2 33864 1 5942
2 33865 1 5942
2 33866 1 5942
2 33867 1 5942
2 33868 1 5943
2 33869 1 5943
2 33870 1 5956
2 33871 1 5956
2 33872 1 5957
2 33873 1 5957
2 33874 1 5962
2 33875 1 5962
2 33876 1 5962
2 33877 1 5962
2 33878 1 5965
2 33879 1 5965
2 33880 1 5965
2 33881 1 5978
2 33882 1 5978
2 33883 1 5978
2 33884 1 5979
2 33885 1 5979
2 33886 1 5979
2 33887 1 5989
2 33888 1 5989
2 33889 1 5992
2 33890 1 5992
2 33891 1 5992
2 33892 1 5993
2 33893 1 5993
2 33894 1 5996
2 33895 1 5996
2 33896 1 5996
2 33897 1 6002
2 33898 1 6002
2 33899 1 6002
2 33900 1 6002
2 33901 1 6002
2 33902 1 6002
2 33903 1 6011
2 33904 1 6011
2 33905 1 6012
2 33906 1 6012
2 33907 1 6020
2 33908 1 6020
2 33909 1 6020
2 33910 1 6020
2 33911 1 6020
2 33912 1 6020
2 33913 1 6020
2 33914 1 6020
2 33915 1 6021
2 33916 1 6021
2 33917 1 6022
2 33918 1 6022
2 33919 1 6022
2 33920 1 6024
2 33921 1 6024
2 33922 1 6024
2 33923 1 6024
2 33924 1 6024
2 33925 1 6024
2 33926 1 6025
2 33927 1 6025
2 33928 1 6027
2 33929 1 6027
2 33930 1 6027
2 33931 1 6027
2 33932 1 6027
2 33933 1 6027
2 33934 1 6027
2 33935 1 6027
2 33936 1 6027
2 33937 1 6027
2 33938 1 6027
2 33939 1 6027
2 33940 1 6028
2 33941 1 6028
2 33942 1 6028
2 33943 1 6028
2 33944 1 6028
2 33945 1 6028
2 33946 1 6028
2 33947 1 6028
2 33948 1 6031
2 33949 1 6031
2 33950 1 6032
2 33951 1 6032
2 33952 1 6034
2 33953 1 6034
2 33954 1 6035
2 33955 1 6035
2 33956 1 6035
2 33957 1 6035
2 33958 1 6035
2 33959 1 6035
2 33960 1 6035
2 33961 1 6035
2 33962 1 6035
2 33963 1 6035
2 33964 1 6035
2 33965 1 6035
2 33966 1 6035
2 33967 1 6035
2 33968 1 6038
2 33969 1 6038
2 33970 1 6039
2 33971 1 6039
2 33972 1 6039
2 33973 1 6042
2 33974 1 6042
2 33975 1 6042
2 33976 1 6042
2 33977 1 6042
2 33978 1 6042
2 33979 1 6042
2 33980 1 6042
2 33981 1 6042
2 33982 1 6042
2 33983 1 6042
2 33984 1 6042
2 33985 1 6042
2 33986 1 6042
2 33987 1 6042
2 33988 1 6042
2 33989 1 6042
2 33990 1 6042
2 33991 1 6042
2 33992 1 6047
2 33993 1 6047
2 33994 1 6047
2 33995 1 6047
2 33996 1 6047
2 33997 1 6047
2 33998 1 6050
2 33999 1 6050
2 34000 1 6050
2 34001 1 6051
2 34002 1 6051
2 34003 1 6058
2 34004 1 6058
2 34005 1 6058
2 34006 1 6058
2 34007 1 6058
2 34008 1 6058
2 34009 1 6058
2 34010 1 6058
2 34011 1 6058
2 34012 1 6058
2 34013 1 6058
2 34014 1 6058
2 34015 1 6058
2 34016 1 6059
2 34017 1 6059
2 34018 1 6064
2 34019 1 6064
2 34020 1 6070
2 34021 1 6070
2 34022 1 6070
2 34023 1 6070
2 34024 1 6070
2 34025 1 6070
2 34026 1 6070
2 34027 1 6070
2 34028 1 6070
2 34029 1 6070
2 34030 1 6070
2 34031 1 6070
2 34032 1 6070
2 34033 1 6070
2 34034 1 6070
2 34035 1 6070
2 34036 1 6070
2 34037 1 6070
2 34038 1 6070
2 34039 1 6071
2 34040 1 6071
2 34041 1 6073
2 34042 1 6073
2 34043 1 6073
2 34044 1 6073
2 34045 1 6074
2 34046 1 6074
2 34047 1 6074
2 34048 1 6074
2 34049 1 6090
2 34050 1 6090
2 34051 1 6095
2 34052 1 6095
2 34053 1 6095
2 34054 1 6095
2 34055 1 6095
2 34056 1 6095
2 34057 1 6095
2 34058 1 6098
2 34059 1 6098
2 34060 1 6111
2 34061 1 6111
2 34062 1 6111
2 34063 1 6111
2 34064 1 6111
2 34065 1 6111
2 34066 1 6111
2 34067 1 6111
2 34068 1 6111
2 34069 1 6111
2 34070 1 6111
2 34071 1 6112
2 34072 1 6112
2 34073 1 6112
2 34074 1 6112
2 34075 1 6112
2 34076 1 6112
2 34077 1 6112
2 34078 1 6112
2 34079 1 6112
2 34080 1 6112
2 34081 1 6112
2 34082 1 6112
2 34083 1 6112
2 34084 1 6113
2 34085 1 6113
2 34086 1 6113
2 34087 1 6113
2 34088 1 6113
2 34089 1 6113
2 34090 1 6113
2 34091 1 6113
2 34092 1 6113
2 34093 1 6115
2 34094 1 6115
2 34095 1 6115
2 34096 1 6115
2 34097 1 6115
2 34098 1 6118
2 34099 1 6118
2 34100 1 6118
2 34101 1 6123
2 34102 1 6123
2 34103 1 6128
2 34104 1 6128
2 34105 1 6128
2 34106 1 6134
2 34107 1 6134
2 34108 1 6140
2 34109 1 6140
2 34110 1 6148
2 34111 1 6148
2 34112 1 6163
2 34113 1 6163
2 34114 1 6163
2 34115 1 6163
2 34116 1 6167
2 34117 1 6167
2 34118 1 6167
2 34119 1 6167
2 34120 1 6170
2 34121 1 6170
2 34122 1 6174
2 34123 1 6174
2 34124 1 6174
2 34125 1 6174
2 34126 1 6174
2 34127 1 6174
2 34128 1 6178
2 34129 1 6178
2 34130 1 6180
2 34131 1 6180
2 34132 1 6180
2 34133 1 6180
2 34134 1 6180
2 34135 1 6180
2 34136 1 6180
2 34137 1 6180
2 34138 1 6180
2 34139 1 6180
2 34140 1 6180
2 34141 1 6180
2 34142 1 6180
2 34143 1 6180
2 34144 1 6180
2 34145 1 6180
2 34146 1 6180
2 34147 1 6180
2 34148 1 6195
2 34149 1 6195
2 34150 1 6195
2 34151 1 6195
2 34152 1 6195
2 34153 1 6203
2 34154 1 6203
2 34155 1 6203
2 34156 1 6203
2 34157 1 6203
2 34158 1 6203
2 34159 1 6203
2 34160 1 6204
2 34161 1 6204
2 34162 1 6204
2 34163 1 6205
2 34164 1 6205
2 34165 1 6205
2 34166 1 6205
2 34167 1 6205
2 34168 1 6205
2 34169 1 6205
2 34170 1 6205
2 34171 1 6206
2 34172 1 6206
2 34173 1 6206
2 34174 1 6206
2 34175 1 6206
2 34176 1 6206
2 34177 1 6207
2 34178 1 6207
2 34179 1 6207
2 34180 1 6207
2 34181 1 6207
2 34182 1 6210
2 34183 1 6210
2 34184 1 6211
2 34185 1 6211
2 34186 1 6211
2 34187 1 6212
2 34188 1 6212
2 34189 1 6214
2 34190 1 6214
2 34191 1 6214
2 34192 1 6214
2 34193 1 6214
2 34194 1 6215
2 34195 1 6215
2 34196 1 6222
2 34197 1 6222
2 34198 1 6222
2 34199 1 6222
2 34200 1 6222
2 34201 1 6223
2 34202 1 6223
2 34203 1 6236
2 34204 1 6236
2 34205 1 6236
2 34206 1 6236
2 34207 1 6236
2 34208 1 6236
2 34209 1 6241
2 34210 1 6241
2 34211 1 6242
2 34212 1 6242
2 34213 1 6244
2 34214 1 6244
2 34215 1 6247
2 34216 1 6247
2 34217 1 6250
2 34218 1 6250
2 34219 1 6250
2 34220 1 6253
2 34221 1 6253
2 34222 1 6256
2 34223 1 6256
2 34224 1 6256
2 34225 1 6256
2 34226 1 6256
2 34227 1 6256
2 34228 1 6257
2 34229 1 6257
2 34230 1 6257
2 34231 1 6258
2 34232 1 6258
2 34233 1 6258
2 34234 1 6258
2 34235 1 6258
2 34236 1 6266
2 34237 1 6266
2 34238 1 6267
2 34239 1 6267
2 34240 1 6274
2 34241 1 6274
2 34242 1 6274
2 34243 1 6276
2 34244 1 6276
2 34245 1 6277
2 34246 1 6277
2 34247 1 6277
2 34248 1 6279
2 34249 1 6279
2 34250 1 6281
2 34251 1 6281
2 34252 1 6281
2 34253 1 6281
2 34254 1 6281
2 34255 1 6282
2 34256 1 6282
2 34257 1 6282
2 34258 1 6294
2 34259 1 6294
2 34260 1 6294
2 34261 1 6294
2 34262 1 6297
2 34263 1 6297
2 34264 1 6315
2 34265 1 6315
2 34266 1 6315
2 34267 1 6316
2 34268 1 6316
2 34269 1 6317
2 34270 1 6317
2 34271 1 6317
2 34272 1 6317
2 34273 1 6317
2 34274 1 6317
2 34275 1 6317
2 34276 1 6317
2 34277 1 6318
2 34278 1 6318
2 34279 1 6318
2 34280 1 6318
2 34281 1 6318
2 34282 1 6318
2 34283 1 6318
2 34284 1 6318
2 34285 1 6319
2 34286 1 6319
2 34287 1 6322
2 34288 1 6322
2 34289 1 6322
2 34290 1 6322
2 34291 1 6335
2 34292 1 6335
2 34293 1 6335
2 34294 1 6335
2 34295 1 6335
2 34296 1 6335
2 34297 1 6336
2 34298 1 6336
2 34299 1 6339
2 34300 1 6339
2 34301 1 6350
2 34302 1 6350
2 34303 1 6350
2 34304 1 6350
2 34305 1 6351
2 34306 1 6351
2 34307 1 6351
2 34308 1 6351
2 34309 1 6351
2 34310 1 6351
2 34311 1 6351
2 34312 1 6351
2 34313 1 6351
2 34314 1 6351
2 34315 1 6353
2 34316 1 6353
2 34317 1 6353
2 34318 1 6354
2 34319 1 6354
2 34320 1 6354
2 34321 1 6354
2 34322 1 6354
2 34323 1 6354
2 34324 1 6354
2 34325 1 6354
2 34326 1 6354
2 34327 1 6354
2 34328 1 6354
2 34329 1 6354
2 34330 1 6354
2 34331 1 6354
2 34332 1 6354
2 34333 1 6354
2 34334 1 6354
2 34335 1 6354
2 34336 1 6354
2 34337 1 6354
2 34338 1 6354
2 34339 1 6354
2 34340 1 6360
2 34341 1 6360
2 34342 1 6371
2 34343 1 6371
2 34344 1 6372
2 34345 1 6372
2 34346 1 6374
2 34347 1 6374
2 34348 1 6374
2 34349 1 6374
2 34350 1 6374
2 34351 1 6374
2 34352 1 6375
2 34353 1 6375
2 34354 1 6379
2 34355 1 6379
2 34356 1 6399
2 34357 1 6399
2 34358 1 6399
2 34359 1 6399
2 34360 1 6449
2 34361 1 6449
2 34362 1 6449
2 34363 1 6449
2 34364 1 6450
2 34365 1 6450
2 34366 1 6467
2 34367 1 6467
2 34368 1 6477
2 34369 1 6477
2 34370 1 6477
2 34371 1 6477
2 34372 1 6478
2 34373 1 6478
2 34374 1 6478
2 34375 1 6479
2 34376 1 6479
2 34377 1 6488
2 34378 1 6488
2 34379 1 6489
2 34380 1 6489
2 34381 1 6497
2 34382 1 6497
2 34383 1 6500
2 34384 1 6500
2 34385 1 6512
2 34386 1 6512
2 34387 1 6520
2 34388 1 6520
2 34389 1 6520
2 34390 1 6520
2 34391 1 6520
2 34392 1 6520
2 34393 1 6520
2 34394 1 6520
2 34395 1 6521
2 34396 1 6521
2 34397 1 6530
2 34398 1 6530
2 34399 1 6553
2 34400 1 6553
2 34401 1 6553
2 34402 1 6553
2 34403 1 6553
2 34404 1 6554
2 34405 1 6554
2 34406 1 6555
2 34407 1 6555
2 34408 1 6558
2 34409 1 6558
2 34410 1 6558
2 34411 1 6561
2 34412 1 6561
2 34413 1 6578
2 34414 1 6578
2 34415 1 6578
2 34416 1 6578
2 34417 1 6578
2 34418 1 6578
2 34419 1 6586
2 34420 1 6586
2 34421 1 6586
2 34422 1 6586
2 34423 1 6586
2 34424 1 6586
2 34425 1 6586
2 34426 1 6586
2 34427 1 6586
2 34428 1 6600
2 34429 1 6600
2 34430 1 6600
2 34431 1 6601
2 34432 1 6601
2 34433 1 6602
2 34434 1 6602
2 34435 1 6605
2 34436 1 6605
2 34437 1 6605
2 34438 1 6605
2 34439 1 6605
2 34440 1 6608
2 34441 1 6608
2 34442 1 6609
2 34443 1 6609
2 34444 1 6610
2 34445 1 6610
2 34446 1 6614
2 34447 1 6614
2 34448 1 6614
2 34449 1 6614
2 34450 1 6614
2 34451 1 6617
2 34452 1 6617
2 34453 1 6617
2 34454 1 6617
2 34455 1 6617
2 34456 1 6617
2 34457 1 6617
2 34458 1 6621
2 34459 1 6621
2 34460 1 6621
2 34461 1 6621
2 34462 1 6621
2 34463 1 6621
2 34464 1 6621
2 34465 1 6621
2 34466 1 6621
2 34467 1 6621
2 34468 1 6621
2 34469 1 6622
2 34470 1 6622
2 34471 1 6633
2 34472 1 6633
2 34473 1 6634
2 34474 1 6634
2 34475 1 6634
2 34476 1 6634
2 34477 1 6634
2 34478 1 6656
2 34479 1 6656
2 34480 1 6656
2 34481 1 6660
2 34482 1 6660
2 34483 1 6660
2 34484 1 6660
2 34485 1 6661
2 34486 1 6661
2 34487 1 6661
2 34488 1 6662
2 34489 1 6662
2 34490 1 6662
2 34491 1 6672
2 34492 1 6672
2 34493 1 6672
2 34494 1 6673
2 34495 1 6673
2 34496 1 6674
2 34497 1 6674
2 34498 1 6693
2 34499 1 6693
2 34500 1 6693
2 34501 1 6693
2 34502 1 6694
2 34503 1 6694
2 34504 1 6694
2 34505 1 6694
2 34506 1 6701
2 34507 1 6701
2 34508 1 6701
2 34509 1 6701
2 34510 1 6708
2 34511 1 6708
2 34512 1 6708
2 34513 1 6708
2 34514 1 6708
2 34515 1 6708
2 34516 1 6708
2 34517 1 6709
2 34518 1 6709
2 34519 1 6711
2 34520 1 6711
2 34521 1 6711
2 34522 1 6712
2 34523 1 6712
2 34524 1 6722
2 34525 1 6722
2 34526 1 6723
2 34527 1 6723
2 34528 1 6723
2 34529 1 6723
2 34530 1 6723
2 34531 1 6734
2 34532 1 6734
2 34533 1 6734
2 34534 1 6739
2 34535 1 6739
2 34536 1 6740
2 34537 1 6740
2 34538 1 6750
2 34539 1 6750
2 34540 1 6750
2 34541 1 6750
2 34542 1 6750
2 34543 1 6754
2 34544 1 6754
2 34545 1 6757
2 34546 1 6757
2 34547 1 6757
2 34548 1 6758
2 34549 1 6758
2 34550 1 6764
2 34551 1 6764
2 34552 1 6764
2 34553 1 6779
2 34554 1 6779
2 34555 1 6779
2 34556 1 6787
2 34557 1 6787
2 34558 1 6787
2 34559 1 6787
2 34560 1 6787
2 34561 1 6787
2 34562 1 6787
2 34563 1 6787
2 34564 1 6787
2 34565 1 6788
2 34566 1 6788
2 34567 1 6788
2 34568 1 6788
2 34569 1 6788
2 34570 1 6788
2 34571 1 6801
2 34572 1 6801
2 34573 1 6801
2 34574 1 6811
2 34575 1 6811
2 34576 1 6811
2 34577 1 6825
2 34578 1 6825
2 34579 1 6825
2 34580 1 6825
2 34581 1 6825
2 34582 1 6826
2 34583 1 6826
2 34584 1 6826
2 34585 1 6826
2 34586 1 6826
2 34587 1 6826
2 34588 1 6842
2 34589 1 6842
2 34590 1 6842
2 34591 1 6842
2 34592 1 6842
2 34593 1 6853
2 34594 1 6853
2 34595 1 6857
2 34596 1 6857
2 34597 1 6857
2 34598 1 6872
2 34599 1 6872
2 34600 1 6872
2 34601 1 6875
2 34602 1 6875
2 34603 1 6875
2 34604 1 6881
2 34605 1 6881
2 34606 1 6881
2 34607 1 6881
2 34608 1 6881
2 34609 1 6891
2 34610 1 6891
2 34611 1 6891
2 34612 1 6891
2 34613 1 6891
2 34614 1 6891
2 34615 1 6893
2 34616 1 6893
2 34617 1 6893
2 34618 1 6902
2 34619 1 6902
2 34620 1 6902
2 34621 1 6902
2 34622 1 6902
2 34623 1 6903
2 34624 1 6903
2 34625 1 6928
2 34626 1 6928
2 34627 1 6936
2 34628 1 6936
2 34629 1 6936
2 34630 1 6936
2 34631 1 6936
2 34632 1 6936
2 34633 1 6945
2 34634 1 6945
2 34635 1 6945
2 34636 1 6986
2 34637 1 6986
2 34638 1 6986
2 34639 1 6986
2 34640 1 6986
2 34641 1 6986
2 34642 1 7024
2 34643 1 7024
2 34644 1 7024
2 34645 1 7024
2 34646 1 7025
2 34647 1 7025
2 34648 1 7025
2 34649 1 7026
2 34650 1 7026
2 34651 1 7037
2 34652 1 7037
2 34653 1 7037
2 34654 1 7044
2 34655 1 7044
2 34656 1 7044
2 34657 1 7055
2 34658 1 7055
2 34659 1 7056
2 34660 1 7056
2 34661 1 7056
2 34662 1 7081
2 34663 1 7081
2 34664 1 7081
2 34665 1 7081
2 34666 1 7084
2 34667 1 7084
2 34668 1 7087
2 34669 1 7087
2 34670 1 7117
2 34671 1 7117
2 34672 1 7117
2 34673 1 7117
2 34674 1 7117
2 34675 1 7118
2 34676 1 7118
2 34677 1 7118
2 34678 1 7118
2 34679 1 7118
2 34680 1 7118
2 34681 1 7118
2 34682 1 7118
2 34683 1 7118
2 34684 1 7118
2 34685 1 7121
2 34686 1 7121
2 34687 1 7121
2 34688 1 7122
2 34689 1 7122
2 34690 1 7122
2 34691 1 7122
2 34692 1 7122
2 34693 1 7122
2 34694 1 7123
2 34695 1 7123
2 34696 1 7131
2 34697 1 7131
2 34698 1 7140
2 34699 1 7140
2 34700 1 7140
2 34701 1 7144
2 34702 1 7144
2 34703 1 7154
2 34704 1 7154
2 34705 1 7154
2 34706 1 7159
2 34707 1 7159
2 34708 1 7168
2 34709 1 7168
2 34710 1 7168
2 34711 1 7168
2 34712 1 7169
2 34713 1 7169
2 34714 1 7171
2 34715 1 7171
2 34716 1 7171
2 34717 1 7178
2 34718 1 7178
2 34719 1 7186
2 34720 1 7186
2 34721 1 7200
2 34722 1 7200
2 34723 1 7200
2 34724 1 7231
2 34725 1 7231
2 34726 1 7239
2 34727 1 7239
2 34728 1 7247
2 34729 1 7247
2 34730 1 7249
2 34731 1 7249
2 34732 1 7255
2 34733 1 7255
2 34734 1 7255
2 34735 1 7263
2 34736 1 7263
2 34737 1 7279
2 34738 1 7279
2 34739 1 7279
2 34740 1 7279
2 34741 1 7279
2 34742 1 7281
2 34743 1 7281
2 34744 1 7287
2 34745 1 7287
2 34746 1 7314
2 34747 1 7314
2 34748 1 7315
2 34749 1 7315
2 34750 1 7322
2 34751 1 7322
2 34752 1 7322
2 34753 1 7322
2 34754 1 7323
2 34755 1 7323
2 34756 1 7326
2 34757 1 7326
2 34758 1 7333
2 34759 1 7333
2 34760 1 7354
2 34761 1 7354
2 34762 1 7355
2 34763 1 7355
2 34764 1 7355
2 34765 1 7378
2 34766 1 7378
2 34767 1 7378
2 34768 1 7379
2 34769 1 7379
2 34770 1 7386
2 34771 1 7386
2 34772 1 7414
2 34773 1 7414
2 34774 1 7417
2 34775 1 7417
2 34776 1 7435
2 34777 1 7435
2 34778 1 7435
2 34779 1 7435
2 34780 1 7444
2 34781 1 7444
2 34782 1 7444
2 34783 1 7444
2 34784 1 7444
2 34785 1 7444
2 34786 1 7444
2 34787 1 7444
2 34788 1 7444
2 34789 1 7444
2 34790 1 7444
2 34791 1 7447
2 34792 1 7447
2 34793 1 7450
2 34794 1 7450
2 34795 1 7450
2 34796 1 7450
2 34797 1 7453
2 34798 1 7453
2 34799 1 7453
2 34800 1 7454
2 34801 1 7454
2 34802 1 7474
2 34803 1 7474
2 34804 1 7474
2 34805 1 7474
2 34806 1 7474
2 34807 1 7474
2 34808 1 7474
2 34809 1 7474
2 34810 1 7474
2 34811 1 7474
2 34812 1 7489
2 34813 1 7489
2 34814 1 7489
2 34815 1 7490
2 34816 1 7490
2 34817 1 7499
2 34818 1 7499
2 34819 1 7499
2 34820 1 7499
2 34821 1 7502
2 34822 1 7502
2 34823 1 7516
2 34824 1 7516
2 34825 1 7530
2 34826 1 7530
2 34827 1 7530
2 34828 1 7531
2 34829 1 7531
2 34830 1 7542
2 34831 1 7542
2 34832 1 7556
2 34833 1 7556
2 34834 1 7559
2 34835 1 7559
2 34836 1 7568
2 34837 1 7568
2 34838 1 7569
2 34839 1 7569
2 34840 1 7577
2 34841 1 7577
2 34842 1 7579
2 34843 1 7579
2 34844 1 7586
2 34845 1 7586
2 34846 1 7617
2 34847 1 7617
2 34848 1 7630
2 34849 1 7630
2 34850 1 7630
2 34851 1 7631
2 34852 1 7631
2 34853 1 7643
2 34854 1 7643
2 34855 1 7643
2 34856 1 7643
2 34857 1 7643
2 34858 1 7643
2 34859 1 7643
2 34860 1 7644
2 34861 1 7644
2 34862 1 7644
2 34863 1 7644
2 34864 1 7644
2 34865 1 7644
2 34866 1 7644
2 34867 1 7644
2 34868 1 7661
2 34869 1 7661
2 34870 1 7661
2 34871 1 7661
2 34872 1 7662
2 34873 1 7662
2 34874 1 7666
2 34875 1 7666
2 34876 1 7666
2 34877 1 7666
2 34878 1 7666
2 34879 1 7666
2 34880 1 7666
2 34881 1 7666
2 34882 1 7666
2 34883 1 7666
2 34884 1 7666
2 34885 1 7666
2 34886 1 7666
2 34887 1 7667
2 34888 1 7667
2 34889 1 7667
2 34890 1 7667
2 34891 1 7667
2 34892 1 7667
2 34893 1 7673
2 34894 1 7673
2 34895 1 7674
2 34896 1 7674
2 34897 1 7682
2 34898 1 7682
2 34899 1 7684
2 34900 1 7684
2 34901 1 7684
2 34902 1 7684
2 34903 1 7684
2 34904 1 7689
2 34905 1 7689
2 34906 1 7703
2 34907 1 7703
2 34908 1 7707
2 34909 1 7707
2 34910 1 7708
2 34911 1 7708
2 34912 1 7708
2 34913 1 7708
2 34914 1 7708
2 34915 1 7723
2 34916 1 7723
2 34917 1 7723
2 34918 1 7723
2 34919 1 7723
2 34920 1 7723
2 34921 1 7723
2 34922 1 7723
2 34923 1 7726
2 34924 1 7726
2 34925 1 7727
2 34926 1 7727
2 34927 1 7734
2 34928 1 7734
2 34929 1 7734
2 34930 1 7734
2 34931 1 7734
2 34932 1 7734
2 34933 1 7734
2 34934 1 7734
2 34935 1 7734
2 34936 1 7734
2 34937 1 7734
2 34938 1 7734
2 34939 1 7734
2 34940 1 7734
2 34941 1 7734
2 34942 1 7734
2 34943 1 7734
2 34944 1 7734
2 34945 1 7734
2 34946 1 7734
2 34947 1 7737
2 34948 1 7737
2 34949 1 7737
2 34950 1 7737
2 34951 1 7737
2 34952 1 7737
2 34953 1 7737
2 34954 1 7737
2 34955 1 7737
2 34956 1 7737
2 34957 1 7737
2 34958 1 7739
2 34959 1 7739
2 34960 1 7739
2 34961 1 7739
2 34962 1 7739
2 34963 1 7740
2 34964 1 7740
2 34965 1 7756
2 34966 1 7756
2 34967 1 7756
2 34968 1 7764
2 34969 1 7764
2 34970 1 7768
2 34971 1 7768
2 34972 1 7768
2 34973 1 7768
2 34974 1 7768
2 34975 1 7771
2 34976 1 7771
2 34977 1 7771
2 34978 1 7771
2 34979 1 7771
2 34980 1 7771
2 34981 1 7771
2 34982 1 7771
2 34983 1 7771
2 34984 1 7771
2 34985 1 7771
2 34986 1 7771
2 34987 1 7771
2 34988 1 7771
2 34989 1 7773
2 34990 1 7773
2 34991 1 7774
2 34992 1 7774
2 34993 1 7777
2 34994 1 7777
2 34995 1 7777
2 34996 1 7777
2 34997 1 7777
2 34998 1 7777
2 34999 1 7783
2 35000 1 7783
2 35001 1 7786
2 35002 1 7786
2 35003 1 7786
2 35004 1 7786
2 35005 1 7821
2 35006 1 7821
2 35007 1 7821
2 35008 1 7821
2 35009 1 7822
2 35010 1 7822
2 35011 1 7822
2 35012 1 7822
2 35013 1 7822
2 35014 1 7822
2 35015 1 7825
2 35016 1 7825
2 35017 1 7826
2 35018 1 7826
2 35019 1 7828
2 35020 1 7828
2 35021 1 7828
2 35022 1 7828
2 35023 1 7863
2 35024 1 7863
2 35025 1 7876
2 35026 1 7876
2 35027 1 7876
2 35028 1 7876
2 35029 1 7876
2 35030 1 7876
2 35031 1 7876
2 35032 1 7878
2 35033 1 7878
2 35034 1 7878
2 35035 1 7880
2 35036 1 7880
2 35037 1 7897
2 35038 1 7897
2 35039 1 7909
2 35040 1 7909
2 35041 1 7921
2 35042 1 7921
2 35043 1 7930
2 35044 1 7930
2 35045 1 7930
2 35046 1 7938
2 35047 1 7938
2 35048 1 7938
2 35049 1 7938
2 35050 1 7948
2 35051 1 7948
2 35052 1 7949
2 35053 1 7949
2 35054 1 7949
2 35055 1 7949
2 35056 1 7949
2 35057 1 7949
2 35058 1 7949
2 35059 1 7949
2 35060 1 7949
2 35061 1 7949
2 35062 1 7949
2 35063 1 7949
2 35064 1 7957
2 35065 1 7957
2 35066 1 7958
2 35067 1 7958
2 35068 1 7958
2 35069 1 7967
2 35070 1 7967
2 35071 1 7976
2 35072 1 7976
2 35073 1 7981
2 35074 1 7981
2 35075 1 7981
2 35076 1 8003
2 35077 1 8003
2 35078 1 8007
2 35079 1 8007
2 35080 1 8007
2 35081 1 8010
2 35082 1 8010
2 35083 1 8010
2 35084 1 8010
2 35085 1 8010
2 35086 1 8010
2 35087 1 8010
2 35088 1 8010
2 35089 1 8010
2 35090 1 8010
2 35091 1 8010
2 35092 1 8017
2 35093 1 8017
2 35094 1 8017
2 35095 1 8017
2 35096 1 8018
2 35097 1 8018
2 35098 1 8025
2 35099 1 8025
2 35100 1 8026
2 35101 1 8026
2 35102 1 8026
2 35103 1 8027
2 35104 1 8027
2 35105 1 8033
2 35106 1 8033
2 35107 1 8033
2 35108 1 8033
2 35109 1 8033
2 35110 1 8036
2 35111 1 8036
2 35112 1 8058
2 35113 1 8058
2 35114 1 8058
2 35115 1 8058
2 35116 1 8059
2 35117 1 8059
2 35118 1 8059
2 35119 1 8059
2 35120 1 8063
2 35121 1 8063
2 35122 1 8068
2 35123 1 8068
2 35124 1 8068
2 35125 1 8073
2 35126 1 8073
2 35127 1 8073
2 35128 1 8073
2 35129 1 8073
2 35130 1 8073
2 35131 1 8073
2 35132 1 8073
2 35133 1 8073
2 35134 1 8074
2 35135 1 8074
2 35136 1 8074
2 35137 1 8076
2 35138 1 8076
2 35139 1 8080
2 35140 1 8080
2 35141 1 8121
2 35142 1 8121
2 35143 1 8121
2 35144 1 8121
2 35145 1 8121
2 35146 1 8121
2 35147 1 8122
2 35148 1 8122
2 35149 1 8125
2 35150 1 8125
2 35151 1 8131
2 35152 1 8131
2 35153 1 8138
2 35154 1 8138
2 35155 1 8138
2 35156 1 8147
2 35157 1 8147
2 35158 1 8148
2 35159 1 8148
2 35160 1 8168
2 35161 1 8168
2 35162 1 8168
2 35163 1 8168
2 35164 1 8168
2 35165 1 8168
2 35166 1 8173
2 35167 1 8173
2 35168 1 8181
2 35169 1 8181
2 35170 1 8181
2 35171 1 8181
2 35172 1 8181
2 35173 1 8194
2 35174 1 8194
2 35175 1 8194
2 35176 1 8194
2 35177 1 8194
2 35178 1 8198
2 35179 1 8198
2 35180 1 8198
2 35181 1 8201
2 35182 1 8201
2 35183 1 8202
2 35184 1 8202
2 35185 1 8222
2 35186 1 8222
2 35187 1 8222
2 35188 1 8235
2 35189 1 8235
2 35190 1 8249
2 35191 1 8249
2 35192 1 8271
2 35193 1 8271
2 35194 1 8289
2 35195 1 8289
2 35196 1 8290
2 35197 1 8290
2 35198 1 8302
2 35199 1 8302
2 35200 1 8333
2 35201 1 8333
2 35202 1 8334
2 35203 1 8334
2 35204 1 8334
2 35205 1 8334
2 35206 1 8335
2 35207 1 8335
2 35208 1 8337
2 35209 1 8337
2 35210 1 8337
2 35211 1 8337
2 35212 1 8337
2 35213 1 8337
2 35214 1 8337
2 35215 1 8342
2 35216 1 8342
2 35217 1 8359
2 35218 1 8359
2 35219 1 8362
2 35220 1 8362
2 35221 1 8362
2 35222 1 8367
2 35223 1 8367
2 35224 1 8376
2 35225 1 8376
2 35226 1 8377
2 35227 1 8377
2 35228 1 8380
2 35229 1 8380
2 35230 1 8381
2 35231 1 8381
2 35232 1 8391
2 35233 1 8391
2 35234 1 8391
2 35235 1 8393
2 35236 1 8393
2 35237 1 8402
2 35238 1 8402
2 35239 1 8402
2 35240 1 8403
2 35241 1 8403
2 35242 1 8404
2 35243 1 8404
2 35244 1 8408
2 35245 1 8408
2 35246 1 8409
2 35247 1 8409
2 35248 1 8409
2 35249 1 8410
2 35250 1 8410
2 35251 1 8424
2 35252 1 8424
2 35253 1 8439
2 35254 1 8439
2 35255 1 8440
2 35256 1 8440
2 35257 1 8440
2 35258 1 8440
2 35259 1 8440
2 35260 1 8440
2 35261 1 8441
2 35262 1 8441
2 35263 1 8441
2 35264 1 8441
2 35265 1 8444
2 35266 1 8444
2 35267 1 8444
2 35268 1 8445
2 35269 1 8445
2 35270 1 8446
2 35271 1 8446
2 35272 1 8448
2 35273 1 8448
2 35274 1 8448
2 35275 1 8448
2 35276 1 8460
2 35277 1 8460
2 35278 1 8460
2 35279 1 8461
2 35280 1 8461
2 35281 1 8461
2 35282 1 8462
2 35283 1 8462
2 35284 1 8462
2 35285 1 8462
2 35286 1 8462
2 35287 1 8472
2 35288 1 8472
2 35289 1 8472
2 35290 1 8472
2 35291 1 8472
2 35292 1 8472
2 35293 1 8473
2 35294 1 8473
2 35295 1 8473
2 35296 1 8473
2 35297 1 8473
2 35298 1 8473
2 35299 1 8477
2 35300 1 8477
2 35301 1 8477
2 35302 1 8478
2 35303 1 8478
2 35304 1 8478
2 35305 1 8478
2 35306 1 8478
2 35307 1 8488
2 35308 1 8488
2 35309 1 8488
2 35310 1 8488
2 35311 1 8505
2 35312 1 8505
2 35313 1 8518
2 35314 1 8518
2 35315 1 8518
2 35316 1 8544
2 35317 1 8544
2 35318 1 8565
2 35319 1 8565
2 35320 1 8565
2 35321 1 8565
2 35322 1 8568
2 35323 1 8568
2 35324 1 8568
2 35325 1 8578
2 35326 1 8578
2 35327 1 8584
2 35328 1 8584
2 35329 1 8587
2 35330 1 8587
2 35331 1 8596
2 35332 1 8596
2 35333 1 8596
2 35334 1 8596
2 35335 1 8596
2 35336 1 8604
2 35337 1 8604
2 35338 1 8607
2 35339 1 8607
2 35340 1 8607
2 35341 1 8611
2 35342 1 8611
2 35343 1 8611
2 35344 1 8635
2 35345 1 8635
2 35346 1 8665
2 35347 1 8665
2 35348 1 8665
2 35349 1 8694
2 35350 1 8694
2 35351 1 8695
2 35352 1 8695
2 35353 1 8695
2 35354 1 8695
2 35355 1 8695
2 35356 1 8695
2 35357 1 8695
2 35358 1 8710
2 35359 1 8710
2 35360 1 8710
2 35361 1 8723
2 35362 1 8723
2 35363 1 8729
2 35364 1 8729
2 35365 1 8734
2 35366 1 8734
2 35367 1 8738
2 35368 1 8738
2 35369 1 8744
2 35370 1 8744
2 35371 1 8756
2 35372 1 8756
2 35373 1 8762
2 35374 1 8762
2 35375 1 8767
2 35376 1 8767
2 35377 1 8770
2 35378 1 8770
2 35379 1 8770
2 35380 1 8771
2 35381 1 8771
2 35382 1 8818
2 35383 1 8818
2 35384 1 8819
2 35385 1 8819
2 35386 1 8819
2 35387 1 8819
2 35388 1 8842
2 35389 1 8842
2 35390 1 8849
2 35391 1 8849
2 35392 1 8876
2 35393 1 8876
2 35394 1 8882
2 35395 1 8882
2 35396 1 8895
2 35397 1 8895
2 35398 1 8895
2 35399 1 8895
2 35400 1 8896
2 35401 1 8896
2 35402 1 8898
2 35403 1 8898
2 35404 1 8898
2 35405 1 8899
2 35406 1 8899
2 35407 1 8916
2 35408 1 8916
2 35409 1 8917
2 35410 1 8917
2 35411 1 8938
2 35412 1 8938
2 35413 1 8938
2 35414 1 8938
2 35415 1 8940
2 35416 1 8940
2 35417 1 8940
2 35418 1 8940
2 35419 1 8940
2 35420 1 8940
2 35421 1 8941
2 35422 1 8941
2 35423 1 8941
2 35424 1 8953
2 35425 1 8953
2 35426 1 8953
2 35427 1 8954
2 35428 1 8954
2 35429 1 8954
2 35430 1 8954
2 35431 1 8955
2 35432 1 8955
2 35433 1 8958
2 35434 1 8958
2 35435 1 8958
2 35436 1 8977
2 35437 1 8977
2 35438 1 8977
2 35439 1 8982
2 35440 1 8982
2 35441 1 8984
2 35442 1 8984
2 35443 1 8984
2 35444 1 8984
2 35445 1 8988
2 35446 1 8988
2 35447 1 8988
2 35448 1 8997
2 35449 1 8997
2 35450 1 9000
2 35451 1 9000
2 35452 1 9007
2 35453 1 9007
2 35454 1 9007
2 35455 1 9014
2 35456 1 9014
2 35457 1 9014
2 35458 1 9014
2 35459 1 9015
2 35460 1 9015
2 35461 1 9023
2 35462 1 9023
2 35463 1 9023
2 35464 1 9025
2 35465 1 9025
2 35466 1 9025
2 35467 1 9028
2 35468 1 9028
2 35469 1 9028
2 35470 1 9028
2 35471 1 9028
2 35472 1 9028
2 35473 1 9029
2 35474 1 9029
2 35475 1 9030
2 35476 1 9030
2 35477 1 9064
2 35478 1 9064
2 35479 1 9065
2 35480 1 9065
2 35481 1 9077
2 35482 1 9077
2 35483 1 9077
2 35484 1 9081
2 35485 1 9081
2 35486 1 9081
2 35487 1 9081
2 35488 1 9081
2 35489 1 9082
2 35490 1 9082
2 35491 1 9086
2 35492 1 9086
2 35493 1 9086
2 35494 1 9087
2 35495 1 9087
2 35496 1 9093
2 35497 1 9093
2 35498 1 9118
2 35499 1 9118
2 35500 1 9118
2 35501 1 9129
2 35502 1 9129
2 35503 1 9131
2 35504 1 9131
2 35505 1 9134
2 35506 1 9134
2 35507 1 9134
2 35508 1 9134
2 35509 1 9134
2 35510 1 9134
2 35511 1 9137
2 35512 1 9137
2 35513 1 9137
2 35514 1 9137
2 35515 1 9139
2 35516 1 9139
2 35517 1 9139
2 35518 1 9139
2 35519 1 9141
2 35520 1 9141
2 35521 1 9188
2 35522 1 9188
2 35523 1 9189
2 35524 1 9189
2 35525 1 9193
2 35526 1 9193
2 35527 1 9193
2 35528 1 9196
2 35529 1 9196
2 35530 1 9214
2 35531 1 9214
2 35532 1 9214
2 35533 1 9226
2 35534 1 9226
2 35535 1 9226
2 35536 1 9226
2 35537 1 9226
2 35538 1 9236
2 35539 1 9236
2 35540 1 9236
2 35541 1 9236
2 35542 1 9237
2 35543 1 9237
2 35544 1 9237
2 35545 1 9237
2 35546 1 9237
2 35547 1 9245
2 35548 1 9245
2 35549 1 9245
2 35550 1 9246
2 35551 1 9246
2 35552 1 9246
2 35553 1 9246
2 35554 1 9246
2 35555 1 9247
2 35556 1 9247
2 35557 1 9255
2 35558 1 9255
2 35559 1 9258
2 35560 1 9258
2 35561 1 9261
2 35562 1 9261
2 35563 1 9261
2 35564 1 9261
2 35565 1 9261
2 35566 1 9261
2 35567 1 9284
2 35568 1 9284
2 35569 1 9323
2 35570 1 9323
2 35571 1 9332
2 35572 1 9332
2 35573 1 9333
2 35574 1 9333
2 35575 1 9333
2 35576 1 9333
2 35577 1 9343
2 35578 1 9343
2 35579 1 9363
2 35580 1 9363
2 35581 1 9368
2 35582 1 9368
2 35583 1 9378
2 35584 1 9378
2 35585 1 9383
2 35586 1 9383
2 35587 1 9383
2 35588 1 9383
2 35589 1 9383
2 35590 1 9383
2 35591 1 9383
2 35592 1 9397
2 35593 1 9397
2 35594 1 9397
2 35595 1 9397
2 35596 1 9397
2 35597 1 9402
2 35598 1 9402
2 35599 1 9405
2 35600 1 9405
2 35601 1 9405
2 35602 1 9428
2 35603 1 9428
2 35604 1 9429
2 35605 1 9429
2 35606 1 9437
2 35607 1 9437
2 35608 1 9437
2 35609 1 9446
2 35610 1 9446
2 35611 1 9455
2 35612 1 9455
2 35613 1 9455
2 35614 1 9455
2 35615 1 9456
2 35616 1 9456
2 35617 1 9466
2 35618 1 9466
2 35619 1 9466
2 35620 1 9467
2 35621 1 9467
2 35622 1 9467
2 35623 1 9487
2 35624 1 9487
2 35625 1 9520
2 35626 1 9520
2 35627 1 9529
2 35628 1 9529
2 35629 1 9529
2 35630 1 9530
2 35631 1 9530
2 35632 1 9530
2 35633 1 9533
2 35634 1 9533
2 35635 1 9533
2 35636 1 9534
2 35637 1 9534
2 35638 1 9561
2 35639 1 9561
2 35640 1 9571
2 35641 1 9571
2 35642 1 9571
2 35643 1 9571
2 35644 1 9571
2 35645 1 9571
2 35646 1 9588
2 35647 1 9588
2 35648 1 9591
2 35649 1 9591
2 35650 1 9603
2 35651 1 9603
2 35652 1 9603
2 35653 1 9603
2 35654 1 9613
2 35655 1 9613
2 35656 1 9622
2 35657 1 9622
2 35658 1 9623
2 35659 1 9623
2 35660 1 9645
2 35661 1 9645
2 35662 1 9678
2 35663 1 9678
2 35664 1 9678
2 35665 1 9678
2 35666 1 9678
2 35667 1 9679
2 35668 1 9679
2 35669 1 9686
2 35670 1 9686
2 35671 1 9694
2 35672 1 9694
2 35673 1 9694
2 35674 1 9703
2 35675 1 9703
2 35676 1 9703
2 35677 1 9703
2 35678 1 9703
2 35679 1 9703
2 35680 1 9705
2 35681 1 9705
2 35682 1 9706
2 35683 1 9706
2 35684 1 9715
2 35685 1 9715
2 35686 1 9718
2 35687 1 9718
2 35688 1 9718
2 35689 1 9718
2 35690 1 9718
2 35691 1 9719
2 35692 1 9719
2 35693 1 9724
2 35694 1 9724
2 35695 1 9737
2 35696 1 9737
2 35697 1 9752
2 35698 1 9752
2 35699 1 9752
2 35700 1 9752
2 35701 1 9756
2 35702 1 9756
2 35703 1 9758
2 35704 1 9758
2 35705 1 9761
2 35706 1 9761
2 35707 1 9761
2 35708 1 9772
2 35709 1 9772
2 35710 1 9772
2 35711 1 9773
2 35712 1 9773
2 35713 1 9773
2 35714 1 9775
2 35715 1 9775
2 35716 1 9808
2 35717 1 9808
2 35718 1 9808
2 35719 1 9811
2 35720 1 9811
2 35721 1 9811
2 35722 1 9811
2 35723 1 9811
2 35724 1 9815
2 35725 1 9815
2 35726 1 9823
2 35727 1 9823
2 35728 1 9834
2 35729 1 9834
2 35730 1 9850
2 35731 1 9850
2 35732 1 9883
2 35733 1 9883
2 35734 1 9883
2 35735 1 9883
2 35736 1 9883
2 35737 1 9883
2 35738 1 9885
2 35739 1 9885
2 35740 1 9885
2 35741 1 9887
2 35742 1 9887
2 35743 1 9925
2 35744 1 9925
2 35745 1 9925
2 35746 1 9925
2 35747 1 9925
2 35748 1 9927
2 35749 1 9927
2 35750 1 9933
2 35751 1 9933
2 35752 1 9933
2 35753 1 9951
2 35754 1 9951
2 35755 1 9951
2 35756 1 9951
2 35757 1 9951
2 35758 1 9991
2 35759 1 9991
2 35760 1 9991
2 35761 1 9991
2 35762 1 9991
2 35763 1 10003
2 35764 1 10003
2 35765 1 10003
2 35766 1 10011
2 35767 1 10011
2 35768 1 10016
2 35769 1 10016
2 35770 1 10016
2 35771 1 10021
2 35772 1 10021
2 35773 1 10026
2 35774 1 10026
2 35775 1 10030
2 35776 1 10030
2 35777 1 10095
2 35778 1 10095
2 35779 1 10095
2 35780 1 10095
2 35781 1 10114
2 35782 1 10114
2 35783 1 10117
2 35784 1 10117
2 35785 1 10140
2 35786 1 10140
2 35787 1 10140
2 35788 1 10147
2 35789 1 10147
2 35790 1 10157
2 35791 1 10157
2 35792 1 10200
2 35793 1 10200
2 35794 1 10201
2 35795 1 10201
2 35796 1 10201
2 35797 1 10201
2 35798 1 10211
2 35799 1 10211
2 35800 1 10214
2 35801 1 10214
2 35802 1 10214
2 35803 1 10221
2 35804 1 10221
2 35805 1 10222
2 35806 1 10222
2 35807 1 10226
2 35808 1 10226
2 35809 1 10227
2 35810 1 10227
2 35811 1 10227
2 35812 1 10227
2 35813 1 10240
2 35814 1 10240
2 35815 1 10240
2 35816 1 10240
2 35817 1 10241
2 35818 1 10241
2 35819 1 10244
2 35820 1 10244
2 35821 1 10277
2 35822 1 10277
2 35823 1 10281
2 35824 1 10281
2 35825 1 10281
2 35826 1 10288
2 35827 1 10288
2 35828 1 10295
2 35829 1 10295
2 35830 1 10304
2 35831 1 10304
2 35832 1 10304
2 35833 1 10305
2 35834 1 10305
2 35835 1 10305
2 35836 1 10315
2 35837 1 10315
2 35838 1 10317
2 35839 1 10317
2 35840 1 10321
2 35841 1 10321
2 35842 1 10321
2 35843 1 10324
2 35844 1 10324
2 35845 1 10324
2 35846 1 10325
2 35847 1 10325
2 35848 1 10342
2 35849 1 10342
2 35850 1 10355
2 35851 1 10355
2 35852 1 10355
2 35853 1 10355
2 35854 1 10355
2 35855 1 10376
2 35856 1 10376
2 35857 1 10376
2 35858 1 10384
2 35859 1 10384
2 35860 1 10384
2 35861 1 10384
2 35862 1 10386
2 35863 1 10386
2 35864 1 10402
2 35865 1 10402
2 35866 1 10415
2 35867 1 10415
2 35868 1 10423
2 35869 1 10423
2 35870 1 10443
2 35871 1 10443
2 35872 1 10445
2 35873 1 10445
2 35874 1 10448
2 35875 1 10448
2 35876 1 10454
2 35877 1 10454
2 35878 1 10455
2 35879 1 10455
2 35880 1 10455
2 35881 1 10464
2 35882 1 10464
2 35883 1 10465
2 35884 1 10465
2 35885 1 10466
2 35886 1 10466
2 35887 1 10497
2 35888 1 10497
2 35889 1 10500
2 35890 1 10500
2 35891 1 10508
2 35892 1 10508
2 35893 1 10508
2 35894 1 10509
2 35895 1 10509
2 35896 1 10517
2 35897 1 10517
2 35898 1 10517
2 35899 1 10517
2 35900 1 10517
2 35901 1 10517
2 35902 1 10517
2 35903 1 10518
2 35904 1 10518
2 35905 1 10518
2 35906 1 10519
2 35907 1 10519
2 35908 1 10526
2 35909 1 10526
2 35910 1 10533
2 35911 1 10533
2 35912 1 10539
2 35913 1 10539
2 35914 1 10594
2 35915 1 10594
2 35916 1 10608
2 35917 1 10608
2 35918 1 10608
2 35919 1 10608
2 35920 1 10608
2 35921 1 10631
2 35922 1 10631
2 35923 1 10632
2 35924 1 10632
2 35925 1 10670
2 35926 1 10670
2 35927 1 10673
2 35928 1 10673
2 35929 1 10700
2 35930 1 10700
2 35931 1 10701
2 35932 1 10701
2 35933 1 10711
2 35934 1 10711
2 35935 1 10712
2 35936 1 10712
2 35937 1 10749
2 35938 1 10749
2 35939 1 10752
2 35940 1 10752
2 35941 1 10753
2 35942 1 10753
2 35943 1 10766
2 35944 1 10766
2 35945 1 10783
2 35946 1 10783
2 35947 1 10791
2 35948 1 10791
2 35949 1 10794
2 35950 1 10794
2 35951 1 10795
2 35952 1 10795
2 35953 1 10796
2 35954 1 10796
2 35955 1 10837
2 35956 1 10837
2 35957 1 10838
2 35958 1 10838
2 35959 1 10852
2 35960 1 10852
2 35961 1 10852
2 35962 1 10876
2 35963 1 10876
2 35964 1 10880
2 35965 1 10880
2 35966 1 10890
2 35967 1 10890
2 35968 1 10890
2 35969 1 10890
2 35970 1 10900
2 35971 1 10900
2 35972 1 10900
2 35973 1 10907
2 35974 1 10907
2 35975 1 10910
2 35976 1 10910
2 35977 1 10913
2 35978 1 10913
2 35979 1 10921
2 35980 1 10921
2 35981 1 10953
2 35982 1 10953
2 35983 1 10975
2 35984 1 10975
2 35985 1 10998
2 35986 1 10998
2 35987 1 11000
2 35988 1 11000
2 35989 1 11002
2 35990 1 11002
2 35991 1 11008
2 35992 1 11008
2 35993 1 11026
2 35994 1 11026
2 35995 1 11026
2 35996 1 11029
2 35997 1 11029
2 35998 1 11030
2 35999 1 11030
2 36000 1 11049
2 36001 1 11049
2 36002 1 11049
2 36003 1 11049
2 36004 1 11070
2 36005 1 11070
2 36006 1 11102
2 36007 1 11102
2 36008 1 11109
2 36009 1 11109
2 36010 1 11109
2 36011 1 11109
2 36012 1 11110
2 36013 1 11110
2 36014 1 11115
2 36015 1 11115
2 36016 1 11115
2 36017 1 11115
2 36018 1 11115
2 36019 1 11115
2 36020 1 11115
2 36021 1 11115
2 36022 1 11132
2 36023 1 11132
2 36024 1 11139
2 36025 1 11139
2 36026 1 11142
2 36027 1 11142
2 36028 1 11145
2 36029 1 11145
2 36030 1 11147
2 36031 1 11147
2 36032 1 11148
2 36033 1 11148
2 36034 1 11152
2 36035 1 11152
2 36036 1 11152
2 36037 1 11152
2 36038 1 11152
2 36039 1 11152
2 36040 1 11152
2 36041 1 11154
2 36042 1 11154
2 36043 1 11155
2 36044 1 11155
2 36045 1 11164
2 36046 1 11164
2 36047 1 11164
2 36048 1 11164
2 36049 1 11164
2 36050 1 11164
2 36051 1 11169
2 36052 1 11169
2 36053 1 11188
2 36054 1 11188
2 36055 1 11188
2 36056 1 11188
2 36057 1 11188
2 36058 1 11198
2 36059 1 11198
2 36060 1 11198
2 36061 1 11205
2 36062 1 11205
2 36063 1 11205
2 36064 1 11205
2 36065 1 11206
2 36066 1 11206
2 36067 1 11207
2 36068 1 11207
2 36069 1 11207
2 36070 1 11228
2 36071 1 11228
2 36072 1 11228
2 36073 1 11234
2 36074 1 11234
2 36075 1 11234
2 36076 1 11234
2 36077 1 11234
2 36078 1 11234
2 36079 1 11236
2 36080 1 11236
2 36081 1 11243
2 36082 1 11243
2 36083 1 11243
2 36084 1 11244
2 36085 1 11244
2 36086 1 11252
2 36087 1 11252
2 36088 1 11252
2 36089 1 11252
2 36090 1 11286
2 36091 1 11286
2 36092 1 11312
2 36093 1 11312
2 36094 1 11312
2 36095 1 11312
2 36096 1 11313
2 36097 1 11313
2 36098 1 11318
2 36099 1 11318
2 36100 1 11326
2 36101 1 11326
2 36102 1 11326
2 36103 1 11330
2 36104 1 11330
2 36105 1 11335
2 36106 1 11335
2 36107 1 11337
2 36108 1 11337
2 36109 1 11340
2 36110 1 11340
2 36111 1 11340
2 36112 1 11340
2 36113 1 11340
2 36114 1 11341
2 36115 1 11341
2 36116 1 11342
2 36117 1 11342
2 36118 1 11361
2 36119 1 11361
2 36120 1 11376
2 36121 1 11376
2 36122 1 11376
2 36123 1 11376
2 36124 1 11376
2 36125 1 11378
2 36126 1 11378
2 36127 1 11379
2 36128 1 11379
2 36129 1 11381
2 36130 1 11381
2 36131 1 11381
2 36132 1 11381
2 36133 1 11381
2 36134 1 11393
2 36135 1 11393
2 36136 1 11400
2 36137 1 11400
2 36138 1 11410
2 36139 1 11410
2 36140 1 11421
2 36141 1 11421
2 36142 1 11435
2 36143 1 11435
2 36144 1 11442
2 36145 1 11442
2 36146 1 11442
2 36147 1 11442
2 36148 1 11466
2 36149 1 11466
2 36150 1 11467
2 36151 1 11467
2 36152 1 11478
2 36153 1 11478
2 36154 1 11478
2 36155 1 11478
2 36156 1 11485
2 36157 1 11485
2 36158 1 11485
2 36159 1 11485
2 36160 1 11491
2 36161 1 11491
2 36162 1 11499
2 36163 1 11499
2 36164 1 11500
2 36165 1 11500
2 36166 1 11500
2 36167 1 11500
2 36168 1 11504
2 36169 1 11504
2 36170 1 11504
2 36171 1 11505
2 36172 1 11505
2 36173 1 11513
2 36174 1 11513
2 36175 1 11563
2 36176 1 11563
2 36177 1 11563
2 36178 1 11563
2 36179 1 11563
2 36180 1 11586
2 36181 1 11586
2 36182 1 11623
2 36183 1 11623
2 36184 1 11623
2 36185 1 11632
2 36186 1 11632
2 36187 1 11640
2 36188 1 11640
2 36189 1 11640
2 36190 1 11646
2 36191 1 11646
2 36192 1 11652
2 36193 1 11652
2 36194 1 11661
2 36195 1 11661
2 36196 1 11662
2 36197 1 11662
2 36198 1 11685
2 36199 1 11685
2 36200 1 11685
2 36201 1 11712
2 36202 1 11712
2 36203 1 11712
2 36204 1 11721
2 36205 1 11721
2 36206 1 11733
2 36207 1 11733
2 36208 1 11734
2 36209 1 11734
2 36210 1 11762
2 36211 1 11762
2 36212 1 11765
2 36213 1 11765
2 36214 1 11777
2 36215 1 11777
2 36216 1 11777
2 36217 1 11777
2 36218 1 11777
2 36219 1 11777
2 36220 1 11781
2 36221 1 11781
2 36222 1 11782
2 36223 1 11782
2 36224 1 11782
2 36225 1 11783
2 36226 1 11783
2 36227 1 11790
2 36228 1 11790
2 36229 1 11799
2 36230 1 11799
2 36231 1 11808
2 36232 1 11808
2 36233 1 11809
2 36234 1 11809
2 36235 1 11809
2 36236 1 11809
2 36237 1 11809
2 36238 1 11809
2 36239 1 11809
2 36240 1 11809
2 36241 1 11812
2 36242 1 11812
2 36243 1 11813
2 36244 1 11813
2 36245 1 11823
2 36246 1 11823
2 36247 1 11823
2 36248 1 11823
2 36249 1 11823
2 36250 1 11827
2 36251 1 11827
2 36252 1 11858
2 36253 1 11858
2 36254 1 11861
2 36255 1 11861
2 36256 1 11862
2 36257 1 11862
2 36258 1 11870
2 36259 1 11870
2 36260 1 11887
2 36261 1 11887
2 36262 1 11902
2 36263 1 11902
2 36264 1 11902
2 36265 1 11903
2 36266 1 11903
2 36267 1 11906
2 36268 1 11906
2 36269 1 11907
2 36270 1 11907
2 36271 1 11907
2 36272 1 11917
2 36273 1 11917
2 36274 1 11917
2 36275 1 11917
2 36276 1 11917
2 36277 1 11917
2 36278 1 11917
2 36279 1 11917
2 36280 1 11922
2 36281 1 11922
2 36282 1 11932
2 36283 1 11932
2 36284 1 11932
2 36285 1 11949
2 36286 1 11949
2 36287 1 11969
2 36288 1 11969
2 36289 1 11969
2 36290 1 12004
2 36291 1 12004
2 36292 1 12012
2 36293 1 12012
2 36294 1 12015
2 36295 1 12015
2 36296 1 12022
2 36297 1 12022
2 36298 1 12035
2 36299 1 12035
2 36300 1 12052
2 36301 1 12052
2 36302 1 12056
2 36303 1 12056
2 36304 1 12080
2 36305 1 12080
2 36306 1 12088
2 36307 1 12088
2 36308 1 12118
2 36309 1 12118
2 36310 1 12119
2 36311 1 12119
2 36312 1 12126
2 36313 1 12126
2 36314 1 12132
2 36315 1 12132
2 36316 1 12135
2 36317 1 12135
2 36318 1 12145
2 36319 1 12145
2 36320 1 12146
2 36321 1 12146
2 36322 1 12153
2 36323 1 12153
2 36324 1 12155
2 36325 1 12155
2 36326 1 12160
2 36327 1 12160
2 36328 1 12160
2 36329 1 12160
2 36330 1 12160
2 36331 1 12160
2 36332 1 12160
2 36333 1 12160
2 36334 1 12160
2 36335 1 12164
2 36336 1 12164
2 36337 1 12164
2 36338 1 12164
2 36339 1 12171
2 36340 1 12171
2 36341 1 12193
2 36342 1 12193
2 36343 1 12204
2 36344 1 12204
2 36345 1 12207
2 36346 1 12207
2 36347 1 12250
2 36348 1 12250
2 36349 1 12253
2 36350 1 12253
2 36351 1 12253
2 36352 1 12300
2 36353 1 12300
2 36354 1 12317
2 36355 1 12317
2 36356 1 12321
2 36357 1 12321
2 36358 1 12321
2 36359 1 12321
2 36360 1 12326
2 36361 1 12326
2 36362 1 12334
2 36363 1 12334
2 36364 1 12344
2 36365 1 12344
2 36366 1 12344
2 36367 1 12354
2 36368 1 12354
2 36369 1 12354
2 36370 1 12354
2 36371 1 12354
2 36372 1 12354
2 36373 1 12354
2 36374 1 12355
2 36375 1 12355
2 36376 1 12355
2 36377 1 12355
2 36378 1 12364
2 36379 1 12364
2 36380 1 12367
2 36381 1 12367
2 36382 1 12367
2 36383 1 12367
2 36384 1 12367
2 36385 1 12393
2 36386 1 12393
2 36387 1 12435
2 36388 1 12435
2 36389 1 12435
2 36390 1 12463
2 36391 1 12463
2 36392 1 12463
2 36393 1 12463
2 36394 1 12466
2 36395 1 12466
2 36396 1 12468
2 36397 1 12468
2 36398 1 12475
2 36399 1 12475
2 36400 1 12480
2 36401 1 12480
2 36402 1 12483
2 36403 1 12483
2 36404 1 12517
2 36405 1 12517
2 36406 1 12547
2 36407 1 12547
2 36408 1 12547
2 36409 1 12548
2 36410 1 12548
2 36411 1 12555
2 36412 1 12555
2 36413 1 12555
2 36414 1 12573
2 36415 1 12573
2 36416 1 12589
2 36417 1 12589
2 36418 1 12589
2 36419 1 12592
2 36420 1 12592
2 36421 1 12644
2 36422 1 12644
2 36423 1 12648
2 36424 1 12648
2 36425 1 12675
2 36426 1 12675
2 36427 1 12675
2 36428 1 12685
2 36429 1 12685
2 36430 1 12696
2 36431 1 12696
2 36432 1 12696
2 36433 1 12701
2 36434 1 12701
2 36435 1 12701
2 36436 1 12701
2 36437 1 12717
2 36438 1 12717
2 36439 1 12746
2 36440 1 12746
2 36441 1 12747
2 36442 1 12747
2 36443 1 12768
2 36444 1 12768
2 36445 1 12770
2 36446 1 12770
2 36447 1 12772
2 36448 1 12772
2 36449 1 12774
2 36450 1 12774
2 36451 1 12774
2 36452 1 12806
2 36453 1 12806
2 36454 1 12832
2 36455 1 12832
2 36456 1 12848
2 36457 1 12848
2 36458 1 12882
2 36459 1 12882
2 36460 1 12959
2 36461 1 12959
2 36462 1 12959
2 36463 1 12978
2 36464 1 12978
2 36465 1 12986
2 36466 1 12986
2 36467 1 13014
2 36468 1 13014
2 36469 1 13014
2 36470 1 13015
2 36471 1 13015
2 36472 1 13016
2 36473 1 13016
2 36474 1 13036
2 36475 1 13036
2 36476 1 13083
2 36477 1 13083
2 36478 1 13083
2 36479 1 13083
2 36480 1 13084
2 36481 1 13084
2 36482 1 13086
2 36483 1 13086
2 36484 1 13086
2 36485 1 13122
2 36486 1 13122
2 36487 1 13122
2 36488 1 13123
2 36489 1 13123
2 36490 1 13132
2 36491 1 13132
2 36492 1 13132
2 36493 1 13133
2 36494 1 13133
2 36495 1 13145
2 36496 1 13145
2 36497 1 13167
2 36498 1 13167
2 36499 1 13170
2 36500 1 13170
2 36501 1 13170
2 36502 1 13178
2 36503 1 13178
2 36504 1 13178
2 36505 1 13179
2 36506 1 13179
2 36507 1 13179
2 36508 1 13196
2 36509 1 13196
2 36510 1 13200
2 36511 1 13200
2 36512 1 13200
2 36513 1 13200
2 36514 1 13201
2 36515 1 13201
2 36516 1 13213
2 36517 1 13213
2 36518 1 13213
2 36519 1 13232
2 36520 1 13232
2 36521 1 13234
2 36522 1 13234
2 36523 1 13237
2 36524 1 13237
2 36525 1 13237
2 36526 1 13237
2 36527 1 13256
2 36528 1 13256
2 36529 1 13279
2 36530 1 13279
2 36531 1 13280
2 36532 1 13280
2 36533 1 13289
2 36534 1 13289
2 36535 1 13294
2 36536 1 13294
2 36537 1 13326
2 36538 1 13326
2 36539 1 13327
2 36540 1 13327
2 36541 1 13341
2 36542 1 13341
2 36543 1 13341
2 36544 1 13341
2 36545 1 13341
2 36546 1 13341
2 36547 1 13342
2 36548 1 13342
2 36549 1 13343
2 36550 1 13343
2 36551 1 13344
2 36552 1 13344
2 36553 1 13344
2 36554 1 13355
2 36555 1 13355
2 36556 1 13364
2 36557 1 13364
2 36558 1 13365
2 36559 1 13365
2 36560 1 13365
2 36561 1 13373
2 36562 1 13373
2 36563 1 13373
2 36564 1 13374
2 36565 1 13374
2 36566 1 13374
2 36567 1 13375
2 36568 1 13375
2 36569 1 13375
2 36570 1 13386
2 36571 1 13386
2 36572 1 13386
2 36573 1 13386
2 36574 1 13386
2 36575 1 13386
2 36576 1 13386
2 36577 1 13386
2 36578 1 13386
2 36579 1 13386
2 36580 1 13387
2 36581 1 13387
2 36582 1 13387
2 36583 1 13397
2 36584 1 13397
2 36585 1 13397
2 36586 1 13400
2 36587 1 13400
2 36588 1 13403
2 36589 1 13403
2 36590 1 13423
2 36591 1 13423
2 36592 1 13424
2 36593 1 13424
2 36594 1 13424
2 36595 1 13424
2 36596 1 13424
2 36597 1 13434
2 36598 1 13434
2 36599 1 13443
2 36600 1 13443
2 36601 1 13443
2 36602 1 13448
2 36603 1 13448
2 36604 1 13465
2 36605 1 13465
2 36606 1 13465
2 36607 1 13466
2 36608 1 13466
2 36609 1 13489
2 36610 1 13489
2 36611 1 13532
2 36612 1 13532
2 36613 1 13541
2 36614 1 13541
2 36615 1 13566
2 36616 1 13566
2 36617 1 13578
2 36618 1 13578
2 36619 1 13582
2 36620 1 13582
2 36621 1 13583
2 36622 1 13583
2 36623 1 13583
2 36624 1 13592
2 36625 1 13592
2 36626 1 13593
2 36627 1 13593
2 36628 1 13593
2 36629 1 13594
2 36630 1 13594
2 36631 1 13602
2 36632 1 13602
2 36633 1 13609
2 36634 1 13609
2 36635 1 13609
2 36636 1 13619
2 36637 1 13619
2 36638 1 13629
2 36639 1 13629
2 36640 1 13639
2 36641 1 13639
2 36642 1 13639
2 36643 1 13639
2 36644 1 13640
2 36645 1 13640
2 36646 1 13674
2 36647 1 13674
2 36648 1 13675
2 36649 1 13675
2 36650 1 13686
2 36651 1 13686
2 36652 1 13689
2 36653 1 13689
2 36654 1 13690
2 36655 1 13690
2 36656 1 13701
2 36657 1 13701
2 36658 1 13713
2 36659 1 13713
2 36660 1 13765
2 36661 1 13765
2 36662 1 13765
2 36663 1 13771
2 36664 1 13771
2 36665 1 13796
2 36666 1 13796
2 36667 1 13799
2 36668 1 13799
2 36669 1 13842
2 36670 1 13842
2 36671 1 13842
2 36672 1 13842
2 36673 1 13842
2 36674 1 13864
2 36675 1 13864
2 36676 1 13864
2 36677 1 13881
2 36678 1 13881
2 36679 1 13881
2 36680 1 13884
2 36681 1 13884
2 36682 1 13890
2 36683 1 13890
2 36684 1 13901
2 36685 1 13901
2 36686 1 13905
2 36687 1 13905
2 36688 1 13905
2 36689 1 13905
2 36690 1 13915
2 36691 1 13915
2 36692 1 13915
2 36693 1 13915
2 36694 1 13932
2 36695 1 13932
2 36696 1 13932
2 36697 1 13932
2 36698 1 13932
2 36699 1 13932
2 36700 1 13932
2 36701 1 13932
2 36702 1 13932
2 36703 1 13932
2 36704 1 13935
2 36705 1 13935
2 36706 1 13936
2 36707 1 13936
2 36708 1 13936
2 36709 1 13936
2 36710 1 13944
2 36711 1 13944
2 36712 1 13945
2 36713 1 13945
2 36714 1 13945
2 36715 1 13945
2 36716 1 13945
2 36717 1 13959
2 36718 1 13959
2 36719 1 13959
2 36720 1 13959
2 36721 1 13959
2 36722 1 13959
2 36723 1 13959
2 36724 1 13959
2 36725 1 13959
2 36726 1 13961
2 36727 1 13961
2 36728 1 13963
2 36729 1 13963
2 36730 1 13970
2 36731 1 13970
2 36732 1 13970
2 36733 1 13979
2 36734 1 13979
2 36735 1 13986
2 36736 1 13986
2 36737 1 13997
2 36738 1 13997
2 36739 1 13999
2 36740 1 13999
2 36741 1 14001
2 36742 1 14001
2 36743 1 14002
2 36744 1 14002
2 36745 1 14002
2 36746 1 14002
2 36747 1 14002
2 36748 1 14002
2 36749 1 14002
2 36750 1 14002
2 36751 1 14002
2 36752 1 14002
2 36753 1 14002
2 36754 1 14002
2 36755 1 14002
2 36756 1 14032
2 36757 1 14032
2 36758 1 14035
2 36759 1 14035
2 36760 1 14035
2 36761 1 14035
2 36762 1 14035
2 36763 1 14035
2 36764 1 14035
2 36765 1 14035
2 36766 1 14036
2 36767 1 14036
2 36768 1 14037
2 36769 1 14037
2 36770 1 14038
2 36771 1 14038
2 36772 1 14038
2 36773 1 14042
2 36774 1 14042
2 36775 1 14042
2 36776 1 14056
2 36777 1 14056
2 36778 1 14056
2 36779 1 14056
2 36780 1 14056
2 36781 1 14056
2 36782 1 14056
2 36783 1 14056
2 36784 1 14056
2 36785 1 14056
2 36786 1 14056
2 36787 1 14056
2 36788 1 14056
2 36789 1 14056
2 36790 1 14056
2 36791 1 14056
2 36792 1 14056
2 36793 1 14056
2 36794 1 14056
2 36795 1 14056
2 36796 1 14061
2 36797 1 14061
2 36798 1 14061
2 36799 1 14061
2 36800 1 14069
2 36801 1 14069
2 36802 1 14069
2 36803 1 14069
2 36804 1 14069
2 36805 1 14069
2 36806 1 14069
2 36807 1 14069
2 36808 1 14069
2 36809 1 14069
2 36810 1 14069
2 36811 1 14069
2 36812 1 14069
2 36813 1 14069
2 36814 1 14069
2 36815 1 14069
2 36816 1 14069
2 36817 1 14069
2 36818 1 14069
2 36819 1 14069
2 36820 1 14069
2 36821 1 14069
2 36822 1 14069
2 36823 1 14069
2 36824 1 14069
2 36825 1 14069
2 36826 1 14069
2 36827 1 14080
2 36828 1 14080
2 36829 1 14080
2 36830 1 14085
2 36831 1 14085
2 36832 1 14098
2 36833 1 14098
2 36834 1 14108
2 36835 1 14108
2 36836 1 14108
2 36837 1 14108
2 36838 1 14108
2 36839 1 14109
2 36840 1 14109
2 36841 1 14111
2 36842 1 14111
2 36843 1 14111
2 36844 1 14113
2 36845 1 14113
2 36846 1 14113
2 36847 1 14119
2 36848 1 14119
2 36849 1 14127
2 36850 1 14127
2 36851 1 14127
2 36852 1 14127
2 36853 1 14127
2 36854 1 14127
2 36855 1 14127
2 36856 1 14127
2 36857 1 14127
2 36858 1 14127
2 36859 1 14142
2 36860 1 14142
2 36861 1 14171
2 36862 1 14171
2 36863 1 14171
2 36864 1 14171
2 36865 1 14172
2 36866 1 14172
2 36867 1 14174
2 36868 1 14174
2 36869 1 14174
2 36870 1 14174
2 36871 1 14175
2 36872 1 14175
2 36873 1 14182
2 36874 1 14182
2 36875 1 14182
2 36876 1 14184
2 36877 1 14184
2 36878 1 14187
2 36879 1 14187
2 36880 1 14187
2 36881 1 14202
2 36882 1 14202
2 36883 1 14202
2 36884 1 14203
2 36885 1 14203
2 36886 1 14203
2 36887 1 14212
2 36888 1 14212
2 36889 1 14229
2 36890 1 14229
2 36891 1 14233
2 36892 1 14233
2 36893 1 14234
2 36894 1 14234
2 36895 1 14234
2 36896 1 14234
2 36897 1 14234
2 36898 1 14234
2 36899 1 14234
2 36900 1 14234
2 36901 1 14253
2 36902 1 14253
2 36903 1 14262
2 36904 1 14262
2 36905 1 14262
2 36906 1 14262
2 36907 1 14262
2 36908 1 14262
2 36909 1 14278
2 36910 1 14278
2 36911 1 14280
2 36912 1 14280
2 36913 1 14280
2 36914 1 14280
2 36915 1 14280
2 36916 1 14280
2 36917 1 14292
2 36918 1 14292
2 36919 1 14294
2 36920 1 14294
2 36921 1 14298
2 36922 1 14298
2 36923 1 14301
2 36924 1 14301
2 36925 1 14301
2 36926 1 14304
2 36927 1 14304
2 36928 1 14305
2 36929 1 14305
2 36930 1 14335
2 36931 1 14335
2 36932 1 14335
2 36933 1 14380
2 36934 1 14380
2 36935 1 14389
2 36936 1 14389
2 36937 1 14390
2 36938 1 14390
2 36939 1 14391
2 36940 1 14391
2 36941 1 14392
2 36942 1 14392
2 36943 1 14392
2 36944 1 14392
2 36945 1 14392
2 36946 1 14392
2 36947 1 14392
2 36948 1 14392
2 36949 1 14392
2 36950 1 14393
2 36951 1 14393
2 36952 1 14396
2 36953 1 14396
2 36954 1 14396
2 36955 1 14396
2 36956 1 14396
2 36957 1 14396
2 36958 1 14396
2 36959 1 14396
2 36960 1 14407
2 36961 1 14407
2 36962 1 14407
2 36963 1 14426
2 36964 1 14426
2 36965 1 14426
2 36966 1 14426
2 36967 1 14426
2 36968 1 14427
2 36969 1 14427
2 36970 1 14446
2 36971 1 14446
2 36972 1 14446
2 36973 1 14448
2 36974 1 14448
2 36975 1 14486
2 36976 1 14486
2 36977 1 14487
2 36978 1 14487
2 36979 1 14487
2 36980 1 14487
2 36981 1 14487
2 36982 1 14487
2 36983 1 14508
2 36984 1 14508
2 36985 1 14513
2 36986 1 14513
2 36987 1 14522
2 36988 1 14522
2 36989 1 14522
2 36990 1 14522
2 36991 1 14523
2 36992 1 14523
2 36993 1 14524
2 36994 1 14524
2 36995 1 14524
2 36996 1 14524
2 36997 1 14536
2 36998 1 14536
2 36999 1 14546
2 37000 1 14546
2 37001 1 14546
2 37002 1 14546
2 37003 1 14553
2 37004 1 14553
2 37005 1 14554
2 37006 1 14554
2 37007 1 14554
2 37008 1 14554
2 37009 1 14554
2 37010 1 14564
2 37011 1 14564
2 37012 1 14564
2 37013 1 14564
2 37014 1 14564
2 37015 1 14564
2 37016 1 14564
2 37017 1 14564
2 37018 1 14566
2 37019 1 14566
2 37020 1 14568
2 37021 1 14568
2 37022 1 14576
2 37023 1 14576
2 37024 1 14576
2 37025 1 14577
2 37026 1 14577
2 37027 1 14579
2 37028 1 14579
2 37029 1 14591
2 37030 1 14591
2 37031 1 14604
2 37032 1 14604
2 37033 1 14604
2 37034 1 14604
2 37035 1 14604
2 37036 1 14617
2 37037 1 14617
2 37038 1 14629
2 37039 1 14629
2 37040 1 14634
2 37041 1 14634
2 37042 1 14655
2 37043 1 14655
2 37044 1 14660
2 37045 1 14660
2 37046 1 14674
2 37047 1 14674
2 37048 1 14676
2 37049 1 14676
2 37050 1 14677
2 37051 1 14677
2 37052 1 14679
2 37053 1 14679
2 37054 1 14685
2 37055 1 14685
2 37056 1 14686
2 37057 1 14686
2 37058 1 14686
2 37059 1 14686
2 37060 1 14694
2 37061 1 14694
2 37062 1 14697
2 37063 1 14697
2 37064 1 14697
2 37065 1 14697
2 37066 1 14702
2 37067 1 14702
2 37068 1 14704
2 37069 1 14704
2 37070 1 14704
2 37071 1 14704
2 37072 1 14720
2 37073 1 14720
2 37074 1 14720
2 37075 1 14755
2 37076 1 14755
2 37077 1 14756
2 37078 1 14756
2 37079 1 14756
2 37080 1 14756
2 37081 1 14756
2 37082 1 14756
2 37083 1 14757
2 37084 1 14757
2 37085 1 14757
2 37086 1 14761
2 37087 1 14761
2 37088 1 14761
2 37089 1 14782
2 37090 1 14782
2 37091 1 14784
2 37092 1 14784
2 37093 1 14815
2 37094 1 14815
2 37095 1 14823
2 37096 1 14823
2 37097 1 14824
2 37098 1 14824
2 37099 1 14846
2 37100 1 14846
2 37101 1 14856
2 37102 1 14856
2 37103 1 14856
2 37104 1 14898
2 37105 1 14898
2 37106 1 14906
2 37107 1 14906
2 37108 1 14926
2 37109 1 14926
2 37110 1 14930
2 37111 1 14930
2 37112 1 14934
2 37113 1 14934
2 37114 1 14934
2 37115 1 14934
2 37116 1 14934
2 37117 1 14934
2 37118 1 14934
2 37119 1 14934
2 37120 1 14934
2 37121 1 14934
2 37122 1 14934
2 37123 1 14934
2 37124 1 14934
2 37125 1 14934
2 37126 1 14934
2 37127 1 14934
2 37128 1 14935
2 37129 1 14935
2 37130 1 14935
2 37131 1 14940
2 37132 1 14940
2 37133 1 14940
2 37134 1 14940
2 37135 1 14941
2 37136 1 14941
2 37137 1 14942
2 37138 1 14942
2 37139 1 14943
2 37140 1 14943
2 37141 1 14955
2 37142 1 14955
2 37143 1 14955
2 37144 1 14956
2 37145 1 14956
2 37146 1 14956
2 37147 1 14999
2 37148 1 14999
2 37149 1 15008
2 37150 1 15008
2 37151 1 15017
2 37152 1 15017
2 37153 1 15037
2 37154 1 15037
2 37155 1 15038
2 37156 1 15038
2 37157 1 15055
2 37158 1 15055
2 37159 1 15064
2 37160 1 15064
2 37161 1 15065
2 37162 1 15065
2 37163 1 15066
2 37164 1 15066
2 37165 1 15067
2 37166 1 15067
2 37167 1 15067
2 37168 1 15067
2 37169 1 15072
2 37170 1 15072
2 37171 1 15080
2 37172 1 15080
2 37173 1 15087
2 37174 1 15087
2 37175 1 15112
2 37176 1 15112
2 37177 1 15122
2 37178 1 15122
2 37179 1 15125
2 37180 1 15125
2 37181 1 15125
2 37182 1 15125
2 37183 1 15125
2 37184 1 15125
2 37185 1 15125
2 37186 1 15125
2 37187 1 15125
2 37188 1 15126
2 37189 1 15126
2 37190 1 15127
2 37191 1 15127
2 37192 1 15127
2 37193 1 15155
2 37194 1 15155
2 37195 1 15159
2 37196 1 15159
2 37197 1 15174
2 37198 1 15174
2 37199 1 15174
2 37200 1 15185
2 37201 1 15185
2 37202 1 15204
2 37203 1 15204
2 37204 1 15220
2 37205 1 15220
2 37206 1 15220
2 37207 1 15220
2 37208 1 15233
2 37209 1 15233
2 37210 1 15233
2 37211 1 15239
2 37212 1 15239
2 37213 1 15245
2 37214 1 15245
2 37215 1 15253
2 37216 1 15253
2 37217 1 15267
2 37218 1 15267
2 37219 1 15302
2 37220 1 15302
2 37221 1 15311
2 37222 1 15311
2 37223 1 15316
2 37224 1 15316
2 37225 1 15317
2 37226 1 15317
2 37227 1 15317
2 37228 1 15317
2 37229 1 15327
2 37230 1 15327
2 37231 1 15331
2 37232 1 15331
2 37233 1 15340
2 37234 1 15340
2 37235 1 15367
2 37236 1 15367
2 37237 1 15367
2 37238 1 15367
2 37239 1 15370
2 37240 1 15370
2 37241 1 15370
2 37242 1 15375
2 37243 1 15375
2 37244 1 15375
2 37245 1 15392
2 37246 1 15392
2 37247 1 15400
2 37248 1 15400
2 37249 1 15400
2 37250 1 15400
2 37251 1 15400
2 37252 1 15423
2 37253 1 15423
2 37254 1 15453
2 37255 1 15453
2 37256 1 15454
2 37257 1 15454
2 37258 1 15454
2 37259 1 15454
2 37260 1 15462
2 37261 1 15462
2 37262 1 15476
2 37263 1 15476
2 37264 1 15484
2 37265 1 15484
2 37266 1 15484
2 37267 1 15485
2 37268 1 15485
2 37269 1 15485
2 37270 1 15485
2 37271 1 15485
2 37272 1 15486
2 37273 1 15486
2 37274 1 15488
2 37275 1 15488
2 37276 1 15507
2 37277 1 15507
2 37278 1 15507
2 37279 1 15510
2 37280 1 15510
2 37281 1 15510
2 37282 1 15518
2 37283 1 15518
2 37284 1 15518
2 37285 1 15519
2 37286 1 15519
2 37287 1 15521
2 37288 1 15521
2 37289 1 15524
2 37290 1 15524
2 37291 1 15524
2 37292 1 15524
2 37293 1 15524
2 37294 1 15524
2 37295 1 15533
2 37296 1 15533
2 37297 1 15533
2 37298 1 15534
2 37299 1 15534
2 37300 1 15534
2 37301 1 15534
2 37302 1 15534
2 37303 1 15536
2 37304 1 15536
2 37305 1 15549
2 37306 1 15549
2 37307 1 15556
2 37308 1 15556
2 37309 1 15564
2 37310 1 15564
2 37311 1 15564
2 37312 1 15564
2 37313 1 15574
2 37314 1 15574
2 37315 1 15575
2 37316 1 15575
2 37317 1 15588
2 37318 1 15588
2 37319 1 15591
2 37320 1 15591
2 37321 1 15599
2 37322 1 15599
2 37323 1 15619
2 37324 1 15619
2 37325 1 15625
2 37326 1 15625
2 37327 1 15625
2 37328 1 15630
2 37329 1 15630
2 37330 1 15630
2 37331 1 15630
2 37332 1 15641
2 37333 1 15641
2 37334 1 15641
2 37335 1 15646
2 37336 1 15646
2 37337 1 15647
2 37338 1 15647
2 37339 1 15687
2 37340 1 15687
2 37341 1 15692
2 37342 1 15692
2 37343 1 15710
2 37344 1 15710
2 37345 1 15745
2 37346 1 15745
2 37347 1 15745
2 37348 1 15745
2 37349 1 15745
2 37350 1 15745
2 37351 1 15745
2 37352 1 15745
2 37353 1 15746
2 37354 1 15746
2 37355 1 15775
2 37356 1 15775
2 37357 1 15802
2 37358 1 15802
2 37359 1 15802
2 37360 1 15802
2 37361 1 15802
2 37362 1 15802
2 37363 1 15802
2 37364 1 15811
2 37365 1 15811
2 37366 1 15847
2 37367 1 15847
2 37368 1 15848
2 37369 1 15848
2 37370 1 15848
2 37371 1 15855
2 37372 1 15855
2 37373 1 15856
2 37374 1 15856
2 37375 1 15856
2 37376 1 15869
2 37377 1 15869
2 37378 1 15870
2 37379 1 15870
2 37380 1 15870
2 37381 1 15873
2 37382 1 15873
2 37383 1 15874
2 37384 1 15874
2 37385 1 15874
2 37386 1 15874
2 37387 1 15875
2 37388 1 15875
2 37389 1 15878
2 37390 1 15878
2 37391 1 15878
2 37392 1 15883
2 37393 1 15883
2 37394 1 15885
2 37395 1 15885
2 37396 1 15885
2 37397 1 15886
2 37398 1 15886
2 37399 1 15893
2 37400 1 15893
2 37401 1 15896
2 37402 1 15896
2 37403 1 15896
2 37404 1 15898
2 37405 1 15898
2 37406 1 15902
2 37407 1 15902
2 37408 1 15913
2 37409 1 15913
2 37410 1 15914
2 37411 1 15914
2 37412 1 15931
2 37413 1 15931
2 37414 1 15948
2 37415 1 15948
2 37416 1 15948
2 37417 1 15948
2 37418 1 15960
2 37419 1 15960
2 37420 1 15967
2 37421 1 15967
2 37422 1 15970
2 37423 1 15970
2 37424 1 15990
2 37425 1 15990
2 37426 1 16027
2 37427 1 16027
2 37428 1 16034
2 37429 1 16034
2 37430 1 16057
2 37431 1 16057
2 37432 1 16081
2 37433 1 16081
2 37434 1 16109
2 37435 1 16109
2 37436 1 16119
2 37437 1 16119
2 37438 1 16129
2 37439 1 16129
2 37440 1 16129
2 37441 1 16129
2 37442 1 16129
2 37443 1 16130
2 37444 1 16130
2 37445 1 16140
2 37446 1 16140
2 37447 1 16140
2 37448 1 16154
2 37449 1 16154
2 37450 1 16154
2 37451 1 16155
2 37452 1 16155
2 37453 1 16164
2 37454 1 16164
2 37455 1 16164
2 37456 1 16164
2 37457 1 16164
2 37458 1 16177
2 37459 1 16177
2 37460 1 16177
2 37461 1 16178
2 37462 1 16178
2 37463 1 16178
2 37464 1 16179
2 37465 1 16179
2 37466 1 16180
2 37467 1 16180
2 37468 1 16180
2 37469 1 16184
2 37470 1 16184
2 37471 1 16187
2 37472 1 16187
2 37473 1 16192
2 37474 1 16192
2 37475 1 16208
2 37476 1 16208
2 37477 1 16250
2 37478 1 16250
2 37479 1 16283
2 37480 1 16283
2 37481 1 16283
2 37482 1 16283
2 37483 1 16309
2 37484 1 16309
2 37485 1 16379
2 37486 1 16379
2 37487 1 16412
2 37488 1 16412
2 37489 1 16419
2 37490 1 16419
2 37491 1 16451
2 37492 1 16451
2 37493 1 16503
2 37494 1 16503
2 37495 1 16506
2 37496 1 16506
2 37497 1 16522
2 37498 1 16522
2 37499 1 16541
2 37500 1 16541
2 37501 1 16565
2 37502 1 16565
2 37503 1 16565
2 37504 1 16566
2 37505 1 16566
2 37506 1 16566
2 37507 1 16574
2 37508 1 16574
2 37509 1 16584
2 37510 1 16584
2 37511 1 16584
2 37512 1 16584
2 37513 1 16588
2 37514 1 16588
2 37515 1 16605
2 37516 1 16605
2 37517 1 16614
2 37518 1 16614
2 37519 1 16616
2 37520 1 16616
2 37521 1 16625
2 37522 1 16625
2 37523 1 16629
2 37524 1 16629
2 37525 1 16629
2 37526 1 16629
2 37527 1 16638
2 37528 1 16638
2 37529 1 16638
2 37530 1 16638
2 37531 1 16653
2 37532 1 16653
2 37533 1 16663
2 37534 1 16663
2 37535 1 16677
2 37536 1 16677
2 37537 1 16703
2 37538 1 16703
2 37539 1 16718
2 37540 1 16718
2 37541 1 16718
2 37542 1 16718
2 37543 1 16787
2 37544 1 16787
2 37545 1 16787
2 37546 1 16787
2 37547 1 16787
2 37548 1 16788
2 37549 1 16788
2 37550 1 16790
2 37551 1 16790
2 37552 1 16817
2 37553 1 16817
2 37554 1 16834
2 37555 1 16834
2 37556 1 16835
2 37557 1 16835
2 37558 1 16837
2 37559 1 16837
2 37560 1 16838
2 37561 1 16838
2 37562 1 16839
2 37563 1 16839
2 37564 1 16840
2 37565 1 16840
2 37566 1 16844
2 37567 1 16844
2 37568 1 16857
2 37569 1 16857
2 37570 1 16857
2 37571 1 16857
2 37572 1 16857
2 37573 1 16857
2 37574 1 16873
2 37575 1 16873
2 37576 1 16882
2 37577 1 16882
2 37578 1 16896
2 37579 1 16896
2 37580 1 16896
2 37581 1 16896
2 37582 1 16896
2 37583 1 16900
2 37584 1 16900
2 37585 1 16900
2 37586 1 16909
2 37587 1 16909
2 37588 1 16909
2 37589 1 16909
2 37590 1 16909
2 37591 1 16910
2 37592 1 16910
2 37593 1 16925
2 37594 1 16925
2 37595 1 16954
2 37596 1 16954
2 37597 1 16957
2 37598 1 16957
2 37599 1 16982
2 37600 1 16982
2 37601 1 17013
2 37602 1 17013
2 37603 1 17019
2 37604 1 17019
2 37605 1 17019
2 37606 1 17025
2 37607 1 17025
2 37608 1 17053
2 37609 1 17053
2 37610 1 17053
2 37611 1 17053
2 37612 1 17054
2 37613 1 17054
2 37614 1 17054
2 37615 1 17054
2 37616 1 17058
2 37617 1 17058
2 37618 1 17067
2 37619 1 17067
2 37620 1 17087
2 37621 1 17087
2 37622 1 17120
2 37623 1 17120
2 37624 1 17120
2 37625 1 17132
2 37626 1 17132
2 37627 1 17150
2 37628 1 17150
2 37629 1 17150
2 37630 1 17158
2 37631 1 17158
2 37632 1 17163
2 37633 1 17163
2 37634 1 17163
2 37635 1 17163
2 37636 1 17163
2 37637 1 17163
2 37638 1 17163
2 37639 1 17178
2 37640 1 17178
2 37641 1 17220
2 37642 1 17220
2 37643 1 17222
2 37644 1 17222
2 37645 1 17226
2 37646 1 17226
2 37647 1 17226
2 37648 1 17226
2 37649 1 17228
2 37650 1 17228
2 37651 1 17239
2 37652 1 17239
2 37653 1 17323
2 37654 1 17323
2 37655 1 17323
2 37656 1 17324
2 37657 1 17324
2 37658 1 17330
2 37659 1 17330
2 37660 1 17340
2 37661 1 17340
2 37662 1 17354
2 37663 1 17354
2 37664 1 17354
2 37665 1 17357
2 37666 1 17357
2 37667 1 17361
2 37668 1 17361
2 37669 1 17362
2 37670 1 17362
2 37671 1 17362
2 37672 1 17362
2 37673 1 17362
2 37674 1 17362
2 37675 1 17362
2 37676 1 17362
2 37677 1 17365
2 37678 1 17365
2 37679 1 17366
2 37680 1 17366
2 37681 1 17367
2 37682 1 17367
2 37683 1 17367
2 37684 1 17370
2 37685 1 17370
2 37686 1 17371
2 37687 1 17371
2 37688 1 17371
2 37689 1 17373
2 37690 1 17373
2 37691 1 17375
2 37692 1 17375
2 37693 1 17382
2 37694 1 17382
2 37695 1 17401
2 37696 1 17401
2 37697 1 17404
2 37698 1 17404
2 37699 1 17404
2 37700 1 17424
2 37701 1 17424
2 37702 1 17424
2 37703 1 17424
2 37704 1 17425
2 37705 1 17425
2 37706 1 17425
2 37707 1 17425
2 37708 1 17428
2 37709 1 17428
2 37710 1 17428
2 37711 1 17428
2 37712 1 17428
2 37713 1 17428
2 37714 1 17428
2 37715 1 17428
2 37716 1 17428
2 37717 1 17428
2 37718 1 17428
2 37719 1 17437
2 37720 1 17437
2 37721 1 17437
2 37722 1 17445
2 37723 1 17445
2 37724 1 17445
2 37725 1 17464
2 37726 1 17464
2 37727 1 17464
2 37728 1 17472
2 37729 1 17472
2 37730 1 17472
2 37731 1 17476
2 37732 1 17476
2 37733 1 17476
2 37734 1 17490
2 37735 1 17490
2 37736 1 17495
2 37737 1 17495
2 37738 1 17495
2 37739 1 17495
2 37740 1 17514
2 37741 1 17514
2 37742 1 17514
2 37743 1 17514
2 37744 1 17515
2 37745 1 17515
2 37746 1 17517
2 37747 1 17517
2 37748 1 17518
2 37749 1 17518
2 37750 1 17518
2 37751 1 17536
2 37752 1 17536
2 37753 1 17536
2 37754 1 17542
2 37755 1 17542
2 37756 1 17551
2 37757 1 17551
2 37758 1 17562
2 37759 1 17562
2 37760 1 17562
2 37761 1 17562
2 37762 1 17562
2 37763 1 17575
2 37764 1 17575
2 37765 1 17575
2 37766 1 17575
2 37767 1 17604
2 37768 1 17604
2 37769 1 17610
2 37770 1 17610
2 37771 1 17614
2 37772 1 17614
2 37773 1 17625
2 37774 1 17625
2 37775 1 17634
2 37776 1 17634
2 37777 1 17640
2 37778 1 17640
2 37779 1 17640
2 37780 1 17640
2 37781 1 17649
2 37782 1 17649
2 37783 1 17649
2 37784 1 17660
2 37785 1 17660
2 37786 1 17660
2 37787 1 17667
2 37788 1 17667
2 37789 1 17668
2 37790 1 17668
2 37791 1 17693
2 37792 1 17693
2 37793 1 17693
2 37794 1 17711
2 37795 1 17711
2 37796 1 17720
2 37797 1 17720
2 37798 1 17720
2 37799 1 17721
2 37800 1 17721
2 37801 1 17732
2 37802 1 17732
2 37803 1 17737
2 37804 1 17737
2 37805 1 17740
2 37806 1 17740
2 37807 1 17745
2 37808 1 17745
2 37809 1 17745
2 37810 1 17755
2 37811 1 17755
2 37812 1 17799
2 37813 1 17799
2 37814 1 17799
2 37815 1 17805
2 37816 1 17805
2 37817 1 17819
2 37818 1 17819
2 37819 1 17835
2 37820 1 17835
2 37821 1 17836
2 37822 1 17836
2 37823 1 17854
2 37824 1 17854
2 37825 1 17863
2 37826 1 17863
2 37827 1 17864
2 37828 1 17864
2 37829 1 17899
2 37830 1 17899
2 37831 1 17909
2 37832 1 17909
2 37833 1 17909
2 37834 1 17910
2 37835 1 17910
2 37836 1 17943
2 37837 1 17943
2 37838 1 17943
2 37839 1 17943
2 37840 1 17965
2 37841 1 17965
2 37842 1 17973
2 37843 1 17973
2 37844 1 17975
2 37845 1 17975
2 37846 1 17978
2 37847 1 17978
2 37848 1 17981
2 37849 1 17981
2 37850 1 17981
2 37851 1 17982
2 37852 1 17982
2 37853 1 17982
2 37854 1 17998
2 37855 1 17998
2 37856 1 18012
2 37857 1 18012
2 37858 1 18028
2 37859 1 18028
2 37860 1 18041
2 37861 1 18041
2 37862 1 18041
2 37863 1 18054
2 37864 1 18054
2 37865 1 18078
2 37866 1 18078
2 37867 1 18080
2 37868 1 18080
2 37869 1 18083
2 37870 1 18083
2 37871 1 18094
2 37872 1 18094
2 37873 1 18097
2 37874 1 18097
2 37875 1 18100
2 37876 1 18100
2 37877 1 18100
2 37878 1 18103
2 37879 1 18103
2 37880 1 18143
2 37881 1 18143
2 37882 1 18155
2 37883 1 18155
2 37884 1 18163
2 37885 1 18163
2 37886 1 18164
2 37887 1 18164
2 37888 1 18237
2 37889 1 18237
2 37890 1 18250
2 37891 1 18250
2 37892 1 18289
2 37893 1 18289
2 37894 1 18289
2 37895 1 18291
2 37896 1 18291
2 37897 1 18292
2 37898 1 18292
2 37899 1 18292
2 37900 1 18299
2 37901 1 18299
2 37902 1 18299
2 37903 1 18303
2 37904 1 18303
2 37905 1 18303
2 37906 1 18306
2 37907 1 18306
2 37908 1 18306
2 37909 1 18313
2 37910 1 18313
2 37911 1 18324
2 37912 1 18324
2 37913 1 18326
2 37914 1 18326
2 37915 1 18351
2 37916 1 18351
2 37917 1 18354
2 37918 1 18354
2 37919 1 18369
2 37920 1 18369
2 37921 1 18403
2 37922 1 18403
2 37923 1 18419
2 37924 1 18419
2 37925 1 18419
2 37926 1 18429
2 37927 1 18429
2 37928 1 18479
2 37929 1 18479
2 37930 1 18536
2 37931 1 18536
2 37932 1 18544
2 37933 1 18544
2 37934 1 18559
2 37935 1 18559
2 37936 1 18559
2 37937 1 18559
2 37938 1 18559
2 37939 1 18586
2 37940 1 18586
2 37941 1 18589
2 37942 1 18589
2 37943 1 18617
2 37944 1 18617
2 37945 1 18637
2 37946 1 18637
2 37947 1 18637
2 37948 1 18637
2 37949 1 18637
2 37950 1 18638
2 37951 1 18638
2 37952 1 18639
2 37953 1 18639
2 37954 1 18649
2 37955 1 18649
2 37956 1 18652
2 37957 1 18652
2 37958 1 18711
2 37959 1 18711
2 37960 1 18721
2 37961 1 18721
2 37962 1 18731
2 37963 1 18731
2 37964 1 18782
2 37965 1 18782
2 37966 1 18799
2 37967 1 18799
2 37968 1 18801
2 37969 1 18801
2 37970 1 18833
2 37971 1 18833
2 37972 1 18833
2 37973 1 18843
2 37974 1 18843
2 37975 1 18847
2 37976 1 18847
2 37977 1 18862
2 37978 1 18862
2 37979 1 18870
2 37980 1 18870
2 37981 1 18871
2 37982 1 18871
2 37983 1 18879
2 37984 1 18879
2 37985 1 18889
2 37986 1 18889
2 37987 1 18907
2 37988 1 18907
2 37989 1 18926
2 37990 1 18926
2 37991 1 18926
2 37992 1 18926
2 37993 1 18926
2 37994 1 18926
2 37995 1 18926
2 37996 1 18939
2 37997 1 18939
2 37998 1 18980
2 37999 1 18980
2 38000 1 18995
2 38001 1 18995
2 38002 1 19030
2 38003 1 19030
2 38004 1 19042
2 38005 1 19042
2 38006 1 19042
2 38007 1 19042
2 38008 1 19043
2 38009 1 19043
2 38010 1 19050
2 38011 1 19050
2 38012 1 19052
2 38013 1 19052
2 38014 1 19052
2 38015 1 19055
2 38016 1 19055
2 38017 1 19055
2 38018 1 19061
2 38019 1 19061
2 38020 1 19061
2 38021 1 19067
2 38022 1 19067
2 38023 1 19067
2 38024 1 19067
2 38025 1 19071
2 38026 1 19071
2 38027 1 19074
2 38028 1 19074
2 38029 1 19082
2 38030 1 19082
2 38031 1 19111
2 38032 1 19111
2 38033 1 19111
2 38034 1 19143
2 38035 1 19143
2 38036 1 19159
2 38037 1 19159
2 38038 1 19159
2 38039 1 19183
2 38040 1 19183
2 38041 1 19183
2 38042 1 19195
2 38043 1 19195
2 38044 1 19195
2 38045 1 19231
2 38046 1 19231
2 38047 1 19251
2 38048 1 19251
2 38049 1 19251
2 38050 1 19251
2 38051 1 19298
2 38052 1 19298
2 38053 1 19304
2 38054 1 19304
2 38055 1 19331
2 38056 1 19331
2 38057 1 19341
2 38058 1 19341
2 38059 1 19342
2 38060 1 19342
2 38061 1 19352
2 38062 1 19352
2 38063 1 19357
2 38064 1 19357
2 38065 1 19358
2 38066 1 19358
2 38067 1 19360
2 38068 1 19360
2 38069 1 19361
2 38070 1 19361
2 38071 1 19392
2 38072 1 19392
2 38073 1 19393
2 38074 1 19393
2 38075 1 19404
2 38076 1 19404
2 38077 1 19412
2 38078 1 19412
2 38079 1 19414
2 38080 1 19414
2 38081 1 19434
2 38082 1 19434
2 38083 1 19499
2 38084 1 19499
2 38085 1 19500
2 38086 1 19500
2 38087 1 19505
2 38088 1 19505
2 38089 1 19505
2 38090 1 19505
2 38091 1 19517
2 38092 1 19517
2 38093 1 19518
2 38094 1 19518
2 38095 1 19539
2 38096 1 19539
2 38097 1 19583
2 38098 1 19583
2 38099 1 19595
2 38100 1 19595
2 38101 1 19600
2 38102 1 19600
2 38103 1 19600
2 38104 1 19646
2 38105 1 19646
2 38106 1 19681
2 38107 1 19681
2 38108 1 19708
2 38109 1 19708
2 38110 1 19726
2 38111 1 19726
2 38112 1 19726
2 38113 1 19732
2 38114 1 19732
2 38115 1 19732
2 38116 1 19758
2 38117 1 19758
2 38118 1 19765
2 38119 1 19765
2 38120 1 19768
2 38121 1 19768
2 38122 1 19802
2 38123 1 19802
2 38124 1 19815
2 38125 1 19815
2 38126 1 19815
2 38127 1 19823
2 38128 1 19823
2 38129 1 19824
2 38130 1 19824
2 38131 1 19869
2 38132 1 19869
2 38133 1 19869
2 38134 1 19869
2 38135 1 19869
2 38136 1 19911
2 38137 1 19911
2 38138 1 19925
2 38139 1 19925
2 38140 1 19949
2 38141 1 19949
2 38142 1 20010
2 38143 1 20010
2 38144 1 20023
2 38145 1 20023
2 38146 1 20024
2 38147 1 20024
2 38148 1 20032
2 38149 1 20032
2 38150 1 20104
2 38151 1 20104
2 38152 1 20134
2 38153 1 20134
2 38154 1 20151
2 38155 1 20151
2 38156 1 20162
2 38157 1 20162
2 38158 1 20172
2 38159 1 20172
2 38160 1 20172
2 38161 1 20172
2 38162 1 20178
2 38163 1 20178
2 38164 1 20179
2 38165 1 20179
2 38166 1 20194
2 38167 1 20194
2 38168 1 20206
2 38169 1 20206
2 38170 1 20228
2 38171 1 20228
2 38172 1 20228
2 38173 1 20257
2 38174 1 20257
2 38175 1 20264
2 38176 1 20264
2 38177 1 20265
2 38178 1 20265
2 38179 1 20274
2 38180 1 20274
2 38181 1 20274
2 38182 1 20275
2 38183 1 20275
2 38184 1 20278
2 38185 1 20278
2 38186 1 20278
2 38187 1 20279
2 38188 1 20279
2 38189 1 20290
2 38190 1 20290
2 38191 1 20312
2 38192 1 20312
2 38193 1 20326
2 38194 1 20326
2 38195 1 20326
2 38196 1 20326
2 38197 1 20332
2 38198 1 20332
2 38199 1 20332
2 38200 1 20346
2 38201 1 20346
2 38202 1 20346
2 38203 1 20358
2 38204 1 20358
2 38205 1 20359
2 38206 1 20359
2 38207 1 20365
2 38208 1 20365
2 38209 1 20365
2 38210 1 20365
2 38211 1 20370
2 38212 1 20370
2 38213 1 20370
2 38214 1 20370
2 38215 1 20377
2 38216 1 20377
2 38217 1 20378
2 38218 1 20378
2 38219 1 20419
2 38220 1 20419
2 38221 1 20419
2 38222 1 20443
2 38223 1 20443
2 38224 1 20443
2 38225 1 20474
2 38226 1 20474
2 38227 1 20506
2 38228 1 20506
2 38229 1 20506
2 38230 1 20517
2 38231 1 20517
2 38232 1 20520
2 38233 1 20520
2 38234 1 20550
2 38235 1 20550
2 38236 1 20604
2 38237 1 20604
2 38238 1 20644
2 38239 1 20644
2 38240 1 20659
2 38241 1 20659
2 38242 1 20680
2 38243 1 20680
2 38244 1 20692
2 38245 1 20692
2 38246 1 20768
2 38247 1 20768
2 38248 1 20768
2 38249 1 20774
2 38250 1 20774
2 38251 1 20785
2 38252 1 20785
2 38253 1 20793
2 38254 1 20793
2 38255 1 20900
2 38256 1 20900
2 38257 1 20908
2 38258 1 20908
2 38259 1 20926
2 38260 1 20926
2 38261 1 20926
2 38262 1 20926
2 38263 1 20938
2 38264 1 20938
2 38265 1 20941
2 38266 1 20941
2 38267 1 20942
2 38268 1 20942
2 38269 1 20960
2 38270 1 20960
2 38271 1 20974
2 38272 1 20974
2 38273 1 20996
2 38274 1 20996
2 38275 1 21008
2 38276 1 21008
2 38277 1 21117
2 38278 1 21117
2 38279 1 21117
2 38280 1 21117
2 38281 1 21175
2 38282 1 21175
2 38283 1 21196
2 38284 1 21196
2 38285 1 21232
2 38286 1 21232
2 38287 1 21284
2 38288 1 21284
2 38289 1 21284
2 38290 1 21321
2 38291 1 21321
2 38292 1 21325
2 38293 1 21325
2 38294 1 21347
2 38295 1 21347
2 38296 1 21361
2 38297 1 21361
2 38298 1 21366
2 38299 1 21366
2 38300 1 21366
2 38301 1 21366
2 38302 1 21393
2 38303 1 21393
2 38304 1 21425
2 38305 1 21425
2 38306 1 21429
2 38307 1 21429
2 38308 1 21429
2 38309 1 21431
2 38310 1 21431
2 38311 1 21432
2 38312 1 21432
2 38313 1 21498
2 38314 1 21498
2 38315 1 21522
2 38316 1 21522
2 38317 1 21522
2 38318 1 21586
2 38319 1 21586
2 38320 1 21589
2 38321 1 21589
2 38322 1 21590
2 38323 1 21590
2 38324 1 21594
2 38325 1 21594
2 38326 1 21612
2 38327 1 21612
2 38328 1 21641
2 38329 1 21641
2 38330 1 21642
2 38331 1 21642
2 38332 1 21644
2 38333 1 21644
2 38334 1 21706
2 38335 1 21706
2 38336 1 21718
2 38337 1 21718
2 38338 1 21763
2 38339 1 21763
2 38340 1 21843
2 38341 1 21843
2 38342 1 21944
2 38343 1 21944
2 38344 1 21944
2 38345 1 22071
2 38346 1 22071
2 38347 1 22146
2 38348 1 22146
2 38349 1 22196
2 38350 1 22196
2 38351 1 22204
2 38352 1 22204
2 38353 1 22260
2 38354 1 22260
2 38355 1 22274
2 38356 1 22274
0 27 5 51 1 25
0 28 5 133 1 22373
0 29 5 102 1 22527
0 30 5 94 1 22663
0 31 5 85 1 22776
0 32 5 126 1 22872
0 33 5 76 1 22990
0 34 5 100 1 23056
0 35 5 56 1 23157
0 36 5 85 1 23207
0 37 5 79 1 23289
0 38 5 69 1 23368
0 39 5 55 1 23438
0 40 5 67 1 23490
0 41 5 71 1 23567
0 42 5 58 1 23596
0 43 5 1 1 23645
0 44 5 74 1 23647
0 45 5 113 1 23750
0 46 5 98 1 23860
0 47 5 89 1 23962
0 48 5 90 1 24048
0 49 5 95 1 24140
0 50 5 77 1 24221
0 51 5 42 1 24309
0 52 7 35 2 22777 23439
0 53 5 1 1 26325
0 54 7 21 2 23369 23963
0 55 5 4 1 26360
0 56 7 4 2 24805 23491
0 57 5 2 1 26385
0 58 7 7 2 22991 25451
0 59 7 21 2 23597 26283
0 60 5 23 1 26398
0 61 7 1 2 26391 26399
0 62 5 2 1 61
0 63 7 1 2 26389 26442
0 64 5 1 1 63
0 65 7 1 2 23057 64
0 66 5 1 1 65
0 67 7 21 2 24806 25452
0 68 5 13 1 26444
0 69 7 3 2 23058 25453
0 70 5 3 1 26478
0 71 7 17 2 25589 24310
0 72 5 24 1 26484
0 73 7 7 2 22992 25007
0 74 7 1 2 26485 26525
0 75 5 2 1 74
0 76 7 1 2 26481 26532
0 77 5 1 1 76
0 78 7 1 2 26465 77
0 79 5 1 1 78
0 80 7 1 2 66 79
0 81 5 1 1 80
0 82 7 1 2 26206 81
0 83 5 1 1 82
0 84 7 9 2 22873 25454
0 85 5 2 1 26534
0 86 7 4 2 23059 26284
0 87 5 3 1 26545
0 88 7 1 2 26535 26546
0 89 5 1 1 88
0 90 7 2 2 23492 24222
0 91 5 1 1 26552
0 92 7 1 2 26526 26553
0 93 5 1 1 92
0 94 7 1 2 89 93
0 95 5 1 1 94
0 96 7 1 2 23598 95
0 97 5 1 1 96
0 98 7 4 2 24931 23493
0 99 5 2 1 26554
0 100 7 8 2 22874 24223
0 101 5 1 1 26560
0 102 7 1 2 26558 101
0 103 5 1 1 102
0 104 7 12 2 24932 24224
0 105 5 27 1 26568
0 106 7 5 2 25008 23599
0 107 5 2 1 26607
0 108 7 8 2 23060 25590
0 109 5 1 1 26614
0 110 7 1 2 26612 109
0 111 5 12 1 110
0 112 7 1 2 26580 26622
0 113 7 1 2 103 112
0 114 5 1 1 113
0 115 7 1 2 97 114
0 116 7 1 2 83 115
0 117 5 1 1 116
0 118 7 1 2 26111 117
0 119 5 1 1 118
0 120 7 7 2 24225 26419
0 121 5 9 1 26634
0 122 7 4 2 23061 26641
0 123 5 1 1 26650
0 124 7 1 2 24141 26651
0 125 5 2 1 124
0 126 7 8 2 24226 26285
0 127 5 2 1 26656
0 128 7 8 2 26207 24311
0 129 7 2 2 25591 26666
0 130 5 4 1 26674
0 131 7 1 2 26664 26676
0 132 5 2 1 131
0 133 7 9 2 25592 24227
0 134 5 1 1 26682
0 135 7 1 2 23062 134
0 136 5 2 1 135
0 137 7 1 2 22993 26691
0 138 7 1 2 26680 137
0 139 5 1 1 138
0 140 7 1 2 26654 139
0 141 5 1 1 140
0 142 7 1 2 23494 141
0 143 5 1 1 142
0 144 7 4 2 24142 26286
0 145 7 8 2 23063 23600
0 146 5 5 1 26697
0 147 7 5 2 26208 26698
0 148 5 1 1 26710
0 149 7 4 2 26693 26711
0 150 7 1 2 22994 26715
0 151 5 1 1 150
0 152 7 1 2 143 151
0 153 5 1 1 152
0 154 7 1 2 22875 153
0 155 5 1 1 154
0 156 7 3 2 23064 26400
0 157 5 2 1 26719
0 158 7 3 2 23495 24143
0 159 5 2 1 26724
0 160 7 19 2 22995 26209
0 161 5 14 1 26729
0 162 7 1 2 26725 26730
0 163 7 1 2 26720 162
0 164 5 1 1 163
0 165 7 1 2 155 164
0 166 7 1 2 119 165
0 167 5 1 1 166
0 168 7 1 2 26361 167
0 169 5 1 1 168
0 170 7 17 2 25327 25932
0 171 5 1 1 26762
0 172 7 5 2 25455 26112
0 173 5 2 1 26779
0 174 7 2 2 26727 26784
0 175 5 20 1 26786
0 176 7 1 2 26748 26420
0 177 5 3 1 176
0 178 7 14 2 26581 26808
0 179 7 5 2 26788 26811
0 180 7 5 2 22876 26825
0 181 7 1 2 26763 26830
0 182 5 1 1 181
0 183 7 1 2 169 182
0 184 5 1 1 183
0 185 7 1 2 26326 184
0 186 5 1 1 185
0 187 7 8 2 23370 25396
0 188 7 14 2 24720 25933
0 189 7 2 2 26835 26843
0 190 5 1 1 26857
0 191 7 1 2 26831 26858
0 192 5 1 1 191
0 193 7 1 2 186 192
0 194 5 1 1 193
0 195 7 1 2 23861 194
0 196 5 1 1 195
0 197 7 8 2 22877 25328
0 198 5 1 1 26859
0 199 7 5 2 24721 25834
0 200 7 5 2 23964 26867
0 201 7 2 2 25397 26872
0 202 5 1 1 26877
0 203 7 1 2 26860 26878
0 204 7 1 2 26826 203
0 205 5 1 1 204
0 206 7 1 2 196 205
0 207 5 1 1 206
0 208 7 1 2 22664 207
0 209 5 1 1 208
0 210 7 19 2 24722 25398
0 211 5 1 1 26879
0 212 7 2 2 26381 171
0 213 5 25 1 26898
0 214 7 5 2 25835 26900
0 215 7 2 2 26880 26925
0 216 5 1 1 26930
0 217 7 24 2 25836 23965
0 218 7 5 2 25329 26932
0 219 5 1 1 26956
0 220 7 18 2 23862 25934
0 221 7 5 2 23371 26961
0 222 5 1 1 26979
0 223 7 1 2 219 222
0 224 5 23 1 223
0 225 7 1 2 26327 26984
0 226 5 1 1 225
0 227 7 1 2 216 226
0 228 5 2 1 227
0 229 7 3 2 24626 27007
0 230 5 1 1 27009
0 231 7 1 2 27010 26832
0 232 5 1 1 231
0 233 7 1 2 209 232
0 234 5 1 1 233
0 235 7 1 2 23290 234
0 236 5 1 1 235
0 237 7 16 2 25248 25837
0 238 5 1 1 27012
0 239 7 12 2 23372 25935
0 240 5 1 1 27028
0 241 7 15 2 25330 23966
0 242 5 2 1 27040
0 243 7 38 2 240 27055
0 244 7 1 2 26328 27057
0 245 5 1 1 244
0 246 7 1 2 190 245
0 247 5 1 1 246
0 248 7 1 2 22665 247
0 249 5 1 1 248
0 250 7 2 2 24627 27029
0 251 5 1 1 27095
0 252 7 1 2 26329 27096
0 253 5 1 1 252
0 254 7 1 2 249 253
0 255 5 2 1 254
0 256 7 3 2 27013 27097
0 257 7 1 2 26833 27099
0 258 5 1 1 257
0 259 7 1 2 236 258
0 260 5 1 1 259
0 261 7 1 2 23751 260
0 262 5 1 1 261
0 263 7 7 2 25249 25721
0 264 7 3 2 23863 27102
0 265 7 1 2 53 26899
0 266 5 1 1 265
0 267 7 1 2 211 27056
0 268 5 1 1 267
0 269 7 1 2 24628 268
0 270 7 1 2 266 269
0 271 5 1 1 270
0 272 7 2 2 22666 26881
0 273 5 1 1 27112
0 274 7 2 2 27113 27041
0 275 5 1 1 27114
0 276 7 1 2 271 275
0 277 5 1 1 276
0 278 7 3 2 27109 277
0 279 7 1 2 26834 27116
0 280 5 1 1 279
0 281 7 1 2 262 280
0 282 5 1 1 281
0 283 7 1 2 22528 282
0 284 5 1 1 283
0 285 7 1 2 24629 26330
0 286 5 1 1 285
0 287 7 1 2 273 286
0 288 5 21 1 287
0 289 7 9 2 23752 25936
0 290 7 10 2 23373 25838
0 291 7 3 2 27140 27149
0 292 5 2 1 27159
0 293 7 8 2 25722 23967
0 294 7 11 2 25331 23864
0 295 7 2 2 27164 27172
0 296 5 1 1 27183
0 297 7 1 2 27162 296
0 298 5 4 1 297
0 299 7 1 2 23291 27185
0 300 5 2 1 299
0 301 7 1 2 27103 26985
0 302 5 1 1 301
0 303 7 1 2 27189 302
0 304 5 1 1 303
0 305 7 1 2 27119 304
0 306 5 2 1 305
0 307 7 32 2 25723 23865
0 308 7 4 2 25250 27193
0 309 5 1 1 27225
0 310 7 21 2 23753 25839
0 311 5 1 1 27229
0 312 7 1 2 23292 27230
0 313 5 2 1 312
0 314 7 1 2 309 27250
0 315 5 12 1 314
0 316 7 8 2 22667 22778
0 317 7 8 2 23440 27264
0 318 7 1 2 27252 27272
0 319 5 2 1 318
0 320 7 8 2 23293 23866
0 321 5 4 1 27282
0 322 7 2 2 238 27290
0 323 5 35 1 27294
0 324 7 16 2 24630 24723
0 325 7 9 2 25399 27331
0 326 7 3 2 27296 27347
0 327 5 1 1 27356
0 328 7 1 2 25724 27357
0 329 5 1 1 328
0 330 7 1 2 27280 329
0 331 5 1 1 330
0 332 7 1 2 27058 331
0 333 5 1 1 332
0 334 7 1 2 27191 333
0 335 5 1 1 334
0 336 7 8 2 24524 22878
0 337 7 1 2 27359 26827
0 338 7 1 2 335 337
0 339 5 1 1 338
0 340 7 1 2 284 339
0 341 5 1 1 340
0 342 7 1 2 23208 341
0 343 5 1 1 342
0 344 7 6 2 22879 25163
0 345 7 1 2 23294 26986
0 346 5 1 1 345
0 347 7 4 2 25251 27030
0 348 5 1 1 27373
0 349 7 1 2 25840 27374
0 350 5 1 1 349
0 351 7 1 2 346 350
0 352 5 2 1 351
0 353 7 1 2 22529 27377
0 354 5 1 1 353
0 355 7 13 2 23295 23374
0 356 5 1 1 27379
0 357 7 10 2 24525 25937
0 358 7 2 2 27380 27392
0 359 5 1 1 27402
0 360 7 1 2 25841 27403
0 361 5 1 1 360
0 362 7 1 2 354 361
0 363 5 1 1 362
0 364 7 1 2 27120 363
0 365 5 1 1 364
0 366 7 1 2 27297 27273
0 367 5 1 1 366
0 368 7 12 2 24631 25842
0 369 7 8 2 24724 23296
0 370 7 2 2 25400 27416
0 371 7 1 2 27404 27424
0 372 5 1 1 371
0 373 7 1 2 367 372
0 374 5 2 1 373
0 375 7 1 2 22530 27426
0 376 5 1 1 375
0 377 7 15 2 23297 25843
0 378 5 2 1 27428
0 379 7 16 2 24526 22668
0 380 7 2 2 27445 26331
0 381 5 1 1 27461
0 382 7 1 2 27429 27462
0 383 5 1 1 382
0 384 7 1 2 376 383
0 385 5 1 1 384
0 386 7 1 2 27059 385
0 387 5 1 1 386
0 388 7 1 2 365 387
0 389 5 1 1 388
0 390 7 1 2 25725 26828
0 391 7 2 2 389 390
0 392 7 1 2 27367 27463
0 393 5 1 1 392
0 394 7 1 2 343 393
0 395 5 1 1 394
0 396 7 1 2 22374 395
0 397 5 1 1 396
0 398 7 6 2 22880 23209
0 399 7 2 2 24391 27465
0 400 7 1 2 27471 27464
0 401 5 1 1 400
0 402 7 1 2 397 401
0 403 5 1 1 402
0 404 7 1 2 24049 403
0 405 5 1 1 404
0 406 7 11 2 26501 26421
0 407 7 13 2 22996 24228
0 408 5 5 1 27484
0 409 7 10 2 24050 26113
0 410 7 4 2 22881 27502
0 411 5 1 1 27512
0 412 7 11 2 26021 24144
0 413 5 1 1 27516
0 414 7 3 2 24807 27517
0 415 5 1 1 27527
0 416 7 1 2 411 415
0 417 5 12 1 416
0 418 7 1 2 27485 27530
0 419 5 1 1 418
0 420 7 12 2 24933 26210
0 421 5 1 1 27542
0 422 7 2 2 23496 27503
0 423 5 2 1 27554
0 424 7 2 2 25456 27518
0 425 5 1 1 27558
0 426 7 1 2 23065 27559
0 427 5 1 1 426
0 428 7 1 2 27556 427
0 429 5 1 1 428
0 430 7 1 2 27543 429
0 431 5 1 1 430
0 432 7 1 2 419 431
0 433 5 1 1 432
0 434 7 1 2 26362 433
0 435 5 1 1 434
0 436 7 3 2 23066 25332
0 437 7 2 2 22882 27560
0 438 7 3 2 27497 421
0 439 5 26 1 27565
0 440 7 3 2 25938 27568
0 441 7 20 2 25457 24145
0 442 5 8 1 27597
0 443 7 3 2 24051 27617
0 444 7 2 2 27594 27625
0 445 7 1 2 27563 27628
0 446 5 1 1 445
0 447 7 1 2 435 446
0 448 5 1 1 447
0 449 7 1 2 26332 448
0 450 5 1 1 449
0 451 7 3 2 24725 26836
0 452 5 1 1 27630
0 453 7 7 2 22883 23067
0 454 7 1 2 27631 27633
0 455 7 1 2 27629 454
0 456 5 1 1 455
0 457 7 1 2 450 456
0 458 5 1 1 457
0 459 7 1 2 23867 458
0 460 5 1 1 459
0 461 7 2 2 27569 27626
0 462 7 10 2 24726 23068
0 463 5 1 1 27642
0 464 7 5 2 22884 25401
0 465 7 1 2 27643 27652
0 466 7 1 2 26957 465
0 467 7 1 2 27640 466
0 468 5 1 1 467
0 469 7 1 2 460 468
0 470 5 1 1 469
0 471 7 1 2 22669 470
0 472 5 1 1 471
0 473 7 8 2 24632 22885
0 474 7 2 2 27570 27657
0 475 7 8 2 23069 24052
0 476 5 1 1 27667
0 477 7 2 2 27618 27668
0 478 7 1 2 27665 27675
0 479 7 1 2 27008 478
0 480 5 1 1 479
0 481 7 1 2 472 480
0 482 5 1 1 481
0 483 7 1 2 23298 482
0 484 5 1 1 483
0 485 7 4 2 22886 27619
0 486 5 1 1 27677
0 487 7 2 2 23070 27571
0 488 7 2 2 27678 27681
0 489 7 2 2 24053 27683
0 490 7 1 2 27100 27685
0 491 5 1 1 490
0 492 7 1 2 484 491
0 493 5 1 1 492
0 494 7 1 2 23754 493
0 495 5 1 1 494
0 496 7 1 2 27117 27686
0 497 5 1 1 496
0 498 7 1 2 495 497
0 499 5 1 1 498
0 500 7 1 2 22531 499
0 501 5 1 1 500
0 502 7 3 2 25402 27194
0 503 7 3 2 24633 27417
0 504 7 1 2 27687 27690
0 505 5 1 1 504
0 506 7 1 2 27281 505
0 507 5 1 1 506
0 508 7 2 2 26901 507
0 509 5 1 1 27693
0 510 7 10 2 24634 23968
0 511 5 3 1 27695
0 512 7 2 2 26868 27696
0 513 7 1 2 26837 27104
0 514 7 1 2 27708 513
0 515 5 1 1 514
0 516 7 1 2 27192 515
0 517 7 1 2 509 516
0 518 5 2 1 517
0 519 7 2 2 27572 27360
0 520 7 1 2 27712 27676
0 521 7 1 2 27710 520
0 522 5 1 1 521
0 523 7 1 2 501 522
0 524 5 1 1 523
0 525 7 1 2 23210 524
0 526 5 1 1 525
0 527 7 14 2 23071 25164
0 528 7 2 2 22887 27714
0 529 7 8 2 27121 26987
0 530 5 1 1 27730
0 531 7 3 2 27150 27697
0 532 5 1 1 27738
0 533 7 1 2 26882 27739
0 534 5 1 1 533
0 535 7 6 2 23441 23868
0 536 7 3 2 27265 27741
0 537 7 1 2 27060 27747
0 538 5 1 1 537
0 539 7 1 2 534 538
0 540 7 1 2 530 539
0 541 5 1 1 540
0 542 7 1 2 23299 541
0 543 5 1 1 542
0 544 7 10 2 25252 23375
0 545 5 1 1 27750
0 546 7 2 2 25844 27751
0 547 7 1 2 23969 27274
0 548 7 1 2 27760 547
0 549 5 1 1 548
0 550 7 1 2 543 549
0 551 5 1 1 550
0 552 7 1 2 22532 551
0 553 5 1 1 552
0 554 7 6 2 23442 27381
0 555 7 6 2 24527 27266
0 556 7 2 2 26933 27768
0 557 7 1 2 27762 27774
0 558 5 1 1 557
0 559 7 1 2 553 558
0 560 5 1 1 559
0 561 7 3 2 25726 27573
0 562 7 1 2 27776 27627
0 563 7 2 2 560 562
0 564 7 1 2 27728 27779
0 565 5 1 1 564
0 566 7 1 2 526 565
0 567 5 1 1 566
0 568 7 1 2 22375 567
0 569 5 1 1 568
0 570 7 9 2 23072 23211
0 571 7 3 2 24392 22888
0 572 7 1 2 27781 27790
0 573 7 1 2 27780 572
0 574 5 1 1 573
0 575 7 1 2 569 574
0 576 5 1 1 575
0 577 7 1 2 27473 576
0 578 5 1 1 577
0 579 7 23 2 24934 25009
0 580 5 4 1 27793
0 581 7 1 2 22533 27348
0 582 5 1 1 581
0 583 7 1 2 381 582
0 584 5 3 1 583
0 585 7 1 2 27253 27820
0 586 5 2 1 585
0 587 7 8 2 24528 27332
0 588 7 3 2 23300 25403
0 589 7 1 2 27195 27833
0 590 7 1 2 27825 589
0 591 5 1 1 590
0 592 7 2 2 27823 591
0 593 7 17 2 22534 22670
0 594 5 1 1 27838
0 595 7 3 2 27839 26333
0 596 7 2 2 23755 27298
0 597 7 1 2 27855 27858
0 598 5 1 1 597
0 599 7 1 2 27836 598
0 600 5 1 1 599
0 601 7 1 2 23212 600
0 602 5 1 1 601
0 603 7 7 2 23301 25727
0 604 7 12 2 22535 25165
0 605 5 1 1 27867
0 606 7 1 2 27860 27868
0 607 7 1 2 27748 606
0 608 5 2 1 607
0 609 7 1 2 602 27879
0 610 5 1 1 609
0 611 7 1 2 22376 610
0 612 5 1 1 611
0 613 7 6 2 22671 23302
0 614 7 2 2 27881 26334
0 615 7 3 2 24393 27887
0 616 5 1 1 27889
0 617 7 8 2 22536 23213
0 618 5 1 1 27892
0 619 7 2 2 27890 27893
0 620 5 1 1 27900
0 621 7 1 2 27196 27901
0 622 5 2 1 621
0 623 7 1 2 612 27902
0 624 5 1 1 623
0 625 7 1 2 27061 624
0 626 5 1 1 625
0 627 7 11 2 24394 23214
0 628 5 1 1 27904
0 629 7 12 2 22377 25166
0 630 5 1 1 27915
0 631 7 7 2 628 630
0 632 5 63 1 27927
0 633 7 4 2 22779 23303
0 634 5 2 1 27997
0 635 7 3 2 24727 23443
0 636 5 2 1 28003
0 637 7 1 2 28001 28006
0 638 7 5 2 22672 25404
0 639 5 1 1 28008
0 640 7 8 2 24635 25253
0 641 5 1 1 28013
0 642 7 1 2 639 641
0 643 7 7 2 637 642
0 644 7 1 2 22537 28021
0 645 5 1 1 644
0 646 7 7 2 23304 23444
0 647 7 4 2 22780 28028
0 648 7 2 2 27446 28035
0 649 5 1 1 28039
0 650 7 1 2 645 649
0 651 5 9 1 650
0 652 7 1 2 27934 28041
0 653 5 1 1 652
0 654 7 12 2 22378 24529
0 655 7 6 2 24636 28050
0 656 7 11 2 23215 25254
0 657 7 3 2 28068 26883
0 658 7 1 2 28062 28079
0 659 5 1 1 658
0 660 7 1 2 653 659
0 661 5 1 1 660
0 662 7 1 2 27165 661
0 663 5 1 1 662
0 664 7 7 2 24530 23305
0 665 5 2 1 28082
0 666 7 8 2 22538 25255
0 667 5 1 1 28091
0 668 7 2 2 28089 667
0 669 5 77 1 28099
0 670 7 11 2 28101 27122
0 671 5 1 1 28178
0 672 7 28 2 22379 23216
0 673 5 7 1 28189
0 674 7 1 2 27141 28190
0 675 7 1 2 28179 674
0 676 5 1 1 675
0 677 7 1 2 663 676
0 678 5 1 1 677
0 679 7 1 2 27151 678
0 680 5 1 1 679
0 681 7 26 2 22539 23306
0 682 5 3 1 28224
0 683 7 12 2 23217 23756
0 684 5 3 1 28253
0 685 7 12 2 25167 25728
0 686 5 1 1 28268
0 687 7 2 2 28265 686
0 688 5 10 1 28280
0 689 7 1 2 28225 28282
0 690 5 1 1 689
0 691 7 27 2 24531 25256
0 692 5 5 1 28292
0 693 7 6 2 25729 28293
0 694 5 1 1 28324
0 695 7 2 2 23218 28325
0 696 5 1 1 28330
0 697 7 1 2 690 696
0 698 5 2 1 697
0 699 7 1 2 22380 28332
0 700 5 1 1 699
0 701 7 19 2 24395 22540
0 702 7 13 2 23219 23307
0 703 5 1 1 28353
0 704 7 4 2 28334 28354
0 705 7 2 2 25730 28366
0 706 5 1 1 28370
0 707 7 1 2 700 706
0 708 5 5 1 707
0 709 7 1 2 26988 28372
0 710 5 1 1 709
0 711 7 3 2 28102 28191
0 712 7 1 2 27184 28377
0 713 5 1 1 712
0 714 7 1 2 710 713
0 715 5 1 1 714
0 716 7 1 2 27123 715
0 717 5 1 1 716
0 718 7 1 2 680 717
0 719 7 1 2 626 718
0 720 5 1 1 719
0 721 7 16 2 24312 26683
0 722 7 1 2 26789 28380
0 723 7 1 2 720 722
0 724 5 1 1 723
0 725 7 6 2 23220 23376
0 726 7 4 2 28029 28396
0 727 7 4 2 22781 24146
0 728 5 2 1 28406
0 729 7 1 2 28402 28407
0 730 7 2 2 25458 23601
0 731 7 15 2 26211 26287
0 732 7 2 2 28412 28414
0 733 5 2 1 28429
0 734 7 18 2 23757 23869
0 735 5 2 1 28433
0 736 7 4 2 23970 28434
0 737 7 6 2 22381 27840
0 738 7 1 2 28453 28457
0 739 7 1 2 28430 738
0 740 7 1 2 729 739
0 741 5 1 1 740
0 742 7 1 2 724 741
0 743 5 1 1 742
0 744 7 1 2 27794 743
0 745 5 1 1 744
0 746 7 7 2 23073 24147
0 747 5 1 1 28463
0 748 7 4 2 25010 26212
0 749 5 1 1 28470
0 750 7 3 2 26486 28471
0 751 5 2 1 28474
0 752 7 1 2 747 28477
0 753 5 1 1 752
0 754 7 1 2 22997 753
0 755 5 1 1 754
0 756 7 2 2 27544 26401
0 757 5 3 1 28479
0 758 7 1 2 25011 28480
0 759 5 1 1 758
0 760 7 1 2 755 759
0 761 5 1 1 760
0 762 7 1 2 25459 761
0 763 5 1 1 762
0 764 7 5 2 25012 24148
0 765 5 1 1 28484
0 766 7 2 2 23497 26487
0 767 5 2 1 28489
0 768 7 1 2 28481 28491
0 769 5 1 1 768
0 770 7 1 2 28485 769
0 771 5 1 1 770
0 772 7 1 2 763 771
0 773 5 1 1 772
0 774 7 1 2 26363 773
0 775 5 1 1 774
0 776 7 22 2 23498 26114
0 777 5 10 1 28493
0 778 7 2 2 24935 26422
0 779 5 4 1 28525
0 780 7 2 2 22998 26502
0 781 5 2 1 28531
0 782 7 3 2 28527 28533
0 783 7 2 2 28515 28535
0 784 7 3 2 28472 28538
0 785 5 1 1 28540
0 786 7 1 2 26764 28541
0 787 5 1 1 786
0 788 7 15 2 22999 23074
0 789 5 1 1 28543
0 790 7 10 2 23971 24149
0 791 5 1 1 28558
0 792 7 3 2 23377 28559
0 793 5 1 1 28568
0 794 7 1 2 28544 28569
0 795 5 1 1 794
0 796 7 7 2 26115 24313
0 797 5 2 1 28571
0 798 7 2 2 27795 28572
0 799 5 1 1 28580
0 800 7 1 2 27062 28581
0 801 5 1 1 800
0 802 7 1 2 795 801
0 803 5 1 1 802
0 804 7 1 2 25593 803
0 805 5 1 1 804
0 806 7 11 2 24936 23075
0 807 5 1 1 28582
0 808 7 1 2 26364 28583
0 809 5 1 1 808
0 810 7 2 2 25013 26765
0 811 5 1 1 28593
0 812 7 1 2 23000 28594
0 813 5 1 1 812
0 814 7 1 2 809 813
0 815 5 1 1 814
0 816 7 2 2 28516 26402
0 817 7 1 2 815 28595
0 818 5 1 1 817
0 819 7 4 2 26790 26423
0 820 5 1 1 28597
0 821 7 6 2 23378 23499
0 822 5 1 1 28601
0 823 7 1 2 27063 822
0 824 7 1 2 28598 823
0 825 5 1 1 824
0 826 7 1 2 818 825
0 827 7 1 2 805 826
0 828 5 1 1 827
0 829 7 1 2 24229 828
0 830 5 1 1 829
0 831 7 1 2 787 830
0 832 7 1 2 775 831
0 833 5 1 1 832
0 834 7 1 2 27749 833
0 835 5 1 1 834
0 836 7 3 2 24937 25594
0 837 7 2 2 28607 28573
0 838 5 1 1 28610
0 839 7 2 2 23001 23602
0 840 7 2 2 26288 28517
0 841 7 1 2 28612 28614
0 842 5 1 1 841
0 843 7 1 2 838 842
0 844 5 4 1 843
0 845 7 1 2 25014 28616
0 846 5 2 1 845
0 847 7 1 2 820 28620
0 848 5 3 1 847
0 849 7 1 2 24230 28622
0 850 5 1 1 849
0 851 7 1 2 785 850
0 852 5 3 1 851
0 853 7 2 2 22673 26989
0 854 5 3 1 28628
0 855 7 1 2 26884 28629
0 856 5 1 1 855
0 857 7 1 2 230 856
0 858 5 1 1 857
0 859 7 1 2 28625 858
0 860 5 1 1 859
0 861 7 1 2 835 860
0 862 5 1 1 861
0 863 7 1 2 23308 862
0 864 5 1 1 863
0 865 7 1 2 27101 28626
0 866 5 1 1 865
0 867 7 1 2 864 866
0 868 5 1 1 867
0 869 7 1 2 23758 868
0 870 5 1 1 869
0 871 7 1 2 27118 28627
0 872 5 1 1 871
0 873 7 1 2 22541 872
0 874 7 1 2 870 873
0 875 5 1 1 874
0 876 7 2 2 27197 27375
0 877 5 1 1 28633
0 878 7 1 2 27190 877
0 879 5 1 1 878
0 880 7 1 2 28623 879
0 881 5 1 1 880
0 882 7 22 2 28518 27620
0 883 7 5 2 23500 25595
0 884 5 2 1 28657
0 885 7 1 2 26289 28662
0 886 5 1 1 885
0 887 7 1 2 28635 886
0 888 5 1 1 887
0 889 7 1 2 28621 888
0 890 5 1 1 889
0 891 7 20 2 25257 25333
0 892 7 2 2 25731 26934
0 893 7 1 2 28664 28684
0 894 7 1 2 890 893
0 895 5 1 1 894
0 896 7 1 2 881 895
0 897 5 1 1 896
0 898 7 1 2 27124 897
0 899 5 1 1 898
0 900 7 1 2 26365 28617
0 901 5 1 1 900
0 902 7 3 2 25939 28599
0 903 7 1 2 25334 28686
0 904 5 1 1 903
0 905 7 1 2 901 904
0 906 5 1 1 905
0 907 7 1 2 25015 906
0 908 5 1 1 907
0 909 7 1 2 28658 28570
0 910 5 1 1 909
0 911 7 5 2 25596 25940
0 912 7 1 2 25335 28689
0 913 5 1 1 912
0 914 7 1 2 26382 913
0 915 5 2 1 914
0 916 7 1 2 24314 26791
0 917 7 1 2 28694 916
0 918 5 1 1 917
0 919 7 1 2 910 918
0 920 7 1 2 908 919
0 921 5 1 1 920
0 922 7 13 2 25732 25845
0 923 5 1 1 28696
0 924 7 2 2 25405 28697
0 925 7 1 2 25258 27333
0 926 7 1 2 28709 925
0 927 7 1 2 921 926
0 928 5 1 1 927
0 929 7 1 2 27694 28624
0 930 5 1 1 929
0 931 7 1 2 928 930
0 932 7 1 2 899 931
0 933 5 1 1 932
0 934 7 1 2 24231 933
0 935 5 1 1 934
0 936 7 1 2 27711 28542
0 937 5 1 1 936
0 938 7 1 2 24532 937
0 939 7 1 2 935 938
0 940 5 1 1 939
0 941 7 1 2 28192 940
0 942 7 1 2 875 941
0 943 5 1 1 942
0 944 7 7 2 25336 23445
0 945 5 1 1 28711
0 946 7 1 2 22782 28712
0 947 5 1 1 946
0 948 7 1 2 452 947
0 949 5 26 1 948
0 950 7 5 2 23309 23972
0 951 7 3 2 24637 28744
0 952 5 1 1 28749
0 953 7 1 2 28618 28750
0 954 5 1 1 953
0 955 7 11 2 22674 25259
0 956 7 1 2 28752 28687
0 957 5 1 1 956
0 958 7 1 2 954 957
0 959 5 1 1 958
0 960 7 1 2 22542 959
0 961 5 1 1 960
0 962 7 13 2 22675 25941
0 963 5 3 1 28763
0 964 7 3 2 28083 28764
0 965 5 1 1 28779
0 966 7 1 2 28780 28600
0 967 5 1 1 966
0 968 7 1 2 961 967
0 969 5 1 1 968
0 970 7 1 2 28718 969
0 971 5 1 1 970
0 972 7 12 2 25337 25406
0 973 7 5 2 23310 28782
0 974 5 1 1 28794
0 975 7 12 2 23379 23446
0 976 7 7 2 22783 28799
0 977 5 1 1 28811
0 978 7 1 2 974 977
0 979 5 1 1 978
0 980 7 12 2 28002 979
0 981 7 1 2 22543 28818
0 982 5 1 1 981
0 983 7 5 2 24533 22784
0 984 7 3 2 23311 28830
0 985 7 1 2 28800 28835
0 986 5 1 1 985
0 987 7 1 2 982 986
0 988 5 6 1 987
0 989 7 21 2 22676 23973
0 990 5 2 1 28844
0 991 7 1 2 28845 28619
0 992 5 1 1 991
0 993 7 1 2 24638 28688
0 994 5 1 1 993
0 995 7 1 2 992 994
0 996 5 1 1 995
0 997 7 1 2 28838 996
0 998 5 1 1 997
0 999 7 1 2 971 998
0 1000 5 1 1 999
0 1001 7 1 2 24232 1000
0 1002 5 1 1 1001
0 1003 7 1 2 22677 28819
0 1004 5 1 1 1003
0 1005 7 13 2 24639 23312
0 1006 7 1 2 28719 28867
0 1007 5 1 1 1006
0 1008 7 1 2 1004 1007
0 1009 5 2 1 1008
0 1010 7 1 2 22544 28880
0 1011 5 1 1 1010
0 1012 7 5 2 23313 28801
0 1013 7 1 2 28882 27769
0 1014 5 1 1 1013
0 1015 7 1 2 1011 1014
0 1016 5 2 1 1015
0 1017 7 4 2 23974 26213
0 1018 7 1 2 28889 28539
0 1019 7 1 2 28887 1018
0 1020 5 1 1 1019
0 1021 7 1 2 1002 1020
0 1022 5 1 1 1021
0 1023 7 1 2 25846 1022
0 1024 5 1 1 1023
0 1025 7 5 2 23603 26657
0 1026 5 2 1 28893
0 1027 7 1 2 28898 26677
0 1028 5 2 1 1027
0 1029 7 1 2 23002 28900
0 1030 5 1 1 1029
0 1031 7 1 2 28482 1030
0 1032 5 2 1 1031
0 1033 7 1 2 28519 28902
0 1034 5 1 1 1033
0 1035 7 2 2 24938 26116
0 1036 5 1 1 28904
0 1037 7 1 2 28905 28381
0 1038 5 2 1 1037
0 1039 7 1 2 1034 28906
0 1040 5 1 1 1039
0 1041 7 4 2 23870 28226
0 1042 5 1 1 28908
0 1043 7 2 2 27098 28909
0 1044 7 1 2 1040 28912
0 1045 5 1 1 1044
0 1046 7 1 2 1024 1045
0 1047 5 1 1 1046
0 1048 7 1 2 25016 1047
0 1049 5 1 1 1048
0 1050 7 1 2 26424 28913
0 1051 5 1 1 1050
0 1052 7 1 2 28042 28695
0 1053 5 1 1 1052
0 1054 7 2 2 23314 27042
0 1055 5 2 1 28914
0 1056 7 1 2 25597 27376
0 1057 5 1 1 1056
0 1058 7 1 2 28916 1057
0 1059 5 1 1 1058
0 1060 7 1 2 22545 1059
0 1061 5 1 1 1060
0 1062 7 4 2 24534 25598
0 1063 7 3 2 23315 27031
0 1064 7 1 2 28918 28922
0 1065 5 1 1 1064
0 1066 7 1 2 1061 1065
0 1067 5 1 1 1066
0 1068 7 1 2 27125 1067
0 1069 5 1 1 1068
0 1070 7 1 2 1053 1069
0 1071 5 1 1 1070
0 1072 7 3 2 25847 24315
0 1073 7 1 2 1071 28925
0 1074 5 1 1 1073
0 1075 7 1 2 1051 1074
0 1076 5 1 1 1075
0 1077 7 1 2 26792 1076
0 1078 5 1 1 1077
0 1079 7 3 2 25848 28560
0 1080 7 1 2 28928 28659
0 1081 7 1 2 28888 1080
0 1082 5 1 1 1081
0 1083 7 1 2 1078 1082
0 1084 5 1 1 1083
0 1085 7 1 2 24233 1084
0 1086 5 1 1 1085
0 1087 7 1 2 1049 1086
0 1088 5 1 1 1087
0 1089 7 1 2 25733 28217
0 1090 7 1 2 1088 1089
0 1091 5 1 1 1090
0 1092 7 1 2 943 1091
0 1093 5 1 1 1092
0 1094 7 24 2 24396 25168
0 1095 5 8 1 28931
0 1096 7 1 2 24808 28955
0 1097 7 1 2 1093 1096
0 1098 5 1 1 1097
0 1099 7 1 2 745 1098
0 1100 5 1 1 1099
0 1101 7 1 2 26022 1100
0 1102 5 1 1 1101
0 1103 7 1 2 578 1102
0 1104 7 1 2 405 1103
0 1105 5 1 1 1104
0 1106 7 1 2 23648 1105
0 1107 5 1 1 1106
0 1108 7 7 2 22785 25407
0 1109 5 1 1 28963
0 1110 7 1 2 28007 1109
0 1111 5 52 1 1110
0 1112 7 5 2 22678 24054
0 1113 7 3 2 25017 28536
0 1114 5 1 1 29027
0 1115 7 10 2 24939 25460
0 1116 5 1 1 29030
0 1117 7 7 2 23076 27474
0 1118 5 1 1 29040
0 1119 7 1 2 29031 29041
0 1120 5 1 1 1119
0 1121 7 1 2 1114 1120
0 1122 5 1 1 1121
0 1123 7 18 2 22889 23501
0 1124 5 8 1 29047
0 1125 7 1 2 26214 29065
0 1126 7 1 2 1122 1125
0 1127 5 1 1 1126
0 1128 7 5 2 25018 26403
0 1129 5 1 1 29073
0 1130 7 1 2 1129 1118
0 1131 5 7 1 1130
0 1132 7 1 2 25461 29078
0 1133 5 1 1 1132
0 1134 7 3 2 24809 26404
0 1135 5 1 1 29085
0 1136 7 1 2 25019 29086
0 1137 5 1 1 1136
0 1138 7 1 2 1133 1137
0 1139 5 1 1 1138
0 1140 7 1 2 23003 1139
0 1141 5 1 1 1140
0 1142 7 4 2 26390 26543
0 1143 5 31 1 29088
0 1144 7 2 2 29092 26425
0 1145 5 1 1 29123
0 1146 7 5 2 25020 26488
0 1147 5 1 1 29125
0 1148 7 1 2 26555 29126
0 1149 5 1 1 1148
0 1150 7 1 2 1145 1149
0 1151 7 1 2 1141 1150
0 1152 5 1 1 1151
0 1153 7 1 2 24234 1152
0 1154 5 1 1 1153
0 1155 7 1 2 1127 1154
0 1156 5 1 1 1155
0 1157 7 1 2 24150 1156
0 1158 5 1 1 1157
0 1159 7 1 2 26445 28903
0 1160 5 1 1 1159
0 1161 7 1 2 28907 1160
0 1162 5 1 1 1161
0 1163 7 1 2 25021 29066
0 1164 7 1 2 1162 1163
0 1165 5 1 1 1164
0 1166 7 1 2 1158 1165
0 1167 5 1 1 1166
0 1168 7 1 2 28373 1167
0 1169 5 1 1 1168
0 1170 7 3 2 24535 27935
0 1171 5 1 1 29130
0 1172 7 1 2 22382 28294
0 1173 5 2 1 1172
0 1174 7 5 2 23316 27936
0 1175 5 1 1 29135
0 1176 7 1 2 29133 1175
0 1177 5 1 1 1176
0 1178 7 36 2 1171 1177
0 1179 7 18 2 26117 24235
0 1180 5 1 1 29176
0 1181 7 2 2 29140 29177
0 1182 7 5 2 25462 25599
0 1183 5 1 1 29196
0 1184 7 1 2 24810 25734
0 1185 7 1 2 29197 1184
0 1186 7 1 2 29194 1185
0 1187 5 1 1 1186
0 1188 7 1 2 1169 1187
0 1189 5 1 1 1188
0 1190 7 1 2 23649 1189
0 1191 5 1 1 1190
0 1192 7 5 2 24536 28069
0 1193 5 1 1 29201
0 1194 7 8 2 25169 23317
0 1195 7 3 2 22546 29206
0 1196 5 1 1 29214
0 1197 7 1 2 1193 1196
0 1198 5 17 1 1197
0 1199 7 3 2 24397 29217
0 1200 5 1 1 29234
0 1201 7 7 2 27916 28295
0 1202 5 1 1 29237
0 1203 7 1 2 1200 1202
0 1204 5 25 1 1203
0 1205 7 18 2 24151 24236
0 1206 5 4 1 29269
0 1207 7 2 2 25647 29270
0 1208 7 2 2 23759 29291
0 1209 7 1 2 23077 26503
0 1210 5 3 1 1209
0 1211 7 1 2 29295 29124
0 1212 7 1 2 29293 1211
0 1213 7 1 2 29244 1212
0 1214 5 1 1 1213
0 1215 7 1 2 1191 1214
0 1216 5 1 1 1215
0 1217 7 1 2 29022 1216
0 1218 5 1 1 1217
0 1219 7 9 2 24640 26023
0 1220 7 4 2 25735 29141
0 1221 7 4 2 23004 26118
0 1222 7 1 2 22890 1147
0 1223 5 1 1 1222
0 1224 7 1 2 29311 1223
0 1225 5 1 1 1224
0 1226 7 5 2 24811 24152
0 1227 5 4 1 29315
0 1228 7 1 2 29320 29042
0 1229 5 1 1 1228
0 1230 7 6 2 25022 26119
0 1231 7 2 2 26405 29324
0 1232 5 1 1 29330
0 1233 7 1 2 1229 1232
0 1234 5 1 1 1233
0 1235 7 1 2 24940 1234
0 1236 5 1 1 1235
0 1237 7 1 2 1225 1236
0 1238 5 1 1 1237
0 1239 7 1 2 26215 1238
0 1240 5 1 1 1239
0 1241 7 1 2 24812 28578
0 1242 5 1 1 1241
0 1243 7 2 2 29043 1242
0 1244 5 1 1 29332
0 1245 7 1 2 27486 29333
0 1246 5 1 1 1245
0 1247 7 1 2 1240 1246
0 1248 5 1 1 1247
0 1249 7 1 2 23502 1248
0 1250 5 1 1 1249
0 1251 7 6 2 22891 26120
0 1252 5 6 1 29334
0 1253 7 3 2 27545 29044
0 1254 5 1 1 29346
0 1255 7 1 2 24316 26699
0 1256 5 2 1 1255
0 1257 7 1 2 24237 29349
0 1258 5 1 1 1257
0 1259 7 4 2 23503 26216
0 1260 5 2 1 29351
0 1261 7 1 2 23005 29355
0 1262 7 1 2 1258 1261
0 1263 5 1 1 1262
0 1264 7 1 2 1254 1263
0 1265 5 1 1 1264
0 1266 7 1 2 29335 1265
0 1267 5 1 1 1266
0 1268 7 1 2 1250 1267
0 1269 5 1 1 1268
0 1270 7 1 2 29307 1269
0 1271 5 1 1 1270
0 1272 7 1 2 26731 29127
0 1273 5 2 1 1272
0 1274 7 1 2 27574 29079
0 1275 5 1 1 1274
0 1276 7 1 2 29357 1275
0 1277 5 1 1 1276
0 1278 7 1 2 28494 1277
0 1279 5 1 1 1278
0 1280 7 1 2 27475 27684
0 1281 5 1 1 1280
0 1282 7 1 2 1279 1281
0 1283 5 1 1 1282
0 1284 7 10 2 23318 23760
0 1285 7 8 2 22383 22547
0 1286 5 2 1 29369
0 1287 7 3 2 23221 29370
0 1288 7 1 2 29359 29379
0 1289 7 1 2 1283 1288
0 1290 5 1 1 1289
0 1291 7 1 2 1271 1290
0 1292 5 1 1 1291
0 1293 7 1 2 23650 1292
0 1294 5 1 1 1293
0 1295 7 8 2 26121 29093
0 1296 5 1 1 29382
0 1297 7 2 2 23761 29383
0 1298 7 13 2 25170 25648
0 1299 7 2 2 28296 29392
0 1300 5 1 1 29405
0 1301 7 19 2 23222 23651
0 1302 7 3 2 28227 29407
0 1303 5 2 1 29426
0 1304 7 1 2 1300 29429
0 1305 5 2 1 1304
0 1306 7 1 2 22384 29431
0 1307 5 1 1 1306
0 1308 7 1 2 25649 29235
0 1309 5 1 1 1308
0 1310 7 1 2 1307 1309
0 1311 5 2 1 1310
0 1312 7 1 2 29390 29433
0 1313 5 1 1 1312
0 1314 7 7 2 22892 24153
0 1315 5 3 1 29435
0 1316 7 2 2 23504 29436
0 1317 5 1 1 29445
0 1318 7 1 2 1296 1317
0 1319 5 1 1 1318
0 1320 7 4 2 25650 28297
0 1321 7 3 2 24398 27715
0 1322 7 3 2 29447 29451
0 1323 5 1 1 29454
0 1324 7 1 2 25736 29455
0 1325 7 1 2 1319 1324
0 1326 5 1 1 1325
0 1327 7 1 2 1313 1326
0 1328 5 1 1 1327
0 1329 7 1 2 26812 1328
0 1330 5 1 1 1329
0 1331 7 1 2 1294 1330
0 1332 5 1 1 1331
0 1333 7 1 2 29298 1332
0 1334 5 1 1 1333
0 1335 7 5 2 25023 25171
0 1336 7 4 2 25651 29457
0 1337 7 2 2 28298 29462
0 1338 5 1 1 29466
0 1339 7 1 2 29430 1338
0 1340 5 3 1 1339
0 1341 7 1 2 22385 29468
0 1342 5 1 1 1341
0 1343 7 29 2 25024 25652
0 1344 7 2 2 29236 29471
0 1345 5 1 1 29500
0 1346 7 1 2 1342 1345
0 1347 5 1 1 1346
0 1348 7 1 2 26426 1347
0 1349 5 1 1 1348
0 1350 7 2 2 25653 26489
0 1351 7 1 2 29245 29502
0 1352 5 1 1 1351
0 1353 7 1 2 1349 1352
0 1354 5 1 1 1353
0 1355 7 1 2 29178 1354
0 1356 5 1 1 1355
0 1357 7 4 2 24154 26813
0 1358 5 2 1 29504
0 1359 7 1 2 29434 29505
0 1360 5 1 1 1359
0 1361 7 1 2 23762 1360
0 1362 7 1 2 1356 1361
0 1363 5 1 1 1362
0 1364 7 12 2 25463 24055
0 1365 7 6 2 22679 24813
0 1366 7 2 2 29510 29522
0 1367 5 1 1 29528
0 1368 7 5 2 23505 26024
0 1369 7 1 2 29530 27658
0 1370 5 1 1 1369
0 1371 7 1 2 1367 1370
0 1372 5 6 1 1371
0 1373 7 2 2 26427 29296
0 1374 5 9 1 29541
0 1375 7 9 2 24238 29542
0 1376 7 5 2 26490 27796
0 1377 5 2 1 29561
0 1378 7 1 2 29552 29566
0 1379 5 1 1 1378
0 1380 7 4 2 28608 26667
0 1381 5 1 1 29568
0 1382 7 1 2 1379 1381
0 1383 5 7 1 1382
0 1384 7 3 2 26122 29572
0 1385 5 1 1 29579
0 1386 7 10 2 25172 25260
0 1387 7 17 2 24399 24537
0 1388 5 1 1 29592
0 1389 7 2 2 25654 29593
0 1390 7 1 2 29582 29609
0 1391 7 1 2 29580 1390
0 1392 5 1 1 1391
0 1393 7 18 2 24239 24317
0 1394 5 1 1 29611
0 1395 7 4 2 26123 29612
0 1396 5 1 1 29629
0 1397 7 1 2 29508 1396
0 1398 5 1 1 1397
0 1399 7 6 2 22386 23652
0 1400 7 5 2 29218 29633
0 1401 5 1 1 29639
0 1402 7 3 2 23319 28335
0 1403 5 1 1 29644
0 1404 7 1 2 29408 29645
0 1405 5 1 1 1404
0 1406 7 1 2 1401 1405
0 1407 5 1 1 1406
0 1408 7 1 2 1398 1407
0 1409 5 1 1 1408
0 1410 7 1 2 25737 1409
0 1411 7 1 2 1392 1410
0 1412 5 1 1 1411
0 1413 7 1 2 29535 1412
0 1414 7 1 2 1363 1413
0 1415 5 1 1 1414
0 1416 7 1 2 1334 1415
0 1417 7 1 2 1218 1416
0 1418 5 1 1 1417
0 1419 7 1 2 26990 1418
0 1420 5 1 1 1419
0 1421 7 4 2 24814 26793
0 1422 5 1 1 29647
0 1423 7 4 2 22893 27598
0 1424 5 2 1 29651
0 1425 7 1 2 1422 29655
0 1426 5 10 1 1425
0 1427 7 8 2 22387 29409
0 1428 5 2 1 29667
0 1429 7 4 2 28932 29472
0 1430 5 1 1 29677
0 1431 7 1 2 29675 1430
0 1432 5 2 1 1431
0 1433 7 1 2 24318 29681
0 1434 5 1 1 1433
0 1435 7 12 2 23653 28193
0 1436 5 1 1 29683
0 1437 7 8 2 25655 28933
0 1438 7 1 2 29695 26549
0 1439 5 1 1 1438
0 1440 7 1 2 1436 1439
0 1441 5 1 1 1440
0 1442 7 1 2 25600 1441
0 1443 5 1 1 1442
0 1444 7 1 2 1434 1443
0 1445 5 2 1 1444
0 1446 7 1 2 29657 29703
0 1447 5 1 1 1446
0 1448 7 5 2 23006 26290
0 1449 7 1 2 29705 28464
0 1450 5 1 1 1449
0 1451 7 1 2 799 1450
0 1452 5 1 1 1451
0 1453 7 1 2 25464 1452
0 1454 5 1 1 1453
0 1455 7 2 2 25025 24319
0 1456 5 4 1 29710
0 1457 7 2 2 29711 29340
0 1458 5 1 1 29716
0 1459 7 1 2 24941 27621
0 1460 7 1 2 29717 1459
0 1461 5 1 1 1460
0 1462 7 1 2 1454 1461
0 1463 5 1 1 1462
0 1464 7 2 2 25601 29684
0 1465 7 1 2 1463 29718
0 1466 5 1 1 1465
0 1467 7 1 2 1447 1466
0 1468 5 1 1 1467
0 1469 7 1 2 29023 1468
0 1470 5 1 1 1469
0 1471 7 1 2 26124 29704
0 1472 5 1 1 1471
0 1473 7 1 2 29706 26615
0 1474 7 1 2 29685 1473
0 1475 5 1 1 1474
0 1476 7 1 2 1472 1475
0 1477 5 1 1 1476
0 1478 7 1 2 23506 1477
0 1479 5 1 1 1478
0 1480 7 5 2 26125 26291
0 1481 7 1 2 28545 29720
0 1482 7 1 2 29719 1481
0 1483 5 1 1 1482
0 1484 7 1 2 1479 1483
0 1485 5 1 1 1484
0 1486 7 1 2 22894 1485
0 1487 5 1 1 1486
0 1488 7 5 2 23654 27782
0 1489 7 3 2 22388 25602
0 1490 7 3 2 23007 23507
0 1491 5 1 1 29733
0 1492 7 1 2 29734 29721
0 1493 7 1 2 29730 1492
0 1494 7 1 2 29725 1493
0 1495 5 1 1 1494
0 1496 7 1 2 1487 1495
0 1497 5 1 1 1496
0 1498 7 1 2 29299 1497
0 1499 5 1 1 1498
0 1500 7 1 2 1470 1499
0 1501 5 1 1 1500
0 1502 7 1 2 23975 1501
0 1503 5 1 1 1502
0 1504 7 4 2 25942 27504
0 1505 7 2 2 26446 29736
0 1506 7 1 2 24320 27797
0 1507 5 1 1 1506
0 1508 7 2 2 26550 1507
0 1509 7 4 2 24641 25656
0 1510 7 2 2 28934 29744
0 1511 7 1 2 25603 29748
0 1512 7 1 2 29742 1511
0 1513 7 1 2 29740 1512
0 1514 5 1 1 1513
0 1515 7 1 2 1503 1514
0 1516 5 1 1 1515
0 1517 7 1 2 23871 1516
0 1518 5 1 1 1517
0 1519 7 21 2 25849 25943
0 1520 7 7 2 23655 29750
0 1521 7 1 2 23604 29712
0 1522 5 1 1 1521
0 1523 7 10 2 26551 1522
0 1524 5 2 1 29778
0 1525 7 1 2 29771 29779
0 1526 7 2 2 26126 27937
0 1527 7 2 2 26025 29048
0 1528 7 2 2 22680 29792
0 1529 7 1 2 29790 29794
0 1530 7 1 2 1525 1529
0 1531 5 1 1 1530
0 1532 7 1 2 1518 1531
0 1533 5 1 1 1532
0 1534 7 1 2 24240 1533
0 1535 5 1 1 1534
0 1536 7 2 2 23976 29531
0 1537 7 3 2 26292 26582
0 1538 7 1 2 29796 29798
0 1539 5 1 1 1538
0 1540 7 3 2 24056 29613
0 1541 7 5 2 25026 25465
0 1542 5 1 1 29804
0 1543 7 1 2 25944 29805
0 1544 7 1 2 29801 1543
0 1545 5 1 1 1544
0 1546 7 1 2 1539 1545
0 1547 5 1 1 1546
0 1548 7 1 2 26127 1547
0 1549 5 1 1 1548
0 1550 7 9 2 24155 26217
0 1551 5 1 1 29809
0 1552 7 20 2 25945 24057
0 1553 7 2 2 29818 26479
0 1554 7 1 2 29810 29838
0 1555 5 1 1 1554
0 1556 7 1 2 1549 1555
0 1557 5 1 1 1556
0 1558 7 1 2 24815 1557
0 1559 5 1 1 1558
0 1560 7 2 2 26026 26794
0 1561 7 3 2 22895 23977
0 1562 7 1 2 29842 29799
0 1563 7 1 2 29840 1562
0 1564 5 1 1 1563
0 1565 7 1 2 1559 1564
0 1566 5 1 1 1565
0 1567 7 1 2 29696 1566
0 1568 5 1 1 1567
0 1569 7 1 2 22896 26795
0 1570 5 2 1 1569
0 1571 7 1 2 24816 28495
0 1572 5 1 1 1571
0 1573 7 1 2 29845 1572
0 1574 5 7 1 1573
0 1575 7 1 2 29847 26583
0 1576 5 1 1 1575
0 1577 7 3 2 25027 27575
0 1578 7 1 2 28496 29854
0 1579 5 1 1 1578
0 1580 7 1 2 1576 1579
0 1581 5 1 1 1580
0 1582 7 1 2 26293 1581
0 1583 5 1 1 1582
0 1584 7 1 2 28520 486
0 1585 5 5 1 1584
0 1586 7 2 2 24321 27682
0 1587 7 1 2 29857 29862
0 1588 5 1 1 1587
0 1589 7 1 2 1583 1588
0 1590 5 1 1 1589
0 1591 7 20 2 23978 26027
0 1592 7 1 2 29864 29668
0 1593 7 1 2 1590 1592
0 1594 5 1 1 1593
0 1595 7 1 2 1568 1594
0 1596 5 1 1 1595
0 1597 7 1 2 24642 1596
0 1598 5 1 1 1597
0 1599 7 21 2 23979 24058
0 1600 7 3 2 22681 29884
0 1601 7 2 2 24817 26584
0 1602 7 4 2 24400 29393
0 1603 5 1 1 29910
0 1604 7 1 2 29676 1603
0 1605 5 3 1 1604
0 1606 7 1 2 29908 29914
0 1607 5 1 1 1606
0 1608 7 1 2 29686 29855
0 1609 5 1 1 1608
0 1610 7 1 2 1607 1609
0 1611 5 1 1 1610
0 1612 7 1 2 26294 1611
0 1613 5 1 1 1612
0 1614 7 1 2 29687 29863
0 1615 5 1 1 1614
0 1616 7 1 2 1613 1615
0 1617 5 1 1 1616
0 1618 7 1 2 27599 1617
0 1619 5 1 1 1618
0 1620 7 6 2 22389 24818
0 1621 7 2 2 29917 29410
0 1622 7 1 2 28615 29923
0 1623 7 1 2 29856 1622
0 1624 5 1 1 1623
0 1625 7 1 2 1619 1624
0 1626 5 1 1 1625
0 1627 7 1 2 29905 1626
0 1628 5 1 1 1627
0 1629 7 1 2 1598 1628
0 1630 5 1 1 1629
0 1631 7 1 2 23872 1630
0 1632 5 1 1 1631
0 1633 7 3 2 26295 27938
0 1634 7 7 2 26028 29751
0 1635 7 5 2 22682 23656
0 1636 7 1 2 29935 26585
0 1637 7 1 2 29928 1636
0 1638 7 1 2 29925 1637
0 1639 7 1 2 29384 1638
0 1640 5 1 1 1639
0 1641 7 1 2 1632 1640
0 1642 5 1 1 1641
0 1643 7 1 2 23605 1642
0 1644 5 1 1 1643
0 1645 7 4 2 23873 26218
0 1646 7 21 2 24059 24156
0 1647 7 16 2 25466 29944
0 1648 7 1 2 29965 29523
0 1649 5 1 1 1648
0 1650 7 8 2 26029 29848
0 1651 7 1 2 24643 29981
0 1652 5 1 1 1651
0 1653 7 1 2 1649 1652
0 1654 5 3 1 1653
0 1655 7 1 2 29989 29915
0 1656 5 1 1 1655
0 1657 7 1 2 28497 29300
0 1658 5 2 1 1657
0 1659 7 1 2 25467 29341
0 1660 5 1 1 1659
0 1661 7 2 2 29321 1660
0 1662 5 5 1 29994
0 1663 7 1 2 29996 29024
0 1664 5 1 1 1663
0 1665 7 1 2 29992 1664
0 1666 5 1 1 1665
0 1667 7 1 2 29128 29688
0 1668 7 1 2 1666 1667
0 1669 5 1 1 1668
0 1670 7 1 2 1656 1669
0 1671 5 1 1 1670
0 1672 7 1 2 23008 1671
0 1673 5 1 1 1672
0 1674 7 4 2 22683 25468
0 1675 7 2 2 29945 30001
0 1676 5 2 1 30005
0 1677 7 1 2 29301 29858
0 1678 5 1 1 1677
0 1679 7 1 2 30007 1678
0 1680 5 1 1 1679
0 1681 7 4 2 22390 24942
0 1682 7 3 2 27783 30009
0 1683 7 1 2 25604 23657
0 1684 7 1 2 26296 1683
0 1685 7 1 2 30013 1684
0 1686 7 1 2 1680 1685
0 1687 5 1 1 1686
0 1688 7 1 2 1673 1687
0 1689 5 1 1 1688
0 1690 7 1 2 23980 1689
0 1691 5 1 1 1690
0 1692 7 3 2 25469 25657
0 1693 7 2 2 25173 30016
0 1694 7 1 2 29819 30019
0 1695 7 15 2 24644 24819
0 1696 5 1 1 30021
0 1697 7 2 2 24401 30022
0 1698 7 1 2 28611 30036
0 1699 7 1 2 1694 1698
0 1700 5 1 1 1699
0 1701 7 1 2 1691 1700
0 1702 5 1 1 1701
0 1703 7 1 2 29940 1702
0 1704 5 1 1 1703
0 1705 7 1 2 1644 1704
0 1706 7 1 2 1535 1705
0 1707 5 1 1 1706
0 1708 7 1 2 28103 1707
0 1709 5 1 1 1708
0 1710 7 3 2 25261 25605
0 1711 7 4 2 24820 24060
0 1712 7 1 2 29271 30041
0 1713 7 1 2 30038 1712
0 1714 7 6 2 23508 27447
0 1715 7 1 2 30045 29678
0 1716 7 1 2 1713 1715
0 1717 5 1 1 1716
0 1718 7 2 2 26219 27798
0 1719 5 1 1 30051
0 1720 7 1 2 26482 1719
0 1721 5 1 1 1720
0 1722 7 1 2 22897 1721
0 1723 5 1 1 1722
0 1724 7 1 2 22898 26586
0 1725 5 3 1 1724
0 1726 7 1 2 23078 23509
0 1727 7 1 2 30053 1726
0 1728 5 1 1 1727
0 1729 7 1 2 1723 1728
0 1730 5 1 1 1729
0 1731 7 1 2 23606 1730
0 1732 5 1 1 1731
0 1733 7 1 2 26466 27487
0 1734 7 1 2 26705 1733
0 1735 5 1 1 1734
0 1736 7 1 2 1732 1735
0 1737 5 1 1 1736
0 1738 7 4 2 26128 29302
0 1739 7 3 2 23658 29142
0 1740 5 1 1 30060
0 1741 7 1 2 30056 30061
0 1742 7 1 2 1737 1741
0 1743 5 1 1 1742
0 1744 7 1 2 1717 1743
0 1745 5 1 1 1744
0 1746 7 1 2 26297 1745
0 1747 5 1 1 1746
0 1748 7 2 2 24241 26608
0 1749 5 1 1 30063
0 1750 7 1 2 27566 807
0 1751 5 1 1 1750
0 1752 7 1 2 25606 1751
0 1753 5 1 1 1752
0 1754 7 1 2 1749 1753
0 1755 5 1 1 1754
0 1756 7 2 2 24157 29594
0 1757 7 12 2 22684 25174
0 1758 7 4 2 24821 25262
0 1759 7 2 2 30067 30079
0 1760 7 2 2 23510 24061
0 1761 7 2 2 25658 24322
0 1762 7 1 2 30085 30087
0 1763 7 1 2 30083 1762
0 1764 7 1 2 30065 1763
0 1765 7 1 2 1755 1764
0 1766 5 1 1 1765
0 1767 7 1 2 1747 1766
0 1768 5 1 1 1767
0 1769 7 1 2 26935 1768
0 1770 5 1 1 1769
0 1771 7 4 2 22899 25607
0 1772 5 3 1 30089
0 1773 7 1 2 29707 26623
0 1774 5 1 1 1773
0 1775 7 1 2 30093 1774
0 1776 5 1 1 1775
0 1777 7 1 2 24158 1776
0 1778 5 1 1 1777
0 1779 7 5 2 24822 26129
0 1780 5 1 1 30096
0 1781 7 1 2 30097 29780
0 1782 5 1 1 1781
0 1783 7 1 2 1778 1782
0 1784 5 1 1 1783
0 1785 7 1 2 24242 1784
0 1786 5 1 1 1785
0 1787 7 2 2 23607 24159
0 1788 7 1 2 24823 30101
0 1789 7 1 2 29800 1788
0 1790 5 1 1 1789
0 1791 7 1 2 1786 1790
0 1792 5 1 1 1791
0 1793 7 3 2 27405 29511
0 1794 7 1 2 29640 30103
0 1795 5 1 1 1794
0 1796 7 13 2 23659 25850
0 1797 7 2 2 23223 30106
0 1798 7 3 2 22548 28868
0 1799 7 3 2 30119 30121
0 1800 7 1 2 24402 29512
0 1801 7 1 2 30124 1800
0 1802 5 1 1 1801
0 1803 7 1 2 1795 1802
0 1804 5 1 1 1803
0 1805 7 1 2 1792 1804
0 1806 5 1 1 1805
0 1807 7 15 2 25659 23874
0 1808 7 3 2 26030 30127
0 1809 7 4 2 24403 23079
0 1810 7 2 2 29583 30145
0 1811 7 2 2 22900 27448
0 1812 7 1 2 30149 30151
0 1813 7 1 2 30142 1812
0 1814 7 1 2 26829 1813
0 1815 5 1 1 1814
0 1816 7 1 2 1806 1815
0 1817 5 1 1 1816
0 1818 7 1 2 25946 1817
0 1819 5 1 1 1818
0 1820 7 1 2 25338 1819
0 1821 7 1 2 1770 1820
0 1822 7 1 2 1709 1821
0 1823 5 1 1 1822
0 1824 7 2 2 24943 29080
0 1825 5 2 1 30153
0 1826 7 1 2 26467 30154
0 1827 5 1 1 1826
0 1828 7 2 2 26527 28490
0 1829 5 1 1 30157
0 1830 7 1 2 1827 1829
0 1831 5 1 1 1830
0 1832 7 1 2 28846 1831
0 1833 5 1 1 1832
0 1834 7 21 2 24645 25947
0 1835 5 1 1 30159
0 1836 7 1 2 30160 29094
0 1837 7 1 2 28528 1836
0 1838 5 1 1 1837
0 1839 7 1 2 1833 1838
0 1840 5 1 1 1839
0 1841 7 1 2 26220 1840
0 1842 5 1 1 1841
0 1843 7 2 2 29095 26406
0 1844 7 3 2 22685 23080
0 1845 7 2 2 23981 30182
0 1846 5 1 1 30185
0 1847 7 1 2 23009 30161
0 1848 5 1 1 1847
0 1849 7 1 2 1846 1848
0 1850 5 1 1 1849
0 1851 7 1 2 30180 1850
0 1852 5 1 1 1851
0 1853 7 1 2 1842 1852
0 1854 5 1 1 1853
0 1855 7 1 2 26130 1854
0 1856 5 1 1 1855
0 1857 7 1 2 28847 29347
0 1858 5 1 1 1857
0 1859 7 1 2 30162 29506
0 1860 5 1 1 1859
0 1861 7 1 2 1858 1860
0 1862 5 1 1 1861
0 1863 7 1 2 29049 1862
0 1864 5 1 1 1863
0 1865 7 1 2 1856 1864
0 1866 5 1 1 1865
0 1867 7 1 2 26031 1866
0 1868 5 1 1 1867
0 1869 7 10 2 25948 24160
0 1870 7 1 2 30187 29529
0 1871 7 1 2 26814 1870
0 1872 5 1 1 1871
0 1873 7 1 2 1868 1872
0 1874 5 1 1 1873
0 1875 7 5 2 25851 27939
0 1876 7 1 2 23660 30197
0 1877 7 1 2 1874 1876
0 1878 5 1 1 1877
0 1879 7 4 2 25175 23982
0 1880 7 6 2 25470 23875
0 1881 7 3 2 23608 25660
0 1882 7 1 2 30206 30212
0 1883 7 1 2 30202 1882
0 1884 7 5 2 24062 26221
0 1885 7 2 2 30215 26694
0 1886 7 1 2 30220 30037
0 1887 7 1 2 1883 1886
0 1888 5 1 1 1887
0 1889 7 1 2 1878 1888
0 1890 5 1 1 1889
0 1891 7 1 2 28104 1890
0 1892 5 1 1 1891
0 1893 7 6 2 25852 28105
0 1894 5 1 1 30222
0 1895 7 3 2 27940 30223
0 1896 7 2 2 26298 26706
0 1897 5 1 1 30231
0 1898 7 1 2 26131 30232
0 1899 5 1 1 1898
0 1900 7 1 2 1244 1899
0 1901 5 1 1 1900
0 1902 7 1 2 23010 1901
0 1903 5 1 1 1902
0 1904 7 1 2 28584 26407
0 1905 5 2 1 1904
0 1906 7 1 2 22901 24323
0 1907 5 1 1 1906
0 1908 7 1 2 30233 1907
0 1909 5 1 1 1908
0 1910 7 1 2 26132 1909
0 1911 5 1 1 1910
0 1912 7 1 2 1903 1911
0 1913 5 1 1 1912
0 1914 7 1 2 29865 1913
0 1915 5 1 1 1914
0 1916 7 4 2 24161 29820
0 1917 7 2 2 24824 26428
0 1918 5 1 1 30239
0 1919 7 1 2 29567 1918
0 1920 5 3 1 1919
0 1921 7 1 2 30235 30241
0 1922 5 1 1 1921
0 1923 7 1 2 1915 1922
0 1924 5 1 1 1923
0 1925 7 1 2 23511 1924
0 1926 5 1 1 1925
0 1927 7 5 2 23011 24162
0 1928 5 1 1 30244
0 1929 7 1 2 30245 29081
0 1930 5 1 1 1929
0 1931 7 12 2 24825 25028
0 1932 7 1 2 26133 30249
0 1933 5 1 1 1932
0 1934 7 1 2 29442 1933
0 1935 5 3 1 1934
0 1936 7 1 2 26429 30261
0 1937 5 1 1 1936
0 1938 7 3 2 24826 25608
0 1939 5 1 1 30264
0 1940 7 2 2 28574 30265
0 1941 5 1 1 30267
0 1942 7 1 2 1937 1941
0 1943 7 1 2 1930 1942
0 1944 5 1 1 1943
0 1945 7 1 2 25471 1944
0 1946 5 1 1 1945
0 1947 7 3 2 24827 23609
0 1948 7 1 2 26695 26528
0 1949 7 1 2 30269 1948
0 1950 5 1 1 1949
0 1951 7 1 2 1946 1950
0 1952 5 1 1 1951
0 1953 7 1 2 29821 1952
0 1954 5 1 1 1953
0 1955 7 1 2 29350 1897
0 1956 5 1 1 1955
0 1957 7 7 2 23983 26134
0 1958 7 2 2 23012 26032
0 1959 7 2 2 30272 30279
0 1960 7 1 2 22902 30281
0 1961 7 1 2 1956 1960
0 1962 5 1 1 1961
0 1963 7 1 2 1954 1962
0 1964 7 1 2 1926 1963
0 1965 5 1 1 1964
0 1966 7 1 2 30228 1965
0 1967 5 1 1 1966
0 1968 7 1 2 22686 1967
0 1969 5 1 1 1968
0 1970 7 9 2 26033 29336
0 1971 7 3 2 26962 30283
0 1972 5 1 1 30292
0 1973 7 1 2 26616 30293
0 1974 5 1 1 1973
0 1975 7 2 2 24828 29885
0 1976 7 5 2 23610 25853
0 1977 7 1 2 29806 30297
0 1978 7 1 2 30295 1977
0 1979 5 1 1 1978
0 1980 7 1 2 1974 1979
0 1981 5 1 1 1980
0 1982 7 1 2 29708 1981
0 1983 5 1 1 1982
0 1984 7 1 2 29067 29562
0 1985 5 1 1 1984
0 1986 7 1 2 25472 30240
0 1987 5 1 1 1986
0 1988 7 1 2 1985 1987
0 1989 5 1 1 1988
0 1990 7 8 2 25854 24063
0 1991 7 1 2 30273 30302
0 1992 7 1 2 1989 1991
0 1993 5 1 1 1992
0 1994 7 1 2 1983 1993
0 1995 5 1 1 1994
0 1996 7 1 2 29143 1995
0 1997 5 1 1 1996
0 1998 7 16 2 28106 27941
0 1999 7 20 2 25949 26034
0 2000 7 4 2 25855 30326
0 2001 7 4 2 30310 30346
0 2002 5 1 1 30350
0 2003 7 8 2 26135 29050
0 2004 5 2 1 30354
0 2005 7 1 2 30355 29781
0 2006 7 1 2 30351 2005
0 2007 5 1 1 2006
0 2008 7 1 2 24646 2007
0 2009 7 1 2 1997 2008
0 2010 5 1 1 2009
0 2011 7 1 2 23661 2010
0 2012 7 1 2 1969 2011
0 2013 5 1 1 2012
0 2014 7 7 2 24163 29096
0 2015 7 3 2 25950 28753
0 2016 5 1 1 30371
0 2017 7 1 2 30364 30372
0 2018 5 1 1 2017
0 2019 7 4 2 24647 25473
0 2020 7 8 2 24829 23320
0 2021 7 1 2 30274 30378
0 2022 7 1 2 30374 2021
0 2023 5 1 1 2022
0 2024 7 1 2 2018 2023
0 2025 5 1 1 2024
0 2026 7 1 2 24538 2025
0 2027 5 1 1 2026
0 2028 7 3 2 22549 30023
0 2029 7 5 2 25263 23984
0 2030 7 1 2 26780 30389
0 2031 7 1 2 30386 2030
0 2032 5 1 1 2031
0 2033 7 1 2 2027 2032
0 2034 5 1 1 2033
0 2035 7 1 2 24064 2034
0 2036 5 1 1 2035
0 2037 7 4 2 29532 30275
0 2038 5 2 1 30394
0 2039 7 8 2 22903 25264
0 2040 7 2 2 27449 30400
0 2041 7 1 2 30395 30408
0 2042 5 1 1 2041
0 2043 7 1 2 2036 2042
0 2044 5 1 1 2043
0 2045 7 2 2 25029 26430
0 2046 5 2 1 30410
0 2047 7 2 2 26504 30412
0 2048 5 1 1 30414
0 2049 7 1 2 28935 30128
0 2050 7 1 2 2048 2049
0 2051 7 1 2 2044 2050
0 2052 5 1 1 2051
0 2053 7 1 2 2013 2052
0 2054 5 1 1 2053
0 2055 7 1 2 24243 2054
0 2056 5 1 1 2055
0 2057 7 4 2 28585 27476
0 2058 7 1 2 27600 30416
0 2059 5 1 1 2058
0 2060 7 1 2 29997 29028
0 2061 5 1 1 2060
0 2062 7 1 2 2059 2061
0 2063 5 1 1 2062
0 2064 7 1 2 24065 30125
0 2065 7 1 2 2063 2064
0 2066 5 1 1 2065
0 2067 7 1 2 28299 30068
0 2068 7 1 2 28529 2067
0 2069 7 1 2 30143 2068
0 2070 7 1 2 29849 2069
0 2071 5 1 1 2070
0 2072 7 1 2 2066 2071
0 2073 5 1 1 2072
0 2074 7 1 2 26222 2073
0 2075 5 1 1 2074
0 2076 7 3 2 27450 29982
0 2077 5 1 1 30420
0 2078 7 4 2 26299 28613
0 2079 7 12 2 25265 23876
0 2080 5 1 1 30427
0 2081 7 1 2 30428 29394
0 2082 7 1 2 30423 2081
0 2083 7 1 2 30421 2082
0 2084 5 1 1 2083
0 2085 7 1 2 2075 2084
0 2086 5 1 1 2085
0 2087 7 1 2 23985 2086
0 2088 5 1 1 2087
0 2089 7 5 2 24539 23013
0 2090 7 1 2 24830 30069
0 2091 7 2 2 30439 2090
0 2092 7 7 2 25266 25661
0 2093 7 1 2 29946 30446
0 2094 7 1 2 30444 2093
0 2095 5 1 1 2094
0 2096 7 1 2 28869 27466
0 2097 7 5 2 22550 23662
0 2098 7 17 2 26035 26136
0 2099 7 1 2 30458 26587
0 2100 7 1 2 30453 2099
0 2101 7 1 2 2096 2100
0 2102 5 1 1 2101
0 2103 7 1 2 2095 2102
0 2104 5 1 1 2103
0 2105 7 1 2 26300 2104
0 2106 5 1 1 2105
0 2107 7 5 2 24066 29811
0 2108 7 2 2 30475 30447
0 2109 7 1 2 24831 27451
0 2110 7 1 2 27716 2109
0 2111 7 1 2 30480 2110
0 2112 5 1 1 2111
0 2113 7 1 2 2106 2112
0 2114 5 1 1 2113
0 2115 7 1 2 23611 2114
0 2116 5 1 1 2115
0 2117 7 1 2 30445 30481
0 2118 5 1 1 2117
0 2119 7 1 2 2116 2118
0 2120 5 1 1 2119
0 2121 7 1 2 25951 30207
0 2122 7 1 2 2120 2121
0 2123 5 1 1 2122
0 2124 7 1 2 2088 2123
0 2125 5 1 1 2124
0 2126 7 1 2 24404 2125
0 2127 5 1 1 2126
0 2128 7 1 2 26588 30294
0 2129 5 1 1 2128
0 2130 7 2 2 23986 27799
0 2131 7 3 2 25856 30216
0 2132 7 1 2 29342 30484
0 2133 7 1 2 30482 2132
0 2134 5 1 1 2133
0 2135 7 1 2 2129 2134
0 2136 5 1 1 2135
0 2137 7 1 2 26301 2136
0 2138 5 1 1 2137
0 2139 7 1 2 29886 28586
0 2140 7 8 2 25857 24164
0 2141 7 1 2 30487 26668
0 2142 7 1 2 2139 2141
0 2143 5 1 1 2142
0 2144 7 1 2 2138 2143
0 2145 5 1 1 2144
0 2146 7 1 2 23612 2145
0 2147 5 1 1 2146
0 2148 7 1 2 23014 1458
0 2149 5 1 1 2148
0 2150 7 2 2 24165 26547
0 2151 5 1 1 30495
0 2152 7 1 2 24944 2151
0 2153 5 1 1 2152
0 2154 7 4 2 25609 26936
0 2155 7 1 2 30217 30497
0 2156 7 1 2 2153 2155
0 2157 7 1 2 2149 2156
0 2158 5 1 1 2157
0 2159 7 1 2 2147 2158
0 2160 5 1 1 2159
0 2161 7 1 2 25474 2160
0 2162 5 1 1 2161
0 2163 7 1 2 26937 30250
0 2164 7 1 2 30476 2163
0 2165 7 1 2 28537 2164
0 2166 5 1 1 2165
0 2167 7 1 2 2162 2166
0 2168 5 1 1 2167
0 2169 7 1 2 24648 29641
0 2170 7 1 2 2168 2169
0 2171 5 1 1 2170
0 2172 7 1 2 23380 2171
0 2173 7 1 2 2127 2172
0 2174 7 1 2 2056 2173
0 2175 7 1 2 1892 2174
0 2176 5 1 1 2175
0 2177 7 1 2 1823 2176
0 2178 5 1 1 2177
0 2179 7 2 2 24649 24067
0 2180 7 9 2 23877 28107
0 2181 7 2 2 25662 29553
0 2182 7 2 2 25176 27791
0 2183 7 1 2 30512 30514
0 2184 5 1 1 2183
0 2185 7 2 2 22904 26635
0 2186 5 3 1 30516
0 2187 7 1 2 30155 1135
0 2188 5 1 1 2187
0 2189 7 1 2 26223 2188
0 2190 5 1 1 2189
0 2191 7 1 2 30518 2190
0 2192 5 2 1 2191
0 2193 7 1 2 29669 30521
0 2194 5 1 1 2193
0 2195 7 1 2 2184 2194
0 2196 5 1 1 2195
0 2197 7 1 2 25475 2196
0 2198 5 1 1 2197
0 2199 7 2 2 23512 28936
0 2200 7 1 2 30513 30523
0 2201 5 1 1 2200
0 2202 7 4 2 23613 23663
0 2203 7 6 2 25030 23224
0 2204 5 1 1 30529
0 2205 7 2 2 30525 30530
0 2206 7 1 2 30010 28415
0 2207 7 1 2 30535 2206
0 2208 5 1 1 2207
0 2209 7 1 2 2201 2208
0 2210 5 1 1 2209
0 2211 7 1 2 24832 2210
0 2212 5 1 1 2211
0 2213 7 1 2 2198 2212
0 2214 5 1 1 2213
0 2215 7 1 2 24166 2214
0 2216 5 1 1 2215
0 2217 7 5 2 26684 28575
0 2218 5 4 1 30537
0 2219 7 1 2 28431 30542
0 2220 5 1 1 2219
0 2221 7 2 2 30011 30251
0 2222 7 1 2 29411 30546
0 2223 7 1 2 2220 2222
0 2224 5 1 1 2223
0 2225 7 1 2 2216 2224
0 2226 5 1 1 2225
0 2227 7 1 2 30503 2226
0 2228 5 1 1 2227
0 2229 7 7 2 22905 25663
0 2230 7 4 2 25177 25476
0 2231 7 2 2 30548 30555
0 2232 7 4 2 25031 24244
0 2233 5 5 1 30561
0 2234 7 1 2 26749 28300
0 2235 7 1 2 30565 2234
0 2236 7 1 2 30559 2235
0 2237 5 1 1 2236
0 2238 7 1 2 30562 26556
0 2239 7 1 2 29427 2238
0 2240 5 1 1 2239
0 2241 7 1 2 2237 2240
0 2242 5 1 1 2241
0 2243 7 1 2 25610 2242
0 2244 5 1 1 2243
0 2245 7 1 2 29097 29428
0 2246 5 1 1 2245
0 2247 7 10 2 24540 25178
0 2248 7 5 2 22906 25032
0 2249 7 2 2 30570 30580
0 2250 7 3 2 25267 23614
0 2251 7 1 2 30017 30587
0 2252 7 1 2 30585 2251
0 2253 5 1 1 2252
0 2254 7 1 2 2246 2253
0 2255 5 1 1 2254
0 2256 7 1 2 24245 2255
0 2257 5 1 1 2256
0 2258 7 1 2 2244 2257
0 2259 5 1 1 2258
0 2260 7 1 2 24324 2259
0 2261 5 1 1 2260
0 2262 7 3 2 23081 24246
0 2263 5 2 1 30590
0 2264 7 1 2 30593 26613
0 2265 7 1 2 1939 30556
0 2266 7 1 2 2264 2265
0 2267 7 9 2 22907 26224
0 2268 5 1 1 30595
0 2269 7 1 2 26302 2268
0 2270 7 1 2 29448 2269
0 2271 7 1 2 2266 2270
0 2272 5 1 1 2271
0 2273 7 2 2 23321 23664
0 2274 7 6 2 23225 30604
0 2275 7 3 2 22551 23513
0 2276 7 1 2 24833 30612
0 2277 7 1 2 26685 2276
0 2278 7 1 2 30606 2277
0 2279 5 1 1 2278
0 2280 7 1 2 2272 2279
0 2281 7 1 2 2261 2280
0 2282 5 1 1 2281
0 2283 7 1 2 24405 2282
0 2284 5 1 1 2283
0 2285 7 1 2 23514 30242
0 2286 5 1 1 2285
0 2287 7 1 2 24325 26536
0 2288 5 1 1 2287
0 2289 7 1 2 2286 2288
0 2290 5 1 1 2289
0 2291 7 1 2 24247 29642
0 2292 7 1 2 2290 2291
0 2293 5 1 1 2292
0 2294 7 1 2 2284 2293
0 2295 5 1 1 2294
0 2296 7 1 2 30488 2295
0 2297 5 1 1 2296
0 2298 7 1 2 2228 2297
0 2299 5 1 1 2298
0 2300 7 1 2 30501 2299
0 2301 5 1 1 2300
0 2302 7 9 2 24650 23226
0 2303 7 4 2 25268 30615
0 2304 7 1 2 29966 30624
0 2305 5 1 1 2304
0 2306 7 4 2 23322 23515
0 2307 7 3 2 30459 30628
0 2308 7 1 2 30070 30632
0 2309 5 1 1 2308
0 2310 7 1 2 2305 2309
0 2311 5 1 1 2310
0 2312 7 1 2 22552 2311
0 2313 5 1 1 2312
0 2314 7 21 2 24541 23227
0 2315 7 1 2 29967 28870
0 2316 5 1 1 2315
0 2317 7 2 2 23516 28754
0 2318 7 1 2 30460 30656
0 2319 5 1 1 2318
0 2320 7 1 2 2316 2319
0 2321 5 1 1 2320
0 2322 7 1 2 30635 2321
0 2323 5 1 1 2322
0 2324 7 1 2 2313 2323
0 2325 5 1 1 2324
0 2326 7 1 2 22391 2325
0 2327 5 1 1 2326
0 2328 7 2 2 22687 23228
0 2329 7 2 2 28336 30658
0 2330 7 1 2 30633 30660
0 2331 5 1 1 2330
0 2332 7 1 2 2327 2331
0 2333 5 1 1 2332
0 2334 7 1 2 24248 29082
0 2335 5 1 1 2334
0 2336 7 1 2 28478 2335
0 2337 5 1 1 2336
0 2338 7 1 2 2333 2337
0 2339 5 1 1 2338
0 2340 7 3 2 22688 29144
0 2341 7 2 2 24249 27477
0 2342 7 8 2 23082 26036
0 2343 5 1 1 30667
0 2344 7 1 2 27679 30668
0 2345 7 1 2 30665 2344
0 2346 7 1 2 30662 2345
0 2347 5 1 1 2346
0 2348 7 1 2 2339 2347
0 2349 5 1 1 2348
0 2350 7 1 2 23878 2349
0 2351 5 1 1 2350
0 2352 7 6 2 23517 30461
0 2353 7 5 2 22689 25858
0 2354 7 1 2 30681 27942
0 2355 7 1 2 30675 2354
0 2356 5 1 1 2355
0 2357 7 13 2 22392 24651
0 2358 7 2 2 30686 30531
0 2359 7 2 2 23879 24068
0 2360 7 1 2 26491 28521
0 2361 7 1 2 30701 2360
0 2362 7 1 2 30699 2361
0 2363 5 1 1 2362
0 2364 7 1 2 2356 2363
0 2365 5 1 1 2364
0 2366 7 1 2 26225 2365
0 2367 5 1 1 2366
0 2368 7 8 2 24069 24250
0 2369 7 2 2 23880 30703
0 2370 7 1 2 30711 28596
0 2371 7 1 2 30700 2370
0 2372 5 1 1 2371
0 2373 7 1 2 2367 2372
0 2374 5 1 1 2373
0 2375 7 1 2 28108 2374
0 2376 5 1 1 2375
0 2377 7 2 2 25477 26226
0 2378 5 1 1 30713
0 2379 7 1 2 25033 28894
0 2380 5 1 1 2379
0 2381 7 1 2 2378 2380
0 2382 5 1 1 2381
0 2383 7 1 2 29947 27406
0 2384 7 1 2 2382 2383
0 2385 7 1 2 29145 2384
0 2386 5 1 1 2385
0 2387 7 1 2 2376 2386
0 2388 5 1 1 2387
0 2389 7 1 2 24834 2388
0 2390 5 1 1 2389
0 2391 7 4 2 26037 26303
0 2392 5 1 1 30715
0 2393 7 2 2 22908 30716
0 2394 7 1 2 30657 30719
0 2395 5 1 1 2394
0 2396 7 3 2 24652 29614
0 2397 7 4 2 23083 23323
0 2398 7 1 2 30724 29513
0 2399 7 1 2 30721 2398
0 2400 5 1 1 2399
0 2401 7 1 2 2395 2400
0 2402 5 1 1 2401
0 2403 7 1 2 22553 2402
0 2404 5 1 1 2403
0 2405 7 1 2 23324 30046
0 2406 7 1 2 30720 2405
0 2407 5 1 1 2406
0 2408 7 1 2 2404 2407
0 2409 5 1 1 2408
0 2410 7 1 2 27943 2409
0 2411 5 1 1 2410
0 2412 7 9 2 23084 25269
0 2413 7 5 2 23229 25478
0 2414 7 1 2 30728 30737
0 2415 7 1 2 28063 2414
0 2416 7 1 2 29802 2415
0 2417 5 1 1 2416
0 2418 7 1 2 2411 2417
0 2419 5 1 1 2418
0 2420 7 1 2 24167 30298
0 2421 7 1 2 2419 2420
0 2422 5 1 1 2421
0 2423 7 1 2 2390 2422
0 2424 7 1 2 2351 2423
0 2425 5 1 1 2424
0 2426 7 1 2 23665 2425
0 2427 5 1 1 2426
0 2428 7 4 2 23666 26038
0 2429 7 2 2 28498 30742
0 2430 7 1 2 30746 30663
0 2431 5 1 1 2430
0 2432 7 2 2 24653 28109
0 2433 7 1 2 29968 30748
0 2434 7 1 2 29916 2433
0 2435 5 1 1 2434
0 2436 7 1 2 2431 2435
0 2437 5 1 1 2436
0 2438 7 1 2 23881 2437
0 2439 5 1 1 2438
0 2440 7 5 2 24168 30303
0 2441 7 2 2 30375 30750
0 2442 7 1 2 30755 29456
0 2443 5 1 1 2442
0 2444 7 1 2 2439 2443
0 2445 5 1 1 2444
0 2446 7 1 2 24835 26642
0 2447 7 1 2 2445 2446
0 2448 5 1 1 2447
0 2449 7 2 2 28014 29595
0 2450 7 1 2 30757 30751
0 2451 7 1 2 28382 30560
0 2452 7 1 2 2450 2451
0 2453 5 1 1 2452
0 2454 7 1 2 2448 2453
0 2455 7 1 2 2427 2454
0 2456 5 1 1 2455
0 2457 7 1 2 23015 2456
0 2458 5 1 1 2457
0 2459 7 7 2 23615 26227
0 2460 7 1 2 29051 30759
0 2461 7 1 2 30489 2460
0 2462 7 1 2 28110 2461
0 2463 7 1 2 29926 2462
0 2464 5 1 1 2463
0 2465 7 1 2 27680 29348
0 2466 5 1 1 2465
0 2467 7 1 2 28499 30522
0 2468 5 1 1 2467
0 2469 7 1 2 2466 2468
0 2470 5 1 1 2469
0 2471 7 1 2 23882 29146
0 2472 7 1 2 2470 2471
0 2473 5 1 1 2472
0 2474 7 1 2 2464 2473
0 2475 5 1 1 2474
0 2476 7 1 2 26039 29936
0 2477 7 1 2 2475 2476
0 2478 5 1 1 2477
0 2479 7 2 2 22690 27944
0 2480 7 2 2 22909 30766
0 2481 7 7 2 25859 26040
0 2482 7 1 2 26732 30770
0 2483 7 1 2 30768 2482
0 2484 5 1 1 2483
0 2485 7 7 2 23230 23883
0 2486 7 2 2 30777 30687
0 2487 7 1 2 30704 30784
0 2488 7 1 2 30243 2487
0 2489 5 1 1 2488
0 2490 7 1 2 2484 2489
0 2491 5 1 1 2490
0 2492 7 1 2 28111 2491
0 2493 5 1 1 2492
0 2494 7 8 2 22691 23884
0 2495 7 3 2 26041 30786
0 2496 7 3 2 22910 30794
0 2497 7 1 2 26815 30797
0 2498 7 1 2 29147 2497
0 2499 5 1 1 2498
0 2500 7 1 2 2493 2499
0 2501 5 1 1 2500
0 2502 7 1 2 23667 2501
0 2503 5 1 1 2502
0 2504 7 6 2 25179 30448
0 2505 7 1 2 30304 29596
0 2506 7 1 2 30024 2505
0 2507 7 1 2 30800 2506
0 2508 7 1 2 29573 2507
0 2509 5 1 1 2508
0 2510 7 1 2 2503 2509
0 2511 5 1 1 2510
0 2512 7 1 2 28636 2511
0 2513 5 1 1 2512
0 2514 7 1 2 2478 2513
0 2515 7 1 2 2458 2514
0 2516 7 1 2 2301 2515
0 2517 5 1 1 2516
0 2518 7 1 2 27064 2517
0 2519 5 1 1 2518
0 2520 7 5 2 26042 26963
0 2521 7 1 2 28500 30806
0 2522 5 1 1 2521
0 2523 7 3 2 25860 29887
0 2524 7 1 2 27601 30811
0 2525 5 1 1 2524
0 2526 7 2 2 2522 2525
0 2527 5 13 1 30814
0 2528 7 1 2 27488 26617
0 2529 5 1 1 2528
0 2530 7 1 2 22911 30566
0 2531 5 2 1 2530
0 2532 7 1 2 23616 26589
0 2533 7 1 2 30829 2532
0 2534 5 1 1 2533
0 2535 7 1 2 2529 2534
0 2536 5 1 1 2535
0 2537 7 1 2 26304 2536
0 2538 5 1 1 2537
0 2539 7 1 2 22912 26686
0 2540 5 1 1 2539
0 2541 7 1 2 2538 2540
0 2542 5 1 1 2541
0 2543 7 9 2 24654 23381
0 2544 5 1 1 30831
0 2545 7 1 2 30832 29643
0 2546 5 1 1 2545
0 2547 7 4 2 23382 23668
0 2548 7 1 2 27905 30840
0 2549 7 1 2 30122 2548
0 2550 5 1 1 2549
0 2551 7 1 2 2546 2550
0 2552 5 1 1 2551
0 2553 7 1 2 2542 2552
0 2554 5 1 1 2553
0 2555 7 1 2 22913 29574
0 2556 5 1 1 2555
0 2557 7 8 2 24836 23085
0 2558 7 1 2 30844 26816
0 2559 5 1 1 2558
0 2560 7 1 2 2556 2559
0 2561 5 1 1 2560
0 2562 7 6 2 22692 25339
0 2563 5 2 1 30852
0 2564 7 1 2 30853 28301
0 2565 7 1 2 29911 2564
0 2566 7 1 2 2561 2565
0 2567 5 1 1 2566
0 2568 7 1 2 2554 2567
0 2569 5 1 1 2568
0 2570 7 1 2 30816 2569
0 2571 5 1 1 2570
0 2572 7 1 2 25738 2571
0 2573 7 1 2 2519 2572
0 2574 7 1 2 2178 2573
0 2575 5 1 1 2574
0 2576 7 3 2 27043 30504
0 2577 5 1 1 30860
0 2578 7 1 2 30861 29990
0 2579 5 1 1 2578
0 2580 7 2 2 29948 27299
0 2581 7 1 2 30376 30863
0 2582 5 1 1 2581
0 2583 7 7 2 23885 28755
0 2584 7 1 2 30865 30676
0 2585 5 1 1 2584
0 2586 7 1 2 2582 2585
0 2587 5 1 1 2586
0 2588 7 1 2 24837 2587
0 2589 5 1 1 2588
0 2590 7 2 2 30401 29841
0 2591 7 1 2 30787 30872
0 2592 5 1 1 2591
0 2593 7 1 2 2589 2592
0 2594 5 1 1 2593
0 2595 7 1 2 24542 2594
0 2596 5 1 1 2595
0 2597 7 3 2 27602 30042
0 2598 7 4 2 24655 23886
0 2599 7 1 2 28092 30877
0 2600 7 1 2 30874 2599
0 2601 5 1 1 2600
0 2602 7 1 2 2596 2601
0 2603 5 1 1 2602
0 2604 7 1 2 27065 2603
0 2605 5 1 1 2604
0 2606 7 1 2 2579 2605
0 2607 5 2 1 2606
0 2608 7 1 2 26817 30881
0 2609 5 1 1 2608
0 2610 7 1 2 30008 29993
0 2611 5 1 1 2610
0 2612 7 1 2 22914 2611
0 2613 5 1 1 2612
0 2614 7 1 2 29648 29025
0 2615 5 1 1 2614
0 2616 7 1 2 2613 2615
0 2617 5 2 1 2616
0 2618 7 1 2 30862 30883
0 2619 5 1 1 2618
0 2620 7 3 2 22554 30429
0 2621 5 2 1 30885
0 2622 7 2 2 24543 27300
0 2623 5 1 1 30890
0 2624 7 2 2 30888 2623
0 2625 5 9 1 30892
0 2626 7 1 2 29658 30502
0 2627 7 1 2 30894 2626
0 2628 5 1 1 2627
0 2629 7 6 2 23518 23887
0 2630 7 2 2 30462 30903
0 2631 7 1 2 30909 30409
0 2632 5 1 1 2631
0 2633 7 1 2 2628 2632
0 2634 5 1 1 2633
0 2635 7 1 2 27066 2634
0 2636 5 1 1 2635
0 2637 7 1 2 2619 2636
0 2638 5 1 1 2637
0 2639 7 1 2 29554 2638
0 2640 5 1 1 2639
0 2641 7 1 2 2609 2640
0 2642 5 1 1 2641
0 2643 7 1 2 29395 2642
0 2644 5 1 1 2643
0 2645 7 2 2 28228 30788
0 2646 7 2 2 24070 29722
0 2647 7 1 2 26700 30913
0 2648 5 2 1 2647
0 2649 7 2 2 25034 26043
0 2650 5 1 1 30917
0 2651 7 2 2 26492 30918
0 2652 5 1 1 30919
0 2653 7 1 2 30915 2652
0 2654 5 2 1 2653
0 2655 7 1 2 23016 30921
0 2656 5 1 1 2655
0 2657 7 5 2 24945 26044
0 2658 7 1 2 30923 29083
0 2659 5 1 1 2658
0 2660 7 1 2 2656 2659
0 2661 5 1 1 2660
0 2662 7 1 2 26366 2661
0 2663 5 1 1 2662
0 2664 7 3 2 26045 26766
0 2665 7 1 2 30928 30417
0 2666 5 1 1 2665
0 2667 7 1 2 2663 2666
0 2668 5 1 1 2667
0 2669 7 1 2 22915 2668
0 2670 5 1 1 2669
0 2671 7 1 2 26533 30156
0 2672 5 2 1 2671
0 2673 7 1 2 26767 30931
0 2674 5 1 1 2673
0 2675 7 1 2 26367 30418
0 2676 5 1 1 2675
0 2677 7 1 2 2674 2676
0 2678 5 1 1 2677
0 2679 7 1 2 30463 2678
0 2680 5 1 1 2679
0 2681 7 1 2 2670 2680
0 2682 5 1 1 2681
0 2683 7 1 2 23519 2682
0 2684 5 1 1 2683
0 2685 7 1 2 24946 26902
0 2686 7 1 2 30284 2685
0 2687 7 1 2 29045 2686
0 2688 5 1 1 2687
0 2689 7 1 2 2684 2688
0 2690 5 1 1 2689
0 2691 7 1 2 30911 2690
0 2692 5 1 1 2691
0 2693 7 1 2 22693 26903
0 2694 5 1 1 2693
0 2695 7 1 2 251 2694
0 2696 5 12 1 2695
0 2697 7 1 2 30933 29983
0 2698 5 1 1 2697
0 2699 7 3 2 27603 29822
0 2700 5 1 1 30945
0 2701 7 7 2 24838 23383
0 2702 5 1 1 30948
0 2703 7 1 2 22694 30949
0 2704 7 1 2 30946 2703
0 2705 5 1 1 2704
0 2706 7 1 2 2698 2705
0 2707 5 2 1 2706
0 2708 7 1 2 28112 30955
0 2709 5 1 1 2708
0 2710 7 5 2 24071 26904
0 2711 7 2 2 24169 30957
0 2712 7 1 2 25479 30123
0 2713 7 2 2 30962 2712
0 2714 5 1 1 30964
0 2715 7 1 2 24839 30965
0 2716 5 1 1 2715
0 2717 7 1 2 2709 2716
0 2718 5 2 1 2717
0 2719 7 1 2 25861 30966
0 2720 5 1 1 2719
0 2721 7 2 2 26046 30912
0 2722 7 1 2 23520 30188
0 2723 7 1 2 26861 2722
0 2724 5 1 1 2723
0 2725 7 1 2 27067 29385
0 2726 5 1 1 2725
0 2727 7 1 2 2724 2726
0 2728 5 1 1 2727
0 2729 7 1 2 30968 2728
0 2730 5 1 1 2729
0 2731 7 1 2 2720 2730
0 2732 5 1 1 2731
0 2733 7 1 2 28530 2732
0 2734 5 1 1 2733
0 2735 7 18 2 22695 23384
0 2736 5 2 1 30970
0 2737 7 8 2 25952 30971
0 2738 7 1 2 29969 30990
0 2739 5 1 1 2738
0 2740 7 1 2 26047 29859
0 2741 7 1 2 30934 2740
0 2742 5 1 1 2741
0 2743 7 1 2 2739 2742
0 2744 5 1 1 2743
0 2745 7 1 2 28113 2744
0 2746 5 1 1 2745
0 2747 7 1 2 2714 2746
0 2748 5 1 1 2747
0 2749 7 1 2 30419 2748
0 2750 5 1 1 2749
0 2751 7 1 2 29823 29998
0 2752 5 1 1 2751
0 2753 7 1 2 30972 30398
0 2754 7 1 2 2752 2753
0 2755 5 1 1 2754
0 2756 7 4 2 30327 28501
0 2757 5 2 1 30998
0 2758 7 1 2 30988 31002
0 2759 5 1 1 2758
0 2760 7 18 2 24656 25340
0 2761 5 2 1 31004
0 2762 7 1 2 28114 31022
0 2763 7 1 2 2759 2762
0 2764 7 1 2 2755 2763
0 2765 5 1 1 2764
0 2766 7 2 2 23325 26905
0 2767 7 14 2 22555 24657
0 2768 7 2 2 24072 31026
0 2769 7 1 2 31024 31040
0 2770 7 1 2 29999 2769
0 2771 5 1 1 2770
0 2772 7 1 2 2765 2771
0 2773 5 1 1 2772
0 2774 7 1 2 29029 2773
0 2775 5 1 1 2774
0 2776 7 1 2 2750 2775
0 2777 5 1 1 2776
0 2778 7 1 2 25862 2777
0 2779 5 1 1 2778
0 2780 7 1 2 2734 2779
0 2781 7 1 2 2692 2780
0 2782 5 1 1 2781
0 2783 7 1 2 26228 2782
0 2784 5 1 1 2783
0 2785 7 2 2 23086 26468
0 2786 7 1 2 31042 28532
0 2787 5 1 1 2786
0 2788 7 1 2 29068 2787
0 2789 5 1 1 2788
0 2790 7 1 2 26636 2789
0 2791 5 1 1 2790
0 2792 7 1 2 29098 30424
0 2793 5 1 1 2792
0 2794 7 1 2 2791 2793
0 2795 5 1 1 2794
0 2796 7 1 2 26906 2795
0 2797 5 1 1 2796
0 2798 7 4 2 23017 25341
0 2799 7 2 2 31044 26408
0 2800 7 5 2 25953 24251
0 2801 7 5 2 25035 23521
0 2802 7 1 2 31050 31055
0 2803 7 1 2 31048 2802
0 2804 5 1 1 2803
0 2805 7 1 2 2797 2804
0 2806 5 1 1 2805
0 2807 7 1 2 26137 2806
0 2808 5 1 1 2807
0 2809 7 1 2 26768 30666
0 2810 5 1 1 2809
0 2811 7 1 2 793 2810
0 2812 5 1 1 2811
0 2813 7 1 2 23018 2812
0 2814 5 1 1 2813
0 2815 7 3 2 26138 26590
0 2816 5 2 1 31060
0 2817 7 4 2 23987 26305
0 2818 7 3 2 23385 23617
0 2819 7 1 2 31065 31069
0 2820 7 1 2 31063 2819
0 2821 5 1 1 2820
0 2822 7 1 2 2814 2821
0 2823 5 1 1 2822
0 2824 7 1 2 23087 2823
0 2825 5 1 1 2824
0 2826 7 1 2 30189 31049
0 2827 5 1 1 2826
0 2828 7 1 2 2825 2827
0 2829 5 1 1 2828
0 2830 7 1 2 29052 2829
0 2831 5 1 1 2830
0 2832 7 1 2 2808 2831
0 2833 5 1 1 2832
0 2834 7 1 2 2833 30969
0 2835 5 1 1 2834
0 2836 7 1 2 30425 30967
0 2837 5 1 1 2836
0 2838 7 1 2 29198 30496
0 2839 5 1 1 2838
0 2840 7 6 2 24170 24326
0 2841 7 1 2 26480 31072
0 2842 5 1 1 2841
0 2843 7 2 2 25036 30000
0 2844 7 1 2 26306 31078
0 2845 5 1 1 2844
0 2846 7 1 2 2842 2845
0 2847 5 1 1 2846
0 2848 7 1 2 23618 2847
0 2849 5 1 1 2848
0 2850 7 1 2 2839 2849
0 2851 5 1 1 2850
0 2852 7 1 2 23019 2851
0 2853 5 1 1 2852
0 2854 7 1 2 29659 26431
0 2855 5 1 1 2854
0 2856 7 2 2 27622 30362
0 2857 7 1 2 31080 29563
0 2858 5 1 1 2857
0 2859 7 1 2 2855 2858
0 2860 7 1 2 2853 2859
0 2861 5 1 1 2860
0 2862 7 1 2 952 2016
0 2863 5 2 1 2862
0 2864 7 1 2 22556 31082
0 2865 5 1 1 2864
0 2866 7 1 2 965 2865
0 2867 5 1 1 2866
0 2868 7 1 2 23386 2867
0 2869 5 1 1 2868
0 2870 7 5 2 22557 31005
0 2871 5 1 1 31084
0 2872 7 6 2 23326 25954
0 2873 7 1 2 31085 31089
0 2874 5 1 1 2873
0 2875 7 1 2 2869 2874
0 2876 5 1 1 2875
0 2877 7 1 2 24073 2876
0 2878 7 1 2 2861 2877
0 2879 5 1 1 2878
0 2880 7 1 2 28502 29074
0 2881 5 1 1 2880
0 2882 7 1 2 29995 29046
0 2883 5 1 1 2882
0 2884 7 1 2 2881 2883
0 2885 5 1 1 2884
0 2886 7 1 2 23020 2885
0 2887 5 1 1 2886
0 2888 7 3 2 26139 26432
0 2889 5 1 1 31095
0 2890 7 1 2 29053 31096
0 2891 5 1 1 2890
0 2892 7 1 2 2887 2891
0 2893 5 1 1 2892
0 2894 7 2 2 28115 30935
0 2895 5 1 1 31098
0 2896 7 1 2 26048 31099
0 2897 7 1 2 2893 2896
0 2898 5 1 1 2897
0 2899 7 1 2 2879 2898
0 2900 5 1 1 2899
0 2901 7 1 2 24252 2900
0 2902 5 1 1 2901
0 2903 7 1 2 2837 2902
0 2904 5 1 1 2903
0 2905 7 1 2 25863 2904
0 2906 5 1 1 2905
0 2907 7 1 2 2835 2906
0 2908 7 1 2 2784 2907
0 2909 5 1 1 2908
0 2910 7 1 2 29412 2909
0 2911 5 1 1 2910
0 2912 7 1 2 2644 2911
0 2913 5 1 1 2912
0 2914 7 1 2 22393 2913
0 2915 5 1 1 2914
0 2916 7 8 2 24406 25664
0 2917 7 22 2 23888 23988
0 2918 7 6 2 23231 25342
0 2919 7 1 2 31108 31130
0 2920 5 1 1 2919
0 2921 7 2 2 25180 25955
0 2922 7 4 2 27152 31136
0 2923 5 1 1 31138
0 2924 7 1 2 2920 2923
0 2925 5 5 1 2924
0 2926 7 1 2 28116 29555
0 2927 7 1 2 30884 2926
0 2928 5 1 1 2927
0 2929 7 1 2 28117 26818
0 2930 7 1 2 29991 2929
0 2931 5 1 1 2930
0 2932 7 1 2 2928 2931
0 2933 5 1 1 2932
0 2934 7 1 2 31142 2933
0 2935 5 1 1 2934
0 2936 7 2 2 23232 30430
0 2937 5 3 1 31147
0 2938 7 3 2 25181 27430
0 2939 5 1 1 31152
0 2940 7 1 2 31149 2939
0 2941 5 12 1 2940
0 2942 7 1 2 31027 30875
0 2943 5 1 1 2942
0 2944 7 1 2 2077 2943
0 2945 5 1 1 2944
0 2946 7 1 2 31155 2945
0 2947 5 1 1 2946
0 2948 7 4 2 25182 27841
0 2949 5 1 1 31167
0 2950 7 1 2 31168 29984
0 2951 5 1 1 2950
0 2952 7 7 2 24074 29316
0 2953 7 1 2 30636 30377
0 2954 7 1 2 31171 2953
0 2955 5 1 1 2954
0 2956 7 1 2 2951 2955
0 2957 5 1 1 2956
0 2958 7 1 2 27301 2957
0 2959 5 1 1 2958
0 2960 7 1 2 2947 2959
0 2961 5 1 1 2960
0 2962 7 1 2 26819 2961
0 2963 5 1 1 2962
0 2964 7 2 2 24544 30616
0 2965 7 1 2 29970 31178
0 2966 5 1 1 2965
0 2967 7 1 2 31169 30677
0 2968 5 1 1 2967
0 2969 7 1 2 2966 2968
0 2970 5 1 1 2969
0 2971 7 1 2 22916 2970
0 2972 5 1 1 2971
0 2973 7 3 2 24075 26796
0 2974 7 17 2 24545 24658
0 2975 7 5 2 24840 23233
0 2976 7 3 2 31183 31200
0 2977 7 1 2 31180 31205
0 2978 5 1 1 2977
0 2979 7 1 2 2972 2978
0 2980 5 1 1 2979
0 2981 7 1 2 27302 2980
0 2982 5 1 1 2981
0 2983 7 1 2 27604 31041
0 2984 5 1 1 2983
0 2985 7 1 2 27452 30678
0 2986 5 1 1 2985
0 2987 7 1 2 2984 2986
0 2988 5 1 1 2987
0 2989 7 1 2 22917 2988
0 2990 5 1 1 2989
0 2991 7 3 2 24841 31181
0 2992 7 1 2 31208 31028
0 2993 5 1 1 2992
0 2994 7 1 2 2990 2993
0 2995 5 1 1 2994
0 2996 7 1 2 31156 2995
0 2997 5 1 1 2996
0 2998 7 1 2 2982 2997
0 2999 5 1 1 2998
0 3000 7 1 2 29556 2999
0 3001 5 1 1 3000
0 3002 7 1 2 2963 3001
0 3003 5 1 1 3002
0 3004 7 1 2 27068 3003
0 3005 5 1 1 3004
0 3006 7 1 2 2935 3005
0 3007 5 1 1 3006
0 3008 7 1 2 31100 3007
0 3009 5 1 1 3008
0 3010 7 1 2 23763 3009
0 3011 7 1 2 2915 3010
0 3012 5 1 1 3011
0 3013 7 1 2 2575 3012
0 3014 5 1 1 3013
0 3015 7 1 2 1420 3014
0 3016 5 1 1 3015
0 3017 7 1 2 28970 3016
0 3018 5 1 1 3017
0 3019 7 12 2 22918 24076
0 3020 7 1 2 31211 26820
0 3021 5 2 1 3020
0 3022 7 7 2 24842 26049
0 3023 7 9 2 25611 29615
0 3024 7 1 2 31225 31232
0 3025 5 1 1 3024
0 3026 7 1 2 31223 3025
0 3027 5 1 1 3026
0 3028 7 2 2 30688 30571
0 3029 7 1 2 26885 31241
0 3030 5 1 1 3029
0 3031 7 1 2 27275 27869
0 3032 5 1 1 3031
0 3033 7 1 2 30637 27349
0 3034 5 1 1 3033
0 3035 7 1 2 3032 3034
0 3036 5 2 1 3035
0 3037 7 1 2 24407 31243
0 3038 5 1 1 3037
0 3039 7 1 2 3030 3038
0 3040 5 1 1 3039
0 3041 7 1 2 27303 3040
0 3042 5 1 1 3041
0 3043 7 1 2 24408 31157
0 3044 5 1 1 3043
0 3045 7 3 2 27917 30431
0 3046 5 2 1 31245
0 3047 7 1 2 3044 31248
0 3048 5 3 1 3047
0 3049 7 1 2 27821 31250
0 3050 5 1 1 3049
0 3051 7 1 2 3042 3050
0 3052 5 1 1 3051
0 3053 7 1 2 23764 3052
0 3054 5 1 1 3053
0 3055 7 3 2 27014 28269
0 3056 5 1 1 31253
0 3057 7 2 2 25408 31254
0 3058 7 3 2 24659 29597
0 3059 7 1 2 27644 31258
0 3060 7 1 2 31256 3059
0 3061 5 1 1 3060
0 3062 7 1 2 3054 3061
0 3063 5 1 1 3062
0 3064 7 1 2 3027 3063
0 3065 5 1 1 3064
0 3066 7 6 2 22558 23765
0 3067 5 2 1 31261
0 3068 7 1 2 25183 27427
0 3069 5 1 1 3068
0 3070 7 3 2 25409 23889
0 3071 7 2 2 25270 31269
0 3072 7 8 2 24728 23234
0 3073 7 2 2 24660 31274
0 3074 7 1 2 31272 31282
0 3075 5 1 1 3074
0 3076 7 1 2 3069 3075
0 3077 5 1 1 3076
0 3078 7 2 2 31262 3077
0 3079 5 2 1 31284
0 3080 7 1 2 23766 27276
0 3081 7 2 2 31158 3080
0 3082 5 2 1 31288
0 3083 7 3 2 27283 28254
0 3084 5 2 1 31292
0 3085 7 1 2 25184 26493
0 3086 5 1 1 3085
0 3087 7 1 2 27015 28283
0 3088 7 1 2 3086 3087
0 3089 5 1 1 3088
0 3090 7 1 2 31295 3089
0 3091 5 1 1 3090
0 3092 7 1 2 27350 3091
0 3093 5 1 1 3092
0 3094 7 1 2 31290 3093
0 3095 5 1 1 3094
0 3096 7 1 2 24546 3095
0 3097 5 1 1 3096
0 3098 7 1 2 31286 3097
0 3099 5 1 1 3098
0 3100 7 1 2 24409 3099
0 3101 5 1 1 3100
0 3102 7 1 2 30432 27277
0 3103 5 1 1 3102
0 3104 7 1 2 327 3103
0 3105 5 1 1 3104
0 3106 7 1 2 24547 3105
0 3107 5 1 1 3106
0 3108 7 4 2 22559 27334
0 3109 7 1 2 31297 31273
0 3110 5 1 1 3109
0 3111 7 1 2 3107 3110
0 3112 5 5 1 3111
0 3113 7 5 2 25185 23767
0 3114 5 2 1 31306
0 3115 7 2 2 22394 31307
0 3116 5 1 1 31313
0 3117 7 1 2 31301 31314
0 3118 5 1 1 3117
0 3119 7 1 2 3101 3118
0 3120 5 1 1 3119
0 3121 7 1 2 30411 3120
0 3122 5 1 1 3121
0 3123 7 11 2 25271 25410
0 3124 5 1 1 31315
0 3125 7 1 2 25612 31316
0 3126 7 2 2 31259 3125
0 3127 7 4 2 23021 25186
0 3128 7 3 2 24729 25739
0 3129 7 1 2 31328 31332
0 3130 7 1 2 28926 3129
0 3131 7 1 2 31326 3130
0 3132 5 1 1 3131
0 3133 7 1 2 3122 3132
0 3134 5 1 1 3133
0 3135 7 1 2 24253 3134
0 3136 5 1 1 3135
0 3137 7 6 2 24947 25740
0 3138 5 1 1 31335
0 3139 7 2 2 24730 31336
0 3140 7 7 2 25187 25864
0 3141 7 1 2 31343 26669
0 3142 7 1 2 31341 3141
0 3143 7 1 2 31327 3142
0 3144 5 1 1 3143
0 3145 7 1 2 3136 3144
0 3146 5 1 1 3145
0 3147 7 1 2 31226 3146
0 3148 5 1 1 3147
0 3149 7 1 2 3065 3148
0 3150 5 1 1 3149
0 3151 7 1 2 27069 3150
0 3152 5 1 1 3151
0 3153 7 2 2 24548 28022
0 3154 5 1 1 31350
0 3155 7 7 2 24731 31029
0 3156 7 1 2 31317 31352
0 3157 5 1 1 3156
0 3158 7 2 2 3154 3157
0 3159 5 5 1 31359
0 3160 7 1 2 31227 29557
0 3161 5 1 1 3160
0 3162 7 1 2 31224 3161
0 3163 5 4 1 3162
0 3164 7 1 2 26368 31366
0 3165 5 1 1 3164
0 3166 7 2 2 26050 29575
0 3167 7 4 2 24843 25343
0 3168 5 1 1 31372
0 3169 7 1 2 25956 31373
0 3170 7 1 2 31370 3169
0 3171 5 1 1 3170
0 3172 7 1 2 3165 3171
0 3173 5 1 1 3172
0 3174 7 1 2 31361 3173
0 3175 5 1 1 3174
0 3176 7 3 2 28180 31367
0 3177 7 1 2 27044 31376
0 3178 5 1 1 3177
0 3179 7 1 2 3175 3178
0 3180 5 1 1 3179
0 3181 7 1 2 23890 3180
0 3182 5 1 1 3181
0 3183 7 2 2 24077 30729
0 3184 7 1 2 26958 27361
0 3185 7 1 2 31379 3184
0 3186 7 1 2 27126 26821
0 3187 7 1 2 3185 3186
0 3188 5 1 1 3187
0 3189 7 1 2 3182 3188
0 3190 5 1 1 3189
0 3191 7 1 2 25741 3190
0 3192 5 1 1 3191
0 3193 7 1 2 27160 31377
0 3194 5 1 1 3193
0 3195 7 1 2 3192 3194
0 3196 5 1 1 3195
0 3197 7 1 2 28937 3196
0 3198 5 1 1 3197
0 3199 7 2 2 23768 29219
0 3200 7 1 2 31368 31381
0 3201 5 1 1 3200
0 3202 7 2 2 25742 30080
0 3203 7 1 2 30572 31383
0 3204 7 1 2 31371 3203
0 3205 5 1 1 3204
0 3206 7 1 2 3201 3205
0 3207 5 1 1 3206
0 3208 7 1 2 24410 3207
0 3209 5 1 1 3208
0 3210 7 5 2 25188 28051
0 3211 7 1 2 25272 23769
0 3212 7 3 2 31385 3211
0 3213 5 1 1 31390
0 3214 7 1 2 31369 31391
0 3215 5 1 1 3214
0 3216 7 1 2 3209 3215
0 3217 5 1 1 3216
0 3218 7 1 2 27731 3217
0 3219 5 1 1 3218
0 3220 7 6 2 23770 23989
0 3221 7 2 2 27173 31393
0 3222 7 1 2 27945 31399
0 3223 7 1 2 31378 3222
0 3224 5 1 1 3223
0 3225 7 1 2 3219 3224
0 3226 7 1 2 3198 3225
0 3227 7 1 2 3152 3226
0 3228 5 1 1 3227
0 3229 7 1 2 26797 3228
0 3230 5 1 1 3229
0 3231 7 1 2 22696 28720
0 3232 5 1 1 3231
0 3233 7 1 2 24661 28812
0 3234 5 1 1 3233
0 3235 7 2 2 3232 3234
0 3236 5 8 1 31401
0 3237 7 1 2 25273 31403
0 3238 5 1 1 3237
0 3239 7 2 2 28795 27335
0 3240 5 1 1 31411
0 3241 7 1 2 3238 3240
0 3242 5 4 1 3241
0 3243 7 2 2 24549 31413
0 3244 5 1 1 31417
0 3245 7 12 2 22560 24732
0 3246 7 3 2 31419 28783
0 3247 5 1 1 31431
0 3248 7 1 2 31432 28015
0 3249 5 1 1 3248
0 3250 7 1 2 3244 3249
0 3251 5 2 1 3250
0 3252 7 1 2 23088 26781
0 3253 5 1 1 3252
0 3254 7 1 2 26728 3253
0 3255 5 2 1 3254
0 3256 7 7 2 23022 26643
0 3257 5 1 1 31438
0 3258 7 1 2 31436 31439
0 3259 5 1 1 3258
0 3260 7 1 2 28637 28579
0 3261 7 1 2 26712 3260
0 3262 5 1 1 3261
0 3263 7 1 2 3259 3262
0 3264 5 1 1 3263
0 3265 7 5 2 24078 26964
0 3266 7 16 2 24411 25743
0 3267 5 1 1 31450
0 3268 7 1 2 27368 31451
0 3269 7 1 2 31445 3268
0 3270 7 1 2 3264 3269
0 3271 7 1 2 31434 3270
0 3272 5 1 1 3271
0 3273 7 1 2 3230 3272
0 3274 5 1 1 3273
0 3275 7 1 2 25665 3274
0 3276 5 1 1 3275
0 3277 7 1 2 27557 425
0 3278 5 23 1 3277
0 3279 7 1 2 29358 30519
0 3280 5 2 1 3279
0 3281 7 2 2 23669 31489
0 3282 7 6 2 22561 27267
0 3283 7 1 2 25274 23447
0 3284 7 1 2 27231 3283
0 3285 7 1 2 31493 3284
0 3286 5 2 1 3285
0 3287 7 1 2 27837 31499
0 3288 5 1 1 3287
0 3289 7 1 2 23235 3288
0 3290 5 1 1 3289
0 3291 7 1 2 27880 3290
0 3292 5 2 1 3291
0 3293 7 1 2 31491 31501
0 3294 5 1 1 3293
0 3295 7 14 2 25666 23771
0 3296 7 5 2 25189 31503
0 3297 5 2 1 31517
0 3298 7 3 2 29297 30517
0 3299 5 1 1 31524
0 3300 7 1 2 31518 31525
0 3301 7 1 2 31302 3300
0 3302 5 1 1 3301
0 3303 7 1 2 22395 3302
0 3304 7 1 2 3294 3303
0 3305 5 1 1 3304
0 3306 7 1 2 27304 31244
0 3307 5 1 1 3306
0 3308 7 1 2 31159 27822
0 3309 5 1 1 3308
0 3310 7 1 2 3307 3309
0 3311 5 2 1 3310
0 3312 7 2 2 23772 31527
0 3313 5 1 1 31529
0 3314 7 1 2 29473 31530
0 3315 5 1 1 3314
0 3316 7 1 2 27198 30607
0 3317 7 1 2 27856 3316
0 3318 5 1 1 3317
0 3319 7 1 2 3315 3318
0 3320 5 1 1 3319
0 3321 7 1 2 26433 3320
0 3322 5 1 1 3321
0 3323 7 2 2 31184 27645
0 3324 7 1 2 31531 31257
0 3325 5 1 1 3324
0 3326 7 1 2 3313 3325
0 3327 5 1 1 3326
0 3328 7 1 2 29503 3327
0 3329 5 1 1 3328
0 3330 7 1 2 3322 3329
0 3331 5 1 1 3330
0 3332 7 1 2 26561 3331
0 3333 5 1 1 3332
0 3334 7 1 2 31494 26670
0 3335 7 3 2 25613 27199
0 3336 7 2 2 23448 26529
0 3337 7 1 2 30608 31536
0 3338 7 1 2 31533 3337
0 3339 7 1 2 3334 3338
0 3340 5 1 1 3339
0 3341 7 1 2 24412 3340
0 3342 7 1 2 3333 3341
0 3343 5 1 1 3342
0 3344 7 1 2 3305 3343
0 3345 5 1 1 3344
0 3346 7 3 2 23089 23670
0 3347 7 3 2 27576 31538
0 3348 7 1 2 22396 31502
0 3349 5 1 1 3348
0 3350 7 1 2 27903 3349
0 3351 5 1 1 3350
0 3352 7 1 2 31541 3351
0 3353 5 1 1 3352
0 3354 7 2 2 25037 28698
0 3355 7 1 2 24413 31544
0 3356 7 5 2 24733 31185
0 3357 7 2 2 24254 30549
0 3358 7 5 2 25190 31318
0 3359 7 1 2 31551 31553
0 3360 7 1 2 31546 3359
0 3361 7 1 2 3355 3360
0 3362 5 1 1 3361
0 3363 7 1 2 3353 3362
0 3364 5 1 1 3363
0 3365 7 1 2 27478 3364
0 3366 5 1 1 3365
0 3367 7 2 2 27882 27894
0 3368 7 5 2 22786 23671
0 3369 7 1 2 27742 31560
0 3370 7 2 2 31558 3369
0 3371 7 1 2 29075 31565
0 3372 5 1 1 3371
0 3373 7 4 2 31319 27826
0 3374 7 2 2 27369 30088
0 3375 7 3 2 25614 25865
0 3376 7 1 2 31571 31573
0 3377 7 1 2 31567 3376
0 3378 5 1 1 3377
0 3379 7 1 2 3372 3378
0 3380 5 1 1 3379
0 3381 7 1 2 31452 3380
0 3382 5 1 1 3381
0 3383 7 2 2 28255 30107
0 3384 7 1 2 28043 31576
0 3385 5 1 1 3384
0 3386 7 4 2 22697 29207
0 3387 7 1 2 26335 31578
0 3388 5 1 1 3387
0 3389 7 1 2 28070 27351
0 3390 5 1 1 3389
0 3391 7 1 2 3388 3390
0 3392 5 4 1 3391
0 3393 7 1 2 22562 31582
0 3394 5 1 1 3393
0 3395 7 1 2 30638 28023
0 3396 5 1 1 3395
0 3397 7 1 2 3394 3396
0 3398 5 3 1 3397
0 3399 7 3 2 23672 27200
0 3400 7 1 2 31586 31589
0 3401 5 1 1 3400
0 3402 7 1 2 3385 3401
0 3403 5 1 1 3402
0 3404 7 1 2 22397 29076
0 3405 7 1 2 3403 3404
0 3406 5 1 1 3405
0 3407 7 1 2 3382 3406
0 3408 5 1 1 3407
0 3409 7 1 2 27577 3408
0 3410 5 1 1 3409
0 3411 7 4 2 26809 29909
0 3412 5 3 1 31592
0 3413 7 13 2 23673 25744
0 3414 7 4 2 23236 31599
0 3415 5 3 1 31612
0 3416 7 1 2 31522 31616
0 3417 5 6 1 3416
0 3418 7 3 2 22398 25866
0 3419 5 1 1 31625
0 3420 7 10 2 22563 23891
0 3421 5 4 1 31628
0 3422 7 1 2 31638 1388
0 3423 7 1 2 3419 3422
0 3424 7 1 2 31619 3423
0 3425 5 1 1 3424
0 3426 7 2 2 22564 30108
0 3427 7 2 2 22399 28284
0 3428 5 1 1 31644
0 3429 7 1 2 31642 31645
0 3430 5 1 1 3429
0 3431 7 6 2 25667 28435
0 3432 7 1 2 24414 30639
0 3433 7 1 2 31646 3432
0 3434 5 1 1 3433
0 3435 7 1 2 3430 3434
0 3436 7 1 2 3425 3435
0 3437 5 1 1 3436
0 3438 7 1 2 28024 3437
0 3439 5 1 1 3438
0 3440 7 15 2 24550 25867
0 3441 5 1 1 31652
0 3442 7 1 2 3441 31639
0 3443 5 25 1 3442
0 3444 7 3 2 22787 23237
0 3445 7 2 2 28030 31692
0 3446 7 4 2 22698 23773
0 3447 7 1 2 31697 29634
0 3448 7 1 2 31695 3447
0 3449 5 1 1 3448
0 3450 7 7 2 24734 25275
0 3451 7 2 2 27717 31701
0 3452 7 5 2 24415 24662
0 3453 7 8 2 25668 25745
0 3454 5 1 1 31715
0 3455 7 2 2 25411 31716
0 3456 7 1 2 31710 31723
0 3457 7 1 2 31708 3456
0 3458 5 1 1 3457
0 3459 7 1 2 3449 3458
0 3460 5 1 1 3459
0 3461 7 1 2 31653 3460
0 3462 5 1 1 3461
0 3463 7 2 2 25412 31702
0 3464 7 2 2 31725 30689
0 3465 5 1 1 31727
0 3466 7 1 2 616 3465
0 3467 5 1 1 3466
0 3468 7 1 2 31620 3467
0 3469 5 1 1 3468
0 3470 7 2 2 23674 27861
0 3471 7 1 2 27918 27278
0 3472 7 1 2 31729 3471
0 3473 5 1 1 3472
0 3474 7 1 2 31711 31504
0 3475 7 1 2 28080 3474
0 3476 5 1 1 3475
0 3477 7 1 2 3473 3476
0 3478 7 1 2 3469 3477
0 3479 7 1 2 3462 3478
0 3480 5 1 1 3479
0 3481 7 1 2 31667 3480
0 3482 5 1 1 3481
0 3483 7 1 2 3439 3482
0 3484 5 1 1 3483
0 3485 7 1 2 31593 3484
0 3486 5 1 1 3485
0 3487 7 1 2 3410 3486
0 3488 7 1 2 3366 3487
0 3489 7 1 2 3345 3488
0 3490 5 1 1 3489
0 3491 7 1 2 27070 3490
0 3492 5 1 1 3491
0 3493 7 3 2 30845 26591
0 3494 7 1 2 31285 31731
0 3495 5 1 1 3494
0 3496 7 1 2 27352 31293
0 3497 5 1 1 3496
0 3498 7 1 2 31291 3497
0 3499 5 1 1 3498
0 3500 7 1 2 31732 3499
0 3501 5 1 1 3500
0 3502 7 3 2 25746 26733
0 3503 5 1 1 31734
0 3504 7 1 2 25191 3503
0 3505 5 1 1 3504
0 3506 7 4 2 23090 23774
0 3507 7 5 2 26592 31737
0 3508 5 1 1 31741
0 3509 7 1 2 23238 3508
0 3510 5 1 1 3509
0 3511 7 3 2 3505 3510
0 3512 7 1 2 24844 31746
0 3513 5 1 1 3512
0 3514 7 4 2 22919 26569
0 3515 5 2 1 31749
0 3516 7 2 2 25747 31750
0 3517 7 1 2 25192 31755
0 3518 5 1 1 3517
0 3519 7 1 2 3513 3518
0 3520 5 1 1 3519
0 3521 7 1 2 27016 27353
0 3522 7 1 2 3520 3521
0 3523 5 1 1 3522
0 3524 7 1 2 3501 3523
0 3525 5 1 1 3524
0 3526 7 1 2 24551 3525
0 3527 5 1 1 3526
0 3528 7 1 2 3495 3527
0 3529 5 1 1 3528
0 3530 7 1 2 24416 3529
0 3531 5 1 1 3530
0 3532 7 2 2 26593 31303
0 3533 7 3 2 25193 29918
0 3534 7 1 2 31738 31759
0 3535 7 1 2 31757 3534
0 3536 5 1 1 3535
0 3537 7 1 2 3531 3536
0 3538 5 1 1 3537
0 3539 7 1 2 27071 3538
0 3540 5 1 1 3539
0 3541 7 3 2 29246 31742
0 3542 5 1 1 31762
0 3543 7 4 2 29598 29584
0 3544 7 1 2 31765 31735
0 3545 5 1 1 3544
0 3546 7 1 2 3542 3545
0 3547 5 1 1 3546
0 3548 7 1 2 24845 3547
0 3549 5 1 1 3548
0 3550 7 1 2 31766 31756
0 3551 5 1 1 3550
0 3552 7 1 2 3549 3551
0 3553 5 1 1 3552
0 3554 7 1 2 27732 3553
0 3555 5 1 1 3554
0 3556 7 1 2 25194 27186
0 3557 5 1 1 3556
0 3558 7 4 2 23990 27174
0 3559 7 1 2 28256 31769
0 3560 5 1 1 3559
0 3561 7 1 2 3557 3560
0 3562 5 1 1 3561
0 3563 7 3 2 26594 28181
0 3564 7 1 2 30846 31773
0 3565 7 1 2 3562 3564
0 3566 5 1 1 3565
0 3567 7 3 2 24846 26734
0 3568 5 5 1 31776
0 3569 7 1 2 31779 31753
0 3570 5 2 1 3569
0 3571 7 1 2 26769 31784
0 3572 5 1 1 3571
0 3573 7 1 2 26369 31733
0 3574 5 1 1 3573
0 3575 7 1 2 3572 3574
0 3576 5 1 1 3575
0 3577 7 1 2 23892 28270
0 3578 7 1 2 31362 3577
0 3579 7 1 2 3576 3578
0 3580 5 1 1 3579
0 3581 7 1 2 3566 3580
0 3582 5 1 1 3581
0 3583 7 1 2 24417 3582
0 3584 5 1 1 3583
0 3585 7 3 2 31774 31400
0 3586 7 1 2 27718 29919
0 3587 7 1 2 31786 3586
0 3588 5 1 1 3587
0 3589 7 1 2 3584 3588
0 3590 7 1 2 3555 3589
0 3591 7 1 2 3540 3590
0 3592 5 1 1 3591
0 3593 7 1 2 25669 3592
0 3594 5 1 1 3593
0 3595 7 5 2 31006 26886
0 3596 5 1 1 31789
0 3597 7 1 2 29148 31790
0 3598 5 1 1 3597
0 3599 7 2 2 28118 31404
0 3600 5 1 1 31794
0 3601 7 1 2 27946 31795
0 3602 5 1 1 3601
0 3603 7 1 2 3598 3602
0 3604 5 1 1 3603
0 3605 7 6 2 25957 28699
0 3606 7 1 2 26595 31796
0 3607 7 2 2 3604 3606
0 3608 7 1 2 24847 31539
0 3609 7 1 2 31802 3608
0 3610 5 1 1 3609
0 3611 7 1 2 3594 3610
0 3612 5 1 1 3611
0 3613 7 1 2 26505 3612
0 3614 5 1 1 3613
0 3615 7 2 2 29599 30039
0 3616 7 1 2 31804 31572
0 3617 5 1 1 3616
0 3618 7 2 2 23675 29077
0 3619 7 1 2 29149 31806
0 3620 5 1 1 3619
0 3621 7 1 2 3617 3620
0 3622 5 1 1 3621
0 3623 7 1 2 25748 3622
0 3624 5 1 1 3623
0 3625 7 5 2 23775 29371
0 3626 7 1 2 23327 26307
0 3627 7 1 2 31808 3626
0 3628 7 1 2 30536 3627
0 3629 5 1 1 3628
0 3630 7 1 2 3624 3629
0 3631 5 1 1 3630
0 3632 7 1 2 27578 3631
0 3633 5 1 1 3632
0 3634 7 1 2 28374 31542
0 3635 5 1 1 3634
0 3636 7 2 2 29600 30581
0 3637 7 3 2 25749 24255
0 3638 7 1 2 31815 30801
0 3639 7 1 2 31813 3638
0 3640 5 1 1 3639
0 3641 7 1 2 3635 3640
0 3642 5 1 1 3641
0 3643 7 1 2 27479 3642
0 3644 5 1 1 3643
0 3645 7 3 2 23776 29247
0 3646 7 1 2 29782 31818
0 3647 5 1 1 3646
0 3648 7 3 2 23091 28271
0 3649 5 1 1 31821
0 3650 7 1 2 24327 31822
0 3651 7 1 2 31805 3650
0 3652 5 1 1 3651
0 3653 7 1 2 3647 3652
0 3654 5 1 1 3653
0 3655 7 1 2 31552 3654
0 3656 5 1 1 3655
0 3657 7 1 2 28375 31492
0 3658 5 1 1 3657
0 3659 7 1 2 23676 28333
0 3660 5 1 1 3659
0 3661 7 1 2 28302 31519
0 3662 5 1 1 3661
0 3663 7 1 2 22400 3662
0 3664 7 1 2 3660 3663
0 3665 5 1 1 3664
0 3666 7 1 2 28229 31621
0 3667 5 1 1 3666
0 3668 7 1 2 28266 3649
0 3669 5 4 1 3668
0 3670 7 1 2 31824 29449
0 3671 5 1 1 3670
0 3672 7 1 2 24418 3671
0 3673 7 1 2 3667 3672
0 3674 5 1 1 3673
0 3675 7 1 2 3674 31594
0 3676 7 1 2 3665 3675
0 3677 5 1 1 3676
0 3678 7 1 2 3658 3677
0 3679 7 1 2 3656 3678
0 3680 7 1 2 3644 3679
0 3681 7 1 2 3633 3680
0 3682 5 1 1 3681
0 3683 7 1 2 27733 3682
0 3684 5 1 1 3683
0 3685 7 4 2 23991 28802
0 3686 7 5 2 23239 27431
0 3687 7 1 2 31828 31832
0 3688 7 1 2 27770 3687
0 3689 7 1 2 31807 3688
0 3690 5 1 1 3689
0 3691 7 6 2 25958 24328
0 3692 7 7 2 25615 25670
0 3693 7 1 2 31270 31843
0 3694 7 1 2 31837 3693
0 3695 7 11 2 25195 25344
0 3696 5 1 1 31850
0 3697 7 2 2 31851 30402
0 3698 7 1 2 31298 31861
0 3699 7 1 2 3694 3698
0 3700 5 1 1 3699
0 3701 7 1 2 3690 3700
0 3702 5 1 1 3701
0 3703 7 1 2 24419 3702
0 3704 5 1 1 3703
0 3705 7 1 2 27175 28182
0 3706 5 1 1 3705
0 3707 7 1 2 27153 31568
0 3708 5 1 1 3707
0 3709 7 1 2 3706 3708
0 3710 5 1 1 3709
0 3711 7 1 2 23240 3710
0 3712 5 1 1 3711
0 3713 7 5 2 27453 27382
0 3714 5 1 1 31863
0 3715 7 2 2 23449 25868
0 3716 7 4 2 22788 25196
0 3717 7 2 2 31868 31870
0 3718 7 1 2 31864 31874
0 3719 5 1 1 3718
0 3720 7 1 2 3712 3719
0 3721 5 1 1 3720
0 3722 7 2 2 22401 3721
0 3723 5 1 1 31876
0 3724 7 2 2 31066 30526
0 3725 7 1 2 25038 31878
0 3726 7 1 2 31877 3725
0 3727 5 1 1 3726
0 3728 7 1 2 3704 3727
0 3729 5 1 1 3728
0 3730 7 1 2 27579 3729
0 3731 5 1 1 3730
0 3732 7 6 2 25039 23387
0 3733 7 2 2 25959 31880
0 3734 7 2 2 30198 31886
0 3735 5 1 1 31888
0 3736 7 5 2 25345 31109
0 3737 7 1 2 28194 31890
0 3738 5 1 1 3737
0 3739 7 1 2 3735 3738
0 3740 5 1 1 3739
0 3741 7 1 2 23677 3740
0 3742 5 1 1 3741
0 3743 7 4 2 24420 29458
0 3744 7 1 2 25671 31895
0 3745 7 1 2 31770 3744
0 3746 5 1 1 3745
0 3747 7 1 2 3742 3746
0 3748 5 1 1 3747
0 3749 7 1 2 26434 3748
0 3750 5 1 1 3749
0 3751 7 2 2 29396 31891
0 3752 5 1 1 31899
0 3753 7 1 2 29772 28397
0 3754 5 1 1 3753
0 3755 7 1 2 3752 3754
0 3756 5 1 1 3755
0 3757 7 1 2 24421 3756
0 3758 5 1 1 3757
0 3759 7 1 2 31139 29635
0 3760 5 1 1 3759
0 3761 7 1 2 3758 3760
0 3762 5 1 1 3761
0 3763 7 1 2 26494 3762
0 3764 5 1 1 3763
0 3765 7 1 2 3750 3764
0 3766 5 1 1 3765
0 3767 7 1 2 26562 3766
0 3768 5 1 1 3767
0 3769 7 2 2 23023 23893
0 3770 7 1 2 27045 31901
0 3771 7 1 2 29670 3770
0 3772 7 1 2 28475 3771
0 3773 5 1 1 3772
0 3774 7 1 2 3768 3773
0 3775 5 1 1 3774
0 3776 7 1 2 28183 3775
0 3777 5 1 1 3776
0 3778 7 1 2 22402 31143
0 3779 5 1 1 3778
0 3780 7 7 2 24422 25869
0 3781 7 2 2 28398 31903
0 3782 7 1 2 25960 31910
0 3783 5 1 1 3782
0 3784 7 1 2 3779 3783
0 3785 5 1 1 3784
0 3786 7 1 2 23678 3785
0 3787 5 1 1 3786
0 3788 7 1 2 29697 31892
0 3789 5 1 1 3788
0 3790 7 1 2 3787 3789
0 3791 5 1 1 3790
0 3792 7 1 2 28184 3791
0 3793 5 1 1 3792
0 3794 7 2 2 23092 26770
0 3795 5 1 1 31912
0 3796 7 1 2 26383 3795
0 3797 5 2 1 3796
0 3798 7 4 2 24423 24735
0 3799 7 3 2 31030 31916
0 3800 7 1 2 30129 31920
0 3801 7 1 2 31554 3800
0 3802 7 1 2 31914 3801
0 3803 5 1 1 3802
0 3804 7 1 2 3793 3803
0 3805 5 1 1 3804
0 3806 7 1 2 31595 3805
0 3807 5 1 1 3806
0 3808 7 1 2 26370 31490
0 3809 5 1 1 3808
0 3810 7 1 2 26771 26563
0 3811 7 1 2 29783 3810
0 3812 5 1 1 3811
0 3813 7 1 2 3809 3812
0 3814 5 2 1 3813
0 3815 7 1 2 22403 31583
0 3816 5 1 1 3815
0 3817 7 1 2 23241 27891
0 3818 5 1 1 3817
0 3819 7 1 2 3816 3818
0 3820 5 2 1 3819
0 3821 7 4 2 23679 31654
0 3822 7 1 2 31925 31927
0 3823 7 1 2 31923 3822
0 3824 5 1 1 3823
0 3825 7 2 2 25616 27561
0 3826 7 1 2 31838 31931
0 3827 5 1 1 3826
0 3828 7 1 2 26371 29784
0 3829 5 1 1 3828
0 3830 7 1 2 3827 3829
0 3831 5 1 1 3830
0 3832 7 3 2 24256 30130
0 3833 7 1 2 31320 27370
0 3834 7 1 2 31933 3833
0 3835 7 1 2 31921 3834
0 3836 7 1 2 3831 3835
0 3837 5 1 1 3836
0 3838 7 1 2 25750 3837
0 3839 7 1 2 3824 3838
0 3840 7 1 2 3807 3839
0 3841 7 1 2 3777 3840
0 3842 7 1 2 3731 3841
0 3843 7 1 2 31596 3299
0 3844 5 2 1 3843
0 3845 7 1 2 26372 31936
0 3846 5 1 1 3845
0 3847 7 2 2 26495 26564
0 3848 5 1 1 31938
0 3849 7 1 2 31597 3848
0 3850 5 1 1 3849
0 3851 7 1 2 31913 3850
0 3852 5 1 1 3851
0 3853 7 1 2 3846 3852
0 3854 5 1 1 3853
0 3855 7 1 2 30131 30573
0 3856 7 1 2 3854 3855
0 3857 5 1 1 3856
0 3858 7 10 2 22565 25870
0 3859 5 3 1 31940
0 3860 7 3 2 31941 29413
0 3861 5 2 1 31953
0 3862 7 1 2 31954 31924
0 3863 5 1 1 3862
0 3864 7 1 2 26772 31934
0 3865 7 1 2 30586 3864
0 3866 5 1 1 3865
0 3867 7 2 2 26938 27580
0 3868 7 3 2 23093 23388
0 3869 7 2 2 31960 29414
0 3870 7 1 2 22566 31963
0 3871 7 1 2 31958 3870
0 3872 5 1 1 3871
0 3873 7 1 2 3866 3872
0 3874 5 1 1 3873
0 3875 7 1 2 27480 3874
0 3876 5 1 1 3875
0 3877 7 5 2 23242 25871
0 3878 7 6 2 22567 25040
0 3879 7 1 2 23389 31970
0 3880 7 1 2 31965 3879
0 3881 7 1 2 31879 3880
0 3882 5 1 1 3881
0 3883 7 4 2 25672 31852
0 3884 7 4 2 25617 23894
0 3885 7 1 2 27362 31839
0 3886 7 1 2 31980 3885
0 3887 7 1 2 31976 3886
0 3888 5 1 1 3887
0 3889 7 1 2 3882 3888
0 3890 5 1 1 3889
0 3891 7 1 2 27581 3890
0 3892 5 1 1 3891
0 3893 7 1 2 3876 3892
0 3894 7 1 2 3863 3893
0 3895 7 1 2 3857 3894
0 3896 5 1 1 3895
0 3897 7 1 2 24424 3896
0 3898 5 1 1 3897
0 3899 7 2 2 22568 27919
0 3900 7 2 2 30109 31984
0 3901 5 1 1 31986
0 3902 7 1 2 26229 30932
0 3903 5 1 1 3902
0 3904 7 1 2 27489 29084
0 3905 5 1 1 3904
0 3906 7 1 2 30520 3905
0 3907 7 2 2 3903 3906
0 3908 5 1 1 31988
0 3909 7 1 2 26373 3908
0 3910 5 1 1 3909
0 3911 7 1 2 26773 31526
0 3912 5 1 1 3911
0 3913 7 1 2 3910 3912
0 3914 5 1 1 3913
0 3915 7 1 2 31987 3914
0 3916 5 1 1 3915
0 3917 7 1 2 3898 3916
0 3918 5 1 1 3917
0 3919 7 1 2 28025 3918
0 3920 5 1 1 3919
0 3921 7 5 2 25276 28784
0 3922 7 2 2 31420 31990
0 3923 5 1 1 31995
0 3924 7 2 2 24257 30163
0 3925 7 5 2 22920 23895
0 3926 7 1 2 31997 31999
0 3927 7 1 2 29679 3926
0 3928 7 1 2 31996 3927
0 3929 5 1 1 3928
0 3930 7 1 2 28040 31911
0 3931 5 1 1 3930
0 3932 7 1 2 3723 3931
0 3933 5 1 1 3932
0 3934 7 1 2 23992 31543
0 3935 7 1 2 3933 3934
0 3936 5 1 1 3935
0 3937 7 1 2 3929 3936
0 3938 5 1 1 3937
0 3939 7 1 2 27481 3938
0 3940 5 1 1 3939
0 3941 7 1 2 3920 3940
0 3942 7 1 2 3842 3941
0 3943 5 1 1 3942
0 3944 7 2 2 28185 31937
0 3945 7 1 2 31900 32004
0 3946 5 1 1 3945
0 3947 7 1 2 31598 31989
0 3948 5 1 1 3947
0 3949 7 2 2 23390 29752
0 3950 7 1 2 32006 28186
0 3951 5 1 1 3950
0 3952 7 5 2 22569 22789
0 3953 7 2 2 27883 32008
0 3954 7 1 2 28713 26965
0 3955 7 1 2 32013 3954
0 3956 5 1 1 3955
0 3957 7 1 2 3951 3956
0 3958 5 1 1 3957
0 3959 7 1 2 3948 3958
0 3960 5 1 1 3959
0 3961 7 12 2 25041 25618
0 3962 5 1 1 32015
0 3963 7 3 2 22921 32016
0 3964 5 1 1 32027
0 3965 7 1 2 23619 27490
0 3966 5 1 1 3965
0 3967 7 1 2 3964 3966
0 3968 5 1 1 3967
0 3969 7 1 2 24329 3968
0 3970 5 1 1 3969
0 3971 7 1 2 23094 29087
0 3972 5 1 1 3971
0 3973 7 2 2 23024 25619
0 3974 7 1 2 29713 32030
0 3975 5 1 1 3974
0 3976 7 1 2 3975 30234
0 3977 5 1 1 3976
0 3978 7 1 2 24258 3977
0 3979 5 1 1 3978
0 3980 7 1 2 3972 3979
0 3981 7 1 2 3970 3980
0 3982 5 1 1 3981
0 3983 7 7 2 23391 27884
0 3984 7 2 2 22570 31110
0 3985 7 2 2 26336 32039
0 3986 5 1 1 32041
0 3987 7 1 2 32032 32042
0 3988 7 1 2 3982 3987
0 3989 5 1 1 3988
0 3990 7 1 2 3960 3989
0 3991 5 1 1 3990
0 3992 7 1 2 29415 3991
0 3993 5 1 1 3992
0 3994 7 1 2 3946 3993
0 3995 5 1 1 3994
0 3996 7 1 2 22404 3995
0 3997 5 1 1 3996
0 3998 7 1 2 31144 31101
0 3999 7 1 2 32005 3998
0 4000 5 1 1 3999
0 4001 7 1 2 23777 4000
0 4002 7 1 2 3997 4001
0 4003 5 1 1 4002
0 4004 7 1 2 3943 4003
0 4005 5 1 1 4004
0 4006 7 1 2 3684 4005
0 4007 7 1 2 3614 4006
0 4008 7 1 2 3492 4007
0 4009 5 1 1 4008
0 4010 7 1 2 31466 4009
0 4011 5 1 1 4010
0 4012 7 21 2 26 23158
0 4013 5 4 1 32043
0 4014 7 2 2 2544 30858
0 4015 5 59 1 32068
0 4016 7 1 2 32070 29985
0 4017 5 1 1 4016
0 4018 7 2 2 29971 30950
0 4019 5 1 1 32129
0 4020 7 1 2 22699 32130
0 4021 5 1 1 4020
0 4022 7 1 2 4017 4021
0 4023 5 1 1 4022
0 4024 7 1 2 28084 4023
0 4025 5 1 1 4024
0 4026 7 1 2 32071 30873
0 4027 5 1 1 4026
0 4028 7 1 2 23392 29972
0 4029 5 1 1 4028
0 4030 7 3 2 25346 26051
0 4031 5 1 1 32131
0 4032 7 2 2 26140 32132
0 4033 7 1 2 23522 32134
0 4034 5 1 1 4033
0 4035 7 1 2 4029 4034
0 4036 5 2 1 4035
0 4037 7 1 2 22700 32136
0 4038 5 1 1 4037
0 4039 7 1 2 28602 30057
0 4040 5 1 1 4039
0 4041 7 2 2 4038 4040
0 4042 5 1 1 32138
0 4043 7 1 2 25277 32139
0 4044 5 1 1 4043
0 4045 7 2 2 29973 31007
0 4046 5 1 1 32140
0 4047 7 1 2 23328 4046
0 4048 5 1 1 4047
0 4049 7 1 2 24848 4048
0 4050 7 1 2 4044 4049
0 4051 5 1 1 4050
0 4052 7 1 2 4027 4051
0 4053 5 1 1 4052
0 4054 7 1 2 22571 4053
0 4055 5 1 1 4054
0 4056 7 1 2 4025 4055
0 4057 5 1 1 4056
0 4058 7 1 2 26230 4057
0 4059 5 1 1 4058
0 4060 7 7 2 28119 32072
0 4061 7 1 2 32142 30280
0 4062 7 1 2 29850 4061
0 4063 5 1 1 4062
0 4064 7 1 2 4059 4063
0 4065 5 1 1 4064
0 4066 7 1 2 27947 4065
0 4067 5 1 1 4066
0 4068 7 1 2 22405 30477
0 4069 7 4 2 25347 25480
0 4070 7 2 2 25278 32149
0 4071 7 1 2 32153 31206
0 4072 7 1 2 4068 4071
0 4073 5 1 1 4072
0 4074 7 1 2 4067 4073
0 4075 5 1 1 4074
0 4076 7 1 2 23095 31797
0 4077 7 1 2 4075 4076
0 4078 5 1 1 4077
0 4079 7 5 2 23243 27383
0 4080 7 6 2 22922 23025
0 4081 7 3 2 32155 32160
0 4082 7 3 2 23523 23993
0 4083 7 2 2 28436 32169
0 4084 7 1 2 27519 32172
0 4085 7 1 2 28458 4084
0 4086 7 1 2 32166 4085
0 4087 5 1 1 4086
0 4088 7 1 2 23680 4087
0 4089 7 1 2 4078 4088
0 4090 5 1 1 4089
0 4091 7 1 2 27232 30936
0 4092 5 1 1 4091
0 4093 7 3 2 27166 30878
0 4094 5 1 1 32174
0 4095 7 1 2 25348 32175
0 4096 5 1 1 4095
0 4097 7 1 2 4092 4096
0 4098 5 2 1 4097
0 4099 7 1 2 25279 32177
0 4100 5 1 1 4099
0 4101 7 3 2 23896 26907
0 4102 7 2 2 23778 27885
0 4103 7 1 2 32179 32182
0 4104 5 1 1 4103
0 4105 7 1 2 4100 4104
0 4106 5 1 1 4105
0 4107 7 1 2 29986 4106
0 4108 5 1 1 4107
0 4109 7 1 2 22701 27187
0 4110 5 1 1 4109
0 4111 7 13 2 25751 31111
0 4112 7 1 2 32184 30833
0 4113 5 1 1 4112
0 4114 7 1 2 4110 4113
0 4115 5 2 1 4114
0 4116 7 1 2 25280 32197
0 4117 5 1 1 4116
0 4118 7 2 2 26908 28871
0 4119 5 1 1 32199
0 4120 7 1 2 27233 32200
0 4121 5 1 1 4120
0 4122 7 1 2 4117 4121
0 4123 5 1 1 4122
0 4124 7 1 2 4123 30876
0 4125 5 1 1 4124
0 4126 7 1 2 4108 4125
0 4127 5 1 1 4126
0 4128 7 1 2 26596 4127
0 4129 5 1 1 4128
0 4130 7 4 2 25961 29949
0 4131 7 1 2 27201 32201
0 4132 7 3 2 25481 30025
0 4133 7 2 2 23026 28665
0 4134 7 1 2 32205 32208
0 4135 7 1 2 4131 4134
0 4136 5 1 1 4135
0 4137 7 1 2 4129 4136
0 4138 5 1 1 4137
0 4139 7 1 2 23096 4138
0 4140 5 1 1 4139
0 4141 7 5 2 24663 24948
0 4142 7 2 2 24259 27505
0 4143 7 2 2 32210 32215
0 4144 7 5 2 25962 27202
0 4145 7 1 2 28666 26447
0 4146 7 1 2 32219 4145
0 4147 7 1 2 32217 4146
0 4148 5 1 1 4147
0 4149 7 1 2 22572 4148
0 4150 7 1 2 4140 4149
0 4151 5 1 1 4150
0 4152 7 1 2 22702 545
0 4153 5 1 1 4152
0 4154 7 10 2 23329 25349
0 4155 5 1 1 32224
0 4156 7 1 2 24664 4155
0 4157 5 1 1 4156
0 4158 7 26 2 4153 4157
0 4159 7 3 2 30190 30043
0 4160 5 1 1 32260
0 4161 7 1 2 26392 32261
0 4162 5 1 1 4161
0 4163 7 1 2 29866 29099
0 4164 7 1 2 31061 4163
0 4165 5 1 1 4164
0 4166 7 1 2 4162 4165
0 4167 5 1 1 4166
0 4168 7 1 2 32234 4167
0 4169 5 1 1 4168
0 4170 7 2 2 28561 26597
0 4171 7 1 2 32225 32263
0 4172 7 1 2 29536 4171
0 4173 5 1 1 4172
0 4174 7 1 2 4169 4173
0 4175 5 1 1 4174
0 4176 7 1 2 23097 4175
0 4177 5 1 1 4176
0 4178 7 1 2 23330 24079
0 4179 7 1 2 32206 4178
0 4180 5 1 1 4179
0 4181 7 1 2 25281 29795
0 4182 5 1 1 4181
0 4183 7 1 2 4180 4182
0 4184 5 2 1 4183
0 4185 7 1 2 31961 32264
0 4186 5 1 1 4185
0 4187 7 3 2 24949 29179
0 4188 5 2 1 32267
0 4189 7 1 2 26774 32268
0 4190 5 1 1 4189
0 4191 7 1 2 4186 4190
0 4192 5 1 1 4191
0 4193 7 1 2 32265 4192
0 4194 5 1 1 4193
0 4195 7 2 2 26735 29851
0 4196 5 1 1 32272
0 4197 7 1 2 28756 30929
0 4198 7 1 2 32273 4197
0 4199 5 1 1 4198
0 4200 7 1 2 4194 4199
0 4201 7 1 2 4177 4200
0 4202 5 1 1 4201
0 4203 7 1 2 23897 4202
0 4204 5 1 1 4203
0 4205 7 4 2 24665 26909
0 4206 5 1 1 32274
0 4207 7 1 2 29812 26393
0 4208 5 3 1 4207
0 4209 7 2 2 26798 26570
0 4210 5 1 1 32281
0 4211 7 1 2 32278 4210
0 4212 5 2 1 4211
0 4213 7 1 2 24849 32283
0 4214 5 1 1 4213
0 4215 7 6 2 24950 29272
0 4216 7 1 2 26537 32285
0 4217 5 1 1 4216
0 4218 7 1 2 4214 4217
0 4219 5 1 1 4218
0 4220 7 1 2 32275 4219
0 4221 5 1 1 4220
0 4222 7 1 2 29100 26598
0 4223 5 1 1 4222
0 4224 7 1 2 31780 29089
0 4225 5 1 1 4224
0 4226 7 1 2 30854 28562
0 4227 7 1 2 4225 4226
0 4228 7 1 2 4223 4227
0 4229 5 1 1 4228
0 4230 7 1 2 4221 4229
0 4231 5 1 1 4230
0 4232 7 1 2 24080 27017
0 4233 7 1 2 4231 4232
0 4234 5 1 1 4233
0 4235 7 1 2 4204 4234
0 4236 5 1 1 4235
0 4237 7 1 2 25752 4236
0 4238 5 1 1 4237
0 4239 7 1 2 27432 31743
0 4240 7 1 2 30956 4239
0 4241 5 1 1 4240
0 4242 7 1 2 24552 4241
0 4243 7 1 2 4238 4242
0 4244 5 1 1 4243
0 4245 7 1 2 28938 4244
0 4246 7 1 2 4151 4245
0 4247 5 1 1 4246
0 4248 7 1 2 24171 31763
0 4249 5 1 1 4248
0 4250 7 3 2 24951 25197
0 4251 7 2 2 29601 32291
0 4252 7 1 2 27105 29180
0 4253 7 1 2 32294 4252
0 4254 5 1 1 4253
0 4255 7 1 2 4249 4254
0 4256 5 1 1 4255
0 4257 7 1 2 29537 4256
0 4258 5 1 1 4257
0 4259 7 1 2 31747 29386
0 4260 5 1 1 4259
0 4261 7 2 2 22923 31329
0 4262 7 2 2 25753 24172
0 4263 7 1 2 29352 32298
0 4264 7 1 2 32296 4263
0 4265 5 1 1 4264
0 4266 7 1 2 4260 4265
0 4267 5 1 1 4266
0 4268 7 1 2 28303 4267
0 4269 5 1 1 4268
0 4270 7 2 2 26599 29391
0 4271 7 2 2 23098 27870
0 4272 7 1 2 23331 32302
0 4273 7 1 2 32300 4272
0 4274 5 1 1 4273
0 4275 7 1 2 4269 4274
0 4276 5 1 1 4275
0 4277 7 1 2 24425 4276
0 4278 5 1 1 4277
0 4279 7 1 2 30730 31386
0 4280 7 1 2 32301 4279
0 4281 5 1 1 4280
0 4282 7 1 2 4278 4281
0 4283 5 1 1 4282
0 4284 7 1 2 29303 4283
0 4285 5 1 1 4284
0 4286 7 1 2 4258 4285
0 4287 5 1 1 4286
0 4288 7 1 2 26991 4287
0 4289 5 1 1 4288
0 4290 7 1 2 27948 31744
0 4291 7 1 2 30882 4290
0 4292 5 1 1 4291
0 4293 7 1 2 25673 4292
0 4294 7 1 2 4289 4293
0 4295 7 1 2 4247 4294
0 4296 5 1 1 4295
0 4297 7 1 2 28971 4296
0 4298 7 1 2 4090 4297
0 4299 5 1 1 4298
0 4300 7 1 2 765 1180
0 4301 7 2 2 28638 4300
0 4302 7 1 2 29824 31717
0 4303 7 2 2 32304 4302
0 4304 7 7 2 25198 28667
0 4305 7 2 2 29602 32308
0 4306 7 1 2 32161 32315
0 4307 7 1 2 32306 4306
0 4308 5 1 1 4307
0 4309 7 1 2 27520 26394
0 4310 5 1 1 4309
0 4311 7 1 2 26231 27555
0 4312 5 1 1 4311
0 4313 7 1 2 4310 4312
0 4314 5 1 1 4313
0 4315 7 6 2 24850 23994
0 4316 7 15 2 22406 23779
0 4317 5 2 1 32323
0 4318 7 1 2 32324 30454
0 4319 7 1 2 32317 4318
0 4320 7 1 2 32156 4319
0 4321 7 1 2 4314 4320
0 4322 5 1 1 4321
0 4323 7 1 2 4308 4322
0 4324 5 1 1 4323
0 4325 7 1 2 26337 4324
0 4326 5 1 1 4325
0 4327 7 2 2 25282 26838
0 4328 7 7 2 24553 24736
0 4329 7 4 2 24426 32342
0 4330 7 1 2 32340 32349
0 4331 7 1 2 32297 4330
0 4332 7 1 2 32307 4331
0 4333 5 1 1 4332
0 4334 7 1 2 4326 4333
0 4335 5 1 1 4334
0 4336 7 1 2 22703 4335
0 4337 5 1 1 4336
0 4338 7 1 2 24554 28820
0 4339 5 1 1 4338
0 4340 7 1 2 4339 3923
0 4341 5 4 1 4340
0 4342 7 3 2 23027 24081
0 4343 5 1 1 32357
0 4344 7 5 2 22924 25963
0 4345 7 1 2 25754 32360
0 4346 7 1 2 32358 4345
0 4347 7 1 2 29749 4346
0 4348 7 1 2 32305 4347
0 4349 7 1 2 32353 4348
0 4350 5 1 1 4349
0 4351 7 1 2 4337 4350
0 4352 5 1 1 4351
0 4353 7 1 2 23898 4352
0 4354 5 1 1 4353
0 4355 7 1 2 23393 31360
0 4356 5 1 1 4355
0 4357 7 1 2 25350 671
0 4358 5 1 1 4357
0 4359 7 6 2 23099 23899
0 4360 7 1 2 32365 26600
0 4361 7 1 2 4358 4360
0 4362 7 1 2 4356 4361
0 4363 5 1 1 4362
0 4364 7 3 2 27127 31045
0 4365 7 2 2 25872 26232
0 4366 7 1 2 28304 32374
0 4367 7 1 2 32371 4366
0 4368 5 1 1 4367
0 4369 7 1 2 4363 4368
0 4370 5 1 1 4369
0 4371 7 1 2 23995 31212
0 4372 7 1 2 4370 4371
0 4373 5 1 1 4372
0 4374 7 3 2 24851 26571
0 4375 7 5 2 23900 26052
0 4376 7 1 2 26775 32379
0 4377 7 1 2 32376 4376
0 4378 7 1 2 31363 4377
0 4379 5 1 1 4378
0 4380 7 1 2 4373 4379
0 4381 5 1 1 4380
0 4382 7 1 2 25755 4381
0 4383 5 1 1 4382
0 4384 7 3 2 24082 27634
0 4385 7 1 2 27161 32384
0 4386 7 1 2 31775 4385
0 4387 5 1 1 4386
0 4388 7 1 2 4383 4387
0 4389 5 1 1 4388
0 4390 7 1 2 25199 4389
0 4391 5 1 1 4390
0 4392 7 1 2 27669 27467
0 4393 7 1 2 31787 4392
0 4394 5 1 1 4393
0 4395 7 1 2 24555 31289
0 4396 5 1 1 4395
0 4397 7 1 2 31287 4396
0 4398 5 1 1 4397
0 4399 7 1 2 26601 32385
0 4400 7 1 2 4398 4399
0 4401 5 1 1 4400
0 4402 7 1 2 31213 31748
0 4403 5 1 1 4402
0 4404 7 8 2 24852 24952
0 4405 5 1 1 32387
0 4406 7 7 2 26053 24260
0 4407 7 1 2 25756 32395
0 4408 7 2 2 32388 4407
0 4409 7 1 2 25200 32402
0 4410 5 1 1 4409
0 4411 7 1 2 4403 4410
0 4412 5 1 1 4411
0 4413 7 1 2 27018 4412
0 4414 5 1 1 4413
0 4415 7 4 2 22925 28355
0 4416 7 1 2 28437 27670
0 4417 7 1 2 26602 4416
0 4418 7 1 2 32404 4417
0 4419 5 1 1 4418
0 4420 7 1 2 4414 4419
0 4421 5 1 1 4420
0 4422 7 1 2 24556 27354
0 4423 7 1 2 4421 4422
0 4424 5 1 1 4423
0 4425 7 1 2 4401 4424
0 4426 5 1 1 4425
0 4427 7 1 2 27072 4426
0 4428 5 1 1 4427
0 4429 7 1 2 4394 4428
0 4430 7 1 2 4391 4429
0 4431 5 1 1 4430
0 4432 7 1 2 24427 4431
0 4433 5 1 1 4432
0 4434 7 1 2 32386 31788
0 4435 5 1 1 4434
0 4436 7 1 2 22926 31739
0 4437 7 1 2 30958 4436
0 4438 7 1 2 31758 4437
0 4439 5 1 1 4438
0 4440 7 1 2 4435 4439
0 4441 5 1 1 4440
0 4442 7 1 2 27920 4441
0 4443 5 1 1 4442
0 4444 7 1 2 31214 31764
0 4445 5 1 1 4444
0 4446 7 1 2 31767 32403
0 4447 5 1 1 4446
0 4448 7 1 2 4445 4447
0 4449 5 1 1 4448
0 4450 7 1 2 27734 4449
0 4451 5 1 1 4450
0 4452 7 1 2 25674 4451
0 4453 7 1 2 4443 4452
0 4454 7 1 2 4433 4453
0 4455 5 1 1 4454
0 4456 7 1 2 23100 31803
0 4457 5 1 1 4456
0 4458 7 1 2 28890 28036
0 4459 7 3 2 23244 28438
0 4460 7 3 2 30973 29372
0 4461 7 1 2 32408 32411
0 4462 7 1 2 4458 4461
0 4463 5 1 1 4462
0 4464 7 1 2 4457 4463
0 4465 5 1 1 4464
0 4466 7 1 2 31215 4465
0 4467 5 1 1 4466
0 4468 7 1 2 23681 4467
0 4469 5 1 1 4468
0 4470 7 1 2 26799 4469
0 4471 7 1 2 4455 4470
0 4472 5 1 1 4471
0 4473 7 1 2 4354 4472
0 4474 7 1 2 4299 4473
0 4475 5 1 1 4474
0 4476 7 1 2 26506 4475
0 4477 5 1 1 4476
0 4478 7 1 2 32044 4477
0 4479 7 1 2 4011 4478
0 4480 7 1 2 3276 4479
0 4481 7 1 2 3018 4480
0 4482 7 1 2 1107 4481
0 4483 5 1 1 4482
0 4484 7 1 2 29360 30937
0 4485 5 1 1 4484
0 4486 7 4 2 25351 27167
0 4487 7 1 2 28016 32414
0 4488 5 1 1 4487
0 4489 7 1 2 4485 4488
0 4490 5 1 1 4489
0 4491 7 1 2 23245 4490
0 4492 5 1 1 4491
0 4493 7 3 2 23394 25757
0 4494 7 3 2 23996 32418
0 4495 7 1 2 31579 32421
0 4496 5 1 1 4495
0 4497 7 1 2 4492 4496
0 4498 5 1 1 4497
0 4499 7 1 2 23901 4498
0 4500 5 1 1 4499
0 4501 7 1 2 25283 30938
0 4502 5 1 1 4501
0 4503 7 1 2 27046 28872
0 4504 5 2 1 4503
0 4505 7 1 2 4502 32424
0 4506 5 1 1 4505
0 4507 7 2 2 23246 27234
0 4508 7 1 2 4506 32426
0 4509 5 1 1 4508
0 4510 7 1 2 4500 4509
0 4511 5 1 1 4510
0 4512 7 1 2 22573 4511
0 4513 5 1 1 4512
0 4514 7 1 2 23332 32178
0 4515 5 1 1 4514
0 4516 7 1 2 30866 32422
0 4517 5 1 1 4516
0 4518 7 1 2 4515 4517
0 4519 5 1 1 4518
0 4520 7 1 2 30640 4519
0 4521 5 1 1 4520
0 4522 7 1 2 4513 4521
0 4523 5 1 1 4522
0 4524 7 1 2 22407 4523
0 4525 5 1 1 4524
0 4526 7 2 2 24428 27842
0 4527 7 3 2 32428 32157
0 4528 5 1 1 32430
0 4529 7 1 2 32185 32431
0 4530 5 1 1 4529
0 4531 7 1 2 4525 4530
0 4532 5 3 1 4531
0 4533 7 6 2 25413 26054
0 4534 5 1 1 32436
0 4535 7 6 2 23450 24083
0 4536 5 2 1 32442
0 4537 7 1 2 4534 32448
0 4538 5 13 1 4537
0 4539 7 3 2 22790 32450
0 4540 5 1 1 32463
0 4541 7 9 2 23451 26055
0 4542 5 2 1 32466
0 4543 7 2 2 24737 32467
0 4544 5 1 1 32477
0 4545 7 1 2 4540 4544
0 4546 5 15 1 4545
0 4547 7 1 2 32433 32479
0 4548 5 1 1 4547
0 4549 7 2 2 28120 32198
0 4550 5 1 1 32494
0 4551 7 3 2 23780 28230
0 4552 5 1 1 32496
0 4553 7 1 2 27407 26910
0 4554 5 1 1 4553
0 4555 7 2 2 28630 4554
0 4556 5 3 1 32499
0 4557 7 1 2 32497 32501
0 4558 5 1 1 4557
0 4559 7 1 2 4550 4558
0 4560 5 2 1 4559
0 4561 7 2 2 24084 28195
0 4562 7 1 2 26887 32506
0 4563 7 1 2 32504 4562
0 4564 5 1 1 4563
0 4565 7 1 2 4548 4564
0 4566 5 1 1 4565
0 4567 7 1 2 29387 4566
0 4568 5 1 1 4567
0 4569 7 12 2 24738 26056
0 4570 5 1 1 32508
0 4571 7 16 2 22791 24085
0 4572 5 1 1 32520
0 4573 7 2 2 4570 4572
0 4574 5 26 1 32536
0 4575 7 5 2 24173 32538
0 4576 7 1 2 28865 1835
0 4577 5 28 1 4576
0 4578 7 4 2 25873 32569
0 4579 7 1 2 31263 32597
0 4580 5 1 1 4579
0 4581 7 1 2 27454 32186
0 4582 5 1 1 4581
0 4583 7 1 2 4580 4582
0 4584 5 5 1 4583
0 4585 7 15 2 25414 25482
0 4586 5 1 1 32606
0 4587 7 6 2 25352 32607
0 4588 7 1 2 30379 32621
0 4589 5 1 1 4588
0 4590 7 16 2 23452 23524
0 4591 5 1 1 32627
0 4592 7 6 2 23395 32628
0 4593 7 1 2 32643 30403
0 4594 5 1 1 4593
0 4595 7 1 2 4589 4594
0 4596 5 11 1 4595
0 4597 7 1 2 32601 32649
0 4598 5 1 1 4597
0 4599 7 5 2 31668 32570
0 4600 7 2 2 23781 32660
0 4601 7 2 2 29054 28883
0 4602 7 1 2 32665 32667
0 4603 5 1 1 4602
0 4604 7 2 2 24853 28668
0 4605 7 1 2 27843 32608
0 4606 7 1 2 32187 4605
0 4607 7 1 2 32669 4606
0 4608 5 1 1 4607
0 4609 7 1 2 4603 4608
0 4610 7 1 2 4598 4609
0 4611 5 1 1 4610
0 4612 7 1 2 28196 4611
0 4613 5 1 1 4612
0 4614 7 3 2 23333 29373
0 4615 7 1 2 30071 32671
0 4616 5 1 1 4615
0 4617 7 2 2 22574 27886
0 4618 7 1 2 27906 32674
0 4619 5 1 1 4618
0 4620 7 1 2 4616 4619
0 4621 5 1 1 4620
0 4622 7 1 2 27168 32000
0 4623 7 1 2 32644 4622
0 4624 7 1 2 4621 4623
0 4625 5 1 1 4624
0 4626 7 1 2 4613 4625
0 4627 5 1 1 4626
0 4628 7 1 2 32564 4627
0 4629 5 1 1 4628
0 4630 7 1 2 4568 4629
0 4631 5 1 1 4630
0 4632 7 1 2 26603 4631
0 4633 5 1 1 4632
0 4634 7 4 2 24854 28071
0 4635 7 1 2 32676 32622
0 4636 5 1 1 4635
0 4637 7 1 2 23334 27371
0 4638 7 1 2 32645 4637
0 4639 5 1 1 4638
0 4640 7 1 2 4636 4639
0 4641 5 5 1 4640
0 4642 7 1 2 22575 32680
0 4643 5 1 1 4642
0 4644 7 1 2 30641 32650
0 4645 5 1 1 4644
0 4646 7 1 2 4643 4645
0 4647 5 1 1 4646
0 4648 7 1 2 22408 4647
0 4649 5 1 1 4648
0 4650 7 5 2 28031 28603
0 4651 7 2 2 27472 32685
0 4652 5 1 1 32690
0 4653 7 1 2 22576 32691
0 4654 5 1 1 4653
0 4655 7 1 2 4649 4654
0 4656 5 2 1 4655
0 4657 7 3 2 26966 29950
0 4658 7 2 2 22792 23028
0 4659 7 5 2 24666 25758
0 4660 7 1 2 32697 32699
0 4661 7 1 2 32694 4660
0 4662 7 1 2 32692 4661
0 4663 5 1 1 4662
0 4664 7 1 2 4633 4663
0 4665 5 1 1 4664
0 4666 7 1 2 23101 4665
0 4667 5 1 1 4666
0 4668 7 6 2 23453 25483
0 4669 7 2 2 24855 32704
0 4670 5 1 1 32710
0 4671 7 5 2 25415 23525
0 4672 7 3 2 22927 32712
0 4673 5 1 1 32717
0 4674 7 1 2 4670 4673
0 4675 5 23 1 4674
0 4676 7 2 2 356 4031
0 4677 7 4 2 25284 24086
0 4678 5 1 1 32745
0 4679 7 1 2 4678 32537
0 4680 7 4 2 32743 4679
0 4681 7 1 2 32602 32749
0 4682 5 1 1 4681
0 4683 7 14 2 22793 26057
0 4684 5 1 1 32753
0 4685 7 4 2 27384 32754
0 4686 7 3 2 23782 32767
0 4687 5 1 1 32771
0 4688 7 1 2 32661 32772
0 4689 5 1 1 4688
0 4690 7 3 2 31421 29888
0 4691 5 1 1 32774
0 4692 7 4 2 25353 25759
0 4693 7 1 2 30867 32777
0 4694 7 1 2 32775 4693
0 4695 5 1 1 4694
0 4696 7 1 2 4689 4695
0 4697 7 2 2 4682 4696
0 4698 5 1 1 32781
0 4699 7 2 2 27142 30682
0 4700 5 1 1 32783
0 4701 7 1 2 4094 4700
0 4702 5 2 1 4701
0 4703 7 1 2 28121 32785
0 4704 5 1 1 4703
0 4705 7 5 2 24667 26939
0 4706 5 1 1 32787
0 4707 7 6 2 22704 26967
0 4708 5 1 1 32792
0 4709 7 1 2 4706 4708
0 4710 5 14 1 4709
0 4711 7 2 2 32798 32498
0 4712 5 1 1 32812
0 4713 7 1 2 4704 4712
0 4714 5 4 1 4713
0 4715 7 6 2 24739 23396
0 4716 7 2 2 24087 32818
0 4717 5 3 1 32824
0 4718 7 2 2 22794 32133
0 4719 5 1 1 32829
0 4720 7 1 2 32826 4719
0 4721 5 6 1 4720
0 4722 7 1 2 32814 32831
0 4723 5 1 1 4722
0 4724 7 1 2 32782 4723
0 4725 5 1 1 4724
0 4726 7 1 2 23247 4725
0 4727 5 1 1 4726
0 4728 7 2 2 29208 31495
0 4729 7 1 2 32380 32423
0 4730 7 1 2 32837 4729
0 4731 5 1 1 4730
0 4732 7 1 2 4727 4731
0 4733 5 1 1 4732
0 4734 7 1 2 22409 4733
0 4735 5 1 1 4734
0 4736 7 2 2 31496 27907
0 4737 7 4 2 23397 23902
0 4738 7 1 2 27862 29867
0 4739 7 1 2 32841 4738
0 4740 7 1 2 32839 4739
0 4741 5 1 1 4740
0 4742 7 1 2 4735 4741
0 4743 5 1 1 4742
0 4744 7 1 2 26604 4743
0 4745 5 1 1 4744
0 4746 7 1 2 31008 28072
0 4747 5 1 1 4746
0 4748 7 1 2 25201 32033
0 4749 5 1 1 4748
0 4750 7 1 2 4747 4749
0 4751 5 9 1 4750
0 4752 7 1 2 22577 32845
0 4753 5 1 1 4752
0 4754 7 1 2 32235 30642
0 4755 5 1 1 4754
0 4756 7 1 2 4753 4755
0 4757 5 3 1 4756
0 4758 7 1 2 22410 32854
0 4759 5 1 1 4758
0 4760 7 1 2 4759 4528
0 4761 5 5 1 4760
0 4762 7 3 2 32857 32220
0 4763 7 1 2 24740 32359
0 4764 7 1 2 32862 4763
0 4765 5 1 1 4764
0 4766 7 1 2 4745 4765
0 4767 5 1 1 4766
0 4768 7 1 2 23102 4767
0 4769 5 1 1 4768
0 4770 7 2 2 24741 23903
0 4771 5 1 1 32865
0 4772 7 5 2 23904 30328
0 4773 5 1 1 32867
0 4774 7 5 2 24742 29889
0 4775 5 1 1 32872
0 4776 7 1 2 4773 4775
0 4777 5 1 1 4776
0 4778 7 7 2 4771 4777
0 4779 7 2 2 29150 32877
0 4780 5 2 1 32884
0 4781 7 4 2 25964 28122
0 4782 7 2 2 32755 32888
0 4783 7 1 2 30199 32892
0 4784 5 1 1 4783
0 4785 7 1 2 32886 4784
0 4786 5 1 1 4785
0 4787 7 1 2 32073 4786
0 4788 5 1 1 4787
0 4789 7 1 2 22578 32236
0 4790 5 1 1 4789
0 4791 7 1 2 3714 4790
0 4792 5 11 1 4791
0 4793 7 1 2 27949 32894
0 4794 5 2 1 4793
0 4795 7 4 2 28669 31186
0 4796 7 1 2 28197 32907
0 4797 5 1 1 4796
0 4798 7 1 2 32905 4797
0 4799 5 5 1 4798
0 4800 7 5 2 22795 29868
0 4801 5 2 1 32916
0 4802 7 4 2 24743 29825
0 4803 5 1 1 32923
0 4804 7 1 2 32921 4803
0 4805 5 12 1 4804
0 4806 7 1 2 25874 32927
0 4807 7 1 2 32911 4806
0 4808 5 1 1 4807
0 4809 7 1 2 4788 4808
0 4810 5 1 1 4809
0 4811 7 1 2 31736 4810
0 4812 5 1 1 4811
0 4813 7 1 2 4769 4812
0 4814 5 1 1 4813
0 4815 7 1 2 24174 4814
0 4816 5 1 1 4815
0 4817 7 1 2 32799 29151
0 4818 5 1 1 4817
0 4819 7 4 2 29753 30767
0 4820 7 1 2 28123 32939
0 4821 5 1 1 4820
0 4822 7 1 2 4818 4821
0 4823 5 4 1 4822
0 4824 7 1 2 32832 32943
0 4825 5 1 1 4824
0 4826 7 2 2 26968 28198
0 4827 7 1 2 31187 32947
0 4828 5 1 1 4827
0 4829 7 2 2 32571 31942
0 4830 7 1 2 27950 32949
0 4831 5 1 1 4830
0 4832 7 1 2 4828 4831
0 4833 5 4 1 4832
0 4834 7 1 2 32750 32951
0 4835 5 1 1 4834
0 4836 7 3 2 31655 32572
0 4837 5 1 1 32955
0 4838 7 3 2 26969 31031
0 4839 5 1 1 32958
0 4840 7 1 2 4837 4839
0 4841 5 6 1 4840
0 4842 7 2 2 25285 31275
0 4843 7 5 2 25354 24088
0 4844 7 1 2 32967 32969
0 4845 5 1 1 4844
0 4846 7 1 2 25202 32768
0 4847 5 1 1 4846
0 4848 7 1 2 4845 4847
0 4849 5 1 1 4848
0 4850 7 1 2 22411 4849
0 4851 5 1 1 4850
0 4852 7 2 2 24429 31693
0 4853 7 3 2 23398 26058
0 4854 7 1 2 23335 32976
0 4855 7 1 2 32974 4854
0 4856 5 1 1 4855
0 4857 7 1 2 4851 4856
0 4858 5 3 1 4857
0 4859 7 1 2 32961 32979
0 4860 5 1 1 4859
0 4861 7 1 2 4835 4860
0 4862 7 1 2 4825 4861
0 4863 5 1 1 4862
0 4864 7 1 2 29181 31337
0 4865 7 1 2 4863 4864
0 4866 5 1 1 4865
0 4867 7 1 2 4816 4866
0 4868 5 1 1 4867
0 4869 7 1 2 32720 4868
0 4870 5 1 1 4869
0 4871 7 17 2 26141 26233
0 4872 7 4 2 23029 32982
0 4873 7 1 2 30807 29152
0 4874 5 1 1 4873
0 4875 7 1 2 2002 4874
0 4876 5 1 1 4875
0 4877 7 1 2 32999 4876
0 4878 5 1 1 4877
0 4879 7 5 2 24089 26940
0 4880 7 1 2 33003 32286
0 4881 7 1 2 29153 4880
0 4882 5 1 1 4881
0 4883 7 1 2 4878 4882
0 4884 5 1 1 4883
0 4885 7 1 2 32074 4884
0 4886 5 1 1 4885
0 4887 7 4 2 26059 26234
0 4888 7 4 2 23997 33008
0 4889 7 2 2 33012 29312
0 4890 5 2 1 33016
0 4891 7 2 2 26572 30236
0 4892 5 1 1 33020
0 4893 7 1 2 33018 4892
0 4894 5 1 1 4893
0 4895 7 1 2 25875 4894
0 4896 7 1 2 32912 4895
0 4897 5 1 1 4896
0 4898 7 1 2 4886 4897
0 4899 5 1 1 4898
0 4900 7 1 2 28972 4899
0 4901 5 1 1 4900
0 4902 7 3 2 1551 27498
0 4903 7 1 2 413 4343
0 4904 5 1 1 4903
0 4905 7 2 2 33022 4904
0 4906 7 1 2 28721 32944
0 4907 5 1 1 4906
0 4908 7 1 2 28821 32952
0 4909 5 1 1 4908
0 4910 7 2 2 31276 31991
0 4911 5 1 1 33027
0 4912 7 4 2 25203 27385
0 4913 7 2 2 26338 33029
0 4914 5 1 1 33033
0 4915 7 1 2 4911 4914
0 4916 5 5 1 4915
0 4917 7 1 2 22412 33035
0 4918 5 1 1 4917
0 4919 7 5 2 24430 22796
0 4920 7 2 2 33040 28403
0 4921 5 1 1 33045
0 4922 7 1 2 4918 4921
0 4923 5 3 1 4922
0 4924 7 1 2 33047 32962
0 4925 5 1 1 4924
0 4926 7 1 2 4909 4925
0 4927 7 1 2 4907 4926
0 4928 5 2 1 4927
0 4929 7 1 2 33025 33050
0 4930 5 1 1 4929
0 4931 7 1 2 4901 4930
0 4932 5 1 1 4931
0 4933 7 1 2 29101 4932
0 4934 5 1 1 4933
0 4935 7 1 2 4591 2702
0 4936 5 1 1 4935
0 4937 7 1 2 4586 198
0 4938 5 1 1 4937
0 4939 7 14 2 4936 4938
0 4940 7 3 2 28124 32539
0 4941 7 3 2 23030 29813
0 4942 5 2 1 33069
0 4943 7 1 2 33072 32270
0 4944 5 6 1 4943
0 4945 7 1 2 32940 33074
0 4946 5 1 1 4945
0 4947 7 2 2 27784 30690
0 4948 7 5 2 24175 31112
0 4949 7 1 2 33082 26605
0 4950 7 1 2 33080 4949
0 4951 5 1 1 4950
0 4952 7 1 2 4946 4951
0 4953 5 1 1 4952
0 4954 7 1 2 33066 4953
0 4955 5 1 1 4954
0 4956 7 1 2 32800 32269
0 4957 5 1 1 4956
0 4958 7 1 2 32788 33070
0 4959 5 1 1 4958
0 4960 7 1 2 4957 4959
0 4961 5 1 1 4960
0 4962 7 1 2 32540 4961
0 4963 5 1 1 4962
0 4964 7 3 2 26235 32509
0 4965 5 1 1 33087
0 4966 7 1 2 22797 27671
0 4967 5 1 1 4966
0 4968 7 1 2 4965 4967
0 4969 5 1 1 4968
0 4970 7 1 2 32793 30246
0 4971 7 1 2 4969 4970
0 4972 5 1 1 4971
0 4973 7 1 2 4963 4972
0 4974 5 1 1 4973
0 4975 7 1 2 29154 4974
0 4976 5 1 1 4975
0 4977 7 1 2 4955 4976
0 4978 5 1 1 4977
0 4979 7 1 2 33052 4978
0 4980 5 1 1 4979
0 4981 7 7 2 22579 27951
0 4982 7 4 2 25876 33090
0 4983 7 7 2 32573 32541
0 4984 7 1 2 33097 33101
0 4985 5 1 1 4984
0 4986 7 2 2 25965 30778
0 4987 7 1 2 26060 30691
0 4988 7 1 2 32343 4987
0 4989 7 1 2 33108 4988
0 4990 5 1 1 4989
0 4991 7 1 2 4985 4990
0 4992 5 1 1 4991
0 4993 7 1 2 32651 4992
0 4994 5 1 1 4993
0 4995 7 1 2 22413 32681
0 4996 5 1 1 4995
0 4997 7 1 2 4652 4996
0 4998 5 4 1 4997
0 4999 7 1 2 30808 31353
0 5000 5 1 1 4999
0 5001 7 1 2 31656 33102
0 5002 5 1 1 5001
0 5003 7 1 2 5000 5002
0 5004 5 1 1 5003
0 5005 7 1 2 33110 5004
0 5006 5 1 1 5005
0 5007 7 1 2 4994 5006
0 5008 5 1 1 5007
0 5009 7 1 2 33075 5008
0 5010 5 1 1 5009
0 5011 7 2 2 22798 23905
0 5012 7 4 2 25966 33114
0 5013 7 1 2 33116 32218
0 5014 7 1 2 32693 5013
0 5015 5 1 1 5014
0 5016 7 1 2 5010 5015
0 5017 7 1 2 4980 5016
0 5018 7 1 2 4934 5017
0 5019 5 1 1 5018
0 5020 7 1 2 25760 5019
0 5021 5 1 1 5020
0 5022 7 1 2 27305 28765
0 5023 5 1 1 5022
0 5024 7 1 2 26941 28873
0 5025 5 2 1 5024
0 5026 7 1 2 5023 33120
0 5027 5 1 1 5026
0 5028 7 1 2 22580 5027
0 5029 5 1 1 5028
0 5030 7 3 2 24557 27433
0 5031 5 1 1 33122
0 5032 7 2 2 28766 33123
0 5033 5 1 1 33125
0 5034 7 1 2 5029 5033
0 5035 5 5 1 5034
0 5036 7 1 2 28199 31745
0 5037 7 1 2 33053 5036
0 5038 7 1 2 32565 5037
0 5039 7 1 2 33127 5038
0 5040 5 1 1 5039
0 5041 7 1 2 5021 5040
0 5042 7 1 2 4870 5041
0 5043 7 1 2 4667 5042
0 5044 5 1 1 5043
0 5045 7 1 2 26507 5044
0 5046 5 1 1 5045
0 5047 7 7 2 24744 24090
0 5048 5 1 1 33132
0 5049 7 15 2 4684 5048
0 5050 7 1 2 26822 28465
0 5051 5 1 1 5050
0 5052 7 1 2 1385 5051
0 5053 5 3 1 5052
0 5054 7 1 2 32956 33154
0 5055 5 1 1 5054
0 5056 7 9 2 25967 26142
0 5057 7 4 2 24668 33157
0 5058 7 1 2 33166 29576
0 5059 5 1 1 5058
0 5060 7 2 2 29785 29182
0 5061 5 1 1 33170
0 5062 7 1 2 29509 5061
0 5063 5 2 1 5062
0 5064 7 2 2 23998 33172
0 5065 7 1 2 22705 33174
0 5066 5 1 1 5065
0 5067 7 1 2 5059 5066
0 5068 5 1 1 5067
0 5069 7 2 2 23906 5068
0 5070 7 1 2 22581 33176
0 5071 5 1 1 5070
0 5072 7 1 2 5055 5071
0 5073 5 1 1 5072
0 5074 7 1 2 33111 5073
0 5075 5 1 1 5074
0 5076 7 5 2 23454 26143
0 5077 5 1 1 33178
0 5078 7 3 2 33179 26823
0 5079 7 2 2 22706 26374
0 5080 5 1 1 33186
0 5081 7 5 2 25968 32075
0 5082 7 1 2 23103 33188
0 5083 5 1 1 5082
0 5084 7 1 2 5080 5083
0 5085 5 3 1 5084
0 5086 7 1 2 25286 33193
0 5087 5 1 1 5086
0 5088 7 1 2 32425 5087
0 5089 5 1 1 5088
0 5090 7 1 2 24558 5089
0 5091 5 1 1 5090
0 5092 7 1 2 31086 30390
0 5093 5 1 1 5092
0 5094 7 1 2 5091 5093
0 5095 5 1 1 5094
0 5096 7 1 2 28200 5095
0 5097 5 1 1 5096
0 5098 7 1 2 22582 29136
0 5099 7 1 2 33194 5098
0 5100 5 1 1 5099
0 5101 7 1 2 5097 5100
0 5102 5 1 1 5101
0 5103 7 1 2 33183 5102
0 5104 5 1 1 5103
0 5105 7 3 2 29273 29786
0 5106 7 4 2 23248 25416
0 5107 7 2 2 22414 33199
0 5108 7 1 2 23999 33203
0 5109 7 1 2 32143 5108
0 5110 7 1 2 33196 5109
0 5111 5 1 1 5110
0 5112 7 1 2 23907 5111
0 5113 7 1 2 5104 5112
0 5114 5 1 1 5113
0 5115 7 2 2 24176 29577
0 5116 7 1 2 24669 25417
0 5117 7 1 2 29155 5116
0 5118 7 1 2 33205 5117
0 5119 5 1 1 5118
0 5120 7 1 2 30311 30183
0 5121 7 1 2 33184 5120
0 5122 5 1 1 5121
0 5123 7 1 2 5119 5122
0 5124 5 1 1 5123
0 5125 7 1 2 27073 5124
0 5126 5 1 1 5125
0 5127 7 1 2 28009 33206
0 5128 5 1 1 5127
0 5129 7 3 2 24670 23104
0 5130 7 1 2 33207 33185
0 5131 5 1 1 5130
0 5132 7 1 2 5128 5131
0 5133 5 1 1 5132
0 5134 7 1 2 348 28917
0 5135 5 5 1 5134
0 5136 7 1 2 22583 33210
0 5137 5 1 1 5136
0 5138 7 1 2 5137 359
0 5139 5 2 1 5138
0 5140 7 1 2 27952 33215
0 5141 5 1 1 5140
0 5142 7 3 2 28073 27047
0 5143 5 1 1 33217
0 5144 7 1 2 28052 33218
0 5145 5 1 1 5144
0 5146 7 1 2 5141 5145
0 5147 5 1 1 5146
0 5148 7 1 2 5133 5147
0 5149 5 1 1 5148
0 5150 7 1 2 25877 5149
0 5151 7 1 2 5126 5150
0 5152 5 1 1 5151
0 5153 7 1 2 29102 5152
0 5154 7 1 2 5114 5153
0 5155 5 1 1 5154
0 5156 7 1 2 5075 5155
0 5157 5 1 1 5156
0 5158 7 1 2 25761 5157
0 5159 5 1 1 5158
0 5160 7 7 2 23783 28201
0 5161 7 2 2 26144 32662
0 5162 7 1 2 33227 32668
0 5163 5 1 1 5162
0 5164 7 1 2 23336 32502
0 5165 5 1 1 5164
0 5166 7 1 2 27019 30991
0 5167 5 1 1 5166
0 5168 7 1 2 5165 5167
0 5169 5 1 1 5168
0 5170 7 1 2 22584 5169
0 5171 5 1 1 5170
0 5172 7 1 2 27154 28781
0 5173 5 1 1 5172
0 5174 7 1 2 5171 5173
0 5175 5 3 1 5174
0 5176 7 2 2 25418 29103
0 5177 7 1 2 24177 33232
0 5178 7 1 2 33229 5177
0 5179 5 1 1 5178
0 5180 7 1 2 5163 5179
0 5181 5 1 1 5180
0 5182 7 1 2 29558 5181
0 5183 5 1 1 5182
0 5184 7 1 2 22585 27306
0 5185 5 1 1 5184
0 5186 7 1 2 5031 5185
0 5187 5 13 1 5186
0 5188 7 1 2 33234 29388
0 5189 5 1 1 5188
0 5190 7 3 2 23337 31669
0 5191 7 1 2 29446 33247
0 5192 5 1 1 5191
0 5193 7 1 2 5189 5192
0 5194 5 1 1 5193
0 5195 7 1 2 23399 32574
0 5196 7 1 2 5194 5195
0 5197 5 1 1 5196
0 5198 7 1 2 25355 29389
0 5199 7 1 2 33128 5198
0 5200 5 1 1 5199
0 5201 7 1 2 5197 5200
0 5202 5 1 1 5201
0 5203 7 1 2 23455 26824
0 5204 7 1 2 5202 5203
0 5205 5 1 1 5204
0 5206 7 1 2 5183 5205
0 5207 5 1 1 5206
0 5208 7 1 2 33220 5207
0 5209 5 1 1 5208
0 5210 7 1 2 5159 5209
0 5211 5 1 1 5210
0 5212 7 1 2 33139 5211
0 5213 5 1 1 5212
0 5214 7 6 2 24745 25042
0 5215 5 1 1 33250
0 5216 7 1 2 5215 31440
0 5217 5 1 1 5216
0 5218 7 3 2 26061 24330
0 5219 5 1 1 33256
0 5220 7 1 2 26713 5219
0 5221 5 1 1 5220
0 5222 7 1 2 5217 5221
0 5223 5 1 1 5222
0 5224 7 1 2 32221 32566
0 5225 7 3 2 5223 5224
0 5226 7 1 2 30664 33259
0 5227 5 1 1 5226
0 5228 7 1 2 32801 29581
0 5229 5 1 1 5228
0 5230 7 2 2 26942 33208
0 5231 7 1 2 29507 33262
0 5232 5 1 1 5231
0 5233 7 1 2 5229 5232
0 5234 5 1 1 5233
0 5235 7 1 2 29156 5234
0 5236 5 1 1 5235
0 5237 7 1 2 30785 33175
0 5238 5 1 1 5237
0 5239 7 2 2 25969 30683
0 5240 7 2 2 27953 33155
0 5241 7 1 2 33264 33266
0 5242 5 1 1 5241
0 5243 7 1 2 5238 5242
0 5244 5 1 1 5243
0 5245 7 1 2 28125 5244
0 5246 5 1 1 5245
0 5247 7 1 2 5236 5246
0 5248 5 1 1 5247
0 5249 7 1 2 25762 5248
0 5250 5 1 1 5249
0 5251 7 3 2 33221 33173
0 5252 5 1 1 33268
0 5253 7 1 2 33129 33269
0 5254 5 1 1 5253
0 5255 7 1 2 5250 5254
0 5256 5 2 1 5255
0 5257 7 1 2 33140 33271
0 5258 5 1 1 5257
0 5259 7 1 2 5227 5258
0 5260 5 1 1 5259
0 5261 7 1 2 33054 5260
0 5262 5 1 1 5261
0 5263 7 1 2 25763 33267
0 5264 5 1 1 5263
0 5265 7 1 2 5252 5264
0 5266 5 1 1 5265
0 5267 7 1 2 32950 5266
0 5268 5 1 1 5267
0 5269 7 6 2 23249 25764
0 5270 5 1 1 33273
0 5271 7 4 2 28053 33274
0 5272 7 1 2 33279 33177
0 5273 5 1 1 5272
0 5274 7 1 2 5268 5273
0 5275 5 2 1 5274
0 5276 7 1 2 32542 33283
0 5277 5 1 1 5276
0 5278 7 7 2 23250 28054
0 5279 7 2 2 24671 33285
0 5280 7 1 2 33292 33260
0 5281 5 1 1 5280
0 5282 7 1 2 5277 5281
0 5283 5 1 1 5282
0 5284 7 1 2 32652 5283
0 5285 5 1 1 5284
0 5286 7 1 2 31032 33112
0 5287 7 1 2 33261 5286
0 5288 5 1 1 5287
0 5289 7 1 2 5285 5288
0 5290 7 1 2 5262 5289
0 5291 7 1 2 5213 5290
0 5292 7 2 2 31062 26810
0 5293 7 3 2 25419 33294
0 5294 5 1 1 33296
0 5295 7 1 2 23456 33197
0 5296 5 1 1 5295
0 5297 7 1 2 5294 5296
0 5298 5 2 1 5297
0 5299 7 2 2 33222 33299
0 5300 5 1 1 33301
0 5301 7 1 2 23105 33297
0 5302 5 1 1 5301
0 5303 7 3 2 23457 24178
0 5304 5 3 1 33303
0 5305 7 1 2 33304 29578
0 5306 5 1 1 5305
0 5307 7 1 2 5302 5306
0 5308 5 2 1 5307
0 5309 7 2 2 27954 33309
0 5310 7 1 2 25765 33311
0 5311 5 1 1 5310
0 5312 7 1 2 5300 5311
0 5313 5 1 1 5312
0 5314 7 1 2 31943 5313
0 5315 5 1 1 5314
0 5316 7 1 2 33280 27743
0 5317 7 1 2 33198 5316
0 5318 5 1 1 5317
0 5319 7 1 2 5315 5318
0 5320 5 1 1 5319
0 5321 7 1 2 32928 5320
0 5322 5 1 1 5321
0 5323 7 1 2 23106 32924
0 5324 5 1 1 5323
0 5325 7 1 2 32922 5324
0 5326 5 1 1 5325
0 5327 7 1 2 33295 5326
0 5328 5 1 1 5327
0 5329 7 1 2 32510 29569
0 5330 5 1 1 5329
0 5331 7 1 2 26062 29564
0 5332 5 1 1 5331
0 5333 7 1 2 32543 5332
0 5334 7 1 2 29559 5333
0 5335 5 1 1 5334
0 5336 7 1 2 5330 5335
0 5337 5 1 1 5336
0 5338 7 1 2 30191 5337
0 5339 5 1 1 5338
0 5340 7 1 2 5328 5339
0 5341 5 1 1 5340
0 5342 7 2 2 23908 5341
0 5343 7 1 2 25420 33281
0 5344 7 1 2 33313 5343
0 5345 5 1 1 5344
0 5346 7 1 2 5322 5345
0 5347 5 1 1 5346
0 5348 7 1 2 32237 5347
0 5349 5 1 1 5348
0 5350 7 2 2 22415 32846
0 5351 5 1 1 33315
0 5352 7 1 2 24431 30974
0 5353 7 2 2 28356 5352
0 5354 5 1 1 33317
0 5355 7 1 2 5351 5354
0 5356 5 8 1 5355
0 5357 7 1 2 31657 29570
0 5358 5 1 1 5357
0 5359 7 1 2 25878 29565
0 5360 5 1 1 5359
0 5361 7 1 2 31670 5360
0 5362 7 1 2 29560 5361
0 5363 5 1 1 5362
0 5364 7 1 2 5358 5363
0 5365 5 1 1 5364
0 5366 7 1 2 33305 5365
0 5367 5 1 1 5366
0 5368 7 6 2 24559 23107
0 5369 7 2 2 25879 33327
0 5370 5 1 1 33333
0 5371 7 1 2 33298 33334
0 5372 5 1 1 5371
0 5373 7 1 2 5367 5372
0 5374 5 1 1 5373
0 5375 7 1 2 32929 5374
0 5376 5 1 1 5375
0 5377 7 3 2 22586 25421
0 5378 7 1 2 33335 33314
0 5379 5 1 1 5378
0 5380 7 1 2 5376 5379
0 5381 5 1 1 5380
0 5382 7 1 2 33319 5381
0 5383 5 1 1 5382
0 5384 7 1 2 32885 33310
0 5385 5 1 1 5384
0 5386 7 1 2 29754 32756
0 5387 7 1 2 33312 5386
0 5388 5 1 1 5387
0 5389 7 4 2 24000 32866
0 5390 7 1 2 33338 32507
0 5391 7 1 2 33300 5390
0 5392 5 1 1 5391
0 5393 7 1 2 5388 5392
0 5394 5 1 1 5393
0 5395 7 1 2 28126 5394
0 5396 5 1 1 5395
0 5397 7 1 2 5385 5396
0 5398 5 1 1 5397
0 5399 7 1 2 32076 5398
0 5400 5 1 1 5399
0 5401 7 1 2 5383 5400
0 5402 5 1 1 5401
0 5403 7 1 2 25766 5402
0 5404 5 1 1 5403
0 5405 7 2 2 29929 28836
0 5406 5 1 1 33342
0 5407 7 1 2 33004 27418
0 5408 5 1 1 5407
0 5409 7 1 2 22799 30329
0 5410 7 1 2 27307 5409
0 5411 5 1 1 5410
0 5412 7 1 2 5408 5411
0 5413 5 1 1 5412
0 5414 7 1 2 22587 5413
0 5415 5 1 1 5414
0 5416 7 1 2 5406 5415
0 5417 5 1 1 5416
0 5418 7 1 2 32077 5417
0 5419 5 1 1 5418
0 5420 7 1 2 30975 32930
0 5421 7 1 2 33248 5420
0 5422 5 1 1 5421
0 5423 7 1 2 5419 5422
0 5424 5 1 1 5423
0 5425 7 1 2 33302 5424
0 5426 5 1 1 5425
0 5427 7 1 2 5404 5426
0 5428 7 1 2 5349 5427
0 5429 5 1 1 5428
0 5430 7 1 2 29104 5429
0 5431 5 1 1 5430
0 5432 7 1 2 32833 33272
0 5433 5 1 1 5432
0 5434 7 4 2 24672 25043
0 5435 7 2 2 25970 33344
0 5436 5 1 1 33348
0 5437 7 1 2 29630 33349
0 5438 5 1 1 5437
0 5439 7 2 2 26308 28848
0 5440 7 1 2 29814 33350
0 5441 5 1 1 5440
0 5442 7 1 2 5438 5441
0 5443 5 1 1 5442
0 5444 7 1 2 23620 5443
0 5445 5 1 1 5444
0 5446 7 1 2 28849 29787
0 5447 5 1 1 5446
0 5448 7 1 2 25620 30164
0 5449 7 1 2 29743 5448
0 5450 5 1 1 5449
0 5451 7 1 2 5447 5450
0 5452 5 1 1 5451
0 5453 7 1 2 24261 5452
0 5454 5 1 1 5453
0 5455 7 1 2 30165 29571
0 5456 5 1 1 5455
0 5457 7 1 2 5454 5456
0 5458 5 1 1 5457
0 5459 7 1 2 26145 5458
0 5460 5 1 1 5459
0 5461 7 1 2 5445 5460
0 5462 5 1 1 5461
0 5463 7 1 2 5462 32980
0 5464 5 1 1 5463
0 5465 7 1 2 32757 33195
0 5466 5 1 1 5465
0 5467 7 2 2 29826 32819
0 5468 5 1 1 33352
0 5469 7 1 2 22707 33353
0 5470 5 1 1 5469
0 5471 7 1 2 5466 5470
0 5472 5 1 1 5471
0 5473 7 1 2 31441 5472
0 5474 5 1 1 5473
0 5475 7 13 2 24673 22800
0 5476 7 3 2 23400 33354
0 5477 7 1 2 33367 30717
0 5478 5 1 1 5477
0 5479 7 9 2 22801 25356
0 5480 7 1 2 33370 30718
0 5481 5 1 1 5480
0 5482 7 1 2 32827 5481
0 5483 5 1 1 5482
0 5484 7 1 2 22708 5483
0 5485 5 1 1 5484
0 5486 7 1 2 5478 5485
0 5487 5 2 1 5486
0 5488 7 4 2 23108 25971
0 5489 7 1 2 33381 30760
0 5490 7 1 2 33379 5489
0 5491 5 1 1 5490
0 5492 7 1 2 5474 5491
0 5493 5 1 1 5492
0 5494 7 1 2 29137 5493
0 5495 5 1 1 5494
0 5496 7 2 2 26236 29827
0 5497 7 4 2 25357 23621
0 5498 7 1 2 31703 33387
0 5499 7 1 2 33385 5498
0 5500 7 1 2 33081 5499
0 5501 5 1 1 5500
0 5502 7 1 2 5495 5501
0 5503 5 1 1 5502
0 5504 7 1 2 24179 5503
0 5505 5 1 1 5504
0 5506 7 1 2 5464 5505
0 5507 5 1 1 5506
0 5508 7 1 2 22588 5507
0 5509 5 1 1 5508
0 5510 7 1 2 33371 30669
0 5511 5 1 1 5510
0 5512 7 1 2 32828 5511
0 5513 5 1 1 5512
0 5514 7 1 2 22709 5513
0 5515 5 1 1 5514
0 5516 7 1 2 33368 30670
0 5517 5 1 1 5516
0 5518 7 1 2 5515 5517
0 5519 5 1 1 5518
0 5520 7 1 2 31442 5519
0 5521 5 1 1 5520
0 5522 7 1 2 26714 33380
0 5523 5 1 1 5522
0 5524 7 1 2 5521 5523
0 5525 5 1 1 5524
0 5526 7 1 2 25287 5525
0 5527 5 1 1 5526
0 5528 7 1 2 148 3257
0 5529 5 1 1 5528
0 5530 7 1 2 27691 32970
0 5531 7 1 2 5529 5530
0 5532 5 1 1 5531
0 5533 7 1 2 5527 5532
0 5534 5 1 1 5533
0 5535 7 1 2 30192 33286
0 5536 7 1 2 5534 5535
0 5537 5 1 1 5536
0 5538 7 1 2 5509 5537
0 5539 5 1 1 5538
0 5540 7 1 2 27203 5539
0 5541 5 1 1 5540
0 5542 7 1 2 32751 33284
0 5543 5 1 1 5542
0 5544 7 1 2 32769 33270
0 5545 5 1 1 5544
0 5546 7 1 2 25767 32981
0 5547 7 1 2 33156 5546
0 5548 5 1 1 5547
0 5549 7 1 2 5545 5548
0 5550 5 1 1 5549
0 5551 7 1 2 31658 5550
0 5552 5 1 1 5551
0 5553 7 1 2 32773 33171
0 5554 5 1 1 5553
0 5555 7 2 2 25768 31704
0 5556 7 1 2 32971 33391
0 5557 5 1 1 5556
0 5558 7 1 2 4687 5557
0 5559 5 1 1 5558
0 5560 7 1 2 31443 5559
0 5561 5 1 1 5560
0 5562 7 5 2 23784 26237
0 5563 7 1 2 33393 26409
0 5564 7 1 2 32770 5563
0 5565 5 1 1 5564
0 5566 7 1 2 5561 5565
0 5567 5 1 1 5566
0 5568 7 1 2 24180 5567
0 5569 5 1 1 5568
0 5570 7 1 2 5554 5569
0 5571 5 1 1 5570
0 5572 7 1 2 31629 28202
0 5573 7 1 2 5571 5572
0 5574 5 1 1 5573
0 5575 7 1 2 5552 5574
0 5576 5 1 1 5575
0 5577 7 1 2 32575 5576
0 5578 5 1 1 5577
0 5579 7 1 2 5543 5578
0 5580 7 1 2 5541 5579
0 5581 7 1 2 5433 5580
0 5582 5 1 1 5581
0 5583 7 1 2 32721 5582
0 5584 5 1 1 5583
0 5585 7 1 2 5431 5584
0 5586 7 1 2 5291 5585
0 5587 7 1 2 5046 5586
0 5588 5 1 1 5587
0 5589 7 1 2 25675 5588
0 5590 5 1 1 5589
0 5591 7 1 2 32064 5590
0 5592 5 1 1 5591
0 5593 7 9 2 24340 25107
0 5594 5 6 1 33398
0 5595 7 1 2 23568 33407
0 5596 7 1 2 5592 5595
0 5597 7 1 2 4483 5596
0 5598 5 1 1 5597
0 5599 7 14 2 25518 24262
0 5600 5 4 1 33413
0 5601 7 2 2 22710 30817
0 5602 5 1 1 33431
0 5603 7 1 2 25972 30756
0 5604 5 1 1 5603
0 5605 7 1 2 5602 5604
0 5606 5 1 1 5605
0 5607 7 1 2 33414 5606
0 5608 5 1 1 5607
0 5609 7 2 2 26063 29815
0 5610 7 4 2 26943 33433
0 5611 7 1 2 24674 23526
0 5612 7 1 2 33435 5611
0 5613 5 1 1 5612
0 5614 7 1 2 5608 5613
0 5615 5 1 1 5614
0 5616 7 1 2 23338 5615
0 5617 5 1 1 5616
0 5618 7 2 2 26064 29183
0 5619 7 1 2 25288 30684
0 5620 7 8 2 23527 25973
0 5621 7 11 2 25044 25519
0 5622 5 1 1 33449
0 5623 7 1 2 33441 33450
0 5624 7 1 2 5619 5623
0 5625 7 1 2 33439 5624
0 5626 5 1 1 5625
0 5627 7 1 2 5617 5626
0 5628 5 1 1 5627
0 5629 7 1 2 29416 5628
0 5630 5 1 1 5629
0 5631 7 4 2 24091 29274
0 5632 7 1 2 25204 28757
0 5633 7 1 2 33460 5632
0 5634 7 3 2 25676 31113
0 5635 7 7 2 25484 25520
0 5636 5 1 1 33467
0 5637 7 2 2 25045 33468
0 5638 7 1 2 33464 33474
0 5639 7 1 2 5633 5638
0 5640 5 1 1 5639
0 5641 7 1 2 5630 5640
0 5642 5 1 1 5641
0 5643 7 1 2 24953 5642
0 5644 5 1 1 5643
0 5645 7 8 2 25521 26238
0 5646 5 1 1 33476
0 5647 7 1 2 27499 5646
0 5648 5 5 1 5647
0 5649 7 1 2 27521 26944
0 5650 7 3 2 33484 5649
0 5651 7 2 2 24675 30629
0 5652 7 1 2 29417 33492
0 5653 7 1 2 33489 5652
0 5654 5 1 1 5653
0 5655 7 1 2 5644 5654
0 5656 5 1 1 5655
0 5657 7 1 2 22589 5656
0 5658 5 1 1 5657
0 5659 7 8 2 23528 23682
0 5660 7 3 2 23251 33494
0 5661 7 5 2 29755 30464
0 5662 7 1 2 33502 33505
0 5663 5 2 1 5662
0 5664 7 6 2 31114 29951
0 5665 7 1 2 33512 30020
0 5666 5 1 1 5665
0 5667 7 1 2 33510 5666
0 5668 5 2 1 5667
0 5669 7 1 2 23339 33518
0 5670 5 1 1 5669
0 5671 7 1 2 30818 30802
0 5672 5 1 1 5671
0 5673 7 1 2 5670 5672
0 5674 5 1 1 5673
0 5675 7 6 2 33415 27800
0 5676 5 1 1 33520
0 5677 7 1 2 27455 33521
0 5678 7 1 2 5674 5677
0 5679 5 1 1 5678
0 5680 7 1 2 5658 5679
0 5681 5 1 1 5680
0 5682 7 1 2 25769 5681
0 5683 5 1 1 5682
0 5684 7 4 2 23529 25880
0 5685 7 4 2 26146 30330
0 5686 7 3 2 33526 33530
0 5687 7 1 2 25205 33534
0 5688 5 1 1 5687
0 5689 7 3 2 23909 29890
0 5690 7 2 2 24181 33537
0 5691 7 1 2 30738 33540
0 5692 5 2 1 5691
0 5693 7 1 2 5688 33542
0 5694 5 1 1 5693
0 5695 7 2 2 28127 5694
0 5696 5 1 1 33544
0 5697 7 18 2 24954 25522
0 5698 5 15 1 33546
0 5699 7 6 2 24263 33547
0 5700 7 1 2 31698 29474
0 5701 7 1 2 33579 5700
0 5702 7 1 2 33545 5701
0 5703 5 1 1 5702
0 5704 7 1 2 5683 5703
0 5705 5 1 1 5704
0 5706 7 1 2 24432 5705
0 5707 5 1 1 5706
0 5708 7 1 2 30819 29469
0 5709 5 1 1 5708
0 5710 7 1 2 23109 33511
0 5711 5 1 1 5710
0 5712 7 1 2 28128 33519
0 5713 7 1 2 5711 5712
0 5714 5 1 1 5713
0 5715 7 1 2 5709 5714
0 5716 5 1 1 5715
0 5717 7 1 2 23785 5716
0 5718 5 1 1 5717
0 5719 7 3 2 25206 23530
0 5720 7 3 2 25046 33585
0 5721 7 1 2 33588 33506
0 5722 5 1 1 5721
0 5723 7 1 2 33543 5722
0 5724 5 1 1 5723
0 5725 7 1 2 28129 31600
0 5726 7 1 2 5724 5725
0 5727 5 1 1 5726
0 5728 7 1 2 5718 5727
0 5729 5 1 1 5728
0 5730 7 3 2 22416 22711
0 5731 7 1 2 33591 33580
0 5732 7 1 2 5729 5731
0 5733 5 1 1 5732
0 5734 7 1 2 5707 5733
0 5735 5 1 1 5734
0 5736 7 1 2 23159 5735
0 5737 5 1 1 5736
0 5738 7 2 2 25677 33416
0 5739 7 1 2 23786 33535
0 5740 5 1 1 5739
0 5741 7 3 2 32188 29974
0 5742 5 1 1 33596
0 5743 7 1 2 5740 5742
0 5744 5 6 1 5743
0 5745 7 1 2 22417 33599
0 5746 5 2 1 5745
0 5747 7 1 2 27928 33605
0 5748 5 1 1 5747
0 5749 7 3 2 28700 30999
0 5750 5 1 1 33607
0 5751 7 1 2 28218 5750
0 5752 5 1 1 5751
0 5753 7 1 2 28130 5752
0 5754 7 1 2 5748 5753
0 5755 5 1 1 5754
0 5756 7 2 2 22590 30820
0 5757 5 2 1 33610
0 5758 7 1 2 32338 3267
0 5759 5 6 1 5758
0 5760 7 1 2 28357 33614
0 5761 7 1 2 33611 5760
0 5762 5 1 1 5761
0 5763 7 1 2 5755 5762
0 5764 5 1 1 5763
0 5765 7 2 2 33594 5764
0 5766 7 4 2 24955 25108
0 5767 7 4 2 22712 25047
0 5768 7 1 2 33622 33626
0 5769 7 1 2 33620 5768
0 5770 5 1 1 5769
0 5771 7 1 2 5737 5770
0 5772 5 1 1 5771
0 5773 7 1 2 22307 5772
0 5774 5 1 1 5773
0 5775 7 12 2 24341 23160
0 5776 5 1 1 33630
0 5777 7 3 2 22713 33631
0 5778 7 1 2 27801 33642
0 5779 7 1 2 33621 5778
0 5780 5 1 1 5779
0 5781 7 1 2 5774 5780
0 5782 5 1 1 5781
0 5783 7 1 2 24856 5782
0 5784 5 1 1 5783
0 5785 7 6 2 22418 25770
0 5786 7 14 2 23161 23683
0 5787 5 4 1 33651
0 5788 7 18 2 25109 25678
0 5789 5 1 1 33669
0 5790 7 2 2 25048 33670
0 5791 5 1 1 33687
0 5792 7 1 2 33665 5791
0 5793 5 6 1 5792
0 5794 7 1 2 33645 33689
0 5795 5 1 1 5794
0 5796 7 3 2 23162 23787
0 5797 5 1 1 33695
0 5798 7 9 2 24433 25049
0 5799 7 2 2 33696 33698
0 5800 5 1 1 33707
0 5801 7 1 2 25679 33708
0 5802 5 1 1 5801
0 5803 7 1 2 5795 5802
0 5804 5 1 1 5803
0 5805 7 1 2 22308 5804
0 5806 5 1 1 5805
0 5807 7 4 2 23163 25680
0 5808 7 5 2 24342 33709
0 5809 5 1 1 33713
0 5810 7 9 2 25050 25771
0 5811 7 4 2 33714 33718
0 5812 7 2 2 22419 33727
0 5813 5 1 1 33731
0 5814 7 1 2 5806 5813
0 5815 5 1 1 5814
0 5816 7 1 2 33432 5815
0 5817 5 1 1 5816
0 5818 7 1 2 23164 25485
0 5819 7 1 2 30237 5818
0 5820 7 8 2 23684 28701
0 5821 7 3 2 22309 30692
0 5822 7 1 2 33733 33741
0 5823 7 1 2 5819 5822
0 5824 5 1 1 5823
0 5825 7 1 2 5817 5824
0 5826 5 1 1 5825
0 5827 7 1 2 33417 5826
0 5828 5 1 1 5827
0 5829 7 3 2 23165 33742
0 5830 7 1 2 25772 33495
0 5831 7 1 2 33436 5830
0 5832 7 1 2 33744 5831
0 5833 5 1 1 5832
0 5834 7 1 2 5828 5833
0 5835 5 1 1 5834
0 5836 7 1 2 24956 5835
0 5837 5 1 1 5836
0 5838 7 2 2 23531 31601
0 5839 7 2 2 33490 33747
0 5840 7 1 2 33745 33749
0 5841 5 1 1 5840
0 5842 7 1 2 5837 5841
0 5843 5 1 1 5842
0 5844 7 1 2 24857 5843
0 5845 5 1 1 5844
0 5846 7 2 2 29869 29275
0 5847 7 2 2 33734 33751
0 5848 7 2 2 25523 33753
0 5849 7 5 2 24957 23166
0 5850 7 2 2 29055 33757
0 5851 7 1 2 33743 33762
0 5852 7 1 2 33755 5851
0 5853 5 1 1 5852
0 5854 7 1 2 5845 5853
0 5855 5 1 1 5854
0 5856 7 1 2 29220 5855
0 5857 5 1 1 5856
0 5858 7 2 2 33758 32405
0 5859 7 6 2 23532 25524
0 5860 5 1 1 33766
0 5861 7 1 2 26945 31033
0 5862 7 1 2 33767 5861
0 5863 7 6 2 26065 29276
0 5864 5 1 1 33772
0 5865 7 8 2 22310 24434
0 5866 7 2 2 31602 33778
0 5867 7 1 2 33773 33786
0 5868 7 1 2 5862 5867
0 5869 7 1 2 33764 5868
0 5870 5 1 1 5869
0 5871 7 1 2 5857 5870
0 5872 7 1 2 5784 5871
0 5873 5 1 1 5872
0 5874 7 1 2 28722 5873
0 5875 5 1 1 5874
0 5876 7 6 2 25422 25881
0 5877 7 3 2 29891 33788
0 5878 5 1 1 33794
0 5879 7 1 2 23458 30809
0 5880 5 1 1 5879
0 5881 7 1 2 5878 5880
0 5882 5 10 1 5881
0 5883 7 1 2 22802 33797
0 5884 5 2 1 5883
0 5885 7 2 2 28004 30812
0 5886 5 1 1 33809
0 5887 7 1 2 33807 5886
0 5888 5 1 1 5887
0 5889 7 1 2 29157 5888
0 5890 5 1 1 5889
0 5891 7 8 2 23459 30331
0 5892 7 5 2 22803 25051
0 5893 7 1 2 33811 33819
0 5894 7 1 2 30229 5893
0 5895 5 1 1 5894
0 5896 7 1 2 5890 5895
0 5897 5 1 1 5896
0 5898 7 1 2 25773 5897
0 5899 5 1 1 5898
0 5900 7 4 2 30332 26339
0 5901 7 2 2 33824 33235
0 5902 7 1 2 33223 33828
0 5903 5 1 1 5902
0 5904 7 1 2 5899 5903
0 5905 5 1 1 5904
0 5906 7 1 2 32078 5905
0 5907 5 1 1 5906
0 5908 7 2 2 24746 29459
0 5909 7 6 2 22591 29756
0 5910 7 3 2 25423 25774
0 5911 7 2 2 33832 33838
0 5912 7 1 2 33830 33841
0 5913 5 1 1 5912
0 5914 7 8 2 24560 23910
0 5915 5 5 1 33843
0 5916 7 1 2 31267 33851
0 5917 5 2 1 5916
0 5918 7 5 2 23460 24001
0 5919 7 1 2 28451 33858
0 5920 7 1 2 31694 5919
0 5921 7 1 2 33856 5920
0 5922 5 1 1 5921
0 5923 7 1 2 5913 5922
0 5924 5 1 1 5923
0 5925 7 1 2 22420 5924
0 5926 5 1 1 5925
0 5927 7 1 2 30532 31917
0 5928 7 1 2 33842 5927
0 5929 5 1 1 5928
0 5930 7 1 2 5926 5929
0 5931 5 1 1 5930
0 5932 7 1 2 32238 5931
0 5933 5 1 1 5932
0 5934 7 1 2 33789 27393
0 5935 7 1 2 33251 5934
0 5936 5 1 1 5935
0 5937 7 1 2 3986 5936
0 5938 5 1 1 5937
0 5939 7 1 2 25775 5938
0 5940 7 1 2 33320 5939
0 5941 5 1 1 5940
0 5942 7 5 2 28037 28399
0 5943 7 2 2 28055 33863
0 5944 7 1 2 28850 27235
0 5945 7 1 2 33868 5944
0 5946 5 1 1 5945
0 5947 7 1 2 5941 5946
0 5948 7 1 2 5933 5947
0 5949 5 1 1 5948
0 5950 7 1 2 26066 5949
0 5951 5 1 1 5950
0 5952 7 1 2 5907 5951
0 5953 5 1 1 5952
0 5954 7 1 2 23685 5953
0 5955 5 1 1 5954
0 5956 7 2 2 23788 31671
0 5957 7 2 2 30693 32309
0 5958 5 1 1 33872
0 5959 7 1 2 24435 32847
0 5960 5 1 1 5959
0 5961 7 1 2 5958 5960
0 5962 5 4 1 5961
0 5963 7 1 2 33870 33874
0 5964 5 1 1 5963
0 5965 7 3 2 28439 31387
0 5966 5 1 1 33878
0 5967 7 1 2 31950 28281
0 5968 5 1 1 5967
0 5969 7 1 2 33852 31311
0 5970 5 1 1 5969
0 5971 7 1 2 24436 5970
0 5972 7 1 2 5968 5971
0 5973 5 1 1 5972
0 5974 7 1 2 5966 5973
0 5975 5 1 1 5974
0 5976 7 1 2 32239 5975
0 5977 5 1 1 5976
0 5978 7 3 2 28017 31853
0 5979 7 3 2 31630 31453
0 5980 5 1 1 33884
0 5981 7 1 2 33881 33885
0 5982 5 1 1 5981
0 5983 7 1 2 5977 5982
0 5984 7 1 2 5964 5983
0 5985 5 1 1 5984
0 5986 7 1 2 24002 5985
0 5987 5 1 1 5986
0 5988 7 1 2 24437 33236
0 5989 5 2 1 5988
0 5990 7 1 2 27929 33887
0 5991 5 1 1 5990
0 5992 7 3 2 24561 30433
0 5993 5 2 1 33889
0 5994 7 1 2 27955 33892
0 5995 5 1 1 5994
0 5996 7 3 2 5991 5995
0 5997 7 1 2 27143 32079
0 5998 7 1 2 33894 5997
0 5999 5 1 1 5998
0 6000 7 1 2 5987 5999
0 6001 5 1 1 6000
0 6002 7 6 2 26067 26340
0 6003 7 1 2 33897 29475
0 6004 7 1 2 6001 6003
0 6005 5 1 1 6004
0 6006 7 1 2 5955 6005
0 6007 5 1 1 6006
0 6008 7 1 2 23167 6007
0 6009 5 1 1 6008
0 6010 7 1 2 25681 32468
0 6011 7 2 2 32434 6010
0 6012 7 2 2 22804 25110
0 6013 7 1 2 25052 33905
0 6014 7 1 2 33903 6013
0 6015 5 1 1 6014
0 6016 7 1 2 6009 6015
0 6017 5 1 1 6016
0 6018 7 1 2 22311 6017
0 6019 5 1 1 6018
0 6020 7 8 2 25424 24092
0 6021 5 2 1 33907
0 6022 7 3 2 22805 33908
0 6023 5 1 1 33917
0 6024 7 6 2 24747 32451
0 6025 5 2 1 33920
0 6026 7 1 2 6023 33926
0 6027 5 12 1 6026
0 6028 7 8 2 23686 32045
0 6029 7 1 2 32863 33940
0 6030 5 1 1 6029
0 6031 7 2 2 25111 23340
0 6032 5 2 1 33948
0 6033 7 1 2 28319 33950
0 6034 5 2 1 6033
0 6035 7 14 2 23168 25207
0 6036 5 1 1 33954
0 6037 7 1 2 618 6036
0 6038 5 2 1 6037
0 6039 7 3 2 33952 33968
0 6040 7 1 2 22421 33970
0 6041 5 1 1 6040
0 6042 7 19 2 24438 23169
0 6043 5 1 1 33973
0 6044 7 1 2 29221 33974
0 6045 5 1 1 6044
0 6046 7 1 2 6041 6045
0 6047 5 6 1 6046
0 6048 7 1 2 29476 33992
0 6049 5 1 1 6048
0 6050 7 3 2 22592 23170
0 6051 7 2 2 22422 33998
0 6052 7 1 2 30609 34001
0 6053 5 1 1 6052
0 6054 7 1 2 6049 6053
0 6055 5 1 1 6054
0 6056 7 1 2 22312 6055
0 6057 5 1 1 6056
0 6058 7 13 2 24343 22423
0 6059 7 2 2 31971 34003
0 6060 7 1 2 28358 33710
0 6061 7 1 2 34016 6060
0 6062 5 1 1 6061
0 6063 7 1 2 6057 6062
0 6064 5 2 1 6063
0 6065 7 1 2 32503 34018
0 6066 5 1 1 6065
0 6067 7 1 2 22714 27048
0 6068 5 1 1 6067
0 6069 7 1 2 4206 6068
0 6070 5 19 1 6069
0 6071 7 2 2 28131 34020
0 6072 5 1 1 34039
0 6073 7 4 2 23911 27956
0 6074 7 4 2 32046 34041
0 6075 7 1 2 34045 29477
0 6076 7 1 2 34040 6075
0 6077 5 1 1 6076
0 6078 7 1 2 6066 6077
0 6079 5 1 1 6078
0 6080 7 1 2 23789 6079
0 6081 5 1 1 6080
0 6082 7 1 2 28203 33690
0 6083 5 1 1 6082
0 6084 7 1 2 33975 29463
0 6085 5 1 1 6084
0 6086 7 1 2 6083 6085
0 6087 5 1 1 6086
0 6088 7 1 2 22313 6087
0 6089 5 1 1 6088
0 6090 7 2 2 25053 33715
0 6091 5 1 1 34049
0 6092 7 1 2 28204 34050
0 6093 5 1 1 6092
0 6094 7 1 2 6089 6093
0 6095 5 7 1 6094
0 6096 7 1 2 32495 34051
0 6097 5 1 1 6096
0 6098 7 2 2 6081 6097
0 6099 7 1 2 6030 34058
0 6100 5 1 1 6099
0 6101 7 1 2 33928 6100
0 6102 5 1 1 6101
0 6103 7 1 2 33632 33820
0 6104 7 1 2 33904 6103
0 6105 5 1 1 6104
0 6106 7 1 2 6102 6105
0 6107 7 1 2 6019 6106
0 6108 5 1 1 6107
0 6109 7 1 2 27491 6108
0 6110 5 1 1 6109
0 6111 7 11 2 23031 23569
0 6112 5 13 1 34060
0 6113 7 9 2 26239 34071
0 6114 5 1 1 34084
0 6115 7 5 2 25974 32469
0 6116 7 1 2 33237 34052
0 6117 5 1 1 6116
0 6118 7 3 2 28305 29478
0 6119 7 1 2 34046 34098
0 6120 5 1 1 6119
0 6121 7 1 2 6117 6120
0 6122 5 1 1 6121
0 6123 7 2 2 23790 6122
0 6124 5 1 1 34101
0 6125 7 1 2 25054 27020
0 6126 5 1 1 6125
0 6127 7 1 2 27291 6126
0 6128 5 3 1 6127
0 6129 7 1 2 22593 34103
0 6130 5 1 1 6129
0 6131 7 1 2 25055 33124
0 6132 5 1 1 6131
0 6133 7 1 2 6130 6132
0 6134 5 2 1 6133
0 6135 7 1 2 27957 34106
0 6136 5 1 1 6135
0 6137 7 1 2 28056 31148
0 6138 5 1 1 6137
0 6139 7 1 2 6136 6138
0 6140 5 2 1 6139
0 6141 7 1 2 32047 31603
0 6142 7 1 2 34108 6141
0 6143 5 1 1 6142
0 6144 7 1 2 6124 6143
0 6145 5 1 1 6144
0 6146 7 1 2 34093 6145
0 6147 5 1 1 6146
0 6148 7 2 2 25776 30062
0 6149 7 1 2 33795 32048
0 6150 7 1 2 34110 6149
0 6151 5 1 1 6150
0 6152 7 1 2 6147 6151
0 6153 5 1 1 6152
0 6154 7 1 2 22806 6153
0 6155 5 1 1 6154
0 6156 7 1 2 32049 33810
0 6157 7 1 2 34111 6156
0 6158 5 1 1 6157
0 6159 7 1 2 6155 6158
0 6160 5 1 1 6159
0 6161 7 1 2 32080 6160
0 6162 5 1 1 6161
0 6163 7 4 2 25358 31188
0 6164 5 1 1 34112
0 6165 7 1 2 2949 6164
0 6166 5 1 1 6165
0 6167 7 4 2 3696 6166
0 6168 7 1 2 22424 34116
0 6169 5 1 1 6168
0 6170 7 2 2 22715 28400
0 6171 7 1 2 28337 34120
0 6172 5 1 1 6171
0 6173 7 1 2 6169 6172
0 6174 5 6 1 6173
0 6175 7 1 2 34122 34104
0 6176 5 1 1 6175
0 6177 7 1 2 24562 30976
0 6178 5 2 1 6177
0 6179 7 1 2 2871 34128
0 6180 5 18 1 6179
0 6181 7 1 2 25056 31153
0 6182 5 1 1 6181
0 6183 7 1 2 31150 6182
0 6184 5 1 1 6183
0 6185 7 1 2 22425 6184
0 6186 5 1 1 6185
0 6187 7 1 2 31833 33699
0 6188 5 1 1 6187
0 6189 7 1 2 6186 6188
0 6190 5 1 1 6189
0 6191 7 1 2 34130 6190
0 6192 5 1 1 6191
0 6193 7 1 2 6176 6192
0 6194 5 1 1 6193
0 6195 7 5 2 25777 25975
0 6196 7 1 2 33941 34148
0 6197 7 1 2 6194 6196
0 6198 5 1 1 6197
0 6199 7 1 2 34059 6198
0 6200 5 1 1 6199
0 6201 7 1 2 33929 6200
0 6202 5 1 1 6201
0 6203 7 7 2 22807 24003
0 6204 7 3 2 32470 34153
0 6205 7 8 2 27386 27844
0 6206 7 6 2 23171 23252
0 6207 7 5 2 34171 34004
0 6208 5 1 1 34177
0 6209 7 1 2 34163 34178
0 6210 5 2 1 6209
0 6211 7 3 2 25289 27958
0 6212 7 2 2 34131 34184
0 6213 5 1 1 34187
0 6214 7 5 2 24439 31189
0 6215 7 2 2 23253 32226
0 6216 7 1 2 34189 34194
0 6217 5 1 1 6216
0 6218 7 1 2 6213 6217
0 6219 5 1 1 6218
0 6220 7 1 2 23172 6219
0 6221 5 1 1 6220
0 6222 7 5 2 25112 23254
0 6223 7 2 2 22426 34196
0 6224 5 1 1 34201
0 6225 7 1 2 34164 34202
0 6226 5 1 1 6225
0 6227 7 1 2 6221 6226
0 6228 5 1 1 6227
0 6229 7 1 2 22314 6228
0 6230 5 1 1 6229
0 6231 7 1 2 34182 6230
0 6232 5 1 1 6231
0 6233 7 1 2 28440 29479
0 6234 7 1 2 6232 6233
0 6235 5 1 1 6234
0 6236 7 6 2 22427 25359
0 6237 5 1 1 34203
0 6238 7 1 2 594 6237
0 6239 5 1 1 6238
0 6240 7 1 2 30859 29377
0 6241 7 2 2 6239 6240
0 6242 7 2 2 23173 31308
0 6243 5 1 1 34211
0 6244 7 2 2 25113 33275
0 6245 5 1 1 34213
0 6246 7 1 2 6243 6245
0 6247 5 2 1 6246
0 6248 7 1 2 29480 34215
0 6249 5 1 1 6248
0 6250 7 3 2 34172 31604
0 6251 5 1 1 34217
0 6252 7 1 2 6249 6251
0 6253 5 2 1 6252
0 6254 7 1 2 27284 34220
0 6255 5 1 1 6254
0 6256 7 6 2 25057 23791
0 6257 7 3 2 25882 34222
0 6258 7 5 2 23174 25290
0 6259 7 1 2 29397 34231
0 6260 7 1 2 34228 6259
0 6261 5 1 1 6260
0 6262 7 1 2 6255 6261
0 6263 5 1 1 6262
0 6264 7 1 2 22315 6263
0 6265 5 1 1 6264
0 6266 7 2 2 27285 31718
0 6267 7 2 2 33633 30533
0 6268 7 1 2 34236 34238
0 6269 5 1 1 6268
0 6270 7 1 2 6265 6269
0 6271 5 1 1 6270
0 6272 7 1 2 34209 6271
0 6273 5 1 1 6272
0 6274 7 3 2 27254 34053
0 6275 7 1 2 34132 34240
0 6276 5 2 1 6275
0 6277 7 3 2 22428 33716
0 6278 7 1 2 27845 31881
0 6279 7 2 2 34245 6278
0 6280 5 1 1 34248
0 6281 7 5 2 23175 25360
0 6282 7 3 2 34190 34250
0 6283 5 1 1 34255
0 6284 7 1 2 34256 29481
0 6285 5 1 1 6284
0 6286 7 1 2 33691 32412
0 6287 5 1 1 6286
0 6288 7 1 2 6285 6287
0 6289 5 1 1 6288
0 6290 7 1 2 22316 6289
0 6291 5 1 1 6290
0 6292 7 1 2 6280 6291
0 6293 5 1 1 6292
0 6294 7 4 2 27292 311
0 6295 5 1 1 34258
0 6296 7 1 2 703 31312
0 6297 7 2 2 6295 6296
0 6298 7 1 2 6293 34262
0 6299 5 1 1 6298
0 6300 7 1 2 34243 6299
0 6301 7 1 2 6273 6300
0 6302 7 1 2 6235 6301
0 6303 5 1 1 6302
0 6304 7 1 2 34160 6303
0 6305 5 1 1 6304
0 6306 7 1 2 6202 6305
0 6307 7 1 2 6162 6306
0 6308 5 1 1 6307
0 6309 7 1 2 34085 6308
0 6310 5 1 1 6309
0 6311 7 1 2 6110 6310
0 6312 5 1 1 6311
0 6313 7 1 2 24858 6312
0 6314 5 1 1 6313
0 6315 7 3 2 25525 31751
0 6316 5 2 1 34264
0 6317 7 8 2 24093 28973
0 6318 7 8 2 22716 25114
0 6319 7 2 2 23401 28702
0 6320 7 1 2 34277 34285
0 6321 5 1 1 6320
0 6322 7 4 2 23176 28441
0 6323 7 1 2 31009 34287
0 6324 5 1 1 6323
0 6325 7 1 2 6321 6324
0 6326 5 1 1 6325
0 6327 7 1 2 22317 6326
0 6328 5 1 1 6327
0 6329 7 1 2 33643 34286
0 6330 5 1 1 6329
0 6331 7 1 2 6328 6330
0 6332 5 1 1 6331
0 6333 7 1 2 30312 6332
0 6334 5 1 1 6333
0 6335 7 6 2 25361 25883
0 6336 7 2 2 24676 34291
0 6337 7 1 2 6043 29378
0 6338 5 1 1 6337
0 6339 7 2 2 33953 6338
0 6340 7 1 2 22318 34299
0 6341 5 1 1 6340
0 6342 7 1 2 23177 28231
0 6343 7 1 2 34005 6342
0 6344 5 1 1 6343
0 6345 7 1 2 6341 6344
0 6346 5 1 1 6345
0 6347 7 1 2 28285 6346
0 6348 5 1 1 6347
0 6349 7 1 2 29134 1403
0 6350 5 4 1 6349
0 6351 7 10 2 22319 25115
0 6352 5 1 1 34305
0 6353 7 3 2 5776 6352
0 6354 5 22 1 34315
0 6355 7 1 2 33276 34318
0 6356 5 1 1 6355
0 6357 7 1 2 22320 34212
0 6358 5 1 1 6357
0 6359 7 1 2 6356 6358
0 6360 5 2 1 6359
0 6361 7 1 2 34301 34340
0 6362 5 1 1 6361
0 6363 7 1 2 6348 6362
0 6364 5 1 1 6363
0 6365 7 1 2 34297 6364
0 6366 5 1 1 6365
0 6367 7 1 2 6334 6366
0 6368 5 1 1 6367
0 6369 7 1 2 29482 6368
0 6370 5 1 1 6369
0 6371 7 2 2 28132 34054
0 6372 7 2 2 27204 31010
0 6373 5 1 1 34344
0 6374 7 6 2 23402 23792
0 6375 7 2 2 25884 34346
0 6376 7 1 2 22717 34352
0 6377 5 1 1 6376
0 6378 7 1 2 6373 6377
0 6379 5 2 1 6378
0 6380 7 1 2 34342 34354
0 6381 5 1 1 6380
0 6382 7 1 2 31264 30110
0 6383 7 1 2 34195 6382
0 6384 7 1 2 33746 6383
0 6385 5 1 1 6384
0 6386 7 1 2 6381 6385
0 6387 7 1 2 6370 6386
0 6388 5 1 1 6387
0 6389 7 1 2 25976 6388
0 6390 5 1 1 6389
0 6391 7 1 2 33976 34099
0 6392 5 1 1 6391
0 6393 7 1 2 32672 33692
0 6394 5 1 1 6393
0 6395 7 1 2 6392 6394
0 6396 5 1 1 6395
0 6397 7 1 2 22321 6396
0 6398 5 1 1 6397
0 6399 7 4 2 23341 31972
0 6400 7 1 2 34006 33711
0 6401 7 1 2 34356 6400
0 6402 5 1 1 6401
0 6403 7 1 2 6398 6402
0 6404 5 1 1 6403
0 6405 7 1 2 28286 6404
0 6406 5 1 1 6405
0 6407 7 1 2 22322 34221
0 6408 5 1 1 6407
0 6409 7 1 2 31719 34239
0 6410 5 1 1 6409
0 6411 7 1 2 6408 6410
0 6412 5 1 1 6411
0 6413 7 1 2 34302 6412
0 6414 5 1 1 6413
0 6415 7 1 2 6406 6414
0 6416 5 1 1 6415
0 6417 7 1 2 28631 532
0 6418 5 1 1 6417
0 6419 7 1 2 6416 6418
0 6420 5 1 1 6419
0 6421 7 1 2 22429 34216
0 6422 5 1 1 6421
0 6423 7 1 2 33977 28287
0 6424 5 1 1 6423
0 6425 7 1 2 6422 6424
0 6426 5 1 1 6425
0 6427 7 1 2 29483 6426
0 6428 5 1 1 6427
0 6429 7 1 2 22430 34218
0 6430 5 1 1 6429
0 6431 7 1 2 6428 6430
0 6432 5 1 1 6431
0 6433 7 1 2 22323 6432
0 6434 5 1 1 6433
0 6435 7 1 2 23255 33732
0 6436 5 1 1 6435
0 6437 7 1 2 6434 6436
0 6438 5 1 1 6437
0 6439 7 1 2 31115 32144
0 6440 7 1 2 6438 6439
0 6441 5 1 1 6440
0 6442 7 1 2 6420 6441
0 6443 7 1 2 6390 6442
0 6444 5 1 1 6443
0 6445 7 1 2 34269 6444
0 6446 5 1 1 6445
0 6447 7 1 2 27959 28839
0 6448 5 1 1 6447
0 6449 7 4 2 22431 32344
0 6450 7 2 2 31321 31131
0 6451 7 1 2 34360 34364
0 6452 5 1 1 6451
0 6453 7 1 2 6448 6452
0 6454 5 1 1 6453
0 6455 7 1 2 31545 6454
0 6456 5 1 1 6455
0 6457 7 1 2 31631 32325
0 6458 7 1 2 33864 6457
0 6459 5 1 1 6458
0 6460 7 1 2 6456 6459
0 6461 5 1 1 6460
0 6462 7 1 2 30166 33942
0 6463 7 1 2 6461 6462
0 6464 5 1 1 6463
0 6465 7 1 2 3056 31296
0 6466 5 1 1 6465
0 6467 7 2 2 28813 29374
0 6468 7 1 2 25116 34366
0 6469 5 1 1 6468
0 6470 7 1 2 23178 28785
0 6471 7 1 2 32350 6470
0 6472 5 1 1 6471
0 6473 7 1 2 6469 6472
0 6474 5 1 1 6473
0 6475 7 1 2 22324 6474
0 6476 5 1 1 6475
0 6477 7 4 2 24344 29375
0 6478 7 3 2 23179 23461
0 6479 7 2 2 22808 34372
0 6480 7 1 2 23403 34375
0 6481 7 1 2 34368 6480
0 6482 5 1 1 6481
0 6483 7 1 2 6476 6482
0 6484 5 1 1 6483
0 6485 7 1 2 6466 6484
0 6486 5 1 1 6485
0 6487 7 1 2 5797 33951
0 6488 5 2 1 6487
0 6489 7 2 2 22325 34377
0 6490 7 1 2 34379 34259
0 6491 5 1 1 6490
0 6492 7 1 2 25778 27434
0 6493 7 1 2 33634 6492
0 6494 5 1 1 6493
0 6495 7 1 2 6491 6494
0 6496 5 1 1 6495
0 6497 7 2 2 24563 28814
0 6498 5 1 1 34381
0 6499 7 1 2 3247 6498
0 6500 5 2 1 6499
0 6501 7 1 2 27960 34383
0 6502 7 1 2 6496 6501
0 6503 5 1 1 6502
0 6504 7 1 2 6486 6503
0 6505 5 1 1 6504
0 6506 7 1 2 29484 6505
0 6507 5 1 1 6506
0 6508 7 1 2 34241 34384
0 6509 5 1 1 6508
0 6510 7 1 2 33693 34367
0 6511 5 1 1 6510
0 6512 7 2 2 26888 29485
0 6513 7 1 2 29603 34251
0 6514 7 1 2 34385 6513
0 6515 5 1 1 6514
0 6516 7 1 2 6511 6515
0 6517 5 1 1 6516
0 6518 7 1 2 22326 6517
0 6519 5 1 1 6518
0 6520 7 8 2 25058 23180
0 6521 7 2 2 34007 34387
0 6522 7 1 2 22594 25682
0 6523 7 1 2 28815 6522
0 6524 7 1 2 34395 6523
0 6525 5 1 1 6524
0 6526 7 1 2 6519 6525
0 6527 5 1 1 6526
0 6528 7 1 2 34263 6527
0 6529 5 1 1 6528
0 6530 7 2 2 28786 34361
0 6531 5 1 1 34397
0 6532 7 1 2 28816 28338
0 6533 5 1 1 6532
0 6534 7 1 2 6531 6533
0 6535 5 1 1 6534
0 6536 7 1 2 22327 27286
0 6537 7 1 2 34219 6536
0 6538 5 1 1 6537
0 6539 7 1 2 27308 29486
0 6540 7 1 2 34341 6539
0 6541 5 1 1 6540
0 6542 7 1 2 6538 6541
0 6543 5 1 1 6542
0 6544 7 1 2 6535 6543
0 6545 5 1 1 6544
0 6546 7 1 2 6529 6545
0 6547 7 1 2 6509 6546
0 6548 7 1 2 6507 6547
0 6549 7 1 2 6464 6548
0 6550 5 1 1 6549
0 6551 7 1 2 32576 6550
0 6552 5 1 1 6551
0 6553 7 5 2 23912 27863
0 6554 7 2 2 23687 33999
0 6555 7 2 2 34399 34404
0 6556 5 1 1 34406
0 6557 7 1 2 33666 5789
0 6558 5 3 1 6557
0 6559 7 1 2 30224 34408
0 6560 5 1 1 6559
0 6561 7 2 2 23913 33671
0 6562 7 1 2 28232 34411
0 6563 5 1 1 6562
0 6564 7 1 2 6560 6563
0 6565 5 1 1 6564
0 6566 7 1 2 25779 6565
0 6567 5 1 1 6566
0 6568 7 1 2 34288 29450
0 6569 5 1 1 6568
0 6570 7 1 2 6567 6569
0 6571 5 1 1 6570
0 6572 7 1 2 25059 6571
0 6573 5 1 1 6572
0 6574 7 1 2 6556 6573
0 6575 5 1 1 6574
0 6576 7 1 2 28767 6575
0 6577 5 1 1 6576
0 6578 7 6 2 24564 23181
0 6579 7 1 2 34413 27859
0 6580 5 1 1 6579
0 6581 7 1 2 22595 34378
0 6582 7 1 2 34260 6581
0 6583 5 1 1 6582
0 6584 7 1 2 6580 6583
0 6585 5 1 1 6584
0 6586 7 9 2 25683 24004
0 6587 7 1 2 34419 33345
0 6588 7 1 2 6585 6587
0 6589 5 1 1 6588
0 6590 7 1 2 6577 6589
0 6591 5 1 1 6590
0 6592 7 1 2 22328 6591
0 6593 5 1 1 6592
0 6594 7 1 2 33728 33130
0 6595 5 1 1 6594
0 6596 7 1 2 6593 6595
0 6597 5 1 1 6596
0 6598 7 1 2 27961 6597
0 6599 5 1 1 6598
0 6600 7 3 2 25977 27456
0 6601 5 2 1 34428
0 6602 7 2 2 24005 31034
0 6603 5 1 1 34433
0 6604 7 1 2 34431 6603
0 6605 5 5 1 6604
0 6606 7 1 2 34435 34242
0 6607 5 1 1 6606
0 6608 7 2 2 28205 32050
0 6609 7 2 2 23688 34440
0 6610 7 2 2 27144 27846
0 6611 5 1 1 34444
0 6612 7 1 2 34442 34445
0 6613 5 1 1 6612
0 6614 7 5 2 24440 33955
0 6615 5 1 1 34446
0 6616 7 1 2 6224 6615
0 6617 5 7 1 6616
0 6618 7 1 2 22329 34451
0 6619 5 1 1 6618
0 6620 7 1 2 6619 6208
0 6621 5 11 1 6620
0 6622 7 2 2 27169 31190
0 6623 5 1 1 34469
0 6624 7 1 2 6611 6623
0 6625 5 1 1 6624
0 6626 7 1 2 29487 6625
0 6627 7 1 2 34458 6626
0 6628 5 1 1 6627
0 6629 7 1 2 6613 6628
0 6630 5 1 1 6629
0 6631 7 1 2 27309 6630
0 6632 5 1 1 6631
0 6633 7 2 2 23342 34443
0 6634 7 5 2 24006 27205
0 6635 7 1 2 31191 34473
0 6636 7 1 2 34471 6635
0 6637 5 1 1 6636
0 6638 7 1 2 6632 6637
0 6639 7 1 2 6607 6638
0 6640 7 1 2 6599 6639
0 6641 5 1 1 6640
0 6642 7 1 2 28723 6641
0 6643 5 1 1 6642
0 6644 7 1 2 6552 6643
0 6645 5 1 1 6644
0 6646 7 1 2 26068 6645
0 6647 5 1 1 6646
0 6648 7 1 2 6446 6647
0 6649 5 1 1 6648
0 6650 7 1 2 34265 6649
0 6651 5 1 1 6650
0 6652 7 1 2 6314 6651
0 6653 5 1 1 6652
0 6654 7 1 2 28639 6653
0 6655 5 1 1 6654
0 6656 7 3 2 26538 30111
0 6657 7 1 2 22596 33956
0 6658 7 1 2 34478 6657
0 6659 5 1 1 6658
0 6660 7 4 2 24565 25684
0 6661 7 3 2 23914 34481
0 6662 7 3 2 25117 23533
0 6663 7 1 2 31201 34488
0 6664 7 1 2 34485 6663
0 6665 5 1 1 6664
0 6666 7 1 2 6659 6665
0 6667 5 1 1 6666
0 6668 7 1 2 22432 6667
0 6669 5 1 1 6668
0 6670 7 1 2 27895 34479
0 6671 5 1 1 6670
0 6672 7 3 2 24859 25685
0 6673 7 2 2 30904 34491
0 6674 7 2 2 24566 34494
0 6675 7 1 2 25208 34496
0 6676 5 1 1 6675
0 6677 7 1 2 6671 6676
0 6678 5 1 1 6677
0 6679 7 1 2 33978 6678
0 6680 5 1 1 6679
0 6681 7 1 2 6669 6680
0 6682 5 1 1 6681
0 6683 7 1 2 22330 6682
0 6684 5 1 1 6683
0 6685 7 1 2 34179 34497
0 6686 5 1 1 6685
0 6687 7 1 2 6684 6686
0 6688 5 1 1 6687
0 6689 7 1 2 32240 6688
0 6690 5 1 1 6689
0 6691 7 1 2 34414 34480
0 6692 5 1 1 6691
0 6693 7 4 2 22597 25118
0 6694 7 4 2 30132 34498
0 6695 7 1 2 26386 34502
0 6696 5 1 1 6695
0 6697 7 1 2 6692 6696
0 6698 5 1 1 6697
0 6699 7 1 2 22331 6698
0 6700 5 1 1 6699
0 6701 7 4 2 24345 34000
0 6702 7 1 2 34506 34495
0 6703 5 1 1 6702
0 6704 7 1 2 6700 6703
0 6705 5 1 1 6704
0 6706 7 1 2 33321 6705
0 6707 5 1 1 6706
0 6708 7 7 2 25362 28018
0 6709 7 2 2 29398 34510
0 6710 5 1 1 34517
0 6711 7 3 2 22332 28339
0 6712 7 2 2 24860 23182
0 6713 7 1 2 30905 34522
0 6714 7 1 2 34519 6713
0 6715 7 1 2 34518 6714
0 6716 5 1 1 6715
0 6717 7 1 2 6707 6716
0 6718 7 1 2 6690 6717
0 6719 5 1 1 6718
0 6720 7 1 2 29952 6719
0 6721 5 1 1 6720
0 6722 7 2 2 32081 30313
0 6723 7 5 2 23689 30771
0 6724 7 1 2 30356 32051
0 6725 7 1 2 34526 6724
0 6726 7 1 2 34524 6725
0 6727 5 1 1 6726
0 6728 7 1 2 6721 6727
0 6729 5 1 1 6728
0 6730 7 1 2 25780 6729
0 6731 5 1 1 6730
0 6732 7 1 2 34459 33238
0 6733 5 1 1 6732
0 6734 7 3 2 28306 32052
0 6735 7 1 2 34042 34531
0 6736 5 1 1 6735
0 6737 7 1 2 6733 6736
0 6738 5 1 1 6737
0 6739 7 2 2 32082 29056
0 6740 7 2 2 30465 31505
0 6741 7 1 2 34534 34536
0 6742 7 1 2 6738 6741
0 6743 5 1 1 6742
0 6744 7 1 2 6731 6743
0 6745 5 1 1 6744
0 6746 7 1 2 25978 6745
0 6747 5 1 1 6746
0 6748 7 1 2 22598 27255
0 6749 5 1 1 6748
0 6750 7 5 2 24567 27206
0 6751 7 1 2 23343 34538
0 6752 5 1 1 6751
0 6753 7 1 2 6749 6752
0 6754 5 2 1 6753
0 6755 7 1 2 34460 34543
0 6756 5 1 1 6755
0 6757 7 3 2 23793 32053
0 6758 7 2 2 27962 30895
0 6759 5 1 1 34548
0 6760 7 1 2 34545 34549
0 6761 5 1 1 6760
0 6762 7 1 2 6756 6761
0 6763 5 1 1 6762
0 6764 7 3 2 24094 32083
0 6765 7 1 2 29652 34420
0 6766 7 1 2 34550 6765
0 6767 7 1 2 6763 6766
0 6768 5 1 1 6767
0 6769 7 1 2 6747 6768
0 6770 5 1 1 6769
0 6771 7 1 2 25060 6770
0 6772 5 1 1 6771
0 6773 7 1 2 30821 28376
0 6774 5 1 1 6773
0 6775 7 1 2 33600 28378
0 6776 5 1 1 6775
0 6777 7 1 2 6774 6776
0 6778 5 1 1 6777
0 6779 7 3 2 22928 32084
0 6780 7 1 2 33943 34553
0 6781 7 1 2 6778 6780
0 6782 5 1 1 6781
0 6783 7 1 2 6772 6782
0 6784 5 1 1 6783
0 6785 7 1 2 34086 6784
0 6786 5 1 1 6785
0 6787 7 9 2 25209 30133
0 6788 7 6 2 24568 25061
0 6789 7 1 2 34556 34565
0 6790 5 1 1 6789
0 6791 7 1 2 6790 31956
0 6792 5 1 1 6791
0 6793 7 1 2 24441 6792
0 6794 5 1 1 6793
0 6795 7 1 2 6794 3901
0 6796 5 1 1 6795
0 6797 7 1 2 32241 6796
0 6798 5 1 1 6797
0 6799 7 1 2 33322 31928
0 6800 5 1 1 6799
0 6801 7 3 2 25062 28670
0 6802 7 1 2 28939 31035
0 6803 7 1 2 30134 6802
0 6804 7 1 2 34571 6803
0 6805 5 1 1 6804
0 6806 7 1 2 6800 6805
0 6807 7 1 2 6798 6806
0 6808 5 1 1 6807
0 6809 7 1 2 31172 6808
0 6810 5 1 1 6809
0 6811 7 3 2 23690 32085
0 6812 7 1 2 30285 34574
0 6813 7 1 2 34109 6812
0 6814 5 1 1 6813
0 6815 7 1 2 6810 6814
0 6816 5 1 1 6815
0 6817 7 1 2 25781 6816
0 6818 5 1 1 6817
0 6819 7 1 2 33239 29682
0 6820 5 1 1 6819
0 6821 7 1 2 34043 34100
0 6822 5 1 1 6821
0 6823 7 1 2 6820 6822
0 6824 5 1 1 6823
0 6825 7 5 2 23794 26069
0 6826 7 6 2 26147 34577
0 6827 7 1 2 34554 34582
0 6828 7 1 2 6824 6827
0 6829 5 1 1 6828
0 6830 7 1 2 6818 6829
0 6831 5 1 1 6830
0 6832 7 1 2 23534 6831
0 6833 5 1 1 6832
0 6834 7 1 2 29514 33735
0 6835 7 1 2 30262 6834
0 6836 7 1 2 32913 6835
0 6837 5 1 1 6836
0 6838 7 1 2 6833 6837
0 6839 5 1 1 6838
0 6840 7 1 2 23032 6839
0 6841 5 1 1 6840
0 6842 7 5 2 22929 33548
0 6843 5 1 1 34588
0 6844 7 1 2 34589 26483
0 6845 7 1 2 33736 6844
0 6846 7 1 2 31182 6845
0 6847 7 1 2 32914 6846
0 6848 5 1 1 6847
0 6849 7 1 2 6841 6848
0 6850 5 1 1 6849
0 6851 7 1 2 25979 6850
0 6852 5 1 1 6851
0 6853 7 2 2 24442 33277
0 6854 5 1 1 34593
0 6855 7 1 2 6854 3428
0 6856 5 1 1 6855
0 6857 7 3 2 23691 6856
0 6858 5 1 1 34595
0 6859 7 1 2 33700 31520
0 6860 5 1 1 6859
0 6861 7 1 2 6858 6860
0 6862 5 1 1 6861
0 6863 7 1 2 27435 6862
0 6864 5 1 1 6863
0 6865 7 1 2 25686 27226
0 6866 7 1 2 31896 6865
0 6867 5 1 1 6866
0 6868 7 1 2 6864 6867
0 6869 5 1 1 6868
0 6870 7 1 2 22599 6869
0 6871 5 1 1 6870
0 6872 7 3 2 30574 33701
0 6873 7 1 2 34598 34237
0 6874 5 1 1 6873
0 6875 7 3 2 31506 29460
0 6876 5 1 1 34601
0 6877 7 1 2 31617 6876
0 6878 5 1 1 6877
0 6879 7 1 2 22433 6878
0 6880 5 1 1 6879
0 6881 7 5 2 25687 33702
0 6882 7 1 2 28257 34604
0 6883 5 1 1 6882
0 6884 7 1 2 6880 6883
0 6885 5 1 1 6884
0 6886 7 1 2 30896 6885
0 6887 5 1 1 6886
0 6888 7 1 2 6874 6887
0 6889 7 1 2 6871 6888
0 6890 5 1 1 6889
0 6891 7 6 2 24007 32086
0 6892 5 1 1 34609
0 6893 7 3 2 24182 34610
0 6894 7 1 2 26395 31216
0 6895 7 1 2 34615 6894
0 6896 7 1 2 6890 6895
0 6897 5 1 1 6896
0 6898 7 1 2 6852 6897
0 6899 5 1 1 6898
0 6900 7 1 2 32054 6899
0 6901 5 1 1 6900
0 6902 7 5 2 25210 23404
0 6903 7 2 2 25782 31173
0 6904 7 1 2 34618 34623
0 6905 5 1 1 6904
0 6906 7 1 2 34578 29337
0 6907 7 1 2 31132 6906
0 6908 5 1 1 6907
0 6909 7 1 2 6905 6908
0 6910 5 1 1 6909
0 6911 7 1 2 22718 6910
0 6912 5 1 1 6911
0 6913 7 1 2 30834 27468
0 6914 7 1 2 34583 6913
0 6915 5 1 1 6914
0 6916 7 1 2 6912 6915
0 6917 5 1 1 6916
0 6918 7 1 2 23344 6917
0 6919 5 1 1 6918
0 6920 7 1 2 29953 28074
0 6921 7 1 2 32778 30026
0 6922 7 1 2 6920 6921
0 6923 5 1 1 6922
0 6924 7 1 2 6919 6923
0 6925 5 1 1 6924
0 6926 7 1 2 23915 6925
0 6927 5 1 1 6926
0 6928 7 2 2 32087 27469
0 6929 7 1 2 27021 34584
0 6930 7 1 2 34625 6929
0 6931 5 1 1 6930
0 6932 7 1 2 6927 6931
0 6933 5 1 1 6932
0 6934 7 1 2 33442 6933
0 6935 5 1 1 6934
0 6936 7 6 2 28563 29515
0 6937 5 1 1 34627
0 6938 7 1 2 27256 34628
0 6939 7 1 2 34626 6938
0 6940 5 1 1 6939
0 6941 7 1 2 6935 6940
0 6942 5 1 1 6941
0 6943 7 1 2 22600 6942
0 6944 5 1 1 6943
0 6945 7 3 2 24861 27207
0 6946 7 1 2 29954 27752
0 6947 7 1 2 34633 6946
0 6948 5 1 1 6947
0 6949 7 1 2 27436 26862
0 6950 7 1 2 34585 6949
0 6951 5 1 1 6950
0 6952 7 1 2 6948 6951
0 6953 5 1 1 6952
0 6954 7 1 2 22719 6953
0 6955 5 1 1 6954
0 6956 7 1 2 30286 34353
0 6957 5 1 1 6956
0 6958 7 1 2 27176 34624
0 6959 5 1 1 6958
0 6960 7 1 2 6957 6959
0 6961 5 1 1 6960
0 6962 7 1 2 28874 6961
0 6963 5 1 1 6962
0 6964 7 1 2 6955 6963
0 6965 5 1 1 6964
0 6966 7 1 2 33443 6965
0 6967 5 1 1 6966
0 6968 7 1 2 22930 29516
0 6969 7 1 2 34400 6968
0 6970 7 1 2 34616 6969
0 6971 5 1 1 6970
0 6972 7 1 2 6967 6971
0 6973 5 1 1 6972
0 6974 7 1 2 30643 6973
0 6975 5 1 1 6974
0 6976 7 1 2 6944 6975
0 6977 5 1 1 6976
0 6978 7 1 2 22434 6977
0 6979 5 1 1 6978
0 6980 7 1 2 25783 26387
0 6981 7 1 2 32695 6980
0 6982 7 1 2 32432 6981
0 6983 5 1 1 6982
0 6984 7 1 2 6979 6983
0 6985 5 1 1 6984
0 6986 7 6 2 25688 34319
0 6987 7 1 2 34636 26530
0 6988 7 1 2 6985 6987
0 6989 5 1 1 6988
0 6990 7 1 2 6901 6989
0 6991 5 1 1 6990
0 6992 7 1 2 24264 6991
0 6993 5 1 1 6992
0 6994 7 1 2 6786 6993
0 6995 5 1 1 6994
0 6996 7 1 2 28974 6995
0 6997 5 1 1 6996
0 6998 7 1 2 30047 33491
0 6999 5 1 1 6998
0 7000 7 1 2 24569 31056
0 7001 7 1 2 33507 7000
0 7002 5 1 1 7001
0 7003 7 1 2 33612 7002
0 7004 5 1 1 7003
0 7005 7 1 2 24677 7004
0 7006 5 1 1 7005
0 7007 7 1 2 29517 30490
0 7008 7 1 2 34429 7007
0 7009 5 1 1 7008
0 7010 7 1 2 7006 7009
0 7011 5 1 1 7010
0 7012 7 1 2 33418 7011
0 7013 5 1 1 7012
0 7014 7 1 2 30048 33437
0 7015 5 1 1 7014
0 7016 7 1 2 7013 7015
0 7017 5 1 1 7016
0 7018 7 1 2 24958 7017
0 7019 5 1 1 7018
0 7020 7 1 2 6999 7019
0 7021 5 1 1 7020
0 7022 7 1 2 31605 7021
0 7023 5 1 1 7022
0 7024 7 4 2 30705 28564
0 7025 7 3 2 34642 31647
0 7026 7 2 2 24570 32211
0 7027 7 1 2 33475 34649
0 7028 7 1 2 34646 7027
0 7029 5 1 1 7028
0 7030 7 1 2 7023 7029
0 7031 5 1 1 7030
0 7032 7 1 2 22435 7031
0 7033 5 1 1 7032
0 7034 7 1 2 31659 31000
0 7035 5 1 1 7034
0 7036 7 1 2 33613 7035
0 7037 5 3 1 7036
0 7038 7 1 2 23795 34651
0 7039 5 1 1 7038
0 7040 7 1 2 24571 33597
0 7041 5 1 1 7040
0 7042 7 1 2 7039 7041
0 7043 5 1 1 7042
0 7044 7 3 2 24443 27802
0 7045 5 1 1 34654
0 7046 7 1 2 33419 29745
0 7047 7 1 2 34655 7046
0 7048 7 1 2 7043 7047
0 7049 5 1 1 7048
0 7050 7 1 2 7033 7049
0 7051 5 1 1 7050
0 7052 7 1 2 23183 7051
0 7053 5 1 1 7052
0 7054 7 1 2 33420 31720
0 7055 7 2 2 34652 7054
0 7056 7 3 2 25119 27803
0 7057 5 1 1 34659
0 7058 7 1 2 30694 34660
0 7059 7 1 2 34657 7058
0 7060 5 1 1 7059
0 7061 7 1 2 7053 7060
0 7062 5 1 1 7061
0 7063 7 1 2 22333 7062
0 7064 5 1 1 7063
0 7065 7 1 2 32212 34396
0 7066 7 1 2 34658 7065
0 7067 5 1 1 7066
0 7068 7 1 2 7064 7067
0 7069 5 1 1 7068
0 7070 7 1 2 24862 7069
0 7071 5 1 1 7070
0 7072 7 1 2 22334 22436
0 7073 7 1 2 27457 7072
0 7074 7 1 2 33763 7073
0 7075 7 1 2 33756 7074
0 7076 5 1 1 7075
0 7077 7 1 2 7071 7076
0 7078 5 1 1 7077
0 7079 7 1 2 33036 7078
0 7080 5 1 1 7079
0 7081 7 4 2 28442 34421
0 7082 7 1 2 29975 34662
0 7083 5 1 1 7082
0 7084 7 2 2 31798 30747
0 7085 5 1 1 34666
0 7086 7 1 2 7083 7085
0 7087 5 2 1 7086
0 7088 7 1 2 22601 34668
0 7089 5 1 1 7088
0 7090 7 1 2 24572 31507
0 7091 7 1 2 30822 7090
0 7092 5 1 1 7091
0 7093 7 1 2 7089 7092
0 7094 5 1 1 7093
0 7095 7 1 2 33346 7094
0 7096 5 1 1 7095
0 7097 7 1 2 33833 31606
0 7098 7 1 2 30006 7097
0 7099 5 1 1 7098
0 7100 7 1 2 7096 7099
0 7101 5 1 1 7100
0 7102 7 1 2 33421 7101
0 7103 5 1 1 7102
0 7104 7 1 2 27847 33748
0 7105 7 1 2 33438 7104
0 7106 5 1 1 7105
0 7107 7 1 2 7103 7106
0 7108 5 1 1 7107
0 7109 7 1 2 24959 7108
0 7110 5 1 1 7109
0 7111 7 1 2 27848 33750
0 7112 5 1 1 7111
0 7113 7 1 2 7110 7112
0 7114 5 1 1 7113
0 7115 7 1 2 23184 7114
0 7116 5 1 1 7115
0 7117 7 5 2 22602 25784
0 7118 7 10 2 25689 25885
0 7119 7 1 2 33768 34675
0 7120 7 1 2 34670 7119
0 7121 7 3 2 30333 29184
0 7122 7 6 2 25063 25120
0 7123 7 2 2 34688 32213
0 7124 7 1 2 34685 34694
0 7125 7 1 2 7120 7124
0 7126 5 1 1 7125
0 7127 7 1 2 7116 7126
0 7128 5 1 1 7127
0 7129 7 1 2 24863 7128
0 7130 5 1 1 7129
0 7131 7 2 2 23185 23535
0 7132 7 1 2 27849 34696
0 7133 7 1 2 34590 7132
0 7134 7 1 2 33754 7133
0 7135 5 1 1 7134
0 7136 7 1 2 7130 7135
0 7137 5 1 1 7136
0 7138 7 1 2 22335 7137
0 7139 5 1 1 7138
0 7140 7 3 2 33635 34492
0 7141 5 1 1 34698
0 7142 7 1 2 33527 31036
0 7143 7 1 2 34699 7142
0 7144 7 2 2 33549 33719
0 7145 7 1 2 34686 34701
0 7146 7 1 2 7143 7145
0 7147 5 1 1 7146
0 7148 7 1 2 7139 7147
0 7149 5 1 1 7148
0 7150 7 1 2 27963 7149
0 7151 5 1 1 7150
0 7152 7 1 2 22603 33601
0 7153 5 1 1 7152
0 7154 7 3 2 24573 25785
0 7155 7 1 2 30823 34703
0 7156 5 1 1 7155
0 7157 7 1 2 7153 7156
0 7158 5 1 1 7157
0 7159 7 2 2 24960 30027
0 7160 7 1 2 33422 34706
0 7161 7 1 2 34055 7160
0 7162 7 1 2 7158 7161
0 7163 5 1 1 7162
0 7164 7 1 2 7151 7163
0 7165 5 1 1 7164
0 7166 7 1 2 28822 7165
0 7167 5 1 1 7166
0 7168 7 4 2 33423 32389
0 7169 7 2 2 28975 34708
0 7170 7 1 2 26384 811
0 7171 5 3 1 7170
0 7172 7 1 2 27408 34714
0 7173 5 1 1 7172
0 7174 7 1 2 28632 7173
0 7175 5 1 1 7174
0 7176 7 1 2 33652 7175
0 7177 5 1 1 7176
0 7178 7 2 2 22720 34689
0 7179 7 1 2 25690 26980
0 7180 7 1 2 34717 7179
0 7181 5 1 1 7180
0 7182 7 1 2 7177 7181
0 7183 5 1 1 7182
0 7184 7 1 2 22336 7183
0 7185 5 1 1 7184
0 7186 7 2 2 27032 33627
0 7187 7 1 2 23916 33717
0 7188 7 1 2 34719 7187
0 7189 5 1 1 7188
0 7190 7 1 2 7185 7189
0 7191 5 1 1 7190
0 7192 7 1 2 29158 7191
0 7193 5 1 1 7192
0 7194 7 1 2 22337 34409
0 7195 5 1 1 7194
0 7196 7 1 2 5809 7195
0 7197 5 1 1 7196
0 7198 7 1 2 7197 30230
0 7199 5 1 1 7198
0 7200 7 3 2 23186 33779
0 7201 7 1 2 28307 34721
0 7202 7 1 2 34557 7201
0 7203 5 1 1 7202
0 7204 7 1 2 7199 7203
0 7205 5 1 1 7204
0 7206 7 1 2 34720 7205
0 7207 5 1 1 7206
0 7208 7 1 2 7193 7207
0 7209 5 1 1 7208
0 7210 7 1 2 25786 7209
0 7211 5 1 1 7210
0 7212 7 1 2 30992 34102
0 7213 5 1 1 7212
0 7214 7 1 2 34056 34544
0 7215 5 1 1 7214
0 7216 7 1 2 27864 34507
0 7217 5 1 1 7216
0 7218 7 1 2 28090 31268
0 7219 7 1 2 34380 7218
0 7220 5 1 1 7219
0 7221 7 1 2 7217 7220
0 7222 5 1 1 7221
0 7223 7 1 2 27964 7222
0 7224 5 1 1 7223
0 7225 7 1 2 34461 28326
0 7226 5 1 1 7225
0 7227 7 1 2 7224 7226
0 7228 5 1 1 7227
0 7229 7 1 2 25886 7228
0 7230 5 1 1 7229
0 7231 7 2 2 23796 28133
0 7232 7 1 2 34047 34724
0 7233 5 1 1 7232
0 7234 7 1 2 7230 7233
0 7235 5 1 1 7234
0 7236 7 1 2 29488 7235
0 7237 5 1 1 7236
0 7238 7 1 2 7215 7237
0 7239 5 2 1 7238
0 7240 7 1 2 34021 34726
0 7241 5 1 1 7240
0 7242 7 1 2 7213 7241
0 7243 7 1 2 7211 7242
0 7244 5 1 1 7243
0 7245 7 1 2 34712 7244
0 7246 5 1 1 7245
0 7247 7 2 2 24574 30779
0 7248 5 1 1 34728
0 7249 7 2 2 25887 27871
0 7250 5 1 1 34730
0 7251 7 1 2 7248 7250
0 7252 5 1 1 7251
0 7253 7 1 2 33979 7252
0 7254 5 1 1 7253
0 7255 7 3 2 25121 25888
0 7256 5 1 1 34732
0 7257 7 1 2 33853 7256
0 7258 5 1 1 7257
0 7259 7 1 2 22437 33969
0 7260 7 1 2 7258 7259
0 7261 5 1 1 7260
0 7262 7 1 2 7254 7261
0 7263 5 2 1 7262
0 7264 7 1 2 29489 34735
0 7265 5 1 1 7264
0 7266 7 1 2 34002 30120
0 7267 5 1 1 7266
0 7268 7 1 2 7265 7267
0 7269 5 1 1 7268
0 7270 7 1 2 22338 7269
0 7271 5 1 1 7270
0 7272 7 1 2 34173 34676
0 7273 7 1 2 34017 7272
0 7274 5 1 1 7273
0 7275 7 1 2 7271 7274
0 7276 5 1 1 7275
0 7277 7 1 2 28026 7276
0 7278 5 1 1 7277
0 7279 7 5 2 24678 25211
0 7280 5 1 1 34737
0 7281 7 2 2 26889 34232
0 7282 7 1 2 34738 34742
0 7283 5 1 1 7282
0 7284 7 1 2 34278 31696
0 7285 5 1 1 7284
0 7286 7 1 2 7283 7285
0 7287 5 2 1 7286
0 7288 7 1 2 22438 34744
0 7289 5 1 1 7288
0 7290 7 1 2 31584 33980
0 7291 5 1 1 7290
0 7292 7 1 2 7289 7291
0 7293 5 1 1 7292
0 7294 7 1 2 22339 7293
0 7295 5 1 1 7294
0 7296 7 1 2 27888 34180
0 7297 5 1 1 7296
0 7298 7 1 2 7295 7297
0 7299 5 1 1 7298
0 7300 7 1 2 31672 29490
0 7301 7 1 2 7299 7300
0 7302 5 1 1 7301
0 7303 7 1 2 31660 27279
0 7304 7 1 2 34472 7303
0 7305 5 1 1 7304
0 7306 7 1 2 7302 7305
0 7307 7 1 2 7278 7306
0 7308 5 1 1 7307
0 7309 7 1 2 23797 7308
0 7310 5 1 1 7309
0 7311 7 1 2 22439 31587
0 7312 5 1 1 7311
0 7313 7 1 2 7312 620
0 7314 5 2 1 7313
0 7315 7 2 2 27208 34746
0 7316 7 1 2 34748 33944
0 7317 5 1 1 7316
0 7318 7 1 2 7310 7317
0 7319 5 1 1 7318
0 7320 7 1 2 27074 7319
0 7321 5 1 1 7320
0 7322 7 4 2 26375 30135
0 7323 7 2 2 24575 34197
0 7324 7 1 2 34750 34754
0 7325 5 1 1 7324
0 7326 7 2 2 31854 33653
0 7327 7 1 2 33834 34756
0 7328 5 1 1 7327
0 7329 7 1 2 7325 7328
0 7330 5 1 1 7329
0 7331 7 1 2 22440 7330
0 7332 5 1 1 7331
0 7333 7 2 2 31116 34482
0 7334 7 1 2 34758 34619
0 7335 5 1 1 7334
0 7336 7 1 2 22604 31133
0 7337 7 1 2 29773 7336
0 7338 5 1 1 7337
0 7339 7 1 2 7335 7338
0 7340 5 1 1 7339
0 7341 7 1 2 33981 7340
0 7342 5 1 1 7341
0 7343 7 1 2 7332 7342
0 7344 5 1 1 7343
0 7345 7 1 2 25064 7344
0 7346 5 1 1 7345
0 7347 7 1 2 26376 34405
0 7348 7 1 2 30200 7347
0 7349 5 1 1 7348
0 7350 7 1 2 7346 7349
0 7351 5 1 1 7350
0 7352 7 1 2 22340 7351
0 7353 5 1 1 7352
0 7354 7 2 2 24576 34388
0 7355 7 3 2 24346 28206
0 7356 7 1 2 34751 34762
0 7357 7 1 2 34760 7356
0 7358 5 1 1 7357
0 7359 7 1 2 7353 7358
0 7360 5 1 1 7359
0 7361 7 1 2 28027 7360
0 7362 5 1 1 7361
0 7363 7 1 2 34499 34752
0 7364 5 1 1 7363
0 7365 7 1 2 25363 34415
0 7366 7 1 2 29774 7365
0 7367 5 1 1 7366
0 7368 7 1 2 7364 7367
0 7369 5 1 1 7368
0 7370 7 1 2 22341 7369
0 7371 5 1 1 7370
0 7372 7 1 2 34508 34753
0 7373 5 1 1 7372
0 7374 7 1 2 7371 7373
0 7375 5 1 1 7374
0 7376 7 1 2 25065 7375
0 7377 5 1 1 7376
0 7378 7 3 2 22342 34416
0 7379 7 2 2 26946 30841
0 7380 7 1 2 34765 34768
0 7381 5 1 1 7380
0 7382 7 1 2 7377 7381
0 7383 5 1 1 7382
0 7384 7 1 2 31926 7383
0 7385 5 1 1 7384
0 7386 7 2 2 31354 31897
0 7387 7 1 2 33465 32341
0 7388 7 1 2 34770 7387
0 7389 5 1 1 7388
0 7390 7 1 2 29159 26992
0 7391 5 1 1 7390
0 7392 7 1 2 28134 31889
0 7393 5 1 1 7392
0 7394 7 1 2 7391 7393
0 7395 5 1 1 7394
0 7396 7 1 2 23692 27128
0 7397 7 1 2 7395 7396
0 7398 5 1 1 7397
0 7399 7 1 2 7389 7398
0 7400 5 1 1 7399
0 7401 7 1 2 32055 7400
0 7402 5 1 1 7401
0 7403 7 1 2 7385 7402
0 7404 7 1 2 7362 7403
0 7405 5 1 1 7404
0 7406 7 1 2 25787 7405
0 7407 5 1 1 7406
0 7408 7 1 2 27129 27188
0 7409 7 1 2 34343 7408
0 7410 5 1 1 7409
0 7411 7 1 2 27735 34019
0 7412 5 1 1 7411
0 7413 7 1 2 24008 27965
0 7414 7 2 2 28187 7413
0 7415 7 1 2 29491 34772
0 7416 5 1 1 7415
0 7417 7 2 2 25980 30610
0 7418 7 1 2 22441 27857
0 7419 7 1 2 34774 7418
0 7420 5 1 1 7419
0 7421 7 1 2 7416 7420
0 7422 5 1 1 7421
0 7423 7 1 2 27177 32056
0 7424 7 1 2 7422 7423
0 7425 5 1 1 7424
0 7426 7 1 2 7412 7425
0 7427 5 1 1 7426
0 7428 7 1 2 23798 7427
0 7429 5 1 1 7428
0 7430 7 1 2 7410 7429
0 7431 7 1 2 7407 7430
0 7432 7 1 2 7321 7431
0 7433 5 1 1 7432
0 7434 7 1 2 27500 6114
0 7435 5 4 1 7434
0 7436 7 1 2 22931 34776
0 7437 7 1 2 7433 7436
0 7438 5 1 1 7437
0 7439 7 1 2 7246 7438
0 7440 5 1 1 7439
0 7441 7 1 2 31467 7440
0 7442 5 1 1 7441
0 7443 7 1 2 30399 2700
0 7444 5 11 1 7443
0 7445 7 1 2 24679 28724
0 7446 5 1 1 7445
0 7447 7 2 2 30855 26890
0 7448 5 1 1 34791
0 7449 7 1 2 7446 7448
0 7450 5 4 1 7449
0 7451 7 1 2 34793 34727
0 7452 5 1 1 7451
0 7453 7 3 2 28803 27268
0 7454 7 2 2 25788 33240
0 7455 7 1 2 34320 34800
0 7456 5 1 1 7455
0 7457 7 1 2 28443 34532
0 7458 5 1 1 7457
0 7459 7 1 2 7456 7458
0 7460 5 1 1 7459
0 7461 7 1 2 29492 7460
0 7462 5 1 1 7461
0 7463 7 1 2 22343 34407
0 7464 5 1 1 7463
0 7465 7 1 2 7462 7464
0 7466 5 1 1 7465
0 7467 7 1 2 27966 7466
0 7468 5 1 1 7467
0 7469 7 1 2 1894 694
0 7470 5 1 1 7469
0 7471 7 1 2 923 7470
0 7472 7 1 2 34057 7471
0 7473 5 1 1 7472
0 7474 7 10 2 23917 31508
0 7475 7 1 2 34357 34802
0 7476 7 1 2 34462 7475
0 7477 5 1 1 7476
0 7478 7 1 2 7473 7477
0 7479 7 1 2 7468 7478
0 7480 5 1 1 7479
0 7481 7 1 2 34797 7480
0 7482 5 1 1 7481
0 7483 7 1 2 7452 7482
0 7484 5 1 1 7483
0 7485 7 1 2 34709 7484
0 7486 5 1 1 7485
0 7487 7 1 2 34113 33957
0 7488 5 1 1 7487
0 7489 7 3 2 22605 34198
0 7490 7 2 2 30977 34812
0 7491 5 1 1 34815
0 7492 7 1 2 7488 7491
0 7493 5 1 1 7492
0 7494 7 1 2 22442 7493
0 7495 5 1 1 7494
0 7496 7 1 2 34117 33982
0 7497 5 1 1 7496
0 7498 7 1 2 7495 7497
0 7499 5 4 1 7498
0 7500 7 1 2 34817 29493
0 7501 5 1 1 7500
0 7502 7 2 2 34174 30842
0 7503 7 1 2 34821 28459
0 7504 5 1 1 7503
0 7505 7 1 2 7501 7504
0 7506 5 1 1 7505
0 7507 7 1 2 22344 7506
0 7508 5 1 1 7507
0 7509 7 1 2 23256 34249
0 7510 5 1 1 7509
0 7511 7 1 2 7508 7510
0 7512 5 1 1 7511
0 7513 7 1 2 27310 7512
0 7514 5 1 1 7513
0 7515 7 1 2 25291 34133
0 7516 7 2 2 34048 7515
0 7517 5 1 1 34823
0 7518 7 1 2 34824 29494
0 7519 5 1 1 7518
0 7520 7 1 2 7514 7519
0 7521 5 1 1 7520
0 7522 7 1 2 23799 7521
0 7523 5 1 1 7522
0 7524 7 1 2 22345 33694
0 7525 5 1 1 7524
0 7526 7 1 2 6091 7525
0 7527 5 1 1 7526
0 7528 7 1 2 34123 7527
0 7529 5 1 1 7528
0 7530 7 3 2 22346 34566
0 7531 7 2 2 31855 31712
0 7532 7 1 2 34828 33712
0 7533 7 1 2 34825 7532
0 7534 5 1 1 7533
0 7535 7 1 2 7529 7534
0 7536 5 1 1 7535
0 7537 7 1 2 34401 7536
0 7538 5 1 1 7537
0 7539 7 1 2 34244 7538
0 7540 7 1 2 7523 7539
0 7541 5 1 1 7540
0 7542 7 2 2 22932 28976
0 7543 7 1 2 34777 34830
0 7544 7 1 2 7541 7543
0 7545 5 1 1 7544
0 7546 7 1 2 7486 7545
0 7547 5 1 1 7546
0 7548 7 1 2 34780 7547
0 7549 5 1 1 7548
0 7550 7 1 2 33615 34653
0 7551 5 1 1 7550
0 7552 7 1 2 33598 28057
0 7553 5 1 1 7552
0 7554 7 1 2 7551 7553
0 7555 5 1 1 7554
0 7556 7 2 2 33595 7555
0 7557 7 1 2 33865 34695
0 7558 5 1 1 7557
0 7559 7 2 2 31856 34233
0 7560 7 1 2 27355 27804
0 7561 7 1 2 34834 7560
0 7562 5 1 1 7561
0 7563 7 1 2 7558 7562
0 7564 5 1 1 7563
0 7565 7 1 2 34832 7564
0 7566 5 1 1 7565
0 7567 7 1 2 31673 32326
0 7568 5 2 1 7567
0 7569 7 2 2 25889 34567
0 7570 5 1 1 34838
0 7571 7 1 2 31640 7570
0 7572 5 1 1 7571
0 7573 7 1 2 31454 7572
0 7574 5 1 1 7573
0 7575 7 1 2 34836 7574
0 7576 5 1 1 7575
0 7577 7 2 2 29185 33769
0 7578 5 1 1 34840
0 7579 7 2 2 25981 32214
0 7580 7 1 2 34841 34842
0 7581 7 1 2 7576 7580
0 7582 5 1 1 7581
0 7583 7 1 2 25789 33528
0 7584 7 1 2 30066 7583
0 7585 5 1 1 7584
0 7586 7 2 2 26148 31809
0 7587 7 1 2 30208 34844
0 7588 5 1 1 7587
0 7589 7 1 2 7585 7588
0 7590 5 1 1 7589
0 7591 7 1 2 28851 34778
0 7592 7 1 2 7590 7591
0 7593 5 1 1 7592
0 7594 7 1 2 7582 7593
0 7595 5 1 1 7594
0 7596 7 1 2 26070 7595
0 7597 5 1 1 7596
0 7598 7 1 2 31904 34436
0 7599 5 1 1 7598
0 7600 7 1 2 31117 28064
0 7601 5 1 1 7600
0 7602 7 1 2 7599 7601
0 7603 5 1 1 7602
0 7604 7 1 2 25790 7603
0 7605 5 1 1 7604
0 7606 7 1 2 32802 31810
0 7607 5 1 1 7606
0 7608 7 1 2 7605 7607
0 7609 5 1 1 7608
0 7610 7 1 2 29976 33581
0 7611 7 1 2 7609 7610
0 7612 5 1 1 7611
0 7613 7 1 2 7597 7612
0 7614 5 1 1 7613
0 7615 7 1 2 23693 7614
0 7616 5 1 1 7615
0 7617 7 2 2 29032 33451
0 7618 7 1 2 34191 34846
0 7619 7 1 2 34647 7618
0 7620 5 1 1 7619
0 7621 7 1 2 7616 7620
0 7622 5 1 1 7621
0 7623 7 1 2 23187 33866
0 7624 7 1 2 7622 7623
0 7625 5 1 1 7624
0 7626 7 1 2 7566 7625
0 7627 5 1 1 7626
0 7628 7 1 2 22347 7627
0 7629 5 1 1 7628
0 7630 7 3 2 22809 24961
0 7631 7 2 2 25066 34848
0 7632 7 1 2 24680 33636
0 7633 7 1 2 28404 7632
0 7634 7 1 2 34851 7633
0 7635 7 1 2 34833 7634
0 7636 5 1 1 7635
0 7637 7 1 2 7629 7636
0 7638 5 1 1 7637
0 7639 7 1 2 24864 7638
0 7640 5 1 1 7639
0 7641 7 1 2 27771 33774
0 7642 7 1 2 28685 7641
0 7643 7 7 2 23536 28804
0 7644 7 8 2 25526 23694
0 7645 7 1 2 34860 33780
0 7646 7 1 2 34853 7645
0 7647 7 1 2 33765 7646
0 7648 7 1 2 7642 7647
0 7649 5 1 1 7648
0 7650 7 1 2 7640 7649
0 7651 7 1 2 7549 7650
0 7652 7 1 2 7442 7651
0 7653 7 1 2 7167 7652
0 7654 7 1 2 7080 7653
0 7655 7 1 2 6997 7654
0 7656 7 1 2 6655 7655
0 7657 7 1 2 5875 7656
0 7658 5 1 1 7657
0 7659 7 1 2 26435 7658
0 7660 5 1 1 7659
0 7661 7 4 2 23570 26240
0 7662 5 2 1 34868
0 7663 7 1 2 24962 34872
0 7664 5 1 1 7663
0 7665 7 1 2 33427 7664
0 7666 5 13 1 7665
0 7667 7 6 2 24865 34874
0 7668 5 1 1 34887
0 7669 7 1 2 7668 5676
0 7670 5 1 1 7669
0 7671 7 1 2 33930 7670
0 7672 5 1 1 7671
0 7673 7 2 2 26736 31217
0 7674 5 2 1 34893
0 7675 7 1 2 26891 34894
0 7676 5 1 1 7675
0 7677 7 1 2 7672 7676
0 7678 5 1 1 7677
0 7679 7 1 2 28640 7678
0 7680 5 1 1 7679
0 7681 7 1 2 22933 34875
0 7682 5 2 1 7681
0 7683 7 1 2 22934 5622
0 7684 5 5 1 7683
0 7685 7 1 2 26737 34899
0 7686 5 1 1 7685
0 7687 7 1 2 34897 7686
0 7688 5 1 1 7687
0 7689 7 2 2 25425 31468
0 7690 5 1 1 34904
0 7691 7 1 2 23462 29977
0 7692 5 1 1 7691
0 7693 7 1 2 7690 7692
0 7694 5 1 1 7693
0 7695 7 1 2 24748 7694
0 7696 5 1 1 7695
0 7697 7 1 2 27605 33918
0 7698 5 1 1 7697
0 7699 7 1 2 7696 7698
0 7700 5 1 1 7699
0 7701 7 1 2 7688 7700
0 7702 5 1 1 7701
0 7703 7 2 2 23537 32983
0 7704 5 1 1 34906
0 7705 7 1 2 25067 29287
0 7706 7 1 2 27567 7705
0 7707 7 2 2 7704 7706
0 7708 7 5 2 24866 25527
0 7709 5 1 1 34910
0 7710 7 1 2 34911 33931
0 7711 7 1 2 34908 7710
0 7712 5 1 1 7711
0 7713 7 1 2 7702 7712
0 7714 7 1 2 7680 7713
0 7715 5 1 1 7714
0 7716 7 1 2 26959 7715
0 7717 5 1 1 7716
0 7718 7 1 2 23405 33909
0 7719 5 1 1 7718
0 7720 7 1 2 25364 32471
0 7721 5 1 1 7720
0 7722 7 1 2 7719 7721
0 7723 5 8 1 7722
0 7724 7 1 2 22810 30365
0 7725 5 1 1 7724
0 7726 7 2 2 24749 29057
0 7727 5 2 1 34923
0 7728 7 1 2 26149 34924
0 7729 5 1 1 7728
0 7730 7 1 2 7725 7729
0 7731 5 1 1 7730
0 7732 7 1 2 34915 7731
0 7733 5 1 1 7732
0 7734 7 20 2 32475 33915
0 7735 7 1 2 32820 30366
0 7736 5 1 1 7735
0 7737 7 11 2 22811 22935
0 7738 5 1 1 34947
0 7739 7 5 2 25365 23538
0 7740 7 2 2 34948 34958
0 7741 7 1 2 26150 34963
0 7742 5 1 1 7741
0 7743 7 1 2 7736 7742
0 7744 5 1 1 7743
0 7745 7 1 2 34927 7744
0 7746 5 1 1 7745
0 7747 7 1 2 7733 7746
0 7748 5 1 1 7747
0 7749 7 1 2 26750 7748
0 7750 5 1 1 7749
0 7751 7 1 2 22812 34916
0 7752 5 1 1 7751
0 7753 7 1 2 32821 32452
0 7754 5 1 1 7753
0 7755 7 1 2 7752 7754
0 7756 5 3 1 7755
0 7757 7 1 2 26448 29186
0 7758 7 1 2 34965 7757
0 7759 5 1 1 7758
0 7760 7 1 2 7750 7759
0 7761 5 1 1 7760
0 7762 7 1 2 25982 7761
0 7763 5 1 1 7762
0 7764 7 2 2 29069 33076
0 7765 5 1 1 34968
0 7766 7 1 2 25426 29828
0 7767 5 1 1 7766
0 7768 7 5 2 23463 29870
0 7769 5 1 1 34970
0 7770 7 1 2 7767 7769
0 7771 5 14 1 7770
0 7772 7 1 2 22813 34975
0 7773 5 2 1 7772
0 7774 7 2 2 26844 32453
0 7775 5 1 1 34991
0 7776 7 1 2 34989 7775
0 7777 5 6 1 7776
0 7778 7 1 2 23406 34993
0 7779 5 1 1 7778
0 7780 7 1 2 25366 33825
0 7781 5 1 1 7780
0 7782 7 1 2 7779 7781
0 7783 5 2 1 7782
0 7784 7 1 2 34969 34999
0 7785 5 1 1 7784
0 7786 7 4 2 24750 23033
0 7787 5 1 1 35001
0 7788 7 1 2 28410 7787
0 7789 5 1 1 7788
0 7790 7 1 2 33023 7789
0 7791 7 1 2 34917 7790
0 7792 5 1 1 7791
0 7793 7 1 2 32822 32287
0 7794 5 1 1 7793
0 7795 7 1 2 33372 33000
0 7796 5 1 1 7795
0 7797 7 1 2 7794 7796
0 7798 5 1 1 7797
0 7799 7 1 2 34928 7798
0 7800 5 1 1 7799
0 7801 7 1 2 7792 7800
0 7802 5 1 1 7801
0 7803 7 1 2 33444 7802
0 7804 5 1 1 7803
0 7805 7 1 2 7785 7804
0 7806 5 1 1 7805
0 7807 7 1 2 25068 7806
0 7808 5 1 1 7807
0 7809 7 1 2 23034 28473
0 7810 5 1 1 7809
0 7811 7 1 2 1036 7810
0 7812 5 1 1 7811
0 7813 7 1 2 29829 26449
0 7814 5 1 1 7813
0 7815 7 1 2 22936 29797
0 7816 5 1 1 7815
0 7817 7 1 2 7814 7816
0 7818 5 1 1 7817
0 7819 7 1 2 28977 7818
0 7820 5 1 1 7819
0 7821 7 4 2 26071 26450
0 7822 7 6 2 25427 25983
0 7823 7 1 2 24751 35009
0 7824 5 1 1 7823
0 7825 7 2 2 22814 33859
0 7826 5 2 1 35015
0 7827 7 1 2 7824 35017
0 7828 5 4 1 7827
0 7829 7 1 2 35005 35019
0 7830 5 1 1 7829
0 7831 7 1 2 7820 7830
0 7832 5 1 1 7831
0 7833 7 1 2 23407 7832
0 7834 5 1 1 7833
0 7835 7 1 2 26451 33373
0 7836 7 1 2 34094 7835
0 7837 5 1 1 7836
0 7838 7 1 2 7834 7837
0 7839 5 1 1 7838
0 7840 7 1 2 7812 7839
0 7841 5 1 1 7840
0 7842 7 1 2 7808 7841
0 7843 7 1 2 7763 7842
0 7844 5 1 1 7843
0 7845 7 1 2 25528 7844
0 7846 5 1 1 7845
0 7847 7 1 2 23408 33021
0 7848 5 1 1 7847
0 7849 7 1 2 26072 26911
0 7850 7 1 2 33001 7849
0 7851 5 1 1 7850
0 7852 7 1 2 7848 7851
0 7853 5 1 1 7852
0 7854 7 1 2 28978 7853
0 7855 5 1 1 7854
0 7856 7 1 2 25984 28725
0 7857 7 1 2 33026 7856
0 7858 5 1 1 7857
0 7859 7 1 2 7855 7858
0 7860 5 1 1 7859
0 7861 7 1 2 29105 7860
0 7862 5 1 1 7861
0 7863 7 2 2 25985 33077
0 7864 7 1 2 32834 35023
0 7865 5 1 1 7864
0 7866 7 1 2 29187 31882
0 7867 7 1 2 32917 7866
0 7868 5 1 1 7867
0 7869 7 1 2 7865 7868
0 7870 5 1 1 7869
0 7871 7 1 2 32722 7870
0 7872 5 1 1 7871
0 7873 7 1 2 32544 33055
0 7874 7 1 2 35024 7873
0 7875 5 1 1 7874
0 7876 7 7 2 24752 22937
0 7877 5 1 1 35025
0 7878 7 3 2 35026 32629
0 7879 5 1 1 35032
0 7880 7 2 2 30466 35033
0 7881 5 1 1 35035
0 7882 7 1 2 26377 30563
0 7883 7 1 2 35036 7882
0 7884 5 1 1 7883
0 7885 7 1 2 7875 7884
0 7886 7 1 2 7872 7885
0 7887 7 1 2 7862 7886
0 7888 7 1 2 7846 7887
0 7889 5 1 1 7888
0 7890 7 1 2 23918 7889
0 7891 5 1 1 7890
0 7892 7 1 2 7717 7891
0 7893 5 1 1 7892
0 7894 7 1 2 26309 7893
0 7895 5 1 1 7894
0 7896 7 1 2 33564 30567
0 7897 5 2 1 7896
0 7898 7 1 2 29106 35037
0 7899 5 1 1 7898
0 7900 7 1 2 23539 33522
0 7901 5 1 1 7900
0 7902 7 1 2 7899 7901
0 7903 5 1 1 7902
0 7904 7 1 2 27522 7903
0 7905 5 1 1 7904
0 7906 7 1 2 23540 29188
0 7907 5 1 1 7906
0 7908 7 1 2 28522 26751
0 7909 5 2 1 7908
0 7910 7 1 2 25529 27623
0 7911 7 1 2 35039 7910
0 7912 5 1 1 7911
0 7913 7 1 2 7907 7912
0 7914 5 1 1 7913
0 7915 7 1 2 25069 7914
0 7916 5 1 1 7915
0 7917 7 1 2 7916 7578
0 7918 5 1 1 7917
0 7919 7 1 2 22938 7918
0 7920 5 1 1 7919
0 7921 7 2 2 29313 33452
0 7922 7 1 2 35041 29353
0 7923 5 1 1 7922
0 7924 7 1 2 7920 7923
0 7925 5 1 1 7924
0 7926 7 1 2 24095 7925
0 7927 5 1 1 7926
0 7928 7 1 2 7905 7927
0 7929 5 1 1 7928
0 7930 7 3 2 23409 31118
0 7931 7 1 2 35043 26341
0 7932 7 1 2 7929 7931
0 7933 5 1 1 7932
0 7934 7 1 2 7895 7933
0 7935 5 1 1 7934
0 7936 7 1 2 22721 7935
0 7937 5 1 1 7936
0 7938 7 4 2 24753 27606
0 7939 7 1 2 26912 35046
0 7940 5 1 1 7939
0 7941 7 1 2 24009 28503
0 7942 7 1 2 33374 7941
0 7943 5 1 1 7942
0 7944 7 1 2 7940 7943
0 7945 5 1 1 7944
0 7946 7 1 2 34900 7945
0 7947 5 1 1 7946
0 7948 7 2 2 28523 33453
0 7949 7 12 2 24754 24867
0 7950 7 1 2 26913 35052
0 7951 7 1 2 35050 7950
0 7952 5 1 1 7951
0 7953 7 1 2 7947 7952
0 7954 5 1 1 7953
0 7955 7 1 2 26738 7954
0 7956 5 1 1 7955
0 7957 7 2 2 24265 26914
0 7958 7 3 2 24755 32390
0 7959 7 1 2 26151 33454
0 7960 7 1 2 35066 7959
0 7961 7 1 2 35064 7960
0 7962 5 1 1 7961
0 7963 7 1 2 7956 7962
0 7964 5 1 1 7963
0 7965 7 1 2 25890 7964
0 7966 5 1 1 7965
0 7967 7 2 2 32984 34901
0 7968 7 1 2 27033 30906
0 7969 7 1 2 32698 7968
0 7970 7 1 2 35069 7969
0 7971 5 1 1 7970
0 7972 7 1 2 7966 7971
0 7973 5 1 1 7972
0 7974 7 1 2 34929 7973
0 7975 5 1 1 7974
0 7976 7 2 2 34976 34292
0 7977 5 1 1 35071
0 7978 7 1 2 23410 33798
0 7979 5 1 1 7978
0 7980 7 1 2 7977 7979
0 7981 5 3 1 7980
0 7982 7 1 2 22815 35073
0 7983 5 1 1 7982
0 7984 7 1 2 26926 33921
0 7985 5 1 1 7984
0 7986 7 1 2 7983 7985
0 7987 5 1 1 7986
0 7988 7 1 2 29660 7987
0 7989 5 1 1 7988
0 7990 7 1 2 26993 32480
0 7991 5 1 1 7990
0 7992 7 1 2 24096 26931
0 7993 5 1 1 7992
0 7994 7 1 2 7991 7993
0 7995 5 1 1 7994
0 7996 7 1 2 30357 7995
0 7997 5 1 1 7996
0 7998 7 1 2 7989 7997
0 7999 5 1 1 7998
0 8000 7 1 2 34876 7999
0 8001 5 1 1 8000
0 8002 7 1 2 22816 27607
0 8003 5 2 1 8002
0 8004 7 1 2 24756 28504
0 8005 5 1 1 8004
0 8006 7 1 2 35076 8005
0 8007 5 3 1 8006
0 8008 7 1 2 34902 35078
0 8009 5 1 1 8008
0 8010 7 11 2 22817 24868
0 8011 7 1 2 35081 35051
0 8012 5 1 1 8011
0 8013 7 1 2 8009 8012
0 8014 5 1 1 8013
0 8015 7 1 2 26739 8014
0 8016 5 1 1 8015
0 8017 7 4 2 33550 30252
0 8018 7 2 2 22818 35092
0 8019 7 1 2 29189 35096
0 8020 5 1 1 8019
0 8021 7 1 2 8016 8020
0 8022 5 1 1 8021
0 8023 7 1 2 35074 8022
0 8024 5 1 1 8023
0 8025 7 2 2 26740 35027
0 8026 5 3 1 35098
0 8027 7 2 2 22819 33523
0 8028 5 1 1 35103
0 8029 7 1 2 35100 8028
0 8030 5 1 1 8029
0 8031 7 1 2 35075 8030
0 8032 5 1 1 8031
0 8033 7 5 2 26741 34949
0 8034 7 1 2 26994 35105
0 8035 5 1 1 8034
0 8036 7 2 2 25530 27805
0 8037 7 1 2 26869 35110
0 8038 7 1 2 35065 8037
0 8039 5 1 1 8038
0 8040 7 1 2 8035 8039
0 8041 5 1 1 8040
0 8042 7 1 2 34930 8041
0 8043 5 1 1 8042
0 8044 7 1 2 8032 8043
0 8045 5 1 1 8044
0 8046 7 1 2 28641 8045
0 8047 5 1 1 8046
0 8048 7 1 2 8024 8047
0 8049 7 1 2 8001 8048
0 8050 7 1 2 7975 8049
0 8051 5 1 1 8050
0 8052 7 1 2 24681 26310
0 8053 7 1 2 8051 8052
0 8054 5 1 1 8053
0 8055 7 1 2 28233 8054
0 8056 7 1 2 7937 8055
0 8057 5 1 1 8056
0 8058 7 4 2 25891 26311
0 8059 7 4 2 24183 26452
0 8060 5 1 1 35116
0 8061 7 1 2 22722 35000
0 8062 5 1 1 8061
0 8063 7 2 2 30334 33369
0 8064 5 1 1 35120
0 8065 7 1 2 23464 35121
0 8066 5 1 1 8065
0 8067 7 1 2 8062 8066
0 8068 5 3 1 8067
0 8069 7 1 2 35117 35122
0 8070 5 1 1 8069
0 8071 7 1 2 30939 32481
0 8072 5 1 1 8071
0 8073 7 9 2 22723 24757
0 8074 7 3 2 24097 35125
0 8075 5 1 1 35134
0 8076 7 2 2 35010 35135
0 8077 7 1 2 23411 35137
0 8078 5 1 1 8077
0 8079 7 1 2 8072 8078
0 8080 5 2 1 8079
0 8081 7 1 2 28505 34903
0 8082 5 1 1 8081
0 8083 7 1 2 29846 8082
0 8084 5 1 1 8083
0 8085 7 1 2 35139 8084
0 8086 5 1 1 8085
0 8087 7 1 2 8070 8086
0 8088 5 1 1 8087
0 8089 7 1 2 26742 8088
0 8090 5 1 1 8089
0 8091 7 1 2 29661 35123
0 8092 5 1 1 8091
0 8093 7 1 2 30358 35140
0 8094 5 1 1 8093
0 8095 7 1 2 8092 8094
0 8096 5 1 1 8095
0 8097 7 1 2 34877 8096
0 8098 5 1 1 8097
0 8099 7 1 2 29277 26557
0 8100 5 1 1 8099
0 8101 7 1 2 25486 31777
0 8102 5 1 1 8101
0 8103 7 1 2 8100 8102
0 8104 7 1 2 7765 8103
0 8105 5 1 1 8104
0 8106 7 1 2 33455 8105
0 8107 7 1 2 35124 8106
0 8108 5 1 1 8107
0 8109 7 1 2 8098 8108
0 8110 7 1 2 8090 8109
0 8111 5 1 1 8110
0 8112 7 1 2 35112 8111
0 8113 5 1 1 8112
0 8114 7 1 2 28250 8113
0 8115 5 1 1 8114
0 8116 7 1 2 28320 29418
0 8117 7 1 2 8115 8116
0 8118 7 1 2 8057 8117
0 8119 5 1 1 8118
0 8120 7 1 2 31781 34898
0 8121 5 6 1 8120
0 8122 7 2 2 28308 26995
0 8123 5 1 1 35147
0 8124 7 1 2 2577 8123
0 8125 5 2 1 8124
0 8126 7 1 2 27130 35149
0 8127 5 1 1 8126
0 8128 7 1 2 27075 31304
0 8129 5 1 1 8128
0 8130 7 1 2 8127 8129
0 8131 5 2 1 8130
0 8132 7 1 2 31469 35151
0 8133 5 1 1 8132
0 8134 7 1 2 31023 33893
0 8135 5 1 1 8134
0 8136 7 1 2 34129 30893
0 8137 5 1 1 8136
0 8138 7 3 2 8135 8137
0 8139 7 1 2 34781 35153
0 8140 5 1 1 8139
0 8141 7 1 2 28093 31119
0 8142 7 1 2 29978 8141
0 8143 5 1 1 8142
0 8144 7 1 2 25292 30815
0 8145 5 1 1 8144
0 8146 7 1 2 23345 6937
0 8147 5 2 1 8146
0 8148 7 2 2 24577 27443
0 8149 5 1 1 35158
0 8150 7 1 2 35156 35159
0 8151 7 1 2 8145 8150
0 8152 5 1 1 8151
0 8153 7 1 2 8143 8152
0 8154 5 1 1 8153
0 8155 7 1 2 32088 8154
0 8156 5 1 1 8155
0 8157 7 1 2 8140 8156
0 8158 5 1 1 8157
0 8159 7 1 2 28979 8158
0 8160 5 1 1 8159
0 8161 7 1 2 8133 8160
0 8162 5 1 1 8161
0 8163 7 1 2 35141 8162
0 8164 5 1 1 8163
0 8165 7 1 2 22820 34888
0 8166 5 1 1 8165
0 8167 7 1 2 35101 8166
0 8168 5 6 1 8167
0 8169 7 1 2 34977 35154
0 8170 5 1 1 8169
0 8171 7 1 2 25293 33799
0 8172 5 1 1 8171
0 8173 7 2 2 33910 28745
0 8174 5 1 1 35166
0 8175 7 1 2 23919 35167
0 8176 5 1 1 8175
0 8177 7 1 2 8172 8176
0 8178 5 1 1 8177
0 8179 7 1 2 24578 8178
0 8180 5 1 1 8179
0 8181 7 5 2 25428 29892
0 8182 7 1 2 30886 35168
0 8183 5 1 1 8182
0 8184 7 1 2 8180 8183
0 8185 5 1 1 8184
0 8186 7 1 2 32089 8185
0 8187 5 1 1 8186
0 8188 7 1 2 8170 8187
0 8189 5 1 1 8188
0 8190 7 1 2 35160 8189
0 8191 5 1 1 8190
0 8192 7 1 2 35126 34889
0 8193 5 1 1 8192
0 8194 7 5 2 26241 32162
0 8195 7 1 2 35173 33355
0 8196 5 1 1 8195
0 8197 7 1 2 8193 8196
0 8198 5 3 1 8197
0 8199 7 1 2 35150 35178
0 8200 5 1 1 8199
0 8201 7 2 2 22821 30596
0 8202 7 2 2 30868 30440
0 8203 7 1 2 35181 35183
0 8204 5 1 1 8203
0 8205 7 1 2 27336 34890
0 8206 7 1 2 30897 8205
0 8207 5 1 1 8206
0 8208 7 1 2 8204 8207
0 8209 5 1 1 8208
0 8210 7 1 2 27076 8209
0 8211 5 1 1 8210
0 8212 7 1 2 8200 8211
0 8213 5 1 1 8212
0 8214 7 1 2 34931 8213
0 8215 5 1 1 8214
0 8216 7 1 2 8191 8215
0 8217 5 1 1 8216
0 8218 7 1 2 28642 8217
0 8219 5 1 1 8218
0 8220 7 1 2 8164 8219
0 8221 5 1 1 8220
0 8222 7 3 2 25691 26312
0 8223 7 1 2 25212 35185
0 8224 7 1 2 8221 8223
0 8225 5 1 1 8224
0 8226 7 1 2 8119 8225
0 8227 5 1 1 8226
0 8228 7 1 2 22443 8227
0 8229 5 1 1 8228
0 8230 7 1 2 26996 29222
0 8231 5 1 1 8230
0 8232 7 1 2 28135 31145
0 8233 5 1 1 8232
0 8234 7 1 2 8231 8233
0 8235 5 2 1 8234
0 8236 7 1 2 27131 35188
0 8237 5 1 1 8236
0 8238 7 1 2 27077 31528
0 8239 5 1 1 8238
0 8240 7 1 2 8237 8239
0 8241 5 1 1 8240
0 8242 7 1 2 31470 8241
0 8243 5 1 1 8242
0 8244 7 1 2 27311 34118
0 8245 5 1 1 8244
0 8246 7 1 2 34134 31160
0 8247 5 1 1 8246
0 8248 7 1 2 8245 8247
0 8249 5 2 1 8248
0 8250 7 1 2 34782 35190
0 8251 5 1 1 8250
0 8252 7 1 2 30824 29223
0 8253 5 1 1 8252
0 8254 7 1 2 5696 8253
0 8255 5 1 1 8254
0 8256 7 1 2 32090 8255
0 8257 5 1 1 8256
0 8258 7 1 2 8251 8257
0 8259 5 1 1 8258
0 8260 7 1 2 28980 8259
0 8261 5 1 1 8260
0 8262 7 1 2 8243 8261
0 8263 5 1 1 8262
0 8264 7 1 2 35142 8263
0 8265 5 1 1 8264
0 8266 7 1 2 34978 35191
0 8267 5 1 1 8266
0 8268 7 1 2 33800 29224
0 8269 5 1 1 8268
0 8270 7 1 2 24010 33911
0 8271 7 2 2 30780 8270
0 8272 5 1 1 35192
0 8273 7 1 2 33812 31344
0 8274 5 1 1 8273
0 8275 7 1 2 8272 8274
0 8276 5 1 1 8275
0 8277 7 1 2 28136 8276
0 8278 5 1 1 8277
0 8279 7 1 2 8269 8278
0 8280 5 1 1 8279
0 8281 7 1 2 32091 8280
0 8282 5 1 1 8281
0 8283 7 1 2 8267 8282
0 8284 5 1 1 8283
0 8285 7 1 2 35161 8284
0 8286 5 1 1 8285
0 8287 7 1 2 35179 35189
0 8288 5 1 1 8287
0 8289 7 2 2 24758 31202
0 8290 7 2 2 31192 35194
0 8291 7 1 2 34878 35196
0 8292 5 1 1 8291
0 8293 7 1 2 30597 31330
0 8294 7 1 2 31497 8293
0 8295 5 1 1 8294
0 8296 7 1 2 8292 8295
0 8297 5 1 1 8296
0 8298 7 1 2 27312 8297
0 8299 5 1 1 8298
0 8300 7 1 2 35174 27772
0 8301 5 1 1 8300
0 8302 7 2 2 34891 31355
0 8303 5 1 1 35198
0 8304 7 1 2 8301 8303
0 8305 5 1 1 8304
0 8306 7 1 2 31161 8305
0 8307 5 1 1 8306
0 8308 7 1 2 8299 8307
0 8309 5 1 1 8308
0 8310 7 1 2 27078 8309
0 8311 5 1 1 8310
0 8312 7 1 2 8288 8311
0 8313 5 1 1 8312
0 8314 7 1 2 34932 8313
0 8315 5 1 1 8314
0 8316 7 1 2 8286 8315
0 8317 5 1 1 8316
0 8318 7 1 2 28643 8317
0 8319 5 1 1 8318
0 8320 7 1 2 8265 8319
0 8321 5 1 1 8320
0 8322 7 1 2 24444 35186
0 8323 7 1 2 8321 8322
0 8324 5 1 1 8323
0 8325 7 1 2 8229 8324
0 8326 5 1 1 8325
0 8327 7 1 2 23622 8326
0 8328 5 1 1 8327
0 8329 7 1 2 30094 28483
0 8330 5 1 1 8329
0 8331 7 1 2 28506 8330
0 8332 5 1 1 8331
0 8333 7 2 2 23035 29860
0 8334 7 4 2 25621 26242
0 8335 5 2 1 35202
0 8336 7 1 2 35206 28899
0 8337 5 7 1 8336
0 8338 7 1 2 35200 35208
0 8339 5 1 1 8338
0 8340 7 1 2 8332 8339
0 8341 5 1 1 8340
0 8342 7 2 2 27763 29419
0 8343 7 1 2 8341 35215
0 8344 5 1 1 8343
0 8345 7 1 2 26508 28787
0 8346 7 1 2 26752 8345
0 8347 7 1 2 30803 8346
0 8348 7 1 2 29662 8347
0 8349 5 1 1 8348
0 8350 7 1 2 8344 8349
0 8351 5 1 1 8350
0 8352 7 1 2 22822 8351
0 8353 5 1 1 8352
0 8354 7 1 2 23465 27608
0 8355 5 1 1 8354
0 8356 7 1 2 25429 28507
0 8357 5 1 1 8356
0 8358 7 1 2 8355 8357
0 8359 5 2 1 8358
0 8360 7 1 2 22939 35217
0 8361 5 1 1 8360
0 8362 7 3 2 24869 23466
0 8363 7 1 2 26800 35219
0 8364 5 1 1 8363
0 8365 7 1 2 8361 8364
0 8366 5 1 1 8365
0 8367 7 2 2 26509 31705
0 8368 7 1 2 26753 31977
0 8369 7 1 2 35222 8368
0 8370 7 1 2 8366 8369
0 8371 5 1 1 8370
0 8372 7 1 2 8353 8371
0 8373 5 1 1 8372
0 8374 7 1 2 25531 8373
0 8375 5 1 1 8374
0 8376 7 2 2 31857 30449
0 8377 7 2 2 26510 35224
0 8378 7 1 2 28964 32288
0 8379 5 1 1 8378
0 8380 7 2 2 23036 25430
0 8381 5 2 1 35228
0 8382 7 1 2 35230 33306
0 8383 5 1 1 8382
0 8384 7 1 2 24759 33024
0 8385 7 1 2 8383 8384
0 8386 5 1 1 8385
0 8387 7 1 2 8379 8386
0 8388 5 1 1 8387
0 8389 7 1 2 35226 8388
0 8390 5 1 1 8389
0 8391 7 3 2 32985 30527
0 8392 7 1 2 26313 35232
0 8393 7 2 2 33867 8392
0 8394 5 1 1 35235
0 8395 7 1 2 25487 8394
0 8396 7 1 2 8390 8395
0 8397 5 1 1 8396
0 8398 7 1 2 25431 31978
0 8399 7 1 2 35223 8398
0 8400 7 1 2 33078 8399
0 8401 5 1 1 8400
0 8402 7 3 2 26696 30761
0 8403 5 2 1 35237
0 8404 7 2 2 25622 26152
0 8405 7 1 2 24266 35242
0 8406 5 1 1 8405
0 8407 7 1 2 35240 8406
0 8408 5 2 1 8407
0 8409 7 3 2 23412 28359
0 8410 7 2 2 35246 31561
0 8411 7 1 2 23467 35249
0 8412 7 1 2 35244 8411
0 8413 5 1 1 8412
0 8414 7 1 2 23541 8413
0 8415 7 1 2 8401 8414
0 8416 5 1 1 8415
0 8417 7 1 2 22940 8416
0 8418 7 1 2 8397 8417
0 8419 5 1 1 8418
0 8420 7 1 2 23542 35236
0 8421 5 1 1 8420
0 8422 7 1 2 28981 32284
0 8423 5 1 1 8422
0 8424 7 2 2 24760 35229
0 8425 7 1 2 34907 35251
0 8426 5 1 1 8425
0 8427 7 1 2 8423 8426
0 8428 5 1 1 8427
0 8429 7 1 2 8428 35227
0 8430 5 1 1 8429
0 8431 7 1 2 8421 8430
0 8432 5 1 1 8431
0 8433 7 1 2 24870 8432
0 8434 5 1 1 8433
0 8435 7 1 2 24098 8434
0 8436 7 1 2 8419 8435
0 8437 7 1 2 8375 8436
0 8438 5 1 1 8437
0 8439 7 2 2 24184 34879
0 8440 7 6 2 25488 28788
0 8441 7 4 2 35255 30804
0 8442 7 1 2 35253 35261
0 8443 5 1 1 8442
0 8444 7 3 2 23468 23695
0 8445 7 2 2 28604 35265
0 8446 7 2 2 28360 35268
0 8447 7 1 2 26153 33428
0 8448 5 4 1 8447
0 8449 7 1 2 35272 29709
0 8450 7 1 2 35270 8449
0 8451 5 1 1 8450
0 8452 7 1 2 8443 8451
0 8453 5 1 1 8452
0 8454 7 1 2 22941 8453
0 8455 5 1 1 8454
0 8456 7 1 2 34880 28644
0 8457 5 1 1 8456
0 8458 7 1 2 32279 8457
0 8459 5 1 1 8458
0 8460 7 3 2 25367 25692
0 8461 7 3 2 31322 35276
0 8462 7 5 2 24871 25213
0 8463 7 1 2 35279 35282
0 8464 7 1 2 8459 8463
0 8465 5 1 1 8464
0 8466 7 1 2 8455 8465
0 8467 5 1 1 8466
0 8468 7 1 2 23623 8467
0 8469 5 1 1 8468
0 8470 7 1 2 34881 29663
0 8471 5 1 1 8470
0 8472 7 6 2 24872 23037
0 8473 7 6 2 26243 35287
0 8474 7 1 2 27609 35293
0 8475 5 1 1 8474
0 8476 7 1 2 8471 8475
0 8477 5 3 1 8476
0 8478 7 5 2 28789 29585
0 8479 7 1 2 35187 35302
0 8480 7 1 2 35299 8479
0 8481 5 1 1 8480
0 8482 7 1 2 8469 8481
0 8483 5 1 1 8482
0 8484 7 1 2 24761 8483
0 8485 5 1 1 8484
0 8486 7 1 2 32713 30426
0 8487 5 1 1 8486
0 8488 7 4 2 24963 23469
0 8489 7 1 2 29199 35307
0 8490 5 1 1 8489
0 8491 7 1 2 8487 8490
0 8492 5 1 1 8491
0 8493 7 1 2 22942 8492
0 8494 5 1 1 8493
0 8495 7 1 2 23543 28609
0 8496 5 1 1 8495
0 8497 7 1 2 26443 8496
0 8498 5 1 1 8497
0 8499 7 1 2 35220 8498
0 8500 5 1 1 8499
0 8501 7 1 2 8494 8500
0 8502 5 1 1 8501
0 8503 7 1 2 35273 8502
0 8504 5 1 1 8503
0 8505 7 2 2 27492 26410
0 8506 5 1 1 35311
0 8507 7 1 2 8506 30095
0 8508 5 1 1 8507
0 8509 7 1 2 25489 8508
0 8510 5 1 1 8509
0 8511 7 1 2 24873 35312
0 8512 5 1 1 8511
0 8513 7 1 2 28660 30054
0 8514 5 1 1 8513
0 8515 7 1 2 8512 8514
0 8516 7 1 2 8510 8515
0 8517 5 1 1 8516
0 8518 7 3 2 23470 25532
0 8519 7 1 2 24185 35313
0 8520 7 1 2 8517 8519
0 8521 5 1 1 8520
0 8522 7 1 2 8504 8521
0 8523 5 1 1 8522
0 8524 7 1 2 35250 8523
0 8525 5 1 1 8524
0 8526 7 1 2 26073 8525
0 8527 7 1 2 8485 8526
0 8528 5 1 1 8527
0 8529 7 1 2 22724 8528
0 8530 7 1 2 8438 8529
0 8531 5 1 1 8530
0 8532 7 1 2 31471 28726
0 8533 5 1 1 8532
0 8534 7 1 2 28982 32137
0 8535 5 1 1 8534
0 8536 7 1 2 8533 8535
0 8537 5 1 1 8536
0 8538 7 1 2 35143 8537
0 8539 5 1 1 8538
0 8540 7 1 2 34918 35162
0 8541 5 1 1 8540
0 8542 7 1 2 25368 35106
0 8543 5 1 1 8542
0 8544 7 2 2 32823 34892
0 8545 5 1 1 35316
0 8546 7 1 2 8543 8545
0 8547 5 1 1 8546
0 8548 7 1 2 34933 8547
0 8549 5 1 1 8548
0 8550 7 1 2 8541 8549
0 8551 5 1 1 8550
0 8552 7 1 2 28645 8551
0 8553 5 1 1 8552
0 8554 7 1 2 8539 8553
0 8555 5 1 1 8554
0 8556 7 1 2 26511 28019
0 8557 7 1 2 29399 8556
0 8558 7 1 2 8555 8557
0 8559 5 1 1 8558
0 8560 7 1 2 8531 8559
0 8561 5 1 1 8560
0 8562 7 1 2 22606 8561
0 8563 5 1 1 8562
0 8564 7 1 2 3124 32449
0 8565 7 4 2 32744 8564
0 8566 7 1 2 22823 35318
0 8567 5 1 1 8566
0 8568 7 3 2 24762 32227
0 8569 7 1 2 32454 35322
0 8570 5 1 1 8569
0 8571 7 1 2 8567 8570
0 8572 5 1 1 8571
0 8573 7 1 2 22725 8572
0 8574 5 1 1 8573
0 8575 7 1 2 28875 34966
0 8576 5 1 1 8575
0 8577 7 1 2 8574 8576
0 8578 5 2 1 8577
0 8579 7 1 2 35300 35325
0 8580 5 1 1 8579
0 8581 7 1 2 34882 30359
0 8582 5 1 1 8581
0 8583 7 1 2 4196 8582
0 8584 5 2 1 8583
0 8585 7 1 2 32242 32482
0 8586 5 1 1 8585
0 8587 7 2 2 25432 34551
0 8588 7 1 2 27419 35329
0 8589 5 1 1 8588
0 8590 7 1 2 8586 8589
0 8591 5 1 1 8590
0 8592 7 1 2 35327 8591
0 8593 5 1 1 8592
0 8594 7 1 2 8580 8593
0 8595 5 1 1 8594
0 8596 7 5 2 25693 26512
0 8597 7 1 2 35331 30575
0 8598 7 1 2 8595 8597
0 8599 5 1 1 8598
0 8600 7 1 2 8563 8599
0 8601 5 1 1 8600
0 8602 7 1 2 22444 8601
0 8603 5 1 1 8602
0 8604 7 2 2 26074 28805
0 8605 7 1 2 29209 35336
0 8606 5 1 1 8605
0 8607 7 3 2 25369 28075
0 8608 7 1 2 33912 35338
0 8609 5 1 1 8608
0 8610 7 1 2 8606 8609
0 8611 5 3 1 8610
0 8612 7 1 2 22824 35341
0 8613 5 1 1 8612
0 8614 7 1 2 23257 28671
0 8615 7 1 2 33922 8614
0 8616 5 1 1 8615
0 8617 7 1 2 8613 8616
0 8618 5 1 1 8617
0 8619 7 1 2 22726 8618
0 8620 5 1 1 8619
0 8621 7 1 2 30625 34967
0 8622 5 1 1 8621
0 8623 7 1 2 8620 8622
0 8624 5 1 1 8623
0 8625 7 1 2 22607 8624
0 8626 5 1 1 8625
0 8627 7 1 2 30644 35326
0 8628 5 1 1 8627
0 8629 7 1 2 8626 8628
0 8630 5 1 1 8629
0 8631 7 1 2 35301 8630
0 8632 5 1 1 8631
0 8633 7 1 2 32855 32483
0 8634 5 1 1 8633
0 8635 7 2 2 33133 32145
0 8636 5 1 1 35344
0 8637 7 1 2 33200 35345
0 8638 5 1 1 8637
0 8639 7 1 2 8634 8638
0 8640 5 1 1 8639
0 8641 7 1 2 35328 8640
0 8642 5 1 1 8641
0 8643 7 1 2 8632 8642
0 8644 5 1 1 8643
0 8645 7 1 2 24445 35332
0 8646 7 1 2 8644 8645
0 8647 5 1 1 8646
0 8648 7 1 2 8603 8647
0 8649 5 1 1 8648
0 8650 7 1 2 24011 8649
0 8651 5 1 1 8650
0 8652 7 1 2 29248 4042
0 8653 5 1 1 8652
0 8654 7 1 2 30314 32141
0 8655 5 1 1 8654
0 8656 7 1 2 8653 8655
0 8657 5 1 1 8656
0 8658 7 1 2 28983 8657
0 8659 5 1 1 8658
0 8660 7 1 2 31405 29249
0 8661 5 1 1 8660
0 8662 7 1 2 30315 31791
0 8663 5 1 1 8662
0 8664 7 1 2 8661 8663
0 8665 5 3 1 8664
0 8666 7 1 2 31472 35346
0 8667 5 1 1 8666
0 8668 7 1 2 8659 8667
0 8669 5 1 1 8668
0 8670 7 1 2 35144 8669
0 8671 5 1 1 8670
0 8672 7 1 2 30989 32476
0 8673 5 1 1 8672
0 8674 7 1 2 32069 33916
0 8675 5 1 1 8674
0 8676 7 1 2 8673 8675
0 8677 7 1 2 29250 8676
0 8678 5 1 1 8677
0 8679 7 1 2 31011 33913
0 8680 7 1 2 30316 8679
0 8681 5 1 1 8680
0 8682 7 1 2 8678 8681
0 8683 5 1 1 8682
0 8684 7 1 2 35163 8683
0 8685 5 1 1 8684
0 8686 7 1 2 32092 35107
0 8687 5 1 1 8686
0 8688 7 1 2 22727 35317
0 8689 5 1 1 8688
0 8690 7 1 2 8687 8689
0 8691 5 1 1 8690
0 8692 7 1 2 29251 8691
0 8693 5 1 1 8692
0 8694 7 2 2 30317 30028
0 8695 7 7 2 24763 25370
0 8696 5 1 1 35351
0 8697 7 1 2 34883 35352
0 8698 7 1 2 35349 8697
0 8699 5 1 1 8698
0 8700 7 1 2 8693 8699
0 8701 5 1 1 8700
0 8702 7 1 2 34934 8701
0 8703 5 1 1 8702
0 8704 7 1 2 8685 8703
0 8705 5 1 1 8704
0 8706 7 1 2 28646 8705
0 8707 5 1 1 8706
0 8708 7 1 2 8671 8707
0 8709 5 1 1 8708
0 8710 7 3 2 25986 26513
0 8711 7 1 2 25694 35358
0 8712 7 1 2 8709 8711
0 8713 5 1 1 8712
0 8714 7 1 2 8651 8713
0 8715 5 1 1 8714
0 8716 7 1 2 23920 8715
0 8717 5 1 1 8716
0 8718 7 1 2 25214 33216
0 8719 5 1 1 8718
0 8720 7 1 2 27049 29202
0 8721 5 1 1 8720
0 8722 7 1 2 8719 8721
0 8723 5 2 1 8722
0 8724 7 1 2 24446 35361
0 8725 5 1 1 8724
0 8726 7 1 2 27050 29238
0 8727 5 1 1 8726
0 8728 7 1 2 8725 8727
0 8729 5 2 1 8728
0 8730 7 1 2 27132 35363
0 8731 5 1 1 8730
0 8732 7 1 2 25215 28044
0 8733 5 1 1 8732
0 8734 7 2 2 23258 31323
0 8735 7 1 2 35365 27827
0 8736 5 1 1 8735
0 8737 7 1 2 8733 8736
0 8738 5 2 1 8737
0 8739 7 1 2 24447 35367
0 8740 5 1 1 8739
0 8741 7 1 2 30576 31728
0 8742 5 1 1 8741
0 8743 7 1 2 8740 8742
0 8744 5 2 1 8743
0 8745 7 1 2 27079 35369
0 8746 5 1 1 8745
0 8747 7 1 2 8731 8746
0 8748 5 1 1 8747
0 8749 7 1 2 31473 8748
0 8750 5 1 1 8749
0 8751 7 1 2 25216 32895
0 8752 5 1 1 8751
0 8753 7 1 2 30645 34511
0 8754 5 1 1 8753
0 8755 7 1 2 8752 8754
0 8756 5 2 1 8755
0 8757 7 1 2 24448 35371
0 8758 5 1 1 8757
0 8759 7 1 2 24579 33873
0 8760 5 1 1 8759
0 8761 7 1 2 8758 8760
0 8762 5 2 1 8761
0 8763 7 1 2 34783 35373
0 8764 5 1 1 8763
0 8765 7 1 2 25294 31003
0 8766 5 1 1 8765
0 8767 7 2 2 35157 8766
0 8768 7 1 2 22608 35375
0 8769 5 1 1 8768
0 8770 7 3 2 25987 30467
0 8771 7 2 2 24580 30630
0 8772 7 1 2 35377 35380
0 8773 5 1 1 8772
0 8774 7 1 2 8769 8773
0 8775 5 1 1 8774
0 8776 7 1 2 25217 8775
0 8777 5 1 1 8776
0 8778 7 1 2 29203 34629
0 8779 5 1 1 8778
0 8780 7 1 2 8777 8779
0 8781 5 1 1 8780
0 8782 7 1 2 24449 8781
0 8783 5 1 1 8782
0 8784 7 1 2 34630 29239
0 8785 5 1 1 8784
0 8786 7 1 2 8783 8785
0 8787 5 1 1 8786
0 8788 7 1 2 32093 8787
0 8789 5 1 1 8788
0 8790 7 1 2 8764 8789
0 8791 5 1 1 8790
0 8792 7 1 2 28984 8791
0 8793 5 1 1 8792
0 8794 7 1 2 8750 8793
0 8795 5 1 1 8794
0 8796 7 1 2 35145 8795
0 8797 5 1 1 8796
0 8798 7 1 2 34979 35374
0 8799 5 1 1 8798
0 8800 7 1 2 29204 35169
0 8801 5 1 1 8800
0 8802 7 1 2 25295 34095
0 8803 5 1 1 8802
0 8804 7 1 2 8174 8803
0 8805 5 1 1 8804
0 8806 7 1 2 22609 8805
0 8807 5 1 1 8806
0 8808 7 1 2 28085 33813
0 8809 5 1 1 8808
0 8810 7 1 2 8807 8809
0 8811 5 1 1 8810
0 8812 7 1 2 25218 8811
0 8813 5 1 1 8812
0 8814 7 1 2 8801 8813
0 8815 5 1 1 8814
0 8816 7 1 2 24450 8815
0 8817 5 1 1 8816
0 8818 7 2 2 24099 30391
0 8819 7 4 2 24581 25433
0 8820 7 1 2 27921 35384
0 8821 7 1 2 35382 8820
0 8822 5 1 1 8821
0 8823 7 1 2 8817 8822
0 8824 5 1 1 8823
0 8825 7 1 2 32094 8824
0 8826 5 1 1 8825
0 8827 7 1 2 8799 8826
0 8828 5 1 1 8827
0 8829 7 1 2 35164 8828
0 8830 5 1 1 8829
0 8831 7 1 2 35180 35364
0 8832 5 1 1 8831
0 8833 7 1 2 23346 35199
0 8834 5 1 1 8833
0 8835 7 1 2 28137 27269
0 8836 7 1 2 35175 8835
0 8837 5 1 1 8836
0 8838 7 1 2 8834 8837
0 8839 5 1 1 8838
0 8840 7 1 2 25219 8839
0 8841 5 1 1 8840
0 8842 7 2 2 25296 34884
0 8843 7 1 2 35197 35388
0 8844 5 1 1 8843
0 8845 7 1 2 8841 8844
0 8846 5 1 1 8845
0 8847 7 1 2 24451 8846
0 8848 5 1 1 8847
0 8849 7 2 2 24874 27337
0 8850 7 1 2 35390 31388
0 8851 7 1 2 35389 8850
0 8852 5 1 1 8851
0 8853 7 1 2 8848 8852
0 8854 5 1 1 8853
0 8855 7 1 2 27080 8854
0 8856 5 1 1 8855
0 8857 7 1 2 8832 8856
0 8858 5 1 1 8857
0 8859 7 1 2 34935 8858
0 8860 5 1 1 8859
0 8861 7 1 2 8830 8860
0 8862 5 1 1 8861
0 8863 7 1 2 28647 8862
0 8864 5 1 1 8863
0 8865 7 1 2 8797 8864
0 8866 5 1 1 8865
0 8867 7 1 2 25892 35333
0 8868 7 1 2 8866 8867
0 8869 5 1 1 8868
0 8870 7 1 2 8717 8869
0 8871 5 1 1 8870
0 8872 7 1 2 23110 8871
0 8873 5 1 1 8872
0 8874 7 1 2 32484 33230
0 8875 5 1 1 8874
0 8876 7 2 2 27420 33336
0 8877 7 1 2 30305 35392
0 8878 7 1 2 30940 8877
0 8879 5 1 1 8878
0 8880 7 1 2 8875 8879
0 8881 5 1 1 8880
0 8882 7 2 2 29278 34861
0 8883 7 1 2 30739 35394
0 8884 7 1 2 30547 8883
0 8885 7 1 2 8881 8884
0 8886 5 1 1 8885
0 8887 7 1 2 8873 8886
0 8888 7 1 2 8328 8887
0 8889 5 1 1 8888
0 8890 7 1 2 23800 8889
0 8891 5 1 1 8890
0 8892 7 1 2 34912 30924
0 8893 5 1 1 8892
0 8894 7 1 2 34895 8893
0 8895 5 4 1 8894
0 8896 7 2 2 30505 35396
0 8897 5 1 1 35400
0 8898 7 3 2 31661 30731
0 8899 7 2 2 32396 34913
0 8900 5 1 1 35405
0 8901 7 1 2 34896 8900
0 8902 5 1 1 8901
0 8903 7 1 2 35402 8902
0 8904 5 1 1 8903
0 8905 7 1 2 8897 8904
0 8906 5 1 1 8905
0 8907 7 1 2 34794 8906
0 8908 5 1 1 8907
0 8909 7 1 2 30869 35397
0 8910 7 1 2 34382 8909
0 8911 5 1 1 8910
0 8912 7 1 2 8908 8911
0 8913 5 1 1 8912
0 8914 7 1 2 24012 8913
0 8915 5 1 1 8914
0 8916 7 2 2 25371 31271
0 8917 7 2 2 27692 35407
0 8918 5 1 1 35409
0 8919 7 1 2 23921 31402
0 8920 5 1 1 8919
0 8921 7 1 2 25893 3596
0 8922 5 1 1 8921
0 8923 7 1 2 25297 8922
0 8924 7 1 2 8920 8923
0 8925 5 1 1 8924
0 8926 7 1 2 8918 8925
0 8927 5 1 1 8926
0 8928 7 1 2 35406 8927
0 8929 5 1 1 8928
0 8930 7 1 2 23038 30404
0 8931 7 1 2 31792 8930
0 8932 7 1 2 30485 8931
0 8933 5 1 1 8932
0 8934 7 1 2 8929 8933
0 8935 5 1 1 8934
0 8936 7 1 2 24582 8935
0 8937 5 1 1 8936
0 8938 7 4 2 23922 32397
0 8939 7 1 2 28094 35411
0 8940 7 6 2 25434 25533
0 8941 7 3 2 25372 35415
0 8942 7 1 2 35421 35391
0 8943 7 1 2 8939 8942
0 8944 5 1 1 8943
0 8945 7 1 2 8937 8944
0 8946 5 1 1 8945
0 8947 7 1 2 33382 8946
0 8948 5 1 1 8947
0 8949 7 1 2 8915 8948
0 8950 5 1 1 8949
0 8951 7 1 2 26801 8950
0 8952 5 1 1 8951
0 8953 7 3 2 23039 30732
0 8954 7 4 2 33009 33158
0 8955 7 2 2 24583 35427
0 8956 7 1 2 35424 35431
0 8957 5 1 1 8956
0 8958 7 3 2 25534 24186
0 8959 7 1 2 24964 29893
0 8960 7 1 2 35433 8959
0 8961 7 1 2 28138 8960
0 8962 5 1 1 8961
0 8963 7 1 2 8957 8962
0 8964 5 1 1 8963
0 8965 7 1 2 29107 8964
0 8966 5 1 1 8965
0 8967 7 1 2 27363 33445
0 8968 7 1 2 35425 8967
0 8969 7 1 2 33434 8968
0 8970 5 1 1 8969
0 8971 7 1 2 8966 8970
0 8972 5 1 1 8971
0 8973 7 1 2 32095 8972
0 8974 5 1 1 8973
0 8975 7 1 2 30951 29518
0 8976 5 1 1 8975
0 8977 7 3 2 29533 26863
0 8978 5 1 1 35436
0 8979 7 1 2 8976 8978
0 8980 5 1 1 8979
0 8981 7 1 2 26154 33551
0 8982 5 2 1 8981
0 8983 7 1 2 35439 33073
0 8984 5 4 1 8983
0 8985 7 1 2 24013 35441
0 8986 7 1 2 30749 8985
0 8987 5 1 1 8986
0 8988 7 3 2 25535 31051
0 8989 7 1 2 26155 28758
0 8990 7 1 2 33328 8989
0 8991 7 1 2 35445 8990
0 8992 5 1 1 8991
0 8993 7 1 2 8987 8992
0 8994 5 1 1 8993
0 8995 7 1 2 8980 8994
0 8996 5 1 1 8995
0 8997 7 2 2 23413 30405
0 8998 7 1 2 29534 35448
0 8999 5 1 1 8998
0 9000 7 2 2 25373 29519
0 9001 7 1 2 30380 35450
0 9002 5 1 1 9001
0 9003 7 1 2 8999 9002
0 9004 5 1 1 9003
0 9005 7 1 2 24584 9004
0 9006 5 1 1 9005
0 9007 7 3 2 22610 30081
0 9008 7 1 2 35451 35452
0 9009 5 1 1 9008
0 9010 7 1 2 9006 9009
0 9011 5 1 1 9010
0 9012 7 1 2 28852 35442
0 9013 5 1 1 9012
0 9014 7 4 2 23111 25536
0 9015 7 2 2 35455 29190
0 9016 5 1 1 35459
0 9017 7 1 2 30167 35460
0 9018 5 1 1 9017
0 9019 7 1 2 9013 9018
0 9020 5 1 1 9019
0 9021 7 1 2 9011 9020
0 9022 5 1 1 9021
0 9023 7 3 2 28095 31012
0 9024 5 1 1 35461
0 9025 7 3 2 24585 32243
0 9026 5 1 1 35464
0 9027 7 1 2 9024 9026
0 9028 5 6 1 9027
0 9029 7 2 2 32202 33552
0 9030 5 2 1 35473
0 9031 7 1 2 35475 33019
0 9032 5 1 1 9031
0 9033 7 1 2 29108 9032
0 9034 7 1 2 35467 9033
0 9035 5 1 1 9034
0 9036 7 1 2 9022 9035
0 9037 7 1 2 8996 9036
0 9038 7 1 2 8974 9037
0 9039 5 1 1 9038
0 9040 7 1 2 23923 9039
0 9041 5 1 1 9040
0 9042 7 1 2 31013 33017
0 9043 5 1 1 9042
0 9044 7 1 2 30706 35434
0 9045 7 1 2 34022 9044
0 9046 5 1 1 9045
0 9047 7 1 2 9043 9046
0 9048 5 1 1 9047
0 9049 7 1 2 29109 9048
0 9050 5 1 1 9049
0 9051 7 1 2 26453 30959
0 9052 5 1 1 9051
0 9053 7 1 2 24014 35437
0 9054 5 1 1 9053
0 9055 7 1 2 9052 9054
0 9056 5 1 1 9055
0 9057 7 1 2 24682 9056
0 9058 5 1 1 9057
0 9059 7 1 2 25374 30002
0 9060 7 1 2 30296 9059
0 9061 5 1 1 9060
0 9062 7 1 2 9058 9061
0 9063 5 1 1 9062
0 9064 7 2 2 24187 26754
0 9065 5 2 1 35477
0 9066 7 1 2 35479 35274
0 9067 7 1 2 9063 9066
0 9068 5 1 1 9067
0 9069 7 1 2 9050 9068
0 9070 5 1 1 9069
0 9071 7 1 2 35403 9070
0 9072 5 1 1 9071
0 9073 7 1 2 9041 9072
0 9074 5 1 1 9073
0 9075 7 1 2 28985 9074
0 9076 5 1 1 9075
0 9077 7 3 2 23924 32354
0 9078 7 1 2 22943 33424
0 9079 5 1 1 9078
0 9080 7 1 2 31782 9079
0 9081 5 5 1 9080
0 9082 7 2 2 25988 35484
0 9083 7 1 2 35489 33209
0 9084 5 1 1 9083
0 9085 7 1 2 31783 6843
0 9086 5 3 1 9085
0 9087 7 2 2 28853 35491
0 9088 5 1 1 35494
0 9089 7 1 2 9084 9088
0 9090 5 1 1 9089
0 9091 7 1 2 35481 9090
0 9092 5 1 1 9091
0 9093 7 2 2 30506 35492
0 9094 5 1 1 35496
0 9095 7 1 2 35485 35404
0 9096 5 1 1 9095
0 9097 7 1 2 9094 9096
0 9098 5 1 1 9097
0 9099 7 1 2 27698 9098
0 9100 5 1 1 9099
0 9101 7 1 2 30870 33329
0 9102 7 1 2 35490 9101
0 9103 5 1 1 9102
0 9104 7 1 2 9100 9103
0 9105 5 1 1 9104
0 9106 7 1 2 28727 9105
0 9107 5 1 1 9106
0 9108 7 1 2 28672 26892
0 9109 7 1 2 33330 9108
0 9110 7 1 2 32598 9109
0 9111 7 1 2 35486 9110
0 9112 5 1 1 9111
0 9113 7 1 2 9107 9112
0 9114 7 1 2 9092 9113
0 9115 5 1 1 9114
0 9116 7 1 2 31474 9115
0 9117 5 1 1 9116
0 9118 7 3 2 30209 29737
0 9119 7 1 2 26743 27635
0 9120 7 1 2 35498 9119
0 9121 7 1 2 31435 9120
0 9122 5 1 1 9121
0 9123 7 1 2 9117 9122
0 9124 7 1 2 9076 9123
0 9125 7 1 2 8952 9124
0 9126 5 1 1 9125
0 9127 7 1 2 26314 9126
0 9128 5 1 1 9127
0 9129 7 2 2 24764 32723
0 9130 5 1 1 35501
0 9131 7 2 2 28965 26454
0 9132 5 1 1 35503
0 9133 7 1 2 9130 9132
0 9134 5 6 1 9133
0 9135 7 1 2 35505 35468
0 9136 5 1 1 9135
0 9137 7 4 2 22944 23471
0 9138 5 1 1 35511
0 9139 7 4 2 23544 35512
0 9140 7 1 2 32096 28831
0 9141 7 2 2 35515 9140
0 9142 5 1 1 35519
0 9143 7 1 2 25298 35520
0 9144 5 1 1 9143
0 9145 7 1 2 9136 9144
0 9146 5 1 1 9145
0 9147 7 1 2 26244 28546
0 9148 7 1 2 32696 9147
0 9149 7 1 2 9146 9148
0 9150 5 1 1 9149
0 9151 7 1 2 9128 9150
0 9152 5 1 1 9151
0 9153 7 1 2 23624 9152
0 9154 5 1 1 9153
0 9155 7 1 2 26915 30306
0 9156 7 1 2 32207 9155
0 9157 5 1 1 9156
0 9158 7 1 2 32794 35438
0 9159 5 1 1 9158
0 9160 7 1 2 26997 29538
0 9161 5 1 1 9160
0 9162 7 1 2 9159 9161
0 9163 7 1 2 9157 9162
0 9164 5 1 1 9163
0 9165 7 1 2 26156 9164
0 9166 5 1 1 9165
0 9167 7 1 2 30307 30367
0 9168 7 1 2 34023 9167
0 9169 5 1 1 9168
0 9170 7 1 2 9166 9169
0 9171 5 1 1 9170
0 9172 7 1 2 25299 9171
0 9173 5 1 1 9172
0 9174 7 1 2 32228 30029
0 9175 7 1 2 35499 9174
0 9176 5 1 1 9175
0 9177 7 1 2 9173 9176
0 9178 5 1 1 9177
0 9179 7 1 2 24586 9178
0 9180 5 1 1 9179
0 9181 7 1 2 31014 35453
0 9182 7 1 2 35500 9181
0 9183 5 1 1 9182
0 9184 7 1 2 9180 9183
0 9185 5 1 1 9184
0 9186 7 1 2 27582 9185
0 9187 5 1 1 9186
0 9188 7 2 2 22945 34784
0 9189 5 2 1 35521
0 9190 7 1 2 26388 32203
0 9191 5 1 1 9190
0 9192 7 1 2 35523 9191
0 9193 5 3 1 9192
0 9194 7 1 2 35525 35469
0 9195 5 1 1 9194
0 9196 7 2 2 29894 29664
0 9197 7 1 2 35528 32146
0 9198 5 1 1 9197
0 9199 7 1 2 9195 9198
0 9200 5 1 1 9199
0 9201 7 1 2 23925 28587
0 9202 7 1 2 9200 9201
0 9203 5 1 1 9202
0 9204 7 1 2 9187 9203
0 9205 5 1 1 9204
0 9206 7 1 2 25537 9205
0 9207 5 1 1 9206
0 9208 7 1 2 25375 29987
0 9209 5 1 1 9208
0 9210 7 1 2 4019 9209
0 9211 5 1 1 9210
0 9212 7 1 2 24683 9211
0 9213 5 1 1 9212
0 9214 7 3 2 29955 29524
0 9215 5 1 1 35530
0 9216 7 1 2 32150 35531
0 9217 5 1 1 9216
0 9218 7 1 2 9213 9217
0 9219 5 1 1 9218
0 9220 7 1 2 28139 9219
0 9221 5 1 1 9220
0 9222 7 1 2 27753 30422
0 9223 5 1 1 9222
0 9224 7 1 2 9221 9223
0 9225 5 1 1 9224
0 9226 7 5 2 23926 28891
0 9227 7 1 2 35533 28547
0 9228 7 1 2 9225 9227
0 9229 5 1 1 9228
0 9230 7 1 2 9207 9229
0 9231 5 1 1 9230
0 9232 7 1 2 28986 9231
0 9233 5 1 1 9232
0 9234 7 1 2 23112 35497
0 9235 5 1 1 9234
0 9236 7 4 2 25538 27583
0 9237 7 5 2 25894 35538
0 9238 7 1 2 25300 27364
0 9239 7 1 2 35542 9238
0 9240 5 1 1 9239
0 9241 7 1 2 9235 9240
0 9242 5 1 1 9241
0 9243 7 1 2 27699 9242
0 9244 5 1 1 9243
0 9245 7 3 2 24587 28759
0 9246 7 5 2 25539 23927
0 9247 7 2 2 35547 35550
0 9248 7 1 2 27584 32361
0 9249 7 1 2 35555 9248
0 9250 5 1 1 9249
0 9251 7 1 2 9244 9250
0 9252 5 1 1 9251
0 9253 7 1 2 28728 9252
0 9254 5 1 1 9253
0 9255 7 2 2 25301 27585
0 9256 7 1 2 25540 35353
0 9257 7 1 2 35557 9256
0 9258 7 2 2 32957 9257
0 9259 7 1 2 27653 35559
0 9260 5 1 1 9259
0 9261 7 6 2 25541 25989
0 9262 7 1 2 27666 35561
0 9263 5 1 1 9262
0 9264 7 1 2 23113 35495
0 9265 5 1 1 9264
0 9266 7 1 2 9263 9265
0 9267 5 1 1 9266
0 9268 7 1 2 35482 9267
0 9269 5 1 1 9268
0 9270 7 1 2 9260 9269
0 9271 7 1 2 9254 9270
0 9272 5 1 1 9271
0 9273 7 1 2 31475 9272
0 9274 5 1 1 9273
0 9275 7 1 2 23114 35401
0 9276 5 1 1 9275
0 9277 7 1 2 28309 31228
0 9278 7 1 2 35543 9277
0 9279 5 1 1 9278
0 9280 7 1 2 9276 9279
0 9281 5 1 1 9280
0 9282 7 1 2 27700 9281
0 9283 5 1 1 9282
0 9284 7 2 2 27595 31229
0 9285 7 1 2 35556 35567
0 9286 5 1 1 9285
0 9287 7 1 2 9283 9286
0 9288 5 1 1 9287
0 9289 7 1 2 28729 9288
0 9290 5 1 1 9289
0 9291 7 1 2 35398 30186
0 9292 5 1 1 9291
0 9293 7 1 2 24684 25542
0 9294 7 1 2 35568 9293
0 9295 5 1 1 9294
0 9296 7 1 2 9292 9295
0 9297 5 1 1 9296
0 9298 7 1 2 35483 9297
0 9299 5 1 1 9298
0 9300 7 1 2 25435 31230
0 9301 7 1 2 35560 9300
0 9302 5 1 1 9301
0 9303 7 1 2 9299 9302
0 9304 7 1 2 9290 9303
0 9305 5 1 1 9304
0 9306 7 1 2 28648 9305
0 9307 5 1 1 9306
0 9308 7 1 2 9274 9307
0 9309 7 1 2 9233 9308
0 9310 7 1 2 9154 9309
0 9311 5 1 1 9310
0 9312 7 1 2 35334 28940
0 9313 7 1 2 9311 9312
0 9314 5 1 1 9313
0 9315 7 1 2 31193 29775
0 9316 7 1 2 33048 9315
0 9317 5 1 1 9316
0 9318 7 1 2 28340 30072
0 9319 7 1 2 33339 9318
0 9320 7 1 2 35280 9319
0 9321 5 1 1 9320
0 9322 7 1 2 9317 9321
0 9323 7 2 2 23696 30617
0 9324 7 1 2 33835 35569
0 9325 5 1 1 9324
0 9326 7 1 2 30073 34759
0 9327 5 1 1 9326
0 9328 7 1 2 9325 9327
0 9329 5 1 1 9328
0 9330 7 1 2 24452 9329
0 9331 5 1 1 9330
0 9332 7 2 2 22445 29757
0 9333 7 4 2 25220 23697
0 9334 7 1 2 31037 35573
0 9335 7 1 2 35571 9334
0 9336 5 1 1 9335
0 9337 7 1 2 9331 9336
0 9338 5 1 1 9337
0 9339 7 1 2 28823 9338
0 9340 5 1 1 9339
0 9341 7 1 2 29776 30659
0 9342 5 1 1 9341
0 9343 7 2 2 34739 34422
0 9344 7 1 2 23928 35577
0 9345 5 1 1 9344
0 9346 7 1 2 9342 9345
0 9347 5 1 1 9346
0 9348 7 1 2 24453 9347
0 9349 5 1 1 9348
0 9350 7 1 2 29758 27922
0 9351 7 1 2 29937 9350
0 9352 5 1 1 9351
0 9353 7 1 2 9349 9352
0 9354 5 1 1 9353
0 9355 7 1 2 28730 28140
0 9356 7 1 2 9354 9355
0 9357 5 1 1 9356
0 9358 7 1 2 9340 9357
0 9359 7 1 2 9322 9358
0 9360 5 1 1 9359
0 9361 7 1 2 26075 9360
0 9362 5 1 1 9361
0 9363 7 2 2 27754 28768
0 9364 7 1 2 24588 35579
0 9365 5 1 1 9364
0 9366 7 1 2 6072 9365
0 9367 5 1 1 9366
0 9368 7 2 2 28987 30702
0 9369 7 1 2 29698 35581
0 9370 7 1 2 9367 9369
0 9371 5 1 1 9370
0 9372 7 1 2 9362 9371
0 9373 5 1 1 9372
0 9374 7 1 2 29110 29543
0 9375 7 1 2 9373 9374
0 9376 5 1 1 9375
0 9377 7 1 2 26839 35127
0 9378 7 2 2 30810 9377
0 9379 5 1 1 35583
0 9380 7 1 2 34936 26873
0 9381 5 1 1 9380
0 9382 7 1 2 33808 9381
0 9383 5 7 1 9382
0 9384 7 1 2 32097 35585
0 9385 5 1 1 9384
0 9386 7 1 2 9379 9385
0 9387 5 1 1 9386
0 9388 7 1 2 29160 9387
0 9389 5 1 1 9388
0 9390 7 1 2 27313 34124
0 9391 5 1 1 9390
0 9392 7 1 2 22446 31162
0 9393 5 1 1 9392
0 9394 7 1 2 24454 31834
0 9395 5 1 1 9394
0 9396 7 1 2 9393 9395
0 9397 5 5 1 9396
0 9398 7 1 2 34135 35592
0 9399 5 1 1 9398
0 9400 7 1 2 9391 9399
0 9401 5 1 1 9400
0 9402 7 2 2 32443 26845
0 9403 5 1 1 35597
0 9404 7 1 2 34990 9403
0 9405 5 3 1 9404
0 9406 7 1 2 9401 35599
0 9407 5 1 1 9406
0 9408 7 1 2 34611 33932
0 9409 5 1 1 9408
0 9410 7 1 2 28790 26846
0 9411 7 1 2 29304 9410
0 9412 5 1 1 9411
0 9413 7 1 2 9409 9412
0 9414 5 1 1 9413
0 9415 7 1 2 23929 28379
0 9416 7 1 2 9414 9415
0 9417 5 1 1 9416
0 9418 7 1 2 9407 9417
0 9419 7 1 2 9389 9418
0 9420 5 1 1 9419
0 9421 7 1 2 23698 30181
0 9422 7 1 2 9420 9421
0 9423 5 1 1 9422
0 9424 7 1 2 9376 9423
0 9425 5 1 1 9424
0 9426 7 1 2 29279 9425
0 9427 5 1 1 9426
0 9428 7 2 2 26315 33844
0 9429 7 2 2 28207 35602
0 9430 5 1 1 35604
0 9431 7 1 2 29714 33098
0 9432 5 1 1 9431
0 9433 7 1 2 9430 9432
0 9434 5 1 1 9433
0 9435 7 1 2 32925 9434
0 9436 5 1 1 9435
0 9437 7 3 2 22447 22825
0 9438 7 1 2 26076 31067
0 9439 7 1 2 35606 9438
0 9440 7 1 2 34729 9439
0 9441 5 1 1 9440
0 9442 7 1 2 9436 9441
0 9443 5 1 1 9442
0 9444 7 1 2 23625 9443
0 9445 5 1 1 9444
0 9446 7 2 2 26316 29759
0 9447 7 1 2 24765 27672
0 9448 7 1 2 35609 9447
0 9449 7 1 2 33091 9448
0 9450 5 1 1 9449
0 9451 7 1 2 9445 9450
0 9452 5 1 1 9451
0 9453 7 1 2 24267 9452
0 9454 5 1 1 9453
0 9455 7 4 2 25623 24015
0 9456 7 2 2 22611 35611
0 9457 7 1 2 25895 32758
0 9458 7 1 2 35615 9457
0 9459 7 1 2 29927 9458
0 9460 5 1 1 9459
0 9461 7 1 2 9454 9460
0 9462 5 1 1 9461
0 9463 7 1 2 23699 9462
0 9464 5 1 1 9463
0 9465 7 1 2 24016 31935
0 9466 7 3 2 29544 9465
0 9467 7 3 2 25221 29604
0 9468 7 1 2 32759 35620
0 9469 7 1 2 35617 9468
0 9470 5 1 1 9469
0 9471 7 1 2 9464 9470
0 9472 5 1 1 9471
0 9473 7 1 2 32244 9472
0 9474 5 1 1 9473
0 9475 7 1 2 32760 35462
0 9476 5 1 1 9475
0 9477 7 1 2 8636 9476
0 9478 5 1 1 9477
0 9479 7 1 2 28941 35618
0 9480 7 1 2 9478 9479
0 9481 5 1 1 9480
0 9482 7 1 2 9474 9481
0 9483 5 1 1 9482
0 9484 7 1 2 32724 9483
0 9485 5 1 1 9484
0 9486 7 1 2 31632 32931
0 9487 5 2 1 9486
0 9488 7 1 2 31662 32926
0 9489 5 1 1 9488
0 9490 7 1 2 35623 9489
0 9491 5 1 1 9490
0 9492 7 1 2 26411 9491
0 9493 5 1 1 9492
0 9494 7 1 2 24589 27646
0 9495 7 1 2 30308 9494
0 9496 7 1 2 35359 9495
0 9497 5 1 1 9496
0 9498 7 1 2 9493 9497
0 9499 5 1 1 9498
0 9500 7 1 2 33323 9499
0 9501 5 1 1 9500
0 9502 7 1 2 28208 32873
0 9503 7 1 2 30507 9502
0 9504 5 1 1 9503
0 9505 7 1 2 32887 9504
0 9506 5 1 1 9505
0 9507 7 1 2 26412 9506
0 9508 5 1 1 9507
0 9509 7 1 2 22826 29788
0 9510 7 1 2 30352 9509
0 9511 5 1 1 9510
0 9512 7 1 2 9508 9511
0 9513 5 1 1 9512
0 9514 7 1 2 32098 9513
0 9515 5 1 1 9514
0 9516 7 1 2 9501 9515
0 9517 5 1 1 9516
0 9518 7 1 2 24268 9517
0 9519 5 1 1 9518
0 9520 7 2 2 29871 35113
0 9521 7 1 2 25624 28832
0 9522 7 1 2 35625 9521
0 9523 7 1 2 33324 9522
0 9524 5 1 1 9523
0 9525 7 1 2 9519 9524
0 9526 5 1 1 9525
0 9527 7 1 2 32725 9526
0 9528 5 1 1 9527
0 9529 7 3 2 24100 26317
0 9530 7 3 2 23626 35627
0 9531 7 1 2 35630 27775
0 9532 5 1 1 9531
0 9533 7 3 2 23930 32577
0 9534 7 2 2 22612 35633
0 9535 5 1 1 35636
0 9536 7 1 2 26413 35637
0 9537 5 1 1 9536
0 9538 7 1 2 27409 27394
0 9539 7 1 2 29789 9538
0 9540 5 1 1 9539
0 9541 7 1 2 9537 9540
0 9542 5 1 1 9541
0 9543 7 1 2 33141 9542
0 9544 5 1 1 9543
0 9545 7 1 2 9532 9544
0 9546 5 1 1 9545
0 9547 7 1 2 24269 9546
0 9548 5 1 1 9547
0 9549 7 1 2 35128 28919
0 9550 7 1 2 35626 9549
0 9551 5 1 1 9550
0 9552 7 1 2 9548 9551
0 9553 5 1 1 9552
0 9554 7 1 2 33113 9553
0 9555 5 1 1 9554
0 9556 7 1 2 29161 34795
0 9557 5 1 1 9556
0 9558 7 1 2 30318 34798
0 9559 5 1 1 9558
0 9560 7 1 2 9557 9559
0 9561 5 2 1 9560
0 9562 7 1 2 26947 26658
0 9563 7 1 2 35006 9562
0 9564 7 1 2 35638 9563
0 9565 5 1 1 9564
0 9566 7 1 2 9555 9565
0 9567 7 1 2 9528 9566
0 9568 5 1 1 9567
0 9569 7 1 2 23700 9568
0 9570 5 1 1 9569
0 9571 7 6 2 23627 24270
0 9572 5 1 1 35640
0 9573 7 1 2 30813 33356
0 9574 5 1 1 9573
0 9575 7 1 2 32795 33142
0 9576 5 1 1 9575
0 9577 7 1 2 9574 9576
0 9578 5 1 1 9577
0 9579 7 1 2 35641 9578
0 9580 5 1 1 9579
0 9581 7 1 2 26077 27338
0 9582 7 1 2 30498 9581
0 9583 5 1 1 9582
0 9584 7 1 2 9580 9583
0 9585 5 1 1 9584
0 9586 7 1 2 29162 9585
0 9587 5 1 1 9586
0 9588 7 2 2 24271 33067
0 9589 7 1 2 3962 32941
0 9590 5 1 1 9589
0 9591 7 2 2 22448 30618
0 9592 7 1 2 23628 31120
0 9593 7 1 2 35648 9592
0 9594 5 1 1 9593
0 9595 7 1 2 9590 9594
0 9596 5 1 1 9595
0 9597 7 1 2 35646 9596
0 9598 5 1 1 9597
0 9599 7 1 2 9587 9598
0 9600 5 1 1 9599
0 9601 7 1 2 26318 9600
0 9602 5 1 1 9601
0 9603 7 4 2 23115 25896
0 9604 7 1 2 35650 28769
0 9605 7 1 2 35642 9604
0 9606 7 1 2 27967 9605
0 9607 7 1 2 33068 9606
0 9608 5 1 1 9607
0 9609 7 1 2 9602 9608
0 9610 5 1 1 9609
0 9611 7 1 2 23701 9610
0 9612 5 1 1 9611
0 9613 7 2 2 24685 31121
0 9614 7 1 2 29699 35654
0 9615 7 1 2 29545 9614
0 9616 7 1 2 35647 9615
0 9617 5 1 1 9616
0 9618 7 1 2 9612 9617
0 9619 5 1 1 9618
0 9620 7 1 2 33056 9619
0 9621 5 1 1 9620
0 9622 7 2 2 24766 25625
0 9623 7 2 2 26078 35656
0 9624 5 1 1 35658
0 9625 7 1 2 32521 35643
0 9626 5 1 1 9625
0 9627 7 1 2 9624 9626
0 9628 5 1 1 9627
0 9629 7 1 2 33351 9628
0 9630 5 1 1 9629
0 9631 7 1 2 32545 31998
0 9632 7 1 2 30415 9631
0 9633 5 1 1 9632
0 9634 7 1 2 9630 9633
0 9635 5 1 1 9634
0 9636 7 1 2 33099 9635
0 9637 5 1 1 9636
0 9638 7 1 2 35605 35644
0 9639 7 1 2 33103 9638
0 9640 5 1 1 9639
0 9641 7 1 2 9637 9640
0 9642 5 1 1 9641
0 9643 7 1 2 23702 9642
0 9644 5 1 1 9643
0 9645 7 2 2 32546 35619
0 9646 7 1 2 30074 29605
0 9647 7 1 2 35660 9646
0 9648 5 1 1 9647
0 9649 7 1 2 9644 9648
0 9650 5 1 1 9649
0 9651 7 1 2 32653 9650
0 9652 5 1 1 9651
0 9653 7 1 2 28341 32623
0 9654 7 1 2 30084 9653
0 9655 7 1 2 35661 9654
0 9656 5 1 1 9655
0 9657 7 1 2 9652 9656
0 9658 7 1 2 9621 9657
0 9659 7 1 2 9570 9658
0 9660 7 1 2 9485 9659
0 9661 5 1 1 9660
0 9662 7 1 2 26157 9661
0 9663 5 1 1 9662
0 9664 7 1 2 9427 9663
0 9665 5 1 1 9664
0 9666 7 1 2 34072 9665
0 9667 5 1 1 9666
0 9668 7 1 2 25302 33531
0 9669 7 1 2 29546 9668
0 9670 5 1 1 9669
0 9671 7 1 2 25070 28746
0 9672 7 1 2 33461 9671
0 9673 5 1 1 9672
0 9674 7 1 2 9670 9673
0 9675 5 1 1 9674
0 9676 7 1 2 24590 9675
0 9677 5 1 1 9676
0 9678 7 5 2 24017 30707
0 9679 7 2 2 28486 35662
0 9680 7 1 2 28096 35667
0 9681 5 1 1 9680
0 9682 7 1 2 9677 9681
0 9683 5 1 1 9682
0 9684 7 1 2 25490 9683
0 9685 5 1 1 9684
0 9686 7 2 2 27523 33446
0 9687 7 1 2 28310 35669
0 9688 7 1 2 29547 9687
0 9689 5 1 1 9688
0 9690 7 1 2 9685 9689
0 9691 5 1 1 9690
0 9692 7 1 2 23259 9691
0 9693 5 1 1 9692
0 9694 7 3 2 25222 30335
0 9695 7 1 2 26802 28234
0 9696 7 1 2 35671 9695
0 9697 7 1 2 29548 9696
0 9698 5 1 1 9697
0 9699 7 1 2 9693 9698
0 9700 5 1 1 9699
0 9701 7 1 2 33553 9700
0 9702 5 1 1 9701
0 9703 7 6 2 25990 26245
0 9704 7 1 2 23040 35674
0 9705 7 2 2 31476 9704
0 9706 7 2 2 29225 29549
0 9707 7 1 2 35680 35682
0 9708 5 1 1 9707
0 9709 7 1 2 9702 9708
0 9710 5 1 1 9709
0 9711 7 1 2 24875 9710
0 9712 5 1 1 9711
0 9713 7 1 2 26787 35440
0 9714 5 1 1 9713
0 9715 7 2 2 35040 9714
0 9716 7 1 2 24101 35684
0 9717 5 1 1 9716
0 9718 7 5 2 25543 26079
0 9719 7 2 2 24188 35686
0 9720 7 1 2 29033 35691
0 9721 5 1 1 9720
0 9722 7 1 2 9717 9721
0 9723 5 1 1 9722
0 9724 7 2 2 32362 9723
0 9725 7 1 2 35693 35683
0 9726 5 1 1 9725
0 9727 7 1 2 9712 9726
0 9728 5 1 1 9727
0 9729 7 1 2 22449 9728
0 9730 5 1 1 9729
0 9731 7 1 2 31477 35493
0 9732 5 1 1 9731
0 9733 7 1 2 28649 35399
0 9734 5 1 1 9733
0 9735 7 1 2 9732 9734
0 9736 5 1 1 9735
0 9737 7 2 2 23260 31090
0 9738 7 1 2 28342 35695
0 9739 7 1 2 29550 9738
0 9740 7 1 2 9736 9739
0 9741 5 1 1 9740
0 9742 7 1 2 9730 9741
0 9743 5 1 1 9742
0 9744 7 1 2 31793 9743
0 9745 5 1 1 9744
0 9746 7 1 2 22946 35685
0 9747 5 1 1 9746
0 9748 7 1 2 28508 31778
0 9749 5 1 1 9748
0 9750 7 1 2 9747 9749
0 9751 5 1 1 9750
0 9752 7 4 2 30319 29551
0 9753 7 1 2 30336 35697
0 9754 7 1 2 9751 9753
0 9755 5 1 1 9754
0 9756 7 2 2 26744 31079
0 9757 5 1 1 35701
0 9758 7 2 2 24876 29191
0 9759 7 1 2 25071 35703
0 9760 5 1 1 9759
0 9761 7 3 2 26803 30830
0 9762 5 1 1 35705
0 9763 7 1 2 29656 9762
0 9764 7 1 2 9760 9763
0 9765 5 1 1 9764
0 9766 7 1 2 24965 9765
0 9767 5 1 1 9766
0 9768 7 1 2 9757 9767
0 9769 5 1 1 9768
0 9770 7 1 2 35631 9769
0 9771 5 1 1 9770
0 9772 7 3 2 25491 26080
0 9773 7 3 2 24877 35708
0 9774 5 1 1 35711
0 9775 7 2 2 29280 27806
0 9776 7 1 2 35712 35714
0 9777 5 1 1 9776
0 9778 7 1 2 9771 9777
0 9779 5 1 1 9778
0 9780 7 1 2 25544 9779
0 9781 5 1 1 9780
0 9782 7 1 2 35288 28413
0 9783 7 1 2 30221 9782
0 9784 5 1 1 9783
0 9785 7 1 2 9781 9784
0 9786 5 1 1 9785
0 9787 7 1 2 24018 29163
0 9788 7 1 2 9786 9787
0 9789 5 1 1 9788
0 9790 7 1 2 9755 9789
0 9791 5 1 1 9790
0 9792 7 1 2 32099 9791
0 9793 5 1 1 9792
0 9794 7 1 2 28673 33293
0 9795 5 1 1 9794
0 9796 7 1 2 32906 9795
0 9797 5 1 1 9796
0 9798 7 1 2 29830 35715
0 9799 5 1 1 9798
0 9800 7 1 2 749 30594
0 9801 5 1 1 9800
0 9802 7 1 2 9801 30282
0 9803 5 1 1 9802
0 9804 7 1 2 9799 9803
0 9805 5 1 1 9804
0 9806 7 1 2 25545 9805
0 9807 5 1 1 9806
0 9808 7 3 2 22947 29872
0 9809 7 1 2 33071 35716
0 9810 5 1 1 9809
0 9811 7 5 2 26158 29873
0 9812 7 1 2 28548 35719
0 9813 5 1 1 9812
0 9814 7 1 2 35476 9813
0 9815 5 2 1 9814
0 9816 7 1 2 24878 35724
0 9817 5 1 1 9816
0 9818 7 1 2 9810 9817
0 9819 7 1 2 9807 9818
0 9820 5 1 1 9819
0 9821 7 1 2 23629 9820
0 9822 5 1 1 9821
0 9823 7 2 2 30468 29843
0 9824 5 1 1 35726
0 9825 7 1 2 35038 35727
0 9826 5 1 1 9825
0 9827 7 1 2 30847 35474
0 9828 5 1 1 9827
0 9829 7 1 2 9826 9828
0 9830 7 1 2 9822 9829
0 9831 5 1 1 9830
0 9832 7 1 2 23545 9831
0 9833 5 1 1 9832
0 9834 7 2 2 24879 35443
0 9835 5 1 1 35728
0 9836 7 1 2 24189 34591
0 9837 5 1 1 9836
0 9838 7 1 2 9835 9837
0 9839 5 1 1 9838
0 9840 7 1 2 29839 9839
0 9841 5 1 1 9840
0 9842 7 1 2 22948 35725
0 9843 5 1 1 9842
0 9844 7 1 2 29831 35729
0 9845 5 1 1 9844
0 9846 7 1 2 9843 9845
0 9847 5 1 1 9846
0 9848 7 1 2 25492 9847
0 9849 5 1 1 9848
0 9850 7 2 2 26246 35717
0 9851 7 1 2 35730 35042
0 9852 5 1 1 9851
0 9853 7 1 2 9849 9852
0 9854 5 1 1 9853
0 9855 7 1 2 23630 9854
0 9856 5 1 1 9855
0 9857 7 1 2 9841 9856
0 9858 7 1 2 9833 9857
0 9859 5 1 1 9858
0 9860 7 1 2 26319 9859
0 9861 5 1 1 9860
0 9862 7 1 2 28650 33554
0 9863 5 1 1 9862
0 9864 7 1 2 32280 9863
0 9865 5 1 1 9864
0 9866 7 1 2 24880 9865
0 9867 5 1 1 9866
0 9868 7 1 2 29653 33555
0 9869 5 1 1 9868
0 9870 7 1 2 9867 9869
0 9871 5 1 1 9870
0 9872 7 1 2 29832 26701
0 9873 7 1 2 9871 9872
0 9874 5 1 1 9873
0 9875 7 1 2 9861 9874
0 9876 5 1 1 9875
0 9877 7 1 2 9797 9876
0 9878 5 1 1 9877
0 9879 7 1 2 9793 9878
0 9880 5 1 1 9879
0 9881 7 1 2 28988 9880
0 9882 5 1 1 9881
0 9883 7 6 2 26159 26514
0 9884 5 1 1 35732
0 9885 7 3 2 26081 35733
0 9886 7 1 2 30413 32889
0 9887 7 2 2 35738 9886
0 9888 5 1 1 35741
0 9889 7 1 2 25223 35742
0 9890 5 1 1 9889
0 9891 7 1 2 29226 35668
0 9892 5 1 1 9891
0 9893 7 1 2 9890 9892
0 9894 5 1 1 9893
0 9895 7 1 2 22450 9894
0 9896 5 1 1 9895
0 9897 7 1 2 34358 34643
0 9898 5 1 1 9897
0 9899 7 1 2 9888 9898
0 9900 5 1 1 9899
0 9901 7 1 2 27908 9900
0 9902 5 1 1 9901
0 9903 7 1 2 9896 9902
0 9904 5 1 1 9903
0 9905 7 1 2 25493 9904
0 9906 5 1 1 9905
0 9907 7 1 2 35698 35670
0 9908 5 1 1 9907
0 9909 7 1 2 9906 9908
0 9910 5 1 1 9909
0 9911 7 1 2 33556 9910
0 9912 5 1 1 9911
0 9913 7 1 2 35699 35681
0 9914 5 1 1 9913
0 9915 7 1 2 9912 9914
0 9916 5 1 1 9915
0 9917 7 1 2 24881 9916
0 9918 5 1 1 9917
0 9919 7 1 2 35700 35694
0 9920 5 1 1 9919
0 9921 7 1 2 9918 9920
0 9922 5 1 1 9921
0 9923 7 1 2 31406 9922
0 9924 5 1 1 9923
0 9925 7 5 2 25546 29281
0 9926 7 1 2 29034 30253
0 9927 7 2 2 35743 9926
0 9928 7 1 2 29833 35748
0 9929 5 1 1 9928
0 9930 7 1 2 23631 35702
0 9931 5 1 1 9930
0 9932 7 1 2 24882 26707
0 9933 5 3 1 9932
0 9934 7 1 2 1183 35750
0 9935 5 1 1 9934
0 9936 7 1 2 29192 9935
0 9937 5 1 1 9936
0 9938 7 1 2 28663 35706
0 9939 5 1 1 9938
0 9940 7 1 2 26539 30102
0 9941 5 1 1 9940
0 9942 7 1 2 9939 9941
0 9943 7 1 2 9937 9942
0 9944 5 1 1 9943
0 9945 7 1 2 24966 9944
0 9946 5 1 1 9945
0 9947 7 1 2 9931 9946
0 9948 5 1 1 9947
0 9949 7 1 2 25547 9948
0 9950 5 1 1 9949
0 9951 7 5 2 23632 26160
0 9952 5 1 1 35753
0 9953 7 1 2 26455 9952
0 9954 7 1 2 35207 9953
0 9955 7 1 2 35480 9954
0 9956 5 1 1 9955
0 9957 7 1 2 26082 9956
0 9958 7 1 2 9950 9957
0 9959 5 1 1 9958
0 9960 7 1 2 22949 35444
0 9961 5 1 1 9960
0 9962 7 1 2 23041 35070
0 9963 5 1 1 9962
0 9964 7 1 2 9961 9963
0 9965 5 1 1 9964
0 9966 7 1 2 23546 9965
0 9967 5 1 1 9966
0 9968 7 1 2 26782 35176
0 9969 5 1 1 9968
0 9970 7 1 2 9967 9969
0 9971 5 1 1 9970
0 9972 7 1 2 23633 9971
0 9973 5 1 1 9972
0 9974 7 1 2 24102 9973
0 9975 5 1 1 9974
0 9976 7 1 2 31068 9975
0 9977 7 1 2 9959 9976
0 9978 5 1 1 9977
0 9979 7 1 2 9929 9978
0 9980 5 1 1 9979
0 9981 7 1 2 35639 9980
0 9982 5 1 1 9981
0 9983 7 1 2 25897 9982
0 9984 7 1 2 9924 9983
0 9985 7 1 2 9882 9984
0 9986 7 1 2 9745 9985
0 9987 5 1 1 9986
0 9988 7 1 2 25224 28923
0 9989 5 1 1 9988
0 9990 7 1 2 5143 9989
0 9991 5 5 1 9990
0 9992 7 1 2 22728 35758
0 9993 5 1 1 9992
0 9994 7 1 2 27081 30626
0 9995 5 1 1 9994
0 9996 7 1 2 9993 9995
0 9997 5 1 1 9996
0 9998 7 1 2 22613 9997
0 9999 5 1 1 9998
0 10000 7 1 2 22729 33211
0 10001 5 1 1 10000
0 10002 7 1 2 10001 4119
0 10003 5 3 1 10002
0 10004 7 1 2 30646 35763
0 10005 5 1 1 10004
0 10006 7 1 2 9999 10005
0 10007 5 1 1 10006
0 10008 7 1 2 22451 10007
0 10009 5 1 1 10008
0 10010 7 1 2 28401 28343
0 10011 7 2 2 31091 10010
0 10012 5 1 1 35766
0 10013 7 1 2 22730 35767
0 10014 5 1 1 10013
0 10015 7 1 2 10009 10014
0 10016 5 3 1 10015
0 10017 7 1 2 33933 35768
0 10018 5 1 1 10017
0 10019 7 1 2 29164 30941
0 10020 5 1 1 10019
0 10021 7 2 2 24019 30695
0 10022 7 1 2 28141 31134
0 10023 7 1 2 35771 10022
0 10024 5 1 1 10023
0 10025 7 1 2 10020 10024
0 10026 5 2 1 10025
0 10027 7 1 2 33898 35773
0 10028 5 1 1 10027
0 10029 7 1 2 10018 10028
0 10030 5 2 1 10029
0 10031 7 1 2 24883 34909
0 10032 5 1 1 10031
0 10033 7 1 2 24967 35707
0 10034 5 1 1 10033
0 10035 7 1 2 10032 10034
0 10036 5 1 1 10035
0 10037 7 1 2 35775 10036
0 10038 5 1 1 10037
0 10039 7 1 2 22614 35759
0 10040 5 1 1 10039
0 10041 7 1 2 30647 33212
0 10042 5 1 1 10041
0 10043 7 1 2 10040 10042
0 10044 5 1 1 10043
0 10045 7 1 2 22452 10044
0 10046 5 1 1 10045
0 10047 7 1 2 10012 10046
0 10048 5 1 1 10047
0 10049 7 1 2 27133 10048
0 10050 5 1 1 10049
0 10051 7 1 2 34747 27082
0 10052 5 1 1 10051
0 10053 7 1 2 10050 10052
0 10054 5 1 1 10053
0 10055 7 1 2 31478 10054
0 10056 5 1 1 10055
0 10057 7 1 2 34785 32858
0 10058 5 1 1 10057
0 10059 7 1 2 31137 30634
0 10060 5 1 1 10059
0 10061 7 1 2 28076 34631
0 10062 5 1 1 10061
0 10063 7 1 2 10060 10062
0 10064 5 1 1 10063
0 10065 7 1 2 22615 10064
0 10066 5 1 1 10065
0 10067 7 1 2 30648 35376
0 10068 5 1 1 10067
0 10069 7 1 2 10066 10068
0 10070 5 1 1 10069
0 10071 7 1 2 22453 10070
0 10072 5 1 1 10071
0 10073 7 1 2 31001 28367
0 10074 5 1 1 10073
0 10075 7 1 2 10072 10074
0 10076 5 1 1 10075
0 10077 7 1 2 32100 10076
0 10078 5 1 1 10077
0 10079 7 1 2 10058 10078
0 10080 5 1 1 10079
0 10081 7 1 2 28989 10080
0 10082 5 1 1 10081
0 10083 7 1 2 10056 10082
0 10084 5 1 1 10083
0 10085 7 1 2 27501 789
0 10086 7 1 2 4405 10085
0 10087 7 1 2 10084 10086
0 10088 5 1 1 10087
0 10089 7 1 2 10038 10088
0 10090 5 1 1 10089
0 10091 7 1 2 25548 10090
0 10092 5 1 1 10091
0 10093 7 1 2 32485 35774
0 10094 5 1 1 10093
0 10095 7 4 2 24103 26893
0 10096 7 1 2 35769 35777
0 10097 5 1 1 10096
0 10098 7 1 2 10094 10097
0 10099 5 1 1 10098
0 10100 7 1 2 29852 10099
0 10101 5 1 1 10100
0 10102 7 1 2 35776 35118
0 10103 5 1 1 10102
0 10104 7 1 2 10101 10103
0 10105 5 1 1 10104
0 10106 7 1 2 26745 10105
0 10107 5 1 1 10106
0 10108 7 1 2 10092 10107
0 10109 5 1 1 10108
0 10110 7 1 2 26414 10109
0 10111 5 1 1 10110
0 10112 7 1 2 32486 35770
0 10113 5 1 1 10112
0 10114 7 2 2 28915 31038
0 10115 5 1 1 35781
0 10116 7 1 2 2895 10115
0 10117 5 2 1 10116
0 10118 7 1 2 33134 33204
0 10119 7 1 2 35783 10118
0 10120 5 1 1 10119
0 10121 7 1 2 10113 10120
0 10122 5 1 1 10121
0 10123 7 1 2 35749 10122
0 10124 5 1 1 10123
0 10125 7 1 2 23931 10124
0 10126 7 1 2 10111 10125
0 10127 5 1 1 10126
0 10128 7 1 2 23703 10127
0 10129 7 1 2 9987 10128
0 10130 5 1 1 10129
0 10131 7 1 2 9667 10130
0 10132 7 1 2 9314 10131
0 10133 5 1 1 10132
0 10134 7 1 2 25791 10133
0 10135 5 1 1 10134
0 10136 7 1 2 23188 10135
0 10137 7 1 2 8891 10136
0 10138 5 1 1 10137
0 10139 7 1 2 27034 29361
0 10140 5 3 1 10139
0 10141 7 1 2 30733 32415
0 10142 5 1 1 10141
0 10143 7 1 2 35785 10142
0 10144 5 1 1 10143
0 10145 7 1 2 24591 10144
0 10146 5 1 1 10145
0 10147 7 2 2 23801 28097
0 10148 7 1 2 27035 35788
0 10149 5 1 1 10148
0 10150 7 1 2 10146 10149
0 10151 5 1 1 10150
0 10152 7 1 2 25898 10151
0 10153 5 1 1 10152
0 10154 7 1 2 25303 32416
0 10155 5 1 1 10154
0 10156 7 1 2 35786 10155
0 10157 5 2 1 10156
0 10158 7 1 2 31633 35790
0 10159 5 1 1 10158
0 10160 7 1 2 10153 10159
0 10161 5 1 1 10160
0 10162 7 1 2 24686 10161
0 10163 5 1 1 10162
0 10164 7 1 2 28674 33836
0 10165 5 1 1 10164
0 10166 7 1 2 31674 31025
0 10167 5 1 1 10166
0 10168 7 1 2 10165 10167
0 10169 5 1 1 10168
0 10170 7 1 2 31699 10169
0 10171 5 1 1 10170
0 10172 7 1 2 10163 10171
0 10173 5 1 1 10172
0 10174 7 1 2 23261 10173
0 10175 5 1 1 10174
0 10176 7 1 2 24020 31865
0 10177 5 1 1 10176
0 10178 7 1 2 28142 33189
0 10179 5 1 1 10178
0 10180 7 1 2 10177 10179
0 10181 5 1 1 10180
0 10182 7 1 2 35651 10181
0 10183 5 1 1 10182
0 10184 7 1 2 32034 32040
0 10185 5 1 1 10184
0 10186 7 1 2 10183 10185
0 10187 5 1 1 10186
0 10188 7 1 2 28272 10187
0 10189 5 1 1 10188
0 10190 7 1 2 10175 10189
0 10191 5 1 1 10190
0 10192 7 1 2 35108 10191
0 10193 5 1 1 10192
0 10194 7 1 2 29227 34612
0 10195 5 1 1 10194
0 10196 7 1 2 32848 27395
0 10197 5 1 1 10196
0 10198 7 1 2 10195 10197
0 10199 5 1 1 10198
0 10200 7 2 2 24272 28703
0 10201 7 4 2 24767 25549
0 10202 7 1 2 35794 30848
0 10203 7 1 2 35792 10202
0 10204 7 1 2 10199 10203
0 10205 5 1 1 10204
0 10206 7 1 2 10193 10205
0 10207 5 1 1 10206
0 10208 7 1 2 22454 10207
0 10209 5 1 1 10208
0 10210 7 1 2 22827 32163
0 10211 7 2 2 35534 10210
0 10212 7 1 2 33282 35798
0 10213 5 1 1 10212
0 10214 7 3 2 23042 23262
0 10215 7 1 2 35800 30598
0 10216 7 1 2 34154 32327
0 10217 7 1 2 10215 10216
0 10218 5 1 1 10217
0 10219 7 1 2 24021 35109
0 10220 5 1 1 10219
0 10221 7 2 2 24884 25991
0 10222 7 2 2 35803 35795
0 10223 7 1 2 24273 35805
0 10224 5 1 1 10223
0 10225 7 1 2 10220 10224
0 10226 5 2 1 10225
0 10227 7 4 2 25792 27968
0 10228 5 1 1 35809
0 10229 7 1 2 23116 35810
0 10230 7 1 2 35807 10229
0 10231 5 1 1 10230
0 10232 7 1 2 10218 10231
0 10233 5 1 1 10232
0 10234 7 1 2 31944 10233
0 10235 5 1 1 10234
0 10236 7 1 2 10213 10235
0 10237 5 1 1 10236
0 10238 7 1 2 32245 10237
0 10239 5 1 1 10238
0 10240 7 4 2 22828 25304
0 10241 7 2 2 35675 32164
0 10242 7 1 2 35813 35817
0 10243 5 1 1 10242
0 10244 7 2 2 24022 24274
0 10245 7 1 2 35796 35819
0 10246 7 1 2 30381 10245
0 10247 5 1 1 10246
0 10248 7 1 2 10243 10247
0 10249 5 1 1 10248
0 10250 7 1 2 22616 10249
0 10251 5 1 1 10250
0 10252 7 1 2 35818 28837
0 10253 5 1 1 10252
0 10254 7 1 2 10251 10253
0 10255 5 1 1 10254
0 10256 7 1 2 32101 10255
0 10257 5 1 1 10256
0 10258 7 1 2 31866 35808
0 10259 5 1 1 10258
0 10260 7 1 2 10257 10259
0 10261 5 1 1 10260
0 10262 7 1 2 35652 10261
0 10263 5 1 1 10262
0 10264 7 1 2 34165 35799
0 10265 5 1 1 10264
0 10266 7 1 2 10263 10265
0 10267 5 1 1 10266
0 10268 7 1 2 34594 10267
0 10269 5 1 1 10268
0 10270 7 1 2 10239 10269
0 10271 7 1 2 10209 10270
0 10272 5 1 1 10271
0 10273 7 1 2 34937 10272
0 10274 5 1 1 10273
0 10275 7 1 2 28258 35099
0 10276 5 1 1 10275
0 10277 7 2 2 33425 35082
0 10278 5 1 1 35821
0 10279 7 1 2 35102 10278
0 10280 5 1 1 10279
0 10281 7 3 2 25793 10280
0 10282 7 1 2 27719 35823
0 10283 5 1 1 10282
0 10284 7 1 2 10276 10283
0 10285 5 1 1 10284
0 10286 7 1 2 32896 10285
0 10287 5 1 1 10286
0 10288 7 2 2 27785 32908
0 10289 7 1 2 35826 35824
0 10290 5 1 1 10289
0 10291 7 1 2 10287 10290
0 10292 5 1 1 10291
0 10293 7 1 2 25899 10292
0 10294 5 1 1 10293
0 10295 7 2 2 23802 29941
0 10296 7 1 2 22731 31422
0 10297 7 1 2 35828 10296
0 10298 7 1 2 32167 10297
0 10299 5 1 1 10298
0 10300 7 1 2 10294 10299
0 10301 5 1 1 10300
0 10302 7 1 2 22455 10301
0 10303 5 1 1 10302
0 10304 7 3 2 23117 35825
0 10305 7 3 2 25900 27909
0 10306 7 1 2 32897 35833
0 10307 7 1 2 35830 10306
0 10308 5 1 1 10307
0 10309 7 1 2 10303 10308
0 10310 5 1 1 10309
0 10311 7 1 2 34980 10310
0 10312 5 1 1 10311
0 10313 7 1 2 27969 35831
0 10314 5 1 1 10313
0 10315 7 2 2 22456 31277
0 10316 7 1 2 32165 33394
0 10317 7 2 2 35836 10316
0 10318 5 1 1 35838
0 10319 7 1 2 10314 10318
0 10320 5 1 1 10319
0 10321 7 3 2 30337 31869
0 10322 7 1 2 10320 35840
0 10323 5 1 1 10322
0 10324 7 3 2 22457 23043
0 10325 7 2 2 29895 35843
0 10326 7 1 2 31278 30599
0 10327 7 1 2 27688 10326
0 10328 7 1 2 35846 10327
0 10329 5 1 1 10328
0 10330 7 1 2 10323 10329
0 10331 5 1 1 10330
0 10332 7 1 2 28143 10331
0 10333 5 1 1 10332
0 10334 7 1 2 28235 35839
0 10335 5 1 1 10334
0 10336 7 1 2 29165 35832
0 10337 5 1 1 10336
0 10338 7 1 2 10335 10337
0 10339 5 1 1 10338
0 10340 7 1 2 10339 33801
0 10341 5 1 1 10340
0 10342 7 2 2 26970 34950
0 10343 7 1 2 23118 26746
0 10344 7 1 2 32437 10343
0 10345 7 1 2 35848 10344
0 10346 7 1 2 29308 10345
0 10347 5 1 1 10346
0 10348 7 1 2 10341 10347
0 10349 7 1 2 10333 10348
0 10350 5 1 1 10349
0 10351 7 1 2 32102 10350
0 10352 5 1 1 10351
0 10353 7 1 2 33860 35177
0 10354 5 1 1 10353
0 10355 7 5 2 23119 25436
0 10356 7 1 2 24885 35850
0 10357 7 1 2 35446 10356
0 10358 5 1 1 10357
0 10359 7 1 2 10354 10358
0 10360 5 1 1 10359
0 10361 7 1 2 27209 32511
0 10362 7 1 2 10360 10361
0 10363 7 1 2 32859 10362
0 10364 5 1 1 10363
0 10365 7 1 2 10352 10364
0 10366 7 1 2 10312 10365
0 10367 7 1 2 10274 10366
0 10368 5 1 1 10367
0 10369 7 1 2 28651 10368
0 10370 5 1 1 10369
0 10371 7 1 2 22950 31479
0 10372 5 1 1 10371
0 10373 7 1 2 26083 29649
0 10374 5 1 1 10373
0 10375 7 1 2 10372 10374
0 10376 5 3 1 10375
0 10377 7 1 2 28824 32603
0 10378 5 1 1 10377
0 10379 7 1 2 28731 32815
0 10380 5 1 1 10379
0 10381 7 1 2 27170 30871
0 10382 7 1 2 31433 10381
0 10383 5 1 1 10382
0 10384 7 4 2 22829 23414
0 10385 5 1 1 35858
0 10386 7 2 2 28032 35859
0 10387 7 1 2 32666 35862
0 10388 5 1 1 10387
0 10389 7 1 2 10383 10388
0 10390 7 1 2 10380 10389
0 10391 7 1 2 10378 10390
0 10392 5 1 1 10391
0 10393 7 1 2 23263 10392
0 10394 5 1 1 10393
0 10395 7 1 2 27210 31829
0 10396 7 1 2 32838 10395
0 10397 5 1 1 10396
0 10398 7 1 2 10394 10397
0 10399 5 1 1 10398
0 10400 7 1 2 22458 10399
0 10401 5 1 1 10400
0 10402 7 2 2 28033 35044
0 10403 7 1 2 25794 32840
0 10404 7 1 2 35864 10403
0 10405 5 1 1 10404
0 10406 7 1 2 10401 10405
0 10407 5 1 1 10406
0 10408 7 1 2 35855 10407
0 10409 5 1 1 10408
0 10410 7 1 2 22951 33602
0 10411 5 1 1 10410
0 10412 7 1 2 32189 31209
0 10413 5 1 1 10412
0 10414 7 1 2 10411 10413
0 10415 5 2 1 10414
0 10416 7 1 2 28086 35866
0 10417 5 1 1 10416
0 10418 7 1 2 22952 30825
0 10419 5 1 1 10418
0 10420 7 1 2 29650 33005
0 10421 5 1 1 10420
0 10422 7 1 2 10419 10421
0 10423 5 2 1 10422
0 10424 7 1 2 23347 35868
0 10425 5 1 1 10424
0 10426 7 1 2 25305 29930
0 10427 7 1 2 30360 10426
0 10428 5 1 1 10427
0 10429 7 1 2 10425 10428
0 10430 5 1 1 10429
0 10431 7 1 2 23803 10430
0 10432 5 1 1 10431
0 10433 7 1 2 35529 27110
0 10434 5 1 1 10433
0 10435 7 1 2 10432 10434
0 10436 5 1 1 10435
0 10437 7 1 2 22617 10436
0 10438 5 1 1 10437
0 10439 7 1 2 10417 10438
0 10440 5 1 1 10439
0 10441 7 1 2 32103 10440
0 10442 5 1 1 10441
0 10443 7 2 2 27314 30978
0 10444 5 1 1 35870
0 10445 7 2 2 32229 27410
0 10446 5 1 1 35872
0 10447 7 1 2 10444 10446
0 10448 5 2 1 10447
0 10449 7 1 2 22618 35874
0 10450 5 1 1 10449
0 10451 7 1 2 25901 31867
0 10452 5 1 1 10451
0 10453 7 1 2 10450 10452
0 10454 5 2 1 10453
0 10455 7 3 2 24104 35804
0 10456 7 1 2 23804 26783
0 10457 7 1 2 35878 10456
0 10458 7 1 2 35876 10457
0 10459 5 1 1 10458
0 10460 7 1 2 10442 10459
0 10461 5 1 1 10460
0 10462 7 1 2 28209 10461
0 10463 5 1 1 10462
0 10464 7 2 2 27257 34136
0 10465 5 2 1 35881
0 10466 7 2 2 27850 34347
0 10467 7 1 2 27315 35885
0 10468 5 1 1 10467
0 10469 7 1 2 28087 34345
0 10470 5 1 1 10469
0 10471 7 1 2 10468 10470
0 10472 7 1 2 35883 10471
0 10473 5 1 1 10472
0 10474 7 1 2 28210 10473
0 10475 5 1 1 10474
0 10476 7 1 2 30979 34402
0 10477 7 1 2 33092 10476
0 10478 5 1 1 10477
0 10479 7 1 2 10475 10478
0 10480 5 1 1 10479
0 10481 7 1 2 35526 10480
0 10482 5 1 1 10481
0 10483 7 1 2 10463 10482
0 10484 5 1 1 10483
0 10485 7 1 2 28990 10484
0 10486 5 1 1 10485
0 10487 7 1 2 10409 10486
0 10488 5 1 1 10487
0 10489 7 1 2 34885 10488
0 10490 5 1 1 10489
0 10491 7 1 2 31825 35294
0 10492 5 1 1 10491
0 10493 7 1 2 25550 31816
0 10494 7 1 2 27729 10493
0 10495 5 1 1 10494
0 10496 7 1 2 10492 10495
0 10497 5 2 1 10496
0 10498 7 1 2 35887 28045
0 10499 5 1 1 10498
0 10500 7 2 2 25795 35487
0 10501 7 1 2 35366 31532
0 10502 7 1 2 35889 10501
0 10503 5 1 1 10502
0 10504 7 1 2 10499 10503
0 10505 5 1 1 10504
0 10506 7 1 2 25902 10505
0 10507 5 1 1 10506
0 10508 7 3 2 22830 27851
0 10509 7 2 2 28034 35891
0 10510 7 1 2 35295 32409
0 10511 7 1 2 35894 10510
0 10512 5 1 1 10511
0 10513 7 1 2 10507 10512
0 10514 5 1 1 10513
0 10515 7 1 2 22459 10514
0 10516 5 1 1 10515
0 10517 7 7 2 23120 25796
0 10518 7 3 2 35488 35896
0 10519 7 2 2 35834 35903
0 10520 7 1 2 35906 28046
0 10521 5 1 1 10520
0 10522 7 1 2 10516 10521
0 10523 5 1 1 10522
0 10524 7 1 2 27083 10523
0 10525 5 1 1 10524
0 10526 7 2 2 35296 33224
0 10527 5 1 1 35908
0 10528 7 1 2 28236 35909
0 10529 5 1 1 10528
0 10530 7 1 2 35904 29166
0 10531 5 1 1 10530
0 10532 7 1 2 10529 10531
0 10533 5 2 1 10532
0 10534 7 1 2 35910 26998
0 10535 5 1 1 10534
0 10536 7 1 2 27970 35905
0 10537 5 1 1 10536
0 10538 7 1 2 10527 10537
0 10539 5 2 1 10538
0 10540 7 1 2 35912 32007
0 10541 5 1 1 10540
0 10542 7 1 2 31203 31046
0 10543 7 1 2 33646 10542
0 10544 7 1 2 35535 10543
0 10545 5 1 1 10544
0 10546 7 1 2 10541 10545
0 10547 5 1 1 10546
0 10548 7 1 2 28144 10547
0 10549 5 1 1 10548
0 10550 7 1 2 10535 10549
0 10551 5 1 1 10550
0 10552 7 1 2 27134 10551
0 10553 5 1 1 10552
0 10554 7 1 2 27564 35447
0 10555 5 1 1 10554
0 10556 7 1 2 35297 31915
0 10557 5 1 1 10556
0 10558 7 1 2 10555 10557
0 10559 5 1 1 10558
0 10560 7 1 2 10559 34749
0 10561 5 1 1 10560
0 10562 7 1 2 10553 10561
0 10563 7 1 2 10525 10562
0 10564 5 1 1 10563
0 10565 7 1 2 31480 10564
0 10566 5 1 1 10565
0 10567 7 1 2 32898 35888
0 10568 5 1 1 10567
0 10569 7 1 2 35827 35890
0 10570 5 1 1 10569
0 10571 7 1 2 10568 10570
0 10572 5 1 1 10571
0 10573 7 1 2 25903 10572
0 10574 5 1 1 10573
0 10575 7 1 2 24886 35801
0 10576 7 1 2 35829 10575
0 10577 7 1 2 34166 10576
0 10578 5 1 1 10577
0 10579 7 1 2 10574 10578
0 10580 5 1 1 10579
0 10581 7 1 2 22460 10580
0 10582 5 1 1 10581
0 10583 7 1 2 32899 35907
0 10584 5 1 1 10583
0 10585 7 1 2 10582 10584
0 10586 5 1 1 10585
0 10587 7 1 2 34786 10586
0 10588 5 1 1 10587
0 10589 7 1 2 30826 35911
0 10590 5 1 1 10589
0 10591 7 1 2 33536 35913
0 10592 5 1 1 10591
0 10593 7 1 2 30478 26396
0 10594 7 2 2 23264 29920
0 10595 7 1 2 35914 34474
0 10596 7 1 2 10593 10595
0 10597 5 1 1 10596
0 10598 7 1 2 10592 10597
0 10599 5 1 1 10598
0 10600 7 1 2 28145 10599
0 10601 5 1 1 10600
0 10602 7 1 2 10590 10601
0 10603 5 1 1 10602
0 10604 7 1 2 32104 10603
0 10605 5 1 1 10604
0 10606 7 1 2 29735 33013
0 10607 5 1 1 10606
0 10608 7 5 2 25992 30708
0 10609 7 1 2 25494 35456
0 10610 7 1 2 35916 10609
0 10611 5 1 1 10610
0 10612 7 1 2 10607 10611
0 10613 5 1 1 10612
0 10614 7 1 2 27211 30098
0 10615 7 1 2 10613 10614
0 10616 7 1 2 32860 10615
0 10617 5 1 1 10616
0 10618 7 1 2 10605 10617
0 10619 7 1 2 10588 10618
0 10620 5 1 1 10619
0 10621 7 1 2 28991 10620
0 10622 5 1 1 10621
0 10623 7 1 2 29167 31407
0 10624 5 1 1 10623
0 10625 7 1 2 27339 34204
0 10626 7 1 2 33201 10625
0 10627 7 1 2 28146 10626
0 10628 5 1 1 10627
0 10629 7 1 2 10624 10628
0 10630 5 1 1 10629
0 10631 7 2 2 35897 31902
0 10632 7 2 2 27506 35676
0 10633 7 1 2 35923 26540
0 10634 7 1 2 35921 10633
0 10635 7 1 2 10630 10634
0 10636 5 1 1 10635
0 10637 7 1 2 10622 10636
0 10638 7 1 2 10566 10637
0 10639 7 1 2 10490 10638
0 10640 7 1 2 10370 10639
0 10641 5 1 1 10640
0 10642 7 1 2 26320 10641
0 10643 5 1 1 10642
0 10644 7 1 2 32861 35506
0 10645 5 1 1 10644
0 10646 7 1 2 26342 34535
0 10647 7 1 2 29168 10646
0 10648 5 1 1 10647
0 10649 7 1 2 10645 10648
0 10650 5 1 1 10649
0 10651 7 1 2 30218 30193
0 10652 7 1 2 35922 10651
0 10653 7 1 2 10650 10652
0 10654 5 1 1 10653
0 10655 7 1 2 10643 10654
0 10656 5 1 1 10655
0 10657 7 1 2 23634 10656
0 10658 5 1 1 10657
0 10659 7 1 2 23415 34981
0 10660 5 1 1 10659
0 10661 7 1 2 23472 30930
0 10662 5 1 1 10661
0 10663 7 1 2 10660 10662
0 10664 5 1 1 10663
0 10665 7 1 2 22732 10664
0 10666 5 1 1 10665
0 10667 7 1 2 30835 33814
0 10668 5 1 1 10667
0 10669 7 1 2 10666 10668
0 10670 5 2 1 10669
0 10671 7 1 2 30225 35925
0 10672 5 1 1 10671
0 10673 7 2 2 32105 33802
0 10674 5 1 1 35927
0 10675 7 1 2 24687 35072
0 10676 5 1 1 10675
0 10677 7 1 2 10674 10676
0 10678 5 1 1 10677
0 10679 7 1 2 28237 10678
0 10680 5 1 1 10679
0 10681 7 1 2 10672 10680
0 10682 5 1 1 10681
0 10683 7 1 2 22831 10682
0 10684 5 1 1 10683
0 10685 7 1 2 28238 35584
0 10686 5 1 1 10685
0 10687 7 1 2 10684 10686
0 10688 5 1 1 10687
0 10689 7 1 2 27586 10688
0 10690 5 1 1 10689
0 10691 7 1 2 26755 32366
0 10692 7 1 2 34167 10691
0 10693 7 1 2 34161 10692
0 10694 5 1 1 10693
0 10695 7 1 2 10690 10694
0 10696 5 1 1 10695
0 10697 7 1 2 25551 10696
0 10698 5 1 1 10697
0 10699 7 1 2 31498 32398
0 10700 7 2 2 24968 30725
0 10701 7 2 2 26378 27744
0 10702 7 1 2 35929 35931
0 10703 7 1 2 10699 10702
0 10704 5 1 1 10703
0 10705 7 1 2 10698 10704
0 10706 5 1 1 10705
0 10707 7 1 2 24887 10706
0 10708 5 1 1 10707
0 10709 7 1 2 26247 30789
0 10710 7 1 2 28884 10709
0 10711 7 2 2 22953 28549
0 10712 7 2 2 31423 29874
0 10713 7 1 2 35933 35935
0 10714 7 1 2 10710 10713
0 10715 5 1 1 10714
0 10716 7 1 2 10708 10715
0 10717 5 1 1 10716
0 10718 7 1 2 35811 10717
0 10719 5 1 1 10718
0 10720 7 1 2 34298 33919
0 10721 5 1 1 10720
0 10722 7 1 2 31408 32381
0 10723 5 1 1 10722
0 10724 7 1 2 10721 10723
0 10725 5 1 1 10724
0 10726 7 1 2 25306 10725
0 10727 5 1 1 10726
0 10728 7 1 2 26084 35410
0 10729 5 1 1 10728
0 10730 7 1 2 10727 10729
0 10731 5 1 1 10730
0 10732 7 1 2 25993 10731
0 10733 5 1 1 10732
0 10734 7 1 2 28760 33375
0 10735 7 1 2 33796 10734
0 10736 5 1 1 10735
0 10737 7 1 2 10733 10736
0 10738 5 1 1 10737
0 10739 7 1 2 24592 10738
0 10740 5 1 1 10739
0 10741 7 1 2 31087 32868
0 10742 7 1 2 31726 10741
0 10743 5 1 1 10742
0 10744 7 1 2 10740 10743
0 10745 5 1 1 10744
0 10746 7 1 2 27777 34914
0 10747 7 1 2 10745 10746
0 10748 5 1 1 10747
0 10749 7 2 2 23121 35165
0 10750 7 1 2 32816 35937
0 10751 5 1 1 10750
0 10752 7 2 2 25552 27106
0 10753 7 2 2 35939 31959
0 10754 7 1 2 31194 35083
0 10755 7 1 2 35941 10754
0 10756 5 1 1 10755
0 10757 7 1 2 10751 10756
0 10758 5 1 1 10757
0 10759 7 1 2 34919 10758
0 10760 5 1 1 10759
0 10761 7 1 2 32604 35319
0 10762 5 1 1 10761
0 10763 7 1 2 27764 34579
0 10764 7 1 2 32663 10763
0 10765 5 1 1 10764
0 10766 7 2 2 29896 27689
0 10767 5 1 1 35943
0 10768 7 1 2 27852 28675
0 10769 7 1 2 35944 10768
0 10770 5 1 1 10769
0 10771 7 1 2 10765 10770
0 10772 7 1 2 10762 10771
0 10773 5 1 1 10772
0 10774 7 1 2 35938 10773
0 10775 5 1 1 10774
0 10776 7 1 2 10760 10775
0 10777 7 1 2 10748 10776
0 10778 5 1 1 10777
0 10779 7 1 2 28211 10778
0 10780 5 1 1 10779
0 10781 7 1 2 29169 34024
0 10782 5 1 1 10781
0 10783 7 2 2 30320 30993
0 10784 5 1 1 35945
0 10785 7 1 2 10782 10784
0 10786 5 1 1 10785
0 10787 7 1 2 27778 10786
0 10788 5 1 1 10787
0 10789 7 1 2 22619 35764
0 10790 5 1 1 10789
0 10791 7 2 2 27387 34430
0 10792 5 1 1 35947
0 10793 7 1 2 10790 10792
0 10794 5 2 1 10793
0 10795 7 2 2 22461 23122
0 10796 7 2 2 26756 35951
0 10797 7 1 2 28259 35953
0 10798 7 1 2 35949 10797
0 10799 5 1 1 10798
0 10800 7 1 2 10788 10799
0 10801 5 1 1 10800
0 10802 7 1 2 25904 10801
0 10803 5 1 1 10802
0 10804 7 1 2 27171 32147
0 10805 5 1 1 10804
0 10806 7 1 2 23805 27036
0 10807 7 1 2 32675 10806
0 10808 5 1 1 10807
0 10809 7 1 2 10805 10808
0 10810 5 1 1 10809
0 10811 7 1 2 35954 30781
0 10812 7 1 2 10810 10811
0 10813 5 1 1 10812
0 10814 7 1 2 10803 10813
0 10815 5 1 1 10814
0 10816 7 1 2 25553 10815
0 10817 5 1 1 10816
0 10818 7 1 2 24275 30014
0 10819 7 1 2 32505 10818
0 10820 5 1 1 10819
0 10821 7 1 2 10817 10820
0 10822 5 1 1 10821
0 10823 7 1 2 35053 10822
0 10824 5 1 1 10823
0 10825 7 1 2 28550 35182
0 10826 7 1 2 32435 10825
0 10827 5 1 1 10826
0 10828 7 1 2 10824 10827
0 10829 5 1 1 10828
0 10830 7 1 2 34938 10829
0 10831 5 1 1 10830
0 10832 7 1 2 10780 10831
0 10833 7 1 2 10719 10832
0 10834 5 1 1 10833
0 10835 7 1 2 28652 10834
0 10836 5 1 1 10835
0 10837 7 2 2 24023 26757
0 10838 7 2 2 31962 35955
0 10839 5 1 1 35957
0 10840 7 1 2 26776 27587
0 10841 5 1 1 10840
0 10842 7 1 2 10839 10841
0 10843 5 1 1 10842
0 10844 7 1 2 27287 10843
0 10845 5 1 1 10844
0 10846 7 1 2 26927 35558
0 10847 5 1 1 10846
0 10848 7 1 2 10845 10847
0 10849 5 1 1 10848
0 10850 7 1 2 25554 10849
0 10851 5 1 1 10850
0 10852 7 3 2 35820 32842
0 10853 7 1 2 35930 35959
0 10854 5 1 1 10853
0 10855 7 1 2 10851 10854
0 10856 5 1 1 10855
0 10857 7 1 2 22733 10856
0 10858 5 1 1 10857
0 10859 7 1 2 24688 35539
0 10860 7 1 2 27378 10859
0 10861 5 1 1 10860
0 10862 7 1 2 10858 10861
0 10863 5 1 1 10862
0 10864 7 1 2 32761 10863
0 10865 5 1 1 10864
0 10866 7 1 2 35544 33135
0 10867 7 1 2 35765 10866
0 10868 5 1 1 10867
0 10869 7 1 2 10865 10868
0 10870 5 1 1 10869
0 10871 7 1 2 22620 10870
0 10872 5 1 1 10871
0 10873 7 1 2 26916 32762
0 10874 5 1 1 10873
0 10875 7 1 2 5468 10874
0 10876 5 2 1 10875
0 10877 7 1 2 22734 35962
0 10878 5 1 1 10877
0 10879 7 1 2 10878 8064
0 10880 5 2 1 10879
0 10881 7 1 2 28088 35545
0 10882 7 1 2 35964 10881
0 10883 5 1 1 10882
0 10884 7 1 2 10872 10883
0 10885 5 1 1 10884
0 10886 7 1 2 22954 10885
0 10887 5 1 1 10886
0 10888 7 1 2 24888 32367
0 10889 7 1 2 33014 10888
0 10890 7 4 2 23044 27388
0 10891 7 1 2 35892 35966
0 10892 7 1 2 10889 10891
0 10893 5 1 1 10892
0 10894 7 1 2 10887 10893
0 10895 5 1 1 10894
0 10896 7 1 2 25797 10895
0 10897 5 1 1 10896
0 10898 7 1 2 28219 10897
0 10899 5 1 1 10898
0 10900 7 3 2 23123 35146
0 10901 7 1 2 32817 35970
0 10902 5 1 1 10901
0 10903 7 1 2 24593 27659
0 10904 7 1 2 35942 10903
0 10905 5 1 1 10904
0 10906 7 1 2 10902 10905
0 10907 5 2 1 10906
0 10908 7 1 2 32835 35973
0 10909 5 1 1 10908
0 10910 7 2 2 27713 35940
0 10911 7 1 2 22735 32878
0 10912 5 1 1 10911
0 10913 7 2 2 27340 30309
0 10914 5 1 1 35977
0 10915 7 1 2 25994 35978
0 10916 5 1 1 10915
0 10917 7 1 2 10912 10916
0 10918 5 1 1 10917
0 10919 7 1 2 25376 10918
0 10920 5 1 1 10919
0 10921 7 2 2 26085 33357
0 10922 5 1 1 35979
0 10923 7 1 2 26981 35980
0 10924 5 1 1 10923
0 10925 7 1 2 10920 10924
0 10926 5 1 1 10925
0 10927 7 1 2 35975 10926
0 10928 5 1 1 10927
0 10929 7 1 2 35971 4698
0 10930 5 1 1 10929
0 10931 7 1 2 28212 10930
0 10932 7 1 2 10928 10931
0 10933 7 1 2 10909 10932
0 10934 5 1 1 10933
0 10935 7 1 2 28956 35218
0 10936 7 1 2 10934 10935
0 10937 7 1 2 10899 10936
0 10938 5 1 1 10937
0 10939 7 1 2 27507 32711
0 10940 5 1 1 10939
0 10941 7 1 2 22955 34905
0 10942 5 1 1 10941
0 10943 7 1 2 10940 10942
0 10944 5 1 1 10943
0 10945 7 1 2 24768 10944
0 10946 5 1 1 10945
0 10947 7 1 2 27508 35504
0 10948 5 1 1 10947
0 10949 7 1 2 10946 10948
0 10950 5 1 1 10949
0 10951 7 1 2 35540 10950
0 10952 5 1 1 10951
0 10953 7 2 2 26758 35435
0 10954 7 1 2 27673 35981
0 10955 5 1 1 10954
0 10956 7 1 2 28588 33462
0 10957 5 1 1 10956
0 10958 7 1 2 10955 10957
0 10959 5 1 1 10958
0 10960 7 1 2 28992 29111
0 10961 7 1 2 10959 10960
0 10962 5 1 1 10961
0 10963 7 1 2 10952 10962
0 10964 5 1 1 10963
0 10965 7 1 2 32864 10964
0 10966 5 1 1 10965
0 10967 7 1 2 22736 35958
0 10968 5 1 1 10967
0 10969 7 1 2 32106 27596
0 10970 5 1 1 10969
0 10971 7 1 2 10968 10970
0 10972 5 1 1 10971
0 10973 7 1 2 23932 10972
0 10974 5 1 1 10973
0 10975 7 2 2 27411 27051
0 10976 5 1 1 35983
0 10977 7 1 2 27588 35984
0 10978 5 1 1 10977
0 10979 7 1 2 10974 10978
0 10980 5 1 1 10979
0 10981 7 1 2 25555 10980
0 10982 5 1 1 10981
0 10983 7 1 2 22737 28589
0 10984 7 1 2 35960 10983
0 10985 5 1 1 10984
0 10986 7 1 2 10982 10985
0 10987 5 1 1 10986
0 10988 7 1 2 26161 32630
0 10989 7 1 2 10987 10988
0 10990 5 1 1 10989
0 10991 7 1 2 27610 33790
0 10992 7 1 2 35541 10991
0 10993 7 1 2 34025 10992
0 10994 5 1 1 10993
0 10995 7 1 2 28239 10994
0 10996 7 1 2 10990 10995
0 10997 5 1 1 10996
0 10998 7 2 2 34854 33167
0 10999 5 1 1 35985
0 11000 7 2 2 30194 32609
0 11001 5 1 1 35987
0 11002 7 2 2 33180 32170
0 11003 5 1 1 35989
0 11004 7 1 2 11001 11003
0 11005 5 1 1 11004
0 11006 7 1 2 23416 11005
0 11007 5 1 1 11006
0 11008 7 2 2 28714 28509
0 11009 5 1 1 35991
0 11010 7 1 2 25995 35992
0 11011 5 1 1 11010
0 11012 7 1 2 11007 11011
0 11013 5 1 1 11012
0 11014 7 1 2 22738 11013
0 11015 5 1 1 11014
0 11016 7 1 2 10999 11015
0 11017 5 1 1 11016
0 11018 7 1 2 35546 11017
0 11019 5 1 1 11018
0 11020 7 1 2 28251 11019
0 11021 5 1 1 11020
0 11022 7 1 2 22956 28321
0 11023 7 1 2 11021 11022
0 11024 7 1 2 10997 11023
0 11025 5 1 1 11024
0 11026 7 3 2 24024 32631
0 11027 7 1 2 30726 30952
0 11028 7 1 2 35993 11027
0 11029 7 2 2 22739 29314
0 11030 7 2 2 26248 31634
0 11031 5 1 1 35998
0 11032 7 1 2 35996 35999
0 11033 7 1 2 11028 11032
0 11034 5 1 1 11033
0 11035 7 1 2 11025 11034
0 11036 5 1 1 11035
0 11037 7 1 2 25798 11036
0 11038 5 1 1 11037
0 11039 7 1 2 28220 11038
0 11040 5 1 1 11039
0 11041 7 1 2 26840 27611
0 11042 5 1 1 11041
0 11043 7 1 2 11042 11009
0 11044 5 1 1 11043
0 11045 7 1 2 35974 11044
0 11046 5 1 1 11045
0 11047 7 1 2 28929 32610
0 11048 5 1 1 11047
0 11049 7 4 2 23933 33159
0 11050 7 1 2 32632 36000
0 11051 5 1 1 11050
0 11052 7 1 2 11048 11051
0 11053 5 1 1 11052
0 11054 7 1 2 22740 11053
0 11055 5 1 1 11054
0 11056 7 1 2 27412 35988
0 11057 5 1 1 11056
0 11058 7 1 2 11055 11057
0 11059 5 1 1 11058
0 11060 7 1 2 25377 11059
0 11061 5 1 1 11060
0 11062 7 1 2 23934 35986
0 11063 5 1 1 11062
0 11064 7 1 2 11061 11063
0 11065 5 1 1 11064
0 11066 7 1 2 35976 11065
0 11067 5 1 1 11066
0 11068 7 1 2 28796 27612
0 11069 5 1 1 11068
0 11070 7 2 2 25307 28806
0 11071 7 1 2 28510 36004
0 11072 5 1 1 11071
0 11073 7 1 2 11069 11072
0 11074 5 1 1 11073
0 11075 7 1 2 32605 11074
0 11076 5 1 1 11075
0 11077 7 1 2 29362 34855
0 11078 7 1 2 33228 11077
0 11079 5 1 1 11078
0 11080 7 1 2 27107 27853
0 11081 7 1 2 35256 11080
0 11082 7 1 2 33083 11081
0 11083 5 1 1 11082
0 11084 7 1 2 11079 11083
0 11085 7 1 2 11076 11084
0 11086 5 1 1 11085
0 11087 7 1 2 35972 11086
0 11088 5 1 1 11087
0 11089 7 1 2 28213 11088
0 11090 7 1 2 11067 11089
0 11091 7 1 2 11046 11090
0 11092 5 1 1 11091
0 11093 7 1 2 28957 32547
0 11094 7 1 2 11092 11093
0 11095 7 1 2 11040 11094
0 11096 5 1 1 11095
0 11097 7 1 2 10966 11096
0 11098 7 1 2 10938 11097
0 11099 7 1 2 10836 11098
0 11100 7 1 2 10658 11099
0 11101 5 1 1 11100
0 11102 7 2 2 35335 11101
0 11103 5 1 1 36006
0 11104 7 1 2 25122 11103
0 11105 5 1 1 11104
0 11106 7 1 2 22348 11105
0 11107 7 1 2 10138 11106
0 11108 5 1 1 11107
0 11109 7 4 2 22462 25123
0 11110 7 2 2 27816 33608
0 11111 7 1 2 36008 36012
0 11112 5 1 1 11111
0 11113 7 1 2 24455 33603
0 11114 5 1 1 11113
0 11115 7 8 2 25495 23806
0 11116 7 1 2 22463 36014
0 11117 7 1 2 33513 11116
0 11118 5 1 1 11117
0 11119 7 1 2 11114 11118
0 11120 5 1 1 11119
0 11121 7 1 2 23189 11120
0 11122 5 1 1 11121
0 11123 7 1 2 11112 11122
0 11124 5 1 1 11123
0 11125 7 1 2 25695 11124
0 11126 5 1 1 11125
0 11127 7 1 2 23190 29636
0 11128 7 1 2 33609 11127
0 11129 5 1 1 11128
0 11130 7 1 2 11126 11129
0 11131 5 1 1 11130
0 11132 7 2 2 26249 28993
0 11133 7 1 2 22957 36022
0 11134 7 1 2 11131 11133
0 11135 5 1 1 11134
0 11136 7 1 2 25437 30600
0 11137 5 1 1 11136
0 11138 7 1 2 26573 35221
0 11139 5 2 1 11138
0 11140 7 1 2 11137 36024
0 11141 5 1 1 11140
0 11142 7 2 2 24769 11141
0 11143 5 1 1 36026
0 11144 7 1 2 28966 32377
0 11145 5 2 1 11144
0 11146 7 1 2 11143 36028
0 11147 5 2 1 11146
0 11148 7 2 2 23807 31122
0 11149 7 1 2 23191 36032
0 11150 7 1 2 36030 11149
0 11151 5 1 1 11150
0 11152 7 7 2 26250 27817
0 11153 5 1 1 36034
0 11154 7 2 2 22958 26343
0 11155 7 2 2 36035 36041
0 11156 5 1 1 36043
0 11157 7 1 2 25124 31799
0 11158 7 1 2 36044 11157
0 11159 5 1 1 11158
0 11160 7 1 2 11151 11159
0 11161 5 1 1 11160
0 11162 7 1 2 22464 11161
0 11163 5 1 1 11162
0 11164 7 6 2 24276 32391
0 11165 5 1 1 36045
0 11166 7 1 2 25438 32190
0 11167 7 1 2 36046 11166
0 11168 5 1 1 11167
0 11169 7 2 2 25905 35677
0 11170 7 1 2 23808 35513
0 11171 7 1 2 36051 11170
0 11172 5 1 1 11171
0 11173 7 1 2 11168 11172
0 11174 5 1 1 11173
0 11175 7 1 2 22832 11174
0 11176 5 1 1 11175
0 11177 7 1 2 32191 36027
0 11178 5 1 1 11177
0 11179 7 1 2 11176 11178
0 11180 5 1 1 11179
0 11181 7 1 2 33983 11180
0 11182 5 1 1 11181
0 11183 7 1 2 11163 11182
0 11184 5 1 1 11183
0 11185 7 1 2 25696 11184
0 11186 5 1 1 11185
0 11187 7 1 2 23192 36042
0 11188 7 5 2 23704 33647
0 11189 7 1 2 36052 36053
0 11190 7 1 2 11187 11189
0 11191 5 1 1 11190
0 11192 7 1 2 11186 11191
0 11193 5 1 1 11192
0 11194 7 1 2 31481 11193
0 11195 5 1 1 11194
0 11196 7 1 2 26344 34669
0 11197 5 1 1 11196
0 11198 7 3 2 34787 26894
0 11199 7 1 2 31648 36058
0 11200 5 1 1 11199
0 11201 7 1 2 11197 11200
0 11202 5 1 1 11201
0 11203 7 1 2 23193 11202
0 11204 5 1 1 11203
0 11205 7 4 2 30338 28704
0 11206 7 2 2 26162 36061
0 11207 7 3 2 22833 32633
0 11208 7 1 2 33672 36067
0 11209 7 1 2 36065 11208
0 11210 5 1 1 11209
0 11211 7 1 2 11204 11210
0 11212 5 1 1 11211
0 11213 7 1 2 22465 11212
0 11214 5 1 1 11213
0 11215 7 1 2 33604 26345
0 11216 5 1 1 11215
0 11217 7 1 2 27212 36059
0 11218 5 1 1 11217
0 11219 7 1 2 11216 11218
0 11220 5 1 1 11219
0 11221 7 1 2 23194 31102
0 11222 7 1 2 11220 11221
0 11223 5 1 1 11222
0 11224 7 1 2 11214 11223
0 11225 5 1 1 11224
0 11226 7 1 2 36047 11225
0 11227 5 1 1 11226
0 11228 7 3 2 33923 33466
0 11229 7 1 2 33616 36070
0 11230 5 1 1 11229
0 11231 7 1 2 27236 34096
0 11232 5 1 1 11231
0 11233 7 1 2 10767 11232
0 11234 5 6 1 11233
0 11235 7 1 2 25697 36073
0 11236 5 2 1 11235
0 11237 7 1 2 24456 36079
0 11238 5 1 1 11237
0 11239 7 1 2 35841 31607
0 11240 5 1 1 11239
0 11241 7 1 2 35170 34803
0 11242 5 1 1 11241
0 11243 7 3 2 11240 11242
0 11244 5 2 1 36081
0 11245 7 1 2 22466 36082
0 11246 5 1 1 11245
0 11247 7 1 2 22834 11246
0 11248 7 1 2 11238 11247
0 11249 5 1 1 11248
0 11250 7 1 2 11230 11249
0 11251 5 1 1 11250
0 11252 7 4 2 24889 26251
0 11253 5 1 1 36086
0 11254 7 1 2 11253 31754
0 11255 5 1 1 11254
0 11256 7 1 2 23195 11255
0 11257 7 1 2 11251 11256
0 11258 5 1 1 11257
0 11259 7 1 2 24890 11153
0 11260 5 1 1 11259
0 11261 7 1 2 22467 26346
0 11262 7 1 2 33673 11261
0 11263 7 1 2 30055 36062
0 11264 7 1 2 11262 11263
0 11265 7 1 2 11260 11264
0 11266 5 1 1 11265
0 11267 7 1 2 11258 11266
0 11268 5 1 1 11267
0 11269 7 1 2 28653 11268
0 11270 5 1 1 11269
0 11271 7 1 2 11227 11270
0 11272 7 1 2 11195 11271
0 11273 7 1 2 11135 11272
0 11274 5 1 1 11273
0 11275 7 1 2 22349 11274
0 11276 5 1 1 11275
0 11277 7 1 2 23473 35856
0 11278 5 1 1 11277
0 11279 7 1 2 27654 30679
0 11280 5 1 1 11279
0 11281 7 1 2 11278 11280
0 11282 5 1 1 11281
0 11283 7 1 2 22835 11282
0 11284 5 1 1 11283
0 11285 7 1 2 7881 11284
0 11286 5 2 1 11285
0 11287 7 1 2 36036 36090
0 11288 5 1 1 11287
0 11289 7 1 2 26347 26574
0 11290 7 1 2 29988 11289
0 11291 5 1 1 11290
0 11292 7 1 2 11288 11291
0 11293 5 1 1 11292
0 11294 7 1 2 31800 34246
0 11295 7 1 2 11293 11294
0 11296 5 1 1 11295
0 11297 7 1 2 11276 11296
0 11298 5 1 1 11297
0 11299 7 1 2 25556 11298
0 11300 5 1 1 11299
0 11301 7 1 2 35844 33383
0 11302 7 1 2 35793 11301
0 11303 7 1 2 34637 11302
0 11304 7 1 2 36091 11303
0 11305 5 1 1 11304
0 11306 7 1 2 11300 11305
0 11307 5 1 1 11306
0 11308 7 1 2 28147 11307
0 11309 5 1 1 11308
0 11310 7 1 2 25072 26759
0 11311 5 1 1 11310
0 11312 7 4 2 33485 11311
0 11313 7 2 2 31455 36092
0 11314 5 1 1 36096
0 11315 7 1 2 32328 33477
0 11316 5 1 1 11315
0 11317 7 1 2 11314 11316
0 11318 5 2 1 11317
0 11319 7 1 2 29665 35586
0 11320 5 1 1 11319
0 11321 7 1 2 26971 32487
0 11322 5 1 1 11321
0 11323 7 1 2 33006 26895
0 11324 5 1 1 11323
0 11325 7 1 2 11322 11324
0 11326 5 3 1 11325
0 11327 7 1 2 30361 36100
0 11328 5 1 1 11327
0 11329 7 1 2 11320 11328
0 11330 5 2 1 11329
0 11331 7 1 2 36098 36103
0 11332 5 1 1 11331
0 11333 7 1 2 35587 29853
0 11334 5 1 1 11333
0 11335 7 2 2 24025 32488
0 11336 5 1 1 36105
0 11337 7 2 2 25996 35778
0 11338 5 1 1 36107
0 11339 7 1 2 11336 11338
0 11340 5 5 1 11339
0 11341 7 2 2 26456 30491
0 11342 7 2 2 36109 36114
0 11343 5 1 1 36116
0 11344 7 1 2 11334 11343
0 11345 5 1 1 11344
0 11346 7 1 2 33617 33582
0 11347 7 1 2 11345 11346
0 11348 5 1 1 11347
0 11349 7 1 2 11332 11348
0 11350 5 1 1 11349
0 11351 7 1 2 22350 34483
0 11352 7 1 2 34234 11351
0 11353 7 1 2 11350 11352
0 11354 5 1 1 11353
0 11355 7 1 2 11309 11354
0 11356 5 1 1 11355
0 11357 7 1 2 25225 11356
0 11358 5 1 1 11357
0 11359 7 1 2 36009 36074
0 11360 5 1 1 11359
0 11361 7 2 2 24457 25439
0 11362 7 1 2 29897 36118
0 11363 7 1 2 34289 11362
0 11364 5 1 1 11363
0 11365 7 1 2 11360 11364
0 11366 5 1 1 11365
0 11367 7 1 2 25698 11366
0 11368 5 1 1 11367
0 11369 7 1 2 35266 33984
0 11370 7 1 2 36063 11369
0 11371 5 1 1 11370
0 11372 7 1 2 11368 11371
0 11373 5 1 1 11372
0 11374 7 1 2 22836 11373
0 11375 5 1 1 11374
0 11376 7 5 2 25799 36010
0 11377 5 1 1 36120
0 11378 7 2 2 24458 33697
0 11379 5 2 1 36125
0 11380 7 1 2 11377 36127
0 11381 5 5 1 11380
0 11382 7 1 2 36071 36129
0 11383 5 1 1 11382
0 11384 7 1 2 11375 11383
0 11385 5 1 1 11384
0 11386 7 1 2 22351 11385
0 11387 5 1 1 11386
0 11388 7 1 2 22837 36075
0 11389 5 1 1 11388
0 11390 7 1 2 32192 33924
0 11391 5 1 1 11390
0 11392 7 1 2 11389 11391
0 11393 5 2 1 11392
0 11394 7 1 2 34247 36134
0 11395 5 1 1 11394
0 11396 7 1 2 11387 11395
0 11397 5 1 1 11396
0 11398 7 1 2 28148 11397
0 11399 5 1 1 11398
0 11400 7 2 2 23348 35588
0 11401 5 1 1 36136
0 11402 7 1 2 34638 31811
0 11403 7 1 2 36137 11402
0 11404 5 1 1 11403
0 11405 7 1 2 11399 11404
0 11406 5 1 1 11405
0 11407 7 1 2 29288 31064
0 11408 7 1 2 11406 11407
0 11409 5 1 1 11408
0 11410 7 2 2 27022 34097
0 11411 5 1 1 36138
0 11412 7 1 2 22838 36139
0 11413 5 1 1 11412
0 11414 7 1 2 11401 11413
0 11415 5 1 1 11414
0 11416 7 1 2 22621 11415
0 11417 5 1 1 11416
0 11418 7 1 2 23474 33343
0 11419 5 1 1 11418
0 11420 7 1 2 11417 11419
0 11421 5 2 1 11420
0 11422 7 1 2 24190 36037
0 11423 5 1 1 11422
0 11424 7 1 2 32271 11423
0 11425 5 1 1 11424
0 11426 7 1 2 31456 34639
0 11427 7 1 2 11425 11426
0 11428 7 1 2 36140 11427
0 11429 5 1 1 11428
0 11430 7 1 2 11409 11429
0 11431 5 1 1 11430
0 11432 7 1 2 25557 11431
0 11433 5 1 1 11432
0 11434 7 1 2 27493 30146
0 11435 7 2 2 34640 11434
0 11436 7 1 2 32299 36142
0 11437 7 1 2 36141 11436
0 11438 5 1 1 11437
0 11439 7 1 2 23547 11438
0 11440 7 1 2 11433 11439
0 11441 5 1 1 11440
0 11442 7 4 2 24026 33934
0 11443 7 1 2 27437 36097
0 11444 5 1 1 11443
0 11445 7 1 2 22468 33478
0 11446 7 1 2 27258 11445
0 11447 5 1 1 11446
0 11448 7 1 2 11444 11447
0 11449 5 1 1 11448
0 11450 7 1 2 22622 11449
0 11451 5 1 1 11450
0 11452 7 1 2 23349 33648
0 11453 7 1 2 33845 33479
0 11454 7 1 2 11452 11453
0 11455 5 1 1 11454
0 11456 7 1 2 11451 11455
0 11457 5 1 1 11456
0 11458 7 1 2 36144 11457
0 11459 5 1 1 11458
0 11460 7 1 2 36099 33829
0 11461 5 1 1 11460
0 11462 7 1 2 11459 11461
0 11463 5 1 1 11462
0 11464 7 1 2 34321 11463
0 11465 5 1 1 11464
0 11466 7 2 2 34290 33781
0 11467 7 2 2 36145 36148
0 11468 5 1 1 36150
0 11469 7 1 2 28149 33480
0 11470 7 1 2 36151 11469
0 11471 5 1 1 11470
0 11472 7 1 2 11465 11471
0 11473 5 1 1 11472
0 11474 7 1 2 26163 11473
0 11475 5 1 1 11474
0 11476 7 1 2 22352 36130
0 11477 5 1 1 11476
0 11478 7 4 2 23196 25800
0 11479 7 1 2 36152 34008
0 11480 5 1 1 11479
0 11481 7 1 2 11477 11480
0 11482 5 1 1 11481
0 11483 7 1 2 30508 11482
0 11484 5 1 1 11483
0 11485 7 4 2 25906 28240
0 11486 7 1 2 34322 33618
0 11487 7 1 2 36156 11486
0 11488 5 1 1 11487
0 11489 7 1 2 11484 11488
0 11490 5 1 1 11489
0 11491 7 2 2 29282 33557
0 11492 7 1 2 36110 36160
0 11493 7 1 2 11490 11492
0 11494 5 1 1 11493
0 11495 7 1 2 11475 11494
0 11496 5 1 1 11495
0 11497 7 1 2 25699 11496
0 11498 5 1 1 11497
0 11499 7 2 2 35254 36111
0 11500 7 4 2 22469 25073
0 11501 7 1 2 23935 36164
0 11502 7 1 2 36162 11501
0 11503 5 1 1 11502
0 11504 7 3 2 26348 31905
0 11505 7 2 2 26164 35562
0 11506 7 1 2 33010 36171
0 11507 7 1 2 36168 11506
0 11508 5 1 1 11507
0 11509 7 1 2 11503 11508
0 11510 5 1 1 11509
0 11511 7 1 2 28150 11510
0 11512 5 1 1 11511
0 11513 7 2 2 24277 34073
0 11514 5 1 1 36173
0 11515 7 1 2 36112 36174
0 11516 5 1 1 11515
0 11517 7 1 2 33558 36106
0 11518 5 1 1 11517
0 11519 7 1 2 11516 11518
0 11520 5 1 1 11519
0 11521 7 1 2 24459 28487
0 11522 7 1 2 36157 11521
0 11523 7 1 2 11520 11522
0 11524 5 1 1 11523
0 11525 7 1 2 11512 11524
0 11526 5 1 1 11525
0 11527 7 1 2 25801 11526
0 11528 5 1 1 11527
0 11529 7 1 2 32673 34229
0 11530 7 1 2 36163 11529
0 11531 5 1 1 11530
0 11532 7 1 2 11528 11531
0 11533 5 1 1 11532
0 11534 7 1 2 33945 11533
0 11535 5 1 1 11534
0 11536 7 1 2 25496 11535
0 11537 7 1 2 11498 11536
0 11538 5 1 1 11537
0 11539 7 1 2 11441 11538
0 11540 5 1 1 11539
0 11541 7 1 2 24891 11540
0 11542 5 1 1 11541
0 11543 7 1 2 22470 36135
0 11544 5 1 1 11543
0 11545 7 1 2 24460 28705
0 11546 7 1 2 33826 11545
0 11547 5 1 1 11546
0 11548 7 1 2 11544 11547
0 11549 5 1 1 11548
0 11550 7 1 2 34323 11549
0 11551 5 1 1 11550
0 11552 7 1 2 11468 11551
0 11553 5 1 1 11552
0 11554 7 1 2 25700 11553
0 11555 5 1 1 11554
0 11556 7 1 2 29931 33787
0 11557 7 1 2 34376 11556
0 11558 5 1 1 11557
0 11559 7 1 2 11555 11558
0 11560 5 1 1 11559
0 11561 7 1 2 32282 11560
0 11562 5 1 1 11561
0 11563 7 5 2 23809 29760
0 11564 7 1 2 26349 36175
0 11565 5 1 1 11564
0 11566 7 1 2 32193 26896
0 11567 5 1 1 11566
0 11568 7 1 2 11565 11567
0 11569 5 1 1 11568
0 11570 7 1 2 22471 11569
0 11571 5 1 1 11570
0 11572 7 1 2 27818 34149
0 11573 7 1 2 36169 11572
0 11574 5 1 1 11573
0 11575 7 1 2 11571 11574
0 11576 5 1 1 11575
0 11577 7 1 2 34324 11576
0 11578 5 1 1 11577
0 11579 7 1 2 33340 36119
0 11580 7 1 2 34546 11579
0 11581 5 1 1 11580
0 11582 7 1 2 11578 11581
0 11583 5 1 1 11582
0 11584 7 1 2 25701 11583
0 11585 5 1 1 11584
0 11586 7 2 2 23475 29761
0 11587 7 1 2 25802 33041
0 11588 7 1 2 33946 11587
0 11589 7 1 2 36180 11588
0 11590 5 1 1 11589
0 11591 7 1 2 11585 11590
0 11592 5 1 1 11591
0 11593 7 1 2 31482 11592
0 11594 5 1 1 11593
0 11595 7 1 2 34632 36149
0 11596 5 1 1 11595
0 11597 7 1 2 24461 36013
0 11598 5 1 1 11597
0 11599 7 1 2 33606 11598
0 11600 5 1 1 11599
0 11601 7 1 2 34325 11600
0 11602 5 1 1 11601
0 11603 7 1 2 11596 11602
0 11604 5 1 1 11603
0 11605 7 1 2 25702 11604
0 11606 5 1 1 11605
0 11607 7 1 2 34667 34722
0 11608 5 1 1 11607
0 11609 7 1 2 11606 11608
0 11610 5 1 1 11609
0 11611 7 1 2 28994 11610
0 11612 5 1 1 11611
0 11613 7 1 2 11594 11612
0 11614 5 1 1 11613
0 11615 7 1 2 26252 11614
0 11616 5 1 1 11615
0 11617 7 1 2 11562 11616
0 11618 5 1 1 11617
0 11619 7 1 2 25558 11618
0 11620 5 1 1 11619
0 11621 7 1 2 28005 30680
0 11622 5 1 1 11621
0 11623 7 3 2 32714 30469
0 11624 5 1 1 36182
0 11625 7 1 2 23476 31483
0 11626 5 1 1 11625
0 11627 7 1 2 11624 11626
0 11628 5 1 1 11627
0 11629 7 1 2 22839 11628
0 11630 5 1 1 11629
0 11631 7 1 2 11622 11630
0 11632 5 2 1 11631
0 11633 7 1 2 31801 36143
0 11634 7 1 2 36185 11633
0 11635 5 1 1 11634
0 11636 7 1 2 11620 11635
0 11637 5 1 1 11636
0 11638 7 1 2 28151 11637
0 11639 5 1 1 11638
0 11640 7 3 2 26804 35589
0 11641 7 1 2 26575 36187
0 11642 5 1 1 11641
0 11643 7 1 2 26972 26350
0 11644 5 1 1 11643
0 11645 7 1 2 202 11644
0 11646 5 2 1 11645
0 11647 7 1 2 31484 36190
0 11648 5 1 1 11647
0 11649 7 1 2 28995 30827
0 11650 5 1 1 11649
0 11651 7 1 2 11648 11650
0 11652 5 2 1 11651
0 11653 7 1 2 26253 7045
0 11654 7 1 2 36192 11653
0 11655 5 1 1 11654
0 11656 7 1 2 11642 11655
0 11657 5 1 1 11656
0 11658 7 1 2 25559 33619
0 11659 7 1 2 11657 11658
0 11660 5 1 1 11659
0 11661 7 2 2 24278 28551
0 11662 7 2 2 36194 36193
0 11663 7 1 2 31457 36196
0 11664 5 1 1 11663
0 11665 7 1 2 11660 11664
0 11666 5 1 1 11665
0 11667 7 1 2 28241 34641
0 11668 7 1 2 11666 11667
0 11669 5 1 1 11668
0 11670 7 1 2 22959 11669
0 11671 7 1 2 11639 11670
0 11672 5 1 1 11671
0 11673 7 1 2 23265 11672
0 11674 7 1 2 11542 11673
0 11675 5 1 1 11674
0 11676 7 1 2 11358 11675
0 11677 5 1 1 11676
0 11678 7 1 2 25626 11677
0 11679 5 1 1 11678
0 11680 7 1 2 30434 33958
0 11681 5 1 1 11680
0 11682 7 1 2 25125 31835
0 11683 5 1 1 11682
0 11684 7 1 2 11681 11683
0 11685 5 3 1 11684
0 11686 7 1 2 22623 36198
0 11687 5 1 1 11686
0 11688 7 1 2 30891 33959
0 11689 5 1 1 11688
0 11690 7 1 2 11687 11689
0 11691 5 1 1 11690
0 11692 7 1 2 11691 34493
0 11693 5 1 1 11692
0 11694 7 1 2 23197 28361
0 11695 7 1 2 33456 11694
0 11696 7 1 2 31643 11695
0 11697 5 1 1 11696
0 11698 7 1 2 11693 11697
0 11699 5 1 1 11698
0 11700 7 1 2 22353 11699
0 11701 5 1 1 11700
0 11702 7 1 2 28242 31966
0 11703 7 1 2 34700 11702
0 11704 5 1 1 11703
0 11705 7 1 2 11701 11704
0 11706 5 1 1 11705
0 11707 7 1 2 36146 11706
0 11708 5 1 1 11707
0 11709 7 1 2 24892 34558
0 11710 7 1 2 34533 11709
0 11711 5 1 1 11710
0 11712 7 3 2 24893 33674
0 11713 5 1 1 36201
0 11714 7 1 2 34862 34389
0 11715 5 1 1 11714
0 11716 7 1 2 11713 11715
0 11717 5 1 1 11716
0 11718 7 1 2 22354 11717
0 11719 5 1 1 11718
0 11720 7 1 2 7141 11719
0 11721 5 2 1 11720
0 11722 7 1 2 23266 33241
0 11723 7 1 2 36204 11722
0 11724 5 1 1 11723
0 11725 7 1 2 11711 11724
0 11726 5 1 1 11725
0 11727 7 1 2 33827 11726
0 11728 5 1 1 11727
0 11729 7 1 2 11708 11728
0 11730 5 1 1 11729
0 11731 7 1 2 23810 11730
0 11732 5 1 1 11731
0 11733 7 2 2 24894 33960
0 11734 7 2 2 22355 22840
0 11735 7 1 2 35267 36208
0 11736 7 1 2 30347 11735
0 11737 7 1 2 36206 11736
0 11738 5 1 1 11737
0 11739 7 1 2 30782 36147
0 11740 7 1 2 36205 11739
0 11741 5 1 1 11740
0 11742 7 1 2 11738 11741
0 11743 5 1 1 11742
0 11744 7 1 2 25803 28152
0 11745 7 1 2 11743 11744
0 11746 5 1 1 11745
0 11747 7 1 2 11732 11746
0 11748 5 1 1 11747
0 11749 7 1 2 22472 11748
0 11750 5 1 1 11749
0 11751 7 1 2 36072 28288
0 11752 5 1 1 11751
0 11753 7 1 2 25226 36080
0 11754 5 1 1 11753
0 11755 7 1 2 23267 36083
0 11756 5 1 1 11755
0 11757 7 1 2 22841 11756
0 11758 7 1 2 11754 11757
0 11759 5 1 1 11758
0 11760 7 1 2 11752 11759
0 11761 5 1 1 11760
0 11762 7 2 2 24895 28153
0 11763 7 1 2 11761 36210
0 11764 5 1 1 11763
0 11765 7 2 2 33278 34359
0 11766 7 1 2 34863 36212
0 11767 7 1 2 35590 11766
0 11768 5 1 1 11767
0 11769 7 1 2 11764 11768
0 11770 5 1 1 11769
0 11771 7 1 2 34723 11770
0 11772 5 1 1 11771
0 11773 7 1 2 11750 11772
0 11774 5 1 1 11773
0 11775 7 1 2 28654 11774
0 11776 5 1 1 11775
0 11777 7 6 2 24770 25497
0 11778 7 1 2 27213 28565
0 11779 7 1 2 36214 11778
0 11780 5 1 1 11779
0 11781 7 2 2 23548 23811
0 11782 7 3 2 25907 33160
0 11783 7 2 2 22842 36222
0 11784 7 1 2 36220 36225
0 11785 5 1 1 11784
0 11786 7 1 2 11780 11785
0 11787 5 1 1 11786
0 11788 7 1 2 34463 11787
0 11789 5 1 1 11788
0 11790 7 2 2 24191 27971
0 11791 7 1 2 32057 36215
0 11792 7 1 2 28454 11791
0 11793 7 1 2 36227 11792
0 11794 5 1 1 11793
0 11795 7 1 2 11789 11794
0 11796 5 1 1 11795
0 11797 7 1 2 25703 11796
0 11798 5 1 1 11797
0 11799 7 2 2 34150 30112
0 11800 7 1 2 36209 34697
0 11801 7 1 2 36229 11800
0 11802 7 1 2 29791 11801
0 11803 5 1 1 11802
0 11804 7 1 2 11798 11803
0 11805 5 1 1 11804
0 11806 7 1 2 22960 11805
0 11807 5 1 1 11806
0 11808 7 2 2 22356 23268
0 11809 7 8 2 22473 24771
0 11810 7 1 2 27214 36233
0 11811 7 1 2 36231 11810
0 11812 7 2 2 24896 34390
0 11813 7 2 2 30276 34864
0 11814 7 1 2 36241 36243
0 11815 7 1 2 11811 11814
0 11816 5 1 1 11815
0 11817 7 1 2 11807 11816
0 11818 5 1 1 11817
0 11819 7 1 2 28154 11818
0 11820 5 1 1 11819
0 11821 7 1 2 22357 33971
0 11822 5 1 1 11821
0 11823 7 5 2 23350 27896
0 11824 7 1 2 33637 36245
0 11825 5 1 1 11824
0 11826 7 1 2 11822 11825
0 11827 5 2 1 11826
0 11828 7 1 2 28511 33117
0 11829 5 1 1 11828
0 11830 7 1 2 26948 35047
0 11831 5 1 1 11830
0 11832 7 1 2 11829 11831
0 11833 5 1 1 11832
0 11834 7 1 2 30550 11833
0 11835 7 1 2 36250 11834
0 11836 5 1 1 11835
0 11837 7 1 2 27438 36232
0 11838 7 1 2 30455 11837
0 11839 7 1 2 30277 35797
0 11840 7 1 2 36242 11839
0 11841 7 1 2 11838 11840
0 11842 5 1 1 11841
0 11843 7 1 2 11836 11842
0 11844 5 1 1 11843
0 11845 7 1 2 32329 11844
0 11846 5 1 1 11845
0 11847 7 1 2 30382 26870
0 11848 7 1 2 36153 30534
0 11849 7 1 2 11847 11848
0 11850 7 1 2 36244 34520
0 11851 7 1 2 11849 11850
0 11852 5 1 1 11851
0 11853 7 1 2 11846 11852
0 11854 7 1 2 11820 11853
0 11855 5 1 1 11854
0 11856 7 1 2 32455 11855
0 11857 5 1 1 11856
0 11858 7 2 2 35079 30551
0 11859 7 1 2 36251 36252
0 11860 5 1 1 11859
0 11861 7 2 2 35084 29325
0 11862 7 2 2 34865 36254
0 11863 7 1 2 32058 36246
0 11864 7 1 2 36256 11863
0 11865 5 1 1 11864
0 11866 7 1 2 11860 11865
0 11867 5 1 1 11866
0 11868 7 1 2 32330 11867
0 11869 5 1 1 11868
0 11870 7 2 2 25560 25804
0 11871 7 1 2 28368 36258
0 11872 7 1 2 33947 36255
0 11873 7 1 2 11871 11872
0 11874 5 1 1 11873
0 11875 7 1 2 11869 11874
0 11876 5 1 1 11875
0 11877 7 1 2 33803 11876
0 11878 5 1 1 11877
0 11879 7 1 2 34464 36253
0 11880 5 1 1 11879
0 11881 7 1 2 36257 34441
0 11882 5 1 1 11881
0 11883 7 1 2 11880 11882
0 11884 5 1 1 11883
0 11885 7 1 2 36076 11884
0 11886 5 1 1 11885
0 11887 7 2 2 27972 36084
0 11888 7 1 2 22961 32059
0 11889 7 1 2 35080 11888
0 11890 7 1 2 36260 11889
0 11891 5 1 1 11890
0 11892 7 1 2 11886 11891
0 11893 5 1 1 11892
0 11894 7 1 2 28155 11893
0 11895 5 1 1 11894
0 11896 7 1 2 11878 11895
0 11897 7 1 2 11857 11896
0 11898 7 1 2 11776 11897
0 11899 5 1 1 11898
0 11900 7 1 2 25627 11899
0 11901 5 1 1 11900
0 11902 7 3 2 26949 30470
0 11903 7 2 2 23198 25440
0 11904 7 1 2 26457 36265
0 11905 7 1 2 36262 11904
0 11906 7 2 2 31424 33782
0 11907 7 3 2 27865 29420
0 11908 7 1 2 36267 36269
0 11909 7 1 2 11905 11908
0 11910 5 1 1 11909
0 11911 7 1 2 11901 11910
0 11912 5 1 1 11911
0 11913 7 1 2 27589 11912
0 11914 5 1 1 11913
0 11915 7 1 2 24969 36126
0 11916 5 1 1 11915
0 11917 7 8 2 23045 25561
0 11918 7 1 2 36272 36121
0 11919 5 1 1 11918
0 11920 7 1 2 11916 11919
0 11921 5 1 1 11920
0 11922 7 2 2 30601 11921
0 11923 7 1 2 36191 36280
0 11924 5 1 1 11923
0 11925 7 1 2 26950 36131
0 11926 7 1 2 34713 11925
0 11927 5 1 1 11926
0 11928 7 1 2 11924 11927
0 11929 5 1 1 11928
0 11930 7 1 2 31485 11929
0 11931 5 1 1 11930
0 11932 7 3 2 24897 25908
0 11933 7 1 2 33583 36282
0 11934 7 1 2 36132 11933
0 11935 7 1 2 36060 11934
0 11936 5 1 1 11935
0 11937 7 1 2 11931 11936
0 11938 7 1 2 28996 36281
0 11939 5 1 1 11938
0 11940 7 1 2 35822 35308
0 11941 7 1 2 36133 11940
0 11942 5 1 1 11941
0 11943 7 1 2 11939 11942
0 11944 5 1 1 11943
0 11945 7 1 2 30828 11944
0 11946 5 1 1 11945
0 11947 7 1 2 36122 31785
0 11948 5 1 1 11947
0 11949 7 2 2 23812 24279
0 11950 7 1 2 36285 27792
0 11951 7 1 2 33759 11950
0 11952 5 1 1 11951
0 11953 7 1 2 11948 11952
0 11954 5 1 1 11953
0 11955 7 1 2 25562 11954
0 11956 5 1 1 11955
0 11957 7 1 2 33395 32392
0 11958 7 1 2 33985 11957
0 11959 5 1 1 11958
0 11960 7 1 2 11956 11959
0 11961 5 1 1 11960
0 11962 7 1 2 36188 11961
0 11963 5 1 1 11962
0 11964 7 1 2 11946 11963
0 11965 7 1 2 11937 11964
0 11966 5 1 1 11965
0 11967 7 1 2 25704 11966
0 11968 5 1 1 11967
0 11969 7 3 2 27590 31081
0 11970 7 1 2 35591 36287
0 11971 5 1 1 11970
0 11972 7 1 2 24280 36108
0 11973 5 1 1 11972
0 11974 7 1 2 35956 32489
0 11975 5 1 1 11974
0 11976 7 1 2 11973 11975
0 11977 5 1 1 11976
0 11978 7 1 2 36115 11977
0 11979 5 1 1 11978
0 11980 7 1 2 11971 11979
0 11981 5 1 1 11980
0 11982 7 1 2 25563 11981
0 11983 5 1 1 11982
0 11984 7 1 2 26576 36117
0 11985 5 1 1 11984
0 11986 7 1 2 11983 11985
0 11987 5 1 1 11986
0 11988 7 1 2 36054 34391
0 11989 7 1 2 11987 11988
0 11990 5 1 1 11989
0 11991 7 1 2 11968 11990
0 11992 5 1 1 11991
0 11993 7 1 2 25628 11992
0 11994 5 1 1 11993
0 11995 7 1 2 35898 36011
0 11996 5 1 1 11995
0 11997 7 1 2 36128 11996
0 11998 5 1 1 11997
0 11999 7 1 2 31844 11998
0 12000 7 1 2 36104 11999
0 12001 5 1 1 12000
0 12002 7 1 2 23199 29921
0 12003 7 1 2 35720 12002
0 12004 7 2 2 24772 32611
0 12005 7 1 2 33737 36290
0 12006 7 1 2 12003 12005
0 12007 5 1 1 12006
0 12008 7 1 2 12001 12007
0 12009 5 1 1 12008
0 12010 7 1 2 33486 12009
0 12011 5 1 1 12010
0 12012 7 2 2 24281 35751
0 12013 7 1 2 33469 36292
0 12014 5 1 1 12013
0 12015 7 2 2 24898 29356
0 12016 7 1 2 24282 5860
0 12017 5 1 1 12016
0 12018 7 1 2 36294 12017
0 12019 5 1 1 12018
0 12020 7 1 2 12014 12019
0 12021 5 1 1 12020
0 12022 7 2 2 35721 30113
0 12023 7 1 2 33760 36234
0 12024 7 1 2 33839 12023
0 12025 7 1 2 36296 12024
0 12026 7 1 2 12021 12025
0 12027 5 1 1 12026
0 12028 7 1 2 12011 12027
0 12029 7 1 2 11994 12028
0 12030 5 1 1 12029
0 12031 7 1 2 22358 12030
0 12032 5 1 1 12031
0 12033 7 1 2 26351 30910
0 12034 5 1 1 12033
0 12035 7 2 2 25909 29956
0 12036 7 1 2 36291 36298
0 12037 5 1 1 12036
0 12038 7 1 2 12034 12037
0 12039 5 1 1 12038
0 12040 7 1 2 32378 12039
0 12041 5 1 1 12040
0 12042 7 1 2 36038 32001
0 12043 7 1 2 36186 12042
0 12044 5 1 1 12043
0 12045 7 1 2 12041 12044
0 12046 5 1 1 12045
0 12047 7 1 2 25997 12046
0 12048 5 1 1 12047
0 12049 7 1 2 27807 36025
0 12050 7 1 2 36029 12049
0 12051 5 1 1 12050
0 12052 7 2 2 36031 12051
0 12053 5 1 1 36300
0 12054 7 1 2 31486 36301
0 12055 5 1 1 12054
0 12056 7 2 2 28997 30479
0 12057 7 1 2 26541 27819
0 12058 7 1 2 36302 12057
0 12059 5 1 1 12058
0 12060 7 1 2 24773 36183
0 12061 5 1 1 12060
0 12062 7 1 2 29979 26352
0 12063 5 1 1 12062
0 12064 7 1 2 12061 12063
0 12065 5 1 1 12064
0 12066 7 1 2 36048 12065
0 12067 5 1 1 12066
0 12068 7 1 2 12059 12067
0 12069 7 1 2 12055 12068
0 12070 5 1 1 12069
0 12071 7 1 2 26951 12070
0 12072 5 1 1 12071
0 12073 7 1 2 12048 12072
0 12074 5 1 1 12073
0 12075 7 1 2 25564 12074
0 12076 5 1 1 12075
0 12077 7 1 2 24899 36093
0 12078 5 1 1 12077
0 12079 7 1 2 34267 12078
0 12080 5 2 1 12079
0 12081 7 1 2 36304 36189
0 12082 5 1 1 12081
0 12083 7 1 2 22962 36197
0 12084 5 1 1 12083
0 12085 7 1 2 12082 12084
0 12086 7 1 2 12076 12085
0 12087 5 1 1 12086
0 12088 7 2 2 33638 31845
0 12089 7 1 2 33649 36306
0 12090 7 1 2 12087 12089
0 12091 5 1 1 12090
0 12092 7 1 2 12032 12091
0 12093 5 1 1 12092
0 12094 7 1 2 29228 12093
0 12095 5 1 1 12094
0 12096 7 1 2 29035 36293
0 12097 5 1 1 12096
0 12098 7 1 2 24283 26559
0 12099 5 1 1 12098
0 12100 7 1 2 36295 12099
0 12101 5 1 1 12100
0 12102 7 1 2 12097 12101
0 12103 5 1 1 12102
0 12104 7 1 2 34175 36259
0 12105 7 1 2 27834 12104
0 12106 7 1 2 36268 12105
0 12107 7 1 2 36297 12106
0 12108 7 1 2 12103 12107
0 12109 5 1 1 12108
0 12110 7 1 2 12095 12109
0 12111 7 1 2 11914 12110
0 12112 7 1 2 11679 12111
0 12113 5 1 1 12112
0 12114 7 1 2 32107 12113
0 12115 5 1 1 12114
0 12116 7 1 2 22359 34818
0 12117 5 1 1 12116
0 12118 7 2 2 23417 33592
0 12119 7 2 2 36308 34509
0 12120 5 1 1 36310
0 12121 7 1 2 23269 36311
0 12122 5 1 1 12121
0 12123 7 1 2 12117 12122
0 12124 5 1 1 12123
0 12125 7 1 2 27316 12124
0 12126 5 2 1 12125
0 12127 7 1 2 22474 36199
0 12128 5 1 1 12127
0 12129 7 1 2 31163 33986
0 12130 5 1 1 12129
0 12131 7 1 2 12128 12130
0 12132 5 2 1 12131
0 12133 7 1 2 22360 36314
0 12134 5 1 1 12133
0 12135 7 2 2 31836 33639
0 12136 5 1 1 36316
0 12137 7 1 2 22475 36317
0 12138 5 1 1 12137
0 12139 7 1 2 12134 12138
0 12140 5 1 1 12139
0 12141 7 1 2 34137 12140
0 12142 5 1 1 12141
0 12143 7 1 2 36312 12142
0 12144 5 1 1 12143
0 12145 7 2 2 23813 12144
0 12146 5 2 1 36318
0 12147 7 1 2 24970 36319
0 12148 5 1 1 12147
0 12149 7 1 2 22361 27413
0 12150 7 1 2 36273 36154
0 12151 7 1 2 12149 12150
0 12152 7 1 2 32316 12151
0 12153 5 2 1 12152
0 12154 7 1 2 12148 36322
0 12155 5 2 1 12154
0 12156 7 1 2 35020 36324
0 12157 5 1 1 12156
0 12158 7 1 2 35470 34465
0 12159 5 1 1 12158
0 12160 7 9 2 27973 34326
0 12161 7 1 2 34168 36326
0 12162 5 1 1 12161
0 12163 7 1 2 12159 12162
0 12164 5 4 1 12163
0 12165 7 1 2 35563 35252
0 12166 5 1 1 12165
0 12167 7 1 2 24971 35016
0 12168 5 1 1 12167
0 12169 7 1 2 12166 12168
0 12170 5 1 1 12169
0 12171 7 2 2 36335 12170
0 12172 7 1 2 27215 36339
0 12173 5 1 1 12172
0 12174 7 1 2 12157 12173
0 12175 5 1 1 12174
0 12176 7 1 2 30602 12175
0 12177 5 1 1 12176
0 12178 7 1 2 23814 34819
0 12179 5 1 1 12178
0 12180 7 1 2 31858 36155
0 12181 7 1 2 34192 12180
0 12182 5 1 1 12181
0 12183 7 1 2 12179 12182
0 12184 5 1 1 12183
0 12185 7 1 2 22362 12184
0 12186 5 1 1 12185
0 12187 7 1 2 35886 34181
0 12188 5 1 1 12187
0 12189 7 1 2 12186 12188
0 12190 5 1 1 12189
0 12191 7 1 2 27317 12190
0 12192 5 1 1 12191
0 12193 7 2 2 34125 34327
0 12194 5 1 1 36341
0 12195 7 1 2 27866 36342
0 12196 5 1 1 12195
0 12197 7 1 2 34188 34547
0 12198 5 1 1 12197
0 12199 7 1 2 12196 12198
0 12200 5 1 1 12199
0 12201 7 1 2 23936 12200
0 12202 5 1 1 12201
0 12203 7 1 2 35882 34466
0 12204 5 2 1 12203
0 12205 7 1 2 12202 36343
0 12206 7 1 2 12192 12205
0 12207 5 2 1 12206
0 12208 7 1 2 28998 35564
0 12209 7 1 2 36049 12208
0 12210 7 1 2 36345 12209
0 12211 5 1 1 12210
0 12212 7 1 2 12177 12211
0 12213 5 1 1 12212
0 12214 7 1 2 31487 12213
0 12215 5 1 1 12214
0 12216 7 1 2 34788 26353
0 12217 5 1 1 12216
0 12218 7 1 2 26847 36184
0 12219 5 1 1 12218
0 12220 7 1 2 12217 12219
0 12221 5 1 1 12220
0 12222 7 1 2 36346 12221
0 12223 5 1 1 12222
0 12224 7 1 2 22363 36200
0 12225 5 1 1 12224
0 12226 7 1 2 12136 12225
0 12227 5 1 1 12226
0 12228 7 1 2 12227 34210
0 12229 5 1 1 12228
0 12230 7 1 2 36309 34500
0 12231 5 1 1 12230
0 12232 7 1 2 12231 6283
0 12233 5 1 1 12232
0 12234 7 1 2 22364 12233
0 12235 5 1 1 12234
0 12236 7 1 2 12120 12235
0 12237 5 1 1 12236
0 12238 7 1 2 31164 12237
0 12239 5 1 1 12238
0 12240 7 1 2 27318 34138
0 12241 7 1 2 34467 12240
0 12242 5 1 1 12241
0 12243 7 1 2 12239 12242
0 12244 7 1 2 12229 12243
0 12245 5 1 1 12244
0 12246 7 1 2 25805 12245
0 12247 5 1 1 12246
0 12248 7 1 2 23200 33882
0 12249 5 1 1 12248
0 12250 7 2 2 35247 34279
0 12251 5 1 1 36347
0 12252 7 1 2 12249 12251
0 12253 5 3 1 12252
0 12254 7 1 2 22624 36349
0 12255 5 1 1 12254
0 12256 7 1 2 35465 33961
0 12257 5 1 1 12256
0 12258 7 1 2 12255 12257
0 12259 5 1 1 12258
0 12260 7 1 2 22476 12259
0 12261 5 1 1 12260
0 12262 7 1 2 32856 33987
0 12263 5 1 1 12262
0 12264 7 1 2 12261 12263
0 12265 5 1 1 12264
0 12266 7 1 2 22365 12265
0 12267 5 1 1 12266
0 12268 7 1 2 34183 12267
0 12269 5 1 1 12268
0 12270 7 1 2 27237 12269
0 12271 5 1 1 12270
0 12272 7 1 2 12247 12271
0 12273 5 1 1 12272
0 12274 7 1 2 35048 35171
0 12275 7 1 2 12273 12274
0 12276 5 1 1 12275
0 12277 7 1 2 12223 12276
0 12278 5 1 1 12277
0 12279 7 1 2 34710 12278
0 12280 5 1 1 12279
0 12281 7 1 2 36313 7517
0 12282 5 1 1 12281
0 12283 7 1 2 23815 12282
0 12284 5 1 1 12283
0 12285 7 1 2 34766 34829
0 12286 5 1 1 12285
0 12287 7 1 2 12194 12286
0 12288 5 1 1 12287
0 12289 7 1 2 34403 12288
0 12290 5 1 1 12289
0 12291 7 1 2 36344 12290
0 12292 7 1 2 12284 12291
0 12293 5 1 1 12292
0 12294 7 1 2 24972 12293
0 12295 5 1 1 12294
0 12296 7 1 2 36323 12295
0 12297 5 1 1 12296
0 12298 7 1 2 35522 12297
0 12299 5 1 1 12298
0 12300 7 2 2 1491 1116
0 12301 7 1 2 32222 34074
0 12302 7 1 2 36352 12301
0 12303 7 1 2 31210 12302
0 12304 7 1 2 36336 12303
0 12305 5 1 1 12304
0 12306 7 1 2 12299 12305
0 12307 5 1 1 12306
0 12308 7 1 2 36023 12307
0 12309 5 1 1 12308
0 12310 7 1 2 12280 12309
0 12311 7 1 2 12215 12310
0 12312 7 1 2 35851 26848
0 12313 5 1 1 12312
0 12314 7 1 2 35018 12313
0 12315 5 1 1 12314
0 12316 7 1 2 27216 12315
0 12317 7 2 2 36337 12316
0 12318 5 1 1 36354
0 12319 7 1 2 25910 32060
0 12320 7 1 2 32700 12319
0 12321 7 4 2 24462 33331
0 12322 7 1 2 32310 36356
0 12323 7 1 2 12320 12322
0 12324 5 1 1 12323
0 12325 7 1 2 36320 12324
0 12326 5 2 1 12325
0 12327 7 1 2 35021 36360
0 12328 5 1 1 12327
0 12329 7 1 2 12318 12328
0 12330 5 1 1 12329
0 12331 7 1 2 28512 31218
0 12332 7 1 2 12330 12331
0 12333 5 1 1 12332
0 12334 7 2 2 31635 36123
0 12335 7 1 2 34789 36362
0 12336 5 1 1 12335
0 12337 7 1 2 30396 33988
0 12338 7 1 2 33871 12337
0 12339 5 1 1 12338
0 12340 7 1 2 12336 12339
0 12341 5 1 1 12340
0 12342 7 1 2 22963 12341
0 12343 5 1 1 12342
0 12344 7 3 2 35879 31437
0 12345 5 1 1 36364
0 12346 7 1 2 36365 36363
0 12347 5 1 1 12346
0 12348 7 1 2 12343 12347
0 12349 5 1 1 12348
0 12350 7 1 2 32849 12349
0 12351 5 1 1 12350
0 12352 7 1 2 28273 34959
0 12353 7 1 2 36263 12352
0 12354 7 7 2 23124 23201
0 12355 7 4 2 22964 36367
0 12356 7 1 2 36374 30758
0 12357 7 1 2 12353 12356
0 12358 5 1 1 12357
0 12359 7 1 2 12351 12358
0 12360 5 1 1 12359
0 12361 7 1 2 22366 12360
0 12362 5 1 1 12361
0 12363 7 1 2 35524 12345
0 12364 5 2 1 12363
0 12365 7 1 2 34539 36378
0 12366 5 1 1 12365
0 12367 7 5 2 22625 22965
0 12368 7 1 2 36221 36380
0 12369 7 1 2 36264 12368
0 12370 5 1 1 12369
0 12371 7 1 2 12366 12370
0 12372 5 1 1 12371
0 12373 7 1 2 34468 12372
0 12374 5 1 1 12373
0 12375 7 1 2 27974 34767
0 12376 7 1 2 30287 32173
0 12377 7 1 2 12375 12376
0 12378 5 1 1 12377
0 12379 7 1 2 12374 12378
0 12380 5 1 1 12379
0 12381 7 1 2 32246 12380
0 12382 5 1 1 12381
0 12383 7 1 2 22367 36350
0 12384 5 1 1 12383
0 12385 7 1 2 32158 33644
0 12386 5 1 1 12385
0 12387 7 1 2 12384 12386
0 12388 5 1 1 12387
0 12389 7 1 2 34837 5980
0 12390 5 1 1 12389
0 12391 7 1 2 30397 12390
0 12392 5 1 1 12391
0 12393 7 2 2 25806 28344
0 12394 7 1 2 27613 36385
0 12395 7 1 2 31446 12394
0 12396 5 1 1 12395
0 12397 7 1 2 12392 12396
0 12398 5 1 1 12397
0 12399 7 1 2 22966 12398
0 12400 5 1 1 12399
0 12401 7 1 2 36366 33886
0 12402 5 1 1 12401
0 12403 7 1 2 12400 12402
0 12404 5 1 1 12403
0 12405 7 1 2 12388 12404
0 12406 5 1 1 12405
0 12407 7 1 2 22626 27217
0 12408 7 1 2 33640 12407
0 12409 7 1 2 33316 12408
0 12410 7 1 2 36379 12409
0 12411 5 1 1 12410
0 12412 7 1 2 12406 12411
0 12413 7 1 2 12382 12412
0 12414 7 1 2 12362 12413
0 12415 5 1 1 12414
0 12416 7 1 2 28999 12415
0 12417 5 1 1 12416
0 12418 7 1 2 34994 36361
0 12419 5 1 1 12418
0 12420 7 1 2 26086 36355
0 12421 5 1 1 12420
0 12422 7 1 2 12419 12421
0 12423 5 1 1 12422
0 12424 7 1 2 29666 12423
0 12425 5 1 1 12424
0 12426 7 1 2 12417 12425
0 12427 7 1 2 12333 12426
0 12428 5 1 1 12427
0 12429 7 1 2 33487 12428
0 12430 5 1 1 12429
0 12431 7 1 2 36325 36087
0 12432 5 1 1 12431
0 12433 7 1 2 23937 36338
0 12434 5 1 1 12433
0 12435 7 3 2 22368 31195
0 12436 7 1 2 36387 31906
0 12437 7 1 2 34835 12436
0 12438 5 1 1 12437
0 12439 7 1 2 12434 12438
0 12440 5 1 1 12439
0 12441 7 1 2 25807 12440
0 12442 5 1 1 12441
0 12443 7 1 2 36321 12442
0 12444 5 1 1 12443
0 12445 7 1 2 12444 34266
0 12446 5 1 1 12445
0 12447 7 1 2 12432 12446
0 12448 5 1 1 12447
0 12449 7 1 2 34995 12448
0 12450 5 1 1 12449
0 12451 7 1 2 33011 34634
0 12452 7 1 2 36340 12451
0 12453 5 1 1 12452
0 12454 7 1 2 12450 12453
0 12455 5 1 1 12454
0 12456 7 1 2 28655 12455
0 12457 5 1 1 12456
0 12458 7 1 2 12430 12457
0 12459 7 1 2 12311 12458
0 12460 5 1 1 12459
0 12461 7 1 2 25705 12460
0 12462 5 1 1 12461
0 12463 7 4 2 34886 27614
0 12464 7 1 2 36101 36390
0 12465 5 1 1 12464
0 12466 7 2 2 27591 34996
0 12467 7 1 2 26165 35551
0 12468 7 2 2 36394 12467
0 12469 5 1 1 36396
0 12470 7 1 2 12465 12469
0 12471 5 1 1 12470
0 12472 7 1 2 24900 12471
0 12473 5 1 1 12472
0 12474 7 1 2 26805 35552
0 12475 7 2 2 36395 12474
0 12476 5 1 1 36398
0 12477 7 1 2 12473 12476
0 12478 5 1 1 12477
0 12479 7 1 2 23351 32419
0 12480 7 2 2 12478 12479
0 12481 7 1 2 31170 36400
0 12482 5 1 1 12481
0 12483 7 2 2 24901 29036
0 12484 7 1 2 33775 36402
0 12485 5 1 1 12484
0 12486 7 1 2 30363 27641
0 12487 5 1 1 12486
0 12488 7 1 2 35007 35478
0 12489 5 1 1 12488
0 12490 7 1 2 12487 12489
0 12491 5 1 1 12490
0 12492 7 1 2 25565 12491
0 12493 5 1 1 12492
0 12494 7 1 2 12485 12493
0 12495 5 1 1 12494
0 12496 7 1 2 35011 12495
0 12497 5 1 1 12496
0 12498 7 1 2 35982 11165
0 12499 5 1 1 12498
0 12500 7 1 2 24902 29289
0 12501 7 1 2 35275 12500
0 12502 5 1 1 12501
0 12503 7 1 2 12499 12502
0 12504 5 1 1 12503
0 12505 7 1 2 26087 12504
0 12506 5 1 1 12505
0 12507 7 1 2 26606 27513
0 12508 5 1 1 12507
0 12509 7 1 2 12506 12508
0 12510 5 1 1 12509
0 12511 7 1 2 23549 12510
0 12512 5 1 1 12511
0 12513 7 1 2 26785 1928
0 12514 5 1 1 12513
0 12515 7 1 2 26565 12514
0 12516 5 1 1 12515
0 12517 7 2 2 24973 29070
0 12518 5 1 1 36404
0 12519 7 1 2 32986 36405
0 12520 5 1 1 12519
0 12521 7 1 2 12516 12520
0 12522 5 1 1 12521
0 12523 7 1 2 25566 12522
0 12524 5 1 1 12523
0 12525 7 1 2 26254 29654
0 12526 5 1 1 12525
0 12527 7 1 2 12524 12526
0 12528 5 1 1 12527
0 12529 7 1 2 26088 12528
0 12530 5 1 1 12529
0 12531 7 1 2 12512 12530
0 12532 5 1 1 12531
0 12533 7 1 2 24027 12532
0 12534 5 1 1 12533
0 12535 7 1 2 35880 36391
0 12536 5 1 1 12535
0 12537 7 1 2 12534 12536
0 12538 5 1 1 12537
0 12539 7 1 2 23477 12538
0 12540 5 1 1 12539
0 12541 7 1 2 12497 12540
0 12542 5 1 1 12541
0 12543 7 1 2 27288 12542
0 12544 5 1 1 12543
0 12545 7 1 2 34982 36288
0 12546 5 1 1 12545
0 12547 7 3 2 26760 35119
0 12548 7 2 2 25998 32456
0 12549 7 1 2 36406 36409
0 12550 5 1 1 12549
0 12551 7 1 2 12546 12550
0 12552 5 1 1 12551
0 12553 7 1 2 25567 12552
0 12554 5 1 1 12553
0 12555 7 3 2 27615 36050
0 12556 5 1 1 36411
0 12557 7 1 2 36412 36410
0 12558 5 1 1 12557
0 12559 7 1 2 12554 12558
0 12560 5 1 1 12559
0 12561 7 1 2 27023 12560
0 12562 5 1 1 12561
0 12563 7 1 2 22843 12562
0 12564 7 1 2 12544 12563
0 12565 5 1 1 12564
0 12566 7 1 2 23352 33804
0 12567 5 1 1 12566
0 12568 7 1 2 12567 11411
0 12569 5 1 1 12568
0 12570 7 1 2 36392 12569
0 12571 5 1 1 12570
0 12572 7 1 2 27319 27592
0 12573 7 2 2 32457 12572
0 12574 7 1 2 36172 36414
0 12575 5 1 1 12574
0 12576 7 1 2 12571 12575
0 12577 5 1 1 12576
0 12578 7 1 2 24903 12577
0 12579 5 1 1 12578
0 12580 7 1 2 26806 35565
0 12581 7 1 2 36415 12580
0 12582 5 1 1 12581
0 12583 7 1 2 24774 12582
0 12584 7 1 2 12579 12583
0 12585 5 1 1 12584
0 12586 7 1 2 30980 12585
0 12587 7 1 2 12565 12586
0 12588 5 1 1 12587
0 12589 7 3 2 25999 32490
0 12590 7 1 2 36413 36416
0 12591 5 1 1 12590
0 12592 7 2 2 34997 36289
0 12593 5 1 1 36419
0 12594 7 1 2 36407 36417
0 12595 5 1 1 12594
0 12596 7 1 2 12593 12595
0 12597 5 1 1 12596
0 12598 7 1 2 25568 12597
0 12599 5 1 1 12598
0 12600 7 1 2 12591 12599
0 12601 5 1 1 12600
0 12602 7 1 2 35873 12601
0 12603 5 1 1 12602
0 12604 7 1 2 23816 12603
0 12605 7 1 2 12588 12604
0 12606 5 1 1 12605
0 12607 7 1 2 25308 36102
0 12608 5 1 1 12607
0 12609 7 1 2 33538 27425
0 12610 5 1 1 12609
0 12611 7 1 2 12608 12610
0 12612 5 1 1 12611
0 12613 7 1 2 31015 12612
0 12614 5 1 1 12613
0 12615 7 1 2 24775 27755
0 12616 7 1 2 28010 12615
0 12617 7 1 2 33539 12616
0 12618 5 1 1 12617
0 12619 7 1 2 12614 12618
0 12620 5 1 1 12619
0 12621 7 1 2 36393 12620
0 12622 5 1 1 12621
0 12623 7 1 2 34512 36397
0 12624 5 1 1 12623
0 12625 7 1 2 12622 12624
0 12626 5 1 1 12625
0 12627 7 1 2 24904 12626
0 12628 5 1 1 12627
0 12629 7 1 2 34513 36399
0 12630 5 1 1 12629
0 12631 7 1 2 25808 12630
0 12632 7 1 2 12628 12631
0 12633 5 1 1 12632
0 12634 7 1 2 12606 12633
0 12635 5 1 1 12634
0 12636 7 1 2 22627 12635
0 12637 5 1 1 12636
0 12638 7 1 2 25569 36408
0 12639 5 1 1 12638
0 12640 7 1 2 12556 12639
0 12641 5 1 1 12640
0 12642 7 1 2 30981 27259
0 12643 5 1 1 12642
0 12644 7 2 2 25378 27218
0 12645 7 1 2 28876 36421
0 12646 5 1 1 12645
0 12647 7 1 2 12643 12646
0 12648 5 2 1 12647
0 12649 7 1 2 36418 36423
0 12650 5 1 1 12649
0 12651 7 1 2 35172 31333
0 12652 7 1 2 35875 12651
0 12653 5 1 1 12652
0 12654 7 1 2 12650 12653
0 12655 5 1 1 12654
0 12656 7 1 2 12641 12655
0 12657 5 1 1 12656
0 12658 7 1 2 25570 36424
0 12659 7 1 2 36420 12658
0 12660 5 1 1 12659
0 12661 7 1 2 24594 12660
0 12662 7 1 2 12657 12661
0 12663 5 1 1 12662
0 12664 7 1 2 23270 12663
0 12665 7 1 2 12637 12664
0 12666 5 1 1 12665
0 12667 7 1 2 12482 12666
0 12668 5 1 1 12667
0 12669 7 1 2 22477 12668
0 12670 5 1 1 12669
0 12671 7 1 2 36401 30661
0 12672 5 1 1 12671
0 12673 7 1 2 12670 12672
0 12674 5 1 1 12673
0 12675 7 3 2 25074 23705
0 12676 7 1 2 32061 36425
0 12677 7 1 2 12674 12676
0 12678 5 1 1 12677
0 12679 7 1 2 12462 12678
0 12680 5 1 1 12679
0 12681 7 1 2 25629 12680
0 12682 5 1 1 12681
0 12683 7 1 2 32726 36039
0 12684 5 1 1 12683
0 12685 7 2 2 24284 29112
0 12686 7 1 2 35309 36428
0 12687 5 1 1 12686
0 12688 7 1 2 12684 12687
0 12689 5 1 1 12688
0 12690 7 1 2 25571 12689
0 12691 5 1 1 12690
0 12692 7 1 2 32727 36195
0 12693 5 1 1 12692
0 12694 7 1 2 12691 12693
0 12695 5 1 1 12694
0 12696 7 3 2 25630 33675
0 12697 7 1 2 12695 36430
0 12698 5 1 1 12697
0 12699 7 1 2 32393 33770
0 12700 5 1 1 12699
0 12701 7 4 2 25631 33457
0 12702 5 1 1 36433
0 12703 7 1 2 26469 12702
0 12704 5 1 1 12703
0 12705 7 1 2 23046 29071
0 12706 7 1 2 12704 12705
0 12707 5 1 1 12706
0 12708 7 1 2 12700 12707
0 12709 5 1 1 12708
0 12710 7 1 2 23478 12709
0 12711 5 1 1 12710
0 12712 7 1 2 24974 26708
0 12713 5 1 1 12712
0 12714 7 1 2 32718 12713
0 12715 5 1 1 12714
0 12716 7 1 2 32705 33559
0 12717 5 2 1 12716
0 12718 7 1 2 12715 36437
0 12719 5 1 1 12718
0 12720 7 1 2 35752 12719
0 12721 5 1 1 12720
0 12722 7 1 2 24285 12721
0 12723 7 1 2 12711 12722
0 12724 5 1 1 12723
0 12725 7 1 2 32728 34075
0 12726 5 1 1 12725
0 12727 7 1 2 29072 35310
0 12728 7 1 2 36434 12727
0 12729 5 1 1 12728
0 12730 7 1 2 26255 12729
0 12731 7 1 2 12726 12730
0 12732 5 1 1 12731
0 12733 7 1 2 33654 12732
0 12734 7 1 2 12724 12733
0 12735 5 1 1 12734
0 12736 7 1 2 12698 12735
0 12737 5 1 1 12736
0 12738 7 1 2 22844 12737
0 12739 5 1 1 12738
0 12740 7 1 2 23125 36431
0 12741 5 1 1 12740
0 12742 7 1 2 33667 12741
0 12743 5 1 1 12742
0 12744 7 1 2 33488 12743
0 12745 5 1 1 12744
0 12746 7 2 2 23706 24286
0 12747 7 2 2 36368 36439
0 12748 5 1 1 36441
0 12749 7 1 2 23635 36442
0 12750 5 1 1 12749
0 12751 7 1 2 36274 36432
0 12752 5 1 1 12751
0 12753 7 1 2 24975 33655
0 12754 5 1 1 12753
0 12755 7 1 2 12752 12754
0 12756 5 1 1 12755
0 12757 7 1 2 26256 12756
0 12758 5 1 1 12757
0 12759 7 1 2 12750 12758
0 12760 7 1 2 12745 12759
0 12761 5 1 1 12760
0 12762 7 1 2 35034 12761
0 12763 5 1 1 12762
0 12764 7 1 2 12739 12763
0 12765 5 1 1 12764
0 12766 7 1 2 24028 12765
0 12767 5 1 1 12766
0 12768 7 2 2 25572 34410
0 12769 7 1 2 29113 26577
0 12770 7 2 2 36443 12769
0 12771 5 1 1 36445
0 12772 7 2 2 27593 33656
0 12773 5 1 1 36447
0 12774 7 3 2 23126 33676
0 12775 5 1 1 36449
0 12776 7 1 2 27494 36450
0 12777 5 1 1 12776
0 12778 7 1 2 12773 12777
0 12779 5 1 1 12778
0 12780 7 1 2 25498 12779
0 12781 5 1 1 12780
0 12782 7 1 2 30714 7057
0 12783 7 1 2 36444 12782
0 12784 5 1 1 12783
0 12785 7 1 2 12781 12784
0 12786 5 1 1 12785
0 12787 7 1 2 24905 12786
0 12788 5 1 1 12787
0 12789 7 1 2 12771 12788
0 12790 5 1 1 12789
0 12791 7 1 2 35657 35012
0 12792 7 1 2 12790 12791
0 12793 5 1 1 12792
0 12794 7 1 2 26089 12793
0 12795 7 1 2 12767 12794
0 12796 5 1 1 12795
0 12797 7 1 2 34779 33657
0 12798 7 1 2 35507 12797
0 12799 5 1 1 12798
0 12800 7 1 2 29000 36446
0 12801 5 1 1 12800
0 12802 7 1 2 12799 12801
0 12803 5 1 1 12802
0 12804 7 1 2 26000 12803
0 12805 5 1 1 12804
0 12806 7 2 2 26458 35013
0 12807 5 1 1 36452
0 12808 7 1 2 22967 35994
0 12809 5 1 1 12808
0 12810 7 1 2 12807 12809
0 12811 5 1 1 12810
0 12812 7 1 2 22845 12811
0 12813 5 1 1 12812
0 12814 7 1 2 32729 26849
0 12815 5 1 1 12814
0 12816 7 1 2 12813 12815
0 12817 5 1 1 12816
0 12818 7 1 2 33677 36094
0 12819 7 1 2 12817 12818
0 12820 5 1 1 12819
0 12821 7 1 2 12805 12820
0 12822 5 1 1 12821
0 12823 7 1 2 25632 12822
0 12824 5 1 1 12823
0 12825 7 1 2 24105 12824
0 12826 5 1 1 12825
0 12827 7 1 2 26166 12826
0 12828 7 1 2 12796 12827
0 12829 5 1 1 12828
0 12830 7 1 2 29114 34087
0 12831 5 1 1 12830
0 12832 7 2 2 25573 31057
0 12833 7 1 2 27495 36454
0 12834 5 1 1 12833
0 12835 7 1 2 12831 12834
0 12836 5 1 1 12835
0 12837 7 1 2 24106 12836
0 12838 5 1 1 12837
0 12839 7 1 2 24287 35687
0 12840 7 1 2 36403 12839
0 12841 5 1 1 12840
0 12842 7 1 2 12838 12841
0 12843 5 1 1 12842
0 12844 7 1 2 29001 12843
0 12845 5 1 1 12844
0 12846 7 1 2 33233 33088
0 12847 5 1 1 12846
0 12848 7 2 2 25499 30709
0 12849 7 1 2 26354 30254
0 12850 7 1 2 36456 12849
0 12851 5 1 1 12850
0 12852 7 1 2 12847 12851
0 12853 5 1 1 12852
0 12854 7 1 2 34076 12853
0 12855 5 1 1 12854
0 12856 7 1 2 29090 33565
0 12857 5 1 1 12856
0 12858 7 1 2 26897 32399
0 12859 7 1 2 12518 12858
0 12860 7 1 2 12857 12859
0 12861 5 1 1 12860
0 12862 7 1 2 12855 12861
0 12863 7 1 2 12845 12862
0 12864 5 1 1 12863
0 12865 7 1 2 33658 12864
0 12866 5 1 1 12865
0 12867 7 1 2 24107 28967
0 12868 5 1 1 12867
0 12869 7 1 2 33927 12868
0 12870 5 1 1 12869
0 12871 7 1 2 29115 36040
0 12872 5 1 1 12871
0 12873 7 1 2 23550 31752
0 12874 5 1 1 12873
0 12875 7 1 2 12872 12874
0 12876 5 1 1 12875
0 12877 7 1 2 25574 12876
0 12878 5 1 1 12877
0 12879 7 1 2 28552 36429
0 12880 5 1 1 12879
0 12881 7 1 2 12878 12880
0 12882 5 2 1 12881
0 12883 7 1 2 12870 36458
0 12884 5 1 1 12883
0 12885 7 1 2 26459 26578
0 12886 7 1 2 32464 12885
0 12887 5 1 1 12886
0 12888 7 1 2 32706 32400
0 12889 7 1 2 35067 12888
0 12890 5 1 1 12889
0 12891 7 1 2 12887 12890
0 12892 5 1 1 12891
0 12893 7 1 2 25575 12892
0 12894 5 1 1 12893
0 12895 7 1 2 12884 12894
0 12896 5 1 1 12895
0 12897 7 1 2 33678 12896
0 12898 5 1 1 12897
0 12899 7 1 2 12866 12898
0 12900 5 1 1 12899
0 12901 7 1 2 26001 12900
0 12902 5 1 1 12901
0 12903 7 1 2 36448 36455
0 12904 5 1 1 12903
0 12905 7 1 2 33679 36459
0 12906 5 1 1 12905
0 12907 7 1 2 12904 12906
0 12908 5 1 1 12907
0 12909 7 1 2 34162 12908
0 12910 5 1 1 12909
0 12911 7 1 2 12902 12910
0 12912 5 1 1 12911
0 12913 7 1 2 25633 24192
0 12914 7 1 2 12912 12913
0 12915 5 1 1 12914
0 12916 7 1 2 12829 12915
0 12917 5 1 1 12916
0 12918 7 1 2 22369 12917
0 12919 5 1 1 12918
0 12920 7 1 2 26002 12053
0 12921 5 1 1 12920
0 12922 7 1 2 24029 11156
0 12923 5 1 1 12922
0 12924 7 1 2 25576 12923
0 12925 7 1 2 12921 12924
0 12926 5 1 1 12925
0 12927 7 1 2 27496 27636
0 12928 7 1 2 35022 12927
0 12929 5 1 1 12928
0 12930 7 1 2 12926 12929
0 12931 5 1 1 12930
0 12932 7 1 2 31488 12931
0 12933 5 1 1 12932
0 12934 7 1 2 26807 34998
0 12935 7 1 2 36305 12934
0 12936 5 1 1 12935
0 12937 7 1 2 36095 34831
0 12938 5 1 1 12937
0 12939 7 1 2 26355 34711
0 12940 5 1 1 12939
0 12941 7 1 2 12938 12940
0 12942 5 1 1 12941
0 12943 7 1 2 34790 12942
0 12944 5 1 1 12943
0 12945 7 1 2 24976 32715
0 12946 7 1 2 35806 12945
0 12947 7 1 2 33440 12946
0 12948 5 1 1 12947
0 12949 7 1 2 12944 12948
0 12950 7 1 2 12936 12949
0 12951 7 1 2 12933 12950
0 12952 5 1 1 12951
0 12953 7 1 2 12952 36307
0 12954 5 1 1 12953
0 12955 7 1 2 12919 12954
0 12956 5 1 1 12955
0 12957 7 1 2 28706 12956
0 12958 5 1 1 12957
0 12959 7 3 2 29037 35416
0 12960 7 1 2 25634 35054
0 12961 7 1 2 32062 12960
0 12962 7 1 2 36460 12961
0 12963 7 1 2 34648 12962
0 12964 5 1 1 12963
0 12965 7 1 2 12958 12964
0 12966 5 1 1 12965
0 12967 7 1 2 32915 12966
0 12968 5 1 1 12967
0 12969 7 1 2 12682 12968
0 12970 7 1 2 12115 12969
0 12971 5 1 1 12970
0 12972 7 1 2 24331 12971
0 12973 5 1 1 12972
0 12974 7 1 2 36007 33641
0 12975 5 1 1 12974
0 12976 7 1 2 31394 34822
0 12977 5 1 1 12976
0 12978 7 2 2 32779 29400
0 12979 7 1 2 35678 34690
0 12980 7 1 2 36463 12979
0 12981 5 1 1 12980
0 12982 7 1 2 12977 12981
0 12983 5 1 1 12982
0 12984 7 1 2 26356 12983
0 12985 5 1 1 12984
0 12986 7 2 2 25809 35679
0 12987 7 1 2 25126 34620
0 12988 7 1 2 34386 12987
0 12989 7 1 2 36465 12988
0 12990 5 1 1 12989
0 12991 7 1 2 12985 12990
0 12992 5 1 1 12991
0 12993 7 1 2 23938 12992
0 12994 5 1 1 12993
0 12995 7 1 2 28892 35354
0 12996 7 1 2 31345 34691
0 12997 7 1 2 12995 12996
0 12998 7 1 2 31724 12997
0 12999 5 1 1 12998
0 13000 7 1 2 12994 12999
0 13001 5 1 1 13000
0 13002 7 1 2 24193 34077
0 13003 7 1 2 13001 13002
0 13004 5 1 1 13003
0 13005 7 1 2 28260 26357
0 13006 7 1 2 33560 33659
0 13007 7 1 2 13005 13006
0 13008 7 1 2 35961 13007
0 13009 5 1 1 13008
0 13010 7 1 2 13004 13009
0 13011 5 1 1 13010
0 13012 7 1 2 22741 13011
0 13013 5 1 1 13012
0 13014 7 3 2 24194 34088
0 13015 7 2 2 25810 36467
0 13016 7 2 2 25127 36470
0 13017 7 1 2 36472 29464
0 13018 7 1 2 27011 13017
0 13019 5 1 1 13018
0 13020 7 1 2 13013 13019
0 13021 5 1 1 13020
0 13022 7 1 2 23353 13021
0 13023 5 1 1 13022
0 13024 7 1 2 31409 31346
0 13025 5 1 1 13024
0 13026 7 1 2 35408 31283
0 13027 5 1 1 13026
0 13028 7 1 2 13025 13027
0 13029 5 1 1 13028
0 13030 7 1 2 26003 13029
0 13031 5 1 1 13030
0 13032 7 1 2 33187 31875
0 13033 5 1 1 13032
0 13034 7 1 2 13031 13033
0 13035 5 1 1 13034
0 13036 7 2 2 25309 33680
0 13037 7 1 2 33720 36474
0 13038 7 1 2 36468 13037
0 13039 7 1 2 13035 13038
0 13040 5 1 1 13039
0 13041 7 1 2 13023 13040
0 13042 5 1 1 13041
0 13043 7 1 2 22628 13042
0 13044 5 1 1 13043
0 13045 7 1 2 27135 35760
0 13046 5 1 1 13045
0 13047 7 1 2 31585 27084
0 13048 5 1 1 13047
0 13049 7 1 2 13046 13048
0 13050 5 1 1 13049
0 13051 7 1 2 25911 13050
0 13052 5 1 1 13051
0 13053 7 1 2 31414 33109
0 13054 5 1 1 13053
0 13055 7 1 2 13052 13054
0 13056 5 1 1 13055
0 13057 7 1 2 25706 34568
0 13058 7 1 2 36473 13057
0 13059 7 1 2 13056 13058
0 13060 5 1 1 13059
0 13061 7 1 2 13044 13060
0 13062 5 1 1 13061
0 13063 7 1 2 22478 13062
0 13064 5 1 1 13063
0 13065 7 1 2 32803 33972
0 13066 5 1 1 13065
0 13067 7 1 2 34280 31967
0 13068 7 1 2 32890 13067
0 13069 5 1 1 13068
0 13070 7 1 2 13066 13069
0 13071 5 1 1 13070
0 13072 7 1 2 28732 13071
0 13073 5 1 1 13072
0 13074 7 1 2 32599 34813
0 13075 5 1 1 13074
0 13076 7 1 2 26973 31196
0 13077 7 1 2 33962 13076
0 13078 5 1 1 13077
0 13079 7 1 2 13075 13078
0 13080 5 1 1 13079
0 13081 7 1 2 28825 13080
0 13082 5 1 1 13081
0 13083 7 4 2 25128 28362
0 13084 7 2 2 28817 36476
0 13085 5 1 1 36480
0 13086 7 3 2 24776 33963
0 13087 7 1 2 31992 36482
0 13088 5 1 1 13087
0 13089 7 1 2 13085 13088
0 13090 5 1 1 13089
0 13091 7 1 2 32963 13090
0 13092 5 1 1 13091
0 13093 7 1 2 13082 13092
0 13094 7 1 2 13073 13093
0 13095 5 1 1 13094
0 13096 7 1 2 36471 34605
0 13097 7 1 2 13095 13096
0 13098 5 1 1 13097
0 13099 7 1 2 13064 13098
0 13100 5 1 1 13099
0 13101 7 1 2 22370 13100
0 13102 5 1 1 13101
0 13103 7 1 2 36469 33729
0 13104 7 1 2 33051 13103
0 13105 5 1 1 13104
0 13106 7 1 2 13102 13105
0 13107 5 1 1 13106
0 13108 7 1 2 26090 13107
0 13109 5 1 1 13108
0 13110 7 1 2 29170 34328
0 13111 5 1 1 13110
0 13112 7 1 2 32063 31768
0 13113 5 1 1 13112
0 13114 7 1 2 13111 13113
0 13115 5 1 1 13114
0 13116 7 1 2 34026 13115
0 13117 5 1 1 13116
0 13118 7 1 2 35946 34329
0 13119 5 1 1 13118
0 13120 7 1 2 13117 13119
0 13121 5 1 1 13120
0 13122 7 3 2 25075 34078
0 13123 7 2 2 25707 28707
0 13124 7 1 2 36485 36488
0 13125 7 1 2 36303 13124
0 13126 7 1 2 13121 13125
0 13127 5 1 1 13126
0 13128 7 1 2 13109 13127
0 13129 5 1 1 13128
0 13130 7 1 2 29116 13129
0 13131 5 1 1 13130
0 13132 7 3 2 25708 26257
0 13133 7 2 2 27808 36490
0 13134 7 1 2 35148 34447
0 13135 5 1 1 13134
0 13136 7 1 2 25129 26982
0 13137 7 1 2 29171 13136
0 13138 5 1 1 13137
0 13139 7 1 2 13135 13138
0 13140 5 1 1 13139
0 13141 7 1 2 29539 13140
0 13142 5 1 1 13141
0 13143 7 1 2 24595 32266
0 13144 5 1 1 13143
0 13145 7 2 2 25310 29520
0 13146 7 1 2 30387 36495
0 13147 5 1 1 13146
0 13148 7 1 2 13144 13147
0 13149 5 1 1 13148
0 13150 7 1 2 34452 13149
0 13151 5 1 1 13150
0 13152 7 1 2 26091 33949
0 13153 7 1 2 30613 13152
0 13154 7 1 2 30769 13153
0 13155 5 1 1 13154
0 13156 7 1 2 13151 13155
0 13157 5 1 1 13156
0 13158 7 1 2 26004 27178
0 13159 7 1 2 13157 13158
0 13160 5 1 1 13159
0 13161 7 1 2 13142 13160
0 13162 5 1 1 13161
0 13163 7 1 2 36493 13162
0 13164 5 1 1 13163
0 13165 7 1 2 22742 23202
0 13166 7 1 2 27637 13165
0 13167 7 2 2 33496 13166
0 13168 7 1 2 35412 36497
0 13169 5 1 1 13168
0 13170 7 3 2 33681 29807
0 13171 7 1 2 30486 34707
0 13172 7 1 2 36499 13171
0 13173 5 1 1 13172
0 13174 7 1 2 13169 13173
0 13175 5 1 1 13174
0 13176 7 1 2 29172 13175
0 13177 5 1 1 13176
0 13178 7 3 2 30052 34677
0 13179 7 3 2 29606 33964
0 13180 7 1 2 30030 36496
0 13181 7 1 2 36505 13180
0 13182 5 1 1 13181
0 13183 7 1 2 34281 29793
0 13184 7 1 2 30321 13183
0 13185 5 1 1 13184
0 13186 7 1 2 13182 13185
0 13187 5 1 1 13186
0 13188 7 1 2 36502 13187
0 13189 5 1 1 13188
0 13190 7 1 2 13177 13189
0 13191 5 1 1 13190
0 13192 7 1 2 27085 13191
0 13193 5 1 1 13192
0 13194 7 1 2 22479 35761
0 13195 5 1 1 13194
0 13196 7 2 2 27910 28924
0 13197 5 1 1 36508
0 13198 7 1 2 13195 13197
0 13199 5 1 1 13198
0 13200 7 4 2 24596 25130
0 13201 7 2 2 29540 36503
0 13202 7 1 2 36510 36514
0 13203 5 1 1 13202
0 13204 7 1 2 31039 33497
0 13205 7 1 2 35413 13204
0 13206 7 1 2 36375 13205
0 13207 5 1 1 13206
0 13208 7 1 2 13203 13207
0 13209 5 1 1 13208
0 13210 7 1 2 13199 13209
0 13211 5 1 1 13210
0 13212 7 1 2 27660 33287
0 13213 7 3 2 36369 33498
0 13214 7 1 2 35414 36516
0 13215 7 1 2 13212 13214
0 13216 5 1 1 13215
0 13217 7 1 2 25131 33093
0 13218 7 1 2 36515 13217
0 13219 5 1 1 13218
0 13220 7 1 2 13216 13219
0 13221 5 1 1 13220
0 13222 7 1 2 33213 13221
0 13223 5 1 1 13222
0 13224 7 1 2 13211 13223
0 13225 7 1 2 13193 13224
0 13226 7 1 2 13164 13225
0 13227 5 1 1 13226
0 13228 7 1 2 29002 13227
0 13229 5 1 1 13228
0 13230 7 1 2 35663 36498
0 13231 5 1 1 13230
0 13232 7 2 2 34661 36491
0 13233 5 1 1 36519
0 13234 7 2 2 22968 30086
0 13235 5 1 1 36521
0 13236 7 1 2 9774 13235
0 13237 5 4 1 13236
0 13238 7 1 2 32578 36523
0 13239 7 1 2 36520 13238
0 13240 5 1 1 13239
0 13241 7 1 2 13231 13240
0 13242 5 1 1 13241
0 13243 7 1 2 33100 13242
0 13244 5 1 1 13243
0 13245 7 1 2 34453 36494
0 13246 7 1 2 36524 13245
0 13247 5 1 1 13246
0 13248 7 1 2 23551 30710
0 13249 7 1 2 36376 13248
0 13250 7 1 2 29671 13249
0 13251 5 1 1 13250
0 13252 7 1 2 13247 13251
0 13253 5 1 1 13252
0 13254 7 1 2 30168 13253
0 13255 5 1 1 13254
0 13256 7 2 2 35664 36377
0 13257 7 1 2 33593 33503
0 13258 7 1 2 36527 13257
0 13259 5 1 1 13258
0 13260 7 1 2 13255 13259
0 13261 5 1 1 13260
0 13262 7 1 2 33846 13261
0 13263 5 1 1 13262
0 13264 7 1 2 13244 13263
0 13265 5 1 1 13264
0 13266 7 1 2 28826 13265
0 13267 5 1 1 13266
0 13268 7 1 2 12748 13233
0 13269 5 1 1 13268
0 13270 7 1 2 36522 13269
0 13271 5 1 1 13270
0 13272 7 1 2 27546 31231
0 13273 7 1 2 36500 13272
0 13274 5 1 1 13273
0 13275 7 1 2 13271 13274
0 13276 5 1 1 13275
0 13277 7 1 2 29173 13276
0 13278 5 1 1 13277
0 13279 7 2 2 26258 36525
0 13280 7 2 2 23203 36529
0 13281 7 1 2 34656 29406
0 13282 7 1 2 36531 13281
0 13283 5 1 1 13282
0 13284 7 1 2 13278 13283
0 13285 5 1 1 13284
0 13286 7 1 2 32804 13285
0 13287 5 1 1 13286
0 13288 7 1 2 29495 33623
0 13289 7 2 2 36530 13288
0 13290 7 1 2 32942 36533
0 13291 5 1 1 13290
0 13292 7 1 2 30696 32002
0 13293 7 1 2 33499 13292
0 13294 7 2 2 23127 34176
0 13295 7 1 2 35665 36535
0 13296 7 1 2 13293 13295
0 13297 5 1 1 13296
0 13298 7 1 2 13291 13297
0 13299 5 1 1 13298
0 13300 7 1 2 28156 13299
0 13301 5 1 1 13300
0 13302 7 1 2 13287 13301
0 13303 5 1 1 13302
0 13304 7 1 2 28733 13303
0 13305 5 1 1 13304
0 13306 7 1 2 36511 36504
0 13307 7 1 2 36526 13306
0 13308 5 1 1 13307
0 13309 7 1 2 36381 36517
0 13310 7 1 2 30712 13309
0 13311 5 1 1 13310
0 13312 7 1 2 13308 13311
0 13313 5 1 1 13312
0 13314 7 1 2 32579 13313
0 13315 5 1 1 13314
0 13316 7 1 2 32959 36534
0 13317 5 1 1 13316
0 13318 7 1 2 30114 30049
0 13319 7 1 2 36528 13318
0 13320 5 1 1 13319
0 13321 7 1 2 13317 13320
0 13322 7 1 2 13315 13321
0 13323 5 1 1 13322
0 13324 7 1 2 33049 13323
0 13325 5 1 1 13324
0 13326 7 2 2 31706 31859
0 13327 7 2 2 25076 25441
0 13328 7 1 2 24977 31103
0 13329 7 1 2 36539 13328
0 13330 7 1 2 36537 13329
0 13331 7 1 2 32964 13330
0 13332 7 1 2 36532 13331
0 13333 5 1 1 13332
0 13334 7 1 2 13325 13333
0 13335 7 1 2 13305 13334
0 13336 7 1 2 13267 13335
0 13337 7 1 2 13229 13336
0 13338 5 1 1 13337
0 13339 7 1 2 26167 13338
0 13340 5 1 1 13339
0 13341 7 6 2 23707 23939
0 13342 7 2 2 26470 36541
0 13343 7 2 2 23047 36370
0 13344 7 3 2 22629 36549
0 13345 7 1 2 36547 36551
0 13346 5 1 1 13345
0 13347 7 1 2 29058 33682
0 13348 7 1 2 34839 13347
0 13349 5 1 1 13348
0 13350 7 1 2 13346 13349
0 13351 5 1 1 13350
0 13352 7 1 2 24777 13351
0 13353 5 1 1 13352
0 13354 7 1 2 31663 30255
0 13355 7 2 2 22846 25500
0 13356 7 1 2 33683 36554
0 13357 7 1 2 13354 13356
0 13358 5 1 1 13357
0 13359 7 1 2 13353 13358
0 13360 5 1 1 13359
0 13361 7 1 2 26168 13360
0 13362 5 1 1 13361
0 13363 7 1 2 35077 34925
0 13364 5 2 1 13363
0 13365 7 3 2 36542 36556
0 13366 7 1 2 36558 36552
0 13367 5 1 1 13366
0 13368 7 1 2 13362 13367
0 13369 5 1 1 13368
0 13370 7 1 2 26259 13369
0 13371 5 1 1 13370
0 13372 7 1 2 24288 28524
0 13373 7 3 2 8060 13372
0 13374 7 3 2 36543 36561
0 13375 7 3 2 36371 34849
0 13376 7 1 2 22630 36567
0 13377 7 1 2 36564 13376
0 13378 5 1 1 13377
0 13379 7 1 2 13371 13378
0 13380 5 1 1 13379
0 13381 7 1 2 33325 13380
0 13382 5 1 1 13381
0 13383 7 1 2 22847 26460
0 13384 5 1 1 13383
0 13385 7 1 2 34926 13384
0 13386 5 10 1 13385
0 13387 7 3 2 32987 36570
0 13388 7 1 2 27414 30450
0 13389 7 1 2 34252 13388
0 13390 7 1 2 34599 13389
0 13391 7 1 2 36580 13390
0 13392 5 1 1 13391
0 13393 7 1 2 13382 13392
0 13394 5 1 1 13393
0 13395 7 1 2 34983 13394
0 13396 5 1 1 13395
0 13397 7 3 2 25709 27975
0 13398 5 1 1 36583
0 13399 7 1 2 34692 36571
0 13400 7 2 2 36584 13399
0 13401 7 1 2 31945 36586
0 13402 5 1 1 13401
0 13403 7 2 2 35002 36372
0 13404 7 1 2 33288 36548
0 13405 7 1 2 36588 13404
0 13406 5 1 1 13405
0 13407 7 1 2 13402 13406
0 13408 5 1 1 13407
0 13409 7 1 2 26169 13408
0 13410 5 1 1 13409
0 13411 7 1 2 33289 36550
0 13412 7 1 2 36559 13411
0 13413 5 1 1 13412
0 13414 7 1 2 13410 13413
0 13415 5 1 1 13414
0 13416 7 1 2 34984 13415
0 13417 5 1 1 13416
0 13418 7 1 2 35385 29496
0 13419 7 1 2 31447 13418
0 13420 7 1 2 34454 13419
0 13421 7 1 2 36572 13420
0 13422 5 1 1 13421
0 13423 7 2 2 23479 30201
0 13424 7 5 2 28553 33660
0 13425 7 1 2 26471 35936
0 13426 7 1 2 36592 13425
0 13427 7 1 2 36590 13426
0 13428 5 1 1 13427
0 13429 7 1 2 13422 13428
0 13430 5 1 1 13429
0 13431 7 1 2 26170 13430
0 13432 5 1 1 13431
0 13433 7 1 2 24030 30743
0 13434 7 2 2 36557 13433
0 13435 7 1 2 36553 36597
0 13436 7 1 2 36591 13435
0 13437 5 1 1 13436
0 13438 7 1 2 13432 13437
0 13439 7 1 2 13417 13438
0 13440 5 1 1 13439
0 13441 7 1 2 26260 13440
0 13442 5 1 1 13441
0 13443 7 3 2 24978 25912
0 13444 5 1 1 36599
0 13445 7 1 2 31562 34373
0 13446 7 1 2 36600 13445
0 13447 7 1 2 31043 33752
0 13448 7 2 2 13446 13447
0 13449 7 1 2 33094 36602
0 13450 5 1 1 13449
0 13451 7 1 2 33290 36568
0 13452 7 1 2 34985 13451
0 13453 7 1 2 36565 13452
0 13454 5 1 1 13453
0 13455 7 1 2 13450 13454
0 13456 7 1 2 13442 13455
0 13457 5 1 1 13456
0 13458 7 1 2 32247 13457
0 13459 5 1 1 13458
0 13460 7 1 2 33337 31448
0 13461 7 1 2 33688 13460
0 13462 7 1 2 36573 13461
0 13463 5 1 1 13462
0 13464 7 1 2 26472 32478
0 13465 7 3 2 23204 31540
0 13466 7 2 2 26952 30441
0 13467 7 1 2 36604 36607
0 13468 7 1 2 13464 13467
0 13469 5 1 1 13468
0 13470 7 1 2 13463 13469
0 13471 5 1 1 13470
0 13472 7 1 2 26171 13471
0 13473 5 1 1 13472
0 13474 7 1 2 35653 30442
0 13475 7 1 2 34374 13474
0 13476 7 1 2 36598 13475
0 13477 5 1 1 13476
0 13478 7 1 2 13473 13477
0 13479 5 1 1 13478
0 13480 7 1 2 26261 13479
0 13481 5 1 1 13480
0 13482 7 1 2 24597 36603
0 13483 5 1 1 13482
0 13484 7 1 2 13481 13483
0 13485 5 1 1 13484
0 13486 7 1 2 33326 13485
0 13487 5 1 1 13486
0 13488 7 1 2 35281 31973
0 13489 7 2 2 33965 31713
0 13490 7 1 2 31449 36609
0 13491 7 1 2 13488 13490
0 13492 7 1 2 36581 13491
0 13493 5 1 1 13492
0 13494 7 1 2 13487 13493
0 13495 7 1 2 13459 13494
0 13496 7 1 2 13396 13495
0 13497 7 1 2 27624 36593
0 13498 5 1 1 13497
0 13499 7 1 2 26172 29497
0 13500 7 1 2 34489 13499
0 13501 5 1 1 13500
0 13502 7 1 2 13498 13501
0 13503 5 1 1 13502
0 13504 7 1 2 22969 13503
0 13505 5 1 1 13504
0 13506 7 1 2 28513 36594
0 13507 5 1 1 13506
0 13508 7 1 2 13505 13507
0 13509 5 1 1 13508
0 13510 7 1 2 24778 13509
0 13511 5 1 1 13510
0 13512 7 1 2 24195 36595
0 13513 5 1 1 13512
0 13514 7 1 2 29326 36202
0 13515 5 1 1 13514
0 13516 7 1 2 13513 13515
0 13517 5 1 1 13516
0 13518 7 1 2 36555 13517
0 13519 5 1 1 13518
0 13520 7 1 2 13511 13519
0 13521 5 1 1 13520
0 13522 7 1 2 26262 13521
0 13523 5 1 1 13522
0 13524 7 1 2 23708 36569
0 13525 7 1 2 36562 13524
0 13526 5 1 1 13525
0 13527 7 1 2 13523 13526
0 13528 5 1 1 13527
0 13529 7 1 2 29174 13528
0 13530 5 1 1 13529
0 13531 7 1 2 30577 34235
0 13532 7 2 2 34606 13531
0 13533 7 1 2 36582 36611
0 13534 5 1 1 13533
0 13535 7 1 2 13530 13534
0 13536 5 1 1 13535
0 13537 7 1 2 33805 13536
0 13538 5 1 1 13537
0 13539 7 1 2 35842 36587
0 13540 5 1 1 13539
0 13541 7 2 2 35193 33661
0 13542 7 1 2 27647 35845
0 13543 7 1 2 26473 13542
0 13544 7 1 2 36613 13543
0 13545 5 1 1 13544
0 13546 7 1 2 13540 13545
0 13547 5 1 1 13546
0 13548 7 1 2 26173 13547
0 13549 5 1 1 13548
0 13550 7 1 2 27786 36266
0 13551 7 1 2 35847 13550
0 13552 7 1 2 36560 13551
0 13553 5 1 1 13552
0 13554 7 1 2 13549 13553
0 13555 5 1 1 13554
0 13556 7 1 2 26263 13555
0 13557 5 1 1 13556
0 13558 7 1 2 28590 35607
0 13559 7 1 2 36563 13558
0 13560 7 1 2 36614 13559
0 13561 5 1 1 13560
0 13562 7 1 2 13557 13561
0 13563 5 1 1 13562
0 13564 7 1 2 28157 13563
0 13565 5 1 1 13564
0 13566 7 2 2 27648 33761
0 13567 7 1 2 23709 32707
0 13568 7 1 2 33007 13567
0 13569 7 1 2 36615 13568
0 13570 7 1 2 29195 13569
0 13571 5 1 1 13570
0 13572 7 1 2 13565 13571
0 13573 7 1 2 13538 13572
0 13574 5 1 1 13573
0 13575 7 1 2 32108 13574
0 13576 5 1 1 13575
0 13577 7 1 2 24689 23710
0 13578 7 2 2 36589 13577
0 13579 7 1 2 27616 30783
0 13580 7 1 2 36617 13579
0 13581 5 1 1 13580
0 13582 7 2 2 34951 34718
0 13583 7 3 2 26174 34678
0 13584 7 1 2 33586 36621
0 13585 7 1 2 36619 13584
0 13586 5 1 1 13585
0 13587 7 1 2 13581 13586
0 13588 5 1 1 13587
0 13589 7 1 2 22480 13588
0 13590 5 1 1 13589
0 13591 7 1 2 34490 36622
0 13592 7 2 2 22848 30582
0 13593 7 3 2 24463 22743
0 13594 7 2 2 23271 36626
0 13595 7 1 2 36624 36629
0 13596 7 1 2 13591 13595
0 13597 5 1 1 13596
0 13598 7 1 2 13590 13597
0 13599 5 1 1 13598
0 13600 7 1 2 26917 13599
0 13601 5 1 1 13600
0 13602 7 2 2 22970 36226
0 13603 7 1 2 30836 33684
0 13604 7 1 2 33589 13603
0 13605 7 1 2 36631 13604
0 13606 5 1 1 13605
0 13607 7 1 2 25379 26397
0 13608 7 1 2 33084 13607
0 13609 7 3 2 23711 35129
0 13610 7 1 2 36536 36633
0 13611 7 1 2 13608 13610
0 13612 5 1 1 13611
0 13613 7 1 2 13606 13612
0 13614 5 1 1 13613
0 13615 7 1 2 22481 13614
0 13616 5 1 1 13615
0 13617 7 1 2 27179 30619
0 13618 5 1 1 13617
0 13619 7 2 2 30685 34621
0 13620 5 1 1 36636
0 13621 7 1 2 13618 13620
0 13622 5 1 1 13621
0 13623 7 1 2 22482 13622
0 13624 5 1 1 13623
0 13625 7 1 2 30982 35835
0 13626 5 1 1 13625
0 13627 7 1 2 13624 13626
0 13628 5 1 1 13627
0 13629 7 2 2 29861 36596
0 13630 7 1 2 34155 36638
0 13631 5 1 1 13630
0 13632 7 1 2 30099 26850
0 13633 7 1 2 36501 13632
0 13634 5 1 1 13633
0 13635 7 1 2 13631 13634
0 13636 5 1 1 13635
0 13637 7 1 2 13628 13636
0 13638 5 1 1 13637
0 13639 7 4 2 34952 28605
0 13640 7 2 2 23272 36640
0 13641 7 1 2 34733 36644
0 13642 5 1 1 13641
0 13643 7 1 2 30210 31374
0 13644 7 1 2 36483 13643
0 13645 5 1 1 13644
0 13646 7 1 2 13642 13645
0 13647 5 1 1 13646
0 13648 7 1 2 33168 34607
0 13649 7 1 2 13647 13648
0 13650 5 1 1 13649
0 13651 7 1 2 13638 13650
0 13652 7 1 2 13616 13651
0 13653 7 1 2 13601 13652
0 13654 5 1 1 13653
0 13655 7 1 2 26264 13654
0 13656 5 1 1 13655
0 13657 7 1 2 24779 23205
0 13658 7 1 2 30015 13657
0 13659 7 1 2 34027 13658
0 13660 7 1 2 36566 13659
0 13661 5 1 1 13660
0 13662 7 1 2 13656 13661
0 13663 5 1 1 13662
0 13664 7 1 2 28158 13663
0 13665 5 1 1 13664
0 13666 7 1 2 35130 32289
0 13667 5 1 1 13666
0 13668 7 1 2 33358 33002
0 13669 5 1 1 13668
0 13670 7 1 2 13667 13669
0 13671 5 1 1 13670
0 13672 7 1 2 26474 13671
0 13673 5 1 1 13672
0 13674 7 2 2 29059 33359
0 13675 5 2 1 36646
0 13676 7 1 2 22744 35049
0 13677 5 1 1 13676
0 13678 7 1 2 36648 13677
0 13679 5 1 1 13678
0 13680 7 1 2 26747 13679
0 13681 5 1 1 13680
0 13682 7 1 2 13673 13681
0 13683 5 1 1 13682
0 13684 7 1 2 36605 13683
0 13685 5 1 1 13684
0 13686 7 2 2 29525 36216
0 13687 5 1 1 36650
0 13688 7 1 2 36649 13687
0 13689 5 2 1 13688
0 13690 7 2 2 25132 29327
0 13691 7 1 2 36492 36654
0 13692 7 1 2 36652 13691
0 13693 5 1 1 13692
0 13694 7 1 2 13685 13693
0 13695 5 1 1 13694
0 13696 7 1 2 26999 13695
0 13697 5 1 1 13696
0 13698 7 1 2 23940 27270
0 13699 7 1 2 36639 13698
0 13700 5 1 1 13699
0 13701 7 2 2 30031 36217
0 13702 7 1 2 34679 36655
0 13703 7 1 2 36656 13702
0 13704 5 1 1 13703
0 13705 7 1 2 13700 13704
0 13706 5 1 1 13705
0 13707 7 1 2 27086 13706
0 13708 5 1 1 13707
0 13709 7 1 2 25710 34960
0 13710 7 1 2 36001 13709
0 13711 7 1 2 36620 13710
0 13712 5 1 1 13711
0 13713 7 2 2 23418 25501
0 13714 5 1 1 36658
0 13715 7 1 2 28930 36659
0 13716 7 1 2 36618 13715
0 13717 5 1 1 13716
0 13718 7 1 2 13712 13717
0 13719 7 1 2 13708 13718
0 13720 5 1 1 13719
0 13721 7 1 2 26265 13720
0 13722 5 1 1 13721
0 13723 7 1 2 36002 30003
0 13724 5 1 1 13723
0 13725 7 1 2 24196 26475
0 13726 7 1 2 32789 13725
0 13727 5 1 1 13726
0 13728 7 1 2 13724 13727
0 13729 5 1 1 13728
0 13730 7 1 2 24289 30843
0 13731 7 1 2 36616 13730
0 13732 7 1 2 13729 13731
0 13733 5 1 1 13732
0 13734 7 1 2 13722 13733
0 13735 7 1 2 13697 13734
0 13736 5 1 1 13735
0 13737 7 1 2 29175 13736
0 13738 5 1 1 13737
0 13739 7 1 2 27000 36653
0 13740 5 1 1 13739
0 13741 7 1 2 26928 36657
0 13742 5 1 1 13741
0 13743 7 1 2 32796 34964
0 13744 5 1 1 13743
0 13745 7 1 2 13742 13744
0 13746 7 1 2 13740 13745
0 13747 5 1 1 13746
0 13748 7 1 2 32988 36612
0 13749 7 1 2 13747 13748
0 13750 5 1 1 13749
0 13751 7 1 2 13738 13750
0 13752 7 1 2 13665 13751
0 13753 5 1 1 13752
0 13754 7 1 2 34939 13753
0 13755 5 1 1 13754
0 13756 7 1 2 13576 13755
0 13757 7 1 2 13496 13756
0 13758 5 1 1 13757
0 13759 7 1 2 25577 13758
0 13760 5 1 1 13759
0 13761 7 1 2 13340 13760
0 13762 5 1 1 13761
0 13763 7 1 2 25811 13762
0 13764 5 1 1 13763
0 13765 7 3 2 26092 29003
0 13766 7 1 2 30942 33242
0 13767 5 1 1 13766
0 13768 7 1 2 25913 35782
0 13769 5 1 1 13768
0 13770 7 1 2 13767 13769
0 13771 5 2 1 13770
0 13772 7 1 2 36660 36663
0 13773 5 1 1 13772
0 13774 7 1 2 32600 28840
0 13775 5 1 1 13774
0 13776 7 1 2 28734 33131
0 13777 5 1 1 13776
0 13778 7 1 2 35863 32960
0 13779 5 1 1 13778
0 13780 7 1 2 13777 13779
0 13781 7 1 2 13775 13780
0 13782 5 1 1 13781
0 13783 7 1 2 24108 13782
0 13784 5 1 1 13783
0 13785 7 1 2 13773 13784
0 13786 5 1 1 13785
0 13787 7 1 2 35201 33481
0 13788 5 1 1 13787
0 13789 7 1 2 28514 26566
0 13790 5 1 1 13789
0 13791 7 1 2 13788 13790
0 13792 5 1 1 13791
0 13793 7 1 2 13786 13792
0 13794 5 1 1 13793
0 13795 7 1 2 33935 33231
0 13796 5 2 1 13795
0 13797 7 1 2 33190 33243
0 13798 5 1 1 13797
0 13799 7 2 2 26953 32900
0 13800 5 1 1 36667
0 13801 7 1 2 13798 13800
0 13802 5 1 1 13801
0 13803 7 1 2 33899 13802
0 13804 5 1 1 13803
0 13805 7 1 2 36665 13804
0 13806 5 1 1 13805
0 13807 7 1 2 26476 32290
0 13808 7 1 2 13806 13807
0 13809 5 1 1 13808
0 13810 7 1 2 33900 36664
0 13811 5 1 1 13810
0 13812 7 1 2 36666 13811
0 13813 5 1 1 13812
0 13814 7 1 2 25502 33079
0 13815 7 1 2 13813 13814
0 13816 5 1 1 13815
0 13817 7 1 2 13809 13816
0 13818 5 1 1 13817
0 13819 7 1 2 25578 13818
0 13820 5 1 1 13819
0 13821 7 1 2 13794 13820
0 13822 5 1 1 13821
0 13823 7 1 2 23128 13822
0 13824 5 1 1 13823
0 13825 7 1 2 29283 30925
0 13826 5 1 1 13825
0 13827 7 1 2 26761 29343
0 13828 5 1 1 13827
0 13829 7 1 2 24109 29322
0 13830 7 1 2 13828 13829
0 13831 5 1 1 13830
0 13832 7 1 2 13826 13831
0 13833 5 1 1 13832
0 13834 7 1 2 25579 13833
0 13835 5 1 1 13834
0 13836 7 1 2 24290 27514
0 13837 5 1 1 13836
0 13838 7 1 2 13835 13837
0 13839 5 1 1 13838
0 13840 7 1 2 23552 13839
0 13841 5 1 1 13840
0 13842 7 5 2 24110 32989
0 13843 7 1 2 22971 36275
0 13844 7 1 2 36669 13843
0 13845 5 1 1 13844
0 13846 7 1 2 13841 13845
0 13847 5 1 1 13846
0 13848 7 1 2 35932 32014
0 13849 7 1 2 13847 13848
0 13850 5 1 1 13849
0 13851 7 1 2 13824 13850
0 13852 5 1 1 13851
0 13853 7 1 2 33225 33662
0 13854 7 1 2 13852 13853
0 13855 5 1 1 13854
0 13856 7 1 2 13764 13855
0 13857 5 1 1 13856
0 13858 7 1 2 22371 13857
0 13859 5 1 1 13858
0 13860 7 1 2 34920 32945
0 13861 5 1 1 13860
0 13862 7 1 2 22483 35342
0 13863 5 1 1 13862
0 13864 7 3 2 24464 28363
0 13865 7 1 2 35337 36674
0 13866 5 1 1 13865
0 13867 7 1 2 13863 13866
0 13868 5 1 1 13867
0 13869 7 1 2 32965 13868
0 13870 5 1 1 13869
0 13871 7 1 2 35320 32953
0 13872 5 1 1 13871
0 13873 7 1 2 13870 13872
0 13874 7 1 2 13861 13873
0 13875 5 1 1 13874
0 13876 7 1 2 36574 13875
0 13877 5 1 1 13876
0 13878 7 1 2 7738 13714
0 13879 5 1 1 13878
0 13880 7 1 2 10385 26544
0 13881 7 3 2 13879 13880
0 13882 7 1 2 32946 36677
0 13883 5 1 1 13882
0 13884 7 2 2 27389 33587
0 13885 7 1 2 34953 36680
0 13886 5 1 1 13885
0 13887 7 1 2 35195 32154
0 13888 5 1 1 13887
0 13889 7 1 2 13886 13888
0 13890 5 2 1 13889
0 13891 7 1 2 22484 36682
0 13892 5 1 1 13891
0 13893 7 1 2 36641 36675
0 13894 5 1 1 13893
0 13895 7 1 2 13892 13894
0 13896 5 1 1 13895
0 13897 7 1 2 32966 13896
0 13898 5 1 1 13897
0 13899 7 1 2 26461 35323
0 13900 5 1 1 13899
0 13901 7 2 2 23419 29060
0 13902 7 1 2 35814 36684
0 13903 5 1 1 13902
0 13904 7 1 2 13900 13903
0 13905 5 4 1 13904
0 13906 7 1 2 32954 36686
0 13907 5 1 1 13906
0 13908 7 1 2 13898 13907
0 13909 7 1 2 13883 13908
0 13910 5 1 1 13909
0 13911 7 1 2 34940 13910
0 13912 5 1 1 13911
0 13913 7 1 2 13877 13912
0 13914 5 1 1 13913
0 13915 7 4 2 26175 34089
0 13916 7 1 2 33730 36690
0 13917 7 1 2 13914 13916
0 13918 5 1 1 13917
0 13919 7 1 2 13859 13918
0 13920 7 1 2 13131 13919
0 13921 5 1 1 13920
0 13922 7 1 2 27482 13921
0 13923 5 1 1 13922
0 13924 7 1 2 12975 13923
0 13925 7 1 2 12973 13924
0 13926 7 1 2 11108 13925
0 13927 7 1 2 7660 13926
0 13928 7 1 2 5598 13927
0 13929 5 1 1 13928
0 13930 7 1 2 23646 13929
0 13931 5 1 1 13930
0 13932 7 10 2 23571 26644
0 13933 7 1 2 32522 36694
0 13934 5 1 1 13933
0 13935 7 2 2 26093 28416
0 13936 7 4 2 25580 23636
0 13937 7 1 2 24780 36706
0 13938 7 1 2 36704 13937
0 13939 5 1 1 13938
0 13940 7 1 2 13934 13939
0 13941 5 1 1 13940
0 13942 7 1 2 23048 13941
0 13943 5 1 1 13942
0 13944 7 2 2 24781 28417
0 13945 7 5 2 23572 23637
0 13946 7 1 2 30926 36712
0 13947 7 1 2 36710 13946
0 13948 5 1 1 13947
0 13949 7 1 2 13943 13948
0 13950 5 1 1 13949
0 13951 7 1 2 23129 13950
0 13952 5 1 1 13951
0 13953 7 1 2 35104 33257
0 13954 5 1 1 13953
0 13955 7 1 2 13952 13954
0 13956 5 1 1 13955
0 13957 7 1 2 26777 13956
0 13958 5 1 1 13957
0 13959 7 9 2 28554 36695
0 13960 5 1 1 36717
0 13961 7 2 2 32548 36718
0 13962 5 1 1 36726
0 13963 7 2 2 24031 36727
0 13964 7 1 2 23420 36728
0 13965 5 1 1 13964
0 13966 7 1 2 13958 13965
0 13967 5 1 1 13966
0 13968 7 1 2 32612 13967
0 13969 5 1 1 13968
0 13970 7 3 2 23573 34856
0 13971 7 1 2 35612 35003
0 13972 7 1 2 29803 13971
0 13973 7 1 2 36730 13972
0 13974 5 1 1 13973
0 13975 7 1 2 13969 13974
0 13976 5 1 1 13975
0 13977 7 1 2 24906 13976
0 13978 5 1 1 13977
0 13979 7 2 2 32634 26864
0 13980 7 1 2 36733 36729
0 13981 5 1 1 13980
0 13982 7 1 2 13978 13981
0 13983 5 1 1 13982
0 13984 7 1 2 24690 13983
0 13985 5 1 1 13984
0 13986 7 2 2 24032 36696
0 13987 7 1 2 35289 30184
0 13988 7 1 2 32549 13987
0 13989 7 1 2 32624 13988
0 13990 7 1 2 36735 13989
0 13991 5 1 1 13990
0 13992 7 1 2 13985 13991
0 13993 5 1 1 13992
0 13994 7 1 2 22631 13993
0 13995 5 1 1 13994
0 13996 7 1 2 26266 29715
0 13997 5 2 1 13996
0 13998 7 1 2 26722 36737
0 13999 5 2 1 13998
0 14000 7 1 2 28854 36739
0 14001 5 2 1 14000
0 14002 7 13 2 23130 35209
0 14003 5 1 1 36743
0 14004 7 1 2 30169 36744
0 14005 5 1 1 14004
0 14006 7 1 2 36741 14005
0 14007 5 1 1 14006
0 14008 7 1 2 35028 14007
0 14009 5 1 1 14008
0 14010 7 1 2 35085 28690
0 14011 7 1 2 30722 14010
0 14012 5 1 1 14011
0 14013 7 1 2 14009 14012
0 14014 5 1 1 14013
0 14015 7 1 2 26094 14014
0 14016 5 1 1 14015
0 14017 7 1 2 30170 28418
0 14018 5 1 1 14017
0 14019 7 1 2 36742 14018
0 14020 5 1 1 14019
0 14021 7 1 2 22849 31219
0 14022 7 1 2 14020 14021
0 14023 5 1 1 14022
0 14024 7 1 2 14016 14023
0 14025 5 1 1 14024
0 14026 7 1 2 30443 36731
0 14027 7 1 2 14025 14026
0 14028 5 1 1 14027
0 14029 7 1 2 24197 14028
0 14030 7 1 2 13995 14029
0 14031 5 1 1 14030
0 14032 7 2 2 24291 26515
0 14033 5 1 1 36756
0 14034 7 1 2 26678 14033
0 14035 5 8 1 14034
0 14036 7 2 2 32550 36758
0 14037 7 2 2 23574 24033
0 14038 7 3 2 22632 24979
0 14039 7 1 2 32613 36770
0 14040 7 1 2 36768 14039
0 14041 5 1 1 14040
0 14042 7 3 2 22633 24034
0 14043 5 1 1 36773
0 14044 7 1 2 32614 36276
0 14045 7 1 2 36774 14044
0 14046 5 1 1 14045
0 14047 7 1 2 14041 14046
0 14048 5 1 1 14047
0 14049 7 1 2 36766 14048
0 14050 5 1 1 14049
0 14051 7 1 2 26267 32523
0 14052 5 1 1 14051
0 14053 7 1 2 26268 26609
0 14054 5 1 1 14053
0 14055 7 1 2 14003 14054
0 14056 5 20 1 14055
0 14057 7 1 2 32512 36776
0 14058 5 1 1 14057
0 14059 7 1 2 14052 14058
0 14060 5 1 1 14059
0 14061 7 4 2 32635 34061
0 14062 7 1 2 27396 36796
0 14063 7 1 2 14060 14062
0 14064 5 1 1 14063
0 14065 7 1 2 14050 14064
0 14066 5 1 1 14065
0 14067 7 1 2 23421 14066
0 14068 5 1 1 14067
0 14069 7 27 2 34079 33566
0 14070 5 1 1 36800
0 14071 7 1 2 32524 26659
0 14072 5 1 1 14071
0 14073 7 1 2 35659 30568
0 14074 7 1 2 36738 14073
0 14075 5 1 1 14074
0 14076 7 1 2 14072 14075
0 14077 5 1 1 14076
0 14078 7 1 2 36801 14077
0 14079 5 1 1 14078
0 14080 7 3 2 35457 28895
0 14081 5 1 1 36827
0 14082 7 1 2 32017 34090
0 14083 5 1 1 14082
0 14084 7 1 2 14081 14083
0 14085 5 2 1 14084
0 14086 7 1 2 32525 36830
0 14087 5 1 1 14086
0 14088 7 1 2 14079 14087
0 14089 5 1 1 14088
0 14090 7 1 2 22634 32151
0 14091 7 1 2 35014 14090
0 14092 7 1 2 14089 14091
0 14093 5 1 1 14092
0 14094 7 1 2 14068 14093
0 14095 5 1 1 14094
0 14096 7 1 2 24907 14095
0 14097 5 1 1 14096
0 14098 7 2 2 22972 36767
0 14099 7 1 2 22635 33861
0 14100 7 1 2 34961 14099
0 14101 7 1 2 36802 14100
0 14102 7 1 2 36832 14101
0 14103 5 1 1 14102
0 14104 7 1 2 14097 14103
0 14105 5 1 1 14104
0 14106 7 1 2 24691 14105
0 14107 5 1 1 14106
0 14108 7 5 2 28855 32551
0 14109 5 2 1 36834
0 14110 7 1 2 22636 28791
0 14111 7 3 2 26462 14110
0 14112 5 1 1 36841
0 14113 7 3 2 27365 32646
0 14114 5 1 1 36844
0 14115 7 1 2 14112 14114
0 14116 5 1 1 14115
0 14117 7 1 2 26681 14116
0 14118 5 1 1 14117
0 14119 7 2 2 28807 29061
0 14120 7 1 2 24598 35645
0 14121 7 1 2 36847 14120
0 14122 5 1 1 14121
0 14123 7 1 2 14118 14122
0 14124 5 1 1 14123
0 14125 7 1 2 36803 14124
0 14126 5 1 1 14125
0 14127 7 10 2 26269 26516
0 14128 5 1 1 36849
0 14129 7 1 2 24599 30953
0 14130 7 1 2 36850 14129
0 14131 7 1 2 36797 14130
0 14132 5 1 1 14131
0 14133 7 1 2 14126 14132
0 14134 5 1 1 14133
0 14135 7 1 2 36835 14134
0 14136 5 1 1 14135
0 14137 7 1 2 26176 14136
0 14138 7 1 2 14107 14137
0 14139 5 1 1 14138
0 14140 7 1 2 14031 14139
0 14141 5 1 1 14140
0 14142 7 2 2 34869 30247
0 14143 5 1 1 36859
0 14144 7 1 2 36860 36845
0 14145 5 1 1 14144
0 14146 7 1 2 29193 36804
0 14147 7 1 2 36842 14146
0 14148 5 1 1 14147
0 14149 7 1 2 14145 14148
0 14150 5 1 1 14149
0 14151 7 1 2 23638 14150
0 14152 5 1 1 14151
0 14153 7 1 2 23575 32031
0 14154 7 1 2 29631 14153
0 14155 7 1 2 36846 14154
0 14156 5 1 1 14155
0 14157 7 1 2 14152 14156
0 14158 5 1 1 14157
0 14159 7 1 2 30171 463
0 14160 7 1 2 33143 14159
0 14161 5 1 1 14160
0 14162 7 1 2 36839 14161
0 14163 5 1 1 14162
0 14164 7 1 2 14158 14163
0 14165 5 1 1 14164
0 14166 7 1 2 22745 33057
0 14167 5 1 1 14166
0 14168 7 1 2 27661 32647
0 14169 5 1 1 14168
0 14170 7 1 2 14167 14169
0 14171 5 4 1 14170
0 14172 7 2 2 35243 36486
0 14173 5 1 1 36865
0 14174 7 4 2 23576 24198
0 14175 5 2 1 36867
0 14176 7 1 2 28555 36868
0 14177 5 1 1 14176
0 14178 7 1 2 14173 14177
0 14179 5 1 1 14178
0 14180 7 1 2 32526 14179
0 14181 5 1 1 14180
0 14182 7 3 2 26496 29328
0 14183 5 1 1 36873
0 14184 7 2 2 26415 28466
0 14185 5 1 1 36876
0 14186 7 1 2 14183 14185
0 14187 5 3 1 14186
0 14188 7 1 2 32513 36805
0 14189 7 1 2 36878 14188
0 14190 5 1 1 14189
0 14191 7 1 2 14181 14190
0 14192 5 1 1 14191
0 14193 7 1 2 26270 14192
0 14194 5 1 1 14193
0 14195 7 1 2 32527 34062
0 14196 7 1 2 36877 14195
0 14197 5 1 1 14196
0 14198 7 1 2 14194 14197
0 14199 5 1 1 14198
0 14200 7 1 2 27397 14199
0 14201 5 1 1 14200
0 14202 7 3 2 26095 27398
0 14203 7 3 2 26177 26624
0 14204 7 1 2 35004 36884
0 14205 5 1 1 14204
0 14206 7 1 2 34852 31073
0 14207 5 1 1 14206
0 14208 7 1 2 14205 14207
0 14209 5 1 1 14208
0 14210 7 1 2 36881 14209
0 14211 5 1 1 14210
0 14212 7 2 2 24199 26436
0 14213 7 1 2 31425 30483
0 14214 7 1 2 36887 14213
0 14215 5 1 1 14214
0 14216 7 1 2 26723 28534
0 14217 5 1 1 14216
0 14218 7 1 2 28833 33161
0 14219 7 1 2 14217 14218
0 14220 5 1 1 14219
0 14221 7 1 2 14215 14220
0 14222 5 1 1 14221
0 14223 7 1 2 24111 14222
0 14224 5 1 1 14223
0 14225 7 1 2 25581 14224
0 14226 7 1 2 14211 14225
0 14227 5 1 1 14226
0 14228 7 1 2 32514 26625
0 14229 5 2 1 14228
0 14230 7 1 2 26517 32528
0 14231 5 1 1 14230
0 14232 7 1 2 36889 14231
0 14233 5 2 1 14232
0 14234 7 8 2 24600 24980
0 14235 5 1 1 36893
0 14236 7 1 2 33162 36894
0 14237 7 1 2 36891 14236
0 14238 5 1 1 14237
0 14239 7 1 2 23577 14238
0 14240 5 1 1 14239
0 14241 7 1 2 24292 14240
0 14242 7 1 2 14227 14241
0 14243 5 1 1 14242
0 14244 7 1 2 14201 14243
0 14245 5 1 1 14244
0 14246 7 1 2 36861 14245
0 14247 5 1 1 14246
0 14248 7 1 2 14165 14247
0 14249 7 1 2 14141 14248
0 14250 5 1 1 14249
0 14251 7 1 2 23354 14250
0 14252 5 1 1 14251
0 14253 7 2 2 26005 36862
0 14254 7 1 2 24293 36892
0 14255 5 1 1 14254
0 14256 7 1 2 33089 29129
0 14257 5 1 1 14256
0 14258 7 1 2 14255 14257
0 14259 5 1 1 14258
0 14260 7 1 2 26178 14259
0 14261 5 1 1 14260
0 14262 7 6 2 23639 26096
0 14263 5 1 1 36903
0 14264 7 1 2 28467 36904
0 14265 7 1 2 36711 14264
0 14266 5 1 1 14265
0 14267 7 1 2 14261 14266
0 14268 5 1 1 14267
0 14269 7 1 2 36901 14268
0 14270 5 1 1 14269
0 14271 7 1 2 30983 35990
0 14272 7 1 2 36833 14271
0 14273 5 1 1 14272
0 14274 7 1 2 14270 14273
0 14275 5 1 1 14274
0 14276 7 1 2 36806 14275
0 14277 5 1 1 14276
0 14278 7 2 2 27509 35203
0 14279 5 1 1 36909
0 14280 7 6 2 24200 29616
0 14281 7 1 2 35688 36911
0 14282 5 1 1 14281
0 14283 7 1 2 14279 14282
0 14284 5 1 1 14283
0 14285 7 1 2 24981 14284
0 14286 5 1 1 14285
0 14287 7 1 2 25582 25635
0 14288 7 1 2 36670 14287
0 14289 5 1 1 14288
0 14290 7 1 2 14286 14289
0 14291 5 1 1 14290
0 14292 7 2 2 25077 14291
0 14293 5 1 1 36917
0 14294 7 2 2 22850 36902
0 14295 7 1 2 36918 36919
0 14296 5 1 1 14295
0 14297 7 1 2 27510 26660
0 14298 7 2 2 36707 14297
0 14299 7 1 2 36920 36921
0 14300 5 1 1 14299
0 14301 7 3 2 29834 33360
0 14302 5 1 1 36923
0 14303 7 1 2 36924 36848
0 14304 5 2 1 14303
0 14305 7 2 2 23422 36453
0 14306 5 1 1 36928
0 14307 7 1 2 32529 36929
0 14308 5 1 1 14307
0 14309 7 1 2 27087 8696
0 14310 7 1 2 32552 35516
0 14311 7 1 2 14309 14310
0 14312 5 1 1 14311
0 14313 7 1 2 14308 14312
0 14314 5 1 1 14313
0 14315 7 1 2 22746 14314
0 14316 5 1 1 14315
0 14317 7 1 2 36926 14316
0 14318 5 1 1 14317
0 14319 7 1 2 30248 36697
0 14320 7 1 2 14318 14319
0 14321 5 1 1 14320
0 14322 7 1 2 14300 14321
0 14323 5 1 1 14322
0 14324 7 1 2 23131 14323
0 14325 5 1 1 14324
0 14326 7 1 2 14296 14325
0 14327 7 1 2 14277 14326
0 14328 5 1 1 14327
0 14329 7 1 2 28098 14328
0 14330 5 1 1 14329
0 14331 7 1 2 24692 26778
0 14332 5 1 1 14331
0 14333 7 1 2 6892 14332
0 14334 5 1 1 14333
0 14335 7 3 2 33426 28526
0 14336 7 1 2 33821 36930
0 14337 7 1 2 14334 14336
0 14338 5 1 1 14337
0 14339 7 1 2 24782 34613
0 14340 7 1 2 36719 14339
0 14341 5 1 1 14340
0 14342 7 1 2 14338 14341
0 14343 5 1 1 14342
0 14344 7 1 2 24201 14343
0 14345 5 1 1 14344
0 14346 7 1 2 33169 35355
0 14347 7 1 2 36831 14346
0 14348 5 1 1 14347
0 14349 7 1 2 14345 14348
0 14350 5 1 1 14349
0 14351 7 1 2 24112 14350
0 14352 5 1 1 14351
0 14353 7 1 2 34614 26437
0 14354 5 1 1 14353
0 14355 7 1 2 31016 31840
0 14356 5 1 1 14355
0 14357 7 1 2 14354 14356
0 14358 5 1 1 14357
0 14359 7 1 2 24783 35111
0 14360 7 1 2 33776 14359
0 14361 7 1 2 14358 14360
0 14362 5 1 1 14361
0 14363 7 1 2 14352 14362
0 14364 5 1 1 14363
0 14365 7 1 2 23355 14364
0 14366 5 1 1 14365
0 14367 7 1 2 24784 36910
0 14368 5 1 1 14367
0 14369 7 1 2 26438 2392
0 14370 7 1 2 33144 14369
0 14371 7 1 2 36161 14370
0 14372 5 1 1 14371
0 14373 7 1 2 14368 14372
0 14374 5 1 1 14373
0 14375 7 1 2 36487 14374
0 14376 5 1 1 14375
0 14377 7 1 2 27649 36922
0 14378 5 1 1 14377
0 14379 7 1 2 14376 14378
0 14380 5 2 1 14379
0 14381 7 1 2 35580 36933
0 14382 5 1 1 14381
0 14383 7 1 2 14366 14382
0 14384 5 1 1 14383
0 14385 7 1 2 22637 14384
0 14386 5 1 1 14385
0 14387 7 1 2 35948 36934
0 14388 5 1 1 14387
0 14389 7 2 2 23132 35245
0 14390 5 2 1 36935
0 14391 7 2 2 9572 26679
0 14392 5 9 1 36939
0 14393 7 2 2 29329 36941
0 14394 5 1 1 36950
0 14395 7 1 2 36937 14394
0 14396 5 8 1 14395
0 14397 7 1 2 32893 36952
0 14398 5 1 1 14397
0 14399 7 1 2 23356 26179
0 14400 7 1 2 32776 14399
0 14401 7 1 2 36759 14400
0 14402 5 1 1 14401
0 14403 7 1 2 14398 14402
0 14404 5 1 1 14403
0 14405 7 1 2 32109 14404
0 14406 5 1 1 14405
0 14407 7 3 2 35204 28576
0 14408 5 1 1 36960
0 14409 7 1 2 32918 36961
0 14410 7 1 2 32901 14409
0 14411 5 1 1 14410
0 14412 7 1 2 14406 14411
0 14413 5 1 1 14412
0 14414 7 1 2 36807 14413
0 14415 5 1 1 14414
0 14416 7 1 2 14388 14415
0 14417 7 1 2 14386 14416
0 14418 5 1 1 14417
0 14419 7 1 2 32730 14418
0 14420 5 1 1 14419
0 14421 7 1 2 14330 14420
0 14422 7 1 2 14252 14421
0 14423 5 1 1 14422
0 14424 7 1 2 29421 14423
0 14425 5 1 1 14424
0 14426 7 5 2 26321 32990
0 14427 7 2 2 32311 36963
0 14428 7 1 2 30339 32615
0 14429 7 1 2 30213 14428
0 14430 7 1 2 35093 27828
0 14431 7 1 2 14429 14430
0 14432 7 1 2 36968 14431
0 14433 5 1 1 14432
0 14434 7 1 2 14425 14433
0 14435 5 1 1 14434
0 14436 7 1 2 31626 14435
0 14437 5 1 1 14436
0 14438 7 1 2 27998 35672
0 14439 5 1 1 14438
0 14440 7 1 2 29898 32968
0 14441 5 1 1 14440
0 14442 7 1 2 14439 14441
0 14443 5 1 1 14442
0 14444 7 1 2 22638 14443
0 14445 5 1 1 14444
0 14446 7 3 2 29899 27421
0 14447 5 1 1 36970
0 14448 7 2 2 30340 35815
0 14449 5 1 1 36973
0 14450 7 1 2 14447 14449
0 14451 5 1 1 14450
0 14452 7 1 2 30649 14451
0 14453 5 1 1 14452
0 14454 7 1 2 14445 14453
0 14455 5 1 1 14454
0 14456 7 1 2 35238 14455
0 14457 5 1 1 14456
0 14458 7 1 2 31279 35613
0 14459 7 1 2 28159 14458
0 14460 7 1 2 32216 14459
0 14461 5 1 1 14460
0 14462 7 1 2 14457 14461
0 14463 5 1 1 14462
0 14464 7 1 2 23133 14463
0 14465 5 1 1 14464
0 14466 7 1 2 29900 31280
0 14467 7 1 2 28160 14466
0 14468 7 1 2 36951 14467
0 14469 5 1 1 14468
0 14470 7 1 2 14465 14469
0 14471 5 1 1 14470
0 14472 7 1 2 32110 32731
0 14473 7 1 2 14471 14472
0 14474 5 1 1 14473
0 14475 7 1 2 29229 36863
0 14476 5 1 1 14475
0 14477 7 1 2 30620 32625
0 14478 7 1 2 36211 14477
0 14479 5 1 1 14478
0 14480 7 1 2 14476 14479
0 14481 5 1 1 14480
0 14482 7 1 2 32553 33384
0 14483 7 1 2 35239 14482
0 14484 5 1 1 14483
0 14485 7 1 2 25078 36940
0 14486 5 2 1 14485
0 14487 7 6 2 26692 36975
0 14488 7 1 2 32530 33163
0 14489 7 1 2 36977 14488
0 14490 5 1 1 14489
0 14491 7 1 2 14484 14490
0 14492 5 1 1 14491
0 14493 7 1 2 14481 14492
0 14494 5 1 1 14493
0 14495 7 1 2 22747 32682
0 14496 5 1 1 14495
0 14497 7 1 2 33058 30627
0 14498 5 1 1 14497
0 14499 7 1 2 14496 14498
0 14500 5 1 1 14499
0 14501 7 1 2 22639 14500
0 14502 5 1 1 14501
0 14503 7 1 2 22748 32654
0 14504 5 1 1 14503
0 14505 7 1 2 28877 33059
0 14506 5 1 1 14505
0 14507 7 1 2 14504 14506
0 14508 5 2 1 14507
0 14509 7 1 2 30650 36983
0 14510 5 1 1 14509
0 14511 7 1 2 14502 14510
0 14512 5 1 1 14511
0 14513 7 2 2 24035 32554
0 14514 7 1 2 36985 36953
0 14515 7 1 2 14512 14514
0 14516 5 1 1 14515
0 14517 7 1 2 14494 14516
0 14518 7 1 2 14474 14517
0 14519 5 1 1 14518
0 14520 7 1 2 36808 14519
0 14521 5 1 1 14520
0 14522 7 4 2 24036 29957
0 14523 7 2 2 24332 36987
0 14524 7 4 2 24294 36991
0 14525 7 1 2 23578 28661
0 14526 7 1 2 30032 32345
0 14527 7 1 2 14525 14526
0 14528 7 1 2 32159 31537
0 14529 7 1 2 14527 14528
0 14530 7 1 2 36993 14529
0 14531 5 1 1 14530
0 14532 7 1 2 14521 14531
0 14533 5 1 1 14532
0 14534 7 1 2 31104 14533
0 14535 5 1 1 14534
0 14536 7 2 2 36809 36760
0 14537 7 1 2 26180 36997
0 14538 5 1 1 14537
0 14539 7 1 2 23049 36869
0 14540 7 1 2 36740 14539
0 14541 5 1 1 14540
0 14542 7 1 2 14538 14541
0 14543 5 1 1 14542
0 14544 7 1 2 24113 14543
0 14545 5 1 1 14544
0 14546 7 4 2 27809 26637
0 14547 7 1 2 35692 36999
0 14548 5 1 1 14547
0 14549 7 1 2 14545 14548
0 14550 5 1 1 14549
0 14551 7 1 2 35271 14550
0 14552 5 1 1 14551
0 14553 7 2 2 24202 35210
0 14554 7 5 2 24982 33470
0 14555 7 1 2 35852 32746
0 14556 7 1 2 31979 14555
0 14557 7 1 2 37005 14556
0 14558 7 1 2 37003 14557
0 14559 5 1 1 14558
0 14560 7 1 2 14552 14559
0 14561 5 1 1 14560
0 14562 7 1 2 22973 14561
0 14563 5 1 1 14562
0 14564 7 8 2 36810 36954
0 14565 5 1 1 37010
0 14566 7 2 2 25583 35211
0 14567 5 1 1 37018
0 14568 7 2 2 28591 37019
0 14569 5 1 1 37020
0 14570 7 1 2 26181 37021
0 14571 5 1 1 14570
0 14572 7 1 2 14565 14571
0 14573 5 1 1 14572
0 14574 7 1 2 35262 14573
0 14575 5 1 1 14574
0 14576 7 3 2 23579 23712
0 14577 7 2 2 28419 37022
0 14578 7 1 2 35802 32686
0 14579 7 2 2 37025 14578
0 14580 5 1 1 37027
0 14581 7 1 2 26182 37028
0 14582 5 1 1 14581
0 14583 7 1 2 14575 14582
0 14584 5 1 1 14583
0 14585 7 1 2 30044 14584
0 14586 5 1 1 14585
0 14587 7 1 2 14563 14586
0 14588 5 1 1 14587
0 14589 7 1 2 30172 14588
0 14590 5 1 1 14589
0 14591 7 2 2 28420 30270
0 14592 5 1 1 37029
0 14593 7 1 2 36277 37030
0 14594 5 1 1 14593
0 14595 7 1 2 14567 14592
0 14596 5 1 1 14595
0 14597 7 1 2 24983 7709
0 14598 7 1 2 14596 14597
0 14599 5 1 1 14598
0 14600 7 1 2 14594 14599
0 14601 5 1 1 14600
0 14602 7 1 2 35263 14601
0 14603 5 1 1 14602
0 14604 7 5 2 29062 34063
0 14605 7 1 2 26645 37031
0 14606 7 1 2 35216 14605
0 14607 5 1 1 14606
0 14608 7 1 2 14603 14607
0 14609 5 1 1 14608
0 14610 7 1 2 23134 14609
0 14611 5 1 1 14610
0 14612 7 1 2 32636 37026
0 14613 7 1 2 32168 14612
0 14614 5 1 1 14613
0 14615 7 1 2 14611 14614
0 14616 5 1 1 14615
0 14617 7 2 2 24203 14616
0 14618 5 1 1 37036
0 14619 7 1 2 36811 36978
0 14620 5 1 1 14619
0 14621 7 1 2 14620 14569
0 14622 5 1 1 14621
0 14623 7 1 2 35264 14622
0 14624 5 1 1 14623
0 14625 7 1 2 14624 14580
0 14626 5 1 1 14625
0 14627 7 1 2 24908 14626
0 14628 5 1 1 14627
0 14629 7 2 2 23713 27470
0 14630 7 1 2 32687 37038
0 14631 7 1 2 36998 14630
0 14632 5 1 1 14631
0 14633 7 1 2 14628 14632
0 14634 5 2 1 14633
0 14635 7 1 2 26183 37040
0 14636 5 1 1 14635
0 14637 7 1 2 14618 14636
0 14638 5 1 1 14637
0 14639 7 1 2 29906 14638
0 14640 5 1 1 14639
0 14641 7 1 2 14590 14640
0 14642 5 1 1 14641
0 14643 7 1 2 22851 14642
0 14644 5 1 1 14643
0 14645 7 1 2 28856 37041
0 14646 5 1 1 14645
0 14647 7 1 2 26567 36812
0 14648 5 1 1 14647
0 14649 7 1 2 23580 35298
0 14650 5 1 1 14649
0 14651 7 1 2 14648 14650
0 14652 5 1 1 14651
0 14653 7 1 2 26518 14652
0 14654 5 1 1 14653
0 14655 7 2 2 30090 26671
0 14656 7 1 2 36813 37042
0 14657 5 1 1 14656
0 14658 7 1 2 14654 14657
0 14659 5 1 1 14658
0 14660 7 2 2 27765 33504
0 14661 7 1 2 30173 37044
0 14662 7 1 2 14659 14661
0 14663 5 1 1 14662
0 14664 7 1 2 14646 14663
0 14665 5 1 1 14664
0 14666 7 1 2 26184 14665
0 14667 5 1 1 14666
0 14668 7 1 2 32580 37037
0 14669 5 1 1 14668
0 14670 7 1 2 14667 14669
0 14671 5 1 1 14670
0 14672 7 1 2 32515 14671
0 14673 5 1 1 14672
0 14674 7 2 2 30219 35754
0 14675 5 1 1 37046
0 14676 7 2 2 26497 33777
0 14677 5 2 1 37048
0 14678 7 1 2 14675 37050
0 14679 5 2 1 14678
0 14680 7 1 2 35086 37052
0 14681 5 1 1 14680
0 14682 7 1 2 23640 29816
0 14683 5 1 1 14682
0 14684 7 1 2 30543 14683
0 14685 5 2 1 14684
0 14686 7 4 2 22974 37054
0 14687 5 1 1 37056
0 14688 7 1 2 33145 37057
0 14689 5 1 1 14688
0 14690 7 1 2 14681 14689
0 14691 5 1 1 14690
0 14692 7 1 2 30174 14691
0 14693 5 1 1 14692
0 14694 7 2 2 35755 36088
0 14695 5 1 1 37060
0 14696 7 1 2 14695 14687
0 14697 5 4 1 14696
0 14698 7 1 2 36836 37062
0 14699 5 1 1 14698
0 14700 7 1 2 14693 14699
0 14701 5 1 1 14700
0 14702 7 2 2 34064 37045
0 14703 5 1 1 37066
0 14704 7 4 2 35417 32152
0 14705 7 1 2 27810 30805
0 14706 7 1 2 37068 14705
0 14707 5 1 1 14706
0 14708 7 1 2 14703 14707
0 14709 5 1 1 14708
0 14710 7 1 2 14701 14709
0 14711 5 1 1 14710
0 14712 7 1 2 14673 14711
0 14713 7 1 2 14644 14712
0 14714 5 1 1 14713
0 14715 7 1 2 22640 14714
0 14716 5 1 1 14715
0 14717 7 1 2 23581 33376
0 14718 7 1 2 35739 14717
0 14719 5 1 1 14718
0 14720 7 3 2 23423 26439
0 14721 7 1 2 33458 37072
0 14722 7 1 2 32567 14721
0 14723 5 1 1 14722
0 14724 7 1 2 14719 14723
0 14725 5 1 1 14724
0 14726 7 1 2 24984 14725
0 14727 5 1 1 14726
0 14728 7 1 2 33377 36278
0 14729 7 1 2 35740 14728
0 14730 5 1 1 14729
0 14731 7 1 2 14727 14730
0 14732 5 1 1 14731
0 14733 7 1 2 24295 14732
0 14734 5 1 1 14733
0 14735 7 1 2 34065 26655
0 14736 5 1 1 14735
0 14737 7 1 2 34080 14408
0 14738 5 1 1 14737
0 14739 7 1 2 32830 33567
0 14740 7 1 2 14738 14739
0 14741 7 1 2 14736 14740
0 14742 5 1 1 14741
0 14743 7 1 2 14734 14742
0 14744 5 1 1 14743
0 14745 7 1 2 34775 14744
0 14746 5 1 1 14745
0 14747 7 1 2 24114 34423
0 14748 7 1 2 36538 14747
0 14749 7 1 2 37011 14748
0 14750 5 1 1 14749
0 14751 7 1 2 14746 14750
0 14752 5 1 1 14751
0 14753 7 1 2 22749 14752
0 14754 5 1 1 14753
0 14755 7 2 2 26185 36814
0 14756 7 6 2 25079 25311
0 14757 7 3 2 29401 37077
0 14758 7 1 2 32874 37083
0 14759 5 1 1 14758
0 14760 7 1 2 23714 32763
0 14761 7 3 2 35696 14760
0 14762 5 1 1 37086
0 14763 7 1 2 14759 14762
0 14764 5 1 1 14763
0 14765 7 1 2 36942 14764
0 14766 5 1 1 14765
0 14767 7 1 2 26322 37087
0 14768 5 1 1 14767
0 14769 7 1 2 29901 31846
0 14770 7 1 2 31709 14769
0 14771 5 1 1 14770
0 14772 7 1 2 14768 14771
0 14773 5 1 1 14772
0 14774 7 1 2 24296 14773
0 14775 5 1 1 14774
0 14776 7 1 2 14766 14775
0 14777 5 1 1 14776
0 14778 7 1 2 37075 14777
0 14779 5 1 1 14778
0 14780 7 1 2 36698 37088
0 14781 5 1 1 14780
0 14782 7 2 2 24785 25227
0 14783 7 1 2 32747 28421
0 14784 7 2 2 37089 14783
0 14785 7 1 2 34424 36708
0 14786 7 1 2 37091 14785
0 14787 5 1 1 14786
0 14788 7 1 2 14781 14787
0 14789 5 1 1 14788
0 14790 7 1 2 23050 14789
0 14791 5 1 1 14790
0 14792 7 1 2 24985 34425
0 14793 7 1 2 36713 14792
0 14794 7 1 2 37092 14793
0 14795 5 1 1 14794
0 14796 7 1 2 14791 14795
0 14797 5 1 1 14796
0 14798 7 1 2 28468 14797
0 14799 5 1 1 14798
0 14800 7 1 2 14779 14799
0 14801 5 1 1 14800
0 14802 7 1 2 30837 14801
0 14803 5 1 1 14802
0 14804 7 1 2 14754 14803
0 14805 5 1 1 14804
0 14806 7 1 2 22641 14805
0 14807 5 1 1 14806
0 14808 7 1 2 36971 36955
0 14809 5 1 1 14808
0 14810 7 1 2 26716 36974
0 14811 5 1 1 14810
0 14812 7 1 2 14809 14811
0 14813 5 1 1 14812
0 14814 7 1 2 25711 30578
0 14815 7 2 2 36815 14814
0 14816 7 1 2 32111 37093
0 14817 7 1 2 14813 14816
0 14818 5 1 1 14817
0 14819 7 1 2 14807 14818
0 14820 5 1 1 14819
0 14821 7 1 2 32732 14820
0 14822 5 1 1 14821
0 14823 7 2 2 27897 29938
0 14824 7 2 2 31092 37095
0 14825 7 1 2 36761 37097
0 14826 5 1 1 14825
0 14827 7 1 2 28161 35578
0 14828 7 1 2 36979 14827
0 14829 5 1 1 14828
0 14830 7 1 2 14826 14829
0 14831 5 1 1 14830
0 14832 7 1 2 26186 14831
0 14833 5 1 1 14832
0 14834 7 1 2 28100 28776
0 14835 5 1 1 14834
0 14836 7 1 2 28322 27705
0 14837 5 1 1 14836
0 14838 7 1 2 29402 14837
0 14839 7 1 2 26717 14838
0 14840 7 1 2 14835 14839
0 14841 5 1 1 14840
0 14842 7 1 2 14833 14841
0 14843 5 1 1 14842
0 14844 7 1 2 32555 14843
0 14845 5 1 1 14844
0 14846 7 2 2 29738 36980
0 14847 7 1 2 27458 30451
0 14848 7 1 2 31871 14847
0 14849 7 1 2 37099 14848
0 14850 5 1 1 14849
0 14851 7 1 2 14845 14850
0 14852 5 1 1 14851
0 14853 7 1 2 36816 14852
0 14854 5 1 1 14853
0 14855 7 1 2 25080 32764
0 14856 7 3 2 26638 14855
0 14857 7 1 2 33561 37101
0 14858 5 1 1 14857
0 14859 7 1 2 13962 14858
0 14860 5 1 1 14859
0 14861 7 1 2 24204 37098
0 14862 7 1 2 14860 14861
0 14863 5 1 1 14862
0 14864 7 1 2 14854 14863
0 14865 5 1 1 14864
0 14866 7 1 2 33060 14865
0 14867 5 1 1 14866
0 14868 7 1 2 33361 37100
0 14869 5 1 1 14868
0 14870 7 1 2 28857 36956
0 14871 5 1 1 14870
0 14872 7 1 2 30175 26718
0 14873 5 1 1 14872
0 14874 7 1 2 14871 14873
0 14875 5 1 1 14874
0 14876 7 1 2 33146 14875
0 14877 5 1 1 14876
0 14878 7 1 2 14869 14877
0 14879 5 1 1 14878
0 14880 7 1 2 32655 37094
0 14881 7 1 2 14879 14880
0 14882 5 1 1 14881
0 14883 7 1 2 14867 14882
0 14884 7 1 2 14822 14883
0 14885 7 1 2 14716 14884
0 14886 5 1 1 14885
0 14887 7 1 2 22485 14886
0 14888 5 1 1 14887
0 14889 7 1 2 14535 14888
0 14890 5 1 1 14889
0 14891 7 1 2 23941 14890
0 14892 5 1 1 14891
0 14893 7 1 2 23817 14892
0 14894 7 1 2 14437 14893
0 14895 5 1 1 14894
0 14896 7 1 2 35762 35517
0 14897 5 1 1 14896
0 14898 7 2 2 26918 32616
0 14899 7 1 2 32677 37104
0 14900 5 1 1 14899
0 14901 7 1 2 14897 14900
0 14902 5 1 1 14901
0 14903 7 1 2 24115 14902
0 14904 5 1 1 14903
0 14905 7 1 2 23424 30341
0 14906 7 2 2 32733 14905
0 14907 7 1 2 29210 37106
0 14908 5 1 1 14907
0 14909 7 1 2 14904 14908
0 14910 5 1 1 14909
0 14911 7 1 2 22486 14910
0 14912 5 1 1 14911
0 14913 7 1 2 29063 32458
0 14914 5 1 1 14913
0 14915 7 1 2 23480 35008
0 14916 5 1 1 14915
0 14917 7 1 2 14914 14916
0 14918 5 1 1 14917
0 14919 7 1 2 36509 14918
0 14920 5 1 1 14919
0 14921 7 1 2 14912 14920
0 14922 5 1 1 14921
0 14923 7 1 2 37012 14922
0 14924 5 1 1 14923
0 14925 7 1 2 27528 28383
0 14926 5 2 1 14925
0 14927 7 1 2 24116 37063
0 14928 5 1 1 14927
0 14929 7 1 2 37108 14928
0 14930 5 2 1 14929
0 14931 7 1 2 25081 37110
0 14932 5 1 1 14931
0 14933 7 1 2 1780 29443
0 14934 5 16 1 14933
0 14935 7 3 2 37112 36745
0 14936 5 1 1 37128
0 14937 7 1 2 24117 37129
0 14938 5 1 1 14937
0 14939 7 1 2 14932 14938
0 14940 5 4 1 14939
0 14941 7 2 2 26006 37131
0 14942 7 2 2 27911 34066
0 14943 7 2 2 28885 37137
0 14944 7 1 2 23553 37139
0 14945 7 1 2 37135 14944
0 14946 5 1 1 14945
0 14947 7 1 2 14924 14946
0 14948 5 1 1 14947
0 14949 7 1 2 31675 14948
0 14950 5 1 1 14949
0 14951 7 1 2 27930 33854
0 14952 5 1 1 14951
0 14953 7 1 2 28221 31951
0 14954 5 1 1 14953
0 14955 7 3 2 14952 14954
0 14956 7 3 2 37141 37013
0 14957 7 1 2 33214 35518
0 14958 5 1 1 14957
0 14959 7 1 2 30383 37105
0 14960 5 1 1 14959
0 14961 7 1 2 14958 14960
0 14962 5 1 1 14961
0 14963 7 1 2 24118 14962
0 14964 5 1 1 14963
0 14965 7 1 2 25312 37107
0 14966 5 1 1 14965
0 14967 7 1 2 14964 14966
0 14968 5 1 1 14967
0 14969 7 1 2 37144 14968
0 14970 5 1 1 14969
0 14971 7 1 2 14950 14970
0 14972 5 1 1 14971
0 14973 7 1 2 31563 14972
0 14974 5 1 1 14973
0 14975 7 1 2 25584 34644
0 14976 7 1 2 34559 14975
0 14977 5 1 1 14976
0 14978 7 1 2 31968 37023
0 14979 7 1 2 35428 14978
0 14980 5 1 1 14979
0 14981 7 1 2 14977 14980
0 14982 5 1 1 14981
0 14983 7 1 2 25636 36165
0 14984 7 1 2 14982 14983
0 14985 5 1 1 14984
0 14986 7 1 2 28942 35566
0 14987 7 1 2 30762 30671
0 14988 7 1 2 14986 14987
0 14989 7 1 2 36623 14988
0 14990 5 1 1 14989
0 14991 7 1 2 14985 14990
0 14992 5 1 1 14991
0 14993 7 1 2 24333 14992
0 14994 5 1 1 14993
0 14995 7 1 2 26187 30064
0 14996 5 1 1 14995
0 14997 7 1 2 36938 14996
0 14998 5 1 1 14997
0 14999 7 2 2 29422 31627
0 15000 7 1 2 23582 30342
0 15001 7 1 2 37147 15000
0 15002 7 1 2 14998 15001
0 15003 5 1 1 15002
0 15004 7 1 2 14994 15003
0 15005 5 1 1 15004
0 15006 7 1 2 25313 15005
0 15007 5 1 1 15006
0 15008 7 2 2 23357 23583
0 15009 7 1 2 30744 37149
0 15010 7 1 2 32948 15009
0 15011 7 1 2 36957 15010
0 15012 5 1 1 15011
0 15013 7 1 2 15007 15012
0 15014 5 1 1 15013
0 15015 7 1 2 24601 15014
0 15016 5 1 1 15015
0 15017 7 2 2 30343 30456
0 15018 7 1 2 23584 37151
0 15019 7 1 2 35593 15018
0 15020 7 1 2 36958 15019
0 15021 5 1 1 15020
0 15022 7 1 2 15016 15021
0 15023 5 1 1 15022
0 15024 7 1 2 25380 15023
0 15025 5 1 1 15024
0 15026 7 1 2 22642 31165
0 15027 5 1 1 15026
0 15028 7 1 2 27320 30651
0 15029 5 1 1 15028
0 15030 7 1 2 15027 15029
0 15031 5 1 1 15030
0 15032 7 1 2 22487 15031
0 15033 5 1 1 15032
0 15034 7 1 2 27912 36158
0 15035 5 1 1 15034
0 15036 7 1 2 15033 15035
0 15037 5 2 1 15036
0 15038 7 2 2 36959 37153
0 15039 7 1 2 23715 32977
0 15040 7 1 2 36769 15039
0 15041 7 1 2 37155 15040
0 15042 5 1 1 15041
0 15043 7 1 2 15025 15042
0 15044 5 1 1 15043
0 15045 7 1 2 24986 15044
0 15046 5 1 1 15045
0 15047 7 1 2 36279 30745
0 15048 7 1 2 26919 15047
0 15049 7 1 2 37156 15048
0 15050 5 1 1 15049
0 15051 7 1 2 15046 15050
0 15052 5 1 1 15051
0 15053 7 1 2 25442 15052
0 15054 5 1 1 15053
0 15055 7 2 2 23716 24119
0 15056 7 1 2 31830 37157
0 15057 7 1 2 37014 15056
0 15058 7 1 2 37154 15057
0 15059 5 1 1 15058
0 15060 7 1 2 15054 15059
0 15061 5 1 1 15060
0 15062 7 1 2 25503 15061
0 15063 5 1 1 15062
0 15064 7 2 2 29958 29617
0 15065 7 2 2 30499 37159
0 15066 5 2 1 37161
0 15067 7 4 2 23641 32991
0 15068 7 1 2 32869 37165
0 15069 5 1 1 15068
0 15070 7 1 2 37163 15069
0 15071 5 1 1 15070
0 15072 7 2 2 22643 15071
0 15073 5 1 1 37169
0 15074 7 1 2 35432 30299
0 15075 5 1 1 15074
0 15076 7 1 2 15073 15075
0 15077 5 1 1 15076
0 15078 7 1 2 24465 15077
0 15079 5 1 1 15078
0 15080 7 2 2 31981 36994
0 15081 7 1 2 28058 37171
0 15082 5 1 1 15081
0 15083 7 1 2 15079 15082
0 15084 5 1 1 15083
0 15085 7 1 2 25082 15084
0 15086 5 1 1 15085
0 15087 7 2 2 31676 30147
0 15088 7 1 2 33532 35212
0 15089 7 1 2 37173 15088
0 15090 5 1 1 15089
0 15091 7 1 2 15086 15090
0 15092 5 1 1 15091
0 15093 7 1 2 37067 15092
0 15094 5 1 1 15093
0 15095 7 1 2 24909 15094
0 15096 7 1 2 15063 15095
0 15097 5 1 1 15096
0 15098 7 1 2 33202 35383
0 15099 5 1 1 15098
0 15100 7 1 2 29211 33815
0 15101 5 1 1 15100
0 15102 7 1 2 15099 15101
0 15103 5 1 1 15102
0 15104 7 1 2 22488 15103
0 15105 5 1 1 15104
0 15106 7 1 2 33816 36676
0 15107 5 1 1 15106
0 15108 7 1 2 15105 15107
0 15109 5 1 1 15108
0 15110 7 1 2 23425 15109
0 15111 5 1 1 15110
0 15112 7 2 2 22489 28715
0 15113 7 1 2 28077 29875
0 15114 7 1 2 37175 15113
0 15115 5 1 1 15114
0 15116 7 1 2 15111 15115
0 15117 5 1 1 15116
0 15118 7 1 2 37015 15117
0 15119 5 1 1 15118
0 15120 7 1 2 24205 36777
0 15121 5 1 1 15120
0 15122 7 2 2 32018 29632
0 15123 5 1 1 37177
0 15124 7 1 2 15121 15123
0 15125 5 9 1 15124
0 15126 7 2 2 26097 37179
0 15127 7 3 2 26007 37188
0 15128 7 1 2 37190 37140
0 15129 5 1 1 15128
0 15130 7 1 2 15119 15129
0 15131 5 1 1 15130
0 15132 7 1 2 31677 15131
0 15133 5 1 1 15132
0 15134 7 1 2 34921 28747
0 15135 5 1 1 15134
0 15136 7 1 2 27756 33817
0 15137 5 1 1 15136
0 15138 7 1 2 15135 15137
0 15139 5 1 1 15138
0 15140 7 1 2 37145 15139
0 15141 5 1 1 15140
0 15142 7 1 2 15133 15141
0 15143 5 1 1 15142
0 15144 7 1 2 33500 15143
0 15145 5 1 1 15144
0 15146 7 1 2 22975 15145
0 15147 5 1 1 15146
0 15148 7 1 2 24786 15147
0 15149 7 1 2 15097 15148
0 15150 5 1 1 15149
0 15151 7 1 2 14974 15150
0 15152 5 1 1 15151
0 15153 7 1 2 24693 15152
0 15154 5 1 1 15153
0 15155 7 2 2 23554 26920
0 15156 7 1 2 35514 37193
0 15157 5 1 1 15156
0 15158 7 1 2 14306 15157
0 15159 5 2 1 15158
0 15160 7 1 2 29138 37195
0 15161 5 1 1 15160
0 15162 7 1 2 35915 30392
0 15163 7 1 2 32626 15162
0 15164 5 1 1 15163
0 15165 7 1 2 15161 15164
0 15166 5 1 1 15165
0 15167 7 1 2 37016 15166
0 15168 5 1 1 15167
0 15169 7 1 2 37113 36778
0 15170 5 1 1 15169
0 15171 7 1 2 22976 37178
0 15172 5 1 1 15171
0 15173 7 1 2 15170 15172
0 15174 5 3 1 15173
0 15175 7 1 2 30631 37138
0 15176 7 1 2 31831 15175
0 15177 7 1 2 37197 15176
0 15178 5 1 1 15177
0 15179 7 1 2 15168 15178
0 15180 5 1 1 15179
0 15181 7 1 2 31678 15180
0 15182 5 1 1 15181
0 15183 7 1 2 25314 37196
0 15184 5 1 1 15183
0 15185 7 2 2 32230 32617
0 15186 7 1 2 32318 37200
0 15187 5 1 1 15186
0 15188 7 1 2 15184 15187
0 15189 5 1 1 15188
0 15190 7 1 2 37146 15189
0 15191 5 1 1 15190
0 15192 7 1 2 15182 15191
0 15193 5 1 1 15192
0 15194 7 1 2 32556 15193
0 15195 5 1 1 15194
0 15196 7 1 2 35673 32009
0 15197 5 1 1 15196
0 15198 7 1 2 30652 32875
0 15199 5 1 1 15198
0 15200 7 1 2 15197 15199
0 15201 5 1 1 15200
0 15202 7 1 2 22490 15201
0 15203 5 1 1 15202
0 15204 7 2 2 26008 32010
0 15205 7 1 2 26098 27913
0 15206 7 1 2 37202 15205
0 15207 5 1 1 15206
0 15208 7 1 2 15203 15207
0 15209 5 1 1 15208
0 15210 7 1 2 27321 15209
0 15211 5 1 1 15210
0 15212 7 1 2 22852 36882
0 15213 5 1 1 15212
0 15214 7 1 2 4691 15213
0 15215 5 1 1 15214
0 15216 7 1 2 35594 15215
0 15217 5 1 1 15216
0 15218 7 1 2 15211 15217
0 15219 5 1 1 15218
0 15220 7 4 2 32734 37017
0 15221 7 1 2 25381 37204
0 15222 7 1 2 15219 15221
0 15223 5 1 1 15222
0 15224 7 1 2 15195 15223
0 15225 5 1 1 15224
0 15226 7 1 2 29939 15225
0 15227 5 1 1 15226
0 15228 7 1 2 25812 15227
0 15229 7 1 2 15154 15228
0 15230 5 1 1 15229
0 15231 7 1 2 14895 15230
0 15232 5 1 1 15231
0 15233 7 3 2 28261 29637
0 15234 7 1 2 36775 37150
0 15235 7 1 2 29004 15234
0 15236 7 1 2 32135 15235
0 15237 7 1 2 31444 15236
0 15238 5 1 1 15237
0 15239 7 2 2 33568 37053
0 15240 5 1 1 37211
0 15241 7 1 2 23051 36714
0 15242 7 1 2 30914 15241
0 15243 5 1 1 15242
0 15244 7 1 2 15240 15243
0 15245 5 2 1 15244
0 15246 7 1 2 26009 28841
0 15247 7 1 2 37213 15246
0 15248 5 1 1 15247
0 15249 7 1 2 15238 15248
0 15250 5 1 1 15249
0 15251 7 1 2 24694 15250
0 15252 5 1 1 15251
0 15253 7 2 2 23426 28162
0 15254 7 1 2 32491 37215
0 15255 5 1 1 15254
0 15256 7 1 2 35393 32972
0 15257 5 1 1 15256
0 15258 7 1 2 15255 15257
0 15259 5 1 1 15258
0 15260 7 1 2 35997 36736
0 15261 7 1 2 15259 15260
0 15262 5 1 1 15261
0 15263 7 1 2 15252 15262
0 15264 5 1 1 15263
0 15265 7 1 2 23135 15264
0 15266 5 1 1 15265
0 15267 7 2 2 33562 31097
0 15268 7 1 2 28858 37217
0 15269 5 1 1 15268
0 15270 7 1 2 30176 31074
0 15271 7 1 2 36715 15270
0 15272 5 1 1 15271
0 15273 7 1 2 15269 15272
0 15274 5 1 1 15273
0 15275 7 1 2 26099 15274
0 15276 7 1 2 28842 15275
0 15277 5 1 1 15276
0 15278 7 1 2 34270 37218
0 15279 7 1 2 35950 15278
0 15280 5 1 1 15279
0 15281 7 1 2 15277 15280
0 15282 5 1 1 15281
0 15283 7 1 2 30564 15282
0 15284 5 1 1 15283
0 15285 7 1 2 15266 15284
0 15286 5 1 1 15285
0 15287 7 1 2 25914 15286
0 15288 5 1 1 15287
0 15289 7 1 2 30790 31093
0 15290 5 1 1 15289
0 15291 7 1 2 33121 15290
0 15292 5 1 1 15291
0 15293 7 1 2 24120 36720
0 15294 5 1 1 15293
0 15295 7 1 2 35689 37000
0 15296 5 1 1 15295
0 15297 7 1 2 15294 15296
0 15298 5 1 1 15297
0 15299 7 1 2 15292 15298
0 15300 5 1 1 15299
0 15301 7 1 2 33569 1394
0 15302 7 2 2 11514 15301
0 15303 7 1 2 28770 30300
0 15304 7 1 2 31380 15303
0 15305 7 1 2 37219 15304
0 15306 5 1 1 15305
0 15307 7 1 2 15300 15306
0 15308 5 1 1 15307
0 15309 7 1 2 26188 15308
0 15310 5 1 1 15309
0 15311 7 2 2 25083 36716
0 15312 5 1 1 37221
0 15313 7 1 2 33570 26618
0 15314 5 1 1 15313
0 15315 7 1 2 15312 15314
0 15316 5 2 1 15315
0 15317 7 4 2 27524 29618
0 15318 7 1 2 27024 28771
0 15319 7 1 2 37225 15318
0 15320 7 1 2 37223 15319
0 15321 5 1 1 15320
0 15322 7 1 2 15310 15321
0 15323 5 1 1 15322
0 15324 7 1 2 22644 15323
0 15325 5 1 1 15324
0 15326 7 1 2 37226 37222
0 15327 5 2 1 15326
0 15328 7 1 2 23136 37214
0 15329 5 1 1 15328
0 15330 7 1 2 37229 15329
0 15331 5 2 1 15330
0 15332 7 1 2 33126 37231
0 15333 5 1 1 15332
0 15334 7 1 2 15325 15333
0 15335 5 1 1 15334
0 15336 7 1 2 28735 15335
0 15337 5 1 1 15336
0 15338 7 1 2 30943 36661
0 15339 5 1 1 15338
0 15340 7 2 2 22853 32581
0 15341 7 1 2 23427 32444
0 15342 7 1 2 37233 15341
0 15343 5 1 1 15342
0 15344 7 1 2 15339 15343
0 15345 5 1 1 15344
0 15346 7 1 2 36721 15345
0 15347 5 1 1 15346
0 15348 7 1 2 22750 35600
0 15349 5 1 1 15348
0 15350 7 1 2 33362 33818
0 15351 5 1 1 15350
0 15352 7 1 2 15349 15351
0 15353 5 1 1 15352
0 15354 7 1 2 31883 36931
0 15355 7 1 2 15353 15354
0 15356 5 1 1 15355
0 15357 7 1 2 15347 15356
0 15358 5 1 1 15357
0 15359 7 1 2 26189 28910
0 15360 7 1 2 15358 15359
0 15361 5 1 1 15360
0 15362 7 1 2 15337 15361
0 15363 7 1 2 15288 15362
0 15364 5 1 1 15363
0 15365 7 1 2 37208 15364
0 15366 5 1 1 15365
0 15367 7 4 2 24466 33721
0 15368 5 1 1 37235
0 15369 7 1 2 32339 15368
0 15370 5 3 1 15369
0 15371 7 1 2 36943 37239
0 15372 5 1 1 15371
0 15373 7 1 2 31458 26619
0 15374 5 1 1 15373
0 15375 7 3 2 23818 26323
0 15376 7 1 2 22491 37242
0 15377 5 1 1 15376
0 15378 7 1 2 15374 15377
0 15379 5 1 1 15378
0 15380 7 1 2 24297 15379
0 15381 5 1 1 15380
0 15382 7 1 2 15372 15381
0 15383 5 1 1 15382
0 15384 7 1 2 32472 32843
0 15385 5 1 1 15384
0 15386 7 1 2 33914 34293
0 15387 5 1 1 15386
0 15388 7 1 2 15385 15387
0 15389 5 1 1 15388
0 15390 7 1 2 22854 15389
0 15391 5 1 1 15390
0 15392 7 2 2 25915 35356
0 15393 7 1 2 32445 37245
0 15394 5 1 1 15393
0 15395 7 1 2 15391 15394
0 15396 5 1 1 15395
0 15397 7 1 2 22645 15396
0 15398 7 1 2 15383 15397
0 15399 5 1 1 15398
0 15400 7 5 2 25813 36981
0 15401 7 1 2 34205 35582
0 15402 5 1 1 15401
0 15403 7 1 2 36170 32978
0 15404 5 1 1 15403
0 15405 7 1 2 15402 15404
0 15406 5 1 1 15405
0 15407 7 1 2 24602 15406
0 15408 7 1 2 37247 15407
0 15409 5 1 1 15408
0 15410 7 1 2 15399 15409
0 15411 5 1 1 15410
0 15412 7 1 2 23358 15411
0 15413 5 1 1 15412
0 15414 7 1 2 34206 32748
0 15415 7 1 2 31679 15414
0 15416 7 1 2 29005 15415
0 15417 7 1 2 37248 15416
0 15418 5 1 1 15417
0 15419 7 1 2 15413 15418
0 15420 5 1 1 15419
0 15421 7 1 2 24206 15420
0 15422 5 1 1 15421
0 15423 7 2 2 28059 30435
0 15424 5 1 1 37252
0 15425 7 1 2 33888 15424
0 15426 5 1 1 15425
0 15427 7 1 2 36662 15426
0 15428 5 1 1 15427
0 15429 7 1 2 32446 33042
0 15430 7 1 2 33249 15429
0 15431 5 1 1 15430
0 15432 7 1 2 15428 15431
0 15433 5 1 1 15432
0 15434 7 1 2 32420 26702
0 15435 7 1 2 36964 15434
0 15436 7 1 2 15433 15435
0 15437 5 1 1 15436
0 15438 7 1 2 15422 15437
0 15439 5 1 1 15438
0 15440 7 1 2 23273 15439
0 15441 5 1 1 15440
0 15442 7 1 2 25382 26687
0 15443 7 1 2 30752 15442
0 15444 5 1 1 15443
0 15445 7 1 2 32844 35756
0 15446 7 1 2 36705 15445
0 15447 5 1 1 15446
0 15448 7 1 2 15444 15447
0 15449 5 1 1 15448
0 15450 7 1 2 23137 15449
0 15451 5 1 1 15450
0 15452 7 1 2 25084 24121
0 15453 7 2 2 36944 15452
0 15454 7 4 2 24207 37254
0 15455 5 1 1 37256
0 15456 7 1 2 34294 37257
0 15457 5 1 1 15456
0 15458 7 1 2 15451 15457
0 15459 5 1 1 15458
0 15460 7 1 2 23359 15459
0 15461 5 1 1 15460
0 15462 7 2 2 30772 36965
0 15463 7 1 2 30734 31070
0 15464 7 1 2 37260 15463
0 15465 5 1 1 15464
0 15466 7 1 2 15461 15465
0 15467 5 1 1 15466
0 15468 7 1 2 22646 15467
0 15469 5 1 1 15468
0 15470 7 1 2 24603 30727
0 15471 7 1 2 31071 15470
0 15472 7 1 2 37261 15471
0 15473 5 1 1 15472
0 15474 7 1 2 15469 15473
0 15475 5 1 1 15474
0 15476 7 2 2 22492 28274
0 15477 7 1 2 29006 37262
0 15478 7 1 2 15475 15477
0 15479 5 1 1 15478
0 15480 7 1 2 15441 15479
0 15481 5 1 1 15480
0 15482 7 1 2 23717 15481
0 15483 5 1 1 15482
0 15484 7 3 2 27180 31509
0 15485 7 5 2 23642 28422
0 15486 7 2 2 27511 37267
0 15487 5 1 1 37272
0 15488 7 2 2 22493 31426
0 15489 7 1 2 27720 31324
0 15490 7 1 2 37274 15489
0 15491 7 1 2 37273 15490
0 15492 5 1 1 15491
0 15493 7 1 2 30322 34271
0 15494 5 1 1 15493
0 15495 7 1 2 32438 29586
0 15496 7 1 2 37275 15495
0 15497 5 1 1 15496
0 15498 7 1 2 15494 15497
0 15499 5 1 1 15498
0 15500 7 1 2 24208 36982
0 15501 7 1 2 15499 15500
0 15502 5 1 1 15501
0 15503 7 1 2 15492 15502
0 15504 5 1 1 15503
0 15505 7 1 2 37264 15504
0 15506 5 1 1 15505
0 15507 7 3 2 26100 36945
0 15508 7 1 2 28488 37276
0 15509 5 1 1 15508
0 15510 7 3 2 30763 29723
0 15511 5 1 1 37279
0 15512 7 1 2 5864 15511
0 15513 5 1 1 15512
0 15514 7 1 2 23138 14263
0 15515 7 1 2 15513 15514
0 15516 5 1 1 15515
0 15517 7 1 2 15509 15516
0 15518 5 3 1 15517
0 15519 7 2 2 28345 34804
0 15520 5 1 1 37285
0 15521 7 2 2 31680 36055
0 15522 5 1 1 37287
0 15523 7 1 2 15520 15522
0 15524 5 6 1 15523
0 15525 7 1 2 33037 37289
0 15526 7 1 2 37282 15525
0 15527 5 1 1 15526
0 15528 7 1 2 15506 15527
0 15529 7 1 2 15483 15528
0 15530 5 1 1 15529
0 15531 7 1 2 32582 15530
0 15532 5 1 1 15531
0 15533 7 3 2 26010 27238
0 15534 7 5 2 26101 37280
0 15535 7 1 2 37295 37298
0 15536 5 2 1 15535
0 15537 7 1 2 34645 31534
0 15538 5 1 1 15537
0 15539 7 1 2 37303 15538
0 15540 5 1 1 15539
0 15541 7 1 2 23139 15540
0 15542 5 1 1 15541
0 15543 7 1 2 34475 37258
0 15544 5 1 1 15543
0 15545 7 1 2 15542 15544
0 15546 5 1 1 15545
0 15547 7 1 2 24695 15546
0 15548 5 1 1 15547
0 15549 7 2 2 29959 36762
0 15550 7 1 2 32784 37305
0 15551 5 1 1 15550
0 15552 7 1 2 15548 15551
0 15553 5 1 1 15552
0 15554 7 1 2 23428 15553
0 15555 5 1 1 15554
0 15556 7 2 2 33388 36966
0 15557 7 1 2 32786 30672
0 15558 7 1 2 37307 15557
0 15559 5 1 1 15558
0 15560 7 1 2 15555 15559
0 15561 5 1 1 15560
0 15562 7 1 2 29689 15561
0 15563 5 1 1 15562
0 15564 7 4 2 24298 29960
0 15565 7 1 2 26620 37309
0 15566 5 1 1 15565
0 15567 7 1 2 15455 15566
0 15568 5 1 1 15567
0 15569 7 1 2 23429 15568
0 15570 5 1 1 15569
0 15571 7 1 2 27562 37299
0 15572 5 1 1 15571
0 15573 7 1 2 15570 15572
0 15574 5 2 1 15573
0 15575 7 2 2 28772 33738
0 15576 5 1 1 37315
0 15577 7 1 2 27701 31649
0 15578 5 1 1 15577
0 15579 7 1 2 15576 15578
0 15580 5 1 1 15579
0 15581 7 1 2 27976 15580
0 15582 7 1 2 37313 15581
0 15583 5 1 1 15582
0 15584 7 1 2 15563 15583
0 15585 5 1 1 15584
0 15586 7 1 2 28163 15585
0 15587 5 1 1 15586
0 15588 7 2 2 23718 32805
0 15589 7 1 2 29309 37314
0 15590 5 1 1 15589
0 15591 7 2 2 35248 31812
0 15592 7 1 2 37319 37306
0 15593 5 1 1 15592
0 15594 7 1 2 15590 15593
0 15595 5 1 1 15594
0 15596 7 1 2 37317 15595
0 15597 5 1 1 15596
0 15598 7 1 2 29876 37281
0 15599 5 2 1 15598
0 15600 7 1 2 33463 28691
0 15601 5 1 1 15600
0 15602 7 1 2 37321 15601
0 15603 5 1 1 15602
0 15604 7 1 2 23140 15603
0 15605 5 1 1 15604
0 15606 7 1 2 26011 37259
0 15607 5 1 1 15606
0 15608 7 1 2 15605 15607
0 15609 5 1 1 15608
0 15610 7 1 2 30984 34805
0 15611 7 1 2 29252 15610
0 15612 7 1 2 15609 15611
0 15613 5 1 1 15612
0 15614 7 1 2 15597 15613
0 15615 7 1 2 15587 15614
0 15616 5 1 1 15615
0 15617 7 1 2 29007 15616
0 15618 5 1 1 15617
0 15619 7 2 2 30115 34671
0 15620 5 1 1 37323
0 15621 7 1 2 24604 34806
0 15622 5 1 1 15621
0 15623 7 1 2 15620 15622
0 15624 5 1 1 15623
0 15625 7 3 2 27977 15624
0 15626 5 1 1 37325
0 15627 7 1 2 33291 31590
0 15628 5 1 1 15627
0 15629 7 1 2 15626 15628
0 15630 5 4 1 15629
0 15631 7 1 2 31083 37328
0 15632 5 1 1 15631
0 15633 7 1 2 30621 30393
0 15634 5 1 1 15633
0 15635 7 1 2 26012 31580
0 15636 5 1 1 15635
0 15637 7 1 2 15634 15636
0 15638 5 1 1 15637
0 15639 7 1 2 37290 15638
0 15640 5 1 1 15639
0 15641 7 3 2 31681 31608
0 15642 7 1 2 26013 28364
0 15643 7 1 2 36627 15642
0 15644 7 1 2 37332 15643
0 15645 5 1 1 15644
0 15646 7 2 2 30697 27872
0 15647 7 2 2 25712 31395
0 15648 7 1 2 30436 37337
0 15649 7 1 2 37335 15648
0 15650 5 1 1 15649
0 15651 7 1 2 15645 15650
0 15652 7 1 2 15640 15651
0 15653 7 1 2 15632 15652
0 15654 5 1 1 15653
0 15655 7 1 2 15654 37283
0 15656 5 1 1 15655
0 15657 7 1 2 28773 34107
0 15658 5 1 1 15657
0 15659 7 1 2 32790 28243
0 15660 5 1 1 15659
0 15661 7 1 2 15658 15660
0 15662 5 1 1 15661
0 15663 7 1 2 36946 15662
0 15664 5 1 1 15663
0 15665 7 1 2 28244 26661
0 15666 7 1 2 32806 15665
0 15667 5 1 1 15666
0 15668 7 1 2 15664 15667
0 15669 5 1 1 15668
0 15670 7 1 2 27525 37209
0 15671 7 1 2 15669 15670
0 15672 5 1 1 15671
0 15673 7 1 2 15656 15672
0 15674 5 1 1 15673
0 15675 7 1 2 28736 15674
0 15676 5 1 1 15675
0 15677 7 1 2 28866 5436
0 15678 5 1 1 15677
0 15679 7 1 2 36947 15678
0 15680 5 1 1 15679
0 15681 7 1 2 28859 26662
0 15682 5 1 1 15681
0 15683 7 1 2 15680 15682
0 15684 5 1 1 15683
0 15685 7 1 2 23819 24209
0 15686 7 1 2 34527 15685
0 15687 7 2 2 15684 15686
0 15688 7 1 2 33869 37339
0 15689 5 1 1 15688
0 15690 7 1 2 29380 37340
0 15691 5 1 1 15690
0 15692 7 2 2 32583 37329
0 15693 7 1 2 37341 37284
0 15694 5 1 1 15693
0 15695 7 1 2 15691 15694
0 15696 5 1 1 15695
0 15697 7 1 2 28827 15696
0 15698 5 1 1 15697
0 15699 7 1 2 15689 15698
0 15700 7 1 2 15676 15699
0 15701 7 1 2 15618 15700
0 15702 7 1 2 15532 15701
0 15703 5 1 1 15702
0 15704 7 1 2 36817 15703
0 15705 5 1 1 15704
0 15706 7 1 2 15366 15705
0 15707 5 1 1 15706
0 15708 7 1 2 29117 15707
0 15709 5 1 1 15708
0 15710 7 2 2 23585 26463
0 15711 7 1 2 35734 37343
0 15712 5 1 1 15711
0 15713 7 1 2 33771 30583
0 15714 7 1 2 36888 15713
0 15715 5 1 1 15714
0 15716 7 1 2 15712 15715
0 15717 5 1 1 15716
0 15718 7 1 2 24987 15717
0 15719 5 1 1 15718
0 15720 7 1 2 9884 36871
0 15721 5 1 1 15720
0 15722 7 1 2 5636 28492
0 15723 5 1 1 15722
0 15724 7 1 2 35290 15723
0 15725 7 1 2 15721 15724
0 15726 5 1 1 15725
0 15727 7 1 2 15719 15726
0 15728 5 1 1 15727
0 15729 7 1 2 32331 15728
0 15730 5 1 1 15729
0 15731 7 1 2 30158 36870
0 15732 5 1 1 15731
0 15733 7 1 2 25504 36818
0 15734 7 1 2 36885 15733
0 15735 5 1 1 15734
0 15736 7 1 2 15732 15735
0 15737 5 1 1 15736
0 15738 7 1 2 24910 31459
0 15739 7 1 2 15737 15738
0 15740 5 1 1 15739
0 15741 7 1 2 15730 15740
0 15742 5 1 1 15741
0 15743 7 1 2 23481 15742
0 15744 5 1 1 15743
0 15745 7 8 2 23820 26519
0 15746 7 2 2 22494 37345
0 15747 5 1 1 37353
0 15748 7 1 2 31460 26626
0 15749 5 1 1 15748
0 15750 7 1 2 15747 15749
0 15751 5 1 1 15750
0 15752 7 1 2 32719 37076
0 15753 7 1 2 15751 15752
0 15754 5 1 1 15753
0 15755 7 1 2 15744 15754
0 15756 5 1 1 15755
0 15757 7 1 2 24299 15756
0 15758 5 1 1 15757
0 15759 7 1 2 32332 36699
0 15760 5 1 1 15759
0 15761 7 1 2 31461 28423
0 15762 7 1 2 36709 15761
0 15763 5 1 1 15762
0 15764 7 1 2 15760 15763
0 15765 5 1 1 15764
0 15766 7 1 2 28469 15765
0 15767 5 1 1 15766
0 15768 7 1 2 33482 31462
0 15769 7 1 2 36874 15768
0 15770 5 1 1 15769
0 15771 7 1 2 15767 15770
0 15772 5 1 1 15771
0 15773 7 1 2 23052 15772
0 15774 5 1 1 15773
0 15775 7 2 2 24988 31463
0 15776 5 1 1 37355
0 15777 7 1 2 34870 37356
0 15778 7 1 2 36879 15777
0 15779 5 1 1 15778
0 15780 7 1 2 15774 15779
0 15781 5 1 1 15780
0 15782 7 1 2 32735 15781
0 15783 5 1 1 15782
0 15784 7 1 2 15758 15783
0 15785 5 1 1 15784
0 15786 7 1 2 23274 15785
0 15787 5 1 1 15786
0 15788 7 1 2 37205 37263
0 15789 5 1 1 15788
0 15790 7 1 2 15787 15789
0 15791 5 1 1 15790
0 15792 7 1 2 32035 15791
0 15793 5 1 1 15792
0 15794 7 1 2 24696 33650
0 15795 7 1 2 35339 15794
0 15796 7 1 2 37206 15795
0 15797 5 1 1 15796
0 15798 7 1 2 15793 15797
0 15799 5 1 1 15798
0 15800 7 1 2 31682 15799
0 15801 5 1 1 15800
0 15802 7 7 2 25585 37001
0 15803 5 1 1 37357
0 15804 7 1 2 37358 36984
0 15805 5 1 1 15804
0 15806 7 1 2 32248 32736
0 15807 7 1 2 36722 15806
0 15808 5 1 1 15807
0 15809 7 1 2 15805 15808
0 15810 5 1 1 15809
0 15811 7 2 2 22495 27239
0 15812 7 1 2 24210 27898
0 15813 7 1 2 37364 15812
0 15814 7 1 2 15810 15813
0 15815 5 1 1 15814
0 15816 7 1 2 26190 37249
0 15817 5 1 1 15816
0 15818 7 1 2 24211 35899
0 15819 7 1 2 37268 15818
0 15820 5 1 1 15819
0 15821 7 1 2 15817 15820
0 15822 5 1 1 15821
0 15823 7 1 2 37142 15822
0 15824 5 1 1 15823
0 15825 7 1 2 31969 36757
0 15826 7 1 2 34845 15825
0 15827 5 1 1 15826
0 15828 7 1 2 15824 15827
0 15829 5 1 1 15828
0 15830 7 1 2 32249 15829
0 15831 5 1 1 15830
0 15832 7 1 2 22496 34169
0 15833 7 1 2 32410 36962
0 15834 7 1 2 15832 15833
0 15835 5 1 1 15834
0 15836 7 1 2 15831 15835
0 15837 5 1 1 15836
0 15838 7 1 2 32737 36819
0 15839 7 1 2 15837 15838
0 15840 5 1 1 15839
0 15841 7 1 2 15815 15840
0 15842 7 1 2 15801 15841
0 15843 5 1 1 15842
0 15844 7 1 2 23719 15843
0 15845 5 1 1 15844
0 15846 7 1 2 27978 35471
0 15847 5 2 1 15846
0 15848 7 3 2 22751 34622
0 15849 7 1 2 29646 37368
0 15850 5 1 1 15849
0 15851 7 1 2 37366 15850
0 15852 5 1 1 15851
0 15853 7 1 2 37207 15852
0 15854 5 1 1 15853
0 15855 7 2 2 29317 31233
0 15856 7 3 2 35303 33471
0 15857 7 1 2 27811 28460
0 15858 7 1 2 37373 15857
0 15859 7 1 2 37371 15858
0 15860 5 1 1 15859
0 15861 7 1 2 15854 15860
0 15862 5 1 1 15861
0 15863 7 1 2 34807 15862
0 15864 5 1 1 15863
0 15865 7 1 2 15845 15864
0 15866 5 1 1 15865
0 15867 7 1 2 32932 15866
0 15868 5 1 1 15867
0 15869 7 2 2 24989 23275
0 15870 7 3 2 25315 37376
0 15871 7 1 2 37378 37069
0 15872 5 1 1 15871
0 15873 7 2 2 23482 23586
0 15874 7 4 2 23053 37381
0 15875 7 2 2 36681 37383
0 15876 5 1 1 37387
0 15877 7 1 2 15872 15876
0 15878 5 3 1 15877
0 15879 7 1 2 32429 34663
0 15880 5 1 1 15879
0 15881 7 1 2 32584 37288
0 15882 5 1 1 15881
0 15883 7 2 2 15880 15882
0 15884 5 1 1 37392
0 15885 7 3 2 26191 35213
0 15886 7 2 2 30673 37394
0 15887 7 1 2 15884 37397
0 15888 5 1 1 15887
0 15889 7 1 2 35233 36064
0 15890 5 1 1 15889
0 15891 7 1 2 31510 37172
0 15892 5 1 1 15891
0 15893 7 2 2 15890 15892
0 15894 7 1 2 22497 37399
0 15895 5 1 1 15894
0 15896 7 3 2 25814 31234
0 15897 7 1 2 33514 37401
0 15898 5 2 1 15897
0 15899 7 1 2 37404 37304
0 15900 5 1 1 15899
0 15901 7 1 2 25713 15900
0 15902 5 2 1 15901
0 15903 7 1 2 24467 37406
0 15904 5 1 1 15903
0 15905 7 1 2 24605 15904
0 15906 7 1 2 15895 15905
0 15907 5 1 1 15906
0 15908 7 1 2 36056 37170
0 15909 5 1 1 15908
0 15910 7 1 2 24697 15909
0 15911 7 1 2 15907 15910
0 15912 5 1 1 15911
0 15913 7 2 2 30238 28384
0 15914 5 2 1 37408
0 15915 7 1 2 35722 30764
0 15916 5 1 1 15915
0 15917 7 1 2 37410 15916
0 15918 5 1 1 15917
0 15919 7 1 2 37291 15918
0 15920 5 1 1 15919
0 15921 7 1 2 22752 15920
0 15922 5 1 1 15921
0 15923 7 1 2 25085 15922
0 15924 7 1 2 15912 15923
0 15925 5 1 1 15924
0 15926 7 1 2 15888 15925
0 15927 5 1 1 15926
0 15928 7 1 2 35055 15927
0 15929 5 1 1 15928
0 15930 7 1 2 22855 37132
0 15931 5 2 1 15930
0 15932 7 1 2 35029 37189
0 15933 5 1 1 15932
0 15934 7 1 2 37412 15933
0 15935 5 1 1 15934
0 15936 7 1 2 32585 37292
0 15937 7 1 2 15935 15936
0 15938 5 1 1 15937
0 15939 7 1 2 15929 15938
0 15940 5 1 1 15939
0 15941 7 1 2 37389 15940
0 15942 5 1 1 15941
0 15943 7 1 2 25133 15942
0 15944 7 1 2 15868 15943
0 15945 7 1 2 15709 15944
0 15946 7 1 2 15232 15945
0 15947 5 1 1 15946
0 15948 7 4 2 25443 37359
0 15949 7 1 2 35340 37414
0 15950 5 1 1 15949
0 15951 7 1 2 123 14128
0 15952 5 1 1 15951
0 15953 7 1 2 33030 37384
0 15954 7 1 2 15952 15953
0 15955 5 1 1 15954
0 15956 7 1 2 15950 15955
0 15957 5 1 1 15956
0 15958 7 1 2 23555 15957
0 15959 5 1 1 15958
0 15960 7 2 2 37070 36851
0 15961 7 1 2 37379 37418
0 15962 5 1 1 15961
0 15963 7 1 2 15959 15962
0 15964 5 1 1 15963
0 15965 7 1 2 22647 15964
0 15966 5 1 1 15965
0 15967 7 2 2 28808 36700
0 15968 7 1 2 35426 37420
0 15969 5 1 1 15968
0 15970 7 2 2 25383 37415
0 15971 7 1 2 23360 37422
0 15972 5 1 1 15971
0 15973 7 1 2 15969 15972
0 15974 5 1 1 15973
0 15975 7 1 2 23556 30653
0 15976 7 1 2 15974 15975
0 15977 5 1 1 15976
0 15978 7 1 2 15966 15977
0 15979 5 1 1 15978
0 15980 7 1 2 23821 15979
0 15981 5 1 1 15980
0 15982 7 1 2 35304 34672
0 15983 7 1 2 37006 15982
0 15984 7 1 2 36779 15983
0 15985 5 1 1 15984
0 15986 7 1 2 15981 15985
0 15987 5 1 1 15986
0 15988 7 1 2 23942 15987
0 15989 5 1 1 15988
0 15990 7 2 2 28708 36780
0 15991 7 1 2 37374 36895
0 15992 7 1 2 37424 15991
0 15993 5 1 1 15992
0 15994 7 1 2 15989 15993
0 15995 5 1 1 15994
0 15996 7 1 2 24468 15995
0 15997 5 1 1 15996
0 15998 7 1 2 37419 36771
0 15999 5 1 1 15998
0 16000 7 1 2 24606 28556
0 16001 7 1 2 37421 16000
0 16002 5 1 1 16001
0 16003 7 1 2 22648 35422
0 16004 7 1 2 37002 16003
0 16005 5 1 1 16004
0 16006 7 1 2 16002 16005
0 16007 5 1 1 16006
0 16008 7 1 2 23557 16007
0 16009 5 1 1 16008
0 16010 7 1 2 15999 16009
0 16011 5 1 1 16010
0 16012 7 1 2 25316 16011
0 16013 5 1 1 16012
0 16014 7 1 2 35381 37423
0 16015 5 1 1 16014
0 16016 7 1 2 16013 16015
0 16017 5 1 1 16016
0 16018 7 1 2 27923 28444
0 16019 7 1 2 16017 16018
0 16020 5 1 1 16019
0 16021 7 1 2 15997 16020
0 16022 5 1 1 16021
0 16023 7 1 2 32586 16022
0 16024 5 1 1 16023
0 16025 7 1 2 33875 26652
0 16026 5 1 1 16025
0 16027 7 2 2 33031 36628
0 16028 7 1 2 37426 36852
0 16029 5 1 1 16028
0 16030 7 1 2 16026 16029
0 16031 5 1 1 16030
0 16032 7 1 2 37385 16031
0 16033 5 1 1 16032
0 16034 7 2 2 32112 27979
0 16035 7 1 2 31325 37428
0 16036 7 1 2 37360 16035
0 16037 5 1 1 16036
0 16038 7 1 2 16033 16037
0 16039 5 1 1 16038
0 16040 7 1 2 23558 16039
0 16041 5 1 1 16040
0 16042 7 1 2 28011 29038
0 16043 7 1 2 33483 16042
0 16044 7 1 2 26520 28676
0 16045 7 1 2 27980 16044
0 16046 7 1 2 16043 16045
0 16047 5 1 1 16046
0 16048 7 1 2 16041 16047
0 16049 5 1 1 16048
0 16050 7 1 2 25916 16049
0 16051 5 1 1 16050
0 16052 7 1 2 28716 36723
0 16053 5 1 1 16052
0 16054 7 1 2 23430 37416
0 16055 5 1 1 16054
0 16056 7 1 2 16053 16055
0 16057 5 2 1 16056
0 16058 7 1 2 34044 33493
0 16059 7 1 2 37430 16058
0 16060 5 1 1 16059
0 16061 7 1 2 16051 16060
0 16062 5 1 1 16061
0 16063 7 1 2 24607 16062
0 16064 5 1 1 16063
0 16065 7 1 2 30838 31166
0 16066 5 1 1 16065
0 16067 7 1 2 31581 34295
0 16068 5 1 1 16067
0 16069 7 1 2 16066 16068
0 16070 5 1 1 16069
0 16071 7 1 2 24469 16070
0 16072 5 1 1 16071
0 16073 7 1 2 30839 31246
0 16074 5 1 1 16073
0 16075 7 1 2 16072 16074
0 16076 5 1 1 16075
0 16077 7 1 2 37417 16076
0 16078 5 1 1 16077
0 16079 7 1 2 31017 31251
0 16080 5 1 1 16079
0 16081 7 2 2 24470 30075
0 16082 7 1 2 27761 37432
0 16083 5 1 1 16082
0 16084 7 1 2 16080 16083
0 16085 5 1 1 16084
0 16086 7 1 2 26653 37386
0 16087 7 1 2 16085 16086
0 16088 5 1 1 16087
0 16089 7 1 2 16078 16088
0 16090 5 1 1 16089
0 16091 7 1 2 30614 16090
0 16092 5 1 1 16091
0 16093 7 1 2 16064 16092
0 16094 5 1 1 16093
0 16095 7 1 2 24037 16094
0 16096 5 1 1 16095
0 16097 7 1 2 30791 33447
0 16098 7 1 2 29253 16097
0 16099 7 1 2 37431 16098
0 16100 5 1 1 16099
0 16101 7 1 2 16096 16100
0 16102 5 1 1 16101
0 16103 7 1 2 23822 16102
0 16104 5 1 1 16103
0 16105 7 1 2 16024 16104
0 16106 5 1 1 16105
0 16107 7 1 2 33147 16106
0 16108 5 1 1 16107
0 16109 7 2 2 28327 26627
0 16110 5 1 1 37434
0 16111 7 1 2 28943 37435
0 16112 5 1 1 16111
0 16113 7 1 2 29254 37346
0 16114 5 1 1 16113
0 16115 7 1 2 16112 16114
0 16116 5 1 1 16115
0 16117 7 1 2 24300 16116
0 16118 5 1 1 16117
0 16119 7 2 2 28311 33722
0 16120 5 1 1 37436
0 16121 7 1 2 28944 26675
0 16122 7 1 2 37437 16121
0 16123 5 1 1 16122
0 16124 7 1 2 16118 16123
0 16125 5 1 1 16124
0 16126 7 1 2 30104 16125
0 16127 5 1 1 16126
0 16128 7 1 2 30050 28424
0 16129 7 5 2 23643 25815
0 16130 7 2 2 32382 37438
0 16131 7 1 2 30150 37443
0 16132 7 1 2 16128 16131
0 16133 5 1 1 16132
0 16134 7 1 2 16127 16133
0 16135 5 1 1 16134
0 16136 7 1 2 29008 16135
0 16137 5 1 1 16136
0 16138 7 1 2 31364 37250
0 16139 5 1 1 16138
0 16140 7 3 2 23823 36763
0 16141 7 1 2 35895 37445
0 16142 5 1 1 16141
0 16143 7 1 2 16139 16142
0 16144 5 1 1 16143
0 16145 7 1 2 23943 16144
0 16146 5 1 1 16145
0 16147 7 1 2 25917 31569
0 16148 7 1 2 37251 16147
0 16149 5 1 1 16148
0 16150 7 1 2 16146 16149
0 16151 5 1 1 16150
0 16152 7 1 2 35709 16151
0 16153 5 1 1 16152
0 16154 7 3 2 23559 37269
0 16155 7 2 2 24122 37448
0 16156 5 1 1 37451
0 16157 7 1 2 35900 37452
0 16158 7 1 2 31305 16157
0 16159 5 1 1 16158
0 16160 7 1 2 16153 16159
0 16161 5 1 1 16160
0 16162 7 1 2 28945 16161
0 16163 5 1 1 16162
0 16164 7 5 2 35710 37446
0 16165 7 1 2 23944 28958
0 16166 7 1 2 31365 16165
0 16167 7 1 2 37453 16166
0 16168 5 1 1 16167
0 16169 7 1 2 16163 16168
0 16170 5 1 1 16169
0 16171 7 1 2 28222 16170
0 16172 5 1 1 16171
0 16173 7 1 2 16137 16172
0 16174 5 1 1 16173
0 16175 7 1 2 27088 16174
0 16176 5 1 1 16175
0 16177 7 3 2 24123 36764
0 16178 7 3 2 36015 37458
0 16179 7 2 2 27924 37461
0 16180 7 3 2 23945 34028
0 16181 5 1 1 37466
0 16182 7 1 2 37464 37467
0 16183 5 1 1 16182
0 16184 7 2 2 29521 26688
0 16185 7 1 2 32194 37469
0 16186 5 1 1 16185
0 16187 7 2 2 33396 35114
0 16188 7 1 2 33448 36905
0 16189 7 1 2 37471 16188
0 16190 5 1 1 16189
0 16191 7 1 2 16186 16190
0 16192 5 2 1 16191
0 16193 7 1 2 23431 37473
0 16194 5 1 1 16193
0 16195 7 1 2 29877 37449
0 16196 5 1 1 16195
0 16197 7 1 2 36457 28692
0 16198 5 1 1 16197
0 16199 7 1 2 16196 16198
0 16200 5 1 1 16199
0 16201 7 1 2 36422 16200
0 16202 5 1 1 16201
0 16203 7 1 2 16194 16202
0 16204 5 1 1 16203
0 16205 7 1 2 23141 16204
0 16206 5 1 1 16205
0 16207 7 1 2 30211 33723
0 16208 7 2 2 36948 16207
0 16209 7 1 2 30960 37475
0 16210 5 1 1 16209
0 16211 7 1 2 16206 16210
0 16212 5 1 1 16211
0 16213 7 1 2 25228 16212
0 16214 5 1 1 16213
0 16215 7 1 2 23276 32180
0 16216 7 1 2 37462 16215
0 16217 5 1 1 16216
0 16218 7 1 2 24698 16217
0 16219 7 1 2 16214 16218
0 16220 5 1 1 16219
0 16221 7 1 2 23142 37474
0 16222 5 1 1 16221
0 16223 7 1 2 29902 37476
0 16224 5 1 1 16223
0 16225 7 1 2 16222 16224
0 16226 5 1 1 16225
0 16227 7 1 2 25229 16226
0 16228 5 1 1 16227
0 16229 7 1 2 30740 28455
0 16230 7 1 2 37459 16229
0 16231 5 1 1 16230
0 16232 7 1 2 16228 16231
0 16233 5 1 1 16232
0 16234 7 1 2 25384 16233
0 16235 5 1 1 16234
0 16236 7 1 2 27155 30557
0 16237 7 1 2 35917 16236
0 16238 7 1 2 37347 16237
0 16239 5 1 1 16238
0 16240 7 1 2 22753 16239
0 16241 7 1 2 16235 16240
0 16242 5 1 1 16241
0 16243 7 1 2 24471 16242
0 16244 7 1 2 16220 16243
0 16245 5 1 1 16244
0 16246 7 1 2 16183 16245
0 16247 5 1 1 16246
0 16248 7 1 2 28164 16247
0 16249 5 1 1 16248
0 16250 7 2 2 28245 30076
0 16251 5 1 1 37477
0 16252 7 1 2 22754 29205
0 16253 5 1 1 16252
0 16254 7 1 2 16251 16253
0 16255 5 1 1 16254
0 16256 7 1 2 37463 16255
0 16257 5 1 1 16256
0 16258 7 1 2 22755 37470
0 16259 5 1 1 16258
0 16260 7 1 2 29305 37450
0 16261 5 1 1 16260
0 16262 7 1 2 16259 16261
0 16263 5 1 1 16262
0 16264 7 1 2 23143 16263
0 16265 5 1 1 16264
0 16266 7 1 2 30004 37255
0 16267 5 1 1 16266
0 16268 7 1 2 16265 16267
0 16269 5 1 1 16268
0 16270 7 1 2 28275 28312
0 16271 7 1 2 16269 16270
0 16272 5 1 1 16271
0 16273 7 1 2 16257 16272
0 16274 5 1 1 16273
0 16275 7 1 2 24472 16274
0 16276 5 1 1 16275
0 16277 7 1 2 35548 37465
0 16278 5 1 1 16277
0 16279 7 1 2 16276 16278
0 16280 5 1 1 16279
0 16281 7 1 2 27001 16280
0 16282 5 1 1 16281
0 16283 7 4 2 25637 23824
0 16284 7 1 2 26379 26672
0 16285 7 1 2 37479 16284
0 16286 7 1 2 30105 16285
0 16287 7 1 2 29255 16286
0 16288 5 1 1 16287
0 16289 7 1 2 16282 16288
0 16290 7 1 2 16249 16289
0 16291 5 1 1 16290
0 16292 7 1 2 29009 16291
0 16293 5 1 1 16292
0 16294 7 1 2 32401 29200
0 16295 5 1 1 16294
0 16296 7 1 2 16156 16295
0 16297 5 1 1 16296
0 16298 7 1 2 23144 16297
0 16299 5 1 1 16298
0 16300 7 1 2 29808 37277
0 16301 5 1 1 16300
0 16302 7 1 2 16299 16301
0 16303 5 1 1 16302
0 16304 7 1 2 28276 16303
0 16305 5 1 1 16304
0 16306 7 1 2 23277 37454
0 16307 5 1 1 16306
0 16308 7 1 2 16305 16307
0 16309 5 2 1 16308
0 16310 7 1 2 28313 37483
0 16311 5 1 1 16310
0 16312 7 1 2 29215 37455
0 16313 5 1 1 16312
0 16314 7 1 2 16311 16313
0 16315 5 1 1 16314
0 16316 7 1 2 24473 16315
0 16317 5 1 1 16316
0 16318 7 1 2 29240 37456
0 16319 5 1 1 16318
0 16320 7 1 2 16317 16319
0 16321 5 1 1 16320
0 16322 7 1 2 27002 16321
0 16323 5 1 1 16322
0 16324 7 1 2 24474 37484
0 16325 5 1 1 16324
0 16326 7 1 2 27925 37457
0 16327 5 1 1 16326
0 16328 7 1 2 16325 16327
0 16329 5 1 1 16328
0 16330 7 1 2 31771 16329
0 16331 5 1 1 16330
0 16332 7 1 2 36016 33703
0 16333 7 1 2 31140 16332
0 16334 7 1 2 37278 16333
0 16335 5 1 1 16334
0 16336 7 1 2 16331 16335
0 16337 5 1 1 16336
0 16338 7 1 2 28165 16337
0 16339 5 1 1 16338
0 16340 7 1 2 16323 16339
0 16341 5 1 1 16340
0 16342 7 1 2 27136 16341
0 16343 5 1 1 16342
0 16344 7 1 2 34715 36949
0 16345 5 1 1 16344
0 16346 7 1 2 26380 26663
0 16347 5 1 1 16346
0 16348 7 1 2 16345 16347
0 16349 5 1 1 16348
0 16350 7 1 2 36017 30773
0 16351 7 1 2 16349 16350
0 16352 7 1 2 35370 16351
0 16353 5 1 1 16352
0 16354 7 1 2 16343 16353
0 16355 7 1 2 16293 16354
0 16356 7 1 2 16176 16355
0 16357 5 1 1 16356
0 16358 7 1 2 36820 16357
0 16359 5 1 1 16358
0 16360 7 1 2 32902 35601
0 16361 5 1 1 16360
0 16362 7 1 2 23361 31427
0 16363 7 1 2 33862 16362
0 16364 7 1 2 34552 16363
0 16365 5 1 1 16364
0 16366 7 1 2 16361 16365
0 16367 5 1 1 16366
0 16368 7 1 2 25918 16367
0 16369 5 1 1 16368
0 16370 7 1 2 28246 27745
0 16371 7 1 2 35965 16370
0 16372 5 1 1 16371
0 16373 7 1 2 16369 16372
0 16374 5 1 1 16373
0 16375 7 1 2 36932 16374
0 16376 5 1 1 16375
0 16377 7 1 2 34871 36906
0 16378 7 1 2 35967 16377
0 16379 7 2 2 36181 31547
0 16380 7 1 2 16378 37485
0 16381 5 1 1 16380
0 16382 7 1 2 16376 16381
0 16383 5 1 1 16382
0 16384 7 1 2 25086 16383
0 16385 5 1 1 16384
0 16386 7 1 2 28012 34156
0 16387 7 1 2 31683 16386
0 16388 7 1 2 26646 16387
0 16389 5 1 1 16388
0 16390 7 1 2 35214 37486
0 16391 5 1 1 16390
0 16392 7 1 2 16389 16391
0 16393 5 1 1 16392
0 16394 7 1 2 26102 16393
0 16395 5 1 1 16394
0 16396 7 1 2 31684 26416
0 16397 5 1 1 16396
0 16398 7 1 2 11031 16397
0 16399 5 1 1 16398
0 16400 7 1 2 35138 16399
0 16401 5 1 1 16400
0 16402 7 1 2 16395 16401
0 16403 5 1 1 16402
0 16404 7 1 2 23432 16403
0 16405 5 1 1 16404
0 16406 7 1 2 26851 35632
0 16407 5 1 1 16406
0 16408 7 1 2 32919 26647
0 16409 5 1 1 16408
0 16410 7 1 2 16407 16409
0 16411 5 1 1 16410
0 16412 7 2 2 33791 16411
0 16413 7 1 2 31088 37487
0 16414 5 1 1 16413
0 16415 7 1 2 16405 16414
0 16416 5 1 1 16415
0 16417 7 1 2 23362 16416
0 16418 5 1 1 16417
0 16419 7 2 2 29762 35628
0 16420 7 1 2 26358 30588
0 16421 7 1 2 37489 16420
0 16422 5 1 1 16421
0 16423 7 1 2 27835 26648
0 16424 7 1 2 32879 16423
0 16425 5 1 1 16424
0 16426 7 1 2 16422 16425
0 16427 5 1 1 16426
0 16428 7 1 2 22649 16427
0 16429 5 1 1 16428
0 16430 7 1 2 27399 35629
0 16431 7 1 2 30301 16430
0 16432 7 1 2 28038 16431
0 16433 5 1 1 16432
0 16434 7 1 2 16429 16433
0 16435 5 1 1 16434
0 16436 7 1 2 32113 16435
0 16437 5 1 1 16436
0 16438 7 1 2 27854 27757
0 16439 7 1 2 37488 16438
0 16440 5 1 1 16439
0 16441 7 1 2 16437 16440
0 16442 7 1 2 16418 16441
0 16443 5 1 1 16442
0 16444 7 1 2 23587 28557
0 16445 7 1 2 16443 16444
0 16446 5 1 1 16445
0 16447 7 1 2 16385 16446
0 16448 5 1 1 16447
0 16449 7 1 2 30524 16448
0 16450 5 1 1 16449
0 16451 7 2 2 32516 32618
0 16452 7 1 2 30765 37491
0 16453 5 1 1 16452
0 16454 7 1 2 23560 26639
0 16455 7 1 2 34272 16454
0 16456 5 1 1 16455
0 16457 7 1 2 16453 16456
0 16458 5 1 1 16457
0 16459 7 1 2 25087 16458
0 16460 5 1 1 16459
0 16461 7 1 2 37492 36746
0 16462 5 1 1 16461
0 16463 7 1 2 16460 16462
0 16464 5 1 1 16463
0 16465 7 1 2 26014 16464
0 16466 5 1 1 16465
0 16467 7 1 2 35995 37102
0 16468 5 1 1 16467
0 16469 7 1 2 16466 16468
0 16470 5 1 1 16469
0 16471 7 1 2 25385 16470
0 16472 5 1 1 16471
0 16473 7 1 2 32637 33252
0 16474 7 1 2 35666 16473
0 16475 7 1 2 37073 16474
0 16476 5 1 1 16475
0 16477 7 1 2 16472 16476
0 16478 5 1 1 16477
0 16479 7 1 2 25919 16478
0 16480 5 1 1 16479
0 16481 7 1 2 26974 34857
0 16482 7 1 2 37103 16481
0 16483 5 1 1 16482
0 16484 7 1 2 16480 16483
0 16485 5 1 1 16484
0 16486 7 1 2 24699 16485
0 16487 5 1 1 16486
0 16488 7 1 2 23946 35963
0 16489 5 1 1 16488
0 16490 7 1 2 29903 37246
0 16491 5 1 1 16490
0 16492 7 1 2 16489 16491
0 16493 5 1 1 16492
0 16494 7 1 2 32638 33628
0 16495 7 1 2 26640 16494
0 16496 7 1 2 16493 16495
0 16497 5 1 1 16496
0 16498 7 1 2 16487 16497
0 16499 5 1 1 16498
0 16500 7 1 2 33563 16499
0 16501 5 1 1 16500
0 16502 7 1 2 10922 8075
0 16503 5 2 1 16502
0 16504 7 1 2 27003 37493
0 16505 5 1 1 16504
0 16506 7 2 2 32765 30792
0 16507 5 1 1 37495
0 16508 7 1 2 27089 37496
0 16509 5 1 1 16508
0 16510 7 1 2 32791 32825
0 16511 5 1 1 16510
0 16512 7 1 2 16509 16511
0 16513 7 1 2 16505 16512
0 16514 5 1 1 16513
0 16515 7 1 2 26649 16514
0 16516 5 1 1 16515
0 16517 7 1 2 27341 33389
0 16518 7 1 2 37490 16517
0 16519 5 1 1 16518
0 16520 7 1 2 16516 16519
0 16521 5 1 1 16520
0 16522 7 2 2 32716 34067
0 16523 5 1 1 37497
0 16524 7 1 2 23145 37498
0 16525 7 1 2 16521 16524
0 16526 5 1 1 16525
0 16527 7 1 2 28314 16526
0 16528 7 1 2 16501 16527
0 16529 5 1 1 16528
0 16530 7 1 2 29878 33378
0 16531 5 1 1 16530
0 16532 7 1 2 24787 30961
0 16533 5 1 1 16532
0 16534 7 1 2 16531 16533
0 16535 5 1 1 16534
0 16536 7 1 2 24700 16535
0 16537 5 1 1 16536
0 16538 7 1 2 27052 35136
0 16539 5 1 1 16538
0 16540 7 1 2 16537 16539
0 16541 5 2 1 16540
0 16542 7 1 2 23483 15803
0 16543 5 1 1 16542
0 16544 7 1 2 25444 13960
0 16545 5 1 1 16544
0 16546 7 1 2 30907 16545
0 16547 7 1 2 16543 16546
0 16548 7 1 2 37499 16547
0 16549 5 1 1 16548
0 16550 7 1 2 28323 16549
0 16551 5 1 1 16550
0 16552 7 1 2 28252 27981
0 16553 7 1 2 16551 16552
0 16554 7 1 2 16529 16553
0 16555 5 1 1 16554
0 16556 7 1 2 16450 16555
0 16557 5 1 1 16556
0 16558 7 1 2 23825 16557
0 16559 5 1 1 16558
0 16560 7 1 2 16359 16559
0 16561 7 1 2 16108 16560
0 16562 5 1 1 16561
0 16563 7 1 2 37114 16562
0 16564 5 1 1 16563
0 16565 7 3 2 31123 29284
0 16566 7 3 2 27787 33571
0 16567 7 1 2 24334 26865
0 16568 7 1 2 37504 16567
0 16569 7 1 2 37501 16568
0 16570 5 1 1 16569
0 16571 7 1 2 24911 34091
0 16572 5 1 1 16571
0 16573 7 1 2 34268 16572
0 16574 5 2 1 16573
0 16575 7 1 2 33164 31884
0 16576 7 1 2 31347 16575
0 16577 7 1 2 37507 16576
0 16578 5 1 1 16577
0 16579 7 1 2 16570 16578
0 16580 5 1 1 16579
0 16581 7 1 2 25638 16580
0 16582 5 1 1 16581
0 16583 7 1 2 25586 26192
0 16584 7 4 2 28896 16583
0 16585 5 1 1 37509
0 16586 7 1 2 31141 37510
0 16587 5 1 1 16586
0 16588 7 2 2 33085 36701
0 16589 7 1 2 23278 31047
0 16590 7 1 2 37513 16589
0 16591 5 1 1 16590
0 16592 7 1 2 16587 16591
0 16593 5 1 1 16592
0 16594 7 1 2 30849 16593
0 16595 5 1 1 16594
0 16596 7 1 2 16582 16595
0 16597 5 1 1 16596
0 16598 7 1 2 24475 16597
0 16599 5 1 1 16598
0 16600 7 1 2 33572 31939
0 16601 5 1 1 16600
0 16602 7 1 2 35291 36702
0 16603 5 1 1 16602
0 16604 7 1 2 16601 16603
0 16605 5 2 1 16604
0 16606 7 1 2 27721 34207
0 16607 7 1 2 33086 16606
0 16608 7 1 2 37515 16607
0 16609 5 1 1 16608
0 16610 7 1 2 16599 16609
0 16611 5 1 1 16610
0 16612 7 1 2 25505 16611
0 16613 5 1 1 16612
0 16614 7 2 2 28566 29619
0 16615 7 1 2 30850 33573
0 16616 7 2 2 37517 16615
0 16617 7 1 2 34962 31982
0 16618 7 1 2 27982 16617
0 16619 7 1 2 37519 16618
0 16620 5 1 1 16619
0 16621 7 1 2 16613 16620
0 16622 5 1 1 16621
0 16623 7 1 2 29010 16622
0 16624 5 1 1 16623
0 16625 7 2 2 27983 26440
0 16626 7 1 2 35094 37502
0 16627 7 1 2 37521 16626
0 16628 5 1 1 16627
0 16629 7 4 2 29763 28946
0 16630 7 1 2 35757 27638
0 16631 7 1 2 37523 16630
0 16632 7 1 2 37220 16631
0 16633 5 1 1 16632
0 16634 7 1 2 16628 16633
0 16635 5 1 1 16634
0 16636 7 1 2 25506 16635
0 16637 5 1 1 16636
0 16638 7 4 2 23146 33574
0 16639 7 1 2 30271 37527
0 16640 5 1 1 16639
0 16641 7 1 2 34081 32028
0 16642 5 1 1 16641
0 16643 7 1 2 16640 16642
0 16644 5 1 1 16643
0 16645 7 1 2 26271 16644
0 16646 5 1 1 16645
0 16647 7 1 2 22977 36828
0 16648 5 1 1 16647
0 16649 7 1 2 16646 16648
0 16650 5 1 1 16649
0 16651 7 1 2 26193 16650
0 16652 5 1 1 16651
0 16653 7 2 2 23588 29817
0 16654 5 1 1 37531
0 16655 7 1 2 35934 37532
0 16656 5 1 1 16655
0 16657 7 1 2 16652 16656
0 16658 5 1 1 16657
0 16659 7 1 2 23561 37524
0 16660 7 1 2 16658 16659
0 16661 5 1 1 16660
0 16662 7 1 2 16637 16661
0 16663 5 2 1 16662
0 16664 7 1 2 28737 37533
0 16665 5 1 1 16664
0 16666 7 1 2 16624 16665
0 16667 5 1 1 16666
0 16668 7 1 2 24124 16667
0 16669 5 1 1 16668
0 16670 7 1 2 29118 37224
0 16671 5 1 1 16670
0 16672 7 1 2 34592 31058
0 16673 5 1 1 16672
0 16674 7 1 2 16671 16673
0 16675 5 1 1 16674
0 16676 7 1 2 37525 37227
0 16677 7 2 2 16675 16676
0 16678 7 1 2 28738 37535
0 16679 5 1 1 16678
0 16680 7 1 2 16669 16679
0 16681 5 1 1 16680
0 16682 7 1 2 32183 16681
0 16683 5 1 1 16682
0 16684 7 1 2 35968 37514
0 16685 5 1 1 16684
0 16686 7 1 2 29764 28677
0 16687 7 1 2 37511 16686
0 16688 5 1 1 16687
0 16689 7 1 2 16685 16688
0 16690 5 1 1 16689
0 16691 7 1 2 23147 16690
0 16692 5 1 1 16691
0 16693 7 1 2 26015 31574
0 16694 7 1 2 34572 16693
0 16695 7 1 2 36691 16694
0 16696 5 1 1 16695
0 16697 7 1 2 16692 16696
0 16698 5 1 1 16697
0 16699 7 1 2 24912 16698
0 16700 5 1 1 16699
0 16701 7 1 2 24301 36435
0 16702 7 1 2 24990 25317
0 16703 7 2 2 26866 16702
0 16704 7 1 2 36223 37537
0 16705 7 1 2 16701 16704
0 16706 5 1 1 16705
0 16707 7 1 2 16700 16706
0 16708 5 1 1 16707
0 16709 7 1 2 29011 16708
0 16710 5 1 1 16709
0 16711 7 1 2 35865 36912
0 16712 7 1 2 35097 16711
0 16713 5 1 1 16712
0 16714 7 1 2 16710 16713
0 16715 5 1 1 16714
0 16716 7 1 2 25507 16715
0 16717 5 1 1 16716
0 16718 7 4 2 24788 23589
0 16719 7 1 2 35292 31983
0 16720 7 1 2 37539 16719
0 16721 7 1 2 32688 37518
0 16722 7 1 2 16720 16721
0 16723 5 1 1 16722
0 16724 7 1 2 16717 16723
0 16725 5 1 1 16724
0 16726 7 1 2 27984 16725
0 16727 5 1 1 16726
0 16728 7 1 2 25508 32394
0 16729 7 1 2 36436 16728
0 16730 7 1 2 37503 16729
0 16731 7 1 2 33046 16730
0 16732 5 1 1 16731
0 16733 7 1 2 23562 37512
0 16734 5 1 1 16733
0 16735 7 1 2 34068 91
0 16736 7 1 2 28656 16735
0 16737 7 1 2 2889 16736
0 16738 5 1 1 16737
0 16739 7 1 2 16734 16738
0 16740 5 1 1 16739
0 16741 7 1 2 23148 16740
0 16742 5 1 1 16741
0 16743 7 1 2 29354 36866
0 16744 5 1 1 16743
0 16745 7 1 2 16742 16744
0 16746 5 1 1 16745
0 16747 7 1 2 26016 33792
0 16748 7 1 2 36235 16747
0 16749 7 1 2 31862 16748
0 16750 7 1 2 16746 16749
0 16751 5 1 1 16750
0 16752 7 1 2 16732 16751
0 16753 7 1 2 16727 16752
0 16754 5 1 1 16753
0 16755 7 1 2 24125 16754
0 16756 5 1 1 16755
0 16757 7 1 2 22978 37232
0 16758 5 1 1 16757
0 16759 7 1 2 25509 16758
0 16760 5 1 1 16759
0 16761 7 1 2 16585 14143
0 16762 5 1 1 16761
0 16763 7 1 2 27674 16762
0 16764 5 1 1 16763
0 16765 7 1 2 29064 16764
0 16766 7 1 2 14293 16765
0 16767 5 1 1 16766
0 16768 7 1 2 23149 37212
0 16769 5 1 1 16768
0 16770 7 1 2 24913 37230
0 16771 7 1 2 16769 16770
0 16772 5 1 1 16771
0 16773 7 1 2 24476 29765
0 16774 7 1 2 16772 16773
0 16775 7 1 2 16767 16774
0 16776 7 1 2 16760 16775
0 16777 5 1 1 16776
0 16778 7 1 2 25510 24302
0 16779 7 1 2 29731 16778
0 16780 7 1 2 35095 16779
0 16781 7 1 2 33515 16780
0 16782 5 1 1 16781
0 16783 7 1 2 16777 16782
0 16784 5 1 1 16783
0 16785 7 1 2 33038 16784
0 16786 5 1 1 16785
0 16787 7 5 2 26689 31075
0 16788 7 2 2 35305 36236
0 16789 5 1 1 37548
0 16790 7 2 2 29766 37549
0 16791 7 1 2 26103 37550
0 16792 5 1 1 16791
0 16793 7 1 2 35045 29139
0 16794 7 1 2 34273 16793
0 16795 5 1 1 16794
0 16796 7 1 2 16792 16795
0 16797 5 1 1 16796
0 16798 7 1 2 37543 16797
0 16799 5 1 1 16798
0 16800 7 1 2 37551 37047
0 16801 5 1 1 16800
0 16802 7 1 2 16799 16801
0 16803 5 1 1 16802
0 16804 7 1 2 37528 16803
0 16805 5 1 1 16804
0 16806 7 1 2 26610 37540
0 16807 7 1 2 35572 16806
0 16808 7 1 2 35306 37228
0 16809 7 1 2 16807 16808
0 16810 5 1 1 16809
0 16811 7 1 2 16805 16810
0 16812 5 1 1 16811
0 16813 7 1 2 29119 16812
0 16814 5 1 1 16813
0 16815 7 1 2 36237 29620
0 16816 7 1 2 29932 16815
0 16817 7 2 2 24212 35418
0 16818 7 1 2 33590 37538
0 16819 7 1 2 37552 16818
0 16820 7 1 2 16816 16819
0 16821 5 1 1 16820
0 16822 7 1 2 16814 16821
0 16823 7 1 2 16786 16822
0 16824 7 1 2 16756 16823
0 16825 5 1 1 16824
0 16826 7 1 2 23826 16825
0 16827 5 1 1 16826
0 16828 7 1 2 24477 37390
0 16829 5 1 1 16828
0 16830 7 1 2 30012 37375
0 16831 5 1 1 16830
0 16832 7 1 2 16829 16831
0 16833 5 1 1 16832
0 16834 7 2 2 25639 31076
0 16835 5 2 1 37554
0 16836 7 1 2 33386 37556
0 16837 7 2 2 37115 16836
0 16838 7 2 2 27240 37558
0 16839 7 2 2 22856 37560
0 16840 5 2 1 37562
0 16841 7 1 2 34635 36988
0 16842 5 1 1 16841
0 16843 7 1 2 25920 32363
0 16844 7 2 2 34586 16843
0 16845 5 1 1 37566
0 16846 7 1 2 16842 16845
0 16847 5 1 1 16846
0 16848 7 1 2 33253 31235
0 16849 7 1 2 16847 16848
0 16850 5 1 1 16849
0 16851 7 1 2 37564 16850
0 16852 5 1 1 16851
0 16853 7 1 2 16833 16852
0 16854 5 1 1 16853
0 16855 7 1 2 29461 31918
0 16856 7 1 2 29621 16855
0 16857 7 6 2 28678 35419
0 16858 7 1 2 29039 30091
0 16859 7 1 2 37568 16858
0 16860 7 1 2 16856 16859
0 16861 7 1 2 36066 16860
0 16862 5 1 1 16861
0 16863 7 1 2 16854 16862
0 16864 7 1 2 16827 16863
0 16865 5 1 1 16864
0 16866 7 1 2 24701 16865
0 16867 5 1 1 16866
0 16868 7 1 2 16683 16867
0 16869 5 1 1 16868
0 16870 7 1 2 24608 16869
0 16871 5 1 1 16870
0 16872 7 1 2 26726 31124
0 16873 7 2 2 37460 16872
0 16874 7 1 2 31204 37574
0 16875 5 1 1 16874
0 16876 7 1 2 23563 26690
0 16877 5 1 1 16876
0 16878 7 1 2 23150 28432
0 16879 7 1 2 16877 16878
0 16880 5 1 1 16879
0 16881 7 1 2 1542 36976
0 16882 7 2 2 16880 16881
0 16883 7 1 2 27372 33508
0 16884 7 1 2 37576 16883
0 16885 5 1 1 16884
0 16886 7 1 2 16875 16885
0 16887 5 1 1 16886
0 16888 7 1 2 24478 16887
0 16889 5 1 1 16888
0 16890 7 1 2 31760 37575
0 16891 5 1 1 16890
0 16892 7 1 2 16889 16891
0 16893 5 1 1 16892
0 16894 7 1 2 28166 16893
0 16895 5 1 1 16894
0 16896 7 5 2 23564 36765
0 16897 7 1 2 30753 32319
0 16898 5 1 1 16897
0 16899 7 1 2 1972 16898
0 16900 5 3 1 16899
0 16901 7 1 2 37578 37583
0 16902 7 1 2 29256 16901
0 16903 5 1 1 16902
0 16904 7 1 2 16895 16903
0 16905 5 1 1 16904
0 16906 7 1 2 32114 16905
0 16907 5 1 1 16906
0 16908 7 1 2 9824 4160
0 16909 5 5 1 16908
0 16910 7 2 2 31685 37586
0 16911 7 1 2 37579 37591
0 16912 5 1 1 16911
0 16913 7 1 2 27366 26673
0 16914 7 1 2 31575 16913
0 16915 7 1 2 30947 16914
0 16916 5 1 1 16915
0 16917 7 1 2 16912 16916
0 16918 5 1 1 16917
0 16919 7 1 2 33876 16918
0 16920 5 1 1 16919
0 16921 7 1 2 16907 16920
0 16922 5 1 1 16921
0 16923 7 1 2 23827 16922
0 16924 5 1 1 16923
0 16925 7 2 2 28277 37577
0 16926 5 1 1 37593
0 16927 7 1 2 28262 37580
0 16928 5 1 1 16927
0 16929 7 1 2 16926 16928
0 16930 5 1 1 16929
0 16931 7 1 2 33847 16930
0 16932 5 1 1 16931
0 16933 7 1 2 33529 27873
0 16934 7 1 2 37447 16933
0 16935 5 1 1 16934
0 16936 7 1 2 16932 16935
0 16937 5 1 1 16936
0 16938 7 1 2 24479 16937
0 16939 5 1 1 16938
0 16940 7 1 2 33879 37581
0 16941 5 1 1 16940
0 16942 7 1 2 16939 16941
0 16943 5 1 1 16942
0 16944 7 1 2 37587 16943
0 16945 5 1 1 16944
0 16946 7 1 2 31265 29980
0 16947 7 1 2 37526 37043
0 16948 7 1 2 16946 16947
0 16949 5 1 1 16948
0 16950 7 1 2 16945 16949
0 16951 5 1 1 16950
0 16952 7 1 2 32250 16951
0 16953 5 1 1 16952
0 16954 7 2 2 24480 37594
0 16955 7 1 2 32320 30864
0 16956 5 1 1 16955
0 16957 7 2 2 30406 35378
0 16958 5 1 1 37597
0 16959 7 1 2 23947 37598
0 16960 5 1 1 16959
0 16961 7 1 2 16956 16960
0 16962 5 1 1 16961
0 16963 7 1 2 24609 16962
0 16964 5 1 1 16963
0 16965 7 1 2 35454 33516
0 16966 5 1 1 16965
0 16967 7 1 2 16964 16966
0 16968 5 1 1 16967
0 16969 7 1 2 32115 16968
0 16970 5 1 1 16969
0 16971 7 1 2 34514 37592
0 16972 5 1 1 16971
0 16973 7 1 2 16970 16972
0 16974 5 1 1 16973
0 16975 7 1 2 37595 16974
0 16976 5 1 1 16975
0 16977 7 1 2 16953 16976
0 16978 7 1 2 16924 16977
0 16979 5 1 1 16978
0 16980 7 1 2 29012 16979
0 16981 5 1 1 16980
0 16982 7 2 2 24213 30256
0 16983 7 1 2 36907 37599
0 16984 5 1 1 16983
0 16985 7 1 2 35735 31220
0 16986 5 1 1 16985
0 16987 7 1 2 16984 16986
0 16988 5 1 1 16987
0 16989 7 1 2 24303 16988
0 16990 5 1 1 16989
0 16991 7 1 2 27529 28476
0 16992 5 1 1 16991
0 16993 7 1 2 16990 16992
0 16994 5 1 1 16993
0 16995 7 1 2 23565 16994
0 16996 5 1 1 16995
0 16997 7 1 2 35713 36936
0 16998 5 1 1 16997
0 16999 7 1 2 16996 16998
0 17000 5 1 1 16999
0 17001 7 1 2 22650 31412
0 17002 5 1 1 17001
0 17003 7 1 2 3600 17002
0 17004 5 1 1 17003
0 17005 7 1 2 25230 17004
0 17006 5 1 1 17005
0 17007 7 1 2 31135 31570
0 17008 5 1 1 17007
0 17009 7 1 2 17006 17008
0 17010 5 1 1 17009
0 17011 7 1 2 24481 17010
0 17012 5 1 1 17011
0 17013 7 2 2 29587 34398
0 17014 5 1 1 37601
0 17015 7 1 2 24702 37602
0 17016 5 1 1 17015
0 17017 7 1 2 17012 17016
0 17018 5 1 1 17017
0 17019 7 3 2 29767 17018
0 17020 7 1 2 17000 37603
0 17021 5 1 1 17020
0 17022 7 1 2 29216 31907
0 17023 5 1 1 17022
0 17024 7 1 2 6759 17023
0 17025 5 2 1 17024
0 17026 7 1 2 34796 37606
0 17027 5 1 1 17026
0 17028 7 1 2 34799 33895
0 17029 5 1 1 17028
0 17030 7 1 2 17027 17029
0 17031 5 1 1 17030
0 17032 7 1 2 24038 17031
0 17033 5 1 1 17032
0 17034 7 1 2 26975 35347
0 17035 5 1 1 17034
0 17036 7 1 2 17033 17035
0 17037 5 1 1 17036
0 17038 7 1 2 27531 37582
0 17039 7 1 2 17037 17038
0 17040 5 1 1 17039
0 17041 7 1 2 17021 17040
0 17042 5 1 1 17041
0 17043 7 1 2 23828 17042
0 17044 5 1 1 17043
0 17045 7 1 2 35152 27532
0 17046 7 1 2 37596 17045
0 17047 5 1 1 17046
0 17048 7 1 2 17044 17047
0 17049 7 1 2 16981 17048
0 17050 5 1 1 17049
0 17051 7 1 2 36821 17050
0 17052 5 1 1 17051
0 17053 7 4 2 32116 29257
0 17054 7 4 2 29013 36724
0 17055 5 1 1 37612
0 17056 7 1 2 37608 37613
0 17057 5 1 1 17056
0 17058 7 2 2 29212 28346
0 17059 7 1 2 31410 37616
0 17060 5 1 1 17059
0 17061 7 1 2 27985 31418
0 17062 5 1 1 17061
0 17063 7 1 2 17060 17062
0 17064 5 1 1 17063
0 17065 7 1 2 26441 17064
0 17066 5 1 1 17065
0 17067 7 2 2 25640 27342
0 17068 7 1 2 31993 37618
0 17069 7 1 2 33095 17068
0 17070 5 1 1 17069
0 17071 7 1 2 17066 17070
0 17072 5 1 1 17071
0 17073 7 1 2 33524 17072
0 17074 5 1 1 17073
0 17075 7 1 2 17057 17074
0 17076 5 1 1 17075
0 17077 7 1 2 23829 17076
0 17078 5 1 1 17077
0 17079 7 1 2 31236 31338
0 17080 7 1 2 37569 17079
0 17081 7 1 2 34771 17080
0 17082 5 1 1 17081
0 17083 7 1 2 17078 17082
0 17084 5 1 1 17083
0 17085 7 1 2 25511 17084
0 17086 5 1 1 17085
0 17087 7 2 2 29622 37480
0 17088 7 1 2 31922 37620
0 17089 7 1 2 37388 17088
0 17090 5 1 1 17089
0 17091 7 1 2 17086 17090
0 17092 5 1 1 17091
0 17093 7 1 2 37584 17092
0 17094 5 1 1 17093
0 17095 7 1 2 28739 37361
0 17096 5 1 1 17095
0 17097 7 1 2 25386 37614
0 17098 5 1 1 17097
0 17099 7 1 2 17096 17098
0 17100 5 1 1 17099
0 17101 7 1 2 24703 17100
0 17102 5 1 1 17101
0 17103 7 1 2 34792 32019
0 17104 7 1 2 33584 17103
0 17105 5 1 1 17104
0 17106 7 1 2 17102 17105
0 17107 5 1 1 17106
0 17108 7 1 2 34185 17107
0 17109 5 1 1 17108
0 17110 7 1 2 26359 37362
0 17111 5 1 1 17110
0 17112 7 1 2 17055 17111
0 17113 5 1 1 17112
0 17114 7 1 2 17113 37427
0 17115 5 1 1 17114
0 17116 7 1 2 17109 17115
0 17117 5 1 1 17116
0 17118 7 1 2 23830 17117
0 17119 5 1 1 17118
0 17120 7 3 2 24482 35131
0 17121 7 1 2 27812 29588
0 17122 7 1 2 35423 17121
0 17123 7 1 2 37622 17122
0 17124 7 1 2 37402 17123
0 17125 5 1 1 17124
0 17126 7 1 2 17119 17125
0 17127 5 1 1 17126
0 17128 7 1 2 25512 17127
0 17129 5 1 1 17128
0 17130 7 1 2 27390 31331
0 17131 7 1 2 37621 17130
0 17132 7 2 2 23590 32639
0 17133 7 1 2 37625 37623
0 17134 7 1 2 17131 17133
0 17135 5 1 1 17134
0 17136 7 1 2 17129 17135
0 17137 5 1 1 17136
0 17138 7 1 2 31686 17137
0 17139 5 1 1 17138
0 17140 7 1 2 32251 37615
0 17141 5 1 1 17140
0 17142 7 1 2 28881 37363
0 17143 5 1 1 17142
0 17144 7 1 2 17141 17143
0 17145 5 1 1 17144
0 17146 7 1 2 27931 31952
0 17147 5 1 1 17146
0 17148 7 1 2 28959 33855
0 17149 5 1 1 17148
0 17150 7 3 2 17147 17149
0 17151 7 1 2 36018 37627
0 17152 7 1 2 17145 17151
0 17153 5 1 1 17152
0 17154 7 1 2 17139 17153
0 17155 5 1 1 17154
0 17156 7 1 2 37588 17155
0 17157 5 1 1 17156
0 17158 7 2 2 33459 36019
0 17159 7 1 2 24789 28717
0 17160 7 1 2 37380 17159
0 17161 7 1 2 37630 17160
0 17162 5 1 1 17161
0 17163 7 7 2 28679 32619
0 17164 7 1 2 34702 37632
0 17165 5 1 1 17164
0 17166 7 1 2 23831 35969
0 17167 7 1 2 37626 17166
0 17168 5 1 1 17167
0 17169 7 1 2 17165 17168
0 17170 5 1 1 17169
0 17171 7 1 2 25641 31872
0 17172 7 1 2 17170 17171
0 17173 5 1 1 17172
0 17174 7 1 2 17162 17173
0 17175 5 1 1 17174
0 17176 7 1 2 24483 17175
0 17177 5 1 1 17176
0 17178 7 2 2 32292 37631
0 17179 7 1 2 31707 37176
0 17180 7 1 2 37639 17179
0 17181 5 1 1 17180
0 17182 7 1 2 17177 17181
0 17183 5 1 1 17182
0 17184 7 1 2 31687 17183
0 17185 5 1 1 17184
0 17186 7 1 2 32231 34223
0 17187 7 1 2 29014 17186
0 17188 7 1 2 37007 17187
0 17189 7 1 2 37628 17188
0 17190 5 1 1 17189
0 17191 7 1 2 17185 17190
0 17192 5 1 1 17191
0 17193 7 1 2 24335 17192
0 17194 5 1 1 17193
0 17195 7 1 2 27181 27813
0 17196 7 1 2 33472 37481
0 17197 7 1 2 17195 17196
0 17198 7 1 2 29015 17197
0 17199 7 1 2 30323 17198
0 17200 5 1 1 17199
0 17201 7 1 2 17194 17200
0 17202 5 1 1 17201
0 17203 7 1 2 24304 17202
0 17204 5 1 1 17203
0 17205 7 1 2 27986 32355
0 17206 5 1 1 17205
0 17207 7 1 2 33034 28347
0 17208 5 1 1 17207
0 17209 7 1 2 17206 17208
0 17210 5 1 1 17209
0 17211 7 1 2 23054 32368
0 17212 7 1 2 36020 17211
0 17213 7 1 2 36703 17212
0 17214 7 1 2 17210 17213
0 17215 5 1 1 17214
0 17216 7 1 2 17204 17215
0 17217 5 1 1 17216
0 17218 7 1 2 32587 17217
0 17219 5 1 1 17218
0 17220 7 2 2 32807 29258
0 17221 5 1 1 37641
0 17222 7 2 2 31125 30324
0 17223 7 1 2 24704 37643
0 17224 5 1 1 17223
0 17225 7 1 2 17221 17224
0 17226 5 4 1 17225
0 17227 7 1 2 28740 37645
0 17228 5 2 1 17227
0 17229 7 1 2 25231 28843
0 17230 5 1 1 17229
0 17231 7 1 2 24610 33028
0 17232 5 1 1 17231
0 17233 7 1 2 17230 17232
0 17234 5 1 1 17233
0 17235 7 1 2 24484 17234
0 17236 5 1 1 17235
0 17237 7 1 2 17014 17236
0 17238 5 1 1 17237
0 17239 7 2 2 26954 17238
0 17240 7 1 2 22756 37651
0 17241 5 1 1 17240
0 17242 7 1 2 37649 17241
0 17243 5 1 1 17242
0 17244 7 1 2 36725 17243
0 17245 5 1 1 17244
0 17246 7 1 2 30856 30500
0 17247 5 1 1 17246
0 17248 7 1 2 32808 37074
0 17249 5 1 1 17248
0 17250 7 1 2 17247 17249
0 17251 5 1 1 17250
0 17252 7 1 2 29259 17251
0 17253 5 1 1 17252
0 17254 7 1 2 35655 37522
0 17255 5 1 1 17254
0 17256 7 1 2 25921 31841
0 17257 7 1 2 37433 17256
0 17258 5 1 1 17257
0 17259 7 1 2 17255 17258
0 17260 5 1 1 17259
0 17261 7 1 2 37216 17260
0 17262 5 1 1 17261
0 17263 7 1 2 17253 17262
0 17264 5 1 1 17263
0 17265 7 1 2 29016 33525
0 17266 7 1 2 17264 17265
0 17267 5 1 1 17266
0 17268 7 1 2 17245 17267
0 17269 5 1 1 17268
0 17270 7 1 2 36021 17269
0 17271 5 1 1 17270
0 17272 7 1 2 17219 17271
0 17273 5 1 1 17272
0 17274 7 1 2 27533 17273
0 17275 5 1 1 17274
0 17276 7 1 2 31415 37534
0 17277 5 1 1 17276
0 17278 7 1 2 32369 34186
0 17279 7 1 2 34617 17278
0 17280 7 1 2 37516 17279
0 17281 5 1 1 17280
0 17282 7 1 2 32020 37508
0 17283 5 1 1 17282
0 17284 7 1 2 24914 36829
0 17285 5 1 1 17284
0 17286 7 1 2 17283 17285
0 17287 5 1 1 17286
0 17288 7 1 2 28947 36224
0 17289 7 1 2 32252 17288
0 17290 7 1 2 17287 17289
0 17291 5 1 1 17290
0 17292 7 1 2 17281 17291
0 17293 5 1 1 17292
0 17294 7 1 2 25513 17293
0 17295 5 1 1 17294
0 17296 7 1 2 30908 30040
0 17297 7 1 2 37520 17296
0 17298 7 1 2 37429 17297
0 17299 5 1 1 17298
0 17300 7 1 2 17295 17299
0 17301 5 1 1 17300
0 17302 7 1 2 29017 17301
0 17303 5 1 1 17302
0 17304 7 1 2 17277 17303
0 17305 5 1 1 17304
0 17306 7 1 2 24126 17305
0 17307 5 1 1 17306
0 17308 7 1 2 31416 37536
0 17309 5 1 1 17308
0 17310 7 1 2 17307 17309
0 17311 5 1 1 17310
0 17312 7 1 2 31266 17311
0 17313 5 1 1 17312
0 17314 7 1 2 17275 17313
0 17315 7 1 2 17157 17314
0 17316 7 1 2 17094 17315
0 17317 7 1 2 17052 17316
0 17318 7 1 2 16871 17317
0 17319 7 1 2 16564 17318
0 17320 5 1 1 17319
0 17321 7 1 2 23720 17320
0 17322 5 1 1 17321
0 17323 7 3 2 33541 29623
0 17324 7 2 2 35056 31260
0 17325 7 1 2 31994 31847
0 17326 7 1 2 37640 17325
0 17327 7 1 2 37656 17326
0 17328 7 1 2 37653 17327
0 17329 5 1 1 17328
0 17330 7 2 2 17322 17329
0 17331 5 1 1 37658
0 17332 7 1 2 23206 37659
0 17333 5 1 1 17332
0 17334 7 1 2 24347 17333
0 17335 7 1 2 15947 17334
0 17336 5 1 1 17335
0 17337 7 1 2 25134 17331
0 17338 5 1 1 17337
0 17339 7 1 2 36461 36033
0 17340 7 2 2 25088 33663
0 17341 5 1 1 37660
0 17342 7 1 2 37661 37310
0 17343 7 1 2 17339 17342
0 17344 7 1 2 25642 32312
0 17345 7 1 2 37657 17344
0 17346 7 1 2 17343 17345
0 17347 5 1 1 17346
0 17348 7 1 2 17338 17347
0 17349 5 1 1 17348
0 17350 7 1 2 22372 17349
0 17351 5 1 1 17350
0 17352 7 1 2 2204 3138
0 17353 5 1 1 17352
0 17354 7 3 2 5270 17353
0 17355 7 1 2 24485 37662
0 17356 5 1 1 17355
0 17357 7 2 2 25089 31309
0 17358 7 1 2 22498 37665
0 17359 5 1 1 17358
0 17360 7 1 2 17356 17359
0 17361 5 2 1 17360
0 17362 7 8 2 23721 34306
0 17363 7 1 2 30437 37669
0 17364 7 1 2 37667 17363
0 17365 5 2 1 17364
0 17366 7 2 2 23832 27987
0 17367 7 3 2 25318 36544
0 17368 7 1 2 34392 37681
0 17369 7 1 2 37679 17368
0 17370 5 2 1 17369
0 17371 7 3 2 25319 23722
0 17372 5 1 1 37686
0 17373 7 2 2 27219 37687
0 17374 7 1 2 34448 37689
0 17375 5 2 1 17374
0 17376 7 1 2 23723 35595
0 17377 5 1 1 17376
0 17378 7 1 2 23948 30452
0 17379 7 1 2 29452 17378
0 17380 5 1 1 17379
0 17381 7 1 2 17377 17380
0 17382 5 2 1 17381
0 17383 7 1 2 25816 37693
0 17384 5 1 1 17383
0 17385 7 1 2 31511 30148
0 17386 7 1 2 31154 17385
0 17387 5 1 1 17386
0 17388 7 1 2 17384 17387
0 17389 5 1 1 17388
0 17390 7 1 2 25135 17389
0 17391 5 1 1 17390
0 17392 7 1 2 37691 17391
0 17393 5 1 1 17392
0 17394 7 1 2 24991 17393
0 17395 5 1 1 17394
0 17396 7 1 2 37684 17395
0 17397 5 1 1 17396
0 17398 7 1 2 24348 17397
0 17399 5 1 1 17398
0 17400 7 1 2 37677 17399
0 17401 5 2 1 17400
0 17402 7 1 2 34437 37695
0 17403 5 1 1 17402
0 17404 7 3 2 22757 24992
0 17405 7 1 2 34501 34151
0 17406 7 1 2 37697 17405
0 17407 5 1 1 17406
0 17408 7 1 2 31197 34393
0 17409 7 1 2 31396 17408
0 17410 5 1 1 17409
0 17411 7 1 2 17407 17410
0 17412 5 1 1 17411
0 17413 7 1 2 24349 17412
0 17414 5 1 1 17413
0 17415 7 1 2 31397 34693
0 17416 7 1 2 36388 17415
0 17417 5 1 1 17416
0 17418 7 1 2 17414 17417
0 17419 5 1 1 17418
0 17420 7 1 2 27988 17419
0 17421 5 1 1 17420
0 17422 7 1 2 24350 34455
0 17423 5 1 1 17422
0 17424 7 4 2 25136 25232
0 17425 7 4 2 33783 37700
0 17426 5 1 1 37704
0 17427 7 1 2 17423 17426
0 17428 5 11 1 17427
0 17429 7 1 2 24993 34470
0 17430 7 1 2 37708 17429
0 17431 5 1 1 17430
0 17432 7 1 2 17421 17431
0 17433 5 1 1 17432
0 17434 7 1 2 23724 17433
0 17435 5 1 1 17434
0 17436 7 1 2 25817 34650
0 17437 7 3 2 34426 33399
0 17438 7 1 2 29453 37719
0 17439 7 1 2 17436 17438
0 17440 5 1 1 17439
0 17441 7 1 2 17435 17440
0 17442 5 1 1 17441
0 17443 7 1 2 27322 17442
0 17444 5 1 1 17443
0 17445 7 3 2 25090 23363
0 17446 5 1 1 37722
0 17447 7 1 2 37723 37318
0 17448 7 1 2 37709 17447
0 17449 5 1 1 17448
0 17450 7 1 2 31126 30622
0 17451 5 1 1 17450
0 17452 7 1 2 23151 28774
0 17453 7 1 2 31348 17452
0 17454 5 1 1 17453
0 17455 7 1 2 17451 17454
0 17456 5 1 1 17455
0 17457 7 1 2 24486 17456
0 17458 5 1 1 17457
0 17459 7 1 2 25233 23949
0 17460 7 1 2 35772 17459
0 17461 5 1 1 17460
0 17462 7 1 2 17458 17461
0 17463 5 1 1 17462
0 17464 7 3 2 24351 24994
0 17465 7 1 2 36475 37725
0 17466 7 1 2 17463 17465
0 17467 5 1 1 17466
0 17468 7 1 2 17449 17467
0 17469 5 1 1 17468
0 17470 7 1 2 22651 17469
0 17471 5 1 1 17470
0 17472 7 3 2 24705 29131
0 17473 7 1 2 23152 27025
0 17474 5 1 1 17473
0 17475 7 1 2 27293 17474
0 17476 5 3 1 17475
0 17477 7 1 2 24995 37720
0 17478 7 1 2 37731 17477
0 17479 7 1 2 37728 17478
0 17480 5 1 1 17479
0 17481 7 1 2 17471 17480
0 17482 5 1 1 17481
0 17483 7 1 2 23833 17482
0 17484 5 1 1 17483
0 17485 7 1 2 17444 17484
0 17486 7 1 2 17403 17485
0 17487 5 1 1 17486
0 17488 7 1 2 32459 17487
0 17489 5 1 1 17488
0 17490 7 2 2 34941 2650
0 17491 7 1 2 30136 33400
0 17492 7 1 2 37734 17491
0 17493 7 1 2 29260 17492
0 17494 5 1 1 17493
0 17495 7 4 2 25445 23725
0 17496 7 1 2 26104 37736
0 17497 7 1 2 30226 17496
0 17498 7 1 2 37710 17497
0 17499 5 1 1 17498
0 17500 7 1 2 17494 17499
0 17501 5 1 1 17500
0 17502 7 1 2 27145 37698
0 17503 7 1 2 17501 17502
0 17504 5 1 1 17503
0 17505 7 1 2 17489 17504
0 17506 5 1 1 17505
0 17507 7 1 2 36678 17506
0 17508 5 1 1 17507
0 17509 7 1 2 24487 34119
0 17510 5 1 1 17509
0 17511 7 1 2 31860 28065
0 17512 5 1 1 17511
0 17513 7 1 2 17510 17512
0 17514 5 4 1 17513
0 17515 7 2 2 37732 37740
0 17516 5 1 1 37744
0 17517 7 2 2 24352 33685
0 17518 7 3 2 23834 37746
0 17519 7 1 2 37745 37748
0 17520 5 1 1 17519
0 17521 7 1 2 23726 34126
0 17522 5 1 1 17521
0 17523 7 1 2 27722 35277
0 17524 7 1 2 34193 17523
0 17525 5 1 1 17524
0 17526 7 1 2 17522 17525
0 17527 5 1 1 17526
0 17528 7 1 2 25137 17527
0 17529 5 1 1 17528
0 17530 7 1 2 35574 34257
0 17531 5 1 1 17530
0 17532 7 1 2 17529 17531
0 17533 5 1 1 17532
0 17534 7 1 2 24353 17533
0 17535 5 1 1 17534
0 17536 7 3 2 28948 37670
0 17537 5 1 1 37751
0 17538 7 1 2 34114 37752
0 17539 5 1 1 17538
0 17540 7 1 2 17535 17539
0 17541 5 1 1 17540
0 17542 7 2 2 27323 17541
0 17543 5 1 1 37754
0 17544 7 1 2 25818 37755
0 17545 5 1 1 17544
0 17546 7 1 2 17520 17545
0 17547 5 1 1 17546
0 17548 7 1 2 24996 17547
0 17549 5 1 1 17548
0 17550 7 1 2 23727 28445
0 17551 7 2 2 37724 17550
0 17552 7 1 2 34330 37741
0 17553 5 1 1 17552
0 17554 7 1 2 34816 34009
0 17555 5 1 1 17554
0 17556 7 1 2 17553 17555
0 17557 5 1 1 17556
0 17558 7 1 2 37756 17557
0 17559 5 1 1 17558
0 17560 7 1 2 27260 27723
0 17561 5 1 1 17560
0 17562 7 5 2 25320 28446
0 17563 7 1 2 23279 37758
0 17564 5 1 1 17563
0 17565 7 1 2 17561 17564
0 17566 5 1 1 17565
0 17567 7 1 2 25714 17566
0 17568 5 1 1 17567
0 17569 7 1 2 27439 31613
0 17570 5 1 1 17569
0 17571 7 1 2 24488 17570
0 17572 7 1 2 17568 17571
0 17573 5 1 1 17572
0 17574 7 1 2 3454 17372
0 17575 7 4 2 34261 17574
0 17576 7 1 2 25234 37763
0 17577 5 1 1 17576
0 17578 7 1 2 28078 31591
0 17579 5 1 1 17578
0 17580 7 1 2 22499 17579
0 17581 7 1 2 17577 17580
0 17582 5 1 1 17581
0 17583 7 1 2 25138 17582
0 17584 7 1 2 17573 17583
0 17585 5 1 1 17584
0 17586 7 1 2 37692 17585
0 17587 5 1 1 17586
0 17588 7 1 2 24997 17587
0 17589 5 1 1 17588
0 17590 7 1 2 17589 37685
0 17591 5 1 1 17590
0 17592 7 1 2 24354 17591
0 17593 5 1 1 17592
0 17594 7 1 2 17593 37678
0 17595 5 1 1 17594
0 17596 7 1 2 34139 17595
0 17597 5 1 1 17596
0 17598 7 1 2 17559 17597
0 17599 7 1 2 17549 17598
0 17600 5 1 1 17599
0 17601 7 1 2 34986 17600
0 17602 5 1 1 17601
0 17603 7 1 2 33668 12775
0 17604 5 2 1 17603
0 17605 7 1 2 28949 37767
0 17606 5 1 1 17605
0 17607 7 1 2 25139 29672
0 17608 5 1 1 17607
0 17609 7 1 2 17606 17608
0 17610 5 2 1 17609
0 17611 7 1 2 24355 37769
0 17612 5 1 1 17611
0 17613 7 1 2 17537 17612
0 17614 5 2 1 17613
0 17615 7 1 2 32148 36077
0 17616 7 1 2 37771 17615
0 17617 5 1 1 17616
0 17618 7 1 2 36085 33401
0 17619 7 1 2 34525 17618
0 17620 5 1 1 17619
0 17621 7 1 2 17617 17620
0 17622 5 1 1 17621
0 17623 7 1 2 24998 17622
0 17624 5 1 1 17623
0 17625 7 2 2 30509 36327
0 17626 5 1 1 37773
0 17627 7 1 2 35330 37774
0 17628 5 1 1 17627
0 17629 7 1 2 32903 37711
0 17630 5 1 1 17629
0 17631 7 1 2 32909 36328
0 17632 5 1 1 17631
0 17633 7 1 2 17630 17632
0 17634 5 2 1 17633
0 17635 7 1 2 23484 30774
0 17636 7 1 2 37775 17635
0 17637 5 1 1 17636
0 17638 7 1 2 17628 17637
0 17639 5 1 1 17638
0 17640 7 4 2 23835 36426
0 17641 7 1 2 24039 37777
0 17642 7 1 2 17639 17641
0 17643 5 1 1 17642
0 17644 7 1 2 17624 17643
0 17645 7 1 2 17602 17644
0 17646 5 1 1 17645
0 17647 7 1 2 36575 17646
0 17648 5 1 1 17647
0 17649 7 3 2 25514 31375
0 17650 7 1 2 31428 37781
0 17651 5 1 1 17650
0 17652 7 1 2 24611 36642
0 17653 5 1 1 17652
0 17654 7 1 2 17651 17653
0 17655 5 1 1 17654
0 17656 7 1 2 37696 17655
0 17657 5 1 1 17656
0 17658 7 1 2 34560 36896
0 17659 5 1 1 17658
0 17660 7 3 2 31974 30116
0 17661 7 1 2 23280 37784
0 17662 5 1 1 17661
0 17663 7 1 2 17659 17662
0 17664 5 1 1 17663
0 17665 7 1 2 22500 17664
0 17666 5 1 1 17665
0 17667 7 2 2 23281 30137
0 17668 7 2 2 24489 36897
0 17669 7 1 2 37787 37789
0 17670 5 1 1 17669
0 17671 7 1 2 17666 17670
0 17672 5 1 1 17671
0 17673 7 1 2 25140 17672
0 17674 5 1 1 17673
0 17675 7 1 2 34449 37785
0 17676 5 1 1 17675
0 17677 7 1 2 17674 17676
0 17678 5 1 1 17677
0 17679 7 1 2 24356 17678
0 17680 5 1 1 17679
0 17681 7 1 2 37705 37786
0 17682 5 1 1 17681
0 17683 7 1 2 17680 17682
0 17684 5 1 1 17683
0 17685 7 1 2 36687 17684
0 17686 5 1 1 17685
0 17687 7 1 2 24490 36683
0 17688 5 1 1 17687
0 17689 7 1 2 29922 36218
0 17690 7 1 2 32313 17689
0 17691 5 1 1 17690
0 17692 7 1 2 17688 17691
0 17693 5 3 1 17692
0 17694 7 1 2 24999 34503
0 17695 5 1 1 17694
0 17696 7 1 2 34394 31929
0 17697 5 1 1 17696
0 17698 7 1 2 17695 17697
0 17699 5 1 1 17698
0 17700 7 1 2 24357 17699
0 17701 5 1 1 17700
0 17702 7 1 2 25141 30117
0 17703 7 1 2 34826 17702
0 17704 5 1 1 17703
0 17705 7 1 2 17701 17704
0 17706 5 1 1 17705
0 17707 7 1 2 37791 17706
0 17708 5 1 1 17707
0 17709 7 1 2 27156 33501
0 17710 7 1 2 36477 17709
0 17711 7 2 2 24358 28060
0 17712 7 1 2 36625 37794
0 17713 7 1 2 17710 17712
0 17714 5 1 1 17713
0 17715 7 1 2 17708 17714
0 17716 7 1 2 17686 17715
0 17717 5 1 1 17716
0 17718 7 1 2 23836 17717
0 17719 5 1 1 17718
0 17720 7 3 2 25515 36203
0 17721 7 2 2 28680 29607
0 17722 7 1 2 24359 25922
0 17723 7 1 2 27724 17722
0 17724 7 1 2 31342 17723
0 17725 7 1 2 37799 17724
0 17726 7 1 2 37796 17725
0 17727 5 1 1 17726
0 17728 7 1 2 17719 17727
0 17729 5 1 1 17728
0 17730 7 1 2 28860 17729
0 17731 5 1 1 17730
0 17732 7 2 2 25235 32232
0 17733 7 1 2 32370 32351
0 17734 7 1 2 37801 17733
0 17735 7 1 2 37797 17734
0 17736 5 1 1 17735
0 17737 7 2 2 36382 31873
0 17738 7 1 2 28606 37803
0 17739 5 1 1 17738
0 17740 7 2 2 24612 35057
0 17741 7 1 2 25387 30741
0 17742 7 1 2 37805 17741
0 17743 5 1 1 17742
0 17744 7 1 2 17739 17743
0 17745 5 3 1 17744
0 17746 7 1 2 22501 37807
0 17747 5 1 1 17746
0 17748 7 1 2 28348 36645
0 17749 5 1 1 17748
0 17750 7 1 2 17747 17749
0 17751 5 1 1 17750
0 17752 7 1 2 25142 17751
0 17753 5 1 1 17752
0 17754 7 1 2 34253 30558
0 17755 7 2 2 37806 17754
0 17756 5 1 1 37810
0 17757 7 1 2 24491 37811
0 17758 5 1 1 17757
0 17759 7 1 2 17753 17758
0 17760 5 1 1 17759
0 17761 7 1 2 23728 27324
0 17762 7 1 2 17760 17761
0 17763 5 1 1 17762
0 17764 7 1 2 17736 17763
0 17765 5 1 1 17764
0 17766 7 1 2 25819 17765
0 17767 5 1 1 17766
0 17768 7 1 2 24492 37808
0 17769 5 1 1 17768
0 17770 7 1 2 25236 34362
0 17771 7 1 2 37782 17770
0 17772 5 1 1 17771
0 17773 7 1 2 17769 17772
0 17774 5 1 1 17773
0 17775 7 1 2 30735 31512
0 17776 7 1 2 34734 17775
0 17777 7 1 2 17774 17776
0 17778 5 1 1 17777
0 17779 7 1 2 17767 17778
0 17780 5 1 1 17779
0 17781 7 1 2 25000 17780
0 17782 5 1 1 17781
0 17783 7 1 2 34814 36643
0 17784 5 1 1 17783
0 17785 7 1 2 17756 17784
0 17786 5 1 1 17785
0 17787 7 1 2 22502 17786
0 17788 5 1 1 17787
0 17789 7 1 2 33989 37809
0 17790 5 1 1 17789
0 17791 7 1 2 17788 17790
0 17792 5 1 1 17791
0 17793 7 1 2 37757 17792
0 17794 5 1 1 17793
0 17795 7 1 2 17782 17794
0 17796 5 1 1 17795
0 17797 7 1 2 24360 17796
0 17798 5 1 1 17797
0 17799 7 3 2 29363 27874
0 17800 5 1 1 37812
0 17801 7 1 2 35860 31059
0 17802 7 1 2 32003 17801
0 17803 7 1 2 37813 17802
0 17804 5 1 1 17803
0 17805 7 2 2 25820 27325
0 17806 7 1 2 32293 37815
0 17807 5 1 1 17806
0 17808 7 1 2 25091 31294
0 17809 5 1 1 17808
0 17810 7 1 2 17807 17809
0 17811 5 1 1 17810
0 17812 7 1 2 32346 37783
0 17813 7 1 2 17811 17812
0 17814 5 1 1 17813
0 17815 7 1 2 17804 17814
0 17816 5 1 1 17815
0 17817 7 1 2 24493 17816
0 17818 5 1 1 17817
0 17819 7 2 2 28447 30257
0 17820 7 1 2 28061 36219
0 17821 7 1 2 37802 17820
0 17822 7 1 2 37817 17821
0 17823 5 1 1 17822
0 17824 7 1 2 17818 17823
0 17825 5 1 1 17824
0 17826 7 1 2 37671 17825
0 17827 5 1 1 17826
0 17828 7 1 2 17798 17827
0 17829 7 1 2 17731 17828
0 17830 7 1 2 17657 17829
0 17831 5 1 1 17830
0 17832 7 1 2 32588 32460
0 17833 7 1 2 17831 17832
0 17834 5 1 1 17833
0 17835 7 2 2 27875 31908
0 17836 7 2 2 33664 37819
0 17837 5 1 1 37821
0 17838 7 1 2 33332 34561
0 17839 5 1 1 17838
0 17840 7 1 2 31957 17839
0 17841 5 1 1 17840
0 17842 7 1 2 22503 17841
0 17843 5 1 1 17842
0 17844 7 1 2 36357 37788
0 17845 5 1 1 17844
0 17846 7 1 2 17843 17845
0 17847 5 1 1 17846
0 17848 7 1 2 25143 17847
0 17849 5 1 1 17848
0 17850 7 1 2 17837 17849
0 17851 5 1 1 17850
0 17852 7 1 2 32439 17851
0 17853 5 1 1 17852
0 17854 7 2 2 24127 27989
0 17855 7 1 2 25715 27746
0 17856 7 1 2 36512 17855
0 17857 7 1 2 37823 17856
0 17858 5 1 1 17857
0 17859 7 1 2 17853 17858
0 17860 5 1 1 17859
0 17861 7 1 2 24361 17860
0 17862 5 1 1 17861
0 17863 7 2 2 34521 37701
0 17864 7 2 2 32440 30118
0 17865 7 1 2 37825 37827
0 17866 5 1 1 17865
0 17867 7 1 2 17862 17866
0 17868 5 1 1 17867
0 17869 7 1 2 36688 17868
0 17870 5 1 1 17869
0 17871 7 1 2 34504 37735
0 17872 5 1 1 17871
0 17873 7 1 2 25446 34417
0 17874 7 1 2 34528 17873
0 17875 5 1 1 17874
0 17876 7 1 2 17872 17875
0 17877 5 1 1 17876
0 17878 7 1 2 24362 17877
0 17879 5 1 1 17878
0 17880 7 1 2 35386 34307
0 17881 7 1 2 34529 17880
0 17882 5 1 1 17881
0 17883 7 1 2 17879 17882
0 17884 5 1 1 17883
0 17885 7 1 2 37792 17884
0 17886 5 1 1 17885
0 17887 7 1 2 27999 34010
0 17888 7 1 2 36685 17887
0 17889 7 1 2 34755 37828
0 17890 7 1 2 17888 17889
0 17891 5 1 1 17890
0 17892 7 1 2 17886 17891
0 17893 7 1 2 17870 17892
0 17894 5 1 1 17893
0 17895 7 1 2 23837 17894
0 17896 5 1 1 17895
0 17897 7 1 2 32708 34680
0 17898 7 1 2 32973 17897
0 17899 7 2 2 30851 37702
0 17900 7 1 2 24363 27108
0 17901 7 1 2 32352 17900
0 17902 7 1 2 37829 17901
0 17903 7 1 2 17898 17902
0 17904 5 1 1 17903
0 17905 7 1 2 17896 17904
0 17906 5 1 1 17905
0 17907 7 1 2 34843 17906
0 17908 5 1 1 17907
0 17909 7 3 2 25144 33784
0 17910 7 2 2 28315 37831
0 17911 5 1 1 37834
0 17912 7 1 2 24364 34300
0 17913 5 1 1 17912
0 17914 7 1 2 17911 17913
0 17915 5 1 1 17914
0 17916 7 1 2 37663 17915
0 17917 5 1 1 17916
0 17918 7 1 2 33966 34224
0 17919 5 1 1 17918
0 17920 7 1 2 25001 34214
0 17921 5 1 1 17920
0 17922 7 1 2 17919 17921
0 17923 5 1 1 17922
0 17924 7 1 2 24365 17923
0 17925 5 1 1 17924
0 17926 7 1 2 34308 37666
0 17927 5 1 1 17926
0 17928 7 1 2 17925 17927
0 17929 5 1 1 17928
0 17930 7 1 2 34303 17929
0 17931 5 1 1 17930
0 17932 7 1 2 17917 17931
0 17933 5 1 1 17932
0 17934 7 1 2 23729 17933
0 17935 5 1 1 17934
0 17936 7 1 2 28316 28289
0 17937 5 1 1 17936
0 17938 7 1 2 17800 17937
0 17939 5 1 1 17938
0 17940 7 1 2 24494 17939
0 17941 5 1 1 17940
0 17942 7 1 2 3213 17941
0 17943 5 4 1 17942
0 17944 7 1 2 36451 37726
0 17945 7 1 2 37836 17944
0 17946 5 1 1 17945
0 17947 7 1 2 17935 17946
0 17948 5 1 1 17947
0 17949 7 1 2 35928 36576
0 17950 7 1 2 17948 17949
0 17951 5 1 1 17950
0 17952 7 1 2 17908 17951
0 17953 7 1 2 17834 17952
0 17954 7 1 2 17648 17953
0 17955 7 1 2 17508 17954
0 17956 5 1 1 17955
0 17957 7 1 2 26194 17956
0 17958 5 1 1 17957
0 17959 7 1 2 23153 30227
0 17960 5 1 1 17959
0 17961 7 1 2 1042 17960
0 17962 5 1 1 17961
0 17963 7 1 2 23838 17962
0 17964 5 1 1 17963
0 17965 7 2 2 35901 28317
0 17966 7 1 2 23950 37840
0 17967 5 1 1 17966
0 17968 7 1 2 17964 17967
0 17969 5 1 1 17968
0 17970 7 1 2 25237 17969
0 17971 5 1 1 17970
0 17972 7 1 2 30654 37759
0 17973 5 2 1 17972
0 17974 7 1 2 17971 37842
0 17975 5 2 1 17974
0 17976 7 1 2 31105 37844
0 17977 5 1 1 17976
0 17978 7 2 2 27990 31609
0 17979 7 1 2 33244 37846
0 17980 5 1 1 17979
0 17981 7 3 2 25821 29423
0 17982 5 3 1 37848
0 17983 7 1 2 31523 37851
0 17984 5 1 1 17983
0 17985 7 1 2 17984 37253
0 17986 5 1 1 17985
0 17987 7 1 2 17980 17986
0 17988 7 1 2 17977 17987
0 17989 5 1 1 17988
0 17990 7 1 2 25145 17989
0 17991 5 1 1 17990
0 17992 7 1 2 36506 37690
0 17993 5 1 1 17992
0 17994 7 1 2 17991 17993
0 17995 5 1 1 17994
0 17996 7 1 2 25002 17995
0 17997 5 1 1 17996
0 17998 7 2 2 36427 33993
0 17999 7 1 2 28448 37854
0 18000 5 1 1 17999
0 18001 7 1 2 17997 18000
0 18002 5 1 1 18001
0 18003 7 1 2 27037 18002
0 18004 5 1 1 18003
0 18005 7 1 2 34296 31398
0 18006 7 1 2 37855 18005
0 18007 5 1 1 18006
0 18008 7 1 2 18004 18007
0 18009 5 1 1 18008
0 18010 7 1 2 24366 18009
0 18011 5 1 1 18010
0 18012 7 2 2 27004 29261
0 18013 5 1 1 37856
0 18014 7 1 2 34225 37857
0 18015 5 1 1 18014
0 18016 7 1 2 28634 32295
0 18017 5 1 1 18016
0 18018 7 1 2 18015 18017
0 18019 5 1 1 18018
0 18020 7 1 2 37672 18019
0 18021 5 1 1 18020
0 18022 7 1 2 18011 18021
0 18023 5 1 1 18022
0 18024 7 1 2 22758 18023
0 18025 5 1 1 18024
0 18026 7 1 2 31339 37770
0 18027 5 1 1 18026
0 18028 7 2 2 25716 33624
0 18029 5 1 1 37858
0 18030 7 1 2 17341 18029
0 18031 5 1 1 18030
0 18032 7 1 2 37680 18031
0 18033 5 1 1 18032
0 18034 7 1 2 18027 18033
0 18035 5 1 1 18034
0 18036 7 1 2 30510 18035
0 18037 5 1 1 18036
0 18038 7 1 2 23154 31521
0 18039 5 1 1 18038
0 18040 7 1 2 37852 18039
0 18041 5 3 1 18040
0 18042 7 1 2 34304 37860
0 18043 5 1 1 18042
0 18044 7 1 2 31985 31730
0 18045 5 1 1 18044
0 18046 7 1 2 30736 28290
0 18047 7 1 2 29610 18046
0 18048 5 1 1 18047
0 18049 7 1 2 18045 18048
0 18050 7 1 2 18043 18049
0 18051 5 1 1 18050
0 18052 7 1 2 25146 18051
0 18053 5 1 1 18052
0 18054 7 2 2 36507 37688
0 18055 5 1 1 37863
0 18056 7 1 2 25822 37864
0 18057 5 1 1 18056
0 18058 7 1 2 18053 18057
0 18059 5 1 1 18058
0 18060 7 1 2 36601 18059
0 18061 5 1 1 18060
0 18062 7 1 2 18037 18061
0 18063 5 1 1 18062
0 18064 7 1 2 24367 18063
0 18065 5 1 1 18064
0 18066 7 1 2 30511 37668
0 18067 5 1 1 18066
0 18068 7 1 2 31255 37790
0 18069 5 1 1 18068
0 18070 7 1 2 18067 18069
0 18071 5 1 1 18070
0 18072 7 1 2 37673 18071
0 18073 5 1 1 18072
0 18074 7 1 2 18065 18073
0 18075 5 1 1 18074
0 18076 7 1 2 34029 18075
0 18077 5 1 1 18076
0 18078 7 2 2 29262 34331
0 18079 5 1 1 37865
0 18080 7 2 2 36478 34369
0 18081 5 1 1 37867
0 18082 7 1 2 18079 18081
0 18083 5 2 1 18082
0 18084 7 1 2 27740 37778
0 18085 7 1 2 37869 18084
0 18086 5 1 1 18085
0 18087 7 1 2 18077 18086
0 18088 7 1 2 18025 18087
0 18089 5 1 1 18088
0 18090 7 1 2 33936 18089
0 18091 5 1 1 18090
0 18092 7 1 2 34736 37779
0 18093 5 1 1 18092
0 18094 7 2 2 27220 35575
0 18095 7 1 2 24495 34418
0 18096 7 1 2 37871 18095
0 18097 5 2 1 18096
0 18098 7 1 2 25238 37324
0 18099 5 1 1 18098
0 18100 7 3 2 23951 31622
0 18101 7 1 2 24613 37875
0 18102 5 1 1 18101
0 18103 7 2 2 18099 18102
0 18104 5 1 1 37878
0 18105 7 1 2 22504 37879
0 18106 5 1 1 18105
0 18107 7 1 2 31946 37861
0 18108 5 1 1 18107
0 18109 7 1 2 31826 34486
0 18110 5 1 1 18109
0 18111 7 1 2 24496 18110
0 18112 7 1 2 18108 18111
0 18113 5 1 1 18112
0 18114 7 1 2 25147 18113
0 18115 7 1 2 18106 18114
0 18116 5 1 1 18115
0 18117 7 1 2 37873 18116
0 18118 5 1 1 18117
0 18119 7 1 2 25003 18118
0 18120 5 1 1 18119
0 18121 7 1 2 18093 18120
0 18122 5 1 1 18121
0 18123 7 1 2 24368 18122
0 18124 5 1 1 18123
0 18125 7 1 2 33848 37664
0 18126 5 1 1 18125
0 18127 7 1 2 34226 34731
0 18128 5 1 1 18127
0 18129 7 1 2 18126 18128
0 18130 5 1 1 18129
0 18131 7 1 2 24497 18130
0 18132 5 1 1 18131
0 18133 7 1 2 25092 33880
0 18134 5 1 1 18133
0 18135 7 1 2 18132 18134
0 18136 5 1 1 18135
0 18137 7 1 2 37674 18136
0 18138 5 1 1 18137
0 18139 7 1 2 18124 18138
0 18140 5 1 1 18139
0 18141 7 1 2 34971 18140
0 18142 5 1 1 18141
0 18143 7 2 2 29835 27241
0 18144 7 1 2 31975 37737
0 18145 7 1 2 37880 18144
0 18146 7 1 2 37712 18145
0 18147 5 1 1 18146
0 18148 7 1 2 18142 18147
0 18149 5 1 1 18148
0 18150 7 1 2 32253 18149
0 18151 5 1 1 18150
0 18152 7 1 2 24498 37845
0 18153 5 1 1 18152
0 18154 7 1 2 31389 37760
0 18155 5 2 1 18154
0 18156 7 1 2 18153 37882
0 18157 5 1 1 18156
0 18158 7 1 2 33191 18157
0 18159 5 1 1 18158
0 18160 7 1 2 25823 37174
0 18161 5 1 1 18160
0 18162 7 1 2 31641 5370
0 18163 5 2 1 18162
0 18164 7 2 2 23839 37884
0 18165 7 1 2 22505 37886
0 18166 5 1 1 18165
0 18167 7 1 2 18161 18166
0 18168 5 1 1 18167
0 18169 7 1 2 34515 30203
0 18170 7 1 2 18168 18169
0 18171 5 1 1 18170
0 18172 7 1 2 18159 18171
0 18173 5 1 1 18172
0 18174 7 1 2 32473 33686
0 18175 7 1 2 37727 18174
0 18176 7 1 2 18173 18175
0 18177 5 1 1 18176
0 18178 7 1 2 24369 36351
0 18179 5 1 1 18178
0 18180 7 1 2 34309 33883
0 18181 5 1 1 18180
0 18182 7 1 2 18179 18181
0 18183 5 1 1 18182
0 18184 7 1 2 35387 36166
0 18185 7 1 2 37881 18184
0 18186 5 1 1 18185
0 18187 7 1 2 23840 36167
0 18188 5 1 1 18187
0 18189 7 1 2 15776 18188
0 18190 5 1 1 18189
0 18191 7 1 2 31688 34972
0 18192 7 1 2 18190 18191
0 18193 5 1 1 18192
0 18194 7 1 2 18186 18193
0 18195 5 1 1 18194
0 18196 7 1 2 18183 18195
0 18197 5 1 1 18196
0 18198 7 1 2 27227 36898
0 18199 5 1 1 18198
0 18200 7 1 2 13444 17446
0 18201 5 1 1 18200
0 18202 7 1 2 27444 18201
0 18203 5 1 1 18202
0 18204 7 1 2 14235 18203
0 18205 5 1 1 18204
0 18206 7 1 2 23841 8149
0 18207 7 1 2 18205 18206
0 18208 5 1 1 18207
0 18209 7 1 2 18199 18208
0 18210 5 1 1 18209
0 18211 7 1 2 37713 18210
0 18212 5 1 1 18211
0 18213 7 1 2 33625 34801
0 18214 5 1 1 18213
0 18215 7 1 2 34761 37761
0 18216 5 1 1 18215
0 18217 7 1 2 18214 18216
0 18218 5 1 1 18217
0 18219 7 1 2 24370 18218
0 18220 5 1 1 18219
0 18221 7 1 2 25148 34827
0 18222 7 1 2 37762 18221
0 18223 5 1 1 18222
0 18224 7 1 2 18220 18223
0 18225 5 1 1 18224
0 18226 7 1 2 27991 18225
0 18227 5 1 1 18226
0 18228 7 1 2 18212 18227
0 18229 5 1 1 18228
0 18230 7 1 2 32474 33192
0 18231 7 1 2 18229 18230
0 18232 5 1 1 18231
0 18233 7 1 2 18197 18232
0 18234 5 1 1 18233
0 18235 7 1 2 23730 18234
0 18236 5 1 1 18235
0 18237 7 2 2 23731 31689
0 18238 7 1 2 25004 36124
0 18239 5 1 1 18238
0 18240 7 1 2 5800 18239
0 18241 5 1 1 18240
0 18242 7 1 2 24371 18241
0 18243 5 1 1 18242
0 18244 7 1 2 34227 37832
0 18245 5 1 1 18244
0 18246 7 1 2 18243 18245
0 18247 5 1 1 18246
0 18248 7 1 2 37888 18247
0 18249 5 1 1 18248
0 18250 7 2 2 24372 24499
0 18251 7 1 2 37890 37859
0 18252 7 1 2 37887 18251
0 18253 5 1 1 18252
0 18254 7 1 2 18249 18253
0 18255 5 1 1 18254
0 18256 7 1 2 34973 18255
0 18257 5 1 1 18256
0 18258 7 1 2 29836 29608
0 18259 7 1 2 37738 18258
0 18260 7 1 2 34332 34230
0 18261 7 1 2 18259 18260
0 18262 5 1 1 18261
0 18263 7 1 2 18257 18262
0 18264 5 1 1 18263
0 18265 7 1 2 32850 18264
0 18266 5 1 1 18265
0 18267 7 1 2 18236 18266
0 18268 7 1 2 18177 18267
0 18269 7 1 2 18151 18268
0 18270 5 1 1 18269
0 18271 7 1 2 22857 18270
0 18272 5 1 1 18271
0 18273 7 1 2 23732 27242
0 18274 7 1 2 476 35231
0 18275 7 1 2 18273 18274
0 18276 7 1 2 34992 18275
0 18277 7 1 2 37776 18276
0 18278 5 1 1 18277
0 18279 7 1 2 18272 18278
0 18280 7 1 2 18091 18279
0 18281 5 1 1 18280
0 18282 7 1 2 30368 18281
0 18283 5 1 1 18282
0 18284 7 1 2 17958 18283
0 18285 5 1 1 18284
0 18286 7 1 2 33429 34873
0 18287 7 1 2 18285 18286
0 18288 5 1 1 18287
0 18289 7 3 2 26105 27146
0 18290 7 1 2 29285 35314
0 18291 5 2 1 18290
0 18292 7 3 2 23591 32992
0 18293 7 1 2 35853 37897
0 18294 5 1 1 18293
0 18295 7 1 2 37895 18294
0 18296 5 1 1 18295
0 18297 7 1 2 22858 18296
0 18298 5 1 1 18297
0 18299 7 3 2 32993 37382
0 18300 7 1 2 27650 37900
0 18301 5 1 1 18300
0 18302 7 1 2 18298 18301
0 18303 5 3 1 18302
0 18304 7 1 2 27758 37903
0 18305 5 1 1 18304
0 18306 7 3 2 25447 35744
0 18307 7 1 2 35324 37906
0 18308 5 1 1 18307
0 18309 7 1 2 18305 18308
0 18310 5 1 1 18309
0 18311 7 1 2 34562 18310
0 18312 5 1 1 18311
0 18313 7 2 2 32994 37024
0 18314 7 1 2 25923 31281
0 18315 7 1 2 28886 18314
0 18316 7 1 2 37909 18315
0 18317 5 1 1 18316
0 18318 7 1 2 18312 18317
0 18319 5 1 1 18318
0 18320 7 1 2 24706 18319
0 18321 5 1 1 18320
0 18322 7 1 2 25388 37904
0 18323 5 1 1 18322
0 18324 7 2 2 26841 35745
0 18325 5 1 1 37911
0 18326 7 2 2 24790 37912
0 18327 5 1 1 37913
0 18328 7 1 2 18323 18327
0 18329 5 1 1 18328
0 18330 7 1 2 28761 34563
0 18331 7 1 2 18329 18330
0 18332 5 1 1 18331
0 18333 7 1 2 18321 18332
0 18334 5 1 1 18333
0 18335 7 1 2 25149 18334
0 18336 5 1 1 18335
0 18337 7 1 2 24707 28681
0 18338 7 1 2 33793 18337
0 18339 7 1 2 35395 36484
0 18340 7 1 2 18338 18339
0 18341 5 1 1 18340
0 18342 7 1 2 18336 18341
0 18343 5 1 1 18342
0 18344 7 1 2 22506 18343
0 18345 5 1 1 18344
0 18346 7 1 2 32117 37905
0 18347 5 1 1 18346
0 18348 7 1 2 22759 37914
0 18349 5 1 1 18348
0 18350 7 1 2 18347 18349
0 18351 5 2 1 18350
0 18352 7 1 2 25321 37915
0 18353 5 1 1 18352
0 18354 7 2 2 28797 35746
0 18355 5 1 1 37917
0 18356 7 1 2 27343 37918
0 18357 5 1 1 18356
0 18358 7 1 2 18353 18357
0 18359 5 1 1 18358
0 18360 7 1 2 27914 34412
0 18361 7 1 2 18359 18360
0 18362 5 1 1 18361
0 18363 7 1 2 18345 18362
0 18364 5 1 1 18363
0 18365 7 1 2 24614 18364
0 18366 5 1 1 18365
0 18367 7 1 2 29213 37916
0 18368 5 1 1 18367
0 18369 7 2 2 35747 34365
0 18370 5 1 1 37919
0 18371 7 1 2 27344 37920
0 18372 5 1 1 18371
0 18373 7 1 2 18368 18372
0 18374 5 1 1 18373
0 18375 7 1 2 24500 34505
0 18376 7 1 2 18374 18375
0 18377 5 1 1 18376
0 18378 7 1 2 18366 18377
0 18379 5 1 1 18378
0 18380 7 1 2 24373 18379
0 18381 5 1 1 18380
0 18382 7 1 2 27926 34310
0 18383 7 1 2 36440 30492
0 18384 7 1 2 18382 18383
0 18385 7 1 2 31548 37570
0 18386 7 1 2 18384 18385
0 18387 5 1 1 18386
0 18388 7 1 2 18381 18387
0 18389 5 1 1 18388
0 18390 7 1 2 37892 18389
0 18391 5 1 1 18390
0 18392 7 1 2 1740 1323
0 18393 5 1 1 18392
0 18394 7 1 2 25150 18393
0 18395 5 1 1 18394
0 18396 7 1 2 18055 18395
0 18397 5 1 1 18396
0 18398 7 1 2 24374 18397
0 18399 5 1 1 18398
0 18400 7 1 2 35576 37835
0 18401 5 1 1 18400
0 18402 7 1 2 18399 18401
0 18403 5 2 1 18402
0 18404 7 1 2 32880 37921
0 18405 5 1 1 18404
0 18406 7 1 2 31564 33402
0 18407 7 1 2 30353 18406
0 18408 5 1 1 18407
0 18409 7 1 2 18405 18408
0 18410 5 1 1 18409
0 18411 7 1 2 25824 18410
0 18412 5 1 1 18411
0 18413 7 1 2 34476 33136
0 18414 5 1 1 18413
0 18415 7 1 2 32766 37296
0 18416 5 1 1 18415
0 18417 7 1 2 18414 18416
0 18418 5 1 1 18417
0 18419 7 3 2 28167 18418
0 18420 5 1 1 37923
0 18421 7 1 2 37772 37924
0 18422 5 1 1 18421
0 18423 7 1 2 24615 37733
0 18424 5 1 1 18423
0 18425 7 1 2 30889 18424
0 18426 5 1 1 18425
0 18427 7 1 2 27992 18426
0 18428 5 1 1 18427
0 18429 7 2 2 27725 27440
0 18430 5 1 1 37926
0 18431 7 1 2 28349 37927
0 18432 5 1 1 18431
0 18433 7 1 2 18428 18432
0 18434 5 1 1 18433
0 18435 7 1 2 23842 33137
0 18436 7 1 2 37721 18435
0 18437 7 1 2 18434 18436
0 18438 5 1 1 18437
0 18439 7 1 2 18422 18438
0 18440 7 1 2 18412 18439
0 18441 5 1 1 18440
0 18442 7 1 2 32118 18441
0 18443 5 1 1 18442
0 18444 7 1 2 25151 37694
0 18445 5 1 1 18444
0 18446 7 1 2 34450 37682
0 18447 5 1 1 18446
0 18448 7 1 2 18445 18447
0 18449 5 1 1 18448
0 18450 7 1 2 24375 18449
0 18451 5 1 1 18450
0 18452 7 1 2 37706 37683
0 18453 5 1 1 18452
0 18454 7 1 2 18451 18453
0 18455 5 1 1 18454
0 18456 7 1 2 34140 18455
0 18457 5 1 1 18456
0 18458 7 1 2 17543 18457
0 18459 5 1 1 18458
0 18460 7 1 2 25825 18459
0 18461 5 1 1 18460
0 18462 7 1 2 31151 18430
0 18463 5 1 1 18462
0 18464 7 1 2 24501 18463
0 18465 5 1 1 18464
0 18466 7 1 2 31249 18465
0 18467 5 1 1 18466
0 18468 7 1 2 34141 18467
0 18469 5 1 1 18468
0 18470 7 1 2 17516 18469
0 18471 5 1 1 18470
0 18472 7 1 2 18471 37749
0 18473 5 1 1 18472
0 18474 7 1 2 18461 18473
0 18475 5 1 1 18474
0 18476 7 1 2 32933 18475
0 18477 5 1 1 18476
0 18478 7 1 2 18443 18477
0 18479 5 2 1 18478
0 18480 7 1 2 25448 37898
0 18481 5 1 1 18480
0 18482 7 1 2 18481 37896
0 18483 5 1 1 18482
0 18484 7 1 2 37928 18483
0 18485 5 1 1 18484
0 18486 7 1 2 25389 37901
0 18487 5 1 1 18486
0 18488 7 1 2 18325 18487
0 18489 5 1 1 18488
0 18490 7 1 2 25826 32809
0 18491 7 1 2 37922 18490
0 18492 5 1 1 18491
0 18493 7 1 2 32176 37753
0 18494 5 1 1 18493
0 18495 7 1 2 27702 37876
0 18496 5 1 1 18495
0 18497 7 1 2 25239 37316
0 18498 5 1 1 18497
0 18499 7 1 2 22507 18498
0 18500 7 1 2 18496 18499
0 18501 5 1 1 18500
0 18502 7 1 2 33265 37862
0 18503 5 1 1 18502
0 18504 7 1 2 30138 27703
0 18505 7 1 2 31827 18504
0 18506 5 1 1 18505
0 18507 7 1 2 24502 18506
0 18508 7 1 2 18503 18507
0 18509 5 1 1 18508
0 18510 7 1 2 25152 18509
0 18511 7 1 2 18501 18510
0 18512 5 1 1 18511
0 18513 7 1 2 31127 31610
0 18514 7 1 2 36610 18513
0 18515 5 1 1 18514
0 18516 7 1 2 18512 18515
0 18517 5 1 1 18516
0 18518 7 1 2 24376 18517
0 18519 5 1 1 18518
0 18520 7 1 2 18494 18519
0 18521 5 1 1 18520
0 18522 7 1 2 28168 18521
0 18523 5 1 1 18522
0 18524 7 1 2 33263 37747
0 18525 7 1 2 31819 18524
0 18526 5 1 1 18525
0 18527 7 1 2 18523 18526
0 18528 7 1 2 18492 18527
0 18529 5 1 1 18528
0 18530 7 1 2 33148 18529
0 18531 5 1 1 18530
0 18532 7 1 2 30348 36634
0 18533 7 1 2 34725 18532
0 18534 7 1 2 37714 18533
0 18535 5 1 1 18534
0 18536 7 2 2 26976 31513
0 18537 7 1 2 24377 32531
0 18538 7 1 2 34282 18537
0 18539 7 1 2 37930 18538
0 18540 7 1 2 29263 18539
0 18541 5 1 1 18540
0 18542 7 1 2 18535 18541
0 18543 7 1 2 18531 18542
0 18544 5 2 1 18543
0 18545 7 1 2 18489 37932
0 18546 5 1 1 18545
0 18547 7 1 2 36005 37899
0 18548 5 1 1 18547
0 18549 7 1 2 18355 18548
0 18550 5 1 1 18549
0 18551 7 1 2 23733 37143
0 18552 5 1 1 18551
0 18553 7 1 2 36358 34564
0 18554 5 1 1 18553
0 18555 7 1 2 18552 18554
0 18556 5 1 1 18555
0 18557 7 1 2 25827 18556
0 18558 5 1 1 18557
0 18559 7 5 2 25924 31514
0 18560 7 1 2 27726 28350
0 18561 7 1 2 37934 18560
0 18562 5 1 1 18561
0 18563 7 1 2 18558 18562
0 18564 5 1 1 18563
0 18565 7 1 2 25153 18564
0 18566 5 1 1 18565
0 18567 7 1 2 18566 37874
0 18568 5 1 1 18567
0 18569 7 1 2 24378 18568
0 18570 5 1 1 18569
0 18571 7 1 2 33785 36513
0 18572 7 1 2 37872 18571
0 18573 5 1 1 18572
0 18574 7 1 2 18570 18573
0 18575 5 1 1 18574
0 18576 7 1 2 32589 18575
0 18577 5 1 1 18576
0 18578 7 1 2 27459 33403
0 18579 7 1 2 28456 18578
0 18580 7 1 2 36585 18579
0 18581 5 1 1 18580
0 18582 7 1 2 18577 18581
0 18583 5 1 1 18582
0 18584 7 1 2 32557 18583
0 18585 5 1 1 18584
0 18586 7 2 2 32532 30139
0 18587 7 1 2 30579 37939
0 18588 5 1 1 18587
0 18589 7 2 2 31429 34530
0 18590 7 1 2 23282 37941
0 18591 5 1 1 18590
0 18592 7 1 2 18588 18591
0 18593 5 1 1 18592
0 18594 7 1 2 22508 18593
0 18595 5 1 1 18594
0 18596 7 1 2 24128 34487
0 18597 7 1 2 32975 18596
0 18598 5 1 1 18597
0 18599 7 1 2 18595 18598
0 18600 5 1 1 18599
0 18601 7 1 2 25154 18600
0 18602 5 1 1 18601
0 18603 7 1 2 32517 37822
0 18604 5 1 1 18603
0 18605 7 1 2 18602 18604
0 18606 5 1 1 18605
0 18607 7 1 2 24379 18606
0 18608 5 1 1 18607
0 18609 7 1 2 37707 37942
0 18610 5 1 1 18609
0 18611 7 1 2 18608 18610
0 18612 5 1 1 18611
0 18613 7 1 2 23843 30177
0 18614 7 1 2 18612 18613
0 18615 5 1 1 18614
0 18616 7 1 2 18585 18615
0 18617 5 2 1 18616
0 18618 7 1 2 18550 37943
0 18619 5 1 1 18618
0 18620 7 1 2 33032 37902
0 18621 5 1 1 18620
0 18622 7 1 2 18370 18621
0 18623 5 1 1 18622
0 18624 7 1 2 36925 37286
0 18625 5 1 1 18624
0 18626 7 1 2 32590 36359
0 18627 7 1 2 37935 18626
0 18628 5 1 1 18627
0 18629 7 1 2 37393 18628
0 18630 5 1 1 18629
0 18631 7 1 2 33149 18630
0 18632 5 1 1 18631
0 18633 7 1 2 18625 18632
0 18634 5 1 1 18633
0 18635 7 1 2 25155 18634
0 18636 5 1 1 18635
0 18637 7 5 2 23734 23844
0 18638 7 2 2 30349 37945
0 18639 7 2 2 27829 37950
0 18640 7 1 2 33990 37952
0 18641 5 1 1 18640
0 18642 7 1 2 18636 18641
0 18643 5 1 1 18642
0 18644 7 1 2 24380 18643
0 18645 5 1 1 18644
0 18646 7 1 2 37833 37953
0 18647 5 1 1 18646
0 18648 7 1 2 18645 18647
0 18649 5 2 1 18648
0 18650 7 1 2 18623 37954
0 18651 5 1 1 18650
0 18652 7 2 2 31690 31464
0 18653 7 1 2 28405 37910
0 18654 5 1 1 18653
0 18655 7 1 2 27727 29292
0 18656 7 1 2 37571 18655
0 18657 5 1 1 18656
0 18658 7 1 2 18654 18657
0 18659 5 1 1 18658
0 18660 7 1 2 25156 18659
0 18661 5 1 1 18660
0 18662 7 1 2 25322 34757
0 18663 7 1 2 37907 18662
0 18664 5 1 1 18663
0 18665 7 1 2 18661 18664
0 18666 5 1 1 18665
0 18667 7 1 2 24381 18666
0 18668 5 1 1 18667
0 18669 7 1 2 32314 37675
0 18670 7 1 2 37908 18669
0 18671 5 1 1 18670
0 18672 7 1 2 18668 18671
0 18673 5 1 1 18672
0 18674 7 1 2 37956 18673
0 18675 5 1 1 18674
0 18676 7 1 2 34011 37703
0 18677 7 1 2 37572 18676
0 18678 7 1 2 29294 18677
0 18679 7 1 2 37885 18678
0 18680 5 1 1 18679
0 18681 7 1 2 18675 18680
0 18682 5 1 1 18681
0 18683 7 1 2 33104 18682
0 18684 5 1 1 18683
0 18685 7 1 2 18651 18684
0 18686 7 1 2 18619 18685
0 18687 7 1 2 18546 18686
0 18688 7 1 2 18485 18687
0 18689 7 1 2 18391 18688
0 18690 5 1 1 18689
0 18691 7 1 2 29120 18690
0 18692 5 1 1 18691
0 18693 7 1 2 32738 37929
0 18694 5 1 1 18693
0 18695 7 1 2 33061 37933
0 18696 5 1 1 18695
0 18697 7 1 2 32656 37944
0 18698 5 1 1 18697
0 18699 7 1 2 32683 37955
0 18700 5 1 1 18699
0 18701 7 1 2 36207 37633
0 18702 5 1 1 18701
0 18703 7 1 2 22979 34199
0 18704 7 1 2 32689 18703
0 18705 5 1 1 18704
0 18706 7 1 2 18702 18705
0 18707 5 1 1 18706
0 18708 7 1 2 32518 31930
0 18709 7 1 2 18707 18708
0 18710 5 1 1 18709
0 18711 7 2 2 25157 29589
0 18712 7 1 2 37958 37940
0 18713 7 1 2 36843 18712
0 18714 5 1 1 18713
0 18715 7 1 2 18710 18714
0 18716 5 1 1 18715
0 18717 7 1 2 24382 18716
0 18718 5 1 1 18717
0 18719 7 1 2 25323 35283
0 18720 7 1 2 35257 18719
0 18721 7 2 2 37676 18720
0 18722 5 1 1 37960
0 18723 7 1 2 30775 32347
0 18724 7 1 2 37961 18723
0 18725 5 1 1 18724
0 18726 7 1 2 18718 18725
0 18727 5 1 1 18726
0 18728 7 1 2 27147 30698
0 18729 7 1 2 18727 18728
0 18730 5 1 1 18729
0 18731 7 2 2 25158 32406
0 18732 7 1 2 35269 37962
0 18733 5 1 1 18732
0 18734 7 1 2 35284 37634
0 18735 7 1 2 37768 18734
0 18736 5 1 1 18735
0 18737 7 1 2 18733 18736
0 18738 5 1 1 18737
0 18739 7 1 2 24383 18738
0 18740 5 1 1 18739
0 18741 7 1 2 18722 18740
0 18742 5 1 1 18741
0 18743 7 1 2 37957 18742
0 18744 5 1 1 18743
0 18745 7 1 2 37635 37936
0 18746 7 1 2 37830 37795
0 18747 7 1 2 18745 18746
0 18748 5 1 1 18747
0 18749 7 1 2 18744 18748
0 18750 5 1 1 18749
0 18751 7 1 2 32591 18750
0 18752 5 1 1 18751
0 18753 7 1 2 35285 34283
0 18754 7 1 2 34664 18753
0 18755 7 1 2 34370 37636
0 18756 7 1 2 18754 18755
0 18757 5 1 1 18756
0 18758 7 1 2 18752 18757
0 18759 5 1 1 18758
0 18760 7 1 2 33150 18759
0 18761 5 1 1 18760
0 18762 7 1 2 18730 18761
0 18763 7 1 2 18700 18762
0 18764 7 1 2 18698 18763
0 18765 7 1 2 18696 18764
0 18766 7 1 2 18694 18765
0 18767 5 1 1 18766
0 18768 7 1 2 33430 36872
0 18769 5 1 1 18768
0 18770 7 1 2 29290 18769
0 18771 7 1 2 18767 18770
0 18772 5 1 1 18771
0 18773 7 1 2 22859 32739
0 18774 5 1 1 18773
0 18775 7 1 2 7879 18774
0 18776 5 1 1 18775
0 18777 7 1 2 37609 18776
0 18778 5 1 1 18777
0 18779 7 1 2 34170 28950
0 18780 5 1 1 18779
0 18781 7 1 2 37367 18780
0 18782 5 2 1 18781
0 18783 7 1 2 32620 35058
0 18784 7 1 2 37964 18783
0 18785 5 1 1 18784
0 18786 7 1 2 18778 18785
0 18787 5 1 1 18786
0 18788 7 1 2 9016 16654
0 18789 5 1 1 18788
0 18790 7 1 2 32870 37750
0 18791 7 1 2 18789 18790
0 18792 7 1 2 18787 18791
0 18793 5 1 1 18792
0 18794 7 1 2 18772 18793
0 18795 7 1 2 18692 18794
0 18796 5 1 1 18795
0 18797 7 1 2 23055 18796
0 18798 5 1 1 18797
0 18799 7 2 2 34284 34763
0 18800 7 1 2 23592 24305
0 18801 7 2 2 29768 18800
0 18802 7 1 2 37966 37968
0 18803 5 1 1 18802
0 18804 7 1 2 30077 37969
0 18805 5 1 1 18804
0 18806 7 1 2 24708 37377
0 18807 7 1 2 35536 18806
0 18808 5 1 1 18807
0 18809 7 1 2 18805 18808
0 18810 5 1 1 18809
0 18811 7 1 2 24503 18810
0 18812 5 1 1 18811
0 18813 7 1 2 22509 30879
0 18814 7 1 2 27547 30204
0 18815 7 1 2 18813 18814
0 18816 5 1 1 18815
0 18817 7 1 2 18812 18816
0 18818 5 1 1 18817
0 18819 7 1 2 34333 18818
0 18820 5 1 1 18819
0 18821 7 1 2 18803 18820
0 18822 5 1 1 18821
0 18823 7 1 2 32533 18822
0 18824 5 1 1 18823
0 18825 7 1 2 27345 30927
0 18826 7 1 2 35537 18825
0 18827 7 1 2 36329 18826
0 18828 5 1 1 18827
0 18829 7 1 2 18824 18828
0 18830 5 1 1 18829
0 18831 7 1 2 28169 18830
0 18832 5 1 1 18831
0 18833 7 3 2 32810 32558
0 18834 7 1 2 27548 37970
0 18835 7 1 2 37870 18834
0 18836 5 1 1 18835
0 18837 7 1 2 18832 18836
0 18838 5 1 1 18837
0 18839 7 1 2 33062 18838
0 18840 5 1 1 18839
0 18841 7 1 2 32881 37866
0 18842 5 1 1 18841
0 18843 7 2 2 25925 34371
0 18844 7 1 2 36479 37973
0 18845 5 1 1 18844
0 18846 7 1 2 17626 18845
0 18847 5 2 1 18846
0 18848 7 1 2 32876 37975
0 18849 5 1 1 18848
0 18850 7 1 2 34012 33906
0 18851 7 1 2 32871 18850
0 18852 7 1 2 36247 18851
0 18853 5 1 1 18852
0 18854 7 1 2 18849 18853
0 18855 7 1 2 18842 18854
0 18856 5 1 1 18855
0 18857 7 1 2 32119 18856
0 18858 5 1 1 18857
0 18859 7 1 2 31664 32920
0 18860 5 1 1 18859
0 18861 7 1 2 35624 18860
0 18862 5 2 1 18861
0 18863 7 1 2 27391 37967
0 18864 7 1 2 37977 18863
0 18865 5 1 1 18864
0 18866 7 1 2 18858 18865
0 18867 5 1 1 18866
0 18868 7 1 2 27549 18867
0 18869 5 1 1 18868
0 18870 7 2 2 31947 37715
0 18871 7 2 2 35918 37541
0 18872 5 1 1 37981
0 18873 7 1 2 33015 34850
0 18874 5 1 1 18873
0 18875 7 1 2 18872 18874
0 18876 5 1 1 18875
0 18877 7 1 2 37979 18876
0 18878 5 1 1 18877
0 18879 7 2 2 29942 36899
0 18880 7 1 2 32934 37983
0 18881 7 1 2 36330 18880
0 18882 5 1 1 18881
0 18883 7 1 2 18878 18882
0 18884 5 1 1 18883
0 18885 7 1 2 32254 18884
0 18886 5 1 1 18885
0 18887 7 1 2 27550 37978
0 18888 5 1 1 18887
0 18889 7 2 2 31665 35919
0 18890 7 1 2 37542 37985
0 18891 5 1 1 18890
0 18892 7 1 2 18888 18891
0 18893 5 1 1 18892
0 18894 7 1 2 34334 33877
0 18895 7 1 2 18893 18894
0 18896 5 1 1 18895
0 18897 7 1 2 31666 34013
0 18898 7 1 2 36348 18897
0 18899 7 1 2 37982 18898
0 18900 5 1 1 18899
0 18901 7 1 2 18896 18900
0 18902 7 1 2 18886 18901
0 18903 7 1 2 18869 18902
0 18904 5 1 1 18903
0 18905 7 1 2 32740 18904
0 18906 5 1 1 18905
0 18907 7 2 2 23593 33363
0 18908 7 1 2 35920 37987
0 18909 5 1 1 18908
0 18910 7 1 2 27551 36837
0 18911 5 1 1 18910
0 18912 7 1 2 18909 18911
0 18913 5 1 1 18912
0 18914 7 1 2 37980 18913
0 18915 5 1 1 18914
0 18916 7 1 2 33105 37984
0 18917 7 1 2 36331 18916
0 18918 5 1 1 18917
0 18919 7 1 2 18915 18918
0 18920 5 1 1 18919
0 18921 7 1 2 32657 18920
0 18922 5 1 1 18921
0 18923 7 1 2 26955 27460
0 18924 5 1 1 18923
0 18925 7 1 2 9535 18924
0 18926 5 7 1 18925
0 18927 7 1 2 27552 32559
0 18928 7 1 2 37989 18927
0 18929 5 1 1 18928
0 18930 7 1 2 37986 37988
0 18931 5 1 1 18930
0 18932 7 1 2 18929 18931
0 18933 5 1 1 18932
0 18934 7 1 2 24504 32684
0 18935 5 1 1 18934
0 18936 7 1 2 31761 37637
0 18937 5 1 1 18936
0 18938 7 1 2 18935 18937
0 18939 5 2 1 18938
0 18940 7 1 2 34335 37996
0 18941 5 1 1 18940
0 18942 7 1 2 34858 34014
0 18943 7 1 2 37963 18942
0 18944 5 1 1 18943
0 18945 7 1 2 18941 18944
0 18946 5 1 1 18945
0 18947 7 1 2 18933 18946
0 18948 5 1 1 18947
0 18949 7 1 2 18922 18948
0 18950 7 1 2 18906 18949
0 18951 7 1 2 18840 18950
0 18952 5 1 1 18951
0 18953 7 1 2 26195 18952
0 18954 5 1 1 18953
0 18955 7 1 2 36159 37716
0 18956 5 1 1 18955
0 18957 7 1 2 30898 36332
0 18958 5 1 1 18957
0 18959 7 1 2 18956 18958
0 18960 5 1 1 18959
0 18961 7 1 2 34030 18960
0 18962 5 1 1 18961
0 18963 7 1 2 33245 37717
0 18964 5 1 1 18963
0 18965 7 1 2 33890 36333
0 18966 5 1 1 18965
0 18967 7 1 2 18964 18966
0 18968 5 1 1 18967
0 18969 7 1 2 30994 18968
0 18970 5 1 1 18969
0 18971 7 1 2 18962 18970
0 18972 5 1 1 18971
0 18973 7 1 2 34274 18972
0 18974 5 1 1 18973
0 18975 7 1 2 24505 33039
0 18976 5 1 1 18975
0 18977 7 1 2 16789 18976
0 18978 5 1 1 18977
0 18979 7 1 2 37990 18978
0 18980 5 2 1 18979
0 18981 7 1 2 28741 37642
0 18982 5 1 1 18981
0 18983 7 1 2 37998 18982
0 18984 5 1 1 18983
0 18985 7 1 2 34336 18984
0 18986 5 1 1 18985
0 18987 7 1 2 34337 37629
0 18988 5 1 1 18987
0 18989 7 1 2 34200 37974
0 18990 5 1 1 18989
0 18991 7 1 2 18988 18990
0 18992 5 1 1 18991
0 18993 7 1 2 28861 18992
0 18994 5 1 1 18993
0 18995 7 2 2 34338 37729
0 18996 7 1 2 26977 38000
0 18997 5 1 1 18996
0 18998 7 1 2 18994 18997
0 18999 5 1 1 18998
0 19000 7 1 2 28828 18999
0 19001 5 1 1 19000
0 19002 7 1 2 27704 37976
0 19003 5 1 1 19002
0 19004 7 1 2 32797 37868
0 19005 5 1 1 19004
0 19006 7 1 2 19003 19005
0 19007 5 1 1 19006
0 19008 7 1 2 28742 19007
0 19009 5 1 1 19008
0 19010 7 1 2 34015 36481
0 19011 7 1 2 37991 19010
0 19012 5 1 1 19011
0 19013 7 1 2 19009 19012
0 19014 7 1 2 19001 19013
0 19015 7 1 2 18986 19014
0 19016 5 1 1 19015
0 19017 7 1 2 26106 19016
0 19018 5 1 1 19017
0 19019 7 1 2 18974 19018
0 19020 5 1 1 19019
0 19021 7 1 2 27553 30369
0 19022 7 1 2 19020 19021
0 19023 5 1 1 19022
0 19024 7 1 2 18954 19023
0 19025 5 1 1 19024
0 19026 7 1 2 37780 19025
0 19027 5 1 1 19026
0 19028 7 1 2 34687 37959
0 19029 7 1 2 37344 19028
0 19030 7 2 2 27830 37891
0 19031 7 1 2 28792 28592
0 19032 7 1 2 36489 19031
0 19033 7 1 2 38002 19032
0 19034 7 1 2 19029 19033
0 19035 5 1 1 19034
0 19036 7 1 2 19027 19035
0 19037 7 1 2 18798 19036
0 19038 7 1 2 18288 19037
0 19039 5 1 1 19038
0 19040 7 1 2 27483 19039
0 19041 5 1 1 19040
0 19042 7 4 2 23845 28425
0 19043 7 2 2 28365 29376
0 19044 7 1 2 38004 38008
0 19045 5 1 1 19044
0 19046 7 1 2 29310 36747
0 19047 5 1 1 19046
0 19048 7 1 2 19045 19047
0 19049 5 1 1 19048
0 19050 7 2 2 37116 19049
0 19051 5 1 1 38010
0 19052 7 3 2 25093 28278
0 19053 5 1 1 38012
0 19054 7 1 2 28267 19053
0 19055 5 3 1 19054
0 19056 7 1 2 28247 38015
0 19057 5 1 1 19056
0 19058 7 1 2 25094 28331
0 19059 5 1 1 19058
0 19060 7 1 2 19057 19059
0 19061 5 3 1 19060
0 19062 7 1 2 22510 38018
0 19063 5 1 1 19062
0 19064 7 1 2 24506 36213
0 19065 5 1 1 19064
0 19066 7 1 2 19063 19065
0 19067 5 4 1 19066
0 19068 7 1 2 37064 38021
0 19069 5 1 1 19068
0 19070 7 1 2 19051 19069
0 19071 5 2 1 19070
0 19072 7 1 2 29306 38025
0 19073 5 1 1 19072
0 19074 7 2 2 24129 37372
0 19075 7 1 2 22760 38027
0 19076 7 1 2 38022 19075
0 19077 5 1 1 19076
0 19078 7 1 2 19073 19077
0 19079 5 1 1 19078
0 19080 7 1 2 23735 19079
0 19081 5 1 1 19080
0 19082 7 2 2 25717 30258
0 19083 7 1 2 29026 37544
0 19084 5 1 1 19083
0 19085 7 1 2 24709 37300
0 19086 5 1 1 19085
0 19087 7 1 2 19084 19086
0 19088 5 1 1 19087
0 19089 7 1 2 38029 19088
0 19090 7 1 2 37837 19089
0 19091 5 1 1 19090
0 19092 7 1 2 19081 19091
0 19093 5 1 1 19092
0 19094 7 1 2 22860 19093
0 19095 5 1 1 19094
0 19096 7 1 2 37111 38023
0 19097 5 1 1 19096
0 19098 7 1 2 24130 38011
0 19099 5 1 1 19098
0 19100 7 1 2 19097 19099
0 19101 5 1 1 19100
0 19102 7 1 2 36635 19101
0 19103 5 1 1 19102
0 19104 7 1 2 19095 19103
0 19105 5 1 1 19104
0 19106 7 1 2 27005 19105
0 19107 5 1 1 19106
0 19108 7 1 2 31221 37055
0 19109 5 1 1 19108
0 19110 7 1 2 37109 19109
0 19111 5 3 1 19110
0 19112 7 1 2 22761 31146
0 19113 5 1 1 19112
0 19114 7 1 2 30623 32181
0 19115 5 1 1 19114
0 19116 7 1 2 19113 19115
0 19117 5 1 1 19116
0 19118 7 1 2 33724 19117
0 19119 5 1 1 19118
0 19120 7 1 2 34121 36176
0 19121 5 1 1 19120
0 19122 7 1 2 19119 19121
0 19123 5 1 1 19122
0 19124 7 1 2 23736 19123
0 19125 5 1 1 19124
0 19126 7 1 2 34602 37468
0 19127 5 1 1 19126
0 19128 7 1 2 19125 19127
0 19129 5 1 1 19128
0 19130 7 1 2 22511 19129
0 19131 5 1 1 19130
0 19132 7 1 2 27038 33739
0 19133 5 1 1 19132
0 19134 7 1 2 27053 34808
0 19135 5 1 1 19134
0 19136 7 1 2 19133 19135
0 19137 5 1 1 19136
0 19138 7 1 2 22762 19137
0 19139 5 1 1 19138
0 19140 7 1 2 32276 34809
0 19141 5 1 1 19140
0 19142 7 1 2 19139 19141
0 19143 5 2 1 19142
0 19144 7 1 2 23283 33704
0 19145 7 1 2 38034 19144
0 19146 5 1 1 19145
0 19147 7 1 2 19131 19146
0 19148 5 1 1 19147
0 19149 7 1 2 38031 19148
0 19150 5 1 1 19149
0 19151 7 1 2 32195 31932
0 19152 5 1 1 19151
0 19153 7 1 2 34348 35610
0 19154 5 1 1 19153
0 19155 7 1 2 19152 19154
0 19156 5 1 1 19155
0 19157 7 1 2 29437 19156
0 19158 5 1 1 19157
0 19159 7 3 2 25828 26628
0 19160 7 1 2 31772 38036
0 19161 5 1 1 19160
0 19162 7 1 2 27163 19161
0 19163 5 1 1 19162
0 19164 7 1 2 30100 19163
0 19165 5 1 1 19164
0 19166 7 1 2 19158 19165
0 19167 5 1 1 19166
0 19168 7 1 2 22763 19167
0 19169 5 1 1 19168
0 19170 7 1 2 29438 26621
0 19171 5 1 1 19170
0 19172 7 1 2 24915 36886
0 19173 5 1 1 19172
0 19174 7 1 2 19171 19173
0 19175 5 1 1 19174
0 19176 7 1 2 27221 32277
0 19177 7 1 2 19175 19176
0 19178 5 1 1 19177
0 19179 7 1 2 19169 19178
0 19180 5 1 1 19179
0 19181 7 1 2 26272 19180
0 19182 5 1 1 19181
0 19183 7 3 2 26417 30591
0 19184 7 1 2 27222 37117
0 19185 7 1 2 38039 19184
0 19186 7 1 2 34031 19185
0 19187 5 1 1 19186
0 19188 7 1 2 19182 19187
0 19189 5 1 1 19188
0 19190 7 1 2 29690 19189
0 19191 5 1 1 19190
0 19192 7 1 2 25095 37061
0 19193 5 1 1 19192
0 19194 7 1 2 14936 19193
0 19195 5 3 1 19194
0 19196 7 1 2 27993 38042
0 19197 7 1 2 38035 19196
0 19198 5 1 1 19197
0 19199 7 1 2 19191 19198
0 19200 5 1 1 19199
0 19201 7 1 2 24131 19200
0 19202 5 1 1 19201
0 19203 7 1 2 19150 19202
0 19204 5 1 1 19203
0 19205 7 1 2 28170 19204
0 19206 5 1 1 19205
0 19207 7 1 2 38032 37240
0 19208 5 1 1 19207
0 19209 7 1 2 31465 38043
0 19210 5 1 1 19209
0 19211 7 1 2 29439 28426
0 19212 5 1 1 19211
0 19213 7 1 2 23433 26498
0 19214 5 1 1 19213
0 19215 7 1 2 24916 32995
0 19216 7 1 2 19214 19215
0 19217 5 1 1 19216
0 19218 7 1 2 19212 19217
0 19219 5 1 1 19218
0 19220 7 1 2 32333 19219
0 19221 5 1 1 19220
0 19222 7 1 2 19210 19221
0 19223 5 1 1 19222
0 19224 7 1 2 24132 19223
0 19225 5 1 1 19224
0 19226 7 1 2 19208 19225
0 19227 5 1 1 19226
0 19228 7 1 2 26921 30126
0 19229 7 1 2 19227 19228
0 19230 5 1 1 19229
0 19231 7 2 2 30995 34810
0 19232 7 1 2 24507 38045
0 19233 5 1 1 19232
0 19234 7 1 2 32701 29638
0 19235 7 1 2 26929 19234
0 19236 5 1 1 19235
0 19237 7 1 2 19233 19236
0 19238 5 1 1 19237
0 19239 7 1 2 29230 19238
0 19240 5 1 1 19239
0 19241 7 1 2 29241 38046
0 19242 5 1 1 19241
0 19243 7 1 2 19240 19242
0 19244 5 1 1 19243
0 19245 7 1 2 37133 19244
0 19246 5 1 1 19245
0 19247 7 1 2 24791 19246
0 19248 7 1 2 19230 19247
0 19249 7 1 2 19206 19248
0 19250 5 1 1 19249
0 19251 7 4 2 27148 30776
0 19252 7 1 2 38047 37166
0 19253 5 1 1 19252
0 19254 7 1 2 37405 19253
0 19255 5 1 1 19254
0 19256 7 1 2 23284 19255
0 19257 5 1 1 19256
0 19258 7 1 2 31349 37439
0 19259 7 1 2 35429 19258
0 19260 5 1 1 19259
0 19261 7 1 2 19257 19260
0 19262 5 1 1 19261
0 19263 7 1 2 23737 19262
0 19264 5 1 1 19263
0 19265 7 1 2 31848 31310
0 19266 7 1 2 37654 19265
0 19267 5 1 1 19266
0 19268 7 1 2 19264 19267
0 19269 5 1 1 19268
0 19270 7 1 2 22512 19269
0 19271 5 1 1 19270
0 19272 7 1 2 23285 37400
0 19273 5 1 1 19272
0 19274 7 1 2 25240 37407
0 19275 5 1 1 19274
0 19276 7 1 2 24508 19275
0 19277 7 1 2 19273 19276
0 19278 5 1 1 19277
0 19279 7 1 2 19271 19278
0 19280 5 1 1 19279
0 19281 7 1 2 25096 19280
0 19282 5 1 1 19281
0 19283 7 1 2 29769 34596
0 19284 7 1 2 37398 19283
0 19285 5 1 1 19284
0 19286 7 1 2 19282 19285
0 19287 5 1 1 19286
0 19288 7 1 2 32120 19287
0 19289 5 1 1 19288
0 19290 7 1 2 31018 37877
0 19291 5 1 1 19290
0 19292 7 1 2 31611 36637
0 19293 5 1 1 19292
0 19294 7 1 2 19291 19293
0 19295 5 1 1 19294
0 19296 7 1 2 36748 19295
0 19297 5 1 1 19296
0 19298 7 2 2 30985 29424
0 19299 7 1 2 37472 38051
0 19300 5 1 1 19299
0 19301 7 1 2 22513 19300
0 19302 7 1 2 19297 19301
0 19303 5 1 1 19302
0 19304 7 2 2 22764 27157
0 19305 7 1 2 31817 29726
0 19306 5 1 1 19305
0 19307 7 1 2 26273 34603
0 19308 5 1 1 19307
0 19309 7 1 2 19306 19308
0 19310 5 1 1 19309
0 19311 7 1 2 38053 19310
0 19312 5 1 1 19311
0 19313 7 1 2 27788 36286
0 19314 5 1 1 19313
0 19315 7 1 2 26274 38013
0 19316 5 1 1 19315
0 19317 7 1 2 19314 19316
0 19318 5 1 1 19317
0 19319 7 1 2 27182 29746
0 19320 7 1 2 19318 19319
0 19321 5 1 1 19320
0 19322 7 1 2 19312 19321
0 19323 5 1 1 19322
0 19324 7 1 2 26418 19323
0 19325 5 1 1 19324
0 19326 7 1 2 31019 31650
0 19327 5 1 1 19326
0 19328 7 1 2 30986 33740
0 19329 5 1 1 19328
0 19330 7 1 2 19327 19329
0 19331 5 2 1 19330
0 19332 7 1 2 27789 35205
0 19333 7 1 2 38055 19332
0 19334 5 1 1 19333
0 19335 7 1 2 24509 19334
0 19336 7 1 2 19325 19335
0 19337 5 1 1 19336
0 19338 7 1 2 35723 19337
0 19339 7 1 2 19303 19338
0 19340 5 1 1 19339
0 19341 7 2 2 32021 31842
0 19342 7 2 2 37311 38057
0 19343 5 1 1 38059
0 19344 7 1 2 29912 38060
0 19345 7 1 2 34355 19344
0 19346 5 1 1 19345
0 19347 7 1 2 19340 19346
0 19348 7 1 2 19289 19347
0 19349 5 1 1 19348
0 19350 7 1 2 24917 19349
0 19351 5 1 1 19350
0 19352 7 2 2 31174 29624
0 19353 7 1 2 28693 38061
0 19354 5 1 1 19353
0 19355 7 1 2 29879 37065
0 19356 5 1 1 19355
0 19357 7 2 2 19354 19356
0 19358 5 2 1 38063
0 19359 7 1 2 25097 38065
0 19360 5 2 1 19359
0 19361 7 2 2 27526 29844
0 19362 7 1 2 36749 38069
0 19363 5 1 1 19362
0 19364 7 1 2 38067 19363
0 19365 5 1 1 19364
0 19366 7 1 2 27994 38056
0 19367 5 1 1 19366
0 19368 7 1 2 32780 36545
0 19369 7 1 2 35649 19368
0 19370 5 1 1 19369
0 19371 7 1 2 19367 19370
0 19372 5 1 1 19371
0 19373 7 1 2 19365 19372
0 19374 5 1 1 19373
0 19375 7 1 2 29933 34555
0 19376 7 1 2 34597 19375
0 19377 7 1 2 37180 19376
0 19378 5 1 1 19377
0 19379 7 1 2 28427 38070
0 19380 5 1 1 19379
0 19381 7 1 2 38064 19380
0 19382 5 1 1 19381
0 19383 7 1 2 37365 38052
0 19384 7 1 2 19382 19383
0 19385 5 1 1 19384
0 19386 7 1 2 19378 19385
0 19387 7 1 2 19374 19386
0 19388 7 1 2 19351 19387
0 19389 5 1 1 19388
0 19390 7 1 2 28171 19389
0 19391 5 1 1 19390
0 19392 7 2 2 24336 28291
0 19393 7 2 2 37312 38071
0 19394 7 1 2 25643 27415
0 19395 7 1 2 38073 19394
0 19396 5 1 1 19395
0 19397 7 1 2 30078 37444
0 19398 7 1 2 36967 19397
0 19399 5 1 1 19398
0 19400 7 1 2 19396 19399
0 19401 5 1 1 19400
0 19402 7 1 2 24918 19401
0 19403 5 1 1 19402
0 19404 7 2 2 30795 37058
0 19405 5 1 1 38075
0 19406 7 1 2 28263 38076
0 19407 5 1 1 19406
0 19408 7 1 2 19403 19407
0 19409 5 1 1 19408
0 19410 7 1 2 28318 19409
0 19411 5 1 1 19410
0 19412 7 2 2 25926 31175
0 19413 7 1 2 24710 28385
0 19414 7 2 2 38077 19413
0 19415 5 1 1 38079
0 19416 7 1 2 19415 19405
0 19417 5 1 1 19416
0 19418 7 1 2 37814 19417
0 19419 5 1 1 19418
0 19420 7 1 2 19411 19419
0 19421 5 1 1 19420
0 19422 7 1 2 25098 19421
0 19423 5 1 1 19422
0 19424 7 1 2 24214 30798
0 19425 7 1 2 31382 19424
0 19426 7 1 2 36750 19425
0 19427 5 1 1 19426
0 19428 7 1 2 19423 19427
0 19429 5 1 1 19428
0 19430 7 1 2 24510 19429
0 19431 5 1 1 19430
0 19432 7 1 2 30799 37181
0 19433 5 1 1 19432
0 19434 7 2 2 32022 30723
0 19435 7 1 2 38078 38081
0 19436 5 1 1 19435
0 19437 7 1 2 19433 19436
0 19438 5 1 1 19437
0 19439 7 1 2 31392 19438
0 19440 5 1 1 19439
0 19441 7 1 2 25718 19440
0 19442 7 1 2 19431 19441
0 19443 5 1 1 19442
0 19444 7 1 2 30796 38026
0 19445 5 1 1 19444
0 19446 7 1 2 38024 38080
0 19447 5 1 1 19446
0 19448 7 1 2 23738 19447
0 19449 7 1 2 19445 19448
0 19450 5 1 1 19449
0 19451 7 1 2 26922 19450
0 19452 7 1 2 19443 19451
0 19453 5 1 1 19452
0 19454 7 1 2 31052 27662
0 19455 7 1 2 36875 19454
0 19456 5 1 1 19455
0 19457 7 1 2 791 28777
0 19458 7 1 2 29344 1696
0 19459 7 1 2 19457 19458
0 19460 7 1 2 36781 19459
0 19461 5 1 1 19460
0 19462 7 1 2 19456 19461
0 19463 5 1 1 19462
0 19464 7 1 2 23434 19463
0 19465 5 1 1 19464
0 19466 7 1 2 28775 30259
0 19467 7 1 2 37308 19466
0 19468 5 1 1 19467
0 19469 7 1 2 19465 19468
0 19470 5 1 1 19469
0 19471 7 1 2 31820 30144
0 19472 7 1 2 19470 19471
0 19473 5 1 1 19472
0 19474 7 1 2 22861 19473
0 19475 7 1 2 19453 19474
0 19476 7 1 2 19391 19475
0 19477 5 1 1 19476
0 19478 7 1 2 19250 19477
0 19479 5 1 1 19478
0 19480 7 1 2 19107 19479
0 19481 5 1 1 19480
0 19482 7 1 2 33404 19481
0 19483 5 1 1 19482
0 19484 7 1 2 22862 37585
0 19485 5 1 1 19484
0 19486 7 1 2 26874 27534
0 19487 5 1 1 19486
0 19488 7 1 2 19485 19487
0 19489 5 1 1 19488
0 19490 7 1 2 23364 19489
0 19491 5 1 1 19490
0 19492 7 1 2 35816 30584
0 19493 7 1 2 33509 19492
0 19494 5 1 1 19493
0 19495 7 1 2 19491 19494
0 19496 5 1 1 19495
0 19497 7 1 2 23846 19496
0 19498 5 1 1 19497
0 19499 7 2 2 34477 37078
0 19500 7 2 2 24792 27535
0 19501 5 1 1 38085
0 19502 7 1 2 29961 35087
0 19503 5 1 1 19502
0 19504 7 1 2 19501 19503
0 19505 5 4 1 19504
0 19506 7 1 2 38083 38087
0 19507 5 1 1 19506
0 19508 7 1 2 19498 19507
0 19509 5 1 1 19508
0 19510 7 1 2 32121 19509
0 19511 5 1 1 19510
0 19512 7 1 2 22863 37589
0 19513 5 1 1 19512
0 19514 7 1 2 26852 27536
0 19515 5 1 1 19514
0 19516 7 1 2 19513 19515
0 19517 5 2 1 19516
0 19518 7 2 2 30987 29364
0 19519 5 1 1 38093
0 19520 7 1 2 32702 34573
0 19521 5 1 1 19520
0 19522 7 1 2 19519 19521
0 19523 5 1 1 19522
0 19524 7 1 2 23952 19523
0 19525 7 1 2 38091 19524
0 19526 5 1 1 19525
0 19527 7 1 2 19511 19526
0 19528 5 1 1 19527
0 19529 7 1 2 31237 19528
0 19530 5 1 1 19529
0 19531 7 1 2 22652 19530
0 19532 5 1 1 19531
0 19533 7 1 2 32417 37079
0 19534 5 1 1 19533
0 19535 7 1 2 35787 19534
0 19536 5 1 1 19535
0 19537 7 1 2 38088 19536
0 19538 5 1 1 19537
0 19539 7 2 2 34954 30471
0 19540 7 1 2 29365 38095
0 19541 7 1 2 34716 19540
0 19542 5 1 1 19541
0 19543 7 1 2 19538 19542
0 19544 5 1 1 19543
0 19545 7 1 2 28386 19544
0 19546 5 1 1 19545
0 19547 7 1 2 34349 27422
0 19548 7 1 2 37559 19547
0 19549 5 1 1 19548
0 19550 7 1 2 19546 19549
0 19551 5 1 1 19550
0 19552 7 1 2 22765 19551
0 19553 5 1 1 19552
0 19554 7 1 2 35791 30288
0 19555 5 1 1 19554
0 19556 7 1 2 31384 30963
0 19557 5 1 1 19556
0 19558 7 1 2 19555 19557
0 19559 5 1 1 19558
0 19560 7 1 2 22864 19559
0 19561 5 1 1 19560
0 19562 7 1 2 26923 33392
0 19563 7 1 2 27537 19562
0 19564 5 1 1 19563
0 19565 7 1 2 19561 19564
0 19566 5 1 1 19565
0 19567 7 1 2 38082 19566
0 19568 5 1 1 19567
0 19569 7 1 2 19553 19568
0 19570 5 1 1 19569
0 19571 7 1 2 25927 19570
0 19572 5 1 1 19571
0 19573 7 1 2 30384 36989
0 19574 5 1 1 19573
0 19575 7 1 2 16958 19574
0 19576 5 1 1 19575
0 19577 7 1 2 22865 19576
0 19578 5 1 1 19577
0 19579 7 1 2 28748 38086
0 19580 5 1 1 19579
0 19581 7 1 2 19578 19580
0 19582 5 1 1 19581
0 19583 7 2 2 27223 32023
0 19584 7 1 2 32122 29625
0 19585 7 1 2 38097 19584
0 19586 7 1 2 19582 19585
0 19587 5 1 1 19586
0 19588 7 1 2 24616 19587
0 19589 7 1 2 19572 19588
0 19590 5 1 1 19589
0 19591 7 1 2 19532 19590
0 19592 5 1 1 19591
0 19593 7 1 2 31430 37561
0 19594 5 1 1 19593
0 19595 7 2 2 22653 27243
0 19596 5 1 1 38099
0 19597 7 1 2 33849 33725
0 19598 5 1 1 19597
0 19599 7 1 2 19596 19598
0 19600 5 3 1 19599
0 19601 7 1 2 28387 38101
0 19602 7 1 2 38092 19601
0 19603 5 1 1 19602
0 19604 7 1 2 19594 19603
0 19605 5 1 1 19604
0 19606 7 1 2 32255 19605
0 19607 5 1 1 19606
0 19608 7 1 2 34516 38037
0 19609 5 1 1 19608
0 19610 7 1 2 26521 38094
0 19611 5 1 1 19610
0 19612 7 1 2 19609 19611
0 19613 5 1 1 19612
0 19614 7 1 2 22654 19613
0 19615 5 1 1 19614
0 19616 7 1 2 35466 38038
0 19617 5 1 1 19616
0 19618 7 1 2 19615 19617
0 19619 5 1 1 19618
0 19620 7 1 2 26275 19619
0 19621 5 1 1 19620
0 19622 7 1 2 25829 38040
0 19623 7 1 2 35472 19622
0 19624 5 1 1 19623
0 19625 7 1 2 19621 19624
0 19626 5 1 1 19625
0 19627 7 1 2 23953 19626
0 19628 5 1 1 19627
0 19629 7 1 2 32910 37425
0 19630 5 1 1 19629
0 19631 7 1 2 19628 19630
0 19632 5 1 1 19631
0 19633 7 1 2 32935 19632
0 19634 5 1 1 19633
0 19635 7 1 2 36782 37925
0 19636 5 1 1 19635
0 19637 7 1 2 28248 37348
0 19638 5 1 1 19637
0 19639 7 1 2 16110 19638
0 19640 5 1 1 19639
0 19641 7 1 2 26276 19640
0 19642 5 1 1 19641
0 19643 7 1 2 28897 37841
0 19644 5 1 1 19643
0 19645 7 1 2 19642 19644
0 19646 5 2 1 19645
0 19647 7 1 2 32882 38104
0 19648 5 1 1 19647
0 19649 7 1 2 19636 19648
0 19650 5 1 1 19649
0 19651 7 1 2 32123 19650
0 19652 5 1 1 19651
0 19653 7 1 2 22866 34580
0 19654 7 1 2 36853 19653
0 19655 7 1 2 36668 19654
0 19656 5 1 1 19655
0 19657 7 1 2 19652 19656
0 19658 7 1 2 19634 19657
0 19659 5 1 1 19658
0 19660 7 1 2 37118 19659
0 19661 5 1 1 19660
0 19662 7 1 2 19607 19661
0 19663 7 1 2 19592 19662
0 19664 5 1 1 19663
0 19665 7 1 2 28951 19664
0 19666 5 1 1 19665
0 19667 7 1 2 30082 29739
0 19668 5 1 1 19667
0 19669 7 1 2 26522 30407
0 19670 7 1 2 32204 19669
0 19671 5 1 1 19670
0 19672 7 1 2 19668 19671
0 19673 5 1 1 19672
0 19674 7 1 2 31020 26871
0 19675 7 1 2 19673 19674
0 19676 5 1 1 19675
0 19677 7 1 2 27295 28778
0 19678 5 1 1 19677
0 19679 7 1 2 2080 27706
0 19680 5 1 1 19679
0 19681 7 2 2 19678 19680
0 19682 7 1 2 32836 38106
0 19683 5 1 1 19682
0 19684 7 1 2 32752 35634
0 19685 5 1 1 19684
0 19686 7 1 2 27026 35357
0 19687 7 1 2 29907 19686
0 19688 5 1 1 19687
0 19689 7 1 2 19685 19688
0 19690 7 1 2 19683 19689
0 19691 5 1 1 19690
0 19692 7 1 2 26523 37119
0 19693 7 1 2 19691 19692
0 19694 5 1 1 19693
0 19695 7 1 2 19676 19694
0 19696 5 1 1 19695
0 19697 7 1 2 26277 19696
0 19698 5 1 1 19697
0 19699 7 1 2 23954 30944
0 19700 5 1 1 19699
0 19701 7 1 2 10976 19700
0 19702 5 1 1 19701
0 19703 7 1 2 25324 19702
0 19704 5 1 1 19703
0 19705 7 1 2 28878 31893
0 19706 5 1 1 19705
0 19707 7 1 2 19704 19706
0 19708 5 2 1 19707
0 19709 7 1 2 38096 38108
0 19710 5 1 1 19709
0 19711 7 1 2 25325 32500
0 19712 5 1 1 19711
0 19713 7 1 2 23365 16181
0 19714 5 1 1 19713
0 19715 7 1 2 38089 19714
0 19716 7 1 2 19712 19715
0 19717 5 1 1 19716
0 19718 7 1 2 19710 19717
0 19719 5 1 1 19718
0 19720 7 1 2 28388 19719
0 19721 5 1 1 19720
0 19722 7 1 2 19698 19721
0 19723 5 1 1 19722
0 19724 7 1 2 24617 19723
0 19725 5 1 1 19724
0 19726 7 3 2 37120 36854
0 19727 5 1 1 38110
0 19728 7 1 2 37500 38111
0 19729 5 1 1 19728
0 19730 7 1 2 34032 38090
0 19731 5 1 1 19730
0 19732 7 3 2 24711 34955
0 19733 7 1 2 27054 30472
0 19734 7 1 2 38113 19733
0 19735 5 1 1 19734
0 19736 7 1 2 19731 19735
0 19737 5 1 1 19736
0 19738 7 1 2 28389 19737
0 19739 5 1 1 19738
0 19740 7 1 2 19729 19739
0 19741 5 1 1 19740
0 19742 7 1 2 30887 19741
0 19743 5 1 1 19742
0 19744 7 1 2 19725 19743
0 19745 5 1 1 19744
0 19746 7 1 2 23847 28960
0 19747 7 1 2 19745 19746
0 19748 5 1 1 19747
0 19749 7 1 2 19666 19748
0 19750 5 1 1 19749
0 19751 7 1 2 23739 28223
0 19752 7 1 2 33408 19751
0 19753 7 1 2 19750 19752
0 19754 5 1 1 19753
0 19755 7 1 2 19483 19754
0 19756 5 1 1 19755
0 19757 7 1 2 36438 16523
0 19758 5 2 1 19757
0 19759 7 1 2 32065 38116
0 19760 7 1 2 19756 19759
0 19761 5 1 1 19760
0 19762 7 1 2 27224 37080
0 19763 5 1 1 19762
0 19764 7 1 2 27251 19763
0 19765 5 2 1 19764
0 19766 7 1 2 38118 38033
0 19767 5 1 1 19766
0 19768 7 2 2 27441 38005
0 19769 5 1 1 38120
0 19770 7 1 2 29440 38121
0 19771 5 1 1 19770
0 19772 7 1 2 27111 38044
0 19773 5 1 1 19772
0 19774 7 1 2 19771 19773
0 19775 5 1 1 19774
0 19776 7 1 2 24133 19775
0 19777 5 1 1 19776
0 19778 7 1 2 19767 19777
0 19779 5 1 1 19778
0 19780 7 1 2 29691 19779
0 19781 5 1 1 19780
0 19782 7 1 2 27995 37764
0 19783 7 1 2 37134 19782
0 19784 5 1 1 19783
0 19785 7 1 2 19781 19784
0 19786 5 1 1 19785
0 19787 7 1 2 34438 19786
0 19788 5 1 1 19787
0 19789 7 1 2 35360 37096
0 19790 5 1 1 19789
0 19791 7 1 2 24040 34484
0 19792 7 1 2 34740 19791
0 19793 7 1 2 26629 19792
0 19794 5 1 1 19793
0 19795 7 1 2 19790 19794
0 19796 5 1 1 19795
0 19797 7 1 2 22514 19796
0 19798 5 1 1 19797
0 19799 7 1 2 27707 605
0 19800 5 1 1 19799
0 19801 7 1 2 7280 14043
0 19802 7 2 2 19800 19801
0 19803 7 1 2 31106 26630
0 19804 7 1 2 38122 19803
0 19805 5 1 1 19804
0 19806 7 1 2 19798 19805
0 19807 5 1 1 19806
0 19808 7 1 2 26278 19807
0 19809 5 1 1 19808
0 19810 7 1 2 24511 38123
0 19811 5 1 1 19810
0 19812 7 1 2 28066 30205
0 19813 5 1 1 19812
0 19814 7 1 2 19811 19813
0 19815 5 3 1 19814
0 19816 7 1 2 25719 38041
0 19817 7 1 2 38124 19816
0 19818 5 1 1 19817
0 19819 7 1 2 19809 19818
0 19820 5 1 1 19819
0 19821 7 1 2 24919 19820
0 19822 5 1 1 19821
0 19823 7 2 2 29626 38125
0 19824 7 2 2 32024 30552
0 19825 7 1 2 38127 38129
0 19826 5 1 1 19825
0 19827 7 1 2 19822 19826
0 19828 5 1 1 19827
0 19829 7 1 2 23955 19828
0 19830 5 1 1 19829
0 19831 7 1 2 26499 34432
0 19832 5 1 1 19831
0 19833 7 1 2 32375 29924
0 19834 7 1 2 34439 19833
0 19835 7 1 2 19832 19834
0 19836 5 1 1 19835
0 19837 7 1 2 19830 19836
0 19838 5 1 1 19837
0 19839 7 1 2 26196 19838
0 19840 5 1 1 19839
0 19841 7 1 2 30140 29441
0 19842 7 1 2 36783 19841
0 19843 7 1 2 38126 19842
0 19844 5 1 1 19843
0 19845 7 1 2 19840 19844
0 19846 5 1 1 19845
0 19847 7 1 2 24134 19846
0 19848 5 1 1 19847
0 19849 7 1 2 32383 31849
0 19850 7 1 2 37600 19849
0 19851 7 1 2 38128 19850
0 19852 5 1 1 19851
0 19853 7 1 2 19848 19852
0 19854 5 1 1 19853
0 19855 7 1 2 23366 19854
0 19856 5 1 1 19855
0 19857 7 1 2 29777 32678
0 19858 7 1 2 36671 28461
0 19859 7 1 2 19857 19858
0 19860 5 1 1 19859
0 19861 7 1 2 19856 19860
0 19862 5 1 1 19861
0 19863 7 1 2 23848 19862
0 19864 5 1 1 19863
0 19865 7 1 2 19788 19864
0 19866 5 1 1 19865
0 19867 7 1 2 22867 19866
0 19868 5 1 1 19867
0 19869 7 5 2 26197 36784
0 19870 5 1 1 38131
0 19871 7 1 2 29880 38132
0 19872 5 1 1 19871
0 19873 7 1 2 19343 19872
0 19874 5 1 1 19873
0 19875 7 1 2 24920 19874
0 19876 5 1 1 19875
0 19877 7 1 2 35718 37182
0 19878 5 1 1 19877
0 19879 7 1 2 19876 19878
0 19880 5 1 1 19879
0 19881 7 1 2 24712 19880
0 19882 5 1 1 19881
0 19883 7 1 2 35614 33629
0 19884 7 1 2 38062 19883
0 19885 5 1 1 19884
0 19886 7 1 2 19882 19885
0 19887 5 1 1 19886
0 19888 7 1 2 22655 19887
0 19889 5 1 1 19888
0 19890 7 1 2 30152 37191
0 19891 5 1 1 19890
0 19892 7 1 2 19889 19891
0 19893 5 1 1 19892
0 19894 7 1 2 37765 19893
0 19895 5 1 1 19894
0 19896 7 1 2 29881 37130
0 19897 5 1 1 19896
0 19898 7 1 2 38068 19897
0 19899 5 1 1 19898
0 19900 7 1 2 28449 29747
0 19901 7 1 2 19899 19900
0 19902 5 1 1 19901
0 19903 7 1 2 30473 29526
0 19904 7 1 2 36230 19903
0 19905 7 1 2 36785 19904
0 19906 5 1 1 19905
0 19907 7 1 2 19902 19906
0 19908 5 1 1 19907
0 19909 7 1 2 23367 19908
0 19910 5 1 1 19909
0 19911 7 2 2 26978 37301
0 19912 5 1 1 38136
0 19913 7 1 2 23849 28762
0 19914 7 1 2 38030 19913
0 19915 7 1 2 38137 19914
0 19916 5 1 1 19915
0 19917 7 1 2 19910 19916
0 19918 5 1 1 19917
0 19919 7 1 2 24618 19918
0 19920 5 1 1 19919
0 19921 7 1 2 19895 19920
0 19922 5 1 1 19921
0 19923 7 1 2 27996 19922
0 19924 5 1 1 19923
0 19925 7 2 2 28214 30457
0 19926 7 1 2 38119 38066
0 19927 5 1 1 19926
0 19928 7 1 2 27228 36751
0 19929 5 1 1 19928
0 19930 7 1 2 19769 19929
0 19931 5 1 1 19930
0 19932 7 1 2 29882 37121
0 19933 7 1 2 19931 19932
0 19934 5 1 1 19933
0 19935 7 1 2 19927 19934
0 19936 5 1 1 19935
0 19937 7 1 2 38138 19936
0 19938 5 1 1 19937
0 19939 7 1 2 24713 19938
0 19940 5 1 1 19939
0 19941 7 1 2 27027 36786
0 19942 5 1 1 19941
0 19943 7 1 2 27289 36855
0 19944 5 1 1 19943
0 19945 7 1 2 19942 19944
0 19946 5 1 1 19945
0 19947 7 1 2 37122 19946
0 19948 5 1 1 19947
0 19949 7 2 2 29338 28390
0 19950 5 1 1 38140
0 19951 7 1 2 34105 38141
0 19952 5 1 1 19951
0 19953 7 1 2 19948 19952
0 19954 5 1 1 19953
0 19955 7 1 2 30344 19954
0 19956 5 1 1 19955
0 19957 7 1 2 30385 37162
0 19958 5 1 1 19957
0 19959 7 1 2 19956 19958
0 19960 5 1 1 19959
0 19961 7 1 2 23850 19960
0 19962 5 1 1 19961
0 19963 7 1 2 38084 38028
0 19964 5 1 1 19963
0 19965 7 1 2 19962 19964
0 19966 5 1 1 19965
0 19967 7 1 2 22656 19966
0 19968 5 1 1 19967
0 19969 7 1 2 27261 36883
0 19970 7 1 2 37198 19969
0 19971 5 1 1 19970
0 19972 7 1 2 19968 19971
0 19973 5 1 1 19972
0 19974 7 1 2 29692 19973
0 19975 5 1 1 19974
0 19976 7 1 2 35616 37160
0 19977 5 1 1 19976
0 19978 7 1 2 27400 37302
0 19979 5 1 1 19978
0 19980 7 1 2 19977 19979
0 19981 5 1 1 19980
0 19982 7 1 2 24921 27262
0 19983 7 1 2 19981 19982
0 19984 5 1 1 19983
0 19985 7 1 2 28911 37893
0 19986 7 1 2 37059 19985
0 19987 5 1 1 19986
0 19988 7 1 2 19984 19987
0 19989 5 1 1 19988
0 19990 7 1 2 25099 19989
0 19991 5 1 1 19990
0 19992 7 1 2 28450 31094
0 19993 7 1 2 36383 30674
0 19994 7 1 2 19992 19993
0 19995 7 1 2 37004 19994
0 19996 5 1 1 19995
0 19997 7 1 2 19991 19996
0 19998 5 1 1 19997
0 19999 7 1 2 29700 19998
0 20000 5 1 1 19999
0 20001 7 1 2 22766 20000
0 20002 7 1 2 19975 20001
0 20003 5 1 1 20002
0 20004 7 1 2 19940 20003
0 20005 5 1 1 20004
0 20006 7 1 2 19924 20005
0 20007 5 1 1 20006
0 20008 7 1 2 24793 20007
0 20009 5 1 1 20008
0 20010 7 2 2 29627 38016
0 20011 7 1 2 28408 38142
0 20012 5 1 1 20011
0 20013 7 1 2 35902 32996
0 20014 7 1 2 37090 20013
0 20015 5 1 1 20014
0 20016 7 1 2 20012 20015
0 20017 5 1 1 20016
0 20018 7 1 2 25644 20017
0 20019 5 1 1 20018
0 20020 7 1 2 23155 26665
0 20021 5 1 1 20020
0 20022 7 1 2 30569 37440
0 20023 7 2 2 20021 20022
0 20024 7 2 2 24794 26198
0 20025 7 1 2 25241 38146
0 20026 7 1 2 38144 20025
0 20027 5 1 1 20026
0 20028 7 1 2 20019 20027
0 20029 5 1 1 20028
0 20030 7 1 2 24922 20029
0 20031 5 1 1 20030
0 20032 7 2 2 25830 37183
0 20033 7 1 2 25242 35030
0 20034 7 1 2 38148 20033
0 20035 5 1 1 20034
0 20036 7 1 2 20031 20035
0 20037 5 1 1 20036
0 20038 7 1 2 37152 20037
0 20039 5 1 1 20038
0 20040 7 1 2 30528 36466
0 20041 7 1 2 37804 20040
0 20042 5 1 1 20041
0 20043 7 1 2 24041 35059
0 20044 7 1 2 28920 29628
0 20045 7 1 2 20043 20044
0 20046 7 1 2 31623 20045
0 20047 5 1 1 20046
0 20048 7 1 2 20042 20047
0 20049 5 1 1 20048
0 20050 7 1 2 25100 20049
0 20051 5 1 1 20050
0 20052 7 1 2 28264 36856
0 20053 5 1 1 20052
0 20054 7 1 2 28279 36752
0 20055 5 1 1 20054
0 20056 7 1 2 20053 20055
0 20057 5 1 1 20056
0 20058 7 1 2 23740 32364
0 20059 7 1 2 32011 20058
0 20060 7 1 2 20057 20059
0 20061 5 1 1 20060
0 20062 7 1 2 20051 20061
0 20063 5 1 1 20062
0 20064 7 1 2 24215 20063
0 20065 5 1 1 20064
0 20066 7 1 2 22980 38143
0 20067 5 1 1 20066
0 20068 7 1 2 31823 36089
0 20069 5 1 1 20068
0 20070 7 1 2 20067 20069
0 20071 5 1 1 20070
0 20072 7 1 2 25645 20071
0 20073 5 1 1 20072
0 20074 7 1 2 35286 38145
0 20075 5 1 1 20074
0 20076 7 1 2 20073 20075
0 20077 5 1 1 20076
0 20078 7 1 2 23741 26199
0 20079 7 1 2 37203 20078
0 20080 7 1 2 20077 20079
0 20081 5 1 1 20080
0 20082 7 1 2 20065 20081
0 20083 5 1 1 20082
0 20084 7 1 2 24135 20083
0 20085 5 1 1 20084
0 20086 7 1 2 22515 20085
0 20087 7 1 2 20039 20086
0 20088 5 1 1 20087
0 20089 7 1 2 34427 28921
0 20090 7 1 2 38074 20089
0 20091 5 1 1 20090
0 20092 7 1 2 29403 37243
0 20093 5 1 1 20092
0 20094 7 1 2 37853 20093
0 20095 5 1 1 20094
0 20096 7 1 2 22657 23644
0 20097 7 1 2 35430 20096
0 20098 7 1 2 20095 20097
0 20099 5 1 1 20098
0 20100 7 1 2 20091 20099
0 20101 5 1 1 20100
0 20102 7 1 2 25101 20101
0 20103 5 1 1 20102
0 20104 7 2 2 29727 37395
0 20105 7 1 2 30345 34673
0 20106 7 1 2 38150 20105
0 20107 5 1 1 20106
0 20108 7 1 2 20103 20107
0 20109 5 1 1 20108
0 20110 7 1 2 24923 20109
0 20111 5 1 1 20110
0 20112 7 1 2 36384 37849
0 20113 7 1 2 37192 20112
0 20114 5 1 1 20113
0 20115 7 1 2 20111 20114
0 20116 5 1 1 20115
0 20117 7 1 2 24795 20116
0 20118 5 1 1 20117
0 20119 7 1 2 32012 37850
0 20120 7 1 2 37136 20119
0 20121 5 1 1 20120
0 20122 7 1 2 24512 20121
0 20123 7 1 2 20118 20122
0 20124 5 1 1 20123
0 20125 7 1 2 22767 20124
0 20126 7 1 2 20088 20125
0 20127 5 1 1 20126
0 20128 7 1 2 32519 37199
0 20129 5 1 1 20128
0 20130 7 1 2 37413 20129
0 20131 5 1 1 20130
0 20132 7 1 2 24042 20131
0 20133 5 1 1 20132
0 20134 7 2 2 24796 37409
0 20135 7 1 2 30260 38152
0 20136 5 1 1 20135
0 20137 7 1 2 20133 20136
0 20138 5 1 1 20137
0 20139 7 1 2 28067 31614
0 20140 7 1 2 20138 20139
0 20141 5 1 1 20140
0 20142 7 1 2 20127 20141
0 20143 5 1 1 20142
0 20144 7 1 2 27326 20143
0 20145 5 1 1 20144
0 20146 7 1 2 33405 20145
0 20147 7 1 2 20009 20146
0 20148 7 1 2 19868 20147
0 20149 5 1 1 20148
0 20150 7 1 2 22868 27538
0 20151 5 2 1 20150
0 20152 7 1 2 30289 33254
0 20153 5 1 1 20152
0 20154 7 1 2 38154 20153
0 20155 5 1 1 20154
0 20156 7 1 2 37297 20155
0 20157 5 1 1 20156
0 20158 7 1 2 32196 33255
0 20159 7 1 2 31176 20158
0 20160 5 1 1 20159
0 20161 7 1 2 20157 20160
0 20162 5 2 1 20161
0 20163 7 1 2 28391 38156
0 20164 5 1 1 20163
0 20165 7 1 2 37565 20164
0 20166 5 1 1 20165
0 20167 7 1 2 22768 20166
0 20168 5 1 1 20167
0 20169 7 1 2 24797 30290
0 20170 5 1 1 20169
0 20171 7 1 2 38155 20170
0 20172 5 4 1 20171
0 20173 7 1 2 24043 38158
0 20174 5 1 1 20173
0 20175 7 1 2 24798 32262
0 20176 5 1 1 20175
0 20177 7 1 2 20174 20176
0 20178 5 2 1 20177
0 20179 7 2 2 23956 32703
0 20180 7 1 2 25102 28392
0 20181 7 1 2 38164 20180
0 20182 7 1 2 38162 20181
0 20183 5 1 1 20182
0 20184 7 1 2 20168 20183
0 20185 5 1 1 20184
0 20186 7 1 2 28172 20185
0 20187 5 1 1 20186
0 20188 7 1 2 38165 36986
0 20189 5 1 1 20188
0 20190 7 1 2 35132 38048
0 20191 5 1 1 20190
0 20192 7 1 2 20189 20191
0 20193 5 1 1 20192
0 20194 7 2 2 28173 20193
0 20195 5 1 1 38166
0 20196 7 1 2 36787 38167
0 20197 5 1 1 20196
0 20198 7 1 2 37971 38105
0 20199 5 1 1 20198
0 20200 7 1 2 20197 20199
0 20201 5 1 1 20200
0 20202 7 1 2 37123 20201
0 20203 5 1 1 20202
0 20204 7 1 2 32811 38159
0 20205 5 1 1 20204
0 20206 7 2 2 32592 35060
0 20207 7 1 2 30754 38168
0 20208 5 1 1 20207
0 20209 7 1 2 20205 20208
0 20210 5 1 1 20209
0 20211 7 1 2 4552 16120
0 20212 5 1 1 20211
0 20213 7 1 2 31238 20212
0 20214 7 1 2 20210 20213
0 20215 5 1 1 20214
0 20216 7 1 2 20203 20215
0 20217 7 1 2 20187 20216
0 20218 5 1 1 20217
0 20219 7 1 2 24513 20218
0 20220 5 1 1 20219
0 20221 7 1 2 27932 20220
0 20222 5 1 1 20221
0 20223 7 1 2 24619 38107
0 20224 5 1 1 20223
0 20225 7 1 2 30438 34434
0 20226 5 1 1 20225
0 20227 7 1 2 20224 20226
0 20228 5 3 1 20227
0 20229 7 1 2 38160 38170
0 20230 5 1 1 20229
0 20231 7 1 2 29962 38169
0 20232 7 1 2 30899 20231
0 20233 5 1 1 20232
0 20234 7 1 2 20230 20233
0 20235 5 1 1 20234
0 20236 7 1 2 28393 20235
0 20237 5 1 1 20236
0 20238 7 1 2 32560 38112
0 20239 7 1 2 38171 20238
0 20240 5 1 1 20239
0 20241 7 1 2 20237 20240
0 20242 5 1 1 20241
0 20243 7 1 2 23851 20242
0 20244 5 1 1 20243
0 20245 7 1 2 28961 20244
0 20246 5 1 1 20245
0 20247 7 1 2 23742 20246
0 20248 7 1 2 20222 20247
0 20249 5 1 1 20248
0 20250 7 1 2 33409 20249
0 20251 5 1 1 20250
0 20252 7 1 2 26842 37008
0 20253 5 1 1 20252
0 20254 7 1 2 25390 36798
0 20255 5 1 1 20254
0 20256 7 1 2 20253 20255
0 20257 5 2 1 20256
0 20258 7 1 2 32066 38173
0 20259 7 1 2 20251 20258
0 20260 7 1 2 20149 20259
0 20261 5 1 1 20260
0 20262 7 1 2 37051 15487
0 20263 5 1 1 20262
0 20264 7 2 2 33705 34681
0 20265 7 2 2 34069 38175
0 20266 7 1 2 27137 35362
0 20267 5 1 1 20266
0 20268 7 1 2 27090 35368
0 20269 5 1 1 20268
0 20270 7 1 2 20267 20269
0 20271 5 1 1 20270
0 20272 7 1 2 38177 20271
0 20273 5 1 1 20272
0 20274 7 3 2 33575 29728
0 20275 7 2 2 28249 38179
0 20276 7 1 2 27006 38182
0 20277 5 1 1 20276
0 20278 7 3 2 25103 29590
0 20279 7 2 2 23594 35278
0 20280 7 1 2 36608 38187
0 20281 7 1 2 38184 20280
0 20282 5 1 1 20281
0 20283 7 1 2 20277 20282
0 20284 5 1 1 20283
0 20285 7 1 2 27138 20284
0 20286 5 1 1 20285
0 20287 7 1 2 31566 37529
0 20288 5 1 1 20287
0 20289 7 1 2 26531 31555
0 20290 7 2 2 23595 34682
0 20291 7 1 2 31549 38189
0 20292 7 1 2 20289 20291
0 20293 5 1 1 20292
0 20294 7 1 2 20288 20293
0 20295 5 1 1 20294
0 20296 7 1 2 26924 20295
0 20297 5 1 1 20296
0 20298 7 1 2 34769 37505
0 20299 7 1 2 28047 20298
0 20300 5 1 1 20299
0 20301 7 1 2 20297 20300
0 20302 7 1 2 20286 20301
0 20303 5 1 1 20302
0 20304 7 1 2 22516 20303
0 20305 5 1 1 20304
0 20306 7 1 2 20273 20305
0 20307 5 1 1 20306
0 20308 7 1 2 23566 20307
0 20309 5 1 1 20308
0 20310 7 1 2 34033 29264
0 20311 5 1 1 20310
0 20312 7 2 2 32891 37369
0 20313 5 1 1 38191
0 20314 7 1 2 24514 38192
0 20315 5 1 1 20314
0 20316 7 1 2 20311 20315
0 20317 5 1 1 20316
0 20318 7 1 2 29018 34683
0 20319 7 1 2 34847 20318
0 20320 7 1 2 20317 20319
0 20321 5 1 1 20320
0 20322 7 1 2 20309 20321
0 20323 5 1 1 20322
0 20324 7 1 2 23852 20323
0 20325 5 1 1 20324
0 20326 7 4 2 29404 37236
0 20327 7 1 2 34034 30900
0 20328 5 1 1 20327
0 20329 7 1 2 26983 35549
0 20330 5 1 1 20329
0 20331 7 1 2 20328 20330
0 20332 5 3 1 20331
0 20333 7 1 2 24799 38117
0 20334 5 1 1 20333
0 20335 7 1 2 28968 37009
0 20336 5 1 1 20335
0 20337 7 1 2 20334 20336
0 20338 5 1 1 20337
0 20339 7 1 2 38197 20338
0 20340 5 1 1 20339
0 20341 7 1 2 24620 38109
0 20342 5 1 1 20341
0 20343 7 1 2 31128 35463
0 20344 5 1 1 20343
0 20345 7 1 2 20342 20344
0 20346 5 3 1 20345
0 20347 7 1 2 34070 36068
0 20348 7 1 2 38200 20347
0 20349 5 1 1 20348
0 20350 7 1 2 20340 20349
0 20351 5 1 1 20350
0 20352 7 1 2 38193 20351
0 20353 5 1 1 20352
0 20354 7 1 2 20325 20353
0 20355 5 1 1 20354
0 20356 7 1 2 25159 20355
0 20357 5 1 1 20356
0 20358 7 2 2 23853 33576
0 20359 7 2 2 36518 38203
0 20360 7 1 2 29132 35635
0 20361 5 1 1 20360
0 20362 7 1 2 28862 37820
0 20363 5 1 1 20362
0 20364 7 1 2 20361 20363
0 20365 5 4 1 20364
0 20366 7 1 2 28829 38207
0 20367 5 1 1 20366
0 20368 7 1 2 37999 20367
0 20369 7 1 2 37650 20368
0 20370 5 4 1 20369
0 20371 7 1 2 38205 38211
0 20372 5 1 1 20371
0 20373 7 1 2 20357 20372
0 20374 5 1 1 20373
0 20375 7 1 2 24924 20374
0 20376 5 1 1 20375
0 20377 7 2 2 37530 37946
0 20378 7 2 2 26542 38215
0 20379 7 1 2 34254 34773
0 20380 5 1 1 20379
0 20381 7 1 2 22658 34745
0 20382 5 1 1 20381
0 20383 7 1 2 33967 31351
0 20384 5 1 1 20383
0 20385 7 1 2 20382 20384
0 20386 5 1 1 20385
0 20387 7 1 2 22517 20386
0 20388 5 1 1 20387
0 20389 7 1 2 31588 33991
0 20390 5 1 1 20389
0 20391 7 1 2 20388 20390
0 20392 5 1 1 20391
0 20393 7 1 2 27091 20392
0 20394 5 1 1 20393
0 20395 7 1 2 20380 20394
0 20396 5 1 1 20395
0 20397 7 1 2 23957 20396
0 20398 5 1 1 20397
0 20399 7 1 2 27736 33994
0 20400 5 1 1 20399
0 20401 7 1 2 28048 34456
0 20402 5 1 1 20401
0 20403 7 1 2 34743 37730
0 20404 5 1 1 20403
0 20405 7 1 2 20402 20404
0 20406 5 1 1 20405
0 20407 7 1 2 24044 27158
0 20408 7 1 2 20406 20407
0 20409 5 1 1 20408
0 20410 7 1 2 20400 20409
0 20411 7 1 2 20398 20410
0 20412 5 1 1 20411
0 20413 7 1 2 38217 20412
0 20414 5 1 1 20413
0 20415 7 1 2 20376 20414
0 20416 5 1 1 20415
0 20417 7 1 2 24384 20416
0 20418 5 1 1 20417
0 20419 7 3 2 29121 38216
0 20420 7 1 2 34311 38219
0 20421 7 1 2 38212 20420
0 20422 5 1 1 20421
0 20423 7 1 2 20418 20422
0 20424 5 1 1 20423
0 20425 7 1 2 20263 20424
0 20426 5 1 1 20425
0 20427 7 1 2 35420 31340
0 20428 7 1 2 29934 20427
0 20429 7 1 2 38003 20428
0 20430 7 1 2 37798 36969
0 20431 7 1 2 20429 20430
0 20432 5 1 1 20431
0 20433 7 1 2 35508 38001
0 20434 5 1 1 20433
0 20435 7 1 2 32640 34312
0 20436 7 1 2 35893 20435
0 20437 7 1 2 30515 20436
0 20438 5 1 1 20437
0 20439 7 1 2 20434 20438
0 20440 5 1 1 20439
0 20441 7 1 2 34092 20440
0 20442 5 1 1 20441
0 20443 7 3 2 24306 36334
0 20444 7 1 2 28834 27663
0 20445 7 1 2 36462 20444
0 20446 7 1 2 38222 20445
0 20447 5 1 1 20446
0 20448 7 1 2 20442 20447
0 20449 5 1 1 20448
0 20450 7 1 2 26200 20449
0 20451 5 1 1 20450
0 20452 7 1 2 36651 36900
0 20453 7 1 2 37553 20452
0 20454 7 1 2 38223 20453
0 20455 5 1 1 20454
0 20456 7 1 2 20451 20455
0 20457 5 1 1 20456
0 20458 7 1 2 25391 20457
0 20459 5 1 1 20458
0 20460 7 1 2 22769 35509
0 20461 5 1 1 20460
0 20462 7 1 2 27664 36069
0 20463 5 1 1 20462
0 20464 7 1 2 20461 20463
0 20465 5 1 1 20464
0 20466 7 1 2 23435 36692
0 20467 7 1 2 37826 20466
0 20468 7 1 2 20465 20467
0 20469 5 1 1 20468
0 20470 7 1 2 26017 20469
0 20471 7 1 2 20459 20470
0 20472 5 1 1 20471
0 20473 7 1 2 25005 35258
0 20474 7 2 2 38224 20473
0 20475 7 1 2 27773 29339
0 20476 5 1 1 20475
0 20477 7 1 2 29318 31356
0 20478 5 1 1 20477
0 20479 7 1 2 20476 20478
0 20480 5 1 1 20479
0 20481 7 1 2 25587 20480
0 20482 7 1 2 38225 20481
0 20483 5 1 1 20482
0 20484 7 1 2 24045 20483
0 20485 5 1 1 20484
0 20486 7 1 2 25928 20485
0 20487 7 1 2 20472 20486
0 20488 5 1 1 20487
0 20489 7 1 2 22869 33063
0 20490 5 1 1 20489
0 20491 7 1 2 23436 35502
0 20492 5 1 1 20491
0 20493 7 1 2 20490 20492
0 20494 5 1 1 20493
0 20495 7 1 2 22770 20494
0 20496 5 1 1 20495
0 20497 7 1 2 32648 38114
0 20498 5 1 1 20497
0 20499 7 1 2 20496 20498
0 20500 5 1 1 20499
0 20501 7 1 2 24385 33837
0 20502 7 1 2 36693 20501
0 20503 7 1 2 20500 20502
0 20504 5 1 1 20503
0 20505 7 1 2 29286 35068
0 20506 7 3 2 25449 33473
0 20507 7 1 2 36389 31894
0 20508 7 1 2 38227 20507
0 20509 7 1 2 20505 20508
0 20510 5 1 1 20509
0 20511 7 1 2 20504 20510
0 20512 5 1 1 20511
0 20513 7 1 2 34457 20512
0 20514 5 1 1 20513
0 20515 7 1 2 30195 35061
0 20516 5 1 1 20515
0 20517 7 2 2 30278 34956
0 20518 5 1 1 38230
0 20519 7 1 2 20516 20518
0 20520 5 2 1 20519
0 20521 7 1 2 22771 38232
0 20522 5 1 1 20521
0 20523 7 1 2 33165 38115
0 20524 5 1 1 20523
0 20525 7 1 2 20522 20524
0 20526 5 1 1 20525
0 20527 7 1 2 33096 34339
0 20528 7 1 2 20526 20527
0 20529 5 1 1 20528
0 20530 7 1 2 28567 34523
0 20531 7 1 2 34764 20530
0 20532 7 1 2 31550 20531
0 20533 5 1 1 20532
0 20534 7 1 2 20529 20533
0 20535 5 1 1 20534
0 20536 7 1 2 35553 26579
0 20537 7 1 2 35259 20536
0 20538 7 1 2 20535 20537
0 20539 5 1 1 20538
0 20540 7 1 2 20514 20539
0 20541 7 1 2 20488 20540
0 20542 5 1 1 20541
0 20543 7 1 2 24136 20542
0 20544 5 1 1 20543
0 20545 7 1 2 7877 28411
0 20546 5 1 1 20545
0 20547 7 1 2 29444 20546
0 20548 7 1 2 37992 20547
0 20549 5 1 1 20548
0 20550 7 2 2 24621 33364
0 20551 7 1 2 30196 36283
0 20552 7 1 2 38234 20551
0 20553 5 1 1 20552
0 20554 7 1 2 20549 20553
0 20555 5 1 1 20554
0 20556 7 1 2 35690 38226
0 20557 7 1 2 20555 20556
0 20558 5 1 1 20557
0 20559 7 1 2 20544 20558
0 20560 5 1 1 20559
0 20561 7 1 2 25326 20560
0 20562 5 1 1 20561
0 20563 7 1 2 34142 35510
0 20564 5 1 1 20563
0 20565 7 1 2 9142 20564
0 20566 5 1 1 20565
0 20567 7 1 2 34082 27442
0 20568 7 1 2 35924 20567
0 20569 7 1 2 37718 20568
0 20570 7 1 2 20566 20569
0 20571 5 1 1 20570
0 20572 7 1 2 20562 20571
0 20573 5 1 1 20572
0 20574 7 1 2 24337 37947
0 20575 7 1 2 20573 20574
0 20576 5 1 1 20575
0 20577 7 1 2 20432 20576
0 20578 5 1 1 20577
0 20579 7 1 2 26709 20578
0 20580 5 1 1 20579
0 20581 7 1 2 38098 36992
0 20582 5 1 1 20581
0 20583 7 1 2 29770 34587
0 20584 7 1 2 26721 20583
0 20585 5 1 1 20584
0 20586 7 1 2 20582 20585
0 20587 5 1 1 20586
0 20588 7 1 2 22659 20587
0 20589 5 1 1 20588
0 20590 7 1 2 32025 28927
0 20591 7 1 2 36990 20590
0 20592 5 1 1 20591
0 20593 7 1 2 26548 36908
0 20594 7 1 2 36003 20593
0 20595 5 1 1 20594
0 20596 7 1 2 20592 20595
0 20597 5 1 1 20596
0 20598 7 1 2 34704 20597
0 20599 5 1 1 20598
0 20600 7 1 2 20589 20599
0 20601 5 1 1 20600
0 20602 7 1 2 23286 20601
0 20603 5 1 1 20602
0 20604 7 2 2 35115 35379
0 20605 7 1 2 32303 37441
0 20606 7 1 2 38236 20605
0 20607 5 1 1 20606
0 20608 7 1 2 20603 20607
0 20609 5 1 1 20608
0 20610 7 1 2 23743 20609
0 20611 5 1 1 20610
0 20612 7 1 2 24137 32026
0 20613 7 1 2 27876 31077
0 20614 7 1 2 20612 20613
0 20615 7 1 2 34665 20614
0 20616 5 1 1 20615
0 20617 7 1 2 20611 20616
0 20618 5 1 1 20617
0 20619 7 1 2 22518 20618
0 20620 5 1 1 20619
0 20621 7 1 2 25646 29498
0 20622 7 1 2 33517 20621
0 20623 7 1 2 38072 20622
0 20624 5 1 1 20623
0 20625 7 1 2 26703 31615
0 20626 7 1 2 38237 20625
0 20627 5 1 1 20626
0 20628 7 1 2 20624 20627
0 20629 5 1 1 20628
0 20630 7 1 2 28351 20629
0 20631 5 1 1 20630
0 20632 7 1 2 24714 20631
0 20633 7 1 2 20620 20632
0 20634 5 1 1 20633
0 20635 7 1 2 29963 38058
0 20636 5 1 1 20635
0 20637 7 1 2 29883 26704
0 20638 7 1 2 29724 20637
0 20639 5 1 1 20638
0 20640 7 1 2 20636 20639
0 20641 5 1 1 20640
0 20642 7 1 2 37330 20641
0 20643 5 1 1 20642
0 20644 7 2 2 29381 37555
0 20645 7 1 2 36177 37158
0 20646 7 1 2 38238 20645
0 20647 5 1 1 20646
0 20648 7 1 2 22772 20647
0 20649 7 1 2 20643 20648
0 20650 5 1 1 20649
0 20651 7 1 2 24800 20650
0 20652 7 1 2 20634 20651
0 20653 5 1 1 20652
0 20654 7 1 2 26201 30916
0 20655 5 1 1 20654
0 20656 7 1 2 30922 20655
0 20657 7 1 2 37331 20656
0 20658 5 1 1 20657
0 20659 7 2 2 37482 38139
0 20660 7 1 2 30493 33258
0 20661 7 1 2 38240 20660
0 20662 5 1 1 20661
0 20663 7 1 2 20658 20662
0 20664 5 1 1 20663
0 20665 7 1 2 37234 20664
0 20666 5 1 1 20665
0 20667 7 1 2 24925 20666
0 20668 7 1 2 20653 20667
0 20669 5 1 1 20668
0 20670 7 1 2 32561 37342
0 20671 5 1 1 20670
0 20672 7 1 2 28215 31299
0 20673 7 1 2 37951 20672
0 20674 5 1 1 20673
0 20675 7 1 2 20671 20674
0 20676 5 1 1 20675
0 20677 7 1 2 36880 20676
0 20678 5 1 1 20677
0 20679 7 1 2 36840 14302
0 20680 5 2 1 20679
0 20681 7 1 2 25929 28577
0 20682 7 1 2 38241 20681
0 20683 7 1 2 38242 20682
0 20684 5 1 1 20683
0 20685 7 1 2 22981 20684
0 20686 7 1 2 20678 20685
0 20687 5 1 1 20686
0 20688 7 1 2 20669 20687
0 20689 5 1 1 20688
0 20690 7 1 2 24307 20689
0 20691 5 1 1 20690
0 20692 7 2 2 33850 26631
0 20693 7 1 2 28863 31624
0 20694 5 1 1 20693
0 20695 7 1 2 35570 34152
0 20696 5 1 1 20695
0 20697 7 1 2 20694 20696
0 20698 5 1 1 20697
0 20699 7 1 2 22519 20698
0 20700 5 1 1 20699
0 20701 7 1 2 36630 37338
0 20702 5 1 1 20701
0 20703 7 1 2 20700 20702
0 20704 5 1 1 20703
0 20705 7 1 2 32562 20704
0 20706 5 1 1 20705
0 20707 7 1 2 26018 33365
0 20708 7 1 2 31515 20707
0 20709 7 1 2 37824 20708
0 20710 5 1 1 20709
0 20711 7 1 2 20706 20710
0 20712 5 1 1 20711
0 20713 7 1 2 37124 20712
0 20714 5 1 1 20713
0 20715 7 1 2 27346 30553
0 20716 7 1 2 37894 20715
0 20717 7 1 2 36228 20716
0 20718 5 1 1 20717
0 20719 7 1 2 20714 20718
0 20720 5 1 1 20719
0 20721 7 1 2 38244 20720
0 20722 5 1 1 20721
0 20723 7 1 2 35812 26632
0 20724 7 1 2 33106 20723
0 20725 5 1 1 20724
0 20726 7 1 2 28216 37349
0 20727 7 1 2 36838 20726
0 20728 5 1 1 20727
0 20729 7 1 2 20725 20728
0 20730 5 1 1 20729
0 20731 7 1 2 23744 20730
0 20732 5 1 1 20731
0 20733 7 1 2 32534 37557
0 20734 5 1 1 20733
0 20735 7 1 2 36890 20734
0 20736 5 1 1 20735
0 20737 7 1 2 30178 37210
0 20738 7 1 2 20736 20737
0 20739 5 1 1 20738
0 20740 7 1 2 20732 20739
0 20741 5 1 1 20740
0 20742 7 1 2 37125 20741
0 20743 5 1 1 20742
0 20744 7 1 2 26019 35062
0 20745 7 1 2 30214 37244
0 20746 7 1 2 20744 20745
0 20747 7 1 2 30058 31898
0 20748 7 1 2 20746 20747
0 20749 5 1 1 20748
0 20750 7 1 2 20743 20749
0 20751 5 1 1 20750
0 20752 7 1 2 31948 20751
0 20753 5 1 1 20752
0 20754 7 1 2 26279 20753
0 20755 7 1 2 20722 20754
0 20756 5 1 1 20755
0 20757 7 1 2 24386 20756
0 20758 7 1 2 20691 20757
0 20759 5 1 1 20758
0 20760 7 1 2 34316 20759
0 20761 5 1 1 20760
0 20762 7 1 2 27759 36799
0 20763 5 1 1 20762
0 20764 7 1 2 25006 32233
0 20765 7 1 2 38228 20764
0 20766 5 1 1 20765
0 20767 7 1 2 20763 20766
0 20768 5 3 1 20767
0 20769 7 1 2 31949 37350
0 20770 5 1 1 20769
0 20771 7 1 2 25831 38245
0 20772 5 1 1 20771
0 20773 7 1 2 20770 20772
0 20774 5 2 1 20773
0 20775 7 1 2 28864 38249
0 20776 5 1 1 20775
0 20777 7 1 2 30179 34540
0 20778 7 1 2 26633 20777
0 20779 5 1 1 20778
0 20780 7 1 2 20776 20779
0 20781 5 1 1 20780
0 20782 7 1 2 26280 20781
0 20783 5 1 1 20782
0 20784 7 1 2 30592 37442
0 20785 7 2 2 35603 20784
0 20786 5 1 1 38251
0 20787 7 1 2 32593 38252
0 20788 5 1 1 20787
0 20789 7 1 2 20783 20788
0 20790 5 1 1 20789
0 20791 7 1 2 32563 20790
0 20792 5 1 1 20791
0 20793 7 2 2 26107 36788
0 20794 7 1 2 31357 36178
0 20795 7 1 2 38253 20794
0 20796 5 1 1 20795
0 20797 7 1 2 20792 20796
0 20798 5 1 1 20797
0 20799 7 1 2 37126 20798
0 20800 5 1 1 20799
0 20801 7 1 2 24715 38157
0 20802 5 1 1 20801
0 20803 7 1 2 22773 27244
0 20804 7 1 2 38163 20803
0 20805 5 1 1 20804
0 20806 7 1 2 20802 20805
0 20807 5 1 1 20806
0 20808 7 1 2 31239 20807
0 20809 5 1 1 20808
0 20810 7 1 2 24716 37563
0 20811 5 1 1 20810
0 20812 7 1 2 20809 20811
0 20813 5 1 1 20812
0 20814 7 1 2 22660 20813
0 20815 5 1 1 20814
0 20816 7 1 2 32594 38161
0 20817 5 1 1 20816
0 20818 7 1 2 26853 35532
0 20819 5 1 1 20818
0 20820 7 1 2 20817 20819
0 20821 5 1 1 20820
0 20822 7 1 2 23958 20821
0 20823 5 1 1 20822
0 20824 7 1 2 31177 27709
0 20825 5 1 1 20824
0 20826 7 1 2 20823 20825
0 20827 5 1 1 20826
0 20828 7 1 2 34569 37403
0 20829 7 1 2 20827 20828
0 20830 5 1 1 20829
0 20831 7 1 2 20815 20830
0 20832 7 1 2 20800 20831
0 20833 5 1 1 20832
0 20834 7 1 2 24515 20833
0 20835 5 1 1 20834
0 20836 7 1 2 27933 20835
0 20837 5 1 1 20836
0 20838 7 1 2 29527 38153
0 20839 5 1 1 20838
0 20840 7 1 2 35088 37049
0 20841 5 1 1 20840
0 20842 7 1 2 19727 19950
0 20843 5 1 1 20842
0 20844 7 1 2 33151 20843
0 20845 5 1 1 20844
0 20846 7 1 2 20841 20845
0 20847 5 1 1 20846
0 20848 7 1 2 32595 20847
0 20849 5 1 1 20848
0 20850 7 1 2 20839 20849
0 20851 5 1 1 20850
0 20852 7 1 2 23959 20851
0 20853 5 1 1 20852
0 20854 7 1 2 36284 37619
0 20855 7 1 2 36995 20854
0 20856 5 1 1 20855
0 20857 7 1 2 20853 20856
0 20858 5 1 1 20857
0 20859 7 1 2 24622 20858
0 20860 5 1 1 20859
0 20861 7 1 2 31358 30266
0 20862 7 1 2 37655 20861
0 20863 5 1 1 20862
0 20864 7 1 2 20860 20863
0 20865 5 1 1 20864
0 20866 7 1 2 23854 20865
0 20867 5 1 1 20866
0 20868 7 1 2 28962 20867
0 20869 5 1 1 20868
0 20870 7 1 2 23745 20869
0 20871 7 1 2 20837 20870
0 20872 5 1 1 20871
0 20873 7 1 2 33410 20872
0 20874 5 1 1 20873
0 20875 7 1 2 38246 20874
0 20876 7 1 2 20761 20875
0 20877 5 1 1 20876
0 20878 7 1 2 32372 29501
0 20879 5 1 1 20878
0 20880 7 1 2 28049 31964
0 20881 5 1 1 20880
0 20882 7 1 2 29467 32373
0 20883 5 1 1 20882
0 20884 7 1 2 20881 20883
0 20885 5 1 1 20884
0 20886 7 1 2 22520 20885
0 20887 5 1 1 20886
0 20888 7 1 2 20879 20887
0 20889 5 1 1 20888
0 20890 7 1 2 25588 20889
0 20891 5 1 1 20890
0 20892 7 1 2 27814 38188
0 20893 7 1 2 27139 20892
0 20894 7 1 2 29265 20893
0 20895 5 1 1 20894
0 20896 7 1 2 20891 20895
0 20897 5 1 1 20896
0 20898 7 1 2 24046 20897
0 20899 5 1 1 20898
0 20900 7 2 2 28188 36822
0 20901 7 1 2 31887 29913
0 20902 7 1 2 38255 20901
0 20903 5 1 1 20902
0 20904 7 1 2 20899 20903
0 20905 5 1 1 20904
0 20906 7 1 2 27245 20905
0 20907 5 1 1 20906
0 20908 7 2 2 27246 31198
0 20909 7 1 2 36238 31556
0 20910 5 1 1 20909
0 20911 7 1 2 24516 28081
0 20912 5 1 1 20911
0 20913 7 1 2 20910 20912
0 20914 5 1 1 20913
0 20915 7 1 2 38257 20914
0 20916 5 1 1 20915
0 20917 7 1 2 27358 34705
0 20918 5 1 1 20917
0 20919 7 1 2 31500 20918
0 20920 7 1 2 27824 20919
0 20921 5 1 1 20920
0 20922 7 1 2 28952 20921
0 20923 5 1 1 20922
0 20924 7 1 2 20916 20923
0 20925 5 1 1 20924
0 20926 7 4 2 29499 36823
0 20927 7 1 2 20925 38259
0 20928 5 1 1 20927
0 20929 7 1 2 29366 35315
0 20930 7 1 2 33115 20929
0 20931 7 1 2 28462 29729
0 20932 7 1 2 20930 20931
0 20933 5 1 1 20932
0 20934 7 1 2 20928 20933
0 20935 5 1 1 20934
0 20936 7 1 2 27092 20935
0 20937 5 1 1 20936
0 20938 7 2 2 27899 35952
0 20939 7 1 2 29367 34866
0 20940 7 1 2 38263 20939
0 20941 5 2 1 20940
0 20942 7 2 2 31721 36824
0 20943 7 1 2 35621 37081
0 20944 7 1 2 38267 20943
0 20945 5 1 1 20944
0 20946 7 1 2 38265 20945
0 20947 5 1 1 20946
0 20948 7 1 2 27737 20947
0 20949 5 1 1 20948
0 20950 7 1 2 31129 33706
0 20951 7 1 2 36464 20950
0 20952 7 1 2 38256 20951
0 20953 5 1 1 20952
0 20954 7 1 2 20949 20953
0 20955 7 1 2 20937 20954
0 20956 7 1 2 20907 20955
0 20957 5 1 1 20956
0 20958 7 1 2 35857 20957
0 20959 5 1 1 20958
0 20960 7 2 2 27247 28682
0 20961 7 1 2 31179 38269
0 20962 5 1 1 20961
0 20963 7 1 2 34115 37816
0 20964 5 1 1 20963
0 20965 7 1 2 35789 38054
0 20966 5 1 1 20965
0 20967 7 1 2 35884 20966
0 20968 7 1 2 20964 20967
0 20969 5 1 1 20968
0 20970 7 1 2 25243 20969
0 20971 5 1 1 20970
0 20972 7 1 2 20962 20971
0 20973 5 1 1 20972
0 20974 7 2 2 24517 20973
0 20975 5 1 1 38271
0 20976 7 1 2 31242 38270
0 20977 5 1 1 20976
0 20978 7 1 2 20975 20977
0 20979 5 1 1 20978
0 20980 7 1 2 38260 20979
0 20981 5 1 1 20980
0 20982 7 1 2 35554 37948
0 20983 7 1 2 32036 20982
0 20984 7 1 2 38264 20983
0 20985 5 1 1 20984
0 20986 7 1 2 20981 20985
0 20987 5 1 1 20986
0 20988 7 1 2 29741 20987
0 20989 5 1 1 20988
0 20990 7 1 2 37838 38261
0 20991 5 1 1 20990
0 20992 7 1 2 38266 20991
0 20993 5 1 1 20992
0 20994 7 1 2 35869 20993
0 20995 5 1 1 20994
0 20996 7 2 2 28953 38262
0 20997 7 1 2 28174 38273
0 20998 7 1 2 35867 20997
0 20999 5 1 1 20998
0 21000 7 1 2 20995 20999
0 21001 5 1 1 21000
0 21002 7 1 2 32124 21001
0 21003 5 1 1 21002
0 21004 7 1 2 36825 37082
0 21005 7 1 2 37937 21004
0 21006 7 1 2 37742 21005
0 21007 5 1 1 21006
0 21008 7 2 2 34867 31740
0 21009 7 1 2 23287 32413
0 21010 7 1 2 38275 21009
0 21011 5 1 1 21010
0 21012 7 1 2 25392 33347
0 21013 7 1 2 35622 21012
0 21014 7 1 2 38268 21013
0 21015 5 1 1 21014
0 21016 7 1 2 21011 21015
0 21017 5 1 1 21016
0 21018 7 1 2 27327 21017
0 21019 5 1 1 21018
0 21020 7 1 2 27263 38274
0 21021 5 1 1 21020
0 21022 7 1 2 35458 29368
0 21023 7 1 2 37148 21022
0 21024 5 1 1 21023
0 21025 7 1 2 21021 21024
0 21026 5 1 1 21025
0 21027 7 1 2 34143 21026
0 21028 5 1 1 21027
0 21029 7 1 2 21019 21028
0 21030 7 1 2 21007 21029
0 21031 5 1 1 21030
0 21032 7 1 2 35527 21031
0 21033 5 1 1 21032
0 21034 7 1 2 21003 21033
0 21035 7 1 2 20989 21034
0 21036 5 1 1 21035
0 21037 7 1 2 29019 21036
0 21038 5 1 1 21037
0 21039 7 1 2 33533 30018
0 21040 7 1 2 36826 37818
0 21041 7 1 2 21039 21040
0 21042 7 1 2 35348 21041
0 21043 5 1 1 21042
0 21044 7 1 2 21038 21043
0 21045 7 1 2 20959 21044
0 21046 5 1 1 21045
0 21047 7 1 2 33406 21046
0 21048 5 1 1 21047
0 21049 7 1 2 34035 37607
0 21050 5 1 1 21049
0 21051 7 1 2 30996 33896
0 21052 5 1 1 21051
0 21053 7 1 2 21050 21052
0 21054 5 1 1 21053
0 21055 7 1 2 34275 21054
0 21056 5 1 1 21055
0 21057 7 1 2 26108 38213
0 21058 5 1 1 21057
0 21059 7 1 2 21056 21058
0 21060 5 1 1 21059
0 21061 7 1 2 30370 21060
0 21062 5 1 1 21061
0 21063 7 1 2 34922 37646
0 21064 5 1 1 21063
0 21065 7 1 2 24518 35343
0 21066 5 1 1 21065
0 21067 7 1 2 24138 34208
0 21068 7 1 2 31557 21067
0 21069 5 1 1 21068
0 21070 7 1 2 21066 21069
0 21071 5 1 1 21070
0 21072 7 1 2 37993 21071
0 21073 5 1 1 21072
0 21074 7 1 2 35321 38208
0 21075 5 1 1 21074
0 21076 7 1 2 21073 21075
0 21077 7 1 2 21064 21076
0 21078 5 1 1 21077
0 21079 7 1 2 36577 21078
0 21080 5 1 1 21079
0 21081 7 1 2 36679 37647
0 21082 5 1 1 21081
0 21083 7 1 2 36689 38209
0 21084 5 1 1 21083
0 21085 7 1 2 37994 37793
0 21086 5 1 1 21085
0 21087 7 1 2 21084 21086
0 21088 7 1 2 21082 21087
0 21089 5 1 1 21088
0 21090 7 1 2 34942 21089
0 21091 5 1 1 21090
0 21092 7 1 2 21080 21091
0 21093 5 1 1 21092
0 21094 7 1 2 26202 21093
0 21095 5 1 1 21094
0 21096 7 1 2 21062 21095
0 21097 5 1 1 21096
0 21098 7 1 2 33411 38276
0 21099 7 1 2 21097 21098
0 21100 5 1 1 21099
0 21101 7 1 2 21048 21100
0 21102 5 1 1 21101
0 21103 7 1 2 32067 28901
0 21104 7 1 2 21102 21103
0 21105 5 1 1 21104
0 21106 7 1 2 20877 21105
0 21107 7 1 2 20580 21106
0 21108 7 1 2 20426 21107
0 21109 7 1 2 20261 21108
0 21110 7 1 2 19761 21109
0 21111 7 1 2 35241 30544
0 21112 5 1 1 21111
0 21113 7 1 2 29091 34083
0 21114 5 1 1 21113
0 21115 7 1 2 26477 33577
0 21116 5 1 1 21115
0 21117 7 4 2 21114 21116
0 21118 7 1 2 33901 38277
0 21119 5 1 1 21118
0 21120 7 1 2 32492 37032
0 21121 5 1 1 21120
0 21122 7 1 2 21119 21121
0 21123 5 1 1 21122
0 21124 7 1 2 25244 35784
0 21125 5 1 1 21124
0 21126 7 1 2 31199 33219
0 21127 5 1 1 21126
0 21128 7 1 2 21125 21127
0 21129 5 1 1 21128
0 21130 7 1 2 21123 21129
0 21131 5 1 1 21130
0 21132 7 1 2 29231 34036
0 21133 5 1 1 21132
0 21134 7 1 2 20313 21133
0 21135 5 1 1 21134
0 21136 7 1 2 33937 38278
0 21137 5 1 1 21136
0 21138 7 1 2 35779 37033
0 21139 5 1 1 21138
0 21140 7 1 2 21137 21139
0 21141 5 1 1 21140
0 21142 7 1 2 21135 21141
0 21143 5 1 1 21142
0 21144 7 1 2 21131 21143
0 21145 5 1 1 21144
0 21146 7 1 2 38176 21145
0 21147 5 1 1 21146
0 21148 7 1 2 34037 33938
0 21149 5 1 1 21148
0 21150 7 1 2 25393 33366
0 21151 7 1 2 34974 21150
0 21152 5 1 1 21151
0 21153 7 1 2 21149 21152
0 21154 5 1 1 21153
0 21155 7 1 2 38279 21154
0 21156 5 1 1 21155
0 21157 7 1 2 25394 36113
0 21158 5 1 1 21157
0 21159 7 1 2 27632 29904
0 21160 5 1 1 21159
0 21161 7 1 2 21158 21160
0 21162 5 1 1 21161
0 21163 7 1 2 24717 21162
0 21164 5 1 1 21163
0 21165 7 1 2 24139 27115
0 21166 5 1 1 21165
0 21167 7 1 2 21164 21166
0 21168 5 1 1 21167
0 21169 7 1 2 37034 21168
0 21170 5 1 1 21169
0 21171 7 1 2 21156 21170
0 21172 5 1 1 21171
0 21173 7 1 2 21172 37084
0 21174 5 1 1 21173
0 21175 7 2 2 22870 29837
0 21176 7 1 2 38281 36734
0 21177 5 1 1 21176
0 21178 7 1 2 22982 32171
0 21179 7 1 2 32465 21178
0 21180 5 1 1 21179
0 21181 7 1 2 34987 36578
0 21182 5 1 1 21181
0 21183 7 1 2 26464 35598
0 21184 5 1 1 21183
0 21185 7 1 2 21182 21184
0 21186 7 1 2 21180 21185
0 21187 5 1 1 21186
0 21188 7 1 2 23437 21187
0 21189 5 1 1 21188
0 21190 7 1 2 21177 21189
0 21191 5 1 1 21190
0 21192 7 1 2 22774 21191
0 21193 5 1 1 21192
0 21194 7 1 2 36927 21193
0 21195 5 1 1 21194
0 21196 7 2 2 30605 37506
0 21197 7 1 2 21195 38283
0 21198 5 1 1 21197
0 21199 7 1 2 24623 21198
0 21200 7 1 2 21174 21199
0 21201 5 1 1 21200
0 21202 7 1 2 32256 32936
0 21203 5 1 1 21202
0 21204 7 1 2 32125 36972
0 21205 5 1 1 21204
0 21206 7 1 2 21203 21205
0 21207 5 1 1 21206
0 21208 7 1 2 32741 21207
0 21209 5 1 1 21208
0 21210 7 1 2 32658 38243
0 21211 5 1 1 21210
0 21212 7 1 2 32535 30373
0 21213 5 1 1 21212
0 21214 7 1 2 33152 28751
0 21215 5 1 1 21214
0 21216 7 1 2 21213 21215
0 21217 5 1 1 21216
0 21218 7 1 2 33064 21217
0 21219 5 1 1 21218
0 21220 7 1 2 21211 21219
0 21221 7 1 2 21209 21220
0 21222 5 1 1 21221
0 21223 7 1 2 38180 21222
0 21224 5 1 1 21223
0 21225 7 1 2 22661 21224
0 21226 5 1 1 21225
0 21227 7 1 2 25930 21226
0 21228 7 1 2 21201 21227
0 21229 5 1 1 21228
0 21230 7 1 2 35926 36579
0 21231 5 1 1 21230
0 21232 7 2 2 30954 26854
0 21233 7 1 2 25516 38285
0 21234 5 1 1 21233
0 21235 7 1 2 34957 37194
0 21236 5 1 1 21235
0 21237 7 1 2 21234 21236
0 21238 5 1 1 21237
0 21239 7 1 2 22775 21238
0 21240 5 1 1 21239
0 21241 7 1 2 27039 36647
0 21242 5 1 1 21241
0 21243 7 1 2 21240 21242
0 21244 5 1 1 21243
0 21245 7 1 2 34943 21244
0 21246 5 1 1 21245
0 21247 7 1 2 21231 21246
0 21248 5 1 1 21247
0 21249 7 1 2 31636 38284
0 21250 7 1 2 21248 21249
0 21251 5 1 1 21250
0 21252 7 1 2 21229 21251
0 21253 5 1 1 21252
0 21254 7 1 2 22521 21253
0 21255 5 1 1 21254
0 21256 7 1 2 21147 21255
0 21257 5 1 1 21256
0 21258 7 1 2 23855 21257
0 21259 5 1 1 21258
0 21260 7 1 2 33939 38198
0 21261 5 1 1 21260
0 21262 7 1 2 33902 38201
0 21263 5 1 1 21262
0 21264 7 1 2 21261 21263
0 21265 5 1 1 21264
0 21266 7 1 2 38280 21265
0 21267 5 1 1 21266
0 21268 7 1 2 32493 38202
0 21269 5 1 1 21268
0 21270 7 1 2 35780 38199
0 21271 5 1 1 21270
0 21272 7 1 2 21269 21271
0 21273 5 1 1 21272
0 21274 7 1 2 37035 21273
0 21275 5 1 1 21274
0 21276 7 1 2 21267 21275
0 21277 5 1 1 21276
0 21278 7 1 2 38194 21277
0 21279 5 1 1 21278
0 21280 7 1 2 21259 21279
0 21281 5 1 1 21280
0 21282 7 1 2 25160 21281
0 21283 5 1 1 21282
0 21284 7 3 2 33578 37949
0 21285 7 1 2 28175 36864
0 21286 5 1 1 21285
0 21287 7 1 2 30388 37201
0 21288 5 1 1 21287
0 21289 7 1 2 21286 21288
0 21290 5 1 1 21289
0 21291 7 1 2 25245 21290
0 21292 5 1 1 21291
0 21293 7 1 2 31207 37638
0 21294 5 1 1 21293
0 21295 7 1 2 21292 21294
0 21296 5 1 1 21295
0 21297 7 1 2 24519 21296
0 21298 5 1 1 21297
0 21299 7 1 2 35260 30033
0 21300 7 1 2 29242 21299
0 21301 5 1 1 21300
0 21302 7 1 2 21298 21301
0 21303 5 1 1 21302
0 21304 7 1 2 25931 38282
0 21305 7 1 2 21303 21304
0 21306 5 1 1 21305
0 21307 7 1 2 10914 16507
0 21308 5 1 1 21307
0 21309 7 1 2 29266 21308
0 21310 5 1 1 21309
0 21311 7 1 2 30880 33138
0 21312 7 1 2 30325 21311
0 21313 5 1 1 21312
0 21314 7 1 2 21310 21313
0 21315 5 1 1 21314
0 21316 7 1 2 27093 21315
0 21317 5 1 1 21316
0 21318 7 1 2 25395 37644
0 21319 5 1 1 21318
0 21320 7 1 2 18013 21319
0 21321 5 2 1 21320
0 21322 7 1 2 37494 38290
0 21323 5 1 1 21322
0 21324 7 1 2 28176 31909
0 21325 7 2 2 37370 21324
0 21326 7 1 2 32937 38292
0 21327 5 1 1 21326
0 21328 7 1 2 21323 21327
0 21329 7 1 2 21317 21328
0 21330 5 1 1 21329
0 21331 7 1 2 32742 21330
0 21332 5 1 1 21331
0 21333 7 1 2 33065 37648
0 21334 5 1 1 21333
0 21335 7 1 2 32659 38210
0 21336 5 1 1 21335
0 21337 7 1 2 37995 37997
0 21338 5 1 1 21337
0 21339 7 1 2 21336 21338
0 21340 7 1 2 21334 21339
0 21341 5 1 1 21340
0 21342 7 1 2 33153 21341
0 21343 5 1 1 21342
0 21344 7 1 2 21332 21343
0 21345 7 1 2 21306 21344
0 21346 5 1 1 21345
0 21347 7 2 2 38287 21346
0 21348 7 1 2 36373 38294
0 21349 5 1 1 21348
0 21350 7 1 2 21283 21349
0 21351 5 1 1 21350
0 21352 7 1 2 24387 21351
0 21353 5 1 1 21352
0 21354 7 1 2 23156 34313
0 21355 7 1 2 38295 21354
0 21356 5 1 1 21355
0 21357 7 1 2 21353 21356
0 21358 5 1 1 21357
0 21359 7 1 2 21112 21358
0 21360 5 1 1 21359
0 21361 7 2 2 24926 37184
0 21362 5 1 1 38296
0 21363 7 1 2 32029 36913
0 21364 5 1 1 21363
0 21365 7 1 2 21362 21364
0 21366 5 4 1 21365
0 21367 7 1 2 13398 31618
0 21368 5 1 1 21367
0 21369 7 1 2 10228 21368
0 21370 7 1 2 38298 21369
0 21371 5 1 1 21370
0 21372 7 1 2 30092 31107
0 21373 7 1 2 36914 21372
0 21374 7 1 2 38014 21373
0 21375 5 1 1 21374
0 21376 7 1 2 21371 21375
0 21377 5 1 1 21376
0 21378 7 1 2 33341 21377
0 21379 5 1 1 21378
0 21380 7 1 2 36789 37847
0 21381 5 1 1 21380
0 21382 7 1 2 29701 26611
0 21383 7 1 2 38006 21382
0 21384 5 1 1 21383
0 21385 7 1 2 21381 21384
0 21386 5 1 1 21385
0 21387 7 1 2 36632 21386
0 21388 5 1 1 21387
0 21389 7 1 2 21379 21388
0 21390 5 1 1 21389
0 21391 7 1 2 32461 21390
0 21392 5 1 1 21391
0 21393 7 2 2 23485 31240
0 21394 5 1 1 38302
0 21395 7 1 2 19870 21394
0 21396 5 1 1 21395
0 21397 7 1 2 26109 5077
0 21398 7 1 2 21396 21397
0 21399 5 1 1 21398
0 21400 7 1 2 23486 36672
0 21401 5 1 1 21400
0 21402 7 1 2 21399 21401
0 21403 5 1 1 21402
0 21404 7 1 2 36179 21403
0 21405 5 1 1 21404
0 21406 7 1 2 36540 31535
0 21407 7 1 2 36996 21406
0 21408 5 1 1 21407
0 21409 7 1 2 21405 21408
0 21410 5 1 1 21409
0 21411 7 1 2 35608 37039
0 21412 7 1 2 21410 21411
0 21413 5 1 1 21412
0 21414 7 1 2 22871 38299
0 21415 5 1 1 21414
0 21416 7 1 2 35031 38133
0 21417 5 1 1 21416
0 21418 7 1 2 21415 21417
0 21419 5 1 1 21418
0 21420 7 1 2 36261 21419
0 21421 5 1 1 21420
0 21422 7 1 2 35837 35234
0 21423 5 1 1 21422
0 21424 7 1 2 28409 28394
0 21425 5 2 1 21424
0 21426 7 1 2 24801 37167
0 21427 5 1 1 21426
0 21428 7 1 2 38304 21427
0 21429 5 3 1 21428
0 21430 7 1 2 24338 38305
0 21431 5 2 1 21430
0 21432 7 2 2 38306 38309
0 21433 7 1 2 29702 38311
0 21434 5 1 1 21433
0 21435 7 1 2 21423 21434
0 21436 5 1 1 21435
0 21437 7 1 2 25104 21436
0 21438 5 1 1 21437
0 21439 7 1 2 36239 38151
0 21440 5 1 1 21439
0 21441 7 1 2 21438 21440
0 21442 5 1 1 21441
0 21443 7 1 2 22983 21442
0 21444 5 1 1 21443
0 21445 7 1 2 35089 29673
0 21446 7 1 2 37185 21445
0 21447 5 1 1 21446
0 21448 7 1 2 21444 21447
0 21449 5 1 1 21448
0 21450 7 1 2 36078 21449
0 21451 5 1 1 21450
0 21452 7 1 2 21421 21451
0 21453 7 1 2 21413 21452
0 21454 7 1 2 21392 21453
0 21455 5 1 1 21454
0 21456 7 1 2 28177 21455
0 21457 5 1 1 21456
0 21458 7 1 2 35849 38134
0 21459 5 1 1 21458
0 21460 7 1 2 26875 38300
0 21461 5 1 1 21460
0 21462 7 1 2 21459 21461
0 21463 5 1 1 21462
0 21464 7 1 2 36057 21463
0 21465 5 1 1 21464
0 21466 7 1 2 24047 27248
0 21467 7 1 2 31919 21466
0 21468 7 1 2 36915 38130
0 21469 7 1 2 21467 21468
0 21470 5 1 1 21469
0 21471 7 1 2 21465 21470
0 21472 5 1 1 21471
0 21473 7 1 2 32462 21472
0 21474 5 1 1 21473
0 21475 7 1 2 27539 36790
0 21476 5 1 1 21475
0 21477 7 1 2 35704 30920
0 21478 5 1 1 21477
0 21479 7 1 2 21476 21478
0 21480 5 1 1 21479
0 21481 7 1 2 23487 21480
0 21482 5 1 1 21481
0 21483 7 1 2 30603 32441
0 21484 7 1 2 29331 21483
0 21485 5 1 1 21484
0 21486 7 1 2 21482 21485
0 21487 5 1 1 21486
0 21488 7 1 2 33043 37931
0 21489 7 1 2 21487 21488
0 21490 5 1 1 21489
0 21491 7 1 2 21474 21490
0 21492 5 1 1 21491
0 21493 7 1 2 29232 21492
0 21494 5 1 1 21493
0 21495 7 1 2 23746 37351
0 21496 7 1 2 38009 21495
0 21497 5 1 1 21496
0 21498 7 2 2 26324 31722
0 21499 7 1 2 34600 30589
0 21500 7 1 2 38313 21499
0 21501 5 1 1 21500
0 21502 7 1 2 21497 21501
0 21503 5 1 1 21502
0 21504 7 1 2 32997 33118
0 21505 7 1 2 21503 21504
0 21506 5 1 1 21505
0 21507 7 1 2 29432 37237
0 21508 5 1 1 21507
0 21509 7 1 2 32334 29470
0 21510 5 1 1 21509
0 21511 7 1 2 21508 21510
0 21512 5 1 1 21511
0 21513 7 1 2 26876 37545
0 21514 7 1 2 21512 21513
0 21515 5 1 1 21514
0 21516 7 1 2 21506 21515
0 21517 5 1 1 21516
0 21518 7 1 2 22984 21517
0 21519 5 1 1 21518
0 21520 7 1 2 30538 37241
0 21521 5 1 1 21520
0 21522 7 3 2 24216 36857
0 21523 5 1 1 38315
0 21524 7 1 2 32335 38316
0 21525 5 1 1 21524
0 21526 7 1 2 21521 21525
0 21527 5 1 1 21526
0 21528 7 1 2 27423 32321
0 21529 7 1 2 31955 21528
0 21530 7 1 2 21527 21529
0 21531 5 1 1 21530
0 21532 7 1 2 21519 21531
0 21533 5 1 1 21532
0 21534 7 1 2 34944 21533
0 21535 5 1 1 21534
0 21536 7 1 2 30474 37739
0 21537 7 1 2 32407 21536
0 21538 5 1 1 21537
0 21539 7 1 2 33181 31222
0 21540 7 1 2 30611 21539
0 21541 5 1 1 21540
0 21542 7 1 2 21538 21541
0 21543 5 1 1 21542
0 21544 7 1 2 36386 21543
0 21545 5 1 1 21544
0 21546 7 1 2 23488 31516
0 21547 7 1 2 29243 21546
0 21548 7 1 2 27540 21547
0 21549 5 1 1 21548
0 21550 7 1 2 21545 21549
0 21551 5 1 1 21550
0 21552 7 1 2 33119 21551
0 21553 5 1 1 21552
0 21554 7 1 2 28352 30494
0 21555 7 1 2 32322 21554
0 21556 7 1 2 36270 21555
0 21557 7 1 2 33925 21556
0 21558 5 1 1 21557
0 21559 7 1 2 21553 21558
0 21560 5 1 1 21559
0 21561 7 1 2 36791 21560
0 21562 5 1 1 21561
0 21563 7 1 2 27655 37270
0 21564 5 1 1 21563
0 21565 7 1 2 24927 38303
0 21566 5 1 1 21565
0 21567 7 1 2 21564 21566
0 21568 5 1 1 21567
0 21569 7 1 2 27401 33822
0 21570 7 1 2 34537 21569
0 21571 7 1 2 31247 21570
0 21572 7 1 2 21568 21571
0 21573 5 1 1 21572
0 21574 7 1 2 21562 21573
0 21575 7 1 2 21535 21574
0 21576 7 1 2 21494 21575
0 21577 7 1 2 21457 21576
0 21578 5 1 1 21577
0 21579 7 1 2 32126 21578
0 21580 5 1 1 21579
0 21581 7 1 2 26855 38301
0 21582 5 1 1 21581
0 21583 7 1 2 36792 38231
0 21584 5 1 1 21583
0 21585 7 1 2 21582 21584
0 21586 5 2 1 21585
0 21587 7 1 2 37326 38318
0 21588 5 1 1 21587
0 21589 7 2 2 26856 37546
0 21590 5 2 1 38320
0 21591 7 1 2 34157 37168
0 21592 5 1 1 21591
0 21593 7 1 2 38322 21592
0 21594 5 2 1 21593
0 21595 7 1 2 38102 38324
0 21596 5 1 1 21595
0 21597 7 1 2 34541 36753
0 21598 5 1 1 21597
0 21599 7 1 2 28428 38100
0 21600 5 1 1 21599
0 21601 7 1 2 21598 21600
0 21602 5 1 1 21601
0 21603 7 1 2 26203 34158
0 21604 7 1 2 21602 21603
0 21605 5 1 1 21604
0 21606 7 1 2 21596 21605
0 21607 5 1 1 21606
0 21608 7 1 2 29693 21607
0 21609 5 1 1 21608
0 21610 7 1 2 24339 38323
0 21611 5 1 1 21610
0 21612 7 2 2 38325 21611
0 21613 7 1 2 28452 29680
0 21614 7 1 2 33857 21613
0 21615 7 1 2 38326 21614
0 21616 5 1 1 21615
0 21617 7 1 2 21609 21616
0 21618 5 1 1 21617
0 21619 7 1 2 22985 21618
0 21620 5 1 1 21619
0 21621 7 1 2 32223 32348
0 21622 7 1 2 29674 21621
0 21623 7 1 2 38297 21622
0 21624 5 1 1 21623
0 21625 7 1 2 21620 21624
0 21626 7 1 2 21588 21625
0 21627 5 1 1 21626
0 21628 7 1 2 32257 21627
0 21629 5 1 1 21628
0 21630 7 1 2 37293 38319
0 21631 5 1 1 21630
0 21632 7 1 2 31814 37938
0 21633 7 1 2 38327 21632
0 21634 5 1 1 21633
0 21635 7 1 2 21631 21634
0 21636 5 1 1 21635
0 21637 7 1 2 32851 21636
0 21638 5 1 1 21637
0 21639 7 1 2 31021 37085
0 21640 5 1 1 21639
0 21641 7 2 2 32037 29425
0 21642 5 2 1 38328
0 21643 7 1 2 21640 38330
0 21644 5 2 1 21643
0 21645 7 1 2 32336 38332
0 21646 5 1 1 21645
0 21647 7 1 2 6710 38331
0 21648 5 1 1 21647
0 21649 7 1 2 37238 21648
0 21650 5 1 1 21649
0 21651 7 1 2 21646 21650
0 21652 5 1 1 21651
0 21653 7 1 2 38321 21652
0 21654 5 1 1 21653
0 21655 7 1 2 38329 37354
0 21656 5 1 1 21655
0 21657 7 1 2 31714 33390
0 21658 7 1 2 38185 21657
0 21659 7 1 2 38314 21658
0 21660 5 1 1 21659
0 21661 7 1 2 21656 21660
0 21662 5 1 1 21661
0 21663 7 1 2 34159 32998
0 21664 7 1 2 21662 21663
0 21665 5 1 1 21664
0 21666 7 1 2 21654 21665
0 21667 5 1 1 21666
0 21668 7 1 2 22986 21667
0 21669 5 1 1 21668
0 21670 7 1 2 31053 31885
0 21671 7 1 2 36271 21670
0 21672 7 1 2 30268 37624
0 21673 7 1 2 21671 21672
0 21674 5 1 1 21673
0 21675 7 1 2 21669 21674
0 21676 5 1 1 21675
0 21677 7 1 2 31691 21676
0 21678 5 1 1 21677
0 21679 7 1 2 26960 30554
0 21680 7 1 2 37271 38235
0 21681 7 1 2 38186 21680
0 21682 7 1 2 21679 21681
0 21683 5 1 1 21682
0 21684 7 1 2 26500 31637
0 21685 7 1 2 31054 35063
0 21686 7 1 2 21684 21685
0 21687 7 1 2 38333 21686
0 21688 5 1 1 21687
0 21689 7 1 2 21683 21688
0 21690 5 1 1 21689
0 21691 7 1 2 26204 21690
0 21692 5 1 1 21691
0 21693 7 1 2 36546 31559
0 21694 7 1 2 38286 21693
0 21695 7 1 2 38317 21694
0 21696 5 1 1 21695
0 21697 7 1 2 21692 21696
0 21698 5 1 1 21697
0 21699 7 1 2 32337 21698
0 21700 5 1 1 21699
0 21701 7 1 2 33318 37333
0 21702 5 1 1 21701
0 21703 7 1 2 28683 34811
0 21704 7 1 2 37336 21703
0 21705 5 1 1 21704
0 21706 7 2 2 21702 21705
0 21707 5 1 1 38334
0 21708 7 1 2 36793 38233
0 21709 7 1 2 21707 21708
0 21710 5 1 1 21709
0 21711 7 1 2 21700 21710
0 21712 7 1 2 21678 21711
0 21713 7 1 2 21638 21712
0 21714 7 1 2 21629 21713
0 21715 5 1 1 21714
0 21716 7 1 2 34945 21715
0 21717 5 1 1 21716
0 21718 7 2 2 25720 38312
0 21719 7 1 2 38272 38336
0 21720 5 1 1 21719
0 21721 7 1 2 32258 18104
0 21722 5 1 1 21721
0 21723 7 1 2 35225 38258
0 21724 7 1 2 38310 21723
0 21725 5 1 1 21724
0 21726 7 1 2 32852 37334
0 21727 5 1 1 21726
0 21728 7 1 2 28020 27877
0 21729 7 1 2 37265 21728
0 21730 5 1 1 21729
0 21731 7 1 2 22522 21730
0 21732 7 1 2 21727 21731
0 21733 7 1 2 21725 21732
0 21734 7 1 2 21722 21733
0 21735 5 1 1 21734
0 21736 7 1 2 23747 34674
0 21737 7 1 2 35871 21736
0 21738 5 1 1 21737
0 21739 7 1 2 34144 37766
0 21740 5 1 1 21739
0 21741 7 1 2 24624 28879
0 21742 7 1 2 37266 21741
0 21743 5 1 1 21742
0 21744 7 1 2 21740 21743
0 21745 7 1 2 21738 21744
0 21746 5 1 1 21745
0 21747 7 1 2 23288 21746
0 21748 5 1 1 21747
0 21749 7 1 2 34350 30141
0 21750 7 1 2 37478 21749
0 21751 5 1 1 21750
0 21752 7 1 2 24520 21751
0 21753 7 1 2 21748 21752
0 21754 5 1 1 21753
0 21755 7 1 2 38307 21754
0 21756 7 1 2 21735 21755
0 21757 5 1 1 21756
0 21758 7 1 2 21720 21757
0 21759 5 1 1 21758
0 21760 7 1 2 25105 21759
0 21761 5 1 1 21760
0 21762 7 1 2 26205 31334
0 21763 7 2 2 36754 21762
0 21764 7 1 2 34127 38338
0 21765 5 1 1 21764
0 21766 7 1 2 24308 27271
0 21767 7 1 2 34351 21766
0 21768 7 1 2 38239 21767
0 21769 5 1 1 21768
0 21770 7 1 2 21765 21769
0 21771 5 1 1 21770
0 21772 7 1 2 27328 21771
0 21773 5 1 1 21772
0 21774 7 1 2 35596 38339
0 21775 5 1 1 21774
0 21776 7 1 2 28000 29732
0 21777 7 1 2 32427 21776
0 21778 7 1 2 36916 21777
0 21779 5 1 1 21778
0 21780 7 1 2 21775 21779
0 21781 5 1 1 21780
0 21782 7 1 2 34145 21781
0 21783 5 1 1 21782
0 21784 7 1 2 29943 35133
0 21785 7 1 2 35736 21784
0 21786 7 1 2 37320 21785
0 21787 5 1 1 21786
0 21788 7 1 2 21783 21787
0 21789 7 1 2 21773 21788
0 21790 5 1 1 21789
0 21791 7 1 2 23748 21790
0 21792 5 1 1 21791
0 21793 7 1 2 27651 31651
0 21794 7 1 2 37396 21793
0 21795 7 1 2 37965 21794
0 21796 5 1 1 21795
0 21797 7 1 2 21792 21796
0 21798 7 1 2 21761 21797
0 21799 5 1 1 21798
0 21800 7 1 2 22987 21799
0 21801 5 1 1 21800
0 21802 7 1 2 37327 37186
0 21803 5 1 1 21802
0 21804 7 1 2 26281 38250
0 21805 5 1 1 21804
0 21806 7 1 2 20786 21805
0 21807 5 1 1 21806
0 21808 7 1 2 24217 21807
0 21809 5 1 1 21808
0 21810 7 1 2 30539 38103
0 21811 5 1 1 21810
0 21812 7 1 2 21809 21811
0 21813 5 1 1 21812
0 21814 7 1 2 29694 21813
0 21815 5 1 1 21814
0 21816 7 1 2 21803 21815
0 21817 5 1 1 21816
0 21818 7 1 2 32259 21817
0 21819 5 1 1 21818
0 21820 7 1 2 32853 37294
0 21821 5 1 1 21820
0 21822 7 1 2 21821 38335
0 21823 5 1 1 21822
0 21824 7 1 2 37187 21823
0 21825 5 1 1 21824
0 21826 7 1 2 30545 21523
0 21827 5 1 1 21826
0 21828 7 1 2 33226 32038
0 21829 7 1 2 37889 21828
0 21830 7 1 2 21827 21829
0 21831 5 1 1 21830
0 21832 7 1 2 21825 21831
0 21833 7 1 2 21819 21832
0 21834 5 1 1 21833
0 21835 7 1 2 35090 21834
0 21836 5 1 1 21835
0 21837 7 1 2 21801 21836
0 21838 5 1 1 21837
0 21839 7 1 2 34988 21838
0 21840 5 1 1 21839
0 21841 7 1 2 38019 38308
0 21842 5 1 1 21841
0 21843 7 2 2 25832 29233
0 21844 7 1 2 36755 38340
0 21845 5 1 1 21844
0 21846 7 1 2 36248 38007
0 21847 5 1 1 21846
0 21848 7 1 2 21845 21847
0 21849 5 1 1 21848
0 21850 7 1 2 38147 21849
0 21851 5 1 1 21850
0 21852 7 1 2 21842 21851
0 21853 5 1 1 21852
0 21854 7 1 2 22523 21853
0 21855 5 1 1 21854
0 21856 7 1 2 33823 37547
0 21857 5 1 1 21856
0 21858 7 1 2 24802 38135
0 21859 5 1 1 21858
0 21860 7 1 2 21857 21859
0 21861 5 1 1 21860
0 21862 7 1 2 28371 21861
0 21863 5 1 1 21862
0 21864 7 1 2 21855 21863
0 21865 5 1 1 21864
0 21866 7 1 2 34575 21865
0 21867 5 1 1 21866
0 21868 7 1 2 25106 32127
0 21869 7 1 2 37839 21868
0 21870 7 1 2 38337 21869
0 21871 5 1 1 21870
0 21872 7 1 2 21867 21871
0 21873 5 1 1 21872
0 21874 7 1 2 22988 21873
0 21875 5 1 1 21874
0 21876 7 1 2 36794 38341
0 21877 5 1 1 21876
0 21878 7 1 2 26282 36249
0 21879 7 1 2 37352 21878
0 21880 5 1 1 21879
0 21881 7 1 2 21877 21880
0 21882 5 1 1 21881
0 21883 7 1 2 24218 21882
0 21884 5 1 1 21883
0 21885 7 1 2 30540 38020
0 21886 5 1 1 21885
0 21887 7 1 2 21884 21886
0 21888 5 1 1 21887
0 21889 7 1 2 22524 21888
0 21890 5 1 1 21889
0 21891 7 1 2 28369 38149
0 21892 5 1 1 21891
0 21893 7 1 2 21890 21892
0 21894 5 1 1 21893
0 21895 7 1 2 35091 34576
0 21896 7 1 2 21894 21895
0 21897 5 1 1 21896
0 21898 7 1 2 21875 21897
0 21899 5 1 1 21898
0 21900 7 1 2 33806 21899
0 21901 5 1 1 21900
0 21902 7 1 2 32447 36858
0 21903 5 1 1 21902
0 21904 7 1 2 25450 38254
0 21905 5 1 1 21904
0 21906 7 1 2 21903 21905
0 21907 5 1 1 21906
0 21908 7 1 2 24219 21907
0 21909 5 1 1 21908
0 21910 7 1 2 34946 2343
0 21911 7 1 2 30541 21910
0 21912 5 1 1 21911
0 21913 7 1 2 21909 21912
0 21914 5 1 1 21913
0 21915 7 1 2 24928 21914
0 21916 5 1 1 21915
0 21917 7 1 2 27656 36673
0 21918 5 1 1 21917
0 21919 7 1 2 21916 21918
0 21920 5 1 1 21919
0 21921 7 1 2 26020 21920
0 21922 5 1 1 21921
0 21923 7 1 2 23489 35737
0 21924 7 1 2 35731 21923
0 21925 5 1 1 21924
0 21926 7 1 2 21922 21925
0 21927 5 1 1 21926
0 21928 7 1 2 36240 31577
0 21929 7 1 2 32904 21928
0 21930 7 1 2 21927 21929
0 21931 5 1 1 21930
0 21932 7 1 2 21901 21931
0 21933 7 1 2 21840 21932
0 21934 7 1 2 21717 21933
0 21935 7 1 2 21580 21934
0 21936 5 1 1 21935
0 21937 7 1 2 24388 21936
0 21938 5 1 1 21937
0 21939 7 1 2 34317 21938
0 21940 5 1 1 21939
0 21941 7 1 2 24521 38017
0 21942 5 1 1 21941
0 21943 7 1 2 3116 21942
0 21944 5 3 1 21943
0 21945 7 1 2 30901 38342
0 21946 5 1 1 21945
0 21947 7 1 2 27249 37617
0 21948 5 1 1 21947
0 21949 7 1 2 21946 21948
0 21950 5 1 1 21949
0 21951 7 1 2 34038 21950
0 21952 5 1 1 21951
0 21953 7 1 2 23856 33246
0 21954 5 1 1 21953
0 21955 7 1 2 33891 33726
0 21956 5 1 1 21955
0 21957 7 1 2 21954 21956
0 21958 5 1 1 21957
0 21959 7 1 2 25246 21958
0 21960 5 1 1 21959
0 21961 7 1 2 37843 21960
0 21962 5 1 1 21961
0 21963 7 1 2 24522 21962
0 21964 5 1 1 21963
0 21965 7 1 2 37883 21964
0 21966 5 1 1 21965
0 21967 7 1 2 30997 21966
0 21968 5 1 1 21967
0 21969 7 1 2 21952 21968
0 21970 5 1 1 21969
0 21971 7 1 2 34276 21970
0 21972 5 1 1 21971
0 21973 7 1 2 31700 37652
0 21974 5 1 1 21973
0 21975 7 1 2 38172 38343
0 21976 5 1 1 21975
0 21977 7 1 2 32813 28954
0 21978 5 1 1 21977
0 21979 7 1 2 21976 21978
0 21980 5 1 1 21979
0 21981 7 1 2 28743 21980
0 21982 5 1 1 21981
0 21983 7 1 2 32356 38344
0 21984 5 1 1 21983
0 21985 7 1 2 23857 33044
0 21986 7 1 2 27878 21985
0 21987 7 1 2 27766 21986
0 21988 5 1 1 21987
0 21989 7 1 2 21984 21988
0 21990 5 1 1 21989
0 21991 7 1 2 23960 21990
0 21992 5 1 1 21991
0 21993 7 1 2 33831 28710
0 21994 7 1 2 37800 21993
0 21995 5 1 1 21994
0 21996 7 1 2 21992 21995
0 21997 5 1 1 21996
0 21998 7 1 2 32596 21997
0 21999 5 1 1 21998
0 22000 7 1 2 21982 21999
0 22001 7 1 2 21974 22000
0 22002 5 1 1 22001
0 22003 7 1 2 26110 22002
0 22004 5 1 1 22003
0 22005 7 1 2 21972 22004
0 22006 5 1 1 22005
0 22007 7 1 2 37127 22006
0 22008 5 1 1 22007
0 22009 7 1 2 34581 30263
0 22010 7 1 2 37604 22009
0 22011 5 1 1 22010
0 22012 7 1 2 22008 22011
0 22013 5 1 1 22012
0 22014 7 1 2 28395 22013
0 22015 5 1 1 22014
0 22016 7 1 2 32883 28328
0 22017 5 1 1 22016
0 22018 7 1 2 18420 22017
0 22019 5 1 1 22018
0 22020 7 1 2 32128 22019
0 22021 5 1 1 22020
0 22022 7 1 2 25833 32938
0 22023 7 1 2 35155 22022
0 22024 5 1 1 22023
0 22025 7 1 2 22021 22024
0 22026 5 1 1 22025
0 22027 7 1 2 29345 33307
0 22028 5 1 1 22027
0 22029 7 1 2 9138 22028
0 22030 7 1 2 22026 22029
0 22031 5 1 1 22030
0 22032 7 1 2 28329 37972
0 22033 5 1 1 22032
0 22034 7 1 2 20195 22033
0 22035 5 1 1 22034
0 22036 7 1 2 945 29323
0 22037 5 1 1 22036
0 22038 7 1 2 33308 3168
0 22039 7 1 2 22037 22038
0 22040 7 1 2 22035 22039
0 22041 5 1 1 22040
0 22042 7 1 2 33107 34542
0 22043 5 1 1 22042
0 22044 7 1 2 31300 38049
0 22045 5 1 1 22044
0 22046 7 1 2 22043 22045
0 22047 5 1 1 22046
0 22048 7 1 2 33182 35449
0 22049 5 1 1 22048
0 22050 7 1 2 28798 29319
0 22051 5 1 1 22050
0 22052 7 1 2 22049 22051
0 22053 5 1 1 22052
0 22054 7 1 2 22047 22053
0 22055 5 1 1 22054
0 22056 7 1 2 27767 27831
0 22057 7 1 2 37567 22056
0 22058 5 1 1 22057
0 22059 7 1 2 33840 32670
0 22060 7 1 2 32664 22059
0 22061 7 1 2 32568 22060
0 22062 5 1 1 22061
0 22063 7 1 2 22058 22062
0 22064 7 1 2 22055 22063
0 22065 7 1 2 22041 22064
0 22066 7 1 2 22031 22065
0 22067 5 1 1 22066
0 22068 7 1 2 25247 22067
0 22069 5 1 1 22068
0 22070 7 1 2 24220 28793
0 22071 7 2 2 38050 22070
0 22072 7 1 2 32679 27832
0 22073 7 1 2 38345 22072
0 22074 5 1 1 22073
0 22075 7 1 2 22069 22074
0 22076 5 1 1 22075
0 22077 7 1 2 24523 22076
0 22078 5 1 1 22077
0 22079 7 1 2 30034 29591
0 22080 7 1 2 34363 22079
0 22081 7 1 2 38346 22080
0 22082 5 1 1 22081
0 22083 7 1 2 22078 22082
0 22084 5 1 1 22083
0 22085 7 1 2 36795 22084
0 22086 5 1 1 22085
0 22087 7 1 2 27541 38214
0 22088 5 1 1 22087
0 22089 7 1 2 30035 36299
0 22090 5 1 1 22089
0 22091 7 1 2 30793 30291
0 22092 5 1 1 22091
0 22093 7 1 2 22090 22092
0 22094 5 1 1 22093
0 22095 7 1 2 29267 22094
0 22096 5 1 1 22095
0 22097 7 1 2 23961 29964
0 22098 7 1 2 35350 22097
0 22099 5 1 1 22098
0 22100 7 1 2 22096 22099
0 22101 5 1 1 22100
0 22102 7 1 2 27094 22101
0 22103 5 1 1 22102
0 22104 7 1 2 22989 30059
0 22105 5 1 1 22104
0 22106 7 1 2 9215 22105
0 22107 5 1 1 22106
0 22108 7 1 2 38291 22107
0 22109 5 1 1 22108
0 22110 7 1 2 37590 38293
0 22111 5 1 1 22110
0 22112 7 1 2 22109 22111
0 22113 7 1 2 22103 22112
0 22114 5 1 1 22113
0 22115 7 1 2 29020 22114
0 22116 5 1 1 22115
0 22117 7 1 2 22088 22116
0 22118 5 1 1 22117
0 22119 7 1 2 26524 22118
0 22120 5 1 1 22119
0 22121 7 1 2 27515 37605
0 22122 5 1 1 22121
0 22123 7 1 2 22120 22122
0 22124 5 1 1 22123
0 22125 7 1 2 33397 22124
0 22126 5 1 1 22125
0 22127 7 1 2 22086 22126
0 22128 7 1 2 22015 22127
0 22129 5 1 1 22128
0 22130 7 1 2 23749 22129
0 22131 5 1 1 22130
0 22132 7 1 2 33412 22131
0 22133 5 1 1 22132
0 22134 7 1 2 36353 14070
0 22135 7 1 2 22133 22134
0 22136 7 1 2 21940 22135
0 22137 5 1 1 22136
0 22138 7 1 2 37164 19912
0 22139 5 1 1 22138
0 22140 7 1 2 24625 38247
0 22141 5 1 1 22140
0 22142 7 1 2 25517 36772
0 22143 7 1 2 37573 22142
0 22144 5 1 1 22143
0 22145 7 1 2 22141 22144
0 22146 5 2 1 22145
0 22147 7 1 2 29465 38347
0 22148 5 1 1 22147
0 22149 7 1 2 34859 38183
0 22150 5 1 1 22149
0 22151 7 1 2 22148 22150
0 22152 5 1 1 22151
0 22153 7 1 2 22525 22152
0 22154 5 1 1 22153
0 22155 7 1 2 22662 37391
0 22156 5 1 1 22155
0 22157 7 1 2 30655 38248
0 22158 5 1 1 22157
0 22159 7 1 2 22156 22158
0 22160 5 1 1 22159
0 22161 7 1 2 34608 22160
0 22162 5 1 1 22161
0 22163 7 1 2 22154 22162
0 22164 5 1 1 22163
0 22165 7 1 2 23858 22164
0 22166 5 1 1 22165
0 22167 7 1 2 38348 38195
0 22168 5 1 1 22167
0 22169 7 1 2 22166 22168
0 22170 5 1 1 22169
0 22171 7 1 2 25161 22170
0 22172 5 1 1 22171
0 22173 7 1 2 28809 38206
0 22174 7 1 2 29268 22173
0 22175 5 1 1 22174
0 22176 7 1 2 22172 22175
0 22177 5 1 1 22176
0 22178 7 1 2 24929 22177
0 22179 5 1 1 22178
0 22180 7 1 2 28810 38218
0 22181 7 1 2 33995 22180
0 22182 5 1 1 22181
0 22183 7 1 2 22179 22182
0 22184 5 1 1 22183
0 22185 7 1 2 24803 22184
0 22186 5 1 1 22185
0 22187 7 1 2 35861 35854
0 22188 7 1 2 29122 22187
0 22189 7 1 2 38288 22188
0 22190 7 1 2 33996 22189
0 22191 5 1 1 22190
0 22192 7 1 2 22186 22191
0 22193 5 1 1 22192
0 22194 7 1 2 24718 22193
0 22195 5 1 1 22194
0 22196 7 2 2 29021 38220
0 22197 7 1 2 30857 33997
0 22198 7 1 2 38349 22197
0 22199 5 1 1 22198
0 22200 7 1 2 22195 22199
0 22201 5 1 1 22200
0 22202 7 1 2 24389 22201
0 22203 5 1 1 22202
0 22204 7 2 2 34314 38350
0 22205 7 1 2 37610 38351
0 22206 5 1 1 22205
0 22207 7 1 2 22203 22206
0 22208 5 1 1 22207
0 22209 7 1 2 22139 22208
0 22210 5 1 1 22209
0 22211 7 1 2 37411 37322
0 22212 5 1 1 22211
0 22213 7 1 2 35877 38181
0 22214 5 1 1 22213
0 22215 7 1 2 34741 34570
0 22216 7 1 2 32209 22215
0 22217 7 1 2 38190 22216
0 22218 5 1 1 22217
0 22219 7 1 2 22214 22218
0 22220 5 1 1 22219
0 22221 7 1 2 22526 22220
0 22222 5 1 1 22221
0 22223 7 1 2 35372 38178
0 22224 5 1 1 22223
0 22225 7 1 2 22222 22224
0 22226 5 1 1 22225
0 22227 7 1 2 32641 22226
0 22228 5 1 1 22227
0 22229 7 1 2 27815 34684
0 22230 7 1 2 38229 22229
0 22231 7 1 2 37611 22230
0 22232 5 1 1 22231
0 22233 7 1 2 22228 22232
0 22234 5 1 1 22233
0 22235 7 1 2 23859 22234
0 22236 5 1 1 22235
0 22237 7 1 2 24719 38174
0 22238 5 1 1 22237
0 22239 7 1 2 37071 37699
0 22240 5 1 1 22239
0 22241 7 1 2 22238 22240
0 22242 5 1 1 22241
0 22243 7 1 2 30902 22242
0 22244 5 1 1 22243
0 22245 7 1 2 35184 36732
0 22246 5 1 1 22245
0 22247 7 1 2 22244 22246
0 22248 5 1 1 22247
0 22249 7 1 2 38196 22248
0 22250 5 1 1 22249
0 22251 7 1 2 22236 22250
0 22252 5 1 1 22251
0 22253 7 1 2 25162 22252
0 22254 5 1 1 22253
0 22255 7 1 2 27329 37743
0 22256 5 1 1 22255
0 22257 7 1 2 34146 31252
0 22258 5 1 1 22257
0 22259 7 1 2 22256 22258
0 22260 5 2 1 22259
0 22261 7 1 2 32642 36606
0 22262 7 1 2 38204 22261
0 22263 7 1 2 38353 22262
0 22264 5 1 1 22263
0 22265 7 1 2 22254 22264
0 22266 5 1 1 22265
0 22267 7 1 2 24930 22266
0 22268 5 1 1 22267
0 22269 7 1 2 27330 34820
0 22270 5 1 1 22269
0 22271 7 1 2 34147 36315
0 22272 5 1 1 22271
0 22273 7 1 2 22270 22272
0 22274 5 2 1 22273
0 22275 7 1 2 32709 27639
0 22276 7 1 2 38289 22275
0 22277 7 1 2 38355 22276
0 22278 5 1 1 22277
0 22279 7 1 2 22268 22278
0 22280 5 1 1 22279
0 22281 7 1 2 24804 22280
0 22282 5 1 1 22281
0 22283 7 1 2 28969 38221
0 22284 7 1 2 38356 22283
0 22285 5 1 1 22284
0 22286 7 1 2 22282 22285
0 22287 5 1 1 22286
0 22288 7 1 2 24390 22287
0 22289 5 1 1 22288
0 22290 7 1 2 38352 38354
0 22291 5 1 1 22290
0 22292 7 1 2 22289 22291
0 22293 5 1 1 22292
0 22294 7 1 2 22212 22293
0 22295 5 1 1 22294
0 22296 7 1 2 22210 22295
0 22297 7 1 2 22137 22296
0 22298 7 1 2 21360 22297
0 22299 7 1 2 21110 22298
0 22300 7 1 2 19041 22299
0 22301 7 1 2 17351 22300
0 22302 7 1 2 17336 22301
0 22303 5 1 1 22302
0 22304 7 1 2 43 22303
0 22305 5 1 1 22304
0 22306 7 1 2 13931 22305
3 49999 5 0 1 22306
