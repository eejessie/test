1 0 0 4 0
2 25 1 0
2 26 1 0
2 929 1 0
2 930 1 0
1 1 0 10 0
2 931 1 1
2 932 1 1
2 933 1 1
2 934 1 1
2 935 1 1
2 936 1 1
2 937 1 1
2 938 1 1
2 939 1 1
2 940 1 1
1 2 0 14 0
2 941 1 2
2 942 1 2
2 943 1 2
2 944 1 2
2 945 1 2
2 946 1 2
2 947 1 2
2 948 1 2
2 949 1 2
2 950 1 2
2 951 1 2
2 952 1 2
2 953 1 2
2 954 1 2
1 3 0 10 0
2 955 1 3
2 956 1 3
2 957 1 3
2 958 1 3
2 959 1 3
2 960 1 3
2 961 1 3
2 962 1 3
2 963 1 3
2 964 1 3
1 4 0 11 0
2 965 1 4
2 966 1 4
2 967 1 4
2 968 1 4
2 969 1 4
2 970 1 4
2 971 1 4
2 972 1 4
2 973 1 4
2 974 1 4
2 975 1 4
1 5 0 12 0
2 976 1 5
2 977 1 5
2 978 1 5
2 979 1 5
2 980 1 5
2 981 1 5
2 982 1 5
2 983 1 5
2 984 1 5
2 985 1 5
2 986 1 5
2 987 1 5
1 6 0 9 0
2 988 1 6
2 989 1 6
2 990 1 6
2 991 1 6
2 992 1 6
2 993 1 6
2 994 1 6
2 995 1 6
2 996 1 6
1 7 0 9 0
2 997 1 7
2 998 1 7
2 999 1 7
2 1000 1 7
2 1001 1 7
2 1002 1 7
2 1003 1 7
2 1004 1 7
2 1005 1 7
1 8 0 2 0
2 1006 1 8
2 1007 1 8
1 9 0 4 0
2 1008 1 9
2 1009 1 9
2 1010 1 9
2 1011 1 9
1 10 0 2 0
2 1012 1 10
2 1013 1 10
1 11 0 2 0
2 1014 1 11
2 1015 1 11
1 12 0 3 0
2 1016 1 12
2 1017 1 12
2 1018 1 12
1 13 0 2 0
2 1019 1 13
2 1020 1 13
1 14 0 2 0
2 1021 1 14
2 1022 1 14
1 15 0 3 0
2 1023 1 15
2 1024 1 15
2 1025 1 15
1 16 0 2 0
2 1026 1 16
2 1027 1 16
1 17 0 5 0
2 1028 1 17
2 1029 1 17
2 1030 1 17
2 1031 1 17
2 1032 1 17
1 18 0 2 0
2 1033 1 18
2 1034 1 18
1 19 0 2 0
2 1035 1 19
2 1036 1 19
1 20 0 3 0
2 1037 1 20
2 1038 1 20
2 1039 1 20
1 21 0 2 0
2 1040 1 21
2 1041 1 21
1 22 0 2 0
2 1042 1 22
2 1043 1 22
1 23 0 2 0
2 1044 1 23
2 1045 1 23
1 24 0 4 0
2 1046 1 24
2 1047 1 24
2 1048 1 24
2 1049 1 24
2 1050 1 27
2 1051 1 27
2 1052 1 27
2 1053 1 27
2 1054 1 27
2 1055 1 27
2 1056 1 27
2 1057 1 28
2 1058 1 28
2 1059 1 28
2 1060 1 28
2 1061 1 28
2 1062 1 28
2 1063 1 28
2 1064 1 28
2 1065 1 28
2 1066 1 28
2 1067 1 28
2 1068 1 28
2 1069 1 29
2 1070 1 29
2 1071 1 29
2 1072 1 29
2 1073 1 29
2 1074 1 29
2 1075 1 29
2 1076 1 29
2 1077 1 29
2 1078 1 30
2 1079 1 30
2 1080 1 30
2 1081 1 30
2 1082 1 30
2 1083 1 30
2 1084 1 30
2 1085 1 30
2 1086 1 31
2 1087 1 31
2 1088 1 31
2 1089 1 31
2 1090 1 31
2 1091 1 31
2 1092 1 31
2 1093 1 31
2 1094 1 32
2 1095 1 32
2 1096 1 32
2 1097 1 32
2 1098 1 32
2 1099 1 32
2 1100 1 32
2 1101 1 32
2 1102 1 32
2 1103 1 33
2 1104 1 33
2 1105 1 33
2 1106 1 33
2 1107 1 33
2 1108 1 33
2 1109 1 33
2 1110 1 33
2 1111 1 34
2 1112 1 34
2 1113 1 34
2 1114 1 34
2 1115 1 34
2 1116 1 36
2 1117 1 36
2 1118 1 36
2 1119 1 39
2 1120 1 39
2 1121 1 44
2 1122 1 44
2 1123 1 44
2 1124 1 47
2 1125 1 47
2 1126 1 50
2 1127 1 50
2 1128 1 51
2 1129 1 51
2 1130 1 51
2 1131 1 52
2 1132 1 52
2 1133 1 52
2 1134 1 52
2 1135 1 53
2 1136 1 53
2 1137 1 54
2 1138 1 54
2 1139 1 54
2 1140 1 54
2 1141 1 55
2 1142 1 55
2 1143 1 56
2 1144 1 56
2 1145 1 56
2 1146 1 56
2 1147 1 56
2 1148 1 57
2 1149 1 57
2 1150 1 57
2 1151 1 57
2 1152 1 58
2 1153 1 58
2 1154 1 58
2 1155 1 58
2 1156 1 59
2 1157 1 59
2 1158 1 59
2 1159 1 60
2 1160 1 60
2 1161 1 60
2 1162 1 60
2 1163 1 61
2 1164 1 61
2 1165 1 61
2 1166 1 61
2 1167 1 61
2 1168 1 61
2 1169 1 61
2 1170 1 63
2 1171 1 63
2 1172 1 67
2 1173 1 67
2 1174 1 67
2 1175 1 72
2 1176 1 72
2 1177 1 72
2 1178 1 72
2 1179 1 72
2 1180 1 72
2 1181 1 72
2 1182 1 72
2 1183 1 72
2 1184 1 73
2 1185 1 73
2 1186 1 73
2 1187 1 74
2 1188 1 74
2 1189 1 74
2 1190 1 74
2 1191 1 77
2 1192 1 77
2 1193 1 77
2 1194 1 78
2 1195 1 78
2 1196 1 78
2 1197 1 78
2 1198 1 81
2 1199 1 81
2 1200 1 84
2 1201 1 84
2 1202 1 84
2 1203 1 84
2 1204 1 84
2 1205 1 84
2 1206 1 84
2 1207 1 88
2 1208 1 88
2 1209 1 88
2 1210 1 92
2 1211 1 92
2 1212 1 92
2 1213 1 92
2 1214 1 92
2 1215 1 92
2 1216 1 92
2 1217 1 92
2 1218 1 92
2 1219 1 92
2 1220 1 92
2 1221 1 97
2 1222 1 97
2 1223 1 97
2 1224 1 97
2 1225 1 97
2 1226 1 97
2 1227 1 97
2 1228 1 97
2 1229 1 98
2 1230 1 98
2 1231 1 98
2 1232 1 98
2 1233 1 98
2 1234 1 99
2 1235 1 99
2 1236 1 99
2 1237 1 101
2 1238 1 101
2 1239 1 101
2 1240 1 101
2 1241 1 104
2 1242 1 104
2 1243 1 104
2 1244 1 105
2 1245 1 105
2 1246 1 105
2 1247 1 107
2 1248 1 107
2 1249 1 107
2 1250 1 107
2 1251 1 114
2 1252 1 114
2 1253 1 114
2 1254 1 114
2 1255 1 114
2 1256 1 114
2 1257 1 114
2 1258 1 114
2 1259 1 114
2 1260 1 116
2 1261 1 116
2 1262 1 116
2 1263 1 116
2 1264 1 117
2 1265 1 117
2 1266 1 118
2 1267 1 118
2 1268 1 118
2 1269 1 118
2 1270 1 121
2 1271 1 121
2 1272 1 121
2 1273 1 121
2 1274 1 122
2 1275 1 122
2 1276 1 122
2 1277 1 123
2 1278 1 123
2 1279 1 130
2 1280 1 130
2 1281 1 130
2 1282 1 130
2 1283 1 147
2 1284 1 147
2 1285 1 147
2 1286 1 150
2 1287 1 150
2 1288 1 176
2 1289 1 176
2 1290 1 176
2 1291 1 180
2 1292 1 180
2 1293 1 180
2 1294 1 180
2 1295 1 180
2 1296 1 181
2 1297 1 181
2 1298 1 181
2 1299 1 181
2 1300 1 185
2 1301 1 185
2 1302 1 185
2 1303 1 185
2 1304 1 196
2 1305 1 196
2 1306 1 196
2 1307 1 196
2 1308 1 207
2 1309 1 207
2 1310 1 207
2 1311 1 207
2 1312 1 218
2 1313 1 218
2 1314 1 218
2 1315 1 218
2 1316 1 219
2 1317 1 219
2 1318 1 221
2 1319 1 221
2 1320 1 236
2 1321 1 236
2 1322 1 240
2 1323 1 240
2 1324 1 240
2 1325 1 240
2 1326 1 240
2 1327 1 245
2 1328 1 245
2 1329 1 245
2 1330 1 249
2 1331 1 249
2 1332 1 250
2 1333 1 250
2 1334 1 250
2 1335 1 250
2 1336 1 250
2 1337 1 250
2 1338 1 251
2 1339 1 251
2 1340 1 251
2 1341 1 251
2 1342 1 251
2 1343 1 251
2 1344 1 252
2 1345 1 252
2 1346 1 253
2 1347 1 253
2 1348 1 256
2 1349 1 256
2 1350 1 256
2 1351 1 257
2 1352 1 257
2 1353 1 259
2 1354 1 259
2 1355 1 260
2 1356 1 260
2 1357 1 262
2 1358 1 262
2 1359 1 265
2 1360 1 265
2 1361 1 269
2 1362 1 269
2 1363 1 272
2 1364 1 272
2 1365 1 272
2 1366 1 273
2 1367 1 273
2 1368 1 276
2 1369 1 276
2 1370 1 276
2 1371 1 276
2 1372 1 276
2 1373 1 277
2 1374 1 277
2 1375 1 277
2 1376 1 278
2 1377 1 278
2 1378 1 278
2 1379 1 278
2 1380 1 278
2 1381 1 278
2 1382 1 278
2 1383 1 278
2 1384 1 279
2 1385 1 279
2 1386 1 280
2 1387 1 280
2 1388 1 283
2 1389 1 283
2 1390 1 284
2 1391 1 284
2 1392 1 284
2 1393 1 284
2 1394 1 288
2 1395 1 288
2 1396 1 288
2 1397 1 288
2 1398 1 288
2 1399 1 288
2 1400 1 289
2 1401 1 289
2 1402 1 289
2 1403 1 300
2 1404 1 300
2 1405 1 302
2 1406 1 302
2 1407 1 302
2 1408 1 309
2 1409 1 309
2 1410 1 309
2 1411 1 309
2 1412 1 311
2 1413 1 311
2 1414 1 312
2 1415 1 312
2 1416 1 312
2 1417 1 312
2 1418 1 319
2 1419 1 319
2 1420 1 319
2 1421 1 319
2 1422 1 319
2 1423 1 327
2 1424 1 327
2 1425 1 327
2 1426 1 339
2 1427 1 339
2 1428 1 340
2 1429 1 340
2 1430 1 340
2 1431 1 340
2 1432 1 341
2 1433 1 341
2 1434 1 341
2 1435 1 342
2 1436 1 342
2 1437 1 342
2 1438 1 342
2 1439 1 344
2 1440 1 344
2 1441 1 346
2 1442 1 346
2 1443 1 346
2 1444 1 348
2 1445 1 348
2 1446 1 348
2 1447 1 348
2 1448 1 356
2 1449 1 356
2 1450 1 372
2 1451 1 372
2 1452 1 385
2 1453 1 385
2 1454 1 401
2 1455 1 401
2 1456 1 401
2 1457 1 404
2 1458 1 404
2 1459 1 405
2 1460 1 405
2 1461 1 413
2 1462 1 413
2 1463 1 413
2 1464 1 427
2 1465 1 427
2 1466 1 432
2 1467 1 432
2 1468 1 432
2 1469 1 432
2 1470 1 432
2 1471 1 432
2 1472 1 441
2 1473 1 441
2 1474 1 441
2 1475 1 451
2 1476 1 451
2 1477 1 451
2 1478 1 452
2 1479 1 452
2 1480 1 452
2 1481 1 468
2 1482 1 468
2 1483 1 504
2 1484 1 504
2 1485 1 507
2 1486 1 507
2 1487 1 540
2 1488 1 540
2 1489 1 540
2 1490 1 541
2 1491 1 541
2 1492 1 541
2 1493 1 574
2 1494 1 574
2 1495 1 605
2 1496 1 605
2 1497 1 605
2 1498 1 606
2 1499 1 606
2 1500 1 607
2 1501 1 607
2 1502 1 607
2 1503 1 607
2 1504 1 608
2 1505 1 608
2 1506 1 614
2 1507 1 614
2 1508 1 616
2 1509 1 616
2 1510 1 647
2 1511 1 647
2 1512 1 647
2 1513 1 647
2 1514 1 648
2 1515 1 648
2 1516 1 648
2 1517 1 648
2 1518 1 648
2 1519 1 649
2 1520 1 649
2 1521 1 651
2 1522 1 651
2 1523 1 651
2 1524 1 662
2 1525 1 662
2 1526 1 663
2 1527 1 663
2 1528 1 663
2 1529 1 663
2 1530 1 664
2 1531 1 664
2 1532 1 664
2 1533 1 664
2 1534 1 664
2 1535 1 674
2 1536 1 674
2 1537 1 674
2 1538 1 674
2 1539 1 674
2 1540 1 744
2 1541 1 744
2 1542 1 750
2 1543 1 750
2 1544 1 759
2 1545 1 759
2 1546 1 759
2 1547 1 767
2 1548 1 767
2 1549 1 775
2 1550 1 775
2 1551 1 778
2 1552 1 778
2 1553 1 788
2 1554 1 788
2 1555 1 833
2 1556 1 833
2 1557 1 836
2 1558 1 836
2 1559 1 844
2 1560 1 844
2 1561 1 853
2 1562 1 853
2 1563 1 883
2 1564 1 883
2 1565 1 887
2 1566 1 887
0 27 5 7 1 25
0 28 5 12 1 931
0 29 5 9 1 941
0 30 5 8 1 955
0 31 5 8 1 965
0 32 5 9 1 976
0 33 5 8 1 988
0 34 5 5 1 997
0 35 5 1 1 1006
0 36 5 3 1 1008
0 37 5 1 1 1012
0 38 5 1 1 1014
0 39 5 2 1 1016
0 40 5 1 1 1019
0 41 5 1 1 1021
0 42 5 1 1 1023
0 43 5 1 1 1026
0 44 5 3 1 1028
0 45 5 1 1 1033
0 46 5 1 1 1035
0 47 5 2 1 1037
0 48 5 1 1 1040
0 49 5 1 1 1042
0 50 5 2 1 1044
0 51 5 3 1 1046
0 52 7 4 2 1119 1038
0 53 5 2 1 1131
0 54 7 4 2 1017 1124
0 55 5 2 1 1137
0 56 7 5 2 1135 1141
0 57 7 4 2 1020 48
0 58 5 4 1 1148
0 59 7 3 2 40 1041
0 60 5 4 1 1156
0 61 7 7 2 1152 1159
0 62 5 1 1 1163
0 63 7 2 2 1024 1126
0 64 5 1 1 1170
0 65 7 1 2 1047 1171
0 66 5 1 1 65
0 67 7 3 2 42 1045
0 68 5 1 1 1172
0 69 7 1 2 1128 1173
0 70 5 1 1 69
0 71 7 1 2 66 70
0 72 5 9 1 71
0 73 7 3 2 1022 49
0 74 5 4 1 1184
0 75 7 1 2 1111 1187
0 76 5 1 1 75
0 77 7 3 2 41 1043
0 78 5 4 1 1191
0 79 7 1 2 998 1194
0 80 5 1 1 79
0 81 7 2 2 76 80
0 82 7 1 2 1175 1198
0 83 5 1 1 82
0 84 7 7 2 1112 1129
0 85 5 1 1 1200
0 86 7 1 2 1188 85
0 87 5 1 1 86
0 88 7 3 2 999 1048
0 89 5 1 1 1207
0 90 7 1 2 1195 89
0 91 5 1 1 90
0 92 7 11 2 64 68
0 93 7 1 2 91 1210
0 94 7 1 2 87 93
0 95 5 1 1 94
0 96 7 1 2 83 95
0 97 5 8 1 96
0 98 7 5 2 38 1036
0 99 5 3 1 1229
0 100 7 1 2 1086 1094
0 101 7 4 2 989 100
0 102 7 1 2 1230 1237
0 103 5 1 1 102
0 104 7 3 2 1015 46
0 105 5 3 1 1241
0 106 7 1 2 966 977
0 107 7 4 2 1103 106
0 108 7 1 2 1242 1247
0 109 5 1 1 108
0 110 7 1 2 103 109
0 111 5 1 1 110
0 112 7 1 2 1221 111
0 113 5 1 1 112
0 114 7 9 2 1189 1196
0 115 5 1 1 1251
0 116 7 4 2 967 1243
0 117 7 2 2 978 990
0 118 7 4 2 1113 1264
0 119 7 1 2 1260 1266
0 120 5 1 1 119
0 121 7 4 2 1095 1104
0 122 7 3 2 1087 1270
0 123 7 2 2 1231 1274
0 124 7 1 2 1000 1277
0 125 5 1 1 124
0 126 7 1 2 120 125
0 127 5 1 1 126
0 128 7 1 2 1176 127
0 129 5 1 1 128
0 130 7 4 2 1208 1265
0 131 7 1 2 1261 1279
0 132 5 1 1 131
0 133 7 1 2 1201 1278
0 134 5 1 1 133
0 135 7 1 2 132 134
0 136 5 1 1 135
0 137 7 1 2 1211 136
0 138 5 1 1 137
0 139 7 1 2 129 138
0 140 5 1 1 139
0 141 7 1 2 1252 140
0 142 5 1 1 141
0 143 7 1 2 113 142
0 144 5 1 1 143
0 145 7 1 2 1164 144
0 146 5 1 1 145
0 147 7 3 2 1105 1157
0 148 7 1 2 1202 1283
0 149 5 1 1 148
0 150 7 2 2 991 1149
0 151 7 1 2 1209 1286
0 152 5 1 1 151
0 153 7 1 2 149 152
0 154 5 1 1 153
0 155 7 1 2 1212 154
0 156 5 1 1 155
0 157 7 1 2 992 1114
0 158 5 1 1 157
0 159 7 1 2 1160 158
0 160 5 1 1 159
0 161 7 1 2 1106 1001
0 162 5 1 1 161
0 163 7 1 2 1153 162
0 164 5 1 1 163
0 165 7 1 2 160 164
0 166 7 1 2 1177 165
0 167 5 1 1 166
0 168 7 1 2 156 167
0 169 5 1 1 168
0 170 7 1 2 1253 169
0 171 5 1 1 170
0 172 7 1 2 1107 1154
0 173 5 1 1 172
0 174 7 1 2 993 1161
0 175 5 1 1 174
0 176 7 3 2 173 175
0 177 7 1 2 1222 1288
0 178 5 1 1 177
0 179 7 1 2 171 178
0 180 5 5 1 179
0 181 7 4 2 968 1096
0 182 5 1 1 1296
0 183 7 1 2 1234 182
0 184 5 1 1 183
0 185 7 4 2 1088 979
0 186 5 1 1 1300
0 187 7 1 2 1244 186
0 188 5 1 1 187
0 189 7 1 2 184 188
0 190 7 1 2 1291 189
0 191 5 1 1 190
0 192 7 1 2 146 191
0 193 5 1 1 192
0 194 7 1 2 1143 193
0 195 5 1 1 194
0 196 7 4 2 1203 1271
0 197 7 1 2 1132 1304
0 198 5 1 1 197
0 199 7 1 2 1138 1280
0 200 5 1 1 199
0 201 7 1 2 198 200
0 202 5 1 1 201
0 203 7 1 2 1213 202
0 204 5 1 1 203
0 205 7 1 2 1139 1267
0 206 5 1 1 205
0 207 7 4 2 1002 1272
0 208 7 1 2 1133 1308
0 209 5 1 1 208
0 210 7 1 2 206 209
0 211 5 1 1 210
0 212 7 1 2 1178 211
0 213 5 1 1 212
0 214 7 1 2 204 213
0 215 5 1 1 214
0 216 7 1 2 1254 215
0 217 5 1 1 216
0 218 7 4 2 1097 994
0 219 7 2 2 1134 1312
0 220 5 1 1 1316
0 221 7 2 2 980 1108
0 222 7 1 2 1140 1318
0 223 5 1 1 222
0 224 7 1 2 220 223
0 225 5 1 1 224
0 226 7 1 2 1223 225
0 227 5 1 1 226
0 228 7 1 2 217 227
0 229 5 1 1 228
0 230 7 1 2 1165 229
0 231 5 1 1 230
0 232 7 1 2 1098 1142
0 233 5 1 1 232
0 234 7 1 2 981 1136
0 235 5 1 1 234
0 236 7 2 2 233 235
0 237 7 1 2 1292 1320
0 238 5 1 1 237
0 239 7 1 2 231 238
0 240 5 5 1 239
0 241 7 1 2 1089 1245
0 242 5 1 1 241
0 243 7 1 2 969 1235
0 244 5 1 1 243
0 245 7 3 2 242 244
0 246 7 1 2 1322 1327
0 247 5 1 1 246
0 248 7 1 2 195 247
0 249 5 2 1 248
0 250 7 6 2 1007 43
0 251 5 6 1 1332
0 252 7 2 2 1057 1116
0 253 5 2 1 1344
0 254 7 1 2 1333 1345
0 255 5 1 1 254
0 256 7 3 2 35 1027
0 257 5 2 1 1348
0 258 7 1 2 1121 1351
0 259 5 2 1 258
0 260 7 2 2 932 1009
0 261 5 1 1 1355
0 262 7 2 2 1346 261
0 263 5 1 1 1357
0 264 7 1 2 1010 1029
0 265 7 2 2 1349 264
0 266 5 1 1 1359
0 267 7 1 2 263 266
0 268 5 1 1 267
0 269 7 2 2 1353 268
0 270 5 1 1 1361
0 271 7 1 2 255 270
0 272 5 3 1 271
0 273 7 2 2 1069 956
0 274 7 1 2 1363 1366
0 275 5 1 1 274
0 276 7 5 2 1011 1122
0 277 5 3 1 1368
0 278 7 8 2 1117 1030
0 279 5 2 1 1376
0 280 7 2 2 933 1384
0 281 5 1 1 1386
0 282 7 1 2 1373 281
0 283 5 2 1 282
0 284 7 4 2 1334 1388
0 285 5 1 1 1390
0 286 7 1 2 1078 285
0 287 5 1 1 286
0 288 7 6 2 1350 1377
0 289 7 3 2 1058 1394
0 290 5 1 1 1400
0 291 7 1 2 957 290
0 292 5 1 1 291
0 293 7 1 2 942 292
0 294 7 1 2 287 293
0 295 5 1 1 294
0 296 7 1 2 275 295
0 297 5 1 1 296
0 298 7 1 2 1050 297
0 299 5 1 1 298
0 300 7 2 2 1367 1378
0 301 5 1 1 1403
0 302 7 3 2 943 1079
0 303 7 1 2 1369 1405
0 304 5 1 1 303
0 305 7 1 2 301 304
0 306 5 1 1 305
0 307 7 1 2 934 306
0 308 5 1 1 307
0 309 7 4 2 1374 1385
0 310 5 1 1 1408
0 311 7 2 2 1059 1070
0 312 7 4 2 1409 1412
0 313 7 1 2 958 1414
0 314 5 1 1 313
0 315 7 1 2 308 314
0 316 5 1 1 315
0 317 7 1 2 1338 316
0 318 5 1 1 317
0 319 7 5 2 26 1352
0 320 7 1 2 1060 1404
0 321 5 1 1 320
0 322 7 1 2 935 1410
0 323 5 1 1 322
0 324 7 1 2 1061 1370
0 325 5 1 1 324
0 326 7 1 2 323 325
0 327 5 3 1 326
0 328 7 1 2 1406 1423
0 329 5 1 1 328
0 330 7 1 2 321 329
0 331 5 1 1 330
0 332 7 1 2 1418 331
0 333 5 1 1 332
0 334 7 1 2 318 333
0 335 7 1 2 299 334
0 336 5 1 1 335
0 337 7 1 2 1330 336
0 338 5 1 1 337
0 339 7 2 2 1236 1246
0 340 7 4 2 1080 1090
0 341 7 3 2 1071 1428
0 342 7 4 2 1379 1432
0 343 5 1 1 1435
0 344 7 2 2 1305 1436
0 345 5 1 1 1439
0 346 7 3 2 959 970
0 347 7 1 2 944 1371
0 348 7 4 2 1441 347
0 349 5 1 1 1444
0 350 7 1 2 1281 1445
0 351 5 1 1 350
0 352 7 1 2 345 351
0 353 5 1 1 352
0 354 7 1 2 936 353
0 355 5 1 1 354
0 356 7 2 2 1415 1429
0 357 7 1 2 1306 1448
0 358 5 1 1 357
0 359 7 1 2 355 358
0 360 5 1 1 359
0 361 7 1 2 1214 360
0 362 5 1 1 361
0 363 7 1 2 1268 1446
0 364 5 1 1 363
0 365 7 1 2 1309 1437
0 366 5 1 1 365
0 367 7 1 2 364 366
0 368 5 1 1 367
0 369 7 1 2 937 368
0 370 5 1 1 369
0 371 7 1 2 1062 1310
0 372 7 2 2 1433 371
0 373 7 1 2 1411 1450
0 374 5 1 1 373
0 375 7 1 2 370 374
0 376 5 1 1 375
0 377 7 1 2 1179 376
0 378 5 1 1 377
0 379 7 1 2 362 378
0 380 5 1 1 379
0 381 7 1 2 1255 380
0 382 5 1 1 381
0 383 7 1 2 1319 1447
0 384 5 1 1 383
0 385 7 2 2 1313 1438
0 386 5 1 1 1452
0 387 7 1 2 384 386
0 388 5 1 1 387
0 389 7 1 2 938 388
0 390 5 1 1 389
0 391 7 1 2 1314 1449
0 392 5 1 1 391
0 393 7 1 2 390 392
0 394 5 1 1 393
0 395 7 1 2 1224 394
0 396 5 1 1 395
0 397 7 1 2 382 396
0 398 5 1 1 397
0 399 7 1 2 1339 398
0 400 5 1 1 399
0 401 7 3 2 1269 1442
0 402 7 1 2 1391 1454
0 403 5 1 1 402
0 404 7 2 2 1063 1081
0 405 7 2 2 1275 1457
0 406 7 1 2 1003 1395
0 407 7 1 2 1459 406
0 408 5 1 1 407
0 409 7 1 2 403 408
0 410 5 1 1 409
0 411 7 1 2 1180 410
0 412 5 1 1 411
0 413 7 3 2 1282 1443
0 414 7 1 2 1392 1461
0 415 5 1 1 414
0 416 7 1 2 1204 1396
0 417 7 1 2 1460 416
0 418 5 1 1 417
0 419 7 1 2 415 418
0 420 5 1 1 419
0 421 7 1 2 1215 420
0 422 5 1 1 421
0 423 7 1 2 412 422
0 424 5 1 1 423
0 425 7 1 2 945 424
0 426 5 1 1 425
0 427 7 2 2 1004 1181
0 428 5 1 1 1464
0 429 7 1 2 1216 1205
0 430 5 1 1 429
0 431 7 1 2 428 430
0 432 5 6 1 431
0 433 7 1 2 1273 1434
0 434 7 1 2 1364 433
0 435 7 1 2 1466 434
0 436 5 1 1 435
0 437 7 1 2 426 436
0 438 5 1 1 437
0 439 7 1 2 1256 438
0 440 5 1 1 439
0 441 7 3 2 960 1393
0 442 7 1 2 1248 1472
0 443 5 1 1 442
0 444 7 1 2 1238 1458
0 445 7 1 2 1397 444
0 446 5 1 1 445
0 447 7 1 2 443 446
0 448 5 1 1 447
0 449 7 1 2 946 448
0 450 5 1 1 449
0 451 7 3 2 1072 1082
0 452 7 3 2 1365 1475
0 453 5 1 1 1478
0 454 7 1 2 1239 1479
0 455 5 1 1 454
0 456 7 1 2 450 455
0 457 5 1 1 456
0 458 7 1 2 1225 457
0 459 5 1 1 458
0 460 7 1 2 440 459
0 461 5 1 1 460
0 462 7 1 2 1051 461
0 463 5 1 1 462
0 464 7 1 2 400 463
0 465 5 1 1 464
0 466 7 1 2 1166 465
0 467 5 1 1 466
0 468 7 2 2 982 1430
0 469 7 1 2 1401 1481
0 470 5 1 1 469
0 471 7 1 2 1297 1473
0 472 5 1 1 471
0 473 7 1 2 470 472
0 474 5 1 1 473
0 475 7 1 2 947 474
0 476 5 1 1 475
0 477 7 1 2 1301 1480
0 478 5 1 1 477
0 479 7 1 2 476 478
0 480 5 1 1 479
0 481 7 1 2 1052 480
0 482 5 1 1 481
0 483 7 1 2 1099 349
0 484 5 1 1 483
0 485 7 1 2 983 343
0 486 5 1 1 485
0 487 7 1 2 939 486
0 488 7 1 2 484 487
0 489 5 1 1 488
0 490 7 1 2 1416 1482
0 491 5 1 1 490
0 492 7 1 2 489 491
0 493 5 1 1 492
0 494 7 1 2 1340 493
0 495 5 1 1 494
0 496 7 1 2 482 495
0 497 5 1 1 496
0 498 7 1 2 1293 497
0 499 5 1 1 498
0 500 7 1 2 467 499
0 501 5 1 1 500
0 502 7 1 2 1144 501
0 503 5 1 1 502
0 504 7 2 2 971 1380
0 505 7 1 2 1476 1483
0 506 5 1 1 505
0 507 7 2 2 948 1091
0 508 7 1 2 961 1372
0 509 7 1 2 1485 508
0 510 5 1 1 509
0 511 7 1 2 506 510
0 512 5 1 1 511
0 513 7 1 2 940 512
0 514 5 1 1 513
0 515 7 1 2 1083 972
0 516 7 1 2 1417 515
0 517 5 1 1 516
0 518 7 1 2 514 517
0 519 5 1 1 518
0 520 7 1 2 1341 519
0 521 5 1 1 520
0 522 7 1 2 1402 1407
0 523 5 1 1 522
0 524 7 1 2 453 523
0 525 5 1 1 524
0 526 7 1 2 973 525
0 527 5 1 1 526
0 528 7 1 2 1474 1486
0 529 5 1 1 528
0 530 7 1 2 527 529
0 531 5 1 1 530
0 532 7 1 2 1053 531
0 533 5 1 1 532
0 534 7 1 2 521 533
0 535 5 1 1 534
0 536 7 1 2 1323 535
0 537 5 1 1 536
0 538 7 1 2 1064 1453
0 539 5 1 1 538
0 540 7 3 2 949 1424
0 541 7 3 2 962 1487
0 542 7 1 2 1249 1490
0 543 5 1 1 542
0 544 7 1 2 539 543
0 545 5 1 1 544
0 546 7 1 2 1226 545
0 547 5 1 1 546
0 548 7 1 2 1065 1440
0 549 5 1 1 548
0 550 7 1 2 1462 1488
0 551 5 1 1 550
0 552 7 1 2 549 551
0 553 5 1 1 552
0 554 7 1 2 1217 553
0 555 5 1 1 554
0 556 7 1 2 1455 1489
0 557 5 1 1 556
0 558 7 1 2 1381 1451
0 559 5 1 1 558
0 560 7 1 2 557 559
0 561 5 1 1 560
0 562 7 1 2 1182 561
0 563 5 1 1 562
0 564 7 1 2 555 563
0 565 5 1 1 564
0 566 7 1 2 1257 565
0 567 5 1 1 566
0 568 7 1 2 547 567
0 569 5 1 1 568
0 570 7 1 2 1167 569
0 571 5 1 1 570
0 572 7 1 2 1298 1491
0 573 5 1 1 572
0 574 7 2 2 1066 1477
0 575 7 1 2 1302 1382
0 576 7 1 2 1493 575
0 577 5 1 1 576
0 578 7 1 2 573 577
0 579 5 1 1 578
0 580 7 1 2 1294 579
0 581 5 1 1 580
0 582 7 1 2 571 581
0 583 5 1 1 582
0 584 7 1 2 1145 583
0 585 5 1 1 584
0 586 7 1 2 1092 1492
0 587 5 1 1 586
0 588 7 1 2 1484 1494
0 589 5 1 1 588
0 590 7 1 2 587 589
0 591 5 1 1 590
0 592 7 1 2 1324 591
0 593 5 1 1 592
0 594 7 1 2 585 593
0 595 5 1 1 594
0 596 7 1 2 1419 595
0 597 5 1 1 596
0 598 7 1 2 537 597
0 599 7 1 2 503 598
0 600 5 1 1 599
0 601 7 1 2 1426 600
0 602 5 1 1 601
0 603 7 1 2 338 602
0 604 5 1 1 603
0 605 7 3 2 37 1034
0 606 5 2 1 1495
0 607 7 4 2 1013 45
0 608 5 2 1 1500
0 609 7 1 2 1498 1504
0 610 7 1 2 604 609
0 611 5 1 1 610
0 612 7 1 2 1073 1389
0 613 5 1 1 612
0 614 7 2 2 1067 950
0 615 7 1 2 1118 1506
0 616 5 2 1 615
0 617 7 1 2 613 1508
0 618 5 1 1 617
0 619 7 1 2 1335 618
0 620 5 1 1 619
0 621 7 1 2 951 1362
0 622 5 1 1 621
0 623 7 1 2 620 622
0 624 5 1 1 623
0 625 7 1 2 1054 624
0 626 5 1 1 625
0 627 7 1 2 1074 1425
0 628 5 1 1 627
0 629 7 1 2 1383 1507
0 630 5 1 1 629
0 631 7 1 2 628 630
0 632 5 1 1 631
0 633 7 1 2 1420 632
0 634 5 1 1 633
0 635 7 1 2 1068 310
0 636 5 1 1 635
0 637 7 1 2 952 1387
0 638 5 1 1 637
0 639 7 1 2 1075 1375
0 640 5 1 1 639
0 641 7 1 2 1342 640
0 642 7 1 2 638 641
0 643 7 1 2 636 642
0 644 5 1 1 643
0 645 7 1 2 634 644
0 646 7 1 2 626 645
0 647 5 4 1 646
0 648 7 5 2 963 1501
0 649 7 2 2 1093 1514
0 650 5 1 1 1519
0 651 7 3 2 1084 1496
0 652 7 1 2 974 1521
0 653 5 1 1 652
0 654 7 1 2 650 653
0 655 5 1 1 654
0 656 7 1 2 1510 655
0 657 5 1 1 656
0 658 7 1 2 1085 1505
0 659 5 1 1 658
0 660 7 1 2 964 1499
0 661 5 1 1 660
0 662 7 2 2 659 661
0 663 7 4 2 1398 1524
0 664 7 5 2 1055 1413
0 665 7 1 2 975 1530
0 666 7 1 2 1526 665
0 667 5 1 1 666
0 668 7 1 2 657 667
0 669 5 1 1 668
0 670 7 1 2 1325 669
0 671 5 1 1 670
0 672 7 1 2 1299 1515
0 673 5 1 1 672
0 674 7 5 2 1431 1497
0 675 7 1 2 984 1535
0 676 5 1 1 675
0 677 7 1 2 673 676
0 678 5 1 1 677
0 679 7 1 2 1511 678
0 680 5 1 1 679
0 681 7 1 2 1303 1531
0 682 7 1 2 1527 681
0 683 5 1 1 682
0 684 7 1 2 680 683
0 685 5 1 1 684
0 686 7 1 2 1295 685
0 687 5 1 1 686
0 688 7 1 2 1463 1502
0 689 5 1 1 688
0 690 7 1 2 1307 1536
0 691 5 1 1 690
0 692 7 1 2 689 691
0 693 5 1 1 692
0 694 7 1 2 1218 693
0 695 5 1 1 694
0 696 7 1 2 1311 1537
0 697 5 1 1 696
0 698 7 1 2 1456 1503
0 699 5 1 1 698
0 700 7 1 2 697 699
0 701 5 1 1 700
0 702 7 1 2 1183 701
0 703 5 1 1 702
0 704 7 1 2 695 703
0 705 5 1 1 704
0 706 7 1 2 1512 705
0 707 5 1 1 706
0 708 7 1 2 1276 1532
0 709 7 1 2 1528 708
0 710 7 1 2 1467 709
0 711 5 1 1 710
0 712 7 1 2 707 711
0 713 5 1 1 712
0 714 7 1 2 1258 713
0 715 5 1 1 714
0 716 7 1 2 1250 1516
0 717 5 1 1 716
0 718 7 1 2 1315 1538
0 719 5 1 1 718
0 720 7 1 2 717 719
0 721 5 1 1 720
0 722 7 1 2 1513 721
0 723 5 1 1 722
0 724 7 1 2 1240 1533
0 725 7 1 2 1529 724
0 726 5 1 1 725
0 727 7 1 2 723 726
0 728 5 1 1 727
0 729 7 1 2 1227 728
0 730 5 1 1 729
0 731 7 1 2 715 730
0 732 5 1 1 731
0 733 7 1 2 1168 732
0 734 5 1 1 733
0 735 7 1 2 687 734
0 736 5 1 1 735
0 737 7 1 2 1146 736
0 738 5 1 1 737
0 739 7 1 2 671 738
0 740 5 1 1 739
0 741 7 1 2 1427 740
0 742 5 1 1 741
0 743 7 1 2 985 1018
0 744 7 2 2 1125 743
0 745 7 1 2 1284 1468
0 746 5 1 1 745
0 747 7 1 2 1005 1219
0 748 5 1 1 747
0 749 7 1 2 1115 1025
0 750 7 2 2 1127 749
0 751 5 1 1 1542
0 752 7 1 2 748 751
0 753 5 1 1 752
0 754 7 1 2 1049 753
0 755 5 1 1 754
0 756 7 1 2 1174 1206
0 757 5 1 1 756
0 758 7 1 2 755 757
0 759 5 3 1 758
0 760 7 1 2 1287 1544
0 761 5 1 1 760
0 762 7 1 2 746 761
0 763 5 1 1 762
0 764 7 1 2 1540 763
0 765 5 1 1 764
0 766 7 1 2 1100 1120
0 767 7 2 2 1039 766
0 768 7 1 2 1289 1547
0 769 7 1 2 1469 768
0 770 5 1 1 769
0 771 7 1 2 765 770
0 772 5 1 1 771
0 773 7 1 2 1259 772
0 774 5 1 1 773
0 775 7 2 2 1109 1192
0 776 5 1 1 1549
0 777 7 1 2 1110 1190
0 778 5 2 1 777
0 779 7 1 2 1197 1551
0 780 5 1 1 779
0 781 7 1 2 776 780
0 782 7 1 2 1470 781
0 783 5 1 1 782
0 784 7 1 2 995 1185
0 785 7 1 2 1545 784
0 786 5 1 1 785
0 787 7 1 2 783 786
0 788 5 2 1 787
0 789 7 1 2 1169 1321
0 790 7 1 2 1553 789
0 791 5 1 1 790
0 792 7 1 2 1290 1541
0 793 5 1 1 792
0 794 7 1 2 1150 1317
0 795 5 1 1 794
0 796 7 1 2 793 795
0 797 5 1 1 796
0 798 7 1 2 1228 797
0 799 5 1 1 798
0 800 7 1 2 1199 1220
0 801 5 1 1 800
0 802 7 1 2 1193 1543
0 803 5 1 1 802
0 804 7 1 2 801 803
0 805 5 1 1 804
0 806 7 1 2 1130 805
0 807 5 1 1 806
0 808 7 1 2 1186 1465
0 809 5 1 1 808
0 810 7 1 2 807 809
0 811 5 1 1 810
0 812 7 1 2 1285 1548
0 813 7 1 2 811 812
0 814 5 1 1 813
0 815 7 1 2 799 814
0 816 7 1 2 791 815
0 817 7 1 2 774 816
0 818 5 1 1 817
0 819 7 1 2 1232 1539
0 820 7 1 2 818 819
0 821 5 1 1 820
0 822 7 1 2 1471 1550
0 823 5 1 1 822
0 824 7 1 2 996 115
0 825 5 1 1 824
0 826 7 1 2 1552 825
0 827 7 1 2 1546 826
0 828 5 1 1 827
0 829 7 1 2 823 828
0 830 5 1 1 829
0 831 7 1 2 986 62
0 832 5 1 1 831
0 833 7 2 2 1262 1517
0 834 5 1 1 1555
0 835 7 1 2 1101 1155
0 836 5 2 1 835
0 837 7 1 2 1556 1557
0 838 7 1 2 832 837
0 839 5 1 1 838
0 840 7 1 2 1328 1522
0 841 5 1 1 840
0 842 7 1 2 1233 1520
0 843 5 1 1 842
0 844 7 2 2 841 843
0 845 5 1 1 1559
0 846 7 1 2 987 1151
0 847 7 1 2 845 846
0 848 5 1 1 847
0 849 7 1 2 839 848
0 850 5 1 1 849
0 851 7 1 2 830 850
0 852 5 1 1 851
0 853 7 2 2 1102 1158
0 854 5 1 1 1561
0 855 7 1 2 1560 854
0 856 5 1 1 855
0 857 7 1 2 1162 1558
0 858 5 1 1 857
0 859 7 1 2 834 1562
0 860 5 1 1 859
0 861 7 1 2 858 860
0 862 7 1 2 856 861
0 863 7 1 2 1554 862
0 864 5 1 1 863
0 865 7 1 2 852 864
0 866 5 1 1 865
0 867 7 1 2 1147 866
0 868 5 1 1 867
0 869 7 1 2 1329 1518
0 870 5 1 1 869
0 871 7 1 2 1263 1523
0 872 5 1 1 871
0 873 7 1 2 870 872
0 874 5 1 1 873
0 875 7 1 2 1326 874
0 876 5 1 1 875
0 877 7 1 2 868 876
0 878 7 1 2 821 877
0 879 5 1 1 878
0 880 7 1 2 1399 1534
0 881 7 1 2 879 880
0 882 5 1 1 881
0 883 7 2 2 1076 1123
0 884 7 1 2 1421 1563
0 885 5 1 1 884
0 886 7 1 2 1031 1343
0 887 5 2 1 886
0 888 7 1 2 929 1565
0 889 5 1 1 888
0 890 7 1 2 953 1354
0 891 7 1 2 889 890
0 892 5 1 1 891
0 893 7 1 2 885 892
0 894 5 1 1 893
0 895 7 1 2 1358 894
0 896 5 1 1 895
0 897 7 1 2 1077 1356
0 898 5 1 1 897
0 899 7 1 2 1509 898
0 900 5 1 1 899
0 901 7 1 2 1032 1422
0 902 5 1 1 901
0 903 7 1 2 930 1336
0 904 5 1 1 903
0 905 7 1 2 1566 904
0 906 5 1 1 905
0 907 7 1 2 902 906
0 908 5 1 1 907
0 909 7 1 2 900 908
0 910 5 1 1 909
0 911 7 1 2 954 1360
0 912 5 1 1 911
0 913 7 1 2 1337 1347
0 914 7 1 2 1564 913
0 915 5 1 1 914
0 916 7 1 2 912 915
0 917 5 1 1 916
0 918 7 1 2 1056 917
0 919 5 1 1 918
0 920 7 1 2 910 919
0 921 7 1 2 896 920
0 922 5 1 1 921
0 923 7 1 2 1525 922
0 924 7 1 2 1331 923
0 925 5 1 1 924
0 926 7 1 2 882 925
0 927 7 1 2 742 926
0 928 7 1 2 611 927
3 1999 5 0 1 928
