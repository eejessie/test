1 0 0 2 0
2 13 1 0
2 173 1 0
1 1 0 2 0
2 174 1 1
2 175 1 1
1 2 0 2 0
2 176 1 2
2 177 1 2
1 3 0 2 0
2 178 1 3
2 179 1 3
1 4 0 2 0
2 180 1 4
2 181 1 4
1 5 0 2 0
2 182 1 5
2 183 1 5
1 6 0 2 0
2 184 1 6
2 185 1 6
1 7 0 2 0
2 186 1 7
2 187 1 7
1 8 0 2 0
2 188 1 8
2 189 1 8
1 9 0 2 0
2 190 1 9
2 191 1 9
1 10 0 2 0
2 192 1 10
2 193 1 10
1 11 0 2 0
2 194 1 11
2 195 1 11
1 12 0 2 0
2 196 1 12
2 197 1 12
2 198 1 28
2 199 1 28
2 200 1 30
2 201 1 30
2 202 1 31
2 203 1 31
2 204 1 34
2 205 1 34
2 206 1 36
2 207 1 36
2 208 1 38
2 209 1 38
2 210 1 40
2 211 1 40
2 212 1 41
2 213 1 41
2 214 1 42
2 215 1 42
2 216 1 42
2 217 1 45
2 218 1 45
2 219 1 46
2 220 1 46
2 221 1 49
2 222 1 49
2 223 1 50
2 224 1 50
2 225 1 55
2 226 1 55
2 227 1 58
2 228 1 58
2 229 1 59
2 230 1 59
2 231 1 65
2 232 1 65
2 233 1 68
2 234 1 68
2 235 1 70
2 236 1 70
2 237 1 70
2 238 1 71
2 239 1 71
2 240 1 77
2 241 1 77
2 242 1 79
2 243 1 79
2 244 1 79
2 245 1 80
2 246 1 80
2 247 1 80
2 248 1 82
2 249 1 82
2 250 1 85
2 251 1 85
2 252 1 87
2 253 1 87
2 254 1 88
2 255 1 88
2 256 1 91
2 257 1 91
2 258 1 92
2 259 1 92
2 260 1 95
2 261 1 95
2 262 1 96
2 263 1 96
2 264 1 97
2 265 1 97
2 266 1 101
2 267 1 101
2 268 1 103
2 269 1 103
2 270 1 105
2 271 1 105
2 272 1 106
2 273 1 106
2 274 1 106
2 275 1 112
2 276 1 112
2 277 1 114
2 278 1 114
2 279 1 117
2 280 1 117
2 281 1 118
2 282 1 118
2 283 1 121
2 284 1 121
2 285 1 121
2 286 1 122
2 287 1 122
2 288 1 129
2 289 1 129
2 290 1 130
2 291 1 130
2 292 1 142
2 293 1 142
2 294 1 142
0 14 5 1 1 13
0 15 5 1 1 174
0 16 5 1 1 176
0 17 5 1 1 178
0 18 5 1 1 180
0 19 5 1 1 182
0 20 5 1 1 184
0 21 5 1 1 186
0 22 5 1 1 188
0 23 5 1 1 190
0 24 5 1 1 192
0 25 5 1 1 194
0 26 5 1 1 196
0 27 7 1 2 17 21
0 28 5 2 1 27
0 29 7 1 2 179 187
0 30 5 2 1 29
0 31 7 2 2 198 200
0 32 5 1 1 202
0 33 7 1 2 16 20
0 34 5 2 1 33
0 35 7 1 2 177 185
0 36 5 2 1 35
0 37 7 1 2 15 19
0 38 5 2 1 37
0 39 7 1 2 175 183
0 40 5 2 1 39
0 41 7 2 2 173 181
0 42 5 3 1 212
0 43 7 1 2 210 214
0 44 5 1 1 43
0 45 7 2 2 208 44
0 46 5 2 1 217
0 47 7 1 2 206 219
0 48 5 1 1 47
0 49 7 2 2 204 48
0 50 5 2 1 221
0 51 7 1 2 32 222
0 52 5 1 1 51
0 53 7 1 2 203 223
0 54 5 1 1 53
0 55 7 2 2 52 54
0 56 5 1 1 225
0 57 7 1 2 25 56
0 58 5 2 1 57
0 59 7 2 2 205 207
0 60 5 1 1 229
0 61 7 1 2 220 230
0 62 5 1 1 61
0 63 7 1 2 218 60
0 64 5 1 1 63
0 65 7 2 2 62 64
0 66 5 1 1 231
0 67 7 1 2 24 66
0 68 5 2 1 67
0 69 7 1 2 193 232
0 70 5 3 1 69
0 71 7 2 2 209 211
0 72 5 1 1 238
0 73 7 1 2 213 72
0 74 5 1 1 73
0 75 7 1 2 215 239
0 76 5 1 1 75
0 77 7 2 2 74 76
0 78 5 1 1 240
0 79 7 3 2 23 78
0 80 5 3 1 242
0 81 7 1 2 191 241
0 82 5 2 1 81
0 83 7 1 2 14 18
0 84 5 1 1 83
0 85 7 2 2 216 84
0 86 5 1 1 250
0 87 7 2 2 189 86
0 88 5 2 1 252
0 89 7 1 2 248 254
0 90 5 1 1 89
0 91 7 2 2 245 90
0 92 5 2 1 256
0 93 7 1 2 235 258
0 94 5 1 1 93
0 95 7 2 2 233 94
0 96 5 2 1 260
0 97 7 2 2 227 261
0 98 5 1 1 264
0 99 7 1 2 201 224
0 100 5 1 1 99
0 101 7 2 2 199 100
0 102 5 1 1 266
0 103 7 2 2 26 267
0 104 5 1 1 268
0 105 7 2 2 195 226
0 106 5 3 1 270
0 107 7 1 2 269 271
0 108 5 1 1 107
0 109 7 1 2 265 108
0 110 5 1 1 109
0 111 7 1 2 197 102
0 112 5 2 1 111
0 113 7 1 2 104 275
0 114 5 2 1 113
0 115 7 1 2 98 277
0 116 5 1 1 115
0 117 7 2 2 228 272
0 118 5 2 1 279
0 119 7 1 2 262 281
0 120 5 1 1 119
0 121 7 3 2 234 236
0 122 5 2 1 283
0 123 7 1 2 257 286
0 124 5 1 1 123
0 125 7 1 2 259 284
0 126 5 1 1 125
0 127 7 1 2 124 126
0 128 5 1 1 127
0 129 7 2 2 246 249
0 130 5 2 1 288
0 131 7 1 2 253 290
0 132 5 1 1 131
0 133 7 1 2 255 289
0 134 5 1 1 133
0 135 7 1 2 132 134
0 136 5 1 1 135
0 137 7 1 2 128 136
0 138 7 1 2 120 137
0 139 7 1 2 116 138
0 140 7 1 2 110 139
0 141 5 1 1 140
0 142 7 3 2 237 243
0 143 5 1 1 292
0 144 7 1 2 280 143
0 145 5 1 1 144
0 146 7 1 2 282 293
0 147 5 1 1 146
0 148 7 1 2 145 147
0 149 5 1 1 148
0 150 7 1 2 276 273
0 151 7 1 2 263 150
0 152 5 1 1 151
0 153 7 1 2 274 294
0 154 5 1 1 153
0 155 7 1 2 278 154
0 156 5 1 1 155
0 157 7 1 2 22 251
0 158 5 1 1 157
0 159 7 1 2 291 158
0 160 5 1 1 159
0 161 7 1 2 244 287
0 162 5 1 1 161
0 163 7 1 2 247 285
0 164 5 1 1 163
0 165 7 1 2 162 164
0 166 5 1 1 165
0 167 7 1 2 160 166
0 168 7 1 2 156 167
0 169 7 1 2 152 168
0 170 7 1 2 149 169
0 171 5 1 1 170
0 172 7 1 2 141 171
3 399 5 0 1 172
