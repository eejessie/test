1 0 0 4 0
2 49 1 0
2 4369 1 0
2 4370 1 0
2 4371 1 0
1 1 0 5 0
2 4372 1 1
2 4373 1 1
2 4374 1 1
2 4375 1 1
2 4376 1 1
1 2 0 6 0
2 4377 1 2
2 4378 1 2
2 4379 1 2
2 4380 1 2
2 4381 1 2
2 4382 1 2
1 3 0 6 0
2 4383 1 3
2 4384 1 3
2 4385 1 3
2 4386 1 3
2 4387 1 3
2 4388 1 3
1 4 0 6 0
2 4389 1 4
2 4390 1 4
2 4391 1 4
2 4392 1 4
2 4393 1 4
2 4394 1 4
1 5 0 7 0
2 4395 1 5
2 4396 1 5
2 4397 1 5
2 4398 1 5
2 4399 1 5
2 4400 1 5
2 4401 1 5
1 6 0 7 0
2 4402 1 6
2 4403 1 6
2 4404 1 6
2 4405 1 6
2 4406 1 6
2 4407 1 6
2 4408 1 6
1 7 0 6 0
2 4409 1 7
2 4410 1 7
2 4411 1 7
2 4412 1 7
2 4413 1 7
2 4414 1 7
1 8 0 7 0
2 4415 1 8
2 4416 1 8
2 4417 1 8
2 4418 1 8
2 4419 1 8
2 4420 1 8
2 4421 1 8
1 9 0 6 0
2 4422 1 9
2 4423 1 9
2 4424 1 9
2 4425 1 9
2 4426 1 9
2 4427 1 9
1 10 0 6 0
2 4428 1 10
2 4429 1 10
2 4430 1 10
2 4431 1 10
2 4432 1 10
2 4433 1 10
1 11 0 7 0
2 4434 1 11
2 4435 1 11
2 4436 1 11
2 4437 1 11
2 4438 1 11
2 4439 1 11
2 4440 1 11
1 12 0 7 0
2 4441 1 12
2 4442 1 12
2 4443 1 12
2 4444 1 12
2 4445 1 12
2 4446 1 12
2 4447 1 12
1 13 0 6 0
2 4448 1 13
2 4449 1 13
2 4450 1 13
2 4451 1 13
2 4452 1 13
2 4453 1 13
1 14 0 7 0
2 4454 1 14
2 4455 1 14
2 4456 1 14
2 4457 1 14
2 4458 1 14
2 4459 1 14
2 4460 1 14
1 15 0 6 0
2 4461 1 15
2 4462 1 15
2 4463 1 15
2 4464 1 15
2 4465 1 15
2 4466 1 15
1 16 0 6 0
2 4467 1 16
2 4468 1 16
2 4469 1 16
2 4470 1 16
2 4471 1 16
2 4472 1 16
1 17 0 7 0
2 4473 1 17
2 4474 1 17
2 4475 1 17
2 4476 1 17
2 4477 1 17
2 4478 1 17
2 4479 1 17
1 18 0 7 0
2 4480 1 18
2 4481 1 18
2 4482 1 18
2 4483 1 18
2 4484 1 18
2 4485 1 18
2 4486 1 18
1 19 0 6 0
2 4487 1 19
2 4488 1 19
2 4489 1 19
2 4490 1 19
2 4491 1 19
2 4492 1 19
1 20 0 7 0
2 4493 1 20
2 4494 1 20
2 4495 1 20
2 4496 1 20
2 4497 1 20
2 4498 1 20
2 4499 1 20
1 21 0 6 0
2 4500 1 21
2 4501 1 21
2 4502 1 21
2 4503 1 21
2 4504 1 21
2 4505 1 21
1 22 0 6 0
2 4506 1 22
2 4507 1 22
2 4508 1 22
2 4509 1 22
2 4510 1 22
2 4511 1 22
1 23 0 7 0
2 4512 1 23
2 4513 1 23
2 4514 1 23
2 4515 1 23
2 4516 1 23
2 4517 1 23
2 4518 1 23
1 24 0 7 0
2 4519 1 24
2 4520 1 24
2 4521 1 24
2 4522 1 24
2 4523 1 24
2 4524 1 24
2 4525 1 24
1 25 0 6 0
2 4526 1 25
2 4527 1 25
2 4528 1 25
2 4529 1 25
2 4530 1 25
2 4531 1 25
1 26 0 7 0
2 4532 1 26
2 4533 1 26
2 4534 1 26
2 4535 1 26
2 4536 1 26
2 4537 1 26
2 4538 1 26
1 27 0 6 0
2 4539 1 27
2 4540 1 27
2 4541 1 27
2 4542 1 27
2 4543 1 27
2 4544 1 27
1 28 0 6 0
2 4545 1 28
2 4546 1 28
2 4547 1 28
2 4548 1 28
2 4549 1 28
2 4550 1 28
1 29 0 7 0
2 4551 1 29
2 4552 1 29
2 4553 1 29
2 4554 1 29
2 4555 1 29
2 4556 1 29
2 4557 1 29
1 30 0 7 0
2 4558 1 30
2 4559 1 30
2 4560 1 30
2 4561 1 30
2 4562 1 30
2 4563 1 30
2 4564 1 30
1 31 0 6 0
2 4565 1 31
2 4566 1 31
2 4567 1 31
2 4568 1 31
2 4569 1 31
2 4570 1 31
1 32 0 7 0
2 4571 1 32
2 4572 1 32
2 4573 1 32
2 4574 1 32
2 4575 1 32
2 4576 1 32
2 4577 1 32
1 33 0 6 0
2 4578 1 33
2 4579 1 33
2 4580 1 33
2 4581 1 33
2 4582 1 33
2 4583 1 33
1 34 0 6 0
2 4584 1 34
2 4585 1 34
2 4586 1 34
2 4587 1 34
2 4588 1 34
2 4589 1 34
1 35 0 7 0
2 4590 1 35
2 4591 1 35
2 4592 1 35
2 4593 1 35
2 4594 1 35
2 4595 1 35
2 4596 1 35
1 36 0 7 0
2 4597 1 36
2 4598 1 36
2 4599 1 36
2 4600 1 36
2 4601 1 36
2 4602 1 36
2 4603 1 36
1 37 0 6 0
2 4604 1 37
2 4605 1 37
2 4606 1 37
2 4607 1 37
2 4608 1 37
2 4609 1 37
1 38 0 7 0
2 4610 1 38
2 4611 1 38
2 4612 1 38
2 4613 1 38
2 4614 1 38
2 4615 1 38
2 4616 1 38
1 39 0 6 0
2 4617 1 39
2 4618 1 39
2 4619 1 39
2 4620 1 39
2 4621 1 39
2 4622 1 39
1 40 0 6 0
2 4623 1 40
2 4624 1 40
2 4625 1 40
2 4626 1 40
2 4627 1 40
2 4628 1 40
1 41 0 7 0
2 4629 1 41
2 4630 1 41
2 4631 1 41
2 4632 1 41
2 4633 1 41
2 4634 1 41
2 4635 1 41
1 42 0 7 0
2 4636 1 42
2 4637 1 42
2 4638 1 42
2 4639 1 42
2 4640 1 42
2 4641 1 42
2 4642 1 42
1 43 0 7 0
2 4643 1 43
2 4644 1 43
2 4645 1 43
2 4646 1 43
2 4647 1 43
2 4648 1 43
2 4649 1 43
1 44 0 7 0
2 4650 1 44
2 4651 1 44
2 4652 1 44
2 4653 1 44
2 4654 1 44
2 4655 1 44
2 4656 1 44
1 45 0 8 0
2 4657 1 45
2 4658 1 45
2 4659 1 45
2 4660 1 45
2 4661 1 45
2 4662 1 45
2 4663 1 45
2 4664 1 45
1 46 0 8 0
2 4665 1 46
2 4666 1 46
2 4667 1 46
2 4668 1 46
2 4669 1 46
2 4670 1 46
2 4671 1 46
2 4672 1 46
1 47 0 7 0
2 4673 1 47
2 4674 1 47
2 4675 1 47
2 4676 1 47
2 4677 1 47
2 4678 1 47
2 4679 1 47
1 48 0 6 0
2 4680 1 48
2 4681 1 48
2 4682 1 48
2 4683 1 48
2 4684 1 48
2 4685 1 48
2 4686 1 50
2 4687 1 50
2 4688 1 50
2 4689 1 50
2 4690 1 50
2 4691 1 51
2 4692 1 51
2 4693 1 51
2 4694 1 51
2 4695 1 51
2 4696 1 51
2 4697 1 52
2 4698 1 52
2 4699 1 52
2 4700 1 52
2 4701 1 52
2 4702 1 52
2 4703 1 53
2 4704 1 53
2 4705 1 53
2 4706 1 53
2 4707 1 53
2 4708 1 53
2 4709 1 54
2 4710 1 54
2 4711 1 54
2 4712 1 54
2 4713 1 54
2 4714 1 54
2 4715 1 55
2 4716 1 55
2 4717 1 55
2 4718 1 55
2 4719 1 55
2 4720 1 56
2 4721 1 56
2 4722 1 56
2 4723 1 56
2 4724 1 56
2 4725 1 56
2 4726 1 57
2 4727 1 57
2 4728 1 57
2 4729 1 57
2 4730 1 57
2 4731 1 57
2 4732 1 58
2 4733 1 58
2 4734 1 58
2 4735 1 58
2 4736 1 58
2 4737 1 59
2 4738 1 59
2 4739 1 59
2 4740 1 59
2 4741 1 59
2 4742 1 59
2 4743 1 60
2 4744 1 60
2 4745 1 60
2 4746 1 60
2 4747 1 60
2 4748 1 60
2 4749 1 61
2 4750 1 61
2 4751 1 61
2 4752 1 61
2 4753 1 61
2 4754 1 62
2 4755 1 62
2 4756 1 62
2 4757 1 62
2 4758 1 62
2 4759 1 62
2 4760 1 63
2 4761 1 63
2 4762 1 63
2 4763 1 63
2 4764 1 63
2 4765 1 63
2 4766 1 64
2 4767 1 64
2 4768 1 64
2 4769 1 64
2 4770 1 64
2 4771 1 65
2 4772 1 65
2 4773 1 65
2 4774 1 65
2 4775 1 65
2 4776 1 65
2 4777 1 66
2 4778 1 66
2 4779 1 66
2 4780 1 66
2 4781 1 66
2 4782 1 66
2 4783 1 67
2 4784 1 67
2 4785 1 67
2 4786 1 67
2 4787 1 67
2 4788 1 68
2 4789 1 68
2 4790 1 68
2 4791 1 68
2 4792 1 68
2 4793 1 68
2 4794 1 69
2 4795 1 69
2 4796 1 69
2 4797 1 69
2 4798 1 69
2 4799 1 69
2 4800 1 69
2 4801 1 70
2 4802 1 70
2 4803 1 70
2 4804 1 70
2 4805 1 70
2 4806 1 70
2 4807 1 71
2 4808 1 71
2 4809 1 71
2 4810 1 71
2 4811 1 71
2 4812 1 71
2 4813 1 71
2 4814 1 72
2 4815 1 72
2 4816 1 72
2 4817 1 72
2 4818 1 72
2 4819 1 72
2 4820 1 72
2 4821 1 73
2 4822 1 73
2 4823 1 73
2 4824 1 73
2 4825 1 73
2 4826 1 73
2 4827 1 74
2 4828 1 74
2 4829 1 74
2 4830 1 74
2 4831 1 74
2 4832 1 74
2 4833 1 74
2 4834 1 75
2 4835 1 75
2 4836 1 75
2 4837 1 75
2 4838 1 75
2 4839 1 75
2 4840 1 75
2 4841 1 76
2 4842 1 76
2 4843 1 76
2 4844 1 76
2 4845 1 76
2 4846 1 76
2 4847 1 77
2 4848 1 77
2 4849 1 77
2 4850 1 77
2 4851 1 77
2 4852 1 77
2 4853 1 77
2 4854 1 78
2 4855 1 78
2 4856 1 78
2 4857 1 78
2 4858 1 78
2 4859 1 78
2 4860 1 78
2 4861 1 79
2 4862 1 79
2 4863 1 79
2 4864 1 79
2 4865 1 79
2 4866 1 79
2 4867 1 80
2 4868 1 80
2 4869 1 80
2 4870 1 80
2 4871 1 80
2 4872 1 80
2 4873 1 80
2 4874 1 81
2 4875 1 81
2 4876 1 81
2 4877 1 81
2 4878 1 81
2 4879 1 81
2 4880 1 81
2 4881 1 82
2 4882 1 82
2 4883 1 82
2 4884 1 82
2 4885 1 82
2 4886 1 83
2 4887 1 83
2 4888 1 83
2 4889 1 83
2 4890 1 83
2 4891 1 83
2 4892 1 84
2 4893 1 84
2 4894 1 84
2 4895 1 84
2 4896 1 84
2 4897 1 84
2 4898 1 85
2 4899 1 85
2 4900 1 85
2 4901 1 85
2 4902 1 85
2 4903 1 86
2 4904 1 86
2 4905 1 86
2 4906 1 86
2 4907 1 86
2 4908 1 86
2 4909 1 87
2 4910 1 87
2 4911 1 87
2 4912 1 87
2 4913 1 87
2 4914 1 87
2 4915 1 88
2 4916 1 88
2 4917 1 88
2 4918 1 88
2 4919 1 88
2 4920 1 89
2 4921 1 89
2 4922 1 89
2 4923 1 89
2 4924 1 89
2 4925 1 89
2 4926 1 90
2 4927 1 90
2 4928 1 90
2 4929 1 90
2 4930 1 90
2 4931 1 90
2 4932 1 91
2 4933 1 91
2 4934 1 91
2 4935 1 91
2 4936 1 91
2 4937 1 92
2 4938 1 92
2 4939 1 92
2 4940 1 92
2 4941 1 92
2 4942 1 92
2 4943 1 93
2 4944 1 93
2 4945 1 93
2 4946 1 93
2 4947 1 93
2 4948 1 94
2 4949 1 94
2 4950 1 94
2 4951 1 94
2 4952 1 94
2 4953 1 94
2 4954 1 95
2 4955 1 95
2 4956 1 95
2 4957 1 95
2 4958 1 95
2 4959 1 95
2 4960 1 96
2 4961 1 96
2 4962 1 96
2 4963 1 96
2 4964 1 96
2 4965 1 97
2 4966 1 97
2 4967 1 97
2 4968 1 98
2 4969 1 98
2 4970 1 98
2 4971 1 98
2 4972 1 103
2 4973 1 103
2 4974 1 104
2 4975 1 104
2 4976 1 105
2 4977 1 105
2 4978 1 109
2 4979 1 109
2 4980 1 111
2 4981 1 111
2 4982 1 112
2 4983 1 112
2 4984 1 115
2 4985 1 115
2 4986 1 116
2 4987 1 116
2 4988 1 120
2 4989 1 120
2 4990 1 123
2 4991 1 123
2 4992 1 126
2 4993 1 126
2 4994 1 128
2 4995 1 128
2 4996 1 129
2 4997 1 129
2 4998 1 132
2 4999 1 132
2 5000 1 133
2 5001 1 133
2 5002 1 134
2 5003 1 134
2 5004 1 138
2 5005 1 138
2 5006 1 141
2 5007 1 141
2 5008 1 142
2 5009 1 142
2 5010 1 145
2 5011 1 145
2 5012 1 148
2 5013 1 148
2 5014 1 150
2 5015 1 150
2 5016 1 151
2 5017 1 151
2 5018 1 156
2 5019 1 156
2 5020 1 159
2 5021 1 159
2 5022 1 164
2 5023 1 164
2 5024 1 164
2 5025 1 170
2 5026 1 170
2 5027 1 170
2 5028 1 172
2 5029 1 172
2 5030 1 175
2 5031 1 175
2 5032 1 178
2 5033 1 178
2 5034 1 180
2 5035 1 180
2 5036 1 181
2 5037 1 181
2 5038 1 186
2 5039 1 186
2 5040 1 189
2 5041 1 189
2 5042 1 190
2 5043 1 190
2 5044 1 193
2 5045 1 193
2 5046 1 196
2 5047 1 196
2 5048 1 198
2 5049 1 198
2 5050 1 199
2 5051 1 199
2 5052 1 204
2 5053 1 204
2 5054 1 207
2 5055 1 207
2 5056 1 212
2 5057 1 212
2 5058 1 212
2 5059 1 218
2 5060 1 218
2 5061 1 218
2 5062 1 220
2 5063 1 220
2 5064 1 223
2 5065 1 223
2 5066 1 226
2 5067 1 226
2 5068 1 228
2 5069 1 228
2 5070 1 229
2 5071 1 229
2 5072 1 234
2 5073 1 234
2 5074 1 237
2 5075 1 237
2 5076 1 238
2 5077 1 238
2 5078 1 241
2 5079 1 241
2 5080 1 244
2 5081 1 244
2 5082 1 246
2 5083 1 246
2 5084 1 247
2 5085 1 247
2 5086 1 252
2 5087 1 252
2 5088 1 255
2 5089 1 255
2 5090 1 260
2 5091 1 260
2 5092 1 260
2 5093 1 266
2 5094 1 266
2 5095 1 266
2 5096 1 268
2 5097 1 268
2 5098 1 271
2 5099 1 271
2 5100 1 274
2 5101 1 274
2 5102 1 276
2 5103 1 276
2 5104 1 277
2 5105 1 277
2 5106 1 282
2 5107 1 282
2 5108 1 285
2 5109 1 285
2 5110 1 286
2 5111 1 286
2 5112 1 289
2 5113 1 289
2 5114 1 292
2 5115 1 292
2 5116 1 294
2 5117 1 294
2 5118 1 295
2 5119 1 295
2 5120 1 300
2 5121 1 300
2 5122 1 303
2 5123 1 303
2 5124 1 308
2 5125 1 308
2 5126 1 308
2 5127 1 314
2 5128 1 314
2 5129 1 314
2 5130 1 316
2 5131 1 316
2 5132 1 319
2 5133 1 319
2 5134 1 322
2 5135 1 322
2 5136 1 324
2 5137 1 324
2 5138 1 325
2 5139 1 325
2 5140 1 330
2 5141 1 330
2 5142 1 333
2 5143 1 333
2 5144 1 334
2 5145 1 334
2 5146 1 337
2 5147 1 337
2 5148 1 340
2 5149 1 340
2 5150 1 342
2 5151 1 342
2 5152 1 343
2 5153 1 343
2 5154 1 348
2 5155 1 348
2 5156 1 351
2 5157 1 351
2 5158 1 356
2 5159 1 356
2 5160 1 356
2 5161 1 362
2 5162 1 362
2 5163 1 362
2 5164 1 364
2 5165 1 364
2 5166 1 367
2 5167 1 367
2 5168 1 370
2 5169 1 370
2 5170 1 372
2 5171 1 372
2 5172 1 373
2 5173 1 373
2 5174 1 378
2 5175 1 378
2 5176 1 381
2 5177 1 381
2 5178 1 382
2 5179 1 382
2 5180 1 385
2 5181 1 385
2 5182 1 388
2 5183 1 388
2 5184 1 390
2 5185 1 390
2 5186 1 391
2 5187 1 391
2 5188 1 396
2 5189 1 396
2 5190 1 399
2 5191 1 399
2 5192 1 404
2 5193 1 404
2 5194 1 404
2 5195 1 410
2 5196 1 410
2 5197 1 410
2 5198 1 412
2 5199 1 412
2 5200 1 415
2 5201 1 415
2 5202 1 418
2 5203 1 418
2 5204 1 420
2 5205 1 420
2 5206 1 421
2 5207 1 421
2 5208 1 426
2 5209 1 426
2 5210 1 429
2 5211 1 429
2 5212 1 430
2 5213 1 430
2 5214 1 433
2 5215 1 433
2 5216 1 436
2 5217 1 436
2 5218 1 438
2 5219 1 438
2 5220 1 439
2 5221 1 439
2 5222 1 444
2 5223 1 444
2 5224 1 447
2 5225 1 447
2 5226 1 452
2 5227 1 452
2 5228 1 452
2 5229 1 458
2 5230 1 458
2 5231 1 458
2 5232 1 460
2 5233 1 460
2 5234 1 463
2 5235 1 463
2 5236 1 466
2 5237 1 466
2 5238 1 468
2 5239 1 468
2 5240 1 469
2 5241 1 469
2 5242 1 474
2 5243 1 474
2 5244 1 477
2 5245 1 477
2 5246 1 478
2 5247 1 478
2 5248 1 481
2 5249 1 481
2 5250 1 484
2 5251 1 484
2 5252 1 486
2 5253 1 486
2 5254 1 487
2 5255 1 487
2 5256 1 492
2 5257 1 492
2 5258 1 495
2 5259 1 495
2 5260 1 500
2 5261 1 500
2 5262 1 500
2 5263 1 506
2 5264 1 506
2 5265 1 506
2 5266 1 508
2 5267 1 508
2 5268 1 511
2 5269 1 511
2 5270 1 514
2 5271 1 514
2 5272 1 516
2 5273 1 516
2 5274 1 517
2 5275 1 517
2 5276 1 522
2 5277 1 522
2 5278 1 525
2 5279 1 525
2 5280 1 526
2 5281 1 526
2 5282 1 529
2 5283 1 529
2 5284 1 532
2 5285 1 532
2 5286 1 534
2 5287 1 534
2 5288 1 535
2 5289 1 535
2 5290 1 540
2 5291 1 540
2 5292 1 543
2 5293 1 543
2 5294 1 548
2 5295 1 548
2 5296 1 548
2 5297 1 554
2 5298 1 554
2 5299 1 554
2 5300 1 556
2 5301 1 556
2 5302 1 559
2 5303 1 559
2 5304 1 562
2 5305 1 562
2 5306 1 564
2 5307 1 564
2 5308 1 565
2 5309 1 565
2 5310 1 570
2 5311 1 570
2 5312 1 573
2 5313 1 573
2 5314 1 574
2 5315 1 574
2 5316 1 577
2 5317 1 577
2 5318 1 580
2 5319 1 580
2 5320 1 582
2 5321 1 582
2 5322 1 583
2 5323 1 583
2 5324 1 588
2 5325 1 588
2 5326 1 591
2 5327 1 591
2 5328 1 596
2 5329 1 596
2 5330 1 596
2 5331 1 602
2 5332 1 602
2 5333 1 602
2 5334 1 604
2 5335 1 604
2 5336 1 607
2 5337 1 607
2 5338 1 610
2 5339 1 610
2 5340 1 612
2 5341 1 612
2 5342 1 613
2 5343 1 613
2 5344 1 618
2 5345 1 618
2 5346 1 621
2 5347 1 621
2 5348 1 622
2 5349 1 622
2 5350 1 625
2 5351 1 625
2 5352 1 628
2 5353 1 628
2 5354 1 630
2 5355 1 630
2 5356 1 631
2 5357 1 631
2 5358 1 636
2 5359 1 636
2 5360 1 639
2 5361 1 639
2 5362 1 644
2 5363 1 644
2 5364 1 644
2 5365 1 650
2 5366 1 650
2 5367 1 650
2 5368 1 652
2 5369 1 652
2 5370 1 655
2 5371 1 655
2 5372 1 658
2 5373 1 658
2 5374 1 660
2 5375 1 660
2 5376 1 661
2 5377 1 661
2 5378 1 666
2 5379 1 666
2 5380 1 669
2 5381 1 669
2 5382 1 670
2 5383 1 670
2 5384 1 673
2 5385 1 673
2 5386 1 676
2 5387 1 676
2 5388 1 678
2 5389 1 678
2 5390 1 679
2 5391 1 679
2 5392 1 684
2 5393 1 684
2 5394 1 687
2 5395 1 687
2 5396 1 692
2 5397 1 692
2 5398 1 692
2 5399 1 698
2 5400 1 698
2 5401 1 698
2 5402 1 700
2 5403 1 700
2 5404 1 703
2 5405 1 703
2 5406 1 706
2 5407 1 706
2 5408 1 708
2 5409 1 708
2 5410 1 709
2 5411 1 709
2 5412 1 714
2 5413 1 714
2 5414 1 717
2 5415 1 717
2 5416 1 718
2 5417 1 718
2 5418 1 721
2 5419 1 721
2 5420 1 724
2 5421 1 724
2 5422 1 726
2 5423 1 726
2 5424 1 727
2 5425 1 727
2 5426 1 732
2 5427 1 732
2 5428 1 735
2 5429 1 735
2 5430 1 740
2 5431 1 740
2 5432 1 740
2 5433 1 746
2 5434 1 746
2 5435 1 746
2 5436 1 748
2 5437 1 748
2 5438 1 751
2 5439 1 751
2 5440 1 754
2 5441 1 754
2 5442 1 756
2 5443 1 756
2 5444 1 757
2 5445 1 757
2 5446 1 762
2 5447 1 762
2 5448 1 765
2 5449 1 765
2 5450 1 766
2 5451 1 766
2 5452 1 769
2 5453 1 769
2 5454 1 772
2 5455 1 772
2 5456 1 774
2 5457 1 774
2 5458 1 775
2 5459 1 775
2 5460 1 780
2 5461 1 780
2 5462 1 783
2 5463 1 783
2 5464 1 788
2 5465 1 788
2 5466 1 788
2 5467 1 794
2 5468 1 794
2 5469 1 794
2 5470 1 796
2 5471 1 796
2 5472 1 799
2 5473 1 799
2 5474 1 802
2 5475 1 802
2 5476 1 804
2 5477 1 804
2 5478 1 805
2 5479 1 805
2 5480 1 810
2 5481 1 810
2 5482 1 813
2 5483 1 813
2 5484 1 814
2 5485 1 814
2 5486 1 817
2 5487 1 817
2 5488 1 820
2 5489 1 820
2 5490 1 822
2 5491 1 822
2 5492 1 823
2 5493 1 823
2 5494 1 828
2 5495 1 828
2 5496 1 831
2 5497 1 831
2 5498 1 836
2 5499 1 836
2 5500 1 836
2 5501 1 842
2 5502 1 842
2 5503 1 842
2 5504 1 844
2 5505 1 844
2 5506 1 847
2 5507 1 847
2 5508 1 850
2 5509 1 850
2 5510 1 852
2 5511 1 852
2 5512 1 853
2 5513 1 853
2 5514 1 858
2 5515 1 858
2 5516 1 861
2 5517 1 861
2 5518 1 862
2 5519 1 862
2 5520 1 865
2 5521 1 865
2 5522 1 868
2 5523 1 868
2 5524 1 870
2 5525 1 870
2 5526 1 871
2 5527 1 871
2 5528 1 876
2 5529 1 876
2 5530 1 879
2 5531 1 879
2 5532 1 884
2 5533 1 884
2 5534 1 884
2 5535 1 890
2 5536 1 890
2 5537 1 890
2 5538 1 892
2 5539 1 892
2 5540 1 895
2 5541 1 895
2 5542 1 898
2 5543 1 898
2 5544 1 900
2 5545 1 900
2 5546 1 901
2 5547 1 901
2 5548 1 906
2 5549 1 906
2 5550 1 909
2 5551 1 909
2 5552 1 910
2 5553 1 910
2 5554 1 913
2 5555 1 913
2 5556 1 916
2 5557 1 916
2 5558 1 918
2 5559 1 918
2 5560 1 919
2 5561 1 919
2 5562 1 924
2 5563 1 924
2 5564 1 927
2 5565 1 927
2 5566 1 932
2 5567 1 932
2 5568 1 932
2 5569 1 938
2 5570 1 938
2 5571 1 938
2 5572 1 940
2 5573 1 940
2 5574 1 943
2 5575 1 943
2 5576 1 946
2 5577 1 946
2 5578 1 948
2 5579 1 948
2 5580 1 949
2 5581 1 949
2 5582 1 954
2 5583 1 954
2 5584 1 957
2 5585 1 957
2 5586 1 958
2 5587 1 958
2 5588 1 961
2 5589 1 961
2 5590 1 964
2 5591 1 964
2 5592 1 966
2 5593 1 966
2 5594 1 967
2 5595 1 967
2 5596 1 972
2 5597 1 972
2 5598 1 975
2 5599 1 975
2 5600 1 980
2 5601 1 980
2 5602 1 980
2 5603 1 986
2 5604 1 986
2 5605 1 986
2 5606 1 988
2 5607 1 988
2 5608 1 991
2 5609 1 991
2 5610 1 994
2 5611 1 994
2 5612 1 996
2 5613 1 996
2 5614 1 997
2 5615 1 997
2 5616 1 1002
2 5617 1 1002
2 5618 1 1005
2 5619 1 1005
2 5620 1 1006
2 5621 1 1006
2 5622 1 1009
2 5623 1 1009
2 5624 1 1012
2 5625 1 1012
2 5626 1 1014
2 5627 1 1014
2 5628 1 1015
2 5629 1 1015
2 5630 1 1020
2 5631 1 1020
2 5632 1 1023
2 5633 1 1023
2 5634 1 1028
2 5635 1 1028
2 5636 1 1028
2 5637 1 1034
2 5638 1 1034
2 5639 1 1034
2 5640 1 1036
2 5641 1 1036
2 5642 1 1039
2 5643 1 1039
2 5644 1 1042
2 5645 1 1042
2 5646 1 1044
2 5647 1 1044
2 5648 1 1045
2 5649 1 1045
2 5650 1 1050
2 5651 1 1050
2 5652 1 1053
2 5653 1 1053
2 5654 1 1054
2 5655 1 1054
2 5656 1 1057
2 5657 1 1057
2 5658 1 1060
2 5659 1 1060
2 5660 1 1062
2 5661 1 1062
2 5662 1 1063
2 5663 1 1063
2 5664 1 1068
2 5665 1 1068
2 5666 1 1071
2 5667 1 1071
2 5668 1 1076
2 5669 1 1076
2 5670 1 1076
2 5671 1 1082
2 5672 1 1082
2 5673 1 1082
2 5674 1 1084
2 5675 1 1084
2 5676 1 1087
2 5677 1 1087
2 5678 1 1090
2 5679 1 1090
2 5680 1 1092
2 5681 1 1092
2 5682 1 1093
2 5683 1 1093
2 5684 1 1098
2 5685 1 1098
2 5686 1 1101
2 5687 1 1101
2 5688 1 1102
2 5689 1 1102
2 5690 1 1105
2 5691 1 1105
2 5692 1 1108
2 5693 1 1108
2 5694 1 1110
2 5695 1 1110
2 5696 1 1111
2 5697 1 1111
2 5698 1 1116
2 5699 1 1116
2 5700 1 1119
2 5701 1 1119
2 5702 1 1124
2 5703 1 1124
2 5704 1 1124
2 5705 1 1126
2 5706 1 1126
2 5707 1 1129
2 5708 1 1129
2 5709 1 1132
2 5710 1 1132
2 5711 1 1132
2 5712 1 1133
2 5713 1 1133
2 5714 1 1135
2 5715 1 1135
2 5716 1 1140
2 5717 1 1140
2 5718 1 1143
2 5719 1 1143
2 5720 1 1148
2 5721 1 1148
2 5722 1 1154
2 5723 1 1154
2 5724 1 1156
2 5725 1 1156
2 5726 1 1159
2 5727 1 1159
2 5728 1 1160
2 5729 1 1160
2 5730 1 1163
2 5731 1 1163
2 5732 1 1163
2 5733 1 1170
2 5734 1 1170
2 5735 1 1189
2 5736 1 1189
2 5737 1 1193
2 5738 1 1193
2 5739 1 1196
2 5740 1 1196
2 5741 1 1199
2 5742 1 1199
2 5743 1 1204
2 5744 1 1204
2 5745 1 1205
2 5746 1 1205
2 5747 1 1212
2 5748 1 1212
2 5749 1 1215
2 5750 1 1215
2 5751 1 1218
2 5752 1 1218
2 5753 1 1219
2 5754 1 1219
2 5755 1 1219
2 5756 1 1227
2 5757 1 1227
2 5758 1 1231
2 5759 1 1231
2 5760 1 1234
2 5761 1 1234
2 5762 1 1240
2 5763 1 1240
2 5764 1 1243
2 5765 1 1243
2 5766 1 1246
2 5767 1 1246
2 5768 1 1247
2 5769 1 1247
2 5770 1 1247
2 5771 1 1253
2 5772 1 1253
2 5773 1 1257
2 5774 1 1257
2 5775 1 1260
2 5776 1 1260
2 5777 1 1261
2 5778 1 1261
2 5779 1 1267
2 5780 1 1267
2 5781 1 1270
2 5782 1 1270
2 5783 1 1276
2 5784 1 1276
2 5785 1 1280
2 5786 1 1280
2 5787 1 1282
2 5788 1 1282
2 5789 1 1285
2 5790 1 1285
2 5791 1 1288
2 5792 1 1288
2 5793 1 1295
2 5794 1 1295
2 5795 1 1299
2 5796 1 1299
2 5797 1 1300
2 5798 1 1300
2 5799 1 1301
2 5800 1 1301
2 5801 1 1302
2 5802 1 1302
2 5803 1 1309
2 5804 1 1309
2 5805 1 1312
2 5806 1 1312
2 5807 1 1318
2 5808 1 1318
2 5809 1 1324
2 5810 1 1324
2 5811 1 1327
2 5812 1 1327
2 5813 1 1330
2 5814 1 1330
2 5815 1 1331
2 5816 1 1331
2 5817 1 1331
2 5818 1 1337
2 5819 1 1337
2 5820 1 1341
2 5821 1 1341
2 5822 1 1344
2 5823 1 1344
2 5824 1 1345
2 5825 1 1345
2 5826 1 1351
2 5827 1 1351
2 5828 1 1354
2 5829 1 1354
2 5830 1 1360
2 5831 1 1360
2 5832 1 1364
2 5833 1 1364
2 5834 1 1366
2 5835 1 1366
2 5836 1 1369
2 5837 1 1369
2 5838 1 1372
2 5839 1 1372
2 5840 1 1379
2 5841 1 1379
2 5842 1 1383
2 5843 1 1383
2 5844 1 1384
2 5845 1 1384
2 5846 1 1385
2 5847 1 1385
2 5848 1 1386
2 5849 1 1386
2 5850 1 1393
2 5851 1 1393
2 5852 1 1396
2 5853 1 1396
2 5854 1 1402
2 5855 1 1402
2 5856 1 1408
2 5857 1 1408
2 5858 1 1411
2 5859 1 1411
2 5860 1 1414
2 5861 1 1414
2 5862 1 1415
2 5863 1 1415
2 5864 1 1415
2 5865 1 1421
2 5866 1 1421
2 5867 1 1425
2 5868 1 1425
2 5869 1 1428
2 5870 1 1428
2 5871 1 1429
2 5872 1 1429
2 5873 1 1435
2 5874 1 1435
2 5875 1 1438
2 5876 1 1438
2 5877 1 1444
2 5878 1 1444
2 5879 1 1448
2 5880 1 1448
2 5881 1 1450
2 5882 1 1450
2 5883 1 1453
2 5884 1 1453
2 5885 1 1456
2 5886 1 1456
2 5887 1 1463
2 5888 1 1463
2 5889 1 1467
2 5890 1 1467
2 5891 1 1468
2 5892 1 1468
2 5893 1 1469
2 5894 1 1469
2 5895 1 1470
2 5896 1 1470
2 5897 1 1477
2 5898 1 1477
2 5899 1 1480
2 5900 1 1480
2 5901 1 1486
2 5902 1 1486
2 5903 1 1492
2 5904 1 1492
2 5905 1 1495
2 5906 1 1495
2 5907 1 1498
2 5908 1 1498
2 5909 1 1499
2 5910 1 1499
2 5911 1 1499
2 5912 1 1505
2 5913 1 1505
2 5914 1 1509
2 5915 1 1509
2 5916 1 1512
2 5917 1 1512
2 5918 1 1513
2 5919 1 1513
2 5920 1 1519
2 5921 1 1519
2 5922 1 1522
2 5923 1 1522
2 5924 1 1528
2 5925 1 1528
2 5926 1 1532
2 5927 1 1532
2 5928 1 1534
2 5929 1 1534
2 5930 1 1537
2 5931 1 1537
2 5932 1 1540
2 5933 1 1540
2 5934 1 1547
2 5935 1 1547
2 5936 1 1551
2 5937 1 1551
2 5938 1 1552
2 5939 1 1552
2 5940 1 1553
2 5941 1 1553
2 5942 1 1554
2 5943 1 1554
2 5944 1 1561
2 5945 1 1561
2 5946 1 1564
2 5947 1 1564
2 5948 1 1570
2 5949 1 1570
2 5950 1 1576
2 5951 1 1576
2 5952 1 1579
2 5953 1 1579
2 5954 1 1582
2 5955 1 1582
2 5956 1 1583
2 5957 1 1583
2 5958 1 1583
2 5959 1 1589
2 5960 1 1589
2 5961 1 1593
2 5962 1 1593
2 5963 1 1596
2 5964 1 1596
2 5965 1 1597
2 5966 1 1597
2 5967 1 1603
2 5968 1 1603
2 5969 1 1606
2 5970 1 1606
2 5971 1 1612
2 5972 1 1612
2 5973 1 1616
2 5974 1 1616
2 5975 1 1618
2 5976 1 1618
2 5977 1 1621
2 5978 1 1621
2 5979 1 1624
2 5980 1 1624
2 5981 1 1631
2 5982 1 1631
2 5983 1 1635
2 5984 1 1635
2 5985 1 1636
2 5986 1 1636
2 5987 1 1637
2 5988 1 1637
2 5989 1 1638
2 5990 1 1638
2 5991 1 1645
2 5992 1 1645
2 5993 1 1648
2 5994 1 1648
2 5995 1 1654
2 5996 1 1654
2 5997 1 1660
2 5998 1 1660
2 5999 1 1663
2 6000 1 1663
2 6001 1 1666
2 6002 1 1666
2 6003 1 1667
2 6004 1 1667
2 6005 1 1667
2 6006 1 1673
2 6007 1 1673
2 6008 1 1677
2 6009 1 1677
2 6010 1 1680
2 6011 1 1680
2 6012 1 1681
2 6013 1 1681
2 6014 1 1687
2 6015 1 1687
2 6016 1 1690
2 6017 1 1690
2 6018 1 1696
2 6019 1 1696
2 6020 1 1700
2 6021 1 1700
2 6022 1 1702
2 6023 1 1702
2 6024 1 1705
2 6025 1 1705
2 6026 1 1708
2 6027 1 1708
2 6028 1 1715
2 6029 1 1715
2 6030 1 1719
2 6031 1 1719
2 6032 1 1720
2 6033 1 1720
2 6034 1 1721
2 6035 1 1721
2 6036 1 1722
2 6037 1 1722
2 6038 1 1729
2 6039 1 1729
2 6040 1 1732
2 6041 1 1732
2 6042 1 1738
2 6043 1 1738
2 6044 1 1744
2 6045 1 1744
2 6046 1 1747
2 6047 1 1747
2 6048 1 1750
2 6049 1 1750
2 6050 1 1751
2 6051 1 1751
2 6052 1 1751
2 6053 1 1759
2 6054 1 1759
2 6055 1 1763
2 6056 1 1763
2 6057 1 1767
2 6058 1 1767
2 6059 1 1772
2 6060 1 1772
2 6061 1 1773
2 6062 1 1773
2 6063 1 1776
2 6064 1 1776
2 6065 1 1778
2 6066 1 1778
2 6067 1 1779
2 6068 1 1779
2 6069 1 1784
2 6070 1 1784
2 6071 1 1787
2 6072 1 1787
2 6073 1 1793
2 6074 1 1793
2 6075 1 1798
2 6076 1 1798
2 6077 1 1799
2 6078 1 1799
2 6079 1 1802
2 6080 1 1802
2 6081 1 1804
2 6082 1 1804
2 6083 1 1820
2 6084 1 1820
2 6085 1 1823
2 6086 1 1823
2 6087 1 1829
2 6088 1 1829
2 6089 1 1829
2 6090 1 1830
2 6091 1 1830
2 6092 1 1830
2 6093 1 1830
2 6094 1 1830
2 6095 1 1832
2 6096 1 1832
2 6097 1 1833
2 6098 1 1833
2 6099 1 1834
2 6100 1 1834
2 6101 1 1841
2 6102 1 1841
2 6103 1 1842
2 6104 1 1842
2 6105 1 1849
2 6106 1 1849
2 6107 1 1849
2 6108 1 1855
2 6109 1 1855
2 6110 1 1856
2 6111 1 1856
2 6112 1 1857
2 6113 1 1857
2 6114 1 1859
2 6115 1 1859
2 6116 1 1861
2 6117 1 1861
2 6118 1 1862
2 6119 1 1862
2 6120 1 1873
2 6121 1 1873
2 6122 1 1875
2 6123 1 1875
2 6124 1 1877
2 6125 1 1877
2 6126 1 1880
2 6127 1 1880
2 6128 1 1880
2 6129 1 1880
2 6130 1 1885
2 6131 1 1885
2 6132 1 1886
2 6133 1 1886
2 6134 1 1890
2 6135 1 1890
2 6136 1 1899
2 6137 1 1899
2 6138 1 1902
2 6139 1 1902
2 6140 1 1903
2 6141 1 1903
2 6142 1 1906
2 6143 1 1906
2 6144 1 1906
2 6145 1 1908
2 6146 1 1908
2 6147 1 1910
2 6148 1 1910
2 6149 1 1912
2 6150 1 1912
2 6151 1 1919
2 6152 1 1919
2 6153 1 1920
2 6154 1 1920
2 6155 1 1926
2 6156 1 1926
2 6157 1 1929
2 6158 1 1929
2 6159 1 1930
2 6160 1 1930
2 6161 1 1935
2 6162 1 1935
2 6163 1 1939
2 6164 1 1939
2 6165 1 1939
2 6166 1 1939
2 6167 1 1943
2 6168 1 1943
2 6169 1 1946
2 6170 1 1946
2 6171 1 1947
2 6172 1 1947
2 6173 1 1950
2 6174 1 1950
2 6175 1 1950
2 6176 1 1953
2 6177 1 1953
2 6178 1 1957
2 6179 1 1957
2 6180 1 1958
2 6181 1 1958
2 6182 1 1960
2 6183 1 1960
2 6184 1 1962
2 6185 1 1962
2 6186 1 1964
2 6187 1 1964
2 6188 1 1967
2 6189 1 1967
2 6190 1 1967
2 6191 1 1967
2 6192 1 1969
2 6193 1 1969
2 6194 1 1971
2 6195 1 1971
2 6196 1 1975
2 6197 1 1975
2 6198 1 1984
2 6199 1 1984
2 6200 1 1985
2 6201 1 1985
2 6202 1 1991
2 6203 1 1991
2 6204 1 1994
2 6205 1 1994
2 6206 1 1995
2 6207 1 1995
2 6208 1 1998
2 6209 1 1998
2 6210 1 2000
2 6211 1 2000
2 6212 1 2002
2 6213 1 2002
2 6214 1 2004
2 6215 1 2004
2 6216 1 2006
2 6217 1 2006
2 6218 1 2009
2 6219 1 2009
2 6220 1 2009
2 6221 1 2009
2 6222 1 2014
2 6223 1 2014
2 6224 1 2015
2 6225 1 2015
2 6226 1 2019
2 6227 1 2019
2 6228 1 2028
2 6229 1 2028
2 6230 1 2031
2 6231 1 2031
2 6232 1 2032
2 6233 1 2032
2 6234 1 2035
2 6235 1 2035
2 6236 1 2035
2 6237 1 2037
2 6238 1 2037
2 6239 1 2039
2 6240 1 2039
2 6241 1 2041
2 6242 1 2041
2 6243 1 2048
2 6244 1 2048
2 6245 1 2049
2 6246 1 2049
2 6247 1 2055
2 6248 1 2055
2 6249 1 2058
2 6250 1 2058
2 6251 1 2059
2 6252 1 2059
2 6253 1 2064
2 6254 1 2064
2 6255 1 2068
2 6256 1 2068
2 6257 1 2068
2 6258 1 2068
2 6259 1 2072
2 6260 1 2072
2 6261 1 2075
2 6262 1 2075
2 6263 1 2076
2 6264 1 2076
2 6265 1 2079
2 6266 1 2079
2 6267 1 2079
2 6268 1 2082
2 6269 1 2082
2 6270 1 2086
2 6271 1 2086
2 6272 1 2087
2 6273 1 2087
2 6274 1 2089
2 6275 1 2089
2 6276 1 2091
2 6277 1 2091
2 6278 1 2093
2 6279 1 2093
2 6280 1 2096
2 6281 1 2096
2 6282 1 2096
2 6283 1 2096
2 6284 1 2098
2 6285 1 2098
2 6286 1 2100
2 6287 1 2100
2 6288 1 2104
2 6289 1 2104
2 6290 1 2113
2 6291 1 2113
2 6292 1 2114
2 6293 1 2114
2 6294 1 2120
2 6295 1 2120
2 6296 1 2123
2 6297 1 2123
2 6298 1 2124
2 6299 1 2124
2 6300 1 2127
2 6301 1 2127
2 6302 1 2127
2 6303 1 2127
2 6304 1 2131
2 6305 1 2131
2 6306 1 2134
2 6307 1 2134
2 6308 1 2135
2 6309 1 2135
2 6310 1 2138
2 6311 1 2138
2 6312 1 2138
2 6313 1 2138
2 6314 1 2142
2 6315 1 2142
2 6316 1 2144
2 6317 1 2144
2 6318 1 2153
2 6319 1 2153
2 6320 1 2156
2 6321 1 2156
2 6322 1 2157
2 6323 1 2157
2 6324 1 2160
2 6325 1 2160
2 6326 1 2160
2 6327 1 2160
2 6328 1 2162
2 6329 1 2162
2 6330 1 2164
2 6331 1 2164
2 6332 1 2168
2 6333 1 2168
2 6334 1 2177
2 6335 1 2177
2 6336 1 2178
2 6337 1 2178
2 6338 1 2184
2 6339 1 2184
2 6340 1 2187
2 6341 1 2187
2 6342 1 2188
2 6343 1 2188
2 6344 1 2191
2 6345 1 2191
2 6346 1 2191
2 6347 1 2193
2 6348 1 2193
2 6349 1 2195
2 6350 1 2195
2 6351 1 2197
2 6352 1 2197
2 6353 1 2199
2 6354 1 2199
2 6355 1 2202
2 6356 1 2202
2 6357 1 2202
2 6358 1 2202
2 6359 1 2206
2 6360 1 2206
2 6361 1 2208
2 6362 1 2208
2 6363 1 2217
2 6364 1 2217
2 6365 1 2220
2 6366 1 2220
2 6367 1 2221
2 6368 1 2221
2 6369 1 2224
2 6370 1 2224
2 6371 1 2224
2 6372 1 2224
2 6373 1 2226
2 6374 1 2226
2 6375 1 2228
2 6376 1 2228
2 6377 1 2232
2 6378 1 2232
2 6379 1 2241
2 6380 1 2241
2 6381 1 2242
2 6382 1 2242
2 6383 1 2248
2 6384 1 2248
2 6385 1 2251
2 6386 1 2251
2 6387 1 2252
2 6388 1 2252
2 6389 1 2255
2 6390 1 2255
2 6391 1 2255
2 6392 1 2255
2 6393 1 2259
2 6394 1 2259
2 6395 1 2262
2 6396 1 2262
2 6397 1 2263
2 6398 1 2263
2 6399 1 2266
2 6400 1 2266
2 6401 1 2266
2 6402 1 2266
2 6403 1 2270
2 6404 1 2270
2 6405 1 2272
2 6406 1 2272
2 6407 1 2281
2 6408 1 2281
2 6409 1 2284
2 6410 1 2284
2 6411 1 2285
2 6412 1 2285
2 6413 1 2288
2 6414 1 2288
2 6415 1 2288
2 6416 1 2288
2 6417 1 2290
2 6418 1 2290
2 6419 1 2292
2 6420 1 2292
2 6421 1 2296
2 6422 1 2296
2 6423 1 2305
2 6424 1 2305
2 6425 1 2306
2 6426 1 2306
2 6427 1 2312
2 6428 1 2312
2 6429 1 2315
2 6430 1 2315
2 6431 1 2316
2 6432 1 2316
2 6433 1 2319
2 6434 1 2319
2 6435 1 2319
2 6436 1 2319
2 6437 1 2323
2 6438 1 2323
2 6439 1 2326
2 6440 1 2326
2 6441 1 2327
2 6442 1 2327
2 6443 1 2330
2 6444 1 2330
2 6445 1 2330
2 6446 1 2332
2 6447 1 2332
2 6448 1 2334
2 6449 1 2334
2 6450 1 2336
2 6451 1 2336
2 6452 1 2345
2 6453 1 2345
2 6454 1 2347
2 6455 1 2347
2 6456 1 2349
2 6457 1 2349
2 6458 1 2352
2 6459 1 2352
2 6460 1 2352
2 6461 1 2352
2 6462 1 2354
2 6463 1 2354
2 6464 1 2356
2 6465 1 2356
2 6466 1 2360
2 6467 1 2360
2 6468 1 2369
2 6469 1 2369
2 6470 1 2370
2 6471 1 2370
2 6472 1 2376
2 6473 1 2376
2 6474 1 2379
2 6475 1 2379
2 6476 1 2380
2 6477 1 2380
2 6478 1 2383
2 6479 1 2383
2 6480 1 2383
2 6481 1 2383
2 6482 1 2387
2 6483 1 2387
2 6484 1 2390
2 6485 1 2390
2 6486 1 2391
2 6487 1 2391
2 6488 1 2394
2 6489 1 2394
2 6490 1 2394
2 6491 1 2394
2 6492 1 2398
2 6493 1 2398
2 6494 1 2400
2 6495 1 2400
2 6496 1 2409
2 6497 1 2409
2 6498 1 2412
2 6499 1 2412
2 6500 1 2413
2 6501 1 2413
2 6502 1 2416
2 6503 1 2416
2 6504 1 2416
2 6505 1 2416
2 6506 1 2418
2 6507 1 2418
2 6508 1 2420
2 6509 1 2420
2 6510 1 2424
2 6511 1 2424
2 6512 1 2433
2 6513 1 2433
2 6514 1 2434
2 6515 1 2434
2 6516 1 2440
2 6517 1 2440
2 6518 1 2443
2 6519 1 2443
2 6520 1 2444
2 6521 1 2444
2 6522 1 2447
2 6523 1 2447
2 6524 1 2447
2 6525 1 2447
2 6526 1 2451
2 6527 1 2451
2 6528 1 2454
2 6529 1 2454
2 6530 1 2455
2 6531 1 2455
2 6532 1 2458
2 6533 1 2458
2 6534 1 2458
2 6535 1 2460
2 6536 1 2460
2 6537 1 2462
2 6538 1 2462
2 6539 1 2464
2 6540 1 2464
2 6541 1 2473
2 6542 1 2473
2 6543 1 2475
2 6544 1 2475
2 6545 1 2477
2 6546 1 2477
2 6547 1 2480
2 6548 1 2480
2 6549 1 2480
2 6550 1 2480
2 6551 1 2482
2 6552 1 2482
2 6553 1 2484
2 6554 1 2484
2 6555 1 2488
2 6556 1 2488
2 6557 1 2497
2 6558 1 2497
2 6559 1 2498
2 6560 1 2498
2 6561 1 2504
2 6562 1 2504
2 6563 1 2507
2 6564 1 2507
2 6565 1 2508
2 6566 1 2508
2 6567 1 2511
2 6568 1 2511
2 6569 1 2511
2 6570 1 2511
2 6571 1 2515
2 6572 1 2515
2 6573 1 2518
2 6574 1 2518
2 6575 1 2519
2 6576 1 2519
2 6577 1 2522
2 6578 1 2522
2 6579 1 2522
2 6580 1 2522
2 6581 1 2526
2 6582 1 2526
2 6583 1 2528
2 6584 1 2528
2 6585 1 2537
2 6586 1 2537
2 6587 1 2540
2 6588 1 2540
2 6589 1 2541
2 6590 1 2541
2 6591 1 2544
2 6592 1 2544
2 6593 1 2544
2 6594 1 2544
2 6595 1 2546
2 6596 1 2546
2 6597 1 2548
2 6598 1 2548
2 6599 1 2552
2 6600 1 2552
2 6601 1 2561
2 6602 1 2561
2 6603 1 2562
2 6604 1 2562
2 6605 1 2568
2 6606 1 2568
2 6607 1 2571
2 6608 1 2571
2 6609 1 2572
2 6610 1 2572
2 6611 1 2575
2 6612 1 2575
2 6613 1 2575
2 6614 1 2575
2 6615 1 2579
2 6616 1 2579
2 6617 1 2582
2 6618 1 2582
2 6619 1 2583
2 6620 1 2583
2 6621 1 2586
2 6622 1 2586
2 6623 1 2586
2 6624 1 2588
2 6625 1 2588
2 6626 1 2590
2 6627 1 2590
2 6628 1 2592
2 6629 1 2592
2 6630 1 2601
2 6631 1 2601
2 6632 1 2603
2 6633 1 2603
2 6634 1 2605
2 6635 1 2605
2 6636 1 2608
2 6637 1 2608
2 6638 1 2608
2 6639 1 2608
2 6640 1 2610
2 6641 1 2610
2 6642 1 2612
2 6643 1 2612
2 6644 1 2616
2 6645 1 2616
2 6646 1 2625
2 6647 1 2625
2 6648 1 2626
2 6649 1 2626
2 6650 1 2632
2 6651 1 2632
2 6652 1 2635
2 6653 1 2635
2 6654 1 2636
2 6655 1 2636
2 6656 1 2639
2 6657 1 2639
2 6658 1 2639
2 6659 1 2639
2 6660 1 2643
2 6661 1 2643
2 6662 1 2646
2 6663 1 2646
2 6664 1 2647
2 6665 1 2647
2 6666 1 2650
2 6667 1 2650
2 6668 1 2650
2 6669 1 2650
2 6670 1 2654
2 6671 1 2654
2 6672 1 2656
2 6673 1 2656
2 6674 1 2665
2 6675 1 2665
2 6676 1 2668
2 6677 1 2668
2 6678 1 2669
2 6679 1 2669
2 6680 1 2672
2 6681 1 2672
2 6682 1 2672
2 6683 1 2672
2 6684 1 2674
2 6685 1 2674
2 6686 1 2676
2 6687 1 2676
2 6688 1 2678
2 6689 1 2678
2 6690 1 2685
2 6691 1 2685
2 6692 1 2686
2 6693 1 2686
2 6694 1 2689
2 6695 1 2689
2 6696 1 2690
2 6697 1 2690
2 6698 1 2693
2 6699 1 2693
2 6700 1 2693
2 6701 1 2693
2 6702 1 2704
2 6703 1 2704
2 6704 1 2707
2 6705 1 2707
2 6706 1 2710
2 6707 1 2710
2 6708 1 2711
2 6709 1 2711
2 6710 1 2714
2 6711 1 2714
2 6712 1 2714
2 6713 1 2716
2 6714 1 2716
2 6715 1 2718
2 6716 1 2718
2 6717 1 2720
2 6718 1 2720
2 6719 1 2733
2 6720 1 2733
2 6721 1 2735
2 6722 1 2735
2 6723 1 2737
2 6724 1 2737
2 6725 1 2740
2 6726 1 2740
2 6727 1 2741
2 6728 1 2741
2 6729 1 2743
2 6730 1 2743
2 6731 1 2746
2 6732 1 2746
2 6733 1 2746
2 6734 1 2746
2 6735 1 2748
2 6736 1 2748
2 6737 1 2750
2 6738 1 2750
2 6739 1 2753
2 6740 1 2753
2 6741 1 2754
2 6742 1 2754
2 6743 1 2757
2 6744 1 2757
2 6745 1 2757
2 6746 1 2768
2 6747 1 2768
2 6748 1 2771
2 6749 1 2771
2 6750 1 2774
2 6751 1 2774
2 6752 1 2775
2 6753 1 2775
2 6754 1 2779
2 6755 1 2779
2 6756 1 2780
2 6757 1 2780
2 6758 1 2797
2 6759 1 2797
2 6760 1 2808
2 6761 1 2808
2 6762 1 2811
2 6763 1 2811
2 6764 1 2813
2 6765 1 2813
2 6766 1 2815
2 6767 1 2815
2 6768 1 2817
2 6769 1 2817
2 6770 1 2818
2 6771 1 2818
2 6772 1 2819
2 6773 1 2819
2 6774 1 2819
2 6775 1 2822
2 6776 1 2822
2 6777 1 2823
2 6778 1 2823
2 6779 1 2826
2 6780 1 2826
2 6781 1 2829
2 6782 1 2829
2 6783 1 2831
2 6784 1 2831
2 6785 1 2834
2 6786 1 2834
2 6787 1 2837
2 6788 1 2837
2 6789 1 2839
2 6790 1 2839
2 6791 1 2842
2 6792 1 2842
2 6793 1 2845
2 6794 1 2845
2 6795 1 2847
2 6796 1 2847
2 6797 1 2850
2 6798 1 2850
2 6799 1 2853
2 6800 1 2853
2 6801 1 2855
2 6802 1 2855
2 6803 1 2858
2 6804 1 2858
2 6805 1 2861
2 6806 1 2861
2 6807 1 2863
2 6808 1 2863
2 6809 1 2866
2 6810 1 2866
2 6811 1 2869
2 6812 1 2869
2 6813 1 2871
2 6814 1 2871
2 6815 1 2874
2 6816 1 2874
2 6817 1 2877
2 6818 1 2877
2 6819 1 2879
2 6820 1 2879
2 6821 1 2882
2 6822 1 2882
2 6823 1 2885
2 6824 1 2885
2 6825 1 2887
2 6826 1 2887
2 6827 1 2890
2 6828 1 2890
2 6829 1 2893
2 6830 1 2893
2 6831 1 2895
2 6832 1 2895
2 6833 1 2898
2 6834 1 2898
2 6835 1 2901
2 6836 1 2901
2 6837 1 2903
2 6838 1 2903
2 6839 1 2906
2 6840 1 2906
2 6841 1 2909
2 6842 1 2909
2 6843 1 2911
2 6844 1 2911
2 6845 1 2914
2 6846 1 2914
2 6847 1 2917
2 6848 1 2917
2 6849 1 2919
2 6850 1 2919
2 6851 1 2922
2 6852 1 2922
2 6853 1 2925
2 6854 1 2925
2 6855 1 2927
2 6856 1 2927
2 6857 1 2930
2 6858 1 2930
2 6859 1 2930
2 6860 1 2930
2 6861 1 2931
2 6862 1 2931
2 6863 1 2931
2 6864 1 2932
2 6865 1 2932
2 6866 1 2938
2 6867 1 2938
2 6868 1 2938
2 6869 1 2938
2 6870 1 2939
2 6871 1 2939
2 6872 1 2939
2 6873 1 2941
2 6874 1 2941
2 6875 1 2941
2 6876 1 2941
2 6877 1 2943
2 6878 1 2943
2 6879 1 2943
2 6880 1 2944
2 6881 1 2944
2 6882 1 2950
2 6883 1 2950
2 6884 1 2950
2 6885 1 2950
2 6886 1 2951
2 6887 1 2951
2 6888 1 2951
2 6889 1 2953
2 6890 1 2953
2 6891 1 2953
2 6892 1 2953
2 6893 1 2955
2 6894 1 2955
2 6895 1 2955
2 6896 1 2956
2 6897 1 2956
2 6898 1 2962
2 6899 1 2962
2 6900 1 2962
2 6901 1 2963
2 6902 1 2963
2 6903 1 2965
2 6904 1 2965
2 6905 1 2965
2 6906 1 2965
2 6907 1 2967
2 6908 1 2967
2 6909 1 2967
2 6910 1 2968
2 6911 1 2968
2 6912 1 2974
2 6913 1 2974
2 6914 1 2975
2 6915 1 2975
2 6916 1 2977
2 6917 1 2977
2 6918 1 2977
2 6919 1 2977
2 6920 1 2979
2 6921 1 2979
2 6922 1 2979
2 6923 1 2980
2 6924 1 2980
2 6925 1 2986
2 6926 1 2986
2 6927 1 2989
2 6928 1 2989
2 6929 1 2989
2 6930 1 2989
2 6931 1 2991
2 6932 1 2991
2 6933 1 2991
2 6934 1 2992
2 6935 1 2992
2 6936 1 2998
2 6937 1 2998
2 6938 1 3001
2 6939 1 3001
2 6940 1 3001
2 6941 1 3003
2 6942 1 3003
2 6943 1 3003
2 6944 1 3006
2 6945 1 3006
2 6946 1 3008
2 6947 1 3008
2 6948 1 3009
2 6949 1 3009
2 6950 1 3009
2 6951 1 3010
2 6952 1 3010
2 6953 1 3012
2 6954 1 3012
2 6955 1 3012
2 6956 1 3016
2 6957 1 3016
2 6958 1 3017
2 6959 1 3017
2 6960 1 3020
2 6961 1 3020
2 6962 1 3021
2 6963 1 3021
2 6964 1 3024
2 6965 1 3024
2 6966 1 3025
2 6967 1 3025
2 6968 1 3028
2 6969 1 3028
2 6970 1 3029
2 6971 1 3029
2 6972 1 3032
2 6973 1 3032
2 6974 1 3033
2 6975 1 3033
2 6976 1 3034
2 6977 1 3034
2 6978 1 3040
2 6979 1 3040
2 6980 1 3040
2 6981 1 3040
2 6982 1 3041
2 6983 1 3041
2 6984 1 3041
2 6985 1 3043
2 6986 1 3043
2 6987 1 3043
2 6988 1 3043
2 6989 1 3045
2 6990 1 3045
2 6991 1 3045
2 6992 1 3046
2 6993 1 3046
2 6994 1 3046
2 6995 1 3047
2 6996 1 3047
2 6997 1 3052
2 6998 1 3052
2 6999 1 3052
2 7000 1 3052
2 7001 1 3053
2 7002 1 3053
2 7003 1 3053
2 7004 1 3054
2 7005 1 3054
2 7006 1 3060
2 7007 1 3060
2 7008 1 3060
2 7009 1 3060
2 7010 1 3061
2 7011 1 3061
2 7012 1 3061
2 7013 1 3063
2 7014 1 3063
2 7015 1 3063
2 7016 1 3063
2 7017 1 3065
2 7018 1 3065
2 7019 1 3065
2 7020 1 3066
2 7021 1 3066
2 7022 1 3072
2 7023 1 3072
2 7024 1 3073
2 7025 1 3073
2 7026 1 3073
2 7027 1 3075
2 7028 1 3075
2 7029 1 3075
2 7030 1 3075
2 7031 1 3077
2 7032 1 3077
2 7033 1 3077
2 7034 1 3078
2 7035 1 3078
2 7036 1 3084
2 7037 1 3084
2 7038 1 3084
2 7039 1 3084
2 7040 1 3085
2 7041 1 3085
2 7042 1 3085
2 7043 1 3087
2 7044 1 3087
2 7045 1 3087
2 7046 1 3087
2 7047 1 3089
2 7048 1 3089
2 7049 1 3089
2 7050 1 3092
2 7051 1 3092
2 7052 1 3093
2 7053 1 3093
2 7054 1 3096
2 7055 1 3096
2 7056 1 3097
2 7057 1 3097
2 7058 1 3100
2 7059 1 3100
2 7060 1 3101
2 7061 1 3101
2 7062 1 3104
2 7063 1 3104
2 7064 1 3105
2 7065 1 3105
2 7066 1 3106
2 7067 1 3106
2 7068 1 3112
2 7069 1 3112
2 7070 1 3113
2 7071 1 3113
2 7072 1 3113
2 7073 1 3115
2 7074 1 3115
2 7075 1 3115
2 7076 1 3115
2 7077 1 3117
2 7078 1 3117
2 7079 1 3117
2 7080 1 3118
2 7081 1 3118
2 7082 1 3118
2 7083 1 3119
2 7084 1 3119
2 7085 1 3124
2 7086 1 3124
2 7087 1 3124
2 7088 1 3124
2 7089 1 3125
2 7090 1 3125
2 7091 1 3125
2 7092 1 3127
2 7093 1 3127
2 7094 1 3130
2 7095 1 3130
2 7096 1 3132
2 7097 1 3132
2 7098 1 3132
2 7099 1 3133
2 7100 1 3133
2 7101 1 3138
2 7102 1 3138
2 7103 1 3138
2 7104 1 3138
2 7105 1 3139
2 7106 1 3139
2 7107 1 3139
2 7108 1 3141
2 7109 1 3141
2 7110 1 3142
2 7111 1 3142
2 7112 1 3144
2 7113 1 3144
2 7114 1 3144
2 7115 1 3145
2 7116 1 3145
2 7117 1 3150
2 7118 1 3150
2 7119 1 3150
2 7120 1 3150
2 7121 1 3151
2 7122 1 3151
2 7123 1 3151
2 7124 1 3152
2 7125 1 3152
2 7126 1 3158
2 7127 1 3158
2 7128 1 3158
2 7129 1 3158
2 7130 1 3159
2 7131 1 3159
2 7132 1 3159
2 7133 1 3161
2 7134 1 3161
2 7135 1 3161
2 7136 1 3163
2 7137 1 3163
2 7138 1 3163
2 7139 1 3163
2 7140 1 3164
2 7141 1 3164
2 7142 1 3164
2 7143 1 3165
2 7144 1 3165
2 7145 1 3168
2 7146 1 3168
2 7147 1 3169
2 7148 1 3169
2 7149 1 3174
2 7150 1 3174
2 7151 1 3174
2 7152 1 3175
2 7153 1 3175
2 7154 1 3177
2 7155 1 3177
2 7156 1 3180
2 7157 1 3180
2 7158 1 3183
2 7159 1 3183
2 7160 1 3186
2 7161 1 3186
2 7162 1 3189
2 7163 1 3189
2 7164 1 3190
2 7165 1 3190
2 7166 1 3190
2 7167 1 3191
2 7168 1 3191
2 7169 1 3196
2 7170 1 3196
2 7171 1 3196
2 7172 1 3196
2 7173 1 3197
2 7174 1 3197
2 7175 1 3197
2 7176 1 3198
2 7177 1 3198
2 7178 1 3198
2 7179 1 3199
2 7180 1 3199
2 7181 1 3204
2 7182 1 3204
2 7183 1 3204
2 7184 1 3204
2 7185 1 3205
2 7186 1 3205
2 7187 1 3205
2 7188 1 3207
2 7189 1 3207
2 7190 1 3210
2 7191 1 3210
2 7192 1 3213
2 7193 1 3213
2 7194 1 3214
2 7195 1 3214
2 7196 1 3218
2 7197 1 3218
2 7198 1 3221
2 7199 1 3221
2 7200 1 3222
2 7201 1 3222
2 7202 1 3222
2 7203 1 3223
2 7204 1 3223
2 7205 1 3228
2 7206 1 3228
2 7207 1 3228
2 7208 1 3228
2 7209 1 3229
2 7210 1 3229
2 7211 1 3229
2 7212 1 3231
2 7213 1 3231
2 7214 1 3234
2 7215 1 3234
2 7216 1 3237
2 7217 1 3237
2 7218 1 3238
2 7219 1 3238
2 7220 1 3242
2 7221 1 3242
2 7222 1 3245
2 7223 1 3245
2 7224 1 3246
2 7225 1 3246
2 7226 1 3246
2 7227 1 3247
2 7228 1 3247
2 7229 1 3252
2 7230 1 3252
2 7231 1 3252
2 7232 1 3252
2 7233 1 3253
2 7234 1 3253
2 7235 1 3253
2 7236 1 3255
2 7237 1 3255
2 7238 1 3258
2 7239 1 3258
2 7240 1 3261
2 7241 1 3261
2 7242 1 3262
2 7243 1 3262
2 7244 1 3266
2 7245 1 3266
2 7246 1 3269
2 7247 1 3269
2 7248 1 3270
2 7249 1 3270
2 7250 1 3270
2 7251 1 3271
2 7252 1 3271
2 7253 1 3276
2 7254 1 3276
2 7255 1 3276
2 7256 1 3276
2 7257 1 3276
2 7258 1 3277
2 7259 1 3277
2 7260 1 3277
2 7261 1 3279
2 7262 1 3279
2 7263 1 3282
2 7264 1 3282
2 7265 1 3285
2 7266 1 3285
2 7267 1 3286
2 7268 1 3286
2 7269 1 3290
2 7270 1 3290
2 7271 1 3293
2 7272 1 3293
2 7273 1 3294
2 7274 1 3294
2 7275 1 3294
2 7276 1 3295
2 7277 1 3295
2 7278 1 3300
2 7279 1 3300
2 7280 1 3300
2 7281 1 3300
2 7282 1 3301
2 7283 1 3301
2 7284 1 3301
2 7285 1 3303
2 7286 1 3303
2 7287 1 3306
2 7288 1 3306
2 7289 1 3309
2 7290 1 3309
2 7291 1 3310
2 7292 1 3310
2 7293 1 3314
2 7294 1 3314
2 7295 1 3317
2 7296 1 3317
2 7297 1 3318
2 7298 1 3318
2 7299 1 3318
2 7300 1 3319
2 7301 1 3319
2 7302 1 3324
2 7303 1 3324
2 7304 1 3324
2 7305 1 3325
2 7306 1 3325
2 7307 1 3325
2 7308 1 3327
2 7309 1 3327
2 7310 1 3330
2 7311 1 3330
2 7312 1 3333
2 7313 1 3333
2 7314 1 3334
2 7315 1 3334
2 7316 1 3338
2 7317 1 3338
2 7318 1 3341
2 7319 1 3341
2 7320 1 3342
2 7321 1 3342
2 7322 1 3343
2 7323 1 3343
2 7324 1 3346
2 7325 1 3346
2 7326 1 3349
2 7327 1 3349
2 7328 1 3352
2 7329 1 3352
2 7330 1 3354
2 7331 1 3354
2 7332 1 3355
2 7333 1 3355
2 7334 1 3355
2 7335 1 3356
2 7336 1 3356
2 7337 1 3356
2 7338 1 3357
2 7339 1 3357
2 7340 1 3357
2 7341 1 3357
2 7342 1 3357
2 7343 1 3360
2 7344 1 3360
2 7345 1 3361
2 7346 1 3361
2 7347 1 3364
2 7348 1 3364
2 7349 1 3367
2 7350 1 3367
2 7351 1 3368
2 7352 1 3368
2 7353 1 3372
2 7354 1 3372
2 7355 1 3375
2 7356 1 3375
2 7357 1 3376
2 7358 1 3376
2 7359 1 3380
2 7360 1 3380
2 7361 1 3383
2 7362 1 3383
2 7363 1 3384
2 7364 1 3384
2 7365 1 3388
2 7366 1 3388
2 7367 1 3391
2 7368 1 3391
2 7369 1 3392
2 7370 1 3392
2 7371 1 3396
2 7372 1 3396
2 7373 1 3399
2 7374 1 3399
2 7375 1 3400
2 7376 1 3400
2 7377 1 3404
2 7378 1 3404
2 7379 1 3407
2 7380 1 3407
2 7381 1 3408
2 7382 1 3408
2 7383 1 3412
2 7384 1 3412
2 7385 1 3415
2 7386 1 3415
2 7387 1 3416
2 7388 1 3416
2 7389 1 3420
2 7390 1 3420
2 7391 1 3423
2 7392 1 3423
2 7393 1 3424
2 7394 1 3424
2 7395 1 3426
2 7396 1 3426
2 7397 1 3430
2 7398 1 3430
2 7399 1 3431
2 7400 1 3431
2 7401 1 3432
2 7402 1 3432
2 7403 1 3438
2 7404 1 3438
2 7405 1 3438
2 7406 1 3438
2 7407 1 3439
2 7408 1 3439
2 7409 1 3439
2 7410 1 3441
2 7411 1 3441
2 7412 1 3441
2 7413 1 3441
2 7414 1 3443
2 7415 1 3443
2 7416 1 3443
2 7417 1 3444
2 7418 1 3444
2 7419 1 3444
2 7420 1 3445
2 7421 1 3445
2 7422 1 3450
2 7423 1 3450
2 7424 1 3450
2 7425 1 3451
2 7426 1 3451
2 7427 1 3453
2 7428 1 3453
2 7429 1 3456
2 7430 1 3456
2 7431 1 3459
2 7432 1 3459
2 7433 1 3462
2 7434 1 3462
2 7435 1 3465
2 7436 1 3465
2 7437 1 3468
2 7438 1 3468
2 7439 1 3471
2 7440 1 3471
2 7441 1 3474
2 7442 1 3474
2 7443 1 3478
2 7444 1 3478
2 7445 1 3484
2 7446 1 3484
2 7447 1 3484
2 7448 1 3484
2 7449 1 3485
2 7450 1 3485
2 7451 1 3485
2 7452 1 3488
2 7453 1 3488
2 7454 1 3492
2 7455 1 3492
2 7456 1 3498
2 7457 1 3498
2 7458 1 3498
2 7459 1 3498
2 7460 1 3499
2 7461 1 3499
2 7462 1 3499
2 7463 1 3502
2 7464 1 3502
2 7465 1 3510
2 7466 1 3510
2 7467 1 3518
2 7468 1 3518
2 7469 1 3522
2 7470 1 3522
2 7471 1 3530
2 7472 1 3530
2 7473 1 3534
2 7474 1 3534
2 7475 1 3540
2 7476 1 3540
2 7477 1 3541
2 7478 1 3541
2 7479 1 3546
2 7480 1 3546
2 7481 1 3554
2 7482 1 3554
2 7483 1 3562
2 7484 1 3562
2 7485 1 3565
2 7486 1 3565
2 7487 1 3567
2 7488 1 3567
2 7489 1 3587
2 7490 1 3587
2 7491 1 3599
2 7492 1 3599
2 7493 1 3614
2 7494 1 3614
2 7495 1 3633
2 7496 1 3633
2 7497 1 3634
2 7498 1 3634
2 7499 1 3634
2 7500 1 3634
2 7501 1 3634
2 7502 1 3636
2 7503 1 3636
2 7504 1 3636
2 7505 1 3636
2 7506 1 3636
2 7507 1 3638
2 7508 1 3638
2 7509 1 3638
2 7510 1 3638
2 7511 1 3640
2 7512 1 3640
2 7513 1 3640
2 7514 1 3642
2 7515 1 3642
2 7516 1 3642
2 7517 1 3642
2 7518 1 3644
2 7519 1 3644
2 7520 1 3644
2 7521 1 3647
2 7522 1 3647
2 7523 1 3648
2 7524 1 3648
2 7525 1 3651
2 7526 1 3651
2 7527 1 3652
2 7528 1 3652
2 7529 1 3655
2 7530 1 3655
2 7531 1 3655
2 7532 1 3656
2 7533 1 3656
2 7534 1 3656
2 7535 1 3659
2 7536 1 3659
2 7537 1 3659
2 7538 1 3660
2 7539 1 3660
2 7540 1 3661
2 7541 1 3661
2 7542 1 3661
2 7543 1 3662
2 7544 1 3662
2 7545 1 3667
2 7546 1 3667
2 7547 1 3667
2 7548 1 3668
2 7549 1 3668
2 7550 1 3671
2 7551 1 3671
2 7552 1 3674
2 7553 1 3674
2 7554 1 3682
2 7555 1 3682
2 7556 1 3682
2 7557 1 3683
2 7558 1 3683
2 7559 1 3688
2 7560 1 3688
2 7561 1 3688
2 7562 1 3688
2 7563 1 3689
2 7564 1 3689
2 7565 1 3694
2 7566 1 3694
2 7567 1 3701
2 7568 1 3701
2 7569 1 3701
2 7570 1 3702
2 7571 1 3702
2 7572 1 3707
2 7573 1 3707
2 7574 1 3710
2 7575 1 3710
2 7576 1 3711
2 7577 1 3711
2 7578 1 3729
2 7579 1 3729
2 7580 1 3730
2 7581 1 3730
2 7582 1 3733
2 7583 1 3733
2 7584 1 3734
2 7585 1 3734
2 7586 1 3737
2 7587 1 3737
2 7588 1 3738
2 7589 1 3738
2 7590 1 3741
2 7591 1 3741
2 7592 1 3742
2 7593 1 3742
2 7594 1 3745
2 7595 1 3745
2 7596 1 3746
2 7597 1 3746
2 7598 1 3749
2 7599 1 3749
2 7600 1 3750
2 7601 1 3750
2 7602 1 3753
2 7603 1 3753
2 7604 1 3754
2 7605 1 3754
2 7606 1 3757
2 7607 1 3757
2 7608 1 3758
2 7609 1 3758
2 7610 1 3761
2 7611 1 3761
2 7612 1 3762
2 7613 1 3762
2 7614 1 3765
2 7615 1 3765
2 7616 1 3766
2 7617 1 3766
2 7618 1 3769
2 7619 1 3769
2 7620 1 3770
2 7621 1 3770
2 7622 1 3773
2 7623 1 3773
2 7624 1 3774
2 7625 1 3774
2 7626 1 3777
2 7627 1 3777
2 7628 1 3778
2 7629 1 3778
2 7630 1 3781
2 7631 1 3781
2 7632 1 3782
2 7633 1 3782
2 7634 1 3785
2 7635 1 3785
2 7636 1 3785
2 7637 1 3786
2 7638 1 3786
2 7639 1 3789
2 7640 1 3789
2 7641 1 3789
2 7642 1 3789
2 7643 1 3789
2 7644 1 3790
2 7645 1 3790
2 7646 1 3790
2 7647 1 3790
2 7648 1 3792
2 7649 1 3792
2 7650 1 3795
2 7651 1 3795
2 7652 1 3798
2 7653 1 3798
2 7654 1 3821
2 7655 1 3821
2 7656 1 3821
2 7657 1 3822
2 7658 1 3822
2 7659 1 3822
2 7660 1 3827
2 7661 1 3827
2 7662 1 3827
2 7663 1 3827
2 7664 1 3828
2 7665 1 3828
2 7666 1 3828
2 7667 1 3830
2 7668 1 3830
2 7669 1 3835
2 7670 1 3835
2 7671 1 3835
2 7672 1 3835
2 7673 1 3836
2 7674 1 3836
2 7675 1 3836
2 7676 1 3839
2 7677 1 3839
2 7678 1 3842
2 7679 1 3842
2 7680 1 3843
2 7681 1 3843
2 7682 1 3849
2 7683 1 3849
2 7684 1 3849
2 7685 1 3850
2 7686 1 3850
2 7687 1 3850
2 7688 1 3852
2 7689 1 3852
2 7690 1 3855
2 7691 1 3855
2 7692 1 3861
2 7693 1 3861
2 7694 1 3861
2 7695 1 3861
2 7696 1 3862
2 7697 1 3862
2 7698 1 3862
2 7699 1 3864
2 7700 1 3864
2 7701 1 3867
2 7702 1 3867
2 7703 1 3870
2 7704 1 3870
2 7705 1 3875
2 7706 1 3875
2 7707 1 3875
2 7708 1 3875
2 7709 1 3876
2 7710 1 3876
2 7711 1 3876
2 7712 1 3881
2 7713 1 3881
2 7714 1 3881
2 7715 1 3881
2 7716 1 3882
2 7717 1 3882
2 7718 1 3882
2 7719 1 3884
2 7720 1 3884
2 7721 1 3887
2 7722 1 3887
2 7723 1 3890
2 7724 1 3890
2 7725 1 3891
2 7726 1 3891
2 7727 1 3895
2 7728 1 3895
2 7729 1 3898
2 7730 1 3898
2 7731 1 3903
2 7732 1 3903
2 7733 1 3903
2 7734 1 3903
2 7735 1 3904
2 7736 1 3904
2 7737 1 3904
2 7738 1 3906
2 7739 1 3906
2 7740 1 3909
2 7741 1 3909
2 7742 1 3912
2 7743 1 3912
2 7744 1 3913
2 7745 1 3913
2 7746 1 3917
2 7747 1 3917
2 7748 1 3920
2 7749 1 3920
2 7750 1 3925
2 7751 1 3925
2 7752 1 3925
2 7753 1 3925
2 7754 1 3926
2 7755 1 3926
2 7756 1 3926
2 7757 1 3928
2 7758 1 3928
2 7759 1 3931
2 7760 1 3931
2 7761 1 3934
2 7762 1 3934
2 7763 1 3935
2 7764 1 3935
2 7765 1 3939
2 7766 1 3939
2 7767 1 3942
2 7768 1 3942
2 7769 1 3947
2 7770 1 3947
2 7771 1 3947
2 7772 1 3947
2 7773 1 3948
2 7774 1 3948
2 7775 1 3948
2 7776 1 3948
2 7777 1 3950
2 7778 1 3950
2 7779 1 3953
2 7780 1 3953
2 7781 1 3956
2 7782 1 3956
2 7783 1 3957
2 7784 1 3957
2 7785 1 3961
2 7786 1 3961
2 7787 1 3964
2 7788 1 3964
2 7789 1 3969
2 7790 1 3969
2 7791 1 3969
2 7792 1 3969
2 7793 1 3970
2 7794 1 3970
2 7795 1 3972
2 7796 1 3972
2 7797 1 3975
2 7798 1 3975
2 7799 1 3978
2 7800 1 3978
2 7801 1 3979
2 7802 1 3979
2 7803 1 3983
2 7804 1 3983
2 7805 1 3986
2 7806 1 3986
2 7807 1 3991
2 7808 1 3991
2 7809 1 3991
2 7810 1 3992
2 7811 1 3992
2 7812 1 3992
2 7813 1 3994
2 7814 1 3994
2 7815 1 3997
2 7816 1 3997
2 7817 1 4000
2 7818 1 4000
2 7819 1 4001
2 7820 1 4001
2 7821 1 4005
2 7822 1 4005
2 7823 1 4008
2 7824 1 4008
2 7825 1 4009
2 7826 1 4009
2 7827 1 4010
2 7828 1 4010
2 7829 1 4013
2 7830 1 4013
2 7831 1 4016
2 7832 1 4016
2 7833 1 4019
2 7834 1 4019
2 7835 1 4023
2 7836 1 4023
2 7837 1 4024
2 7838 1 4024
2 7839 1 4027
2 7840 1 4027
2 7841 1 4030
2 7842 1 4030
2 7843 1 4031
2 7844 1 4031
2 7845 1 4035
2 7846 1 4035
2 7847 1 4038
2 7848 1 4038
2 7849 1 4039
2 7850 1 4039
2 7851 1 4043
2 7852 1 4043
2 7853 1 4046
2 7854 1 4046
2 7855 1 4047
2 7856 1 4047
2 7857 1 4051
2 7858 1 4051
2 7859 1 4054
2 7860 1 4054
2 7861 1 4055
2 7862 1 4055
2 7863 1 4059
2 7864 1 4059
2 7865 1 4062
2 7866 1 4062
2 7867 1 4063
2 7868 1 4063
2 7869 1 4067
2 7870 1 4067
2 7871 1 4070
2 7872 1 4070
2 7873 1 4071
2 7874 1 4071
2 7875 1 4075
2 7876 1 4075
2 7877 1 4078
2 7878 1 4078
2 7879 1 4079
2 7880 1 4079
2 7881 1 4083
2 7882 1 4083
2 7883 1 4086
2 7884 1 4086
2 7885 1 4087
2 7886 1 4087
2 7887 1 4089
2 7888 1 4089
2 7889 1 4095
2 7890 1 4095
2 7891 1 4096
2 7892 1 4096
2 7893 1 4098
2 7894 1 4098
2 7895 1 4101
2 7896 1 4101
2 7897 1 4104
2 7898 1 4104
2 7899 1 4107
2 7900 1 4107
2 7901 1 4110
2 7902 1 4110
2 7903 1 4113
2 7904 1 4113
2 7905 1 4116
2 7906 1 4116
2 7907 1 4119
2 7908 1 4119
2 7909 1 4125
2 7910 1 4125
2 7911 1 4131
2 7912 1 4131
2 7913 1 4139
2 7914 1 4139
2 7915 1 4147
2 7916 1 4147
2 7917 1 4151
2 7918 1 4151
2 7919 1 4159
2 7920 1 4159
2 7921 1 4163
2 7922 1 4163
2 7923 1 4169
2 7924 1 4169
2 7925 1 4170
2 7926 1 4170
2 7927 1 4175
2 7928 1 4175
2 7929 1 4183
2 7930 1 4183
2 7931 1 4191
2 7932 1 4191
2 7933 1 4211
2 7934 1 4211
2 7935 1 4223
2 7936 1 4223
2 7937 1 4238
2 7938 1 4238
2 7939 1 4261
2 7940 1 4261
2 7941 1 4269
2 7942 1 4269
2 7943 1 4269
2 7944 1 4270
2 7945 1 4270
2 7946 1 4270
2 7947 1 4281
2 7948 1 4281
2 7949 1 4281
2 7950 1 4281
2 7951 1 4281
2 7952 1 4282
2 7953 1 4282
2 7954 1 4282
2 7955 1 4284
2 7956 1 4284
2 7957 1 4287
2 7958 1 4287
2 7959 1 4290
2 7960 1 4290
2 7961 1 4306
2 7962 1 4306
2 7963 1 4310
2 7964 1 4310
2 7965 1 4313
2 7966 1 4313
2 7967 1 4322
2 7968 1 4322
0 50 5 5 1 49
0 51 5 6 1 4372
0 52 5 6 1 4377
0 53 5 6 1 4383
0 54 5 6 1 4389
0 55 5 5 1 4395
0 56 5 6 1 4402
0 57 5 6 1 4409
0 58 5 5 1 4415
0 59 5 6 1 4422
0 60 5 6 1 4428
0 61 5 5 1 4434
0 62 5 6 1 4441
0 63 5 6 1 4448
0 64 5 5 1 4454
0 65 5 6 1 4461
0 66 5 6 1 4467
0 67 5 5 1 4473
0 68 5 6 1 4480
0 69 5 7 1 4487
0 70 5 6 1 4493
0 71 5 7 1 4500
0 72 5 7 1 4506
0 73 5 6 1 4512
0 74 5 7 1 4519
0 75 5 7 1 4526
0 76 5 6 1 4532
0 77 5 7 1 4539
0 78 5 7 1 4545
0 79 5 6 1 4551
0 80 5 7 1 4558
0 81 5 7 1 4565
0 82 5 5 1 4571
0 83 5 6 1 4578
0 84 5 6 1 4584
0 85 5 5 1 4590
0 86 5 6 1 4597
0 87 5 6 1 4604
0 88 5 5 1 4610
0 89 5 6 1 4617
0 90 5 6 1 4623
0 91 5 5 1 4629
0 92 5 6 1 4636
0 93 5 5 1 4643
0 94 5 6 1 4650
0 95 5 6 1 4657
0 96 5 5 1 4665
0 97 5 3 1 4673
0 98 5 4 1 4680
0 99 7 1 2 4666 4968
0 100 5 1 1 99
0 101 7 1 2 4960 4674
0 102 7 1 2 4681 101
0 103 5 2 1 102
0 104 7 2 2 100 4972
0 105 7 2 2 4954 4974
0 106 5 1 1 4976
0 107 7 1 2 4675 4977
0 108 5 1 1 107
0 109 7 2 2 4965 4682
0 110 5 1 1 4978
0 111 7 2 2 4961 4979
0 112 5 2 1 4980
0 113 7 1 2 4658 4981
0 114 5 1 1 113
0 115 7 2 2 108 114
0 116 5 2 1 4984
0 117 7 1 2 4676 4973
0 118 7 1 2 106 117
0 119 5 1 1 118
0 120 7 2 2 4982 119
0 121 5 1 1 4988
0 122 7 1 2 4955 121
0 123 5 2 1 122
0 124 7 1 2 4659 4989
0 125 5 1 1 124
0 126 7 2 2 4990 125
0 127 5 1 1 4992
0 128 7 2 2 4948 4993
0 129 5 2 1 4994
0 130 7 1 2 4975 4991
0 131 5 1 1 130
0 132 7 2 2 4677 4969
0 133 5 2 1 4998
0 134 7 2 2 4667 4999
0 135 5 1 1 5002
0 136 7 1 2 4956 5003
0 137 5 1 1 136
0 138 7 2 2 131 137
0 139 5 1 1 5004
0 140 7 1 2 4996 5005
0 141 5 2 1 140
0 142 7 2 2 4985 5006
0 143 5 1 1 5008
0 144 7 1 2 4949 143
0 145 5 2 1 144
0 146 7 1 2 4651 5009
0 147 5 1 1 146
0 148 7 2 2 5010 147
0 149 5 1 1 5012
0 150 7 2 2 4943 5013
0 151 5 2 1 5014
0 152 7 1 2 127 5011
0 153 5 1 1 152
0 154 7 1 2 4986 4995
0 155 5 1 1 154
0 156 7 2 2 153 155
0 157 5 1 1 5018
0 158 7 1 2 5016 157
0 159 5 2 1 158
0 160 7 1 2 4987 4997
0 161 5 1 1 160
0 162 7 1 2 139 161
0 163 5 1 1 162
0 164 7 3 2 5007 163
0 165 5 1 1 5022
0 166 7 1 2 5017 5023
0 167 5 1 1 166
0 168 7 1 2 5019 167
0 169 5 1 1 168
0 170 7 3 2 5020 169
0 171 5 1 1 5025
0 172 7 2 2 5021 165
0 173 5 1 1 5028
0 174 7 1 2 4944 173
0 175 5 2 1 174
0 176 7 1 2 4644 5029
0 177 5 1 1 176
0 178 7 2 2 5030 177
0 179 5 1 1 5032
0 180 7 2 2 4937 5033
0 181 5 2 1 5034
0 182 7 1 2 149 5031
0 183 5 1 1 182
0 184 7 1 2 5015 5024
0 185 5 1 1 184
0 186 7 2 2 183 185
0 187 5 1 1 5038
0 188 7 1 2 5036 187
0 189 5 2 1 188
0 190 7 2 2 171 5040
0 191 5 1 1 5042
0 192 7 1 2 4938 191
0 193 5 2 1 192
0 194 7 1 2 4637 5043
0 195 5 1 1 194
0 196 7 2 2 5044 195
0 197 5 1 1 5046
0 198 7 2 2 4932 5047
0 199 5 2 1 5048
0 200 7 1 2 179 5045
0 201 5 1 1 200
0 202 7 1 2 5026 5035
0 203 5 1 1 202
0 204 7 2 2 201 203
0 205 5 1 1 5052
0 206 7 1 2 5050 205
0 207 5 2 1 206
0 208 7 1 2 5027 5037
0 209 5 1 1 208
0 210 7 1 2 5039 209
0 211 5 1 1 210
0 212 7 3 2 5041 211
0 213 5 1 1 5056
0 214 7 1 2 5051 5057
0 215 5 1 1 214
0 216 7 1 2 5053 215
0 217 5 1 1 216
0 218 7 3 2 5054 217
0 219 5 1 1 5059
0 220 7 2 2 5055 213
0 221 5 1 1 5062
0 222 7 1 2 4933 221
0 223 5 2 1 222
0 224 7 1 2 4630 5063
0 225 5 1 1 224
0 226 7 2 2 5064 225
0 227 5 1 1 5066
0 228 7 2 2 4926 5067
0 229 5 2 1 5068
0 230 7 1 2 197 5065
0 231 5 1 1 230
0 232 7 1 2 5049 5058
0 233 5 1 1 232
0 234 7 2 2 231 233
0 235 5 1 1 5072
0 236 7 1 2 5070 235
0 237 5 2 1 236
0 238 7 2 2 219 5074
0 239 5 1 1 5076
0 240 7 1 2 4927 239
0 241 5 2 1 240
0 242 7 1 2 4624 5077
0 243 5 1 1 242
0 244 7 2 2 5078 243
0 245 5 1 1 5080
0 246 7 2 2 4920 5081
0 247 5 2 1 5082
0 248 7 1 2 227 5079
0 249 5 1 1 248
0 250 7 1 2 5060 5069
0 251 5 1 1 250
0 252 7 2 2 249 251
0 253 5 1 1 5086
0 254 7 1 2 5084 253
0 255 5 2 1 254
0 256 7 1 2 5061 5071
0 257 5 1 1 256
0 258 7 1 2 5073 257
0 259 5 1 1 258
0 260 7 3 2 5075 259
0 261 5 1 1 5090
0 262 7 1 2 5085 5091
0 263 5 1 1 262
0 264 7 1 2 5087 263
0 265 5 1 1 264
0 266 7 3 2 5088 265
0 267 5 1 1 5093
0 268 7 2 2 5089 261
0 269 5 1 1 5096
0 270 7 1 2 4921 269
0 271 5 2 1 270
0 272 7 1 2 4618 5097
0 273 5 1 1 272
0 274 7 2 2 5098 273
0 275 5 1 1 5100
0 276 7 2 2 4915 5101
0 277 5 2 1 5102
0 278 7 1 2 245 5099
0 279 5 1 1 278
0 280 7 1 2 5083 5092
0 281 5 1 1 280
0 282 7 2 2 279 281
0 283 5 1 1 5106
0 284 7 1 2 5104 283
0 285 5 2 1 284
0 286 7 2 2 267 5108
0 287 5 1 1 5110
0 288 7 1 2 4916 287
0 289 5 2 1 288
0 290 7 1 2 4611 5111
0 291 5 1 1 290
0 292 7 2 2 5112 291
0 293 5 1 1 5114
0 294 7 2 2 4909 5115
0 295 5 2 1 5116
0 296 7 1 2 275 5113
0 297 5 1 1 296
0 298 7 1 2 5094 5103
0 299 5 1 1 298
0 300 7 2 2 297 299
0 301 5 1 1 5120
0 302 7 1 2 5118 301
0 303 5 2 1 302
0 304 7 1 2 5095 5105
0 305 5 1 1 304
0 306 7 1 2 5107 305
0 307 5 1 1 306
0 308 7 3 2 5109 307
0 309 5 1 1 5124
0 310 7 1 2 5119 5125
0 311 5 1 1 310
0 312 7 1 2 5121 311
0 313 5 1 1 312
0 314 7 3 2 5122 313
0 315 5 1 1 5127
0 316 7 2 2 5123 309
0 317 5 1 1 5130
0 318 7 1 2 4910 317
0 319 5 2 1 318
0 320 7 1 2 4605 5131
0 321 5 1 1 320
0 322 7 2 2 5132 321
0 323 5 1 1 5134
0 324 7 2 2 4903 5135
0 325 5 2 1 5136
0 326 7 1 2 293 5133
0 327 5 1 1 326
0 328 7 1 2 5117 5126
0 329 5 1 1 328
0 330 7 2 2 327 329
0 331 5 1 1 5140
0 332 7 1 2 5138 331
0 333 5 2 1 332
0 334 7 2 2 315 5142
0 335 5 1 1 5144
0 336 7 1 2 4904 335
0 337 5 2 1 336
0 338 7 1 2 4598 5145
0 339 5 1 1 338
0 340 7 2 2 5146 339
0 341 5 1 1 5148
0 342 7 2 2 4898 5149
0 343 5 2 1 5150
0 344 7 1 2 323 5147
0 345 5 1 1 344
0 346 7 1 2 5128 5137
0 347 5 1 1 346
0 348 7 2 2 345 347
0 349 5 1 1 5154
0 350 7 1 2 5152 349
0 351 5 2 1 350
0 352 7 1 2 5129 5139
0 353 5 1 1 352
0 354 7 1 2 5141 353
0 355 5 1 1 354
0 356 7 3 2 5143 355
0 357 5 1 1 5158
0 358 7 1 2 5153 5159
0 359 5 1 1 358
0 360 7 1 2 5155 359
0 361 5 1 1 360
0 362 7 3 2 5156 361
0 363 5 1 1 5161
0 364 7 2 2 5157 357
0 365 5 1 1 5164
0 366 7 1 2 4899 365
0 367 5 2 1 366
0 368 7 1 2 4591 5165
0 369 5 1 1 368
0 370 7 2 2 5166 369
0 371 5 1 1 5168
0 372 7 2 2 4892 5169
0 373 5 2 1 5170
0 374 7 1 2 341 5167
0 375 5 1 1 374
0 376 7 1 2 5151 5160
0 377 5 1 1 376
0 378 7 2 2 375 377
0 379 5 1 1 5174
0 380 7 1 2 5172 379
0 381 5 2 1 380
0 382 7 2 2 363 5176
0 383 5 1 1 5178
0 384 7 1 2 4893 383
0 385 5 2 1 384
0 386 7 1 2 4585 5179
0 387 5 1 1 386
0 388 7 2 2 5180 387
0 389 5 1 1 5182
0 390 7 2 2 4886 5183
0 391 5 2 1 5184
0 392 7 1 2 371 5181
0 393 5 1 1 392
0 394 7 1 2 5162 5171
0 395 5 1 1 394
0 396 7 2 2 393 395
0 397 5 1 1 5188
0 398 7 1 2 5186 397
0 399 5 2 1 398
0 400 7 1 2 5163 5173
0 401 5 1 1 400
0 402 7 1 2 5175 401
0 403 5 1 1 402
0 404 7 3 2 5177 403
0 405 5 1 1 5192
0 406 7 1 2 5187 5193
0 407 5 1 1 406
0 408 7 1 2 5189 407
0 409 5 1 1 408
0 410 7 3 2 5190 409
0 411 5 1 1 5195
0 412 7 2 2 5191 405
0 413 5 1 1 5198
0 414 7 1 2 4887 413
0 415 5 2 1 414
0 416 7 1 2 4579 5199
0 417 5 1 1 416
0 418 7 2 2 5200 417
0 419 5 1 1 5202
0 420 7 2 2 4881 5203
0 421 5 2 1 5204
0 422 7 1 2 389 5201
0 423 5 1 1 422
0 424 7 1 2 5185 5194
0 425 5 1 1 424
0 426 7 2 2 423 425
0 427 5 1 1 5208
0 428 7 1 2 5206 427
0 429 5 2 1 428
0 430 7 2 2 411 5210
0 431 5 1 1 5212
0 432 7 1 2 4882 431
0 433 5 2 1 432
0 434 7 1 2 4572 5213
0 435 5 1 1 434
0 436 7 2 2 5214 435
0 437 5 1 1 5216
0 438 7 2 2 4874 5217
0 439 5 2 1 5218
0 440 7 1 2 419 5215
0 441 5 1 1 440
0 442 7 1 2 5196 5205
0 443 5 1 1 442
0 444 7 2 2 441 443
0 445 5 1 1 5222
0 446 7 1 2 5220 445
0 447 5 2 1 446
0 448 7 1 2 5197 5207
0 449 5 1 1 448
0 450 7 1 2 5209 449
0 451 5 1 1 450
0 452 7 3 2 5211 451
0 453 5 1 1 5226
0 454 7 1 2 5221 5227
0 455 5 1 1 454
0 456 7 1 2 5223 455
0 457 5 1 1 456
0 458 7 3 2 5224 457
0 459 5 1 1 5229
0 460 7 2 2 5225 453
0 461 5 1 1 5232
0 462 7 1 2 4875 461
0 463 5 2 1 462
0 464 7 1 2 4566 5233
0 465 5 1 1 464
0 466 7 2 2 5234 465
0 467 5 1 1 5236
0 468 7 2 2 4867 5237
0 469 5 2 1 5238
0 470 7 1 2 437 5235
0 471 5 1 1 470
0 472 7 1 2 5219 5228
0 473 5 1 1 472
0 474 7 2 2 471 473
0 475 5 1 1 5242
0 476 7 1 2 5240 475
0 477 5 2 1 476
0 478 7 2 2 459 5244
0 479 5 1 1 5246
0 480 7 1 2 4868 479
0 481 5 2 1 480
0 482 7 1 2 4559 5247
0 483 5 1 1 482
0 484 7 2 2 5248 483
0 485 5 1 1 5250
0 486 7 2 2 4861 5251
0 487 5 2 1 5252
0 488 7 1 2 467 5249
0 489 5 1 1 488
0 490 7 1 2 5230 5239
0 491 5 1 1 490
0 492 7 2 2 489 491
0 493 5 1 1 5256
0 494 7 1 2 5254 493
0 495 5 2 1 494
0 496 7 1 2 5231 5241
0 497 5 1 1 496
0 498 7 1 2 5243 497
0 499 5 1 1 498
0 500 7 3 2 5245 499
0 501 5 1 1 5260
0 502 7 1 2 5255 5261
0 503 5 1 1 502
0 504 7 1 2 5257 503
0 505 5 1 1 504
0 506 7 3 2 5258 505
0 507 5 1 1 5263
0 508 7 2 2 5259 501
0 509 5 1 1 5266
0 510 7 1 2 4862 509
0 511 5 2 1 510
0 512 7 1 2 4552 5267
0 513 5 1 1 512
0 514 7 2 2 5268 513
0 515 5 1 1 5270
0 516 7 2 2 4854 5271
0 517 5 2 1 5272
0 518 7 1 2 485 5269
0 519 5 1 1 518
0 520 7 1 2 5253 5262
0 521 5 1 1 520
0 522 7 2 2 519 521
0 523 5 1 1 5276
0 524 7 1 2 5274 523
0 525 5 2 1 524
0 526 7 2 2 507 5278
0 527 5 1 1 5280
0 528 7 1 2 4855 527
0 529 5 2 1 528
0 530 7 1 2 4546 5281
0 531 5 1 1 530
0 532 7 2 2 5282 531
0 533 5 1 1 5284
0 534 7 2 2 4847 5285
0 535 5 2 1 5286
0 536 7 1 2 515 5283
0 537 5 1 1 536
0 538 7 1 2 5264 5273
0 539 5 1 1 538
0 540 7 2 2 537 539
0 541 5 1 1 5290
0 542 7 1 2 5288 541
0 543 5 2 1 542
0 544 7 1 2 5265 5275
0 545 5 1 1 544
0 546 7 1 2 5277 545
0 547 5 1 1 546
0 548 7 3 2 5279 547
0 549 5 1 1 5294
0 550 7 1 2 5289 5295
0 551 5 1 1 550
0 552 7 1 2 5291 551
0 553 5 1 1 552
0 554 7 3 2 5292 553
0 555 5 1 1 5297
0 556 7 2 2 5293 549
0 557 5 1 1 5300
0 558 7 1 2 4848 557
0 559 5 2 1 558
0 560 7 1 2 4540 5301
0 561 5 1 1 560
0 562 7 2 2 5302 561
0 563 5 1 1 5304
0 564 7 2 2 4841 5305
0 565 5 2 1 5306
0 566 7 1 2 533 5303
0 567 5 1 1 566
0 568 7 1 2 5287 5296
0 569 5 1 1 568
0 570 7 2 2 567 569
0 571 5 1 1 5310
0 572 7 1 2 5308 571
0 573 5 2 1 572
0 574 7 2 2 555 5312
0 575 5 1 1 5314
0 576 7 1 2 4842 575
0 577 5 2 1 576
0 578 7 1 2 4533 5315
0 579 5 1 1 578
0 580 7 2 2 5316 579
0 581 5 1 1 5318
0 582 7 2 2 4834 5319
0 583 5 2 1 5320
0 584 7 1 2 563 5317
0 585 5 1 1 584
0 586 7 1 2 5298 5307
0 587 5 1 1 586
0 588 7 2 2 585 587
0 589 5 1 1 5324
0 590 7 1 2 5322 589
0 591 5 2 1 590
0 592 7 1 2 5299 5309
0 593 5 1 1 592
0 594 7 1 2 5311 593
0 595 5 1 1 594
0 596 7 3 2 5313 595
0 597 5 1 1 5328
0 598 7 1 2 5323 5329
0 599 5 1 1 598
0 600 7 1 2 5325 599
0 601 5 1 1 600
0 602 7 3 2 5326 601
0 603 5 1 1 5331
0 604 7 2 2 5327 597
0 605 5 1 1 5334
0 606 7 1 2 4835 605
0 607 5 2 1 606
0 608 7 1 2 4527 5335
0 609 5 1 1 608
0 610 7 2 2 5336 609
0 611 5 1 1 5338
0 612 7 2 2 4827 5339
0 613 5 2 1 5340
0 614 7 1 2 581 5337
0 615 5 1 1 614
0 616 7 1 2 5321 5330
0 617 5 1 1 616
0 618 7 2 2 615 617
0 619 5 1 1 5344
0 620 7 1 2 5342 619
0 621 5 2 1 620
0 622 7 2 2 603 5346
0 623 5 1 1 5348
0 624 7 1 2 4828 623
0 625 5 2 1 624
0 626 7 1 2 4520 5349
0 627 5 1 1 626
0 628 7 2 2 5350 627
0 629 5 1 1 5352
0 630 7 2 2 4821 5353
0 631 5 2 1 5354
0 632 7 1 2 611 5351
0 633 5 1 1 632
0 634 7 1 2 5332 5341
0 635 5 1 1 634
0 636 7 2 2 633 635
0 637 5 1 1 5358
0 638 7 1 2 5356 637
0 639 5 2 1 638
0 640 7 1 2 5333 5343
0 641 5 1 1 640
0 642 7 1 2 5345 641
0 643 5 1 1 642
0 644 7 3 2 5347 643
0 645 5 1 1 5362
0 646 7 1 2 5357 5363
0 647 5 1 1 646
0 648 7 1 2 5359 647
0 649 5 1 1 648
0 650 7 3 2 5360 649
0 651 5 1 1 5365
0 652 7 2 2 5361 645
0 653 5 1 1 5368
0 654 7 1 2 4822 653
0 655 5 2 1 654
0 656 7 1 2 4513 5369
0 657 5 1 1 656
0 658 7 2 2 5370 657
0 659 5 1 1 5372
0 660 7 2 2 4814 5373
0 661 5 2 1 5374
0 662 7 1 2 629 5371
0 663 5 1 1 662
0 664 7 1 2 5355 5364
0 665 5 1 1 664
0 666 7 2 2 663 665
0 667 5 1 1 5378
0 668 7 1 2 5376 667
0 669 5 2 1 668
0 670 7 2 2 651 5380
0 671 5 1 1 5382
0 672 7 1 2 4815 671
0 673 5 2 1 672
0 674 7 1 2 4507 5383
0 675 5 1 1 674
0 676 7 2 2 5384 675
0 677 5 1 1 5386
0 678 7 2 2 4807 5387
0 679 5 2 1 5388
0 680 7 1 2 659 5385
0 681 5 1 1 680
0 682 7 1 2 5366 5375
0 683 5 1 1 682
0 684 7 2 2 681 683
0 685 5 1 1 5392
0 686 7 1 2 5390 685
0 687 5 2 1 686
0 688 7 1 2 5367 5377
0 689 5 1 1 688
0 690 7 1 2 5379 689
0 691 5 1 1 690
0 692 7 3 2 5381 691
0 693 5 1 1 5396
0 694 7 1 2 5391 5397
0 695 5 1 1 694
0 696 7 1 2 5393 695
0 697 5 1 1 696
0 698 7 3 2 5394 697
0 699 5 1 1 5399
0 700 7 2 2 5395 693
0 701 5 1 1 5402
0 702 7 1 2 4808 701
0 703 5 2 1 702
0 704 7 1 2 4501 5403
0 705 5 1 1 704
0 706 7 2 2 5404 705
0 707 5 1 1 5406
0 708 7 2 2 4801 5407
0 709 5 2 1 5408
0 710 7 1 2 677 5405
0 711 5 1 1 710
0 712 7 1 2 5389 5398
0 713 5 1 1 712
0 714 7 2 2 711 713
0 715 5 1 1 5412
0 716 7 1 2 5410 715
0 717 5 2 1 716
0 718 7 2 2 699 5414
0 719 5 1 1 5416
0 720 7 1 2 4802 719
0 721 5 2 1 720
0 722 7 1 2 4494 5417
0 723 5 1 1 722
0 724 7 2 2 5418 723
0 725 5 1 1 5420
0 726 7 2 2 4794 5421
0 727 5 2 1 5422
0 728 7 1 2 707 5419
0 729 5 1 1 728
0 730 7 1 2 5400 5409
0 731 5 1 1 730
0 732 7 2 2 729 731
0 733 5 1 1 5426
0 734 7 1 2 5424 733
0 735 5 2 1 734
0 736 7 1 2 5401 5411
0 737 5 1 1 736
0 738 7 1 2 5413 737
0 739 5 1 1 738
0 740 7 3 2 5415 739
0 741 5 1 1 5430
0 742 7 1 2 5425 5431
0 743 5 1 1 742
0 744 7 1 2 5427 743
0 745 5 1 1 744
0 746 7 3 2 5428 745
0 747 5 1 1 5433
0 748 7 2 2 5429 741
0 749 5 1 1 5436
0 750 7 1 2 4795 749
0 751 5 2 1 750
0 752 7 1 2 4488 5437
0 753 5 1 1 752
0 754 7 2 2 5438 753
0 755 5 1 1 5440
0 756 7 2 2 4788 5441
0 757 5 2 1 5442
0 758 7 1 2 725 5439
0 759 5 1 1 758
0 760 7 1 2 5423 5432
0 761 5 1 1 760
0 762 7 2 2 759 761
0 763 5 1 1 5446
0 764 7 1 2 5444 763
0 765 5 2 1 764
0 766 7 2 2 747 5448
0 767 5 1 1 5450
0 768 7 1 2 4789 767
0 769 5 2 1 768
0 770 7 1 2 4481 5451
0 771 5 1 1 770
0 772 7 2 2 5452 771
0 773 5 1 1 5454
0 774 7 2 2 4783 5455
0 775 5 2 1 5456
0 776 7 1 2 755 5453
0 777 5 1 1 776
0 778 7 1 2 5434 5443
0 779 5 1 1 778
0 780 7 2 2 777 779
0 781 5 1 1 5460
0 782 7 1 2 5458 781
0 783 5 2 1 782
0 784 7 1 2 5435 5445
0 785 5 1 1 784
0 786 7 1 2 5447 785
0 787 5 1 1 786
0 788 7 3 2 5449 787
0 789 5 1 1 5464
0 790 7 1 2 5459 5465
0 791 5 1 1 790
0 792 7 1 2 5461 791
0 793 5 1 1 792
0 794 7 3 2 5462 793
0 795 5 1 1 5467
0 796 7 2 2 5463 789
0 797 5 1 1 5470
0 798 7 1 2 4784 797
0 799 5 2 1 798
0 800 7 1 2 4474 5471
0 801 5 1 1 800
0 802 7 2 2 5472 801
0 803 5 1 1 5474
0 804 7 2 2 4777 5475
0 805 5 2 1 5476
0 806 7 1 2 773 5473
0 807 5 1 1 806
0 808 7 1 2 5457 5466
0 809 5 1 1 808
0 810 7 2 2 807 809
0 811 5 1 1 5480
0 812 7 1 2 5478 811
0 813 5 2 1 812
0 814 7 2 2 795 5482
0 815 5 1 1 5484
0 816 7 1 2 4778 815
0 817 5 2 1 816
0 818 7 1 2 4468 5485
0 819 5 1 1 818
0 820 7 2 2 5486 819
0 821 5 1 1 5488
0 822 7 2 2 4771 5489
0 823 5 2 1 5490
0 824 7 1 2 803 5487
0 825 5 1 1 824
0 826 7 1 2 5468 5477
0 827 5 1 1 826
0 828 7 2 2 825 827
0 829 5 1 1 5494
0 830 7 1 2 5492 829
0 831 5 2 1 830
0 832 7 1 2 5469 5479
0 833 5 1 1 832
0 834 7 1 2 5481 833
0 835 5 1 1 834
0 836 7 3 2 5483 835
0 837 5 1 1 5498
0 838 7 1 2 5493 5499
0 839 5 1 1 838
0 840 7 1 2 5495 839
0 841 5 1 1 840
0 842 7 3 2 5496 841
0 843 5 1 1 5501
0 844 7 2 2 5497 837
0 845 5 1 1 5504
0 846 7 1 2 4772 845
0 847 5 2 1 846
0 848 7 1 2 4462 5505
0 849 5 1 1 848
0 850 7 2 2 5506 849
0 851 5 1 1 5508
0 852 7 2 2 4766 5509
0 853 5 2 1 5510
0 854 7 1 2 821 5507
0 855 5 1 1 854
0 856 7 1 2 5491 5500
0 857 5 1 1 856
0 858 7 2 2 855 857
0 859 5 1 1 5514
0 860 7 1 2 5512 859
0 861 5 2 1 860
0 862 7 2 2 843 5516
0 863 5 1 1 5518
0 864 7 1 2 4767 863
0 865 5 2 1 864
0 866 7 1 2 4455 5519
0 867 5 1 1 866
0 868 7 2 2 5520 867
0 869 5 1 1 5522
0 870 7 2 2 4760 5523
0 871 5 2 1 5524
0 872 7 1 2 851 5521
0 873 5 1 1 872
0 874 7 1 2 5502 5511
0 875 5 1 1 874
0 876 7 2 2 873 875
0 877 5 1 1 5528
0 878 7 1 2 5526 877
0 879 5 2 1 878
0 880 7 1 2 5503 5513
0 881 5 1 1 880
0 882 7 1 2 5515 881
0 883 5 1 1 882
0 884 7 3 2 5517 883
0 885 5 1 1 5532
0 886 7 1 2 5527 5533
0 887 5 1 1 886
0 888 7 1 2 5529 887
0 889 5 1 1 888
0 890 7 3 2 5530 889
0 891 5 1 1 5535
0 892 7 2 2 5531 885
0 893 5 1 1 5538
0 894 7 1 2 4761 893
0 895 5 2 1 894
0 896 7 1 2 4449 5539
0 897 5 1 1 896
0 898 7 2 2 5540 897
0 899 5 1 1 5542
0 900 7 2 2 4754 5543
0 901 5 2 1 5544
0 902 7 1 2 869 5541
0 903 5 1 1 902
0 904 7 1 2 5525 5534
0 905 5 1 1 904
0 906 7 2 2 903 905
0 907 5 1 1 5548
0 908 7 1 2 5546 907
0 909 5 2 1 908
0 910 7 2 2 891 5550
0 911 5 1 1 5552
0 912 7 1 2 4755 911
0 913 5 2 1 912
0 914 7 1 2 4442 5553
0 915 5 1 1 914
0 916 7 2 2 5554 915
0 917 5 1 1 5556
0 918 7 2 2 4749 5557
0 919 5 2 1 5558
0 920 7 1 2 899 5555
0 921 5 1 1 920
0 922 7 1 2 5536 5545
0 923 5 1 1 922
0 924 7 2 2 921 923
0 925 5 1 1 5562
0 926 7 1 2 5560 925
0 927 5 2 1 926
0 928 7 1 2 5537 5547
0 929 5 1 1 928
0 930 7 1 2 5549 929
0 931 5 1 1 930
0 932 7 3 2 5551 931
0 933 5 1 1 5566
0 934 7 1 2 5561 5567
0 935 5 1 1 934
0 936 7 1 2 5563 935
0 937 5 1 1 936
0 938 7 3 2 5564 937
0 939 5 1 1 5569
0 940 7 2 2 5565 933
0 941 5 1 1 5572
0 942 7 1 2 4750 941
0 943 5 2 1 942
0 944 7 1 2 4435 5573
0 945 5 1 1 944
0 946 7 2 2 5574 945
0 947 5 1 1 5576
0 948 7 2 2 4743 5577
0 949 5 2 1 5578
0 950 7 1 2 917 5575
0 951 5 1 1 950
0 952 7 1 2 5559 5568
0 953 5 1 1 952
0 954 7 2 2 951 953
0 955 5 1 1 5582
0 956 7 1 2 5580 955
0 957 5 2 1 956
0 958 7 2 2 939 5584
0 959 5 1 1 5586
0 960 7 1 2 4744 959
0 961 5 2 1 960
0 962 7 1 2 4429 5587
0 963 5 1 1 962
0 964 7 2 2 5588 963
0 965 5 1 1 5590
0 966 7 2 2 4737 5591
0 967 5 2 1 5592
0 968 7 1 2 947 5589
0 969 5 1 1 968
0 970 7 1 2 5570 5579
0 971 5 1 1 970
0 972 7 2 2 969 971
0 973 5 1 1 5596
0 974 7 1 2 5594 973
0 975 5 2 1 974
0 976 7 1 2 5571 5581
0 977 5 1 1 976
0 978 7 1 2 5583 977
0 979 5 1 1 978
0 980 7 3 2 5585 979
0 981 5 1 1 5600
0 982 7 1 2 5595 5601
0 983 5 1 1 982
0 984 7 1 2 5597 983
0 985 5 1 1 984
0 986 7 3 2 5598 985
0 987 5 1 1 5603
0 988 7 2 2 5599 981
0 989 5 1 1 5606
0 990 7 1 2 4738 989
0 991 5 2 1 990
0 992 7 1 2 4423 5607
0 993 5 1 1 992
0 994 7 2 2 5608 993
0 995 5 1 1 5610
0 996 7 2 2 4732 5611
0 997 5 2 1 5612
0 998 7 1 2 965 5609
0 999 5 1 1 998
0 1000 7 1 2 5593 5602
0 1001 5 1 1 1000
0 1002 7 2 2 999 1001
0 1003 5 1 1 5616
0 1004 7 1 2 5614 1003
0 1005 5 2 1 1004
0 1006 7 2 2 987 5618
0 1007 5 1 1 5620
0 1008 7 1 2 4733 1007
0 1009 5 2 1 1008
0 1010 7 1 2 4416 5621
0 1011 5 1 1 1010
0 1012 7 2 2 5622 1011
0 1013 5 1 1 5624
0 1014 7 2 2 4726 5625
0 1015 5 2 1 5626
0 1016 7 1 2 995 5623
0 1017 5 1 1 1016
0 1018 7 1 2 5604 5613
0 1019 5 1 1 1018
0 1020 7 2 2 1017 1019
0 1021 5 1 1 5630
0 1022 7 1 2 5628 1021
0 1023 5 2 1 1022
0 1024 7 1 2 5605 5615
0 1025 5 1 1 1024
0 1026 7 1 2 5617 1025
0 1027 5 1 1 1026
0 1028 7 3 2 5619 1027
0 1029 5 1 1 5634
0 1030 7 1 2 5629 5635
0 1031 5 1 1 1030
0 1032 7 1 2 5631 1031
0 1033 5 1 1 1032
0 1034 7 3 2 5632 1033
0 1035 5 1 1 5637
0 1036 7 2 2 5633 1029
0 1037 5 1 1 5640
0 1038 7 1 2 4727 1037
0 1039 5 2 1 1038
0 1040 7 1 2 4410 5641
0 1041 5 1 1 1040
0 1042 7 2 2 5642 1041
0 1043 5 1 1 5644
0 1044 7 2 2 4720 5645
0 1045 5 2 1 5646
0 1046 7 1 2 1013 5643
0 1047 5 1 1 1046
0 1048 7 1 2 5627 5636
0 1049 5 1 1 1048
0 1050 7 2 2 1047 1049
0 1051 5 1 1 5650
0 1052 7 1 2 5648 1051
0 1053 5 2 1 1052
0 1054 7 2 2 1035 5652
0 1055 5 1 1 5654
0 1056 7 1 2 4721 1055
0 1057 5 2 1 1056
0 1058 7 1 2 4403 5655
0 1059 5 1 1 1058
0 1060 7 2 2 5656 1059
0 1061 5 1 1 5658
0 1062 7 2 2 4715 5659
0 1063 5 2 1 5660
0 1064 7 1 2 1043 5657
0 1065 5 1 1 1064
0 1066 7 1 2 5638 5647
0 1067 5 1 1 1066
0 1068 7 2 2 1065 1067
0 1069 5 1 1 5664
0 1070 7 1 2 5662 1069
0 1071 5 2 1 1070
0 1072 7 1 2 5639 5649
0 1073 5 1 1 1072
0 1074 7 1 2 5651 1073
0 1075 5 1 1 1074
0 1076 7 3 2 5653 1075
0 1077 5 1 1 5668
0 1078 7 1 2 5663 5669
0 1079 5 1 1 1078
0 1080 7 1 2 5665 1079
0 1081 5 1 1 1080
0 1082 7 3 2 5666 1081
0 1083 5 1 1 5671
0 1084 7 2 2 5667 1077
0 1085 5 1 1 5674
0 1086 7 1 2 4716 1085
0 1087 5 2 1 1086
0 1088 7 1 2 4396 5675
0 1089 5 1 1 1088
0 1090 7 2 2 5676 1089
0 1091 5 1 1 5678
0 1092 7 2 2 4709 5679
0 1093 5 2 1 5680
0 1094 7 1 2 1061 5677
0 1095 5 1 1 1094
0 1096 7 1 2 5661 5670
0 1097 5 1 1 1096
0 1098 7 2 2 1095 1097
0 1099 5 1 1 5684
0 1100 7 1 2 5682 1099
0 1101 5 2 1 1100
0 1102 7 2 2 1083 5686
0 1103 5 1 1 5688
0 1104 7 1 2 4710 1103
0 1105 5 2 1 1104
0 1106 7 1 2 4390 5689
0 1107 5 1 1 1106
0 1108 7 2 2 5690 1107
0 1109 5 1 1 5692
0 1110 7 2 2 4703 5693
0 1111 5 2 1 5694
0 1112 7 1 2 1091 5691
0 1113 5 1 1 1112
0 1114 7 1 2 5672 5681
0 1115 5 1 1 1114
0 1116 7 2 2 1113 1115
0 1117 5 1 1 5698
0 1118 7 1 2 5696 1117
0 1119 5 2 1 1118
0 1120 7 1 2 5673 5683
0 1121 5 1 1 1120
0 1122 7 1 2 5685 1121
0 1123 5 1 1 1122
0 1124 7 3 2 5687 1123
0 1125 5 1 1 5702
0 1126 7 2 2 5700 1125
0 1127 5 1 1 5705
0 1128 7 1 2 4704 1127
0 1129 5 2 1 1128
0 1130 7 1 2 4384 5706
0 1131 5 1 1 1130
0 1132 7 3 2 5707 1131
0 1133 5 2 1 5709
0 1134 7 1 2 4697 5710
0 1135 5 2 1 1134
0 1136 7 1 2 1109 5708
0 1137 5 1 1 1136
0 1138 7 1 2 5695 5703
0 1139 5 1 1 1138
0 1140 7 2 2 1137 1139
0 1141 5 1 1 5716
0 1142 7 1 2 5714 1141
0 1143 5 2 1 1142
0 1144 7 1 2 5697 5704
0 1145 5 1 1 1144
0 1146 7 1 2 5699 1145
0 1147 5 1 1 1146
0 1148 7 2 2 5701 1147
0 1149 5 1 1 5720
0 1150 7 1 2 5715 5721
0 1151 5 1 1 1150
0 1152 7 1 2 5717 1151
0 1153 5 1 1 1152
0 1154 7 2 2 5718 1153
0 1155 5 1 1 5722
0 1156 7 2 2 5719 1149
0 1157 5 1 1 5724
0 1158 7 1 2 4378 5725
0 1159 5 2 1 1158
0 1160 7 2 2 5711 5726
0 1161 5 1 1 5728
0 1162 7 1 2 4698 1157
0 1163 5 3 1 1162
0 1164 7 1 2 5712 5730
0 1165 5 1 1 1164
0 1166 7 1 2 4686 4373
0 1167 7 1 2 1165 1166
0 1168 7 1 2 1161 1167
0 1169 5 1 1 1168
0 1170 7 2 2 4369 4691
0 1171 5 1 1 5733
0 1172 7 1 2 5731 5734
0 1173 7 1 2 5729 1172
0 1174 5 1 1 1173
0 1175 7 1 2 1169 1174
0 1176 5 1 1 1175
0 1177 7 1 2 1155 1176
0 1178 5 1 1 1177
0 1179 7 1 2 4370 5713
0 1180 5 1 1 1179
0 1181 7 1 2 4692 5723
0 1182 5 1 1 1181
0 1183 7 1 2 1180 1182
0 1184 5 1 1 1183
0 1185 7 1 2 5732 1171
0 1186 7 1 2 5727 1185
0 1187 7 1 2 1184 1186
0 1188 5 1 1 1187
0 1189 7 2 2 4668 110
0 1190 5 1 1 5735
0 1191 7 1 2 4962 5000
0 1192 5 1 1 1191
0 1193 7 2 2 1190 1192
0 1194 5 1 1 5737
0 1195 7 1 2 4660 5738
0 1196 5 2 1 1195
0 1197 7 1 2 5001 5736
0 1198 5 1 1 1197
0 1199 7 2 2 4983 1198
0 1200 5 1 1 5741
0 1201 7 1 2 5739 5742
0 1202 5 1 1 1201
0 1203 7 1 2 4661 1200
0 1204 5 2 1 1203
0 1205 7 2 2 1202 5743
0 1206 5 1 1 5745
0 1207 7 1 2 4950 5746
0 1208 5 1 1 1207
0 1209 7 1 2 4957 1194
0 1210 5 1 1 1209
0 1211 7 1 2 5740 1210
0 1212 7 2 2 5744 1211
0 1213 5 1 1 5747
0 1214 7 1 2 4652 5748
0 1215 5 2 1 1214
0 1216 7 1 2 4653 1206
0 1217 7 1 2 5749 1216
0 1218 5 2 1 1217
0 1219 7 3 2 1208 5751
0 1220 5 1 1 5753
0 1221 7 1 2 4645 1220
0 1222 5 1 1 1221
0 1223 7 1 2 4951 1213
0 1224 5 1 1 1223
0 1225 7 1 2 5750 1224
0 1226 7 1 2 5752 1225
0 1227 5 2 1 1226
0 1228 7 1 2 5754 5756
0 1229 5 1 1 1228
0 1230 7 1 2 4646 1229
0 1231 5 2 1 1230
0 1232 7 1 2 5755 5758
0 1233 5 1 1 1232
0 1234 7 2 2 1222 1233
0 1235 5 1 1 5760
0 1236 7 1 2 4939 5761
0 1237 5 1 1 1236
0 1238 7 1 2 4945 5757
0 1239 5 1 1 1238
0 1240 7 2 2 5759 1239
0 1241 5 1 1 5762
0 1242 7 1 2 4638 5763
0 1243 5 2 1 1242
0 1244 7 1 2 4639 1235
0 1245 7 1 2 5764 1244
0 1246 5 2 1 1245
0 1247 7 3 2 1237 5766
0 1248 5 1 1 5768
0 1249 7 1 2 4940 1241
0 1250 5 1 1 1249
0 1251 7 1 2 5765 1250
0 1252 7 1 2 5767 1251
0 1253 5 2 1 1252
0 1254 7 1 2 5769 5771
0 1255 5 1 1 1254
0 1256 7 1 2 4631 1255
0 1257 5 2 1 1256
0 1258 7 1 2 4934 5772
0 1259 5 1 1 1258
0 1260 7 2 2 5773 1259
0 1261 5 2 1 5775
0 1262 7 1 2 4632 1248
0 1263 5 1 1 1262
0 1264 7 1 2 5770 5774
0 1265 5 1 1 1264
0 1266 7 1 2 1263 1265
0 1267 5 2 1 1266
0 1268 7 1 2 5777 5779
0 1269 5 1 1 1268
0 1270 7 2 2 4625 1269
0 1271 5 1 1 5781
0 1272 7 1 2 5778 5782
0 1273 5 1 1 1272
0 1274 7 1 2 4928 5776
0 1275 5 1 1 1274
0 1276 7 2 2 1273 1275
0 1277 5 1 1 5783
0 1278 7 1 2 4929 5780
0 1279 5 1 1 1278
0 1280 7 2 2 1271 1279
0 1281 5 1 1 5785
0 1282 7 2 2 4619 1281
0 1283 5 1 1 5787
0 1284 7 1 2 5784 5788
0 1285 5 2 1 1284
0 1286 7 1 2 4922 5786
0 1287 5 1 1 1286
0 1288 7 2 2 1283 1287
0 1289 5 1 1 5791
0 1290 7 1 2 5789 1289
0 1291 5 1 1 1290
0 1292 7 1 2 4917 1291
0 1293 5 1 1 1292
0 1294 7 1 2 4923 1277
0 1295 5 2 1 1294
0 1296 7 1 2 5792 5793
0 1297 5 1 1 1296
0 1298 7 1 2 4612 1297
0 1299 5 2 1 1298
0 1300 7 2 2 1293 5795
0 1301 5 2 1 5797
0 1302 7 2 2 5790 5794
0 1303 5 1 1 5801
0 1304 7 1 2 4613 1303
0 1305 5 1 1 1304
0 1306 7 1 2 5796 5802
0 1307 5 1 1 1306
0 1308 7 1 2 1305 1307
0 1309 5 2 1 1308
0 1310 7 1 2 5799 5803
0 1311 5 1 1 1310
0 1312 7 2 2 4606 1311
0 1313 5 1 1 5805
0 1314 7 1 2 5800 5806
0 1315 5 1 1 1314
0 1316 7 1 2 4911 5798
0 1317 5 1 1 1316
0 1318 7 2 2 1315 1317
0 1319 5 1 1 5807
0 1320 7 1 2 4905 1319
0 1321 5 1 1 1320
0 1322 7 1 2 4912 5804
0 1323 5 1 1 1322
0 1324 7 2 2 1313 1323
0 1325 5 1 1 5809
0 1326 7 1 2 4599 5810
0 1327 5 2 1 1326
0 1328 7 1 2 4600 5808
0 1329 7 1 2 5811 1328
0 1330 5 2 1 1329
0 1331 7 3 2 1321 5813
0 1332 5 1 1 5815
0 1333 7 1 2 4906 1325
0 1334 5 1 1 1333
0 1335 7 1 2 5812 1334
0 1336 7 1 2 5814 1335
0 1337 5 2 1 1336
0 1338 7 1 2 5816 5818
0 1339 5 1 1 1338
0 1340 7 1 2 4592 1339
0 1341 5 2 1 1340
0 1342 7 1 2 4900 5819
0 1343 5 1 1 1342
0 1344 7 2 2 5820 1343
0 1345 5 2 1 5822
0 1346 7 1 2 4593 1332
0 1347 5 1 1 1346
0 1348 7 1 2 5817 5821
0 1349 5 1 1 1348
0 1350 7 1 2 1347 1349
0 1351 5 2 1 1350
0 1352 7 1 2 5824 5826
0 1353 5 1 1 1352
0 1354 7 2 2 4586 1353
0 1355 5 1 1 5828
0 1356 7 1 2 5825 5829
0 1357 5 1 1 1356
0 1358 7 1 2 4894 5823
0 1359 5 1 1 1358
0 1360 7 2 2 1357 1359
0 1361 5 1 1 5830
0 1362 7 1 2 4895 5827
0 1363 5 1 1 1362
0 1364 7 2 2 1355 1363
0 1365 5 1 1 5832
0 1366 7 2 2 4580 1365
0 1367 5 1 1 5834
0 1368 7 1 2 5831 5835
0 1369 5 2 1 1368
0 1370 7 1 2 4888 5833
0 1371 5 1 1 1370
0 1372 7 2 2 1367 1371
0 1373 5 1 1 5838
0 1374 7 1 2 5836 1373
0 1375 5 1 1 1374
0 1376 7 1 2 4883 1375
0 1377 5 1 1 1376
0 1378 7 1 2 4889 1361
0 1379 5 2 1 1378
0 1380 7 1 2 5839 5840
0 1381 5 1 1 1380
0 1382 7 1 2 4573 1381
0 1383 5 2 1 1382
0 1384 7 2 2 1377 5842
0 1385 5 2 1 5844
0 1386 7 2 2 5837 5841
0 1387 5 1 1 5848
0 1388 7 1 2 4574 1387
0 1389 5 1 1 1388
0 1390 7 1 2 5843 5849
0 1391 5 1 1 1390
0 1392 7 1 2 1389 1391
0 1393 5 2 1 1392
0 1394 7 1 2 5846 5850
0 1395 5 1 1 1394
0 1396 7 2 2 4567 1395
0 1397 5 1 1 5852
0 1398 7 1 2 5847 5853
0 1399 5 1 1 1398
0 1400 7 1 2 4876 5845
0 1401 5 1 1 1400
0 1402 7 2 2 1399 1401
0 1403 5 1 1 5854
0 1404 7 1 2 4869 1403
0 1405 5 1 1 1404
0 1406 7 1 2 4877 5851
0 1407 5 1 1 1406
0 1408 7 2 2 1397 1407
0 1409 5 1 1 5856
0 1410 7 1 2 4560 5857
0 1411 5 2 1 1410
0 1412 7 1 2 4561 5855
0 1413 7 1 2 5858 1412
0 1414 5 2 1 1413
0 1415 7 3 2 1405 5860
0 1416 5 1 1 5862
0 1417 7 1 2 4870 1409
0 1418 5 1 1 1417
0 1419 7 1 2 5859 1418
0 1420 7 1 2 5861 1419
0 1421 5 2 1 1420
0 1422 7 1 2 5863 5865
0 1423 5 1 1 1422
0 1424 7 1 2 4553 1423
0 1425 5 2 1 1424
0 1426 7 1 2 4863 5866
0 1427 5 1 1 1426
0 1428 7 2 2 5867 1427
0 1429 5 2 1 5869
0 1430 7 1 2 4554 1416
0 1431 5 1 1 1430
0 1432 7 1 2 5864 5868
0 1433 5 1 1 1432
0 1434 7 1 2 1431 1433
0 1435 5 2 1 1434
0 1436 7 1 2 5871 5873
0 1437 5 1 1 1436
0 1438 7 2 2 4547 1437
0 1439 5 1 1 5875
0 1440 7 1 2 5872 5876
0 1441 5 1 1 1440
0 1442 7 1 2 4856 5870
0 1443 5 1 1 1442
0 1444 7 2 2 1441 1443
0 1445 5 1 1 5877
0 1446 7 1 2 4857 5874
0 1447 5 1 1 1446
0 1448 7 2 2 1439 1447
0 1449 5 1 1 5879
0 1450 7 2 2 4541 1449
0 1451 5 1 1 5881
0 1452 7 1 2 5878 5882
0 1453 5 2 1 1452
0 1454 7 1 2 4849 5880
0 1455 5 1 1 1454
0 1456 7 2 2 1451 1455
0 1457 5 1 1 5885
0 1458 7 1 2 5883 1457
0 1459 5 1 1 1458
0 1460 7 1 2 4843 1459
0 1461 5 1 1 1460
0 1462 7 1 2 4850 1445
0 1463 5 2 1 1462
0 1464 7 1 2 5886 5887
0 1465 5 1 1 1464
0 1466 7 1 2 4534 1465
0 1467 5 2 1 1466
0 1468 7 2 2 1461 5889
0 1469 5 2 1 5891
0 1470 7 2 2 5884 5888
0 1471 5 1 1 5895
0 1472 7 1 2 4535 1471
0 1473 5 1 1 1472
0 1474 7 1 2 5890 5896
0 1475 5 1 1 1474
0 1476 7 1 2 1473 1475
0 1477 5 2 1 1476
0 1478 7 1 2 5893 5897
0 1479 5 1 1 1478
0 1480 7 2 2 4528 1479
0 1481 5 1 1 5899
0 1482 7 1 2 5894 5900
0 1483 5 1 1 1482
0 1484 7 1 2 4836 5892
0 1485 5 1 1 1484
0 1486 7 2 2 1483 1485
0 1487 5 1 1 5901
0 1488 7 1 2 4829 1487
0 1489 5 1 1 1488
0 1490 7 1 2 4837 5898
0 1491 5 1 1 1490
0 1492 7 2 2 1481 1491
0 1493 5 1 1 5903
0 1494 7 1 2 4521 5904
0 1495 5 2 1 1494
0 1496 7 1 2 4522 5902
0 1497 7 1 2 5905 1496
0 1498 5 2 1 1497
0 1499 7 3 2 1489 5907
0 1500 5 1 1 5909
0 1501 7 1 2 4830 1493
0 1502 5 1 1 1501
0 1503 7 1 2 5906 1502
0 1504 7 1 2 5908 1503
0 1505 5 2 1 1504
0 1506 7 1 2 5910 5912
0 1507 5 1 1 1506
0 1508 7 1 2 4514 1507
0 1509 5 2 1 1508
0 1510 7 1 2 4823 5913
0 1511 5 1 1 1510
0 1512 7 2 2 5914 1511
0 1513 5 2 1 5916
0 1514 7 1 2 4515 1500
0 1515 5 1 1 1514
0 1516 7 1 2 5911 5915
0 1517 5 1 1 1516
0 1518 7 1 2 1515 1517
0 1519 5 2 1 1518
0 1520 7 1 2 5918 5920
0 1521 5 1 1 1520
0 1522 7 2 2 4508 1521
0 1523 5 1 1 5922
0 1524 7 1 2 5919 5923
0 1525 5 1 1 1524
0 1526 7 1 2 4816 5917
0 1527 5 1 1 1526
0 1528 7 2 2 1525 1527
0 1529 5 1 1 5924
0 1530 7 1 2 4817 5921
0 1531 5 1 1 1530
0 1532 7 2 2 1523 1531
0 1533 5 1 1 5926
0 1534 7 2 2 4502 1533
0 1535 5 1 1 5928
0 1536 7 1 2 5925 5929
0 1537 5 2 1 1536
0 1538 7 1 2 4809 5927
0 1539 5 1 1 1538
0 1540 7 2 2 1535 1539
0 1541 5 1 1 5932
0 1542 7 1 2 5930 1541
0 1543 5 1 1 1542
0 1544 7 1 2 4803 1543
0 1545 5 1 1 1544
0 1546 7 1 2 4810 1529
0 1547 5 2 1 1546
0 1548 7 1 2 5933 5934
0 1549 5 1 1 1548
0 1550 7 1 2 4495 1549
0 1551 5 2 1 1550
0 1552 7 2 2 1545 5936
0 1553 5 2 1 5938
0 1554 7 2 2 5931 5935
0 1555 5 1 1 5942
0 1556 7 1 2 4496 1555
0 1557 5 1 1 1556
0 1558 7 1 2 5937 5943
0 1559 5 1 1 1558
0 1560 7 1 2 1557 1559
0 1561 5 2 1 1560
0 1562 7 1 2 5940 5944
0 1563 5 1 1 1562
0 1564 7 2 2 4489 1563
0 1565 5 1 1 5946
0 1566 7 1 2 5941 5947
0 1567 5 1 1 1566
0 1568 7 1 2 4796 5939
0 1569 5 1 1 1568
0 1570 7 2 2 1567 1569
0 1571 5 1 1 5948
0 1572 7 1 2 4790 1571
0 1573 5 1 1 1572
0 1574 7 1 2 4797 5945
0 1575 5 1 1 1574
0 1576 7 2 2 1565 1575
0 1577 5 1 1 5950
0 1578 7 1 2 4482 5951
0 1579 5 2 1 1578
0 1580 7 1 2 4483 5949
0 1581 7 1 2 5952 1580
0 1582 5 2 1 1581
0 1583 7 3 2 1573 5954
0 1584 5 1 1 5956
0 1585 7 1 2 4791 1577
0 1586 5 1 1 1585
0 1587 7 1 2 5953 1586
0 1588 7 1 2 5955 1587
0 1589 5 2 1 1588
0 1590 7 1 2 5957 5959
0 1591 5 1 1 1590
0 1592 7 1 2 4475 1591
0 1593 5 2 1 1592
0 1594 7 1 2 4785 5960
0 1595 5 1 1 1594
0 1596 7 2 2 5961 1595
0 1597 5 2 1 5963
0 1598 7 1 2 4476 1584
0 1599 5 1 1 1598
0 1600 7 1 2 5958 5962
0 1601 5 1 1 1600
0 1602 7 1 2 1599 1601
0 1603 5 2 1 1602
0 1604 7 1 2 5965 5967
0 1605 5 1 1 1604
0 1606 7 2 2 4469 1605
0 1607 5 1 1 5969
0 1608 7 1 2 5966 5970
0 1609 5 1 1 1608
0 1610 7 1 2 4779 5964
0 1611 5 1 1 1610
0 1612 7 2 2 1609 1611
0 1613 5 1 1 5971
0 1614 7 1 2 4780 5968
0 1615 5 1 1 1614
0 1616 7 2 2 1607 1615
0 1617 5 1 1 5973
0 1618 7 2 2 4463 1617
0 1619 5 1 1 5975
0 1620 7 1 2 5972 5976
0 1621 5 2 1 1620
0 1622 7 1 2 4773 5974
0 1623 5 1 1 1622
0 1624 7 2 2 1619 1623
0 1625 5 1 1 5979
0 1626 7 1 2 5977 1625
0 1627 5 1 1 1626
0 1628 7 1 2 4768 1627
0 1629 5 1 1 1628
0 1630 7 1 2 4774 1613
0 1631 5 2 1 1630
0 1632 7 1 2 5980 5981
0 1633 5 1 1 1632
0 1634 7 1 2 4456 1633
0 1635 5 2 1 1634
0 1636 7 2 2 1629 5983
0 1637 5 2 1 5985
0 1638 7 2 2 5978 5982
0 1639 5 1 1 5989
0 1640 7 1 2 4457 1639
0 1641 5 1 1 1640
0 1642 7 1 2 5984 5990
0 1643 5 1 1 1642
0 1644 7 1 2 1641 1643
0 1645 5 2 1 1644
0 1646 7 1 2 5987 5991
0 1647 5 1 1 1646
0 1648 7 2 2 4450 1647
0 1649 5 1 1 5993
0 1650 7 1 2 5988 5994
0 1651 5 1 1 1650
0 1652 7 1 2 4762 5986
0 1653 5 1 1 1652
0 1654 7 2 2 1651 1653
0 1655 5 1 1 5995
0 1656 7 1 2 4756 1655
0 1657 5 1 1 1656
0 1658 7 1 2 4763 5992
0 1659 5 1 1 1658
0 1660 7 2 2 1649 1659
0 1661 5 1 1 5997
0 1662 7 1 2 4443 5998
0 1663 5 2 1 1662
0 1664 7 1 2 4444 5996
0 1665 7 1 2 5999 1664
0 1666 5 2 1 1665
0 1667 7 3 2 1657 6001
0 1668 5 1 1 6003
0 1669 7 1 2 4757 1661
0 1670 5 1 1 1669
0 1671 7 1 2 6000 1670
0 1672 7 1 2 6002 1671
0 1673 5 2 1 1672
0 1674 7 1 2 6004 6006
0 1675 5 1 1 1674
0 1676 7 1 2 4436 1675
0 1677 5 2 1 1676
0 1678 7 1 2 4751 6007
0 1679 5 1 1 1678
0 1680 7 2 2 6008 1679
0 1681 5 2 1 6010
0 1682 7 1 2 4437 1668
0 1683 5 1 1 1682
0 1684 7 1 2 6005 6009
0 1685 5 1 1 1684
0 1686 7 1 2 1683 1685
0 1687 5 2 1 1686
0 1688 7 1 2 6012 6014
0 1689 5 1 1 1688
0 1690 7 2 2 4430 1689
0 1691 5 1 1 6016
0 1692 7 1 2 6013 6017
0 1693 5 1 1 1692
0 1694 7 1 2 4745 6011
0 1695 5 1 1 1694
0 1696 7 2 2 1693 1695
0 1697 5 1 1 6018
0 1698 7 1 2 4746 6015
0 1699 5 1 1 1698
0 1700 7 2 2 1691 1699
0 1701 5 1 1 6020
0 1702 7 2 2 4424 1701
0 1703 5 1 1 6022
0 1704 7 1 2 6019 6023
0 1705 5 2 1 1704
0 1706 7 1 2 4739 6021
0 1707 5 1 1 1706
0 1708 7 2 2 1703 1707
0 1709 5 1 1 6026
0 1710 7 1 2 6024 1709
0 1711 5 1 1 1710
0 1712 7 1 2 4734 1711
0 1713 5 1 1 1712
0 1714 7 1 2 4740 1697
0 1715 5 2 1 1714
0 1716 7 1 2 6027 6028
0 1717 5 1 1 1716
0 1718 7 1 2 4417 1717
0 1719 5 2 1 1718
0 1720 7 2 2 1713 6030
0 1721 5 2 1 6032
0 1722 7 2 2 6025 6029
0 1723 5 1 1 6036
0 1724 7 1 2 4418 1723
0 1725 5 1 1 1724
0 1726 7 1 2 6031 6037
0 1727 5 1 1 1726
0 1728 7 1 2 1725 1727
0 1729 5 2 1 1728
0 1730 7 1 2 6034 6038
0 1731 5 1 1 1730
0 1732 7 2 2 4411 1731
0 1733 5 1 1 6040
0 1734 7 1 2 6035 6041
0 1735 5 1 1 1734
0 1736 7 1 2 4728 6033
0 1737 5 1 1 1736
0 1738 7 2 2 1735 1737
0 1739 5 1 1 6042
0 1740 7 1 2 4722 1739
0 1741 5 1 1 1740
0 1742 7 1 2 4729 6039
0 1743 5 1 1 1742
0 1744 7 2 2 1733 1743
0 1745 5 1 1 6044
0 1746 7 1 2 4404 6045
0 1747 5 2 1 1746
0 1748 7 1 2 4405 6043
0 1749 7 1 2 6046 1748
0 1750 5 2 1 1749
0 1751 7 3 2 1741 6048
0 1752 5 1 1 6050
0 1753 7 1 2 4397 1752
0 1754 5 1 1 1753
0 1755 7 1 2 4723 1745
0 1756 5 1 1 1755
0 1757 7 1 2 6047 1756
0 1758 7 1 2 6049 1757
0 1759 5 2 1 1758
0 1760 7 1 2 6051 6053
0 1761 5 1 1 1760
0 1762 7 1 2 4398 1761
0 1763 5 2 1 1762
0 1764 7 1 2 6052 6055
0 1765 5 1 1 1764
0 1766 7 1 2 1754 1765
0 1767 5 2 1 1766
0 1768 7 1 2 4711 6057
0 1769 5 1 1 1768
0 1770 7 1 2 4717 6054
0 1771 5 1 1 1770
0 1772 7 2 2 6056 1771
0 1773 5 2 1 6059
0 1774 7 1 2 6058 6061
0 1775 5 1 1 1774
0 1776 7 2 2 4391 1775
0 1777 5 1 1 6063
0 1778 7 2 2 1769 1777
0 1779 5 2 1 6065
0 1780 7 1 2 6062 6064
0 1781 5 1 1 1780
0 1782 7 1 2 4712 6060
0 1783 5 1 1 1782
0 1784 7 2 2 1781 1783
0 1785 7 1 2 6067 6069
0 1786 5 1 1 1785
0 1787 7 2 2 4385 1786
0 1788 5 1 1 6071
0 1789 7 1 2 6068 6072
0 1790 5 1 1 1789
0 1791 7 1 2 4705 6066
0 1792 5 1 1 1791
0 1793 7 2 2 1790 1792
0 1794 7 1 2 4699 6073
0 1795 5 1 1 1794
0 1796 7 1 2 4706 6070
0 1797 5 1 1 1796
0 1798 7 2 2 1788 1797
0 1799 5 2 1 6075
0 1800 7 1 2 6074 6077
0 1801 5 1 1 1800
0 1802 7 2 2 4379 1801
0 1803 5 1 1 6079
0 1804 7 2 2 1795 1803
0 1805 5 1 1 6081
0 1806 7 1 2 6078 6080
0 1807 5 1 1 1806
0 1808 7 1 2 4700 6076
0 1809 5 1 1 1808
0 1810 7 1 2 4693 1809
0 1811 7 1 2 1807 1810
0 1812 5 1 1 1811
0 1813 7 1 2 1805 1812
0 1814 5 1 1 1813
0 1815 7 1 2 4694 6082
0 1816 5 1 1 1815
0 1817 7 1 2 4687 1816
0 1818 7 1 2 1814 1817
0 1819 5 1 1 1818
0 1820 7 2 2 4669 4678
0 1821 5 1 1 6083
0 1822 7 1 2 4683 1821
0 1823 5 2 1 1822
0 1824 7 1 2 4958 6085
0 1825 5 1 1 1824
0 1826 7 1 2 135 6086
0 1827 5 1 1 1826
0 1828 7 1 2 4662 1827
0 1829 5 3 1 1828
0 1830 7 5 2 1825 6087
0 1831 5 1 1 6090
0 1832 7 2 2 4684 6084
0 1833 5 2 1 6095
0 1834 7 2 2 4663 4670
0 1835 5 1 1 6099
0 1836 7 1 2 4966 1835
0 1837 5 1 1 1836
0 1838 7 1 2 4970 6100
0 1839 5 1 1 1838
0 1840 7 1 2 1837 1839
0 1841 7 2 2 6097 1840
0 1842 5 2 1 6101
0 1843 7 1 2 4952 6103
0 1844 5 1 1 1843
0 1845 7 1 2 4963 6098
0 1846 5 1 1 1845
0 1847 7 1 2 4671 6096
0 1848 5 1 1 1847
0 1849 7 3 2 1846 1848
0 1850 5 1 1 6105
0 1851 7 1 2 6091 6106
0 1852 5 1 1 1851
0 1853 7 1 2 6104 1852
0 1854 5 1 1 1853
0 1855 7 2 2 4654 1854
0 1856 5 2 1 6108
0 1857 7 2 2 1844 6110
0 1858 5 1 1 6112
0 1859 7 2 2 4647 6113
0 1860 7 1 2 6092 6114
0 1861 5 2 1 1860
0 1862 7 2 2 4655 6093
0 1863 5 1 1 6118
0 1864 7 1 2 6102 6119
0 1865 5 1 1 1864
0 1866 7 1 2 6088 1865
0 1867 5 1 1 1866
0 1868 7 1 2 1850 1867
0 1869 5 1 1 1868
0 1870 7 1 2 6089 6107
0 1871 7 1 2 1863 1870
0 1872 5 1 1 1871
0 1873 7 2 2 1869 1872
0 1874 7 1 2 6116 6120
0 1875 5 2 1 1874
0 1876 7 1 2 4648 6122
0 1877 5 2 1 1876
0 1878 7 1 2 4946 6121
0 1879 5 1 1 1878
0 1880 7 4 2 6124 1879
0 1881 5 1 1 6126
0 1882 7 1 2 1858 6125
0 1883 5 1 1 1882
0 1884 7 1 2 6115 6123
0 1885 5 2 1 1884
0 1886 7 2 2 1883 6130
0 1887 5 1 1 6132
0 1888 7 1 2 4640 6127
0 1889 7 1 2 6133 1888
0 1890 5 2 1 1889
0 1891 7 1 2 6094 6111
0 1892 5 1 1 1891
0 1893 7 1 2 1831 6109
0 1894 5 1 1 1893
0 1895 7 1 2 1892 1894
0 1896 7 1 2 6131 1895
0 1897 5 1 1 1896
0 1898 7 1 2 6117 1897
0 1899 5 2 1 1898
0 1900 7 1 2 6134 6136
0 1901 5 1 1 1900
0 1902 7 2 2 4641 1901
0 1903 5 2 1 6138
0 1904 7 1 2 4941 6137
0 1905 5 1 1 1904
0 1906 7 3 2 6140 1905
0 1907 5 1 1 6142
0 1908 7 2 2 4633 6143
0 1909 7 1 2 6128 6145
0 1910 5 2 1 1909
0 1911 7 1 2 6129 6139
0 1912 5 2 1 1911
0 1913 7 1 2 1881 6141
0 1914 5 1 1 1913
0 1915 7 1 2 6149 1914
0 1916 5 1 1 1915
0 1917 7 1 2 1887 6150
0 1918 5 1 1 1917
0 1919 7 2 2 6135 1918
0 1920 5 2 1 6151
0 1921 7 1 2 6146 6152
0 1922 5 1 1 1921
0 1923 7 1 2 1916 1922
0 1924 5 1 1 1923
0 1925 7 1 2 6147 1924
0 1926 5 2 1 1925
0 1927 7 1 2 6148 6153
0 1928 5 1 1 1927
0 1929 7 2 2 4634 1928
0 1930 5 2 1 6157
0 1931 7 1 2 6144 6159
0 1932 5 1 1 1931
0 1933 7 1 2 1907 6158
0 1934 5 1 1 1933
0 1935 7 2 2 1932 1934
0 1936 5 1 1 6161
0 1937 7 1 2 4935 6154
0 1938 5 1 1 1937
0 1939 7 4 2 6160 1938
0 1940 5 1 1 6163
0 1941 7 1 2 4626 6164
0 1942 7 1 2 1936 1941
0 1943 5 2 1 1942
0 1944 7 1 2 6155 6167
0 1945 5 1 1 1944
0 1946 7 2 2 4627 1945
0 1947 5 2 1 6169
0 1948 7 1 2 4930 6156
0 1949 5 1 1 1948
0 1950 7 3 2 6171 1949
0 1951 5 1 1 6173
0 1952 7 1 2 6165 6170
0 1953 5 2 1 1952
0 1954 7 1 2 6162 6176
0 1955 5 1 1 1954
0 1956 7 1 2 6168 1955
0 1957 5 2 1 1956
0 1958 7 2 2 4620 6174
0 1959 7 1 2 6166 6180
0 1960 5 2 1 1959
0 1961 7 1 2 6178 6182
0 1962 5 2 1 1961
0 1963 7 1 2 4621 6184
0 1964 5 2 1 1963
0 1965 7 1 2 4924 6179
0 1966 5 1 1 1965
0 1967 7 4 2 6186 1966
0 1968 5 1 1 6188
0 1969 7 2 2 4614 6189
0 1970 7 1 2 6175 6192
0 1971 5 2 1 1970
0 1972 7 1 2 1951 6187
0 1973 5 1 1 1972
0 1974 7 1 2 6181 6185
0 1975 5 2 1 1974
0 1976 7 1 2 1973 6196
0 1977 5 1 1 1976
0 1978 7 1 2 1940 6172
0 1979 5 1 1 1978
0 1980 7 1 2 6177 1979
0 1981 5 1 1 1980
0 1982 7 1 2 6197 1981
0 1983 5 1 1 1982
0 1984 7 2 2 6183 1983
0 1985 5 2 1 6198
0 1986 7 1 2 6193 6199
0 1987 5 1 1 1986
0 1988 7 1 2 1977 1987
0 1989 5 1 1 1988
0 1990 7 1 2 6194 1989
0 1991 5 2 1 1990
0 1992 7 1 2 6195 6200
0 1993 5 1 1 1992
0 1994 7 2 2 4615 1993
0 1995 5 2 1 6204
0 1996 7 1 2 4918 6201
0 1997 5 1 1 1996
0 1998 7 2 2 6206 1997
0 1999 5 1 1 6208
0 2000 7 2 2 4607 6209
0 2001 7 1 2 6190 6210
0 2002 5 2 1 2001
0 2003 7 1 2 6202 6212
0 2004 5 2 1 2003
0 2005 7 1 2 4608 6214
0 2006 5 2 1 2005
0 2007 7 1 2 4913 6203
0 2008 5 1 1 2007
0 2009 7 4 2 6216 2008
0 2010 5 1 1 6218
0 2011 7 1 2 1999 6217
0 2012 5 1 1 2011
0 2013 7 1 2 6211 6215
0 2014 5 2 1 2013
0 2015 7 2 2 2012 6222
0 2016 5 1 1 6224
0 2017 7 1 2 4601 6219
0 2018 7 1 2 6225 2017
0 2019 5 2 1 2018
0 2020 7 1 2 6191 6207
0 2021 5 1 1 2020
0 2022 7 1 2 1968 6205
0 2023 5 1 1 2022
0 2024 7 1 2 2021 2023
0 2025 7 1 2 6223 2024
0 2026 5 1 1 2025
0 2027 7 1 2 6213 2026
0 2028 5 2 1 2027
0 2029 7 1 2 6226 6228
0 2030 5 1 1 2029
0 2031 7 2 2 4602 2030
0 2032 5 2 1 6230
0 2033 7 1 2 4907 6229
0 2034 5 1 1 2033
0 2035 7 3 2 6232 2034
0 2036 5 1 1 6234
0 2037 7 2 2 4594 6235
0 2038 7 1 2 6220 6237
0 2039 5 2 1 2038
0 2040 7 1 2 6221 6231
0 2041 5 2 1 2040
0 2042 7 1 2 2010 6233
0 2043 5 1 1 2042
0 2044 7 1 2 6241 2043
0 2045 5 1 1 2044
0 2046 7 1 2 2016 6242
0 2047 5 1 1 2046
0 2048 7 2 2 6227 2047
0 2049 5 2 1 6243
0 2050 7 1 2 6238 6244
0 2051 5 1 1 2050
0 2052 7 1 2 2045 2051
0 2053 5 1 1 2052
0 2054 7 1 2 6239 2053
0 2055 5 2 1 2054
0 2056 7 1 2 6240 6245
0 2057 5 1 1 2056
0 2058 7 2 2 4595 2057
0 2059 5 2 1 6249
0 2060 7 1 2 6236 6251
0 2061 5 1 1 2060
0 2062 7 1 2 2036 6250
0 2063 5 1 1 2062
0 2064 7 2 2 2061 2063
0 2065 5 1 1 6253
0 2066 7 1 2 4901 6246
0 2067 5 1 1 2066
0 2068 7 4 2 6252 2067
0 2069 5 1 1 6255
0 2070 7 1 2 4587 6256
0 2071 7 1 2 2065 2070
0 2072 5 2 1 2071
0 2073 7 1 2 6247 6259
0 2074 5 1 1 2073
0 2075 7 2 2 4588 2074
0 2076 5 2 1 6261
0 2077 7 1 2 4896 6248
0 2078 5 1 1 2077
0 2079 7 3 2 6263 2078
0 2080 5 1 1 6265
0 2081 7 1 2 6257 6262
0 2082 5 2 1 2081
0 2083 7 1 2 6254 6268
0 2084 5 1 1 2083
0 2085 7 1 2 6260 2084
0 2086 5 2 1 2085
0 2087 7 2 2 4581 6266
0 2088 7 1 2 6258 6272
0 2089 5 2 1 2088
0 2090 7 1 2 6270 6274
0 2091 5 2 1 2090
0 2092 7 1 2 4582 6276
0 2093 5 2 1 2092
0 2094 7 1 2 4890 6271
0 2095 5 1 1 2094
0 2096 7 4 2 6278 2095
0 2097 5 1 1 6280
0 2098 7 2 2 4575 6281
0 2099 7 1 2 6267 6284
0 2100 5 2 1 2099
0 2101 7 1 2 2080 6279
0 2102 5 1 1 2101
0 2103 7 1 2 6273 6277
0 2104 5 2 1 2103
0 2105 7 1 2 2102 6288
0 2106 5 1 1 2105
0 2107 7 1 2 2069 6264
0 2108 5 1 1 2107
0 2109 7 1 2 6269 2108
0 2110 5 1 1 2109
0 2111 7 1 2 6289 2110
0 2112 5 1 1 2111
0 2113 7 2 2 6275 2112
0 2114 5 2 1 6290
0 2115 7 1 2 6285 6291
0 2116 5 1 1 2115
0 2117 7 1 2 2106 2116
0 2118 5 1 1 2117
0 2119 7 1 2 6286 2118
0 2120 5 2 1 2119
0 2121 7 1 2 6287 6292
0 2122 5 1 1 2121
0 2123 7 2 2 4576 2122
0 2124 5 2 1 6296
0 2125 7 1 2 4884 6293
0 2126 5 1 1 2125
0 2127 7 4 2 6298 2126
0 2128 5 1 1 6300
0 2129 7 1 2 4568 6282
0 2130 7 1 2 6301 2129
0 2131 5 2 1 2130
0 2132 7 1 2 6294 6304
0 2133 5 1 1 2132
0 2134 7 2 2 4569 2133
0 2135 5 2 1 6306
0 2136 7 1 2 4878 6295
0 2137 5 1 1 2136
0 2138 7 4 2 6308 2137
0 2139 5 1 1 6310
0 2140 7 1 2 4562 6302
0 2141 7 1 2 6311 2140
0 2142 5 2 1 2141
0 2143 7 1 2 6303 6307
0 2144 5 2 1 2143
0 2145 7 1 2 6283 6299
0 2146 5 1 1 2145
0 2147 7 1 2 2097 6297
0 2148 5 1 1 2147
0 2149 7 1 2 2146 2148
0 2150 7 1 2 6316 2149
0 2151 5 1 1 2150
0 2152 7 1 2 6305 2151
0 2153 5 2 1 2152
0 2154 7 1 2 6314 6318
0 2155 5 1 1 2154
0 2156 7 2 2 4563 2155
0 2157 5 2 1 6320
0 2158 7 1 2 4871 6319
0 2159 5 1 1 2158
0 2160 7 4 2 6322 2159
0 2161 5 1 1 6324
0 2162 7 2 2 4555 6325
0 2163 7 1 2 6312 6328
0 2164 5 2 1 2163
0 2165 7 1 2 2139 6323
0 2166 5 1 1 2165
0 2167 7 1 2 6313 6321
0 2168 5 2 1 2167
0 2169 7 1 2 2166 6332
0 2170 5 1 1 2169
0 2171 7 1 2 2128 6309
0 2172 5 1 1 2171
0 2173 7 1 2 6317 2172
0 2174 5 1 1 2173
0 2175 7 1 2 6333 2174
0 2176 5 1 1 2175
0 2177 7 2 2 6315 2176
0 2178 5 2 1 6334
0 2179 7 1 2 6329 6335
0 2180 5 1 1 2179
0 2181 7 1 2 2170 2180
0 2182 5 1 1 2181
0 2183 7 1 2 6330 2182
0 2184 5 2 1 2183
0 2185 7 1 2 6331 6336
0 2186 5 1 1 2185
0 2187 7 2 2 4556 2186
0 2188 5 2 1 6340
0 2189 7 1 2 4864 6337
0 2190 5 1 1 2189
0 2191 7 3 2 6342 2190
0 2192 5 1 1 6344
0 2193 7 2 2 4548 6345
0 2194 7 1 2 6326 6347
0 2195 5 2 1 2194
0 2196 7 1 2 6338 6349
0 2197 5 2 1 2196
0 2198 7 1 2 4549 6351
0 2199 5 2 1 2198
0 2200 7 1 2 4858 6339
0 2201 5 1 1 2200
0 2202 7 4 2 6353 2201
0 2203 5 1 1 6355
0 2204 7 1 2 4542 6346
0 2205 7 1 2 6356 2204
0 2206 5 2 1 2205
0 2207 7 1 2 6348 6352
0 2208 5 2 1 2207
0 2209 7 1 2 6327 6343
0 2210 5 1 1 2209
0 2211 7 1 2 2161 6341
0 2212 5 1 1 2211
0 2213 7 1 2 2210 2212
0 2214 7 1 2 6361 2213
0 2215 5 1 1 2214
0 2216 7 1 2 6350 2215
0 2217 5 2 1 2216
0 2218 7 1 2 6359 6363
0 2219 5 1 1 2218
0 2220 7 2 2 4543 2219
0 2221 5 2 1 6365
0 2222 7 1 2 4851 6364
0 2223 5 1 1 2222
0 2224 7 4 2 6367 2223
0 2225 5 1 1 6369
0 2226 7 2 2 4536 6370
0 2227 7 1 2 6357 6373
0 2228 5 2 1 2227
0 2229 7 1 2 2203 6368
0 2230 5 1 1 2229
0 2231 7 1 2 6358 6366
0 2232 5 2 1 2231
0 2233 7 1 2 2230 6377
0 2234 5 1 1 2233
0 2235 7 1 2 2192 6354
0 2236 5 1 1 2235
0 2237 7 1 2 6362 2236
0 2238 5 1 1 2237
0 2239 7 1 2 6378 2238
0 2240 5 1 1 2239
0 2241 7 2 2 6360 2240
0 2242 5 2 1 6379
0 2243 7 1 2 6374 6380
0 2244 5 1 1 2243
0 2245 7 1 2 2234 2244
0 2246 5 1 1 2245
0 2247 7 1 2 6375 2246
0 2248 5 2 1 2247
0 2249 7 1 2 6376 6381
0 2250 5 1 1 2249
0 2251 7 2 2 4537 2250
0 2252 5 2 1 6385
0 2253 7 1 2 4844 6382
0 2254 5 1 1 2253
0 2255 7 4 2 6387 2254
0 2256 5 1 1 6389
0 2257 7 1 2 4529 6371
0 2258 7 1 2 6390 2257
0 2259 5 2 1 2258
0 2260 7 1 2 6383 6393
0 2261 5 1 1 2260
0 2262 7 2 2 4530 2261
0 2263 5 2 1 6395
0 2264 7 1 2 4838 6384
0 2265 5 1 1 2264
0 2266 7 4 2 6397 2265
0 2267 5 1 1 6399
0 2268 7 1 2 4523 6391
0 2269 7 1 2 6400 2268
0 2270 5 2 1 2269
0 2271 7 1 2 6392 6396
0 2272 5 2 1 2271
0 2273 7 1 2 6372 6388
0 2274 5 1 1 2273
0 2275 7 1 2 2225 6386
0 2276 5 1 1 2275
0 2277 7 1 2 2274 2276
0 2278 7 1 2 6405 2277
0 2279 5 1 1 2278
0 2280 7 1 2 6394 2279
0 2281 5 2 1 2280
0 2282 7 1 2 6403 6407
0 2283 5 1 1 2282
0 2284 7 2 2 4524 2283
0 2285 5 2 1 6409
0 2286 7 1 2 4831 6408
0 2287 5 1 1 2286
0 2288 7 4 2 6411 2287
0 2289 5 1 1 6413
0 2290 7 2 2 4516 6414
0 2291 7 1 2 6401 6417
0 2292 5 2 1 2291
0 2293 7 1 2 2267 6412
0 2294 5 1 1 2293
0 2295 7 1 2 6402 6410
0 2296 5 2 1 2295
0 2297 7 1 2 2294 6421
0 2298 5 1 1 2297
0 2299 7 1 2 2256 6398
0 2300 5 1 1 2299
0 2301 7 1 2 6406 2300
0 2302 5 1 1 2301
0 2303 7 1 2 6422 2302
0 2304 5 1 1 2303
0 2305 7 2 2 6404 2304
0 2306 5 2 1 6423
0 2307 7 1 2 6418 6424
0 2308 5 1 1 2307
0 2309 7 1 2 2298 2308
0 2310 5 1 1 2309
0 2311 7 1 2 6419 2310
0 2312 5 2 1 2311
0 2313 7 1 2 6420 6425
0 2314 5 1 1 2313
0 2315 7 2 2 4517 2314
0 2316 5 2 1 6429
0 2317 7 1 2 4824 6426
0 2318 5 1 1 2317
0 2319 7 4 2 6431 2318
0 2320 5 1 1 6433
0 2321 7 1 2 4509 6415
0 2322 7 1 2 6434 2321
0 2323 5 2 1 2322
0 2324 7 1 2 6427 6437
0 2325 5 1 1 2324
0 2326 7 2 2 4510 2325
0 2327 5 2 1 6439
0 2328 7 1 2 4818 6428
0 2329 5 1 1 2328
0 2330 7 3 2 6441 2329
0 2331 5 1 1 6443
0 2332 7 2 2 4503 6444
0 2333 7 1 2 6435 6446
0 2334 5 2 1 2333
0 2335 7 1 2 6436 6440
0 2336 5 2 1 2335
0 2337 7 1 2 6416 6432
0 2338 5 1 1 2337
0 2339 7 1 2 2289 6430
0 2340 5 1 1 2339
0 2341 7 1 2 2338 2340
0 2342 7 1 2 6450 2341
0 2343 5 1 1 2342
0 2344 7 1 2 6438 2343
0 2345 5 2 1 2344
0 2346 7 1 2 6448 6452
0 2347 5 2 1 2346
0 2348 7 1 2 4504 6454
0 2349 5 2 1 2348
0 2350 7 1 2 4811 6453
0 2351 5 1 1 2350
0 2352 7 4 2 6456 2351
0 2353 5 1 1 6458
0 2354 7 2 2 4497 6459
0 2355 7 1 2 6445 6462
0 2356 5 2 1 2355
0 2357 7 1 2 2331 6457
0 2358 5 1 1 2357
0 2359 7 1 2 6447 6455
0 2360 5 2 1 2359
0 2361 7 1 2 2358 6466
0 2362 5 1 1 2361
0 2363 7 1 2 2320 6442
0 2364 5 1 1 2363
0 2365 7 1 2 6451 2364
0 2366 5 1 1 2365
0 2367 7 1 2 6467 2366
0 2368 5 1 1 2367
0 2369 7 2 2 6449 2368
0 2370 5 2 1 6468
0 2371 7 1 2 6463 6469
0 2372 5 1 1 2371
0 2373 7 1 2 2362 2372
0 2374 5 1 1 2373
0 2375 7 1 2 6464 2374
0 2376 5 2 1 2375
0 2377 7 1 2 6465 6470
0 2378 5 1 1 2377
0 2379 7 2 2 4498 2378
0 2380 5 2 1 6474
0 2381 7 1 2 4804 6471
0 2382 5 1 1 2381
0 2383 7 4 2 6476 2382
0 2384 5 1 1 6478
0 2385 7 1 2 4490 6460
0 2386 7 1 2 6479 2385
0 2387 5 2 1 2386
0 2388 7 1 2 6472 6482
0 2389 5 1 1 2388
0 2390 7 2 2 4491 2389
0 2391 5 2 1 6484
0 2392 7 1 2 4798 6473
0 2393 5 1 1 2392
0 2394 7 4 2 6486 2393
0 2395 5 1 1 6488
0 2396 7 1 2 4484 6480
0 2397 7 1 2 6489 2396
0 2398 5 2 1 2397
0 2399 7 1 2 6481 6485
0 2400 5 2 1 2399
0 2401 7 1 2 6461 6477
0 2402 5 1 1 2401
0 2403 7 1 2 2353 6475
0 2404 5 1 1 2403
0 2405 7 1 2 2402 2404
0 2406 7 1 2 6494 2405
0 2407 5 1 1 2406
0 2408 7 1 2 6483 2407
0 2409 5 2 1 2408
0 2410 7 1 2 6492 6496
0 2411 5 1 1 2410
0 2412 7 2 2 4485 2411
0 2413 5 2 1 6498
0 2414 7 1 2 4792 6497
0 2415 5 1 1 2414
0 2416 7 4 2 6500 2415
0 2417 5 1 1 6502
0 2418 7 2 2 4477 6503
0 2419 7 1 2 6490 6506
0 2420 5 2 1 2419
0 2421 7 1 2 2395 6501
0 2422 5 1 1 2421
0 2423 7 1 2 6491 6499
0 2424 5 2 1 2423
0 2425 7 1 2 2422 6510
0 2426 5 1 1 2425
0 2427 7 1 2 2384 6487
0 2428 5 1 1 2427
0 2429 7 1 2 6495 2428
0 2430 5 1 1 2429
0 2431 7 1 2 6511 2430
0 2432 5 1 1 2431
0 2433 7 2 2 6493 2432
0 2434 5 2 1 6512
0 2435 7 1 2 6507 6513
0 2436 5 1 1 2435
0 2437 7 1 2 2426 2436
0 2438 5 1 1 2437
0 2439 7 1 2 6508 2438
0 2440 5 2 1 2439
0 2441 7 1 2 6509 6514
0 2442 5 1 1 2441
0 2443 7 2 2 4478 2442
0 2444 5 2 1 6518
0 2445 7 1 2 4786 6515
0 2446 5 1 1 2445
0 2447 7 4 2 6520 2446
0 2448 5 1 1 6522
0 2449 7 1 2 4470 6504
0 2450 7 1 2 6523 2449
0 2451 5 2 1 2450
0 2452 7 1 2 6516 6526
0 2453 5 1 1 2452
0 2454 7 2 2 4471 2453
0 2455 5 2 1 6528
0 2456 7 1 2 4781 6517
0 2457 5 1 1 2456
0 2458 7 3 2 6530 2457
0 2459 5 1 1 6532
0 2460 7 2 2 4464 6533
0 2461 7 1 2 6524 6535
0 2462 5 2 1 2461
0 2463 7 1 2 6525 6529
0 2464 5 2 1 2463
0 2465 7 1 2 6505 6521
0 2466 5 1 1 2465
0 2467 7 1 2 2417 6519
0 2468 5 1 1 2467
0 2469 7 1 2 2466 2468
0 2470 7 1 2 6539 2469
0 2471 5 1 1 2470
0 2472 7 1 2 6527 2471
0 2473 5 2 1 2472
0 2474 7 1 2 6537 6541
0 2475 5 2 1 2474
0 2476 7 1 2 4465 6543
0 2477 5 2 1 2476
0 2478 7 1 2 4775 6542
0 2479 5 1 1 2478
0 2480 7 4 2 6545 2479
0 2481 5 1 1 6547
0 2482 7 2 2 4458 6548
0 2483 7 1 2 6534 6551
0 2484 5 2 1 2483
0 2485 7 1 2 2459 6546
0 2486 5 1 1 2485
0 2487 7 1 2 6536 6544
0 2488 5 2 1 2487
0 2489 7 1 2 2486 6555
0 2490 5 1 1 2489
0 2491 7 1 2 2448 6531
0 2492 5 1 1 2491
0 2493 7 1 2 6540 2492
0 2494 5 1 1 2493
0 2495 7 1 2 6556 2494
0 2496 5 1 1 2495
0 2497 7 2 2 6538 2496
0 2498 5 2 1 6557
0 2499 7 1 2 6552 6558
0 2500 5 1 1 2499
0 2501 7 1 2 2490 2500
0 2502 5 1 1 2501
0 2503 7 1 2 6553 2502
0 2504 5 2 1 2503
0 2505 7 1 2 6554 6559
0 2506 5 1 1 2505
0 2507 7 2 2 4459 2506
0 2508 5 2 1 6563
0 2509 7 1 2 4769 6560
0 2510 5 1 1 2509
0 2511 7 4 2 6565 2510
0 2512 5 1 1 6567
0 2513 7 1 2 4451 6549
0 2514 7 1 2 6568 2513
0 2515 5 2 1 2514
0 2516 7 1 2 6561 6571
0 2517 5 1 1 2516
0 2518 7 2 2 4452 2517
0 2519 5 2 1 6573
0 2520 7 1 2 4764 6562
0 2521 5 1 1 2520
0 2522 7 4 2 6575 2521
0 2523 5 1 1 6577
0 2524 7 1 2 4445 6569
0 2525 7 1 2 6578 2524
0 2526 5 2 1 2525
0 2527 7 1 2 6570 6574
0 2528 5 2 1 2527
0 2529 7 1 2 6550 6566
0 2530 5 1 1 2529
0 2531 7 1 2 2481 6564
0 2532 5 1 1 2531
0 2533 7 1 2 2530 2532
0 2534 7 1 2 6583 2533
0 2535 5 1 1 2534
0 2536 7 1 2 6572 2535
0 2537 5 2 1 2536
0 2538 7 1 2 6581 6585
0 2539 5 1 1 2538
0 2540 7 2 2 4446 2539
0 2541 5 2 1 6587
0 2542 7 1 2 4758 6586
0 2543 5 1 1 2542
0 2544 7 4 2 6589 2543
0 2545 5 1 1 6591
0 2546 7 2 2 4438 6592
0 2547 7 1 2 6579 6595
0 2548 5 2 1 2547
0 2549 7 1 2 2523 6590
0 2550 5 1 1 2549
0 2551 7 1 2 6580 6588
0 2552 5 2 1 2551
0 2553 7 1 2 2550 6599
0 2554 5 1 1 2553
0 2555 7 1 2 2512 6576
0 2556 5 1 1 2555
0 2557 7 1 2 6584 2556
0 2558 5 1 1 2557
0 2559 7 1 2 6600 2558
0 2560 5 1 1 2559
0 2561 7 2 2 6582 2560
0 2562 5 2 1 6601
0 2563 7 1 2 6596 6602
0 2564 5 1 1 2563
0 2565 7 1 2 2554 2564
0 2566 5 1 1 2565
0 2567 7 1 2 6597 2566
0 2568 5 2 1 2567
0 2569 7 1 2 6598 6603
0 2570 5 1 1 2569
0 2571 7 2 2 4439 2570
0 2572 5 2 1 6607
0 2573 7 1 2 4752 6604
0 2574 5 1 1 2573
0 2575 7 4 2 6609 2574
0 2576 5 1 1 6611
0 2577 7 1 2 4431 6593
0 2578 7 1 2 6612 2577
0 2579 5 2 1 2578
0 2580 7 1 2 6605 6615
0 2581 5 1 1 2580
0 2582 7 2 2 4432 2581
0 2583 5 2 1 6617
0 2584 7 1 2 4747 6606
0 2585 5 1 1 2584
0 2586 7 3 2 6619 2585
0 2587 5 1 1 6621
0 2588 7 2 2 4425 6622
0 2589 7 1 2 6613 6624
0 2590 5 2 1 2589
0 2591 7 1 2 6614 6618
0 2592 5 2 1 2591
0 2593 7 1 2 6594 6610
0 2594 5 1 1 2593
0 2595 7 1 2 2545 6608
0 2596 5 1 1 2595
0 2597 7 1 2 2594 2596
0 2598 7 1 2 6628 2597
0 2599 5 1 1 2598
0 2600 7 1 2 6616 2599
0 2601 5 2 1 2600
0 2602 7 1 2 6626 6630
0 2603 5 2 1 2602
0 2604 7 1 2 4426 6632
0 2605 5 2 1 2604
0 2606 7 1 2 4741 6631
0 2607 5 1 1 2606
0 2608 7 4 2 6634 2607
0 2609 5 1 1 6636
0 2610 7 2 2 4419 6637
0 2611 7 1 2 6623 6640
0 2612 5 2 1 2611
0 2613 7 1 2 2587 6635
0 2614 5 1 1 2613
0 2615 7 1 2 6625 6633
0 2616 5 2 1 2615
0 2617 7 1 2 2614 6644
0 2618 5 1 1 2617
0 2619 7 1 2 2576 6620
0 2620 5 1 1 2619
0 2621 7 1 2 6629 2620
0 2622 5 1 1 2621
0 2623 7 1 2 6645 2622
0 2624 5 1 1 2623
0 2625 7 2 2 6627 2624
0 2626 5 2 1 6646
0 2627 7 1 2 6641 6647
0 2628 5 1 1 2627
0 2629 7 1 2 2618 2628
0 2630 5 1 1 2629
0 2631 7 1 2 6642 2630
0 2632 5 2 1 2631
0 2633 7 1 2 6643 6648
0 2634 5 1 1 2633
0 2635 7 2 2 4420 2634
0 2636 5 2 1 6652
0 2637 7 1 2 4735 6649
0 2638 5 1 1 2637
0 2639 7 4 2 6654 2638
0 2640 5 1 1 6656
0 2641 7 1 2 4412 6638
0 2642 7 1 2 6657 2641
0 2643 5 2 1 2642
0 2644 7 1 2 6650 6660
0 2645 5 1 1 2644
0 2646 7 2 2 4413 2645
0 2647 5 2 1 6662
0 2648 7 1 2 4730 6651
0 2649 5 1 1 2648
0 2650 7 4 2 6664 2649
0 2651 5 1 1 6666
0 2652 7 1 2 4406 6658
0 2653 7 1 2 6667 2652
0 2654 5 2 1 2653
0 2655 7 1 2 6659 6663
0 2656 5 2 1 2655
0 2657 7 1 2 6639 6655
0 2658 5 1 1 2657
0 2659 7 1 2 2609 6653
0 2660 5 1 1 2659
0 2661 7 1 2 2658 2660
0 2662 7 1 2 6672 2661
0 2663 5 1 1 2662
0 2664 7 1 2 6661 2663
0 2665 5 2 1 2664
0 2666 7 1 2 6670 6674
0 2667 5 1 1 2666
0 2668 7 2 2 4407 2667
0 2669 5 2 1 6676
0 2670 7 1 2 4724 6675
0 2671 5 1 1 2670
0 2672 7 4 2 6678 2671
0 2673 5 1 1 6680
0 2674 7 2 2 4399 6681
0 2675 7 1 2 6668 6684
0 2676 5 2 1 2675
0 2677 7 1 2 6669 6677
0 2678 5 2 1 2677
0 2679 7 1 2 2640 6665
0 2680 5 1 1 2679
0 2681 7 1 2 6673 2680
0 2682 5 1 1 2681
0 2683 7 1 2 6688 2682
0 2684 5 1 1 2683
0 2685 7 2 2 6671 2684
0 2686 5 2 1 6690
0 2687 7 1 2 6686 6692
0 2688 5 1 1 2687
0 2689 7 2 2 4400 2688
0 2690 5 2 1 6694
0 2691 7 1 2 4718 6693
0 2692 5 1 1 2691
0 2693 7 4 2 6696 2692
0 2694 5 1 1 6698
0 2695 7 1 2 2651 6679
0 2696 5 1 1 2695
0 2697 7 1 2 6689 2696
0 2698 5 1 1 2697
0 2699 7 1 2 6685 6691
0 2700 5 1 1 2699
0 2701 7 1 2 2698 2700
0 2702 5 1 1 2701
0 2703 7 1 2 6687 2702
0 2704 5 2 1 2703
0 2705 7 1 2 4392 6682
0 2706 7 1 2 6699 2705
0 2707 5 2 1 2706
0 2708 7 1 2 6702 6704
0 2709 5 1 1 2708
0 2710 7 2 2 4393 2709
0 2711 5 2 1 6706
0 2712 7 1 2 4713 6703
0 2713 5 1 1 2712
0 2714 7 3 2 6708 2713
0 2715 5 1 1 6710
0 2716 7 2 2 4386 6711
0 2717 7 1 2 6700 6713
0 2718 5 2 1 2717
0 2719 7 1 2 6701 6707
0 2720 5 2 1 2719
0 2721 7 1 2 2694 6709
0 2722 5 1 1 2721
0 2723 7 1 2 6717 2722
0 2724 5 1 1 2723
0 2725 7 1 2 6683 6697
0 2726 5 1 1 2725
0 2727 7 1 2 2673 6695
0 2728 5 1 1 2727
0 2729 7 1 2 2726 2728
0 2730 7 1 2 6718 2729
0 2731 5 1 1 2730
0 2732 7 1 2 6705 2731
0 2733 5 2 1 2732
0 2734 7 1 2 6715 6719
0 2735 5 2 1 2734
0 2736 7 1 2 6714 6721
0 2737 5 2 1 2736
0 2738 7 1 2 2724 6723
0 2739 5 1 1 2738
0 2740 7 2 2 6716 2739
0 2741 5 2 1 6725
0 2742 7 1 2 4387 6722
0 2743 5 2 1 2742
0 2744 7 1 2 4707 6720
0 2745 5 1 1 2744
0 2746 7 4 2 6729 2745
0 2747 5 1 1 6731
0 2748 7 2 2 4380 6732
0 2749 7 1 2 6712 6735
0 2750 5 2 1 2749
0 2751 7 1 2 6727 6737
0 2752 5 1 1 2751
0 2753 7 2 2 4381 2752
0 2754 5 2 1 6739
0 2755 7 1 2 4701 6728
0 2756 5 1 1 2755
0 2757 7 3 2 6741 2756
0 2758 5 1 1 6743
0 2759 7 1 2 2715 6730
0 2760 5 1 1 2759
0 2761 7 1 2 6724 2760
0 2762 5 1 1 2761
0 2763 7 1 2 6726 6736
0 2764 5 1 1 2763
0 2765 7 1 2 2762 2764
0 2766 5 1 1 2765
0 2767 7 1 2 6738 2766
0 2768 5 2 1 2767
0 2769 7 1 2 4374 6733
0 2770 7 1 2 6744 2769
0 2771 5 2 1 2770
0 2772 7 1 2 6746 6748
0 2773 5 1 1 2772
0 2774 7 2 2 4375 2773
0 2775 5 2 1 6750
0 2776 7 1 2 2758 6752
0 2777 5 1 1 2776
0 2778 7 1 2 6745 6751
0 2779 5 2 1 2778
0 2780 7 2 2 2777 6754
0 2781 5 1 1 6756
0 2782 7 1 2 6734 6742
0 2783 5 1 1 2782
0 2784 7 1 2 2747 6740
0 2785 5 1 1 2784
0 2786 7 1 2 2783 2785
0 2787 7 1 2 6755 2786
0 2788 5 1 1 2787
0 2789 7 1 2 6749 2788
0 2790 5 1 1 2789
0 2791 7 1 2 4688 2790
0 2792 5 1 1 2791
0 2793 7 1 2 2781 2792
0 2794 5 1 1 2793
0 2795 7 1 2 4695 6747
0 2796 5 1 1 2795
0 2797 7 2 2 6753 2796
0 2798 5 1 1 6758
0 2799 7 1 2 6757 2798
0 2800 5 1 1 2799
0 2801 7 1 2 4689 6759
0 2802 5 1 1 2801
0 2803 7 1 2 2800 2802
0 2804 7 1 2 2794 2803
0 2805 5 1 1 2804
0 2806 7 1 2 1819 2805
0 2807 7 1 2 1188 2806
0 2808 7 2 2 1178 2807
0 2809 5 1 1 6760
0 2810 7 1 2 4702 4793
0 2811 5 2 1 2810
0 2812 7 1 2 4382 4486
0 2813 5 2 1 2812
0 2814 7 1 2 4696 4787
0 2815 5 2 1 2814
0 2816 7 1 2 4376 4479
0 2817 5 2 1 2816
0 2818 7 2 2 4371 4472
0 2819 5 3 1 6770
0 2820 7 1 2 6768 6772
0 2821 5 1 1 2820
0 2822 7 2 2 6766 2821
0 2823 5 2 1 6775
0 2824 7 1 2 6764 6777
0 2825 5 1 1 2824
0 2826 7 2 2 6762 2825
0 2827 5 1 1 6779
0 2828 7 1 2 4708 2827
0 2829 5 2 1 2828
0 2830 7 1 2 4388 6780
0 2831 5 2 1 2830
0 2832 7 1 2 4799 6783
0 2833 5 1 1 2832
0 2834 7 2 2 6781 2833
0 2835 5 1 1 6785
0 2836 7 1 2 4714 2835
0 2837 5 2 1 2836
0 2838 7 1 2 4394 6786
0 2839 5 2 1 2838
0 2840 7 1 2 4805 6789
0 2841 5 1 1 2840
0 2842 7 2 2 6787 2841
0 2843 5 1 1 6791
0 2844 7 1 2 4719 2843
0 2845 5 2 1 2844
0 2846 7 1 2 4401 6792
0 2847 5 2 1 2846
0 2848 7 1 2 4812 6795
0 2849 5 1 1 2848
0 2850 7 2 2 6793 2849
0 2851 5 1 1 6797
0 2852 7 1 2 4725 2851
0 2853 5 2 1 2852
0 2854 7 1 2 4408 6798
0 2855 5 2 1 2854
0 2856 7 1 2 4819 6801
0 2857 5 1 1 2856
0 2858 7 2 2 6799 2857
0 2859 5 1 1 6803
0 2860 7 1 2 4731 2859
0 2861 5 2 1 2860
0 2862 7 1 2 4414 6804
0 2863 5 2 1 2862
0 2864 7 1 2 4825 6807
0 2865 5 1 1 2864
0 2866 7 2 2 6805 2865
0 2867 5 1 1 6809
0 2868 7 1 2 4736 2867
0 2869 5 2 1 2868
0 2870 7 1 2 4421 6810
0 2871 5 2 1 2870
0 2872 7 1 2 4832 6813
0 2873 5 1 1 2872
0 2874 7 2 2 6811 2873
0 2875 5 1 1 6815
0 2876 7 1 2 4742 2875
0 2877 5 2 1 2876
0 2878 7 1 2 4427 6816
0 2879 5 2 1 2878
0 2880 7 1 2 4839 6819
0 2881 5 1 1 2880
0 2882 7 2 2 6817 2881
0 2883 5 1 1 6821
0 2884 7 1 2 4748 2883
0 2885 5 2 1 2884
0 2886 7 1 2 4433 6822
0 2887 5 2 1 2886
0 2888 7 1 2 4845 6825
0 2889 5 1 1 2888
0 2890 7 2 2 6823 2889
0 2891 5 1 1 6827
0 2892 7 1 2 4753 2891
0 2893 5 2 1 2892
0 2894 7 1 2 4440 6828
0 2895 5 2 1 2894
0 2896 7 1 2 4852 6831
0 2897 5 1 1 2896
0 2898 7 2 2 6829 2897
0 2899 5 1 1 6833
0 2900 7 1 2 4759 2899
0 2901 5 2 1 2900
0 2902 7 1 2 4447 6834
0 2903 5 2 1 2902
0 2904 7 1 2 4859 6837
0 2905 5 1 1 2904
0 2906 7 2 2 6835 2905
0 2907 5 1 1 6839
0 2908 7 1 2 4765 2907
0 2909 5 2 1 2908
0 2910 7 1 2 4453 6840
0 2911 5 2 1 2910
0 2912 7 1 2 4865 6843
0 2913 5 1 1 2912
0 2914 7 2 2 6841 2913
0 2915 5 1 1 6845
0 2916 7 1 2 4770 2915
0 2917 5 2 1 2916
0 2918 7 1 2 4460 6846
0 2919 5 2 1 2918
0 2920 7 1 2 4872 6849
0 2921 5 1 1 2920
0 2922 7 2 2 6847 2921
0 2923 5 1 1 6851
0 2924 7 1 2 4776 2923
0 2925 5 2 1 2924
0 2926 7 1 2 4466 6852
0 2927 5 2 1 2926
0 2928 7 1 2 4879 6855
0 2929 5 1 1 2928
0 2930 7 4 2 6853 2929
0 2931 5 3 1 6857
0 2932 7 2 2 6800 6802
0 2933 5 1 1 6864
0 2934 7 1 2 4511 6865
0 2935 5 1 1 2934
0 2936 7 1 2 4820 2933
0 2937 5 1 1 2936
0 2938 7 4 2 2935 2937
0 2939 5 3 1 6866
0 2940 7 1 2 4919 6867
0 2941 5 4 1 2940
0 2942 7 1 2 4616 6870
0 2943 5 3 1 2942
0 2944 7 2 2 6794 6796
0 2945 5 1 1 6880
0 2946 7 1 2 4505 6881
0 2947 5 1 1 2946
0 2948 7 1 2 4813 2945
0 2949 5 1 1 2948
0 2950 7 4 2 2947 2949
0 2951 5 3 1 6882
0 2952 7 1 2 4914 6883
0 2953 5 4 1 2952
0 2954 7 1 2 4609 6886
0 2955 5 3 1 2954
0 2956 7 2 2 6788 6790
0 2957 5 1 1 6896
0 2958 7 1 2 4499 6897
0 2959 5 1 1 2958
0 2960 7 1 2 4806 2957
0 2961 5 1 1 2960
0 2962 7 3 2 2959 2961
0 2963 5 2 1 6898
0 2964 7 1 2 4908 6899
0 2965 5 4 1 2964
0 2966 7 1 2 4603 6901
0 2967 5 3 1 2966
0 2968 7 2 2 6782 6784
0 2969 5 1 1 6910
0 2970 7 1 2 4492 6911
0 2971 5 1 1 2970
0 2972 7 1 2 4800 2969
0 2973 5 1 1 2972
0 2974 7 2 2 2971 2973
0 2975 5 2 1 6912
0 2976 7 1 2 4902 6913
0 2977 5 4 1 2976
0 2978 7 1 2 4596 6914
0 2979 5 3 1 2978
0 2980 7 2 2 6763 6765
0 2981 5 1 1 6923
0 2982 7 1 2 6776 2981
0 2983 5 1 1 2982
0 2984 7 1 2 6778 6924
0 2985 5 1 1 2984
0 2986 7 2 2 2983 2985
0 2987 5 1 1 6925
0 2988 7 1 2 4897 2987
0 2989 5 4 1 2988
0 2990 7 1 2 4589 6926
0 2991 5 3 1 2990
0 2992 7 2 2 6767 6769
0 2993 5 1 1 6934
0 2994 7 1 2 6771 2993
0 2995 5 1 1 2994
0 2996 7 1 2 6773 6935
0 2997 5 1 1 2996
0 2998 7 2 2 2995 2997
0 2999 5 1 1 6936
0 3000 7 1 2 4583 6937
0 3001 5 3 1 3000
0 3002 7 1 2 4891 2999
0 3003 5 3 1 3002
0 3004 7 1 2 4690 4782
0 3005 5 1 1 3004
0 3006 7 2 2 6774 3005
0 3007 5 1 1 6944
0 3008 7 2 2 4885 6945
0 3009 5 3 1 6946
0 3010 7 2 2 6941 6948
0 3011 5 1 1 6951
0 3012 7 3 2 6938 3011
0 3013 5 1 1 6953
0 3014 7 1 2 6931 6954
0 3015 5 1 1 3014
0 3016 7 2 2 6927 3015
0 3017 5 2 1 6956
0 3018 7 1 2 6920 6958
0 3019 5 1 1 3018
0 3020 7 2 2 6916 3019
0 3021 5 2 1 6960
0 3022 7 1 2 6907 6962
0 3023 5 1 1 3022
0 3024 7 2 2 6903 3023
0 3025 5 2 1 6964
0 3026 7 1 2 6893 6966
0 3027 5 1 1 3026
0 3028 7 2 2 6889 3027
0 3029 5 2 1 6968
0 3030 7 1 2 6877 6970
0 3031 5 1 1 3030
0 3032 7 2 2 6873 3031
0 3033 5 2 1 6972
0 3034 7 2 2 6806 6808
0 3035 5 1 1 6976
0 3036 7 1 2 4518 6977
0 3037 5 1 1 3036
0 3038 7 1 2 4826 3035
0 3039 5 1 1 3038
0 3040 7 4 2 3037 3039
0 3041 5 3 1 6978
0 3042 7 1 2 4925 6979
0 3043 5 4 1 3042
0 3044 7 1 2 4622 6982
0 3045 5 3 1 3044
0 3046 7 3 2 6985 6989
0 3047 5 2 1 6992
0 3048 7 1 2 6973 6995
0 3049 5 1 1 3048
0 3050 7 1 2 6974 6993
0 3051 5 1 1 3050
0 3052 7 4 2 3049 3051
0 3053 5 3 1 6997
0 3054 7 2 2 6824 6826
0 3055 5 1 1 7004
0 3056 7 1 2 4538 7005
0 3057 5 1 1 3056
0 3058 7 1 2 4846 3055
0 3059 5 1 1 3058
0 3060 7 4 2 3057 3059
0 3061 5 3 1 7006
0 3062 7 1 2 4942 7007
0 3063 5 4 1 3062
0 3064 7 1 2 4642 7010
0 3065 5 3 1 3064
0 3066 7 2 2 6818 6820
0 3067 5 1 1 7020
0 3068 7 1 2 4531 7021
0 3069 5 1 1 3068
0 3070 7 1 2 4840 3067
0 3071 5 1 1 3070
0 3072 7 2 2 3069 3071
0 3073 5 3 1 7022
0 3074 7 1 2 4936 7023
0 3075 5 4 1 3074
0 3076 7 1 2 4635 7024
0 3077 5 3 1 3076
0 3078 7 2 2 6812 6814
0 3079 5 1 1 7034
0 3080 7 1 2 4525 7035
0 3081 5 1 1 3080
0 3082 7 1 2 4833 3079
0 3083 5 1 1 3082
0 3084 7 4 2 3081 3083
0 3085 5 3 1 7036
0 3086 7 1 2 4931 7037
0 3087 5 4 1 3086
0 3088 7 1 2 4628 7040
0 3089 5 3 1 3088
0 3090 7 1 2 6990 6975
0 3091 5 1 1 3090
0 3092 7 2 2 6986 3091
0 3093 5 2 1 7050
0 3094 7 1 2 7047 7052
0 3095 5 1 1 3094
0 3096 7 2 2 7043 3095
0 3097 5 2 1 7054
0 3098 7 1 2 7031 7056
0 3099 5 1 1 3098
0 3100 7 2 2 7027 3099
0 3101 5 2 1 7058
0 3102 7 1 2 7017 7060
0 3103 5 1 1 3102
0 3104 7 2 2 7013 3103
0 3105 5 2 1 7062
0 3106 7 2 2 6830 6832
0 3107 5 1 1 7066
0 3108 7 1 2 4544 7067
0 3109 5 1 1 3108
0 3110 7 1 2 4853 3107
0 3111 5 1 1 3110
0 3112 7 2 2 3109 3111
0 3113 5 3 1 7068
0 3114 7 1 2 4947 7069
0 3115 5 4 1 3114
0 3116 7 1 2 4649 7070
0 3117 5 3 1 3116
0 3118 7 3 2 7073 7077
0 3119 5 2 1 7080
0 3120 7 1 2 7063 7083
0 3121 5 1 1 3120
0 3122 7 1 2 7064 7081
0 3123 5 1 1 3122
0 3124 7 4 2 3121 3123
0 3125 5 3 1 7085
0 3126 7 1 2 7001 7089
0 3127 5 2 1 3126
0 3128 7 1 2 6998 7086
0 3129 5 1 1 3128
0 3130 7 2 2 7092 3129
0 3131 5 1 1 7094
0 3132 7 3 2 7044 7048
0 3133 5 2 1 7096
0 3134 7 1 2 7051 7099
0 3135 5 1 1 3134
0 3136 7 1 2 7053 7097
0 3137 5 1 1 3136
0 3138 7 4 2 3135 3137
0 3139 5 3 1 7101
0 3140 7 1 2 7095 7105
0 3141 5 2 1 3140
0 3142 7 2 2 7093 7108
0 3143 5 1 1 7110
0 3144 7 3 2 7028 7032
0 3145 5 2 1 7112
0 3146 7 1 2 7055 7115
0 3147 5 1 1 3146
0 3148 7 1 2 7057 7113
0 3149 5 1 1 3148
0 3150 7 4 2 3147 3149
0 3151 5 3 1 7117
0 3152 7 2 2 6836 6838
0 3153 5 1 1 7124
0 3154 7 1 2 4550 7125
0 3155 5 1 1 3154
0 3156 7 1 2 4860 3153
0 3157 5 1 1 3156
0 3158 7 4 2 3155 3157
0 3159 5 3 1 7126
0 3160 7 1 2 4656 7130
0 3161 5 3 1 3160
0 3162 7 1 2 4953 7127
0 3163 5 4 1 3162
0 3164 7 3 2 7133 7136
0 3165 5 2 1 7140
0 3166 7 1 2 7078 7065
0 3167 5 1 1 3166
0 3168 7 2 2 7074 3167
0 3169 5 2 1 7145
0 3170 7 1 2 7143 7146
0 3171 5 1 1 3170
0 3172 7 1 2 7141 7147
0 3173 5 1 1 3172
0 3174 7 3 2 3171 3173
0 3175 5 2 1 7149
0 3176 7 1 2 7152 7106
0 3177 5 2 1 3176
0 3178 7 1 2 7150 7102
0 3179 5 1 1 3178
0 3180 7 2 2 7154 3179
0 3181 5 1 1 7156
0 3182 7 1 2 7121 7157
0 3183 5 2 1 3182
0 3184 7 1 2 7118 3181
0 3185 5 1 1 3184
0 3186 7 2 2 7158 3185
0 3187 5 1 1 7160
0 3188 7 1 2 3143 7161
0 3189 5 2 1 3188
0 3190 7 3 2 7014 7018
0 3191 5 2 1 7164
0 3192 7 1 2 7059 7167
0 3193 5 1 1 3192
0 3194 7 1 2 7061 7165
0 3195 5 1 1 3194
0 3196 7 4 2 3193 3195
0 3197 5 3 1 7169
0 3198 7 3 2 6874 6878
0 3199 5 2 1 7176
0 3200 7 1 2 6969 7179
0 3201 5 1 1 3200
0 3202 7 1 2 6971 7177
0 3203 5 1 1 3202
0 3204 7 4 2 3201 3203
0 3205 5 3 1 7181
0 3206 7 1 2 7173 7185
0 3207 5 2 1 3206
0 3208 7 1 2 7170 7182
0 3209 5 1 1 3208
0 3210 7 2 2 7188 3209
0 3211 5 1 1 7190
0 3212 7 1 2 7191 7002
0 3213 5 2 1 3212
0 3214 7 2 2 7189 7192
0 3215 5 1 1 7194
0 3216 7 1 2 3131 7103
0 3217 5 1 1 3216
0 3218 7 2 2 7109 3217
0 3219 5 1 1 7196
0 3220 7 1 2 3215 7197
0 3221 5 2 1 3220
0 3222 7 3 2 6890 6894
0 3223 5 2 1 7200
0 3224 7 1 2 6965 7203
0 3225 5 1 1 3224
0 3226 7 1 2 6967 7201
0 3227 5 1 1 3226
0 3228 7 4 2 3225 3227
0 3229 5 3 1 7205
0 3230 7 1 2 7122 7209
0 3231 5 2 1 3230
0 3232 7 1 2 7119 7206
0 3233 5 1 1 3232
0 3234 7 2 2 7212 3233
0 3235 5 1 1 7214
0 3236 7 1 2 7186 7215
0 3237 5 2 1 3236
0 3238 7 2 2 7213 7216
0 3239 5 1 1 7218
0 3240 7 1 2 3211 6999
0 3241 5 1 1 3240
0 3242 7 2 2 7193 3241
0 3243 5 1 1 7220
0 3244 7 1 2 3239 7221
0 3245 5 2 1 3244
0 3246 7 3 2 6904 6908
0 3247 5 2 1 7224
0 3248 7 1 2 6961 7227
0 3249 5 1 1 3248
0 3250 7 1 2 6963 7225
0 3251 5 1 1 3250
0 3252 7 4 2 3249 3251
0 3253 5 3 1 7229
0 3254 7 1 2 7107 7233
0 3255 5 2 1 3254
0 3256 7 1 2 7104 7230
0 3257 5 1 1 3256
0 3258 7 2 2 7236 3257
0 3259 5 1 1 7238
0 3260 7 1 2 7210 7239
0 3261 5 2 1 3260
0 3262 7 2 2 7237 7240
0 3263 5 1 1 7242
0 3264 7 1 2 7183 3235
0 3265 5 1 1 3264
0 3266 7 2 2 7217 3265
0 3267 5 1 1 7244
0 3268 7 1 2 3263 7245
0 3269 5 2 1 3268
0 3270 7 3 2 6917 6921
0 3271 5 2 1 7248
0 3272 7 1 2 6957 7251
0 3273 5 1 1 3272
0 3274 7 1 2 6959 7249
0 3275 5 1 1 3274
0 3276 7 5 2 3273 3275
0 3277 5 3 1 7253
0 3278 7 1 2 7003 7258
0 3279 5 2 1 3278
0 3280 7 1 2 7000 7254
0 3281 5 1 1 3280
0 3282 7 2 2 7261 3281
0 3283 5 1 1 7263
0 3284 7 1 2 7234 7264
0 3285 5 2 1 3284
0 3286 7 2 2 7262 7265
0 3287 5 1 1 7267
0 3288 7 1 2 7207 3259
0 3289 5 1 1 3288
0 3290 7 2 2 7241 3289
0 3291 5 1 1 7269
0 3292 7 1 2 3287 7270
0 3293 5 2 1 3292
0 3294 7 3 2 6928 6932
0 3295 5 2 1 7273
0 3296 7 1 2 6955 7274
0 3297 5 1 1 3296
0 3298 7 1 2 3013 7276
0 3299 5 1 1 3298
0 3300 7 4 2 3297 3299
0 3301 5 3 1 7278
0 3302 7 1 2 7187 7282
0 3303 5 2 1 3302
0 3304 7 1 2 7184 7279
0 3305 5 1 1 3304
0 3306 7 2 2 7285 3305
0 3307 5 1 1 7287
0 3308 7 1 2 7259 7288
0 3309 5 2 1 3308
0 3310 7 2 2 7286 7289
0 3311 5 1 1 7291
0 3312 7 1 2 7231 3283
0 3313 5 1 1 3312
0 3314 7 2 2 7266 3313
0 3315 5 1 1 7293
0 3316 7 1 2 3311 7294
0 3317 5 2 1 3316
0 3318 7 3 2 6939 6942
0 3319 5 2 1 7297
0 3320 7 1 2 6947 7300
0 3321 5 1 1 3320
0 3322 7 1 2 6949 7298
0 3323 5 1 1 3322
0 3324 7 3 2 3321 3323
0 3325 5 3 1 7302
0 3326 7 1 2 7211 7303
0 3327 5 2 1 3326
0 3328 7 1 2 7208 7305
0 3329 5 1 1 3328
0 3330 7 2 2 7308 3329
0 3331 5 1 1 7310
0 3332 7 1 2 7283 7311
0 3333 5 2 1 3332
0 3334 7 2 2 7309 7312
0 3335 5 1 1 7314
0 3336 7 1 2 7255 3307
0 3337 5 1 1 3336
0 3338 7 2 2 7290 3337
0 3339 5 1 1 7316
0 3340 7 1 2 3335 7317
0 3341 5 2 1 3340
0 3342 7 2 2 7235 7304
0 3343 5 2 1 7320
0 3344 7 1 2 7280 3331
0 3345 5 1 1 3344
0 3346 7 2 2 7313 3345
0 3347 5 1 1 7324
0 3348 7 1 2 7321 7325
0 3349 5 2 1 3348
0 3350 7 1 2 7322 3347
0 3351 5 1 1 3350
0 3352 7 2 2 7326 3351
0 3353 5 1 1 7328
0 3354 7 2 2 4577 3007
0 3355 5 3 1 7330
0 3356 7 3 2 6950 7332
0 3357 5 5 1 7335
0 3358 7 1 2 7232 7306
0 3359 5 1 1 3358
0 3360 7 2 2 7323 3359
0 3361 5 2 1 7343
0 3362 7 1 2 7256 7345
0 3363 5 1 1 3362
0 3364 7 2 2 7338 3363
0 3365 5 1 1 7347
0 3366 7 1 2 7329 7348
0 3367 5 2 1 3366
0 3368 7 2 2 7327 7349
0 3369 5 1 1 7351
0 3370 7 1 2 7315 3339
0 3371 5 1 1 3370
0 3372 7 2 2 7318 3371
0 3373 5 1 1 7353
0 3374 7 1 2 3369 7354
0 3375 5 2 1 3374
0 3376 7 2 2 7319 7355
0 3377 5 1 1 7357
0 3378 7 1 2 7292 3315
0 3379 5 1 1 3378
0 3380 7 2 2 7295 3379
0 3381 5 1 1 7359
0 3382 7 1 2 3377 7360
0 3383 5 2 1 3382
0 3384 7 2 2 7296 7361
0 3385 5 1 1 7363
0 3386 7 1 2 7268 3291
0 3387 5 1 1 3386
0 3388 7 2 2 7271 3387
0 3389 5 1 1 7365
0 3390 7 1 2 3385 7366
0 3391 5 2 1 3390
0 3392 7 2 2 7272 7367
0 3393 5 1 1 7369
0 3394 7 1 2 7243 3267
0 3395 5 1 1 3394
0 3396 7 2 2 7246 3395
0 3397 5 1 1 7371
0 3398 7 1 2 3393 7372
0 3399 5 2 1 3398
0 3400 7 2 2 7247 7373
0 3401 5 1 1 7375
0 3402 7 1 2 7219 3243
0 3403 5 1 1 3402
0 3404 7 2 2 7222 3403
0 3405 5 1 1 7377
0 3406 7 1 2 3401 7378
0 3407 5 2 1 3406
0 3408 7 2 2 7223 7379
0 3409 5 1 1 7381
0 3410 7 1 2 7195 3219
0 3411 5 1 1 3410
0 3412 7 2 2 7198 3411
0 3413 5 1 1 7383
0 3414 7 1 2 3409 7384
0 3415 5 2 1 3414
0 3416 7 2 2 7199 7385
0 3417 5 1 1 7387
0 3418 7 1 2 7111 3187
0 3419 5 1 1 3418
0 3420 7 2 2 7162 3419
0 3421 5 1 1 7389
0 3422 7 1 2 3417 7390
0 3423 5 2 1 3422
0 3424 7 2 2 7163 7391
0 3425 5 1 1 7393
0 3426 7 2 2 7155 7159
0 3427 5 1 1 7395
0 3428 7 1 2 7134 7148
0 3429 5 1 1 3428
0 3430 7 2 2 7137 3429
0 3431 5 2 1 7397
0 3432 7 2 2 6842 6844
0 3433 5 1 1 7401
0 3434 7 1 2 4557 7402
0 3435 5 1 1 3434
0 3436 7 1 2 4866 3433
0 3437 5 1 1 3436
0 3438 7 4 2 3435 3437
0 3439 5 3 1 7403
0 3440 7 1 2 4959 7404
0 3441 5 4 1 3440
0 3442 7 1 2 4664 7407
0 3443 5 3 1 3442
0 3444 7 3 2 7410 7414
0 3445 5 2 1 7417
0 3446 7 1 2 7398 7420
0 3447 5 1 1 3446
0 3448 7 1 2 7399 7418
0 3449 5 1 1 3448
0 3450 7 3 2 3447 3449
0 3451 5 2 1 7422
0 3452 7 1 2 7425 7123
0 3453 5 2 1 3452
0 3454 7 1 2 7423 7120
0 3455 5 1 1 3454
0 3456 7 2 2 7427 3455
0 3457 5 1 1 7429
0 3458 7 1 2 7174 7430
0 3459 5 2 1 3458
0 3460 7 1 2 7171 3457
0 3461 5 1 1 3460
0 3462 7 2 2 7431 3461
0 3463 5 1 1 7433
0 3464 7 1 2 3427 7434
0 3465 5 2 1 3464
0 3466 7 1 2 7396 3463
0 3467 5 1 1 3466
0 3468 7 2 2 7435 3467
0 3469 5 1 1 7437
0 3470 7 1 2 3425 7438
0 3471 5 2 1 3470
0 3472 7 1 2 7394 3469
0 3473 5 1 1 3472
0 3474 7 2 2 7439 3473
0 3475 5 1 1 7441
0 3476 7 1 2 6858 3475
0 3477 5 1 1 3476
0 3478 7 2 2 6854 6856
0 3479 5 1 1 7443
0 3480 7 1 2 4570 7444
0 3481 5 1 1 3480
0 3482 7 1 2 4880 3479
0 3483 5 1 1 3482
0 3484 7 4 2 3481 3483
0 3485 5 3 1 7445
0 3486 7 1 2 7388 3421
0 3487 5 1 1 3486
0 3488 7 2 2 7392 3487
0 3489 5 1 1 7452
0 3490 7 1 2 7449 7453
0 3491 5 1 1 3490
0 3492 7 2 2 6848 6850
0 3493 5 1 1 7454
0 3494 7 1 2 4564 7455
0 3495 5 1 1 3494
0 3496 7 1 2 4873 3493
0 3497 5 1 1 3496
0 3498 7 4 2 3495 3497
0 3499 5 3 1 7456
0 3500 7 1 2 7376 3405
0 3501 5 1 1 3500
0 3502 7 2 2 7380 3501
0 3503 5 1 1 7463
0 3504 7 1 2 7405 3503
0 3505 5 1 1 3504
0 3506 7 1 2 7408 7464
0 3507 5 1 1 3506
0 3508 7 1 2 7370 3397
0 3509 5 1 1 3508
0 3510 7 2 2 7374 3509
0 3511 5 1 1 7465
0 3512 7 1 2 7128 3511
0 3513 5 1 1 3512
0 3514 7 1 2 7131 7466
0 3515 5 1 1 3514
0 3516 7 1 2 7364 3389
0 3517 5 1 1 3516
0 3518 7 2 2 7368 3517
0 3519 5 1 1 7467
0 3520 7 1 2 7358 3381
0 3521 5 1 1 3520
0 3522 7 2 2 7362 3521
0 3523 5 1 1 7469
0 3524 7 1 2 7011 7470
0 3525 5 1 1 3524
0 3526 7 1 2 7008 3523
0 3527 5 1 1 3526
0 3528 7 1 2 7352 3373
0 3529 5 1 1 3528
0 3530 7 2 2 7356 3529
0 3531 5 1 1 7471
0 3532 7 1 2 3353 3365
0 3533 5 1 1 3532
0 3534 7 2 2 7350 3533
0 3535 5 1 1 7473
0 3536 7 1 2 7041 7474
0 3537 5 1 1 3536
0 3538 7 1 2 7038 3535
0 3539 5 1 1 3538
0 3540 7 2 2 7257 7339
0 3541 5 2 1 7475
0 3542 7 1 2 7344 7477
0 3543 5 1 1 3542
0 3544 7 1 2 7346 7476
0 3545 5 1 1 3544
0 3546 7 2 2 3543 3545
0 3547 5 1 1 7479
0 3548 7 1 2 6983 3547
0 3549 5 1 1 3548
0 3550 7 1 2 6980 7480
0 3551 5 1 1 3550
0 3552 7 1 2 7260 7336
0 3553 5 1 1 3552
0 3554 7 2 2 7478 3553
0 3555 5 1 1 7481
0 3556 7 1 2 6868 7482
0 3557 5 1 1 3556
0 3558 7 1 2 6884 7281
0 3559 5 1 1 3558
0 3560 7 1 2 6887 7284
0 3561 5 1 1 3560
0 3562 7 2 2 6915 7340
0 3563 5 1 1 7483
0 3564 7 1 2 6900 3563
0 3565 5 2 1 3564
0 3566 7 1 2 6902 7484
0 3567 5 2 1 3566
0 3568 7 1 2 7307 7487
0 3569 5 1 1 3568
0 3570 7 1 2 7485 3569
0 3571 5 1 1 3570
0 3572 7 1 2 3561 3571
0 3573 5 1 1 3572
0 3574 7 1 2 3559 3573
0 3575 7 1 2 3557 3574
0 3576 5 1 1 3575
0 3577 7 1 2 6871 3555
0 3578 5 1 1 3577
0 3579 7 1 2 3576 3578
0 3580 5 1 1 3579
0 3581 7 1 2 3551 3580
0 3582 5 1 1 3581
0 3583 7 1 2 3549 3582
0 3584 5 1 1 3583
0 3585 7 1 2 3539 3584
0 3586 5 1 1 3585
0 3587 7 2 2 3537 3586
0 3588 5 1 1 7489
0 3589 7 1 2 7472 3588
0 3590 5 1 1 3589
0 3591 7 1 2 3531 7490
0 3592 5 1 1 3591
0 3593 7 1 2 7025 3592
0 3594 5 1 1 3593
0 3595 7 1 2 3590 3594
0 3596 5 1 1 3595
0 3597 7 1 2 3527 3596
0 3598 5 1 1 3597
0 3599 7 2 2 3525 3598
0 3600 5 1 1 7491
0 3601 7 1 2 7468 3600
0 3602 5 1 1 3601
0 3603 7 1 2 3519 7492
0 3604 5 1 1 3603
0 3605 7 1 2 7071 3604
0 3606 5 1 1 3605
0 3607 7 1 2 3602 3606
0 3608 7 1 2 3515 3607
0 3609 5 1 1 3608
0 3610 7 1 2 3513 3609
0 3611 5 1 1 3610
0 3612 7 1 2 3507 3611
0 3613 5 1 1 3612
0 3614 7 2 2 3505 3613
0 3615 5 1 1 7493
0 3616 7 1 2 7460 7494
0 3617 5 1 1 3616
0 3618 7 1 2 7457 3615
0 3619 5 1 1 3618
0 3620 7 1 2 7382 3413
0 3621 5 1 1 3620
0 3622 7 1 2 7386 3621
0 3623 7 1 2 3619 3622
0 3624 5 1 1 3623
0 3625 7 1 2 3617 3624
0 3626 7 1 2 3491 3625
0 3627 5 1 1 3626
0 3628 7 1 2 7446 3489
0 3629 5 1 1 3628
0 3630 7 1 2 3627 3629
0 3631 7 1 2 3477 3630
0 3632 5 1 1 3631
0 3633 7 2 2 4971 6859
0 3634 5 5 1 7495
0 3635 7 1 2 4685 6861
0 3636 5 5 1 3635
0 3637 7 1 2 4967 7447
0 3638 5 4 1 3637
0 3639 7 1 2 4679 7450
0 3640 5 3 1 3639
0 3641 7 1 2 4964 7458
0 3642 5 4 1 3641
0 3643 7 1 2 4672 7461
0 3644 5 3 1 3643
0 3645 7 1 2 7415 7400
0 3646 5 1 1 3645
0 3647 7 2 2 7411 3646
0 3648 5 2 1 7521
0 3649 7 1 2 7518 7523
0 3650 5 1 1 3649
0 3651 7 2 2 7514 3650
0 3652 5 2 1 7525
0 3653 7 1 2 7511 7527
0 3654 5 1 1 3653
0 3655 7 3 2 7507 3654
0 3656 5 3 1 7529
0 3657 7 1 2 7502 7532
0 3658 5 1 1 3657
0 3659 7 3 2 7497 3658
0 3660 5 2 1 7535
0 3661 7 3 2 7508 7512
0 3662 5 2 1 7540
0 3663 7 1 2 7526 7543
0 3664 5 1 1 3663
0 3665 7 1 2 7528 7541
0 3666 5 1 1 3665
0 3667 7 3 2 3664 3666
0 3668 5 2 1 7545
0 3669 7 1 2 7538 7548
0 3670 5 1 1 3669
0 3671 7 2 2 7536 7546
0 3672 5 1 1 7550
0 3673 7 1 2 3670 3672
0 3674 5 2 1 3673
0 3675 7 1 2 7498 7533
0 3676 5 1 1 3675
0 3677 7 1 2 7503 7530
0 3678 5 1 1 3677
0 3679 7 1 2 3676 3678
0 3680 7 1 2 7552 3679
0 3681 5 1 1 3680
0 3682 7 3 2 7515 7519
0 3683 5 2 1 7554
0 3684 7 1 2 7522 7557
0 3685 5 1 1 3684
0 3686 7 1 2 7524 7555
0 3687 5 1 1 3686
0 3688 7 4 2 3685 3687
0 3689 5 2 1 7559
0 3690 7 1 2 7539 7560
0 3691 5 1 1 3690
0 3692 7 1 2 7537 7563
0 3693 5 1 1 3692
0 3694 7 2 2 3691 3693
0 3695 5 1 1 7565
0 3696 7 1 2 7426 3695
0 3697 5 1 1 3696
0 3698 7 1 2 3681 3697
0 3699 7 1 2 3632 3698
0 3700 7 1 2 7553 7566
0 3701 7 3 2 7504 7499
0 3702 5 2 1 7567
0 3703 7 1 2 7570 7531
0 3704 5 1 1 3703
0 3705 7 1 2 7568 7534
0 3706 5 1 1 3705
0 3707 7 2 2 3704 3706
0 3708 5 1 1 7572
0 3709 7 1 2 7153 3708
0 3710 5 2 1 3709
0 3711 7 2 2 7151 7573
0 3712 5 1 1 7576
0 3713 7 1 2 7574 3712
0 3714 5 1 1 3713
0 3715 7 1 2 6862 7442
0 3716 5 1 1 3715
0 3717 7 1 2 3714 3716
0 3718 7 1 2 3700 3717
0 3719 7 1 2 7549 7090
0 3720 5 1 1 3719
0 3721 7 1 2 7547 7087
0 3722 5 1 1 3721
0 3723 7 1 2 3720 3722
0 3724 5 1 1 3723
0 3725 7 1 2 7551 7577
0 3726 7 1 2 3724 3725
0 3727 7 1 2 6940 7333
0 3728 5 1 1 3727
0 3729 7 2 2 6943 3728
0 3730 5 2 1 7578
0 3731 7 1 2 6933 7580
0 3732 5 1 1 3731
0 3733 7 2 2 6929 3732
0 3734 5 2 1 7582
0 3735 7 1 2 6922 7584
0 3736 5 1 1 3735
0 3737 7 2 2 6918 3736
0 3738 5 2 1 7586
0 3739 7 1 2 6909 7588
0 3740 5 1 1 3739
0 3741 7 2 2 6905 3740
0 3742 5 2 1 7590
0 3743 7 1 2 6895 7592
0 3744 5 1 1 3743
0 3745 7 2 2 6891 3744
0 3746 5 2 1 7594
0 3747 7 1 2 6879 7596
0 3748 5 1 1 3747
0 3749 7 2 2 6875 3748
0 3750 5 2 1 7598
0 3751 7 1 2 6991 7600
0 3752 5 1 1 3751
0 3753 7 2 2 6987 3752
0 3754 5 2 1 7602
0 3755 7 1 2 7049 7604
0 3756 5 1 1 3755
0 3757 7 2 2 7045 3756
0 3758 5 2 1 7606
0 3759 7 1 2 7033 7608
0 3760 5 1 1 3759
0 3761 7 2 2 7029 3760
0 3762 5 2 1 7610
0 3763 7 1 2 7019 7612
0 3764 5 1 1 3763
0 3765 7 2 2 7015 3764
0 3766 5 2 1 7614
0 3767 7 1 2 7079 7616
0 3768 5 1 1 3767
0 3769 7 2 2 7075 3768
0 3770 5 2 1 7618
0 3771 7 1 2 7135 7620
0 3772 5 1 1 3771
0 3773 7 2 2 7138 3772
0 3774 5 2 1 7622
0 3775 7 1 2 7416 7624
0 3776 5 1 1 3775
0 3777 7 2 2 7412 3776
0 3778 5 2 1 7626
0 3779 7 1 2 7520 7628
0 3780 5 1 1 3779
0 3781 7 2 2 7516 3780
0 3782 5 2 1 7630
0 3783 7 1 2 7513 7632
0 3784 5 1 1 3783
0 3785 7 3 2 7509 3784
0 3786 5 2 1 7634
0 3787 7 1 2 7505 7637
0 3788 5 1 1 3787
0 3789 7 5 2 7500 3788
0 3790 5 4 1 7639
0 3791 7 1 2 7564 7175
0 3792 5 2 1 3791
0 3793 7 1 2 7561 7172
0 3794 5 1 1 3793
0 3795 7 2 2 7648 3794
0 3796 5 1 1 7650
0 3797 7 1 2 7091 7651
0 3798 5 2 1 3797
0 3799 7 1 2 7088 3796
0 3800 5 1 1 3799
0 3801 7 1 2 7652 3800
0 3802 5 1 1 3801
0 3803 7 1 2 7440 3802
0 3804 7 1 2 7640 3803
0 3805 7 1 2 7424 7428
0 3806 7 1 2 7562 3805
0 3807 7 1 2 7432 3806
0 3808 7 1 2 7649 3807
0 3809 7 1 2 7436 3808
0 3810 7 1 2 7653 3809
0 3811 7 1 2 7575 3810
0 3812 7 1 2 3804 3811
0 3813 7 1 2 3726 3812
0 3814 7 1 2 3718 3813
0 3815 7 1 2 3699 3814
0 3816 5 1 1 3815
0 3817 7 1 2 7084 7615
0 3818 5 1 1 3817
0 3819 7 1 2 7082 7617
0 3820 5 1 1 3819
0 3821 7 3 2 3818 3820
0 3822 5 3 1 7654
0 3823 7 1 2 6996 7599
0 3824 5 1 1 3823
0 3825 7 1 2 6994 7601
0 3826 5 1 1 3825
0 3827 7 4 2 3824 3826
0 3828 5 3 1 7660
0 3829 7 1 2 7655 7661
0 3830 5 2 1 3829
0 3831 7 1 2 7100 7603
0 3832 5 1 1 3831
0 3833 7 1 2 7098 7605
0 3834 5 1 1 3833
0 3835 7 4 2 3832 3834
0 3836 5 3 1 7669
0 3837 7 1 2 7657 7664
0 3838 5 1 1 3837
0 3839 7 2 2 7667 3838
0 3840 5 1 1 7676
0 3841 7 1 2 7670 7677
0 3842 5 2 1 3841
0 3843 7 2 2 7668 7678
0 3844 5 1 1 7680
0 3845 7 1 2 7144 7619
0 3846 5 1 1 3845
0 3847 7 1 2 7142 7621
0 3848 5 1 1 3847
0 3849 7 3 2 3846 3848
0 3850 5 3 1 7682
0 3851 7 1 2 7683 7671
0 3852 5 2 1 3851
0 3853 7 1 2 7685 7673
0 3854 5 1 1 3853
0 3855 7 2 2 7688 3854
0 3856 5 1 1 7690
0 3857 7 1 2 7116 7607
0 3858 5 1 1 3857
0 3859 7 1 2 7114 7609
0 3860 5 1 1 3859
0 3861 7 4 2 3858 3860
0 3862 5 3 1 7692
0 3863 7 1 2 7691 7693
0 3864 5 2 1 3863
0 3865 7 1 2 3856 7696
0 3866 5 1 1 3865
0 3867 7 2 2 7699 3866
0 3868 5 1 1 7701
0 3869 7 1 2 3844 7702
0 3870 5 2 1 3869
0 3871 7 1 2 7168 7611
0 3872 5 1 1 3871
0 3873 7 1 2 7166 7613
0 3874 5 1 1 3873
0 3875 7 4 2 3872 3874
0 3876 5 3 1 7705
0 3877 7 1 2 7180 7595
0 3878 5 1 1 3877
0 3879 7 1 2 7178 7597
0 3880 5 1 1 3879
0 3881 7 4 2 3878 3880
0 3882 5 3 1 7712
0 3883 7 1 2 7706 7713
0 3884 5 2 1 3883
0 3885 7 1 2 7709 7716
0 3886 5 1 1 3885
0 3887 7 2 2 7719 3886
0 3888 5 1 1 7721
0 3889 7 1 2 7662 7722
0 3890 5 2 1 3889
0 3891 7 2 2 7720 7723
0 3892 5 1 1 7725
0 3893 7 1 2 7674 3840
0 3894 5 1 1 3893
0 3895 7 2 2 7679 3894
0 3896 5 1 1 7727
0 3897 7 1 2 3892 7728
0 3898 5 2 1 3897
0 3899 7 1 2 7204 7591
0 3900 5 1 1 3899
0 3901 7 1 2 7202 7593
0 3902 5 1 1 3901
0 3903 7 4 2 3900 3902
0 3904 5 3 1 7731
0 3905 7 1 2 7694 7732
0 3906 5 2 1 3905
0 3907 7 1 2 7697 7735
0 3908 5 1 1 3907
0 3909 7 2 2 7738 3908
0 3910 5 1 1 7740
0 3911 7 1 2 7714 7741
0 3912 5 2 1 3911
0 3913 7 2 2 7739 7742
0 3914 5 1 1 7744
0 3915 7 1 2 7665 3888
0 3916 5 1 1 3915
0 3917 7 2 2 7724 3916
0 3918 5 1 1 7746
0 3919 7 1 2 3914 7747
0 3920 5 2 1 3919
0 3921 7 1 2 7228 7587
0 3922 5 1 1 3921
0 3923 7 1 2 7226 7589
0 3924 5 1 1 3923
0 3925 7 4 2 3922 3924
0 3926 5 3 1 7750
0 3927 7 1 2 7672 7751
0 3928 5 2 1 3927
0 3929 7 1 2 7675 7754
0 3930 5 1 1 3929
0 3931 7 2 2 7757 3930
0 3932 5 1 1 7759
0 3933 7 1 2 7733 7760
0 3934 5 2 1 3933
0 3935 7 2 2 7758 7761
0 3936 5 1 1 7763
0 3937 7 1 2 7717 3910
0 3938 5 1 1 3937
0 3939 7 2 2 7743 3938
0 3940 5 1 1 7765
0 3941 7 1 2 3936 7766
0 3942 5 2 1 3941
0 3943 7 1 2 7250 7585
0 3944 5 1 1 3943
0 3945 7 1 2 7252 7583
0 3946 5 1 1 3945
0 3947 7 4 2 3944 3946
0 3948 5 4 1 7769
0 3949 7 1 2 7663 7770
0 3950 5 2 1 3949
0 3951 7 1 2 7666 7773
0 3952 5 1 1 3951
0 3953 7 2 2 7777 3952
0 3954 5 1 1 7779
0 3955 7 1 2 7752 7780
0 3956 5 2 1 3955
0 3957 7 2 2 7778 7781
0 3958 5 1 1 7783
0 3959 7 1 2 7736 3932
0 3960 5 1 1 3959
0 3961 7 2 2 7762 3960
0 3962 5 1 1 7785
0 3963 7 1 2 3958 7786
0 3964 5 2 1 3963
0 3965 7 1 2 7275 7581
0 3966 5 1 1 3965
0 3967 7 1 2 7277 7579
0 3968 5 1 1 3967
0 3969 7 4 2 3966 3968
0 3970 5 2 1 7789
0 3971 7 1 2 7715 7790
0 3972 5 2 1 3971
0 3973 7 1 2 7718 7793
0 3974 5 1 1 3973
0 3975 7 2 2 7795 3974
0 3976 5 1 1 7797
0 3977 7 1 2 7771 7798
0 3978 5 2 1 3977
0 3979 7 2 2 7796 7799
0 3980 5 1 1 7801
0 3981 7 1 2 7755 3954
0 3982 5 1 1 3981
0 3983 7 2 2 7782 3982
0 3984 5 1 1 7803
0 3985 7 1 2 3980 7804
0 3986 5 2 1 3985
0 3987 7 1 2 7299 7334
0 3988 5 1 1 3987
0 3989 7 1 2 7301 7331
0 3990 5 1 1 3989
0 3991 7 3 2 3988 3990
0 3992 5 3 1 7807
0 3993 7 1 2 7734 7808
0 3994 5 2 1 3993
0 3995 7 1 2 7737 7810
0 3996 5 1 1 3995
0 3997 7 2 2 7813 3996
0 3998 5 1 1 7815
0 3999 7 1 2 7791 7816
0 4000 5 2 1 3999
0 4001 7 2 2 7814 7817
0 4002 5 1 1 7819
0 4003 7 1 2 7774 3976
0 4004 5 1 1 4003
0 4005 7 2 2 7800 4004
0 4006 5 1 1 7821
0 4007 7 1 2 4002 7822
0 4008 5 2 1 4007
0 4009 7 2 2 7753 7809
0 4010 5 2 1 7825
0 4011 7 1 2 7794 3998
0 4012 5 1 1 4011
0 4013 7 2 2 7818 4012
0 4014 5 1 1 7829
0 4015 7 1 2 7826 7830
0 4016 5 2 1 4015
0 4017 7 1 2 7827 4014
0 4018 5 1 1 4017
0 4019 7 2 2 7831 4018
0 4020 5 1 1 7833
0 4021 7 1 2 7756 7811
0 4022 5 1 1 4021
0 4023 7 2 2 7828 4022
0 4024 5 2 1 7835
0 4025 7 1 2 7775 7837
0 4026 5 1 1 4025
0 4027 7 2 2 7341 4026
0 4028 5 1 1 7839
0 4029 7 1 2 7834 7840
0 4030 5 2 1 4029
0 4031 7 2 2 7832 7841
0 4032 5 1 1 7843
0 4033 7 1 2 7820 4006
0 4034 5 1 1 4033
0 4035 7 2 2 7823 4034
0 4036 5 1 1 7845
0 4037 7 1 2 4032 7846
0 4038 5 2 1 4037
0 4039 7 2 2 7824 7847
0 4040 5 1 1 7849
0 4041 7 1 2 7802 3984
0 4042 5 1 1 4041
0 4043 7 2 2 7805 4042
0 4044 5 1 1 7851
0 4045 7 1 2 4040 7852
0 4046 5 2 1 4045
0 4047 7 2 2 7806 7853
0 4048 5 1 1 7855
0 4049 7 1 2 7784 3962
0 4050 5 1 1 4049
0 4051 7 2 2 7787 4050
0 4052 5 1 1 7857
0 4053 7 1 2 4048 7858
0 4054 5 2 1 4053
0 4055 7 2 2 7788 7859
0 4056 5 1 1 7861
0 4057 7 1 2 7764 3940
0 4058 5 1 1 4057
0 4059 7 2 2 7767 4058
0 4060 5 1 1 7863
0 4061 7 1 2 4056 7864
0 4062 5 2 1 4061
0 4063 7 2 2 7768 7865
0 4064 5 1 1 7867
0 4065 7 1 2 7745 3918
0 4066 5 1 1 4065
0 4067 7 2 2 7748 4066
0 4068 5 1 1 7869
0 4069 7 1 2 4064 7870
0 4070 5 2 1 4069
0 4071 7 2 2 7749 7871
0 4072 5 1 1 7873
0 4073 7 1 2 7726 3896
0 4074 5 1 1 4073
0 4075 7 2 2 7729 4074
0 4076 5 1 1 7875
0 4077 7 1 2 4072 7876
0 4078 5 2 1 4077
0 4079 7 2 2 7730 7877
0 4080 5 1 1 7879
0 4081 7 1 2 7681 3868
0 4082 5 1 1 4081
0 4083 7 2 2 7703 4082
0 4084 5 1 1 7881
0 4085 7 1 2 4080 7882
0 4086 5 2 1 4085
0 4087 7 2 2 7704 7883
0 4088 5 1 1 7885
0 4089 7 2 2 7689 7700
0 4090 5 1 1 7887
0 4091 7 1 2 7421 7623
0 4092 5 1 1 4091
0 4093 7 1 2 7419 7625
0 4094 5 1 1 4093
0 4095 7 2 2 4092 4094
0 4096 5 2 1 7889
0 4097 7 1 2 7695 7890
0 4098 5 2 1 4097
0 4099 7 1 2 7698 7891
0 4100 5 1 1 4099
0 4101 7 2 2 7893 4100
0 4102 5 1 1 7895
0 4103 7 1 2 7896 7707
0 4104 5 2 1 4103
0 4105 7 1 2 4102 7710
0 4106 5 1 1 4105
0 4107 7 2 2 7897 4106
0 4108 5 1 1 7899
0 4109 7 1 2 4090 7900
0 4110 5 2 1 4109
0 4111 7 1 2 7888 4108
0 4112 5 1 1 4111
0 4113 7 2 2 7901 4112
0 4114 5 1 1 7903
0 4115 7 1 2 4088 7904
0 4116 5 2 1 4115
0 4117 7 1 2 7886 4114
0 4118 5 1 1 4117
0 4119 7 2 2 7905 4118
0 4120 5 1 1 7907
0 4121 7 1 2 6860 4120
0 4122 5 1 1 4121
0 4123 7 1 2 7880 4084
0 4124 5 1 1 4123
0 4125 7 2 2 7884 4124
0 4126 5 1 1 7909
0 4127 7 1 2 7451 7910
0 4128 5 1 1 4127
0 4129 7 1 2 7868 4068
0 4130 5 1 1 4129
0 4131 7 2 2 7872 4130
0 4132 5 1 1 7911
0 4133 7 1 2 7406 4132
0 4134 5 1 1 4133
0 4135 7 1 2 7409 7912
0 4136 5 1 1 4135
0 4137 7 1 2 7862 4060
0 4138 5 1 1 4137
0 4139 7 2 2 7866 4138
0 4140 5 1 1 7913
0 4141 7 1 2 7129 4140
0 4142 5 1 1 4141
0 4143 7 1 2 7132 7914
0 4144 5 1 1 4143
0 4145 7 1 2 7856 4052
0 4146 5 1 1 4145
0 4147 7 2 2 7860 4146
0 4148 5 1 1 7915
0 4149 7 1 2 7850 4044
0 4150 5 1 1 4149
0 4151 7 2 2 7854 4150
0 4152 5 1 1 7917
0 4153 7 1 2 7012 7918
0 4154 5 1 1 4153
0 4155 7 1 2 7009 4152
0 4156 5 1 1 4155
0 4157 7 1 2 7844 4036
0 4158 5 1 1 4157
0 4159 7 2 2 7848 4158
0 4160 5 1 1 7919
0 4161 7 1 2 4020 4028
0 4162 5 1 1 4161
0 4163 7 2 2 7842 4162
0 4164 5 1 1 7921
0 4165 7 1 2 7042 7922
0 4166 5 1 1 4165
0 4167 7 1 2 7039 4164
0 4168 5 1 1 4167
0 4169 7 2 2 7342 7776
0 4170 5 2 1 7923
0 4171 7 1 2 7836 7925
0 4172 5 1 1 4171
0 4173 7 1 2 7838 7924
0 4174 5 1 1 4173
0 4175 7 2 2 4172 4174
0 4176 5 1 1 7927
0 4177 7 1 2 6984 4176
0 4178 5 1 1 4177
0 4179 7 1 2 6981 7928
0 4180 5 1 1 4179
0 4181 7 1 2 7337 7772
0 4182 5 1 1 4181
0 4183 7 2 2 7926 4182
0 4184 5 1 1 7929
0 4185 7 1 2 6872 4184
0 4186 5 1 1 4185
0 4187 7 1 2 6869 7930
0 4188 5 1 1 4187
0 4189 7 1 2 7488 7812
0 4190 5 1 1 4189
0 4191 7 2 2 7486 4190
0 4192 5 1 1 7931
0 4193 7 1 2 6885 4192
0 4194 5 1 1 4193
0 4195 7 1 2 7792 4194
0 4196 5 1 1 4195
0 4197 7 1 2 6888 7932
0 4198 5 1 1 4197
0 4199 7 1 2 4196 4198
0 4200 5 1 1 4199
0 4201 7 1 2 4188 4200
0 4202 5 1 1 4201
0 4203 7 1 2 4186 4202
0 4204 5 1 1 4203
0 4205 7 1 2 4180 4204
0 4206 5 1 1 4205
0 4207 7 1 2 4178 4206
0 4208 5 1 1 4207
0 4209 7 1 2 4168 4208
0 4210 5 1 1 4209
0 4211 7 2 2 4166 4210
0 4212 5 1 1 7933
0 4213 7 1 2 7920 4212
0 4214 5 1 1 4213
0 4215 7 1 2 4160 7934
0 4216 5 1 1 4215
0 4217 7 1 2 7026 4216
0 4218 5 1 1 4217
0 4219 7 1 2 4214 4218
0 4220 5 1 1 4219
0 4221 7 1 2 4156 4220
0 4222 5 1 1 4221
0 4223 7 2 2 4154 4222
0 4224 5 1 1 7935
0 4225 7 1 2 7916 4224
0 4226 5 1 1 4225
0 4227 7 1 2 4148 7936
0 4228 5 1 1 4227
0 4229 7 1 2 7072 4228
0 4230 5 1 1 4229
0 4231 7 1 2 4226 4230
0 4232 7 1 2 4144 4231
0 4233 5 1 1 4232
0 4234 7 1 2 4142 4233
0 4235 5 1 1 4234
0 4236 7 1 2 4136 4235
0 4237 5 1 1 4236
0 4238 7 2 2 4134 4237
0 4239 5 1 1 7937
0 4240 7 1 2 7462 7938
0 4241 5 1 1 4240
0 4242 7 1 2 7459 4239
0 4243 5 1 1 4242
0 4244 7 1 2 7874 4076
0 4245 5 1 1 4244
0 4246 7 1 2 7878 4245
0 4247 7 1 2 4243 4246
0 4248 5 1 1 4247
0 4249 7 1 2 4241 4248
0 4250 7 1 2 4128 4249
0 4251 5 1 1 4250
0 4252 7 1 2 7448 4126
0 4253 5 1 1 4252
0 4254 7 1 2 4251 4253
0 4255 7 1 2 4122 4254
0 4256 5 1 1 4255
0 4257 7 1 2 7571 7635
0 4258 5 1 1 4257
0 4259 7 1 2 7569 7638
0 4260 5 1 1 4259
0 4261 7 2 2 4258 4260
0 4262 5 1 1 7939
0 4263 7 1 2 7686 7940
0 4264 5 1 1 4263
0 4265 7 1 2 7544 7631
0 4266 5 1 1 4265
0 4267 7 1 2 7542 7633
0 4268 5 1 1 4267
0 4269 7 3 2 4266 4268
0 4270 5 3 1 7941
0 4271 7 1 2 7641 7944
0 4272 5 1 1 4271
0 4273 7 1 2 7684 4262
0 4274 5 1 1 4273
0 4275 7 1 2 4272 4274
0 4276 7 1 2 4264 4275
0 4277 7 1 2 7558 7627
0 4278 5 1 1 4277
0 4279 7 1 2 7556 7629
0 4280 5 1 1 4279
0 4281 7 5 2 4278 4280
0 4282 5 3 1 7947
0 4283 7 1 2 7948 7708
0 4284 5 2 1 4283
0 4285 7 1 2 7952 7711
0 4286 5 1 1 4285
0 4287 7 2 2 7955 4286
0 4288 5 1 1 7957
0 4289 7 1 2 7958 7656
0 4290 5 2 1 4289
0 4291 7 1 2 7687 7658
0 4292 7 1 2 7892 4291
0 4293 7 1 2 7956 4292
0 4294 7 1 2 7902 4293
0 4295 7 1 2 7945 4294
0 4296 7 1 2 7959 4295
0 4297 7 1 2 7644 7906
0 4298 7 1 2 4296 4297
0 4299 7 1 2 7949 7942
0 4300 5 1 1 4299
0 4301 7 1 2 7506 7636
0 4302 5 1 1 4301
0 4303 7 1 2 7496 4302
0 4304 7 1 2 4300 4303
0 4305 5 1 1 4304
0 4306 7 2 2 7894 7898
0 4307 5 1 1 7961
0 4308 7 1 2 4288 7659
0 4309 5 1 1 4308
0 4310 7 2 2 7960 4309
0 4311 5 1 1 7963
0 4312 7 1 2 4307 7964
0 4313 5 2 1 4312
0 4314 7 1 2 4305 7965
0 4315 7 1 2 4298 4314
0 4316 7 1 2 4276 4315
0 4317 7 1 2 4256 4316
0 4318 7 1 2 7642 7943
0 4319 5 1 1 4318
0 4320 7 1 2 7645 7946
0 4321 5 1 1 4320
0 4322 7 2 2 4319 4321
0 4323 5 1 1 7967
0 4324 7 1 2 7950 7968
0 4325 5 1 1 4324
0 4326 7 1 2 7953 4323
0 4327 5 1 1 4326
0 4328 7 1 2 4325 4327
0 4329 5 1 1 4328
0 4330 7 1 2 7646 7954
0 4331 5 1 1 4330
0 4332 7 1 2 7643 7951
0 4333 5 1 1 4332
0 4334 7 1 2 4331 4333
0 4335 5 1 1 4334
0 4336 7 1 2 7962 4311
0 4337 5 1 1 4336
0 4338 7 1 2 7966 4337
0 4339 5 1 1 4338
0 4340 7 1 2 6863 7908
0 4341 5 1 1 4340
0 4342 7 1 2 4339 4341
0 4343 7 1 2 4335 4342
0 4344 7 1 2 4329 4343
0 4345 7 1 2 4317 4344
0 4346 5 1 1 4345
0 4347 7 1 2 3816 4346
0 4348 7 1 2 2809 4347
0 4349 5 1 1 4348
0 4350 7 1 2 6930 6952
0 4351 7 1 2 6919 4350
0 4352 7 1 2 6906 4351
0 4353 7 1 2 6892 4352
0 4354 7 1 2 6876 4353
0 4355 7 1 2 6988 4354
0 4356 7 1 2 7046 4355
0 4357 7 1 2 7030 4356
0 4358 7 1 2 7016 4357
0 4359 7 1 2 7076 4358
0 4360 7 1 2 7139 4359
0 4361 7 1 2 7413 4360
0 4362 7 1 2 7517 4361
0 4363 7 1 2 7501 4362
0 4364 7 1 2 7510 4363
0 4365 7 1 2 7647 4364
0 4366 5 1 1 4365
0 4367 7 1 2 6761 4366
0 4368 5 1 1 4367
3 9999 7 0 2 4349 4368
