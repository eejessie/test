1 0 0 8 0
2 16 1 0
2 17 1 0
2 18 1 0
2 19 1 0
2 20 1 0
2 21 1 0
2 22 1 0
2 23 1 0
1 1 0 8 0
2 24 1 1
2 25 1 1
2 26 1 1
2 27 1 1
2 28 1 1
2 29 1 1
2 30 1 1
2 31 1 1
1 2 0 8 0
2 32 1 2
2 41 1 2
2 64 1 2
2 103 1 2
2 158 1 2
2 230 1 2
2 327 1 2
2 436 1 2
1 3 0 8 0
2 541 1 3
2 631 1 3
2 712 1 3
2 777 1 3
2 830 1 3
2 869 1 3
2 887 1 3
2 895 1 3
1 4 0 8 0
2 896 1 4
2 897 1 4
2 898 1 4
2 899 1 4
2 900 1 4
2 901 1 4
2 902 1 4
2 903 1 4
1 5 0 8 0
2 904 1 5
2 905 1 5
2 906 1 5
2 907 1 5
2 908 1 5
2 909 1 5
2 910 1 5
2 911 1 5
1 6 0 8 0
2 912 1 6
2 913 1 6
2 914 1 6
2 915 1 6
2 916 1 6
2 917 1 6
2 918 1 6
2 919 1 6
1 7 0 8 0
2 920 1 7
2 921 1 7
2 922 1 7
2 923 1 7
2 924 1 7
2 925 1 7
2 926 1 7
2 927 1 7
1 8 0 8 0
2 928 1 8
2 929 1 8
2 930 1 8
2 931 1 8
2 932 1 8
2 933 1 8
2 934 1 8
2 935 1 8
1 9 0 8 0
2 936 1 9
2 937 1 9
2 938 1 9
2 939 1 9
2 940 1 9
2 941 1 9
2 942 1 9
2 943 1 9
1 10 0 8 0
2 944 1 10
2 945 1 10
2 946 1 10
2 947 1 10
2 948 1 10
2 949 1 10
2 950 1 10
2 951 1 10
1 11 0 8 0
2 952 1 11
2 953 1 11
2 954 1 11
2 955 1 11
2 956 1 11
2 957 1 11
2 958 1 11
2 959 1 11
1 12 0 8 0
2 960 1 12
2 961 1 12
2 962 1 12
2 963 1 12
2 964 1 12
2 965 1 12
2 966 1 12
2 967 1 12
1 13 0 8 0
2 968 1 13
2 969 1 13
2 970 1 13
2 971 1 13
2 972 1 13
2 973 1 13
2 974 1 13
2 975 1 13
1 14 0 9 0
2 976 1 14
2 977 1 14
2 978 1 14
2 979 1 14
2 980 1 14
2 981 1 14
2 982 1 14
2 983 1 14
2 984 1 14
1 15 0 8 0
2 985 1 15
2 986 1 15
2 987 1 15
2 988 1 15
2 989 1 15
2 990 1 15
2 991 1 15
2 992 1 15
2 993 1 33
2 994 1 33
2 995 1 35
2 996 1 35
2 997 1 39
2 998 1 39
2 999 1 40
2 1000 1 40
2 1001 1 42
2 1002 1 42
2 1003 1 44
2 1004 1 44
2 1005 1 46
2 1006 1 46
2 1007 1 51
2 1008 1 51
2 1009 1 52
2 1010 1 52
2 1011 1 55
2 1012 1 55
2 1013 1 58
2 1014 1 58
2 1015 1 60
2 1016 1 60
2 1017 1 61
2 1018 1 61
2 1019 1 65
2 1020 1 65
2 1021 1 67
2 1022 1 67
2 1023 1 69
2 1024 1 69
2 1025 1 71
2 1026 1 71
2 1027 1 73
2 1028 1 73
2 1029 1 78
2 1030 1 78
2 1031 1 79
2 1032 1 79
2 1033 1 82
2 1034 1 82
2 1035 1 85
2 1036 1 85
2 1037 1 88
2 1038 1 88
2 1039 1 91
2 1040 1 91
2 1041 1 94
2 1042 1 94
2 1043 1 97
2 1044 1 97
2 1045 1 99
2 1046 1 99
2 1047 1 100
2 1048 1 100
2 1049 1 104
2 1050 1 104
2 1051 1 106
2 1052 1 106
2 1053 1 108
2 1054 1 108
2 1055 1 110
2 1056 1 110
2 1057 1 112
2 1058 1 112
2 1059 1 117
2 1060 1 117
2 1061 1 118
2 1062 1 118
2 1063 1 121
2 1064 1 121
2 1065 1 124
2 1066 1 124
2 1067 1 127
2 1068 1 127
2 1069 1 130
2 1070 1 130
2 1071 1 132
2 1072 1 132
2 1073 1 134
2 1074 1 134
2 1075 1 138
2 1076 1 138
2 1077 1 139
2 1078 1 139
2 1079 1 140
2 1080 1 140
2 1081 1 143
2 1082 1 143
2 1083 1 146
2 1084 1 146
2 1085 1 148
2 1086 1 148
2 1087 1 149
2 1088 1 149
2 1089 1 152
2 1090 1 152
2 1091 1 154
2 1092 1 154
2 1093 1 155
2 1094 1 155
2 1095 1 159
2 1096 1 159
2 1097 1 161
2 1098 1 161
2 1099 1 163
2 1100 1 163
2 1101 1 165
2 1102 1 165
2 1103 1 170
2 1104 1 170
2 1105 1 171
2 1106 1 171
2 1107 1 174
2 1108 1 174
2 1109 1 177
2 1110 1 177
2 1111 1 179
2 1112 1 179
2 1113 1 181
2 1114 1 181
2 1115 1 183
2 1116 1 183
2 1117 1 185
2 1118 1 185
2 1119 1 190
2 1120 1 190
2 1121 1 191
2 1122 1 191
2 1123 1 194
2 1124 1 194
2 1125 1 197
2 1126 1 197
2 1127 1 200
2 1128 1 200
2 1129 1 203
2 1130 1 203
2 1131 1 206
2 1132 1 206
2 1133 1 209
2 1134 1 209
2 1135 1 212
2 1136 1 212
2 1137 1 215
2 1138 1 215
2 1139 1 218
2 1140 1 218
2 1141 1 221
2 1142 1 221
2 1143 1 221
2 1144 1 221
2 1145 1 223
2 1146 1 223
2 1147 1 231
2 1148 1 231
2 1149 1 233
2 1150 1 233
2 1151 1 235
2 1152 1 235
2 1153 1 237
2 1154 1 237
2 1155 1 239
2 1156 1 239
2 1157 1 240
2 1158 1 240
2 1159 1 243
2 1160 1 243
2 1161 1 245
2 1162 1 245
2 1163 1 247
2 1164 1 247
2 1165 1 249
2 1166 1 249
2 1167 1 251
2 1168 1 251
2 1169 1 256
2 1170 1 256
2 1171 1 257
2 1172 1 257
2 1173 1 260
2 1174 1 260
2 1175 1 263
2 1176 1 263
2 1177 1 265
2 1178 1 265
2 1179 1 267
2 1180 1 267
2 1181 1 269
2 1182 1 269
2 1183 1 271
2 1184 1 271
2 1185 1 276
2 1186 1 276
2 1187 1 277
2 1188 1 277
2 1189 1 280
2 1190 1 280
2 1191 1 283
2 1192 1 283
2 1193 1 286
2 1194 1 286
2 1195 1 289
2 1196 1 289
2 1197 1 292
2 1198 1 292
2 1199 1 295
2 1200 1 295
2 1201 1 298
2 1202 1 298
2 1203 1 301
2 1204 1 301
2 1205 1 304
2 1206 1 304
2 1207 1 307
2 1208 1 307
2 1209 1 309
2 1210 1 309
2 1211 1 310
2 1212 1 310
2 1213 1 313
2 1214 1 313
2 1215 1 316
2 1216 1 316
2 1217 1 319
2 1218 1 319
2 1219 1 321
2 1220 1 321
2 1221 1 324
2 1222 1 324
2 1223 1 328
2 1224 1 328
2 1225 1 330
2 1226 1 330
2 1227 1 332
2 1228 1 332
2 1229 1 334
2 1230 1 334
2 1231 1 336
2 1232 1 336
2 1233 1 339
2 1234 1 339
2 1235 1 342
2 1236 1 342
2 1237 1 345
2 1238 1 345
2 1239 1 348
2 1240 1 348
2 1241 1 350
2 1242 1 350
2 1243 1 352
2 1244 1 352
2 1245 1 354
2 1246 1 354
2 1247 1 356
2 1248 1 356
2 1249 1 361
2 1250 1 361
2 1251 1 362
2 1252 1 362
2 1253 1 365
2 1254 1 365
2 1255 1 368
2 1256 1 368
2 1257 1 370
2 1258 1 370
2 1259 1 372
2 1260 1 372
2 1261 1 374
2 1262 1 374
2 1263 1 375
2 1264 1 375
2 1265 1 376
2 1266 1 376
2 1267 1 381
2 1268 1 381
2 1269 1 382
2 1270 1 382
2 1271 1 385
2 1272 1 385
2 1273 1 388
2 1274 1 388
2 1275 1 391
2 1276 1 391
2 1277 1 394
2 1278 1 394
2 1279 1 397
2 1280 1 397
2 1281 1 400
2 1282 1 400
2 1283 1 403
2 1284 1 403
2 1285 1 406
2 1286 1 406
2 1287 1 409
2 1288 1 409
2 1289 1 412
2 1290 1 412
2 1291 1 415
2 1292 1 415
2 1293 1 418
2 1294 1 418
2 1295 1 421
2 1296 1 421
2 1297 1 424
2 1298 1 424
2 1299 1 427
2 1300 1 427
2 1301 1 430
2 1302 1 430
2 1303 1 433
2 1304 1 433
2 1305 1 437
2 1306 1 437
2 1307 1 439
2 1308 1 439
2 1309 1 441
2 1310 1 441
2 1311 1 443
2 1312 1 443
2 1313 1 445
2 1314 1 445
2 1315 1 447
2 1316 1 447
2 1317 1 449
2 1318 1 449
2 1319 1 452
2 1320 1 452
2 1321 1 455
2 1322 1 455
2 1323 1 458
2 1324 1 458
2 1325 1 461
2 1326 1 461
2 1327 1 463
2 1328 1 463
2 1329 1 465
2 1330 1 465
2 1331 1 467
2 1332 1 467
2 1333 1 469
2 1334 1 469
2 1335 1 474
2 1336 1 474
2 1337 1 475
2 1338 1 475
2 1339 1 478
2 1340 1 478
2 1341 1 481
2 1342 1 481
2 1343 1 483
2 1344 1 483
2 1345 1 485
2 1346 1 485
2 1347 1 487
2 1348 1 487
2 1349 1 492
2 1350 1 492
2 1351 1 493
2 1352 1 493
2 1353 1 496
2 1354 1 496
2 1355 1 499
2 1356 1 499
2 1357 1 502
2 1358 1 502
2 1359 1 505
2 1360 1 505
2 1361 1 508
2 1362 1 508
2 1363 1 511
2 1364 1 511
2 1365 1 514
2 1366 1 514
2 1367 1 517
2 1368 1 517
2 1369 1 520
2 1370 1 520
2 1371 1 523
2 1372 1 523
2 1373 1 526
2 1374 1 526
2 1375 1 529
2 1376 1 529
2 1377 1 532
2 1378 1 532
2 1379 1 535
2 1380 1 535
2 1381 1 538
2 1382 1 538
2 1383 1 542
2 1384 1 542
2 1385 1 544
2 1386 1 544
2 1387 1 546
2 1388 1 546
2 1389 1 548
2 1390 1 548
2 1391 1 550
2 1392 1 550
2 1393 1 552
2 1394 1 552
2 1395 1 554
2 1396 1 554
2 1397 1 557
2 1398 1 557
2 1399 1 560
2 1400 1 560
2 1401 1 563
2 1402 1 563
2 1403 1 566
2 1404 1 566
2 1405 1 568
2 1406 1 568
2 1407 1 570
2 1408 1 570
2 1409 1 572
2 1410 1 572
2 1411 1 574
2 1412 1 574
2 1413 1 579
2 1414 1 579
2 1415 1 580
2 1416 1 580
2 1417 1 583
2 1418 1 583
2 1419 1 586
2 1420 1 586
2 1421 1 589
2 1422 1 589
2 1423 1 592
2 1424 1 592
2 1425 1 595
2 1426 1 595
2 1427 1 598
2 1428 1 598
2 1429 1 601
2 1430 1 601
2 1431 1 604
2 1432 1 604
2 1433 1 607
2 1434 1 607
2 1435 1 610
2 1436 1 610
2 1437 1 613
2 1438 1 613
2 1439 1 616
2 1440 1 616
2 1441 1 619
2 1442 1 619
2 1443 1 622
2 1444 1 622
2 1445 1 625
2 1446 1 625
2 1447 1 628
2 1448 1 628
2 1449 1 632
2 1450 1 632
2 1451 1 634
2 1452 1 634
2 1453 1 636
2 1454 1 636
2 1455 1 638
2 1456 1 638
2 1457 1 640
2 1458 1 640
2 1459 1 642
2 1460 1 642
2 1461 1 644
2 1462 1 644
2 1463 1 647
2 1464 1 647
2 1465 1 650
2 1466 1 650
2 1467 1 653
2 1468 1 653
2 1469 1 656
2 1470 1 656
2 1471 1 658
2 1472 1 658
2 1473 1 660
2 1474 1 660
2 1475 1 662
2 1476 1 662
2 1477 1 664
2 1478 1 664
2 1479 1 669
2 1480 1 669
2 1481 1 670
2 1482 1 670
2 1483 1 673
2 1484 1 673
2 1485 1 676
2 1486 1 676
2 1487 1 679
2 1488 1 679
2 1489 1 682
2 1490 1 682
2 1491 1 685
2 1492 1 685
2 1493 1 688
2 1494 1 688
2 1495 1 691
2 1496 1 691
2 1497 1 694
2 1498 1 694
2 1499 1 697
2 1500 1 697
2 1501 1 700
2 1502 1 700
2 1503 1 703
2 1504 1 703
2 1505 1 706
2 1506 1 706
2 1507 1 709
2 1508 1 709
2 1509 1 713
2 1510 1 713
2 1511 1 715
2 1512 1 715
2 1513 1 717
2 1514 1 717
2 1515 1 719
2 1516 1 719
2 1517 1 721
2 1518 1 721
2 1519 1 723
2 1520 1 723
2 1521 1 725
2 1522 1 725
2 1523 1 728
2 1524 1 728
2 1525 1 731
2 1526 1 731
2 1527 1 734
2 1528 1 734
2 1529 1 737
2 1530 1 737
2 1531 1 739
2 1532 1 739
2 1533 1 741
2 1534 1 741
2 1535 1 745
2 1536 1 745
2 1537 1 746
2 1538 1 746
2 1539 1 747
2 1540 1 747
2 1541 1 749
2 1542 1 749
2 1543 1 750
2 1544 1 750
2 1545 1 753
2 1546 1 753
2 1547 1 756
2 1548 1 756
2 1549 1 759
2 1550 1 759
2 1551 1 762
2 1552 1 762
2 1553 1 765
2 1554 1 765
2 1555 1 768
2 1556 1 768
2 1557 1 771
2 1558 1 771
2 1559 1 774
2 1560 1 774
2 1561 1 778
2 1562 1 778
2 1563 1 780
2 1564 1 780
2 1565 1 782
2 1566 1 782
2 1567 1 784
2 1568 1 784
2 1569 1 786
2 1570 1 786
2 1571 1 789
2 1572 1 789
2 1573 1 793
2 1574 1 793
2 1575 1 794
2 1576 1 794
2 1577 1 797
2 1578 1 797
2 1579 1 800
2 1580 1 800
2 1581 1 802
2 1582 1 802
2 1583 1 803
2 1584 1 803
2 1585 1 806
2 1586 1 806
2 1587 1 809
2 1588 1 809
2 1589 1 812
2 1590 1 812
2 1591 1 815
2 1592 1 815
2 1593 1 818
2 1594 1 818
2 1595 1 821
2 1596 1 821
2 1597 1 824
2 1598 1 824
2 1599 1 827
2 1600 1 827
2 1601 1 831
2 1602 1 831
2 1603 1 833
2 1604 1 833
2 1605 1 835
2 1606 1 835
2 1607 1 837
2 1608 1 837
2 1609 1 839
2 1610 1 839
2 1611 1 844
2 1612 1 844
2 1613 1 844
2 1614 1 845
2 1615 1 845
2 1616 1 848
2 1617 1 848
2 1618 1 851
2 1619 1 851
2 1620 1 854
2 1621 1 854
2 1622 1 857
2 1623 1 857
2 1624 1 860
2 1625 1 860
2 1626 1 863
2 1627 1 863
2 1628 1 866
2 1629 1 866
2 1630 1 870
2 1631 1 870
2 1632 1 872
2 1633 1 872
2 1634 1 875
2 1635 1 875
2 1636 1 878
2 1637 1 878
2 1638 1 881
2 1639 1 881
2 1640 1 883
2 1641 1 883
2 1642 1 884
2 1643 1 884
3 1784 7 0 2 16 928
0 33 7 2 2 17 936
0 34 5 1 1 993
0 35 7 2 2 24 929
0 36 5 1 1 995
0 37 7 1 2 34 36
0 38 5 1 1 37
0 39 7 2 2 994 996
0 40 5 2 1 997
3 1785 7 0 2 38 999
0 42 7 2 2 18 944
0 43 5 1 1 1001
0 44 7 2 2 25 937
0 45 5 1 1 1003
0 46 7 2 2 32 930
0 47 5 1 1 1005
0 48 7 1 2 45 47
0 49 5 1 1 48
0 50 7 1 2 1004 1006
0 51 5 2 1 50
0 52 7 2 2 49 1007
0 53 5 1 1 1009
0 54 7 1 2 1002 1010
0 55 5 2 1 54
0 56 7 1 2 43 53
0 57 5 1 1 56
0 58 7 2 2 1011 57
0 59 5 1 1 1013
0 60 7 2 2 998 1014
0 61 5 2 1 1015
0 62 7 1 2 1000 59
0 63 5 1 1 62
3 1786 7 0 2 1017 63
0 65 7 2 2 19 952
0 66 5 1 1 1019
0 67 7 2 2 1008 1012
0 68 5 1 1 1021
0 69 7 2 2 26 945
0 70 5 1 1 1023
0 71 7 2 2 41 938
0 72 5 1 1 1025
0 73 7 2 2 541 931
0 74 5 1 1 1027
0 75 7 1 2 72 74
0 76 5 1 1 75
0 77 7 1 2 1026 1028
0 78 5 2 1 77
0 79 7 2 2 76 1029
0 80 5 1 1 1031
0 81 7 1 2 1024 1032
0 82 5 2 1 81
0 83 7 1 2 70 80
0 84 5 1 1 83
0 85 7 2 2 1033 84
0 86 5 1 1 1035
0 87 7 1 2 68 1036
0 88 5 2 1 87
0 89 7 1 2 1022 86
0 90 5 1 1 89
0 91 7 2 2 1037 90
0 92 5 1 1 1039
0 93 7 1 2 1020 1040
0 94 5 2 1 93
0 95 7 1 2 66 92
0 96 5 1 1 95
0 97 7 2 2 1041 96
0 98 5 1 1 1043
0 99 7 2 2 1016 1044
0 100 5 2 1 1045
0 101 7 1 2 1018 98
0 102 5 1 1 101
3 1787 7 0 2 1047 102
0 104 7 2 2 1038 1042
0 105 5 1 1 1049
0 106 7 2 2 1030 1034
0 107 5 1 1 1051
0 108 7 2 2 64 946
0 109 5 1 1 1053
0 110 7 2 2 631 939
0 111 5 1 1 1055
0 112 7 2 2 896 932
0 113 5 1 1 1057
0 114 7 1 2 111 113
0 115 5 1 1 114
0 116 7 1 2 1056 1058
0 117 5 2 1 116
0 118 7 2 2 115 1059
0 119 5 1 1 1061
0 120 7 1 2 1054 1062
0 121 5 2 1 120
0 122 7 1 2 109 119
0 123 5 1 1 122
0 124 7 2 2 1063 123
0 125 5 1 1 1065
0 126 7 1 2 107 1066
0 127 5 2 1 126
0 128 7 1 2 1052 125
0 129 5 1 1 128
0 130 7 2 2 1067 129
0 131 5 1 1 1069
0 132 7 2 2 20 960
0 133 5 1 1 1071
0 134 7 2 2 27 953
0 135 5 1 1 1073
0 136 7 1 2 133 135
0 137 5 1 1 136
0 138 7 2 2 1072 1074
0 139 5 2 1 1075
0 140 7 2 2 137 1077
0 141 5 1 1 1079
0 142 7 1 2 1070 1080
0 143 5 2 1 142
0 144 7 1 2 131 141
0 145 5 1 1 144
0 146 7 2 2 1081 145
0 147 5 1 1 1083
0 148 7 2 2 105 1084
0 149 5 2 1 1085
0 150 7 1 2 1050 147
0 151 5 1 1 150
0 152 7 2 2 1087 151
0 153 5 1 1 1089
0 154 7 2 2 1046 1090
0 155 5 2 1 1091
0 156 7 1 2 1048 153
0 157 5 1 1 156
3 1788 7 0 2 1093 157
0 159 7 2 2 1068 1082
0 160 5 1 1 1095
0 161 7 2 2 21 968
0 162 5 1 1 1097
0 163 7 2 2 28 961
0 164 5 1 1 1099
0 165 7 2 2 103 954
0 166 5 1 1 1101
0 167 7 1 2 164 166
0 168 5 1 1 167
0 169 7 1 2 1100 1102
0 170 5 2 1 169
0 171 7 2 2 168 1103
0 172 5 1 1 1105
0 173 7 1 2 1098 1106
0 174 5 2 1 173
0 175 7 1 2 162 172
0 176 5 1 1 175
0 177 7 2 2 1107 176
0 178 5 1 1 1109
0 179 7 2 2 1060 1064
0 180 5 1 1 1111
0 181 7 2 2 712 947
0 182 5 1 1 1113
0 183 7 2 2 897 940
0 184 5 1 1 1115
0 185 7 2 2 904 933
0 186 5 1 1 1117
0 187 7 1 2 184 186
0 188 5 1 1 187
0 189 7 1 2 1116 1118
0 190 5 2 1 189
0 191 7 2 2 188 1119
0 192 5 1 1 1121
0 193 7 1 2 1114 1122
0 194 5 2 1 193
0 195 7 1 2 182 192
0 196 5 1 1 195
0 197 7 2 2 1123 196
0 198 5 1 1 1125
0 199 7 1 2 180 1126
0 200 5 2 1 199
0 201 7 1 2 1112 198
0 202 5 1 1 201
0 203 7 2 2 1127 202
0 204 5 1 1 1129
0 205 7 1 2 1110 1130
0 206 5 2 1 205
0 207 7 1 2 178 204
0 208 5 1 1 207
0 209 7 2 2 1131 208
0 210 5 1 1 1133
0 211 7 1 2 160 1134
0 212 5 2 1 211
0 213 7 1 2 1096 210
0 214 5 1 1 213
0 215 7 2 2 1135 214
0 216 5 1 1 1137
0 217 7 1 2 1076 1138
0 218 5 2 1 217
0 219 7 1 2 1078 216
0 220 5 1 1 219
0 221 7 4 2 1139 220
0 222 5 1 1 1141
0 223 7 2 2 1088 1094
0 224 5 1 1 1145
0 225 7 1 2 1142 1146
0 226 5 1 1 225
0 227 7 1 2 222 224
0 228 5 1 1 227
0 229 7 1 2 226 228
3 1789 5 0 1 229
0 231 7 2 2 1086 1143
0 232 5 1 1 1147
0 233 7 2 2 1136 1140
0 234 5 1 1 1149
0 235 7 2 2 22 976
0 236 5 1 1 1151
0 237 7 2 2 1104 1108
0 238 5 1 1 1153
0 239 7 2 2 1152 238
0 240 5 2 1 1155
0 241 7 1 2 236 1154
0 242 5 1 1 241
0 243 7 2 2 1157 242
0 244 5 1 1 1159
0 245 7 2 2 1128 1132
0 246 5 1 1 1161
0 247 7 2 2 29 969
0 248 5 1 1 1163
0 249 7 2 2 158 962
0 250 5 1 1 1165
0 251 7 2 2 777 955
0 252 5 1 1 1167
0 253 7 1 2 250 252
0 254 5 1 1 253
0 255 7 1 2 1166 1168
0 256 5 2 1 255
0 257 7 2 2 254 1169
0 258 5 1 1 1171
0 259 7 1 2 1164 1172
0 260 5 2 1 259
0 261 7 1 2 248 258
0 262 5 1 1 261
0 263 7 2 2 1173 262
0 264 5 1 1 1175
0 265 7 2 2 1120 1124
0 266 5 1 1 1177
0 267 7 2 2 898 948
0 268 5 1 1 1179
0 269 7 2 2 905 941
0 270 5 1 1 1181
0 271 7 2 2 912 934
0 272 5 1 1 1183
0 273 7 1 2 270 272
0 274 5 1 1 273
0 275 7 1 2 1182 1184
0 276 5 2 1 275
0 277 7 2 2 274 1185
0 278 5 1 1 1187
0 279 7 1 2 1180 1188
0 280 5 2 1 279
0 281 7 1 2 268 278
0 282 5 1 1 281
0 283 7 2 2 1189 282
0 284 5 1 1 1191
0 285 7 1 2 266 1192
0 286 5 2 1 285
0 287 7 1 2 1178 284
0 288 5 1 1 287
0 289 7 2 2 1193 288
0 290 5 1 1 1195
0 291 7 1 2 1176 1196
0 292 5 2 1 291
0 293 7 1 2 264 290
0 294 5 1 1 293
0 295 7 2 2 1197 294
0 296 5 1 1 1199
0 297 7 1 2 246 1200
0 298 5 2 1 297
0 299 7 1 2 1162 296
0 300 5 1 1 299
0 301 7 2 2 1201 300
0 302 5 1 1 1203
0 303 7 1 2 1160 1204
0 304 5 2 1 303
0 305 7 1 2 244 302
0 306 5 1 1 305
0 307 7 2 2 1205 306
0 308 5 1 1 1207
0 309 7 2 2 234 1208
0 310 5 2 1 1209
0 311 7 1 2 1150 308
0 312 5 1 1 311
0 313 7 2 2 1211 312
0 314 5 1 1 1213
0 315 7 1 2 1148 1214
0 316 5 2 1 315
0 317 7 1 2 232 314
0 318 5 1 1 317
0 319 7 2 2 1215 318
0 320 5 1 1 1217
0 321 7 2 2 1092 1144
0 322 5 1 1 1219
0 323 7 1 2 1218 1220
0 324 5 2 1 323
0 325 7 1 2 320 322
0 326 5 1 1 325
3 1790 7 0 2 1221 326
0 328 7 2 2 1216 1222
0 329 5 1 1 1223
0 330 7 2 2 1202 1206
0 331 5 1 1 1225
0 332 7 2 2 23 985
0 333 5 1 1 1227
0 334 7 2 2 1170 1174
0 335 5 1 1 1229
0 336 7 2 2 30 977
0 337 5 1 1 1231
0 338 7 1 2 335 1232
0 339 5 2 1 338
0 340 7 1 2 1230 337
0 341 5 1 1 340
0 342 7 2 2 1233 341
0 343 5 1 1 1235
0 344 7 1 2 1228 1236
0 345 5 2 1 344
0 346 7 1 2 333 343
0 347 5 1 1 346
0 348 7 2 2 1237 347
0 349 5 1 1 1239
0 350 7 2 2 1194 1198
0 351 5 1 1 1241
0 352 7 2 2 230 970
0 353 5 1 1 1243
0 354 7 2 2 830 963
0 355 5 1 1 1245
0 356 7 2 2 899 956
0 357 5 1 1 1247
0 358 7 1 2 355 357
0 359 5 1 1 358
0 360 7 1 2 1246 1248
0 361 5 2 1 360
0 362 7 2 2 359 1249
0 363 5 1 1 1251
0 364 7 1 2 1244 1252
0 365 5 2 1 364
0 366 7 1 2 353 363
0 367 5 1 1 366
0 368 7 2 2 1253 367
0 369 5 1 1 1255
0 370 7 2 2 1186 1190
0 371 5 1 1 1257
0 372 7 2 2 906 949
0 373 5 1 1 1259
0 374 7 2 2 913 942
0 375 5 2 1 1261
0 376 7 2 2 920 935
0 377 5 1 1 1265
0 378 7 1 2 1263 377
0 379 5 1 1 378
0 380 7 1 2 1262 1266
0 381 5 2 1 380
0 382 7 2 2 379 1267
0 383 5 1 1 1269
0 384 7 1 2 1260 1270
0 385 5 2 1 384
0 386 7 1 2 373 383
0 387 5 1 1 386
0 388 7 2 2 1271 387
0 389 5 1 1 1273
0 390 7 1 2 371 1274
0 391 5 2 1 390
0 392 7 1 2 1258 389
0 393 5 1 1 392
0 394 7 2 2 1275 393
0 395 5 1 1 1277
0 396 7 1 2 1256 1278
0 397 5 2 1 396
0 398 7 1 2 369 395
0 399 5 1 1 398
0 400 7 2 2 1279 399
0 401 5 1 1 1281
0 402 7 1 2 351 1282
0 403 5 2 1 402
0 404 7 1 2 1242 401
0 405 5 1 1 404
0 406 7 2 2 1283 405
0 407 5 1 1 1285
0 408 7 1 2 1240 1286
0 409 5 2 1 408
0 410 7 1 2 349 407
0 411 5 1 1 410
0 412 7 2 2 1287 411
0 413 5 1 1 1289
0 414 7 1 2 331 1290
0 415 5 2 1 414
0 416 7 1 2 1226 413
0 417 5 1 1 416
0 418 7 2 2 1291 417
0 419 5 1 1 1293
0 420 7 1 2 1156 1294
0 421 5 2 1 420
0 422 7 1 2 1158 419
0 423 5 1 1 422
0 424 7 2 2 1295 423
0 425 5 1 1 1297
0 426 7 1 2 1210 1298
0 427 5 2 1 426
0 428 7 1 2 1212 425
0 429 5 1 1 428
0 430 7 2 2 1299 429
0 431 5 1 1 1301
0 432 7 1 2 329 1302
0 433 5 2 1 432
0 434 7 1 2 1224 431
0 435 5 1 1 434
3 1791 7 0 2 1303 435
0 437 7 2 2 1300 1304
0 438 5 1 1 1305
0 439 7 2 2 1292 1296
0 440 5 1 1 1307
0 441 7 2 2 1234 1238
0 442 5 1 1 1309
0 443 7 2 2 1284 1288
0 444 5 1 1 1311
0 445 7 2 2 31 986
0 446 5 1 1 1313
0 447 7 2 2 1250 1254
0 448 5 1 1 1315
0 449 7 2 2 327 978
0 450 5 1 1 1317
0 451 7 1 2 448 1318
0 452 5 2 1 451
0 453 7 1 2 1316 450
0 454 5 1 1 453
0 455 7 2 2 1319 454
0 456 5 1 1 1321
0 457 7 1 2 1314 1322
0 458 5 2 1 457
0 459 7 1 2 446 456
0 460 5 1 1 459
0 461 7 2 2 1323 460
0 462 5 1 1 1325
0 463 7 2 2 1276 1280
0 464 5 1 1 1327
0 465 7 2 2 869 971
0 466 5 1 1 1329
0 467 7 2 2 900 964
0 468 5 1 1 1331
0 469 7 2 2 907 957
0 470 5 1 1 1333
0 471 7 1 2 468 470
0 472 5 1 1 471
0 473 7 1 2 1332 1334
0 474 5 2 1 473
0 475 7 2 2 472 1335
0 476 5 1 1 1337
0 477 7 1 2 1330 1338
0 478 5 2 1 477
0 479 7 1 2 466 476
0 480 5 1 1 479
0 481 7 2 2 1339 480
0 482 5 1 1 1341
0 483 7 2 2 1268 1272
0 484 5 1 1 1343
0 485 7 2 2 921 943
0 486 5 1 1 1345
0 487 7 2 2 914 950
0 488 5 1 1 1347
0 489 7 1 2 486 488
0 490 5 1 1 489
0 491 7 1 2 1346 1348
0 492 5 2 1 491
0 493 7 2 2 490 1349
0 494 5 1 1 1351
0 495 7 1 2 484 1352
0 496 5 2 1 495
0 497 7 1 2 1344 494
0 498 5 1 1 497
0 499 7 2 2 1353 498
0 500 5 1 1 1355
0 501 7 1 2 1342 1356
0 502 5 2 1 501
0 503 7 1 2 482 500
0 504 5 1 1 503
0 505 7 2 2 1357 504
0 506 5 1 1 1359
0 507 7 1 2 464 1360
0 508 5 2 1 507
0 509 7 1 2 1328 506
0 510 5 1 1 509
0 511 7 2 2 1361 510
0 512 5 1 1 1363
0 513 7 1 2 1326 1364
0 514 5 2 1 513
0 515 7 1 2 462 512
0 516 5 1 1 515
0 517 7 2 2 1365 516
0 518 5 1 1 1367
0 519 7 1 2 444 1368
0 520 5 2 1 519
0 521 7 1 2 1312 518
0 522 5 1 1 521
0 523 7 2 2 1369 522
0 524 5 1 1 1371
0 525 7 1 2 442 1372
0 526 5 2 1 525
0 527 7 1 2 1310 524
0 528 5 1 1 527
0 529 7 2 2 1373 528
0 530 5 1 1 1375
0 531 7 1 2 440 1376
0 532 5 2 1 531
0 533 7 1 2 1308 530
0 534 5 1 1 533
0 535 7 2 2 1377 534
0 536 5 1 1 1379
0 537 7 1 2 438 1380
0 538 5 2 1 537
0 539 7 1 2 1306 536
0 540 5 1 1 539
3 1792 7 0 2 1381 540
0 542 7 2 2 1378 1382
0 543 5 1 1 1383
0 544 7 2 2 1370 1374
0 545 5 1 1 1385
0 546 7 2 2 1320 1324
0 547 5 1 1 1387
0 548 7 2 2 1362 1366
0 549 5 1 1 1389
0 550 7 2 2 436 987
0 551 5 1 1 1391
0 552 7 2 2 1336 1340
0 553 5 1 1 1393
0 554 7 2 2 887 979
0 555 5 1 1 1395
0 556 7 1 2 553 1396
0 557 5 2 1 556
0 558 7 1 2 1394 555
0 559 5 1 1 558
0 560 7 2 2 1397 559
0 561 5 1 1 1399
0 562 7 1 2 1392 1400
0 563 5 2 1 562
0 564 7 1 2 551 561
0 565 5 1 1 564
0 566 7 2 2 1401 565
0 567 5 1 1 1403
0 568 7 2 2 1354 1358
0 569 5 1 1 1405
0 570 7 2 2 901 972
0 571 5 1 1 1407
0 572 7 2 2 908 965
0 573 5 1 1 1409
0 574 7 2 2 915 958
0 575 5 1 1 1411
0 576 7 1 2 573 575
0 577 5 1 1 576
0 578 7 1 2 1410 1412
0 579 5 2 1 578
0 580 7 2 2 577 1413
0 581 5 1 1 1415
0 582 7 1 2 1408 1416
0 583 5 2 1 582
0 584 7 1 2 571 581
0 585 5 1 1 584
0 586 7 2 2 1417 585
0 587 5 1 1 1419
0 588 7 1 2 922 951
0 589 7 2 2 1264 588
0 590 5 1 1 1421
0 591 7 1 2 1420 1422
0 592 5 2 1 591
0 593 7 1 2 587 590
0 594 5 1 1 593
0 595 7 2 2 1423 594
0 596 5 1 1 1425
0 597 7 1 2 569 1426
0 598 5 2 1 597
0 599 7 1 2 1406 596
0 600 5 1 1 599
0 601 7 2 2 1427 600
0 602 5 1 1 1429
0 603 7 1 2 1404 1430
0 604 5 2 1 603
0 605 7 1 2 567 602
0 606 5 1 1 605
0 607 7 2 2 1431 606
0 608 5 1 1 1433
0 609 7 1 2 549 1434
0 610 5 2 1 609
0 611 7 1 2 1390 608
0 612 5 1 1 611
0 613 7 2 2 1435 612
0 614 5 1 1 1437
0 615 7 1 2 547 1438
0 616 5 2 1 615
0 617 7 1 2 1388 614
0 618 5 1 1 617
0 619 7 2 2 1439 618
0 620 5 1 1 1441
0 621 7 1 2 545 1442
0 622 5 2 1 621
0 623 7 1 2 1386 620
0 624 5 1 1 623
0 625 7 2 2 1443 624
0 626 5 1 1 1445
0 627 7 1 2 543 1446
0 628 5 2 1 627
0 629 7 1 2 1384 626
0 630 5 1 1 629
3 1793 7 0 2 1447 630
0 632 7 2 2 1444 1448
0 633 5 1 1 1449
0 634 7 2 2 1436 1440
0 635 5 1 1 1451
0 636 7 2 2 1398 1402
0 637 5 1 1 1453
0 638 7 2 2 1428 1432
0 639 5 1 1 1455
0 640 7 2 2 895 988
0 641 5 1 1 1457
0 642 7 2 2 1414 1418
0 643 5 1 1 1459
0 644 7 2 2 902 980
0 645 5 1 1 1461
0 646 7 1 2 643 1462
0 647 5 2 1 646
0 648 7 1 2 1460 645
0 649 5 1 1 648
0 650 7 2 2 1463 649
0 651 5 1 1 1465
0 652 7 1 2 1458 1466
0 653 5 2 1 652
0 654 7 1 2 641 651
0 655 5 1 1 654
0 656 7 2 2 1467 655
0 657 5 1 1 1469
0 658 7 2 2 1350 1424
0 659 5 1 1 1471
0 660 7 2 2 909 973
0 661 5 1 1 1473
0 662 7 2 2 916 966
0 663 5 1 1 1475
0 664 7 2 2 923 959
0 665 5 1 1 1477
0 666 7 1 2 663 665
0 667 5 1 1 666
0 668 7 1 2 1476 1478
0 669 5 2 1 668
0 670 7 2 2 667 1479
0 671 5 1 1 1481
0 672 7 1 2 1474 1482
0 673 5 2 1 672
0 674 7 1 2 661 671
0 675 5 1 1 674
0 676 7 2 2 1483 675
0 677 5 1 1 1485
0 678 7 1 2 659 1486
0 679 5 2 1 678
0 680 7 1 2 1472 677
0 681 5 1 1 680
0 682 7 2 2 1487 681
0 683 5 1 1 1489
0 684 7 1 2 1470 1490
0 685 5 2 1 684
0 686 7 1 2 657 683
0 687 5 1 1 686
0 688 7 2 2 1491 687
0 689 5 1 1 1493
0 690 7 1 2 639 1494
0 691 5 2 1 690
0 692 7 1 2 1456 689
0 693 5 1 1 692
0 694 7 2 2 1495 693
0 695 5 1 1 1497
0 696 7 1 2 637 1498
0 697 5 2 1 696
0 698 7 1 2 1454 695
0 699 5 1 1 698
0 700 7 2 2 1499 699
0 701 5 1 1 1501
0 702 7 1 2 635 1502
0 703 5 2 1 702
0 704 7 1 2 1452 701
0 705 5 1 1 704
0 706 7 2 2 1503 705
0 707 5 1 1 1505
0 708 7 1 2 633 1506
0 709 5 2 1 708
0 710 7 1 2 1450 707
0 711 5 1 1 710
3 1794 7 0 2 1507 711
0 713 7 2 2 1504 1508
0 714 5 1 1 1509
0 715 7 2 2 1496 1500
0 716 5 1 1 1511
0 717 7 2 2 1464 1468
0 718 5 1 1 1513
0 719 7 2 2 1488 1492
0 720 5 1 1 1515
0 721 7 2 2 903 989
0 722 5 1 1 1517
0 723 7 2 2 1480 1484
0 724 5 1 1 1519
0 725 7 2 2 910 981
0 726 5 1 1 1521
0 727 7 1 2 724 1522
0 728 5 2 1 727
0 729 7 1 2 1520 726
0 730 5 1 1 729
0 731 7 2 2 1523 730
0 732 5 1 1 1525
0 733 7 1 2 1518 1526
0 734 5 2 1 733
0 735 7 1 2 722 732
0 736 5 1 1 735
0 737 7 2 2 1527 736
0 738 5 1 1 1529
0 739 7 2 2 924 967
0 740 5 1 1 1531
0 741 7 2 2 917 974
0 742 5 1 1 1533
0 743 7 1 2 740 742
0 744 5 1 1 743
0 745 7 2 2 1532 1534
0 746 5 2 1 1535
0 747 7 2 2 744 1537
0 748 5 1 1 1539
0 749 7 2 2 1530 1540
0 750 5 2 1 1541
0 751 7 1 2 738 748
0 752 5 1 1 751
0 753 7 2 2 1543 752
0 754 5 1 1 1545
0 755 7 1 2 720 1546
0 756 5 2 1 755
0 757 7 1 2 1516 754
0 758 5 1 1 757
0 759 7 2 2 1547 758
0 760 5 1 1 1549
0 761 7 1 2 718 1550
0 762 5 2 1 761
0 763 7 1 2 1514 760
0 764 5 1 1 763
0 765 7 2 2 1551 764
0 766 5 1 1 1553
0 767 7 1 2 716 1554
0 768 5 2 1 767
0 769 7 1 2 1512 766
0 770 5 1 1 769
0 771 7 2 2 1555 770
0 772 5 1 1 1557
0 773 7 1 2 714 1558
0 774 5 2 1 773
0 775 7 1 2 1510 772
0 776 5 1 1 775
3 1795 7 0 2 1559 776
0 778 7 2 2 1556 1560
0 779 5 1 1 1561
0 780 7 2 2 1548 1552
0 781 5 1 1 1563
0 782 7 2 2 1524 1528
0 783 5 1 1 1565
0 784 7 2 2 925 975
0 785 5 1 1 1567
0 786 7 2 2 911 990
0 787 5 1 1 1569
0 788 7 1 2 918 982
0 789 5 2 1 788
0 790 7 1 2 1538 1571
0 791 5 1 1 790
0 792 7 1 2 983 1536
0 793 5 2 1 792
0 794 7 2 2 791 1573
0 795 5 1 1 1575
0 796 7 1 2 1570 1576
0 797 5 2 1 796
0 798 7 1 2 787 795
0 799 5 1 1 798
0 800 7 2 2 1577 799
0 801 5 1 1 1579
0 802 7 2 2 1568 1580
0 803 5 2 1 1581
0 804 7 1 2 785 801
0 805 5 1 1 804
0 806 7 2 2 1583 805
0 807 5 1 1 1585
0 808 7 1 2 1542 1586
0 809 5 2 1 808
0 810 7 1 2 1544 807
0 811 5 1 1 810
0 812 7 2 2 1587 811
0 813 5 1 1 1589
0 814 7 1 2 783 1590
0 815 5 2 1 814
0 816 7 1 2 1566 813
0 817 5 1 1 816
0 818 7 2 2 1591 817
0 819 5 1 1 1593
0 820 7 1 2 781 1594
0 821 5 2 1 820
0 822 7 1 2 1564 819
0 823 5 1 1 822
0 824 7 2 2 1595 823
0 825 5 1 1 1597
0 826 7 1 2 779 1598
0 827 5 2 1 826
0 828 7 1 2 1562 825
0 829 5 1 1 828
3 1796 7 0 2 1599 829
0 831 7 2 2 1596 1600
0 832 5 1 1 1601
0 833 7 2 2 1588 1592
0 834 5 1 1 1603
0 835 7 2 2 1574 1578
0 836 5 1 1 1605
0 837 7 2 2 919 991
0 838 5 1 1 1607
0 839 7 2 2 926 984
0 840 5 1 1 1609
0 841 7 1 2 838 840
0 842 5 1 1 841
0 843 7 1 2 1608 1610
0 844 5 3 1 843
0 845 7 2 2 842 1611
0 846 5 1 1 1614
0 847 7 1 2 1582 1615
0 848 5 2 1 847
0 849 7 1 2 1584 846
0 850 5 1 1 849
0 851 7 2 2 1616 850
0 852 5 1 1 1618
0 853 7 1 2 836 1619
0 854 5 2 1 853
0 855 7 1 2 1606 852
0 856 5 1 1 855
0 857 7 2 2 1620 856
0 858 5 1 1 1622
0 859 7 1 2 834 1623
0 860 5 2 1 859
0 861 7 1 2 1604 858
0 862 5 1 1 861
0 863 7 2 2 1624 862
0 864 5 1 1 1626
0 865 7 1 2 832 1627
0 866 5 2 1 865
0 867 7 1 2 1602 864
0 868 5 1 1 867
3 1797 7 0 2 1628 868
0 870 7 2 2 1625 1629
0 871 5 1 1 1630
0 872 7 2 2 1617 1621
0 873 5 1 1 1632
0 874 7 1 2 927 992
0 875 7 2 2 1572 874
0 876 5 1 1 1634
0 877 7 1 2 873 1635
0 878 5 2 1 877
0 879 7 1 2 1633 876
0 880 5 1 1 879
0 881 7 2 2 1636 880
0 882 5 1 1 1638
0 883 7 2 2 871 1639
0 884 5 2 1 1640
0 885 7 1 2 1631 882
0 886 5 1 1 885
3 1798 7 0 2 1642 886
0 888 7 1 2 1612 1641
0 889 5 1 1 888
0 890 7 1 2 1613 1637
0 891 5 1 1 890
0 892 7 1 2 1643 891
0 893 5 1 1 892
0 894 7 1 2 889 893
3 1799 5 0 1 894
